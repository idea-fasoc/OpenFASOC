* NGSPICE file created from diff_pair_sample_0943.ext - technology: sky130A

.subckt diff_pair_sample_0943 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=0 ps=0 w=14.11 l=3.76
X1 VTAIL.t7 VN.t0 VDD2.t3 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=2.32815 ps=14.44 w=14.11 l=3.76
X2 VTAIL.t6 VN.t1 VDD2.t2 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=2.32815 ps=14.44 w=14.11 l=3.76
X3 VDD1.t3 VP.t0 VTAIL.t3 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=2.32815 pd=14.44 as=5.5029 ps=29 w=14.11 l=3.76
X4 B.t8 B.t6 B.t7 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=0 ps=0 w=14.11 l=3.76
X5 VTAIL.t0 VP.t1 VDD1.t2 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=2.32815 ps=14.44 w=14.11 l=3.76
X6 B.t5 B.t3 B.t4 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=0 ps=0 w=14.11 l=3.76
X7 VDD1.t1 VP.t2 VTAIL.t1 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=2.32815 pd=14.44 as=5.5029 ps=29 w=14.11 l=3.76
X8 VDD2.t0 VN.t2 VTAIL.t5 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=2.32815 pd=14.44 as=5.5029 ps=29 w=14.11 l=3.76
X9 B.t2 B.t0 B.t1 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=0 ps=0 w=14.11 l=3.76
X10 VTAIL.t2 VP.t3 VDD1.t0 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=5.5029 pd=29 as=2.32815 ps=14.44 w=14.11 l=3.76
X11 VDD2.t1 VN.t3 VTAIL.t4 w_n3424_n3790# sky130_fd_pr__pfet_01v8 ad=2.32815 pd=14.44 as=5.5029 ps=29 w=14.11 l=3.76
R0 B.n562 B.n561 585
R1 B.n563 B.n80 585
R2 B.n565 B.n564 585
R3 B.n566 B.n79 585
R4 B.n568 B.n567 585
R5 B.n569 B.n78 585
R6 B.n571 B.n570 585
R7 B.n572 B.n77 585
R8 B.n574 B.n573 585
R9 B.n575 B.n76 585
R10 B.n577 B.n576 585
R11 B.n578 B.n75 585
R12 B.n580 B.n579 585
R13 B.n581 B.n74 585
R14 B.n583 B.n582 585
R15 B.n584 B.n73 585
R16 B.n586 B.n585 585
R17 B.n587 B.n72 585
R18 B.n589 B.n588 585
R19 B.n590 B.n71 585
R20 B.n592 B.n591 585
R21 B.n593 B.n70 585
R22 B.n595 B.n594 585
R23 B.n596 B.n69 585
R24 B.n598 B.n597 585
R25 B.n599 B.n68 585
R26 B.n601 B.n600 585
R27 B.n602 B.n67 585
R28 B.n604 B.n603 585
R29 B.n605 B.n66 585
R30 B.n607 B.n606 585
R31 B.n608 B.n65 585
R32 B.n610 B.n609 585
R33 B.n611 B.n64 585
R34 B.n613 B.n612 585
R35 B.n614 B.n63 585
R36 B.n616 B.n615 585
R37 B.n617 B.n62 585
R38 B.n619 B.n618 585
R39 B.n620 B.n61 585
R40 B.n622 B.n621 585
R41 B.n623 B.n60 585
R42 B.n625 B.n624 585
R43 B.n626 B.n59 585
R44 B.n628 B.n627 585
R45 B.n629 B.n58 585
R46 B.n631 B.n630 585
R47 B.n632 B.n55 585
R48 B.n635 B.n634 585
R49 B.n636 B.n54 585
R50 B.n638 B.n637 585
R51 B.n639 B.n53 585
R52 B.n641 B.n640 585
R53 B.n642 B.n52 585
R54 B.n644 B.n643 585
R55 B.n645 B.n51 585
R56 B.n647 B.n646 585
R57 B.n649 B.n648 585
R58 B.n650 B.n47 585
R59 B.n652 B.n651 585
R60 B.n653 B.n46 585
R61 B.n655 B.n654 585
R62 B.n656 B.n45 585
R63 B.n658 B.n657 585
R64 B.n659 B.n44 585
R65 B.n661 B.n660 585
R66 B.n662 B.n43 585
R67 B.n664 B.n663 585
R68 B.n665 B.n42 585
R69 B.n667 B.n666 585
R70 B.n668 B.n41 585
R71 B.n670 B.n669 585
R72 B.n671 B.n40 585
R73 B.n673 B.n672 585
R74 B.n674 B.n39 585
R75 B.n676 B.n675 585
R76 B.n677 B.n38 585
R77 B.n679 B.n678 585
R78 B.n680 B.n37 585
R79 B.n682 B.n681 585
R80 B.n683 B.n36 585
R81 B.n685 B.n684 585
R82 B.n686 B.n35 585
R83 B.n688 B.n687 585
R84 B.n689 B.n34 585
R85 B.n691 B.n690 585
R86 B.n692 B.n33 585
R87 B.n694 B.n693 585
R88 B.n695 B.n32 585
R89 B.n697 B.n696 585
R90 B.n698 B.n31 585
R91 B.n700 B.n699 585
R92 B.n701 B.n30 585
R93 B.n703 B.n702 585
R94 B.n704 B.n29 585
R95 B.n706 B.n705 585
R96 B.n707 B.n28 585
R97 B.n709 B.n708 585
R98 B.n710 B.n27 585
R99 B.n712 B.n711 585
R100 B.n713 B.n26 585
R101 B.n715 B.n714 585
R102 B.n716 B.n25 585
R103 B.n718 B.n717 585
R104 B.n719 B.n24 585
R105 B.n560 B.n81 585
R106 B.n559 B.n558 585
R107 B.n557 B.n82 585
R108 B.n556 B.n555 585
R109 B.n554 B.n83 585
R110 B.n553 B.n552 585
R111 B.n551 B.n84 585
R112 B.n550 B.n549 585
R113 B.n548 B.n85 585
R114 B.n547 B.n546 585
R115 B.n545 B.n86 585
R116 B.n544 B.n543 585
R117 B.n542 B.n87 585
R118 B.n541 B.n540 585
R119 B.n539 B.n88 585
R120 B.n538 B.n537 585
R121 B.n536 B.n89 585
R122 B.n535 B.n534 585
R123 B.n533 B.n90 585
R124 B.n532 B.n531 585
R125 B.n530 B.n91 585
R126 B.n529 B.n528 585
R127 B.n527 B.n92 585
R128 B.n526 B.n525 585
R129 B.n524 B.n93 585
R130 B.n523 B.n522 585
R131 B.n521 B.n94 585
R132 B.n520 B.n519 585
R133 B.n518 B.n95 585
R134 B.n517 B.n516 585
R135 B.n515 B.n96 585
R136 B.n514 B.n513 585
R137 B.n512 B.n97 585
R138 B.n511 B.n510 585
R139 B.n509 B.n98 585
R140 B.n508 B.n507 585
R141 B.n506 B.n99 585
R142 B.n505 B.n504 585
R143 B.n503 B.n100 585
R144 B.n502 B.n501 585
R145 B.n500 B.n101 585
R146 B.n499 B.n498 585
R147 B.n497 B.n102 585
R148 B.n496 B.n495 585
R149 B.n494 B.n103 585
R150 B.n493 B.n492 585
R151 B.n491 B.n104 585
R152 B.n490 B.n489 585
R153 B.n488 B.n105 585
R154 B.n487 B.n486 585
R155 B.n485 B.n106 585
R156 B.n484 B.n483 585
R157 B.n482 B.n107 585
R158 B.n481 B.n480 585
R159 B.n479 B.n108 585
R160 B.n478 B.n477 585
R161 B.n476 B.n109 585
R162 B.n475 B.n474 585
R163 B.n473 B.n110 585
R164 B.n472 B.n471 585
R165 B.n470 B.n111 585
R166 B.n469 B.n468 585
R167 B.n467 B.n112 585
R168 B.n466 B.n465 585
R169 B.n464 B.n113 585
R170 B.n463 B.n462 585
R171 B.n461 B.n114 585
R172 B.n460 B.n459 585
R173 B.n458 B.n115 585
R174 B.n457 B.n456 585
R175 B.n455 B.n116 585
R176 B.n454 B.n453 585
R177 B.n452 B.n117 585
R178 B.n451 B.n450 585
R179 B.n449 B.n118 585
R180 B.n448 B.n447 585
R181 B.n446 B.n119 585
R182 B.n445 B.n444 585
R183 B.n443 B.n120 585
R184 B.n442 B.n441 585
R185 B.n440 B.n121 585
R186 B.n439 B.n438 585
R187 B.n437 B.n122 585
R188 B.n436 B.n435 585
R189 B.n434 B.n123 585
R190 B.n433 B.n432 585
R191 B.n431 B.n124 585
R192 B.n430 B.n429 585
R193 B.n428 B.n125 585
R194 B.n269 B.n182 585
R195 B.n271 B.n270 585
R196 B.n272 B.n181 585
R197 B.n274 B.n273 585
R198 B.n275 B.n180 585
R199 B.n277 B.n276 585
R200 B.n278 B.n179 585
R201 B.n280 B.n279 585
R202 B.n281 B.n178 585
R203 B.n283 B.n282 585
R204 B.n284 B.n177 585
R205 B.n286 B.n285 585
R206 B.n287 B.n176 585
R207 B.n289 B.n288 585
R208 B.n290 B.n175 585
R209 B.n292 B.n291 585
R210 B.n293 B.n174 585
R211 B.n295 B.n294 585
R212 B.n296 B.n173 585
R213 B.n298 B.n297 585
R214 B.n299 B.n172 585
R215 B.n301 B.n300 585
R216 B.n302 B.n171 585
R217 B.n304 B.n303 585
R218 B.n305 B.n170 585
R219 B.n307 B.n306 585
R220 B.n308 B.n169 585
R221 B.n310 B.n309 585
R222 B.n311 B.n168 585
R223 B.n313 B.n312 585
R224 B.n314 B.n167 585
R225 B.n316 B.n315 585
R226 B.n317 B.n166 585
R227 B.n319 B.n318 585
R228 B.n320 B.n165 585
R229 B.n322 B.n321 585
R230 B.n323 B.n164 585
R231 B.n325 B.n324 585
R232 B.n326 B.n163 585
R233 B.n328 B.n327 585
R234 B.n329 B.n162 585
R235 B.n331 B.n330 585
R236 B.n332 B.n161 585
R237 B.n334 B.n333 585
R238 B.n335 B.n160 585
R239 B.n337 B.n336 585
R240 B.n338 B.n159 585
R241 B.n340 B.n339 585
R242 B.n342 B.n341 585
R243 B.n343 B.n155 585
R244 B.n345 B.n344 585
R245 B.n346 B.n154 585
R246 B.n348 B.n347 585
R247 B.n349 B.n153 585
R248 B.n351 B.n350 585
R249 B.n352 B.n152 585
R250 B.n354 B.n353 585
R251 B.n356 B.n149 585
R252 B.n358 B.n357 585
R253 B.n359 B.n148 585
R254 B.n361 B.n360 585
R255 B.n362 B.n147 585
R256 B.n364 B.n363 585
R257 B.n365 B.n146 585
R258 B.n367 B.n366 585
R259 B.n368 B.n145 585
R260 B.n370 B.n369 585
R261 B.n371 B.n144 585
R262 B.n373 B.n372 585
R263 B.n374 B.n143 585
R264 B.n376 B.n375 585
R265 B.n377 B.n142 585
R266 B.n379 B.n378 585
R267 B.n380 B.n141 585
R268 B.n382 B.n381 585
R269 B.n383 B.n140 585
R270 B.n385 B.n384 585
R271 B.n386 B.n139 585
R272 B.n388 B.n387 585
R273 B.n389 B.n138 585
R274 B.n391 B.n390 585
R275 B.n392 B.n137 585
R276 B.n394 B.n393 585
R277 B.n395 B.n136 585
R278 B.n397 B.n396 585
R279 B.n398 B.n135 585
R280 B.n400 B.n399 585
R281 B.n401 B.n134 585
R282 B.n403 B.n402 585
R283 B.n404 B.n133 585
R284 B.n406 B.n405 585
R285 B.n407 B.n132 585
R286 B.n409 B.n408 585
R287 B.n410 B.n131 585
R288 B.n412 B.n411 585
R289 B.n413 B.n130 585
R290 B.n415 B.n414 585
R291 B.n416 B.n129 585
R292 B.n418 B.n417 585
R293 B.n419 B.n128 585
R294 B.n421 B.n420 585
R295 B.n422 B.n127 585
R296 B.n424 B.n423 585
R297 B.n425 B.n126 585
R298 B.n427 B.n426 585
R299 B.n268 B.n267 585
R300 B.n266 B.n183 585
R301 B.n265 B.n264 585
R302 B.n263 B.n184 585
R303 B.n262 B.n261 585
R304 B.n260 B.n185 585
R305 B.n259 B.n258 585
R306 B.n257 B.n186 585
R307 B.n256 B.n255 585
R308 B.n254 B.n187 585
R309 B.n253 B.n252 585
R310 B.n251 B.n188 585
R311 B.n250 B.n249 585
R312 B.n248 B.n189 585
R313 B.n247 B.n246 585
R314 B.n245 B.n190 585
R315 B.n244 B.n243 585
R316 B.n242 B.n191 585
R317 B.n241 B.n240 585
R318 B.n239 B.n192 585
R319 B.n238 B.n237 585
R320 B.n236 B.n193 585
R321 B.n235 B.n234 585
R322 B.n233 B.n194 585
R323 B.n232 B.n231 585
R324 B.n230 B.n195 585
R325 B.n229 B.n228 585
R326 B.n227 B.n196 585
R327 B.n226 B.n225 585
R328 B.n224 B.n197 585
R329 B.n223 B.n222 585
R330 B.n221 B.n198 585
R331 B.n220 B.n219 585
R332 B.n218 B.n199 585
R333 B.n217 B.n216 585
R334 B.n215 B.n200 585
R335 B.n214 B.n213 585
R336 B.n212 B.n201 585
R337 B.n211 B.n210 585
R338 B.n209 B.n202 585
R339 B.n208 B.n207 585
R340 B.n206 B.n203 585
R341 B.n205 B.n204 585
R342 B.n2 B.n0 585
R343 B.n785 B.n1 585
R344 B.n784 B.n783 585
R345 B.n782 B.n3 585
R346 B.n781 B.n780 585
R347 B.n779 B.n4 585
R348 B.n778 B.n777 585
R349 B.n776 B.n5 585
R350 B.n775 B.n774 585
R351 B.n773 B.n6 585
R352 B.n772 B.n771 585
R353 B.n770 B.n7 585
R354 B.n769 B.n768 585
R355 B.n767 B.n8 585
R356 B.n766 B.n765 585
R357 B.n764 B.n9 585
R358 B.n763 B.n762 585
R359 B.n761 B.n10 585
R360 B.n760 B.n759 585
R361 B.n758 B.n11 585
R362 B.n757 B.n756 585
R363 B.n755 B.n12 585
R364 B.n754 B.n753 585
R365 B.n752 B.n13 585
R366 B.n751 B.n750 585
R367 B.n749 B.n14 585
R368 B.n748 B.n747 585
R369 B.n746 B.n15 585
R370 B.n745 B.n744 585
R371 B.n743 B.n16 585
R372 B.n742 B.n741 585
R373 B.n740 B.n17 585
R374 B.n739 B.n738 585
R375 B.n737 B.n18 585
R376 B.n736 B.n735 585
R377 B.n734 B.n19 585
R378 B.n733 B.n732 585
R379 B.n731 B.n20 585
R380 B.n730 B.n729 585
R381 B.n728 B.n21 585
R382 B.n727 B.n726 585
R383 B.n725 B.n22 585
R384 B.n724 B.n723 585
R385 B.n722 B.n23 585
R386 B.n721 B.n720 585
R387 B.n787 B.n786 585
R388 B.n269 B.n268 550.159
R389 B.n720 B.n719 550.159
R390 B.n426 B.n125 550.159
R391 B.n562 B.n81 550.159
R392 B.n150 B.t11 492.95
R393 B.n56 B.t4 492.95
R394 B.n156 B.t2 492.95
R395 B.n48 B.t7 492.95
R396 B.n151 B.t10 413.63
R397 B.n57 B.t5 413.63
R398 B.n157 B.t1 413.63
R399 B.n49 B.t8 413.63
R400 B.n150 B.t9 299.752
R401 B.n156 B.t0 299.752
R402 B.n48 B.t6 299.752
R403 B.n56 B.t3 299.752
R404 B.n268 B.n183 163.367
R405 B.n264 B.n183 163.367
R406 B.n264 B.n263 163.367
R407 B.n263 B.n262 163.367
R408 B.n262 B.n185 163.367
R409 B.n258 B.n185 163.367
R410 B.n258 B.n257 163.367
R411 B.n257 B.n256 163.367
R412 B.n256 B.n187 163.367
R413 B.n252 B.n187 163.367
R414 B.n252 B.n251 163.367
R415 B.n251 B.n250 163.367
R416 B.n250 B.n189 163.367
R417 B.n246 B.n189 163.367
R418 B.n246 B.n245 163.367
R419 B.n245 B.n244 163.367
R420 B.n244 B.n191 163.367
R421 B.n240 B.n191 163.367
R422 B.n240 B.n239 163.367
R423 B.n239 B.n238 163.367
R424 B.n238 B.n193 163.367
R425 B.n234 B.n193 163.367
R426 B.n234 B.n233 163.367
R427 B.n233 B.n232 163.367
R428 B.n232 B.n195 163.367
R429 B.n228 B.n195 163.367
R430 B.n228 B.n227 163.367
R431 B.n227 B.n226 163.367
R432 B.n226 B.n197 163.367
R433 B.n222 B.n197 163.367
R434 B.n222 B.n221 163.367
R435 B.n221 B.n220 163.367
R436 B.n220 B.n199 163.367
R437 B.n216 B.n199 163.367
R438 B.n216 B.n215 163.367
R439 B.n215 B.n214 163.367
R440 B.n214 B.n201 163.367
R441 B.n210 B.n201 163.367
R442 B.n210 B.n209 163.367
R443 B.n209 B.n208 163.367
R444 B.n208 B.n203 163.367
R445 B.n204 B.n203 163.367
R446 B.n204 B.n2 163.367
R447 B.n786 B.n2 163.367
R448 B.n786 B.n785 163.367
R449 B.n785 B.n784 163.367
R450 B.n784 B.n3 163.367
R451 B.n780 B.n3 163.367
R452 B.n780 B.n779 163.367
R453 B.n779 B.n778 163.367
R454 B.n778 B.n5 163.367
R455 B.n774 B.n5 163.367
R456 B.n774 B.n773 163.367
R457 B.n773 B.n772 163.367
R458 B.n772 B.n7 163.367
R459 B.n768 B.n7 163.367
R460 B.n768 B.n767 163.367
R461 B.n767 B.n766 163.367
R462 B.n766 B.n9 163.367
R463 B.n762 B.n9 163.367
R464 B.n762 B.n761 163.367
R465 B.n761 B.n760 163.367
R466 B.n760 B.n11 163.367
R467 B.n756 B.n11 163.367
R468 B.n756 B.n755 163.367
R469 B.n755 B.n754 163.367
R470 B.n754 B.n13 163.367
R471 B.n750 B.n13 163.367
R472 B.n750 B.n749 163.367
R473 B.n749 B.n748 163.367
R474 B.n748 B.n15 163.367
R475 B.n744 B.n15 163.367
R476 B.n744 B.n743 163.367
R477 B.n743 B.n742 163.367
R478 B.n742 B.n17 163.367
R479 B.n738 B.n17 163.367
R480 B.n738 B.n737 163.367
R481 B.n737 B.n736 163.367
R482 B.n736 B.n19 163.367
R483 B.n732 B.n19 163.367
R484 B.n732 B.n731 163.367
R485 B.n731 B.n730 163.367
R486 B.n730 B.n21 163.367
R487 B.n726 B.n21 163.367
R488 B.n726 B.n725 163.367
R489 B.n725 B.n724 163.367
R490 B.n724 B.n23 163.367
R491 B.n720 B.n23 163.367
R492 B.n270 B.n269 163.367
R493 B.n270 B.n181 163.367
R494 B.n274 B.n181 163.367
R495 B.n275 B.n274 163.367
R496 B.n276 B.n275 163.367
R497 B.n276 B.n179 163.367
R498 B.n280 B.n179 163.367
R499 B.n281 B.n280 163.367
R500 B.n282 B.n281 163.367
R501 B.n282 B.n177 163.367
R502 B.n286 B.n177 163.367
R503 B.n287 B.n286 163.367
R504 B.n288 B.n287 163.367
R505 B.n288 B.n175 163.367
R506 B.n292 B.n175 163.367
R507 B.n293 B.n292 163.367
R508 B.n294 B.n293 163.367
R509 B.n294 B.n173 163.367
R510 B.n298 B.n173 163.367
R511 B.n299 B.n298 163.367
R512 B.n300 B.n299 163.367
R513 B.n300 B.n171 163.367
R514 B.n304 B.n171 163.367
R515 B.n305 B.n304 163.367
R516 B.n306 B.n305 163.367
R517 B.n306 B.n169 163.367
R518 B.n310 B.n169 163.367
R519 B.n311 B.n310 163.367
R520 B.n312 B.n311 163.367
R521 B.n312 B.n167 163.367
R522 B.n316 B.n167 163.367
R523 B.n317 B.n316 163.367
R524 B.n318 B.n317 163.367
R525 B.n318 B.n165 163.367
R526 B.n322 B.n165 163.367
R527 B.n323 B.n322 163.367
R528 B.n324 B.n323 163.367
R529 B.n324 B.n163 163.367
R530 B.n328 B.n163 163.367
R531 B.n329 B.n328 163.367
R532 B.n330 B.n329 163.367
R533 B.n330 B.n161 163.367
R534 B.n334 B.n161 163.367
R535 B.n335 B.n334 163.367
R536 B.n336 B.n335 163.367
R537 B.n336 B.n159 163.367
R538 B.n340 B.n159 163.367
R539 B.n341 B.n340 163.367
R540 B.n341 B.n155 163.367
R541 B.n345 B.n155 163.367
R542 B.n346 B.n345 163.367
R543 B.n347 B.n346 163.367
R544 B.n347 B.n153 163.367
R545 B.n351 B.n153 163.367
R546 B.n352 B.n351 163.367
R547 B.n353 B.n352 163.367
R548 B.n353 B.n149 163.367
R549 B.n358 B.n149 163.367
R550 B.n359 B.n358 163.367
R551 B.n360 B.n359 163.367
R552 B.n360 B.n147 163.367
R553 B.n364 B.n147 163.367
R554 B.n365 B.n364 163.367
R555 B.n366 B.n365 163.367
R556 B.n366 B.n145 163.367
R557 B.n370 B.n145 163.367
R558 B.n371 B.n370 163.367
R559 B.n372 B.n371 163.367
R560 B.n372 B.n143 163.367
R561 B.n376 B.n143 163.367
R562 B.n377 B.n376 163.367
R563 B.n378 B.n377 163.367
R564 B.n378 B.n141 163.367
R565 B.n382 B.n141 163.367
R566 B.n383 B.n382 163.367
R567 B.n384 B.n383 163.367
R568 B.n384 B.n139 163.367
R569 B.n388 B.n139 163.367
R570 B.n389 B.n388 163.367
R571 B.n390 B.n389 163.367
R572 B.n390 B.n137 163.367
R573 B.n394 B.n137 163.367
R574 B.n395 B.n394 163.367
R575 B.n396 B.n395 163.367
R576 B.n396 B.n135 163.367
R577 B.n400 B.n135 163.367
R578 B.n401 B.n400 163.367
R579 B.n402 B.n401 163.367
R580 B.n402 B.n133 163.367
R581 B.n406 B.n133 163.367
R582 B.n407 B.n406 163.367
R583 B.n408 B.n407 163.367
R584 B.n408 B.n131 163.367
R585 B.n412 B.n131 163.367
R586 B.n413 B.n412 163.367
R587 B.n414 B.n413 163.367
R588 B.n414 B.n129 163.367
R589 B.n418 B.n129 163.367
R590 B.n419 B.n418 163.367
R591 B.n420 B.n419 163.367
R592 B.n420 B.n127 163.367
R593 B.n424 B.n127 163.367
R594 B.n425 B.n424 163.367
R595 B.n426 B.n425 163.367
R596 B.n430 B.n125 163.367
R597 B.n431 B.n430 163.367
R598 B.n432 B.n431 163.367
R599 B.n432 B.n123 163.367
R600 B.n436 B.n123 163.367
R601 B.n437 B.n436 163.367
R602 B.n438 B.n437 163.367
R603 B.n438 B.n121 163.367
R604 B.n442 B.n121 163.367
R605 B.n443 B.n442 163.367
R606 B.n444 B.n443 163.367
R607 B.n444 B.n119 163.367
R608 B.n448 B.n119 163.367
R609 B.n449 B.n448 163.367
R610 B.n450 B.n449 163.367
R611 B.n450 B.n117 163.367
R612 B.n454 B.n117 163.367
R613 B.n455 B.n454 163.367
R614 B.n456 B.n455 163.367
R615 B.n456 B.n115 163.367
R616 B.n460 B.n115 163.367
R617 B.n461 B.n460 163.367
R618 B.n462 B.n461 163.367
R619 B.n462 B.n113 163.367
R620 B.n466 B.n113 163.367
R621 B.n467 B.n466 163.367
R622 B.n468 B.n467 163.367
R623 B.n468 B.n111 163.367
R624 B.n472 B.n111 163.367
R625 B.n473 B.n472 163.367
R626 B.n474 B.n473 163.367
R627 B.n474 B.n109 163.367
R628 B.n478 B.n109 163.367
R629 B.n479 B.n478 163.367
R630 B.n480 B.n479 163.367
R631 B.n480 B.n107 163.367
R632 B.n484 B.n107 163.367
R633 B.n485 B.n484 163.367
R634 B.n486 B.n485 163.367
R635 B.n486 B.n105 163.367
R636 B.n490 B.n105 163.367
R637 B.n491 B.n490 163.367
R638 B.n492 B.n491 163.367
R639 B.n492 B.n103 163.367
R640 B.n496 B.n103 163.367
R641 B.n497 B.n496 163.367
R642 B.n498 B.n497 163.367
R643 B.n498 B.n101 163.367
R644 B.n502 B.n101 163.367
R645 B.n503 B.n502 163.367
R646 B.n504 B.n503 163.367
R647 B.n504 B.n99 163.367
R648 B.n508 B.n99 163.367
R649 B.n509 B.n508 163.367
R650 B.n510 B.n509 163.367
R651 B.n510 B.n97 163.367
R652 B.n514 B.n97 163.367
R653 B.n515 B.n514 163.367
R654 B.n516 B.n515 163.367
R655 B.n516 B.n95 163.367
R656 B.n520 B.n95 163.367
R657 B.n521 B.n520 163.367
R658 B.n522 B.n521 163.367
R659 B.n522 B.n93 163.367
R660 B.n526 B.n93 163.367
R661 B.n527 B.n526 163.367
R662 B.n528 B.n527 163.367
R663 B.n528 B.n91 163.367
R664 B.n532 B.n91 163.367
R665 B.n533 B.n532 163.367
R666 B.n534 B.n533 163.367
R667 B.n534 B.n89 163.367
R668 B.n538 B.n89 163.367
R669 B.n539 B.n538 163.367
R670 B.n540 B.n539 163.367
R671 B.n540 B.n87 163.367
R672 B.n544 B.n87 163.367
R673 B.n545 B.n544 163.367
R674 B.n546 B.n545 163.367
R675 B.n546 B.n85 163.367
R676 B.n550 B.n85 163.367
R677 B.n551 B.n550 163.367
R678 B.n552 B.n551 163.367
R679 B.n552 B.n83 163.367
R680 B.n556 B.n83 163.367
R681 B.n557 B.n556 163.367
R682 B.n558 B.n557 163.367
R683 B.n558 B.n81 163.367
R684 B.n719 B.n718 163.367
R685 B.n718 B.n25 163.367
R686 B.n714 B.n25 163.367
R687 B.n714 B.n713 163.367
R688 B.n713 B.n712 163.367
R689 B.n712 B.n27 163.367
R690 B.n708 B.n27 163.367
R691 B.n708 B.n707 163.367
R692 B.n707 B.n706 163.367
R693 B.n706 B.n29 163.367
R694 B.n702 B.n29 163.367
R695 B.n702 B.n701 163.367
R696 B.n701 B.n700 163.367
R697 B.n700 B.n31 163.367
R698 B.n696 B.n31 163.367
R699 B.n696 B.n695 163.367
R700 B.n695 B.n694 163.367
R701 B.n694 B.n33 163.367
R702 B.n690 B.n33 163.367
R703 B.n690 B.n689 163.367
R704 B.n689 B.n688 163.367
R705 B.n688 B.n35 163.367
R706 B.n684 B.n35 163.367
R707 B.n684 B.n683 163.367
R708 B.n683 B.n682 163.367
R709 B.n682 B.n37 163.367
R710 B.n678 B.n37 163.367
R711 B.n678 B.n677 163.367
R712 B.n677 B.n676 163.367
R713 B.n676 B.n39 163.367
R714 B.n672 B.n39 163.367
R715 B.n672 B.n671 163.367
R716 B.n671 B.n670 163.367
R717 B.n670 B.n41 163.367
R718 B.n666 B.n41 163.367
R719 B.n666 B.n665 163.367
R720 B.n665 B.n664 163.367
R721 B.n664 B.n43 163.367
R722 B.n660 B.n43 163.367
R723 B.n660 B.n659 163.367
R724 B.n659 B.n658 163.367
R725 B.n658 B.n45 163.367
R726 B.n654 B.n45 163.367
R727 B.n654 B.n653 163.367
R728 B.n653 B.n652 163.367
R729 B.n652 B.n47 163.367
R730 B.n648 B.n47 163.367
R731 B.n648 B.n647 163.367
R732 B.n647 B.n51 163.367
R733 B.n643 B.n51 163.367
R734 B.n643 B.n642 163.367
R735 B.n642 B.n641 163.367
R736 B.n641 B.n53 163.367
R737 B.n637 B.n53 163.367
R738 B.n637 B.n636 163.367
R739 B.n636 B.n635 163.367
R740 B.n635 B.n55 163.367
R741 B.n630 B.n55 163.367
R742 B.n630 B.n629 163.367
R743 B.n629 B.n628 163.367
R744 B.n628 B.n59 163.367
R745 B.n624 B.n59 163.367
R746 B.n624 B.n623 163.367
R747 B.n623 B.n622 163.367
R748 B.n622 B.n61 163.367
R749 B.n618 B.n61 163.367
R750 B.n618 B.n617 163.367
R751 B.n617 B.n616 163.367
R752 B.n616 B.n63 163.367
R753 B.n612 B.n63 163.367
R754 B.n612 B.n611 163.367
R755 B.n611 B.n610 163.367
R756 B.n610 B.n65 163.367
R757 B.n606 B.n65 163.367
R758 B.n606 B.n605 163.367
R759 B.n605 B.n604 163.367
R760 B.n604 B.n67 163.367
R761 B.n600 B.n67 163.367
R762 B.n600 B.n599 163.367
R763 B.n599 B.n598 163.367
R764 B.n598 B.n69 163.367
R765 B.n594 B.n69 163.367
R766 B.n594 B.n593 163.367
R767 B.n593 B.n592 163.367
R768 B.n592 B.n71 163.367
R769 B.n588 B.n71 163.367
R770 B.n588 B.n587 163.367
R771 B.n587 B.n586 163.367
R772 B.n586 B.n73 163.367
R773 B.n582 B.n73 163.367
R774 B.n582 B.n581 163.367
R775 B.n581 B.n580 163.367
R776 B.n580 B.n75 163.367
R777 B.n576 B.n75 163.367
R778 B.n576 B.n575 163.367
R779 B.n575 B.n574 163.367
R780 B.n574 B.n77 163.367
R781 B.n570 B.n77 163.367
R782 B.n570 B.n569 163.367
R783 B.n569 B.n568 163.367
R784 B.n568 B.n79 163.367
R785 B.n564 B.n79 163.367
R786 B.n564 B.n563 163.367
R787 B.n563 B.n562 163.367
R788 B.n151 B.n150 79.3217
R789 B.n157 B.n156 79.3217
R790 B.n49 B.n48 79.3217
R791 B.n57 B.n56 79.3217
R792 B.n355 B.n151 59.5399
R793 B.n158 B.n157 59.5399
R794 B.n50 B.n49 59.5399
R795 B.n633 B.n57 59.5399
R796 B.n561 B.n560 35.7468
R797 B.n721 B.n24 35.7468
R798 B.n428 B.n427 35.7468
R799 B.n267 B.n182 35.7468
R800 B B.n787 18.0485
R801 B.n717 B.n24 10.6151
R802 B.n717 B.n716 10.6151
R803 B.n716 B.n715 10.6151
R804 B.n715 B.n26 10.6151
R805 B.n711 B.n26 10.6151
R806 B.n711 B.n710 10.6151
R807 B.n710 B.n709 10.6151
R808 B.n709 B.n28 10.6151
R809 B.n705 B.n28 10.6151
R810 B.n705 B.n704 10.6151
R811 B.n704 B.n703 10.6151
R812 B.n703 B.n30 10.6151
R813 B.n699 B.n30 10.6151
R814 B.n699 B.n698 10.6151
R815 B.n698 B.n697 10.6151
R816 B.n697 B.n32 10.6151
R817 B.n693 B.n32 10.6151
R818 B.n693 B.n692 10.6151
R819 B.n692 B.n691 10.6151
R820 B.n691 B.n34 10.6151
R821 B.n687 B.n34 10.6151
R822 B.n687 B.n686 10.6151
R823 B.n686 B.n685 10.6151
R824 B.n685 B.n36 10.6151
R825 B.n681 B.n36 10.6151
R826 B.n681 B.n680 10.6151
R827 B.n680 B.n679 10.6151
R828 B.n679 B.n38 10.6151
R829 B.n675 B.n38 10.6151
R830 B.n675 B.n674 10.6151
R831 B.n674 B.n673 10.6151
R832 B.n673 B.n40 10.6151
R833 B.n669 B.n40 10.6151
R834 B.n669 B.n668 10.6151
R835 B.n668 B.n667 10.6151
R836 B.n667 B.n42 10.6151
R837 B.n663 B.n42 10.6151
R838 B.n663 B.n662 10.6151
R839 B.n662 B.n661 10.6151
R840 B.n661 B.n44 10.6151
R841 B.n657 B.n44 10.6151
R842 B.n657 B.n656 10.6151
R843 B.n656 B.n655 10.6151
R844 B.n655 B.n46 10.6151
R845 B.n651 B.n46 10.6151
R846 B.n651 B.n650 10.6151
R847 B.n650 B.n649 10.6151
R848 B.n646 B.n645 10.6151
R849 B.n645 B.n644 10.6151
R850 B.n644 B.n52 10.6151
R851 B.n640 B.n52 10.6151
R852 B.n640 B.n639 10.6151
R853 B.n639 B.n638 10.6151
R854 B.n638 B.n54 10.6151
R855 B.n634 B.n54 10.6151
R856 B.n632 B.n631 10.6151
R857 B.n631 B.n58 10.6151
R858 B.n627 B.n58 10.6151
R859 B.n627 B.n626 10.6151
R860 B.n626 B.n625 10.6151
R861 B.n625 B.n60 10.6151
R862 B.n621 B.n60 10.6151
R863 B.n621 B.n620 10.6151
R864 B.n620 B.n619 10.6151
R865 B.n619 B.n62 10.6151
R866 B.n615 B.n62 10.6151
R867 B.n615 B.n614 10.6151
R868 B.n614 B.n613 10.6151
R869 B.n613 B.n64 10.6151
R870 B.n609 B.n64 10.6151
R871 B.n609 B.n608 10.6151
R872 B.n608 B.n607 10.6151
R873 B.n607 B.n66 10.6151
R874 B.n603 B.n66 10.6151
R875 B.n603 B.n602 10.6151
R876 B.n602 B.n601 10.6151
R877 B.n601 B.n68 10.6151
R878 B.n597 B.n68 10.6151
R879 B.n597 B.n596 10.6151
R880 B.n596 B.n595 10.6151
R881 B.n595 B.n70 10.6151
R882 B.n591 B.n70 10.6151
R883 B.n591 B.n590 10.6151
R884 B.n590 B.n589 10.6151
R885 B.n589 B.n72 10.6151
R886 B.n585 B.n72 10.6151
R887 B.n585 B.n584 10.6151
R888 B.n584 B.n583 10.6151
R889 B.n583 B.n74 10.6151
R890 B.n579 B.n74 10.6151
R891 B.n579 B.n578 10.6151
R892 B.n578 B.n577 10.6151
R893 B.n577 B.n76 10.6151
R894 B.n573 B.n76 10.6151
R895 B.n573 B.n572 10.6151
R896 B.n572 B.n571 10.6151
R897 B.n571 B.n78 10.6151
R898 B.n567 B.n78 10.6151
R899 B.n567 B.n566 10.6151
R900 B.n566 B.n565 10.6151
R901 B.n565 B.n80 10.6151
R902 B.n561 B.n80 10.6151
R903 B.n429 B.n428 10.6151
R904 B.n429 B.n124 10.6151
R905 B.n433 B.n124 10.6151
R906 B.n434 B.n433 10.6151
R907 B.n435 B.n434 10.6151
R908 B.n435 B.n122 10.6151
R909 B.n439 B.n122 10.6151
R910 B.n440 B.n439 10.6151
R911 B.n441 B.n440 10.6151
R912 B.n441 B.n120 10.6151
R913 B.n445 B.n120 10.6151
R914 B.n446 B.n445 10.6151
R915 B.n447 B.n446 10.6151
R916 B.n447 B.n118 10.6151
R917 B.n451 B.n118 10.6151
R918 B.n452 B.n451 10.6151
R919 B.n453 B.n452 10.6151
R920 B.n453 B.n116 10.6151
R921 B.n457 B.n116 10.6151
R922 B.n458 B.n457 10.6151
R923 B.n459 B.n458 10.6151
R924 B.n459 B.n114 10.6151
R925 B.n463 B.n114 10.6151
R926 B.n464 B.n463 10.6151
R927 B.n465 B.n464 10.6151
R928 B.n465 B.n112 10.6151
R929 B.n469 B.n112 10.6151
R930 B.n470 B.n469 10.6151
R931 B.n471 B.n470 10.6151
R932 B.n471 B.n110 10.6151
R933 B.n475 B.n110 10.6151
R934 B.n476 B.n475 10.6151
R935 B.n477 B.n476 10.6151
R936 B.n477 B.n108 10.6151
R937 B.n481 B.n108 10.6151
R938 B.n482 B.n481 10.6151
R939 B.n483 B.n482 10.6151
R940 B.n483 B.n106 10.6151
R941 B.n487 B.n106 10.6151
R942 B.n488 B.n487 10.6151
R943 B.n489 B.n488 10.6151
R944 B.n489 B.n104 10.6151
R945 B.n493 B.n104 10.6151
R946 B.n494 B.n493 10.6151
R947 B.n495 B.n494 10.6151
R948 B.n495 B.n102 10.6151
R949 B.n499 B.n102 10.6151
R950 B.n500 B.n499 10.6151
R951 B.n501 B.n500 10.6151
R952 B.n501 B.n100 10.6151
R953 B.n505 B.n100 10.6151
R954 B.n506 B.n505 10.6151
R955 B.n507 B.n506 10.6151
R956 B.n507 B.n98 10.6151
R957 B.n511 B.n98 10.6151
R958 B.n512 B.n511 10.6151
R959 B.n513 B.n512 10.6151
R960 B.n513 B.n96 10.6151
R961 B.n517 B.n96 10.6151
R962 B.n518 B.n517 10.6151
R963 B.n519 B.n518 10.6151
R964 B.n519 B.n94 10.6151
R965 B.n523 B.n94 10.6151
R966 B.n524 B.n523 10.6151
R967 B.n525 B.n524 10.6151
R968 B.n525 B.n92 10.6151
R969 B.n529 B.n92 10.6151
R970 B.n530 B.n529 10.6151
R971 B.n531 B.n530 10.6151
R972 B.n531 B.n90 10.6151
R973 B.n535 B.n90 10.6151
R974 B.n536 B.n535 10.6151
R975 B.n537 B.n536 10.6151
R976 B.n537 B.n88 10.6151
R977 B.n541 B.n88 10.6151
R978 B.n542 B.n541 10.6151
R979 B.n543 B.n542 10.6151
R980 B.n543 B.n86 10.6151
R981 B.n547 B.n86 10.6151
R982 B.n548 B.n547 10.6151
R983 B.n549 B.n548 10.6151
R984 B.n549 B.n84 10.6151
R985 B.n553 B.n84 10.6151
R986 B.n554 B.n553 10.6151
R987 B.n555 B.n554 10.6151
R988 B.n555 B.n82 10.6151
R989 B.n559 B.n82 10.6151
R990 B.n560 B.n559 10.6151
R991 B.n271 B.n182 10.6151
R992 B.n272 B.n271 10.6151
R993 B.n273 B.n272 10.6151
R994 B.n273 B.n180 10.6151
R995 B.n277 B.n180 10.6151
R996 B.n278 B.n277 10.6151
R997 B.n279 B.n278 10.6151
R998 B.n279 B.n178 10.6151
R999 B.n283 B.n178 10.6151
R1000 B.n284 B.n283 10.6151
R1001 B.n285 B.n284 10.6151
R1002 B.n285 B.n176 10.6151
R1003 B.n289 B.n176 10.6151
R1004 B.n290 B.n289 10.6151
R1005 B.n291 B.n290 10.6151
R1006 B.n291 B.n174 10.6151
R1007 B.n295 B.n174 10.6151
R1008 B.n296 B.n295 10.6151
R1009 B.n297 B.n296 10.6151
R1010 B.n297 B.n172 10.6151
R1011 B.n301 B.n172 10.6151
R1012 B.n302 B.n301 10.6151
R1013 B.n303 B.n302 10.6151
R1014 B.n303 B.n170 10.6151
R1015 B.n307 B.n170 10.6151
R1016 B.n308 B.n307 10.6151
R1017 B.n309 B.n308 10.6151
R1018 B.n309 B.n168 10.6151
R1019 B.n313 B.n168 10.6151
R1020 B.n314 B.n313 10.6151
R1021 B.n315 B.n314 10.6151
R1022 B.n315 B.n166 10.6151
R1023 B.n319 B.n166 10.6151
R1024 B.n320 B.n319 10.6151
R1025 B.n321 B.n320 10.6151
R1026 B.n321 B.n164 10.6151
R1027 B.n325 B.n164 10.6151
R1028 B.n326 B.n325 10.6151
R1029 B.n327 B.n326 10.6151
R1030 B.n327 B.n162 10.6151
R1031 B.n331 B.n162 10.6151
R1032 B.n332 B.n331 10.6151
R1033 B.n333 B.n332 10.6151
R1034 B.n333 B.n160 10.6151
R1035 B.n337 B.n160 10.6151
R1036 B.n338 B.n337 10.6151
R1037 B.n339 B.n338 10.6151
R1038 B.n343 B.n342 10.6151
R1039 B.n344 B.n343 10.6151
R1040 B.n344 B.n154 10.6151
R1041 B.n348 B.n154 10.6151
R1042 B.n349 B.n348 10.6151
R1043 B.n350 B.n349 10.6151
R1044 B.n350 B.n152 10.6151
R1045 B.n354 B.n152 10.6151
R1046 B.n357 B.n356 10.6151
R1047 B.n357 B.n148 10.6151
R1048 B.n361 B.n148 10.6151
R1049 B.n362 B.n361 10.6151
R1050 B.n363 B.n362 10.6151
R1051 B.n363 B.n146 10.6151
R1052 B.n367 B.n146 10.6151
R1053 B.n368 B.n367 10.6151
R1054 B.n369 B.n368 10.6151
R1055 B.n369 B.n144 10.6151
R1056 B.n373 B.n144 10.6151
R1057 B.n374 B.n373 10.6151
R1058 B.n375 B.n374 10.6151
R1059 B.n375 B.n142 10.6151
R1060 B.n379 B.n142 10.6151
R1061 B.n380 B.n379 10.6151
R1062 B.n381 B.n380 10.6151
R1063 B.n381 B.n140 10.6151
R1064 B.n385 B.n140 10.6151
R1065 B.n386 B.n385 10.6151
R1066 B.n387 B.n386 10.6151
R1067 B.n387 B.n138 10.6151
R1068 B.n391 B.n138 10.6151
R1069 B.n392 B.n391 10.6151
R1070 B.n393 B.n392 10.6151
R1071 B.n393 B.n136 10.6151
R1072 B.n397 B.n136 10.6151
R1073 B.n398 B.n397 10.6151
R1074 B.n399 B.n398 10.6151
R1075 B.n399 B.n134 10.6151
R1076 B.n403 B.n134 10.6151
R1077 B.n404 B.n403 10.6151
R1078 B.n405 B.n404 10.6151
R1079 B.n405 B.n132 10.6151
R1080 B.n409 B.n132 10.6151
R1081 B.n410 B.n409 10.6151
R1082 B.n411 B.n410 10.6151
R1083 B.n411 B.n130 10.6151
R1084 B.n415 B.n130 10.6151
R1085 B.n416 B.n415 10.6151
R1086 B.n417 B.n416 10.6151
R1087 B.n417 B.n128 10.6151
R1088 B.n421 B.n128 10.6151
R1089 B.n422 B.n421 10.6151
R1090 B.n423 B.n422 10.6151
R1091 B.n423 B.n126 10.6151
R1092 B.n427 B.n126 10.6151
R1093 B.n267 B.n266 10.6151
R1094 B.n266 B.n265 10.6151
R1095 B.n265 B.n184 10.6151
R1096 B.n261 B.n184 10.6151
R1097 B.n261 B.n260 10.6151
R1098 B.n260 B.n259 10.6151
R1099 B.n259 B.n186 10.6151
R1100 B.n255 B.n186 10.6151
R1101 B.n255 B.n254 10.6151
R1102 B.n254 B.n253 10.6151
R1103 B.n253 B.n188 10.6151
R1104 B.n249 B.n188 10.6151
R1105 B.n249 B.n248 10.6151
R1106 B.n248 B.n247 10.6151
R1107 B.n247 B.n190 10.6151
R1108 B.n243 B.n190 10.6151
R1109 B.n243 B.n242 10.6151
R1110 B.n242 B.n241 10.6151
R1111 B.n241 B.n192 10.6151
R1112 B.n237 B.n192 10.6151
R1113 B.n237 B.n236 10.6151
R1114 B.n236 B.n235 10.6151
R1115 B.n235 B.n194 10.6151
R1116 B.n231 B.n194 10.6151
R1117 B.n231 B.n230 10.6151
R1118 B.n230 B.n229 10.6151
R1119 B.n229 B.n196 10.6151
R1120 B.n225 B.n196 10.6151
R1121 B.n225 B.n224 10.6151
R1122 B.n224 B.n223 10.6151
R1123 B.n223 B.n198 10.6151
R1124 B.n219 B.n198 10.6151
R1125 B.n219 B.n218 10.6151
R1126 B.n218 B.n217 10.6151
R1127 B.n217 B.n200 10.6151
R1128 B.n213 B.n200 10.6151
R1129 B.n213 B.n212 10.6151
R1130 B.n212 B.n211 10.6151
R1131 B.n211 B.n202 10.6151
R1132 B.n207 B.n202 10.6151
R1133 B.n207 B.n206 10.6151
R1134 B.n206 B.n205 10.6151
R1135 B.n205 B.n0 10.6151
R1136 B.n783 B.n1 10.6151
R1137 B.n783 B.n782 10.6151
R1138 B.n782 B.n781 10.6151
R1139 B.n781 B.n4 10.6151
R1140 B.n777 B.n4 10.6151
R1141 B.n777 B.n776 10.6151
R1142 B.n776 B.n775 10.6151
R1143 B.n775 B.n6 10.6151
R1144 B.n771 B.n6 10.6151
R1145 B.n771 B.n770 10.6151
R1146 B.n770 B.n769 10.6151
R1147 B.n769 B.n8 10.6151
R1148 B.n765 B.n8 10.6151
R1149 B.n765 B.n764 10.6151
R1150 B.n764 B.n763 10.6151
R1151 B.n763 B.n10 10.6151
R1152 B.n759 B.n10 10.6151
R1153 B.n759 B.n758 10.6151
R1154 B.n758 B.n757 10.6151
R1155 B.n757 B.n12 10.6151
R1156 B.n753 B.n12 10.6151
R1157 B.n753 B.n752 10.6151
R1158 B.n752 B.n751 10.6151
R1159 B.n751 B.n14 10.6151
R1160 B.n747 B.n14 10.6151
R1161 B.n747 B.n746 10.6151
R1162 B.n746 B.n745 10.6151
R1163 B.n745 B.n16 10.6151
R1164 B.n741 B.n16 10.6151
R1165 B.n741 B.n740 10.6151
R1166 B.n740 B.n739 10.6151
R1167 B.n739 B.n18 10.6151
R1168 B.n735 B.n18 10.6151
R1169 B.n735 B.n734 10.6151
R1170 B.n734 B.n733 10.6151
R1171 B.n733 B.n20 10.6151
R1172 B.n729 B.n20 10.6151
R1173 B.n729 B.n728 10.6151
R1174 B.n728 B.n727 10.6151
R1175 B.n727 B.n22 10.6151
R1176 B.n723 B.n22 10.6151
R1177 B.n723 B.n722 10.6151
R1178 B.n722 B.n721 10.6151
R1179 B.n646 B.n50 6.5566
R1180 B.n634 B.n633 6.5566
R1181 B.n342 B.n158 6.5566
R1182 B.n355 B.n354 6.5566
R1183 B.n649 B.n50 4.05904
R1184 B.n633 B.n632 4.05904
R1185 B.n339 B.n158 4.05904
R1186 B.n356 B.n355 4.05904
R1187 B.n787 B.n0 2.81026
R1188 B.n787 B.n1 2.81026
R1189 VN.n0 VN.t0 124.126
R1190 VN.n1 VN.t2 124.126
R1191 VN.n0 VN.t3 122.784
R1192 VN.n1 VN.t1 122.784
R1193 VN VN.n1 53.5439
R1194 VN VN.n0 1.88864
R1195 VDD2.n2 VDD2.n0 121.475
R1196 VDD2.n2 VDD2.n1 75.019
R1197 VDD2.n1 VDD2.t2 2.30419
R1198 VDD2.n1 VDD2.t0 2.30419
R1199 VDD2.n0 VDD2.t3 2.30419
R1200 VDD2.n0 VDD2.t1 2.30419
R1201 VDD2 VDD2.n2 0.0586897
R1202 VTAIL.n618 VTAIL.n546 756.745
R1203 VTAIL.n72 VTAIL.n0 756.745
R1204 VTAIL.n150 VTAIL.n78 756.745
R1205 VTAIL.n228 VTAIL.n156 756.745
R1206 VTAIL.n540 VTAIL.n468 756.745
R1207 VTAIL.n462 VTAIL.n390 756.745
R1208 VTAIL.n384 VTAIL.n312 756.745
R1209 VTAIL.n306 VTAIL.n234 756.745
R1210 VTAIL.n570 VTAIL.n569 585
R1211 VTAIL.n575 VTAIL.n574 585
R1212 VTAIL.n577 VTAIL.n576 585
R1213 VTAIL.n566 VTAIL.n565 585
R1214 VTAIL.n583 VTAIL.n582 585
R1215 VTAIL.n585 VTAIL.n584 585
R1216 VTAIL.n562 VTAIL.n561 585
R1217 VTAIL.n591 VTAIL.n590 585
R1218 VTAIL.n593 VTAIL.n592 585
R1219 VTAIL.n558 VTAIL.n557 585
R1220 VTAIL.n599 VTAIL.n598 585
R1221 VTAIL.n601 VTAIL.n600 585
R1222 VTAIL.n554 VTAIL.n553 585
R1223 VTAIL.n607 VTAIL.n606 585
R1224 VTAIL.n609 VTAIL.n608 585
R1225 VTAIL.n550 VTAIL.n549 585
R1226 VTAIL.n616 VTAIL.n615 585
R1227 VTAIL.n617 VTAIL.n548 585
R1228 VTAIL.n619 VTAIL.n618 585
R1229 VTAIL.n24 VTAIL.n23 585
R1230 VTAIL.n29 VTAIL.n28 585
R1231 VTAIL.n31 VTAIL.n30 585
R1232 VTAIL.n20 VTAIL.n19 585
R1233 VTAIL.n37 VTAIL.n36 585
R1234 VTAIL.n39 VTAIL.n38 585
R1235 VTAIL.n16 VTAIL.n15 585
R1236 VTAIL.n45 VTAIL.n44 585
R1237 VTAIL.n47 VTAIL.n46 585
R1238 VTAIL.n12 VTAIL.n11 585
R1239 VTAIL.n53 VTAIL.n52 585
R1240 VTAIL.n55 VTAIL.n54 585
R1241 VTAIL.n8 VTAIL.n7 585
R1242 VTAIL.n61 VTAIL.n60 585
R1243 VTAIL.n63 VTAIL.n62 585
R1244 VTAIL.n4 VTAIL.n3 585
R1245 VTAIL.n70 VTAIL.n69 585
R1246 VTAIL.n71 VTAIL.n2 585
R1247 VTAIL.n73 VTAIL.n72 585
R1248 VTAIL.n102 VTAIL.n101 585
R1249 VTAIL.n107 VTAIL.n106 585
R1250 VTAIL.n109 VTAIL.n108 585
R1251 VTAIL.n98 VTAIL.n97 585
R1252 VTAIL.n115 VTAIL.n114 585
R1253 VTAIL.n117 VTAIL.n116 585
R1254 VTAIL.n94 VTAIL.n93 585
R1255 VTAIL.n123 VTAIL.n122 585
R1256 VTAIL.n125 VTAIL.n124 585
R1257 VTAIL.n90 VTAIL.n89 585
R1258 VTAIL.n131 VTAIL.n130 585
R1259 VTAIL.n133 VTAIL.n132 585
R1260 VTAIL.n86 VTAIL.n85 585
R1261 VTAIL.n139 VTAIL.n138 585
R1262 VTAIL.n141 VTAIL.n140 585
R1263 VTAIL.n82 VTAIL.n81 585
R1264 VTAIL.n148 VTAIL.n147 585
R1265 VTAIL.n149 VTAIL.n80 585
R1266 VTAIL.n151 VTAIL.n150 585
R1267 VTAIL.n180 VTAIL.n179 585
R1268 VTAIL.n185 VTAIL.n184 585
R1269 VTAIL.n187 VTAIL.n186 585
R1270 VTAIL.n176 VTAIL.n175 585
R1271 VTAIL.n193 VTAIL.n192 585
R1272 VTAIL.n195 VTAIL.n194 585
R1273 VTAIL.n172 VTAIL.n171 585
R1274 VTAIL.n201 VTAIL.n200 585
R1275 VTAIL.n203 VTAIL.n202 585
R1276 VTAIL.n168 VTAIL.n167 585
R1277 VTAIL.n209 VTAIL.n208 585
R1278 VTAIL.n211 VTAIL.n210 585
R1279 VTAIL.n164 VTAIL.n163 585
R1280 VTAIL.n217 VTAIL.n216 585
R1281 VTAIL.n219 VTAIL.n218 585
R1282 VTAIL.n160 VTAIL.n159 585
R1283 VTAIL.n226 VTAIL.n225 585
R1284 VTAIL.n227 VTAIL.n158 585
R1285 VTAIL.n229 VTAIL.n228 585
R1286 VTAIL.n541 VTAIL.n540 585
R1287 VTAIL.n539 VTAIL.n470 585
R1288 VTAIL.n538 VTAIL.n537 585
R1289 VTAIL.n473 VTAIL.n471 585
R1290 VTAIL.n532 VTAIL.n531 585
R1291 VTAIL.n530 VTAIL.n529 585
R1292 VTAIL.n477 VTAIL.n476 585
R1293 VTAIL.n524 VTAIL.n523 585
R1294 VTAIL.n522 VTAIL.n521 585
R1295 VTAIL.n481 VTAIL.n480 585
R1296 VTAIL.n516 VTAIL.n515 585
R1297 VTAIL.n514 VTAIL.n513 585
R1298 VTAIL.n485 VTAIL.n484 585
R1299 VTAIL.n508 VTAIL.n507 585
R1300 VTAIL.n506 VTAIL.n505 585
R1301 VTAIL.n489 VTAIL.n488 585
R1302 VTAIL.n500 VTAIL.n499 585
R1303 VTAIL.n498 VTAIL.n497 585
R1304 VTAIL.n493 VTAIL.n492 585
R1305 VTAIL.n463 VTAIL.n462 585
R1306 VTAIL.n461 VTAIL.n392 585
R1307 VTAIL.n460 VTAIL.n459 585
R1308 VTAIL.n395 VTAIL.n393 585
R1309 VTAIL.n454 VTAIL.n453 585
R1310 VTAIL.n452 VTAIL.n451 585
R1311 VTAIL.n399 VTAIL.n398 585
R1312 VTAIL.n446 VTAIL.n445 585
R1313 VTAIL.n444 VTAIL.n443 585
R1314 VTAIL.n403 VTAIL.n402 585
R1315 VTAIL.n438 VTAIL.n437 585
R1316 VTAIL.n436 VTAIL.n435 585
R1317 VTAIL.n407 VTAIL.n406 585
R1318 VTAIL.n430 VTAIL.n429 585
R1319 VTAIL.n428 VTAIL.n427 585
R1320 VTAIL.n411 VTAIL.n410 585
R1321 VTAIL.n422 VTAIL.n421 585
R1322 VTAIL.n420 VTAIL.n419 585
R1323 VTAIL.n415 VTAIL.n414 585
R1324 VTAIL.n385 VTAIL.n384 585
R1325 VTAIL.n383 VTAIL.n314 585
R1326 VTAIL.n382 VTAIL.n381 585
R1327 VTAIL.n317 VTAIL.n315 585
R1328 VTAIL.n376 VTAIL.n375 585
R1329 VTAIL.n374 VTAIL.n373 585
R1330 VTAIL.n321 VTAIL.n320 585
R1331 VTAIL.n368 VTAIL.n367 585
R1332 VTAIL.n366 VTAIL.n365 585
R1333 VTAIL.n325 VTAIL.n324 585
R1334 VTAIL.n360 VTAIL.n359 585
R1335 VTAIL.n358 VTAIL.n357 585
R1336 VTAIL.n329 VTAIL.n328 585
R1337 VTAIL.n352 VTAIL.n351 585
R1338 VTAIL.n350 VTAIL.n349 585
R1339 VTAIL.n333 VTAIL.n332 585
R1340 VTAIL.n344 VTAIL.n343 585
R1341 VTAIL.n342 VTAIL.n341 585
R1342 VTAIL.n337 VTAIL.n336 585
R1343 VTAIL.n307 VTAIL.n306 585
R1344 VTAIL.n305 VTAIL.n236 585
R1345 VTAIL.n304 VTAIL.n303 585
R1346 VTAIL.n239 VTAIL.n237 585
R1347 VTAIL.n298 VTAIL.n297 585
R1348 VTAIL.n296 VTAIL.n295 585
R1349 VTAIL.n243 VTAIL.n242 585
R1350 VTAIL.n290 VTAIL.n289 585
R1351 VTAIL.n288 VTAIL.n287 585
R1352 VTAIL.n247 VTAIL.n246 585
R1353 VTAIL.n282 VTAIL.n281 585
R1354 VTAIL.n280 VTAIL.n279 585
R1355 VTAIL.n251 VTAIL.n250 585
R1356 VTAIL.n274 VTAIL.n273 585
R1357 VTAIL.n272 VTAIL.n271 585
R1358 VTAIL.n255 VTAIL.n254 585
R1359 VTAIL.n266 VTAIL.n265 585
R1360 VTAIL.n264 VTAIL.n263 585
R1361 VTAIL.n259 VTAIL.n258 585
R1362 VTAIL.n571 VTAIL.t4 327.466
R1363 VTAIL.n25 VTAIL.t7 327.466
R1364 VTAIL.n103 VTAIL.t1 327.466
R1365 VTAIL.n181 VTAIL.t2 327.466
R1366 VTAIL.n494 VTAIL.t3 327.466
R1367 VTAIL.n416 VTAIL.t0 327.466
R1368 VTAIL.n338 VTAIL.t5 327.466
R1369 VTAIL.n260 VTAIL.t6 327.466
R1370 VTAIL.n575 VTAIL.n569 171.744
R1371 VTAIL.n576 VTAIL.n575 171.744
R1372 VTAIL.n576 VTAIL.n565 171.744
R1373 VTAIL.n583 VTAIL.n565 171.744
R1374 VTAIL.n584 VTAIL.n583 171.744
R1375 VTAIL.n584 VTAIL.n561 171.744
R1376 VTAIL.n591 VTAIL.n561 171.744
R1377 VTAIL.n592 VTAIL.n591 171.744
R1378 VTAIL.n592 VTAIL.n557 171.744
R1379 VTAIL.n599 VTAIL.n557 171.744
R1380 VTAIL.n600 VTAIL.n599 171.744
R1381 VTAIL.n600 VTAIL.n553 171.744
R1382 VTAIL.n607 VTAIL.n553 171.744
R1383 VTAIL.n608 VTAIL.n607 171.744
R1384 VTAIL.n608 VTAIL.n549 171.744
R1385 VTAIL.n616 VTAIL.n549 171.744
R1386 VTAIL.n617 VTAIL.n616 171.744
R1387 VTAIL.n618 VTAIL.n617 171.744
R1388 VTAIL.n29 VTAIL.n23 171.744
R1389 VTAIL.n30 VTAIL.n29 171.744
R1390 VTAIL.n30 VTAIL.n19 171.744
R1391 VTAIL.n37 VTAIL.n19 171.744
R1392 VTAIL.n38 VTAIL.n37 171.744
R1393 VTAIL.n38 VTAIL.n15 171.744
R1394 VTAIL.n45 VTAIL.n15 171.744
R1395 VTAIL.n46 VTAIL.n45 171.744
R1396 VTAIL.n46 VTAIL.n11 171.744
R1397 VTAIL.n53 VTAIL.n11 171.744
R1398 VTAIL.n54 VTAIL.n53 171.744
R1399 VTAIL.n54 VTAIL.n7 171.744
R1400 VTAIL.n61 VTAIL.n7 171.744
R1401 VTAIL.n62 VTAIL.n61 171.744
R1402 VTAIL.n62 VTAIL.n3 171.744
R1403 VTAIL.n70 VTAIL.n3 171.744
R1404 VTAIL.n71 VTAIL.n70 171.744
R1405 VTAIL.n72 VTAIL.n71 171.744
R1406 VTAIL.n107 VTAIL.n101 171.744
R1407 VTAIL.n108 VTAIL.n107 171.744
R1408 VTAIL.n108 VTAIL.n97 171.744
R1409 VTAIL.n115 VTAIL.n97 171.744
R1410 VTAIL.n116 VTAIL.n115 171.744
R1411 VTAIL.n116 VTAIL.n93 171.744
R1412 VTAIL.n123 VTAIL.n93 171.744
R1413 VTAIL.n124 VTAIL.n123 171.744
R1414 VTAIL.n124 VTAIL.n89 171.744
R1415 VTAIL.n131 VTAIL.n89 171.744
R1416 VTAIL.n132 VTAIL.n131 171.744
R1417 VTAIL.n132 VTAIL.n85 171.744
R1418 VTAIL.n139 VTAIL.n85 171.744
R1419 VTAIL.n140 VTAIL.n139 171.744
R1420 VTAIL.n140 VTAIL.n81 171.744
R1421 VTAIL.n148 VTAIL.n81 171.744
R1422 VTAIL.n149 VTAIL.n148 171.744
R1423 VTAIL.n150 VTAIL.n149 171.744
R1424 VTAIL.n185 VTAIL.n179 171.744
R1425 VTAIL.n186 VTAIL.n185 171.744
R1426 VTAIL.n186 VTAIL.n175 171.744
R1427 VTAIL.n193 VTAIL.n175 171.744
R1428 VTAIL.n194 VTAIL.n193 171.744
R1429 VTAIL.n194 VTAIL.n171 171.744
R1430 VTAIL.n201 VTAIL.n171 171.744
R1431 VTAIL.n202 VTAIL.n201 171.744
R1432 VTAIL.n202 VTAIL.n167 171.744
R1433 VTAIL.n209 VTAIL.n167 171.744
R1434 VTAIL.n210 VTAIL.n209 171.744
R1435 VTAIL.n210 VTAIL.n163 171.744
R1436 VTAIL.n217 VTAIL.n163 171.744
R1437 VTAIL.n218 VTAIL.n217 171.744
R1438 VTAIL.n218 VTAIL.n159 171.744
R1439 VTAIL.n226 VTAIL.n159 171.744
R1440 VTAIL.n227 VTAIL.n226 171.744
R1441 VTAIL.n228 VTAIL.n227 171.744
R1442 VTAIL.n540 VTAIL.n539 171.744
R1443 VTAIL.n539 VTAIL.n538 171.744
R1444 VTAIL.n538 VTAIL.n471 171.744
R1445 VTAIL.n531 VTAIL.n471 171.744
R1446 VTAIL.n531 VTAIL.n530 171.744
R1447 VTAIL.n530 VTAIL.n476 171.744
R1448 VTAIL.n523 VTAIL.n476 171.744
R1449 VTAIL.n523 VTAIL.n522 171.744
R1450 VTAIL.n522 VTAIL.n480 171.744
R1451 VTAIL.n515 VTAIL.n480 171.744
R1452 VTAIL.n515 VTAIL.n514 171.744
R1453 VTAIL.n514 VTAIL.n484 171.744
R1454 VTAIL.n507 VTAIL.n484 171.744
R1455 VTAIL.n507 VTAIL.n506 171.744
R1456 VTAIL.n506 VTAIL.n488 171.744
R1457 VTAIL.n499 VTAIL.n488 171.744
R1458 VTAIL.n499 VTAIL.n498 171.744
R1459 VTAIL.n498 VTAIL.n492 171.744
R1460 VTAIL.n462 VTAIL.n461 171.744
R1461 VTAIL.n461 VTAIL.n460 171.744
R1462 VTAIL.n460 VTAIL.n393 171.744
R1463 VTAIL.n453 VTAIL.n393 171.744
R1464 VTAIL.n453 VTAIL.n452 171.744
R1465 VTAIL.n452 VTAIL.n398 171.744
R1466 VTAIL.n445 VTAIL.n398 171.744
R1467 VTAIL.n445 VTAIL.n444 171.744
R1468 VTAIL.n444 VTAIL.n402 171.744
R1469 VTAIL.n437 VTAIL.n402 171.744
R1470 VTAIL.n437 VTAIL.n436 171.744
R1471 VTAIL.n436 VTAIL.n406 171.744
R1472 VTAIL.n429 VTAIL.n406 171.744
R1473 VTAIL.n429 VTAIL.n428 171.744
R1474 VTAIL.n428 VTAIL.n410 171.744
R1475 VTAIL.n421 VTAIL.n410 171.744
R1476 VTAIL.n421 VTAIL.n420 171.744
R1477 VTAIL.n420 VTAIL.n414 171.744
R1478 VTAIL.n384 VTAIL.n383 171.744
R1479 VTAIL.n383 VTAIL.n382 171.744
R1480 VTAIL.n382 VTAIL.n315 171.744
R1481 VTAIL.n375 VTAIL.n315 171.744
R1482 VTAIL.n375 VTAIL.n374 171.744
R1483 VTAIL.n374 VTAIL.n320 171.744
R1484 VTAIL.n367 VTAIL.n320 171.744
R1485 VTAIL.n367 VTAIL.n366 171.744
R1486 VTAIL.n366 VTAIL.n324 171.744
R1487 VTAIL.n359 VTAIL.n324 171.744
R1488 VTAIL.n359 VTAIL.n358 171.744
R1489 VTAIL.n358 VTAIL.n328 171.744
R1490 VTAIL.n351 VTAIL.n328 171.744
R1491 VTAIL.n351 VTAIL.n350 171.744
R1492 VTAIL.n350 VTAIL.n332 171.744
R1493 VTAIL.n343 VTAIL.n332 171.744
R1494 VTAIL.n343 VTAIL.n342 171.744
R1495 VTAIL.n342 VTAIL.n336 171.744
R1496 VTAIL.n306 VTAIL.n305 171.744
R1497 VTAIL.n305 VTAIL.n304 171.744
R1498 VTAIL.n304 VTAIL.n237 171.744
R1499 VTAIL.n297 VTAIL.n237 171.744
R1500 VTAIL.n297 VTAIL.n296 171.744
R1501 VTAIL.n296 VTAIL.n242 171.744
R1502 VTAIL.n289 VTAIL.n242 171.744
R1503 VTAIL.n289 VTAIL.n288 171.744
R1504 VTAIL.n288 VTAIL.n246 171.744
R1505 VTAIL.n281 VTAIL.n246 171.744
R1506 VTAIL.n281 VTAIL.n280 171.744
R1507 VTAIL.n280 VTAIL.n250 171.744
R1508 VTAIL.n273 VTAIL.n250 171.744
R1509 VTAIL.n273 VTAIL.n272 171.744
R1510 VTAIL.n272 VTAIL.n254 171.744
R1511 VTAIL.n265 VTAIL.n254 171.744
R1512 VTAIL.n265 VTAIL.n264 171.744
R1513 VTAIL.n264 VTAIL.n258 171.744
R1514 VTAIL.t4 VTAIL.n569 85.8723
R1515 VTAIL.t7 VTAIL.n23 85.8723
R1516 VTAIL.t1 VTAIL.n101 85.8723
R1517 VTAIL.t2 VTAIL.n179 85.8723
R1518 VTAIL.t3 VTAIL.n492 85.8723
R1519 VTAIL.t0 VTAIL.n414 85.8723
R1520 VTAIL.t5 VTAIL.n336 85.8723
R1521 VTAIL.t6 VTAIL.n258 85.8723
R1522 VTAIL.n623 VTAIL.n622 35.8702
R1523 VTAIL.n77 VTAIL.n76 35.8702
R1524 VTAIL.n155 VTAIL.n154 35.8702
R1525 VTAIL.n233 VTAIL.n232 35.8702
R1526 VTAIL.n545 VTAIL.n544 35.8702
R1527 VTAIL.n467 VTAIL.n466 35.8702
R1528 VTAIL.n389 VTAIL.n388 35.8702
R1529 VTAIL.n311 VTAIL.n310 35.8702
R1530 VTAIL.n623 VTAIL.n545 28.0565
R1531 VTAIL.n311 VTAIL.n233 28.0565
R1532 VTAIL.n571 VTAIL.n570 16.3895
R1533 VTAIL.n25 VTAIL.n24 16.3895
R1534 VTAIL.n103 VTAIL.n102 16.3895
R1535 VTAIL.n181 VTAIL.n180 16.3895
R1536 VTAIL.n494 VTAIL.n493 16.3895
R1537 VTAIL.n416 VTAIL.n415 16.3895
R1538 VTAIL.n338 VTAIL.n337 16.3895
R1539 VTAIL.n260 VTAIL.n259 16.3895
R1540 VTAIL.n619 VTAIL.n548 13.1884
R1541 VTAIL.n73 VTAIL.n2 13.1884
R1542 VTAIL.n151 VTAIL.n80 13.1884
R1543 VTAIL.n229 VTAIL.n158 13.1884
R1544 VTAIL.n541 VTAIL.n470 13.1884
R1545 VTAIL.n463 VTAIL.n392 13.1884
R1546 VTAIL.n385 VTAIL.n314 13.1884
R1547 VTAIL.n307 VTAIL.n236 13.1884
R1548 VTAIL.n574 VTAIL.n573 12.8005
R1549 VTAIL.n615 VTAIL.n614 12.8005
R1550 VTAIL.n620 VTAIL.n546 12.8005
R1551 VTAIL.n28 VTAIL.n27 12.8005
R1552 VTAIL.n69 VTAIL.n68 12.8005
R1553 VTAIL.n74 VTAIL.n0 12.8005
R1554 VTAIL.n106 VTAIL.n105 12.8005
R1555 VTAIL.n147 VTAIL.n146 12.8005
R1556 VTAIL.n152 VTAIL.n78 12.8005
R1557 VTAIL.n184 VTAIL.n183 12.8005
R1558 VTAIL.n225 VTAIL.n224 12.8005
R1559 VTAIL.n230 VTAIL.n156 12.8005
R1560 VTAIL.n542 VTAIL.n468 12.8005
R1561 VTAIL.n537 VTAIL.n472 12.8005
R1562 VTAIL.n497 VTAIL.n496 12.8005
R1563 VTAIL.n464 VTAIL.n390 12.8005
R1564 VTAIL.n459 VTAIL.n394 12.8005
R1565 VTAIL.n419 VTAIL.n418 12.8005
R1566 VTAIL.n386 VTAIL.n312 12.8005
R1567 VTAIL.n381 VTAIL.n316 12.8005
R1568 VTAIL.n341 VTAIL.n340 12.8005
R1569 VTAIL.n308 VTAIL.n234 12.8005
R1570 VTAIL.n303 VTAIL.n238 12.8005
R1571 VTAIL.n263 VTAIL.n262 12.8005
R1572 VTAIL.n577 VTAIL.n568 12.0247
R1573 VTAIL.n613 VTAIL.n550 12.0247
R1574 VTAIL.n31 VTAIL.n22 12.0247
R1575 VTAIL.n67 VTAIL.n4 12.0247
R1576 VTAIL.n109 VTAIL.n100 12.0247
R1577 VTAIL.n145 VTAIL.n82 12.0247
R1578 VTAIL.n187 VTAIL.n178 12.0247
R1579 VTAIL.n223 VTAIL.n160 12.0247
R1580 VTAIL.n536 VTAIL.n473 12.0247
R1581 VTAIL.n500 VTAIL.n491 12.0247
R1582 VTAIL.n458 VTAIL.n395 12.0247
R1583 VTAIL.n422 VTAIL.n413 12.0247
R1584 VTAIL.n380 VTAIL.n317 12.0247
R1585 VTAIL.n344 VTAIL.n335 12.0247
R1586 VTAIL.n302 VTAIL.n239 12.0247
R1587 VTAIL.n266 VTAIL.n257 12.0247
R1588 VTAIL.n578 VTAIL.n566 11.249
R1589 VTAIL.n610 VTAIL.n609 11.249
R1590 VTAIL.n32 VTAIL.n20 11.249
R1591 VTAIL.n64 VTAIL.n63 11.249
R1592 VTAIL.n110 VTAIL.n98 11.249
R1593 VTAIL.n142 VTAIL.n141 11.249
R1594 VTAIL.n188 VTAIL.n176 11.249
R1595 VTAIL.n220 VTAIL.n219 11.249
R1596 VTAIL.n533 VTAIL.n532 11.249
R1597 VTAIL.n501 VTAIL.n489 11.249
R1598 VTAIL.n455 VTAIL.n454 11.249
R1599 VTAIL.n423 VTAIL.n411 11.249
R1600 VTAIL.n377 VTAIL.n376 11.249
R1601 VTAIL.n345 VTAIL.n333 11.249
R1602 VTAIL.n299 VTAIL.n298 11.249
R1603 VTAIL.n267 VTAIL.n255 11.249
R1604 VTAIL.n582 VTAIL.n581 10.4732
R1605 VTAIL.n606 VTAIL.n552 10.4732
R1606 VTAIL.n36 VTAIL.n35 10.4732
R1607 VTAIL.n60 VTAIL.n6 10.4732
R1608 VTAIL.n114 VTAIL.n113 10.4732
R1609 VTAIL.n138 VTAIL.n84 10.4732
R1610 VTAIL.n192 VTAIL.n191 10.4732
R1611 VTAIL.n216 VTAIL.n162 10.4732
R1612 VTAIL.n529 VTAIL.n475 10.4732
R1613 VTAIL.n505 VTAIL.n504 10.4732
R1614 VTAIL.n451 VTAIL.n397 10.4732
R1615 VTAIL.n427 VTAIL.n426 10.4732
R1616 VTAIL.n373 VTAIL.n319 10.4732
R1617 VTAIL.n349 VTAIL.n348 10.4732
R1618 VTAIL.n295 VTAIL.n241 10.4732
R1619 VTAIL.n271 VTAIL.n270 10.4732
R1620 VTAIL.n585 VTAIL.n564 9.69747
R1621 VTAIL.n605 VTAIL.n554 9.69747
R1622 VTAIL.n39 VTAIL.n18 9.69747
R1623 VTAIL.n59 VTAIL.n8 9.69747
R1624 VTAIL.n117 VTAIL.n96 9.69747
R1625 VTAIL.n137 VTAIL.n86 9.69747
R1626 VTAIL.n195 VTAIL.n174 9.69747
R1627 VTAIL.n215 VTAIL.n164 9.69747
R1628 VTAIL.n528 VTAIL.n477 9.69747
R1629 VTAIL.n508 VTAIL.n487 9.69747
R1630 VTAIL.n450 VTAIL.n399 9.69747
R1631 VTAIL.n430 VTAIL.n409 9.69747
R1632 VTAIL.n372 VTAIL.n321 9.69747
R1633 VTAIL.n352 VTAIL.n331 9.69747
R1634 VTAIL.n294 VTAIL.n243 9.69747
R1635 VTAIL.n274 VTAIL.n253 9.69747
R1636 VTAIL.n622 VTAIL.n621 9.45567
R1637 VTAIL.n76 VTAIL.n75 9.45567
R1638 VTAIL.n154 VTAIL.n153 9.45567
R1639 VTAIL.n232 VTAIL.n231 9.45567
R1640 VTAIL.n544 VTAIL.n543 9.45567
R1641 VTAIL.n466 VTAIL.n465 9.45567
R1642 VTAIL.n388 VTAIL.n387 9.45567
R1643 VTAIL.n310 VTAIL.n309 9.45567
R1644 VTAIL.n621 VTAIL.n620 9.3005
R1645 VTAIL.n560 VTAIL.n559 9.3005
R1646 VTAIL.n589 VTAIL.n588 9.3005
R1647 VTAIL.n587 VTAIL.n586 9.3005
R1648 VTAIL.n564 VTAIL.n563 9.3005
R1649 VTAIL.n581 VTAIL.n580 9.3005
R1650 VTAIL.n579 VTAIL.n578 9.3005
R1651 VTAIL.n568 VTAIL.n567 9.3005
R1652 VTAIL.n573 VTAIL.n572 9.3005
R1653 VTAIL.n595 VTAIL.n594 9.3005
R1654 VTAIL.n597 VTAIL.n596 9.3005
R1655 VTAIL.n556 VTAIL.n555 9.3005
R1656 VTAIL.n603 VTAIL.n602 9.3005
R1657 VTAIL.n605 VTAIL.n604 9.3005
R1658 VTAIL.n552 VTAIL.n551 9.3005
R1659 VTAIL.n611 VTAIL.n610 9.3005
R1660 VTAIL.n613 VTAIL.n612 9.3005
R1661 VTAIL.n614 VTAIL.n547 9.3005
R1662 VTAIL.n75 VTAIL.n74 9.3005
R1663 VTAIL.n14 VTAIL.n13 9.3005
R1664 VTAIL.n43 VTAIL.n42 9.3005
R1665 VTAIL.n41 VTAIL.n40 9.3005
R1666 VTAIL.n18 VTAIL.n17 9.3005
R1667 VTAIL.n35 VTAIL.n34 9.3005
R1668 VTAIL.n33 VTAIL.n32 9.3005
R1669 VTAIL.n22 VTAIL.n21 9.3005
R1670 VTAIL.n27 VTAIL.n26 9.3005
R1671 VTAIL.n49 VTAIL.n48 9.3005
R1672 VTAIL.n51 VTAIL.n50 9.3005
R1673 VTAIL.n10 VTAIL.n9 9.3005
R1674 VTAIL.n57 VTAIL.n56 9.3005
R1675 VTAIL.n59 VTAIL.n58 9.3005
R1676 VTAIL.n6 VTAIL.n5 9.3005
R1677 VTAIL.n65 VTAIL.n64 9.3005
R1678 VTAIL.n67 VTAIL.n66 9.3005
R1679 VTAIL.n68 VTAIL.n1 9.3005
R1680 VTAIL.n153 VTAIL.n152 9.3005
R1681 VTAIL.n92 VTAIL.n91 9.3005
R1682 VTAIL.n121 VTAIL.n120 9.3005
R1683 VTAIL.n119 VTAIL.n118 9.3005
R1684 VTAIL.n96 VTAIL.n95 9.3005
R1685 VTAIL.n113 VTAIL.n112 9.3005
R1686 VTAIL.n111 VTAIL.n110 9.3005
R1687 VTAIL.n100 VTAIL.n99 9.3005
R1688 VTAIL.n105 VTAIL.n104 9.3005
R1689 VTAIL.n127 VTAIL.n126 9.3005
R1690 VTAIL.n129 VTAIL.n128 9.3005
R1691 VTAIL.n88 VTAIL.n87 9.3005
R1692 VTAIL.n135 VTAIL.n134 9.3005
R1693 VTAIL.n137 VTAIL.n136 9.3005
R1694 VTAIL.n84 VTAIL.n83 9.3005
R1695 VTAIL.n143 VTAIL.n142 9.3005
R1696 VTAIL.n145 VTAIL.n144 9.3005
R1697 VTAIL.n146 VTAIL.n79 9.3005
R1698 VTAIL.n231 VTAIL.n230 9.3005
R1699 VTAIL.n170 VTAIL.n169 9.3005
R1700 VTAIL.n199 VTAIL.n198 9.3005
R1701 VTAIL.n197 VTAIL.n196 9.3005
R1702 VTAIL.n174 VTAIL.n173 9.3005
R1703 VTAIL.n191 VTAIL.n190 9.3005
R1704 VTAIL.n189 VTAIL.n188 9.3005
R1705 VTAIL.n178 VTAIL.n177 9.3005
R1706 VTAIL.n183 VTAIL.n182 9.3005
R1707 VTAIL.n205 VTAIL.n204 9.3005
R1708 VTAIL.n207 VTAIL.n206 9.3005
R1709 VTAIL.n166 VTAIL.n165 9.3005
R1710 VTAIL.n213 VTAIL.n212 9.3005
R1711 VTAIL.n215 VTAIL.n214 9.3005
R1712 VTAIL.n162 VTAIL.n161 9.3005
R1713 VTAIL.n221 VTAIL.n220 9.3005
R1714 VTAIL.n223 VTAIL.n222 9.3005
R1715 VTAIL.n224 VTAIL.n157 9.3005
R1716 VTAIL.n520 VTAIL.n519 9.3005
R1717 VTAIL.n479 VTAIL.n478 9.3005
R1718 VTAIL.n526 VTAIL.n525 9.3005
R1719 VTAIL.n528 VTAIL.n527 9.3005
R1720 VTAIL.n475 VTAIL.n474 9.3005
R1721 VTAIL.n534 VTAIL.n533 9.3005
R1722 VTAIL.n536 VTAIL.n535 9.3005
R1723 VTAIL.n472 VTAIL.n469 9.3005
R1724 VTAIL.n543 VTAIL.n542 9.3005
R1725 VTAIL.n518 VTAIL.n517 9.3005
R1726 VTAIL.n483 VTAIL.n482 9.3005
R1727 VTAIL.n512 VTAIL.n511 9.3005
R1728 VTAIL.n510 VTAIL.n509 9.3005
R1729 VTAIL.n487 VTAIL.n486 9.3005
R1730 VTAIL.n504 VTAIL.n503 9.3005
R1731 VTAIL.n502 VTAIL.n501 9.3005
R1732 VTAIL.n491 VTAIL.n490 9.3005
R1733 VTAIL.n496 VTAIL.n495 9.3005
R1734 VTAIL.n442 VTAIL.n441 9.3005
R1735 VTAIL.n401 VTAIL.n400 9.3005
R1736 VTAIL.n448 VTAIL.n447 9.3005
R1737 VTAIL.n450 VTAIL.n449 9.3005
R1738 VTAIL.n397 VTAIL.n396 9.3005
R1739 VTAIL.n456 VTAIL.n455 9.3005
R1740 VTAIL.n458 VTAIL.n457 9.3005
R1741 VTAIL.n394 VTAIL.n391 9.3005
R1742 VTAIL.n465 VTAIL.n464 9.3005
R1743 VTAIL.n440 VTAIL.n439 9.3005
R1744 VTAIL.n405 VTAIL.n404 9.3005
R1745 VTAIL.n434 VTAIL.n433 9.3005
R1746 VTAIL.n432 VTAIL.n431 9.3005
R1747 VTAIL.n409 VTAIL.n408 9.3005
R1748 VTAIL.n426 VTAIL.n425 9.3005
R1749 VTAIL.n424 VTAIL.n423 9.3005
R1750 VTAIL.n413 VTAIL.n412 9.3005
R1751 VTAIL.n418 VTAIL.n417 9.3005
R1752 VTAIL.n364 VTAIL.n363 9.3005
R1753 VTAIL.n323 VTAIL.n322 9.3005
R1754 VTAIL.n370 VTAIL.n369 9.3005
R1755 VTAIL.n372 VTAIL.n371 9.3005
R1756 VTAIL.n319 VTAIL.n318 9.3005
R1757 VTAIL.n378 VTAIL.n377 9.3005
R1758 VTAIL.n380 VTAIL.n379 9.3005
R1759 VTAIL.n316 VTAIL.n313 9.3005
R1760 VTAIL.n387 VTAIL.n386 9.3005
R1761 VTAIL.n362 VTAIL.n361 9.3005
R1762 VTAIL.n327 VTAIL.n326 9.3005
R1763 VTAIL.n356 VTAIL.n355 9.3005
R1764 VTAIL.n354 VTAIL.n353 9.3005
R1765 VTAIL.n331 VTAIL.n330 9.3005
R1766 VTAIL.n348 VTAIL.n347 9.3005
R1767 VTAIL.n346 VTAIL.n345 9.3005
R1768 VTAIL.n335 VTAIL.n334 9.3005
R1769 VTAIL.n340 VTAIL.n339 9.3005
R1770 VTAIL.n286 VTAIL.n285 9.3005
R1771 VTAIL.n245 VTAIL.n244 9.3005
R1772 VTAIL.n292 VTAIL.n291 9.3005
R1773 VTAIL.n294 VTAIL.n293 9.3005
R1774 VTAIL.n241 VTAIL.n240 9.3005
R1775 VTAIL.n300 VTAIL.n299 9.3005
R1776 VTAIL.n302 VTAIL.n301 9.3005
R1777 VTAIL.n238 VTAIL.n235 9.3005
R1778 VTAIL.n309 VTAIL.n308 9.3005
R1779 VTAIL.n284 VTAIL.n283 9.3005
R1780 VTAIL.n249 VTAIL.n248 9.3005
R1781 VTAIL.n278 VTAIL.n277 9.3005
R1782 VTAIL.n276 VTAIL.n275 9.3005
R1783 VTAIL.n253 VTAIL.n252 9.3005
R1784 VTAIL.n270 VTAIL.n269 9.3005
R1785 VTAIL.n268 VTAIL.n267 9.3005
R1786 VTAIL.n257 VTAIL.n256 9.3005
R1787 VTAIL.n262 VTAIL.n261 9.3005
R1788 VTAIL.n586 VTAIL.n562 8.92171
R1789 VTAIL.n602 VTAIL.n601 8.92171
R1790 VTAIL.n40 VTAIL.n16 8.92171
R1791 VTAIL.n56 VTAIL.n55 8.92171
R1792 VTAIL.n118 VTAIL.n94 8.92171
R1793 VTAIL.n134 VTAIL.n133 8.92171
R1794 VTAIL.n196 VTAIL.n172 8.92171
R1795 VTAIL.n212 VTAIL.n211 8.92171
R1796 VTAIL.n525 VTAIL.n524 8.92171
R1797 VTAIL.n509 VTAIL.n485 8.92171
R1798 VTAIL.n447 VTAIL.n446 8.92171
R1799 VTAIL.n431 VTAIL.n407 8.92171
R1800 VTAIL.n369 VTAIL.n368 8.92171
R1801 VTAIL.n353 VTAIL.n329 8.92171
R1802 VTAIL.n291 VTAIL.n290 8.92171
R1803 VTAIL.n275 VTAIL.n251 8.92171
R1804 VTAIL.n590 VTAIL.n589 8.14595
R1805 VTAIL.n598 VTAIL.n556 8.14595
R1806 VTAIL.n44 VTAIL.n43 8.14595
R1807 VTAIL.n52 VTAIL.n10 8.14595
R1808 VTAIL.n122 VTAIL.n121 8.14595
R1809 VTAIL.n130 VTAIL.n88 8.14595
R1810 VTAIL.n200 VTAIL.n199 8.14595
R1811 VTAIL.n208 VTAIL.n166 8.14595
R1812 VTAIL.n521 VTAIL.n479 8.14595
R1813 VTAIL.n513 VTAIL.n512 8.14595
R1814 VTAIL.n443 VTAIL.n401 8.14595
R1815 VTAIL.n435 VTAIL.n434 8.14595
R1816 VTAIL.n365 VTAIL.n323 8.14595
R1817 VTAIL.n357 VTAIL.n356 8.14595
R1818 VTAIL.n287 VTAIL.n245 8.14595
R1819 VTAIL.n279 VTAIL.n278 8.14595
R1820 VTAIL.n593 VTAIL.n560 7.3702
R1821 VTAIL.n597 VTAIL.n558 7.3702
R1822 VTAIL.n47 VTAIL.n14 7.3702
R1823 VTAIL.n51 VTAIL.n12 7.3702
R1824 VTAIL.n125 VTAIL.n92 7.3702
R1825 VTAIL.n129 VTAIL.n90 7.3702
R1826 VTAIL.n203 VTAIL.n170 7.3702
R1827 VTAIL.n207 VTAIL.n168 7.3702
R1828 VTAIL.n520 VTAIL.n481 7.3702
R1829 VTAIL.n516 VTAIL.n483 7.3702
R1830 VTAIL.n442 VTAIL.n403 7.3702
R1831 VTAIL.n438 VTAIL.n405 7.3702
R1832 VTAIL.n364 VTAIL.n325 7.3702
R1833 VTAIL.n360 VTAIL.n327 7.3702
R1834 VTAIL.n286 VTAIL.n247 7.3702
R1835 VTAIL.n282 VTAIL.n249 7.3702
R1836 VTAIL.n594 VTAIL.n593 6.59444
R1837 VTAIL.n594 VTAIL.n558 6.59444
R1838 VTAIL.n48 VTAIL.n47 6.59444
R1839 VTAIL.n48 VTAIL.n12 6.59444
R1840 VTAIL.n126 VTAIL.n125 6.59444
R1841 VTAIL.n126 VTAIL.n90 6.59444
R1842 VTAIL.n204 VTAIL.n203 6.59444
R1843 VTAIL.n204 VTAIL.n168 6.59444
R1844 VTAIL.n517 VTAIL.n481 6.59444
R1845 VTAIL.n517 VTAIL.n516 6.59444
R1846 VTAIL.n439 VTAIL.n403 6.59444
R1847 VTAIL.n439 VTAIL.n438 6.59444
R1848 VTAIL.n361 VTAIL.n325 6.59444
R1849 VTAIL.n361 VTAIL.n360 6.59444
R1850 VTAIL.n283 VTAIL.n247 6.59444
R1851 VTAIL.n283 VTAIL.n282 6.59444
R1852 VTAIL.n590 VTAIL.n560 5.81868
R1853 VTAIL.n598 VTAIL.n597 5.81868
R1854 VTAIL.n44 VTAIL.n14 5.81868
R1855 VTAIL.n52 VTAIL.n51 5.81868
R1856 VTAIL.n122 VTAIL.n92 5.81868
R1857 VTAIL.n130 VTAIL.n129 5.81868
R1858 VTAIL.n200 VTAIL.n170 5.81868
R1859 VTAIL.n208 VTAIL.n207 5.81868
R1860 VTAIL.n521 VTAIL.n520 5.81868
R1861 VTAIL.n513 VTAIL.n483 5.81868
R1862 VTAIL.n443 VTAIL.n442 5.81868
R1863 VTAIL.n435 VTAIL.n405 5.81868
R1864 VTAIL.n365 VTAIL.n364 5.81868
R1865 VTAIL.n357 VTAIL.n327 5.81868
R1866 VTAIL.n287 VTAIL.n286 5.81868
R1867 VTAIL.n279 VTAIL.n249 5.81868
R1868 VTAIL.n589 VTAIL.n562 5.04292
R1869 VTAIL.n601 VTAIL.n556 5.04292
R1870 VTAIL.n43 VTAIL.n16 5.04292
R1871 VTAIL.n55 VTAIL.n10 5.04292
R1872 VTAIL.n121 VTAIL.n94 5.04292
R1873 VTAIL.n133 VTAIL.n88 5.04292
R1874 VTAIL.n199 VTAIL.n172 5.04292
R1875 VTAIL.n211 VTAIL.n166 5.04292
R1876 VTAIL.n524 VTAIL.n479 5.04292
R1877 VTAIL.n512 VTAIL.n485 5.04292
R1878 VTAIL.n446 VTAIL.n401 5.04292
R1879 VTAIL.n434 VTAIL.n407 5.04292
R1880 VTAIL.n368 VTAIL.n323 5.04292
R1881 VTAIL.n356 VTAIL.n329 5.04292
R1882 VTAIL.n290 VTAIL.n245 5.04292
R1883 VTAIL.n278 VTAIL.n251 5.04292
R1884 VTAIL.n586 VTAIL.n585 4.26717
R1885 VTAIL.n602 VTAIL.n554 4.26717
R1886 VTAIL.n40 VTAIL.n39 4.26717
R1887 VTAIL.n56 VTAIL.n8 4.26717
R1888 VTAIL.n118 VTAIL.n117 4.26717
R1889 VTAIL.n134 VTAIL.n86 4.26717
R1890 VTAIL.n196 VTAIL.n195 4.26717
R1891 VTAIL.n212 VTAIL.n164 4.26717
R1892 VTAIL.n525 VTAIL.n477 4.26717
R1893 VTAIL.n509 VTAIL.n508 4.26717
R1894 VTAIL.n447 VTAIL.n399 4.26717
R1895 VTAIL.n431 VTAIL.n430 4.26717
R1896 VTAIL.n369 VTAIL.n321 4.26717
R1897 VTAIL.n353 VTAIL.n352 4.26717
R1898 VTAIL.n291 VTAIL.n243 4.26717
R1899 VTAIL.n275 VTAIL.n274 4.26717
R1900 VTAIL.n572 VTAIL.n571 3.70982
R1901 VTAIL.n26 VTAIL.n25 3.70982
R1902 VTAIL.n104 VTAIL.n103 3.70982
R1903 VTAIL.n182 VTAIL.n181 3.70982
R1904 VTAIL.n495 VTAIL.n494 3.70982
R1905 VTAIL.n417 VTAIL.n416 3.70982
R1906 VTAIL.n339 VTAIL.n338 3.70982
R1907 VTAIL.n261 VTAIL.n260 3.70982
R1908 VTAIL.n389 VTAIL.n311 3.52636
R1909 VTAIL.n545 VTAIL.n467 3.52636
R1910 VTAIL.n233 VTAIL.n155 3.52636
R1911 VTAIL.n582 VTAIL.n564 3.49141
R1912 VTAIL.n606 VTAIL.n605 3.49141
R1913 VTAIL.n36 VTAIL.n18 3.49141
R1914 VTAIL.n60 VTAIL.n59 3.49141
R1915 VTAIL.n114 VTAIL.n96 3.49141
R1916 VTAIL.n138 VTAIL.n137 3.49141
R1917 VTAIL.n192 VTAIL.n174 3.49141
R1918 VTAIL.n216 VTAIL.n215 3.49141
R1919 VTAIL.n529 VTAIL.n528 3.49141
R1920 VTAIL.n505 VTAIL.n487 3.49141
R1921 VTAIL.n451 VTAIL.n450 3.49141
R1922 VTAIL.n427 VTAIL.n409 3.49141
R1923 VTAIL.n373 VTAIL.n372 3.49141
R1924 VTAIL.n349 VTAIL.n331 3.49141
R1925 VTAIL.n295 VTAIL.n294 3.49141
R1926 VTAIL.n271 VTAIL.n253 3.49141
R1927 VTAIL.n581 VTAIL.n566 2.71565
R1928 VTAIL.n609 VTAIL.n552 2.71565
R1929 VTAIL.n35 VTAIL.n20 2.71565
R1930 VTAIL.n63 VTAIL.n6 2.71565
R1931 VTAIL.n113 VTAIL.n98 2.71565
R1932 VTAIL.n141 VTAIL.n84 2.71565
R1933 VTAIL.n191 VTAIL.n176 2.71565
R1934 VTAIL.n219 VTAIL.n162 2.71565
R1935 VTAIL.n532 VTAIL.n475 2.71565
R1936 VTAIL.n504 VTAIL.n489 2.71565
R1937 VTAIL.n454 VTAIL.n397 2.71565
R1938 VTAIL.n426 VTAIL.n411 2.71565
R1939 VTAIL.n376 VTAIL.n319 2.71565
R1940 VTAIL.n348 VTAIL.n333 2.71565
R1941 VTAIL.n298 VTAIL.n241 2.71565
R1942 VTAIL.n270 VTAIL.n255 2.71565
R1943 VTAIL.n578 VTAIL.n577 1.93989
R1944 VTAIL.n610 VTAIL.n550 1.93989
R1945 VTAIL.n32 VTAIL.n31 1.93989
R1946 VTAIL.n64 VTAIL.n4 1.93989
R1947 VTAIL.n110 VTAIL.n109 1.93989
R1948 VTAIL.n142 VTAIL.n82 1.93989
R1949 VTAIL.n188 VTAIL.n187 1.93989
R1950 VTAIL.n220 VTAIL.n160 1.93989
R1951 VTAIL.n533 VTAIL.n473 1.93989
R1952 VTAIL.n501 VTAIL.n500 1.93989
R1953 VTAIL.n455 VTAIL.n395 1.93989
R1954 VTAIL.n423 VTAIL.n422 1.93989
R1955 VTAIL.n377 VTAIL.n317 1.93989
R1956 VTAIL.n345 VTAIL.n344 1.93989
R1957 VTAIL.n299 VTAIL.n239 1.93989
R1958 VTAIL.n267 VTAIL.n266 1.93989
R1959 VTAIL VTAIL.n77 1.82162
R1960 VTAIL VTAIL.n623 1.70524
R1961 VTAIL.n574 VTAIL.n568 1.16414
R1962 VTAIL.n615 VTAIL.n613 1.16414
R1963 VTAIL.n622 VTAIL.n546 1.16414
R1964 VTAIL.n28 VTAIL.n22 1.16414
R1965 VTAIL.n69 VTAIL.n67 1.16414
R1966 VTAIL.n76 VTAIL.n0 1.16414
R1967 VTAIL.n106 VTAIL.n100 1.16414
R1968 VTAIL.n147 VTAIL.n145 1.16414
R1969 VTAIL.n154 VTAIL.n78 1.16414
R1970 VTAIL.n184 VTAIL.n178 1.16414
R1971 VTAIL.n225 VTAIL.n223 1.16414
R1972 VTAIL.n232 VTAIL.n156 1.16414
R1973 VTAIL.n544 VTAIL.n468 1.16414
R1974 VTAIL.n537 VTAIL.n536 1.16414
R1975 VTAIL.n497 VTAIL.n491 1.16414
R1976 VTAIL.n466 VTAIL.n390 1.16414
R1977 VTAIL.n459 VTAIL.n458 1.16414
R1978 VTAIL.n419 VTAIL.n413 1.16414
R1979 VTAIL.n388 VTAIL.n312 1.16414
R1980 VTAIL.n381 VTAIL.n380 1.16414
R1981 VTAIL.n341 VTAIL.n335 1.16414
R1982 VTAIL.n310 VTAIL.n234 1.16414
R1983 VTAIL.n303 VTAIL.n302 1.16414
R1984 VTAIL.n263 VTAIL.n257 1.16414
R1985 VTAIL.n467 VTAIL.n389 0.470328
R1986 VTAIL.n155 VTAIL.n77 0.470328
R1987 VTAIL.n573 VTAIL.n570 0.388379
R1988 VTAIL.n614 VTAIL.n548 0.388379
R1989 VTAIL.n620 VTAIL.n619 0.388379
R1990 VTAIL.n27 VTAIL.n24 0.388379
R1991 VTAIL.n68 VTAIL.n2 0.388379
R1992 VTAIL.n74 VTAIL.n73 0.388379
R1993 VTAIL.n105 VTAIL.n102 0.388379
R1994 VTAIL.n146 VTAIL.n80 0.388379
R1995 VTAIL.n152 VTAIL.n151 0.388379
R1996 VTAIL.n183 VTAIL.n180 0.388379
R1997 VTAIL.n224 VTAIL.n158 0.388379
R1998 VTAIL.n230 VTAIL.n229 0.388379
R1999 VTAIL.n542 VTAIL.n541 0.388379
R2000 VTAIL.n472 VTAIL.n470 0.388379
R2001 VTAIL.n496 VTAIL.n493 0.388379
R2002 VTAIL.n464 VTAIL.n463 0.388379
R2003 VTAIL.n394 VTAIL.n392 0.388379
R2004 VTAIL.n418 VTAIL.n415 0.388379
R2005 VTAIL.n386 VTAIL.n385 0.388379
R2006 VTAIL.n316 VTAIL.n314 0.388379
R2007 VTAIL.n340 VTAIL.n337 0.388379
R2008 VTAIL.n308 VTAIL.n307 0.388379
R2009 VTAIL.n238 VTAIL.n236 0.388379
R2010 VTAIL.n262 VTAIL.n259 0.388379
R2011 VTAIL.n572 VTAIL.n567 0.155672
R2012 VTAIL.n579 VTAIL.n567 0.155672
R2013 VTAIL.n580 VTAIL.n579 0.155672
R2014 VTAIL.n580 VTAIL.n563 0.155672
R2015 VTAIL.n587 VTAIL.n563 0.155672
R2016 VTAIL.n588 VTAIL.n587 0.155672
R2017 VTAIL.n588 VTAIL.n559 0.155672
R2018 VTAIL.n595 VTAIL.n559 0.155672
R2019 VTAIL.n596 VTAIL.n595 0.155672
R2020 VTAIL.n596 VTAIL.n555 0.155672
R2021 VTAIL.n603 VTAIL.n555 0.155672
R2022 VTAIL.n604 VTAIL.n603 0.155672
R2023 VTAIL.n604 VTAIL.n551 0.155672
R2024 VTAIL.n611 VTAIL.n551 0.155672
R2025 VTAIL.n612 VTAIL.n611 0.155672
R2026 VTAIL.n612 VTAIL.n547 0.155672
R2027 VTAIL.n621 VTAIL.n547 0.155672
R2028 VTAIL.n26 VTAIL.n21 0.155672
R2029 VTAIL.n33 VTAIL.n21 0.155672
R2030 VTAIL.n34 VTAIL.n33 0.155672
R2031 VTAIL.n34 VTAIL.n17 0.155672
R2032 VTAIL.n41 VTAIL.n17 0.155672
R2033 VTAIL.n42 VTAIL.n41 0.155672
R2034 VTAIL.n42 VTAIL.n13 0.155672
R2035 VTAIL.n49 VTAIL.n13 0.155672
R2036 VTAIL.n50 VTAIL.n49 0.155672
R2037 VTAIL.n50 VTAIL.n9 0.155672
R2038 VTAIL.n57 VTAIL.n9 0.155672
R2039 VTAIL.n58 VTAIL.n57 0.155672
R2040 VTAIL.n58 VTAIL.n5 0.155672
R2041 VTAIL.n65 VTAIL.n5 0.155672
R2042 VTAIL.n66 VTAIL.n65 0.155672
R2043 VTAIL.n66 VTAIL.n1 0.155672
R2044 VTAIL.n75 VTAIL.n1 0.155672
R2045 VTAIL.n104 VTAIL.n99 0.155672
R2046 VTAIL.n111 VTAIL.n99 0.155672
R2047 VTAIL.n112 VTAIL.n111 0.155672
R2048 VTAIL.n112 VTAIL.n95 0.155672
R2049 VTAIL.n119 VTAIL.n95 0.155672
R2050 VTAIL.n120 VTAIL.n119 0.155672
R2051 VTAIL.n120 VTAIL.n91 0.155672
R2052 VTAIL.n127 VTAIL.n91 0.155672
R2053 VTAIL.n128 VTAIL.n127 0.155672
R2054 VTAIL.n128 VTAIL.n87 0.155672
R2055 VTAIL.n135 VTAIL.n87 0.155672
R2056 VTAIL.n136 VTAIL.n135 0.155672
R2057 VTAIL.n136 VTAIL.n83 0.155672
R2058 VTAIL.n143 VTAIL.n83 0.155672
R2059 VTAIL.n144 VTAIL.n143 0.155672
R2060 VTAIL.n144 VTAIL.n79 0.155672
R2061 VTAIL.n153 VTAIL.n79 0.155672
R2062 VTAIL.n182 VTAIL.n177 0.155672
R2063 VTAIL.n189 VTAIL.n177 0.155672
R2064 VTAIL.n190 VTAIL.n189 0.155672
R2065 VTAIL.n190 VTAIL.n173 0.155672
R2066 VTAIL.n197 VTAIL.n173 0.155672
R2067 VTAIL.n198 VTAIL.n197 0.155672
R2068 VTAIL.n198 VTAIL.n169 0.155672
R2069 VTAIL.n205 VTAIL.n169 0.155672
R2070 VTAIL.n206 VTAIL.n205 0.155672
R2071 VTAIL.n206 VTAIL.n165 0.155672
R2072 VTAIL.n213 VTAIL.n165 0.155672
R2073 VTAIL.n214 VTAIL.n213 0.155672
R2074 VTAIL.n214 VTAIL.n161 0.155672
R2075 VTAIL.n221 VTAIL.n161 0.155672
R2076 VTAIL.n222 VTAIL.n221 0.155672
R2077 VTAIL.n222 VTAIL.n157 0.155672
R2078 VTAIL.n231 VTAIL.n157 0.155672
R2079 VTAIL.n543 VTAIL.n469 0.155672
R2080 VTAIL.n535 VTAIL.n469 0.155672
R2081 VTAIL.n535 VTAIL.n534 0.155672
R2082 VTAIL.n534 VTAIL.n474 0.155672
R2083 VTAIL.n527 VTAIL.n474 0.155672
R2084 VTAIL.n527 VTAIL.n526 0.155672
R2085 VTAIL.n526 VTAIL.n478 0.155672
R2086 VTAIL.n519 VTAIL.n478 0.155672
R2087 VTAIL.n519 VTAIL.n518 0.155672
R2088 VTAIL.n518 VTAIL.n482 0.155672
R2089 VTAIL.n511 VTAIL.n482 0.155672
R2090 VTAIL.n511 VTAIL.n510 0.155672
R2091 VTAIL.n510 VTAIL.n486 0.155672
R2092 VTAIL.n503 VTAIL.n486 0.155672
R2093 VTAIL.n503 VTAIL.n502 0.155672
R2094 VTAIL.n502 VTAIL.n490 0.155672
R2095 VTAIL.n495 VTAIL.n490 0.155672
R2096 VTAIL.n465 VTAIL.n391 0.155672
R2097 VTAIL.n457 VTAIL.n391 0.155672
R2098 VTAIL.n457 VTAIL.n456 0.155672
R2099 VTAIL.n456 VTAIL.n396 0.155672
R2100 VTAIL.n449 VTAIL.n396 0.155672
R2101 VTAIL.n449 VTAIL.n448 0.155672
R2102 VTAIL.n448 VTAIL.n400 0.155672
R2103 VTAIL.n441 VTAIL.n400 0.155672
R2104 VTAIL.n441 VTAIL.n440 0.155672
R2105 VTAIL.n440 VTAIL.n404 0.155672
R2106 VTAIL.n433 VTAIL.n404 0.155672
R2107 VTAIL.n433 VTAIL.n432 0.155672
R2108 VTAIL.n432 VTAIL.n408 0.155672
R2109 VTAIL.n425 VTAIL.n408 0.155672
R2110 VTAIL.n425 VTAIL.n424 0.155672
R2111 VTAIL.n424 VTAIL.n412 0.155672
R2112 VTAIL.n417 VTAIL.n412 0.155672
R2113 VTAIL.n387 VTAIL.n313 0.155672
R2114 VTAIL.n379 VTAIL.n313 0.155672
R2115 VTAIL.n379 VTAIL.n378 0.155672
R2116 VTAIL.n378 VTAIL.n318 0.155672
R2117 VTAIL.n371 VTAIL.n318 0.155672
R2118 VTAIL.n371 VTAIL.n370 0.155672
R2119 VTAIL.n370 VTAIL.n322 0.155672
R2120 VTAIL.n363 VTAIL.n322 0.155672
R2121 VTAIL.n363 VTAIL.n362 0.155672
R2122 VTAIL.n362 VTAIL.n326 0.155672
R2123 VTAIL.n355 VTAIL.n326 0.155672
R2124 VTAIL.n355 VTAIL.n354 0.155672
R2125 VTAIL.n354 VTAIL.n330 0.155672
R2126 VTAIL.n347 VTAIL.n330 0.155672
R2127 VTAIL.n347 VTAIL.n346 0.155672
R2128 VTAIL.n346 VTAIL.n334 0.155672
R2129 VTAIL.n339 VTAIL.n334 0.155672
R2130 VTAIL.n309 VTAIL.n235 0.155672
R2131 VTAIL.n301 VTAIL.n235 0.155672
R2132 VTAIL.n301 VTAIL.n300 0.155672
R2133 VTAIL.n300 VTAIL.n240 0.155672
R2134 VTAIL.n293 VTAIL.n240 0.155672
R2135 VTAIL.n293 VTAIL.n292 0.155672
R2136 VTAIL.n292 VTAIL.n244 0.155672
R2137 VTAIL.n285 VTAIL.n244 0.155672
R2138 VTAIL.n285 VTAIL.n284 0.155672
R2139 VTAIL.n284 VTAIL.n248 0.155672
R2140 VTAIL.n277 VTAIL.n248 0.155672
R2141 VTAIL.n277 VTAIL.n276 0.155672
R2142 VTAIL.n276 VTAIL.n252 0.155672
R2143 VTAIL.n269 VTAIL.n252 0.155672
R2144 VTAIL.n269 VTAIL.n268 0.155672
R2145 VTAIL.n268 VTAIL.n256 0.155672
R2146 VTAIL.n261 VTAIL.n256 0.155672
R2147 VP.n21 VP.n20 161.3
R2148 VP.n19 VP.n1 161.3
R2149 VP.n18 VP.n17 161.3
R2150 VP.n16 VP.n2 161.3
R2151 VP.n15 VP.n14 161.3
R2152 VP.n13 VP.n3 161.3
R2153 VP.n12 VP.n11 161.3
R2154 VP.n10 VP.n4 161.3
R2155 VP.n9 VP.n8 161.3
R2156 VP.n5 VP.t1 124.124
R2157 VP.n5 VP.t0 122.784
R2158 VP.n7 VP.t3 90.4396
R2159 VP.n0 VP.t2 90.4396
R2160 VP.n7 VP.n6 87.8654
R2161 VP.n22 VP.n0 87.8654
R2162 VP.n6 VP.n5 53.3786
R2163 VP.n14 VP.n13 40.4934
R2164 VP.n14 VP.n2 40.4934
R2165 VP.n8 VP.n4 24.4675
R2166 VP.n12 VP.n4 24.4675
R2167 VP.n13 VP.n12 24.4675
R2168 VP.n18 VP.n2 24.4675
R2169 VP.n19 VP.n18 24.4675
R2170 VP.n20 VP.n19 24.4675
R2171 VP.n8 VP.n7 2.20253
R2172 VP.n20 VP.n0 2.20253
R2173 VP.n9 VP.n6 0.354971
R2174 VP.n22 VP.n21 0.354971
R2175 VP VP.n22 0.26696
R2176 VP.n10 VP.n9 0.189894
R2177 VP.n11 VP.n10 0.189894
R2178 VP.n11 VP.n3 0.189894
R2179 VP.n15 VP.n3 0.189894
R2180 VP.n16 VP.n15 0.189894
R2181 VP.n17 VP.n16 0.189894
R2182 VP.n17 VP.n1 0.189894
R2183 VP.n21 VP.n1 0.189894
R2184 VDD1 VDD1.n1 121.999
R2185 VDD1 VDD1.n0 75.0772
R2186 VDD1.n0 VDD1.t2 2.30419
R2187 VDD1.n0 VDD1.t3 2.30419
R2188 VDD1.n1 VDD1.t0 2.30419
R2189 VDD1.n1 VDD1.t1 2.30419
C0 B w_n3424_n3790# 11.2638f
C1 VP w_n3424_n3790# 6.50131f
C2 VTAIL w_n3424_n3790# 4.46922f
C3 VP B 2.09422f
C4 VN w_n3424_n3790# 6.05821f
C5 VDD1 w_n3424_n3790# 1.72376f
C6 VTAIL B 6.14329f
C7 VDD2 w_n3424_n3790# 1.80545f
C8 VN B 1.35352f
C9 VDD1 B 1.52419f
C10 VTAIL VP 5.84745f
C11 VDD2 B 1.59554f
C12 VN VP 7.41952f
C13 VDD1 VP 6.17304f
C14 VDD2 VP 0.467972f
C15 VN VTAIL 5.83334f
C16 VDD1 VTAIL 6.17396f
C17 VDD1 VN 0.149902f
C18 VDD2 VTAIL 6.23594f
C19 VN VDD2 5.856f
C20 VDD1 VDD2 1.30724f
C21 VDD2 VSUBS 1.183351f
C22 VDD1 VSUBS 6.686389f
C23 VTAIL VSUBS 1.462144f
C24 VN VSUBS 6.15704f
C25 VP VSUBS 2.969713f
C26 B VSUBS 5.452732f
C27 w_n3424_n3790# VSUBS 0.159298p
C28 VDD1.t2 VSUBS 0.306958f
C29 VDD1.t3 VSUBS 0.306958f
C30 VDD1.n0 VSUBS 2.48425f
C31 VDD1.t0 VSUBS 0.306958f
C32 VDD1.t1 VSUBS 0.306958f
C33 VDD1.n1 VSUBS 3.36077f
C34 VP.t2 VSUBS 4.1562f
C35 VP.n0 VSUBS 1.55063f
C36 VP.n1 VSUBS 0.02863f
C37 VP.n2 VSUBS 0.056902f
C38 VP.n3 VSUBS 0.02863f
C39 VP.n4 VSUBS 0.053359f
C40 VP.t1 VSUBS 4.6122f
C41 VP.t0 VSUBS 4.59485f
C42 VP.n5 VSUBS 4.72038f
C43 VP.n6 VSUBS 1.81166f
C44 VP.t3 VSUBS 4.1562f
C45 VP.n7 VSUBS 1.55063f
C46 VP.n8 VSUBS 0.029385f
C47 VP.n9 VSUBS 0.046209f
C48 VP.n10 VSUBS 0.02863f
C49 VP.n11 VSUBS 0.02863f
C50 VP.n12 VSUBS 0.053359f
C51 VP.n13 VSUBS 0.056902f
C52 VP.n14 VSUBS 0.023145f
C53 VP.n15 VSUBS 0.02863f
C54 VP.n16 VSUBS 0.02863f
C55 VP.n17 VSUBS 0.02863f
C56 VP.n18 VSUBS 0.053359f
C57 VP.n19 VSUBS 0.053359f
C58 VP.n20 VSUBS 0.029385f
C59 VP.n21 VSUBS 0.046209f
C60 VP.n22 VSUBS 0.087876f
C61 VTAIL.n0 VSUBS 0.025525f
C62 VTAIL.n1 VSUBS 0.02378f
C63 VTAIL.n2 VSUBS 0.013154f
C64 VTAIL.n3 VSUBS 0.030203f
C65 VTAIL.n4 VSUBS 0.01353f
C66 VTAIL.n5 VSUBS 0.02378f
C67 VTAIL.n6 VSUBS 0.012778f
C68 VTAIL.n7 VSUBS 0.030203f
C69 VTAIL.n8 VSUBS 0.01353f
C70 VTAIL.n9 VSUBS 0.02378f
C71 VTAIL.n10 VSUBS 0.012778f
C72 VTAIL.n11 VSUBS 0.030203f
C73 VTAIL.n12 VSUBS 0.01353f
C74 VTAIL.n13 VSUBS 0.02378f
C75 VTAIL.n14 VSUBS 0.012778f
C76 VTAIL.n15 VSUBS 0.030203f
C77 VTAIL.n16 VSUBS 0.01353f
C78 VTAIL.n17 VSUBS 0.02378f
C79 VTAIL.n18 VSUBS 0.012778f
C80 VTAIL.n19 VSUBS 0.030203f
C81 VTAIL.n20 VSUBS 0.01353f
C82 VTAIL.n21 VSUBS 0.02378f
C83 VTAIL.n22 VSUBS 0.012778f
C84 VTAIL.n23 VSUBS 0.022652f
C85 VTAIL.n24 VSUBS 0.019214f
C86 VTAIL.t7 VSUBS 0.064606f
C87 VTAIL.n25 VSUBS 0.161384f
C88 VTAIL.n26 VSUBS 1.4223f
C89 VTAIL.n27 VSUBS 0.012778f
C90 VTAIL.n28 VSUBS 0.01353f
C91 VTAIL.n29 VSUBS 0.030203f
C92 VTAIL.n30 VSUBS 0.030203f
C93 VTAIL.n31 VSUBS 0.01353f
C94 VTAIL.n32 VSUBS 0.012778f
C95 VTAIL.n33 VSUBS 0.02378f
C96 VTAIL.n34 VSUBS 0.02378f
C97 VTAIL.n35 VSUBS 0.012778f
C98 VTAIL.n36 VSUBS 0.01353f
C99 VTAIL.n37 VSUBS 0.030203f
C100 VTAIL.n38 VSUBS 0.030203f
C101 VTAIL.n39 VSUBS 0.01353f
C102 VTAIL.n40 VSUBS 0.012778f
C103 VTAIL.n41 VSUBS 0.02378f
C104 VTAIL.n42 VSUBS 0.02378f
C105 VTAIL.n43 VSUBS 0.012778f
C106 VTAIL.n44 VSUBS 0.01353f
C107 VTAIL.n45 VSUBS 0.030203f
C108 VTAIL.n46 VSUBS 0.030203f
C109 VTAIL.n47 VSUBS 0.01353f
C110 VTAIL.n48 VSUBS 0.012778f
C111 VTAIL.n49 VSUBS 0.02378f
C112 VTAIL.n50 VSUBS 0.02378f
C113 VTAIL.n51 VSUBS 0.012778f
C114 VTAIL.n52 VSUBS 0.01353f
C115 VTAIL.n53 VSUBS 0.030203f
C116 VTAIL.n54 VSUBS 0.030203f
C117 VTAIL.n55 VSUBS 0.01353f
C118 VTAIL.n56 VSUBS 0.012778f
C119 VTAIL.n57 VSUBS 0.02378f
C120 VTAIL.n58 VSUBS 0.02378f
C121 VTAIL.n59 VSUBS 0.012778f
C122 VTAIL.n60 VSUBS 0.01353f
C123 VTAIL.n61 VSUBS 0.030203f
C124 VTAIL.n62 VSUBS 0.030203f
C125 VTAIL.n63 VSUBS 0.01353f
C126 VTAIL.n64 VSUBS 0.012778f
C127 VTAIL.n65 VSUBS 0.02378f
C128 VTAIL.n66 VSUBS 0.02378f
C129 VTAIL.n67 VSUBS 0.012778f
C130 VTAIL.n68 VSUBS 0.012778f
C131 VTAIL.n69 VSUBS 0.01353f
C132 VTAIL.n70 VSUBS 0.030203f
C133 VTAIL.n71 VSUBS 0.030203f
C134 VTAIL.n72 VSUBS 0.071063f
C135 VTAIL.n73 VSUBS 0.013154f
C136 VTAIL.n74 VSUBS 0.012778f
C137 VTAIL.n75 VSUBS 0.061138f
C138 VTAIL.n76 VSUBS 0.035826f
C139 VTAIL.n77 VSUBS 0.199342f
C140 VTAIL.n78 VSUBS 0.025525f
C141 VTAIL.n79 VSUBS 0.02378f
C142 VTAIL.n80 VSUBS 0.013154f
C143 VTAIL.n81 VSUBS 0.030203f
C144 VTAIL.n82 VSUBS 0.01353f
C145 VTAIL.n83 VSUBS 0.02378f
C146 VTAIL.n84 VSUBS 0.012778f
C147 VTAIL.n85 VSUBS 0.030203f
C148 VTAIL.n86 VSUBS 0.01353f
C149 VTAIL.n87 VSUBS 0.02378f
C150 VTAIL.n88 VSUBS 0.012778f
C151 VTAIL.n89 VSUBS 0.030203f
C152 VTAIL.n90 VSUBS 0.01353f
C153 VTAIL.n91 VSUBS 0.02378f
C154 VTAIL.n92 VSUBS 0.012778f
C155 VTAIL.n93 VSUBS 0.030203f
C156 VTAIL.n94 VSUBS 0.01353f
C157 VTAIL.n95 VSUBS 0.02378f
C158 VTAIL.n96 VSUBS 0.012778f
C159 VTAIL.n97 VSUBS 0.030203f
C160 VTAIL.n98 VSUBS 0.01353f
C161 VTAIL.n99 VSUBS 0.02378f
C162 VTAIL.n100 VSUBS 0.012778f
C163 VTAIL.n101 VSUBS 0.022652f
C164 VTAIL.n102 VSUBS 0.019214f
C165 VTAIL.t1 VSUBS 0.064606f
C166 VTAIL.n103 VSUBS 0.161384f
C167 VTAIL.n104 VSUBS 1.4223f
C168 VTAIL.n105 VSUBS 0.012778f
C169 VTAIL.n106 VSUBS 0.01353f
C170 VTAIL.n107 VSUBS 0.030203f
C171 VTAIL.n108 VSUBS 0.030203f
C172 VTAIL.n109 VSUBS 0.01353f
C173 VTAIL.n110 VSUBS 0.012778f
C174 VTAIL.n111 VSUBS 0.02378f
C175 VTAIL.n112 VSUBS 0.02378f
C176 VTAIL.n113 VSUBS 0.012778f
C177 VTAIL.n114 VSUBS 0.01353f
C178 VTAIL.n115 VSUBS 0.030203f
C179 VTAIL.n116 VSUBS 0.030203f
C180 VTAIL.n117 VSUBS 0.01353f
C181 VTAIL.n118 VSUBS 0.012778f
C182 VTAIL.n119 VSUBS 0.02378f
C183 VTAIL.n120 VSUBS 0.02378f
C184 VTAIL.n121 VSUBS 0.012778f
C185 VTAIL.n122 VSUBS 0.01353f
C186 VTAIL.n123 VSUBS 0.030203f
C187 VTAIL.n124 VSUBS 0.030203f
C188 VTAIL.n125 VSUBS 0.01353f
C189 VTAIL.n126 VSUBS 0.012778f
C190 VTAIL.n127 VSUBS 0.02378f
C191 VTAIL.n128 VSUBS 0.02378f
C192 VTAIL.n129 VSUBS 0.012778f
C193 VTAIL.n130 VSUBS 0.01353f
C194 VTAIL.n131 VSUBS 0.030203f
C195 VTAIL.n132 VSUBS 0.030203f
C196 VTAIL.n133 VSUBS 0.01353f
C197 VTAIL.n134 VSUBS 0.012778f
C198 VTAIL.n135 VSUBS 0.02378f
C199 VTAIL.n136 VSUBS 0.02378f
C200 VTAIL.n137 VSUBS 0.012778f
C201 VTAIL.n138 VSUBS 0.01353f
C202 VTAIL.n139 VSUBS 0.030203f
C203 VTAIL.n140 VSUBS 0.030203f
C204 VTAIL.n141 VSUBS 0.01353f
C205 VTAIL.n142 VSUBS 0.012778f
C206 VTAIL.n143 VSUBS 0.02378f
C207 VTAIL.n144 VSUBS 0.02378f
C208 VTAIL.n145 VSUBS 0.012778f
C209 VTAIL.n146 VSUBS 0.012778f
C210 VTAIL.n147 VSUBS 0.01353f
C211 VTAIL.n148 VSUBS 0.030203f
C212 VTAIL.n149 VSUBS 0.030203f
C213 VTAIL.n150 VSUBS 0.071063f
C214 VTAIL.n151 VSUBS 0.013154f
C215 VTAIL.n152 VSUBS 0.012778f
C216 VTAIL.n153 VSUBS 0.061138f
C217 VTAIL.n154 VSUBS 0.035826f
C218 VTAIL.n155 VSUBS 0.329966f
C219 VTAIL.n156 VSUBS 0.025525f
C220 VTAIL.n157 VSUBS 0.02378f
C221 VTAIL.n158 VSUBS 0.013154f
C222 VTAIL.n159 VSUBS 0.030203f
C223 VTAIL.n160 VSUBS 0.01353f
C224 VTAIL.n161 VSUBS 0.02378f
C225 VTAIL.n162 VSUBS 0.012778f
C226 VTAIL.n163 VSUBS 0.030203f
C227 VTAIL.n164 VSUBS 0.01353f
C228 VTAIL.n165 VSUBS 0.02378f
C229 VTAIL.n166 VSUBS 0.012778f
C230 VTAIL.n167 VSUBS 0.030203f
C231 VTAIL.n168 VSUBS 0.01353f
C232 VTAIL.n169 VSUBS 0.02378f
C233 VTAIL.n170 VSUBS 0.012778f
C234 VTAIL.n171 VSUBS 0.030203f
C235 VTAIL.n172 VSUBS 0.01353f
C236 VTAIL.n173 VSUBS 0.02378f
C237 VTAIL.n174 VSUBS 0.012778f
C238 VTAIL.n175 VSUBS 0.030203f
C239 VTAIL.n176 VSUBS 0.01353f
C240 VTAIL.n177 VSUBS 0.02378f
C241 VTAIL.n178 VSUBS 0.012778f
C242 VTAIL.n179 VSUBS 0.022652f
C243 VTAIL.n180 VSUBS 0.019214f
C244 VTAIL.t2 VSUBS 0.064606f
C245 VTAIL.n181 VSUBS 0.161384f
C246 VTAIL.n182 VSUBS 1.4223f
C247 VTAIL.n183 VSUBS 0.012778f
C248 VTAIL.n184 VSUBS 0.01353f
C249 VTAIL.n185 VSUBS 0.030203f
C250 VTAIL.n186 VSUBS 0.030203f
C251 VTAIL.n187 VSUBS 0.01353f
C252 VTAIL.n188 VSUBS 0.012778f
C253 VTAIL.n189 VSUBS 0.02378f
C254 VTAIL.n190 VSUBS 0.02378f
C255 VTAIL.n191 VSUBS 0.012778f
C256 VTAIL.n192 VSUBS 0.01353f
C257 VTAIL.n193 VSUBS 0.030203f
C258 VTAIL.n194 VSUBS 0.030203f
C259 VTAIL.n195 VSUBS 0.01353f
C260 VTAIL.n196 VSUBS 0.012778f
C261 VTAIL.n197 VSUBS 0.02378f
C262 VTAIL.n198 VSUBS 0.02378f
C263 VTAIL.n199 VSUBS 0.012778f
C264 VTAIL.n200 VSUBS 0.01353f
C265 VTAIL.n201 VSUBS 0.030203f
C266 VTAIL.n202 VSUBS 0.030203f
C267 VTAIL.n203 VSUBS 0.01353f
C268 VTAIL.n204 VSUBS 0.012778f
C269 VTAIL.n205 VSUBS 0.02378f
C270 VTAIL.n206 VSUBS 0.02378f
C271 VTAIL.n207 VSUBS 0.012778f
C272 VTAIL.n208 VSUBS 0.01353f
C273 VTAIL.n209 VSUBS 0.030203f
C274 VTAIL.n210 VSUBS 0.030203f
C275 VTAIL.n211 VSUBS 0.01353f
C276 VTAIL.n212 VSUBS 0.012778f
C277 VTAIL.n213 VSUBS 0.02378f
C278 VTAIL.n214 VSUBS 0.02378f
C279 VTAIL.n215 VSUBS 0.012778f
C280 VTAIL.n216 VSUBS 0.01353f
C281 VTAIL.n217 VSUBS 0.030203f
C282 VTAIL.n218 VSUBS 0.030203f
C283 VTAIL.n219 VSUBS 0.01353f
C284 VTAIL.n220 VSUBS 0.012778f
C285 VTAIL.n221 VSUBS 0.02378f
C286 VTAIL.n222 VSUBS 0.02378f
C287 VTAIL.n223 VSUBS 0.012778f
C288 VTAIL.n224 VSUBS 0.012778f
C289 VTAIL.n225 VSUBS 0.01353f
C290 VTAIL.n226 VSUBS 0.030203f
C291 VTAIL.n227 VSUBS 0.030203f
C292 VTAIL.n228 VSUBS 0.071063f
C293 VTAIL.n229 VSUBS 0.013154f
C294 VTAIL.n230 VSUBS 0.012778f
C295 VTAIL.n231 VSUBS 0.061138f
C296 VTAIL.n232 VSUBS 0.035826f
C297 VTAIL.n233 VSUBS 1.81918f
C298 VTAIL.n234 VSUBS 0.025525f
C299 VTAIL.n235 VSUBS 0.02378f
C300 VTAIL.n236 VSUBS 0.013154f
C301 VTAIL.n237 VSUBS 0.030203f
C302 VTAIL.n238 VSUBS 0.012778f
C303 VTAIL.n239 VSUBS 0.01353f
C304 VTAIL.n240 VSUBS 0.02378f
C305 VTAIL.n241 VSUBS 0.012778f
C306 VTAIL.n242 VSUBS 0.030203f
C307 VTAIL.n243 VSUBS 0.01353f
C308 VTAIL.n244 VSUBS 0.02378f
C309 VTAIL.n245 VSUBS 0.012778f
C310 VTAIL.n246 VSUBS 0.030203f
C311 VTAIL.n247 VSUBS 0.01353f
C312 VTAIL.n248 VSUBS 0.02378f
C313 VTAIL.n249 VSUBS 0.012778f
C314 VTAIL.n250 VSUBS 0.030203f
C315 VTAIL.n251 VSUBS 0.01353f
C316 VTAIL.n252 VSUBS 0.02378f
C317 VTAIL.n253 VSUBS 0.012778f
C318 VTAIL.n254 VSUBS 0.030203f
C319 VTAIL.n255 VSUBS 0.01353f
C320 VTAIL.n256 VSUBS 0.02378f
C321 VTAIL.n257 VSUBS 0.012778f
C322 VTAIL.n258 VSUBS 0.022652f
C323 VTAIL.n259 VSUBS 0.019214f
C324 VTAIL.t6 VSUBS 0.064606f
C325 VTAIL.n260 VSUBS 0.161384f
C326 VTAIL.n261 VSUBS 1.4223f
C327 VTAIL.n262 VSUBS 0.012778f
C328 VTAIL.n263 VSUBS 0.01353f
C329 VTAIL.n264 VSUBS 0.030203f
C330 VTAIL.n265 VSUBS 0.030203f
C331 VTAIL.n266 VSUBS 0.01353f
C332 VTAIL.n267 VSUBS 0.012778f
C333 VTAIL.n268 VSUBS 0.02378f
C334 VTAIL.n269 VSUBS 0.02378f
C335 VTAIL.n270 VSUBS 0.012778f
C336 VTAIL.n271 VSUBS 0.01353f
C337 VTAIL.n272 VSUBS 0.030203f
C338 VTAIL.n273 VSUBS 0.030203f
C339 VTAIL.n274 VSUBS 0.01353f
C340 VTAIL.n275 VSUBS 0.012778f
C341 VTAIL.n276 VSUBS 0.02378f
C342 VTAIL.n277 VSUBS 0.02378f
C343 VTAIL.n278 VSUBS 0.012778f
C344 VTAIL.n279 VSUBS 0.01353f
C345 VTAIL.n280 VSUBS 0.030203f
C346 VTAIL.n281 VSUBS 0.030203f
C347 VTAIL.n282 VSUBS 0.01353f
C348 VTAIL.n283 VSUBS 0.012778f
C349 VTAIL.n284 VSUBS 0.02378f
C350 VTAIL.n285 VSUBS 0.02378f
C351 VTAIL.n286 VSUBS 0.012778f
C352 VTAIL.n287 VSUBS 0.01353f
C353 VTAIL.n288 VSUBS 0.030203f
C354 VTAIL.n289 VSUBS 0.030203f
C355 VTAIL.n290 VSUBS 0.01353f
C356 VTAIL.n291 VSUBS 0.012778f
C357 VTAIL.n292 VSUBS 0.02378f
C358 VTAIL.n293 VSUBS 0.02378f
C359 VTAIL.n294 VSUBS 0.012778f
C360 VTAIL.n295 VSUBS 0.01353f
C361 VTAIL.n296 VSUBS 0.030203f
C362 VTAIL.n297 VSUBS 0.030203f
C363 VTAIL.n298 VSUBS 0.01353f
C364 VTAIL.n299 VSUBS 0.012778f
C365 VTAIL.n300 VSUBS 0.02378f
C366 VTAIL.n301 VSUBS 0.02378f
C367 VTAIL.n302 VSUBS 0.012778f
C368 VTAIL.n303 VSUBS 0.01353f
C369 VTAIL.n304 VSUBS 0.030203f
C370 VTAIL.n305 VSUBS 0.030203f
C371 VTAIL.n306 VSUBS 0.071063f
C372 VTAIL.n307 VSUBS 0.013154f
C373 VTAIL.n308 VSUBS 0.012778f
C374 VTAIL.n309 VSUBS 0.061138f
C375 VTAIL.n310 VSUBS 0.035826f
C376 VTAIL.n311 VSUBS 1.81918f
C377 VTAIL.n312 VSUBS 0.025525f
C378 VTAIL.n313 VSUBS 0.02378f
C379 VTAIL.n314 VSUBS 0.013154f
C380 VTAIL.n315 VSUBS 0.030203f
C381 VTAIL.n316 VSUBS 0.012778f
C382 VTAIL.n317 VSUBS 0.01353f
C383 VTAIL.n318 VSUBS 0.02378f
C384 VTAIL.n319 VSUBS 0.012778f
C385 VTAIL.n320 VSUBS 0.030203f
C386 VTAIL.n321 VSUBS 0.01353f
C387 VTAIL.n322 VSUBS 0.02378f
C388 VTAIL.n323 VSUBS 0.012778f
C389 VTAIL.n324 VSUBS 0.030203f
C390 VTAIL.n325 VSUBS 0.01353f
C391 VTAIL.n326 VSUBS 0.02378f
C392 VTAIL.n327 VSUBS 0.012778f
C393 VTAIL.n328 VSUBS 0.030203f
C394 VTAIL.n329 VSUBS 0.01353f
C395 VTAIL.n330 VSUBS 0.02378f
C396 VTAIL.n331 VSUBS 0.012778f
C397 VTAIL.n332 VSUBS 0.030203f
C398 VTAIL.n333 VSUBS 0.01353f
C399 VTAIL.n334 VSUBS 0.02378f
C400 VTAIL.n335 VSUBS 0.012778f
C401 VTAIL.n336 VSUBS 0.022652f
C402 VTAIL.n337 VSUBS 0.019214f
C403 VTAIL.t5 VSUBS 0.064606f
C404 VTAIL.n338 VSUBS 0.161384f
C405 VTAIL.n339 VSUBS 1.4223f
C406 VTAIL.n340 VSUBS 0.012778f
C407 VTAIL.n341 VSUBS 0.01353f
C408 VTAIL.n342 VSUBS 0.030203f
C409 VTAIL.n343 VSUBS 0.030203f
C410 VTAIL.n344 VSUBS 0.01353f
C411 VTAIL.n345 VSUBS 0.012778f
C412 VTAIL.n346 VSUBS 0.02378f
C413 VTAIL.n347 VSUBS 0.02378f
C414 VTAIL.n348 VSUBS 0.012778f
C415 VTAIL.n349 VSUBS 0.01353f
C416 VTAIL.n350 VSUBS 0.030203f
C417 VTAIL.n351 VSUBS 0.030203f
C418 VTAIL.n352 VSUBS 0.01353f
C419 VTAIL.n353 VSUBS 0.012778f
C420 VTAIL.n354 VSUBS 0.02378f
C421 VTAIL.n355 VSUBS 0.02378f
C422 VTAIL.n356 VSUBS 0.012778f
C423 VTAIL.n357 VSUBS 0.01353f
C424 VTAIL.n358 VSUBS 0.030203f
C425 VTAIL.n359 VSUBS 0.030203f
C426 VTAIL.n360 VSUBS 0.01353f
C427 VTAIL.n361 VSUBS 0.012778f
C428 VTAIL.n362 VSUBS 0.02378f
C429 VTAIL.n363 VSUBS 0.02378f
C430 VTAIL.n364 VSUBS 0.012778f
C431 VTAIL.n365 VSUBS 0.01353f
C432 VTAIL.n366 VSUBS 0.030203f
C433 VTAIL.n367 VSUBS 0.030203f
C434 VTAIL.n368 VSUBS 0.01353f
C435 VTAIL.n369 VSUBS 0.012778f
C436 VTAIL.n370 VSUBS 0.02378f
C437 VTAIL.n371 VSUBS 0.02378f
C438 VTAIL.n372 VSUBS 0.012778f
C439 VTAIL.n373 VSUBS 0.01353f
C440 VTAIL.n374 VSUBS 0.030203f
C441 VTAIL.n375 VSUBS 0.030203f
C442 VTAIL.n376 VSUBS 0.01353f
C443 VTAIL.n377 VSUBS 0.012778f
C444 VTAIL.n378 VSUBS 0.02378f
C445 VTAIL.n379 VSUBS 0.02378f
C446 VTAIL.n380 VSUBS 0.012778f
C447 VTAIL.n381 VSUBS 0.01353f
C448 VTAIL.n382 VSUBS 0.030203f
C449 VTAIL.n383 VSUBS 0.030203f
C450 VTAIL.n384 VSUBS 0.071063f
C451 VTAIL.n385 VSUBS 0.013154f
C452 VTAIL.n386 VSUBS 0.012778f
C453 VTAIL.n387 VSUBS 0.061138f
C454 VTAIL.n388 VSUBS 0.035826f
C455 VTAIL.n389 VSUBS 0.329966f
C456 VTAIL.n390 VSUBS 0.025525f
C457 VTAIL.n391 VSUBS 0.02378f
C458 VTAIL.n392 VSUBS 0.013154f
C459 VTAIL.n393 VSUBS 0.030203f
C460 VTAIL.n394 VSUBS 0.012778f
C461 VTAIL.n395 VSUBS 0.01353f
C462 VTAIL.n396 VSUBS 0.02378f
C463 VTAIL.n397 VSUBS 0.012778f
C464 VTAIL.n398 VSUBS 0.030203f
C465 VTAIL.n399 VSUBS 0.01353f
C466 VTAIL.n400 VSUBS 0.02378f
C467 VTAIL.n401 VSUBS 0.012778f
C468 VTAIL.n402 VSUBS 0.030203f
C469 VTAIL.n403 VSUBS 0.01353f
C470 VTAIL.n404 VSUBS 0.02378f
C471 VTAIL.n405 VSUBS 0.012778f
C472 VTAIL.n406 VSUBS 0.030203f
C473 VTAIL.n407 VSUBS 0.01353f
C474 VTAIL.n408 VSUBS 0.02378f
C475 VTAIL.n409 VSUBS 0.012778f
C476 VTAIL.n410 VSUBS 0.030203f
C477 VTAIL.n411 VSUBS 0.01353f
C478 VTAIL.n412 VSUBS 0.02378f
C479 VTAIL.n413 VSUBS 0.012778f
C480 VTAIL.n414 VSUBS 0.022652f
C481 VTAIL.n415 VSUBS 0.019214f
C482 VTAIL.t0 VSUBS 0.064606f
C483 VTAIL.n416 VSUBS 0.161384f
C484 VTAIL.n417 VSUBS 1.4223f
C485 VTAIL.n418 VSUBS 0.012778f
C486 VTAIL.n419 VSUBS 0.01353f
C487 VTAIL.n420 VSUBS 0.030203f
C488 VTAIL.n421 VSUBS 0.030203f
C489 VTAIL.n422 VSUBS 0.01353f
C490 VTAIL.n423 VSUBS 0.012778f
C491 VTAIL.n424 VSUBS 0.02378f
C492 VTAIL.n425 VSUBS 0.02378f
C493 VTAIL.n426 VSUBS 0.012778f
C494 VTAIL.n427 VSUBS 0.01353f
C495 VTAIL.n428 VSUBS 0.030203f
C496 VTAIL.n429 VSUBS 0.030203f
C497 VTAIL.n430 VSUBS 0.01353f
C498 VTAIL.n431 VSUBS 0.012778f
C499 VTAIL.n432 VSUBS 0.02378f
C500 VTAIL.n433 VSUBS 0.02378f
C501 VTAIL.n434 VSUBS 0.012778f
C502 VTAIL.n435 VSUBS 0.01353f
C503 VTAIL.n436 VSUBS 0.030203f
C504 VTAIL.n437 VSUBS 0.030203f
C505 VTAIL.n438 VSUBS 0.01353f
C506 VTAIL.n439 VSUBS 0.012778f
C507 VTAIL.n440 VSUBS 0.02378f
C508 VTAIL.n441 VSUBS 0.02378f
C509 VTAIL.n442 VSUBS 0.012778f
C510 VTAIL.n443 VSUBS 0.01353f
C511 VTAIL.n444 VSUBS 0.030203f
C512 VTAIL.n445 VSUBS 0.030203f
C513 VTAIL.n446 VSUBS 0.01353f
C514 VTAIL.n447 VSUBS 0.012778f
C515 VTAIL.n448 VSUBS 0.02378f
C516 VTAIL.n449 VSUBS 0.02378f
C517 VTAIL.n450 VSUBS 0.012778f
C518 VTAIL.n451 VSUBS 0.01353f
C519 VTAIL.n452 VSUBS 0.030203f
C520 VTAIL.n453 VSUBS 0.030203f
C521 VTAIL.n454 VSUBS 0.01353f
C522 VTAIL.n455 VSUBS 0.012778f
C523 VTAIL.n456 VSUBS 0.02378f
C524 VTAIL.n457 VSUBS 0.02378f
C525 VTAIL.n458 VSUBS 0.012778f
C526 VTAIL.n459 VSUBS 0.01353f
C527 VTAIL.n460 VSUBS 0.030203f
C528 VTAIL.n461 VSUBS 0.030203f
C529 VTAIL.n462 VSUBS 0.071063f
C530 VTAIL.n463 VSUBS 0.013154f
C531 VTAIL.n464 VSUBS 0.012778f
C532 VTAIL.n465 VSUBS 0.061138f
C533 VTAIL.n466 VSUBS 0.035826f
C534 VTAIL.n467 VSUBS 0.329966f
C535 VTAIL.n468 VSUBS 0.025525f
C536 VTAIL.n469 VSUBS 0.02378f
C537 VTAIL.n470 VSUBS 0.013154f
C538 VTAIL.n471 VSUBS 0.030203f
C539 VTAIL.n472 VSUBS 0.012778f
C540 VTAIL.n473 VSUBS 0.01353f
C541 VTAIL.n474 VSUBS 0.02378f
C542 VTAIL.n475 VSUBS 0.012778f
C543 VTAIL.n476 VSUBS 0.030203f
C544 VTAIL.n477 VSUBS 0.01353f
C545 VTAIL.n478 VSUBS 0.02378f
C546 VTAIL.n479 VSUBS 0.012778f
C547 VTAIL.n480 VSUBS 0.030203f
C548 VTAIL.n481 VSUBS 0.01353f
C549 VTAIL.n482 VSUBS 0.02378f
C550 VTAIL.n483 VSUBS 0.012778f
C551 VTAIL.n484 VSUBS 0.030203f
C552 VTAIL.n485 VSUBS 0.01353f
C553 VTAIL.n486 VSUBS 0.02378f
C554 VTAIL.n487 VSUBS 0.012778f
C555 VTAIL.n488 VSUBS 0.030203f
C556 VTAIL.n489 VSUBS 0.01353f
C557 VTAIL.n490 VSUBS 0.02378f
C558 VTAIL.n491 VSUBS 0.012778f
C559 VTAIL.n492 VSUBS 0.022652f
C560 VTAIL.n493 VSUBS 0.019214f
C561 VTAIL.t3 VSUBS 0.064606f
C562 VTAIL.n494 VSUBS 0.161384f
C563 VTAIL.n495 VSUBS 1.4223f
C564 VTAIL.n496 VSUBS 0.012778f
C565 VTAIL.n497 VSUBS 0.01353f
C566 VTAIL.n498 VSUBS 0.030203f
C567 VTAIL.n499 VSUBS 0.030203f
C568 VTAIL.n500 VSUBS 0.01353f
C569 VTAIL.n501 VSUBS 0.012778f
C570 VTAIL.n502 VSUBS 0.02378f
C571 VTAIL.n503 VSUBS 0.02378f
C572 VTAIL.n504 VSUBS 0.012778f
C573 VTAIL.n505 VSUBS 0.01353f
C574 VTAIL.n506 VSUBS 0.030203f
C575 VTAIL.n507 VSUBS 0.030203f
C576 VTAIL.n508 VSUBS 0.01353f
C577 VTAIL.n509 VSUBS 0.012778f
C578 VTAIL.n510 VSUBS 0.02378f
C579 VTAIL.n511 VSUBS 0.02378f
C580 VTAIL.n512 VSUBS 0.012778f
C581 VTAIL.n513 VSUBS 0.01353f
C582 VTAIL.n514 VSUBS 0.030203f
C583 VTAIL.n515 VSUBS 0.030203f
C584 VTAIL.n516 VSUBS 0.01353f
C585 VTAIL.n517 VSUBS 0.012778f
C586 VTAIL.n518 VSUBS 0.02378f
C587 VTAIL.n519 VSUBS 0.02378f
C588 VTAIL.n520 VSUBS 0.012778f
C589 VTAIL.n521 VSUBS 0.01353f
C590 VTAIL.n522 VSUBS 0.030203f
C591 VTAIL.n523 VSUBS 0.030203f
C592 VTAIL.n524 VSUBS 0.01353f
C593 VTAIL.n525 VSUBS 0.012778f
C594 VTAIL.n526 VSUBS 0.02378f
C595 VTAIL.n527 VSUBS 0.02378f
C596 VTAIL.n528 VSUBS 0.012778f
C597 VTAIL.n529 VSUBS 0.01353f
C598 VTAIL.n530 VSUBS 0.030203f
C599 VTAIL.n531 VSUBS 0.030203f
C600 VTAIL.n532 VSUBS 0.01353f
C601 VTAIL.n533 VSUBS 0.012778f
C602 VTAIL.n534 VSUBS 0.02378f
C603 VTAIL.n535 VSUBS 0.02378f
C604 VTAIL.n536 VSUBS 0.012778f
C605 VTAIL.n537 VSUBS 0.01353f
C606 VTAIL.n538 VSUBS 0.030203f
C607 VTAIL.n539 VSUBS 0.030203f
C608 VTAIL.n540 VSUBS 0.071063f
C609 VTAIL.n541 VSUBS 0.013154f
C610 VTAIL.n542 VSUBS 0.012778f
C611 VTAIL.n543 VSUBS 0.061138f
C612 VTAIL.n544 VSUBS 0.035826f
C613 VTAIL.n545 VSUBS 1.81918f
C614 VTAIL.n546 VSUBS 0.025525f
C615 VTAIL.n547 VSUBS 0.02378f
C616 VTAIL.n548 VSUBS 0.013154f
C617 VTAIL.n549 VSUBS 0.030203f
C618 VTAIL.n550 VSUBS 0.01353f
C619 VTAIL.n551 VSUBS 0.02378f
C620 VTAIL.n552 VSUBS 0.012778f
C621 VTAIL.n553 VSUBS 0.030203f
C622 VTAIL.n554 VSUBS 0.01353f
C623 VTAIL.n555 VSUBS 0.02378f
C624 VTAIL.n556 VSUBS 0.012778f
C625 VTAIL.n557 VSUBS 0.030203f
C626 VTAIL.n558 VSUBS 0.01353f
C627 VTAIL.n559 VSUBS 0.02378f
C628 VTAIL.n560 VSUBS 0.012778f
C629 VTAIL.n561 VSUBS 0.030203f
C630 VTAIL.n562 VSUBS 0.01353f
C631 VTAIL.n563 VSUBS 0.02378f
C632 VTAIL.n564 VSUBS 0.012778f
C633 VTAIL.n565 VSUBS 0.030203f
C634 VTAIL.n566 VSUBS 0.01353f
C635 VTAIL.n567 VSUBS 0.02378f
C636 VTAIL.n568 VSUBS 0.012778f
C637 VTAIL.n569 VSUBS 0.022652f
C638 VTAIL.n570 VSUBS 0.019214f
C639 VTAIL.t4 VSUBS 0.064606f
C640 VTAIL.n571 VSUBS 0.161384f
C641 VTAIL.n572 VSUBS 1.4223f
C642 VTAIL.n573 VSUBS 0.012778f
C643 VTAIL.n574 VSUBS 0.01353f
C644 VTAIL.n575 VSUBS 0.030203f
C645 VTAIL.n576 VSUBS 0.030203f
C646 VTAIL.n577 VSUBS 0.01353f
C647 VTAIL.n578 VSUBS 0.012778f
C648 VTAIL.n579 VSUBS 0.02378f
C649 VTAIL.n580 VSUBS 0.02378f
C650 VTAIL.n581 VSUBS 0.012778f
C651 VTAIL.n582 VSUBS 0.01353f
C652 VTAIL.n583 VSUBS 0.030203f
C653 VTAIL.n584 VSUBS 0.030203f
C654 VTAIL.n585 VSUBS 0.01353f
C655 VTAIL.n586 VSUBS 0.012778f
C656 VTAIL.n587 VSUBS 0.02378f
C657 VTAIL.n588 VSUBS 0.02378f
C658 VTAIL.n589 VSUBS 0.012778f
C659 VTAIL.n590 VSUBS 0.01353f
C660 VTAIL.n591 VSUBS 0.030203f
C661 VTAIL.n592 VSUBS 0.030203f
C662 VTAIL.n593 VSUBS 0.01353f
C663 VTAIL.n594 VSUBS 0.012778f
C664 VTAIL.n595 VSUBS 0.02378f
C665 VTAIL.n596 VSUBS 0.02378f
C666 VTAIL.n597 VSUBS 0.012778f
C667 VTAIL.n598 VSUBS 0.01353f
C668 VTAIL.n599 VSUBS 0.030203f
C669 VTAIL.n600 VSUBS 0.030203f
C670 VTAIL.n601 VSUBS 0.01353f
C671 VTAIL.n602 VSUBS 0.012778f
C672 VTAIL.n603 VSUBS 0.02378f
C673 VTAIL.n604 VSUBS 0.02378f
C674 VTAIL.n605 VSUBS 0.012778f
C675 VTAIL.n606 VSUBS 0.01353f
C676 VTAIL.n607 VSUBS 0.030203f
C677 VTAIL.n608 VSUBS 0.030203f
C678 VTAIL.n609 VSUBS 0.01353f
C679 VTAIL.n610 VSUBS 0.012778f
C680 VTAIL.n611 VSUBS 0.02378f
C681 VTAIL.n612 VSUBS 0.02378f
C682 VTAIL.n613 VSUBS 0.012778f
C683 VTAIL.n614 VSUBS 0.012778f
C684 VTAIL.n615 VSUBS 0.01353f
C685 VTAIL.n616 VSUBS 0.030203f
C686 VTAIL.n617 VSUBS 0.030203f
C687 VTAIL.n618 VSUBS 0.071063f
C688 VTAIL.n619 VSUBS 0.013154f
C689 VTAIL.n620 VSUBS 0.012778f
C690 VTAIL.n621 VSUBS 0.061138f
C691 VTAIL.n622 VSUBS 0.035826f
C692 VTAIL.n623 VSUBS 1.67964f
C693 VDD2.t3 VSUBS 0.302008f
C694 VDD2.t1 VSUBS 0.302008f
C695 VDD2.n0 VSUBS 3.2803f
C696 VDD2.t2 VSUBS 0.302008f
C697 VDD2.t0 VSUBS 0.302008f
C698 VDD2.n1 VSUBS 2.44355f
C699 VDD2.n2 VSUBS 4.85457f
C700 VN.t3 VSUBS 4.12943f
C701 VN.t0 VSUBS 4.14502f
C702 VN.n0 VSUBS 2.49906f
C703 VN.t1 VSUBS 4.12943f
C704 VN.t2 VSUBS 4.14502f
C705 VN.n1 VSUBS 4.2525f
C706 B.n0 VSUBS 0.004152f
C707 B.n1 VSUBS 0.004152f
C708 B.n2 VSUBS 0.006567f
C709 B.n3 VSUBS 0.006567f
C710 B.n4 VSUBS 0.006567f
C711 B.n5 VSUBS 0.006567f
C712 B.n6 VSUBS 0.006567f
C713 B.n7 VSUBS 0.006567f
C714 B.n8 VSUBS 0.006567f
C715 B.n9 VSUBS 0.006567f
C716 B.n10 VSUBS 0.006567f
C717 B.n11 VSUBS 0.006567f
C718 B.n12 VSUBS 0.006567f
C719 B.n13 VSUBS 0.006567f
C720 B.n14 VSUBS 0.006567f
C721 B.n15 VSUBS 0.006567f
C722 B.n16 VSUBS 0.006567f
C723 B.n17 VSUBS 0.006567f
C724 B.n18 VSUBS 0.006567f
C725 B.n19 VSUBS 0.006567f
C726 B.n20 VSUBS 0.006567f
C727 B.n21 VSUBS 0.006567f
C728 B.n22 VSUBS 0.006567f
C729 B.n23 VSUBS 0.006567f
C730 B.n24 VSUBS 0.016709f
C731 B.n25 VSUBS 0.006567f
C732 B.n26 VSUBS 0.006567f
C733 B.n27 VSUBS 0.006567f
C734 B.n28 VSUBS 0.006567f
C735 B.n29 VSUBS 0.006567f
C736 B.n30 VSUBS 0.006567f
C737 B.n31 VSUBS 0.006567f
C738 B.n32 VSUBS 0.006567f
C739 B.n33 VSUBS 0.006567f
C740 B.n34 VSUBS 0.006567f
C741 B.n35 VSUBS 0.006567f
C742 B.n36 VSUBS 0.006567f
C743 B.n37 VSUBS 0.006567f
C744 B.n38 VSUBS 0.006567f
C745 B.n39 VSUBS 0.006567f
C746 B.n40 VSUBS 0.006567f
C747 B.n41 VSUBS 0.006567f
C748 B.n42 VSUBS 0.006567f
C749 B.n43 VSUBS 0.006567f
C750 B.n44 VSUBS 0.006567f
C751 B.n45 VSUBS 0.006567f
C752 B.n46 VSUBS 0.006567f
C753 B.n47 VSUBS 0.006567f
C754 B.t8 VSUBS 0.242885f
C755 B.t7 VSUBS 0.284403f
C756 B.t6 VSUBS 2.29925f
C757 B.n48 VSUBS 0.453286f
C758 B.n49 VSUBS 0.267382f
C759 B.n50 VSUBS 0.015214f
C760 B.n51 VSUBS 0.006567f
C761 B.n52 VSUBS 0.006567f
C762 B.n53 VSUBS 0.006567f
C763 B.n54 VSUBS 0.006567f
C764 B.n55 VSUBS 0.006567f
C765 B.t5 VSUBS 0.242888f
C766 B.t4 VSUBS 0.284405f
C767 B.t3 VSUBS 2.29925f
C768 B.n56 VSUBS 0.453283f
C769 B.n57 VSUBS 0.267379f
C770 B.n58 VSUBS 0.006567f
C771 B.n59 VSUBS 0.006567f
C772 B.n60 VSUBS 0.006567f
C773 B.n61 VSUBS 0.006567f
C774 B.n62 VSUBS 0.006567f
C775 B.n63 VSUBS 0.006567f
C776 B.n64 VSUBS 0.006567f
C777 B.n65 VSUBS 0.006567f
C778 B.n66 VSUBS 0.006567f
C779 B.n67 VSUBS 0.006567f
C780 B.n68 VSUBS 0.006567f
C781 B.n69 VSUBS 0.006567f
C782 B.n70 VSUBS 0.006567f
C783 B.n71 VSUBS 0.006567f
C784 B.n72 VSUBS 0.006567f
C785 B.n73 VSUBS 0.006567f
C786 B.n74 VSUBS 0.006567f
C787 B.n75 VSUBS 0.006567f
C788 B.n76 VSUBS 0.006567f
C789 B.n77 VSUBS 0.006567f
C790 B.n78 VSUBS 0.006567f
C791 B.n79 VSUBS 0.006567f
C792 B.n80 VSUBS 0.006567f
C793 B.n81 VSUBS 0.015931f
C794 B.n82 VSUBS 0.006567f
C795 B.n83 VSUBS 0.006567f
C796 B.n84 VSUBS 0.006567f
C797 B.n85 VSUBS 0.006567f
C798 B.n86 VSUBS 0.006567f
C799 B.n87 VSUBS 0.006567f
C800 B.n88 VSUBS 0.006567f
C801 B.n89 VSUBS 0.006567f
C802 B.n90 VSUBS 0.006567f
C803 B.n91 VSUBS 0.006567f
C804 B.n92 VSUBS 0.006567f
C805 B.n93 VSUBS 0.006567f
C806 B.n94 VSUBS 0.006567f
C807 B.n95 VSUBS 0.006567f
C808 B.n96 VSUBS 0.006567f
C809 B.n97 VSUBS 0.006567f
C810 B.n98 VSUBS 0.006567f
C811 B.n99 VSUBS 0.006567f
C812 B.n100 VSUBS 0.006567f
C813 B.n101 VSUBS 0.006567f
C814 B.n102 VSUBS 0.006567f
C815 B.n103 VSUBS 0.006567f
C816 B.n104 VSUBS 0.006567f
C817 B.n105 VSUBS 0.006567f
C818 B.n106 VSUBS 0.006567f
C819 B.n107 VSUBS 0.006567f
C820 B.n108 VSUBS 0.006567f
C821 B.n109 VSUBS 0.006567f
C822 B.n110 VSUBS 0.006567f
C823 B.n111 VSUBS 0.006567f
C824 B.n112 VSUBS 0.006567f
C825 B.n113 VSUBS 0.006567f
C826 B.n114 VSUBS 0.006567f
C827 B.n115 VSUBS 0.006567f
C828 B.n116 VSUBS 0.006567f
C829 B.n117 VSUBS 0.006567f
C830 B.n118 VSUBS 0.006567f
C831 B.n119 VSUBS 0.006567f
C832 B.n120 VSUBS 0.006567f
C833 B.n121 VSUBS 0.006567f
C834 B.n122 VSUBS 0.006567f
C835 B.n123 VSUBS 0.006567f
C836 B.n124 VSUBS 0.006567f
C837 B.n125 VSUBS 0.015931f
C838 B.n126 VSUBS 0.006567f
C839 B.n127 VSUBS 0.006567f
C840 B.n128 VSUBS 0.006567f
C841 B.n129 VSUBS 0.006567f
C842 B.n130 VSUBS 0.006567f
C843 B.n131 VSUBS 0.006567f
C844 B.n132 VSUBS 0.006567f
C845 B.n133 VSUBS 0.006567f
C846 B.n134 VSUBS 0.006567f
C847 B.n135 VSUBS 0.006567f
C848 B.n136 VSUBS 0.006567f
C849 B.n137 VSUBS 0.006567f
C850 B.n138 VSUBS 0.006567f
C851 B.n139 VSUBS 0.006567f
C852 B.n140 VSUBS 0.006567f
C853 B.n141 VSUBS 0.006567f
C854 B.n142 VSUBS 0.006567f
C855 B.n143 VSUBS 0.006567f
C856 B.n144 VSUBS 0.006567f
C857 B.n145 VSUBS 0.006567f
C858 B.n146 VSUBS 0.006567f
C859 B.n147 VSUBS 0.006567f
C860 B.n148 VSUBS 0.006567f
C861 B.n149 VSUBS 0.006567f
C862 B.t10 VSUBS 0.242888f
C863 B.t11 VSUBS 0.284405f
C864 B.t9 VSUBS 2.29925f
C865 B.n150 VSUBS 0.453283f
C866 B.n151 VSUBS 0.267379f
C867 B.n152 VSUBS 0.006567f
C868 B.n153 VSUBS 0.006567f
C869 B.n154 VSUBS 0.006567f
C870 B.n155 VSUBS 0.006567f
C871 B.t1 VSUBS 0.242885f
C872 B.t2 VSUBS 0.284403f
C873 B.t0 VSUBS 2.29925f
C874 B.n156 VSUBS 0.453286f
C875 B.n157 VSUBS 0.267382f
C876 B.n158 VSUBS 0.015214f
C877 B.n159 VSUBS 0.006567f
C878 B.n160 VSUBS 0.006567f
C879 B.n161 VSUBS 0.006567f
C880 B.n162 VSUBS 0.006567f
C881 B.n163 VSUBS 0.006567f
C882 B.n164 VSUBS 0.006567f
C883 B.n165 VSUBS 0.006567f
C884 B.n166 VSUBS 0.006567f
C885 B.n167 VSUBS 0.006567f
C886 B.n168 VSUBS 0.006567f
C887 B.n169 VSUBS 0.006567f
C888 B.n170 VSUBS 0.006567f
C889 B.n171 VSUBS 0.006567f
C890 B.n172 VSUBS 0.006567f
C891 B.n173 VSUBS 0.006567f
C892 B.n174 VSUBS 0.006567f
C893 B.n175 VSUBS 0.006567f
C894 B.n176 VSUBS 0.006567f
C895 B.n177 VSUBS 0.006567f
C896 B.n178 VSUBS 0.006567f
C897 B.n179 VSUBS 0.006567f
C898 B.n180 VSUBS 0.006567f
C899 B.n181 VSUBS 0.006567f
C900 B.n182 VSUBS 0.016709f
C901 B.n183 VSUBS 0.006567f
C902 B.n184 VSUBS 0.006567f
C903 B.n185 VSUBS 0.006567f
C904 B.n186 VSUBS 0.006567f
C905 B.n187 VSUBS 0.006567f
C906 B.n188 VSUBS 0.006567f
C907 B.n189 VSUBS 0.006567f
C908 B.n190 VSUBS 0.006567f
C909 B.n191 VSUBS 0.006567f
C910 B.n192 VSUBS 0.006567f
C911 B.n193 VSUBS 0.006567f
C912 B.n194 VSUBS 0.006567f
C913 B.n195 VSUBS 0.006567f
C914 B.n196 VSUBS 0.006567f
C915 B.n197 VSUBS 0.006567f
C916 B.n198 VSUBS 0.006567f
C917 B.n199 VSUBS 0.006567f
C918 B.n200 VSUBS 0.006567f
C919 B.n201 VSUBS 0.006567f
C920 B.n202 VSUBS 0.006567f
C921 B.n203 VSUBS 0.006567f
C922 B.n204 VSUBS 0.006567f
C923 B.n205 VSUBS 0.006567f
C924 B.n206 VSUBS 0.006567f
C925 B.n207 VSUBS 0.006567f
C926 B.n208 VSUBS 0.006567f
C927 B.n209 VSUBS 0.006567f
C928 B.n210 VSUBS 0.006567f
C929 B.n211 VSUBS 0.006567f
C930 B.n212 VSUBS 0.006567f
C931 B.n213 VSUBS 0.006567f
C932 B.n214 VSUBS 0.006567f
C933 B.n215 VSUBS 0.006567f
C934 B.n216 VSUBS 0.006567f
C935 B.n217 VSUBS 0.006567f
C936 B.n218 VSUBS 0.006567f
C937 B.n219 VSUBS 0.006567f
C938 B.n220 VSUBS 0.006567f
C939 B.n221 VSUBS 0.006567f
C940 B.n222 VSUBS 0.006567f
C941 B.n223 VSUBS 0.006567f
C942 B.n224 VSUBS 0.006567f
C943 B.n225 VSUBS 0.006567f
C944 B.n226 VSUBS 0.006567f
C945 B.n227 VSUBS 0.006567f
C946 B.n228 VSUBS 0.006567f
C947 B.n229 VSUBS 0.006567f
C948 B.n230 VSUBS 0.006567f
C949 B.n231 VSUBS 0.006567f
C950 B.n232 VSUBS 0.006567f
C951 B.n233 VSUBS 0.006567f
C952 B.n234 VSUBS 0.006567f
C953 B.n235 VSUBS 0.006567f
C954 B.n236 VSUBS 0.006567f
C955 B.n237 VSUBS 0.006567f
C956 B.n238 VSUBS 0.006567f
C957 B.n239 VSUBS 0.006567f
C958 B.n240 VSUBS 0.006567f
C959 B.n241 VSUBS 0.006567f
C960 B.n242 VSUBS 0.006567f
C961 B.n243 VSUBS 0.006567f
C962 B.n244 VSUBS 0.006567f
C963 B.n245 VSUBS 0.006567f
C964 B.n246 VSUBS 0.006567f
C965 B.n247 VSUBS 0.006567f
C966 B.n248 VSUBS 0.006567f
C967 B.n249 VSUBS 0.006567f
C968 B.n250 VSUBS 0.006567f
C969 B.n251 VSUBS 0.006567f
C970 B.n252 VSUBS 0.006567f
C971 B.n253 VSUBS 0.006567f
C972 B.n254 VSUBS 0.006567f
C973 B.n255 VSUBS 0.006567f
C974 B.n256 VSUBS 0.006567f
C975 B.n257 VSUBS 0.006567f
C976 B.n258 VSUBS 0.006567f
C977 B.n259 VSUBS 0.006567f
C978 B.n260 VSUBS 0.006567f
C979 B.n261 VSUBS 0.006567f
C980 B.n262 VSUBS 0.006567f
C981 B.n263 VSUBS 0.006567f
C982 B.n264 VSUBS 0.006567f
C983 B.n265 VSUBS 0.006567f
C984 B.n266 VSUBS 0.006567f
C985 B.n267 VSUBS 0.015931f
C986 B.n268 VSUBS 0.015931f
C987 B.n269 VSUBS 0.016709f
C988 B.n270 VSUBS 0.006567f
C989 B.n271 VSUBS 0.006567f
C990 B.n272 VSUBS 0.006567f
C991 B.n273 VSUBS 0.006567f
C992 B.n274 VSUBS 0.006567f
C993 B.n275 VSUBS 0.006567f
C994 B.n276 VSUBS 0.006567f
C995 B.n277 VSUBS 0.006567f
C996 B.n278 VSUBS 0.006567f
C997 B.n279 VSUBS 0.006567f
C998 B.n280 VSUBS 0.006567f
C999 B.n281 VSUBS 0.006567f
C1000 B.n282 VSUBS 0.006567f
C1001 B.n283 VSUBS 0.006567f
C1002 B.n284 VSUBS 0.006567f
C1003 B.n285 VSUBS 0.006567f
C1004 B.n286 VSUBS 0.006567f
C1005 B.n287 VSUBS 0.006567f
C1006 B.n288 VSUBS 0.006567f
C1007 B.n289 VSUBS 0.006567f
C1008 B.n290 VSUBS 0.006567f
C1009 B.n291 VSUBS 0.006567f
C1010 B.n292 VSUBS 0.006567f
C1011 B.n293 VSUBS 0.006567f
C1012 B.n294 VSUBS 0.006567f
C1013 B.n295 VSUBS 0.006567f
C1014 B.n296 VSUBS 0.006567f
C1015 B.n297 VSUBS 0.006567f
C1016 B.n298 VSUBS 0.006567f
C1017 B.n299 VSUBS 0.006567f
C1018 B.n300 VSUBS 0.006567f
C1019 B.n301 VSUBS 0.006567f
C1020 B.n302 VSUBS 0.006567f
C1021 B.n303 VSUBS 0.006567f
C1022 B.n304 VSUBS 0.006567f
C1023 B.n305 VSUBS 0.006567f
C1024 B.n306 VSUBS 0.006567f
C1025 B.n307 VSUBS 0.006567f
C1026 B.n308 VSUBS 0.006567f
C1027 B.n309 VSUBS 0.006567f
C1028 B.n310 VSUBS 0.006567f
C1029 B.n311 VSUBS 0.006567f
C1030 B.n312 VSUBS 0.006567f
C1031 B.n313 VSUBS 0.006567f
C1032 B.n314 VSUBS 0.006567f
C1033 B.n315 VSUBS 0.006567f
C1034 B.n316 VSUBS 0.006567f
C1035 B.n317 VSUBS 0.006567f
C1036 B.n318 VSUBS 0.006567f
C1037 B.n319 VSUBS 0.006567f
C1038 B.n320 VSUBS 0.006567f
C1039 B.n321 VSUBS 0.006567f
C1040 B.n322 VSUBS 0.006567f
C1041 B.n323 VSUBS 0.006567f
C1042 B.n324 VSUBS 0.006567f
C1043 B.n325 VSUBS 0.006567f
C1044 B.n326 VSUBS 0.006567f
C1045 B.n327 VSUBS 0.006567f
C1046 B.n328 VSUBS 0.006567f
C1047 B.n329 VSUBS 0.006567f
C1048 B.n330 VSUBS 0.006567f
C1049 B.n331 VSUBS 0.006567f
C1050 B.n332 VSUBS 0.006567f
C1051 B.n333 VSUBS 0.006567f
C1052 B.n334 VSUBS 0.006567f
C1053 B.n335 VSUBS 0.006567f
C1054 B.n336 VSUBS 0.006567f
C1055 B.n337 VSUBS 0.006567f
C1056 B.n338 VSUBS 0.006567f
C1057 B.n339 VSUBS 0.004539f
C1058 B.n340 VSUBS 0.006567f
C1059 B.n341 VSUBS 0.006567f
C1060 B.n342 VSUBS 0.005311f
C1061 B.n343 VSUBS 0.006567f
C1062 B.n344 VSUBS 0.006567f
C1063 B.n345 VSUBS 0.006567f
C1064 B.n346 VSUBS 0.006567f
C1065 B.n347 VSUBS 0.006567f
C1066 B.n348 VSUBS 0.006567f
C1067 B.n349 VSUBS 0.006567f
C1068 B.n350 VSUBS 0.006567f
C1069 B.n351 VSUBS 0.006567f
C1070 B.n352 VSUBS 0.006567f
C1071 B.n353 VSUBS 0.006567f
C1072 B.n354 VSUBS 0.005311f
C1073 B.n355 VSUBS 0.015214f
C1074 B.n356 VSUBS 0.004539f
C1075 B.n357 VSUBS 0.006567f
C1076 B.n358 VSUBS 0.006567f
C1077 B.n359 VSUBS 0.006567f
C1078 B.n360 VSUBS 0.006567f
C1079 B.n361 VSUBS 0.006567f
C1080 B.n362 VSUBS 0.006567f
C1081 B.n363 VSUBS 0.006567f
C1082 B.n364 VSUBS 0.006567f
C1083 B.n365 VSUBS 0.006567f
C1084 B.n366 VSUBS 0.006567f
C1085 B.n367 VSUBS 0.006567f
C1086 B.n368 VSUBS 0.006567f
C1087 B.n369 VSUBS 0.006567f
C1088 B.n370 VSUBS 0.006567f
C1089 B.n371 VSUBS 0.006567f
C1090 B.n372 VSUBS 0.006567f
C1091 B.n373 VSUBS 0.006567f
C1092 B.n374 VSUBS 0.006567f
C1093 B.n375 VSUBS 0.006567f
C1094 B.n376 VSUBS 0.006567f
C1095 B.n377 VSUBS 0.006567f
C1096 B.n378 VSUBS 0.006567f
C1097 B.n379 VSUBS 0.006567f
C1098 B.n380 VSUBS 0.006567f
C1099 B.n381 VSUBS 0.006567f
C1100 B.n382 VSUBS 0.006567f
C1101 B.n383 VSUBS 0.006567f
C1102 B.n384 VSUBS 0.006567f
C1103 B.n385 VSUBS 0.006567f
C1104 B.n386 VSUBS 0.006567f
C1105 B.n387 VSUBS 0.006567f
C1106 B.n388 VSUBS 0.006567f
C1107 B.n389 VSUBS 0.006567f
C1108 B.n390 VSUBS 0.006567f
C1109 B.n391 VSUBS 0.006567f
C1110 B.n392 VSUBS 0.006567f
C1111 B.n393 VSUBS 0.006567f
C1112 B.n394 VSUBS 0.006567f
C1113 B.n395 VSUBS 0.006567f
C1114 B.n396 VSUBS 0.006567f
C1115 B.n397 VSUBS 0.006567f
C1116 B.n398 VSUBS 0.006567f
C1117 B.n399 VSUBS 0.006567f
C1118 B.n400 VSUBS 0.006567f
C1119 B.n401 VSUBS 0.006567f
C1120 B.n402 VSUBS 0.006567f
C1121 B.n403 VSUBS 0.006567f
C1122 B.n404 VSUBS 0.006567f
C1123 B.n405 VSUBS 0.006567f
C1124 B.n406 VSUBS 0.006567f
C1125 B.n407 VSUBS 0.006567f
C1126 B.n408 VSUBS 0.006567f
C1127 B.n409 VSUBS 0.006567f
C1128 B.n410 VSUBS 0.006567f
C1129 B.n411 VSUBS 0.006567f
C1130 B.n412 VSUBS 0.006567f
C1131 B.n413 VSUBS 0.006567f
C1132 B.n414 VSUBS 0.006567f
C1133 B.n415 VSUBS 0.006567f
C1134 B.n416 VSUBS 0.006567f
C1135 B.n417 VSUBS 0.006567f
C1136 B.n418 VSUBS 0.006567f
C1137 B.n419 VSUBS 0.006567f
C1138 B.n420 VSUBS 0.006567f
C1139 B.n421 VSUBS 0.006567f
C1140 B.n422 VSUBS 0.006567f
C1141 B.n423 VSUBS 0.006567f
C1142 B.n424 VSUBS 0.006567f
C1143 B.n425 VSUBS 0.006567f
C1144 B.n426 VSUBS 0.016709f
C1145 B.n427 VSUBS 0.016709f
C1146 B.n428 VSUBS 0.015931f
C1147 B.n429 VSUBS 0.006567f
C1148 B.n430 VSUBS 0.006567f
C1149 B.n431 VSUBS 0.006567f
C1150 B.n432 VSUBS 0.006567f
C1151 B.n433 VSUBS 0.006567f
C1152 B.n434 VSUBS 0.006567f
C1153 B.n435 VSUBS 0.006567f
C1154 B.n436 VSUBS 0.006567f
C1155 B.n437 VSUBS 0.006567f
C1156 B.n438 VSUBS 0.006567f
C1157 B.n439 VSUBS 0.006567f
C1158 B.n440 VSUBS 0.006567f
C1159 B.n441 VSUBS 0.006567f
C1160 B.n442 VSUBS 0.006567f
C1161 B.n443 VSUBS 0.006567f
C1162 B.n444 VSUBS 0.006567f
C1163 B.n445 VSUBS 0.006567f
C1164 B.n446 VSUBS 0.006567f
C1165 B.n447 VSUBS 0.006567f
C1166 B.n448 VSUBS 0.006567f
C1167 B.n449 VSUBS 0.006567f
C1168 B.n450 VSUBS 0.006567f
C1169 B.n451 VSUBS 0.006567f
C1170 B.n452 VSUBS 0.006567f
C1171 B.n453 VSUBS 0.006567f
C1172 B.n454 VSUBS 0.006567f
C1173 B.n455 VSUBS 0.006567f
C1174 B.n456 VSUBS 0.006567f
C1175 B.n457 VSUBS 0.006567f
C1176 B.n458 VSUBS 0.006567f
C1177 B.n459 VSUBS 0.006567f
C1178 B.n460 VSUBS 0.006567f
C1179 B.n461 VSUBS 0.006567f
C1180 B.n462 VSUBS 0.006567f
C1181 B.n463 VSUBS 0.006567f
C1182 B.n464 VSUBS 0.006567f
C1183 B.n465 VSUBS 0.006567f
C1184 B.n466 VSUBS 0.006567f
C1185 B.n467 VSUBS 0.006567f
C1186 B.n468 VSUBS 0.006567f
C1187 B.n469 VSUBS 0.006567f
C1188 B.n470 VSUBS 0.006567f
C1189 B.n471 VSUBS 0.006567f
C1190 B.n472 VSUBS 0.006567f
C1191 B.n473 VSUBS 0.006567f
C1192 B.n474 VSUBS 0.006567f
C1193 B.n475 VSUBS 0.006567f
C1194 B.n476 VSUBS 0.006567f
C1195 B.n477 VSUBS 0.006567f
C1196 B.n478 VSUBS 0.006567f
C1197 B.n479 VSUBS 0.006567f
C1198 B.n480 VSUBS 0.006567f
C1199 B.n481 VSUBS 0.006567f
C1200 B.n482 VSUBS 0.006567f
C1201 B.n483 VSUBS 0.006567f
C1202 B.n484 VSUBS 0.006567f
C1203 B.n485 VSUBS 0.006567f
C1204 B.n486 VSUBS 0.006567f
C1205 B.n487 VSUBS 0.006567f
C1206 B.n488 VSUBS 0.006567f
C1207 B.n489 VSUBS 0.006567f
C1208 B.n490 VSUBS 0.006567f
C1209 B.n491 VSUBS 0.006567f
C1210 B.n492 VSUBS 0.006567f
C1211 B.n493 VSUBS 0.006567f
C1212 B.n494 VSUBS 0.006567f
C1213 B.n495 VSUBS 0.006567f
C1214 B.n496 VSUBS 0.006567f
C1215 B.n497 VSUBS 0.006567f
C1216 B.n498 VSUBS 0.006567f
C1217 B.n499 VSUBS 0.006567f
C1218 B.n500 VSUBS 0.006567f
C1219 B.n501 VSUBS 0.006567f
C1220 B.n502 VSUBS 0.006567f
C1221 B.n503 VSUBS 0.006567f
C1222 B.n504 VSUBS 0.006567f
C1223 B.n505 VSUBS 0.006567f
C1224 B.n506 VSUBS 0.006567f
C1225 B.n507 VSUBS 0.006567f
C1226 B.n508 VSUBS 0.006567f
C1227 B.n509 VSUBS 0.006567f
C1228 B.n510 VSUBS 0.006567f
C1229 B.n511 VSUBS 0.006567f
C1230 B.n512 VSUBS 0.006567f
C1231 B.n513 VSUBS 0.006567f
C1232 B.n514 VSUBS 0.006567f
C1233 B.n515 VSUBS 0.006567f
C1234 B.n516 VSUBS 0.006567f
C1235 B.n517 VSUBS 0.006567f
C1236 B.n518 VSUBS 0.006567f
C1237 B.n519 VSUBS 0.006567f
C1238 B.n520 VSUBS 0.006567f
C1239 B.n521 VSUBS 0.006567f
C1240 B.n522 VSUBS 0.006567f
C1241 B.n523 VSUBS 0.006567f
C1242 B.n524 VSUBS 0.006567f
C1243 B.n525 VSUBS 0.006567f
C1244 B.n526 VSUBS 0.006567f
C1245 B.n527 VSUBS 0.006567f
C1246 B.n528 VSUBS 0.006567f
C1247 B.n529 VSUBS 0.006567f
C1248 B.n530 VSUBS 0.006567f
C1249 B.n531 VSUBS 0.006567f
C1250 B.n532 VSUBS 0.006567f
C1251 B.n533 VSUBS 0.006567f
C1252 B.n534 VSUBS 0.006567f
C1253 B.n535 VSUBS 0.006567f
C1254 B.n536 VSUBS 0.006567f
C1255 B.n537 VSUBS 0.006567f
C1256 B.n538 VSUBS 0.006567f
C1257 B.n539 VSUBS 0.006567f
C1258 B.n540 VSUBS 0.006567f
C1259 B.n541 VSUBS 0.006567f
C1260 B.n542 VSUBS 0.006567f
C1261 B.n543 VSUBS 0.006567f
C1262 B.n544 VSUBS 0.006567f
C1263 B.n545 VSUBS 0.006567f
C1264 B.n546 VSUBS 0.006567f
C1265 B.n547 VSUBS 0.006567f
C1266 B.n548 VSUBS 0.006567f
C1267 B.n549 VSUBS 0.006567f
C1268 B.n550 VSUBS 0.006567f
C1269 B.n551 VSUBS 0.006567f
C1270 B.n552 VSUBS 0.006567f
C1271 B.n553 VSUBS 0.006567f
C1272 B.n554 VSUBS 0.006567f
C1273 B.n555 VSUBS 0.006567f
C1274 B.n556 VSUBS 0.006567f
C1275 B.n557 VSUBS 0.006567f
C1276 B.n558 VSUBS 0.006567f
C1277 B.n559 VSUBS 0.006567f
C1278 B.n560 VSUBS 0.01664f
C1279 B.n561 VSUBS 0.016f
C1280 B.n562 VSUBS 0.016709f
C1281 B.n563 VSUBS 0.006567f
C1282 B.n564 VSUBS 0.006567f
C1283 B.n565 VSUBS 0.006567f
C1284 B.n566 VSUBS 0.006567f
C1285 B.n567 VSUBS 0.006567f
C1286 B.n568 VSUBS 0.006567f
C1287 B.n569 VSUBS 0.006567f
C1288 B.n570 VSUBS 0.006567f
C1289 B.n571 VSUBS 0.006567f
C1290 B.n572 VSUBS 0.006567f
C1291 B.n573 VSUBS 0.006567f
C1292 B.n574 VSUBS 0.006567f
C1293 B.n575 VSUBS 0.006567f
C1294 B.n576 VSUBS 0.006567f
C1295 B.n577 VSUBS 0.006567f
C1296 B.n578 VSUBS 0.006567f
C1297 B.n579 VSUBS 0.006567f
C1298 B.n580 VSUBS 0.006567f
C1299 B.n581 VSUBS 0.006567f
C1300 B.n582 VSUBS 0.006567f
C1301 B.n583 VSUBS 0.006567f
C1302 B.n584 VSUBS 0.006567f
C1303 B.n585 VSUBS 0.006567f
C1304 B.n586 VSUBS 0.006567f
C1305 B.n587 VSUBS 0.006567f
C1306 B.n588 VSUBS 0.006567f
C1307 B.n589 VSUBS 0.006567f
C1308 B.n590 VSUBS 0.006567f
C1309 B.n591 VSUBS 0.006567f
C1310 B.n592 VSUBS 0.006567f
C1311 B.n593 VSUBS 0.006567f
C1312 B.n594 VSUBS 0.006567f
C1313 B.n595 VSUBS 0.006567f
C1314 B.n596 VSUBS 0.006567f
C1315 B.n597 VSUBS 0.006567f
C1316 B.n598 VSUBS 0.006567f
C1317 B.n599 VSUBS 0.006567f
C1318 B.n600 VSUBS 0.006567f
C1319 B.n601 VSUBS 0.006567f
C1320 B.n602 VSUBS 0.006567f
C1321 B.n603 VSUBS 0.006567f
C1322 B.n604 VSUBS 0.006567f
C1323 B.n605 VSUBS 0.006567f
C1324 B.n606 VSUBS 0.006567f
C1325 B.n607 VSUBS 0.006567f
C1326 B.n608 VSUBS 0.006567f
C1327 B.n609 VSUBS 0.006567f
C1328 B.n610 VSUBS 0.006567f
C1329 B.n611 VSUBS 0.006567f
C1330 B.n612 VSUBS 0.006567f
C1331 B.n613 VSUBS 0.006567f
C1332 B.n614 VSUBS 0.006567f
C1333 B.n615 VSUBS 0.006567f
C1334 B.n616 VSUBS 0.006567f
C1335 B.n617 VSUBS 0.006567f
C1336 B.n618 VSUBS 0.006567f
C1337 B.n619 VSUBS 0.006567f
C1338 B.n620 VSUBS 0.006567f
C1339 B.n621 VSUBS 0.006567f
C1340 B.n622 VSUBS 0.006567f
C1341 B.n623 VSUBS 0.006567f
C1342 B.n624 VSUBS 0.006567f
C1343 B.n625 VSUBS 0.006567f
C1344 B.n626 VSUBS 0.006567f
C1345 B.n627 VSUBS 0.006567f
C1346 B.n628 VSUBS 0.006567f
C1347 B.n629 VSUBS 0.006567f
C1348 B.n630 VSUBS 0.006567f
C1349 B.n631 VSUBS 0.006567f
C1350 B.n632 VSUBS 0.004539f
C1351 B.n633 VSUBS 0.015214f
C1352 B.n634 VSUBS 0.005311f
C1353 B.n635 VSUBS 0.006567f
C1354 B.n636 VSUBS 0.006567f
C1355 B.n637 VSUBS 0.006567f
C1356 B.n638 VSUBS 0.006567f
C1357 B.n639 VSUBS 0.006567f
C1358 B.n640 VSUBS 0.006567f
C1359 B.n641 VSUBS 0.006567f
C1360 B.n642 VSUBS 0.006567f
C1361 B.n643 VSUBS 0.006567f
C1362 B.n644 VSUBS 0.006567f
C1363 B.n645 VSUBS 0.006567f
C1364 B.n646 VSUBS 0.005311f
C1365 B.n647 VSUBS 0.006567f
C1366 B.n648 VSUBS 0.006567f
C1367 B.n649 VSUBS 0.004539f
C1368 B.n650 VSUBS 0.006567f
C1369 B.n651 VSUBS 0.006567f
C1370 B.n652 VSUBS 0.006567f
C1371 B.n653 VSUBS 0.006567f
C1372 B.n654 VSUBS 0.006567f
C1373 B.n655 VSUBS 0.006567f
C1374 B.n656 VSUBS 0.006567f
C1375 B.n657 VSUBS 0.006567f
C1376 B.n658 VSUBS 0.006567f
C1377 B.n659 VSUBS 0.006567f
C1378 B.n660 VSUBS 0.006567f
C1379 B.n661 VSUBS 0.006567f
C1380 B.n662 VSUBS 0.006567f
C1381 B.n663 VSUBS 0.006567f
C1382 B.n664 VSUBS 0.006567f
C1383 B.n665 VSUBS 0.006567f
C1384 B.n666 VSUBS 0.006567f
C1385 B.n667 VSUBS 0.006567f
C1386 B.n668 VSUBS 0.006567f
C1387 B.n669 VSUBS 0.006567f
C1388 B.n670 VSUBS 0.006567f
C1389 B.n671 VSUBS 0.006567f
C1390 B.n672 VSUBS 0.006567f
C1391 B.n673 VSUBS 0.006567f
C1392 B.n674 VSUBS 0.006567f
C1393 B.n675 VSUBS 0.006567f
C1394 B.n676 VSUBS 0.006567f
C1395 B.n677 VSUBS 0.006567f
C1396 B.n678 VSUBS 0.006567f
C1397 B.n679 VSUBS 0.006567f
C1398 B.n680 VSUBS 0.006567f
C1399 B.n681 VSUBS 0.006567f
C1400 B.n682 VSUBS 0.006567f
C1401 B.n683 VSUBS 0.006567f
C1402 B.n684 VSUBS 0.006567f
C1403 B.n685 VSUBS 0.006567f
C1404 B.n686 VSUBS 0.006567f
C1405 B.n687 VSUBS 0.006567f
C1406 B.n688 VSUBS 0.006567f
C1407 B.n689 VSUBS 0.006567f
C1408 B.n690 VSUBS 0.006567f
C1409 B.n691 VSUBS 0.006567f
C1410 B.n692 VSUBS 0.006567f
C1411 B.n693 VSUBS 0.006567f
C1412 B.n694 VSUBS 0.006567f
C1413 B.n695 VSUBS 0.006567f
C1414 B.n696 VSUBS 0.006567f
C1415 B.n697 VSUBS 0.006567f
C1416 B.n698 VSUBS 0.006567f
C1417 B.n699 VSUBS 0.006567f
C1418 B.n700 VSUBS 0.006567f
C1419 B.n701 VSUBS 0.006567f
C1420 B.n702 VSUBS 0.006567f
C1421 B.n703 VSUBS 0.006567f
C1422 B.n704 VSUBS 0.006567f
C1423 B.n705 VSUBS 0.006567f
C1424 B.n706 VSUBS 0.006567f
C1425 B.n707 VSUBS 0.006567f
C1426 B.n708 VSUBS 0.006567f
C1427 B.n709 VSUBS 0.006567f
C1428 B.n710 VSUBS 0.006567f
C1429 B.n711 VSUBS 0.006567f
C1430 B.n712 VSUBS 0.006567f
C1431 B.n713 VSUBS 0.006567f
C1432 B.n714 VSUBS 0.006567f
C1433 B.n715 VSUBS 0.006567f
C1434 B.n716 VSUBS 0.006567f
C1435 B.n717 VSUBS 0.006567f
C1436 B.n718 VSUBS 0.006567f
C1437 B.n719 VSUBS 0.016709f
C1438 B.n720 VSUBS 0.015931f
C1439 B.n721 VSUBS 0.015931f
C1440 B.n722 VSUBS 0.006567f
C1441 B.n723 VSUBS 0.006567f
C1442 B.n724 VSUBS 0.006567f
C1443 B.n725 VSUBS 0.006567f
C1444 B.n726 VSUBS 0.006567f
C1445 B.n727 VSUBS 0.006567f
C1446 B.n728 VSUBS 0.006567f
C1447 B.n729 VSUBS 0.006567f
C1448 B.n730 VSUBS 0.006567f
C1449 B.n731 VSUBS 0.006567f
C1450 B.n732 VSUBS 0.006567f
C1451 B.n733 VSUBS 0.006567f
C1452 B.n734 VSUBS 0.006567f
C1453 B.n735 VSUBS 0.006567f
C1454 B.n736 VSUBS 0.006567f
C1455 B.n737 VSUBS 0.006567f
C1456 B.n738 VSUBS 0.006567f
C1457 B.n739 VSUBS 0.006567f
C1458 B.n740 VSUBS 0.006567f
C1459 B.n741 VSUBS 0.006567f
C1460 B.n742 VSUBS 0.006567f
C1461 B.n743 VSUBS 0.006567f
C1462 B.n744 VSUBS 0.006567f
C1463 B.n745 VSUBS 0.006567f
C1464 B.n746 VSUBS 0.006567f
C1465 B.n747 VSUBS 0.006567f
C1466 B.n748 VSUBS 0.006567f
C1467 B.n749 VSUBS 0.006567f
C1468 B.n750 VSUBS 0.006567f
C1469 B.n751 VSUBS 0.006567f
C1470 B.n752 VSUBS 0.006567f
C1471 B.n753 VSUBS 0.006567f
C1472 B.n754 VSUBS 0.006567f
C1473 B.n755 VSUBS 0.006567f
C1474 B.n756 VSUBS 0.006567f
C1475 B.n757 VSUBS 0.006567f
C1476 B.n758 VSUBS 0.006567f
C1477 B.n759 VSUBS 0.006567f
C1478 B.n760 VSUBS 0.006567f
C1479 B.n761 VSUBS 0.006567f
C1480 B.n762 VSUBS 0.006567f
C1481 B.n763 VSUBS 0.006567f
C1482 B.n764 VSUBS 0.006567f
C1483 B.n765 VSUBS 0.006567f
C1484 B.n766 VSUBS 0.006567f
C1485 B.n767 VSUBS 0.006567f
C1486 B.n768 VSUBS 0.006567f
C1487 B.n769 VSUBS 0.006567f
C1488 B.n770 VSUBS 0.006567f
C1489 B.n771 VSUBS 0.006567f
C1490 B.n772 VSUBS 0.006567f
C1491 B.n773 VSUBS 0.006567f
C1492 B.n774 VSUBS 0.006567f
C1493 B.n775 VSUBS 0.006567f
C1494 B.n776 VSUBS 0.006567f
C1495 B.n777 VSUBS 0.006567f
C1496 B.n778 VSUBS 0.006567f
C1497 B.n779 VSUBS 0.006567f
C1498 B.n780 VSUBS 0.006567f
C1499 B.n781 VSUBS 0.006567f
C1500 B.n782 VSUBS 0.006567f
C1501 B.n783 VSUBS 0.006567f
C1502 B.n784 VSUBS 0.006567f
C1503 B.n785 VSUBS 0.006567f
C1504 B.n786 VSUBS 0.006567f
C1505 B.n787 VSUBS 0.014869f
.ends

