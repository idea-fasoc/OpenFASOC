* NGSPICE file created from diff_pair_sample_1308.ext - technology: sky130A

.subckt diff_pair_sample_1308 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=1.75725 ps=10.98 w=10.65 l=0.33
X1 VDD1.t5 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=1.75725 ps=10.98 w=10.65 l=0.33
X2 VTAIL.t5 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=1.75725 ps=10.98 w=10.65 l=0.33
X3 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=1.75725 ps=10.98 w=10.65 l=0.33
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=0 ps=0 w=10.65 l=0.33
X5 VDD2.t4 VN.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=1.75725 ps=10.98 w=10.65 l=0.33
X6 VTAIL.t8 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=1.75725 ps=10.98 w=10.65 l=0.33
X7 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=1.75725 ps=10.98 w=10.65 l=0.33
X8 VDD2.t2 VN.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=4.1535 ps=22.08 w=10.65 l=0.33
X9 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=4.1535 ps=22.08 w=10.65 l=0.33
X10 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=0 ps=0 w=10.65 l=0.33
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=0 ps=0 w=10.65 l=0.33
X12 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=4.1535 ps=22.08 w=10.65 l=0.33
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.1535 pd=22.08 as=0 ps=0 w=10.65 l=0.33
X14 VTAIL.t9 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=1.75725 ps=10.98 w=10.65 l=0.33
X15 VDD2.t0 VN.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.75725 pd=10.98 as=4.1535 ps=22.08 w=10.65 l=0.33
R0 VN.n0 VN.t0 926.609
R1 VN.n4 VN.t3 926.609
R2 VN.n2 VN.t5 896.812
R3 VN.n6 VN.t1 896.812
R4 VN.n1 VN.t2 873.442
R5 VN.n5 VN.t4 873.442
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 73.0308
R9 VN.n6 VN.n5 73.0308
R10 VN.n7 VN.n4 65.9987
R11 VN.n3 VN.n0 65.9987
R12 VN VN.n7 39.116
R13 VN.n5 VN.n4 29.7615
R14 VN.n1 VN.n0 29.7615
R15 VN VN.n3 0.0516364
R16 VTAIL.n234 VTAIL.n182 289.615
R17 VTAIL.n54 VTAIL.n2 289.615
R18 VTAIL.n176 VTAIL.n124 289.615
R19 VTAIL.n116 VTAIL.n64 289.615
R20 VTAIL.n201 VTAIL.n200 185
R21 VTAIL.n198 VTAIL.n197 185
R22 VTAIL.n207 VTAIL.n206 185
R23 VTAIL.n209 VTAIL.n208 185
R24 VTAIL.n194 VTAIL.n193 185
R25 VTAIL.n215 VTAIL.n214 185
R26 VTAIL.n218 VTAIL.n217 185
R27 VTAIL.n216 VTAIL.n190 185
R28 VTAIL.n223 VTAIL.n189 185
R29 VTAIL.n225 VTAIL.n224 185
R30 VTAIL.n227 VTAIL.n226 185
R31 VTAIL.n186 VTAIL.n185 185
R32 VTAIL.n233 VTAIL.n232 185
R33 VTAIL.n235 VTAIL.n234 185
R34 VTAIL.n21 VTAIL.n20 185
R35 VTAIL.n18 VTAIL.n17 185
R36 VTAIL.n27 VTAIL.n26 185
R37 VTAIL.n29 VTAIL.n28 185
R38 VTAIL.n14 VTAIL.n13 185
R39 VTAIL.n35 VTAIL.n34 185
R40 VTAIL.n38 VTAIL.n37 185
R41 VTAIL.n36 VTAIL.n10 185
R42 VTAIL.n43 VTAIL.n9 185
R43 VTAIL.n45 VTAIL.n44 185
R44 VTAIL.n47 VTAIL.n46 185
R45 VTAIL.n6 VTAIL.n5 185
R46 VTAIL.n53 VTAIL.n52 185
R47 VTAIL.n55 VTAIL.n54 185
R48 VTAIL.n177 VTAIL.n176 185
R49 VTAIL.n175 VTAIL.n174 185
R50 VTAIL.n128 VTAIL.n127 185
R51 VTAIL.n169 VTAIL.n168 185
R52 VTAIL.n167 VTAIL.n166 185
R53 VTAIL.n165 VTAIL.n131 185
R54 VTAIL.n135 VTAIL.n132 185
R55 VTAIL.n160 VTAIL.n159 185
R56 VTAIL.n158 VTAIL.n157 185
R57 VTAIL.n137 VTAIL.n136 185
R58 VTAIL.n152 VTAIL.n151 185
R59 VTAIL.n150 VTAIL.n149 185
R60 VTAIL.n141 VTAIL.n140 185
R61 VTAIL.n144 VTAIL.n143 185
R62 VTAIL.n117 VTAIL.n116 185
R63 VTAIL.n115 VTAIL.n114 185
R64 VTAIL.n68 VTAIL.n67 185
R65 VTAIL.n109 VTAIL.n108 185
R66 VTAIL.n107 VTAIL.n106 185
R67 VTAIL.n105 VTAIL.n71 185
R68 VTAIL.n75 VTAIL.n72 185
R69 VTAIL.n100 VTAIL.n99 185
R70 VTAIL.n98 VTAIL.n97 185
R71 VTAIL.n77 VTAIL.n76 185
R72 VTAIL.n92 VTAIL.n91 185
R73 VTAIL.n90 VTAIL.n89 185
R74 VTAIL.n81 VTAIL.n80 185
R75 VTAIL.n84 VTAIL.n83 185
R76 VTAIL.t6 VTAIL.n199 149.524
R77 VTAIL.t3 VTAIL.n19 149.524
R78 VTAIL.t2 VTAIL.n142 149.524
R79 VTAIL.t11 VTAIL.n82 149.524
R80 VTAIL.n200 VTAIL.n197 104.615
R81 VTAIL.n207 VTAIL.n197 104.615
R82 VTAIL.n208 VTAIL.n207 104.615
R83 VTAIL.n208 VTAIL.n193 104.615
R84 VTAIL.n215 VTAIL.n193 104.615
R85 VTAIL.n217 VTAIL.n215 104.615
R86 VTAIL.n217 VTAIL.n216 104.615
R87 VTAIL.n216 VTAIL.n189 104.615
R88 VTAIL.n225 VTAIL.n189 104.615
R89 VTAIL.n226 VTAIL.n225 104.615
R90 VTAIL.n226 VTAIL.n185 104.615
R91 VTAIL.n233 VTAIL.n185 104.615
R92 VTAIL.n234 VTAIL.n233 104.615
R93 VTAIL.n20 VTAIL.n17 104.615
R94 VTAIL.n27 VTAIL.n17 104.615
R95 VTAIL.n28 VTAIL.n27 104.615
R96 VTAIL.n28 VTAIL.n13 104.615
R97 VTAIL.n35 VTAIL.n13 104.615
R98 VTAIL.n37 VTAIL.n35 104.615
R99 VTAIL.n37 VTAIL.n36 104.615
R100 VTAIL.n36 VTAIL.n9 104.615
R101 VTAIL.n45 VTAIL.n9 104.615
R102 VTAIL.n46 VTAIL.n45 104.615
R103 VTAIL.n46 VTAIL.n5 104.615
R104 VTAIL.n53 VTAIL.n5 104.615
R105 VTAIL.n54 VTAIL.n53 104.615
R106 VTAIL.n176 VTAIL.n175 104.615
R107 VTAIL.n175 VTAIL.n127 104.615
R108 VTAIL.n168 VTAIL.n127 104.615
R109 VTAIL.n168 VTAIL.n167 104.615
R110 VTAIL.n167 VTAIL.n131 104.615
R111 VTAIL.n135 VTAIL.n131 104.615
R112 VTAIL.n159 VTAIL.n135 104.615
R113 VTAIL.n159 VTAIL.n158 104.615
R114 VTAIL.n158 VTAIL.n136 104.615
R115 VTAIL.n151 VTAIL.n136 104.615
R116 VTAIL.n151 VTAIL.n150 104.615
R117 VTAIL.n150 VTAIL.n140 104.615
R118 VTAIL.n143 VTAIL.n140 104.615
R119 VTAIL.n116 VTAIL.n115 104.615
R120 VTAIL.n115 VTAIL.n67 104.615
R121 VTAIL.n108 VTAIL.n67 104.615
R122 VTAIL.n108 VTAIL.n107 104.615
R123 VTAIL.n107 VTAIL.n71 104.615
R124 VTAIL.n75 VTAIL.n71 104.615
R125 VTAIL.n99 VTAIL.n75 104.615
R126 VTAIL.n99 VTAIL.n98 104.615
R127 VTAIL.n98 VTAIL.n76 104.615
R128 VTAIL.n91 VTAIL.n76 104.615
R129 VTAIL.n91 VTAIL.n90 104.615
R130 VTAIL.n90 VTAIL.n80 104.615
R131 VTAIL.n83 VTAIL.n80 104.615
R132 VTAIL.n200 VTAIL.t6 52.3082
R133 VTAIL.n20 VTAIL.t3 52.3082
R134 VTAIL.n143 VTAIL.t2 52.3082
R135 VTAIL.n83 VTAIL.t11 52.3082
R136 VTAIL.n123 VTAIL.n122 45.0797
R137 VTAIL.n63 VTAIL.n62 45.0797
R138 VTAIL.n1 VTAIL.n0 45.0795
R139 VTAIL.n61 VTAIL.n60 45.0795
R140 VTAIL.n239 VTAIL.n238 31.6035
R141 VTAIL.n59 VTAIL.n58 31.6035
R142 VTAIL.n181 VTAIL.n180 31.6035
R143 VTAIL.n121 VTAIL.n120 31.6035
R144 VTAIL.n63 VTAIL.n61 22.6858
R145 VTAIL.n239 VTAIL.n181 22.1169
R146 VTAIL.n224 VTAIL.n223 13.1884
R147 VTAIL.n44 VTAIL.n43 13.1884
R148 VTAIL.n166 VTAIL.n165 13.1884
R149 VTAIL.n106 VTAIL.n105 13.1884
R150 VTAIL.n222 VTAIL.n190 12.8005
R151 VTAIL.n227 VTAIL.n188 12.8005
R152 VTAIL.n42 VTAIL.n10 12.8005
R153 VTAIL.n47 VTAIL.n8 12.8005
R154 VTAIL.n169 VTAIL.n130 12.8005
R155 VTAIL.n164 VTAIL.n132 12.8005
R156 VTAIL.n109 VTAIL.n70 12.8005
R157 VTAIL.n104 VTAIL.n72 12.8005
R158 VTAIL.n219 VTAIL.n218 12.0247
R159 VTAIL.n228 VTAIL.n186 12.0247
R160 VTAIL.n39 VTAIL.n38 12.0247
R161 VTAIL.n48 VTAIL.n6 12.0247
R162 VTAIL.n170 VTAIL.n128 12.0247
R163 VTAIL.n161 VTAIL.n160 12.0247
R164 VTAIL.n110 VTAIL.n68 12.0247
R165 VTAIL.n101 VTAIL.n100 12.0247
R166 VTAIL.n214 VTAIL.n192 11.249
R167 VTAIL.n232 VTAIL.n231 11.249
R168 VTAIL.n34 VTAIL.n12 11.249
R169 VTAIL.n52 VTAIL.n51 11.249
R170 VTAIL.n174 VTAIL.n173 11.249
R171 VTAIL.n157 VTAIL.n134 11.249
R172 VTAIL.n114 VTAIL.n113 11.249
R173 VTAIL.n97 VTAIL.n74 11.249
R174 VTAIL.n213 VTAIL.n194 10.4732
R175 VTAIL.n235 VTAIL.n184 10.4732
R176 VTAIL.n33 VTAIL.n14 10.4732
R177 VTAIL.n55 VTAIL.n4 10.4732
R178 VTAIL.n177 VTAIL.n126 10.4732
R179 VTAIL.n156 VTAIL.n137 10.4732
R180 VTAIL.n117 VTAIL.n66 10.4732
R181 VTAIL.n96 VTAIL.n77 10.4732
R182 VTAIL.n201 VTAIL.n199 10.2747
R183 VTAIL.n21 VTAIL.n19 10.2747
R184 VTAIL.n144 VTAIL.n142 10.2747
R185 VTAIL.n84 VTAIL.n82 10.2747
R186 VTAIL.n210 VTAIL.n209 9.69747
R187 VTAIL.n236 VTAIL.n182 9.69747
R188 VTAIL.n30 VTAIL.n29 9.69747
R189 VTAIL.n56 VTAIL.n2 9.69747
R190 VTAIL.n178 VTAIL.n124 9.69747
R191 VTAIL.n153 VTAIL.n152 9.69747
R192 VTAIL.n118 VTAIL.n64 9.69747
R193 VTAIL.n93 VTAIL.n92 9.69747
R194 VTAIL.n238 VTAIL.n237 9.45567
R195 VTAIL.n58 VTAIL.n57 9.45567
R196 VTAIL.n180 VTAIL.n179 9.45567
R197 VTAIL.n120 VTAIL.n119 9.45567
R198 VTAIL.n237 VTAIL.n236 9.3005
R199 VTAIL.n184 VTAIL.n183 9.3005
R200 VTAIL.n231 VTAIL.n230 9.3005
R201 VTAIL.n229 VTAIL.n228 9.3005
R202 VTAIL.n188 VTAIL.n187 9.3005
R203 VTAIL.n203 VTAIL.n202 9.3005
R204 VTAIL.n205 VTAIL.n204 9.3005
R205 VTAIL.n196 VTAIL.n195 9.3005
R206 VTAIL.n211 VTAIL.n210 9.3005
R207 VTAIL.n213 VTAIL.n212 9.3005
R208 VTAIL.n192 VTAIL.n191 9.3005
R209 VTAIL.n220 VTAIL.n219 9.3005
R210 VTAIL.n222 VTAIL.n221 9.3005
R211 VTAIL.n57 VTAIL.n56 9.3005
R212 VTAIL.n4 VTAIL.n3 9.3005
R213 VTAIL.n51 VTAIL.n50 9.3005
R214 VTAIL.n49 VTAIL.n48 9.3005
R215 VTAIL.n8 VTAIL.n7 9.3005
R216 VTAIL.n23 VTAIL.n22 9.3005
R217 VTAIL.n25 VTAIL.n24 9.3005
R218 VTAIL.n16 VTAIL.n15 9.3005
R219 VTAIL.n31 VTAIL.n30 9.3005
R220 VTAIL.n33 VTAIL.n32 9.3005
R221 VTAIL.n12 VTAIL.n11 9.3005
R222 VTAIL.n40 VTAIL.n39 9.3005
R223 VTAIL.n42 VTAIL.n41 9.3005
R224 VTAIL.n146 VTAIL.n145 9.3005
R225 VTAIL.n148 VTAIL.n147 9.3005
R226 VTAIL.n139 VTAIL.n138 9.3005
R227 VTAIL.n154 VTAIL.n153 9.3005
R228 VTAIL.n156 VTAIL.n155 9.3005
R229 VTAIL.n134 VTAIL.n133 9.3005
R230 VTAIL.n162 VTAIL.n161 9.3005
R231 VTAIL.n164 VTAIL.n163 9.3005
R232 VTAIL.n179 VTAIL.n178 9.3005
R233 VTAIL.n126 VTAIL.n125 9.3005
R234 VTAIL.n173 VTAIL.n172 9.3005
R235 VTAIL.n171 VTAIL.n170 9.3005
R236 VTAIL.n130 VTAIL.n129 9.3005
R237 VTAIL.n86 VTAIL.n85 9.3005
R238 VTAIL.n88 VTAIL.n87 9.3005
R239 VTAIL.n79 VTAIL.n78 9.3005
R240 VTAIL.n94 VTAIL.n93 9.3005
R241 VTAIL.n96 VTAIL.n95 9.3005
R242 VTAIL.n74 VTAIL.n73 9.3005
R243 VTAIL.n102 VTAIL.n101 9.3005
R244 VTAIL.n104 VTAIL.n103 9.3005
R245 VTAIL.n119 VTAIL.n118 9.3005
R246 VTAIL.n66 VTAIL.n65 9.3005
R247 VTAIL.n113 VTAIL.n112 9.3005
R248 VTAIL.n111 VTAIL.n110 9.3005
R249 VTAIL.n70 VTAIL.n69 9.3005
R250 VTAIL.n206 VTAIL.n196 8.92171
R251 VTAIL.n26 VTAIL.n16 8.92171
R252 VTAIL.n149 VTAIL.n139 8.92171
R253 VTAIL.n89 VTAIL.n79 8.92171
R254 VTAIL.n205 VTAIL.n198 8.14595
R255 VTAIL.n25 VTAIL.n18 8.14595
R256 VTAIL.n148 VTAIL.n141 8.14595
R257 VTAIL.n88 VTAIL.n81 8.14595
R258 VTAIL.n202 VTAIL.n201 7.3702
R259 VTAIL.n22 VTAIL.n21 7.3702
R260 VTAIL.n145 VTAIL.n144 7.3702
R261 VTAIL.n85 VTAIL.n84 7.3702
R262 VTAIL.n202 VTAIL.n198 5.81868
R263 VTAIL.n22 VTAIL.n18 5.81868
R264 VTAIL.n145 VTAIL.n141 5.81868
R265 VTAIL.n85 VTAIL.n81 5.81868
R266 VTAIL.n206 VTAIL.n205 5.04292
R267 VTAIL.n26 VTAIL.n25 5.04292
R268 VTAIL.n149 VTAIL.n148 5.04292
R269 VTAIL.n89 VTAIL.n88 5.04292
R270 VTAIL.n209 VTAIL.n196 4.26717
R271 VTAIL.n238 VTAIL.n182 4.26717
R272 VTAIL.n29 VTAIL.n16 4.26717
R273 VTAIL.n58 VTAIL.n2 4.26717
R274 VTAIL.n180 VTAIL.n124 4.26717
R275 VTAIL.n152 VTAIL.n139 4.26717
R276 VTAIL.n120 VTAIL.n64 4.26717
R277 VTAIL.n92 VTAIL.n79 4.26717
R278 VTAIL.n210 VTAIL.n194 3.49141
R279 VTAIL.n236 VTAIL.n235 3.49141
R280 VTAIL.n30 VTAIL.n14 3.49141
R281 VTAIL.n56 VTAIL.n55 3.49141
R282 VTAIL.n178 VTAIL.n177 3.49141
R283 VTAIL.n153 VTAIL.n137 3.49141
R284 VTAIL.n118 VTAIL.n117 3.49141
R285 VTAIL.n93 VTAIL.n77 3.49141
R286 VTAIL.n203 VTAIL.n199 2.84303
R287 VTAIL.n23 VTAIL.n19 2.84303
R288 VTAIL.n146 VTAIL.n142 2.84303
R289 VTAIL.n86 VTAIL.n82 2.84303
R290 VTAIL.n214 VTAIL.n213 2.71565
R291 VTAIL.n232 VTAIL.n184 2.71565
R292 VTAIL.n34 VTAIL.n33 2.71565
R293 VTAIL.n52 VTAIL.n4 2.71565
R294 VTAIL.n174 VTAIL.n126 2.71565
R295 VTAIL.n157 VTAIL.n156 2.71565
R296 VTAIL.n114 VTAIL.n66 2.71565
R297 VTAIL.n97 VTAIL.n96 2.71565
R298 VTAIL.n218 VTAIL.n192 1.93989
R299 VTAIL.n231 VTAIL.n186 1.93989
R300 VTAIL.n38 VTAIL.n12 1.93989
R301 VTAIL.n51 VTAIL.n6 1.93989
R302 VTAIL.n173 VTAIL.n128 1.93989
R303 VTAIL.n160 VTAIL.n134 1.93989
R304 VTAIL.n113 VTAIL.n68 1.93989
R305 VTAIL.n100 VTAIL.n74 1.93989
R306 VTAIL.n0 VTAIL.t7 1.85965
R307 VTAIL.n0 VTAIL.t8 1.85965
R308 VTAIL.n60 VTAIL.t0 1.85965
R309 VTAIL.n60 VTAIL.t5 1.85965
R310 VTAIL.n122 VTAIL.t4 1.85965
R311 VTAIL.n122 VTAIL.t1 1.85965
R312 VTAIL.n62 VTAIL.t10 1.85965
R313 VTAIL.n62 VTAIL.t9 1.85965
R314 VTAIL.n219 VTAIL.n190 1.16414
R315 VTAIL.n228 VTAIL.n227 1.16414
R316 VTAIL.n39 VTAIL.n10 1.16414
R317 VTAIL.n48 VTAIL.n47 1.16414
R318 VTAIL.n170 VTAIL.n169 1.16414
R319 VTAIL.n161 VTAIL.n132 1.16414
R320 VTAIL.n110 VTAIL.n109 1.16414
R321 VTAIL.n101 VTAIL.n72 1.16414
R322 VTAIL.n123 VTAIL.n121 0.75481
R323 VTAIL.n59 VTAIL.n1 0.75481
R324 VTAIL.n121 VTAIL.n63 0.569465
R325 VTAIL.n181 VTAIL.n123 0.569465
R326 VTAIL.n61 VTAIL.n59 0.569465
R327 VTAIL.n223 VTAIL.n222 0.388379
R328 VTAIL.n224 VTAIL.n188 0.388379
R329 VTAIL.n43 VTAIL.n42 0.388379
R330 VTAIL.n44 VTAIL.n8 0.388379
R331 VTAIL.n166 VTAIL.n130 0.388379
R332 VTAIL.n165 VTAIL.n164 0.388379
R333 VTAIL.n106 VTAIL.n70 0.388379
R334 VTAIL.n105 VTAIL.n104 0.388379
R335 VTAIL VTAIL.n239 0.369034
R336 VTAIL VTAIL.n1 0.200931
R337 VTAIL.n204 VTAIL.n203 0.155672
R338 VTAIL.n204 VTAIL.n195 0.155672
R339 VTAIL.n211 VTAIL.n195 0.155672
R340 VTAIL.n212 VTAIL.n211 0.155672
R341 VTAIL.n212 VTAIL.n191 0.155672
R342 VTAIL.n220 VTAIL.n191 0.155672
R343 VTAIL.n221 VTAIL.n220 0.155672
R344 VTAIL.n221 VTAIL.n187 0.155672
R345 VTAIL.n229 VTAIL.n187 0.155672
R346 VTAIL.n230 VTAIL.n229 0.155672
R347 VTAIL.n230 VTAIL.n183 0.155672
R348 VTAIL.n237 VTAIL.n183 0.155672
R349 VTAIL.n24 VTAIL.n23 0.155672
R350 VTAIL.n24 VTAIL.n15 0.155672
R351 VTAIL.n31 VTAIL.n15 0.155672
R352 VTAIL.n32 VTAIL.n31 0.155672
R353 VTAIL.n32 VTAIL.n11 0.155672
R354 VTAIL.n40 VTAIL.n11 0.155672
R355 VTAIL.n41 VTAIL.n40 0.155672
R356 VTAIL.n41 VTAIL.n7 0.155672
R357 VTAIL.n49 VTAIL.n7 0.155672
R358 VTAIL.n50 VTAIL.n49 0.155672
R359 VTAIL.n50 VTAIL.n3 0.155672
R360 VTAIL.n57 VTAIL.n3 0.155672
R361 VTAIL.n179 VTAIL.n125 0.155672
R362 VTAIL.n172 VTAIL.n125 0.155672
R363 VTAIL.n172 VTAIL.n171 0.155672
R364 VTAIL.n171 VTAIL.n129 0.155672
R365 VTAIL.n163 VTAIL.n129 0.155672
R366 VTAIL.n163 VTAIL.n162 0.155672
R367 VTAIL.n162 VTAIL.n133 0.155672
R368 VTAIL.n155 VTAIL.n133 0.155672
R369 VTAIL.n155 VTAIL.n154 0.155672
R370 VTAIL.n154 VTAIL.n138 0.155672
R371 VTAIL.n147 VTAIL.n138 0.155672
R372 VTAIL.n147 VTAIL.n146 0.155672
R373 VTAIL.n119 VTAIL.n65 0.155672
R374 VTAIL.n112 VTAIL.n65 0.155672
R375 VTAIL.n112 VTAIL.n111 0.155672
R376 VTAIL.n111 VTAIL.n69 0.155672
R377 VTAIL.n103 VTAIL.n69 0.155672
R378 VTAIL.n103 VTAIL.n102 0.155672
R379 VTAIL.n102 VTAIL.n73 0.155672
R380 VTAIL.n95 VTAIL.n73 0.155672
R381 VTAIL.n95 VTAIL.n94 0.155672
R382 VTAIL.n94 VTAIL.n78 0.155672
R383 VTAIL.n87 VTAIL.n78 0.155672
R384 VTAIL.n87 VTAIL.n86 0.155672
R385 VDD2.n111 VDD2.n59 289.615
R386 VDD2.n52 VDD2.n0 289.615
R387 VDD2.n112 VDD2.n111 185
R388 VDD2.n110 VDD2.n109 185
R389 VDD2.n63 VDD2.n62 185
R390 VDD2.n104 VDD2.n103 185
R391 VDD2.n102 VDD2.n101 185
R392 VDD2.n100 VDD2.n66 185
R393 VDD2.n70 VDD2.n67 185
R394 VDD2.n95 VDD2.n94 185
R395 VDD2.n93 VDD2.n92 185
R396 VDD2.n72 VDD2.n71 185
R397 VDD2.n87 VDD2.n86 185
R398 VDD2.n85 VDD2.n84 185
R399 VDD2.n76 VDD2.n75 185
R400 VDD2.n79 VDD2.n78 185
R401 VDD2.n19 VDD2.n18 185
R402 VDD2.n16 VDD2.n15 185
R403 VDD2.n25 VDD2.n24 185
R404 VDD2.n27 VDD2.n26 185
R405 VDD2.n12 VDD2.n11 185
R406 VDD2.n33 VDD2.n32 185
R407 VDD2.n36 VDD2.n35 185
R408 VDD2.n34 VDD2.n8 185
R409 VDD2.n41 VDD2.n7 185
R410 VDD2.n43 VDD2.n42 185
R411 VDD2.n45 VDD2.n44 185
R412 VDD2.n4 VDD2.n3 185
R413 VDD2.n51 VDD2.n50 185
R414 VDD2.n53 VDD2.n52 185
R415 VDD2.t4 VDD2.n77 149.524
R416 VDD2.t5 VDD2.n17 149.524
R417 VDD2.n111 VDD2.n110 104.615
R418 VDD2.n110 VDD2.n62 104.615
R419 VDD2.n103 VDD2.n62 104.615
R420 VDD2.n103 VDD2.n102 104.615
R421 VDD2.n102 VDD2.n66 104.615
R422 VDD2.n70 VDD2.n66 104.615
R423 VDD2.n94 VDD2.n70 104.615
R424 VDD2.n94 VDD2.n93 104.615
R425 VDD2.n93 VDD2.n71 104.615
R426 VDD2.n86 VDD2.n71 104.615
R427 VDD2.n86 VDD2.n85 104.615
R428 VDD2.n85 VDD2.n75 104.615
R429 VDD2.n78 VDD2.n75 104.615
R430 VDD2.n18 VDD2.n15 104.615
R431 VDD2.n25 VDD2.n15 104.615
R432 VDD2.n26 VDD2.n25 104.615
R433 VDD2.n26 VDD2.n11 104.615
R434 VDD2.n33 VDD2.n11 104.615
R435 VDD2.n35 VDD2.n33 104.615
R436 VDD2.n35 VDD2.n34 104.615
R437 VDD2.n34 VDD2.n7 104.615
R438 VDD2.n43 VDD2.n7 104.615
R439 VDD2.n44 VDD2.n43 104.615
R440 VDD2.n44 VDD2.n3 104.615
R441 VDD2.n51 VDD2.n3 104.615
R442 VDD2.n52 VDD2.n51 104.615
R443 VDD2.n58 VDD2.n57 61.8452
R444 VDD2 VDD2.n117 61.8424
R445 VDD2.n78 VDD2.t4 52.3082
R446 VDD2.n18 VDD2.t5 52.3082
R447 VDD2.n58 VDD2.n56 48.6537
R448 VDD2.n116 VDD2.n115 48.2823
R449 VDD2.n116 VDD2.n58 34.7455
R450 VDD2.n101 VDD2.n100 13.1884
R451 VDD2.n42 VDD2.n41 13.1884
R452 VDD2.n104 VDD2.n65 12.8005
R453 VDD2.n99 VDD2.n67 12.8005
R454 VDD2.n40 VDD2.n8 12.8005
R455 VDD2.n45 VDD2.n6 12.8005
R456 VDD2.n105 VDD2.n63 12.0247
R457 VDD2.n96 VDD2.n95 12.0247
R458 VDD2.n37 VDD2.n36 12.0247
R459 VDD2.n46 VDD2.n4 12.0247
R460 VDD2.n109 VDD2.n108 11.249
R461 VDD2.n92 VDD2.n69 11.249
R462 VDD2.n32 VDD2.n10 11.249
R463 VDD2.n50 VDD2.n49 11.249
R464 VDD2.n112 VDD2.n61 10.4732
R465 VDD2.n91 VDD2.n72 10.4732
R466 VDD2.n31 VDD2.n12 10.4732
R467 VDD2.n53 VDD2.n2 10.4732
R468 VDD2.n79 VDD2.n77 10.2747
R469 VDD2.n19 VDD2.n17 10.2747
R470 VDD2.n113 VDD2.n59 9.69747
R471 VDD2.n88 VDD2.n87 9.69747
R472 VDD2.n28 VDD2.n27 9.69747
R473 VDD2.n54 VDD2.n0 9.69747
R474 VDD2.n115 VDD2.n114 9.45567
R475 VDD2.n56 VDD2.n55 9.45567
R476 VDD2.n81 VDD2.n80 9.3005
R477 VDD2.n83 VDD2.n82 9.3005
R478 VDD2.n74 VDD2.n73 9.3005
R479 VDD2.n89 VDD2.n88 9.3005
R480 VDD2.n91 VDD2.n90 9.3005
R481 VDD2.n69 VDD2.n68 9.3005
R482 VDD2.n97 VDD2.n96 9.3005
R483 VDD2.n99 VDD2.n98 9.3005
R484 VDD2.n114 VDD2.n113 9.3005
R485 VDD2.n61 VDD2.n60 9.3005
R486 VDD2.n108 VDD2.n107 9.3005
R487 VDD2.n106 VDD2.n105 9.3005
R488 VDD2.n65 VDD2.n64 9.3005
R489 VDD2.n55 VDD2.n54 9.3005
R490 VDD2.n2 VDD2.n1 9.3005
R491 VDD2.n49 VDD2.n48 9.3005
R492 VDD2.n47 VDD2.n46 9.3005
R493 VDD2.n6 VDD2.n5 9.3005
R494 VDD2.n21 VDD2.n20 9.3005
R495 VDD2.n23 VDD2.n22 9.3005
R496 VDD2.n14 VDD2.n13 9.3005
R497 VDD2.n29 VDD2.n28 9.3005
R498 VDD2.n31 VDD2.n30 9.3005
R499 VDD2.n10 VDD2.n9 9.3005
R500 VDD2.n38 VDD2.n37 9.3005
R501 VDD2.n40 VDD2.n39 9.3005
R502 VDD2.n84 VDD2.n74 8.92171
R503 VDD2.n24 VDD2.n14 8.92171
R504 VDD2.n83 VDD2.n76 8.14595
R505 VDD2.n23 VDD2.n16 8.14595
R506 VDD2.n80 VDD2.n79 7.3702
R507 VDD2.n20 VDD2.n19 7.3702
R508 VDD2.n80 VDD2.n76 5.81868
R509 VDD2.n20 VDD2.n16 5.81868
R510 VDD2.n84 VDD2.n83 5.04292
R511 VDD2.n24 VDD2.n23 5.04292
R512 VDD2.n115 VDD2.n59 4.26717
R513 VDD2.n87 VDD2.n74 4.26717
R514 VDD2.n27 VDD2.n14 4.26717
R515 VDD2.n56 VDD2.n0 4.26717
R516 VDD2.n113 VDD2.n112 3.49141
R517 VDD2.n88 VDD2.n72 3.49141
R518 VDD2.n28 VDD2.n12 3.49141
R519 VDD2.n54 VDD2.n53 3.49141
R520 VDD2.n81 VDD2.n77 2.84303
R521 VDD2.n21 VDD2.n17 2.84303
R522 VDD2.n109 VDD2.n61 2.71565
R523 VDD2.n92 VDD2.n91 2.71565
R524 VDD2.n32 VDD2.n31 2.71565
R525 VDD2.n50 VDD2.n2 2.71565
R526 VDD2.n108 VDD2.n63 1.93989
R527 VDD2.n95 VDD2.n69 1.93989
R528 VDD2.n36 VDD2.n10 1.93989
R529 VDD2.n49 VDD2.n4 1.93989
R530 VDD2.n117 VDD2.t1 1.85965
R531 VDD2.n117 VDD2.t2 1.85965
R532 VDD2.n57 VDD2.t3 1.85965
R533 VDD2.n57 VDD2.t0 1.85965
R534 VDD2.n105 VDD2.n104 1.16414
R535 VDD2.n96 VDD2.n67 1.16414
R536 VDD2.n37 VDD2.n8 1.16414
R537 VDD2.n46 VDD2.n45 1.16414
R538 VDD2 VDD2.n116 0.485414
R539 VDD2.n101 VDD2.n65 0.388379
R540 VDD2.n100 VDD2.n99 0.388379
R541 VDD2.n41 VDD2.n40 0.388379
R542 VDD2.n42 VDD2.n6 0.388379
R543 VDD2.n114 VDD2.n60 0.155672
R544 VDD2.n107 VDD2.n60 0.155672
R545 VDD2.n107 VDD2.n106 0.155672
R546 VDD2.n106 VDD2.n64 0.155672
R547 VDD2.n98 VDD2.n64 0.155672
R548 VDD2.n98 VDD2.n97 0.155672
R549 VDD2.n97 VDD2.n68 0.155672
R550 VDD2.n90 VDD2.n68 0.155672
R551 VDD2.n90 VDD2.n89 0.155672
R552 VDD2.n89 VDD2.n73 0.155672
R553 VDD2.n82 VDD2.n73 0.155672
R554 VDD2.n82 VDD2.n81 0.155672
R555 VDD2.n22 VDD2.n21 0.155672
R556 VDD2.n22 VDD2.n13 0.155672
R557 VDD2.n29 VDD2.n13 0.155672
R558 VDD2.n30 VDD2.n29 0.155672
R559 VDD2.n30 VDD2.n9 0.155672
R560 VDD2.n38 VDD2.n9 0.155672
R561 VDD2.n39 VDD2.n38 0.155672
R562 VDD2.n39 VDD2.n5 0.155672
R563 VDD2.n47 VDD2.n5 0.155672
R564 VDD2.n48 VDD2.n47 0.155672
R565 VDD2.n48 VDD2.n1 0.155672
R566 VDD2.n55 VDD2.n1 0.155672
R567 B.n296 B.t13 990.389
R568 B.n394 B.t17 990.389
R569 B.n79 B.t6 990.389
R570 B.n77 B.t10 990.389
R571 B.n566 B.n565 585
R572 B.n567 B.n566 585
R573 B.n247 B.n76 585
R574 B.n246 B.n245 585
R575 B.n244 B.n243 585
R576 B.n242 B.n241 585
R577 B.n240 B.n239 585
R578 B.n238 B.n237 585
R579 B.n236 B.n235 585
R580 B.n234 B.n233 585
R581 B.n232 B.n231 585
R582 B.n230 B.n229 585
R583 B.n228 B.n227 585
R584 B.n226 B.n225 585
R585 B.n224 B.n223 585
R586 B.n222 B.n221 585
R587 B.n220 B.n219 585
R588 B.n218 B.n217 585
R589 B.n216 B.n215 585
R590 B.n214 B.n213 585
R591 B.n212 B.n211 585
R592 B.n210 B.n209 585
R593 B.n208 B.n207 585
R594 B.n206 B.n205 585
R595 B.n204 B.n203 585
R596 B.n202 B.n201 585
R597 B.n200 B.n199 585
R598 B.n198 B.n197 585
R599 B.n196 B.n195 585
R600 B.n194 B.n193 585
R601 B.n192 B.n191 585
R602 B.n190 B.n189 585
R603 B.n188 B.n187 585
R604 B.n186 B.n185 585
R605 B.n184 B.n183 585
R606 B.n182 B.n181 585
R607 B.n180 B.n179 585
R608 B.n178 B.n177 585
R609 B.n176 B.n175 585
R610 B.n173 B.n172 585
R611 B.n171 B.n170 585
R612 B.n169 B.n168 585
R613 B.n167 B.n166 585
R614 B.n165 B.n164 585
R615 B.n163 B.n162 585
R616 B.n161 B.n160 585
R617 B.n159 B.n158 585
R618 B.n157 B.n156 585
R619 B.n155 B.n154 585
R620 B.n153 B.n152 585
R621 B.n151 B.n150 585
R622 B.n149 B.n148 585
R623 B.n147 B.n146 585
R624 B.n145 B.n144 585
R625 B.n143 B.n142 585
R626 B.n141 B.n140 585
R627 B.n139 B.n138 585
R628 B.n137 B.n136 585
R629 B.n135 B.n134 585
R630 B.n133 B.n132 585
R631 B.n131 B.n130 585
R632 B.n129 B.n128 585
R633 B.n127 B.n126 585
R634 B.n125 B.n124 585
R635 B.n123 B.n122 585
R636 B.n121 B.n120 585
R637 B.n119 B.n118 585
R638 B.n117 B.n116 585
R639 B.n115 B.n114 585
R640 B.n113 B.n112 585
R641 B.n111 B.n110 585
R642 B.n109 B.n108 585
R643 B.n107 B.n106 585
R644 B.n105 B.n104 585
R645 B.n103 B.n102 585
R646 B.n101 B.n100 585
R647 B.n99 B.n98 585
R648 B.n97 B.n96 585
R649 B.n95 B.n94 585
R650 B.n93 B.n92 585
R651 B.n91 B.n90 585
R652 B.n89 B.n88 585
R653 B.n87 B.n86 585
R654 B.n85 B.n84 585
R655 B.n83 B.n82 585
R656 B.n32 B.n31 585
R657 B.n564 B.n33 585
R658 B.n568 B.n33 585
R659 B.n563 B.n562 585
R660 B.n562 B.n29 585
R661 B.n561 B.n28 585
R662 B.n574 B.n28 585
R663 B.n560 B.n27 585
R664 B.n575 B.n27 585
R665 B.n559 B.n26 585
R666 B.n576 B.n26 585
R667 B.n558 B.n557 585
R668 B.n557 B.n22 585
R669 B.n556 B.n21 585
R670 B.n582 B.n21 585
R671 B.n555 B.n20 585
R672 B.n583 B.n20 585
R673 B.n554 B.n19 585
R674 B.n584 B.n19 585
R675 B.n553 B.n552 585
R676 B.n552 B.n18 585
R677 B.n551 B.n14 585
R678 B.n590 B.n14 585
R679 B.n550 B.n13 585
R680 B.n591 B.n13 585
R681 B.n549 B.n12 585
R682 B.n592 B.n12 585
R683 B.n548 B.n547 585
R684 B.n547 B.n11 585
R685 B.n546 B.n7 585
R686 B.n598 B.n7 585
R687 B.n545 B.n6 585
R688 B.n599 B.n6 585
R689 B.n544 B.n5 585
R690 B.n600 B.n5 585
R691 B.n543 B.n542 585
R692 B.n542 B.n4 585
R693 B.n541 B.n248 585
R694 B.n541 B.n540 585
R695 B.n530 B.n249 585
R696 B.n533 B.n249 585
R697 B.n532 B.n531 585
R698 B.n534 B.n532 585
R699 B.n529 B.n253 585
R700 B.n256 B.n253 585
R701 B.n528 B.n527 585
R702 B.n527 B.n526 585
R703 B.n255 B.n254 585
R704 B.n519 B.n255 585
R705 B.n518 B.n517 585
R706 B.n520 B.n518 585
R707 B.n516 B.n261 585
R708 B.n261 B.n260 585
R709 B.n515 B.n514 585
R710 B.n514 B.n513 585
R711 B.n263 B.n262 585
R712 B.n264 B.n263 585
R713 B.n506 B.n505 585
R714 B.n507 B.n506 585
R715 B.n504 B.n269 585
R716 B.n269 B.n268 585
R717 B.n503 B.n502 585
R718 B.n502 B.n501 585
R719 B.n271 B.n270 585
R720 B.n272 B.n271 585
R721 B.n494 B.n493 585
R722 B.n495 B.n494 585
R723 B.n275 B.n274 585
R724 B.n324 B.n322 585
R725 B.n325 B.n321 585
R726 B.n325 B.n276 585
R727 B.n328 B.n327 585
R728 B.n329 B.n320 585
R729 B.n331 B.n330 585
R730 B.n333 B.n319 585
R731 B.n336 B.n335 585
R732 B.n337 B.n318 585
R733 B.n339 B.n338 585
R734 B.n341 B.n317 585
R735 B.n344 B.n343 585
R736 B.n345 B.n316 585
R737 B.n347 B.n346 585
R738 B.n349 B.n315 585
R739 B.n352 B.n351 585
R740 B.n353 B.n314 585
R741 B.n355 B.n354 585
R742 B.n357 B.n313 585
R743 B.n360 B.n359 585
R744 B.n361 B.n312 585
R745 B.n363 B.n362 585
R746 B.n365 B.n311 585
R747 B.n368 B.n367 585
R748 B.n369 B.n310 585
R749 B.n371 B.n370 585
R750 B.n373 B.n309 585
R751 B.n376 B.n375 585
R752 B.n377 B.n308 585
R753 B.n379 B.n378 585
R754 B.n381 B.n307 585
R755 B.n384 B.n383 585
R756 B.n385 B.n306 585
R757 B.n387 B.n386 585
R758 B.n389 B.n305 585
R759 B.n392 B.n391 585
R760 B.n393 B.n304 585
R761 B.n398 B.n397 585
R762 B.n400 B.n303 585
R763 B.n403 B.n402 585
R764 B.n404 B.n302 585
R765 B.n406 B.n405 585
R766 B.n408 B.n301 585
R767 B.n411 B.n410 585
R768 B.n412 B.n300 585
R769 B.n414 B.n413 585
R770 B.n416 B.n299 585
R771 B.n419 B.n418 585
R772 B.n420 B.n295 585
R773 B.n422 B.n421 585
R774 B.n424 B.n294 585
R775 B.n427 B.n426 585
R776 B.n428 B.n293 585
R777 B.n430 B.n429 585
R778 B.n432 B.n292 585
R779 B.n435 B.n434 585
R780 B.n436 B.n291 585
R781 B.n438 B.n437 585
R782 B.n440 B.n290 585
R783 B.n443 B.n442 585
R784 B.n444 B.n289 585
R785 B.n446 B.n445 585
R786 B.n448 B.n288 585
R787 B.n451 B.n450 585
R788 B.n452 B.n287 585
R789 B.n454 B.n453 585
R790 B.n456 B.n286 585
R791 B.n459 B.n458 585
R792 B.n460 B.n285 585
R793 B.n462 B.n461 585
R794 B.n464 B.n284 585
R795 B.n467 B.n466 585
R796 B.n468 B.n283 585
R797 B.n470 B.n469 585
R798 B.n472 B.n282 585
R799 B.n475 B.n474 585
R800 B.n476 B.n281 585
R801 B.n478 B.n477 585
R802 B.n480 B.n280 585
R803 B.n483 B.n482 585
R804 B.n484 B.n279 585
R805 B.n486 B.n485 585
R806 B.n488 B.n278 585
R807 B.n491 B.n490 585
R808 B.n492 B.n277 585
R809 B.n497 B.n496 585
R810 B.n496 B.n495 585
R811 B.n498 B.n273 585
R812 B.n273 B.n272 585
R813 B.n500 B.n499 585
R814 B.n501 B.n500 585
R815 B.n267 B.n266 585
R816 B.n268 B.n267 585
R817 B.n509 B.n508 585
R818 B.n508 B.n507 585
R819 B.n510 B.n265 585
R820 B.n265 B.n264 585
R821 B.n512 B.n511 585
R822 B.n513 B.n512 585
R823 B.n259 B.n258 585
R824 B.n260 B.n259 585
R825 B.n522 B.n521 585
R826 B.n521 B.n520 585
R827 B.n523 B.n257 585
R828 B.n519 B.n257 585
R829 B.n525 B.n524 585
R830 B.n526 B.n525 585
R831 B.n252 B.n251 585
R832 B.n256 B.n252 585
R833 B.n536 B.n535 585
R834 B.n535 B.n534 585
R835 B.n537 B.n250 585
R836 B.n533 B.n250 585
R837 B.n539 B.n538 585
R838 B.n540 B.n539 585
R839 B.n2 B.n0 585
R840 B.n4 B.n2 585
R841 B.n3 B.n1 585
R842 B.n599 B.n3 585
R843 B.n597 B.n596 585
R844 B.n598 B.n597 585
R845 B.n595 B.n8 585
R846 B.n11 B.n8 585
R847 B.n594 B.n593 585
R848 B.n593 B.n592 585
R849 B.n10 B.n9 585
R850 B.n591 B.n10 585
R851 B.n589 B.n588 585
R852 B.n590 B.n589 585
R853 B.n587 B.n15 585
R854 B.n18 B.n15 585
R855 B.n586 B.n585 585
R856 B.n585 B.n584 585
R857 B.n17 B.n16 585
R858 B.n583 B.n17 585
R859 B.n581 B.n580 585
R860 B.n582 B.n581 585
R861 B.n579 B.n23 585
R862 B.n23 B.n22 585
R863 B.n578 B.n577 585
R864 B.n577 B.n576 585
R865 B.n25 B.n24 585
R866 B.n575 B.n25 585
R867 B.n573 B.n572 585
R868 B.n574 B.n573 585
R869 B.n571 B.n30 585
R870 B.n30 B.n29 585
R871 B.n570 B.n569 585
R872 B.n569 B.n568 585
R873 B.n602 B.n601 585
R874 B.n601 B.n600 585
R875 B.n496 B.n275 468.476
R876 B.n569 B.n32 468.476
R877 B.n494 B.n277 468.476
R878 B.n566 B.n33 468.476
R879 B.n296 B.t16 271.577
R880 B.n77 B.t11 271.577
R881 B.n394 B.t19 271.577
R882 B.n79 B.t8 271.577
R883 B.n297 B.t15 258.777
R884 B.n78 B.t12 258.777
R885 B.n395 B.t18 258.777
R886 B.n80 B.t9 258.777
R887 B.n567 B.n75 256.663
R888 B.n567 B.n74 256.663
R889 B.n567 B.n73 256.663
R890 B.n567 B.n72 256.663
R891 B.n567 B.n71 256.663
R892 B.n567 B.n70 256.663
R893 B.n567 B.n69 256.663
R894 B.n567 B.n68 256.663
R895 B.n567 B.n67 256.663
R896 B.n567 B.n66 256.663
R897 B.n567 B.n65 256.663
R898 B.n567 B.n64 256.663
R899 B.n567 B.n63 256.663
R900 B.n567 B.n62 256.663
R901 B.n567 B.n61 256.663
R902 B.n567 B.n60 256.663
R903 B.n567 B.n59 256.663
R904 B.n567 B.n58 256.663
R905 B.n567 B.n57 256.663
R906 B.n567 B.n56 256.663
R907 B.n567 B.n55 256.663
R908 B.n567 B.n54 256.663
R909 B.n567 B.n53 256.663
R910 B.n567 B.n52 256.663
R911 B.n567 B.n51 256.663
R912 B.n567 B.n50 256.663
R913 B.n567 B.n49 256.663
R914 B.n567 B.n48 256.663
R915 B.n567 B.n47 256.663
R916 B.n567 B.n46 256.663
R917 B.n567 B.n45 256.663
R918 B.n567 B.n44 256.663
R919 B.n567 B.n43 256.663
R920 B.n567 B.n42 256.663
R921 B.n567 B.n41 256.663
R922 B.n567 B.n40 256.663
R923 B.n567 B.n39 256.663
R924 B.n567 B.n38 256.663
R925 B.n567 B.n37 256.663
R926 B.n567 B.n36 256.663
R927 B.n567 B.n35 256.663
R928 B.n567 B.n34 256.663
R929 B.n323 B.n276 256.663
R930 B.n326 B.n276 256.663
R931 B.n332 B.n276 256.663
R932 B.n334 B.n276 256.663
R933 B.n340 B.n276 256.663
R934 B.n342 B.n276 256.663
R935 B.n348 B.n276 256.663
R936 B.n350 B.n276 256.663
R937 B.n356 B.n276 256.663
R938 B.n358 B.n276 256.663
R939 B.n364 B.n276 256.663
R940 B.n366 B.n276 256.663
R941 B.n372 B.n276 256.663
R942 B.n374 B.n276 256.663
R943 B.n380 B.n276 256.663
R944 B.n382 B.n276 256.663
R945 B.n388 B.n276 256.663
R946 B.n390 B.n276 256.663
R947 B.n399 B.n276 256.663
R948 B.n401 B.n276 256.663
R949 B.n407 B.n276 256.663
R950 B.n409 B.n276 256.663
R951 B.n415 B.n276 256.663
R952 B.n417 B.n276 256.663
R953 B.n423 B.n276 256.663
R954 B.n425 B.n276 256.663
R955 B.n431 B.n276 256.663
R956 B.n433 B.n276 256.663
R957 B.n439 B.n276 256.663
R958 B.n441 B.n276 256.663
R959 B.n447 B.n276 256.663
R960 B.n449 B.n276 256.663
R961 B.n455 B.n276 256.663
R962 B.n457 B.n276 256.663
R963 B.n463 B.n276 256.663
R964 B.n465 B.n276 256.663
R965 B.n471 B.n276 256.663
R966 B.n473 B.n276 256.663
R967 B.n479 B.n276 256.663
R968 B.n481 B.n276 256.663
R969 B.n487 B.n276 256.663
R970 B.n489 B.n276 256.663
R971 B.n496 B.n273 163.367
R972 B.n500 B.n273 163.367
R973 B.n500 B.n267 163.367
R974 B.n508 B.n267 163.367
R975 B.n508 B.n265 163.367
R976 B.n512 B.n265 163.367
R977 B.n512 B.n259 163.367
R978 B.n521 B.n259 163.367
R979 B.n521 B.n257 163.367
R980 B.n525 B.n257 163.367
R981 B.n525 B.n252 163.367
R982 B.n535 B.n252 163.367
R983 B.n535 B.n250 163.367
R984 B.n539 B.n250 163.367
R985 B.n539 B.n2 163.367
R986 B.n601 B.n2 163.367
R987 B.n601 B.n3 163.367
R988 B.n597 B.n3 163.367
R989 B.n597 B.n8 163.367
R990 B.n593 B.n8 163.367
R991 B.n593 B.n10 163.367
R992 B.n589 B.n10 163.367
R993 B.n589 B.n15 163.367
R994 B.n585 B.n15 163.367
R995 B.n585 B.n17 163.367
R996 B.n581 B.n17 163.367
R997 B.n581 B.n23 163.367
R998 B.n577 B.n23 163.367
R999 B.n577 B.n25 163.367
R1000 B.n573 B.n25 163.367
R1001 B.n573 B.n30 163.367
R1002 B.n569 B.n30 163.367
R1003 B.n325 B.n324 163.367
R1004 B.n327 B.n325 163.367
R1005 B.n331 B.n320 163.367
R1006 B.n335 B.n333 163.367
R1007 B.n339 B.n318 163.367
R1008 B.n343 B.n341 163.367
R1009 B.n347 B.n316 163.367
R1010 B.n351 B.n349 163.367
R1011 B.n355 B.n314 163.367
R1012 B.n359 B.n357 163.367
R1013 B.n363 B.n312 163.367
R1014 B.n367 B.n365 163.367
R1015 B.n371 B.n310 163.367
R1016 B.n375 B.n373 163.367
R1017 B.n379 B.n308 163.367
R1018 B.n383 B.n381 163.367
R1019 B.n387 B.n306 163.367
R1020 B.n391 B.n389 163.367
R1021 B.n398 B.n304 163.367
R1022 B.n402 B.n400 163.367
R1023 B.n406 B.n302 163.367
R1024 B.n410 B.n408 163.367
R1025 B.n414 B.n300 163.367
R1026 B.n418 B.n416 163.367
R1027 B.n422 B.n295 163.367
R1028 B.n426 B.n424 163.367
R1029 B.n430 B.n293 163.367
R1030 B.n434 B.n432 163.367
R1031 B.n438 B.n291 163.367
R1032 B.n442 B.n440 163.367
R1033 B.n446 B.n289 163.367
R1034 B.n450 B.n448 163.367
R1035 B.n454 B.n287 163.367
R1036 B.n458 B.n456 163.367
R1037 B.n462 B.n285 163.367
R1038 B.n466 B.n464 163.367
R1039 B.n470 B.n283 163.367
R1040 B.n474 B.n472 163.367
R1041 B.n478 B.n281 163.367
R1042 B.n482 B.n480 163.367
R1043 B.n486 B.n279 163.367
R1044 B.n490 B.n488 163.367
R1045 B.n494 B.n271 163.367
R1046 B.n502 B.n271 163.367
R1047 B.n502 B.n269 163.367
R1048 B.n506 B.n269 163.367
R1049 B.n506 B.n263 163.367
R1050 B.n514 B.n263 163.367
R1051 B.n514 B.n261 163.367
R1052 B.n518 B.n261 163.367
R1053 B.n518 B.n255 163.367
R1054 B.n527 B.n255 163.367
R1055 B.n527 B.n253 163.367
R1056 B.n532 B.n253 163.367
R1057 B.n532 B.n249 163.367
R1058 B.n541 B.n249 163.367
R1059 B.n542 B.n541 163.367
R1060 B.n542 B.n5 163.367
R1061 B.n6 B.n5 163.367
R1062 B.n7 B.n6 163.367
R1063 B.n547 B.n7 163.367
R1064 B.n547 B.n12 163.367
R1065 B.n13 B.n12 163.367
R1066 B.n14 B.n13 163.367
R1067 B.n552 B.n14 163.367
R1068 B.n552 B.n19 163.367
R1069 B.n20 B.n19 163.367
R1070 B.n21 B.n20 163.367
R1071 B.n557 B.n21 163.367
R1072 B.n557 B.n26 163.367
R1073 B.n27 B.n26 163.367
R1074 B.n28 B.n27 163.367
R1075 B.n562 B.n28 163.367
R1076 B.n562 B.n33 163.367
R1077 B.n84 B.n83 163.367
R1078 B.n88 B.n87 163.367
R1079 B.n92 B.n91 163.367
R1080 B.n96 B.n95 163.367
R1081 B.n100 B.n99 163.367
R1082 B.n104 B.n103 163.367
R1083 B.n108 B.n107 163.367
R1084 B.n112 B.n111 163.367
R1085 B.n116 B.n115 163.367
R1086 B.n120 B.n119 163.367
R1087 B.n124 B.n123 163.367
R1088 B.n128 B.n127 163.367
R1089 B.n132 B.n131 163.367
R1090 B.n136 B.n135 163.367
R1091 B.n140 B.n139 163.367
R1092 B.n144 B.n143 163.367
R1093 B.n148 B.n147 163.367
R1094 B.n152 B.n151 163.367
R1095 B.n156 B.n155 163.367
R1096 B.n160 B.n159 163.367
R1097 B.n164 B.n163 163.367
R1098 B.n168 B.n167 163.367
R1099 B.n172 B.n171 163.367
R1100 B.n177 B.n176 163.367
R1101 B.n181 B.n180 163.367
R1102 B.n185 B.n184 163.367
R1103 B.n189 B.n188 163.367
R1104 B.n193 B.n192 163.367
R1105 B.n197 B.n196 163.367
R1106 B.n201 B.n200 163.367
R1107 B.n205 B.n204 163.367
R1108 B.n209 B.n208 163.367
R1109 B.n213 B.n212 163.367
R1110 B.n217 B.n216 163.367
R1111 B.n221 B.n220 163.367
R1112 B.n225 B.n224 163.367
R1113 B.n229 B.n228 163.367
R1114 B.n233 B.n232 163.367
R1115 B.n237 B.n236 163.367
R1116 B.n241 B.n240 163.367
R1117 B.n245 B.n244 163.367
R1118 B.n566 B.n76 163.367
R1119 B.n495 B.n276 79.4354
R1120 B.n568 B.n567 79.4354
R1121 B.n323 B.n275 71.676
R1122 B.n327 B.n326 71.676
R1123 B.n332 B.n331 71.676
R1124 B.n335 B.n334 71.676
R1125 B.n340 B.n339 71.676
R1126 B.n343 B.n342 71.676
R1127 B.n348 B.n347 71.676
R1128 B.n351 B.n350 71.676
R1129 B.n356 B.n355 71.676
R1130 B.n359 B.n358 71.676
R1131 B.n364 B.n363 71.676
R1132 B.n367 B.n366 71.676
R1133 B.n372 B.n371 71.676
R1134 B.n375 B.n374 71.676
R1135 B.n380 B.n379 71.676
R1136 B.n383 B.n382 71.676
R1137 B.n388 B.n387 71.676
R1138 B.n391 B.n390 71.676
R1139 B.n399 B.n398 71.676
R1140 B.n402 B.n401 71.676
R1141 B.n407 B.n406 71.676
R1142 B.n410 B.n409 71.676
R1143 B.n415 B.n414 71.676
R1144 B.n418 B.n417 71.676
R1145 B.n423 B.n422 71.676
R1146 B.n426 B.n425 71.676
R1147 B.n431 B.n430 71.676
R1148 B.n434 B.n433 71.676
R1149 B.n439 B.n438 71.676
R1150 B.n442 B.n441 71.676
R1151 B.n447 B.n446 71.676
R1152 B.n450 B.n449 71.676
R1153 B.n455 B.n454 71.676
R1154 B.n458 B.n457 71.676
R1155 B.n463 B.n462 71.676
R1156 B.n466 B.n465 71.676
R1157 B.n471 B.n470 71.676
R1158 B.n474 B.n473 71.676
R1159 B.n479 B.n478 71.676
R1160 B.n482 B.n481 71.676
R1161 B.n487 B.n486 71.676
R1162 B.n490 B.n489 71.676
R1163 B.n34 B.n32 71.676
R1164 B.n84 B.n35 71.676
R1165 B.n88 B.n36 71.676
R1166 B.n92 B.n37 71.676
R1167 B.n96 B.n38 71.676
R1168 B.n100 B.n39 71.676
R1169 B.n104 B.n40 71.676
R1170 B.n108 B.n41 71.676
R1171 B.n112 B.n42 71.676
R1172 B.n116 B.n43 71.676
R1173 B.n120 B.n44 71.676
R1174 B.n124 B.n45 71.676
R1175 B.n128 B.n46 71.676
R1176 B.n132 B.n47 71.676
R1177 B.n136 B.n48 71.676
R1178 B.n140 B.n49 71.676
R1179 B.n144 B.n50 71.676
R1180 B.n148 B.n51 71.676
R1181 B.n152 B.n52 71.676
R1182 B.n156 B.n53 71.676
R1183 B.n160 B.n54 71.676
R1184 B.n164 B.n55 71.676
R1185 B.n168 B.n56 71.676
R1186 B.n172 B.n57 71.676
R1187 B.n177 B.n58 71.676
R1188 B.n181 B.n59 71.676
R1189 B.n185 B.n60 71.676
R1190 B.n189 B.n61 71.676
R1191 B.n193 B.n62 71.676
R1192 B.n197 B.n63 71.676
R1193 B.n201 B.n64 71.676
R1194 B.n205 B.n65 71.676
R1195 B.n209 B.n66 71.676
R1196 B.n213 B.n67 71.676
R1197 B.n217 B.n68 71.676
R1198 B.n221 B.n69 71.676
R1199 B.n225 B.n70 71.676
R1200 B.n229 B.n71 71.676
R1201 B.n233 B.n72 71.676
R1202 B.n237 B.n73 71.676
R1203 B.n241 B.n74 71.676
R1204 B.n245 B.n75 71.676
R1205 B.n76 B.n75 71.676
R1206 B.n244 B.n74 71.676
R1207 B.n240 B.n73 71.676
R1208 B.n236 B.n72 71.676
R1209 B.n232 B.n71 71.676
R1210 B.n228 B.n70 71.676
R1211 B.n224 B.n69 71.676
R1212 B.n220 B.n68 71.676
R1213 B.n216 B.n67 71.676
R1214 B.n212 B.n66 71.676
R1215 B.n208 B.n65 71.676
R1216 B.n204 B.n64 71.676
R1217 B.n200 B.n63 71.676
R1218 B.n196 B.n62 71.676
R1219 B.n192 B.n61 71.676
R1220 B.n188 B.n60 71.676
R1221 B.n184 B.n59 71.676
R1222 B.n180 B.n58 71.676
R1223 B.n176 B.n57 71.676
R1224 B.n171 B.n56 71.676
R1225 B.n167 B.n55 71.676
R1226 B.n163 B.n54 71.676
R1227 B.n159 B.n53 71.676
R1228 B.n155 B.n52 71.676
R1229 B.n151 B.n51 71.676
R1230 B.n147 B.n50 71.676
R1231 B.n143 B.n49 71.676
R1232 B.n139 B.n48 71.676
R1233 B.n135 B.n47 71.676
R1234 B.n131 B.n46 71.676
R1235 B.n127 B.n45 71.676
R1236 B.n123 B.n44 71.676
R1237 B.n119 B.n43 71.676
R1238 B.n115 B.n42 71.676
R1239 B.n111 B.n41 71.676
R1240 B.n107 B.n40 71.676
R1241 B.n103 B.n39 71.676
R1242 B.n99 B.n38 71.676
R1243 B.n95 B.n37 71.676
R1244 B.n91 B.n36 71.676
R1245 B.n87 B.n35 71.676
R1246 B.n83 B.n34 71.676
R1247 B.n324 B.n323 71.676
R1248 B.n326 B.n320 71.676
R1249 B.n333 B.n332 71.676
R1250 B.n334 B.n318 71.676
R1251 B.n341 B.n340 71.676
R1252 B.n342 B.n316 71.676
R1253 B.n349 B.n348 71.676
R1254 B.n350 B.n314 71.676
R1255 B.n357 B.n356 71.676
R1256 B.n358 B.n312 71.676
R1257 B.n365 B.n364 71.676
R1258 B.n366 B.n310 71.676
R1259 B.n373 B.n372 71.676
R1260 B.n374 B.n308 71.676
R1261 B.n381 B.n380 71.676
R1262 B.n382 B.n306 71.676
R1263 B.n389 B.n388 71.676
R1264 B.n390 B.n304 71.676
R1265 B.n400 B.n399 71.676
R1266 B.n401 B.n302 71.676
R1267 B.n408 B.n407 71.676
R1268 B.n409 B.n300 71.676
R1269 B.n416 B.n415 71.676
R1270 B.n417 B.n295 71.676
R1271 B.n424 B.n423 71.676
R1272 B.n425 B.n293 71.676
R1273 B.n432 B.n431 71.676
R1274 B.n433 B.n291 71.676
R1275 B.n440 B.n439 71.676
R1276 B.n441 B.n289 71.676
R1277 B.n448 B.n447 71.676
R1278 B.n449 B.n287 71.676
R1279 B.n456 B.n455 71.676
R1280 B.n457 B.n285 71.676
R1281 B.n464 B.n463 71.676
R1282 B.n465 B.n283 71.676
R1283 B.n472 B.n471 71.676
R1284 B.n473 B.n281 71.676
R1285 B.n480 B.n479 71.676
R1286 B.n481 B.n279 71.676
R1287 B.n488 B.n487 71.676
R1288 B.n489 B.n277 71.676
R1289 B.n298 B.n297 59.5399
R1290 B.n396 B.n395 59.5399
R1291 B.n81 B.n80 59.5399
R1292 B.n174 B.n78 59.5399
R1293 B.n495 B.n272 46.9707
R1294 B.n501 B.n272 46.9707
R1295 B.n501 B.n268 46.9707
R1296 B.n507 B.n268 46.9707
R1297 B.n513 B.n264 46.9707
R1298 B.n513 B.n260 46.9707
R1299 B.n520 B.n260 46.9707
R1300 B.n520 B.n519 46.9707
R1301 B.n526 B.n256 46.9707
R1302 B.n534 B.n533 46.9707
R1303 B.n540 B.n4 46.9707
R1304 B.n600 B.n4 46.9707
R1305 B.n600 B.n599 46.9707
R1306 B.n599 B.n598 46.9707
R1307 B.n592 B.n11 46.9707
R1308 B.n591 B.n590 46.9707
R1309 B.n584 B.n18 46.9707
R1310 B.n584 B.n583 46.9707
R1311 B.n583 B.n582 46.9707
R1312 B.n582 B.n22 46.9707
R1313 B.n576 B.n575 46.9707
R1314 B.n575 B.n574 46.9707
R1315 B.n574 B.n29 46.9707
R1316 B.n568 B.n29 46.9707
R1317 B.n570 B.n31 30.4395
R1318 B.n565 B.n564 30.4395
R1319 B.n493 B.n492 30.4395
R1320 B.n497 B.n274 30.4395
R1321 B.t14 B.n264 28.3208
R1322 B.t7 B.n22 28.3208
R1323 B.n540 B.t3 26.9393
R1324 B.n598 B.t4 26.9393
R1325 B.n519 B.t0 25.5578
R1326 B.n18 B.t2 25.5578
R1327 B.n534 B.t5 24.1763
R1328 B.n592 B.t1 24.1763
R1329 B.n256 B.t5 22.7948
R1330 B.t1 B.n591 22.7948
R1331 B.n526 B.t0 21.4134
R1332 B.n590 B.t2 21.4134
R1333 B.n533 B.t3 20.0319
R1334 B.n11 B.t4 20.0319
R1335 B.n507 B.t14 18.6504
R1336 B.n576 B.t7 18.6504
R1337 B B.n602 18.0485
R1338 B.n297 B.n296 12.8005
R1339 B.n395 B.n394 12.8005
R1340 B.n80 B.n79 12.8005
R1341 B.n78 B.n77 12.8005
R1342 B.n82 B.n31 10.6151
R1343 B.n85 B.n82 10.6151
R1344 B.n86 B.n85 10.6151
R1345 B.n89 B.n86 10.6151
R1346 B.n90 B.n89 10.6151
R1347 B.n93 B.n90 10.6151
R1348 B.n94 B.n93 10.6151
R1349 B.n97 B.n94 10.6151
R1350 B.n98 B.n97 10.6151
R1351 B.n101 B.n98 10.6151
R1352 B.n102 B.n101 10.6151
R1353 B.n105 B.n102 10.6151
R1354 B.n106 B.n105 10.6151
R1355 B.n109 B.n106 10.6151
R1356 B.n110 B.n109 10.6151
R1357 B.n113 B.n110 10.6151
R1358 B.n114 B.n113 10.6151
R1359 B.n117 B.n114 10.6151
R1360 B.n118 B.n117 10.6151
R1361 B.n121 B.n118 10.6151
R1362 B.n122 B.n121 10.6151
R1363 B.n125 B.n122 10.6151
R1364 B.n126 B.n125 10.6151
R1365 B.n129 B.n126 10.6151
R1366 B.n130 B.n129 10.6151
R1367 B.n133 B.n130 10.6151
R1368 B.n134 B.n133 10.6151
R1369 B.n137 B.n134 10.6151
R1370 B.n138 B.n137 10.6151
R1371 B.n141 B.n138 10.6151
R1372 B.n142 B.n141 10.6151
R1373 B.n145 B.n142 10.6151
R1374 B.n146 B.n145 10.6151
R1375 B.n149 B.n146 10.6151
R1376 B.n150 B.n149 10.6151
R1377 B.n153 B.n150 10.6151
R1378 B.n154 B.n153 10.6151
R1379 B.n158 B.n157 10.6151
R1380 B.n161 B.n158 10.6151
R1381 B.n162 B.n161 10.6151
R1382 B.n165 B.n162 10.6151
R1383 B.n166 B.n165 10.6151
R1384 B.n169 B.n166 10.6151
R1385 B.n170 B.n169 10.6151
R1386 B.n173 B.n170 10.6151
R1387 B.n178 B.n175 10.6151
R1388 B.n179 B.n178 10.6151
R1389 B.n182 B.n179 10.6151
R1390 B.n183 B.n182 10.6151
R1391 B.n186 B.n183 10.6151
R1392 B.n187 B.n186 10.6151
R1393 B.n190 B.n187 10.6151
R1394 B.n191 B.n190 10.6151
R1395 B.n194 B.n191 10.6151
R1396 B.n195 B.n194 10.6151
R1397 B.n198 B.n195 10.6151
R1398 B.n199 B.n198 10.6151
R1399 B.n202 B.n199 10.6151
R1400 B.n203 B.n202 10.6151
R1401 B.n206 B.n203 10.6151
R1402 B.n207 B.n206 10.6151
R1403 B.n210 B.n207 10.6151
R1404 B.n211 B.n210 10.6151
R1405 B.n214 B.n211 10.6151
R1406 B.n215 B.n214 10.6151
R1407 B.n218 B.n215 10.6151
R1408 B.n219 B.n218 10.6151
R1409 B.n222 B.n219 10.6151
R1410 B.n223 B.n222 10.6151
R1411 B.n226 B.n223 10.6151
R1412 B.n227 B.n226 10.6151
R1413 B.n230 B.n227 10.6151
R1414 B.n231 B.n230 10.6151
R1415 B.n234 B.n231 10.6151
R1416 B.n235 B.n234 10.6151
R1417 B.n238 B.n235 10.6151
R1418 B.n239 B.n238 10.6151
R1419 B.n242 B.n239 10.6151
R1420 B.n243 B.n242 10.6151
R1421 B.n246 B.n243 10.6151
R1422 B.n247 B.n246 10.6151
R1423 B.n565 B.n247 10.6151
R1424 B.n493 B.n270 10.6151
R1425 B.n503 B.n270 10.6151
R1426 B.n504 B.n503 10.6151
R1427 B.n505 B.n504 10.6151
R1428 B.n505 B.n262 10.6151
R1429 B.n515 B.n262 10.6151
R1430 B.n516 B.n515 10.6151
R1431 B.n517 B.n516 10.6151
R1432 B.n517 B.n254 10.6151
R1433 B.n528 B.n254 10.6151
R1434 B.n529 B.n528 10.6151
R1435 B.n531 B.n529 10.6151
R1436 B.n531 B.n530 10.6151
R1437 B.n530 B.n248 10.6151
R1438 B.n543 B.n248 10.6151
R1439 B.n544 B.n543 10.6151
R1440 B.n545 B.n544 10.6151
R1441 B.n546 B.n545 10.6151
R1442 B.n548 B.n546 10.6151
R1443 B.n549 B.n548 10.6151
R1444 B.n550 B.n549 10.6151
R1445 B.n551 B.n550 10.6151
R1446 B.n553 B.n551 10.6151
R1447 B.n554 B.n553 10.6151
R1448 B.n555 B.n554 10.6151
R1449 B.n556 B.n555 10.6151
R1450 B.n558 B.n556 10.6151
R1451 B.n559 B.n558 10.6151
R1452 B.n560 B.n559 10.6151
R1453 B.n561 B.n560 10.6151
R1454 B.n563 B.n561 10.6151
R1455 B.n564 B.n563 10.6151
R1456 B.n322 B.n274 10.6151
R1457 B.n322 B.n321 10.6151
R1458 B.n328 B.n321 10.6151
R1459 B.n329 B.n328 10.6151
R1460 B.n330 B.n329 10.6151
R1461 B.n330 B.n319 10.6151
R1462 B.n336 B.n319 10.6151
R1463 B.n337 B.n336 10.6151
R1464 B.n338 B.n337 10.6151
R1465 B.n338 B.n317 10.6151
R1466 B.n344 B.n317 10.6151
R1467 B.n345 B.n344 10.6151
R1468 B.n346 B.n345 10.6151
R1469 B.n346 B.n315 10.6151
R1470 B.n352 B.n315 10.6151
R1471 B.n353 B.n352 10.6151
R1472 B.n354 B.n353 10.6151
R1473 B.n354 B.n313 10.6151
R1474 B.n360 B.n313 10.6151
R1475 B.n361 B.n360 10.6151
R1476 B.n362 B.n361 10.6151
R1477 B.n362 B.n311 10.6151
R1478 B.n368 B.n311 10.6151
R1479 B.n369 B.n368 10.6151
R1480 B.n370 B.n369 10.6151
R1481 B.n370 B.n309 10.6151
R1482 B.n376 B.n309 10.6151
R1483 B.n377 B.n376 10.6151
R1484 B.n378 B.n377 10.6151
R1485 B.n378 B.n307 10.6151
R1486 B.n384 B.n307 10.6151
R1487 B.n385 B.n384 10.6151
R1488 B.n386 B.n385 10.6151
R1489 B.n386 B.n305 10.6151
R1490 B.n392 B.n305 10.6151
R1491 B.n393 B.n392 10.6151
R1492 B.n397 B.n393 10.6151
R1493 B.n403 B.n303 10.6151
R1494 B.n404 B.n403 10.6151
R1495 B.n405 B.n404 10.6151
R1496 B.n405 B.n301 10.6151
R1497 B.n411 B.n301 10.6151
R1498 B.n412 B.n411 10.6151
R1499 B.n413 B.n412 10.6151
R1500 B.n413 B.n299 10.6151
R1501 B.n420 B.n419 10.6151
R1502 B.n421 B.n420 10.6151
R1503 B.n421 B.n294 10.6151
R1504 B.n427 B.n294 10.6151
R1505 B.n428 B.n427 10.6151
R1506 B.n429 B.n428 10.6151
R1507 B.n429 B.n292 10.6151
R1508 B.n435 B.n292 10.6151
R1509 B.n436 B.n435 10.6151
R1510 B.n437 B.n436 10.6151
R1511 B.n437 B.n290 10.6151
R1512 B.n443 B.n290 10.6151
R1513 B.n444 B.n443 10.6151
R1514 B.n445 B.n444 10.6151
R1515 B.n445 B.n288 10.6151
R1516 B.n451 B.n288 10.6151
R1517 B.n452 B.n451 10.6151
R1518 B.n453 B.n452 10.6151
R1519 B.n453 B.n286 10.6151
R1520 B.n459 B.n286 10.6151
R1521 B.n460 B.n459 10.6151
R1522 B.n461 B.n460 10.6151
R1523 B.n461 B.n284 10.6151
R1524 B.n467 B.n284 10.6151
R1525 B.n468 B.n467 10.6151
R1526 B.n469 B.n468 10.6151
R1527 B.n469 B.n282 10.6151
R1528 B.n475 B.n282 10.6151
R1529 B.n476 B.n475 10.6151
R1530 B.n477 B.n476 10.6151
R1531 B.n477 B.n280 10.6151
R1532 B.n483 B.n280 10.6151
R1533 B.n484 B.n483 10.6151
R1534 B.n485 B.n484 10.6151
R1535 B.n485 B.n278 10.6151
R1536 B.n491 B.n278 10.6151
R1537 B.n492 B.n491 10.6151
R1538 B.n498 B.n497 10.6151
R1539 B.n499 B.n498 10.6151
R1540 B.n499 B.n266 10.6151
R1541 B.n509 B.n266 10.6151
R1542 B.n510 B.n509 10.6151
R1543 B.n511 B.n510 10.6151
R1544 B.n511 B.n258 10.6151
R1545 B.n522 B.n258 10.6151
R1546 B.n523 B.n522 10.6151
R1547 B.n524 B.n523 10.6151
R1548 B.n524 B.n251 10.6151
R1549 B.n536 B.n251 10.6151
R1550 B.n537 B.n536 10.6151
R1551 B.n538 B.n537 10.6151
R1552 B.n538 B.n0 10.6151
R1553 B.n596 B.n1 10.6151
R1554 B.n596 B.n595 10.6151
R1555 B.n595 B.n594 10.6151
R1556 B.n594 B.n9 10.6151
R1557 B.n588 B.n9 10.6151
R1558 B.n588 B.n587 10.6151
R1559 B.n587 B.n586 10.6151
R1560 B.n586 B.n16 10.6151
R1561 B.n580 B.n16 10.6151
R1562 B.n580 B.n579 10.6151
R1563 B.n579 B.n578 10.6151
R1564 B.n578 B.n24 10.6151
R1565 B.n572 B.n24 10.6151
R1566 B.n572 B.n571 10.6151
R1567 B.n571 B.n570 10.6151
R1568 B.n157 B.n81 6.5566
R1569 B.n174 B.n173 6.5566
R1570 B.n396 B.n303 6.5566
R1571 B.n299 B.n298 6.5566
R1572 B.n154 B.n81 4.05904
R1573 B.n175 B.n174 4.05904
R1574 B.n397 B.n396 4.05904
R1575 B.n419 B.n298 4.05904
R1576 B.n602 B.n0 2.81026
R1577 B.n602 B.n1 2.81026
R1578 VP.n1 VP.t2 926.609
R1579 VP.n8 VP.t4 896.812
R1580 VP.n6 VP.t0 896.812
R1581 VP.n3 VP.t5 896.812
R1582 VP.n7 VP.t1 873.442
R1583 VP.n2 VP.t3 873.442
R1584 VP.n9 VP.n8 161.3
R1585 VP.n4 VP.n3 161.3
R1586 VP.n7 VP.n0 161.3
R1587 VP.n6 VP.n5 161.3
R1588 VP.n7 VP.n6 73.0308
R1589 VP.n8 VP.n7 73.0308
R1590 VP.n3 VP.n2 73.0308
R1591 VP.n4 VP.n1 65.9987
R1592 VP.n5 VP.n4 38.7353
R1593 VP.n2 VP.n1 29.7615
R1594 VP.n5 VP.n0 0.189894
R1595 VP.n9 VP.n0 0.189894
R1596 VP VP.n9 0.0516364
R1597 VDD1.n52 VDD1.n0 289.615
R1598 VDD1.n109 VDD1.n57 289.615
R1599 VDD1.n53 VDD1.n52 185
R1600 VDD1.n51 VDD1.n50 185
R1601 VDD1.n4 VDD1.n3 185
R1602 VDD1.n45 VDD1.n44 185
R1603 VDD1.n43 VDD1.n42 185
R1604 VDD1.n41 VDD1.n7 185
R1605 VDD1.n11 VDD1.n8 185
R1606 VDD1.n36 VDD1.n35 185
R1607 VDD1.n34 VDD1.n33 185
R1608 VDD1.n13 VDD1.n12 185
R1609 VDD1.n28 VDD1.n27 185
R1610 VDD1.n26 VDD1.n25 185
R1611 VDD1.n17 VDD1.n16 185
R1612 VDD1.n20 VDD1.n19 185
R1613 VDD1.n76 VDD1.n75 185
R1614 VDD1.n73 VDD1.n72 185
R1615 VDD1.n82 VDD1.n81 185
R1616 VDD1.n84 VDD1.n83 185
R1617 VDD1.n69 VDD1.n68 185
R1618 VDD1.n90 VDD1.n89 185
R1619 VDD1.n93 VDD1.n92 185
R1620 VDD1.n91 VDD1.n65 185
R1621 VDD1.n98 VDD1.n64 185
R1622 VDD1.n100 VDD1.n99 185
R1623 VDD1.n102 VDD1.n101 185
R1624 VDD1.n61 VDD1.n60 185
R1625 VDD1.n108 VDD1.n107 185
R1626 VDD1.n110 VDD1.n109 185
R1627 VDD1.t3 VDD1.n18 149.524
R1628 VDD1.t5 VDD1.n74 149.524
R1629 VDD1.n52 VDD1.n51 104.615
R1630 VDD1.n51 VDD1.n3 104.615
R1631 VDD1.n44 VDD1.n3 104.615
R1632 VDD1.n44 VDD1.n43 104.615
R1633 VDD1.n43 VDD1.n7 104.615
R1634 VDD1.n11 VDD1.n7 104.615
R1635 VDD1.n35 VDD1.n11 104.615
R1636 VDD1.n35 VDD1.n34 104.615
R1637 VDD1.n34 VDD1.n12 104.615
R1638 VDD1.n27 VDD1.n12 104.615
R1639 VDD1.n27 VDD1.n26 104.615
R1640 VDD1.n26 VDD1.n16 104.615
R1641 VDD1.n19 VDD1.n16 104.615
R1642 VDD1.n75 VDD1.n72 104.615
R1643 VDD1.n82 VDD1.n72 104.615
R1644 VDD1.n83 VDD1.n82 104.615
R1645 VDD1.n83 VDD1.n68 104.615
R1646 VDD1.n90 VDD1.n68 104.615
R1647 VDD1.n92 VDD1.n90 104.615
R1648 VDD1.n92 VDD1.n91 104.615
R1649 VDD1.n91 VDD1.n64 104.615
R1650 VDD1.n100 VDD1.n64 104.615
R1651 VDD1.n101 VDD1.n100 104.615
R1652 VDD1.n101 VDD1.n60 104.615
R1653 VDD1.n108 VDD1.n60 104.615
R1654 VDD1.n109 VDD1.n108 104.615
R1655 VDD1.n115 VDD1.n114 61.8452
R1656 VDD1.n117 VDD1.n116 61.7583
R1657 VDD1.n19 VDD1.t3 52.3082
R1658 VDD1.n75 VDD1.t5 52.3082
R1659 VDD1 VDD1.n56 48.7672
R1660 VDD1.n115 VDD1.n113 48.6537
R1661 VDD1.n117 VDD1.n115 35.613
R1662 VDD1.n42 VDD1.n41 13.1884
R1663 VDD1.n99 VDD1.n98 13.1884
R1664 VDD1.n45 VDD1.n6 12.8005
R1665 VDD1.n40 VDD1.n8 12.8005
R1666 VDD1.n97 VDD1.n65 12.8005
R1667 VDD1.n102 VDD1.n63 12.8005
R1668 VDD1.n46 VDD1.n4 12.0247
R1669 VDD1.n37 VDD1.n36 12.0247
R1670 VDD1.n94 VDD1.n93 12.0247
R1671 VDD1.n103 VDD1.n61 12.0247
R1672 VDD1.n50 VDD1.n49 11.249
R1673 VDD1.n33 VDD1.n10 11.249
R1674 VDD1.n89 VDD1.n67 11.249
R1675 VDD1.n107 VDD1.n106 11.249
R1676 VDD1.n53 VDD1.n2 10.4732
R1677 VDD1.n32 VDD1.n13 10.4732
R1678 VDD1.n88 VDD1.n69 10.4732
R1679 VDD1.n110 VDD1.n59 10.4732
R1680 VDD1.n20 VDD1.n18 10.2747
R1681 VDD1.n76 VDD1.n74 10.2747
R1682 VDD1.n54 VDD1.n0 9.69747
R1683 VDD1.n29 VDD1.n28 9.69747
R1684 VDD1.n85 VDD1.n84 9.69747
R1685 VDD1.n111 VDD1.n57 9.69747
R1686 VDD1.n56 VDD1.n55 9.45567
R1687 VDD1.n113 VDD1.n112 9.45567
R1688 VDD1.n22 VDD1.n21 9.3005
R1689 VDD1.n24 VDD1.n23 9.3005
R1690 VDD1.n15 VDD1.n14 9.3005
R1691 VDD1.n30 VDD1.n29 9.3005
R1692 VDD1.n32 VDD1.n31 9.3005
R1693 VDD1.n10 VDD1.n9 9.3005
R1694 VDD1.n38 VDD1.n37 9.3005
R1695 VDD1.n40 VDD1.n39 9.3005
R1696 VDD1.n55 VDD1.n54 9.3005
R1697 VDD1.n2 VDD1.n1 9.3005
R1698 VDD1.n49 VDD1.n48 9.3005
R1699 VDD1.n47 VDD1.n46 9.3005
R1700 VDD1.n6 VDD1.n5 9.3005
R1701 VDD1.n112 VDD1.n111 9.3005
R1702 VDD1.n59 VDD1.n58 9.3005
R1703 VDD1.n106 VDD1.n105 9.3005
R1704 VDD1.n104 VDD1.n103 9.3005
R1705 VDD1.n63 VDD1.n62 9.3005
R1706 VDD1.n78 VDD1.n77 9.3005
R1707 VDD1.n80 VDD1.n79 9.3005
R1708 VDD1.n71 VDD1.n70 9.3005
R1709 VDD1.n86 VDD1.n85 9.3005
R1710 VDD1.n88 VDD1.n87 9.3005
R1711 VDD1.n67 VDD1.n66 9.3005
R1712 VDD1.n95 VDD1.n94 9.3005
R1713 VDD1.n97 VDD1.n96 9.3005
R1714 VDD1.n25 VDD1.n15 8.92171
R1715 VDD1.n81 VDD1.n71 8.92171
R1716 VDD1.n24 VDD1.n17 8.14595
R1717 VDD1.n80 VDD1.n73 8.14595
R1718 VDD1.n21 VDD1.n20 7.3702
R1719 VDD1.n77 VDD1.n76 7.3702
R1720 VDD1.n21 VDD1.n17 5.81868
R1721 VDD1.n77 VDD1.n73 5.81868
R1722 VDD1.n25 VDD1.n24 5.04292
R1723 VDD1.n81 VDD1.n80 5.04292
R1724 VDD1.n56 VDD1.n0 4.26717
R1725 VDD1.n28 VDD1.n15 4.26717
R1726 VDD1.n84 VDD1.n71 4.26717
R1727 VDD1.n113 VDD1.n57 4.26717
R1728 VDD1.n54 VDD1.n53 3.49141
R1729 VDD1.n29 VDD1.n13 3.49141
R1730 VDD1.n85 VDD1.n69 3.49141
R1731 VDD1.n111 VDD1.n110 3.49141
R1732 VDD1.n22 VDD1.n18 2.84303
R1733 VDD1.n78 VDD1.n74 2.84303
R1734 VDD1.n50 VDD1.n2 2.71565
R1735 VDD1.n33 VDD1.n32 2.71565
R1736 VDD1.n89 VDD1.n88 2.71565
R1737 VDD1.n107 VDD1.n59 2.71565
R1738 VDD1.n49 VDD1.n4 1.93989
R1739 VDD1.n36 VDD1.n10 1.93989
R1740 VDD1.n93 VDD1.n67 1.93989
R1741 VDD1.n106 VDD1.n61 1.93989
R1742 VDD1.n116 VDD1.t2 1.85965
R1743 VDD1.n116 VDD1.t0 1.85965
R1744 VDD1.n114 VDD1.t4 1.85965
R1745 VDD1.n114 VDD1.t1 1.85965
R1746 VDD1.n46 VDD1.n45 1.16414
R1747 VDD1.n37 VDD1.n8 1.16414
R1748 VDD1.n94 VDD1.n65 1.16414
R1749 VDD1.n103 VDD1.n102 1.16414
R1750 VDD1.n42 VDD1.n6 0.388379
R1751 VDD1.n41 VDD1.n40 0.388379
R1752 VDD1.n98 VDD1.n97 0.388379
R1753 VDD1.n99 VDD1.n63 0.388379
R1754 VDD1.n55 VDD1.n1 0.155672
R1755 VDD1.n48 VDD1.n1 0.155672
R1756 VDD1.n48 VDD1.n47 0.155672
R1757 VDD1.n47 VDD1.n5 0.155672
R1758 VDD1.n39 VDD1.n5 0.155672
R1759 VDD1.n39 VDD1.n38 0.155672
R1760 VDD1.n38 VDD1.n9 0.155672
R1761 VDD1.n31 VDD1.n9 0.155672
R1762 VDD1.n31 VDD1.n30 0.155672
R1763 VDD1.n30 VDD1.n14 0.155672
R1764 VDD1.n23 VDD1.n14 0.155672
R1765 VDD1.n23 VDD1.n22 0.155672
R1766 VDD1.n79 VDD1.n78 0.155672
R1767 VDD1.n79 VDD1.n70 0.155672
R1768 VDD1.n86 VDD1.n70 0.155672
R1769 VDD1.n87 VDD1.n86 0.155672
R1770 VDD1.n87 VDD1.n66 0.155672
R1771 VDD1.n95 VDD1.n66 0.155672
R1772 VDD1.n96 VDD1.n95 0.155672
R1773 VDD1.n96 VDD1.n62 0.155672
R1774 VDD1.n104 VDD1.n62 0.155672
R1775 VDD1.n105 VDD1.n104 0.155672
R1776 VDD1.n105 VDD1.n58 0.155672
R1777 VDD1.n112 VDD1.n58 0.155672
R1778 VDD1 VDD1.n117 0.0845517
C0 VN VTAIL 2.18301f
C1 VN VDD1 0.147689f
C2 VTAIL VDD2 12.1141f
C3 VDD2 VDD1 0.580626f
C4 VN VP 4.47404f
C5 VTAIL VDD1 12.0832f
C6 VP VDD2 0.266282f
C7 VTAIL VP 2.19769f
C8 VP VDD1 2.69103f
C9 VN VDD2 2.57694f
C10 VDD2 B 3.983615f
C11 VDD1 B 3.939879f
C12 VTAIL B 5.557331f
C13 VN B 6.72213f
C14 VP B 4.556145f
C15 VDD1.n0 B 0.036173f
C16 VDD1.n1 B 0.02717f
C17 VDD1.n2 B 0.0146f
C18 VDD1.n3 B 0.034509f
C19 VDD1.n4 B 0.015459f
C20 VDD1.n5 B 0.02717f
C21 VDD1.n6 B 0.0146f
C22 VDD1.n7 B 0.034509f
C23 VDD1.n8 B 0.015459f
C24 VDD1.n9 B 0.02717f
C25 VDD1.n10 B 0.0146f
C26 VDD1.n11 B 0.034509f
C27 VDD1.n12 B 0.034509f
C28 VDD1.n13 B 0.015459f
C29 VDD1.n14 B 0.02717f
C30 VDD1.n15 B 0.0146f
C31 VDD1.n16 B 0.034509f
C32 VDD1.n17 B 0.015459f
C33 VDD1.n18 B 0.181812f
C34 VDD1.t3 B 0.058087f
C35 VDD1.n19 B 0.025882f
C36 VDD1.n20 B 0.024395f
C37 VDD1.n21 B 0.0146f
C38 VDD1.n22 B 1.20753f
C39 VDD1.n23 B 0.02717f
C40 VDD1.n24 B 0.0146f
C41 VDD1.n25 B 0.015459f
C42 VDD1.n26 B 0.034509f
C43 VDD1.n27 B 0.034509f
C44 VDD1.n28 B 0.015459f
C45 VDD1.n29 B 0.0146f
C46 VDD1.n30 B 0.02717f
C47 VDD1.n31 B 0.02717f
C48 VDD1.n32 B 0.0146f
C49 VDD1.n33 B 0.015459f
C50 VDD1.n34 B 0.034509f
C51 VDD1.n35 B 0.034509f
C52 VDD1.n36 B 0.015459f
C53 VDD1.n37 B 0.0146f
C54 VDD1.n38 B 0.02717f
C55 VDD1.n39 B 0.02717f
C56 VDD1.n40 B 0.0146f
C57 VDD1.n41 B 0.015029f
C58 VDD1.n42 B 0.015029f
C59 VDD1.n43 B 0.034509f
C60 VDD1.n44 B 0.034509f
C61 VDD1.n45 B 0.015459f
C62 VDD1.n46 B 0.0146f
C63 VDD1.n47 B 0.02717f
C64 VDD1.n48 B 0.02717f
C65 VDD1.n49 B 0.0146f
C66 VDD1.n50 B 0.015459f
C67 VDD1.n51 B 0.034509f
C68 VDD1.n52 B 0.07114f
C69 VDD1.n53 B 0.015459f
C70 VDD1.n54 B 0.0146f
C71 VDD1.n55 B 0.061688f
C72 VDD1.n56 B 0.05911f
C73 VDD1.n57 B 0.036173f
C74 VDD1.n58 B 0.02717f
C75 VDD1.n59 B 0.0146f
C76 VDD1.n60 B 0.034509f
C77 VDD1.n61 B 0.015459f
C78 VDD1.n62 B 0.02717f
C79 VDD1.n63 B 0.0146f
C80 VDD1.n64 B 0.034509f
C81 VDD1.n65 B 0.015459f
C82 VDD1.n66 B 0.02717f
C83 VDD1.n67 B 0.0146f
C84 VDD1.n68 B 0.034509f
C85 VDD1.n69 B 0.015459f
C86 VDD1.n70 B 0.02717f
C87 VDD1.n71 B 0.0146f
C88 VDD1.n72 B 0.034509f
C89 VDD1.n73 B 0.015459f
C90 VDD1.n74 B 0.181812f
C91 VDD1.t5 B 0.058087f
C92 VDD1.n75 B 0.025882f
C93 VDD1.n76 B 0.024395f
C94 VDD1.n77 B 0.0146f
C95 VDD1.n78 B 1.20753f
C96 VDD1.n79 B 0.02717f
C97 VDD1.n80 B 0.0146f
C98 VDD1.n81 B 0.015459f
C99 VDD1.n82 B 0.034509f
C100 VDD1.n83 B 0.034509f
C101 VDD1.n84 B 0.015459f
C102 VDD1.n85 B 0.0146f
C103 VDD1.n86 B 0.02717f
C104 VDD1.n87 B 0.02717f
C105 VDD1.n88 B 0.0146f
C106 VDD1.n89 B 0.015459f
C107 VDD1.n90 B 0.034509f
C108 VDD1.n91 B 0.034509f
C109 VDD1.n92 B 0.034509f
C110 VDD1.n93 B 0.015459f
C111 VDD1.n94 B 0.0146f
C112 VDD1.n95 B 0.02717f
C113 VDD1.n96 B 0.02717f
C114 VDD1.n97 B 0.0146f
C115 VDD1.n98 B 0.015029f
C116 VDD1.n99 B 0.015029f
C117 VDD1.n100 B 0.034509f
C118 VDD1.n101 B 0.034509f
C119 VDD1.n102 B 0.015459f
C120 VDD1.n103 B 0.0146f
C121 VDD1.n104 B 0.02717f
C122 VDD1.n105 B 0.02717f
C123 VDD1.n106 B 0.0146f
C124 VDD1.n107 B 0.015459f
C125 VDD1.n108 B 0.034509f
C126 VDD1.n109 B 0.07114f
C127 VDD1.n110 B 0.015459f
C128 VDD1.n111 B 0.0146f
C129 VDD1.n112 B 0.061688f
C130 VDD1.n113 B 0.058829f
C131 VDD1.t4 B 0.228661f
C132 VDD1.t1 B 0.228661f
C133 VDD1.n114 B 2.02183f
C134 VDD1.n115 B 1.82214f
C135 VDD1.t2 B 0.228661f
C136 VDD1.t0 B 0.228661f
C137 VDD1.n116 B 2.02141f
C138 VDD1.n117 B 2.21985f
C139 VP.n0 B 0.05768f
C140 VP.t1 B 0.57362f
C141 VP.t0 B 0.579616f
C142 VP.t2 B 0.587622f
C143 VP.n1 B 0.24133f
C144 VP.t3 B 0.57362f
C145 VP.n2 B 0.249578f
C146 VP.t5 B 0.579616f
C147 VP.n3 B 0.248917f
C148 VP.n4 B 2.19255f
C149 VP.n5 B 2.12581f
C150 VP.n6 B 0.248917f
C151 VP.n7 B 0.249578f
C152 VP.t4 B 0.579616f
C153 VP.n8 B 0.248917f
C154 VP.n9 B 0.0447f
C155 VDD2.n0 B 0.036174f
C156 VDD2.n1 B 0.027171f
C157 VDD2.n2 B 0.0146f
C158 VDD2.n3 B 0.03451f
C159 VDD2.n4 B 0.015459f
C160 VDD2.n5 B 0.027171f
C161 VDD2.n6 B 0.0146f
C162 VDD2.n7 B 0.03451f
C163 VDD2.n8 B 0.015459f
C164 VDD2.n9 B 0.027171f
C165 VDD2.n10 B 0.0146f
C166 VDD2.n11 B 0.03451f
C167 VDD2.n12 B 0.015459f
C168 VDD2.n13 B 0.027171f
C169 VDD2.n14 B 0.0146f
C170 VDD2.n15 B 0.03451f
C171 VDD2.n16 B 0.015459f
C172 VDD2.n17 B 0.181816f
C173 VDD2.t5 B 0.058088f
C174 VDD2.n18 B 0.025882f
C175 VDD2.n19 B 0.024396f
C176 VDD2.n20 B 0.0146f
C177 VDD2.n21 B 1.20756f
C178 VDD2.n22 B 0.027171f
C179 VDD2.n23 B 0.0146f
C180 VDD2.n24 B 0.015459f
C181 VDD2.n25 B 0.03451f
C182 VDD2.n26 B 0.03451f
C183 VDD2.n27 B 0.015459f
C184 VDD2.n28 B 0.0146f
C185 VDD2.n29 B 0.027171f
C186 VDD2.n30 B 0.027171f
C187 VDD2.n31 B 0.0146f
C188 VDD2.n32 B 0.015459f
C189 VDD2.n33 B 0.03451f
C190 VDD2.n34 B 0.03451f
C191 VDD2.n35 B 0.03451f
C192 VDD2.n36 B 0.015459f
C193 VDD2.n37 B 0.0146f
C194 VDD2.n38 B 0.027171f
C195 VDD2.n39 B 0.027171f
C196 VDD2.n40 B 0.0146f
C197 VDD2.n41 B 0.01503f
C198 VDD2.n42 B 0.01503f
C199 VDD2.n43 B 0.03451f
C200 VDD2.n44 B 0.03451f
C201 VDD2.n45 B 0.015459f
C202 VDD2.n46 B 0.0146f
C203 VDD2.n47 B 0.027171f
C204 VDD2.n48 B 0.027171f
C205 VDD2.n49 B 0.0146f
C206 VDD2.n50 B 0.015459f
C207 VDD2.n51 B 0.03451f
C208 VDD2.n52 B 0.071142f
C209 VDD2.n53 B 0.015459f
C210 VDD2.n54 B 0.0146f
C211 VDD2.n55 B 0.06169f
C212 VDD2.n56 B 0.058831f
C213 VDD2.t3 B 0.228666f
C214 VDD2.t0 B 0.228666f
C215 VDD2.n57 B 2.02188f
C216 VDD2.n58 B 1.74788f
C217 VDD2.n59 B 0.036174f
C218 VDD2.n60 B 0.027171f
C219 VDD2.n61 B 0.0146f
C220 VDD2.n62 B 0.03451f
C221 VDD2.n63 B 0.015459f
C222 VDD2.n64 B 0.027171f
C223 VDD2.n65 B 0.0146f
C224 VDD2.n66 B 0.03451f
C225 VDD2.n67 B 0.015459f
C226 VDD2.n68 B 0.027171f
C227 VDD2.n69 B 0.0146f
C228 VDD2.n70 B 0.03451f
C229 VDD2.n71 B 0.03451f
C230 VDD2.n72 B 0.015459f
C231 VDD2.n73 B 0.027171f
C232 VDD2.n74 B 0.0146f
C233 VDD2.n75 B 0.03451f
C234 VDD2.n76 B 0.015459f
C235 VDD2.n77 B 0.181816f
C236 VDD2.t4 B 0.058088f
C237 VDD2.n78 B 0.025882f
C238 VDD2.n79 B 0.024396f
C239 VDD2.n80 B 0.0146f
C240 VDD2.n81 B 1.20756f
C241 VDD2.n82 B 0.027171f
C242 VDD2.n83 B 0.0146f
C243 VDD2.n84 B 0.015459f
C244 VDD2.n85 B 0.03451f
C245 VDD2.n86 B 0.03451f
C246 VDD2.n87 B 0.015459f
C247 VDD2.n88 B 0.0146f
C248 VDD2.n89 B 0.027171f
C249 VDD2.n90 B 0.027171f
C250 VDD2.n91 B 0.0146f
C251 VDD2.n92 B 0.015459f
C252 VDD2.n93 B 0.03451f
C253 VDD2.n94 B 0.03451f
C254 VDD2.n95 B 0.015459f
C255 VDD2.n96 B 0.0146f
C256 VDD2.n97 B 0.027171f
C257 VDD2.n98 B 0.027171f
C258 VDD2.n99 B 0.0146f
C259 VDD2.n100 B 0.01503f
C260 VDD2.n101 B 0.01503f
C261 VDD2.n102 B 0.03451f
C262 VDD2.n103 B 0.03451f
C263 VDD2.n104 B 0.015459f
C264 VDD2.n105 B 0.0146f
C265 VDD2.n106 B 0.027171f
C266 VDD2.n107 B 0.027171f
C267 VDD2.n108 B 0.0146f
C268 VDD2.n109 B 0.015459f
C269 VDD2.n110 B 0.03451f
C270 VDD2.n111 B 0.071142f
C271 VDD2.n112 B 0.015459f
C272 VDD2.n113 B 0.0146f
C273 VDD2.n114 B 0.06169f
C274 VDD2.n115 B 0.058175f
C275 VDD2.n116 B 1.9964f
C276 VDD2.t1 B 0.228666f
C277 VDD2.t2 B 0.228666f
C278 VDD2.n117 B 2.02185f
C279 VTAIL.t7 B 0.236601f
C280 VTAIL.t8 B 0.236601f
C281 VTAIL.n0 B 2.00803f
C282 VTAIL.n1 B 0.363075f
C283 VTAIL.n2 B 0.037429f
C284 VTAIL.n3 B 0.028113f
C285 VTAIL.n4 B 0.015107f
C286 VTAIL.n5 B 0.035707f
C287 VTAIL.n6 B 0.015995f
C288 VTAIL.n7 B 0.028113f
C289 VTAIL.n8 B 0.015107f
C290 VTAIL.n9 B 0.035707f
C291 VTAIL.n10 B 0.015995f
C292 VTAIL.n11 B 0.028113f
C293 VTAIL.n12 B 0.015107f
C294 VTAIL.n13 B 0.035707f
C295 VTAIL.n14 B 0.015995f
C296 VTAIL.n15 B 0.028113f
C297 VTAIL.n16 B 0.015107f
C298 VTAIL.n17 B 0.035707f
C299 VTAIL.n18 B 0.015995f
C300 VTAIL.n19 B 0.188124f
C301 VTAIL.t3 B 0.060103f
C302 VTAIL.n20 B 0.02678f
C303 VTAIL.n21 B 0.025242f
C304 VTAIL.n22 B 0.015107f
C305 VTAIL.n23 B 1.24946f
C306 VTAIL.n24 B 0.028113f
C307 VTAIL.n25 B 0.015107f
C308 VTAIL.n26 B 0.015995f
C309 VTAIL.n27 B 0.035707f
C310 VTAIL.n28 B 0.035707f
C311 VTAIL.n29 B 0.015995f
C312 VTAIL.n30 B 0.015107f
C313 VTAIL.n31 B 0.028113f
C314 VTAIL.n32 B 0.028113f
C315 VTAIL.n33 B 0.015107f
C316 VTAIL.n34 B 0.015995f
C317 VTAIL.n35 B 0.035707f
C318 VTAIL.n36 B 0.035707f
C319 VTAIL.n37 B 0.035707f
C320 VTAIL.n38 B 0.015995f
C321 VTAIL.n39 B 0.015107f
C322 VTAIL.n40 B 0.028113f
C323 VTAIL.n41 B 0.028113f
C324 VTAIL.n42 B 0.015107f
C325 VTAIL.n43 B 0.015551f
C326 VTAIL.n44 B 0.015551f
C327 VTAIL.n45 B 0.035707f
C328 VTAIL.n46 B 0.035707f
C329 VTAIL.n47 B 0.015995f
C330 VTAIL.n48 B 0.015107f
C331 VTAIL.n49 B 0.028113f
C332 VTAIL.n50 B 0.028113f
C333 VTAIL.n51 B 0.015107f
C334 VTAIL.n52 B 0.015995f
C335 VTAIL.n53 B 0.035707f
C336 VTAIL.n54 B 0.07361f
C337 VTAIL.n55 B 0.015995f
C338 VTAIL.n56 B 0.015107f
C339 VTAIL.n57 B 0.063831f
C340 VTAIL.n58 B 0.040773f
C341 VTAIL.n59 B 0.143233f
C342 VTAIL.t0 B 0.236601f
C343 VTAIL.t5 B 0.236601f
C344 VTAIL.n60 B 2.00803f
C345 VTAIL.n61 B 1.64478f
C346 VTAIL.t10 B 0.236601f
C347 VTAIL.t9 B 0.236601f
C348 VTAIL.n62 B 2.00804f
C349 VTAIL.n63 B 1.64477f
C350 VTAIL.n64 B 0.037429f
C351 VTAIL.n65 B 0.028113f
C352 VTAIL.n66 B 0.015107f
C353 VTAIL.n67 B 0.035707f
C354 VTAIL.n68 B 0.015995f
C355 VTAIL.n69 B 0.028113f
C356 VTAIL.n70 B 0.015107f
C357 VTAIL.n71 B 0.035707f
C358 VTAIL.n72 B 0.015995f
C359 VTAIL.n73 B 0.028113f
C360 VTAIL.n74 B 0.015107f
C361 VTAIL.n75 B 0.035707f
C362 VTAIL.n76 B 0.035707f
C363 VTAIL.n77 B 0.015995f
C364 VTAIL.n78 B 0.028113f
C365 VTAIL.n79 B 0.015107f
C366 VTAIL.n80 B 0.035707f
C367 VTAIL.n81 B 0.015995f
C368 VTAIL.n82 B 0.188124f
C369 VTAIL.t11 B 0.060103f
C370 VTAIL.n83 B 0.02678f
C371 VTAIL.n84 B 0.025242f
C372 VTAIL.n85 B 0.015107f
C373 VTAIL.n86 B 1.24946f
C374 VTAIL.n87 B 0.028113f
C375 VTAIL.n88 B 0.015107f
C376 VTAIL.n89 B 0.015995f
C377 VTAIL.n90 B 0.035707f
C378 VTAIL.n91 B 0.035707f
C379 VTAIL.n92 B 0.015995f
C380 VTAIL.n93 B 0.015107f
C381 VTAIL.n94 B 0.028113f
C382 VTAIL.n95 B 0.028113f
C383 VTAIL.n96 B 0.015107f
C384 VTAIL.n97 B 0.015995f
C385 VTAIL.n98 B 0.035707f
C386 VTAIL.n99 B 0.035707f
C387 VTAIL.n100 B 0.015995f
C388 VTAIL.n101 B 0.015107f
C389 VTAIL.n102 B 0.028113f
C390 VTAIL.n103 B 0.028113f
C391 VTAIL.n104 B 0.015107f
C392 VTAIL.n105 B 0.015551f
C393 VTAIL.n106 B 0.015551f
C394 VTAIL.n107 B 0.035707f
C395 VTAIL.n108 B 0.035707f
C396 VTAIL.n109 B 0.015995f
C397 VTAIL.n110 B 0.015107f
C398 VTAIL.n111 B 0.028113f
C399 VTAIL.n112 B 0.028113f
C400 VTAIL.n113 B 0.015107f
C401 VTAIL.n114 B 0.015995f
C402 VTAIL.n115 B 0.035707f
C403 VTAIL.n116 B 0.07361f
C404 VTAIL.n117 B 0.015995f
C405 VTAIL.n118 B 0.015107f
C406 VTAIL.n119 B 0.063831f
C407 VTAIL.n120 B 0.040773f
C408 VTAIL.n121 B 0.143233f
C409 VTAIL.t4 B 0.236601f
C410 VTAIL.t1 B 0.236601f
C411 VTAIL.n122 B 2.00804f
C412 VTAIL.n123 B 0.396448f
C413 VTAIL.n124 B 0.037429f
C414 VTAIL.n125 B 0.028113f
C415 VTAIL.n126 B 0.015107f
C416 VTAIL.n127 B 0.035707f
C417 VTAIL.n128 B 0.015995f
C418 VTAIL.n129 B 0.028113f
C419 VTAIL.n130 B 0.015107f
C420 VTAIL.n131 B 0.035707f
C421 VTAIL.n132 B 0.015995f
C422 VTAIL.n133 B 0.028113f
C423 VTAIL.n134 B 0.015107f
C424 VTAIL.n135 B 0.035707f
C425 VTAIL.n136 B 0.035707f
C426 VTAIL.n137 B 0.015995f
C427 VTAIL.n138 B 0.028113f
C428 VTAIL.n139 B 0.015107f
C429 VTAIL.n140 B 0.035707f
C430 VTAIL.n141 B 0.015995f
C431 VTAIL.n142 B 0.188124f
C432 VTAIL.t2 B 0.060103f
C433 VTAIL.n143 B 0.02678f
C434 VTAIL.n144 B 0.025242f
C435 VTAIL.n145 B 0.015107f
C436 VTAIL.n146 B 1.24946f
C437 VTAIL.n147 B 0.028113f
C438 VTAIL.n148 B 0.015107f
C439 VTAIL.n149 B 0.015995f
C440 VTAIL.n150 B 0.035707f
C441 VTAIL.n151 B 0.035707f
C442 VTAIL.n152 B 0.015995f
C443 VTAIL.n153 B 0.015107f
C444 VTAIL.n154 B 0.028113f
C445 VTAIL.n155 B 0.028113f
C446 VTAIL.n156 B 0.015107f
C447 VTAIL.n157 B 0.015995f
C448 VTAIL.n158 B 0.035707f
C449 VTAIL.n159 B 0.035707f
C450 VTAIL.n160 B 0.015995f
C451 VTAIL.n161 B 0.015107f
C452 VTAIL.n162 B 0.028113f
C453 VTAIL.n163 B 0.028113f
C454 VTAIL.n164 B 0.015107f
C455 VTAIL.n165 B 0.015551f
C456 VTAIL.n166 B 0.015551f
C457 VTAIL.n167 B 0.035707f
C458 VTAIL.n168 B 0.035707f
C459 VTAIL.n169 B 0.015995f
C460 VTAIL.n170 B 0.015107f
C461 VTAIL.n171 B 0.028113f
C462 VTAIL.n172 B 0.028113f
C463 VTAIL.n173 B 0.015107f
C464 VTAIL.n174 B 0.015995f
C465 VTAIL.n175 B 0.035707f
C466 VTAIL.n176 B 0.07361f
C467 VTAIL.n177 B 0.015995f
C468 VTAIL.n178 B 0.015107f
C469 VTAIL.n179 B 0.063831f
C470 VTAIL.n180 B 0.040773f
C471 VTAIL.n181 B 1.34002f
C472 VTAIL.n182 B 0.037429f
C473 VTAIL.n183 B 0.028113f
C474 VTAIL.n184 B 0.015107f
C475 VTAIL.n185 B 0.035707f
C476 VTAIL.n186 B 0.015995f
C477 VTAIL.n187 B 0.028113f
C478 VTAIL.n188 B 0.015107f
C479 VTAIL.n189 B 0.035707f
C480 VTAIL.n190 B 0.015995f
C481 VTAIL.n191 B 0.028113f
C482 VTAIL.n192 B 0.015107f
C483 VTAIL.n193 B 0.035707f
C484 VTAIL.n194 B 0.015995f
C485 VTAIL.n195 B 0.028113f
C486 VTAIL.n196 B 0.015107f
C487 VTAIL.n197 B 0.035707f
C488 VTAIL.n198 B 0.015995f
C489 VTAIL.n199 B 0.188124f
C490 VTAIL.t6 B 0.060103f
C491 VTAIL.n200 B 0.02678f
C492 VTAIL.n201 B 0.025242f
C493 VTAIL.n202 B 0.015107f
C494 VTAIL.n203 B 1.24946f
C495 VTAIL.n204 B 0.028113f
C496 VTAIL.n205 B 0.015107f
C497 VTAIL.n206 B 0.015995f
C498 VTAIL.n207 B 0.035707f
C499 VTAIL.n208 B 0.035707f
C500 VTAIL.n209 B 0.015995f
C501 VTAIL.n210 B 0.015107f
C502 VTAIL.n211 B 0.028113f
C503 VTAIL.n212 B 0.028113f
C504 VTAIL.n213 B 0.015107f
C505 VTAIL.n214 B 0.015995f
C506 VTAIL.n215 B 0.035707f
C507 VTAIL.n216 B 0.035707f
C508 VTAIL.n217 B 0.035707f
C509 VTAIL.n218 B 0.015995f
C510 VTAIL.n219 B 0.015107f
C511 VTAIL.n220 B 0.028113f
C512 VTAIL.n221 B 0.028113f
C513 VTAIL.n222 B 0.015107f
C514 VTAIL.n223 B 0.015551f
C515 VTAIL.n224 B 0.015551f
C516 VTAIL.n225 B 0.035707f
C517 VTAIL.n226 B 0.035707f
C518 VTAIL.n227 B 0.015995f
C519 VTAIL.n228 B 0.015107f
C520 VTAIL.n229 B 0.028113f
C521 VTAIL.n230 B 0.028113f
C522 VTAIL.n231 B 0.015107f
C523 VTAIL.n232 B 0.015995f
C524 VTAIL.n233 B 0.035707f
C525 VTAIL.n234 B 0.07361f
C526 VTAIL.n235 B 0.015995f
C527 VTAIL.n236 B 0.015107f
C528 VTAIL.n237 B 0.063831f
C529 VTAIL.n238 B 0.040773f
C530 VTAIL.n239 B 1.32186f
C531 VN.t0 B 0.576399f
C532 VN.n0 B 0.236721f
C533 VN.t2 B 0.562664f
C534 VN.n1 B 0.244811f
C535 VN.t5 B 0.568545f
C536 VN.n2 B 0.244163f
C537 VN.n3 B 0.161824f
C538 VN.t3 B 0.576399f
C539 VN.n4 B 0.236721f
C540 VN.t1 B 0.568545f
C541 VN.t4 B 0.562664f
C542 VN.n5 B 0.244811f
C543 VN.n6 B 0.244163f
C544 VN.n7 B 2.18801f
.ends

