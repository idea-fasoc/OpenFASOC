* NGSPICE file created from diff_pair_sample_0355.ext - technology: sky130A

.subckt diff_pair_sample_0355 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=1.2636 ps=7.26 w=3.24 l=0.88
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=1.2636 ps=7.26 w=3.24 l=0.88
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=1.2636 ps=7.26 w=3.24 l=0.88
X3 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=1.2636 ps=7.26 w=3.24 l=0.88
X4 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=0 ps=0 w=3.24 l=0.88
X5 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=0 ps=0 w=3.24 l=0.88
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=0 ps=0 w=3.24 l=0.88
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2636 pd=7.26 as=0 ps=0 w=3.24 l=0.88
R0 VN VN.t0 328.526
R1 VN VN.t1 294.724
R2 VTAIL.n58 VTAIL.n48 289.615
R3 VTAIL.n10 VTAIL.n0 289.615
R4 VTAIL.n42 VTAIL.n32 289.615
R5 VTAIL.n26 VTAIL.n16 289.615
R6 VTAIL.n52 VTAIL.n51 185
R7 VTAIL.n57 VTAIL.n56 185
R8 VTAIL.n59 VTAIL.n58 185
R9 VTAIL.n4 VTAIL.n3 185
R10 VTAIL.n9 VTAIL.n8 185
R11 VTAIL.n11 VTAIL.n10 185
R12 VTAIL.n43 VTAIL.n42 185
R13 VTAIL.n41 VTAIL.n40 185
R14 VTAIL.n36 VTAIL.n35 185
R15 VTAIL.n27 VTAIL.n26 185
R16 VTAIL.n25 VTAIL.n24 185
R17 VTAIL.n20 VTAIL.n19 185
R18 VTAIL.n53 VTAIL.t0 148.606
R19 VTAIL.n5 VTAIL.t2 148.606
R20 VTAIL.n37 VTAIL.t3 148.606
R21 VTAIL.n21 VTAIL.t1 148.606
R22 VTAIL.n57 VTAIL.n51 104.615
R23 VTAIL.n58 VTAIL.n57 104.615
R24 VTAIL.n9 VTAIL.n3 104.615
R25 VTAIL.n10 VTAIL.n9 104.615
R26 VTAIL.n42 VTAIL.n41 104.615
R27 VTAIL.n41 VTAIL.n35 104.615
R28 VTAIL.n26 VTAIL.n25 104.615
R29 VTAIL.n25 VTAIL.n19 104.615
R30 VTAIL.t0 VTAIL.n51 52.3082
R31 VTAIL.t2 VTAIL.n3 52.3082
R32 VTAIL.t3 VTAIL.n35 52.3082
R33 VTAIL.t1 VTAIL.n19 52.3082
R34 VTAIL.n63 VTAIL.n62 34.5126
R35 VTAIL.n15 VTAIL.n14 34.5126
R36 VTAIL.n47 VTAIL.n46 34.5126
R37 VTAIL.n31 VTAIL.n30 34.5126
R38 VTAIL.n31 VTAIL.n15 17.2634
R39 VTAIL.n63 VTAIL.n47 16.2203
R40 VTAIL.n53 VTAIL.n52 15.5966
R41 VTAIL.n5 VTAIL.n4 15.5966
R42 VTAIL.n37 VTAIL.n36 15.5966
R43 VTAIL.n21 VTAIL.n20 15.5966
R44 VTAIL.n56 VTAIL.n55 12.8005
R45 VTAIL.n8 VTAIL.n7 12.8005
R46 VTAIL.n40 VTAIL.n39 12.8005
R47 VTAIL.n24 VTAIL.n23 12.8005
R48 VTAIL.n59 VTAIL.n50 12.0247
R49 VTAIL.n11 VTAIL.n2 12.0247
R50 VTAIL.n43 VTAIL.n34 12.0247
R51 VTAIL.n27 VTAIL.n18 12.0247
R52 VTAIL.n60 VTAIL.n48 11.249
R53 VTAIL.n12 VTAIL.n0 11.249
R54 VTAIL.n44 VTAIL.n32 11.249
R55 VTAIL.n28 VTAIL.n16 11.249
R56 VTAIL.n62 VTAIL.n61 9.45567
R57 VTAIL.n14 VTAIL.n13 9.45567
R58 VTAIL.n46 VTAIL.n45 9.45567
R59 VTAIL.n30 VTAIL.n29 9.45567
R60 VTAIL.n61 VTAIL.n60 9.3005
R61 VTAIL.n50 VTAIL.n49 9.3005
R62 VTAIL.n55 VTAIL.n54 9.3005
R63 VTAIL.n13 VTAIL.n12 9.3005
R64 VTAIL.n2 VTAIL.n1 9.3005
R65 VTAIL.n7 VTAIL.n6 9.3005
R66 VTAIL.n45 VTAIL.n44 9.3005
R67 VTAIL.n34 VTAIL.n33 9.3005
R68 VTAIL.n39 VTAIL.n38 9.3005
R69 VTAIL.n29 VTAIL.n28 9.3005
R70 VTAIL.n18 VTAIL.n17 9.3005
R71 VTAIL.n23 VTAIL.n22 9.3005
R72 VTAIL.n54 VTAIL.n53 4.46457
R73 VTAIL.n6 VTAIL.n5 4.46457
R74 VTAIL.n38 VTAIL.n37 4.46457
R75 VTAIL.n22 VTAIL.n21 4.46457
R76 VTAIL.n62 VTAIL.n48 2.71565
R77 VTAIL.n14 VTAIL.n0 2.71565
R78 VTAIL.n46 VTAIL.n32 2.71565
R79 VTAIL.n30 VTAIL.n16 2.71565
R80 VTAIL.n60 VTAIL.n59 1.93989
R81 VTAIL.n12 VTAIL.n11 1.93989
R82 VTAIL.n44 VTAIL.n43 1.93989
R83 VTAIL.n28 VTAIL.n27 1.93989
R84 VTAIL.n56 VTAIL.n50 1.16414
R85 VTAIL.n8 VTAIL.n2 1.16414
R86 VTAIL.n40 VTAIL.n34 1.16414
R87 VTAIL.n24 VTAIL.n18 1.16414
R88 VTAIL.n47 VTAIL.n31 0.991879
R89 VTAIL VTAIL.n15 0.789293
R90 VTAIL.n55 VTAIL.n52 0.388379
R91 VTAIL.n7 VTAIL.n4 0.388379
R92 VTAIL.n39 VTAIL.n36 0.388379
R93 VTAIL.n23 VTAIL.n20 0.388379
R94 VTAIL VTAIL.n63 0.203086
R95 VTAIL.n54 VTAIL.n49 0.155672
R96 VTAIL.n61 VTAIL.n49 0.155672
R97 VTAIL.n6 VTAIL.n1 0.155672
R98 VTAIL.n13 VTAIL.n1 0.155672
R99 VTAIL.n45 VTAIL.n33 0.155672
R100 VTAIL.n38 VTAIL.n33 0.155672
R101 VTAIL.n29 VTAIL.n17 0.155672
R102 VTAIL.n22 VTAIL.n17 0.155672
R103 VDD2.n25 VDD2.n15 289.615
R104 VDD2.n10 VDD2.n0 289.615
R105 VDD2.n26 VDD2.n25 185
R106 VDD2.n24 VDD2.n23 185
R107 VDD2.n19 VDD2.n18 185
R108 VDD2.n4 VDD2.n3 185
R109 VDD2.n9 VDD2.n8 185
R110 VDD2.n11 VDD2.n10 185
R111 VDD2.n20 VDD2.t1 148.606
R112 VDD2.n5 VDD2.t0 148.606
R113 VDD2.n25 VDD2.n24 104.615
R114 VDD2.n24 VDD2.n18 104.615
R115 VDD2.n9 VDD2.n3 104.615
R116 VDD2.n10 VDD2.n9 104.615
R117 VDD2.n30 VDD2.n14 79.7474
R118 VDD2.t1 VDD2.n18 52.3082
R119 VDD2.t0 VDD2.n3 52.3082
R120 VDD2.n30 VDD2.n29 51.1914
R121 VDD2.n20 VDD2.n19 15.5966
R122 VDD2.n5 VDD2.n4 15.5966
R123 VDD2.n23 VDD2.n22 12.8005
R124 VDD2.n8 VDD2.n7 12.8005
R125 VDD2.n26 VDD2.n17 12.0247
R126 VDD2.n11 VDD2.n2 12.0247
R127 VDD2.n27 VDD2.n15 11.249
R128 VDD2.n12 VDD2.n0 11.249
R129 VDD2.n29 VDD2.n28 9.45567
R130 VDD2.n14 VDD2.n13 9.45567
R131 VDD2.n28 VDD2.n27 9.3005
R132 VDD2.n17 VDD2.n16 9.3005
R133 VDD2.n22 VDD2.n21 9.3005
R134 VDD2.n13 VDD2.n12 9.3005
R135 VDD2.n2 VDD2.n1 9.3005
R136 VDD2.n7 VDD2.n6 9.3005
R137 VDD2.n21 VDD2.n20 4.46457
R138 VDD2.n6 VDD2.n5 4.46457
R139 VDD2.n29 VDD2.n15 2.71565
R140 VDD2.n14 VDD2.n0 2.71565
R141 VDD2.n27 VDD2.n26 1.93989
R142 VDD2.n12 VDD2.n11 1.93989
R143 VDD2.n23 VDD2.n17 1.16414
R144 VDD2.n8 VDD2.n2 1.16414
R145 VDD2.n22 VDD2.n19 0.388379
R146 VDD2.n7 VDD2.n4 0.388379
R147 VDD2 VDD2.n30 0.319466
R148 VDD2.n28 VDD2.n16 0.155672
R149 VDD2.n21 VDD2.n16 0.155672
R150 VDD2.n6 VDD2.n1 0.155672
R151 VDD2.n13 VDD2.n1 0.155672
R152 B.n336 B.n335 585
R153 B.n337 B.n336 585
R154 B.n134 B.n52 585
R155 B.n133 B.n132 585
R156 B.n131 B.n130 585
R157 B.n129 B.n128 585
R158 B.n127 B.n126 585
R159 B.n125 B.n124 585
R160 B.n123 B.n122 585
R161 B.n121 B.n120 585
R162 B.n119 B.n118 585
R163 B.n117 B.n116 585
R164 B.n115 B.n114 585
R165 B.n113 B.n112 585
R166 B.n111 B.n110 585
R167 B.n109 B.n108 585
R168 B.n107 B.n106 585
R169 B.n104 B.n103 585
R170 B.n102 B.n101 585
R171 B.n100 B.n99 585
R172 B.n98 B.n97 585
R173 B.n96 B.n95 585
R174 B.n94 B.n93 585
R175 B.n92 B.n91 585
R176 B.n90 B.n89 585
R177 B.n88 B.n87 585
R178 B.n86 B.n85 585
R179 B.n84 B.n83 585
R180 B.n82 B.n81 585
R181 B.n80 B.n79 585
R182 B.n78 B.n77 585
R183 B.n76 B.n75 585
R184 B.n74 B.n73 585
R185 B.n72 B.n71 585
R186 B.n70 B.n69 585
R187 B.n68 B.n67 585
R188 B.n66 B.n65 585
R189 B.n64 B.n63 585
R190 B.n62 B.n61 585
R191 B.n60 B.n59 585
R192 B.n32 B.n31 585
R193 B.n340 B.n339 585
R194 B.n334 B.n53 585
R195 B.n53 B.n29 585
R196 B.n333 B.n28 585
R197 B.n344 B.n28 585
R198 B.n332 B.n27 585
R199 B.n345 B.n27 585
R200 B.n331 B.n26 585
R201 B.n346 B.n26 585
R202 B.n330 B.n329 585
R203 B.n329 B.n25 585
R204 B.n328 B.n21 585
R205 B.n352 B.n21 585
R206 B.n327 B.n20 585
R207 B.n353 B.n20 585
R208 B.n326 B.n19 585
R209 B.n354 B.n19 585
R210 B.n325 B.n324 585
R211 B.n324 B.n15 585
R212 B.n323 B.n14 585
R213 B.n360 B.n14 585
R214 B.n322 B.n13 585
R215 B.n361 B.n13 585
R216 B.n321 B.n12 585
R217 B.n362 B.n12 585
R218 B.n320 B.n319 585
R219 B.n319 B.n8 585
R220 B.n318 B.n7 585
R221 B.n368 B.n7 585
R222 B.n317 B.n6 585
R223 B.n369 B.n6 585
R224 B.n316 B.n5 585
R225 B.n370 B.n5 585
R226 B.n315 B.n314 585
R227 B.n314 B.n4 585
R228 B.n313 B.n135 585
R229 B.n313 B.n312 585
R230 B.n303 B.n136 585
R231 B.n137 B.n136 585
R232 B.n305 B.n304 585
R233 B.n306 B.n305 585
R234 B.n302 B.n142 585
R235 B.n142 B.n141 585
R236 B.n301 B.n300 585
R237 B.n300 B.n299 585
R238 B.n144 B.n143 585
R239 B.n145 B.n144 585
R240 B.n292 B.n291 585
R241 B.n293 B.n292 585
R242 B.n290 B.n150 585
R243 B.n150 B.n149 585
R244 B.n289 B.n288 585
R245 B.n288 B.n287 585
R246 B.n152 B.n151 585
R247 B.n280 B.n152 585
R248 B.n279 B.n278 585
R249 B.n281 B.n279 585
R250 B.n277 B.n157 585
R251 B.n157 B.n156 585
R252 B.n276 B.n275 585
R253 B.n275 B.n274 585
R254 B.n159 B.n158 585
R255 B.n160 B.n159 585
R256 B.n270 B.n269 585
R257 B.n163 B.n162 585
R258 B.n266 B.n265 585
R259 B.n267 B.n266 585
R260 B.n264 B.n183 585
R261 B.n263 B.n262 585
R262 B.n261 B.n260 585
R263 B.n259 B.n258 585
R264 B.n257 B.n256 585
R265 B.n255 B.n254 585
R266 B.n253 B.n252 585
R267 B.n251 B.n250 585
R268 B.n249 B.n248 585
R269 B.n247 B.n246 585
R270 B.n245 B.n244 585
R271 B.n243 B.n242 585
R272 B.n241 B.n240 585
R273 B.n238 B.n237 585
R274 B.n236 B.n235 585
R275 B.n234 B.n233 585
R276 B.n232 B.n231 585
R277 B.n230 B.n229 585
R278 B.n228 B.n227 585
R279 B.n226 B.n225 585
R280 B.n224 B.n223 585
R281 B.n222 B.n221 585
R282 B.n220 B.n219 585
R283 B.n218 B.n217 585
R284 B.n216 B.n215 585
R285 B.n214 B.n213 585
R286 B.n212 B.n211 585
R287 B.n210 B.n209 585
R288 B.n208 B.n207 585
R289 B.n206 B.n205 585
R290 B.n204 B.n203 585
R291 B.n202 B.n201 585
R292 B.n200 B.n199 585
R293 B.n198 B.n197 585
R294 B.n196 B.n195 585
R295 B.n194 B.n193 585
R296 B.n192 B.n191 585
R297 B.n190 B.n189 585
R298 B.n271 B.n161 585
R299 B.n161 B.n160 585
R300 B.n273 B.n272 585
R301 B.n274 B.n273 585
R302 B.n155 B.n154 585
R303 B.n156 B.n155 585
R304 B.n283 B.n282 585
R305 B.n282 B.n281 585
R306 B.n284 B.n153 585
R307 B.n280 B.n153 585
R308 B.n286 B.n285 585
R309 B.n287 B.n286 585
R310 B.n148 B.n147 585
R311 B.n149 B.n148 585
R312 B.n295 B.n294 585
R313 B.n294 B.n293 585
R314 B.n296 B.n146 585
R315 B.n146 B.n145 585
R316 B.n298 B.n297 585
R317 B.n299 B.n298 585
R318 B.n140 B.n139 585
R319 B.n141 B.n140 585
R320 B.n308 B.n307 585
R321 B.n307 B.n306 585
R322 B.n309 B.n138 585
R323 B.n138 B.n137 585
R324 B.n311 B.n310 585
R325 B.n312 B.n311 585
R326 B.n2 B.n0 585
R327 B.n4 B.n2 585
R328 B.n3 B.n1 585
R329 B.n369 B.n3 585
R330 B.n367 B.n366 585
R331 B.n368 B.n367 585
R332 B.n365 B.n9 585
R333 B.n9 B.n8 585
R334 B.n364 B.n363 585
R335 B.n363 B.n362 585
R336 B.n11 B.n10 585
R337 B.n361 B.n11 585
R338 B.n359 B.n358 585
R339 B.n360 B.n359 585
R340 B.n357 B.n16 585
R341 B.n16 B.n15 585
R342 B.n356 B.n355 585
R343 B.n355 B.n354 585
R344 B.n18 B.n17 585
R345 B.n353 B.n18 585
R346 B.n351 B.n350 585
R347 B.n352 B.n351 585
R348 B.n349 B.n22 585
R349 B.n25 B.n22 585
R350 B.n348 B.n347 585
R351 B.n347 B.n346 585
R352 B.n24 B.n23 585
R353 B.n345 B.n24 585
R354 B.n343 B.n342 585
R355 B.n344 B.n343 585
R356 B.n341 B.n30 585
R357 B.n30 B.n29 585
R358 B.n372 B.n371 585
R359 B.n371 B.n370 585
R360 B.n269 B.n161 569.379
R361 B.n339 B.n30 569.379
R362 B.n189 B.n159 569.379
R363 B.n336 B.n53 569.379
R364 B.n186 B.t2 290.769
R365 B.n184 B.t6 290.769
R366 B.n56 B.t13 290.769
R367 B.n54 B.t9 290.769
R368 B.n337 B.n51 256.663
R369 B.n337 B.n50 256.663
R370 B.n337 B.n49 256.663
R371 B.n337 B.n48 256.663
R372 B.n337 B.n47 256.663
R373 B.n337 B.n46 256.663
R374 B.n337 B.n45 256.663
R375 B.n337 B.n44 256.663
R376 B.n337 B.n43 256.663
R377 B.n337 B.n42 256.663
R378 B.n337 B.n41 256.663
R379 B.n337 B.n40 256.663
R380 B.n337 B.n39 256.663
R381 B.n337 B.n38 256.663
R382 B.n337 B.n37 256.663
R383 B.n337 B.n36 256.663
R384 B.n337 B.n35 256.663
R385 B.n337 B.n34 256.663
R386 B.n337 B.n33 256.663
R387 B.n338 B.n337 256.663
R388 B.n268 B.n267 256.663
R389 B.n267 B.n164 256.663
R390 B.n267 B.n165 256.663
R391 B.n267 B.n166 256.663
R392 B.n267 B.n167 256.663
R393 B.n267 B.n168 256.663
R394 B.n267 B.n169 256.663
R395 B.n267 B.n170 256.663
R396 B.n267 B.n171 256.663
R397 B.n267 B.n172 256.663
R398 B.n267 B.n173 256.663
R399 B.n267 B.n174 256.663
R400 B.n267 B.n175 256.663
R401 B.n267 B.n176 256.663
R402 B.n267 B.n177 256.663
R403 B.n267 B.n178 256.663
R404 B.n267 B.n179 256.663
R405 B.n267 B.n180 256.663
R406 B.n267 B.n181 256.663
R407 B.n267 B.n182 256.663
R408 B.n267 B.n160 179.145
R409 B.n337 B.n29 179.145
R410 B.n273 B.n161 163.367
R411 B.n273 B.n155 163.367
R412 B.n282 B.n155 163.367
R413 B.n282 B.n153 163.367
R414 B.n286 B.n153 163.367
R415 B.n286 B.n148 163.367
R416 B.n294 B.n148 163.367
R417 B.n294 B.n146 163.367
R418 B.n298 B.n146 163.367
R419 B.n298 B.n140 163.367
R420 B.n307 B.n140 163.367
R421 B.n307 B.n138 163.367
R422 B.n311 B.n138 163.367
R423 B.n311 B.n2 163.367
R424 B.n371 B.n2 163.367
R425 B.n371 B.n3 163.367
R426 B.n367 B.n3 163.367
R427 B.n367 B.n9 163.367
R428 B.n363 B.n9 163.367
R429 B.n363 B.n11 163.367
R430 B.n359 B.n11 163.367
R431 B.n359 B.n16 163.367
R432 B.n355 B.n16 163.367
R433 B.n355 B.n18 163.367
R434 B.n351 B.n18 163.367
R435 B.n351 B.n22 163.367
R436 B.n347 B.n22 163.367
R437 B.n347 B.n24 163.367
R438 B.n343 B.n24 163.367
R439 B.n343 B.n30 163.367
R440 B.n266 B.n163 163.367
R441 B.n266 B.n183 163.367
R442 B.n262 B.n261 163.367
R443 B.n258 B.n257 163.367
R444 B.n254 B.n253 163.367
R445 B.n250 B.n249 163.367
R446 B.n246 B.n245 163.367
R447 B.n242 B.n241 163.367
R448 B.n237 B.n236 163.367
R449 B.n233 B.n232 163.367
R450 B.n229 B.n228 163.367
R451 B.n225 B.n224 163.367
R452 B.n221 B.n220 163.367
R453 B.n217 B.n216 163.367
R454 B.n213 B.n212 163.367
R455 B.n209 B.n208 163.367
R456 B.n205 B.n204 163.367
R457 B.n201 B.n200 163.367
R458 B.n197 B.n196 163.367
R459 B.n193 B.n192 163.367
R460 B.n275 B.n159 163.367
R461 B.n275 B.n157 163.367
R462 B.n279 B.n157 163.367
R463 B.n279 B.n152 163.367
R464 B.n288 B.n152 163.367
R465 B.n288 B.n150 163.367
R466 B.n292 B.n150 163.367
R467 B.n292 B.n144 163.367
R468 B.n300 B.n144 163.367
R469 B.n300 B.n142 163.367
R470 B.n305 B.n142 163.367
R471 B.n305 B.n136 163.367
R472 B.n313 B.n136 163.367
R473 B.n314 B.n313 163.367
R474 B.n314 B.n5 163.367
R475 B.n6 B.n5 163.367
R476 B.n7 B.n6 163.367
R477 B.n319 B.n7 163.367
R478 B.n319 B.n12 163.367
R479 B.n13 B.n12 163.367
R480 B.n14 B.n13 163.367
R481 B.n324 B.n14 163.367
R482 B.n324 B.n19 163.367
R483 B.n20 B.n19 163.367
R484 B.n21 B.n20 163.367
R485 B.n329 B.n21 163.367
R486 B.n329 B.n26 163.367
R487 B.n27 B.n26 163.367
R488 B.n28 B.n27 163.367
R489 B.n53 B.n28 163.367
R490 B.n59 B.n32 163.367
R491 B.n63 B.n62 163.367
R492 B.n67 B.n66 163.367
R493 B.n71 B.n70 163.367
R494 B.n75 B.n74 163.367
R495 B.n79 B.n78 163.367
R496 B.n83 B.n82 163.367
R497 B.n87 B.n86 163.367
R498 B.n91 B.n90 163.367
R499 B.n95 B.n94 163.367
R500 B.n99 B.n98 163.367
R501 B.n103 B.n102 163.367
R502 B.n108 B.n107 163.367
R503 B.n112 B.n111 163.367
R504 B.n116 B.n115 163.367
R505 B.n120 B.n119 163.367
R506 B.n124 B.n123 163.367
R507 B.n128 B.n127 163.367
R508 B.n132 B.n131 163.367
R509 B.n336 B.n52 163.367
R510 B.n186 B.t5 156.422
R511 B.n54 B.t11 156.422
R512 B.n184 B.t8 156.422
R513 B.n56 B.t14 156.422
R514 B.n187 B.t4 132.956
R515 B.n55 B.t12 132.956
R516 B.n185 B.t7 132.954
R517 B.n57 B.t15 132.954
R518 B.n274 B.n160 87.6396
R519 B.n274 B.n156 87.6396
R520 B.n281 B.n156 87.6396
R521 B.n281 B.n280 87.6396
R522 B.n287 B.n149 87.6396
R523 B.n293 B.n149 87.6396
R524 B.n293 B.n145 87.6396
R525 B.n299 B.n145 87.6396
R526 B.n299 B.n141 87.6396
R527 B.n306 B.n141 87.6396
R528 B.n312 B.n137 87.6396
R529 B.n312 B.n4 87.6396
R530 B.n370 B.n4 87.6396
R531 B.n370 B.n369 87.6396
R532 B.n369 B.n368 87.6396
R533 B.n368 B.n8 87.6396
R534 B.n362 B.n361 87.6396
R535 B.n361 B.n360 87.6396
R536 B.n360 B.n15 87.6396
R537 B.n354 B.n15 87.6396
R538 B.n354 B.n353 87.6396
R539 B.n353 B.n352 87.6396
R540 B.n346 B.n25 87.6396
R541 B.n346 B.n345 87.6396
R542 B.n345 B.n344 87.6396
R543 B.n344 B.n29 87.6396
R544 B.n280 B.t3 74.7515
R545 B.n25 B.t10 74.7515
R546 B.n269 B.n268 71.676
R547 B.n183 B.n164 71.676
R548 B.n261 B.n165 71.676
R549 B.n257 B.n166 71.676
R550 B.n253 B.n167 71.676
R551 B.n249 B.n168 71.676
R552 B.n245 B.n169 71.676
R553 B.n241 B.n170 71.676
R554 B.n236 B.n171 71.676
R555 B.n232 B.n172 71.676
R556 B.n228 B.n173 71.676
R557 B.n224 B.n174 71.676
R558 B.n220 B.n175 71.676
R559 B.n216 B.n176 71.676
R560 B.n212 B.n177 71.676
R561 B.n208 B.n178 71.676
R562 B.n204 B.n179 71.676
R563 B.n200 B.n180 71.676
R564 B.n196 B.n181 71.676
R565 B.n192 B.n182 71.676
R566 B.n339 B.n338 71.676
R567 B.n59 B.n33 71.676
R568 B.n63 B.n34 71.676
R569 B.n67 B.n35 71.676
R570 B.n71 B.n36 71.676
R571 B.n75 B.n37 71.676
R572 B.n79 B.n38 71.676
R573 B.n83 B.n39 71.676
R574 B.n87 B.n40 71.676
R575 B.n91 B.n41 71.676
R576 B.n95 B.n42 71.676
R577 B.n99 B.n43 71.676
R578 B.n103 B.n44 71.676
R579 B.n108 B.n45 71.676
R580 B.n112 B.n46 71.676
R581 B.n116 B.n47 71.676
R582 B.n120 B.n48 71.676
R583 B.n124 B.n49 71.676
R584 B.n128 B.n50 71.676
R585 B.n132 B.n51 71.676
R586 B.n52 B.n51 71.676
R587 B.n131 B.n50 71.676
R588 B.n127 B.n49 71.676
R589 B.n123 B.n48 71.676
R590 B.n119 B.n47 71.676
R591 B.n115 B.n46 71.676
R592 B.n111 B.n45 71.676
R593 B.n107 B.n44 71.676
R594 B.n102 B.n43 71.676
R595 B.n98 B.n42 71.676
R596 B.n94 B.n41 71.676
R597 B.n90 B.n40 71.676
R598 B.n86 B.n39 71.676
R599 B.n82 B.n38 71.676
R600 B.n78 B.n37 71.676
R601 B.n74 B.n36 71.676
R602 B.n70 B.n35 71.676
R603 B.n66 B.n34 71.676
R604 B.n62 B.n33 71.676
R605 B.n338 B.n32 71.676
R606 B.n268 B.n163 71.676
R607 B.n262 B.n164 71.676
R608 B.n258 B.n165 71.676
R609 B.n254 B.n166 71.676
R610 B.n250 B.n167 71.676
R611 B.n246 B.n168 71.676
R612 B.n242 B.n169 71.676
R613 B.n237 B.n170 71.676
R614 B.n233 B.n171 71.676
R615 B.n229 B.n172 71.676
R616 B.n225 B.n173 71.676
R617 B.n221 B.n174 71.676
R618 B.n217 B.n175 71.676
R619 B.n213 B.n176 71.676
R620 B.n209 B.n177 71.676
R621 B.n205 B.n178 71.676
R622 B.n201 B.n179 71.676
R623 B.n197 B.n180 71.676
R624 B.n193 B.n181 71.676
R625 B.n189 B.n182 71.676
R626 B.n188 B.n187 59.5399
R627 B.n239 B.n185 59.5399
R628 B.n58 B.n57 59.5399
R629 B.n105 B.n55 59.5399
R630 B.n306 B.t1 54.1306
R631 B.n362 B.t0 54.1306
R632 B.n341 B.n340 36.9956
R633 B.n335 B.n334 36.9956
R634 B.n190 B.n158 36.9956
R635 B.n271 B.n270 36.9956
R636 B.t1 B.n137 33.5096
R637 B.t0 B.n8 33.5096
R638 B.n187 B.n186 23.4672
R639 B.n185 B.n184 23.4672
R640 B.n57 B.n56 23.4672
R641 B.n55 B.n54 23.4672
R642 B B.n372 18.0485
R643 B.n287 B.t3 12.8886
R644 B.n352 B.t10 12.8886
R645 B.n340 B.n31 10.6151
R646 B.n60 B.n31 10.6151
R647 B.n61 B.n60 10.6151
R648 B.n64 B.n61 10.6151
R649 B.n65 B.n64 10.6151
R650 B.n68 B.n65 10.6151
R651 B.n69 B.n68 10.6151
R652 B.n72 B.n69 10.6151
R653 B.n73 B.n72 10.6151
R654 B.n76 B.n73 10.6151
R655 B.n77 B.n76 10.6151
R656 B.n80 B.n77 10.6151
R657 B.n81 B.n80 10.6151
R658 B.n84 B.n81 10.6151
R659 B.n85 B.n84 10.6151
R660 B.n89 B.n88 10.6151
R661 B.n92 B.n89 10.6151
R662 B.n93 B.n92 10.6151
R663 B.n96 B.n93 10.6151
R664 B.n97 B.n96 10.6151
R665 B.n100 B.n97 10.6151
R666 B.n101 B.n100 10.6151
R667 B.n104 B.n101 10.6151
R668 B.n109 B.n106 10.6151
R669 B.n110 B.n109 10.6151
R670 B.n113 B.n110 10.6151
R671 B.n114 B.n113 10.6151
R672 B.n117 B.n114 10.6151
R673 B.n118 B.n117 10.6151
R674 B.n121 B.n118 10.6151
R675 B.n122 B.n121 10.6151
R676 B.n125 B.n122 10.6151
R677 B.n126 B.n125 10.6151
R678 B.n129 B.n126 10.6151
R679 B.n130 B.n129 10.6151
R680 B.n133 B.n130 10.6151
R681 B.n134 B.n133 10.6151
R682 B.n335 B.n134 10.6151
R683 B.n276 B.n158 10.6151
R684 B.n277 B.n276 10.6151
R685 B.n278 B.n277 10.6151
R686 B.n278 B.n151 10.6151
R687 B.n289 B.n151 10.6151
R688 B.n290 B.n289 10.6151
R689 B.n291 B.n290 10.6151
R690 B.n291 B.n143 10.6151
R691 B.n301 B.n143 10.6151
R692 B.n302 B.n301 10.6151
R693 B.n304 B.n302 10.6151
R694 B.n304 B.n303 10.6151
R695 B.n303 B.n135 10.6151
R696 B.n315 B.n135 10.6151
R697 B.n316 B.n315 10.6151
R698 B.n317 B.n316 10.6151
R699 B.n318 B.n317 10.6151
R700 B.n320 B.n318 10.6151
R701 B.n321 B.n320 10.6151
R702 B.n322 B.n321 10.6151
R703 B.n323 B.n322 10.6151
R704 B.n325 B.n323 10.6151
R705 B.n326 B.n325 10.6151
R706 B.n327 B.n326 10.6151
R707 B.n328 B.n327 10.6151
R708 B.n330 B.n328 10.6151
R709 B.n331 B.n330 10.6151
R710 B.n332 B.n331 10.6151
R711 B.n333 B.n332 10.6151
R712 B.n334 B.n333 10.6151
R713 B.n270 B.n162 10.6151
R714 B.n265 B.n162 10.6151
R715 B.n265 B.n264 10.6151
R716 B.n264 B.n263 10.6151
R717 B.n263 B.n260 10.6151
R718 B.n260 B.n259 10.6151
R719 B.n259 B.n256 10.6151
R720 B.n256 B.n255 10.6151
R721 B.n255 B.n252 10.6151
R722 B.n252 B.n251 10.6151
R723 B.n251 B.n248 10.6151
R724 B.n248 B.n247 10.6151
R725 B.n247 B.n244 10.6151
R726 B.n244 B.n243 10.6151
R727 B.n243 B.n240 10.6151
R728 B.n238 B.n235 10.6151
R729 B.n235 B.n234 10.6151
R730 B.n234 B.n231 10.6151
R731 B.n231 B.n230 10.6151
R732 B.n230 B.n227 10.6151
R733 B.n227 B.n226 10.6151
R734 B.n226 B.n223 10.6151
R735 B.n223 B.n222 10.6151
R736 B.n219 B.n218 10.6151
R737 B.n218 B.n215 10.6151
R738 B.n215 B.n214 10.6151
R739 B.n214 B.n211 10.6151
R740 B.n211 B.n210 10.6151
R741 B.n210 B.n207 10.6151
R742 B.n207 B.n206 10.6151
R743 B.n206 B.n203 10.6151
R744 B.n203 B.n202 10.6151
R745 B.n202 B.n199 10.6151
R746 B.n199 B.n198 10.6151
R747 B.n198 B.n195 10.6151
R748 B.n195 B.n194 10.6151
R749 B.n194 B.n191 10.6151
R750 B.n191 B.n190 10.6151
R751 B.n272 B.n271 10.6151
R752 B.n272 B.n154 10.6151
R753 B.n283 B.n154 10.6151
R754 B.n284 B.n283 10.6151
R755 B.n285 B.n284 10.6151
R756 B.n285 B.n147 10.6151
R757 B.n295 B.n147 10.6151
R758 B.n296 B.n295 10.6151
R759 B.n297 B.n296 10.6151
R760 B.n297 B.n139 10.6151
R761 B.n308 B.n139 10.6151
R762 B.n309 B.n308 10.6151
R763 B.n310 B.n309 10.6151
R764 B.n310 B.n0 10.6151
R765 B.n366 B.n1 10.6151
R766 B.n366 B.n365 10.6151
R767 B.n365 B.n364 10.6151
R768 B.n364 B.n10 10.6151
R769 B.n358 B.n10 10.6151
R770 B.n358 B.n357 10.6151
R771 B.n357 B.n356 10.6151
R772 B.n356 B.n17 10.6151
R773 B.n350 B.n17 10.6151
R774 B.n350 B.n349 10.6151
R775 B.n349 B.n348 10.6151
R776 B.n348 B.n23 10.6151
R777 B.n342 B.n23 10.6151
R778 B.n342 B.n341 10.6151
R779 B.n88 B.n58 7.18099
R780 B.n105 B.n104 7.18099
R781 B.n239 B.n238 7.18099
R782 B.n222 B.n188 7.18099
R783 B.n85 B.n58 3.43465
R784 B.n106 B.n105 3.43465
R785 B.n240 B.n239 3.43465
R786 B.n219 B.n188 3.43465
R787 B.n372 B.n0 2.81026
R788 B.n372 B.n1 2.81026
R789 VP.n0 VP.t0 328.146
R790 VP.n0 VP.t1 294.673
R791 VP VP.n0 0.0516364
R792 VDD1.n10 VDD1.n0 289.615
R793 VDD1.n25 VDD1.n15 289.615
R794 VDD1.n11 VDD1.n10 185
R795 VDD1.n9 VDD1.n8 185
R796 VDD1.n4 VDD1.n3 185
R797 VDD1.n19 VDD1.n18 185
R798 VDD1.n24 VDD1.n23 185
R799 VDD1.n26 VDD1.n25 185
R800 VDD1.n5 VDD1.t1 148.606
R801 VDD1.n20 VDD1.t0 148.606
R802 VDD1.n10 VDD1.n9 104.615
R803 VDD1.n9 VDD1.n3 104.615
R804 VDD1.n24 VDD1.n18 104.615
R805 VDD1.n25 VDD1.n24 104.615
R806 VDD1 VDD1.n29 80.533
R807 VDD1.t1 VDD1.n3 52.3082
R808 VDD1.t0 VDD1.n18 52.3082
R809 VDD1 VDD1.n14 51.5104
R810 VDD1.n5 VDD1.n4 15.5966
R811 VDD1.n20 VDD1.n19 15.5966
R812 VDD1.n8 VDD1.n7 12.8005
R813 VDD1.n23 VDD1.n22 12.8005
R814 VDD1.n11 VDD1.n2 12.0247
R815 VDD1.n26 VDD1.n17 12.0247
R816 VDD1.n12 VDD1.n0 11.249
R817 VDD1.n27 VDD1.n15 11.249
R818 VDD1.n14 VDD1.n13 9.45567
R819 VDD1.n29 VDD1.n28 9.45567
R820 VDD1.n13 VDD1.n12 9.3005
R821 VDD1.n2 VDD1.n1 9.3005
R822 VDD1.n7 VDD1.n6 9.3005
R823 VDD1.n28 VDD1.n27 9.3005
R824 VDD1.n17 VDD1.n16 9.3005
R825 VDD1.n22 VDD1.n21 9.3005
R826 VDD1.n6 VDD1.n5 4.46457
R827 VDD1.n21 VDD1.n20 4.46457
R828 VDD1.n14 VDD1.n0 2.71565
R829 VDD1.n29 VDD1.n15 2.71565
R830 VDD1.n12 VDD1.n11 1.93989
R831 VDD1.n27 VDD1.n26 1.93989
R832 VDD1.n8 VDD1.n2 1.16414
R833 VDD1.n23 VDD1.n17 1.16414
R834 VDD1.n7 VDD1.n4 0.388379
R835 VDD1.n22 VDD1.n19 0.388379
R836 VDD1.n13 VDD1.n1 0.155672
R837 VDD1.n6 VDD1.n1 0.155672
R838 VDD1.n21 VDD1.n16 0.155672
R839 VDD1.n28 VDD1.n16 0.155672
C0 VP VTAIL 0.744978f
C1 VDD2 VDD1 0.477633f
C2 VDD2 VN 0.755168f
C3 VP VDD1 0.866482f
C4 VP VN 3.02481f
C5 VDD1 VTAIL 2.40387f
C6 VTAIL VN 0.73075f
C7 VDD2 VP 0.266838f
C8 VDD2 VTAIL 2.444f
C9 VDD1 VN 0.15385f
C10 VDD2 B 2.217465f
C11 VDD1 B 3.50141f
C12 VTAIL B 2.956477f
C13 VN B 5.7362f
C14 VP B 3.540668f
C15 VDD1.n0 B 0.021488f
C16 VDD1.n1 B 0.015587f
C17 VDD1.n2 B 0.008376f
C18 VDD1.n3 B 0.014848f
C19 VDD1.n4 B 0.011544f
C20 VDD1.t1 B 0.033496f
C21 VDD1.n5 B 0.058022f
C22 VDD1.n6 B 0.170379f
C23 VDD1.n7 B 0.008376f
C24 VDD1.n8 B 0.008868f
C25 VDD1.n9 B 0.019797f
C26 VDD1.n10 B 0.042113f
C27 VDD1.n11 B 0.008868f
C28 VDD1.n12 B 0.008376f
C29 VDD1.n13 B 0.038583f
C30 VDD1.n14 B 0.034602f
C31 VDD1.n15 B 0.021488f
C32 VDD1.n16 B 0.015587f
C33 VDD1.n17 B 0.008376f
C34 VDD1.n18 B 0.014848f
C35 VDD1.n19 B 0.011544f
C36 VDD1.t0 B 0.033496f
C37 VDD1.n20 B 0.058022f
C38 VDD1.n21 B 0.170379f
C39 VDD1.n22 B 0.008376f
C40 VDD1.n23 B 0.008868f
C41 VDD1.n24 B 0.019797f
C42 VDD1.n25 B 0.042113f
C43 VDD1.n26 B 0.008868f
C44 VDD1.n27 B 0.008376f
C45 VDD1.n28 B 0.038583f
C46 VDD1.n29 B 0.237651f
C47 VP.t0 B 0.511463f
C48 VP.t1 B 0.401425f
C49 VP.n0 B 2.07036f
C50 VDD2.n0 B 0.022016f
C51 VDD2.n1 B 0.01597f
C52 VDD2.n2 B 0.008582f
C53 VDD2.n3 B 0.015213f
C54 VDD2.n4 B 0.011828f
C55 VDD2.t0 B 0.034319f
C56 VDD2.n5 B 0.059448f
C57 VDD2.n6 B 0.174567f
C58 VDD2.n7 B 0.008582f
C59 VDD2.n8 B 0.009086f
C60 VDD2.n9 B 0.020284f
C61 VDD2.n10 B 0.043148f
C62 VDD2.n11 B 0.009086f
C63 VDD2.n12 B 0.008582f
C64 VDD2.n13 B 0.039531f
C65 VDD2.n14 B 0.225636f
C66 VDD2.n15 B 0.022016f
C67 VDD2.n16 B 0.01597f
C68 VDD2.n17 B 0.008582f
C69 VDD2.n18 B 0.015213f
C70 VDD2.n19 B 0.011828f
C71 VDD2.t1 B 0.034319f
C72 VDD2.n20 B 0.059448f
C73 VDD2.n21 B 0.174567f
C74 VDD2.n22 B 0.008582f
C75 VDD2.n23 B 0.009086f
C76 VDD2.n24 B 0.020284f
C77 VDD2.n25 B 0.043148f
C78 VDD2.n26 B 0.009086f
C79 VDD2.n27 B 0.008582f
C80 VDD2.n28 B 0.039531f
C81 VDD2.n29 B 0.035151f
C82 VDD2.n30 B 1.13504f
C83 VTAIL.n0 B 0.026091f
C84 VTAIL.n1 B 0.018926f
C85 VTAIL.n2 B 0.01017f
C86 VTAIL.n3 B 0.018028f
C87 VTAIL.n4 B 0.014017f
C88 VTAIL.t2 B 0.040671f
C89 VTAIL.n5 B 0.070451f
C90 VTAIL.n6 B 0.206878f
C91 VTAIL.n7 B 0.01017f
C92 VTAIL.n8 B 0.010768f
C93 VTAIL.n9 B 0.024038f
C94 VTAIL.n10 B 0.051135f
C95 VTAIL.n11 B 0.010768f
C96 VTAIL.n12 B 0.01017f
C97 VTAIL.n13 B 0.046848f
C98 VTAIL.n14 B 0.028611f
C99 VTAIL.n15 B 0.621711f
C100 VTAIL.n16 B 0.026091f
C101 VTAIL.n17 B 0.018926f
C102 VTAIL.n18 B 0.01017f
C103 VTAIL.n19 B 0.018028f
C104 VTAIL.n20 B 0.014017f
C105 VTAIL.t1 B 0.040671f
C106 VTAIL.n21 B 0.070451f
C107 VTAIL.n22 B 0.206878f
C108 VTAIL.n23 B 0.01017f
C109 VTAIL.n24 B 0.010768f
C110 VTAIL.n25 B 0.024038f
C111 VTAIL.n26 B 0.051135f
C112 VTAIL.n27 B 0.010768f
C113 VTAIL.n28 B 0.01017f
C114 VTAIL.n29 B 0.046848f
C115 VTAIL.n30 B 0.028611f
C116 VTAIL.n31 B 0.634065f
C117 VTAIL.n32 B 0.026091f
C118 VTAIL.n33 B 0.018926f
C119 VTAIL.n34 B 0.01017f
C120 VTAIL.n35 B 0.018028f
C121 VTAIL.n36 B 0.014017f
C122 VTAIL.t3 B 0.040671f
C123 VTAIL.n37 B 0.070451f
C124 VTAIL.n38 B 0.206878f
C125 VTAIL.n39 B 0.01017f
C126 VTAIL.n40 B 0.010768f
C127 VTAIL.n41 B 0.024038f
C128 VTAIL.n42 B 0.051135f
C129 VTAIL.n43 B 0.010768f
C130 VTAIL.n44 B 0.01017f
C131 VTAIL.n45 B 0.046848f
C132 VTAIL.n46 B 0.028611f
C133 VTAIL.n47 B 0.570454f
C134 VTAIL.n48 B 0.026091f
C135 VTAIL.n49 B 0.018926f
C136 VTAIL.n50 B 0.01017f
C137 VTAIL.n51 B 0.018028f
C138 VTAIL.n52 B 0.014017f
C139 VTAIL.t0 B 0.040671f
C140 VTAIL.n53 B 0.070451f
C141 VTAIL.n54 B 0.206878f
C142 VTAIL.n55 B 0.01017f
C143 VTAIL.n56 B 0.010768f
C144 VTAIL.n57 B 0.024038f
C145 VTAIL.n58 B 0.051135f
C146 VTAIL.n59 B 0.010768f
C147 VTAIL.n60 B 0.01017f
C148 VTAIL.n61 B 0.046848f
C149 VTAIL.n62 B 0.028611f
C150 VTAIL.n63 B 0.522351f
C151 VN.t1 B 0.394701f
C152 VN.t0 B 0.506439f
.ends

