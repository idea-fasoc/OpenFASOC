* NGSPICE file created from diff_pair_sample_1169.ext - technology: sky130A

.subckt diff_pair_sample_1169 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=2.48985 ps=15.42 w=15.09 l=2.62
X1 VTAIL.t6 VP.t1 VDD1.t3 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=2.48985 ps=15.42 w=15.09 l=2.62
X2 B.t11 B.t9 B.t10 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=0 ps=0 w=15.09 l=2.62
X3 VDD2.t3 VN.t0 VTAIL.t0 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=2.48985 pd=15.42 as=5.8851 ps=30.96 w=15.09 l=2.62
X4 VDD1.t1 VP.t2 VTAIL.t5 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=2.48985 pd=15.42 as=5.8851 ps=30.96 w=15.09 l=2.62
X5 VDD1.t2 VP.t3 VTAIL.t4 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=2.48985 pd=15.42 as=5.8851 ps=30.96 w=15.09 l=2.62
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=2.48985 pd=15.42 as=5.8851 ps=30.96 w=15.09 l=2.62
X7 VTAIL.t2 VN.t2 VDD2.t1 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=2.48985 ps=15.42 w=15.09 l=2.62
X8 B.t8 B.t6 B.t7 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=0 ps=0 w=15.09 l=2.62
X9 B.t5 B.t3 B.t4 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=0 ps=0 w=15.09 l=2.62
X10 VTAIL.t3 VN.t3 VDD2.t0 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=2.48985 ps=15.42 w=15.09 l=2.62
X11 B.t2 B.t0 B.t1 w_n2740_n3986# sky130_fd_pr__pfet_01v8 ad=5.8851 pd=30.96 as=0 ps=0 w=15.09 l=2.62
R0 VP.n4 VP.t0 175.141
R1 VP.n4 VP.t3 174.363
R2 VP.n14 VP.n0 161.3
R3 VP.n13 VP.n12 161.3
R4 VP.n11 VP.n1 161.3
R5 VP.n10 VP.n9 161.3
R6 VP.n8 VP.n2 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n3 VP.t1 138.805
R9 VP.n15 VP.t2 138.805
R10 VP.n5 VP.n3 99.7463
R11 VP.n16 VP.n15 99.7463
R12 VP.n9 VP.n1 56.5193
R13 VP.n5 VP.n4 53.0403
R14 VP.n8 VP.n7 24.4675
R15 VP.n9 VP.n8 24.4675
R16 VP.n13 VP.n1 24.4675
R17 VP.n14 VP.n13 24.4675
R18 VP.n7 VP.n3 11.0107
R19 VP.n15 VP.n14 11.0107
R20 VP.n6 VP.n5 0.278367
R21 VP.n16 VP.n0 0.278367
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153454
R28 VDD1 VDD1.n1 117.127
R29 VDD1 VDD1.n0 72.3086
R30 VDD1.n0 VDD1.t0 2.15458
R31 VDD1.n0 VDD1.t2 2.15458
R32 VDD1.n1 VDD1.t3 2.15458
R33 VDD1.n1 VDD1.t1 2.15458
R34 VTAIL.n5 VTAIL.t7 57.7259
R35 VTAIL.n4 VTAIL.t1 57.7259
R36 VTAIL.n3 VTAIL.t3 57.7259
R37 VTAIL.n7 VTAIL.t0 57.7256
R38 VTAIL.n0 VTAIL.t2 57.7256
R39 VTAIL.n1 VTAIL.t5 57.7256
R40 VTAIL.n2 VTAIL.t6 57.7256
R41 VTAIL.n6 VTAIL.t4 57.7256
R42 VTAIL.n7 VTAIL.n6 27.9186
R43 VTAIL.n3 VTAIL.n2 27.9186
R44 VTAIL.n4 VTAIL.n3 2.5436
R45 VTAIL.n6 VTAIL.n5 2.5436
R46 VTAIL.n2 VTAIL.n1 2.5436
R47 VTAIL VTAIL.n0 1.33024
R48 VTAIL VTAIL.n7 1.21386
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 B.n512 B.n79 585
R52 B.n514 B.n513 585
R53 B.n515 B.n78 585
R54 B.n517 B.n516 585
R55 B.n518 B.n77 585
R56 B.n520 B.n519 585
R57 B.n521 B.n76 585
R58 B.n523 B.n522 585
R59 B.n524 B.n75 585
R60 B.n526 B.n525 585
R61 B.n527 B.n74 585
R62 B.n529 B.n528 585
R63 B.n530 B.n73 585
R64 B.n532 B.n531 585
R65 B.n533 B.n72 585
R66 B.n535 B.n534 585
R67 B.n536 B.n71 585
R68 B.n538 B.n537 585
R69 B.n539 B.n70 585
R70 B.n541 B.n540 585
R71 B.n542 B.n69 585
R72 B.n544 B.n543 585
R73 B.n545 B.n68 585
R74 B.n547 B.n546 585
R75 B.n548 B.n67 585
R76 B.n550 B.n549 585
R77 B.n551 B.n66 585
R78 B.n553 B.n552 585
R79 B.n554 B.n65 585
R80 B.n556 B.n555 585
R81 B.n557 B.n64 585
R82 B.n559 B.n558 585
R83 B.n560 B.n63 585
R84 B.n562 B.n561 585
R85 B.n563 B.n62 585
R86 B.n565 B.n564 585
R87 B.n566 B.n61 585
R88 B.n568 B.n567 585
R89 B.n569 B.n60 585
R90 B.n571 B.n570 585
R91 B.n572 B.n59 585
R92 B.n574 B.n573 585
R93 B.n575 B.n58 585
R94 B.n577 B.n576 585
R95 B.n578 B.n57 585
R96 B.n580 B.n579 585
R97 B.n581 B.n56 585
R98 B.n583 B.n582 585
R99 B.n584 B.n55 585
R100 B.n586 B.n585 585
R101 B.n587 B.n52 585
R102 B.n590 B.n589 585
R103 B.n591 B.n51 585
R104 B.n593 B.n592 585
R105 B.n594 B.n50 585
R106 B.n596 B.n595 585
R107 B.n597 B.n49 585
R108 B.n599 B.n598 585
R109 B.n600 B.n45 585
R110 B.n602 B.n601 585
R111 B.n603 B.n44 585
R112 B.n605 B.n604 585
R113 B.n606 B.n43 585
R114 B.n608 B.n607 585
R115 B.n609 B.n42 585
R116 B.n611 B.n610 585
R117 B.n612 B.n41 585
R118 B.n614 B.n613 585
R119 B.n615 B.n40 585
R120 B.n617 B.n616 585
R121 B.n618 B.n39 585
R122 B.n620 B.n619 585
R123 B.n621 B.n38 585
R124 B.n623 B.n622 585
R125 B.n624 B.n37 585
R126 B.n626 B.n625 585
R127 B.n627 B.n36 585
R128 B.n629 B.n628 585
R129 B.n630 B.n35 585
R130 B.n632 B.n631 585
R131 B.n633 B.n34 585
R132 B.n635 B.n634 585
R133 B.n636 B.n33 585
R134 B.n638 B.n637 585
R135 B.n639 B.n32 585
R136 B.n641 B.n640 585
R137 B.n642 B.n31 585
R138 B.n644 B.n643 585
R139 B.n645 B.n30 585
R140 B.n647 B.n646 585
R141 B.n648 B.n29 585
R142 B.n650 B.n649 585
R143 B.n651 B.n28 585
R144 B.n653 B.n652 585
R145 B.n654 B.n27 585
R146 B.n656 B.n655 585
R147 B.n657 B.n26 585
R148 B.n659 B.n658 585
R149 B.n660 B.n25 585
R150 B.n662 B.n661 585
R151 B.n663 B.n24 585
R152 B.n665 B.n664 585
R153 B.n666 B.n23 585
R154 B.n668 B.n667 585
R155 B.n669 B.n22 585
R156 B.n671 B.n670 585
R157 B.n672 B.n21 585
R158 B.n674 B.n673 585
R159 B.n675 B.n20 585
R160 B.n677 B.n676 585
R161 B.n678 B.n19 585
R162 B.n511 B.n510 585
R163 B.n509 B.n80 585
R164 B.n508 B.n507 585
R165 B.n506 B.n81 585
R166 B.n505 B.n504 585
R167 B.n503 B.n82 585
R168 B.n502 B.n501 585
R169 B.n500 B.n83 585
R170 B.n499 B.n498 585
R171 B.n497 B.n84 585
R172 B.n496 B.n495 585
R173 B.n494 B.n85 585
R174 B.n493 B.n492 585
R175 B.n491 B.n86 585
R176 B.n490 B.n489 585
R177 B.n488 B.n87 585
R178 B.n487 B.n486 585
R179 B.n485 B.n88 585
R180 B.n484 B.n483 585
R181 B.n482 B.n89 585
R182 B.n481 B.n480 585
R183 B.n479 B.n90 585
R184 B.n478 B.n477 585
R185 B.n476 B.n91 585
R186 B.n475 B.n474 585
R187 B.n473 B.n92 585
R188 B.n472 B.n471 585
R189 B.n470 B.n93 585
R190 B.n469 B.n468 585
R191 B.n467 B.n94 585
R192 B.n466 B.n465 585
R193 B.n464 B.n95 585
R194 B.n463 B.n462 585
R195 B.n461 B.n96 585
R196 B.n460 B.n459 585
R197 B.n458 B.n97 585
R198 B.n457 B.n456 585
R199 B.n455 B.n98 585
R200 B.n454 B.n453 585
R201 B.n452 B.n99 585
R202 B.n451 B.n450 585
R203 B.n449 B.n100 585
R204 B.n448 B.n447 585
R205 B.n446 B.n101 585
R206 B.n445 B.n444 585
R207 B.n443 B.n102 585
R208 B.n442 B.n441 585
R209 B.n440 B.n103 585
R210 B.n439 B.n438 585
R211 B.n437 B.n104 585
R212 B.n436 B.n435 585
R213 B.n434 B.n105 585
R214 B.n433 B.n432 585
R215 B.n431 B.n106 585
R216 B.n430 B.n429 585
R217 B.n428 B.n107 585
R218 B.n427 B.n426 585
R219 B.n425 B.n108 585
R220 B.n424 B.n423 585
R221 B.n422 B.n109 585
R222 B.n421 B.n420 585
R223 B.n419 B.n110 585
R224 B.n418 B.n417 585
R225 B.n416 B.n111 585
R226 B.n415 B.n414 585
R227 B.n413 B.n112 585
R228 B.n412 B.n411 585
R229 B.n410 B.n113 585
R230 B.n409 B.n408 585
R231 B.n238 B.n171 585
R232 B.n240 B.n239 585
R233 B.n241 B.n170 585
R234 B.n243 B.n242 585
R235 B.n244 B.n169 585
R236 B.n246 B.n245 585
R237 B.n247 B.n168 585
R238 B.n249 B.n248 585
R239 B.n250 B.n167 585
R240 B.n252 B.n251 585
R241 B.n253 B.n166 585
R242 B.n255 B.n254 585
R243 B.n256 B.n165 585
R244 B.n258 B.n257 585
R245 B.n259 B.n164 585
R246 B.n261 B.n260 585
R247 B.n262 B.n163 585
R248 B.n264 B.n263 585
R249 B.n265 B.n162 585
R250 B.n267 B.n266 585
R251 B.n268 B.n161 585
R252 B.n270 B.n269 585
R253 B.n271 B.n160 585
R254 B.n273 B.n272 585
R255 B.n274 B.n159 585
R256 B.n276 B.n275 585
R257 B.n277 B.n158 585
R258 B.n279 B.n278 585
R259 B.n280 B.n157 585
R260 B.n282 B.n281 585
R261 B.n283 B.n156 585
R262 B.n285 B.n284 585
R263 B.n286 B.n155 585
R264 B.n288 B.n287 585
R265 B.n289 B.n154 585
R266 B.n291 B.n290 585
R267 B.n292 B.n153 585
R268 B.n294 B.n293 585
R269 B.n295 B.n152 585
R270 B.n297 B.n296 585
R271 B.n298 B.n151 585
R272 B.n300 B.n299 585
R273 B.n301 B.n150 585
R274 B.n303 B.n302 585
R275 B.n304 B.n149 585
R276 B.n306 B.n305 585
R277 B.n307 B.n148 585
R278 B.n309 B.n308 585
R279 B.n310 B.n147 585
R280 B.n312 B.n311 585
R281 B.n313 B.n144 585
R282 B.n316 B.n315 585
R283 B.n317 B.n143 585
R284 B.n319 B.n318 585
R285 B.n320 B.n142 585
R286 B.n322 B.n321 585
R287 B.n323 B.n141 585
R288 B.n325 B.n324 585
R289 B.n326 B.n140 585
R290 B.n331 B.n330 585
R291 B.n332 B.n139 585
R292 B.n334 B.n333 585
R293 B.n335 B.n138 585
R294 B.n337 B.n336 585
R295 B.n338 B.n137 585
R296 B.n340 B.n339 585
R297 B.n341 B.n136 585
R298 B.n343 B.n342 585
R299 B.n344 B.n135 585
R300 B.n346 B.n345 585
R301 B.n347 B.n134 585
R302 B.n349 B.n348 585
R303 B.n350 B.n133 585
R304 B.n352 B.n351 585
R305 B.n353 B.n132 585
R306 B.n355 B.n354 585
R307 B.n356 B.n131 585
R308 B.n358 B.n357 585
R309 B.n359 B.n130 585
R310 B.n361 B.n360 585
R311 B.n362 B.n129 585
R312 B.n364 B.n363 585
R313 B.n365 B.n128 585
R314 B.n367 B.n366 585
R315 B.n368 B.n127 585
R316 B.n370 B.n369 585
R317 B.n371 B.n126 585
R318 B.n373 B.n372 585
R319 B.n374 B.n125 585
R320 B.n376 B.n375 585
R321 B.n377 B.n124 585
R322 B.n379 B.n378 585
R323 B.n380 B.n123 585
R324 B.n382 B.n381 585
R325 B.n383 B.n122 585
R326 B.n385 B.n384 585
R327 B.n386 B.n121 585
R328 B.n388 B.n387 585
R329 B.n389 B.n120 585
R330 B.n391 B.n390 585
R331 B.n392 B.n119 585
R332 B.n394 B.n393 585
R333 B.n395 B.n118 585
R334 B.n397 B.n396 585
R335 B.n398 B.n117 585
R336 B.n400 B.n399 585
R337 B.n401 B.n116 585
R338 B.n403 B.n402 585
R339 B.n404 B.n115 585
R340 B.n406 B.n405 585
R341 B.n407 B.n114 585
R342 B.n237 B.n236 585
R343 B.n235 B.n172 585
R344 B.n234 B.n233 585
R345 B.n232 B.n173 585
R346 B.n231 B.n230 585
R347 B.n229 B.n174 585
R348 B.n228 B.n227 585
R349 B.n226 B.n175 585
R350 B.n225 B.n224 585
R351 B.n223 B.n176 585
R352 B.n222 B.n221 585
R353 B.n220 B.n177 585
R354 B.n219 B.n218 585
R355 B.n217 B.n178 585
R356 B.n216 B.n215 585
R357 B.n214 B.n179 585
R358 B.n213 B.n212 585
R359 B.n211 B.n180 585
R360 B.n210 B.n209 585
R361 B.n208 B.n181 585
R362 B.n207 B.n206 585
R363 B.n205 B.n182 585
R364 B.n204 B.n203 585
R365 B.n202 B.n183 585
R366 B.n201 B.n200 585
R367 B.n199 B.n184 585
R368 B.n198 B.n197 585
R369 B.n196 B.n185 585
R370 B.n195 B.n194 585
R371 B.n193 B.n186 585
R372 B.n192 B.n191 585
R373 B.n190 B.n187 585
R374 B.n189 B.n188 585
R375 B.n2 B.n0 585
R376 B.n729 B.n1 585
R377 B.n728 B.n727 585
R378 B.n726 B.n3 585
R379 B.n725 B.n724 585
R380 B.n723 B.n4 585
R381 B.n722 B.n721 585
R382 B.n720 B.n5 585
R383 B.n719 B.n718 585
R384 B.n717 B.n6 585
R385 B.n716 B.n715 585
R386 B.n714 B.n7 585
R387 B.n713 B.n712 585
R388 B.n711 B.n8 585
R389 B.n710 B.n709 585
R390 B.n708 B.n9 585
R391 B.n707 B.n706 585
R392 B.n705 B.n10 585
R393 B.n704 B.n703 585
R394 B.n702 B.n11 585
R395 B.n701 B.n700 585
R396 B.n699 B.n12 585
R397 B.n698 B.n697 585
R398 B.n696 B.n13 585
R399 B.n695 B.n694 585
R400 B.n693 B.n14 585
R401 B.n692 B.n691 585
R402 B.n690 B.n15 585
R403 B.n689 B.n688 585
R404 B.n687 B.n16 585
R405 B.n686 B.n685 585
R406 B.n684 B.n17 585
R407 B.n683 B.n682 585
R408 B.n681 B.n18 585
R409 B.n680 B.n679 585
R410 B.n731 B.n730 585
R411 B.n238 B.n237 521.33
R412 B.n680 B.n19 521.33
R413 B.n409 B.n114 521.33
R414 B.n512 B.n511 521.33
R415 B.n327 B.t6 346.882
R416 B.n145 B.t0 346.882
R417 B.n46 B.t9 346.882
R418 B.n53 B.t3 346.882
R419 B.n327 B.t8 166.281
R420 B.n53 B.t4 166.281
R421 B.n145 B.t2 166.262
R422 B.n46 B.t10 166.262
R423 B.n237 B.n172 163.367
R424 B.n233 B.n172 163.367
R425 B.n233 B.n232 163.367
R426 B.n232 B.n231 163.367
R427 B.n231 B.n174 163.367
R428 B.n227 B.n174 163.367
R429 B.n227 B.n226 163.367
R430 B.n226 B.n225 163.367
R431 B.n225 B.n176 163.367
R432 B.n221 B.n176 163.367
R433 B.n221 B.n220 163.367
R434 B.n220 B.n219 163.367
R435 B.n219 B.n178 163.367
R436 B.n215 B.n178 163.367
R437 B.n215 B.n214 163.367
R438 B.n214 B.n213 163.367
R439 B.n213 B.n180 163.367
R440 B.n209 B.n180 163.367
R441 B.n209 B.n208 163.367
R442 B.n208 B.n207 163.367
R443 B.n207 B.n182 163.367
R444 B.n203 B.n182 163.367
R445 B.n203 B.n202 163.367
R446 B.n202 B.n201 163.367
R447 B.n201 B.n184 163.367
R448 B.n197 B.n184 163.367
R449 B.n197 B.n196 163.367
R450 B.n196 B.n195 163.367
R451 B.n195 B.n186 163.367
R452 B.n191 B.n186 163.367
R453 B.n191 B.n190 163.367
R454 B.n190 B.n189 163.367
R455 B.n189 B.n2 163.367
R456 B.n730 B.n2 163.367
R457 B.n730 B.n729 163.367
R458 B.n729 B.n728 163.367
R459 B.n728 B.n3 163.367
R460 B.n724 B.n3 163.367
R461 B.n724 B.n723 163.367
R462 B.n723 B.n722 163.367
R463 B.n722 B.n5 163.367
R464 B.n718 B.n5 163.367
R465 B.n718 B.n717 163.367
R466 B.n717 B.n716 163.367
R467 B.n716 B.n7 163.367
R468 B.n712 B.n7 163.367
R469 B.n712 B.n711 163.367
R470 B.n711 B.n710 163.367
R471 B.n710 B.n9 163.367
R472 B.n706 B.n9 163.367
R473 B.n706 B.n705 163.367
R474 B.n705 B.n704 163.367
R475 B.n704 B.n11 163.367
R476 B.n700 B.n11 163.367
R477 B.n700 B.n699 163.367
R478 B.n699 B.n698 163.367
R479 B.n698 B.n13 163.367
R480 B.n694 B.n13 163.367
R481 B.n694 B.n693 163.367
R482 B.n693 B.n692 163.367
R483 B.n692 B.n15 163.367
R484 B.n688 B.n15 163.367
R485 B.n688 B.n687 163.367
R486 B.n687 B.n686 163.367
R487 B.n686 B.n17 163.367
R488 B.n682 B.n17 163.367
R489 B.n682 B.n681 163.367
R490 B.n681 B.n680 163.367
R491 B.n239 B.n238 163.367
R492 B.n239 B.n170 163.367
R493 B.n243 B.n170 163.367
R494 B.n244 B.n243 163.367
R495 B.n245 B.n244 163.367
R496 B.n245 B.n168 163.367
R497 B.n249 B.n168 163.367
R498 B.n250 B.n249 163.367
R499 B.n251 B.n250 163.367
R500 B.n251 B.n166 163.367
R501 B.n255 B.n166 163.367
R502 B.n256 B.n255 163.367
R503 B.n257 B.n256 163.367
R504 B.n257 B.n164 163.367
R505 B.n261 B.n164 163.367
R506 B.n262 B.n261 163.367
R507 B.n263 B.n262 163.367
R508 B.n263 B.n162 163.367
R509 B.n267 B.n162 163.367
R510 B.n268 B.n267 163.367
R511 B.n269 B.n268 163.367
R512 B.n269 B.n160 163.367
R513 B.n273 B.n160 163.367
R514 B.n274 B.n273 163.367
R515 B.n275 B.n274 163.367
R516 B.n275 B.n158 163.367
R517 B.n279 B.n158 163.367
R518 B.n280 B.n279 163.367
R519 B.n281 B.n280 163.367
R520 B.n281 B.n156 163.367
R521 B.n285 B.n156 163.367
R522 B.n286 B.n285 163.367
R523 B.n287 B.n286 163.367
R524 B.n287 B.n154 163.367
R525 B.n291 B.n154 163.367
R526 B.n292 B.n291 163.367
R527 B.n293 B.n292 163.367
R528 B.n293 B.n152 163.367
R529 B.n297 B.n152 163.367
R530 B.n298 B.n297 163.367
R531 B.n299 B.n298 163.367
R532 B.n299 B.n150 163.367
R533 B.n303 B.n150 163.367
R534 B.n304 B.n303 163.367
R535 B.n305 B.n304 163.367
R536 B.n305 B.n148 163.367
R537 B.n309 B.n148 163.367
R538 B.n310 B.n309 163.367
R539 B.n311 B.n310 163.367
R540 B.n311 B.n144 163.367
R541 B.n316 B.n144 163.367
R542 B.n317 B.n316 163.367
R543 B.n318 B.n317 163.367
R544 B.n318 B.n142 163.367
R545 B.n322 B.n142 163.367
R546 B.n323 B.n322 163.367
R547 B.n324 B.n323 163.367
R548 B.n324 B.n140 163.367
R549 B.n331 B.n140 163.367
R550 B.n332 B.n331 163.367
R551 B.n333 B.n332 163.367
R552 B.n333 B.n138 163.367
R553 B.n337 B.n138 163.367
R554 B.n338 B.n337 163.367
R555 B.n339 B.n338 163.367
R556 B.n339 B.n136 163.367
R557 B.n343 B.n136 163.367
R558 B.n344 B.n343 163.367
R559 B.n345 B.n344 163.367
R560 B.n345 B.n134 163.367
R561 B.n349 B.n134 163.367
R562 B.n350 B.n349 163.367
R563 B.n351 B.n350 163.367
R564 B.n351 B.n132 163.367
R565 B.n355 B.n132 163.367
R566 B.n356 B.n355 163.367
R567 B.n357 B.n356 163.367
R568 B.n357 B.n130 163.367
R569 B.n361 B.n130 163.367
R570 B.n362 B.n361 163.367
R571 B.n363 B.n362 163.367
R572 B.n363 B.n128 163.367
R573 B.n367 B.n128 163.367
R574 B.n368 B.n367 163.367
R575 B.n369 B.n368 163.367
R576 B.n369 B.n126 163.367
R577 B.n373 B.n126 163.367
R578 B.n374 B.n373 163.367
R579 B.n375 B.n374 163.367
R580 B.n375 B.n124 163.367
R581 B.n379 B.n124 163.367
R582 B.n380 B.n379 163.367
R583 B.n381 B.n380 163.367
R584 B.n381 B.n122 163.367
R585 B.n385 B.n122 163.367
R586 B.n386 B.n385 163.367
R587 B.n387 B.n386 163.367
R588 B.n387 B.n120 163.367
R589 B.n391 B.n120 163.367
R590 B.n392 B.n391 163.367
R591 B.n393 B.n392 163.367
R592 B.n393 B.n118 163.367
R593 B.n397 B.n118 163.367
R594 B.n398 B.n397 163.367
R595 B.n399 B.n398 163.367
R596 B.n399 B.n116 163.367
R597 B.n403 B.n116 163.367
R598 B.n404 B.n403 163.367
R599 B.n405 B.n404 163.367
R600 B.n405 B.n114 163.367
R601 B.n410 B.n409 163.367
R602 B.n411 B.n410 163.367
R603 B.n411 B.n112 163.367
R604 B.n415 B.n112 163.367
R605 B.n416 B.n415 163.367
R606 B.n417 B.n416 163.367
R607 B.n417 B.n110 163.367
R608 B.n421 B.n110 163.367
R609 B.n422 B.n421 163.367
R610 B.n423 B.n422 163.367
R611 B.n423 B.n108 163.367
R612 B.n427 B.n108 163.367
R613 B.n428 B.n427 163.367
R614 B.n429 B.n428 163.367
R615 B.n429 B.n106 163.367
R616 B.n433 B.n106 163.367
R617 B.n434 B.n433 163.367
R618 B.n435 B.n434 163.367
R619 B.n435 B.n104 163.367
R620 B.n439 B.n104 163.367
R621 B.n440 B.n439 163.367
R622 B.n441 B.n440 163.367
R623 B.n441 B.n102 163.367
R624 B.n445 B.n102 163.367
R625 B.n446 B.n445 163.367
R626 B.n447 B.n446 163.367
R627 B.n447 B.n100 163.367
R628 B.n451 B.n100 163.367
R629 B.n452 B.n451 163.367
R630 B.n453 B.n452 163.367
R631 B.n453 B.n98 163.367
R632 B.n457 B.n98 163.367
R633 B.n458 B.n457 163.367
R634 B.n459 B.n458 163.367
R635 B.n459 B.n96 163.367
R636 B.n463 B.n96 163.367
R637 B.n464 B.n463 163.367
R638 B.n465 B.n464 163.367
R639 B.n465 B.n94 163.367
R640 B.n469 B.n94 163.367
R641 B.n470 B.n469 163.367
R642 B.n471 B.n470 163.367
R643 B.n471 B.n92 163.367
R644 B.n475 B.n92 163.367
R645 B.n476 B.n475 163.367
R646 B.n477 B.n476 163.367
R647 B.n477 B.n90 163.367
R648 B.n481 B.n90 163.367
R649 B.n482 B.n481 163.367
R650 B.n483 B.n482 163.367
R651 B.n483 B.n88 163.367
R652 B.n487 B.n88 163.367
R653 B.n488 B.n487 163.367
R654 B.n489 B.n488 163.367
R655 B.n489 B.n86 163.367
R656 B.n493 B.n86 163.367
R657 B.n494 B.n493 163.367
R658 B.n495 B.n494 163.367
R659 B.n495 B.n84 163.367
R660 B.n499 B.n84 163.367
R661 B.n500 B.n499 163.367
R662 B.n501 B.n500 163.367
R663 B.n501 B.n82 163.367
R664 B.n505 B.n82 163.367
R665 B.n506 B.n505 163.367
R666 B.n507 B.n506 163.367
R667 B.n507 B.n80 163.367
R668 B.n511 B.n80 163.367
R669 B.n676 B.n19 163.367
R670 B.n676 B.n675 163.367
R671 B.n675 B.n674 163.367
R672 B.n674 B.n21 163.367
R673 B.n670 B.n21 163.367
R674 B.n670 B.n669 163.367
R675 B.n669 B.n668 163.367
R676 B.n668 B.n23 163.367
R677 B.n664 B.n23 163.367
R678 B.n664 B.n663 163.367
R679 B.n663 B.n662 163.367
R680 B.n662 B.n25 163.367
R681 B.n658 B.n25 163.367
R682 B.n658 B.n657 163.367
R683 B.n657 B.n656 163.367
R684 B.n656 B.n27 163.367
R685 B.n652 B.n27 163.367
R686 B.n652 B.n651 163.367
R687 B.n651 B.n650 163.367
R688 B.n650 B.n29 163.367
R689 B.n646 B.n29 163.367
R690 B.n646 B.n645 163.367
R691 B.n645 B.n644 163.367
R692 B.n644 B.n31 163.367
R693 B.n640 B.n31 163.367
R694 B.n640 B.n639 163.367
R695 B.n639 B.n638 163.367
R696 B.n638 B.n33 163.367
R697 B.n634 B.n33 163.367
R698 B.n634 B.n633 163.367
R699 B.n633 B.n632 163.367
R700 B.n632 B.n35 163.367
R701 B.n628 B.n35 163.367
R702 B.n628 B.n627 163.367
R703 B.n627 B.n626 163.367
R704 B.n626 B.n37 163.367
R705 B.n622 B.n37 163.367
R706 B.n622 B.n621 163.367
R707 B.n621 B.n620 163.367
R708 B.n620 B.n39 163.367
R709 B.n616 B.n39 163.367
R710 B.n616 B.n615 163.367
R711 B.n615 B.n614 163.367
R712 B.n614 B.n41 163.367
R713 B.n610 B.n41 163.367
R714 B.n610 B.n609 163.367
R715 B.n609 B.n608 163.367
R716 B.n608 B.n43 163.367
R717 B.n604 B.n43 163.367
R718 B.n604 B.n603 163.367
R719 B.n603 B.n602 163.367
R720 B.n602 B.n45 163.367
R721 B.n598 B.n45 163.367
R722 B.n598 B.n597 163.367
R723 B.n597 B.n596 163.367
R724 B.n596 B.n50 163.367
R725 B.n592 B.n50 163.367
R726 B.n592 B.n591 163.367
R727 B.n591 B.n590 163.367
R728 B.n590 B.n52 163.367
R729 B.n585 B.n52 163.367
R730 B.n585 B.n584 163.367
R731 B.n584 B.n583 163.367
R732 B.n583 B.n56 163.367
R733 B.n579 B.n56 163.367
R734 B.n579 B.n578 163.367
R735 B.n578 B.n577 163.367
R736 B.n577 B.n58 163.367
R737 B.n573 B.n58 163.367
R738 B.n573 B.n572 163.367
R739 B.n572 B.n571 163.367
R740 B.n571 B.n60 163.367
R741 B.n567 B.n60 163.367
R742 B.n567 B.n566 163.367
R743 B.n566 B.n565 163.367
R744 B.n565 B.n62 163.367
R745 B.n561 B.n62 163.367
R746 B.n561 B.n560 163.367
R747 B.n560 B.n559 163.367
R748 B.n559 B.n64 163.367
R749 B.n555 B.n64 163.367
R750 B.n555 B.n554 163.367
R751 B.n554 B.n553 163.367
R752 B.n553 B.n66 163.367
R753 B.n549 B.n66 163.367
R754 B.n549 B.n548 163.367
R755 B.n548 B.n547 163.367
R756 B.n547 B.n68 163.367
R757 B.n543 B.n68 163.367
R758 B.n543 B.n542 163.367
R759 B.n542 B.n541 163.367
R760 B.n541 B.n70 163.367
R761 B.n537 B.n70 163.367
R762 B.n537 B.n536 163.367
R763 B.n536 B.n535 163.367
R764 B.n535 B.n72 163.367
R765 B.n531 B.n72 163.367
R766 B.n531 B.n530 163.367
R767 B.n530 B.n529 163.367
R768 B.n529 B.n74 163.367
R769 B.n525 B.n74 163.367
R770 B.n525 B.n524 163.367
R771 B.n524 B.n523 163.367
R772 B.n523 B.n76 163.367
R773 B.n519 B.n76 163.367
R774 B.n519 B.n518 163.367
R775 B.n518 B.n517 163.367
R776 B.n517 B.n78 163.367
R777 B.n513 B.n78 163.367
R778 B.n513 B.n512 163.367
R779 B.n328 B.t7 109.07
R780 B.n54 B.t5 109.07
R781 B.n146 B.t1 109.05
R782 B.n47 B.t11 109.05
R783 B.n329 B.n328 59.5399
R784 B.n314 B.n146 59.5399
R785 B.n48 B.n47 59.5399
R786 B.n588 B.n54 59.5399
R787 B.n328 B.n327 57.2126
R788 B.n146 B.n145 57.2126
R789 B.n47 B.n46 57.2126
R790 B.n54 B.n53 57.2126
R791 B.n679 B.n678 33.8737
R792 B.n510 B.n79 33.8737
R793 B.n408 B.n407 33.8737
R794 B.n236 B.n171 33.8737
R795 B B.n731 18.0485
R796 B.n678 B.n677 10.6151
R797 B.n677 B.n20 10.6151
R798 B.n673 B.n20 10.6151
R799 B.n673 B.n672 10.6151
R800 B.n672 B.n671 10.6151
R801 B.n671 B.n22 10.6151
R802 B.n667 B.n22 10.6151
R803 B.n667 B.n666 10.6151
R804 B.n666 B.n665 10.6151
R805 B.n665 B.n24 10.6151
R806 B.n661 B.n24 10.6151
R807 B.n661 B.n660 10.6151
R808 B.n660 B.n659 10.6151
R809 B.n659 B.n26 10.6151
R810 B.n655 B.n26 10.6151
R811 B.n655 B.n654 10.6151
R812 B.n654 B.n653 10.6151
R813 B.n653 B.n28 10.6151
R814 B.n649 B.n28 10.6151
R815 B.n649 B.n648 10.6151
R816 B.n648 B.n647 10.6151
R817 B.n647 B.n30 10.6151
R818 B.n643 B.n30 10.6151
R819 B.n643 B.n642 10.6151
R820 B.n642 B.n641 10.6151
R821 B.n641 B.n32 10.6151
R822 B.n637 B.n32 10.6151
R823 B.n637 B.n636 10.6151
R824 B.n636 B.n635 10.6151
R825 B.n635 B.n34 10.6151
R826 B.n631 B.n34 10.6151
R827 B.n631 B.n630 10.6151
R828 B.n630 B.n629 10.6151
R829 B.n629 B.n36 10.6151
R830 B.n625 B.n36 10.6151
R831 B.n625 B.n624 10.6151
R832 B.n624 B.n623 10.6151
R833 B.n623 B.n38 10.6151
R834 B.n619 B.n38 10.6151
R835 B.n619 B.n618 10.6151
R836 B.n618 B.n617 10.6151
R837 B.n617 B.n40 10.6151
R838 B.n613 B.n40 10.6151
R839 B.n613 B.n612 10.6151
R840 B.n612 B.n611 10.6151
R841 B.n611 B.n42 10.6151
R842 B.n607 B.n42 10.6151
R843 B.n607 B.n606 10.6151
R844 B.n606 B.n605 10.6151
R845 B.n605 B.n44 10.6151
R846 B.n601 B.n600 10.6151
R847 B.n600 B.n599 10.6151
R848 B.n599 B.n49 10.6151
R849 B.n595 B.n49 10.6151
R850 B.n595 B.n594 10.6151
R851 B.n594 B.n593 10.6151
R852 B.n593 B.n51 10.6151
R853 B.n589 B.n51 10.6151
R854 B.n587 B.n586 10.6151
R855 B.n586 B.n55 10.6151
R856 B.n582 B.n55 10.6151
R857 B.n582 B.n581 10.6151
R858 B.n581 B.n580 10.6151
R859 B.n580 B.n57 10.6151
R860 B.n576 B.n57 10.6151
R861 B.n576 B.n575 10.6151
R862 B.n575 B.n574 10.6151
R863 B.n574 B.n59 10.6151
R864 B.n570 B.n59 10.6151
R865 B.n570 B.n569 10.6151
R866 B.n569 B.n568 10.6151
R867 B.n568 B.n61 10.6151
R868 B.n564 B.n61 10.6151
R869 B.n564 B.n563 10.6151
R870 B.n563 B.n562 10.6151
R871 B.n562 B.n63 10.6151
R872 B.n558 B.n63 10.6151
R873 B.n558 B.n557 10.6151
R874 B.n557 B.n556 10.6151
R875 B.n556 B.n65 10.6151
R876 B.n552 B.n65 10.6151
R877 B.n552 B.n551 10.6151
R878 B.n551 B.n550 10.6151
R879 B.n550 B.n67 10.6151
R880 B.n546 B.n67 10.6151
R881 B.n546 B.n545 10.6151
R882 B.n545 B.n544 10.6151
R883 B.n544 B.n69 10.6151
R884 B.n540 B.n69 10.6151
R885 B.n540 B.n539 10.6151
R886 B.n539 B.n538 10.6151
R887 B.n538 B.n71 10.6151
R888 B.n534 B.n71 10.6151
R889 B.n534 B.n533 10.6151
R890 B.n533 B.n532 10.6151
R891 B.n532 B.n73 10.6151
R892 B.n528 B.n73 10.6151
R893 B.n528 B.n527 10.6151
R894 B.n527 B.n526 10.6151
R895 B.n526 B.n75 10.6151
R896 B.n522 B.n75 10.6151
R897 B.n522 B.n521 10.6151
R898 B.n521 B.n520 10.6151
R899 B.n520 B.n77 10.6151
R900 B.n516 B.n77 10.6151
R901 B.n516 B.n515 10.6151
R902 B.n515 B.n514 10.6151
R903 B.n514 B.n79 10.6151
R904 B.n408 B.n113 10.6151
R905 B.n412 B.n113 10.6151
R906 B.n413 B.n412 10.6151
R907 B.n414 B.n413 10.6151
R908 B.n414 B.n111 10.6151
R909 B.n418 B.n111 10.6151
R910 B.n419 B.n418 10.6151
R911 B.n420 B.n419 10.6151
R912 B.n420 B.n109 10.6151
R913 B.n424 B.n109 10.6151
R914 B.n425 B.n424 10.6151
R915 B.n426 B.n425 10.6151
R916 B.n426 B.n107 10.6151
R917 B.n430 B.n107 10.6151
R918 B.n431 B.n430 10.6151
R919 B.n432 B.n431 10.6151
R920 B.n432 B.n105 10.6151
R921 B.n436 B.n105 10.6151
R922 B.n437 B.n436 10.6151
R923 B.n438 B.n437 10.6151
R924 B.n438 B.n103 10.6151
R925 B.n442 B.n103 10.6151
R926 B.n443 B.n442 10.6151
R927 B.n444 B.n443 10.6151
R928 B.n444 B.n101 10.6151
R929 B.n448 B.n101 10.6151
R930 B.n449 B.n448 10.6151
R931 B.n450 B.n449 10.6151
R932 B.n450 B.n99 10.6151
R933 B.n454 B.n99 10.6151
R934 B.n455 B.n454 10.6151
R935 B.n456 B.n455 10.6151
R936 B.n456 B.n97 10.6151
R937 B.n460 B.n97 10.6151
R938 B.n461 B.n460 10.6151
R939 B.n462 B.n461 10.6151
R940 B.n462 B.n95 10.6151
R941 B.n466 B.n95 10.6151
R942 B.n467 B.n466 10.6151
R943 B.n468 B.n467 10.6151
R944 B.n468 B.n93 10.6151
R945 B.n472 B.n93 10.6151
R946 B.n473 B.n472 10.6151
R947 B.n474 B.n473 10.6151
R948 B.n474 B.n91 10.6151
R949 B.n478 B.n91 10.6151
R950 B.n479 B.n478 10.6151
R951 B.n480 B.n479 10.6151
R952 B.n480 B.n89 10.6151
R953 B.n484 B.n89 10.6151
R954 B.n485 B.n484 10.6151
R955 B.n486 B.n485 10.6151
R956 B.n486 B.n87 10.6151
R957 B.n490 B.n87 10.6151
R958 B.n491 B.n490 10.6151
R959 B.n492 B.n491 10.6151
R960 B.n492 B.n85 10.6151
R961 B.n496 B.n85 10.6151
R962 B.n497 B.n496 10.6151
R963 B.n498 B.n497 10.6151
R964 B.n498 B.n83 10.6151
R965 B.n502 B.n83 10.6151
R966 B.n503 B.n502 10.6151
R967 B.n504 B.n503 10.6151
R968 B.n504 B.n81 10.6151
R969 B.n508 B.n81 10.6151
R970 B.n509 B.n508 10.6151
R971 B.n510 B.n509 10.6151
R972 B.n240 B.n171 10.6151
R973 B.n241 B.n240 10.6151
R974 B.n242 B.n241 10.6151
R975 B.n242 B.n169 10.6151
R976 B.n246 B.n169 10.6151
R977 B.n247 B.n246 10.6151
R978 B.n248 B.n247 10.6151
R979 B.n248 B.n167 10.6151
R980 B.n252 B.n167 10.6151
R981 B.n253 B.n252 10.6151
R982 B.n254 B.n253 10.6151
R983 B.n254 B.n165 10.6151
R984 B.n258 B.n165 10.6151
R985 B.n259 B.n258 10.6151
R986 B.n260 B.n259 10.6151
R987 B.n260 B.n163 10.6151
R988 B.n264 B.n163 10.6151
R989 B.n265 B.n264 10.6151
R990 B.n266 B.n265 10.6151
R991 B.n266 B.n161 10.6151
R992 B.n270 B.n161 10.6151
R993 B.n271 B.n270 10.6151
R994 B.n272 B.n271 10.6151
R995 B.n272 B.n159 10.6151
R996 B.n276 B.n159 10.6151
R997 B.n277 B.n276 10.6151
R998 B.n278 B.n277 10.6151
R999 B.n278 B.n157 10.6151
R1000 B.n282 B.n157 10.6151
R1001 B.n283 B.n282 10.6151
R1002 B.n284 B.n283 10.6151
R1003 B.n284 B.n155 10.6151
R1004 B.n288 B.n155 10.6151
R1005 B.n289 B.n288 10.6151
R1006 B.n290 B.n289 10.6151
R1007 B.n290 B.n153 10.6151
R1008 B.n294 B.n153 10.6151
R1009 B.n295 B.n294 10.6151
R1010 B.n296 B.n295 10.6151
R1011 B.n296 B.n151 10.6151
R1012 B.n300 B.n151 10.6151
R1013 B.n301 B.n300 10.6151
R1014 B.n302 B.n301 10.6151
R1015 B.n302 B.n149 10.6151
R1016 B.n306 B.n149 10.6151
R1017 B.n307 B.n306 10.6151
R1018 B.n308 B.n307 10.6151
R1019 B.n308 B.n147 10.6151
R1020 B.n312 B.n147 10.6151
R1021 B.n313 B.n312 10.6151
R1022 B.n315 B.n143 10.6151
R1023 B.n319 B.n143 10.6151
R1024 B.n320 B.n319 10.6151
R1025 B.n321 B.n320 10.6151
R1026 B.n321 B.n141 10.6151
R1027 B.n325 B.n141 10.6151
R1028 B.n326 B.n325 10.6151
R1029 B.n330 B.n326 10.6151
R1030 B.n334 B.n139 10.6151
R1031 B.n335 B.n334 10.6151
R1032 B.n336 B.n335 10.6151
R1033 B.n336 B.n137 10.6151
R1034 B.n340 B.n137 10.6151
R1035 B.n341 B.n340 10.6151
R1036 B.n342 B.n341 10.6151
R1037 B.n342 B.n135 10.6151
R1038 B.n346 B.n135 10.6151
R1039 B.n347 B.n346 10.6151
R1040 B.n348 B.n347 10.6151
R1041 B.n348 B.n133 10.6151
R1042 B.n352 B.n133 10.6151
R1043 B.n353 B.n352 10.6151
R1044 B.n354 B.n353 10.6151
R1045 B.n354 B.n131 10.6151
R1046 B.n358 B.n131 10.6151
R1047 B.n359 B.n358 10.6151
R1048 B.n360 B.n359 10.6151
R1049 B.n360 B.n129 10.6151
R1050 B.n364 B.n129 10.6151
R1051 B.n365 B.n364 10.6151
R1052 B.n366 B.n365 10.6151
R1053 B.n366 B.n127 10.6151
R1054 B.n370 B.n127 10.6151
R1055 B.n371 B.n370 10.6151
R1056 B.n372 B.n371 10.6151
R1057 B.n372 B.n125 10.6151
R1058 B.n376 B.n125 10.6151
R1059 B.n377 B.n376 10.6151
R1060 B.n378 B.n377 10.6151
R1061 B.n378 B.n123 10.6151
R1062 B.n382 B.n123 10.6151
R1063 B.n383 B.n382 10.6151
R1064 B.n384 B.n383 10.6151
R1065 B.n384 B.n121 10.6151
R1066 B.n388 B.n121 10.6151
R1067 B.n389 B.n388 10.6151
R1068 B.n390 B.n389 10.6151
R1069 B.n390 B.n119 10.6151
R1070 B.n394 B.n119 10.6151
R1071 B.n395 B.n394 10.6151
R1072 B.n396 B.n395 10.6151
R1073 B.n396 B.n117 10.6151
R1074 B.n400 B.n117 10.6151
R1075 B.n401 B.n400 10.6151
R1076 B.n402 B.n401 10.6151
R1077 B.n402 B.n115 10.6151
R1078 B.n406 B.n115 10.6151
R1079 B.n407 B.n406 10.6151
R1080 B.n236 B.n235 10.6151
R1081 B.n235 B.n234 10.6151
R1082 B.n234 B.n173 10.6151
R1083 B.n230 B.n173 10.6151
R1084 B.n230 B.n229 10.6151
R1085 B.n229 B.n228 10.6151
R1086 B.n228 B.n175 10.6151
R1087 B.n224 B.n175 10.6151
R1088 B.n224 B.n223 10.6151
R1089 B.n223 B.n222 10.6151
R1090 B.n222 B.n177 10.6151
R1091 B.n218 B.n177 10.6151
R1092 B.n218 B.n217 10.6151
R1093 B.n217 B.n216 10.6151
R1094 B.n216 B.n179 10.6151
R1095 B.n212 B.n179 10.6151
R1096 B.n212 B.n211 10.6151
R1097 B.n211 B.n210 10.6151
R1098 B.n210 B.n181 10.6151
R1099 B.n206 B.n181 10.6151
R1100 B.n206 B.n205 10.6151
R1101 B.n205 B.n204 10.6151
R1102 B.n204 B.n183 10.6151
R1103 B.n200 B.n183 10.6151
R1104 B.n200 B.n199 10.6151
R1105 B.n199 B.n198 10.6151
R1106 B.n198 B.n185 10.6151
R1107 B.n194 B.n185 10.6151
R1108 B.n194 B.n193 10.6151
R1109 B.n193 B.n192 10.6151
R1110 B.n192 B.n187 10.6151
R1111 B.n188 B.n187 10.6151
R1112 B.n188 B.n0 10.6151
R1113 B.n727 B.n1 10.6151
R1114 B.n727 B.n726 10.6151
R1115 B.n726 B.n725 10.6151
R1116 B.n725 B.n4 10.6151
R1117 B.n721 B.n4 10.6151
R1118 B.n721 B.n720 10.6151
R1119 B.n720 B.n719 10.6151
R1120 B.n719 B.n6 10.6151
R1121 B.n715 B.n6 10.6151
R1122 B.n715 B.n714 10.6151
R1123 B.n714 B.n713 10.6151
R1124 B.n713 B.n8 10.6151
R1125 B.n709 B.n8 10.6151
R1126 B.n709 B.n708 10.6151
R1127 B.n708 B.n707 10.6151
R1128 B.n707 B.n10 10.6151
R1129 B.n703 B.n10 10.6151
R1130 B.n703 B.n702 10.6151
R1131 B.n702 B.n701 10.6151
R1132 B.n701 B.n12 10.6151
R1133 B.n697 B.n12 10.6151
R1134 B.n697 B.n696 10.6151
R1135 B.n696 B.n695 10.6151
R1136 B.n695 B.n14 10.6151
R1137 B.n691 B.n14 10.6151
R1138 B.n691 B.n690 10.6151
R1139 B.n690 B.n689 10.6151
R1140 B.n689 B.n16 10.6151
R1141 B.n685 B.n16 10.6151
R1142 B.n685 B.n684 10.6151
R1143 B.n684 B.n683 10.6151
R1144 B.n683 B.n18 10.6151
R1145 B.n679 B.n18 10.6151
R1146 B.n601 B.n48 6.5566
R1147 B.n589 B.n588 6.5566
R1148 B.n315 B.n314 6.5566
R1149 B.n330 B.n329 6.5566
R1150 B.n48 B.n44 4.05904
R1151 B.n588 B.n587 4.05904
R1152 B.n314 B.n313 4.05904
R1153 B.n329 B.n139 4.05904
R1154 B.n731 B.n0 2.81026
R1155 B.n731 B.n1 2.81026
R1156 VN.n0 VN.t2 175.141
R1157 VN.n1 VN.t1 175.141
R1158 VN.n0 VN.t0 174.363
R1159 VN.n1 VN.t3 174.363
R1160 VN VN.n1 53.3191
R1161 VN VN.n0 4.29263
R1162 VDD2.n2 VDD2.n0 116.603
R1163 VDD2.n2 VDD2.n1 72.2504
R1164 VDD2.n1 VDD2.t0 2.15458
R1165 VDD2.n1 VDD2.t2 2.15458
R1166 VDD2.n0 VDD2.t1 2.15458
R1167 VDD2.n0 VDD2.t3 2.15458
R1168 VDD2 VDD2.n2 0.0586897
C0 B VDD2 1.40007f
C1 VDD2 w_n2740_n3986# 1.59924f
C2 B VP 1.73343f
C3 VP w_n2740_n3986# 5.04615f
C4 VN VTAIL 5.67472f
C5 VN VDD1 0.149154f
C6 VTAIL VDD1 6.14331f
C7 B w_n2740_n3986# 10.1373f
C8 VN VDD2 5.89746f
C9 VDD2 VTAIL 6.19766f
C10 VDD2 VDD1 1.02554f
C11 VN VP 6.77523f
C12 VP VTAIL 5.68883f
C13 VP VDD1 6.14328f
C14 VN B 1.14873f
C15 VN w_n2740_n3986# 4.69386f
C16 B VTAIL 5.97096f
C17 VP VDD2 0.395714f
C18 VTAIL w_n2740_n3986# 4.66956f
C19 B VDD1 1.3476f
C20 w_n2740_n3986# VDD1 1.54268f
C21 VDD2 VSUBS 1.031147f
C22 VDD1 VSUBS 6.1009f
C23 VTAIL VSUBS 1.362166f
C24 VN VSUBS 5.5731f
C25 VP VSUBS 2.407638f
C26 B VSUBS 4.55539f
C27 w_n2740_n3986# VSUBS 0.13392p
C28 VDD2.t1 VSUBS 0.317689f
C29 VDD2.t3 VSUBS 0.317689f
C30 VDD2.n0 VSUBS 3.40592f
C31 VDD2.t0 VSUBS 0.317689f
C32 VDD2.t2 VSUBS 0.317689f
C33 VDD2.n1 VSUBS 2.58659f
C34 VDD2.n2 VSUBS 4.61269f
C35 VN.t2 VSUBS 3.63888f
C36 VN.t0 VSUBS 3.63293f
C37 VN.n0 VSUBS 2.31528f
C38 VN.t1 VSUBS 3.63888f
C39 VN.t3 VSUBS 3.63293f
C40 VN.n1 VSUBS 4.10975f
C41 B.n0 VSUBS 0.003986f
C42 B.n1 VSUBS 0.003986f
C43 B.n2 VSUBS 0.006304f
C44 B.n3 VSUBS 0.006304f
C45 B.n4 VSUBS 0.006304f
C46 B.n5 VSUBS 0.006304f
C47 B.n6 VSUBS 0.006304f
C48 B.n7 VSUBS 0.006304f
C49 B.n8 VSUBS 0.006304f
C50 B.n9 VSUBS 0.006304f
C51 B.n10 VSUBS 0.006304f
C52 B.n11 VSUBS 0.006304f
C53 B.n12 VSUBS 0.006304f
C54 B.n13 VSUBS 0.006304f
C55 B.n14 VSUBS 0.006304f
C56 B.n15 VSUBS 0.006304f
C57 B.n16 VSUBS 0.006304f
C58 B.n17 VSUBS 0.006304f
C59 B.n18 VSUBS 0.006304f
C60 B.n19 VSUBS 0.01554f
C61 B.n20 VSUBS 0.006304f
C62 B.n21 VSUBS 0.006304f
C63 B.n22 VSUBS 0.006304f
C64 B.n23 VSUBS 0.006304f
C65 B.n24 VSUBS 0.006304f
C66 B.n25 VSUBS 0.006304f
C67 B.n26 VSUBS 0.006304f
C68 B.n27 VSUBS 0.006304f
C69 B.n28 VSUBS 0.006304f
C70 B.n29 VSUBS 0.006304f
C71 B.n30 VSUBS 0.006304f
C72 B.n31 VSUBS 0.006304f
C73 B.n32 VSUBS 0.006304f
C74 B.n33 VSUBS 0.006304f
C75 B.n34 VSUBS 0.006304f
C76 B.n35 VSUBS 0.006304f
C77 B.n36 VSUBS 0.006304f
C78 B.n37 VSUBS 0.006304f
C79 B.n38 VSUBS 0.006304f
C80 B.n39 VSUBS 0.006304f
C81 B.n40 VSUBS 0.006304f
C82 B.n41 VSUBS 0.006304f
C83 B.n42 VSUBS 0.006304f
C84 B.n43 VSUBS 0.006304f
C85 B.n44 VSUBS 0.004357f
C86 B.n45 VSUBS 0.006304f
C87 B.t11 VSUBS 0.452607f
C88 B.t10 VSUBS 0.471846f
C89 B.t9 VSUBS 1.59897f
C90 B.n46 VSUBS 0.252483f
C91 B.n47 VSUBS 0.0649f
C92 B.n48 VSUBS 0.014605f
C93 B.n49 VSUBS 0.006304f
C94 B.n50 VSUBS 0.006304f
C95 B.n51 VSUBS 0.006304f
C96 B.n52 VSUBS 0.006304f
C97 B.t5 VSUBS 0.452594f
C98 B.t4 VSUBS 0.471835f
C99 B.t3 VSUBS 1.59897f
C100 B.n53 VSUBS 0.252494f
C101 B.n54 VSUBS 0.064913f
C102 B.n55 VSUBS 0.006304f
C103 B.n56 VSUBS 0.006304f
C104 B.n57 VSUBS 0.006304f
C105 B.n58 VSUBS 0.006304f
C106 B.n59 VSUBS 0.006304f
C107 B.n60 VSUBS 0.006304f
C108 B.n61 VSUBS 0.006304f
C109 B.n62 VSUBS 0.006304f
C110 B.n63 VSUBS 0.006304f
C111 B.n64 VSUBS 0.006304f
C112 B.n65 VSUBS 0.006304f
C113 B.n66 VSUBS 0.006304f
C114 B.n67 VSUBS 0.006304f
C115 B.n68 VSUBS 0.006304f
C116 B.n69 VSUBS 0.006304f
C117 B.n70 VSUBS 0.006304f
C118 B.n71 VSUBS 0.006304f
C119 B.n72 VSUBS 0.006304f
C120 B.n73 VSUBS 0.006304f
C121 B.n74 VSUBS 0.006304f
C122 B.n75 VSUBS 0.006304f
C123 B.n76 VSUBS 0.006304f
C124 B.n77 VSUBS 0.006304f
C125 B.n78 VSUBS 0.006304f
C126 B.n79 VSUBS 0.014822f
C127 B.n80 VSUBS 0.006304f
C128 B.n81 VSUBS 0.006304f
C129 B.n82 VSUBS 0.006304f
C130 B.n83 VSUBS 0.006304f
C131 B.n84 VSUBS 0.006304f
C132 B.n85 VSUBS 0.006304f
C133 B.n86 VSUBS 0.006304f
C134 B.n87 VSUBS 0.006304f
C135 B.n88 VSUBS 0.006304f
C136 B.n89 VSUBS 0.006304f
C137 B.n90 VSUBS 0.006304f
C138 B.n91 VSUBS 0.006304f
C139 B.n92 VSUBS 0.006304f
C140 B.n93 VSUBS 0.006304f
C141 B.n94 VSUBS 0.006304f
C142 B.n95 VSUBS 0.006304f
C143 B.n96 VSUBS 0.006304f
C144 B.n97 VSUBS 0.006304f
C145 B.n98 VSUBS 0.006304f
C146 B.n99 VSUBS 0.006304f
C147 B.n100 VSUBS 0.006304f
C148 B.n101 VSUBS 0.006304f
C149 B.n102 VSUBS 0.006304f
C150 B.n103 VSUBS 0.006304f
C151 B.n104 VSUBS 0.006304f
C152 B.n105 VSUBS 0.006304f
C153 B.n106 VSUBS 0.006304f
C154 B.n107 VSUBS 0.006304f
C155 B.n108 VSUBS 0.006304f
C156 B.n109 VSUBS 0.006304f
C157 B.n110 VSUBS 0.006304f
C158 B.n111 VSUBS 0.006304f
C159 B.n112 VSUBS 0.006304f
C160 B.n113 VSUBS 0.006304f
C161 B.n114 VSUBS 0.01554f
C162 B.n115 VSUBS 0.006304f
C163 B.n116 VSUBS 0.006304f
C164 B.n117 VSUBS 0.006304f
C165 B.n118 VSUBS 0.006304f
C166 B.n119 VSUBS 0.006304f
C167 B.n120 VSUBS 0.006304f
C168 B.n121 VSUBS 0.006304f
C169 B.n122 VSUBS 0.006304f
C170 B.n123 VSUBS 0.006304f
C171 B.n124 VSUBS 0.006304f
C172 B.n125 VSUBS 0.006304f
C173 B.n126 VSUBS 0.006304f
C174 B.n127 VSUBS 0.006304f
C175 B.n128 VSUBS 0.006304f
C176 B.n129 VSUBS 0.006304f
C177 B.n130 VSUBS 0.006304f
C178 B.n131 VSUBS 0.006304f
C179 B.n132 VSUBS 0.006304f
C180 B.n133 VSUBS 0.006304f
C181 B.n134 VSUBS 0.006304f
C182 B.n135 VSUBS 0.006304f
C183 B.n136 VSUBS 0.006304f
C184 B.n137 VSUBS 0.006304f
C185 B.n138 VSUBS 0.006304f
C186 B.n139 VSUBS 0.004357f
C187 B.n140 VSUBS 0.006304f
C188 B.n141 VSUBS 0.006304f
C189 B.n142 VSUBS 0.006304f
C190 B.n143 VSUBS 0.006304f
C191 B.n144 VSUBS 0.006304f
C192 B.t1 VSUBS 0.452607f
C193 B.t2 VSUBS 0.471846f
C194 B.t0 VSUBS 1.59897f
C195 B.n145 VSUBS 0.252483f
C196 B.n146 VSUBS 0.0649f
C197 B.n147 VSUBS 0.006304f
C198 B.n148 VSUBS 0.006304f
C199 B.n149 VSUBS 0.006304f
C200 B.n150 VSUBS 0.006304f
C201 B.n151 VSUBS 0.006304f
C202 B.n152 VSUBS 0.006304f
C203 B.n153 VSUBS 0.006304f
C204 B.n154 VSUBS 0.006304f
C205 B.n155 VSUBS 0.006304f
C206 B.n156 VSUBS 0.006304f
C207 B.n157 VSUBS 0.006304f
C208 B.n158 VSUBS 0.006304f
C209 B.n159 VSUBS 0.006304f
C210 B.n160 VSUBS 0.006304f
C211 B.n161 VSUBS 0.006304f
C212 B.n162 VSUBS 0.006304f
C213 B.n163 VSUBS 0.006304f
C214 B.n164 VSUBS 0.006304f
C215 B.n165 VSUBS 0.006304f
C216 B.n166 VSUBS 0.006304f
C217 B.n167 VSUBS 0.006304f
C218 B.n168 VSUBS 0.006304f
C219 B.n169 VSUBS 0.006304f
C220 B.n170 VSUBS 0.006304f
C221 B.n171 VSUBS 0.01554f
C222 B.n172 VSUBS 0.006304f
C223 B.n173 VSUBS 0.006304f
C224 B.n174 VSUBS 0.006304f
C225 B.n175 VSUBS 0.006304f
C226 B.n176 VSUBS 0.006304f
C227 B.n177 VSUBS 0.006304f
C228 B.n178 VSUBS 0.006304f
C229 B.n179 VSUBS 0.006304f
C230 B.n180 VSUBS 0.006304f
C231 B.n181 VSUBS 0.006304f
C232 B.n182 VSUBS 0.006304f
C233 B.n183 VSUBS 0.006304f
C234 B.n184 VSUBS 0.006304f
C235 B.n185 VSUBS 0.006304f
C236 B.n186 VSUBS 0.006304f
C237 B.n187 VSUBS 0.006304f
C238 B.n188 VSUBS 0.006304f
C239 B.n189 VSUBS 0.006304f
C240 B.n190 VSUBS 0.006304f
C241 B.n191 VSUBS 0.006304f
C242 B.n192 VSUBS 0.006304f
C243 B.n193 VSUBS 0.006304f
C244 B.n194 VSUBS 0.006304f
C245 B.n195 VSUBS 0.006304f
C246 B.n196 VSUBS 0.006304f
C247 B.n197 VSUBS 0.006304f
C248 B.n198 VSUBS 0.006304f
C249 B.n199 VSUBS 0.006304f
C250 B.n200 VSUBS 0.006304f
C251 B.n201 VSUBS 0.006304f
C252 B.n202 VSUBS 0.006304f
C253 B.n203 VSUBS 0.006304f
C254 B.n204 VSUBS 0.006304f
C255 B.n205 VSUBS 0.006304f
C256 B.n206 VSUBS 0.006304f
C257 B.n207 VSUBS 0.006304f
C258 B.n208 VSUBS 0.006304f
C259 B.n209 VSUBS 0.006304f
C260 B.n210 VSUBS 0.006304f
C261 B.n211 VSUBS 0.006304f
C262 B.n212 VSUBS 0.006304f
C263 B.n213 VSUBS 0.006304f
C264 B.n214 VSUBS 0.006304f
C265 B.n215 VSUBS 0.006304f
C266 B.n216 VSUBS 0.006304f
C267 B.n217 VSUBS 0.006304f
C268 B.n218 VSUBS 0.006304f
C269 B.n219 VSUBS 0.006304f
C270 B.n220 VSUBS 0.006304f
C271 B.n221 VSUBS 0.006304f
C272 B.n222 VSUBS 0.006304f
C273 B.n223 VSUBS 0.006304f
C274 B.n224 VSUBS 0.006304f
C275 B.n225 VSUBS 0.006304f
C276 B.n226 VSUBS 0.006304f
C277 B.n227 VSUBS 0.006304f
C278 B.n228 VSUBS 0.006304f
C279 B.n229 VSUBS 0.006304f
C280 B.n230 VSUBS 0.006304f
C281 B.n231 VSUBS 0.006304f
C282 B.n232 VSUBS 0.006304f
C283 B.n233 VSUBS 0.006304f
C284 B.n234 VSUBS 0.006304f
C285 B.n235 VSUBS 0.006304f
C286 B.n236 VSUBS 0.014681f
C287 B.n237 VSUBS 0.014681f
C288 B.n238 VSUBS 0.01554f
C289 B.n239 VSUBS 0.006304f
C290 B.n240 VSUBS 0.006304f
C291 B.n241 VSUBS 0.006304f
C292 B.n242 VSUBS 0.006304f
C293 B.n243 VSUBS 0.006304f
C294 B.n244 VSUBS 0.006304f
C295 B.n245 VSUBS 0.006304f
C296 B.n246 VSUBS 0.006304f
C297 B.n247 VSUBS 0.006304f
C298 B.n248 VSUBS 0.006304f
C299 B.n249 VSUBS 0.006304f
C300 B.n250 VSUBS 0.006304f
C301 B.n251 VSUBS 0.006304f
C302 B.n252 VSUBS 0.006304f
C303 B.n253 VSUBS 0.006304f
C304 B.n254 VSUBS 0.006304f
C305 B.n255 VSUBS 0.006304f
C306 B.n256 VSUBS 0.006304f
C307 B.n257 VSUBS 0.006304f
C308 B.n258 VSUBS 0.006304f
C309 B.n259 VSUBS 0.006304f
C310 B.n260 VSUBS 0.006304f
C311 B.n261 VSUBS 0.006304f
C312 B.n262 VSUBS 0.006304f
C313 B.n263 VSUBS 0.006304f
C314 B.n264 VSUBS 0.006304f
C315 B.n265 VSUBS 0.006304f
C316 B.n266 VSUBS 0.006304f
C317 B.n267 VSUBS 0.006304f
C318 B.n268 VSUBS 0.006304f
C319 B.n269 VSUBS 0.006304f
C320 B.n270 VSUBS 0.006304f
C321 B.n271 VSUBS 0.006304f
C322 B.n272 VSUBS 0.006304f
C323 B.n273 VSUBS 0.006304f
C324 B.n274 VSUBS 0.006304f
C325 B.n275 VSUBS 0.006304f
C326 B.n276 VSUBS 0.006304f
C327 B.n277 VSUBS 0.006304f
C328 B.n278 VSUBS 0.006304f
C329 B.n279 VSUBS 0.006304f
C330 B.n280 VSUBS 0.006304f
C331 B.n281 VSUBS 0.006304f
C332 B.n282 VSUBS 0.006304f
C333 B.n283 VSUBS 0.006304f
C334 B.n284 VSUBS 0.006304f
C335 B.n285 VSUBS 0.006304f
C336 B.n286 VSUBS 0.006304f
C337 B.n287 VSUBS 0.006304f
C338 B.n288 VSUBS 0.006304f
C339 B.n289 VSUBS 0.006304f
C340 B.n290 VSUBS 0.006304f
C341 B.n291 VSUBS 0.006304f
C342 B.n292 VSUBS 0.006304f
C343 B.n293 VSUBS 0.006304f
C344 B.n294 VSUBS 0.006304f
C345 B.n295 VSUBS 0.006304f
C346 B.n296 VSUBS 0.006304f
C347 B.n297 VSUBS 0.006304f
C348 B.n298 VSUBS 0.006304f
C349 B.n299 VSUBS 0.006304f
C350 B.n300 VSUBS 0.006304f
C351 B.n301 VSUBS 0.006304f
C352 B.n302 VSUBS 0.006304f
C353 B.n303 VSUBS 0.006304f
C354 B.n304 VSUBS 0.006304f
C355 B.n305 VSUBS 0.006304f
C356 B.n306 VSUBS 0.006304f
C357 B.n307 VSUBS 0.006304f
C358 B.n308 VSUBS 0.006304f
C359 B.n309 VSUBS 0.006304f
C360 B.n310 VSUBS 0.006304f
C361 B.n311 VSUBS 0.006304f
C362 B.n312 VSUBS 0.006304f
C363 B.n313 VSUBS 0.004357f
C364 B.n314 VSUBS 0.014605f
C365 B.n315 VSUBS 0.005099f
C366 B.n316 VSUBS 0.006304f
C367 B.n317 VSUBS 0.006304f
C368 B.n318 VSUBS 0.006304f
C369 B.n319 VSUBS 0.006304f
C370 B.n320 VSUBS 0.006304f
C371 B.n321 VSUBS 0.006304f
C372 B.n322 VSUBS 0.006304f
C373 B.n323 VSUBS 0.006304f
C374 B.n324 VSUBS 0.006304f
C375 B.n325 VSUBS 0.006304f
C376 B.n326 VSUBS 0.006304f
C377 B.t7 VSUBS 0.452594f
C378 B.t8 VSUBS 0.471835f
C379 B.t6 VSUBS 1.59897f
C380 B.n327 VSUBS 0.252494f
C381 B.n328 VSUBS 0.064913f
C382 B.n329 VSUBS 0.014605f
C383 B.n330 VSUBS 0.005099f
C384 B.n331 VSUBS 0.006304f
C385 B.n332 VSUBS 0.006304f
C386 B.n333 VSUBS 0.006304f
C387 B.n334 VSUBS 0.006304f
C388 B.n335 VSUBS 0.006304f
C389 B.n336 VSUBS 0.006304f
C390 B.n337 VSUBS 0.006304f
C391 B.n338 VSUBS 0.006304f
C392 B.n339 VSUBS 0.006304f
C393 B.n340 VSUBS 0.006304f
C394 B.n341 VSUBS 0.006304f
C395 B.n342 VSUBS 0.006304f
C396 B.n343 VSUBS 0.006304f
C397 B.n344 VSUBS 0.006304f
C398 B.n345 VSUBS 0.006304f
C399 B.n346 VSUBS 0.006304f
C400 B.n347 VSUBS 0.006304f
C401 B.n348 VSUBS 0.006304f
C402 B.n349 VSUBS 0.006304f
C403 B.n350 VSUBS 0.006304f
C404 B.n351 VSUBS 0.006304f
C405 B.n352 VSUBS 0.006304f
C406 B.n353 VSUBS 0.006304f
C407 B.n354 VSUBS 0.006304f
C408 B.n355 VSUBS 0.006304f
C409 B.n356 VSUBS 0.006304f
C410 B.n357 VSUBS 0.006304f
C411 B.n358 VSUBS 0.006304f
C412 B.n359 VSUBS 0.006304f
C413 B.n360 VSUBS 0.006304f
C414 B.n361 VSUBS 0.006304f
C415 B.n362 VSUBS 0.006304f
C416 B.n363 VSUBS 0.006304f
C417 B.n364 VSUBS 0.006304f
C418 B.n365 VSUBS 0.006304f
C419 B.n366 VSUBS 0.006304f
C420 B.n367 VSUBS 0.006304f
C421 B.n368 VSUBS 0.006304f
C422 B.n369 VSUBS 0.006304f
C423 B.n370 VSUBS 0.006304f
C424 B.n371 VSUBS 0.006304f
C425 B.n372 VSUBS 0.006304f
C426 B.n373 VSUBS 0.006304f
C427 B.n374 VSUBS 0.006304f
C428 B.n375 VSUBS 0.006304f
C429 B.n376 VSUBS 0.006304f
C430 B.n377 VSUBS 0.006304f
C431 B.n378 VSUBS 0.006304f
C432 B.n379 VSUBS 0.006304f
C433 B.n380 VSUBS 0.006304f
C434 B.n381 VSUBS 0.006304f
C435 B.n382 VSUBS 0.006304f
C436 B.n383 VSUBS 0.006304f
C437 B.n384 VSUBS 0.006304f
C438 B.n385 VSUBS 0.006304f
C439 B.n386 VSUBS 0.006304f
C440 B.n387 VSUBS 0.006304f
C441 B.n388 VSUBS 0.006304f
C442 B.n389 VSUBS 0.006304f
C443 B.n390 VSUBS 0.006304f
C444 B.n391 VSUBS 0.006304f
C445 B.n392 VSUBS 0.006304f
C446 B.n393 VSUBS 0.006304f
C447 B.n394 VSUBS 0.006304f
C448 B.n395 VSUBS 0.006304f
C449 B.n396 VSUBS 0.006304f
C450 B.n397 VSUBS 0.006304f
C451 B.n398 VSUBS 0.006304f
C452 B.n399 VSUBS 0.006304f
C453 B.n400 VSUBS 0.006304f
C454 B.n401 VSUBS 0.006304f
C455 B.n402 VSUBS 0.006304f
C456 B.n403 VSUBS 0.006304f
C457 B.n404 VSUBS 0.006304f
C458 B.n405 VSUBS 0.006304f
C459 B.n406 VSUBS 0.006304f
C460 B.n407 VSUBS 0.01554f
C461 B.n408 VSUBS 0.014681f
C462 B.n409 VSUBS 0.014681f
C463 B.n410 VSUBS 0.006304f
C464 B.n411 VSUBS 0.006304f
C465 B.n412 VSUBS 0.006304f
C466 B.n413 VSUBS 0.006304f
C467 B.n414 VSUBS 0.006304f
C468 B.n415 VSUBS 0.006304f
C469 B.n416 VSUBS 0.006304f
C470 B.n417 VSUBS 0.006304f
C471 B.n418 VSUBS 0.006304f
C472 B.n419 VSUBS 0.006304f
C473 B.n420 VSUBS 0.006304f
C474 B.n421 VSUBS 0.006304f
C475 B.n422 VSUBS 0.006304f
C476 B.n423 VSUBS 0.006304f
C477 B.n424 VSUBS 0.006304f
C478 B.n425 VSUBS 0.006304f
C479 B.n426 VSUBS 0.006304f
C480 B.n427 VSUBS 0.006304f
C481 B.n428 VSUBS 0.006304f
C482 B.n429 VSUBS 0.006304f
C483 B.n430 VSUBS 0.006304f
C484 B.n431 VSUBS 0.006304f
C485 B.n432 VSUBS 0.006304f
C486 B.n433 VSUBS 0.006304f
C487 B.n434 VSUBS 0.006304f
C488 B.n435 VSUBS 0.006304f
C489 B.n436 VSUBS 0.006304f
C490 B.n437 VSUBS 0.006304f
C491 B.n438 VSUBS 0.006304f
C492 B.n439 VSUBS 0.006304f
C493 B.n440 VSUBS 0.006304f
C494 B.n441 VSUBS 0.006304f
C495 B.n442 VSUBS 0.006304f
C496 B.n443 VSUBS 0.006304f
C497 B.n444 VSUBS 0.006304f
C498 B.n445 VSUBS 0.006304f
C499 B.n446 VSUBS 0.006304f
C500 B.n447 VSUBS 0.006304f
C501 B.n448 VSUBS 0.006304f
C502 B.n449 VSUBS 0.006304f
C503 B.n450 VSUBS 0.006304f
C504 B.n451 VSUBS 0.006304f
C505 B.n452 VSUBS 0.006304f
C506 B.n453 VSUBS 0.006304f
C507 B.n454 VSUBS 0.006304f
C508 B.n455 VSUBS 0.006304f
C509 B.n456 VSUBS 0.006304f
C510 B.n457 VSUBS 0.006304f
C511 B.n458 VSUBS 0.006304f
C512 B.n459 VSUBS 0.006304f
C513 B.n460 VSUBS 0.006304f
C514 B.n461 VSUBS 0.006304f
C515 B.n462 VSUBS 0.006304f
C516 B.n463 VSUBS 0.006304f
C517 B.n464 VSUBS 0.006304f
C518 B.n465 VSUBS 0.006304f
C519 B.n466 VSUBS 0.006304f
C520 B.n467 VSUBS 0.006304f
C521 B.n468 VSUBS 0.006304f
C522 B.n469 VSUBS 0.006304f
C523 B.n470 VSUBS 0.006304f
C524 B.n471 VSUBS 0.006304f
C525 B.n472 VSUBS 0.006304f
C526 B.n473 VSUBS 0.006304f
C527 B.n474 VSUBS 0.006304f
C528 B.n475 VSUBS 0.006304f
C529 B.n476 VSUBS 0.006304f
C530 B.n477 VSUBS 0.006304f
C531 B.n478 VSUBS 0.006304f
C532 B.n479 VSUBS 0.006304f
C533 B.n480 VSUBS 0.006304f
C534 B.n481 VSUBS 0.006304f
C535 B.n482 VSUBS 0.006304f
C536 B.n483 VSUBS 0.006304f
C537 B.n484 VSUBS 0.006304f
C538 B.n485 VSUBS 0.006304f
C539 B.n486 VSUBS 0.006304f
C540 B.n487 VSUBS 0.006304f
C541 B.n488 VSUBS 0.006304f
C542 B.n489 VSUBS 0.006304f
C543 B.n490 VSUBS 0.006304f
C544 B.n491 VSUBS 0.006304f
C545 B.n492 VSUBS 0.006304f
C546 B.n493 VSUBS 0.006304f
C547 B.n494 VSUBS 0.006304f
C548 B.n495 VSUBS 0.006304f
C549 B.n496 VSUBS 0.006304f
C550 B.n497 VSUBS 0.006304f
C551 B.n498 VSUBS 0.006304f
C552 B.n499 VSUBS 0.006304f
C553 B.n500 VSUBS 0.006304f
C554 B.n501 VSUBS 0.006304f
C555 B.n502 VSUBS 0.006304f
C556 B.n503 VSUBS 0.006304f
C557 B.n504 VSUBS 0.006304f
C558 B.n505 VSUBS 0.006304f
C559 B.n506 VSUBS 0.006304f
C560 B.n507 VSUBS 0.006304f
C561 B.n508 VSUBS 0.006304f
C562 B.n509 VSUBS 0.006304f
C563 B.n510 VSUBS 0.0154f
C564 B.n511 VSUBS 0.014681f
C565 B.n512 VSUBS 0.01554f
C566 B.n513 VSUBS 0.006304f
C567 B.n514 VSUBS 0.006304f
C568 B.n515 VSUBS 0.006304f
C569 B.n516 VSUBS 0.006304f
C570 B.n517 VSUBS 0.006304f
C571 B.n518 VSUBS 0.006304f
C572 B.n519 VSUBS 0.006304f
C573 B.n520 VSUBS 0.006304f
C574 B.n521 VSUBS 0.006304f
C575 B.n522 VSUBS 0.006304f
C576 B.n523 VSUBS 0.006304f
C577 B.n524 VSUBS 0.006304f
C578 B.n525 VSUBS 0.006304f
C579 B.n526 VSUBS 0.006304f
C580 B.n527 VSUBS 0.006304f
C581 B.n528 VSUBS 0.006304f
C582 B.n529 VSUBS 0.006304f
C583 B.n530 VSUBS 0.006304f
C584 B.n531 VSUBS 0.006304f
C585 B.n532 VSUBS 0.006304f
C586 B.n533 VSUBS 0.006304f
C587 B.n534 VSUBS 0.006304f
C588 B.n535 VSUBS 0.006304f
C589 B.n536 VSUBS 0.006304f
C590 B.n537 VSUBS 0.006304f
C591 B.n538 VSUBS 0.006304f
C592 B.n539 VSUBS 0.006304f
C593 B.n540 VSUBS 0.006304f
C594 B.n541 VSUBS 0.006304f
C595 B.n542 VSUBS 0.006304f
C596 B.n543 VSUBS 0.006304f
C597 B.n544 VSUBS 0.006304f
C598 B.n545 VSUBS 0.006304f
C599 B.n546 VSUBS 0.006304f
C600 B.n547 VSUBS 0.006304f
C601 B.n548 VSUBS 0.006304f
C602 B.n549 VSUBS 0.006304f
C603 B.n550 VSUBS 0.006304f
C604 B.n551 VSUBS 0.006304f
C605 B.n552 VSUBS 0.006304f
C606 B.n553 VSUBS 0.006304f
C607 B.n554 VSUBS 0.006304f
C608 B.n555 VSUBS 0.006304f
C609 B.n556 VSUBS 0.006304f
C610 B.n557 VSUBS 0.006304f
C611 B.n558 VSUBS 0.006304f
C612 B.n559 VSUBS 0.006304f
C613 B.n560 VSUBS 0.006304f
C614 B.n561 VSUBS 0.006304f
C615 B.n562 VSUBS 0.006304f
C616 B.n563 VSUBS 0.006304f
C617 B.n564 VSUBS 0.006304f
C618 B.n565 VSUBS 0.006304f
C619 B.n566 VSUBS 0.006304f
C620 B.n567 VSUBS 0.006304f
C621 B.n568 VSUBS 0.006304f
C622 B.n569 VSUBS 0.006304f
C623 B.n570 VSUBS 0.006304f
C624 B.n571 VSUBS 0.006304f
C625 B.n572 VSUBS 0.006304f
C626 B.n573 VSUBS 0.006304f
C627 B.n574 VSUBS 0.006304f
C628 B.n575 VSUBS 0.006304f
C629 B.n576 VSUBS 0.006304f
C630 B.n577 VSUBS 0.006304f
C631 B.n578 VSUBS 0.006304f
C632 B.n579 VSUBS 0.006304f
C633 B.n580 VSUBS 0.006304f
C634 B.n581 VSUBS 0.006304f
C635 B.n582 VSUBS 0.006304f
C636 B.n583 VSUBS 0.006304f
C637 B.n584 VSUBS 0.006304f
C638 B.n585 VSUBS 0.006304f
C639 B.n586 VSUBS 0.006304f
C640 B.n587 VSUBS 0.004357f
C641 B.n588 VSUBS 0.014605f
C642 B.n589 VSUBS 0.005099f
C643 B.n590 VSUBS 0.006304f
C644 B.n591 VSUBS 0.006304f
C645 B.n592 VSUBS 0.006304f
C646 B.n593 VSUBS 0.006304f
C647 B.n594 VSUBS 0.006304f
C648 B.n595 VSUBS 0.006304f
C649 B.n596 VSUBS 0.006304f
C650 B.n597 VSUBS 0.006304f
C651 B.n598 VSUBS 0.006304f
C652 B.n599 VSUBS 0.006304f
C653 B.n600 VSUBS 0.006304f
C654 B.n601 VSUBS 0.005099f
C655 B.n602 VSUBS 0.006304f
C656 B.n603 VSUBS 0.006304f
C657 B.n604 VSUBS 0.006304f
C658 B.n605 VSUBS 0.006304f
C659 B.n606 VSUBS 0.006304f
C660 B.n607 VSUBS 0.006304f
C661 B.n608 VSUBS 0.006304f
C662 B.n609 VSUBS 0.006304f
C663 B.n610 VSUBS 0.006304f
C664 B.n611 VSUBS 0.006304f
C665 B.n612 VSUBS 0.006304f
C666 B.n613 VSUBS 0.006304f
C667 B.n614 VSUBS 0.006304f
C668 B.n615 VSUBS 0.006304f
C669 B.n616 VSUBS 0.006304f
C670 B.n617 VSUBS 0.006304f
C671 B.n618 VSUBS 0.006304f
C672 B.n619 VSUBS 0.006304f
C673 B.n620 VSUBS 0.006304f
C674 B.n621 VSUBS 0.006304f
C675 B.n622 VSUBS 0.006304f
C676 B.n623 VSUBS 0.006304f
C677 B.n624 VSUBS 0.006304f
C678 B.n625 VSUBS 0.006304f
C679 B.n626 VSUBS 0.006304f
C680 B.n627 VSUBS 0.006304f
C681 B.n628 VSUBS 0.006304f
C682 B.n629 VSUBS 0.006304f
C683 B.n630 VSUBS 0.006304f
C684 B.n631 VSUBS 0.006304f
C685 B.n632 VSUBS 0.006304f
C686 B.n633 VSUBS 0.006304f
C687 B.n634 VSUBS 0.006304f
C688 B.n635 VSUBS 0.006304f
C689 B.n636 VSUBS 0.006304f
C690 B.n637 VSUBS 0.006304f
C691 B.n638 VSUBS 0.006304f
C692 B.n639 VSUBS 0.006304f
C693 B.n640 VSUBS 0.006304f
C694 B.n641 VSUBS 0.006304f
C695 B.n642 VSUBS 0.006304f
C696 B.n643 VSUBS 0.006304f
C697 B.n644 VSUBS 0.006304f
C698 B.n645 VSUBS 0.006304f
C699 B.n646 VSUBS 0.006304f
C700 B.n647 VSUBS 0.006304f
C701 B.n648 VSUBS 0.006304f
C702 B.n649 VSUBS 0.006304f
C703 B.n650 VSUBS 0.006304f
C704 B.n651 VSUBS 0.006304f
C705 B.n652 VSUBS 0.006304f
C706 B.n653 VSUBS 0.006304f
C707 B.n654 VSUBS 0.006304f
C708 B.n655 VSUBS 0.006304f
C709 B.n656 VSUBS 0.006304f
C710 B.n657 VSUBS 0.006304f
C711 B.n658 VSUBS 0.006304f
C712 B.n659 VSUBS 0.006304f
C713 B.n660 VSUBS 0.006304f
C714 B.n661 VSUBS 0.006304f
C715 B.n662 VSUBS 0.006304f
C716 B.n663 VSUBS 0.006304f
C717 B.n664 VSUBS 0.006304f
C718 B.n665 VSUBS 0.006304f
C719 B.n666 VSUBS 0.006304f
C720 B.n667 VSUBS 0.006304f
C721 B.n668 VSUBS 0.006304f
C722 B.n669 VSUBS 0.006304f
C723 B.n670 VSUBS 0.006304f
C724 B.n671 VSUBS 0.006304f
C725 B.n672 VSUBS 0.006304f
C726 B.n673 VSUBS 0.006304f
C727 B.n674 VSUBS 0.006304f
C728 B.n675 VSUBS 0.006304f
C729 B.n676 VSUBS 0.006304f
C730 B.n677 VSUBS 0.006304f
C731 B.n678 VSUBS 0.01554f
C732 B.n679 VSUBS 0.014681f
C733 B.n680 VSUBS 0.014681f
C734 B.n681 VSUBS 0.006304f
C735 B.n682 VSUBS 0.006304f
C736 B.n683 VSUBS 0.006304f
C737 B.n684 VSUBS 0.006304f
C738 B.n685 VSUBS 0.006304f
C739 B.n686 VSUBS 0.006304f
C740 B.n687 VSUBS 0.006304f
C741 B.n688 VSUBS 0.006304f
C742 B.n689 VSUBS 0.006304f
C743 B.n690 VSUBS 0.006304f
C744 B.n691 VSUBS 0.006304f
C745 B.n692 VSUBS 0.006304f
C746 B.n693 VSUBS 0.006304f
C747 B.n694 VSUBS 0.006304f
C748 B.n695 VSUBS 0.006304f
C749 B.n696 VSUBS 0.006304f
C750 B.n697 VSUBS 0.006304f
C751 B.n698 VSUBS 0.006304f
C752 B.n699 VSUBS 0.006304f
C753 B.n700 VSUBS 0.006304f
C754 B.n701 VSUBS 0.006304f
C755 B.n702 VSUBS 0.006304f
C756 B.n703 VSUBS 0.006304f
C757 B.n704 VSUBS 0.006304f
C758 B.n705 VSUBS 0.006304f
C759 B.n706 VSUBS 0.006304f
C760 B.n707 VSUBS 0.006304f
C761 B.n708 VSUBS 0.006304f
C762 B.n709 VSUBS 0.006304f
C763 B.n710 VSUBS 0.006304f
C764 B.n711 VSUBS 0.006304f
C765 B.n712 VSUBS 0.006304f
C766 B.n713 VSUBS 0.006304f
C767 B.n714 VSUBS 0.006304f
C768 B.n715 VSUBS 0.006304f
C769 B.n716 VSUBS 0.006304f
C770 B.n717 VSUBS 0.006304f
C771 B.n718 VSUBS 0.006304f
C772 B.n719 VSUBS 0.006304f
C773 B.n720 VSUBS 0.006304f
C774 B.n721 VSUBS 0.006304f
C775 B.n722 VSUBS 0.006304f
C776 B.n723 VSUBS 0.006304f
C777 B.n724 VSUBS 0.006304f
C778 B.n725 VSUBS 0.006304f
C779 B.n726 VSUBS 0.006304f
C780 B.n727 VSUBS 0.006304f
C781 B.n728 VSUBS 0.006304f
C782 B.n729 VSUBS 0.006304f
C783 B.n730 VSUBS 0.006304f
C784 B.n731 VSUBS 0.014274f
C785 VTAIL.t2 VSUBS 2.74071f
C786 VTAIL.n0 VSUBS 0.758621f
C787 VTAIL.t5 VSUBS 2.74071f
C788 VTAIL.n1 VSUBS 0.84806f
C789 VTAIL.t6 VSUBS 2.74071f
C790 VTAIL.n2 VSUBS 2.27051f
C791 VTAIL.t3 VSUBS 2.74072f
C792 VTAIL.n3 VSUBS 2.27051f
C793 VTAIL.t1 VSUBS 2.74072f
C794 VTAIL.n4 VSUBS 0.848056f
C795 VTAIL.t7 VSUBS 2.74072f
C796 VTAIL.n5 VSUBS 0.848056f
C797 VTAIL.t4 VSUBS 2.74071f
C798 VTAIL.n6 VSUBS 2.27051f
C799 VTAIL.t0 VSUBS 2.74071f
C800 VTAIL.n7 VSUBS 2.1725f
C801 VDD1.t0 VSUBS 0.31773f
C802 VDD1.t2 VSUBS 0.31773f
C803 VDD1.n0 VSUBS 2.58752f
C804 VDD1.t3 VSUBS 0.31773f
C805 VDD1.t1 VSUBS 0.31773f
C806 VDD1.n1 VSUBS 3.43253f
C807 VP.n0 VSUBS 0.04177f
C808 VP.t2 VSUBS 3.43276f
C809 VP.n1 VSUBS 0.04625f
C810 VP.n2 VSUBS 0.031682f
C811 VP.t1 VSUBS 3.43276f
C812 VP.n3 VSUBS 1.3083f
C813 VP.t3 VSUBS 3.71857f
C814 VP.t0 VSUBS 3.72465f
C815 VP.n4 VSUBS 4.19006f
C816 VP.n5 VSUBS 1.88414f
C817 VP.n6 VSUBS 0.04177f
C818 VP.n7 VSUBS 0.043012f
C819 VP.n8 VSUBS 0.059047f
C820 VP.n9 VSUBS 0.04625f
C821 VP.n10 VSUBS 0.031682f
C822 VP.n11 VSUBS 0.031682f
C823 VP.n12 VSUBS 0.031682f
C824 VP.n13 VSUBS 0.059047f
C825 VP.n14 VSUBS 0.043012f
C826 VP.n15 VSUBS 1.3083f
C827 VP.n16 VSUBS 0.050873f
.ends

