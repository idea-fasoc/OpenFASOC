* NGSPICE file created from diff_pair_sample_0378.ext - technology: sky130A

.subckt diff_pair_sample_0378 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X1 VDD1.t7 VP.t0 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=1.8057 ps=10.04 w=4.63 l=1.24
X2 VDD1.t6 VP.t1 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X3 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0 ps=0 w=4.63 l=1.24
X4 VTAIL.t12 VN.t1 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X5 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X6 VDD1.t4 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X7 VTAIL.t8 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X8 VTAIL.t13 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0.76395 ps=4.96 w=4.63 l=1.24
X9 VTAIL.t11 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0.76395 ps=4.96 w=4.63 l=1.24
X10 VDD2.t3 VN.t4 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=1.8057 ps=10.04 w=4.63 l=1.24
X11 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0.76395 ps=4.96 w=4.63 l=1.24
X12 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X13 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0 ps=0 w=4.63 l=1.24
X14 VDD2.t2 VN.t5 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=1.8057 ps=10.04 w=4.63 l=1.24
X15 VTAIL.t6 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0.76395 ps=4.96 w=4.63 l=1.24
X16 VDD2.t0 VN.t7 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=0.76395 ps=4.96 w=4.63 l=1.24
X17 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0 ps=0 w=4.63 l=1.24
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8057 pd=10.04 as=0 ps=0 w=4.63 l=1.24
X19 VDD1.t0 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76395 pd=4.96 as=1.8057 ps=10.04 w=4.63 l=1.24
R0 VN.n27 VN.n15 161.3
R1 VN.n26 VN.n25 161.3
R2 VN.n24 VN.n23 161.3
R3 VN.n22 VN.n17 161.3
R4 VN.n21 VN.n20 161.3
R5 VN.n12 VN.n0 161.3
R6 VN.n11 VN.n10 161.3
R7 VN.n9 VN.n8 161.3
R8 VN.n7 VN.n2 161.3
R9 VN.n6 VN.n5 161.3
R10 VN.n4 VN.t6 141.601
R11 VN.n19 VN.t5 141.601
R12 VN.n13 VN.t4 121.861
R13 VN.n28 VN.t3 121.861
R14 VN.n3 VN.t0 89.9868
R15 VN.n1 VN.t2 89.9868
R16 VN.n18 VN.t1 89.9868
R17 VN.n16 VN.t7 89.9868
R18 VN.n29 VN.n28 80.6037
R19 VN.n14 VN.n13 80.6037
R20 VN.n4 VN.n3 43.5433
R21 VN.n19 VN.n18 43.5433
R22 VN.n7 VN.n6 40.4934
R23 VN.n8 VN.n7 40.4934
R24 VN.n22 VN.n21 40.4934
R25 VN.n23 VN.n22 40.4934
R26 VN VN.n29 39.4006
R27 VN.n13 VN.n12 34.3247
R28 VN.n28 VN.n27 34.3247
R29 VN.n12 VN.n11 33.6945
R30 VN.n27 VN.n26 33.6945
R31 VN.n20 VN.n19 29.3131
R32 VN.n5 VN.n4 29.3131
R33 VN.n6 VN.n3 13.9467
R34 VN.n8 VN.n1 13.9467
R35 VN.n21 VN.n18 13.9467
R36 VN.n23 VN.n16 13.9467
R37 VN.n11 VN.n1 10.5213
R38 VN.n26 VN.n16 10.5213
R39 VN.n29 VN.n15 0.285035
R40 VN.n14 VN.n0 0.285035
R41 VN.n25 VN.n15 0.189894
R42 VN.n25 VN.n24 0.189894
R43 VN.n24 VN.n17 0.189894
R44 VN.n20 VN.n17 0.189894
R45 VN.n5 VN.n2 0.189894
R46 VN.n9 VN.n2 0.189894
R47 VN.n10 VN.n9 0.189894
R48 VN.n10 VN.n0 0.189894
R49 VN VN.n14 0.146778
R50 VTAIL.n194 VTAIL.n176 289.615
R51 VTAIL.n20 VTAIL.n2 289.615
R52 VTAIL.n44 VTAIL.n26 289.615
R53 VTAIL.n70 VTAIL.n52 289.615
R54 VTAIL.n170 VTAIL.n152 289.615
R55 VTAIL.n144 VTAIL.n126 289.615
R56 VTAIL.n120 VTAIL.n102 289.615
R57 VTAIL.n94 VTAIL.n76 289.615
R58 VTAIL.n185 VTAIL.n184 185
R59 VTAIL.n187 VTAIL.n186 185
R60 VTAIL.n180 VTAIL.n179 185
R61 VTAIL.n193 VTAIL.n192 185
R62 VTAIL.n195 VTAIL.n194 185
R63 VTAIL.n11 VTAIL.n10 185
R64 VTAIL.n13 VTAIL.n12 185
R65 VTAIL.n6 VTAIL.n5 185
R66 VTAIL.n19 VTAIL.n18 185
R67 VTAIL.n21 VTAIL.n20 185
R68 VTAIL.n35 VTAIL.n34 185
R69 VTAIL.n37 VTAIL.n36 185
R70 VTAIL.n30 VTAIL.n29 185
R71 VTAIL.n43 VTAIL.n42 185
R72 VTAIL.n45 VTAIL.n44 185
R73 VTAIL.n61 VTAIL.n60 185
R74 VTAIL.n63 VTAIL.n62 185
R75 VTAIL.n56 VTAIL.n55 185
R76 VTAIL.n69 VTAIL.n68 185
R77 VTAIL.n71 VTAIL.n70 185
R78 VTAIL.n171 VTAIL.n170 185
R79 VTAIL.n169 VTAIL.n168 185
R80 VTAIL.n156 VTAIL.n155 185
R81 VTAIL.n163 VTAIL.n162 185
R82 VTAIL.n161 VTAIL.n160 185
R83 VTAIL.n145 VTAIL.n144 185
R84 VTAIL.n143 VTAIL.n142 185
R85 VTAIL.n130 VTAIL.n129 185
R86 VTAIL.n137 VTAIL.n136 185
R87 VTAIL.n135 VTAIL.n134 185
R88 VTAIL.n121 VTAIL.n120 185
R89 VTAIL.n119 VTAIL.n118 185
R90 VTAIL.n106 VTAIL.n105 185
R91 VTAIL.n113 VTAIL.n112 185
R92 VTAIL.n111 VTAIL.n110 185
R93 VTAIL.n95 VTAIL.n94 185
R94 VTAIL.n93 VTAIL.n92 185
R95 VTAIL.n80 VTAIL.n79 185
R96 VTAIL.n87 VTAIL.n86 185
R97 VTAIL.n85 VTAIL.n84 185
R98 VTAIL.n183 VTAIL.t10 147.714
R99 VTAIL.n9 VTAIL.t6 147.714
R100 VTAIL.n33 VTAIL.t2 147.714
R101 VTAIL.n59 VTAIL.t4 147.714
R102 VTAIL.n159 VTAIL.t15 147.714
R103 VTAIL.n133 VTAIL.t13 147.714
R104 VTAIL.n109 VTAIL.t7 147.714
R105 VTAIL.n83 VTAIL.t11 147.714
R106 VTAIL.n186 VTAIL.n185 104.615
R107 VTAIL.n186 VTAIL.n179 104.615
R108 VTAIL.n193 VTAIL.n179 104.615
R109 VTAIL.n194 VTAIL.n193 104.615
R110 VTAIL.n12 VTAIL.n11 104.615
R111 VTAIL.n12 VTAIL.n5 104.615
R112 VTAIL.n19 VTAIL.n5 104.615
R113 VTAIL.n20 VTAIL.n19 104.615
R114 VTAIL.n36 VTAIL.n35 104.615
R115 VTAIL.n36 VTAIL.n29 104.615
R116 VTAIL.n43 VTAIL.n29 104.615
R117 VTAIL.n44 VTAIL.n43 104.615
R118 VTAIL.n62 VTAIL.n61 104.615
R119 VTAIL.n62 VTAIL.n55 104.615
R120 VTAIL.n69 VTAIL.n55 104.615
R121 VTAIL.n70 VTAIL.n69 104.615
R122 VTAIL.n170 VTAIL.n169 104.615
R123 VTAIL.n169 VTAIL.n155 104.615
R124 VTAIL.n162 VTAIL.n155 104.615
R125 VTAIL.n162 VTAIL.n161 104.615
R126 VTAIL.n144 VTAIL.n143 104.615
R127 VTAIL.n143 VTAIL.n129 104.615
R128 VTAIL.n136 VTAIL.n129 104.615
R129 VTAIL.n136 VTAIL.n135 104.615
R130 VTAIL.n120 VTAIL.n119 104.615
R131 VTAIL.n119 VTAIL.n105 104.615
R132 VTAIL.n112 VTAIL.n105 104.615
R133 VTAIL.n112 VTAIL.n111 104.615
R134 VTAIL.n94 VTAIL.n93 104.615
R135 VTAIL.n93 VTAIL.n79 104.615
R136 VTAIL.n86 VTAIL.n79 104.615
R137 VTAIL.n86 VTAIL.n85 104.615
R138 VTAIL.n151 VTAIL.n150 55.3206
R139 VTAIL.n101 VTAIL.n100 55.3206
R140 VTAIL.n1 VTAIL.n0 55.3204
R141 VTAIL.n51 VTAIL.n50 55.3204
R142 VTAIL.n185 VTAIL.t10 52.3082
R143 VTAIL.n11 VTAIL.t6 52.3082
R144 VTAIL.n35 VTAIL.t2 52.3082
R145 VTAIL.n61 VTAIL.t4 52.3082
R146 VTAIL.n161 VTAIL.t15 52.3082
R147 VTAIL.n135 VTAIL.t13 52.3082
R148 VTAIL.n111 VTAIL.t7 52.3082
R149 VTAIL.n85 VTAIL.t11 52.3082
R150 VTAIL.n199 VTAIL.n198 33.5429
R151 VTAIL.n25 VTAIL.n24 33.5429
R152 VTAIL.n49 VTAIL.n48 33.5429
R153 VTAIL.n75 VTAIL.n74 33.5429
R154 VTAIL.n175 VTAIL.n174 33.5429
R155 VTAIL.n149 VTAIL.n148 33.5429
R156 VTAIL.n125 VTAIL.n124 33.5429
R157 VTAIL.n99 VTAIL.n98 33.5429
R158 VTAIL.n199 VTAIL.n175 17.7117
R159 VTAIL.n99 VTAIL.n75 17.7117
R160 VTAIL.n184 VTAIL.n183 15.6631
R161 VTAIL.n10 VTAIL.n9 15.6631
R162 VTAIL.n34 VTAIL.n33 15.6631
R163 VTAIL.n60 VTAIL.n59 15.6631
R164 VTAIL.n160 VTAIL.n159 15.6631
R165 VTAIL.n134 VTAIL.n133 15.6631
R166 VTAIL.n110 VTAIL.n109 15.6631
R167 VTAIL.n84 VTAIL.n83 15.6631
R168 VTAIL.n187 VTAIL.n182 12.8005
R169 VTAIL.n13 VTAIL.n8 12.8005
R170 VTAIL.n37 VTAIL.n32 12.8005
R171 VTAIL.n63 VTAIL.n58 12.8005
R172 VTAIL.n163 VTAIL.n158 12.8005
R173 VTAIL.n137 VTAIL.n132 12.8005
R174 VTAIL.n113 VTAIL.n108 12.8005
R175 VTAIL.n87 VTAIL.n82 12.8005
R176 VTAIL.n188 VTAIL.n180 12.0247
R177 VTAIL.n14 VTAIL.n6 12.0247
R178 VTAIL.n38 VTAIL.n30 12.0247
R179 VTAIL.n64 VTAIL.n56 12.0247
R180 VTAIL.n164 VTAIL.n156 12.0247
R181 VTAIL.n138 VTAIL.n130 12.0247
R182 VTAIL.n114 VTAIL.n106 12.0247
R183 VTAIL.n88 VTAIL.n80 12.0247
R184 VTAIL.n192 VTAIL.n191 11.249
R185 VTAIL.n18 VTAIL.n17 11.249
R186 VTAIL.n42 VTAIL.n41 11.249
R187 VTAIL.n68 VTAIL.n67 11.249
R188 VTAIL.n168 VTAIL.n167 11.249
R189 VTAIL.n142 VTAIL.n141 11.249
R190 VTAIL.n118 VTAIL.n117 11.249
R191 VTAIL.n92 VTAIL.n91 11.249
R192 VTAIL.n195 VTAIL.n178 10.4732
R193 VTAIL.n21 VTAIL.n4 10.4732
R194 VTAIL.n45 VTAIL.n28 10.4732
R195 VTAIL.n71 VTAIL.n54 10.4732
R196 VTAIL.n171 VTAIL.n154 10.4732
R197 VTAIL.n145 VTAIL.n128 10.4732
R198 VTAIL.n121 VTAIL.n104 10.4732
R199 VTAIL.n95 VTAIL.n78 10.4732
R200 VTAIL.n196 VTAIL.n176 9.69747
R201 VTAIL.n22 VTAIL.n2 9.69747
R202 VTAIL.n46 VTAIL.n26 9.69747
R203 VTAIL.n72 VTAIL.n52 9.69747
R204 VTAIL.n172 VTAIL.n152 9.69747
R205 VTAIL.n146 VTAIL.n126 9.69747
R206 VTAIL.n122 VTAIL.n102 9.69747
R207 VTAIL.n96 VTAIL.n76 9.69747
R208 VTAIL.n198 VTAIL.n197 9.45567
R209 VTAIL.n24 VTAIL.n23 9.45567
R210 VTAIL.n48 VTAIL.n47 9.45567
R211 VTAIL.n74 VTAIL.n73 9.45567
R212 VTAIL.n174 VTAIL.n173 9.45567
R213 VTAIL.n148 VTAIL.n147 9.45567
R214 VTAIL.n124 VTAIL.n123 9.45567
R215 VTAIL.n98 VTAIL.n97 9.45567
R216 VTAIL.n197 VTAIL.n196 9.3005
R217 VTAIL.n178 VTAIL.n177 9.3005
R218 VTAIL.n191 VTAIL.n190 9.3005
R219 VTAIL.n189 VTAIL.n188 9.3005
R220 VTAIL.n182 VTAIL.n181 9.3005
R221 VTAIL.n23 VTAIL.n22 9.3005
R222 VTAIL.n4 VTAIL.n3 9.3005
R223 VTAIL.n17 VTAIL.n16 9.3005
R224 VTAIL.n15 VTAIL.n14 9.3005
R225 VTAIL.n8 VTAIL.n7 9.3005
R226 VTAIL.n47 VTAIL.n46 9.3005
R227 VTAIL.n28 VTAIL.n27 9.3005
R228 VTAIL.n41 VTAIL.n40 9.3005
R229 VTAIL.n39 VTAIL.n38 9.3005
R230 VTAIL.n32 VTAIL.n31 9.3005
R231 VTAIL.n73 VTAIL.n72 9.3005
R232 VTAIL.n54 VTAIL.n53 9.3005
R233 VTAIL.n67 VTAIL.n66 9.3005
R234 VTAIL.n65 VTAIL.n64 9.3005
R235 VTAIL.n58 VTAIL.n57 9.3005
R236 VTAIL.n173 VTAIL.n172 9.3005
R237 VTAIL.n154 VTAIL.n153 9.3005
R238 VTAIL.n167 VTAIL.n166 9.3005
R239 VTAIL.n165 VTAIL.n164 9.3005
R240 VTAIL.n158 VTAIL.n157 9.3005
R241 VTAIL.n147 VTAIL.n146 9.3005
R242 VTAIL.n128 VTAIL.n127 9.3005
R243 VTAIL.n141 VTAIL.n140 9.3005
R244 VTAIL.n139 VTAIL.n138 9.3005
R245 VTAIL.n132 VTAIL.n131 9.3005
R246 VTAIL.n123 VTAIL.n122 9.3005
R247 VTAIL.n104 VTAIL.n103 9.3005
R248 VTAIL.n117 VTAIL.n116 9.3005
R249 VTAIL.n115 VTAIL.n114 9.3005
R250 VTAIL.n108 VTAIL.n107 9.3005
R251 VTAIL.n97 VTAIL.n96 9.3005
R252 VTAIL.n78 VTAIL.n77 9.3005
R253 VTAIL.n91 VTAIL.n90 9.3005
R254 VTAIL.n89 VTAIL.n88 9.3005
R255 VTAIL.n82 VTAIL.n81 9.3005
R256 VTAIL.n183 VTAIL.n181 4.39059
R257 VTAIL.n9 VTAIL.n7 4.39059
R258 VTAIL.n33 VTAIL.n31 4.39059
R259 VTAIL.n59 VTAIL.n57 4.39059
R260 VTAIL.n159 VTAIL.n157 4.39059
R261 VTAIL.n133 VTAIL.n131 4.39059
R262 VTAIL.n109 VTAIL.n107 4.39059
R263 VTAIL.n83 VTAIL.n81 4.39059
R264 VTAIL.n0 VTAIL.t9 4.27696
R265 VTAIL.n0 VTAIL.t8 4.27696
R266 VTAIL.n50 VTAIL.t0 4.27696
R267 VTAIL.n50 VTAIL.t1 4.27696
R268 VTAIL.n150 VTAIL.t14 4.27696
R269 VTAIL.n150 VTAIL.t3 4.27696
R270 VTAIL.n100 VTAIL.t5 4.27696
R271 VTAIL.n100 VTAIL.t12 4.27696
R272 VTAIL.n198 VTAIL.n176 4.26717
R273 VTAIL.n24 VTAIL.n2 4.26717
R274 VTAIL.n48 VTAIL.n26 4.26717
R275 VTAIL.n74 VTAIL.n52 4.26717
R276 VTAIL.n174 VTAIL.n152 4.26717
R277 VTAIL.n148 VTAIL.n126 4.26717
R278 VTAIL.n124 VTAIL.n102 4.26717
R279 VTAIL.n98 VTAIL.n76 4.26717
R280 VTAIL.n196 VTAIL.n195 3.49141
R281 VTAIL.n22 VTAIL.n21 3.49141
R282 VTAIL.n46 VTAIL.n45 3.49141
R283 VTAIL.n72 VTAIL.n71 3.49141
R284 VTAIL.n172 VTAIL.n171 3.49141
R285 VTAIL.n146 VTAIL.n145 3.49141
R286 VTAIL.n122 VTAIL.n121 3.49141
R287 VTAIL.n96 VTAIL.n95 3.49141
R288 VTAIL.n192 VTAIL.n178 2.71565
R289 VTAIL.n18 VTAIL.n4 2.71565
R290 VTAIL.n42 VTAIL.n28 2.71565
R291 VTAIL.n68 VTAIL.n54 2.71565
R292 VTAIL.n168 VTAIL.n154 2.71565
R293 VTAIL.n142 VTAIL.n128 2.71565
R294 VTAIL.n118 VTAIL.n104 2.71565
R295 VTAIL.n92 VTAIL.n78 2.71565
R296 VTAIL.n191 VTAIL.n180 1.93989
R297 VTAIL.n17 VTAIL.n6 1.93989
R298 VTAIL.n41 VTAIL.n30 1.93989
R299 VTAIL.n67 VTAIL.n56 1.93989
R300 VTAIL.n167 VTAIL.n156 1.93989
R301 VTAIL.n141 VTAIL.n130 1.93989
R302 VTAIL.n117 VTAIL.n106 1.93989
R303 VTAIL.n91 VTAIL.n80 1.93989
R304 VTAIL.n101 VTAIL.n99 1.35395
R305 VTAIL.n125 VTAIL.n101 1.35395
R306 VTAIL.n151 VTAIL.n149 1.35395
R307 VTAIL.n175 VTAIL.n151 1.35395
R308 VTAIL.n75 VTAIL.n51 1.35395
R309 VTAIL.n51 VTAIL.n49 1.35395
R310 VTAIL.n25 VTAIL.n1 1.35395
R311 VTAIL VTAIL.n199 1.29576
R312 VTAIL.n188 VTAIL.n187 1.16414
R313 VTAIL.n14 VTAIL.n13 1.16414
R314 VTAIL.n38 VTAIL.n37 1.16414
R315 VTAIL.n64 VTAIL.n63 1.16414
R316 VTAIL.n164 VTAIL.n163 1.16414
R317 VTAIL.n138 VTAIL.n137 1.16414
R318 VTAIL.n114 VTAIL.n113 1.16414
R319 VTAIL.n88 VTAIL.n87 1.16414
R320 VTAIL.n149 VTAIL.n125 0.470328
R321 VTAIL.n49 VTAIL.n25 0.470328
R322 VTAIL.n184 VTAIL.n182 0.388379
R323 VTAIL.n10 VTAIL.n8 0.388379
R324 VTAIL.n34 VTAIL.n32 0.388379
R325 VTAIL.n60 VTAIL.n58 0.388379
R326 VTAIL.n160 VTAIL.n158 0.388379
R327 VTAIL.n134 VTAIL.n132 0.388379
R328 VTAIL.n110 VTAIL.n108 0.388379
R329 VTAIL.n84 VTAIL.n82 0.388379
R330 VTAIL.n189 VTAIL.n181 0.155672
R331 VTAIL.n190 VTAIL.n189 0.155672
R332 VTAIL.n190 VTAIL.n177 0.155672
R333 VTAIL.n197 VTAIL.n177 0.155672
R334 VTAIL.n15 VTAIL.n7 0.155672
R335 VTAIL.n16 VTAIL.n15 0.155672
R336 VTAIL.n16 VTAIL.n3 0.155672
R337 VTAIL.n23 VTAIL.n3 0.155672
R338 VTAIL.n39 VTAIL.n31 0.155672
R339 VTAIL.n40 VTAIL.n39 0.155672
R340 VTAIL.n40 VTAIL.n27 0.155672
R341 VTAIL.n47 VTAIL.n27 0.155672
R342 VTAIL.n65 VTAIL.n57 0.155672
R343 VTAIL.n66 VTAIL.n65 0.155672
R344 VTAIL.n66 VTAIL.n53 0.155672
R345 VTAIL.n73 VTAIL.n53 0.155672
R346 VTAIL.n173 VTAIL.n153 0.155672
R347 VTAIL.n166 VTAIL.n153 0.155672
R348 VTAIL.n166 VTAIL.n165 0.155672
R349 VTAIL.n165 VTAIL.n157 0.155672
R350 VTAIL.n147 VTAIL.n127 0.155672
R351 VTAIL.n140 VTAIL.n127 0.155672
R352 VTAIL.n140 VTAIL.n139 0.155672
R353 VTAIL.n139 VTAIL.n131 0.155672
R354 VTAIL.n123 VTAIL.n103 0.155672
R355 VTAIL.n116 VTAIL.n103 0.155672
R356 VTAIL.n116 VTAIL.n115 0.155672
R357 VTAIL.n115 VTAIL.n107 0.155672
R358 VTAIL.n97 VTAIL.n77 0.155672
R359 VTAIL.n90 VTAIL.n77 0.155672
R360 VTAIL.n90 VTAIL.n89 0.155672
R361 VTAIL.n89 VTAIL.n81 0.155672
R362 VTAIL VTAIL.n1 0.0586897
R363 VDD2.n2 VDD2.n1 72.6206
R364 VDD2.n2 VDD2.n0 72.6206
R365 VDD2 VDD2.n5 72.6178
R366 VDD2.n4 VDD2.n3 71.9994
R367 VDD2.n4 VDD2.n2 33.7972
R368 VDD2.n5 VDD2.t6 4.27696
R369 VDD2.n5 VDD2.t2 4.27696
R370 VDD2.n3 VDD2.t4 4.27696
R371 VDD2.n3 VDD2.t0 4.27696
R372 VDD2.n1 VDD2.t5 4.27696
R373 VDD2.n1 VDD2.t3 4.27696
R374 VDD2.n0 VDD2.t1 4.27696
R375 VDD2.n0 VDD2.t7 4.27696
R376 VDD2 VDD2.n4 0.735414
R377 B.n504 B.n503 585
R378 B.n505 B.n504 585
R379 B.n182 B.n84 585
R380 B.n181 B.n180 585
R381 B.n179 B.n178 585
R382 B.n177 B.n176 585
R383 B.n175 B.n174 585
R384 B.n173 B.n172 585
R385 B.n171 B.n170 585
R386 B.n169 B.n168 585
R387 B.n167 B.n166 585
R388 B.n165 B.n164 585
R389 B.n163 B.n162 585
R390 B.n161 B.n160 585
R391 B.n159 B.n158 585
R392 B.n157 B.n156 585
R393 B.n155 B.n154 585
R394 B.n153 B.n152 585
R395 B.n151 B.n150 585
R396 B.n149 B.n148 585
R397 B.n147 B.n146 585
R398 B.n144 B.n143 585
R399 B.n142 B.n141 585
R400 B.n140 B.n139 585
R401 B.n138 B.n137 585
R402 B.n136 B.n135 585
R403 B.n134 B.n133 585
R404 B.n132 B.n131 585
R405 B.n130 B.n129 585
R406 B.n128 B.n127 585
R407 B.n126 B.n125 585
R408 B.n124 B.n123 585
R409 B.n122 B.n121 585
R410 B.n120 B.n119 585
R411 B.n118 B.n117 585
R412 B.n116 B.n115 585
R413 B.n114 B.n113 585
R414 B.n112 B.n111 585
R415 B.n110 B.n109 585
R416 B.n108 B.n107 585
R417 B.n106 B.n105 585
R418 B.n104 B.n103 585
R419 B.n102 B.n101 585
R420 B.n100 B.n99 585
R421 B.n98 B.n97 585
R422 B.n96 B.n95 585
R423 B.n94 B.n93 585
R424 B.n92 B.n91 585
R425 B.n60 B.n59 585
R426 B.n508 B.n507 585
R427 B.n502 B.n85 585
R428 B.n85 B.n57 585
R429 B.n501 B.n56 585
R430 B.n512 B.n56 585
R431 B.n500 B.n55 585
R432 B.n513 B.n55 585
R433 B.n499 B.n54 585
R434 B.n514 B.n54 585
R435 B.n498 B.n497 585
R436 B.n497 B.n50 585
R437 B.n496 B.n49 585
R438 B.n520 B.n49 585
R439 B.n495 B.n48 585
R440 B.n521 B.n48 585
R441 B.n494 B.n47 585
R442 B.n522 B.n47 585
R443 B.n493 B.n492 585
R444 B.n492 B.n43 585
R445 B.n491 B.n42 585
R446 B.n528 B.n42 585
R447 B.n490 B.n41 585
R448 B.n529 B.n41 585
R449 B.n489 B.n40 585
R450 B.n530 B.n40 585
R451 B.n488 B.n487 585
R452 B.n487 B.n36 585
R453 B.n486 B.n35 585
R454 B.n536 B.n35 585
R455 B.n485 B.n34 585
R456 B.n537 B.n34 585
R457 B.n484 B.n33 585
R458 B.n538 B.n33 585
R459 B.n483 B.n482 585
R460 B.n482 B.n29 585
R461 B.n481 B.n28 585
R462 B.n544 B.n28 585
R463 B.n480 B.n27 585
R464 B.n545 B.n27 585
R465 B.n479 B.n26 585
R466 B.n546 B.n26 585
R467 B.n478 B.n477 585
R468 B.n477 B.n22 585
R469 B.n476 B.n21 585
R470 B.n552 B.n21 585
R471 B.n475 B.n20 585
R472 B.n553 B.n20 585
R473 B.n474 B.n19 585
R474 B.n554 B.n19 585
R475 B.n473 B.n472 585
R476 B.n472 B.n15 585
R477 B.n471 B.n14 585
R478 B.n560 B.n14 585
R479 B.n470 B.n13 585
R480 B.n561 B.n13 585
R481 B.n469 B.n12 585
R482 B.n562 B.n12 585
R483 B.n468 B.n467 585
R484 B.n467 B.n8 585
R485 B.n466 B.n7 585
R486 B.n568 B.n7 585
R487 B.n465 B.n6 585
R488 B.n569 B.n6 585
R489 B.n464 B.n5 585
R490 B.n570 B.n5 585
R491 B.n463 B.n462 585
R492 B.n462 B.n4 585
R493 B.n461 B.n183 585
R494 B.n461 B.n460 585
R495 B.n451 B.n184 585
R496 B.n185 B.n184 585
R497 B.n453 B.n452 585
R498 B.n454 B.n453 585
R499 B.n450 B.n190 585
R500 B.n190 B.n189 585
R501 B.n449 B.n448 585
R502 B.n448 B.n447 585
R503 B.n192 B.n191 585
R504 B.n193 B.n192 585
R505 B.n440 B.n439 585
R506 B.n441 B.n440 585
R507 B.n438 B.n197 585
R508 B.n201 B.n197 585
R509 B.n437 B.n436 585
R510 B.n436 B.n435 585
R511 B.n199 B.n198 585
R512 B.n200 B.n199 585
R513 B.n428 B.n427 585
R514 B.n429 B.n428 585
R515 B.n426 B.n206 585
R516 B.n206 B.n205 585
R517 B.n425 B.n424 585
R518 B.n424 B.n423 585
R519 B.n208 B.n207 585
R520 B.n209 B.n208 585
R521 B.n416 B.n415 585
R522 B.n417 B.n416 585
R523 B.n414 B.n214 585
R524 B.n214 B.n213 585
R525 B.n413 B.n412 585
R526 B.n412 B.n411 585
R527 B.n216 B.n215 585
R528 B.n217 B.n216 585
R529 B.n404 B.n403 585
R530 B.n405 B.n404 585
R531 B.n402 B.n222 585
R532 B.n222 B.n221 585
R533 B.n401 B.n400 585
R534 B.n400 B.n399 585
R535 B.n224 B.n223 585
R536 B.n225 B.n224 585
R537 B.n392 B.n391 585
R538 B.n393 B.n392 585
R539 B.n390 B.n230 585
R540 B.n230 B.n229 585
R541 B.n389 B.n388 585
R542 B.n388 B.n387 585
R543 B.n232 B.n231 585
R544 B.n233 B.n232 585
R545 B.n380 B.n379 585
R546 B.n381 B.n380 585
R547 B.n378 B.n238 585
R548 B.n238 B.n237 585
R549 B.n377 B.n376 585
R550 B.n376 B.n375 585
R551 B.n240 B.n239 585
R552 B.n241 B.n240 585
R553 B.n371 B.n370 585
R554 B.n244 B.n243 585
R555 B.n367 B.n366 585
R556 B.n368 B.n367 585
R557 B.n365 B.n268 585
R558 B.n364 B.n363 585
R559 B.n362 B.n361 585
R560 B.n360 B.n359 585
R561 B.n358 B.n357 585
R562 B.n356 B.n355 585
R563 B.n354 B.n353 585
R564 B.n352 B.n351 585
R565 B.n350 B.n349 585
R566 B.n348 B.n347 585
R567 B.n346 B.n345 585
R568 B.n344 B.n343 585
R569 B.n342 B.n341 585
R570 B.n340 B.n339 585
R571 B.n338 B.n337 585
R572 B.n336 B.n335 585
R573 B.n334 B.n333 585
R574 B.n331 B.n330 585
R575 B.n329 B.n328 585
R576 B.n327 B.n326 585
R577 B.n325 B.n324 585
R578 B.n323 B.n322 585
R579 B.n321 B.n320 585
R580 B.n319 B.n318 585
R581 B.n317 B.n316 585
R582 B.n315 B.n314 585
R583 B.n313 B.n312 585
R584 B.n311 B.n310 585
R585 B.n309 B.n308 585
R586 B.n307 B.n306 585
R587 B.n305 B.n304 585
R588 B.n303 B.n302 585
R589 B.n301 B.n300 585
R590 B.n299 B.n298 585
R591 B.n297 B.n296 585
R592 B.n295 B.n294 585
R593 B.n293 B.n292 585
R594 B.n291 B.n290 585
R595 B.n289 B.n288 585
R596 B.n287 B.n286 585
R597 B.n285 B.n284 585
R598 B.n283 B.n282 585
R599 B.n281 B.n280 585
R600 B.n279 B.n278 585
R601 B.n277 B.n276 585
R602 B.n275 B.n274 585
R603 B.n372 B.n242 585
R604 B.n242 B.n241 585
R605 B.n374 B.n373 585
R606 B.n375 B.n374 585
R607 B.n236 B.n235 585
R608 B.n237 B.n236 585
R609 B.n383 B.n382 585
R610 B.n382 B.n381 585
R611 B.n384 B.n234 585
R612 B.n234 B.n233 585
R613 B.n386 B.n385 585
R614 B.n387 B.n386 585
R615 B.n228 B.n227 585
R616 B.n229 B.n228 585
R617 B.n395 B.n394 585
R618 B.n394 B.n393 585
R619 B.n396 B.n226 585
R620 B.n226 B.n225 585
R621 B.n398 B.n397 585
R622 B.n399 B.n398 585
R623 B.n220 B.n219 585
R624 B.n221 B.n220 585
R625 B.n407 B.n406 585
R626 B.n406 B.n405 585
R627 B.n408 B.n218 585
R628 B.n218 B.n217 585
R629 B.n410 B.n409 585
R630 B.n411 B.n410 585
R631 B.n212 B.n211 585
R632 B.n213 B.n212 585
R633 B.n419 B.n418 585
R634 B.n418 B.n417 585
R635 B.n420 B.n210 585
R636 B.n210 B.n209 585
R637 B.n422 B.n421 585
R638 B.n423 B.n422 585
R639 B.n204 B.n203 585
R640 B.n205 B.n204 585
R641 B.n431 B.n430 585
R642 B.n430 B.n429 585
R643 B.n432 B.n202 585
R644 B.n202 B.n200 585
R645 B.n434 B.n433 585
R646 B.n435 B.n434 585
R647 B.n196 B.n195 585
R648 B.n201 B.n196 585
R649 B.n443 B.n442 585
R650 B.n442 B.n441 585
R651 B.n444 B.n194 585
R652 B.n194 B.n193 585
R653 B.n446 B.n445 585
R654 B.n447 B.n446 585
R655 B.n188 B.n187 585
R656 B.n189 B.n188 585
R657 B.n456 B.n455 585
R658 B.n455 B.n454 585
R659 B.n457 B.n186 585
R660 B.n186 B.n185 585
R661 B.n459 B.n458 585
R662 B.n460 B.n459 585
R663 B.n2 B.n0 585
R664 B.n4 B.n2 585
R665 B.n3 B.n1 585
R666 B.n569 B.n3 585
R667 B.n567 B.n566 585
R668 B.n568 B.n567 585
R669 B.n565 B.n9 585
R670 B.n9 B.n8 585
R671 B.n564 B.n563 585
R672 B.n563 B.n562 585
R673 B.n11 B.n10 585
R674 B.n561 B.n11 585
R675 B.n559 B.n558 585
R676 B.n560 B.n559 585
R677 B.n557 B.n16 585
R678 B.n16 B.n15 585
R679 B.n556 B.n555 585
R680 B.n555 B.n554 585
R681 B.n18 B.n17 585
R682 B.n553 B.n18 585
R683 B.n551 B.n550 585
R684 B.n552 B.n551 585
R685 B.n549 B.n23 585
R686 B.n23 B.n22 585
R687 B.n548 B.n547 585
R688 B.n547 B.n546 585
R689 B.n25 B.n24 585
R690 B.n545 B.n25 585
R691 B.n543 B.n542 585
R692 B.n544 B.n543 585
R693 B.n541 B.n30 585
R694 B.n30 B.n29 585
R695 B.n540 B.n539 585
R696 B.n539 B.n538 585
R697 B.n32 B.n31 585
R698 B.n537 B.n32 585
R699 B.n535 B.n534 585
R700 B.n536 B.n535 585
R701 B.n533 B.n37 585
R702 B.n37 B.n36 585
R703 B.n532 B.n531 585
R704 B.n531 B.n530 585
R705 B.n39 B.n38 585
R706 B.n529 B.n39 585
R707 B.n527 B.n526 585
R708 B.n528 B.n527 585
R709 B.n525 B.n44 585
R710 B.n44 B.n43 585
R711 B.n524 B.n523 585
R712 B.n523 B.n522 585
R713 B.n46 B.n45 585
R714 B.n521 B.n46 585
R715 B.n519 B.n518 585
R716 B.n520 B.n519 585
R717 B.n517 B.n51 585
R718 B.n51 B.n50 585
R719 B.n516 B.n515 585
R720 B.n515 B.n514 585
R721 B.n53 B.n52 585
R722 B.n513 B.n53 585
R723 B.n511 B.n510 585
R724 B.n512 B.n511 585
R725 B.n509 B.n58 585
R726 B.n58 B.n57 585
R727 B.n572 B.n571 585
R728 B.n571 B.n570 585
R729 B.n370 B.n242 569.379
R730 B.n507 B.n58 569.379
R731 B.n274 B.n240 569.379
R732 B.n504 B.n85 569.379
R733 B.n271 B.t8 294.308
R734 B.n269 B.t12 294.308
R735 B.n88 B.t19 294.308
R736 B.n86 B.t15 294.308
R737 B.n505 B.n83 256.663
R738 B.n505 B.n82 256.663
R739 B.n505 B.n81 256.663
R740 B.n505 B.n80 256.663
R741 B.n505 B.n79 256.663
R742 B.n505 B.n78 256.663
R743 B.n505 B.n77 256.663
R744 B.n505 B.n76 256.663
R745 B.n505 B.n75 256.663
R746 B.n505 B.n74 256.663
R747 B.n505 B.n73 256.663
R748 B.n505 B.n72 256.663
R749 B.n505 B.n71 256.663
R750 B.n505 B.n70 256.663
R751 B.n505 B.n69 256.663
R752 B.n505 B.n68 256.663
R753 B.n505 B.n67 256.663
R754 B.n505 B.n66 256.663
R755 B.n505 B.n65 256.663
R756 B.n505 B.n64 256.663
R757 B.n505 B.n63 256.663
R758 B.n505 B.n62 256.663
R759 B.n505 B.n61 256.663
R760 B.n506 B.n505 256.663
R761 B.n369 B.n368 256.663
R762 B.n368 B.n245 256.663
R763 B.n368 B.n246 256.663
R764 B.n368 B.n247 256.663
R765 B.n368 B.n248 256.663
R766 B.n368 B.n249 256.663
R767 B.n368 B.n250 256.663
R768 B.n368 B.n251 256.663
R769 B.n368 B.n252 256.663
R770 B.n368 B.n253 256.663
R771 B.n368 B.n254 256.663
R772 B.n368 B.n255 256.663
R773 B.n368 B.n256 256.663
R774 B.n368 B.n257 256.663
R775 B.n368 B.n258 256.663
R776 B.n368 B.n259 256.663
R777 B.n368 B.n260 256.663
R778 B.n368 B.n261 256.663
R779 B.n368 B.n262 256.663
R780 B.n368 B.n263 256.663
R781 B.n368 B.n264 256.663
R782 B.n368 B.n265 256.663
R783 B.n368 B.n266 256.663
R784 B.n368 B.n267 256.663
R785 B.n271 B.t11 186.06
R786 B.n86 B.t17 186.06
R787 B.n269 B.t14 186.06
R788 B.n88 B.t20 186.06
R789 B.n374 B.n242 163.367
R790 B.n374 B.n236 163.367
R791 B.n382 B.n236 163.367
R792 B.n382 B.n234 163.367
R793 B.n386 B.n234 163.367
R794 B.n386 B.n228 163.367
R795 B.n394 B.n228 163.367
R796 B.n394 B.n226 163.367
R797 B.n398 B.n226 163.367
R798 B.n398 B.n220 163.367
R799 B.n406 B.n220 163.367
R800 B.n406 B.n218 163.367
R801 B.n410 B.n218 163.367
R802 B.n410 B.n212 163.367
R803 B.n418 B.n212 163.367
R804 B.n418 B.n210 163.367
R805 B.n422 B.n210 163.367
R806 B.n422 B.n204 163.367
R807 B.n430 B.n204 163.367
R808 B.n430 B.n202 163.367
R809 B.n434 B.n202 163.367
R810 B.n434 B.n196 163.367
R811 B.n442 B.n196 163.367
R812 B.n442 B.n194 163.367
R813 B.n446 B.n194 163.367
R814 B.n446 B.n188 163.367
R815 B.n455 B.n188 163.367
R816 B.n455 B.n186 163.367
R817 B.n459 B.n186 163.367
R818 B.n459 B.n2 163.367
R819 B.n571 B.n2 163.367
R820 B.n571 B.n3 163.367
R821 B.n567 B.n3 163.367
R822 B.n567 B.n9 163.367
R823 B.n563 B.n9 163.367
R824 B.n563 B.n11 163.367
R825 B.n559 B.n11 163.367
R826 B.n559 B.n16 163.367
R827 B.n555 B.n16 163.367
R828 B.n555 B.n18 163.367
R829 B.n551 B.n18 163.367
R830 B.n551 B.n23 163.367
R831 B.n547 B.n23 163.367
R832 B.n547 B.n25 163.367
R833 B.n543 B.n25 163.367
R834 B.n543 B.n30 163.367
R835 B.n539 B.n30 163.367
R836 B.n539 B.n32 163.367
R837 B.n535 B.n32 163.367
R838 B.n535 B.n37 163.367
R839 B.n531 B.n37 163.367
R840 B.n531 B.n39 163.367
R841 B.n527 B.n39 163.367
R842 B.n527 B.n44 163.367
R843 B.n523 B.n44 163.367
R844 B.n523 B.n46 163.367
R845 B.n519 B.n46 163.367
R846 B.n519 B.n51 163.367
R847 B.n515 B.n51 163.367
R848 B.n515 B.n53 163.367
R849 B.n511 B.n53 163.367
R850 B.n511 B.n58 163.367
R851 B.n367 B.n244 163.367
R852 B.n367 B.n268 163.367
R853 B.n363 B.n362 163.367
R854 B.n359 B.n358 163.367
R855 B.n355 B.n354 163.367
R856 B.n351 B.n350 163.367
R857 B.n347 B.n346 163.367
R858 B.n343 B.n342 163.367
R859 B.n339 B.n338 163.367
R860 B.n335 B.n334 163.367
R861 B.n330 B.n329 163.367
R862 B.n326 B.n325 163.367
R863 B.n322 B.n321 163.367
R864 B.n318 B.n317 163.367
R865 B.n314 B.n313 163.367
R866 B.n310 B.n309 163.367
R867 B.n306 B.n305 163.367
R868 B.n302 B.n301 163.367
R869 B.n298 B.n297 163.367
R870 B.n294 B.n293 163.367
R871 B.n290 B.n289 163.367
R872 B.n286 B.n285 163.367
R873 B.n282 B.n281 163.367
R874 B.n278 B.n277 163.367
R875 B.n376 B.n240 163.367
R876 B.n376 B.n238 163.367
R877 B.n380 B.n238 163.367
R878 B.n380 B.n232 163.367
R879 B.n388 B.n232 163.367
R880 B.n388 B.n230 163.367
R881 B.n392 B.n230 163.367
R882 B.n392 B.n224 163.367
R883 B.n400 B.n224 163.367
R884 B.n400 B.n222 163.367
R885 B.n404 B.n222 163.367
R886 B.n404 B.n216 163.367
R887 B.n412 B.n216 163.367
R888 B.n412 B.n214 163.367
R889 B.n416 B.n214 163.367
R890 B.n416 B.n208 163.367
R891 B.n424 B.n208 163.367
R892 B.n424 B.n206 163.367
R893 B.n428 B.n206 163.367
R894 B.n428 B.n199 163.367
R895 B.n436 B.n199 163.367
R896 B.n436 B.n197 163.367
R897 B.n440 B.n197 163.367
R898 B.n440 B.n192 163.367
R899 B.n448 B.n192 163.367
R900 B.n448 B.n190 163.367
R901 B.n453 B.n190 163.367
R902 B.n453 B.n184 163.367
R903 B.n461 B.n184 163.367
R904 B.n462 B.n461 163.367
R905 B.n462 B.n5 163.367
R906 B.n6 B.n5 163.367
R907 B.n7 B.n6 163.367
R908 B.n467 B.n7 163.367
R909 B.n467 B.n12 163.367
R910 B.n13 B.n12 163.367
R911 B.n14 B.n13 163.367
R912 B.n472 B.n14 163.367
R913 B.n472 B.n19 163.367
R914 B.n20 B.n19 163.367
R915 B.n21 B.n20 163.367
R916 B.n477 B.n21 163.367
R917 B.n477 B.n26 163.367
R918 B.n27 B.n26 163.367
R919 B.n28 B.n27 163.367
R920 B.n482 B.n28 163.367
R921 B.n482 B.n33 163.367
R922 B.n34 B.n33 163.367
R923 B.n35 B.n34 163.367
R924 B.n487 B.n35 163.367
R925 B.n487 B.n40 163.367
R926 B.n41 B.n40 163.367
R927 B.n42 B.n41 163.367
R928 B.n492 B.n42 163.367
R929 B.n492 B.n47 163.367
R930 B.n48 B.n47 163.367
R931 B.n49 B.n48 163.367
R932 B.n497 B.n49 163.367
R933 B.n497 B.n54 163.367
R934 B.n55 B.n54 163.367
R935 B.n56 B.n55 163.367
R936 B.n85 B.n56 163.367
R937 B.n91 B.n60 163.367
R938 B.n95 B.n94 163.367
R939 B.n99 B.n98 163.367
R940 B.n103 B.n102 163.367
R941 B.n107 B.n106 163.367
R942 B.n111 B.n110 163.367
R943 B.n115 B.n114 163.367
R944 B.n119 B.n118 163.367
R945 B.n123 B.n122 163.367
R946 B.n127 B.n126 163.367
R947 B.n131 B.n130 163.367
R948 B.n135 B.n134 163.367
R949 B.n139 B.n138 163.367
R950 B.n143 B.n142 163.367
R951 B.n148 B.n147 163.367
R952 B.n152 B.n151 163.367
R953 B.n156 B.n155 163.367
R954 B.n160 B.n159 163.367
R955 B.n164 B.n163 163.367
R956 B.n168 B.n167 163.367
R957 B.n172 B.n171 163.367
R958 B.n176 B.n175 163.367
R959 B.n180 B.n179 163.367
R960 B.n504 B.n84 163.367
R961 B.n272 B.t10 155.613
R962 B.n87 B.t18 155.613
R963 B.n270 B.t13 155.613
R964 B.n89 B.t21 155.613
R965 B.n368 B.n241 152.145
R966 B.n505 B.n57 152.145
R967 B.n375 B.n241 75.5179
R968 B.n375 B.n237 75.5179
R969 B.n381 B.n237 75.5179
R970 B.n381 B.n233 75.5179
R971 B.n387 B.n233 75.5179
R972 B.n393 B.n229 75.5179
R973 B.n393 B.n225 75.5179
R974 B.n399 B.n225 75.5179
R975 B.n399 B.n221 75.5179
R976 B.n405 B.n221 75.5179
R977 B.n405 B.n217 75.5179
R978 B.n411 B.n217 75.5179
R979 B.n417 B.n213 75.5179
R980 B.n417 B.n209 75.5179
R981 B.n423 B.n209 75.5179
R982 B.n429 B.n205 75.5179
R983 B.n429 B.n200 75.5179
R984 B.n435 B.n200 75.5179
R985 B.n435 B.n201 75.5179
R986 B.n441 B.n193 75.5179
R987 B.n447 B.n193 75.5179
R988 B.n447 B.n189 75.5179
R989 B.n454 B.n189 75.5179
R990 B.n460 B.n185 75.5179
R991 B.n460 B.n4 75.5179
R992 B.n570 B.n4 75.5179
R993 B.n570 B.n569 75.5179
R994 B.n569 B.n568 75.5179
R995 B.n568 B.n8 75.5179
R996 B.n562 B.n561 75.5179
R997 B.n561 B.n560 75.5179
R998 B.n560 B.n15 75.5179
R999 B.n554 B.n15 75.5179
R1000 B.n553 B.n552 75.5179
R1001 B.n552 B.n22 75.5179
R1002 B.n546 B.n22 75.5179
R1003 B.n546 B.n545 75.5179
R1004 B.n544 B.n29 75.5179
R1005 B.n538 B.n29 75.5179
R1006 B.n538 B.n537 75.5179
R1007 B.n536 B.n36 75.5179
R1008 B.n530 B.n36 75.5179
R1009 B.n530 B.n529 75.5179
R1010 B.n529 B.n528 75.5179
R1011 B.n528 B.n43 75.5179
R1012 B.n522 B.n43 75.5179
R1013 B.n522 B.n521 75.5179
R1014 B.n520 B.n50 75.5179
R1015 B.n514 B.n50 75.5179
R1016 B.n514 B.n513 75.5179
R1017 B.n513 B.n512 75.5179
R1018 B.n512 B.n57 75.5179
R1019 B.n370 B.n369 71.676
R1020 B.n268 B.n245 71.676
R1021 B.n362 B.n246 71.676
R1022 B.n358 B.n247 71.676
R1023 B.n354 B.n248 71.676
R1024 B.n350 B.n249 71.676
R1025 B.n346 B.n250 71.676
R1026 B.n342 B.n251 71.676
R1027 B.n338 B.n252 71.676
R1028 B.n334 B.n253 71.676
R1029 B.n329 B.n254 71.676
R1030 B.n325 B.n255 71.676
R1031 B.n321 B.n256 71.676
R1032 B.n317 B.n257 71.676
R1033 B.n313 B.n258 71.676
R1034 B.n309 B.n259 71.676
R1035 B.n305 B.n260 71.676
R1036 B.n301 B.n261 71.676
R1037 B.n297 B.n262 71.676
R1038 B.n293 B.n263 71.676
R1039 B.n289 B.n264 71.676
R1040 B.n285 B.n265 71.676
R1041 B.n281 B.n266 71.676
R1042 B.n277 B.n267 71.676
R1043 B.n507 B.n506 71.676
R1044 B.n91 B.n61 71.676
R1045 B.n95 B.n62 71.676
R1046 B.n99 B.n63 71.676
R1047 B.n103 B.n64 71.676
R1048 B.n107 B.n65 71.676
R1049 B.n111 B.n66 71.676
R1050 B.n115 B.n67 71.676
R1051 B.n119 B.n68 71.676
R1052 B.n123 B.n69 71.676
R1053 B.n127 B.n70 71.676
R1054 B.n131 B.n71 71.676
R1055 B.n135 B.n72 71.676
R1056 B.n139 B.n73 71.676
R1057 B.n143 B.n74 71.676
R1058 B.n148 B.n75 71.676
R1059 B.n152 B.n76 71.676
R1060 B.n156 B.n77 71.676
R1061 B.n160 B.n78 71.676
R1062 B.n164 B.n79 71.676
R1063 B.n168 B.n80 71.676
R1064 B.n172 B.n81 71.676
R1065 B.n176 B.n82 71.676
R1066 B.n180 B.n83 71.676
R1067 B.n84 B.n83 71.676
R1068 B.n179 B.n82 71.676
R1069 B.n175 B.n81 71.676
R1070 B.n171 B.n80 71.676
R1071 B.n167 B.n79 71.676
R1072 B.n163 B.n78 71.676
R1073 B.n159 B.n77 71.676
R1074 B.n155 B.n76 71.676
R1075 B.n151 B.n75 71.676
R1076 B.n147 B.n74 71.676
R1077 B.n142 B.n73 71.676
R1078 B.n138 B.n72 71.676
R1079 B.n134 B.n71 71.676
R1080 B.n130 B.n70 71.676
R1081 B.n126 B.n69 71.676
R1082 B.n122 B.n68 71.676
R1083 B.n118 B.n67 71.676
R1084 B.n114 B.n66 71.676
R1085 B.n110 B.n65 71.676
R1086 B.n106 B.n64 71.676
R1087 B.n102 B.n63 71.676
R1088 B.n98 B.n62 71.676
R1089 B.n94 B.n61 71.676
R1090 B.n506 B.n60 71.676
R1091 B.n369 B.n244 71.676
R1092 B.n363 B.n245 71.676
R1093 B.n359 B.n246 71.676
R1094 B.n355 B.n247 71.676
R1095 B.n351 B.n248 71.676
R1096 B.n347 B.n249 71.676
R1097 B.n343 B.n250 71.676
R1098 B.n339 B.n251 71.676
R1099 B.n335 B.n252 71.676
R1100 B.n330 B.n253 71.676
R1101 B.n326 B.n254 71.676
R1102 B.n322 B.n255 71.676
R1103 B.n318 B.n256 71.676
R1104 B.n314 B.n257 71.676
R1105 B.n310 B.n258 71.676
R1106 B.n306 B.n259 71.676
R1107 B.n302 B.n260 71.676
R1108 B.n298 B.n261 71.676
R1109 B.n294 B.n262 71.676
R1110 B.n290 B.n263 71.676
R1111 B.n286 B.n264 71.676
R1112 B.n282 B.n265 71.676
R1113 B.n278 B.n266 71.676
R1114 B.n274 B.n267 71.676
R1115 B.t2 B.n185 68.8546
R1116 B.t5 B.n8 68.8546
R1117 B.n423 B.t0 64.4124
R1118 B.t3 B.n544 64.4124
R1119 B.n273 B.n272 59.5399
R1120 B.n332 B.n270 59.5399
R1121 B.n90 B.n89 59.5399
R1122 B.n145 B.n87 59.5399
R1123 B.t4 B.n213 57.7491
R1124 B.n537 B.t6 57.7491
R1125 B.t9 B.n229 44.4225
R1126 B.n521 B.t16 44.4225
R1127 B.n441 B.t1 39.9803
R1128 B.n554 B.t7 39.9803
R1129 B.n509 B.n508 36.9956
R1130 B.n503 B.n502 36.9956
R1131 B.n275 B.n239 36.9956
R1132 B.n372 B.n371 36.9956
R1133 B.n201 B.t1 35.5381
R1134 B.t7 B.n553 35.5381
R1135 B.n387 B.t9 31.0959
R1136 B.t16 B.n520 31.0959
R1137 B.n272 B.n271 30.449
R1138 B.n270 B.n269 30.449
R1139 B.n89 B.n88 30.449
R1140 B.n87 B.n86 30.449
R1141 B B.n572 18.0485
R1142 B.n411 B.t4 17.7693
R1143 B.t6 B.n536 17.7693
R1144 B.t0 B.n205 11.106
R1145 B.n545 B.t3 11.106
R1146 B.n508 B.n59 10.6151
R1147 B.n92 B.n59 10.6151
R1148 B.n93 B.n92 10.6151
R1149 B.n96 B.n93 10.6151
R1150 B.n97 B.n96 10.6151
R1151 B.n100 B.n97 10.6151
R1152 B.n101 B.n100 10.6151
R1153 B.n104 B.n101 10.6151
R1154 B.n105 B.n104 10.6151
R1155 B.n108 B.n105 10.6151
R1156 B.n109 B.n108 10.6151
R1157 B.n112 B.n109 10.6151
R1158 B.n113 B.n112 10.6151
R1159 B.n116 B.n113 10.6151
R1160 B.n117 B.n116 10.6151
R1161 B.n120 B.n117 10.6151
R1162 B.n121 B.n120 10.6151
R1163 B.n124 B.n121 10.6151
R1164 B.n125 B.n124 10.6151
R1165 B.n129 B.n128 10.6151
R1166 B.n132 B.n129 10.6151
R1167 B.n133 B.n132 10.6151
R1168 B.n136 B.n133 10.6151
R1169 B.n137 B.n136 10.6151
R1170 B.n140 B.n137 10.6151
R1171 B.n141 B.n140 10.6151
R1172 B.n144 B.n141 10.6151
R1173 B.n149 B.n146 10.6151
R1174 B.n150 B.n149 10.6151
R1175 B.n153 B.n150 10.6151
R1176 B.n154 B.n153 10.6151
R1177 B.n157 B.n154 10.6151
R1178 B.n158 B.n157 10.6151
R1179 B.n161 B.n158 10.6151
R1180 B.n162 B.n161 10.6151
R1181 B.n165 B.n162 10.6151
R1182 B.n166 B.n165 10.6151
R1183 B.n169 B.n166 10.6151
R1184 B.n170 B.n169 10.6151
R1185 B.n173 B.n170 10.6151
R1186 B.n174 B.n173 10.6151
R1187 B.n177 B.n174 10.6151
R1188 B.n178 B.n177 10.6151
R1189 B.n181 B.n178 10.6151
R1190 B.n182 B.n181 10.6151
R1191 B.n503 B.n182 10.6151
R1192 B.n377 B.n239 10.6151
R1193 B.n378 B.n377 10.6151
R1194 B.n379 B.n378 10.6151
R1195 B.n379 B.n231 10.6151
R1196 B.n389 B.n231 10.6151
R1197 B.n390 B.n389 10.6151
R1198 B.n391 B.n390 10.6151
R1199 B.n391 B.n223 10.6151
R1200 B.n401 B.n223 10.6151
R1201 B.n402 B.n401 10.6151
R1202 B.n403 B.n402 10.6151
R1203 B.n403 B.n215 10.6151
R1204 B.n413 B.n215 10.6151
R1205 B.n414 B.n413 10.6151
R1206 B.n415 B.n414 10.6151
R1207 B.n415 B.n207 10.6151
R1208 B.n425 B.n207 10.6151
R1209 B.n426 B.n425 10.6151
R1210 B.n427 B.n426 10.6151
R1211 B.n427 B.n198 10.6151
R1212 B.n437 B.n198 10.6151
R1213 B.n438 B.n437 10.6151
R1214 B.n439 B.n438 10.6151
R1215 B.n439 B.n191 10.6151
R1216 B.n449 B.n191 10.6151
R1217 B.n450 B.n449 10.6151
R1218 B.n452 B.n450 10.6151
R1219 B.n452 B.n451 10.6151
R1220 B.n451 B.n183 10.6151
R1221 B.n463 B.n183 10.6151
R1222 B.n464 B.n463 10.6151
R1223 B.n465 B.n464 10.6151
R1224 B.n466 B.n465 10.6151
R1225 B.n468 B.n466 10.6151
R1226 B.n469 B.n468 10.6151
R1227 B.n470 B.n469 10.6151
R1228 B.n471 B.n470 10.6151
R1229 B.n473 B.n471 10.6151
R1230 B.n474 B.n473 10.6151
R1231 B.n475 B.n474 10.6151
R1232 B.n476 B.n475 10.6151
R1233 B.n478 B.n476 10.6151
R1234 B.n479 B.n478 10.6151
R1235 B.n480 B.n479 10.6151
R1236 B.n481 B.n480 10.6151
R1237 B.n483 B.n481 10.6151
R1238 B.n484 B.n483 10.6151
R1239 B.n485 B.n484 10.6151
R1240 B.n486 B.n485 10.6151
R1241 B.n488 B.n486 10.6151
R1242 B.n489 B.n488 10.6151
R1243 B.n490 B.n489 10.6151
R1244 B.n491 B.n490 10.6151
R1245 B.n493 B.n491 10.6151
R1246 B.n494 B.n493 10.6151
R1247 B.n495 B.n494 10.6151
R1248 B.n496 B.n495 10.6151
R1249 B.n498 B.n496 10.6151
R1250 B.n499 B.n498 10.6151
R1251 B.n500 B.n499 10.6151
R1252 B.n501 B.n500 10.6151
R1253 B.n502 B.n501 10.6151
R1254 B.n371 B.n243 10.6151
R1255 B.n366 B.n243 10.6151
R1256 B.n366 B.n365 10.6151
R1257 B.n365 B.n364 10.6151
R1258 B.n364 B.n361 10.6151
R1259 B.n361 B.n360 10.6151
R1260 B.n360 B.n357 10.6151
R1261 B.n357 B.n356 10.6151
R1262 B.n356 B.n353 10.6151
R1263 B.n353 B.n352 10.6151
R1264 B.n352 B.n349 10.6151
R1265 B.n349 B.n348 10.6151
R1266 B.n348 B.n345 10.6151
R1267 B.n345 B.n344 10.6151
R1268 B.n344 B.n341 10.6151
R1269 B.n341 B.n340 10.6151
R1270 B.n340 B.n337 10.6151
R1271 B.n337 B.n336 10.6151
R1272 B.n336 B.n333 10.6151
R1273 B.n331 B.n328 10.6151
R1274 B.n328 B.n327 10.6151
R1275 B.n327 B.n324 10.6151
R1276 B.n324 B.n323 10.6151
R1277 B.n323 B.n320 10.6151
R1278 B.n320 B.n319 10.6151
R1279 B.n319 B.n316 10.6151
R1280 B.n316 B.n315 10.6151
R1281 B.n312 B.n311 10.6151
R1282 B.n311 B.n308 10.6151
R1283 B.n308 B.n307 10.6151
R1284 B.n307 B.n304 10.6151
R1285 B.n304 B.n303 10.6151
R1286 B.n303 B.n300 10.6151
R1287 B.n300 B.n299 10.6151
R1288 B.n299 B.n296 10.6151
R1289 B.n296 B.n295 10.6151
R1290 B.n295 B.n292 10.6151
R1291 B.n292 B.n291 10.6151
R1292 B.n291 B.n288 10.6151
R1293 B.n288 B.n287 10.6151
R1294 B.n287 B.n284 10.6151
R1295 B.n284 B.n283 10.6151
R1296 B.n283 B.n280 10.6151
R1297 B.n280 B.n279 10.6151
R1298 B.n279 B.n276 10.6151
R1299 B.n276 B.n275 10.6151
R1300 B.n373 B.n372 10.6151
R1301 B.n373 B.n235 10.6151
R1302 B.n383 B.n235 10.6151
R1303 B.n384 B.n383 10.6151
R1304 B.n385 B.n384 10.6151
R1305 B.n385 B.n227 10.6151
R1306 B.n395 B.n227 10.6151
R1307 B.n396 B.n395 10.6151
R1308 B.n397 B.n396 10.6151
R1309 B.n397 B.n219 10.6151
R1310 B.n407 B.n219 10.6151
R1311 B.n408 B.n407 10.6151
R1312 B.n409 B.n408 10.6151
R1313 B.n409 B.n211 10.6151
R1314 B.n419 B.n211 10.6151
R1315 B.n420 B.n419 10.6151
R1316 B.n421 B.n420 10.6151
R1317 B.n421 B.n203 10.6151
R1318 B.n431 B.n203 10.6151
R1319 B.n432 B.n431 10.6151
R1320 B.n433 B.n432 10.6151
R1321 B.n433 B.n195 10.6151
R1322 B.n443 B.n195 10.6151
R1323 B.n444 B.n443 10.6151
R1324 B.n445 B.n444 10.6151
R1325 B.n445 B.n187 10.6151
R1326 B.n456 B.n187 10.6151
R1327 B.n457 B.n456 10.6151
R1328 B.n458 B.n457 10.6151
R1329 B.n458 B.n0 10.6151
R1330 B.n566 B.n1 10.6151
R1331 B.n566 B.n565 10.6151
R1332 B.n565 B.n564 10.6151
R1333 B.n564 B.n10 10.6151
R1334 B.n558 B.n10 10.6151
R1335 B.n558 B.n557 10.6151
R1336 B.n557 B.n556 10.6151
R1337 B.n556 B.n17 10.6151
R1338 B.n550 B.n17 10.6151
R1339 B.n550 B.n549 10.6151
R1340 B.n549 B.n548 10.6151
R1341 B.n548 B.n24 10.6151
R1342 B.n542 B.n24 10.6151
R1343 B.n542 B.n541 10.6151
R1344 B.n541 B.n540 10.6151
R1345 B.n540 B.n31 10.6151
R1346 B.n534 B.n31 10.6151
R1347 B.n534 B.n533 10.6151
R1348 B.n533 B.n532 10.6151
R1349 B.n532 B.n38 10.6151
R1350 B.n526 B.n38 10.6151
R1351 B.n526 B.n525 10.6151
R1352 B.n525 B.n524 10.6151
R1353 B.n524 B.n45 10.6151
R1354 B.n518 B.n45 10.6151
R1355 B.n518 B.n517 10.6151
R1356 B.n517 B.n516 10.6151
R1357 B.n516 B.n52 10.6151
R1358 B.n510 B.n52 10.6151
R1359 B.n510 B.n509 10.6151
R1360 B.n454 B.t2 6.6638
R1361 B.n562 B.t5 6.6638
R1362 B.n128 B.n90 6.5566
R1363 B.n145 B.n144 6.5566
R1364 B.n332 B.n331 6.5566
R1365 B.n315 B.n273 6.5566
R1366 B.n125 B.n90 4.05904
R1367 B.n146 B.n145 4.05904
R1368 B.n333 B.n332 4.05904
R1369 B.n312 B.n273 4.05904
R1370 B.n572 B.n0 2.81026
R1371 B.n572 B.n1 2.81026
R1372 VP.n11 VP.n10 161.3
R1373 VP.n12 VP.n7 161.3
R1374 VP.n14 VP.n13 161.3
R1375 VP.n16 VP.n15 161.3
R1376 VP.n17 VP.n5 161.3
R1377 VP.n32 VP.n0 161.3
R1378 VP.n31 VP.n30 161.3
R1379 VP.n29 VP.n28 161.3
R1380 VP.n27 VP.n2 161.3
R1381 VP.n26 VP.n25 161.3
R1382 VP.n24 VP.n23 161.3
R1383 VP.n22 VP.n4 161.3
R1384 VP.n9 VP.t4 141.601
R1385 VP.n21 VP.t5 121.861
R1386 VP.n33 VP.t7 121.861
R1387 VP.n18 VP.t0 121.861
R1388 VP.n3 VP.t3 89.9868
R1389 VP.n1 VP.t2 89.9868
R1390 VP.n6 VP.t6 89.9868
R1391 VP.n8 VP.t1 89.9868
R1392 VP.n19 VP.n18 80.6037
R1393 VP.n34 VP.n33 80.6037
R1394 VP.n21 VP.n20 80.6037
R1395 VP.n9 VP.n8 43.5433
R1396 VP.n27 VP.n26 40.4934
R1397 VP.n28 VP.n27 40.4934
R1398 VP.n13 VP.n12 40.4934
R1399 VP.n12 VP.n11 40.4934
R1400 VP.n20 VP.n19 39.115
R1401 VP.n22 VP.n21 34.3247
R1402 VP.n33 VP.n32 34.3247
R1403 VP.n18 VP.n17 34.3247
R1404 VP.n23 VP.n22 33.6945
R1405 VP.n32 VP.n31 33.6945
R1406 VP.n17 VP.n16 33.6945
R1407 VP.n10 VP.n9 29.3131
R1408 VP.n26 VP.n3 13.9467
R1409 VP.n28 VP.n1 13.9467
R1410 VP.n13 VP.n6 13.9467
R1411 VP.n11 VP.n8 13.9467
R1412 VP.n23 VP.n3 10.5213
R1413 VP.n31 VP.n1 10.5213
R1414 VP.n16 VP.n6 10.5213
R1415 VP.n19 VP.n5 0.285035
R1416 VP.n20 VP.n4 0.285035
R1417 VP.n34 VP.n0 0.285035
R1418 VP.n10 VP.n7 0.189894
R1419 VP.n14 VP.n7 0.189894
R1420 VP.n15 VP.n14 0.189894
R1421 VP.n15 VP.n5 0.189894
R1422 VP.n24 VP.n4 0.189894
R1423 VP.n25 VP.n24 0.189894
R1424 VP.n25 VP.n2 0.189894
R1425 VP.n29 VP.n2 0.189894
R1426 VP.n30 VP.n29 0.189894
R1427 VP.n30 VP.n0 0.189894
R1428 VP VP.n34 0.146778
R1429 VDD1 VDD1.n0 72.7343
R1430 VDD1.n3 VDD1.n2 72.6206
R1431 VDD1.n3 VDD1.n1 72.6206
R1432 VDD1.n5 VDD1.n4 71.9992
R1433 VDD1.n5 VDD1.n3 34.3802
R1434 VDD1.n4 VDD1.t1 4.27696
R1435 VDD1.n4 VDD1.t7 4.27696
R1436 VDD1.n0 VDD1.t3 4.27696
R1437 VDD1.n0 VDD1.t6 4.27696
R1438 VDD1.n2 VDD1.t5 4.27696
R1439 VDD1.n2 VDD1.t0 4.27696
R1440 VDD1.n1 VDD1.t2 4.27696
R1441 VDD1.n1 VDD1.t4 4.27696
R1442 VDD1 VDD1.n5 0.619035
C0 VDD1 VDD2 1.09481f
C1 VP VDD1 3.21779f
C2 VTAIL VDD1 5.06528f
C3 VP VDD2 0.378989f
C4 VTAIL VDD2 5.11058f
C5 VN VDD1 0.152943f
C6 VTAIL VP 3.36099f
C7 VN VDD2 2.99286f
C8 VN VP 4.63336f
C9 VN VTAIL 3.34689f
C10 VDD2 B 3.416244f
C11 VDD1 B 3.711509f
C12 VTAIL B 4.942329f
C13 VN B 9.61953f
C14 VP B 8.139984f
C15 VDD1.t3 B 0.092931f
C16 VDD1.t6 B 0.092931f
C17 VDD1.n0 B 0.752048f
C18 VDD1.t2 B 0.092931f
C19 VDD1.t4 B 0.092931f
C20 VDD1.n1 B 0.751382f
C21 VDD1.t5 B 0.092931f
C22 VDD1.t0 B 0.092931f
C23 VDD1.n2 B 0.751382f
C24 VDD1.n3 B 2.11518f
C25 VDD1.t1 B 0.092931f
C26 VDD1.t7 B 0.092931f
C27 VDD1.n4 B 0.748186f
C28 VDD1.n5 B 1.94961f
C29 VP.n0 B 0.050528f
C30 VP.t2 B 0.565392f
C31 VP.n1 B 0.237924f
C32 VP.n2 B 0.037867f
C33 VP.t3 B 0.565392f
C34 VP.n3 B 0.237924f
C35 VP.n4 B 0.050528f
C36 VP.n5 B 0.050528f
C37 VP.t0 B 0.637327f
C38 VP.t6 B 0.565392f
C39 VP.n6 B 0.237924f
C40 VP.n7 B 0.037867f
C41 VP.t1 B 0.565392f
C42 VP.n8 B 0.288357f
C43 VP.t4 B 0.681924f
C44 VP.n9 B 0.301119f
C45 VP.n10 B 0.198043f
C46 VP.n11 B 0.060275f
C47 VP.n12 B 0.030612f
C48 VP.n13 B 0.060275f
C49 VP.n14 B 0.037867f
C50 VP.n15 B 0.037867f
C51 VP.n16 B 0.056625f
C52 VP.n17 B 0.026496f
C53 VP.n18 B 0.311232f
C54 VP.n19 B 1.39748f
C55 VP.n20 B 1.43228f
C56 VP.t5 B 0.637327f
C57 VP.n21 B 0.311232f
C58 VP.n22 B 0.026496f
C59 VP.n23 B 0.056625f
C60 VP.n24 B 0.037867f
C61 VP.n25 B 0.037867f
C62 VP.n26 B 0.060275f
C63 VP.n27 B 0.030612f
C64 VP.n28 B 0.060275f
C65 VP.n29 B 0.037867f
C66 VP.n30 B 0.037867f
C67 VP.n31 B 0.056625f
C68 VP.n32 B 0.026496f
C69 VP.t7 B 0.637327f
C70 VP.n33 B 0.311232f
C71 VP.n34 B 0.035464f
C72 VDD2.t1 B 0.091729f
C73 VDD2.t7 B 0.091729f
C74 VDD2.n0 B 0.74166f
C75 VDD2.t5 B 0.091729f
C76 VDD2.t3 B 0.091729f
C77 VDD2.n1 B 0.74166f
C78 VDD2.n2 B 2.03449f
C79 VDD2.t4 B 0.091729f
C80 VDD2.t0 B 0.091729f
C81 VDD2.n3 B 0.738509f
C82 VDD2.n4 B 1.8945f
C83 VDD2.t6 B 0.091729f
C84 VDD2.t2 B 0.091729f
C85 VDD2.n5 B 0.741635f
C86 VTAIL.t9 B 0.083542f
C87 VTAIL.t8 B 0.083542f
C88 VTAIL.n0 B 0.619507f
C89 VTAIL.n1 B 0.306334f
C90 VTAIL.n2 B 0.03194f
C91 VTAIL.n3 B 0.022833f
C92 VTAIL.n4 B 0.01227f
C93 VTAIL.n5 B 0.029001f
C94 VTAIL.n6 B 0.012991f
C95 VTAIL.n7 B 0.39865f
C96 VTAIL.n8 B 0.01227f
C97 VTAIL.t6 B 0.047616f
C98 VTAIL.n9 B 0.090712f
C99 VTAIL.n10 B 0.017115f
C100 VTAIL.n11 B 0.021751f
C101 VTAIL.n12 B 0.029001f
C102 VTAIL.n13 B 0.012991f
C103 VTAIL.n14 B 0.01227f
C104 VTAIL.n15 B 0.022833f
C105 VTAIL.n16 B 0.022833f
C106 VTAIL.n17 B 0.01227f
C107 VTAIL.n18 B 0.012991f
C108 VTAIL.n19 B 0.029001f
C109 VTAIL.n20 B 0.06251f
C110 VTAIL.n21 B 0.012991f
C111 VTAIL.n22 B 0.01227f
C112 VTAIL.n23 B 0.054962f
C113 VTAIL.n24 B 0.035015f
C114 VTAIL.n25 B 0.154881f
C115 VTAIL.n26 B 0.03194f
C116 VTAIL.n27 B 0.022833f
C117 VTAIL.n28 B 0.01227f
C118 VTAIL.n29 B 0.029001f
C119 VTAIL.n30 B 0.012991f
C120 VTAIL.n31 B 0.39865f
C121 VTAIL.n32 B 0.01227f
C122 VTAIL.t2 B 0.047616f
C123 VTAIL.n33 B 0.090712f
C124 VTAIL.n34 B 0.017115f
C125 VTAIL.n35 B 0.021751f
C126 VTAIL.n36 B 0.029001f
C127 VTAIL.n37 B 0.012991f
C128 VTAIL.n38 B 0.01227f
C129 VTAIL.n39 B 0.022833f
C130 VTAIL.n40 B 0.022833f
C131 VTAIL.n41 B 0.01227f
C132 VTAIL.n42 B 0.012991f
C133 VTAIL.n43 B 0.029001f
C134 VTAIL.n44 B 0.06251f
C135 VTAIL.n45 B 0.012991f
C136 VTAIL.n46 B 0.01227f
C137 VTAIL.n47 B 0.054962f
C138 VTAIL.n48 B 0.035015f
C139 VTAIL.n49 B 0.154881f
C140 VTAIL.t0 B 0.083542f
C141 VTAIL.t1 B 0.083542f
C142 VTAIL.n50 B 0.619507f
C143 VTAIL.n51 B 0.401632f
C144 VTAIL.n52 B 0.03194f
C145 VTAIL.n53 B 0.022833f
C146 VTAIL.n54 B 0.01227f
C147 VTAIL.n55 B 0.029001f
C148 VTAIL.n56 B 0.012991f
C149 VTAIL.n57 B 0.39865f
C150 VTAIL.n58 B 0.01227f
C151 VTAIL.t4 B 0.047616f
C152 VTAIL.n59 B 0.090712f
C153 VTAIL.n60 B 0.017115f
C154 VTAIL.n61 B 0.021751f
C155 VTAIL.n62 B 0.029001f
C156 VTAIL.n63 B 0.012991f
C157 VTAIL.n64 B 0.01227f
C158 VTAIL.n65 B 0.022833f
C159 VTAIL.n66 B 0.022833f
C160 VTAIL.n67 B 0.01227f
C161 VTAIL.n68 B 0.012991f
C162 VTAIL.n69 B 0.029001f
C163 VTAIL.n70 B 0.06251f
C164 VTAIL.n71 B 0.012991f
C165 VTAIL.n72 B 0.01227f
C166 VTAIL.n73 B 0.054962f
C167 VTAIL.n74 B 0.035015f
C168 VTAIL.n75 B 0.82372f
C169 VTAIL.n76 B 0.03194f
C170 VTAIL.n77 B 0.022833f
C171 VTAIL.n78 B 0.01227f
C172 VTAIL.n79 B 0.029001f
C173 VTAIL.n80 B 0.012991f
C174 VTAIL.n81 B 0.39865f
C175 VTAIL.n82 B 0.01227f
C176 VTAIL.t11 B 0.047616f
C177 VTAIL.n83 B 0.090712f
C178 VTAIL.n84 B 0.017115f
C179 VTAIL.n85 B 0.021751f
C180 VTAIL.n86 B 0.029001f
C181 VTAIL.n87 B 0.012991f
C182 VTAIL.n88 B 0.01227f
C183 VTAIL.n89 B 0.022833f
C184 VTAIL.n90 B 0.022833f
C185 VTAIL.n91 B 0.01227f
C186 VTAIL.n92 B 0.012991f
C187 VTAIL.n93 B 0.029001f
C188 VTAIL.n94 B 0.06251f
C189 VTAIL.n95 B 0.012991f
C190 VTAIL.n96 B 0.01227f
C191 VTAIL.n97 B 0.054962f
C192 VTAIL.n98 B 0.035015f
C193 VTAIL.n99 B 0.82372f
C194 VTAIL.t5 B 0.083542f
C195 VTAIL.t12 B 0.083542f
C196 VTAIL.n100 B 0.619511f
C197 VTAIL.n101 B 0.401628f
C198 VTAIL.n102 B 0.03194f
C199 VTAIL.n103 B 0.022833f
C200 VTAIL.n104 B 0.01227f
C201 VTAIL.n105 B 0.029001f
C202 VTAIL.n106 B 0.012991f
C203 VTAIL.n107 B 0.39865f
C204 VTAIL.n108 B 0.01227f
C205 VTAIL.t7 B 0.047616f
C206 VTAIL.n109 B 0.090712f
C207 VTAIL.n110 B 0.017115f
C208 VTAIL.n111 B 0.021751f
C209 VTAIL.n112 B 0.029001f
C210 VTAIL.n113 B 0.012991f
C211 VTAIL.n114 B 0.01227f
C212 VTAIL.n115 B 0.022833f
C213 VTAIL.n116 B 0.022833f
C214 VTAIL.n117 B 0.01227f
C215 VTAIL.n118 B 0.012991f
C216 VTAIL.n119 B 0.029001f
C217 VTAIL.n120 B 0.06251f
C218 VTAIL.n121 B 0.012991f
C219 VTAIL.n122 B 0.01227f
C220 VTAIL.n123 B 0.054962f
C221 VTAIL.n124 B 0.035015f
C222 VTAIL.n125 B 0.154881f
C223 VTAIL.n126 B 0.03194f
C224 VTAIL.n127 B 0.022833f
C225 VTAIL.n128 B 0.01227f
C226 VTAIL.n129 B 0.029001f
C227 VTAIL.n130 B 0.012991f
C228 VTAIL.n131 B 0.39865f
C229 VTAIL.n132 B 0.01227f
C230 VTAIL.t13 B 0.047616f
C231 VTAIL.n133 B 0.090712f
C232 VTAIL.n134 B 0.017115f
C233 VTAIL.n135 B 0.021751f
C234 VTAIL.n136 B 0.029001f
C235 VTAIL.n137 B 0.012991f
C236 VTAIL.n138 B 0.01227f
C237 VTAIL.n139 B 0.022833f
C238 VTAIL.n140 B 0.022833f
C239 VTAIL.n141 B 0.01227f
C240 VTAIL.n142 B 0.012991f
C241 VTAIL.n143 B 0.029001f
C242 VTAIL.n144 B 0.06251f
C243 VTAIL.n145 B 0.012991f
C244 VTAIL.n146 B 0.01227f
C245 VTAIL.n147 B 0.054962f
C246 VTAIL.n148 B 0.035015f
C247 VTAIL.n149 B 0.154881f
C248 VTAIL.t14 B 0.083542f
C249 VTAIL.t3 B 0.083542f
C250 VTAIL.n150 B 0.619511f
C251 VTAIL.n151 B 0.401628f
C252 VTAIL.n152 B 0.03194f
C253 VTAIL.n153 B 0.022833f
C254 VTAIL.n154 B 0.01227f
C255 VTAIL.n155 B 0.029001f
C256 VTAIL.n156 B 0.012991f
C257 VTAIL.n157 B 0.39865f
C258 VTAIL.n158 B 0.01227f
C259 VTAIL.t15 B 0.047616f
C260 VTAIL.n159 B 0.090712f
C261 VTAIL.n160 B 0.017115f
C262 VTAIL.n161 B 0.021751f
C263 VTAIL.n162 B 0.029001f
C264 VTAIL.n163 B 0.012991f
C265 VTAIL.n164 B 0.01227f
C266 VTAIL.n165 B 0.022833f
C267 VTAIL.n166 B 0.022833f
C268 VTAIL.n167 B 0.01227f
C269 VTAIL.n168 B 0.012991f
C270 VTAIL.n169 B 0.029001f
C271 VTAIL.n170 B 0.06251f
C272 VTAIL.n171 B 0.012991f
C273 VTAIL.n172 B 0.01227f
C274 VTAIL.n173 B 0.054962f
C275 VTAIL.n174 B 0.035015f
C276 VTAIL.n175 B 0.82372f
C277 VTAIL.n176 B 0.03194f
C278 VTAIL.n177 B 0.022833f
C279 VTAIL.n178 B 0.01227f
C280 VTAIL.n179 B 0.029001f
C281 VTAIL.n180 B 0.012991f
C282 VTAIL.n181 B 0.39865f
C283 VTAIL.n182 B 0.01227f
C284 VTAIL.t10 B 0.047616f
C285 VTAIL.n183 B 0.090712f
C286 VTAIL.n184 B 0.017115f
C287 VTAIL.n185 B 0.021751f
C288 VTAIL.n186 B 0.029001f
C289 VTAIL.n187 B 0.012991f
C290 VTAIL.n188 B 0.01227f
C291 VTAIL.n189 B 0.022833f
C292 VTAIL.n190 B 0.022833f
C293 VTAIL.n191 B 0.01227f
C294 VTAIL.n192 B 0.012991f
C295 VTAIL.n193 B 0.029001f
C296 VTAIL.n194 B 0.06251f
C297 VTAIL.n195 B 0.012991f
C298 VTAIL.n196 B 0.01227f
C299 VTAIL.n197 B 0.054962f
C300 VTAIL.n198 B 0.035015f
C301 VTAIL.n199 B 0.819439f
C302 VN.n0 B 0.048942f
C303 VN.t2 B 0.547644f
C304 VN.n1 B 0.230456f
C305 VN.n2 B 0.036678f
C306 VN.t0 B 0.547644f
C307 VN.n3 B 0.279306f
C308 VN.t6 B 0.660519f
C309 VN.n4 B 0.291667f
C310 VN.n5 B 0.191826f
C311 VN.n6 B 0.058383f
C312 VN.n7 B 0.029651f
C313 VN.n8 B 0.058383f
C314 VN.n9 B 0.036678f
C315 VN.n10 B 0.036678f
C316 VN.n11 B 0.054848f
C317 VN.n12 B 0.025664f
C318 VN.t4 B 0.617321f
C319 VN.n13 B 0.301463f
C320 VN.n14 B 0.03435f
C321 VN.n15 B 0.048942f
C322 VN.t7 B 0.547644f
C323 VN.n16 B 0.230456f
C324 VN.n17 B 0.036678f
C325 VN.t1 B 0.547644f
C326 VN.n18 B 0.279306f
C327 VN.t5 B 0.660519f
C328 VN.n19 B 0.291667f
C329 VN.n20 B 0.191826f
C330 VN.n21 B 0.058383f
C331 VN.n22 B 0.029651f
C332 VN.n23 B 0.058383f
C333 VN.n24 B 0.036678f
C334 VN.n25 B 0.036678f
C335 VN.n26 B 0.054848f
C336 VN.n27 B 0.025664f
C337 VN.t3 B 0.617321f
C338 VN.n28 B 0.301463f
C339 VN.n29 B 1.37446f
.ends

