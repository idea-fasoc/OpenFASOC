* NGSPICE file created from diff_pair_sample_0035.ext - technology: sky130A

.subckt diff_pair_sample_0035 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=2.72
X1 VTAIL.t15 VP.t0 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=2.72
X2 VTAIL.t1 VN.t0 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=2.72
X3 VTAIL.t2 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X4 VDD2.t5 VN.t2 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X5 VDD1.t1 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=2.72
X6 VDD1.t6 VP.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=2.72
X7 VTAIL.t4 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=2.72
X8 VDD1.t0 VP.t3 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X9 VTAIL.t6 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X10 VDD2.t2 VN.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X11 VTAIL.t11 VP.t4 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X12 VDD2.t1 VN.t6 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=2.72
X13 VTAIL.t10 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=2.72
X14 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=2.72
X15 VTAIL.t9 VP.t6 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X16 VDD1.t5 VP.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=2.72
X17 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=2.72
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=2.72
X19 VDD2.t0 VN.t7 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=2.72
R0 B.n596 B.n595 585
R1 B.n180 B.n113 585
R2 B.n179 B.n178 585
R3 B.n177 B.n176 585
R4 B.n175 B.n174 585
R5 B.n173 B.n172 585
R6 B.n171 B.n170 585
R7 B.n169 B.n168 585
R8 B.n167 B.n166 585
R9 B.n165 B.n164 585
R10 B.n163 B.n162 585
R11 B.n160 B.n159 585
R12 B.n158 B.n157 585
R13 B.n156 B.n155 585
R14 B.n154 B.n153 585
R15 B.n152 B.n151 585
R16 B.n150 B.n149 585
R17 B.n148 B.n147 585
R18 B.n146 B.n145 585
R19 B.n144 B.n143 585
R20 B.n142 B.n141 585
R21 B.n139 B.n138 585
R22 B.n137 B.n136 585
R23 B.n135 B.n134 585
R24 B.n133 B.n132 585
R25 B.n131 B.n130 585
R26 B.n129 B.n128 585
R27 B.n127 B.n126 585
R28 B.n125 B.n124 585
R29 B.n123 B.n122 585
R30 B.n121 B.n120 585
R31 B.n119 B.n118 585
R32 B.n594 B.n97 585
R33 B.n599 B.n97 585
R34 B.n593 B.n96 585
R35 B.n600 B.n96 585
R36 B.n592 B.n591 585
R37 B.n591 B.n92 585
R38 B.n590 B.n91 585
R39 B.n606 B.n91 585
R40 B.n589 B.n90 585
R41 B.n607 B.n90 585
R42 B.n588 B.n89 585
R43 B.n608 B.n89 585
R44 B.n587 B.n586 585
R45 B.n586 B.n85 585
R46 B.n585 B.n84 585
R47 B.n614 B.n84 585
R48 B.n584 B.n83 585
R49 B.n615 B.n83 585
R50 B.n583 B.n82 585
R51 B.n616 B.n82 585
R52 B.n582 B.n581 585
R53 B.n581 B.n78 585
R54 B.n580 B.n77 585
R55 B.n622 B.n77 585
R56 B.n579 B.n76 585
R57 B.n623 B.n76 585
R58 B.n578 B.n75 585
R59 B.n624 B.n75 585
R60 B.n577 B.n576 585
R61 B.n576 B.n71 585
R62 B.n575 B.n70 585
R63 B.n630 B.n70 585
R64 B.n574 B.n69 585
R65 B.n631 B.n69 585
R66 B.n573 B.n68 585
R67 B.n632 B.n68 585
R68 B.n572 B.n571 585
R69 B.n571 B.n64 585
R70 B.n570 B.n63 585
R71 B.n638 B.n63 585
R72 B.n569 B.n62 585
R73 B.t3 B.n62 585
R74 B.n568 B.n61 585
R75 B.n639 B.n61 585
R76 B.n567 B.n566 585
R77 B.n566 B.n57 585
R78 B.n565 B.n56 585
R79 B.n645 B.n56 585
R80 B.n564 B.n55 585
R81 B.n646 B.n55 585
R82 B.n563 B.n54 585
R83 B.n647 B.n54 585
R84 B.n562 B.n561 585
R85 B.n561 B.n50 585
R86 B.n560 B.n49 585
R87 B.n653 B.n49 585
R88 B.n559 B.n48 585
R89 B.n654 B.n48 585
R90 B.n558 B.n47 585
R91 B.n655 B.n47 585
R92 B.n557 B.n556 585
R93 B.n556 B.n43 585
R94 B.n555 B.n42 585
R95 B.n661 B.n42 585
R96 B.n554 B.n41 585
R97 B.n662 B.n41 585
R98 B.n553 B.n40 585
R99 B.n663 B.n40 585
R100 B.n552 B.n551 585
R101 B.n551 B.n36 585
R102 B.n550 B.n35 585
R103 B.n669 B.n35 585
R104 B.n549 B.n34 585
R105 B.n670 B.n34 585
R106 B.n548 B.n33 585
R107 B.n671 B.n33 585
R108 B.n547 B.n546 585
R109 B.n546 B.n29 585
R110 B.n545 B.n28 585
R111 B.n677 B.n28 585
R112 B.n544 B.n27 585
R113 B.n678 B.n27 585
R114 B.n543 B.n26 585
R115 B.n679 B.n26 585
R116 B.n542 B.n541 585
R117 B.n541 B.n22 585
R118 B.n540 B.n21 585
R119 B.n685 B.n21 585
R120 B.n539 B.n20 585
R121 B.n686 B.n20 585
R122 B.n538 B.n19 585
R123 B.n687 B.n19 585
R124 B.n537 B.n536 585
R125 B.n536 B.n18 585
R126 B.n535 B.n14 585
R127 B.n693 B.n14 585
R128 B.n534 B.n13 585
R129 B.n694 B.n13 585
R130 B.n533 B.n12 585
R131 B.n695 B.n12 585
R132 B.n532 B.n531 585
R133 B.n531 B.n8 585
R134 B.n530 B.n7 585
R135 B.n701 B.n7 585
R136 B.n529 B.n6 585
R137 B.n702 B.n6 585
R138 B.n528 B.n5 585
R139 B.n703 B.n5 585
R140 B.n527 B.n526 585
R141 B.n526 B.n4 585
R142 B.n525 B.n181 585
R143 B.n525 B.n524 585
R144 B.n515 B.n182 585
R145 B.n183 B.n182 585
R146 B.n517 B.n516 585
R147 B.n518 B.n517 585
R148 B.n514 B.n188 585
R149 B.n188 B.n187 585
R150 B.n513 B.n512 585
R151 B.n512 B.n511 585
R152 B.n190 B.n189 585
R153 B.n504 B.n190 585
R154 B.n503 B.n502 585
R155 B.n505 B.n503 585
R156 B.n501 B.n195 585
R157 B.n195 B.n194 585
R158 B.n500 B.n499 585
R159 B.n499 B.n498 585
R160 B.n197 B.n196 585
R161 B.n198 B.n197 585
R162 B.n491 B.n490 585
R163 B.n492 B.n491 585
R164 B.n489 B.n203 585
R165 B.n203 B.n202 585
R166 B.n488 B.n487 585
R167 B.n487 B.n486 585
R168 B.n205 B.n204 585
R169 B.n206 B.n205 585
R170 B.n479 B.n478 585
R171 B.n480 B.n479 585
R172 B.n477 B.n211 585
R173 B.n211 B.n210 585
R174 B.n476 B.n475 585
R175 B.n475 B.n474 585
R176 B.n213 B.n212 585
R177 B.n214 B.n213 585
R178 B.n467 B.n466 585
R179 B.n468 B.n467 585
R180 B.n465 B.n219 585
R181 B.n219 B.n218 585
R182 B.n464 B.n463 585
R183 B.n463 B.n462 585
R184 B.n221 B.n220 585
R185 B.n222 B.n221 585
R186 B.n455 B.n454 585
R187 B.n456 B.n455 585
R188 B.n453 B.n226 585
R189 B.n230 B.n226 585
R190 B.n452 B.n451 585
R191 B.n451 B.n450 585
R192 B.n228 B.n227 585
R193 B.n229 B.n228 585
R194 B.n443 B.n442 585
R195 B.n444 B.n443 585
R196 B.n441 B.n235 585
R197 B.n235 B.n234 585
R198 B.n440 B.n439 585
R199 B.n439 B.n438 585
R200 B.n237 B.n236 585
R201 B.n238 B.n237 585
R202 B.n431 B.n430 585
R203 B.n432 B.n431 585
R204 B.n429 B.n242 585
R205 B.n242 B.t5 585
R206 B.n428 B.n427 585
R207 B.n427 B.n426 585
R208 B.n244 B.n243 585
R209 B.n245 B.n244 585
R210 B.n419 B.n418 585
R211 B.n420 B.n419 585
R212 B.n417 B.n250 585
R213 B.n250 B.n249 585
R214 B.n416 B.n415 585
R215 B.n415 B.n414 585
R216 B.n252 B.n251 585
R217 B.n253 B.n252 585
R218 B.n407 B.n406 585
R219 B.n408 B.n407 585
R220 B.n405 B.n258 585
R221 B.n258 B.n257 585
R222 B.n404 B.n403 585
R223 B.n403 B.n402 585
R224 B.n260 B.n259 585
R225 B.n261 B.n260 585
R226 B.n395 B.n394 585
R227 B.n396 B.n395 585
R228 B.n393 B.n266 585
R229 B.n266 B.n265 585
R230 B.n392 B.n391 585
R231 B.n391 B.n390 585
R232 B.n268 B.n267 585
R233 B.n269 B.n268 585
R234 B.n383 B.n382 585
R235 B.n384 B.n383 585
R236 B.n381 B.n274 585
R237 B.n274 B.n273 585
R238 B.n380 B.n379 585
R239 B.n379 B.n378 585
R240 B.n276 B.n275 585
R241 B.n277 B.n276 585
R242 B.n371 B.n370 585
R243 B.n372 B.n371 585
R244 B.n369 B.n282 585
R245 B.n282 B.n281 585
R246 B.n364 B.n363 585
R247 B.n362 B.n300 585
R248 B.n361 B.n299 585
R249 B.n366 B.n299 585
R250 B.n360 B.n359 585
R251 B.n358 B.n357 585
R252 B.n356 B.n355 585
R253 B.n354 B.n353 585
R254 B.n352 B.n351 585
R255 B.n350 B.n349 585
R256 B.n348 B.n347 585
R257 B.n346 B.n345 585
R258 B.n344 B.n343 585
R259 B.n342 B.n341 585
R260 B.n340 B.n339 585
R261 B.n338 B.n337 585
R262 B.n336 B.n335 585
R263 B.n334 B.n333 585
R264 B.n332 B.n331 585
R265 B.n330 B.n329 585
R266 B.n328 B.n327 585
R267 B.n326 B.n325 585
R268 B.n324 B.n323 585
R269 B.n322 B.n321 585
R270 B.n320 B.n319 585
R271 B.n318 B.n317 585
R272 B.n316 B.n315 585
R273 B.n314 B.n313 585
R274 B.n312 B.n311 585
R275 B.n310 B.n309 585
R276 B.n308 B.n307 585
R277 B.n284 B.n283 585
R278 B.n368 B.n367 585
R279 B.n367 B.n366 585
R280 B.n280 B.n279 585
R281 B.n281 B.n280 585
R282 B.n374 B.n373 585
R283 B.n373 B.n372 585
R284 B.n375 B.n278 585
R285 B.n278 B.n277 585
R286 B.n377 B.n376 585
R287 B.n378 B.n377 585
R288 B.n272 B.n271 585
R289 B.n273 B.n272 585
R290 B.n386 B.n385 585
R291 B.n385 B.n384 585
R292 B.n387 B.n270 585
R293 B.n270 B.n269 585
R294 B.n389 B.n388 585
R295 B.n390 B.n389 585
R296 B.n264 B.n263 585
R297 B.n265 B.n264 585
R298 B.n398 B.n397 585
R299 B.n397 B.n396 585
R300 B.n399 B.n262 585
R301 B.n262 B.n261 585
R302 B.n401 B.n400 585
R303 B.n402 B.n401 585
R304 B.n256 B.n255 585
R305 B.n257 B.n256 585
R306 B.n410 B.n409 585
R307 B.n409 B.n408 585
R308 B.n411 B.n254 585
R309 B.n254 B.n253 585
R310 B.n413 B.n412 585
R311 B.n414 B.n413 585
R312 B.n248 B.n247 585
R313 B.n249 B.n248 585
R314 B.n422 B.n421 585
R315 B.n421 B.n420 585
R316 B.n423 B.n246 585
R317 B.n246 B.n245 585
R318 B.n425 B.n424 585
R319 B.n426 B.n425 585
R320 B.n241 B.n240 585
R321 B.t5 B.n241 585
R322 B.n434 B.n433 585
R323 B.n433 B.n432 585
R324 B.n435 B.n239 585
R325 B.n239 B.n238 585
R326 B.n437 B.n436 585
R327 B.n438 B.n437 585
R328 B.n233 B.n232 585
R329 B.n234 B.n233 585
R330 B.n446 B.n445 585
R331 B.n445 B.n444 585
R332 B.n447 B.n231 585
R333 B.n231 B.n229 585
R334 B.n449 B.n448 585
R335 B.n450 B.n449 585
R336 B.n225 B.n224 585
R337 B.n230 B.n225 585
R338 B.n458 B.n457 585
R339 B.n457 B.n456 585
R340 B.n459 B.n223 585
R341 B.n223 B.n222 585
R342 B.n461 B.n460 585
R343 B.n462 B.n461 585
R344 B.n217 B.n216 585
R345 B.n218 B.n217 585
R346 B.n470 B.n469 585
R347 B.n469 B.n468 585
R348 B.n471 B.n215 585
R349 B.n215 B.n214 585
R350 B.n473 B.n472 585
R351 B.n474 B.n473 585
R352 B.n209 B.n208 585
R353 B.n210 B.n209 585
R354 B.n482 B.n481 585
R355 B.n481 B.n480 585
R356 B.n483 B.n207 585
R357 B.n207 B.n206 585
R358 B.n485 B.n484 585
R359 B.n486 B.n485 585
R360 B.n201 B.n200 585
R361 B.n202 B.n201 585
R362 B.n494 B.n493 585
R363 B.n493 B.n492 585
R364 B.n495 B.n199 585
R365 B.n199 B.n198 585
R366 B.n497 B.n496 585
R367 B.n498 B.n497 585
R368 B.n193 B.n192 585
R369 B.n194 B.n193 585
R370 B.n507 B.n506 585
R371 B.n506 B.n505 585
R372 B.n508 B.n191 585
R373 B.n504 B.n191 585
R374 B.n510 B.n509 585
R375 B.n511 B.n510 585
R376 B.n186 B.n185 585
R377 B.n187 B.n186 585
R378 B.n520 B.n519 585
R379 B.n519 B.n518 585
R380 B.n521 B.n184 585
R381 B.n184 B.n183 585
R382 B.n523 B.n522 585
R383 B.n524 B.n523 585
R384 B.n2 B.n0 585
R385 B.n4 B.n2 585
R386 B.n3 B.n1 585
R387 B.n702 B.n3 585
R388 B.n700 B.n699 585
R389 B.n701 B.n700 585
R390 B.n698 B.n9 585
R391 B.n9 B.n8 585
R392 B.n697 B.n696 585
R393 B.n696 B.n695 585
R394 B.n11 B.n10 585
R395 B.n694 B.n11 585
R396 B.n692 B.n691 585
R397 B.n693 B.n692 585
R398 B.n690 B.n15 585
R399 B.n18 B.n15 585
R400 B.n689 B.n688 585
R401 B.n688 B.n687 585
R402 B.n17 B.n16 585
R403 B.n686 B.n17 585
R404 B.n684 B.n683 585
R405 B.n685 B.n684 585
R406 B.n682 B.n23 585
R407 B.n23 B.n22 585
R408 B.n681 B.n680 585
R409 B.n680 B.n679 585
R410 B.n25 B.n24 585
R411 B.n678 B.n25 585
R412 B.n676 B.n675 585
R413 B.n677 B.n676 585
R414 B.n674 B.n30 585
R415 B.n30 B.n29 585
R416 B.n673 B.n672 585
R417 B.n672 B.n671 585
R418 B.n32 B.n31 585
R419 B.n670 B.n32 585
R420 B.n668 B.n667 585
R421 B.n669 B.n668 585
R422 B.n666 B.n37 585
R423 B.n37 B.n36 585
R424 B.n665 B.n664 585
R425 B.n664 B.n663 585
R426 B.n39 B.n38 585
R427 B.n662 B.n39 585
R428 B.n660 B.n659 585
R429 B.n661 B.n660 585
R430 B.n658 B.n44 585
R431 B.n44 B.n43 585
R432 B.n657 B.n656 585
R433 B.n656 B.n655 585
R434 B.n46 B.n45 585
R435 B.n654 B.n46 585
R436 B.n652 B.n651 585
R437 B.n653 B.n652 585
R438 B.n650 B.n51 585
R439 B.n51 B.n50 585
R440 B.n649 B.n648 585
R441 B.n648 B.n647 585
R442 B.n53 B.n52 585
R443 B.n646 B.n53 585
R444 B.n644 B.n643 585
R445 B.n645 B.n644 585
R446 B.n642 B.n58 585
R447 B.n58 B.n57 585
R448 B.n641 B.n640 585
R449 B.n640 B.n639 585
R450 B.n60 B.n59 585
R451 B.t3 B.n60 585
R452 B.n637 B.n636 585
R453 B.n638 B.n637 585
R454 B.n635 B.n65 585
R455 B.n65 B.n64 585
R456 B.n634 B.n633 585
R457 B.n633 B.n632 585
R458 B.n67 B.n66 585
R459 B.n631 B.n67 585
R460 B.n629 B.n628 585
R461 B.n630 B.n629 585
R462 B.n627 B.n72 585
R463 B.n72 B.n71 585
R464 B.n626 B.n625 585
R465 B.n625 B.n624 585
R466 B.n74 B.n73 585
R467 B.n623 B.n74 585
R468 B.n621 B.n620 585
R469 B.n622 B.n621 585
R470 B.n619 B.n79 585
R471 B.n79 B.n78 585
R472 B.n618 B.n617 585
R473 B.n617 B.n616 585
R474 B.n81 B.n80 585
R475 B.n615 B.n81 585
R476 B.n613 B.n612 585
R477 B.n614 B.n613 585
R478 B.n611 B.n86 585
R479 B.n86 B.n85 585
R480 B.n610 B.n609 585
R481 B.n609 B.n608 585
R482 B.n88 B.n87 585
R483 B.n607 B.n88 585
R484 B.n605 B.n604 585
R485 B.n606 B.n605 585
R486 B.n603 B.n93 585
R487 B.n93 B.n92 585
R488 B.n602 B.n601 585
R489 B.n601 B.n600 585
R490 B.n95 B.n94 585
R491 B.n599 B.n95 585
R492 B.n705 B.n704 585
R493 B.n704 B.n703 585
R494 B.n364 B.n280 463.671
R495 B.n118 B.n95 463.671
R496 B.n367 B.n282 463.671
R497 B.n596 B.n97 463.671
R498 B.n598 B.n597 256.663
R499 B.n598 B.n112 256.663
R500 B.n598 B.n111 256.663
R501 B.n598 B.n110 256.663
R502 B.n598 B.n109 256.663
R503 B.n598 B.n108 256.663
R504 B.n598 B.n107 256.663
R505 B.n598 B.n106 256.663
R506 B.n598 B.n105 256.663
R507 B.n598 B.n104 256.663
R508 B.n598 B.n103 256.663
R509 B.n598 B.n102 256.663
R510 B.n598 B.n101 256.663
R511 B.n598 B.n100 256.663
R512 B.n598 B.n99 256.663
R513 B.n598 B.n98 256.663
R514 B.n366 B.n365 256.663
R515 B.n366 B.n285 256.663
R516 B.n366 B.n286 256.663
R517 B.n366 B.n287 256.663
R518 B.n366 B.n288 256.663
R519 B.n366 B.n289 256.663
R520 B.n366 B.n290 256.663
R521 B.n366 B.n291 256.663
R522 B.n366 B.n292 256.663
R523 B.n366 B.n293 256.663
R524 B.n366 B.n294 256.663
R525 B.n366 B.n295 256.663
R526 B.n366 B.n296 256.663
R527 B.n366 B.n297 256.663
R528 B.n366 B.n298 256.663
R529 B.n304 B.t12 222.398
R530 B.n301 B.t19 222.398
R531 B.n116 B.t16 222.398
R532 B.n114 B.t8 222.398
R533 B.n366 B.n281 193.601
R534 B.n599 B.n598 193.601
R535 B.n304 B.t15 167.606
R536 B.n114 B.t10 167.606
R537 B.n301 B.t21 167.605
R538 B.n116 B.t17 167.605
R539 B.n373 B.n280 163.367
R540 B.n373 B.n278 163.367
R541 B.n377 B.n278 163.367
R542 B.n377 B.n272 163.367
R543 B.n385 B.n272 163.367
R544 B.n385 B.n270 163.367
R545 B.n389 B.n270 163.367
R546 B.n389 B.n264 163.367
R547 B.n397 B.n264 163.367
R548 B.n397 B.n262 163.367
R549 B.n401 B.n262 163.367
R550 B.n401 B.n256 163.367
R551 B.n409 B.n256 163.367
R552 B.n409 B.n254 163.367
R553 B.n413 B.n254 163.367
R554 B.n413 B.n248 163.367
R555 B.n421 B.n248 163.367
R556 B.n421 B.n246 163.367
R557 B.n425 B.n246 163.367
R558 B.n425 B.n241 163.367
R559 B.n433 B.n241 163.367
R560 B.n433 B.n239 163.367
R561 B.n437 B.n239 163.367
R562 B.n437 B.n233 163.367
R563 B.n445 B.n233 163.367
R564 B.n445 B.n231 163.367
R565 B.n449 B.n231 163.367
R566 B.n449 B.n225 163.367
R567 B.n457 B.n225 163.367
R568 B.n457 B.n223 163.367
R569 B.n461 B.n223 163.367
R570 B.n461 B.n217 163.367
R571 B.n469 B.n217 163.367
R572 B.n469 B.n215 163.367
R573 B.n473 B.n215 163.367
R574 B.n473 B.n209 163.367
R575 B.n481 B.n209 163.367
R576 B.n481 B.n207 163.367
R577 B.n485 B.n207 163.367
R578 B.n485 B.n201 163.367
R579 B.n493 B.n201 163.367
R580 B.n493 B.n199 163.367
R581 B.n497 B.n199 163.367
R582 B.n497 B.n193 163.367
R583 B.n506 B.n193 163.367
R584 B.n506 B.n191 163.367
R585 B.n510 B.n191 163.367
R586 B.n510 B.n186 163.367
R587 B.n519 B.n186 163.367
R588 B.n519 B.n184 163.367
R589 B.n523 B.n184 163.367
R590 B.n523 B.n2 163.367
R591 B.n704 B.n2 163.367
R592 B.n704 B.n3 163.367
R593 B.n700 B.n3 163.367
R594 B.n700 B.n9 163.367
R595 B.n696 B.n9 163.367
R596 B.n696 B.n11 163.367
R597 B.n692 B.n11 163.367
R598 B.n692 B.n15 163.367
R599 B.n688 B.n15 163.367
R600 B.n688 B.n17 163.367
R601 B.n684 B.n17 163.367
R602 B.n684 B.n23 163.367
R603 B.n680 B.n23 163.367
R604 B.n680 B.n25 163.367
R605 B.n676 B.n25 163.367
R606 B.n676 B.n30 163.367
R607 B.n672 B.n30 163.367
R608 B.n672 B.n32 163.367
R609 B.n668 B.n32 163.367
R610 B.n668 B.n37 163.367
R611 B.n664 B.n37 163.367
R612 B.n664 B.n39 163.367
R613 B.n660 B.n39 163.367
R614 B.n660 B.n44 163.367
R615 B.n656 B.n44 163.367
R616 B.n656 B.n46 163.367
R617 B.n652 B.n46 163.367
R618 B.n652 B.n51 163.367
R619 B.n648 B.n51 163.367
R620 B.n648 B.n53 163.367
R621 B.n644 B.n53 163.367
R622 B.n644 B.n58 163.367
R623 B.n640 B.n58 163.367
R624 B.n640 B.n60 163.367
R625 B.n637 B.n60 163.367
R626 B.n637 B.n65 163.367
R627 B.n633 B.n65 163.367
R628 B.n633 B.n67 163.367
R629 B.n629 B.n67 163.367
R630 B.n629 B.n72 163.367
R631 B.n625 B.n72 163.367
R632 B.n625 B.n74 163.367
R633 B.n621 B.n74 163.367
R634 B.n621 B.n79 163.367
R635 B.n617 B.n79 163.367
R636 B.n617 B.n81 163.367
R637 B.n613 B.n81 163.367
R638 B.n613 B.n86 163.367
R639 B.n609 B.n86 163.367
R640 B.n609 B.n88 163.367
R641 B.n605 B.n88 163.367
R642 B.n605 B.n93 163.367
R643 B.n601 B.n93 163.367
R644 B.n601 B.n95 163.367
R645 B.n300 B.n299 163.367
R646 B.n359 B.n299 163.367
R647 B.n357 B.n356 163.367
R648 B.n353 B.n352 163.367
R649 B.n349 B.n348 163.367
R650 B.n345 B.n344 163.367
R651 B.n341 B.n340 163.367
R652 B.n337 B.n336 163.367
R653 B.n333 B.n332 163.367
R654 B.n329 B.n328 163.367
R655 B.n325 B.n324 163.367
R656 B.n321 B.n320 163.367
R657 B.n317 B.n316 163.367
R658 B.n313 B.n312 163.367
R659 B.n309 B.n308 163.367
R660 B.n367 B.n284 163.367
R661 B.n371 B.n282 163.367
R662 B.n371 B.n276 163.367
R663 B.n379 B.n276 163.367
R664 B.n379 B.n274 163.367
R665 B.n383 B.n274 163.367
R666 B.n383 B.n268 163.367
R667 B.n391 B.n268 163.367
R668 B.n391 B.n266 163.367
R669 B.n395 B.n266 163.367
R670 B.n395 B.n260 163.367
R671 B.n403 B.n260 163.367
R672 B.n403 B.n258 163.367
R673 B.n407 B.n258 163.367
R674 B.n407 B.n252 163.367
R675 B.n415 B.n252 163.367
R676 B.n415 B.n250 163.367
R677 B.n419 B.n250 163.367
R678 B.n419 B.n244 163.367
R679 B.n427 B.n244 163.367
R680 B.n427 B.n242 163.367
R681 B.n431 B.n242 163.367
R682 B.n431 B.n237 163.367
R683 B.n439 B.n237 163.367
R684 B.n439 B.n235 163.367
R685 B.n443 B.n235 163.367
R686 B.n443 B.n228 163.367
R687 B.n451 B.n228 163.367
R688 B.n451 B.n226 163.367
R689 B.n455 B.n226 163.367
R690 B.n455 B.n221 163.367
R691 B.n463 B.n221 163.367
R692 B.n463 B.n219 163.367
R693 B.n467 B.n219 163.367
R694 B.n467 B.n213 163.367
R695 B.n475 B.n213 163.367
R696 B.n475 B.n211 163.367
R697 B.n479 B.n211 163.367
R698 B.n479 B.n205 163.367
R699 B.n487 B.n205 163.367
R700 B.n487 B.n203 163.367
R701 B.n491 B.n203 163.367
R702 B.n491 B.n197 163.367
R703 B.n499 B.n197 163.367
R704 B.n499 B.n195 163.367
R705 B.n503 B.n195 163.367
R706 B.n503 B.n190 163.367
R707 B.n512 B.n190 163.367
R708 B.n512 B.n188 163.367
R709 B.n517 B.n188 163.367
R710 B.n517 B.n182 163.367
R711 B.n525 B.n182 163.367
R712 B.n526 B.n525 163.367
R713 B.n526 B.n5 163.367
R714 B.n6 B.n5 163.367
R715 B.n7 B.n6 163.367
R716 B.n531 B.n7 163.367
R717 B.n531 B.n12 163.367
R718 B.n13 B.n12 163.367
R719 B.n14 B.n13 163.367
R720 B.n536 B.n14 163.367
R721 B.n536 B.n19 163.367
R722 B.n20 B.n19 163.367
R723 B.n21 B.n20 163.367
R724 B.n541 B.n21 163.367
R725 B.n541 B.n26 163.367
R726 B.n27 B.n26 163.367
R727 B.n28 B.n27 163.367
R728 B.n546 B.n28 163.367
R729 B.n546 B.n33 163.367
R730 B.n34 B.n33 163.367
R731 B.n35 B.n34 163.367
R732 B.n551 B.n35 163.367
R733 B.n551 B.n40 163.367
R734 B.n41 B.n40 163.367
R735 B.n42 B.n41 163.367
R736 B.n556 B.n42 163.367
R737 B.n556 B.n47 163.367
R738 B.n48 B.n47 163.367
R739 B.n49 B.n48 163.367
R740 B.n561 B.n49 163.367
R741 B.n561 B.n54 163.367
R742 B.n55 B.n54 163.367
R743 B.n56 B.n55 163.367
R744 B.n566 B.n56 163.367
R745 B.n566 B.n61 163.367
R746 B.n62 B.n61 163.367
R747 B.n63 B.n62 163.367
R748 B.n571 B.n63 163.367
R749 B.n571 B.n68 163.367
R750 B.n69 B.n68 163.367
R751 B.n70 B.n69 163.367
R752 B.n576 B.n70 163.367
R753 B.n576 B.n75 163.367
R754 B.n76 B.n75 163.367
R755 B.n77 B.n76 163.367
R756 B.n581 B.n77 163.367
R757 B.n581 B.n82 163.367
R758 B.n83 B.n82 163.367
R759 B.n84 B.n83 163.367
R760 B.n586 B.n84 163.367
R761 B.n586 B.n89 163.367
R762 B.n90 B.n89 163.367
R763 B.n91 B.n90 163.367
R764 B.n591 B.n91 163.367
R765 B.n591 B.n96 163.367
R766 B.n97 B.n96 163.367
R767 B.n122 B.n121 163.367
R768 B.n126 B.n125 163.367
R769 B.n130 B.n129 163.367
R770 B.n134 B.n133 163.367
R771 B.n138 B.n137 163.367
R772 B.n143 B.n142 163.367
R773 B.n147 B.n146 163.367
R774 B.n151 B.n150 163.367
R775 B.n155 B.n154 163.367
R776 B.n159 B.n158 163.367
R777 B.n164 B.n163 163.367
R778 B.n168 B.n167 163.367
R779 B.n172 B.n171 163.367
R780 B.n176 B.n175 163.367
R781 B.n178 B.n113 163.367
R782 B.n372 B.n281 108.8
R783 B.n372 B.n277 108.8
R784 B.n378 B.n277 108.8
R785 B.n378 B.n273 108.8
R786 B.n384 B.n273 108.8
R787 B.n384 B.n269 108.8
R788 B.n390 B.n269 108.8
R789 B.n396 B.n265 108.8
R790 B.n396 B.n261 108.8
R791 B.n402 B.n261 108.8
R792 B.n402 B.n257 108.8
R793 B.n408 B.n257 108.8
R794 B.n408 B.n253 108.8
R795 B.n414 B.n253 108.8
R796 B.n414 B.n249 108.8
R797 B.n420 B.n249 108.8
R798 B.n420 B.n245 108.8
R799 B.n426 B.n245 108.8
R800 B.n426 B.t5 108.8
R801 B.n432 B.t5 108.8
R802 B.n432 B.n238 108.8
R803 B.n438 B.n238 108.8
R804 B.n438 B.n234 108.8
R805 B.n444 B.n234 108.8
R806 B.n444 B.n229 108.8
R807 B.n450 B.n229 108.8
R808 B.n450 B.n230 108.8
R809 B.n456 B.n222 108.8
R810 B.n462 B.n222 108.8
R811 B.n462 B.n218 108.8
R812 B.n468 B.n218 108.8
R813 B.n468 B.n214 108.8
R814 B.n474 B.n214 108.8
R815 B.n474 B.n210 108.8
R816 B.n480 B.n210 108.8
R817 B.n486 B.n206 108.8
R818 B.n486 B.n202 108.8
R819 B.n492 B.n202 108.8
R820 B.n492 B.n198 108.8
R821 B.n498 B.n198 108.8
R822 B.n498 B.n194 108.8
R823 B.n505 B.n194 108.8
R824 B.n505 B.n504 108.8
R825 B.n511 B.n187 108.8
R826 B.n518 B.n187 108.8
R827 B.n518 B.n183 108.8
R828 B.n524 B.n183 108.8
R829 B.n524 B.n4 108.8
R830 B.n703 B.n4 108.8
R831 B.n703 B.n702 108.8
R832 B.n702 B.n701 108.8
R833 B.n701 B.n8 108.8
R834 B.n695 B.n8 108.8
R835 B.n695 B.n694 108.8
R836 B.n694 B.n693 108.8
R837 B.n687 B.n18 108.8
R838 B.n687 B.n686 108.8
R839 B.n686 B.n685 108.8
R840 B.n685 B.n22 108.8
R841 B.n679 B.n22 108.8
R842 B.n679 B.n678 108.8
R843 B.n678 B.n677 108.8
R844 B.n677 B.n29 108.8
R845 B.n671 B.n670 108.8
R846 B.n670 B.n669 108.8
R847 B.n669 B.n36 108.8
R848 B.n663 B.n36 108.8
R849 B.n663 B.n662 108.8
R850 B.n662 B.n661 108.8
R851 B.n661 B.n43 108.8
R852 B.n655 B.n43 108.8
R853 B.n654 B.n653 108.8
R854 B.n653 B.n50 108.8
R855 B.n647 B.n50 108.8
R856 B.n647 B.n646 108.8
R857 B.n646 B.n645 108.8
R858 B.n645 B.n57 108.8
R859 B.n639 B.n57 108.8
R860 B.n639 B.t3 108.8
R861 B.t3 B.n638 108.8
R862 B.n638 B.n64 108.8
R863 B.n632 B.n64 108.8
R864 B.n632 B.n631 108.8
R865 B.n631 B.n630 108.8
R866 B.n630 B.n71 108.8
R867 B.n624 B.n71 108.8
R868 B.n624 B.n623 108.8
R869 B.n623 B.n622 108.8
R870 B.n622 B.n78 108.8
R871 B.n616 B.n78 108.8
R872 B.n616 B.n615 108.8
R873 B.n614 B.n85 108.8
R874 B.n608 B.n85 108.8
R875 B.n608 B.n607 108.8
R876 B.n607 B.n606 108.8
R877 B.n606 B.n92 108.8
R878 B.n600 B.n92 108.8
R879 B.n600 B.n599 108.8
R880 B.n305 B.t14 108.454
R881 B.n115 B.t11 108.454
R882 B.n302 B.t20 108.454
R883 B.n117 B.t18 108.454
R884 B.n230 B.t2 105.6
R885 B.t0 B.n654 105.6
R886 B.n480 B.t7 102.4
R887 B.n671 B.t6 102.4
R888 B.n504 B.t1 99.2005
R889 B.n18 B.t4 99.2005
R890 B.n390 B.t13 89.6005
R891 B.t9 B.n614 89.6005
R892 B.n365 B.n364 71.676
R893 B.n359 B.n285 71.676
R894 B.n356 B.n286 71.676
R895 B.n352 B.n287 71.676
R896 B.n348 B.n288 71.676
R897 B.n344 B.n289 71.676
R898 B.n340 B.n290 71.676
R899 B.n336 B.n291 71.676
R900 B.n332 B.n292 71.676
R901 B.n328 B.n293 71.676
R902 B.n324 B.n294 71.676
R903 B.n320 B.n295 71.676
R904 B.n316 B.n296 71.676
R905 B.n312 B.n297 71.676
R906 B.n308 B.n298 71.676
R907 B.n118 B.n98 71.676
R908 B.n122 B.n99 71.676
R909 B.n126 B.n100 71.676
R910 B.n130 B.n101 71.676
R911 B.n134 B.n102 71.676
R912 B.n138 B.n103 71.676
R913 B.n143 B.n104 71.676
R914 B.n147 B.n105 71.676
R915 B.n151 B.n106 71.676
R916 B.n155 B.n107 71.676
R917 B.n159 B.n108 71.676
R918 B.n164 B.n109 71.676
R919 B.n168 B.n110 71.676
R920 B.n172 B.n111 71.676
R921 B.n176 B.n112 71.676
R922 B.n597 B.n113 71.676
R923 B.n597 B.n596 71.676
R924 B.n178 B.n112 71.676
R925 B.n175 B.n111 71.676
R926 B.n171 B.n110 71.676
R927 B.n167 B.n109 71.676
R928 B.n163 B.n108 71.676
R929 B.n158 B.n107 71.676
R930 B.n154 B.n106 71.676
R931 B.n150 B.n105 71.676
R932 B.n146 B.n104 71.676
R933 B.n142 B.n103 71.676
R934 B.n137 B.n102 71.676
R935 B.n133 B.n101 71.676
R936 B.n129 B.n100 71.676
R937 B.n125 B.n99 71.676
R938 B.n121 B.n98 71.676
R939 B.n365 B.n300 71.676
R940 B.n357 B.n285 71.676
R941 B.n353 B.n286 71.676
R942 B.n349 B.n287 71.676
R943 B.n345 B.n288 71.676
R944 B.n341 B.n289 71.676
R945 B.n337 B.n290 71.676
R946 B.n333 B.n291 71.676
R947 B.n329 B.n292 71.676
R948 B.n325 B.n293 71.676
R949 B.n321 B.n294 71.676
R950 B.n317 B.n295 71.676
R951 B.n313 B.n296 71.676
R952 B.n309 B.n297 71.676
R953 B.n298 B.n284 71.676
R954 B.n306 B.n305 59.5399
R955 B.n303 B.n302 59.5399
R956 B.n140 B.n117 59.5399
R957 B.n161 B.n115 59.5399
R958 B.n305 B.n304 59.152
R959 B.n302 B.n301 59.152
R960 B.n117 B.n116 59.152
R961 B.n115 B.n114 59.152
R962 B.n119 B.n94 30.1273
R963 B.n595 B.n594 30.1273
R964 B.n369 B.n368 30.1273
R965 B.n363 B.n279 30.1273
R966 B.t13 B.n265 19.2005
R967 B.n615 B.t9 19.2005
R968 B B.n705 18.0485
R969 B.n120 B.n119 10.6151
R970 B.n123 B.n120 10.6151
R971 B.n124 B.n123 10.6151
R972 B.n127 B.n124 10.6151
R973 B.n128 B.n127 10.6151
R974 B.n131 B.n128 10.6151
R975 B.n132 B.n131 10.6151
R976 B.n135 B.n132 10.6151
R977 B.n136 B.n135 10.6151
R978 B.n139 B.n136 10.6151
R979 B.n144 B.n141 10.6151
R980 B.n145 B.n144 10.6151
R981 B.n148 B.n145 10.6151
R982 B.n149 B.n148 10.6151
R983 B.n152 B.n149 10.6151
R984 B.n153 B.n152 10.6151
R985 B.n156 B.n153 10.6151
R986 B.n157 B.n156 10.6151
R987 B.n160 B.n157 10.6151
R988 B.n165 B.n162 10.6151
R989 B.n166 B.n165 10.6151
R990 B.n169 B.n166 10.6151
R991 B.n170 B.n169 10.6151
R992 B.n173 B.n170 10.6151
R993 B.n174 B.n173 10.6151
R994 B.n177 B.n174 10.6151
R995 B.n179 B.n177 10.6151
R996 B.n180 B.n179 10.6151
R997 B.n595 B.n180 10.6151
R998 B.n370 B.n369 10.6151
R999 B.n370 B.n275 10.6151
R1000 B.n380 B.n275 10.6151
R1001 B.n381 B.n380 10.6151
R1002 B.n382 B.n381 10.6151
R1003 B.n382 B.n267 10.6151
R1004 B.n392 B.n267 10.6151
R1005 B.n393 B.n392 10.6151
R1006 B.n394 B.n393 10.6151
R1007 B.n394 B.n259 10.6151
R1008 B.n404 B.n259 10.6151
R1009 B.n405 B.n404 10.6151
R1010 B.n406 B.n405 10.6151
R1011 B.n406 B.n251 10.6151
R1012 B.n416 B.n251 10.6151
R1013 B.n417 B.n416 10.6151
R1014 B.n418 B.n417 10.6151
R1015 B.n418 B.n243 10.6151
R1016 B.n428 B.n243 10.6151
R1017 B.n429 B.n428 10.6151
R1018 B.n430 B.n429 10.6151
R1019 B.n430 B.n236 10.6151
R1020 B.n440 B.n236 10.6151
R1021 B.n441 B.n440 10.6151
R1022 B.n442 B.n441 10.6151
R1023 B.n442 B.n227 10.6151
R1024 B.n452 B.n227 10.6151
R1025 B.n453 B.n452 10.6151
R1026 B.n454 B.n453 10.6151
R1027 B.n454 B.n220 10.6151
R1028 B.n464 B.n220 10.6151
R1029 B.n465 B.n464 10.6151
R1030 B.n466 B.n465 10.6151
R1031 B.n466 B.n212 10.6151
R1032 B.n476 B.n212 10.6151
R1033 B.n477 B.n476 10.6151
R1034 B.n478 B.n477 10.6151
R1035 B.n478 B.n204 10.6151
R1036 B.n488 B.n204 10.6151
R1037 B.n489 B.n488 10.6151
R1038 B.n490 B.n489 10.6151
R1039 B.n490 B.n196 10.6151
R1040 B.n500 B.n196 10.6151
R1041 B.n501 B.n500 10.6151
R1042 B.n502 B.n501 10.6151
R1043 B.n502 B.n189 10.6151
R1044 B.n513 B.n189 10.6151
R1045 B.n514 B.n513 10.6151
R1046 B.n516 B.n514 10.6151
R1047 B.n516 B.n515 10.6151
R1048 B.n515 B.n181 10.6151
R1049 B.n527 B.n181 10.6151
R1050 B.n528 B.n527 10.6151
R1051 B.n529 B.n528 10.6151
R1052 B.n530 B.n529 10.6151
R1053 B.n532 B.n530 10.6151
R1054 B.n533 B.n532 10.6151
R1055 B.n534 B.n533 10.6151
R1056 B.n535 B.n534 10.6151
R1057 B.n537 B.n535 10.6151
R1058 B.n538 B.n537 10.6151
R1059 B.n539 B.n538 10.6151
R1060 B.n540 B.n539 10.6151
R1061 B.n542 B.n540 10.6151
R1062 B.n543 B.n542 10.6151
R1063 B.n544 B.n543 10.6151
R1064 B.n545 B.n544 10.6151
R1065 B.n547 B.n545 10.6151
R1066 B.n548 B.n547 10.6151
R1067 B.n549 B.n548 10.6151
R1068 B.n550 B.n549 10.6151
R1069 B.n552 B.n550 10.6151
R1070 B.n553 B.n552 10.6151
R1071 B.n554 B.n553 10.6151
R1072 B.n555 B.n554 10.6151
R1073 B.n557 B.n555 10.6151
R1074 B.n558 B.n557 10.6151
R1075 B.n559 B.n558 10.6151
R1076 B.n560 B.n559 10.6151
R1077 B.n562 B.n560 10.6151
R1078 B.n563 B.n562 10.6151
R1079 B.n564 B.n563 10.6151
R1080 B.n565 B.n564 10.6151
R1081 B.n567 B.n565 10.6151
R1082 B.n568 B.n567 10.6151
R1083 B.n569 B.n568 10.6151
R1084 B.n570 B.n569 10.6151
R1085 B.n572 B.n570 10.6151
R1086 B.n573 B.n572 10.6151
R1087 B.n574 B.n573 10.6151
R1088 B.n575 B.n574 10.6151
R1089 B.n577 B.n575 10.6151
R1090 B.n578 B.n577 10.6151
R1091 B.n579 B.n578 10.6151
R1092 B.n580 B.n579 10.6151
R1093 B.n582 B.n580 10.6151
R1094 B.n583 B.n582 10.6151
R1095 B.n584 B.n583 10.6151
R1096 B.n585 B.n584 10.6151
R1097 B.n587 B.n585 10.6151
R1098 B.n588 B.n587 10.6151
R1099 B.n589 B.n588 10.6151
R1100 B.n590 B.n589 10.6151
R1101 B.n592 B.n590 10.6151
R1102 B.n593 B.n592 10.6151
R1103 B.n594 B.n593 10.6151
R1104 B.n363 B.n362 10.6151
R1105 B.n362 B.n361 10.6151
R1106 B.n361 B.n360 10.6151
R1107 B.n360 B.n358 10.6151
R1108 B.n358 B.n355 10.6151
R1109 B.n355 B.n354 10.6151
R1110 B.n354 B.n351 10.6151
R1111 B.n351 B.n350 10.6151
R1112 B.n350 B.n347 10.6151
R1113 B.n347 B.n346 10.6151
R1114 B.n343 B.n342 10.6151
R1115 B.n342 B.n339 10.6151
R1116 B.n339 B.n338 10.6151
R1117 B.n338 B.n335 10.6151
R1118 B.n335 B.n334 10.6151
R1119 B.n334 B.n331 10.6151
R1120 B.n331 B.n330 10.6151
R1121 B.n330 B.n327 10.6151
R1122 B.n327 B.n326 10.6151
R1123 B.n323 B.n322 10.6151
R1124 B.n322 B.n319 10.6151
R1125 B.n319 B.n318 10.6151
R1126 B.n318 B.n315 10.6151
R1127 B.n315 B.n314 10.6151
R1128 B.n314 B.n311 10.6151
R1129 B.n311 B.n310 10.6151
R1130 B.n310 B.n307 10.6151
R1131 B.n307 B.n283 10.6151
R1132 B.n368 B.n283 10.6151
R1133 B.n374 B.n279 10.6151
R1134 B.n375 B.n374 10.6151
R1135 B.n376 B.n375 10.6151
R1136 B.n376 B.n271 10.6151
R1137 B.n386 B.n271 10.6151
R1138 B.n387 B.n386 10.6151
R1139 B.n388 B.n387 10.6151
R1140 B.n388 B.n263 10.6151
R1141 B.n398 B.n263 10.6151
R1142 B.n399 B.n398 10.6151
R1143 B.n400 B.n399 10.6151
R1144 B.n400 B.n255 10.6151
R1145 B.n410 B.n255 10.6151
R1146 B.n411 B.n410 10.6151
R1147 B.n412 B.n411 10.6151
R1148 B.n412 B.n247 10.6151
R1149 B.n422 B.n247 10.6151
R1150 B.n423 B.n422 10.6151
R1151 B.n424 B.n423 10.6151
R1152 B.n424 B.n240 10.6151
R1153 B.n434 B.n240 10.6151
R1154 B.n435 B.n434 10.6151
R1155 B.n436 B.n435 10.6151
R1156 B.n436 B.n232 10.6151
R1157 B.n446 B.n232 10.6151
R1158 B.n447 B.n446 10.6151
R1159 B.n448 B.n447 10.6151
R1160 B.n448 B.n224 10.6151
R1161 B.n458 B.n224 10.6151
R1162 B.n459 B.n458 10.6151
R1163 B.n460 B.n459 10.6151
R1164 B.n460 B.n216 10.6151
R1165 B.n470 B.n216 10.6151
R1166 B.n471 B.n470 10.6151
R1167 B.n472 B.n471 10.6151
R1168 B.n472 B.n208 10.6151
R1169 B.n482 B.n208 10.6151
R1170 B.n483 B.n482 10.6151
R1171 B.n484 B.n483 10.6151
R1172 B.n484 B.n200 10.6151
R1173 B.n494 B.n200 10.6151
R1174 B.n495 B.n494 10.6151
R1175 B.n496 B.n495 10.6151
R1176 B.n496 B.n192 10.6151
R1177 B.n507 B.n192 10.6151
R1178 B.n508 B.n507 10.6151
R1179 B.n509 B.n508 10.6151
R1180 B.n509 B.n185 10.6151
R1181 B.n520 B.n185 10.6151
R1182 B.n521 B.n520 10.6151
R1183 B.n522 B.n521 10.6151
R1184 B.n522 B.n0 10.6151
R1185 B.n699 B.n1 10.6151
R1186 B.n699 B.n698 10.6151
R1187 B.n698 B.n697 10.6151
R1188 B.n697 B.n10 10.6151
R1189 B.n691 B.n10 10.6151
R1190 B.n691 B.n690 10.6151
R1191 B.n690 B.n689 10.6151
R1192 B.n689 B.n16 10.6151
R1193 B.n683 B.n16 10.6151
R1194 B.n683 B.n682 10.6151
R1195 B.n682 B.n681 10.6151
R1196 B.n681 B.n24 10.6151
R1197 B.n675 B.n24 10.6151
R1198 B.n675 B.n674 10.6151
R1199 B.n674 B.n673 10.6151
R1200 B.n673 B.n31 10.6151
R1201 B.n667 B.n31 10.6151
R1202 B.n667 B.n666 10.6151
R1203 B.n666 B.n665 10.6151
R1204 B.n665 B.n38 10.6151
R1205 B.n659 B.n38 10.6151
R1206 B.n659 B.n658 10.6151
R1207 B.n658 B.n657 10.6151
R1208 B.n657 B.n45 10.6151
R1209 B.n651 B.n45 10.6151
R1210 B.n651 B.n650 10.6151
R1211 B.n650 B.n649 10.6151
R1212 B.n649 B.n52 10.6151
R1213 B.n643 B.n52 10.6151
R1214 B.n643 B.n642 10.6151
R1215 B.n642 B.n641 10.6151
R1216 B.n641 B.n59 10.6151
R1217 B.n636 B.n59 10.6151
R1218 B.n636 B.n635 10.6151
R1219 B.n635 B.n634 10.6151
R1220 B.n634 B.n66 10.6151
R1221 B.n628 B.n66 10.6151
R1222 B.n628 B.n627 10.6151
R1223 B.n627 B.n626 10.6151
R1224 B.n626 B.n73 10.6151
R1225 B.n620 B.n73 10.6151
R1226 B.n620 B.n619 10.6151
R1227 B.n619 B.n618 10.6151
R1228 B.n618 B.n80 10.6151
R1229 B.n612 B.n80 10.6151
R1230 B.n612 B.n611 10.6151
R1231 B.n611 B.n610 10.6151
R1232 B.n610 B.n87 10.6151
R1233 B.n604 B.n87 10.6151
R1234 B.n604 B.n603 10.6151
R1235 B.n603 B.n602 10.6151
R1236 B.n602 B.n94 10.6151
R1237 B.n511 B.t1 9.6005
R1238 B.n693 B.t4 9.6005
R1239 B.n140 B.n139 9.36635
R1240 B.n162 B.n161 9.36635
R1241 B.n346 B.n303 9.36635
R1242 B.n323 B.n306 9.36635
R1243 B.t7 B.n206 6.4005
R1244 B.t6 B.n29 6.4005
R1245 B.n456 B.t2 3.2005
R1246 B.n655 B.t0 3.2005
R1247 B.n705 B.n0 2.81026
R1248 B.n705 B.n1 2.81026
R1249 B.n141 B.n140 1.24928
R1250 B.n161 B.n160 1.24928
R1251 B.n343 B.n303 1.24928
R1252 B.n326 B.n306 1.24928
R1253 VP.n21 VP.n20 161.3
R1254 VP.n22 VP.n17 161.3
R1255 VP.n24 VP.n23 161.3
R1256 VP.n25 VP.n16 161.3
R1257 VP.n27 VP.n26 161.3
R1258 VP.n28 VP.n15 161.3
R1259 VP.n30 VP.n29 161.3
R1260 VP.n32 VP.n31 161.3
R1261 VP.n33 VP.n13 161.3
R1262 VP.n35 VP.n34 161.3
R1263 VP.n36 VP.n12 161.3
R1264 VP.n38 VP.n37 161.3
R1265 VP.n39 VP.n11 161.3
R1266 VP.n72 VP.n0 161.3
R1267 VP.n71 VP.n70 161.3
R1268 VP.n69 VP.n1 161.3
R1269 VP.n68 VP.n67 161.3
R1270 VP.n66 VP.n2 161.3
R1271 VP.n65 VP.n64 161.3
R1272 VP.n63 VP.n62 161.3
R1273 VP.n61 VP.n4 161.3
R1274 VP.n60 VP.n59 161.3
R1275 VP.n58 VP.n5 161.3
R1276 VP.n57 VP.n56 161.3
R1277 VP.n55 VP.n6 161.3
R1278 VP.n54 VP.n53 161.3
R1279 VP.n52 VP.n51 161.3
R1280 VP.n50 VP.n8 161.3
R1281 VP.n49 VP.n48 161.3
R1282 VP.n47 VP.n9 161.3
R1283 VP.n46 VP.n45 161.3
R1284 VP.n44 VP.n10 161.3
R1285 VP.n43 VP.n42 106.954
R1286 VP.n74 VP.n73 106.954
R1287 VP.n41 VP.n40 106.954
R1288 VP.n19 VP.n18 71.8269
R1289 VP.n19 VP.t5 45.4874
R1290 VP.n49 VP.n9 45.2793
R1291 VP.n67 VP.n1 45.2793
R1292 VP.n34 VP.n12 45.2793
R1293 VP.n42 VP.n41 43.5298
R1294 VP.n56 VP.n5 40.4106
R1295 VP.n60 VP.n5 40.4106
R1296 VP.n27 VP.n16 40.4106
R1297 VP.n23 VP.n16 40.4106
R1298 VP.n50 VP.n49 35.5419
R1299 VP.n67 VP.n66 35.5419
R1300 VP.n34 VP.n33 35.5419
R1301 VP.n45 VP.n44 24.3439
R1302 VP.n45 VP.n9 24.3439
R1303 VP.n51 VP.n50 24.3439
R1304 VP.n55 VP.n54 24.3439
R1305 VP.n56 VP.n55 24.3439
R1306 VP.n61 VP.n60 24.3439
R1307 VP.n62 VP.n61 24.3439
R1308 VP.n66 VP.n65 24.3439
R1309 VP.n71 VP.n1 24.3439
R1310 VP.n72 VP.n71 24.3439
R1311 VP.n38 VP.n12 24.3439
R1312 VP.n39 VP.n38 24.3439
R1313 VP.n28 VP.n27 24.3439
R1314 VP.n29 VP.n28 24.3439
R1315 VP.n33 VP.n32 24.3439
R1316 VP.n22 VP.n21 24.3439
R1317 VP.n23 VP.n22 24.3439
R1318 VP.n51 VP.n7 23.1268
R1319 VP.n65 VP.n3 23.1268
R1320 VP.n32 VP.n14 23.1268
R1321 VP.n43 VP.t0 14.177
R1322 VP.n7 VP.t7 14.177
R1323 VP.n3 VP.t4 14.177
R1324 VP.n73 VP.t1 14.177
R1325 VP.n40 VP.t2 14.177
R1326 VP.n14 VP.t6 14.177
R1327 VP.n18 VP.t3 14.177
R1328 VP.n20 VP.n19 7.28005
R1329 VP.n44 VP.n43 3.65202
R1330 VP.n73 VP.n72 3.65202
R1331 VP.n40 VP.n39 3.65202
R1332 VP.n54 VP.n7 1.21767
R1333 VP.n62 VP.n3 1.21767
R1334 VP.n29 VP.n14 1.21767
R1335 VP.n21 VP.n18 1.21767
R1336 VP.n41 VP.n11 0.278398
R1337 VP.n42 VP.n10 0.278398
R1338 VP.n74 VP.n0 0.278398
R1339 VP.n20 VP.n17 0.189894
R1340 VP.n24 VP.n17 0.189894
R1341 VP.n25 VP.n24 0.189894
R1342 VP.n26 VP.n25 0.189894
R1343 VP.n26 VP.n15 0.189894
R1344 VP.n30 VP.n15 0.189894
R1345 VP.n31 VP.n30 0.189894
R1346 VP.n31 VP.n13 0.189894
R1347 VP.n35 VP.n13 0.189894
R1348 VP.n36 VP.n35 0.189894
R1349 VP.n37 VP.n36 0.189894
R1350 VP.n37 VP.n11 0.189894
R1351 VP.n46 VP.n10 0.189894
R1352 VP.n47 VP.n46 0.189894
R1353 VP.n48 VP.n47 0.189894
R1354 VP.n48 VP.n8 0.189894
R1355 VP.n52 VP.n8 0.189894
R1356 VP.n53 VP.n52 0.189894
R1357 VP.n53 VP.n6 0.189894
R1358 VP.n57 VP.n6 0.189894
R1359 VP.n58 VP.n57 0.189894
R1360 VP.n59 VP.n58 0.189894
R1361 VP.n59 VP.n4 0.189894
R1362 VP.n63 VP.n4 0.189894
R1363 VP.n64 VP.n63 0.189894
R1364 VP.n64 VP.n2 0.189894
R1365 VP.n68 VP.n2 0.189894
R1366 VP.n69 VP.n68 0.189894
R1367 VP.n70 VP.n69 0.189894
R1368 VP.n70 VP.n0 0.189894
R1369 VP VP.n74 0.153422
R1370 VDD1 VDD1.n0 116.573
R1371 VDD1.n3 VDD1.n2 116.46
R1372 VDD1.n3 VDD1.n1 116.46
R1373 VDD1.n5 VDD1.n4 115.201
R1374 VDD1.n5 VDD1.n3 37.5095
R1375 VDD1.n4 VDD1.t2 12.3755
R1376 VDD1.n4 VDD1.t6 12.3755
R1377 VDD1.n0 VDD1.t4 12.3755
R1378 VDD1.n0 VDD1.t0 12.3755
R1379 VDD1.n2 VDD1.t7 12.3755
R1380 VDD1.n2 VDD1.t1 12.3755
R1381 VDD1.n1 VDD1.t3 12.3755
R1382 VDD1.n1 VDD1.t5 12.3755
R1383 VDD1 VDD1.n5 1.25697
R1384 VTAIL.n15 VTAIL.t7 110.897
R1385 VTAIL.n2 VTAIL.t1 110.897
R1386 VTAIL.n3 VTAIL.t14 110.897
R1387 VTAIL.n6 VTAIL.t15 110.897
R1388 VTAIL.n14 VTAIL.t13 110.897
R1389 VTAIL.n11 VTAIL.t10 110.897
R1390 VTAIL.n10 VTAIL.t5 110.897
R1391 VTAIL.n7 VTAIL.t4 110.897
R1392 VTAIL.n1 VTAIL.n0 98.5218
R1393 VTAIL.n5 VTAIL.n4 98.5218
R1394 VTAIL.n13 VTAIL.n12 98.5218
R1395 VTAIL.n9 VTAIL.n8 98.5218
R1396 VTAIL.n15 VTAIL.n14 16.3755
R1397 VTAIL.n7 VTAIL.n6 16.3755
R1398 VTAIL.n0 VTAIL.t3 12.3755
R1399 VTAIL.n0 VTAIL.t2 12.3755
R1400 VTAIL.n4 VTAIL.t8 12.3755
R1401 VTAIL.n4 VTAIL.t11 12.3755
R1402 VTAIL.n12 VTAIL.t12 12.3755
R1403 VTAIL.n12 VTAIL.t9 12.3755
R1404 VTAIL.n8 VTAIL.t0 12.3755
R1405 VTAIL.n8 VTAIL.t6 12.3755
R1406 VTAIL.n9 VTAIL.n7 2.62981
R1407 VTAIL.n10 VTAIL.n9 2.62981
R1408 VTAIL.n13 VTAIL.n11 2.62981
R1409 VTAIL.n14 VTAIL.n13 2.62981
R1410 VTAIL.n6 VTAIL.n5 2.62981
R1411 VTAIL.n5 VTAIL.n3 2.62981
R1412 VTAIL.n2 VTAIL.n1 2.62981
R1413 VTAIL VTAIL.n15 2.57162
R1414 VTAIL.n11 VTAIL.n10 0.470328
R1415 VTAIL.n3 VTAIL.n2 0.470328
R1416 VTAIL VTAIL.n1 0.0586897
R1417 VN.n59 VN.n31 161.3
R1418 VN.n58 VN.n57 161.3
R1419 VN.n56 VN.n32 161.3
R1420 VN.n55 VN.n54 161.3
R1421 VN.n53 VN.n33 161.3
R1422 VN.n52 VN.n51 161.3
R1423 VN.n50 VN.n49 161.3
R1424 VN.n48 VN.n35 161.3
R1425 VN.n47 VN.n46 161.3
R1426 VN.n45 VN.n36 161.3
R1427 VN.n44 VN.n43 161.3
R1428 VN.n42 VN.n37 161.3
R1429 VN.n41 VN.n40 161.3
R1430 VN.n28 VN.n0 161.3
R1431 VN.n27 VN.n26 161.3
R1432 VN.n25 VN.n1 161.3
R1433 VN.n24 VN.n23 161.3
R1434 VN.n22 VN.n2 161.3
R1435 VN.n21 VN.n20 161.3
R1436 VN.n19 VN.n18 161.3
R1437 VN.n17 VN.n4 161.3
R1438 VN.n16 VN.n15 161.3
R1439 VN.n14 VN.n5 161.3
R1440 VN.n13 VN.n12 161.3
R1441 VN.n11 VN.n6 161.3
R1442 VN.n10 VN.n9 161.3
R1443 VN.n30 VN.n29 106.954
R1444 VN.n61 VN.n60 106.954
R1445 VN.n8 VN.n7 71.8269
R1446 VN.n39 VN.n38 71.8269
R1447 VN.n8 VN.t0 45.4874
R1448 VN.n39 VN.t6 45.4874
R1449 VN.n23 VN.n1 45.2793
R1450 VN.n54 VN.n32 45.2793
R1451 VN VN.n61 43.8087
R1452 VN.n12 VN.n5 40.4106
R1453 VN.n16 VN.n5 40.4106
R1454 VN.n43 VN.n36 40.4106
R1455 VN.n47 VN.n36 40.4106
R1456 VN.n23 VN.n22 35.5419
R1457 VN.n54 VN.n53 35.5419
R1458 VN.n11 VN.n10 24.3439
R1459 VN.n12 VN.n11 24.3439
R1460 VN.n17 VN.n16 24.3439
R1461 VN.n18 VN.n17 24.3439
R1462 VN.n22 VN.n21 24.3439
R1463 VN.n27 VN.n1 24.3439
R1464 VN.n28 VN.n27 24.3439
R1465 VN.n43 VN.n42 24.3439
R1466 VN.n42 VN.n41 24.3439
R1467 VN.n53 VN.n52 24.3439
R1468 VN.n49 VN.n48 24.3439
R1469 VN.n48 VN.n47 24.3439
R1470 VN.n59 VN.n58 24.3439
R1471 VN.n58 VN.n32 24.3439
R1472 VN.n21 VN.n3 23.1268
R1473 VN.n52 VN.n34 23.1268
R1474 VN.n7 VN.t2 14.177
R1475 VN.n3 VN.t1 14.177
R1476 VN.n29 VN.t7 14.177
R1477 VN.n38 VN.t4 14.177
R1478 VN.n34 VN.t5 14.177
R1479 VN.n60 VN.t3 14.177
R1480 VN.n40 VN.n39 7.28005
R1481 VN.n9 VN.n8 7.28005
R1482 VN.n29 VN.n28 3.65202
R1483 VN.n60 VN.n59 3.65202
R1484 VN.n10 VN.n7 1.21767
R1485 VN.n18 VN.n3 1.21767
R1486 VN.n41 VN.n38 1.21767
R1487 VN.n49 VN.n34 1.21767
R1488 VN.n61 VN.n31 0.278398
R1489 VN.n30 VN.n0 0.278398
R1490 VN.n57 VN.n31 0.189894
R1491 VN.n57 VN.n56 0.189894
R1492 VN.n56 VN.n55 0.189894
R1493 VN.n55 VN.n33 0.189894
R1494 VN.n51 VN.n33 0.189894
R1495 VN.n51 VN.n50 0.189894
R1496 VN.n50 VN.n35 0.189894
R1497 VN.n46 VN.n35 0.189894
R1498 VN.n46 VN.n45 0.189894
R1499 VN.n45 VN.n44 0.189894
R1500 VN.n44 VN.n37 0.189894
R1501 VN.n40 VN.n37 0.189894
R1502 VN.n9 VN.n6 0.189894
R1503 VN.n13 VN.n6 0.189894
R1504 VN.n14 VN.n13 0.189894
R1505 VN.n15 VN.n14 0.189894
R1506 VN.n15 VN.n4 0.189894
R1507 VN.n19 VN.n4 0.189894
R1508 VN.n20 VN.n19 0.189894
R1509 VN.n20 VN.n2 0.189894
R1510 VN.n24 VN.n2 0.189894
R1511 VN.n25 VN.n24 0.189894
R1512 VN.n26 VN.n25 0.189894
R1513 VN.n26 VN.n0 0.189894
R1514 VN VN.n30 0.153422
R1515 VDD2.n2 VDD2.n1 116.46
R1516 VDD2.n2 VDD2.n0 116.46
R1517 VDD2 VDD2.n5 116.457
R1518 VDD2.n4 VDD2.n3 115.201
R1519 VDD2.n4 VDD2.n2 36.9265
R1520 VDD2.n5 VDD2.t3 12.3755
R1521 VDD2.n5 VDD2.t1 12.3755
R1522 VDD2.n3 VDD2.t4 12.3755
R1523 VDD2.n3 VDD2.t2 12.3755
R1524 VDD2.n1 VDD2.t6 12.3755
R1525 VDD2.n1 VDD2.t0 12.3755
R1526 VDD2.n0 VDD2.t7 12.3755
R1527 VDD2.n0 VDD2.t5 12.3755
R1528 VDD2 VDD2.n4 1.37334
C0 VDD1 VDD2 1.83766f
C1 VDD1 VTAIL 4.68812f
C2 VN VP 5.8989f
C3 VDD2 VP 0.539483f
C4 VDD2 VN 1.57452f
C5 VTAIL VP 2.81545f
C6 VTAIL VN 2.80135f
C7 VDD2 VTAIL 4.74334f
C8 VDD1 VP 1.95324f
C9 VDD1 VN 0.157569f
C10 VDD2 B 4.440573f
C11 VDD1 B 4.872541f
C12 VTAIL B 3.842754f
C13 VN B 14.950311f
C14 VP B 13.58422f
C15 VDD2.t7 B 0.022704f
C16 VDD2.t5 B 0.022704f
C17 VDD2.n0 B 0.134265f
C18 VDD2.t6 B 0.022704f
C19 VDD2.t0 B 0.022704f
C20 VDD2.n1 B 0.134265f
C21 VDD2.n2 B 1.92354f
C22 VDD2.t4 B 0.022704f
C23 VDD2.t2 B 0.022704f
C24 VDD2.n3 B 0.13033f
C25 VDD2.n4 B 1.55005f
C26 VDD2.t3 B 0.022704f
C27 VDD2.t1 B 0.022704f
C28 VDD2.n5 B 0.134251f
C29 VN.n0 B 0.035039f
C30 VN.t7 B 0.256595f
C31 VN.n1 B 0.051369f
C32 VN.n2 B 0.026575f
C33 VN.t1 B 0.256595f
C34 VN.n3 B 0.132617f
C35 VN.n4 B 0.026575f
C36 VN.n5 B 0.021505f
C37 VN.n6 B 0.026575f
C38 VN.t2 B 0.256595f
C39 VN.n7 B 0.202835f
C40 VN.t0 B 0.463313f
C41 VN.n8 B 0.209915f
C42 VN.n9 B 0.259981f
C43 VN.n10 B 0.02643f
C44 VN.n11 B 0.049778f
C45 VN.n12 B 0.0531f
C46 VN.n13 B 0.026575f
C47 VN.n14 B 0.026575f
C48 VN.n15 B 0.026575f
C49 VN.n16 B 0.0531f
C50 VN.n17 B 0.049778f
C51 VN.n18 B 0.02643f
C52 VN.n19 B 0.026575f
C53 VN.n20 B 0.026575f
C54 VN.n21 B 0.048549f
C55 VN.n22 B 0.053959f
C56 VN.n23 B 0.022378f
C57 VN.n24 B 0.026575f
C58 VN.n25 B 0.026575f
C59 VN.n26 B 0.026575f
C60 VN.n27 B 0.049778f
C61 VN.n28 B 0.028887f
C62 VN.n29 B 0.217419f
C63 VN.n30 B 0.04832f
C64 VN.n31 B 0.035039f
C65 VN.t3 B 0.256595f
C66 VN.n32 B 0.051369f
C67 VN.n33 B 0.026575f
C68 VN.t5 B 0.256595f
C69 VN.n34 B 0.132617f
C70 VN.n35 B 0.026575f
C71 VN.n36 B 0.021505f
C72 VN.n37 B 0.026575f
C73 VN.t4 B 0.256595f
C74 VN.n38 B 0.202835f
C75 VN.t6 B 0.463313f
C76 VN.n39 B 0.209915f
C77 VN.n40 B 0.259981f
C78 VN.n41 B 0.02643f
C79 VN.n42 B 0.049778f
C80 VN.n43 B 0.0531f
C81 VN.n44 B 0.026575f
C82 VN.n45 B 0.026575f
C83 VN.n46 B 0.026575f
C84 VN.n47 B 0.0531f
C85 VN.n48 B 0.049778f
C86 VN.n49 B 0.02643f
C87 VN.n50 B 0.026575f
C88 VN.n51 B 0.026575f
C89 VN.n52 B 0.048549f
C90 VN.n53 B 0.053959f
C91 VN.n54 B 0.022378f
C92 VN.n55 B 0.026575f
C93 VN.n56 B 0.026575f
C94 VN.n57 B 0.026575f
C95 VN.n58 B 0.049778f
C96 VN.n59 B 0.028887f
C97 VN.n60 B 0.217419f
C98 VN.n61 B 1.21672f
C99 VTAIL.t3 B 0.042724f
C100 VTAIL.t2 B 0.042724f
C101 VTAIL.n0 B 0.204484f
C102 VTAIL.n1 B 0.534717f
C103 VTAIL.t1 B 0.289951f
C104 VTAIL.n2 B 0.610591f
C105 VTAIL.t14 B 0.289951f
C106 VTAIL.n3 B 0.610591f
C107 VTAIL.t8 B 0.042724f
C108 VTAIL.t11 B 0.042724f
C109 VTAIL.n4 B 0.204484f
C110 VTAIL.n5 B 0.814666f
C111 VTAIL.t15 B 0.289951f
C112 VTAIL.n6 B 1.45491f
C113 VTAIL.t4 B 0.289951f
C114 VTAIL.n7 B 1.45491f
C115 VTAIL.t0 B 0.042724f
C116 VTAIL.t6 B 0.042724f
C117 VTAIL.n8 B 0.204484f
C118 VTAIL.n9 B 0.814665f
C119 VTAIL.t5 B 0.289951f
C120 VTAIL.n10 B 0.61059f
C121 VTAIL.t10 B 0.289951f
C122 VTAIL.n11 B 0.61059f
C123 VTAIL.t12 B 0.042724f
C124 VTAIL.t9 B 0.042724f
C125 VTAIL.n12 B 0.204484f
C126 VTAIL.n13 B 0.814665f
C127 VTAIL.t13 B 0.289951f
C128 VTAIL.n14 B 1.45491f
C129 VTAIL.t7 B 0.289951f
C130 VTAIL.n15 B 1.44858f
C131 VDD1.t4 B 0.022388f
C132 VDD1.t0 B 0.022388f
C133 VDD1.n0 B 0.132815f
C134 VDD1.t3 B 0.022388f
C135 VDD1.t5 B 0.022388f
C136 VDD1.n1 B 0.132397f
C137 VDD1.t7 B 0.022388f
C138 VDD1.t1 B 0.022388f
C139 VDD1.n2 B 0.132397f
C140 VDD1.n3 B 1.93375f
C141 VDD1.t2 B 0.022388f
C142 VDD1.t6 B 0.022388f
C143 VDD1.n4 B 0.128516f
C144 VDD1.n5 B 1.55026f
C145 VP.n0 B 0.03519f
C146 VP.t1 B 0.257702f
C147 VP.n1 B 0.05159f
C148 VP.n2 B 0.02669f
C149 VP.t4 B 0.257702f
C150 VP.n3 B 0.133189f
C151 VP.n4 B 0.02669f
C152 VP.n5 B 0.021598f
C153 VP.n6 B 0.02669f
C154 VP.t7 B 0.257702f
C155 VP.n7 B 0.133189f
C156 VP.n8 B 0.02669f
C157 VP.n9 B 0.05159f
C158 VP.n10 B 0.03519f
C159 VP.t0 B 0.257702f
C160 VP.n11 B 0.03519f
C161 VP.t2 B 0.257702f
C162 VP.n12 B 0.05159f
C163 VP.n13 B 0.02669f
C164 VP.t6 B 0.257702f
C165 VP.n14 B 0.133189f
C166 VP.n15 B 0.02669f
C167 VP.n16 B 0.021598f
C168 VP.n17 B 0.02669f
C169 VP.t3 B 0.257702f
C170 VP.n18 B 0.20371f
C171 VP.t5 B 0.465311f
C172 VP.n19 B 0.21082f
C173 VP.n20 B 0.261102f
C174 VP.n21 B 0.026544f
C175 VP.n22 B 0.049992f
C176 VP.n23 B 0.053329f
C177 VP.n24 B 0.02669f
C178 VP.n25 B 0.02669f
C179 VP.n26 B 0.02669f
C180 VP.n27 B 0.053329f
C181 VP.n28 B 0.049992f
C182 VP.n29 B 0.026544f
C183 VP.n30 B 0.02669f
C184 VP.n31 B 0.02669f
C185 VP.n32 B 0.048758f
C186 VP.n33 B 0.054192f
C187 VP.n34 B 0.022474f
C188 VP.n35 B 0.02669f
C189 VP.n36 B 0.02669f
C190 VP.n37 B 0.02669f
C191 VP.n38 B 0.049992f
C192 VP.n39 B 0.029012f
C193 VP.n40 B 0.218357f
C194 VP.n41 B 1.20729f
C195 VP.n42 B 1.22927f
C196 VP.n43 B 0.218357f
C197 VP.n44 B 0.029012f
C198 VP.n45 B 0.049992f
C199 VP.n46 B 0.02669f
C200 VP.n47 B 0.02669f
C201 VP.n48 B 0.02669f
C202 VP.n49 B 0.022474f
C203 VP.n50 B 0.054192f
C204 VP.n51 B 0.048758f
C205 VP.n52 B 0.02669f
C206 VP.n53 B 0.02669f
C207 VP.n54 B 0.026544f
C208 VP.n55 B 0.049992f
C209 VP.n56 B 0.053329f
C210 VP.n57 B 0.02669f
C211 VP.n58 B 0.02669f
C212 VP.n59 B 0.02669f
C213 VP.n60 B 0.053329f
C214 VP.n61 B 0.049992f
C215 VP.n62 B 0.026544f
C216 VP.n63 B 0.02669f
C217 VP.n64 B 0.02669f
C218 VP.n65 B 0.048758f
C219 VP.n66 B 0.054192f
C220 VP.n67 B 0.022474f
C221 VP.n68 B 0.02669f
C222 VP.n69 B 0.02669f
C223 VP.n70 B 0.02669f
C224 VP.n71 B 0.049992f
C225 VP.n72 B 0.029012f
C226 VP.n73 B 0.218357f
C227 VP.n74 B 0.048529f
.ends

