* NGSPICE file created from diff_pair_sample_1081.ext - technology: sky130A

.subckt diff_pair_sample_1081 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=1.0461 pd=6.67 as=2.4726 ps=13.46 w=6.34 l=2.15
X1 B.t11 B.t9 B.t10 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=0 ps=0 w=6.34 l=2.15
X2 VTAIL.t7 VN.t0 VDD2.t3 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=1.0461 ps=6.67 w=6.34 l=2.15
X3 VDD1.t2 VP.t1 VTAIL.t4 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=1.0461 pd=6.67 as=2.4726 ps=13.46 w=6.34 l=2.15
X4 VTAIL.t3 VP.t2 VDD1.t1 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=1.0461 ps=6.67 w=6.34 l=2.15
X5 VTAIL.t5 VP.t3 VDD1.t0 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=1.0461 ps=6.67 w=6.34 l=2.15
X6 VDD2.t2 VN.t1 VTAIL.t2 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=1.0461 pd=6.67 as=2.4726 ps=13.46 w=6.34 l=2.15
X7 VDD2.t1 VN.t2 VTAIL.t0 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=1.0461 pd=6.67 as=2.4726 ps=13.46 w=6.34 l=2.15
X8 B.t8 B.t6 B.t7 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=0 ps=0 w=6.34 l=2.15
X9 VTAIL.t1 VN.t3 VDD2.t0 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=1.0461 ps=6.67 w=6.34 l=2.15
X10 B.t5 B.t3 B.t4 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=0 ps=0 w=6.34 l=2.15
X11 B.t2 B.t0 B.t1 w_n2458_n2236# sky130_fd_pr__pfet_01v8 ad=2.4726 pd=13.46 as=0 ps=0 w=6.34 l=2.15
R0 VP.n12 VP.n0 161.3
R1 VP.n11 VP.n10 161.3
R2 VP.n9 VP.n1 161.3
R3 VP.n8 VP.n7 161.3
R4 VP.n6 VP.n2 161.3
R5 VP.n3 VP.t3 106.466
R6 VP.n3 VP.t0 105.838
R7 VP.n5 VP.n4 99.1042
R8 VP.n14 VP.n13 99.1042
R9 VP.n5 VP.t2 71.0675
R10 VP.n13 VP.t1 71.0675
R11 VP.n4 VP.n3 46.4927
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 11.8046
R17 VP.n13 VP.n12 11.8046
R18 VP.n4 VP.n2 0.278335
R19 VP.n14 VP.n0 0.278335
R20 VP.n8 VP.n2 0.189894
R21 VP.n9 VP.n8 0.189894
R22 VP.n10 VP.n9 0.189894
R23 VP.n10 VP.n0 0.189894
R24 VP VP.n14 0.153485
R25 VTAIL.n5 VTAIL.t5 78.2887
R26 VTAIL.n4 VTAIL.t2 78.2887
R27 VTAIL.n3 VTAIL.t7 78.2887
R28 VTAIL.n7 VTAIL.t0 78.2886
R29 VTAIL.n0 VTAIL.t1 78.2886
R30 VTAIL.n1 VTAIL.t4 78.2886
R31 VTAIL.n2 VTAIL.t3 78.2886
R32 VTAIL.n6 VTAIL.t6 78.2886
R33 VTAIL.n7 VTAIL.n6 19.9703
R34 VTAIL.n3 VTAIL.n2 19.9703
R35 VTAIL.n4 VTAIL.n3 2.13843
R36 VTAIL.n6 VTAIL.n5 2.13843
R37 VTAIL.n2 VTAIL.n1 2.13843
R38 VTAIL VTAIL.n0 1.12766
R39 VTAIL VTAIL.n7 1.01128
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 125.96
R43 VDD1 VDD1.n0 89.8986
R44 VDD1.n0 VDD1.t0 5.12747
R45 VDD1.n0 VDD1.t3 5.12747
R46 VDD1.n1 VDD1.t1 5.12747
R47 VDD1.n1 VDD1.t2 5.12747
R48 B.n356 B.n355 585
R49 B.n357 B.n50 585
R50 B.n359 B.n358 585
R51 B.n360 B.n49 585
R52 B.n362 B.n361 585
R53 B.n363 B.n48 585
R54 B.n365 B.n364 585
R55 B.n366 B.n47 585
R56 B.n368 B.n367 585
R57 B.n369 B.n46 585
R58 B.n371 B.n370 585
R59 B.n372 B.n45 585
R60 B.n374 B.n373 585
R61 B.n375 B.n44 585
R62 B.n377 B.n376 585
R63 B.n378 B.n43 585
R64 B.n380 B.n379 585
R65 B.n381 B.n42 585
R66 B.n383 B.n382 585
R67 B.n384 B.n41 585
R68 B.n386 B.n385 585
R69 B.n387 B.n40 585
R70 B.n389 B.n388 585
R71 B.n390 B.n39 585
R72 B.n392 B.n391 585
R73 B.n394 B.n393 585
R74 B.n395 B.n35 585
R75 B.n397 B.n396 585
R76 B.n398 B.n34 585
R77 B.n400 B.n399 585
R78 B.n401 B.n33 585
R79 B.n403 B.n402 585
R80 B.n404 B.n32 585
R81 B.n406 B.n405 585
R82 B.n408 B.n29 585
R83 B.n410 B.n409 585
R84 B.n411 B.n28 585
R85 B.n413 B.n412 585
R86 B.n414 B.n27 585
R87 B.n416 B.n415 585
R88 B.n417 B.n26 585
R89 B.n419 B.n418 585
R90 B.n420 B.n25 585
R91 B.n422 B.n421 585
R92 B.n423 B.n24 585
R93 B.n425 B.n424 585
R94 B.n426 B.n23 585
R95 B.n428 B.n427 585
R96 B.n429 B.n22 585
R97 B.n431 B.n430 585
R98 B.n432 B.n21 585
R99 B.n434 B.n433 585
R100 B.n435 B.n20 585
R101 B.n437 B.n436 585
R102 B.n438 B.n19 585
R103 B.n440 B.n439 585
R104 B.n441 B.n18 585
R105 B.n443 B.n442 585
R106 B.n444 B.n17 585
R107 B.n354 B.n51 585
R108 B.n353 B.n352 585
R109 B.n351 B.n52 585
R110 B.n350 B.n349 585
R111 B.n348 B.n53 585
R112 B.n347 B.n346 585
R113 B.n345 B.n54 585
R114 B.n344 B.n343 585
R115 B.n342 B.n55 585
R116 B.n341 B.n340 585
R117 B.n339 B.n56 585
R118 B.n338 B.n337 585
R119 B.n336 B.n57 585
R120 B.n335 B.n334 585
R121 B.n333 B.n58 585
R122 B.n332 B.n331 585
R123 B.n330 B.n59 585
R124 B.n329 B.n328 585
R125 B.n327 B.n60 585
R126 B.n326 B.n325 585
R127 B.n324 B.n61 585
R128 B.n323 B.n322 585
R129 B.n321 B.n62 585
R130 B.n320 B.n319 585
R131 B.n318 B.n63 585
R132 B.n317 B.n316 585
R133 B.n315 B.n64 585
R134 B.n314 B.n313 585
R135 B.n312 B.n65 585
R136 B.n311 B.n310 585
R137 B.n309 B.n66 585
R138 B.n308 B.n307 585
R139 B.n306 B.n67 585
R140 B.n305 B.n304 585
R141 B.n303 B.n68 585
R142 B.n302 B.n301 585
R143 B.n300 B.n69 585
R144 B.n299 B.n298 585
R145 B.n297 B.n70 585
R146 B.n296 B.n295 585
R147 B.n294 B.n71 585
R148 B.n293 B.n292 585
R149 B.n291 B.n72 585
R150 B.n290 B.n289 585
R151 B.n288 B.n73 585
R152 B.n287 B.n286 585
R153 B.n285 B.n74 585
R154 B.n284 B.n283 585
R155 B.n282 B.n75 585
R156 B.n281 B.n280 585
R157 B.n279 B.n76 585
R158 B.n278 B.n277 585
R159 B.n276 B.n77 585
R160 B.n275 B.n274 585
R161 B.n273 B.n78 585
R162 B.n272 B.n271 585
R163 B.n270 B.n79 585
R164 B.n269 B.n268 585
R165 B.n267 B.n80 585
R166 B.n266 B.n265 585
R167 B.n264 B.n81 585
R168 B.n174 B.n115 585
R169 B.n176 B.n175 585
R170 B.n177 B.n114 585
R171 B.n179 B.n178 585
R172 B.n180 B.n113 585
R173 B.n182 B.n181 585
R174 B.n183 B.n112 585
R175 B.n185 B.n184 585
R176 B.n186 B.n111 585
R177 B.n188 B.n187 585
R178 B.n189 B.n110 585
R179 B.n191 B.n190 585
R180 B.n192 B.n109 585
R181 B.n194 B.n193 585
R182 B.n195 B.n108 585
R183 B.n197 B.n196 585
R184 B.n198 B.n107 585
R185 B.n200 B.n199 585
R186 B.n201 B.n106 585
R187 B.n203 B.n202 585
R188 B.n204 B.n105 585
R189 B.n206 B.n205 585
R190 B.n207 B.n104 585
R191 B.n209 B.n208 585
R192 B.n210 B.n101 585
R193 B.n213 B.n212 585
R194 B.n214 B.n100 585
R195 B.n216 B.n215 585
R196 B.n217 B.n99 585
R197 B.n219 B.n218 585
R198 B.n220 B.n98 585
R199 B.n222 B.n221 585
R200 B.n223 B.n97 585
R201 B.n225 B.n224 585
R202 B.n227 B.n226 585
R203 B.n228 B.n93 585
R204 B.n230 B.n229 585
R205 B.n231 B.n92 585
R206 B.n233 B.n232 585
R207 B.n234 B.n91 585
R208 B.n236 B.n235 585
R209 B.n237 B.n90 585
R210 B.n239 B.n238 585
R211 B.n240 B.n89 585
R212 B.n242 B.n241 585
R213 B.n243 B.n88 585
R214 B.n245 B.n244 585
R215 B.n246 B.n87 585
R216 B.n248 B.n247 585
R217 B.n249 B.n86 585
R218 B.n251 B.n250 585
R219 B.n252 B.n85 585
R220 B.n254 B.n253 585
R221 B.n255 B.n84 585
R222 B.n257 B.n256 585
R223 B.n258 B.n83 585
R224 B.n260 B.n259 585
R225 B.n261 B.n82 585
R226 B.n263 B.n262 585
R227 B.n173 B.n172 585
R228 B.n171 B.n116 585
R229 B.n170 B.n169 585
R230 B.n168 B.n117 585
R231 B.n167 B.n166 585
R232 B.n165 B.n118 585
R233 B.n164 B.n163 585
R234 B.n162 B.n119 585
R235 B.n161 B.n160 585
R236 B.n159 B.n120 585
R237 B.n158 B.n157 585
R238 B.n156 B.n121 585
R239 B.n155 B.n154 585
R240 B.n153 B.n122 585
R241 B.n152 B.n151 585
R242 B.n150 B.n123 585
R243 B.n149 B.n148 585
R244 B.n147 B.n124 585
R245 B.n146 B.n145 585
R246 B.n144 B.n125 585
R247 B.n143 B.n142 585
R248 B.n141 B.n126 585
R249 B.n140 B.n139 585
R250 B.n138 B.n127 585
R251 B.n137 B.n136 585
R252 B.n135 B.n128 585
R253 B.n134 B.n133 585
R254 B.n132 B.n129 585
R255 B.n131 B.n130 585
R256 B.n2 B.n0 585
R257 B.n489 B.n1 585
R258 B.n488 B.n487 585
R259 B.n486 B.n3 585
R260 B.n485 B.n484 585
R261 B.n483 B.n4 585
R262 B.n482 B.n481 585
R263 B.n480 B.n5 585
R264 B.n479 B.n478 585
R265 B.n477 B.n6 585
R266 B.n476 B.n475 585
R267 B.n474 B.n7 585
R268 B.n473 B.n472 585
R269 B.n471 B.n8 585
R270 B.n470 B.n469 585
R271 B.n468 B.n9 585
R272 B.n467 B.n466 585
R273 B.n465 B.n10 585
R274 B.n464 B.n463 585
R275 B.n462 B.n11 585
R276 B.n461 B.n460 585
R277 B.n459 B.n12 585
R278 B.n458 B.n457 585
R279 B.n456 B.n13 585
R280 B.n455 B.n454 585
R281 B.n453 B.n14 585
R282 B.n452 B.n451 585
R283 B.n450 B.n15 585
R284 B.n449 B.n448 585
R285 B.n447 B.n16 585
R286 B.n446 B.n445 585
R287 B.n491 B.n490 585
R288 B.n172 B.n115 540.549
R289 B.n446 B.n17 540.549
R290 B.n262 B.n81 540.549
R291 B.n356 B.n51 540.549
R292 B.n94 B.t0 278.317
R293 B.n102 B.t3 278.317
R294 B.n30 B.t6 278.317
R295 B.n36 B.t9 278.317
R296 B.n172 B.n171 163.367
R297 B.n171 B.n170 163.367
R298 B.n170 B.n117 163.367
R299 B.n166 B.n117 163.367
R300 B.n166 B.n165 163.367
R301 B.n165 B.n164 163.367
R302 B.n164 B.n119 163.367
R303 B.n160 B.n119 163.367
R304 B.n160 B.n159 163.367
R305 B.n159 B.n158 163.367
R306 B.n158 B.n121 163.367
R307 B.n154 B.n121 163.367
R308 B.n154 B.n153 163.367
R309 B.n153 B.n152 163.367
R310 B.n152 B.n123 163.367
R311 B.n148 B.n123 163.367
R312 B.n148 B.n147 163.367
R313 B.n147 B.n146 163.367
R314 B.n146 B.n125 163.367
R315 B.n142 B.n125 163.367
R316 B.n142 B.n141 163.367
R317 B.n141 B.n140 163.367
R318 B.n140 B.n127 163.367
R319 B.n136 B.n127 163.367
R320 B.n136 B.n135 163.367
R321 B.n135 B.n134 163.367
R322 B.n134 B.n129 163.367
R323 B.n130 B.n129 163.367
R324 B.n130 B.n2 163.367
R325 B.n490 B.n2 163.367
R326 B.n490 B.n489 163.367
R327 B.n489 B.n488 163.367
R328 B.n488 B.n3 163.367
R329 B.n484 B.n3 163.367
R330 B.n484 B.n483 163.367
R331 B.n483 B.n482 163.367
R332 B.n482 B.n5 163.367
R333 B.n478 B.n5 163.367
R334 B.n478 B.n477 163.367
R335 B.n477 B.n476 163.367
R336 B.n476 B.n7 163.367
R337 B.n472 B.n7 163.367
R338 B.n472 B.n471 163.367
R339 B.n471 B.n470 163.367
R340 B.n470 B.n9 163.367
R341 B.n466 B.n9 163.367
R342 B.n466 B.n465 163.367
R343 B.n465 B.n464 163.367
R344 B.n464 B.n11 163.367
R345 B.n460 B.n11 163.367
R346 B.n460 B.n459 163.367
R347 B.n459 B.n458 163.367
R348 B.n458 B.n13 163.367
R349 B.n454 B.n13 163.367
R350 B.n454 B.n453 163.367
R351 B.n453 B.n452 163.367
R352 B.n452 B.n15 163.367
R353 B.n448 B.n15 163.367
R354 B.n448 B.n447 163.367
R355 B.n447 B.n446 163.367
R356 B.n176 B.n115 163.367
R357 B.n177 B.n176 163.367
R358 B.n178 B.n177 163.367
R359 B.n178 B.n113 163.367
R360 B.n182 B.n113 163.367
R361 B.n183 B.n182 163.367
R362 B.n184 B.n183 163.367
R363 B.n184 B.n111 163.367
R364 B.n188 B.n111 163.367
R365 B.n189 B.n188 163.367
R366 B.n190 B.n189 163.367
R367 B.n190 B.n109 163.367
R368 B.n194 B.n109 163.367
R369 B.n195 B.n194 163.367
R370 B.n196 B.n195 163.367
R371 B.n196 B.n107 163.367
R372 B.n200 B.n107 163.367
R373 B.n201 B.n200 163.367
R374 B.n202 B.n201 163.367
R375 B.n202 B.n105 163.367
R376 B.n206 B.n105 163.367
R377 B.n207 B.n206 163.367
R378 B.n208 B.n207 163.367
R379 B.n208 B.n101 163.367
R380 B.n213 B.n101 163.367
R381 B.n214 B.n213 163.367
R382 B.n215 B.n214 163.367
R383 B.n215 B.n99 163.367
R384 B.n219 B.n99 163.367
R385 B.n220 B.n219 163.367
R386 B.n221 B.n220 163.367
R387 B.n221 B.n97 163.367
R388 B.n225 B.n97 163.367
R389 B.n226 B.n225 163.367
R390 B.n226 B.n93 163.367
R391 B.n230 B.n93 163.367
R392 B.n231 B.n230 163.367
R393 B.n232 B.n231 163.367
R394 B.n232 B.n91 163.367
R395 B.n236 B.n91 163.367
R396 B.n237 B.n236 163.367
R397 B.n238 B.n237 163.367
R398 B.n238 B.n89 163.367
R399 B.n242 B.n89 163.367
R400 B.n243 B.n242 163.367
R401 B.n244 B.n243 163.367
R402 B.n244 B.n87 163.367
R403 B.n248 B.n87 163.367
R404 B.n249 B.n248 163.367
R405 B.n250 B.n249 163.367
R406 B.n250 B.n85 163.367
R407 B.n254 B.n85 163.367
R408 B.n255 B.n254 163.367
R409 B.n256 B.n255 163.367
R410 B.n256 B.n83 163.367
R411 B.n260 B.n83 163.367
R412 B.n261 B.n260 163.367
R413 B.n262 B.n261 163.367
R414 B.n266 B.n81 163.367
R415 B.n267 B.n266 163.367
R416 B.n268 B.n267 163.367
R417 B.n268 B.n79 163.367
R418 B.n272 B.n79 163.367
R419 B.n273 B.n272 163.367
R420 B.n274 B.n273 163.367
R421 B.n274 B.n77 163.367
R422 B.n278 B.n77 163.367
R423 B.n279 B.n278 163.367
R424 B.n280 B.n279 163.367
R425 B.n280 B.n75 163.367
R426 B.n284 B.n75 163.367
R427 B.n285 B.n284 163.367
R428 B.n286 B.n285 163.367
R429 B.n286 B.n73 163.367
R430 B.n290 B.n73 163.367
R431 B.n291 B.n290 163.367
R432 B.n292 B.n291 163.367
R433 B.n292 B.n71 163.367
R434 B.n296 B.n71 163.367
R435 B.n297 B.n296 163.367
R436 B.n298 B.n297 163.367
R437 B.n298 B.n69 163.367
R438 B.n302 B.n69 163.367
R439 B.n303 B.n302 163.367
R440 B.n304 B.n303 163.367
R441 B.n304 B.n67 163.367
R442 B.n308 B.n67 163.367
R443 B.n309 B.n308 163.367
R444 B.n310 B.n309 163.367
R445 B.n310 B.n65 163.367
R446 B.n314 B.n65 163.367
R447 B.n315 B.n314 163.367
R448 B.n316 B.n315 163.367
R449 B.n316 B.n63 163.367
R450 B.n320 B.n63 163.367
R451 B.n321 B.n320 163.367
R452 B.n322 B.n321 163.367
R453 B.n322 B.n61 163.367
R454 B.n326 B.n61 163.367
R455 B.n327 B.n326 163.367
R456 B.n328 B.n327 163.367
R457 B.n328 B.n59 163.367
R458 B.n332 B.n59 163.367
R459 B.n333 B.n332 163.367
R460 B.n334 B.n333 163.367
R461 B.n334 B.n57 163.367
R462 B.n338 B.n57 163.367
R463 B.n339 B.n338 163.367
R464 B.n340 B.n339 163.367
R465 B.n340 B.n55 163.367
R466 B.n344 B.n55 163.367
R467 B.n345 B.n344 163.367
R468 B.n346 B.n345 163.367
R469 B.n346 B.n53 163.367
R470 B.n350 B.n53 163.367
R471 B.n351 B.n350 163.367
R472 B.n352 B.n351 163.367
R473 B.n352 B.n51 163.367
R474 B.n442 B.n17 163.367
R475 B.n442 B.n441 163.367
R476 B.n441 B.n440 163.367
R477 B.n440 B.n19 163.367
R478 B.n436 B.n19 163.367
R479 B.n436 B.n435 163.367
R480 B.n435 B.n434 163.367
R481 B.n434 B.n21 163.367
R482 B.n430 B.n21 163.367
R483 B.n430 B.n429 163.367
R484 B.n429 B.n428 163.367
R485 B.n428 B.n23 163.367
R486 B.n424 B.n23 163.367
R487 B.n424 B.n423 163.367
R488 B.n423 B.n422 163.367
R489 B.n422 B.n25 163.367
R490 B.n418 B.n25 163.367
R491 B.n418 B.n417 163.367
R492 B.n417 B.n416 163.367
R493 B.n416 B.n27 163.367
R494 B.n412 B.n27 163.367
R495 B.n412 B.n411 163.367
R496 B.n411 B.n410 163.367
R497 B.n410 B.n29 163.367
R498 B.n405 B.n29 163.367
R499 B.n405 B.n404 163.367
R500 B.n404 B.n403 163.367
R501 B.n403 B.n33 163.367
R502 B.n399 B.n33 163.367
R503 B.n399 B.n398 163.367
R504 B.n398 B.n397 163.367
R505 B.n397 B.n35 163.367
R506 B.n393 B.n35 163.367
R507 B.n393 B.n392 163.367
R508 B.n392 B.n39 163.367
R509 B.n388 B.n39 163.367
R510 B.n388 B.n387 163.367
R511 B.n387 B.n386 163.367
R512 B.n386 B.n41 163.367
R513 B.n382 B.n41 163.367
R514 B.n382 B.n381 163.367
R515 B.n381 B.n380 163.367
R516 B.n380 B.n43 163.367
R517 B.n376 B.n43 163.367
R518 B.n376 B.n375 163.367
R519 B.n375 B.n374 163.367
R520 B.n374 B.n45 163.367
R521 B.n370 B.n45 163.367
R522 B.n370 B.n369 163.367
R523 B.n369 B.n368 163.367
R524 B.n368 B.n47 163.367
R525 B.n364 B.n47 163.367
R526 B.n364 B.n363 163.367
R527 B.n363 B.n362 163.367
R528 B.n362 B.n49 163.367
R529 B.n358 B.n49 163.367
R530 B.n358 B.n357 163.367
R531 B.n357 B.n356 163.367
R532 B.n94 B.t2 162.952
R533 B.n36 B.t10 162.952
R534 B.n102 B.t5 162.946
R535 B.n30 B.t7 162.946
R536 B.n95 B.t1 114.856
R537 B.n37 B.t11 114.856
R538 B.n103 B.t4 114.849
R539 B.n31 B.t8 114.849
R540 B.n96 B.n95 59.5399
R541 B.n211 B.n103 59.5399
R542 B.n407 B.n31 59.5399
R543 B.n38 B.n37 59.5399
R544 B.n95 B.n94 48.0975
R545 B.n103 B.n102 48.0975
R546 B.n31 B.n30 48.0975
R547 B.n37 B.n36 48.0975
R548 B.n445 B.n444 35.1225
R549 B.n355 B.n354 35.1225
R550 B.n264 B.n263 35.1225
R551 B.n174 B.n173 35.1225
R552 B B.n491 18.0485
R553 B.n444 B.n443 10.6151
R554 B.n443 B.n18 10.6151
R555 B.n439 B.n18 10.6151
R556 B.n439 B.n438 10.6151
R557 B.n438 B.n437 10.6151
R558 B.n437 B.n20 10.6151
R559 B.n433 B.n20 10.6151
R560 B.n433 B.n432 10.6151
R561 B.n432 B.n431 10.6151
R562 B.n431 B.n22 10.6151
R563 B.n427 B.n22 10.6151
R564 B.n427 B.n426 10.6151
R565 B.n426 B.n425 10.6151
R566 B.n425 B.n24 10.6151
R567 B.n421 B.n24 10.6151
R568 B.n421 B.n420 10.6151
R569 B.n420 B.n419 10.6151
R570 B.n419 B.n26 10.6151
R571 B.n415 B.n26 10.6151
R572 B.n415 B.n414 10.6151
R573 B.n414 B.n413 10.6151
R574 B.n413 B.n28 10.6151
R575 B.n409 B.n28 10.6151
R576 B.n409 B.n408 10.6151
R577 B.n406 B.n32 10.6151
R578 B.n402 B.n32 10.6151
R579 B.n402 B.n401 10.6151
R580 B.n401 B.n400 10.6151
R581 B.n400 B.n34 10.6151
R582 B.n396 B.n34 10.6151
R583 B.n396 B.n395 10.6151
R584 B.n395 B.n394 10.6151
R585 B.n391 B.n390 10.6151
R586 B.n390 B.n389 10.6151
R587 B.n389 B.n40 10.6151
R588 B.n385 B.n40 10.6151
R589 B.n385 B.n384 10.6151
R590 B.n384 B.n383 10.6151
R591 B.n383 B.n42 10.6151
R592 B.n379 B.n42 10.6151
R593 B.n379 B.n378 10.6151
R594 B.n378 B.n377 10.6151
R595 B.n377 B.n44 10.6151
R596 B.n373 B.n44 10.6151
R597 B.n373 B.n372 10.6151
R598 B.n372 B.n371 10.6151
R599 B.n371 B.n46 10.6151
R600 B.n367 B.n46 10.6151
R601 B.n367 B.n366 10.6151
R602 B.n366 B.n365 10.6151
R603 B.n365 B.n48 10.6151
R604 B.n361 B.n48 10.6151
R605 B.n361 B.n360 10.6151
R606 B.n360 B.n359 10.6151
R607 B.n359 B.n50 10.6151
R608 B.n355 B.n50 10.6151
R609 B.n265 B.n264 10.6151
R610 B.n265 B.n80 10.6151
R611 B.n269 B.n80 10.6151
R612 B.n270 B.n269 10.6151
R613 B.n271 B.n270 10.6151
R614 B.n271 B.n78 10.6151
R615 B.n275 B.n78 10.6151
R616 B.n276 B.n275 10.6151
R617 B.n277 B.n276 10.6151
R618 B.n277 B.n76 10.6151
R619 B.n281 B.n76 10.6151
R620 B.n282 B.n281 10.6151
R621 B.n283 B.n282 10.6151
R622 B.n283 B.n74 10.6151
R623 B.n287 B.n74 10.6151
R624 B.n288 B.n287 10.6151
R625 B.n289 B.n288 10.6151
R626 B.n289 B.n72 10.6151
R627 B.n293 B.n72 10.6151
R628 B.n294 B.n293 10.6151
R629 B.n295 B.n294 10.6151
R630 B.n295 B.n70 10.6151
R631 B.n299 B.n70 10.6151
R632 B.n300 B.n299 10.6151
R633 B.n301 B.n300 10.6151
R634 B.n301 B.n68 10.6151
R635 B.n305 B.n68 10.6151
R636 B.n306 B.n305 10.6151
R637 B.n307 B.n306 10.6151
R638 B.n307 B.n66 10.6151
R639 B.n311 B.n66 10.6151
R640 B.n312 B.n311 10.6151
R641 B.n313 B.n312 10.6151
R642 B.n313 B.n64 10.6151
R643 B.n317 B.n64 10.6151
R644 B.n318 B.n317 10.6151
R645 B.n319 B.n318 10.6151
R646 B.n319 B.n62 10.6151
R647 B.n323 B.n62 10.6151
R648 B.n324 B.n323 10.6151
R649 B.n325 B.n324 10.6151
R650 B.n325 B.n60 10.6151
R651 B.n329 B.n60 10.6151
R652 B.n330 B.n329 10.6151
R653 B.n331 B.n330 10.6151
R654 B.n331 B.n58 10.6151
R655 B.n335 B.n58 10.6151
R656 B.n336 B.n335 10.6151
R657 B.n337 B.n336 10.6151
R658 B.n337 B.n56 10.6151
R659 B.n341 B.n56 10.6151
R660 B.n342 B.n341 10.6151
R661 B.n343 B.n342 10.6151
R662 B.n343 B.n54 10.6151
R663 B.n347 B.n54 10.6151
R664 B.n348 B.n347 10.6151
R665 B.n349 B.n348 10.6151
R666 B.n349 B.n52 10.6151
R667 B.n353 B.n52 10.6151
R668 B.n354 B.n353 10.6151
R669 B.n175 B.n174 10.6151
R670 B.n175 B.n114 10.6151
R671 B.n179 B.n114 10.6151
R672 B.n180 B.n179 10.6151
R673 B.n181 B.n180 10.6151
R674 B.n181 B.n112 10.6151
R675 B.n185 B.n112 10.6151
R676 B.n186 B.n185 10.6151
R677 B.n187 B.n186 10.6151
R678 B.n187 B.n110 10.6151
R679 B.n191 B.n110 10.6151
R680 B.n192 B.n191 10.6151
R681 B.n193 B.n192 10.6151
R682 B.n193 B.n108 10.6151
R683 B.n197 B.n108 10.6151
R684 B.n198 B.n197 10.6151
R685 B.n199 B.n198 10.6151
R686 B.n199 B.n106 10.6151
R687 B.n203 B.n106 10.6151
R688 B.n204 B.n203 10.6151
R689 B.n205 B.n204 10.6151
R690 B.n205 B.n104 10.6151
R691 B.n209 B.n104 10.6151
R692 B.n210 B.n209 10.6151
R693 B.n212 B.n100 10.6151
R694 B.n216 B.n100 10.6151
R695 B.n217 B.n216 10.6151
R696 B.n218 B.n217 10.6151
R697 B.n218 B.n98 10.6151
R698 B.n222 B.n98 10.6151
R699 B.n223 B.n222 10.6151
R700 B.n224 B.n223 10.6151
R701 B.n228 B.n227 10.6151
R702 B.n229 B.n228 10.6151
R703 B.n229 B.n92 10.6151
R704 B.n233 B.n92 10.6151
R705 B.n234 B.n233 10.6151
R706 B.n235 B.n234 10.6151
R707 B.n235 B.n90 10.6151
R708 B.n239 B.n90 10.6151
R709 B.n240 B.n239 10.6151
R710 B.n241 B.n240 10.6151
R711 B.n241 B.n88 10.6151
R712 B.n245 B.n88 10.6151
R713 B.n246 B.n245 10.6151
R714 B.n247 B.n246 10.6151
R715 B.n247 B.n86 10.6151
R716 B.n251 B.n86 10.6151
R717 B.n252 B.n251 10.6151
R718 B.n253 B.n252 10.6151
R719 B.n253 B.n84 10.6151
R720 B.n257 B.n84 10.6151
R721 B.n258 B.n257 10.6151
R722 B.n259 B.n258 10.6151
R723 B.n259 B.n82 10.6151
R724 B.n263 B.n82 10.6151
R725 B.n173 B.n116 10.6151
R726 B.n169 B.n116 10.6151
R727 B.n169 B.n168 10.6151
R728 B.n168 B.n167 10.6151
R729 B.n167 B.n118 10.6151
R730 B.n163 B.n118 10.6151
R731 B.n163 B.n162 10.6151
R732 B.n162 B.n161 10.6151
R733 B.n161 B.n120 10.6151
R734 B.n157 B.n120 10.6151
R735 B.n157 B.n156 10.6151
R736 B.n156 B.n155 10.6151
R737 B.n155 B.n122 10.6151
R738 B.n151 B.n122 10.6151
R739 B.n151 B.n150 10.6151
R740 B.n150 B.n149 10.6151
R741 B.n149 B.n124 10.6151
R742 B.n145 B.n124 10.6151
R743 B.n145 B.n144 10.6151
R744 B.n144 B.n143 10.6151
R745 B.n143 B.n126 10.6151
R746 B.n139 B.n126 10.6151
R747 B.n139 B.n138 10.6151
R748 B.n138 B.n137 10.6151
R749 B.n137 B.n128 10.6151
R750 B.n133 B.n128 10.6151
R751 B.n133 B.n132 10.6151
R752 B.n132 B.n131 10.6151
R753 B.n131 B.n0 10.6151
R754 B.n487 B.n1 10.6151
R755 B.n487 B.n486 10.6151
R756 B.n486 B.n485 10.6151
R757 B.n485 B.n4 10.6151
R758 B.n481 B.n4 10.6151
R759 B.n481 B.n480 10.6151
R760 B.n480 B.n479 10.6151
R761 B.n479 B.n6 10.6151
R762 B.n475 B.n6 10.6151
R763 B.n475 B.n474 10.6151
R764 B.n474 B.n473 10.6151
R765 B.n473 B.n8 10.6151
R766 B.n469 B.n8 10.6151
R767 B.n469 B.n468 10.6151
R768 B.n468 B.n467 10.6151
R769 B.n467 B.n10 10.6151
R770 B.n463 B.n10 10.6151
R771 B.n463 B.n462 10.6151
R772 B.n462 B.n461 10.6151
R773 B.n461 B.n12 10.6151
R774 B.n457 B.n12 10.6151
R775 B.n457 B.n456 10.6151
R776 B.n456 B.n455 10.6151
R777 B.n455 B.n14 10.6151
R778 B.n451 B.n14 10.6151
R779 B.n451 B.n450 10.6151
R780 B.n450 B.n449 10.6151
R781 B.n449 B.n16 10.6151
R782 B.n445 B.n16 10.6151
R783 B.n407 B.n406 6.5566
R784 B.n394 B.n38 6.5566
R785 B.n212 B.n211 6.5566
R786 B.n224 B.n96 6.5566
R787 B.n408 B.n407 4.05904
R788 B.n391 B.n38 4.05904
R789 B.n211 B.n210 4.05904
R790 B.n227 B.n96 4.05904
R791 B.n491 B.n0 2.81026
R792 B.n491 B.n1 2.81026
R793 VN.n0 VN.t3 106.466
R794 VN.n1 VN.t1 106.466
R795 VN.n0 VN.t2 105.838
R796 VN.n1 VN.t0 105.838
R797 VN VN.n1 46.7716
R798 VN VN.n0 5.96475
R799 VDD2.n2 VDD2.n0 125.434
R800 VDD2.n2 VDD2.n1 89.8404
R801 VDD2.n1 VDD2.t3 5.12747
R802 VDD2.n1 VDD2.t2 5.12747
R803 VDD2.n0 VDD2.t0 5.12747
R804 VDD2.n0 VDD2.t1 5.12747
R805 VDD2 VDD2.n2 0.0586897
C0 VTAIL w_n2458_n2236# 2.67476f
C1 B w_n2458_n2236# 7.11207f
C2 w_n2458_n2236# VDD2 1.25707f
C3 VDD1 VP 2.78816f
C4 VN VTAIL 2.7532f
C5 VN B 0.957554f
C6 B VTAIL 2.92327f
C7 VN VDD2 2.57171f
C8 VP w_n2458_n2236# 4.29912f
C9 VTAIL VDD2 3.97099f
C10 B VDD2 1.07602f
C11 VDD1 w_n2458_n2236# 1.21101f
C12 VN VP 4.8195f
C13 VTAIL VP 2.76731f
C14 VN VDD1 0.148755f
C15 B VP 1.47794f
C16 VTAIL VDD1 3.9198f
C17 VP VDD2 0.365833f
C18 B VDD1 1.03126f
C19 VN w_n2458_n2236# 3.98427f
C20 VDD1 VDD2 0.919287f
C21 VDD2 VSUBS 0.7323f
C22 VDD1 VSUBS 4.718259f
C23 VTAIL VSUBS 0.681542f
C24 VN VSUBS 5.07621f
C25 VP VSUBS 1.73251f
C26 B VSUBS 3.405947f
C27 w_n2458_n2236# VSUBS 68.5192f
C28 VDD2.t0 VSUBS 0.137894f
C29 VDD2.t1 VSUBS 0.137894f
C30 VDD2.n0 VSUBS 1.36166f
C31 VDD2.t3 VSUBS 0.137894f
C32 VDD2.t2 VSUBS 0.137894f
C33 VDD2.n1 VSUBS 0.926639f
C34 VDD2.n2 VSUBS 3.5646f
C35 VN.t3 VSUBS 1.86226f
C36 VN.t2 VSUBS 1.85729f
C37 VN.n0 VSUBS 1.24618f
C38 VN.t1 VSUBS 1.86226f
C39 VN.t0 VSUBS 1.85729f
C40 VN.n1 VSUBS 3.09142f
C41 B.n0 VSUBS 0.005245f
C42 B.n1 VSUBS 0.005245f
C43 B.n2 VSUBS 0.008294f
C44 B.n3 VSUBS 0.008294f
C45 B.n4 VSUBS 0.008294f
C46 B.n5 VSUBS 0.008294f
C47 B.n6 VSUBS 0.008294f
C48 B.n7 VSUBS 0.008294f
C49 B.n8 VSUBS 0.008294f
C50 B.n9 VSUBS 0.008294f
C51 B.n10 VSUBS 0.008294f
C52 B.n11 VSUBS 0.008294f
C53 B.n12 VSUBS 0.008294f
C54 B.n13 VSUBS 0.008294f
C55 B.n14 VSUBS 0.008294f
C56 B.n15 VSUBS 0.008294f
C57 B.n16 VSUBS 0.008294f
C58 B.n17 VSUBS 0.020604f
C59 B.n18 VSUBS 0.008294f
C60 B.n19 VSUBS 0.008294f
C61 B.n20 VSUBS 0.008294f
C62 B.n21 VSUBS 0.008294f
C63 B.n22 VSUBS 0.008294f
C64 B.n23 VSUBS 0.008294f
C65 B.n24 VSUBS 0.008294f
C66 B.n25 VSUBS 0.008294f
C67 B.n26 VSUBS 0.008294f
C68 B.n27 VSUBS 0.008294f
C69 B.n28 VSUBS 0.008294f
C70 B.n29 VSUBS 0.008294f
C71 B.t8 VSUBS 0.221789f
C72 B.t7 VSUBS 0.242493f
C73 B.t6 VSUBS 0.754229f
C74 B.n30 VSUBS 0.137093f
C75 B.n31 VSUBS 0.081973f
C76 B.n32 VSUBS 0.008294f
C77 B.n33 VSUBS 0.008294f
C78 B.n34 VSUBS 0.008294f
C79 B.n35 VSUBS 0.008294f
C80 B.t11 VSUBS 0.221788f
C81 B.t10 VSUBS 0.242492f
C82 B.t9 VSUBS 0.754229f
C83 B.n36 VSUBS 0.137094f
C84 B.n37 VSUBS 0.081974f
C85 B.n38 VSUBS 0.019217f
C86 B.n39 VSUBS 0.008294f
C87 B.n40 VSUBS 0.008294f
C88 B.n41 VSUBS 0.008294f
C89 B.n42 VSUBS 0.008294f
C90 B.n43 VSUBS 0.008294f
C91 B.n44 VSUBS 0.008294f
C92 B.n45 VSUBS 0.008294f
C93 B.n46 VSUBS 0.008294f
C94 B.n47 VSUBS 0.008294f
C95 B.n48 VSUBS 0.008294f
C96 B.n49 VSUBS 0.008294f
C97 B.n50 VSUBS 0.008294f
C98 B.n51 VSUBS 0.020137f
C99 B.n52 VSUBS 0.008294f
C100 B.n53 VSUBS 0.008294f
C101 B.n54 VSUBS 0.008294f
C102 B.n55 VSUBS 0.008294f
C103 B.n56 VSUBS 0.008294f
C104 B.n57 VSUBS 0.008294f
C105 B.n58 VSUBS 0.008294f
C106 B.n59 VSUBS 0.008294f
C107 B.n60 VSUBS 0.008294f
C108 B.n61 VSUBS 0.008294f
C109 B.n62 VSUBS 0.008294f
C110 B.n63 VSUBS 0.008294f
C111 B.n64 VSUBS 0.008294f
C112 B.n65 VSUBS 0.008294f
C113 B.n66 VSUBS 0.008294f
C114 B.n67 VSUBS 0.008294f
C115 B.n68 VSUBS 0.008294f
C116 B.n69 VSUBS 0.008294f
C117 B.n70 VSUBS 0.008294f
C118 B.n71 VSUBS 0.008294f
C119 B.n72 VSUBS 0.008294f
C120 B.n73 VSUBS 0.008294f
C121 B.n74 VSUBS 0.008294f
C122 B.n75 VSUBS 0.008294f
C123 B.n76 VSUBS 0.008294f
C124 B.n77 VSUBS 0.008294f
C125 B.n78 VSUBS 0.008294f
C126 B.n79 VSUBS 0.008294f
C127 B.n80 VSUBS 0.008294f
C128 B.n81 VSUBS 0.020137f
C129 B.n82 VSUBS 0.008294f
C130 B.n83 VSUBS 0.008294f
C131 B.n84 VSUBS 0.008294f
C132 B.n85 VSUBS 0.008294f
C133 B.n86 VSUBS 0.008294f
C134 B.n87 VSUBS 0.008294f
C135 B.n88 VSUBS 0.008294f
C136 B.n89 VSUBS 0.008294f
C137 B.n90 VSUBS 0.008294f
C138 B.n91 VSUBS 0.008294f
C139 B.n92 VSUBS 0.008294f
C140 B.n93 VSUBS 0.008294f
C141 B.t1 VSUBS 0.221788f
C142 B.t2 VSUBS 0.242492f
C143 B.t0 VSUBS 0.754229f
C144 B.n94 VSUBS 0.137094f
C145 B.n95 VSUBS 0.081974f
C146 B.n96 VSUBS 0.019217f
C147 B.n97 VSUBS 0.008294f
C148 B.n98 VSUBS 0.008294f
C149 B.n99 VSUBS 0.008294f
C150 B.n100 VSUBS 0.008294f
C151 B.n101 VSUBS 0.008294f
C152 B.t4 VSUBS 0.221789f
C153 B.t5 VSUBS 0.242493f
C154 B.t3 VSUBS 0.754229f
C155 B.n102 VSUBS 0.137093f
C156 B.n103 VSUBS 0.081973f
C157 B.n104 VSUBS 0.008294f
C158 B.n105 VSUBS 0.008294f
C159 B.n106 VSUBS 0.008294f
C160 B.n107 VSUBS 0.008294f
C161 B.n108 VSUBS 0.008294f
C162 B.n109 VSUBS 0.008294f
C163 B.n110 VSUBS 0.008294f
C164 B.n111 VSUBS 0.008294f
C165 B.n112 VSUBS 0.008294f
C166 B.n113 VSUBS 0.008294f
C167 B.n114 VSUBS 0.008294f
C168 B.n115 VSUBS 0.020604f
C169 B.n116 VSUBS 0.008294f
C170 B.n117 VSUBS 0.008294f
C171 B.n118 VSUBS 0.008294f
C172 B.n119 VSUBS 0.008294f
C173 B.n120 VSUBS 0.008294f
C174 B.n121 VSUBS 0.008294f
C175 B.n122 VSUBS 0.008294f
C176 B.n123 VSUBS 0.008294f
C177 B.n124 VSUBS 0.008294f
C178 B.n125 VSUBS 0.008294f
C179 B.n126 VSUBS 0.008294f
C180 B.n127 VSUBS 0.008294f
C181 B.n128 VSUBS 0.008294f
C182 B.n129 VSUBS 0.008294f
C183 B.n130 VSUBS 0.008294f
C184 B.n131 VSUBS 0.008294f
C185 B.n132 VSUBS 0.008294f
C186 B.n133 VSUBS 0.008294f
C187 B.n134 VSUBS 0.008294f
C188 B.n135 VSUBS 0.008294f
C189 B.n136 VSUBS 0.008294f
C190 B.n137 VSUBS 0.008294f
C191 B.n138 VSUBS 0.008294f
C192 B.n139 VSUBS 0.008294f
C193 B.n140 VSUBS 0.008294f
C194 B.n141 VSUBS 0.008294f
C195 B.n142 VSUBS 0.008294f
C196 B.n143 VSUBS 0.008294f
C197 B.n144 VSUBS 0.008294f
C198 B.n145 VSUBS 0.008294f
C199 B.n146 VSUBS 0.008294f
C200 B.n147 VSUBS 0.008294f
C201 B.n148 VSUBS 0.008294f
C202 B.n149 VSUBS 0.008294f
C203 B.n150 VSUBS 0.008294f
C204 B.n151 VSUBS 0.008294f
C205 B.n152 VSUBS 0.008294f
C206 B.n153 VSUBS 0.008294f
C207 B.n154 VSUBS 0.008294f
C208 B.n155 VSUBS 0.008294f
C209 B.n156 VSUBS 0.008294f
C210 B.n157 VSUBS 0.008294f
C211 B.n158 VSUBS 0.008294f
C212 B.n159 VSUBS 0.008294f
C213 B.n160 VSUBS 0.008294f
C214 B.n161 VSUBS 0.008294f
C215 B.n162 VSUBS 0.008294f
C216 B.n163 VSUBS 0.008294f
C217 B.n164 VSUBS 0.008294f
C218 B.n165 VSUBS 0.008294f
C219 B.n166 VSUBS 0.008294f
C220 B.n167 VSUBS 0.008294f
C221 B.n168 VSUBS 0.008294f
C222 B.n169 VSUBS 0.008294f
C223 B.n170 VSUBS 0.008294f
C224 B.n171 VSUBS 0.008294f
C225 B.n172 VSUBS 0.020137f
C226 B.n173 VSUBS 0.020137f
C227 B.n174 VSUBS 0.020604f
C228 B.n175 VSUBS 0.008294f
C229 B.n176 VSUBS 0.008294f
C230 B.n177 VSUBS 0.008294f
C231 B.n178 VSUBS 0.008294f
C232 B.n179 VSUBS 0.008294f
C233 B.n180 VSUBS 0.008294f
C234 B.n181 VSUBS 0.008294f
C235 B.n182 VSUBS 0.008294f
C236 B.n183 VSUBS 0.008294f
C237 B.n184 VSUBS 0.008294f
C238 B.n185 VSUBS 0.008294f
C239 B.n186 VSUBS 0.008294f
C240 B.n187 VSUBS 0.008294f
C241 B.n188 VSUBS 0.008294f
C242 B.n189 VSUBS 0.008294f
C243 B.n190 VSUBS 0.008294f
C244 B.n191 VSUBS 0.008294f
C245 B.n192 VSUBS 0.008294f
C246 B.n193 VSUBS 0.008294f
C247 B.n194 VSUBS 0.008294f
C248 B.n195 VSUBS 0.008294f
C249 B.n196 VSUBS 0.008294f
C250 B.n197 VSUBS 0.008294f
C251 B.n198 VSUBS 0.008294f
C252 B.n199 VSUBS 0.008294f
C253 B.n200 VSUBS 0.008294f
C254 B.n201 VSUBS 0.008294f
C255 B.n202 VSUBS 0.008294f
C256 B.n203 VSUBS 0.008294f
C257 B.n204 VSUBS 0.008294f
C258 B.n205 VSUBS 0.008294f
C259 B.n206 VSUBS 0.008294f
C260 B.n207 VSUBS 0.008294f
C261 B.n208 VSUBS 0.008294f
C262 B.n209 VSUBS 0.008294f
C263 B.n210 VSUBS 0.005733f
C264 B.n211 VSUBS 0.019217f
C265 B.n212 VSUBS 0.006709f
C266 B.n213 VSUBS 0.008294f
C267 B.n214 VSUBS 0.008294f
C268 B.n215 VSUBS 0.008294f
C269 B.n216 VSUBS 0.008294f
C270 B.n217 VSUBS 0.008294f
C271 B.n218 VSUBS 0.008294f
C272 B.n219 VSUBS 0.008294f
C273 B.n220 VSUBS 0.008294f
C274 B.n221 VSUBS 0.008294f
C275 B.n222 VSUBS 0.008294f
C276 B.n223 VSUBS 0.008294f
C277 B.n224 VSUBS 0.006709f
C278 B.n225 VSUBS 0.008294f
C279 B.n226 VSUBS 0.008294f
C280 B.n227 VSUBS 0.005733f
C281 B.n228 VSUBS 0.008294f
C282 B.n229 VSUBS 0.008294f
C283 B.n230 VSUBS 0.008294f
C284 B.n231 VSUBS 0.008294f
C285 B.n232 VSUBS 0.008294f
C286 B.n233 VSUBS 0.008294f
C287 B.n234 VSUBS 0.008294f
C288 B.n235 VSUBS 0.008294f
C289 B.n236 VSUBS 0.008294f
C290 B.n237 VSUBS 0.008294f
C291 B.n238 VSUBS 0.008294f
C292 B.n239 VSUBS 0.008294f
C293 B.n240 VSUBS 0.008294f
C294 B.n241 VSUBS 0.008294f
C295 B.n242 VSUBS 0.008294f
C296 B.n243 VSUBS 0.008294f
C297 B.n244 VSUBS 0.008294f
C298 B.n245 VSUBS 0.008294f
C299 B.n246 VSUBS 0.008294f
C300 B.n247 VSUBS 0.008294f
C301 B.n248 VSUBS 0.008294f
C302 B.n249 VSUBS 0.008294f
C303 B.n250 VSUBS 0.008294f
C304 B.n251 VSUBS 0.008294f
C305 B.n252 VSUBS 0.008294f
C306 B.n253 VSUBS 0.008294f
C307 B.n254 VSUBS 0.008294f
C308 B.n255 VSUBS 0.008294f
C309 B.n256 VSUBS 0.008294f
C310 B.n257 VSUBS 0.008294f
C311 B.n258 VSUBS 0.008294f
C312 B.n259 VSUBS 0.008294f
C313 B.n260 VSUBS 0.008294f
C314 B.n261 VSUBS 0.008294f
C315 B.n262 VSUBS 0.020604f
C316 B.n263 VSUBS 0.020604f
C317 B.n264 VSUBS 0.020137f
C318 B.n265 VSUBS 0.008294f
C319 B.n266 VSUBS 0.008294f
C320 B.n267 VSUBS 0.008294f
C321 B.n268 VSUBS 0.008294f
C322 B.n269 VSUBS 0.008294f
C323 B.n270 VSUBS 0.008294f
C324 B.n271 VSUBS 0.008294f
C325 B.n272 VSUBS 0.008294f
C326 B.n273 VSUBS 0.008294f
C327 B.n274 VSUBS 0.008294f
C328 B.n275 VSUBS 0.008294f
C329 B.n276 VSUBS 0.008294f
C330 B.n277 VSUBS 0.008294f
C331 B.n278 VSUBS 0.008294f
C332 B.n279 VSUBS 0.008294f
C333 B.n280 VSUBS 0.008294f
C334 B.n281 VSUBS 0.008294f
C335 B.n282 VSUBS 0.008294f
C336 B.n283 VSUBS 0.008294f
C337 B.n284 VSUBS 0.008294f
C338 B.n285 VSUBS 0.008294f
C339 B.n286 VSUBS 0.008294f
C340 B.n287 VSUBS 0.008294f
C341 B.n288 VSUBS 0.008294f
C342 B.n289 VSUBS 0.008294f
C343 B.n290 VSUBS 0.008294f
C344 B.n291 VSUBS 0.008294f
C345 B.n292 VSUBS 0.008294f
C346 B.n293 VSUBS 0.008294f
C347 B.n294 VSUBS 0.008294f
C348 B.n295 VSUBS 0.008294f
C349 B.n296 VSUBS 0.008294f
C350 B.n297 VSUBS 0.008294f
C351 B.n298 VSUBS 0.008294f
C352 B.n299 VSUBS 0.008294f
C353 B.n300 VSUBS 0.008294f
C354 B.n301 VSUBS 0.008294f
C355 B.n302 VSUBS 0.008294f
C356 B.n303 VSUBS 0.008294f
C357 B.n304 VSUBS 0.008294f
C358 B.n305 VSUBS 0.008294f
C359 B.n306 VSUBS 0.008294f
C360 B.n307 VSUBS 0.008294f
C361 B.n308 VSUBS 0.008294f
C362 B.n309 VSUBS 0.008294f
C363 B.n310 VSUBS 0.008294f
C364 B.n311 VSUBS 0.008294f
C365 B.n312 VSUBS 0.008294f
C366 B.n313 VSUBS 0.008294f
C367 B.n314 VSUBS 0.008294f
C368 B.n315 VSUBS 0.008294f
C369 B.n316 VSUBS 0.008294f
C370 B.n317 VSUBS 0.008294f
C371 B.n318 VSUBS 0.008294f
C372 B.n319 VSUBS 0.008294f
C373 B.n320 VSUBS 0.008294f
C374 B.n321 VSUBS 0.008294f
C375 B.n322 VSUBS 0.008294f
C376 B.n323 VSUBS 0.008294f
C377 B.n324 VSUBS 0.008294f
C378 B.n325 VSUBS 0.008294f
C379 B.n326 VSUBS 0.008294f
C380 B.n327 VSUBS 0.008294f
C381 B.n328 VSUBS 0.008294f
C382 B.n329 VSUBS 0.008294f
C383 B.n330 VSUBS 0.008294f
C384 B.n331 VSUBS 0.008294f
C385 B.n332 VSUBS 0.008294f
C386 B.n333 VSUBS 0.008294f
C387 B.n334 VSUBS 0.008294f
C388 B.n335 VSUBS 0.008294f
C389 B.n336 VSUBS 0.008294f
C390 B.n337 VSUBS 0.008294f
C391 B.n338 VSUBS 0.008294f
C392 B.n339 VSUBS 0.008294f
C393 B.n340 VSUBS 0.008294f
C394 B.n341 VSUBS 0.008294f
C395 B.n342 VSUBS 0.008294f
C396 B.n343 VSUBS 0.008294f
C397 B.n344 VSUBS 0.008294f
C398 B.n345 VSUBS 0.008294f
C399 B.n346 VSUBS 0.008294f
C400 B.n347 VSUBS 0.008294f
C401 B.n348 VSUBS 0.008294f
C402 B.n349 VSUBS 0.008294f
C403 B.n350 VSUBS 0.008294f
C404 B.n351 VSUBS 0.008294f
C405 B.n352 VSUBS 0.008294f
C406 B.n353 VSUBS 0.008294f
C407 B.n354 VSUBS 0.021048f
C408 B.n355 VSUBS 0.019692f
C409 B.n356 VSUBS 0.020604f
C410 B.n357 VSUBS 0.008294f
C411 B.n358 VSUBS 0.008294f
C412 B.n359 VSUBS 0.008294f
C413 B.n360 VSUBS 0.008294f
C414 B.n361 VSUBS 0.008294f
C415 B.n362 VSUBS 0.008294f
C416 B.n363 VSUBS 0.008294f
C417 B.n364 VSUBS 0.008294f
C418 B.n365 VSUBS 0.008294f
C419 B.n366 VSUBS 0.008294f
C420 B.n367 VSUBS 0.008294f
C421 B.n368 VSUBS 0.008294f
C422 B.n369 VSUBS 0.008294f
C423 B.n370 VSUBS 0.008294f
C424 B.n371 VSUBS 0.008294f
C425 B.n372 VSUBS 0.008294f
C426 B.n373 VSUBS 0.008294f
C427 B.n374 VSUBS 0.008294f
C428 B.n375 VSUBS 0.008294f
C429 B.n376 VSUBS 0.008294f
C430 B.n377 VSUBS 0.008294f
C431 B.n378 VSUBS 0.008294f
C432 B.n379 VSUBS 0.008294f
C433 B.n380 VSUBS 0.008294f
C434 B.n381 VSUBS 0.008294f
C435 B.n382 VSUBS 0.008294f
C436 B.n383 VSUBS 0.008294f
C437 B.n384 VSUBS 0.008294f
C438 B.n385 VSUBS 0.008294f
C439 B.n386 VSUBS 0.008294f
C440 B.n387 VSUBS 0.008294f
C441 B.n388 VSUBS 0.008294f
C442 B.n389 VSUBS 0.008294f
C443 B.n390 VSUBS 0.008294f
C444 B.n391 VSUBS 0.005733f
C445 B.n392 VSUBS 0.008294f
C446 B.n393 VSUBS 0.008294f
C447 B.n394 VSUBS 0.006709f
C448 B.n395 VSUBS 0.008294f
C449 B.n396 VSUBS 0.008294f
C450 B.n397 VSUBS 0.008294f
C451 B.n398 VSUBS 0.008294f
C452 B.n399 VSUBS 0.008294f
C453 B.n400 VSUBS 0.008294f
C454 B.n401 VSUBS 0.008294f
C455 B.n402 VSUBS 0.008294f
C456 B.n403 VSUBS 0.008294f
C457 B.n404 VSUBS 0.008294f
C458 B.n405 VSUBS 0.008294f
C459 B.n406 VSUBS 0.006709f
C460 B.n407 VSUBS 0.019217f
C461 B.n408 VSUBS 0.005733f
C462 B.n409 VSUBS 0.008294f
C463 B.n410 VSUBS 0.008294f
C464 B.n411 VSUBS 0.008294f
C465 B.n412 VSUBS 0.008294f
C466 B.n413 VSUBS 0.008294f
C467 B.n414 VSUBS 0.008294f
C468 B.n415 VSUBS 0.008294f
C469 B.n416 VSUBS 0.008294f
C470 B.n417 VSUBS 0.008294f
C471 B.n418 VSUBS 0.008294f
C472 B.n419 VSUBS 0.008294f
C473 B.n420 VSUBS 0.008294f
C474 B.n421 VSUBS 0.008294f
C475 B.n422 VSUBS 0.008294f
C476 B.n423 VSUBS 0.008294f
C477 B.n424 VSUBS 0.008294f
C478 B.n425 VSUBS 0.008294f
C479 B.n426 VSUBS 0.008294f
C480 B.n427 VSUBS 0.008294f
C481 B.n428 VSUBS 0.008294f
C482 B.n429 VSUBS 0.008294f
C483 B.n430 VSUBS 0.008294f
C484 B.n431 VSUBS 0.008294f
C485 B.n432 VSUBS 0.008294f
C486 B.n433 VSUBS 0.008294f
C487 B.n434 VSUBS 0.008294f
C488 B.n435 VSUBS 0.008294f
C489 B.n436 VSUBS 0.008294f
C490 B.n437 VSUBS 0.008294f
C491 B.n438 VSUBS 0.008294f
C492 B.n439 VSUBS 0.008294f
C493 B.n440 VSUBS 0.008294f
C494 B.n441 VSUBS 0.008294f
C495 B.n442 VSUBS 0.008294f
C496 B.n443 VSUBS 0.008294f
C497 B.n444 VSUBS 0.020604f
C498 B.n445 VSUBS 0.020137f
C499 B.n446 VSUBS 0.020137f
C500 B.n447 VSUBS 0.008294f
C501 B.n448 VSUBS 0.008294f
C502 B.n449 VSUBS 0.008294f
C503 B.n450 VSUBS 0.008294f
C504 B.n451 VSUBS 0.008294f
C505 B.n452 VSUBS 0.008294f
C506 B.n453 VSUBS 0.008294f
C507 B.n454 VSUBS 0.008294f
C508 B.n455 VSUBS 0.008294f
C509 B.n456 VSUBS 0.008294f
C510 B.n457 VSUBS 0.008294f
C511 B.n458 VSUBS 0.008294f
C512 B.n459 VSUBS 0.008294f
C513 B.n460 VSUBS 0.008294f
C514 B.n461 VSUBS 0.008294f
C515 B.n462 VSUBS 0.008294f
C516 B.n463 VSUBS 0.008294f
C517 B.n464 VSUBS 0.008294f
C518 B.n465 VSUBS 0.008294f
C519 B.n466 VSUBS 0.008294f
C520 B.n467 VSUBS 0.008294f
C521 B.n468 VSUBS 0.008294f
C522 B.n469 VSUBS 0.008294f
C523 B.n470 VSUBS 0.008294f
C524 B.n471 VSUBS 0.008294f
C525 B.n472 VSUBS 0.008294f
C526 B.n473 VSUBS 0.008294f
C527 B.n474 VSUBS 0.008294f
C528 B.n475 VSUBS 0.008294f
C529 B.n476 VSUBS 0.008294f
C530 B.n477 VSUBS 0.008294f
C531 B.n478 VSUBS 0.008294f
C532 B.n479 VSUBS 0.008294f
C533 B.n480 VSUBS 0.008294f
C534 B.n481 VSUBS 0.008294f
C535 B.n482 VSUBS 0.008294f
C536 B.n483 VSUBS 0.008294f
C537 B.n484 VSUBS 0.008294f
C538 B.n485 VSUBS 0.008294f
C539 B.n486 VSUBS 0.008294f
C540 B.n487 VSUBS 0.008294f
C541 B.n488 VSUBS 0.008294f
C542 B.n489 VSUBS 0.008294f
C543 B.n490 VSUBS 0.008294f
C544 B.n491 VSUBS 0.018781f
C545 VDD1.t0 VSUBS 0.13786f
C546 VDD1.t3 VSUBS 0.13786f
C547 VDD1.n0 VSUBS 0.926838f
C548 VDD1.t1 VSUBS 0.13786f
C549 VDD1.t2 VSUBS 0.13786f
C550 VDD1.n1 VSUBS 1.38184f
C551 VTAIL.t1 VSUBS 1.09929f
C552 VTAIL.n0 VSUBS 0.711684f
C553 VTAIL.t4 VSUBS 1.09929f
C554 VTAIL.n1 VSUBS 0.79885f
C555 VTAIL.t3 VSUBS 1.09929f
C556 VTAIL.n2 VSUBS 1.77758f
C557 VTAIL.t7 VSUBS 1.09929f
C558 VTAIL.n3 VSUBS 1.77757f
C559 VTAIL.t2 VSUBS 1.09929f
C560 VTAIL.n4 VSUBS 0.798844f
C561 VTAIL.t5 VSUBS 1.09929f
C562 VTAIL.n5 VSUBS 0.798844f
C563 VTAIL.t6 VSUBS 1.09929f
C564 VTAIL.n6 VSUBS 1.77758f
C565 VTAIL.t0 VSUBS 1.09929f
C566 VTAIL.n7 VSUBS 1.68038f
C567 VP.n0 VSUBS 0.05999f
C568 VP.t1 VSUBS 1.6469f
C569 VP.n1 VSUBS 0.036752f
C570 VP.n2 VSUBS 0.05999f
C571 VP.t2 VSUBS 1.6469f
C572 VP.t0 VSUBS 1.93106f
C573 VP.t3 VSUBS 1.93622f
C574 VP.n3 VSUBS 3.19038f
C575 VP.n4 VSUBS 2.13994f
C576 VP.n5 VSUBS 0.749127f
C577 VP.n6 VSUBS 0.062722f
C578 VP.n7 VSUBS 0.089964f
C579 VP.n8 VSUBS 0.045505f
C580 VP.n9 VSUBS 0.045505f
C581 VP.n10 VSUBS 0.045505f
C582 VP.n11 VSUBS 0.089964f
C583 VP.n12 VSUBS 0.062722f
C584 VP.n13 VSUBS 0.749127f
C585 VP.n14 VSUBS 0.065986f
.ends

