* NGSPICE file created from diff_pair_sample_0464.ext - technology: sky130A

.subckt diff_pair_sample_0464 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=2.5116 ps=13.66 w=6.44 l=2.88
X1 VTAIL.t10 VN.t1 VDD2.t4 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=1.0626 ps=6.77 w=6.44 l=2.88
X2 B.t11 B.t9 B.t10 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=0 ps=0 w=6.44 l=2.88
X3 VDD1.t5 VP.t0 VTAIL.t2 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=2.5116 ps=13.66 w=6.44 l=2.88
X4 VDD2.t3 VN.t2 VTAIL.t6 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=1.0626 ps=6.77 w=6.44 l=2.88
X5 VDD1.t4 VP.t1 VTAIL.t3 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=1.0626 ps=6.77 w=6.44 l=2.88
X6 B.t8 B.t6 B.t7 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=0 ps=0 w=6.44 l=2.88
X7 VDD2.t2 VN.t3 VTAIL.t11 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=2.5116 ps=13.66 w=6.44 l=2.88
X8 VTAIL.t4 VP.t2 VDD1.t3 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=1.0626 ps=6.77 w=6.44 l=2.88
X9 VDD1.t2 VP.t3 VTAIL.t5 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=1.0626 ps=6.77 w=6.44 l=2.88
X10 VDD1.t1 VP.t4 VTAIL.t0 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=2.5116 ps=13.66 w=6.44 l=2.88
X11 B.t5 B.t3 B.t4 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=0 ps=0 w=6.44 l=2.88
X12 VTAIL.t1 VP.t5 VDD1.t0 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=1.0626 ps=6.77 w=6.44 l=2.88
X13 VDD2.t1 VN.t4 VTAIL.t9 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=1.0626 ps=6.77 w=6.44 l=2.88
X14 B.t2 B.t0 B.t1 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=2.5116 pd=13.66 as=0 ps=0 w=6.44 l=2.88
X15 VTAIL.t7 VN.t5 VDD2.t0 w_n3538_n2256# sky130_fd_pr__pfet_01v8 ad=1.0626 pd=6.77 as=1.0626 ps=6.77 w=6.44 l=2.88
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t3 85.789
R13 VN.n4 VN.t2 85.789
R14 VN.n15 VN.n0 67.6211
R15 VN.n31 VN.n16 67.6211
R16 VN.n5 VN.n4 61.7085
R17 VN.n21 VN.n20 61.7085
R18 VN.n11 VN.n2 54.6242
R19 VN.n27 VN.n18 54.6242
R20 VN.n5 VN.t1 53.8908
R21 VN.n0 VN.t0 53.8908
R22 VN.n21 VN.t5 53.8908
R23 VN.n16 VN.t4 53.8908
R24 VN VN.n31 45.858
R25 VN.n12 VN.n11 26.5299
R26 VN.n28 VN.n27 26.5299
R27 VN.n7 VN.n6 24.5923
R28 VN.n7 VN.n2 24.5923
R29 VN.n13 VN.n12 24.5923
R30 VN.n23 VN.n18 24.5923
R31 VN.n23 VN.n22 24.5923
R32 VN.n29 VN.n28 24.5923
R33 VN.n13 VN.n0 22.625
R34 VN.n29 VN.n16 22.625
R35 VN.n6 VN.n5 12.2964
R36 VN.n22 VN.n21 12.2964
R37 VN.n4 VN.n3 5.34748
R38 VN.n20 VN.n19 5.34748
R39 VN.n31 VN.n30 0.354861
R40 VN.n15 VN.n14 0.354861
R41 VN VN.n15 0.267071
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n7 VTAIL.t11 80.1485
R53 VTAIL.n11 VTAIL.t8 80.1484
R54 VTAIL.n2 VTAIL.t0 80.1484
R55 VTAIL.n10 VTAIL.t2 80.1484
R56 VTAIL.n9 VTAIL.n8 75.1012
R57 VTAIL.n6 VTAIL.n5 75.1012
R58 VTAIL.n1 VTAIL.n0 75.101
R59 VTAIL.n4 VTAIL.n3 75.101
R60 VTAIL.n6 VTAIL.n4 23.4531
R61 VTAIL.n11 VTAIL.n10 20.6858
R62 VTAIL.n0 VTAIL.t6 5.04786
R63 VTAIL.n0 VTAIL.t10 5.04786
R64 VTAIL.n3 VTAIL.t5 5.04786
R65 VTAIL.n3 VTAIL.t4 5.04786
R66 VTAIL.n8 VTAIL.t3 5.04786
R67 VTAIL.n8 VTAIL.t1 5.04786
R68 VTAIL.n5 VTAIL.t9 5.04786
R69 VTAIL.n5 VTAIL.t7 5.04786
R70 VTAIL.n7 VTAIL.n6 2.76774
R71 VTAIL.n10 VTAIL.n9 2.76774
R72 VTAIL.n4 VTAIL.n2 2.76774
R73 VTAIL VTAIL.n11 2.01774
R74 VTAIL.n9 VTAIL.n7 1.85395
R75 VTAIL.n2 VTAIL.n1 1.85395
R76 VTAIL VTAIL.n1 0.7505
R77 VDD2.n1 VDD2.t3 98.8472
R78 VDD2.n2 VDD2.t1 96.8273
R79 VDD2.n1 VDD2.n0 92.4162
R80 VDD2 VDD2.n3 92.4134
R81 VDD2.n2 VDD2.n1 38.2606
R82 VDD2.n3 VDD2.t0 5.04786
R83 VDD2.n3 VDD2.t2 5.04786
R84 VDD2.n0 VDD2.t4 5.04786
R85 VDD2.n0 VDD2.t5 5.04786
R86 VDD2 VDD2.n2 2.13412
R87 B.n463 B.n462 585
R88 B.n464 B.n59 585
R89 B.n466 B.n465 585
R90 B.n467 B.n58 585
R91 B.n469 B.n468 585
R92 B.n470 B.n57 585
R93 B.n472 B.n471 585
R94 B.n473 B.n56 585
R95 B.n475 B.n474 585
R96 B.n476 B.n55 585
R97 B.n478 B.n477 585
R98 B.n479 B.n54 585
R99 B.n481 B.n480 585
R100 B.n482 B.n53 585
R101 B.n484 B.n483 585
R102 B.n485 B.n52 585
R103 B.n487 B.n486 585
R104 B.n488 B.n51 585
R105 B.n490 B.n489 585
R106 B.n491 B.n50 585
R107 B.n493 B.n492 585
R108 B.n494 B.n49 585
R109 B.n496 B.n495 585
R110 B.n497 B.n45 585
R111 B.n499 B.n498 585
R112 B.n500 B.n44 585
R113 B.n502 B.n501 585
R114 B.n503 B.n43 585
R115 B.n505 B.n504 585
R116 B.n506 B.n42 585
R117 B.n508 B.n507 585
R118 B.n509 B.n41 585
R119 B.n511 B.n510 585
R120 B.n512 B.n40 585
R121 B.n514 B.n513 585
R122 B.n516 B.n37 585
R123 B.n518 B.n517 585
R124 B.n519 B.n36 585
R125 B.n521 B.n520 585
R126 B.n522 B.n35 585
R127 B.n524 B.n523 585
R128 B.n525 B.n34 585
R129 B.n527 B.n526 585
R130 B.n528 B.n33 585
R131 B.n530 B.n529 585
R132 B.n531 B.n32 585
R133 B.n533 B.n532 585
R134 B.n534 B.n31 585
R135 B.n536 B.n535 585
R136 B.n537 B.n30 585
R137 B.n539 B.n538 585
R138 B.n540 B.n29 585
R139 B.n542 B.n541 585
R140 B.n543 B.n28 585
R141 B.n545 B.n544 585
R142 B.n546 B.n27 585
R143 B.n548 B.n547 585
R144 B.n549 B.n26 585
R145 B.n551 B.n550 585
R146 B.n552 B.n25 585
R147 B.n461 B.n60 585
R148 B.n460 B.n459 585
R149 B.n458 B.n61 585
R150 B.n457 B.n456 585
R151 B.n455 B.n62 585
R152 B.n454 B.n453 585
R153 B.n452 B.n63 585
R154 B.n451 B.n450 585
R155 B.n449 B.n64 585
R156 B.n448 B.n447 585
R157 B.n446 B.n65 585
R158 B.n445 B.n444 585
R159 B.n443 B.n66 585
R160 B.n442 B.n441 585
R161 B.n440 B.n67 585
R162 B.n439 B.n438 585
R163 B.n437 B.n68 585
R164 B.n436 B.n435 585
R165 B.n434 B.n69 585
R166 B.n433 B.n432 585
R167 B.n431 B.n70 585
R168 B.n430 B.n429 585
R169 B.n428 B.n71 585
R170 B.n427 B.n426 585
R171 B.n425 B.n72 585
R172 B.n424 B.n423 585
R173 B.n422 B.n73 585
R174 B.n421 B.n420 585
R175 B.n419 B.n74 585
R176 B.n418 B.n417 585
R177 B.n416 B.n75 585
R178 B.n415 B.n414 585
R179 B.n413 B.n76 585
R180 B.n412 B.n411 585
R181 B.n410 B.n77 585
R182 B.n409 B.n408 585
R183 B.n407 B.n78 585
R184 B.n406 B.n405 585
R185 B.n404 B.n79 585
R186 B.n403 B.n402 585
R187 B.n401 B.n80 585
R188 B.n400 B.n399 585
R189 B.n398 B.n81 585
R190 B.n397 B.n396 585
R191 B.n395 B.n82 585
R192 B.n394 B.n393 585
R193 B.n392 B.n83 585
R194 B.n391 B.n390 585
R195 B.n389 B.n84 585
R196 B.n388 B.n387 585
R197 B.n386 B.n85 585
R198 B.n385 B.n384 585
R199 B.n383 B.n86 585
R200 B.n382 B.n381 585
R201 B.n380 B.n87 585
R202 B.n379 B.n378 585
R203 B.n377 B.n88 585
R204 B.n376 B.n375 585
R205 B.n374 B.n89 585
R206 B.n373 B.n372 585
R207 B.n371 B.n90 585
R208 B.n370 B.n369 585
R209 B.n368 B.n91 585
R210 B.n367 B.n366 585
R211 B.n365 B.n92 585
R212 B.n364 B.n363 585
R213 B.n362 B.n93 585
R214 B.n361 B.n360 585
R215 B.n359 B.n94 585
R216 B.n358 B.n357 585
R217 B.n356 B.n95 585
R218 B.n355 B.n354 585
R219 B.n353 B.n96 585
R220 B.n352 B.n351 585
R221 B.n350 B.n97 585
R222 B.n349 B.n348 585
R223 B.n347 B.n98 585
R224 B.n346 B.n345 585
R225 B.n344 B.n99 585
R226 B.n343 B.n342 585
R227 B.n341 B.n100 585
R228 B.n340 B.n339 585
R229 B.n338 B.n101 585
R230 B.n337 B.n336 585
R231 B.n335 B.n102 585
R232 B.n334 B.n333 585
R233 B.n332 B.n103 585
R234 B.n331 B.n330 585
R235 B.n329 B.n104 585
R236 B.n328 B.n327 585
R237 B.n326 B.n105 585
R238 B.n325 B.n324 585
R239 B.n323 B.n106 585
R240 B.n232 B.n231 585
R241 B.n233 B.n140 585
R242 B.n235 B.n234 585
R243 B.n236 B.n139 585
R244 B.n238 B.n237 585
R245 B.n239 B.n138 585
R246 B.n241 B.n240 585
R247 B.n242 B.n137 585
R248 B.n244 B.n243 585
R249 B.n245 B.n136 585
R250 B.n247 B.n246 585
R251 B.n248 B.n135 585
R252 B.n250 B.n249 585
R253 B.n251 B.n134 585
R254 B.n253 B.n252 585
R255 B.n254 B.n133 585
R256 B.n256 B.n255 585
R257 B.n257 B.n132 585
R258 B.n259 B.n258 585
R259 B.n260 B.n131 585
R260 B.n262 B.n261 585
R261 B.n263 B.n130 585
R262 B.n265 B.n264 585
R263 B.n266 B.n129 585
R264 B.n268 B.n267 585
R265 B.n270 B.n126 585
R266 B.n272 B.n271 585
R267 B.n273 B.n125 585
R268 B.n275 B.n274 585
R269 B.n276 B.n124 585
R270 B.n278 B.n277 585
R271 B.n279 B.n123 585
R272 B.n281 B.n280 585
R273 B.n282 B.n122 585
R274 B.n284 B.n283 585
R275 B.n286 B.n285 585
R276 B.n287 B.n118 585
R277 B.n289 B.n288 585
R278 B.n290 B.n117 585
R279 B.n292 B.n291 585
R280 B.n293 B.n116 585
R281 B.n295 B.n294 585
R282 B.n296 B.n115 585
R283 B.n298 B.n297 585
R284 B.n299 B.n114 585
R285 B.n301 B.n300 585
R286 B.n302 B.n113 585
R287 B.n304 B.n303 585
R288 B.n305 B.n112 585
R289 B.n307 B.n306 585
R290 B.n308 B.n111 585
R291 B.n310 B.n309 585
R292 B.n311 B.n110 585
R293 B.n313 B.n312 585
R294 B.n314 B.n109 585
R295 B.n316 B.n315 585
R296 B.n317 B.n108 585
R297 B.n319 B.n318 585
R298 B.n320 B.n107 585
R299 B.n322 B.n321 585
R300 B.n230 B.n141 585
R301 B.n229 B.n228 585
R302 B.n227 B.n142 585
R303 B.n226 B.n225 585
R304 B.n224 B.n143 585
R305 B.n223 B.n222 585
R306 B.n221 B.n144 585
R307 B.n220 B.n219 585
R308 B.n218 B.n145 585
R309 B.n217 B.n216 585
R310 B.n215 B.n146 585
R311 B.n214 B.n213 585
R312 B.n212 B.n147 585
R313 B.n211 B.n210 585
R314 B.n209 B.n148 585
R315 B.n208 B.n207 585
R316 B.n206 B.n149 585
R317 B.n205 B.n204 585
R318 B.n203 B.n150 585
R319 B.n202 B.n201 585
R320 B.n200 B.n151 585
R321 B.n199 B.n198 585
R322 B.n197 B.n152 585
R323 B.n196 B.n195 585
R324 B.n194 B.n153 585
R325 B.n193 B.n192 585
R326 B.n191 B.n154 585
R327 B.n190 B.n189 585
R328 B.n188 B.n155 585
R329 B.n187 B.n186 585
R330 B.n185 B.n156 585
R331 B.n184 B.n183 585
R332 B.n182 B.n157 585
R333 B.n181 B.n180 585
R334 B.n179 B.n158 585
R335 B.n178 B.n177 585
R336 B.n176 B.n159 585
R337 B.n175 B.n174 585
R338 B.n173 B.n160 585
R339 B.n172 B.n171 585
R340 B.n170 B.n161 585
R341 B.n169 B.n168 585
R342 B.n167 B.n162 585
R343 B.n166 B.n165 585
R344 B.n164 B.n163 585
R345 B.n2 B.n0 585
R346 B.n621 B.n1 585
R347 B.n620 B.n619 585
R348 B.n618 B.n3 585
R349 B.n617 B.n616 585
R350 B.n615 B.n4 585
R351 B.n614 B.n613 585
R352 B.n612 B.n5 585
R353 B.n611 B.n610 585
R354 B.n609 B.n6 585
R355 B.n608 B.n607 585
R356 B.n606 B.n7 585
R357 B.n605 B.n604 585
R358 B.n603 B.n8 585
R359 B.n602 B.n601 585
R360 B.n600 B.n9 585
R361 B.n599 B.n598 585
R362 B.n597 B.n10 585
R363 B.n596 B.n595 585
R364 B.n594 B.n11 585
R365 B.n593 B.n592 585
R366 B.n591 B.n12 585
R367 B.n590 B.n589 585
R368 B.n588 B.n13 585
R369 B.n587 B.n586 585
R370 B.n585 B.n14 585
R371 B.n584 B.n583 585
R372 B.n582 B.n15 585
R373 B.n581 B.n580 585
R374 B.n579 B.n16 585
R375 B.n578 B.n577 585
R376 B.n576 B.n17 585
R377 B.n575 B.n574 585
R378 B.n573 B.n18 585
R379 B.n572 B.n571 585
R380 B.n570 B.n19 585
R381 B.n569 B.n568 585
R382 B.n567 B.n20 585
R383 B.n566 B.n565 585
R384 B.n564 B.n21 585
R385 B.n563 B.n562 585
R386 B.n561 B.n22 585
R387 B.n560 B.n559 585
R388 B.n558 B.n23 585
R389 B.n557 B.n556 585
R390 B.n555 B.n24 585
R391 B.n554 B.n553 585
R392 B.n623 B.n622 585
R393 B.n231 B.n230 487.695
R394 B.n554 B.n25 487.695
R395 B.n321 B.n106 487.695
R396 B.n463 B.n60 487.695
R397 B.n119 B.t9 262.325
R398 B.n127 B.t3 262.325
R399 B.n38 B.t6 262.325
R400 B.n46 B.t0 262.325
R401 B.n119 B.t11 178.97
R402 B.n46 B.t1 178.97
R403 B.n127 B.t5 178.964
R404 B.n38 B.t7 178.964
R405 B.n230 B.n229 163.367
R406 B.n229 B.n142 163.367
R407 B.n225 B.n142 163.367
R408 B.n225 B.n224 163.367
R409 B.n224 B.n223 163.367
R410 B.n223 B.n144 163.367
R411 B.n219 B.n144 163.367
R412 B.n219 B.n218 163.367
R413 B.n218 B.n217 163.367
R414 B.n217 B.n146 163.367
R415 B.n213 B.n146 163.367
R416 B.n213 B.n212 163.367
R417 B.n212 B.n211 163.367
R418 B.n211 B.n148 163.367
R419 B.n207 B.n148 163.367
R420 B.n207 B.n206 163.367
R421 B.n206 B.n205 163.367
R422 B.n205 B.n150 163.367
R423 B.n201 B.n150 163.367
R424 B.n201 B.n200 163.367
R425 B.n200 B.n199 163.367
R426 B.n199 B.n152 163.367
R427 B.n195 B.n152 163.367
R428 B.n195 B.n194 163.367
R429 B.n194 B.n193 163.367
R430 B.n193 B.n154 163.367
R431 B.n189 B.n154 163.367
R432 B.n189 B.n188 163.367
R433 B.n188 B.n187 163.367
R434 B.n187 B.n156 163.367
R435 B.n183 B.n156 163.367
R436 B.n183 B.n182 163.367
R437 B.n182 B.n181 163.367
R438 B.n181 B.n158 163.367
R439 B.n177 B.n158 163.367
R440 B.n177 B.n176 163.367
R441 B.n176 B.n175 163.367
R442 B.n175 B.n160 163.367
R443 B.n171 B.n160 163.367
R444 B.n171 B.n170 163.367
R445 B.n170 B.n169 163.367
R446 B.n169 B.n162 163.367
R447 B.n165 B.n162 163.367
R448 B.n165 B.n164 163.367
R449 B.n164 B.n2 163.367
R450 B.n622 B.n2 163.367
R451 B.n622 B.n621 163.367
R452 B.n621 B.n620 163.367
R453 B.n620 B.n3 163.367
R454 B.n616 B.n3 163.367
R455 B.n616 B.n615 163.367
R456 B.n615 B.n614 163.367
R457 B.n614 B.n5 163.367
R458 B.n610 B.n5 163.367
R459 B.n610 B.n609 163.367
R460 B.n609 B.n608 163.367
R461 B.n608 B.n7 163.367
R462 B.n604 B.n7 163.367
R463 B.n604 B.n603 163.367
R464 B.n603 B.n602 163.367
R465 B.n602 B.n9 163.367
R466 B.n598 B.n9 163.367
R467 B.n598 B.n597 163.367
R468 B.n597 B.n596 163.367
R469 B.n596 B.n11 163.367
R470 B.n592 B.n11 163.367
R471 B.n592 B.n591 163.367
R472 B.n591 B.n590 163.367
R473 B.n590 B.n13 163.367
R474 B.n586 B.n13 163.367
R475 B.n586 B.n585 163.367
R476 B.n585 B.n584 163.367
R477 B.n584 B.n15 163.367
R478 B.n580 B.n15 163.367
R479 B.n580 B.n579 163.367
R480 B.n579 B.n578 163.367
R481 B.n578 B.n17 163.367
R482 B.n574 B.n17 163.367
R483 B.n574 B.n573 163.367
R484 B.n573 B.n572 163.367
R485 B.n572 B.n19 163.367
R486 B.n568 B.n19 163.367
R487 B.n568 B.n567 163.367
R488 B.n567 B.n566 163.367
R489 B.n566 B.n21 163.367
R490 B.n562 B.n21 163.367
R491 B.n562 B.n561 163.367
R492 B.n561 B.n560 163.367
R493 B.n560 B.n23 163.367
R494 B.n556 B.n23 163.367
R495 B.n556 B.n555 163.367
R496 B.n555 B.n554 163.367
R497 B.n231 B.n140 163.367
R498 B.n235 B.n140 163.367
R499 B.n236 B.n235 163.367
R500 B.n237 B.n236 163.367
R501 B.n237 B.n138 163.367
R502 B.n241 B.n138 163.367
R503 B.n242 B.n241 163.367
R504 B.n243 B.n242 163.367
R505 B.n243 B.n136 163.367
R506 B.n247 B.n136 163.367
R507 B.n248 B.n247 163.367
R508 B.n249 B.n248 163.367
R509 B.n249 B.n134 163.367
R510 B.n253 B.n134 163.367
R511 B.n254 B.n253 163.367
R512 B.n255 B.n254 163.367
R513 B.n255 B.n132 163.367
R514 B.n259 B.n132 163.367
R515 B.n260 B.n259 163.367
R516 B.n261 B.n260 163.367
R517 B.n261 B.n130 163.367
R518 B.n265 B.n130 163.367
R519 B.n266 B.n265 163.367
R520 B.n267 B.n266 163.367
R521 B.n267 B.n126 163.367
R522 B.n272 B.n126 163.367
R523 B.n273 B.n272 163.367
R524 B.n274 B.n273 163.367
R525 B.n274 B.n124 163.367
R526 B.n278 B.n124 163.367
R527 B.n279 B.n278 163.367
R528 B.n280 B.n279 163.367
R529 B.n280 B.n122 163.367
R530 B.n284 B.n122 163.367
R531 B.n285 B.n284 163.367
R532 B.n285 B.n118 163.367
R533 B.n289 B.n118 163.367
R534 B.n290 B.n289 163.367
R535 B.n291 B.n290 163.367
R536 B.n291 B.n116 163.367
R537 B.n295 B.n116 163.367
R538 B.n296 B.n295 163.367
R539 B.n297 B.n296 163.367
R540 B.n297 B.n114 163.367
R541 B.n301 B.n114 163.367
R542 B.n302 B.n301 163.367
R543 B.n303 B.n302 163.367
R544 B.n303 B.n112 163.367
R545 B.n307 B.n112 163.367
R546 B.n308 B.n307 163.367
R547 B.n309 B.n308 163.367
R548 B.n309 B.n110 163.367
R549 B.n313 B.n110 163.367
R550 B.n314 B.n313 163.367
R551 B.n315 B.n314 163.367
R552 B.n315 B.n108 163.367
R553 B.n319 B.n108 163.367
R554 B.n320 B.n319 163.367
R555 B.n321 B.n320 163.367
R556 B.n325 B.n106 163.367
R557 B.n326 B.n325 163.367
R558 B.n327 B.n326 163.367
R559 B.n327 B.n104 163.367
R560 B.n331 B.n104 163.367
R561 B.n332 B.n331 163.367
R562 B.n333 B.n332 163.367
R563 B.n333 B.n102 163.367
R564 B.n337 B.n102 163.367
R565 B.n338 B.n337 163.367
R566 B.n339 B.n338 163.367
R567 B.n339 B.n100 163.367
R568 B.n343 B.n100 163.367
R569 B.n344 B.n343 163.367
R570 B.n345 B.n344 163.367
R571 B.n345 B.n98 163.367
R572 B.n349 B.n98 163.367
R573 B.n350 B.n349 163.367
R574 B.n351 B.n350 163.367
R575 B.n351 B.n96 163.367
R576 B.n355 B.n96 163.367
R577 B.n356 B.n355 163.367
R578 B.n357 B.n356 163.367
R579 B.n357 B.n94 163.367
R580 B.n361 B.n94 163.367
R581 B.n362 B.n361 163.367
R582 B.n363 B.n362 163.367
R583 B.n363 B.n92 163.367
R584 B.n367 B.n92 163.367
R585 B.n368 B.n367 163.367
R586 B.n369 B.n368 163.367
R587 B.n369 B.n90 163.367
R588 B.n373 B.n90 163.367
R589 B.n374 B.n373 163.367
R590 B.n375 B.n374 163.367
R591 B.n375 B.n88 163.367
R592 B.n379 B.n88 163.367
R593 B.n380 B.n379 163.367
R594 B.n381 B.n380 163.367
R595 B.n381 B.n86 163.367
R596 B.n385 B.n86 163.367
R597 B.n386 B.n385 163.367
R598 B.n387 B.n386 163.367
R599 B.n387 B.n84 163.367
R600 B.n391 B.n84 163.367
R601 B.n392 B.n391 163.367
R602 B.n393 B.n392 163.367
R603 B.n393 B.n82 163.367
R604 B.n397 B.n82 163.367
R605 B.n398 B.n397 163.367
R606 B.n399 B.n398 163.367
R607 B.n399 B.n80 163.367
R608 B.n403 B.n80 163.367
R609 B.n404 B.n403 163.367
R610 B.n405 B.n404 163.367
R611 B.n405 B.n78 163.367
R612 B.n409 B.n78 163.367
R613 B.n410 B.n409 163.367
R614 B.n411 B.n410 163.367
R615 B.n411 B.n76 163.367
R616 B.n415 B.n76 163.367
R617 B.n416 B.n415 163.367
R618 B.n417 B.n416 163.367
R619 B.n417 B.n74 163.367
R620 B.n421 B.n74 163.367
R621 B.n422 B.n421 163.367
R622 B.n423 B.n422 163.367
R623 B.n423 B.n72 163.367
R624 B.n427 B.n72 163.367
R625 B.n428 B.n427 163.367
R626 B.n429 B.n428 163.367
R627 B.n429 B.n70 163.367
R628 B.n433 B.n70 163.367
R629 B.n434 B.n433 163.367
R630 B.n435 B.n434 163.367
R631 B.n435 B.n68 163.367
R632 B.n439 B.n68 163.367
R633 B.n440 B.n439 163.367
R634 B.n441 B.n440 163.367
R635 B.n441 B.n66 163.367
R636 B.n445 B.n66 163.367
R637 B.n446 B.n445 163.367
R638 B.n447 B.n446 163.367
R639 B.n447 B.n64 163.367
R640 B.n451 B.n64 163.367
R641 B.n452 B.n451 163.367
R642 B.n453 B.n452 163.367
R643 B.n453 B.n62 163.367
R644 B.n457 B.n62 163.367
R645 B.n458 B.n457 163.367
R646 B.n459 B.n458 163.367
R647 B.n459 B.n60 163.367
R648 B.n550 B.n25 163.367
R649 B.n550 B.n549 163.367
R650 B.n549 B.n548 163.367
R651 B.n548 B.n27 163.367
R652 B.n544 B.n27 163.367
R653 B.n544 B.n543 163.367
R654 B.n543 B.n542 163.367
R655 B.n542 B.n29 163.367
R656 B.n538 B.n29 163.367
R657 B.n538 B.n537 163.367
R658 B.n537 B.n536 163.367
R659 B.n536 B.n31 163.367
R660 B.n532 B.n31 163.367
R661 B.n532 B.n531 163.367
R662 B.n531 B.n530 163.367
R663 B.n530 B.n33 163.367
R664 B.n526 B.n33 163.367
R665 B.n526 B.n525 163.367
R666 B.n525 B.n524 163.367
R667 B.n524 B.n35 163.367
R668 B.n520 B.n35 163.367
R669 B.n520 B.n519 163.367
R670 B.n519 B.n518 163.367
R671 B.n518 B.n37 163.367
R672 B.n513 B.n37 163.367
R673 B.n513 B.n512 163.367
R674 B.n512 B.n511 163.367
R675 B.n511 B.n41 163.367
R676 B.n507 B.n41 163.367
R677 B.n507 B.n506 163.367
R678 B.n506 B.n505 163.367
R679 B.n505 B.n43 163.367
R680 B.n501 B.n43 163.367
R681 B.n501 B.n500 163.367
R682 B.n500 B.n499 163.367
R683 B.n499 B.n45 163.367
R684 B.n495 B.n45 163.367
R685 B.n495 B.n494 163.367
R686 B.n494 B.n493 163.367
R687 B.n493 B.n50 163.367
R688 B.n489 B.n50 163.367
R689 B.n489 B.n488 163.367
R690 B.n488 B.n487 163.367
R691 B.n487 B.n52 163.367
R692 B.n483 B.n52 163.367
R693 B.n483 B.n482 163.367
R694 B.n482 B.n481 163.367
R695 B.n481 B.n54 163.367
R696 B.n477 B.n54 163.367
R697 B.n477 B.n476 163.367
R698 B.n476 B.n475 163.367
R699 B.n475 B.n56 163.367
R700 B.n471 B.n56 163.367
R701 B.n471 B.n470 163.367
R702 B.n470 B.n469 163.367
R703 B.n469 B.n58 163.367
R704 B.n465 B.n58 163.367
R705 B.n465 B.n464 163.367
R706 B.n464 B.n463 163.367
R707 B.n120 B.t10 116.716
R708 B.n47 B.t2 116.716
R709 B.n128 B.t4 116.709
R710 B.n39 B.t8 116.709
R711 B.n120 B.n119 62.255
R712 B.n128 B.n127 62.255
R713 B.n39 B.n38 62.255
R714 B.n47 B.n46 62.255
R715 B.n121 B.n120 59.5399
R716 B.n269 B.n128 59.5399
R717 B.n515 B.n39 59.5399
R718 B.n48 B.n47 59.5399
R719 B.n553 B.n552 31.6883
R720 B.n462 B.n461 31.6883
R721 B.n323 B.n322 31.6883
R722 B.n232 B.n141 31.6883
R723 B B.n623 18.0485
R724 B.n552 B.n551 10.6151
R725 B.n551 B.n26 10.6151
R726 B.n547 B.n26 10.6151
R727 B.n547 B.n546 10.6151
R728 B.n546 B.n545 10.6151
R729 B.n545 B.n28 10.6151
R730 B.n541 B.n28 10.6151
R731 B.n541 B.n540 10.6151
R732 B.n540 B.n539 10.6151
R733 B.n539 B.n30 10.6151
R734 B.n535 B.n30 10.6151
R735 B.n535 B.n534 10.6151
R736 B.n534 B.n533 10.6151
R737 B.n533 B.n32 10.6151
R738 B.n529 B.n32 10.6151
R739 B.n529 B.n528 10.6151
R740 B.n528 B.n527 10.6151
R741 B.n527 B.n34 10.6151
R742 B.n523 B.n34 10.6151
R743 B.n523 B.n522 10.6151
R744 B.n522 B.n521 10.6151
R745 B.n521 B.n36 10.6151
R746 B.n517 B.n36 10.6151
R747 B.n517 B.n516 10.6151
R748 B.n514 B.n40 10.6151
R749 B.n510 B.n40 10.6151
R750 B.n510 B.n509 10.6151
R751 B.n509 B.n508 10.6151
R752 B.n508 B.n42 10.6151
R753 B.n504 B.n42 10.6151
R754 B.n504 B.n503 10.6151
R755 B.n503 B.n502 10.6151
R756 B.n502 B.n44 10.6151
R757 B.n498 B.n497 10.6151
R758 B.n497 B.n496 10.6151
R759 B.n496 B.n49 10.6151
R760 B.n492 B.n49 10.6151
R761 B.n492 B.n491 10.6151
R762 B.n491 B.n490 10.6151
R763 B.n490 B.n51 10.6151
R764 B.n486 B.n51 10.6151
R765 B.n486 B.n485 10.6151
R766 B.n485 B.n484 10.6151
R767 B.n484 B.n53 10.6151
R768 B.n480 B.n53 10.6151
R769 B.n480 B.n479 10.6151
R770 B.n479 B.n478 10.6151
R771 B.n478 B.n55 10.6151
R772 B.n474 B.n55 10.6151
R773 B.n474 B.n473 10.6151
R774 B.n473 B.n472 10.6151
R775 B.n472 B.n57 10.6151
R776 B.n468 B.n57 10.6151
R777 B.n468 B.n467 10.6151
R778 B.n467 B.n466 10.6151
R779 B.n466 B.n59 10.6151
R780 B.n462 B.n59 10.6151
R781 B.n324 B.n323 10.6151
R782 B.n324 B.n105 10.6151
R783 B.n328 B.n105 10.6151
R784 B.n329 B.n328 10.6151
R785 B.n330 B.n329 10.6151
R786 B.n330 B.n103 10.6151
R787 B.n334 B.n103 10.6151
R788 B.n335 B.n334 10.6151
R789 B.n336 B.n335 10.6151
R790 B.n336 B.n101 10.6151
R791 B.n340 B.n101 10.6151
R792 B.n341 B.n340 10.6151
R793 B.n342 B.n341 10.6151
R794 B.n342 B.n99 10.6151
R795 B.n346 B.n99 10.6151
R796 B.n347 B.n346 10.6151
R797 B.n348 B.n347 10.6151
R798 B.n348 B.n97 10.6151
R799 B.n352 B.n97 10.6151
R800 B.n353 B.n352 10.6151
R801 B.n354 B.n353 10.6151
R802 B.n354 B.n95 10.6151
R803 B.n358 B.n95 10.6151
R804 B.n359 B.n358 10.6151
R805 B.n360 B.n359 10.6151
R806 B.n360 B.n93 10.6151
R807 B.n364 B.n93 10.6151
R808 B.n365 B.n364 10.6151
R809 B.n366 B.n365 10.6151
R810 B.n366 B.n91 10.6151
R811 B.n370 B.n91 10.6151
R812 B.n371 B.n370 10.6151
R813 B.n372 B.n371 10.6151
R814 B.n372 B.n89 10.6151
R815 B.n376 B.n89 10.6151
R816 B.n377 B.n376 10.6151
R817 B.n378 B.n377 10.6151
R818 B.n378 B.n87 10.6151
R819 B.n382 B.n87 10.6151
R820 B.n383 B.n382 10.6151
R821 B.n384 B.n383 10.6151
R822 B.n384 B.n85 10.6151
R823 B.n388 B.n85 10.6151
R824 B.n389 B.n388 10.6151
R825 B.n390 B.n389 10.6151
R826 B.n390 B.n83 10.6151
R827 B.n394 B.n83 10.6151
R828 B.n395 B.n394 10.6151
R829 B.n396 B.n395 10.6151
R830 B.n396 B.n81 10.6151
R831 B.n400 B.n81 10.6151
R832 B.n401 B.n400 10.6151
R833 B.n402 B.n401 10.6151
R834 B.n402 B.n79 10.6151
R835 B.n406 B.n79 10.6151
R836 B.n407 B.n406 10.6151
R837 B.n408 B.n407 10.6151
R838 B.n408 B.n77 10.6151
R839 B.n412 B.n77 10.6151
R840 B.n413 B.n412 10.6151
R841 B.n414 B.n413 10.6151
R842 B.n414 B.n75 10.6151
R843 B.n418 B.n75 10.6151
R844 B.n419 B.n418 10.6151
R845 B.n420 B.n419 10.6151
R846 B.n420 B.n73 10.6151
R847 B.n424 B.n73 10.6151
R848 B.n425 B.n424 10.6151
R849 B.n426 B.n425 10.6151
R850 B.n426 B.n71 10.6151
R851 B.n430 B.n71 10.6151
R852 B.n431 B.n430 10.6151
R853 B.n432 B.n431 10.6151
R854 B.n432 B.n69 10.6151
R855 B.n436 B.n69 10.6151
R856 B.n437 B.n436 10.6151
R857 B.n438 B.n437 10.6151
R858 B.n438 B.n67 10.6151
R859 B.n442 B.n67 10.6151
R860 B.n443 B.n442 10.6151
R861 B.n444 B.n443 10.6151
R862 B.n444 B.n65 10.6151
R863 B.n448 B.n65 10.6151
R864 B.n449 B.n448 10.6151
R865 B.n450 B.n449 10.6151
R866 B.n450 B.n63 10.6151
R867 B.n454 B.n63 10.6151
R868 B.n455 B.n454 10.6151
R869 B.n456 B.n455 10.6151
R870 B.n456 B.n61 10.6151
R871 B.n460 B.n61 10.6151
R872 B.n461 B.n460 10.6151
R873 B.n233 B.n232 10.6151
R874 B.n234 B.n233 10.6151
R875 B.n234 B.n139 10.6151
R876 B.n238 B.n139 10.6151
R877 B.n239 B.n238 10.6151
R878 B.n240 B.n239 10.6151
R879 B.n240 B.n137 10.6151
R880 B.n244 B.n137 10.6151
R881 B.n245 B.n244 10.6151
R882 B.n246 B.n245 10.6151
R883 B.n246 B.n135 10.6151
R884 B.n250 B.n135 10.6151
R885 B.n251 B.n250 10.6151
R886 B.n252 B.n251 10.6151
R887 B.n252 B.n133 10.6151
R888 B.n256 B.n133 10.6151
R889 B.n257 B.n256 10.6151
R890 B.n258 B.n257 10.6151
R891 B.n258 B.n131 10.6151
R892 B.n262 B.n131 10.6151
R893 B.n263 B.n262 10.6151
R894 B.n264 B.n263 10.6151
R895 B.n264 B.n129 10.6151
R896 B.n268 B.n129 10.6151
R897 B.n271 B.n270 10.6151
R898 B.n271 B.n125 10.6151
R899 B.n275 B.n125 10.6151
R900 B.n276 B.n275 10.6151
R901 B.n277 B.n276 10.6151
R902 B.n277 B.n123 10.6151
R903 B.n281 B.n123 10.6151
R904 B.n282 B.n281 10.6151
R905 B.n283 B.n282 10.6151
R906 B.n287 B.n286 10.6151
R907 B.n288 B.n287 10.6151
R908 B.n288 B.n117 10.6151
R909 B.n292 B.n117 10.6151
R910 B.n293 B.n292 10.6151
R911 B.n294 B.n293 10.6151
R912 B.n294 B.n115 10.6151
R913 B.n298 B.n115 10.6151
R914 B.n299 B.n298 10.6151
R915 B.n300 B.n299 10.6151
R916 B.n300 B.n113 10.6151
R917 B.n304 B.n113 10.6151
R918 B.n305 B.n304 10.6151
R919 B.n306 B.n305 10.6151
R920 B.n306 B.n111 10.6151
R921 B.n310 B.n111 10.6151
R922 B.n311 B.n310 10.6151
R923 B.n312 B.n311 10.6151
R924 B.n312 B.n109 10.6151
R925 B.n316 B.n109 10.6151
R926 B.n317 B.n316 10.6151
R927 B.n318 B.n317 10.6151
R928 B.n318 B.n107 10.6151
R929 B.n322 B.n107 10.6151
R930 B.n228 B.n141 10.6151
R931 B.n228 B.n227 10.6151
R932 B.n227 B.n226 10.6151
R933 B.n226 B.n143 10.6151
R934 B.n222 B.n143 10.6151
R935 B.n222 B.n221 10.6151
R936 B.n221 B.n220 10.6151
R937 B.n220 B.n145 10.6151
R938 B.n216 B.n145 10.6151
R939 B.n216 B.n215 10.6151
R940 B.n215 B.n214 10.6151
R941 B.n214 B.n147 10.6151
R942 B.n210 B.n147 10.6151
R943 B.n210 B.n209 10.6151
R944 B.n209 B.n208 10.6151
R945 B.n208 B.n149 10.6151
R946 B.n204 B.n149 10.6151
R947 B.n204 B.n203 10.6151
R948 B.n203 B.n202 10.6151
R949 B.n202 B.n151 10.6151
R950 B.n198 B.n151 10.6151
R951 B.n198 B.n197 10.6151
R952 B.n197 B.n196 10.6151
R953 B.n196 B.n153 10.6151
R954 B.n192 B.n153 10.6151
R955 B.n192 B.n191 10.6151
R956 B.n191 B.n190 10.6151
R957 B.n190 B.n155 10.6151
R958 B.n186 B.n155 10.6151
R959 B.n186 B.n185 10.6151
R960 B.n185 B.n184 10.6151
R961 B.n184 B.n157 10.6151
R962 B.n180 B.n157 10.6151
R963 B.n180 B.n179 10.6151
R964 B.n179 B.n178 10.6151
R965 B.n178 B.n159 10.6151
R966 B.n174 B.n159 10.6151
R967 B.n174 B.n173 10.6151
R968 B.n173 B.n172 10.6151
R969 B.n172 B.n161 10.6151
R970 B.n168 B.n161 10.6151
R971 B.n168 B.n167 10.6151
R972 B.n167 B.n166 10.6151
R973 B.n166 B.n163 10.6151
R974 B.n163 B.n0 10.6151
R975 B.n619 B.n1 10.6151
R976 B.n619 B.n618 10.6151
R977 B.n618 B.n617 10.6151
R978 B.n617 B.n4 10.6151
R979 B.n613 B.n4 10.6151
R980 B.n613 B.n612 10.6151
R981 B.n612 B.n611 10.6151
R982 B.n611 B.n6 10.6151
R983 B.n607 B.n6 10.6151
R984 B.n607 B.n606 10.6151
R985 B.n606 B.n605 10.6151
R986 B.n605 B.n8 10.6151
R987 B.n601 B.n8 10.6151
R988 B.n601 B.n600 10.6151
R989 B.n600 B.n599 10.6151
R990 B.n599 B.n10 10.6151
R991 B.n595 B.n10 10.6151
R992 B.n595 B.n594 10.6151
R993 B.n594 B.n593 10.6151
R994 B.n593 B.n12 10.6151
R995 B.n589 B.n12 10.6151
R996 B.n589 B.n588 10.6151
R997 B.n588 B.n587 10.6151
R998 B.n587 B.n14 10.6151
R999 B.n583 B.n14 10.6151
R1000 B.n583 B.n582 10.6151
R1001 B.n582 B.n581 10.6151
R1002 B.n581 B.n16 10.6151
R1003 B.n577 B.n16 10.6151
R1004 B.n577 B.n576 10.6151
R1005 B.n576 B.n575 10.6151
R1006 B.n575 B.n18 10.6151
R1007 B.n571 B.n18 10.6151
R1008 B.n571 B.n570 10.6151
R1009 B.n570 B.n569 10.6151
R1010 B.n569 B.n20 10.6151
R1011 B.n565 B.n20 10.6151
R1012 B.n565 B.n564 10.6151
R1013 B.n564 B.n563 10.6151
R1014 B.n563 B.n22 10.6151
R1015 B.n559 B.n22 10.6151
R1016 B.n559 B.n558 10.6151
R1017 B.n558 B.n557 10.6151
R1018 B.n557 B.n24 10.6151
R1019 B.n553 B.n24 10.6151
R1020 B.n516 B.n515 9.36635
R1021 B.n498 B.n48 9.36635
R1022 B.n269 B.n268 9.36635
R1023 B.n286 B.n121 9.36635
R1024 B.n623 B.n0 2.81026
R1025 B.n623 B.n1 2.81026
R1026 B.n515 B.n514 1.24928
R1027 B.n48 B.n44 1.24928
R1028 B.n270 B.n269 1.24928
R1029 B.n283 B.n121 1.24928
R1030 VP.n13 VP.n10 161.3
R1031 VP.n15 VP.n14 161.3
R1032 VP.n16 VP.n9 161.3
R1033 VP.n18 VP.n17 161.3
R1034 VP.n19 VP.n8 161.3
R1035 VP.n21 VP.n20 161.3
R1036 VP.n43 VP.n42 161.3
R1037 VP.n41 VP.n1 161.3
R1038 VP.n40 VP.n39 161.3
R1039 VP.n38 VP.n2 161.3
R1040 VP.n37 VP.n36 161.3
R1041 VP.n35 VP.n3 161.3
R1042 VP.n33 VP.n32 161.3
R1043 VP.n31 VP.n4 161.3
R1044 VP.n30 VP.n29 161.3
R1045 VP.n28 VP.n5 161.3
R1046 VP.n27 VP.n26 161.3
R1047 VP.n25 VP.n6 161.3
R1048 VP.n11 VP.t1 85.7888
R1049 VP.n24 VP.n23 67.6211
R1050 VP.n44 VP.n0 67.6211
R1051 VP.n22 VP.n7 67.6211
R1052 VP.n12 VP.n11 61.7085
R1053 VP.n29 VP.n28 54.6242
R1054 VP.n40 VP.n2 54.6242
R1055 VP.n18 VP.n9 54.6242
R1056 VP.n23 VP.t3 53.8908
R1057 VP.n34 VP.t2 53.8908
R1058 VP.n0 VP.t4 53.8908
R1059 VP.n7 VP.t0 53.8908
R1060 VP.n12 VP.t5 53.8908
R1061 VP.n24 VP.n22 45.6927
R1062 VP.n28 VP.n27 26.5299
R1063 VP.n41 VP.n40 26.5299
R1064 VP.n19 VP.n18 26.5299
R1065 VP.n27 VP.n6 24.5923
R1066 VP.n29 VP.n4 24.5923
R1067 VP.n33 VP.n4 24.5923
R1068 VP.n36 VP.n35 24.5923
R1069 VP.n36 VP.n2 24.5923
R1070 VP.n42 VP.n41 24.5923
R1071 VP.n20 VP.n19 24.5923
R1072 VP.n14 VP.n13 24.5923
R1073 VP.n14 VP.n9 24.5923
R1074 VP.n23 VP.n6 22.625
R1075 VP.n42 VP.n0 22.625
R1076 VP.n20 VP.n7 22.625
R1077 VP.n34 VP.n33 12.2964
R1078 VP.n35 VP.n34 12.2964
R1079 VP.n13 VP.n12 12.2964
R1080 VP.n11 VP.n10 5.34744
R1081 VP.n22 VP.n21 0.354861
R1082 VP.n25 VP.n24 0.354861
R1083 VP.n44 VP.n43 0.354861
R1084 VP VP.n44 0.267071
R1085 VP.n15 VP.n10 0.189894
R1086 VP.n16 VP.n15 0.189894
R1087 VP.n17 VP.n16 0.189894
R1088 VP.n17 VP.n8 0.189894
R1089 VP.n21 VP.n8 0.189894
R1090 VP.n26 VP.n25 0.189894
R1091 VP.n26 VP.n5 0.189894
R1092 VP.n30 VP.n5 0.189894
R1093 VP.n31 VP.n30 0.189894
R1094 VP.n32 VP.n31 0.189894
R1095 VP.n32 VP.n3 0.189894
R1096 VP.n37 VP.n3 0.189894
R1097 VP.n38 VP.n37 0.189894
R1098 VP.n39 VP.n38 0.189894
R1099 VP.n39 VP.n1 0.189894
R1100 VP.n43 VP.n1 0.189894
R1101 VDD1 VDD1.t4 98.9609
R1102 VDD1.n1 VDD1.t2 98.8472
R1103 VDD1.n1 VDD1.n0 92.4162
R1104 VDD1.n3 VDD1.n2 91.7798
R1105 VDD1.n3 VDD1.n1 40.2272
R1106 VDD1.n2 VDD1.t0 5.04786
R1107 VDD1.n2 VDD1.t5 5.04786
R1108 VDD1.n0 VDD1.t3 5.04786
R1109 VDD1.n0 VDD1.t1 5.04786
R1110 VDD1 VDD1.n3 0.634121
C0 VN w_n3538_n2256# 6.66462f
C1 B VN 1.16194f
C2 VDD2 VN 3.85791f
C3 VP VN 6.16632f
C4 B w_n3538_n2256# 8.51189f
C5 VDD2 w_n3538_n2256# 2.06941f
C6 B VDD2 1.80538f
C7 VTAIL VDD1 5.85136f
C8 VP w_n3538_n2256# 7.12281f
C9 B VP 1.92835f
C10 VP VDD2 0.482021f
C11 VN VDD1 0.151496f
C12 VDD1 w_n3538_n2256# 1.97541f
C13 B VDD1 1.72458f
C14 VDD2 VDD1 1.51586f
C15 VP VDD1 4.18619f
C16 VTAIL VN 4.48846f
C17 VTAIL w_n3538_n2256# 2.22801f
C18 B VTAIL 2.53017f
C19 VTAIL VDD2 5.90551f
C20 VTAIL VP 4.50265f
C21 VDD2 VSUBS 1.695924f
C22 VDD1 VSUBS 2.037599f
C23 VTAIL VSUBS 0.726077f
C24 VN VSUBS 5.8737f
C25 VP VSUBS 2.796976f
C26 B VSUBS 4.443712f
C27 w_n3538_n2256# VSUBS 99.474396f
C28 VDD1.t4 VSUBS 1.04277f
C29 VDD1.t2 VSUBS 1.04195f
C30 VDD1.t3 VSUBS 0.113768f
C31 VDD1.t1 VSUBS 0.113768f
C32 VDD1.n0 VSUBS 0.774635f
C33 VDD1.n1 VSUBS 2.87963f
C34 VDD1.t0 VSUBS 0.113768f
C35 VDD1.t5 VSUBS 0.113768f
C36 VDD1.n2 VSUBS 0.770336f
C37 VDD1.n3 VSUBS 2.36668f
C38 VP.t4 VSUBS 1.82599f
C39 VP.n0 VSUBS 0.822511f
C40 VP.n1 VSUBS 0.037048f
C41 VP.n2 VSUBS 0.064226f
C42 VP.n3 VSUBS 0.037048f
C43 VP.t2 VSUBS 1.82599f
C44 VP.n4 VSUBS 0.068701f
C45 VP.n5 VSUBS 0.037048f
C46 VP.n6 VSUBS 0.065988f
C47 VP.t0 VSUBS 1.82599f
C48 VP.n7 VSUBS 0.822511f
C49 VP.n8 VSUBS 0.037048f
C50 VP.n9 VSUBS 0.064226f
C51 VP.n10 VSUBS 0.393699f
C52 VP.t5 VSUBS 1.82599f
C53 VP.t1 VSUBS 2.16807f
C54 VP.n11 VSUBS 0.760882f
C55 VP.n12 VSUBS 0.790373f
C56 VP.n13 VSUBS 0.051743f
C57 VP.n14 VSUBS 0.068701f
C58 VP.n15 VSUBS 0.037048f
C59 VP.n16 VSUBS 0.037048f
C60 VP.n17 VSUBS 0.037048f
C61 VP.n18 VSUBS 0.041204f
C62 VP.n19 VSUBS 0.07098f
C63 VP.n20 VSUBS 0.065988f
C64 VP.n21 VSUBS 0.059785f
C65 VP.n22 VSUBS 1.82705f
C66 VP.t3 VSUBS 1.82599f
C67 VP.n23 VSUBS 0.822511f
C68 VP.n24 VSUBS 1.85628f
C69 VP.n25 VSUBS 0.059785f
C70 VP.n26 VSUBS 0.037048f
C71 VP.n27 VSUBS 0.07098f
C72 VP.n28 VSUBS 0.041204f
C73 VP.n29 VSUBS 0.064226f
C74 VP.n30 VSUBS 0.037048f
C75 VP.n31 VSUBS 0.037048f
C76 VP.n32 VSUBS 0.037048f
C77 VP.n33 VSUBS 0.051743f
C78 VP.n34 VSUBS 0.675804f
C79 VP.n35 VSUBS 0.051743f
C80 VP.n36 VSUBS 0.068701f
C81 VP.n37 VSUBS 0.037048f
C82 VP.n38 VSUBS 0.037048f
C83 VP.n39 VSUBS 0.037048f
C84 VP.n40 VSUBS 0.041204f
C85 VP.n41 VSUBS 0.07098f
C86 VP.n42 VSUBS 0.065988f
C87 VP.n43 VSUBS 0.059785f
C88 VP.n44 VSUBS 0.071336f
C89 B.n0 VSUBS 0.004677f
C90 B.n1 VSUBS 0.004677f
C91 B.n2 VSUBS 0.007397f
C92 B.n3 VSUBS 0.007397f
C93 B.n4 VSUBS 0.007397f
C94 B.n5 VSUBS 0.007397f
C95 B.n6 VSUBS 0.007397f
C96 B.n7 VSUBS 0.007397f
C97 B.n8 VSUBS 0.007397f
C98 B.n9 VSUBS 0.007397f
C99 B.n10 VSUBS 0.007397f
C100 B.n11 VSUBS 0.007397f
C101 B.n12 VSUBS 0.007397f
C102 B.n13 VSUBS 0.007397f
C103 B.n14 VSUBS 0.007397f
C104 B.n15 VSUBS 0.007397f
C105 B.n16 VSUBS 0.007397f
C106 B.n17 VSUBS 0.007397f
C107 B.n18 VSUBS 0.007397f
C108 B.n19 VSUBS 0.007397f
C109 B.n20 VSUBS 0.007397f
C110 B.n21 VSUBS 0.007397f
C111 B.n22 VSUBS 0.007397f
C112 B.n23 VSUBS 0.007397f
C113 B.n24 VSUBS 0.007397f
C114 B.n25 VSUBS 0.017265f
C115 B.n26 VSUBS 0.007397f
C116 B.n27 VSUBS 0.007397f
C117 B.n28 VSUBS 0.007397f
C118 B.n29 VSUBS 0.007397f
C119 B.n30 VSUBS 0.007397f
C120 B.n31 VSUBS 0.007397f
C121 B.n32 VSUBS 0.007397f
C122 B.n33 VSUBS 0.007397f
C123 B.n34 VSUBS 0.007397f
C124 B.n35 VSUBS 0.007397f
C125 B.n36 VSUBS 0.007397f
C126 B.n37 VSUBS 0.007397f
C127 B.t8 VSUBS 0.201451f
C128 B.t7 VSUBS 0.224375f
C129 B.t6 VSUBS 0.928513f
C130 B.n38 VSUBS 0.132475f
C131 B.n39 VSUBS 0.07645f
C132 B.n40 VSUBS 0.007397f
C133 B.n41 VSUBS 0.007397f
C134 B.n42 VSUBS 0.007397f
C135 B.n43 VSUBS 0.007397f
C136 B.n44 VSUBS 0.004133f
C137 B.n45 VSUBS 0.007397f
C138 B.t2 VSUBS 0.20145f
C139 B.t1 VSUBS 0.224374f
C140 B.t0 VSUBS 0.928513f
C141 B.n46 VSUBS 0.132476f
C142 B.n47 VSUBS 0.076451f
C143 B.n48 VSUBS 0.017137f
C144 B.n49 VSUBS 0.007397f
C145 B.n50 VSUBS 0.007397f
C146 B.n51 VSUBS 0.007397f
C147 B.n52 VSUBS 0.007397f
C148 B.n53 VSUBS 0.007397f
C149 B.n54 VSUBS 0.007397f
C150 B.n55 VSUBS 0.007397f
C151 B.n56 VSUBS 0.007397f
C152 B.n57 VSUBS 0.007397f
C153 B.n58 VSUBS 0.007397f
C154 B.n59 VSUBS 0.007397f
C155 B.n60 VSUBS 0.016672f
C156 B.n61 VSUBS 0.007397f
C157 B.n62 VSUBS 0.007397f
C158 B.n63 VSUBS 0.007397f
C159 B.n64 VSUBS 0.007397f
C160 B.n65 VSUBS 0.007397f
C161 B.n66 VSUBS 0.007397f
C162 B.n67 VSUBS 0.007397f
C163 B.n68 VSUBS 0.007397f
C164 B.n69 VSUBS 0.007397f
C165 B.n70 VSUBS 0.007397f
C166 B.n71 VSUBS 0.007397f
C167 B.n72 VSUBS 0.007397f
C168 B.n73 VSUBS 0.007397f
C169 B.n74 VSUBS 0.007397f
C170 B.n75 VSUBS 0.007397f
C171 B.n76 VSUBS 0.007397f
C172 B.n77 VSUBS 0.007397f
C173 B.n78 VSUBS 0.007397f
C174 B.n79 VSUBS 0.007397f
C175 B.n80 VSUBS 0.007397f
C176 B.n81 VSUBS 0.007397f
C177 B.n82 VSUBS 0.007397f
C178 B.n83 VSUBS 0.007397f
C179 B.n84 VSUBS 0.007397f
C180 B.n85 VSUBS 0.007397f
C181 B.n86 VSUBS 0.007397f
C182 B.n87 VSUBS 0.007397f
C183 B.n88 VSUBS 0.007397f
C184 B.n89 VSUBS 0.007397f
C185 B.n90 VSUBS 0.007397f
C186 B.n91 VSUBS 0.007397f
C187 B.n92 VSUBS 0.007397f
C188 B.n93 VSUBS 0.007397f
C189 B.n94 VSUBS 0.007397f
C190 B.n95 VSUBS 0.007397f
C191 B.n96 VSUBS 0.007397f
C192 B.n97 VSUBS 0.007397f
C193 B.n98 VSUBS 0.007397f
C194 B.n99 VSUBS 0.007397f
C195 B.n100 VSUBS 0.007397f
C196 B.n101 VSUBS 0.007397f
C197 B.n102 VSUBS 0.007397f
C198 B.n103 VSUBS 0.007397f
C199 B.n104 VSUBS 0.007397f
C200 B.n105 VSUBS 0.007397f
C201 B.n106 VSUBS 0.016672f
C202 B.n107 VSUBS 0.007397f
C203 B.n108 VSUBS 0.007397f
C204 B.n109 VSUBS 0.007397f
C205 B.n110 VSUBS 0.007397f
C206 B.n111 VSUBS 0.007397f
C207 B.n112 VSUBS 0.007397f
C208 B.n113 VSUBS 0.007397f
C209 B.n114 VSUBS 0.007397f
C210 B.n115 VSUBS 0.007397f
C211 B.n116 VSUBS 0.007397f
C212 B.n117 VSUBS 0.007397f
C213 B.n118 VSUBS 0.007397f
C214 B.t10 VSUBS 0.20145f
C215 B.t11 VSUBS 0.224374f
C216 B.t9 VSUBS 0.928513f
C217 B.n119 VSUBS 0.132476f
C218 B.n120 VSUBS 0.076451f
C219 B.n121 VSUBS 0.017137f
C220 B.n122 VSUBS 0.007397f
C221 B.n123 VSUBS 0.007397f
C222 B.n124 VSUBS 0.007397f
C223 B.n125 VSUBS 0.007397f
C224 B.n126 VSUBS 0.007397f
C225 B.t4 VSUBS 0.201451f
C226 B.t5 VSUBS 0.224375f
C227 B.t3 VSUBS 0.928513f
C228 B.n127 VSUBS 0.132475f
C229 B.n128 VSUBS 0.07645f
C230 B.n129 VSUBS 0.007397f
C231 B.n130 VSUBS 0.007397f
C232 B.n131 VSUBS 0.007397f
C233 B.n132 VSUBS 0.007397f
C234 B.n133 VSUBS 0.007397f
C235 B.n134 VSUBS 0.007397f
C236 B.n135 VSUBS 0.007397f
C237 B.n136 VSUBS 0.007397f
C238 B.n137 VSUBS 0.007397f
C239 B.n138 VSUBS 0.007397f
C240 B.n139 VSUBS 0.007397f
C241 B.n140 VSUBS 0.007397f
C242 B.n141 VSUBS 0.016672f
C243 B.n142 VSUBS 0.007397f
C244 B.n143 VSUBS 0.007397f
C245 B.n144 VSUBS 0.007397f
C246 B.n145 VSUBS 0.007397f
C247 B.n146 VSUBS 0.007397f
C248 B.n147 VSUBS 0.007397f
C249 B.n148 VSUBS 0.007397f
C250 B.n149 VSUBS 0.007397f
C251 B.n150 VSUBS 0.007397f
C252 B.n151 VSUBS 0.007397f
C253 B.n152 VSUBS 0.007397f
C254 B.n153 VSUBS 0.007397f
C255 B.n154 VSUBS 0.007397f
C256 B.n155 VSUBS 0.007397f
C257 B.n156 VSUBS 0.007397f
C258 B.n157 VSUBS 0.007397f
C259 B.n158 VSUBS 0.007397f
C260 B.n159 VSUBS 0.007397f
C261 B.n160 VSUBS 0.007397f
C262 B.n161 VSUBS 0.007397f
C263 B.n162 VSUBS 0.007397f
C264 B.n163 VSUBS 0.007397f
C265 B.n164 VSUBS 0.007397f
C266 B.n165 VSUBS 0.007397f
C267 B.n166 VSUBS 0.007397f
C268 B.n167 VSUBS 0.007397f
C269 B.n168 VSUBS 0.007397f
C270 B.n169 VSUBS 0.007397f
C271 B.n170 VSUBS 0.007397f
C272 B.n171 VSUBS 0.007397f
C273 B.n172 VSUBS 0.007397f
C274 B.n173 VSUBS 0.007397f
C275 B.n174 VSUBS 0.007397f
C276 B.n175 VSUBS 0.007397f
C277 B.n176 VSUBS 0.007397f
C278 B.n177 VSUBS 0.007397f
C279 B.n178 VSUBS 0.007397f
C280 B.n179 VSUBS 0.007397f
C281 B.n180 VSUBS 0.007397f
C282 B.n181 VSUBS 0.007397f
C283 B.n182 VSUBS 0.007397f
C284 B.n183 VSUBS 0.007397f
C285 B.n184 VSUBS 0.007397f
C286 B.n185 VSUBS 0.007397f
C287 B.n186 VSUBS 0.007397f
C288 B.n187 VSUBS 0.007397f
C289 B.n188 VSUBS 0.007397f
C290 B.n189 VSUBS 0.007397f
C291 B.n190 VSUBS 0.007397f
C292 B.n191 VSUBS 0.007397f
C293 B.n192 VSUBS 0.007397f
C294 B.n193 VSUBS 0.007397f
C295 B.n194 VSUBS 0.007397f
C296 B.n195 VSUBS 0.007397f
C297 B.n196 VSUBS 0.007397f
C298 B.n197 VSUBS 0.007397f
C299 B.n198 VSUBS 0.007397f
C300 B.n199 VSUBS 0.007397f
C301 B.n200 VSUBS 0.007397f
C302 B.n201 VSUBS 0.007397f
C303 B.n202 VSUBS 0.007397f
C304 B.n203 VSUBS 0.007397f
C305 B.n204 VSUBS 0.007397f
C306 B.n205 VSUBS 0.007397f
C307 B.n206 VSUBS 0.007397f
C308 B.n207 VSUBS 0.007397f
C309 B.n208 VSUBS 0.007397f
C310 B.n209 VSUBS 0.007397f
C311 B.n210 VSUBS 0.007397f
C312 B.n211 VSUBS 0.007397f
C313 B.n212 VSUBS 0.007397f
C314 B.n213 VSUBS 0.007397f
C315 B.n214 VSUBS 0.007397f
C316 B.n215 VSUBS 0.007397f
C317 B.n216 VSUBS 0.007397f
C318 B.n217 VSUBS 0.007397f
C319 B.n218 VSUBS 0.007397f
C320 B.n219 VSUBS 0.007397f
C321 B.n220 VSUBS 0.007397f
C322 B.n221 VSUBS 0.007397f
C323 B.n222 VSUBS 0.007397f
C324 B.n223 VSUBS 0.007397f
C325 B.n224 VSUBS 0.007397f
C326 B.n225 VSUBS 0.007397f
C327 B.n226 VSUBS 0.007397f
C328 B.n227 VSUBS 0.007397f
C329 B.n228 VSUBS 0.007397f
C330 B.n229 VSUBS 0.007397f
C331 B.n230 VSUBS 0.016672f
C332 B.n231 VSUBS 0.017265f
C333 B.n232 VSUBS 0.017265f
C334 B.n233 VSUBS 0.007397f
C335 B.n234 VSUBS 0.007397f
C336 B.n235 VSUBS 0.007397f
C337 B.n236 VSUBS 0.007397f
C338 B.n237 VSUBS 0.007397f
C339 B.n238 VSUBS 0.007397f
C340 B.n239 VSUBS 0.007397f
C341 B.n240 VSUBS 0.007397f
C342 B.n241 VSUBS 0.007397f
C343 B.n242 VSUBS 0.007397f
C344 B.n243 VSUBS 0.007397f
C345 B.n244 VSUBS 0.007397f
C346 B.n245 VSUBS 0.007397f
C347 B.n246 VSUBS 0.007397f
C348 B.n247 VSUBS 0.007397f
C349 B.n248 VSUBS 0.007397f
C350 B.n249 VSUBS 0.007397f
C351 B.n250 VSUBS 0.007397f
C352 B.n251 VSUBS 0.007397f
C353 B.n252 VSUBS 0.007397f
C354 B.n253 VSUBS 0.007397f
C355 B.n254 VSUBS 0.007397f
C356 B.n255 VSUBS 0.007397f
C357 B.n256 VSUBS 0.007397f
C358 B.n257 VSUBS 0.007397f
C359 B.n258 VSUBS 0.007397f
C360 B.n259 VSUBS 0.007397f
C361 B.n260 VSUBS 0.007397f
C362 B.n261 VSUBS 0.007397f
C363 B.n262 VSUBS 0.007397f
C364 B.n263 VSUBS 0.007397f
C365 B.n264 VSUBS 0.007397f
C366 B.n265 VSUBS 0.007397f
C367 B.n266 VSUBS 0.007397f
C368 B.n267 VSUBS 0.007397f
C369 B.n268 VSUBS 0.006962f
C370 B.n269 VSUBS 0.017137f
C371 B.n270 VSUBS 0.004133f
C372 B.n271 VSUBS 0.007397f
C373 B.n272 VSUBS 0.007397f
C374 B.n273 VSUBS 0.007397f
C375 B.n274 VSUBS 0.007397f
C376 B.n275 VSUBS 0.007397f
C377 B.n276 VSUBS 0.007397f
C378 B.n277 VSUBS 0.007397f
C379 B.n278 VSUBS 0.007397f
C380 B.n279 VSUBS 0.007397f
C381 B.n280 VSUBS 0.007397f
C382 B.n281 VSUBS 0.007397f
C383 B.n282 VSUBS 0.007397f
C384 B.n283 VSUBS 0.004133f
C385 B.n284 VSUBS 0.007397f
C386 B.n285 VSUBS 0.007397f
C387 B.n286 VSUBS 0.006962f
C388 B.n287 VSUBS 0.007397f
C389 B.n288 VSUBS 0.007397f
C390 B.n289 VSUBS 0.007397f
C391 B.n290 VSUBS 0.007397f
C392 B.n291 VSUBS 0.007397f
C393 B.n292 VSUBS 0.007397f
C394 B.n293 VSUBS 0.007397f
C395 B.n294 VSUBS 0.007397f
C396 B.n295 VSUBS 0.007397f
C397 B.n296 VSUBS 0.007397f
C398 B.n297 VSUBS 0.007397f
C399 B.n298 VSUBS 0.007397f
C400 B.n299 VSUBS 0.007397f
C401 B.n300 VSUBS 0.007397f
C402 B.n301 VSUBS 0.007397f
C403 B.n302 VSUBS 0.007397f
C404 B.n303 VSUBS 0.007397f
C405 B.n304 VSUBS 0.007397f
C406 B.n305 VSUBS 0.007397f
C407 B.n306 VSUBS 0.007397f
C408 B.n307 VSUBS 0.007397f
C409 B.n308 VSUBS 0.007397f
C410 B.n309 VSUBS 0.007397f
C411 B.n310 VSUBS 0.007397f
C412 B.n311 VSUBS 0.007397f
C413 B.n312 VSUBS 0.007397f
C414 B.n313 VSUBS 0.007397f
C415 B.n314 VSUBS 0.007397f
C416 B.n315 VSUBS 0.007397f
C417 B.n316 VSUBS 0.007397f
C418 B.n317 VSUBS 0.007397f
C419 B.n318 VSUBS 0.007397f
C420 B.n319 VSUBS 0.007397f
C421 B.n320 VSUBS 0.007397f
C422 B.n321 VSUBS 0.017265f
C423 B.n322 VSUBS 0.017265f
C424 B.n323 VSUBS 0.016672f
C425 B.n324 VSUBS 0.007397f
C426 B.n325 VSUBS 0.007397f
C427 B.n326 VSUBS 0.007397f
C428 B.n327 VSUBS 0.007397f
C429 B.n328 VSUBS 0.007397f
C430 B.n329 VSUBS 0.007397f
C431 B.n330 VSUBS 0.007397f
C432 B.n331 VSUBS 0.007397f
C433 B.n332 VSUBS 0.007397f
C434 B.n333 VSUBS 0.007397f
C435 B.n334 VSUBS 0.007397f
C436 B.n335 VSUBS 0.007397f
C437 B.n336 VSUBS 0.007397f
C438 B.n337 VSUBS 0.007397f
C439 B.n338 VSUBS 0.007397f
C440 B.n339 VSUBS 0.007397f
C441 B.n340 VSUBS 0.007397f
C442 B.n341 VSUBS 0.007397f
C443 B.n342 VSUBS 0.007397f
C444 B.n343 VSUBS 0.007397f
C445 B.n344 VSUBS 0.007397f
C446 B.n345 VSUBS 0.007397f
C447 B.n346 VSUBS 0.007397f
C448 B.n347 VSUBS 0.007397f
C449 B.n348 VSUBS 0.007397f
C450 B.n349 VSUBS 0.007397f
C451 B.n350 VSUBS 0.007397f
C452 B.n351 VSUBS 0.007397f
C453 B.n352 VSUBS 0.007397f
C454 B.n353 VSUBS 0.007397f
C455 B.n354 VSUBS 0.007397f
C456 B.n355 VSUBS 0.007397f
C457 B.n356 VSUBS 0.007397f
C458 B.n357 VSUBS 0.007397f
C459 B.n358 VSUBS 0.007397f
C460 B.n359 VSUBS 0.007397f
C461 B.n360 VSUBS 0.007397f
C462 B.n361 VSUBS 0.007397f
C463 B.n362 VSUBS 0.007397f
C464 B.n363 VSUBS 0.007397f
C465 B.n364 VSUBS 0.007397f
C466 B.n365 VSUBS 0.007397f
C467 B.n366 VSUBS 0.007397f
C468 B.n367 VSUBS 0.007397f
C469 B.n368 VSUBS 0.007397f
C470 B.n369 VSUBS 0.007397f
C471 B.n370 VSUBS 0.007397f
C472 B.n371 VSUBS 0.007397f
C473 B.n372 VSUBS 0.007397f
C474 B.n373 VSUBS 0.007397f
C475 B.n374 VSUBS 0.007397f
C476 B.n375 VSUBS 0.007397f
C477 B.n376 VSUBS 0.007397f
C478 B.n377 VSUBS 0.007397f
C479 B.n378 VSUBS 0.007397f
C480 B.n379 VSUBS 0.007397f
C481 B.n380 VSUBS 0.007397f
C482 B.n381 VSUBS 0.007397f
C483 B.n382 VSUBS 0.007397f
C484 B.n383 VSUBS 0.007397f
C485 B.n384 VSUBS 0.007397f
C486 B.n385 VSUBS 0.007397f
C487 B.n386 VSUBS 0.007397f
C488 B.n387 VSUBS 0.007397f
C489 B.n388 VSUBS 0.007397f
C490 B.n389 VSUBS 0.007397f
C491 B.n390 VSUBS 0.007397f
C492 B.n391 VSUBS 0.007397f
C493 B.n392 VSUBS 0.007397f
C494 B.n393 VSUBS 0.007397f
C495 B.n394 VSUBS 0.007397f
C496 B.n395 VSUBS 0.007397f
C497 B.n396 VSUBS 0.007397f
C498 B.n397 VSUBS 0.007397f
C499 B.n398 VSUBS 0.007397f
C500 B.n399 VSUBS 0.007397f
C501 B.n400 VSUBS 0.007397f
C502 B.n401 VSUBS 0.007397f
C503 B.n402 VSUBS 0.007397f
C504 B.n403 VSUBS 0.007397f
C505 B.n404 VSUBS 0.007397f
C506 B.n405 VSUBS 0.007397f
C507 B.n406 VSUBS 0.007397f
C508 B.n407 VSUBS 0.007397f
C509 B.n408 VSUBS 0.007397f
C510 B.n409 VSUBS 0.007397f
C511 B.n410 VSUBS 0.007397f
C512 B.n411 VSUBS 0.007397f
C513 B.n412 VSUBS 0.007397f
C514 B.n413 VSUBS 0.007397f
C515 B.n414 VSUBS 0.007397f
C516 B.n415 VSUBS 0.007397f
C517 B.n416 VSUBS 0.007397f
C518 B.n417 VSUBS 0.007397f
C519 B.n418 VSUBS 0.007397f
C520 B.n419 VSUBS 0.007397f
C521 B.n420 VSUBS 0.007397f
C522 B.n421 VSUBS 0.007397f
C523 B.n422 VSUBS 0.007397f
C524 B.n423 VSUBS 0.007397f
C525 B.n424 VSUBS 0.007397f
C526 B.n425 VSUBS 0.007397f
C527 B.n426 VSUBS 0.007397f
C528 B.n427 VSUBS 0.007397f
C529 B.n428 VSUBS 0.007397f
C530 B.n429 VSUBS 0.007397f
C531 B.n430 VSUBS 0.007397f
C532 B.n431 VSUBS 0.007397f
C533 B.n432 VSUBS 0.007397f
C534 B.n433 VSUBS 0.007397f
C535 B.n434 VSUBS 0.007397f
C536 B.n435 VSUBS 0.007397f
C537 B.n436 VSUBS 0.007397f
C538 B.n437 VSUBS 0.007397f
C539 B.n438 VSUBS 0.007397f
C540 B.n439 VSUBS 0.007397f
C541 B.n440 VSUBS 0.007397f
C542 B.n441 VSUBS 0.007397f
C543 B.n442 VSUBS 0.007397f
C544 B.n443 VSUBS 0.007397f
C545 B.n444 VSUBS 0.007397f
C546 B.n445 VSUBS 0.007397f
C547 B.n446 VSUBS 0.007397f
C548 B.n447 VSUBS 0.007397f
C549 B.n448 VSUBS 0.007397f
C550 B.n449 VSUBS 0.007397f
C551 B.n450 VSUBS 0.007397f
C552 B.n451 VSUBS 0.007397f
C553 B.n452 VSUBS 0.007397f
C554 B.n453 VSUBS 0.007397f
C555 B.n454 VSUBS 0.007397f
C556 B.n455 VSUBS 0.007397f
C557 B.n456 VSUBS 0.007397f
C558 B.n457 VSUBS 0.007397f
C559 B.n458 VSUBS 0.007397f
C560 B.n459 VSUBS 0.007397f
C561 B.n460 VSUBS 0.007397f
C562 B.n461 VSUBS 0.017573f
C563 B.n462 VSUBS 0.016365f
C564 B.n463 VSUBS 0.017265f
C565 B.n464 VSUBS 0.007397f
C566 B.n465 VSUBS 0.007397f
C567 B.n466 VSUBS 0.007397f
C568 B.n467 VSUBS 0.007397f
C569 B.n468 VSUBS 0.007397f
C570 B.n469 VSUBS 0.007397f
C571 B.n470 VSUBS 0.007397f
C572 B.n471 VSUBS 0.007397f
C573 B.n472 VSUBS 0.007397f
C574 B.n473 VSUBS 0.007397f
C575 B.n474 VSUBS 0.007397f
C576 B.n475 VSUBS 0.007397f
C577 B.n476 VSUBS 0.007397f
C578 B.n477 VSUBS 0.007397f
C579 B.n478 VSUBS 0.007397f
C580 B.n479 VSUBS 0.007397f
C581 B.n480 VSUBS 0.007397f
C582 B.n481 VSUBS 0.007397f
C583 B.n482 VSUBS 0.007397f
C584 B.n483 VSUBS 0.007397f
C585 B.n484 VSUBS 0.007397f
C586 B.n485 VSUBS 0.007397f
C587 B.n486 VSUBS 0.007397f
C588 B.n487 VSUBS 0.007397f
C589 B.n488 VSUBS 0.007397f
C590 B.n489 VSUBS 0.007397f
C591 B.n490 VSUBS 0.007397f
C592 B.n491 VSUBS 0.007397f
C593 B.n492 VSUBS 0.007397f
C594 B.n493 VSUBS 0.007397f
C595 B.n494 VSUBS 0.007397f
C596 B.n495 VSUBS 0.007397f
C597 B.n496 VSUBS 0.007397f
C598 B.n497 VSUBS 0.007397f
C599 B.n498 VSUBS 0.006962f
C600 B.n499 VSUBS 0.007397f
C601 B.n500 VSUBS 0.007397f
C602 B.n501 VSUBS 0.007397f
C603 B.n502 VSUBS 0.007397f
C604 B.n503 VSUBS 0.007397f
C605 B.n504 VSUBS 0.007397f
C606 B.n505 VSUBS 0.007397f
C607 B.n506 VSUBS 0.007397f
C608 B.n507 VSUBS 0.007397f
C609 B.n508 VSUBS 0.007397f
C610 B.n509 VSUBS 0.007397f
C611 B.n510 VSUBS 0.007397f
C612 B.n511 VSUBS 0.007397f
C613 B.n512 VSUBS 0.007397f
C614 B.n513 VSUBS 0.007397f
C615 B.n514 VSUBS 0.004133f
C616 B.n515 VSUBS 0.017137f
C617 B.n516 VSUBS 0.006962f
C618 B.n517 VSUBS 0.007397f
C619 B.n518 VSUBS 0.007397f
C620 B.n519 VSUBS 0.007397f
C621 B.n520 VSUBS 0.007397f
C622 B.n521 VSUBS 0.007397f
C623 B.n522 VSUBS 0.007397f
C624 B.n523 VSUBS 0.007397f
C625 B.n524 VSUBS 0.007397f
C626 B.n525 VSUBS 0.007397f
C627 B.n526 VSUBS 0.007397f
C628 B.n527 VSUBS 0.007397f
C629 B.n528 VSUBS 0.007397f
C630 B.n529 VSUBS 0.007397f
C631 B.n530 VSUBS 0.007397f
C632 B.n531 VSUBS 0.007397f
C633 B.n532 VSUBS 0.007397f
C634 B.n533 VSUBS 0.007397f
C635 B.n534 VSUBS 0.007397f
C636 B.n535 VSUBS 0.007397f
C637 B.n536 VSUBS 0.007397f
C638 B.n537 VSUBS 0.007397f
C639 B.n538 VSUBS 0.007397f
C640 B.n539 VSUBS 0.007397f
C641 B.n540 VSUBS 0.007397f
C642 B.n541 VSUBS 0.007397f
C643 B.n542 VSUBS 0.007397f
C644 B.n543 VSUBS 0.007397f
C645 B.n544 VSUBS 0.007397f
C646 B.n545 VSUBS 0.007397f
C647 B.n546 VSUBS 0.007397f
C648 B.n547 VSUBS 0.007397f
C649 B.n548 VSUBS 0.007397f
C650 B.n549 VSUBS 0.007397f
C651 B.n550 VSUBS 0.007397f
C652 B.n551 VSUBS 0.007397f
C653 B.n552 VSUBS 0.017265f
C654 B.n553 VSUBS 0.016672f
C655 B.n554 VSUBS 0.016672f
C656 B.n555 VSUBS 0.007397f
C657 B.n556 VSUBS 0.007397f
C658 B.n557 VSUBS 0.007397f
C659 B.n558 VSUBS 0.007397f
C660 B.n559 VSUBS 0.007397f
C661 B.n560 VSUBS 0.007397f
C662 B.n561 VSUBS 0.007397f
C663 B.n562 VSUBS 0.007397f
C664 B.n563 VSUBS 0.007397f
C665 B.n564 VSUBS 0.007397f
C666 B.n565 VSUBS 0.007397f
C667 B.n566 VSUBS 0.007397f
C668 B.n567 VSUBS 0.007397f
C669 B.n568 VSUBS 0.007397f
C670 B.n569 VSUBS 0.007397f
C671 B.n570 VSUBS 0.007397f
C672 B.n571 VSUBS 0.007397f
C673 B.n572 VSUBS 0.007397f
C674 B.n573 VSUBS 0.007397f
C675 B.n574 VSUBS 0.007397f
C676 B.n575 VSUBS 0.007397f
C677 B.n576 VSUBS 0.007397f
C678 B.n577 VSUBS 0.007397f
C679 B.n578 VSUBS 0.007397f
C680 B.n579 VSUBS 0.007397f
C681 B.n580 VSUBS 0.007397f
C682 B.n581 VSUBS 0.007397f
C683 B.n582 VSUBS 0.007397f
C684 B.n583 VSUBS 0.007397f
C685 B.n584 VSUBS 0.007397f
C686 B.n585 VSUBS 0.007397f
C687 B.n586 VSUBS 0.007397f
C688 B.n587 VSUBS 0.007397f
C689 B.n588 VSUBS 0.007397f
C690 B.n589 VSUBS 0.007397f
C691 B.n590 VSUBS 0.007397f
C692 B.n591 VSUBS 0.007397f
C693 B.n592 VSUBS 0.007397f
C694 B.n593 VSUBS 0.007397f
C695 B.n594 VSUBS 0.007397f
C696 B.n595 VSUBS 0.007397f
C697 B.n596 VSUBS 0.007397f
C698 B.n597 VSUBS 0.007397f
C699 B.n598 VSUBS 0.007397f
C700 B.n599 VSUBS 0.007397f
C701 B.n600 VSUBS 0.007397f
C702 B.n601 VSUBS 0.007397f
C703 B.n602 VSUBS 0.007397f
C704 B.n603 VSUBS 0.007397f
C705 B.n604 VSUBS 0.007397f
C706 B.n605 VSUBS 0.007397f
C707 B.n606 VSUBS 0.007397f
C708 B.n607 VSUBS 0.007397f
C709 B.n608 VSUBS 0.007397f
C710 B.n609 VSUBS 0.007397f
C711 B.n610 VSUBS 0.007397f
C712 B.n611 VSUBS 0.007397f
C713 B.n612 VSUBS 0.007397f
C714 B.n613 VSUBS 0.007397f
C715 B.n614 VSUBS 0.007397f
C716 B.n615 VSUBS 0.007397f
C717 B.n616 VSUBS 0.007397f
C718 B.n617 VSUBS 0.007397f
C719 B.n618 VSUBS 0.007397f
C720 B.n619 VSUBS 0.007397f
C721 B.n620 VSUBS 0.007397f
C722 B.n621 VSUBS 0.007397f
C723 B.n622 VSUBS 0.007397f
C724 B.n623 VSUBS 0.016749f
C725 VDD2.t3 VSUBS 1.23776f
C726 VDD2.t4 VSUBS 0.135148f
C727 VDD2.t5 VSUBS 0.135148f
C728 VDD2.n0 VSUBS 0.920211f
C729 VDD2.n1 VSUBS 3.28685f
C730 VDD2.t1 VSUBS 1.22382f
C731 VDD2.n2 VSUBS 2.79873f
C732 VDD2.t0 VSUBS 0.135148f
C733 VDD2.t2 VSUBS 0.135148f
C734 VDD2.n3 VSUBS 0.920179f
C735 VTAIL.t6 VSUBS 0.169037f
C736 VTAIL.t10 VSUBS 0.169037f
C737 VTAIL.n0 VSUBS 1.02419f
C738 VTAIL.n1 VSUBS 0.90223f
C739 VTAIL.t0 VSUBS 1.40231f
C740 VTAIL.n2 VSUBS 1.20102f
C741 VTAIL.t5 VSUBS 0.169037f
C742 VTAIL.t4 VSUBS 0.169037f
C743 VTAIL.n3 VSUBS 1.02419f
C744 VTAIL.n4 VSUBS 2.55749f
C745 VTAIL.t9 VSUBS 0.169037f
C746 VTAIL.t7 VSUBS 0.169037f
C747 VTAIL.n5 VSUBS 1.0242f
C748 VTAIL.n6 VSUBS 2.55748f
C749 VTAIL.t11 VSUBS 1.40232f
C750 VTAIL.n7 VSUBS 1.20101f
C751 VTAIL.t3 VSUBS 0.169037f
C752 VTAIL.t1 VSUBS 0.169037f
C753 VTAIL.n8 VSUBS 1.0242f
C754 VTAIL.n9 VSUBS 1.11812f
C755 VTAIL.t2 VSUBS 1.40231f
C756 VTAIL.n10 VSUBS 2.3442f
C757 VTAIL.t8 VSUBS 1.40231f
C758 VTAIL.n11 VSUBS 2.26393f
C759 VN.t0 VSUBS 1.76372f
C760 VN.n0 VSUBS 0.79446f
C761 VN.n1 VSUBS 0.035784f
C762 VN.n2 VSUBS 0.062036f
C763 VN.n3 VSUBS 0.380272f
C764 VN.t1 VSUBS 1.76372f
C765 VN.t2 VSUBS 2.09413f
C766 VN.n4 VSUBS 0.734931f
C767 VN.n5 VSUBS 0.763418f
C768 VN.n6 VSUBS 0.049979f
C769 VN.n7 VSUBS 0.066358f
C770 VN.n8 VSUBS 0.035784f
C771 VN.n9 VSUBS 0.035784f
C772 VN.n10 VSUBS 0.035784f
C773 VN.n11 VSUBS 0.039799f
C774 VN.n12 VSUBS 0.06856f
C775 VN.n13 VSUBS 0.063738f
C776 VN.n14 VSUBS 0.057746f
C777 VN.n15 VSUBS 0.068904f
C778 VN.t4 VSUBS 1.76372f
C779 VN.n16 VSUBS 0.79446f
C780 VN.n17 VSUBS 0.035784f
C781 VN.n18 VSUBS 0.062036f
C782 VN.n19 VSUBS 0.380272f
C783 VN.t5 VSUBS 1.76372f
C784 VN.t3 VSUBS 2.09413f
C785 VN.n20 VSUBS 0.734931f
C786 VN.n21 VSUBS 0.763418f
C787 VN.n22 VSUBS 0.049979f
C788 VN.n23 VSUBS 0.066358f
C789 VN.n24 VSUBS 0.035784f
C790 VN.n25 VSUBS 0.035784f
C791 VN.n26 VSUBS 0.035784f
C792 VN.n27 VSUBS 0.039799f
C793 VN.n28 VSUBS 0.06856f
C794 VN.n29 VSUBS 0.063738f
C795 VN.n30 VSUBS 0.057746f
C796 VN.n31 VSUBS 1.77986f
.ends

