* NGSPICE file created from diff_pair_sample_0542.ext - technology: sky130A

.subckt diff_pair_sample_0542 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=1.419 ps=8.93 w=8.6 l=3.66
X1 VTAIL.t14 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X2 VDD2.t7 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=3.354 ps=17.98 w=8.6 l=3.66
X3 VDD1.t6 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=3.354 ps=17.98 w=8.6 l=3.66
X4 VDD1.t7 VP.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X5 VDD1.t3 VP.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=3.354 ps=17.98 w=8.6 l=3.66
X6 VTAIL.t10 VP.t5 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X7 VDD2.t6 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X8 VTAIL.t3 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=1.419 ps=8.93 w=8.6 l=3.66
X9 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X10 VDD2.t3 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X11 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=0 ps=0 w=8.6 l=3.66
X12 VTAIL.t6 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=1.419 ps=8.93 w=8.6 l=3.66
X13 VDD2.t1 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=3.354 ps=17.98 w=8.6 l=3.66
X14 VTAIL.t9 VP.t6 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=1.419 ps=8.93 w=8.6 l=3.66
X15 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=0 ps=0 w=8.6 l=3.66
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=0 ps=0 w=8.6 l=3.66
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.354 pd=17.98 as=0 ps=0 w=8.6 l=3.66
X18 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
X19 VDD1.t4 VP.t7 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.419 pd=8.93 as=1.419 ps=8.93 w=8.6 l=3.66
R0 VP.n22 VP.n19 161.3
R1 VP.n24 VP.n23 161.3
R2 VP.n25 VP.n18 161.3
R3 VP.n27 VP.n26 161.3
R4 VP.n28 VP.n17 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n31 VP.n16 161.3
R7 VP.n34 VP.n33 161.3
R8 VP.n35 VP.n15 161.3
R9 VP.n37 VP.n36 161.3
R10 VP.n38 VP.n14 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n41 VP.n13 161.3
R13 VP.n43 VP.n42 161.3
R14 VP.n44 VP.n12 161.3
R15 VP.n84 VP.n0 161.3
R16 VP.n83 VP.n82 161.3
R17 VP.n81 VP.n1 161.3
R18 VP.n80 VP.n79 161.3
R19 VP.n78 VP.n2 161.3
R20 VP.n77 VP.n76 161.3
R21 VP.n75 VP.n3 161.3
R22 VP.n74 VP.n73 161.3
R23 VP.n71 VP.n4 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n68 VP.n5 161.3
R26 VP.n67 VP.n66 161.3
R27 VP.n65 VP.n6 161.3
R28 VP.n64 VP.n63 161.3
R29 VP.n62 VP.n7 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n58 VP.n8 161.3
R32 VP.n57 VP.n56 161.3
R33 VP.n55 VP.n9 161.3
R34 VP.n54 VP.n53 161.3
R35 VP.n52 VP.n10 161.3
R36 VP.n51 VP.n50 161.3
R37 VP.n49 VP.n11 161.3
R38 VP.n21 VP.t0 88.8824
R39 VP.n48 VP.n47 58.5258
R40 VP.n86 VP.n85 58.5258
R41 VP.n46 VP.n45 58.5258
R42 VP.n47 VP.t6 56.6289
R43 VP.n59 VP.t7 56.6289
R44 VP.n72 VP.t1 56.6289
R45 VP.n85 VP.t2 56.6289
R46 VP.n45 VP.t4 56.6289
R47 VP.n32 VP.t5 56.6289
R48 VP.n20 VP.t3 56.6289
R49 VP.n48 VP.n46 53.4969
R50 VP.n21 VP.n20 50.8254
R51 VP.n53 VP.n9 41.5458
R52 VP.n79 VP.n78 41.5458
R53 VP.n39 VP.n38 41.5458
R54 VP.n66 VP.n65 40.577
R55 VP.n66 VP.n5 40.577
R56 VP.n26 VP.n17 40.577
R57 VP.n26 VP.n25 40.577
R58 VP.n53 VP.n52 39.6083
R59 VP.n79 VP.n1 39.6083
R60 VP.n39 VP.n13 39.6083
R61 VP.n51 VP.n11 24.5923
R62 VP.n52 VP.n51 24.5923
R63 VP.n57 VP.n9 24.5923
R64 VP.n58 VP.n57 24.5923
R65 VP.n60 VP.n58 24.5923
R66 VP.n64 VP.n7 24.5923
R67 VP.n65 VP.n64 24.5923
R68 VP.n70 VP.n5 24.5923
R69 VP.n71 VP.n70 24.5923
R70 VP.n73 VP.n3 24.5923
R71 VP.n77 VP.n3 24.5923
R72 VP.n78 VP.n77 24.5923
R73 VP.n83 VP.n1 24.5923
R74 VP.n84 VP.n83 24.5923
R75 VP.n43 VP.n13 24.5923
R76 VP.n44 VP.n43 24.5923
R77 VP.n30 VP.n17 24.5923
R78 VP.n31 VP.n30 24.5923
R79 VP.n33 VP.n15 24.5923
R80 VP.n37 VP.n15 24.5923
R81 VP.n38 VP.n37 24.5923
R82 VP.n24 VP.n19 24.5923
R83 VP.n25 VP.n24 24.5923
R84 VP.n59 VP.n7 24.3464
R85 VP.n72 VP.n71 24.3464
R86 VP.n32 VP.n31 24.3464
R87 VP.n20 VP.n19 24.3464
R88 VP.n47 VP.n11 23.8546
R89 VP.n85 VP.n84 23.8546
R90 VP.n45 VP.n44 23.8546
R91 VP.n22 VP.n21 2.54064
R92 VP.n46 VP.n12 0.417304
R93 VP.n49 VP.n48 0.417304
R94 VP.n86 VP.n0 0.417304
R95 VP VP.n86 0.394524
R96 VP.n60 VP.n59 0.246418
R97 VP.n73 VP.n72 0.246418
R98 VP.n33 VP.n32 0.246418
R99 VP.n23 VP.n22 0.189894
R100 VP.n23 VP.n18 0.189894
R101 VP.n27 VP.n18 0.189894
R102 VP.n28 VP.n27 0.189894
R103 VP.n29 VP.n28 0.189894
R104 VP.n29 VP.n16 0.189894
R105 VP.n34 VP.n16 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n14 0.189894
R109 VP.n40 VP.n14 0.189894
R110 VP.n41 VP.n40 0.189894
R111 VP.n42 VP.n41 0.189894
R112 VP.n42 VP.n12 0.189894
R113 VP.n50 VP.n49 0.189894
R114 VP.n50 VP.n10 0.189894
R115 VP.n54 VP.n10 0.189894
R116 VP.n55 VP.n54 0.189894
R117 VP.n56 VP.n55 0.189894
R118 VP.n56 VP.n8 0.189894
R119 VP.n61 VP.n8 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n63 VP.n62 0.189894
R122 VP.n63 VP.n6 0.189894
R123 VP.n67 VP.n6 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n69 VP.n68 0.189894
R126 VP.n69 VP.n4 0.189894
R127 VP.n74 VP.n4 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n76 VP.n75 0.189894
R130 VP.n76 VP.n2 0.189894
R131 VP.n80 VP.n2 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n82 VP.n81 0.189894
R134 VP.n82 VP.n0 0.189894
R135 VDD1 VDD1.n0 66.7707
R136 VDD1.n3 VDD1.n2 66.657
R137 VDD1.n3 VDD1.n1 66.657
R138 VDD1.n5 VDD1.n4 64.9925
R139 VDD1.n5 VDD1.n3 47.1905
R140 VDD1.n4 VDD1.t1 2.30283
R141 VDD1.n4 VDD1.t3 2.30283
R142 VDD1.n0 VDD1.t0 2.30283
R143 VDD1.n0 VDD1.t7 2.30283
R144 VDD1.n2 VDD1.t2 2.30283
R145 VDD1.n2 VDD1.t6 2.30283
R146 VDD1.n1 VDD1.t5 2.30283
R147 VDD1.n1 VDD1.t4 2.30283
R148 VDD1 VDD1.n5 1.66214
R149 VTAIL.n370 VTAIL.n330 289.615
R150 VTAIL.n42 VTAIL.n2 289.615
R151 VTAIL.n88 VTAIL.n48 289.615
R152 VTAIL.n136 VTAIL.n96 289.615
R153 VTAIL.n324 VTAIL.n284 289.615
R154 VTAIL.n276 VTAIL.n236 289.615
R155 VTAIL.n230 VTAIL.n190 289.615
R156 VTAIL.n182 VTAIL.n142 289.615
R157 VTAIL.n345 VTAIL.n344 185
R158 VTAIL.n342 VTAIL.n341 185
R159 VTAIL.n351 VTAIL.n350 185
R160 VTAIL.n353 VTAIL.n352 185
R161 VTAIL.n338 VTAIL.n337 185
R162 VTAIL.n359 VTAIL.n358 185
R163 VTAIL.n362 VTAIL.n361 185
R164 VTAIL.n360 VTAIL.n334 185
R165 VTAIL.n367 VTAIL.n333 185
R166 VTAIL.n369 VTAIL.n368 185
R167 VTAIL.n371 VTAIL.n370 185
R168 VTAIL.n17 VTAIL.n16 185
R169 VTAIL.n14 VTAIL.n13 185
R170 VTAIL.n23 VTAIL.n22 185
R171 VTAIL.n25 VTAIL.n24 185
R172 VTAIL.n10 VTAIL.n9 185
R173 VTAIL.n31 VTAIL.n30 185
R174 VTAIL.n34 VTAIL.n33 185
R175 VTAIL.n32 VTAIL.n6 185
R176 VTAIL.n39 VTAIL.n5 185
R177 VTAIL.n41 VTAIL.n40 185
R178 VTAIL.n43 VTAIL.n42 185
R179 VTAIL.n63 VTAIL.n62 185
R180 VTAIL.n60 VTAIL.n59 185
R181 VTAIL.n69 VTAIL.n68 185
R182 VTAIL.n71 VTAIL.n70 185
R183 VTAIL.n56 VTAIL.n55 185
R184 VTAIL.n77 VTAIL.n76 185
R185 VTAIL.n80 VTAIL.n79 185
R186 VTAIL.n78 VTAIL.n52 185
R187 VTAIL.n85 VTAIL.n51 185
R188 VTAIL.n87 VTAIL.n86 185
R189 VTAIL.n89 VTAIL.n88 185
R190 VTAIL.n111 VTAIL.n110 185
R191 VTAIL.n108 VTAIL.n107 185
R192 VTAIL.n117 VTAIL.n116 185
R193 VTAIL.n119 VTAIL.n118 185
R194 VTAIL.n104 VTAIL.n103 185
R195 VTAIL.n125 VTAIL.n124 185
R196 VTAIL.n128 VTAIL.n127 185
R197 VTAIL.n126 VTAIL.n100 185
R198 VTAIL.n133 VTAIL.n99 185
R199 VTAIL.n135 VTAIL.n134 185
R200 VTAIL.n137 VTAIL.n136 185
R201 VTAIL.n325 VTAIL.n324 185
R202 VTAIL.n323 VTAIL.n322 185
R203 VTAIL.n321 VTAIL.n287 185
R204 VTAIL.n291 VTAIL.n288 185
R205 VTAIL.n316 VTAIL.n315 185
R206 VTAIL.n314 VTAIL.n313 185
R207 VTAIL.n293 VTAIL.n292 185
R208 VTAIL.n308 VTAIL.n307 185
R209 VTAIL.n306 VTAIL.n305 185
R210 VTAIL.n297 VTAIL.n296 185
R211 VTAIL.n300 VTAIL.n299 185
R212 VTAIL.n277 VTAIL.n276 185
R213 VTAIL.n275 VTAIL.n274 185
R214 VTAIL.n273 VTAIL.n239 185
R215 VTAIL.n243 VTAIL.n240 185
R216 VTAIL.n268 VTAIL.n267 185
R217 VTAIL.n266 VTAIL.n265 185
R218 VTAIL.n245 VTAIL.n244 185
R219 VTAIL.n260 VTAIL.n259 185
R220 VTAIL.n258 VTAIL.n257 185
R221 VTAIL.n249 VTAIL.n248 185
R222 VTAIL.n252 VTAIL.n251 185
R223 VTAIL.n231 VTAIL.n230 185
R224 VTAIL.n229 VTAIL.n228 185
R225 VTAIL.n227 VTAIL.n193 185
R226 VTAIL.n197 VTAIL.n194 185
R227 VTAIL.n222 VTAIL.n221 185
R228 VTAIL.n220 VTAIL.n219 185
R229 VTAIL.n199 VTAIL.n198 185
R230 VTAIL.n214 VTAIL.n213 185
R231 VTAIL.n212 VTAIL.n211 185
R232 VTAIL.n203 VTAIL.n202 185
R233 VTAIL.n206 VTAIL.n205 185
R234 VTAIL.n183 VTAIL.n182 185
R235 VTAIL.n181 VTAIL.n180 185
R236 VTAIL.n179 VTAIL.n145 185
R237 VTAIL.n149 VTAIL.n146 185
R238 VTAIL.n174 VTAIL.n173 185
R239 VTAIL.n172 VTAIL.n171 185
R240 VTAIL.n151 VTAIL.n150 185
R241 VTAIL.n166 VTAIL.n165 185
R242 VTAIL.n164 VTAIL.n163 185
R243 VTAIL.n155 VTAIL.n154 185
R244 VTAIL.n158 VTAIL.n157 185
R245 VTAIL.t2 VTAIL.n343 149.524
R246 VTAIL.t6 VTAIL.n15 149.524
R247 VTAIL.t13 VTAIL.n61 149.524
R248 VTAIL.t9 VTAIL.n109 149.524
R249 VTAIL.t11 VTAIL.n298 149.524
R250 VTAIL.t15 VTAIL.n250 149.524
R251 VTAIL.t5 VTAIL.n204 149.524
R252 VTAIL.t3 VTAIL.n156 149.524
R253 VTAIL.n344 VTAIL.n341 104.615
R254 VTAIL.n351 VTAIL.n341 104.615
R255 VTAIL.n352 VTAIL.n351 104.615
R256 VTAIL.n352 VTAIL.n337 104.615
R257 VTAIL.n359 VTAIL.n337 104.615
R258 VTAIL.n361 VTAIL.n359 104.615
R259 VTAIL.n361 VTAIL.n360 104.615
R260 VTAIL.n360 VTAIL.n333 104.615
R261 VTAIL.n369 VTAIL.n333 104.615
R262 VTAIL.n370 VTAIL.n369 104.615
R263 VTAIL.n16 VTAIL.n13 104.615
R264 VTAIL.n23 VTAIL.n13 104.615
R265 VTAIL.n24 VTAIL.n23 104.615
R266 VTAIL.n24 VTAIL.n9 104.615
R267 VTAIL.n31 VTAIL.n9 104.615
R268 VTAIL.n33 VTAIL.n31 104.615
R269 VTAIL.n33 VTAIL.n32 104.615
R270 VTAIL.n32 VTAIL.n5 104.615
R271 VTAIL.n41 VTAIL.n5 104.615
R272 VTAIL.n42 VTAIL.n41 104.615
R273 VTAIL.n62 VTAIL.n59 104.615
R274 VTAIL.n69 VTAIL.n59 104.615
R275 VTAIL.n70 VTAIL.n69 104.615
R276 VTAIL.n70 VTAIL.n55 104.615
R277 VTAIL.n77 VTAIL.n55 104.615
R278 VTAIL.n79 VTAIL.n77 104.615
R279 VTAIL.n79 VTAIL.n78 104.615
R280 VTAIL.n78 VTAIL.n51 104.615
R281 VTAIL.n87 VTAIL.n51 104.615
R282 VTAIL.n88 VTAIL.n87 104.615
R283 VTAIL.n110 VTAIL.n107 104.615
R284 VTAIL.n117 VTAIL.n107 104.615
R285 VTAIL.n118 VTAIL.n117 104.615
R286 VTAIL.n118 VTAIL.n103 104.615
R287 VTAIL.n125 VTAIL.n103 104.615
R288 VTAIL.n127 VTAIL.n125 104.615
R289 VTAIL.n127 VTAIL.n126 104.615
R290 VTAIL.n126 VTAIL.n99 104.615
R291 VTAIL.n135 VTAIL.n99 104.615
R292 VTAIL.n136 VTAIL.n135 104.615
R293 VTAIL.n324 VTAIL.n323 104.615
R294 VTAIL.n323 VTAIL.n287 104.615
R295 VTAIL.n291 VTAIL.n287 104.615
R296 VTAIL.n315 VTAIL.n291 104.615
R297 VTAIL.n315 VTAIL.n314 104.615
R298 VTAIL.n314 VTAIL.n292 104.615
R299 VTAIL.n307 VTAIL.n292 104.615
R300 VTAIL.n307 VTAIL.n306 104.615
R301 VTAIL.n306 VTAIL.n296 104.615
R302 VTAIL.n299 VTAIL.n296 104.615
R303 VTAIL.n276 VTAIL.n275 104.615
R304 VTAIL.n275 VTAIL.n239 104.615
R305 VTAIL.n243 VTAIL.n239 104.615
R306 VTAIL.n267 VTAIL.n243 104.615
R307 VTAIL.n267 VTAIL.n266 104.615
R308 VTAIL.n266 VTAIL.n244 104.615
R309 VTAIL.n259 VTAIL.n244 104.615
R310 VTAIL.n259 VTAIL.n258 104.615
R311 VTAIL.n258 VTAIL.n248 104.615
R312 VTAIL.n251 VTAIL.n248 104.615
R313 VTAIL.n230 VTAIL.n229 104.615
R314 VTAIL.n229 VTAIL.n193 104.615
R315 VTAIL.n197 VTAIL.n193 104.615
R316 VTAIL.n221 VTAIL.n197 104.615
R317 VTAIL.n221 VTAIL.n220 104.615
R318 VTAIL.n220 VTAIL.n198 104.615
R319 VTAIL.n213 VTAIL.n198 104.615
R320 VTAIL.n213 VTAIL.n212 104.615
R321 VTAIL.n212 VTAIL.n202 104.615
R322 VTAIL.n205 VTAIL.n202 104.615
R323 VTAIL.n182 VTAIL.n181 104.615
R324 VTAIL.n181 VTAIL.n145 104.615
R325 VTAIL.n149 VTAIL.n145 104.615
R326 VTAIL.n173 VTAIL.n149 104.615
R327 VTAIL.n173 VTAIL.n172 104.615
R328 VTAIL.n172 VTAIL.n150 104.615
R329 VTAIL.n165 VTAIL.n150 104.615
R330 VTAIL.n165 VTAIL.n164 104.615
R331 VTAIL.n164 VTAIL.n154 104.615
R332 VTAIL.n157 VTAIL.n154 104.615
R333 VTAIL.n344 VTAIL.t2 52.3082
R334 VTAIL.n16 VTAIL.t6 52.3082
R335 VTAIL.n62 VTAIL.t13 52.3082
R336 VTAIL.n110 VTAIL.t9 52.3082
R337 VTAIL.n299 VTAIL.t11 52.3082
R338 VTAIL.n251 VTAIL.t15 52.3082
R339 VTAIL.n205 VTAIL.t5 52.3082
R340 VTAIL.n157 VTAIL.t3 52.3082
R341 VTAIL.n283 VTAIL.n282 48.3139
R342 VTAIL.n189 VTAIL.n188 48.3139
R343 VTAIL.n1 VTAIL.n0 48.3137
R344 VTAIL.n95 VTAIL.n94 48.3137
R345 VTAIL.n375 VTAIL.n374 33.7369
R346 VTAIL.n47 VTAIL.n46 33.7369
R347 VTAIL.n93 VTAIL.n92 33.7369
R348 VTAIL.n141 VTAIL.n140 33.7369
R349 VTAIL.n329 VTAIL.n328 33.7369
R350 VTAIL.n281 VTAIL.n280 33.7369
R351 VTAIL.n235 VTAIL.n234 33.7369
R352 VTAIL.n187 VTAIL.n186 33.7369
R353 VTAIL.n375 VTAIL.n329 23.2203
R354 VTAIL.n187 VTAIL.n141 23.2203
R355 VTAIL.n368 VTAIL.n367 13.1884
R356 VTAIL.n40 VTAIL.n39 13.1884
R357 VTAIL.n86 VTAIL.n85 13.1884
R358 VTAIL.n134 VTAIL.n133 13.1884
R359 VTAIL.n322 VTAIL.n321 13.1884
R360 VTAIL.n274 VTAIL.n273 13.1884
R361 VTAIL.n228 VTAIL.n227 13.1884
R362 VTAIL.n180 VTAIL.n179 13.1884
R363 VTAIL.n366 VTAIL.n334 12.8005
R364 VTAIL.n371 VTAIL.n332 12.8005
R365 VTAIL.n38 VTAIL.n6 12.8005
R366 VTAIL.n43 VTAIL.n4 12.8005
R367 VTAIL.n84 VTAIL.n52 12.8005
R368 VTAIL.n89 VTAIL.n50 12.8005
R369 VTAIL.n132 VTAIL.n100 12.8005
R370 VTAIL.n137 VTAIL.n98 12.8005
R371 VTAIL.n325 VTAIL.n286 12.8005
R372 VTAIL.n320 VTAIL.n288 12.8005
R373 VTAIL.n277 VTAIL.n238 12.8005
R374 VTAIL.n272 VTAIL.n240 12.8005
R375 VTAIL.n231 VTAIL.n192 12.8005
R376 VTAIL.n226 VTAIL.n194 12.8005
R377 VTAIL.n183 VTAIL.n144 12.8005
R378 VTAIL.n178 VTAIL.n146 12.8005
R379 VTAIL.n363 VTAIL.n362 12.0247
R380 VTAIL.n372 VTAIL.n330 12.0247
R381 VTAIL.n35 VTAIL.n34 12.0247
R382 VTAIL.n44 VTAIL.n2 12.0247
R383 VTAIL.n81 VTAIL.n80 12.0247
R384 VTAIL.n90 VTAIL.n48 12.0247
R385 VTAIL.n129 VTAIL.n128 12.0247
R386 VTAIL.n138 VTAIL.n96 12.0247
R387 VTAIL.n326 VTAIL.n284 12.0247
R388 VTAIL.n317 VTAIL.n316 12.0247
R389 VTAIL.n278 VTAIL.n236 12.0247
R390 VTAIL.n269 VTAIL.n268 12.0247
R391 VTAIL.n232 VTAIL.n190 12.0247
R392 VTAIL.n223 VTAIL.n222 12.0247
R393 VTAIL.n184 VTAIL.n142 12.0247
R394 VTAIL.n175 VTAIL.n174 12.0247
R395 VTAIL.n358 VTAIL.n336 11.249
R396 VTAIL.n30 VTAIL.n8 11.249
R397 VTAIL.n76 VTAIL.n54 11.249
R398 VTAIL.n124 VTAIL.n102 11.249
R399 VTAIL.n313 VTAIL.n290 11.249
R400 VTAIL.n265 VTAIL.n242 11.249
R401 VTAIL.n219 VTAIL.n196 11.249
R402 VTAIL.n171 VTAIL.n148 11.249
R403 VTAIL.n357 VTAIL.n338 10.4732
R404 VTAIL.n29 VTAIL.n10 10.4732
R405 VTAIL.n75 VTAIL.n56 10.4732
R406 VTAIL.n123 VTAIL.n104 10.4732
R407 VTAIL.n312 VTAIL.n293 10.4732
R408 VTAIL.n264 VTAIL.n245 10.4732
R409 VTAIL.n218 VTAIL.n199 10.4732
R410 VTAIL.n170 VTAIL.n151 10.4732
R411 VTAIL.n345 VTAIL.n343 10.2747
R412 VTAIL.n17 VTAIL.n15 10.2747
R413 VTAIL.n63 VTAIL.n61 10.2747
R414 VTAIL.n111 VTAIL.n109 10.2747
R415 VTAIL.n300 VTAIL.n298 10.2747
R416 VTAIL.n252 VTAIL.n250 10.2747
R417 VTAIL.n206 VTAIL.n204 10.2747
R418 VTAIL.n158 VTAIL.n156 10.2747
R419 VTAIL.n354 VTAIL.n353 9.69747
R420 VTAIL.n26 VTAIL.n25 9.69747
R421 VTAIL.n72 VTAIL.n71 9.69747
R422 VTAIL.n120 VTAIL.n119 9.69747
R423 VTAIL.n309 VTAIL.n308 9.69747
R424 VTAIL.n261 VTAIL.n260 9.69747
R425 VTAIL.n215 VTAIL.n214 9.69747
R426 VTAIL.n167 VTAIL.n166 9.69747
R427 VTAIL.n374 VTAIL.n373 9.45567
R428 VTAIL.n46 VTAIL.n45 9.45567
R429 VTAIL.n92 VTAIL.n91 9.45567
R430 VTAIL.n140 VTAIL.n139 9.45567
R431 VTAIL.n328 VTAIL.n327 9.45567
R432 VTAIL.n280 VTAIL.n279 9.45567
R433 VTAIL.n234 VTAIL.n233 9.45567
R434 VTAIL.n186 VTAIL.n185 9.45567
R435 VTAIL.n373 VTAIL.n372 9.3005
R436 VTAIL.n332 VTAIL.n331 9.3005
R437 VTAIL.n347 VTAIL.n346 9.3005
R438 VTAIL.n349 VTAIL.n348 9.3005
R439 VTAIL.n340 VTAIL.n339 9.3005
R440 VTAIL.n355 VTAIL.n354 9.3005
R441 VTAIL.n357 VTAIL.n356 9.3005
R442 VTAIL.n336 VTAIL.n335 9.3005
R443 VTAIL.n364 VTAIL.n363 9.3005
R444 VTAIL.n366 VTAIL.n365 9.3005
R445 VTAIL.n45 VTAIL.n44 9.3005
R446 VTAIL.n4 VTAIL.n3 9.3005
R447 VTAIL.n19 VTAIL.n18 9.3005
R448 VTAIL.n21 VTAIL.n20 9.3005
R449 VTAIL.n12 VTAIL.n11 9.3005
R450 VTAIL.n27 VTAIL.n26 9.3005
R451 VTAIL.n29 VTAIL.n28 9.3005
R452 VTAIL.n8 VTAIL.n7 9.3005
R453 VTAIL.n36 VTAIL.n35 9.3005
R454 VTAIL.n38 VTAIL.n37 9.3005
R455 VTAIL.n91 VTAIL.n90 9.3005
R456 VTAIL.n50 VTAIL.n49 9.3005
R457 VTAIL.n65 VTAIL.n64 9.3005
R458 VTAIL.n67 VTAIL.n66 9.3005
R459 VTAIL.n58 VTAIL.n57 9.3005
R460 VTAIL.n73 VTAIL.n72 9.3005
R461 VTAIL.n75 VTAIL.n74 9.3005
R462 VTAIL.n54 VTAIL.n53 9.3005
R463 VTAIL.n82 VTAIL.n81 9.3005
R464 VTAIL.n84 VTAIL.n83 9.3005
R465 VTAIL.n139 VTAIL.n138 9.3005
R466 VTAIL.n98 VTAIL.n97 9.3005
R467 VTAIL.n113 VTAIL.n112 9.3005
R468 VTAIL.n115 VTAIL.n114 9.3005
R469 VTAIL.n106 VTAIL.n105 9.3005
R470 VTAIL.n121 VTAIL.n120 9.3005
R471 VTAIL.n123 VTAIL.n122 9.3005
R472 VTAIL.n102 VTAIL.n101 9.3005
R473 VTAIL.n130 VTAIL.n129 9.3005
R474 VTAIL.n132 VTAIL.n131 9.3005
R475 VTAIL.n302 VTAIL.n301 9.3005
R476 VTAIL.n304 VTAIL.n303 9.3005
R477 VTAIL.n295 VTAIL.n294 9.3005
R478 VTAIL.n310 VTAIL.n309 9.3005
R479 VTAIL.n312 VTAIL.n311 9.3005
R480 VTAIL.n290 VTAIL.n289 9.3005
R481 VTAIL.n318 VTAIL.n317 9.3005
R482 VTAIL.n320 VTAIL.n319 9.3005
R483 VTAIL.n327 VTAIL.n326 9.3005
R484 VTAIL.n286 VTAIL.n285 9.3005
R485 VTAIL.n254 VTAIL.n253 9.3005
R486 VTAIL.n256 VTAIL.n255 9.3005
R487 VTAIL.n247 VTAIL.n246 9.3005
R488 VTAIL.n262 VTAIL.n261 9.3005
R489 VTAIL.n264 VTAIL.n263 9.3005
R490 VTAIL.n242 VTAIL.n241 9.3005
R491 VTAIL.n270 VTAIL.n269 9.3005
R492 VTAIL.n272 VTAIL.n271 9.3005
R493 VTAIL.n279 VTAIL.n278 9.3005
R494 VTAIL.n238 VTAIL.n237 9.3005
R495 VTAIL.n208 VTAIL.n207 9.3005
R496 VTAIL.n210 VTAIL.n209 9.3005
R497 VTAIL.n201 VTAIL.n200 9.3005
R498 VTAIL.n216 VTAIL.n215 9.3005
R499 VTAIL.n218 VTAIL.n217 9.3005
R500 VTAIL.n196 VTAIL.n195 9.3005
R501 VTAIL.n224 VTAIL.n223 9.3005
R502 VTAIL.n226 VTAIL.n225 9.3005
R503 VTAIL.n233 VTAIL.n232 9.3005
R504 VTAIL.n192 VTAIL.n191 9.3005
R505 VTAIL.n160 VTAIL.n159 9.3005
R506 VTAIL.n162 VTAIL.n161 9.3005
R507 VTAIL.n153 VTAIL.n152 9.3005
R508 VTAIL.n168 VTAIL.n167 9.3005
R509 VTAIL.n170 VTAIL.n169 9.3005
R510 VTAIL.n148 VTAIL.n147 9.3005
R511 VTAIL.n176 VTAIL.n175 9.3005
R512 VTAIL.n178 VTAIL.n177 9.3005
R513 VTAIL.n185 VTAIL.n184 9.3005
R514 VTAIL.n144 VTAIL.n143 9.3005
R515 VTAIL.n350 VTAIL.n340 8.92171
R516 VTAIL.n22 VTAIL.n12 8.92171
R517 VTAIL.n68 VTAIL.n58 8.92171
R518 VTAIL.n116 VTAIL.n106 8.92171
R519 VTAIL.n305 VTAIL.n295 8.92171
R520 VTAIL.n257 VTAIL.n247 8.92171
R521 VTAIL.n211 VTAIL.n201 8.92171
R522 VTAIL.n163 VTAIL.n153 8.92171
R523 VTAIL.n349 VTAIL.n342 8.14595
R524 VTAIL.n21 VTAIL.n14 8.14595
R525 VTAIL.n67 VTAIL.n60 8.14595
R526 VTAIL.n115 VTAIL.n108 8.14595
R527 VTAIL.n304 VTAIL.n297 8.14595
R528 VTAIL.n256 VTAIL.n249 8.14595
R529 VTAIL.n210 VTAIL.n203 8.14595
R530 VTAIL.n162 VTAIL.n155 8.14595
R531 VTAIL.n346 VTAIL.n345 7.3702
R532 VTAIL.n18 VTAIL.n17 7.3702
R533 VTAIL.n64 VTAIL.n63 7.3702
R534 VTAIL.n112 VTAIL.n111 7.3702
R535 VTAIL.n301 VTAIL.n300 7.3702
R536 VTAIL.n253 VTAIL.n252 7.3702
R537 VTAIL.n207 VTAIL.n206 7.3702
R538 VTAIL.n159 VTAIL.n158 7.3702
R539 VTAIL.n346 VTAIL.n342 5.81868
R540 VTAIL.n18 VTAIL.n14 5.81868
R541 VTAIL.n64 VTAIL.n60 5.81868
R542 VTAIL.n112 VTAIL.n108 5.81868
R543 VTAIL.n301 VTAIL.n297 5.81868
R544 VTAIL.n253 VTAIL.n249 5.81868
R545 VTAIL.n207 VTAIL.n203 5.81868
R546 VTAIL.n159 VTAIL.n155 5.81868
R547 VTAIL.n350 VTAIL.n349 5.04292
R548 VTAIL.n22 VTAIL.n21 5.04292
R549 VTAIL.n68 VTAIL.n67 5.04292
R550 VTAIL.n116 VTAIL.n115 5.04292
R551 VTAIL.n305 VTAIL.n304 5.04292
R552 VTAIL.n257 VTAIL.n256 5.04292
R553 VTAIL.n211 VTAIL.n210 5.04292
R554 VTAIL.n163 VTAIL.n162 5.04292
R555 VTAIL.n353 VTAIL.n340 4.26717
R556 VTAIL.n25 VTAIL.n12 4.26717
R557 VTAIL.n71 VTAIL.n58 4.26717
R558 VTAIL.n119 VTAIL.n106 4.26717
R559 VTAIL.n308 VTAIL.n295 4.26717
R560 VTAIL.n260 VTAIL.n247 4.26717
R561 VTAIL.n214 VTAIL.n201 4.26717
R562 VTAIL.n166 VTAIL.n153 4.26717
R563 VTAIL.n354 VTAIL.n338 3.49141
R564 VTAIL.n26 VTAIL.n10 3.49141
R565 VTAIL.n72 VTAIL.n56 3.49141
R566 VTAIL.n120 VTAIL.n104 3.49141
R567 VTAIL.n309 VTAIL.n293 3.49141
R568 VTAIL.n261 VTAIL.n245 3.49141
R569 VTAIL.n215 VTAIL.n199 3.49141
R570 VTAIL.n167 VTAIL.n151 3.49141
R571 VTAIL.n189 VTAIL.n187 3.44016
R572 VTAIL.n235 VTAIL.n189 3.44016
R573 VTAIL.n283 VTAIL.n281 3.44016
R574 VTAIL.n329 VTAIL.n283 3.44016
R575 VTAIL.n141 VTAIL.n95 3.44016
R576 VTAIL.n95 VTAIL.n93 3.44016
R577 VTAIL.n47 VTAIL.n1 3.44016
R578 VTAIL VTAIL.n375 3.38197
R579 VTAIL.n347 VTAIL.n343 2.84303
R580 VTAIL.n19 VTAIL.n15 2.84303
R581 VTAIL.n65 VTAIL.n61 2.84303
R582 VTAIL.n113 VTAIL.n109 2.84303
R583 VTAIL.n302 VTAIL.n298 2.84303
R584 VTAIL.n254 VTAIL.n250 2.84303
R585 VTAIL.n208 VTAIL.n204 2.84303
R586 VTAIL.n160 VTAIL.n156 2.84303
R587 VTAIL.n358 VTAIL.n357 2.71565
R588 VTAIL.n30 VTAIL.n29 2.71565
R589 VTAIL.n76 VTAIL.n75 2.71565
R590 VTAIL.n124 VTAIL.n123 2.71565
R591 VTAIL.n313 VTAIL.n312 2.71565
R592 VTAIL.n265 VTAIL.n264 2.71565
R593 VTAIL.n219 VTAIL.n218 2.71565
R594 VTAIL.n171 VTAIL.n170 2.71565
R595 VTAIL.n0 VTAIL.t7 2.30283
R596 VTAIL.n0 VTAIL.t1 2.30283
R597 VTAIL.n94 VTAIL.t8 2.30283
R598 VTAIL.n94 VTAIL.t14 2.30283
R599 VTAIL.n282 VTAIL.t12 2.30283
R600 VTAIL.n282 VTAIL.t10 2.30283
R601 VTAIL.n188 VTAIL.t4 2.30283
R602 VTAIL.n188 VTAIL.t0 2.30283
R603 VTAIL.n362 VTAIL.n336 1.93989
R604 VTAIL.n374 VTAIL.n330 1.93989
R605 VTAIL.n34 VTAIL.n8 1.93989
R606 VTAIL.n46 VTAIL.n2 1.93989
R607 VTAIL.n80 VTAIL.n54 1.93989
R608 VTAIL.n92 VTAIL.n48 1.93989
R609 VTAIL.n128 VTAIL.n102 1.93989
R610 VTAIL.n140 VTAIL.n96 1.93989
R611 VTAIL.n328 VTAIL.n284 1.93989
R612 VTAIL.n316 VTAIL.n290 1.93989
R613 VTAIL.n280 VTAIL.n236 1.93989
R614 VTAIL.n268 VTAIL.n242 1.93989
R615 VTAIL.n234 VTAIL.n190 1.93989
R616 VTAIL.n222 VTAIL.n196 1.93989
R617 VTAIL.n186 VTAIL.n142 1.93989
R618 VTAIL.n174 VTAIL.n148 1.93989
R619 VTAIL.n363 VTAIL.n334 1.16414
R620 VTAIL.n372 VTAIL.n371 1.16414
R621 VTAIL.n35 VTAIL.n6 1.16414
R622 VTAIL.n44 VTAIL.n43 1.16414
R623 VTAIL.n81 VTAIL.n52 1.16414
R624 VTAIL.n90 VTAIL.n89 1.16414
R625 VTAIL.n129 VTAIL.n100 1.16414
R626 VTAIL.n138 VTAIL.n137 1.16414
R627 VTAIL.n326 VTAIL.n325 1.16414
R628 VTAIL.n317 VTAIL.n288 1.16414
R629 VTAIL.n278 VTAIL.n277 1.16414
R630 VTAIL.n269 VTAIL.n240 1.16414
R631 VTAIL.n232 VTAIL.n231 1.16414
R632 VTAIL.n223 VTAIL.n194 1.16414
R633 VTAIL.n184 VTAIL.n183 1.16414
R634 VTAIL.n175 VTAIL.n146 1.16414
R635 VTAIL.n281 VTAIL.n235 0.470328
R636 VTAIL.n93 VTAIL.n47 0.470328
R637 VTAIL.n367 VTAIL.n366 0.388379
R638 VTAIL.n368 VTAIL.n332 0.388379
R639 VTAIL.n39 VTAIL.n38 0.388379
R640 VTAIL.n40 VTAIL.n4 0.388379
R641 VTAIL.n85 VTAIL.n84 0.388379
R642 VTAIL.n86 VTAIL.n50 0.388379
R643 VTAIL.n133 VTAIL.n132 0.388379
R644 VTAIL.n134 VTAIL.n98 0.388379
R645 VTAIL.n322 VTAIL.n286 0.388379
R646 VTAIL.n321 VTAIL.n320 0.388379
R647 VTAIL.n274 VTAIL.n238 0.388379
R648 VTAIL.n273 VTAIL.n272 0.388379
R649 VTAIL.n228 VTAIL.n192 0.388379
R650 VTAIL.n227 VTAIL.n226 0.388379
R651 VTAIL.n180 VTAIL.n144 0.388379
R652 VTAIL.n179 VTAIL.n178 0.388379
R653 VTAIL.n348 VTAIL.n347 0.155672
R654 VTAIL.n348 VTAIL.n339 0.155672
R655 VTAIL.n355 VTAIL.n339 0.155672
R656 VTAIL.n356 VTAIL.n355 0.155672
R657 VTAIL.n356 VTAIL.n335 0.155672
R658 VTAIL.n364 VTAIL.n335 0.155672
R659 VTAIL.n365 VTAIL.n364 0.155672
R660 VTAIL.n365 VTAIL.n331 0.155672
R661 VTAIL.n373 VTAIL.n331 0.155672
R662 VTAIL.n20 VTAIL.n19 0.155672
R663 VTAIL.n20 VTAIL.n11 0.155672
R664 VTAIL.n27 VTAIL.n11 0.155672
R665 VTAIL.n28 VTAIL.n27 0.155672
R666 VTAIL.n28 VTAIL.n7 0.155672
R667 VTAIL.n36 VTAIL.n7 0.155672
R668 VTAIL.n37 VTAIL.n36 0.155672
R669 VTAIL.n37 VTAIL.n3 0.155672
R670 VTAIL.n45 VTAIL.n3 0.155672
R671 VTAIL.n66 VTAIL.n65 0.155672
R672 VTAIL.n66 VTAIL.n57 0.155672
R673 VTAIL.n73 VTAIL.n57 0.155672
R674 VTAIL.n74 VTAIL.n73 0.155672
R675 VTAIL.n74 VTAIL.n53 0.155672
R676 VTAIL.n82 VTAIL.n53 0.155672
R677 VTAIL.n83 VTAIL.n82 0.155672
R678 VTAIL.n83 VTAIL.n49 0.155672
R679 VTAIL.n91 VTAIL.n49 0.155672
R680 VTAIL.n114 VTAIL.n113 0.155672
R681 VTAIL.n114 VTAIL.n105 0.155672
R682 VTAIL.n121 VTAIL.n105 0.155672
R683 VTAIL.n122 VTAIL.n121 0.155672
R684 VTAIL.n122 VTAIL.n101 0.155672
R685 VTAIL.n130 VTAIL.n101 0.155672
R686 VTAIL.n131 VTAIL.n130 0.155672
R687 VTAIL.n131 VTAIL.n97 0.155672
R688 VTAIL.n139 VTAIL.n97 0.155672
R689 VTAIL.n327 VTAIL.n285 0.155672
R690 VTAIL.n319 VTAIL.n285 0.155672
R691 VTAIL.n319 VTAIL.n318 0.155672
R692 VTAIL.n318 VTAIL.n289 0.155672
R693 VTAIL.n311 VTAIL.n289 0.155672
R694 VTAIL.n311 VTAIL.n310 0.155672
R695 VTAIL.n310 VTAIL.n294 0.155672
R696 VTAIL.n303 VTAIL.n294 0.155672
R697 VTAIL.n303 VTAIL.n302 0.155672
R698 VTAIL.n279 VTAIL.n237 0.155672
R699 VTAIL.n271 VTAIL.n237 0.155672
R700 VTAIL.n271 VTAIL.n270 0.155672
R701 VTAIL.n270 VTAIL.n241 0.155672
R702 VTAIL.n263 VTAIL.n241 0.155672
R703 VTAIL.n263 VTAIL.n262 0.155672
R704 VTAIL.n262 VTAIL.n246 0.155672
R705 VTAIL.n255 VTAIL.n246 0.155672
R706 VTAIL.n255 VTAIL.n254 0.155672
R707 VTAIL.n233 VTAIL.n191 0.155672
R708 VTAIL.n225 VTAIL.n191 0.155672
R709 VTAIL.n225 VTAIL.n224 0.155672
R710 VTAIL.n224 VTAIL.n195 0.155672
R711 VTAIL.n217 VTAIL.n195 0.155672
R712 VTAIL.n217 VTAIL.n216 0.155672
R713 VTAIL.n216 VTAIL.n200 0.155672
R714 VTAIL.n209 VTAIL.n200 0.155672
R715 VTAIL.n209 VTAIL.n208 0.155672
R716 VTAIL.n185 VTAIL.n143 0.155672
R717 VTAIL.n177 VTAIL.n143 0.155672
R718 VTAIL.n177 VTAIL.n176 0.155672
R719 VTAIL.n176 VTAIL.n147 0.155672
R720 VTAIL.n169 VTAIL.n147 0.155672
R721 VTAIL.n169 VTAIL.n168 0.155672
R722 VTAIL.n168 VTAIL.n152 0.155672
R723 VTAIL.n161 VTAIL.n152 0.155672
R724 VTAIL.n161 VTAIL.n160 0.155672
R725 VTAIL VTAIL.n1 0.0586897
R726 B.n912 B.n911 585
R727 B.n913 B.n912 585
R728 B.n305 B.n159 585
R729 B.n304 B.n303 585
R730 B.n302 B.n301 585
R731 B.n300 B.n299 585
R732 B.n298 B.n297 585
R733 B.n296 B.n295 585
R734 B.n294 B.n293 585
R735 B.n292 B.n291 585
R736 B.n290 B.n289 585
R737 B.n288 B.n287 585
R738 B.n286 B.n285 585
R739 B.n284 B.n283 585
R740 B.n282 B.n281 585
R741 B.n280 B.n279 585
R742 B.n278 B.n277 585
R743 B.n276 B.n275 585
R744 B.n274 B.n273 585
R745 B.n272 B.n271 585
R746 B.n270 B.n269 585
R747 B.n268 B.n267 585
R748 B.n266 B.n265 585
R749 B.n264 B.n263 585
R750 B.n262 B.n261 585
R751 B.n260 B.n259 585
R752 B.n258 B.n257 585
R753 B.n256 B.n255 585
R754 B.n254 B.n253 585
R755 B.n252 B.n251 585
R756 B.n250 B.n249 585
R757 B.n248 B.n247 585
R758 B.n246 B.n245 585
R759 B.n243 B.n242 585
R760 B.n241 B.n240 585
R761 B.n239 B.n238 585
R762 B.n237 B.n236 585
R763 B.n235 B.n234 585
R764 B.n233 B.n232 585
R765 B.n231 B.n230 585
R766 B.n229 B.n228 585
R767 B.n227 B.n226 585
R768 B.n225 B.n224 585
R769 B.n223 B.n222 585
R770 B.n221 B.n220 585
R771 B.n219 B.n218 585
R772 B.n217 B.n216 585
R773 B.n215 B.n214 585
R774 B.n213 B.n212 585
R775 B.n211 B.n210 585
R776 B.n209 B.n208 585
R777 B.n207 B.n206 585
R778 B.n205 B.n204 585
R779 B.n203 B.n202 585
R780 B.n201 B.n200 585
R781 B.n199 B.n198 585
R782 B.n197 B.n196 585
R783 B.n195 B.n194 585
R784 B.n193 B.n192 585
R785 B.n191 B.n190 585
R786 B.n189 B.n188 585
R787 B.n187 B.n186 585
R788 B.n185 B.n184 585
R789 B.n183 B.n182 585
R790 B.n181 B.n180 585
R791 B.n179 B.n178 585
R792 B.n177 B.n176 585
R793 B.n175 B.n174 585
R794 B.n173 B.n172 585
R795 B.n171 B.n170 585
R796 B.n169 B.n168 585
R797 B.n167 B.n166 585
R798 B.n123 B.n122 585
R799 B.n916 B.n915 585
R800 B.n910 B.n160 585
R801 B.n160 B.n120 585
R802 B.n909 B.n119 585
R803 B.n920 B.n119 585
R804 B.n908 B.n118 585
R805 B.n921 B.n118 585
R806 B.n907 B.n117 585
R807 B.n922 B.n117 585
R808 B.n906 B.n905 585
R809 B.n905 B.n113 585
R810 B.n904 B.n112 585
R811 B.n928 B.n112 585
R812 B.n903 B.n111 585
R813 B.n929 B.n111 585
R814 B.n902 B.n110 585
R815 B.n930 B.n110 585
R816 B.n901 B.n900 585
R817 B.n900 B.n106 585
R818 B.n899 B.n105 585
R819 B.n936 B.n105 585
R820 B.n898 B.n104 585
R821 B.n937 B.n104 585
R822 B.n897 B.n103 585
R823 B.n938 B.n103 585
R824 B.n896 B.n895 585
R825 B.n895 B.n99 585
R826 B.n894 B.n98 585
R827 B.n944 B.n98 585
R828 B.n893 B.n97 585
R829 B.n945 B.n97 585
R830 B.n892 B.n96 585
R831 B.n946 B.n96 585
R832 B.n891 B.n890 585
R833 B.n890 B.n92 585
R834 B.n889 B.n91 585
R835 B.n952 B.n91 585
R836 B.n888 B.n90 585
R837 B.n953 B.n90 585
R838 B.n887 B.n89 585
R839 B.n954 B.n89 585
R840 B.n886 B.n885 585
R841 B.n885 B.n85 585
R842 B.n884 B.n84 585
R843 B.n960 B.n84 585
R844 B.n883 B.n83 585
R845 B.n961 B.n83 585
R846 B.n882 B.n82 585
R847 B.n962 B.n82 585
R848 B.n881 B.n880 585
R849 B.n880 B.n81 585
R850 B.n879 B.n77 585
R851 B.n968 B.n77 585
R852 B.n878 B.n76 585
R853 B.n969 B.n76 585
R854 B.n877 B.n75 585
R855 B.n970 B.n75 585
R856 B.n876 B.n875 585
R857 B.n875 B.n71 585
R858 B.n874 B.n70 585
R859 B.n976 B.n70 585
R860 B.n873 B.n69 585
R861 B.n977 B.n69 585
R862 B.n872 B.n68 585
R863 B.n978 B.n68 585
R864 B.n871 B.n870 585
R865 B.n870 B.n64 585
R866 B.n869 B.n63 585
R867 B.n984 B.n63 585
R868 B.n868 B.n62 585
R869 B.n985 B.n62 585
R870 B.n867 B.n61 585
R871 B.n986 B.n61 585
R872 B.n866 B.n865 585
R873 B.n865 B.n60 585
R874 B.n864 B.n56 585
R875 B.n992 B.n56 585
R876 B.n863 B.n55 585
R877 B.n993 B.n55 585
R878 B.n862 B.n54 585
R879 B.n994 B.n54 585
R880 B.n861 B.n860 585
R881 B.n860 B.n50 585
R882 B.n859 B.n49 585
R883 B.n1000 B.n49 585
R884 B.n858 B.n48 585
R885 B.n1001 B.n48 585
R886 B.n857 B.n47 585
R887 B.n1002 B.n47 585
R888 B.n856 B.n855 585
R889 B.n855 B.n43 585
R890 B.n854 B.n42 585
R891 B.n1008 B.n42 585
R892 B.n853 B.n41 585
R893 B.n1009 B.n41 585
R894 B.n852 B.n40 585
R895 B.n1010 B.n40 585
R896 B.n851 B.n850 585
R897 B.n850 B.n36 585
R898 B.n849 B.n35 585
R899 B.n1016 B.n35 585
R900 B.n848 B.n34 585
R901 B.n1017 B.n34 585
R902 B.n847 B.n33 585
R903 B.n1018 B.n33 585
R904 B.n846 B.n845 585
R905 B.n845 B.n29 585
R906 B.n844 B.n28 585
R907 B.n1024 B.n28 585
R908 B.n843 B.n27 585
R909 B.n1025 B.n27 585
R910 B.n842 B.n26 585
R911 B.n1026 B.n26 585
R912 B.n841 B.n840 585
R913 B.n840 B.n22 585
R914 B.n839 B.n21 585
R915 B.n1032 B.n21 585
R916 B.n838 B.n20 585
R917 B.n1033 B.n20 585
R918 B.n837 B.n19 585
R919 B.n1034 B.n19 585
R920 B.n836 B.n835 585
R921 B.n835 B.n15 585
R922 B.n834 B.n14 585
R923 B.n1040 B.n14 585
R924 B.n833 B.n13 585
R925 B.n1041 B.n13 585
R926 B.n832 B.n12 585
R927 B.n1042 B.n12 585
R928 B.n831 B.n830 585
R929 B.n830 B.n8 585
R930 B.n829 B.n7 585
R931 B.n1048 B.n7 585
R932 B.n828 B.n6 585
R933 B.n1049 B.n6 585
R934 B.n827 B.n5 585
R935 B.n1050 B.n5 585
R936 B.n826 B.n825 585
R937 B.n825 B.n4 585
R938 B.n824 B.n306 585
R939 B.n824 B.n823 585
R940 B.n814 B.n307 585
R941 B.n308 B.n307 585
R942 B.n816 B.n815 585
R943 B.n817 B.n816 585
R944 B.n813 B.n313 585
R945 B.n313 B.n312 585
R946 B.n812 B.n811 585
R947 B.n811 B.n810 585
R948 B.n315 B.n314 585
R949 B.n316 B.n315 585
R950 B.n803 B.n802 585
R951 B.n804 B.n803 585
R952 B.n801 B.n321 585
R953 B.n321 B.n320 585
R954 B.n800 B.n799 585
R955 B.n799 B.n798 585
R956 B.n323 B.n322 585
R957 B.n324 B.n323 585
R958 B.n791 B.n790 585
R959 B.n792 B.n791 585
R960 B.n789 B.n329 585
R961 B.n329 B.n328 585
R962 B.n788 B.n787 585
R963 B.n787 B.n786 585
R964 B.n331 B.n330 585
R965 B.n332 B.n331 585
R966 B.n779 B.n778 585
R967 B.n780 B.n779 585
R968 B.n777 B.n337 585
R969 B.n337 B.n336 585
R970 B.n776 B.n775 585
R971 B.n775 B.n774 585
R972 B.n339 B.n338 585
R973 B.n340 B.n339 585
R974 B.n767 B.n766 585
R975 B.n768 B.n767 585
R976 B.n765 B.n345 585
R977 B.n345 B.n344 585
R978 B.n764 B.n763 585
R979 B.n763 B.n762 585
R980 B.n347 B.n346 585
R981 B.n348 B.n347 585
R982 B.n755 B.n754 585
R983 B.n756 B.n755 585
R984 B.n753 B.n353 585
R985 B.n353 B.n352 585
R986 B.n752 B.n751 585
R987 B.n751 B.n750 585
R988 B.n355 B.n354 585
R989 B.n356 B.n355 585
R990 B.n743 B.n742 585
R991 B.n744 B.n743 585
R992 B.n741 B.n361 585
R993 B.n361 B.n360 585
R994 B.n740 B.n739 585
R995 B.n739 B.n738 585
R996 B.n363 B.n362 585
R997 B.n731 B.n363 585
R998 B.n730 B.n729 585
R999 B.n732 B.n730 585
R1000 B.n728 B.n368 585
R1001 B.n368 B.n367 585
R1002 B.n727 B.n726 585
R1003 B.n726 B.n725 585
R1004 B.n370 B.n369 585
R1005 B.n371 B.n370 585
R1006 B.n718 B.n717 585
R1007 B.n719 B.n718 585
R1008 B.n716 B.n376 585
R1009 B.n376 B.n375 585
R1010 B.n715 B.n714 585
R1011 B.n714 B.n713 585
R1012 B.n378 B.n377 585
R1013 B.n379 B.n378 585
R1014 B.n706 B.n705 585
R1015 B.n707 B.n706 585
R1016 B.n704 B.n384 585
R1017 B.n384 B.n383 585
R1018 B.n703 B.n702 585
R1019 B.n702 B.n701 585
R1020 B.n386 B.n385 585
R1021 B.n694 B.n386 585
R1022 B.n693 B.n692 585
R1023 B.n695 B.n693 585
R1024 B.n691 B.n391 585
R1025 B.n391 B.n390 585
R1026 B.n690 B.n689 585
R1027 B.n689 B.n688 585
R1028 B.n393 B.n392 585
R1029 B.n394 B.n393 585
R1030 B.n681 B.n680 585
R1031 B.n682 B.n681 585
R1032 B.n679 B.n399 585
R1033 B.n399 B.n398 585
R1034 B.n678 B.n677 585
R1035 B.n677 B.n676 585
R1036 B.n401 B.n400 585
R1037 B.n402 B.n401 585
R1038 B.n669 B.n668 585
R1039 B.n670 B.n669 585
R1040 B.n667 B.n407 585
R1041 B.n407 B.n406 585
R1042 B.n666 B.n665 585
R1043 B.n665 B.n664 585
R1044 B.n409 B.n408 585
R1045 B.n410 B.n409 585
R1046 B.n657 B.n656 585
R1047 B.n658 B.n657 585
R1048 B.n655 B.n415 585
R1049 B.n415 B.n414 585
R1050 B.n654 B.n653 585
R1051 B.n653 B.n652 585
R1052 B.n417 B.n416 585
R1053 B.n418 B.n417 585
R1054 B.n645 B.n644 585
R1055 B.n646 B.n645 585
R1056 B.n643 B.n423 585
R1057 B.n423 B.n422 585
R1058 B.n642 B.n641 585
R1059 B.n641 B.n640 585
R1060 B.n425 B.n424 585
R1061 B.n426 B.n425 585
R1062 B.n633 B.n632 585
R1063 B.n634 B.n633 585
R1064 B.n631 B.n431 585
R1065 B.n431 B.n430 585
R1066 B.n630 B.n629 585
R1067 B.n629 B.n628 585
R1068 B.n433 B.n432 585
R1069 B.n434 B.n433 585
R1070 B.n624 B.n623 585
R1071 B.n437 B.n436 585
R1072 B.n620 B.n619 585
R1073 B.n621 B.n620 585
R1074 B.n618 B.n473 585
R1075 B.n617 B.n616 585
R1076 B.n615 B.n614 585
R1077 B.n613 B.n612 585
R1078 B.n611 B.n610 585
R1079 B.n609 B.n608 585
R1080 B.n607 B.n606 585
R1081 B.n605 B.n604 585
R1082 B.n603 B.n602 585
R1083 B.n601 B.n600 585
R1084 B.n599 B.n598 585
R1085 B.n597 B.n596 585
R1086 B.n595 B.n594 585
R1087 B.n593 B.n592 585
R1088 B.n591 B.n590 585
R1089 B.n589 B.n588 585
R1090 B.n587 B.n586 585
R1091 B.n585 B.n584 585
R1092 B.n583 B.n582 585
R1093 B.n581 B.n580 585
R1094 B.n579 B.n578 585
R1095 B.n577 B.n576 585
R1096 B.n575 B.n574 585
R1097 B.n573 B.n572 585
R1098 B.n571 B.n570 585
R1099 B.n569 B.n568 585
R1100 B.n567 B.n566 585
R1101 B.n565 B.n564 585
R1102 B.n563 B.n562 585
R1103 B.n560 B.n559 585
R1104 B.n558 B.n557 585
R1105 B.n556 B.n555 585
R1106 B.n554 B.n553 585
R1107 B.n552 B.n551 585
R1108 B.n550 B.n549 585
R1109 B.n548 B.n547 585
R1110 B.n546 B.n545 585
R1111 B.n544 B.n543 585
R1112 B.n542 B.n541 585
R1113 B.n540 B.n539 585
R1114 B.n538 B.n537 585
R1115 B.n536 B.n535 585
R1116 B.n534 B.n533 585
R1117 B.n532 B.n531 585
R1118 B.n530 B.n529 585
R1119 B.n528 B.n527 585
R1120 B.n526 B.n525 585
R1121 B.n524 B.n523 585
R1122 B.n522 B.n521 585
R1123 B.n520 B.n519 585
R1124 B.n518 B.n517 585
R1125 B.n516 B.n515 585
R1126 B.n514 B.n513 585
R1127 B.n512 B.n511 585
R1128 B.n510 B.n509 585
R1129 B.n508 B.n507 585
R1130 B.n506 B.n505 585
R1131 B.n504 B.n503 585
R1132 B.n502 B.n501 585
R1133 B.n500 B.n499 585
R1134 B.n498 B.n497 585
R1135 B.n496 B.n495 585
R1136 B.n494 B.n493 585
R1137 B.n492 B.n491 585
R1138 B.n490 B.n489 585
R1139 B.n488 B.n487 585
R1140 B.n486 B.n485 585
R1141 B.n484 B.n483 585
R1142 B.n482 B.n481 585
R1143 B.n480 B.n479 585
R1144 B.n625 B.n435 585
R1145 B.n435 B.n434 585
R1146 B.n627 B.n626 585
R1147 B.n628 B.n627 585
R1148 B.n429 B.n428 585
R1149 B.n430 B.n429 585
R1150 B.n636 B.n635 585
R1151 B.n635 B.n634 585
R1152 B.n637 B.n427 585
R1153 B.n427 B.n426 585
R1154 B.n639 B.n638 585
R1155 B.n640 B.n639 585
R1156 B.n421 B.n420 585
R1157 B.n422 B.n421 585
R1158 B.n648 B.n647 585
R1159 B.n647 B.n646 585
R1160 B.n649 B.n419 585
R1161 B.n419 B.n418 585
R1162 B.n651 B.n650 585
R1163 B.n652 B.n651 585
R1164 B.n413 B.n412 585
R1165 B.n414 B.n413 585
R1166 B.n660 B.n659 585
R1167 B.n659 B.n658 585
R1168 B.n661 B.n411 585
R1169 B.n411 B.n410 585
R1170 B.n663 B.n662 585
R1171 B.n664 B.n663 585
R1172 B.n405 B.n404 585
R1173 B.n406 B.n405 585
R1174 B.n672 B.n671 585
R1175 B.n671 B.n670 585
R1176 B.n673 B.n403 585
R1177 B.n403 B.n402 585
R1178 B.n675 B.n674 585
R1179 B.n676 B.n675 585
R1180 B.n397 B.n396 585
R1181 B.n398 B.n397 585
R1182 B.n684 B.n683 585
R1183 B.n683 B.n682 585
R1184 B.n685 B.n395 585
R1185 B.n395 B.n394 585
R1186 B.n687 B.n686 585
R1187 B.n688 B.n687 585
R1188 B.n389 B.n388 585
R1189 B.n390 B.n389 585
R1190 B.n697 B.n696 585
R1191 B.n696 B.n695 585
R1192 B.n698 B.n387 585
R1193 B.n694 B.n387 585
R1194 B.n700 B.n699 585
R1195 B.n701 B.n700 585
R1196 B.n382 B.n381 585
R1197 B.n383 B.n382 585
R1198 B.n709 B.n708 585
R1199 B.n708 B.n707 585
R1200 B.n710 B.n380 585
R1201 B.n380 B.n379 585
R1202 B.n712 B.n711 585
R1203 B.n713 B.n712 585
R1204 B.n374 B.n373 585
R1205 B.n375 B.n374 585
R1206 B.n721 B.n720 585
R1207 B.n720 B.n719 585
R1208 B.n722 B.n372 585
R1209 B.n372 B.n371 585
R1210 B.n724 B.n723 585
R1211 B.n725 B.n724 585
R1212 B.n366 B.n365 585
R1213 B.n367 B.n366 585
R1214 B.n734 B.n733 585
R1215 B.n733 B.n732 585
R1216 B.n735 B.n364 585
R1217 B.n731 B.n364 585
R1218 B.n737 B.n736 585
R1219 B.n738 B.n737 585
R1220 B.n359 B.n358 585
R1221 B.n360 B.n359 585
R1222 B.n746 B.n745 585
R1223 B.n745 B.n744 585
R1224 B.n747 B.n357 585
R1225 B.n357 B.n356 585
R1226 B.n749 B.n748 585
R1227 B.n750 B.n749 585
R1228 B.n351 B.n350 585
R1229 B.n352 B.n351 585
R1230 B.n758 B.n757 585
R1231 B.n757 B.n756 585
R1232 B.n759 B.n349 585
R1233 B.n349 B.n348 585
R1234 B.n761 B.n760 585
R1235 B.n762 B.n761 585
R1236 B.n343 B.n342 585
R1237 B.n344 B.n343 585
R1238 B.n770 B.n769 585
R1239 B.n769 B.n768 585
R1240 B.n771 B.n341 585
R1241 B.n341 B.n340 585
R1242 B.n773 B.n772 585
R1243 B.n774 B.n773 585
R1244 B.n335 B.n334 585
R1245 B.n336 B.n335 585
R1246 B.n782 B.n781 585
R1247 B.n781 B.n780 585
R1248 B.n783 B.n333 585
R1249 B.n333 B.n332 585
R1250 B.n785 B.n784 585
R1251 B.n786 B.n785 585
R1252 B.n327 B.n326 585
R1253 B.n328 B.n327 585
R1254 B.n794 B.n793 585
R1255 B.n793 B.n792 585
R1256 B.n795 B.n325 585
R1257 B.n325 B.n324 585
R1258 B.n797 B.n796 585
R1259 B.n798 B.n797 585
R1260 B.n319 B.n318 585
R1261 B.n320 B.n319 585
R1262 B.n806 B.n805 585
R1263 B.n805 B.n804 585
R1264 B.n807 B.n317 585
R1265 B.n317 B.n316 585
R1266 B.n809 B.n808 585
R1267 B.n810 B.n809 585
R1268 B.n311 B.n310 585
R1269 B.n312 B.n311 585
R1270 B.n819 B.n818 585
R1271 B.n818 B.n817 585
R1272 B.n820 B.n309 585
R1273 B.n309 B.n308 585
R1274 B.n822 B.n821 585
R1275 B.n823 B.n822 585
R1276 B.n2 B.n0 585
R1277 B.n4 B.n2 585
R1278 B.n3 B.n1 585
R1279 B.n1049 B.n3 585
R1280 B.n1047 B.n1046 585
R1281 B.n1048 B.n1047 585
R1282 B.n1045 B.n9 585
R1283 B.n9 B.n8 585
R1284 B.n1044 B.n1043 585
R1285 B.n1043 B.n1042 585
R1286 B.n11 B.n10 585
R1287 B.n1041 B.n11 585
R1288 B.n1039 B.n1038 585
R1289 B.n1040 B.n1039 585
R1290 B.n1037 B.n16 585
R1291 B.n16 B.n15 585
R1292 B.n1036 B.n1035 585
R1293 B.n1035 B.n1034 585
R1294 B.n18 B.n17 585
R1295 B.n1033 B.n18 585
R1296 B.n1031 B.n1030 585
R1297 B.n1032 B.n1031 585
R1298 B.n1029 B.n23 585
R1299 B.n23 B.n22 585
R1300 B.n1028 B.n1027 585
R1301 B.n1027 B.n1026 585
R1302 B.n25 B.n24 585
R1303 B.n1025 B.n25 585
R1304 B.n1023 B.n1022 585
R1305 B.n1024 B.n1023 585
R1306 B.n1021 B.n30 585
R1307 B.n30 B.n29 585
R1308 B.n1020 B.n1019 585
R1309 B.n1019 B.n1018 585
R1310 B.n32 B.n31 585
R1311 B.n1017 B.n32 585
R1312 B.n1015 B.n1014 585
R1313 B.n1016 B.n1015 585
R1314 B.n1013 B.n37 585
R1315 B.n37 B.n36 585
R1316 B.n1012 B.n1011 585
R1317 B.n1011 B.n1010 585
R1318 B.n39 B.n38 585
R1319 B.n1009 B.n39 585
R1320 B.n1007 B.n1006 585
R1321 B.n1008 B.n1007 585
R1322 B.n1005 B.n44 585
R1323 B.n44 B.n43 585
R1324 B.n1004 B.n1003 585
R1325 B.n1003 B.n1002 585
R1326 B.n46 B.n45 585
R1327 B.n1001 B.n46 585
R1328 B.n999 B.n998 585
R1329 B.n1000 B.n999 585
R1330 B.n997 B.n51 585
R1331 B.n51 B.n50 585
R1332 B.n996 B.n995 585
R1333 B.n995 B.n994 585
R1334 B.n53 B.n52 585
R1335 B.n993 B.n53 585
R1336 B.n991 B.n990 585
R1337 B.n992 B.n991 585
R1338 B.n989 B.n57 585
R1339 B.n60 B.n57 585
R1340 B.n988 B.n987 585
R1341 B.n987 B.n986 585
R1342 B.n59 B.n58 585
R1343 B.n985 B.n59 585
R1344 B.n983 B.n982 585
R1345 B.n984 B.n983 585
R1346 B.n981 B.n65 585
R1347 B.n65 B.n64 585
R1348 B.n980 B.n979 585
R1349 B.n979 B.n978 585
R1350 B.n67 B.n66 585
R1351 B.n977 B.n67 585
R1352 B.n975 B.n974 585
R1353 B.n976 B.n975 585
R1354 B.n973 B.n72 585
R1355 B.n72 B.n71 585
R1356 B.n972 B.n971 585
R1357 B.n971 B.n970 585
R1358 B.n74 B.n73 585
R1359 B.n969 B.n74 585
R1360 B.n967 B.n966 585
R1361 B.n968 B.n967 585
R1362 B.n965 B.n78 585
R1363 B.n81 B.n78 585
R1364 B.n964 B.n963 585
R1365 B.n963 B.n962 585
R1366 B.n80 B.n79 585
R1367 B.n961 B.n80 585
R1368 B.n959 B.n958 585
R1369 B.n960 B.n959 585
R1370 B.n957 B.n86 585
R1371 B.n86 B.n85 585
R1372 B.n956 B.n955 585
R1373 B.n955 B.n954 585
R1374 B.n88 B.n87 585
R1375 B.n953 B.n88 585
R1376 B.n951 B.n950 585
R1377 B.n952 B.n951 585
R1378 B.n949 B.n93 585
R1379 B.n93 B.n92 585
R1380 B.n948 B.n947 585
R1381 B.n947 B.n946 585
R1382 B.n95 B.n94 585
R1383 B.n945 B.n95 585
R1384 B.n943 B.n942 585
R1385 B.n944 B.n943 585
R1386 B.n941 B.n100 585
R1387 B.n100 B.n99 585
R1388 B.n940 B.n939 585
R1389 B.n939 B.n938 585
R1390 B.n102 B.n101 585
R1391 B.n937 B.n102 585
R1392 B.n935 B.n934 585
R1393 B.n936 B.n935 585
R1394 B.n933 B.n107 585
R1395 B.n107 B.n106 585
R1396 B.n932 B.n931 585
R1397 B.n931 B.n930 585
R1398 B.n109 B.n108 585
R1399 B.n929 B.n109 585
R1400 B.n927 B.n926 585
R1401 B.n928 B.n927 585
R1402 B.n925 B.n114 585
R1403 B.n114 B.n113 585
R1404 B.n924 B.n923 585
R1405 B.n923 B.n922 585
R1406 B.n116 B.n115 585
R1407 B.n921 B.n116 585
R1408 B.n919 B.n918 585
R1409 B.n920 B.n919 585
R1410 B.n917 B.n121 585
R1411 B.n121 B.n120 585
R1412 B.n1052 B.n1051 585
R1413 B.n1051 B.n1050 585
R1414 B.n623 B.n435 449.257
R1415 B.n915 B.n121 449.257
R1416 B.n479 B.n433 449.257
R1417 B.n912 B.n160 449.257
R1418 B.n476 B.t21 300.83
R1419 B.n161 B.t10 300.83
R1420 B.n474 B.t15 300.83
R1421 B.n163 B.t17 300.83
R1422 B.n476 B.t19 265.861
R1423 B.n474 B.t12 265.861
R1424 B.n163 B.t16 265.861
R1425 B.n161 B.t8 265.861
R1426 B.n913 B.n158 256.663
R1427 B.n913 B.n157 256.663
R1428 B.n913 B.n156 256.663
R1429 B.n913 B.n155 256.663
R1430 B.n913 B.n154 256.663
R1431 B.n913 B.n153 256.663
R1432 B.n913 B.n152 256.663
R1433 B.n913 B.n151 256.663
R1434 B.n913 B.n150 256.663
R1435 B.n913 B.n149 256.663
R1436 B.n913 B.n148 256.663
R1437 B.n913 B.n147 256.663
R1438 B.n913 B.n146 256.663
R1439 B.n913 B.n145 256.663
R1440 B.n913 B.n144 256.663
R1441 B.n913 B.n143 256.663
R1442 B.n913 B.n142 256.663
R1443 B.n913 B.n141 256.663
R1444 B.n913 B.n140 256.663
R1445 B.n913 B.n139 256.663
R1446 B.n913 B.n138 256.663
R1447 B.n913 B.n137 256.663
R1448 B.n913 B.n136 256.663
R1449 B.n913 B.n135 256.663
R1450 B.n913 B.n134 256.663
R1451 B.n913 B.n133 256.663
R1452 B.n913 B.n132 256.663
R1453 B.n913 B.n131 256.663
R1454 B.n913 B.n130 256.663
R1455 B.n913 B.n129 256.663
R1456 B.n913 B.n128 256.663
R1457 B.n913 B.n127 256.663
R1458 B.n913 B.n126 256.663
R1459 B.n913 B.n125 256.663
R1460 B.n913 B.n124 256.663
R1461 B.n914 B.n913 256.663
R1462 B.n622 B.n621 256.663
R1463 B.n621 B.n438 256.663
R1464 B.n621 B.n439 256.663
R1465 B.n621 B.n440 256.663
R1466 B.n621 B.n441 256.663
R1467 B.n621 B.n442 256.663
R1468 B.n621 B.n443 256.663
R1469 B.n621 B.n444 256.663
R1470 B.n621 B.n445 256.663
R1471 B.n621 B.n446 256.663
R1472 B.n621 B.n447 256.663
R1473 B.n621 B.n448 256.663
R1474 B.n621 B.n449 256.663
R1475 B.n621 B.n450 256.663
R1476 B.n621 B.n451 256.663
R1477 B.n621 B.n452 256.663
R1478 B.n621 B.n453 256.663
R1479 B.n621 B.n454 256.663
R1480 B.n621 B.n455 256.663
R1481 B.n621 B.n456 256.663
R1482 B.n621 B.n457 256.663
R1483 B.n621 B.n458 256.663
R1484 B.n621 B.n459 256.663
R1485 B.n621 B.n460 256.663
R1486 B.n621 B.n461 256.663
R1487 B.n621 B.n462 256.663
R1488 B.n621 B.n463 256.663
R1489 B.n621 B.n464 256.663
R1490 B.n621 B.n465 256.663
R1491 B.n621 B.n466 256.663
R1492 B.n621 B.n467 256.663
R1493 B.n621 B.n468 256.663
R1494 B.n621 B.n469 256.663
R1495 B.n621 B.n470 256.663
R1496 B.n621 B.n471 256.663
R1497 B.n621 B.n472 256.663
R1498 B.n477 B.t20 223.448
R1499 B.n162 B.t11 223.448
R1500 B.n475 B.t14 223.448
R1501 B.n164 B.t18 223.448
R1502 B.n627 B.n435 163.367
R1503 B.n627 B.n429 163.367
R1504 B.n635 B.n429 163.367
R1505 B.n635 B.n427 163.367
R1506 B.n639 B.n427 163.367
R1507 B.n639 B.n421 163.367
R1508 B.n647 B.n421 163.367
R1509 B.n647 B.n419 163.367
R1510 B.n651 B.n419 163.367
R1511 B.n651 B.n413 163.367
R1512 B.n659 B.n413 163.367
R1513 B.n659 B.n411 163.367
R1514 B.n663 B.n411 163.367
R1515 B.n663 B.n405 163.367
R1516 B.n671 B.n405 163.367
R1517 B.n671 B.n403 163.367
R1518 B.n675 B.n403 163.367
R1519 B.n675 B.n397 163.367
R1520 B.n683 B.n397 163.367
R1521 B.n683 B.n395 163.367
R1522 B.n687 B.n395 163.367
R1523 B.n687 B.n389 163.367
R1524 B.n696 B.n389 163.367
R1525 B.n696 B.n387 163.367
R1526 B.n700 B.n387 163.367
R1527 B.n700 B.n382 163.367
R1528 B.n708 B.n382 163.367
R1529 B.n708 B.n380 163.367
R1530 B.n712 B.n380 163.367
R1531 B.n712 B.n374 163.367
R1532 B.n720 B.n374 163.367
R1533 B.n720 B.n372 163.367
R1534 B.n724 B.n372 163.367
R1535 B.n724 B.n366 163.367
R1536 B.n733 B.n366 163.367
R1537 B.n733 B.n364 163.367
R1538 B.n737 B.n364 163.367
R1539 B.n737 B.n359 163.367
R1540 B.n745 B.n359 163.367
R1541 B.n745 B.n357 163.367
R1542 B.n749 B.n357 163.367
R1543 B.n749 B.n351 163.367
R1544 B.n757 B.n351 163.367
R1545 B.n757 B.n349 163.367
R1546 B.n761 B.n349 163.367
R1547 B.n761 B.n343 163.367
R1548 B.n769 B.n343 163.367
R1549 B.n769 B.n341 163.367
R1550 B.n773 B.n341 163.367
R1551 B.n773 B.n335 163.367
R1552 B.n781 B.n335 163.367
R1553 B.n781 B.n333 163.367
R1554 B.n785 B.n333 163.367
R1555 B.n785 B.n327 163.367
R1556 B.n793 B.n327 163.367
R1557 B.n793 B.n325 163.367
R1558 B.n797 B.n325 163.367
R1559 B.n797 B.n319 163.367
R1560 B.n805 B.n319 163.367
R1561 B.n805 B.n317 163.367
R1562 B.n809 B.n317 163.367
R1563 B.n809 B.n311 163.367
R1564 B.n818 B.n311 163.367
R1565 B.n818 B.n309 163.367
R1566 B.n822 B.n309 163.367
R1567 B.n822 B.n2 163.367
R1568 B.n1051 B.n2 163.367
R1569 B.n1051 B.n3 163.367
R1570 B.n1047 B.n3 163.367
R1571 B.n1047 B.n9 163.367
R1572 B.n1043 B.n9 163.367
R1573 B.n1043 B.n11 163.367
R1574 B.n1039 B.n11 163.367
R1575 B.n1039 B.n16 163.367
R1576 B.n1035 B.n16 163.367
R1577 B.n1035 B.n18 163.367
R1578 B.n1031 B.n18 163.367
R1579 B.n1031 B.n23 163.367
R1580 B.n1027 B.n23 163.367
R1581 B.n1027 B.n25 163.367
R1582 B.n1023 B.n25 163.367
R1583 B.n1023 B.n30 163.367
R1584 B.n1019 B.n30 163.367
R1585 B.n1019 B.n32 163.367
R1586 B.n1015 B.n32 163.367
R1587 B.n1015 B.n37 163.367
R1588 B.n1011 B.n37 163.367
R1589 B.n1011 B.n39 163.367
R1590 B.n1007 B.n39 163.367
R1591 B.n1007 B.n44 163.367
R1592 B.n1003 B.n44 163.367
R1593 B.n1003 B.n46 163.367
R1594 B.n999 B.n46 163.367
R1595 B.n999 B.n51 163.367
R1596 B.n995 B.n51 163.367
R1597 B.n995 B.n53 163.367
R1598 B.n991 B.n53 163.367
R1599 B.n991 B.n57 163.367
R1600 B.n987 B.n57 163.367
R1601 B.n987 B.n59 163.367
R1602 B.n983 B.n59 163.367
R1603 B.n983 B.n65 163.367
R1604 B.n979 B.n65 163.367
R1605 B.n979 B.n67 163.367
R1606 B.n975 B.n67 163.367
R1607 B.n975 B.n72 163.367
R1608 B.n971 B.n72 163.367
R1609 B.n971 B.n74 163.367
R1610 B.n967 B.n74 163.367
R1611 B.n967 B.n78 163.367
R1612 B.n963 B.n78 163.367
R1613 B.n963 B.n80 163.367
R1614 B.n959 B.n80 163.367
R1615 B.n959 B.n86 163.367
R1616 B.n955 B.n86 163.367
R1617 B.n955 B.n88 163.367
R1618 B.n951 B.n88 163.367
R1619 B.n951 B.n93 163.367
R1620 B.n947 B.n93 163.367
R1621 B.n947 B.n95 163.367
R1622 B.n943 B.n95 163.367
R1623 B.n943 B.n100 163.367
R1624 B.n939 B.n100 163.367
R1625 B.n939 B.n102 163.367
R1626 B.n935 B.n102 163.367
R1627 B.n935 B.n107 163.367
R1628 B.n931 B.n107 163.367
R1629 B.n931 B.n109 163.367
R1630 B.n927 B.n109 163.367
R1631 B.n927 B.n114 163.367
R1632 B.n923 B.n114 163.367
R1633 B.n923 B.n116 163.367
R1634 B.n919 B.n116 163.367
R1635 B.n919 B.n121 163.367
R1636 B.n620 B.n437 163.367
R1637 B.n620 B.n473 163.367
R1638 B.n616 B.n615 163.367
R1639 B.n612 B.n611 163.367
R1640 B.n608 B.n607 163.367
R1641 B.n604 B.n603 163.367
R1642 B.n600 B.n599 163.367
R1643 B.n596 B.n595 163.367
R1644 B.n592 B.n591 163.367
R1645 B.n588 B.n587 163.367
R1646 B.n584 B.n583 163.367
R1647 B.n580 B.n579 163.367
R1648 B.n576 B.n575 163.367
R1649 B.n572 B.n571 163.367
R1650 B.n568 B.n567 163.367
R1651 B.n564 B.n563 163.367
R1652 B.n559 B.n558 163.367
R1653 B.n555 B.n554 163.367
R1654 B.n551 B.n550 163.367
R1655 B.n547 B.n546 163.367
R1656 B.n543 B.n542 163.367
R1657 B.n539 B.n538 163.367
R1658 B.n535 B.n534 163.367
R1659 B.n531 B.n530 163.367
R1660 B.n527 B.n526 163.367
R1661 B.n523 B.n522 163.367
R1662 B.n519 B.n518 163.367
R1663 B.n515 B.n514 163.367
R1664 B.n511 B.n510 163.367
R1665 B.n507 B.n506 163.367
R1666 B.n503 B.n502 163.367
R1667 B.n499 B.n498 163.367
R1668 B.n495 B.n494 163.367
R1669 B.n491 B.n490 163.367
R1670 B.n487 B.n486 163.367
R1671 B.n483 B.n482 163.367
R1672 B.n629 B.n433 163.367
R1673 B.n629 B.n431 163.367
R1674 B.n633 B.n431 163.367
R1675 B.n633 B.n425 163.367
R1676 B.n641 B.n425 163.367
R1677 B.n641 B.n423 163.367
R1678 B.n645 B.n423 163.367
R1679 B.n645 B.n417 163.367
R1680 B.n653 B.n417 163.367
R1681 B.n653 B.n415 163.367
R1682 B.n657 B.n415 163.367
R1683 B.n657 B.n409 163.367
R1684 B.n665 B.n409 163.367
R1685 B.n665 B.n407 163.367
R1686 B.n669 B.n407 163.367
R1687 B.n669 B.n401 163.367
R1688 B.n677 B.n401 163.367
R1689 B.n677 B.n399 163.367
R1690 B.n681 B.n399 163.367
R1691 B.n681 B.n393 163.367
R1692 B.n689 B.n393 163.367
R1693 B.n689 B.n391 163.367
R1694 B.n693 B.n391 163.367
R1695 B.n693 B.n386 163.367
R1696 B.n702 B.n386 163.367
R1697 B.n702 B.n384 163.367
R1698 B.n706 B.n384 163.367
R1699 B.n706 B.n378 163.367
R1700 B.n714 B.n378 163.367
R1701 B.n714 B.n376 163.367
R1702 B.n718 B.n376 163.367
R1703 B.n718 B.n370 163.367
R1704 B.n726 B.n370 163.367
R1705 B.n726 B.n368 163.367
R1706 B.n730 B.n368 163.367
R1707 B.n730 B.n363 163.367
R1708 B.n739 B.n363 163.367
R1709 B.n739 B.n361 163.367
R1710 B.n743 B.n361 163.367
R1711 B.n743 B.n355 163.367
R1712 B.n751 B.n355 163.367
R1713 B.n751 B.n353 163.367
R1714 B.n755 B.n353 163.367
R1715 B.n755 B.n347 163.367
R1716 B.n763 B.n347 163.367
R1717 B.n763 B.n345 163.367
R1718 B.n767 B.n345 163.367
R1719 B.n767 B.n339 163.367
R1720 B.n775 B.n339 163.367
R1721 B.n775 B.n337 163.367
R1722 B.n779 B.n337 163.367
R1723 B.n779 B.n331 163.367
R1724 B.n787 B.n331 163.367
R1725 B.n787 B.n329 163.367
R1726 B.n791 B.n329 163.367
R1727 B.n791 B.n323 163.367
R1728 B.n799 B.n323 163.367
R1729 B.n799 B.n321 163.367
R1730 B.n803 B.n321 163.367
R1731 B.n803 B.n315 163.367
R1732 B.n811 B.n315 163.367
R1733 B.n811 B.n313 163.367
R1734 B.n816 B.n313 163.367
R1735 B.n816 B.n307 163.367
R1736 B.n824 B.n307 163.367
R1737 B.n825 B.n824 163.367
R1738 B.n825 B.n5 163.367
R1739 B.n6 B.n5 163.367
R1740 B.n7 B.n6 163.367
R1741 B.n830 B.n7 163.367
R1742 B.n830 B.n12 163.367
R1743 B.n13 B.n12 163.367
R1744 B.n14 B.n13 163.367
R1745 B.n835 B.n14 163.367
R1746 B.n835 B.n19 163.367
R1747 B.n20 B.n19 163.367
R1748 B.n21 B.n20 163.367
R1749 B.n840 B.n21 163.367
R1750 B.n840 B.n26 163.367
R1751 B.n27 B.n26 163.367
R1752 B.n28 B.n27 163.367
R1753 B.n845 B.n28 163.367
R1754 B.n845 B.n33 163.367
R1755 B.n34 B.n33 163.367
R1756 B.n35 B.n34 163.367
R1757 B.n850 B.n35 163.367
R1758 B.n850 B.n40 163.367
R1759 B.n41 B.n40 163.367
R1760 B.n42 B.n41 163.367
R1761 B.n855 B.n42 163.367
R1762 B.n855 B.n47 163.367
R1763 B.n48 B.n47 163.367
R1764 B.n49 B.n48 163.367
R1765 B.n860 B.n49 163.367
R1766 B.n860 B.n54 163.367
R1767 B.n55 B.n54 163.367
R1768 B.n56 B.n55 163.367
R1769 B.n865 B.n56 163.367
R1770 B.n865 B.n61 163.367
R1771 B.n62 B.n61 163.367
R1772 B.n63 B.n62 163.367
R1773 B.n870 B.n63 163.367
R1774 B.n870 B.n68 163.367
R1775 B.n69 B.n68 163.367
R1776 B.n70 B.n69 163.367
R1777 B.n875 B.n70 163.367
R1778 B.n875 B.n75 163.367
R1779 B.n76 B.n75 163.367
R1780 B.n77 B.n76 163.367
R1781 B.n880 B.n77 163.367
R1782 B.n880 B.n82 163.367
R1783 B.n83 B.n82 163.367
R1784 B.n84 B.n83 163.367
R1785 B.n885 B.n84 163.367
R1786 B.n885 B.n89 163.367
R1787 B.n90 B.n89 163.367
R1788 B.n91 B.n90 163.367
R1789 B.n890 B.n91 163.367
R1790 B.n890 B.n96 163.367
R1791 B.n97 B.n96 163.367
R1792 B.n98 B.n97 163.367
R1793 B.n895 B.n98 163.367
R1794 B.n895 B.n103 163.367
R1795 B.n104 B.n103 163.367
R1796 B.n105 B.n104 163.367
R1797 B.n900 B.n105 163.367
R1798 B.n900 B.n110 163.367
R1799 B.n111 B.n110 163.367
R1800 B.n112 B.n111 163.367
R1801 B.n905 B.n112 163.367
R1802 B.n905 B.n117 163.367
R1803 B.n118 B.n117 163.367
R1804 B.n119 B.n118 163.367
R1805 B.n160 B.n119 163.367
R1806 B.n166 B.n123 163.367
R1807 B.n170 B.n169 163.367
R1808 B.n174 B.n173 163.367
R1809 B.n178 B.n177 163.367
R1810 B.n182 B.n181 163.367
R1811 B.n186 B.n185 163.367
R1812 B.n190 B.n189 163.367
R1813 B.n194 B.n193 163.367
R1814 B.n198 B.n197 163.367
R1815 B.n202 B.n201 163.367
R1816 B.n206 B.n205 163.367
R1817 B.n210 B.n209 163.367
R1818 B.n214 B.n213 163.367
R1819 B.n218 B.n217 163.367
R1820 B.n222 B.n221 163.367
R1821 B.n226 B.n225 163.367
R1822 B.n230 B.n229 163.367
R1823 B.n234 B.n233 163.367
R1824 B.n238 B.n237 163.367
R1825 B.n242 B.n241 163.367
R1826 B.n247 B.n246 163.367
R1827 B.n251 B.n250 163.367
R1828 B.n255 B.n254 163.367
R1829 B.n259 B.n258 163.367
R1830 B.n263 B.n262 163.367
R1831 B.n267 B.n266 163.367
R1832 B.n271 B.n270 163.367
R1833 B.n275 B.n274 163.367
R1834 B.n279 B.n278 163.367
R1835 B.n283 B.n282 163.367
R1836 B.n287 B.n286 163.367
R1837 B.n291 B.n290 163.367
R1838 B.n295 B.n294 163.367
R1839 B.n299 B.n298 163.367
R1840 B.n303 B.n302 163.367
R1841 B.n912 B.n159 163.367
R1842 B.n621 B.n434 86.4149
R1843 B.n913 B.n120 86.4149
R1844 B.n477 B.n476 77.3823
R1845 B.n475 B.n474 77.3823
R1846 B.n164 B.n163 77.3823
R1847 B.n162 B.n161 77.3823
R1848 B.n623 B.n622 71.676
R1849 B.n473 B.n438 71.676
R1850 B.n615 B.n439 71.676
R1851 B.n611 B.n440 71.676
R1852 B.n607 B.n441 71.676
R1853 B.n603 B.n442 71.676
R1854 B.n599 B.n443 71.676
R1855 B.n595 B.n444 71.676
R1856 B.n591 B.n445 71.676
R1857 B.n587 B.n446 71.676
R1858 B.n583 B.n447 71.676
R1859 B.n579 B.n448 71.676
R1860 B.n575 B.n449 71.676
R1861 B.n571 B.n450 71.676
R1862 B.n567 B.n451 71.676
R1863 B.n563 B.n452 71.676
R1864 B.n558 B.n453 71.676
R1865 B.n554 B.n454 71.676
R1866 B.n550 B.n455 71.676
R1867 B.n546 B.n456 71.676
R1868 B.n542 B.n457 71.676
R1869 B.n538 B.n458 71.676
R1870 B.n534 B.n459 71.676
R1871 B.n530 B.n460 71.676
R1872 B.n526 B.n461 71.676
R1873 B.n522 B.n462 71.676
R1874 B.n518 B.n463 71.676
R1875 B.n514 B.n464 71.676
R1876 B.n510 B.n465 71.676
R1877 B.n506 B.n466 71.676
R1878 B.n502 B.n467 71.676
R1879 B.n498 B.n468 71.676
R1880 B.n494 B.n469 71.676
R1881 B.n490 B.n470 71.676
R1882 B.n486 B.n471 71.676
R1883 B.n482 B.n472 71.676
R1884 B.n915 B.n914 71.676
R1885 B.n166 B.n124 71.676
R1886 B.n170 B.n125 71.676
R1887 B.n174 B.n126 71.676
R1888 B.n178 B.n127 71.676
R1889 B.n182 B.n128 71.676
R1890 B.n186 B.n129 71.676
R1891 B.n190 B.n130 71.676
R1892 B.n194 B.n131 71.676
R1893 B.n198 B.n132 71.676
R1894 B.n202 B.n133 71.676
R1895 B.n206 B.n134 71.676
R1896 B.n210 B.n135 71.676
R1897 B.n214 B.n136 71.676
R1898 B.n218 B.n137 71.676
R1899 B.n222 B.n138 71.676
R1900 B.n226 B.n139 71.676
R1901 B.n230 B.n140 71.676
R1902 B.n234 B.n141 71.676
R1903 B.n238 B.n142 71.676
R1904 B.n242 B.n143 71.676
R1905 B.n247 B.n144 71.676
R1906 B.n251 B.n145 71.676
R1907 B.n255 B.n146 71.676
R1908 B.n259 B.n147 71.676
R1909 B.n263 B.n148 71.676
R1910 B.n267 B.n149 71.676
R1911 B.n271 B.n150 71.676
R1912 B.n275 B.n151 71.676
R1913 B.n279 B.n152 71.676
R1914 B.n283 B.n153 71.676
R1915 B.n287 B.n154 71.676
R1916 B.n291 B.n155 71.676
R1917 B.n295 B.n156 71.676
R1918 B.n299 B.n157 71.676
R1919 B.n303 B.n158 71.676
R1920 B.n159 B.n158 71.676
R1921 B.n302 B.n157 71.676
R1922 B.n298 B.n156 71.676
R1923 B.n294 B.n155 71.676
R1924 B.n290 B.n154 71.676
R1925 B.n286 B.n153 71.676
R1926 B.n282 B.n152 71.676
R1927 B.n278 B.n151 71.676
R1928 B.n274 B.n150 71.676
R1929 B.n270 B.n149 71.676
R1930 B.n266 B.n148 71.676
R1931 B.n262 B.n147 71.676
R1932 B.n258 B.n146 71.676
R1933 B.n254 B.n145 71.676
R1934 B.n250 B.n144 71.676
R1935 B.n246 B.n143 71.676
R1936 B.n241 B.n142 71.676
R1937 B.n237 B.n141 71.676
R1938 B.n233 B.n140 71.676
R1939 B.n229 B.n139 71.676
R1940 B.n225 B.n138 71.676
R1941 B.n221 B.n137 71.676
R1942 B.n217 B.n136 71.676
R1943 B.n213 B.n135 71.676
R1944 B.n209 B.n134 71.676
R1945 B.n205 B.n133 71.676
R1946 B.n201 B.n132 71.676
R1947 B.n197 B.n131 71.676
R1948 B.n193 B.n130 71.676
R1949 B.n189 B.n129 71.676
R1950 B.n185 B.n128 71.676
R1951 B.n181 B.n127 71.676
R1952 B.n177 B.n126 71.676
R1953 B.n173 B.n125 71.676
R1954 B.n169 B.n124 71.676
R1955 B.n914 B.n123 71.676
R1956 B.n622 B.n437 71.676
R1957 B.n616 B.n438 71.676
R1958 B.n612 B.n439 71.676
R1959 B.n608 B.n440 71.676
R1960 B.n604 B.n441 71.676
R1961 B.n600 B.n442 71.676
R1962 B.n596 B.n443 71.676
R1963 B.n592 B.n444 71.676
R1964 B.n588 B.n445 71.676
R1965 B.n584 B.n446 71.676
R1966 B.n580 B.n447 71.676
R1967 B.n576 B.n448 71.676
R1968 B.n572 B.n449 71.676
R1969 B.n568 B.n450 71.676
R1970 B.n564 B.n451 71.676
R1971 B.n559 B.n452 71.676
R1972 B.n555 B.n453 71.676
R1973 B.n551 B.n454 71.676
R1974 B.n547 B.n455 71.676
R1975 B.n543 B.n456 71.676
R1976 B.n539 B.n457 71.676
R1977 B.n535 B.n458 71.676
R1978 B.n531 B.n459 71.676
R1979 B.n527 B.n460 71.676
R1980 B.n523 B.n461 71.676
R1981 B.n519 B.n462 71.676
R1982 B.n515 B.n463 71.676
R1983 B.n511 B.n464 71.676
R1984 B.n507 B.n465 71.676
R1985 B.n503 B.n466 71.676
R1986 B.n499 B.n467 71.676
R1987 B.n495 B.n468 71.676
R1988 B.n491 B.n469 71.676
R1989 B.n487 B.n470 71.676
R1990 B.n483 B.n471 71.676
R1991 B.n479 B.n472 71.676
R1992 B.n478 B.n477 59.5399
R1993 B.n561 B.n475 59.5399
R1994 B.n165 B.n164 59.5399
R1995 B.n244 B.n162 59.5399
R1996 B.n628 B.n434 53.9104
R1997 B.n628 B.n430 53.9104
R1998 B.n634 B.n430 53.9104
R1999 B.n634 B.n426 53.9104
R2000 B.n640 B.n426 53.9104
R2001 B.n640 B.n422 53.9104
R2002 B.n646 B.n422 53.9104
R2003 B.n646 B.n418 53.9104
R2004 B.n652 B.n418 53.9104
R2005 B.n658 B.n414 53.9104
R2006 B.n658 B.n410 53.9104
R2007 B.n664 B.n410 53.9104
R2008 B.n664 B.n406 53.9104
R2009 B.n670 B.n406 53.9104
R2010 B.n670 B.n402 53.9104
R2011 B.n676 B.n402 53.9104
R2012 B.n676 B.n398 53.9104
R2013 B.n682 B.n398 53.9104
R2014 B.n682 B.n394 53.9104
R2015 B.n688 B.n394 53.9104
R2016 B.n688 B.n390 53.9104
R2017 B.n695 B.n390 53.9104
R2018 B.n695 B.n694 53.9104
R2019 B.n701 B.n383 53.9104
R2020 B.n707 B.n383 53.9104
R2021 B.n707 B.n379 53.9104
R2022 B.n713 B.n379 53.9104
R2023 B.n713 B.n375 53.9104
R2024 B.n719 B.n375 53.9104
R2025 B.n719 B.n371 53.9104
R2026 B.n725 B.n371 53.9104
R2027 B.n725 B.n367 53.9104
R2028 B.n732 B.n367 53.9104
R2029 B.n732 B.n731 53.9104
R2030 B.n738 B.n360 53.9104
R2031 B.n744 B.n360 53.9104
R2032 B.n744 B.n356 53.9104
R2033 B.n750 B.n356 53.9104
R2034 B.n750 B.n352 53.9104
R2035 B.n756 B.n352 53.9104
R2036 B.n756 B.n348 53.9104
R2037 B.n762 B.n348 53.9104
R2038 B.n762 B.n344 53.9104
R2039 B.n768 B.n344 53.9104
R2040 B.n774 B.n340 53.9104
R2041 B.n774 B.n336 53.9104
R2042 B.n780 B.n336 53.9104
R2043 B.n780 B.n332 53.9104
R2044 B.n786 B.n332 53.9104
R2045 B.n786 B.n328 53.9104
R2046 B.n792 B.n328 53.9104
R2047 B.n792 B.n324 53.9104
R2048 B.n798 B.n324 53.9104
R2049 B.n798 B.n320 53.9104
R2050 B.n804 B.n320 53.9104
R2051 B.n810 B.n316 53.9104
R2052 B.n810 B.n312 53.9104
R2053 B.n817 B.n312 53.9104
R2054 B.n817 B.n308 53.9104
R2055 B.n823 B.n308 53.9104
R2056 B.n823 B.n4 53.9104
R2057 B.n1050 B.n4 53.9104
R2058 B.n1050 B.n1049 53.9104
R2059 B.n1049 B.n1048 53.9104
R2060 B.n1048 B.n8 53.9104
R2061 B.n1042 B.n8 53.9104
R2062 B.n1042 B.n1041 53.9104
R2063 B.n1041 B.n1040 53.9104
R2064 B.n1040 B.n15 53.9104
R2065 B.n1034 B.n1033 53.9104
R2066 B.n1033 B.n1032 53.9104
R2067 B.n1032 B.n22 53.9104
R2068 B.n1026 B.n22 53.9104
R2069 B.n1026 B.n1025 53.9104
R2070 B.n1025 B.n1024 53.9104
R2071 B.n1024 B.n29 53.9104
R2072 B.n1018 B.n29 53.9104
R2073 B.n1018 B.n1017 53.9104
R2074 B.n1017 B.n1016 53.9104
R2075 B.n1016 B.n36 53.9104
R2076 B.n1010 B.n1009 53.9104
R2077 B.n1009 B.n1008 53.9104
R2078 B.n1008 B.n43 53.9104
R2079 B.n1002 B.n43 53.9104
R2080 B.n1002 B.n1001 53.9104
R2081 B.n1001 B.n1000 53.9104
R2082 B.n1000 B.n50 53.9104
R2083 B.n994 B.n50 53.9104
R2084 B.n994 B.n993 53.9104
R2085 B.n993 B.n992 53.9104
R2086 B.n986 B.n60 53.9104
R2087 B.n986 B.n985 53.9104
R2088 B.n985 B.n984 53.9104
R2089 B.n984 B.n64 53.9104
R2090 B.n978 B.n64 53.9104
R2091 B.n978 B.n977 53.9104
R2092 B.n977 B.n976 53.9104
R2093 B.n976 B.n71 53.9104
R2094 B.n970 B.n71 53.9104
R2095 B.n970 B.n969 53.9104
R2096 B.n969 B.n968 53.9104
R2097 B.n962 B.n81 53.9104
R2098 B.n962 B.n961 53.9104
R2099 B.n961 B.n960 53.9104
R2100 B.n960 B.n85 53.9104
R2101 B.n954 B.n85 53.9104
R2102 B.n954 B.n953 53.9104
R2103 B.n953 B.n952 53.9104
R2104 B.n952 B.n92 53.9104
R2105 B.n946 B.n92 53.9104
R2106 B.n946 B.n945 53.9104
R2107 B.n945 B.n944 53.9104
R2108 B.n944 B.n99 53.9104
R2109 B.n938 B.n99 53.9104
R2110 B.n938 B.n937 53.9104
R2111 B.n936 B.n106 53.9104
R2112 B.n930 B.n106 53.9104
R2113 B.n930 B.n929 53.9104
R2114 B.n929 B.n928 53.9104
R2115 B.n928 B.n113 53.9104
R2116 B.n922 B.n113 53.9104
R2117 B.n922 B.n921 53.9104
R2118 B.n921 B.n920 53.9104
R2119 B.n920 B.n120 53.9104
R2120 B.n738 B.t4 50.7392
R2121 B.n992 B.t1 50.7392
R2122 B.n768 B.t0 42.8113
R2123 B.n1010 B.t7 42.8113
R2124 B.n701 B.t3 36.469
R2125 B.n968 B.t2 36.469
R2126 B.t13 B.n414 33.2978
R2127 B.n937 B.t9 33.2978
R2128 B.n917 B.n916 29.1907
R2129 B.n480 B.n432 29.1907
R2130 B.n625 B.n624 29.1907
R2131 B.n911 B.n910 29.1907
R2132 B.n804 B.t5 28.541
R2133 B.n1034 B.t6 28.541
R2134 B.t5 B.n316 25.3699
R2135 B.t6 B.n15 25.3699
R2136 B.n652 B.t13 20.6131
R2137 B.t9 B.n936 20.6131
R2138 B B.n1052 18.0485
R2139 B.n694 B.t3 17.4419
R2140 B.n81 B.t2 17.4419
R2141 B.t0 B.n340 11.0996
R2142 B.t7 B.n36 11.0996
R2143 B.n916 B.n122 10.6151
R2144 B.n167 B.n122 10.6151
R2145 B.n168 B.n167 10.6151
R2146 B.n171 B.n168 10.6151
R2147 B.n172 B.n171 10.6151
R2148 B.n175 B.n172 10.6151
R2149 B.n176 B.n175 10.6151
R2150 B.n179 B.n176 10.6151
R2151 B.n180 B.n179 10.6151
R2152 B.n183 B.n180 10.6151
R2153 B.n184 B.n183 10.6151
R2154 B.n187 B.n184 10.6151
R2155 B.n188 B.n187 10.6151
R2156 B.n191 B.n188 10.6151
R2157 B.n192 B.n191 10.6151
R2158 B.n195 B.n192 10.6151
R2159 B.n196 B.n195 10.6151
R2160 B.n199 B.n196 10.6151
R2161 B.n200 B.n199 10.6151
R2162 B.n203 B.n200 10.6151
R2163 B.n204 B.n203 10.6151
R2164 B.n207 B.n204 10.6151
R2165 B.n208 B.n207 10.6151
R2166 B.n211 B.n208 10.6151
R2167 B.n212 B.n211 10.6151
R2168 B.n215 B.n212 10.6151
R2169 B.n216 B.n215 10.6151
R2170 B.n219 B.n216 10.6151
R2171 B.n220 B.n219 10.6151
R2172 B.n223 B.n220 10.6151
R2173 B.n224 B.n223 10.6151
R2174 B.n228 B.n227 10.6151
R2175 B.n231 B.n228 10.6151
R2176 B.n232 B.n231 10.6151
R2177 B.n235 B.n232 10.6151
R2178 B.n236 B.n235 10.6151
R2179 B.n239 B.n236 10.6151
R2180 B.n240 B.n239 10.6151
R2181 B.n243 B.n240 10.6151
R2182 B.n248 B.n245 10.6151
R2183 B.n249 B.n248 10.6151
R2184 B.n252 B.n249 10.6151
R2185 B.n253 B.n252 10.6151
R2186 B.n256 B.n253 10.6151
R2187 B.n257 B.n256 10.6151
R2188 B.n260 B.n257 10.6151
R2189 B.n261 B.n260 10.6151
R2190 B.n264 B.n261 10.6151
R2191 B.n265 B.n264 10.6151
R2192 B.n268 B.n265 10.6151
R2193 B.n269 B.n268 10.6151
R2194 B.n272 B.n269 10.6151
R2195 B.n273 B.n272 10.6151
R2196 B.n276 B.n273 10.6151
R2197 B.n277 B.n276 10.6151
R2198 B.n280 B.n277 10.6151
R2199 B.n281 B.n280 10.6151
R2200 B.n284 B.n281 10.6151
R2201 B.n285 B.n284 10.6151
R2202 B.n288 B.n285 10.6151
R2203 B.n289 B.n288 10.6151
R2204 B.n292 B.n289 10.6151
R2205 B.n293 B.n292 10.6151
R2206 B.n296 B.n293 10.6151
R2207 B.n297 B.n296 10.6151
R2208 B.n300 B.n297 10.6151
R2209 B.n301 B.n300 10.6151
R2210 B.n304 B.n301 10.6151
R2211 B.n305 B.n304 10.6151
R2212 B.n911 B.n305 10.6151
R2213 B.n630 B.n432 10.6151
R2214 B.n631 B.n630 10.6151
R2215 B.n632 B.n631 10.6151
R2216 B.n632 B.n424 10.6151
R2217 B.n642 B.n424 10.6151
R2218 B.n643 B.n642 10.6151
R2219 B.n644 B.n643 10.6151
R2220 B.n644 B.n416 10.6151
R2221 B.n654 B.n416 10.6151
R2222 B.n655 B.n654 10.6151
R2223 B.n656 B.n655 10.6151
R2224 B.n656 B.n408 10.6151
R2225 B.n666 B.n408 10.6151
R2226 B.n667 B.n666 10.6151
R2227 B.n668 B.n667 10.6151
R2228 B.n668 B.n400 10.6151
R2229 B.n678 B.n400 10.6151
R2230 B.n679 B.n678 10.6151
R2231 B.n680 B.n679 10.6151
R2232 B.n680 B.n392 10.6151
R2233 B.n690 B.n392 10.6151
R2234 B.n691 B.n690 10.6151
R2235 B.n692 B.n691 10.6151
R2236 B.n692 B.n385 10.6151
R2237 B.n703 B.n385 10.6151
R2238 B.n704 B.n703 10.6151
R2239 B.n705 B.n704 10.6151
R2240 B.n705 B.n377 10.6151
R2241 B.n715 B.n377 10.6151
R2242 B.n716 B.n715 10.6151
R2243 B.n717 B.n716 10.6151
R2244 B.n717 B.n369 10.6151
R2245 B.n727 B.n369 10.6151
R2246 B.n728 B.n727 10.6151
R2247 B.n729 B.n728 10.6151
R2248 B.n729 B.n362 10.6151
R2249 B.n740 B.n362 10.6151
R2250 B.n741 B.n740 10.6151
R2251 B.n742 B.n741 10.6151
R2252 B.n742 B.n354 10.6151
R2253 B.n752 B.n354 10.6151
R2254 B.n753 B.n752 10.6151
R2255 B.n754 B.n753 10.6151
R2256 B.n754 B.n346 10.6151
R2257 B.n764 B.n346 10.6151
R2258 B.n765 B.n764 10.6151
R2259 B.n766 B.n765 10.6151
R2260 B.n766 B.n338 10.6151
R2261 B.n776 B.n338 10.6151
R2262 B.n777 B.n776 10.6151
R2263 B.n778 B.n777 10.6151
R2264 B.n778 B.n330 10.6151
R2265 B.n788 B.n330 10.6151
R2266 B.n789 B.n788 10.6151
R2267 B.n790 B.n789 10.6151
R2268 B.n790 B.n322 10.6151
R2269 B.n800 B.n322 10.6151
R2270 B.n801 B.n800 10.6151
R2271 B.n802 B.n801 10.6151
R2272 B.n802 B.n314 10.6151
R2273 B.n812 B.n314 10.6151
R2274 B.n813 B.n812 10.6151
R2275 B.n815 B.n813 10.6151
R2276 B.n815 B.n814 10.6151
R2277 B.n814 B.n306 10.6151
R2278 B.n826 B.n306 10.6151
R2279 B.n827 B.n826 10.6151
R2280 B.n828 B.n827 10.6151
R2281 B.n829 B.n828 10.6151
R2282 B.n831 B.n829 10.6151
R2283 B.n832 B.n831 10.6151
R2284 B.n833 B.n832 10.6151
R2285 B.n834 B.n833 10.6151
R2286 B.n836 B.n834 10.6151
R2287 B.n837 B.n836 10.6151
R2288 B.n838 B.n837 10.6151
R2289 B.n839 B.n838 10.6151
R2290 B.n841 B.n839 10.6151
R2291 B.n842 B.n841 10.6151
R2292 B.n843 B.n842 10.6151
R2293 B.n844 B.n843 10.6151
R2294 B.n846 B.n844 10.6151
R2295 B.n847 B.n846 10.6151
R2296 B.n848 B.n847 10.6151
R2297 B.n849 B.n848 10.6151
R2298 B.n851 B.n849 10.6151
R2299 B.n852 B.n851 10.6151
R2300 B.n853 B.n852 10.6151
R2301 B.n854 B.n853 10.6151
R2302 B.n856 B.n854 10.6151
R2303 B.n857 B.n856 10.6151
R2304 B.n858 B.n857 10.6151
R2305 B.n859 B.n858 10.6151
R2306 B.n861 B.n859 10.6151
R2307 B.n862 B.n861 10.6151
R2308 B.n863 B.n862 10.6151
R2309 B.n864 B.n863 10.6151
R2310 B.n866 B.n864 10.6151
R2311 B.n867 B.n866 10.6151
R2312 B.n868 B.n867 10.6151
R2313 B.n869 B.n868 10.6151
R2314 B.n871 B.n869 10.6151
R2315 B.n872 B.n871 10.6151
R2316 B.n873 B.n872 10.6151
R2317 B.n874 B.n873 10.6151
R2318 B.n876 B.n874 10.6151
R2319 B.n877 B.n876 10.6151
R2320 B.n878 B.n877 10.6151
R2321 B.n879 B.n878 10.6151
R2322 B.n881 B.n879 10.6151
R2323 B.n882 B.n881 10.6151
R2324 B.n883 B.n882 10.6151
R2325 B.n884 B.n883 10.6151
R2326 B.n886 B.n884 10.6151
R2327 B.n887 B.n886 10.6151
R2328 B.n888 B.n887 10.6151
R2329 B.n889 B.n888 10.6151
R2330 B.n891 B.n889 10.6151
R2331 B.n892 B.n891 10.6151
R2332 B.n893 B.n892 10.6151
R2333 B.n894 B.n893 10.6151
R2334 B.n896 B.n894 10.6151
R2335 B.n897 B.n896 10.6151
R2336 B.n898 B.n897 10.6151
R2337 B.n899 B.n898 10.6151
R2338 B.n901 B.n899 10.6151
R2339 B.n902 B.n901 10.6151
R2340 B.n903 B.n902 10.6151
R2341 B.n904 B.n903 10.6151
R2342 B.n906 B.n904 10.6151
R2343 B.n907 B.n906 10.6151
R2344 B.n908 B.n907 10.6151
R2345 B.n909 B.n908 10.6151
R2346 B.n910 B.n909 10.6151
R2347 B.n624 B.n436 10.6151
R2348 B.n619 B.n436 10.6151
R2349 B.n619 B.n618 10.6151
R2350 B.n618 B.n617 10.6151
R2351 B.n617 B.n614 10.6151
R2352 B.n614 B.n613 10.6151
R2353 B.n613 B.n610 10.6151
R2354 B.n610 B.n609 10.6151
R2355 B.n609 B.n606 10.6151
R2356 B.n606 B.n605 10.6151
R2357 B.n605 B.n602 10.6151
R2358 B.n602 B.n601 10.6151
R2359 B.n601 B.n598 10.6151
R2360 B.n598 B.n597 10.6151
R2361 B.n597 B.n594 10.6151
R2362 B.n594 B.n593 10.6151
R2363 B.n593 B.n590 10.6151
R2364 B.n590 B.n589 10.6151
R2365 B.n589 B.n586 10.6151
R2366 B.n586 B.n585 10.6151
R2367 B.n585 B.n582 10.6151
R2368 B.n582 B.n581 10.6151
R2369 B.n581 B.n578 10.6151
R2370 B.n578 B.n577 10.6151
R2371 B.n577 B.n574 10.6151
R2372 B.n574 B.n573 10.6151
R2373 B.n573 B.n570 10.6151
R2374 B.n570 B.n569 10.6151
R2375 B.n569 B.n566 10.6151
R2376 B.n566 B.n565 10.6151
R2377 B.n565 B.n562 10.6151
R2378 B.n560 B.n557 10.6151
R2379 B.n557 B.n556 10.6151
R2380 B.n556 B.n553 10.6151
R2381 B.n553 B.n552 10.6151
R2382 B.n552 B.n549 10.6151
R2383 B.n549 B.n548 10.6151
R2384 B.n548 B.n545 10.6151
R2385 B.n545 B.n544 10.6151
R2386 B.n541 B.n540 10.6151
R2387 B.n540 B.n537 10.6151
R2388 B.n537 B.n536 10.6151
R2389 B.n536 B.n533 10.6151
R2390 B.n533 B.n532 10.6151
R2391 B.n532 B.n529 10.6151
R2392 B.n529 B.n528 10.6151
R2393 B.n528 B.n525 10.6151
R2394 B.n525 B.n524 10.6151
R2395 B.n524 B.n521 10.6151
R2396 B.n521 B.n520 10.6151
R2397 B.n520 B.n517 10.6151
R2398 B.n517 B.n516 10.6151
R2399 B.n516 B.n513 10.6151
R2400 B.n513 B.n512 10.6151
R2401 B.n512 B.n509 10.6151
R2402 B.n509 B.n508 10.6151
R2403 B.n508 B.n505 10.6151
R2404 B.n505 B.n504 10.6151
R2405 B.n504 B.n501 10.6151
R2406 B.n501 B.n500 10.6151
R2407 B.n500 B.n497 10.6151
R2408 B.n497 B.n496 10.6151
R2409 B.n496 B.n493 10.6151
R2410 B.n493 B.n492 10.6151
R2411 B.n492 B.n489 10.6151
R2412 B.n489 B.n488 10.6151
R2413 B.n488 B.n485 10.6151
R2414 B.n485 B.n484 10.6151
R2415 B.n484 B.n481 10.6151
R2416 B.n481 B.n480 10.6151
R2417 B.n626 B.n625 10.6151
R2418 B.n626 B.n428 10.6151
R2419 B.n636 B.n428 10.6151
R2420 B.n637 B.n636 10.6151
R2421 B.n638 B.n637 10.6151
R2422 B.n638 B.n420 10.6151
R2423 B.n648 B.n420 10.6151
R2424 B.n649 B.n648 10.6151
R2425 B.n650 B.n649 10.6151
R2426 B.n650 B.n412 10.6151
R2427 B.n660 B.n412 10.6151
R2428 B.n661 B.n660 10.6151
R2429 B.n662 B.n661 10.6151
R2430 B.n662 B.n404 10.6151
R2431 B.n672 B.n404 10.6151
R2432 B.n673 B.n672 10.6151
R2433 B.n674 B.n673 10.6151
R2434 B.n674 B.n396 10.6151
R2435 B.n684 B.n396 10.6151
R2436 B.n685 B.n684 10.6151
R2437 B.n686 B.n685 10.6151
R2438 B.n686 B.n388 10.6151
R2439 B.n697 B.n388 10.6151
R2440 B.n698 B.n697 10.6151
R2441 B.n699 B.n698 10.6151
R2442 B.n699 B.n381 10.6151
R2443 B.n709 B.n381 10.6151
R2444 B.n710 B.n709 10.6151
R2445 B.n711 B.n710 10.6151
R2446 B.n711 B.n373 10.6151
R2447 B.n721 B.n373 10.6151
R2448 B.n722 B.n721 10.6151
R2449 B.n723 B.n722 10.6151
R2450 B.n723 B.n365 10.6151
R2451 B.n734 B.n365 10.6151
R2452 B.n735 B.n734 10.6151
R2453 B.n736 B.n735 10.6151
R2454 B.n736 B.n358 10.6151
R2455 B.n746 B.n358 10.6151
R2456 B.n747 B.n746 10.6151
R2457 B.n748 B.n747 10.6151
R2458 B.n748 B.n350 10.6151
R2459 B.n758 B.n350 10.6151
R2460 B.n759 B.n758 10.6151
R2461 B.n760 B.n759 10.6151
R2462 B.n760 B.n342 10.6151
R2463 B.n770 B.n342 10.6151
R2464 B.n771 B.n770 10.6151
R2465 B.n772 B.n771 10.6151
R2466 B.n772 B.n334 10.6151
R2467 B.n782 B.n334 10.6151
R2468 B.n783 B.n782 10.6151
R2469 B.n784 B.n783 10.6151
R2470 B.n784 B.n326 10.6151
R2471 B.n794 B.n326 10.6151
R2472 B.n795 B.n794 10.6151
R2473 B.n796 B.n795 10.6151
R2474 B.n796 B.n318 10.6151
R2475 B.n806 B.n318 10.6151
R2476 B.n807 B.n806 10.6151
R2477 B.n808 B.n807 10.6151
R2478 B.n808 B.n310 10.6151
R2479 B.n819 B.n310 10.6151
R2480 B.n820 B.n819 10.6151
R2481 B.n821 B.n820 10.6151
R2482 B.n821 B.n0 10.6151
R2483 B.n1046 B.n1 10.6151
R2484 B.n1046 B.n1045 10.6151
R2485 B.n1045 B.n1044 10.6151
R2486 B.n1044 B.n10 10.6151
R2487 B.n1038 B.n10 10.6151
R2488 B.n1038 B.n1037 10.6151
R2489 B.n1037 B.n1036 10.6151
R2490 B.n1036 B.n17 10.6151
R2491 B.n1030 B.n17 10.6151
R2492 B.n1030 B.n1029 10.6151
R2493 B.n1029 B.n1028 10.6151
R2494 B.n1028 B.n24 10.6151
R2495 B.n1022 B.n24 10.6151
R2496 B.n1022 B.n1021 10.6151
R2497 B.n1021 B.n1020 10.6151
R2498 B.n1020 B.n31 10.6151
R2499 B.n1014 B.n31 10.6151
R2500 B.n1014 B.n1013 10.6151
R2501 B.n1013 B.n1012 10.6151
R2502 B.n1012 B.n38 10.6151
R2503 B.n1006 B.n38 10.6151
R2504 B.n1006 B.n1005 10.6151
R2505 B.n1005 B.n1004 10.6151
R2506 B.n1004 B.n45 10.6151
R2507 B.n998 B.n45 10.6151
R2508 B.n998 B.n997 10.6151
R2509 B.n997 B.n996 10.6151
R2510 B.n996 B.n52 10.6151
R2511 B.n990 B.n52 10.6151
R2512 B.n990 B.n989 10.6151
R2513 B.n989 B.n988 10.6151
R2514 B.n988 B.n58 10.6151
R2515 B.n982 B.n58 10.6151
R2516 B.n982 B.n981 10.6151
R2517 B.n981 B.n980 10.6151
R2518 B.n980 B.n66 10.6151
R2519 B.n974 B.n66 10.6151
R2520 B.n974 B.n973 10.6151
R2521 B.n973 B.n972 10.6151
R2522 B.n972 B.n73 10.6151
R2523 B.n966 B.n73 10.6151
R2524 B.n966 B.n965 10.6151
R2525 B.n965 B.n964 10.6151
R2526 B.n964 B.n79 10.6151
R2527 B.n958 B.n79 10.6151
R2528 B.n958 B.n957 10.6151
R2529 B.n957 B.n956 10.6151
R2530 B.n956 B.n87 10.6151
R2531 B.n950 B.n87 10.6151
R2532 B.n950 B.n949 10.6151
R2533 B.n949 B.n948 10.6151
R2534 B.n948 B.n94 10.6151
R2535 B.n942 B.n94 10.6151
R2536 B.n942 B.n941 10.6151
R2537 B.n941 B.n940 10.6151
R2538 B.n940 B.n101 10.6151
R2539 B.n934 B.n101 10.6151
R2540 B.n934 B.n933 10.6151
R2541 B.n933 B.n932 10.6151
R2542 B.n932 B.n108 10.6151
R2543 B.n926 B.n108 10.6151
R2544 B.n926 B.n925 10.6151
R2545 B.n925 B.n924 10.6151
R2546 B.n924 B.n115 10.6151
R2547 B.n918 B.n115 10.6151
R2548 B.n918 B.n917 10.6151
R2549 B.n227 B.n165 6.5566
R2550 B.n244 B.n243 6.5566
R2551 B.n561 B.n560 6.5566
R2552 B.n544 B.n478 6.5566
R2553 B.n224 B.n165 4.05904
R2554 B.n245 B.n244 4.05904
R2555 B.n562 B.n561 4.05904
R2556 B.n541 B.n478 4.05904
R2557 B.n731 B.t4 3.17167
R2558 B.n60 B.t1 3.17167
R2559 B.n1052 B.n0 2.81026
R2560 B.n1052 B.n1 2.81026
R2561 VN.n67 VN.n35 161.3
R2562 VN.n66 VN.n65 161.3
R2563 VN.n64 VN.n36 161.3
R2564 VN.n63 VN.n62 161.3
R2565 VN.n61 VN.n37 161.3
R2566 VN.n60 VN.n59 161.3
R2567 VN.n58 VN.n38 161.3
R2568 VN.n57 VN.n56 161.3
R2569 VN.n54 VN.n39 161.3
R2570 VN.n53 VN.n52 161.3
R2571 VN.n51 VN.n40 161.3
R2572 VN.n50 VN.n49 161.3
R2573 VN.n48 VN.n41 161.3
R2574 VN.n47 VN.n46 161.3
R2575 VN.n45 VN.n42 161.3
R2576 VN.n32 VN.n0 161.3
R2577 VN.n31 VN.n30 161.3
R2578 VN.n29 VN.n1 161.3
R2579 VN.n28 VN.n27 161.3
R2580 VN.n26 VN.n2 161.3
R2581 VN.n25 VN.n24 161.3
R2582 VN.n23 VN.n3 161.3
R2583 VN.n22 VN.n21 161.3
R2584 VN.n19 VN.n4 161.3
R2585 VN.n18 VN.n17 161.3
R2586 VN.n16 VN.n5 161.3
R2587 VN.n15 VN.n14 161.3
R2588 VN.n13 VN.n6 161.3
R2589 VN.n12 VN.n11 161.3
R2590 VN.n10 VN.n7 161.3
R2591 VN.n9 VN.t5 88.8828
R2592 VN.n44 VN.t6 88.8828
R2593 VN.n34 VN.n33 58.5258
R2594 VN.n69 VN.n68 58.5258
R2595 VN.n8 VN.t4 56.6289
R2596 VN.n20 VN.t3 56.6289
R2597 VN.n33 VN.t0 56.6289
R2598 VN.n43 VN.t7 56.6289
R2599 VN.n55 VN.t1 56.6289
R2600 VN.n68 VN.t2 56.6289
R2601 VN VN.n69 53.5347
R2602 VN.n9 VN.n8 50.8254
R2603 VN.n44 VN.n43 50.8254
R2604 VN.n27 VN.n26 41.5458
R2605 VN.n62 VN.n61 41.5458
R2606 VN.n14 VN.n13 40.577
R2607 VN.n14 VN.n5 40.577
R2608 VN.n49 VN.n48 40.577
R2609 VN.n49 VN.n40 40.577
R2610 VN.n27 VN.n1 39.6083
R2611 VN.n62 VN.n36 39.6083
R2612 VN.n12 VN.n7 24.5923
R2613 VN.n13 VN.n12 24.5923
R2614 VN.n18 VN.n5 24.5923
R2615 VN.n19 VN.n18 24.5923
R2616 VN.n21 VN.n3 24.5923
R2617 VN.n25 VN.n3 24.5923
R2618 VN.n26 VN.n25 24.5923
R2619 VN.n31 VN.n1 24.5923
R2620 VN.n32 VN.n31 24.5923
R2621 VN.n48 VN.n47 24.5923
R2622 VN.n47 VN.n42 24.5923
R2623 VN.n61 VN.n60 24.5923
R2624 VN.n60 VN.n38 24.5923
R2625 VN.n56 VN.n38 24.5923
R2626 VN.n54 VN.n53 24.5923
R2627 VN.n53 VN.n40 24.5923
R2628 VN.n67 VN.n66 24.5923
R2629 VN.n66 VN.n36 24.5923
R2630 VN.n8 VN.n7 24.3464
R2631 VN.n20 VN.n19 24.3464
R2632 VN.n43 VN.n42 24.3464
R2633 VN.n55 VN.n54 24.3464
R2634 VN.n33 VN.n32 23.8546
R2635 VN.n68 VN.n67 23.8546
R2636 VN.n45 VN.n44 2.54067
R2637 VN.n10 VN.n9 2.54067
R2638 VN.n69 VN.n35 0.417304
R2639 VN.n34 VN.n0 0.417304
R2640 VN VN.n34 0.394524
R2641 VN.n21 VN.n20 0.246418
R2642 VN.n56 VN.n55 0.246418
R2643 VN.n65 VN.n35 0.189894
R2644 VN.n65 VN.n64 0.189894
R2645 VN.n64 VN.n63 0.189894
R2646 VN.n63 VN.n37 0.189894
R2647 VN.n59 VN.n37 0.189894
R2648 VN.n59 VN.n58 0.189894
R2649 VN.n58 VN.n57 0.189894
R2650 VN.n57 VN.n39 0.189894
R2651 VN.n52 VN.n39 0.189894
R2652 VN.n52 VN.n51 0.189894
R2653 VN.n51 VN.n50 0.189894
R2654 VN.n50 VN.n41 0.189894
R2655 VN.n46 VN.n41 0.189894
R2656 VN.n46 VN.n45 0.189894
R2657 VN.n11 VN.n10 0.189894
R2658 VN.n11 VN.n6 0.189894
R2659 VN.n15 VN.n6 0.189894
R2660 VN.n16 VN.n15 0.189894
R2661 VN.n17 VN.n16 0.189894
R2662 VN.n17 VN.n4 0.189894
R2663 VN.n22 VN.n4 0.189894
R2664 VN.n23 VN.n22 0.189894
R2665 VN.n24 VN.n23 0.189894
R2666 VN.n24 VN.n2 0.189894
R2667 VN.n28 VN.n2 0.189894
R2668 VN.n29 VN.n28 0.189894
R2669 VN.n30 VN.n29 0.189894
R2670 VN.n30 VN.n0 0.189894
R2671 VDD2.n2 VDD2.n1 66.657
R2672 VDD2.n2 VDD2.n0 66.657
R2673 VDD2 VDD2.n5 66.6542
R2674 VDD2.n4 VDD2.n3 64.9927
R2675 VDD2.n4 VDD2.n2 46.6075
R2676 VDD2.n5 VDD2.t0 2.30283
R2677 VDD2.n5 VDD2.t1 2.30283
R2678 VDD2.n3 VDD2.t5 2.30283
R2679 VDD2.n3 VDD2.t6 2.30283
R2680 VDD2.n1 VDD2.t4 2.30283
R2681 VDD2.n1 VDD2.t7 2.30283
R2682 VDD2.n0 VDD2.t2 2.30283
R2683 VDD2.n0 VDD2.t3 2.30283
R2684 VDD2 VDD2.n4 1.77852
C0 VP VTAIL 7.66402f
C1 VDD1 VDD2 2.32426f
C2 VP VN 8.32753f
C3 VTAIL VDD1 7.56067f
C4 VTAIL VDD2 7.62219f
C5 VN VDD1 0.153555f
C6 VN VDD2 6.74248f
C7 VP VDD1 7.21937f
C8 VN VTAIL 7.64992f
C9 VP VDD2 0.632377f
C10 VDD2 B 6.214278f
C11 VDD1 B 6.77614f
C12 VTAIL B 9.139993f
C13 VN B 19.37973f
C14 VP B 18.050463f
C15 VDD2.t2 B 0.188905f
C16 VDD2.t3 B 0.188905f
C17 VDD2.n0 B 1.66307f
C18 VDD2.t4 B 0.188905f
C19 VDD2.t7 B 0.188905f
C20 VDD2.n1 B 1.66307f
C21 VDD2.n2 B 4.07763f
C22 VDD2.t5 B 0.188905f
C23 VDD2.t6 B 0.188905f
C24 VDD2.n3 B 1.64582f
C25 VDD2.n4 B 3.3948f
C26 VDD2.t0 B 0.188905f
C27 VDD2.t1 B 0.188905f
C28 VDD2.n5 B 1.66302f
C29 VN.n0 B 0.035273f
C30 VN.t0 B 1.59048f
C31 VN.n1 B 0.037258f
C32 VN.n2 B 0.018758f
C33 VN.n3 B 0.034784f
C34 VN.n4 B 0.018758f
C35 VN.t3 B 1.59048f
C36 VN.n5 B 0.037084f
C37 VN.n6 B 0.018758f
C38 VN.n7 B 0.034612f
C39 VN.t5 B 1.84938f
C40 VN.t4 B 1.59048f
C41 VN.n8 B 0.644455f
C42 VN.n9 B 0.612856f
C43 VN.n10 B 0.239239f
C44 VN.n11 B 0.018758f
C45 VN.n12 B 0.034784f
C46 VN.n13 B 0.037084f
C47 VN.n14 B 0.01515f
C48 VN.n15 B 0.018758f
C49 VN.n16 B 0.018758f
C50 VN.n17 B 0.018758f
C51 VN.n18 B 0.034784f
C52 VN.n19 B 0.034612f
C53 VN.n20 B 0.568711f
C54 VN.n21 B 0.017784f
C55 VN.n22 B 0.018758f
C56 VN.n23 B 0.018758f
C57 VN.n24 B 0.018758f
C58 VN.n25 B 0.034784f
C59 VN.n26 B 0.036886f
C60 VN.n27 B 0.015174f
C61 VN.n28 B 0.018758f
C62 VN.n29 B 0.018758f
C63 VN.n30 B 0.018758f
C64 VN.n31 B 0.034784f
C65 VN.n32 B 0.034269f
C66 VN.n33 B 0.650082f
C67 VN.n34 B 0.053476f
C68 VN.n35 B 0.035273f
C69 VN.t2 B 1.59048f
C70 VN.n36 B 0.037258f
C71 VN.n37 B 0.018758f
C72 VN.n38 B 0.034784f
C73 VN.n39 B 0.018758f
C74 VN.t1 B 1.59048f
C75 VN.n40 B 0.037084f
C76 VN.n41 B 0.018758f
C77 VN.n42 B 0.034612f
C78 VN.t6 B 1.84938f
C79 VN.t7 B 1.59048f
C80 VN.n43 B 0.644455f
C81 VN.n44 B 0.612856f
C82 VN.n45 B 0.239239f
C83 VN.n46 B 0.018758f
C84 VN.n47 B 0.034784f
C85 VN.n48 B 0.037084f
C86 VN.n49 B 0.01515f
C87 VN.n50 B 0.018758f
C88 VN.n51 B 0.018758f
C89 VN.n52 B 0.018758f
C90 VN.n53 B 0.034784f
C91 VN.n54 B 0.034612f
C92 VN.n55 B 0.568711f
C93 VN.n56 B 0.017784f
C94 VN.n57 B 0.018758f
C95 VN.n58 B 0.018758f
C96 VN.n59 B 0.018758f
C97 VN.n60 B 0.034784f
C98 VN.n61 B 0.036886f
C99 VN.n62 B 0.015174f
C100 VN.n63 B 0.018758f
C101 VN.n64 B 0.018758f
C102 VN.n65 B 0.018758f
C103 VN.n66 B 0.034784f
C104 VN.n67 B 0.034269f
C105 VN.n68 B 0.650082f
C106 VN.n69 B 1.19604f
C107 VTAIL.t7 B 0.151247f
C108 VTAIL.t1 B 0.151247f
C109 VTAIL.n0 B 1.25771f
C110 VTAIL.n1 B 0.458637f
C111 VTAIL.n2 B 0.02948f
C112 VTAIL.n3 B 0.022255f
C113 VTAIL.n4 B 0.011959f
C114 VTAIL.n5 B 0.028267f
C115 VTAIL.n6 B 0.012663f
C116 VTAIL.n7 B 0.022255f
C117 VTAIL.n8 B 0.011959f
C118 VTAIL.n9 B 0.028267f
C119 VTAIL.n10 B 0.012663f
C120 VTAIL.n11 B 0.022255f
C121 VTAIL.n12 B 0.011959f
C122 VTAIL.n13 B 0.028267f
C123 VTAIL.n14 B 0.012663f
C124 VTAIL.n15 B 0.13142f
C125 VTAIL.t6 B 0.04734f
C126 VTAIL.n16 B 0.0212f
C127 VTAIL.n17 B 0.019983f
C128 VTAIL.n18 B 0.011959f
C129 VTAIL.n19 B 0.786162f
C130 VTAIL.n20 B 0.022255f
C131 VTAIL.n21 B 0.011959f
C132 VTAIL.n22 B 0.012663f
C133 VTAIL.n23 B 0.028267f
C134 VTAIL.n24 B 0.028267f
C135 VTAIL.n25 B 0.012663f
C136 VTAIL.n26 B 0.011959f
C137 VTAIL.n27 B 0.022255f
C138 VTAIL.n28 B 0.022255f
C139 VTAIL.n29 B 0.011959f
C140 VTAIL.n30 B 0.012663f
C141 VTAIL.n31 B 0.028267f
C142 VTAIL.n32 B 0.028267f
C143 VTAIL.n33 B 0.028267f
C144 VTAIL.n34 B 0.012663f
C145 VTAIL.n35 B 0.011959f
C146 VTAIL.n36 B 0.022255f
C147 VTAIL.n37 B 0.022255f
C148 VTAIL.n38 B 0.011959f
C149 VTAIL.n39 B 0.012311f
C150 VTAIL.n40 B 0.012311f
C151 VTAIL.n41 B 0.028267f
C152 VTAIL.n42 B 0.058006f
C153 VTAIL.n43 B 0.012663f
C154 VTAIL.n44 B 0.011959f
C155 VTAIL.n45 B 0.053874f
C156 VTAIL.n46 B 0.032203f
C157 VTAIL.n47 B 0.300737f
C158 VTAIL.n48 B 0.02948f
C159 VTAIL.n49 B 0.022255f
C160 VTAIL.n50 B 0.011959f
C161 VTAIL.n51 B 0.028267f
C162 VTAIL.n52 B 0.012663f
C163 VTAIL.n53 B 0.022255f
C164 VTAIL.n54 B 0.011959f
C165 VTAIL.n55 B 0.028267f
C166 VTAIL.n56 B 0.012663f
C167 VTAIL.n57 B 0.022255f
C168 VTAIL.n58 B 0.011959f
C169 VTAIL.n59 B 0.028267f
C170 VTAIL.n60 B 0.012663f
C171 VTAIL.n61 B 0.13142f
C172 VTAIL.t13 B 0.04734f
C173 VTAIL.n62 B 0.0212f
C174 VTAIL.n63 B 0.019983f
C175 VTAIL.n64 B 0.011959f
C176 VTAIL.n65 B 0.786162f
C177 VTAIL.n66 B 0.022255f
C178 VTAIL.n67 B 0.011959f
C179 VTAIL.n68 B 0.012663f
C180 VTAIL.n69 B 0.028267f
C181 VTAIL.n70 B 0.028267f
C182 VTAIL.n71 B 0.012663f
C183 VTAIL.n72 B 0.011959f
C184 VTAIL.n73 B 0.022255f
C185 VTAIL.n74 B 0.022255f
C186 VTAIL.n75 B 0.011959f
C187 VTAIL.n76 B 0.012663f
C188 VTAIL.n77 B 0.028267f
C189 VTAIL.n78 B 0.028267f
C190 VTAIL.n79 B 0.028267f
C191 VTAIL.n80 B 0.012663f
C192 VTAIL.n81 B 0.011959f
C193 VTAIL.n82 B 0.022255f
C194 VTAIL.n83 B 0.022255f
C195 VTAIL.n84 B 0.011959f
C196 VTAIL.n85 B 0.012311f
C197 VTAIL.n86 B 0.012311f
C198 VTAIL.n87 B 0.028267f
C199 VTAIL.n88 B 0.058006f
C200 VTAIL.n89 B 0.012663f
C201 VTAIL.n90 B 0.011959f
C202 VTAIL.n91 B 0.053874f
C203 VTAIL.n92 B 0.032203f
C204 VTAIL.n93 B 0.300737f
C205 VTAIL.t8 B 0.151247f
C206 VTAIL.t14 B 0.151247f
C207 VTAIL.n94 B 1.25771f
C208 VTAIL.n95 B 0.701128f
C209 VTAIL.n96 B 0.02948f
C210 VTAIL.n97 B 0.022255f
C211 VTAIL.n98 B 0.011959f
C212 VTAIL.n99 B 0.028267f
C213 VTAIL.n100 B 0.012663f
C214 VTAIL.n101 B 0.022255f
C215 VTAIL.n102 B 0.011959f
C216 VTAIL.n103 B 0.028267f
C217 VTAIL.n104 B 0.012663f
C218 VTAIL.n105 B 0.022255f
C219 VTAIL.n106 B 0.011959f
C220 VTAIL.n107 B 0.028267f
C221 VTAIL.n108 B 0.012663f
C222 VTAIL.n109 B 0.13142f
C223 VTAIL.t9 B 0.04734f
C224 VTAIL.n110 B 0.0212f
C225 VTAIL.n111 B 0.019983f
C226 VTAIL.n112 B 0.011959f
C227 VTAIL.n113 B 0.786162f
C228 VTAIL.n114 B 0.022255f
C229 VTAIL.n115 B 0.011959f
C230 VTAIL.n116 B 0.012663f
C231 VTAIL.n117 B 0.028267f
C232 VTAIL.n118 B 0.028267f
C233 VTAIL.n119 B 0.012663f
C234 VTAIL.n120 B 0.011959f
C235 VTAIL.n121 B 0.022255f
C236 VTAIL.n122 B 0.022255f
C237 VTAIL.n123 B 0.011959f
C238 VTAIL.n124 B 0.012663f
C239 VTAIL.n125 B 0.028267f
C240 VTAIL.n126 B 0.028267f
C241 VTAIL.n127 B 0.028267f
C242 VTAIL.n128 B 0.012663f
C243 VTAIL.n129 B 0.011959f
C244 VTAIL.n130 B 0.022255f
C245 VTAIL.n131 B 0.022255f
C246 VTAIL.n132 B 0.011959f
C247 VTAIL.n133 B 0.012311f
C248 VTAIL.n134 B 0.012311f
C249 VTAIL.n135 B 0.028267f
C250 VTAIL.n136 B 0.058006f
C251 VTAIL.n137 B 0.012663f
C252 VTAIL.n138 B 0.011959f
C253 VTAIL.n139 B 0.053874f
C254 VTAIL.n140 B 0.032203f
C255 VTAIL.n141 B 1.34768f
C256 VTAIL.n142 B 0.02948f
C257 VTAIL.n143 B 0.022255f
C258 VTAIL.n144 B 0.011959f
C259 VTAIL.n145 B 0.028267f
C260 VTAIL.n146 B 0.012663f
C261 VTAIL.n147 B 0.022255f
C262 VTAIL.n148 B 0.011959f
C263 VTAIL.n149 B 0.028267f
C264 VTAIL.n150 B 0.028267f
C265 VTAIL.n151 B 0.012663f
C266 VTAIL.n152 B 0.022255f
C267 VTAIL.n153 B 0.011959f
C268 VTAIL.n154 B 0.028267f
C269 VTAIL.n155 B 0.012663f
C270 VTAIL.n156 B 0.13142f
C271 VTAIL.t3 B 0.04734f
C272 VTAIL.n157 B 0.0212f
C273 VTAIL.n158 B 0.019983f
C274 VTAIL.n159 B 0.011959f
C275 VTAIL.n160 B 0.786162f
C276 VTAIL.n161 B 0.022255f
C277 VTAIL.n162 B 0.011959f
C278 VTAIL.n163 B 0.012663f
C279 VTAIL.n164 B 0.028267f
C280 VTAIL.n165 B 0.028267f
C281 VTAIL.n166 B 0.012663f
C282 VTAIL.n167 B 0.011959f
C283 VTAIL.n168 B 0.022255f
C284 VTAIL.n169 B 0.022255f
C285 VTAIL.n170 B 0.011959f
C286 VTAIL.n171 B 0.012663f
C287 VTAIL.n172 B 0.028267f
C288 VTAIL.n173 B 0.028267f
C289 VTAIL.n174 B 0.012663f
C290 VTAIL.n175 B 0.011959f
C291 VTAIL.n176 B 0.022255f
C292 VTAIL.n177 B 0.022255f
C293 VTAIL.n178 B 0.011959f
C294 VTAIL.n179 B 0.012311f
C295 VTAIL.n180 B 0.012311f
C296 VTAIL.n181 B 0.028267f
C297 VTAIL.n182 B 0.058006f
C298 VTAIL.n183 B 0.012663f
C299 VTAIL.n184 B 0.011959f
C300 VTAIL.n185 B 0.053874f
C301 VTAIL.n186 B 0.032203f
C302 VTAIL.n187 B 1.34768f
C303 VTAIL.t4 B 0.151247f
C304 VTAIL.t0 B 0.151247f
C305 VTAIL.n188 B 1.25772f
C306 VTAIL.n189 B 0.70112f
C307 VTAIL.n190 B 0.02948f
C308 VTAIL.n191 B 0.022255f
C309 VTAIL.n192 B 0.011959f
C310 VTAIL.n193 B 0.028267f
C311 VTAIL.n194 B 0.012663f
C312 VTAIL.n195 B 0.022255f
C313 VTAIL.n196 B 0.011959f
C314 VTAIL.n197 B 0.028267f
C315 VTAIL.n198 B 0.028267f
C316 VTAIL.n199 B 0.012663f
C317 VTAIL.n200 B 0.022255f
C318 VTAIL.n201 B 0.011959f
C319 VTAIL.n202 B 0.028267f
C320 VTAIL.n203 B 0.012663f
C321 VTAIL.n204 B 0.13142f
C322 VTAIL.t5 B 0.04734f
C323 VTAIL.n205 B 0.0212f
C324 VTAIL.n206 B 0.019983f
C325 VTAIL.n207 B 0.011959f
C326 VTAIL.n208 B 0.786162f
C327 VTAIL.n209 B 0.022255f
C328 VTAIL.n210 B 0.011959f
C329 VTAIL.n211 B 0.012663f
C330 VTAIL.n212 B 0.028267f
C331 VTAIL.n213 B 0.028267f
C332 VTAIL.n214 B 0.012663f
C333 VTAIL.n215 B 0.011959f
C334 VTAIL.n216 B 0.022255f
C335 VTAIL.n217 B 0.022255f
C336 VTAIL.n218 B 0.011959f
C337 VTAIL.n219 B 0.012663f
C338 VTAIL.n220 B 0.028267f
C339 VTAIL.n221 B 0.028267f
C340 VTAIL.n222 B 0.012663f
C341 VTAIL.n223 B 0.011959f
C342 VTAIL.n224 B 0.022255f
C343 VTAIL.n225 B 0.022255f
C344 VTAIL.n226 B 0.011959f
C345 VTAIL.n227 B 0.012311f
C346 VTAIL.n228 B 0.012311f
C347 VTAIL.n229 B 0.028267f
C348 VTAIL.n230 B 0.058006f
C349 VTAIL.n231 B 0.012663f
C350 VTAIL.n232 B 0.011959f
C351 VTAIL.n233 B 0.053874f
C352 VTAIL.n234 B 0.032203f
C353 VTAIL.n235 B 0.300737f
C354 VTAIL.n236 B 0.02948f
C355 VTAIL.n237 B 0.022255f
C356 VTAIL.n238 B 0.011959f
C357 VTAIL.n239 B 0.028267f
C358 VTAIL.n240 B 0.012663f
C359 VTAIL.n241 B 0.022255f
C360 VTAIL.n242 B 0.011959f
C361 VTAIL.n243 B 0.028267f
C362 VTAIL.n244 B 0.028267f
C363 VTAIL.n245 B 0.012663f
C364 VTAIL.n246 B 0.022255f
C365 VTAIL.n247 B 0.011959f
C366 VTAIL.n248 B 0.028267f
C367 VTAIL.n249 B 0.012663f
C368 VTAIL.n250 B 0.13142f
C369 VTAIL.t15 B 0.04734f
C370 VTAIL.n251 B 0.0212f
C371 VTAIL.n252 B 0.019983f
C372 VTAIL.n253 B 0.011959f
C373 VTAIL.n254 B 0.786162f
C374 VTAIL.n255 B 0.022255f
C375 VTAIL.n256 B 0.011959f
C376 VTAIL.n257 B 0.012663f
C377 VTAIL.n258 B 0.028267f
C378 VTAIL.n259 B 0.028267f
C379 VTAIL.n260 B 0.012663f
C380 VTAIL.n261 B 0.011959f
C381 VTAIL.n262 B 0.022255f
C382 VTAIL.n263 B 0.022255f
C383 VTAIL.n264 B 0.011959f
C384 VTAIL.n265 B 0.012663f
C385 VTAIL.n266 B 0.028267f
C386 VTAIL.n267 B 0.028267f
C387 VTAIL.n268 B 0.012663f
C388 VTAIL.n269 B 0.011959f
C389 VTAIL.n270 B 0.022255f
C390 VTAIL.n271 B 0.022255f
C391 VTAIL.n272 B 0.011959f
C392 VTAIL.n273 B 0.012311f
C393 VTAIL.n274 B 0.012311f
C394 VTAIL.n275 B 0.028267f
C395 VTAIL.n276 B 0.058006f
C396 VTAIL.n277 B 0.012663f
C397 VTAIL.n278 B 0.011959f
C398 VTAIL.n279 B 0.053874f
C399 VTAIL.n280 B 0.032203f
C400 VTAIL.n281 B 0.300737f
C401 VTAIL.t12 B 0.151247f
C402 VTAIL.t10 B 0.151247f
C403 VTAIL.n282 B 1.25772f
C404 VTAIL.n283 B 0.70112f
C405 VTAIL.n284 B 0.02948f
C406 VTAIL.n285 B 0.022255f
C407 VTAIL.n286 B 0.011959f
C408 VTAIL.n287 B 0.028267f
C409 VTAIL.n288 B 0.012663f
C410 VTAIL.n289 B 0.022255f
C411 VTAIL.n290 B 0.011959f
C412 VTAIL.n291 B 0.028267f
C413 VTAIL.n292 B 0.028267f
C414 VTAIL.n293 B 0.012663f
C415 VTAIL.n294 B 0.022255f
C416 VTAIL.n295 B 0.011959f
C417 VTAIL.n296 B 0.028267f
C418 VTAIL.n297 B 0.012663f
C419 VTAIL.n298 B 0.13142f
C420 VTAIL.t11 B 0.04734f
C421 VTAIL.n299 B 0.0212f
C422 VTAIL.n300 B 0.019983f
C423 VTAIL.n301 B 0.011959f
C424 VTAIL.n302 B 0.786162f
C425 VTAIL.n303 B 0.022255f
C426 VTAIL.n304 B 0.011959f
C427 VTAIL.n305 B 0.012663f
C428 VTAIL.n306 B 0.028267f
C429 VTAIL.n307 B 0.028267f
C430 VTAIL.n308 B 0.012663f
C431 VTAIL.n309 B 0.011959f
C432 VTAIL.n310 B 0.022255f
C433 VTAIL.n311 B 0.022255f
C434 VTAIL.n312 B 0.011959f
C435 VTAIL.n313 B 0.012663f
C436 VTAIL.n314 B 0.028267f
C437 VTAIL.n315 B 0.028267f
C438 VTAIL.n316 B 0.012663f
C439 VTAIL.n317 B 0.011959f
C440 VTAIL.n318 B 0.022255f
C441 VTAIL.n319 B 0.022255f
C442 VTAIL.n320 B 0.011959f
C443 VTAIL.n321 B 0.012311f
C444 VTAIL.n322 B 0.012311f
C445 VTAIL.n323 B 0.028267f
C446 VTAIL.n324 B 0.058006f
C447 VTAIL.n325 B 0.012663f
C448 VTAIL.n326 B 0.011959f
C449 VTAIL.n327 B 0.053874f
C450 VTAIL.n328 B 0.032203f
C451 VTAIL.n329 B 1.34768f
C452 VTAIL.n330 B 0.02948f
C453 VTAIL.n331 B 0.022255f
C454 VTAIL.n332 B 0.011959f
C455 VTAIL.n333 B 0.028267f
C456 VTAIL.n334 B 0.012663f
C457 VTAIL.n335 B 0.022255f
C458 VTAIL.n336 B 0.011959f
C459 VTAIL.n337 B 0.028267f
C460 VTAIL.n338 B 0.012663f
C461 VTAIL.n339 B 0.022255f
C462 VTAIL.n340 B 0.011959f
C463 VTAIL.n341 B 0.028267f
C464 VTAIL.n342 B 0.012663f
C465 VTAIL.n343 B 0.13142f
C466 VTAIL.t2 B 0.04734f
C467 VTAIL.n344 B 0.0212f
C468 VTAIL.n345 B 0.019983f
C469 VTAIL.n346 B 0.011959f
C470 VTAIL.n347 B 0.786162f
C471 VTAIL.n348 B 0.022255f
C472 VTAIL.n349 B 0.011959f
C473 VTAIL.n350 B 0.012663f
C474 VTAIL.n351 B 0.028267f
C475 VTAIL.n352 B 0.028267f
C476 VTAIL.n353 B 0.012663f
C477 VTAIL.n354 B 0.011959f
C478 VTAIL.n355 B 0.022255f
C479 VTAIL.n356 B 0.022255f
C480 VTAIL.n357 B 0.011959f
C481 VTAIL.n358 B 0.012663f
C482 VTAIL.n359 B 0.028267f
C483 VTAIL.n360 B 0.028267f
C484 VTAIL.n361 B 0.028267f
C485 VTAIL.n362 B 0.012663f
C486 VTAIL.n363 B 0.011959f
C487 VTAIL.n364 B 0.022255f
C488 VTAIL.n365 B 0.022255f
C489 VTAIL.n366 B 0.011959f
C490 VTAIL.n367 B 0.012311f
C491 VTAIL.n368 B 0.012311f
C492 VTAIL.n369 B 0.028267f
C493 VTAIL.n370 B 0.058006f
C494 VTAIL.n371 B 0.012663f
C495 VTAIL.n372 B 0.011959f
C496 VTAIL.n373 B 0.053874f
C497 VTAIL.n374 B 0.032203f
C498 VTAIL.n375 B 1.3435f
C499 VDD1.t0 B 0.193399f
C500 VDD1.t7 B 0.193399f
C501 VDD1.n0 B 1.70408f
C502 VDD1.t5 B 0.193399f
C503 VDD1.t4 B 0.193399f
C504 VDD1.n1 B 1.70263f
C505 VDD1.t2 B 0.193399f
C506 VDD1.t6 B 0.193399f
C507 VDD1.n2 B 1.70263f
C508 VDD1.n3 B 4.23339f
C509 VDD1.t1 B 0.193399f
C510 VDD1.t3 B 0.193399f
C511 VDD1.n4 B 1.68496f
C512 VDD1.n5 B 3.51124f
C513 VP.n0 B 0.036251f
C514 VP.t2 B 1.63462f
C515 VP.n1 B 0.038292f
C516 VP.n2 B 0.019278f
C517 VP.n3 B 0.035749f
C518 VP.n4 B 0.019278f
C519 VP.t1 B 1.63462f
C520 VP.n5 B 0.038113f
C521 VP.n6 B 0.019278f
C522 VP.n7 B 0.035573f
C523 VP.n8 B 0.019278f
C524 VP.n9 B 0.03791f
C525 VP.n10 B 0.019278f
C526 VP.n11 B 0.03522f
C527 VP.n12 B 0.036251f
C528 VP.t4 B 1.63462f
C529 VP.n13 B 0.038292f
C530 VP.n14 B 0.019278f
C531 VP.n15 B 0.035749f
C532 VP.n16 B 0.019278f
C533 VP.t5 B 1.63462f
C534 VP.n17 B 0.038113f
C535 VP.n18 B 0.019278f
C536 VP.n19 B 0.035573f
C537 VP.t0 B 1.90069f
C538 VP.t3 B 1.63462f
C539 VP.n20 B 0.662337f
C540 VP.n21 B 0.629863f
C541 VP.n22 B 0.245877f
C542 VP.n23 B 0.019278f
C543 VP.n24 B 0.035749f
C544 VP.n25 B 0.038113f
C545 VP.n26 B 0.01557f
C546 VP.n27 B 0.019278f
C547 VP.n28 B 0.019278f
C548 VP.n29 B 0.019278f
C549 VP.n30 B 0.035749f
C550 VP.n31 B 0.035573f
C551 VP.n32 B 0.584491f
C552 VP.n33 B 0.018277f
C553 VP.n34 B 0.019278f
C554 VP.n35 B 0.019278f
C555 VP.n36 B 0.019278f
C556 VP.n37 B 0.035749f
C557 VP.n38 B 0.03791f
C558 VP.n39 B 0.015595f
C559 VP.n40 B 0.019278f
C560 VP.n41 B 0.019278f
C561 VP.n42 B 0.019278f
C562 VP.n43 B 0.035749f
C563 VP.n44 B 0.03522f
C564 VP.n45 B 0.66812f
C565 VP.n46 B 1.22443f
C566 VP.t6 B 1.63462f
C567 VP.n47 B 0.66812f
C568 VP.n48 B 1.23742f
C569 VP.n49 B 0.036251f
C570 VP.n50 B 0.019278f
C571 VP.n51 B 0.035749f
C572 VP.n52 B 0.038292f
C573 VP.n53 B 0.015595f
C574 VP.n54 B 0.019278f
C575 VP.n55 B 0.019278f
C576 VP.n56 B 0.019278f
C577 VP.n57 B 0.035749f
C578 VP.n58 B 0.035749f
C579 VP.t7 B 1.63462f
C580 VP.n59 B 0.584491f
C581 VP.n60 B 0.018277f
C582 VP.n61 B 0.019278f
C583 VP.n62 B 0.019278f
C584 VP.n63 B 0.019278f
C585 VP.n64 B 0.035749f
C586 VP.n65 B 0.038113f
C587 VP.n66 B 0.01557f
C588 VP.n67 B 0.019278f
C589 VP.n68 B 0.019278f
C590 VP.n69 B 0.019278f
C591 VP.n70 B 0.035749f
C592 VP.n71 B 0.035573f
C593 VP.n72 B 0.584491f
C594 VP.n73 B 0.018277f
C595 VP.n74 B 0.019278f
C596 VP.n75 B 0.019278f
C597 VP.n76 B 0.019278f
C598 VP.n77 B 0.035749f
C599 VP.n78 B 0.03791f
C600 VP.n79 B 0.015595f
C601 VP.n80 B 0.019278f
C602 VP.n81 B 0.019278f
C603 VP.n82 B 0.019278f
C604 VP.n83 B 0.035749f
C605 VP.n84 B 0.03522f
C606 VP.n85 B 0.66812f
C607 VP.n86 B 0.05496f
.ends

