* NGSPICE file created from diff_pair_sample_1757.ext - technology: sky130A

.subckt diff_pair_sample_1757 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X1 VDD1.t9 VP.t0 VTAIL.t0 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X2 B.t11 B.t9 B.t10 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=0 ps=0 w=17.24 l=1.29
X3 VDD1.t8 VP.t1 VTAIL.t1 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=6.7236 ps=35.26 w=17.24 l=1.29
X4 VDD1.t7 VP.t2 VTAIL.t2 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=6.7236 ps=35.26 w=17.24 l=1.29
X5 VTAIL.t5 VP.t3 VDD1.t6 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X6 VTAIL.t8 VP.t4 VDD1.t5 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X7 VDD1.t4 VP.t5 VTAIL.t3 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=2.8446 ps=17.57 w=17.24 l=1.29
X8 VTAIL.t6 VP.t6 VDD1.t3 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X9 VDD2.t8 VN.t1 VTAIL.t12 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=6.7236 ps=35.26 w=17.24 l=1.29
X10 VDD1.t2 VP.t7 VTAIL.t7 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X11 VTAIL.t14 VN.t2 VDD2.t7 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X12 VTAIL.t17 VN.t3 VDD2.t6 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X13 VDD2.t5 VN.t4 VTAIL.t16 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=6.7236 ps=35.26 w=17.24 l=1.29
X14 VDD2.t4 VN.t5 VTAIL.t10 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=2.8446 ps=17.57 w=17.24 l=1.29
X15 VTAIL.t15 VN.t6 VDD2.t3 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X16 B.t8 B.t6 B.t7 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=0 ps=0 w=17.24 l=1.29
X17 VDD2.t2 VN.t7 VTAIL.t19 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X18 VTAIL.t18 VN.t8 VDD2.t1 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X19 VDD1.t1 VP.t8 VTAIL.t9 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=2.8446 ps=17.57 w=17.24 l=1.29
X20 VTAIL.t4 VP.t9 VDD1.t0 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=2.8446 pd=17.57 as=2.8446 ps=17.57 w=17.24 l=1.29
X21 B.t5 B.t3 B.t4 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=0 ps=0 w=17.24 l=1.29
X22 VDD2.t0 VN.t9 VTAIL.t13 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=2.8446 ps=17.57 w=17.24 l=1.29
X23 B.t2 B.t0 B.t1 w_n2914_n4416# sky130_fd_pr__pfet_01v8 ad=6.7236 pd=35.26 as=0 ps=0 w=17.24 l=1.29
R0 VN.n6 VN.t5 351.041
R1 VN.n32 VN.t1 351.041
R2 VN.n3 VN.t7 322.082
R3 VN.n5 VN.t8 322.082
R4 VN.n16 VN.t3 322.082
R5 VN.n23 VN.t4 322.082
R6 VN.n29 VN.t0 322.082
R7 VN.n31 VN.t6 322.082
R8 VN.n28 VN.t2 322.082
R9 VN.n48 VN.t9 322.082
R10 VN.n24 VN.n23 174.089
R11 VN.n49 VN.n48 174.089
R12 VN.n47 VN.n25 161.3
R13 VN.n46 VN.n45 161.3
R14 VN.n44 VN.n26 161.3
R15 VN.n43 VN.n42 161.3
R16 VN.n41 VN.n27 161.3
R17 VN.n40 VN.n39 161.3
R18 VN.n38 VN.n29 161.3
R19 VN.n37 VN.n36 161.3
R20 VN.n35 VN.n30 161.3
R21 VN.n34 VN.n33 161.3
R22 VN.n22 VN.n0 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n19 VN.n1 161.3
R25 VN.n18 VN.n17 161.3
R26 VN.n15 VN.n2 161.3
R27 VN.n14 VN.n13 161.3
R28 VN.n12 VN.n3 161.3
R29 VN.n11 VN.n10 161.3
R30 VN.n9 VN.n4 161.3
R31 VN.n8 VN.n7 161.3
R32 VN.n6 VN.n5 59.2496
R33 VN.n32 VN.n31 59.2496
R34 VN.n10 VN.n9 56.5617
R35 VN.n15 VN.n14 56.5617
R36 VN.n36 VN.n35 56.5617
R37 VN.n41 VN.n40 56.5617
R38 VN VN.n49 50.2448
R39 VN.n21 VN.n1 47.3584
R40 VN.n46 VN.n26 47.3584
R41 VN.n22 VN.n21 33.7956
R42 VN.n47 VN.n46 33.7956
R43 VN.n33 VN.n32 27.2704
R44 VN.n7 VN.n6 27.2704
R45 VN.n9 VN.n8 24.5923
R46 VN.n10 VN.n3 24.5923
R47 VN.n14 VN.n3 24.5923
R48 VN.n17 VN.n15 24.5923
R49 VN.n35 VN.n34 24.5923
R50 VN.n40 VN.n29 24.5923
R51 VN.n36 VN.n29 24.5923
R52 VN.n42 VN.n41 24.5923
R53 VN.n16 VN.n1 18.6903
R54 VN.n28 VN.n26 18.6903
R55 VN.n23 VN.n22 11.8046
R56 VN.n48 VN.n47 11.8046
R57 VN.n8 VN.n5 5.90254
R58 VN.n17 VN.n16 5.90254
R59 VN.n34 VN.n31 5.90254
R60 VN.n42 VN.n28 5.90254
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n30 0.189894
R70 VN.n33 VN.n30 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n11 VN.n4 0.189894
R73 VN.n12 VN.n11 0.189894
R74 VN.n13 VN.n12 0.189894
R75 VN.n13 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VTAIL.n11 VTAIL.t12 55.9603
R83 VTAIL.n17 VTAIL.t16 55.9602
R84 VTAIL.n2 VTAIL.t1 55.9602
R85 VTAIL.n16 VTAIL.t2 55.9602
R86 VTAIL.n15 VTAIL.n14 54.0749
R87 VTAIL.n13 VTAIL.n12 54.0749
R88 VTAIL.n10 VTAIL.n9 54.0749
R89 VTAIL.n8 VTAIL.n7 54.0749
R90 VTAIL.n19 VTAIL.n18 54.0747
R91 VTAIL.n1 VTAIL.n0 54.0747
R92 VTAIL.n4 VTAIL.n3 54.0747
R93 VTAIL.n6 VTAIL.n5 54.0747
R94 VTAIL.n8 VTAIL.n6 30.0221
R95 VTAIL.n17 VTAIL.n16 28.6255
R96 VTAIL.n18 VTAIL.t19 1.88594
R97 VTAIL.n18 VTAIL.t17 1.88594
R98 VTAIL.n0 VTAIL.t10 1.88594
R99 VTAIL.n0 VTAIL.t18 1.88594
R100 VTAIL.n3 VTAIL.t0 1.88594
R101 VTAIL.n3 VTAIL.t8 1.88594
R102 VTAIL.n5 VTAIL.t3 1.88594
R103 VTAIL.n5 VTAIL.t5 1.88594
R104 VTAIL.n14 VTAIL.t7 1.88594
R105 VTAIL.n14 VTAIL.t4 1.88594
R106 VTAIL.n12 VTAIL.t9 1.88594
R107 VTAIL.n12 VTAIL.t6 1.88594
R108 VTAIL.n9 VTAIL.t11 1.88594
R109 VTAIL.n9 VTAIL.t15 1.88594
R110 VTAIL.n7 VTAIL.t13 1.88594
R111 VTAIL.n7 VTAIL.t14 1.88594
R112 VTAIL.n10 VTAIL.n8 1.39705
R113 VTAIL.n11 VTAIL.n10 1.39705
R114 VTAIL.n15 VTAIL.n13 1.39705
R115 VTAIL.n16 VTAIL.n15 1.39705
R116 VTAIL.n6 VTAIL.n4 1.39705
R117 VTAIL.n4 VTAIL.n2 1.39705
R118 VTAIL.n19 VTAIL.n17 1.39705
R119 VTAIL.n13 VTAIL.n11 1.1686
R120 VTAIL.n2 VTAIL.n1 1.1686
R121 VTAIL VTAIL.n1 1.1061
R122 VTAIL VTAIL.n19 0.291448
R123 VDD2.n1 VDD2.t4 74.0355
R124 VDD2.n4 VDD2.t0 72.6391
R125 VDD2.n3 VDD2.n2 71.7455
R126 VDD2 VDD2.n7 71.7427
R127 VDD2.n6 VDD2.n5 70.7537
R128 VDD2.n1 VDD2.n0 70.7535
R129 VDD2.n4 VDD2.n3 45.211
R130 VDD2.n7 VDD2.t3 1.88594
R131 VDD2.n7 VDD2.t8 1.88594
R132 VDD2.n5 VDD2.t7 1.88594
R133 VDD2.n5 VDD2.t9 1.88594
R134 VDD2.n2 VDD2.t6 1.88594
R135 VDD2.n2 VDD2.t5 1.88594
R136 VDD2.n0 VDD2.t1 1.88594
R137 VDD2.n0 VDD2.t2 1.88594
R138 VDD2.n6 VDD2.n4 1.39705
R139 VDD2 VDD2.n6 0.407828
R140 VDD2.n3 VDD2.n1 0.294292
R141 VP.n14 VP.t8 351.041
R142 VP.n3 VP.t0 322.082
R143 VP.n7 VP.t5 322.082
R144 VP.n5 VP.t3 322.082
R145 VP.n48 VP.t4 322.082
R146 VP.n55 VP.t1 322.082
R147 VP.n11 VP.t7 322.082
R148 VP.n31 VP.t2 322.082
R149 VP.n24 VP.t9 322.082
R150 VP.n13 VP.t6 322.082
R151 VP.n33 VP.n7 174.089
R152 VP.n56 VP.n55 174.089
R153 VP.n32 VP.n31 174.089
R154 VP.n16 VP.n15 161.3
R155 VP.n17 VP.n12 161.3
R156 VP.n19 VP.n18 161.3
R157 VP.n20 VP.n11 161.3
R158 VP.n22 VP.n21 161.3
R159 VP.n23 VP.n10 161.3
R160 VP.n26 VP.n25 161.3
R161 VP.n27 VP.n9 161.3
R162 VP.n29 VP.n28 161.3
R163 VP.n30 VP.n8 161.3
R164 VP.n54 VP.n0 161.3
R165 VP.n53 VP.n52 161.3
R166 VP.n51 VP.n1 161.3
R167 VP.n50 VP.n49 161.3
R168 VP.n47 VP.n2 161.3
R169 VP.n46 VP.n45 161.3
R170 VP.n44 VP.n3 161.3
R171 VP.n43 VP.n42 161.3
R172 VP.n41 VP.n4 161.3
R173 VP.n40 VP.n39 161.3
R174 VP.n38 VP.n37 161.3
R175 VP.n36 VP.n6 161.3
R176 VP.n35 VP.n34 161.3
R177 VP.n14 VP.n13 59.2496
R178 VP.n42 VP.n41 56.5617
R179 VP.n47 VP.n46 56.5617
R180 VP.n23 VP.n22 56.5617
R181 VP.n18 VP.n17 56.5617
R182 VP.n33 VP.n32 49.8641
R183 VP.n37 VP.n36 47.3584
R184 VP.n53 VP.n1 47.3584
R185 VP.n29 VP.n9 47.3584
R186 VP.n36 VP.n35 33.7956
R187 VP.n54 VP.n53 33.7956
R188 VP.n30 VP.n29 33.7956
R189 VP.n15 VP.n14 27.2704
R190 VP.n41 VP.n40 24.5923
R191 VP.n42 VP.n3 24.5923
R192 VP.n46 VP.n3 24.5923
R193 VP.n49 VP.n47 24.5923
R194 VP.n25 VP.n23 24.5923
R195 VP.n18 VP.n11 24.5923
R196 VP.n22 VP.n11 24.5923
R197 VP.n17 VP.n16 24.5923
R198 VP.n37 VP.n5 18.6903
R199 VP.n48 VP.n1 18.6903
R200 VP.n24 VP.n9 18.6903
R201 VP.n35 VP.n7 11.8046
R202 VP.n55 VP.n54 11.8046
R203 VP.n31 VP.n30 11.8046
R204 VP.n40 VP.n5 5.90254
R205 VP.n49 VP.n48 5.90254
R206 VP.n25 VP.n24 5.90254
R207 VP.n16 VP.n13 5.90254
R208 VP.n15 VP.n12 0.189894
R209 VP.n19 VP.n12 0.189894
R210 VP.n20 VP.n19 0.189894
R211 VP.n21 VP.n20 0.189894
R212 VP.n21 VP.n10 0.189894
R213 VP.n26 VP.n10 0.189894
R214 VP.n27 VP.n26 0.189894
R215 VP.n28 VP.n27 0.189894
R216 VP.n28 VP.n8 0.189894
R217 VP.n32 VP.n8 0.189894
R218 VP.n34 VP.n33 0.189894
R219 VP.n34 VP.n6 0.189894
R220 VP.n38 VP.n6 0.189894
R221 VP.n39 VP.n38 0.189894
R222 VP.n39 VP.n4 0.189894
R223 VP.n43 VP.n4 0.189894
R224 VP.n44 VP.n43 0.189894
R225 VP.n45 VP.n44 0.189894
R226 VP.n45 VP.n2 0.189894
R227 VP.n50 VP.n2 0.189894
R228 VP.n51 VP.n50 0.189894
R229 VP.n52 VP.n51 0.189894
R230 VP.n52 VP.n0 0.189894
R231 VP.n56 VP.n0 0.189894
R232 VP VP.n56 0.0516364
R233 VDD1.n1 VDD1.t1 74.0356
R234 VDD1.n3 VDD1.t4 74.0355
R235 VDD1.n5 VDD1.n4 71.7455
R236 VDD1.n1 VDD1.n0 70.7537
R237 VDD1.n7 VDD1.n6 70.7535
R238 VDD1.n3 VDD1.n2 70.7535
R239 VDD1.n7 VDD1.n5 46.4923
R240 VDD1.n6 VDD1.t0 1.88594
R241 VDD1.n6 VDD1.t7 1.88594
R242 VDD1.n0 VDD1.t3 1.88594
R243 VDD1.n0 VDD1.t2 1.88594
R244 VDD1.n4 VDD1.t5 1.88594
R245 VDD1.n4 VDD1.t8 1.88594
R246 VDD1.n2 VDD1.t6 1.88594
R247 VDD1.n2 VDD1.t9 1.88594
R248 VDD1 VDD1.n7 0.989724
R249 VDD1 VDD1.n1 0.407828
R250 VDD1.n5 VDD1.n3 0.294292
R251 B.n447 B.n124 585
R252 B.n446 B.n445 585
R253 B.n444 B.n125 585
R254 B.n443 B.n442 585
R255 B.n441 B.n126 585
R256 B.n440 B.n439 585
R257 B.n438 B.n127 585
R258 B.n437 B.n436 585
R259 B.n435 B.n128 585
R260 B.n434 B.n433 585
R261 B.n432 B.n129 585
R262 B.n431 B.n430 585
R263 B.n429 B.n130 585
R264 B.n428 B.n427 585
R265 B.n426 B.n131 585
R266 B.n425 B.n424 585
R267 B.n423 B.n132 585
R268 B.n422 B.n421 585
R269 B.n420 B.n133 585
R270 B.n419 B.n418 585
R271 B.n417 B.n134 585
R272 B.n416 B.n415 585
R273 B.n414 B.n135 585
R274 B.n413 B.n412 585
R275 B.n411 B.n136 585
R276 B.n410 B.n409 585
R277 B.n408 B.n137 585
R278 B.n407 B.n406 585
R279 B.n405 B.n138 585
R280 B.n404 B.n403 585
R281 B.n402 B.n139 585
R282 B.n401 B.n400 585
R283 B.n399 B.n140 585
R284 B.n398 B.n397 585
R285 B.n396 B.n141 585
R286 B.n395 B.n394 585
R287 B.n393 B.n142 585
R288 B.n392 B.n391 585
R289 B.n390 B.n143 585
R290 B.n389 B.n388 585
R291 B.n387 B.n144 585
R292 B.n386 B.n385 585
R293 B.n384 B.n145 585
R294 B.n383 B.n382 585
R295 B.n381 B.n146 585
R296 B.n380 B.n379 585
R297 B.n378 B.n147 585
R298 B.n377 B.n376 585
R299 B.n375 B.n148 585
R300 B.n374 B.n373 585
R301 B.n372 B.n149 585
R302 B.n371 B.n370 585
R303 B.n369 B.n150 585
R304 B.n368 B.n367 585
R305 B.n366 B.n151 585
R306 B.n365 B.n364 585
R307 B.n363 B.n152 585
R308 B.n361 B.n360 585
R309 B.n359 B.n155 585
R310 B.n358 B.n357 585
R311 B.n356 B.n156 585
R312 B.n355 B.n354 585
R313 B.n353 B.n157 585
R314 B.n352 B.n351 585
R315 B.n350 B.n158 585
R316 B.n349 B.n348 585
R317 B.n347 B.n159 585
R318 B.n346 B.n345 585
R319 B.n341 B.n160 585
R320 B.n340 B.n339 585
R321 B.n338 B.n161 585
R322 B.n337 B.n336 585
R323 B.n335 B.n162 585
R324 B.n334 B.n333 585
R325 B.n332 B.n163 585
R326 B.n331 B.n330 585
R327 B.n329 B.n164 585
R328 B.n328 B.n327 585
R329 B.n326 B.n165 585
R330 B.n325 B.n324 585
R331 B.n323 B.n166 585
R332 B.n322 B.n321 585
R333 B.n320 B.n167 585
R334 B.n319 B.n318 585
R335 B.n317 B.n168 585
R336 B.n316 B.n315 585
R337 B.n314 B.n169 585
R338 B.n313 B.n312 585
R339 B.n311 B.n170 585
R340 B.n310 B.n309 585
R341 B.n308 B.n171 585
R342 B.n307 B.n306 585
R343 B.n305 B.n172 585
R344 B.n304 B.n303 585
R345 B.n302 B.n173 585
R346 B.n301 B.n300 585
R347 B.n299 B.n174 585
R348 B.n298 B.n297 585
R349 B.n296 B.n175 585
R350 B.n295 B.n294 585
R351 B.n293 B.n176 585
R352 B.n292 B.n291 585
R353 B.n290 B.n177 585
R354 B.n289 B.n288 585
R355 B.n287 B.n178 585
R356 B.n286 B.n285 585
R357 B.n284 B.n179 585
R358 B.n283 B.n282 585
R359 B.n281 B.n180 585
R360 B.n280 B.n279 585
R361 B.n278 B.n181 585
R362 B.n277 B.n276 585
R363 B.n275 B.n182 585
R364 B.n274 B.n273 585
R365 B.n272 B.n183 585
R366 B.n271 B.n270 585
R367 B.n269 B.n184 585
R368 B.n268 B.n267 585
R369 B.n266 B.n185 585
R370 B.n265 B.n264 585
R371 B.n263 B.n186 585
R372 B.n262 B.n261 585
R373 B.n260 B.n187 585
R374 B.n259 B.n258 585
R375 B.n449 B.n448 585
R376 B.n450 B.n123 585
R377 B.n452 B.n451 585
R378 B.n453 B.n122 585
R379 B.n455 B.n454 585
R380 B.n456 B.n121 585
R381 B.n458 B.n457 585
R382 B.n459 B.n120 585
R383 B.n461 B.n460 585
R384 B.n462 B.n119 585
R385 B.n464 B.n463 585
R386 B.n465 B.n118 585
R387 B.n467 B.n466 585
R388 B.n468 B.n117 585
R389 B.n470 B.n469 585
R390 B.n471 B.n116 585
R391 B.n473 B.n472 585
R392 B.n474 B.n115 585
R393 B.n476 B.n475 585
R394 B.n477 B.n114 585
R395 B.n479 B.n478 585
R396 B.n480 B.n113 585
R397 B.n482 B.n481 585
R398 B.n483 B.n112 585
R399 B.n485 B.n484 585
R400 B.n486 B.n111 585
R401 B.n488 B.n487 585
R402 B.n489 B.n110 585
R403 B.n491 B.n490 585
R404 B.n492 B.n109 585
R405 B.n494 B.n493 585
R406 B.n495 B.n108 585
R407 B.n497 B.n496 585
R408 B.n498 B.n107 585
R409 B.n500 B.n499 585
R410 B.n501 B.n106 585
R411 B.n503 B.n502 585
R412 B.n504 B.n105 585
R413 B.n506 B.n505 585
R414 B.n507 B.n104 585
R415 B.n509 B.n508 585
R416 B.n510 B.n103 585
R417 B.n512 B.n511 585
R418 B.n513 B.n102 585
R419 B.n515 B.n514 585
R420 B.n516 B.n101 585
R421 B.n518 B.n517 585
R422 B.n519 B.n100 585
R423 B.n521 B.n520 585
R424 B.n522 B.n99 585
R425 B.n524 B.n523 585
R426 B.n525 B.n98 585
R427 B.n527 B.n526 585
R428 B.n528 B.n97 585
R429 B.n530 B.n529 585
R430 B.n531 B.n96 585
R431 B.n533 B.n532 585
R432 B.n534 B.n95 585
R433 B.n536 B.n535 585
R434 B.n537 B.n94 585
R435 B.n539 B.n538 585
R436 B.n540 B.n93 585
R437 B.n542 B.n541 585
R438 B.n543 B.n92 585
R439 B.n545 B.n544 585
R440 B.n546 B.n91 585
R441 B.n548 B.n547 585
R442 B.n549 B.n90 585
R443 B.n551 B.n550 585
R444 B.n552 B.n89 585
R445 B.n554 B.n553 585
R446 B.n555 B.n88 585
R447 B.n557 B.n556 585
R448 B.n558 B.n87 585
R449 B.n745 B.n20 585
R450 B.n744 B.n743 585
R451 B.n742 B.n21 585
R452 B.n741 B.n740 585
R453 B.n739 B.n22 585
R454 B.n738 B.n737 585
R455 B.n736 B.n23 585
R456 B.n735 B.n734 585
R457 B.n733 B.n24 585
R458 B.n732 B.n731 585
R459 B.n730 B.n25 585
R460 B.n729 B.n728 585
R461 B.n727 B.n26 585
R462 B.n726 B.n725 585
R463 B.n724 B.n27 585
R464 B.n723 B.n722 585
R465 B.n721 B.n28 585
R466 B.n720 B.n719 585
R467 B.n718 B.n29 585
R468 B.n717 B.n716 585
R469 B.n715 B.n30 585
R470 B.n714 B.n713 585
R471 B.n712 B.n31 585
R472 B.n711 B.n710 585
R473 B.n709 B.n32 585
R474 B.n708 B.n707 585
R475 B.n706 B.n33 585
R476 B.n705 B.n704 585
R477 B.n703 B.n34 585
R478 B.n702 B.n701 585
R479 B.n700 B.n35 585
R480 B.n699 B.n698 585
R481 B.n697 B.n36 585
R482 B.n696 B.n695 585
R483 B.n694 B.n37 585
R484 B.n693 B.n692 585
R485 B.n691 B.n38 585
R486 B.n690 B.n689 585
R487 B.n688 B.n39 585
R488 B.n687 B.n686 585
R489 B.n685 B.n40 585
R490 B.n684 B.n683 585
R491 B.n682 B.n41 585
R492 B.n681 B.n680 585
R493 B.n679 B.n42 585
R494 B.n678 B.n677 585
R495 B.n676 B.n43 585
R496 B.n675 B.n674 585
R497 B.n673 B.n44 585
R498 B.n672 B.n671 585
R499 B.n670 B.n45 585
R500 B.n669 B.n668 585
R501 B.n667 B.n46 585
R502 B.n666 B.n665 585
R503 B.n664 B.n47 585
R504 B.n663 B.n662 585
R505 B.n661 B.n48 585
R506 B.n660 B.n659 585
R507 B.n658 B.n49 585
R508 B.n657 B.n656 585
R509 B.n655 B.n53 585
R510 B.n654 B.n653 585
R511 B.n652 B.n54 585
R512 B.n651 B.n650 585
R513 B.n649 B.n55 585
R514 B.n648 B.n647 585
R515 B.n646 B.n56 585
R516 B.n644 B.n643 585
R517 B.n642 B.n59 585
R518 B.n641 B.n640 585
R519 B.n639 B.n60 585
R520 B.n638 B.n637 585
R521 B.n636 B.n61 585
R522 B.n635 B.n634 585
R523 B.n633 B.n62 585
R524 B.n632 B.n631 585
R525 B.n630 B.n63 585
R526 B.n629 B.n628 585
R527 B.n627 B.n64 585
R528 B.n626 B.n625 585
R529 B.n624 B.n65 585
R530 B.n623 B.n622 585
R531 B.n621 B.n66 585
R532 B.n620 B.n619 585
R533 B.n618 B.n67 585
R534 B.n617 B.n616 585
R535 B.n615 B.n68 585
R536 B.n614 B.n613 585
R537 B.n612 B.n69 585
R538 B.n611 B.n610 585
R539 B.n609 B.n70 585
R540 B.n608 B.n607 585
R541 B.n606 B.n71 585
R542 B.n605 B.n604 585
R543 B.n603 B.n72 585
R544 B.n602 B.n601 585
R545 B.n600 B.n73 585
R546 B.n599 B.n598 585
R547 B.n597 B.n74 585
R548 B.n596 B.n595 585
R549 B.n594 B.n75 585
R550 B.n593 B.n592 585
R551 B.n591 B.n76 585
R552 B.n590 B.n589 585
R553 B.n588 B.n77 585
R554 B.n587 B.n586 585
R555 B.n585 B.n78 585
R556 B.n584 B.n583 585
R557 B.n582 B.n79 585
R558 B.n581 B.n580 585
R559 B.n579 B.n80 585
R560 B.n578 B.n577 585
R561 B.n576 B.n81 585
R562 B.n575 B.n574 585
R563 B.n573 B.n82 585
R564 B.n572 B.n571 585
R565 B.n570 B.n83 585
R566 B.n569 B.n568 585
R567 B.n567 B.n84 585
R568 B.n566 B.n565 585
R569 B.n564 B.n85 585
R570 B.n563 B.n562 585
R571 B.n561 B.n86 585
R572 B.n560 B.n559 585
R573 B.n747 B.n746 585
R574 B.n748 B.n19 585
R575 B.n750 B.n749 585
R576 B.n751 B.n18 585
R577 B.n753 B.n752 585
R578 B.n754 B.n17 585
R579 B.n756 B.n755 585
R580 B.n757 B.n16 585
R581 B.n759 B.n758 585
R582 B.n760 B.n15 585
R583 B.n762 B.n761 585
R584 B.n763 B.n14 585
R585 B.n765 B.n764 585
R586 B.n766 B.n13 585
R587 B.n768 B.n767 585
R588 B.n769 B.n12 585
R589 B.n771 B.n770 585
R590 B.n772 B.n11 585
R591 B.n774 B.n773 585
R592 B.n775 B.n10 585
R593 B.n777 B.n776 585
R594 B.n778 B.n9 585
R595 B.n780 B.n779 585
R596 B.n781 B.n8 585
R597 B.n783 B.n782 585
R598 B.n784 B.n7 585
R599 B.n786 B.n785 585
R600 B.n787 B.n6 585
R601 B.n789 B.n788 585
R602 B.n790 B.n5 585
R603 B.n792 B.n791 585
R604 B.n793 B.n4 585
R605 B.n795 B.n794 585
R606 B.n796 B.n3 585
R607 B.n798 B.n797 585
R608 B.n799 B.n0 585
R609 B.n2 B.n1 585
R610 B.n206 B.n205 585
R611 B.n208 B.n207 585
R612 B.n209 B.n204 585
R613 B.n211 B.n210 585
R614 B.n212 B.n203 585
R615 B.n214 B.n213 585
R616 B.n215 B.n202 585
R617 B.n217 B.n216 585
R618 B.n218 B.n201 585
R619 B.n220 B.n219 585
R620 B.n221 B.n200 585
R621 B.n223 B.n222 585
R622 B.n224 B.n199 585
R623 B.n226 B.n225 585
R624 B.n227 B.n198 585
R625 B.n229 B.n228 585
R626 B.n230 B.n197 585
R627 B.n232 B.n231 585
R628 B.n233 B.n196 585
R629 B.n235 B.n234 585
R630 B.n236 B.n195 585
R631 B.n238 B.n237 585
R632 B.n239 B.n194 585
R633 B.n241 B.n240 585
R634 B.n242 B.n193 585
R635 B.n244 B.n243 585
R636 B.n245 B.n192 585
R637 B.n247 B.n246 585
R638 B.n248 B.n191 585
R639 B.n250 B.n249 585
R640 B.n251 B.n190 585
R641 B.n253 B.n252 585
R642 B.n254 B.n189 585
R643 B.n256 B.n255 585
R644 B.n257 B.n188 585
R645 B.n342 B.t9 526.644
R646 B.n153 B.t3 526.644
R647 B.n57 B.t0 526.644
R648 B.n50 B.t6 526.644
R649 B.n259 B.n188 502.111
R650 B.n449 B.n124 502.111
R651 B.n559 B.n558 502.111
R652 B.n746 B.n745 502.111
R653 B.n801 B.n800 256.663
R654 B.n800 B.n799 235.042
R655 B.n800 B.n2 235.042
R656 B.n260 B.n259 163.367
R657 B.n261 B.n260 163.367
R658 B.n261 B.n186 163.367
R659 B.n265 B.n186 163.367
R660 B.n266 B.n265 163.367
R661 B.n267 B.n266 163.367
R662 B.n267 B.n184 163.367
R663 B.n271 B.n184 163.367
R664 B.n272 B.n271 163.367
R665 B.n273 B.n272 163.367
R666 B.n273 B.n182 163.367
R667 B.n277 B.n182 163.367
R668 B.n278 B.n277 163.367
R669 B.n279 B.n278 163.367
R670 B.n279 B.n180 163.367
R671 B.n283 B.n180 163.367
R672 B.n284 B.n283 163.367
R673 B.n285 B.n284 163.367
R674 B.n285 B.n178 163.367
R675 B.n289 B.n178 163.367
R676 B.n290 B.n289 163.367
R677 B.n291 B.n290 163.367
R678 B.n291 B.n176 163.367
R679 B.n295 B.n176 163.367
R680 B.n296 B.n295 163.367
R681 B.n297 B.n296 163.367
R682 B.n297 B.n174 163.367
R683 B.n301 B.n174 163.367
R684 B.n302 B.n301 163.367
R685 B.n303 B.n302 163.367
R686 B.n303 B.n172 163.367
R687 B.n307 B.n172 163.367
R688 B.n308 B.n307 163.367
R689 B.n309 B.n308 163.367
R690 B.n309 B.n170 163.367
R691 B.n313 B.n170 163.367
R692 B.n314 B.n313 163.367
R693 B.n315 B.n314 163.367
R694 B.n315 B.n168 163.367
R695 B.n319 B.n168 163.367
R696 B.n320 B.n319 163.367
R697 B.n321 B.n320 163.367
R698 B.n321 B.n166 163.367
R699 B.n325 B.n166 163.367
R700 B.n326 B.n325 163.367
R701 B.n327 B.n326 163.367
R702 B.n327 B.n164 163.367
R703 B.n331 B.n164 163.367
R704 B.n332 B.n331 163.367
R705 B.n333 B.n332 163.367
R706 B.n333 B.n162 163.367
R707 B.n337 B.n162 163.367
R708 B.n338 B.n337 163.367
R709 B.n339 B.n338 163.367
R710 B.n339 B.n160 163.367
R711 B.n346 B.n160 163.367
R712 B.n347 B.n346 163.367
R713 B.n348 B.n347 163.367
R714 B.n348 B.n158 163.367
R715 B.n352 B.n158 163.367
R716 B.n353 B.n352 163.367
R717 B.n354 B.n353 163.367
R718 B.n354 B.n156 163.367
R719 B.n358 B.n156 163.367
R720 B.n359 B.n358 163.367
R721 B.n360 B.n359 163.367
R722 B.n360 B.n152 163.367
R723 B.n365 B.n152 163.367
R724 B.n366 B.n365 163.367
R725 B.n367 B.n366 163.367
R726 B.n367 B.n150 163.367
R727 B.n371 B.n150 163.367
R728 B.n372 B.n371 163.367
R729 B.n373 B.n372 163.367
R730 B.n373 B.n148 163.367
R731 B.n377 B.n148 163.367
R732 B.n378 B.n377 163.367
R733 B.n379 B.n378 163.367
R734 B.n379 B.n146 163.367
R735 B.n383 B.n146 163.367
R736 B.n384 B.n383 163.367
R737 B.n385 B.n384 163.367
R738 B.n385 B.n144 163.367
R739 B.n389 B.n144 163.367
R740 B.n390 B.n389 163.367
R741 B.n391 B.n390 163.367
R742 B.n391 B.n142 163.367
R743 B.n395 B.n142 163.367
R744 B.n396 B.n395 163.367
R745 B.n397 B.n396 163.367
R746 B.n397 B.n140 163.367
R747 B.n401 B.n140 163.367
R748 B.n402 B.n401 163.367
R749 B.n403 B.n402 163.367
R750 B.n403 B.n138 163.367
R751 B.n407 B.n138 163.367
R752 B.n408 B.n407 163.367
R753 B.n409 B.n408 163.367
R754 B.n409 B.n136 163.367
R755 B.n413 B.n136 163.367
R756 B.n414 B.n413 163.367
R757 B.n415 B.n414 163.367
R758 B.n415 B.n134 163.367
R759 B.n419 B.n134 163.367
R760 B.n420 B.n419 163.367
R761 B.n421 B.n420 163.367
R762 B.n421 B.n132 163.367
R763 B.n425 B.n132 163.367
R764 B.n426 B.n425 163.367
R765 B.n427 B.n426 163.367
R766 B.n427 B.n130 163.367
R767 B.n431 B.n130 163.367
R768 B.n432 B.n431 163.367
R769 B.n433 B.n432 163.367
R770 B.n433 B.n128 163.367
R771 B.n437 B.n128 163.367
R772 B.n438 B.n437 163.367
R773 B.n439 B.n438 163.367
R774 B.n439 B.n126 163.367
R775 B.n443 B.n126 163.367
R776 B.n444 B.n443 163.367
R777 B.n445 B.n444 163.367
R778 B.n445 B.n124 163.367
R779 B.n558 B.n557 163.367
R780 B.n557 B.n88 163.367
R781 B.n553 B.n88 163.367
R782 B.n553 B.n552 163.367
R783 B.n552 B.n551 163.367
R784 B.n551 B.n90 163.367
R785 B.n547 B.n90 163.367
R786 B.n547 B.n546 163.367
R787 B.n546 B.n545 163.367
R788 B.n545 B.n92 163.367
R789 B.n541 B.n92 163.367
R790 B.n541 B.n540 163.367
R791 B.n540 B.n539 163.367
R792 B.n539 B.n94 163.367
R793 B.n535 B.n94 163.367
R794 B.n535 B.n534 163.367
R795 B.n534 B.n533 163.367
R796 B.n533 B.n96 163.367
R797 B.n529 B.n96 163.367
R798 B.n529 B.n528 163.367
R799 B.n528 B.n527 163.367
R800 B.n527 B.n98 163.367
R801 B.n523 B.n98 163.367
R802 B.n523 B.n522 163.367
R803 B.n522 B.n521 163.367
R804 B.n521 B.n100 163.367
R805 B.n517 B.n100 163.367
R806 B.n517 B.n516 163.367
R807 B.n516 B.n515 163.367
R808 B.n515 B.n102 163.367
R809 B.n511 B.n102 163.367
R810 B.n511 B.n510 163.367
R811 B.n510 B.n509 163.367
R812 B.n509 B.n104 163.367
R813 B.n505 B.n104 163.367
R814 B.n505 B.n504 163.367
R815 B.n504 B.n503 163.367
R816 B.n503 B.n106 163.367
R817 B.n499 B.n106 163.367
R818 B.n499 B.n498 163.367
R819 B.n498 B.n497 163.367
R820 B.n497 B.n108 163.367
R821 B.n493 B.n108 163.367
R822 B.n493 B.n492 163.367
R823 B.n492 B.n491 163.367
R824 B.n491 B.n110 163.367
R825 B.n487 B.n110 163.367
R826 B.n487 B.n486 163.367
R827 B.n486 B.n485 163.367
R828 B.n485 B.n112 163.367
R829 B.n481 B.n112 163.367
R830 B.n481 B.n480 163.367
R831 B.n480 B.n479 163.367
R832 B.n479 B.n114 163.367
R833 B.n475 B.n114 163.367
R834 B.n475 B.n474 163.367
R835 B.n474 B.n473 163.367
R836 B.n473 B.n116 163.367
R837 B.n469 B.n116 163.367
R838 B.n469 B.n468 163.367
R839 B.n468 B.n467 163.367
R840 B.n467 B.n118 163.367
R841 B.n463 B.n118 163.367
R842 B.n463 B.n462 163.367
R843 B.n462 B.n461 163.367
R844 B.n461 B.n120 163.367
R845 B.n457 B.n120 163.367
R846 B.n457 B.n456 163.367
R847 B.n456 B.n455 163.367
R848 B.n455 B.n122 163.367
R849 B.n451 B.n122 163.367
R850 B.n451 B.n450 163.367
R851 B.n450 B.n449 163.367
R852 B.n745 B.n744 163.367
R853 B.n744 B.n21 163.367
R854 B.n740 B.n21 163.367
R855 B.n740 B.n739 163.367
R856 B.n739 B.n738 163.367
R857 B.n738 B.n23 163.367
R858 B.n734 B.n23 163.367
R859 B.n734 B.n733 163.367
R860 B.n733 B.n732 163.367
R861 B.n732 B.n25 163.367
R862 B.n728 B.n25 163.367
R863 B.n728 B.n727 163.367
R864 B.n727 B.n726 163.367
R865 B.n726 B.n27 163.367
R866 B.n722 B.n27 163.367
R867 B.n722 B.n721 163.367
R868 B.n721 B.n720 163.367
R869 B.n720 B.n29 163.367
R870 B.n716 B.n29 163.367
R871 B.n716 B.n715 163.367
R872 B.n715 B.n714 163.367
R873 B.n714 B.n31 163.367
R874 B.n710 B.n31 163.367
R875 B.n710 B.n709 163.367
R876 B.n709 B.n708 163.367
R877 B.n708 B.n33 163.367
R878 B.n704 B.n33 163.367
R879 B.n704 B.n703 163.367
R880 B.n703 B.n702 163.367
R881 B.n702 B.n35 163.367
R882 B.n698 B.n35 163.367
R883 B.n698 B.n697 163.367
R884 B.n697 B.n696 163.367
R885 B.n696 B.n37 163.367
R886 B.n692 B.n37 163.367
R887 B.n692 B.n691 163.367
R888 B.n691 B.n690 163.367
R889 B.n690 B.n39 163.367
R890 B.n686 B.n39 163.367
R891 B.n686 B.n685 163.367
R892 B.n685 B.n684 163.367
R893 B.n684 B.n41 163.367
R894 B.n680 B.n41 163.367
R895 B.n680 B.n679 163.367
R896 B.n679 B.n678 163.367
R897 B.n678 B.n43 163.367
R898 B.n674 B.n43 163.367
R899 B.n674 B.n673 163.367
R900 B.n673 B.n672 163.367
R901 B.n672 B.n45 163.367
R902 B.n668 B.n45 163.367
R903 B.n668 B.n667 163.367
R904 B.n667 B.n666 163.367
R905 B.n666 B.n47 163.367
R906 B.n662 B.n47 163.367
R907 B.n662 B.n661 163.367
R908 B.n661 B.n660 163.367
R909 B.n660 B.n49 163.367
R910 B.n656 B.n49 163.367
R911 B.n656 B.n655 163.367
R912 B.n655 B.n654 163.367
R913 B.n654 B.n54 163.367
R914 B.n650 B.n54 163.367
R915 B.n650 B.n649 163.367
R916 B.n649 B.n648 163.367
R917 B.n648 B.n56 163.367
R918 B.n643 B.n56 163.367
R919 B.n643 B.n642 163.367
R920 B.n642 B.n641 163.367
R921 B.n641 B.n60 163.367
R922 B.n637 B.n60 163.367
R923 B.n637 B.n636 163.367
R924 B.n636 B.n635 163.367
R925 B.n635 B.n62 163.367
R926 B.n631 B.n62 163.367
R927 B.n631 B.n630 163.367
R928 B.n630 B.n629 163.367
R929 B.n629 B.n64 163.367
R930 B.n625 B.n64 163.367
R931 B.n625 B.n624 163.367
R932 B.n624 B.n623 163.367
R933 B.n623 B.n66 163.367
R934 B.n619 B.n66 163.367
R935 B.n619 B.n618 163.367
R936 B.n618 B.n617 163.367
R937 B.n617 B.n68 163.367
R938 B.n613 B.n68 163.367
R939 B.n613 B.n612 163.367
R940 B.n612 B.n611 163.367
R941 B.n611 B.n70 163.367
R942 B.n607 B.n70 163.367
R943 B.n607 B.n606 163.367
R944 B.n606 B.n605 163.367
R945 B.n605 B.n72 163.367
R946 B.n601 B.n72 163.367
R947 B.n601 B.n600 163.367
R948 B.n600 B.n599 163.367
R949 B.n599 B.n74 163.367
R950 B.n595 B.n74 163.367
R951 B.n595 B.n594 163.367
R952 B.n594 B.n593 163.367
R953 B.n593 B.n76 163.367
R954 B.n589 B.n76 163.367
R955 B.n589 B.n588 163.367
R956 B.n588 B.n587 163.367
R957 B.n587 B.n78 163.367
R958 B.n583 B.n78 163.367
R959 B.n583 B.n582 163.367
R960 B.n582 B.n581 163.367
R961 B.n581 B.n80 163.367
R962 B.n577 B.n80 163.367
R963 B.n577 B.n576 163.367
R964 B.n576 B.n575 163.367
R965 B.n575 B.n82 163.367
R966 B.n571 B.n82 163.367
R967 B.n571 B.n570 163.367
R968 B.n570 B.n569 163.367
R969 B.n569 B.n84 163.367
R970 B.n565 B.n84 163.367
R971 B.n565 B.n564 163.367
R972 B.n564 B.n563 163.367
R973 B.n563 B.n86 163.367
R974 B.n559 B.n86 163.367
R975 B.n746 B.n19 163.367
R976 B.n750 B.n19 163.367
R977 B.n751 B.n750 163.367
R978 B.n752 B.n751 163.367
R979 B.n752 B.n17 163.367
R980 B.n756 B.n17 163.367
R981 B.n757 B.n756 163.367
R982 B.n758 B.n757 163.367
R983 B.n758 B.n15 163.367
R984 B.n762 B.n15 163.367
R985 B.n763 B.n762 163.367
R986 B.n764 B.n763 163.367
R987 B.n764 B.n13 163.367
R988 B.n768 B.n13 163.367
R989 B.n769 B.n768 163.367
R990 B.n770 B.n769 163.367
R991 B.n770 B.n11 163.367
R992 B.n774 B.n11 163.367
R993 B.n775 B.n774 163.367
R994 B.n776 B.n775 163.367
R995 B.n776 B.n9 163.367
R996 B.n780 B.n9 163.367
R997 B.n781 B.n780 163.367
R998 B.n782 B.n781 163.367
R999 B.n782 B.n7 163.367
R1000 B.n786 B.n7 163.367
R1001 B.n787 B.n786 163.367
R1002 B.n788 B.n787 163.367
R1003 B.n788 B.n5 163.367
R1004 B.n792 B.n5 163.367
R1005 B.n793 B.n792 163.367
R1006 B.n794 B.n793 163.367
R1007 B.n794 B.n3 163.367
R1008 B.n798 B.n3 163.367
R1009 B.n799 B.n798 163.367
R1010 B.n206 B.n2 163.367
R1011 B.n207 B.n206 163.367
R1012 B.n207 B.n204 163.367
R1013 B.n211 B.n204 163.367
R1014 B.n212 B.n211 163.367
R1015 B.n213 B.n212 163.367
R1016 B.n213 B.n202 163.367
R1017 B.n217 B.n202 163.367
R1018 B.n218 B.n217 163.367
R1019 B.n219 B.n218 163.367
R1020 B.n219 B.n200 163.367
R1021 B.n223 B.n200 163.367
R1022 B.n224 B.n223 163.367
R1023 B.n225 B.n224 163.367
R1024 B.n225 B.n198 163.367
R1025 B.n229 B.n198 163.367
R1026 B.n230 B.n229 163.367
R1027 B.n231 B.n230 163.367
R1028 B.n231 B.n196 163.367
R1029 B.n235 B.n196 163.367
R1030 B.n236 B.n235 163.367
R1031 B.n237 B.n236 163.367
R1032 B.n237 B.n194 163.367
R1033 B.n241 B.n194 163.367
R1034 B.n242 B.n241 163.367
R1035 B.n243 B.n242 163.367
R1036 B.n243 B.n192 163.367
R1037 B.n247 B.n192 163.367
R1038 B.n248 B.n247 163.367
R1039 B.n249 B.n248 163.367
R1040 B.n249 B.n190 163.367
R1041 B.n253 B.n190 163.367
R1042 B.n254 B.n253 163.367
R1043 B.n255 B.n254 163.367
R1044 B.n255 B.n188 163.367
R1045 B.n153 B.t4 142.356
R1046 B.n57 B.t2 142.356
R1047 B.n342 B.t10 142.333
R1048 B.n50 B.t8 142.333
R1049 B.n154 B.t5 110.936
R1050 B.n58 B.t1 110.936
R1051 B.n343 B.t11 110.915
R1052 B.n51 B.t7 110.915
R1053 B.n344 B.n343 59.5399
R1054 B.n362 B.n154 59.5399
R1055 B.n645 B.n58 59.5399
R1056 B.n52 B.n51 59.5399
R1057 B.n747 B.n20 32.6249
R1058 B.n560 B.n87 32.6249
R1059 B.n448 B.n447 32.6249
R1060 B.n258 B.n257 32.6249
R1061 B.n343 B.n342 31.4187
R1062 B.n154 B.n153 31.4187
R1063 B.n58 B.n57 31.4187
R1064 B.n51 B.n50 31.4187
R1065 B B.n801 18.0485
R1066 B.n748 B.n747 10.6151
R1067 B.n749 B.n748 10.6151
R1068 B.n749 B.n18 10.6151
R1069 B.n753 B.n18 10.6151
R1070 B.n754 B.n753 10.6151
R1071 B.n755 B.n754 10.6151
R1072 B.n755 B.n16 10.6151
R1073 B.n759 B.n16 10.6151
R1074 B.n760 B.n759 10.6151
R1075 B.n761 B.n760 10.6151
R1076 B.n761 B.n14 10.6151
R1077 B.n765 B.n14 10.6151
R1078 B.n766 B.n765 10.6151
R1079 B.n767 B.n766 10.6151
R1080 B.n767 B.n12 10.6151
R1081 B.n771 B.n12 10.6151
R1082 B.n772 B.n771 10.6151
R1083 B.n773 B.n772 10.6151
R1084 B.n773 B.n10 10.6151
R1085 B.n777 B.n10 10.6151
R1086 B.n778 B.n777 10.6151
R1087 B.n779 B.n778 10.6151
R1088 B.n779 B.n8 10.6151
R1089 B.n783 B.n8 10.6151
R1090 B.n784 B.n783 10.6151
R1091 B.n785 B.n784 10.6151
R1092 B.n785 B.n6 10.6151
R1093 B.n789 B.n6 10.6151
R1094 B.n790 B.n789 10.6151
R1095 B.n791 B.n790 10.6151
R1096 B.n791 B.n4 10.6151
R1097 B.n795 B.n4 10.6151
R1098 B.n796 B.n795 10.6151
R1099 B.n797 B.n796 10.6151
R1100 B.n797 B.n0 10.6151
R1101 B.n743 B.n20 10.6151
R1102 B.n743 B.n742 10.6151
R1103 B.n742 B.n741 10.6151
R1104 B.n741 B.n22 10.6151
R1105 B.n737 B.n22 10.6151
R1106 B.n737 B.n736 10.6151
R1107 B.n736 B.n735 10.6151
R1108 B.n735 B.n24 10.6151
R1109 B.n731 B.n24 10.6151
R1110 B.n731 B.n730 10.6151
R1111 B.n730 B.n729 10.6151
R1112 B.n729 B.n26 10.6151
R1113 B.n725 B.n26 10.6151
R1114 B.n725 B.n724 10.6151
R1115 B.n724 B.n723 10.6151
R1116 B.n723 B.n28 10.6151
R1117 B.n719 B.n28 10.6151
R1118 B.n719 B.n718 10.6151
R1119 B.n718 B.n717 10.6151
R1120 B.n717 B.n30 10.6151
R1121 B.n713 B.n30 10.6151
R1122 B.n713 B.n712 10.6151
R1123 B.n712 B.n711 10.6151
R1124 B.n711 B.n32 10.6151
R1125 B.n707 B.n32 10.6151
R1126 B.n707 B.n706 10.6151
R1127 B.n706 B.n705 10.6151
R1128 B.n705 B.n34 10.6151
R1129 B.n701 B.n34 10.6151
R1130 B.n701 B.n700 10.6151
R1131 B.n700 B.n699 10.6151
R1132 B.n699 B.n36 10.6151
R1133 B.n695 B.n36 10.6151
R1134 B.n695 B.n694 10.6151
R1135 B.n694 B.n693 10.6151
R1136 B.n693 B.n38 10.6151
R1137 B.n689 B.n38 10.6151
R1138 B.n689 B.n688 10.6151
R1139 B.n688 B.n687 10.6151
R1140 B.n687 B.n40 10.6151
R1141 B.n683 B.n40 10.6151
R1142 B.n683 B.n682 10.6151
R1143 B.n682 B.n681 10.6151
R1144 B.n681 B.n42 10.6151
R1145 B.n677 B.n42 10.6151
R1146 B.n677 B.n676 10.6151
R1147 B.n676 B.n675 10.6151
R1148 B.n675 B.n44 10.6151
R1149 B.n671 B.n44 10.6151
R1150 B.n671 B.n670 10.6151
R1151 B.n670 B.n669 10.6151
R1152 B.n669 B.n46 10.6151
R1153 B.n665 B.n46 10.6151
R1154 B.n665 B.n664 10.6151
R1155 B.n664 B.n663 10.6151
R1156 B.n663 B.n48 10.6151
R1157 B.n659 B.n658 10.6151
R1158 B.n658 B.n657 10.6151
R1159 B.n657 B.n53 10.6151
R1160 B.n653 B.n53 10.6151
R1161 B.n653 B.n652 10.6151
R1162 B.n652 B.n651 10.6151
R1163 B.n651 B.n55 10.6151
R1164 B.n647 B.n55 10.6151
R1165 B.n647 B.n646 10.6151
R1166 B.n644 B.n59 10.6151
R1167 B.n640 B.n59 10.6151
R1168 B.n640 B.n639 10.6151
R1169 B.n639 B.n638 10.6151
R1170 B.n638 B.n61 10.6151
R1171 B.n634 B.n61 10.6151
R1172 B.n634 B.n633 10.6151
R1173 B.n633 B.n632 10.6151
R1174 B.n632 B.n63 10.6151
R1175 B.n628 B.n63 10.6151
R1176 B.n628 B.n627 10.6151
R1177 B.n627 B.n626 10.6151
R1178 B.n626 B.n65 10.6151
R1179 B.n622 B.n65 10.6151
R1180 B.n622 B.n621 10.6151
R1181 B.n621 B.n620 10.6151
R1182 B.n620 B.n67 10.6151
R1183 B.n616 B.n67 10.6151
R1184 B.n616 B.n615 10.6151
R1185 B.n615 B.n614 10.6151
R1186 B.n614 B.n69 10.6151
R1187 B.n610 B.n69 10.6151
R1188 B.n610 B.n609 10.6151
R1189 B.n609 B.n608 10.6151
R1190 B.n608 B.n71 10.6151
R1191 B.n604 B.n71 10.6151
R1192 B.n604 B.n603 10.6151
R1193 B.n603 B.n602 10.6151
R1194 B.n602 B.n73 10.6151
R1195 B.n598 B.n73 10.6151
R1196 B.n598 B.n597 10.6151
R1197 B.n597 B.n596 10.6151
R1198 B.n596 B.n75 10.6151
R1199 B.n592 B.n75 10.6151
R1200 B.n592 B.n591 10.6151
R1201 B.n591 B.n590 10.6151
R1202 B.n590 B.n77 10.6151
R1203 B.n586 B.n77 10.6151
R1204 B.n586 B.n585 10.6151
R1205 B.n585 B.n584 10.6151
R1206 B.n584 B.n79 10.6151
R1207 B.n580 B.n79 10.6151
R1208 B.n580 B.n579 10.6151
R1209 B.n579 B.n578 10.6151
R1210 B.n578 B.n81 10.6151
R1211 B.n574 B.n81 10.6151
R1212 B.n574 B.n573 10.6151
R1213 B.n573 B.n572 10.6151
R1214 B.n572 B.n83 10.6151
R1215 B.n568 B.n83 10.6151
R1216 B.n568 B.n567 10.6151
R1217 B.n567 B.n566 10.6151
R1218 B.n566 B.n85 10.6151
R1219 B.n562 B.n85 10.6151
R1220 B.n562 B.n561 10.6151
R1221 B.n561 B.n560 10.6151
R1222 B.n556 B.n87 10.6151
R1223 B.n556 B.n555 10.6151
R1224 B.n555 B.n554 10.6151
R1225 B.n554 B.n89 10.6151
R1226 B.n550 B.n89 10.6151
R1227 B.n550 B.n549 10.6151
R1228 B.n549 B.n548 10.6151
R1229 B.n548 B.n91 10.6151
R1230 B.n544 B.n91 10.6151
R1231 B.n544 B.n543 10.6151
R1232 B.n543 B.n542 10.6151
R1233 B.n542 B.n93 10.6151
R1234 B.n538 B.n93 10.6151
R1235 B.n538 B.n537 10.6151
R1236 B.n537 B.n536 10.6151
R1237 B.n536 B.n95 10.6151
R1238 B.n532 B.n95 10.6151
R1239 B.n532 B.n531 10.6151
R1240 B.n531 B.n530 10.6151
R1241 B.n530 B.n97 10.6151
R1242 B.n526 B.n97 10.6151
R1243 B.n526 B.n525 10.6151
R1244 B.n525 B.n524 10.6151
R1245 B.n524 B.n99 10.6151
R1246 B.n520 B.n99 10.6151
R1247 B.n520 B.n519 10.6151
R1248 B.n519 B.n518 10.6151
R1249 B.n518 B.n101 10.6151
R1250 B.n514 B.n101 10.6151
R1251 B.n514 B.n513 10.6151
R1252 B.n513 B.n512 10.6151
R1253 B.n512 B.n103 10.6151
R1254 B.n508 B.n103 10.6151
R1255 B.n508 B.n507 10.6151
R1256 B.n507 B.n506 10.6151
R1257 B.n506 B.n105 10.6151
R1258 B.n502 B.n105 10.6151
R1259 B.n502 B.n501 10.6151
R1260 B.n501 B.n500 10.6151
R1261 B.n500 B.n107 10.6151
R1262 B.n496 B.n107 10.6151
R1263 B.n496 B.n495 10.6151
R1264 B.n495 B.n494 10.6151
R1265 B.n494 B.n109 10.6151
R1266 B.n490 B.n109 10.6151
R1267 B.n490 B.n489 10.6151
R1268 B.n489 B.n488 10.6151
R1269 B.n488 B.n111 10.6151
R1270 B.n484 B.n111 10.6151
R1271 B.n484 B.n483 10.6151
R1272 B.n483 B.n482 10.6151
R1273 B.n482 B.n113 10.6151
R1274 B.n478 B.n113 10.6151
R1275 B.n478 B.n477 10.6151
R1276 B.n477 B.n476 10.6151
R1277 B.n476 B.n115 10.6151
R1278 B.n472 B.n115 10.6151
R1279 B.n472 B.n471 10.6151
R1280 B.n471 B.n470 10.6151
R1281 B.n470 B.n117 10.6151
R1282 B.n466 B.n117 10.6151
R1283 B.n466 B.n465 10.6151
R1284 B.n465 B.n464 10.6151
R1285 B.n464 B.n119 10.6151
R1286 B.n460 B.n119 10.6151
R1287 B.n460 B.n459 10.6151
R1288 B.n459 B.n458 10.6151
R1289 B.n458 B.n121 10.6151
R1290 B.n454 B.n121 10.6151
R1291 B.n454 B.n453 10.6151
R1292 B.n453 B.n452 10.6151
R1293 B.n452 B.n123 10.6151
R1294 B.n448 B.n123 10.6151
R1295 B.n205 B.n1 10.6151
R1296 B.n208 B.n205 10.6151
R1297 B.n209 B.n208 10.6151
R1298 B.n210 B.n209 10.6151
R1299 B.n210 B.n203 10.6151
R1300 B.n214 B.n203 10.6151
R1301 B.n215 B.n214 10.6151
R1302 B.n216 B.n215 10.6151
R1303 B.n216 B.n201 10.6151
R1304 B.n220 B.n201 10.6151
R1305 B.n221 B.n220 10.6151
R1306 B.n222 B.n221 10.6151
R1307 B.n222 B.n199 10.6151
R1308 B.n226 B.n199 10.6151
R1309 B.n227 B.n226 10.6151
R1310 B.n228 B.n227 10.6151
R1311 B.n228 B.n197 10.6151
R1312 B.n232 B.n197 10.6151
R1313 B.n233 B.n232 10.6151
R1314 B.n234 B.n233 10.6151
R1315 B.n234 B.n195 10.6151
R1316 B.n238 B.n195 10.6151
R1317 B.n239 B.n238 10.6151
R1318 B.n240 B.n239 10.6151
R1319 B.n240 B.n193 10.6151
R1320 B.n244 B.n193 10.6151
R1321 B.n245 B.n244 10.6151
R1322 B.n246 B.n245 10.6151
R1323 B.n246 B.n191 10.6151
R1324 B.n250 B.n191 10.6151
R1325 B.n251 B.n250 10.6151
R1326 B.n252 B.n251 10.6151
R1327 B.n252 B.n189 10.6151
R1328 B.n256 B.n189 10.6151
R1329 B.n257 B.n256 10.6151
R1330 B.n258 B.n187 10.6151
R1331 B.n262 B.n187 10.6151
R1332 B.n263 B.n262 10.6151
R1333 B.n264 B.n263 10.6151
R1334 B.n264 B.n185 10.6151
R1335 B.n268 B.n185 10.6151
R1336 B.n269 B.n268 10.6151
R1337 B.n270 B.n269 10.6151
R1338 B.n270 B.n183 10.6151
R1339 B.n274 B.n183 10.6151
R1340 B.n275 B.n274 10.6151
R1341 B.n276 B.n275 10.6151
R1342 B.n276 B.n181 10.6151
R1343 B.n280 B.n181 10.6151
R1344 B.n281 B.n280 10.6151
R1345 B.n282 B.n281 10.6151
R1346 B.n282 B.n179 10.6151
R1347 B.n286 B.n179 10.6151
R1348 B.n287 B.n286 10.6151
R1349 B.n288 B.n287 10.6151
R1350 B.n288 B.n177 10.6151
R1351 B.n292 B.n177 10.6151
R1352 B.n293 B.n292 10.6151
R1353 B.n294 B.n293 10.6151
R1354 B.n294 B.n175 10.6151
R1355 B.n298 B.n175 10.6151
R1356 B.n299 B.n298 10.6151
R1357 B.n300 B.n299 10.6151
R1358 B.n300 B.n173 10.6151
R1359 B.n304 B.n173 10.6151
R1360 B.n305 B.n304 10.6151
R1361 B.n306 B.n305 10.6151
R1362 B.n306 B.n171 10.6151
R1363 B.n310 B.n171 10.6151
R1364 B.n311 B.n310 10.6151
R1365 B.n312 B.n311 10.6151
R1366 B.n312 B.n169 10.6151
R1367 B.n316 B.n169 10.6151
R1368 B.n317 B.n316 10.6151
R1369 B.n318 B.n317 10.6151
R1370 B.n318 B.n167 10.6151
R1371 B.n322 B.n167 10.6151
R1372 B.n323 B.n322 10.6151
R1373 B.n324 B.n323 10.6151
R1374 B.n324 B.n165 10.6151
R1375 B.n328 B.n165 10.6151
R1376 B.n329 B.n328 10.6151
R1377 B.n330 B.n329 10.6151
R1378 B.n330 B.n163 10.6151
R1379 B.n334 B.n163 10.6151
R1380 B.n335 B.n334 10.6151
R1381 B.n336 B.n335 10.6151
R1382 B.n336 B.n161 10.6151
R1383 B.n340 B.n161 10.6151
R1384 B.n341 B.n340 10.6151
R1385 B.n345 B.n341 10.6151
R1386 B.n349 B.n159 10.6151
R1387 B.n350 B.n349 10.6151
R1388 B.n351 B.n350 10.6151
R1389 B.n351 B.n157 10.6151
R1390 B.n355 B.n157 10.6151
R1391 B.n356 B.n355 10.6151
R1392 B.n357 B.n356 10.6151
R1393 B.n357 B.n155 10.6151
R1394 B.n361 B.n155 10.6151
R1395 B.n364 B.n363 10.6151
R1396 B.n364 B.n151 10.6151
R1397 B.n368 B.n151 10.6151
R1398 B.n369 B.n368 10.6151
R1399 B.n370 B.n369 10.6151
R1400 B.n370 B.n149 10.6151
R1401 B.n374 B.n149 10.6151
R1402 B.n375 B.n374 10.6151
R1403 B.n376 B.n375 10.6151
R1404 B.n376 B.n147 10.6151
R1405 B.n380 B.n147 10.6151
R1406 B.n381 B.n380 10.6151
R1407 B.n382 B.n381 10.6151
R1408 B.n382 B.n145 10.6151
R1409 B.n386 B.n145 10.6151
R1410 B.n387 B.n386 10.6151
R1411 B.n388 B.n387 10.6151
R1412 B.n388 B.n143 10.6151
R1413 B.n392 B.n143 10.6151
R1414 B.n393 B.n392 10.6151
R1415 B.n394 B.n393 10.6151
R1416 B.n394 B.n141 10.6151
R1417 B.n398 B.n141 10.6151
R1418 B.n399 B.n398 10.6151
R1419 B.n400 B.n399 10.6151
R1420 B.n400 B.n139 10.6151
R1421 B.n404 B.n139 10.6151
R1422 B.n405 B.n404 10.6151
R1423 B.n406 B.n405 10.6151
R1424 B.n406 B.n137 10.6151
R1425 B.n410 B.n137 10.6151
R1426 B.n411 B.n410 10.6151
R1427 B.n412 B.n411 10.6151
R1428 B.n412 B.n135 10.6151
R1429 B.n416 B.n135 10.6151
R1430 B.n417 B.n416 10.6151
R1431 B.n418 B.n417 10.6151
R1432 B.n418 B.n133 10.6151
R1433 B.n422 B.n133 10.6151
R1434 B.n423 B.n422 10.6151
R1435 B.n424 B.n423 10.6151
R1436 B.n424 B.n131 10.6151
R1437 B.n428 B.n131 10.6151
R1438 B.n429 B.n428 10.6151
R1439 B.n430 B.n429 10.6151
R1440 B.n430 B.n129 10.6151
R1441 B.n434 B.n129 10.6151
R1442 B.n435 B.n434 10.6151
R1443 B.n436 B.n435 10.6151
R1444 B.n436 B.n127 10.6151
R1445 B.n440 B.n127 10.6151
R1446 B.n441 B.n440 10.6151
R1447 B.n442 B.n441 10.6151
R1448 B.n442 B.n125 10.6151
R1449 B.n446 B.n125 10.6151
R1450 B.n447 B.n446 10.6151
R1451 B.n52 B.n48 9.36635
R1452 B.n645 B.n644 9.36635
R1453 B.n345 B.n344 9.36635
R1454 B.n363 B.n362 9.36635
R1455 B.n801 B.n0 8.11757
R1456 B.n801 B.n1 8.11757
R1457 B.n659 B.n52 1.24928
R1458 B.n646 B.n645 1.24928
R1459 B.n344 B.n159 1.24928
R1460 B.n362 B.n361 1.24928
C0 VDD1 VTAIL 14.886401f
C1 VP VTAIL 12.333599f
C2 VN VTAIL 12.319f
C3 VDD2 VTAIL 14.9243f
C4 VDD1 B 2.35003f
C5 B VP 1.63799f
C6 B VN 1.01405f
C7 VDD2 B 2.41694f
C8 VDD1 w_n2914_n4416# 2.66266f
C9 VP w_n2914_n4416# 6.30442f
C10 B VTAIL 4.12934f
C11 w_n2914_n4416# VN 5.92908f
C12 VDD2 w_n2914_n4416# 2.73817f
C13 w_n2914_n4416# VTAIL 3.83402f
C14 VDD1 VP 12.6876f
C15 VDD1 VN 0.150658f
C16 VP VN 7.43493f
C17 VDD2 VDD1 1.33857f
C18 B w_n2914_n4416# 9.81283f
C19 VDD2 VP 0.41756f
C20 VDD2 VN 12.426299f
C21 VDD2 VSUBS 1.818583f
C22 VDD1 VSUBS 1.562246f
C23 VTAIL VSUBS 1.151576f
C24 VN VSUBS 5.95002f
C25 VP VSUBS 2.754188f
C26 B VSUBS 4.185533f
C27 w_n2914_n4416# VSUBS 0.157461p
C28 B.n0 VSUBS 0.007483f
C29 B.n1 VSUBS 0.007483f
C30 B.n2 VSUBS 0.011067f
C31 B.n3 VSUBS 0.008481f
C32 B.n4 VSUBS 0.008481f
C33 B.n5 VSUBS 0.008481f
C34 B.n6 VSUBS 0.008481f
C35 B.n7 VSUBS 0.008481f
C36 B.n8 VSUBS 0.008481f
C37 B.n9 VSUBS 0.008481f
C38 B.n10 VSUBS 0.008481f
C39 B.n11 VSUBS 0.008481f
C40 B.n12 VSUBS 0.008481f
C41 B.n13 VSUBS 0.008481f
C42 B.n14 VSUBS 0.008481f
C43 B.n15 VSUBS 0.008481f
C44 B.n16 VSUBS 0.008481f
C45 B.n17 VSUBS 0.008481f
C46 B.n18 VSUBS 0.008481f
C47 B.n19 VSUBS 0.008481f
C48 B.n20 VSUBS 0.020625f
C49 B.n21 VSUBS 0.008481f
C50 B.n22 VSUBS 0.008481f
C51 B.n23 VSUBS 0.008481f
C52 B.n24 VSUBS 0.008481f
C53 B.n25 VSUBS 0.008481f
C54 B.n26 VSUBS 0.008481f
C55 B.n27 VSUBS 0.008481f
C56 B.n28 VSUBS 0.008481f
C57 B.n29 VSUBS 0.008481f
C58 B.n30 VSUBS 0.008481f
C59 B.n31 VSUBS 0.008481f
C60 B.n32 VSUBS 0.008481f
C61 B.n33 VSUBS 0.008481f
C62 B.n34 VSUBS 0.008481f
C63 B.n35 VSUBS 0.008481f
C64 B.n36 VSUBS 0.008481f
C65 B.n37 VSUBS 0.008481f
C66 B.n38 VSUBS 0.008481f
C67 B.n39 VSUBS 0.008481f
C68 B.n40 VSUBS 0.008481f
C69 B.n41 VSUBS 0.008481f
C70 B.n42 VSUBS 0.008481f
C71 B.n43 VSUBS 0.008481f
C72 B.n44 VSUBS 0.008481f
C73 B.n45 VSUBS 0.008481f
C74 B.n46 VSUBS 0.008481f
C75 B.n47 VSUBS 0.008481f
C76 B.n48 VSUBS 0.007982f
C77 B.n49 VSUBS 0.008481f
C78 B.t7 VSUBS 0.702983f
C79 B.t8 VSUBS 0.718134f
C80 B.t6 VSUBS 1.13593f
C81 B.n50 VSUBS 0.293435f
C82 B.n51 VSUBS 0.080734f
C83 B.n52 VSUBS 0.019649f
C84 B.n53 VSUBS 0.008481f
C85 B.n54 VSUBS 0.008481f
C86 B.n55 VSUBS 0.008481f
C87 B.n56 VSUBS 0.008481f
C88 B.t1 VSUBS 0.702959f
C89 B.t2 VSUBS 0.718113f
C90 B.t0 VSUBS 1.13593f
C91 B.n57 VSUBS 0.293456f
C92 B.n58 VSUBS 0.080758f
C93 B.n59 VSUBS 0.008481f
C94 B.n60 VSUBS 0.008481f
C95 B.n61 VSUBS 0.008481f
C96 B.n62 VSUBS 0.008481f
C97 B.n63 VSUBS 0.008481f
C98 B.n64 VSUBS 0.008481f
C99 B.n65 VSUBS 0.008481f
C100 B.n66 VSUBS 0.008481f
C101 B.n67 VSUBS 0.008481f
C102 B.n68 VSUBS 0.008481f
C103 B.n69 VSUBS 0.008481f
C104 B.n70 VSUBS 0.008481f
C105 B.n71 VSUBS 0.008481f
C106 B.n72 VSUBS 0.008481f
C107 B.n73 VSUBS 0.008481f
C108 B.n74 VSUBS 0.008481f
C109 B.n75 VSUBS 0.008481f
C110 B.n76 VSUBS 0.008481f
C111 B.n77 VSUBS 0.008481f
C112 B.n78 VSUBS 0.008481f
C113 B.n79 VSUBS 0.008481f
C114 B.n80 VSUBS 0.008481f
C115 B.n81 VSUBS 0.008481f
C116 B.n82 VSUBS 0.008481f
C117 B.n83 VSUBS 0.008481f
C118 B.n84 VSUBS 0.008481f
C119 B.n85 VSUBS 0.008481f
C120 B.n86 VSUBS 0.008481f
C121 B.n87 VSUBS 0.019035f
C122 B.n88 VSUBS 0.008481f
C123 B.n89 VSUBS 0.008481f
C124 B.n90 VSUBS 0.008481f
C125 B.n91 VSUBS 0.008481f
C126 B.n92 VSUBS 0.008481f
C127 B.n93 VSUBS 0.008481f
C128 B.n94 VSUBS 0.008481f
C129 B.n95 VSUBS 0.008481f
C130 B.n96 VSUBS 0.008481f
C131 B.n97 VSUBS 0.008481f
C132 B.n98 VSUBS 0.008481f
C133 B.n99 VSUBS 0.008481f
C134 B.n100 VSUBS 0.008481f
C135 B.n101 VSUBS 0.008481f
C136 B.n102 VSUBS 0.008481f
C137 B.n103 VSUBS 0.008481f
C138 B.n104 VSUBS 0.008481f
C139 B.n105 VSUBS 0.008481f
C140 B.n106 VSUBS 0.008481f
C141 B.n107 VSUBS 0.008481f
C142 B.n108 VSUBS 0.008481f
C143 B.n109 VSUBS 0.008481f
C144 B.n110 VSUBS 0.008481f
C145 B.n111 VSUBS 0.008481f
C146 B.n112 VSUBS 0.008481f
C147 B.n113 VSUBS 0.008481f
C148 B.n114 VSUBS 0.008481f
C149 B.n115 VSUBS 0.008481f
C150 B.n116 VSUBS 0.008481f
C151 B.n117 VSUBS 0.008481f
C152 B.n118 VSUBS 0.008481f
C153 B.n119 VSUBS 0.008481f
C154 B.n120 VSUBS 0.008481f
C155 B.n121 VSUBS 0.008481f
C156 B.n122 VSUBS 0.008481f
C157 B.n123 VSUBS 0.008481f
C158 B.n124 VSUBS 0.020625f
C159 B.n125 VSUBS 0.008481f
C160 B.n126 VSUBS 0.008481f
C161 B.n127 VSUBS 0.008481f
C162 B.n128 VSUBS 0.008481f
C163 B.n129 VSUBS 0.008481f
C164 B.n130 VSUBS 0.008481f
C165 B.n131 VSUBS 0.008481f
C166 B.n132 VSUBS 0.008481f
C167 B.n133 VSUBS 0.008481f
C168 B.n134 VSUBS 0.008481f
C169 B.n135 VSUBS 0.008481f
C170 B.n136 VSUBS 0.008481f
C171 B.n137 VSUBS 0.008481f
C172 B.n138 VSUBS 0.008481f
C173 B.n139 VSUBS 0.008481f
C174 B.n140 VSUBS 0.008481f
C175 B.n141 VSUBS 0.008481f
C176 B.n142 VSUBS 0.008481f
C177 B.n143 VSUBS 0.008481f
C178 B.n144 VSUBS 0.008481f
C179 B.n145 VSUBS 0.008481f
C180 B.n146 VSUBS 0.008481f
C181 B.n147 VSUBS 0.008481f
C182 B.n148 VSUBS 0.008481f
C183 B.n149 VSUBS 0.008481f
C184 B.n150 VSUBS 0.008481f
C185 B.n151 VSUBS 0.008481f
C186 B.n152 VSUBS 0.008481f
C187 B.t5 VSUBS 0.702959f
C188 B.t4 VSUBS 0.718113f
C189 B.t3 VSUBS 1.13593f
C190 B.n153 VSUBS 0.293456f
C191 B.n154 VSUBS 0.080758f
C192 B.n155 VSUBS 0.008481f
C193 B.n156 VSUBS 0.008481f
C194 B.n157 VSUBS 0.008481f
C195 B.n158 VSUBS 0.008481f
C196 B.n159 VSUBS 0.004739f
C197 B.n160 VSUBS 0.008481f
C198 B.n161 VSUBS 0.008481f
C199 B.n162 VSUBS 0.008481f
C200 B.n163 VSUBS 0.008481f
C201 B.n164 VSUBS 0.008481f
C202 B.n165 VSUBS 0.008481f
C203 B.n166 VSUBS 0.008481f
C204 B.n167 VSUBS 0.008481f
C205 B.n168 VSUBS 0.008481f
C206 B.n169 VSUBS 0.008481f
C207 B.n170 VSUBS 0.008481f
C208 B.n171 VSUBS 0.008481f
C209 B.n172 VSUBS 0.008481f
C210 B.n173 VSUBS 0.008481f
C211 B.n174 VSUBS 0.008481f
C212 B.n175 VSUBS 0.008481f
C213 B.n176 VSUBS 0.008481f
C214 B.n177 VSUBS 0.008481f
C215 B.n178 VSUBS 0.008481f
C216 B.n179 VSUBS 0.008481f
C217 B.n180 VSUBS 0.008481f
C218 B.n181 VSUBS 0.008481f
C219 B.n182 VSUBS 0.008481f
C220 B.n183 VSUBS 0.008481f
C221 B.n184 VSUBS 0.008481f
C222 B.n185 VSUBS 0.008481f
C223 B.n186 VSUBS 0.008481f
C224 B.n187 VSUBS 0.008481f
C225 B.n188 VSUBS 0.019035f
C226 B.n189 VSUBS 0.008481f
C227 B.n190 VSUBS 0.008481f
C228 B.n191 VSUBS 0.008481f
C229 B.n192 VSUBS 0.008481f
C230 B.n193 VSUBS 0.008481f
C231 B.n194 VSUBS 0.008481f
C232 B.n195 VSUBS 0.008481f
C233 B.n196 VSUBS 0.008481f
C234 B.n197 VSUBS 0.008481f
C235 B.n198 VSUBS 0.008481f
C236 B.n199 VSUBS 0.008481f
C237 B.n200 VSUBS 0.008481f
C238 B.n201 VSUBS 0.008481f
C239 B.n202 VSUBS 0.008481f
C240 B.n203 VSUBS 0.008481f
C241 B.n204 VSUBS 0.008481f
C242 B.n205 VSUBS 0.008481f
C243 B.n206 VSUBS 0.008481f
C244 B.n207 VSUBS 0.008481f
C245 B.n208 VSUBS 0.008481f
C246 B.n209 VSUBS 0.008481f
C247 B.n210 VSUBS 0.008481f
C248 B.n211 VSUBS 0.008481f
C249 B.n212 VSUBS 0.008481f
C250 B.n213 VSUBS 0.008481f
C251 B.n214 VSUBS 0.008481f
C252 B.n215 VSUBS 0.008481f
C253 B.n216 VSUBS 0.008481f
C254 B.n217 VSUBS 0.008481f
C255 B.n218 VSUBS 0.008481f
C256 B.n219 VSUBS 0.008481f
C257 B.n220 VSUBS 0.008481f
C258 B.n221 VSUBS 0.008481f
C259 B.n222 VSUBS 0.008481f
C260 B.n223 VSUBS 0.008481f
C261 B.n224 VSUBS 0.008481f
C262 B.n225 VSUBS 0.008481f
C263 B.n226 VSUBS 0.008481f
C264 B.n227 VSUBS 0.008481f
C265 B.n228 VSUBS 0.008481f
C266 B.n229 VSUBS 0.008481f
C267 B.n230 VSUBS 0.008481f
C268 B.n231 VSUBS 0.008481f
C269 B.n232 VSUBS 0.008481f
C270 B.n233 VSUBS 0.008481f
C271 B.n234 VSUBS 0.008481f
C272 B.n235 VSUBS 0.008481f
C273 B.n236 VSUBS 0.008481f
C274 B.n237 VSUBS 0.008481f
C275 B.n238 VSUBS 0.008481f
C276 B.n239 VSUBS 0.008481f
C277 B.n240 VSUBS 0.008481f
C278 B.n241 VSUBS 0.008481f
C279 B.n242 VSUBS 0.008481f
C280 B.n243 VSUBS 0.008481f
C281 B.n244 VSUBS 0.008481f
C282 B.n245 VSUBS 0.008481f
C283 B.n246 VSUBS 0.008481f
C284 B.n247 VSUBS 0.008481f
C285 B.n248 VSUBS 0.008481f
C286 B.n249 VSUBS 0.008481f
C287 B.n250 VSUBS 0.008481f
C288 B.n251 VSUBS 0.008481f
C289 B.n252 VSUBS 0.008481f
C290 B.n253 VSUBS 0.008481f
C291 B.n254 VSUBS 0.008481f
C292 B.n255 VSUBS 0.008481f
C293 B.n256 VSUBS 0.008481f
C294 B.n257 VSUBS 0.019035f
C295 B.n258 VSUBS 0.020625f
C296 B.n259 VSUBS 0.020625f
C297 B.n260 VSUBS 0.008481f
C298 B.n261 VSUBS 0.008481f
C299 B.n262 VSUBS 0.008481f
C300 B.n263 VSUBS 0.008481f
C301 B.n264 VSUBS 0.008481f
C302 B.n265 VSUBS 0.008481f
C303 B.n266 VSUBS 0.008481f
C304 B.n267 VSUBS 0.008481f
C305 B.n268 VSUBS 0.008481f
C306 B.n269 VSUBS 0.008481f
C307 B.n270 VSUBS 0.008481f
C308 B.n271 VSUBS 0.008481f
C309 B.n272 VSUBS 0.008481f
C310 B.n273 VSUBS 0.008481f
C311 B.n274 VSUBS 0.008481f
C312 B.n275 VSUBS 0.008481f
C313 B.n276 VSUBS 0.008481f
C314 B.n277 VSUBS 0.008481f
C315 B.n278 VSUBS 0.008481f
C316 B.n279 VSUBS 0.008481f
C317 B.n280 VSUBS 0.008481f
C318 B.n281 VSUBS 0.008481f
C319 B.n282 VSUBS 0.008481f
C320 B.n283 VSUBS 0.008481f
C321 B.n284 VSUBS 0.008481f
C322 B.n285 VSUBS 0.008481f
C323 B.n286 VSUBS 0.008481f
C324 B.n287 VSUBS 0.008481f
C325 B.n288 VSUBS 0.008481f
C326 B.n289 VSUBS 0.008481f
C327 B.n290 VSUBS 0.008481f
C328 B.n291 VSUBS 0.008481f
C329 B.n292 VSUBS 0.008481f
C330 B.n293 VSUBS 0.008481f
C331 B.n294 VSUBS 0.008481f
C332 B.n295 VSUBS 0.008481f
C333 B.n296 VSUBS 0.008481f
C334 B.n297 VSUBS 0.008481f
C335 B.n298 VSUBS 0.008481f
C336 B.n299 VSUBS 0.008481f
C337 B.n300 VSUBS 0.008481f
C338 B.n301 VSUBS 0.008481f
C339 B.n302 VSUBS 0.008481f
C340 B.n303 VSUBS 0.008481f
C341 B.n304 VSUBS 0.008481f
C342 B.n305 VSUBS 0.008481f
C343 B.n306 VSUBS 0.008481f
C344 B.n307 VSUBS 0.008481f
C345 B.n308 VSUBS 0.008481f
C346 B.n309 VSUBS 0.008481f
C347 B.n310 VSUBS 0.008481f
C348 B.n311 VSUBS 0.008481f
C349 B.n312 VSUBS 0.008481f
C350 B.n313 VSUBS 0.008481f
C351 B.n314 VSUBS 0.008481f
C352 B.n315 VSUBS 0.008481f
C353 B.n316 VSUBS 0.008481f
C354 B.n317 VSUBS 0.008481f
C355 B.n318 VSUBS 0.008481f
C356 B.n319 VSUBS 0.008481f
C357 B.n320 VSUBS 0.008481f
C358 B.n321 VSUBS 0.008481f
C359 B.n322 VSUBS 0.008481f
C360 B.n323 VSUBS 0.008481f
C361 B.n324 VSUBS 0.008481f
C362 B.n325 VSUBS 0.008481f
C363 B.n326 VSUBS 0.008481f
C364 B.n327 VSUBS 0.008481f
C365 B.n328 VSUBS 0.008481f
C366 B.n329 VSUBS 0.008481f
C367 B.n330 VSUBS 0.008481f
C368 B.n331 VSUBS 0.008481f
C369 B.n332 VSUBS 0.008481f
C370 B.n333 VSUBS 0.008481f
C371 B.n334 VSUBS 0.008481f
C372 B.n335 VSUBS 0.008481f
C373 B.n336 VSUBS 0.008481f
C374 B.n337 VSUBS 0.008481f
C375 B.n338 VSUBS 0.008481f
C376 B.n339 VSUBS 0.008481f
C377 B.n340 VSUBS 0.008481f
C378 B.n341 VSUBS 0.008481f
C379 B.t11 VSUBS 0.702983f
C380 B.t10 VSUBS 0.718134f
C381 B.t9 VSUBS 1.13593f
C382 B.n342 VSUBS 0.293435f
C383 B.n343 VSUBS 0.080734f
C384 B.n344 VSUBS 0.019649f
C385 B.n345 VSUBS 0.007982f
C386 B.n346 VSUBS 0.008481f
C387 B.n347 VSUBS 0.008481f
C388 B.n348 VSUBS 0.008481f
C389 B.n349 VSUBS 0.008481f
C390 B.n350 VSUBS 0.008481f
C391 B.n351 VSUBS 0.008481f
C392 B.n352 VSUBS 0.008481f
C393 B.n353 VSUBS 0.008481f
C394 B.n354 VSUBS 0.008481f
C395 B.n355 VSUBS 0.008481f
C396 B.n356 VSUBS 0.008481f
C397 B.n357 VSUBS 0.008481f
C398 B.n358 VSUBS 0.008481f
C399 B.n359 VSUBS 0.008481f
C400 B.n360 VSUBS 0.008481f
C401 B.n361 VSUBS 0.004739f
C402 B.n362 VSUBS 0.019649f
C403 B.n363 VSUBS 0.007982f
C404 B.n364 VSUBS 0.008481f
C405 B.n365 VSUBS 0.008481f
C406 B.n366 VSUBS 0.008481f
C407 B.n367 VSUBS 0.008481f
C408 B.n368 VSUBS 0.008481f
C409 B.n369 VSUBS 0.008481f
C410 B.n370 VSUBS 0.008481f
C411 B.n371 VSUBS 0.008481f
C412 B.n372 VSUBS 0.008481f
C413 B.n373 VSUBS 0.008481f
C414 B.n374 VSUBS 0.008481f
C415 B.n375 VSUBS 0.008481f
C416 B.n376 VSUBS 0.008481f
C417 B.n377 VSUBS 0.008481f
C418 B.n378 VSUBS 0.008481f
C419 B.n379 VSUBS 0.008481f
C420 B.n380 VSUBS 0.008481f
C421 B.n381 VSUBS 0.008481f
C422 B.n382 VSUBS 0.008481f
C423 B.n383 VSUBS 0.008481f
C424 B.n384 VSUBS 0.008481f
C425 B.n385 VSUBS 0.008481f
C426 B.n386 VSUBS 0.008481f
C427 B.n387 VSUBS 0.008481f
C428 B.n388 VSUBS 0.008481f
C429 B.n389 VSUBS 0.008481f
C430 B.n390 VSUBS 0.008481f
C431 B.n391 VSUBS 0.008481f
C432 B.n392 VSUBS 0.008481f
C433 B.n393 VSUBS 0.008481f
C434 B.n394 VSUBS 0.008481f
C435 B.n395 VSUBS 0.008481f
C436 B.n396 VSUBS 0.008481f
C437 B.n397 VSUBS 0.008481f
C438 B.n398 VSUBS 0.008481f
C439 B.n399 VSUBS 0.008481f
C440 B.n400 VSUBS 0.008481f
C441 B.n401 VSUBS 0.008481f
C442 B.n402 VSUBS 0.008481f
C443 B.n403 VSUBS 0.008481f
C444 B.n404 VSUBS 0.008481f
C445 B.n405 VSUBS 0.008481f
C446 B.n406 VSUBS 0.008481f
C447 B.n407 VSUBS 0.008481f
C448 B.n408 VSUBS 0.008481f
C449 B.n409 VSUBS 0.008481f
C450 B.n410 VSUBS 0.008481f
C451 B.n411 VSUBS 0.008481f
C452 B.n412 VSUBS 0.008481f
C453 B.n413 VSUBS 0.008481f
C454 B.n414 VSUBS 0.008481f
C455 B.n415 VSUBS 0.008481f
C456 B.n416 VSUBS 0.008481f
C457 B.n417 VSUBS 0.008481f
C458 B.n418 VSUBS 0.008481f
C459 B.n419 VSUBS 0.008481f
C460 B.n420 VSUBS 0.008481f
C461 B.n421 VSUBS 0.008481f
C462 B.n422 VSUBS 0.008481f
C463 B.n423 VSUBS 0.008481f
C464 B.n424 VSUBS 0.008481f
C465 B.n425 VSUBS 0.008481f
C466 B.n426 VSUBS 0.008481f
C467 B.n427 VSUBS 0.008481f
C468 B.n428 VSUBS 0.008481f
C469 B.n429 VSUBS 0.008481f
C470 B.n430 VSUBS 0.008481f
C471 B.n431 VSUBS 0.008481f
C472 B.n432 VSUBS 0.008481f
C473 B.n433 VSUBS 0.008481f
C474 B.n434 VSUBS 0.008481f
C475 B.n435 VSUBS 0.008481f
C476 B.n436 VSUBS 0.008481f
C477 B.n437 VSUBS 0.008481f
C478 B.n438 VSUBS 0.008481f
C479 B.n439 VSUBS 0.008481f
C480 B.n440 VSUBS 0.008481f
C481 B.n441 VSUBS 0.008481f
C482 B.n442 VSUBS 0.008481f
C483 B.n443 VSUBS 0.008481f
C484 B.n444 VSUBS 0.008481f
C485 B.n445 VSUBS 0.008481f
C486 B.n446 VSUBS 0.008481f
C487 B.n447 VSUBS 0.019622f
C488 B.n448 VSUBS 0.020038f
C489 B.n449 VSUBS 0.019035f
C490 B.n450 VSUBS 0.008481f
C491 B.n451 VSUBS 0.008481f
C492 B.n452 VSUBS 0.008481f
C493 B.n453 VSUBS 0.008481f
C494 B.n454 VSUBS 0.008481f
C495 B.n455 VSUBS 0.008481f
C496 B.n456 VSUBS 0.008481f
C497 B.n457 VSUBS 0.008481f
C498 B.n458 VSUBS 0.008481f
C499 B.n459 VSUBS 0.008481f
C500 B.n460 VSUBS 0.008481f
C501 B.n461 VSUBS 0.008481f
C502 B.n462 VSUBS 0.008481f
C503 B.n463 VSUBS 0.008481f
C504 B.n464 VSUBS 0.008481f
C505 B.n465 VSUBS 0.008481f
C506 B.n466 VSUBS 0.008481f
C507 B.n467 VSUBS 0.008481f
C508 B.n468 VSUBS 0.008481f
C509 B.n469 VSUBS 0.008481f
C510 B.n470 VSUBS 0.008481f
C511 B.n471 VSUBS 0.008481f
C512 B.n472 VSUBS 0.008481f
C513 B.n473 VSUBS 0.008481f
C514 B.n474 VSUBS 0.008481f
C515 B.n475 VSUBS 0.008481f
C516 B.n476 VSUBS 0.008481f
C517 B.n477 VSUBS 0.008481f
C518 B.n478 VSUBS 0.008481f
C519 B.n479 VSUBS 0.008481f
C520 B.n480 VSUBS 0.008481f
C521 B.n481 VSUBS 0.008481f
C522 B.n482 VSUBS 0.008481f
C523 B.n483 VSUBS 0.008481f
C524 B.n484 VSUBS 0.008481f
C525 B.n485 VSUBS 0.008481f
C526 B.n486 VSUBS 0.008481f
C527 B.n487 VSUBS 0.008481f
C528 B.n488 VSUBS 0.008481f
C529 B.n489 VSUBS 0.008481f
C530 B.n490 VSUBS 0.008481f
C531 B.n491 VSUBS 0.008481f
C532 B.n492 VSUBS 0.008481f
C533 B.n493 VSUBS 0.008481f
C534 B.n494 VSUBS 0.008481f
C535 B.n495 VSUBS 0.008481f
C536 B.n496 VSUBS 0.008481f
C537 B.n497 VSUBS 0.008481f
C538 B.n498 VSUBS 0.008481f
C539 B.n499 VSUBS 0.008481f
C540 B.n500 VSUBS 0.008481f
C541 B.n501 VSUBS 0.008481f
C542 B.n502 VSUBS 0.008481f
C543 B.n503 VSUBS 0.008481f
C544 B.n504 VSUBS 0.008481f
C545 B.n505 VSUBS 0.008481f
C546 B.n506 VSUBS 0.008481f
C547 B.n507 VSUBS 0.008481f
C548 B.n508 VSUBS 0.008481f
C549 B.n509 VSUBS 0.008481f
C550 B.n510 VSUBS 0.008481f
C551 B.n511 VSUBS 0.008481f
C552 B.n512 VSUBS 0.008481f
C553 B.n513 VSUBS 0.008481f
C554 B.n514 VSUBS 0.008481f
C555 B.n515 VSUBS 0.008481f
C556 B.n516 VSUBS 0.008481f
C557 B.n517 VSUBS 0.008481f
C558 B.n518 VSUBS 0.008481f
C559 B.n519 VSUBS 0.008481f
C560 B.n520 VSUBS 0.008481f
C561 B.n521 VSUBS 0.008481f
C562 B.n522 VSUBS 0.008481f
C563 B.n523 VSUBS 0.008481f
C564 B.n524 VSUBS 0.008481f
C565 B.n525 VSUBS 0.008481f
C566 B.n526 VSUBS 0.008481f
C567 B.n527 VSUBS 0.008481f
C568 B.n528 VSUBS 0.008481f
C569 B.n529 VSUBS 0.008481f
C570 B.n530 VSUBS 0.008481f
C571 B.n531 VSUBS 0.008481f
C572 B.n532 VSUBS 0.008481f
C573 B.n533 VSUBS 0.008481f
C574 B.n534 VSUBS 0.008481f
C575 B.n535 VSUBS 0.008481f
C576 B.n536 VSUBS 0.008481f
C577 B.n537 VSUBS 0.008481f
C578 B.n538 VSUBS 0.008481f
C579 B.n539 VSUBS 0.008481f
C580 B.n540 VSUBS 0.008481f
C581 B.n541 VSUBS 0.008481f
C582 B.n542 VSUBS 0.008481f
C583 B.n543 VSUBS 0.008481f
C584 B.n544 VSUBS 0.008481f
C585 B.n545 VSUBS 0.008481f
C586 B.n546 VSUBS 0.008481f
C587 B.n547 VSUBS 0.008481f
C588 B.n548 VSUBS 0.008481f
C589 B.n549 VSUBS 0.008481f
C590 B.n550 VSUBS 0.008481f
C591 B.n551 VSUBS 0.008481f
C592 B.n552 VSUBS 0.008481f
C593 B.n553 VSUBS 0.008481f
C594 B.n554 VSUBS 0.008481f
C595 B.n555 VSUBS 0.008481f
C596 B.n556 VSUBS 0.008481f
C597 B.n557 VSUBS 0.008481f
C598 B.n558 VSUBS 0.019035f
C599 B.n559 VSUBS 0.020625f
C600 B.n560 VSUBS 0.020625f
C601 B.n561 VSUBS 0.008481f
C602 B.n562 VSUBS 0.008481f
C603 B.n563 VSUBS 0.008481f
C604 B.n564 VSUBS 0.008481f
C605 B.n565 VSUBS 0.008481f
C606 B.n566 VSUBS 0.008481f
C607 B.n567 VSUBS 0.008481f
C608 B.n568 VSUBS 0.008481f
C609 B.n569 VSUBS 0.008481f
C610 B.n570 VSUBS 0.008481f
C611 B.n571 VSUBS 0.008481f
C612 B.n572 VSUBS 0.008481f
C613 B.n573 VSUBS 0.008481f
C614 B.n574 VSUBS 0.008481f
C615 B.n575 VSUBS 0.008481f
C616 B.n576 VSUBS 0.008481f
C617 B.n577 VSUBS 0.008481f
C618 B.n578 VSUBS 0.008481f
C619 B.n579 VSUBS 0.008481f
C620 B.n580 VSUBS 0.008481f
C621 B.n581 VSUBS 0.008481f
C622 B.n582 VSUBS 0.008481f
C623 B.n583 VSUBS 0.008481f
C624 B.n584 VSUBS 0.008481f
C625 B.n585 VSUBS 0.008481f
C626 B.n586 VSUBS 0.008481f
C627 B.n587 VSUBS 0.008481f
C628 B.n588 VSUBS 0.008481f
C629 B.n589 VSUBS 0.008481f
C630 B.n590 VSUBS 0.008481f
C631 B.n591 VSUBS 0.008481f
C632 B.n592 VSUBS 0.008481f
C633 B.n593 VSUBS 0.008481f
C634 B.n594 VSUBS 0.008481f
C635 B.n595 VSUBS 0.008481f
C636 B.n596 VSUBS 0.008481f
C637 B.n597 VSUBS 0.008481f
C638 B.n598 VSUBS 0.008481f
C639 B.n599 VSUBS 0.008481f
C640 B.n600 VSUBS 0.008481f
C641 B.n601 VSUBS 0.008481f
C642 B.n602 VSUBS 0.008481f
C643 B.n603 VSUBS 0.008481f
C644 B.n604 VSUBS 0.008481f
C645 B.n605 VSUBS 0.008481f
C646 B.n606 VSUBS 0.008481f
C647 B.n607 VSUBS 0.008481f
C648 B.n608 VSUBS 0.008481f
C649 B.n609 VSUBS 0.008481f
C650 B.n610 VSUBS 0.008481f
C651 B.n611 VSUBS 0.008481f
C652 B.n612 VSUBS 0.008481f
C653 B.n613 VSUBS 0.008481f
C654 B.n614 VSUBS 0.008481f
C655 B.n615 VSUBS 0.008481f
C656 B.n616 VSUBS 0.008481f
C657 B.n617 VSUBS 0.008481f
C658 B.n618 VSUBS 0.008481f
C659 B.n619 VSUBS 0.008481f
C660 B.n620 VSUBS 0.008481f
C661 B.n621 VSUBS 0.008481f
C662 B.n622 VSUBS 0.008481f
C663 B.n623 VSUBS 0.008481f
C664 B.n624 VSUBS 0.008481f
C665 B.n625 VSUBS 0.008481f
C666 B.n626 VSUBS 0.008481f
C667 B.n627 VSUBS 0.008481f
C668 B.n628 VSUBS 0.008481f
C669 B.n629 VSUBS 0.008481f
C670 B.n630 VSUBS 0.008481f
C671 B.n631 VSUBS 0.008481f
C672 B.n632 VSUBS 0.008481f
C673 B.n633 VSUBS 0.008481f
C674 B.n634 VSUBS 0.008481f
C675 B.n635 VSUBS 0.008481f
C676 B.n636 VSUBS 0.008481f
C677 B.n637 VSUBS 0.008481f
C678 B.n638 VSUBS 0.008481f
C679 B.n639 VSUBS 0.008481f
C680 B.n640 VSUBS 0.008481f
C681 B.n641 VSUBS 0.008481f
C682 B.n642 VSUBS 0.008481f
C683 B.n643 VSUBS 0.008481f
C684 B.n644 VSUBS 0.007982f
C685 B.n645 VSUBS 0.019649f
C686 B.n646 VSUBS 0.004739f
C687 B.n647 VSUBS 0.008481f
C688 B.n648 VSUBS 0.008481f
C689 B.n649 VSUBS 0.008481f
C690 B.n650 VSUBS 0.008481f
C691 B.n651 VSUBS 0.008481f
C692 B.n652 VSUBS 0.008481f
C693 B.n653 VSUBS 0.008481f
C694 B.n654 VSUBS 0.008481f
C695 B.n655 VSUBS 0.008481f
C696 B.n656 VSUBS 0.008481f
C697 B.n657 VSUBS 0.008481f
C698 B.n658 VSUBS 0.008481f
C699 B.n659 VSUBS 0.004739f
C700 B.n660 VSUBS 0.008481f
C701 B.n661 VSUBS 0.008481f
C702 B.n662 VSUBS 0.008481f
C703 B.n663 VSUBS 0.008481f
C704 B.n664 VSUBS 0.008481f
C705 B.n665 VSUBS 0.008481f
C706 B.n666 VSUBS 0.008481f
C707 B.n667 VSUBS 0.008481f
C708 B.n668 VSUBS 0.008481f
C709 B.n669 VSUBS 0.008481f
C710 B.n670 VSUBS 0.008481f
C711 B.n671 VSUBS 0.008481f
C712 B.n672 VSUBS 0.008481f
C713 B.n673 VSUBS 0.008481f
C714 B.n674 VSUBS 0.008481f
C715 B.n675 VSUBS 0.008481f
C716 B.n676 VSUBS 0.008481f
C717 B.n677 VSUBS 0.008481f
C718 B.n678 VSUBS 0.008481f
C719 B.n679 VSUBS 0.008481f
C720 B.n680 VSUBS 0.008481f
C721 B.n681 VSUBS 0.008481f
C722 B.n682 VSUBS 0.008481f
C723 B.n683 VSUBS 0.008481f
C724 B.n684 VSUBS 0.008481f
C725 B.n685 VSUBS 0.008481f
C726 B.n686 VSUBS 0.008481f
C727 B.n687 VSUBS 0.008481f
C728 B.n688 VSUBS 0.008481f
C729 B.n689 VSUBS 0.008481f
C730 B.n690 VSUBS 0.008481f
C731 B.n691 VSUBS 0.008481f
C732 B.n692 VSUBS 0.008481f
C733 B.n693 VSUBS 0.008481f
C734 B.n694 VSUBS 0.008481f
C735 B.n695 VSUBS 0.008481f
C736 B.n696 VSUBS 0.008481f
C737 B.n697 VSUBS 0.008481f
C738 B.n698 VSUBS 0.008481f
C739 B.n699 VSUBS 0.008481f
C740 B.n700 VSUBS 0.008481f
C741 B.n701 VSUBS 0.008481f
C742 B.n702 VSUBS 0.008481f
C743 B.n703 VSUBS 0.008481f
C744 B.n704 VSUBS 0.008481f
C745 B.n705 VSUBS 0.008481f
C746 B.n706 VSUBS 0.008481f
C747 B.n707 VSUBS 0.008481f
C748 B.n708 VSUBS 0.008481f
C749 B.n709 VSUBS 0.008481f
C750 B.n710 VSUBS 0.008481f
C751 B.n711 VSUBS 0.008481f
C752 B.n712 VSUBS 0.008481f
C753 B.n713 VSUBS 0.008481f
C754 B.n714 VSUBS 0.008481f
C755 B.n715 VSUBS 0.008481f
C756 B.n716 VSUBS 0.008481f
C757 B.n717 VSUBS 0.008481f
C758 B.n718 VSUBS 0.008481f
C759 B.n719 VSUBS 0.008481f
C760 B.n720 VSUBS 0.008481f
C761 B.n721 VSUBS 0.008481f
C762 B.n722 VSUBS 0.008481f
C763 B.n723 VSUBS 0.008481f
C764 B.n724 VSUBS 0.008481f
C765 B.n725 VSUBS 0.008481f
C766 B.n726 VSUBS 0.008481f
C767 B.n727 VSUBS 0.008481f
C768 B.n728 VSUBS 0.008481f
C769 B.n729 VSUBS 0.008481f
C770 B.n730 VSUBS 0.008481f
C771 B.n731 VSUBS 0.008481f
C772 B.n732 VSUBS 0.008481f
C773 B.n733 VSUBS 0.008481f
C774 B.n734 VSUBS 0.008481f
C775 B.n735 VSUBS 0.008481f
C776 B.n736 VSUBS 0.008481f
C777 B.n737 VSUBS 0.008481f
C778 B.n738 VSUBS 0.008481f
C779 B.n739 VSUBS 0.008481f
C780 B.n740 VSUBS 0.008481f
C781 B.n741 VSUBS 0.008481f
C782 B.n742 VSUBS 0.008481f
C783 B.n743 VSUBS 0.008481f
C784 B.n744 VSUBS 0.008481f
C785 B.n745 VSUBS 0.020625f
C786 B.n746 VSUBS 0.019035f
C787 B.n747 VSUBS 0.019035f
C788 B.n748 VSUBS 0.008481f
C789 B.n749 VSUBS 0.008481f
C790 B.n750 VSUBS 0.008481f
C791 B.n751 VSUBS 0.008481f
C792 B.n752 VSUBS 0.008481f
C793 B.n753 VSUBS 0.008481f
C794 B.n754 VSUBS 0.008481f
C795 B.n755 VSUBS 0.008481f
C796 B.n756 VSUBS 0.008481f
C797 B.n757 VSUBS 0.008481f
C798 B.n758 VSUBS 0.008481f
C799 B.n759 VSUBS 0.008481f
C800 B.n760 VSUBS 0.008481f
C801 B.n761 VSUBS 0.008481f
C802 B.n762 VSUBS 0.008481f
C803 B.n763 VSUBS 0.008481f
C804 B.n764 VSUBS 0.008481f
C805 B.n765 VSUBS 0.008481f
C806 B.n766 VSUBS 0.008481f
C807 B.n767 VSUBS 0.008481f
C808 B.n768 VSUBS 0.008481f
C809 B.n769 VSUBS 0.008481f
C810 B.n770 VSUBS 0.008481f
C811 B.n771 VSUBS 0.008481f
C812 B.n772 VSUBS 0.008481f
C813 B.n773 VSUBS 0.008481f
C814 B.n774 VSUBS 0.008481f
C815 B.n775 VSUBS 0.008481f
C816 B.n776 VSUBS 0.008481f
C817 B.n777 VSUBS 0.008481f
C818 B.n778 VSUBS 0.008481f
C819 B.n779 VSUBS 0.008481f
C820 B.n780 VSUBS 0.008481f
C821 B.n781 VSUBS 0.008481f
C822 B.n782 VSUBS 0.008481f
C823 B.n783 VSUBS 0.008481f
C824 B.n784 VSUBS 0.008481f
C825 B.n785 VSUBS 0.008481f
C826 B.n786 VSUBS 0.008481f
C827 B.n787 VSUBS 0.008481f
C828 B.n788 VSUBS 0.008481f
C829 B.n789 VSUBS 0.008481f
C830 B.n790 VSUBS 0.008481f
C831 B.n791 VSUBS 0.008481f
C832 B.n792 VSUBS 0.008481f
C833 B.n793 VSUBS 0.008481f
C834 B.n794 VSUBS 0.008481f
C835 B.n795 VSUBS 0.008481f
C836 B.n796 VSUBS 0.008481f
C837 B.n797 VSUBS 0.008481f
C838 B.n798 VSUBS 0.008481f
C839 B.n799 VSUBS 0.011067f
C840 B.n800 VSUBS 0.011789f
C841 B.n801 VSUBS 0.023444f
C842 VDD1.t1 VSUBS 3.96355f
C843 VDD1.t3 VSUBS 0.36743f
C844 VDD1.t2 VSUBS 0.36743f
C845 VDD1.n0 VSUBS 3.04277f
C846 VDD1.n1 VSUBS 1.41432f
C847 VDD1.t4 VSUBS 3.96353f
C848 VDD1.t6 VSUBS 0.36743f
C849 VDD1.t9 VSUBS 0.36743f
C850 VDD1.n2 VSUBS 3.04277f
C851 VDD1.n3 VSUBS 1.4066f
C852 VDD1.t5 VSUBS 0.36743f
C853 VDD1.t8 VSUBS 0.36743f
C854 VDD1.n4 VSUBS 3.05302f
C855 VDD1.n5 VSUBS 3.13955f
C856 VDD1.t0 VSUBS 0.36743f
C857 VDD1.t7 VSUBS 0.36743f
C858 VDD1.n6 VSUBS 3.04276f
C859 VDD1.n7 VSUBS 3.57031f
C860 VP.n0 VSUBS 0.038412f
C861 VP.t1 VSUBS 2.34776f
C862 VP.n1 VSUBS 0.063806f
C863 VP.n2 VSUBS 0.038412f
C864 VP.t0 VSUBS 2.34776f
C865 VP.n3 VSUBS 0.869248f
C866 VP.n4 VSUBS 0.038412f
C867 VP.t3 VSUBS 2.34776f
C868 VP.n5 VSUBS 0.833182f
C869 VP.n6 VSUBS 0.038412f
C870 VP.t5 VSUBS 2.34776f
C871 VP.n7 VSUBS 0.901136f
C872 VP.n8 VSUBS 0.038412f
C873 VP.t2 VSUBS 2.34776f
C874 VP.n9 VSUBS 0.063806f
C875 VP.n10 VSUBS 0.038412f
C876 VP.t7 VSUBS 2.34776f
C877 VP.n11 VSUBS 0.869248f
C878 VP.n12 VSUBS 0.038412f
C879 VP.t6 VSUBS 2.34776f
C880 VP.n13 VSUBS 0.886055f
C881 VP.t8 VSUBS 2.42641f
C882 VP.n14 VSUBS 0.927718f
C883 VP.n15 VSUBS 0.201921f
C884 VP.n16 VSUBS 0.044506f
C885 VP.n17 VSUBS 0.049461f
C886 VP.n18 VSUBS 0.062214f
C887 VP.n19 VSUBS 0.038412f
C888 VP.n20 VSUBS 0.038412f
C889 VP.n21 VSUBS 0.038412f
C890 VP.n22 VSUBS 0.062214f
C891 VP.n23 VSUBS 0.049461f
C892 VP.t9 VSUBS 2.34776f
C893 VP.n24 VSUBS 0.833182f
C894 VP.n25 VSUBS 0.044506f
C895 VP.n26 VSUBS 0.038412f
C896 VP.n27 VSUBS 0.038412f
C897 VP.n28 VSUBS 0.038412f
C898 VP.n29 VSUBS 0.033492f
C899 VP.n30 VSUBS 0.058883f
C900 VP.n31 VSUBS 0.901136f
C901 VP.n32 VSUBS 2.08515f
C902 VP.n33 VSUBS 2.11292f
C903 VP.n34 VSUBS 0.038412f
C904 VP.n35 VSUBS 0.058883f
C905 VP.n36 VSUBS 0.033492f
C906 VP.n37 VSUBS 0.063806f
C907 VP.n38 VSUBS 0.038412f
C908 VP.n39 VSUBS 0.038412f
C909 VP.n40 VSUBS 0.044506f
C910 VP.n41 VSUBS 0.049461f
C911 VP.n42 VSUBS 0.062214f
C912 VP.n43 VSUBS 0.038412f
C913 VP.n44 VSUBS 0.038412f
C914 VP.n45 VSUBS 0.038412f
C915 VP.n46 VSUBS 0.062214f
C916 VP.n47 VSUBS 0.049461f
C917 VP.t4 VSUBS 2.34776f
C918 VP.n48 VSUBS 0.833182f
C919 VP.n49 VSUBS 0.044506f
C920 VP.n50 VSUBS 0.038412f
C921 VP.n51 VSUBS 0.038412f
C922 VP.n52 VSUBS 0.038412f
C923 VP.n53 VSUBS 0.033492f
C924 VP.n54 VSUBS 0.058883f
C925 VP.n55 VSUBS 0.901136f
C926 VP.n56 VSUBS 0.035155f
C927 VDD2.t4 VSUBS 3.93917f
C928 VDD2.t1 VSUBS 0.365172f
C929 VDD2.t2 VSUBS 0.365172f
C930 VDD2.n0 VSUBS 3.02407f
C931 VDD2.n1 VSUBS 1.39796f
C932 VDD2.t6 VSUBS 0.365172f
C933 VDD2.t5 VSUBS 0.365172f
C934 VDD2.n2 VSUBS 3.03425f
C935 VDD2.n3 VSUBS 3.02023f
C936 VDD2.t0 VSUBS 3.92514f
C937 VDD2.n4 VSUBS 3.55879f
C938 VDD2.t7 VSUBS 0.365172f
C939 VDD2.t9 VSUBS 0.365172f
C940 VDD2.n5 VSUBS 3.02407f
C941 VDD2.n6 VSUBS 0.674603f
C942 VDD2.t3 VSUBS 0.365172f
C943 VDD2.t8 VSUBS 0.365172f
C944 VDD2.n7 VSUBS 3.0342f
C945 VTAIL.t10 VSUBS 0.36961f
C946 VTAIL.t18 VSUBS 0.36961f
C947 VTAIL.n0 VSUBS 2.90045f
C948 VTAIL.n1 VSUBS 0.847376f
C949 VTAIL.t1 VSUBS 3.78923f
C950 VTAIL.n2 VSUBS 0.992057f
C951 VTAIL.t0 VSUBS 0.36961f
C952 VTAIL.t8 VSUBS 0.36961f
C953 VTAIL.n3 VSUBS 2.90045f
C954 VTAIL.n4 VSUBS 0.892782f
C955 VTAIL.t3 VSUBS 0.36961f
C956 VTAIL.t5 VSUBS 0.36961f
C957 VTAIL.n5 VSUBS 2.90045f
C958 VTAIL.n6 VSUBS 2.68264f
C959 VTAIL.t13 VSUBS 0.36961f
C960 VTAIL.t14 VSUBS 0.36961f
C961 VTAIL.n7 VSUBS 2.90045f
C962 VTAIL.n8 VSUBS 2.68263f
C963 VTAIL.t11 VSUBS 0.36961f
C964 VTAIL.t15 VSUBS 0.36961f
C965 VTAIL.n9 VSUBS 2.90045f
C966 VTAIL.n10 VSUBS 0.892776f
C967 VTAIL.t12 VSUBS 3.78926f
C968 VTAIL.n11 VSUBS 0.992028f
C969 VTAIL.t9 VSUBS 0.36961f
C970 VTAIL.t6 VSUBS 0.36961f
C971 VTAIL.n12 VSUBS 2.90045f
C972 VTAIL.n13 VSUBS 0.872805f
C973 VTAIL.t7 VSUBS 0.36961f
C974 VTAIL.t4 VSUBS 0.36961f
C975 VTAIL.n14 VSUBS 2.90045f
C976 VTAIL.n15 VSUBS 0.892776f
C977 VTAIL.t2 VSUBS 3.78923f
C978 VTAIL.n16 VSUBS 2.6798f
C979 VTAIL.t16 VSUBS 3.78923f
C980 VTAIL.n17 VSUBS 2.6798f
C981 VTAIL.t19 VSUBS 0.36961f
C982 VTAIL.t17 VSUBS 0.36961f
C983 VTAIL.n18 VSUBS 2.90045f
C984 VTAIL.n19 VSUBS 0.79613f
C985 VN.n0 VSUBS 0.037665f
C986 VN.t4 VSUBS 2.30208f
C987 VN.n1 VSUBS 0.062565f
C988 VN.n2 VSUBS 0.037665f
C989 VN.t7 VSUBS 2.30208f
C990 VN.n3 VSUBS 0.852336f
C991 VN.n4 VSUBS 0.037665f
C992 VN.t8 VSUBS 2.30208f
C993 VN.n5 VSUBS 0.868816f
C994 VN.t5 VSUBS 2.3792f
C995 VN.n6 VSUBS 0.909668f
C996 VN.n7 VSUBS 0.197993f
C997 VN.n8 VSUBS 0.04364f
C998 VN.n9 VSUBS 0.048499f
C999 VN.n10 VSUBS 0.061004f
C1000 VN.n11 VSUBS 0.037665f
C1001 VN.n12 VSUBS 0.037665f
C1002 VN.n13 VSUBS 0.037665f
C1003 VN.n14 VSUBS 0.061004f
C1004 VN.n15 VSUBS 0.048499f
C1005 VN.t3 VSUBS 2.30208f
C1006 VN.n16 VSUBS 0.816972f
C1007 VN.n17 VSUBS 0.04364f
C1008 VN.n18 VSUBS 0.037665f
C1009 VN.n19 VSUBS 0.037665f
C1010 VN.n20 VSUBS 0.037665f
C1011 VN.n21 VSUBS 0.032841f
C1012 VN.n22 VSUBS 0.057737f
C1013 VN.n23 VSUBS 0.883603f
C1014 VN.n24 VSUBS 0.034471f
C1015 VN.n25 VSUBS 0.037665f
C1016 VN.t9 VSUBS 2.30208f
C1017 VN.n26 VSUBS 0.062565f
C1018 VN.n27 VSUBS 0.037665f
C1019 VN.t2 VSUBS 2.30208f
C1020 VN.n28 VSUBS 0.816972f
C1021 VN.t0 VSUBS 2.30208f
C1022 VN.n29 VSUBS 0.852336f
C1023 VN.n30 VSUBS 0.037665f
C1024 VN.t6 VSUBS 2.30208f
C1025 VN.n31 VSUBS 0.868816f
C1026 VN.t1 VSUBS 2.3792f
C1027 VN.n32 VSUBS 0.909668f
C1028 VN.n33 VSUBS 0.197993f
C1029 VN.n34 VSUBS 0.04364f
C1030 VN.n35 VSUBS 0.048499f
C1031 VN.n36 VSUBS 0.061004f
C1032 VN.n37 VSUBS 0.037665f
C1033 VN.n38 VSUBS 0.037665f
C1034 VN.n39 VSUBS 0.037665f
C1035 VN.n40 VSUBS 0.061004f
C1036 VN.n41 VSUBS 0.048499f
C1037 VN.n42 VSUBS 0.04364f
C1038 VN.n43 VSUBS 0.037665f
C1039 VN.n44 VSUBS 0.037665f
C1040 VN.n45 VSUBS 0.037665f
C1041 VN.n46 VSUBS 0.032841f
C1042 VN.n47 VSUBS 0.057737f
C1043 VN.n48 VSUBS 0.883603f
C1044 VN.n49 VSUBS 2.06907f
.ends

