* NGSPICE file created from diff_pair_sample_1300.ext - technology: sky130A

.subckt diff_pair_sample_1300 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X1 VTAIL.t18 VN.t1 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X2 VTAIL.t9 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X3 VTAIL.t8 VP.t1 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X4 VDD1.t7 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=2.14005 ps=13.3 w=12.97 l=0.87
X5 VDD1.t6 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=5.0583 ps=26.72 w=12.97 l=0.87
X6 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X7 VDD1.t4 VP.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=5.0583 ps=26.72 w=12.97 l=0.87
X8 VDD1.t3 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=0 ps=0 w=12.97 l=0.87
X10 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=2.14005 ps=13.3 w=12.97 l=0.87
X11 VDD2.t2 VN.t2 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=5.0583 ps=26.72 w=12.97 l=0.87
X12 VDD2.t3 VN.t3 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X13 VDD2.t6 VN.t4 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=5.0583 ps=26.72 w=12.97 l=0.87
X14 VDD2.t1 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X15 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=0 ps=0 w=12.97 l=0.87
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=0 ps=0 w=12.97 l=0.87
X17 VTAIL.t13 VN.t6 VDD2.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X18 VTAIL.t12 VN.t7 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X19 VTAIL.t4 VP.t8 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X20 VDD2.t0 VN.t8 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=2.14005 ps=13.3 w=12.97 l=0.87
X21 VTAIL.t5 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.14005 pd=13.3 as=2.14005 ps=13.3 w=12.97 l=0.87
X22 VDD2.t5 VN.t9 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=2.14005 ps=13.3 w=12.97 l=0.87
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0583 pd=26.72 as=0 ps=0 w=12.97 l=0.87
R0 VN.n4 VN.t9 419.642
R1 VN.n21 VN.t4 419.642
R2 VN.n15 VN.t2 404.714
R3 VN.n32 VN.t8 404.714
R4 VN.n8 VN.t3 359.284
R5 VN.n3 VN.t7 359.284
R6 VN.n13 VN.t6 359.284
R7 VN.n25 VN.t5 359.284
R8 VN.n20 VN.t0 359.284
R9 VN.n30 VN.t1 359.284
R10 VN.n31 VN.n17 161.3
R11 VN.n29 VN.n28 161.3
R12 VN.n27 VN.n18 161.3
R13 VN.n26 VN.n25 161.3
R14 VN.n24 VN.n19 161.3
R15 VN.n23 VN.n22 161.3
R16 VN.n14 VN.n0 161.3
R17 VN.n12 VN.n11 161.3
R18 VN.n10 VN.n1 161.3
R19 VN.n9 VN.n8 161.3
R20 VN.n7 VN.n2 161.3
R21 VN.n6 VN.n5 161.3
R22 VN.n33 VN.n32 80.6037
R23 VN.n16 VN.n15 80.6037
R24 VN.n15 VN.n14 54.8066
R25 VN.n32 VN.n31 54.8066
R26 VN.n7 VN.n6 50.2061
R27 VN.n12 VN.n1 50.2061
R28 VN.n24 VN.n23 50.2061
R29 VN.n29 VN.n18 50.2061
R30 VN VN.n33 44.84
R31 VN.n4 VN.n3 44.4469
R32 VN.n21 VN.n20 44.4469
R33 VN.n22 VN.n21 44.1212
R34 VN.n5 VN.n4 44.1212
R35 VN.n8 VN.n7 30.7807
R36 VN.n8 VN.n1 30.7807
R37 VN.n25 VN.n24 30.7807
R38 VN.n25 VN.n18 30.7807
R39 VN.n14 VN.n13 14.6807
R40 VN.n31 VN.n30 14.6807
R41 VN.n6 VN.n3 9.7873
R42 VN.n13 VN.n12 9.7873
R43 VN.n23 VN.n20 9.7873
R44 VN.n30 VN.n29 9.7873
R45 VN.n33 VN.n17 0.285035
R46 VN.n16 VN.n0 0.285035
R47 VN.n28 VN.n17 0.189894
R48 VN.n28 VN.n27 0.189894
R49 VN.n27 VN.n26 0.189894
R50 VN.n26 VN.n19 0.189894
R51 VN.n22 VN.n19 0.189894
R52 VN.n5 VN.n2 0.189894
R53 VN.n9 VN.n2 0.189894
R54 VN.n10 VN.n9 0.189894
R55 VN.n11 VN.n10 0.189894
R56 VN.n11 VN.n0 0.189894
R57 VN VN.n16 0.146778
R58 VDD2.n1 VDD2.t5 66.2581
R59 VDD2.n4 VDD2.t0 65.2247
R60 VDD2.n3 VDD2.n2 64.4175
R61 VDD2 VDD2.n7 64.4147
R62 VDD2.n6 VDD2.n5 63.6982
R63 VDD2.n1 VDD2.n0 63.697
R64 VDD2.n4 VDD2.n3 39.8101
R65 VDD2.n7 VDD2.t4 1.5271
R66 VDD2.n7 VDD2.t6 1.5271
R67 VDD2.n5 VDD2.t7 1.5271
R68 VDD2.n5 VDD2.t1 1.5271
R69 VDD2.n2 VDD2.t9 1.5271
R70 VDD2.n2 VDD2.t2 1.5271
R71 VDD2.n0 VDD2.t8 1.5271
R72 VDD2.n0 VDD2.t3 1.5271
R73 VDD2.n6 VDD2.n4 1.03498
R74 VDD2 VDD2.n6 0.31731
R75 VDD2.n3 VDD2.n1 0.203775
R76 VTAIL.n11 VTAIL.t15 48.546
R77 VTAIL.n17 VTAIL.t17 48.5448
R78 VTAIL.n2 VTAIL.t7 48.5448
R79 VTAIL.n16 VTAIL.t3 48.5448
R80 VTAIL.n15 VTAIL.n14 47.0194
R81 VTAIL.n13 VTAIL.n12 47.0194
R82 VTAIL.n10 VTAIL.n9 47.0194
R83 VTAIL.n8 VTAIL.n7 47.0194
R84 VTAIL.n19 VTAIL.n18 47.0182
R85 VTAIL.n1 VTAIL.n0 47.0182
R86 VTAIL.n4 VTAIL.n3 47.0182
R87 VTAIL.n6 VTAIL.n5 47.0182
R88 VTAIL.n8 VTAIL.n6 25.6169
R89 VTAIL.n17 VTAIL.n16 24.5824
R90 VTAIL.n18 VTAIL.t16 1.5271
R91 VTAIL.n18 VTAIL.t13 1.5271
R92 VTAIL.n0 VTAIL.t10 1.5271
R93 VTAIL.n0 VTAIL.t12 1.5271
R94 VTAIL.n3 VTAIL.t1 1.5271
R95 VTAIL.n3 VTAIL.t9 1.5271
R96 VTAIL.n5 VTAIL.t6 1.5271
R97 VTAIL.n5 VTAIL.t8 1.5271
R98 VTAIL.n14 VTAIL.t2 1.5271
R99 VTAIL.n14 VTAIL.t4 1.5271
R100 VTAIL.n12 VTAIL.t0 1.5271
R101 VTAIL.n12 VTAIL.t5 1.5271
R102 VTAIL.n9 VTAIL.t14 1.5271
R103 VTAIL.n9 VTAIL.t19 1.5271
R104 VTAIL.n7 VTAIL.t11 1.5271
R105 VTAIL.n7 VTAIL.t18 1.5271
R106 VTAIL.n10 VTAIL.n8 1.03498
R107 VTAIL.n11 VTAIL.n10 1.03498
R108 VTAIL.n15 VTAIL.n13 1.03498
R109 VTAIL.n16 VTAIL.n15 1.03498
R110 VTAIL.n6 VTAIL.n4 1.03498
R111 VTAIL.n4 VTAIL.n2 1.03498
R112 VTAIL.n19 VTAIL.n17 1.03498
R113 VTAIL.n13 VTAIL.n11 0.987569
R114 VTAIL.n2 VTAIL.n1 0.987569
R115 VTAIL VTAIL.n1 0.834552
R116 VTAIL VTAIL.n19 0.200931
R117 B.n604 B.n355 588.598
R118 B.n111 B.n53 588.598
R119 B.n607 B.n357 588.598
R120 B.n735 B.n55 588.598
R121 B.n735 B.n734 585
R122 B.n303 B.n104 585
R123 B.n302 B.n301 585
R124 B.n300 B.n299 585
R125 B.n298 B.n297 585
R126 B.n296 B.n295 585
R127 B.n294 B.n293 585
R128 B.n292 B.n291 585
R129 B.n290 B.n289 585
R130 B.n288 B.n287 585
R131 B.n286 B.n285 585
R132 B.n284 B.n283 585
R133 B.n282 B.n281 585
R134 B.n280 B.n279 585
R135 B.n278 B.n277 585
R136 B.n276 B.n275 585
R137 B.n274 B.n273 585
R138 B.n272 B.n271 585
R139 B.n270 B.n269 585
R140 B.n268 B.n267 585
R141 B.n266 B.n265 585
R142 B.n264 B.n263 585
R143 B.n262 B.n261 585
R144 B.n260 B.n259 585
R145 B.n258 B.n257 585
R146 B.n256 B.n255 585
R147 B.n254 B.n253 585
R148 B.n252 B.n251 585
R149 B.n250 B.n249 585
R150 B.n248 B.n247 585
R151 B.n246 B.n245 585
R152 B.n244 B.n243 585
R153 B.n242 B.n241 585
R154 B.n240 B.n239 585
R155 B.n238 B.n237 585
R156 B.n236 B.n235 585
R157 B.n234 B.n233 585
R158 B.n232 B.n231 585
R159 B.n230 B.n229 585
R160 B.n228 B.n227 585
R161 B.n226 B.n225 585
R162 B.n224 B.n223 585
R163 B.n222 B.n221 585
R164 B.n220 B.n219 585
R165 B.n218 B.n217 585
R166 B.n216 B.n215 585
R167 B.n214 B.n213 585
R168 B.n212 B.n211 585
R169 B.n210 B.n209 585
R170 B.n208 B.n207 585
R171 B.n206 B.n205 585
R172 B.n204 B.n203 585
R173 B.n202 B.n201 585
R174 B.n200 B.n199 585
R175 B.n198 B.n197 585
R176 B.n196 B.n195 585
R177 B.n194 B.n193 585
R178 B.n192 B.n191 585
R179 B.n190 B.n189 585
R180 B.n188 B.n187 585
R181 B.n186 B.n185 585
R182 B.n184 B.n183 585
R183 B.n182 B.n181 585
R184 B.n180 B.n179 585
R185 B.n178 B.n177 585
R186 B.n176 B.n175 585
R187 B.n174 B.n173 585
R188 B.n172 B.n171 585
R189 B.n170 B.n169 585
R190 B.n168 B.n167 585
R191 B.n166 B.n165 585
R192 B.n164 B.n163 585
R193 B.n162 B.n161 585
R194 B.n160 B.n159 585
R195 B.n158 B.n157 585
R196 B.n156 B.n155 585
R197 B.n154 B.n153 585
R198 B.n152 B.n151 585
R199 B.n150 B.n149 585
R200 B.n148 B.n147 585
R201 B.n146 B.n145 585
R202 B.n144 B.n143 585
R203 B.n142 B.n141 585
R204 B.n140 B.n139 585
R205 B.n138 B.n137 585
R206 B.n136 B.n135 585
R207 B.n134 B.n133 585
R208 B.n132 B.n131 585
R209 B.n130 B.n129 585
R210 B.n128 B.n127 585
R211 B.n126 B.n125 585
R212 B.n124 B.n123 585
R213 B.n122 B.n121 585
R214 B.n120 B.n119 585
R215 B.n118 B.n117 585
R216 B.n116 B.n115 585
R217 B.n114 B.n113 585
R218 B.n112 B.n111 585
R219 B.n733 B.n55 585
R220 B.n738 B.n55 585
R221 B.n732 B.n54 585
R222 B.n739 B.n54 585
R223 B.n731 B.n730 585
R224 B.n730 B.n50 585
R225 B.n729 B.n49 585
R226 B.n745 B.n49 585
R227 B.n728 B.n48 585
R228 B.n746 B.n48 585
R229 B.n727 B.n47 585
R230 B.n747 B.n47 585
R231 B.n726 B.n725 585
R232 B.n725 B.n43 585
R233 B.n724 B.n42 585
R234 B.n753 B.n42 585
R235 B.n723 B.n41 585
R236 B.n754 B.n41 585
R237 B.n722 B.n40 585
R238 B.n755 B.n40 585
R239 B.n721 B.n720 585
R240 B.n720 B.n36 585
R241 B.n719 B.n35 585
R242 B.n761 B.n35 585
R243 B.n718 B.n34 585
R244 B.n762 B.n34 585
R245 B.n717 B.n33 585
R246 B.n763 B.n33 585
R247 B.n716 B.n715 585
R248 B.n715 B.n29 585
R249 B.n714 B.n28 585
R250 B.n769 B.n28 585
R251 B.n713 B.n27 585
R252 B.n770 B.n27 585
R253 B.n712 B.n26 585
R254 B.n771 B.n26 585
R255 B.n711 B.n710 585
R256 B.n710 B.n25 585
R257 B.n709 B.n21 585
R258 B.n777 B.n21 585
R259 B.n708 B.n20 585
R260 B.n778 B.n20 585
R261 B.n707 B.n19 585
R262 B.n779 B.n19 585
R263 B.n706 B.n705 585
R264 B.n705 B.n18 585
R265 B.n704 B.n14 585
R266 B.n785 B.n14 585
R267 B.n703 B.n13 585
R268 B.n786 B.n13 585
R269 B.n702 B.n12 585
R270 B.n787 B.n12 585
R271 B.n701 B.n700 585
R272 B.n700 B.n8 585
R273 B.n699 B.n7 585
R274 B.n793 B.n7 585
R275 B.n698 B.n6 585
R276 B.n794 B.n6 585
R277 B.n697 B.n5 585
R278 B.n795 B.n5 585
R279 B.n696 B.n695 585
R280 B.n695 B.n4 585
R281 B.n694 B.n304 585
R282 B.n694 B.n693 585
R283 B.n684 B.n305 585
R284 B.n306 B.n305 585
R285 B.n686 B.n685 585
R286 B.n687 B.n686 585
R287 B.n683 B.n311 585
R288 B.n311 B.n310 585
R289 B.n682 B.n681 585
R290 B.n681 B.n680 585
R291 B.n313 B.n312 585
R292 B.n673 B.n313 585
R293 B.n672 B.n671 585
R294 B.n674 B.n672 585
R295 B.n670 B.n318 585
R296 B.n318 B.n317 585
R297 B.n669 B.n668 585
R298 B.n668 B.n667 585
R299 B.n320 B.n319 585
R300 B.n660 B.n320 585
R301 B.n659 B.n658 585
R302 B.n661 B.n659 585
R303 B.n657 B.n325 585
R304 B.n325 B.n324 585
R305 B.n656 B.n655 585
R306 B.n655 B.n654 585
R307 B.n327 B.n326 585
R308 B.n328 B.n327 585
R309 B.n647 B.n646 585
R310 B.n648 B.n647 585
R311 B.n645 B.n333 585
R312 B.n333 B.n332 585
R313 B.n644 B.n643 585
R314 B.n643 B.n642 585
R315 B.n335 B.n334 585
R316 B.n336 B.n335 585
R317 B.n635 B.n634 585
R318 B.n636 B.n635 585
R319 B.n633 B.n341 585
R320 B.n341 B.n340 585
R321 B.n632 B.n631 585
R322 B.n631 B.n630 585
R323 B.n343 B.n342 585
R324 B.n344 B.n343 585
R325 B.n623 B.n622 585
R326 B.n624 B.n623 585
R327 B.n621 B.n348 585
R328 B.n352 B.n348 585
R329 B.n620 B.n619 585
R330 B.n619 B.n618 585
R331 B.n350 B.n349 585
R332 B.n351 B.n350 585
R333 B.n611 B.n610 585
R334 B.n612 B.n611 585
R335 B.n609 B.n357 585
R336 B.n357 B.n356 585
R337 B.n604 B.n603 585
R338 B.n602 B.n408 585
R339 B.n601 B.n407 585
R340 B.n606 B.n407 585
R341 B.n600 B.n599 585
R342 B.n598 B.n597 585
R343 B.n596 B.n595 585
R344 B.n594 B.n593 585
R345 B.n592 B.n591 585
R346 B.n590 B.n589 585
R347 B.n588 B.n587 585
R348 B.n586 B.n585 585
R349 B.n584 B.n583 585
R350 B.n582 B.n581 585
R351 B.n580 B.n579 585
R352 B.n578 B.n577 585
R353 B.n576 B.n575 585
R354 B.n574 B.n573 585
R355 B.n572 B.n571 585
R356 B.n570 B.n569 585
R357 B.n568 B.n567 585
R358 B.n566 B.n565 585
R359 B.n564 B.n563 585
R360 B.n562 B.n561 585
R361 B.n560 B.n559 585
R362 B.n558 B.n557 585
R363 B.n556 B.n555 585
R364 B.n554 B.n553 585
R365 B.n552 B.n551 585
R366 B.n550 B.n549 585
R367 B.n548 B.n547 585
R368 B.n546 B.n545 585
R369 B.n544 B.n543 585
R370 B.n542 B.n541 585
R371 B.n540 B.n539 585
R372 B.n538 B.n537 585
R373 B.n536 B.n535 585
R374 B.n534 B.n533 585
R375 B.n532 B.n531 585
R376 B.n530 B.n529 585
R377 B.n528 B.n527 585
R378 B.n526 B.n525 585
R379 B.n524 B.n523 585
R380 B.n522 B.n521 585
R381 B.n520 B.n519 585
R382 B.n517 B.n516 585
R383 B.n515 B.n514 585
R384 B.n513 B.n512 585
R385 B.n511 B.n510 585
R386 B.n509 B.n508 585
R387 B.n507 B.n506 585
R388 B.n505 B.n504 585
R389 B.n503 B.n502 585
R390 B.n501 B.n500 585
R391 B.n499 B.n498 585
R392 B.n496 B.n495 585
R393 B.n494 B.n493 585
R394 B.n492 B.n491 585
R395 B.n490 B.n489 585
R396 B.n488 B.n487 585
R397 B.n486 B.n485 585
R398 B.n484 B.n483 585
R399 B.n482 B.n481 585
R400 B.n480 B.n479 585
R401 B.n478 B.n477 585
R402 B.n476 B.n475 585
R403 B.n474 B.n473 585
R404 B.n472 B.n471 585
R405 B.n470 B.n469 585
R406 B.n468 B.n467 585
R407 B.n466 B.n465 585
R408 B.n464 B.n463 585
R409 B.n462 B.n461 585
R410 B.n460 B.n459 585
R411 B.n458 B.n457 585
R412 B.n456 B.n455 585
R413 B.n454 B.n453 585
R414 B.n452 B.n451 585
R415 B.n450 B.n449 585
R416 B.n448 B.n447 585
R417 B.n446 B.n445 585
R418 B.n444 B.n443 585
R419 B.n442 B.n441 585
R420 B.n440 B.n439 585
R421 B.n438 B.n437 585
R422 B.n436 B.n435 585
R423 B.n434 B.n433 585
R424 B.n432 B.n431 585
R425 B.n430 B.n429 585
R426 B.n428 B.n427 585
R427 B.n426 B.n425 585
R428 B.n424 B.n423 585
R429 B.n422 B.n421 585
R430 B.n420 B.n419 585
R431 B.n418 B.n417 585
R432 B.n416 B.n415 585
R433 B.n414 B.n413 585
R434 B.n359 B.n358 585
R435 B.n608 B.n607 585
R436 B.n607 B.n606 585
R437 B.n355 B.n354 585
R438 B.n356 B.n355 585
R439 B.n614 B.n613 585
R440 B.n613 B.n612 585
R441 B.n615 B.n353 585
R442 B.n353 B.n351 585
R443 B.n617 B.n616 585
R444 B.n618 B.n617 585
R445 B.n347 B.n346 585
R446 B.n352 B.n347 585
R447 B.n626 B.n625 585
R448 B.n625 B.n624 585
R449 B.n627 B.n345 585
R450 B.n345 B.n344 585
R451 B.n629 B.n628 585
R452 B.n630 B.n629 585
R453 B.n339 B.n338 585
R454 B.n340 B.n339 585
R455 B.n638 B.n637 585
R456 B.n637 B.n636 585
R457 B.n639 B.n337 585
R458 B.n337 B.n336 585
R459 B.n641 B.n640 585
R460 B.n642 B.n641 585
R461 B.n331 B.n330 585
R462 B.n332 B.n331 585
R463 B.n650 B.n649 585
R464 B.n649 B.n648 585
R465 B.n651 B.n329 585
R466 B.n329 B.n328 585
R467 B.n653 B.n652 585
R468 B.n654 B.n653 585
R469 B.n323 B.n322 585
R470 B.n324 B.n323 585
R471 B.n663 B.n662 585
R472 B.n662 B.n661 585
R473 B.n664 B.n321 585
R474 B.n660 B.n321 585
R475 B.n666 B.n665 585
R476 B.n667 B.n666 585
R477 B.n316 B.n315 585
R478 B.n317 B.n316 585
R479 B.n676 B.n675 585
R480 B.n675 B.n674 585
R481 B.n677 B.n314 585
R482 B.n673 B.n314 585
R483 B.n679 B.n678 585
R484 B.n680 B.n679 585
R485 B.n309 B.n308 585
R486 B.n310 B.n309 585
R487 B.n689 B.n688 585
R488 B.n688 B.n687 585
R489 B.n690 B.n307 585
R490 B.n307 B.n306 585
R491 B.n692 B.n691 585
R492 B.n693 B.n692 585
R493 B.n2 B.n0 585
R494 B.n4 B.n2 585
R495 B.n3 B.n1 585
R496 B.n794 B.n3 585
R497 B.n792 B.n791 585
R498 B.n793 B.n792 585
R499 B.n790 B.n9 585
R500 B.n9 B.n8 585
R501 B.n789 B.n788 585
R502 B.n788 B.n787 585
R503 B.n11 B.n10 585
R504 B.n786 B.n11 585
R505 B.n784 B.n783 585
R506 B.n785 B.n784 585
R507 B.n782 B.n15 585
R508 B.n18 B.n15 585
R509 B.n781 B.n780 585
R510 B.n780 B.n779 585
R511 B.n17 B.n16 585
R512 B.n778 B.n17 585
R513 B.n776 B.n775 585
R514 B.n777 B.n776 585
R515 B.n774 B.n22 585
R516 B.n25 B.n22 585
R517 B.n773 B.n772 585
R518 B.n772 B.n771 585
R519 B.n24 B.n23 585
R520 B.n770 B.n24 585
R521 B.n768 B.n767 585
R522 B.n769 B.n768 585
R523 B.n766 B.n30 585
R524 B.n30 B.n29 585
R525 B.n765 B.n764 585
R526 B.n764 B.n763 585
R527 B.n32 B.n31 585
R528 B.n762 B.n32 585
R529 B.n760 B.n759 585
R530 B.n761 B.n760 585
R531 B.n758 B.n37 585
R532 B.n37 B.n36 585
R533 B.n757 B.n756 585
R534 B.n756 B.n755 585
R535 B.n39 B.n38 585
R536 B.n754 B.n39 585
R537 B.n752 B.n751 585
R538 B.n753 B.n752 585
R539 B.n750 B.n44 585
R540 B.n44 B.n43 585
R541 B.n749 B.n748 585
R542 B.n748 B.n747 585
R543 B.n46 B.n45 585
R544 B.n746 B.n46 585
R545 B.n744 B.n743 585
R546 B.n745 B.n744 585
R547 B.n742 B.n51 585
R548 B.n51 B.n50 585
R549 B.n741 B.n740 585
R550 B.n740 B.n739 585
R551 B.n53 B.n52 585
R552 B.n738 B.n53 585
R553 B.n797 B.n796 585
R554 B.n796 B.n795 585
R555 B.n411 B.t10 561.24
R556 B.n409 B.t18 561.24
R557 B.n108 B.t21 561.24
R558 B.n105 B.t14 561.24
R559 B.n737 B.n736 256.663
R560 B.n737 B.n103 256.663
R561 B.n737 B.n102 256.663
R562 B.n737 B.n101 256.663
R563 B.n737 B.n100 256.663
R564 B.n737 B.n99 256.663
R565 B.n737 B.n98 256.663
R566 B.n737 B.n97 256.663
R567 B.n737 B.n96 256.663
R568 B.n737 B.n95 256.663
R569 B.n737 B.n94 256.663
R570 B.n737 B.n93 256.663
R571 B.n737 B.n92 256.663
R572 B.n737 B.n91 256.663
R573 B.n737 B.n90 256.663
R574 B.n737 B.n89 256.663
R575 B.n737 B.n88 256.663
R576 B.n737 B.n87 256.663
R577 B.n737 B.n86 256.663
R578 B.n737 B.n85 256.663
R579 B.n737 B.n84 256.663
R580 B.n737 B.n83 256.663
R581 B.n737 B.n82 256.663
R582 B.n737 B.n81 256.663
R583 B.n737 B.n80 256.663
R584 B.n737 B.n79 256.663
R585 B.n737 B.n78 256.663
R586 B.n737 B.n77 256.663
R587 B.n737 B.n76 256.663
R588 B.n737 B.n75 256.663
R589 B.n737 B.n74 256.663
R590 B.n737 B.n73 256.663
R591 B.n737 B.n72 256.663
R592 B.n737 B.n71 256.663
R593 B.n737 B.n70 256.663
R594 B.n737 B.n69 256.663
R595 B.n737 B.n68 256.663
R596 B.n737 B.n67 256.663
R597 B.n737 B.n66 256.663
R598 B.n737 B.n65 256.663
R599 B.n737 B.n64 256.663
R600 B.n737 B.n63 256.663
R601 B.n737 B.n62 256.663
R602 B.n737 B.n61 256.663
R603 B.n737 B.n60 256.663
R604 B.n737 B.n59 256.663
R605 B.n737 B.n58 256.663
R606 B.n737 B.n57 256.663
R607 B.n737 B.n56 256.663
R608 B.n606 B.n605 256.663
R609 B.n606 B.n360 256.663
R610 B.n606 B.n361 256.663
R611 B.n606 B.n362 256.663
R612 B.n606 B.n363 256.663
R613 B.n606 B.n364 256.663
R614 B.n606 B.n365 256.663
R615 B.n606 B.n366 256.663
R616 B.n606 B.n367 256.663
R617 B.n606 B.n368 256.663
R618 B.n606 B.n369 256.663
R619 B.n606 B.n370 256.663
R620 B.n606 B.n371 256.663
R621 B.n606 B.n372 256.663
R622 B.n606 B.n373 256.663
R623 B.n606 B.n374 256.663
R624 B.n606 B.n375 256.663
R625 B.n606 B.n376 256.663
R626 B.n606 B.n377 256.663
R627 B.n606 B.n378 256.663
R628 B.n606 B.n379 256.663
R629 B.n606 B.n380 256.663
R630 B.n606 B.n381 256.663
R631 B.n606 B.n382 256.663
R632 B.n606 B.n383 256.663
R633 B.n606 B.n384 256.663
R634 B.n606 B.n385 256.663
R635 B.n606 B.n386 256.663
R636 B.n606 B.n387 256.663
R637 B.n606 B.n388 256.663
R638 B.n606 B.n389 256.663
R639 B.n606 B.n390 256.663
R640 B.n606 B.n391 256.663
R641 B.n606 B.n392 256.663
R642 B.n606 B.n393 256.663
R643 B.n606 B.n394 256.663
R644 B.n606 B.n395 256.663
R645 B.n606 B.n396 256.663
R646 B.n606 B.n397 256.663
R647 B.n606 B.n398 256.663
R648 B.n606 B.n399 256.663
R649 B.n606 B.n400 256.663
R650 B.n606 B.n401 256.663
R651 B.n606 B.n402 256.663
R652 B.n606 B.n403 256.663
R653 B.n606 B.n404 256.663
R654 B.n606 B.n405 256.663
R655 B.n606 B.n406 256.663
R656 B.n613 B.n355 163.367
R657 B.n613 B.n353 163.367
R658 B.n617 B.n353 163.367
R659 B.n617 B.n347 163.367
R660 B.n625 B.n347 163.367
R661 B.n625 B.n345 163.367
R662 B.n629 B.n345 163.367
R663 B.n629 B.n339 163.367
R664 B.n637 B.n339 163.367
R665 B.n637 B.n337 163.367
R666 B.n641 B.n337 163.367
R667 B.n641 B.n331 163.367
R668 B.n649 B.n331 163.367
R669 B.n649 B.n329 163.367
R670 B.n653 B.n329 163.367
R671 B.n653 B.n323 163.367
R672 B.n662 B.n323 163.367
R673 B.n662 B.n321 163.367
R674 B.n666 B.n321 163.367
R675 B.n666 B.n316 163.367
R676 B.n675 B.n316 163.367
R677 B.n675 B.n314 163.367
R678 B.n679 B.n314 163.367
R679 B.n679 B.n309 163.367
R680 B.n688 B.n309 163.367
R681 B.n688 B.n307 163.367
R682 B.n692 B.n307 163.367
R683 B.n692 B.n2 163.367
R684 B.n796 B.n2 163.367
R685 B.n796 B.n3 163.367
R686 B.n792 B.n3 163.367
R687 B.n792 B.n9 163.367
R688 B.n788 B.n9 163.367
R689 B.n788 B.n11 163.367
R690 B.n784 B.n11 163.367
R691 B.n784 B.n15 163.367
R692 B.n780 B.n15 163.367
R693 B.n780 B.n17 163.367
R694 B.n776 B.n17 163.367
R695 B.n776 B.n22 163.367
R696 B.n772 B.n22 163.367
R697 B.n772 B.n24 163.367
R698 B.n768 B.n24 163.367
R699 B.n768 B.n30 163.367
R700 B.n764 B.n30 163.367
R701 B.n764 B.n32 163.367
R702 B.n760 B.n32 163.367
R703 B.n760 B.n37 163.367
R704 B.n756 B.n37 163.367
R705 B.n756 B.n39 163.367
R706 B.n752 B.n39 163.367
R707 B.n752 B.n44 163.367
R708 B.n748 B.n44 163.367
R709 B.n748 B.n46 163.367
R710 B.n744 B.n46 163.367
R711 B.n744 B.n51 163.367
R712 B.n740 B.n51 163.367
R713 B.n740 B.n53 163.367
R714 B.n408 B.n407 163.367
R715 B.n599 B.n407 163.367
R716 B.n597 B.n596 163.367
R717 B.n593 B.n592 163.367
R718 B.n589 B.n588 163.367
R719 B.n585 B.n584 163.367
R720 B.n581 B.n580 163.367
R721 B.n577 B.n576 163.367
R722 B.n573 B.n572 163.367
R723 B.n569 B.n568 163.367
R724 B.n565 B.n564 163.367
R725 B.n561 B.n560 163.367
R726 B.n557 B.n556 163.367
R727 B.n553 B.n552 163.367
R728 B.n549 B.n548 163.367
R729 B.n545 B.n544 163.367
R730 B.n541 B.n540 163.367
R731 B.n537 B.n536 163.367
R732 B.n533 B.n532 163.367
R733 B.n529 B.n528 163.367
R734 B.n525 B.n524 163.367
R735 B.n521 B.n520 163.367
R736 B.n516 B.n515 163.367
R737 B.n512 B.n511 163.367
R738 B.n508 B.n507 163.367
R739 B.n504 B.n503 163.367
R740 B.n500 B.n499 163.367
R741 B.n495 B.n494 163.367
R742 B.n491 B.n490 163.367
R743 B.n487 B.n486 163.367
R744 B.n483 B.n482 163.367
R745 B.n479 B.n478 163.367
R746 B.n475 B.n474 163.367
R747 B.n471 B.n470 163.367
R748 B.n467 B.n466 163.367
R749 B.n463 B.n462 163.367
R750 B.n459 B.n458 163.367
R751 B.n455 B.n454 163.367
R752 B.n451 B.n450 163.367
R753 B.n447 B.n446 163.367
R754 B.n443 B.n442 163.367
R755 B.n439 B.n438 163.367
R756 B.n435 B.n434 163.367
R757 B.n431 B.n430 163.367
R758 B.n427 B.n426 163.367
R759 B.n423 B.n422 163.367
R760 B.n419 B.n418 163.367
R761 B.n415 B.n414 163.367
R762 B.n607 B.n359 163.367
R763 B.n611 B.n357 163.367
R764 B.n611 B.n350 163.367
R765 B.n619 B.n350 163.367
R766 B.n619 B.n348 163.367
R767 B.n623 B.n348 163.367
R768 B.n623 B.n343 163.367
R769 B.n631 B.n343 163.367
R770 B.n631 B.n341 163.367
R771 B.n635 B.n341 163.367
R772 B.n635 B.n335 163.367
R773 B.n643 B.n335 163.367
R774 B.n643 B.n333 163.367
R775 B.n647 B.n333 163.367
R776 B.n647 B.n327 163.367
R777 B.n655 B.n327 163.367
R778 B.n655 B.n325 163.367
R779 B.n659 B.n325 163.367
R780 B.n659 B.n320 163.367
R781 B.n668 B.n320 163.367
R782 B.n668 B.n318 163.367
R783 B.n672 B.n318 163.367
R784 B.n672 B.n313 163.367
R785 B.n681 B.n313 163.367
R786 B.n681 B.n311 163.367
R787 B.n686 B.n311 163.367
R788 B.n686 B.n305 163.367
R789 B.n694 B.n305 163.367
R790 B.n695 B.n694 163.367
R791 B.n695 B.n5 163.367
R792 B.n6 B.n5 163.367
R793 B.n7 B.n6 163.367
R794 B.n700 B.n7 163.367
R795 B.n700 B.n12 163.367
R796 B.n13 B.n12 163.367
R797 B.n14 B.n13 163.367
R798 B.n705 B.n14 163.367
R799 B.n705 B.n19 163.367
R800 B.n20 B.n19 163.367
R801 B.n21 B.n20 163.367
R802 B.n710 B.n21 163.367
R803 B.n710 B.n26 163.367
R804 B.n27 B.n26 163.367
R805 B.n28 B.n27 163.367
R806 B.n715 B.n28 163.367
R807 B.n715 B.n33 163.367
R808 B.n34 B.n33 163.367
R809 B.n35 B.n34 163.367
R810 B.n720 B.n35 163.367
R811 B.n720 B.n40 163.367
R812 B.n41 B.n40 163.367
R813 B.n42 B.n41 163.367
R814 B.n725 B.n42 163.367
R815 B.n725 B.n47 163.367
R816 B.n48 B.n47 163.367
R817 B.n49 B.n48 163.367
R818 B.n730 B.n49 163.367
R819 B.n730 B.n54 163.367
R820 B.n55 B.n54 163.367
R821 B.n115 B.n114 163.367
R822 B.n119 B.n118 163.367
R823 B.n123 B.n122 163.367
R824 B.n127 B.n126 163.367
R825 B.n131 B.n130 163.367
R826 B.n135 B.n134 163.367
R827 B.n139 B.n138 163.367
R828 B.n143 B.n142 163.367
R829 B.n147 B.n146 163.367
R830 B.n151 B.n150 163.367
R831 B.n155 B.n154 163.367
R832 B.n159 B.n158 163.367
R833 B.n163 B.n162 163.367
R834 B.n167 B.n166 163.367
R835 B.n171 B.n170 163.367
R836 B.n175 B.n174 163.367
R837 B.n179 B.n178 163.367
R838 B.n183 B.n182 163.367
R839 B.n187 B.n186 163.367
R840 B.n191 B.n190 163.367
R841 B.n195 B.n194 163.367
R842 B.n199 B.n198 163.367
R843 B.n203 B.n202 163.367
R844 B.n207 B.n206 163.367
R845 B.n211 B.n210 163.367
R846 B.n215 B.n214 163.367
R847 B.n219 B.n218 163.367
R848 B.n223 B.n222 163.367
R849 B.n227 B.n226 163.367
R850 B.n231 B.n230 163.367
R851 B.n235 B.n234 163.367
R852 B.n239 B.n238 163.367
R853 B.n243 B.n242 163.367
R854 B.n247 B.n246 163.367
R855 B.n251 B.n250 163.367
R856 B.n255 B.n254 163.367
R857 B.n259 B.n258 163.367
R858 B.n263 B.n262 163.367
R859 B.n267 B.n266 163.367
R860 B.n271 B.n270 163.367
R861 B.n275 B.n274 163.367
R862 B.n279 B.n278 163.367
R863 B.n283 B.n282 163.367
R864 B.n287 B.n286 163.367
R865 B.n291 B.n290 163.367
R866 B.n295 B.n294 163.367
R867 B.n299 B.n298 163.367
R868 B.n301 B.n104 163.367
R869 B.n411 B.t13 91.9104
R870 B.n105 B.t16 91.9104
R871 B.n409 B.t20 91.8937
R872 B.n108 B.t22 91.8937
R873 B.n606 B.n356 86.2159
R874 B.n738 B.n737 86.2159
R875 B.n605 B.n604 71.676
R876 B.n599 B.n360 71.676
R877 B.n596 B.n361 71.676
R878 B.n592 B.n362 71.676
R879 B.n588 B.n363 71.676
R880 B.n584 B.n364 71.676
R881 B.n580 B.n365 71.676
R882 B.n576 B.n366 71.676
R883 B.n572 B.n367 71.676
R884 B.n568 B.n368 71.676
R885 B.n564 B.n369 71.676
R886 B.n560 B.n370 71.676
R887 B.n556 B.n371 71.676
R888 B.n552 B.n372 71.676
R889 B.n548 B.n373 71.676
R890 B.n544 B.n374 71.676
R891 B.n540 B.n375 71.676
R892 B.n536 B.n376 71.676
R893 B.n532 B.n377 71.676
R894 B.n528 B.n378 71.676
R895 B.n524 B.n379 71.676
R896 B.n520 B.n380 71.676
R897 B.n515 B.n381 71.676
R898 B.n511 B.n382 71.676
R899 B.n507 B.n383 71.676
R900 B.n503 B.n384 71.676
R901 B.n499 B.n385 71.676
R902 B.n494 B.n386 71.676
R903 B.n490 B.n387 71.676
R904 B.n486 B.n388 71.676
R905 B.n482 B.n389 71.676
R906 B.n478 B.n390 71.676
R907 B.n474 B.n391 71.676
R908 B.n470 B.n392 71.676
R909 B.n466 B.n393 71.676
R910 B.n462 B.n394 71.676
R911 B.n458 B.n395 71.676
R912 B.n454 B.n396 71.676
R913 B.n450 B.n397 71.676
R914 B.n446 B.n398 71.676
R915 B.n442 B.n399 71.676
R916 B.n438 B.n400 71.676
R917 B.n434 B.n401 71.676
R918 B.n430 B.n402 71.676
R919 B.n426 B.n403 71.676
R920 B.n422 B.n404 71.676
R921 B.n418 B.n405 71.676
R922 B.n414 B.n406 71.676
R923 B.n111 B.n56 71.676
R924 B.n115 B.n57 71.676
R925 B.n119 B.n58 71.676
R926 B.n123 B.n59 71.676
R927 B.n127 B.n60 71.676
R928 B.n131 B.n61 71.676
R929 B.n135 B.n62 71.676
R930 B.n139 B.n63 71.676
R931 B.n143 B.n64 71.676
R932 B.n147 B.n65 71.676
R933 B.n151 B.n66 71.676
R934 B.n155 B.n67 71.676
R935 B.n159 B.n68 71.676
R936 B.n163 B.n69 71.676
R937 B.n167 B.n70 71.676
R938 B.n171 B.n71 71.676
R939 B.n175 B.n72 71.676
R940 B.n179 B.n73 71.676
R941 B.n183 B.n74 71.676
R942 B.n187 B.n75 71.676
R943 B.n191 B.n76 71.676
R944 B.n195 B.n77 71.676
R945 B.n199 B.n78 71.676
R946 B.n203 B.n79 71.676
R947 B.n207 B.n80 71.676
R948 B.n211 B.n81 71.676
R949 B.n215 B.n82 71.676
R950 B.n219 B.n83 71.676
R951 B.n223 B.n84 71.676
R952 B.n227 B.n85 71.676
R953 B.n231 B.n86 71.676
R954 B.n235 B.n87 71.676
R955 B.n239 B.n88 71.676
R956 B.n243 B.n89 71.676
R957 B.n247 B.n90 71.676
R958 B.n251 B.n91 71.676
R959 B.n255 B.n92 71.676
R960 B.n259 B.n93 71.676
R961 B.n263 B.n94 71.676
R962 B.n267 B.n95 71.676
R963 B.n271 B.n96 71.676
R964 B.n275 B.n97 71.676
R965 B.n279 B.n98 71.676
R966 B.n283 B.n99 71.676
R967 B.n287 B.n100 71.676
R968 B.n291 B.n101 71.676
R969 B.n295 B.n102 71.676
R970 B.n299 B.n103 71.676
R971 B.n736 B.n104 71.676
R972 B.n736 B.n735 71.676
R973 B.n301 B.n103 71.676
R974 B.n298 B.n102 71.676
R975 B.n294 B.n101 71.676
R976 B.n290 B.n100 71.676
R977 B.n286 B.n99 71.676
R978 B.n282 B.n98 71.676
R979 B.n278 B.n97 71.676
R980 B.n274 B.n96 71.676
R981 B.n270 B.n95 71.676
R982 B.n266 B.n94 71.676
R983 B.n262 B.n93 71.676
R984 B.n258 B.n92 71.676
R985 B.n254 B.n91 71.676
R986 B.n250 B.n90 71.676
R987 B.n246 B.n89 71.676
R988 B.n242 B.n88 71.676
R989 B.n238 B.n87 71.676
R990 B.n234 B.n86 71.676
R991 B.n230 B.n85 71.676
R992 B.n226 B.n84 71.676
R993 B.n222 B.n83 71.676
R994 B.n218 B.n82 71.676
R995 B.n214 B.n81 71.676
R996 B.n210 B.n80 71.676
R997 B.n206 B.n79 71.676
R998 B.n202 B.n78 71.676
R999 B.n198 B.n77 71.676
R1000 B.n194 B.n76 71.676
R1001 B.n190 B.n75 71.676
R1002 B.n186 B.n74 71.676
R1003 B.n182 B.n73 71.676
R1004 B.n178 B.n72 71.676
R1005 B.n174 B.n71 71.676
R1006 B.n170 B.n70 71.676
R1007 B.n166 B.n69 71.676
R1008 B.n162 B.n68 71.676
R1009 B.n158 B.n67 71.676
R1010 B.n154 B.n66 71.676
R1011 B.n150 B.n65 71.676
R1012 B.n146 B.n64 71.676
R1013 B.n142 B.n63 71.676
R1014 B.n138 B.n62 71.676
R1015 B.n134 B.n61 71.676
R1016 B.n130 B.n60 71.676
R1017 B.n126 B.n59 71.676
R1018 B.n122 B.n58 71.676
R1019 B.n118 B.n57 71.676
R1020 B.n114 B.n56 71.676
R1021 B.n605 B.n408 71.676
R1022 B.n597 B.n360 71.676
R1023 B.n593 B.n361 71.676
R1024 B.n589 B.n362 71.676
R1025 B.n585 B.n363 71.676
R1026 B.n581 B.n364 71.676
R1027 B.n577 B.n365 71.676
R1028 B.n573 B.n366 71.676
R1029 B.n569 B.n367 71.676
R1030 B.n565 B.n368 71.676
R1031 B.n561 B.n369 71.676
R1032 B.n557 B.n370 71.676
R1033 B.n553 B.n371 71.676
R1034 B.n549 B.n372 71.676
R1035 B.n545 B.n373 71.676
R1036 B.n541 B.n374 71.676
R1037 B.n537 B.n375 71.676
R1038 B.n533 B.n376 71.676
R1039 B.n529 B.n377 71.676
R1040 B.n525 B.n378 71.676
R1041 B.n521 B.n379 71.676
R1042 B.n516 B.n380 71.676
R1043 B.n512 B.n381 71.676
R1044 B.n508 B.n382 71.676
R1045 B.n504 B.n383 71.676
R1046 B.n500 B.n384 71.676
R1047 B.n495 B.n385 71.676
R1048 B.n491 B.n386 71.676
R1049 B.n487 B.n387 71.676
R1050 B.n483 B.n388 71.676
R1051 B.n479 B.n389 71.676
R1052 B.n475 B.n390 71.676
R1053 B.n471 B.n391 71.676
R1054 B.n467 B.n392 71.676
R1055 B.n463 B.n393 71.676
R1056 B.n459 B.n394 71.676
R1057 B.n455 B.n395 71.676
R1058 B.n451 B.n396 71.676
R1059 B.n447 B.n397 71.676
R1060 B.n443 B.n398 71.676
R1061 B.n439 B.n399 71.676
R1062 B.n435 B.n400 71.676
R1063 B.n431 B.n401 71.676
R1064 B.n427 B.n402 71.676
R1065 B.n423 B.n403 71.676
R1066 B.n419 B.n404 71.676
R1067 B.n415 B.n405 71.676
R1068 B.n406 B.n359 71.676
R1069 B.n412 B.t12 68.6377
R1070 B.n106 B.t17 68.6377
R1071 B.n410 B.t19 68.621
R1072 B.n109 B.t23 68.621
R1073 B.n497 B.n412 59.5399
R1074 B.n518 B.n410 59.5399
R1075 B.n110 B.n109 59.5399
R1076 B.n107 B.n106 59.5399
R1077 B.n612 B.n356 40.998
R1078 B.n612 B.n351 40.998
R1079 B.n618 B.n351 40.998
R1080 B.n618 B.n352 40.998
R1081 B.n624 B.n344 40.998
R1082 B.n630 B.n344 40.998
R1083 B.n630 B.n340 40.998
R1084 B.n636 B.n340 40.998
R1085 B.n636 B.n336 40.998
R1086 B.n642 B.n336 40.998
R1087 B.n648 B.n332 40.998
R1088 B.n648 B.n328 40.998
R1089 B.n654 B.n328 40.998
R1090 B.n661 B.n324 40.998
R1091 B.n661 B.n660 40.998
R1092 B.n667 B.n317 40.998
R1093 B.n674 B.n317 40.998
R1094 B.n674 B.n673 40.998
R1095 B.n680 B.n310 40.998
R1096 B.n687 B.n310 40.998
R1097 B.n693 B.n306 40.998
R1098 B.n693 B.n4 40.998
R1099 B.n795 B.n4 40.998
R1100 B.n795 B.n794 40.998
R1101 B.n794 B.n793 40.998
R1102 B.n793 B.n8 40.998
R1103 B.n787 B.n786 40.998
R1104 B.n786 B.n785 40.998
R1105 B.n779 B.n18 40.998
R1106 B.n779 B.n778 40.998
R1107 B.n778 B.n777 40.998
R1108 B.n771 B.n25 40.998
R1109 B.n771 B.n770 40.998
R1110 B.n769 B.n29 40.998
R1111 B.n763 B.n29 40.998
R1112 B.n763 B.n762 40.998
R1113 B.n761 B.n36 40.998
R1114 B.n755 B.n36 40.998
R1115 B.n755 B.n754 40.998
R1116 B.n754 B.n753 40.998
R1117 B.n753 B.n43 40.998
R1118 B.n747 B.n43 40.998
R1119 B.n746 B.n745 40.998
R1120 B.n745 B.n50 40.998
R1121 B.n739 B.n50 40.998
R1122 B.n739 B.n738 40.998
R1123 B.t8 B.n324 39.1893
R1124 B.n770 B.t4 39.1893
R1125 B.n112 B.n52 38.2444
R1126 B.n734 B.n733 38.2444
R1127 B.n609 B.n608 38.2444
R1128 B.n603 B.n354 38.2444
R1129 B.n680 B.t9 36.7777
R1130 B.n785 B.t5 36.7777
R1131 B.n352 B.t11 31.9545
R1132 B.t15 B.n746 31.9545
R1133 B.n687 B.t7 25.9254
R1134 B.n787 B.t0 25.9254
R1135 B.n660 B.t1 23.5138
R1136 B.n25 B.t2 23.5138
R1137 B.n412 B.n411 23.2732
R1138 B.n410 B.n409 23.2732
R1139 B.n109 B.n108 23.2732
R1140 B.n106 B.n105 23.2732
R1141 B.n642 B.t6 21.1022
R1142 B.t3 B.n761 21.1022
R1143 B.t6 B.n332 19.8964
R1144 B.n762 B.t3 19.8964
R1145 B B.n797 18.0485
R1146 B.n667 B.t1 17.4847
R1147 B.n777 B.t2 17.4847
R1148 B.t7 B.n306 15.0731
R1149 B.t0 B.n8 15.0731
R1150 B.n113 B.n112 10.6151
R1151 B.n116 B.n113 10.6151
R1152 B.n117 B.n116 10.6151
R1153 B.n120 B.n117 10.6151
R1154 B.n121 B.n120 10.6151
R1155 B.n124 B.n121 10.6151
R1156 B.n125 B.n124 10.6151
R1157 B.n128 B.n125 10.6151
R1158 B.n129 B.n128 10.6151
R1159 B.n132 B.n129 10.6151
R1160 B.n133 B.n132 10.6151
R1161 B.n136 B.n133 10.6151
R1162 B.n137 B.n136 10.6151
R1163 B.n140 B.n137 10.6151
R1164 B.n141 B.n140 10.6151
R1165 B.n144 B.n141 10.6151
R1166 B.n145 B.n144 10.6151
R1167 B.n148 B.n145 10.6151
R1168 B.n149 B.n148 10.6151
R1169 B.n152 B.n149 10.6151
R1170 B.n153 B.n152 10.6151
R1171 B.n156 B.n153 10.6151
R1172 B.n157 B.n156 10.6151
R1173 B.n160 B.n157 10.6151
R1174 B.n161 B.n160 10.6151
R1175 B.n164 B.n161 10.6151
R1176 B.n165 B.n164 10.6151
R1177 B.n168 B.n165 10.6151
R1178 B.n169 B.n168 10.6151
R1179 B.n172 B.n169 10.6151
R1180 B.n173 B.n172 10.6151
R1181 B.n176 B.n173 10.6151
R1182 B.n177 B.n176 10.6151
R1183 B.n180 B.n177 10.6151
R1184 B.n181 B.n180 10.6151
R1185 B.n184 B.n181 10.6151
R1186 B.n185 B.n184 10.6151
R1187 B.n188 B.n185 10.6151
R1188 B.n189 B.n188 10.6151
R1189 B.n192 B.n189 10.6151
R1190 B.n193 B.n192 10.6151
R1191 B.n196 B.n193 10.6151
R1192 B.n197 B.n196 10.6151
R1193 B.n201 B.n200 10.6151
R1194 B.n204 B.n201 10.6151
R1195 B.n205 B.n204 10.6151
R1196 B.n208 B.n205 10.6151
R1197 B.n209 B.n208 10.6151
R1198 B.n212 B.n209 10.6151
R1199 B.n213 B.n212 10.6151
R1200 B.n216 B.n213 10.6151
R1201 B.n217 B.n216 10.6151
R1202 B.n221 B.n220 10.6151
R1203 B.n224 B.n221 10.6151
R1204 B.n225 B.n224 10.6151
R1205 B.n228 B.n225 10.6151
R1206 B.n229 B.n228 10.6151
R1207 B.n232 B.n229 10.6151
R1208 B.n233 B.n232 10.6151
R1209 B.n236 B.n233 10.6151
R1210 B.n237 B.n236 10.6151
R1211 B.n240 B.n237 10.6151
R1212 B.n241 B.n240 10.6151
R1213 B.n244 B.n241 10.6151
R1214 B.n245 B.n244 10.6151
R1215 B.n248 B.n245 10.6151
R1216 B.n249 B.n248 10.6151
R1217 B.n252 B.n249 10.6151
R1218 B.n253 B.n252 10.6151
R1219 B.n256 B.n253 10.6151
R1220 B.n257 B.n256 10.6151
R1221 B.n260 B.n257 10.6151
R1222 B.n261 B.n260 10.6151
R1223 B.n264 B.n261 10.6151
R1224 B.n265 B.n264 10.6151
R1225 B.n268 B.n265 10.6151
R1226 B.n269 B.n268 10.6151
R1227 B.n272 B.n269 10.6151
R1228 B.n273 B.n272 10.6151
R1229 B.n276 B.n273 10.6151
R1230 B.n277 B.n276 10.6151
R1231 B.n280 B.n277 10.6151
R1232 B.n281 B.n280 10.6151
R1233 B.n284 B.n281 10.6151
R1234 B.n285 B.n284 10.6151
R1235 B.n288 B.n285 10.6151
R1236 B.n289 B.n288 10.6151
R1237 B.n292 B.n289 10.6151
R1238 B.n293 B.n292 10.6151
R1239 B.n296 B.n293 10.6151
R1240 B.n297 B.n296 10.6151
R1241 B.n300 B.n297 10.6151
R1242 B.n302 B.n300 10.6151
R1243 B.n303 B.n302 10.6151
R1244 B.n734 B.n303 10.6151
R1245 B.n610 B.n609 10.6151
R1246 B.n610 B.n349 10.6151
R1247 B.n620 B.n349 10.6151
R1248 B.n621 B.n620 10.6151
R1249 B.n622 B.n621 10.6151
R1250 B.n622 B.n342 10.6151
R1251 B.n632 B.n342 10.6151
R1252 B.n633 B.n632 10.6151
R1253 B.n634 B.n633 10.6151
R1254 B.n634 B.n334 10.6151
R1255 B.n644 B.n334 10.6151
R1256 B.n645 B.n644 10.6151
R1257 B.n646 B.n645 10.6151
R1258 B.n646 B.n326 10.6151
R1259 B.n656 B.n326 10.6151
R1260 B.n657 B.n656 10.6151
R1261 B.n658 B.n657 10.6151
R1262 B.n658 B.n319 10.6151
R1263 B.n669 B.n319 10.6151
R1264 B.n670 B.n669 10.6151
R1265 B.n671 B.n670 10.6151
R1266 B.n671 B.n312 10.6151
R1267 B.n682 B.n312 10.6151
R1268 B.n683 B.n682 10.6151
R1269 B.n685 B.n683 10.6151
R1270 B.n685 B.n684 10.6151
R1271 B.n684 B.n304 10.6151
R1272 B.n696 B.n304 10.6151
R1273 B.n697 B.n696 10.6151
R1274 B.n698 B.n697 10.6151
R1275 B.n699 B.n698 10.6151
R1276 B.n701 B.n699 10.6151
R1277 B.n702 B.n701 10.6151
R1278 B.n703 B.n702 10.6151
R1279 B.n704 B.n703 10.6151
R1280 B.n706 B.n704 10.6151
R1281 B.n707 B.n706 10.6151
R1282 B.n708 B.n707 10.6151
R1283 B.n709 B.n708 10.6151
R1284 B.n711 B.n709 10.6151
R1285 B.n712 B.n711 10.6151
R1286 B.n713 B.n712 10.6151
R1287 B.n714 B.n713 10.6151
R1288 B.n716 B.n714 10.6151
R1289 B.n717 B.n716 10.6151
R1290 B.n718 B.n717 10.6151
R1291 B.n719 B.n718 10.6151
R1292 B.n721 B.n719 10.6151
R1293 B.n722 B.n721 10.6151
R1294 B.n723 B.n722 10.6151
R1295 B.n724 B.n723 10.6151
R1296 B.n726 B.n724 10.6151
R1297 B.n727 B.n726 10.6151
R1298 B.n728 B.n727 10.6151
R1299 B.n729 B.n728 10.6151
R1300 B.n731 B.n729 10.6151
R1301 B.n732 B.n731 10.6151
R1302 B.n733 B.n732 10.6151
R1303 B.n603 B.n602 10.6151
R1304 B.n602 B.n601 10.6151
R1305 B.n601 B.n600 10.6151
R1306 B.n600 B.n598 10.6151
R1307 B.n598 B.n595 10.6151
R1308 B.n595 B.n594 10.6151
R1309 B.n594 B.n591 10.6151
R1310 B.n591 B.n590 10.6151
R1311 B.n590 B.n587 10.6151
R1312 B.n587 B.n586 10.6151
R1313 B.n586 B.n583 10.6151
R1314 B.n583 B.n582 10.6151
R1315 B.n582 B.n579 10.6151
R1316 B.n579 B.n578 10.6151
R1317 B.n578 B.n575 10.6151
R1318 B.n575 B.n574 10.6151
R1319 B.n574 B.n571 10.6151
R1320 B.n571 B.n570 10.6151
R1321 B.n570 B.n567 10.6151
R1322 B.n567 B.n566 10.6151
R1323 B.n566 B.n563 10.6151
R1324 B.n563 B.n562 10.6151
R1325 B.n562 B.n559 10.6151
R1326 B.n559 B.n558 10.6151
R1327 B.n558 B.n555 10.6151
R1328 B.n555 B.n554 10.6151
R1329 B.n554 B.n551 10.6151
R1330 B.n551 B.n550 10.6151
R1331 B.n550 B.n547 10.6151
R1332 B.n547 B.n546 10.6151
R1333 B.n546 B.n543 10.6151
R1334 B.n543 B.n542 10.6151
R1335 B.n542 B.n539 10.6151
R1336 B.n539 B.n538 10.6151
R1337 B.n538 B.n535 10.6151
R1338 B.n535 B.n534 10.6151
R1339 B.n534 B.n531 10.6151
R1340 B.n531 B.n530 10.6151
R1341 B.n530 B.n527 10.6151
R1342 B.n527 B.n526 10.6151
R1343 B.n526 B.n523 10.6151
R1344 B.n523 B.n522 10.6151
R1345 B.n522 B.n519 10.6151
R1346 B.n517 B.n514 10.6151
R1347 B.n514 B.n513 10.6151
R1348 B.n513 B.n510 10.6151
R1349 B.n510 B.n509 10.6151
R1350 B.n509 B.n506 10.6151
R1351 B.n506 B.n505 10.6151
R1352 B.n505 B.n502 10.6151
R1353 B.n502 B.n501 10.6151
R1354 B.n501 B.n498 10.6151
R1355 B.n496 B.n493 10.6151
R1356 B.n493 B.n492 10.6151
R1357 B.n492 B.n489 10.6151
R1358 B.n489 B.n488 10.6151
R1359 B.n488 B.n485 10.6151
R1360 B.n485 B.n484 10.6151
R1361 B.n484 B.n481 10.6151
R1362 B.n481 B.n480 10.6151
R1363 B.n480 B.n477 10.6151
R1364 B.n477 B.n476 10.6151
R1365 B.n476 B.n473 10.6151
R1366 B.n473 B.n472 10.6151
R1367 B.n472 B.n469 10.6151
R1368 B.n469 B.n468 10.6151
R1369 B.n468 B.n465 10.6151
R1370 B.n465 B.n464 10.6151
R1371 B.n464 B.n461 10.6151
R1372 B.n461 B.n460 10.6151
R1373 B.n460 B.n457 10.6151
R1374 B.n457 B.n456 10.6151
R1375 B.n456 B.n453 10.6151
R1376 B.n453 B.n452 10.6151
R1377 B.n452 B.n449 10.6151
R1378 B.n449 B.n448 10.6151
R1379 B.n448 B.n445 10.6151
R1380 B.n445 B.n444 10.6151
R1381 B.n444 B.n441 10.6151
R1382 B.n441 B.n440 10.6151
R1383 B.n440 B.n437 10.6151
R1384 B.n437 B.n436 10.6151
R1385 B.n436 B.n433 10.6151
R1386 B.n433 B.n432 10.6151
R1387 B.n432 B.n429 10.6151
R1388 B.n429 B.n428 10.6151
R1389 B.n428 B.n425 10.6151
R1390 B.n425 B.n424 10.6151
R1391 B.n424 B.n421 10.6151
R1392 B.n421 B.n420 10.6151
R1393 B.n420 B.n417 10.6151
R1394 B.n417 B.n416 10.6151
R1395 B.n416 B.n413 10.6151
R1396 B.n413 B.n358 10.6151
R1397 B.n608 B.n358 10.6151
R1398 B.n614 B.n354 10.6151
R1399 B.n615 B.n614 10.6151
R1400 B.n616 B.n615 10.6151
R1401 B.n616 B.n346 10.6151
R1402 B.n626 B.n346 10.6151
R1403 B.n627 B.n626 10.6151
R1404 B.n628 B.n627 10.6151
R1405 B.n628 B.n338 10.6151
R1406 B.n638 B.n338 10.6151
R1407 B.n639 B.n638 10.6151
R1408 B.n640 B.n639 10.6151
R1409 B.n640 B.n330 10.6151
R1410 B.n650 B.n330 10.6151
R1411 B.n651 B.n650 10.6151
R1412 B.n652 B.n651 10.6151
R1413 B.n652 B.n322 10.6151
R1414 B.n663 B.n322 10.6151
R1415 B.n664 B.n663 10.6151
R1416 B.n665 B.n664 10.6151
R1417 B.n665 B.n315 10.6151
R1418 B.n676 B.n315 10.6151
R1419 B.n677 B.n676 10.6151
R1420 B.n678 B.n677 10.6151
R1421 B.n678 B.n308 10.6151
R1422 B.n689 B.n308 10.6151
R1423 B.n690 B.n689 10.6151
R1424 B.n691 B.n690 10.6151
R1425 B.n691 B.n0 10.6151
R1426 B.n791 B.n1 10.6151
R1427 B.n791 B.n790 10.6151
R1428 B.n790 B.n789 10.6151
R1429 B.n789 B.n10 10.6151
R1430 B.n783 B.n10 10.6151
R1431 B.n783 B.n782 10.6151
R1432 B.n782 B.n781 10.6151
R1433 B.n781 B.n16 10.6151
R1434 B.n775 B.n16 10.6151
R1435 B.n775 B.n774 10.6151
R1436 B.n774 B.n773 10.6151
R1437 B.n773 B.n23 10.6151
R1438 B.n767 B.n23 10.6151
R1439 B.n767 B.n766 10.6151
R1440 B.n766 B.n765 10.6151
R1441 B.n765 B.n31 10.6151
R1442 B.n759 B.n31 10.6151
R1443 B.n759 B.n758 10.6151
R1444 B.n758 B.n757 10.6151
R1445 B.n757 B.n38 10.6151
R1446 B.n751 B.n38 10.6151
R1447 B.n751 B.n750 10.6151
R1448 B.n750 B.n749 10.6151
R1449 B.n749 B.n45 10.6151
R1450 B.n743 B.n45 10.6151
R1451 B.n743 B.n742 10.6151
R1452 B.n742 B.n741 10.6151
R1453 B.n741 B.n52 10.6151
R1454 B.n197 B.n110 9.36635
R1455 B.n220 B.n107 9.36635
R1456 B.n519 B.n518 9.36635
R1457 B.n497 B.n496 9.36635
R1458 B.n624 B.t11 9.04407
R1459 B.n747 B.t15 9.04407
R1460 B.n673 B.t9 4.22083
R1461 B.n18 B.t5 4.22083
R1462 B.n797 B.n0 2.81026
R1463 B.n797 B.n1 2.81026
R1464 B.n654 B.t8 1.80921
R1465 B.t4 B.n769 1.80921
R1466 B.n200 B.n110 1.24928
R1467 B.n217 B.n107 1.24928
R1468 B.n518 B.n517 1.24928
R1469 B.n498 B.n497 1.24928
R1470 VP.n8 VP.t7 419.642
R1471 VP.n22 VP.t2 404.714
R1472 VP.n35 VP.t5 404.714
R1473 VP.n19 VP.t3 404.714
R1474 VP.n28 VP.t6 359.284
R1475 VP.n3 VP.t1 359.284
R1476 VP.n33 VP.t0 359.284
R1477 VP.n12 VP.t4 359.284
R1478 VP.n17 VP.t8 359.284
R1479 VP.n7 VP.t9 359.284
R1480 VP.n10 VP.n9 161.3
R1481 VP.n11 VP.n6 161.3
R1482 VP.n13 VP.n12 161.3
R1483 VP.n14 VP.n5 161.3
R1484 VP.n16 VP.n15 161.3
R1485 VP.n18 VP.n4 161.3
R1486 VP.n34 VP.n0 161.3
R1487 VP.n32 VP.n31 161.3
R1488 VP.n30 VP.n1 161.3
R1489 VP.n29 VP.n28 161.3
R1490 VP.n27 VP.n2 161.3
R1491 VP.n26 VP.n25 161.3
R1492 VP.n24 VP.n23 161.3
R1493 VP.n20 VP.n19 80.6037
R1494 VP.n36 VP.n35 80.6037
R1495 VP.n22 VP.n21 80.6037
R1496 VP.n23 VP.n22 54.8066
R1497 VP.n35 VP.n34 54.8066
R1498 VP.n19 VP.n18 54.8066
R1499 VP.n27 VP.n26 50.2061
R1500 VP.n32 VP.n1 50.2061
R1501 VP.n16 VP.n5 50.2061
R1502 VP.n11 VP.n10 50.2061
R1503 VP.n21 VP.n20 44.5544
R1504 VP.n8 VP.n7 44.4469
R1505 VP.n9 VP.n8 44.1212
R1506 VP.n28 VP.n27 30.7807
R1507 VP.n28 VP.n1 30.7807
R1508 VP.n12 VP.n5 30.7807
R1509 VP.n12 VP.n11 30.7807
R1510 VP.n23 VP.n3 14.6807
R1511 VP.n34 VP.n33 14.6807
R1512 VP.n18 VP.n17 14.6807
R1513 VP.n26 VP.n3 9.7873
R1514 VP.n33 VP.n32 9.7873
R1515 VP.n17 VP.n16 9.7873
R1516 VP.n10 VP.n7 9.7873
R1517 VP.n20 VP.n4 0.285035
R1518 VP.n24 VP.n21 0.285035
R1519 VP.n36 VP.n0 0.285035
R1520 VP.n9 VP.n6 0.189894
R1521 VP.n13 VP.n6 0.189894
R1522 VP.n14 VP.n13 0.189894
R1523 VP.n15 VP.n14 0.189894
R1524 VP.n15 VP.n4 0.189894
R1525 VP.n25 VP.n24 0.189894
R1526 VP.n25 VP.n2 0.189894
R1527 VP.n29 VP.n2 0.189894
R1528 VP.n30 VP.n29 0.189894
R1529 VP.n31 VP.n30 0.189894
R1530 VP.n31 VP.n0 0.189894
R1531 VP VP.n36 0.146778
R1532 VDD1.n1 VDD1.t2 66.2592
R1533 VDD1.n3 VDD1.t7 66.2581
R1534 VDD1.n5 VDD1.n4 64.4175
R1535 VDD1.n1 VDD1.n0 63.6982
R1536 VDD1.n7 VDD1.n6 63.697
R1537 VDD1.n3 VDD1.n2 63.697
R1538 VDD1.n7 VDD1.n5 40.9104
R1539 VDD1.n6 VDD1.t1 1.5271
R1540 VDD1.n6 VDD1.t6 1.5271
R1541 VDD1.n0 VDD1.t0 1.5271
R1542 VDD1.n0 VDD1.t5 1.5271
R1543 VDD1.n4 VDD1.t9 1.5271
R1544 VDD1.n4 VDD1.t4 1.5271
R1545 VDD1.n2 VDD1.t8 1.5271
R1546 VDD1.n2 VDD1.t3 1.5271
R1547 VDD1 VDD1.n7 0.718172
R1548 VDD1 VDD1.n1 0.31731
R1549 VDD1.n5 VDD1.n3 0.203775
C0 VDD1 VP 8.232961f
C1 VN VP 6.03088f
C2 VDD2 VP 0.363335f
C3 VDD1 VTAIL 13.811999f
C4 VN VTAIL 7.901609f
C5 VDD2 VTAIL 13.847401f
C6 VN VDD1 0.149412f
C7 VDD2 VDD1 1.07949f
C8 VTAIL VP 7.91621f
C9 VDD2 VN 8.02388f
C10 VDD2 B 5.336816f
C11 VDD1 B 5.282138f
C12 VTAIL B 7.045303f
C13 VN B 10.317441f
C14 VP B 8.407204f
C15 VDD1.t2 B 2.79034f
C16 VDD1.t0 B 0.242995f
C17 VDD1.t5 B 0.242995f
C18 VDD1.n0 B 2.18326f
C19 VDD1.n1 B 0.625852f
C20 VDD1.t7 B 2.79033f
C21 VDD1.t8 B 0.242995f
C22 VDD1.t3 B 0.242995f
C23 VDD1.n2 B 2.18325f
C24 VDD1.n3 B 0.6199f
C25 VDD1.t9 B 0.242995f
C26 VDD1.t4 B 0.242995f
C27 VDD1.n4 B 2.18699f
C28 VDD1.n5 B 2.01858f
C29 VDD1.t1 B 0.242995f
C30 VDD1.t6 B 0.242995f
C31 VDD1.n6 B 2.18325f
C32 VDD1.n7 B 2.39525f
C33 VP.n0 B 0.052602f
C34 VP.t0 B 1.21456f
C35 VP.n1 B 0.03724f
C36 VP.n2 B 0.039421f
C37 VP.t6 B 1.21456f
C38 VP.t1 B 1.21456f
C39 VP.n3 B 0.451805f
C40 VP.n4 B 0.052602f
C41 VP.t3 B 1.2671f
C42 VP.t8 B 1.21456f
C43 VP.n5 B 0.03724f
C44 VP.n6 B 0.039421f
C45 VP.t4 B 1.21456f
C46 VP.t9 B 1.21456f
C47 VP.n7 B 0.484049f
C48 VP.t7 B 1.28494f
C49 VP.n8 B 0.50007f
C50 VP.n9 B 0.161046f
C51 VP.n10 B 0.050588f
C52 VP.n11 B 0.03724f
C53 VP.n12 B 0.500009f
C54 VP.n13 B 0.039421f
C55 VP.n14 B 0.039421f
C56 VP.n15 B 0.039421f
C57 VP.n16 B 0.050588f
C58 VP.n17 B 0.451805f
C59 VP.n18 B 0.048146f
C60 VP.n19 B 0.501237f
C61 VP.n20 B 1.80607f
C62 VP.n21 B 1.83788f
C63 VP.t2 B 1.2671f
C64 VP.n22 B 0.501237f
C65 VP.n23 B 0.048146f
C66 VP.n24 B 0.052602f
C67 VP.n25 B 0.039421f
C68 VP.n26 B 0.050588f
C69 VP.n27 B 0.03724f
C70 VP.n28 B 0.500009f
C71 VP.n29 B 0.039421f
C72 VP.n30 B 0.039421f
C73 VP.n31 B 0.039421f
C74 VP.n32 B 0.050588f
C75 VP.n33 B 0.451805f
C76 VP.n34 B 0.048146f
C77 VP.t5 B 1.2671f
C78 VP.n35 B 0.501237f
C79 VP.n36 B 0.036919f
C80 VTAIL.t10 B 0.254939f
C81 VTAIL.t12 B 0.254939f
C82 VTAIL.n0 B 2.22182f
C83 VTAIL.n1 B 0.379402f
C84 VTAIL.t7 B 2.83339f
C85 VTAIL.n2 B 0.479188f
C86 VTAIL.t1 B 0.254939f
C87 VTAIL.t9 B 0.254939f
C88 VTAIL.n3 B 2.22182f
C89 VTAIL.n4 B 0.399267f
C90 VTAIL.t6 B 0.254939f
C91 VTAIL.t8 B 0.254939f
C92 VTAIL.n5 B 2.22182f
C93 VTAIL.n6 B 1.71621f
C94 VTAIL.t11 B 0.254939f
C95 VTAIL.t18 B 0.254939f
C96 VTAIL.n7 B 2.22183f
C97 VTAIL.n8 B 1.7162f
C98 VTAIL.t14 B 0.254939f
C99 VTAIL.t19 B 0.254939f
C100 VTAIL.n9 B 2.22183f
C101 VTAIL.n10 B 0.399256f
C102 VTAIL.t15 B 2.83341f
C103 VTAIL.n11 B 0.479171f
C104 VTAIL.t0 B 0.254939f
C105 VTAIL.t5 B 0.254939f
C106 VTAIL.n12 B 2.22183f
C107 VTAIL.n13 B 0.395456f
C108 VTAIL.t2 B 0.254939f
C109 VTAIL.t4 B 0.254939f
C110 VTAIL.n14 B 2.22183f
C111 VTAIL.n15 B 0.399256f
C112 VTAIL.t3 B 2.83339f
C113 VTAIL.n16 B 1.71702f
C114 VTAIL.t17 B 2.83339f
C115 VTAIL.n17 B 1.71702f
C116 VTAIL.t16 B 0.254939f
C117 VTAIL.t13 B 0.254939f
C118 VTAIL.n18 B 2.22182f
C119 VTAIL.n19 B 0.332418f
C120 VDD2.t5 B 2.77601f
C121 VDD2.t8 B 0.241749f
C122 VDD2.t3 B 0.241749f
C123 VDD2.n0 B 2.17205f
C124 VDD2.n1 B 0.616719f
C125 VDD2.t9 B 0.241749f
C126 VDD2.t2 B 0.241749f
C127 VDD2.n2 B 2.17576f
C128 VDD2.n3 B 1.93146f
C129 VDD2.t0 B 2.77076f
C130 VDD2.n4 B 2.37866f
C131 VDD2.t7 B 0.241749f
C132 VDD2.t1 B 0.241749f
C133 VDD2.n5 B 2.17206f
C134 VDD2.n6 B 0.290935f
C135 VDD2.t4 B 0.241749f
C136 VDD2.t6 B 0.241749f
C137 VDD2.n7 B 2.17574f
C138 VN.n0 B 0.051996f
C139 VN.t6 B 1.20056f
C140 VN.n1 B 0.036811f
C141 VN.n2 B 0.038966f
C142 VN.t3 B 1.20056f
C143 VN.t7 B 1.20056f
C144 VN.n3 B 0.478469f
C145 VN.t9 B 1.27013f
C146 VN.n4 B 0.494306f
C147 VN.n5 B 0.159189f
C148 VN.n6 B 0.050005f
C149 VN.n7 B 0.036811f
C150 VN.n8 B 0.494245f
C151 VN.n9 B 0.038966f
C152 VN.n10 B 0.038966f
C153 VN.n11 B 0.038966f
C154 VN.n12 B 0.050005f
C155 VN.n13 B 0.446597f
C156 VN.n14 B 0.047591f
C157 VN.t2 B 1.25249f
C158 VN.n15 B 0.495459f
C159 VN.n16 B 0.036494f
C160 VN.n17 B 0.051996f
C161 VN.t1 B 1.20056f
C162 VN.n18 B 0.036811f
C163 VN.n19 B 0.038966f
C164 VN.t5 B 1.20056f
C165 VN.t0 B 1.20056f
C166 VN.n20 B 0.478469f
C167 VN.t4 B 1.27013f
C168 VN.n21 B 0.494306f
C169 VN.n22 B 0.159189f
C170 VN.n23 B 0.050005f
C171 VN.n24 B 0.036811f
C172 VN.n25 B 0.494245f
C173 VN.n26 B 0.038966f
C174 VN.n27 B 0.038966f
C175 VN.n28 B 0.038966f
C176 VN.n29 B 0.050005f
C177 VN.n30 B 0.446597f
C178 VN.n31 B 0.047591f
C179 VN.t8 B 1.25249f
C180 VN.n32 B 0.495459f
C181 VN.n33 B 1.80689f
.ends

