* NGSPICE file created from diff_pair_sample_0705.ext - technology: sky130A

.subckt diff_pair_sample_0705 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=2.21925 pd=13.78 as=5.2455 ps=27.68 w=13.45 l=3.96
X1 B.t11 B.t9 B.t10 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=0 ps=0 w=13.45 l=3.96
X2 VDD1.t2 VP.t1 VTAIL.t4 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=2.21925 pd=13.78 as=5.2455 ps=27.68 w=13.45 l=3.96
X3 VTAIL.t2 VN.t0 VDD2.t3 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=2.21925 ps=13.78 w=13.45 l=3.96
X4 VDD2.t2 VN.t1 VTAIL.t0 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=2.21925 pd=13.78 as=5.2455 ps=27.68 w=13.45 l=3.96
X5 B.t8 B.t6 B.t7 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=0 ps=0 w=13.45 l=3.96
X6 VTAIL.t3 VN.t2 VDD2.t1 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=2.21925 ps=13.78 w=13.45 l=3.96
X7 B.t5 B.t3 B.t4 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=0 ps=0 w=13.45 l=3.96
X8 VTAIL.t5 VP.t2 VDD1.t1 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=2.21925 ps=13.78 w=13.45 l=3.96
X9 B.t2 B.t0 B.t1 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=0 ps=0 w=13.45 l=3.96
X10 VTAIL.t7 VP.t3 VDD1.t0 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=5.2455 pd=27.68 as=2.21925 ps=13.78 w=13.45 l=3.96
X11 VDD2.t0 VN.t3 VTAIL.t1 w_n3544_n3658# sky130_fd_pr__pfet_01v8 ad=2.21925 pd=13.78 as=5.2455 ps=27.68 w=13.45 l=3.96
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t2 115.666
R9 VP.n4 VP.t1 114.231
R10 VP.n6 VP.t3 81.8553
R11 VP.n19 VP.t0 81.8553
R12 VP.n6 VP.n5 62.8529
R13 VP.n20 VP.n19 62.8529
R14 VP.n13 VP.n12 56.5193
R15 VP.n5 VP.n4 53.444
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 19.3294
R23 VP.n19 VP.n18 19.3294
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n586 VTAIL.n518 756.745
R35 VTAIL.n68 VTAIL.n0 756.745
R36 VTAIL.n142 VTAIL.n74 756.745
R37 VTAIL.n216 VTAIL.n148 756.745
R38 VTAIL.n512 VTAIL.n444 756.745
R39 VTAIL.n438 VTAIL.n370 756.745
R40 VTAIL.n364 VTAIL.n296 756.745
R41 VTAIL.n290 VTAIL.n222 756.745
R42 VTAIL.n543 VTAIL.n542 585
R43 VTAIL.n545 VTAIL.n544 585
R44 VTAIL.n538 VTAIL.n537 585
R45 VTAIL.n551 VTAIL.n550 585
R46 VTAIL.n553 VTAIL.n552 585
R47 VTAIL.n534 VTAIL.n533 585
R48 VTAIL.n560 VTAIL.n559 585
R49 VTAIL.n561 VTAIL.n532 585
R50 VTAIL.n563 VTAIL.n562 585
R51 VTAIL.n530 VTAIL.n529 585
R52 VTAIL.n569 VTAIL.n568 585
R53 VTAIL.n571 VTAIL.n570 585
R54 VTAIL.n526 VTAIL.n525 585
R55 VTAIL.n577 VTAIL.n576 585
R56 VTAIL.n579 VTAIL.n578 585
R57 VTAIL.n522 VTAIL.n521 585
R58 VTAIL.n585 VTAIL.n584 585
R59 VTAIL.n587 VTAIL.n586 585
R60 VTAIL.n25 VTAIL.n24 585
R61 VTAIL.n27 VTAIL.n26 585
R62 VTAIL.n20 VTAIL.n19 585
R63 VTAIL.n33 VTAIL.n32 585
R64 VTAIL.n35 VTAIL.n34 585
R65 VTAIL.n16 VTAIL.n15 585
R66 VTAIL.n42 VTAIL.n41 585
R67 VTAIL.n43 VTAIL.n14 585
R68 VTAIL.n45 VTAIL.n44 585
R69 VTAIL.n12 VTAIL.n11 585
R70 VTAIL.n51 VTAIL.n50 585
R71 VTAIL.n53 VTAIL.n52 585
R72 VTAIL.n8 VTAIL.n7 585
R73 VTAIL.n59 VTAIL.n58 585
R74 VTAIL.n61 VTAIL.n60 585
R75 VTAIL.n4 VTAIL.n3 585
R76 VTAIL.n67 VTAIL.n66 585
R77 VTAIL.n69 VTAIL.n68 585
R78 VTAIL.n99 VTAIL.n98 585
R79 VTAIL.n101 VTAIL.n100 585
R80 VTAIL.n94 VTAIL.n93 585
R81 VTAIL.n107 VTAIL.n106 585
R82 VTAIL.n109 VTAIL.n108 585
R83 VTAIL.n90 VTAIL.n89 585
R84 VTAIL.n116 VTAIL.n115 585
R85 VTAIL.n117 VTAIL.n88 585
R86 VTAIL.n119 VTAIL.n118 585
R87 VTAIL.n86 VTAIL.n85 585
R88 VTAIL.n125 VTAIL.n124 585
R89 VTAIL.n127 VTAIL.n126 585
R90 VTAIL.n82 VTAIL.n81 585
R91 VTAIL.n133 VTAIL.n132 585
R92 VTAIL.n135 VTAIL.n134 585
R93 VTAIL.n78 VTAIL.n77 585
R94 VTAIL.n141 VTAIL.n140 585
R95 VTAIL.n143 VTAIL.n142 585
R96 VTAIL.n173 VTAIL.n172 585
R97 VTAIL.n175 VTAIL.n174 585
R98 VTAIL.n168 VTAIL.n167 585
R99 VTAIL.n181 VTAIL.n180 585
R100 VTAIL.n183 VTAIL.n182 585
R101 VTAIL.n164 VTAIL.n163 585
R102 VTAIL.n190 VTAIL.n189 585
R103 VTAIL.n191 VTAIL.n162 585
R104 VTAIL.n193 VTAIL.n192 585
R105 VTAIL.n160 VTAIL.n159 585
R106 VTAIL.n199 VTAIL.n198 585
R107 VTAIL.n201 VTAIL.n200 585
R108 VTAIL.n156 VTAIL.n155 585
R109 VTAIL.n207 VTAIL.n206 585
R110 VTAIL.n209 VTAIL.n208 585
R111 VTAIL.n152 VTAIL.n151 585
R112 VTAIL.n215 VTAIL.n214 585
R113 VTAIL.n217 VTAIL.n216 585
R114 VTAIL.n513 VTAIL.n512 585
R115 VTAIL.n511 VTAIL.n510 585
R116 VTAIL.n448 VTAIL.n447 585
R117 VTAIL.n505 VTAIL.n504 585
R118 VTAIL.n503 VTAIL.n502 585
R119 VTAIL.n452 VTAIL.n451 585
R120 VTAIL.n497 VTAIL.n496 585
R121 VTAIL.n495 VTAIL.n494 585
R122 VTAIL.n456 VTAIL.n455 585
R123 VTAIL.n460 VTAIL.n458 585
R124 VTAIL.n489 VTAIL.n488 585
R125 VTAIL.n487 VTAIL.n486 585
R126 VTAIL.n462 VTAIL.n461 585
R127 VTAIL.n481 VTAIL.n480 585
R128 VTAIL.n479 VTAIL.n478 585
R129 VTAIL.n466 VTAIL.n465 585
R130 VTAIL.n473 VTAIL.n472 585
R131 VTAIL.n471 VTAIL.n470 585
R132 VTAIL.n439 VTAIL.n438 585
R133 VTAIL.n437 VTAIL.n436 585
R134 VTAIL.n374 VTAIL.n373 585
R135 VTAIL.n431 VTAIL.n430 585
R136 VTAIL.n429 VTAIL.n428 585
R137 VTAIL.n378 VTAIL.n377 585
R138 VTAIL.n423 VTAIL.n422 585
R139 VTAIL.n421 VTAIL.n420 585
R140 VTAIL.n382 VTAIL.n381 585
R141 VTAIL.n386 VTAIL.n384 585
R142 VTAIL.n415 VTAIL.n414 585
R143 VTAIL.n413 VTAIL.n412 585
R144 VTAIL.n388 VTAIL.n387 585
R145 VTAIL.n407 VTAIL.n406 585
R146 VTAIL.n405 VTAIL.n404 585
R147 VTAIL.n392 VTAIL.n391 585
R148 VTAIL.n399 VTAIL.n398 585
R149 VTAIL.n397 VTAIL.n396 585
R150 VTAIL.n365 VTAIL.n364 585
R151 VTAIL.n363 VTAIL.n362 585
R152 VTAIL.n300 VTAIL.n299 585
R153 VTAIL.n357 VTAIL.n356 585
R154 VTAIL.n355 VTAIL.n354 585
R155 VTAIL.n304 VTAIL.n303 585
R156 VTAIL.n349 VTAIL.n348 585
R157 VTAIL.n347 VTAIL.n346 585
R158 VTAIL.n308 VTAIL.n307 585
R159 VTAIL.n312 VTAIL.n310 585
R160 VTAIL.n341 VTAIL.n340 585
R161 VTAIL.n339 VTAIL.n338 585
R162 VTAIL.n314 VTAIL.n313 585
R163 VTAIL.n333 VTAIL.n332 585
R164 VTAIL.n331 VTAIL.n330 585
R165 VTAIL.n318 VTAIL.n317 585
R166 VTAIL.n325 VTAIL.n324 585
R167 VTAIL.n323 VTAIL.n322 585
R168 VTAIL.n291 VTAIL.n290 585
R169 VTAIL.n289 VTAIL.n288 585
R170 VTAIL.n226 VTAIL.n225 585
R171 VTAIL.n283 VTAIL.n282 585
R172 VTAIL.n281 VTAIL.n280 585
R173 VTAIL.n230 VTAIL.n229 585
R174 VTAIL.n275 VTAIL.n274 585
R175 VTAIL.n273 VTAIL.n272 585
R176 VTAIL.n234 VTAIL.n233 585
R177 VTAIL.n238 VTAIL.n236 585
R178 VTAIL.n267 VTAIL.n266 585
R179 VTAIL.n265 VTAIL.n264 585
R180 VTAIL.n240 VTAIL.n239 585
R181 VTAIL.n259 VTAIL.n258 585
R182 VTAIL.n257 VTAIL.n256 585
R183 VTAIL.n244 VTAIL.n243 585
R184 VTAIL.n251 VTAIL.n250 585
R185 VTAIL.n249 VTAIL.n248 585
R186 VTAIL.n541 VTAIL.t1 329.036
R187 VTAIL.n23 VTAIL.t2 329.036
R188 VTAIL.n97 VTAIL.t6 329.036
R189 VTAIL.n171 VTAIL.t7 329.036
R190 VTAIL.n469 VTAIL.t4 329.036
R191 VTAIL.n395 VTAIL.t5 329.036
R192 VTAIL.n321 VTAIL.t0 329.036
R193 VTAIL.n247 VTAIL.t3 329.036
R194 VTAIL.n544 VTAIL.n543 171.744
R195 VTAIL.n544 VTAIL.n537 171.744
R196 VTAIL.n551 VTAIL.n537 171.744
R197 VTAIL.n552 VTAIL.n551 171.744
R198 VTAIL.n552 VTAIL.n533 171.744
R199 VTAIL.n560 VTAIL.n533 171.744
R200 VTAIL.n561 VTAIL.n560 171.744
R201 VTAIL.n562 VTAIL.n561 171.744
R202 VTAIL.n562 VTAIL.n529 171.744
R203 VTAIL.n569 VTAIL.n529 171.744
R204 VTAIL.n570 VTAIL.n569 171.744
R205 VTAIL.n570 VTAIL.n525 171.744
R206 VTAIL.n577 VTAIL.n525 171.744
R207 VTAIL.n578 VTAIL.n577 171.744
R208 VTAIL.n578 VTAIL.n521 171.744
R209 VTAIL.n585 VTAIL.n521 171.744
R210 VTAIL.n586 VTAIL.n585 171.744
R211 VTAIL.n26 VTAIL.n25 171.744
R212 VTAIL.n26 VTAIL.n19 171.744
R213 VTAIL.n33 VTAIL.n19 171.744
R214 VTAIL.n34 VTAIL.n33 171.744
R215 VTAIL.n34 VTAIL.n15 171.744
R216 VTAIL.n42 VTAIL.n15 171.744
R217 VTAIL.n43 VTAIL.n42 171.744
R218 VTAIL.n44 VTAIL.n43 171.744
R219 VTAIL.n44 VTAIL.n11 171.744
R220 VTAIL.n51 VTAIL.n11 171.744
R221 VTAIL.n52 VTAIL.n51 171.744
R222 VTAIL.n52 VTAIL.n7 171.744
R223 VTAIL.n59 VTAIL.n7 171.744
R224 VTAIL.n60 VTAIL.n59 171.744
R225 VTAIL.n60 VTAIL.n3 171.744
R226 VTAIL.n67 VTAIL.n3 171.744
R227 VTAIL.n68 VTAIL.n67 171.744
R228 VTAIL.n100 VTAIL.n99 171.744
R229 VTAIL.n100 VTAIL.n93 171.744
R230 VTAIL.n107 VTAIL.n93 171.744
R231 VTAIL.n108 VTAIL.n107 171.744
R232 VTAIL.n108 VTAIL.n89 171.744
R233 VTAIL.n116 VTAIL.n89 171.744
R234 VTAIL.n117 VTAIL.n116 171.744
R235 VTAIL.n118 VTAIL.n117 171.744
R236 VTAIL.n118 VTAIL.n85 171.744
R237 VTAIL.n125 VTAIL.n85 171.744
R238 VTAIL.n126 VTAIL.n125 171.744
R239 VTAIL.n126 VTAIL.n81 171.744
R240 VTAIL.n133 VTAIL.n81 171.744
R241 VTAIL.n134 VTAIL.n133 171.744
R242 VTAIL.n134 VTAIL.n77 171.744
R243 VTAIL.n141 VTAIL.n77 171.744
R244 VTAIL.n142 VTAIL.n141 171.744
R245 VTAIL.n174 VTAIL.n173 171.744
R246 VTAIL.n174 VTAIL.n167 171.744
R247 VTAIL.n181 VTAIL.n167 171.744
R248 VTAIL.n182 VTAIL.n181 171.744
R249 VTAIL.n182 VTAIL.n163 171.744
R250 VTAIL.n190 VTAIL.n163 171.744
R251 VTAIL.n191 VTAIL.n190 171.744
R252 VTAIL.n192 VTAIL.n191 171.744
R253 VTAIL.n192 VTAIL.n159 171.744
R254 VTAIL.n199 VTAIL.n159 171.744
R255 VTAIL.n200 VTAIL.n199 171.744
R256 VTAIL.n200 VTAIL.n155 171.744
R257 VTAIL.n207 VTAIL.n155 171.744
R258 VTAIL.n208 VTAIL.n207 171.744
R259 VTAIL.n208 VTAIL.n151 171.744
R260 VTAIL.n215 VTAIL.n151 171.744
R261 VTAIL.n216 VTAIL.n215 171.744
R262 VTAIL.n512 VTAIL.n511 171.744
R263 VTAIL.n511 VTAIL.n447 171.744
R264 VTAIL.n504 VTAIL.n447 171.744
R265 VTAIL.n504 VTAIL.n503 171.744
R266 VTAIL.n503 VTAIL.n451 171.744
R267 VTAIL.n496 VTAIL.n451 171.744
R268 VTAIL.n496 VTAIL.n495 171.744
R269 VTAIL.n495 VTAIL.n455 171.744
R270 VTAIL.n460 VTAIL.n455 171.744
R271 VTAIL.n488 VTAIL.n460 171.744
R272 VTAIL.n488 VTAIL.n487 171.744
R273 VTAIL.n487 VTAIL.n461 171.744
R274 VTAIL.n480 VTAIL.n461 171.744
R275 VTAIL.n480 VTAIL.n479 171.744
R276 VTAIL.n479 VTAIL.n465 171.744
R277 VTAIL.n472 VTAIL.n465 171.744
R278 VTAIL.n472 VTAIL.n471 171.744
R279 VTAIL.n438 VTAIL.n437 171.744
R280 VTAIL.n437 VTAIL.n373 171.744
R281 VTAIL.n430 VTAIL.n373 171.744
R282 VTAIL.n430 VTAIL.n429 171.744
R283 VTAIL.n429 VTAIL.n377 171.744
R284 VTAIL.n422 VTAIL.n377 171.744
R285 VTAIL.n422 VTAIL.n421 171.744
R286 VTAIL.n421 VTAIL.n381 171.744
R287 VTAIL.n386 VTAIL.n381 171.744
R288 VTAIL.n414 VTAIL.n386 171.744
R289 VTAIL.n414 VTAIL.n413 171.744
R290 VTAIL.n413 VTAIL.n387 171.744
R291 VTAIL.n406 VTAIL.n387 171.744
R292 VTAIL.n406 VTAIL.n405 171.744
R293 VTAIL.n405 VTAIL.n391 171.744
R294 VTAIL.n398 VTAIL.n391 171.744
R295 VTAIL.n398 VTAIL.n397 171.744
R296 VTAIL.n364 VTAIL.n363 171.744
R297 VTAIL.n363 VTAIL.n299 171.744
R298 VTAIL.n356 VTAIL.n299 171.744
R299 VTAIL.n356 VTAIL.n355 171.744
R300 VTAIL.n355 VTAIL.n303 171.744
R301 VTAIL.n348 VTAIL.n303 171.744
R302 VTAIL.n348 VTAIL.n347 171.744
R303 VTAIL.n347 VTAIL.n307 171.744
R304 VTAIL.n312 VTAIL.n307 171.744
R305 VTAIL.n340 VTAIL.n312 171.744
R306 VTAIL.n340 VTAIL.n339 171.744
R307 VTAIL.n339 VTAIL.n313 171.744
R308 VTAIL.n332 VTAIL.n313 171.744
R309 VTAIL.n332 VTAIL.n331 171.744
R310 VTAIL.n331 VTAIL.n317 171.744
R311 VTAIL.n324 VTAIL.n317 171.744
R312 VTAIL.n324 VTAIL.n323 171.744
R313 VTAIL.n290 VTAIL.n289 171.744
R314 VTAIL.n289 VTAIL.n225 171.744
R315 VTAIL.n282 VTAIL.n225 171.744
R316 VTAIL.n282 VTAIL.n281 171.744
R317 VTAIL.n281 VTAIL.n229 171.744
R318 VTAIL.n274 VTAIL.n229 171.744
R319 VTAIL.n274 VTAIL.n273 171.744
R320 VTAIL.n273 VTAIL.n233 171.744
R321 VTAIL.n238 VTAIL.n233 171.744
R322 VTAIL.n266 VTAIL.n238 171.744
R323 VTAIL.n266 VTAIL.n265 171.744
R324 VTAIL.n265 VTAIL.n239 171.744
R325 VTAIL.n258 VTAIL.n239 171.744
R326 VTAIL.n258 VTAIL.n257 171.744
R327 VTAIL.n257 VTAIL.n243 171.744
R328 VTAIL.n250 VTAIL.n243 171.744
R329 VTAIL.n250 VTAIL.n249 171.744
R330 VTAIL.n543 VTAIL.t1 85.8723
R331 VTAIL.n25 VTAIL.t2 85.8723
R332 VTAIL.n99 VTAIL.t6 85.8723
R333 VTAIL.n173 VTAIL.t7 85.8723
R334 VTAIL.n471 VTAIL.t4 85.8723
R335 VTAIL.n397 VTAIL.t5 85.8723
R336 VTAIL.n323 VTAIL.t0 85.8723
R337 VTAIL.n249 VTAIL.t3 85.8723
R338 VTAIL.n591 VTAIL.n590 30.052
R339 VTAIL.n73 VTAIL.n72 30.052
R340 VTAIL.n147 VTAIL.n146 30.052
R341 VTAIL.n221 VTAIL.n220 30.052
R342 VTAIL.n517 VTAIL.n516 30.052
R343 VTAIL.n443 VTAIL.n442 30.052
R344 VTAIL.n369 VTAIL.n368 30.052
R345 VTAIL.n295 VTAIL.n294 30.052
R346 VTAIL.n591 VTAIL.n517 27.66
R347 VTAIL.n295 VTAIL.n221 27.66
R348 VTAIL.n563 VTAIL.n530 13.1884
R349 VTAIL.n45 VTAIL.n12 13.1884
R350 VTAIL.n119 VTAIL.n86 13.1884
R351 VTAIL.n193 VTAIL.n160 13.1884
R352 VTAIL.n458 VTAIL.n456 13.1884
R353 VTAIL.n384 VTAIL.n382 13.1884
R354 VTAIL.n310 VTAIL.n308 13.1884
R355 VTAIL.n236 VTAIL.n234 13.1884
R356 VTAIL.n564 VTAIL.n532 12.8005
R357 VTAIL.n568 VTAIL.n567 12.8005
R358 VTAIL.n46 VTAIL.n14 12.8005
R359 VTAIL.n50 VTAIL.n49 12.8005
R360 VTAIL.n120 VTAIL.n88 12.8005
R361 VTAIL.n124 VTAIL.n123 12.8005
R362 VTAIL.n194 VTAIL.n162 12.8005
R363 VTAIL.n198 VTAIL.n197 12.8005
R364 VTAIL.n494 VTAIL.n493 12.8005
R365 VTAIL.n490 VTAIL.n489 12.8005
R366 VTAIL.n420 VTAIL.n419 12.8005
R367 VTAIL.n416 VTAIL.n415 12.8005
R368 VTAIL.n346 VTAIL.n345 12.8005
R369 VTAIL.n342 VTAIL.n341 12.8005
R370 VTAIL.n272 VTAIL.n271 12.8005
R371 VTAIL.n268 VTAIL.n267 12.8005
R372 VTAIL.n559 VTAIL.n558 12.0247
R373 VTAIL.n571 VTAIL.n528 12.0247
R374 VTAIL.n41 VTAIL.n40 12.0247
R375 VTAIL.n53 VTAIL.n10 12.0247
R376 VTAIL.n115 VTAIL.n114 12.0247
R377 VTAIL.n127 VTAIL.n84 12.0247
R378 VTAIL.n189 VTAIL.n188 12.0247
R379 VTAIL.n201 VTAIL.n158 12.0247
R380 VTAIL.n497 VTAIL.n454 12.0247
R381 VTAIL.n486 VTAIL.n459 12.0247
R382 VTAIL.n423 VTAIL.n380 12.0247
R383 VTAIL.n412 VTAIL.n385 12.0247
R384 VTAIL.n349 VTAIL.n306 12.0247
R385 VTAIL.n338 VTAIL.n311 12.0247
R386 VTAIL.n275 VTAIL.n232 12.0247
R387 VTAIL.n264 VTAIL.n237 12.0247
R388 VTAIL.n557 VTAIL.n534 11.249
R389 VTAIL.n572 VTAIL.n526 11.249
R390 VTAIL.n39 VTAIL.n16 11.249
R391 VTAIL.n54 VTAIL.n8 11.249
R392 VTAIL.n113 VTAIL.n90 11.249
R393 VTAIL.n128 VTAIL.n82 11.249
R394 VTAIL.n187 VTAIL.n164 11.249
R395 VTAIL.n202 VTAIL.n156 11.249
R396 VTAIL.n498 VTAIL.n452 11.249
R397 VTAIL.n485 VTAIL.n462 11.249
R398 VTAIL.n424 VTAIL.n378 11.249
R399 VTAIL.n411 VTAIL.n388 11.249
R400 VTAIL.n350 VTAIL.n304 11.249
R401 VTAIL.n337 VTAIL.n314 11.249
R402 VTAIL.n276 VTAIL.n230 11.249
R403 VTAIL.n263 VTAIL.n240 11.249
R404 VTAIL.n542 VTAIL.n541 10.7239
R405 VTAIL.n24 VTAIL.n23 10.7239
R406 VTAIL.n98 VTAIL.n97 10.7239
R407 VTAIL.n172 VTAIL.n171 10.7239
R408 VTAIL.n470 VTAIL.n469 10.7239
R409 VTAIL.n396 VTAIL.n395 10.7239
R410 VTAIL.n322 VTAIL.n321 10.7239
R411 VTAIL.n248 VTAIL.n247 10.7239
R412 VTAIL.n554 VTAIL.n553 10.4732
R413 VTAIL.n576 VTAIL.n575 10.4732
R414 VTAIL.n36 VTAIL.n35 10.4732
R415 VTAIL.n58 VTAIL.n57 10.4732
R416 VTAIL.n110 VTAIL.n109 10.4732
R417 VTAIL.n132 VTAIL.n131 10.4732
R418 VTAIL.n184 VTAIL.n183 10.4732
R419 VTAIL.n206 VTAIL.n205 10.4732
R420 VTAIL.n502 VTAIL.n501 10.4732
R421 VTAIL.n482 VTAIL.n481 10.4732
R422 VTAIL.n428 VTAIL.n427 10.4732
R423 VTAIL.n408 VTAIL.n407 10.4732
R424 VTAIL.n354 VTAIL.n353 10.4732
R425 VTAIL.n334 VTAIL.n333 10.4732
R426 VTAIL.n280 VTAIL.n279 10.4732
R427 VTAIL.n260 VTAIL.n259 10.4732
R428 VTAIL.n550 VTAIL.n536 9.69747
R429 VTAIL.n579 VTAIL.n524 9.69747
R430 VTAIL.n32 VTAIL.n18 9.69747
R431 VTAIL.n61 VTAIL.n6 9.69747
R432 VTAIL.n106 VTAIL.n92 9.69747
R433 VTAIL.n135 VTAIL.n80 9.69747
R434 VTAIL.n180 VTAIL.n166 9.69747
R435 VTAIL.n209 VTAIL.n154 9.69747
R436 VTAIL.n505 VTAIL.n450 9.69747
R437 VTAIL.n478 VTAIL.n464 9.69747
R438 VTAIL.n431 VTAIL.n376 9.69747
R439 VTAIL.n404 VTAIL.n390 9.69747
R440 VTAIL.n357 VTAIL.n302 9.69747
R441 VTAIL.n330 VTAIL.n316 9.69747
R442 VTAIL.n283 VTAIL.n228 9.69747
R443 VTAIL.n256 VTAIL.n242 9.69747
R444 VTAIL.n590 VTAIL.n589 9.45567
R445 VTAIL.n72 VTAIL.n71 9.45567
R446 VTAIL.n146 VTAIL.n145 9.45567
R447 VTAIL.n220 VTAIL.n219 9.45567
R448 VTAIL.n516 VTAIL.n515 9.45567
R449 VTAIL.n442 VTAIL.n441 9.45567
R450 VTAIL.n368 VTAIL.n367 9.45567
R451 VTAIL.n294 VTAIL.n293 9.45567
R452 VTAIL.n589 VTAIL.n588 9.3005
R453 VTAIL.n583 VTAIL.n582 9.3005
R454 VTAIL.n581 VTAIL.n580 9.3005
R455 VTAIL.n524 VTAIL.n523 9.3005
R456 VTAIL.n575 VTAIL.n574 9.3005
R457 VTAIL.n573 VTAIL.n572 9.3005
R458 VTAIL.n528 VTAIL.n527 9.3005
R459 VTAIL.n567 VTAIL.n566 9.3005
R460 VTAIL.n540 VTAIL.n539 9.3005
R461 VTAIL.n547 VTAIL.n546 9.3005
R462 VTAIL.n549 VTAIL.n548 9.3005
R463 VTAIL.n536 VTAIL.n535 9.3005
R464 VTAIL.n555 VTAIL.n554 9.3005
R465 VTAIL.n557 VTAIL.n556 9.3005
R466 VTAIL.n558 VTAIL.n531 9.3005
R467 VTAIL.n565 VTAIL.n564 9.3005
R468 VTAIL.n520 VTAIL.n519 9.3005
R469 VTAIL.n71 VTAIL.n70 9.3005
R470 VTAIL.n65 VTAIL.n64 9.3005
R471 VTAIL.n63 VTAIL.n62 9.3005
R472 VTAIL.n6 VTAIL.n5 9.3005
R473 VTAIL.n57 VTAIL.n56 9.3005
R474 VTAIL.n55 VTAIL.n54 9.3005
R475 VTAIL.n10 VTAIL.n9 9.3005
R476 VTAIL.n49 VTAIL.n48 9.3005
R477 VTAIL.n22 VTAIL.n21 9.3005
R478 VTAIL.n29 VTAIL.n28 9.3005
R479 VTAIL.n31 VTAIL.n30 9.3005
R480 VTAIL.n18 VTAIL.n17 9.3005
R481 VTAIL.n37 VTAIL.n36 9.3005
R482 VTAIL.n39 VTAIL.n38 9.3005
R483 VTAIL.n40 VTAIL.n13 9.3005
R484 VTAIL.n47 VTAIL.n46 9.3005
R485 VTAIL.n2 VTAIL.n1 9.3005
R486 VTAIL.n145 VTAIL.n144 9.3005
R487 VTAIL.n139 VTAIL.n138 9.3005
R488 VTAIL.n137 VTAIL.n136 9.3005
R489 VTAIL.n80 VTAIL.n79 9.3005
R490 VTAIL.n131 VTAIL.n130 9.3005
R491 VTAIL.n129 VTAIL.n128 9.3005
R492 VTAIL.n84 VTAIL.n83 9.3005
R493 VTAIL.n123 VTAIL.n122 9.3005
R494 VTAIL.n96 VTAIL.n95 9.3005
R495 VTAIL.n103 VTAIL.n102 9.3005
R496 VTAIL.n105 VTAIL.n104 9.3005
R497 VTAIL.n92 VTAIL.n91 9.3005
R498 VTAIL.n111 VTAIL.n110 9.3005
R499 VTAIL.n113 VTAIL.n112 9.3005
R500 VTAIL.n114 VTAIL.n87 9.3005
R501 VTAIL.n121 VTAIL.n120 9.3005
R502 VTAIL.n76 VTAIL.n75 9.3005
R503 VTAIL.n219 VTAIL.n218 9.3005
R504 VTAIL.n213 VTAIL.n212 9.3005
R505 VTAIL.n211 VTAIL.n210 9.3005
R506 VTAIL.n154 VTAIL.n153 9.3005
R507 VTAIL.n205 VTAIL.n204 9.3005
R508 VTAIL.n203 VTAIL.n202 9.3005
R509 VTAIL.n158 VTAIL.n157 9.3005
R510 VTAIL.n197 VTAIL.n196 9.3005
R511 VTAIL.n170 VTAIL.n169 9.3005
R512 VTAIL.n177 VTAIL.n176 9.3005
R513 VTAIL.n179 VTAIL.n178 9.3005
R514 VTAIL.n166 VTAIL.n165 9.3005
R515 VTAIL.n185 VTAIL.n184 9.3005
R516 VTAIL.n187 VTAIL.n186 9.3005
R517 VTAIL.n188 VTAIL.n161 9.3005
R518 VTAIL.n195 VTAIL.n194 9.3005
R519 VTAIL.n150 VTAIL.n149 9.3005
R520 VTAIL.n468 VTAIL.n467 9.3005
R521 VTAIL.n475 VTAIL.n474 9.3005
R522 VTAIL.n477 VTAIL.n476 9.3005
R523 VTAIL.n464 VTAIL.n463 9.3005
R524 VTAIL.n483 VTAIL.n482 9.3005
R525 VTAIL.n485 VTAIL.n484 9.3005
R526 VTAIL.n459 VTAIL.n457 9.3005
R527 VTAIL.n491 VTAIL.n490 9.3005
R528 VTAIL.n515 VTAIL.n514 9.3005
R529 VTAIL.n446 VTAIL.n445 9.3005
R530 VTAIL.n509 VTAIL.n508 9.3005
R531 VTAIL.n507 VTAIL.n506 9.3005
R532 VTAIL.n450 VTAIL.n449 9.3005
R533 VTAIL.n501 VTAIL.n500 9.3005
R534 VTAIL.n499 VTAIL.n498 9.3005
R535 VTAIL.n454 VTAIL.n453 9.3005
R536 VTAIL.n493 VTAIL.n492 9.3005
R537 VTAIL.n394 VTAIL.n393 9.3005
R538 VTAIL.n401 VTAIL.n400 9.3005
R539 VTAIL.n403 VTAIL.n402 9.3005
R540 VTAIL.n390 VTAIL.n389 9.3005
R541 VTAIL.n409 VTAIL.n408 9.3005
R542 VTAIL.n411 VTAIL.n410 9.3005
R543 VTAIL.n385 VTAIL.n383 9.3005
R544 VTAIL.n417 VTAIL.n416 9.3005
R545 VTAIL.n441 VTAIL.n440 9.3005
R546 VTAIL.n372 VTAIL.n371 9.3005
R547 VTAIL.n435 VTAIL.n434 9.3005
R548 VTAIL.n433 VTAIL.n432 9.3005
R549 VTAIL.n376 VTAIL.n375 9.3005
R550 VTAIL.n427 VTAIL.n426 9.3005
R551 VTAIL.n425 VTAIL.n424 9.3005
R552 VTAIL.n380 VTAIL.n379 9.3005
R553 VTAIL.n419 VTAIL.n418 9.3005
R554 VTAIL.n320 VTAIL.n319 9.3005
R555 VTAIL.n327 VTAIL.n326 9.3005
R556 VTAIL.n329 VTAIL.n328 9.3005
R557 VTAIL.n316 VTAIL.n315 9.3005
R558 VTAIL.n335 VTAIL.n334 9.3005
R559 VTAIL.n337 VTAIL.n336 9.3005
R560 VTAIL.n311 VTAIL.n309 9.3005
R561 VTAIL.n343 VTAIL.n342 9.3005
R562 VTAIL.n367 VTAIL.n366 9.3005
R563 VTAIL.n298 VTAIL.n297 9.3005
R564 VTAIL.n361 VTAIL.n360 9.3005
R565 VTAIL.n359 VTAIL.n358 9.3005
R566 VTAIL.n302 VTAIL.n301 9.3005
R567 VTAIL.n353 VTAIL.n352 9.3005
R568 VTAIL.n351 VTAIL.n350 9.3005
R569 VTAIL.n306 VTAIL.n305 9.3005
R570 VTAIL.n345 VTAIL.n344 9.3005
R571 VTAIL.n246 VTAIL.n245 9.3005
R572 VTAIL.n253 VTAIL.n252 9.3005
R573 VTAIL.n255 VTAIL.n254 9.3005
R574 VTAIL.n242 VTAIL.n241 9.3005
R575 VTAIL.n261 VTAIL.n260 9.3005
R576 VTAIL.n263 VTAIL.n262 9.3005
R577 VTAIL.n237 VTAIL.n235 9.3005
R578 VTAIL.n269 VTAIL.n268 9.3005
R579 VTAIL.n293 VTAIL.n292 9.3005
R580 VTAIL.n224 VTAIL.n223 9.3005
R581 VTAIL.n287 VTAIL.n286 9.3005
R582 VTAIL.n285 VTAIL.n284 9.3005
R583 VTAIL.n228 VTAIL.n227 9.3005
R584 VTAIL.n279 VTAIL.n278 9.3005
R585 VTAIL.n277 VTAIL.n276 9.3005
R586 VTAIL.n232 VTAIL.n231 9.3005
R587 VTAIL.n271 VTAIL.n270 9.3005
R588 VTAIL.n549 VTAIL.n538 8.92171
R589 VTAIL.n580 VTAIL.n522 8.92171
R590 VTAIL.n31 VTAIL.n20 8.92171
R591 VTAIL.n62 VTAIL.n4 8.92171
R592 VTAIL.n105 VTAIL.n94 8.92171
R593 VTAIL.n136 VTAIL.n78 8.92171
R594 VTAIL.n179 VTAIL.n168 8.92171
R595 VTAIL.n210 VTAIL.n152 8.92171
R596 VTAIL.n506 VTAIL.n448 8.92171
R597 VTAIL.n477 VTAIL.n466 8.92171
R598 VTAIL.n432 VTAIL.n374 8.92171
R599 VTAIL.n403 VTAIL.n392 8.92171
R600 VTAIL.n358 VTAIL.n300 8.92171
R601 VTAIL.n329 VTAIL.n318 8.92171
R602 VTAIL.n284 VTAIL.n226 8.92171
R603 VTAIL.n255 VTAIL.n244 8.92171
R604 VTAIL.n546 VTAIL.n545 8.14595
R605 VTAIL.n584 VTAIL.n583 8.14595
R606 VTAIL.n28 VTAIL.n27 8.14595
R607 VTAIL.n66 VTAIL.n65 8.14595
R608 VTAIL.n102 VTAIL.n101 8.14595
R609 VTAIL.n140 VTAIL.n139 8.14595
R610 VTAIL.n176 VTAIL.n175 8.14595
R611 VTAIL.n214 VTAIL.n213 8.14595
R612 VTAIL.n510 VTAIL.n509 8.14595
R613 VTAIL.n474 VTAIL.n473 8.14595
R614 VTAIL.n436 VTAIL.n435 8.14595
R615 VTAIL.n400 VTAIL.n399 8.14595
R616 VTAIL.n362 VTAIL.n361 8.14595
R617 VTAIL.n326 VTAIL.n325 8.14595
R618 VTAIL.n288 VTAIL.n287 8.14595
R619 VTAIL.n252 VTAIL.n251 8.14595
R620 VTAIL.n542 VTAIL.n540 7.3702
R621 VTAIL.n587 VTAIL.n520 7.3702
R622 VTAIL.n590 VTAIL.n518 7.3702
R623 VTAIL.n24 VTAIL.n22 7.3702
R624 VTAIL.n69 VTAIL.n2 7.3702
R625 VTAIL.n72 VTAIL.n0 7.3702
R626 VTAIL.n98 VTAIL.n96 7.3702
R627 VTAIL.n143 VTAIL.n76 7.3702
R628 VTAIL.n146 VTAIL.n74 7.3702
R629 VTAIL.n172 VTAIL.n170 7.3702
R630 VTAIL.n217 VTAIL.n150 7.3702
R631 VTAIL.n220 VTAIL.n148 7.3702
R632 VTAIL.n516 VTAIL.n444 7.3702
R633 VTAIL.n513 VTAIL.n446 7.3702
R634 VTAIL.n470 VTAIL.n468 7.3702
R635 VTAIL.n442 VTAIL.n370 7.3702
R636 VTAIL.n439 VTAIL.n372 7.3702
R637 VTAIL.n396 VTAIL.n394 7.3702
R638 VTAIL.n368 VTAIL.n296 7.3702
R639 VTAIL.n365 VTAIL.n298 7.3702
R640 VTAIL.n322 VTAIL.n320 7.3702
R641 VTAIL.n294 VTAIL.n222 7.3702
R642 VTAIL.n291 VTAIL.n224 7.3702
R643 VTAIL.n248 VTAIL.n246 7.3702
R644 VTAIL.n588 VTAIL.n587 6.59444
R645 VTAIL.n588 VTAIL.n518 6.59444
R646 VTAIL.n70 VTAIL.n69 6.59444
R647 VTAIL.n70 VTAIL.n0 6.59444
R648 VTAIL.n144 VTAIL.n143 6.59444
R649 VTAIL.n144 VTAIL.n74 6.59444
R650 VTAIL.n218 VTAIL.n217 6.59444
R651 VTAIL.n218 VTAIL.n148 6.59444
R652 VTAIL.n514 VTAIL.n444 6.59444
R653 VTAIL.n514 VTAIL.n513 6.59444
R654 VTAIL.n440 VTAIL.n370 6.59444
R655 VTAIL.n440 VTAIL.n439 6.59444
R656 VTAIL.n366 VTAIL.n296 6.59444
R657 VTAIL.n366 VTAIL.n365 6.59444
R658 VTAIL.n292 VTAIL.n222 6.59444
R659 VTAIL.n292 VTAIL.n291 6.59444
R660 VTAIL.n545 VTAIL.n540 5.81868
R661 VTAIL.n584 VTAIL.n520 5.81868
R662 VTAIL.n27 VTAIL.n22 5.81868
R663 VTAIL.n66 VTAIL.n2 5.81868
R664 VTAIL.n101 VTAIL.n96 5.81868
R665 VTAIL.n140 VTAIL.n76 5.81868
R666 VTAIL.n175 VTAIL.n170 5.81868
R667 VTAIL.n214 VTAIL.n150 5.81868
R668 VTAIL.n510 VTAIL.n446 5.81868
R669 VTAIL.n473 VTAIL.n468 5.81868
R670 VTAIL.n436 VTAIL.n372 5.81868
R671 VTAIL.n399 VTAIL.n394 5.81868
R672 VTAIL.n362 VTAIL.n298 5.81868
R673 VTAIL.n325 VTAIL.n320 5.81868
R674 VTAIL.n288 VTAIL.n224 5.81868
R675 VTAIL.n251 VTAIL.n246 5.81868
R676 VTAIL.n546 VTAIL.n538 5.04292
R677 VTAIL.n583 VTAIL.n522 5.04292
R678 VTAIL.n28 VTAIL.n20 5.04292
R679 VTAIL.n65 VTAIL.n4 5.04292
R680 VTAIL.n102 VTAIL.n94 5.04292
R681 VTAIL.n139 VTAIL.n78 5.04292
R682 VTAIL.n176 VTAIL.n168 5.04292
R683 VTAIL.n213 VTAIL.n152 5.04292
R684 VTAIL.n509 VTAIL.n448 5.04292
R685 VTAIL.n474 VTAIL.n466 5.04292
R686 VTAIL.n435 VTAIL.n374 5.04292
R687 VTAIL.n400 VTAIL.n392 5.04292
R688 VTAIL.n361 VTAIL.n300 5.04292
R689 VTAIL.n326 VTAIL.n318 5.04292
R690 VTAIL.n287 VTAIL.n226 5.04292
R691 VTAIL.n252 VTAIL.n244 5.04292
R692 VTAIL.n550 VTAIL.n549 4.26717
R693 VTAIL.n580 VTAIL.n579 4.26717
R694 VTAIL.n32 VTAIL.n31 4.26717
R695 VTAIL.n62 VTAIL.n61 4.26717
R696 VTAIL.n106 VTAIL.n105 4.26717
R697 VTAIL.n136 VTAIL.n135 4.26717
R698 VTAIL.n180 VTAIL.n179 4.26717
R699 VTAIL.n210 VTAIL.n209 4.26717
R700 VTAIL.n506 VTAIL.n505 4.26717
R701 VTAIL.n478 VTAIL.n477 4.26717
R702 VTAIL.n432 VTAIL.n431 4.26717
R703 VTAIL.n404 VTAIL.n403 4.26717
R704 VTAIL.n358 VTAIL.n357 4.26717
R705 VTAIL.n330 VTAIL.n329 4.26717
R706 VTAIL.n284 VTAIL.n283 4.26717
R707 VTAIL.n256 VTAIL.n255 4.26717
R708 VTAIL.n369 VTAIL.n295 3.69878
R709 VTAIL.n517 VTAIL.n443 3.69878
R710 VTAIL.n221 VTAIL.n147 3.69878
R711 VTAIL.n553 VTAIL.n536 3.49141
R712 VTAIL.n576 VTAIL.n524 3.49141
R713 VTAIL.n35 VTAIL.n18 3.49141
R714 VTAIL.n58 VTAIL.n6 3.49141
R715 VTAIL.n109 VTAIL.n92 3.49141
R716 VTAIL.n132 VTAIL.n80 3.49141
R717 VTAIL.n183 VTAIL.n166 3.49141
R718 VTAIL.n206 VTAIL.n154 3.49141
R719 VTAIL.n502 VTAIL.n450 3.49141
R720 VTAIL.n481 VTAIL.n464 3.49141
R721 VTAIL.n428 VTAIL.n376 3.49141
R722 VTAIL.n407 VTAIL.n390 3.49141
R723 VTAIL.n354 VTAIL.n302 3.49141
R724 VTAIL.n333 VTAIL.n316 3.49141
R725 VTAIL.n280 VTAIL.n228 3.49141
R726 VTAIL.n259 VTAIL.n242 3.49141
R727 VTAIL.n554 VTAIL.n534 2.71565
R728 VTAIL.n575 VTAIL.n526 2.71565
R729 VTAIL.n36 VTAIL.n16 2.71565
R730 VTAIL.n57 VTAIL.n8 2.71565
R731 VTAIL.n110 VTAIL.n90 2.71565
R732 VTAIL.n131 VTAIL.n82 2.71565
R733 VTAIL.n184 VTAIL.n164 2.71565
R734 VTAIL.n205 VTAIL.n156 2.71565
R735 VTAIL.n501 VTAIL.n452 2.71565
R736 VTAIL.n482 VTAIL.n462 2.71565
R737 VTAIL.n427 VTAIL.n378 2.71565
R738 VTAIL.n408 VTAIL.n388 2.71565
R739 VTAIL.n353 VTAIL.n304 2.71565
R740 VTAIL.n334 VTAIL.n314 2.71565
R741 VTAIL.n279 VTAIL.n230 2.71565
R742 VTAIL.n260 VTAIL.n240 2.71565
R743 VTAIL.n541 VTAIL.n539 2.41282
R744 VTAIL.n23 VTAIL.n21 2.41282
R745 VTAIL.n97 VTAIL.n95 2.41282
R746 VTAIL.n171 VTAIL.n169 2.41282
R747 VTAIL.n469 VTAIL.n467 2.41282
R748 VTAIL.n395 VTAIL.n393 2.41282
R749 VTAIL.n321 VTAIL.n319 2.41282
R750 VTAIL.n247 VTAIL.n245 2.41282
R751 VTAIL.n559 VTAIL.n557 1.93989
R752 VTAIL.n572 VTAIL.n571 1.93989
R753 VTAIL.n41 VTAIL.n39 1.93989
R754 VTAIL.n54 VTAIL.n53 1.93989
R755 VTAIL.n115 VTAIL.n113 1.93989
R756 VTAIL.n128 VTAIL.n127 1.93989
R757 VTAIL.n189 VTAIL.n187 1.93989
R758 VTAIL.n202 VTAIL.n201 1.93989
R759 VTAIL.n498 VTAIL.n497 1.93989
R760 VTAIL.n486 VTAIL.n485 1.93989
R761 VTAIL.n424 VTAIL.n423 1.93989
R762 VTAIL.n412 VTAIL.n411 1.93989
R763 VTAIL.n350 VTAIL.n349 1.93989
R764 VTAIL.n338 VTAIL.n337 1.93989
R765 VTAIL.n276 VTAIL.n275 1.93989
R766 VTAIL.n264 VTAIL.n263 1.93989
R767 VTAIL VTAIL.n73 1.90783
R768 VTAIL VTAIL.n591 1.79145
R769 VTAIL.n558 VTAIL.n532 1.16414
R770 VTAIL.n568 VTAIL.n528 1.16414
R771 VTAIL.n40 VTAIL.n14 1.16414
R772 VTAIL.n50 VTAIL.n10 1.16414
R773 VTAIL.n114 VTAIL.n88 1.16414
R774 VTAIL.n124 VTAIL.n84 1.16414
R775 VTAIL.n188 VTAIL.n162 1.16414
R776 VTAIL.n198 VTAIL.n158 1.16414
R777 VTAIL.n494 VTAIL.n454 1.16414
R778 VTAIL.n489 VTAIL.n459 1.16414
R779 VTAIL.n420 VTAIL.n380 1.16414
R780 VTAIL.n415 VTAIL.n385 1.16414
R781 VTAIL.n346 VTAIL.n306 1.16414
R782 VTAIL.n341 VTAIL.n311 1.16414
R783 VTAIL.n272 VTAIL.n232 1.16414
R784 VTAIL.n267 VTAIL.n237 1.16414
R785 VTAIL.n443 VTAIL.n369 0.470328
R786 VTAIL.n147 VTAIL.n73 0.470328
R787 VTAIL.n564 VTAIL.n563 0.388379
R788 VTAIL.n567 VTAIL.n530 0.388379
R789 VTAIL.n46 VTAIL.n45 0.388379
R790 VTAIL.n49 VTAIL.n12 0.388379
R791 VTAIL.n120 VTAIL.n119 0.388379
R792 VTAIL.n123 VTAIL.n86 0.388379
R793 VTAIL.n194 VTAIL.n193 0.388379
R794 VTAIL.n197 VTAIL.n160 0.388379
R795 VTAIL.n493 VTAIL.n456 0.388379
R796 VTAIL.n490 VTAIL.n458 0.388379
R797 VTAIL.n419 VTAIL.n382 0.388379
R798 VTAIL.n416 VTAIL.n384 0.388379
R799 VTAIL.n345 VTAIL.n308 0.388379
R800 VTAIL.n342 VTAIL.n310 0.388379
R801 VTAIL.n271 VTAIL.n234 0.388379
R802 VTAIL.n268 VTAIL.n236 0.388379
R803 VTAIL.n547 VTAIL.n539 0.155672
R804 VTAIL.n548 VTAIL.n547 0.155672
R805 VTAIL.n548 VTAIL.n535 0.155672
R806 VTAIL.n555 VTAIL.n535 0.155672
R807 VTAIL.n556 VTAIL.n555 0.155672
R808 VTAIL.n556 VTAIL.n531 0.155672
R809 VTAIL.n565 VTAIL.n531 0.155672
R810 VTAIL.n566 VTAIL.n565 0.155672
R811 VTAIL.n566 VTAIL.n527 0.155672
R812 VTAIL.n573 VTAIL.n527 0.155672
R813 VTAIL.n574 VTAIL.n573 0.155672
R814 VTAIL.n574 VTAIL.n523 0.155672
R815 VTAIL.n581 VTAIL.n523 0.155672
R816 VTAIL.n582 VTAIL.n581 0.155672
R817 VTAIL.n582 VTAIL.n519 0.155672
R818 VTAIL.n589 VTAIL.n519 0.155672
R819 VTAIL.n29 VTAIL.n21 0.155672
R820 VTAIL.n30 VTAIL.n29 0.155672
R821 VTAIL.n30 VTAIL.n17 0.155672
R822 VTAIL.n37 VTAIL.n17 0.155672
R823 VTAIL.n38 VTAIL.n37 0.155672
R824 VTAIL.n38 VTAIL.n13 0.155672
R825 VTAIL.n47 VTAIL.n13 0.155672
R826 VTAIL.n48 VTAIL.n47 0.155672
R827 VTAIL.n48 VTAIL.n9 0.155672
R828 VTAIL.n55 VTAIL.n9 0.155672
R829 VTAIL.n56 VTAIL.n55 0.155672
R830 VTAIL.n56 VTAIL.n5 0.155672
R831 VTAIL.n63 VTAIL.n5 0.155672
R832 VTAIL.n64 VTAIL.n63 0.155672
R833 VTAIL.n64 VTAIL.n1 0.155672
R834 VTAIL.n71 VTAIL.n1 0.155672
R835 VTAIL.n103 VTAIL.n95 0.155672
R836 VTAIL.n104 VTAIL.n103 0.155672
R837 VTAIL.n104 VTAIL.n91 0.155672
R838 VTAIL.n111 VTAIL.n91 0.155672
R839 VTAIL.n112 VTAIL.n111 0.155672
R840 VTAIL.n112 VTAIL.n87 0.155672
R841 VTAIL.n121 VTAIL.n87 0.155672
R842 VTAIL.n122 VTAIL.n121 0.155672
R843 VTAIL.n122 VTAIL.n83 0.155672
R844 VTAIL.n129 VTAIL.n83 0.155672
R845 VTAIL.n130 VTAIL.n129 0.155672
R846 VTAIL.n130 VTAIL.n79 0.155672
R847 VTAIL.n137 VTAIL.n79 0.155672
R848 VTAIL.n138 VTAIL.n137 0.155672
R849 VTAIL.n138 VTAIL.n75 0.155672
R850 VTAIL.n145 VTAIL.n75 0.155672
R851 VTAIL.n177 VTAIL.n169 0.155672
R852 VTAIL.n178 VTAIL.n177 0.155672
R853 VTAIL.n178 VTAIL.n165 0.155672
R854 VTAIL.n185 VTAIL.n165 0.155672
R855 VTAIL.n186 VTAIL.n185 0.155672
R856 VTAIL.n186 VTAIL.n161 0.155672
R857 VTAIL.n195 VTAIL.n161 0.155672
R858 VTAIL.n196 VTAIL.n195 0.155672
R859 VTAIL.n196 VTAIL.n157 0.155672
R860 VTAIL.n203 VTAIL.n157 0.155672
R861 VTAIL.n204 VTAIL.n203 0.155672
R862 VTAIL.n204 VTAIL.n153 0.155672
R863 VTAIL.n211 VTAIL.n153 0.155672
R864 VTAIL.n212 VTAIL.n211 0.155672
R865 VTAIL.n212 VTAIL.n149 0.155672
R866 VTAIL.n219 VTAIL.n149 0.155672
R867 VTAIL.n515 VTAIL.n445 0.155672
R868 VTAIL.n508 VTAIL.n445 0.155672
R869 VTAIL.n508 VTAIL.n507 0.155672
R870 VTAIL.n507 VTAIL.n449 0.155672
R871 VTAIL.n500 VTAIL.n449 0.155672
R872 VTAIL.n500 VTAIL.n499 0.155672
R873 VTAIL.n499 VTAIL.n453 0.155672
R874 VTAIL.n492 VTAIL.n453 0.155672
R875 VTAIL.n492 VTAIL.n491 0.155672
R876 VTAIL.n491 VTAIL.n457 0.155672
R877 VTAIL.n484 VTAIL.n457 0.155672
R878 VTAIL.n484 VTAIL.n483 0.155672
R879 VTAIL.n483 VTAIL.n463 0.155672
R880 VTAIL.n476 VTAIL.n463 0.155672
R881 VTAIL.n476 VTAIL.n475 0.155672
R882 VTAIL.n475 VTAIL.n467 0.155672
R883 VTAIL.n441 VTAIL.n371 0.155672
R884 VTAIL.n434 VTAIL.n371 0.155672
R885 VTAIL.n434 VTAIL.n433 0.155672
R886 VTAIL.n433 VTAIL.n375 0.155672
R887 VTAIL.n426 VTAIL.n375 0.155672
R888 VTAIL.n426 VTAIL.n425 0.155672
R889 VTAIL.n425 VTAIL.n379 0.155672
R890 VTAIL.n418 VTAIL.n379 0.155672
R891 VTAIL.n418 VTAIL.n417 0.155672
R892 VTAIL.n417 VTAIL.n383 0.155672
R893 VTAIL.n410 VTAIL.n383 0.155672
R894 VTAIL.n410 VTAIL.n409 0.155672
R895 VTAIL.n409 VTAIL.n389 0.155672
R896 VTAIL.n402 VTAIL.n389 0.155672
R897 VTAIL.n402 VTAIL.n401 0.155672
R898 VTAIL.n401 VTAIL.n393 0.155672
R899 VTAIL.n367 VTAIL.n297 0.155672
R900 VTAIL.n360 VTAIL.n297 0.155672
R901 VTAIL.n360 VTAIL.n359 0.155672
R902 VTAIL.n359 VTAIL.n301 0.155672
R903 VTAIL.n352 VTAIL.n301 0.155672
R904 VTAIL.n352 VTAIL.n351 0.155672
R905 VTAIL.n351 VTAIL.n305 0.155672
R906 VTAIL.n344 VTAIL.n305 0.155672
R907 VTAIL.n344 VTAIL.n343 0.155672
R908 VTAIL.n343 VTAIL.n309 0.155672
R909 VTAIL.n336 VTAIL.n309 0.155672
R910 VTAIL.n336 VTAIL.n335 0.155672
R911 VTAIL.n335 VTAIL.n315 0.155672
R912 VTAIL.n328 VTAIL.n315 0.155672
R913 VTAIL.n328 VTAIL.n327 0.155672
R914 VTAIL.n327 VTAIL.n319 0.155672
R915 VTAIL.n293 VTAIL.n223 0.155672
R916 VTAIL.n286 VTAIL.n223 0.155672
R917 VTAIL.n286 VTAIL.n285 0.155672
R918 VTAIL.n285 VTAIL.n227 0.155672
R919 VTAIL.n278 VTAIL.n227 0.155672
R920 VTAIL.n278 VTAIL.n277 0.155672
R921 VTAIL.n277 VTAIL.n231 0.155672
R922 VTAIL.n270 VTAIL.n231 0.155672
R923 VTAIL.n270 VTAIL.n269 0.155672
R924 VTAIL.n269 VTAIL.n235 0.155672
R925 VTAIL.n262 VTAIL.n235 0.155672
R926 VTAIL.n262 VTAIL.n261 0.155672
R927 VTAIL.n261 VTAIL.n241 0.155672
R928 VTAIL.n254 VTAIL.n241 0.155672
R929 VTAIL.n254 VTAIL.n253 0.155672
R930 VTAIL.n253 VTAIL.n245 0.155672
R931 VDD1 VDD1.n1 117.076
R932 VDD1 VDD1.n0 70.2055
R933 VDD1.n0 VDD1.t1 2.41723
R934 VDD1.n0 VDD1.t2 2.41723
R935 VDD1.n1 VDD1.t0 2.41723
R936 VDD1.n1 VDD1.t3 2.41723
R937 B.n565 B.n564 585
R938 B.n566 B.n79 585
R939 B.n568 B.n567 585
R940 B.n569 B.n78 585
R941 B.n571 B.n570 585
R942 B.n572 B.n77 585
R943 B.n574 B.n573 585
R944 B.n575 B.n76 585
R945 B.n577 B.n576 585
R946 B.n578 B.n75 585
R947 B.n580 B.n579 585
R948 B.n581 B.n74 585
R949 B.n583 B.n582 585
R950 B.n584 B.n73 585
R951 B.n586 B.n585 585
R952 B.n587 B.n72 585
R953 B.n589 B.n588 585
R954 B.n590 B.n71 585
R955 B.n592 B.n591 585
R956 B.n593 B.n70 585
R957 B.n595 B.n594 585
R958 B.n596 B.n69 585
R959 B.n598 B.n597 585
R960 B.n599 B.n68 585
R961 B.n601 B.n600 585
R962 B.n602 B.n67 585
R963 B.n604 B.n603 585
R964 B.n605 B.n66 585
R965 B.n607 B.n606 585
R966 B.n608 B.n65 585
R967 B.n610 B.n609 585
R968 B.n611 B.n64 585
R969 B.n613 B.n612 585
R970 B.n614 B.n63 585
R971 B.n616 B.n615 585
R972 B.n617 B.n62 585
R973 B.n619 B.n618 585
R974 B.n620 B.n61 585
R975 B.n622 B.n621 585
R976 B.n623 B.n60 585
R977 B.n625 B.n624 585
R978 B.n626 B.n59 585
R979 B.n628 B.n627 585
R980 B.n629 B.n58 585
R981 B.n631 B.n630 585
R982 B.n632 B.n55 585
R983 B.n635 B.n634 585
R984 B.n636 B.n54 585
R985 B.n638 B.n637 585
R986 B.n639 B.n53 585
R987 B.n641 B.n640 585
R988 B.n642 B.n52 585
R989 B.n644 B.n643 585
R990 B.n645 B.n51 585
R991 B.n647 B.n646 585
R992 B.n649 B.n648 585
R993 B.n650 B.n47 585
R994 B.n652 B.n651 585
R995 B.n653 B.n46 585
R996 B.n655 B.n654 585
R997 B.n656 B.n45 585
R998 B.n658 B.n657 585
R999 B.n659 B.n44 585
R1000 B.n661 B.n660 585
R1001 B.n662 B.n43 585
R1002 B.n664 B.n663 585
R1003 B.n665 B.n42 585
R1004 B.n667 B.n666 585
R1005 B.n668 B.n41 585
R1006 B.n670 B.n669 585
R1007 B.n671 B.n40 585
R1008 B.n673 B.n672 585
R1009 B.n674 B.n39 585
R1010 B.n676 B.n675 585
R1011 B.n677 B.n38 585
R1012 B.n679 B.n678 585
R1013 B.n680 B.n37 585
R1014 B.n682 B.n681 585
R1015 B.n683 B.n36 585
R1016 B.n685 B.n684 585
R1017 B.n686 B.n35 585
R1018 B.n688 B.n687 585
R1019 B.n689 B.n34 585
R1020 B.n691 B.n690 585
R1021 B.n692 B.n33 585
R1022 B.n694 B.n693 585
R1023 B.n695 B.n32 585
R1024 B.n697 B.n696 585
R1025 B.n698 B.n31 585
R1026 B.n700 B.n699 585
R1027 B.n701 B.n30 585
R1028 B.n703 B.n702 585
R1029 B.n704 B.n29 585
R1030 B.n706 B.n705 585
R1031 B.n707 B.n28 585
R1032 B.n709 B.n708 585
R1033 B.n710 B.n27 585
R1034 B.n712 B.n711 585
R1035 B.n713 B.n26 585
R1036 B.n715 B.n714 585
R1037 B.n716 B.n25 585
R1038 B.n563 B.n80 585
R1039 B.n562 B.n561 585
R1040 B.n560 B.n81 585
R1041 B.n559 B.n558 585
R1042 B.n557 B.n82 585
R1043 B.n556 B.n555 585
R1044 B.n554 B.n83 585
R1045 B.n553 B.n552 585
R1046 B.n551 B.n84 585
R1047 B.n550 B.n549 585
R1048 B.n548 B.n85 585
R1049 B.n547 B.n546 585
R1050 B.n545 B.n86 585
R1051 B.n544 B.n543 585
R1052 B.n542 B.n87 585
R1053 B.n541 B.n540 585
R1054 B.n539 B.n88 585
R1055 B.n538 B.n537 585
R1056 B.n536 B.n89 585
R1057 B.n535 B.n534 585
R1058 B.n533 B.n90 585
R1059 B.n532 B.n531 585
R1060 B.n530 B.n91 585
R1061 B.n529 B.n528 585
R1062 B.n527 B.n92 585
R1063 B.n526 B.n525 585
R1064 B.n524 B.n93 585
R1065 B.n523 B.n522 585
R1066 B.n521 B.n94 585
R1067 B.n520 B.n519 585
R1068 B.n518 B.n95 585
R1069 B.n517 B.n516 585
R1070 B.n515 B.n96 585
R1071 B.n514 B.n513 585
R1072 B.n512 B.n97 585
R1073 B.n511 B.n510 585
R1074 B.n509 B.n98 585
R1075 B.n508 B.n507 585
R1076 B.n506 B.n99 585
R1077 B.n505 B.n504 585
R1078 B.n503 B.n100 585
R1079 B.n502 B.n501 585
R1080 B.n500 B.n101 585
R1081 B.n499 B.n498 585
R1082 B.n497 B.n102 585
R1083 B.n496 B.n495 585
R1084 B.n494 B.n103 585
R1085 B.n493 B.n492 585
R1086 B.n491 B.n104 585
R1087 B.n490 B.n489 585
R1088 B.n488 B.n105 585
R1089 B.n487 B.n486 585
R1090 B.n485 B.n106 585
R1091 B.n484 B.n483 585
R1092 B.n482 B.n107 585
R1093 B.n481 B.n480 585
R1094 B.n479 B.n108 585
R1095 B.n478 B.n477 585
R1096 B.n476 B.n109 585
R1097 B.n475 B.n474 585
R1098 B.n473 B.n110 585
R1099 B.n472 B.n471 585
R1100 B.n470 B.n111 585
R1101 B.n469 B.n468 585
R1102 B.n467 B.n112 585
R1103 B.n466 B.n465 585
R1104 B.n464 B.n113 585
R1105 B.n463 B.n462 585
R1106 B.n461 B.n114 585
R1107 B.n460 B.n459 585
R1108 B.n458 B.n115 585
R1109 B.n457 B.n456 585
R1110 B.n455 B.n116 585
R1111 B.n454 B.n453 585
R1112 B.n452 B.n117 585
R1113 B.n451 B.n450 585
R1114 B.n449 B.n118 585
R1115 B.n448 B.n447 585
R1116 B.n446 B.n119 585
R1117 B.n445 B.n444 585
R1118 B.n443 B.n120 585
R1119 B.n442 B.n441 585
R1120 B.n440 B.n121 585
R1121 B.n439 B.n438 585
R1122 B.n437 B.n122 585
R1123 B.n436 B.n435 585
R1124 B.n434 B.n123 585
R1125 B.n433 B.n432 585
R1126 B.n431 B.n124 585
R1127 B.n430 B.n429 585
R1128 B.n428 B.n125 585
R1129 B.n427 B.n426 585
R1130 B.n425 B.n126 585
R1131 B.n272 B.n181 585
R1132 B.n274 B.n273 585
R1133 B.n275 B.n180 585
R1134 B.n277 B.n276 585
R1135 B.n278 B.n179 585
R1136 B.n280 B.n279 585
R1137 B.n281 B.n178 585
R1138 B.n283 B.n282 585
R1139 B.n284 B.n177 585
R1140 B.n286 B.n285 585
R1141 B.n287 B.n176 585
R1142 B.n289 B.n288 585
R1143 B.n290 B.n175 585
R1144 B.n292 B.n291 585
R1145 B.n293 B.n174 585
R1146 B.n295 B.n294 585
R1147 B.n296 B.n173 585
R1148 B.n298 B.n297 585
R1149 B.n299 B.n172 585
R1150 B.n301 B.n300 585
R1151 B.n302 B.n171 585
R1152 B.n304 B.n303 585
R1153 B.n305 B.n170 585
R1154 B.n307 B.n306 585
R1155 B.n308 B.n169 585
R1156 B.n310 B.n309 585
R1157 B.n311 B.n168 585
R1158 B.n313 B.n312 585
R1159 B.n314 B.n167 585
R1160 B.n316 B.n315 585
R1161 B.n317 B.n166 585
R1162 B.n319 B.n318 585
R1163 B.n320 B.n165 585
R1164 B.n322 B.n321 585
R1165 B.n323 B.n164 585
R1166 B.n325 B.n324 585
R1167 B.n326 B.n163 585
R1168 B.n328 B.n327 585
R1169 B.n329 B.n162 585
R1170 B.n331 B.n330 585
R1171 B.n332 B.n161 585
R1172 B.n334 B.n333 585
R1173 B.n335 B.n160 585
R1174 B.n337 B.n336 585
R1175 B.n338 B.n159 585
R1176 B.n340 B.n339 585
R1177 B.n342 B.n341 585
R1178 B.n343 B.n155 585
R1179 B.n345 B.n344 585
R1180 B.n346 B.n154 585
R1181 B.n348 B.n347 585
R1182 B.n349 B.n153 585
R1183 B.n351 B.n350 585
R1184 B.n352 B.n152 585
R1185 B.n354 B.n353 585
R1186 B.n356 B.n149 585
R1187 B.n358 B.n357 585
R1188 B.n359 B.n148 585
R1189 B.n361 B.n360 585
R1190 B.n362 B.n147 585
R1191 B.n364 B.n363 585
R1192 B.n365 B.n146 585
R1193 B.n367 B.n366 585
R1194 B.n368 B.n145 585
R1195 B.n370 B.n369 585
R1196 B.n371 B.n144 585
R1197 B.n373 B.n372 585
R1198 B.n374 B.n143 585
R1199 B.n376 B.n375 585
R1200 B.n377 B.n142 585
R1201 B.n379 B.n378 585
R1202 B.n380 B.n141 585
R1203 B.n382 B.n381 585
R1204 B.n383 B.n140 585
R1205 B.n385 B.n384 585
R1206 B.n386 B.n139 585
R1207 B.n388 B.n387 585
R1208 B.n389 B.n138 585
R1209 B.n391 B.n390 585
R1210 B.n392 B.n137 585
R1211 B.n394 B.n393 585
R1212 B.n395 B.n136 585
R1213 B.n397 B.n396 585
R1214 B.n398 B.n135 585
R1215 B.n400 B.n399 585
R1216 B.n401 B.n134 585
R1217 B.n403 B.n402 585
R1218 B.n404 B.n133 585
R1219 B.n406 B.n405 585
R1220 B.n407 B.n132 585
R1221 B.n409 B.n408 585
R1222 B.n410 B.n131 585
R1223 B.n412 B.n411 585
R1224 B.n413 B.n130 585
R1225 B.n415 B.n414 585
R1226 B.n416 B.n129 585
R1227 B.n418 B.n417 585
R1228 B.n419 B.n128 585
R1229 B.n421 B.n420 585
R1230 B.n422 B.n127 585
R1231 B.n424 B.n423 585
R1232 B.n271 B.n270 585
R1233 B.n269 B.n182 585
R1234 B.n268 B.n267 585
R1235 B.n266 B.n183 585
R1236 B.n265 B.n264 585
R1237 B.n263 B.n184 585
R1238 B.n262 B.n261 585
R1239 B.n260 B.n185 585
R1240 B.n259 B.n258 585
R1241 B.n257 B.n186 585
R1242 B.n256 B.n255 585
R1243 B.n254 B.n187 585
R1244 B.n253 B.n252 585
R1245 B.n251 B.n188 585
R1246 B.n250 B.n249 585
R1247 B.n248 B.n189 585
R1248 B.n247 B.n246 585
R1249 B.n245 B.n190 585
R1250 B.n244 B.n243 585
R1251 B.n242 B.n191 585
R1252 B.n241 B.n240 585
R1253 B.n239 B.n192 585
R1254 B.n238 B.n237 585
R1255 B.n236 B.n193 585
R1256 B.n235 B.n234 585
R1257 B.n233 B.n194 585
R1258 B.n232 B.n231 585
R1259 B.n230 B.n195 585
R1260 B.n229 B.n228 585
R1261 B.n227 B.n196 585
R1262 B.n226 B.n225 585
R1263 B.n224 B.n197 585
R1264 B.n223 B.n222 585
R1265 B.n221 B.n198 585
R1266 B.n220 B.n219 585
R1267 B.n218 B.n199 585
R1268 B.n217 B.n216 585
R1269 B.n215 B.n200 585
R1270 B.n214 B.n213 585
R1271 B.n212 B.n201 585
R1272 B.n211 B.n210 585
R1273 B.n209 B.n202 585
R1274 B.n208 B.n207 585
R1275 B.n206 B.n203 585
R1276 B.n205 B.n204 585
R1277 B.n2 B.n0 585
R1278 B.n785 B.n1 585
R1279 B.n784 B.n783 585
R1280 B.n782 B.n3 585
R1281 B.n781 B.n780 585
R1282 B.n779 B.n4 585
R1283 B.n778 B.n777 585
R1284 B.n776 B.n5 585
R1285 B.n775 B.n774 585
R1286 B.n773 B.n6 585
R1287 B.n772 B.n771 585
R1288 B.n770 B.n7 585
R1289 B.n769 B.n768 585
R1290 B.n767 B.n8 585
R1291 B.n766 B.n765 585
R1292 B.n764 B.n9 585
R1293 B.n763 B.n762 585
R1294 B.n761 B.n10 585
R1295 B.n760 B.n759 585
R1296 B.n758 B.n11 585
R1297 B.n757 B.n756 585
R1298 B.n755 B.n12 585
R1299 B.n754 B.n753 585
R1300 B.n752 B.n13 585
R1301 B.n751 B.n750 585
R1302 B.n749 B.n14 585
R1303 B.n748 B.n747 585
R1304 B.n746 B.n15 585
R1305 B.n745 B.n744 585
R1306 B.n743 B.n16 585
R1307 B.n742 B.n741 585
R1308 B.n740 B.n17 585
R1309 B.n739 B.n738 585
R1310 B.n737 B.n18 585
R1311 B.n736 B.n735 585
R1312 B.n734 B.n19 585
R1313 B.n733 B.n732 585
R1314 B.n731 B.n20 585
R1315 B.n730 B.n729 585
R1316 B.n728 B.n21 585
R1317 B.n727 B.n726 585
R1318 B.n725 B.n22 585
R1319 B.n724 B.n723 585
R1320 B.n722 B.n23 585
R1321 B.n721 B.n720 585
R1322 B.n719 B.n24 585
R1323 B.n718 B.n717 585
R1324 B.n787 B.n786 585
R1325 B.n270 B.n181 521.33
R1326 B.n718 B.n25 521.33
R1327 B.n425 B.n424 521.33
R1328 B.n564 B.n563 521.33
R1329 B.n150 B.t11 484.969
R1330 B.n56 B.t4 484.969
R1331 B.n156 B.t2 484.969
R1332 B.n48 B.t7 484.969
R1333 B.n151 B.t10 401.769
R1334 B.n57 B.t5 401.769
R1335 B.n157 B.t1 401.769
R1336 B.n49 B.t8 401.769
R1337 B.n150 B.t9 291.318
R1338 B.n156 B.t0 291.318
R1339 B.n48 B.t6 291.318
R1340 B.n56 B.t3 291.318
R1341 B.n270 B.n269 163.367
R1342 B.n269 B.n268 163.367
R1343 B.n268 B.n183 163.367
R1344 B.n264 B.n183 163.367
R1345 B.n264 B.n263 163.367
R1346 B.n263 B.n262 163.367
R1347 B.n262 B.n185 163.367
R1348 B.n258 B.n185 163.367
R1349 B.n258 B.n257 163.367
R1350 B.n257 B.n256 163.367
R1351 B.n256 B.n187 163.367
R1352 B.n252 B.n187 163.367
R1353 B.n252 B.n251 163.367
R1354 B.n251 B.n250 163.367
R1355 B.n250 B.n189 163.367
R1356 B.n246 B.n189 163.367
R1357 B.n246 B.n245 163.367
R1358 B.n245 B.n244 163.367
R1359 B.n244 B.n191 163.367
R1360 B.n240 B.n191 163.367
R1361 B.n240 B.n239 163.367
R1362 B.n239 B.n238 163.367
R1363 B.n238 B.n193 163.367
R1364 B.n234 B.n193 163.367
R1365 B.n234 B.n233 163.367
R1366 B.n233 B.n232 163.367
R1367 B.n232 B.n195 163.367
R1368 B.n228 B.n195 163.367
R1369 B.n228 B.n227 163.367
R1370 B.n227 B.n226 163.367
R1371 B.n226 B.n197 163.367
R1372 B.n222 B.n197 163.367
R1373 B.n222 B.n221 163.367
R1374 B.n221 B.n220 163.367
R1375 B.n220 B.n199 163.367
R1376 B.n216 B.n199 163.367
R1377 B.n216 B.n215 163.367
R1378 B.n215 B.n214 163.367
R1379 B.n214 B.n201 163.367
R1380 B.n210 B.n201 163.367
R1381 B.n210 B.n209 163.367
R1382 B.n209 B.n208 163.367
R1383 B.n208 B.n203 163.367
R1384 B.n204 B.n203 163.367
R1385 B.n204 B.n2 163.367
R1386 B.n786 B.n2 163.367
R1387 B.n786 B.n785 163.367
R1388 B.n785 B.n784 163.367
R1389 B.n784 B.n3 163.367
R1390 B.n780 B.n3 163.367
R1391 B.n780 B.n779 163.367
R1392 B.n779 B.n778 163.367
R1393 B.n778 B.n5 163.367
R1394 B.n774 B.n5 163.367
R1395 B.n774 B.n773 163.367
R1396 B.n773 B.n772 163.367
R1397 B.n772 B.n7 163.367
R1398 B.n768 B.n7 163.367
R1399 B.n768 B.n767 163.367
R1400 B.n767 B.n766 163.367
R1401 B.n766 B.n9 163.367
R1402 B.n762 B.n9 163.367
R1403 B.n762 B.n761 163.367
R1404 B.n761 B.n760 163.367
R1405 B.n760 B.n11 163.367
R1406 B.n756 B.n11 163.367
R1407 B.n756 B.n755 163.367
R1408 B.n755 B.n754 163.367
R1409 B.n754 B.n13 163.367
R1410 B.n750 B.n13 163.367
R1411 B.n750 B.n749 163.367
R1412 B.n749 B.n748 163.367
R1413 B.n748 B.n15 163.367
R1414 B.n744 B.n15 163.367
R1415 B.n744 B.n743 163.367
R1416 B.n743 B.n742 163.367
R1417 B.n742 B.n17 163.367
R1418 B.n738 B.n17 163.367
R1419 B.n738 B.n737 163.367
R1420 B.n737 B.n736 163.367
R1421 B.n736 B.n19 163.367
R1422 B.n732 B.n19 163.367
R1423 B.n732 B.n731 163.367
R1424 B.n731 B.n730 163.367
R1425 B.n730 B.n21 163.367
R1426 B.n726 B.n21 163.367
R1427 B.n726 B.n725 163.367
R1428 B.n725 B.n724 163.367
R1429 B.n724 B.n23 163.367
R1430 B.n720 B.n23 163.367
R1431 B.n720 B.n719 163.367
R1432 B.n719 B.n718 163.367
R1433 B.n274 B.n181 163.367
R1434 B.n275 B.n274 163.367
R1435 B.n276 B.n275 163.367
R1436 B.n276 B.n179 163.367
R1437 B.n280 B.n179 163.367
R1438 B.n281 B.n280 163.367
R1439 B.n282 B.n281 163.367
R1440 B.n282 B.n177 163.367
R1441 B.n286 B.n177 163.367
R1442 B.n287 B.n286 163.367
R1443 B.n288 B.n287 163.367
R1444 B.n288 B.n175 163.367
R1445 B.n292 B.n175 163.367
R1446 B.n293 B.n292 163.367
R1447 B.n294 B.n293 163.367
R1448 B.n294 B.n173 163.367
R1449 B.n298 B.n173 163.367
R1450 B.n299 B.n298 163.367
R1451 B.n300 B.n299 163.367
R1452 B.n300 B.n171 163.367
R1453 B.n304 B.n171 163.367
R1454 B.n305 B.n304 163.367
R1455 B.n306 B.n305 163.367
R1456 B.n306 B.n169 163.367
R1457 B.n310 B.n169 163.367
R1458 B.n311 B.n310 163.367
R1459 B.n312 B.n311 163.367
R1460 B.n312 B.n167 163.367
R1461 B.n316 B.n167 163.367
R1462 B.n317 B.n316 163.367
R1463 B.n318 B.n317 163.367
R1464 B.n318 B.n165 163.367
R1465 B.n322 B.n165 163.367
R1466 B.n323 B.n322 163.367
R1467 B.n324 B.n323 163.367
R1468 B.n324 B.n163 163.367
R1469 B.n328 B.n163 163.367
R1470 B.n329 B.n328 163.367
R1471 B.n330 B.n329 163.367
R1472 B.n330 B.n161 163.367
R1473 B.n334 B.n161 163.367
R1474 B.n335 B.n334 163.367
R1475 B.n336 B.n335 163.367
R1476 B.n336 B.n159 163.367
R1477 B.n340 B.n159 163.367
R1478 B.n341 B.n340 163.367
R1479 B.n341 B.n155 163.367
R1480 B.n345 B.n155 163.367
R1481 B.n346 B.n345 163.367
R1482 B.n347 B.n346 163.367
R1483 B.n347 B.n153 163.367
R1484 B.n351 B.n153 163.367
R1485 B.n352 B.n351 163.367
R1486 B.n353 B.n352 163.367
R1487 B.n353 B.n149 163.367
R1488 B.n358 B.n149 163.367
R1489 B.n359 B.n358 163.367
R1490 B.n360 B.n359 163.367
R1491 B.n360 B.n147 163.367
R1492 B.n364 B.n147 163.367
R1493 B.n365 B.n364 163.367
R1494 B.n366 B.n365 163.367
R1495 B.n366 B.n145 163.367
R1496 B.n370 B.n145 163.367
R1497 B.n371 B.n370 163.367
R1498 B.n372 B.n371 163.367
R1499 B.n372 B.n143 163.367
R1500 B.n376 B.n143 163.367
R1501 B.n377 B.n376 163.367
R1502 B.n378 B.n377 163.367
R1503 B.n378 B.n141 163.367
R1504 B.n382 B.n141 163.367
R1505 B.n383 B.n382 163.367
R1506 B.n384 B.n383 163.367
R1507 B.n384 B.n139 163.367
R1508 B.n388 B.n139 163.367
R1509 B.n389 B.n388 163.367
R1510 B.n390 B.n389 163.367
R1511 B.n390 B.n137 163.367
R1512 B.n394 B.n137 163.367
R1513 B.n395 B.n394 163.367
R1514 B.n396 B.n395 163.367
R1515 B.n396 B.n135 163.367
R1516 B.n400 B.n135 163.367
R1517 B.n401 B.n400 163.367
R1518 B.n402 B.n401 163.367
R1519 B.n402 B.n133 163.367
R1520 B.n406 B.n133 163.367
R1521 B.n407 B.n406 163.367
R1522 B.n408 B.n407 163.367
R1523 B.n408 B.n131 163.367
R1524 B.n412 B.n131 163.367
R1525 B.n413 B.n412 163.367
R1526 B.n414 B.n413 163.367
R1527 B.n414 B.n129 163.367
R1528 B.n418 B.n129 163.367
R1529 B.n419 B.n418 163.367
R1530 B.n420 B.n419 163.367
R1531 B.n420 B.n127 163.367
R1532 B.n424 B.n127 163.367
R1533 B.n426 B.n425 163.367
R1534 B.n426 B.n125 163.367
R1535 B.n430 B.n125 163.367
R1536 B.n431 B.n430 163.367
R1537 B.n432 B.n431 163.367
R1538 B.n432 B.n123 163.367
R1539 B.n436 B.n123 163.367
R1540 B.n437 B.n436 163.367
R1541 B.n438 B.n437 163.367
R1542 B.n438 B.n121 163.367
R1543 B.n442 B.n121 163.367
R1544 B.n443 B.n442 163.367
R1545 B.n444 B.n443 163.367
R1546 B.n444 B.n119 163.367
R1547 B.n448 B.n119 163.367
R1548 B.n449 B.n448 163.367
R1549 B.n450 B.n449 163.367
R1550 B.n450 B.n117 163.367
R1551 B.n454 B.n117 163.367
R1552 B.n455 B.n454 163.367
R1553 B.n456 B.n455 163.367
R1554 B.n456 B.n115 163.367
R1555 B.n460 B.n115 163.367
R1556 B.n461 B.n460 163.367
R1557 B.n462 B.n461 163.367
R1558 B.n462 B.n113 163.367
R1559 B.n466 B.n113 163.367
R1560 B.n467 B.n466 163.367
R1561 B.n468 B.n467 163.367
R1562 B.n468 B.n111 163.367
R1563 B.n472 B.n111 163.367
R1564 B.n473 B.n472 163.367
R1565 B.n474 B.n473 163.367
R1566 B.n474 B.n109 163.367
R1567 B.n478 B.n109 163.367
R1568 B.n479 B.n478 163.367
R1569 B.n480 B.n479 163.367
R1570 B.n480 B.n107 163.367
R1571 B.n484 B.n107 163.367
R1572 B.n485 B.n484 163.367
R1573 B.n486 B.n485 163.367
R1574 B.n486 B.n105 163.367
R1575 B.n490 B.n105 163.367
R1576 B.n491 B.n490 163.367
R1577 B.n492 B.n491 163.367
R1578 B.n492 B.n103 163.367
R1579 B.n496 B.n103 163.367
R1580 B.n497 B.n496 163.367
R1581 B.n498 B.n497 163.367
R1582 B.n498 B.n101 163.367
R1583 B.n502 B.n101 163.367
R1584 B.n503 B.n502 163.367
R1585 B.n504 B.n503 163.367
R1586 B.n504 B.n99 163.367
R1587 B.n508 B.n99 163.367
R1588 B.n509 B.n508 163.367
R1589 B.n510 B.n509 163.367
R1590 B.n510 B.n97 163.367
R1591 B.n514 B.n97 163.367
R1592 B.n515 B.n514 163.367
R1593 B.n516 B.n515 163.367
R1594 B.n516 B.n95 163.367
R1595 B.n520 B.n95 163.367
R1596 B.n521 B.n520 163.367
R1597 B.n522 B.n521 163.367
R1598 B.n522 B.n93 163.367
R1599 B.n526 B.n93 163.367
R1600 B.n527 B.n526 163.367
R1601 B.n528 B.n527 163.367
R1602 B.n528 B.n91 163.367
R1603 B.n532 B.n91 163.367
R1604 B.n533 B.n532 163.367
R1605 B.n534 B.n533 163.367
R1606 B.n534 B.n89 163.367
R1607 B.n538 B.n89 163.367
R1608 B.n539 B.n538 163.367
R1609 B.n540 B.n539 163.367
R1610 B.n540 B.n87 163.367
R1611 B.n544 B.n87 163.367
R1612 B.n545 B.n544 163.367
R1613 B.n546 B.n545 163.367
R1614 B.n546 B.n85 163.367
R1615 B.n550 B.n85 163.367
R1616 B.n551 B.n550 163.367
R1617 B.n552 B.n551 163.367
R1618 B.n552 B.n83 163.367
R1619 B.n556 B.n83 163.367
R1620 B.n557 B.n556 163.367
R1621 B.n558 B.n557 163.367
R1622 B.n558 B.n81 163.367
R1623 B.n562 B.n81 163.367
R1624 B.n563 B.n562 163.367
R1625 B.n714 B.n25 163.367
R1626 B.n714 B.n713 163.367
R1627 B.n713 B.n712 163.367
R1628 B.n712 B.n27 163.367
R1629 B.n708 B.n27 163.367
R1630 B.n708 B.n707 163.367
R1631 B.n707 B.n706 163.367
R1632 B.n706 B.n29 163.367
R1633 B.n702 B.n29 163.367
R1634 B.n702 B.n701 163.367
R1635 B.n701 B.n700 163.367
R1636 B.n700 B.n31 163.367
R1637 B.n696 B.n31 163.367
R1638 B.n696 B.n695 163.367
R1639 B.n695 B.n694 163.367
R1640 B.n694 B.n33 163.367
R1641 B.n690 B.n33 163.367
R1642 B.n690 B.n689 163.367
R1643 B.n689 B.n688 163.367
R1644 B.n688 B.n35 163.367
R1645 B.n684 B.n35 163.367
R1646 B.n684 B.n683 163.367
R1647 B.n683 B.n682 163.367
R1648 B.n682 B.n37 163.367
R1649 B.n678 B.n37 163.367
R1650 B.n678 B.n677 163.367
R1651 B.n677 B.n676 163.367
R1652 B.n676 B.n39 163.367
R1653 B.n672 B.n39 163.367
R1654 B.n672 B.n671 163.367
R1655 B.n671 B.n670 163.367
R1656 B.n670 B.n41 163.367
R1657 B.n666 B.n41 163.367
R1658 B.n666 B.n665 163.367
R1659 B.n665 B.n664 163.367
R1660 B.n664 B.n43 163.367
R1661 B.n660 B.n43 163.367
R1662 B.n660 B.n659 163.367
R1663 B.n659 B.n658 163.367
R1664 B.n658 B.n45 163.367
R1665 B.n654 B.n45 163.367
R1666 B.n654 B.n653 163.367
R1667 B.n653 B.n652 163.367
R1668 B.n652 B.n47 163.367
R1669 B.n648 B.n47 163.367
R1670 B.n648 B.n647 163.367
R1671 B.n647 B.n51 163.367
R1672 B.n643 B.n51 163.367
R1673 B.n643 B.n642 163.367
R1674 B.n642 B.n641 163.367
R1675 B.n641 B.n53 163.367
R1676 B.n637 B.n53 163.367
R1677 B.n637 B.n636 163.367
R1678 B.n636 B.n635 163.367
R1679 B.n635 B.n55 163.367
R1680 B.n630 B.n55 163.367
R1681 B.n630 B.n629 163.367
R1682 B.n629 B.n628 163.367
R1683 B.n628 B.n59 163.367
R1684 B.n624 B.n59 163.367
R1685 B.n624 B.n623 163.367
R1686 B.n623 B.n622 163.367
R1687 B.n622 B.n61 163.367
R1688 B.n618 B.n61 163.367
R1689 B.n618 B.n617 163.367
R1690 B.n617 B.n616 163.367
R1691 B.n616 B.n63 163.367
R1692 B.n612 B.n63 163.367
R1693 B.n612 B.n611 163.367
R1694 B.n611 B.n610 163.367
R1695 B.n610 B.n65 163.367
R1696 B.n606 B.n65 163.367
R1697 B.n606 B.n605 163.367
R1698 B.n605 B.n604 163.367
R1699 B.n604 B.n67 163.367
R1700 B.n600 B.n67 163.367
R1701 B.n600 B.n599 163.367
R1702 B.n599 B.n598 163.367
R1703 B.n598 B.n69 163.367
R1704 B.n594 B.n69 163.367
R1705 B.n594 B.n593 163.367
R1706 B.n593 B.n592 163.367
R1707 B.n592 B.n71 163.367
R1708 B.n588 B.n71 163.367
R1709 B.n588 B.n587 163.367
R1710 B.n587 B.n586 163.367
R1711 B.n586 B.n73 163.367
R1712 B.n582 B.n73 163.367
R1713 B.n582 B.n581 163.367
R1714 B.n581 B.n580 163.367
R1715 B.n580 B.n75 163.367
R1716 B.n576 B.n75 163.367
R1717 B.n576 B.n575 163.367
R1718 B.n575 B.n574 163.367
R1719 B.n574 B.n77 163.367
R1720 B.n570 B.n77 163.367
R1721 B.n570 B.n569 163.367
R1722 B.n569 B.n568 163.367
R1723 B.n568 B.n79 163.367
R1724 B.n564 B.n79 163.367
R1725 B.n151 B.n150 83.2005
R1726 B.n157 B.n156 83.2005
R1727 B.n49 B.n48 83.2005
R1728 B.n57 B.n56 83.2005
R1729 B.n355 B.n151 59.5399
R1730 B.n158 B.n157 59.5399
R1731 B.n50 B.n49 59.5399
R1732 B.n633 B.n57 59.5399
R1733 B.n717 B.n716 33.8737
R1734 B.n565 B.n80 33.8737
R1735 B.n423 B.n126 33.8737
R1736 B.n272 B.n271 33.8737
R1737 B B.n787 18.0485
R1738 B.n716 B.n715 10.6151
R1739 B.n715 B.n26 10.6151
R1740 B.n711 B.n26 10.6151
R1741 B.n711 B.n710 10.6151
R1742 B.n710 B.n709 10.6151
R1743 B.n709 B.n28 10.6151
R1744 B.n705 B.n28 10.6151
R1745 B.n705 B.n704 10.6151
R1746 B.n704 B.n703 10.6151
R1747 B.n703 B.n30 10.6151
R1748 B.n699 B.n30 10.6151
R1749 B.n699 B.n698 10.6151
R1750 B.n698 B.n697 10.6151
R1751 B.n697 B.n32 10.6151
R1752 B.n693 B.n32 10.6151
R1753 B.n693 B.n692 10.6151
R1754 B.n692 B.n691 10.6151
R1755 B.n691 B.n34 10.6151
R1756 B.n687 B.n34 10.6151
R1757 B.n687 B.n686 10.6151
R1758 B.n686 B.n685 10.6151
R1759 B.n685 B.n36 10.6151
R1760 B.n681 B.n36 10.6151
R1761 B.n681 B.n680 10.6151
R1762 B.n680 B.n679 10.6151
R1763 B.n679 B.n38 10.6151
R1764 B.n675 B.n38 10.6151
R1765 B.n675 B.n674 10.6151
R1766 B.n674 B.n673 10.6151
R1767 B.n673 B.n40 10.6151
R1768 B.n669 B.n40 10.6151
R1769 B.n669 B.n668 10.6151
R1770 B.n668 B.n667 10.6151
R1771 B.n667 B.n42 10.6151
R1772 B.n663 B.n42 10.6151
R1773 B.n663 B.n662 10.6151
R1774 B.n662 B.n661 10.6151
R1775 B.n661 B.n44 10.6151
R1776 B.n657 B.n44 10.6151
R1777 B.n657 B.n656 10.6151
R1778 B.n656 B.n655 10.6151
R1779 B.n655 B.n46 10.6151
R1780 B.n651 B.n46 10.6151
R1781 B.n651 B.n650 10.6151
R1782 B.n650 B.n649 10.6151
R1783 B.n646 B.n645 10.6151
R1784 B.n645 B.n644 10.6151
R1785 B.n644 B.n52 10.6151
R1786 B.n640 B.n52 10.6151
R1787 B.n640 B.n639 10.6151
R1788 B.n639 B.n638 10.6151
R1789 B.n638 B.n54 10.6151
R1790 B.n634 B.n54 10.6151
R1791 B.n632 B.n631 10.6151
R1792 B.n631 B.n58 10.6151
R1793 B.n627 B.n58 10.6151
R1794 B.n627 B.n626 10.6151
R1795 B.n626 B.n625 10.6151
R1796 B.n625 B.n60 10.6151
R1797 B.n621 B.n60 10.6151
R1798 B.n621 B.n620 10.6151
R1799 B.n620 B.n619 10.6151
R1800 B.n619 B.n62 10.6151
R1801 B.n615 B.n62 10.6151
R1802 B.n615 B.n614 10.6151
R1803 B.n614 B.n613 10.6151
R1804 B.n613 B.n64 10.6151
R1805 B.n609 B.n64 10.6151
R1806 B.n609 B.n608 10.6151
R1807 B.n608 B.n607 10.6151
R1808 B.n607 B.n66 10.6151
R1809 B.n603 B.n66 10.6151
R1810 B.n603 B.n602 10.6151
R1811 B.n602 B.n601 10.6151
R1812 B.n601 B.n68 10.6151
R1813 B.n597 B.n68 10.6151
R1814 B.n597 B.n596 10.6151
R1815 B.n596 B.n595 10.6151
R1816 B.n595 B.n70 10.6151
R1817 B.n591 B.n70 10.6151
R1818 B.n591 B.n590 10.6151
R1819 B.n590 B.n589 10.6151
R1820 B.n589 B.n72 10.6151
R1821 B.n585 B.n72 10.6151
R1822 B.n585 B.n584 10.6151
R1823 B.n584 B.n583 10.6151
R1824 B.n583 B.n74 10.6151
R1825 B.n579 B.n74 10.6151
R1826 B.n579 B.n578 10.6151
R1827 B.n578 B.n577 10.6151
R1828 B.n577 B.n76 10.6151
R1829 B.n573 B.n76 10.6151
R1830 B.n573 B.n572 10.6151
R1831 B.n572 B.n571 10.6151
R1832 B.n571 B.n78 10.6151
R1833 B.n567 B.n78 10.6151
R1834 B.n567 B.n566 10.6151
R1835 B.n566 B.n565 10.6151
R1836 B.n427 B.n126 10.6151
R1837 B.n428 B.n427 10.6151
R1838 B.n429 B.n428 10.6151
R1839 B.n429 B.n124 10.6151
R1840 B.n433 B.n124 10.6151
R1841 B.n434 B.n433 10.6151
R1842 B.n435 B.n434 10.6151
R1843 B.n435 B.n122 10.6151
R1844 B.n439 B.n122 10.6151
R1845 B.n440 B.n439 10.6151
R1846 B.n441 B.n440 10.6151
R1847 B.n441 B.n120 10.6151
R1848 B.n445 B.n120 10.6151
R1849 B.n446 B.n445 10.6151
R1850 B.n447 B.n446 10.6151
R1851 B.n447 B.n118 10.6151
R1852 B.n451 B.n118 10.6151
R1853 B.n452 B.n451 10.6151
R1854 B.n453 B.n452 10.6151
R1855 B.n453 B.n116 10.6151
R1856 B.n457 B.n116 10.6151
R1857 B.n458 B.n457 10.6151
R1858 B.n459 B.n458 10.6151
R1859 B.n459 B.n114 10.6151
R1860 B.n463 B.n114 10.6151
R1861 B.n464 B.n463 10.6151
R1862 B.n465 B.n464 10.6151
R1863 B.n465 B.n112 10.6151
R1864 B.n469 B.n112 10.6151
R1865 B.n470 B.n469 10.6151
R1866 B.n471 B.n470 10.6151
R1867 B.n471 B.n110 10.6151
R1868 B.n475 B.n110 10.6151
R1869 B.n476 B.n475 10.6151
R1870 B.n477 B.n476 10.6151
R1871 B.n477 B.n108 10.6151
R1872 B.n481 B.n108 10.6151
R1873 B.n482 B.n481 10.6151
R1874 B.n483 B.n482 10.6151
R1875 B.n483 B.n106 10.6151
R1876 B.n487 B.n106 10.6151
R1877 B.n488 B.n487 10.6151
R1878 B.n489 B.n488 10.6151
R1879 B.n489 B.n104 10.6151
R1880 B.n493 B.n104 10.6151
R1881 B.n494 B.n493 10.6151
R1882 B.n495 B.n494 10.6151
R1883 B.n495 B.n102 10.6151
R1884 B.n499 B.n102 10.6151
R1885 B.n500 B.n499 10.6151
R1886 B.n501 B.n500 10.6151
R1887 B.n501 B.n100 10.6151
R1888 B.n505 B.n100 10.6151
R1889 B.n506 B.n505 10.6151
R1890 B.n507 B.n506 10.6151
R1891 B.n507 B.n98 10.6151
R1892 B.n511 B.n98 10.6151
R1893 B.n512 B.n511 10.6151
R1894 B.n513 B.n512 10.6151
R1895 B.n513 B.n96 10.6151
R1896 B.n517 B.n96 10.6151
R1897 B.n518 B.n517 10.6151
R1898 B.n519 B.n518 10.6151
R1899 B.n519 B.n94 10.6151
R1900 B.n523 B.n94 10.6151
R1901 B.n524 B.n523 10.6151
R1902 B.n525 B.n524 10.6151
R1903 B.n525 B.n92 10.6151
R1904 B.n529 B.n92 10.6151
R1905 B.n530 B.n529 10.6151
R1906 B.n531 B.n530 10.6151
R1907 B.n531 B.n90 10.6151
R1908 B.n535 B.n90 10.6151
R1909 B.n536 B.n535 10.6151
R1910 B.n537 B.n536 10.6151
R1911 B.n537 B.n88 10.6151
R1912 B.n541 B.n88 10.6151
R1913 B.n542 B.n541 10.6151
R1914 B.n543 B.n542 10.6151
R1915 B.n543 B.n86 10.6151
R1916 B.n547 B.n86 10.6151
R1917 B.n548 B.n547 10.6151
R1918 B.n549 B.n548 10.6151
R1919 B.n549 B.n84 10.6151
R1920 B.n553 B.n84 10.6151
R1921 B.n554 B.n553 10.6151
R1922 B.n555 B.n554 10.6151
R1923 B.n555 B.n82 10.6151
R1924 B.n559 B.n82 10.6151
R1925 B.n560 B.n559 10.6151
R1926 B.n561 B.n560 10.6151
R1927 B.n561 B.n80 10.6151
R1928 B.n273 B.n272 10.6151
R1929 B.n273 B.n180 10.6151
R1930 B.n277 B.n180 10.6151
R1931 B.n278 B.n277 10.6151
R1932 B.n279 B.n278 10.6151
R1933 B.n279 B.n178 10.6151
R1934 B.n283 B.n178 10.6151
R1935 B.n284 B.n283 10.6151
R1936 B.n285 B.n284 10.6151
R1937 B.n285 B.n176 10.6151
R1938 B.n289 B.n176 10.6151
R1939 B.n290 B.n289 10.6151
R1940 B.n291 B.n290 10.6151
R1941 B.n291 B.n174 10.6151
R1942 B.n295 B.n174 10.6151
R1943 B.n296 B.n295 10.6151
R1944 B.n297 B.n296 10.6151
R1945 B.n297 B.n172 10.6151
R1946 B.n301 B.n172 10.6151
R1947 B.n302 B.n301 10.6151
R1948 B.n303 B.n302 10.6151
R1949 B.n303 B.n170 10.6151
R1950 B.n307 B.n170 10.6151
R1951 B.n308 B.n307 10.6151
R1952 B.n309 B.n308 10.6151
R1953 B.n309 B.n168 10.6151
R1954 B.n313 B.n168 10.6151
R1955 B.n314 B.n313 10.6151
R1956 B.n315 B.n314 10.6151
R1957 B.n315 B.n166 10.6151
R1958 B.n319 B.n166 10.6151
R1959 B.n320 B.n319 10.6151
R1960 B.n321 B.n320 10.6151
R1961 B.n321 B.n164 10.6151
R1962 B.n325 B.n164 10.6151
R1963 B.n326 B.n325 10.6151
R1964 B.n327 B.n326 10.6151
R1965 B.n327 B.n162 10.6151
R1966 B.n331 B.n162 10.6151
R1967 B.n332 B.n331 10.6151
R1968 B.n333 B.n332 10.6151
R1969 B.n333 B.n160 10.6151
R1970 B.n337 B.n160 10.6151
R1971 B.n338 B.n337 10.6151
R1972 B.n339 B.n338 10.6151
R1973 B.n343 B.n342 10.6151
R1974 B.n344 B.n343 10.6151
R1975 B.n344 B.n154 10.6151
R1976 B.n348 B.n154 10.6151
R1977 B.n349 B.n348 10.6151
R1978 B.n350 B.n349 10.6151
R1979 B.n350 B.n152 10.6151
R1980 B.n354 B.n152 10.6151
R1981 B.n357 B.n356 10.6151
R1982 B.n357 B.n148 10.6151
R1983 B.n361 B.n148 10.6151
R1984 B.n362 B.n361 10.6151
R1985 B.n363 B.n362 10.6151
R1986 B.n363 B.n146 10.6151
R1987 B.n367 B.n146 10.6151
R1988 B.n368 B.n367 10.6151
R1989 B.n369 B.n368 10.6151
R1990 B.n369 B.n144 10.6151
R1991 B.n373 B.n144 10.6151
R1992 B.n374 B.n373 10.6151
R1993 B.n375 B.n374 10.6151
R1994 B.n375 B.n142 10.6151
R1995 B.n379 B.n142 10.6151
R1996 B.n380 B.n379 10.6151
R1997 B.n381 B.n380 10.6151
R1998 B.n381 B.n140 10.6151
R1999 B.n385 B.n140 10.6151
R2000 B.n386 B.n385 10.6151
R2001 B.n387 B.n386 10.6151
R2002 B.n387 B.n138 10.6151
R2003 B.n391 B.n138 10.6151
R2004 B.n392 B.n391 10.6151
R2005 B.n393 B.n392 10.6151
R2006 B.n393 B.n136 10.6151
R2007 B.n397 B.n136 10.6151
R2008 B.n398 B.n397 10.6151
R2009 B.n399 B.n398 10.6151
R2010 B.n399 B.n134 10.6151
R2011 B.n403 B.n134 10.6151
R2012 B.n404 B.n403 10.6151
R2013 B.n405 B.n404 10.6151
R2014 B.n405 B.n132 10.6151
R2015 B.n409 B.n132 10.6151
R2016 B.n410 B.n409 10.6151
R2017 B.n411 B.n410 10.6151
R2018 B.n411 B.n130 10.6151
R2019 B.n415 B.n130 10.6151
R2020 B.n416 B.n415 10.6151
R2021 B.n417 B.n416 10.6151
R2022 B.n417 B.n128 10.6151
R2023 B.n421 B.n128 10.6151
R2024 B.n422 B.n421 10.6151
R2025 B.n423 B.n422 10.6151
R2026 B.n271 B.n182 10.6151
R2027 B.n267 B.n182 10.6151
R2028 B.n267 B.n266 10.6151
R2029 B.n266 B.n265 10.6151
R2030 B.n265 B.n184 10.6151
R2031 B.n261 B.n184 10.6151
R2032 B.n261 B.n260 10.6151
R2033 B.n260 B.n259 10.6151
R2034 B.n259 B.n186 10.6151
R2035 B.n255 B.n186 10.6151
R2036 B.n255 B.n254 10.6151
R2037 B.n254 B.n253 10.6151
R2038 B.n253 B.n188 10.6151
R2039 B.n249 B.n188 10.6151
R2040 B.n249 B.n248 10.6151
R2041 B.n248 B.n247 10.6151
R2042 B.n247 B.n190 10.6151
R2043 B.n243 B.n190 10.6151
R2044 B.n243 B.n242 10.6151
R2045 B.n242 B.n241 10.6151
R2046 B.n241 B.n192 10.6151
R2047 B.n237 B.n192 10.6151
R2048 B.n237 B.n236 10.6151
R2049 B.n236 B.n235 10.6151
R2050 B.n235 B.n194 10.6151
R2051 B.n231 B.n194 10.6151
R2052 B.n231 B.n230 10.6151
R2053 B.n230 B.n229 10.6151
R2054 B.n229 B.n196 10.6151
R2055 B.n225 B.n196 10.6151
R2056 B.n225 B.n224 10.6151
R2057 B.n224 B.n223 10.6151
R2058 B.n223 B.n198 10.6151
R2059 B.n219 B.n198 10.6151
R2060 B.n219 B.n218 10.6151
R2061 B.n218 B.n217 10.6151
R2062 B.n217 B.n200 10.6151
R2063 B.n213 B.n200 10.6151
R2064 B.n213 B.n212 10.6151
R2065 B.n212 B.n211 10.6151
R2066 B.n211 B.n202 10.6151
R2067 B.n207 B.n202 10.6151
R2068 B.n207 B.n206 10.6151
R2069 B.n206 B.n205 10.6151
R2070 B.n205 B.n0 10.6151
R2071 B.n783 B.n1 10.6151
R2072 B.n783 B.n782 10.6151
R2073 B.n782 B.n781 10.6151
R2074 B.n781 B.n4 10.6151
R2075 B.n777 B.n4 10.6151
R2076 B.n777 B.n776 10.6151
R2077 B.n776 B.n775 10.6151
R2078 B.n775 B.n6 10.6151
R2079 B.n771 B.n6 10.6151
R2080 B.n771 B.n770 10.6151
R2081 B.n770 B.n769 10.6151
R2082 B.n769 B.n8 10.6151
R2083 B.n765 B.n8 10.6151
R2084 B.n765 B.n764 10.6151
R2085 B.n764 B.n763 10.6151
R2086 B.n763 B.n10 10.6151
R2087 B.n759 B.n10 10.6151
R2088 B.n759 B.n758 10.6151
R2089 B.n758 B.n757 10.6151
R2090 B.n757 B.n12 10.6151
R2091 B.n753 B.n12 10.6151
R2092 B.n753 B.n752 10.6151
R2093 B.n752 B.n751 10.6151
R2094 B.n751 B.n14 10.6151
R2095 B.n747 B.n14 10.6151
R2096 B.n747 B.n746 10.6151
R2097 B.n746 B.n745 10.6151
R2098 B.n745 B.n16 10.6151
R2099 B.n741 B.n16 10.6151
R2100 B.n741 B.n740 10.6151
R2101 B.n740 B.n739 10.6151
R2102 B.n739 B.n18 10.6151
R2103 B.n735 B.n18 10.6151
R2104 B.n735 B.n734 10.6151
R2105 B.n734 B.n733 10.6151
R2106 B.n733 B.n20 10.6151
R2107 B.n729 B.n20 10.6151
R2108 B.n729 B.n728 10.6151
R2109 B.n728 B.n727 10.6151
R2110 B.n727 B.n22 10.6151
R2111 B.n723 B.n22 10.6151
R2112 B.n723 B.n722 10.6151
R2113 B.n722 B.n721 10.6151
R2114 B.n721 B.n24 10.6151
R2115 B.n717 B.n24 10.6151
R2116 B.n646 B.n50 6.5566
R2117 B.n634 B.n633 6.5566
R2118 B.n342 B.n158 6.5566
R2119 B.n355 B.n354 6.5566
R2120 B.n649 B.n50 4.05904
R2121 B.n633 B.n632 4.05904
R2122 B.n339 B.n158 4.05904
R2123 B.n356 B.n355 4.05904
R2124 B.n787 B.n0 2.81026
R2125 B.n787 B.n1 2.81026
R2126 VN.n0 VN.t0 115.668
R2127 VN.n1 VN.t1 115.668
R2128 VN.n0 VN.t3 114.231
R2129 VN.n1 VN.t2 114.231
R2130 VN VN.n1 53.4821
R2131 VN VN.n0 1.75857
R2132 VDD2.n2 VDD2.n0 116.552
R2133 VDD2.n2 VDD2.n1 70.1474
R2134 VDD2.n1 VDD2.t1 2.41723
R2135 VDD2.n1 VDD2.t2 2.41723
R2136 VDD2.n0 VDD2.t3 2.41723
R2137 VDD2.n0 VDD2.t0 2.41723
R2138 VDD2 VDD2.n2 0.0586897
C0 B w_n3544_n3658# 11.3248f
C1 VP B 2.15172f
C2 B VDD2 1.61669f
C3 B VN 1.38364f
C4 VTAIL B 5.9898f
C5 VP w_n3544_n3658# 6.74538f
C6 B VDD1 1.54204f
C7 VDD2 w_n3544_n3658# 1.83387f
C8 VN w_n3544_n3658# 6.28634f
C9 VP VDD2 0.481003f
C10 VP VN 7.44318f
C11 VTAIL w_n3544_n3658# 4.32887f
C12 VDD2 VN 5.62662f
C13 VTAIL VP 5.68646f
C14 VDD1 w_n3544_n3658# 1.74778f
C15 VTAIL VDD2 6.17081f
C16 VTAIL VN 5.67235f
C17 VP VDD1 5.95615f
C18 VDD2 VDD1 1.36149f
C19 VDD1 VN 0.150387f
C20 VTAIL VDD1 6.10748f
C21 VDD2 VSUBS 1.196307f
C22 VDD1 VSUBS 6.7278f
C23 VTAIL VSUBS 1.466549f
C24 VN VSUBS 6.26143f
C25 VP VSUBS 3.075146f
C26 B VSUBS 5.568861f
C27 w_n3544_n3658# VSUBS 0.159267p
C28 VDD2.t3 VSUBS 0.289092f
C29 VDD2.t0 VSUBS 0.289092f
C30 VDD2.n0 VSUBS 3.16253f
C31 VDD2.t1 VSUBS 0.289092f
C32 VDD2.t2 VSUBS 0.289092f
C33 VDD2.n1 VSUBS 2.28815f
C34 VDD2.n2 VSUBS 4.86296f
C35 VN.t0 VSUBS 4.12448f
C36 VN.t3 VSUBS 4.10679f
C37 VN.n0 VSUBS 2.4598f
C38 VN.t1 VSUBS 4.12448f
C39 VN.t2 VSUBS 4.10679f
C40 VN.n1 VSUBS 4.20075f
C41 B.n0 VSUBS 0.004182f
C42 B.n1 VSUBS 0.004182f
C43 B.n2 VSUBS 0.006613f
C44 B.n3 VSUBS 0.006613f
C45 B.n4 VSUBS 0.006613f
C46 B.n5 VSUBS 0.006613f
C47 B.n6 VSUBS 0.006613f
C48 B.n7 VSUBS 0.006613f
C49 B.n8 VSUBS 0.006613f
C50 B.n9 VSUBS 0.006613f
C51 B.n10 VSUBS 0.006613f
C52 B.n11 VSUBS 0.006613f
C53 B.n12 VSUBS 0.006613f
C54 B.n13 VSUBS 0.006613f
C55 B.n14 VSUBS 0.006613f
C56 B.n15 VSUBS 0.006613f
C57 B.n16 VSUBS 0.006613f
C58 B.n17 VSUBS 0.006613f
C59 B.n18 VSUBS 0.006613f
C60 B.n19 VSUBS 0.006613f
C61 B.n20 VSUBS 0.006613f
C62 B.n21 VSUBS 0.006613f
C63 B.n22 VSUBS 0.006613f
C64 B.n23 VSUBS 0.006613f
C65 B.n24 VSUBS 0.006613f
C66 B.n25 VSUBS 0.016081f
C67 B.n26 VSUBS 0.006613f
C68 B.n27 VSUBS 0.006613f
C69 B.n28 VSUBS 0.006613f
C70 B.n29 VSUBS 0.006613f
C71 B.n30 VSUBS 0.006613f
C72 B.n31 VSUBS 0.006613f
C73 B.n32 VSUBS 0.006613f
C74 B.n33 VSUBS 0.006613f
C75 B.n34 VSUBS 0.006613f
C76 B.n35 VSUBS 0.006613f
C77 B.n36 VSUBS 0.006613f
C78 B.n37 VSUBS 0.006613f
C79 B.n38 VSUBS 0.006613f
C80 B.n39 VSUBS 0.006613f
C81 B.n40 VSUBS 0.006613f
C82 B.n41 VSUBS 0.006613f
C83 B.n42 VSUBS 0.006613f
C84 B.n43 VSUBS 0.006613f
C85 B.n44 VSUBS 0.006613f
C86 B.n45 VSUBS 0.006613f
C87 B.n46 VSUBS 0.006613f
C88 B.n47 VSUBS 0.006613f
C89 B.t8 VSUBS 0.230294f
C90 B.t7 VSUBS 0.273592f
C91 B.t6 VSUBS 2.33799f
C92 B.n48 VSUBS 0.436479f
C93 B.n49 VSUBS 0.261813f
C94 B.n50 VSUBS 0.015321f
C95 B.n51 VSUBS 0.006613f
C96 B.n52 VSUBS 0.006613f
C97 B.n53 VSUBS 0.006613f
C98 B.n54 VSUBS 0.006613f
C99 B.n55 VSUBS 0.006613f
C100 B.t5 VSUBS 0.230297f
C101 B.t4 VSUBS 0.273595f
C102 B.t3 VSUBS 2.33799f
C103 B.n56 VSUBS 0.436476f
C104 B.n57 VSUBS 0.26181f
C105 B.n58 VSUBS 0.006613f
C106 B.n59 VSUBS 0.006613f
C107 B.n60 VSUBS 0.006613f
C108 B.n61 VSUBS 0.006613f
C109 B.n62 VSUBS 0.006613f
C110 B.n63 VSUBS 0.006613f
C111 B.n64 VSUBS 0.006613f
C112 B.n65 VSUBS 0.006613f
C113 B.n66 VSUBS 0.006613f
C114 B.n67 VSUBS 0.006613f
C115 B.n68 VSUBS 0.006613f
C116 B.n69 VSUBS 0.006613f
C117 B.n70 VSUBS 0.006613f
C118 B.n71 VSUBS 0.006613f
C119 B.n72 VSUBS 0.006613f
C120 B.n73 VSUBS 0.006613f
C121 B.n74 VSUBS 0.006613f
C122 B.n75 VSUBS 0.006613f
C123 B.n76 VSUBS 0.006613f
C124 B.n77 VSUBS 0.006613f
C125 B.n78 VSUBS 0.006613f
C126 B.n79 VSUBS 0.006613f
C127 B.n80 VSUBS 0.016375f
C128 B.n81 VSUBS 0.006613f
C129 B.n82 VSUBS 0.006613f
C130 B.n83 VSUBS 0.006613f
C131 B.n84 VSUBS 0.006613f
C132 B.n85 VSUBS 0.006613f
C133 B.n86 VSUBS 0.006613f
C134 B.n87 VSUBS 0.006613f
C135 B.n88 VSUBS 0.006613f
C136 B.n89 VSUBS 0.006613f
C137 B.n90 VSUBS 0.006613f
C138 B.n91 VSUBS 0.006613f
C139 B.n92 VSUBS 0.006613f
C140 B.n93 VSUBS 0.006613f
C141 B.n94 VSUBS 0.006613f
C142 B.n95 VSUBS 0.006613f
C143 B.n96 VSUBS 0.006613f
C144 B.n97 VSUBS 0.006613f
C145 B.n98 VSUBS 0.006613f
C146 B.n99 VSUBS 0.006613f
C147 B.n100 VSUBS 0.006613f
C148 B.n101 VSUBS 0.006613f
C149 B.n102 VSUBS 0.006613f
C150 B.n103 VSUBS 0.006613f
C151 B.n104 VSUBS 0.006613f
C152 B.n105 VSUBS 0.006613f
C153 B.n106 VSUBS 0.006613f
C154 B.n107 VSUBS 0.006613f
C155 B.n108 VSUBS 0.006613f
C156 B.n109 VSUBS 0.006613f
C157 B.n110 VSUBS 0.006613f
C158 B.n111 VSUBS 0.006613f
C159 B.n112 VSUBS 0.006613f
C160 B.n113 VSUBS 0.006613f
C161 B.n114 VSUBS 0.006613f
C162 B.n115 VSUBS 0.006613f
C163 B.n116 VSUBS 0.006613f
C164 B.n117 VSUBS 0.006613f
C165 B.n118 VSUBS 0.006613f
C166 B.n119 VSUBS 0.006613f
C167 B.n120 VSUBS 0.006613f
C168 B.n121 VSUBS 0.006613f
C169 B.n122 VSUBS 0.006613f
C170 B.n123 VSUBS 0.006613f
C171 B.n124 VSUBS 0.006613f
C172 B.n125 VSUBS 0.006613f
C173 B.n126 VSUBS 0.015622f
C174 B.n127 VSUBS 0.006613f
C175 B.n128 VSUBS 0.006613f
C176 B.n129 VSUBS 0.006613f
C177 B.n130 VSUBS 0.006613f
C178 B.n131 VSUBS 0.006613f
C179 B.n132 VSUBS 0.006613f
C180 B.n133 VSUBS 0.006613f
C181 B.n134 VSUBS 0.006613f
C182 B.n135 VSUBS 0.006613f
C183 B.n136 VSUBS 0.006613f
C184 B.n137 VSUBS 0.006613f
C185 B.n138 VSUBS 0.006613f
C186 B.n139 VSUBS 0.006613f
C187 B.n140 VSUBS 0.006613f
C188 B.n141 VSUBS 0.006613f
C189 B.n142 VSUBS 0.006613f
C190 B.n143 VSUBS 0.006613f
C191 B.n144 VSUBS 0.006613f
C192 B.n145 VSUBS 0.006613f
C193 B.n146 VSUBS 0.006613f
C194 B.n147 VSUBS 0.006613f
C195 B.n148 VSUBS 0.006613f
C196 B.n149 VSUBS 0.006613f
C197 B.t10 VSUBS 0.230297f
C198 B.t11 VSUBS 0.273595f
C199 B.t9 VSUBS 2.33799f
C200 B.n150 VSUBS 0.436476f
C201 B.n151 VSUBS 0.26181f
C202 B.n152 VSUBS 0.006613f
C203 B.n153 VSUBS 0.006613f
C204 B.n154 VSUBS 0.006613f
C205 B.n155 VSUBS 0.006613f
C206 B.t1 VSUBS 0.230294f
C207 B.t2 VSUBS 0.273592f
C208 B.t0 VSUBS 2.33799f
C209 B.n156 VSUBS 0.436479f
C210 B.n157 VSUBS 0.261813f
C211 B.n158 VSUBS 0.015321f
C212 B.n159 VSUBS 0.006613f
C213 B.n160 VSUBS 0.006613f
C214 B.n161 VSUBS 0.006613f
C215 B.n162 VSUBS 0.006613f
C216 B.n163 VSUBS 0.006613f
C217 B.n164 VSUBS 0.006613f
C218 B.n165 VSUBS 0.006613f
C219 B.n166 VSUBS 0.006613f
C220 B.n167 VSUBS 0.006613f
C221 B.n168 VSUBS 0.006613f
C222 B.n169 VSUBS 0.006613f
C223 B.n170 VSUBS 0.006613f
C224 B.n171 VSUBS 0.006613f
C225 B.n172 VSUBS 0.006613f
C226 B.n173 VSUBS 0.006613f
C227 B.n174 VSUBS 0.006613f
C228 B.n175 VSUBS 0.006613f
C229 B.n176 VSUBS 0.006613f
C230 B.n177 VSUBS 0.006613f
C231 B.n178 VSUBS 0.006613f
C232 B.n179 VSUBS 0.006613f
C233 B.n180 VSUBS 0.006613f
C234 B.n181 VSUBS 0.016081f
C235 B.n182 VSUBS 0.006613f
C236 B.n183 VSUBS 0.006613f
C237 B.n184 VSUBS 0.006613f
C238 B.n185 VSUBS 0.006613f
C239 B.n186 VSUBS 0.006613f
C240 B.n187 VSUBS 0.006613f
C241 B.n188 VSUBS 0.006613f
C242 B.n189 VSUBS 0.006613f
C243 B.n190 VSUBS 0.006613f
C244 B.n191 VSUBS 0.006613f
C245 B.n192 VSUBS 0.006613f
C246 B.n193 VSUBS 0.006613f
C247 B.n194 VSUBS 0.006613f
C248 B.n195 VSUBS 0.006613f
C249 B.n196 VSUBS 0.006613f
C250 B.n197 VSUBS 0.006613f
C251 B.n198 VSUBS 0.006613f
C252 B.n199 VSUBS 0.006613f
C253 B.n200 VSUBS 0.006613f
C254 B.n201 VSUBS 0.006613f
C255 B.n202 VSUBS 0.006613f
C256 B.n203 VSUBS 0.006613f
C257 B.n204 VSUBS 0.006613f
C258 B.n205 VSUBS 0.006613f
C259 B.n206 VSUBS 0.006613f
C260 B.n207 VSUBS 0.006613f
C261 B.n208 VSUBS 0.006613f
C262 B.n209 VSUBS 0.006613f
C263 B.n210 VSUBS 0.006613f
C264 B.n211 VSUBS 0.006613f
C265 B.n212 VSUBS 0.006613f
C266 B.n213 VSUBS 0.006613f
C267 B.n214 VSUBS 0.006613f
C268 B.n215 VSUBS 0.006613f
C269 B.n216 VSUBS 0.006613f
C270 B.n217 VSUBS 0.006613f
C271 B.n218 VSUBS 0.006613f
C272 B.n219 VSUBS 0.006613f
C273 B.n220 VSUBS 0.006613f
C274 B.n221 VSUBS 0.006613f
C275 B.n222 VSUBS 0.006613f
C276 B.n223 VSUBS 0.006613f
C277 B.n224 VSUBS 0.006613f
C278 B.n225 VSUBS 0.006613f
C279 B.n226 VSUBS 0.006613f
C280 B.n227 VSUBS 0.006613f
C281 B.n228 VSUBS 0.006613f
C282 B.n229 VSUBS 0.006613f
C283 B.n230 VSUBS 0.006613f
C284 B.n231 VSUBS 0.006613f
C285 B.n232 VSUBS 0.006613f
C286 B.n233 VSUBS 0.006613f
C287 B.n234 VSUBS 0.006613f
C288 B.n235 VSUBS 0.006613f
C289 B.n236 VSUBS 0.006613f
C290 B.n237 VSUBS 0.006613f
C291 B.n238 VSUBS 0.006613f
C292 B.n239 VSUBS 0.006613f
C293 B.n240 VSUBS 0.006613f
C294 B.n241 VSUBS 0.006613f
C295 B.n242 VSUBS 0.006613f
C296 B.n243 VSUBS 0.006613f
C297 B.n244 VSUBS 0.006613f
C298 B.n245 VSUBS 0.006613f
C299 B.n246 VSUBS 0.006613f
C300 B.n247 VSUBS 0.006613f
C301 B.n248 VSUBS 0.006613f
C302 B.n249 VSUBS 0.006613f
C303 B.n250 VSUBS 0.006613f
C304 B.n251 VSUBS 0.006613f
C305 B.n252 VSUBS 0.006613f
C306 B.n253 VSUBS 0.006613f
C307 B.n254 VSUBS 0.006613f
C308 B.n255 VSUBS 0.006613f
C309 B.n256 VSUBS 0.006613f
C310 B.n257 VSUBS 0.006613f
C311 B.n258 VSUBS 0.006613f
C312 B.n259 VSUBS 0.006613f
C313 B.n260 VSUBS 0.006613f
C314 B.n261 VSUBS 0.006613f
C315 B.n262 VSUBS 0.006613f
C316 B.n263 VSUBS 0.006613f
C317 B.n264 VSUBS 0.006613f
C318 B.n265 VSUBS 0.006613f
C319 B.n266 VSUBS 0.006613f
C320 B.n267 VSUBS 0.006613f
C321 B.n268 VSUBS 0.006613f
C322 B.n269 VSUBS 0.006613f
C323 B.n270 VSUBS 0.015622f
C324 B.n271 VSUBS 0.015622f
C325 B.n272 VSUBS 0.016081f
C326 B.n273 VSUBS 0.006613f
C327 B.n274 VSUBS 0.006613f
C328 B.n275 VSUBS 0.006613f
C329 B.n276 VSUBS 0.006613f
C330 B.n277 VSUBS 0.006613f
C331 B.n278 VSUBS 0.006613f
C332 B.n279 VSUBS 0.006613f
C333 B.n280 VSUBS 0.006613f
C334 B.n281 VSUBS 0.006613f
C335 B.n282 VSUBS 0.006613f
C336 B.n283 VSUBS 0.006613f
C337 B.n284 VSUBS 0.006613f
C338 B.n285 VSUBS 0.006613f
C339 B.n286 VSUBS 0.006613f
C340 B.n287 VSUBS 0.006613f
C341 B.n288 VSUBS 0.006613f
C342 B.n289 VSUBS 0.006613f
C343 B.n290 VSUBS 0.006613f
C344 B.n291 VSUBS 0.006613f
C345 B.n292 VSUBS 0.006613f
C346 B.n293 VSUBS 0.006613f
C347 B.n294 VSUBS 0.006613f
C348 B.n295 VSUBS 0.006613f
C349 B.n296 VSUBS 0.006613f
C350 B.n297 VSUBS 0.006613f
C351 B.n298 VSUBS 0.006613f
C352 B.n299 VSUBS 0.006613f
C353 B.n300 VSUBS 0.006613f
C354 B.n301 VSUBS 0.006613f
C355 B.n302 VSUBS 0.006613f
C356 B.n303 VSUBS 0.006613f
C357 B.n304 VSUBS 0.006613f
C358 B.n305 VSUBS 0.006613f
C359 B.n306 VSUBS 0.006613f
C360 B.n307 VSUBS 0.006613f
C361 B.n308 VSUBS 0.006613f
C362 B.n309 VSUBS 0.006613f
C363 B.n310 VSUBS 0.006613f
C364 B.n311 VSUBS 0.006613f
C365 B.n312 VSUBS 0.006613f
C366 B.n313 VSUBS 0.006613f
C367 B.n314 VSUBS 0.006613f
C368 B.n315 VSUBS 0.006613f
C369 B.n316 VSUBS 0.006613f
C370 B.n317 VSUBS 0.006613f
C371 B.n318 VSUBS 0.006613f
C372 B.n319 VSUBS 0.006613f
C373 B.n320 VSUBS 0.006613f
C374 B.n321 VSUBS 0.006613f
C375 B.n322 VSUBS 0.006613f
C376 B.n323 VSUBS 0.006613f
C377 B.n324 VSUBS 0.006613f
C378 B.n325 VSUBS 0.006613f
C379 B.n326 VSUBS 0.006613f
C380 B.n327 VSUBS 0.006613f
C381 B.n328 VSUBS 0.006613f
C382 B.n329 VSUBS 0.006613f
C383 B.n330 VSUBS 0.006613f
C384 B.n331 VSUBS 0.006613f
C385 B.n332 VSUBS 0.006613f
C386 B.n333 VSUBS 0.006613f
C387 B.n334 VSUBS 0.006613f
C388 B.n335 VSUBS 0.006613f
C389 B.n336 VSUBS 0.006613f
C390 B.n337 VSUBS 0.006613f
C391 B.n338 VSUBS 0.006613f
C392 B.n339 VSUBS 0.004571f
C393 B.n340 VSUBS 0.006613f
C394 B.n341 VSUBS 0.006613f
C395 B.n342 VSUBS 0.005349f
C396 B.n343 VSUBS 0.006613f
C397 B.n344 VSUBS 0.006613f
C398 B.n345 VSUBS 0.006613f
C399 B.n346 VSUBS 0.006613f
C400 B.n347 VSUBS 0.006613f
C401 B.n348 VSUBS 0.006613f
C402 B.n349 VSUBS 0.006613f
C403 B.n350 VSUBS 0.006613f
C404 B.n351 VSUBS 0.006613f
C405 B.n352 VSUBS 0.006613f
C406 B.n353 VSUBS 0.006613f
C407 B.n354 VSUBS 0.005349f
C408 B.n355 VSUBS 0.015321f
C409 B.n356 VSUBS 0.004571f
C410 B.n357 VSUBS 0.006613f
C411 B.n358 VSUBS 0.006613f
C412 B.n359 VSUBS 0.006613f
C413 B.n360 VSUBS 0.006613f
C414 B.n361 VSUBS 0.006613f
C415 B.n362 VSUBS 0.006613f
C416 B.n363 VSUBS 0.006613f
C417 B.n364 VSUBS 0.006613f
C418 B.n365 VSUBS 0.006613f
C419 B.n366 VSUBS 0.006613f
C420 B.n367 VSUBS 0.006613f
C421 B.n368 VSUBS 0.006613f
C422 B.n369 VSUBS 0.006613f
C423 B.n370 VSUBS 0.006613f
C424 B.n371 VSUBS 0.006613f
C425 B.n372 VSUBS 0.006613f
C426 B.n373 VSUBS 0.006613f
C427 B.n374 VSUBS 0.006613f
C428 B.n375 VSUBS 0.006613f
C429 B.n376 VSUBS 0.006613f
C430 B.n377 VSUBS 0.006613f
C431 B.n378 VSUBS 0.006613f
C432 B.n379 VSUBS 0.006613f
C433 B.n380 VSUBS 0.006613f
C434 B.n381 VSUBS 0.006613f
C435 B.n382 VSUBS 0.006613f
C436 B.n383 VSUBS 0.006613f
C437 B.n384 VSUBS 0.006613f
C438 B.n385 VSUBS 0.006613f
C439 B.n386 VSUBS 0.006613f
C440 B.n387 VSUBS 0.006613f
C441 B.n388 VSUBS 0.006613f
C442 B.n389 VSUBS 0.006613f
C443 B.n390 VSUBS 0.006613f
C444 B.n391 VSUBS 0.006613f
C445 B.n392 VSUBS 0.006613f
C446 B.n393 VSUBS 0.006613f
C447 B.n394 VSUBS 0.006613f
C448 B.n395 VSUBS 0.006613f
C449 B.n396 VSUBS 0.006613f
C450 B.n397 VSUBS 0.006613f
C451 B.n398 VSUBS 0.006613f
C452 B.n399 VSUBS 0.006613f
C453 B.n400 VSUBS 0.006613f
C454 B.n401 VSUBS 0.006613f
C455 B.n402 VSUBS 0.006613f
C456 B.n403 VSUBS 0.006613f
C457 B.n404 VSUBS 0.006613f
C458 B.n405 VSUBS 0.006613f
C459 B.n406 VSUBS 0.006613f
C460 B.n407 VSUBS 0.006613f
C461 B.n408 VSUBS 0.006613f
C462 B.n409 VSUBS 0.006613f
C463 B.n410 VSUBS 0.006613f
C464 B.n411 VSUBS 0.006613f
C465 B.n412 VSUBS 0.006613f
C466 B.n413 VSUBS 0.006613f
C467 B.n414 VSUBS 0.006613f
C468 B.n415 VSUBS 0.006613f
C469 B.n416 VSUBS 0.006613f
C470 B.n417 VSUBS 0.006613f
C471 B.n418 VSUBS 0.006613f
C472 B.n419 VSUBS 0.006613f
C473 B.n420 VSUBS 0.006613f
C474 B.n421 VSUBS 0.006613f
C475 B.n422 VSUBS 0.006613f
C476 B.n423 VSUBS 0.016081f
C477 B.n424 VSUBS 0.016081f
C478 B.n425 VSUBS 0.015622f
C479 B.n426 VSUBS 0.006613f
C480 B.n427 VSUBS 0.006613f
C481 B.n428 VSUBS 0.006613f
C482 B.n429 VSUBS 0.006613f
C483 B.n430 VSUBS 0.006613f
C484 B.n431 VSUBS 0.006613f
C485 B.n432 VSUBS 0.006613f
C486 B.n433 VSUBS 0.006613f
C487 B.n434 VSUBS 0.006613f
C488 B.n435 VSUBS 0.006613f
C489 B.n436 VSUBS 0.006613f
C490 B.n437 VSUBS 0.006613f
C491 B.n438 VSUBS 0.006613f
C492 B.n439 VSUBS 0.006613f
C493 B.n440 VSUBS 0.006613f
C494 B.n441 VSUBS 0.006613f
C495 B.n442 VSUBS 0.006613f
C496 B.n443 VSUBS 0.006613f
C497 B.n444 VSUBS 0.006613f
C498 B.n445 VSUBS 0.006613f
C499 B.n446 VSUBS 0.006613f
C500 B.n447 VSUBS 0.006613f
C501 B.n448 VSUBS 0.006613f
C502 B.n449 VSUBS 0.006613f
C503 B.n450 VSUBS 0.006613f
C504 B.n451 VSUBS 0.006613f
C505 B.n452 VSUBS 0.006613f
C506 B.n453 VSUBS 0.006613f
C507 B.n454 VSUBS 0.006613f
C508 B.n455 VSUBS 0.006613f
C509 B.n456 VSUBS 0.006613f
C510 B.n457 VSUBS 0.006613f
C511 B.n458 VSUBS 0.006613f
C512 B.n459 VSUBS 0.006613f
C513 B.n460 VSUBS 0.006613f
C514 B.n461 VSUBS 0.006613f
C515 B.n462 VSUBS 0.006613f
C516 B.n463 VSUBS 0.006613f
C517 B.n464 VSUBS 0.006613f
C518 B.n465 VSUBS 0.006613f
C519 B.n466 VSUBS 0.006613f
C520 B.n467 VSUBS 0.006613f
C521 B.n468 VSUBS 0.006613f
C522 B.n469 VSUBS 0.006613f
C523 B.n470 VSUBS 0.006613f
C524 B.n471 VSUBS 0.006613f
C525 B.n472 VSUBS 0.006613f
C526 B.n473 VSUBS 0.006613f
C527 B.n474 VSUBS 0.006613f
C528 B.n475 VSUBS 0.006613f
C529 B.n476 VSUBS 0.006613f
C530 B.n477 VSUBS 0.006613f
C531 B.n478 VSUBS 0.006613f
C532 B.n479 VSUBS 0.006613f
C533 B.n480 VSUBS 0.006613f
C534 B.n481 VSUBS 0.006613f
C535 B.n482 VSUBS 0.006613f
C536 B.n483 VSUBS 0.006613f
C537 B.n484 VSUBS 0.006613f
C538 B.n485 VSUBS 0.006613f
C539 B.n486 VSUBS 0.006613f
C540 B.n487 VSUBS 0.006613f
C541 B.n488 VSUBS 0.006613f
C542 B.n489 VSUBS 0.006613f
C543 B.n490 VSUBS 0.006613f
C544 B.n491 VSUBS 0.006613f
C545 B.n492 VSUBS 0.006613f
C546 B.n493 VSUBS 0.006613f
C547 B.n494 VSUBS 0.006613f
C548 B.n495 VSUBS 0.006613f
C549 B.n496 VSUBS 0.006613f
C550 B.n497 VSUBS 0.006613f
C551 B.n498 VSUBS 0.006613f
C552 B.n499 VSUBS 0.006613f
C553 B.n500 VSUBS 0.006613f
C554 B.n501 VSUBS 0.006613f
C555 B.n502 VSUBS 0.006613f
C556 B.n503 VSUBS 0.006613f
C557 B.n504 VSUBS 0.006613f
C558 B.n505 VSUBS 0.006613f
C559 B.n506 VSUBS 0.006613f
C560 B.n507 VSUBS 0.006613f
C561 B.n508 VSUBS 0.006613f
C562 B.n509 VSUBS 0.006613f
C563 B.n510 VSUBS 0.006613f
C564 B.n511 VSUBS 0.006613f
C565 B.n512 VSUBS 0.006613f
C566 B.n513 VSUBS 0.006613f
C567 B.n514 VSUBS 0.006613f
C568 B.n515 VSUBS 0.006613f
C569 B.n516 VSUBS 0.006613f
C570 B.n517 VSUBS 0.006613f
C571 B.n518 VSUBS 0.006613f
C572 B.n519 VSUBS 0.006613f
C573 B.n520 VSUBS 0.006613f
C574 B.n521 VSUBS 0.006613f
C575 B.n522 VSUBS 0.006613f
C576 B.n523 VSUBS 0.006613f
C577 B.n524 VSUBS 0.006613f
C578 B.n525 VSUBS 0.006613f
C579 B.n526 VSUBS 0.006613f
C580 B.n527 VSUBS 0.006613f
C581 B.n528 VSUBS 0.006613f
C582 B.n529 VSUBS 0.006613f
C583 B.n530 VSUBS 0.006613f
C584 B.n531 VSUBS 0.006613f
C585 B.n532 VSUBS 0.006613f
C586 B.n533 VSUBS 0.006613f
C587 B.n534 VSUBS 0.006613f
C588 B.n535 VSUBS 0.006613f
C589 B.n536 VSUBS 0.006613f
C590 B.n537 VSUBS 0.006613f
C591 B.n538 VSUBS 0.006613f
C592 B.n539 VSUBS 0.006613f
C593 B.n540 VSUBS 0.006613f
C594 B.n541 VSUBS 0.006613f
C595 B.n542 VSUBS 0.006613f
C596 B.n543 VSUBS 0.006613f
C597 B.n544 VSUBS 0.006613f
C598 B.n545 VSUBS 0.006613f
C599 B.n546 VSUBS 0.006613f
C600 B.n547 VSUBS 0.006613f
C601 B.n548 VSUBS 0.006613f
C602 B.n549 VSUBS 0.006613f
C603 B.n550 VSUBS 0.006613f
C604 B.n551 VSUBS 0.006613f
C605 B.n552 VSUBS 0.006613f
C606 B.n553 VSUBS 0.006613f
C607 B.n554 VSUBS 0.006613f
C608 B.n555 VSUBS 0.006613f
C609 B.n556 VSUBS 0.006613f
C610 B.n557 VSUBS 0.006613f
C611 B.n558 VSUBS 0.006613f
C612 B.n559 VSUBS 0.006613f
C613 B.n560 VSUBS 0.006613f
C614 B.n561 VSUBS 0.006613f
C615 B.n562 VSUBS 0.006613f
C616 B.n563 VSUBS 0.015622f
C617 B.n564 VSUBS 0.016081f
C618 B.n565 VSUBS 0.015328f
C619 B.n566 VSUBS 0.006613f
C620 B.n567 VSUBS 0.006613f
C621 B.n568 VSUBS 0.006613f
C622 B.n569 VSUBS 0.006613f
C623 B.n570 VSUBS 0.006613f
C624 B.n571 VSUBS 0.006613f
C625 B.n572 VSUBS 0.006613f
C626 B.n573 VSUBS 0.006613f
C627 B.n574 VSUBS 0.006613f
C628 B.n575 VSUBS 0.006613f
C629 B.n576 VSUBS 0.006613f
C630 B.n577 VSUBS 0.006613f
C631 B.n578 VSUBS 0.006613f
C632 B.n579 VSUBS 0.006613f
C633 B.n580 VSUBS 0.006613f
C634 B.n581 VSUBS 0.006613f
C635 B.n582 VSUBS 0.006613f
C636 B.n583 VSUBS 0.006613f
C637 B.n584 VSUBS 0.006613f
C638 B.n585 VSUBS 0.006613f
C639 B.n586 VSUBS 0.006613f
C640 B.n587 VSUBS 0.006613f
C641 B.n588 VSUBS 0.006613f
C642 B.n589 VSUBS 0.006613f
C643 B.n590 VSUBS 0.006613f
C644 B.n591 VSUBS 0.006613f
C645 B.n592 VSUBS 0.006613f
C646 B.n593 VSUBS 0.006613f
C647 B.n594 VSUBS 0.006613f
C648 B.n595 VSUBS 0.006613f
C649 B.n596 VSUBS 0.006613f
C650 B.n597 VSUBS 0.006613f
C651 B.n598 VSUBS 0.006613f
C652 B.n599 VSUBS 0.006613f
C653 B.n600 VSUBS 0.006613f
C654 B.n601 VSUBS 0.006613f
C655 B.n602 VSUBS 0.006613f
C656 B.n603 VSUBS 0.006613f
C657 B.n604 VSUBS 0.006613f
C658 B.n605 VSUBS 0.006613f
C659 B.n606 VSUBS 0.006613f
C660 B.n607 VSUBS 0.006613f
C661 B.n608 VSUBS 0.006613f
C662 B.n609 VSUBS 0.006613f
C663 B.n610 VSUBS 0.006613f
C664 B.n611 VSUBS 0.006613f
C665 B.n612 VSUBS 0.006613f
C666 B.n613 VSUBS 0.006613f
C667 B.n614 VSUBS 0.006613f
C668 B.n615 VSUBS 0.006613f
C669 B.n616 VSUBS 0.006613f
C670 B.n617 VSUBS 0.006613f
C671 B.n618 VSUBS 0.006613f
C672 B.n619 VSUBS 0.006613f
C673 B.n620 VSUBS 0.006613f
C674 B.n621 VSUBS 0.006613f
C675 B.n622 VSUBS 0.006613f
C676 B.n623 VSUBS 0.006613f
C677 B.n624 VSUBS 0.006613f
C678 B.n625 VSUBS 0.006613f
C679 B.n626 VSUBS 0.006613f
C680 B.n627 VSUBS 0.006613f
C681 B.n628 VSUBS 0.006613f
C682 B.n629 VSUBS 0.006613f
C683 B.n630 VSUBS 0.006613f
C684 B.n631 VSUBS 0.006613f
C685 B.n632 VSUBS 0.004571f
C686 B.n633 VSUBS 0.015321f
C687 B.n634 VSUBS 0.005349f
C688 B.n635 VSUBS 0.006613f
C689 B.n636 VSUBS 0.006613f
C690 B.n637 VSUBS 0.006613f
C691 B.n638 VSUBS 0.006613f
C692 B.n639 VSUBS 0.006613f
C693 B.n640 VSUBS 0.006613f
C694 B.n641 VSUBS 0.006613f
C695 B.n642 VSUBS 0.006613f
C696 B.n643 VSUBS 0.006613f
C697 B.n644 VSUBS 0.006613f
C698 B.n645 VSUBS 0.006613f
C699 B.n646 VSUBS 0.005349f
C700 B.n647 VSUBS 0.006613f
C701 B.n648 VSUBS 0.006613f
C702 B.n649 VSUBS 0.004571f
C703 B.n650 VSUBS 0.006613f
C704 B.n651 VSUBS 0.006613f
C705 B.n652 VSUBS 0.006613f
C706 B.n653 VSUBS 0.006613f
C707 B.n654 VSUBS 0.006613f
C708 B.n655 VSUBS 0.006613f
C709 B.n656 VSUBS 0.006613f
C710 B.n657 VSUBS 0.006613f
C711 B.n658 VSUBS 0.006613f
C712 B.n659 VSUBS 0.006613f
C713 B.n660 VSUBS 0.006613f
C714 B.n661 VSUBS 0.006613f
C715 B.n662 VSUBS 0.006613f
C716 B.n663 VSUBS 0.006613f
C717 B.n664 VSUBS 0.006613f
C718 B.n665 VSUBS 0.006613f
C719 B.n666 VSUBS 0.006613f
C720 B.n667 VSUBS 0.006613f
C721 B.n668 VSUBS 0.006613f
C722 B.n669 VSUBS 0.006613f
C723 B.n670 VSUBS 0.006613f
C724 B.n671 VSUBS 0.006613f
C725 B.n672 VSUBS 0.006613f
C726 B.n673 VSUBS 0.006613f
C727 B.n674 VSUBS 0.006613f
C728 B.n675 VSUBS 0.006613f
C729 B.n676 VSUBS 0.006613f
C730 B.n677 VSUBS 0.006613f
C731 B.n678 VSUBS 0.006613f
C732 B.n679 VSUBS 0.006613f
C733 B.n680 VSUBS 0.006613f
C734 B.n681 VSUBS 0.006613f
C735 B.n682 VSUBS 0.006613f
C736 B.n683 VSUBS 0.006613f
C737 B.n684 VSUBS 0.006613f
C738 B.n685 VSUBS 0.006613f
C739 B.n686 VSUBS 0.006613f
C740 B.n687 VSUBS 0.006613f
C741 B.n688 VSUBS 0.006613f
C742 B.n689 VSUBS 0.006613f
C743 B.n690 VSUBS 0.006613f
C744 B.n691 VSUBS 0.006613f
C745 B.n692 VSUBS 0.006613f
C746 B.n693 VSUBS 0.006613f
C747 B.n694 VSUBS 0.006613f
C748 B.n695 VSUBS 0.006613f
C749 B.n696 VSUBS 0.006613f
C750 B.n697 VSUBS 0.006613f
C751 B.n698 VSUBS 0.006613f
C752 B.n699 VSUBS 0.006613f
C753 B.n700 VSUBS 0.006613f
C754 B.n701 VSUBS 0.006613f
C755 B.n702 VSUBS 0.006613f
C756 B.n703 VSUBS 0.006613f
C757 B.n704 VSUBS 0.006613f
C758 B.n705 VSUBS 0.006613f
C759 B.n706 VSUBS 0.006613f
C760 B.n707 VSUBS 0.006613f
C761 B.n708 VSUBS 0.006613f
C762 B.n709 VSUBS 0.006613f
C763 B.n710 VSUBS 0.006613f
C764 B.n711 VSUBS 0.006613f
C765 B.n712 VSUBS 0.006613f
C766 B.n713 VSUBS 0.006613f
C767 B.n714 VSUBS 0.006613f
C768 B.n715 VSUBS 0.006613f
C769 B.n716 VSUBS 0.016081f
C770 B.n717 VSUBS 0.015622f
C771 B.n718 VSUBS 0.015622f
C772 B.n719 VSUBS 0.006613f
C773 B.n720 VSUBS 0.006613f
C774 B.n721 VSUBS 0.006613f
C775 B.n722 VSUBS 0.006613f
C776 B.n723 VSUBS 0.006613f
C777 B.n724 VSUBS 0.006613f
C778 B.n725 VSUBS 0.006613f
C779 B.n726 VSUBS 0.006613f
C780 B.n727 VSUBS 0.006613f
C781 B.n728 VSUBS 0.006613f
C782 B.n729 VSUBS 0.006613f
C783 B.n730 VSUBS 0.006613f
C784 B.n731 VSUBS 0.006613f
C785 B.n732 VSUBS 0.006613f
C786 B.n733 VSUBS 0.006613f
C787 B.n734 VSUBS 0.006613f
C788 B.n735 VSUBS 0.006613f
C789 B.n736 VSUBS 0.006613f
C790 B.n737 VSUBS 0.006613f
C791 B.n738 VSUBS 0.006613f
C792 B.n739 VSUBS 0.006613f
C793 B.n740 VSUBS 0.006613f
C794 B.n741 VSUBS 0.006613f
C795 B.n742 VSUBS 0.006613f
C796 B.n743 VSUBS 0.006613f
C797 B.n744 VSUBS 0.006613f
C798 B.n745 VSUBS 0.006613f
C799 B.n746 VSUBS 0.006613f
C800 B.n747 VSUBS 0.006613f
C801 B.n748 VSUBS 0.006613f
C802 B.n749 VSUBS 0.006613f
C803 B.n750 VSUBS 0.006613f
C804 B.n751 VSUBS 0.006613f
C805 B.n752 VSUBS 0.006613f
C806 B.n753 VSUBS 0.006613f
C807 B.n754 VSUBS 0.006613f
C808 B.n755 VSUBS 0.006613f
C809 B.n756 VSUBS 0.006613f
C810 B.n757 VSUBS 0.006613f
C811 B.n758 VSUBS 0.006613f
C812 B.n759 VSUBS 0.006613f
C813 B.n760 VSUBS 0.006613f
C814 B.n761 VSUBS 0.006613f
C815 B.n762 VSUBS 0.006613f
C816 B.n763 VSUBS 0.006613f
C817 B.n764 VSUBS 0.006613f
C818 B.n765 VSUBS 0.006613f
C819 B.n766 VSUBS 0.006613f
C820 B.n767 VSUBS 0.006613f
C821 B.n768 VSUBS 0.006613f
C822 B.n769 VSUBS 0.006613f
C823 B.n770 VSUBS 0.006613f
C824 B.n771 VSUBS 0.006613f
C825 B.n772 VSUBS 0.006613f
C826 B.n773 VSUBS 0.006613f
C827 B.n774 VSUBS 0.006613f
C828 B.n775 VSUBS 0.006613f
C829 B.n776 VSUBS 0.006613f
C830 B.n777 VSUBS 0.006613f
C831 B.n778 VSUBS 0.006613f
C832 B.n779 VSUBS 0.006613f
C833 B.n780 VSUBS 0.006613f
C834 B.n781 VSUBS 0.006613f
C835 B.n782 VSUBS 0.006613f
C836 B.n783 VSUBS 0.006613f
C837 B.n784 VSUBS 0.006613f
C838 B.n785 VSUBS 0.006613f
C839 B.n786 VSUBS 0.006613f
C840 B.n787 VSUBS 0.014974f
C841 VDD1.t1 VSUBS 0.29394f
C842 VDD1.t2 VSUBS 0.29394f
C843 VDD1.n0 VSUBS 2.32725f
C844 VDD1.t0 VSUBS 0.29394f
C845 VDD1.t3 VSUBS 0.29394f
C846 VDD1.n1 VSUBS 3.24332f
C847 VTAIL.n0 VSUBS 0.026213f
C848 VTAIL.n1 VSUBS 0.024229f
C849 VTAIL.n2 VSUBS 0.01302f
C850 VTAIL.n3 VSUBS 0.030774f
C851 VTAIL.n4 VSUBS 0.013785f
C852 VTAIL.n5 VSUBS 0.024229f
C853 VTAIL.n6 VSUBS 0.01302f
C854 VTAIL.n7 VSUBS 0.030774f
C855 VTAIL.n8 VSUBS 0.013785f
C856 VTAIL.n9 VSUBS 0.024229f
C857 VTAIL.n10 VSUBS 0.01302f
C858 VTAIL.n11 VSUBS 0.030774f
C859 VTAIL.n12 VSUBS 0.013403f
C860 VTAIL.n13 VSUBS 0.024229f
C861 VTAIL.n14 VSUBS 0.013785f
C862 VTAIL.n15 VSUBS 0.030774f
C863 VTAIL.n16 VSUBS 0.013785f
C864 VTAIL.n17 VSUBS 0.024229f
C865 VTAIL.n18 VSUBS 0.01302f
C866 VTAIL.n19 VSUBS 0.030774f
C867 VTAIL.n20 VSUBS 0.013785f
C868 VTAIL.n21 VSUBS 1.34439f
C869 VTAIL.n22 VSUBS 0.01302f
C870 VTAIL.t2 VSUBS 0.06643f
C871 VTAIL.n23 VSUBS 0.2067f
C872 VTAIL.n24 VSUBS 0.02315f
C873 VTAIL.n25 VSUBS 0.02308f
C874 VTAIL.n26 VSUBS 0.030774f
C875 VTAIL.n27 VSUBS 0.013785f
C876 VTAIL.n28 VSUBS 0.01302f
C877 VTAIL.n29 VSUBS 0.024229f
C878 VTAIL.n30 VSUBS 0.024229f
C879 VTAIL.n31 VSUBS 0.01302f
C880 VTAIL.n32 VSUBS 0.013785f
C881 VTAIL.n33 VSUBS 0.030774f
C882 VTAIL.n34 VSUBS 0.030774f
C883 VTAIL.n35 VSUBS 0.013785f
C884 VTAIL.n36 VSUBS 0.01302f
C885 VTAIL.n37 VSUBS 0.024229f
C886 VTAIL.n38 VSUBS 0.024229f
C887 VTAIL.n39 VSUBS 0.01302f
C888 VTAIL.n40 VSUBS 0.01302f
C889 VTAIL.n41 VSUBS 0.013785f
C890 VTAIL.n42 VSUBS 0.030774f
C891 VTAIL.n43 VSUBS 0.030774f
C892 VTAIL.n44 VSUBS 0.030774f
C893 VTAIL.n45 VSUBS 0.013403f
C894 VTAIL.n46 VSUBS 0.01302f
C895 VTAIL.n47 VSUBS 0.024229f
C896 VTAIL.n48 VSUBS 0.024229f
C897 VTAIL.n49 VSUBS 0.01302f
C898 VTAIL.n50 VSUBS 0.013785f
C899 VTAIL.n51 VSUBS 0.030774f
C900 VTAIL.n52 VSUBS 0.030774f
C901 VTAIL.n53 VSUBS 0.013785f
C902 VTAIL.n54 VSUBS 0.01302f
C903 VTAIL.n55 VSUBS 0.024229f
C904 VTAIL.n56 VSUBS 0.024229f
C905 VTAIL.n57 VSUBS 0.01302f
C906 VTAIL.n58 VSUBS 0.013785f
C907 VTAIL.n59 VSUBS 0.030774f
C908 VTAIL.n60 VSUBS 0.030774f
C909 VTAIL.n61 VSUBS 0.013785f
C910 VTAIL.n62 VSUBS 0.01302f
C911 VTAIL.n63 VSUBS 0.024229f
C912 VTAIL.n64 VSUBS 0.024229f
C913 VTAIL.n65 VSUBS 0.01302f
C914 VTAIL.n66 VSUBS 0.013785f
C915 VTAIL.n67 VSUBS 0.030774f
C916 VTAIL.n68 VSUBS 0.073105f
C917 VTAIL.n69 VSUBS 0.013785f
C918 VTAIL.n70 VSUBS 0.01302f
C919 VTAIL.n71 VSUBS 0.052363f
C920 VTAIL.n72 VSUBS 0.036586f
C921 VTAIL.n73 VSUBS 0.20423f
C922 VTAIL.n74 VSUBS 0.026213f
C923 VTAIL.n75 VSUBS 0.024229f
C924 VTAIL.n76 VSUBS 0.01302f
C925 VTAIL.n77 VSUBS 0.030774f
C926 VTAIL.n78 VSUBS 0.013785f
C927 VTAIL.n79 VSUBS 0.024229f
C928 VTAIL.n80 VSUBS 0.01302f
C929 VTAIL.n81 VSUBS 0.030774f
C930 VTAIL.n82 VSUBS 0.013785f
C931 VTAIL.n83 VSUBS 0.024229f
C932 VTAIL.n84 VSUBS 0.01302f
C933 VTAIL.n85 VSUBS 0.030774f
C934 VTAIL.n86 VSUBS 0.013403f
C935 VTAIL.n87 VSUBS 0.024229f
C936 VTAIL.n88 VSUBS 0.013785f
C937 VTAIL.n89 VSUBS 0.030774f
C938 VTAIL.n90 VSUBS 0.013785f
C939 VTAIL.n91 VSUBS 0.024229f
C940 VTAIL.n92 VSUBS 0.01302f
C941 VTAIL.n93 VSUBS 0.030774f
C942 VTAIL.n94 VSUBS 0.013785f
C943 VTAIL.n95 VSUBS 1.34439f
C944 VTAIL.n96 VSUBS 0.01302f
C945 VTAIL.t6 VSUBS 0.06643f
C946 VTAIL.n97 VSUBS 0.2067f
C947 VTAIL.n98 VSUBS 0.02315f
C948 VTAIL.n99 VSUBS 0.02308f
C949 VTAIL.n100 VSUBS 0.030774f
C950 VTAIL.n101 VSUBS 0.013785f
C951 VTAIL.n102 VSUBS 0.01302f
C952 VTAIL.n103 VSUBS 0.024229f
C953 VTAIL.n104 VSUBS 0.024229f
C954 VTAIL.n105 VSUBS 0.01302f
C955 VTAIL.n106 VSUBS 0.013785f
C956 VTAIL.n107 VSUBS 0.030774f
C957 VTAIL.n108 VSUBS 0.030774f
C958 VTAIL.n109 VSUBS 0.013785f
C959 VTAIL.n110 VSUBS 0.01302f
C960 VTAIL.n111 VSUBS 0.024229f
C961 VTAIL.n112 VSUBS 0.024229f
C962 VTAIL.n113 VSUBS 0.01302f
C963 VTAIL.n114 VSUBS 0.01302f
C964 VTAIL.n115 VSUBS 0.013785f
C965 VTAIL.n116 VSUBS 0.030774f
C966 VTAIL.n117 VSUBS 0.030774f
C967 VTAIL.n118 VSUBS 0.030774f
C968 VTAIL.n119 VSUBS 0.013403f
C969 VTAIL.n120 VSUBS 0.01302f
C970 VTAIL.n121 VSUBS 0.024229f
C971 VTAIL.n122 VSUBS 0.024229f
C972 VTAIL.n123 VSUBS 0.01302f
C973 VTAIL.n124 VSUBS 0.013785f
C974 VTAIL.n125 VSUBS 0.030774f
C975 VTAIL.n126 VSUBS 0.030774f
C976 VTAIL.n127 VSUBS 0.013785f
C977 VTAIL.n128 VSUBS 0.01302f
C978 VTAIL.n129 VSUBS 0.024229f
C979 VTAIL.n130 VSUBS 0.024229f
C980 VTAIL.n131 VSUBS 0.01302f
C981 VTAIL.n132 VSUBS 0.013785f
C982 VTAIL.n133 VSUBS 0.030774f
C983 VTAIL.n134 VSUBS 0.030774f
C984 VTAIL.n135 VSUBS 0.013785f
C985 VTAIL.n136 VSUBS 0.01302f
C986 VTAIL.n137 VSUBS 0.024229f
C987 VTAIL.n138 VSUBS 0.024229f
C988 VTAIL.n139 VSUBS 0.01302f
C989 VTAIL.n140 VSUBS 0.013785f
C990 VTAIL.n141 VSUBS 0.030774f
C991 VTAIL.n142 VSUBS 0.073105f
C992 VTAIL.n143 VSUBS 0.013785f
C993 VTAIL.n144 VSUBS 0.01302f
C994 VTAIL.n145 VSUBS 0.052363f
C995 VTAIL.n146 VSUBS 0.036586f
C996 VTAIL.n147 VSUBS 0.344051f
C997 VTAIL.n148 VSUBS 0.026213f
C998 VTAIL.n149 VSUBS 0.024229f
C999 VTAIL.n150 VSUBS 0.01302f
C1000 VTAIL.n151 VSUBS 0.030774f
C1001 VTAIL.n152 VSUBS 0.013785f
C1002 VTAIL.n153 VSUBS 0.024229f
C1003 VTAIL.n154 VSUBS 0.01302f
C1004 VTAIL.n155 VSUBS 0.030774f
C1005 VTAIL.n156 VSUBS 0.013785f
C1006 VTAIL.n157 VSUBS 0.024229f
C1007 VTAIL.n158 VSUBS 0.01302f
C1008 VTAIL.n159 VSUBS 0.030774f
C1009 VTAIL.n160 VSUBS 0.013403f
C1010 VTAIL.n161 VSUBS 0.024229f
C1011 VTAIL.n162 VSUBS 0.013785f
C1012 VTAIL.n163 VSUBS 0.030774f
C1013 VTAIL.n164 VSUBS 0.013785f
C1014 VTAIL.n165 VSUBS 0.024229f
C1015 VTAIL.n166 VSUBS 0.01302f
C1016 VTAIL.n167 VSUBS 0.030774f
C1017 VTAIL.n168 VSUBS 0.013785f
C1018 VTAIL.n169 VSUBS 1.34439f
C1019 VTAIL.n170 VSUBS 0.01302f
C1020 VTAIL.t7 VSUBS 0.06643f
C1021 VTAIL.n171 VSUBS 0.2067f
C1022 VTAIL.n172 VSUBS 0.02315f
C1023 VTAIL.n173 VSUBS 0.02308f
C1024 VTAIL.n174 VSUBS 0.030774f
C1025 VTAIL.n175 VSUBS 0.013785f
C1026 VTAIL.n176 VSUBS 0.01302f
C1027 VTAIL.n177 VSUBS 0.024229f
C1028 VTAIL.n178 VSUBS 0.024229f
C1029 VTAIL.n179 VSUBS 0.01302f
C1030 VTAIL.n180 VSUBS 0.013785f
C1031 VTAIL.n181 VSUBS 0.030774f
C1032 VTAIL.n182 VSUBS 0.030774f
C1033 VTAIL.n183 VSUBS 0.013785f
C1034 VTAIL.n184 VSUBS 0.01302f
C1035 VTAIL.n185 VSUBS 0.024229f
C1036 VTAIL.n186 VSUBS 0.024229f
C1037 VTAIL.n187 VSUBS 0.01302f
C1038 VTAIL.n188 VSUBS 0.01302f
C1039 VTAIL.n189 VSUBS 0.013785f
C1040 VTAIL.n190 VSUBS 0.030774f
C1041 VTAIL.n191 VSUBS 0.030774f
C1042 VTAIL.n192 VSUBS 0.030774f
C1043 VTAIL.n193 VSUBS 0.013403f
C1044 VTAIL.n194 VSUBS 0.01302f
C1045 VTAIL.n195 VSUBS 0.024229f
C1046 VTAIL.n196 VSUBS 0.024229f
C1047 VTAIL.n197 VSUBS 0.01302f
C1048 VTAIL.n198 VSUBS 0.013785f
C1049 VTAIL.n199 VSUBS 0.030774f
C1050 VTAIL.n200 VSUBS 0.030774f
C1051 VTAIL.n201 VSUBS 0.013785f
C1052 VTAIL.n202 VSUBS 0.01302f
C1053 VTAIL.n203 VSUBS 0.024229f
C1054 VTAIL.n204 VSUBS 0.024229f
C1055 VTAIL.n205 VSUBS 0.01302f
C1056 VTAIL.n206 VSUBS 0.013785f
C1057 VTAIL.n207 VSUBS 0.030774f
C1058 VTAIL.n208 VSUBS 0.030774f
C1059 VTAIL.n209 VSUBS 0.013785f
C1060 VTAIL.n210 VSUBS 0.01302f
C1061 VTAIL.n211 VSUBS 0.024229f
C1062 VTAIL.n212 VSUBS 0.024229f
C1063 VTAIL.n213 VSUBS 0.01302f
C1064 VTAIL.n214 VSUBS 0.013785f
C1065 VTAIL.n215 VSUBS 0.030774f
C1066 VTAIL.n216 VSUBS 0.073105f
C1067 VTAIL.n217 VSUBS 0.013785f
C1068 VTAIL.n218 VSUBS 0.01302f
C1069 VTAIL.n219 VSUBS 0.052363f
C1070 VTAIL.n220 VSUBS 0.036586f
C1071 VTAIL.n221 VSUBS 1.83045f
C1072 VTAIL.n222 VSUBS 0.026213f
C1073 VTAIL.n223 VSUBS 0.024229f
C1074 VTAIL.n224 VSUBS 0.01302f
C1075 VTAIL.n225 VSUBS 0.030774f
C1076 VTAIL.n226 VSUBS 0.013785f
C1077 VTAIL.n227 VSUBS 0.024229f
C1078 VTAIL.n228 VSUBS 0.01302f
C1079 VTAIL.n229 VSUBS 0.030774f
C1080 VTAIL.n230 VSUBS 0.013785f
C1081 VTAIL.n231 VSUBS 0.024229f
C1082 VTAIL.n232 VSUBS 0.01302f
C1083 VTAIL.n233 VSUBS 0.030774f
C1084 VTAIL.n234 VSUBS 0.013403f
C1085 VTAIL.n235 VSUBS 0.024229f
C1086 VTAIL.n236 VSUBS 0.013403f
C1087 VTAIL.n237 VSUBS 0.01302f
C1088 VTAIL.n238 VSUBS 0.030774f
C1089 VTAIL.n239 VSUBS 0.030774f
C1090 VTAIL.n240 VSUBS 0.013785f
C1091 VTAIL.n241 VSUBS 0.024229f
C1092 VTAIL.n242 VSUBS 0.01302f
C1093 VTAIL.n243 VSUBS 0.030774f
C1094 VTAIL.n244 VSUBS 0.013785f
C1095 VTAIL.n245 VSUBS 1.34439f
C1096 VTAIL.n246 VSUBS 0.01302f
C1097 VTAIL.t3 VSUBS 0.06643f
C1098 VTAIL.n247 VSUBS 0.2067f
C1099 VTAIL.n248 VSUBS 0.02315f
C1100 VTAIL.n249 VSUBS 0.02308f
C1101 VTAIL.n250 VSUBS 0.030774f
C1102 VTAIL.n251 VSUBS 0.013785f
C1103 VTAIL.n252 VSUBS 0.01302f
C1104 VTAIL.n253 VSUBS 0.024229f
C1105 VTAIL.n254 VSUBS 0.024229f
C1106 VTAIL.n255 VSUBS 0.01302f
C1107 VTAIL.n256 VSUBS 0.013785f
C1108 VTAIL.n257 VSUBS 0.030774f
C1109 VTAIL.n258 VSUBS 0.030774f
C1110 VTAIL.n259 VSUBS 0.013785f
C1111 VTAIL.n260 VSUBS 0.01302f
C1112 VTAIL.n261 VSUBS 0.024229f
C1113 VTAIL.n262 VSUBS 0.024229f
C1114 VTAIL.n263 VSUBS 0.01302f
C1115 VTAIL.n264 VSUBS 0.013785f
C1116 VTAIL.n265 VSUBS 0.030774f
C1117 VTAIL.n266 VSUBS 0.030774f
C1118 VTAIL.n267 VSUBS 0.013785f
C1119 VTAIL.n268 VSUBS 0.01302f
C1120 VTAIL.n269 VSUBS 0.024229f
C1121 VTAIL.n270 VSUBS 0.024229f
C1122 VTAIL.n271 VSUBS 0.01302f
C1123 VTAIL.n272 VSUBS 0.013785f
C1124 VTAIL.n273 VSUBS 0.030774f
C1125 VTAIL.n274 VSUBS 0.030774f
C1126 VTAIL.n275 VSUBS 0.013785f
C1127 VTAIL.n276 VSUBS 0.01302f
C1128 VTAIL.n277 VSUBS 0.024229f
C1129 VTAIL.n278 VSUBS 0.024229f
C1130 VTAIL.n279 VSUBS 0.01302f
C1131 VTAIL.n280 VSUBS 0.013785f
C1132 VTAIL.n281 VSUBS 0.030774f
C1133 VTAIL.n282 VSUBS 0.030774f
C1134 VTAIL.n283 VSUBS 0.013785f
C1135 VTAIL.n284 VSUBS 0.01302f
C1136 VTAIL.n285 VSUBS 0.024229f
C1137 VTAIL.n286 VSUBS 0.024229f
C1138 VTAIL.n287 VSUBS 0.01302f
C1139 VTAIL.n288 VSUBS 0.013785f
C1140 VTAIL.n289 VSUBS 0.030774f
C1141 VTAIL.n290 VSUBS 0.073105f
C1142 VTAIL.n291 VSUBS 0.013785f
C1143 VTAIL.n292 VSUBS 0.01302f
C1144 VTAIL.n293 VSUBS 0.052363f
C1145 VTAIL.n294 VSUBS 0.036586f
C1146 VTAIL.n295 VSUBS 1.83045f
C1147 VTAIL.n296 VSUBS 0.026213f
C1148 VTAIL.n297 VSUBS 0.024229f
C1149 VTAIL.n298 VSUBS 0.01302f
C1150 VTAIL.n299 VSUBS 0.030774f
C1151 VTAIL.n300 VSUBS 0.013785f
C1152 VTAIL.n301 VSUBS 0.024229f
C1153 VTAIL.n302 VSUBS 0.01302f
C1154 VTAIL.n303 VSUBS 0.030774f
C1155 VTAIL.n304 VSUBS 0.013785f
C1156 VTAIL.n305 VSUBS 0.024229f
C1157 VTAIL.n306 VSUBS 0.01302f
C1158 VTAIL.n307 VSUBS 0.030774f
C1159 VTAIL.n308 VSUBS 0.013403f
C1160 VTAIL.n309 VSUBS 0.024229f
C1161 VTAIL.n310 VSUBS 0.013403f
C1162 VTAIL.n311 VSUBS 0.01302f
C1163 VTAIL.n312 VSUBS 0.030774f
C1164 VTAIL.n313 VSUBS 0.030774f
C1165 VTAIL.n314 VSUBS 0.013785f
C1166 VTAIL.n315 VSUBS 0.024229f
C1167 VTAIL.n316 VSUBS 0.01302f
C1168 VTAIL.n317 VSUBS 0.030774f
C1169 VTAIL.n318 VSUBS 0.013785f
C1170 VTAIL.n319 VSUBS 1.34439f
C1171 VTAIL.n320 VSUBS 0.01302f
C1172 VTAIL.t0 VSUBS 0.06643f
C1173 VTAIL.n321 VSUBS 0.2067f
C1174 VTAIL.n322 VSUBS 0.02315f
C1175 VTAIL.n323 VSUBS 0.02308f
C1176 VTAIL.n324 VSUBS 0.030774f
C1177 VTAIL.n325 VSUBS 0.013785f
C1178 VTAIL.n326 VSUBS 0.01302f
C1179 VTAIL.n327 VSUBS 0.024229f
C1180 VTAIL.n328 VSUBS 0.024229f
C1181 VTAIL.n329 VSUBS 0.01302f
C1182 VTAIL.n330 VSUBS 0.013785f
C1183 VTAIL.n331 VSUBS 0.030774f
C1184 VTAIL.n332 VSUBS 0.030774f
C1185 VTAIL.n333 VSUBS 0.013785f
C1186 VTAIL.n334 VSUBS 0.01302f
C1187 VTAIL.n335 VSUBS 0.024229f
C1188 VTAIL.n336 VSUBS 0.024229f
C1189 VTAIL.n337 VSUBS 0.01302f
C1190 VTAIL.n338 VSUBS 0.013785f
C1191 VTAIL.n339 VSUBS 0.030774f
C1192 VTAIL.n340 VSUBS 0.030774f
C1193 VTAIL.n341 VSUBS 0.013785f
C1194 VTAIL.n342 VSUBS 0.01302f
C1195 VTAIL.n343 VSUBS 0.024229f
C1196 VTAIL.n344 VSUBS 0.024229f
C1197 VTAIL.n345 VSUBS 0.01302f
C1198 VTAIL.n346 VSUBS 0.013785f
C1199 VTAIL.n347 VSUBS 0.030774f
C1200 VTAIL.n348 VSUBS 0.030774f
C1201 VTAIL.n349 VSUBS 0.013785f
C1202 VTAIL.n350 VSUBS 0.01302f
C1203 VTAIL.n351 VSUBS 0.024229f
C1204 VTAIL.n352 VSUBS 0.024229f
C1205 VTAIL.n353 VSUBS 0.01302f
C1206 VTAIL.n354 VSUBS 0.013785f
C1207 VTAIL.n355 VSUBS 0.030774f
C1208 VTAIL.n356 VSUBS 0.030774f
C1209 VTAIL.n357 VSUBS 0.013785f
C1210 VTAIL.n358 VSUBS 0.01302f
C1211 VTAIL.n359 VSUBS 0.024229f
C1212 VTAIL.n360 VSUBS 0.024229f
C1213 VTAIL.n361 VSUBS 0.01302f
C1214 VTAIL.n362 VSUBS 0.013785f
C1215 VTAIL.n363 VSUBS 0.030774f
C1216 VTAIL.n364 VSUBS 0.073105f
C1217 VTAIL.n365 VSUBS 0.013785f
C1218 VTAIL.n366 VSUBS 0.01302f
C1219 VTAIL.n367 VSUBS 0.052363f
C1220 VTAIL.n368 VSUBS 0.036586f
C1221 VTAIL.n369 VSUBS 0.344051f
C1222 VTAIL.n370 VSUBS 0.026213f
C1223 VTAIL.n371 VSUBS 0.024229f
C1224 VTAIL.n372 VSUBS 0.01302f
C1225 VTAIL.n373 VSUBS 0.030774f
C1226 VTAIL.n374 VSUBS 0.013785f
C1227 VTAIL.n375 VSUBS 0.024229f
C1228 VTAIL.n376 VSUBS 0.01302f
C1229 VTAIL.n377 VSUBS 0.030774f
C1230 VTAIL.n378 VSUBS 0.013785f
C1231 VTAIL.n379 VSUBS 0.024229f
C1232 VTAIL.n380 VSUBS 0.01302f
C1233 VTAIL.n381 VSUBS 0.030774f
C1234 VTAIL.n382 VSUBS 0.013403f
C1235 VTAIL.n383 VSUBS 0.024229f
C1236 VTAIL.n384 VSUBS 0.013403f
C1237 VTAIL.n385 VSUBS 0.01302f
C1238 VTAIL.n386 VSUBS 0.030774f
C1239 VTAIL.n387 VSUBS 0.030774f
C1240 VTAIL.n388 VSUBS 0.013785f
C1241 VTAIL.n389 VSUBS 0.024229f
C1242 VTAIL.n390 VSUBS 0.01302f
C1243 VTAIL.n391 VSUBS 0.030774f
C1244 VTAIL.n392 VSUBS 0.013785f
C1245 VTAIL.n393 VSUBS 1.34439f
C1246 VTAIL.n394 VSUBS 0.01302f
C1247 VTAIL.t5 VSUBS 0.06643f
C1248 VTAIL.n395 VSUBS 0.2067f
C1249 VTAIL.n396 VSUBS 0.02315f
C1250 VTAIL.n397 VSUBS 0.02308f
C1251 VTAIL.n398 VSUBS 0.030774f
C1252 VTAIL.n399 VSUBS 0.013785f
C1253 VTAIL.n400 VSUBS 0.01302f
C1254 VTAIL.n401 VSUBS 0.024229f
C1255 VTAIL.n402 VSUBS 0.024229f
C1256 VTAIL.n403 VSUBS 0.01302f
C1257 VTAIL.n404 VSUBS 0.013785f
C1258 VTAIL.n405 VSUBS 0.030774f
C1259 VTAIL.n406 VSUBS 0.030774f
C1260 VTAIL.n407 VSUBS 0.013785f
C1261 VTAIL.n408 VSUBS 0.01302f
C1262 VTAIL.n409 VSUBS 0.024229f
C1263 VTAIL.n410 VSUBS 0.024229f
C1264 VTAIL.n411 VSUBS 0.01302f
C1265 VTAIL.n412 VSUBS 0.013785f
C1266 VTAIL.n413 VSUBS 0.030774f
C1267 VTAIL.n414 VSUBS 0.030774f
C1268 VTAIL.n415 VSUBS 0.013785f
C1269 VTAIL.n416 VSUBS 0.01302f
C1270 VTAIL.n417 VSUBS 0.024229f
C1271 VTAIL.n418 VSUBS 0.024229f
C1272 VTAIL.n419 VSUBS 0.01302f
C1273 VTAIL.n420 VSUBS 0.013785f
C1274 VTAIL.n421 VSUBS 0.030774f
C1275 VTAIL.n422 VSUBS 0.030774f
C1276 VTAIL.n423 VSUBS 0.013785f
C1277 VTAIL.n424 VSUBS 0.01302f
C1278 VTAIL.n425 VSUBS 0.024229f
C1279 VTAIL.n426 VSUBS 0.024229f
C1280 VTAIL.n427 VSUBS 0.01302f
C1281 VTAIL.n428 VSUBS 0.013785f
C1282 VTAIL.n429 VSUBS 0.030774f
C1283 VTAIL.n430 VSUBS 0.030774f
C1284 VTAIL.n431 VSUBS 0.013785f
C1285 VTAIL.n432 VSUBS 0.01302f
C1286 VTAIL.n433 VSUBS 0.024229f
C1287 VTAIL.n434 VSUBS 0.024229f
C1288 VTAIL.n435 VSUBS 0.01302f
C1289 VTAIL.n436 VSUBS 0.013785f
C1290 VTAIL.n437 VSUBS 0.030774f
C1291 VTAIL.n438 VSUBS 0.073105f
C1292 VTAIL.n439 VSUBS 0.013785f
C1293 VTAIL.n440 VSUBS 0.01302f
C1294 VTAIL.n441 VSUBS 0.052363f
C1295 VTAIL.n442 VSUBS 0.036586f
C1296 VTAIL.n443 VSUBS 0.344051f
C1297 VTAIL.n444 VSUBS 0.026213f
C1298 VTAIL.n445 VSUBS 0.024229f
C1299 VTAIL.n446 VSUBS 0.01302f
C1300 VTAIL.n447 VSUBS 0.030774f
C1301 VTAIL.n448 VSUBS 0.013785f
C1302 VTAIL.n449 VSUBS 0.024229f
C1303 VTAIL.n450 VSUBS 0.01302f
C1304 VTAIL.n451 VSUBS 0.030774f
C1305 VTAIL.n452 VSUBS 0.013785f
C1306 VTAIL.n453 VSUBS 0.024229f
C1307 VTAIL.n454 VSUBS 0.01302f
C1308 VTAIL.n455 VSUBS 0.030774f
C1309 VTAIL.n456 VSUBS 0.013403f
C1310 VTAIL.n457 VSUBS 0.024229f
C1311 VTAIL.n458 VSUBS 0.013403f
C1312 VTAIL.n459 VSUBS 0.01302f
C1313 VTAIL.n460 VSUBS 0.030774f
C1314 VTAIL.n461 VSUBS 0.030774f
C1315 VTAIL.n462 VSUBS 0.013785f
C1316 VTAIL.n463 VSUBS 0.024229f
C1317 VTAIL.n464 VSUBS 0.01302f
C1318 VTAIL.n465 VSUBS 0.030774f
C1319 VTAIL.n466 VSUBS 0.013785f
C1320 VTAIL.n467 VSUBS 1.34439f
C1321 VTAIL.n468 VSUBS 0.01302f
C1322 VTAIL.t4 VSUBS 0.06643f
C1323 VTAIL.n469 VSUBS 0.2067f
C1324 VTAIL.n470 VSUBS 0.02315f
C1325 VTAIL.n471 VSUBS 0.02308f
C1326 VTAIL.n472 VSUBS 0.030774f
C1327 VTAIL.n473 VSUBS 0.013785f
C1328 VTAIL.n474 VSUBS 0.01302f
C1329 VTAIL.n475 VSUBS 0.024229f
C1330 VTAIL.n476 VSUBS 0.024229f
C1331 VTAIL.n477 VSUBS 0.01302f
C1332 VTAIL.n478 VSUBS 0.013785f
C1333 VTAIL.n479 VSUBS 0.030774f
C1334 VTAIL.n480 VSUBS 0.030774f
C1335 VTAIL.n481 VSUBS 0.013785f
C1336 VTAIL.n482 VSUBS 0.01302f
C1337 VTAIL.n483 VSUBS 0.024229f
C1338 VTAIL.n484 VSUBS 0.024229f
C1339 VTAIL.n485 VSUBS 0.01302f
C1340 VTAIL.n486 VSUBS 0.013785f
C1341 VTAIL.n487 VSUBS 0.030774f
C1342 VTAIL.n488 VSUBS 0.030774f
C1343 VTAIL.n489 VSUBS 0.013785f
C1344 VTAIL.n490 VSUBS 0.01302f
C1345 VTAIL.n491 VSUBS 0.024229f
C1346 VTAIL.n492 VSUBS 0.024229f
C1347 VTAIL.n493 VSUBS 0.01302f
C1348 VTAIL.n494 VSUBS 0.013785f
C1349 VTAIL.n495 VSUBS 0.030774f
C1350 VTAIL.n496 VSUBS 0.030774f
C1351 VTAIL.n497 VSUBS 0.013785f
C1352 VTAIL.n498 VSUBS 0.01302f
C1353 VTAIL.n499 VSUBS 0.024229f
C1354 VTAIL.n500 VSUBS 0.024229f
C1355 VTAIL.n501 VSUBS 0.01302f
C1356 VTAIL.n502 VSUBS 0.013785f
C1357 VTAIL.n503 VSUBS 0.030774f
C1358 VTAIL.n504 VSUBS 0.030774f
C1359 VTAIL.n505 VSUBS 0.013785f
C1360 VTAIL.n506 VSUBS 0.01302f
C1361 VTAIL.n507 VSUBS 0.024229f
C1362 VTAIL.n508 VSUBS 0.024229f
C1363 VTAIL.n509 VSUBS 0.01302f
C1364 VTAIL.n510 VSUBS 0.013785f
C1365 VTAIL.n511 VSUBS 0.030774f
C1366 VTAIL.n512 VSUBS 0.073105f
C1367 VTAIL.n513 VSUBS 0.013785f
C1368 VTAIL.n514 VSUBS 0.01302f
C1369 VTAIL.n515 VSUBS 0.052363f
C1370 VTAIL.n516 VSUBS 0.036586f
C1371 VTAIL.n517 VSUBS 1.83045f
C1372 VTAIL.n518 VSUBS 0.026213f
C1373 VTAIL.n519 VSUBS 0.024229f
C1374 VTAIL.n520 VSUBS 0.01302f
C1375 VTAIL.n521 VSUBS 0.030774f
C1376 VTAIL.n522 VSUBS 0.013785f
C1377 VTAIL.n523 VSUBS 0.024229f
C1378 VTAIL.n524 VSUBS 0.01302f
C1379 VTAIL.n525 VSUBS 0.030774f
C1380 VTAIL.n526 VSUBS 0.013785f
C1381 VTAIL.n527 VSUBS 0.024229f
C1382 VTAIL.n528 VSUBS 0.01302f
C1383 VTAIL.n529 VSUBS 0.030774f
C1384 VTAIL.n530 VSUBS 0.013403f
C1385 VTAIL.n531 VSUBS 0.024229f
C1386 VTAIL.n532 VSUBS 0.013785f
C1387 VTAIL.n533 VSUBS 0.030774f
C1388 VTAIL.n534 VSUBS 0.013785f
C1389 VTAIL.n535 VSUBS 0.024229f
C1390 VTAIL.n536 VSUBS 0.01302f
C1391 VTAIL.n537 VSUBS 0.030774f
C1392 VTAIL.n538 VSUBS 0.013785f
C1393 VTAIL.n539 VSUBS 1.34439f
C1394 VTAIL.n540 VSUBS 0.01302f
C1395 VTAIL.t1 VSUBS 0.06643f
C1396 VTAIL.n541 VSUBS 0.2067f
C1397 VTAIL.n542 VSUBS 0.02315f
C1398 VTAIL.n543 VSUBS 0.02308f
C1399 VTAIL.n544 VSUBS 0.030774f
C1400 VTAIL.n545 VSUBS 0.013785f
C1401 VTAIL.n546 VSUBS 0.01302f
C1402 VTAIL.n547 VSUBS 0.024229f
C1403 VTAIL.n548 VSUBS 0.024229f
C1404 VTAIL.n549 VSUBS 0.01302f
C1405 VTAIL.n550 VSUBS 0.013785f
C1406 VTAIL.n551 VSUBS 0.030774f
C1407 VTAIL.n552 VSUBS 0.030774f
C1408 VTAIL.n553 VSUBS 0.013785f
C1409 VTAIL.n554 VSUBS 0.01302f
C1410 VTAIL.n555 VSUBS 0.024229f
C1411 VTAIL.n556 VSUBS 0.024229f
C1412 VTAIL.n557 VSUBS 0.01302f
C1413 VTAIL.n558 VSUBS 0.01302f
C1414 VTAIL.n559 VSUBS 0.013785f
C1415 VTAIL.n560 VSUBS 0.030774f
C1416 VTAIL.n561 VSUBS 0.030774f
C1417 VTAIL.n562 VSUBS 0.030774f
C1418 VTAIL.n563 VSUBS 0.013403f
C1419 VTAIL.n564 VSUBS 0.01302f
C1420 VTAIL.n565 VSUBS 0.024229f
C1421 VTAIL.n566 VSUBS 0.024229f
C1422 VTAIL.n567 VSUBS 0.01302f
C1423 VTAIL.n568 VSUBS 0.013785f
C1424 VTAIL.n569 VSUBS 0.030774f
C1425 VTAIL.n570 VSUBS 0.030774f
C1426 VTAIL.n571 VSUBS 0.013785f
C1427 VTAIL.n572 VSUBS 0.01302f
C1428 VTAIL.n573 VSUBS 0.024229f
C1429 VTAIL.n574 VSUBS 0.024229f
C1430 VTAIL.n575 VSUBS 0.01302f
C1431 VTAIL.n576 VSUBS 0.013785f
C1432 VTAIL.n577 VSUBS 0.030774f
C1433 VTAIL.n578 VSUBS 0.030774f
C1434 VTAIL.n579 VSUBS 0.013785f
C1435 VTAIL.n580 VSUBS 0.01302f
C1436 VTAIL.n581 VSUBS 0.024229f
C1437 VTAIL.n582 VSUBS 0.024229f
C1438 VTAIL.n583 VSUBS 0.01302f
C1439 VTAIL.n584 VSUBS 0.013785f
C1440 VTAIL.n585 VSUBS 0.030774f
C1441 VTAIL.n586 VSUBS 0.073105f
C1442 VTAIL.n587 VSUBS 0.013785f
C1443 VTAIL.n588 VSUBS 0.01302f
C1444 VTAIL.n589 VSUBS 0.052363f
C1445 VTAIL.n590 VSUBS 0.036586f
C1446 VTAIL.n591 VSUBS 1.68154f
C1447 VP.n0 VSUBS 0.053446f
C1448 VP.t0 VSUBS 4.13603f
C1449 VP.n1 VSUBS 0.052956f
C1450 VP.n2 VSUBS 0.028413f
C1451 VP.n3 VSUBS 0.052956f
C1452 VP.t1 VSUBS 4.60616f
C1453 VP.t2 VSUBS 4.626f
C1454 VP.n4 VSUBS 4.7045f
C1455 VP.n5 VSUBS 1.8247f
C1456 VP.t3 VSUBS 4.13603f
C1457 VP.n6 VSUBS 1.5624f
C1458 VP.n7 VSUBS 0.047464f
C1459 VP.n8 VSUBS 0.053446f
C1460 VP.n9 VSUBS 0.028413f
C1461 VP.n10 VSUBS 0.028413f
C1462 VP.n11 VSUBS 0.052956f
C1463 VP.n12 VSUBS 0.041479f
C1464 VP.n13 VSUBS 0.041479f
C1465 VP.n14 VSUBS 0.028413f
C1466 VP.n15 VSUBS 0.028413f
C1467 VP.n16 VSUBS 0.028413f
C1468 VP.n17 VSUBS 0.052956f
C1469 VP.n18 VSUBS 0.047464f
C1470 VP.n19 VSUBS 1.5624f
C1471 VP.n20 VSUBS 0.091781f
.ends

