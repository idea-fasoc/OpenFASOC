* NGSPICE file created from diff_pair_sample_0149.ext - technology: sky130A

.subckt diff_pair_sample_0149 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=2.99
X1 VDD1.t8 VP.t1 VTAIL.t18 B.t2 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X2 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X3 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X4 VDD1.t7 VP.t2 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X5 VTAIL.t14 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X6 VTAIL.t1 VN.t2 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X7 VDD2.t6 VN.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=2.99
X8 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=2.99
X9 VDD1.t5 VP.t4 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=2.99
X10 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=2.99
X11 VDD2.t5 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=2.99
X12 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=2.99
X13 VDD2.t3 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=2.99
X14 VTAIL.t17 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X15 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X16 VDD1.t3 VP.t6 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=2.99
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=2.99
X18 VTAIL.t3 VN.t8 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=2.99
X20 VDD1.t2 VP.t7 VTAIL.t19 B.t4 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=2.99
X21 VTAIL.t15 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X22 VDD2.t0 VN.t9 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
X23 VTAIL.t13 VP.t9 VDD1.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=2.99
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t4 92.6706
R47 VP.n61 VP.n60 70.9831
R48 VP.n104 VP.n0 70.9831
R49 VP.n59 VP.n14 70.9831
R50 VP.n26 VP.n25 70.1652
R51 VP.n61 VP.t0 61.0162
R52 VP.n69 VP.t3 61.0162
R53 VP.n82 VP.t2 61.0162
R54 VP.n94 VP.t8 61.0162
R55 VP.n0 VP.t6 61.0162
R56 VP.n14 VP.t7 61.0162
R57 VP.n49 VP.t5 61.0162
R58 VP.n37 VP.t1 61.0162
R59 VP.n25 VP.t9 61.0162
R60 VP.n67 VP.n12 56.5193
R61 VP.n100 VP.n2 56.5193
R62 VP.n55 VP.n16 56.5193
R63 VP.n60 VP.n59 51.9842
R64 VP.n76 VP.n8 49.2348
R65 VP.n88 VP.n87 49.2348
R66 VP.n43 VP.n42 49.2348
R67 VP.n31 VP.n22 49.2348
R68 VP.n76 VP.n75 31.752
R69 VP.n89 VP.n88 31.752
R70 VP.n44 VP.n43 31.752
R71 VP.n31 VP.n30 31.752
R72 VP.n63 VP.n62 24.4675
R73 VP.n63 VP.n12 24.4675
R74 VP.n68 VP.n67 24.4675
R75 VP.n70 VP.n68 24.4675
R76 VP.n74 VP.n10 24.4675
R77 VP.n75 VP.n74 24.4675
R78 VP.n80 VP.n8 24.4675
R79 VP.n81 VP.n80 24.4675
R80 VP.n83 VP.n6 24.4675
R81 VP.n87 VP.n6 24.4675
R82 VP.n89 VP.n4 24.4675
R83 VP.n93 VP.n4 24.4675
R84 VP.n96 VP.n95 24.4675
R85 VP.n96 VP.n2 24.4675
R86 VP.n101 VP.n100 24.4675
R87 VP.n102 VP.n101 24.4675
R88 VP.n56 VP.n55 24.4675
R89 VP.n57 VP.n56 24.4675
R90 VP.n44 VP.n18 24.4675
R91 VP.n48 VP.n18 24.4675
R92 VP.n51 VP.n50 24.4675
R93 VP.n51 VP.n16 24.4675
R94 VP.n35 VP.n22 24.4675
R95 VP.n36 VP.n35 24.4675
R96 VP.n38 VP.n20 24.4675
R97 VP.n42 VP.n20 24.4675
R98 VP.n29 VP.n24 24.4675
R99 VP.n30 VP.n29 24.4675
R100 VP.n70 VP.n69 21.0421
R101 VP.n95 VP.n94 21.0421
R102 VP.n50 VP.n49 21.0421
R103 VP.n62 VP.n61 19.0848
R104 VP.n102 VP.n0 19.0848
R105 VP.n57 VP.n14 19.0848
R106 VP.n82 VP.n81 12.234
R107 VP.n83 VP.n82 12.234
R108 VP.n37 VP.n36 12.234
R109 VP.n38 VP.n37 12.234
R110 VP.n27 VP.n26 5.61939
R111 VP.n69 VP.n10 3.42588
R112 VP.n94 VP.n93 3.42588
R113 VP.n49 VP.n48 3.42588
R114 VP.n25 VP.n24 3.42588
R115 VP.n59 VP.n58 0.354971
R116 VP.n60 VP.n13 0.354971
R117 VP.n104 VP.n103 0.354971
R118 VP VP.n104 0.26696
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VTAIL.n11 VTAIL.t7 52.7493
R164 VTAIL.n17 VTAIL.t4 52.7491
R165 VTAIL.n2 VTAIL.t11 52.7491
R166 VTAIL.n16 VTAIL.t19 52.7491
R167 VTAIL.n15 VTAIL.n14 50.1337
R168 VTAIL.n13 VTAIL.n12 50.1337
R169 VTAIL.n10 VTAIL.n9 50.1337
R170 VTAIL.n8 VTAIL.n7 50.1337
R171 VTAIL.n19 VTAIL.n18 50.1335
R172 VTAIL.n1 VTAIL.n0 50.1335
R173 VTAIL.n4 VTAIL.n3 50.1335
R174 VTAIL.n6 VTAIL.n5 50.1335
R175 VTAIL.n8 VTAIL.n6 24.6169
R176 VTAIL.n17 VTAIL.n16 21.7548
R177 VTAIL.n10 VTAIL.n8 2.86257
R178 VTAIL.n11 VTAIL.n10 2.86257
R179 VTAIL.n15 VTAIL.n13 2.86257
R180 VTAIL.n16 VTAIL.n15 2.86257
R181 VTAIL.n6 VTAIL.n4 2.86257
R182 VTAIL.n4 VTAIL.n2 2.86257
R183 VTAIL.n19 VTAIL.n17 2.86257
R184 VTAIL.n18 VTAIL.t2 2.61609
R185 VTAIL.n18 VTAIL.t3 2.61609
R186 VTAIL.n0 VTAIL.t9 2.61609
R187 VTAIL.n0 VTAIL.t8 2.61609
R188 VTAIL.n3 VTAIL.t16 2.61609
R189 VTAIL.n3 VTAIL.t15 2.61609
R190 VTAIL.n5 VTAIL.t10 2.61609
R191 VTAIL.n5 VTAIL.t14 2.61609
R192 VTAIL.n14 VTAIL.t18 2.61609
R193 VTAIL.n14 VTAIL.t17 2.61609
R194 VTAIL.n12 VTAIL.t12 2.61609
R195 VTAIL.n12 VTAIL.t13 2.61609
R196 VTAIL.n9 VTAIL.t6 2.61609
R197 VTAIL.n9 VTAIL.t1 2.61609
R198 VTAIL.n7 VTAIL.t0 2.61609
R199 VTAIL.n7 VTAIL.t5 2.61609
R200 VTAIL VTAIL.n1 2.20524
R201 VTAIL.n13 VTAIL.n11 1.90136
R202 VTAIL.n2 VTAIL.n1 1.90136
R203 VTAIL VTAIL.n19 0.657828
R204 VDD1.n1 VDD1.t5 72.2901
R205 VDD1.n3 VDD1.t9 72.29
R206 VDD1.n5 VDD1.n4 68.9035
R207 VDD1.n1 VDD1.n0 66.8125
R208 VDD1.n7 VDD1.n6 66.8123
R209 VDD1.n3 VDD1.n2 66.8123
R210 VDD1.n7 VDD1.n5 45.85
R211 VDD1.n6 VDD1.t4 2.61609
R212 VDD1.n6 VDD1.t2 2.61609
R213 VDD1.n0 VDD1.t0 2.61609
R214 VDD1.n0 VDD1.t8 2.61609
R215 VDD1.n4 VDD1.t1 2.61609
R216 VDD1.n4 VDD1.t3 2.61609
R217 VDD1.n2 VDD1.t6 2.61609
R218 VDD1.n2 VDD1.t7 2.61609
R219 VDD1 VDD1.n7 2.08886
R220 VDD1 VDD1.n1 0.774207
R221 VDD1.n5 VDD1.n3 0.660671
R222 B.n747 B.n160 585
R223 B.n160 B.n121 585
R224 B.n749 B.n748 585
R225 B.n751 B.n159 585
R226 B.n754 B.n753 585
R227 B.n755 B.n158 585
R228 B.n757 B.n756 585
R229 B.n759 B.n157 585
R230 B.n762 B.n761 585
R231 B.n763 B.n156 585
R232 B.n765 B.n764 585
R233 B.n767 B.n155 585
R234 B.n770 B.n769 585
R235 B.n771 B.n154 585
R236 B.n773 B.n772 585
R237 B.n775 B.n153 585
R238 B.n778 B.n777 585
R239 B.n779 B.n152 585
R240 B.n781 B.n780 585
R241 B.n783 B.n151 585
R242 B.n786 B.n785 585
R243 B.n787 B.n150 585
R244 B.n789 B.n788 585
R245 B.n791 B.n149 585
R246 B.n794 B.n793 585
R247 B.n795 B.n148 585
R248 B.n797 B.n796 585
R249 B.n799 B.n147 585
R250 B.n801 B.n800 585
R251 B.n803 B.n802 585
R252 B.n806 B.n805 585
R253 B.n807 B.n142 585
R254 B.n809 B.n808 585
R255 B.n811 B.n141 585
R256 B.n814 B.n813 585
R257 B.n815 B.n140 585
R258 B.n817 B.n816 585
R259 B.n819 B.n139 585
R260 B.n822 B.n821 585
R261 B.n824 B.n136 585
R262 B.n826 B.n825 585
R263 B.n828 B.n135 585
R264 B.n831 B.n830 585
R265 B.n832 B.n134 585
R266 B.n834 B.n833 585
R267 B.n836 B.n133 585
R268 B.n839 B.n838 585
R269 B.n840 B.n132 585
R270 B.n842 B.n841 585
R271 B.n844 B.n131 585
R272 B.n847 B.n846 585
R273 B.n848 B.n130 585
R274 B.n850 B.n849 585
R275 B.n852 B.n129 585
R276 B.n855 B.n854 585
R277 B.n856 B.n128 585
R278 B.n858 B.n857 585
R279 B.n860 B.n127 585
R280 B.n863 B.n862 585
R281 B.n864 B.n126 585
R282 B.n866 B.n865 585
R283 B.n868 B.n125 585
R284 B.n871 B.n870 585
R285 B.n872 B.n124 585
R286 B.n874 B.n873 585
R287 B.n876 B.n123 585
R288 B.n879 B.n878 585
R289 B.n880 B.n122 585
R290 B.n746 B.n120 585
R291 B.n883 B.n120 585
R292 B.n745 B.n119 585
R293 B.n884 B.n119 585
R294 B.n744 B.n118 585
R295 B.n885 B.n118 585
R296 B.n743 B.n742 585
R297 B.n742 B.n114 585
R298 B.n741 B.n113 585
R299 B.n891 B.n113 585
R300 B.n740 B.n112 585
R301 B.n892 B.n112 585
R302 B.n739 B.n111 585
R303 B.n893 B.n111 585
R304 B.n738 B.n737 585
R305 B.n737 B.n110 585
R306 B.n736 B.n106 585
R307 B.n899 B.n106 585
R308 B.n735 B.n105 585
R309 B.n900 B.n105 585
R310 B.n734 B.n104 585
R311 B.n901 B.n104 585
R312 B.n733 B.n732 585
R313 B.n732 B.n100 585
R314 B.n731 B.n99 585
R315 B.n907 B.n99 585
R316 B.n730 B.n98 585
R317 B.n908 B.n98 585
R318 B.n729 B.n97 585
R319 B.n909 B.n97 585
R320 B.n728 B.n727 585
R321 B.n727 B.n93 585
R322 B.n726 B.n92 585
R323 B.n915 B.n92 585
R324 B.n725 B.n91 585
R325 B.n916 B.n91 585
R326 B.n724 B.n90 585
R327 B.n917 B.n90 585
R328 B.n723 B.n722 585
R329 B.n722 B.n86 585
R330 B.n721 B.n85 585
R331 B.n923 B.n85 585
R332 B.n720 B.n84 585
R333 B.n924 B.n84 585
R334 B.n719 B.n83 585
R335 B.n925 B.n83 585
R336 B.n718 B.n717 585
R337 B.n717 B.n79 585
R338 B.n716 B.n78 585
R339 B.n931 B.n78 585
R340 B.n715 B.n77 585
R341 B.n932 B.n77 585
R342 B.n714 B.n76 585
R343 B.n933 B.n76 585
R344 B.n713 B.n712 585
R345 B.n712 B.n72 585
R346 B.n711 B.n71 585
R347 B.n939 B.n71 585
R348 B.n710 B.n70 585
R349 B.n940 B.n70 585
R350 B.n709 B.n69 585
R351 B.n941 B.n69 585
R352 B.n708 B.n707 585
R353 B.n707 B.n65 585
R354 B.n706 B.n64 585
R355 B.n947 B.n64 585
R356 B.n705 B.n63 585
R357 B.n948 B.n63 585
R358 B.n704 B.n62 585
R359 B.n949 B.n62 585
R360 B.n703 B.n702 585
R361 B.n702 B.n58 585
R362 B.n701 B.n57 585
R363 B.n955 B.n57 585
R364 B.n700 B.n56 585
R365 B.n956 B.n56 585
R366 B.n699 B.n55 585
R367 B.n957 B.n55 585
R368 B.n698 B.n697 585
R369 B.n697 B.n51 585
R370 B.n696 B.n50 585
R371 B.n963 B.n50 585
R372 B.n695 B.n49 585
R373 B.n964 B.n49 585
R374 B.n694 B.n48 585
R375 B.n965 B.n48 585
R376 B.n693 B.n692 585
R377 B.n692 B.n44 585
R378 B.n691 B.n43 585
R379 B.n971 B.n43 585
R380 B.n690 B.n42 585
R381 B.n972 B.n42 585
R382 B.n689 B.n41 585
R383 B.n973 B.n41 585
R384 B.n688 B.n687 585
R385 B.n687 B.n37 585
R386 B.n686 B.n36 585
R387 B.n979 B.n36 585
R388 B.n685 B.n35 585
R389 B.n980 B.n35 585
R390 B.n684 B.n34 585
R391 B.n981 B.n34 585
R392 B.n683 B.n682 585
R393 B.n682 B.n30 585
R394 B.n681 B.n29 585
R395 B.n987 B.n29 585
R396 B.n680 B.n28 585
R397 B.n988 B.n28 585
R398 B.n679 B.n27 585
R399 B.n989 B.n27 585
R400 B.n678 B.n677 585
R401 B.n677 B.n23 585
R402 B.n676 B.n22 585
R403 B.n995 B.n22 585
R404 B.n675 B.n21 585
R405 B.n996 B.n21 585
R406 B.n674 B.n20 585
R407 B.n997 B.n20 585
R408 B.n673 B.n672 585
R409 B.n672 B.n16 585
R410 B.n671 B.n15 585
R411 B.n1003 B.n15 585
R412 B.n670 B.n14 585
R413 B.n1004 B.n14 585
R414 B.n669 B.n13 585
R415 B.n1005 B.n13 585
R416 B.n668 B.n667 585
R417 B.n667 B.n12 585
R418 B.n666 B.n665 585
R419 B.n666 B.n8 585
R420 B.n664 B.n7 585
R421 B.n1012 B.n7 585
R422 B.n663 B.n6 585
R423 B.n1013 B.n6 585
R424 B.n662 B.n5 585
R425 B.n1014 B.n5 585
R426 B.n661 B.n660 585
R427 B.n660 B.n4 585
R428 B.n659 B.n161 585
R429 B.n659 B.n658 585
R430 B.n649 B.n162 585
R431 B.n163 B.n162 585
R432 B.n651 B.n650 585
R433 B.n652 B.n651 585
R434 B.n648 B.n168 585
R435 B.n168 B.n167 585
R436 B.n647 B.n646 585
R437 B.n646 B.n645 585
R438 B.n170 B.n169 585
R439 B.n171 B.n170 585
R440 B.n638 B.n637 585
R441 B.n639 B.n638 585
R442 B.n636 B.n176 585
R443 B.n176 B.n175 585
R444 B.n635 B.n634 585
R445 B.n634 B.n633 585
R446 B.n178 B.n177 585
R447 B.n179 B.n178 585
R448 B.n626 B.n625 585
R449 B.n627 B.n626 585
R450 B.n624 B.n184 585
R451 B.n184 B.n183 585
R452 B.n623 B.n622 585
R453 B.n622 B.n621 585
R454 B.n186 B.n185 585
R455 B.n187 B.n186 585
R456 B.n614 B.n613 585
R457 B.n615 B.n614 585
R458 B.n612 B.n192 585
R459 B.n192 B.n191 585
R460 B.n611 B.n610 585
R461 B.n610 B.n609 585
R462 B.n194 B.n193 585
R463 B.n195 B.n194 585
R464 B.n602 B.n601 585
R465 B.n603 B.n602 585
R466 B.n600 B.n200 585
R467 B.n200 B.n199 585
R468 B.n599 B.n598 585
R469 B.n598 B.n597 585
R470 B.n202 B.n201 585
R471 B.n203 B.n202 585
R472 B.n590 B.n589 585
R473 B.n591 B.n590 585
R474 B.n588 B.n208 585
R475 B.n208 B.n207 585
R476 B.n587 B.n586 585
R477 B.n586 B.n585 585
R478 B.n210 B.n209 585
R479 B.n211 B.n210 585
R480 B.n578 B.n577 585
R481 B.n579 B.n578 585
R482 B.n576 B.n216 585
R483 B.n216 B.n215 585
R484 B.n575 B.n574 585
R485 B.n574 B.n573 585
R486 B.n218 B.n217 585
R487 B.n219 B.n218 585
R488 B.n566 B.n565 585
R489 B.n567 B.n566 585
R490 B.n564 B.n224 585
R491 B.n224 B.n223 585
R492 B.n563 B.n562 585
R493 B.n562 B.n561 585
R494 B.n226 B.n225 585
R495 B.n227 B.n226 585
R496 B.n554 B.n553 585
R497 B.n555 B.n554 585
R498 B.n552 B.n232 585
R499 B.n232 B.n231 585
R500 B.n551 B.n550 585
R501 B.n550 B.n549 585
R502 B.n234 B.n233 585
R503 B.n235 B.n234 585
R504 B.n542 B.n541 585
R505 B.n543 B.n542 585
R506 B.n540 B.n240 585
R507 B.n240 B.n239 585
R508 B.n539 B.n538 585
R509 B.n538 B.n537 585
R510 B.n242 B.n241 585
R511 B.n243 B.n242 585
R512 B.n530 B.n529 585
R513 B.n531 B.n530 585
R514 B.n528 B.n248 585
R515 B.n248 B.n247 585
R516 B.n527 B.n526 585
R517 B.n526 B.n525 585
R518 B.n250 B.n249 585
R519 B.n251 B.n250 585
R520 B.n518 B.n517 585
R521 B.n519 B.n518 585
R522 B.n516 B.n256 585
R523 B.n256 B.n255 585
R524 B.n515 B.n514 585
R525 B.n514 B.n513 585
R526 B.n258 B.n257 585
R527 B.n259 B.n258 585
R528 B.n506 B.n505 585
R529 B.n507 B.n506 585
R530 B.n504 B.n264 585
R531 B.n264 B.n263 585
R532 B.n503 B.n502 585
R533 B.n502 B.n501 585
R534 B.n266 B.n265 585
R535 B.n267 B.n266 585
R536 B.n494 B.n493 585
R537 B.n495 B.n494 585
R538 B.n492 B.n272 585
R539 B.n272 B.n271 585
R540 B.n491 B.n490 585
R541 B.n490 B.n489 585
R542 B.n274 B.n273 585
R543 B.n482 B.n274 585
R544 B.n481 B.n480 585
R545 B.n483 B.n481 585
R546 B.n479 B.n279 585
R547 B.n279 B.n278 585
R548 B.n478 B.n477 585
R549 B.n477 B.n476 585
R550 B.n281 B.n280 585
R551 B.n282 B.n281 585
R552 B.n469 B.n468 585
R553 B.n470 B.n469 585
R554 B.n467 B.n287 585
R555 B.n287 B.n286 585
R556 B.n466 B.n465 585
R557 B.n465 B.n464 585
R558 B.n461 B.n291 585
R559 B.n460 B.n459 585
R560 B.n457 B.n292 585
R561 B.n457 B.n290 585
R562 B.n456 B.n455 585
R563 B.n454 B.n453 585
R564 B.n452 B.n294 585
R565 B.n450 B.n449 585
R566 B.n448 B.n295 585
R567 B.n447 B.n446 585
R568 B.n444 B.n296 585
R569 B.n442 B.n441 585
R570 B.n440 B.n297 585
R571 B.n439 B.n438 585
R572 B.n436 B.n298 585
R573 B.n434 B.n433 585
R574 B.n432 B.n299 585
R575 B.n431 B.n430 585
R576 B.n428 B.n300 585
R577 B.n426 B.n425 585
R578 B.n424 B.n301 585
R579 B.n423 B.n422 585
R580 B.n420 B.n302 585
R581 B.n418 B.n417 585
R582 B.n416 B.n303 585
R583 B.n415 B.n414 585
R584 B.n412 B.n304 585
R585 B.n410 B.n409 585
R586 B.n408 B.n305 585
R587 B.n407 B.n406 585
R588 B.n404 B.n403 585
R589 B.n402 B.n401 585
R590 B.n400 B.n310 585
R591 B.n398 B.n397 585
R592 B.n396 B.n311 585
R593 B.n395 B.n394 585
R594 B.n392 B.n312 585
R595 B.n390 B.n389 585
R596 B.n388 B.n313 585
R597 B.n386 B.n385 585
R598 B.n383 B.n316 585
R599 B.n381 B.n380 585
R600 B.n379 B.n317 585
R601 B.n378 B.n377 585
R602 B.n375 B.n318 585
R603 B.n373 B.n372 585
R604 B.n371 B.n319 585
R605 B.n370 B.n369 585
R606 B.n367 B.n320 585
R607 B.n365 B.n364 585
R608 B.n363 B.n321 585
R609 B.n362 B.n361 585
R610 B.n359 B.n322 585
R611 B.n357 B.n356 585
R612 B.n355 B.n323 585
R613 B.n354 B.n353 585
R614 B.n351 B.n324 585
R615 B.n349 B.n348 585
R616 B.n347 B.n325 585
R617 B.n346 B.n345 585
R618 B.n343 B.n326 585
R619 B.n341 B.n340 585
R620 B.n339 B.n327 585
R621 B.n338 B.n337 585
R622 B.n335 B.n328 585
R623 B.n333 B.n332 585
R624 B.n331 B.n330 585
R625 B.n289 B.n288 585
R626 B.n463 B.n462 585
R627 B.n464 B.n463 585
R628 B.n285 B.n284 585
R629 B.n286 B.n285 585
R630 B.n472 B.n471 585
R631 B.n471 B.n470 585
R632 B.n473 B.n283 585
R633 B.n283 B.n282 585
R634 B.n475 B.n474 585
R635 B.n476 B.n475 585
R636 B.n277 B.n276 585
R637 B.n278 B.n277 585
R638 B.n485 B.n484 585
R639 B.n484 B.n483 585
R640 B.n486 B.n275 585
R641 B.n482 B.n275 585
R642 B.n488 B.n487 585
R643 B.n489 B.n488 585
R644 B.n270 B.n269 585
R645 B.n271 B.n270 585
R646 B.n497 B.n496 585
R647 B.n496 B.n495 585
R648 B.n498 B.n268 585
R649 B.n268 B.n267 585
R650 B.n500 B.n499 585
R651 B.n501 B.n500 585
R652 B.n262 B.n261 585
R653 B.n263 B.n262 585
R654 B.n509 B.n508 585
R655 B.n508 B.n507 585
R656 B.n510 B.n260 585
R657 B.n260 B.n259 585
R658 B.n512 B.n511 585
R659 B.n513 B.n512 585
R660 B.n254 B.n253 585
R661 B.n255 B.n254 585
R662 B.n521 B.n520 585
R663 B.n520 B.n519 585
R664 B.n522 B.n252 585
R665 B.n252 B.n251 585
R666 B.n524 B.n523 585
R667 B.n525 B.n524 585
R668 B.n246 B.n245 585
R669 B.n247 B.n246 585
R670 B.n533 B.n532 585
R671 B.n532 B.n531 585
R672 B.n534 B.n244 585
R673 B.n244 B.n243 585
R674 B.n536 B.n535 585
R675 B.n537 B.n536 585
R676 B.n238 B.n237 585
R677 B.n239 B.n238 585
R678 B.n545 B.n544 585
R679 B.n544 B.n543 585
R680 B.n546 B.n236 585
R681 B.n236 B.n235 585
R682 B.n548 B.n547 585
R683 B.n549 B.n548 585
R684 B.n230 B.n229 585
R685 B.n231 B.n230 585
R686 B.n557 B.n556 585
R687 B.n556 B.n555 585
R688 B.n558 B.n228 585
R689 B.n228 B.n227 585
R690 B.n560 B.n559 585
R691 B.n561 B.n560 585
R692 B.n222 B.n221 585
R693 B.n223 B.n222 585
R694 B.n569 B.n568 585
R695 B.n568 B.n567 585
R696 B.n570 B.n220 585
R697 B.n220 B.n219 585
R698 B.n572 B.n571 585
R699 B.n573 B.n572 585
R700 B.n214 B.n213 585
R701 B.n215 B.n214 585
R702 B.n581 B.n580 585
R703 B.n580 B.n579 585
R704 B.n582 B.n212 585
R705 B.n212 B.n211 585
R706 B.n584 B.n583 585
R707 B.n585 B.n584 585
R708 B.n206 B.n205 585
R709 B.n207 B.n206 585
R710 B.n593 B.n592 585
R711 B.n592 B.n591 585
R712 B.n594 B.n204 585
R713 B.n204 B.n203 585
R714 B.n596 B.n595 585
R715 B.n597 B.n596 585
R716 B.n198 B.n197 585
R717 B.n199 B.n198 585
R718 B.n605 B.n604 585
R719 B.n604 B.n603 585
R720 B.n606 B.n196 585
R721 B.n196 B.n195 585
R722 B.n608 B.n607 585
R723 B.n609 B.n608 585
R724 B.n190 B.n189 585
R725 B.n191 B.n190 585
R726 B.n617 B.n616 585
R727 B.n616 B.n615 585
R728 B.n618 B.n188 585
R729 B.n188 B.n187 585
R730 B.n620 B.n619 585
R731 B.n621 B.n620 585
R732 B.n182 B.n181 585
R733 B.n183 B.n182 585
R734 B.n629 B.n628 585
R735 B.n628 B.n627 585
R736 B.n630 B.n180 585
R737 B.n180 B.n179 585
R738 B.n632 B.n631 585
R739 B.n633 B.n632 585
R740 B.n174 B.n173 585
R741 B.n175 B.n174 585
R742 B.n641 B.n640 585
R743 B.n640 B.n639 585
R744 B.n642 B.n172 585
R745 B.n172 B.n171 585
R746 B.n644 B.n643 585
R747 B.n645 B.n644 585
R748 B.n166 B.n165 585
R749 B.n167 B.n166 585
R750 B.n654 B.n653 585
R751 B.n653 B.n652 585
R752 B.n655 B.n164 585
R753 B.n164 B.n163 585
R754 B.n657 B.n656 585
R755 B.n658 B.n657 585
R756 B.n3 B.n0 585
R757 B.n4 B.n3 585
R758 B.n1011 B.n1 585
R759 B.n1012 B.n1011 585
R760 B.n1010 B.n1009 585
R761 B.n1010 B.n8 585
R762 B.n1008 B.n9 585
R763 B.n12 B.n9 585
R764 B.n1007 B.n1006 585
R765 B.n1006 B.n1005 585
R766 B.n11 B.n10 585
R767 B.n1004 B.n11 585
R768 B.n1002 B.n1001 585
R769 B.n1003 B.n1002 585
R770 B.n1000 B.n17 585
R771 B.n17 B.n16 585
R772 B.n999 B.n998 585
R773 B.n998 B.n997 585
R774 B.n19 B.n18 585
R775 B.n996 B.n19 585
R776 B.n994 B.n993 585
R777 B.n995 B.n994 585
R778 B.n992 B.n24 585
R779 B.n24 B.n23 585
R780 B.n991 B.n990 585
R781 B.n990 B.n989 585
R782 B.n26 B.n25 585
R783 B.n988 B.n26 585
R784 B.n986 B.n985 585
R785 B.n987 B.n986 585
R786 B.n984 B.n31 585
R787 B.n31 B.n30 585
R788 B.n983 B.n982 585
R789 B.n982 B.n981 585
R790 B.n33 B.n32 585
R791 B.n980 B.n33 585
R792 B.n978 B.n977 585
R793 B.n979 B.n978 585
R794 B.n976 B.n38 585
R795 B.n38 B.n37 585
R796 B.n975 B.n974 585
R797 B.n974 B.n973 585
R798 B.n40 B.n39 585
R799 B.n972 B.n40 585
R800 B.n970 B.n969 585
R801 B.n971 B.n970 585
R802 B.n968 B.n45 585
R803 B.n45 B.n44 585
R804 B.n967 B.n966 585
R805 B.n966 B.n965 585
R806 B.n47 B.n46 585
R807 B.n964 B.n47 585
R808 B.n962 B.n961 585
R809 B.n963 B.n962 585
R810 B.n960 B.n52 585
R811 B.n52 B.n51 585
R812 B.n959 B.n958 585
R813 B.n958 B.n957 585
R814 B.n54 B.n53 585
R815 B.n956 B.n54 585
R816 B.n954 B.n953 585
R817 B.n955 B.n954 585
R818 B.n952 B.n59 585
R819 B.n59 B.n58 585
R820 B.n951 B.n950 585
R821 B.n950 B.n949 585
R822 B.n61 B.n60 585
R823 B.n948 B.n61 585
R824 B.n946 B.n945 585
R825 B.n947 B.n946 585
R826 B.n944 B.n66 585
R827 B.n66 B.n65 585
R828 B.n943 B.n942 585
R829 B.n942 B.n941 585
R830 B.n68 B.n67 585
R831 B.n940 B.n68 585
R832 B.n938 B.n937 585
R833 B.n939 B.n938 585
R834 B.n936 B.n73 585
R835 B.n73 B.n72 585
R836 B.n935 B.n934 585
R837 B.n934 B.n933 585
R838 B.n75 B.n74 585
R839 B.n932 B.n75 585
R840 B.n930 B.n929 585
R841 B.n931 B.n930 585
R842 B.n928 B.n80 585
R843 B.n80 B.n79 585
R844 B.n927 B.n926 585
R845 B.n926 B.n925 585
R846 B.n82 B.n81 585
R847 B.n924 B.n82 585
R848 B.n922 B.n921 585
R849 B.n923 B.n922 585
R850 B.n920 B.n87 585
R851 B.n87 B.n86 585
R852 B.n919 B.n918 585
R853 B.n918 B.n917 585
R854 B.n89 B.n88 585
R855 B.n916 B.n89 585
R856 B.n914 B.n913 585
R857 B.n915 B.n914 585
R858 B.n912 B.n94 585
R859 B.n94 B.n93 585
R860 B.n911 B.n910 585
R861 B.n910 B.n909 585
R862 B.n96 B.n95 585
R863 B.n908 B.n96 585
R864 B.n906 B.n905 585
R865 B.n907 B.n906 585
R866 B.n904 B.n101 585
R867 B.n101 B.n100 585
R868 B.n903 B.n902 585
R869 B.n902 B.n901 585
R870 B.n103 B.n102 585
R871 B.n900 B.n103 585
R872 B.n898 B.n897 585
R873 B.n899 B.n898 585
R874 B.n896 B.n107 585
R875 B.n110 B.n107 585
R876 B.n895 B.n894 585
R877 B.n894 B.n893 585
R878 B.n109 B.n108 585
R879 B.n892 B.n109 585
R880 B.n890 B.n889 585
R881 B.n891 B.n890 585
R882 B.n888 B.n115 585
R883 B.n115 B.n114 585
R884 B.n887 B.n886 585
R885 B.n886 B.n885 585
R886 B.n117 B.n116 585
R887 B.n884 B.n117 585
R888 B.n882 B.n881 585
R889 B.n883 B.n882 585
R890 B.n1015 B.n1014 585
R891 B.n1013 B.n2 585
R892 B.n882 B.n122 511.721
R893 B.n160 B.n120 511.721
R894 B.n465 B.n289 511.721
R895 B.n463 B.n291 511.721
R896 B.n137 B.t14 269.584
R897 B.n143 B.t18 269.584
R898 B.n314 B.t10 269.584
R899 B.n306 B.t21 269.584
R900 B.n750 B.n121 256.663
R901 B.n752 B.n121 256.663
R902 B.n758 B.n121 256.663
R903 B.n760 B.n121 256.663
R904 B.n766 B.n121 256.663
R905 B.n768 B.n121 256.663
R906 B.n774 B.n121 256.663
R907 B.n776 B.n121 256.663
R908 B.n782 B.n121 256.663
R909 B.n784 B.n121 256.663
R910 B.n790 B.n121 256.663
R911 B.n792 B.n121 256.663
R912 B.n798 B.n121 256.663
R913 B.n146 B.n121 256.663
R914 B.n804 B.n121 256.663
R915 B.n810 B.n121 256.663
R916 B.n812 B.n121 256.663
R917 B.n818 B.n121 256.663
R918 B.n820 B.n121 256.663
R919 B.n827 B.n121 256.663
R920 B.n829 B.n121 256.663
R921 B.n835 B.n121 256.663
R922 B.n837 B.n121 256.663
R923 B.n843 B.n121 256.663
R924 B.n845 B.n121 256.663
R925 B.n851 B.n121 256.663
R926 B.n853 B.n121 256.663
R927 B.n859 B.n121 256.663
R928 B.n861 B.n121 256.663
R929 B.n867 B.n121 256.663
R930 B.n869 B.n121 256.663
R931 B.n875 B.n121 256.663
R932 B.n877 B.n121 256.663
R933 B.n458 B.n290 256.663
R934 B.n293 B.n290 256.663
R935 B.n451 B.n290 256.663
R936 B.n445 B.n290 256.663
R937 B.n443 B.n290 256.663
R938 B.n437 B.n290 256.663
R939 B.n435 B.n290 256.663
R940 B.n429 B.n290 256.663
R941 B.n427 B.n290 256.663
R942 B.n421 B.n290 256.663
R943 B.n419 B.n290 256.663
R944 B.n413 B.n290 256.663
R945 B.n411 B.n290 256.663
R946 B.n405 B.n290 256.663
R947 B.n309 B.n290 256.663
R948 B.n399 B.n290 256.663
R949 B.n393 B.n290 256.663
R950 B.n391 B.n290 256.663
R951 B.n384 B.n290 256.663
R952 B.n382 B.n290 256.663
R953 B.n376 B.n290 256.663
R954 B.n374 B.n290 256.663
R955 B.n368 B.n290 256.663
R956 B.n366 B.n290 256.663
R957 B.n360 B.n290 256.663
R958 B.n358 B.n290 256.663
R959 B.n352 B.n290 256.663
R960 B.n350 B.n290 256.663
R961 B.n344 B.n290 256.663
R962 B.n342 B.n290 256.663
R963 B.n336 B.n290 256.663
R964 B.n334 B.n290 256.663
R965 B.n329 B.n290 256.663
R966 B.n1017 B.n1016 256.663
R967 B.n878 B.n876 163.367
R968 B.n874 B.n124 163.367
R969 B.n870 B.n868 163.367
R970 B.n866 B.n126 163.367
R971 B.n862 B.n860 163.367
R972 B.n858 B.n128 163.367
R973 B.n854 B.n852 163.367
R974 B.n850 B.n130 163.367
R975 B.n846 B.n844 163.367
R976 B.n842 B.n132 163.367
R977 B.n838 B.n836 163.367
R978 B.n834 B.n134 163.367
R979 B.n830 B.n828 163.367
R980 B.n826 B.n136 163.367
R981 B.n821 B.n819 163.367
R982 B.n817 B.n140 163.367
R983 B.n813 B.n811 163.367
R984 B.n809 B.n142 163.367
R985 B.n805 B.n803 163.367
R986 B.n800 B.n799 163.367
R987 B.n797 B.n148 163.367
R988 B.n793 B.n791 163.367
R989 B.n789 B.n150 163.367
R990 B.n785 B.n783 163.367
R991 B.n781 B.n152 163.367
R992 B.n777 B.n775 163.367
R993 B.n773 B.n154 163.367
R994 B.n769 B.n767 163.367
R995 B.n765 B.n156 163.367
R996 B.n761 B.n759 163.367
R997 B.n757 B.n158 163.367
R998 B.n753 B.n751 163.367
R999 B.n749 B.n160 163.367
R1000 B.n465 B.n287 163.367
R1001 B.n469 B.n287 163.367
R1002 B.n469 B.n281 163.367
R1003 B.n477 B.n281 163.367
R1004 B.n477 B.n279 163.367
R1005 B.n481 B.n279 163.367
R1006 B.n481 B.n274 163.367
R1007 B.n490 B.n274 163.367
R1008 B.n490 B.n272 163.367
R1009 B.n494 B.n272 163.367
R1010 B.n494 B.n266 163.367
R1011 B.n502 B.n266 163.367
R1012 B.n502 B.n264 163.367
R1013 B.n506 B.n264 163.367
R1014 B.n506 B.n258 163.367
R1015 B.n514 B.n258 163.367
R1016 B.n514 B.n256 163.367
R1017 B.n518 B.n256 163.367
R1018 B.n518 B.n250 163.367
R1019 B.n526 B.n250 163.367
R1020 B.n526 B.n248 163.367
R1021 B.n530 B.n248 163.367
R1022 B.n530 B.n242 163.367
R1023 B.n538 B.n242 163.367
R1024 B.n538 B.n240 163.367
R1025 B.n542 B.n240 163.367
R1026 B.n542 B.n234 163.367
R1027 B.n550 B.n234 163.367
R1028 B.n550 B.n232 163.367
R1029 B.n554 B.n232 163.367
R1030 B.n554 B.n226 163.367
R1031 B.n562 B.n226 163.367
R1032 B.n562 B.n224 163.367
R1033 B.n566 B.n224 163.367
R1034 B.n566 B.n218 163.367
R1035 B.n574 B.n218 163.367
R1036 B.n574 B.n216 163.367
R1037 B.n578 B.n216 163.367
R1038 B.n578 B.n210 163.367
R1039 B.n586 B.n210 163.367
R1040 B.n586 B.n208 163.367
R1041 B.n590 B.n208 163.367
R1042 B.n590 B.n202 163.367
R1043 B.n598 B.n202 163.367
R1044 B.n598 B.n200 163.367
R1045 B.n602 B.n200 163.367
R1046 B.n602 B.n194 163.367
R1047 B.n610 B.n194 163.367
R1048 B.n610 B.n192 163.367
R1049 B.n614 B.n192 163.367
R1050 B.n614 B.n186 163.367
R1051 B.n622 B.n186 163.367
R1052 B.n622 B.n184 163.367
R1053 B.n626 B.n184 163.367
R1054 B.n626 B.n178 163.367
R1055 B.n634 B.n178 163.367
R1056 B.n634 B.n176 163.367
R1057 B.n638 B.n176 163.367
R1058 B.n638 B.n170 163.367
R1059 B.n646 B.n170 163.367
R1060 B.n646 B.n168 163.367
R1061 B.n651 B.n168 163.367
R1062 B.n651 B.n162 163.367
R1063 B.n659 B.n162 163.367
R1064 B.n660 B.n659 163.367
R1065 B.n660 B.n5 163.367
R1066 B.n6 B.n5 163.367
R1067 B.n7 B.n6 163.367
R1068 B.n666 B.n7 163.367
R1069 B.n667 B.n666 163.367
R1070 B.n667 B.n13 163.367
R1071 B.n14 B.n13 163.367
R1072 B.n15 B.n14 163.367
R1073 B.n672 B.n15 163.367
R1074 B.n672 B.n20 163.367
R1075 B.n21 B.n20 163.367
R1076 B.n22 B.n21 163.367
R1077 B.n677 B.n22 163.367
R1078 B.n677 B.n27 163.367
R1079 B.n28 B.n27 163.367
R1080 B.n29 B.n28 163.367
R1081 B.n682 B.n29 163.367
R1082 B.n682 B.n34 163.367
R1083 B.n35 B.n34 163.367
R1084 B.n36 B.n35 163.367
R1085 B.n687 B.n36 163.367
R1086 B.n687 B.n41 163.367
R1087 B.n42 B.n41 163.367
R1088 B.n43 B.n42 163.367
R1089 B.n692 B.n43 163.367
R1090 B.n692 B.n48 163.367
R1091 B.n49 B.n48 163.367
R1092 B.n50 B.n49 163.367
R1093 B.n697 B.n50 163.367
R1094 B.n697 B.n55 163.367
R1095 B.n56 B.n55 163.367
R1096 B.n57 B.n56 163.367
R1097 B.n702 B.n57 163.367
R1098 B.n702 B.n62 163.367
R1099 B.n63 B.n62 163.367
R1100 B.n64 B.n63 163.367
R1101 B.n707 B.n64 163.367
R1102 B.n707 B.n69 163.367
R1103 B.n70 B.n69 163.367
R1104 B.n71 B.n70 163.367
R1105 B.n712 B.n71 163.367
R1106 B.n712 B.n76 163.367
R1107 B.n77 B.n76 163.367
R1108 B.n78 B.n77 163.367
R1109 B.n717 B.n78 163.367
R1110 B.n717 B.n83 163.367
R1111 B.n84 B.n83 163.367
R1112 B.n85 B.n84 163.367
R1113 B.n722 B.n85 163.367
R1114 B.n722 B.n90 163.367
R1115 B.n91 B.n90 163.367
R1116 B.n92 B.n91 163.367
R1117 B.n727 B.n92 163.367
R1118 B.n727 B.n97 163.367
R1119 B.n98 B.n97 163.367
R1120 B.n99 B.n98 163.367
R1121 B.n732 B.n99 163.367
R1122 B.n732 B.n104 163.367
R1123 B.n105 B.n104 163.367
R1124 B.n106 B.n105 163.367
R1125 B.n737 B.n106 163.367
R1126 B.n737 B.n111 163.367
R1127 B.n112 B.n111 163.367
R1128 B.n113 B.n112 163.367
R1129 B.n742 B.n113 163.367
R1130 B.n742 B.n118 163.367
R1131 B.n119 B.n118 163.367
R1132 B.n120 B.n119 163.367
R1133 B.n459 B.n457 163.367
R1134 B.n457 B.n456 163.367
R1135 B.n453 B.n452 163.367
R1136 B.n450 B.n295 163.367
R1137 B.n446 B.n444 163.367
R1138 B.n442 B.n297 163.367
R1139 B.n438 B.n436 163.367
R1140 B.n434 B.n299 163.367
R1141 B.n430 B.n428 163.367
R1142 B.n426 B.n301 163.367
R1143 B.n422 B.n420 163.367
R1144 B.n418 B.n303 163.367
R1145 B.n414 B.n412 163.367
R1146 B.n410 B.n305 163.367
R1147 B.n406 B.n404 163.367
R1148 B.n401 B.n400 163.367
R1149 B.n398 B.n311 163.367
R1150 B.n394 B.n392 163.367
R1151 B.n390 B.n313 163.367
R1152 B.n385 B.n383 163.367
R1153 B.n381 B.n317 163.367
R1154 B.n377 B.n375 163.367
R1155 B.n373 B.n319 163.367
R1156 B.n369 B.n367 163.367
R1157 B.n365 B.n321 163.367
R1158 B.n361 B.n359 163.367
R1159 B.n357 B.n323 163.367
R1160 B.n353 B.n351 163.367
R1161 B.n349 B.n325 163.367
R1162 B.n345 B.n343 163.367
R1163 B.n341 B.n327 163.367
R1164 B.n337 B.n335 163.367
R1165 B.n333 B.n330 163.367
R1166 B.n463 B.n285 163.367
R1167 B.n471 B.n285 163.367
R1168 B.n471 B.n283 163.367
R1169 B.n475 B.n283 163.367
R1170 B.n475 B.n277 163.367
R1171 B.n484 B.n277 163.367
R1172 B.n484 B.n275 163.367
R1173 B.n488 B.n275 163.367
R1174 B.n488 B.n270 163.367
R1175 B.n496 B.n270 163.367
R1176 B.n496 B.n268 163.367
R1177 B.n500 B.n268 163.367
R1178 B.n500 B.n262 163.367
R1179 B.n508 B.n262 163.367
R1180 B.n508 B.n260 163.367
R1181 B.n512 B.n260 163.367
R1182 B.n512 B.n254 163.367
R1183 B.n520 B.n254 163.367
R1184 B.n520 B.n252 163.367
R1185 B.n524 B.n252 163.367
R1186 B.n524 B.n246 163.367
R1187 B.n532 B.n246 163.367
R1188 B.n532 B.n244 163.367
R1189 B.n536 B.n244 163.367
R1190 B.n536 B.n238 163.367
R1191 B.n544 B.n238 163.367
R1192 B.n544 B.n236 163.367
R1193 B.n548 B.n236 163.367
R1194 B.n548 B.n230 163.367
R1195 B.n556 B.n230 163.367
R1196 B.n556 B.n228 163.367
R1197 B.n560 B.n228 163.367
R1198 B.n560 B.n222 163.367
R1199 B.n568 B.n222 163.367
R1200 B.n568 B.n220 163.367
R1201 B.n572 B.n220 163.367
R1202 B.n572 B.n214 163.367
R1203 B.n580 B.n214 163.367
R1204 B.n580 B.n212 163.367
R1205 B.n584 B.n212 163.367
R1206 B.n584 B.n206 163.367
R1207 B.n592 B.n206 163.367
R1208 B.n592 B.n204 163.367
R1209 B.n596 B.n204 163.367
R1210 B.n596 B.n198 163.367
R1211 B.n604 B.n198 163.367
R1212 B.n604 B.n196 163.367
R1213 B.n608 B.n196 163.367
R1214 B.n608 B.n190 163.367
R1215 B.n616 B.n190 163.367
R1216 B.n616 B.n188 163.367
R1217 B.n620 B.n188 163.367
R1218 B.n620 B.n182 163.367
R1219 B.n628 B.n182 163.367
R1220 B.n628 B.n180 163.367
R1221 B.n632 B.n180 163.367
R1222 B.n632 B.n174 163.367
R1223 B.n640 B.n174 163.367
R1224 B.n640 B.n172 163.367
R1225 B.n644 B.n172 163.367
R1226 B.n644 B.n166 163.367
R1227 B.n653 B.n166 163.367
R1228 B.n653 B.n164 163.367
R1229 B.n657 B.n164 163.367
R1230 B.n657 B.n3 163.367
R1231 B.n1015 B.n3 163.367
R1232 B.n1011 B.n2 163.367
R1233 B.n1011 B.n1010 163.367
R1234 B.n1010 B.n9 163.367
R1235 B.n1006 B.n9 163.367
R1236 B.n1006 B.n11 163.367
R1237 B.n1002 B.n11 163.367
R1238 B.n1002 B.n17 163.367
R1239 B.n998 B.n17 163.367
R1240 B.n998 B.n19 163.367
R1241 B.n994 B.n19 163.367
R1242 B.n994 B.n24 163.367
R1243 B.n990 B.n24 163.367
R1244 B.n990 B.n26 163.367
R1245 B.n986 B.n26 163.367
R1246 B.n986 B.n31 163.367
R1247 B.n982 B.n31 163.367
R1248 B.n982 B.n33 163.367
R1249 B.n978 B.n33 163.367
R1250 B.n978 B.n38 163.367
R1251 B.n974 B.n38 163.367
R1252 B.n974 B.n40 163.367
R1253 B.n970 B.n40 163.367
R1254 B.n970 B.n45 163.367
R1255 B.n966 B.n45 163.367
R1256 B.n966 B.n47 163.367
R1257 B.n962 B.n47 163.367
R1258 B.n962 B.n52 163.367
R1259 B.n958 B.n52 163.367
R1260 B.n958 B.n54 163.367
R1261 B.n954 B.n54 163.367
R1262 B.n954 B.n59 163.367
R1263 B.n950 B.n59 163.367
R1264 B.n950 B.n61 163.367
R1265 B.n946 B.n61 163.367
R1266 B.n946 B.n66 163.367
R1267 B.n942 B.n66 163.367
R1268 B.n942 B.n68 163.367
R1269 B.n938 B.n68 163.367
R1270 B.n938 B.n73 163.367
R1271 B.n934 B.n73 163.367
R1272 B.n934 B.n75 163.367
R1273 B.n930 B.n75 163.367
R1274 B.n930 B.n80 163.367
R1275 B.n926 B.n80 163.367
R1276 B.n926 B.n82 163.367
R1277 B.n922 B.n82 163.367
R1278 B.n922 B.n87 163.367
R1279 B.n918 B.n87 163.367
R1280 B.n918 B.n89 163.367
R1281 B.n914 B.n89 163.367
R1282 B.n914 B.n94 163.367
R1283 B.n910 B.n94 163.367
R1284 B.n910 B.n96 163.367
R1285 B.n906 B.n96 163.367
R1286 B.n906 B.n101 163.367
R1287 B.n902 B.n101 163.367
R1288 B.n902 B.n103 163.367
R1289 B.n898 B.n103 163.367
R1290 B.n898 B.n107 163.367
R1291 B.n894 B.n107 163.367
R1292 B.n894 B.n109 163.367
R1293 B.n890 B.n109 163.367
R1294 B.n890 B.n115 163.367
R1295 B.n886 B.n115 163.367
R1296 B.n886 B.n117 163.367
R1297 B.n882 B.n117 163.367
R1298 B.n143 B.t19 134.883
R1299 B.n314 B.t13 134.883
R1300 B.n137 B.t16 134.875
R1301 B.n306 B.t23 134.875
R1302 B.n464 B.n290 117.323
R1303 B.n883 B.n121 117.323
R1304 B.n877 B.n122 71.676
R1305 B.n876 B.n875 71.676
R1306 B.n869 B.n124 71.676
R1307 B.n868 B.n867 71.676
R1308 B.n861 B.n126 71.676
R1309 B.n860 B.n859 71.676
R1310 B.n853 B.n128 71.676
R1311 B.n852 B.n851 71.676
R1312 B.n845 B.n130 71.676
R1313 B.n844 B.n843 71.676
R1314 B.n837 B.n132 71.676
R1315 B.n836 B.n835 71.676
R1316 B.n829 B.n134 71.676
R1317 B.n828 B.n827 71.676
R1318 B.n820 B.n136 71.676
R1319 B.n819 B.n818 71.676
R1320 B.n812 B.n140 71.676
R1321 B.n811 B.n810 71.676
R1322 B.n804 B.n142 71.676
R1323 B.n803 B.n146 71.676
R1324 B.n799 B.n798 71.676
R1325 B.n792 B.n148 71.676
R1326 B.n791 B.n790 71.676
R1327 B.n784 B.n150 71.676
R1328 B.n783 B.n782 71.676
R1329 B.n776 B.n152 71.676
R1330 B.n775 B.n774 71.676
R1331 B.n768 B.n154 71.676
R1332 B.n767 B.n766 71.676
R1333 B.n760 B.n156 71.676
R1334 B.n759 B.n758 71.676
R1335 B.n752 B.n158 71.676
R1336 B.n751 B.n750 71.676
R1337 B.n750 B.n749 71.676
R1338 B.n753 B.n752 71.676
R1339 B.n758 B.n757 71.676
R1340 B.n761 B.n760 71.676
R1341 B.n766 B.n765 71.676
R1342 B.n769 B.n768 71.676
R1343 B.n774 B.n773 71.676
R1344 B.n777 B.n776 71.676
R1345 B.n782 B.n781 71.676
R1346 B.n785 B.n784 71.676
R1347 B.n790 B.n789 71.676
R1348 B.n793 B.n792 71.676
R1349 B.n798 B.n797 71.676
R1350 B.n800 B.n146 71.676
R1351 B.n805 B.n804 71.676
R1352 B.n810 B.n809 71.676
R1353 B.n813 B.n812 71.676
R1354 B.n818 B.n817 71.676
R1355 B.n821 B.n820 71.676
R1356 B.n827 B.n826 71.676
R1357 B.n830 B.n829 71.676
R1358 B.n835 B.n834 71.676
R1359 B.n838 B.n837 71.676
R1360 B.n843 B.n842 71.676
R1361 B.n846 B.n845 71.676
R1362 B.n851 B.n850 71.676
R1363 B.n854 B.n853 71.676
R1364 B.n859 B.n858 71.676
R1365 B.n862 B.n861 71.676
R1366 B.n867 B.n866 71.676
R1367 B.n870 B.n869 71.676
R1368 B.n875 B.n874 71.676
R1369 B.n878 B.n877 71.676
R1370 B.n458 B.n291 71.676
R1371 B.n456 B.n293 71.676
R1372 B.n452 B.n451 71.676
R1373 B.n445 B.n295 71.676
R1374 B.n444 B.n443 71.676
R1375 B.n437 B.n297 71.676
R1376 B.n436 B.n435 71.676
R1377 B.n429 B.n299 71.676
R1378 B.n428 B.n427 71.676
R1379 B.n421 B.n301 71.676
R1380 B.n420 B.n419 71.676
R1381 B.n413 B.n303 71.676
R1382 B.n412 B.n411 71.676
R1383 B.n405 B.n305 71.676
R1384 B.n404 B.n309 71.676
R1385 B.n400 B.n399 71.676
R1386 B.n393 B.n311 71.676
R1387 B.n392 B.n391 71.676
R1388 B.n384 B.n313 71.676
R1389 B.n383 B.n382 71.676
R1390 B.n376 B.n317 71.676
R1391 B.n375 B.n374 71.676
R1392 B.n368 B.n319 71.676
R1393 B.n367 B.n366 71.676
R1394 B.n360 B.n321 71.676
R1395 B.n359 B.n358 71.676
R1396 B.n352 B.n323 71.676
R1397 B.n351 B.n350 71.676
R1398 B.n344 B.n325 71.676
R1399 B.n343 B.n342 71.676
R1400 B.n336 B.n327 71.676
R1401 B.n335 B.n334 71.676
R1402 B.n330 B.n329 71.676
R1403 B.n459 B.n458 71.676
R1404 B.n453 B.n293 71.676
R1405 B.n451 B.n450 71.676
R1406 B.n446 B.n445 71.676
R1407 B.n443 B.n442 71.676
R1408 B.n438 B.n437 71.676
R1409 B.n435 B.n434 71.676
R1410 B.n430 B.n429 71.676
R1411 B.n427 B.n426 71.676
R1412 B.n422 B.n421 71.676
R1413 B.n419 B.n418 71.676
R1414 B.n414 B.n413 71.676
R1415 B.n411 B.n410 71.676
R1416 B.n406 B.n405 71.676
R1417 B.n401 B.n309 71.676
R1418 B.n399 B.n398 71.676
R1419 B.n394 B.n393 71.676
R1420 B.n391 B.n390 71.676
R1421 B.n385 B.n384 71.676
R1422 B.n382 B.n381 71.676
R1423 B.n377 B.n376 71.676
R1424 B.n374 B.n373 71.676
R1425 B.n369 B.n368 71.676
R1426 B.n366 B.n365 71.676
R1427 B.n361 B.n360 71.676
R1428 B.n358 B.n357 71.676
R1429 B.n353 B.n352 71.676
R1430 B.n350 B.n349 71.676
R1431 B.n345 B.n344 71.676
R1432 B.n342 B.n341 71.676
R1433 B.n337 B.n336 71.676
R1434 B.n334 B.n333 71.676
R1435 B.n329 B.n289 71.676
R1436 B.n1016 B.n1015 71.676
R1437 B.n1016 B.n2 71.676
R1438 B.n144 B.t20 70.4958
R1439 B.n315 B.t12 70.4958
R1440 B.n138 B.t17 70.4871
R1441 B.n307 B.t22 70.4871
R1442 B.n138 B.n137 64.3884
R1443 B.n144 B.n143 64.3884
R1444 B.n315 B.n314 64.3884
R1445 B.n307 B.n306 64.3884
R1446 B.n823 B.n138 59.5399
R1447 B.n145 B.n144 59.5399
R1448 B.n387 B.n315 59.5399
R1449 B.n308 B.n307 59.5399
R1450 B.n464 B.n286 58.2333
R1451 B.n470 B.n286 58.2333
R1452 B.n470 B.n282 58.2333
R1453 B.n476 B.n282 58.2333
R1454 B.n476 B.n278 58.2333
R1455 B.n483 B.n278 58.2333
R1456 B.n483 B.n482 58.2333
R1457 B.n489 B.n271 58.2333
R1458 B.n495 B.n271 58.2333
R1459 B.n495 B.n267 58.2333
R1460 B.n501 B.n267 58.2333
R1461 B.n501 B.n263 58.2333
R1462 B.n507 B.n263 58.2333
R1463 B.n507 B.n259 58.2333
R1464 B.n513 B.n259 58.2333
R1465 B.n513 B.n255 58.2333
R1466 B.n519 B.n255 58.2333
R1467 B.n519 B.n251 58.2333
R1468 B.n525 B.n251 58.2333
R1469 B.n531 B.n247 58.2333
R1470 B.n531 B.n243 58.2333
R1471 B.n537 B.n243 58.2333
R1472 B.n537 B.n239 58.2333
R1473 B.n543 B.n239 58.2333
R1474 B.n543 B.n235 58.2333
R1475 B.n549 B.n235 58.2333
R1476 B.n549 B.n231 58.2333
R1477 B.n555 B.n231 58.2333
R1478 B.n561 B.n227 58.2333
R1479 B.n561 B.n223 58.2333
R1480 B.n567 B.n223 58.2333
R1481 B.n567 B.n219 58.2333
R1482 B.n573 B.n219 58.2333
R1483 B.n573 B.n215 58.2333
R1484 B.n579 B.n215 58.2333
R1485 B.n579 B.n211 58.2333
R1486 B.n585 B.n211 58.2333
R1487 B.n591 B.n207 58.2333
R1488 B.n591 B.n203 58.2333
R1489 B.n597 B.n203 58.2333
R1490 B.n597 B.n199 58.2333
R1491 B.n603 B.n199 58.2333
R1492 B.n603 B.n195 58.2333
R1493 B.n609 B.n195 58.2333
R1494 B.n609 B.n191 58.2333
R1495 B.n615 B.n191 58.2333
R1496 B.n621 B.n187 58.2333
R1497 B.n621 B.n183 58.2333
R1498 B.n627 B.n183 58.2333
R1499 B.n627 B.n179 58.2333
R1500 B.n633 B.n179 58.2333
R1501 B.n633 B.n175 58.2333
R1502 B.n639 B.n175 58.2333
R1503 B.n639 B.n171 58.2333
R1504 B.n645 B.n171 58.2333
R1505 B.n652 B.n167 58.2333
R1506 B.n652 B.n163 58.2333
R1507 B.n658 B.n163 58.2333
R1508 B.n658 B.n4 58.2333
R1509 B.n1014 B.n4 58.2333
R1510 B.n1014 B.n1013 58.2333
R1511 B.n1013 B.n1012 58.2333
R1512 B.n1012 B.n8 58.2333
R1513 B.n12 B.n8 58.2333
R1514 B.n1005 B.n12 58.2333
R1515 B.n1005 B.n1004 58.2333
R1516 B.n1003 B.n16 58.2333
R1517 B.n997 B.n16 58.2333
R1518 B.n997 B.n996 58.2333
R1519 B.n996 B.n995 58.2333
R1520 B.n995 B.n23 58.2333
R1521 B.n989 B.n23 58.2333
R1522 B.n989 B.n988 58.2333
R1523 B.n988 B.n987 58.2333
R1524 B.n987 B.n30 58.2333
R1525 B.n981 B.n980 58.2333
R1526 B.n980 B.n979 58.2333
R1527 B.n979 B.n37 58.2333
R1528 B.n973 B.n37 58.2333
R1529 B.n973 B.n972 58.2333
R1530 B.n972 B.n971 58.2333
R1531 B.n971 B.n44 58.2333
R1532 B.n965 B.n44 58.2333
R1533 B.n965 B.n964 58.2333
R1534 B.n963 B.n51 58.2333
R1535 B.n957 B.n51 58.2333
R1536 B.n957 B.n956 58.2333
R1537 B.n956 B.n955 58.2333
R1538 B.n955 B.n58 58.2333
R1539 B.n949 B.n58 58.2333
R1540 B.n949 B.n948 58.2333
R1541 B.n948 B.n947 58.2333
R1542 B.n947 B.n65 58.2333
R1543 B.n941 B.n940 58.2333
R1544 B.n940 B.n939 58.2333
R1545 B.n939 B.n72 58.2333
R1546 B.n933 B.n72 58.2333
R1547 B.n933 B.n932 58.2333
R1548 B.n932 B.n931 58.2333
R1549 B.n931 B.n79 58.2333
R1550 B.n925 B.n79 58.2333
R1551 B.n925 B.n924 58.2333
R1552 B.n923 B.n86 58.2333
R1553 B.n917 B.n86 58.2333
R1554 B.n917 B.n916 58.2333
R1555 B.n916 B.n915 58.2333
R1556 B.n915 B.n93 58.2333
R1557 B.n909 B.n93 58.2333
R1558 B.n909 B.n908 58.2333
R1559 B.n908 B.n907 58.2333
R1560 B.n907 B.n100 58.2333
R1561 B.n901 B.n100 58.2333
R1562 B.n901 B.n900 58.2333
R1563 B.n900 B.n899 58.2333
R1564 B.n893 B.n110 58.2333
R1565 B.n893 B.n892 58.2333
R1566 B.n892 B.n891 58.2333
R1567 B.n891 B.n114 58.2333
R1568 B.n885 B.n114 58.2333
R1569 B.n885 B.n884 58.2333
R1570 B.n884 B.n883 58.2333
R1571 B.n482 B.t11 57.3769
R1572 B.t7 B.n167 57.3769
R1573 B.n1004 B.t9 57.3769
R1574 B.n110 B.t15 57.3769
R1575 B.n525 B.t0 55.6642
R1576 B.t4 B.n923 55.6642
R1577 B.t1 B.n187 43.6751
R1578 B.t8 B.n30 43.6751
R1579 B.n555 B.t5 41.9624
R1580 B.n941 B.t3 41.9624
R1581 B.n462 B.n461 33.2493
R1582 B.n466 B.n288 33.2493
R1583 B.n747 B.n746 33.2493
R1584 B.n881 B.n880 33.2493
R1585 B.t6 B.n207 29.9733
R1586 B.n964 B.t2 29.9733
R1587 B.n585 B.t6 28.2605
R1588 B.t2 B.n963 28.2605
R1589 B B.n1017 18.0485
R1590 B.t5 B.n227 16.2714
R1591 B.t3 B.n65 16.2714
R1592 B.n615 B.t1 14.5587
R1593 B.n981 B.t8 14.5587
R1594 B.n462 B.n284 10.6151
R1595 B.n472 B.n284 10.6151
R1596 B.n473 B.n472 10.6151
R1597 B.n474 B.n473 10.6151
R1598 B.n474 B.n276 10.6151
R1599 B.n485 B.n276 10.6151
R1600 B.n486 B.n485 10.6151
R1601 B.n487 B.n486 10.6151
R1602 B.n487 B.n269 10.6151
R1603 B.n497 B.n269 10.6151
R1604 B.n498 B.n497 10.6151
R1605 B.n499 B.n498 10.6151
R1606 B.n499 B.n261 10.6151
R1607 B.n509 B.n261 10.6151
R1608 B.n510 B.n509 10.6151
R1609 B.n511 B.n510 10.6151
R1610 B.n511 B.n253 10.6151
R1611 B.n521 B.n253 10.6151
R1612 B.n522 B.n521 10.6151
R1613 B.n523 B.n522 10.6151
R1614 B.n523 B.n245 10.6151
R1615 B.n533 B.n245 10.6151
R1616 B.n534 B.n533 10.6151
R1617 B.n535 B.n534 10.6151
R1618 B.n535 B.n237 10.6151
R1619 B.n545 B.n237 10.6151
R1620 B.n546 B.n545 10.6151
R1621 B.n547 B.n546 10.6151
R1622 B.n547 B.n229 10.6151
R1623 B.n557 B.n229 10.6151
R1624 B.n558 B.n557 10.6151
R1625 B.n559 B.n558 10.6151
R1626 B.n559 B.n221 10.6151
R1627 B.n569 B.n221 10.6151
R1628 B.n570 B.n569 10.6151
R1629 B.n571 B.n570 10.6151
R1630 B.n571 B.n213 10.6151
R1631 B.n581 B.n213 10.6151
R1632 B.n582 B.n581 10.6151
R1633 B.n583 B.n582 10.6151
R1634 B.n583 B.n205 10.6151
R1635 B.n593 B.n205 10.6151
R1636 B.n594 B.n593 10.6151
R1637 B.n595 B.n594 10.6151
R1638 B.n595 B.n197 10.6151
R1639 B.n605 B.n197 10.6151
R1640 B.n606 B.n605 10.6151
R1641 B.n607 B.n606 10.6151
R1642 B.n607 B.n189 10.6151
R1643 B.n617 B.n189 10.6151
R1644 B.n618 B.n617 10.6151
R1645 B.n619 B.n618 10.6151
R1646 B.n619 B.n181 10.6151
R1647 B.n629 B.n181 10.6151
R1648 B.n630 B.n629 10.6151
R1649 B.n631 B.n630 10.6151
R1650 B.n631 B.n173 10.6151
R1651 B.n641 B.n173 10.6151
R1652 B.n642 B.n641 10.6151
R1653 B.n643 B.n642 10.6151
R1654 B.n643 B.n165 10.6151
R1655 B.n654 B.n165 10.6151
R1656 B.n655 B.n654 10.6151
R1657 B.n656 B.n655 10.6151
R1658 B.n656 B.n0 10.6151
R1659 B.n461 B.n460 10.6151
R1660 B.n460 B.n292 10.6151
R1661 B.n455 B.n292 10.6151
R1662 B.n455 B.n454 10.6151
R1663 B.n454 B.n294 10.6151
R1664 B.n449 B.n294 10.6151
R1665 B.n449 B.n448 10.6151
R1666 B.n448 B.n447 10.6151
R1667 B.n447 B.n296 10.6151
R1668 B.n441 B.n296 10.6151
R1669 B.n441 B.n440 10.6151
R1670 B.n440 B.n439 10.6151
R1671 B.n439 B.n298 10.6151
R1672 B.n433 B.n298 10.6151
R1673 B.n433 B.n432 10.6151
R1674 B.n432 B.n431 10.6151
R1675 B.n431 B.n300 10.6151
R1676 B.n425 B.n300 10.6151
R1677 B.n425 B.n424 10.6151
R1678 B.n424 B.n423 10.6151
R1679 B.n423 B.n302 10.6151
R1680 B.n417 B.n302 10.6151
R1681 B.n417 B.n416 10.6151
R1682 B.n416 B.n415 10.6151
R1683 B.n415 B.n304 10.6151
R1684 B.n409 B.n304 10.6151
R1685 B.n409 B.n408 10.6151
R1686 B.n408 B.n407 10.6151
R1687 B.n403 B.n402 10.6151
R1688 B.n402 B.n310 10.6151
R1689 B.n397 B.n310 10.6151
R1690 B.n397 B.n396 10.6151
R1691 B.n396 B.n395 10.6151
R1692 B.n395 B.n312 10.6151
R1693 B.n389 B.n312 10.6151
R1694 B.n389 B.n388 10.6151
R1695 B.n386 B.n316 10.6151
R1696 B.n380 B.n316 10.6151
R1697 B.n380 B.n379 10.6151
R1698 B.n379 B.n378 10.6151
R1699 B.n378 B.n318 10.6151
R1700 B.n372 B.n318 10.6151
R1701 B.n372 B.n371 10.6151
R1702 B.n371 B.n370 10.6151
R1703 B.n370 B.n320 10.6151
R1704 B.n364 B.n320 10.6151
R1705 B.n364 B.n363 10.6151
R1706 B.n363 B.n362 10.6151
R1707 B.n362 B.n322 10.6151
R1708 B.n356 B.n322 10.6151
R1709 B.n356 B.n355 10.6151
R1710 B.n355 B.n354 10.6151
R1711 B.n354 B.n324 10.6151
R1712 B.n348 B.n324 10.6151
R1713 B.n348 B.n347 10.6151
R1714 B.n347 B.n346 10.6151
R1715 B.n346 B.n326 10.6151
R1716 B.n340 B.n326 10.6151
R1717 B.n340 B.n339 10.6151
R1718 B.n339 B.n338 10.6151
R1719 B.n338 B.n328 10.6151
R1720 B.n332 B.n328 10.6151
R1721 B.n332 B.n331 10.6151
R1722 B.n331 B.n288 10.6151
R1723 B.n467 B.n466 10.6151
R1724 B.n468 B.n467 10.6151
R1725 B.n468 B.n280 10.6151
R1726 B.n478 B.n280 10.6151
R1727 B.n479 B.n478 10.6151
R1728 B.n480 B.n479 10.6151
R1729 B.n480 B.n273 10.6151
R1730 B.n491 B.n273 10.6151
R1731 B.n492 B.n491 10.6151
R1732 B.n493 B.n492 10.6151
R1733 B.n493 B.n265 10.6151
R1734 B.n503 B.n265 10.6151
R1735 B.n504 B.n503 10.6151
R1736 B.n505 B.n504 10.6151
R1737 B.n505 B.n257 10.6151
R1738 B.n515 B.n257 10.6151
R1739 B.n516 B.n515 10.6151
R1740 B.n517 B.n516 10.6151
R1741 B.n517 B.n249 10.6151
R1742 B.n527 B.n249 10.6151
R1743 B.n528 B.n527 10.6151
R1744 B.n529 B.n528 10.6151
R1745 B.n529 B.n241 10.6151
R1746 B.n539 B.n241 10.6151
R1747 B.n540 B.n539 10.6151
R1748 B.n541 B.n540 10.6151
R1749 B.n541 B.n233 10.6151
R1750 B.n551 B.n233 10.6151
R1751 B.n552 B.n551 10.6151
R1752 B.n553 B.n552 10.6151
R1753 B.n553 B.n225 10.6151
R1754 B.n563 B.n225 10.6151
R1755 B.n564 B.n563 10.6151
R1756 B.n565 B.n564 10.6151
R1757 B.n565 B.n217 10.6151
R1758 B.n575 B.n217 10.6151
R1759 B.n576 B.n575 10.6151
R1760 B.n577 B.n576 10.6151
R1761 B.n577 B.n209 10.6151
R1762 B.n587 B.n209 10.6151
R1763 B.n588 B.n587 10.6151
R1764 B.n589 B.n588 10.6151
R1765 B.n589 B.n201 10.6151
R1766 B.n599 B.n201 10.6151
R1767 B.n600 B.n599 10.6151
R1768 B.n601 B.n600 10.6151
R1769 B.n601 B.n193 10.6151
R1770 B.n611 B.n193 10.6151
R1771 B.n612 B.n611 10.6151
R1772 B.n613 B.n612 10.6151
R1773 B.n613 B.n185 10.6151
R1774 B.n623 B.n185 10.6151
R1775 B.n624 B.n623 10.6151
R1776 B.n625 B.n624 10.6151
R1777 B.n625 B.n177 10.6151
R1778 B.n635 B.n177 10.6151
R1779 B.n636 B.n635 10.6151
R1780 B.n637 B.n636 10.6151
R1781 B.n637 B.n169 10.6151
R1782 B.n647 B.n169 10.6151
R1783 B.n648 B.n647 10.6151
R1784 B.n650 B.n648 10.6151
R1785 B.n650 B.n649 10.6151
R1786 B.n649 B.n161 10.6151
R1787 B.n661 B.n161 10.6151
R1788 B.n662 B.n661 10.6151
R1789 B.n663 B.n662 10.6151
R1790 B.n664 B.n663 10.6151
R1791 B.n665 B.n664 10.6151
R1792 B.n668 B.n665 10.6151
R1793 B.n669 B.n668 10.6151
R1794 B.n670 B.n669 10.6151
R1795 B.n671 B.n670 10.6151
R1796 B.n673 B.n671 10.6151
R1797 B.n674 B.n673 10.6151
R1798 B.n675 B.n674 10.6151
R1799 B.n676 B.n675 10.6151
R1800 B.n678 B.n676 10.6151
R1801 B.n679 B.n678 10.6151
R1802 B.n680 B.n679 10.6151
R1803 B.n681 B.n680 10.6151
R1804 B.n683 B.n681 10.6151
R1805 B.n684 B.n683 10.6151
R1806 B.n685 B.n684 10.6151
R1807 B.n686 B.n685 10.6151
R1808 B.n688 B.n686 10.6151
R1809 B.n689 B.n688 10.6151
R1810 B.n690 B.n689 10.6151
R1811 B.n691 B.n690 10.6151
R1812 B.n693 B.n691 10.6151
R1813 B.n694 B.n693 10.6151
R1814 B.n695 B.n694 10.6151
R1815 B.n696 B.n695 10.6151
R1816 B.n698 B.n696 10.6151
R1817 B.n699 B.n698 10.6151
R1818 B.n700 B.n699 10.6151
R1819 B.n701 B.n700 10.6151
R1820 B.n703 B.n701 10.6151
R1821 B.n704 B.n703 10.6151
R1822 B.n705 B.n704 10.6151
R1823 B.n706 B.n705 10.6151
R1824 B.n708 B.n706 10.6151
R1825 B.n709 B.n708 10.6151
R1826 B.n710 B.n709 10.6151
R1827 B.n711 B.n710 10.6151
R1828 B.n713 B.n711 10.6151
R1829 B.n714 B.n713 10.6151
R1830 B.n715 B.n714 10.6151
R1831 B.n716 B.n715 10.6151
R1832 B.n718 B.n716 10.6151
R1833 B.n719 B.n718 10.6151
R1834 B.n720 B.n719 10.6151
R1835 B.n721 B.n720 10.6151
R1836 B.n723 B.n721 10.6151
R1837 B.n724 B.n723 10.6151
R1838 B.n725 B.n724 10.6151
R1839 B.n726 B.n725 10.6151
R1840 B.n728 B.n726 10.6151
R1841 B.n729 B.n728 10.6151
R1842 B.n730 B.n729 10.6151
R1843 B.n731 B.n730 10.6151
R1844 B.n733 B.n731 10.6151
R1845 B.n734 B.n733 10.6151
R1846 B.n735 B.n734 10.6151
R1847 B.n736 B.n735 10.6151
R1848 B.n738 B.n736 10.6151
R1849 B.n739 B.n738 10.6151
R1850 B.n740 B.n739 10.6151
R1851 B.n741 B.n740 10.6151
R1852 B.n743 B.n741 10.6151
R1853 B.n744 B.n743 10.6151
R1854 B.n745 B.n744 10.6151
R1855 B.n746 B.n745 10.6151
R1856 B.n1009 B.n1 10.6151
R1857 B.n1009 B.n1008 10.6151
R1858 B.n1008 B.n1007 10.6151
R1859 B.n1007 B.n10 10.6151
R1860 B.n1001 B.n10 10.6151
R1861 B.n1001 B.n1000 10.6151
R1862 B.n1000 B.n999 10.6151
R1863 B.n999 B.n18 10.6151
R1864 B.n993 B.n18 10.6151
R1865 B.n993 B.n992 10.6151
R1866 B.n992 B.n991 10.6151
R1867 B.n991 B.n25 10.6151
R1868 B.n985 B.n25 10.6151
R1869 B.n985 B.n984 10.6151
R1870 B.n984 B.n983 10.6151
R1871 B.n983 B.n32 10.6151
R1872 B.n977 B.n32 10.6151
R1873 B.n977 B.n976 10.6151
R1874 B.n976 B.n975 10.6151
R1875 B.n975 B.n39 10.6151
R1876 B.n969 B.n39 10.6151
R1877 B.n969 B.n968 10.6151
R1878 B.n968 B.n967 10.6151
R1879 B.n967 B.n46 10.6151
R1880 B.n961 B.n46 10.6151
R1881 B.n961 B.n960 10.6151
R1882 B.n960 B.n959 10.6151
R1883 B.n959 B.n53 10.6151
R1884 B.n953 B.n53 10.6151
R1885 B.n953 B.n952 10.6151
R1886 B.n952 B.n951 10.6151
R1887 B.n951 B.n60 10.6151
R1888 B.n945 B.n60 10.6151
R1889 B.n945 B.n944 10.6151
R1890 B.n944 B.n943 10.6151
R1891 B.n943 B.n67 10.6151
R1892 B.n937 B.n67 10.6151
R1893 B.n937 B.n936 10.6151
R1894 B.n936 B.n935 10.6151
R1895 B.n935 B.n74 10.6151
R1896 B.n929 B.n74 10.6151
R1897 B.n929 B.n928 10.6151
R1898 B.n928 B.n927 10.6151
R1899 B.n927 B.n81 10.6151
R1900 B.n921 B.n81 10.6151
R1901 B.n921 B.n920 10.6151
R1902 B.n920 B.n919 10.6151
R1903 B.n919 B.n88 10.6151
R1904 B.n913 B.n88 10.6151
R1905 B.n913 B.n912 10.6151
R1906 B.n912 B.n911 10.6151
R1907 B.n911 B.n95 10.6151
R1908 B.n905 B.n95 10.6151
R1909 B.n905 B.n904 10.6151
R1910 B.n904 B.n903 10.6151
R1911 B.n903 B.n102 10.6151
R1912 B.n897 B.n102 10.6151
R1913 B.n897 B.n896 10.6151
R1914 B.n896 B.n895 10.6151
R1915 B.n895 B.n108 10.6151
R1916 B.n889 B.n108 10.6151
R1917 B.n889 B.n888 10.6151
R1918 B.n888 B.n887 10.6151
R1919 B.n887 B.n116 10.6151
R1920 B.n881 B.n116 10.6151
R1921 B.n880 B.n879 10.6151
R1922 B.n879 B.n123 10.6151
R1923 B.n873 B.n123 10.6151
R1924 B.n873 B.n872 10.6151
R1925 B.n872 B.n871 10.6151
R1926 B.n871 B.n125 10.6151
R1927 B.n865 B.n125 10.6151
R1928 B.n865 B.n864 10.6151
R1929 B.n864 B.n863 10.6151
R1930 B.n863 B.n127 10.6151
R1931 B.n857 B.n127 10.6151
R1932 B.n857 B.n856 10.6151
R1933 B.n856 B.n855 10.6151
R1934 B.n855 B.n129 10.6151
R1935 B.n849 B.n129 10.6151
R1936 B.n849 B.n848 10.6151
R1937 B.n848 B.n847 10.6151
R1938 B.n847 B.n131 10.6151
R1939 B.n841 B.n131 10.6151
R1940 B.n841 B.n840 10.6151
R1941 B.n840 B.n839 10.6151
R1942 B.n839 B.n133 10.6151
R1943 B.n833 B.n133 10.6151
R1944 B.n833 B.n832 10.6151
R1945 B.n832 B.n831 10.6151
R1946 B.n831 B.n135 10.6151
R1947 B.n825 B.n135 10.6151
R1948 B.n825 B.n824 10.6151
R1949 B.n822 B.n139 10.6151
R1950 B.n816 B.n139 10.6151
R1951 B.n816 B.n815 10.6151
R1952 B.n815 B.n814 10.6151
R1953 B.n814 B.n141 10.6151
R1954 B.n808 B.n141 10.6151
R1955 B.n808 B.n807 10.6151
R1956 B.n807 B.n806 10.6151
R1957 B.n802 B.n801 10.6151
R1958 B.n801 B.n147 10.6151
R1959 B.n796 B.n147 10.6151
R1960 B.n796 B.n795 10.6151
R1961 B.n795 B.n794 10.6151
R1962 B.n794 B.n149 10.6151
R1963 B.n788 B.n149 10.6151
R1964 B.n788 B.n787 10.6151
R1965 B.n787 B.n786 10.6151
R1966 B.n786 B.n151 10.6151
R1967 B.n780 B.n151 10.6151
R1968 B.n780 B.n779 10.6151
R1969 B.n779 B.n778 10.6151
R1970 B.n778 B.n153 10.6151
R1971 B.n772 B.n153 10.6151
R1972 B.n772 B.n771 10.6151
R1973 B.n771 B.n770 10.6151
R1974 B.n770 B.n155 10.6151
R1975 B.n764 B.n155 10.6151
R1976 B.n764 B.n763 10.6151
R1977 B.n763 B.n762 10.6151
R1978 B.n762 B.n157 10.6151
R1979 B.n756 B.n157 10.6151
R1980 B.n756 B.n755 10.6151
R1981 B.n755 B.n754 10.6151
R1982 B.n754 B.n159 10.6151
R1983 B.n748 B.n159 10.6151
R1984 B.n748 B.n747 10.6151
R1985 B.n1017 B.n0 8.11757
R1986 B.n1017 B.n1 8.11757
R1987 B.n403 B.n308 6.5566
R1988 B.n388 B.n387 6.5566
R1989 B.n823 B.n822 6.5566
R1990 B.n806 B.n145 6.5566
R1991 B.n407 B.n308 4.05904
R1992 B.n387 B.n386 4.05904
R1993 B.n824 B.n823 4.05904
R1994 B.n802 B.n145 4.05904
R1995 B.t0 B.n247 2.56959
R1996 B.n924 B.t4 2.56959
R1997 B.n489 B.t11 0.856864
R1998 B.n645 B.t7 0.856864
R1999 B.t9 B.n1003 0.856864
R2000 B.n899 B.t15 0.856864
R2001 VN.n90 VN.n89 161.3
R2002 VN.n88 VN.n47 161.3
R2003 VN.n87 VN.n86 161.3
R2004 VN.n85 VN.n48 161.3
R2005 VN.n84 VN.n83 161.3
R2006 VN.n82 VN.n49 161.3
R2007 VN.n80 VN.n79 161.3
R2008 VN.n78 VN.n50 161.3
R2009 VN.n77 VN.n76 161.3
R2010 VN.n75 VN.n51 161.3
R2011 VN.n74 VN.n73 161.3
R2012 VN.n72 VN.n52 161.3
R2013 VN.n71 VN.n70 161.3
R2014 VN.n68 VN.n53 161.3
R2015 VN.n67 VN.n66 161.3
R2016 VN.n65 VN.n54 161.3
R2017 VN.n64 VN.n63 161.3
R2018 VN.n62 VN.n55 161.3
R2019 VN.n61 VN.n60 161.3
R2020 VN.n59 VN.n56 161.3
R2021 VN.n44 VN.n43 161.3
R2022 VN.n42 VN.n1 161.3
R2023 VN.n41 VN.n40 161.3
R2024 VN.n39 VN.n2 161.3
R2025 VN.n38 VN.n37 161.3
R2026 VN.n36 VN.n3 161.3
R2027 VN.n34 VN.n33 161.3
R2028 VN.n32 VN.n4 161.3
R2029 VN.n31 VN.n30 161.3
R2030 VN.n29 VN.n5 161.3
R2031 VN.n28 VN.n27 161.3
R2032 VN.n26 VN.n6 161.3
R2033 VN.n25 VN.n24 161.3
R2034 VN.n22 VN.n7 161.3
R2035 VN.n21 VN.n20 161.3
R2036 VN.n19 VN.n8 161.3
R2037 VN.n18 VN.n17 161.3
R2038 VN.n16 VN.n9 161.3
R2039 VN.n15 VN.n14 161.3
R2040 VN.n13 VN.n10 161.3
R2041 VN.n58 VN.t6 92.6708
R2042 VN.n12 VN.t3 92.6708
R2043 VN.n45 VN.n0 70.9831
R2044 VN.n91 VN.n46 70.9831
R2045 VN.n12 VN.n11 70.1651
R2046 VN.n58 VN.n57 70.1651
R2047 VN.n11 VN.t1 61.0162
R2048 VN.n23 VN.t9 61.0162
R2049 VN.n35 VN.t8 61.0162
R2050 VN.n0 VN.t4 61.0162
R2051 VN.n57 VN.t2 61.0162
R2052 VN.n69 VN.t7 61.0162
R2053 VN.n81 VN.t0 61.0162
R2054 VN.n46 VN.t5 61.0162
R2055 VN.n41 VN.n2 56.5193
R2056 VN.n87 VN.n48 56.5193
R2057 VN VN.n91 52.1495
R2058 VN.n17 VN.n8 49.2348
R2059 VN.n29 VN.n28 49.2348
R2060 VN.n63 VN.n54 49.2348
R2061 VN.n75 VN.n74 49.2348
R2062 VN.n17 VN.n16 31.752
R2063 VN.n30 VN.n29 31.752
R2064 VN.n63 VN.n62 31.752
R2065 VN.n76 VN.n75 31.752
R2066 VN.n15 VN.n10 24.4675
R2067 VN.n16 VN.n15 24.4675
R2068 VN.n21 VN.n8 24.4675
R2069 VN.n22 VN.n21 24.4675
R2070 VN.n24 VN.n6 24.4675
R2071 VN.n28 VN.n6 24.4675
R2072 VN.n30 VN.n4 24.4675
R2073 VN.n34 VN.n4 24.4675
R2074 VN.n37 VN.n36 24.4675
R2075 VN.n37 VN.n2 24.4675
R2076 VN.n42 VN.n41 24.4675
R2077 VN.n43 VN.n42 24.4675
R2078 VN.n62 VN.n61 24.4675
R2079 VN.n61 VN.n56 24.4675
R2080 VN.n74 VN.n52 24.4675
R2081 VN.n70 VN.n52 24.4675
R2082 VN.n68 VN.n67 24.4675
R2083 VN.n67 VN.n54 24.4675
R2084 VN.n83 VN.n48 24.4675
R2085 VN.n83 VN.n82 24.4675
R2086 VN.n80 VN.n50 24.4675
R2087 VN.n76 VN.n50 24.4675
R2088 VN.n89 VN.n88 24.4675
R2089 VN.n88 VN.n87 24.4675
R2090 VN.n36 VN.n35 21.0421
R2091 VN.n82 VN.n81 21.0421
R2092 VN.n43 VN.n0 19.0848
R2093 VN.n89 VN.n46 19.0848
R2094 VN.n23 VN.n22 12.234
R2095 VN.n24 VN.n23 12.234
R2096 VN.n70 VN.n69 12.234
R2097 VN.n69 VN.n68 12.234
R2098 VN.n59 VN.n58 5.61943
R2099 VN.n13 VN.n12 5.61943
R2100 VN.n11 VN.n10 3.42588
R2101 VN.n35 VN.n34 3.42588
R2102 VN.n57 VN.n56 3.42588
R2103 VN.n81 VN.n80 3.42588
R2104 VN.n91 VN.n90 0.354971
R2105 VN.n45 VN.n44 0.354971
R2106 VN VN.n45 0.26696
R2107 VN.n90 VN.n47 0.189894
R2108 VN.n86 VN.n47 0.189894
R2109 VN.n86 VN.n85 0.189894
R2110 VN.n85 VN.n84 0.189894
R2111 VN.n84 VN.n49 0.189894
R2112 VN.n79 VN.n49 0.189894
R2113 VN.n79 VN.n78 0.189894
R2114 VN.n78 VN.n77 0.189894
R2115 VN.n77 VN.n51 0.189894
R2116 VN.n73 VN.n51 0.189894
R2117 VN.n73 VN.n72 0.189894
R2118 VN.n72 VN.n71 0.189894
R2119 VN.n71 VN.n53 0.189894
R2120 VN.n66 VN.n53 0.189894
R2121 VN.n66 VN.n65 0.189894
R2122 VN.n65 VN.n64 0.189894
R2123 VN.n64 VN.n55 0.189894
R2124 VN.n60 VN.n55 0.189894
R2125 VN.n60 VN.n59 0.189894
R2126 VN.n14 VN.n13 0.189894
R2127 VN.n14 VN.n9 0.189894
R2128 VN.n18 VN.n9 0.189894
R2129 VN.n19 VN.n18 0.189894
R2130 VN.n20 VN.n19 0.189894
R2131 VN.n20 VN.n7 0.189894
R2132 VN.n25 VN.n7 0.189894
R2133 VN.n26 VN.n25 0.189894
R2134 VN.n27 VN.n26 0.189894
R2135 VN.n27 VN.n5 0.189894
R2136 VN.n31 VN.n5 0.189894
R2137 VN.n32 VN.n31 0.189894
R2138 VN.n33 VN.n32 0.189894
R2139 VN.n33 VN.n3 0.189894
R2140 VN.n38 VN.n3 0.189894
R2141 VN.n39 VN.n38 0.189894
R2142 VN.n40 VN.n39 0.189894
R2143 VN.n40 VN.n1 0.189894
R2144 VN.n44 VN.n1 0.189894
R2145 VDD2.n1 VDD2.t6 72.29
R2146 VDD2.n4 VDD2.t4 69.4281
R2147 VDD2.n3 VDD2.n2 68.9035
R2148 VDD2 VDD2.n7 68.9007
R2149 VDD2.n6 VDD2.n5 66.8125
R2150 VDD2.n1 VDD2.n0 66.8123
R2151 VDD2.n4 VDD2.n3 43.836
R2152 VDD2.n6 VDD2.n4 2.86257
R2153 VDD2.n7 VDD2.t7 2.61609
R2154 VDD2.n7 VDD2.t3 2.61609
R2155 VDD2.n5 VDD2.t9 2.61609
R2156 VDD2.n5 VDD2.t2 2.61609
R2157 VDD2.n2 VDD2.t1 2.61609
R2158 VDD2.n2 VDD2.t5 2.61609
R2159 VDD2.n0 VDD2.t8 2.61609
R2160 VDD2.n0 VDD2.t0 2.61609
R2161 VDD2 VDD2.n6 0.774207
R2162 VDD2.n3 VDD2.n1 0.660671
C0 VTAIL VDD2 8.66535f
C1 VDD2 VDD1 2.4281f
C2 VTAIL VN 8.113529f
C3 VN VDD1 0.154276f
C4 VTAIL VDD1 8.61051f
C5 VDD2 VP 0.63304f
C6 VN VP 8.15609f
C7 VN VDD2 7.10054f
C8 VTAIL VP 8.12773f
C9 VDD1 VP 7.576129f
C10 VDD2 B 6.921974f
C11 VDD1 B 6.865047f
C12 VTAIL B 6.745031f
C13 VN B 19.688461f
C14 VP B 18.268923f
C15 VDD2.t6 B 1.70539f
C16 VDD2.t8 B 0.153767f
C17 VDD2.t0 B 0.153767f
C18 VDD2.n0 B 1.32578f
C19 VDD2.n1 B 0.985276f
C20 VDD2.t1 B 0.153767f
C21 VDD2.t5 B 0.153767f
C22 VDD2.n2 B 1.34471f
C23 VDD2.n3 B 2.90937f
C24 VDD2.t4 B 1.6852f
C25 VDD2.n4 B 2.99853f
C26 VDD2.t9 B 0.153767f
C27 VDD2.t2 B 0.153767f
C28 VDD2.n5 B 1.32579f
C29 VDD2.n6 B 0.503872f
C30 VDD2.t7 B 0.153767f
C31 VDD2.t3 B 0.153767f
C32 VDD2.n7 B 1.34467f
C33 VN.t4 B 1.27732f
C34 VN.n0 B 0.54643f
C35 VN.n1 B 0.021064f
C36 VN.n2 B 0.029576f
C37 VN.n3 B 0.021064f
C38 VN.t8 B 1.27732f
C39 VN.n4 B 0.039259f
C40 VN.n5 B 0.021064f
C41 VN.n6 B 0.039259f
C42 VN.n7 B 0.021064f
C43 VN.t9 B 1.27732f
C44 VN.n8 B 0.039062f
C45 VN.n9 B 0.021064f
C46 VN.n10 B 0.02259f
C47 VN.t1 B 1.27732f
C48 VN.n11 B 0.525018f
C49 VN.t3 B 1.48379f
C50 VN.n12 B 0.508993f
C51 VN.n13 B 0.227878f
C52 VN.n14 B 0.021064f
C53 VN.n15 B 0.039259f
C54 VN.n16 B 0.04237f
C55 VN.n17 B 0.019327f
C56 VN.n18 B 0.021064f
C57 VN.n19 B 0.021064f
C58 VN.n20 B 0.021064f
C59 VN.n21 B 0.039259f
C60 VN.n22 B 0.029568f
C61 VN.n23 B 0.464767f
C62 VN.n24 B 0.029568f
C63 VN.n25 B 0.021064f
C64 VN.n26 B 0.021064f
C65 VN.n27 B 0.021064f
C66 VN.n28 B 0.039062f
C67 VN.n29 B 0.019327f
C68 VN.n30 B 0.04237f
C69 VN.n31 B 0.021064f
C70 VN.n32 B 0.021064f
C71 VN.n33 B 0.021064f
C72 VN.n34 B 0.02259f
C73 VN.n35 B 0.464767f
C74 VN.n36 B 0.036545f
C75 VN.n37 B 0.039259f
C76 VN.n38 B 0.021064f
C77 VN.n39 B 0.021064f
C78 VN.n40 B 0.021064f
C79 VN.n41 B 0.031924f
C80 VN.n42 B 0.039259f
C81 VN.n43 B 0.034995f
C82 VN.n44 B 0.033998f
C83 VN.n45 B 0.044623f
C84 VN.t5 B 1.27732f
C85 VN.n46 B 0.54643f
C86 VN.n47 B 0.021064f
C87 VN.n48 B 0.029576f
C88 VN.n49 B 0.021064f
C89 VN.t0 B 1.27732f
C90 VN.n50 B 0.039259f
C91 VN.n51 B 0.021064f
C92 VN.n52 B 0.039259f
C93 VN.n53 B 0.021064f
C94 VN.t7 B 1.27732f
C95 VN.n54 B 0.039062f
C96 VN.n55 B 0.021064f
C97 VN.n56 B 0.02259f
C98 VN.t6 B 1.48379f
C99 VN.t2 B 1.27732f
C100 VN.n57 B 0.525018f
C101 VN.n58 B 0.508993f
C102 VN.n59 B 0.227878f
C103 VN.n60 B 0.021064f
C104 VN.n61 B 0.039259f
C105 VN.n62 B 0.04237f
C106 VN.n63 B 0.019327f
C107 VN.n64 B 0.021064f
C108 VN.n65 B 0.021064f
C109 VN.n66 B 0.021064f
C110 VN.n67 B 0.039259f
C111 VN.n68 B 0.029568f
C112 VN.n69 B 0.464767f
C113 VN.n70 B 0.029568f
C114 VN.n71 B 0.021064f
C115 VN.n72 B 0.021064f
C116 VN.n73 B 0.021064f
C117 VN.n74 B 0.039062f
C118 VN.n75 B 0.019327f
C119 VN.n76 B 0.04237f
C120 VN.n77 B 0.021064f
C121 VN.n78 B 0.021064f
C122 VN.n79 B 0.021064f
C123 VN.n80 B 0.02259f
C124 VN.n81 B 0.464767f
C125 VN.n82 B 0.036545f
C126 VN.n83 B 0.039259f
C127 VN.n84 B 0.021064f
C128 VN.n85 B 0.021064f
C129 VN.n86 B 0.021064f
C130 VN.n87 B 0.031924f
C131 VN.n88 B 0.039259f
C132 VN.n89 B 0.034995f
C133 VN.n90 B 0.033998f
C134 VN.n91 B 1.26792f
C135 VDD1.t5 B 1.73383f
C136 VDD1.t0 B 0.156331f
C137 VDD1.t8 B 0.156331f
C138 VDD1.n0 B 1.34789f
C139 VDD1.n1 B 1.01034f
C140 VDD1.t9 B 1.73383f
C141 VDD1.t6 B 0.156331f
C142 VDD1.t7 B 0.156331f
C143 VDD1.n2 B 1.34789f
C144 VDD1.n3 B 1.0017f
C145 VDD1.t1 B 0.156331f
C146 VDD1.t3 B 0.156331f
C147 VDD1.n4 B 1.36713f
C148 VDD1.n5 B 3.09587f
C149 VDD1.t4 B 0.156331f
C150 VDD1.t2 B 0.156331f
C151 VDD1.n6 B 1.34789f
C152 VDD1.n7 B 3.12197f
C153 VTAIL.t9 B 0.163715f
C154 VTAIL.t8 B 0.163715f
C155 VTAIL.n0 B 1.34148f
C156 VTAIL.n1 B 0.610785f
C157 VTAIL.t11 B 1.70743f
C158 VTAIL.n2 B 0.749292f
C159 VTAIL.t16 B 0.163715f
C160 VTAIL.t15 B 0.163715f
C161 VTAIL.n3 B 1.34148f
C162 VTAIL.n4 B 0.753515f
C163 VTAIL.t10 B 0.163715f
C164 VTAIL.t14 B 0.163715f
C165 VTAIL.n5 B 1.34148f
C166 VTAIL.n6 B 1.95315f
C167 VTAIL.t0 B 0.163715f
C168 VTAIL.t5 B 0.163715f
C169 VTAIL.n7 B 1.34148f
C170 VTAIL.n8 B 1.95314f
C171 VTAIL.t6 B 0.163715f
C172 VTAIL.t1 B 0.163715f
C173 VTAIL.n9 B 1.34148f
C174 VTAIL.n10 B 0.753512f
C175 VTAIL.t7 B 1.70743f
C176 VTAIL.n11 B 0.749288f
C177 VTAIL.t12 B 0.163715f
C178 VTAIL.t13 B 0.163715f
C179 VTAIL.n12 B 1.34148f
C180 VTAIL.n13 B 0.668748f
C181 VTAIL.t18 B 0.163715f
C182 VTAIL.t17 B 0.163715f
C183 VTAIL.n14 B 1.34148f
C184 VTAIL.n15 B 0.753512f
C185 VTAIL.t19 B 1.70743f
C186 VTAIL.n16 B 1.7813f
C187 VTAIL.t4 B 1.70743f
C188 VTAIL.n17 B 1.7813f
C189 VTAIL.t2 B 0.163715f
C190 VTAIL.t3 B 0.163715f
C191 VTAIL.n18 B 1.34148f
C192 VTAIL.n19 B 0.559091f
C193 VP.t6 B 1.30626f
C194 VP.n0 B 0.558813f
C195 VP.n1 B 0.021542f
C196 VP.n2 B 0.030247f
C197 VP.n3 B 0.021542f
C198 VP.t8 B 1.30626f
C199 VP.n4 B 0.040148f
C200 VP.n5 B 0.021542f
C201 VP.n6 B 0.040148f
C202 VP.n7 B 0.021542f
C203 VP.t2 B 1.30626f
C204 VP.n8 B 0.039947f
C205 VP.n9 B 0.021542f
C206 VP.n10 B 0.023102f
C207 VP.n11 B 0.021542f
C208 VP.n12 B 0.032648f
C209 VP.n13 B 0.034768f
C210 VP.t0 B 1.30626f
C211 VP.t7 B 1.30626f
C212 VP.n14 B 0.558813f
C213 VP.n15 B 0.021542f
C214 VP.n16 B 0.030247f
C215 VP.n17 B 0.021542f
C216 VP.t5 B 1.30626f
C217 VP.n18 B 0.040148f
C218 VP.n19 B 0.021542f
C219 VP.n20 B 0.040148f
C220 VP.n21 B 0.021542f
C221 VP.t1 B 1.30626f
C222 VP.n22 B 0.039947f
C223 VP.n23 B 0.021542f
C224 VP.n24 B 0.023102f
C225 VP.t4 B 1.51742f
C226 VP.t9 B 1.30626f
C227 VP.n25 B 0.536916f
C228 VP.n26 B 0.520529f
C229 VP.n27 B 0.233043f
C230 VP.n28 B 0.021542f
C231 VP.n29 B 0.040148f
C232 VP.n30 B 0.04333f
C233 VP.n31 B 0.019765f
C234 VP.n32 B 0.021542f
C235 VP.n33 B 0.021542f
C236 VP.n34 B 0.021542f
C237 VP.n35 B 0.040148f
C238 VP.n36 B 0.030238f
C239 VP.n37 B 0.475299f
C240 VP.n38 B 0.030238f
C241 VP.n39 B 0.021542f
C242 VP.n40 B 0.021542f
C243 VP.n41 B 0.021542f
C244 VP.n42 B 0.039947f
C245 VP.n43 B 0.019765f
C246 VP.n44 B 0.04333f
C247 VP.n45 B 0.021542f
C248 VP.n46 B 0.021542f
C249 VP.n47 B 0.021542f
C250 VP.n48 B 0.023102f
C251 VP.n49 B 0.475299f
C252 VP.n50 B 0.037373f
C253 VP.n51 B 0.040148f
C254 VP.n52 B 0.021542f
C255 VP.n53 B 0.021542f
C256 VP.n54 B 0.021542f
C257 VP.n55 B 0.032648f
C258 VP.n56 B 0.040148f
C259 VP.n57 B 0.035788f
C260 VP.n58 B 0.034768f
C261 VP.n59 B 1.28795f
C262 VP.n60 B 1.30285f
C263 VP.n61 B 0.558813f
C264 VP.n62 B 0.035788f
C265 VP.n63 B 0.040148f
C266 VP.n64 B 0.021542f
C267 VP.n65 B 0.021542f
C268 VP.n66 B 0.021542f
C269 VP.n67 B 0.030247f
C270 VP.n68 B 0.040148f
C271 VP.t3 B 1.30626f
C272 VP.n69 B 0.475299f
C273 VP.n70 B 0.037373f
C274 VP.n71 B 0.021542f
C275 VP.n72 B 0.021542f
C276 VP.n73 B 0.021542f
C277 VP.n74 B 0.040148f
C278 VP.n75 B 0.04333f
C279 VP.n76 B 0.019765f
C280 VP.n77 B 0.021542f
C281 VP.n78 B 0.021542f
C282 VP.n79 B 0.021542f
C283 VP.n80 B 0.040148f
C284 VP.n81 B 0.030238f
C285 VP.n82 B 0.475299f
C286 VP.n83 B 0.030238f
C287 VP.n84 B 0.021542f
C288 VP.n85 B 0.021542f
C289 VP.n86 B 0.021542f
C290 VP.n87 B 0.039947f
C291 VP.n88 B 0.019765f
C292 VP.n89 B 0.04333f
C293 VP.n90 B 0.021542f
C294 VP.n91 B 0.021542f
C295 VP.n92 B 0.021542f
C296 VP.n93 B 0.023102f
C297 VP.n94 B 0.475299f
C298 VP.n95 B 0.037373f
C299 VP.n96 B 0.040148f
C300 VP.n97 B 0.021542f
C301 VP.n98 B 0.021542f
C302 VP.n99 B 0.021542f
C303 VP.n100 B 0.032648f
C304 VP.n101 B 0.040148f
C305 VP.n102 B 0.035788f
C306 VP.n103 B 0.034768f
C307 VP.n104 B 0.045635f
.ends

