* NGSPICE file created from diff_pair_sample_0443.ext - technology: sky130A

.subckt diff_pair_sample_0443 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=0 ps=0 w=17.6 l=0.27
X1 VTAIL.t7 VN.t0 VDD2.t2 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=2.904 ps=17.93 w=17.6 l=0.27
X2 VTAIL.t6 VN.t1 VDD2.t1 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=2.904 ps=17.93 w=17.6 l=0.27
X3 B.t8 B.t6 B.t7 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=0 ps=0 w=17.6 l=0.27
X4 VDD1.t3 VP.t0 VTAIL.t2 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=2.904 pd=17.93 as=6.864 ps=35.98 w=17.6 l=0.27
X5 VTAIL.t3 VP.t1 VDD1.t2 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=2.904 ps=17.93 w=17.6 l=0.27
X6 B.t5 B.t3 B.t4 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=0 ps=0 w=17.6 l=0.27
X7 B.t2 B.t0 B.t1 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=0 ps=0 w=17.6 l=0.27
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=6.864 pd=35.98 as=2.904 ps=17.93 w=17.6 l=0.27
X9 VDD1.t0 VP.t3 VTAIL.t1 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=2.904 pd=17.93 as=6.864 ps=35.98 w=17.6 l=0.27
X10 VDD2.t0 VN.t2 VTAIL.t5 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=2.904 pd=17.93 as=6.864 ps=35.98 w=17.6 l=0.27
X11 VDD2.t3 VN.t3 VTAIL.t4 w_n1330_n4492# sky130_fd_pr__pfet_01v8 ad=2.904 pd=17.93 as=6.864 ps=35.98 w=17.6 l=0.27
R0 B.n125 B.t0 1791.69
R1 B.n281 B.t6 1791.69
R2 B.n46 B.t3 1791.69
R3 B.n38 B.t9 1791.69
R4 B.n372 B.n371 585
R5 B.n370 B.n91 585
R6 B.n369 B.n368 585
R7 B.n367 B.n92 585
R8 B.n366 B.n365 585
R9 B.n364 B.n93 585
R10 B.n363 B.n362 585
R11 B.n361 B.n94 585
R12 B.n360 B.n359 585
R13 B.n358 B.n95 585
R14 B.n357 B.n356 585
R15 B.n355 B.n96 585
R16 B.n354 B.n353 585
R17 B.n352 B.n97 585
R18 B.n351 B.n350 585
R19 B.n349 B.n98 585
R20 B.n348 B.n347 585
R21 B.n346 B.n99 585
R22 B.n345 B.n344 585
R23 B.n343 B.n100 585
R24 B.n342 B.n341 585
R25 B.n340 B.n101 585
R26 B.n339 B.n338 585
R27 B.n337 B.n102 585
R28 B.n336 B.n335 585
R29 B.n334 B.n103 585
R30 B.n333 B.n332 585
R31 B.n331 B.n104 585
R32 B.n330 B.n329 585
R33 B.n328 B.n105 585
R34 B.n327 B.n326 585
R35 B.n325 B.n106 585
R36 B.n324 B.n323 585
R37 B.n322 B.n107 585
R38 B.n321 B.n320 585
R39 B.n319 B.n108 585
R40 B.n318 B.n317 585
R41 B.n316 B.n109 585
R42 B.n315 B.n314 585
R43 B.n313 B.n110 585
R44 B.n312 B.n311 585
R45 B.n310 B.n111 585
R46 B.n309 B.n308 585
R47 B.n307 B.n112 585
R48 B.n306 B.n305 585
R49 B.n304 B.n113 585
R50 B.n303 B.n302 585
R51 B.n301 B.n114 585
R52 B.n300 B.n299 585
R53 B.n298 B.n115 585
R54 B.n297 B.n296 585
R55 B.n295 B.n116 585
R56 B.n294 B.n293 585
R57 B.n292 B.n117 585
R58 B.n291 B.n290 585
R59 B.n289 B.n118 585
R60 B.n288 B.n287 585
R61 B.n286 B.n119 585
R62 B.n285 B.n284 585
R63 B.n280 B.n120 585
R64 B.n279 B.n278 585
R65 B.n277 B.n121 585
R66 B.n276 B.n275 585
R67 B.n274 B.n122 585
R68 B.n273 B.n272 585
R69 B.n271 B.n123 585
R70 B.n270 B.n269 585
R71 B.n268 B.n124 585
R72 B.n266 B.n265 585
R73 B.n264 B.n127 585
R74 B.n263 B.n262 585
R75 B.n261 B.n128 585
R76 B.n260 B.n259 585
R77 B.n258 B.n129 585
R78 B.n257 B.n256 585
R79 B.n255 B.n130 585
R80 B.n254 B.n253 585
R81 B.n252 B.n131 585
R82 B.n251 B.n250 585
R83 B.n249 B.n132 585
R84 B.n248 B.n247 585
R85 B.n246 B.n133 585
R86 B.n245 B.n244 585
R87 B.n243 B.n134 585
R88 B.n242 B.n241 585
R89 B.n240 B.n135 585
R90 B.n239 B.n238 585
R91 B.n237 B.n136 585
R92 B.n236 B.n235 585
R93 B.n234 B.n137 585
R94 B.n233 B.n232 585
R95 B.n231 B.n138 585
R96 B.n230 B.n229 585
R97 B.n228 B.n139 585
R98 B.n227 B.n226 585
R99 B.n225 B.n140 585
R100 B.n224 B.n223 585
R101 B.n222 B.n141 585
R102 B.n221 B.n220 585
R103 B.n219 B.n142 585
R104 B.n218 B.n217 585
R105 B.n216 B.n143 585
R106 B.n215 B.n214 585
R107 B.n213 B.n144 585
R108 B.n212 B.n211 585
R109 B.n210 B.n145 585
R110 B.n209 B.n208 585
R111 B.n207 B.n146 585
R112 B.n206 B.n205 585
R113 B.n204 B.n147 585
R114 B.n203 B.n202 585
R115 B.n201 B.n148 585
R116 B.n200 B.n199 585
R117 B.n198 B.n149 585
R118 B.n197 B.n196 585
R119 B.n195 B.n150 585
R120 B.n194 B.n193 585
R121 B.n192 B.n151 585
R122 B.n191 B.n190 585
R123 B.n189 B.n152 585
R124 B.n188 B.n187 585
R125 B.n186 B.n153 585
R126 B.n185 B.n184 585
R127 B.n183 B.n154 585
R128 B.n182 B.n181 585
R129 B.n180 B.n155 585
R130 B.n373 B.n90 585
R131 B.n375 B.n374 585
R132 B.n376 B.n89 585
R133 B.n378 B.n377 585
R134 B.n379 B.n88 585
R135 B.n381 B.n380 585
R136 B.n382 B.n87 585
R137 B.n384 B.n383 585
R138 B.n385 B.n86 585
R139 B.n387 B.n386 585
R140 B.n388 B.n85 585
R141 B.n390 B.n389 585
R142 B.n391 B.n84 585
R143 B.n393 B.n392 585
R144 B.n394 B.n83 585
R145 B.n396 B.n395 585
R146 B.n397 B.n82 585
R147 B.n399 B.n398 585
R148 B.n400 B.n81 585
R149 B.n402 B.n401 585
R150 B.n403 B.n80 585
R151 B.n405 B.n404 585
R152 B.n406 B.n79 585
R153 B.n408 B.n407 585
R154 B.n409 B.n78 585
R155 B.n411 B.n410 585
R156 B.n412 B.n77 585
R157 B.n414 B.n413 585
R158 B.n604 B.n603 585
R159 B.n602 B.n9 585
R160 B.n601 B.n600 585
R161 B.n599 B.n10 585
R162 B.n598 B.n597 585
R163 B.n596 B.n11 585
R164 B.n595 B.n594 585
R165 B.n593 B.n12 585
R166 B.n592 B.n591 585
R167 B.n590 B.n13 585
R168 B.n589 B.n588 585
R169 B.n587 B.n14 585
R170 B.n586 B.n585 585
R171 B.n584 B.n15 585
R172 B.n583 B.n582 585
R173 B.n581 B.n16 585
R174 B.n580 B.n579 585
R175 B.n578 B.n17 585
R176 B.n577 B.n576 585
R177 B.n575 B.n18 585
R178 B.n574 B.n573 585
R179 B.n572 B.n19 585
R180 B.n571 B.n570 585
R181 B.n569 B.n20 585
R182 B.n568 B.n567 585
R183 B.n566 B.n21 585
R184 B.n565 B.n564 585
R185 B.n563 B.n22 585
R186 B.n562 B.n561 585
R187 B.n560 B.n23 585
R188 B.n559 B.n558 585
R189 B.n557 B.n24 585
R190 B.n556 B.n555 585
R191 B.n554 B.n25 585
R192 B.n553 B.n552 585
R193 B.n551 B.n26 585
R194 B.n550 B.n549 585
R195 B.n548 B.n27 585
R196 B.n547 B.n546 585
R197 B.n545 B.n28 585
R198 B.n544 B.n543 585
R199 B.n542 B.n29 585
R200 B.n541 B.n540 585
R201 B.n539 B.n30 585
R202 B.n538 B.n537 585
R203 B.n536 B.n31 585
R204 B.n535 B.n534 585
R205 B.n533 B.n32 585
R206 B.n532 B.n531 585
R207 B.n530 B.n33 585
R208 B.n529 B.n528 585
R209 B.n527 B.n34 585
R210 B.n526 B.n525 585
R211 B.n524 B.n35 585
R212 B.n523 B.n522 585
R213 B.n521 B.n36 585
R214 B.n520 B.n519 585
R215 B.n518 B.n37 585
R216 B.n516 B.n515 585
R217 B.n514 B.n40 585
R218 B.n513 B.n512 585
R219 B.n511 B.n41 585
R220 B.n510 B.n509 585
R221 B.n508 B.n42 585
R222 B.n507 B.n506 585
R223 B.n505 B.n43 585
R224 B.n504 B.n503 585
R225 B.n502 B.n44 585
R226 B.n501 B.n500 585
R227 B.n499 B.n45 585
R228 B.n498 B.n497 585
R229 B.n496 B.n49 585
R230 B.n495 B.n494 585
R231 B.n493 B.n50 585
R232 B.n492 B.n491 585
R233 B.n490 B.n51 585
R234 B.n489 B.n488 585
R235 B.n487 B.n52 585
R236 B.n486 B.n485 585
R237 B.n484 B.n53 585
R238 B.n483 B.n482 585
R239 B.n481 B.n54 585
R240 B.n480 B.n479 585
R241 B.n478 B.n55 585
R242 B.n477 B.n476 585
R243 B.n475 B.n56 585
R244 B.n474 B.n473 585
R245 B.n472 B.n57 585
R246 B.n471 B.n470 585
R247 B.n469 B.n58 585
R248 B.n468 B.n467 585
R249 B.n466 B.n59 585
R250 B.n465 B.n464 585
R251 B.n463 B.n60 585
R252 B.n462 B.n461 585
R253 B.n460 B.n61 585
R254 B.n459 B.n458 585
R255 B.n457 B.n62 585
R256 B.n456 B.n455 585
R257 B.n454 B.n63 585
R258 B.n453 B.n452 585
R259 B.n451 B.n64 585
R260 B.n450 B.n449 585
R261 B.n448 B.n65 585
R262 B.n447 B.n446 585
R263 B.n445 B.n66 585
R264 B.n444 B.n443 585
R265 B.n442 B.n67 585
R266 B.n441 B.n440 585
R267 B.n439 B.n68 585
R268 B.n438 B.n437 585
R269 B.n436 B.n69 585
R270 B.n435 B.n434 585
R271 B.n433 B.n70 585
R272 B.n432 B.n431 585
R273 B.n430 B.n71 585
R274 B.n429 B.n428 585
R275 B.n427 B.n72 585
R276 B.n426 B.n425 585
R277 B.n424 B.n73 585
R278 B.n423 B.n422 585
R279 B.n421 B.n74 585
R280 B.n420 B.n419 585
R281 B.n418 B.n75 585
R282 B.n417 B.n416 585
R283 B.n415 B.n76 585
R284 B.n605 B.n8 585
R285 B.n607 B.n606 585
R286 B.n608 B.n7 585
R287 B.n610 B.n609 585
R288 B.n611 B.n6 585
R289 B.n613 B.n612 585
R290 B.n614 B.n5 585
R291 B.n616 B.n615 585
R292 B.n617 B.n4 585
R293 B.n619 B.n618 585
R294 B.n620 B.n3 585
R295 B.n622 B.n621 585
R296 B.n623 B.n0 585
R297 B.n2 B.n1 585
R298 B.n162 B.n161 585
R299 B.n164 B.n163 585
R300 B.n165 B.n160 585
R301 B.n167 B.n166 585
R302 B.n168 B.n159 585
R303 B.n170 B.n169 585
R304 B.n171 B.n158 585
R305 B.n173 B.n172 585
R306 B.n174 B.n157 585
R307 B.n176 B.n175 585
R308 B.n177 B.n156 585
R309 B.n179 B.n178 585
R310 B.n281 B.t7 488.252
R311 B.n46 B.t5 488.252
R312 B.n125 B.t1 488.252
R313 B.n38 B.t11 488.252
R314 B.n282 B.t8 476.616
R315 B.n47 B.t4 476.616
R316 B.n126 B.t2 476.616
R317 B.n39 B.t10 476.616
R318 B.n180 B.n179 473.281
R319 B.n371 B.n90 473.281
R320 B.n413 B.n76 473.281
R321 B.n605 B.n604 473.281
R322 B.n625 B.n624 256.663
R323 B.n624 B.n623 235.042
R324 B.n624 B.n2 235.042
R325 B.n181 B.n180 163.367
R326 B.n181 B.n154 163.367
R327 B.n185 B.n154 163.367
R328 B.n186 B.n185 163.367
R329 B.n187 B.n186 163.367
R330 B.n187 B.n152 163.367
R331 B.n191 B.n152 163.367
R332 B.n192 B.n191 163.367
R333 B.n193 B.n192 163.367
R334 B.n193 B.n150 163.367
R335 B.n197 B.n150 163.367
R336 B.n198 B.n197 163.367
R337 B.n199 B.n198 163.367
R338 B.n199 B.n148 163.367
R339 B.n203 B.n148 163.367
R340 B.n204 B.n203 163.367
R341 B.n205 B.n204 163.367
R342 B.n205 B.n146 163.367
R343 B.n209 B.n146 163.367
R344 B.n210 B.n209 163.367
R345 B.n211 B.n210 163.367
R346 B.n211 B.n144 163.367
R347 B.n215 B.n144 163.367
R348 B.n216 B.n215 163.367
R349 B.n217 B.n216 163.367
R350 B.n217 B.n142 163.367
R351 B.n221 B.n142 163.367
R352 B.n222 B.n221 163.367
R353 B.n223 B.n222 163.367
R354 B.n223 B.n140 163.367
R355 B.n227 B.n140 163.367
R356 B.n228 B.n227 163.367
R357 B.n229 B.n228 163.367
R358 B.n229 B.n138 163.367
R359 B.n233 B.n138 163.367
R360 B.n234 B.n233 163.367
R361 B.n235 B.n234 163.367
R362 B.n235 B.n136 163.367
R363 B.n239 B.n136 163.367
R364 B.n240 B.n239 163.367
R365 B.n241 B.n240 163.367
R366 B.n241 B.n134 163.367
R367 B.n245 B.n134 163.367
R368 B.n246 B.n245 163.367
R369 B.n247 B.n246 163.367
R370 B.n247 B.n132 163.367
R371 B.n251 B.n132 163.367
R372 B.n252 B.n251 163.367
R373 B.n253 B.n252 163.367
R374 B.n253 B.n130 163.367
R375 B.n257 B.n130 163.367
R376 B.n258 B.n257 163.367
R377 B.n259 B.n258 163.367
R378 B.n259 B.n128 163.367
R379 B.n263 B.n128 163.367
R380 B.n264 B.n263 163.367
R381 B.n265 B.n264 163.367
R382 B.n265 B.n124 163.367
R383 B.n270 B.n124 163.367
R384 B.n271 B.n270 163.367
R385 B.n272 B.n271 163.367
R386 B.n272 B.n122 163.367
R387 B.n276 B.n122 163.367
R388 B.n277 B.n276 163.367
R389 B.n278 B.n277 163.367
R390 B.n278 B.n120 163.367
R391 B.n285 B.n120 163.367
R392 B.n286 B.n285 163.367
R393 B.n287 B.n286 163.367
R394 B.n287 B.n118 163.367
R395 B.n291 B.n118 163.367
R396 B.n292 B.n291 163.367
R397 B.n293 B.n292 163.367
R398 B.n293 B.n116 163.367
R399 B.n297 B.n116 163.367
R400 B.n298 B.n297 163.367
R401 B.n299 B.n298 163.367
R402 B.n299 B.n114 163.367
R403 B.n303 B.n114 163.367
R404 B.n304 B.n303 163.367
R405 B.n305 B.n304 163.367
R406 B.n305 B.n112 163.367
R407 B.n309 B.n112 163.367
R408 B.n310 B.n309 163.367
R409 B.n311 B.n310 163.367
R410 B.n311 B.n110 163.367
R411 B.n315 B.n110 163.367
R412 B.n316 B.n315 163.367
R413 B.n317 B.n316 163.367
R414 B.n317 B.n108 163.367
R415 B.n321 B.n108 163.367
R416 B.n322 B.n321 163.367
R417 B.n323 B.n322 163.367
R418 B.n323 B.n106 163.367
R419 B.n327 B.n106 163.367
R420 B.n328 B.n327 163.367
R421 B.n329 B.n328 163.367
R422 B.n329 B.n104 163.367
R423 B.n333 B.n104 163.367
R424 B.n334 B.n333 163.367
R425 B.n335 B.n334 163.367
R426 B.n335 B.n102 163.367
R427 B.n339 B.n102 163.367
R428 B.n340 B.n339 163.367
R429 B.n341 B.n340 163.367
R430 B.n341 B.n100 163.367
R431 B.n345 B.n100 163.367
R432 B.n346 B.n345 163.367
R433 B.n347 B.n346 163.367
R434 B.n347 B.n98 163.367
R435 B.n351 B.n98 163.367
R436 B.n352 B.n351 163.367
R437 B.n353 B.n352 163.367
R438 B.n353 B.n96 163.367
R439 B.n357 B.n96 163.367
R440 B.n358 B.n357 163.367
R441 B.n359 B.n358 163.367
R442 B.n359 B.n94 163.367
R443 B.n363 B.n94 163.367
R444 B.n364 B.n363 163.367
R445 B.n365 B.n364 163.367
R446 B.n365 B.n92 163.367
R447 B.n369 B.n92 163.367
R448 B.n370 B.n369 163.367
R449 B.n371 B.n370 163.367
R450 B.n413 B.n412 163.367
R451 B.n412 B.n411 163.367
R452 B.n411 B.n78 163.367
R453 B.n407 B.n78 163.367
R454 B.n407 B.n406 163.367
R455 B.n406 B.n405 163.367
R456 B.n405 B.n80 163.367
R457 B.n401 B.n80 163.367
R458 B.n401 B.n400 163.367
R459 B.n400 B.n399 163.367
R460 B.n399 B.n82 163.367
R461 B.n395 B.n82 163.367
R462 B.n395 B.n394 163.367
R463 B.n394 B.n393 163.367
R464 B.n393 B.n84 163.367
R465 B.n389 B.n84 163.367
R466 B.n389 B.n388 163.367
R467 B.n388 B.n387 163.367
R468 B.n387 B.n86 163.367
R469 B.n383 B.n86 163.367
R470 B.n383 B.n382 163.367
R471 B.n382 B.n381 163.367
R472 B.n381 B.n88 163.367
R473 B.n377 B.n88 163.367
R474 B.n377 B.n376 163.367
R475 B.n376 B.n375 163.367
R476 B.n375 B.n90 163.367
R477 B.n604 B.n9 163.367
R478 B.n600 B.n9 163.367
R479 B.n600 B.n599 163.367
R480 B.n599 B.n598 163.367
R481 B.n598 B.n11 163.367
R482 B.n594 B.n11 163.367
R483 B.n594 B.n593 163.367
R484 B.n593 B.n592 163.367
R485 B.n592 B.n13 163.367
R486 B.n588 B.n13 163.367
R487 B.n588 B.n587 163.367
R488 B.n587 B.n586 163.367
R489 B.n586 B.n15 163.367
R490 B.n582 B.n15 163.367
R491 B.n582 B.n581 163.367
R492 B.n581 B.n580 163.367
R493 B.n580 B.n17 163.367
R494 B.n576 B.n17 163.367
R495 B.n576 B.n575 163.367
R496 B.n575 B.n574 163.367
R497 B.n574 B.n19 163.367
R498 B.n570 B.n19 163.367
R499 B.n570 B.n569 163.367
R500 B.n569 B.n568 163.367
R501 B.n568 B.n21 163.367
R502 B.n564 B.n21 163.367
R503 B.n564 B.n563 163.367
R504 B.n563 B.n562 163.367
R505 B.n562 B.n23 163.367
R506 B.n558 B.n23 163.367
R507 B.n558 B.n557 163.367
R508 B.n557 B.n556 163.367
R509 B.n556 B.n25 163.367
R510 B.n552 B.n25 163.367
R511 B.n552 B.n551 163.367
R512 B.n551 B.n550 163.367
R513 B.n550 B.n27 163.367
R514 B.n546 B.n27 163.367
R515 B.n546 B.n545 163.367
R516 B.n545 B.n544 163.367
R517 B.n544 B.n29 163.367
R518 B.n540 B.n29 163.367
R519 B.n540 B.n539 163.367
R520 B.n539 B.n538 163.367
R521 B.n538 B.n31 163.367
R522 B.n534 B.n31 163.367
R523 B.n534 B.n533 163.367
R524 B.n533 B.n532 163.367
R525 B.n532 B.n33 163.367
R526 B.n528 B.n33 163.367
R527 B.n528 B.n527 163.367
R528 B.n527 B.n526 163.367
R529 B.n526 B.n35 163.367
R530 B.n522 B.n35 163.367
R531 B.n522 B.n521 163.367
R532 B.n521 B.n520 163.367
R533 B.n520 B.n37 163.367
R534 B.n515 B.n37 163.367
R535 B.n515 B.n514 163.367
R536 B.n514 B.n513 163.367
R537 B.n513 B.n41 163.367
R538 B.n509 B.n41 163.367
R539 B.n509 B.n508 163.367
R540 B.n508 B.n507 163.367
R541 B.n507 B.n43 163.367
R542 B.n503 B.n43 163.367
R543 B.n503 B.n502 163.367
R544 B.n502 B.n501 163.367
R545 B.n501 B.n45 163.367
R546 B.n497 B.n45 163.367
R547 B.n497 B.n496 163.367
R548 B.n496 B.n495 163.367
R549 B.n495 B.n50 163.367
R550 B.n491 B.n50 163.367
R551 B.n491 B.n490 163.367
R552 B.n490 B.n489 163.367
R553 B.n489 B.n52 163.367
R554 B.n485 B.n52 163.367
R555 B.n485 B.n484 163.367
R556 B.n484 B.n483 163.367
R557 B.n483 B.n54 163.367
R558 B.n479 B.n54 163.367
R559 B.n479 B.n478 163.367
R560 B.n478 B.n477 163.367
R561 B.n477 B.n56 163.367
R562 B.n473 B.n56 163.367
R563 B.n473 B.n472 163.367
R564 B.n472 B.n471 163.367
R565 B.n471 B.n58 163.367
R566 B.n467 B.n58 163.367
R567 B.n467 B.n466 163.367
R568 B.n466 B.n465 163.367
R569 B.n465 B.n60 163.367
R570 B.n461 B.n60 163.367
R571 B.n461 B.n460 163.367
R572 B.n460 B.n459 163.367
R573 B.n459 B.n62 163.367
R574 B.n455 B.n62 163.367
R575 B.n455 B.n454 163.367
R576 B.n454 B.n453 163.367
R577 B.n453 B.n64 163.367
R578 B.n449 B.n64 163.367
R579 B.n449 B.n448 163.367
R580 B.n448 B.n447 163.367
R581 B.n447 B.n66 163.367
R582 B.n443 B.n66 163.367
R583 B.n443 B.n442 163.367
R584 B.n442 B.n441 163.367
R585 B.n441 B.n68 163.367
R586 B.n437 B.n68 163.367
R587 B.n437 B.n436 163.367
R588 B.n436 B.n435 163.367
R589 B.n435 B.n70 163.367
R590 B.n431 B.n70 163.367
R591 B.n431 B.n430 163.367
R592 B.n430 B.n429 163.367
R593 B.n429 B.n72 163.367
R594 B.n425 B.n72 163.367
R595 B.n425 B.n424 163.367
R596 B.n424 B.n423 163.367
R597 B.n423 B.n74 163.367
R598 B.n419 B.n74 163.367
R599 B.n419 B.n418 163.367
R600 B.n418 B.n417 163.367
R601 B.n417 B.n76 163.367
R602 B.n606 B.n605 163.367
R603 B.n606 B.n7 163.367
R604 B.n610 B.n7 163.367
R605 B.n611 B.n610 163.367
R606 B.n612 B.n611 163.367
R607 B.n612 B.n5 163.367
R608 B.n616 B.n5 163.367
R609 B.n617 B.n616 163.367
R610 B.n618 B.n617 163.367
R611 B.n618 B.n3 163.367
R612 B.n622 B.n3 163.367
R613 B.n623 B.n622 163.367
R614 B.n162 B.n2 163.367
R615 B.n163 B.n162 163.367
R616 B.n163 B.n160 163.367
R617 B.n167 B.n160 163.367
R618 B.n168 B.n167 163.367
R619 B.n169 B.n168 163.367
R620 B.n169 B.n158 163.367
R621 B.n173 B.n158 163.367
R622 B.n174 B.n173 163.367
R623 B.n175 B.n174 163.367
R624 B.n175 B.n156 163.367
R625 B.n179 B.n156 163.367
R626 B.n267 B.n126 59.5399
R627 B.n283 B.n282 59.5399
R628 B.n48 B.n47 59.5399
R629 B.n517 B.n39 59.5399
R630 B.n603 B.n8 30.7517
R631 B.n415 B.n414 30.7517
R632 B.n373 B.n372 30.7517
R633 B.n178 B.n155 30.7517
R634 B B.n625 18.0485
R635 B.n126 B.n125 11.6369
R636 B.n282 B.n281 11.6369
R637 B.n47 B.n46 11.6369
R638 B.n39 B.n38 11.6369
R639 B.n607 B.n8 10.6151
R640 B.n608 B.n607 10.6151
R641 B.n609 B.n608 10.6151
R642 B.n609 B.n6 10.6151
R643 B.n613 B.n6 10.6151
R644 B.n614 B.n613 10.6151
R645 B.n615 B.n614 10.6151
R646 B.n615 B.n4 10.6151
R647 B.n619 B.n4 10.6151
R648 B.n620 B.n619 10.6151
R649 B.n621 B.n620 10.6151
R650 B.n621 B.n0 10.6151
R651 B.n603 B.n602 10.6151
R652 B.n602 B.n601 10.6151
R653 B.n601 B.n10 10.6151
R654 B.n597 B.n10 10.6151
R655 B.n597 B.n596 10.6151
R656 B.n596 B.n595 10.6151
R657 B.n595 B.n12 10.6151
R658 B.n591 B.n12 10.6151
R659 B.n591 B.n590 10.6151
R660 B.n590 B.n589 10.6151
R661 B.n589 B.n14 10.6151
R662 B.n585 B.n14 10.6151
R663 B.n585 B.n584 10.6151
R664 B.n584 B.n583 10.6151
R665 B.n583 B.n16 10.6151
R666 B.n579 B.n16 10.6151
R667 B.n579 B.n578 10.6151
R668 B.n578 B.n577 10.6151
R669 B.n577 B.n18 10.6151
R670 B.n573 B.n18 10.6151
R671 B.n573 B.n572 10.6151
R672 B.n572 B.n571 10.6151
R673 B.n571 B.n20 10.6151
R674 B.n567 B.n20 10.6151
R675 B.n567 B.n566 10.6151
R676 B.n566 B.n565 10.6151
R677 B.n565 B.n22 10.6151
R678 B.n561 B.n22 10.6151
R679 B.n561 B.n560 10.6151
R680 B.n560 B.n559 10.6151
R681 B.n559 B.n24 10.6151
R682 B.n555 B.n24 10.6151
R683 B.n555 B.n554 10.6151
R684 B.n554 B.n553 10.6151
R685 B.n553 B.n26 10.6151
R686 B.n549 B.n26 10.6151
R687 B.n549 B.n548 10.6151
R688 B.n548 B.n547 10.6151
R689 B.n547 B.n28 10.6151
R690 B.n543 B.n28 10.6151
R691 B.n543 B.n542 10.6151
R692 B.n542 B.n541 10.6151
R693 B.n541 B.n30 10.6151
R694 B.n537 B.n30 10.6151
R695 B.n537 B.n536 10.6151
R696 B.n536 B.n535 10.6151
R697 B.n535 B.n32 10.6151
R698 B.n531 B.n32 10.6151
R699 B.n531 B.n530 10.6151
R700 B.n530 B.n529 10.6151
R701 B.n529 B.n34 10.6151
R702 B.n525 B.n34 10.6151
R703 B.n525 B.n524 10.6151
R704 B.n524 B.n523 10.6151
R705 B.n523 B.n36 10.6151
R706 B.n519 B.n36 10.6151
R707 B.n519 B.n518 10.6151
R708 B.n516 B.n40 10.6151
R709 B.n512 B.n40 10.6151
R710 B.n512 B.n511 10.6151
R711 B.n511 B.n510 10.6151
R712 B.n510 B.n42 10.6151
R713 B.n506 B.n42 10.6151
R714 B.n506 B.n505 10.6151
R715 B.n505 B.n504 10.6151
R716 B.n504 B.n44 10.6151
R717 B.n500 B.n499 10.6151
R718 B.n499 B.n498 10.6151
R719 B.n498 B.n49 10.6151
R720 B.n494 B.n49 10.6151
R721 B.n494 B.n493 10.6151
R722 B.n493 B.n492 10.6151
R723 B.n492 B.n51 10.6151
R724 B.n488 B.n51 10.6151
R725 B.n488 B.n487 10.6151
R726 B.n487 B.n486 10.6151
R727 B.n486 B.n53 10.6151
R728 B.n482 B.n53 10.6151
R729 B.n482 B.n481 10.6151
R730 B.n481 B.n480 10.6151
R731 B.n480 B.n55 10.6151
R732 B.n476 B.n55 10.6151
R733 B.n476 B.n475 10.6151
R734 B.n475 B.n474 10.6151
R735 B.n474 B.n57 10.6151
R736 B.n470 B.n57 10.6151
R737 B.n470 B.n469 10.6151
R738 B.n469 B.n468 10.6151
R739 B.n468 B.n59 10.6151
R740 B.n464 B.n59 10.6151
R741 B.n464 B.n463 10.6151
R742 B.n463 B.n462 10.6151
R743 B.n462 B.n61 10.6151
R744 B.n458 B.n61 10.6151
R745 B.n458 B.n457 10.6151
R746 B.n457 B.n456 10.6151
R747 B.n456 B.n63 10.6151
R748 B.n452 B.n63 10.6151
R749 B.n452 B.n451 10.6151
R750 B.n451 B.n450 10.6151
R751 B.n450 B.n65 10.6151
R752 B.n446 B.n65 10.6151
R753 B.n446 B.n445 10.6151
R754 B.n445 B.n444 10.6151
R755 B.n444 B.n67 10.6151
R756 B.n440 B.n67 10.6151
R757 B.n440 B.n439 10.6151
R758 B.n439 B.n438 10.6151
R759 B.n438 B.n69 10.6151
R760 B.n434 B.n69 10.6151
R761 B.n434 B.n433 10.6151
R762 B.n433 B.n432 10.6151
R763 B.n432 B.n71 10.6151
R764 B.n428 B.n71 10.6151
R765 B.n428 B.n427 10.6151
R766 B.n427 B.n426 10.6151
R767 B.n426 B.n73 10.6151
R768 B.n422 B.n73 10.6151
R769 B.n422 B.n421 10.6151
R770 B.n421 B.n420 10.6151
R771 B.n420 B.n75 10.6151
R772 B.n416 B.n75 10.6151
R773 B.n416 B.n415 10.6151
R774 B.n414 B.n77 10.6151
R775 B.n410 B.n77 10.6151
R776 B.n410 B.n409 10.6151
R777 B.n409 B.n408 10.6151
R778 B.n408 B.n79 10.6151
R779 B.n404 B.n79 10.6151
R780 B.n404 B.n403 10.6151
R781 B.n403 B.n402 10.6151
R782 B.n402 B.n81 10.6151
R783 B.n398 B.n81 10.6151
R784 B.n398 B.n397 10.6151
R785 B.n397 B.n396 10.6151
R786 B.n396 B.n83 10.6151
R787 B.n392 B.n83 10.6151
R788 B.n392 B.n391 10.6151
R789 B.n391 B.n390 10.6151
R790 B.n390 B.n85 10.6151
R791 B.n386 B.n85 10.6151
R792 B.n386 B.n385 10.6151
R793 B.n385 B.n384 10.6151
R794 B.n384 B.n87 10.6151
R795 B.n380 B.n87 10.6151
R796 B.n380 B.n379 10.6151
R797 B.n379 B.n378 10.6151
R798 B.n378 B.n89 10.6151
R799 B.n374 B.n89 10.6151
R800 B.n374 B.n373 10.6151
R801 B.n161 B.n1 10.6151
R802 B.n164 B.n161 10.6151
R803 B.n165 B.n164 10.6151
R804 B.n166 B.n165 10.6151
R805 B.n166 B.n159 10.6151
R806 B.n170 B.n159 10.6151
R807 B.n171 B.n170 10.6151
R808 B.n172 B.n171 10.6151
R809 B.n172 B.n157 10.6151
R810 B.n176 B.n157 10.6151
R811 B.n177 B.n176 10.6151
R812 B.n178 B.n177 10.6151
R813 B.n182 B.n155 10.6151
R814 B.n183 B.n182 10.6151
R815 B.n184 B.n183 10.6151
R816 B.n184 B.n153 10.6151
R817 B.n188 B.n153 10.6151
R818 B.n189 B.n188 10.6151
R819 B.n190 B.n189 10.6151
R820 B.n190 B.n151 10.6151
R821 B.n194 B.n151 10.6151
R822 B.n195 B.n194 10.6151
R823 B.n196 B.n195 10.6151
R824 B.n196 B.n149 10.6151
R825 B.n200 B.n149 10.6151
R826 B.n201 B.n200 10.6151
R827 B.n202 B.n201 10.6151
R828 B.n202 B.n147 10.6151
R829 B.n206 B.n147 10.6151
R830 B.n207 B.n206 10.6151
R831 B.n208 B.n207 10.6151
R832 B.n208 B.n145 10.6151
R833 B.n212 B.n145 10.6151
R834 B.n213 B.n212 10.6151
R835 B.n214 B.n213 10.6151
R836 B.n214 B.n143 10.6151
R837 B.n218 B.n143 10.6151
R838 B.n219 B.n218 10.6151
R839 B.n220 B.n219 10.6151
R840 B.n220 B.n141 10.6151
R841 B.n224 B.n141 10.6151
R842 B.n225 B.n224 10.6151
R843 B.n226 B.n225 10.6151
R844 B.n226 B.n139 10.6151
R845 B.n230 B.n139 10.6151
R846 B.n231 B.n230 10.6151
R847 B.n232 B.n231 10.6151
R848 B.n232 B.n137 10.6151
R849 B.n236 B.n137 10.6151
R850 B.n237 B.n236 10.6151
R851 B.n238 B.n237 10.6151
R852 B.n238 B.n135 10.6151
R853 B.n242 B.n135 10.6151
R854 B.n243 B.n242 10.6151
R855 B.n244 B.n243 10.6151
R856 B.n244 B.n133 10.6151
R857 B.n248 B.n133 10.6151
R858 B.n249 B.n248 10.6151
R859 B.n250 B.n249 10.6151
R860 B.n250 B.n131 10.6151
R861 B.n254 B.n131 10.6151
R862 B.n255 B.n254 10.6151
R863 B.n256 B.n255 10.6151
R864 B.n256 B.n129 10.6151
R865 B.n260 B.n129 10.6151
R866 B.n261 B.n260 10.6151
R867 B.n262 B.n261 10.6151
R868 B.n262 B.n127 10.6151
R869 B.n266 B.n127 10.6151
R870 B.n269 B.n268 10.6151
R871 B.n269 B.n123 10.6151
R872 B.n273 B.n123 10.6151
R873 B.n274 B.n273 10.6151
R874 B.n275 B.n274 10.6151
R875 B.n275 B.n121 10.6151
R876 B.n279 B.n121 10.6151
R877 B.n280 B.n279 10.6151
R878 B.n284 B.n280 10.6151
R879 B.n288 B.n119 10.6151
R880 B.n289 B.n288 10.6151
R881 B.n290 B.n289 10.6151
R882 B.n290 B.n117 10.6151
R883 B.n294 B.n117 10.6151
R884 B.n295 B.n294 10.6151
R885 B.n296 B.n295 10.6151
R886 B.n296 B.n115 10.6151
R887 B.n300 B.n115 10.6151
R888 B.n301 B.n300 10.6151
R889 B.n302 B.n301 10.6151
R890 B.n302 B.n113 10.6151
R891 B.n306 B.n113 10.6151
R892 B.n307 B.n306 10.6151
R893 B.n308 B.n307 10.6151
R894 B.n308 B.n111 10.6151
R895 B.n312 B.n111 10.6151
R896 B.n313 B.n312 10.6151
R897 B.n314 B.n313 10.6151
R898 B.n314 B.n109 10.6151
R899 B.n318 B.n109 10.6151
R900 B.n319 B.n318 10.6151
R901 B.n320 B.n319 10.6151
R902 B.n320 B.n107 10.6151
R903 B.n324 B.n107 10.6151
R904 B.n325 B.n324 10.6151
R905 B.n326 B.n325 10.6151
R906 B.n326 B.n105 10.6151
R907 B.n330 B.n105 10.6151
R908 B.n331 B.n330 10.6151
R909 B.n332 B.n331 10.6151
R910 B.n332 B.n103 10.6151
R911 B.n336 B.n103 10.6151
R912 B.n337 B.n336 10.6151
R913 B.n338 B.n337 10.6151
R914 B.n338 B.n101 10.6151
R915 B.n342 B.n101 10.6151
R916 B.n343 B.n342 10.6151
R917 B.n344 B.n343 10.6151
R918 B.n344 B.n99 10.6151
R919 B.n348 B.n99 10.6151
R920 B.n349 B.n348 10.6151
R921 B.n350 B.n349 10.6151
R922 B.n350 B.n97 10.6151
R923 B.n354 B.n97 10.6151
R924 B.n355 B.n354 10.6151
R925 B.n356 B.n355 10.6151
R926 B.n356 B.n95 10.6151
R927 B.n360 B.n95 10.6151
R928 B.n361 B.n360 10.6151
R929 B.n362 B.n361 10.6151
R930 B.n362 B.n93 10.6151
R931 B.n366 B.n93 10.6151
R932 B.n367 B.n366 10.6151
R933 B.n368 B.n367 10.6151
R934 B.n368 B.n91 10.6151
R935 B.n372 B.n91 10.6151
R936 B.n518 B.n517 8.74196
R937 B.n500 B.n48 8.74196
R938 B.n267 B.n266 8.74196
R939 B.n283 B.n119 8.74196
R940 B.n625 B.n0 8.11757
R941 B.n625 B.n1 8.11757
R942 B.n517 B.n516 1.87367
R943 B.n48 B.n44 1.87367
R944 B.n268 B.n267 1.87367
R945 B.n284 B.n283 1.87367
R946 VN.n0 VN.t2 1732.6
R947 VN.n0 VN.t0 1732.6
R948 VN.n1 VN.t1 1732.6
R949 VN.n1 VN.t3 1732.6
R950 VN VN.n1 205.097
R951 VN VN.n0 161.351
R952 VDD2.n2 VDD2.n0 111.029
R953 VDD2.n2 VDD2.n1 70.5736
R954 VDD2.n1 VDD2.t1 1.84737
R955 VDD2.n1 VDD2.t3 1.84737
R956 VDD2.n0 VDD2.t2 1.84737
R957 VDD2.n0 VDD2.t0 1.84737
R958 VDD2 VDD2.n2 0.0586897
R959 VTAIL.n778 VTAIL.n686 756.745
R960 VTAIL.n92 VTAIL.n0 756.745
R961 VTAIL.n190 VTAIL.n98 756.745
R962 VTAIL.n288 VTAIL.n196 756.745
R963 VTAIL.n680 VTAIL.n588 756.745
R964 VTAIL.n582 VTAIL.n490 756.745
R965 VTAIL.n484 VTAIL.n392 756.745
R966 VTAIL.n386 VTAIL.n294 756.745
R967 VTAIL.n719 VTAIL.n718 585
R968 VTAIL.n721 VTAIL.n720 585
R969 VTAIL.n714 VTAIL.n713 585
R970 VTAIL.n727 VTAIL.n726 585
R971 VTAIL.n729 VTAIL.n728 585
R972 VTAIL.n710 VTAIL.n709 585
R973 VTAIL.n735 VTAIL.n734 585
R974 VTAIL.n737 VTAIL.n736 585
R975 VTAIL.n706 VTAIL.n705 585
R976 VTAIL.n743 VTAIL.n742 585
R977 VTAIL.n745 VTAIL.n744 585
R978 VTAIL.n702 VTAIL.n701 585
R979 VTAIL.n751 VTAIL.n750 585
R980 VTAIL.n753 VTAIL.n752 585
R981 VTAIL.n698 VTAIL.n697 585
R982 VTAIL.n760 VTAIL.n759 585
R983 VTAIL.n761 VTAIL.n696 585
R984 VTAIL.n763 VTAIL.n762 585
R985 VTAIL.n694 VTAIL.n693 585
R986 VTAIL.n769 VTAIL.n768 585
R987 VTAIL.n771 VTAIL.n770 585
R988 VTAIL.n690 VTAIL.n689 585
R989 VTAIL.n777 VTAIL.n776 585
R990 VTAIL.n779 VTAIL.n778 585
R991 VTAIL.n33 VTAIL.n32 585
R992 VTAIL.n35 VTAIL.n34 585
R993 VTAIL.n28 VTAIL.n27 585
R994 VTAIL.n41 VTAIL.n40 585
R995 VTAIL.n43 VTAIL.n42 585
R996 VTAIL.n24 VTAIL.n23 585
R997 VTAIL.n49 VTAIL.n48 585
R998 VTAIL.n51 VTAIL.n50 585
R999 VTAIL.n20 VTAIL.n19 585
R1000 VTAIL.n57 VTAIL.n56 585
R1001 VTAIL.n59 VTAIL.n58 585
R1002 VTAIL.n16 VTAIL.n15 585
R1003 VTAIL.n65 VTAIL.n64 585
R1004 VTAIL.n67 VTAIL.n66 585
R1005 VTAIL.n12 VTAIL.n11 585
R1006 VTAIL.n74 VTAIL.n73 585
R1007 VTAIL.n75 VTAIL.n10 585
R1008 VTAIL.n77 VTAIL.n76 585
R1009 VTAIL.n8 VTAIL.n7 585
R1010 VTAIL.n83 VTAIL.n82 585
R1011 VTAIL.n85 VTAIL.n84 585
R1012 VTAIL.n4 VTAIL.n3 585
R1013 VTAIL.n91 VTAIL.n90 585
R1014 VTAIL.n93 VTAIL.n92 585
R1015 VTAIL.n131 VTAIL.n130 585
R1016 VTAIL.n133 VTAIL.n132 585
R1017 VTAIL.n126 VTAIL.n125 585
R1018 VTAIL.n139 VTAIL.n138 585
R1019 VTAIL.n141 VTAIL.n140 585
R1020 VTAIL.n122 VTAIL.n121 585
R1021 VTAIL.n147 VTAIL.n146 585
R1022 VTAIL.n149 VTAIL.n148 585
R1023 VTAIL.n118 VTAIL.n117 585
R1024 VTAIL.n155 VTAIL.n154 585
R1025 VTAIL.n157 VTAIL.n156 585
R1026 VTAIL.n114 VTAIL.n113 585
R1027 VTAIL.n163 VTAIL.n162 585
R1028 VTAIL.n165 VTAIL.n164 585
R1029 VTAIL.n110 VTAIL.n109 585
R1030 VTAIL.n172 VTAIL.n171 585
R1031 VTAIL.n173 VTAIL.n108 585
R1032 VTAIL.n175 VTAIL.n174 585
R1033 VTAIL.n106 VTAIL.n105 585
R1034 VTAIL.n181 VTAIL.n180 585
R1035 VTAIL.n183 VTAIL.n182 585
R1036 VTAIL.n102 VTAIL.n101 585
R1037 VTAIL.n189 VTAIL.n188 585
R1038 VTAIL.n191 VTAIL.n190 585
R1039 VTAIL.n229 VTAIL.n228 585
R1040 VTAIL.n231 VTAIL.n230 585
R1041 VTAIL.n224 VTAIL.n223 585
R1042 VTAIL.n237 VTAIL.n236 585
R1043 VTAIL.n239 VTAIL.n238 585
R1044 VTAIL.n220 VTAIL.n219 585
R1045 VTAIL.n245 VTAIL.n244 585
R1046 VTAIL.n247 VTAIL.n246 585
R1047 VTAIL.n216 VTAIL.n215 585
R1048 VTAIL.n253 VTAIL.n252 585
R1049 VTAIL.n255 VTAIL.n254 585
R1050 VTAIL.n212 VTAIL.n211 585
R1051 VTAIL.n261 VTAIL.n260 585
R1052 VTAIL.n263 VTAIL.n262 585
R1053 VTAIL.n208 VTAIL.n207 585
R1054 VTAIL.n270 VTAIL.n269 585
R1055 VTAIL.n271 VTAIL.n206 585
R1056 VTAIL.n273 VTAIL.n272 585
R1057 VTAIL.n204 VTAIL.n203 585
R1058 VTAIL.n279 VTAIL.n278 585
R1059 VTAIL.n281 VTAIL.n280 585
R1060 VTAIL.n200 VTAIL.n199 585
R1061 VTAIL.n287 VTAIL.n286 585
R1062 VTAIL.n289 VTAIL.n288 585
R1063 VTAIL.n681 VTAIL.n680 585
R1064 VTAIL.n679 VTAIL.n678 585
R1065 VTAIL.n592 VTAIL.n591 585
R1066 VTAIL.n673 VTAIL.n672 585
R1067 VTAIL.n671 VTAIL.n670 585
R1068 VTAIL.n596 VTAIL.n595 585
R1069 VTAIL.n600 VTAIL.n598 585
R1070 VTAIL.n665 VTAIL.n664 585
R1071 VTAIL.n663 VTAIL.n662 585
R1072 VTAIL.n602 VTAIL.n601 585
R1073 VTAIL.n657 VTAIL.n656 585
R1074 VTAIL.n655 VTAIL.n654 585
R1075 VTAIL.n606 VTAIL.n605 585
R1076 VTAIL.n649 VTAIL.n648 585
R1077 VTAIL.n647 VTAIL.n646 585
R1078 VTAIL.n610 VTAIL.n609 585
R1079 VTAIL.n641 VTAIL.n640 585
R1080 VTAIL.n639 VTAIL.n638 585
R1081 VTAIL.n614 VTAIL.n613 585
R1082 VTAIL.n633 VTAIL.n632 585
R1083 VTAIL.n631 VTAIL.n630 585
R1084 VTAIL.n618 VTAIL.n617 585
R1085 VTAIL.n625 VTAIL.n624 585
R1086 VTAIL.n623 VTAIL.n622 585
R1087 VTAIL.n583 VTAIL.n582 585
R1088 VTAIL.n581 VTAIL.n580 585
R1089 VTAIL.n494 VTAIL.n493 585
R1090 VTAIL.n575 VTAIL.n574 585
R1091 VTAIL.n573 VTAIL.n572 585
R1092 VTAIL.n498 VTAIL.n497 585
R1093 VTAIL.n502 VTAIL.n500 585
R1094 VTAIL.n567 VTAIL.n566 585
R1095 VTAIL.n565 VTAIL.n564 585
R1096 VTAIL.n504 VTAIL.n503 585
R1097 VTAIL.n559 VTAIL.n558 585
R1098 VTAIL.n557 VTAIL.n556 585
R1099 VTAIL.n508 VTAIL.n507 585
R1100 VTAIL.n551 VTAIL.n550 585
R1101 VTAIL.n549 VTAIL.n548 585
R1102 VTAIL.n512 VTAIL.n511 585
R1103 VTAIL.n543 VTAIL.n542 585
R1104 VTAIL.n541 VTAIL.n540 585
R1105 VTAIL.n516 VTAIL.n515 585
R1106 VTAIL.n535 VTAIL.n534 585
R1107 VTAIL.n533 VTAIL.n532 585
R1108 VTAIL.n520 VTAIL.n519 585
R1109 VTAIL.n527 VTAIL.n526 585
R1110 VTAIL.n525 VTAIL.n524 585
R1111 VTAIL.n485 VTAIL.n484 585
R1112 VTAIL.n483 VTAIL.n482 585
R1113 VTAIL.n396 VTAIL.n395 585
R1114 VTAIL.n477 VTAIL.n476 585
R1115 VTAIL.n475 VTAIL.n474 585
R1116 VTAIL.n400 VTAIL.n399 585
R1117 VTAIL.n404 VTAIL.n402 585
R1118 VTAIL.n469 VTAIL.n468 585
R1119 VTAIL.n467 VTAIL.n466 585
R1120 VTAIL.n406 VTAIL.n405 585
R1121 VTAIL.n461 VTAIL.n460 585
R1122 VTAIL.n459 VTAIL.n458 585
R1123 VTAIL.n410 VTAIL.n409 585
R1124 VTAIL.n453 VTAIL.n452 585
R1125 VTAIL.n451 VTAIL.n450 585
R1126 VTAIL.n414 VTAIL.n413 585
R1127 VTAIL.n445 VTAIL.n444 585
R1128 VTAIL.n443 VTAIL.n442 585
R1129 VTAIL.n418 VTAIL.n417 585
R1130 VTAIL.n437 VTAIL.n436 585
R1131 VTAIL.n435 VTAIL.n434 585
R1132 VTAIL.n422 VTAIL.n421 585
R1133 VTAIL.n429 VTAIL.n428 585
R1134 VTAIL.n427 VTAIL.n426 585
R1135 VTAIL.n387 VTAIL.n386 585
R1136 VTAIL.n385 VTAIL.n384 585
R1137 VTAIL.n298 VTAIL.n297 585
R1138 VTAIL.n379 VTAIL.n378 585
R1139 VTAIL.n377 VTAIL.n376 585
R1140 VTAIL.n302 VTAIL.n301 585
R1141 VTAIL.n306 VTAIL.n304 585
R1142 VTAIL.n371 VTAIL.n370 585
R1143 VTAIL.n369 VTAIL.n368 585
R1144 VTAIL.n308 VTAIL.n307 585
R1145 VTAIL.n363 VTAIL.n362 585
R1146 VTAIL.n361 VTAIL.n360 585
R1147 VTAIL.n312 VTAIL.n311 585
R1148 VTAIL.n355 VTAIL.n354 585
R1149 VTAIL.n353 VTAIL.n352 585
R1150 VTAIL.n316 VTAIL.n315 585
R1151 VTAIL.n347 VTAIL.n346 585
R1152 VTAIL.n345 VTAIL.n344 585
R1153 VTAIL.n320 VTAIL.n319 585
R1154 VTAIL.n339 VTAIL.n338 585
R1155 VTAIL.n337 VTAIL.n336 585
R1156 VTAIL.n324 VTAIL.n323 585
R1157 VTAIL.n331 VTAIL.n330 585
R1158 VTAIL.n329 VTAIL.n328 585
R1159 VTAIL.n717 VTAIL.t5 327.466
R1160 VTAIL.n31 VTAIL.t7 327.466
R1161 VTAIL.n129 VTAIL.t2 327.466
R1162 VTAIL.n227 VTAIL.t0 327.466
R1163 VTAIL.n621 VTAIL.t1 327.466
R1164 VTAIL.n523 VTAIL.t3 327.466
R1165 VTAIL.n425 VTAIL.t4 327.466
R1166 VTAIL.n327 VTAIL.t6 327.466
R1167 VTAIL.n720 VTAIL.n719 171.744
R1168 VTAIL.n720 VTAIL.n713 171.744
R1169 VTAIL.n727 VTAIL.n713 171.744
R1170 VTAIL.n728 VTAIL.n727 171.744
R1171 VTAIL.n728 VTAIL.n709 171.744
R1172 VTAIL.n735 VTAIL.n709 171.744
R1173 VTAIL.n736 VTAIL.n735 171.744
R1174 VTAIL.n736 VTAIL.n705 171.744
R1175 VTAIL.n743 VTAIL.n705 171.744
R1176 VTAIL.n744 VTAIL.n743 171.744
R1177 VTAIL.n744 VTAIL.n701 171.744
R1178 VTAIL.n751 VTAIL.n701 171.744
R1179 VTAIL.n752 VTAIL.n751 171.744
R1180 VTAIL.n752 VTAIL.n697 171.744
R1181 VTAIL.n760 VTAIL.n697 171.744
R1182 VTAIL.n761 VTAIL.n760 171.744
R1183 VTAIL.n762 VTAIL.n761 171.744
R1184 VTAIL.n762 VTAIL.n693 171.744
R1185 VTAIL.n769 VTAIL.n693 171.744
R1186 VTAIL.n770 VTAIL.n769 171.744
R1187 VTAIL.n770 VTAIL.n689 171.744
R1188 VTAIL.n777 VTAIL.n689 171.744
R1189 VTAIL.n778 VTAIL.n777 171.744
R1190 VTAIL.n34 VTAIL.n33 171.744
R1191 VTAIL.n34 VTAIL.n27 171.744
R1192 VTAIL.n41 VTAIL.n27 171.744
R1193 VTAIL.n42 VTAIL.n41 171.744
R1194 VTAIL.n42 VTAIL.n23 171.744
R1195 VTAIL.n49 VTAIL.n23 171.744
R1196 VTAIL.n50 VTAIL.n49 171.744
R1197 VTAIL.n50 VTAIL.n19 171.744
R1198 VTAIL.n57 VTAIL.n19 171.744
R1199 VTAIL.n58 VTAIL.n57 171.744
R1200 VTAIL.n58 VTAIL.n15 171.744
R1201 VTAIL.n65 VTAIL.n15 171.744
R1202 VTAIL.n66 VTAIL.n65 171.744
R1203 VTAIL.n66 VTAIL.n11 171.744
R1204 VTAIL.n74 VTAIL.n11 171.744
R1205 VTAIL.n75 VTAIL.n74 171.744
R1206 VTAIL.n76 VTAIL.n75 171.744
R1207 VTAIL.n76 VTAIL.n7 171.744
R1208 VTAIL.n83 VTAIL.n7 171.744
R1209 VTAIL.n84 VTAIL.n83 171.744
R1210 VTAIL.n84 VTAIL.n3 171.744
R1211 VTAIL.n91 VTAIL.n3 171.744
R1212 VTAIL.n92 VTAIL.n91 171.744
R1213 VTAIL.n132 VTAIL.n131 171.744
R1214 VTAIL.n132 VTAIL.n125 171.744
R1215 VTAIL.n139 VTAIL.n125 171.744
R1216 VTAIL.n140 VTAIL.n139 171.744
R1217 VTAIL.n140 VTAIL.n121 171.744
R1218 VTAIL.n147 VTAIL.n121 171.744
R1219 VTAIL.n148 VTAIL.n147 171.744
R1220 VTAIL.n148 VTAIL.n117 171.744
R1221 VTAIL.n155 VTAIL.n117 171.744
R1222 VTAIL.n156 VTAIL.n155 171.744
R1223 VTAIL.n156 VTAIL.n113 171.744
R1224 VTAIL.n163 VTAIL.n113 171.744
R1225 VTAIL.n164 VTAIL.n163 171.744
R1226 VTAIL.n164 VTAIL.n109 171.744
R1227 VTAIL.n172 VTAIL.n109 171.744
R1228 VTAIL.n173 VTAIL.n172 171.744
R1229 VTAIL.n174 VTAIL.n173 171.744
R1230 VTAIL.n174 VTAIL.n105 171.744
R1231 VTAIL.n181 VTAIL.n105 171.744
R1232 VTAIL.n182 VTAIL.n181 171.744
R1233 VTAIL.n182 VTAIL.n101 171.744
R1234 VTAIL.n189 VTAIL.n101 171.744
R1235 VTAIL.n190 VTAIL.n189 171.744
R1236 VTAIL.n230 VTAIL.n229 171.744
R1237 VTAIL.n230 VTAIL.n223 171.744
R1238 VTAIL.n237 VTAIL.n223 171.744
R1239 VTAIL.n238 VTAIL.n237 171.744
R1240 VTAIL.n238 VTAIL.n219 171.744
R1241 VTAIL.n245 VTAIL.n219 171.744
R1242 VTAIL.n246 VTAIL.n245 171.744
R1243 VTAIL.n246 VTAIL.n215 171.744
R1244 VTAIL.n253 VTAIL.n215 171.744
R1245 VTAIL.n254 VTAIL.n253 171.744
R1246 VTAIL.n254 VTAIL.n211 171.744
R1247 VTAIL.n261 VTAIL.n211 171.744
R1248 VTAIL.n262 VTAIL.n261 171.744
R1249 VTAIL.n262 VTAIL.n207 171.744
R1250 VTAIL.n270 VTAIL.n207 171.744
R1251 VTAIL.n271 VTAIL.n270 171.744
R1252 VTAIL.n272 VTAIL.n271 171.744
R1253 VTAIL.n272 VTAIL.n203 171.744
R1254 VTAIL.n279 VTAIL.n203 171.744
R1255 VTAIL.n280 VTAIL.n279 171.744
R1256 VTAIL.n280 VTAIL.n199 171.744
R1257 VTAIL.n287 VTAIL.n199 171.744
R1258 VTAIL.n288 VTAIL.n287 171.744
R1259 VTAIL.n680 VTAIL.n679 171.744
R1260 VTAIL.n679 VTAIL.n591 171.744
R1261 VTAIL.n672 VTAIL.n591 171.744
R1262 VTAIL.n672 VTAIL.n671 171.744
R1263 VTAIL.n671 VTAIL.n595 171.744
R1264 VTAIL.n600 VTAIL.n595 171.744
R1265 VTAIL.n664 VTAIL.n600 171.744
R1266 VTAIL.n664 VTAIL.n663 171.744
R1267 VTAIL.n663 VTAIL.n601 171.744
R1268 VTAIL.n656 VTAIL.n601 171.744
R1269 VTAIL.n656 VTAIL.n655 171.744
R1270 VTAIL.n655 VTAIL.n605 171.744
R1271 VTAIL.n648 VTAIL.n605 171.744
R1272 VTAIL.n648 VTAIL.n647 171.744
R1273 VTAIL.n647 VTAIL.n609 171.744
R1274 VTAIL.n640 VTAIL.n609 171.744
R1275 VTAIL.n640 VTAIL.n639 171.744
R1276 VTAIL.n639 VTAIL.n613 171.744
R1277 VTAIL.n632 VTAIL.n613 171.744
R1278 VTAIL.n632 VTAIL.n631 171.744
R1279 VTAIL.n631 VTAIL.n617 171.744
R1280 VTAIL.n624 VTAIL.n617 171.744
R1281 VTAIL.n624 VTAIL.n623 171.744
R1282 VTAIL.n582 VTAIL.n581 171.744
R1283 VTAIL.n581 VTAIL.n493 171.744
R1284 VTAIL.n574 VTAIL.n493 171.744
R1285 VTAIL.n574 VTAIL.n573 171.744
R1286 VTAIL.n573 VTAIL.n497 171.744
R1287 VTAIL.n502 VTAIL.n497 171.744
R1288 VTAIL.n566 VTAIL.n502 171.744
R1289 VTAIL.n566 VTAIL.n565 171.744
R1290 VTAIL.n565 VTAIL.n503 171.744
R1291 VTAIL.n558 VTAIL.n503 171.744
R1292 VTAIL.n558 VTAIL.n557 171.744
R1293 VTAIL.n557 VTAIL.n507 171.744
R1294 VTAIL.n550 VTAIL.n507 171.744
R1295 VTAIL.n550 VTAIL.n549 171.744
R1296 VTAIL.n549 VTAIL.n511 171.744
R1297 VTAIL.n542 VTAIL.n511 171.744
R1298 VTAIL.n542 VTAIL.n541 171.744
R1299 VTAIL.n541 VTAIL.n515 171.744
R1300 VTAIL.n534 VTAIL.n515 171.744
R1301 VTAIL.n534 VTAIL.n533 171.744
R1302 VTAIL.n533 VTAIL.n519 171.744
R1303 VTAIL.n526 VTAIL.n519 171.744
R1304 VTAIL.n526 VTAIL.n525 171.744
R1305 VTAIL.n484 VTAIL.n483 171.744
R1306 VTAIL.n483 VTAIL.n395 171.744
R1307 VTAIL.n476 VTAIL.n395 171.744
R1308 VTAIL.n476 VTAIL.n475 171.744
R1309 VTAIL.n475 VTAIL.n399 171.744
R1310 VTAIL.n404 VTAIL.n399 171.744
R1311 VTAIL.n468 VTAIL.n404 171.744
R1312 VTAIL.n468 VTAIL.n467 171.744
R1313 VTAIL.n467 VTAIL.n405 171.744
R1314 VTAIL.n460 VTAIL.n405 171.744
R1315 VTAIL.n460 VTAIL.n459 171.744
R1316 VTAIL.n459 VTAIL.n409 171.744
R1317 VTAIL.n452 VTAIL.n409 171.744
R1318 VTAIL.n452 VTAIL.n451 171.744
R1319 VTAIL.n451 VTAIL.n413 171.744
R1320 VTAIL.n444 VTAIL.n413 171.744
R1321 VTAIL.n444 VTAIL.n443 171.744
R1322 VTAIL.n443 VTAIL.n417 171.744
R1323 VTAIL.n436 VTAIL.n417 171.744
R1324 VTAIL.n436 VTAIL.n435 171.744
R1325 VTAIL.n435 VTAIL.n421 171.744
R1326 VTAIL.n428 VTAIL.n421 171.744
R1327 VTAIL.n428 VTAIL.n427 171.744
R1328 VTAIL.n386 VTAIL.n385 171.744
R1329 VTAIL.n385 VTAIL.n297 171.744
R1330 VTAIL.n378 VTAIL.n297 171.744
R1331 VTAIL.n378 VTAIL.n377 171.744
R1332 VTAIL.n377 VTAIL.n301 171.744
R1333 VTAIL.n306 VTAIL.n301 171.744
R1334 VTAIL.n370 VTAIL.n306 171.744
R1335 VTAIL.n370 VTAIL.n369 171.744
R1336 VTAIL.n369 VTAIL.n307 171.744
R1337 VTAIL.n362 VTAIL.n307 171.744
R1338 VTAIL.n362 VTAIL.n361 171.744
R1339 VTAIL.n361 VTAIL.n311 171.744
R1340 VTAIL.n354 VTAIL.n311 171.744
R1341 VTAIL.n354 VTAIL.n353 171.744
R1342 VTAIL.n353 VTAIL.n315 171.744
R1343 VTAIL.n346 VTAIL.n315 171.744
R1344 VTAIL.n346 VTAIL.n345 171.744
R1345 VTAIL.n345 VTAIL.n319 171.744
R1346 VTAIL.n338 VTAIL.n319 171.744
R1347 VTAIL.n338 VTAIL.n337 171.744
R1348 VTAIL.n337 VTAIL.n323 171.744
R1349 VTAIL.n330 VTAIL.n323 171.744
R1350 VTAIL.n330 VTAIL.n329 171.744
R1351 VTAIL.n719 VTAIL.t5 85.8723
R1352 VTAIL.n33 VTAIL.t7 85.8723
R1353 VTAIL.n131 VTAIL.t2 85.8723
R1354 VTAIL.n229 VTAIL.t0 85.8723
R1355 VTAIL.n623 VTAIL.t1 85.8723
R1356 VTAIL.n525 VTAIL.t3 85.8723
R1357 VTAIL.n427 VTAIL.t4 85.8723
R1358 VTAIL.n329 VTAIL.t6 85.8723
R1359 VTAIL.n783 VTAIL.n782 33.7369
R1360 VTAIL.n97 VTAIL.n96 33.7369
R1361 VTAIL.n195 VTAIL.n194 33.7369
R1362 VTAIL.n293 VTAIL.n292 33.7369
R1363 VTAIL.n685 VTAIL.n684 33.7369
R1364 VTAIL.n587 VTAIL.n586 33.7369
R1365 VTAIL.n489 VTAIL.n488 33.7369
R1366 VTAIL.n391 VTAIL.n390 33.7369
R1367 VTAIL.n783 VTAIL.n685 28.0738
R1368 VTAIL.n391 VTAIL.n293 28.0738
R1369 VTAIL.n718 VTAIL.n717 16.3895
R1370 VTAIL.n32 VTAIL.n31 16.3895
R1371 VTAIL.n130 VTAIL.n129 16.3895
R1372 VTAIL.n228 VTAIL.n227 16.3895
R1373 VTAIL.n622 VTAIL.n621 16.3895
R1374 VTAIL.n524 VTAIL.n523 16.3895
R1375 VTAIL.n426 VTAIL.n425 16.3895
R1376 VTAIL.n328 VTAIL.n327 16.3895
R1377 VTAIL.n763 VTAIL.n694 13.1884
R1378 VTAIL.n77 VTAIL.n8 13.1884
R1379 VTAIL.n175 VTAIL.n106 13.1884
R1380 VTAIL.n273 VTAIL.n204 13.1884
R1381 VTAIL.n598 VTAIL.n596 13.1884
R1382 VTAIL.n500 VTAIL.n498 13.1884
R1383 VTAIL.n402 VTAIL.n400 13.1884
R1384 VTAIL.n304 VTAIL.n302 13.1884
R1385 VTAIL.n721 VTAIL.n716 12.8005
R1386 VTAIL.n764 VTAIL.n696 12.8005
R1387 VTAIL.n768 VTAIL.n767 12.8005
R1388 VTAIL.n35 VTAIL.n30 12.8005
R1389 VTAIL.n78 VTAIL.n10 12.8005
R1390 VTAIL.n82 VTAIL.n81 12.8005
R1391 VTAIL.n133 VTAIL.n128 12.8005
R1392 VTAIL.n176 VTAIL.n108 12.8005
R1393 VTAIL.n180 VTAIL.n179 12.8005
R1394 VTAIL.n231 VTAIL.n226 12.8005
R1395 VTAIL.n274 VTAIL.n206 12.8005
R1396 VTAIL.n278 VTAIL.n277 12.8005
R1397 VTAIL.n670 VTAIL.n669 12.8005
R1398 VTAIL.n666 VTAIL.n665 12.8005
R1399 VTAIL.n625 VTAIL.n620 12.8005
R1400 VTAIL.n572 VTAIL.n571 12.8005
R1401 VTAIL.n568 VTAIL.n567 12.8005
R1402 VTAIL.n527 VTAIL.n522 12.8005
R1403 VTAIL.n474 VTAIL.n473 12.8005
R1404 VTAIL.n470 VTAIL.n469 12.8005
R1405 VTAIL.n429 VTAIL.n424 12.8005
R1406 VTAIL.n376 VTAIL.n375 12.8005
R1407 VTAIL.n372 VTAIL.n371 12.8005
R1408 VTAIL.n331 VTAIL.n326 12.8005
R1409 VTAIL.n722 VTAIL.n714 12.0247
R1410 VTAIL.n759 VTAIL.n758 12.0247
R1411 VTAIL.n771 VTAIL.n692 12.0247
R1412 VTAIL.n36 VTAIL.n28 12.0247
R1413 VTAIL.n73 VTAIL.n72 12.0247
R1414 VTAIL.n85 VTAIL.n6 12.0247
R1415 VTAIL.n134 VTAIL.n126 12.0247
R1416 VTAIL.n171 VTAIL.n170 12.0247
R1417 VTAIL.n183 VTAIL.n104 12.0247
R1418 VTAIL.n232 VTAIL.n224 12.0247
R1419 VTAIL.n269 VTAIL.n268 12.0247
R1420 VTAIL.n281 VTAIL.n202 12.0247
R1421 VTAIL.n673 VTAIL.n594 12.0247
R1422 VTAIL.n662 VTAIL.n599 12.0247
R1423 VTAIL.n626 VTAIL.n618 12.0247
R1424 VTAIL.n575 VTAIL.n496 12.0247
R1425 VTAIL.n564 VTAIL.n501 12.0247
R1426 VTAIL.n528 VTAIL.n520 12.0247
R1427 VTAIL.n477 VTAIL.n398 12.0247
R1428 VTAIL.n466 VTAIL.n403 12.0247
R1429 VTAIL.n430 VTAIL.n422 12.0247
R1430 VTAIL.n379 VTAIL.n300 12.0247
R1431 VTAIL.n368 VTAIL.n305 12.0247
R1432 VTAIL.n332 VTAIL.n324 12.0247
R1433 VTAIL.n726 VTAIL.n725 11.249
R1434 VTAIL.n757 VTAIL.n698 11.249
R1435 VTAIL.n772 VTAIL.n690 11.249
R1436 VTAIL.n40 VTAIL.n39 11.249
R1437 VTAIL.n71 VTAIL.n12 11.249
R1438 VTAIL.n86 VTAIL.n4 11.249
R1439 VTAIL.n138 VTAIL.n137 11.249
R1440 VTAIL.n169 VTAIL.n110 11.249
R1441 VTAIL.n184 VTAIL.n102 11.249
R1442 VTAIL.n236 VTAIL.n235 11.249
R1443 VTAIL.n267 VTAIL.n208 11.249
R1444 VTAIL.n282 VTAIL.n200 11.249
R1445 VTAIL.n674 VTAIL.n592 11.249
R1446 VTAIL.n661 VTAIL.n602 11.249
R1447 VTAIL.n630 VTAIL.n629 11.249
R1448 VTAIL.n576 VTAIL.n494 11.249
R1449 VTAIL.n563 VTAIL.n504 11.249
R1450 VTAIL.n532 VTAIL.n531 11.249
R1451 VTAIL.n478 VTAIL.n396 11.249
R1452 VTAIL.n465 VTAIL.n406 11.249
R1453 VTAIL.n434 VTAIL.n433 11.249
R1454 VTAIL.n380 VTAIL.n298 11.249
R1455 VTAIL.n367 VTAIL.n308 11.249
R1456 VTAIL.n336 VTAIL.n335 11.249
R1457 VTAIL.n729 VTAIL.n712 10.4732
R1458 VTAIL.n754 VTAIL.n753 10.4732
R1459 VTAIL.n776 VTAIL.n775 10.4732
R1460 VTAIL.n43 VTAIL.n26 10.4732
R1461 VTAIL.n68 VTAIL.n67 10.4732
R1462 VTAIL.n90 VTAIL.n89 10.4732
R1463 VTAIL.n141 VTAIL.n124 10.4732
R1464 VTAIL.n166 VTAIL.n165 10.4732
R1465 VTAIL.n188 VTAIL.n187 10.4732
R1466 VTAIL.n239 VTAIL.n222 10.4732
R1467 VTAIL.n264 VTAIL.n263 10.4732
R1468 VTAIL.n286 VTAIL.n285 10.4732
R1469 VTAIL.n678 VTAIL.n677 10.4732
R1470 VTAIL.n658 VTAIL.n657 10.4732
R1471 VTAIL.n633 VTAIL.n616 10.4732
R1472 VTAIL.n580 VTAIL.n579 10.4732
R1473 VTAIL.n560 VTAIL.n559 10.4732
R1474 VTAIL.n535 VTAIL.n518 10.4732
R1475 VTAIL.n482 VTAIL.n481 10.4732
R1476 VTAIL.n462 VTAIL.n461 10.4732
R1477 VTAIL.n437 VTAIL.n420 10.4732
R1478 VTAIL.n384 VTAIL.n383 10.4732
R1479 VTAIL.n364 VTAIL.n363 10.4732
R1480 VTAIL.n339 VTAIL.n322 10.4732
R1481 VTAIL.n730 VTAIL.n710 9.69747
R1482 VTAIL.n750 VTAIL.n700 9.69747
R1483 VTAIL.n779 VTAIL.n688 9.69747
R1484 VTAIL.n44 VTAIL.n24 9.69747
R1485 VTAIL.n64 VTAIL.n14 9.69747
R1486 VTAIL.n93 VTAIL.n2 9.69747
R1487 VTAIL.n142 VTAIL.n122 9.69747
R1488 VTAIL.n162 VTAIL.n112 9.69747
R1489 VTAIL.n191 VTAIL.n100 9.69747
R1490 VTAIL.n240 VTAIL.n220 9.69747
R1491 VTAIL.n260 VTAIL.n210 9.69747
R1492 VTAIL.n289 VTAIL.n198 9.69747
R1493 VTAIL.n681 VTAIL.n590 9.69747
R1494 VTAIL.n654 VTAIL.n604 9.69747
R1495 VTAIL.n634 VTAIL.n614 9.69747
R1496 VTAIL.n583 VTAIL.n492 9.69747
R1497 VTAIL.n556 VTAIL.n506 9.69747
R1498 VTAIL.n536 VTAIL.n516 9.69747
R1499 VTAIL.n485 VTAIL.n394 9.69747
R1500 VTAIL.n458 VTAIL.n408 9.69747
R1501 VTAIL.n438 VTAIL.n418 9.69747
R1502 VTAIL.n387 VTAIL.n296 9.69747
R1503 VTAIL.n360 VTAIL.n310 9.69747
R1504 VTAIL.n340 VTAIL.n320 9.69747
R1505 VTAIL.n782 VTAIL.n781 9.45567
R1506 VTAIL.n96 VTAIL.n95 9.45567
R1507 VTAIL.n194 VTAIL.n193 9.45567
R1508 VTAIL.n292 VTAIL.n291 9.45567
R1509 VTAIL.n684 VTAIL.n683 9.45567
R1510 VTAIL.n586 VTAIL.n585 9.45567
R1511 VTAIL.n488 VTAIL.n487 9.45567
R1512 VTAIL.n390 VTAIL.n389 9.45567
R1513 VTAIL.n781 VTAIL.n780 9.3005
R1514 VTAIL.n688 VTAIL.n687 9.3005
R1515 VTAIL.n775 VTAIL.n774 9.3005
R1516 VTAIL.n773 VTAIL.n772 9.3005
R1517 VTAIL.n692 VTAIL.n691 9.3005
R1518 VTAIL.n767 VTAIL.n766 9.3005
R1519 VTAIL.n739 VTAIL.n738 9.3005
R1520 VTAIL.n708 VTAIL.n707 9.3005
R1521 VTAIL.n733 VTAIL.n732 9.3005
R1522 VTAIL.n731 VTAIL.n730 9.3005
R1523 VTAIL.n712 VTAIL.n711 9.3005
R1524 VTAIL.n725 VTAIL.n724 9.3005
R1525 VTAIL.n723 VTAIL.n722 9.3005
R1526 VTAIL.n716 VTAIL.n715 9.3005
R1527 VTAIL.n741 VTAIL.n740 9.3005
R1528 VTAIL.n704 VTAIL.n703 9.3005
R1529 VTAIL.n747 VTAIL.n746 9.3005
R1530 VTAIL.n749 VTAIL.n748 9.3005
R1531 VTAIL.n700 VTAIL.n699 9.3005
R1532 VTAIL.n755 VTAIL.n754 9.3005
R1533 VTAIL.n757 VTAIL.n756 9.3005
R1534 VTAIL.n758 VTAIL.n695 9.3005
R1535 VTAIL.n765 VTAIL.n764 9.3005
R1536 VTAIL.n95 VTAIL.n94 9.3005
R1537 VTAIL.n2 VTAIL.n1 9.3005
R1538 VTAIL.n89 VTAIL.n88 9.3005
R1539 VTAIL.n87 VTAIL.n86 9.3005
R1540 VTAIL.n6 VTAIL.n5 9.3005
R1541 VTAIL.n81 VTAIL.n80 9.3005
R1542 VTAIL.n53 VTAIL.n52 9.3005
R1543 VTAIL.n22 VTAIL.n21 9.3005
R1544 VTAIL.n47 VTAIL.n46 9.3005
R1545 VTAIL.n45 VTAIL.n44 9.3005
R1546 VTAIL.n26 VTAIL.n25 9.3005
R1547 VTAIL.n39 VTAIL.n38 9.3005
R1548 VTAIL.n37 VTAIL.n36 9.3005
R1549 VTAIL.n30 VTAIL.n29 9.3005
R1550 VTAIL.n55 VTAIL.n54 9.3005
R1551 VTAIL.n18 VTAIL.n17 9.3005
R1552 VTAIL.n61 VTAIL.n60 9.3005
R1553 VTAIL.n63 VTAIL.n62 9.3005
R1554 VTAIL.n14 VTAIL.n13 9.3005
R1555 VTAIL.n69 VTAIL.n68 9.3005
R1556 VTAIL.n71 VTAIL.n70 9.3005
R1557 VTAIL.n72 VTAIL.n9 9.3005
R1558 VTAIL.n79 VTAIL.n78 9.3005
R1559 VTAIL.n193 VTAIL.n192 9.3005
R1560 VTAIL.n100 VTAIL.n99 9.3005
R1561 VTAIL.n187 VTAIL.n186 9.3005
R1562 VTAIL.n185 VTAIL.n184 9.3005
R1563 VTAIL.n104 VTAIL.n103 9.3005
R1564 VTAIL.n179 VTAIL.n178 9.3005
R1565 VTAIL.n151 VTAIL.n150 9.3005
R1566 VTAIL.n120 VTAIL.n119 9.3005
R1567 VTAIL.n145 VTAIL.n144 9.3005
R1568 VTAIL.n143 VTAIL.n142 9.3005
R1569 VTAIL.n124 VTAIL.n123 9.3005
R1570 VTAIL.n137 VTAIL.n136 9.3005
R1571 VTAIL.n135 VTAIL.n134 9.3005
R1572 VTAIL.n128 VTAIL.n127 9.3005
R1573 VTAIL.n153 VTAIL.n152 9.3005
R1574 VTAIL.n116 VTAIL.n115 9.3005
R1575 VTAIL.n159 VTAIL.n158 9.3005
R1576 VTAIL.n161 VTAIL.n160 9.3005
R1577 VTAIL.n112 VTAIL.n111 9.3005
R1578 VTAIL.n167 VTAIL.n166 9.3005
R1579 VTAIL.n169 VTAIL.n168 9.3005
R1580 VTAIL.n170 VTAIL.n107 9.3005
R1581 VTAIL.n177 VTAIL.n176 9.3005
R1582 VTAIL.n291 VTAIL.n290 9.3005
R1583 VTAIL.n198 VTAIL.n197 9.3005
R1584 VTAIL.n285 VTAIL.n284 9.3005
R1585 VTAIL.n283 VTAIL.n282 9.3005
R1586 VTAIL.n202 VTAIL.n201 9.3005
R1587 VTAIL.n277 VTAIL.n276 9.3005
R1588 VTAIL.n249 VTAIL.n248 9.3005
R1589 VTAIL.n218 VTAIL.n217 9.3005
R1590 VTAIL.n243 VTAIL.n242 9.3005
R1591 VTAIL.n241 VTAIL.n240 9.3005
R1592 VTAIL.n222 VTAIL.n221 9.3005
R1593 VTAIL.n235 VTAIL.n234 9.3005
R1594 VTAIL.n233 VTAIL.n232 9.3005
R1595 VTAIL.n226 VTAIL.n225 9.3005
R1596 VTAIL.n251 VTAIL.n250 9.3005
R1597 VTAIL.n214 VTAIL.n213 9.3005
R1598 VTAIL.n257 VTAIL.n256 9.3005
R1599 VTAIL.n259 VTAIL.n258 9.3005
R1600 VTAIL.n210 VTAIL.n209 9.3005
R1601 VTAIL.n265 VTAIL.n264 9.3005
R1602 VTAIL.n267 VTAIL.n266 9.3005
R1603 VTAIL.n268 VTAIL.n205 9.3005
R1604 VTAIL.n275 VTAIL.n274 9.3005
R1605 VTAIL.n608 VTAIL.n607 9.3005
R1606 VTAIL.n651 VTAIL.n650 9.3005
R1607 VTAIL.n653 VTAIL.n652 9.3005
R1608 VTAIL.n604 VTAIL.n603 9.3005
R1609 VTAIL.n659 VTAIL.n658 9.3005
R1610 VTAIL.n661 VTAIL.n660 9.3005
R1611 VTAIL.n599 VTAIL.n597 9.3005
R1612 VTAIL.n667 VTAIL.n666 9.3005
R1613 VTAIL.n683 VTAIL.n682 9.3005
R1614 VTAIL.n590 VTAIL.n589 9.3005
R1615 VTAIL.n677 VTAIL.n676 9.3005
R1616 VTAIL.n675 VTAIL.n674 9.3005
R1617 VTAIL.n594 VTAIL.n593 9.3005
R1618 VTAIL.n669 VTAIL.n668 9.3005
R1619 VTAIL.n645 VTAIL.n644 9.3005
R1620 VTAIL.n643 VTAIL.n642 9.3005
R1621 VTAIL.n612 VTAIL.n611 9.3005
R1622 VTAIL.n637 VTAIL.n636 9.3005
R1623 VTAIL.n635 VTAIL.n634 9.3005
R1624 VTAIL.n616 VTAIL.n615 9.3005
R1625 VTAIL.n629 VTAIL.n628 9.3005
R1626 VTAIL.n627 VTAIL.n626 9.3005
R1627 VTAIL.n620 VTAIL.n619 9.3005
R1628 VTAIL.n510 VTAIL.n509 9.3005
R1629 VTAIL.n553 VTAIL.n552 9.3005
R1630 VTAIL.n555 VTAIL.n554 9.3005
R1631 VTAIL.n506 VTAIL.n505 9.3005
R1632 VTAIL.n561 VTAIL.n560 9.3005
R1633 VTAIL.n563 VTAIL.n562 9.3005
R1634 VTAIL.n501 VTAIL.n499 9.3005
R1635 VTAIL.n569 VTAIL.n568 9.3005
R1636 VTAIL.n585 VTAIL.n584 9.3005
R1637 VTAIL.n492 VTAIL.n491 9.3005
R1638 VTAIL.n579 VTAIL.n578 9.3005
R1639 VTAIL.n577 VTAIL.n576 9.3005
R1640 VTAIL.n496 VTAIL.n495 9.3005
R1641 VTAIL.n571 VTAIL.n570 9.3005
R1642 VTAIL.n547 VTAIL.n546 9.3005
R1643 VTAIL.n545 VTAIL.n544 9.3005
R1644 VTAIL.n514 VTAIL.n513 9.3005
R1645 VTAIL.n539 VTAIL.n538 9.3005
R1646 VTAIL.n537 VTAIL.n536 9.3005
R1647 VTAIL.n518 VTAIL.n517 9.3005
R1648 VTAIL.n531 VTAIL.n530 9.3005
R1649 VTAIL.n529 VTAIL.n528 9.3005
R1650 VTAIL.n522 VTAIL.n521 9.3005
R1651 VTAIL.n412 VTAIL.n411 9.3005
R1652 VTAIL.n455 VTAIL.n454 9.3005
R1653 VTAIL.n457 VTAIL.n456 9.3005
R1654 VTAIL.n408 VTAIL.n407 9.3005
R1655 VTAIL.n463 VTAIL.n462 9.3005
R1656 VTAIL.n465 VTAIL.n464 9.3005
R1657 VTAIL.n403 VTAIL.n401 9.3005
R1658 VTAIL.n471 VTAIL.n470 9.3005
R1659 VTAIL.n487 VTAIL.n486 9.3005
R1660 VTAIL.n394 VTAIL.n393 9.3005
R1661 VTAIL.n481 VTAIL.n480 9.3005
R1662 VTAIL.n479 VTAIL.n478 9.3005
R1663 VTAIL.n398 VTAIL.n397 9.3005
R1664 VTAIL.n473 VTAIL.n472 9.3005
R1665 VTAIL.n449 VTAIL.n448 9.3005
R1666 VTAIL.n447 VTAIL.n446 9.3005
R1667 VTAIL.n416 VTAIL.n415 9.3005
R1668 VTAIL.n441 VTAIL.n440 9.3005
R1669 VTAIL.n439 VTAIL.n438 9.3005
R1670 VTAIL.n420 VTAIL.n419 9.3005
R1671 VTAIL.n433 VTAIL.n432 9.3005
R1672 VTAIL.n431 VTAIL.n430 9.3005
R1673 VTAIL.n424 VTAIL.n423 9.3005
R1674 VTAIL.n314 VTAIL.n313 9.3005
R1675 VTAIL.n357 VTAIL.n356 9.3005
R1676 VTAIL.n359 VTAIL.n358 9.3005
R1677 VTAIL.n310 VTAIL.n309 9.3005
R1678 VTAIL.n365 VTAIL.n364 9.3005
R1679 VTAIL.n367 VTAIL.n366 9.3005
R1680 VTAIL.n305 VTAIL.n303 9.3005
R1681 VTAIL.n373 VTAIL.n372 9.3005
R1682 VTAIL.n389 VTAIL.n388 9.3005
R1683 VTAIL.n296 VTAIL.n295 9.3005
R1684 VTAIL.n383 VTAIL.n382 9.3005
R1685 VTAIL.n381 VTAIL.n380 9.3005
R1686 VTAIL.n300 VTAIL.n299 9.3005
R1687 VTAIL.n375 VTAIL.n374 9.3005
R1688 VTAIL.n351 VTAIL.n350 9.3005
R1689 VTAIL.n349 VTAIL.n348 9.3005
R1690 VTAIL.n318 VTAIL.n317 9.3005
R1691 VTAIL.n343 VTAIL.n342 9.3005
R1692 VTAIL.n341 VTAIL.n340 9.3005
R1693 VTAIL.n322 VTAIL.n321 9.3005
R1694 VTAIL.n335 VTAIL.n334 9.3005
R1695 VTAIL.n333 VTAIL.n332 9.3005
R1696 VTAIL.n326 VTAIL.n325 9.3005
R1697 VTAIL.n734 VTAIL.n733 8.92171
R1698 VTAIL.n749 VTAIL.n702 8.92171
R1699 VTAIL.n780 VTAIL.n686 8.92171
R1700 VTAIL.n48 VTAIL.n47 8.92171
R1701 VTAIL.n63 VTAIL.n16 8.92171
R1702 VTAIL.n94 VTAIL.n0 8.92171
R1703 VTAIL.n146 VTAIL.n145 8.92171
R1704 VTAIL.n161 VTAIL.n114 8.92171
R1705 VTAIL.n192 VTAIL.n98 8.92171
R1706 VTAIL.n244 VTAIL.n243 8.92171
R1707 VTAIL.n259 VTAIL.n212 8.92171
R1708 VTAIL.n290 VTAIL.n196 8.92171
R1709 VTAIL.n682 VTAIL.n588 8.92171
R1710 VTAIL.n653 VTAIL.n606 8.92171
R1711 VTAIL.n638 VTAIL.n637 8.92171
R1712 VTAIL.n584 VTAIL.n490 8.92171
R1713 VTAIL.n555 VTAIL.n508 8.92171
R1714 VTAIL.n540 VTAIL.n539 8.92171
R1715 VTAIL.n486 VTAIL.n392 8.92171
R1716 VTAIL.n457 VTAIL.n410 8.92171
R1717 VTAIL.n442 VTAIL.n441 8.92171
R1718 VTAIL.n388 VTAIL.n294 8.92171
R1719 VTAIL.n359 VTAIL.n312 8.92171
R1720 VTAIL.n344 VTAIL.n343 8.92171
R1721 VTAIL.n737 VTAIL.n708 8.14595
R1722 VTAIL.n746 VTAIL.n745 8.14595
R1723 VTAIL.n51 VTAIL.n22 8.14595
R1724 VTAIL.n60 VTAIL.n59 8.14595
R1725 VTAIL.n149 VTAIL.n120 8.14595
R1726 VTAIL.n158 VTAIL.n157 8.14595
R1727 VTAIL.n247 VTAIL.n218 8.14595
R1728 VTAIL.n256 VTAIL.n255 8.14595
R1729 VTAIL.n650 VTAIL.n649 8.14595
R1730 VTAIL.n641 VTAIL.n612 8.14595
R1731 VTAIL.n552 VTAIL.n551 8.14595
R1732 VTAIL.n543 VTAIL.n514 8.14595
R1733 VTAIL.n454 VTAIL.n453 8.14595
R1734 VTAIL.n445 VTAIL.n416 8.14595
R1735 VTAIL.n356 VTAIL.n355 8.14595
R1736 VTAIL.n347 VTAIL.n318 8.14595
R1737 VTAIL.n738 VTAIL.n706 7.3702
R1738 VTAIL.n742 VTAIL.n704 7.3702
R1739 VTAIL.n52 VTAIL.n20 7.3702
R1740 VTAIL.n56 VTAIL.n18 7.3702
R1741 VTAIL.n150 VTAIL.n118 7.3702
R1742 VTAIL.n154 VTAIL.n116 7.3702
R1743 VTAIL.n248 VTAIL.n216 7.3702
R1744 VTAIL.n252 VTAIL.n214 7.3702
R1745 VTAIL.n646 VTAIL.n608 7.3702
R1746 VTAIL.n642 VTAIL.n610 7.3702
R1747 VTAIL.n548 VTAIL.n510 7.3702
R1748 VTAIL.n544 VTAIL.n512 7.3702
R1749 VTAIL.n450 VTAIL.n412 7.3702
R1750 VTAIL.n446 VTAIL.n414 7.3702
R1751 VTAIL.n352 VTAIL.n314 7.3702
R1752 VTAIL.n348 VTAIL.n316 7.3702
R1753 VTAIL.n741 VTAIL.n706 6.59444
R1754 VTAIL.n742 VTAIL.n741 6.59444
R1755 VTAIL.n55 VTAIL.n20 6.59444
R1756 VTAIL.n56 VTAIL.n55 6.59444
R1757 VTAIL.n153 VTAIL.n118 6.59444
R1758 VTAIL.n154 VTAIL.n153 6.59444
R1759 VTAIL.n251 VTAIL.n216 6.59444
R1760 VTAIL.n252 VTAIL.n251 6.59444
R1761 VTAIL.n646 VTAIL.n645 6.59444
R1762 VTAIL.n645 VTAIL.n610 6.59444
R1763 VTAIL.n548 VTAIL.n547 6.59444
R1764 VTAIL.n547 VTAIL.n512 6.59444
R1765 VTAIL.n450 VTAIL.n449 6.59444
R1766 VTAIL.n449 VTAIL.n414 6.59444
R1767 VTAIL.n352 VTAIL.n351 6.59444
R1768 VTAIL.n351 VTAIL.n316 6.59444
R1769 VTAIL.n738 VTAIL.n737 5.81868
R1770 VTAIL.n745 VTAIL.n704 5.81868
R1771 VTAIL.n52 VTAIL.n51 5.81868
R1772 VTAIL.n59 VTAIL.n18 5.81868
R1773 VTAIL.n150 VTAIL.n149 5.81868
R1774 VTAIL.n157 VTAIL.n116 5.81868
R1775 VTAIL.n248 VTAIL.n247 5.81868
R1776 VTAIL.n255 VTAIL.n214 5.81868
R1777 VTAIL.n649 VTAIL.n608 5.81868
R1778 VTAIL.n642 VTAIL.n641 5.81868
R1779 VTAIL.n551 VTAIL.n510 5.81868
R1780 VTAIL.n544 VTAIL.n543 5.81868
R1781 VTAIL.n453 VTAIL.n412 5.81868
R1782 VTAIL.n446 VTAIL.n445 5.81868
R1783 VTAIL.n355 VTAIL.n314 5.81868
R1784 VTAIL.n348 VTAIL.n347 5.81868
R1785 VTAIL.n734 VTAIL.n708 5.04292
R1786 VTAIL.n746 VTAIL.n702 5.04292
R1787 VTAIL.n782 VTAIL.n686 5.04292
R1788 VTAIL.n48 VTAIL.n22 5.04292
R1789 VTAIL.n60 VTAIL.n16 5.04292
R1790 VTAIL.n96 VTAIL.n0 5.04292
R1791 VTAIL.n146 VTAIL.n120 5.04292
R1792 VTAIL.n158 VTAIL.n114 5.04292
R1793 VTAIL.n194 VTAIL.n98 5.04292
R1794 VTAIL.n244 VTAIL.n218 5.04292
R1795 VTAIL.n256 VTAIL.n212 5.04292
R1796 VTAIL.n292 VTAIL.n196 5.04292
R1797 VTAIL.n684 VTAIL.n588 5.04292
R1798 VTAIL.n650 VTAIL.n606 5.04292
R1799 VTAIL.n638 VTAIL.n612 5.04292
R1800 VTAIL.n586 VTAIL.n490 5.04292
R1801 VTAIL.n552 VTAIL.n508 5.04292
R1802 VTAIL.n540 VTAIL.n514 5.04292
R1803 VTAIL.n488 VTAIL.n392 5.04292
R1804 VTAIL.n454 VTAIL.n410 5.04292
R1805 VTAIL.n442 VTAIL.n416 5.04292
R1806 VTAIL.n390 VTAIL.n294 5.04292
R1807 VTAIL.n356 VTAIL.n312 5.04292
R1808 VTAIL.n344 VTAIL.n318 5.04292
R1809 VTAIL.n733 VTAIL.n710 4.26717
R1810 VTAIL.n750 VTAIL.n749 4.26717
R1811 VTAIL.n780 VTAIL.n779 4.26717
R1812 VTAIL.n47 VTAIL.n24 4.26717
R1813 VTAIL.n64 VTAIL.n63 4.26717
R1814 VTAIL.n94 VTAIL.n93 4.26717
R1815 VTAIL.n145 VTAIL.n122 4.26717
R1816 VTAIL.n162 VTAIL.n161 4.26717
R1817 VTAIL.n192 VTAIL.n191 4.26717
R1818 VTAIL.n243 VTAIL.n220 4.26717
R1819 VTAIL.n260 VTAIL.n259 4.26717
R1820 VTAIL.n290 VTAIL.n289 4.26717
R1821 VTAIL.n682 VTAIL.n681 4.26717
R1822 VTAIL.n654 VTAIL.n653 4.26717
R1823 VTAIL.n637 VTAIL.n614 4.26717
R1824 VTAIL.n584 VTAIL.n583 4.26717
R1825 VTAIL.n556 VTAIL.n555 4.26717
R1826 VTAIL.n539 VTAIL.n516 4.26717
R1827 VTAIL.n486 VTAIL.n485 4.26717
R1828 VTAIL.n458 VTAIL.n457 4.26717
R1829 VTAIL.n441 VTAIL.n418 4.26717
R1830 VTAIL.n388 VTAIL.n387 4.26717
R1831 VTAIL.n360 VTAIL.n359 4.26717
R1832 VTAIL.n343 VTAIL.n320 4.26717
R1833 VTAIL.n717 VTAIL.n715 3.70982
R1834 VTAIL.n31 VTAIL.n29 3.70982
R1835 VTAIL.n129 VTAIL.n127 3.70982
R1836 VTAIL.n227 VTAIL.n225 3.70982
R1837 VTAIL.n621 VTAIL.n619 3.70982
R1838 VTAIL.n523 VTAIL.n521 3.70982
R1839 VTAIL.n425 VTAIL.n423 3.70982
R1840 VTAIL.n327 VTAIL.n325 3.70982
R1841 VTAIL.n730 VTAIL.n729 3.49141
R1842 VTAIL.n753 VTAIL.n700 3.49141
R1843 VTAIL.n776 VTAIL.n688 3.49141
R1844 VTAIL.n44 VTAIL.n43 3.49141
R1845 VTAIL.n67 VTAIL.n14 3.49141
R1846 VTAIL.n90 VTAIL.n2 3.49141
R1847 VTAIL.n142 VTAIL.n141 3.49141
R1848 VTAIL.n165 VTAIL.n112 3.49141
R1849 VTAIL.n188 VTAIL.n100 3.49141
R1850 VTAIL.n240 VTAIL.n239 3.49141
R1851 VTAIL.n263 VTAIL.n210 3.49141
R1852 VTAIL.n286 VTAIL.n198 3.49141
R1853 VTAIL.n678 VTAIL.n590 3.49141
R1854 VTAIL.n657 VTAIL.n604 3.49141
R1855 VTAIL.n634 VTAIL.n633 3.49141
R1856 VTAIL.n580 VTAIL.n492 3.49141
R1857 VTAIL.n559 VTAIL.n506 3.49141
R1858 VTAIL.n536 VTAIL.n535 3.49141
R1859 VTAIL.n482 VTAIL.n394 3.49141
R1860 VTAIL.n461 VTAIL.n408 3.49141
R1861 VTAIL.n438 VTAIL.n437 3.49141
R1862 VTAIL.n384 VTAIL.n296 3.49141
R1863 VTAIL.n363 VTAIL.n310 3.49141
R1864 VTAIL.n340 VTAIL.n339 3.49141
R1865 VTAIL.n726 VTAIL.n712 2.71565
R1866 VTAIL.n754 VTAIL.n698 2.71565
R1867 VTAIL.n775 VTAIL.n690 2.71565
R1868 VTAIL.n40 VTAIL.n26 2.71565
R1869 VTAIL.n68 VTAIL.n12 2.71565
R1870 VTAIL.n89 VTAIL.n4 2.71565
R1871 VTAIL.n138 VTAIL.n124 2.71565
R1872 VTAIL.n166 VTAIL.n110 2.71565
R1873 VTAIL.n187 VTAIL.n102 2.71565
R1874 VTAIL.n236 VTAIL.n222 2.71565
R1875 VTAIL.n264 VTAIL.n208 2.71565
R1876 VTAIL.n285 VTAIL.n200 2.71565
R1877 VTAIL.n677 VTAIL.n592 2.71565
R1878 VTAIL.n658 VTAIL.n602 2.71565
R1879 VTAIL.n630 VTAIL.n616 2.71565
R1880 VTAIL.n579 VTAIL.n494 2.71565
R1881 VTAIL.n560 VTAIL.n504 2.71565
R1882 VTAIL.n532 VTAIL.n518 2.71565
R1883 VTAIL.n481 VTAIL.n396 2.71565
R1884 VTAIL.n462 VTAIL.n406 2.71565
R1885 VTAIL.n434 VTAIL.n420 2.71565
R1886 VTAIL.n383 VTAIL.n298 2.71565
R1887 VTAIL.n364 VTAIL.n308 2.71565
R1888 VTAIL.n336 VTAIL.n322 2.71565
R1889 VTAIL.n725 VTAIL.n714 1.93989
R1890 VTAIL.n759 VTAIL.n757 1.93989
R1891 VTAIL.n772 VTAIL.n771 1.93989
R1892 VTAIL.n39 VTAIL.n28 1.93989
R1893 VTAIL.n73 VTAIL.n71 1.93989
R1894 VTAIL.n86 VTAIL.n85 1.93989
R1895 VTAIL.n137 VTAIL.n126 1.93989
R1896 VTAIL.n171 VTAIL.n169 1.93989
R1897 VTAIL.n184 VTAIL.n183 1.93989
R1898 VTAIL.n235 VTAIL.n224 1.93989
R1899 VTAIL.n269 VTAIL.n267 1.93989
R1900 VTAIL.n282 VTAIL.n281 1.93989
R1901 VTAIL.n674 VTAIL.n673 1.93989
R1902 VTAIL.n662 VTAIL.n661 1.93989
R1903 VTAIL.n629 VTAIL.n618 1.93989
R1904 VTAIL.n576 VTAIL.n575 1.93989
R1905 VTAIL.n564 VTAIL.n563 1.93989
R1906 VTAIL.n531 VTAIL.n520 1.93989
R1907 VTAIL.n478 VTAIL.n477 1.93989
R1908 VTAIL.n466 VTAIL.n465 1.93989
R1909 VTAIL.n433 VTAIL.n422 1.93989
R1910 VTAIL.n380 VTAIL.n379 1.93989
R1911 VTAIL.n368 VTAIL.n367 1.93989
R1912 VTAIL.n335 VTAIL.n324 1.93989
R1913 VTAIL.n722 VTAIL.n721 1.16414
R1914 VTAIL.n758 VTAIL.n696 1.16414
R1915 VTAIL.n768 VTAIL.n692 1.16414
R1916 VTAIL.n36 VTAIL.n35 1.16414
R1917 VTAIL.n72 VTAIL.n10 1.16414
R1918 VTAIL.n82 VTAIL.n6 1.16414
R1919 VTAIL.n134 VTAIL.n133 1.16414
R1920 VTAIL.n170 VTAIL.n108 1.16414
R1921 VTAIL.n180 VTAIL.n104 1.16414
R1922 VTAIL.n232 VTAIL.n231 1.16414
R1923 VTAIL.n268 VTAIL.n206 1.16414
R1924 VTAIL.n278 VTAIL.n202 1.16414
R1925 VTAIL.n670 VTAIL.n594 1.16414
R1926 VTAIL.n665 VTAIL.n599 1.16414
R1927 VTAIL.n626 VTAIL.n625 1.16414
R1928 VTAIL.n572 VTAIL.n496 1.16414
R1929 VTAIL.n567 VTAIL.n501 1.16414
R1930 VTAIL.n528 VTAIL.n527 1.16414
R1931 VTAIL.n474 VTAIL.n398 1.16414
R1932 VTAIL.n469 VTAIL.n403 1.16414
R1933 VTAIL.n430 VTAIL.n429 1.16414
R1934 VTAIL.n376 VTAIL.n300 1.16414
R1935 VTAIL.n371 VTAIL.n305 1.16414
R1936 VTAIL.n332 VTAIL.n331 1.16414
R1937 VTAIL.n489 VTAIL.n391 0.517741
R1938 VTAIL.n685 VTAIL.n587 0.517741
R1939 VTAIL.n293 VTAIL.n195 0.517741
R1940 VTAIL.n587 VTAIL.n489 0.470328
R1941 VTAIL.n195 VTAIL.n97 0.470328
R1942 VTAIL.n718 VTAIL.n716 0.388379
R1943 VTAIL.n764 VTAIL.n763 0.388379
R1944 VTAIL.n767 VTAIL.n694 0.388379
R1945 VTAIL.n32 VTAIL.n30 0.388379
R1946 VTAIL.n78 VTAIL.n77 0.388379
R1947 VTAIL.n81 VTAIL.n8 0.388379
R1948 VTAIL.n130 VTAIL.n128 0.388379
R1949 VTAIL.n176 VTAIL.n175 0.388379
R1950 VTAIL.n179 VTAIL.n106 0.388379
R1951 VTAIL.n228 VTAIL.n226 0.388379
R1952 VTAIL.n274 VTAIL.n273 0.388379
R1953 VTAIL.n277 VTAIL.n204 0.388379
R1954 VTAIL.n669 VTAIL.n596 0.388379
R1955 VTAIL.n666 VTAIL.n598 0.388379
R1956 VTAIL.n622 VTAIL.n620 0.388379
R1957 VTAIL.n571 VTAIL.n498 0.388379
R1958 VTAIL.n568 VTAIL.n500 0.388379
R1959 VTAIL.n524 VTAIL.n522 0.388379
R1960 VTAIL.n473 VTAIL.n400 0.388379
R1961 VTAIL.n470 VTAIL.n402 0.388379
R1962 VTAIL.n426 VTAIL.n424 0.388379
R1963 VTAIL.n375 VTAIL.n302 0.388379
R1964 VTAIL.n372 VTAIL.n304 0.388379
R1965 VTAIL.n328 VTAIL.n326 0.388379
R1966 VTAIL VTAIL.n97 0.31731
R1967 VTAIL VTAIL.n783 0.200931
R1968 VTAIL.n723 VTAIL.n715 0.155672
R1969 VTAIL.n724 VTAIL.n723 0.155672
R1970 VTAIL.n724 VTAIL.n711 0.155672
R1971 VTAIL.n731 VTAIL.n711 0.155672
R1972 VTAIL.n732 VTAIL.n731 0.155672
R1973 VTAIL.n732 VTAIL.n707 0.155672
R1974 VTAIL.n739 VTAIL.n707 0.155672
R1975 VTAIL.n740 VTAIL.n739 0.155672
R1976 VTAIL.n740 VTAIL.n703 0.155672
R1977 VTAIL.n747 VTAIL.n703 0.155672
R1978 VTAIL.n748 VTAIL.n747 0.155672
R1979 VTAIL.n748 VTAIL.n699 0.155672
R1980 VTAIL.n755 VTAIL.n699 0.155672
R1981 VTAIL.n756 VTAIL.n755 0.155672
R1982 VTAIL.n756 VTAIL.n695 0.155672
R1983 VTAIL.n765 VTAIL.n695 0.155672
R1984 VTAIL.n766 VTAIL.n765 0.155672
R1985 VTAIL.n766 VTAIL.n691 0.155672
R1986 VTAIL.n773 VTAIL.n691 0.155672
R1987 VTAIL.n774 VTAIL.n773 0.155672
R1988 VTAIL.n774 VTAIL.n687 0.155672
R1989 VTAIL.n781 VTAIL.n687 0.155672
R1990 VTAIL.n37 VTAIL.n29 0.155672
R1991 VTAIL.n38 VTAIL.n37 0.155672
R1992 VTAIL.n38 VTAIL.n25 0.155672
R1993 VTAIL.n45 VTAIL.n25 0.155672
R1994 VTAIL.n46 VTAIL.n45 0.155672
R1995 VTAIL.n46 VTAIL.n21 0.155672
R1996 VTAIL.n53 VTAIL.n21 0.155672
R1997 VTAIL.n54 VTAIL.n53 0.155672
R1998 VTAIL.n54 VTAIL.n17 0.155672
R1999 VTAIL.n61 VTAIL.n17 0.155672
R2000 VTAIL.n62 VTAIL.n61 0.155672
R2001 VTAIL.n62 VTAIL.n13 0.155672
R2002 VTAIL.n69 VTAIL.n13 0.155672
R2003 VTAIL.n70 VTAIL.n69 0.155672
R2004 VTAIL.n70 VTAIL.n9 0.155672
R2005 VTAIL.n79 VTAIL.n9 0.155672
R2006 VTAIL.n80 VTAIL.n79 0.155672
R2007 VTAIL.n80 VTAIL.n5 0.155672
R2008 VTAIL.n87 VTAIL.n5 0.155672
R2009 VTAIL.n88 VTAIL.n87 0.155672
R2010 VTAIL.n88 VTAIL.n1 0.155672
R2011 VTAIL.n95 VTAIL.n1 0.155672
R2012 VTAIL.n135 VTAIL.n127 0.155672
R2013 VTAIL.n136 VTAIL.n135 0.155672
R2014 VTAIL.n136 VTAIL.n123 0.155672
R2015 VTAIL.n143 VTAIL.n123 0.155672
R2016 VTAIL.n144 VTAIL.n143 0.155672
R2017 VTAIL.n144 VTAIL.n119 0.155672
R2018 VTAIL.n151 VTAIL.n119 0.155672
R2019 VTAIL.n152 VTAIL.n151 0.155672
R2020 VTAIL.n152 VTAIL.n115 0.155672
R2021 VTAIL.n159 VTAIL.n115 0.155672
R2022 VTAIL.n160 VTAIL.n159 0.155672
R2023 VTAIL.n160 VTAIL.n111 0.155672
R2024 VTAIL.n167 VTAIL.n111 0.155672
R2025 VTAIL.n168 VTAIL.n167 0.155672
R2026 VTAIL.n168 VTAIL.n107 0.155672
R2027 VTAIL.n177 VTAIL.n107 0.155672
R2028 VTAIL.n178 VTAIL.n177 0.155672
R2029 VTAIL.n178 VTAIL.n103 0.155672
R2030 VTAIL.n185 VTAIL.n103 0.155672
R2031 VTAIL.n186 VTAIL.n185 0.155672
R2032 VTAIL.n186 VTAIL.n99 0.155672
R2033 VTAIL.n193 VTAIL.n99 0.155672
R2034 VTAIL.n233 VTAIL.n225 0.155672
R2035 VTAIL.n234 VTAIL.n233 0.155672
R2036 VTAIL.n234 VTAIL.n221 0.155672
R2037 VTAIL.n241 VTAIL.n221 0.155672
R2038 VTAIL.n242 VTAIL.n241 0.155672
R2039 VTAIL.n242 VTAIL.n217 0.155672
R2040 VTAIL.n249 VTAIL.n217 0.155672
R2041 VTAIL.n250 VTAIL.n249 0.155672
R2042 VTAIL.n250 VTAIL.n213 0.155672
R2043 VTAIL.n257 VTAIL.n213 0.155672
R2044 VTAIL.n258 VTAIL.n257 0.155672
R2045 VTAIL.n258 VTAIL.n209 0.155672
R2046 VTAIL.n265 VTAIL.n209 0.155672
R2047 VTAIL.n266 VTAIL.n265 0.155672
R2048 VTAIL.n266 VTAIL.n205 0.155672
R2049 VTAIL.n275 VTAIL.n205 0.155672
R2050 VTAIL.n276 VTAIL.n275 0.155672
R2051 VTAIL.n276 VTAIL.n201 0.155672
R2052 VTAIL.n283 VTAIL.n201 0.155672
R2053 VTAIL.n284 VTAIL.n283 0.155672
R2054 VTAIL.n284 VTAIL.n197 0.155672
R2055 VTAIL.n291 VTAIL.n197 0.155672
R2056 VTAIL.n683 VTAIL.n589 0.155672
R2057 VTAIL.n676 VTAIL.n589 0.155672
R2058 VTAIL.n676 VTAIL.n675 0.155672
R2059 VTAIL.n675 VTAIL.n593 0.155672
R2060 VTAIL.n668 VTAIL.n593 0.155672
R2061 VTAIL.n668 VTAIL.n667 0.155672
R2062 VTAIL.n667 VTAIL.n597 0.155672
R2063 VTAIL.n660 VTAIL.n597 0.155672
R2064 VTAIL.n660 VTAIL.n659 0.155672
R2065 VTAIL.n659 VTAIL.n603 0.155672
R2066 VTAIL.n652 VTAIL.n603 0.155672
R2067 VTAIL.n652 VTAIL.n651 0.155672
R2068 VTAIL.n651 VTAIL.n607 0.155672
R2069 VTAIL.n644 VTAIL.n607 0.155672
R2070 VTAIL.n644 VTAIL.n643 0.155672
R2071 VTAIL.n643 VTAIL.n611 0.155672
R2072 VTAIL.n636 VTAIL.n611 0.155672
R2073 VTAIL.n636 VTAIL.n635 0.155672
R2074 VTAIL.n635 VTAIL.n615 0.155672
R2075 VTAIL.n628 VTAIL.n615 0.155672
R2076 VTAIL.n628 VTAIL.n627 0.155672
R2077 VTAIL.n627 VTAIL.n619 0.155672
R2078 VTAIL.n585 VTAIL.n491 0.155672
R2079 VTAIL.n578 VTAIL.n491 0.155672
R2080 VTAIL.n578 VTAIL.n577 0.155672
R2081 VTAIL.n577 VTAIL.n495 0.155672
R2082 VTAIL.n570 VTAIL.n495 0.155672
R2083 VTAIL.n570 VTAIL.n569 0.155672
R2084 VTAIL.n569 VTAIL.n499 0.155672
R2085 VTAIL.n562 VTAIL.n499 0.155672
R2086 VTAIL.n562 VTAIL.n561 0.155672
R2087 VTAIL.n561 VTAIL.n505 0.155672
R2088 VTAIL.n554 VTAIL.n505 0.155672
R2089 VTAIL.n554 VTAIL.n553 0.155672
R2090 VTAIL.n553 VTAIL.n509 0.155672
R2091 VTAIL.n546 VTAIL.n509 0.155672
R2092 VTAIL.n546 VTAIL.n545 0.155672
R2093 VTAIL.n545 VTAIL.n513 0.155672
R2094 VTAIL.n538 VTAIL.n513 0.155672
R2095 VTAIL.n538 VTAIL.n537 0.155672
R2096 VTAIL.n537 VTAIL.n517 0.155672
R2097 VTAIL.n530 VTAIL.n517 0.155672
R2098 VTAIL.n530 VTAIL.n529 0.155672
R2099 VTAIL.n529 VTAIL.n521 0.155672
R2100 VTAIL.n487 VTAIL.n393 0.155672
R2101 VTAIL.n480 VTAIL.n393 0.155672
R2102 VTAIL.n480 VTAIL.n479 0.155672
R2103 VTAIL.n479 VTAIL.n397 0.155672
R2104 VTAIL.n472 VTAIL.n397 0.155672
R2105 VTAIL.n472 VTAIL.n471 0.155672
R2106 VTAIL.n471 VTAIL.n401 0.155672
R2107 VTAIL.n464 VTAIL.n401 0.155672
R2108 VTAIL.n464 VTAIL.n463 0.155672
R2109 VTAIL.n463 VTAIL.n407 0.155672
R2110 VTAIL.n456 VTAIL.n407 0.155672
R2111 VTAIL.n456 VTAIL.n455 0.155672
R2112 VTAIL.n455 VTAIL.n411 0.155672
R2113 VTAIL.n448 VTAIL.n411 0.155672
R2114 VTAIL.n448 VTAIL.n447 0.155672
R2115 VTAIL.n447 VTAIL.n415 0.155672
R2116 VTAIL.n440 VTAIL.n415 0.155672
R2117 VTAIL.n440 VTAIL.n439 0.155672
R2118 VTAIL.n439 VTAIL.n419 0.155672
R2119 VTAIL.n432 VTAIL.n419 0.155672
R2120 VTAIL.n432 VTAIL.n431 0.155672
R2121 VTAIL.n431 VTAIL.n423 0.155672
R2122 VTAIL.n389 VTAIL.n295 0.155672
R2123 VTAIL.n382 VTAIL.n295 0.155672
R2124 VTAIL.n382 VTAIL.n381 0.155672
R2125 VTAIL.n381 VTAIL.n299 0.155672
R2126 VTAIL.n374 VTAIL.n299 0.155672
R2127 VTAIL.n374 VTAIL.n373 0.155672
R2128 VTAIL.n373 VTAIL.n303 0.155672
R2129 VTAIL.n366 VTAIL.n303 0.155672
R2130 VTAIL.n366 VTAIL.n365 0.155672
R2131 VTAIL.n365 VTAIL.n309 0.155672
R2132 VTAIL.n358 VTAIL.n309 0.155672
R2133 VTAIL.n358 VTAIL.n357 0.155672
R2134 VTAIL.n357 VTAIL.n313 0.155672
R2135 VTAIL.n350 VTAIL.n313 0.155672
R2136 VTAIL.n350 VTAIL.n349 0.155672
R2137 VTAIL.n349 VTAIL.n317 0.155672
R2138 VTAIL.n342 VTAIL.n317 0.155672
R2139 VTAIL.n342 VTAIL.n341 0.155672
R2140 VTAIL.n341 VTAIL.n321 0.155672
R2141 VTAIL.n334 VTAIL.n321 0.155672
R2142 VTAIL.n334 VTAIL.n333 0.155672
R2143 VTAIL.n333 VTAIL.n325 0.155672
R2144 VP.n1 VP.t0 1732.6
R2145 VP.n1 VP.t2 1732.6
R2146 VP.n0 VP.t1 1732.6
R2147 VP.n0 VP.t3 1732.6
R2148 VP.n2 VP.n0 204.718
R2149 VP.n2 VP.n1 161.3
R2150 VP VP.n2 0.0516364
R2151 VDD1 VDD1.n1 111.555
R2152 VDD1 VDD1.n0 70.6317
R2153 VDD1.n0 VDD1.t2 1.84737
R2154 VDD1.n0 VDD1.t0 1.84737
R2155 VDD1.n1 VDD1.t1 1.84737
R2156 VDD1.n1 VDD1.t3 1.84737
C0 VDD2 VTAIL 13.862401f
C1 VDD2 VP 0.246849f
C2 w_n1330_n4492# B 7.980649f
C3 VDD2 VN 2.76959f
C4 VDD1 w_n1330_n4492# 1.11109f
C5 w_n1330_n4492# VTAIL 5.79679f
C6 w_n1330_n4492# VP 2.09706f
C7 w_n1330_n4492# VN 1.93197f
C8 VDD2 w_n1330_n4492# 1.11732f
C9 VDD1 B 1.00061f
C10 VTAIL B 4.89351f
C11 VP B 0.98907f
C12 VN B 0.725965f
C13 VDD1 VTAIL 13.8238f
C14 VDD1 VP 2.86859f
C15 VDD1 VN 0.1477f
C16 VDD2 B 1.01623f
C17 VDD2 VDD1 0.472338f
C18 VP VTAIL 1.99194f
C19 VN VTAIL 1.97784f
C20 VP VN 5.54661f
C21 VDD2 VSUBS 0.765539f
C22 VDD1 VSUBS 6.626601f
C23 VTAIL VSUBS 0.919521f
C24 VN VSUBS 5.82916f
C25 VP VSUBS 1.285128f
C26 B VSUBS 2.727343f
C27 w_n1330_n4492# VSUBS 73.080795f
C28 VDD1.t2 VSUBS 0.478927f
C29 VDD1.t0 VSUBS 0.478927f
C30 VDD1.n0 VSUBS 3.97673f
C31 VDD1.t1 VSUBS 0.478927f
C32 VDD1.t3 VSUBS 0.478927f
C33 VDD1.n1 VSUBS 5.03579f
C34 VP.t1 VSUBS 0.869532f
C35 VP.t3 VSUBS 0.869532f
C36 VP.n0 VSUBS 1.26468f
C37 VP.t2 VSUBS 0.869532f
C38 VP.t0 VSUBS 0.869532f
C39 VP.n1 VSUBS 0.667285f
C40 VP.n2 VSUBS 5.06078f
C41 VTAIL.n0 VSUBS 0.025904f
C42 VTAIL.n1 VSUBS 0.023304f
C43 VTAIL.n2 VSUBS 0.012523f
C44 VTAIL.n3 VSUBS 0.029599f
C45 VTAIL.n4 VSUBS 0.013259f
C46 VTAIL.n5 VSUBS 0.023304f
C47 VTAIL.n6 VSUBS 0.012523f
C48 VTAIL.n7 VSUBS 0.029599f
C49 VTAIL.n8 VSUBS 0.012891f
C50 VTAIL.n9 VSUBS 0.023304f
C51 VTAIL.n10 VSUBS 0.013259f
C52 VTAIL.n11 VSUBS 0.029599f
C53 VTAIL.n12 VSUBS 0.013259f
C54 VTAIL.n13 VSUBS 0.023304f
C55 VTAIL.n14 VSUBS 0.012523f
C56 VTAIL.n15 VSUBS 0.029599f
C57 VTAIL.n16 VSUBS 0.013259f
C58 VTAIL.n17 VSUBS 0.023304f
C59 VTAIL.n18 VSUBS 0.012523f
C60 VTAIL.n19 VSUBS 0.029599f
C61 VTAIL.n20 VSUBS 0.013259f
C62 VTAIL.n21 VSUBS 0.023304f
C63 VTAIL.n22 VSUBS 0.012523f
C64 VTAIL.n23 VSUBS 0.029599f
C65 VTAIL.n24 VSUBS 0.013259f
C66 VTAIL.n25 VSUBS 0.023304f
C67 VTAIL.n26 VSUBS 0.012523f
C68 VTAIL.n27 VSUBS 0.029599f
C69 VTAIL.n28 VSUBS 0.013259f
C70 VTAIL.n29 VSUBS 1.76306f
C71 VTAIL.n30 VSUBS 0.012523f
C72 VTAIL.t7 VSUBS 0.063515f
C73 VTAIL.n31 VSUBS 0.182143f
C74 VTAIL.n32 VSUBS 0.018829f
C75 VTAIL.n33 VSUBS 0.022199f
C76 VTAIL.n34 VSUBS 0.029599f
C77 VTAIL.n35 VSUBS 0.013259f
C78 VTAIL.n36 VSUBS 0.012523f
C79 VTAIL.n37 VSUBS 0.023304f
C80 VTAIL.n38 VSUBS 0.023304f
C81 VTAIL.n39 VSUBS 0.012523f
C82 VTAIL.n40 VSUBS 0.013259f
C83 VTAIL.n41 VSUBS 0.029599f
C84 VTAIL.n42 VSUBS 0.029599f
C85 VTAIL.n43 VSUBS 0.013259f
C86 VTAIL.n44 VSUBS 0.012523f
C87 VTAIL.n45 VSUBS 0.023304f
C88 VTAIL.n46 VSUBS 0.023304f
C89 VTAIL.n47 VSUBS 0.012523f
C90 VTAIL.n48 VSUBS 0.013259f
C91 VTAIL.n49 VSUBS 0.029599f
C92 VTAIL.n50 VSUBS 0.029599f
C93 VTAIL.n51 VSUBS 0.013259f
C94 VTAIL.n52 VSUBS 0.012523f
C95 VTAIL.n53 VSUBS 0.023304f
C96 VTAIL.n54 VSUBS 0.023304f
C97 VTAIL.n55 VSUBS 0.012523f
C98 VTAIL.n56 VSUBS 0.013259f
C99 VTAIL.n57 VSUBS 0.029599f
C100 VTAIL.n58 VSUBS 0.029599f
C101 VTAIL.n59 VSUBS 0.013259f
C102 VTAIL.n60 VSUBS 0.012523f
C103 VTAIL.n61 VSUBS 0.023304f
C104 VTAIL.n62 VSUBS 0.023304f
C105 VTAIL.n63 VSUBS 0.012523f
C106 VTAIL.n64 VSUBS 0.013259f
C107 VTAIL.n65 VSUBS 0.029599f
C108 VTAIL.n66 VSUBS 0.029599f
C109 VTAIL.n67 VSUBS 0.013259f
C110 VTAIL.n68 VSUBS 0.012523f
C111 VTAIL.n69 VSUBS 0.023304f
C112 VTAIL.n70 VSUBS 0.023304f
C113 VTAIL.n71 VSUBS 0.012523f
C114 VTAIL.n72 VSUBS 0.012523f
C115 VTAIL.n73 VSUBS 0.013259f
C116 VTAIL.n74 VSUBS 0.029599f
C117 VTAIL.n75 VSUBS 0.029599f
C118 VTAIL.n76 VSUBS 0.029599f
C119 VTAIL.n77 VSUBS 0.012891f
C120 VTAIL.n78 VSUBS 0.012523f
C121 VTAIL.n79 VSUBS 0.023304f
C122 VTAIL.n80 VSUBS 0.023304f
C123 VTAIL.n81 VSUBS 0.012523f
C124 VTAIL.n82 VSUBS 0.013259f
C125 VTAIL.n83 VSUBS 0.029599f
C126 VTAIL.n84 VSUBS 0.029599f
C127 VTAIL.n85 VSUBS 0.013259f
C128 VTAIL.n86 VSUBS 0.012523f
C129 VTAIL.n87 VSUBS 0.023304f
C130 VTAIL.n88 VSUBS 0.023304f
C131 VTAIL.n89 VSUBS 0.012523f
C132 VTAIL.n90 VSUBS 0.013259f
C133 VTAIL.n91 VSUBS 0.029599f
C134 VTAIL.n92 VSUBS 0.072669f
C135 VTAIL.n93 VSUBS 0.013259f
C136 VTAIL.n94 VSUBS 0.012523f
C137 VTAIL.n95 VSUBS 0.056412f
C138 VTAIL.n96 VSUBS 0.036666f
C139 VTAIL.n97 VSUBS 0.080411f
C140 VTAIL.n98 VSUBS 0.025904f
C141 VTAIL.n99 VSUBS 0.023304f
C142 VTAIL.n100 VSUBS 0.012523f
C143 VTAIL.n101 VSUBS 0.029599f
C144 VTAIL.n102 VSUBS 0.013259f
C145 VTAIL.n103 VSUBS 0.023304f
C146 VTAIL.n104 VSUBS 0.012523f
C147 VTAIL.n105 VSUBS 0.029599f
C148 VTAIL.n106 VSUBS 0.012891f
C149 VTAIL.n107 VSUBS 0.023304f
C150 VTAIL.n108 VSUBS 0.013259f
C151 VTAIL.n109 VSUBS 0.029599f
C152 VTAIL.n110 VSUBS 0.013259f
C153 VTAIL.n111 VSUBS 0.023304f
C154 VTAIL.n112 VSUBS 0.012523f
C155 VTAIL.n113 VSUBS 0.029599f
C156 VTAIL.n114 VSUBS 0.013259f
C157 VTAIL.n115 VSUBS 0.023304f
C158 VTAIL.n116 VSUBS 0.012523f
C159 VTAIL.n117 VSUBS 0.029599f
C160 VTAIL.n118 VSUBS 0.013259f
C161 VTAIL.n119 VSUBS 0.023304f
C162 VTAIL.n120 VSUBS 0.012523f
C163 VTAIL.n121 VSUBS 0.029599f
C164 VTAIL.n122 VSUBS 0.013259f
C165 VTAIL.n123 VSUBS 0.023304f
C166 VTAIL.n124 VSUBS 0.012523f
C167 VTAIL.n125 VSUBS 0.029599f
C168 VTAIL.n126 VSUBS 0.013259f
C169 VTAIL.n127 VSUBS 1.76306f
C170 VTAIL.n128 VSUBS 0.012523f
C171 VTAIL.t2 VSUBS 0.063515f
C172 VTAIL.n129 VSUBS 0.182143f
C173 VTAIL.n130 VSUBS 0.018829f
C174 VTAIL.n131 VSUBS 0.022199f
C175 VTAIL.n132 VSUBS 0.029599f
C176 VTAIL.n133 VSUBS 0.013259f
C177 VTAIL.n134 VSUBS 0.012523f
C178 VTAIL.n135 VSUBS 0.023304f
C179 VTAIL.n136 VSUBS 0.023304f
C180 VTAIL.n137 VSUBS 0.012523f
C181 VTAIL.n138 VSUBS 0.013259f
C182 VTAIL.n139 VSUBS 0.029599f
C183 VTAIL.n140 VSUBS 0.029599f
C184 VTAIL.n141 VSUBS 0.013259f
C185 VTAIL.n142 VSUBS 0.012523f
C186 VTAIL.n143 VSUBS 0.023304f
C187 VTAIL.n144 VSUBS 0.023304f
C188 VTAIL.n145 VSUBS 0.012523f
C189 VTAIL.n146 VSUBS 0.013259f
C190 VTAIL.n147 VSUBS 0.029599f
C191 VTAIL.n148 VSUBS 0.029599f
C192 VTAIL.n149 VSUBS 0.013259f
C193 VTAIL.n150 VSUBS 0.012523f
C194 VTAIL.n151 VSUBS 0.023304f
C195 VTAIL.n152 VSUBS 0.023304f
C196 VTAIL.n153 VSUBS 0.012523f
C197 VTAIL.n154 VSUBS 0.013259f
C198 VTAIL.n155 VSUBS 0.029599f
C199 VTAIL.n156 VSUBS 0.029599f
C200 VTAIL.n157 VSUBS 0.013259f
C201 VTAIL.n158 VSUBS 0.012523f
C202 VTAIL.n159 VSUBS 0.023304f
C203 VTAIL.n160 VSUBS 0.023304f
C204 VTAIL.n161 VSUBS 0.012523f
C205 VTAIL.n162 VSUBS 0.013259f
C206 VTAIL.n163 VSUBS 0.029599f
C207 VTAIL.n164 VSUBS 0.029599f
C208 VTAIL.n165 VSUBS 0.013259f
C209 VTAIL.n166 VSUBS 0.012523f
C210 VTAIL.n167 VSUBS 0.023304f
C211 VTAIL.n168 VSUBS 0.023304f
C212 VTAIL.n169 VSUBS 0.012523f
C213 VTAIL.n170 VSUBS 0.012523f
C214 VTAIL.n171 VSUBS 0.013259f
C215 VTAIL.n172 VSUBS 0.029599f
C216 VTAIL.n173 VSUBS 0.029599f
C217 VTAIL.n174 VSUBS 0.029599f
C218 VTAIL.n175 VSUBS 0.012891f
C219 VTAIL.n176 VSUBS 0.012523f
C220 VTAIL.n177 VSUBS 0.023304f
C221 VTAIL.n178 VSUBS 0.023304f
C222 VTAIL.n179 VSUBS 0.012523f
C223 VTAIL.n180 VSUBS 0.013259f
C224 VTAIL.n181 VSUBS 0.029599f
C225 VTAIL.n182 VSUBS 0.029599f
C226 VTAIL.n183 VSUBS 0.013259f
C227 VTAIL.n184 VSUBS 0.012523f
C228 VTAIL.n185 VSUBS 0.023304f
C229 VTAIL.n186 VSUBS 0.023304f
C230 VTAIL.n187 VSUBS 0.012523f
C231 VTAIL.n188 VSUBS 0.013259f
C232 VTAIL.n189 VSUBS 0.029599f
C233 VTAIL.n190 VSUBS 0.072669f
C234 VTAIL.n191 VSUBS 0.013259f
C235 VTAIL.n192 VSUBS 0.012523f
C236 VTAIL.n193 VSUBS 0.056412f
C237 VTAIL.n194 VSUBS 0.036666f
C238 VTAIL.n195 VSUBS 0.095461f
C239 VTAIL.n196 VSUBS 0.025904f
C240 VTAIL.n197 VSUBS 0.023304f
C241 VTAIL.n198 VSUBS 0.012523f
C242 VTAIL.n199 VSUBS 0.029599f
C243 VTAIL.n200 VSUBS 0.013259f
C244 VTAIL.n201 VSUBS 0.023304f
C245 VTAIL.n202 VSUBS 0.012523f
C246 VTAIL.n203 VSUBS 0.029599f
C247 VTAIL.n204 VSUBS 0.012891f
C248 VTAIL.n205 VSUBS 0.023304f
C249 VTAIL.n206 VSUBS 0.013259f
C250 VTAIL.n207 VSUBS 0.029599f
C251 VTAIL.n208 VSUBS 0.013259f
C252 VTAIL.n209 VSUBS 0.023304f
C253 VTAIL.n210 VSUBS 0.012523f
C254 VTAIL.n211 VSUBS 0.029599f
C255 VTAIL.n212 VSUBS 0.013259f
C256 VTAIL.n213 VSUBS 0.023304f
C257 VTAIL.n214 VSUBS 0.012523f
C258 VTAIL.n215 VSUBS 0.029599f
C259 VTAIL.n216 VSUBS 0.013259f
C260 VTAIL.n217 VSUBS 0.023304f
C261 VTAIL.n218 VSUBS 0.012523f
C262 VTAIL.n219 VSUBS 0.029599f
C263 VTAIL.n220 VSUBS 0.013259f
C264 VTAIL.n221 VSUBS 0.023304f
C265 VTAIL.n222 VSUBS 0.012523f
C266 VTAIL.n223 VSUBS 0.029599f
C267 VTAIL.n224 VSUBS 0.013259f
C268 VTAIL.n225 VSUBS 1.76306f
C269 VTAIL.n226 VSUBS 0.012523f
C270 VTAIL.t0 VSUBS 0.063515f
C271 VTAIL.n227 VSUBS 0.182143f
C272 VTAIL.n228 VSUBS 0.018829f
C273 VTAIL.n229 VSUBS 0.022199f
C274 VTAIL.n230 VSUBS 0.029599f
C275 VTAIL.n231 VSUBS 0.013259f
C276 VTAIL.n232 VSUBS 0.012523f
C277 VTAIL.n233 VSUBS 0.023304f
C278 VTAIL.n234 VSUBS 0.023304f
C279 VTAIL.n235 VSUBS 0.012523f
C280 VTAIL.n236 VSUBS 0.013259f
C281 VTAIL.n237 VSUBS 0.029599f
C282 VTAIL.n238 VSUBS 0.029599f
C283 VTAIL.n239 VSUBS 0.013259f
C284 VTAIL.n240 VSUBS 0.012523f
C285 VTAIL.n241 VSUBS 0.023304f
C286 VTAIL.n242 VSUBS 0.023304f
C287 VTAIL.n243 VSUBS 0.012523f
C288 VTAIL.n244 VSUBS 0.013259f
C289 VTAIL.n245 VSUBS 0.029599f
C290 VTAIL.n246 VSUBS 0.029599f
C291 VTAIL.n247 VSUBS 0.013259f
C292 VTAIL.n248 VSUBS 0.012523f
C293 VTAIL.n249 VSUBS 0.023304f
C294 VTAIL.n250 VSUBS 0.023304f
C295 VTAIL.n251 VSUBS 0.012523f
C296 VTAIL.n252 VSUBS 0.013259f
C297 VTAIL.n253 VSUBS 0.029599f
C298 VTAIL.n254 VSUBS 0.029599f
C299 VTAIL.n255 VSUBS 0.013259f
C300 VTAIL.n256 VSUBS 0.012523f
C301 VTAIL.n257 VSUBS 0.023304f
C302 VTAIL.n258 VSUBS 0.023304f
C303 VTAIL.n259 VSUBS 0.012523f
C304 VTAIL.n260 VSUBS 0.013259f
C305 VTAIL.n261 VSUBS 0.029599f
C306 VTAIL.n262 VSUBS 0.029599f
C307 VTAIL.n263 VSUBS 0.013259f
C308 VTAIL.n264 VSUBS 0.012523f
C309 VTAIL.n265 VSUBS 0.023304f
C310 VTAIL.n266 VSUBS 0.023304f
C311 VTAIL.n267 VSUBS 0.012523f
C312 VTAIL.n268 VSUBS 0.012523f
C313 VTAIL.n269 VSUBS 0.013259f
C314 VTAIL.n270 VSUBS 0.029599f
C315 VTAIL.n271 VSUBS 0.029599f
C316 VTAIL.n272 VSUBS 0.029599f
C317 VTAIL.n273 VSUBS 0.012891f
C318 VTAIL.n274 VSUBS 0.012523f
C319 VTAIL.n275 VSUBS 0.023304f
C320 VTAIL.n276 VSUBS 0.023304f
C321 VTAIL.n277 VSUBS 0.012523f
C322 VTAIL.n278 VSUBS 0.013259f
C323 VTAIL.n279 VSUBS 0.029599f
C324 VTAIL.n280 VSUBS 0.029599f
C325 VTAIL.n281 VSUBS 0.013259f
C326 VTAIL.n282 VSUBS 0.012523f
C327 VTAIL.n283 VSUBS 0.023304f
C328 VTAIL.n284 VSUBS 0.023304f
C329 VTAIL.n285 VSUBS 0.012523f
C330 VTAIL.n286 VSUBS 0.013259f
C331 VTAIL.n287 VSUBS 0.029599f
C332 VTAIL.n288 VSUBS 0.072669f
C333 VTAIL.n289 VSUBS 0.013259f
C334 VTAIL.n290 VSUBS 0.012523f
C335 VTAIL.n291 VSUBS 0.056412f
C336 VTAIL.n292 VSUBS 0.036666f
C337 VTAIL.n293 VSUBS 1.55617f
C338 VTAIL.n294 VSUBS 0.025904f
C339 VTAIL.n295 VSUBS 0.023304f
C340 VTAIL.n296 VSUBS 0.012523f
C341 VTAIL.n297 VSUBS 0.029599f
C342 VTAIL.n298 VSUBS 0.013259f
C343 VTAIL.n299 VSUBS 0.023304f
C344 VTAIL.n300 VSUBS 0.012523f
C345 VTAIL.n301 VSUBS 0.029599f
C346 VTAIL.n302 VSUBS 0.012891f
C347 VTAIL.n303 VSUBS 0.023304f
C348 VTAIL.n304 VSUBS 0.012891f
C349 VTAIL.n305 VSUBS 0.012523f
C350 VTAIL.n306 VSUBS 0.029599f
C351 VTAIL.n307 VSUBS 0.029599f
C352 VTAIL.n308 VSUBS 0.013259f
C353 VTAIL.n309 VSUBS 0.023304f
C354 VTAIL.n310 VSUBS 0.012523f
C355 VTAIL.n311 VSUBS 0.029599f
C356 VTAIL.n312 VSUBS 0.013259f
C357 VTAIL.n313 VSUBS 0.023304f
C358 VTAIL.n314 VSUBS 0.012523f
C359 VTAIL.n315 VSUBS 0.029599f
C360 VTAIL.n316 VSUBS 0.013259f
C361 VTAIL.n317 VSUBS 0.023304f
C362 VTAIL.n318 VSUBS 0.012523f
C363 VTAIL.n319 VSUBS 0.029599f
C364 VTAIL.n320 VSUBS 0.013259f
C365 VTAIL.n321 VSUBS 0.023304f
C366 VTAIL.n322 VSUBS 0.012523f
C367 VTAIL.n323 VSUBS 0.029599f
C368 VTAIL.n324 VSUBS 0.013259f
C369 VTAIL.n325 VSUBS 1.76306f
C370 VTAIL.n326 VSUBS 0.012523f
C371 VTAIL.t6 VSUBS 0.063515f
C372 VTAIL.n327 VSUBS 0.182143f
C373 VTAIL.n328 VSUBS 0.018829f
C374 VTAIL.n329 VSUBS 0.022199f
C375 VTAIL.n330 VSUBS 0.029599f
C376 VTAIL.n331 VSUBS 0.013259f
C377 VTAIL.n332 VSUBS 0.012523f
C378 VTAIL.n333 VSUBS 0.023304f
C379 VTAIL.n334 VSUBS 0.023304f
C380 VTAIL.n335 VSUBS 0.012523f
C381 VTAIL.n336 VSUBS 0.013259f
C382 VTAIL.n337 VSUBS 0.029599f
C383 VTAIL.n338 VSUBS 0.029599f
C384 VTAIL.n339 VSUBS 0.013259f
C385 VTAIL.n340 VSUBS 0.012523f
C386 VTAIL.n341 VSUBS 0.023304f
C387 VTAIL.n342 VSUBS 0.023304f
C388 VTAIL.n343 VSUBS 0.012523f
C389 VTAIL.n344 VSUBS 0.013259f
C390 VTAIL.n345 VSUBS 0.029599f
C391 VTAIL.n346 VSUBS 0.029599f
C392 VTAIL.n347 VSUBS 0.013259f
C393 VTAIL.n348 VSUBS 0.012523f
C394 VTAIL.n349 VSUBS 0.023304f
C395 VTAIL.n350 VSUBS 0.023304f
C396 VTAIL.n351 VSUBS 0.012523f
C397 VTAIL.n352 VSUBS 0.013259f
C398 VTAIL.n353 VSUBS 0.029599f
C399 VTAIL.n354 VSUBS 0.029599f
C400 VTAIL.n355 VSUBS 0.013259f
C401 VTAIL.n356 VSUBS 0.012523f
C402 VTAIL.n357 VSUBS 0.023304f
C403 VTAIL.n358 VSUBS 0.023304f
C404 VTAIL.n359 VSUBS 0.012523f
C405 VTAIL.n360 VSUBS 0.013259f
C406 VTAIL.n361 VSUBS 0.029599f
C407 VTAIL.n362 VSUBS 0.029599f
C408 VTAIL.n363 VSUBS 0.013259f
C409 VTAIL.n364 VSUBS 0.012523f
C410 VTAIL.n365 VSUBS 0.023304f
C411 VTAIL.n366 VSUBS 0.023304f
C412 VTAIL.n367 VSUBS 0.012523f
C413 VTAIL.n368 VSUBS 0.013259f
C414 VTAIL.n369 VSUBS 0.029599f
C415 VTAIL.n370 VSUBS 0.029599f
C416 VTAIL.n371 VSUBS 0.013259f
C417 VTAIL.n372 VSUBS 0.012523f
C418 VTAIL.n373 VSUBS 0.023304f
C419 VTAIL.n374 VSUBS 0.023304f
C420 VTAIL.n375 VSUBS 0.012523f
C421 VTAIL.n376 VSUBS 0.013259f
C422 VTAIL.n377 VSUBS 0.029599f
C423 VTAIL.n378 VSUBS 0.029599f
C424 VTAIL.n379 VSUBS 0.013259f
C425 VTAIL.n380 VSUBS 0.012523f
C426 VTAIL.n381 VSUBS 0.023304f
C427 VTAIL.n382 VSUBS 0.023304f
C428 VTAIL.n383 VSUBS 0.012523f
C429 VTAIL.n384 VSUBS 0.013259f
C430 VTAIL.n385 VSUBS 0.029599f
C431 VTAIL.n386 VSUBS 0.072669f
C432 VTAIL.n387 VSUBS 0.013259f
C433 VTAIL.n388 VSUBS 0.012523f
C434 VTAIL.n389 VSUBS 0.056412f
C435 VTAIL.n390 VSUBS 0.036666f
C436 VTAIL.n391 VSUBS 1.55617f
C437 VTAIL.n392 VSUBS 0.025904f
C438 VTAIL.n393 VSUBS 0.023304f
C439 VTAIL.n394 VSUBS 0.012523f
C440 VTAIL.n395 VSUBS 0.029599f
C441 VTAIL.n396 VSUBS 0.013259f
C442 VTAIL.n397 VSUBS 0.023304f
C443 VTAIL.n398 VSUBS 0.012523f
C444 VTAIL.n399 VSUBS 0.029599f
C445 VTAIL.n400 VSUBS 0.012891f
C446 VTAIL.n401 VSUBS 0.023304f
C447 VTAIL.n402 VSUBS 0.012891f
C448 VTAIL.n403 VSUBS 0.012523f
C449 VTAIL.n404 VSUBS 0.029599f
C450 VTAIL.n405 VSUBS 0.029599f
C451 VTAIL.n406 VSUBS 0.013259f
C452 VTAIL.n407 VSUBS 0.023304f
C453 VTAIL.n408 VSUBS 0.012523f
C454 VTAIL.n409 VSUBS 0.029599f
C455 VTAIL.n410 VSUBS 0.013259f
C456 VTAIL.n411 VSUBS 0.023304f
C457 VTAIL.n412 VSUBS 0.012523f
C458 VTAIL.n413 VSUBS 0.029599f
C459 VTAIL.n414 VSUBS 0.013259f
C460 VTAIL.n415 VSUBS 0.023304f
C461 VTAIL.n416 VSUBS 0.012523f
C462 VTAIL.n417 VSUBS 0.029599f
C463 VTAIL.n418 VSUBS 0.013259f
C464 VTAIL.n419 VSUBS 0.023304f
C465 VTAIL.n420 VSUBS 0.012523f
C466 VTAIL.n421 VSUBS 0.029599f
C467 VTAIL.n422 VSUBS 0.013259f
C468 VTAIL.n423 VSUBS 1.76306f
C469 VTAIL.n424 VSUBS 0.012523f
C470 VTAIL.t4 VSUBS 0.063515f
C471 VTAIL.n425 VSUBS 0.182143f
C472 VTAIL.n426 VSUBS 0.018829f
C473 VTAIL.n427 VSUBS 0.022199f
C474 VTAIL.n428 VSUBS 0.029599f
C475 VTAIL.n429 VSUBS 0.013259f
C476 VTAIL.n430 VSUBS 0.012523f
C477 VTAIL.n431 VSUBS 0.023304f
C478 VTAIL.n432 VSUBS 0.023304f
C479 VTAIL.n433 VSUBS 0.012523f
C480 VTAIL.n434 VSUBS 0.013259f
C481 VTAIL.n435 VSUBS 0.029599f
C482 VTAIL.n436 VSUBS 0.029599f
C483 VTAIL.n437 VSUBS 0.013259f
C484 VTAIL.n438 VSUBS 0.012523f
C485 VTAIL.n439 VSUBS 0.023304f
C486 VTAIL.n440 VSUBS 0.023304f
C487 VTAIL.n441 VSUBS 0.012523f
C488 VTAIL.n442 VSUBS 0.013259f
C489 VTAIL.n443 VSUBS 0.029599f
C490 VTAIL.n444 VSUBS 0.029599f
C491 VTAIL.n445 VSUBS 0.013259f
C492 VTAIL.n446 VSUBS 0.012523f
C493 VTAIL.n447 VSUBS 0.023304f
C494 VTAIL.n448 VSUBS 0.023304f
C495 VTAIL.n449 VSUBS 0.012523f
C496 VTAIL.n450 VSUBS 0.013259f
C497 VTAIL.n451 VSUBS 0.029599f
C498 VTAIL.n452 VSUBS 0.029599f
C499 VTAIL.n453 VSUBS 0.013259f
C500 VTAIL.n454 VSUBS 0.012523f
C501 VTAIL.n455 VSUBS 0.023304f
C502 VTAIL.n456 VSUBS 0.023304f
C503 VTAIL.n457 VSUBS 0.012523f
C504 VTAIL.n458 VSUBS 0.013259f
C505 VTAIL.n459 VSUBS 0.029599f
C506 VTAIL.n460 VSUBS 0.029599f
C507 VTAIL.n461 VSUBS 0.013259f
C508 VTAIL.n462 VSUBS 0.012523f
C509 VTAIL.n463 VSUBS 0.023304f
C510 VTAIL.n464 VSUBS 0.023304f
C511 VTAIL.n465 VSUBS 0.012523f
C512 VTAIL.n466 VSUBS 0.013259f
C513 VTAIL.n467 VSUBS 0.029599f
C514 VTAIL.n468 VSUBS 0.029599f
C515 VTAIL.n469 VSUBS 0.013259f
C516 VTAIL.n470 VSUBS 0.012523f
C517 VTAIL.n471 VSUBS 0.023304f
C518 VTAIL.n472 VSUBS 0.023304f
C519 VTAIL.n473 VSUBS 0.012523f
C520 VTAIL.n474 VSUBS 0.013259f
C521 VTAIL.n475 VSUBS 0.029599f
C522 VTAIL.n476 VSUBS 0.029599f
C523 VTAIL.n477 VSUBS 0.013259f
C524 VTAIL.n478 VSUBS 0.012523f
C525 VTAIL.n479 VSUBS 0.023304f
C526 VTAIL.n480 VSUBS 0.023304f
C527 VTAIL.n481 VSUBS 0.012523f
C528 VTAIL.n482 VSUBS 0.013259f
C529 VTAIL.n483 VSUBS 0.029599f
C530 VTAIL.n484 VSUBS 0.072669f
C531 VTAIL.n485 VSUBS 0.013259f
C532 VTAIL.n486 VSUBS 0.012523f
C533 VTAIL.n487 VSUBS 0.056412f
C534 VTAIL.n488 VSUBS 0.036666f
C535 VTAIL.n489 VSUBS 0.095461f
C536 VTAIL.n490 VSUBS 0.025904f
C537 VTAIL.n491 VSUBS 0.023304f
C538 VTAIL.n492 VSUBS 0.012523f
C539 VTAIL.n493 VSUBS 0.029599f
C540 VTAIL.n494 VSUBS 0.013259f
C541 VTAIL.n495 VSUBS 0.023304f
C542 VTAIL.n496 VSUBS 0.012523f
C543 VTAIL.n497 VSUBS 0.029599f
C544 VTAIL.n498 VSUBS 0.012891f
C545 VTAIL.n499 VSUBS 0.023304f
C546 VTAIL.n500 VSUBS 0.012891f
C547 VTAIL.n501 VSUBS 0.012523f
C548 VTAIL.n502 VSUBS 0.029599f
C549 VTAIL.n503 VSUBS 0.029599f
C550 VTAIL.n504 VSUBS 0.013259f
C551 VTAIL.n505 VSUBS 0.023304f
C552 VTAIL.n506 VSUBS 0.012523f
C553 VTAIL.n507 VSUBS 0.029599f
C554 VTAIL.n508 VSUBS 0.013259f
C555 VTAIL.n509 VSUBS 0.023304f
C556 VTAIL.n510 VSUBS 0.012523f
C557 VTAIL.n511 VSUBS 0.029599f
C558 VTAIL.n512 VSUBS 0.013259f
C559 VTAIL.n513 VSUBS 0.023304f
C560 VTAIL.n514 VSUBS 0.012523f
C561 VTAIL.n515 VSUBS 0.029599f
C562 VTAIL.n516 VSUBS 0.013259f
C563 VTAIL.n517 VSUBS 0.023304f
C564 VTAIL.n518 VSUBS 0.012523f
C565 VTAIL.n519 VSUBS 0.029599f
C566 VTAIL.n520 VSUBS 0.013259f
C567 VTAIL.n521 VSUBS 1.76306f
C568 VTAIL.n522 VSUBS 0.012523f
C569 VTAIL.t3 VSUBS 0.063515f
C570 VTAIL.n523 VSUBS 0.182143f
C571 VTAIL.n524 VSUBS 0.018829f
C572 VTAIL.n525 VSUBS 0.022199f
C573 VTAIL.n526 VSUBS 0.029599f
C574 VTAIL.n527 VSUBS 0.013259f
C575 VTAIL.n528 VSUBS 0.012523f
C576 VTAIL.n529 VSUBS 0.023304f
C577 VTAIL.n530 VSUBS 0.023304f
C578 VTAIL.n531 VSUBS 0.012523f
C579 VTAIL.n532 VSUBS 0.013259f
C580 VTAIL.n533 VSUBS 0.029599f
C581 VTAIL.n534 VSUBS 0.029599f
C582 VTAIL.n535 VSUBS 0.013259f
C583 VTAIL.n536 VSUBS 0.012523f
C584 VTAIL.n537 VSUBS 0.023304f
C585 VTAIL.n538 VSUBS 0.023304f
C586 VTAIL.n539 VSUBS 0.012523f
C587 VTAIL.n540 VSUBS 0.013259f
C588 VTAIL.n541 VSUBS 0.029599f
C589 VTAIL.n542 VSUBS 0.029599f
C590 VTAIL.n543 VSUBS 0.013259f
C591 VTAIL.n544 VSUBS 0.012523f
C592 VTAIL.n545 VSUBS 0.023304f
C593 VTAIL.n546 VSUBS 0.023304f
C594 VTAIL.n547 VSUBS 0.012523f
C595 VTAIL.n548 VSUBS 0.013259f
C596 VTAIL.n549 VSUBS 0.029599f
C597 VTAIL.n550 VSUBS 0.029599f
C598 VTAIL.n551 VSUBS 0.013259f
C599 VTAIL.n552 VSUBS 0.012523f
C600 VTAIL.n553 VSUBS 0.023304f
C601 VTAIL.n554 VSUBS 0.023304f
C602 VTAIL.n555 VSUBS 0.012523f
C603 VTAIL.n556 VSUBS 0.013259f
C604 VTAIL.n557 VSUBS 0.029599f
C605 VTAIL.n558 VSUBS 0.029599f
C606 VTAIL.n559 VSUBS 0.013259f
C607 VTAIL.n560 VSUBS 0.012523f
C608 VTAIL.n561 VSUBS 0.023304f
C609 VTAIL.n562 VSUBS 0.023304f
C610 VTAIL.n563 VSUBS 0.012523f
C611 VTAIL.n564 VSUBS 0.013259f
C612 VTAIL.n565 VSUBS 0.029599f
C613 VTAIL.n566 VSUBS 0.029599f
C614 VTAIL.n567 VSUBS 0.013259f
C615 VTAIL.n568 VSUBS 0.012523f
C616 VTAIL.n569 VSUBS 0.023304f
C617 VTAIL.n570 VSUBS 0.023304f
C618 VTAIL.n571 VSUBS 0.012523f
C619 VTAIL.n572 VSUBS 0.013259f
C620 VTAIL.n573 VSUBS 0.029599f
C621 VTAIL.n574 VSUBS 0.029599f
C622 VTAIL.n575 VSUBS 0.013259f
C623 VTAIL.n576 VSUBS 0.012523f
C624 VTAIL.n577 VSUBS 0.023304f
C625 VTAIL.n578 VSUBS 0.023304f
C626 VTAIL.n579 VSUBS 0.012523f
C627 VTAIL.n580 VSUBS 0.013259f
C628 VTAIL.n581 VSUBS 0.029599f
C629 VTAIL.n582 VSUBS 0.072669f
C630 VTAIL.n583 VSUBS 0.013259f
C631 VTAIL.n584 VSUBS 0.012523f
C632 VTAIL.n585 VSUBS 0.056412f
C633 VTAIL.n586 VSUBS 0.036666f
C634 VTAIL.n587 VSUBS 0.095461f
C635 VTAIL.n588 VSUBS 0.025904f
C636 VTAIL.n589 VSUBS 0.023304f
C637 VTAIL.n590 VSUBS 0.012523f
C638 VTAIL.n591 VSUBS 0.029599f
C639 VTAIL.n592 VSUBS 0.013259f
C640 VTAIL.n593 VSUBS 0.023304f
C641 VTAIL.n594 VSUBS 0.012523f
C642 VTAIL.n595 VSUBS 0.029599f
C643 VTAIL.n596 VSUBS 0.012891f
C644 VTAIL.n597 VSUBS 0.023304f
C645 VTAIL.n598 VSUBS 0.012891f
C646 VTAIL.n599 VSUBS 0.012523f
C647 VTAIL.n600 VSUBS 0.029599f
C648 VTAIL.n601 VSUBS 0.029599f
C649 VTAIL.n602 VSUBS 0.013259f
C650 VTAIL.n603 VSUBS 0.023304f
C651 VTAIL.n604 VSUBS 0.012523f
C652 VTAIL.n605 VSUBS 0.029599f
C653 VTAIL.n606 VSUBS 0.013259f
C654 VTAIL.n607 VSUBS 0.023304f
C655 VTAIL.n608 VSUBS 0.012523f
C656 VTAIL.n609 VSUBS 0.029599f
C657 VTAIL.n610 VSUBS 0.013259f
C658 VTAIL.n611 VSUBS 0.023304f
C659 VTAIL.n612 VSUBS 0.012523f
C660 VTAIL.n613 VSUBS 0.029599f
C661 VTAIL.n614 VSUBS 0.013259f
C662 VTAIL.n615 VSUBS 0.023304f
C663 VTAIL.n616 VSUBS 0.012523f
C664 VTAIL.n617 VSUBS 0.029599f
C665 VTAIL.n618 VSUBS 0.013259f
C666 VTAIL.n619 VSUBS 1.76306f
C667 VTAIL.n620 VSUBS 0.012523f
C668 VTAIL.t1 VSUBS 0.063515f
C669 VTAIL.n621 VSUBS 0.182143f
C670 VTAIL.n622 VSUBS 0.018829f
C671 VTAIL.n623 VSUBS 0.022199f
C672 VTAIL.n624 VSUBS 0.029599f
C673 VTAIL.n625 VSUBS 0.013259f
C674 VTAIL.n626 VSUBS 0.012523f
C675 VTAIL.n627 VSUBS 0.023304f
C676 VTAIL.n628 VSUBS 0.023304f
C677 VTAIL.n629 VSUBS 0.012523f
C678 VTAIL.n630 VSUBS 0.013259f
C679 VTAIL.n631 VSUBS 0.029599f
C680 VTAIL.n632 VSUBS 0.029599f
C681 VTAIL.n633 VSUBS 0.013259f
C682 VTAIL.n634 VSUBS 0.012523f
C683 VTAIL.n635 VSUBS 0.023304f
C684 VTAIL.n636 VSUBS 0.023304f
C685 VTAIL.n637 VSUBS 0.012523f
C686 VTAIL.n638 VSUBS 0.013259f
C687 VTAIL.n639 VSUBS 0.029599f
C688 VTAIL.n640 VSUBS 0.029599f
C689 VTAIL.n641 VSUBS 0.013259f
C690 VTAIL.n642 VSUBS 0.012523f
C691 VTAIL.n643 VSUBS 0.023304f
C692 VTAIL.n644 VSUBS 0.023304f
C693 VTAIL.n645 VSUBS 0.012523f
C694 VTAIL.n646 VSUBS 0.013259f
C695 VTAIL.n647 VSUBS 0.029599f
C696 VTAIL.n648 VSUBS 0.029599f
C697 VTAIL.n649 VSUBS 0.013259f
C698 VTAIL.n650 VSUBS 0.012523f
C699 VTAIL.n651 VSUBS 0.023304f
C700 VTAIL.n652 VSUBS 0.023304f
C701 VTAIL.n653 VSUBS 0.012523f
C702 VTAIL.n654 VSUBS 0.013259f
C703 VTAIL.n655 VSUBS 0.029599f
C704 VTAIL.n656 VSUBS 0.029599f
C705 VTAIL.n657 VSUBS 0.013259f
C706 VTAIL.n658 VSUBS 0.012523f
C707 VTAIL.n659 VSUBS 0.023304f
C708 VTAIL.n660 VSUBS 0.023304f
C709 VTAIL.n661 VSUBS 0.012523f
C710 VTAIL.n662 VSUBS 0.013259f
C711 VTAIL.n663 VSUBS 0.029599f
C712 VTAIL.n664 VSUBS 0.029599f
C713 VTAIL.n665 VSUBS 0.013259f
C714 VTAIL.n666 VSUBS 0.012523f
C715 VTAIL.n667 VSUBS 0.023304f
C716 VTAIL.n668 VSUBS 0.023304f
C717 VTAIL.n669 VSUBS 0.012523f
C718 VTAIL.n670 VSUBS 0.013259f
C719 VTAIL.n671 VSUBS 0.029599f
C720 VTAIL.n672 VSUBS 0.029599f
C721 VTAIL.n673 VSUBS 0.013259f
C722 VTAIL.n674 VSUBS 0.012523f
C723 VTAIL.n675 VSUBS 0.023304f
C724 VTAIL.n676 VSUBS 0.023304f
C725 VTAIL.n677 VSUBS 0.012523f
C726 VTAIL.n678 VSUBS 0.013259f
C727 VTAIL.n679 VSUBS 0.029599f
C728 VTAIL.n680 VSUBS 0.072669f
C729 VTAIL.n681 VSUBS 0.013259f
C730 VTAIL.n682 VSUBS 0.012523f
C731 VTAIL.n683 VSUBS 0.056412f
C732 VTAIL.n684 VSUBS 0.036666f
C733 VTAIL.n685 VSUBS 1.55617f
C734 VTAIL.n686 VSUBS 0.025904f
C735 VTAIL.n687 VSUBS 0.023304f
C736 VTAIL.n688 VSUBS 0.012523f
C737 VTAIL.n689 VSUBS 0.029599f
C738 VTAIL.n690 VSUBS 0.013259f
C739 VTAIL.n691 VSUBS 0.023304f
C740 VTAIL.n692 VSUBS 0.012523f
C741 VTAIL.n693 VSUBS 0.029599f
C742 VTAIL.n694 VSUBS 0.012891f
C743 VTAIL.n695 VSUBS 0.023304f
C744 VTAIL.n696 VSUBS 0.013259f
C745 VTAIL.n697 VSUBS 0.029599f
C746 VTAIL.n698 VSUBS 0.013259f
C747 VTAIL.n699 VSUBS 0.023304f
C748 VTAIL.n700 VSUBS 0.012523f
C749 VTAIL.n701 VSUBS 0.029599f
C750 VTAIL.n702 VSUBS 0.013259f
C751 VTAIL.n703 VSUBS 0.023304f
C752 VTAIL.n704 VSUBS 0.012523f
C753 VTAIL.n705 VSUBS 0.029599f
C754 VTAIL.n706 VSUBS 0.013259f
C755 VTAIL.n707 VSUBS 0.023304f
C756 VTAIL.n708 VSUBS 0.012523f
C757 VTAIL.n709 VSUBS 0.029599f
C758 VTAIL.n710 VSUBS 0.013259f
C759 VTAIL.n711 VSUBS 0.023304f
C760 VTAIL.n712 VSUBS 0.012523f
C761 VTAIL.n713 VSUBS 0.029599f
C762 VTAIL.n714 VSUBS 0.013259f
C763 VTAIL.n715 VSUBS 1.76306f
C764 VTAIL.n716 VSUBS 0.012523f
C765 VTAIL.t5 VSUBS 0.063515f
C766 VTAIL.n717 VSUBS 0.182143f
C767 VTAIL.n718 VSUBS 0.018829f
C768 VTAIL.n719 VSUBS 0.022199f
C769 VTAIL.n720 VSUBS 0.029599f
C770 VTAIL.n721 VSUBS 0.013259f
C771 VTAIL.n722 VSUBS 0.012523f
C772 VTAIL.n723 VSUBS 0.023304f
C773 VTAIL.n724 VSUBS 0.023304f
C774 VTAIL.n725 VSUBS 0.012523f
C775 VTAIL.n726 VSUBS 0.013259f
C776 VTAIL.n727 VSUBS 0.029599f
C777 VTAIL.n728 VSUBS 0.029599f
C778 VTAIL.n729 VSUBS 0.013259f
C779 VTAIL.n730 VSUBS 0.012523f
C780 VTAIL.n731 VSUBS 0.023304f
C781 VTAIL.n732 VSUBS 0.023304f
C782 VTAIL.n733 VSUBS 0.012523f
C783 VTAIL.n734 VSUBS 0.013259f
C784 VTAIL.n735 VSUBS 0.029599f
C785 VTAIL.n736 VSUBS 0.029599f
C786 VTAIL.n737 VSUBS 0.013259f
C787 VTAIL.n738 VSUBS 0.012523f
C788 VTAIL.n739 VSUBS 0.023304f
C789 VTAIL.n740 VSUBS 0.023304f
C790 VTAIL.n741 VSUBS 0.012523f
C791 VTAIL.n742 VSUBS 0.013259f
C792 VTAIL.n743 VSUBS 0.029599f
C793 VTAIL.n744 VSUBS 0.029599f
C794 VTAIL.n745 VSUBS 0.013259f
C795 VTAIL.n746 VSUBS 0.012523f
C796 VTAIL.n747 VSUBS 0.023304f
C797 VTAIL.n748 VSUBS 0.023304f
C798 VTAIL.n749 VSUBS 0.012523f
C799 VTAIL.n750 VSUBS 0.013259f
C800 VTAIL.n751 VSUBS 0.029599f
C801 VTAIL.n752 VSUBS 0.029599f
C802 VTAIL.n753 VSUBS 0.013259f
C803 VTAIL.n754 VSUBS 0.012523f
C804 VTAIL.n755 VSUBS 0.023304f
C805 VTAIL.n756 VSUBS 0.023304f
C806 VTAIL.n757 VSUBS 0.012523f
C807 VTAIL.n758 VSUBS 0.012523f
C808 VTAIL.n759 VSUBS 0.013259f
C809 VTAIL.n760 VSUBS 0.029599f
C810 VTAIL.n761 VSUBS 0.029599f
C811 VTAIL.n762 VSUBS 0.029599f
C812 VTAIL.n763 VSUBS 0.012891f
C813 VTAIL.n764 VSUBS 0.012523f
C814 VTAIL.n765 VSUBS 0.023304f
C815 VTAIL.n766 VSUBS 0.023304f
C816 VTAIL.n767 VSUBS 0.012523f
C817 VTAIL.n768 VSUBS 0.013259f
C818 VTAIL.n769 VSUBS 0.029599f
C819 VTAIL.n770 VSUBS 0.029599f
C820 VTAIL.n771 VSUBS 0.013259f
C821 VTAIL.n772 VSUBS 0.012523f
C822 VTAIL.n773 VSUBS 0.023304f
C823 VTAIL.n774 VSUBS 0.023304f
C824 VTAIL.n775 VSUBS 0.012523f
C825 VTAIL.n776 VSUBS 0.013259f
C826 VTAIL.n777 VSUBS 0.029599f
C827 VTAIL.n778 VSUBS 0.072669f
C828 VTAIL.n779 VSUBS 0.013259f
C829 VTAIL.n780 VSUBS 0.012523f
C830 VTAIL.n781 VSUBS 0.056412f
C831 VTAIL.n782 VSUBS 0.036666f
C832 VTAIL.n783 VSUBS 1.53238f
C833 VDD2.t2 VSUBS 0.482602f
C834 VDD2.t0 VSUBS 0.482602f
C835 VDD2.n0 VSUBS 5.04031f
C836 VDD2.t1 VSUBS 0.482602f
C837 VDD2.t3 VSUBS 0.482602f
C838 VDD2.n1 VSUBS 4.00663f
C839 VDD2.n2 VSUBS 5.65734f
C840 VN.t0 VSUBS 0.68148f
C841 VN.t2 VSUBS 0.68148f
C842 VN.n0 VSUBS 0.522988f
C843 VN.t1 VSUBS 0.68148f
C844 VN.t3 VSUBS 0.68148f
C845 VN.n1 VSUBS 1.00145f
C846 B.n0 VSUBS 0.007434f
C847 B.n1 VSUBS 0.007434f
C848 B.n2 VSUBS 0.010995f
C849 B.n3 VSUBS 0.008426f
C850 B.n4 VSUBS 0.008426f
C851 B.n5 VSUBS 0.008426f
C852 B.n6 VSUBS 0.008426f
C853 B.n7 VSUBS 0.008426f
C854 B.n8 VSUBS 0.018481f
C855 B.n9 VSUBS 0.008426f
C856 B.n10 VSUBS 0.008426f
C857 B.n11 VSUBS 0.008426f
C858 B.n12 VSUBS 0.008426f
C859 B.n13 VSUBS 0.008426f
C860 B.n14 VSUBS 0.008426f
C861 B.n15 VSUBS 0.008426f
C862 B.n16 VSUBS 0.008426f
C863 B.n17 VSUBS 0.008426f
C864 B.n18 VSUBS 0.008426f
C865 B.n19 VSUBS 0.008426f
C866 B.n20 VSUBS 0.008426f
C867 B.n21 VSUBS 0.008426f
C868 B.n22 VSUBS 0.008426f
C869 B.n23 VSUBS 0.008426f
C870 B.n24 VSUBS 0.008426f
C871 B.n25 VSUBS 0.008426f
C872 B.n26 VSUBS 0.008426f
C873 B.n27 VSUBS 0.008426f
C874 B.n28 VSUBS 0.008426f
C875 B.n29 VSUBS 0.008426f
C876 B.n30 VSUBS 0.008426f
C877 B.n31 VSUBS 0.008426f
C878 B.n32 VSUBS 0.008426f
C879 B.n33 VSUBS 0.008426f
C880 B.n34 VSUBS 0.008426f
C881 B.n35 VSUBS 0.008426f
C882 B.n36 VSUBS 0.008426f
C883 B.n37 VSUBS 0.008426f
C884 B.t10 VSUBS 0.411113f
C885 B.t11 VSUBS 0.419838f
C886 B.t9 VSUBS 0.221218f
C887 B.n38 VSUBS 0.43594f
C888 B.n39 VSUBS 0.378109f
C889 B.n40 VSUBS 0.008426f
C890 B.n41 VSUBS 0.008426f
C891 B.n42 VSUBS 0.008426f
C892 B.n43 VSUBS 0.008426f
C893 B.n44 VSUBS 0.004956f
C894 B.n45 VSUBS 0.008426f
C895 B.t4 VSUBS 0.411117f
C896 B.t5 VSUBS 0.419842f
C897 B.t3 VSUBS 0.221218f
C898 B.n46 VSUBS 0.435936f
C899 B.n47 VSUBS 0.378104f
C900 B.n48 VSUBS 0.019522f
C901 B.n49 VSUBS 0.008426f
C902 B.n50 VSUBS 0.008426f
C903 B.n51 VSUBS 0.008426f
C904 B.n52 VSUBS 0.008426f
C905 B.n53 VSUBS 0.008426f
C906 B.n54 VSUBS 0.008426f
C907 B.n55 VSUBS 0.008426f
C908 B.n56 VSUBS 0.008426f
C909 B.n57 VSUBS 0.008426f
C910 B.n58 VSUBS 0.008426f
C911 B.n59 VSUBS 0.008426f
C912 B.n60 VSUBS 0.008426f
C913 B.n61 VSUBS 0.008426f
C914 B.n62 VSUBS 0.008426f
C915 B.n63 VSUBS 0.008426f
C916 B.n64 VSUBS 0.008426f
C917 B.n65 VSUBS 0.008426f
C918 B.n66 VSUBS 0.008426f
C919 B.n67 VSUBS 0.008426f
C920 B.n68 VSUBS 0.008426f
C921 B.n69 VSUBS 0.008426f
C922 B.n70 VSUBS 0.008426f
C923 B.n71 VSUBS 0.008426f
C924 B.n72 VSUBS 0.008426f
C925 B.n73 VSUBS 0.008426f
C926 B.n74 VSUBS 0.008426f
C927 B.n75 VSUBS 0.008426f
C928 B.n76 VSUBS 0.019435f
C929 B.n77 VSUBS 0.008426f
C930 B.n78 VSUBS 0.008426f
C931 B.n79 VSUBS 0.008426f
C932 B.n80 VSUBS 0.008426f
C933 B.n81 VSUBS 0.008426f
C934 B.n82 VSUBS 0.008426f
C935 B.n83 VSUBS 0.008426f
C936 B.n84 VSUBS 0.008426f
C937 B.n85 VSUBS 0.008426f
C938 B.n86 VSUBS 0.008426f
C939 B.n87 VSUBS 0.008426f
C940 B.n88 VSUBS 0.008426f
C941 B.n89 VSUBS 0.008426f
C942 B.n90 VSUBS 0.018481f
C943 B.n91 VSUBS 0.008426f
C944 B.n92 VSUBS 0.008426f
C945 B.n93 VSUBS 0.008426f
C946 B.n94 VSUBS 0.008426f
C947 B.n95 VSUBS 0.008426f
C948 B.n96 VSUBS 0.008426f
C949 B.n97 VSUBS 0.008426f
C950 B.n98 VSUBS 0.008426f
C951 B.n99 VSUBS 0.008426f
C952 B.n100 VSUBS 0.008426f
C953 B.n101 VSUBS 0.008426f
C954 B.n102 VSUBS 0.008426f
C955 B.n103 VSUBS 0.008426f
C956 B.n104 VSUBS 0.008426f
C957 B.n105 VSUBS 0.008426f
C958 B.n106 VSUBS 0.008426f
C959 B.n107 VSUBS 0.008426f
C960 B.n108 VSUBS 0.008426f
C961 B.n109 VSUBS 0.008426f
C962 B.n110 VSUBS 0.008426f
C963 B.n111 VSUBS 0.008426f
C964 B.n112 VSUBS 0.008426f
C965 B.n113 VSUBS 0.008426f
C966 B.n114 VSUBS 0.008426f
C967 B.n115 VSUBS 0.008426f
C968 B.n116 VSUBS 0.008426f
C969 B.n117 VSUBS 0.008426f
C970 B.n118 VSUBS 0.008426f
C971 B.n119 VSUBS 0.007682f
C972 B.n120 VSUBS 0.008426f
C973 B.n121 VSUBS 0.008426f
C974 B.n122 VSUBS 0.008426f
C975 B.n123 VSUBS 0.008426f
C976 B.n124 VSUBS 0.008426f
C977 B.t2 VSUBS 0.411113f
C978 B.t1 VSUBS 0.419838f
C979 B.t0 VSUBS 0.221218f
C980 B.n125 VSUBS 0.43594f
C981 B.n126 VSUBS 0.378109f
C982 B.n127 VSUBS 0.008426f
C983 B.n128 VSUBS 0.008426f
C984 B.n129 VSUBS 0.008426f
C985 B.n130 VSUBS 0.008426f
C986 B.n131 VSUBS 0.008426f
C987 B.n132 VSUBS 0.008426f
C988 B.n133 VSUBS 0.008426f
C989 B.n134 VSUBS 0.008426f
C990 B.n135 VSUBS 0.008426f
C991 B.n136 VSUBS 0.008426f
C992 B.n137 VSUBS 0.008426f
C993 B.n138 VSUBS 0.008426f
C994 B.n139 VSUBS 0.008426f
C995 B.n140 VSUBS 0.008426f
C996 B.n141 VSUBS 0.008426f
C997 B.n142 VSUBS 0.008426f
C998 B.n143 VSUBS 0.008426f
C999 B.n144 VSUBS 0.008426f
C1000 B.n145 VSUBS 0.008426f
C1001 B.n146 VSUBS 0.008426f
C1002 B.n147 VSUBS 0.008426f
C1003 B.n148 VSUBS 0.008426f
C1004 B.n149 VSUBS 0.008426f
C1005 B.n150 VSUBS 0.008426f
C1006 B.n151 VSUBS 0.008426f
C1007 B.n152 VSUBS 0.008426f
C1008 B.n153 VSUBS 0.008426f
C1009 B.n154 VSUBS 0.008426f
C1010 B.n155 VSUBS 0.019435f
C1011 B.n156 VSUBS 0.008426f
C1012 B.n157 VSUBS 0.008426f
C1013 B.n158 VSUBS 0.008426f
C1014 B.n159 VSUBS 0.008426f
C1015 B.n160 VSUBS 0.008426f
C1016 B.n161 VSUBS 0.008426f
C1017 B.n162 VSUBS 0.008426f
C1018 B.n163 VSUBS 0.008426f
C1019 B.n164 VSUBS 0.008426f
C1020 B.n165 VSUBS 0.008426f
C1021 B.n166 VSUBS 0.008426f
C1022 B.n167 VSUBS 0.008426f
C1023 B.n168 VSUBS 0.008426f
C1024 B.n169 VSUBS 0.008426f
C1025 B.n170 VSUBS 0.008426f
C1026 B.n171 VSUBS 0.008426f
C1027 B.n172 VSUBS 0.008426f
C1028 B.n173 VSUBS 0.008426f
C1029 B.n174 VSUBS 0.008426f
C1030 B.n175 VSUBS 0.008426f
C1031 B.n176 VSUBS 0.008426f
C1032 B.n177 VSUBS 0.008426f
C1033 B.n178 VSUBS 0.018481f
C1034 B.n179 VSUBS 0.018481f
C1035 B.n180 VSUBS 0.019435f
C1036 B.n181 VSUBS 0.008426f
C1037 B.n182 VSUBS 0.008426f
C1038 B.n183 VSUBS 0.008426f
C1039 B.n184 VSUBS 0.008426f
C1040 B.n185 VSUBS 0.008426f
C1041 B.n186 VSUBS 0.008426f
C1042 B.n187 VSUBS 0.008426f
C1043 B.n188 VSUBS 0.008426f
C1044 B.n189 VSUBS 0.008426f
C1045 B.n190 VSUBS 0.008426f
C1046 B.n191 VSUBS 0.008426f
C1047 B.n192 VSUBS 0.008426f
C1048 B.n193 VSUBS 0.008426f
C1049 B.n194 VSUBS 0.008426f
C1050 B.n195 VSUBS 0.008426f
C1051 B.n196 VSUBS 0.008426f
C1052 B.n197 VSUBS 0.008426f
C1053 B.n198 VSUBS 0.008426f
C1054 B.n199 VSUBS 0.008426f
C1055 B.n200 VSUBS 0.008426f
C1056 B.n201 VSUBS 0.008426f
C1057 B.n202 VSUBS 0.008426f
C1058 B.n203 VSUBS 0.008426f
C1059 B.n204 VSUBS 0.008426f
C1060 B.n205 VSUBS 0.008426f
C1061 B.n206 VSUBS 0.008426f
C1062 B.n207 VSUBS 0.008426f
C1063 B.n208 VSUBS 0.008426f
C1064 B.n209 VSUBS 0.008426f
C1065 B.n210 VSUBS 0.008426f
C1066 B.n211 VSUBS 0.008426f
C1067 B.n212 VSUBS 0.008426f
C1068 B.n213 VSUBS 0.008426f
C1069 B.n214 VSUBS 0.008426f
C1070 B.n215 VSUBS 0.008426f
C1071 B.n216 VSUBS 0.008426f
C1072 B.n217 VSUBS 0.008426f
C1073 B.n218 VSUBS 0.008426f
C1074 B.n219 VSUBS 0.008426f
C1075 B.n220 VSUBS 0.008426f
C1076 B.n221 VSUBS 0.008426f
C1077 B.n222 VSUBS 0.008426f
C1078 B.n223 VSUBS 0.008426f
C1079 B.n224 VSUBS 0.008426f
C1080 B.n225 VSUBS 0.008426f
C1081 B.n226 VSUBS 0.008426f
C1082 B.n227 VSUBS 0.008426f
C1083 B.n228 VSUBS 0.008426f
C1084 B.n229 VSUBS 0.008426f
C1085 B.n230 VSUBS 0.008426f
C1086 B.n231 VSUBS 0.008426f
C1087 B.n232 VSUBS 0.008426f
C1088 B.n233 VSUBS 0.008426f
C1089 B.n234 VSUBS 0.008426f
C1090 B.n235 VSUBS 0.008426f
C1091 B.n236 VSUBS 0.008426f
C1092 B.n237 VSUBS 0.008426f
C1093 B.n238 VSUBS 0.008426f
C1094 B.n239 VSUBS 0.008426f
C1095 B.n240 VSUBS 0.008426f
C1096 B.n241 VSUBS 0.008426f
C1097 B.n242 VSUBS 0.008426f
C1098 B.n243 VSUBS 0.008426f
C1099 B.n244 VSUBS 0.008426f
C1100 B.n245 VSUBS 0.008426f
C1101 B.n246 VSUBS 0.008426f
C1102 B.n247 VSUBS 0.008426f
C1103 B.n248 VSUBS 0.008426f
C1104 B.n249 VSUBS 0.008426f
C1105 B.n250 VSUBS 0.008426f
C1106 B.n251 VSUBS 0.008426f
C1107 B.n252 VSUBS 0.008426f
C1108 B.n253 VSUBS 0.008426f
C1109 B.n254 VSUBS 0.008426f
C1110 B.n255 VSUBS 0.008426f
C1111 B.n256 VSUBS 0.008426f
C1112 B.n257 VSUBS 0.008426f
C1113 B.n258 VSUBS 0.008426f
C1114 B.n259 VSUBS 0.008426f
C1115 B.n260 VSUBS 0.008426f
C1116 B.n261 VSUBS 0.008426f
C1117 B.n262 VSUBS 0.008426f
C1118 B.n263 VSUBS 0.008426f
C1119 B.n264 VSUBS 0.008426f
C1120 B.n265 VSUBS 0.008426f
C1121 B.n266 VSUBS 0.007682f
C1122 B.n267 VSUBS 0.019522f
C1123 B.n268 VSUBS 0.004956f
C1124 B.n269 VSUBS 0.008426f
C1125 B.n270 VSUBS 0.008426f
C1126 B.n271 VSUBS 0.008426f
C1127 B.n272 VSUBS 0.008426f
C1128 B.n273 VSUBS 0.008426f
C1129 B.n274 VSUBS 0.008426f
C1130 B.n275 VSUBS 0.008426f
C1131 B.n276 VSUBS 0.008426f
C1132 B.n277 VSUBS 0.008426f
C1133 B.n278 VSUBS 0.008426f
C1134 B.n279 VSUBS 0.008426f
C1135 B.n280 VSUBS 0.008426f
C1136 B.t8 VSUBS 0.411117f
C1137 B.t7 VSUBS 0.419842f
C1138 B.t6 VSUBS 0.221218f
C1139 B.n281 VSUBS 0.435936f
C1140 B.n282 VSUBS 0.378104f
C1141 B.n283 VSUBS 0.019522f
C1142 B.n284 VSUBS 0.004956f
C1143 B.n285 VSUBS 0.008426f
C1144 B.n286 VSUBS 0.008426f
C1145 B.n287 VSUBS 0.008426f
C1146 B.n288 VSUBS 0.008426f
C1147 B.n289 VSUBS 0.008426f
C1148 B.n290 VSUBS 0.008426f
C1149 B.n291 VSUBS 0.008426f
C1150 B.n292 VSUBS 0.008426f
C1151 B.n293 VSUBS 0.008426f
C1152 B.n294 VSUBS 0.008426f
C1153 B.n295 VSUBS 0.008426f
C1154 B.n296 VSUBS 0.008426f
C1155 B.n297 VSUBS 0.008426f
C1156 B.n298 VSUBS 0.008426f
C1157 B.n299 VSUBS 0.008426f
C1158 B.n300 VSUBS 0.008426f
C1159 B.n301 VSUBS 0.008426f
C1160 B.n302 VSUBS 0.008426f
C1161 B.n303 VSUBS 0.008426f
C1162 B.n304 VSUBS 0.008426f
C1163 B.n305 VSUBS 0.008426f
C1164 B.n306 VSUBS 0.008426f
C1165 B.n307 VSUBS 0.008426f
C1166 B.n308 VSUBS 0.008426f
C1167 B.n309 VSUBS 0.008426f
C1168 B.n310 VSUBS 0.008426f
C1169 B.n311 VSUBS 0.008426f
C1170 B.n312 VSUBS 0.008426f
C1171 B.n313 VSUBS 0.008426f
C1172 B.n314 VSUBS 0.008426f
C1173 B.n315 VSUBS 0.008426f
C1174 B.n316 VSUBS 0.008426f
C1175 B.n317 VSUBS 0.008426f
C1176 B.n318 VSUBS 0.008426f
C1177 B.n319 VSUBS 0.008426f
C1178 B.n320 VSUBS 0.008426f
C1179 B.n321 VSUBS 0.008426f
C1180 B.n322 VSUBS 0.008426f
C1181 B.n323 VSUBS 0.008426f
C1182 B.n324 VSUBS 0.008426f
C1183 B.n325 VSUBS 0.008426f
C1184 B.n326 VSUBS 0.008426f
C1185 B.n327 VSUBS 0.008426f
C1186 B.n328 VSUBS 0.008426f
C1187 B.n329 VSUBS 0.008426f
C1188 B.n330 VSUBS 0.008426f
C1189 B.n331 VSUBS 0.008426f
C1190 B.n332 VSUBS 0.008426f
C1191 B.n333 VSUBS 0.008426f
C1192 B.n334 VSUBS 0.008426f
C1193 B.n335 VSUBS 0.008426f
C1194 B.n336 VSUBS 0.008426f
C1195 B.n337 VSUBS 0.008426f
C1196 B.n338 VSUBS 0.008426f
C1197 B.n339 VSUBS 0.008426f
C1198 B.n340 VSUBS 0.008426f
C1199 B.n341 VSUBS 0.008426f
C1200 B.n342 VSUBS 0.008426f
C1201 B.n343 VSUBS 0.008426f
C1202 B.n344 VSUBS 0.008426f
C1203 B.n345 VSUBS 0.008426f
C1204 B.n346 VSUBS 0.008426f
C1205 B.n347 VSUBS 0.008426f
C1206 B.n348 VSUBS 0.008426f
C1207 B.n349 VSUBS 0.008426f
C1208 B.n350 VSUBS 0.008426f
C1209 B.n351 VSUBS 0.008426f
C1210 B.n352 VSUBS 0.008426f
C1211 B.n353 VSUBS 0.008426f
C1212 B.n354 VSUBS 0.008426f
C1213 B.n355 VSUBS 0.008426f
C1214 B.n356 VSUBS 0.008426f
C1215 B.n357 VSUBS 0.008426f
C1216 B.n358 VSUBS 0.008426f
C1217 B.n359 VSUBS 0.008426f
C1218 B.n360 VSUBS 0.008426f
C1219 B.n361 VSUBS 0.008426f
C1220 B.n362 VSUBS 0.008426f
C1221 B.n363 VSUBS 0.008426f
C1222 B.n364 VSUBS 0.008426f
C1223 B.n365 VSUBS 0.008426f
C1224 B.n366 VSUBS 0.008426f
C1225 B.n367 VSUBS 0.008426f
C1226 B.n368 VSUBS 0.008426f
C1227 B.n369 VSUBS 0.008426f
C1228 B.n370 VSUBS 0.008426f
C1229 B.n371 VSUBS 0.019435f
C1230 B.n372 VSUBS 0.018378f
C1231 B.n373 VSUBS 0.019538f
C1232 B.n374 VSUBS 0.008426f
C1233 B.n375 VSUBS 0.008426f
C1234 B.n376 VSUBS 0.008426f
C1235 B.n377 VSUBS 0.008426f
C1236 B.n378 VSUBS 0.008426f
C1237 B.n379 VSUBS 0.008426f
C1238 B.n380 VSUBS 0.008426f
C1239 B.n381 VSUBS 0.008426f
C1240 B.n382 VSUBS 0.008426f
C1241 B.n383 VSUBS 0.008426f
C1242 B.n384 VSUBS 0.008426f
C1243 B.n385 VSUBS 0.008426f
C1244 B.n386 VSUBS 0.008426f
C1245 B.n387 VSUBS 0.008426f
C1246 B.n388 VSUBS 0.008426f
C1247 B.n389 VSUBS 0.008426f
C1248 B.n390 VSUBS 0.008426f
C1249 B.n391 VSUBS 0.008426f
C1250 B.n392 VSUBS 0.008426f
C1251 B.n393 VSUBS 0.008426f
C1252 B.n394 VSUBS 0.008426f
C1253 B.n395 VSUBS 0.008426f
C1254 B.n396 VSUBS 0.008426f
C1255 B.n397 VSUBS 0.008426f
C1256 B.n398 VSUBS 0.008426f
C1257 B.n399 VSUBS 0.008426f
C1258 B.n400 VSUBS 0.008426f
C1259 B.n401 VSUBS 0.008426f
C1260 B.n402 VSUBS 0.008426f
C1261 B.n403 VSUBS 0.008426f
C1262 B.n404 VSUBS 0.008426f
C1263 B.n405 VSUBS 0.008426f
C1264 B.n406 VSUBS 0.008426f
C1265 B.n407 VSUBS 0.008426f
C1266 B.n408 VSUBS 0.008426f
C1267 B.n409 VSUBS 0.008426f
C1268 B.n410 VSUBS 0.008426f
C1269 B.n411 VSUBS 0.008426f
C1270 B.n412 VSUBS 0.008426f
C1271 B.n413 VSUBS 0.018481f
C1272 B.n414 VSUBS 0.018481f
C1273 B.n415 VSUBS 0.019435f
C1274 B.n416 VSUBS 0.008426f
C1275 B.n417 VSUBS 0.008426f
C1276 B.n418 VSUBS 0.008426f
C1277 B.n419 VSUBS 0.008426f
C1278 B.n420 VSUBS 0.008426f
C1279 B.n421 VSUBS 0.008426f
C1280 B.n422 VSUBS 0.008426f
C1281 B.n423 VSUBS 0.008426f
C1282 B.n424 VSUBS 0.008426f
C1283 B.n425 VSUBS 0.008426f
C1284 B.n426 VSUBS 0.008426f
C1285 B.n427 VSUBS 0.008426f
C1286 B.n428 VSUBS 0.008426f
C1287 B.n429 VSUBS 0.008426f
C1288 B.n430 VSUBS 0.008426f
C1289 B.n431 VSUBS 0.008426f
C1290 B.n432 VSUBS 0.008426f
C1291 B.n433 VSUBS 0.008426f
C1292 B.n434 VSUBS 0.008426f
C1293 B.n435 VSUBS 0.008426f
C1294 B.n436 VSUBS 0.008426f
C1295 B.n437 VSUBS 0.008426f
C1296 B.n438 VSUBS 0.008426f
C1297 B.n439 VSUBS 0.008426f
C1298 B.n440 VSUBS 0.008426f
C1299 B.n441 VSUBS 0.008426f
C1300 B.n442 VSUBS 0.008426f
C1301 B.n443 VSUBS 0.008426f
C1302 B.n444 VSUBS 0.008426f
C1303 B.n445 VSUBS 0.008426f
C1304 B.n446 VSUBS 0.008426f
C1305 B.n447 VSUBS 0.008426f
C1306 B.n448 VSUBS 0.008426f
C1307 B.n449 VSUBS 0.008426f
C1308 B.n450 VSUBS 0.008426f
C1309 B.n451 VSUBS 0.008426f
C1310 B.n452 VSUBS 0.008426f
C1311 B.n453 VSUBS 0.008426f
C1312 B.n454 VSUBS 0.008426f
C1313 B.n455 VSUBS 0.008426f
C1314 B.n456 VSUBS 0.008426f
C1315 B.n457 VSUBS 0.008426f
C1316 B.n458 VSUBS 0.008426f
C1317 B.n459 VSUBS 0.008426f
C1318 B.n460 VSUBS 0.008426f
C1319 B.n461 VSUBS 0.008426f
C1320 B.n462 VSUBS 0.008426f
C1321 B.n463 VSUBS 0.008426f
C1322 B.n464 VSUBS 0.008426f
C1323 B.n465 VSUBS 0.008426f
C1324 B.n466 VSUBS 0.008426f
C1325 B.n467 VSUBS 0.008426f
C1326 B.n468 VSUBS 0.008426f
C1327 B.n469 VSUBS 0.008426f
C1328 B.n470 VSUBS 0.008426f
C1329 B.n471 VSUBS 0.008426f
C1330 B.n472 VSUBS 0.008426f
C1331 B.n473 VSUBS 0.008426f
C1332 B.n474 VSUBS 0.008426f
C1333 B.n475 VSUBS 0.008426f
C1334 B.n476 VSUBS 0.008426f
C1335 B.n477 VSUBS 0.008426f
C1336 B.n478 VSUBS 0.008426f
C1337 B.n479 VSUBS 0.008426f
C1338 B.n480 VSUBS 0.008426f
C1339 B.n481 VSUBS 0.008426f
C1340 B.n482 VSUBS 0.008426f
C1341 B.n483 VSUBS 0.008426f
C1342 B.n484 VSUBS 0.008426f
C1343 B.n485 VSUBS 0.008426f
C1344 B.n486 VSUBS 0.008426f
C1345 B.n487 VSUBS 0.008426f
C1346 B.n488 VSUBS 0.008426f
C1347 B.n489 VSUBS 0.008426f
C1348 B.n490 VSUBS 0.008426f
C1349 B.n491 VSUBS 0.008426f
C1350 B.n492 VSUBS 0.008426f
C1351 B.n493 VSUBS 0.008426f
C1352 B.n494 VSUBS 0.008426f
C1353 B.n495 VSUBS 0.008426f
C1354 B.n496 VSUBS 0.008426f
C1355 B.n497 VSUBS 0.008426f
C1356 B.n498 VSUBS 0.008426f
C1357 B.n499 VSUBS 0.008426f
C1358 B.n500 VSUBS 0.007682f
C1359 B.n501 VSUBS 0.008426f
C1360 B.n502 VSUBS 0.008426f
C1361 B.n503 VSUBS 0.008426f
C1362 B.n504 VSUBS 0.008426f
C1363 B.n505 VSUBS 0.008426f
C1364 B.n506 VSUBS 0.008426f
C1365 B.n507 VSUBS 0.008426f
C1366 B.n508 VSUBS 0.008426f
C1367 B.n509 VSUBS 0.008426f
C1368 B.n510 VSUBS 0.008426f
C1369 B.n511 VSUBS 0.008426f
C1370 B.n512 VSUBS 0.008426f
C1371 B.n513 VSUBS 0.008426f
C1372 B.n514 VSUBS 0.008426f
C1373 B.n515 VSUBS 0.008426f
C1374 B.n516 VSUBS 0.004956f
C1375 B.n517 VSUBS 0.019522f
C1376 B.n518 VSUBS 0.007682f
C1377 B.n519 VSUBS 0.008426f
C1378 B.n520 VSUBS 0.008426f
C1379 B.n521 VSUBS 0.008426f
C1380 B.n522 VSUBS 0.008426f
C1381 B.n523 VSUBS 0.008426f
C1382 B.n524 VSUBS 0.008426f
C1383 B.n525 VSUBS 0.008426f
C1384 B.n526 VSUBS 0.008426f
C1385 B.n527 VSUBS 0.008426f
C1386 B.n528 VSUBS 0.008426f
C1387 B.n529 VSUBS 0.008426f
C1388 B.n530 VSUBS 0.008426f
C1389 B.n531 VSUBS 0.008426f
C1390 B.n532 VSUBS 0.008426f
C1391 B.n533 VSUBS 0.008426f
C1392 B.n534 VSUBS 0.008426f
C1393 B.n535 VSUBS 0.008426f
C1394 B.n536 VSUBS 0.008426f
C1395 B.n537 VSUBS 0.008426f
C1396 B.n538 VSUBS 0.008426f
C1397 B.n539 VSUBS 0.008426f
C1398 B.n540 VSUBS 0.008426f
C1399 B.n541 VSUBS 0.008426f
C1400 B.n542 VSUBS 0.008426f
C1401 B.n543 VSUBS 0.008426f
C1402 B.n544 VSUBS 0.008426f
C1403 B.n545 VSUBS 0.008426f
C1404 B.n546 VSUBS 0.008426f
C1405 B.n547 VSUBS 0.008426f
C1406 B.n548 VSUBS 0.008426f
C1407 B.n549 VSUBS 0.008426f
C1408 B.n550 VSUBS 0.008426f
C1409 B.n551 VSUBS 0.008426f
C1410 B.n552 VSUBS 0.008426f
C1411 B.n553 VSUBS 0.008426f
C1412 B.n554 VSUBS 0.008426f
C1413 B.n555 VSUBS 0.008426f
C1414 B.n556 VSUBS 0.008426f
C1415 B.n557 VSUBS 0.008426f
C1416 B.n558 VSUBS 0.008426f
C1417 B.n559 VSUBS 0.008426f
C1418 B.n560 VSUBS 0.008426f
C1419 B.n561 VSUBS 0.008426f
C1420 B.n562 VSUBS 0.008426f
C1421 B.n563 VSUBS 0.008426f
C1422 B.n564 VSUBS 0.008426f
C1423 B.n565 VSUBS 0.008426f
C1424 B.n566 VSUBS 0.008426f
C1425 B.n567 VSUBS 0.008426f
C1426 B.n568 VSUBS 0.008426f
C1427 B.n569 VSUBS 0.008426f
C1428 B.n570 VSUBS 0.008426f
C1429 B.n571 VSUBS 0.008426f
C1430 B.n572 VSUBS 0.008426f
C1431 B.n573 VSUBS 0.008426f
C1432 B.n574 VSUBS 0.008426f
C1433 B.n575 VSUBS 0.008426f
C1434 B.n576 VSUBS 0.008426f
C1435 B.n577 VSUBS 0.008426f
C1436 B.n578 VSUBS 0.008426f
C1437 B.n579 VSUBS 0.008426f
C1438 B.n580 VSUBS 0.008426f
C1439 B.n581 VSUBS 0.008426f
C1440 B.n582 VSUBS 0.008426f
C1441 B.n583 VSUBS 0.008426f
C1442 B.n584 VSUBS 0.008426f
C1443 B.n585 VSUBS 0.008426f
C1444 B.n586 VSUBS 0.008426f
C1445 B.n587 VSUBS 0.008426f
C1446 B.n588 VSUBS 0.008426f
C1447 B.n589 VSUBS 0.008426f
C1448 B.n590 VSUBS 0.008426f
C1449 B.n591 VSUBS 0.008426f
C1450 B.n592 VSUBS 0.008426f
C1451 B.n593 VSUBS 0.008426f
C1452 B.n594 VSUBS 0.008426f
C1453 B.n595 VSUBS 0.008426f
C1454 B.n596 VSUBS 0.008426f
C1455 B.n597 VSUBS 0.008426f
C1456 B.n598 VSUBS 0.008426f
C1457 B.n599 VSUBS 0.008426f
C1458 B.n600 VSUBS 0.008426f
C1459 B.n601 VSUBS 0.008426f
C1460 B.n602 VSUBS 0.008426f
C1461 B.n603 VSUBS 0.019435f
C1462 B.n604 VSUBS 0.019435f
C1463 B.n605 VSUBS 0.018481f
C1464 B.n606 VSUBS 0.008426f
C1465 B.n607 VSUBS 0.008426f
C1466 B.n608 VSUBS 0.008426f
C1467 B.n609 VSUBS 0.008426f
C1468 B.n610 VSUBS 0.008426f
C1469 B.n611 VSUBS 0.008426f
C1470 B.n612 VSUBS 0.008426f
C1471 B.n613 VSUBS 0.008426f
C1472 B.n614 VSUBS 0.008426f
C1473 B.n615 VSUBS 0.008426f
C1474 B.n616 VSUBS 0.008426f
C1475 B.n617 VSUBS 0.008426f
C1476 B.n618 VSUBS 0.008426f
C1477 B.n619 VSUBS 0.008426f
C1478 B.n620 VSUBS 0.008426f
C1479 B.n621 VSUBS 0.008426f
C1480 B.n622 VSUBS 0.008426f
C1481 B.n623 VSUBS 0.010995f
C1482 B.n624 VSUBS 0.011713f
C1483 B.n625 VSUBS 0.023292f
.ends

