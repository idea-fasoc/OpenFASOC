* NGSPICE file created from diff_pair_sample_1054.ext - technology: sky130A

.subckt diff_pair_sample_1054 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X1 VTAIL.t18 VP.t1 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=0 ps=0 w=17.62 l=2.35
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=0 ps=0 w=17.62 l=2.35
X4 VDD1.t5 VP.t2 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X5 VDD1.t4 VP.t3 VTAIL.t16 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X6 VTAIL.t0 VN.t0 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X7 VDD1.t1 VP.t4 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=6.8718 ps=36.02 w=17.62 l=2.35
X8 VTAIL.t14 VP.t5 VDD1.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X9 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X10 VTAIL.t13 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X11 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X12 VDD2.t6 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=6.8718 ps=36.02 w=17.62 l=2.35
X13 VDD2.t5 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=6.8718 ps=36.02 w=17.62 l=2.35
X14 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X15 VDD1.t2 VP.t7 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=2.9073 ps=17.95 w=17.62 l=2.35
X16 VDD1.t7 VP.t8 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=6.8718 ps=36.02 w=17.62 l=2.35
X17 VDD2.t3 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=2.9073 ps=17.95 w=17.62 l=2.35
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=0 ps=0 w=17.62 l=2.35
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=0 ps=0 w=17.62 l=2.35
X20 VTAIL.t5 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X21 VTAIL.t4 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9073 pd=17.95 as=2.9073 ps=17.95 w=17.62 l=2.35
X22 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=2.9073 ps=17.95 w=17.62 l=2.35
X23 VDD1.t6 VP.t9 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8718 pd=36.02 as=2.9073 ps=17.95 w=17.62 l=2.35
R0 VP.n19 VP.t7 214.102
R1 VP.n5 VP.t2 180.7
R2 VP.n49 VP.t9 180.7
R3 VP.n57 VP.t0 180.7
R4 VP.n75 VP.t5 180.7
R5 VP.n83 VP.t4 180.7
R6 VP.n16 VP.t3 180.7
R7 VP.n46 VP.t8 180.7
R8 VP.n38 VP.t1 180.7
R9 VP.n20 VP.t6 180.7
R10 VP.n22 VP.n21 161.3
R11 VP.n23 VP.n18 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n26 VP.n17 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n29 VP.n16 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n32 VP.n15 161.3
R18 VP.n34 VP.n33 161.3
R19 VP.n35 VP.n14 161.3
R20 VP.n37 VP.n36 161.3
R21 VP.n39 VP.n13 161.3
R22 VP.n41 VP.n40 161.3
R23 VP.n42 VP.n12 161.3
R24 VP.n44 VP.n43 161.3
R25 VP.n45 VP.n11 161.3
R26 VP.n82 VP.n0 161.3
R27 VP.n81 VP.n80 161.3
R28 VP.n79 VP.n1 161.3
R29 VP.n78 VP.n77 161.3
R30 VP.n76 VP.n2 161.3
R31 VP.n74 VP.n73 161.3
R32 VP.n72 VP.n3 161.3
R33 VP.n71 VP.n70 161.3
R34 VP.n69 VP.n4 161.3
R35 VP.n68 VP.n67 161.3
R36 VP.n66 VP.n5 161.3
R37 VP.n65 VP.n64 161.3
R38 VP.n63 VP.n6 161.3
R39 VP.n62 VP.n61 161.3
R40 VP.n60 VP.n7 161.3
R41 VP.n59 VP.n58 161.3
R42 VP.n56 VP.n8 161.3
R43 VP.n55 VP.n54 161.3
R44 VP.n53 VP.n9 161.3
R45 VP.n52 VP.n51 161.3
R46 VP.n50 VP.n10 161.3
R47 VP.n49 VP.n48 93.2021
R48 VP.n84 VP.n83 93.2021
R49 VP.n47 VP.n46 93.2021
R50 VP.n20 VP.n19 63.1823
R51 VP.n48 VP.n47 56.0906
R52 VP.n63 VP.n62 56.0773
R53 VP.n70 VP.n69 56.0773
R54 VP.n33 VP.n32 56.0773
R55 VP.n26 VP.n25 56.0773
R56 VP.n51 VP.n9 42.5146
R57 VP.n81 VP.n1 42.5146
R58 VP.n44 VP.n12 42.5146
R59 VP.n55 VP.n9 38.6395
R60 VP.n77 VP.n1 38.6395
R61 VP.n40 VP.n12 38.6395
R62 VP.n62 VP.n7 25.0767
R63 VP.n70 VP.n3 25.0767
R64 VP.n33 VP.n14 25.0767
R65 VP.n25 VP.n18 25.0767
R66 VP.n51 VP.n50 24.5923
R67 VP.n56 VP.n55 24.5923
R68 VP.n58 VP.n7 24.5923
R69 VP.n64 VP.n63 24.5923
R70 VP.n64 VP.n5 24.5923
R71 VP.n68 VP.n5 24.5923
R72 VP.n69 VP.n68 24.5923
R73 VP.n74 VP.n3 24.5923
R74 VP.n77 VP.n76 24.5923
R75 VP.n82 VP.n81 24.5923
R76 VP.n45 VP.n44 24.5923
R77 VP.n37 VP.n14 24.5923
R78 VP.n40 VP.n39 24.5923
R79 VP.n27 VP.n26 24.5923
R80 VP.n27 VP.n16 24.5923
R81 VP.n31 VP.n16 24.5923
R82 VP.n32 VP.n31 24.5923
R83 VP.n21 VP.n18 24.5923
R84 VP.n50 VP.n49 17.7066
R85 VP.n83 VP.n82 17.7066
R86 VP.n46 VP.n45 17.7066
R87 VP.n57 VP.n56 15.7393
R88 VP.n76 VP.n75 15.7393
R89 VP.n39 VP.n38 15.7393
R90 VP.n22 VP.n19 9.19198
R91 VP.n58 VP.n57 8.85356
R92 VP.n75 VP.n74 8.85356
R93 VP.n38 VP.n37 8.85356
R94 VP.n21 VP.n20 8.85356
R95 VP.n47 VP.n11 0.278335
R96 VP.n48 VP.n10 0.278335
R97 VP.n84 VP.n0 0.278335
R98 VP.n23 VP.n22 0.189894
R99 VP.n24 VP.n23 0.189894
R100 VP.n24 VP.n17 0.189894
R101 VP.n28 VP.n17 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n30 VP.n29 0.189894
R104 VP.n30 VP.n15 0.189894
R105 VP.n34 VP.n15 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n13 0.189894
R109 VP.n41 VP.n13 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n43 VP.n11 0.189894
R113 VP.n52 VP.n10 0.189894
R114 VP.n53 VP.n52 0.189894
R115 VP.n54 VP.n53 0.189894
R116 VP.n54 VP.n8 0.189894
R117 VP.n59 VP.n8 0.189894
R118 VP.n60 VP.n59 0.189894
R119 VP.n61 VP.n60 0.189894
R120 VP.n61 VP.n6 0.189894
R121 VP.n65 VP.n6 0.189894
R122 VP.n66 VP.n65 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n67 VP.n4 0.189894
R125 VP.n71 VP.n4 0.189894
R126 VP.n72 VP.n71 0.189894
R127 VP.n73 VP.n72 0.189894
R128 VP.n73 VP.n2 0.189894
R129 VP.n78 VP.n2 0.189894
R130 VP.n79 VP.n78 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n80 VP.n0 0.189894
R133 VP VP.n84 0.153485
R134 VDD1.n92 VDD1.n0 289.615
R135 VDD1.n191 VDD1.n99 289.615
R136 VDD1.n93 VDD1.n92 185
R137 VDD1.n91 VDD1.n90 185
R138 VDD1.n4 VDD1.n3 185
R139 VDD1.n85 VDD1.n84 185
R140 VDD1.n83 VDD1.n82 185
R141 VDD1.n8 VDD1.n7 185
R142 VDD1.n12 VDD1.n10 185
R143 VDD1.n77 VDD1.n76 185
R144 VDD1.n75 VDD1.n74 185
R145 VDD1.n14 VDD1.n13 185
R146 VDD1.n69 VDD1.n68 185
R147 VDD1.n67 VDD1.n66 185
R148 VDD1.n18 VDD1.n17 185
R149 VDD1.n61 VDD1.n60 185
R150 VDD1.n59 VDD1.n58 185
R151 VDD1.n22 VDD1.n21 185
R152 VDD1.n53 VDD1.n52 185
R153 VDD1.n51 VDD1.n50 185
R154 VDD1.n26 VDD1.n25 185
R155 VDD1.n45 VDD1.n44 185
R156 VDD1.n43 VDD1.n42 185
R157 VDD1.n30 VDD1.n29 185
R158 VDD1.n37 VDD1.n36 185
R159 VDD1.n35 VDD1.n34 185
R160 VDD1.n132 VDD1.n131 185
R161 VDD1.n134 VDD1.n133 185
R162 VDD1.n127 VDD1.n126 185
R163 VDD1.n140 VDD1.n139 185
R164 VDD1.n142 VDD1.n141 185
R165 VDD1.n123 VDD1.n122 185
R166 VDD1.n148 VDD1.n147 185
R167 VDD1.n150 VDD1.n149 185
R168 VDD1.n119 VDD1.n118 185
R169 VDD1.n156 VDD1.n155 185
R170 VDD1.n158 VDD1.n157 185
R171 VDD1.n115 VDD1.n114 185
R172 VDD1.n164 VDD1.n163 185
R173 VDD1.n166 VDD1.n165 185
R174 VDD1.n111 VDD1.n110 185
R175 VDD1.n173 VDD1.n172 185
R176 VDD1.n174 VDD1.n109 185
R177 VDD1.n176 VDD1.n175 185
R178 VDD1.n107 VDD1.n106 185
R179 VDD1.n182 VDD1.n181 185
R180 VDD1.n184 VDD1.n183 185
R181 VDD1.n103 VDD1.n102 185
R182 VDD1.n190 VDD1.n189 185
R183 VDD1.n192 VDD1.n191 185
R184 VDD1.n33 VDD1.t2 147.659
R185 VDD1.n130 VDD1.t6 147.659
R186 VDD1.n92 VDD1.n91 104.615
R187 VDD1.n91 VDD1.n3 104.615
R188 VDD1.n84 VDD1.n3 104.615
R189 VDD1.n84 VDD1.n83 104.615
R190 VDD1.n83 VDD1.n7 104.615
R191 VDD1.n12 VDD1.n7 104.615
R192 VDD1.n76 VDD1.n12 104.615
R193 VDD1.n76 VDD1.n75 104.615
R194 VDD1.n75 VDD1.n13 104.615
R195 VDD1.n68 VDD1.n13 104.615
R196 VDD1.n68 VDD1.n67 104.615
R197 VDD1.n67 VDD1.n17 104.615
R198 VDD1.n60 VDD1.n17 104.615
R199 VDD1.n60 VDD1.n59 104.615
R200 VDD1.n59 VDD1.n21 104.615
R201 VDD1.n52 VDD1.n21 104.615
R202 VDD1.n52 VDD1.n51 104.615
R203 VDD1.n51 VDD1.n25 104.615
R204 VDD1.n44 VDD1.n25 104.615
R205 VDD1.n44 VDD1.n43 104.615
R206 VDD1.n43 VDD1.n29 104.615
R207 VDD1.n36 VDD1.n29 104.615
R208 VDD1.n36 VDD1.n35 104.615
R209 VDD1.n133 VDD1.n132 104.615
R210 VDD1.n133 VDD1.n126 104.615
R211 VDD1.n140 VDD1.n126 104.615
R212 VDD1.n141 VDD1.n140 104.615
R213 VDD1.n141 VDD1.n122 104.615
R214 VDD1.n148 VDD1.n122 104.615
R215 VDD1.n149 VDD1.n148 104.615
R216 VDD1.n149 VDD1.n118 104.615
R217 VDD1.n156 VDD1.n118 104.615
R218 VDD1.n157 VDD1.n156 104.615
R219 VDD1.n157 VDD1.n114 104.615
R220 VDD1.n164 VDD1.n114 104.615
R221 VDD1.n165 VDD1.n164 104.615
R222 VDD1.n165 VDD1.n110 104.615
R223 VDD1.n173 VDD1.n110 104.615
R224 VDD1.n174 VDD1.n173 104.615
R225 VDD1.n175 VDD1.n174 104.615
R226 VDD1.n175 VDD1.n106 104.615
R227 VDD1.n182 VDD1.n106 104.615
R228 VDD1.n183 VDD1.n182 104.615
R229 VDD1.n183 VDD1.n102 104.615
R230 VDD1.n190 VDD1.n102 104.615
R231 VDD1.n191 VDD1.n190 104.615
R232 VDD1.n199 VDD1.n198 64.2988
R233 VDD1.n98 VDD1.n97 62.6215
R234 VDD1.n197 VDD1.n196 62.6214
R235 VDD1.n201 VDD1.n200 62.6214
R236 VDD1.n98 VDD1.n96 53.1139
R237 VDD1.n197 VDD1.n195 53.1139
R238 VDD1.n35 VDD1.t2 52.3082
R239 VDD1.n132 VDD1.t6 52.3082
R240 VDD1.n201 VDD1.n199 51.6173
R241 VDD1.n34 VDD1.n33 15.6677
R242 VDD1.n131 VDD1.n130 15.6677
R243 VDD1.n10 VDD1.n8 13.1884
R244 VDD1.n176 VDD1.n107 13.1884
R245 VDD1.n82 VDD1.n81 12.8005
R246 VDD1.n78 VDD1.n77 12.8005
R247 VDD1.n37 VDD1.n32 12.8005
R248 VDD1.n134 VDD1.n129 12.8005
R249 VDD1.n177 VDD1.n109 12.8005
R250 VDD1.n181 VDD1.n180 12.8005
R251 VDD1.n85 VDD1.n6 12.0247
R252 VDD1.n74 VDD1.n11 12.0247
R253 VDD1.n38 VDD1.n30 12.0247
R254 VDD1.n135 VDD1.n127 12.0247
R255 VDD1.n172 VDD1.n171 12.0247
R256 VDD1.n184 VDD1.n105 12.0247
R257 VDD1.n86 VDD1.n4 11.249
R258 VDD1.n73 VDD1.n14 11.249
R259 VDD1.n42 VDD1.n41 11.249
R260 VDD1.n139 VDD1.n138 11.249
R261 VDD1.n170 VDD1.n111 11.249
R262 VDD1.n185 VDD1.n103 11.249
R263 VDD1.n90 VDD1.n89 10.4732
R264 VDD1.n70 VDD1.n69 10.4732
R265 VDD1.n45 VDD1.n28 10.4732
R266 VDD1.n142 VDD1.n125 10.4732
R267 VDD1.n167 VDD1.n166 10.4732
R268 VDD1.n189 VDD1.n188 10.4732
R269 VDD1.n93 VDD1.n2 9.69747
R270 VDD1.n66 VDD1.n16 9.69747
R271 VDD1.n46 VDD1.n26 9.69747
R272 VDD1.n143 VDD1.n123 9.69747
R273 VDD1.n163 VDD1.n113 9.69747
R274 VDD1.n192 VDD1.n101 9.69747
R275 VDD1.n96 VDD1.n95 9.45567
R276 VDD1.n195 VDD1.n194 9.45567
R277 VDD1.n20 VDD1.n19 9.3005
R278 VDD1.n63 VDD1.n62 9.3005
R279 VDD1.n65 VDD1.n64 9.3005
R280 VDD1.n16 VDD1.n15 9.3005
R281 VDD1.n71 VDD1.n70 9.3005
R282 VDD1.n73 VDD1.n72 9.3005
R283 VDD1.n11 VDD1.n9 9.3005
R284 VDD1.n79 VDD1.n78 9.3005
R285 VDD1.n95 VDD1.n94 9.3005
R286 VDD1.n2 VDD1.n1 9.3005
R287 VDD1.n89 VDD1.n88 9.3005
R288 VDD1.n87 VDD1.n86 9.3005
R289 VDD1.n6 VDD1.n5 9.3005
R290 VDD1.n81 VDD1.n80 9.3005
R291 VDD1.n57 VDD1.n56 9.3005
R292 VDD1.n55 VDD1.n54 9.3005
R293 VDD1.n24 VDD1.n23 9.3005
R294 VDD1.n49 VDD1.n48 9.3005
R295 VDD1.n47 VDD1.n46 9.3005
R296 VDD1.n28 VDD1.n27 9.3005
R297 VDD1.n41 VDD1.n40 9.3005
R298 VDD1.n39 VDD1.n38 9.3005
R299 VDD1.n32 VDD1.n31 9.3005
R300 VDD1.n194 VDD1.n193 9.3005
R301 VDD1.n101 VDD1.n100 9.3005
R302 VDD1.n188 VDD1.n187 9.3005
R303 VDD1.n186 VDD1.n185 9.3005
R304 VDD1.n105 VDD1.n104 9.3005
R305 VDD1.n180 VDD1.n179 9.3005
R306 VDD1.n152 VDD1.n151 9.3005
R307 VDD1.n121 VDD1.n120 9.3005
R308 VDD1.n146 VDD1.n145 9.3005
R309 VDD1.n144 VDD1.n143 9.3005
R310 VDD1.n125 VDD1.n124 9.3005
R311 VDD1.n138 VDD1.n137 9.3005
R312 VDD1.n136 VDD1.n135 9.3005
R313 VDD1.n129 VDD1.n128 9.3005
R314 VDD1.n154 VDD1.n153 9.3005
R315 VDD1.n117 VDD1.n116 9.3005
R316 VDD1.n160 VDD1.n159 9.3005
R317 VDD1.n162 VDD1.n161 9.3005
R318 VDD1.n113 VDD1.n112 9.3005
R319 VDD1.n168 VDD1.n167 9.3005
R320 VDD1.n170 VDD1.n169 9.3005
R321 VDD1.n171 VDD1.n108 9.3005
R322 VDD1.n178 VDD1.n177 9.3005
R323 VDD1.n94 VDD1.n0 8.92171
R324 VDD1.n65 VDD1.n18 8.92171
R325 VDD1.n50 VDD1.n49 8.92171
R326 VDD1.n147 VDD1.n146 8.92171
R327 VDD1.n162 VDD1.n115 8.92171
R328 VDD1.n193 VDD1.n99 8.92171
R329 VDD1.n62 VDD1.n61 8.14595
R330 VDD1.n53 VDD1.n24 8.14595
R331 VDD1.n150 VDD1.n121 8.14595
R332 VDD1.n159 VDD1.n158 8.14595
R333 VDD1.n58 VDD1.n20 7.3702
R334 VDD1.n54 VDD1.n22 7.3702
R335 VDD1.n151 VDD1.n119 7.3702
R336 VDD1.n155 VDD1.n117 7.3702
R337 VDD1.n58 VDD1.n57 6.59444
R338 VDD1.n57 VDD1.n22 6.59444
R339 VDD1.n154 VDD1.n119 6.59444
R340 VDD1.n155 VDD1.n154 6.59444
R341 VDD1.n61 VDD1.n20 5.81868
R342 VDD1.n54 VDD1.n53 5.81868
R343 VDD1.n151 VDD1.n150 5.81868
R344 VDD1.n158 VDD1.n117 5.81868
R345 VDD1.n96 VDD1.n0 5.04292
R346 VDD1.n62 VDD1.n18 5.04292
R347 VDD1.n50 VDD1.n24 5.04292
R348 VDD1.n147 VDD1.n121 5.04292
R349 VDD1.n159 VDD1.n115 5.04292
R350 VDD1.n195 VDD1.n99 5.04292
R351 VDD1.n33 VDD1.n31 4.38563
R352 VDD1.n130 VDD1.n128 4.38563
R353 VDD1.n94 VDD1.n93 4.26717
R354 VDD1.n66 VDD1.n65 4.26717
R355 VDD1.n49 VDD1.n26 4.26717
R356 VDD1.n146 VDD1.n123 4.26717
R357 VDD1.n163 VDD1.n162 4.26717
R358 VDD1.n193 VDD1.n192 4.26717
R359 VDD1.n90 VDD1.n2 3.49141
R360 VDD1.n69 VDD1.n16 3.49141
R361 VDD1.n46 VDD1.n45 3.49141
R362 VDD1.n143 VDD1.n142 3.49141
R363 VDD1.n166 VDD1.n113 3.49141
R364 VDD1.n189 VDD1.n101 3.49141
R365 VDD1.n89 VDD1.n4 2.71565
R366 VDD1.n70 VDD1.n14 2.71565
R367 VDD1.n42 VDD1.n28 2.71565
R368 VDD1.n139 VDD1.n125 2.71565
R369 VDD1.n167 VDD1.n111 2.71565
R370 VDD1.n188 VDD1.n103 2.71565
R371 VDD1.n86 VDD1.n85 1.93989
R372 VDD1.n74 VDD1.n73 1.93989
R373 VDD1.n41 VDD1.n30 1.93989
R374 VDD1.n138 VDD1.n127 1.93989
R375 VDD1.n172 VDD1.n170 1.93989
R376 VDD1.n185 VDD1.n184 1.93989
R377 VDD1 VDD1.n201 1.67507
R378 VDD1.n82 VDD1.n6 1.16414
R379 VDD1.n77 VDD1.n11 1.16414
R380 VDD1.n38 VDD1.n37 1.16414
R381 VDD1.n135 VDD1.n134 1.16414
R382 VDD1.n171 VDD1.n109 1.16414
R383 VDD1.n181 VDD1.n105 1.16414
R384 VDD1.n200 VDD1.t8 1.12422
R385 VDD1.n200 VDD1.t7 1.12422
R386 VDD1.n97 VDD1.t3 1.12422
R387 VDD1.n97 VDD1.t4 1.12422
R388 VDD1.n198 VDD1.t0 1.12422
R389 VDD1.n198 VDD1.t1 1.12422
R390 VDD1.n196 VDD1.t9 1.12422
R391 VDD1.n196 VDD1.t5 1.12422
R392 VDD1 VDD1.n98 0.636276
R393 VDD1.n199 VDD1.n197 0.52274
R394 VDD1.n81 VDD1.n8 0.388379
R395 VDD1.n78 VDD1.n10 0.388379
R396 VDD1.n34 VDD1.n32 0.388379
R397 VDD1.n131 VDD1.n129 0.388379
R398 VDD1.n177 VDD1.n176 0.388379
R399 VDD1.n180 VDD1.n107 0.388379
R400 VDD1.n95 VDD1.n1 0.155672
R401 VDD1.n88 VDD1.n1 0.155672
R402 VDD1.n88 VDD1.n87 0.155672
R403 VDD1.n87 VDD1.n5 0.155672
R404 VDD1.n80 VDD1.n5 0.155672
R405 VDD1.n80 VDD1.n79 0.155672
R406 VDD1.n79 VDD1.n9 0.155672
R407 VDD1.n72 VDD1.n9 0.155672
R408 VDD1.n72 VDD1.n71 0.155672
R409 VDD1.n71 VDD1.n15 0.155672
R410 VDD1.n64 VDD1.n15 0.155672
R411 VDD1.n64 VDD1.n63 0.155672
R412 VDD1.n63 VDD1.n19 0.155672
R413 VDD1.n56 VDD1.n19 0.155672
R414 VDD1.n56 VDD1.n55 0.155672
R415 VDD1.n55 VDD1.n23 0.155672
R416 VDD1.n48 VDD1.n23 0.155672
R417 VDD1.n48 VDD1.n47 0.155672
R418 VDD1.n47 VDD1.n27 0.155672
R419 VDD1.n40 VDD1.n27 0.155672
R420 VDD1.n40 VDD1.n39 0.155672
R421 VDD1.n39 VDD1.n31 0.155672
R422 VDD1.n136 VDD1.n128 0.155672
R423 VDD1.n137 VDD1.n136 0.155672
R424 VDD1.n137 VDD1.n124 0.155672
R425 VDD1.n144 VDD1.n124 0.155672
R426 VDD1.n145 VDD1.n144 0.155672
R427 VDD1.n145 VDD1.n120 0.155672
R428 VDD1.n152 VDD1.n120 0.155672
R429 VDD1.n153 VDD1.n152 0.155672
R430 VDD1.n153 VDD1.n116 0.155672
R431 VDD1.n160 VDD1.n116 0.155672
R432 VDD1.n161 VDD1.n160 0.155672
R433 VDD1.n161 VDD1.n112 0.155672
R434 VDD1.n168 VDD1.n112 0.155672
R435 VDD1.n169 VDD1.n168 0.155672
R436 VDD1.n169 VDD1.n108 0.155672
R437 VDD1.n178 VDD1.n108 0.155672
R438 VDD1.n179 VDD1.n178 0.155672
R439 VDD1.n179 VDD1.n104 0.155672
R440 VDD1.n186 VDD1.n104 0.155672
R441 VDD1.n187 VDD1.n186 0.155672
R442 VDD1.n187 VDD1.n100 0.155672
R443 VDD1.n194 VDD1.n100 0.155672
R444 VTAIL.n400 VTAIL.n308 289.615
R445 VTAIL.n94 VTAIL.n2 289.615
R446 VTAIL.n302 VTAIL.n210 289.615
R447 VTAIL.n200 VTAIL.n108 289.615
R448 VTAIL.n341 VTAIL.n340 185
R449 VTAIL.n343 VTAIL.n342 185
R450 VTAIL.n336 VTAIL.n335 185
R451 VTAIL.n349 VTAIL.n348 185
R452 VTAIL.n351 VTAIL.n350 185
R453 VTAIL.n332 VTAIL.n331 185
R454 VTAIL.n357 VTAIL.n356 185
R455 VTAIL.n359 VTAIL.n358 185
R456 VTAIL.n328 VTAIL.n327 185
R457 VTAIL.n365 VTAIL.n364 185
R458 VTAIL.n367 VTAIL.n366 185
R459 VTAIL.n324 VTAIL.n323 185
R460 VTAIL.n373 VTAIL.n372 185
R461 VTAIL.n375 VTAIL.n374 185
R462 VTAIL.n320 VTAIL.n319 185
R463 VTAIL.n382 VTAIL.n381 185
R464 VTAIL.n383 VTAIL.n318 185
R465 VTAIL.n385 VTAIL.n384 185
R466 VTAIL.n316 VTAIL.n315 185
R467 VTAIL.n391 VTAIL.n390 185
R468 VTAIL.n393 VTAIL.n392 185
R469 VTAIL.n312 VTAIL.n311 185
R470 VTAIL.n399 VTAIL.n398 185
R471 VTAIL.n401 VTAIL.n400 185
R472 VTAIL.n35 VTAIL.n34 185
R473 VTAIL.n37 VTAIL.n36 185
R474 VTAIL.n30 VTAIL.n29 185
R475 VTAIL.n43 VTAIL.n42 185
R476 VTAIL.n45 VTAIL.n44 185
R477 VTAIL.n26 VTAIL.n25 185
R478 VTAIL.n51 VTAIL.n50 185
R479 VTAIL.n53 VTAIL.n52 185
R480 VTAIL.n22 VTAIL.n21 185
R481 VTAIL.n59 VTAIL.n58 185
R482 VTAIL.n61 VTAIL.n60 185
R483 VTAIL.n18 VTAIL.n17 185
R484 VTAIL.n67 VTAIL.n66 185
R485 VTAIL.n69 VTAIL.n68 185
R486 VTAIL.n14 VTAIL.n13 185
R487 VTAIL.n76 VTAIL.n75 185
R488 VTAIL.n77 VTAIL.n12 185
R489 VTAIL.n79 VTAIL.n78 185
R490 VTAIL.n10 VTAIL.n9 185
R491 VTAIL.n85 VTAIL.n84 185
R492 VTAIL.n87 VTAIL.n86 185
R493 VTAIL.n6 VTAIL.n5 185
R494 VTAIL.n93 VTAIL.n92 185
R495 VTAIL.n95 VTAIL.n94 185
R496 VTAIL.n303 VTAIL.n302 185
R497 VTAIL.n301 VTAIL.n300 185
R498 VTAIL.n214 VTAIL.n213 185
R499 VTAIL.n295 VTAIL.n294 185
R500 VTAIL.n293 VTAIL.n292 185
R501 VTAIL.n218 VTAIL.n217 185
R502 VTAIL.n222 VTAIL.n220 185
R503 VTAIL.n287 VTAIL.n286 185
R504 VTAIL.n285 VTAIL.n284 185
R505 VTAIL.n224 VTAIL.n223 185
R506 VTAIL.n279 VTAIL.n278 185
R507 VTAIL.n277 VTAIL.n276 185
R508 VTAIL.n228 VTAIL.n227 185
R509 VTAIL.n271 VTAIL.n270 185
R510 VTAIL.n269 VTAIL.n268 185
R511 VTAIL.n232 VTAIL.n231 185
R512 VTAIL.n263 VTAIL.n262 185
R513 VTAIL.n261 VTAIL.n260 185
R514 VTAIL.n236 VTAIL.n235 185
R515 VTAIL.n255 VTAIL.n254 185
R516 VTAIL.n253 VTAIL.n252 185
R517 VTAIL.n240 VTAIL.n239 185
R518 VTAIL.n247 VTAIL.n246 185
R519 VTAIL.n245 VTAIL.n244 185
R520 VTAIL.n201 VTAIL.n200 185
R521 VTAIL.n199 VTAIL.n198 185
R522 VTAIL.n112 VTAIL.n111 185
R523 VTAIL.n193 VTAIL.n192 185
R524 VTAIL.n191 VTAIL.n190 185
R525 VTAIL.n116 VTAIL.n115 185
R526 VTAIL.n120 VTAIL.n118 185
R527 VTAIL.n185 VTAIL.n184 185
R528 VTAIL.n183 VTAIL.n182 185
R529 VTAIL.n122 VTAIL.n121 185
R530 VTAIL.n177 VTAIL.n176 185
R531 VTAIL.n175 VTAIL.n174 185
R532 VTAIL.n126 VTAIL.n125 185
R533 VTAIL.n169 VTAIL.n168 185
R534 VTAIL.n167 VTAIL.n166 185
R535 VTAIL.n130 VTAIL.n129 185
R536 VTAIL.n161 VTAIL.n160 185
R537 VTAIL.n159 VTAIL.n158 185
R538 VTAIL.n134 VTAIL.n133 185
R539 VTAIL.n153 VTAIL.n152 185
R540 VTAIL.n151 VTAIL.n150 185
R541 VTAIL.n138 VTAIL.n137 185
R542 VTAIL.n145 VTAIL.n144 185
R543 VTAIL.n143 VTAIL.n142 185
R544 VTAIL.n339 VTAIL.t2 147.659
R545 VTAIL.n33 VTAIL.t15 147.659
R546 VTAIL.n243 VTAIL.t11 147.659
R547 VTAIL.n141 VTAIL.t3 147.659
R548 VTAIL.n342 VTAIL.n341 104.615
R549 VTAIL.n342 VTAIL.n335 104.615
R550 VTAIL.n349 VTAIL.n335 104.615
R551 VTAIL.n350 VTAIL.n349 104.615
R552 VTAIL.n350 VTAIL.n331 104.615
R553 VTAIL.n357 VTAIL.n331 104.615
R554 VTAIL.n358 VTAIL.n357 104.615
R555 VTAIL.n358 VTAIL.n327 104.615
R556 VTAIL.n365 VTAIL.n327 104.615
R557 VTAIL.n366 VTAIL.n365 104.615
R558 VTAIL.n366 VTAIL.n323 104.615
R559 VTAIL.n373 VTAIL.n323 104.615
R560 VTAIL.n374 VTAIL.n373 104.615
R561 VTAIL.n374 VTAIL.n319 104.615
R562 VTAIL.n382 VTAIL.n319 104.615
R563 VTAIL.n383 VTAIL.n382 104.615
R564 VTAIL.n384 VTAIL.n383 104.615
R565 VTAIL.n384 VTAIL.n315 104.615
R566 VTAIL.n391 VTAIL.n315 104.615
R567 VTAIL.n392 VTAIL.n391 104.615
R568 VTAIL.n392 VTAIL.n311 104.615
R569 VTAIL.n399 VTAIL.n311 104.615
R570 VTAIL.n400 VTAIL.n399 104.615
R571 VTAIL.n36 VTAIL.n35 104.615
R572 VTAIL.n36 VTAIL.n29 104.615
R573 VTAIL.n43 VTAIL.n29 104.615
R574 VTAIL.n44 VTAIL.n43 104.615
R575 VTAIL.n44 VTAIL.n25 104.615
R576 VTAIL.n51 VTAIL.n25 104.615
R577 VTAIL.n52 VTAIL.n51 104.615
R578 VTAIL.n52 VTAIL.n21 104.615
R579 VTAIL.n59 VTAIL.n21 104.615
R580 VTAIL.n60 VTAIL.n59 104.615
R581 VTAIL.n60 VTAIL.n17 104.615
R582 VTAIL.n67 VTAIL.n17 104.615
R583 VTAIL.n68 VTAIL.n67 104.615
R584 VTAIL.n68 VTAIL.n13 104.615
R585 VTAIL.n76 VTAIL.n13 104.615
R586 VTAIL.n77 VTAIL.n76 104.615
R587 VTAIL.n78 VTAIL.n77 104.615
R588 VTAIL.n78 VTAIL.n9 104.615
R589 VTAIL.n85 VTAIL.n9 104.615
R590 VTAIL.n86 VTAIL.n85 104.615
R591 VTAIL.n86 VTAIL.n5 104.615
R592 VTAIL.n93 VTAIL.n5 104.615
R593 VTAIL.n94 VTAIL.n93 104.615
R594 VTAIL.n302 VTAIL.n301 104.615
R595 VTAIL.n301 VTAIL.n213 104.615
R596 VTAIL.n294 VTAIL.n213 104.615
R597 VTAIL.n294 VTAIL.n293 104.615
R598 VTAIL.n293 VTAIL.n217 104.615
R599 VTAIL.n222 VTAIL.n217 104.615
R600 VTAIL.n286 VTAIL.n222 104.615
R601 VTAIL.n286 VTAIL.n285 104.615
R602 VTAIL.n285 VTAIL.n223 104.615
R603 VTAIL.n278 VTAIL.n223 104.615
R604 VTAIL.n278 VTAIL.n277 104.615
R605 VTAIL.n277 VTAIL.n227 104.615
R606 VTAIL.n270 VTAIL.n227 104.615
R607 VTAIL.n270 VTAIL.n269 104.615
R608 VTAIL.n269 VTAIL.n231 104.615
R609 VTAIL.n262 VTAIL.n231 104.615
R610 VTAIL.n262 VTAIL.n261 104.615
R611 VTAIL.n261 VTAIL.n235 104.615
R612 VTAIL.n254 VTAIL.n235 104.615
R613 VTAIL.n254 VTAIL.n253 104.615
R614 VTAIL.n253 VTAIL.n239 104.615
R615 VTAIL.n246 VTAIL.n239 104.615
R616 VTAIL.n246 VTAIL.n245 104.615
R617 VTAIL.n200 VTAIL.n199 104.615
R618 VTAIL.n199 VTAIL.n111 104.615
R619 VTAIL.n192 VTAIL.n111 104.615
R620 VTAIL.n192 VTAIL.n191 104.615
R621 VTAIL.n191 VTAIL.n115 104.615
R622 VTAIL.n120 VTAIL.n115 104.615
R623 VTAIL.n184 VTAIL.n120 104.615
R624 VTAIL.n184 VTAIL.n183 104.615
R625 VTAIL.n183 VTAIL.n121 104.615
R626 VTAIL.n176 VTAIL.n121 104.615
R627 VTAIL.n176 VTAIL.n175 104.615
R628 VTAIL.n175 VTAIL.n125 104.615
R629 VTAIL.n168 VTAIL.n125 104.615
R630 VTAIL.n168 VTAIL.n167 104.615
R631 VTAIL.n167 VTAIL.n129 104.615
R632 VTAIL.n160 VTAIL.n129 104.615
R633 VTAIL.n160 VTAIL.n159 104.615
R634 VTAIL.n159 VTAIL.n133 104.615
R635 VTAIL.n152 VTAIL.n133 104.615
R636 VTAIL.n152 VTAIL.n151 104.615
R637 VTAIL.n151 VTAIL.n137 104.615
R638 VTAIL.n144 VTAIL.n137 104.615
R639 VTAIL.n144 VTAIL.n143 104.615
R640 VTAIL.n341 VTAIL.t2 52.3082
R641 VTAIL.n35 VTAIL.t15 52.3082
R642 VTAIL.n245 VTAIL.t11 52.3082
R643 VTAIL.n143 VTAIL.t3 52.3082
R644 VTAIL.n209 VTAIL.n208 45.9428
R645 VTAIL.n207 VTAIL.n206 45.9428
R646 VTAIL.n107 VTAIL.n106 45.9428
R647 VTAIL.n105 VTAIL.n104 45.9428
R648 VTAIL.n407 VTAIL.n406 45.9426
R649 VTAIL.n1 VTAIL.n0 45.9426
R650 VTAIL.n101 VTAIL.n100 45.9426
R651 VTAIL.n103 VTAIL.n102 45.9426
R652 VTAIL.n405 VTAIL.n404 34.1247
R653 VTAIL.n99 VTAIL.n98 34.1247
R654 VTAIL.n307 VTAIL.n306 34.1247
R655 VTAIL.n205 VTAIL.n204 34.1247
R656 VTAIL.n105 VTAIL.n103 32.1772
R657 VTAIL.n405 VTAIL.n307 29.8669
R658 VTAIL.n340 VTAIL.n339 15.6677
R659 VTAIL.n34 VTAIL.n33 15.6677
R660 VTAIL.n244 VTAIL.n243 15.6677
R661 VTAIL.n142 VTAIL.n141 15.6677
R662 VTAIL.n385 VTAIL.n316 13.1884
R663 VTAIL.n79 VTAIL.n10 13.1884
R664 VTAIL.n220 VTAIL.n218 13.1884
R665 VTAIL.n118 VTAIL.n116 13.1884
R666 VTAIL.n343 VTAIL.n338 12.8005
R667 VTAIL.n386 VTAIL.n318 12.8005
R668 VTAIL.n390 VTAIL.n389 12.8005
R669 VTAIL.n37 VTAIL.n32 12.8005
R670 VTAIL.n80 VTAIL.n12 12.8005
R671 VTAIL.n84 VTAIL.n83 12.8005
R672 VTAIL.n292 VTAIL.n291 12.8005
R673 VTAIL.n288 VTAIL.n287 12.8005
R674 VTAIL.n247 VTAIL.n242 12.8005
R675 VTAIL.n190 VTAIL.n189 12.8005
R676 VTAIL.n186 VTAIL.n185 12.8005
R677 VTAIL.n145 VTAIL.n140 12.8005
R678 VTAIL.n344 VTAIL.n336 12.0247
R679 VTAIL.n381 VTAIL.n380 12.0247
R680 VTAIL.n393 VTAIL.n314 12.0247
R681 VTAIL.n38 VTAIL.n30 12.0247
R682 VTAIL.n75 VTAIL.n74 12.0247
R683 VTAIL.n87 VTAIL.n8 12.0247
R684 VTAIL.n295 VTAIL.n216 12.0247
R685 VTAIL.n284 VTAIL.n221 12.0247
R686 VTAIL.n248 VTAIL.n240 12.0247
R687 VTAIL.n193 VTAIL.n114 12.0247
R688 VTAIL.n182 VTAIL.n119 12.0247
R689 VTAIL.n146 VTAIL.n138 12.0247
R690 VTAIL.n348 VTAIL.n347 11.249
R691 VTAIL.n379 VTAIL.n320 11.249
R692 VTAIL.n394 VTAIL.n312 11.249
R693 VTAIL.n42 VTAIL.n41 11.249
R694 VTAIL.n73 VTAIL.n14 11.249
R695 VTAIL.n88 VTAIL.n6 11.249
R696 VTAIL.n296 VTAIL.n214 11.249
R697 VTAIL.n283 VTAIL.n224 11.249
R698 VTAIL.n252 VTAIL.n251 11.249
R699 VTAIL.n194 VTAIL.n112 11.249
R700 VTAIL.n181 VTAIL.n122 11.249
R701 VTAIL.n150 VTAIL.n149 11.249
R702 VTAIL.n351 VTAIL.n334 10.4732
R703 VTAIL.n376 VTAIL.n375 10.4732
R704 VTAIL.n398 VTAIL.n397 10.4732
R705 VTAIL.n45 VTAIL.n28 10.4732
R706 VTAIL.n70 VTAIL.n69 10.4732
R707 VTAIL.n92 VTAIL.n91 10.4732
R708 VTAIL.n300 VTAIL.n299 10.4732
R709 VTAIL.n280 VTAIL.n279 10.4732
R710 VTAIL.n255 VTAIL.n238 10.4732
R711 VTAIL.n198 VTAIL.n197 10.4732
R712 VTAIL.n178 VTAIL.n177 10.4732
R713 VTAIL.n153 VTAIL.n136 10.4732
R714 VTAIL.n352 VTAIL.n332 9.69747
R715 VTAIL.n372 VTAIL.n322 9.69747
R716 VTAIL.n401 VTAIL.n310 9.69747
R717 VTAIL.n46 VTAIL.n26 9.69747
R718 VTAIL.n66 VTAIL.n16 9.69747
R719 VTAIL.n95 VTAIL.n4 9.69747
R720 VTAIL.n303 VTAIL.n212 9.69747
R721 VTAIL.n276 VTAIL.n226 9.69747
R722 VTAIL.n256 VTAIL.n236 9.69747
R723 VTAIL.n201 VTAIL.n110 9.69747
R724 VTAIL.n174 VTAIL.n124 9.69747
R725 VTAIL.n154 VTAIL.n134 9.69747
R726 VTAIL.n404 VTAIL.n403 9.45567
R727 VTAIL.n98 VTAIL.n97 9.45567
R728 VTAIL.n306 VTAIL.n305 9.45567
R729 VTAIL.n204 VTAIL.n203 9.45567
R730 VTAIL.n403 VTAIL.n402 9.3005
R731 VTAIL.n310 VTAIL.n309 9.3005
R732 VTAIL.n397 VTAIL.n396 9.3005
R733 VTAIL.n395 VTAIL.n394 9.3005
R734 VTAIL.n314 VTAIL.n313 9.3005
R735 VTAIL.n389 VTAIL.n388 9.3005
R736 VTAIL.n361 VTAIL.n360 9.3005
R737 VTAIL.n330 VTAIL.n329 9.3005
R738 VTAIL.n355 VTAIL.n354 9.3005
R739 VTAIL.n353 VTAIL.n352 9.3005
R740 VTAIL.n334 VTAIL.n333 9.3005
R741 VTAIL.n347 VTAIL.n346 9.3005
R742 VTAIL.n345 VTAIL.n344 9.3005
R743 VTAIL.n338 VTAIL.n337 9.3005
R744 VTAIL.n363 VTAIL.n362 9.3005
R745 VTAIL.n326 VTAIL.n325 9.3005
R746 VTAIL.n369 VTAIL.n368 9.3005
R747 VTAIL.n371 VTAIL.n370 9.3005
R748 VTAIL.n322 VTAIL.n321 9.3005
R749 VTAIL.n377 VTAIL.n376 9.3005
R750 VTAIL.n379 VTAIL.n378 9.3005
R751 VTAIL.n380 VTAIL.n317 9.3005
R752 VTAIL.n387 VTAIL.n386 9.3005
R753 VTAIL.n97 VTAIL.n96 9.3005
R754 VTAIL.n4 VTAIL.n3 9.3005
R755 VTAIL.n91 VTAIL.n90 9.3005
R756 VTAIL.n89 VTAIL.n88 9.3005
R757 VTAIL.n8 VTAIL.n7 9.3005
R758 VTAIL.n83 VTAIL.n82 9.3005
R759 VTAIL.n55 VTAIL.n54 9.3005
R760 VTAIL.n24 VTAIL.n23 9.3005
R761 VTAIL.n49 VTAIL.n48 9.3005
R762 VTAIL.n47 VTAIL.n46 9.3005
R763 VTAIL.n28 VTAIL.n27 9.3005
R764 VTAIL.n41 VTAIL.n40 9.3005
R765 VTAIL.n39 VTAIL.n38 9.3005
R766 VTAIL.n32 VTAIL.n31 9.3005
R767 VTAIL.n57 VTAIL.n56 9.3005
R768 VTAIL.n20 VTAIL.n19 9.3005
R769 VTAIL.n63 VTAIL.n62 9.3005
R770 VTAIL.n65 VTAIL.n64 9.3005
R771 VTAIL.n16 VTAIL.n15 9.3005
R772 VTAIL.n71 VTAIL.n70 9.3005
R773 VTAIL.n73 VTAIL.n72 9.3005
R774 VTAIL.n74 VTAIL.n11 9.3005
R775 VTAIL.n81 VTAIL.n80 9.3005
R776 VTAIL.n230 VTAIL.n229 9.3005
R777 VTAIL.n273 VTAIL.n272 9.3005
R778 VTAIL.n275 VTAIL.n274 9.3005
R779 VTAIL.n226 VTAIL.n225 9.3005
R780 VTAIL.n281 VTAIL.n280 9.3005
R781 VTAIL.n283 VTAIL.n282 9.3005
R782 VTAIL.n221 VTAIL.n219 9.3005
R783 VTAIL.n289 VTAIL.n288 9.3005
R784 VTAIL.n305 VTAIL.n304 9.3005
R785 VTAIL.n212 VTAIL.n211 9.3005
R786 VTAIL.n299 VTAIL.n298 9.3005
R787 VTAIL.n297 VTAIL.n296 9.3005
R788 VTAIL.n216 VTAIL.n215 9.3005
R789 VTAIL.n291 VTAIL.n290 9.3005
R790 VTAIL.n267 VTAIL.n266 9.3005
R791 VTAIL.n265 VTAIL.n264 9.3005
R792 VTAIL.n234 VTAIL.n233 9.3005
R793 VTAIL.n259 VTAIL.n258 9.3005
R794 VTAIL.n257 VTAIL.n256 9.3005
R795 VTAIL.n238 VTAIL.n237 9.3005
R796 VTAIL.n251 VTAIL.n250 9.3005
R797 VTAIL.n249 VTAIL.n248 9.3005
R798 VTAIL.n242 VTAIL.n241 9.3005
R799 VTAIL.n128 VTAIL.n127 9.3005
R800 VTAIL.n171 VTAIL.n170 9.3005
R801 VTAIL.n173 VTAIL.n172 9.3005
R802 VTAIL.n124 VTAIL.n123 9.3005
R803 VTAIL.n179 VTAIL.n178 9.3005
R804 VTAIL.n181 VTAIL.n180 9.3005
R805 VTAIL.n119 VTAIL.n117 9.3005
R806 VTAIL.n187 VTAIL.n186 9.3005
R807 VTAIL.n203 VTAIL.n202 9.3005
R808 VTAIL.n110 VTAIL.n109 9.3005
R809 VTAIL.n197 VTAIL.n196 9.3005
R810 VTAIL.n195 VTAIL.n194 9.3005
R811 VTAIL.n114 VTAIL.n113 9.3005
R812 VTAIL.n189 VTAIL.n188 9.3005
R813 VTAIL.n165 VTAIL.n164 9.3005
R814 VTAIL.n163 VTAIL.n162 9.3005
R815 VTAIL.n132 VTAIL.n131 9.3005
R816 VTAIL.n157 VTAIL.n156 9.3005
R817 VTAIL.n155 VTAIL.n154 9.3005
R818 VTAIL.n136 VTAIL.n135 9.3005
R819 VTAIL.n149 VTAIL.n148 9.3005
R820 VTAIL.n147 VTAIL.n146 9.3005
R821 VTAIL.n140 VTAIL.n139 9.3005
R822 VTAIL.n356 VTAIL.n355 8.92171
R823 VTAIL.n371 VTAIL.n324 8.92171
R824 VTAIL.n402 VTAIL.n308 8.92171
R825 VTAIL.n50 VTAIL.n49 8.92171
R826 VTAIL.n65 VTAIL.n18 8.92171
R827 VTAIL.n96 VTAIL.n2 8.92171
R828 VTAIL.n304 VTAIL.n210 8.92171
R829 VTAIL.n275 VTAIL.n228 8.92171
R830 VTAIL.n260 VTAIL.n259 8.92171
R831 VTAIL.n202 VTAIL.n108 8.92171
R832 VTAIL.n173 VTAIL.n126 8.92171
R833 VTAIL.n158 VTAIL.n157 8.92171
R834 VTAIL.n359 VTAIL.n330 8.14595
R835 VTAIL.n368 VTAIL.n367 8.14595
R836 VTAIL.n53 VTAIL.n24 8.14595
R837 VTAIL.n62 VTAIL.n61 8.14595
R838 VTAIL.n272 VTAIL.n271 8.14595
R839 VTAIL.n263 VTAIL.n234 8.14595
R840 VTAIL.n170 VTAIL.n169 8.14595
R841 VTAIL.n161 VTAIL.n132 8.14595
R842 VTAIL.n360 VTAIL.n328 7.3702
R843 VTAIL.n364 VTAIL.n326 7.3702
R844 VTAIL.n54 VTAIL.n22 7.3702
R845 VTAIL.n58 VTAIL.n20 7.3702
R846 VTAIL.n268 VTAIL.n230 7.3702
R847 VTAIL.n264 VTAIL.n232 7.3702
R848 VTAIL.n166 VTAIL.n128 7.3702
R849 VTAIL.n162 VTAIL.n130 7.3702
R850 VTAIL.n363 VTAIL.n328 6.59444
R851 VTAIL.n364 VTAIL.n363 6.59444
R852 VTAIL.n57 VTAIL.n22 6.59444
R853 VTAIL.n58 VTAIL.n57 6.59444
R854 VTAIL.n268 VTAIL.n267 6.59444
R855 VTAIL.n267 VTAIL.n232 6.59444
R856 VTAIL.n166 VTAIL.n165 6.59444
R857 VTAIL.n165 VTAIL.n130 6.59444
R858 VTAIL.n360 VTAIL.n359 5.81868
R859 VTAIL.n367 VTAIL.n326 5.81868
R860 VTAIL.n54 VTAIL.n53 5.81868
R861 VTAIL.n61 VTAIL.n20 5.81868
R862 VTAIL.n271 VTAIL.n230 5.81868
R863 VTAIL.n264 VTAIL.n263 5.81868
R864 VTAIL.n169 VTAIL.n128 5.81868
R865 VTAIL.n162 VTAIL.n161 5.81868
R866 VTAIL.n356 VTAIL.n330 5.04292
R867 VTAIL.n368 VTAIL.n324 5.04292
R868 VTAIL.n404 VTAIL.n308 5.04292
R869 VTAIL.n50 VTAIL.n24 5.04292
R870 VTAIL.n62 VTAIL.n18 5.04292
R871 VTAIL.n98 VTAIL.n2 5.04292
R872 VTAIL.n306 VTAIL.n210 5.04292
R873 VTAIL.n272 VTAIL.n228 5.04292
R874 VTAIL.n260 VTAIL.n234 5.04292
R875 VTAIL.n204 VTAIL.n108 5.04292
R876 VTAIL.n170 VTAIL.n126 5.04292
R877 VTAIL.n158 VTAIL.n132 5.04292
R878 VTAIL.n339 VTAIL.n337 4.38563
R879 VTAIL.n33 VTAIL.n31 4.38563
R880 VTAIL.n243 VTAIL.n241 4.38563
R881 VTAIL.n141 VTAIL.n139 4.38563
R882 VTAIL.n355 VTAIL.n332 4.26717
R883 VTAIL.n372 VTAIL.n371 4.26717
R884 VTAIL.n402 VTAIL.n401 4.26717
R885 VTAIL.n49 VTAIL.n26 4.26717
R886 VTAIL.n66 VTAIL.n65 4.26717
R887 VTAIL.n96 VTAIL.n95 4.26717
R888 VTAIL.n304 VTAIL.n303 4.26717
R889 VTAIL.n276 VTAIL.n275 4.26717
R890 VTAIL.n259 VTAIL.n236 4.26717
R891 VTAIL.n202 VTAIL.n201 4.26717
R892 VTAIL.n174 VTAIL.n173 4.26717
R893 VTAIL.n157 VTAIL.n134 4.26717
R894 VTAIL.n352 VTAIL.n351 3.49141
R895 VTAIL.n375 VTAIL.n322 3.49141
R896 VTAIL.n398 VTAIL.n310 3.49141
R897 VTAIL.n46 VTAIL.n45 3.49141
R898 VTAIL.n69 VTAIL.n16 3.49141
R899 VTAIL.n92 VTAIL.n4 3.49141
R900 VTAIL.n300 VTAIL.n212 3.49141
R901 VTAIL.n279 VTAIL.n226 3.49141
R902 VTAIL.n256 VTAIL.n255 3.49141
R903 VTAIL.n198 VTAIL.n110 3.49141
R904 VTAIL.n177 VTAIL.n124 3.49141
R905 VTAIL.n154 VTAIL.n153 3.49141
R906 VTAIL.n348 VTAIL.n334 2.71565
R907 VTAIL.n376 VTAIL.n320 2.71565
R908 VTAIL.n397 VTAIL.n312 2.71565
R909 VTAIL.n42 VTAIL.n28 2.71565
R910 VTAIL.n70 VTAIL.n14 2.71565
R911 VTAIL.n91 VTAIL.n6 2.71565
R912 VTAIL.n299 VTAIL.n214 2.71565
R913 VTAIL.n280 VTAIL.n224 2.71565
R914 VTAIL.n252 VTAIL.n238 2.71565
R915 VTAIL.n197 VTAIL.n112 2.71565
R916 VTAIL.n178 VTAIL.n122 2.71565
R917 VTAIL.n150 VTAIL.n136 2.71565
R918 VTAIL.n107 VTAIL.n105 2.31084
R919 VTAIL.n205 VTAIL.n107 2.31084
R920 VTAIL.n209 VTAIL.n207 2.31084
R921 VTAIL.n307 VTAIL.n209 2.31084
R922 VTAIL.n103 VTAIL.n101 2.31084
R923 VTAIL.n101 VTAIL.n99 2.31084
R924 VTAIL.n407 VTAIL.n405 2.31084
R925 VTAIL.n347 VTAIL.n336 1.93989
R926 VTAIL.n381 VTAIL.n379 1.93989
R927 VTAIL.n394 VTAIL.n393 1.93989
R928 VTAIL.n41 VTAIL.n30 1.93989
R929 VTAIL.n75 VTAIL.n73 1.93989
R930 VTAIL.n88 VTAIL.n87 1.93989
R931 VTAIL.n296 VTAIL.n295 1.93989
R932 VTAIL.n284 VTAIL.n283 1.93989
R933 VTAIL.n251 VTAIL.n240 1.93989
R934 VTAIL.n194 VTAIL.n193 1.93989
R935 VTAIL.n182 VTAIL.n181 1.93989
R936 VTAIL.n149 VTAIL.n138 1.93989
R937 VTAIL VTAIL.n1 1.79145
R938 VTAIL.n207 VTAIL.n205 1.6255
R939 VTAIL.n99 VTAIL.n1 1.6255
R940 VTAIL.n344 VTAIL.n343 1.16414
R941 VTAIL.n380 VTAIL.n318 1.16414
R942 VTAIL.n390 VTAIL.n314 1.16414
R943 VTAIL.n38 VTAIL.n37 1.16414
R944 VTAIL.n74 VTAIL.n12 1.16414
R945 VTAIL.n84 VTAIL.n8 1.16414
R946 VTAIL.n292 VTAIL.n216 1.16414
R947 VTAIL.n287 VTAIL.n221 1.16414
R948 VTAIL.n248 VTAIL.n247 1.16414
R949 VTAIL.n190 VTAIL.n114 1.16414
R950 VTAIL.n185 VTAIL.n119 1.16414
R951 VTAIL.n146 VTAIL.n145 1.16414
R952 VTAIL.n406 VTAIL.t1 1.12422
R953 VTAIL.n406 VTAIL.t5 1.12422
R954 VTAIL.n0 VTAIL.t9 1.12422
R955 VTAIL.n0 VTAIL.t4 1.12422
R956 VTAIL.n100 VTAIL.t17 1.12422
R957 VTAIL.n100 VTAIL.t14 1.12422
R958 VTAIL.n102 VTAIL.t10 1.12422
R959 VTAIL.n102 VTAIL.t19 1.12422
R960 VTAIL.n208 VTAIL.t16 1.12422
R961 VTAIL.n208 VTAIL.t18 1.12422
R962 VTAIL.n206 VTAIL.t12 1.12422
R963 VTAIL.n206 VTAIL.t13 1.12422
R964 VTAIL.n106 VTAIL.t6 1.12422
R965 VTAIL.n106 VTAIL.t8 1.12422
R966 VTAIL.n104 VTAIL.t7 1.12422
R967 VTAIL.n104 VTAIL.t0 1.12422
R968 VTAIL VTAIL.n407 0.519897
R969 VTAIL.n340 VTAIL.n338 0.388379
R970 VTAIL.n386 VTAIL.n385 0.388379
R971 VTAIL.n389 VTAIL.n316 0.388379
R972 VTAIL.n34 VTAIL.n32 0.388379
R973 VTAIL.n80 VTAIL.n79 0.388379
R974 VTAIL.n83 VTAIL.n10 0.388379
R975 VTAIL.n291 VTAIL.n218 0.388379
R976 VTAIL.n288 VTAIL.n220 0.388379
R977 VTAIL.n244 VTAIL.n242 0.388379
R978 VTAIL.n189 VTAIL.n116 0.388379
R979 VTAIL.n186 VTAIL.n118 0.388379
R980 VTAIL.n142 VTAIL.n140 0.388379
R981 VTAIL.n345 VTAIL.n337 0.155672
R982 VTAIL.n346 VTAIL.n345 0.155672
R983 VTAIL.n346 VTAIL.n333 0.155672
R984 VTAIL.n353 VTAIL.n333 0.155672
R985 VTAIL.n354 VTAIL.n353 0.155672
R986 VTAIL.n354 VTAIL.n329 0.155672
R987 VTAIL.n361 VTAIL.n329 0.155672
R988 VTAIL.n362 VTAIL.n361 0.155672
R989 VTAIL.n362 VTAIL.n325 0.155672
R990 VTAIL.n369 VTAIL.n325 0.155672
R991 VTAIL.n370 VTAIL.n369 0.155672
R992 VTAIL.n370 VTAIL.n321 0.155672
R993 VTAIL.n377 VTAIL.n321 0.155672
R994 VTAIL.n378 VTAIL.n377 0.155672
R995 VTAIL.n378 VTAIL.n317 0.155672
R996 VTAIL.n387 VTAIL.n317 0.155672
R997 VTAIL.n388 VTAIL.n387 0.155672
R998 VTAIL.n388 VTAIL.n313 0.155672
R999 VTAIL.n395 VTAIL.n313 0.155672
R1000 VTAIL.n396 VTAIL.n395 0.155672
R1001 VTAIL.n396 VTAIL.n309 0.155672
R1002 VTAIL.n403 VTAIL.n309 0.155672
R1003 VTAIL.n39 VTAIL.n31 0.155672
R1004 VTAIL.n40 VTAIL.n39 0.155672
R1005 VTAIL.n40 VTAIL.n27 0.155672
R1006 VTAIL.n47 VTAIL.n27 0.155672
R1007 VTAIL.n48 VTAIL.n47 0.155672
R1008 VTAIL.n48 VTAIL.n23 0.155672
R1009 VTAIL.n55 VTAIL.n23 0.155672
R1010 VTAIL.n56 VTAIL.n55 0.155672
R1011 VTAIL.n56 VTAIL.n19 0.155672
R1012 VTAIL.n63 VTAIL.n19 0.155672
R1013 VTAIL.n64 VTAIL.n63 0.155672
R1014 VTAIL.n64 VTAIL.n15 0.155672
R1015 VTAIL.n71 VTAIL.n15 0.155672
R1016 VTAIL.n72 VTAIL.n71 0.155672
R1017 VTAIL.n72 VTAIL.n11 0.155672
R1018 VTAIL.n81 VTAIL.n11 0.155672
R1019 VTAIL.n82 VTAIL.n81 0.155672
R1020 VTAIL.n82 VTAIL.n7 0.155672
R1021 VTAIL.n89 VTAIL.n7 0.155672
R1022 VTAIL.n90 VTAIL.n89 0.155672
R1023 VTAIL.n90 VTAIL.n3 0.155672
R1024 VTAIL.n97 VTAIL.n3 0.155672
R1025 VTAIL.n305 VTAIL.n211 0.155672
R1026 VTAIL.n298 VTAIL.n211 0.155672
R1027 VTAIL.n298 VTAIL.n297 0.155672
R1028 VTAIL.n297 VTAIL.n215 0.155672
R1029 VTAIL.n290 VTAIL.n215 0.155672
R1030 VTAIL.n290 VTAIL.n289 0.155672
R1031 VTAIL.n289 VTAIL.n219 0.155672
R1032 VTAIL.n282 VTAIL.n219 0.155672
R1033 VTAIL.n282 VTAIL.n281 0.155672
R1034 VTAIL.n281 VTAIL.n225 0.155672
R1035 VTAIL.n274 VTAIL.n225 0.155672
R1036 VTAIL.n274 VTAIL.n273 0.155672
R1037 VTAIL.n273 VTAIL.n229 0.155672
R1038 VTAIL.n266 VTAIL.n229 0.155672
R1039 VTAIL.n266 VTAIL.n265 0.155672
R1040 VTAIL.n265 VTAIL.n233 0.155672
R1041 VTAIL.n258 VTAIL.n233 0.155672
R1042 VTAIL.n258 VTAIL.n257 0.155672
R1043 VTAIL.n257 VTAIL.n237 0.155672
R1044 VTAIL.n250 VTAIL.n237 0.155672
R1045 VTAIL.n250 VTAIL.n249 0.155672
R1046 VTAIL.n249 VTAIL.n241 0.155672
R1047 VTAIL.n203 VTAIL.n109 0.155672
R1048 VTAIL.n196 VTAIL.n109 0.155672
R1049 VTAIL.n196 VTAIL.n195 0.155672
R1050 VTAIL.n195 VTAIL.n113 0.155672
R1051 VTAIL.n188 VTAIL.n113 0.155672
R1052 VTAIL.n188 VTAIL.n187 0.155672
R1053 VTAIL.n187 VTAIL.n117 0.155672
R1054 VTAIL.n180 VTAIL.n117 0.155672
R1055 VTAIL.n180 VTAIL.n179 0.155672
R1056 VTAIL.n179 VTAIL.n123 0.155672
R1057 VTAIL.n172 VTAIL.n123 0.155672
R1058 VTAIL.n172 VTAIL.n171 0.155672
R1059 VTAIL.n171 VTAIL.n127 0.155672
R1060 VTAIL.n164 VTAIL.n127 0.155672
R1061 VTAIL.n164 VTAIL.n163 0.155672
R1062 VTAIL.n163 VTAIL.n131 0.155672
R1063 VTAIL.n156 VTAIL.n131 0.155672
R1064 VTAIL.n156 VTAIL.n155 0.155672
R1065 VTAIL.n155 VTAIL.n135 0.155672
R1066 VTAIL.n148 VTAIL.n135 0.155672
R1067 VTAIL.n148 VTAIL.n147 0.155672
R1068 VTAIL.n147 VTAIL.n139 0.155672
R1069 B.n1083 B.n1082 585
R1070 B.n417 B.n165 585
R1071 B.n416 B.n415 585
R1072 B.n414 B.n413 585
R1073 B.n412 B.n411 585
R1074 B.n410 B.n409 585
R1075 B.n408 B.n407 585
R1076 B.n406 B.n405 585
R1077 B.n404 B.n403 585
R1078 B.n402 B.n401 585
R1079 B.n400 B.n399 585
R1080 B.n398 B.n397 585
R1081 B.n396 B.n395 585
R1082 B.n394 B.n393 585
R1083 B.n392 B.n391 585
R1084 B.n390 B.n389 585
R1085 B.n388 B.n387 585
R1086 B.n386 B.n385 585
R1087 B.n384 B.n383 585
R1088 B.n382 B.n381 585
R1089 B.n380 B.n379 585
R1090 B.n378 B.n377 585
R1091 B.n376 B.n375 585
R1092 B.n374 B.n373 585
R1093 B.n372 B.n371 585
R1094 B.n370 B.n369 585
R1095 B.n368 B.n367 585
R1096 B.n366 B.n365 585
R1097 B.n364 B.n363 585
R1098 B.n362 B.n361 585
R1099 B.n360 B.n359 585
R1100 B.n358 B.n357 585
R1101 B.n356 B.n355 585
R1102 B.n354 B.n353 585
R1103 B.n352 B.n351 585
R1104 B.n350 B.n349 585
R1105 B.n348 B.n347 585
R1106 B.n346 B.n345 585
R1107 B.n344 B.n343 585
R1108 B.n342 B.n341 585
R1109 B.n340 B.n339 585
R1110 B.n338 B.n337 585
R1111 B.n336 B.n335 585
R1112 B.n334 B.n333 585
R1113 B.n332 B.n331 585
R1114 B.n330 B.n329 585
R1115 B.n328 B.n327 585
R1116 B.n326 B.n325 585
R1117 B.n324 B.n323 585
R1118 B.n322 B.n321 585
R1119 B.n320 B.n319 585
R1120 B.n318 B.n317 585
R1121 B.n316 B.n315 585
R1122 B.n314 B.n313 585
R1123 B.n312 B.n311 585
R1124 B.n310 B.n309 585
R1125 B.n308 B.n307 585
R1126 B.n306 B.n305 585
R1127 B.n304 B.n303 585
R1128 B.n302 B.n301 585
R1129 B.n300 B.n299 585
R1130 B.n298 B.n297 585
R1131 B.n296 B.n295 585
R1132 B.n294 B.n293 585
R1133 B.n292 B.n291 585
R1134 B.n290 B.n289 585
R1135 B.n288 B.n287 585
R1136 B.n286 B.n285 585
R1137 B.n284 B.n283 585
R1138 B.n282 B.n281 585
R1139 B.n280 B.n279 585
R1140 B.n278 B.n277 585
R1141 B.n276 B.n275 585
R1142 B.n274 B.n273 585
R1143 B.n272 B.n271 585
R1144 B.n270 B.n269 585
R1145 B.n268 B.n267 585
R1146 B.n266 B.n265 585
R1147 B.n264 B.n263 585
R1148 B.n262 B.n261 585
R1149 B.n260 B.n259 585
R1150 B.n258 B.n257 585
R1151 B.n256 B.n255 585
R1152 B.n254 B.n253 585
R1153 B.n252 B.n251 585
R1154 B.n250 B.n249 585
R1155 B.n248 B.n247 585
R1156 B.n246 B.n245 585
R1157 B.n244 B.n243 585
R1158 B.n242 B.n241 585
R1159 B.n240 B.n239 585
R1160 B.n238 B.n237 585
R1161 B.n236 B.n235 585
R1162 B.n234 B.n233 585
R1163 B.n232 B.n231 585
R1164 B.n230 B.n229 585
R1165 B.n228 B.n227 585
R1166 B.n226 B.n225 585
R1167 B.n224 B.n223 585
R1168 B.n222 B.n221 585
R1169 B.n220 B.n219 585
R1170 B.n218 B.n217 585
R1171 B.n216 B.n215 585
R1172 B.n214 B.n213 585
R1173 B.n212 B.n211 585
R1174 B.n210 B.n209 585
R1175 B.n208 B.n207 585
R1176 B.n206 B.n205 585
R1177 B.n204 B.n203 585
R1178 B.n202 B.n201 585
R1179 B.n200 B.n199 585
R1180 B.n198 B.n197 585
R1181 B.n196 B.n195 585
R1182 B.n194 B.n193 585
R1183 B.n192 B.n191 585
R1184 B.n190 B.n189 585
R1185 B.n188 B.n187 585
R1186 B.n186 B.n185 585
R1187 B.n184 B.n183 585
R1188 B.n182 B.n181 585
R1189 B.n180 B.n179 585
R1190 B.n178 B.n177 585
R1191 B.n176 B.n175 585
R1192 B.n174 B.n173 585
R1193 B.n103 B.n102 585
R1194 B.n1088 B.n1087 585
R1195 B.n1081 B.n166 585
R1196 B.n166 B.n100 585
R1197 B.n1080 B.n99 585
R1198 B.n1092 B.n99 585
R1199 B.n1079 B.n98 585
R1200 B.n1093 B.n98 585
R1201 B.n1078 B.n97 585
R1202 B.n1094 B.n97 585
R1203 B.n1077 B.n1076 585
R1204 B.n1076 B.n93 585
R1205 B.n1075 B.n92 585
R1206 B.n1100 B.n92 585
R1207 B.n1074 B.n91 585
R1208 B.n1101 B.n91 585
R1209 B.n1073 B.n90 585
R1210 B.n1102 B.n90 585
R1211 B.n1072 B.n1071 585
R1212 B.n1071 B.n86 585
R1213 B.n1070 B.n85 585
R1214 B.n1108 B.n85 585
R1215 B.n1069 B.n84 585
R1216 B.n1109 B.n84 585
R1217 B.n1068 B.n83 585
R1218 B.n1110 B.n83 585
R1219 B.n1067 B.n1066 585
R1220 B.n1066 B.n79 585
R1221 B.n1065 B.n78 585
R1222 B.n1116 B.n78 585
R1223 B.n1064 B.n77 585
R1224 B.n1117 B.n77 585
R1225 B.n1063 B.n76 585
R1226 B.n1118 B.n76 585
R1227 B.n1062 B.n1061 585
R1228 B.n1061 B.n72 585
R1229 B.n1060 B.n71 585
R1230 B.n1124 B.n71 585
R1231 B.n1059 B.n70 585
R1232 B.n1125 B.n70 585
R1233 B.n1058 B.n69 585
R1234 B.n1126 B.n69 585
R1235 B.n1057 B.n1056 585
R1236 B.n1056 B.n65 585
R1237 B.n1055 B.n64 585
R1238 B.n1132 B.n64 585
R1239 B.n1054 B.n63 585
R1240 B.n1133 B.n63 585
R1241 B.n1053 B.n62 585
R1242 B.n1134 B.n62 585
R1243 B.n1052 B.n1051 585
R1244 B.n1051 B.n58 585
R1245 B.n1050 B.n57 585
R1246 B.n1140 B.n57 585
R1247 B.n1049 B.n56 585
R1248 B.n1141 B.n56 585
R1249 B.n1048 B.n55 585
R1250 B.n1142 B.n55 585
R1251 B.n1047 B.n1046 585
R1252 B.n1046 B.n51 585
R1253 B.n1045 B.n50 585
R1254 B.n1148 B.n50 585
R1255 B.n1044 B.n49 585
R1256 B.n1149 B.n49 585
R1257 B.n1043 B.n48 585
R1258 B.n1150 B.n48 585
R1259 B.n1042 B.n1041 585
R1260 B.n1041 B.n44 585
R1261 B.n1040 B.n43 585
R1262 B.n1156 B.n43 585
R1263 B.n1039 B.n42 585
R1264 B.n1157 B.n42 585
R1265 B.n1038 B.n41 585
R1266 B.n1158 B.n41 585
R1267 B.n1037 B.n1036 585
R1268 B.n1036 B.n37 585
R1269 B.n1035 B.n36 585
R1270 B.n1164 B.n36 585
R1271 B.n1034 B.n35 585
R1272 B.n1165 B.n35 585
R1273 B.n1033 B.n34 585
R1274 B.n1166 B.n34 585
R1275 B.n1032 B.n1031 585
R1276 B.n1031 B.n30 585
R1277 B.n1030 B.n29 585
R1278 B.n1172 B.n29 585
R1279 B.n1029 B.n28 585
R1280 B.n1173 B.n28 585
R1281 B.n1028 B.n27 585
R1282 B.n1174 B.n27 585
R1283 B.n1027 B.n1026 585
R1284 B.n1026 B.n23 585
R1285 B.n1025 B.n22 585
R1286 B.n1180 B.n22 585
R1287 B.n1024 B.n21 585
R1288 B.n1181 B.n21 585
R1289 B.n1023 B.n20 585
R1290 B.n1182 B.n20 585
R1291 B.n1022 B.n1021 585
R1292 B.n1021 B.n16 585
R1293 B.n1020 B.n15 585
R1294 B.n1188 B.n15 585
R1295 B.n1019 B.n14 585
R1296 B.n1189 B.n14 585
R1297 B.n1018 B.n13 585
R1298 B.n1190 B.n13 585
R1299 B.n1017 B.n1016 585
R1300 B.n1016 B.n12 585
R1301 B.n1015 B.n1014 585
R1302 B.n1015 B.n8 585
R1303 B.n1013 B.n7 585
R1304 B.n1197 B.n7 585
R1305 B.n1012 B.n6 585
R1306 B.n1198 B.n6 585
R1307 B.n1011 B.n5 585
R1308 B.n1199 B.n5 585
R1309 B.n1010 B.n1009 585
R1310 B.n1009 B.n4 585
R1311 B.n1008 B.n418 585
R1312 B.n1008 B.n1007 585
R1313 B.n998 B.n419 585
R1314 B.n420 B.n419 585
R1315 B.n1000 B.n999 585
R1316 B.n1001 B.n1000 585
R1317 B.n997 B.n425 585
R1318 B.n425 B.n424 585
R1319 B.n996 B.n995 585
R1320 B.n995 B.n994 585
R1321 B.n427 B.n426 585
R1322 B.n428 B.n427 585
R1323 B.n987 B.n986 585
R1324 B.n988 B.n987 585
R1325 B.n985 B.n433 585
R1326 B.n433 B.n432 585
R1327 B.n984 B.n983 585
R1328 B.n983 B.n982 585
R1329 B.n435 B.n434 585
R1330 B.n436 B.n435 585
R1331 B.n975 B.n974 585
R1332 B.n976 B.n975 585
R1333 B.n973 B.n440 585
R1334 B.n444 B.n440 585
R1335 B.n972 B.n971 585
R1336 B.n971 B.n970 585
R1337 B.n442 B.n441 585
R1338 B.n443 B.n442 585
R1339 B.n963 B.n962 585
R1340 B.n964 B.n963 585
R1341 B.n961 B.n449 585
R1342 B.n449 B.n448 585
R1343 B.n960 B.n959 585
R1344 B.n959 B.n958 585
R1345 B.n451 B.n450 585
R1346 B.n452 B.n451 585
R1347 B.n951 B.n950 585
R1348 B.n952 B.n951 585
R1349 B.n949 B.n456 585
R1350 B.n460 B.n456 585
R1351 B.n948 B.n947 585
R1352 B.n947 B.n946 585
R1353 B.n458 B.n457 585
R1354 B.n459 B.n458 585
R1355 B.n939 B.n938 585
R1356 B.n940 B.n939 585
R1357 B.n937 B.n465 585
R1358 B.n465 B.n464 585
R1359 B.n936 B.n935 585
R1360 B.n935 B.n934 585
R1361 B.n467 B.n466 585
R1362 B.n468 B.n467 585
R1363 B.n927 B.n926 585
R1364 B.n928 B.n927 585
R1365 B.n925 B.n472 585
R1366 B.n476 B.n472 585
R1367 B.n924 B.n923 585
R1368 B.n923 B.n922 585
R1369 B.n474 B.n473 585
R1370 B.n475 B.n474 585
R1371 B.n915 B.n914 585
R1372 B.n916 B.n915 585
R1373 B.n913 B.n481 585
R1374 B.n481 B.n480 585
R1375 B.n912 B.n911 585
R1376 B.n911 B.n910 585
R1377 B.n483 B.n482 585
R1378 B.n484 B.n483 585
R1379 B.n903 B.n902 585
R1380 B.n904 B.n903 585
R1381 B.n901 B.n488 585
R1382 B.n492 B.n488 585
R1383 B.n900 B.n899 585
R1384 B.n899 B.n898 585
R1385 B.n490 B.n489 585
R1386 B.n491 B.n490 585
R1387 B.n891 B.n890 585
R1388 B.n892 B.n891 585
R1389 B.n889 B.n497 585
R1390 B.n497 B.n496 585
R1391 B.n888 B.n887 585
R1392 B.n887 B.n886 585
R1393 B.n499 B.n498 585
R1394 B.n500 B.n499 585
R1395 B.n879 B.n878 585
R1396 B.n880 B.n879 585
R1397 B.n877 B.n505 585
R1398 B.n505 B.n504 585
R1399 B.n876 B.n875 585
R1400 B.n875 B.n874 585
R1401 B.n507 B.n506 585
R1402 B.n508 B.n507 585
R1403 B.n867 B.n866 585
R1404 B.n868 B.n867 585
R1405 B.n865 B.n513 585
R1406 B.n513 B.n512 585
R1407 B.n864 B.n863 585
R1408 B.n863 B.n862 585
R1409 B.n515 B.n514 585
R1410 B.n516 B.n515 585
R1411 B.n855 B.n854 585
R1412 B.n856 B.n855 585
R1413 B.n853 B.n521 585
R1414 B.n521 B.n520 585
R1415 B.n852 B.n851 585
R1416 B.n851 B.n850 585
R1417 B.n523 B.n522 585
R1418 B.n524 B.n523 585
R1419 B.n846 B.n845 585
R1420 B.n527 B.n526 585
R1421 B.n842 B.n841 585
R1422 B.n843 B.n842 585
R1423 B.n840 B.n590 585
R1424 B.n839 B.n838 585
R1425 B.n837 B.n836 585
R1426 B.n835 B.n834 585
R1427 B.n833 B.n832 585
R1428 B.n831 B.n830 585
R1429 B.n829 B.n828 585
R1430 B.n827 B.n826 585
R1431 B.n825 B.n824 585
R1432 B.n823 B.n822 585
R1433 B.n821 B.n820 585
R1434 B.n819 B.n818 585
R1435 B.n817 B.n816 585
R1436 B.n815 B.n814 585
R1437 B.n813 B.n812 585
R1438 B.n811 B.n810 585
R1439 B.n809 B.n808 585
R1440 B.n807 B.n806 585
R1441 B.n805 B.n804 585
R1442 B.n803 B.n802 585
R1443 B.n801 B.n800 585
R1444 B.n799 B.n798 585
R1445 B.n797 B.n796 585
R1446 B.n795 B.n794 585
R1447 B.n793 B.n792 585
R1448 B.n791 B.n790 585
R1449 B.n789 B.n788 585
R1450 B.n787 B.n786 585
R1451 B.n785 B.n784 585
R1452 B.n783 B.n782 585
R1453 B.n781 B.n780 585
R1454 B.n779 B.n778 585
R1455 B.n777 B.n776 585
R1456 B.n775 B.n774 585
R1457 B.n773 B.n772 585
R1458 B.n771 B.n770 585
R1459 B.n769 B.n768 585
R1460 B.n767 B.n766 585
R1461 B.n765 B.n764 585
R1462 B.n763 B.n762 585
R1463 B.n761 B.n760 585
R1464 B.n759 B.n758 585
R1465 B.n757 B.n756 585
R1466 B.n755 B.n754 585
R1467 B.n753 B.n752 585
R1468 B.n751 B.n750 585
R1469 B.n749 B.n748 585
R1470 B.n747 B.n746 585
R1471 B.n745 B.n744 585
R1472 B.n743 B.n742 585
R1473 B.n741 B.n740 585
R1474 B.n739 B.n738 585
R1475 B.n737 B.n736 585
R1476 B.n735 B.n734 585
R1477 B.n733 B.n732 585
R1478 B.n730 B.n729 585
R1479 B.n728 B.n727 585
R1480 B.n726 B.n725 585
R1481 B.n724 B.n723 585
R1482 B.n722 B.n721 585
R1483 B.n720 B.n719 585
R1484 B.n718 B.n717 585
R1485 B.n716 B.n715 585
R1486 B.n714 B.n713 585
R1487 B.n712 B.n711 585
R1488 B.n709 B.n708 585
R1489 B.n707 B.n706 585
R1490 B.n705 B.n704 585
R1491 B.n703 B.n702 585
R1492 B.n701 B.n700 585
R1493 B.n699 B.n698 585
R1494 B.n697 B.n696 585
R1495 B.n695 B.n694 585
R1496 B.n693 B.n692 585
R1497 B.n691 B.n690 585
R1498 B.n689 B.n688 585
R1499 B.n687 B.n686 585
R1500 B.n685 B.n684 585
R1501 B.n683 B.n682 585
R1502 B.n681 B.n680 585
R1503 B.n679 B.n678 585
R1504 B.n677 B.n676 585
R1505 B.n675 B.n674 585
R1506 B.n673 B.n672 585
R1507 B.n671 B.n670 585
R1508 B.n669 B.n668 585
R1509 B.n667 B.n666 585
R1510 B.n665 B.n664 585
R1511 B.n663 B.n662 585
R1512 B.n661 B.n660 585
R1513 B.n659 B.n658 585
R1514 B.n657 B.n656 585
R1515 B.n655 B.n654 585
R1516 B.n653 B.n652 585
R1517 B.n651 B.n650 585
R1518 B.n649 B.n648 585
R1519 B.n647 B.n646 585
R1520 B.n645 B.n644 585
R1521 B.n643 B.n642 585
R1522 B.n641 B.n640 585
R1523 B.n639 B.n638 585
R1524 B.n637 B.n636 585
R1525 B.n635 B.n634 585
R1526 B.n633 B.n632 585
R1527 B.n631 B.n630 585
R1528 B.n629 B.n628 585
R1529 B.n627 B.n626 585
R1530 B.n625 B.n624 585
R1531 B.n623 B.n622 585
R1532 B.n621 B.n620 585
R1533 B.n619 B.n618 585
R1534 B.n617 B.n616 585
R1535 B.n615 B.n614 585
R1536 B.n613 B.n612 585
R1537 B.n611 B.n610 585
R1538 B.n609 B.n608 585
R1539 B.n607 B.n606 585
R1540 B.n605 B.n604 585
R1541 B.n603 B.n602 585
R1542 B.n601 B.n600 585
R1543 B.n599 B.n598 585
R1544 B.n597 B.n596 585
R1545 B.n595 B.n589 585
R1546 B.n843 B.n589 585
R1547 B.n847 B.n525 585
R1548 B.n525 B.n524 585
R1549 B.n849 B.n848 585
R1550 B.n850 B.n849 585
R1551 B.n519 B.n518 585
R1552 B.n520 B.n519 585
R1553 B.n858 B.n857 585
R1554 B.n857 B.n856 585
R1555 B.n859 B.n517 585
R1556 B.n517 B.n516 585
R1557 B.n861 B.n860 585
R1558 B.n862 B.n861 585
R1559 B.n511 B.n510 585
R1560 B.n512 B.n511 585
R1561 B.n870 B.n869 585
R1562 B.n869 B.n868 585
R1563 B.n871 B.n509 585
R1564 B.n509 B.n508 585
R1565 B.n873 B.n872 585
R1566 B.n874 B.n873 585
R1567 B.n503 B.n502 585
R1568 B.n504 B.n503 585
R1569 B.n882 B.n881 585
R1570 B.n881 B.n880 585
R1571 B.n883 B.n501 585
R1572 B.n501 B.n500 585
R1573 B.n885 B.n884 585
R1574 B.n886 B.n885 585
R1575 B.n495 B.n494 585
R1576 B.n496 B.n495 585
R1577 B.n894 B.n893 585
R1578 B.n893 B.n892 585
R1579 B.n895 B.n493 585
R1580 B.n493 B.n491 585
R1581 B.n897 B.n896 585
R1582 B.n898 B.n897 585
R1583 B.n487 B.n486 585
R1584 B.n492 B.n487 585
R1585 B.n906 B.n905 585
R1586 B.n905 B.n904 585
R1587 B.n907 B.n485 585
R1588 B.n485 B.n484 585
R1589 B.n909 B.n908 585
R1590 B.n910 B.n909 585
R1591 B.n479 B.n478 585
R1592 B.n480 B.n479 585
R1593 B.n918 B.n917 585
R1594 B.n917 B.n916 585
R1595 B.n919 B.n477 585
R1596 B.n477 B.n475 585
R1597 B.n921 B.n920 585
R1598 B.n922 B.n921 585
R1599 B.n471 B.n470 585
R1600 B.n476 B.n471 585
R1601 B.n930 B.n929 585
R1602 B.n929 B.n928 585
R1603 B.n931 B.n469 585
R1604 B.n469 B.n468 585
R1605 B.n933 B.n932 585
R1606 B.n934 B.n933 585
R1607 B.n463 B.n462 585
R1608 B.n464 B.n463 585
R1609 B.n942 B.n941 585
R1610 B.n941 B.n940 585
R1611 B.n943 B.n461 585
R1612 B.n461 B.n459 585
R1613 B.n945 B.n944 585
R1614 B.n946 B.n945 585
R1615 B.n455 B.n454 585
R1616 B.n460 B.n455 585
R1617 B.n954 B.n953 585
R1618 B.n953 B.n952 585
R1619 B.n955 B.n453 585
R1620 B.n453 B.n452 585
R1621 B.n957 B.n956 585
R1622 B.n958 B.n957 585
R1623 B.n447 B.n446 585
R1624 B.n448 B.n447 585
R1625 B.n966 B.n965 585
R1626 B.n965 B.n964 585
R1627 B.n967 B.n445 585
R1628 B.n445 B.n443 585
R1629 B.n969 B.n968 585
R1630 B.n970 B.n969 585
R1631 B.n439 B.n438 585
R1632 B.n444 B.n439 585
R1633 B.n978 B.n977 585
R1634 B.n977 B.n976 585
R1635 B.n979 B.n437 585
R1636 B.n437 B.n436 585
R1637 B.n981 B.n980 585
R1638 B.n982 B.n981 585
R1639 B.n431 B.n430 585
R1640 B.n432 B.n431 585
R1641 B.n990 B.n989 585
R1642 B.n989 B.n988 585
R1643 B.n991 B.n429 585
R1644 B.n429 B.n428 585
R1645 B.n993 B.n992 585
R1646 B.n994 B.n993 585
R1647 B.n423 B.n422 585
R1648 B.n424 B.n423 585
R1649 B.n1003 B.n1002 585
R1650 B.n1002 B.n1001 585
R1651 B.n1004 B.n421 585
R1652 B.n421 B.n420 585
R1653 B.n1006 B.n1005 585
R1654 B.n1007 B.n1006 585
R1655 B.n3 B.n0 585
R1656 B.n4 B.n3 585
R1657 B.n1196 B.n1 585
R1658 B.n1197 B.n1196 585
R1659 B.n1195 B.n1194 585
R1660 B.n1195 B.n8 585
R1661 B.n1193 B.n9 585
R1662 B.n12 B.n9 585
R1663 B.n1192 B.n1191 585
R1664 B.n1191 B.n1190 585
R1665 B.n11 B.n10 585
R1666 B.n1189 B.n11 585
R1667 B.n1187 B.n1186 585
R1668 B.n1188 B.n1187 585
R1669 B.n1185 B.n17 585
R1670 B.n17 B.n16 585
R1671 B.n1184 B.n1183 585
R1672 B.n1183 B.n1182 585
R1673 B.n19 B.n18 585
R1674 B.n1181 B.n19 585
R1675 B.n1179 B.n1178 585
R1676 B.n1180 B.n1179 585
R1677 B.n1177 B.n24 585
R1678 B.n24 B.n23 585
R1679 B.n1176 B.n1175 585
R1680 B.n1175 B.n1174 585
R1681 B.n26 B.n25 585
R1682 B.n1173 B.n26 585
R1683 B.n1171 B.n1170 585
R1684 B.n1172 B.n1171 585
R1685 B.n1169 B.n31 585
R1686 B.n31 B.n30 585
R1687 B.n1168 B.n1167 585
R1688 B.n1167 B.n1166 585
R1689 B.n33 B.n32 585
R1690 B.n1165 B.n33 585
R1691 B.n1163 B.n1162 585
R1692 B.n1164 B.n1163 585
R1693 B.n1161 B.n38 585
R1694 B.n38 B.n37 585
R1695 B.n1160 B.n1159 585
R1696 B.n1159 B.n1158 585
R1697 B.n40 B.n39 585
R1698 B.n1157 B.n40 585
R1699 B.n1155 B.n1154 585
R1700 B.n1156 B.n1155 585
R1701 B.n1153 B.n45 585
R1702 B.n45 B.n44 585
R1703 B.n1152 B.n1151 585
R1704 B.n1151 B.n1150 585
R1705 B.n47 B.n46 585
R1706 B.n1149 B.n47 585
R1707 B.n1147 B.n1146 585
R1708 B.n1148 B.n1147 585
R1709 B.n1145 B.n52 585
R1710 B.n52 B.n51 585
R1711 B.n1144 B.n1143 585
R1712 B.n1143 B.n1142 585
R1713 B.n54 B.n53 585
R1714 B.n1141 B.n54 585
R1715 B.n1139 B.n1138 585
R1716 B.n1140 B.n1139 585
R1717 B.n1137 B.n59 585
R1718 B.n59 B.n58 585
R1719 B.n1136 B.n1135 585
R1720 B.n1135 B.n1134 585
R1721 B.n61 B.n60 585
R1722 B.n1133 B.n61 585
R1723 B.n1131 B.n1130 585
R1724 B.n1132 B.n1131 585
R1725 B.n1129 B.n66 585
R1726 B.n66 B.n65 585
R1727 B.n1128 B.n1127 585
R1728 B.n1127 B.n1126 585
R1729 B.n68 B.n67 585
R1730 B.n1125 B.n68 585
R1731 B.n1123 B.n1122 585
R1732 B.n1124 B.n1123 585
R1733 B.n1121 B.n73 585
R1734 B.n73 B.n72 585
R1735 B.n1120 B.n1119 585
R1736 B.n1119 B.n1118 585
R1737 B.n75 B.n74 585
R1738 B.n1117 B.n75 585
R1739 B.n1115 B.n1114 585
R1740 B.n1116 B.n1115 585
R1741 B.n1113 B.n80 585
R1742 B.n80 B.n79 585
R1743 B.n1112 B.n1111 585
R1744 B.n1111 B.n1110 585
R1745 B.n82 B.n81 585
R1746 B.n1109 B.n82 585
R1747 B.n1107 B.n1106 585
R1748 B.n1108 B.n1107 585
R1749 B.n1105 B.n87 585
R1750 B.n87 B.n86 585
R1751 B.n1104 B.n1103 585
R1752 B.n1103 B.n1102 585
R1753 B.n89 B.n88 585
R1754 B.n1101 B.n89 585
R1755 B.n1099 B.n1098 585
R1756 B.n1100 B.n1099 585
R1757 B.n1097 B.n94 585
R1758 B.n94 B.n93 585
R1759 B.n1096 B.n1095 585
R1760 B.n1095 B.n1094 585
R1761 B.n96 B.n95 585
R1762 B.n1093 B.n96 585
R1763 B.n1091 B.n1090 585
R1764 B.n1092 B.n1091 585
R1765 B.n1089 B.n101 585
R1766 B.n101 B.n100 585
R1767 B.n1200 B.n1199 585
R1768 B.n1198 B.n2 585
R1769 B.n1087 B.n101 473.281
R1770 B.n1083 B.n166 473.281
R1771 B.n589 B.n523 473.281
R1772 B.n845 B.n525 473.281
R1773 B.n167 B.t16 431.175
R1774 B.n593 B.t13 431.175
R1775 B.n170 B.t19 431.175
R1776 B.n591 B.t23 431.175
R1777 B.n170 B.t18 388.334
R1778 B.n167 B.t14 388.334
R1779 B.n593 B.t10 388.334
R1780 B.n591 B.t21 388.334
R1781 B.n168 B.t17 379.199
R1782 B.n594 B.t12 379.199
R1783 B.n171 B.t20 379.199
R1784 B.n592 B.t22 379.199
R1785 B.n1085 B.n1084 256.663
R1786 B.n1085 B.n164 256.663
R1787 B.n1085 B.n163 256.663
R1788 B.n1085 B.n162 256.663
R1789 B.n1085 B.n161 256.663
R1790 B.n1085 B.n160 256.663
R1791 B.n1085 B.n159 256.663
R1792 B.n1085 B.n158 256.663
R1793 B.n1085 B.n157 256.663
R1794 B.n1085 B.n156 256.663
R1795 B.n1085 B.n155 256.663
R1796 B.n1085 B.n154 256.663
R1797 B.n1085 B.n153 256.663
R1798 B.n1085 B.n152 256.663
R1799 B.n1085 B.n151 256.663
R1800 B.n1085 B.n150 256.663
R1801 B.n1085 B.n149 256.663
R1802 B.n1085 B.n148 256.663
R1803 B.n1085 B.n147 256.663
R1804 B.n1085 B.n146 256.663
R1805 B.n1085 B.n145 256.663
R1806 B.n1085 B.n144 256.663
R1807 B.n1085 B.n143 256.663
R1808 B.n1085 B.n142 256.663
R1809 B.n1085 B.n141 256.663
R1810 B.n1085 B.n140 256.663
R1811 B.n1085 B.n139 256.663
R1812 B.n1085 B.n138 256.663
R1813 B.n1085 B.n137 256.663
R1814 B.n1085 B.n136 256.663
R1815 B.n1085 B.n135 256.663
R1816 B.n1085 B.n134 256.663
R1817 B.n1085 B.n133 256.663
R1818 B.n1085 B.n132 256.663
R1819 B.n1085 B.n131 256.663
R1820 B.n1085 B.n130 256.663
R1821 B.n1085 B.n129 256.663
R1822 B.n1085 B.n128 256.663
R1823 B.n1085 B.n127 256.663
R1824 B.n1085 B.n126 256.663
R1825 B.n1085 B.n125 256.663
R1826 B.n1085 B.n124 256.663
R1827 B.n1085 B.n123 256.663
R1828 B.n1085 B.n122 256.663
R1829 B.n1085 B.n121 256.663
R1830 B.n1085 B.n120 256.663
R1831 B.n1085 B.n119 256.663
R1832 B.n1085 B.n118 256.663
R1833 B.n1085 B.n117 256.663
R1834 B.n1085 B.n116 256.663
R1835 B.n1085 B.n115 256.663
R1836 B.n1085 B.n114 256.663
R1837 B.n1085 B.n113 256.663
R1838 B.n1085 B.n112 256.663
R1839 B.n1085 B.n111 256.663
R1840 B.n1085 B.n110 256.663
R1841 B.n1085 B.n109 256.663
R1842 B.n1085 B.n108 256.663
R1843 B.n1085 B.n107 256.663
R1844 B.n1085 B.n106 256.663
R1845 B.n1085 B.n105 256.663
R1846 B.n1085 B.n104 256.663
R1847 B.n1086 B.n1085 256.663
R1848 B.n844 B.n843 256.663
R1849 B.n843 B.n528 256.663
R1850 B.n843 B.n529 256.663
R1851 B.n843 B.n530 256.663
R1852 B.n843 B.n531 256.663
R1853 B.n843 B.n532 256.663
R1854 B.n843 B.n533 256.663
R1855 B.n843 B.n534 256.663
R1856 B.n843 B.n535 256.663
R1857 B.n843 B.n536 256.663
R1858 B.n843 B.n537 256.663
R1859 B.n843 B.n538 256.663
R1860 B.n843 B.n539 256.663
R1861 B.n843 B.n540 256.663
R1862 B.n843 B.n541 256.663
R1863 B.n843 B.n542 256.663
R1864 B.n843 B.n543 256.663
R1865 B.n843 B.n544 256.663
R1866 B.n843 B.n545 256.663
R1867 B.n843 B.n546 256.663
R1868 B.n843 B.n547 256.663
R1869 B.n843 B.n548 256.663
R1870 B.n843 B.n549 256.663
R1871 B.n843 B.n550 256.663
R1872 B.n843 B.n551 256.663
R1873 B.n843 B.n552 256.663
R1874 B.n843 B.n553 256.663
R1875 B.n843 B.n554 256.663
R1876 B.n843 B.n555 256.663
R1877 B.n843 B.n556 256.663
R1878 B.n843 B.n557 256.663
R1879 B.n843 B.n558 256.663
R1880 B.n843 B.n559 256.663
R1881 B.n843 B.n560 256.663
R1882 B.n843 B.n561 256.663
R1883 B.n843 B.n562 256.663
R1884 B.n843 B.n563 256.663
R1885 B.n843 B.n564 256.663
R1886 B.n843 B.n565 256.663
R1887 B.n843 B.n566 256.663
R1888 B.n843 B.n567 256.663
R1889 B.n843 B.n568 256.663
R1890 B.n843 B.n569 256.663
R1891 B.n843 B.n570 256.663
R1892 B.n843 B.n571 256.663
R1893 B.n843 B.n572 256.663
R1894 B.n843 B.n573 256.663
R1895 B.n843 B.n574 256.663
R1896 B.n843 B.n575 256.663
R1897 B.n843 B.n576 256.663
R1898 B.n843 B.n577 256.663
R1899 B.n843 B.n578 256.663
R1900 B.n843 B.n579 256.663
R1901 B.n843 B.n580 256.663
R1902 B.n843 B.n581 256.663
R1903 B.n843 B.n582 256.663
R1904 B.n843 B.n583 256.663
R1905 B.n843 B.n584 256.663
R1906 B.n843 B.n585 256.663
R1907 B.n843 B.n586 256.663
R1908 B.n843 B.n587 256.663
R1909 B.n843 B.n588 256.663
R1910 B.n1202 B.n1201 256.663
R1911 B.n173 B.n103 163.367
R1912 B.n177 B.n176 163.367
R1913 B.n181 B.n180 163.367
R1914 B.n185 B.n184 163.367
R1915 B.n189 B.n188 163.367
R1916 B.n193 B.n192 163.367
R1917 B.n197 B.n196 163.367
R1918 B.n201 B.n200 163.367
R1919 B.n205 B.n204 163.367
R1920 B.n209 B.n208 163.367
R1921 B.n213 B.n212 163.367
R1922 B.n217 B.n216 163.367
R1923 B.n221 B.n220 163.367
R1924 B.n225 B.n224 163.367
R1925 B.n229 B.n228 163.367
R1926 B.n233 B.n232 163.367
R1927 B.n237 B.n236 163.367
R1928 B.n241 B.n240 163.367
R1929 B.n245 B.n244 163.367
R1930 B.n249 B.n248 163.367
R1931 B.n253 B.n252 163.367
R1932 B.n257 B.n256 163.367
R1933 B.n261 B.n260 163.367
R1934 B.n265 B.n264 163.367
R1935 B.n269 B.n268 163.367
R1936 B.n273 B.n272 163.367
R1937 B.n277 B.n276 163.367
R1938 B.n281 B.n280 163.367
R1939 B.n285 B.n284 163.367
R1940 B.n289 B.n288 163.367
R1941 B.n293 B.n292 163.367
R1942 B.n297 B.n296 163.367
R1943 B.n301 B.n300 163.367
R1944 B.n305 B.n304 163.367
R1945 B.n309 B.n308 163.367
R1946 B.n313 B.n312 163.367
R1947 B.n317 B.n316 163.367
R1948 B.n321 B.n320 163.367
R1949 B.n325 B.n324 163.367
R1950 B.n329 B.n328 163.367
R1951 B.n333 B.n332 163.367
R1952 B.n337 B.n336 163.367
R1953 B.n341 B.n340 163.367
R1954 B.n345 B.n344 163.367
R1955 B.n349 B.n348 163.367
R1956 B.n353 B.n352 163.367
R1957 B.n357 B.n356 163.367
R1958 B.n361 B.n360 163.367
R1959 B.n365 B.n364 163.367
R1960 B.n369 B.n368 163.367
R1961 B.n373 B.n372 163.367
R1962 B.n377 B.n376 163.367
R1963 B.n381 B.n380 163.367
R1964 B.n385 B.n384 163.367
R1965 B.n389 B.n388 163.367
R1966 B.n393 B.n392 163.367
R1967 B.n397 B.n396 163.367
R1968 B.n401 B.n400 163.367
R1969 B.n405 B.n404 163.367
R1970 B.n409 B.n408 163.367
R1971 B.n413 B.n412 163.367
R1972 B.n415 B.n165 163.367
R1973 B.n851 B.n523 163.367
R1974 B.n851 B.n521 163.367
R1975 B.n855 B.n521 163.367
R1976 B.n855 B.n515 163.367
R1977 B.n863 B.n515 163.367
R1978 B.n863 B.n513 163.367
R1979 B.n867 B.n513 163.367
R1980 B.n867 B.n507 163.367
R1981 B.n875 B.n507 163.367
R1982 B.n875 B.n505 163.367
R1983 B.n879 B.n505 163.367
R1984 B.n879 B.n499 163.367
R1985 B.n887 B.n499 163.367
R1986 B.n887 B.n497 163.367
R1987 B.n891 B.n497 163.367
R1988 B.n891 B.n490 163.367
R1989 B.n899 B.n490 163.367
R1990 B.n899 B.n488 163.367
R1991 B.n903 B.n488 163.367
R1992 B.n903 B.n483 163.367
R1993 B.n911 B.n483 163.367
R1994 B.n911 B.n481 163.367
R1995 B.n915 B.n481 163.367
R1996 B.n915 B.n474 163.367
R1997 B.n923 B.n474 163.367
R1998 B.n923 B.n472 163.367
R1999 B.n927 B.n472 163.367
R2000 B.n927 B.n467 163.367
R2001 B.n935 B.n467 163.367
R2002 B.n935 B.n465 163.367
R2003 B.n939 B.n465 163.367
R2004 B.n939 B.n458 163.367
R2005 B.n947 B.n458 163.367
R2006 B.n947 B.n456 163.367
R2007 B.n951 B.n456 163.367
R2008 B.n951 B.n451 163.367
R2009 B.n959 B.n451 163.367
R2010 B.n959 B.n449 163.367
R2011 B.n963 B.n449 163.367
R2012 B.n963 B.n442 163.367
R2013 B.n971 B.n442 163.367
R2014 B.n971 B.n440 163.367
R2015 B.n975 B.n440 163.367
R2016 B.n975 B.n435 163.367
R2017 B.n983 B.n435 163.367
R2018 B.n983 B.n433 163.367
R2019 B.n987 B.n433 163.367
R2020 B.n987 B.n427 163.367
R2021 B.n995 B.n427 163.367
R2022 B.n995 B.n425 163.367
R2023 B.n1000 B.n425 163.367
R2024 B.n1000 B.n419 163.367
R2025 B.n1008 B.n419 163.367
R2026 B.n1009 B.n1008 163.367
R2027 B.n1009 B.n5 163.367
R2028 B.n6 B.n5 163.367
R2029 B.n7 B.n6 163.367
R2030 B.n1015 B.n7 163.367
R2031 B.n1016 B.n1015 163.367
R2032 B.n1016 B.n13 163.367
R2033 B.n14 B.n13 163.367
R2034 B.n15 B.n14 163.367
R2035 B.n1021 B.n15 163.367
R2036 B.n1021 B.n20 163.367
R2037 B.n21 B.n20 163.367
R2038 B.n22 B.n21 163.367
R2039 B.n1026 B.n22 163.367
R2040 B.n1026 B.n27 163.367
R2041 B.n28 B.n27 163.367
R2042 B.n29 B.n28 163.367
R2043 B.n1031 B.n29 163.367
R2044 B.n1031 B.n34 163.367
R2045 B.n35 B.n34 163.367
R2046 B.n36 B.n35 163.367
R2047 B.n1036 B.n36 163.367
R2048 B.n1036 B.n41 163.367
R2049 B.n42 B.n41 163.367
R2050 B.n43 B.n42 163.367
R2051 B.n1041 B.n43 163.367
R2052 B.n1041 B.n48 163.367
R2053 B.n49 B.n48 163.367
R2054 B.n50 B.n49 163.367
R2055 B.n1046 B.n50 163.367
R2056 B.n1046 B.n55 163.367
R2057 B.n56 B.n55 163.367
R2058 B.n57 B.n56 163.367
R2059 B.n1051 B.n57 163.367
R2060 B.n1051 B.n62 163.367
R2061 B.n63 B.n62 163.367
R2062 B.n64 B.n63 163.367
R2063 B.n1056 B.n64 163.367
R2064 B.n1056 B.n69 163.367
R2065 B.n70 B.n69 163.367
R2066 B.n71 B.n70 163.367
R2067 B.n1061 B.n71 163.367
R2068 B.n1061 B.n76 163.367
R2069 B.n77 B.n76 163.367
R2070 B.n78 B.n77 163.367
R2071 B.n1066 B.n78 163.367
R2072 B.n1066 B.n83 163.367
R2073 B.n84 B.n83 163.367
R2074 B.n85 B.n84 163.367
R2075 B.n1071 B.n85 163.367
R2076 B.n1071 B.n90 163.367
R2077 B.n91 B.n90 163.367
R2078 B.n92 B.n91 163.367
R2079 B.n1076 B.n92 163.367
R2080 B.n1076 B.n97 163.367
R2081 B.n98 B.n97 163.367
R2082 B.n99 B.n98 163.367
R2083 B.n166 B.n99 163.367
R2084 B.n842 B.n527 163.367
R2085 B.n842 B.n590 163.367
R2086 B.n838 B.n837 163.367
R2087 B.n834 B.n833 163.367
R2088 B.n830 B.n829 163.367
R2089 B.n826 B.n825 163.367
R2090 B.n822 B.n821 163.367
R2091 B.n818 B.n817 163.367
R2092 B.n814 B.n813 163.367
R2093 B.n810 B.n809 163.367
R2094 B.n806 B.n805 163.367
R2095 B.n802 B.n801 163.367
R2096 B.n798 B.n797 163.367
R2097 B.n794 B.n793 163.367
R2098 B.n790 B.n789 163.367
R2099 B.n786 B.n785 163.367
R2100 B.n782 B.n781 163.367
R2101 B.n778 B.n777 163.367
R2102 B.n774 B.n773 163.367
R2103 B.n770 B.n769 163.367
R2104 B.n766 B.n765 163.367
R2105 B.n762 B.n761 163.367
R2106 B.n758 B.n757 163.367
R2107 B.n754 B.n753 163.367
R2108 B.n750 B.n749 163.367
R2109 B.n746 B.n745 163.367
R2110 B.n742 B.n741 163.367
R2111 B.n738 B.n737 163.367
R2112 B.n734 B.n733 163.367
R2113 B.n729 B.n728 163.367
R2114 B.n725 B.n724 163.367
R2115 B.n721 B.n720 163.367
R2116 B.n717 B.n716 163.367
R2117 B.n713 B.n712 163.367
R2118 B.n708 B.n707 163.367
R2119 B.n704 B.n703 163.367
R2120 B.n700 B.n699 163.367
R2121 B.n696 B.n695 163.367
R2122 B.n692 B.n691 163.367
R2123 B.n688 B.n687 163.367
R2124 B.n684 B.n683 163.367
R2125 B.n680 B.n679 163.367
R2126 B.n676 B.n675 163.367
R2127 B.n672 B.n671 163.367
R2128 B.n668 B.n667 163.367
R2129 B.n664 B.n663 163.367
R2130 B.n660 B.n659 163.367
R2131 B.n656 B.n655 163.367
R2132 B.n652 B.n651 163.367
R2133 B.n648 B.n647 163.367
R2134 B.n644 B.n643 163.367
R2135 B.n640 B.n639 163.367
R2136 B.n636 B.n635 163.367
R2137 B.n632 B.n631 163.367
R2138 B.n628 B.n627 163.367
R2139 B.n624 B.n623 163.367
R2140 B.n620 B.n619 163.367
R2141 B.n616 B.n615 163.367
R2142 B.n612 B.n611 163.367
R2143 B.n608 B.n607 163.367
R2144 B.n604 B.n603 163.367
R2145 B.n600 B.n599 163.367
R2146 B.n596 B.n589 163.367
R2147 B.n849 B.n525 163.367
R2148 B.n849 B.n519 163.367
R2149 B.n857 B.n519 163.367
R2150 B.n857 B.n517 163.367
R2151 B.n861 B.n517 163.367
R2152 B.n861 B.n511 163.367
R2153 B.n869 B.n511 163.367
R2154 B.n869 B.n509 163.367
R2155 B.n873 B.n509 163.367
R2156 B.n873 B.n503 163.367
R2157 B.n881 B.n503 163.367
R2158 B.n881 B.n501 163.367
R2159 B.n885 B.n501 163.367
R2160 B.n885 B.n495 163.367
R2161 B.n893 B.n495 163.367
R2162 B.n893 B.n493 163.367
R2163 B.n897 B.n493 163.367
R2164 B.n897 B.n487 163.367
R2165 B.n905 B.n487 163.367
R2166 B.n905 B.n485 163.367
R2167 B.n909 B.n485 163.367
R2168 B.n909 B.n479 163.367
R2169 B.n917 B.n479 163.367
R2170 B.n917 B.n477 163.367
R2171 B.n921 B.n477 163.367
R2172 B.n921 B.n471 163.367
R2173 B.n929 B.n471 163.367
R2174 B.n929 B.n469 163.367
R2175 B.n933 B.n469 163.367
R2176 B.n933 B.n463 163.367
R2177 B.n941 B.n463 163.367
R2178 B.n941 B.n461 163.367
R2179 B.n945 B.n461 163.367
R2180 B.n945 B.n455 163.367
R2181 B.n953 B.n455 163.367
R2182 B.n953 B.n453 163.367
R2183 B.n957 B.n453 163.367
R2184 B.n957 B.n447 163.367
R2185 B.n965 B.n447 163.367
R2186 B.n965 B.n445 163.367
R2187 B.n969 B.n445 163.367
R2188 B.n969 B.n439 163.367
R2189 B.n977 B.n439 163.367
R2190 B.n977 B.n437 163.367
R2191 B.n981 B.n437 163.367
R2192 B.n981 B.n431 163.367
R2193 B.n989 B.n431 163.367
R2194 B.n989 B.n429 163.367
R2195 B.n993 B.n429 163.367
R2196 B.n993 B.n423 163.367
R2197 B.n1002 B.n423 163.367
R2198 B.n1002 B.n421 163.367
R2199 B.n1006 B.n421 163.367
R2200 B.n1006 B.n3 163.367
R2201 B.n1200 B.n3 163.367
R2202 B.n1196 B.n2 163.367
R2203 B.n1196 B.n1195 163.367
R2204 B.n1195 B.n9 163.367
R2205 B.n1191 B.n9 163.367
R2206 B.n1191 B.n11 163.367
R2207 B.n1187 B.n11 163.367
R2208 B.n1187 B.n17 163.367
R2209 B.n1183 B.n17 163.367
R2210 B.n1183 B.n19 163.367
R2211 B.n1179 B.n19 163.367
R2212 B.n1179 B.n24 163.367
R2213 B.n1175 B.n24 163.367
R2214 B.n1175 B.n26 163.367
R2215 B.n1171 B.n26 163.367
R2216 B.n1171 B.n31 163.367
R2217 B.n1167 B.n31 163.367
R2218 B.n1167 B.n33 163.367
R2219 B.n1163 B.n33 163.367
R2220 B.n1163 B.n38 163.367
R2221 B.n1159 B.n38 163.367
R2222 B.n1159 B.n40 163.367
R2223 B.n1155 B.n40 163.367
R2224 B.n1155 B.n45 163.367
R2225 B.n1151 B.n45 163.367
R2226 B.n1151 B.n47 163.367
R2227 B.n1147 B.n47 163.367
R2228 B.n1147 B.n52 163.367
R2229 B.n1143 B.n52 163.367
R2230 B.n1143 B.n54 163.367
R2231 B.n1139 B.n54 163.367
R2232 B.n1139 B.n59 163.367
R2233 B.n1135 B.n59 163.367
R2234 B.n1135 B.n61 163.367
R2235 B.n1131 B.n61 163.367
R2236 B.n1131 B.n66 163.367
R2237 B.n1127 B.n66 163.367
R2238 B.n1127 B.n68 163.367
R2239 B.n1123 B.n68 163.367
R2240 B.n1123 B.n73 163.367
R2241 B.n1119 B.n73 163.367
R2242 B.n1119 B.n75 163.367
R2243 B.n1115 B.n75 163.367
R2244 B.n1115 B.n80 163.367
R2245 B.n1111 B.n80 163.367
R2246 B.n1111 B.n82 163.367
R2247 B.n1107 B.n82 163.367
R2248 B.n1107 B.n87 163.367
R2249 B.n1103 B.n87 163.367
R2250 B.n1103 B.n89 163.367
R2251 B.n1099 B.n89 163.367
R2252 B.n1099 B.n94 163.367
R2253 B.n1095 B.n94 163.367
R2254 B.n1095 B.n96 163.367
R2255 B.n1091 B.n96 163.367
R2256 B.n1091 B.n101 163.367
R2257 B.n1087 B.n1086 71.676
R2258 B.n173 B.n104 71.676
R2259 B.n177 B.n105 71.676
R2260 B.n181 B.n106 71.676
R2261 B.n185 B.n107 71.676
R2262 B.n189 B.n108 71.676
R2263 B.n193 B.n109 71.676
R2264 B.n197 B.n110 71.676
R2265 B.n201 B.n111 71.676
R2266 B.n205 B.n112 71.676
R2267 B.n209 B.n113 71.676
R2268 B.n213 B.n114 71.676
R2269 B.n217 B.n115 71.676
R2270 B.n221 B.n116 71.676
R2271 B.n225 B.n117 71.676
R2272 B.n229 B.n118 71.676
R2273 B.n233 B.n119 71.676
R2274 B.n237 B.n120 71.676
R2275 B.n241 B.n121 71.676
R2276 B.n245 B.n122 71.676
R2277 B.n249 B.n123 71.676
R2278 B.n253 B.n124 71.676
R2279 B.n257 B.n125 71.676
R2280 B.n261 B.n126 71.676
R2281 B.n265 B.n127 71.676
R2282 B.n269 B.n128 71.676
R2283 B.n273 B.n129 71.676
R2284 B.n277 B.n130 71.676
R2285 B.n281 B.n131 71.676
R2286 B.n285 B.n132 71.676
R2287 B.n289 B.n133 71.676
R2288 B.n293 B.n134 71.676
R2289 B.n297 B.n135 71.676
R2290 B.n301 B.n136 71.676
R2291 B.n305 B.n137 71.676
R2292 B.n309 B.n138 71.676
R2293 B.n313 B.n139 71.676
R2294 B.n317 B.n140 71.676
R2295 B.n321 B.n141 71.676
R2296 B.n325 B.n142 71.676
R2297 B.n329 B.n143 71.676
R2298 B.n333 B.n144 71.676
R2299 B.n337 B.n145 71.676
R2300 B.n341 B.n146 71.676
R2301 B.n345 B.n147 71.676
R2302 B.n349 B.n148 71.676
R2303 B.n353 B.n149 71.676
R2304 B.n357 B.n150 71.676
R2305 B.n361 B.n151 71.676
R2306 B.n365 B.n152 71.676
R2307 B.n369 B.n153 71.676
R2308 B.n373 B.n154 71.676
R2309 B.n377 B.n155 71.676
R2310 B.n381 B.n156 71.676
R2311 B.n385 B.n157 71.676
R2312 B.n389 B.n158 71.676
R2313 B.n393 B.n159 71.676
R2314 B.n397 B.n160 71.676
R2315 B.n401 B.n161 71.676
R2316 B.n405 B.n162 71.676
R2317 B.n409 B.n163 71.676
R2318 B.n413 B.n164 71.676
R2319 B.n1084 B.n165 71.676
R2320 B.n1084 B.n1083 71.676
R2321 B.n415 B.n164 71.676
R2322 B.n412 B.n163 71.676
R2323 B.n408 B.n162 71.676
R2324 B.n404 B.n161 71.676
R2325 B.n400 B.n160 71.676
R2326 B.n396 B.n159 71.676
R2327 B.n392 B.n158 71.676
R2328 B.n388 B.n157 71.676
R2329 B.n384 B.n156 71.676
R2330 B.n380 B.n155 71.676
R2331 B.n376 B.n154 71.676
R2332 B.n372 B.n153 71.676
R2333 B.n368 B.n152 71.676
R2334 B.n364 B.n151 71.676
R2335 B.n360 B.n150 71.676
R2336 B.n356 B.n149 71.676
R2337 B.n352 B.n148 71.676
R2338 B.n348 B.n147 71.676
R2339 B.n344 B.n146 71.676
R2340 B.n340 B.n145 71.676
R2341 B.n336 B.n144 71.676
R2342 B.n332 B.n143 71.676
R2343 B.n328 B.n142 71.676
R2344 B.n324 B.n141 71.676
R2345 B.n320 B.n140 71.676
R2346 B.n316 B.n139 71.676
R2347 B.n312 B.n138 71.676
R2348 B.n308 B.n137 71.676
R2349 B.n304 B.n136 71.676
R2350 B.n300 B.n135 71.676
R2351 B.n296 B.n134 71.676
R2352 B.n292 B.n133 71.676
R2353 B.n288 B.n132 71.676
R2354 B.n284 B.n131 71.676
R2355 B.n280 B.n130 71.676
R2356 B.n276 B.n129 71.676
R2357 B.n272 B.n128 71.676
R2358 B.n268 B.n127 71.676
R2359 B.n264 B.n126 71.676
R2360 B.n260 B.n125 71.676
R2361 B.n256 B.n124 71.676
R2362 B.n252 B.n123 71.676
R2363 B.n248 B.n122 71.676
R2364 B.n244 B.n121 71.676
R2365 B.n240 B.n120 71.676
R2366 B.n236 B.n119 71.676
R2367 B.n232 B.n118 71.676
R2368 B.n228 B.n117 71.676
R2369 B.n224 B.n116 71.676
R2370 B.n220 B.n115 71.676
R2371 B.n216 B.n114 71.676
R2372 B.n212 B.n113 71.676
R2373 B.n208 B.n112 71.676
R2374 B.n204 B.n111 71.676
R2375 B.n200 B.n110 71.676
R2376 B.n196 B.n109 71.676
R2377 B.n192 B.n108 71.676
R2378 B.n188 B.n107 71.676
R2379 B.n184 B.n106 71.676
R2380 B.n180 B.n105 71.676
R2381 B.n176 B.n104 71.676
R2382 B.n1086 B.n103 71.676
R2383 B.n845 B.n844 71.676
R2384 B.n590 B.n528 71.676
R2385 B.n837 B.n529 71.676
R2386 B.n833 B.n530 71.676
R2387 B.n829 B.n531 71.676
R2388 B.n825 B.n532 71.676
R2389 B.n821 B.n533 71.676
R2390 B.n817 B.n534 71.676
R2391 B.n813 B.n535 71.676
R2392 B.n809 B.n536 71.676
R2393 B.n805 B.n537 71.676
R2394 B.n801 B.n538 71.676
R2395 B.n797 B.n539 71.676
R2396 B.n793 B.n540 71.676
R2397 B.n789 B.n541 71.676
R2398 B.n785 B.n542 71.676
R2399 B.n781 B.n543 71.676
R2400 B.n777 B.n544 71.676
R2401 B.n773 B.n545 71.676
R2402 B.n769 B.n546 71.676
R2403 B.n765 B.n547 71.676
R2404 B.n761 B.n548 71.676
R2405 B.n757 B.n549 71.676
R2406 B.n753 B.n550 71.676
R2407 B.n749 B.n551 71.676
R2408 B.n745 B.n552 71.676
R2409 B.n741 B.n553 71.676
R2410 B.n737 B.n554 71.676
R2411 B.n733 B.n555 71.676
R2412 B.n728 B.n556 71.676
R2413 B.n724 B.n557 71.676
R2414 B.n720 B.n558 71.676
R2415 B.n716 B.n559 71.676
R2416 B.n712 B.n560 71.676
R2417 B.n707 B.n561 71.676
R2418 B.n703 B.n562 71.676
R2419 B.n699 B.n563 71.676
R2420 B.n695 B.n564 71.676
R2421 B.n691 B.n565 71.676
R2422 B.n687 B.n566 71.676
R2423 B.n683 B.n567 71.676
R2424 B.n679 B.n568 71.676
R2425 B.n675 B.n569 71.676
R2426 B.n671 B.n570 71.676
R2427 B.n667 B.n571 71.676
R2428 B.n663 B.n572 71.676
R2429 B.n659 B.n573 71.676
R2430 B.n655 B.n574 71.676
R2431 B.n651 B.n575 71.676
R2432 B.n647 B.n576 71.676
R2433 B.n643 B.n577 71.676
R2434 B.n639 B.n578 71.676
R2435 B.n635 B.n579 71.676
R2436 B.n631 B.n580 71.676
R2437 B.n627 B.n581 71.676
R2438 B.n623 B.n582 71.676
R2439 B.n619 B.n583 71.676
R2440 B.n615 B.n584 71.676
R2441 B.n611 B.n585 71.676
R2442 B.n607 B.n586 71.676
R2443 B.n603 B.n587 71.676
R2444 B.n599 B.n588 71.676
R2445 B.n844 B.n527 71.676
R2446 B.n838 B.n528 71.676
R2447 B.n834 B.n529 71.676
R2448 B.n830 B.n530 71.676
R2449 B.n826 B.n531 71.676
R2450 B.n822 B.n532 71.676
R2451 B.n818 B.n533 71.676
R2452 B.n814 B.n534 71.676
R2453 B.n810 B.n535 71.676
R2454 B.n806 B.n536 71.676
R2455 B.n802 B.n537 71.676
R2456 B.n798 B.n538 71.676
R2457 B.n794 B.n539 71.676
R2458 B.n790 B.n540 71.676
R2459 B.n786 B.n541 71.676
R2460 B.n782 B.n542 71.676
R2461 B.n778 B.n543 71.676
R2462 B.n774 B.n544 71.676
R2463 B.n770 B.n545 71.676
R2464 B.n766 B.n546 71.676
R2465 B.n762 B.n547 71.676
R2466 B.n758 B.n548 71.676
R2467 B.n754 B.n549 71.676
R2468 B.n750 B.n550 71.676
R2469 B.n746 B.n551 71.676
R2470 B.n742 B.n552 71.676
R2471 B.n738 B.n553 71.676
R2472 B.n734 B.n554 71.676
R2473 B.n729 B.n555 71.676
R2474 B.n725 B.n556 71.676
R2475 B.n721 B.n557 71.676
R2476 B.n717 B.n558 71.676
R2477 B.n713 B.n559 71.676
R2478 B.n708 B.n560 71.676
R2479 B.n704 B.n561 71.676
R2480 B.n700 B.n562 71.676
R2481 B.n696 B.n563 71.676
R2482 B.n692 B.n564 71.676
R2483 B.n688 B.n565 71.676
R2484 B.n684 B.n566 71.676
R2485 B.n680 B.n567 71.676
R2486 B.n676 B.n568 71.676
R2487 B.n672 B.n569 71.676
R2488 B.n668 B.n570 71.676
R2489 B.n664 B.n571 71.676
R2490 B.n660 B.n572 71.676
R2491 B.n656 B.n573 71.676
R2492 B.n652 B.n574 71.676
R2493 B.n648 B.n575 71.676
R2494 B.n644 B.n576 71.676
R2495 B.n640 B.n577 71.676
R2496 B.n636 B.n578 71.676
R2497 B.n632 B.n579 71.676
R2498 B.n628 B.n580 71.676
R2499 B.n624 B.n581 71.676
R2500 B.n620 B.n582 71.676
R2501 B.n616 B.n583 71.676
R2502 B.n612 B.n584 71.676
R2503 B.n608 B.n585 71.676
R2504 B.n604 B.n586 71.676
R2505 B.n600 B.n587 71.676
R2506 B.n596 B.n588 71.676
R2507 B.n1201 B.n1200 71.676
R2508 B.n1201 B.n2 71.676
R2509 B.n172 B.n171 59.5399
R2510 B.n169 B.n168 59.5399
R2511 B.n710 B.n594 59.5399
R2512 B.n731 B.n592 59.5399
R2513 B.n843 B.n524 56.2137
R2514 B.n1085 B.n100 56.2137
R2515 B.n171 B.n170 51.9763
R2516 B.n168 B.n167 51.9763
R2517 B.n594 B.n593 51.9763
R2518 B.n592 B.n591 51.9763
R2519 B.n850 B.n524 32.6714
R2520 B.n850 B.n520 32.6714
R2521 B.n856 B.n520 32.6714
R2522 B.n856 B.n516 32.6714
R2523 B.n862 B.n516 32.6714
R2524 B.n862 B.n512 32.6714
R2525 B.n868 B.n512 32.6714
R2526 B.n874 B.n508 32.6714
R2527 B.n874 B.n504 32.6714
R2528 B.n880 B.n504 32.6714
R2529 B.n880 B.n500 32.6714
R2530 B.n886 B.n500 32.6714
R2531 B.n886 B.n496 32.6714
R2532 B.n892 B.n496 32.6714
R2533 B.n892 B.n491 32.6714
R2534 B.n898 B.n491 32.6714
R2535 B.n898 B.n492 32.6714
R2536 B.n904 B.n484 32.6714
R2537 B.n910 B.n484 32.6714
R2538 B.n910 B.n480 32.6714
R2539 B.n916 B.n480 32.6714
R2540 B.n916 B.n475 32.6714
R2541 B.n922 B.n475 32.6714
R2542 B.n922 B.n476 32.6714
R2543 B.n928 B.n468 32.6714
R2544 B.n934 B.n468 32.6714
R2545 B.n934 B.n464 32.6714
R2546 B.n940 B.n464 32.6714
R2547 B.n940 B.n459 32.6714
R2548 B.n946 B.n459 32.6714
R2549 B.n946 B.n460 32.6714
R2550 B.n952 B.n452 32.6714
R2551 B.n958 B.n452 32.6714
R2552 B.n958 B.n448 32.6714
R2553 B.n964 B.n448 32.6714
R2554 B.n964 B.n443 32.6714
R2555 B.n970 B.n443 32.6714
R2556 B.n970 B.n444 32.6714
R2557 B.n976 B.n436 32.6714
R2558 B.n982 B.n436 32.6714
R2559 B.n982 B.n432 32.6714
R2560 B.n988 B.n432 32.6714
R2561 B.n988 B.n428 32.6714
R2562 B.n994 B.n428 32.6714
R2563 B.n1001 B.n424 32.6714
R2564 B.n1001 B.n420 32.6714
R2565 B.n1007 B.n420 32.6714
R2566 B.n1007 B.n4 32.6714
R2567 B.n1199 B.n4 32.6714
R2568 B.n1199 B.n1198 32.6714
R2569 B.n1198 B.n1197 32.6714
R2570 B.n1197 B.n8 32.6714
R2571 B.n12 B.n8 32.6714
R2572 B.n1190 B.n12 32.6714
R2573 B.n1190 B.n1189 32.6714
R2574 B.n1188 B.n16 32.6714
R2575 B.n1182 B.n16 32.6714
R2576 B.n1182 B.n1181 32.6714
R2577 B.n1181 B.n1180 32.6714
R2578 B.n1180 B.n23 32.6714
R2579 B.n1174 B.n23 32.6714
R2580 B.n1173 B.n1172 32.6714
R2581 B.n1172 B.n30 32.6714
R2582 B.n1166 B.n30 32.6714
R2583 B.n1166 B.n1165 32.6714
R2584 B.n1165 B.n1164 32.6714
R2585 B.n1164 B.n37 32.6714
R2586 B.n1158 B.n37 32.6714
R2587 B.n1157 B.n1156 32.6714
R2588 B.n1156 B.n44 32.6714
R2589 B.n1150 B.n44 32.6714
R2590 B.n1150 B.n1149 32.6714
R2591 B.n1149 B.n1148 32.6714
R2592 B.n1148 B.n51 32.6714
R2593 B.n1142 B.n51 32.6714
R2594 B.n1141 B.n1140 32.6714
R2595 B.n1140 B.n58 32.6714
R2596 B.n1134 B.n58 32.6714
R2597 B.n1134 B.n1133 32.6714
R2598 B.n1133 B.n1132 32.6714
R2599 B.n1132 B.n65 32.6714
R2600 B.n1126 B.n65 32.6714
R2601 B.n1125 B.n1124 32.6714
R2602 B.n1124 B.n72 32.6714
R2603 B.n1118 B.n72 32.6714
R2604 B.n1118 B.n1117 32.6714
R2605 B.n1117 B.n1116 32.6714
R2606 B.n1116 B.n79 32.6714
R2607 B.n1110 B.n79 32.6714
R2608 B.n1110 B.n1109 32.6714
R2609 B.n1109 B.n1108 32.6714
R2610 B.n1108 B.n86 32.6714
R2611 B.n1102 B.n1101 32.6714
R2612 B.n1101 B.n1100 32.6714
R2613 B.n1100 B.n93 32.6714
R2614 B.n1094 B.n93 32.6714
R2615 B.n1094 B.n1093 32.6714
R2616 B.n1093 B.n1092 32.6714
R2617 B.n1092 B.n100 32.6714
R2618 B.n994 B.t3 31.23
R2619 B.t9 B.n1188 31.23
R2620 B.n847 B.n846 30.7517
R2621 B.n595 B.n522 30.7517
R2622 B.n1082 B.n1081 30.7517
R2623 B.n1089 B.n1088 30.7517
R2624 B.n976 B.t8 30.2691
R2625 B.n1174 B.t4 30.2691
R2626 B.n952 B.t6 26.4255
R2627 B.n1158 B.t1 26.4255
R2628 B.n928 B.t0 22.5819
R2629 B.n1142 B.t5 22.5819
R2630 B.t11 B.n508 21.6209
R2631 B.t15 B.n86 21.6209
R2632 B.n904 B.t7 18.7382
R2633 B.n1126 B.t2 18.7382
R2634 B B.n1202 18.0485
R2635 B.n492 B.t7 13.9337
R2636 B.t2 B.n1125 13.9337
R2637 B.n868 B.t11 11.0509
R2638 B.n1102 B.t15 11.0509
R2639 B.n848 B.n847 10.6151
R2640 B.n848 B.n518 10.6151
R2641 B.n858 B.n518 10.6151
R2642 B.n859 B.n858 10.6151
R2643 B.n860 B.n859 10.6151
R2644 B.n860 B.n510 10.6151
R2645 B.n870 B.n510 10.6151
R2646 B.n871 B.n870 10.6151
R2647 B.n872 B.n871 10.6151
R2648 B.n872 B.n502 10.6151
R2649 B.n882 B.n502 10.6151
R2650 B.n883 B.n882 10.6151
R2651 B.n884 B.n883 10.6151
R2652 B.n884 B.n494 10.6151
R2653 B.n894 B.n494 10.6151
R2654 B.n895 B.n894 10.6151
R2655 B.n896 B.n895 10.6151
R2656 B.n896 B.n486 10.6151
R2657 B.n906 B.n486 10.6151
R2658 B.n907 B.n906 10.6151
R2659 B.n908 B.n907 10.6151
R2660 B.n908 B.n478 10.6151
R2661 B.n918 B.n478 10.6151
R2662 B.n919 B.n918 10.6151
R2663 B.n920 B.n919 10.6151
R2664 B.n920 B.n470 10.6151
R2665 B.n930 B.n470 10.6151
R2666 B.n931 B.n930 10.6151
R2667 B.n932 B.n931 10.6151
R2668 B.n932 B.n462 10.6151
R2669 B.n942 B.n462 10.6151
R2670 B.n943 B.n942 10.6151
R2671 B.n944 B.n943 10.6151
R2672 B.n944 B.n454 10.6151
R2673 B.n954 B.n454 10.6151
R2674 B.n955 B.n954 10.6151
R2675 B.n956 B.n955 10.6151
R2676 B.n956 B.n446 10.6151
R2677 B.n966 B.n446 10.6151
R2678 B.n967 B.n966 10.6151
R2679 B.n968 B.n967 10.6151
R2680 B.n968 B.n438 10.6151
R2681 B.n978 B.n438 10.6151
R2682 B.n979 B.n978 10.6151
R2683 B.n980 B.n979 10.6151
R2684 B.n980 B.n430 10.6151
R2685 B.n990 B.n430 10.6151
R2686 B.n991 B.n990 10.6151
R2687 B.n992 B.n991 10.6151
R2688 B.n992 B.n422 10.6151
R2689 B.n1003 B.n422 10.6151
R2690 B.n1004 B.n1003 10.6151
R2691 B.n1005 B.n1004 10.6151
R2692 B.n1005 B.n0 10.6151
R2693 B.n846 B.n526 10.6151
R2694 B.n841 B.n526 10.6151
R2695 B.n841 B.n840 10.6151
R2696 B.n840 B.n839 10.6151
R2697 B.n839 B.n836 10.6151
R2698 B.n836 B.n835 10.6151
R2699 B.n835 B.n832 10.6151
R2700 B.n832 B.n831 10.6151
R2701 B.n831 B.n828 10.6151
R2702 B.n828 B.n827 10.6151
R2703 B.n827 B.n824 10.6151
R2704 B.n824 B.n823 10.6151
R2705 B.n823 B.n820 10.6151
R2706 B.n820 B.n819 10.6151
R2707 B.n819 B.n816 10.6151
R2708 B.n816 B.n815 10.6151
R2709 B.n815 B.n812 10.6151
R2710 B.n812 B.n811 10.6151
R2711 B.n811 B.n808 10.6151
R2712 B.n808 B.n807 10.6151
R2713 B.n807 B.n804 10.6151
R2714 B.n804 B.n803 10.6151
R2715 B.n803 B.n800 10.6151
R2716 B.n800 B.n799 10.6151
R2717 B.n799 B.n796 10.6151
R2718 B.n796 B.n795 10.6151
R2719 B.n795 B.n792 10.6151
R2720 B.n792 B.n791 10.6151
R2721 B.n791 B.n788 10.6151
R2722 B.n788 B.n787 10.6151
R2723 B.n787 B.n784 10.6151
R2724 B.n784 B.n783 10.6151
R2725 B.n783 B.n780 10.6151
R2726 B.n780 B.n779 10.6151
R2727 B.n779 B.n776 10.6151
R2728 B.n776 B.n775 10.6151
R2729 B.n775 B.n772 10.6151
R2730 B.n772 B.n771 10.6151
R2731 B.n771 B.n768 10.6151
R2732 B.n768 B.n767 10.6151
R2733 B.n767 B.n764 10.6151
R2734 B.n764 B.n763 10.6151
R2735 B.n763 B.n760 10.6151
R2736 B.n760 B.n759 10.6151
R2737 B.n759 B.n756 10.6151
R2738 B.n756 B.n755 10.6151
R2739 B.n755 B.n752 10.6151
R2740 B.n752 B.n751 10.6151
R2741 B.n751 B.n748 10.6151
R2742 B.n748 B.n747 10.6151
R2743 B.n747 B.n744 10.6151
R2744 B.n744 B.n743 10.6151
R2745 B.n743 B.n740 10.6151
R2746 B.n740 B.n739 10.6151
R2747 B.n739 B.n736 10.6151
R2748 B.n736 B.n735 10.6151
R2749 B.n735 B.n732 10.6151
R2750 B.n730 B.n727 10.6151
R2751 B.n727 B.n726 10.6151
R2752 B.n726 B.n723 10.6151
R2753 B.n723 B.n722 10.6151
R2754 B.n722 B.n719 10.6151
R2755 B.n719 B.n718 10.6151
R2756 B.n718 B.n715 10.6151
R2757 B.n715 B.n714 10.6151
R2758 B.n714 B.n711 10.6151
R2759 B.n709 B.n706 10.6151
R2760 B.n706 B.n705 10.6151
R2761 B.n705 B.n702 10.6151
R2762 B.n702 B.n701 10.6151
R2763 B.n701 B.n698 10.6151
R2764 B.n698 B.n697 10.6151
R2765 B.n697 B.n694 10.6151
R2766 B.n694 B.n693 10.6151
R2767 B.n693 B.n690 10.6151
R2768 B.n690 B.n689 10.6151
R2769 B.n689 B.n686 10.6151
R2770 B.n686 B.n685 10.6151
R2771 B.n685 B.n682 10.6151
R2772 B.n682 B.n681 10.6151
R2773 B.n681 B.n678 10.6151
R2774 B.n678 B.n677 10.6151
R2775 B.n677 B.n674 10.6151
R2776 B.n674 B.n673 10.6151
R2777 B.n673 B.n670 10.6151
R2778 B.n670 B.n669 10.6151
R2779 B.n669 B.n666 10.6151
R2780 B.n666 B.n665 10.6151
R2781 B.n665 B.n662 10.6151
R2782 B.n662 B.n661 10.6151
R2783 B.n661 B.n658 10.6151
R2784 B.n658 B.n657 10.6151
R2785 B.n657 B.n654 10.6151
R2786 B.n654 B.n653 10.6151
R2787 B.n653 B.n650 10.6151
R2788 B.n650 B.n649 10.6151
R2789 B.n649 B.n646 10.6151
R2790 B.n646 B.n645 10.6151
R2791 B.n645 B.n642 10.6151
R2792 B.n642 B.n641 10.6151
R2793 B.n641 B.n638 10.6151
R2794 B.n638 B.n637 10.6151
R2795 B.n637 B.n634 10.6151
R2796 B.n634 B.n633 10.6151
R2797 B.n633 B.n630 10.6151
R2798 B.n630 B.n629 10.6151
R2799 B.n629 B.n626 10.6151
R2800 B.n626 B.n625 10.6151
R2801 B.n625 B.n622 10.6151
R2802 B.n622 B.n621 10.6151
R2803 B.n621 B.n618 10.6151
R2804 B.n618 B.n617 10.6151
R2805 B.n617 B.n614 10.6151
R2806 B.n614 B.n613 10.6151
R2807 B.n613 B.n610 10.6151
R2808 B.n610 B.n609 10.6151
R2809 B.n609 B.n606 10.6151
R2810 B.n606 B.n605 10.6151
R2811 B.n605 B.n602 10.6151
R2812 B.n602 B.n601 10.6151
R2813 B.n601 B.n598 10.6151
R2814 B.n598 B.n597 10.6151
R2815 B.n597 B.n595 10.6151
R2816 B.n852 B.n522 10.6151
R2817 B.n853 B.n852 10.6151
R2818 B.n854 B.n853 10.6151
R2819 B.n854 B.n514 10.6151
R2820 B.n864 B.n514 10.6151
R2821 B.n865 B.n864 10.6151
R2822 B.n866 B.n865 10.6151
R2823 B.n866 B.n506 10.6151
R2824 B.n876 B.n506 10.6151
R2825 B.n877 B.n876 10.6151
R2826 B.n878 B.n877 10.6151
R2827 B.n878 B.n498 10.6151
R2828 B.n888 B.n498 10.6151
R2829 B.n889 B.n888 10.6151
R2830 B.n890 B.n889 10.6151
R2831 B.n890 B.n489 10.6151
R2832 B.n900 B.n489 10.6151
R2833 B.n901 B.n900 10.6151
R2834 B.n902 B.n901 10.6151
R2835 B.n902 B.n482 10.6151
R2836 B.n912 B.n482 10.6151
R2837 B.n913 B.n912 10.6151
R2838 B.n914 B.n913 10.6151
R2839 B.n914 B.n473 10.6151
R2840 B.n924 B.n473 10.6151
R2841 B.n925 B.n924 10.6151
R2842 B.n926 B.n925 10.6151
R2843 B.n926 B.n466 10.6151
R2844 B.n936 B.n466 10.6151
R2845 B.n937 B.n936 10.6151
R2846 B.n938 B.n937 10.6151
R2847 B.n938 B.n457 10.6151
R2848 B.n948 B.n457 10.6151
R2849 B.n949 B.n948 10.6151
R2850 B.n950 B.n949 10.6151
R2851 B.n950 B.n450 10.6151
R2852 B.n960 B.n450 10.6151
R2853 B.n961 B.n960 10.6151
R2854 B.n962 B.n961 10.6151
R2855 B.n962 B.n441 10.6151
R2856 B.n972 B.n441 10.6151
R2857 B.n973 B.n972 10.6151
R2858 B.n974 B.n973 10.6151
R2859 B.n974 B.n434 10.6151
R2860 B.n984 B.n434 10.6151
R2861 B.n985 B.n984 10.6151
R2862 B.n986 B.n985 10.6151
R2863 B.n986 B.n426 10.6151
R2864 B.n996 B.n426 10.6151
R2865 B.n997 B.n996 10.6151
R2866 B.n999 B.n997 10.6151
R2867 B.n999 B.n998 10.6151
R2868 B.n998 B.n418 10.6151
R2869 B.n1010 B.n418 10.6151
R2870 B.n1011 B.n1010 10.6151
R2871 B.n1012 B.n1011 10.6151
R2872 B.n1013 B.n1012 10.6151
R2873 B.n1014 B.n1013 10.6151
R2874 B.n1017 B.n1014 10.6151
R2875 B.n1018 B.n1017 10.6151
R2876 B.n1019 B.n1018 10.6151
R2877 B.n1020 B.n1019 10.6151
R2878 B.n1022 B.n1020 10.6151
R2879 B.n1023 B.n1022 10.6151
R2880 B.n1024 B.n1023 10.6151
R2881 B.n1025 B.n1024 10.6151
R2882 B.n1027 B.n1025 10.6151
R2883 B.n1028 B.n1027 10.6151
R2884 B.n1029 B.n1028 10.6151
R2885 B.n1030 B.n1029 10.6151
R2886 B.n1032 B.n1030 10.6151
R2887 B.n1033 B.n1032 10.6151
R2888 B.n1034 B.n1033 10.6151
R2889 B.n1035 B.n1034 10.6151
R2890 B.n1037 B.n1035 10.6151
R2891 B.n1038 B.n1037 10.6151
R2892 B.n1039 B.n1038 10.6151
R2893 B.n1040 B.n1039 10.6151
R2894 B.n1042 B.n1040 10.6151
R2895 B.n1043 B.n1042 10.6151
R2896 B.n1044 B.n1043 10.6151
R2897 B.n1045 B.n1044 10.6151
R2898 B.n1047 B.n1045 10.6151
R2899 B.n1048 B.n1047 10.6151
R2900 B.n1049 B.n1048 10.6151
R2901 B.n1050 B.n1049 10.6151
R2902 B.n1052 B.n1050 10.6151
R2903 B.n1053 B.n1052 10.6151
R2904 B.n1054 B.n1053 10.6151
R2905 B.n1055 B.n1054 10.6151
R2906 B.n1057 B.n1055 10.6151
R2907 B.n1058 B.n1057 10.6151
R2908 B.n1059 B.n1058 10.6151
R2909 B.n1060 B.n1059 10.6151
R2910 B.n1062 B.n1060 10.6151
R2911 B.n1063 B.n1062 10.6151
R2912 B.n1064 B.n1063 10.6151
R2913 B.n1065 B.n1064 10.6151
R2914 B.n1067 B.n1065 10.6151
R2915 B.n1068 B.n1067 10.6151
R2916 B.n1069 B.n1068 10.6151
R2917 B.n1070 B.n1069 10.6151
R2918 B.n1072 B.n1070 10.6151
R2919 B.n1073 B.n1072 10.6151
R2920 B.n1074 B.n1073 10.6151
R2921 B.n1075 B.n1074 10.6151
R2922 B.n1077 B.n1075 10.6151
R2923 B.n1078 B.n1077 10.6151
R2924 B.n1079 B.n1078 10.6151
R2925 B.n1080 B.n1079 10.6151
R2926 B.n1081 B.n1080 10.6151
R2927 B.n1194 B.n1 10.6151
R2928 B.n1194 B.n1193 10.6151
R2929 B.n1193 B.n1192 10.6151
R2930 B.n1192 B.n10 10.6151
R2931 B.n1186 B.n10 10.6151
R2932 B.n1186 B.n1185 10.6151
R2933 B.n1185 B.n1184 10.6151
R2934 B.n1184 B.n18 10.6151
R2935 B.n1178 B.n18 10.6151
R2936 B.n1178 B.n1177 10.6151
R2937 B.n1177 B.n1176 10.6151
R2938 B.n1176 B.n25 10.6151
R2939 B.n1170 B.n25 10.6151
R2940 B.n1170 B.n1169 10.6151
R2941 B.n1169 B.n1168 10.6151
R2942 B.n1168 B.n32 10.6151
R2943 B.n1162 B.n32 10.6151
R2944 B.n1162 B.n1161 10.6151
R2945 B.n1161 B.n1160 10.6151
R2946 B.n1160 B.n39 10.6151
R2947 B.n1154 B.n39 10.6151
R2948 B.n1154 B.n1153 10.6151
R2949 B.n1153 B.n1152 10.6151
R2950 B.n1152 B.n46 10.6151
R2951 B.n1146 B.n46 10.6151
R2952 B.n1146 B.n1145 10.6151
R2953 B.n1145 B.n1144 10.6151
R2954 B.n1144 B.n53 10.6151
R2955 B.n1138 B.n53 10.6151
R2956 B.n1138 B.n1137 10.6151
R2957 B.n1137 B.n1136 10.6151
R2958 B.n1136 B.n60 10.6151
R2959 B.n1130 B.n60 10.6151
R2960 B.n1130 B.n1129 10.6151
R2961 B.n1129 B.n1128 10.6151
R2962 B.n1128 B.n67 10.6151
R2963 B.n1122 B.n67 10.6151
R2964 B.n1122 B.n1121 10.6151
R2965 B.n1121 B.n1120 10.6151
R2966 B.n1120 B.n74 10.6151
R2967 B.n1114 B.n74 10.6151
R2968 B.n1114 B.n1113 10.6151
R2969 B.n1113 B.n1112 10.6151
R2970 B.n1112 B.n81 10.6151
R2971 B.n1106 B.n81 10.6151
R2972 B.n1106 B.n1105 10.6151
R2973 B.n1105 B.n1104 10.6151
R2974 B.n1104 B.n88 10.6151
R2975 B.n1098 B.n88 10.6151
R2976 B.n1098 B.n1097 10.6151
R2977 B.n1097 B.n1096 10.6151
R2978 B.n1096 B.n95 10.6151
R2979 B.n1090 B.n95 10.6151
R2980 B.n1090 B.n1089 10.6151
R2981 B.n1088 B.n102 10.6151
R2982 B.n174 B.n102 10.6151
R2983 B.n175 B.n174 10.6151
R2984 B.n178 B.n175 10.6151
R2985 B.n179 B.n178 10.6151
R2986 B.n182 B.n179 10.6151
R2987 B.n183 B.n182 10.6151
R2988 B.n186 B.n183 10.6151
R2989 B.n187 B.n186 10.6151
R2990 B.n190 B.n187 10.6151
R2991 B.n191 B.n190 10.6151
R2992 B.n194 B.n191 10.6151
R2993 B.n195 B.n194 10.6151
R2994 B.n198 B.n195 10.6151
R2995 B.n199 B.n198 10.6151
R2996 B.n202 B.n199 10.6151
R2997 B.n203 B.n202 10.6151
R2998 B.n206 B.n203 10.6151
R2999 B.n207 B.n206 10.6151
R3000 B.n210 B.n207 10.6151
R3001 B.n211 B.n210 10.6151
R3002 B.n214 B.n211 10.6151
R3003 B.n215 B.n214 10.6151
R3004 B.n218 B.n215 10.6151
R3005 B.n219 B.n218 10.6151
R3006 B.n222 B.n219 10.6151
R3007 B.n223 B.n222 10.6151
R3008 B.n226 B.n223 10.6151
R3009 B.n227 B.n226 10.6151
R3010 B.n230 B.n227 10.6151
R3011 B.n231 B.n230 10.6151
R3012 B.n234 B.n231 10.6151
R3013 B.n235 B.n234 10.6151
R3014 B.n238 B.n235 10.6151
R3015 B.n239 B.n238 10.6151
R3016 B.n242 B.n239 10.6151
R3017 B.n243 B.n242 10.6151
R3018 B.n246 B.n243 10.6151
R3019 B.n247 B.n246 10.6151
R3020 B.n250 B.n247 10.6151
R3021 B.n251 B.n250 10.6151
R3022 B.n254 B.n251 10.6151
R3023 B.n255 B.n254 10.6151
R3024 B.n258 B.n255 10.6151
R3025 B.n259 B.n258 10.6151
R3026 B.n262 B.n259 10.6151
R3027 B.n263 B.n262 10.6151
R3028 B.n266 B.n263 10.6151
R3029 B.n267 B.n266 10.6151
R3030 B.n270 B.n267 10.6151
R3031 B.n271 B.n270 10.6151
R3032 B.n274 B.n271 10.6151
R3033 B.n275 B.n274 10.6151
R3034 B.n278 B.n275 10.6151
R3035 B.n279 B.n278 10.6151
R3036 B.n282 B.n279 10.6151
R3037 B.n283 B.n282 10.6151
R3038 B.n287 B.n286 10.6151
R3039 B.n290 B.n287 10.6151
R3040 B.n291 B.n290 10.6151
R3041 B.n294 B.n291 10.6151
R3042 B.n295 B.n294 10.6151
R3043 B.n298 B.n295 10.6151
R3044 B.n299 B.n298 10.6151
R3045 B.n302 B.n299 10.6151
R3046 B.n303 B.n302 10.6151
R3047 B.n307 B.n306 10.6151
R3048 B.n310 B.n307 10.6151
R3049 B.n311 B.n310 10.6151
R3050 B.n314 B.n311 10.6151
R3051 B.n315 B.n314 10.6151
R3052 B.n318 B.n315 10.6151
R3053 B.n319 B.n318 10.6151
R3054 B.n322 B.n319 10.6151
R3055 B.n323 B.n322 10.6151
R3056 B.n326 B.n323 10.6151
R3057 B.n327 B.n326 10.6151
R3058 B.n330 B.n327 10.6151
R3059 B.n331 B.n330 10.6151
R3060 B.n334 B.n331 10.6151
R3061 B.n335 B.n334 10.6151
R3062 B.n338 B.n335 10.6151
R3063 B.n339 B.n338 10.6151
R3064 B.n342 B.n339 10.6151
R3065 B.n343 B.n342 10.6151
R3066 B.n346 B.n343 10.6151
R3067 B.n347 B.n346 10.6151
R3068 B.n350 B.n347 10.6151
R3069 B.n351 B.n350 10.6151
R3070 B.n354 B.n351 10.6151
R3071 B.n355 B.n354 10.6151
R3072 B.n358 B.n355 10.6151
R3073 B.n359 B.n358 10.6151
R3074 B.n362 B.n359 10.6151
R3075 B.n363 B.n362 10.6151
R3076 B.n366 B.n363 10.6151
R3077 B.n367 B.n366 10.6151
R3078 B.n370 B.n367 10.6151
R3079 B.n371 B.n370 10.6151
R3080 B.n374 B.n371 10.6151
R3081 B.n375 B.n374 10.6151
R3082 B.n378 B.n375 10.6151
R3083 B.n379 B.n378 10.6151
R3084 B.n382 B.n379 10.6151
R3085 B.n383 B.n382 10.6151
R3086 B.n386 B.n383 10.6151
R3087 B.n387 B.n386 10.6151
R3088 B.n390 B.n387 10.6151
R3089 B.n391 B.n390 10.6151
R3090 B.n394 B.n391 10.6151
R3091 B.n395 B.n394 10.6151
R3092 B.n398 B.n395 10.6151
R3093 B.n399 B.n398 10.6151
R3094 B.n402 B.n399 10.6151
R3095 B.n403 B.n402 10.6151
R3096 B.n406 B.n403 10.6151
R3097 B.n407 B.n406 10.6151
R3098 B.n410 B.n407 10.6151
R3099 B.n411 B.n410 10.6151
R3100 B.n414 B.n411 10.6151
R3101 B.n416 B.n414 10.6151
R3102 B.n417 B.n416 10.6151
R3103 B.n1082 B.n417 10.6151
R3104 B.n476 B.t0 10.09
R3105 B.t5 B.n1141 10.09
R3106 B.n732 B.n731 9.36635
R3107 B.n710 B.n709 9.36635
R3108 B.n283 B.n172 9.36635
R3109 B.n306 B.n169 9.36635
R3110 B.n1202 B.n0 8.11757
R3111 B.n1202 B.n1 8.11757
R3112 B.n460 B.t6 6.24641
R3113 B.t1 B.n1157 6.24641
R3114 B.n444 B.t8 2.40277
R3115 B.t4 B.n1173 2.40277
R3116 B.t3 B.n424 1.44186
R3117 B.n1189 B.t9 1.44186
R3118 B.n731 B.n730 1.24928
R3119 B.n711 B.n710 1.24928
R3120 B.n286 B.n172 1.24928
R3121 B.n303 B.n169 1.24928
R3122 VN.n8 VN.t9 214.102
R3123 VN.n45 VN.t3 214.102
R3124 VN.n5 VN.t5 180.7
R3125 VN.n9 VN.t8 180.7
R3126 VN.n27 VN.t7 180.7
R3127 VN.n35 VN.t4 180.7
R3128 VN.n42 VN.t2 180.7
R3129 VN.n46 VN.t1 180.7
R3130 VN.n64 VN.t0 180.7
R3131 VN.n72 VN.t6 180.7
R3132 VN.n71 VN.n37 161.3
R3133 VN.n70 VN.n69 161.3
R3134 VN.n68 VN.n38 161.3
R3135 VN.n67 VN.n66 161.3
R3136 VN.n65 VN.n39 161.3
R3137 VN.n63 VN.n62 161.3
R3138 VN.n61 VN.n40 161.3
R3139 VN.n60 VN.n59 161.3
R3140 VN.n58 VN.n41 161.3
R3141 VN.n57 VN.n56 161.3
R3142 VN.n55 VN.n42 161.3
R3143 VN.n54 VN.n53 161.3
R3144 VN.n52 VN.n43 161.3
R3145 VN.n51 VN.n50 161.3
R3146 VN.n49 VN.n44 161.3
R3147 VN.n48 VN.n47 161.3
R3148 VN.n34 VN.n0 161.3
R3149 VN.n33 VN.n32 161.3
R3150 VN.n31 VN.n1 161.3
R3151 VN.n30 VN.n29 161.3
R3152 VN.n28 VN.n2 161.3
R3153 VN.n26 VN.n25 161.3
R3154 VN.n24 VN.n3 161.3
R3155 VN.n23 VN.n22 161.3
R3156 VN.n21 VN.n4 161.3
R3157 VN.n20 VN.n19 161.3
R3158 VN.n18 VN.n5 161.3
R3159 VN.n17 VN.n16 161.3
R3160 VN.n15 VN.n6 161.3
R3161 VN.n14 VN.n13 161.3
R3162 VN.n12 VN.n7 161.3
R3163 VN.n11 VN.n10 161.3
R3164 VN.n36 VN.n35 93.2021
R3165 VN.n73 VN.n72 93.2021
R3166 VN.n9 VN.n8 63.1823
R3167 VN.n46 VN.n45 63.1823
R3168 VN VN.n73 56.3694
R3169 VN.n15 VN.n14 56.0773
R3170 VN.n22 VN.n21 56.0773
R3171 VN.n52 VN.n51 56.0773
R3172 VN.n59 VN.n58 56.0773
R3173 VN.n33 VN.n1 42.5146
R3174 VN.n70 VN.n38 42.5146
R3175 VN.n29 VN.n1 38.6395
R3176 VN.n66 VN.n38 38.6395
R3177 VN.n14 VN.n7 25.0767
R3178 VN.n22 VN.n3 25.0767
R3179 VN.n51 VN.n44 25.0767
R3180 VN.n59 VN.n40 25.0767
R3181 VN.n10 VN.n7 24.5923
R3182 VN.n16 VN.n15 24.5923
R3183 VN.n16 VN.n5 24.5923
R3184 VN.n20 VN.n5 24.5923
R3185 VN.n21 VN.n20 24.5923
R3186 VN.n26 VN.n3 24.5923
R3187 VN.n29 VN.n28 24.5923
R3188 VN.n34 VN.n33 24.5923
R3189 VN.n47 VN.n44 24.5923
R3190 VN.n58 VN.n57 24.5923
R3191 VN.n57 VN.n42 24.5923
R3192 VN.n53 VN.n42 24.5923
R3193 VN.n53 VN.n52 24.5923
R3194 VN.n66 VN.n65 24.5923
R3195 VN.n63 VN.n40 24.5923
R3196 VN.n71 VN.n70 24.5923
R3197 VN.n35 VN.n34 17.7066
R3198 VN.n72 VN.n71 17.7066
R3199 VN.n28 VN.n27 15.7393
R3200 VN.n65 VN.n64 15.7393
R3201 VN.n48 VN.n45 9.19198
R3202 VN.n11 VN.n8 9.19198
R3203 VN.n10 VN.n9 8.85356
R3204 VN.n27 VN.n26 8.85356
R3205 VN.n47 VN.n46 8.85356
R3206 VN.n64 VN.n63 8.85356
R3207 VN.n73 VN.n37 0.278335
R3208 VN.n36 VN.n0 0.278335
R3209 VN.n69 VN.n37 0.189894
R3210 VN.n69 VN.n68 0.189894
R3211 VN.n68 VN.n67 0.189894
R3212 VN.n67 VN.n39 0.189894
R3213 VN.n62 VN.n39 0.189894
R3214 VN.n62 VN.n61 0.189894
R3215 VN.n61 VN.n60 0.189894
R3216 VN.n60 VN.n41 0.189894
R3217 VN.n56 VN.n41 0.189894
R3218 VN.n56 VN.n55 0.189894
R3219 VN.n55 VN.n54 0.189894
R3220 VN.n54 VN.n43 0.189894
R3221 VN.n50 VN.n43 0.189894
R3222 VN.n50 VN.n49 0.189894
R3223 VN.n49 VN.n48 0.189894
R3224 VN.n12 VN.n11 0.189894
R3225 VN.n13 VN.n12 0.189894
R3226 VN.n13 VN.n6 0.189894
R3227 VN.n17 VN.n6 0.189894
R3228 VN.n18 VN.n17 0.189894
R3229 VN.n19 VN.n18 0.189894
R3230 VN.n19 VN.n4 0.189894
R3231 VN.n23 VN.n4 0.189894
R3232 VN.n24 VN.n23 0.189894
R3233 VN.n25 VN.n24 0.189894
R3234 VN.n25 VN.n2 0.189894
R3235 VN.n30 VN.n2 0.189894
R3236 VN.n31 VN.n30 0.189894
R3237 VN.n32 VN.n31 0.189894
R3238 VN.n32 VN.n0 0.189894
R3239 VN VN.n36 0.153485
R3240 VDD2.n193 VDD2.n101 289.615
R3241 VDD2.n92 VDD2.n0 289.615
R3242 VDD2.n194 VDD2.n193 185
R3243 VDD2.n192 VDD2.n191 185
R3244 VDD2.n105 VDD2.n104 185
R3245 VDD2.n186 VDD2.n185 185
R3246 VDD2.n184 VDD2.n183 185
R3247 VDD2.n109 VDD2.n108 185
R3248 VDD2.n113 VDD2.n111 185
R3249 VDD2.n178 VDD2.n177 185
R3250 VDD2.n176 VDD2.n175 185
R3251 VDD2.n115 VDD2.n114 185
R3252 VDD2.n170 VDD2.n169 185
R3253 VDD2.n168 VDD2.n167 185
R3254 VDD2.n119 VDD2.n118 185
R3255 VDD2.n162 VDD2.n161 185
R3256 VDD2.n160 VDD2.n159 185
R3257 VDD2.n123 VDD2.n122 185
R3258 VDD2.n154 VDD2.n153 185
R3259 VDD2.n152 VDD2.n151 185
R3260 VDD2.n127 VDD2.n126 185
R3261 VDD2.n146 VDD2.n145 185
R3262 VDD2.n144 VDD2.n143 185
R3263 VDD2.n131 VDD2.n130 185
R3264 VDD2.n138 VDD2.n137 185
R3265 VDD2.n136 VDD2.n135 185
R3266 VDD2.n33 VDD2.n32 185
R3267 VDD2.n35 VDD2.n34 185
R3268 VDD2.n28 VDD2.n27 185
R3269 VDD2.n41 VDD2.n40 185
R3270 VDD2.n43 VDD2.n42 185
R3271 VDD2.n24 VDD2.n23 185
R3272 VDD2.n49 VDD2.n48 185
R3273 VDD2.n51 VDD2.n50 185
R3274 VDD2.n20 VDD2.n19 185
R3275 VDD2.n57 VDD2.n56 185
R3276 VDD2.n59 VDD2.n58 185
R3277 VDD2.n16 VDD2.n15 185
R3278 VDD2.n65 VDD2.n64 185
R3279 VDD2.n67 VDD2.n66 185
R3280 VDD2.n12 VDD2.n11 185
R3281 VDD2.n74 VDD2.n73 185
R3282 VDD2.n75 VDD2.n10 185
R3283 VDD2.n77 VDD2.n76 185
R3284 VDD2.n8 VDD2.n7 185
R3285 VDD2.n83 VDD2.n82 185
R3286 VDD2.n85 VDD2.n84 185
R3287 VDD2.n4 VDD2.n3 185
R3288 VDD2.n91 VDD2.n90 185
R3289 VDD2.n93 VDD2.n92 185
R3290 VDD2.n134 VDD2.t3 147.659
R3291 VDD2.n31 VDD2.t0 147.659
R3292 VDD2.n193 VDD2.n192 104.615
R3293 VDD2.n192 VDD2.n104 104.615
R3294 VDD2.n185 VDD2.n104 104.615
R3295 VDD2.n185 VDD2.n184 104.615
R3296 VDD2.n184 VDD2.n108 104.615
R3297 VDD2.n113 VDD2.n108 104.615
R3298 VDD2.n177 VDD2.n113 104.615
R3299 VDD2.n177 VDD2.n176 104.615
R3300 VDD2.n176 VDD2.n114 104.615
R3301 VDD2.n169 VDD2.n114 104.615
R3302 VDD2.n169 VDD2.n168 104.615
R3303 VDD2.n168 VDD2.n118 104.615
R3304 VDD2.n161 VDD2.n118 104.615
R3305 VDD2.n161 VDD2.n160 104.615
R3306 VDD2.n160 VDD2.n122 104.615
R3307 VDD2.n153 VDD2.n122 104.615
R3308 VDD2.n153 VDD2.n152 104.615
R3309 VDD2.n152 VDD2.n126 104.615
R3310 VDD2.n145 VDD2.n126 104.615
R3311 VDD2.n145 VDD2.n144 104.615
R3312 VDD2.n144 VDD2.n130 104.615
R3313 VDD2.n137 VDD2.n130 104.615
R3314 VDD2.n137 VDD2.n136 104.615
R3315 VDD2.n34 VDD2.n33 104.615
R3316 VDD2.n34 VDD2.n27 104.615
R3317 VDD2.n41 VDD2.n27 104.615
R3318 VDD2.n42 VDD2.n41 104.615
R3319 VDD2.n42 VDD2.n23 104.615
R3320 VDD2.n49 VDD2.n23 104.615
R3321 VDD2.n50 VDD2.n49 104.615
R3322 VDD2.n50 VDD2.n19 104.615
R3323 VDD2.n57 VDD2.n19 104.615
R3324 VDD2.n58 VDD2.n57 104.615
R3325 VDD2.n58 VDD2.n15 104.615
R3326 VDD2.n65 VDD2.n15 104.615
R3327 VDD2.n66 VDD2.n65 104.615
R3328 VDD2.n66 VDD2.n11 104.615
R3329 VDD2.n74 VDD2.n11 104.615
R3330 VDD2.n75 VDD2.n74 104.615
R3331 VDD2.n76 VDD2.n75 104.615
R3332 VDD2.n76 VDD2.n7 104.615
R3333 VDD2.n83 VDD2.n7 104.615
R3334 VDD2.n84 VDD2.n83 104.615
R3335 VDD2.n84 VDD2.n3 104.615
R3336 VDD2.n91 VDD2.n3 104.615
R3337 VDD2.n92 VDD2.n91 104.615
R3338 VDD2.n100 VDD2.n99 64.2988
R3339 VDD2 VDD2.n201 64.2959
R3340 VDD2.n200 VDD2.n199 62.6215
R3341 VDD2.n98 VDD2.n97 62.6214
R3342 VDD2.n98 VDD2.n96 53.1139
R3343 VDD2.n136 VDD2.t3 52.3082
R3344 VDD2.n33 VDD2.t0 52.3082
R3345 VDD2.n198 VDD2.n197 50.8035
R3346 VDD2.n198 VDD2.n100 49.8791
R3347 VDD2.n135 VDD2.n134 15.6677
R3348 VDD2.n32 VDD2.n31 15.6677
R3349 VDD2.n111 VDD2.n109 13.1884
R3350 VDD2.n77 VDD2.n8 13.1884
R3351 VDD2.n183 VDD2.n182 12.8005
R3352 VDD2.n179 VDD2.n178 12.8005
R3353 VDD2.n138 VDD2.n133 12.8005
R3354 VDD2.n35 VDD2.n30 12.8005
R3355 VDD2.n78 VDD2.n10 12.8005
R3356 VDD2.n82 VDD2.n81 12.8005
R3357 VDD2.n186 VDD2.n107 12.0247
R3358 VDD2.n175 VDD2.n112 12.0247
R3359 VDD2.n139 VDD2.n131 12.0247
R3360 VDD2.n36 VDD2.n28 12.0247
R3361 VDD2.n73 VDD2.n72 12.0247
R3362 VDD2.n85 VDD2.n6 12.0247
R3363 VDD2.n187 VDD2.n105 11.249
R3364 VDD2.n174 VDD2.n115 11.249
R3365 VDD2.n143 VDD2.n142 11.249
R3366 VDD2.n40 VDD2.n39 11.249
R3367 VDD2.n71 VDD2.n12 11.249
R3368 VDD2.n86 VDD2.n4 11.249
R3369 VDD2.n191 VDD2.n190 10.4732
R3370 VDD2.n171 VDD2.n170 10.4732
R3371 VDD2.n146 VDD2.n129 10.4732
R3372 VDD2.n43 VDD2.n26 10.4732
R3373 VDD2.n68 VDD2.n67 10.4732
R3374 VDD2.n90 VDD2.n89 10.4732
R3375 VDD2.n194 VDD2.n103 9.69747
R3376 VDD2.n167 VDD2.n117 9.69747
R3377 VDD2.n147 VDD2.n127 9.69747
R3378 VDD2.n44 VDD2.n24 9.69747
R3379 VDD2.n64 VDD2.n14 9.69747
R3380 VDD2.n93 VDD2.n2 9.69747
R3381 VDD2.n197 VDD2.n196 9.45567
R3382 VDD2.n96 VDD2.n95 9.45567
R3383 VDD2.n121 VDD2.n120 9.3005
R3384 VDD2.n164 VDD2.n163 9.3005
R3385 VDD2.n166 VDD2.n165 9.3005
R3386 VDD2.n117 VDD2.n116 9.3005
R3387 VDD2.n172 VDD2.n171 9.3005
R3388 VDD2.n174 VDD2.n173 9.3005
R3389 VDD2.n112 VDD2.n110 9.3005
R3390 VDD2.n180 VDD2.n179 9.3005
R3391 VDD2.n196 VDD2.n195 9.3005
R3392 VDD2.n103 VDD2.n102 9.3005
R3393 VDD2.n190 VDD2.n189 9.3005
R3394 VDD2.n188 VDD2.n187 9.3005
R3395 VDD2.n107 VDD2.n106 9.3005
R3396 VDD2.n182 VDD2.n181 9.3005
R3397 VDD2.n158 VDD2.n157 9.3005
R3398 VDD2.n156 VDD2.n155 9.3005
R3399 VDD2.n125 VDD2.n124 9.3005
R3400 VDD2.n150 VDD2.n149 9.3005
R3401 VDD2.n148 VDD2.n147 9.3005
R3402 VDD2.n129 VDD2.n128 9.3005
R3403 VDD2.n142 VDD2.n141 9.3005
R3404 VDD2.n140 VDD2.n139 9.3005
R3405 VDD2.n133 VDD2.n132 9.3005
R3406 VDD2.n95 VDD2.n94 9.3005
R3407 VDD2.n2 VDD2.n1 9.3005
R3408 VDD2.n89 VDD2.n88 9.3005
R3409 VDD2.n87 VDD2.n86 9.3005
R3410 VDD2.n6 VDD2.n5 9.3005
R3411 VDD2.n81 VDD2.n80 9.3005
R3412 VDD2.n53 VDD2.n52 9.3005
R3413 VDD2.n22 VDD2.n21 9.3005
R3414 VDD2.n47 VDD2.n46 9.3005
R3415 VDD2.n45 VDD2.n44 9.3005
R3416 VDD2.n26 VDD2.n25 9.3005
R3417 VDD2.n39 VDD2.n38 9.3005
R3418 VDD2.n37 VDD2.n36 9.3005
R3419 VDD2.n30 VDD2.n29 9.3005
R3420 VDD2.n55 VDD2.n54 9.3005
R3421 VDD2.n18 VDD2.n17 9.3005
R3422 VDD2.n61 VDD2.n60 9.3005
R3423 VDD2.n63 VDD2.n62 9.3005
R3424 VDD2.n14 VDD2.n13 9.3005
R3425 VDD2.n69 VDD2.n68 9.3005
R3426 VDD2.n71 VDD2.n70 9.3005
R3427 VDD2.n72 VDD2.n9 9.3005
R3428 VDD2.n79 VDD2.n78 9.3005
R3429 VDD2.n195 VDD2.n101 8.92171
R3430 VDD2.n166 VDD2.n119 8.92171
R3431 VDD2.n151 VDD2.n150 8.92171
R3432 VDD2.n48 VDD2.n47 8.92171
R3433 VDD2.n63 VDD2.n16 8.92171
R3434 VDD2.n94 VDD2.n0 8.92171
R3435 VDD2.n163 VDD2.n162 8.14595
R3436 VDD2.n154 VDD2.n125 8.14595
R3437 VDD2.n51 VDD2.n22 8.14595
R3438 VDD2.n60 VDD2.n59 8.14595
R3439 VDD2.n159 VDD2.n121 7.3702
R3440 VDD2.n155 VDD2.n123 7.3702
R3441 VDD2.n52 VDD2.n20 7.3702
R3442 VDD2.n56 VDD2.n18 7.3702
R3443 VDD2.n159 VDD2.n158 6.59444
R3444 VDD2.n158 VDD2.n123 6.59444
R3445 VDD2.n55 VDD2.n20 6.59444
R3446 VDD2.n56 VDD2.n55 6.59444
R3447 VDD2.n162 VDD2.n121 5.81868
R3448 VDD2.n155 VDD2.n154 5.81868
R3449 VDD2.n52 VDD2.n51 5.81868
R3450 VDD2.n59 VDD2.n18 5.81868
R3451 VDD2.n197 VDD2.n101 5.04292
R3452 VDD2.n163 VDD2.n119 5.04292
R3453 VDD2.n151 VDD2.n125 5.04292
R3454 VDD2.n48 VDD2.n22 5.04292
R3455 VDD2.n60 VDD2.n16 5.04292
R3456 VDD2.n96 VDD2.n0 5.04292
R3457 VDD2.n134 VDD2.n132 4.38563
R3458 VDD2.n31 VDD2.n29 4.38563
R3459 VDD2.n195 VDD2.n194 4.26717
R3460 VDD2.n167 VDD2.n166 4.26717
R3461 VDD2.n150 VDD2.n127 4.26717
R3462 VDD2.n47 VDD2.n24 4.26717
R3463 VDD2.n64 VDD2.n63 4.26717
R3464 VDD2.n94 VDD2.n93 4.26717
R3465 VDD2.n191 VDD2.n103 3.49141
R3466 VDD2.n170 VDD2.n117 3.49141
R3467 VDD2.n147 VDD2.n146 3.49141
R3468 VDD2.n44 VDD2.n43 3.49141
R3469 VDD2.n67 VDD2.n14 3.49141
R3470 VDD2.n90 VDD2.n2 3.49141
R3471 VDD2.n190 VDD2.n105 2.71565
R3472 VDD2.n171 VDD2.n115 2.71565
R3473 VDD2.n143 VDD2.n129 2.71565
R3474 VDD2.n40 VDD2.n26 2.71565
R3475 VDD2.n68 VDD2.n12 2.71565
R3476 VDD2.n89 VDD2.n4 2.71565
R3477 VDD2.n200 VDD2.n198 2.31084
R3478 VDD2.n187 VDD2.n186 1.93989
R3479 VDD2.n175 VDD2.n174 1.93989
R3480 VDD2.n142 VDD2.n131 1.93989
R3481 VDD2.n39 VDD2.n28 1.93989
R3482 VDD2.n73 VDD2.n71 1.93989
R3483 VDD2.n86 VDD2.n85 1.93989
R3484 VDD2.n183 VDD2.n107 1.16414
R3485 VDD2.n178 VDD2.n112 1.16414
R3486 VDD2.n139 VDD2.n138 1.16414
R3487 VDD2.n36 VDD2.n35 1.16414
R3488 VDD2.n72 VDD2.n10 1.16414
R3489 VDD2.n82 VDD2.n6 1.16414
R3490 VDD2.n201 VDD2.t8 1.12422
R3491 VDD2.n201 VDD2.t6 1.12422
R3492 VDD2.n199 VDD2.t9 1.12422
R3493 VDD2.n199 VDD2.t7 1.12422
R3494 VDD2.n99 VDD2.t2 1.12422
R3495 VDD2.n99 VDD2.t5 1.12422
R3496 VDD2.n97 VDD2.t1 1.12422
R3497 VDD2.n97 VDD2.t4 1.12422
R3498 VDD2 VDD2.n200 0.636276
R3499 VDD2.n100 VDD2.n98 0.52274
R3500 VDD2.n182 VDD2.n109 0.388379
R3501 VDD2.n179 VDD2.n111 0.388379
R3502 VDD2.n135 VDD2.n133 0.388379
R3503 VDD2.n32 VDD2.n30 0.388379
R3504 VDD2.n78 VDD2.n77 0.388379
R3505 VDD2.n81 VDD2.n8 0.388379
R3506 VDD2.n196 VDD2.n102 0.155672
R3507 VDD2.n189 VDD2.n102 0.155672
R3508 VDD2.n189 VDD2.n188 0.155672
R3509 VDD2.n188 VDD2.n106 0.155672
R3510 VDD2.n181 VDD2.n106 0.155672
R3511 VDD2.n181 VDD2.n180 0.155672
R3512 VDD2.n180 VDD2.n110 0.155672
R3513 VDD2.n173 VDD2.n110 0.155672
R3514 VDD2.n173 VDD2.n172 0.155672
R3515 VDD2.n172 VDD2.n116 0.155672
R3516 VDD2.n165 VDD2.n116 0.155672
R3517 VDD2.n165 VDD2.n164 0.155672
R3518 VDD2.n164 VDD2.n120 0.155672
R3519 VDD2.n157 VDD2.n120 0.155672
R3520 VDD2.n157 VDD2.n156 0.155672
R3521 VDD2.n156 VDD2.n124 0.155672
R3522 VDD2.n149 VDD2.n124 0.155672
R3523 VDD2.n149 VDD2.n148 0.155672
R3524 VDD2.n148 VDD2.n128 0.155672
R3525 VDD2.n141 VDD2.n128 0.155672
R3526 VDD2.n141 VDD2.n140 0.155672
R3527 VDD2.n140 VDD2.n132 0.155672
R3528 VDD2.n37 VDD2.n29 0.155672
R3529 VDD2.n38 VDD2.n37 0.155672
R3530 VDD2.n38 VDD2.n25 0.155672
R3531 VDD2.n45 VDD2.n25 0.155672
R3532 VDD2.n46 VDD2.n45 0.155672
R3533 VDD2.n46 VDD2.n21 0.155672
R3534 VDD2.n53 VDD2.n21 0.155672
R3535 VDD2.n54 VDD2.n53 0.155672
R3536 VDD2.n54 VDD2.n17 0.155672
R3537 VDD2.n61 VDD2.n17 0.155672
R3538 VDD2.n62 VDD2.n61 0.155672
R3539 VDD2.n62 VDD2.n13 0.155672
R3540 VDD2.n69 VDD2.n13 0.155672
R3541 VDD2.n70 VDD2.n69 0.155672
R3542 VDD2.n70 VDD2.n9 0.155672
R3543 VDD2.n79 VDD2.n9 0.155672
R3544 VDD2.n80 VDD2.n79 0.155672
R3545 VDD2.n80 VDD2.n5 0.155672
R3546 VDD2.n87 VDD2.n5 0.155672
R3547 VDD2.n88 VDD2.n87 0.155672
R3548 VDD2.n88 VDD2.n1 0.155672
R3549 VDD2.n95 VDD2.n1 0.155672
C0 VP VN 9.06185f
C1 VDD1 VDD2 2.01155f
C2 VP VTAIL 15.407598f
C3 VDD1 VN 0.152993f
C4 VDD1 VTAIL 13.096f
C5 VDD2 VN 15.101901f
C6 VDD2 VTAIL 13.1435f
C7 VN VTAIL 15.393201f
C8 VDD1 VP 15.4964f
C9 VDD2 VP 0.552384f
C10 VDD2 B 7.909934f
C11 VDD1 B 7.883769f
C12 VTAIL B 10.23061f
C13 VN B 17.43451f
C14 VP B 15.832864f
C15 VDD2.n0 B 0.033868f
C16 VDD2.n1 B 0.02342f
C17 VDD2.n2 B 0.012585f
C18 VDD2.n3 B 0.029747f
C19 VDD2.n4 B 0.013325f
C20 VDD2.n5 B 0.02342f
C21 VDD2.n6 B 0.012585f
C22 VDD2.n7 B 0.029747f
C23 VDD2.n8 B 0.012955f
C24 VDD2.n9 B 0.02342f
C25 VDD2.n10 B 0.013325f
C26 VDD2.n11 B 0.029747f
C27 VDD2.n12 B 0.013325f
C28 VDD2.n13 B 0.02342f
C29 VDD2.n14 B 0.012585f
C30 VDD2.n15 B 0.029747f
C31 VDD2.n16 B 0.013325f
C32 VDD2.n17 B 0.02342f
C33 VDD2.n18 B 0.012585f
C34 VDD2.n19 B 0.029747f
C35 VDD2.n20 B 0.013325f
C36 VDD2.n21 B 0.02342f
C37 VDD2.n22 B 0.012585f
C38 VDD2.n23 B 0.029747f
C39 VDD2.n24 B 0.013325f
C40 VDD2.n25 B 0.02342f
C41 VDD2.n26 B 0.012585f
C42 VDD2.n27 B 0.029747f
C43 VDD2.n28 B 0.013325f
C44 VDD2.n29 B 1.805f
C45 VDD2.n30 B 0.012585f
C46 VDD2.t0 B 0.049259f
C47 VDD2.n31 B 0.168139f
C48 VDD2.n32 B 0.017572f
C49 VDD2.n33 B 0.02231f
C50 VDD2.n34 B 0.029747f
C51 VDD2.n35 B 0.013325f
C52 VDD2.n36 B 0.012585f
C53 VDD2.n37 B 0.02342f
C54 VDD2.n38 B 0.02342f
C55 VDD2.n39 B 0.012585f
C56 VDD2.n40 B 0.013325f
C57 VDD2.n41 B 0.029747f
C58 VDD2.n42 B 0.029747f
C59 VDD2.n43 B 0.013325f
C60 VDD2.n44 B 0.012585f
C61 VDD2.n45 B 0.02342f
C62 VDD2.n46 B 0.02342f
C63 VDD2.n47 B 0.012585f
C64 VDD2.n48 B 0.013325f
C65 VDD2.n49 B 0.029747f
C66 VDD2.n50 B 0.029747f
C67 VDD2.n51 B 0.013325f
C68 VDD2.n52 B 0.012585f
C69 VDD2.n53 B 0.02342f
C70 VDD2.n54 B 0.02342f
C71 VDD2.n55 B 0.012585f
C72 VDD2.n56 B 0.013325f
C73 VDD2.n57 B 0.029747f
C74 VDD2.n58 B 0.029747f
C75 VDD2.n59 B 0.013325f
C76 VDD2.n60 B 0.012585f
C77 VDD2.n61 B 0.02342f
C78 VDD2.n62 B 0.02342f
C79 VDD2.n63 B 0.012585f
C80 VDD2.n64 B 0.013325f
C81 VDD2.n65 B 0.029747f
C82 VDD2.n66 B 0.029747f
C83 VDD2.n67 B 0.013325f
C84 VDD2.n68 B 0.012585f
C85 VDD2.n69 B 0.02342f
C86 VDD2.n70 B 0.02342f
C87 VDD2.n71 B 0.012585f
C88 VDD2.n72 B 0.012585f
C89 VDD2.n73 B 0.013325f
C90 VDD2.n74 B 0.029747f
C91 VDD2.n75 B 0.029747f
C92 VDD2.n76 B 0.029747f
C93 VDD2.n77 B 0.012955f
C94 VDD2.n78 B 0.012585f
C95 VDD2.n79 B 0.02342f
C96 VDD2.n80 B 0.02342f
C97 VDD2.n81 B 0.012585f
C98 VDD2.n82 B 0.013325f
C99 VDD2.n83 B 0.029747f
C100 VDD2.n84 B 0.029747f
C101 VDD2.n85 B 0.013325f
C102 VDD2.n86 B 0.012585f
C103 VDD2.n87 B 0.02342f
C104 VDD2.n88 B 0.02342f
C105 VDD2.n89 B 0.012585f
C106 VDD2.n90 B 0.013325f
C107 VDD2.n91 B 0.029747f
C108 VDD2.n92 B 0.066073f
C109 VDD2.n93 B 0.013325f
C110 VDD2.n94 B 0.012585f
C111 VDD2.n95 B 0.057335f
C112 VDD2.n96 B 0.063012f
C113 VDD2.t1 B 0.326104f
C114 VDD2.t4 B 0.326104f
C115 VDD2.n97 B 2.97023f
C116 VDD2.n98 B 0.61876f
C117 VDD2.t2 B 0.326104f
C118 VDD2.t5 B 0.326104f
C119 VDD2.n99 B 2.98335f
C120 VDD2.n100 B 2.92792f
C121 VDD2.n101 B 0.033868f
C122 VDD2.n102 B 0.02342f
C123 VDD2.n103 B 0.012585f
C124 VDD2.n104 B 0.029747f
C125 VDD2.n105 B 0.013325f
C126 VDD2.n106 B 0.02342f
C127 VDD2.n107 B 0.012585f
C128 VDD2.n108 B 0.029747f
C129 VDD2.n109 B 0.012955f
C130 VDD2.n110 B 0.02342f
C131 VDD2.n111 B 0.012955f
C132 VDD2.n112 B 0.012585f
C133 VDD2.n113 B 0.029747f
C134 VDD2.n114 B 0.029747f
C135 VDD2.n115 B 0.013325f
C136 VDD2.n116 B 0.02342f
C137 VDD2.n117 B 0.012585f
C138 VDD2.n118 B 0.029747f
C139 VDD2.n119 B 0.013325f
C140 VDD2.n120 B 0.02342f
C141 VDD2.n121 B 0.012585f
C142 VDD2.n122 B 0.029747f
C143 VDD2.n123 B 0.013325f
C144 VDD2.n124 B 0.02342f
C145 VDD2.n125 B 0.012585f
C146 VDD2.n126 B 0.029747f
C147 VDD2.n127 B 0.013325f
C148 VDD2.n128 B 0.02342f
C149 VDD2.n129 B 0.012585f
C150 VDD2.n130 B 0.029747f
C151 VDD2.n131 B 0.013325f
C152 VDD2.n132 B 1.805f
C153 VDD2.n133 B 0.012585f
C154 VDD2.t3 B 0.049259f
C155 VDD2.n134 B 0.168139f
C156 VDD2.n135 B 0.017572f
C157 VDD2.n136 B 0.02231f
C158 VDD2.n137 B 0.029747f
C159 VDD2.n138 B 0.013325f
C160 VDD2.n139 B 0.012585f
C161 VDD2.n140 B 0.02342f
C162 VDD2.n141 B 0.02342f
C163 VDD2.n142 B 0.012585f
C164 VDD2.n143 B 0.013325f
C165 VDD2.n144 B 0.029747f
C166 VDD2.n145 B 0.029747f
C167 VDD2.n146 B 0.013325f
C168 VDD2.n147 B 0.012585f
C169 VDD2.n148 B 0.02342f
C170 VDD2.n149 B 0.02342f
C171 VDD2.n150 B 0.012585f
C172 VDD2.n151 B 0.013325f
C173 VDD2.n152 B 0.029747f
C174 VDD2.n153 B 0.029747f
C175 VDD2.n154 B 0.013325f
C176 VDD2.n155 B 0.012585f
C177 VDD2.n156 B 0.02342f
C178 VDD2.n157 B 0.02342f
C179 VDD2.n158 B 0.012585f
C180 VDD2.n159 B 0.013325f
C181 VDD2.n160 B 0.029747f
C182 VDD2.n161 B 0.029747f
C183 VDD2.n162 B 0.013325f
C184 VDD2.n163 B 0.012585f
C185 VDD2.n164 B 0.02342f
C186 VDD2.n165 B 0.02342f
C187 VDD2.n166 B 0.012585f
C188 VDD2.n167 B 0.013325f
C189 VDD2.n168 B 0.029747f
C190 VDD2.n169 B 0.029747f
C191 VDD2.n170 B 0.013325f
C192 VDD2.n171 B 0.012585f
C193 VDD2.n172 B 0.02342f
C194 VDD2.n173 B 0.02342f
C195 VDD2.n174 B 0.012585f
C196 VDD2.n175 B 0.013325f
C197 VDD2.n176 B 0.029747f
C198 VDD2.n177 B 0.029747f
C199 VDD2.n178 B 0.013325f
C200 VDD2.n179 B 0.012585f
C201 VDD2.n180 B 0.02342f
C202 VDD2.n181 B 0.02342f
C203 VDD2.n182 B 0.012585f
C204 VDD2.n183 B 0.013325f
C205 VDD2.n184 B 0.029747f
C206 VDD2.n185 B 0.029747f
C207 VDD2.n186 B 0.013325f
C208 VDD2.n187 B 0.012585f
C209 VDD2.n188 B 0.02342f
C210 VDD2.n189 B 0.02342f
C211 VDD2.n190 B 0.012585f
C212 VDD2.n191 B 0.013325f
C213 VDD2.n192 B 0.029747f
C214 VDD2.n193 B 0.066073f
C215 VDD2.n194 B 0.013325f
C216 VDD2.n195 B 0.012585f
C217 VDD2.n196 B 0.057335f
C218 VDD2.n197 B 0.053386f
C219 VDD2.n198 B 3.02059f
C220 VDD2.t9 B 0.326104f
C221 VDD2.t7 B 0.326104f
C222 VDD2.n199 B 2.97024f
C223 VDD2.n200 B 0.414622f
C224 VDD2.t8 B 0.326104f
C225 VDD2.t6 B 0.326104f
C226 VDD2.n201 B 2.98331f
C227 VN.n0 B 0.029092f
C228 VN.t4 B 2.51233f
C229 VN.n1 B 0.017936f
C230 VN.n2 B 0.022068f
C231 VN.t7 B 2.51233f
C232 VN.n3 B 0.041305f
C233 VN.n4 B 0.022068f
C234 VN.t5 B 2.51233f
C235 VN.n5 B 0.894514f
C236 VN.n6 B 0.022068f
C237 VN.n7 B 0.041305f
C238 VN.t9 B 2.66837f
C239 VN.n8 B 0.918975f
C240 VN.t8 B 2.51233f
C241 VN.n9 B 0.930212f
C242 VN.n10 B 0.027993f
C243 VN.n11 B 0.190983f
C244 VN.n12 B 0.022068f
C245 VN.n13 B 0.022068f
C246 VN.n14 B 0.026255f
C247 VN.n15 B 0.03752f
C248 VN.n16 B 0.040923f
C249 VN.n17 B 0.022068f
C250 VN.n18 B 0.022068f
C251 VN.n19 B 0.022068f
C252 VN.n20 B 0.040923f
C253 VN.n21 B 0.03752f
C254 VN.n22 B 0.026255f
C255 VN.n23 B 0.022068f
C256 VN.n24 B 0.022068f
C257 VN.n25 B 0.022068f
C258 VN.n26 B 0.027993f
C259 VN.n27 B 0.873794f
C260 VN.n28 B 0.03365f
C261 VN.n29 B 0.044007f
C262 VN.n30 B 0.022068f
C263 VN.n31 B 0.022068f
C264 VN.n32 B 0.022068f
C265 VN.n33 B 0.043137f
C266 VN.n34 B 0.035266f
C267 VN.n35 B 0.949615f
C268 VN.n36 B 0.029636f
C269 VN.n37 B 0.029092f
C270 VN.t6 B 2.51233f
C271 VN.n38 B 0.017936f
C272 VN.n39 B 0.022068f
C273 VN.t0 B 2.51233f
C274 VN.n40 B 0.041305f
C275 VN.n41 B 0.022068f
C276 VN.t2 B 2.51233f
C277 VN.n42 B 0.894514f
C278 VN.n43 B 0.022068f
C279 VN.n44 B 0.041305f
C280 VN.t3 B 2.66837f
C281 VN.n45 B 0.918975f
C282 VN.t1 B 2.51233f
C283 VN.n46 B 0.930212f
C284 VN.n47 B 0.027993f
C285 VN.n48 B 0.190983f
C286 VN.n49 B 0.022068f
C287 VN.n50 B 0.022068f
C288 VN.n51 B 0.026255f
C289 VN.n52 B 0.03752f
C290 VN.n53 B 0.040923f
C291 VN.n54 B 0.022068f
C292 VN.n55 B 0.022068f
C293 VN.n56 B 0.022068f
C294 VN.n57 B 0.040923f
C295 VN.n58 B 0.03752f
C296 VN.n59 B 0.026255f
C297 VN.n60 B 0.022068f
C298 VN.n61 B 0.022068f
C299 VN.n62 B 0.022068f
C300 VN.n63 B 0.027993f
C301 VN.n64 B 0.873794f
C302 VN.n65 B 0.03365f
C303 VN.n66 B 0.044007f
C304 VN.n67 B 0.022068f
C305 VN.n68 B 0.022068f
C306 VN.n69 B 0.022068f
C307 VN.n70 B 0.043137f
C308 VN.n71 B 0.035266f
C309 VN.n72 B 0.949615f
C310 VN.n73 B 1.45324f
C311 VTAIL.t9 B 0.32883f
C312 VTAIL.t4 B 0.32883f
C313 VTAIL.n0 B 2.92629f
C314 VTAIL.n1 B 0.490513f
C315 VTAIL.n2 B 0.034151f
C316 VTAIL.n3 B 0.023616f
C317 VTAIL.n4 B 0.01269f
C318 VTAIL.n5 B 0.029995f
C319 VTAIL.n6 B 0.013437f
C320 VTAIL.n7 B 0.023616f
C321 VTAIL.n8 B 0.01269f
C322 VTAIL.n9 B 0.029995f
C323 VTAIL.n10 B 0.013064f
C324 VTAIL.n11 B 0.023616f
C325 VTAIL.n12 B 0.013437f
C326 VTAIL.n13 B 0.029995f
C327 VTAIL.n14 B 0.013437f
C328 VTAIL.n15 B 0.023616f
C329 VTAIL.n16 B 0.01269f
C330 VTAIL.n17 B 0.029995f
C331 VTAIL.n18 B 0.013437f
C332 VTAIL.n19 B 0.023616f
C333 VTAIL.n20 B 0.01269f
C334 VTAIL.n21 B 0.029995f
C335 VTAIL.n22 B 0.013437f
C336 VTAIL.n23 B 0.023616f
C337 VTAIL.n24 B 0.01269f
C338 VTAIL.n25 B 0.029995f
C339 VTAIL.n26 B 0.013437f
C340 VTAIL.n27 B 0.023616f
C341 VTAIL.n28 B 0.01269f
C342 VTAIL.n29 B 0.029995f
C343 VTAIL.n30 B 0.013437f
C344 VTAIL.n31 B 1.82008f
C345 VTAIL.n32 B 0.01269f
C346 VTAIL.t15 B 0.049671f
C347 VTAIL.n33 B 0.169544f
C348 VTAIL.n34 B 0.017719f
C349 VTAIL.n35 B 0.022497f
C350 VTAIL.n36 B 0.029995f
C351 VTAIL.n37 B 0.013437f
C352 VTAIL.n38 B 0.01269f
C353 VTAIL.n39 B 0.023616f
C354 VTAIL.n40 B 0.023616f
C355 VTAIL.n41 B 0.01269f
C356 VTAIL.n42 B 0.013437f
C357 VTAIL.n43 B 0.029995f
C358 VTAIL.n44 B 0.029995f
C359 VTAIL.n45 B 0.013437f
C360 VTAIL.n46 B 0.01269f
C361 VTAIL.n47 B 0.023616f
C362 VTAIL.n48 B 0.023616f
C363 VTAIL.n49 B 0.01269f
C364 VTAIL.n50 B 0.013437f
C365 VTAIL.n51 B 0.029995f
C366 VTAIL.n52 B 0.029995f
C367 VTAIL.n53 B 0.013437f
C368 VTAIL.n54 B 0.01269f
C369 VTAIL.n55 B 0.023616f
C370 VTAIL.n56 B 0.023616f
C371 VTAIL.n57 B 0.01269f
C372 VTAIL.n58 B 0.013437f
C373 VTAIL.n59 B 0.029995f
C374 VTAIL.n60 B 0.029995f
C375 VTAIL.n61 B 0.013437f
C376 VTAIL.n62 B 0.01269f
C377 VTAIL.n63 B 0.023616f
C378 VTAIL.n64 B 0.023616f
C379 VTAIL.n65 B 0.01269f
C380 VTAIL.n66 B 0.013437f
C381 VTAIL.n67 B 0.029995f
C382 VTAIL.n68 B 0.029995f
C383 VTAIL.n69 B 0.013437f
C384 VTAIL.n70 B 0.01269f
C385 VTAIL.n71 B 0.023616f
C386 VTAIL.n72 B 0.023616f
C387 VTAIL.n73 B 0.01269f
C388 VTAIL.n74 B 0.01269f
C389 VTAIL.n75 B 0.013437f
C390 VTAIL.n76 B 0.029995f
C391 VTAIL.n77 B 0.029995f
C392 VTAIL.n78 B 0.029995f
C393 VTAIL.n79 B 0.013064f
C394 VTAIL.n80 B 0.01269f
C395 VTAIL.n81 B 0.023616f
C396 VTAIL.n82 B 0.023616f
C397 VTAIL.n83 B 0.01269f
C398 VTAIL.n84 B 0.013437f
C399 VTAIL.n85 B 0.029995f
C400 VTAIL.n86 B 0.029995f
C401 VTAIL.n87 B 0.013437f
C402 VTAIL.n88 B 0.01269f
C403 VTAIL.n89 B 0.023616f
C404 VTAIL.n90 B 0.023616f
C405 VTAIL.n91 B 0.01269f
C406 VTAIL.n92 B 0.013437f
C407 VTAIL.n93 B 0.029995f
C408 VTAIL.n94 B 0.066626f
C409 VTAIL.n95 B 0.013437f
C410 VTAIL.n96 B 0.01269f
C411 VTAIL.n97 B 0.057814f
C412 VTAIL.n98 B 0.03755f
C413 VTAIL.n99 B 0.321461f
C414 VTAIL.t17 B 0.32883f
C415 VTAIL.t14 B 0.32883f
C416 VTAIL.n100 B 2.92629f
C417 VTAIL.n101 B 0.58219f
C418 VTAIL.t10 B 0.32883f
C419 VTAIL.t19 B 0.32883f
C420 VTAIL.n102 B 2.92629f
C421 VTAIL.n103 B 2.23469f
C422 VTAIL.t7 B 0.32883f
C423 VTAIL.t0 B 0.32883f
C424 VTAIL.n104 B 2.9263f
C425 VTAIL.n105 B 2.23467f
C426 VTAIL.t6 B 0.32883f
C427 VTAIL.t8 B 0.32883f
C428 VTAIL.n106 B 2.9263f
C429 VTAIL.n107 B 0.582177f
C430 VTAIL.n108 B 0.034151f
C431 VTAIL.n109 B 0.023616f
C432 VTAIL.n110 B 0.01269f
C433 VTAIL.n111 B 0.029995f
C434 VTAIL.n112 B 0.013437f
C435 VTAIL.n113 B 0.023616f
C436 VTAIL.n114 B 0.01269f
C437 VTAIL.n115 B 0.029995f
C438 VTAIL.n116 B 0.013064f
C439 VTAIL.n117 B 0.023616f
C440 VTAIL.n118 B 0.013064f
C441 VTAIL.n119 B 0.01269f
C442 VTAIL.n120 B 0.029995f
C443 VTAIL.n121 B 0.029995f
C444 VTAIL.n122 B 0.013437f
C445 VTAIL.n123 B 0.023616f
C446 VTAIL.n124 B 0.01269f
C447 VTAIL.n125 B 0.029995f
C448 VTAIL.n126 B 0.013437f
C449 VTAIL.n127 B 0.023616f
C450 VTAIL.n128 B 0.01269f
C451 VTAIL.n129 B 0.029995f
C452 VTAIL.n130 B 0.013437f
C453 VTAIL.n131 B 0.023616f
C454 VTAIL.n132 B 0.01269f
C455 VTAIL.n133 B 0.029995f
C456 VTAIL.n134 B 0.013437f
C457 VTAIL.n135 B 0.023616f
C458 VTAIL.n136 B 0.01269f
C459 VTAIL.n137 B 0.029995f
C460 VTAIL.n138 B 0.013437f
C461 VTAIL.n139 B 1.82008f
C462 VTAIL.n140 B 0.01269f
C463 VTAIL.t3 B 0.049671f
C464 VTAIL.n141 B 0.169544f
C465 VTAIL.n142 B 0.017719f
C466 VTAIL.n143 B 0.022497f
C467 VTAIL.n144 B 0.029995f
C468 VTAIL.n145 B 0.013437f
C469 VTAIL.n146 B 0.01269f
C470 VTAIL.n147 B 0.023616f
C471 VTAIL.n148 B 0.023616f
C472 VTAIL.n149 B 0.01269f
C473 VTAIL.n150 B 0.013437f
C474 VTAIL.n151 B 0.029995f
C475 VTAIL.n152 B 0.029995f
C476 VTAIL.n153 B 0.013437f
C477 VTAIL.n154 B 0.01269f
C478 VTAIL.n155 B 0.023616f
C479 VTAIL.n156 B 0.023616f
C480 VTAIL.n157 B 0.01269f
C481 VTAIL.n158 B 0.013437f
C482 VTAIL.n159 B 0.029995f
C483 VTAIL.n160 B 0.029995f
C484 VTAIL.n161 B 0.013437f
C485 VTAIL.n162 B 0.01269f
C486 VTAIL.n163 B 0.023616f
C487 VTAIL.n164 B 0.023616f
C488 VTAIL.n165 B 0.01269f
C489 VTAIL.n166 B 0.013437f
C490 VTAIL.n167 B 0.029995f
C491 VTAIL.n168 B 0.029995f
C492 VTAIL.n169 B 0.013437f
C493 VTAIL.n170 B 0.01269f
C494 VTAIL.n171 B 0.023616f
C495 VTAIL.n172 B 0.023616f
C496 VTAIL.n173 B 0.01269f
C497 VTAIL.n174 B 0.013437f
C498 VTAIL.n175 B 0.029995f
C499 VTAIL.n176 B 0.029995f
C500 VTAIL.n177 B 0.013437f
C501 VTAIL.n178 B 0.01269f
C502 VTAIL.n179 B 0.023616f
C503 VTAIL.n180 B 0.023616f
C504 VTAIL.n181 B 0.01269f
C505 VTAIL.n182 B 0.013437f
C506 VTAIL.n183 B 0.029995f
C507 VTAIL.n184 B 0.029995f
C508 VTAIL.n185 B 0.013437f
C509 VTAIL.n186 B 0.01269f
C510 VTAIL.n187 B 0.023616f
C511 VTAIL.n188 B 0.023616f
C512 VTAIL.n189 B 0.01269f
C513 VTAIL.n190 B 0.013437f
C514 VTAIL.n191 B 0.029995f
C515 VTAIL.n192 B 0.029995f
C516 VTAIL.n193 B 0.013437f
C517 VTAIL.n194 B 0.01269f
C518 VTAIL.n195 B 0.023616f
C519 VTAIL.n196 B 0.023616f
C520 VTAIL.n197 B 0.01269f
C521 VTAIL.n198 B 0.013437f
C522 VTAIL.n199 B 0.029995f
C523 VTAIL.n200 B 0.066626f
C524 VTAIL.n201 B 0.013437f
C525 VTAIL.n202 B 0.01269f
C526 VTAIL.n203 B 0.057814f
C527 VTAIL.n204 B 0.03755f
C528 VTAIL.n205 B 0.321461f
C529 VTAIL.t12 B 0.32883f
C530 VTAIL.t13 B 0.32883f
C531 VTAIL.n206 B 2.9263f
C532 VTAIL.n207 B 0.530024f
C533 VTAIL.t16 B 0.32883f
C534 VTAIL.t18 B 0.32883f
C535 VTAIL.n208 B 2.9263f
C536 VTAIL.n209 B 0.582177f
C537 VTAIL.n210 B 0.034151f
C538 VTAIL.n211 B 0.023616f
C539 VTAIL.n212 B 0.01269f
C540 VTAIL.n213 B 0.029995f
C541 VTAIL.n214 B 0.013437f
C542 VTAIL.n215 B 0.023616f
C543 VTAIL.n216 B 0.01269f
C544 VTAIL.n217 B 0.029995f
C545 VTAIL.n218 B 0.013064f
C546 VTAIL.n219 B 0.023616f
C547 VTAIL.n220 B 0.013064f
C548 VTAIL.n221 B 0.01269f
C549 VTAIL.n222 B 0.029995f
C550 VTAIL.n223 B 0.029995f
C551 VTAIL.n224 B 0.013437f
C552 VTAIL.n225 B 0.023616f
C553 VTAIL.n226 B 0.01269f
C554 VTAIL.n227 B 0.029995f
C555 VTAIL.n228 B 0.013437f
C556 VTAIL.n229 B 0.023616f
C557 VTAIL.n230 B 0.01269f
C558 VTAIL.n231 B 0.029995f
C559 VTAIL.n232 B 0.013437f
C560 VTAIL.n233 B 0.023616f
C561 VTAIL.n234 B 0.01269f
C562 VTAIL.n235 B 0.029995f
C563 VTAIL.n236 B 0.013437f
C564 VTAIL.n237 B 0.023616f
C565 VTAIL.n238 B 0.01269f
C566 VTAIL.n239 B 0.029995f
C567 VTAIL.n240 B 0.013437f
C568 VTAIL.n241 B 1.82008f
C569 VTAIL.n242 B 0.01269f
C570 VTAIL.t11 B 0.049671f
C571 VTAIL.n243 B 0.169544f
C572 VTAIL.n244 B 0.017719f
C573 VTAIL.n245 B 0.022497f
C574 VTAIL.n246 B 0.029995f
C575 VTAIL.n247 B 0.013437f
C576 VTAIL.n248 B 0.01269f
C577 VTAIL.n249 B 0.023616f
C578 VTAIL.n250 B 0.023616f
C579 VTAIL.n251 B 0.01269f
C580 VTAIL.n252 B 0.013437f
C581 VTAIL.n253 B 0.029995f
C582 VTAIL.n254 B 0.029995f
C583 VTAIL.n255 B 0.013437f
C584 VTAIL.n256 B 0.01269f
C585 VTAIL.n257 B 0.023616f
C586 VTAIL.n258 B 0.023616f
C587 VTAIL.n259 B 0.01269f
C588 VTAIL.n260 B 0.013437f
C589 VTAIL.n261 B 0.029995f
C590 VTAIL.n262 B 0.029995f
C591 VTAIL.n263 B 0.013437f
C592 VTAIL.n264 B 0.01269f
C593 VTAIL.n265 B 0.023616f
C594 VTAIL.n266 B 0.023616f
C595 VTAIL.n267 B 0.01269f
C596 VTAIL.n268 B 0.013437f
C597 VTAIL.n269 B 0.029995f
C598 VTAIL.n270 B 0.029995f
C599 VTAIL.n271 B 0.013437f
C600 VTAIL.n272 B 0.01269f
C601 VTAIL.n273 B 0.023616f
C602 VTAIL.n274 B 0.023616f
C603 VTAIL.n275 B 0.01269f
C604 VTAIL.n276 B 0.013437f
C605 VTAIL.n277 B 0.029995f
C606 VTAIL.n278 B 0.029995f
C607 VTAIL.n279 B 0.013437f
C608 VTAIL.n280 B 0.01269f
C609 VTAIL.n281 B 0.023616f
C610 VTAIL.n282 B 0.023616f
C611 VTAIL.n283 B 0.01269f
C612 VTAIL.n284 B 0.013437f
C613 VTAIL.n285 B 0.029995f
C614 VTAIL.n286 B 0.029995f
C615 VTAIL.n287 B 0.013437f
C616 VTAIL.n288 B 0.01269f
C617 VTAIL.n289 B 0.023616f
C618 VTAIL.n290 B 0.023616f
C619 VTAIL.n291 B 0.01269f
C620 VTAIL.n292 B 0.013437f
C621 VTAIL.n293 B 0.029995f
C622 VTAIL.n294 B 0.029995f
C623 VTAIL.n295 B 0.013437f
C624 VTAIL.n296 B 0.01269f
C625 VTAIL.n297 B 0.023616f
C626 VTAIL.n298 B 0.023616f
C627 VTAIL.n299 B 0.01269f
C628 VTAIL.n300 B 0.013437f
C629 VTAIL.n301 B 0.029995f
C630 VTAIL.n302 B 0.066626f
C631 VTAIL.n303 B 0.013437f
C632 VTAIL.n304 B 0.01269f
C633 VTAIL.n305 B 0.057814f
C634 VTAIL.n306 B 0.03755f
C635 VTAIL.n307 B 1.8503f
C636 VTAIL.n308 B 0.034151f
C637 VTAIL.n309 B 0.023616f
C638 VTAIL.n310 B 0.01269f
C639 VTAIL.n311 B 0.029995f
C640 VTAIL.n312 B 0.013437f
C641 VTAIL.n313 B 0.023616f
C642 VTAIL.n314 B 0.01269f
C643 VTAIL.n315 B 0.029995f
C644 VTAIL.n316 B 0.013064f
C645 VTAIL.n317 B 0.023616f
C646 VTAIL.n318 B 0.013437f
C647 VTAIL.n319 B 0.029995f
C648 VTAIL.n320 B 0.013437f
C649 VTAIL.n321 B 0.023616f
C650 VTAIL.n322 B 0.01269f
C651 VTAIL.n323 B 0.029995f
C652 VTAIL.n324 B 0.013437f
C653 VTAIL.n325 B 0.023616f
C654 VTAIL.n326 B 0.01269f
C655 VTAIL.n327 B 0.029995f
C656 VTAIL.n328 B 0.013437f
C657 VTAIL.n329 B 0.023616f
C658 VTAIL.n330 B 0.01269f
C659 VTAIL.n331 B 0.029995f
C660 VTAIL.n332 B 0.013437f
C661 VTAIL.n333 B 0.023616f
C662 VTAIL.n334 B 0.01269f
C663 VTAIL.n335 B 0.029995f
C664 VTAIL.n336 B 0.013437f
C665 VTAIL.n337 B 1.82008f
C666 VTAIL.n338 B 0.01269f
C667 VTAIL.t2 B 0.049671f
C668 VTAIL.n339 B 0.169544f
C669 VTAIL.n340 B 0.017719f
C670 VTAIL.n341 B 0.022497f
C671 VTAIL.n342 B 0.029995f
C672 VTAIL.n343 B 0.013437f
C673 VTAIL.n344 B 0.01269f
C674 VTAIL.n345 B 0.023616f
C675 VTAIL.n346 B 0.023616f
C676 VTAIL.n347 B 0.01269f
C677 VTAIL.n348 B 0.013437f
C678 VTAIL.n349 B 0.029995f
C679 VTAIL.n350 B 0.029995f
C680 VTAIL.n351 B 0.013437f
C681 VTAIL.n352 B 0.01269f
C682 VTAIL.n353 B 0.023616f
C683 VTAIL.n354 B 0.023616f
C684 VTAIL.n355 B 0.01269f
C685 VTAIL.n356 B 0.013437f
C686 VTAIL.n357 B 0.029995f
C687 VTAIL.n358 B 0.029995f
C688 VTAIL.n359 B 0.013437f
C689 VTAIL.n360 B 0.01269f
C690 VTAIL.n361 B 0.023616f
C691 VTAIL.n362 B 0.023616f
C692 VTAIL.n363 B 0.01269f
C693 VTAIL.n364 B 0.013437f
C694 VTAIL.n365 B 0.029995f
C695 VTAIL.n366 B 0.029995f
C696 VTAIL.n367 B 0.013437f
C697 VTAIL.n368 B 0.01269f
C698 VTAIL.n369 B 0.023616f
C699 VTAIL.n370 B 0.023616f
C700 VTAIL.n371 B 0.01269f
C701 VTAIL.n372 B 0.013437f
C702 VTAIL.n373 B 0.029995f
C703 VTAIL.n374 B 0.029995f
C704 VTAIL.n375 B 0.013437f
C705 VTAIL.n376 B 0.01269f
C706 VTAIL.n377 B 0.023616f
C707 VTAIL.n378 B 0.023616f
C708 VTAIL.n379 B 0.01269f
C709 VTAIL.n380 B 0.01269f
C710 VTAIL.n381 B 0.013437f
C711 VTAIL.n382 B 0.029995f
C712 VTAIL.n383 B 0.029995f
C713 VTAIL.n384 B 0.029995f
C714 VTAIL.n385 B 0.013064f
C715 VTAIL.n386 B 0.01269f
C716 VTAIL.n387 B 0.023616f
C717 VTAIL.n388 B 0.023616f
C718 VTAIL.n389 B 0.01269f
C719 VTAIL.n390 B 0.013437f
C720 VTAIL.n391 B 0.029995f
C721 VTAIL.n392 B 0.029995f
C722 VTAIL.n393 B 0.013437f
C723 VTAIL.n394 B 0.01269f
C724 VTAIL.n395 B 0.023616f
C725 VTAIL.n396 B 0.023616f
C726 VTAIL.n397 B 0.01269f
C727 VTAIL.n398 B 0.013437f
C728 VTAIL.n399 B 0.029995f
C729 VTAIL.n400 B 0.066626f
C730 VTAIL.n401 B 0.013437f
C731 VTAIL.n402 B 0.01269f
C732 VTAIL.n403 B 0.057814f
C733 VTAIL.n404 B 0.03755f
C734 VTAIL.n405 B 1.8503f
C735 VTAIL.t1 B 0.32883f
C736 VTAIL.t5 B 0.32883f
C737 VTAIL.n406 B 2.92629f
C738 VTAIL.n407 B 0.445904f
C739 VDD1.n0 B 0.034218f
C740 VDD1.n1 B 0.023663f
C741 VDD1.n2 B 0.012715f
C742 VDD1.n3 B 0.030055f
C743 VDD1.n4 B 0.013463f
C744 VDD1.n5 B 0.023663f
C745 VDD1.n6 B 0.012715f
C746 VDD1.n7 B 0.030055f
C747 VDD1.n8 B 0.013089f
C748 VDD1.n9 B 0.023663f
C749 VDD1.n10 B 0.013089f
C750 VDD1.n11 B 0.012715f
C751 VDD1.n12 B 0.030055f
C752 VDD1.n13 B 0.030055f
C753 VDD1.n14 B 0.013463f
C754 VDD1.n15 B 0.023663f
C755 VDD1.n16 B 0.012715f
C756 VDD1.n17 B 0.030055f
C757 VDD1.n18 B 0.013463f
C758 VDD1.n19 B 0.023663f
C759 VDD1.n20 B 0.012715f
C760 VDD1.n21 B 0.030055f
C761 VDD1.n22 B 0.013463f
C762 VDD1.n23 B 0.023663f
C763 VDD1.n24 B 0.012715f
C764 VDD1.n25 B 0.030055f
C765 VDD1.n26 B 0.013463f
C766 VDD1.n27 B 0.023663f
C767 VDD1.n28 B 0.012715f
C768 VDD1.n29 B 0.030055f
C769 VDD1.n30 B 0.013463f
C770 VDD1.n31 B 1.82368f
C771 VDD1.n32 B 0.012715f
C772 VDD1.t2 B 0.049769f
C773 VDD1.n33 B 0.169879f
C774 VDD1.n34 B 0.017754f
C775 VDD1.n35 B 0.022541f
C776 VDD1.n36 B 0.030055f
C777 VDD1.n37 B 0.013463f
C778 VDD1.n38 B 0.012715f
C779 VDD1.n39 B 0.023663f
C780 VDD1.n40 B 0.023663f
C781 VDD1.n41 B 0.012715f
C782 VDD1.n42 B 0.013463f
C783 VDD1.n43 B 0.030055f
C784 VDD1.n44 B 0.030055f
C785 VDD1.n45 B 0.013463f
C786 VDD1.n46 B 0.012715f
C787 VDD1.n47 B 0.023663f
C788 VDD1.n48 B 0.023663f
C789 VDD1.n49 B 0.012715f
C790 VDD1.n50 B 0.013463f
C791 VDD1.n51 B 0.030055f
C792 VDD1.n52 B 0.030055f
C793 VDD1.n53 B 0.013463f
C794 VDD1.n54 B 0.012715f
C795 VDD1.n55 B 0.023663f
C796 VDD1.n56 B 0.023663f
C797 VDD1.n57 B 0.012715f
C798 VDD1.n58 B 0.013463f
C799 VDD1.n59 B 0.030055f
C800 VDD1.n60 B 0.030055f
C801 VDD1.n61 B 0.013463f
C802 VDD1.n62 B 0.012715f
C803 VDD1.n63 B 0.023663f
C804 VDD1.n64 B 0.023663f
C805 VDD1.n65 B 0.012715f
C806 VDD1.n66 B 0.013463f
C807 VDD1.n67 B 0.030055f
C808 VDD1.n68 B 0.030055f
C809 VDD1.n69 B 0.013463f
C810 VDD1.n70 B 0.012715f
C811 VDD1.n71 B 0.023663f
C812 VDD1.n72 B 0.023663f
C813 VDD1.n73 B 0.012715f
C814 VDD1.n74 B 0.013463f
C815 VDD1.n75 B 0.030055f
C816 VDD1.n76 B 0.030055f
C817 VDD1.n77 B 0.013463f
C818 VDD1.n78 B 0.012715f
C819 VDD1.n79 B 0.023663f
C820 VDD1.n80 B 0.023663f
C821 VDD1.n81 B 0.012715f
C822 VDD1.n82 B 0.013463f
C823 VDD1.n83 B 0.030055f
C824 VDD1.n84 B 0.030055f
C825 VDD1.n85 B 0.013463f
C826 VDD1.n86 B 0.012715f
C827 VDD1.n87 B 0.023663f
C828 VDD1.n88 B 0.023663f
C829 VDD1.n89 B 0.012715f
C830 VDD1.n90 B 0.013463f
C831 VDD1.n91 B 0.030055f
C832 VDD1.n92 B 0.066757f
C833 VDD1.n93 B 0.013463f
C834 VDD1.n94 B 0.012715f
C835 VDD1.n95 B 0.057928f
C836 VDD1.n96 B 0.063664f
C837 VDD1.t3 B 0.32948f
C838 VDD1.t4 B 0.32948f
C839 VDD1.n97 B 3.00098f
C840 VDD1.n98 B 0.632762f
C841 VDD1.n99 B 0.034218f
C842 VDD1.n100 B 0.023663f
C843 VDD1.n101 B 0.012715f
C844 VDD1.n102 B 0.030055f
C845 VDD1.n103 B 0.013463f
C846 VDD1.n104 B 0.023663f
C847 VDD1.n105 B 0.012715f
C848 VDD1.n106 B 0.030055f
C849 VDD1.n107 B 0.013089f
C850 VDD1.n108 B 0.023663f
C851 VDD1.n109 B 0.013463f
C852 VDD1.n110 B 0.030055f
C853 VDD1.n111 B 0.013463f
C854 VDD1.n112 B 0.023663f
C855 VDD1.n113 B 0.012715f
C856 VDD1.n114 B 0.030055f
C857 VDD1.n115 B 0.013463f
C858 VDD1.n116 B 0.023663f
C859 VDD1.n117 B 0.012715f
C860 VDD1.n118 B 0.030055f
C861 VDD1.n119 B 0.013463f
C862 VDD1.n120 B 0.023663f
C863 VDD1.n121 B 0.012715f
C864 VDD1.n122 B 0.030055f
C865 VDD1.n123 B 0.013463f
C866 VDD1.n124 B 0.023663f
C867 VDD1.n125 B 0.012715f
C868 VDD1.n126 B 0.030055f
C869 VDD1.n127 B 0.013463f
C870 VDD1.n128 B 1.82368f
C871 VDD1.n129 B 0.012715f
C872 VDD1.t6 B 0.049769f
C873 VDD1.n130 B 0.169879f
C874 VDD1.n131 B 0.017754f
C875 VDD1.n132 B 0.022541f
C876 VDD1.n133 B 0.030055f
C877 VDD1.n134 B 0.013463f
C878 VDD1.n135 B 0.012715f
C879 VDD1.n136 B 0.023663f
C880 VDD1.n137 B 0.023663f
C881 VDD1.n138 B 0.012715f
C882 VDD1.n139 B 0.013463f
C883 VDD1.n140 B 0.030055f
C884 VDD1.n141 B 0.030055f
C885 VDD1.n142 B 0.013463f
C886 VDD1.n143 B 0.012715f
C887 VDD1.n144 B 0.023663f
C888 VDD1.n145 B 0.023663f
C889 VDD1.n146 B 0.012715f
C890 VDD1.n147 B 0.013463f
C891 VDD1.n148 B 0.030055f
C892 VDD1.n149 B 0.030055f
C893 VDD1.n150 B 0.013463f
C894 VDD1.n151 B 0.012715f
C895 VDD1.n152 B 0.023663f
C896 VDD1.n153 B 0.023663f
C897 VDD1.n154 B 0.012715f
C898 VDD1.n155 B 0.013463f
C899 VDD1.n156 B 0.030055f
C900 VDD1.n157 B 0.030055f
C901 VDD1.n158 B 0.013463f
C902 VDD1.n159 B 0.012715f
C903 VDD1.n160 B 0.023663f
C904 VDD1.n161 B 0.023663f
C905 VDD1.n162 B 0.012715f
C906 VDD1.n163 B 0.013463f
C907 VDD1.n164 B 0.030055f
C908 VDD1.n165 B 0.030055f
C909 VDD1.n166 B 0.013463f
C910 VDD1.n167 B 0.012715f
C911 VDD1.n168 B 0.023663f
C912 VDD1.n169 B 0.023663f
C913 VDD1.n170 B 0.012715f
C914 VDD1.n171 B 0.012715f
C915 VDD1.n172 B 0.013463f
C916 VDD1.n173 B 0.030055f
C917 VDD1.n174 B 0.030055f
C918 VDD1.n175 B 0.030055f
C919 VDD1.n176 B 0.013089f
C920 VDD1.n177 B 0.012715f
C921 VDD1.n178 B 0.023663f
C922 VDD1.n179 B 0.023663f
C923 VDD1.n180 B 0.012715f
C924 VDD1.n181 B 0.013463f
C925 VDD1.n182 B 0.030055f
C926 VDD1.n183 B 0.030055f
C927 VDD1.n184 B 0.013463f
C928 VDD1.n185 B 0.012715f
C929 VDD1.n186 B 0.023663f
C930 VDD1.n187 B 0.023663f
C931 VDD1.n188 B 0.012715f
C932 VDD1.n189 B 0.013463f
C933 VDD1.n190 B 0.030055f
C934 VDD1.n191 B 0.066757f
C935 VDD1.n192 B 0.013463f
C936 VDD1.n193 B 0.012715f
C937 VDD1.n194 B 0.057928f
C938 VDD1.n195 B 0.063664f
C939 VDD1.t9 B 0.32948f
C940 VDD1.t5 B 0.32948f
C941 VDD1.n196 B 3.00097f
C942 VDD1.n197 B 0.625164f
C943 VDD1.t0 B 0.32948f
C944 VDD1.t1 B 0.32948f
C945 VDD1.n198 B 3.01423f
C946 VDD1.n199 B 3.07332f
C947 VDD1.t8 B 0.32948f
C948 VDD1.t7 B 0.32948f
C949 VDD1.n200 B 3.00097f
C950 VDD1.n201 B 3.30825f
C951 VP.n0 B 0.029409f
C952 VP.t4 B 2.5397f
C953 VP.n1 B 0.018132f
C954 VP.n2 B 0.022308f
C955 VP.t5 B 2.5397f
C956 VP.n3 B 0.041755f
C957 VP.n4 B 0.022308f
C958 VP.t2 B 2.5397f
C959 VP.n5 B 0.904258f
C960 VP.n6 B 0.022308f
C961 VP.n7 B 0.041755f
C962 VP.n8 B 0.022308f
C963 VP.t0 B 2.5397f
C964 VP.n9 B 0.018132f
C965 VP.n10 B 0.029409f
C966 VP.t9 B 2.5397f
C967 VP.n11 B 0.029409f
C968 VP.t8 B 2.5397f
C969 VP.n12 B 0.018132f
C970 VP.n13 B 0.022308f
C971 VP.t1 B 2.5397f
C972 VP.n14 B 0.041755f
C973 VP.n15 B 0.022308f
C974 VP.t3 B 2.5397f
C975 VP.n16 B 0.904258f
C976 VP.n17 B 0.022308f
C977 VP.n18 B 0.041755f
C978 VP.t7 B 2.69743f
C979 VP.n19 B 0.928986f
C980 VP.t6 B 2.5397f
C981 VP.n20 B 0.940345f
C982 VP.n21 B 0.028298f
C983 VP.n22 B 0.193063f
C984 VP.n23 B 0.022308f
C985 VP.n24 B 0.022308f
C986 VP.n25 B 0.026541f
C987 VP.n26 B 0.037928f
C988 VP.n27 B 0.041368f
C989 VP.n28 B 0.022308f
C990 VP.n29 B 0.022308f
C991 VP.n30 B 0.022308f
C992 VP.n31 B 0.041368f
C993 VP.n32 B 0.037928f
C994 VP.n33 B 0.026541f
C995 VP.n34 B 0.022308f
C996 VP.n35 B 0.022308f
C997 VP.n36 B 0.022308f
C998 VP.n37 B 0.028298f
C999 VP.n38 B 0.883312f
C1000 VP.n39 B 0.034016f
C1001 VP.n40 B 0.044487f
C1002 VP.n41 B 0.022308f
C1003 VP.n42 B 0.022308f
C1004 VP.n43 B 0.022308f
C1005 VP.n44 B 0.043607f
C1006 VP.n45 B 0.03565f
C1007 VP.n46 B 0.959959f
C1008 VP.n47 B 1.45729f
C1009 VP.n48 B 1.47163f
C1010 VP.n49 B 0.959959f
C1011 VP.n50 B 0.03565f
C1012 VP.n51 B 0.043607f
C1013 VP.n52 B 0.022308f
C1014 VP.n53 B 0.022308f
C1015 VP.n54 B 0.022308f
C1016 VP.n55 B 0.044487f
C1017 VP.n56 B 0.034016f
C1018 VP.n57 B 0.883312f
C1019 VP.n58 B 0.028298f
C1020 VP.n59 B 0.022308f
C1021 VP.n60 B 0.022308f
C1022 VP.n61 B 0.022308f
C1023 VP.n62 B 0.026541f
C1024 VP.n63 B 0.037928f
C1025 VP.n64 B 0.041368f
C1026 VP.n65 B 0.022308f
C1027 VP.n66 B 0.022308f
C1028 VP.n67 B 0.022308f
C1029 VP.n68 B 0.041368f
C1030 VP.n69 B 0.037928f
C1031 VP.n70 B 0.026541f
C1032 VP.n71 B 0.022308f
C1033 VP.n72 B 0.022308f
C1034 VP.n73 B 0.022308f
C1035 VP.n74 B 0.028298f
C1036 VP.n75 B 0.883312f
C1037 VP.n76 B 0.034016f
C1038 VP.n77 B 0.044487f
C1039 VP.n78 B 0.022308f
C1040 VP.n79 B 0.022308f
C1041 VP.n80 B 0.022308f
C1042 VP.n81 B 0.043607f
C1043 VP.n82 B 0.03565f
C1044 VP.n83 B 0.959959f
C1045 VP.n84 B 0.029959f
.ends

