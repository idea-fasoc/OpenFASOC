* NGSPICE file created from diff_pair_sample_0833.ext - technology: sky130A

.subckt diff_pair_sample_0833 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X1 VDD1.t9 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=0 ps=0 w=18.37 l=0.32
X3 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=0 ps=0 w=18.37 l=0.32
X4 VTAIL.t5 VP.t1 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X5 VDD2.t7 VN.t1 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=3.03105 ps=18.7 w=18.37 l=0.32
X6 VDD1.t7 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=7.1643 ps=37.52 w=18.37 l=0.32
X7 VTAIL.t14 VN.t2 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X8 VDD2.t2 VN.t3 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=7.1643 ps=37.52 w=18.37 l=0.32
X9 VDD1.t6 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=3.03105 ps=18.7 w=18.37 l=0.32
X10 VDD2.t1 VN.t4 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=3.03105 ps=18.7 w=18.37 l=0.32
X11 VDD2.t4 VN.t5 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=7.1643 ps=37.52 w=18.37 l=0.32
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=0 ps=0 w=18.37 l=0.32
X13 VTAIL.t10 VN.t6 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X14 VTAIL.t9 VN.t7 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X15 VTAIL.t4 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X16 VTAIL.t0 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X17 VDD2.t8 VN.t8 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X18 VDD1.t3 VP.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X19 VDD2.t5 VN.t9 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=0 ps=0 w=18.37 l=0.32
X21 VTAIL.t17 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=3.03105 ps=18.7 w=18.37 l=0.32
X22 VDD1.t1 VP.t8 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=3.03105 pd=18.7 as=7.1643 ps=37.52 w=18.37 l=0.32
X23 VDD1.t0 VP.t9 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1643 pd=37.52 as=3.03105 ps=18.7 w=18.37 l=0.32
R0 VN.n9 VN.t3 1525.97
R1 VN.n3 VN.t1 1525.97
R2 VN.n20 VN.t4 1525.97
R3 VN.n14 VN.t5 1525.97
R4 VN.n6 VN.t9 1482.15
R5 VN.n8 VN.t0 1482.15
R6 VN.n2 VN.t6 1482.15
R7 VN.n17 VN.t8 1482.15
R8 VN.n19 VN.t7 1482.15
R9 VN.n13 VN.t2 1482.15
R10 VN.n15 VN.n14 161.489
R11 VN.n4 VN.n3 161.489
R12 VN.n10 VN.n9 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n18 VN.n11 161.3
R15 VN.n17 VN.n16 161.3
R16 VN.n15 VN.n12 161.3
R17 VN.n7 VN.n0 161.3
R18 VN.n6 VN.n5 161.3
R19 VN.n4 VN.n1 161.3
R20 VN.n6 VN.n1 73.0308
R21 VN.n7 VN.n6 73.0308
R22 VN.n18 VN.n17 73.0308
R23 VN.n17 VN.n12 73.0308
R24 VN.n3 VN.n2 51.1217
R25 VN.n9 VN.n8 51.1217
R26 VN.n20 VN.n19 51.1217
R27 VN.n14 VN.n13 51.1217
R28 VN VN.n21 46.0138
R29 VN.n2 VN.n1 21.9096
R30 VN.n8 VN.n7 21.9096
R31 VN.n19 VN.n18 21.9096
R32 VN.n13 VN.n12 21.9096
R33 VN.n21 VN.n11 0.189894
R34 VN.n16 VN.n11 0.189894
R35 VN.n16 VN.n15 0.189894
R36 VN.n5 VN.n4 0.189894
R37 VN.n5 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VDD2.n1 VDD2.t7 64.2962
R41 VDD2.n4 VDD2.t1 63.7368
R42 VDD2.n3 VDD2.n2 63.0237
R43 VDD2 VDD2.n7 63.02
R44 VDD2.n6 VDD2.n5 62.659
R45 VDD2.n1 VDD2.n0 62.6588
R46 VDD2.n4 VDD2.n3 42.2131
R47 VDD2.n7 VDD2.t6 1.07834
R48 VDD2.n7 VDD2.t4 1.07834
R49 VDD2.n5 VDD2.t9 1.07834
R50 VDD2.n5 VDD2.t8 1.07834
R51 VDD2.n2 VDD2.t0 1.07834
R52 VDD2.n2 VDD2.t2 1.07834
R53 VDD2.n0 VDD2.t3 1.07834
R54 VDD2.n0 VDD2.t5 1.07834
R55 VDD2.n6 VDD2.n4 0.560845
R56 VDD2 VDD2.n6 0.198776
R57 VDD2.n3 VDD2.n1 0.0852402
R58 VTAIL.n11 VTAIL.t11 47.0581
R59 VTAIL.n17 VTAIL.t13 47.057
R60 VTAIL.n2 VTAIL.t1 47.057
R61 VTAIL.n16 VTAIL.t18 47.057
R62 VTAIL.n15 VTAIL.n14 45.9802
R63 VTAIL.n13 VTAIL.n12 45.9802
R64 VTAIL.n10 VTAIL.n9 45.9802
R65 VTAIL.n8 VTAIL.n7 45.9802
R66 VTAIL.n19 VTAIL.n18 45.98
R67 VTAIL.n1 VTAIL.n0 45.98
R68 VTAIL.n4 VTAIL.n3 45.98
R69 VTAIL.n6 VTAIL.n5 45.98
R70 VTAIL.n8 VTAIL.n6 29.3238
R71 VTAIL.n17 VTAIL.n16 28.7634
R72 VTAIL.n18 VTAIL.t7 1.07834
R73 VTAIL.n18 VTAIL.t16 1.07834
R74 VTAIL.n0 VTAIL.t15 1.07834
R75 VTAIL.n0 VTAIL.t10 1.07834
R76 VTAIL.n3 VTAIL.t6 1.07834
R77 VTAIL.n3 VTAIL.t4 1.07834
R78 VTAIL.n5 VTAIL.t3 1.07834
R79 VTAIL.n5 VTAIL.t5 1.07834
R80 VTAIL.n14 VTAIL.t2 1.07834
R81 VTAIL.n14 VTAIL.t0 1.07834
R82 VTAIL.n12 VTAIL.t19 1.07834
R83 VTAIL.n12 VTAIL.t17 1.07834
R84 VTAIL.n9 VTAIL.t8 1.07834
R85 VTAIL.n9 VTAIL.t14 1.07834
R86 VTAIL.n7 VTAIL.t12 1.07834
R87 VTAIL.n7 VTAIL.t9 1.07834
R88 VTAIL.n13 VTAIL.n11 0.7505
R89 VTAIL.n2 VTAIL.n1 0.7505
R90 VTAIL.n10 VTAIL.n8 0.560845
R91 VTAIL.n11 VTAIL.n10 0.560845
R92 VTAIL.n15 VTAIL.n13 0.560845
R93 VTAIL.n16 VTAIL.n15 0.560845
R94 VTAIL.n6 VTAIL.n4 0.560845
R95 VTAIL.n4 VTAIL.n2 0.560845
R96 VTAIL.n19 VTAIL.n17 0.560845
R97 VTAIL VTAIL.n1 0.478948
R98 VTAIL VTAIL.n19 0.0823966
R99 B.n108 B.t21 1597.25
R100 B.n105 B.t14 1597.25
R101 B.n467 B.t10 1597.25
R102 B.n465 B.t18 1597.25
R103 B.n815 B.n814 585
R104 B.n363 B.n103 585
R105 B.n362 B.n361 585
R106 B.n360 B.n359 585
R107 B.n358 B.n357 585
R108 B.n356 B.n355 585
R109 B.n354 B.n353 585
R110 B.n352 B.n351 585
R111 B.n350 B.n349 585
R112 B.n348 B.n347 585
R113 B.n346 B.n345 585
R114 B.n344 B.n343 585
R115 B.n342 B.n341 585
R116 B.n340 B.n339 585
R117 B.n338 B.n337 585
R118 B.n336 B.n335 585
R119 B.n334 B.n333 585
R120 B.n332 B.n331 585
R121 B.n330 B.n329 585
R122 B.n328 B.n327 585
R123 B.n326 B.n325 585
R124 B.n324 B.n323 585
R125 B.n322 B.n321 585
R126 B.n320 B.n319 585
R127 B.n318 B.n317 585
R128 B.n316 B.n315 585
R129 B.n314 B.n313 585
R130 B.n312 B.n311 585
R131 B.n310 B.n309 585
R132 B.n308 B.n307 585
R133 B.n306 B.n305 585
R134 B.n304 B.n303 585
R135 B.n302 B.n301 585
R136 B.n300 B.n299 585
R137 B.n298 B.n297 585
R138 B.n296 B.n295 585
R139 B.n294 B.n293 585
R140 B.n292 B.n291 585
R141 B.n290 B.n289 585
R142 B.n288 B.n287 585
R143 B.n286 B.n285 585
R144 B.n284 B.n283 585
R145 B.n282 B.n281 585
R146 B.n280 B.n279 585
R147 B.n278 B.n277 585
R148 B.n276 B.n275 585
R149 B.n274 B.n273 585
R150 B.n272 B.n271 585
R151 B.n270 B.n269 585
R152 B.n268 B.n267 585
R153 B.n266 B.n265 585
R154 B.n264 B.n263 585
R155 B.n262 B.n261 585
R156 B.n260 B.n259 585
R157 B.n258 B.n257 585
R158 B.n256 B.n255 585
R159 B.n254 B.n253 585
R160 B.n252 B.n251 585
R161 B.n250 B.n249 585
R162 B.n248 B.n247 585
R163 B.n246 B.n245 585
R164 B.n244 B.n243 585
R165 B.n242 B.n241 585
R166 B.n240 B.n239 585
R167 B.n238 B.n237 585
R168 B.n236 B.n235 585
R169 B.n234 B.n233 585
R170 B.n232 B.n231 585
R171 B.n230 B.n229 585
R172 B.n228 B.n227 585
R173 B.n226 B.n225 585
R174 B.n224 B.n223 585
R175 B.n222 B.n221 585
R176 B.n220 B.n219 585
R177 B.n218 B.n217 585
R178 B.n216 B.n215 585
R179 B.n214 B.n213 585
R180 B.n212 B.n211 585
R181 B.n210 B.n209 585
R182 B.n208 B.n207 585
R183 B.n206 B.n205 585
R184 B.n204 B.n203 585
R185 B.n202 B.n201 585
R186 B.n200 B.n199 585
R187 B.n198 B.n197 585
R188 B.n196 B.n195 585
R189 B.n194 B.n193 585
R190 B.n192 B.n191 585
R191 B.n190 B.n189 585
R192 B.n188 B.n187 585
R193 B.n186 B.n185 585
R194 B.n184 B.n183 585
R195 B.n182 B.n181 585
R196 B.n180 B.n179 585
R197 B.n178 B.n177 585
R198 B.n176 B.n175 585
R199 B.n174 B.n173 585
R200 B.n172 B.n171 585
R201 B.n170 B.n169 585
R202 B.n168 B.n167 585
R203 B.n166 B.n165 585
R204 B.n164 B.n163 585
R205 B.n162 B.n161 585
R206 B.n160 B.n159 585
R207 B.n158 B.n157 585
R208 B.n156 B.n155 585
R209 B.n154 B.n153 585
R210 B.n152 B.n151 585
R211 B.n150 B.n149 585
R212 B.n148 B.n147 585
R213 B.n146 B.n145 585
R214 B.n144 B.n143 585
R215 B.n142 B.n141 585
R216 B.n140 B.n139 585
R217 B.n138 B.n137 585
R218 B.n136 B.n135 585
R219 B.n134 B.n133 585
R220 B.n132 B.n131 585
R221 B.n130 B.n129 585
R222 B.n128 B.n127 585
R223 B.n126 B.n125 585
R224 B.n124 B.n123 585
R225 B.n122 B.n121 585
R226 B.n120 B.n119 585
R227 B.n118 B.n117 585
R228 B.n116 B.n115 585
R229 B.n114 B.n113 585
R230 B.n112 B.n111 585
R231 B.n39 B.n38 585
R232 B.n820 B.n819 585
R233 B.n813 B.n104 585
R234 B.n104 B.n36 585
R235 B.n812 B.n35 585
R236 B.n824 B.n35 585
R237 B.n811 B.n34 585
R238 B.n825 B.n34 585
R239 B.n810 B.n33 585
R240 B.n826 B.n33 585
R241 B.n809 B.n808 585
R242 B.n808 B.n32 585
R243 B.n807 B.n28 585
R244 B.n832 B.n28 585
R245 B.n806 B.n27 585
R246 B.n833 B.n27 585
R247 B.n805 B.n26 585
R248 B.n834 B.n26 585
R249 B.n804 B.n803 585
R250 B.n803 B.n22 585
R251 B.n802 B.n21 585
R252 B.n840 B.n21 585
R253 B.n801 B.n20 585
R254 B.n841 B.n20 585
R255 B.n800 B.n19 585
R256 B.n842 B.n19 585
R257 B.n799 B.n798 585
R258 B.n798 B.n15 585
R259 B.n797 B.n14 585
R260 B.n848 B.n14 585
R261 B.n796 B.n13 585
R262 B.n849 B.n13 585
R263 B.n795 B.n12 585
R264 B.n850 B.n12 585
R265 B.n794 B.n793 585
R266 B.n793 B.n792 585
R267 B.n791 B.n790 585
R268 B.n791 B.n8 585
R269 B.n789 B.n7 585
R270 B.n857 B.n7 585
R271 B.n788 B.n6 585
R272 B.n858 B.n6 585
R273 B.n787 B.n5 585
R274 B.n859 B.n5 585
R275 B.n786 B.n785 585
R276 B.n785 B.n4 585
R277 B.n784 B.n364 585
R278 B.n784 B.n783 585
R279 B.n773 B.n365 585
R280 B.n776 B.n365 585
R281 B.n775 B.n774 585
R282 B.n777 B.n775 585
R283 B.n772 B.n370 585
R284 B.n370 B.n369 585
R285 B.n771 B.n770 585
R286 B.n770 B.n769 585
R287 B.n372 B.n371 585
R288 B.n373 B.n372 585
R289 B.n762 B.n761 585
R290 B.n763 B.n762 585
R291 B.n760 B.n378 585
R292 B.n378 B.n377 585
R293 B.n759 B.n758 585
R294 B.n758 B.n757 585
R295 B.n380 B.n379 585
R296 B.n381 B.n380 585
R297 B.n750 B.n749 585
R298 B.n751 B.n750 585
R299 B.n748 B.n386 585
R300 B.n386 B.n385 585
R301 B.n747 B.n746 585
R302 B.n746 B.n745 585
R303 B.n388 B.n387 585
R304 B.n738 B.n388 585
R305 B.n737 B.n736 585
R306 B.n739 B.n737 585
R307 B.n735 B.n393 585
R308 B.n393 B.n392 585
R309 B.n734 B.n733 585
R310 B.n733 B.n732 585
R311 B.n395 B.n394 585
R312 B.n396 B.n395 585
R313 B.n728 B.n727 585
R314 B.n399 B.n398 585
R315 B.n724 B.n723 585
R316 B.n725 B.n724 585
R317 B.n722 B.n464 585
R318 B.n721 B.n720 585
R319 B.n719 B.n718 585
R320 B.n717 B.n716 585
R321 B.n715 B.n714 585
R322 B.n713 B.n712 585
R323 B.n711 B.n710 585
R324 B.n709 B.n708 585
R325 B.n707 B.n706 585
R326 B.n705 B.n704 585
R327 B.n703 B.n702 585
R328 B.n701 B.n700 585
R329 B.n699 B.n698 585
R330 B.n697 B.n696 585
R331 B.n695 B.n694 585
R332 B.n693 B.n692 585
R333 B.n691 B.n690 585
R334 B.n689 B.n688 585
R335 B.n687 B.n686 585
R336 B.n685 B.n684 585
R337 B.n683 B.n682 585
R338 B.n681 B.n680 585
R339 B.n679 B.n678 585
R340 B.n677 B.n676 585
R341 B.n675 B.n674 585
R342 B.n673 B.n672 585
R343 B.n671 B.n670 585
R344 B.n669 B.n668 585
R345 B.n667 B.n666 585
R346 B.n665 B.n664 585
R347 B.n663 B.n662 585
R348 B.n661 B.n660 585
R349 B.n659 B.n658 585
R350 B.n657 B.n656 585
R351 B.n655 B.n654 585
R352 B.n653 B.n652 585
R353 B.n651 B.n650 585
R354 B.n649 B.n648 585
R355 B.n647 B.n646 585
R356 B.n645 B.n644 585
R357 B.n643 B.n642 585
R358 B.n641 B.n640 585
R359 B.n639 B.n638 585
R360 B.n637 B.n636 585
R361 B.n635 B.n634 585
R362 B.n633 B.n632 585
R363 B.n631 B.n630 585
R364 B.n629 B.n628 585
R365 B.n627 B.n626 585
R366 B.n625 B.n624 585
R367 B.n623 B.n622 585
R368 B.n621 B.n620 585
R369 B.n619 B.n618 585
R370 B.n617 B.n616 585
R371 B.n615 B.n614 585
R372 B.n613 B.n612 585
R373 B.n611 B.n610 585
R374 B.n608 B.n607 585
R375 B.n606 B.n605 585
R376 B.n604 B.n603 585
R377 B.n602 B.n601 585
R378 B.n600 B.n599 585
R379 B.n598 B.n597 585
R380 B.n596 B.n595 585
R381 B.n594 B.n593 585
R382 B.n592 B.n591 585
R383 B.n590 B.n589 585
R384 B.n587 B.n586 585
R385 B.n585 B.n584 585
R386 B.n583 B.n582 585
R387 B.n581 B.n580 585
R388 B.n579 B.n578 585
R389 B.n577 B.n576 585
R390 B.n575 B.n574 585
R391 B.n573 B.n572 585
R392 B.n571 B.n570 585
R393 B.n569 B.n568 585
R394 B.n567 B.n566 585
R395 B.n565 B.n564 585
R396 B.n563 B.n562 585
R397 B.n561 B.n560 585
R398 B.n559 B.n558 585
R399 B.n557 B.n556 585
R400 B.n555 B.n554 585
R401 B.n553 B.n552 585
R402 B.n551 B.n550 585
R403 B.n549 B.n548 585
R404 B.n547 B.n546 585
R405 B.n545 B.n544 585
R406 B.n543 B.n542 585
R407 B.n541 B.n540 585
R408 B.n539 B.n538 585
R409 B.n537 B.n536 585
R410 B.n535 B.n534 585
R411 B.n533 B.n532 585
R412 B.n531 B.n530 585
R413 B.n529 B.n528 585
R414 B.n527 B.n526 585
R415 B.n525 B.n524 585
R416 B.n523 B.n522 585
R417 B.n521 B.n520 585
R418 B.n519 B.n518 585
R419 B.n517 B.n516 585
R420 B.n515 B.n514 585
R421 B.n513 B.n512 585
R422 B.n511 B.n510 585
R423 B.n509 B.n508 585
R424 B.n507 B.n506 585
R425 B.n505 B.n504 585
R426 B.n503 B.n502 585
R427 B.n501 B.n500 585
R428 B.n499 B.n498 585
R429 B.n497 B.n496 585
R430 B.n495 B.n494 585
R431 B.n493 B.n492 585
R432 B.n491 B.n490 585
R433 B.n489 B.n488 585
R434 B.n487 B.n486 585
R435 B.n485 B.n484 585
R436 B.n483 B.n482 585
R437 B.n481 B.n480 585
R438 B.n479 B.n478 585
R439 B.n477 B.n476 585
R440 B.n475 B.n474 585
R441 B.n473 B.n472 585
R442 B.n471 B.n470 585
R443 B.n469 B.n463 585
R444 B.n725 B.n463 585
R445 B.n729 B.n397 585
R446 B.n397 B.n396 585
R447 B.n731 B.n730 585
R448 B.n732 B.n731 585
R449 B.n391 B.n390 585
R450 B.n392 B.n391 585
R451 B.n741 B.n740 585
R452 B.n740 B.n739 585
R453 B.n742 B.n389 585
R454 B.n738 B.n389 585
R455 B.n744 B.n743 585
R456 B.n745 B.n744 585
R457 B.n384 B.n383 585
R458 B.n385 B.n384 585
R459 B.n753 B.n752 585
R460 B.n752 B.n751 585
R461 B.n754 B.n382 585
R462 B.n382 B.n381 585
R463 B.n756 B.n755 585
R464 B.n757 B.n756 585
R465 B.n376 B.n375 585
R466 B.n377 B.n376 585
R467 B.n765 B.n764 585
R468 B.n764 B.n763 585
R469 B.n766 B.n374 585
R470 B.n374 B.n373 585
R471 B.n768 B.n767 585
R472 B.n769 B.n768 585
R473 B.n368 B.n367 585
R474 B.n369 B.n368 585
R475 B.n779 B.n778 585
R476 B.n778 B.n777 585
R477 B.n780 B.n366 585
R478 B.n776 B.n366 585
R479 B.n782 B.n781 585
R480 B.n783 B.n782 585
R481 B.n3 B.n0 585
R482 B.n4 B.n3 585
R483 B.n856 B.n1 585
R484 B.n857 B.n856 585
R485 B.n855 B.n854 585
R486 B.n855 B.n8 585
R487 B.n853 B.n9 585
R488 B.n792 B.n9 585
R489 B.n852 B.n851 585
R490 B.n851 B.n850 585
R491 B.n11 B.n10 585
R492 B.n849 B.n11 585
R493 B.n847 B.n846 585
R494 B.n848 B.n847 585
R495 B.n845 B.n16 585
R496 B.n16 B.n15 585
R497 B.n844 B.n843 585
R498 B.n843 B.n842 585
R499 B.n18 B.n17 585
R500 B.n841 B.n18 585
R501 B.n839 B.n838 585
R502 B.n840 B.n839 585
R503 B.n837 B.n23 585
R504 B.n23 B.n22 585
R505 B.n836 B.n835 585
R506 B.n835 B.n834 585
R507 B.n25 B.n24 585
R508 B.n833 B.n25 585
R509 B.n831 B.n830 585
R510 B.n832 B.n831 585
R511 B.n829 B.n29 585
R512 B.n32 B.n29 585
R513 B.n828 B.n827 585
R514 B.n827 B.n826 585
R515 B.n31 B.n30 585
R516 B.n825 B.n31 585
R517 B.n823 B.n822 585
R518 B.n824 B.n823 585
R519 B.n821 B.n37 585
R520 B.n37 B.n36 585
R521 B.n860 B.n859 585
R522 B.n858 B.n2 585
R523 B.n819 B.n37 535.745
R524 B.n815 B.n104 535.745
R525 B.n463 B.n395 535.745
R526 B.n727 B.n397 535.745
R527 B.n817 B.n816 256.663
R528 B.n817 B.n102 256.663
R529 B.n817 B.n101 256.663
R530 B.n817 B.n100 256.663
R531 B.n817 B.n99 256.663
R532 B.n817 B.n98 256.663
R533 B.n817 B.n97 256.663
R534 B.n817 B.n96 256.663
R535 B.n817 B.n95 256.663
R536 B.n817 B.n94 256.663
R537 B.n817 B.n93 256.663
R538 B.n817 B.n92 256.663
R539 B.n817 B.n91 256.663
R540 B.n817 B.n90 256.663
R541 B.n817 B.n89 256.663
R542 B.n817 B.n88 256.663
R543 B.n817 B.n87 256.663
R544 B.n817 B.n86 256.663
R545 B.n817 B.n85 256.663
R546 B.n817 B.n84 256.663
R547 B.n817 B.n83 256.663
R548 B.n817 B.n82 256.663
R549 B.n817 B.n81 256.663
R550 B.n817 B.n80 256.663
R551 B.n817 B.n79 256.663
R552 B.n817 B.n78 256.663
R553 B.n817 B.n77 256.663
R554 B.n817 B.n76 256.663
R555 B.n817 B.n75 256.663
R556 B.n817 B.n74 256.663
R557 B.n817 B.n73 256.663
R558 B.n817 B.n72 256.663
R559 B.n817 B.n71 256.663
R560 B.n817 B.n70 256.663
R561 B.n817 B.n69 256.663
R562 B.n817 B.n68 256.663
R563 B.n817 B.n67 256.663
R564 B.n817 B.n66 256.663
R565 B.n817 B.n65 256.663
R566 B.n817 B.n64 256.663
R567 B.n817 B.n63 256.663
R568 B.n817 B.n62 256.663
R569 B.n817 B.n61 256.663
R570 B.n817 B.n60 256.663
R571 B.n817 B.n59 256.663
R572 B.n817 B.n58 256.663
R573 B.n817 B.n57 256.663
R574 B.n817 B.n56 256.663
R575 B.n817 B.n55 256.663
R576 B.n817 B.n54 256.663
R577 B.n817 B.n53 256.663
R578 B.n817 B.n52 256.663
R579 B.n817 B.n51 256.663
R580 B.n817 B.n50 256.663
R581 B.n817 B.n49 256.663
R582 B.n817 B.n48 256.663
R583 B.n817 B.n47 256.663
R584 B.n817 B.n46 256.663
R585 B.n817 B.n45 256.663
R586 B.n817 B.n44 256.663
R587 B.n817 B.n43 256.663
R588 B.n817 B.n42 256.663
R589 B.n817 B.n41 256.663
R590 B.n817 B.n40 256.663
R591 B.n818 B.n817 256.663
R592 B.n726 B.n725 256.663
R593 B.n725 B.n400 256.663
R594 B.n725 B.n401 256.663
R595 B.n725 B.n402 256.663
R596 B.n725 B.n403 256.663
R597 B.n725 B.n404 256.663
R598 B.n725 B.n405 256.663
R599 B.n725 B.n406 256.663
R600 B.n725 B.n407 256.663
R601 B.n725 B.n408 256.663
R602 B.n725 B.n409 256.663
R603 B.n725 B.n410 256.663
R604 B.n725 B.n411 256.663
R605 B.n725 B.n412 256.663
R606 B.n725 B.n413 256.663
R607 B.n725 B.n414 256.663
R608 B.n725 B.n415 256.663
R609 B.n725 B.n416 256.663
R610 B.n725 B.n417 256.663
R611 B.n725 B.n418 256.663
R612 B.n725 B.n419 256.663
R613 B.n725 B.n420 256.663
R614 B.n725 B.n421 256.663
R615 B.n725 B.n422 256.663
R616 B.n725 B.n423 256.663
R617 B.n725 B.n424 256.663
R618 B.n725 B.n425 256.663
R619 B.n725 B.n426 256.663
R620 B.n725 B.n427 256.663
R621 B.n725 B.n428 256.663
R622 B.n725 B.n429 256.663
R623 B.n725 B.n430 256.663
R624 B.n725 B.n431 256.663
R625 B.n725 B.n432 256.663
R626 B.n725 B.n433 256.663
R627 B.n725 B.n434 256.663
R628 B.n725 B.n435 256.663
R629 B.n725 B.n436 256.663
R630 B.n725 B.n437 256.663
R631 B.n725 B.n438 256.663
R632 B.n725 B.n439 256.663
R633 B.n725 B.n440 256.663
R634 B.n725 B.n441 256.663
R635 B.n725 B.n442 256.663
R636 B.n725 B.n443 256.663
R637 B.n725 B.n444 256.663
R638 B.n725 B.n445 256.663
R639 B.n725 B.n446 256.663
R640 B.n725 B.n447 256.663
R641 B.n725 B.n448 256.663
R642 B.n725 B.n449 256.663
R643 B.n725 B.n450 256.663
R644 B.n725 B.n451 256.663
R645 B.n725 B.n452 256.663
R646 B.n725 B.n453 256.663
R647 B.n725 B.n454 256.663
R648 B.n725 B.n455 256.663
R649 B.n725 B.n456 256.663
R650 B.n725 B.n457 256.663
R651 B.n725 B.n458 256.663
R652 B.n725 B.n459 256.663
R653 B.n725 B.n460 256.663
R654 B.n725 B.n461 256.663
R655 B.n725 B.n462 256.663
R656 B.n862 B.n861 256.663
R657 B.n111 B.n39 163.367
R658 B.n115 B.n114 163.367
R659 B.n119 B.n118 163.367
R660 B.n123 B.n122 163.367
R661 B.n127 B.n126 163.367
R662 B.n131 B.n130 163.367
R663 B.n135 B.n134 163.367
R664 B.n139 B.n138 163.367
R665 B.n143 B.n142 163.367
R666 B.n147 B.n146 163.367
R667 B.n151 B.n150 163.367
R668 B.n155 B.n154 163.367
R669 B.n159 B.n158 163.367
R670 B.n163 B.n162 163.367
R671 B.n167 B.n166 163.367
R672 B.n171 B.n170 163.367
R673 B.n175 B.n174 163.367
R674 B.n179 B.n178 163.367
R675 B.n183 B.n182 163.367
R676 B.n187 B.n186 163.367
R677 B.n191 B.n190 163.367
R678 B.n195 B.n194 163.367
R679 B.n199 B.n198 163.367
R680 B.n203 B.n202 163.367
R681 B.n207 B.n206 163.367
R682 B.n211 B.n210 163.367
R683 B.n215 B.n214 163.367
R684 B.n219 B.n218 163.367
R685 B.n223 B.n222 163.367
R686 B.n227 B.n226 163.367
R687 B.n231 B.n230 163.367
R688 B.n235 B.n234 163.367
R689 B.n239 B.n238 163.367
R690 B.n243 B.n242 163.367
R691 B.n247 B.n246 163.367
R692 B.n251 B.n250 163.367
R693 B.n255 B.n254 163.367
R694 B.n259 B.n258 163.367
R695 B.n263 B.n262 163.367
R696 B.n267 B.n266 163.367
R697 B.n271 B.n270 163.367
R698 B.n275 B.n274 163.367
R699 B.n279 B.n278 163.367
R700 B.n283 B.n282 163.367
R701 B.n287 B.n286 163.367
R702 B.n291 B.n290 163.367
R703 B.n295 B.n294 163.367
R704 B.n299 B.n298 163.367
R705 B.n303 B.n302 163.367
R706 B.n307 B.n306 163.367
R707 B.n311 B.n310 163.367
R708 B.n315 B.n314 163.367
R709 B.n319 B.n318 163.367
R710 B.n323 B.n322 163.367
R711 B.n327 B.n326 163.367
R712 B.n331 B.n330 163.367
R713 B.n335 B.n334 163.367
R714 B.n339 B.n338 163.367
R715 B.n343 B.n342 163.367
R716 B.n347 B.n346 163.367
R717 B.n351 B.n350 163.367
R718 B.n355 B.n354 163.367
R719 B.n359 B.n358 163.367
R720 B.n361 B.n103 163.367
R721 B.n733 B.n395 163.367
R722 B.n733 B.n393 163.367
R723 B.n737 B.n393 163.367
R724 B.n737 B.n388 163.367
R725 B.n746 B.n388 163.367
R726 B.n746 B.n386 163.367
R727 B.n750 B.n386 163.367
R728 B.n750 B.n380 163.367
R729 B.n758 B.n380 163.367
R730 B.n758 B.n378 163.367
R731 B.n762 B.n378 163.367
R732 B.n762 B.n372 163.367
R733 B.n770 B.n372 163.367
R734 B.n770 B.n370 163.367
R735 B.n775 B.n370 163.367
R736 B.n775 B.n365 163.367
R737 B.n784 B.n365 163.367
R738 B.n785 B.n784 163.367
R739 B.n785 B.n5 163.367
R740 B.n6 B.n5 163.367
R741 B.n7 B.n6 163.367
R742 B.n791 B.n7 163.367
R743 B.n793 B.n791 163.367
R744 B.n793 B.n12 163.367
R745 B.n13 B.n12 163.367
R746 B.n14 B.n13 163.367
R747 B.n798 B.n14 163.367
R748 B.n798 B.n19 163.367
R749 B.n20 B.n19 163.367
R750 B.n21 B.n20 163.367
R751 B.n803 B.n21 163.367
R752 B.n803 B.n26 163.367
R753 B.n27 B.n26 163.367
R754 B.n28 B.n27 163.367
R755 B.n808 B.n28 163.367
R756 B.n808 B.n33 163.367
R757 B.n34 B.n33 163.367
R758 B.n35 B.n34 163.367
R759 B.n104 B.n35 163.367
R760 B.n724 B.n399 163.367
R761 B.n724 B.n464 163.367
R762 B.n720 B.n719 163.367
R763 B.n716 B.n715 163.367
R764 B.n712 B.n711 163.367
R765 B.n708 B.n707 163.367
R766 B.n704 B.n703 163.367
R767 B.n700 B.n699 163.367
R768 B.n696 B.n695 163.367
R769 B.n692 B.n691 163.367
R770 B.n688 B.n687 163.367
R771 B.n684 B.n683 163.367
R772 B.n680 B.n679 163.367
R773 B.n676 B.n675 163.367
R774 B.n672 B.n671 163.367
R775 B.n668 B.n667 163.367
R776 B.n664 B.n663 163.367
R777 B.n660 B.n659 163.367
R778 B.n656 B.n655 163.367
R779 B.n652 B.n651 163.367
R780 B.n648 B.n647 163.367
R781 B.n644 B.n643 163.367
R782 B.n640 B.n639 163.367
R783 B.n636 B.n635 163.367
R784 B.n632 B.n631 163.367
R785 B.n628 B.n627 163.367
R786 B.n624 B.n623 163.367
R787 B.n620 B.n619 163.367
R788 B.n616 B.n615 163.367
R789 B.n612 B.n611 163.367
R790 B.n607 B.n606 163.367
R791 B.n603 B.n602 163.367
R792 B.n599 B.n598 163.367
R793 B.n595 B.n594 163.367
R794 B.n591 B.n590 163.367
R795 B.n586 B.n585 163.367
R796 B.n582 B.n581 163.367
R797 B.n578 B.n577 163.367
R798 B.n574 B.n573 163.367
R799 B.n570 B.n569 163.367
R800 B.n566 B.n565 163.367
R801 B.n562 B.n561 163.367
R802 B.n558 B.n557 163.367
R803 B.n554 B.n553 163.367
R804 B.n550 B.n549 163.367
R805 B.n546 B.n545 163.367
R806 B.n542 B.n541 163.367
R807 B.n538 B.n537 163.367
R808 B.n534 B.n533 163.367
R809 B.n530 B.n529 163.367
R810 B.n526 B.n525 163.367
R811 B.n522 B.n521 163.367
R812 B.n518 B.n517 163.367
R813 B.n514 B.n513 163.367
R814 B.n510 B.n509 163.367
R815 B.n506 B.n505 163.367
R816 B.n502 B.n501 163.367
R817 B.n498 B.n497 163.367
R818 B.n494 B.n493 163.367
R819 B.n490 B.n489 163.367
R820 B.n486 B.n485 163.367
R821 B.n482 B.n481 163.367
R822 B.n478 B.n477 163.367
R823 B.n474 B.n473 163.367
R824 B.n470 B.n463 163.367
R825 B.n731 B.n397 163.367
R826 B.n731 B.n391 163.367
R827 B.n740 B.n391 163.367
R828 B.n740 B.n389 163.367
R829 B.n744 B.n389 163.367
R830 B.n744 B.n384 163.367
R831 B.n752 B.n384 163.367
R832 B.n752 B.n382 163.367
R833 B.n756 B.n382 163.367
R834 B.n756 B.n376 163.367
R835 B.n764 B.n376 163.367
R836 B.n764 B.n374 163.367
R837 B.n768 B.n374 163.367
R838 B.n768 B.n368 163.367
R839 B.n778 B.n368 163.367
R840 B.n778 B.n366 163.367
R841 B.n782 B.n366 163.367
R842 B.n782 B.n3 163.367
R843 B.n860 B.n3 163.367
R844 B.n856 B.n2 163.367
R845 B.n856 B.n855 163.367
R846 B.n855 B.n9 163.367
R847 B.n851 B.n9 163.367
R848 B.n851 B.n11 163.367
R849 B.n847 B.n11 163.367
R850 B.n847 B.n16 163.367
R851 B.n843 B.n16 163.367
R852 B.n843 B.n18 163.367
R853 B.n839 B.n18 163.367
R854 B.n839 B.n23 163.367
R855 B.n835 B.n23 163.367
R856 B.n835 B.n25 163.367
R857 B.n831 B.n25 163.367
R858 B.n831 B.n29 163.367
R859 B.n827 B.n29 163.367
R860 B.n827 B.n31 163.367
R861 B.n823 B.n31 163.367
R862 B.n823 B.n37 163.367
R863 B.n105 B.t16 80.0272
R864 B.n467 B.t13 80.0272
R865 B.n108 B.t22 80.0025
R866 B.n465 B.t20 80.0025
R867 B.n819 B.n818 71.676
R868 B.n111 B.n40 71.676
R869 B.n115 B.n41 71.676
R870 B.n119 B.n42 71.676
R871 B.n123 B.n43 71.676
R872 B.n127 B.n44 71.676
R873 B.n131 B.n45 71.676
R874 B.n135 B.n46 71.676
R875 B.n139 B.n47 71.676
R876 B.n143 B.n48 71.676
R877 B.n147 B.n49 71.676
R878 B.n151 B.n50 71.676
R879 B.n155 B.n51 71.676
R880 B.n159 B.n52 71.676
R881 B.n163 B.n53 71.676
R882 B.n167 B.n54 71.676
R883 B.n171 B.n55 71.676
R884 B.n175 B.n56 71.676
R885 B.n179 B.n57 71.676
R886 B.n183 B.n58 71.676
R887 B.n187 B.n59 71.676
R888 B.n191 B.n60 71.676
R889 B.n195 B.n61 71.676
R890 B.n199 B.n62 71.676
R891 B.n203 B.n63 71.676
R892 B.n207 B.n64 71.676
R893 B.n211 B.n65 71.676
R894 B.n215 B.n66 71.676
R895 B.n219 B.n67 71.676
R896 B.n223 B.n68 71.676
R897 B.n227 B.n69 71.676
R898 B.n231 B.n70 71.676
R899 B.n235 B.n71 71.676
R900 B.n239 B.n72 71.676
R901 B.n243 B.n73 71.676
R902 B.n247 B.n74 71.676
R903 B.n251 B.n75 71.676
R904 B.n255 B.n76 71.676
R905 B.n259 B.n77 71.676
R906 B.n263 B.n78 71.676
R907 B.n267 B.n79 71.676
R908 B.n271 B.n80 71.676
R909 B.n275 B.n81 71.676
R910 B.n279 B.n82 71.676
R911 B.n283 B.n83 71.676
R912 B.n287 B.n84 71.676
R913 B.n291 B.n85 71.676
R914 B.n295 B.n86 71.676
R915 B.n299 B.n87 71.676
R916 B.n303 B.n88 71.676
R917 B.n307 B.n89 71.676
R918 B.n311 B.n90 71.676
R919 B.n315 B.n91 71.676
R920 B.n319 B.n92 71.676
R921 B.n323 B.n93 71.676
R922 B.n327 B.n94 71.676
R923 B.n331 B.n95 71.676
R924 B.n335 B.n96 71.676
R925 B.n339 B.n97 71.676
R926 B.n343 B.n98 71.676
R927 B.n347 B.n99 71.676
R928 B.n351 B.n100 71.676
R929 B.n355 B.n101 71.676
R930 B.n359 B.n102 71.676
R931 B.n816 B.n103 71.676
R932 B.n816 B.n815 71.676
R933 B.n361 B.n102 71.676
R934 B.n358 B.n101 71.676
R935 B.n354 B.n100 71.676
R936 B.n350 B.n99 71.676
R937 B.n346 B.n98 71.676
R938 B.n342 B.n97 71.676
R939 B.n338 B.n96 71.676
R940 B.n334 B.n95 71.676
R941 B.n330 B.n94 71.676
R942 B.n326 B.n93 71.676
R943 B.n322 B.n92 71.676
R944 B.n318 B.n91 71.676
R945 B.n314 B.n90 71.676
R946 B.n310 B.n89 71.676
R947 B.n306 B.n88 71.676
R948 B.n302 B.n87 71.676
R949 B.n298 B.n86 71.676
R950 B.n294 B.n85 71.676
R951 B.n290 B.n84 71.676
R952 B.n286 B.n83 71.676
R953 B.n282 B.n82 71.676
R954 B.n278 B.n81 71.676
R955 B.n274 B.n80 71.676
R956 B.n270 B.n79 71.676
R957 B.n266 B.n78 71.676
R958 B.n262 B.n77 71.676
R959 B.n258 B.n76 71.676
R960 B.n254 B.n75 71.676
R961 B.n250 B.n74 71.676
R962 B.n246 B.n73 71.676
R963 B.n242 B.n72 71.676
R964 B.n238 B.n71 71.676
R965 B.n234 B.n70 71.676
R966 B.n230 B.n69 71.676
R967 B.n226 B.n68 71.676
R968 B.n222 B.n67 71.676
R969 B.n218 B.n66 71.676
R970 B.n214 B.n65 71.676
R971 B.n210 B.n64 71.676
R972 B.n206 B.n63 71.676
R973 B.n202 B.n62 71.676
R974 B.n198 B.n61 71.676
R975 B.n194 B.n60 71.676
R976 B.n190 B.n59 71.676
R977 B.n186 B.n58 71.676
R978 B.n182 B.n57 71.676
R979 B.n178 B.n56 71.676
R980 B.n174 B.n55 71.676
R981 B.n170 B.n54 71.676
R982 B.n166 B.n53 71.676
R983 B.n162 B.n52 71.676
R984 B.n158 B.n51 71.676
R985 B.n154 B.n50 71.676
R986 B.n150 B.n49 71.676
R987 B.n146 B.n48 71.676
R988 B.n142 B.n47 71.676
R989 B.n138 B.n46 71.676
R990 B.n134 B.n45 71.676
R991 B.n130 B.n44 71.676
R992 B.n126 B.n43 71.676
R993 B.n122 B.n42 71.676
R994 B.n118 B.n41 71.676
R995 B.n114 B.n40 71.676
R996 B.n818 B.n39 71.676
R997 B.n727 B.n726 71.676
R998 B.n464 B.n400 71.676
R999 B.n719 B.n401 71.676
R1000 B.n715 B.n402 71.676
R1001 B.n711 B.n403 71.676
R1002 B.n707 B.n404 71.676
R1003 B.n703 B.n405 71.676
R1004 B.n699 B.n406 71.676
R1005 B.n695 B.n407 71.676
R1006 B.n691 B.n408 71.676
R1007 B.n687 B.n409 71.676
R1008 B.n683 B.n410 71.676
R1009 B.n679 B.n411 71.676
R1010 B.n675 B.n412 71.676
R1011 B.n671 B.n413 71.676
R1012 B.n667 B.n414 71.676
R1013 B.n663 B.n415 71.676
R1014 B.n659 B.n416 71.676
R1015 B.n655 B.n417 71.676
R1016 B.n651 B.n418 71.676
R1017 B.n647 B.n419 71.676
R1018 B.n643 B.n420 71.676
R1019 B.n639 B.n421 71.676
R1020 B.n635 B.n422 71.676
R1021 B.n631 B.n423 71.676
R1022 B.n627 B.n424 71.676
R1023 B.n623 B.n425 71.676
R1024 B.n619 B.n426 71.676
R1025 B.n615 B.n427 71.676
R1026 B.n611 B.n428 71.676
R1027 B.n606 B.n429 71.676
R1028 B.n602 B.n430 71.676
R1029 B.n598 B.n431 71.676
R1030 B.n594 B.n432 71.676
R1031 B.n590 B.n433 71.676
R1032 B.n585 B.n434 71.676
R1033 B.n581 B.n435 71.676
R1034 B.n577 B.n436 71.676
R1035 B.n573 B.n437 71.676
R1036 B.n569 B.n438 71.676
R1037 B.n565 B.n439 71.676
R1038 B.n561 B.n440 71.676
R1039 B.n557 B.n441 71.676
R1040 B.n553 B.n442 71.676
R1041 B.n549 B.n443 71.676
R1042 B.n545 B.n444 71.676
R1043 B.n541 B.n445 71.676
R1044 B.n537 B.n446 71.676
R1045 B.n533 B.n447 71.676
R1046 B.n529 B.n448 71.676
R1047 B.n525 B.n449 71.676
R1048 B.n521 B.n450 71.676
R1049 B.n517 B.n451 71.676
R1050 B.n513 B.n452 71.676
R1051 B.n509 B.n453 71.676
R1052 B.n505 B.n454 71.676
R1053 B.n501 B.n455 71.676
R1054 B.n497 B.n456 71.676
R1055 B.n493 B.n457 71.676
R1056 B.n489 B.n458 71.676
R1057 B.n485 B.n459 71.676
R1058 B.n481 B.n460 71.676
R1059 B.n477 B.n461 71.676
R1060 B.n473 B.n462 71.676
R1061 B.n726 B.n399 71.676
R1062 B.n720 B.n400 71.676
R1063 B.n716 B.n401 71.676
R1064 B.n712 B.n402 71.676
R1065 B.n708 B.n403 71.676
R1066 B.n704 B.n404 71.676
R1067 B.n700 B.n405 71.676
R1068 B.n696 B.n406 71.676
R1069 B.n692 B.n407 71.676
R1070 B.n688 B.n408 71.676
R1071 B.n684 B.n409 71.676
R1072 B.n680 B.n410 71.676
R1073 B.n676 B.n411 71.676
R1074 B.n672 B.n412 71.676
R1075 B.n668 B.n413 71.676
R1076 B.n664 B.n414 71.676
R1077 B.n660 B.n415 71.676
R1078 B.n656 B.n416 71.676
R1079 B.n652 B.n417 71.676
R1080 B.n648 B.n418 71.676
R1081 B.n644 B.n419 71.676
R1082 B.n640 B.n420 71.676
R1083 B.n636 B.n421 71.676
R1084 B.n632 B.n422 71.676
R1085 B.n628 B.n423 71.676
R1086 B.n624 B.n424 71.676
R1087 B.n620 B.n425 71.676
R1088 B.n616 B.n426 71.676
R1089 B.n612 B.n427 71.676
R1090 B.n607 B.n428 71.676
R1091 B.n603 B.n429 71.676
R1092 B.n599 B.n430 71.676
R1093 B.n595 B.n431 71.676
R1094 B.n591 B.n432 71.676
R1095 B.n586 B.n433 71.676
R1096 B.n582 B.n434 71.676
R1097 B.n578 B.n435 71.676
R1098 B.n574 B.n436 71.676
R1099 B.n570 B.n437 71.676
R1100 B.n566 B.n438 71.676
R1101 B.n562 B.n439 71.676
R1102 B.n558 B.n440 71.676
R1103 B.n554 B.n441 71.676
R1104 B.n550 B.n442 71.676
R1105 B.n546 B.n443 71.676
R1106 B.n542 B.n444 71.676
R1107 B.n538 B.n445 71.676
R1108 B.n534 B.n446 71.676
R1109 B.n530 B.n447 71.676
R1110 B.n526 B.n448 71.676
R1111 B.n522 B.n449 71.676
R1112 B.n518 B.n450 71.676
R1113 B.n514 B.n451 71.676
R1114 B.n510 B.n452 71.676
R1115 B.n506 B.n453 71.676
R1116 B.n502 B.n454 71.676
R1117 B.n498 B.n455 71.676
R1118 B.n494 B.n456 71.676
R1119 B.n490 B.n457 71.676
R1120 B.n486 B.n458 71.676
R1121 B.n482 B.n459 71.676
R1122 B.n478 B.n460 71.676
R1123 B.n474 B.n461 71.676
R1124 B.n470 B.n462 71.676
R1125 B.n861 B.n860 71.676
R1126 B.n861 B.n2 71.676
R1127 B.n106 B.t17 67.4212
R1128 B.n468 B.t12 67.4212
R1129 B.n109 B.t23 67.3964
R1130 B.n466 B.t19 67.3964
R1131 B.n725 B.n396 60.0132
R1132 B.n817 B.n36 60.0132
R1133 B.n110 B.n109 59.5399
R1134 B.n107 B.n106 59.5399
R1135 B.n588 B.n468 59.5399
R1136 B.n609 B.n466 59.5399
R1137 B.n729 B.n728 34.8103
R1138 B.n469 B.n394 34.8103
R1139 B.n821 B.n820 34.8103
R1140 B.n814 B.n813 34.8103
R1141 B.n732 B.n396 31.6351
R1142 B.n732 B.n392 31.6351
R1143 B.n739 B.n392 31.6351
R1144 B.n739 B.n738 31.6351
R1145 B.n745 B.n385 31.6351
R1146 B.n751 B.n385 31.6351
R1147 B.n751 B.n381 31.6351
R1148 B.n757 B.n381 31.6351
R1149 B.n763 B.n377 31.6351
R1150 B.n769 B.n373 31.6351
R1151 B.n777 B.n369 31.6351
R1152 B.n783 B.n4 31.6351
R1153 B.n859 B.n4 31.6351
R1154 B.n859 B.n858 31.6351
R1155 B.n858 B.n857 31.6351
R1156 B.n857 B.n8 31.6351
R1157 B.n850 B.n849 31.6351
R1158 B.n848 B.n15 31.6351
R1159 B.n842 B.n841 31.6351
R1160 B.n840 B.n22 31.6351
R1161 B.n834 B.n22 31.6351
R1162 B.n834 B.n833 31.6351
R1163 B.n833 B.n832 31.6351
R1164 B.n826 B.n32 31.6351
R1165 B.n826 B.n825 31.6351
R1166 B.n825 B.n824 31.6351
R1167 B.n824 B.n36 31.6351
R1168 B.t4 B.n776 30.7047
R1169 B.n792 B.t7 30.7047
R1170 B.n776 B.t1 29.7742
R1171 B.n792 B.t9 29.7742
R1172 B.t6 B.n369 27.9134
R1173 B.n849 B.t2 27.9134
R1174 B.n745 B.t11 26.0525
R1175 B.n832 B.t15 26.0525
R1176 B.t5 B.n373 25.1221
R1177 B.t0 B.n15 25.1221
R1178 B.t3 B.n377 22.3308
R1179 B.n841 B.t8 22.3308
R1180 B B.n862 18.0485
R1181 B.n109 B.n108 12.6066
R1182 B.n106 B.n105 12.6066
R1183 B.n468 B.n467 12.6066
R1184 B.n466 B.n465 12.6066
R1185 B.n730 B.n729 10.6151
R1186 B.n730 B.n390 10.6151
R1187 B.n741 B.n390 10.6151
R1188 B.n742 B.n741 10.6151
R1189 B.n743 B.n742 10.6151
R1190 B.n743 B.n383 10.6151
R1191 B.n753 B.n383 10.6151
R1192 B.n754 B.n753 10.6151
R1193 B.n755 B.n754 10.6151
R1194 B.n755 B.n375 10.6151
R1195 B.n765 B.n375 10.6151
R1196 B.n766 B.n765 10.6151
R1197 B.n767 B.n766 10.6151
R1198 B.n767 B.n367 10.6151
R1199 B.n779 B.n367 10.6151
R1200 B.n780 B.n779 10.6151
R1201 B.n781 B.n780 10.6151
R1202 B.n781 B.n0 10.6151
R1203 B.n728 B.n398 10.6151
R1204 B.n723 B.n398 10.6151
R1205 B.n723 B.n722 10.6151
R1206 B.n722 B.n721 10.6151
R1207 B.n721 B.n718 10.6151
R1208 B.n718 B.n717 10.6151
R1209 B.n717 B.n714 10.6151
R1210 B.n714 B.n713 10.6151
R1211 B.n713 B.n710 10.6151
R1212 B.n710 B.n709 10.6151
R1213 B.n709 B.n706 10.6151
R1214 B.n706 B.n705 10.6151
R1215 B.n705 B.n702 10.6151
R1216 B.n702 B.n701 10.6151
R1217 B.n701 B.n698 10.6151
R1218 B.n698 B.n697 10.6151
R1219 B.n697 B.n694 10.6151
R1220 B.n694 B.n693 10.6151
R1221 B.n693 B.n690 10.6151
R1222 B.n690 B.n689 10.6151
R1223 B.n689 B.n686 10.6151
R1224 B.n686 B.n685 10.6151
R1225 B.n685 B.n682 10.6151
R1226 B.n682 B.n681 10.6151
R1227 B.n681 B.n678 10.6151
R1228 B.n678 B.n677 10.6151
R1229 B.n677 B.n674 10.6151
R1230 B.n674 B.n673 10.6151
R1231 B.n673 B.n670 10.6151
R1232 B.n670 B.n669 10.6151
R1233 B.n669 B.n666 10.6151
R1234 B.n666 B.n665 10.6151
R1235 B.n665 B.n662 10.6151
R1236 B.n662 B.n661 10.6151
R1237 B.n661 B.n658 10.6151
R1238 B.n658 B.n657 10.6151
R1239 B.n657 B.n654 10.6151
R1240 B.n654 B.n653 10.6151
R1241 B.n653 B.n650 10.6151
R1242 B.n650 B.n649 10.6151
R1243 B.n649 B.n646 10.6151
R1244 B.n646 B.n645 10.6151
R1245 B.n645 B.n642 10.6151
R1246 B.n642 B.n641 10.6151
R1247 B.n641 B.n638 10.6151
R1248 B.n638 B.n637 10.6151
R1249 B.n637 B.n634 10.6151
R1250 B.n634 B.n633 10.6151
R1251 B.n633 B.n630 10.6151
R1252 B.n630 B.n629 10.6151
R1253 B.n629 B.n626 10.6151
R1254 B.n626 B.n625 10.6151
R1255 B.n625 B.n622 10.6151
R1256 B.n622 B.n621 10.6151
R1257 B.n621 B.n618 10.6151
R1258 B.n618 B.n617 10.6151
R1259 B.n617 B.n614 10.6151
R1260 B.n614 B.n613 10.6151
R1261 B.n613 B.n610 10.6151
R1262 B.n608 B.n605 10.6151
R1263 B.n605 B.n604 10.6151
R1264 B.n604 B.n601 10.6151
R1265 B.n601 B.n600 10.6151
R1266 B.n600 B.n597 10.6151
R1267 B.n597 B.n596 10.6151
R1268 B.n596 B.n593 10.6151
R1269 B.n593 B.n592 10.6151
R1270 B.n592 B.n589 10.6151
R1271 B.n587 B.n584 10.6151
R1272 B.n584 B.n583 10.6151
R1273 B.n583 B.n580 10.6151
R1274 B.n580 B.n579 10.6151
R1275 B.n579 B.n576 10.6151
R1276 B.n576 B.n575 10.6151
R1277 B.n575 B.n572 10.6151
R1278 B.n572 B.n571 10.6151
R1279 B.n571 B.n568 10.6151
R1280 B.n568 B.n567 10.6151
R1281 B.n567 B.n564 10.6151
R1282 B.n564 B.n563 10.6151
R1283 B.n563 B.n560 10.6151
R1284 B.n560 B.n559 10.6151
R1285 B.n559 B.n556 10.6151
R1286 B.n556 B.n555 10.6151
R1287 B.n555 B.n552 10.6151
R1288 B.n552 B.n551 10.6151
R1289 B.n551 B.n548 10.6151
R1290 B.n548 B.n547 10.6151
R1291 B.n547 B.n544 10.6151
R1292 B.n544 B.n543 10.6151
R1293 B.n543 B.n540 10.6151
R1294 B.n540 B.n539 10.6151
R1295 B.n539 B.n536 10.6151
R1296 B.n536 B.n535 10.6151
R1297 B.n535 B.n532 10.6151
R1298 B.n532 B.n531 10.6151
R1299 B.n531 B.n528 10.6151
R1300 B.n528 B.n527 10.6151
R1301 B.n527 B.n524 10.6151
R1302 B.n524 B.n523 10.6151
R1303 B.n523 B.n520 10.6151
R1304 B.n520 B.n519 10.6151
R1305 B.n519 B.n516 10.6151
R1306 B.n516 B.n515 10.6151
R1307 B.n515 B.n512 10.6151
R1308 B.n512 B.n511 10.6151
R1309 B.n511 B.n508 10.6151
R1310 B.n508 B.n507 10.6151
R1311 B.n507 B.n504 10.6151
R1312 B.n504 B.n503 10.6151
R1313 B.n503 B.n500 10.6151
R1314 B.n500 B.n499 10.6151
R1315 B.n499 B.n496 10.6151
R1316 B.n496 B.n495 10.6151
R1317 B.n495 B.n492 10.6151
R1318 B.n492 B.n491 10.6151
R1319 B.n491 B.n488 10.6151
R1320 B.n488 B.n487 10.6151
R1321 B.n487 B.n484 10.6151
R1322 B.n484 B.n483 10.6151
R1323 B.n483 B.n480 10.6151
R1324 B.n480 B.n479 10.6151
R1325 B.n479 B.n476 10.6151
R1326 B.n476 B.n475 10.6151
R1327 B.n475 B.n472 10.6151
R1328 B.n472 B.n471 10.6151
R1329 B.n471 B.n469 10.6151
R1330 B.n734 B.n394 10.6151
R1331 B.n735 B.n734 10.6151
R1332 B.n736 B.n735 10.6151
R1333 B.n736 B.n387 10.6151
R1334 B.n747 B.n387 10.6151
R1335 B.n748 B.n747 10.6151
R1336 B.n749 B.n748 10.6151
R1337 B.n749 B.n379 10.6151
R1338 B.n759 B.n379 10.6151
R1339 B.n760 B.n759 10.6151
R1340 B.n761 B.n760 10.6151
R1341 B.n761 B.n371 10.6151
R1342 B.n771 B.n371 10.6151
R1343 B.n772 B.n771 10.6151
R1344 B.n774 B.n772 10.6151
R1345 B.n774 B.n773 10.6151
R1346 B.n773 B.n364 10.6151
R1347 B.n786 B.n364 10.6151
R1348 B.n787 B.n786 10.6151
R1349 B.n788 B.n787 10.6151
R1350 B.n789 B.n788 10.6151
R1351 B.n790 B.n789 10.6151
R1352 B.n794 B.n790 10.6151
R1353 B.n795 B.n794 10.6151
R1354 B.n796 B.n795 10.6151
R1355 B.n797 B.n796 10.6151
R1356 B.n799 B.n797 10.6151
R1357 B.n800 B.n799 10.6151
R1358 B.n801 B.n800 10.6151
R1359 B.n802 B.n801 10.6151
R1360 B.n804 B.n802 10.6151
R1361 B.n805 B.n804 10.6151
R1362 B.n806 B.n805 10.6151
R1363 B.n807 B.n806 10.6151
R1364 B.n809 B.n807 10.6151
R1365 B.n810 B.n809 10.6151
R1366 B.n811 B.n810 10.6151
R1367 B.n812 B.n811 10.6151
R1368 B.n813 B.n812 10.6151
R1369 B.n854 B.n1 10.6151
R1370 B.n854 B.n853 10.6151
R1371 B.n853 B.n852 10.6151
R1372 B.n852 B.n10 10.6151
R1373 B.n846 B.n10 10.6151
R1374 B.n846 B.n845 10.6151
R1375 B.n845 B.n844 10.6151
R1376 B.n844 B.n17 10.6151
R1377 B.n838 B.n17 10.6151
R1378 B.n838 B.n837 10.6151
R1379 B.n837 B.n836 10.6151
R1380 B.n836 B.n24 10.6151
R1381 B.n830 B.n24 10.6151
R1382 B.n830 B.n829 10.6151
R1383 B.n829 B.n828 10.6151
R1384 B.n828 B.n30 10.6151
R1385 B.n822 B.n30 10.6151
R1386 B.n822 B.n821 10.6151
R1387 B.n820 B.n38 10.6151
R1388 B.n112 B.n38 10.6151
R1389 B.n113 B.n112 10.6151
R1390 B.n116 B.n113 10.6151
R1391 B.n117 B.n116 10.6151
R1392 B.n120 B.n117 10.6151
R1393 B.n121 B.n120 10.6151
R1394 B.n124 B.n121 10.6151
R1395 B.n125 B.n124 10.6151
R1396 B.n128 B.n125 10.6151
R1397 B.n129 B.n128 10.6151
R1398 B.n132 B.n129 10.6151
R1399 B.n133 B.n132 10.6151
R1400 B.n136 B.n133 10.6151
R1401 B.n137 B.n136 10.6151
R1402 B.n140 B.n137 10.6151
R1403 B.n141 B.n140 10.6151
R1404 B.n144 B.n141 10.6151
R1405 B.n145 B.n144 10.6151
R1406 B.n148 B.n145 10.6151
R1407 B.n149 B.n148 10.6151
R1408 B.n152 B.n149 10.6151
R1409 B.n153 B.n152 10.6151
R1410 B.n156 B.n153 10.6151
R1411 B.n157 B.n156 10.6151
R1412 B.n160 B.n157 10.6151
R1413 B.n161 B.n160 10.6151
R1414 B.n164 B.n161 10.6151
R1415 B.n165 B.n164 10.6151
R1416 B.n168 B.n165 10.6151
R1417 B.n169 B.n168 10.6151
R1418 B.n172 B.n169 10.6151
R1419 B.n173 B.n172 10.6151
R1420 B.n176 B.n173 10.6151
R1421 B.n177 B.n176 10.6151
R1422 B.n180 B.n177 10.6151
R1423 B.n181 B.n180 10.6151
R1424 B.n184 B.n181 10.6151
R1425 B.n185 B.n184 10.6151
R1426 B.n188 B.n185 10.6151
R1427 B.n189 B.n188 10.6151
R1428 B.n192 B.n189 10.6151
R1429 B.n193 B.n192 10.6151
R1430 B.n196 B.n193 10.6151
R1431 B.n197 B.n196 10.6151
R1432 B.n200 B.n197 10.6151
R1433 B.n201 B.n200 10.6151
R1434 B.n204 B.n201 10.6151
R1435 B.n205 B.n204 10.6151
R1436 B.n208 B.n205 10.6151
R1437 B.n209 B.n208 10.6151
R1438 B.n212 B.n209 10.6151
R1439 B.n213 B.n212 10.6151
R1440 B.n216 B.n213 10.6151
R1441 B.n217 B.n216 10.6151
R1442 B.n220 B.n217 10.6151
R1443 B.n221 B.n220 10.6151
R1444 B.n224 B.n221 10.6151
R1445 B.n225 B.n224 10.6151
R1446 B.n229 B.n228 10.6151
R1447 B.n232 B.n229 10.6151
R1448 B.n233 B.n232 10.6151
R1449 B.n236 B.n233 10.6151
R1450 B.n237 B.n236 10.6151
R1451 B.n240 B.n237 10.6151
R1452 B.n241 B.n240 10.6151
R1453 B.n244 B.n241 10.6151
R1454 B.n245 B.n244 10.6151
R1455 B.n249 B.n248 10.6151
R1456 B.n252 B.n249 10.6151
R1457 B.n253 B.n252 10.6151
R1458 B.n256 B.n253 10.6151
R1459 B.n257 B.n256 10.6151
R1460 B.n260 B.n257 10.6151
R1461 B.n261 B.n260 10.6151
R1462 B.n264 B.n261 10.6151
R1463 B.n265 B.n264 10.6151
R1464 B.n268 B.n265 10.6151
R1465 B.n269 B.n268 10.6151
R1466 B.n272 B.n269 10.6151
R1467 B.n273 B.n272 10.6151
R1468 B.n276 B.n273 10.6151
R1469 B.n277 B.n276 10.6151
R1470 B.n280 B.n277 10.6151
R1471 B.n281 B.n280 10.6151
R1472 B.n284 B.n281 10.6151
R1473 B.n285 B.n284 10.6151
R1474 B.n288 B.n285 10.6151
R1475 B.n289 B.n288 10.6151
R1476 B.n292 B.n289 10.6151
R1477 B.n293 B.n292 10.6151
R1478 B.n296 B.n293 10.6151
R1479 B.n297 B.n296 10.6151
R1480 B.n300 B.n297 10.6151
R1481 B.n301 B.n300 10.6151
R1482 B.n304 B.n301 10.6151
R1483 B.n305 B.n304 10.6151
R1484 B.n308 B.n305 10.6151
R1485 B.n309 B.n308 10.6151
R1486 B.n312 B.n309 10.6151
R1487 B.n313 B.n312 10.6151
R1488 B.n316 B.n313 10.6151
R1489 B.n317 B.n316 10.6151
R1490 B.n320 B.n317 10.6151
R1491 B.n321 B.n320 10.6151
R1492 B.n324 B.n321 10.6151
R1493 B.n325 B.n324 10.6151
R1494 B.n328 B.n325 10.6151
R1495 B.n329 B.n328 10.6151
R1496 B.n332 B.n329 10.6151
R1497 B.n333 B.n332 10.6151
R1498 B.n336 B.n333 10.6151
R1499 B.n337 B.n336 10.6151
R1500 B.n340 B.n337 10.6151
R1501 B.n341 B.n340 10.6151
R1502 B.n344 B.n341 10.6151
R1503 B.n345 B.n344 10.6151
R1504 B.n348 B.n345 10.6151
R1505 B.n349 B.n348 10.6151
R1506 B.n352 B.n349 10.6151
R1507 B.n353 B.n352 10.6151
R1508 B.n356 B.n353 10.6151
R1509 B.n357 B.n356 10.6151
R1510 B.n360 B.n357 10.6151
R1511 B.n362 B.n360 10.6151
R1512 B.n363 B.n362 10.6151
R1513 B.n814 B.n363 10.6151
R1514 B.n610 B.n609 9.36635
R1515 B.n588 B.n587 9.36635
R1516 B.n225 B.n110 9.36635
R1517 B.n248 B.n107 9.36635
R1518 B.n757 B.t3 9.30479
R1519 B.t8 B.n840 9.30479
R1520 B.n862 B.n0 8.11757
R1521 B.n862 B.n1 8.11757
R1522 B.n763 B.t5 6.5135
R1523 B.n842 B.t0 6.5135
R1524 B.n738 B.t11 5.58308
R1525 B.n32 B.t15 5.58308
R1526 B.n769 B.t6 3.72222
R1527 B.t2 B.n848 3.72222
R1528 B.n783 B.t1 1.86136
R1529 B.t9 B.n8 1.86136
R1530 B.n609 B.n608 1.24928
R1531 B.n589 B.n588 1.24928
R1532 B.n228 B.n110 1.24928
R1533 B.n245 B.n107 1.24928
R1534 B.n777 B.t4 0.930929
R1535 B.n850 B.t7 0.930929
R1536 VP.n21 VP.t2 1525.97
R1537 VP.n14 VP.t3 1525.97
R1538 VP.n5 VP.t9 1525.97
R1539 VP.n11 VP.t8 1525.97
R1540 VP.n18 VP.t0 1482.15
R1541 VP.n20 VP.t4 1482.15
R1542 VP.n13 VP.t1 1482.15
R1543 VP.n8 VP.t6 1482.15
R1544 VP.n4 VP.t7 1482.15
R1545 VP.n10 VP.t5 1482.15
R1546 VP.n6 VP.n5 161.489
R1547 VP.n22 VP.n21 161.3
R1548 VP.n6 VP.n3 161.3
R1549 VP.n8 VP.n7 161.3
R1550 VP.n9 VP.n2 161.3
R1551 VP.n12 VP.n11 161.3
R1552 VP.n19 VP.n0 161.3
R1553 VP.n18 VP.n17 161.3
R1554 VP.n16 VP.n1 161.3
R1555 VP.n15 VP.n14 161.3
R1556 VP.n18 VP.n1 73.0308
R1557 VP.n19 VP.n18 73.0308
R1558 VP.n8 VP.n3 73.0308
R1559 VP.n9 VP.n8 73.0308
R1560 VP.n14 VP.n13 51.1217
R1561 VP.n21 VP.n20 51.1217
R1562 VP.n5 VP.n4 51.1217
R1563 VP.n11 VP.n10 51.1217
R1564 VP.n15 VP.n12 45.6331
R1565 VP.n13 VP.n1 21.9096
R1566 VP.n20 VP.n19 21.9096
R1567 VP.n4 VP.n3 21.9096
R1568 VP.n10 VP.n9 21.9096
R1569 VP.n7 VP.n6 0.189894
R1570 VP.n7 VP.n2 0.189894
R1571 VP.n12 VP.n2 0.189894
R1572 VP.n16 VP.n15 0.189894
R1573 VP.n17 VP.n16 0.189894
R1574 VP.n17 VP.n0 0.189894
R1575 VP.n22 VP.n0 0.189894
R1576 VP VP.n22 0.0516364
R1577 VDD1.n1 VDD1.t0 64.2972
R1578 VDD1.n3 VDD1.t6 64.2962
R1579 VDD1.n5 VDD1.n4 63.0237
R1580 VDD1.n1 VDD1.n0 62.659
R1581 VDD1.n3 VDD1.n2 62.6588
R1582 VDD1.n7 VDD1.n6 62.658
R1583 VDD1.n7 VDD1.n5 43.0763
R1584 VDD1.n6 VDD1.t4 1.07834
R1585 VDD1.n6 VDD1.t1 1.07834
R1586 VDD1.n0 VDD1.t2 1.07834
R1587 VDD1.n0 VDD1.t3 1.07834
R1588 VDD1.n4 VDD1.t5 1.07834
R1589 VDD1.n4 VDD1.t7 1.07834
R1590 VDD1.n2 VDD1.t8 1.07834
R1591 VDD1.n2 VDD1.t9 1.07834
R1592 VDD1 VDD1.n7 0.362569
R1593 VDD1 VDD1.n1 0.198776
R1594 VDD1.n5 VDD1.n3 0.0852402
C0 VTAIL VN 5.51168f
C1 VDD1 VDD2 0.739534f
C2 VP VDD2 0.294318f
C3 VTAIL VDD1 29.960701f
C4 VP VTAIL 5.52678f
C5 VDD1 VN 0.148015f
C6 VP VN 6.21558f
C7 VP VDD1 6.29476f
C8 VTAIL VDD2 29.9862f
C9 VN VDD2 6.15622f
C10 VDD2 B 5.687092f
C11 VDD1 B 5.555562f
C12 VTAIL B 8.284466f
C13 VN B 8.73159f
C14 VP B 6.100422f
C15 VDD1.t0 B 5.01219f
C16 VDD1.t2 B 0.428701f
C17 VDD1.t3 B 0.428701f
C18 VDD1.n0 B 3.91848f
C19 VDD1.n1 B 0.684518f
C20 VDD1.t6 B 5.0122f
C21 VDD1.t8 B 0.428701f
C22 VDD1.t9 B 0.428701f
C23 VDD1.n2 B 3.91848f
C24 VDD1.n3 B 0.681784f
C25 VDD1.t5 B 0.428701f
C26 VDD1.t7 B 0.428701f
C27 VDD1.n4 B 3.92043f
C28 VDD1.n5 B 2.54478f
C29 VDD1.t4 B 0.428701f
C30 VDD1.t1 B 0.428701f
C31 VDD1.n6 B 3.91848f
C32 VDD1.n7 B 3.20574f
C33 VP.n0 B 0.053621f
C34 VP.t4 B 0.88833f
C35 VP.t0 B 0.88833f
C36 VP.n1 B 0.022747f
C37 VP.n2 B 0.053621f
C38 VP.t5 B 0.88833f
C39 VP.t6 B 0.88833f
C40 VP.n3 B 0.022747f
C41 VP.t9 B 0.897977f
C42 VP.t7 B 0.88833f
C43 VP.n4 B 0.331982f
C44 VP.n5 B 0.349128f
C45 VP.n6 B 0.121049f
C46 VP.n7 B 0.053621f
C47 VP.n8 B 0.34977f
C48 VP.n9 B 0.022747f
C49 VP.n10 B 0.331982f
C50 VP.t8 B 0.897977f
C51 VP.n11 B 0.349049f
C52 VP.n12 B 2.53224f
C53 VP.t3 B 0.897977f
C54 VP.t1 B 0.88833f
C55 VP.n13 B 0.331982f
C56 VP.n14 B 0.349049f
C57 VP.n15 B 2.57448f
C58 VP.n16 B 0.053621f
C59 VP.n17 B 0.053621f
C60 VP.n18 B 0.34977f
C61 VP.n19 B 0.022747f
C62 VP.n20 B 0.331982f
C63 VP.t2 B 0.897977f
C64 VP.n21 B 0.349049f
C65 VP.n22 B 0.041554f
C66 VTAIL.t15 B 0.434845f
C67 VTAIL.t10 B 0.434845f
C68 VTAIL.n0 B 3.88994f
C69 VTAIL.n1 B 0.401756f
C70 VTAIL.t1 B 4.96959f
C71 VTAIL.n2 B 0.515946f
C72 VTAIL.t6 B 0.434845f
C73 VTAIL.t4 B 0.434845f
C74 VTAIL.n3 B 3.88994f
C75 VTAIL.n4 B 0.391355f
C76 VTAIL.t3 B 0.434845f
C77 VTAIL.t5 B 0.434845f
C78 VTAIL.n5 B 3.88994f
C79 VTAIL.n6 B 2.38089f
C80 VTAIL.t12 B 0.434845f
C81 VTAIL.t9 B 0.434845f
C82 VTAIL.n7 B 3.88994f
C83 VTAIL.n8 B 2.38089f
C84 VTAIL.t8 B 0.434845f
C85 VTAIL.t14 B 0.434845f
C86 VTAIL.n9 B 3.88994f
C87 VTAIL.n10 B 0.391352f
C88 VTAIL.t11 B 4.96958f
C89 VTAIL.n11 B 0.51596f
C90 VTAIL.t19 B 0.434845f
C91 VTAIL.t17 B 0.434845f
C92 VTAIL.n12 B 3.88994f
C93 VTAIL.n13 B 0.409658f
C94 VTAIL.t2 B 0.434845f
C95 VTAIL.t0 B 0.434845f
C96 VTAIL.n14 B 3.88994f
C97 VTAIL.n15 B 0.391352f
C98 VTAIL.t18 B 4.96958f
C99 VTAIL.n16 B 2.43311f
C100 VTAIL.t13 B 4.96959f
C101 VTAIL.n17 B 2.43309f
C102 VTAIL.t7 B 0.434845f
C103 VTAIL.t16 B 0.434845f
C104 VTAIL.n18 B 3.88994f
C105 VTAIL.n19 B 0.345174f
C106 VDD2.t7 B 5.01345f
C107 VDD2.t3 B 0.428808f
C108 VDD2.t5 B 0.428808f
C109 VDD2.n0 B 3.91946f
C110 VDD2.n1 B 0.681955f
C111 VDD2.t0 B 0.428808f
C112 VDD2.t2 B 0.428808f
C113 VDD2.n2 B 3.92142f
C114 VDD2.n3 B 2.46364f
C115 VDD2.t1 B 5.01013f
C116 VDD2.n4 B 3.22356f
C117 VDD2.t9 B 0.428808f
C118 VDD2.t8 B 0.428808f
C119 VDD2.n5 B 3.91946f
C120 VDD2.n6 B 0.308084f
C121 VDD2.t6 B 0.428808f
C122 VDD2.t4 B 0.428808f
C123 VDD2.n7 B 3.92139f
C124 VN.n0 B 0.053101f
C125 VN.t0 B 0.879711f
C126 VN.t9 B 0.879711f
C127 VN.n1 B 0.022526f
C128 VN.t1 B 0.889264f
C129 VN.t6 B 0.879711f
C130 VN.n2 B 0.328761f
C131 VN.n3 B 0.345741f
C132 VN.n4 B 0.119874f
C133 VN.n5 B 0.053101f
C134 VN.n6 B 0.346376f
C135 VN.n7 B 0.022526f
C136 VN.n8 B 0.328761f
C137 VN.t3 B 0.889264f
C138 VN.n9 B 0.345662f
C139 VN.n10 B 0.041151f
C140 VN.n11 B 0.053101f
C141 VN.t4 B 0.889264f
C142 VN.t7 B 0.879711f
C143 VN.t8 B 0.879711f
C144 VN.n12 B 0.022526f
C145 VN.t2 B 0.879711f
C146 VN.n13 B 0.328761f
C147 VN.t5 B 0.889264f
C148 VN.n14 B 0.345741f
C149 VN.n15 B 0.119874f
C150 VN.n16 B 0.053101f
C151 VN.n17 B 0.346376f
C152 VN.n18 B 0.022526f
C153 VN.n19 B 0.328761f
C154 VN.n20 B 0.345662f
C155 VN.n21 B 2.54236f
.ends

