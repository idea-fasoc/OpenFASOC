* NGSPICE file created from diff_pair_sample_1002.ext - technology: sky130A

.subckt diff_pair_sample_1002 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t2 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=1.37115 ps=8.64 w=8.31 l=3.21
X1 VDD2.t5 VN.t0 VTAIL.t4 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=1.37115 ps=8.64 w=8.31 l=3.21
X2 VDD1.t3 VP.t1 VTAIL.t10 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=3.2409 ps=17.4 w=8.31 l=3.21
X3 VDD1.t5 VP.t2 VTAIL.t9 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=1.37115 ps=8.64 w=8.31 l=3.21
X4 B.t11 B.t9 B.t10 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=0 ps=0 w=8.31 l=3.21
X5 VDD2.t4 VN.t1 VTAIL.t0 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=3.2409 ps=17.4 w=8.31 l=3.21
X6 VDD2.t3 VN.t2 VTAIL.t5 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=3.2409 ps=17.4 w=8.31 l=3.21
X7 VTAIL.t8 VP.t3 VDD1.t0 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=1.37115 ps=8.64 w=8.31 l=3.21
X8 VTAIL.t1 VN.t3 VDD2.t2 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=1.37115 ps=8.64 w=8.31 l=3.21
X9 VTAIL.t2 VN.t4 VDD2.t1 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=1.37115 ps=8.64 w=8.31 l=3.21
X10 B.t8 B.t6 B.t7 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=0 ps=0 w=8.31 l=3.21
X11 VDD1.t4 VP.t4 VTAIL.t7 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=1.37115 pd=8.64 as=3.2409 ps=17.4 w=8.31 l=3.21
X12 B.t5 B.t3 B.t4 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=0 ps=0 w=8.31 l=3.21
X13 VDD1.t1 VP.t5 VTAIL.t6 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=1.37115 ps=8.64 w=8.31 l=3.21
X14 VDD2.t0 VN.t5 VTAIL.t3 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=1.37115 ps=8.64 w=8.31 l=3.21
X15 B.t2 B.t0 B.t1 w_n3802_n2630# sky130_fd_pr__pfet_01v8 ad=3.2409 pd=17.4 as=0 ps=0 w=8.31 l=3.21
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t5 95.2861
R22 VP.n27 VP.n8 75.8765
R23 VP.n50 VP.n0 75.8765
R24 VP.n26 VP.n9 75.8765
R25 VP.n8 VP.t2 62.3902
R26 VP.n4 VP.t3 62.3902
R27 VP.n0 VP.t4 62.3902
R28 VP.n9 VP.t1 62.3902
R29 VP.n13 VP.t0 62.3902
R30 VP.n14 VP.n13 62.0429
R31 VP.n27 VP.n26 48.3554
R32 VP.n31 VP.n6 42.4359
R33 VP.n46 VP.n2 42.4359
R34 VP.n22 VP.n11 42.4359
R35 VP.n35 VP.n6 38.5509
R36 VP.n42 VP.n2 38.5509
R37 VP.n18 VP.n11 38.5509
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 14.1914
R51 VP.n48 VP.n0 14.1914
R52 VP.n24 VP.n9 14.1914
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 4.18228
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1 VDD1.t1 90.4524
R81 VDD1.n1 VDD1.t5 90.3388
R82 VDD1.n1 VDD1.n0 84.9013
R83 VDD1.n3 VDD1.n2 84.1938
R84 VDD1.n3 VDD1.n1 42.9061
R85 VDD1.n2 VDD1.t2 3.91205
R86 VDD1.n2 VDD1.t3 3.91205
R87 VDD1.n0 VDD1.t0 3.91205
R88 VDD1.n0 VDD1.t4 3.91205
R89 VDD1 VDD1.n3 0.705241
R90 VTAIL.n7 VTAIL.t0 71.4266
R91 VTAIL.n11 VTAIL.t5 71.4265
R92 VTAIL.n2 VTAIL.t7 71.4265
R93 VTAIL.n10 VTAIL.t10 71.4265
R94 VTAIL.n9 VTAIL.n8 67.5152
R95 VTAIL.n6 VTAIL.n5 67.5152
R96 VTAIL.n1 VTAIL.n0 67.5149
R97 VTAIL.n4 VTAIL.n3 67.5149
R98 VTAIL.n6 VTAIL.n4 25.6341
R99 VTAIL.n11 VTAIL.n10 22.5824
R100 VTAIL.n0 VTAIL.t3 3.91205
R101 VTAIL.n0 VTAIL.t1 3.91205
R102 VTAIL.n3 VTAIL.t9 3.91205
R103 VTAIL.n3 VTAIL.t8 3.91205
R104 VTAIL.n8 VTAIL.t6 3.91205
R105 VTAIL.n8 VTAIL.t11 3.91205
R106 VTAIL.n5 VTAIL.t4 3.91205
R107 VTAIL.n5 VTAIL.t2 3.91205
R108 VTAIL.n7 VTAIL.n6 3.05222
R109 VTAIL.n10 VTAIL.n9 3.05222
R110 VTAIL.n4 VTAIL.n2 3.05222
R111 VTAIL VTAIL.n11 2.2311
R112 VTAIL.n9 VTAIL.n7 1.99619
R113 VTAIL.n2 VTAIL.n1 1.99619
R114 VTAIL VTAIL.n1 0.821621
R115 VN.n34 VN.n33 161.3
R116 VN.n32 VN.n19 161.3
R117 VN.n31 VN.n30 161.3
R118 VN.n29 VN.n20 161.3
R119 VN.n28 VN.n27 161.3
R120 VN.n26 VN.n21 161.3
R121 VN.n25 VN.n24 161.3
R122 VN.n16 VN.n15 161.3
R123 VN.n14 VN.n1 161.3
R124 VN.n13 VN.n12 161.3
R125 VN.n11 VN.n2 161.3
R126 VN.n10 VN.n9 161.3
R127 VN.n8 VN.n3 161.3
R128 VN.n7 VN.n6 161.3
R129 VN.n5 VN.t5 95.2863
R130 VN.n23 VN.t1 95.2862
R131 VN.n17 VN.n0 75.8765
R132 VN.n35 VN.n18 75.8765
R133 VN.n4 VN.t3 62.3902
R134 VN.n0 VN.t2 62.3902
R135 VN.n22 VN.t4 62.3902
R136 VN.n18 VN.t0 62.3902
R137 VN.n5 VN.n4 62.0429
R138 VN.n23 VN.n22 62.0429
R139 VN VN.n35 48.5207
R140 VN.n13 VN.n2 42.4359
R141 VN.n31 VN.n20 42.4359
R142 VN.n9 VN.n2 38.5509
R143 VN.n27 VN.n20 38.5509
R144 VN.n8 VN.n7 24.4675
R145 VN.n9 VN.n8 24.4675
R146 VN.n14 VN.n13 24.4675
R147 VN.n15 VN.n14 24.4675
R148 VN.n27 VN.n26 24.4675
R149 VN.n26 VN.n25 24.4675
R150 VN.n33 VN.n32 24.4675
R151 VN.n32 VN.n31 24.4675
R152 VN.n15 VN.n0 14.1914
R153 VN.n33 VN.n18 14.1914
R154 VN.n7 VN.n4 12.234
R155 VN.n25 VN.n22 12.234
R156 VN.n24 VN.n23 4.18231
R157 VN.n6 VN.n5 4.18231
R158 VN.n35 VN.n34 0.354971
R159 VN.n17 VN.n16 0.354971
R160 VN VN.n17 0.26696
R161 VN.n34 VN.n19 0.189894
R162 VN.n30 VN.n19 0.189894
R163 VN.n30 VN.n29 0.189894
R164 VN.n29 VN.n28 0.189894
R165 VN.n28 VN.n21 0.189894
R166 VN.n24 VN.n21 0.189894
R167 VN.n6 VN.n3 0.189894
R168 VN.n10 VN.n3 0.189894
R169 VN.n11 VN.n10 0.189894
R170 VN.n12 VN.n11 0.189894
R171 VN.n12 VN.n1 0.189894
R172 VN.n16 VN.n1 0.189894
R173 VDD2.n1 VDD2.t0 90.3388
R174 VDD2.n2 VDD2.t5 88.1054
R175 VDD2.n1 VDD2.n0 84.9013
R176 VDD2 VDD2.n3 84.8985
R177 VDD2.n2 VDD2.n1 40.7972
R178 VDD2.n3 VDD2.t1 3.91205
R179 VDD2.n3 VDD2.t4 3.91205
R180 VDD2.n0 VDD2.t2 3.91205
R181 VDD2.n0 VDD2.t3 3.91205
R182 VDD2 VDD2.n2 2.34748
R183 B.n360 B.n359 585
R184 B.n358 B.n117 585
R185 B.n357 B.n356 585
R186 B.n355 B.n118 585
R187 B.n354 B.n353 585
R188 B.n352 B.n119 585
R189 B.n351 B.n350 585
R190 B.n349 B.n120 585
R191 B.n348 B.n347 585
R192 B.n346 B.n121 585
R193 B.n345 B.n344 585
R194 B.n343 B.n122 585
R195 B.n342 B.n341 585
R196 B.n340 B.n123 585
R197 B.n339 B.n338 585
R198 B.n337 B.n124 585
R199 B.n336 B.n335 585
R200 B.n334 B.n125 585
R201 B.n333 B.n332 585
R202 B.n331 B.n126 585
R203 B.n330 B.n329 585
R204 B.n328 B.n127 585
R205 B.n327 B.n326 585
R206 B.n325 B.n128 585
R207 B.n324 B.n323 585
R208 B.n322 B.n129 585
R209 B.n321 B.n320 585
R210 B.n319 B.n130 585
R211 B.n318 B.n317 585
R212 B.n316 B.n131 585
R213 B.n315 B.n314 585
R214 B.n313 B.n312 585
R215 B.n311 B.n135 585
R216 B.n310 B.n309 585
R217 B.n308 B.n136 585
R218 B.n307 B.n306 585
R219 B.n305 B.n137 585
R220 B.n304 B.n303 585
R221 B.n302 B.n138 585
R222 B.n301 B.n300 585
R223 B.n298 B.n139 585
R224 B.n297 B.n296 585
R225 B.n295 B.n142 585
R226 B.n294 B.n293 585
R227 B.n292 B.n143 585
R228 B.n291 B.n290 585
R229 B.n289 B.n144 585
R230 B.n288 B.n287 585
R231 B.n286 B.n145 585
R232 B.n285 B.n284 585
R233 B.n283 B.n146 585
R234 B.n282 B.n281 585
R235 B.n280 B.n147 585
R236 B.n279 B.n278 585
R237 B.n277 B.n148 585
R238 B.n276 B.n275 585
R239 B.n274 B.n149 585
R240 B.n273 B.n272 585
R241 B.n271 B.n150 585
R242 B.n270 B.n269 585
R243 B.n268 B.n151 585
R244 B.n267 B.n266 585
R245 B.n265 B.n152 585
R246 B.n264 B.n263 585
R247 B.n262 B.n153 585
R248 B.n261 B.n260 585
R249 B.n259 B.n154 585
R250 B.n258 B.n257 585
R251 B.n256 B.n155 585
R252 B.n255 B.n254 585
R253 B.n253 B.n156 585
R254 B.n361 B.n116 585
R255 B.n363 B.n362 585
R256 B.n364 B.n115 585
R257 B.n366 B.n365 585
R258 B.n367 B.n114 585
R259 B.n369 B.n368 585
R260 B.n370 B.n113 585
R261 B.n372 B.n371 585
R262 B.n373 B.n112 585
R263 B.n375 B.n374 585
R264 B.n376 B.n111 585
R265 B.n378 B.n377 585
R266 B.n379 B.n110 585
R267 B.n381 B.n380 585
R268 B.n382 B.n109 585
R269 B.n384 B.n383 585
R270 B.n385 B.n108 585
R271 B.n387 B.n386 585
R272 B.n388 B.n107 585
R273 B.n390 B.n389 585
R274 B.n391 B.n106 585
R275 B.n393 B.n392 585
R276 B.n394 B.n105 585
R277 B.n396 B.n395 585
R278 B.n397 B.n104 585
R279 B.n399 B.n398 585
R280 B.n400 B.n103 585
R281 B.n402 B.n401 585
R282 B.n403 B.n102 585
R283 B.n405 B.n404 585
R284 B.n406 B.n101 585
R285 B.n408 B.n407 585
R286 B.n409 B.n100 585
R287 B.n411 B.n410 585
R288 B.n412 B.n99 585
R289 B.n414 B.n413 585
R290 B.n415 B.n98 585
R291 B.n417 B.n416 585
R292 B.n418 B.n97 585
R293 B.n420 B.n419 585
R294 B.n421 B.n96 585
R295 B.n423 B.n422 585
R296 B.n424 B.n95 585
R297 B.n426 B.n425 585
R298 B.n427 B.n94 585
R299 B.n429 B.n428 585
R300 B.n430 B.n93 585
R301 B.n432 B.n431 585
R302 B.n433 B.n92 585
R303 B.n435 B.n434 585
R304 B.n436 B.n91 585
R305 B.n438 B.n437 585
R306 B.n439 B.n90 585
R307 B.n441 B.n440 585
R308 B.n442 B.n89 585
R309 B.n444 B.n443 585
R310 B.n445 B.n88 585
R311 B.n447 B.n446 585
R312 B.n448 B.n87 585
R313 B.n450 B.n449 585
R314 B.n451 B.n86 585
R315 B.n453 B.n452 585
R316 B.n454 B.n85 585
R317 B.n456 B.n455 585
R318 B.n457 B.n84 585
R319 B.n459 B.n458 585
R320 B.n460 B.n83 585
R321 B.n462 B.n461 585
R322 B.n463 B.n82 585
R323 B.n465 B.n464 585
R324 B.n466 B.n81 585
R325 B.n468 B.n467 585
R326 B.n469 B.n80 585
R327 B.n471 B.n470 585
R328 B.n472 B.n79 585
R329 B.n474 B.n473 585
R330 B.n475 B.n78 585
R331 B.n477 B.n476 585
R332 B.n478 B.n77 585
R333 B.n480 B.n479 585
R334 B.n481 B.n76 585
R335 B.n483 B.n482 585
R336 B.n484 B.n75 585
R337 B.n486 B.n485 585
R338 B.n487 B.n74 585
R339 B.n489 B.n488 585
R340 B.n490 B.n73 585
R341 B.n492 B.n491 585
R342 B.n493 B.n72 585
R343 B.n495 B.n494 585
R344 B.n496 B.n71 585
R345 B.n498 B.n497 585
R346 B.n499 B.n70 585
R347 B.n501 B.n500 585
R348 B.n502 B.n69 585
R349 B.n504 B.n503 585
R350 B.n505 B.n68 585
R351 B.n507 B.n506 585
R352 B.n508 B.n67 585
R353 B.n510 B.n509 585
R354 B.n618 B.n617 585
R355 B.n616 B.n27 585
R356 B.n615 B.n614 585
R357 B.n613 B.n28 585
R358 B.n612 B.n611 585
R359 B.n610 B.n29 585
R360 B.n609 B.n608 585
R361 B.n607 B.n30 585
R362 B.n606 B.n605 585
R363 B.n604 B.n31 585
R364 B.n603 B.n602 585
R365 B.n601 B.n32 585
R366 B.n600 B.n599 585
R367 B.n598 B.n33 585
R368 B.n597 B.n596 585
R369 B.n595 B.n34 585
R370 B.n594 B.n593 585
R371 B.n592 B.n35 585
R372 B.n591 B.n590 585
R373 B.n589 B.n36 585
R374 B.n588 B.n587 585
R375 B.n586 B.n37 585
R376 B.n585 B.n584 585
R377 B.n583 B.n38 585
R378 B.n582 B.n581 585
R379 B.n580 B.n39 585
R380 B.n579 B.n578 585
R381 B.n577 B.n40 585
R382 B.n576 B.n575 585
R383 B.n574 B.n41 585
R384 B.n573 B.n572 585
R385 B.n571 B.n570 585
R386 B.n569 B.n45 585
R387 B.n568 B.n567 585
R388 B.n566 B.n46 585
R389 B.n565 B.n564 585
R390 B.n563 B.n47 585
R391 B.n562 B.n561 585
R392 B.n560 B.n48 585
R393 B.n559 B.n558 585
R394 B.n556 B.n49 585
R395 B.n555 B.n554 585
R396 B.n553 B.n52 585
R397 B.n552 B.n551 585
R398 B.n550 B.n53 585
R399 B.n549 B.n548 585
R400 B.n547 B.n54 585
R401 B.n546 B.n545 585
R402 B.n544 B.n55 585
R403 B.n543 B.n542 585
R404 B.n541 B.n56 585
R405 B.n540 B.n539 585
R406 B.n538 B.n57 585
R407 B.n537 B.n536 585
R408 B.n535 B.n58 585
R409 B.n534 B.n533 585
R410 B.n532 B.n59 585
R411 B.n531 B.n530 585
R412 B.n529 B.n60 585
R413 B.n528 B.n527 585
R414 B.n526 B.n61 585
R415 B.n525 B.n524 585
R416 B.n523 B.n62 585
R417 B.n522 B.n521 585
R418 B.n520 B.n63 585
R419 B.n519 B.n518 585
R420 B.n517 B.n64 585
R421 B.n516 B.n515 585
R422 B.n514 B.n65 585
R423 B.n513 B.n512 585
R424 B.n511 B.n66 585
R425 B.n619 B.n26 585
R426 B.n621 B.n620 585
R427 B.n622 B.n25 585
R428 B.n624 B.n623 585
R429 B.n625 B.n24 585
R430 B.n627 B.n626 585
R431 B.n628 B.n23 585
R432 B.n630 B.n629 585
R433 B.n631 B.n22 585
R434 B.n633 B.n632 585
R435 B.n634 B.n21 585
R436 B.n636 B.n635 585
R437 B.n637 B.n20 585
R438 B.n639 B.n638 585
R439 B.n640 B.n19 585
R440 B.n642 B.n641 585
R441 B.n643 B.n18 585
R442 B.n645 B.n644 585
R443 B.n646 B.n17 585
R444 B.n648 B.n647 585
R445 B.n649 B.n16 585
R446 B.n651 B.n650 585
R447 B.n652 B.n15 585
R448 B.n654 B.n653 585
R449 B.n655 B.n14 585
R450 B.n657 B.n656 585
R451 B.n658 B.n13 585
R452 B.n660 B.n659 585
R453 B.n661 B.n12 585
R454 B.n663 B.n662 585
R455 B.n664 B.n11 585
R456 B.n666 B.n665 585
R457 B.n667 B.n10 585
R458 B.n669 B.n668 585
R459 B.n670 B.n9 585
R460 B.n672 B.n671 585
R461 B.n673 B.n8 585
R462 B.n675 B.n674 585
R463 B.n676 B.n7 585
R464 B.n678 B.n677 585
R465 B.n679 B.n6 585
R466 B.n681 B.n680 585
R467 B.n682 B.n5 585
R468 B.n684 B.n683 585
R469 B.n685 B.n4 585
R470 B.n687 B.n686 585
R471 B.n688 B.n3 585
R472 B.n690 B.n689 585
R473 B.n691 B.n0 585
R474 B.n2 B.n1 585
R475 B.n181 B.n180 585
R476 B.n183 B.n182 585
R477 B.n184 B.n179 585
R478 B.n186 B.n185 585
R479 B.n187 B.n178 585
R480 B.n189 B.n188 585
R481 B.n190 B.n177 585
R482 B.n192 B.n191 585
R483 B.n193 B.n176 585
R484 B.n195 B.n194 585
R485 B.n196 B.n175 585
R486 B.n198 B.n197 585
R487 B.n199 B.n174 585
R488 B.n201 B.n200 585
R489 B.n202 B.n173 585
R490 B.n204 B.n203 585
R491 B.n205 B.n172 585
R492 B.n207 B.n206 585
R493 B.n208 B.n171 585
R494 B.n210 B.n209 585
R495 B.n211 B.n170 585
R496 B.n213 B.n212 585
R497 B.n214 B.n169 585
R498 B.n216 B.n215 585
R499 B.n217 B.n168 585
R500 B.n219 B.n218 585
R501 B.n220 B.n167 585
R502 B.n222 B.n221 585
R503 B.n223 B.n166 585
R504 B.n225 B.n224 585
R505 B.n226 B.n165 585
R506 B.n228 B.n227 585
R507 B.n229 B.n164 585
R508 B.n231 B.n230 585
R509 B.n232 B.n163 585
R510 B.n234 B.n233 585
R511 B.n235 B.n162 585
R512 B.n237 B.n236 585
R513 B.n238 B.n161 585
R514 B.n240 B.n239 585
R515 B.n241 B.n160 585
R516 B.n243 B.n242 585
R517 B.n244 B.n159 585
R518 B.n246 B.n245 585
R519 B.n247 B.n158 585
R520 B.n249 B.n248 585
R521 B.n250 B.n157 585
R522 B.n252 B.n251 585
R523 B.n253 B.n252 550.159
R524 B.n361 B.n360 550.159
R525 B.n511 B.n510 550.159
R526 B.n619 B.n618 550.159
R527 B.n140 B.t0 271.202
R528 B.n132 B.t9 271.202
R529 B.n50 B.t3 271.202
R530 B.n42 B.t6 271.202
R531 B.n693 B.n692 256.663
R532 B.n692 B.n691 235.042
R533 B.n692 B.n2 235.042
R534 B.n132 B.t10 180.036
R535 B.n50 B.t5 180.036
R536 B.n140 B.t1 180.028
R537 B.n42 B.t8 180.028
R538 B.n254 B.n253 163.367
R539 B.n254 B.n155 163.367
R540 B.n258 B.n155 163.367
R541 B.n259 B.n258 163.367
R542 B.n260 B.n259 163.367
R543 B.n260 B.n153 163.367
R544 B.n264 B.n153 163.367
R545 B.n265 B.n264 163.367
R546 B.n266 B.n265 163.367
R547 B.n266 B.n151 163.367
R548 B.n270 B.n151 163.367
R549 B.n271 B.n270 163.367
R550 B.n272 B.n271 163.367
R551 B.n272 B.n149 163.367
R552 B.n276 B.n149 163.367
R553 B.n277 B.n276 163.367
R554 B.n278 B.n277 163.367
R555 B.n278 B.n147 163.367
R556 B.n282 B.n147 163.367
R557 B.n283 B.n282 163.367
R558 B.n284 B.n283 163.367
R559 B.n284 B.n145 163.367
R560 B.n288 B.n145 163.367
R561 B.n289 B.n288 163.367
R562 B.n290 B.n289 163.367
R563 B.n290 B.n143 163.367
R564 B.n294 B.n143 163.367
R565 B.n295 B.n294 163.367
R566 B.n296 B.n295 163.367
R567 B.n296 B.n139 163.367
R568 B.n301 B.n139 163.367
R569 B.n302 B.n301 163.367
R570 B.n303 B.n302 163.367
R571 B.n303 B.n137 163.367
R572 B.n307 B.n137 163.367
R573 B.n308 B.n307 163.367
R574 B.n309 B.n308 163.367
R575 B.n309 B.n135 163.367
R576 B.n313 B.n135 163.367
R577 B.n314 B.n313 163.367
R578 B.n314 B.n131 163.367
R579 B.n318 B.n131 163.367
R580 B.n319 B.n318 163.367
R581 B.n320 B.n319 163.367
R582 B.n320 B.n129 163.367
R583 B.n324 B.n129 163.367
R584 B.n325 B.n324 163.367
R585 B.n326 B.n325 163.367
R586 B.n326 B.n127 163.367
R587 B.n330 B.n127 163.367
R588 B.n331 B.n330 163.367
R589 B.n332 B.n331 163.367
R590 B.n332 B.n125 163.367
R591 B.n336 B.n125 163.367
R592 B.n337 B.n336 163.367
R593 B.n338 B.n337 163.367
R594 B.n338 B.n123 163.367
R595 B.n342 B.n123 163.367
R596 B.n343 B.n342 163.367
R597 B.n344 B.n343 163.367
R598 B.n344 B.n121 163.367
R599 B.n348 B.n121 163.367
R600 B.n349 B.n348 163.367
R601 B.n350 B.n349 163.367
R602 B.n350 B.n119 163.367
R603 B.n354 B.n119 163.367
R604 B.n355 B.n354 163.367
R605 B.n356 B.n355 163.367
R606 B.n356 B.n117 163.367
R607 B.n360 B.n117 163.367
R608 B.n510 B.n67 163.367
R609 B.n506 B.n67 163.367
R610 B.n506 B.n505 163.367
R611 B.n505 B.n504 163.367
R612 B.n504 B.n69 163.367
R613 B.n500 B.n69 163.367
R614 B.n500 B.n499 163.367
R615 B.n499 B.n498 163.367
R616 B.n498 B.n71 163.367
R617 B.n494 B.n71 163.367
R618 B.n494 B.n493 163.367
R619 B.n493 B.n492 163.367
R620 B.n492 B.n73 163.367
R621 B.n488 B.n73 163.367
R622 B.n488 B.n487 163.367
R623 B.n487 B.n486 163.367
R624 B.n486 B.n75 163.367
R625 B.n482 B.n75 163.367
R626 B.n482 B.n481 163.367
R627 B.n481 B.n480 163.367
R628 B.n480 B.n77 163.367
R629 B.n476 B.n77 163.367
R630 B.n476 B.n475 163.367
R631 B.n475 B.n474 163.367
R632 B.n474 B.n79 163.367
R633 B.n470 B.n79 163.367
R634 B.n470 B.n469 163.367
R635 B.n469 B.n468 163.367
R636 B.n468 B.n81 163.367
R637 B.n464 B.n81 163.367
R638 B.n464 B.n463 163.367
R639 B.n463 B.n462 163.367
R640 B.n462 B.n83 163.367
R641 B.n458 B.n83 163.367
R642 B.n458 B.n457 163.367
R643 B.n457 B.n456 163.367
R644 B.n456 B.n85 163.367
R645 B.n452 B.n85 163.367
R646 B.n452 B.n451 163.367
R647 B.n451 B.n450 163.367
R648 B.n450 B.n87 163.367
R649 B.n446 B.n87 163.367
R650 B.n446 B.n445 163.367
R651 B.n445 B.n444 163.367
R652 B.n444 B.n89 163.367
R653 B.n440 B.n89 163.367
R654 B.n440 B.n439 163.367
R655 B.n439 B.n438 163.367
R656 B.n438 B.n91 163.367
R657 B.n434 B.n91 163.367
R658 B.n434 B.n433 163.367
R659 B.n433 B.n432 163.367
R660 B.n432 B.n93 163.367
R661 B.n428 B.n93 163.367
R662 B.n428 B.n427 163.367
R663 B.n427 B.n426 163.367
R664 B.n426 B.n95 163.367
R665 B.n422 B.n95 163.367
R666 B.n422 B.n421 163.367
R667 B.n421 B.n420 163.367
R668 B.n420 B.n97 163.367
R669 B.n416 B.n97 163.367
R670 B.n416 B.n415 163.367
R671 B.n415 B.n414 163.367
R672 B.n414 B.n99 163.367
R673 B.n410 B.n99 163.367
R674 B.n410 B.n409 163.367
R675 B.n409 B.n408 163.367
R676 B.n408 B.n101 163.367
R677 B.n404 B.n101 163.367
R678 B.n404 B.n403 163.367
R679 B.n403 B.n402 163.367
R680 B.n402 B.n103 163.367
R681 B.n398 B.n103 163.367
R682 B.n398 B.n397 163.367
R683 B.n397 B.n396 163.367
R684 B.n396 B.n105 163.367
R685 B.n392 B.n105 163.367
R686 B.n392 B.n391 163.367
R687 B.n391 B.n390 163.367
R688 B.n390 B.n107 163.367
R689 B.n386 B.n107 163.367
R690 B.n386 B.n385 163.367
R691 B.n385 B.n384 163.367
R692 B.n384 B.n109 163.367
R693 B.n380 B.n109 163.367
R694 B.n380 B.n379 163.367
R695 B.n379 B.n378 163.367
R696 B.n378 B.n111 163.367
R697 B.n374 B.n111 163.367
R698 B.n374 B.n373 163.367
R699 B.n373 B.n372 163.367
R700 B.n372 B.n113 163.367
R701 B.n368 B.n113 163.367
R702 B.n368 B.n367 163.367
R703 B.n367 B.n366 163.367
R704 B.n366 B.n115 163.367
R705 B.n362 B.n115 163.367
R706 B.n362 B.n361 163.367
R707 B.n618 B.n27 163.367
R708 B.n614 B.n27 163.367
R709 B.n614 B.n613 163.367
R710 B.n613 B.n612 163.367
R711 B.n612 B.n29 163.367
R712 B.n608 B.n29 163.367
R713 B.n608 B.n607 163.367
R714 B.n607 B.n606 163.367
R715 B.n606 B.n31 163.367
R716 B.n602 B.n31 163.367
R717 B.n602 B.n601 163.367
R718 B.n601 B.n600 163.367
R719 B.n600 B.n33 163.367
R720 B.n596 B.n33 163.367
R721 B.n596 B.n595 163.367
R722 B.n595 B.n594 163.367
R723 B.n594 B.n35 163.367
R724 B.n590 B.n35 163.367
R725 B.n590 B.n589 163.367
R726 B.n589 B.n588 163.367
R727 B.n588 B.n37 163.367
R728 B.n584 B.n37 163.367
R729 B.n584 B.n583 163.367
R730 B.n583 B.n582 163.367
R731 B.n582 B.n39 163.367
R732 B.n578 B.n39 163.367
R733 B.n578 B.n577 163.367
R734 B.n577 B.n576 163.367
R735 B.n576 B.n41 163.367
R736 B.n572 B.n41 163.367
R737 B.n572 B.n571 163.367
R738 B.n571 B.n45 163.367
R739 B.n567 B.n45 163.367
R740 B.n567 B.n566 163.367
R741 B.n566 B.n565 163.367
R742 B.n565 B.n47 163.367
R743 B.n561 B.n47 163.367
R744 B.n561 B.n560 163.367
R745 B.n560 B.n559 163.367
R746 B.n559 B.n49 163.367
R747 B.n554 B.n49 163.367
R748 B.n554 B.n553 163.367
R749 B.n553 B.n552 163.367
R750 B.n552 B.n53 163.367
R751 B.n548 B.n53 163.367
R752 B.n548 B.n547 163.367
R753 B.n547 B.n546 163.367
R754 B.n546 B.n55 163.367
R755 B.n542 B.n55 163.367
R756 B.n542 B.n541 163.367
R757 B.n541 B.n540 163.367
R758 B.n540 B.n57 163.367
R759 B.n536 B.n57 163.367
R760 B.n536 B.n535 163.367
R761 B.n535 B.n534 163.367
R762 B.n534 B.n59 163.367
R763 B.n530 B.n59 163.367
R764 B.n530 B.n529 163.367
R765 B.n529 B.n528 163.367
R766 B.n528 B.n61 163.367
R767 B.n524 B.n61 163.367
R768 B.n524 B.n523 163.367
R769 B.n523 B.n522 163.367
R770 B.n522 B.n63 163.367
R771 B.n518 B.n63 163.367
R772 B.n518 B.n517 163.367
R773 B.n517 B.n516 163.367
R774 B.n516 B.n65 163.367
R775 B.n512 B.n65 163.367
R776 B.n512 B.n511 163.367
R777 B.n620 B.n619 163.367
R778 B.n620 B.n25 163.367
R779 B.n624 B.n25 163.367
R780 B.n625 B.n624 163.367
R781 B.n626 B.n625 163.367
R782 B.n626 B.n23 163.367
R783 B.n630 B.n23 163.367
R784 B.n631 B.n630 163.367
R785 B.n632 B.n631 163.367
R786 B.n632 B.n21 163.367
R787 B.n636 B.n21 163.367
R788 B.n637 B.n636 163.367
R789 B.n638 B.n637 163.367
R790 B.n638 B.n19 163.367
R791 B.n642 B.n19 163.367
R792 B.n643 B.n642 163.367
R793 B.n644 B.n643 163.367
R794 B.n644 B.n17 163.367
R795 B.n648 B.n17 163.367
R796 B.n649 B.n648 163.367
R797 B.n650 B.n649 163.367
R798 B.n650 B.n15 163.367
R799 B.n654 B.n15 163.367
R800 B.n655 B.n654 163.367
R801 B.n656 B.n655 163.367
R802 B.n656 B.n13 163.367
R803 B.n660 B.n13 163.367
R804 B.n661 B.n660 163.367
R805 B.n662 B.n661 163.367
R806 B.n662 B.n11 163.367
R807 B.n666 B.n11 163.367
R808 B.n667 B.n666 163.367
R809 B.n668 B.n667 163.367
R810 B.n668 B.n9 163.367
R811 B.n672 B.n9 163.367
R812 B.n673 B.n672 163.367
R813 B.n674 B.n673 163.367
R814 B.n674 B.n7 163.367
R815 B.n678 B.n7 163.367
R816 B.n679 B.n678 163.367
R817 B.n680 B.n679 163.367
R818 B.n680 B.n5 163.367
R819 B.n684 B.n5 163.367
R820 B.n685 B.n684 163.367
R821 B.n686 B.n685 163.367
R822 B.n686 B.n3 163.367
R823 B.n690 B.n3 163.367
R824 B.n691 B.n690 163.367
R825 B.n181 B.n2 163.367
R826 B.n182 B.n181 163.367
R827 B.n182 B.n179 163.367
R828 B.n186 B.n179 163.367
R829 B.n187 B.n186 163.367
R830 B.n188 B.n187 163.367
R831 B.n188 B.n177 163.367
R832 B.n192 B.n177 163.367
R833 B.n193 B.n192 163.367
R834 B.n194 B.n193 163.367
R835 B.n194 B.n175 163.367
R836 B.n198 B.n175 163.367
R837 B.n199 B.n198 163.367
R838 B.n200 B.n199 163.367
R839 B.n200 B.n173 163.367
R840 B.n204 B.n173 163.367
R841 B.n205 B.n204 163.367
R842 B.n206 B.n205 163.367
R843 B.n206 B.n171 163.367
R844 B.n210 B.n171 163.367
R845 B.n211 B.n210 163.367
R846 B.n212 B.n211 163.367
R847 B.n212 B.n169 163.367
R848 B.n216 B.n169 163.367
R849 B.n217 B.n216 163.367
R850 B.n218 B.n217 163.367
R851 B.n218 B.n167 163.367
R852 B.n222 B.n167 163.367
R853 B.n223 B.n222 163.367
R854 B.n224 B.n223 163.367
R855 B.n224 B.n165 163.367
R856 B.n228 B.n165 163.367
R857 B.n229 B.n228 163.367
R858 B.n230 B.n229 163.367
R859 B.n230 B.n163 163.367
R860 B.n234 B.n163 163.367
R861 B.n235 B.n234 163.367
R862 B.n236 B.n235 163.367
R863 B.n236 B.n161 163.367
R864 B.n240 B.n161 163.367
R865 B.n241 B.n240 163.367
R866 B.n242 B.n241 163.367
R867 B.n242 B.n159 163.367
R868 B.n246 B.n159 163.367
R869 B.n247 B.n246 163.367
R870 B.n248 B.n247 163.367
R871 B.n248 B.n157 163.367
R872 B.n252 B.n157 163.367
R873 B.n133 B.t11 111.382
R874 B.n51 B.t4 111.382
R875 B.n141 B.t2 111.374
R876 B.n43 B.t7 111.374
R877 B.n141 B.n140 68.655
R878 B.n133 B.n132 68.655
R879 B.n51 B.n50 68.655
R880 B.n43 B.n42 68.655
R881 B.n299 B.n141 59.5399
R882 B.n134 B.n133 59.5399
R883 B.n557 B.n51 59.5399
R884 B.n44 B.n43 59.5399
R885 B.n359 B.n116 35.7468
R886 B.n617 B.n26 35.7468
R887 B.n509 B.n66 35.7468
R888 B.n251 B.n156 35.7468
R889 B B.n693 18.0485
R890 B.n621 B.n26 10.6151
R891 B.n622 B.n621 10.6151
R892 B.n623 B.n622 10.6151
R893 B.n623 B.n24 10.6151
R894 B.n627 B.n24 10.6151
R895 B.n628 B.n627 10.6151
R896 B.n629 B.n628 10.6151
R897 B.n629 B.n22 10.6151
R898 B.n633 B.n22 10.6151
R899 B.n634 B.n633 10.6151
R900 B.n635 B.n634 10.6151
R901 B.n635 B.n20 10.6151
R902 B.n639 B.n20 10.6151
R903 B.n640 B.n639 10.6151
R904 B.n641 B.n640 10.6151
R905 B.n641 B.n18 10.6151
R906 B.n645 B.n18 10.6151
R907 B.n646 B.n645 10.6151
R908 B.n647 B.n646 10.6151
R909 B.n647 B.n16 10.6151
R910 B.n651 B.n16 10.6151
R911 B.n652 B.n651 10.6151
R912 B.n653 B.n652 10.6151
R913 B.n653 B.n14 10.6151
R914 B.n657 B.n14 10.6151
R915 B.n658 B.n657 10.6151
R916 B.n659 B.n658 10.6151
R917 B.n659 B.n12 10.6151
R918 B.n663 B.n12 10.6151
R919 B.n664 B.n663 10.6151
R920 B.n665 B.n664 10.6151
R921 B.n665 B.n10 10.6151
R922 B.n669 B.n10 10.6151
R923 B.n670 B.n669 10.6151
R924 B.n671 B.n670 10.6151
R925 B.n671 B.n8 10.6151
R926 B.n675 B.n8 10.6151
R927 B.n676 B.n675 10.6151
R928 B.n677 B.n676 10.6151
R929 B.n677 B.n6 10.6151
R930 B.n681 B.n6 10.6151
R931 B.n682 B.n681 10.6151
R932 B.n683 B.n682 10.6151
R933 B.n683 B.n4 10.6151
R934 B.n687 B.n4 10.6151
R935 B.n688 B.n687 10.6151
R936 B.n689 B.n688 10.6151
R937 B.n689 B.n0 10.6151
R938 B.n617 B.n616 10.6151
R939 B.n616 B.n615 10.6151
R940 B.n615 B.n28 10.6151
R941 B.n611 B.n28 10.6151
R942 B.n611 B.n610 10.6151
R943 B.n610 B.n609 10.6151
R944 B.n609 B.n30 10.6151
R945 B.n605 B.n30 10.6151
R946 B.n605 B.n604 10.6151
R947 B.n604 B.n603 10.6151
R948 B.n603 B.n32 10.6151
R949 B.n599 B.n32 10.6151
R950 B.n599 B.n598 10.6151
R951 B.n598 B.n597 10.6151
R952 B.n597 B.n34 10.6151
R953 B.n593 B.n34 10.6151
R954 B.n593 B.n592 10.6151
R955 B.n592 B.n591 10.6151
R956 B.n591 B.n36 10.6151
R957 B.n587 B.n36 10.6151
R958 B.n587 B.n586 10.6151
R959 B.n586 B.n585 10.6151
R960 B.n585 B.n38 10.6151
R961 B.n581 B.n38 10.6151
R962 B.n581 B.n580 10.6151
R963 B.n580 B.n579 10.6151
R964 B.n579 B.n40 10.6151
R965 B.n575 B.n40 10.6151
R966 B.n575 B.n574 10.6151
R967 B.n574 B.n573 10.6151
R968 B.n570 B.n569 10.6151
R969 B.n569 B.n568 10.6151
R970 B.n568 B.n46 10.6151
R971 B.n564 B.n46 10.6151
R972 B.n564 B.n563 10.6151
R973 B.n563 B.n562 10.6151
R974 B.n562 B.n48 10.6151
R975 B.n558 B.n48 10.6151
R976 B.n556 B.n555 10.6151
R977 B.n555 B.n52 10.6151
R978 B.n551 B.n52 10.6151
R979 B.n551 B.n550 10.6151
R980 B.n550 B.n549 10.6151
R981 B.n549 B.n54 10.6151
R982 B.n545 B.n54 10.6151
R983 B.n545 B.n544 10.6151
R984 B.n544 B.n543 10.6151
R985 B.n543 B.n56 10.6151
R986 B.n539 B.n56 10.6151
R987 B.n539 B.n538 10.6151
R988 B.n538 B.n537 10.6151
R989 B.n537 B.n58 10.6151
R990 B.n533 B.n58 10.6151
R991 B.n533 B.n532 10.6151
R992 B.n532 B.n531 10.6151
R993 B.n531 B.n60 10.6151
R994 B.n527 B.n60 10.6151
R995 B.n527 B.n526 10.6151
R996 B.n526 B.n525 10.6151
R997 B.n525 B.n62 10.6151
R998 B.n521 B.n62 10.6151
R999 B.n521 B.n520 10.6151
R1000 B.n520 B.n519 10.6151
R1001 B.n519 B.n64 10.6151
R1002 B.n515 B.n64 10.6151
R1003 B.n515 B.n514 10.6151
R1004 B.n514 B.n513 10.6151
R1005 B.n513 B.n66 10.6151
R1006 B.n509 B.n508 10.6151
R1007 B.n508 B.n507 10.6151
R1008 B.n507 B.n68 10.6151
R1009 B.n503 B.n68 10.6151
R1010 B.n503 B.n502 10.6151
R1011 B.n502 B.n501 10.6151
R1012 B.n501 B.n70 10.6151
R1013 B.n497 B.n70 10.6151
R1014 B.n497 B.n496 10.6151
R1015 B.n496 B.n495 10.6151
R1016 B.n495 B.n72 10.6151
R1017 B.n491 B.n72 10.6151
R1018 B.n491 B.n490 10.6151
R1019 B.n490 B.n489 10.6151
R1020 B.n489 B.n74 10.6151
R1021 B.n485 B.n74 10.6151
R1022 B.n485 B.n484 10.6151
R1023 B.n484 B.n483 10.6151
R1024 B.n483 B.n76 10.6151
R1025 B.n479 B.n76 10.6151
R1026 B.n479 B.n478 10.6151
R1027 B.n478 B.n477 10.6151
R1028 B.n477 B.n78 10.6151
R1029 B.n473 B.n78 10.6151
R1030 B.n473 B.n472 10.6151
R1031 B.n472 B.n471 10.6151
R1032 B.n471 B.n80 10.6151
R1033 B.n467 B.n80 10.6151
R1034 B.n467 B.n466 10.6151
R1035 B.n466 B.n465 10.6151
R1036 B.n465 B.n82 10.6151
R1037 B.n461 B.n82 10.6151
R1038 B.n461 B.n460 10.6151
R1039 B.n460 B.n459 10.6151
R1040 B.n459 B.n84 10.6151
R1041 B.n455 B.n84 10.6151
R1042 B.n455 B.n454 10.6151
R1043 B.n454 B.n453 10.6151
R1044 B.n453 B.n86 10.6151
R1045 B.n449 B.n86 10.6151
R1046 B.n449 B.n448 10.6151
R1047 B.n448 B.n447 10.6151
R1048 B.n447 B.n88 10.6151
R1049 B.n443 B.n88 10.6151
R1050 B.n443 B.n442 10.6151
R1051 B.n442 B.n441 10.6151
R1052 B.n441 B.n90 10.6151
R1053 B.n437 B.n90 10.6151
R1054 B.n437 B.n436 10.6151
R1055 B.n436 B.n435 10.6151
R1056 B.n435 B.n92 10.6151
R1057 B.n431 B.n92 10.6151
R1058 B.n431 B.n430 10.6151
R1059 B.n430 B.n429 10.6151
R1060 B.n429 B.n94 10.6151
R1061 B.n425 B.n94 10.6151
R1062 B.n425 B.n424 10.6151
R1063 B.n424 B.n423 10.6151
R1064 B.n423 B.n96 10.6151
R1065 B.n419 B.n96 10.6151
R1066 B.n419 B.n418 10.6151
R1067 B.n418 B.n417 10.6151
R1068 B.n417 B.n98 10.6151
R1069 B.n413 B.n98 10.6151
R1070 B.n413 B.n412 10.6151
R1071 B.n412 B.n411 10.6151
R1072 B.n411 B.n100 10.6151
R1073 B.n407 B.n100 10.6151
R1074 B.n407 B.n406 10.6151
R1075 B.n406 B.n405 10.6151
R1076 B.n405 B.n102 10.6151
R1077 B.n401 B.n102 10.6151
R1078 B.n401 B.n400 10.6151
R1079 B.n400 B.n399 10.6151
R1080 B.n399 B.n104 10.6151
R1081 B.n395 B.n104 10.6151
R1082 B.n395 B.n394 10.6151
R1083 B.n394 B.n393 10.6151
R1084 B.n393 B.n106 10.6151
R1085 B.n389 B.n106 10.6151
R1086 B.n389 B.n388 10.6151
R1087 B.n388 B.n387 10.6151
R1088 B.n387 B.n108 10.6151
R1089 B.n383 B.n108 10.6151
R1090 B.n383 B.n382 10.6151
R1091 B.n382 B.n381 10.6151
R1092 B.n381 B.n110 10.6151
R1093 B.n377 B.n110 10.6151
R1094 B.n377 B.n376 10.6151
R1095 B.n376 B.n375 10.6151
R1096 B.n375 B.n112 10.6151
R1097 B.n371 B.n112 10.6151
R1098 B.n371 B.n370 10.6151
R1099 B.n370 B.n369 10.6151
R1100 B.n369 B.n114 10.6151
R1101 B.n365 B.n114 10.6151
R1102 B.n365 B.n364 10.6151
R1103 B.n364 B.n363 10.6151
R1104 B.n363 B.n116 10.6151
R1105 B.n180 B.n1 10.6151
R1106 B.n183 B.n180 10.6151
R1107 B.n184 B.n183 10.6151
R1108 B.n185 B.n184 10.6151
R1109 B.n185 B.n178 10.6151
R1110 B.n189 B.n178 10.6151
R1111 B.n190 B.n189 10.6151
R1112 B.n191 B.n190 10.6151
R1113 B.n191 B.n176 10.6151
R1114 B.n195 B.n176 10.6151
R1115 B.n196 B.n195 10.6151
R1116 B.n197 B.n196 10.6151
R1117 B.n197 B.n174 10.6151
R1118 B.n201 B.n174 10.6151
R1119 B.n202 B.n201 10.6151
R1120 B.n203 B.n202 10.6151
R1121 B.n203 B.n172 10.6151
R1122 B.n207 B.n172 10.6151
R1123 B.n208 B.n207 10.6151
R1124 B.n209 B.n208 10.6151
R1125 B.n209 B.n170 10.6151
R1126 B.n213 B.n170 10.6151
R1127 B.n214 B.n213 10.6151
R1128 B.n215 B.n214 10.6151
R1129 B.n215 B.n168 10.6151
R1130 B.n219 B.n168 10.6151
R1131 B.n220 B.n219 10.6151
R1132 B.n221 B.n220 10.6151
R1133 B.n221 B.n166 10.6151
R1134 B.n225 B.n166 10.6151
R1135 B.n226 B.n225 10.6151
R1136 B.n227 B.n226 10.6151
R1137 B.n227 B.n164 10.6151
R1138 B.n231 B.n164 10.6151
R1139 B.n232 B.n231 10.6151
R1140 B.n233 B.n232 10.6151
R1141 B.n233 B.n162 10.6151
R1142 B.n237 B.n162 10.6151
R1143 B.n238 B.n237 10.6151
R1144 B.n239 B.n238 10.6151
R1145 B.n239 B.n160 10.6151
R1146 B.n243 B.n160 10.6151
R1147 B.n244 B.n243 10.6151
R1148 B.n245 B.n244 10.6151
R1149 B.n245 B.n158 10.6151
R1150 B.n249 B.n158 10.6151
R1151 B.n250 B.n249 10.6151
R1152 B.n251 B.n250 10.6151
R1153 B.n255 B.n156 10.6151
R1154 B.n256 B.n255 10.6151
R1155 B.n257 B.n256 10.6151
R1156 B.n257 B.n154 10.6151
R1157 B.n261 B.n154 10.6151
R1158 B.n262 B.n261 10.6151
R1159 B.n263 B.n262 10.6151
R1160 B.n263 B.n152 10.6151
R1161 B.n267 B.n152 10.6151
R1162 B.n268 B.n267 10.6151
R1163 B.n269 B.n268 10.6151
R1164 B.n269 B.n150 10.6151
R1165 B.n273 B.n150 10.6151
R1166 B.n274 B.n273 10.6151
R1167 B.n275 B.n274 10.6151
R1168 B.n275 B.n148 10.6151
R1169 B.n279 B.n148 10.6151
R1170 B.n280 B.n279 10.6151
R1171 B.n281 B.n280 10.6151
R1172 B.n281 B.n146 10.6151
R1173 B.n285 B.n146 10.6151
R1174 B.n286 B.n285 10.6151
R1175 B.n287 B.n286 10.6151
R1176 B.n287 B.n144 10.6151
R1177 B.n291 B.n144 10.6151
R1178 B.n292 B.n291 10.6151
R1179 B.n293 B.n292 10.6151
R1180 B.n293 B.n142 10.6151
R1181 B.n297 B.n142 10.6151
R1182 B.n298 B.n297 10.6151
R1183 B.n300 B.n138 10.6151
R1184 B.n304 B.n138 10.6151
R1185 B.n305 B.n304 10.6151
R1186 B.n306 B.n305 10.6151
R1187 B.n306 B.n136 10.6151
R1188 B.n310 B.n136 10.6151
R1189 B.n311 B.n310 10.6151
R1190 B.n312 B.n311 10.6151
R1191 B.n316 B.n315 10.6151
R1192 B.n317 B.n316 10.6151
R1193 B.n317 B.n130 10.6151
R1194 B.n321 B.n130 10.6151
R1195 B.n322 B.n321 10.6151
R1196 B.n323 B.n322 10.6151
R1197 B.n323 B.n128 10.6151
R1198 B.n327 B.n128 10.6151
R1199 B.n328 B.n327 10.6151
R1200 B.n329 B.n328 10.6151
R1201 B.n329 B.n126 10.6151
R1202 B.n333 B.n126 10.6151
R1203 B.n334 B.n333 10.6151
R1204 B.n335 B.n334 10.6151
R1205 B.n335 B.n124 10.6151
R1206 B.n339 B.n124 10.6151
R1207 B.n340 B.n339 10.6151
R1208 B.n341 B.n340 10.6151
R1209 B.n341 B.n122 10.6151
R1210 B.n345 B.n122 10.6151
R1211 B.n346 B.n345 10.6151
R1212 B.n347 B.n346 10.6151
R1213 B.n347 B.n120 10.6151
R1214 B.n351 B.n120 10.6151
R1215 B.n352 B.n351 10.6151
R1216 B.n353 B.n352 10.6151
R1217 B.n353 B.n118 10.6151
R1218 B.n357 B.n118 10.6151
R1219 B.n358 B.n357 10.6151
R1220 B.n359 B.n358 10.6151
R1221 B.n693 B.n0 8.11757
R1222 B.n693 B.n1 8.11757
R1223 B.n570 B.n44 6.5566
R1224 B.n558 B.n557 6.5566
R1225 B.n300 B.n299 6.5566
R1226 B.n312 B.n134 6.5566
R1227 B.n573 B.n44 4.05904
R1228 B.n557 B.n556 4.05904
R1229 B.n299 B.n298 4.05904
R1230 B.n315 B.n134 4.05904
C0 w_n3802_n2630# VDD1 2.18279f
C1 VN VDD1 0.151398f
C2 VDD2 VDD1 1.64333f
C3 w_n3802_n2630# B 9.48416f
C4 VP VDD1 5.30939f
C5 VN B 1.25255f
C6 VTAIL VDD1 6.66185f
C7 VN w_n3802_n2630# 7.291669f
C8 VDD2 B 2.04592f
C9 VDD2 w_n3802_n2630# 2.28735f
C10 VN VDD2 4.95371f
C11 VP B 2.07914f
C12 VTAIL B 3.0721f
C13 VP w_n3802_n2630# 7.78492f
C14 VP VN 6.83898f
C15 VTAIL w_n3802_n2630# 2.5163f
C16 VN VTAIL 5.43035f
C17 VP VDD2 0.509618f
C18 VDD2 VTAIL 6.718029f
C19 VP VTAIL 5.44455f
C20 B VDD1 1.9572f
C21 VDD2 VSUBS 1.966607f
C22 VDD1 VSUBS 2.356054f
C23 VTAIL VSUBS 1.185358f
C24 VN VSUBS 6.35798f
C25 VP VSUBS 3.285486f
C26 B VSUBS 4.929176f
C27 w_n3802_n2630# VSUBS 0.12396p
C28 B.n0 VSUBS 0.007855f
C29 B.n1 VSUBS 0.007855f
C30 B.n2 VSUBS 0.011618f
C31 B.n3 VSUBS 0.008903f
C32 B.n4 VSUBS 0.008903f
C33 B.n5 VSUBS 0.008903f
C34 B.n6 VSUBS 0.008903f
C35 B.n7 VSUBS 0.008903f
C36 B.n8 VSUBS 0.008903f
C37 B.n9 VSUBS 0.008903f
C38 B.n10 VSUBS 0.008903f
C39 B.n11 VSUBS 0.008903f
C40 B.n12 VSUBS 0.008903f
C41 B.n13 VSUBS 0.008903f
C42 B.n14 VSUBS 0.008903f
C43 B.n15 VSUBS 0.008903f
C44 B.n16 VSUBS 0.008903f
C45 B.n17 VSUBS 0.008903f
C46 B.n18 VSUBS 0.008903f
C47 B.n19 VSUBS 0.008903f
C48 B.n20 VSUBS 0.008903f
C49 B.n21 VSUBS 0.008903f
C50 B.n22 VSUBS 0.008903f
C51 B.n23 VSUBS 0.008903f
C52 B.n24 VSUBS 0.008903f
C53 B.n25 VSUBS 0.008903f
C54 B.n26 VSUBS 0.021505f
C55 B.n27 VSUBS 0.008903f
C56 B.n28 VSUBS 0.008903f
C57 B.n29 VSUBS 0.008903f
C58 B.n30 VSUBS 0.008903f
C59 B.n31 VSUBS 0.008903f
C60 B.n32 VSUBS 0.008903f
C61 B.n33 VSUBS 0.008903f
C62 B.n34 VSUBS 0.008903f
C63 B.n35 VSUBS 0.008903f
C64 B.n36 VSUBS 0.008903f
C65 B.n37 VSUBS 0.008903f
C66 B.n38 VSUBS 0.008903f
C67 B.n39 VSUBS 0.008903f
C68 B.n40 VSUBS 0.008903f
C69 B.n41 VSUBS 0.008903f
C70 B.t7 VSUBS 0.328145f
C71 B.t8 VSUBS 0.359175f
C72 B.t6 VSUBS 1.59697f
C73 B.n42 VSUBS 0.201223f
C74 B.n43 VSUBS 0.094065f
C75 B.n44 VSUBS 0.020627f
C76 B.n45 VSUBS 0.008903f
C77 B.n46 VSUBS 0.008903f
C78 B.n47 VSUBS 0.008903f
C79 B.n48 VSUBS 0.008903f
C80 B.n49 VSUBS 0.008903f
C81 B.t4 VSUBS 0.328142f
C82 B.t5 VSUBS 0.359172f
C83 B.t3 VSUBS 1.59697f
C84 B.n50 VSUBS 0.201226f
C85 B.n51 VSUBS 0.094068f
C86 B.n52 VSUBS 0.008903f
C87 B.n53 VSUBS 0.008903f
C88 B.n54 VSUBS 0.008903f
C89 B.n55 VSUBS 0.008903f
C90 B.n56 VSUBS 0.008903f
C91 B.n57 VSUBS 0.008903f
C92 B.n58 VSUBS 0.008903f
C93 B.n59 VSUBS 0.008903f
C94 B.n60 VSUBS 0.008903f
C95 B.n61 VSUBS 0.008903f
C96 B.n62 VSUBS 0.008903f
C97 B.n63 VSUBS 0.008903f
C98 B.n64 VSUBS 0.008903f
C99 B.n65 VSUBS 0.008903f
C100 B.n66 VSUBS 0.022747f
C101 B.n67 VSUBS 0.008903f
C102 B.n68 VSUBS 0.008903f
C103 B.n69 VSUBS 0.008903f
C104 B.n70 VSUBS 0.008903f
C105 B.n71 VSUBS 0.008903f
C106 B.n72 VSUBS 0.008903f
C107 B.n73 VSUBS 0.008903f
C108 B.n74 VSUBS 0.008903f
C109 B.n75 VSUBS 0.008903f
C110 B.n76 VSUBS 0.008903f
C111 B.n77 VSUBS 0.008903f
C112 B.n78 VSUBS 0.008903f
C113 B.n79 VSUBS 0.008903f
C114 B.n80 VSUBS 0.008903f
C115 B.n81 VSUBS 0.008903f
C116 B.n82 VSUBS 0.008903f
C117 B.n83 VSUBS 0.008903f
C118 B.n84 VSUBS 0.008903f
C119 B.n85 VSUBS 0.008903f
C120 B.n86 VSUBS 0.008903f
C121 B.n87 VSUBS 0.008903f
C122 B.n88 VSUBS 0.008903f
C123 B.n89 VSUBS 0.008903f
C124 B.n90 VSUBS 0.008903f
C125 B.n91 VSUBS 0.008903f
C126 B.n92 VSUBS 0.008903f
C127 B.n93 VSUBS 0.008903f
C128 B.n94 VSUBS 0.008903f
C129 B.n95 VSUBS 0.008903f
C130 B.n96 VSUBS 0.008903f
C131 B.n97 VSUBS 0.008903f
C132 B.n98 VSUBS 0.008903f
C133 B.n99 VSUBS 0.008903f
C134 B.n100 VSUBS 0.008903f
C135 B.n101 VSUBS 0.008903f
C136 B.n102 VSUBS 0.008903f
C137 B.n103 VSUBS 0.008903f
C138 B.n104 VSUBS 0.008903f
C139 B.n105 VSUBS 0.008903f
C140 B.n106 VSUBS 0.008903f
C141 B.n107 VSUBS 0.008903f
C142 B.n108 VSUBS 0.008903f
C143 B.n109 VSUBS 0.008903f
C144 B.n110 VSUBS 0.008903f
C145 B.n111 VSUBS 0.008903f
C146 B.n112 VSUBS 0.008903f
C147 B.n113 VSUBS 0.008903f
C148 B.n114 VSUBS 0.008903f
C149 B.n115 VSUBS 0.008903f
C150 B.n116 VSUBS 0.022466f
C151 B.n117 VSUBS 0.008903f
C152 B.n118 VSUBS 0.008903f
C153 B.n119 VSUBS 0.008903f
C154 B.n120 VSUBS 0.008903f
C155 B.n121 VSUBS 0.008903f
C156 B.n122 VSUBS 0.008903f
C157 B.n123 VSUBS 0.008903f
C158 B.n124 VSUBS 0.008903f
C159 B.n125 VSUBS 0.008903f
C160 B.n126 VSUBS 0.008903f
C161 B.n127 VSUBS 0.008903f
C162 B.n128 VSUBS 0.008903f
C163 B.n129 VSUBS 0.008903f
C164 B.n130 VSUBS 0.008903f
C165 B.n131 VSUBS 0.008903f
C166 B.t11 VSUBS 0.328142f
C167 B.t10 VSUBS 0.359172f
C168 B.t9 VSUBS 1.59697f
C169 B.n132 VSUBS 0.201226f
C170 B.n133 VSUBS 0.094068f
C171 B.n134 VSUBS 0.020627f
C172 B.n135 VSUBS 0.008903f
C173 B.n136 VSUBS 0.008903f
C174 B.n137 VSUBS 0.008903f
C175 B.n138 VSUBS 0.008903f
C176 B.n139 VSUBS 0.008903f
C177 B.t2 VSUBS 0.328145f
C178 B.t1 VSUBS 0.359175f
C179 B.t0 VSUBS 1.59697f
C180 B.n140 VSUBS 0.201223f
C181 B.n141 VSUBS 0.094065f
C182 B.n142 VSUBS 0.008903f
C183 B.n143 VSUBS 0.008903f
C184 B.n144 VSUBS 0.008903f
C185 B.n145 VSUBS 0.008903f
C186 B.n146 VSUBS 0.008903f
C187 B.n147 VSUBS 0.008903f
C188 B.n148 VSUBS 0.008903f
C189 B.n149 VSUBS 0.008903f
C190 B.n150 VSUBS 0.008903f
C191 B.n151 VSUBS 0.008903f
C192 B.n152 VSUBS 0.008903f
C193 B.n153 VSUBS 0.008903f
C194 B.n154 VSUBS 0.008903f
C195 B.n155 VSUBS 0.008903f
C196 B.n156 VSUBS 0.022747f
C197 B.n157 VSUBS 0.008903f
C198 B.n158 VSUBS 0.008903f
C199 B.n159 VSUBS 0.008903f
C200 B.n160 VSUBS 0.008903f
C201 B.n161 VSUBS 0.008903f
C202 B.n162 VSUBS 0.008903f
C203 B.n163 VSUBS 0.008903f
C204 B.n164 VSUBS 0.008903f
C205 B.n165 VSUBS 0.008903f
C206 B.n166 VSUBS 0.008903f
C207 B.n167 VSUBS 0.008903f
C208 B.n168 VSUBS 0.008903f
C209 B.n169 VSUBS 0.008903f
C210 B.n170 VSUBS 0.008903f
C211 B.n171 VSUBS 0.008903f
C212 B.n172 VSUBS 0.008903f
C213 B.n173 VSUBS 0.008903f
C214 B.n174 VSUBS 0.008903f
C215 B.n175 VSUBS 0.008903f
C216 B.n176 VSUBS 0.008903f
C217 B.n177 VSUBS 0.008903f
C218 B.n178 VSUBS 0.008903f
C219 B.n179 VSUBS 0.008903f
C220 B.n180 VSUBS 0.008903f
C221 B.n181 VSUBS 0.008903f
C222 B.n182 VSUBS 0.008903f
C223 B.n183 VSUBS 0.008903f
C224 B.n184 VSUBS 0.008903f
C225 B.n185 VSUBS 0.008903f
C226 B.n186 VSUBS 0.008903f
C227 B.n187 VSUBS 0.008903f
C228 B.n188 VSUBS 0.008903f
C229 B.n189 VSUBS 0.008903f
C230 B.n190 VSUBS 0.008903f
C231 B.n191 VSUBS 0.008903f
C232 B.n192 VSUBS 0.008903f
C233 B.n193 VSUBS 0.008903f
C234 B.n194 VSUBS 0.008903f
C235 B.n195 VSUBS 0.008903f
C236 B.n196 VSUBS 0.008903f
C237 B.n197 VSUBS 0.008903f
C238 B.n198 VSUBS 0.008903f
C239 B.n199 VSUBS 0.008903f
C240 B.n200 VSUBS 0.008903f
C241 B.n201 VSUBS 0.008903f
C242 B.n202 VSUBS 0.008903f
C243 B.n203 VSUBS 0.008903f
C244 B.n204 VSUBS 0.008903f
C245 B.n205 VSUBS 0.008903f
C246 B.n206 VSUBS 0.008903f
C247 B.n207 VSUBS 0.008903f
C248 B.n208 VSUBS 0.008903f
C249 B.n209 VSUBS 0.008903f
C250 B.n210 VSUBS 0.008903f
C251 B.n211 VSUBS 0.008903f
C252 B.n212 VSUBS 0.008903f
C253 B.n213 VSUBS 0.008903f
C254 B.n214 VSUBS 0.008903f
C255 B.n215 VSUBS 0.008903f
C256 B.n216 VSUBS 0.008903f
C257 B.n217 VSUBS 0.008903f
C258 B.n218 VSUBS 0.008903f
C259 B.n219 VSUBS 0.008903f
C260 B.n220 VSUBS 0.008903f
C261 B.n221 VSUBS 0.008903f
C262 B.n222 VSUBS 0.008903f
C263 B.n223 VSUBS 0.008903f
C264 B.n224 VSUBS 0.008903f
C265 B.n225 VSUBS 0.008903f
C266 B.n226 VSUBS 0.008903f
C267 B.n227 VSUBS 0.008903f
C268 B.n228 VSUBS 0.008903f
C269 B.n229 VSUBS 0.008903f
C270 B.n230 VSUBS 0.008903f
C271 B.n231 VSUBS 0.008903f
C272 B.n232 VSUBS 0.008903f
C273 B.n233 VSUBS 0.008903f
C274 B.n234 VSUBS 0.008903f
C275 B.n235 VSUBS 0.008903f
C276 B.n236 VSUBS 0.008903f
C277 B.n237 VSUBS 0.008903f
C278 B.n238 VSUBS 0.008903f
C279 B.n239 VSUBS 0.008903f
C280 B.n240 VSUBS 0.008903f
C281 B.n241 VSUBS 0.008903f
C282 B.n242 VSUBS 0.008903f
C283 B.n243 VSUBS 0.008903f
C284 B.n244 VSUBS 0.008903f
C285 B.n245 VSUBS 0.008903f
C286 B.n246 VSUBS 0.008903f
C287 B.n247 VSUBS 0.008903f
C288 B.n248 VSUBS 0.008903f
C289 B.n249 VSUBS 0.008903f
C290 B.n250 VSUBS 0.008903f
C291 B.n251 VSUBS 0.021505f
C292 B.n252 VSUBS 0.021505f
C293 B.n253 VSUBS 0.022747f
C294 B.n254 VSUBS 0.008903f
C295 B.n255 VSUBS 0.008903f
C296 B.n256 VSUBS 0.008903f
C297 B.n257 VSUBS 0.008903f
C298 B.n258 VSUBS 0.008903f
C299 B.n259 VSUBS 0.008903f
C300 B.n260 VSUBS 0.008903f
C301 B.n261 VSUBS 0.008903f
C302 B.n262 VSUBS 0.008903f
C303 B.n263 VSUBS 0.008903f
C304 B.n264 VSUBS 0.008903f
C305 B.n265 VSUBS 0.008903f
C306 B.n266 VSUBS 0.008903f
C307 B.n267 VSUBS 0.008903f
C308 B.n268 VSUBS 0.008903f
C309 B.n269 VSUBS 0.008903f
C310 B.n270 VSUBS 0.008903f
C311 B.n271 VSUBS 0.008903f
C312 B.n272 VSUBS 0.008903f
C313 B.n273 VSUBS 0.008903f
C314 B.n274 VSUBS 0.008903f
C315 B.n275 VSUBS 0.008903f
C316 B.n276 VSUBS 0.008903f
C317 B.n277 VSUBS 0.008903f
C318 B.n278 VSUBS 0.008903f
C319 B.n279 VSUBS 0.008903f
C320 B.n280 VSUBS 0.008903f
C321 B.n281 VSUBS 0.008903f
C322 B.n282 VSUBS 0.008903f
C323 B.n283 VSUBS 0.008903f
C324 B.n284 VSUBS 0.008903f
C325 B.n285 VSUBS 0.008903f
C326 B.n286 VSUBS 0.008903f
C327 B.n287 VSUBS 0.008903f
C328 B.n288 VSUBS 0.008903f
C329 B.n289 VSUBS 0.008903f
C330 B.n290 VSUBS 0.008903f
C331 B.n291 VSUBS 0.008903f
C332 B.n292 VSUBS 0.008903f
C333 B.n293 VSUBS 0.008903f
C334 B.n294 VSUBS 0.008903f
C335 B.n295 VSUBS 0.008903f
C336 B.n296 VSUBS 0.008903f
C337 B.n297 VSUBS 0.008903f
C338 B.n298 VSUBS 0.006153f
C339 B.n299 VSUBS 0.020627f
C340 B.n300 VSUBS 0.007201f
C341 B.n301 VSUBS 0.008903f
C342 B.n302 VSUBS 0.008903f
C343 B.n303 VSUBS 0.008903f
C344 B.n304 VSUBS 0.008903f
C345 B.n305 VSUBS 0.008903f
C346 B.n306 VSUBS 0.008903f
C347 B.n307 VSUBS 0.008903f
C348 B.n308 VSUBS 0.008903f
C349 B.n309 VSUBS 0.008903f
C350 B.n310 VSUBS 0.008903f
C351 B.n311 VSUBS 0.008903f
C352 B.n312 VSUBS 0.007201f
C353 B.n313 VSUBS 0.008903f
C354 B.n314 VSUBS 0.008903f
C355 B.n315 VSUBS 0.006153f
C356 B.n316 VSUBS 0.008903f
C357 B.n317 VSUBS 0.008903f
C358 B.n318 VSUBS 0.008903f
C359 B.n319 VSUBS 0.008903f
C360 B.n320 VSUBS 0.008903f
C361 B.n321 VSUBS 0.008903f
C362 B.n322 VSUBS 0.008903f
C363 B.n323 VSUBS 0.008903f
C364 B.n324 VSUBS 0.008903f
C365 B.n325 VSUBS 0.008903f
C366 B.n326 VSUBS 0.008903f
C367 B.n327 VSUBS 0.008903f
C368 B.n328 VSUBS 0.008903f
C369 B.n329 VSUBS 0.008903f
C370 B.n330 VSUBS 0.008903f
C371 B.n331 VSUBS 0.008903f
C372 B.n332 VSUBS 0.008903f
C373 B.n333 VSUBS 0.008903f
C374 B.n334 VSUBS 0.008903f
C375 B.n335 VSUBS 0.008903f
C376 B.n336 VSUBS 0.008903f
C377 B.n337 VSUBS 0.008903f
C378 B.n338 VSUBS 0.008903f
C379 B.n339 VSUBS 0.008903f
C380 B.n340 VSUBS 0.008903f
C381 B.n341 VSUBS 0.008903f
C382 B.n342 VSUBS 0.008903f
C383 B.n343 VSUBS 0.008903f
C384 B.n344 VSUBS 0.008903f
C385 B.n345 VSUBS 0.008903f
C386 B.n346 VSUBS 0.008903f
C387 B.n347 VSUBS 0.008903f
C388 B.n348 VSUBS 0.008903f
C389 B.n349 VSUBS 0.008903f
C390 B.n350 VSUBS 0.008903f
C391 B.n351 VSUBS 0.008903f
C392 B.n352 VSUBS 0.008903f
C393 B.n353 VSUBS 0.008903f
C394 B.n354 VSUBS 0.008903f
C395 B.n355 VSUBS 0.008903f
C396 B.n356 VSUBS 0.008903f
C397 B.n357 VSUBS 0.008903f
C398 B.n358 VSUBS 0.008903f
C399 B.n359 VSUBS 0.021786f
C400 B.n360 VSUBS 0.022747f
C401 B.n361 VSUBS 0.021505f
C402 B.n362 VSUBS 0.008903f
C403 B.n363 VSUBS 0.008903f
C404 B.n364 VSUBS 0.008903f
C405 B.n365 VSUBS 0.008903f
C406 B.n366 VSUBS 0.008903f
C407 B.n367 VSUBS 0.008903f
C408 B.n368 VSUBS 0.008903f
C409 B.n369 VSUBS 0.008903f
C410 B.n370 VSUBS 0.008903f
C411 B.n371 VSUBS 0.008903f
C412 B.n372 VSUBS 0.008903f
C413 B.n373 VSUBS 0.008903f
C414 B.n374 VSUBS 0.008903f
C415 B.n375 VSUBS 0.008903f
C416 B.n376 VSUBS 0.008903f
C417 B.n377 VSUBS 0.008903f
C418 B.n378 VSUBS 0.008903f
C419 B.n379 VSUBS 0.008903f
C420 B.n380 VSUBS 0.008903f
C421 B.n381 VSUBS 0.008903f
C422 B.n382 VSUBS 0.008903f
C423 B.n383 VSUBS 0.008903f
C424 B.n384 VSUBS 0.008903f
C425 B.n385 VSUBS 0.008903f
C426 B.n386 VSUBS 0.008903f
C427 B.n387 VSUBS 0.008903f
C428 B.n388 VSUBS 0.008903f
C429 B.n389 VSUBS 0.008903f
C430 B.n390 VSUBS 0.008903f
C431 B.n391 VSUBS 0.008903f
C432 B.n392 VSUBS 0.008903f
C433 B.n393 VSUBS 0.008903f
C434 B.n394 VSUBS 0.008903f
C435 B.n395 VSUBS 0.008903f
C436 B.n396 VSUBS 0.008903f
C437 B.n397 VSUBS 0.008903f
C438 B.n398 VSUBS 0.008903f
C439 B.n399 VSUBS 0.008903f
C440 B.n400 VSUBS 0.008903f
C441 B.n401 VSUBS 0.008903f
C442 B.n402 VSUBS 0.008903f
C443 B.n403 VSUBS 0.008903f
C444 B.n404 VSUBS 0.008903f
C445 B.n405 VSUBS 0.008903f
C446 B.n406 VSUBS 0.008903f
C447 B.n407 VSUBS 0.008903f
C448 B.n408 VSUBS 0.008903f
C449 B.n409 VSUBS 0.008903f
C450 B.n410 VSUBS 0.008903f
C451 B.n411 VSUBS 0.008903f
C452 B.n412 VSUBS 0.008903f
C453 B.n413 VSUBS 0.008903f
C454 B.n414 VSUBS 0.008903f
C455 B.n415 VSUBS 0.008903f
C456 B.n416 VSUBS 0.008903f
C457 B.n417 VSUBS 0.008903f
C458 B.n418 VSUBS 0.008903f
C459 B.n419 VSUBS 0.008903f
C460 B.n420 VSUBS 0.008903f
C461 B.n421 VSUBS 0.008903f
C462 B.n422 VSUBS 0.008903f
C463 B.n423 VSUBS 0.008903f
C464 B.n424 VSUBS 0.008903f
C465 B.n425 VSUBS 0.008903f
C466 B.n426 VSUBS 0.008903f
C467 B.n427 VSUBS 0.008903f
C468 B.n428 VSUBS 0.008903f
C469 B.n429 VSUBS 0.008903f
C470 B.n430 VSUBS 0.008903f
C471 B.n431 VSUBS 0.008903f
C472 B.n432 VSUBS 0.008903f
C473 B.n433 VSUBS 0.008903f
C474 B.n434 VSUBS 0.008903f
C475 B.n435 VSUBS 0.008903f
C476 B.n436 VSUBS 0.008903f
C477 B.n437 VSUBS 0.008903f
C478 B.n438 VSUBS 0.008903f
C479 B.n439 VSUBS 0.008903f
C480 B.n440 VSUBS 0.008903f
C481 B.n441 VSUBS 0.008903f
C482 B.n442 VSUBS 0.008903f
C483 B.n443 VSUBS 0.008903f
C484 B.n444 VSUBS 0.008903f
C485 B.n445 VSUBS 0.008903f
C486 B.n446 VSUBS 0.008903f
C487 B.n447 VSUBS 0.008903f
C488 B.n448 VSUBS 0.008903f
C489 B.n449 VSUBS 0.008903f
C490 B.n450 VSUBS 0.008903f
C491 B.n451 VSUBS 0.008903f
C492 B.n452 VSUBS 0.008903f
C493 B.n453 VSUBS 0.008903f
C494 B.n454 VSUBS 0.008903f
C495 B.n455 VSUBS 0.008903f
C496 B.n456 VSUBS 0.008903f
C497 B.n457 VSUBS 0.008903f
C498 B.n458 VSUBS 0.008903f
C499 B.n459 VSUBS 0.008903f
C500 B.n460 VSUBS 0.008903f
C501 B.n461 VSUBS 0.008903f
C502 B.n462 VSUBS 0.008903f
C503 B.n463 VSUBS 0.008903f
C504 B.n464 VSUBS 0.008903f
C505 B.n465 VSUBS 0.008903f
C506 B.n466 VSUBS 0.008903f
C507 B.n467 VSUBS 0.008903f
C508 B.n468 VSUBS 0.008903f
C509 B.n469 VSUBS 0.008903f
C510 B.n470 VSUBS 0.008903f
C511 B.n471 VSUBS 0.008903f
C512 B.n472 VSUBS 0.008903f
C513 B.n473 VSUBS 0.008903f
C514 B.n474 VSUBS 0.008903f
C515 B.n475 VSUBS 0.008903f
C516 B.n476 VSUBS 0.008903f
C517 B.n477 VSUBS 0.008903f
C518 B.n478 VSUBS 0.008903f
C519 B.n479 VSUBS 0.008903f
C520 B.n480 VSUBS 0.008903f
C521 B.n481 VSUBS 0.008903f
C522 B.n482 VSUBS 0.008903f
C523 B.n483 VSUBS 0.008903f
C524 B.n484 VSUBS 0.008903f
C525 B.n485 VSUBS 0.008903f
C526 B.n486 VSUBS 0.008903f
C527 B.n487 VSUBS 0.008903f
C528 B.n488 VSUBS 0.008903f
C529 B.n489 VSUBS 0.008903f
C530 B.n490 VSUBS 0.008903f
C531 B.n491 VSUBS 0.008903f
C532 B.n492 VSUBS 0.008903f
C533 B.n493 VSUBS 0.008903f
C534 B.n494 VSUBS 0.008903f
C535 B.n495 VSUBS 0.008903f
C536 B.n496 VSUBS 0.008903f
C537 B.n497 VSUBS 0.008903f
C538 B.n498 VSUBS 0.008903f
C539 B.n499 VSUBS 0.008903f
C540 B.n500 VSUBS 0.008903f
C541 B.n501 VSUBS 0.008903f
C542 B.n502 VSUBS 0.008903f
C543 B.n503 VSUBS 0.008903f
C544 B.n504 VSUBS 0.008903f
C545 B.n505 VSUBS 0.008903f
C546 B.n506 VSUBS 0.008903f
C547 B.n507 VSUBS 0.008903f
C548 B.n508 VSUBS 0.008903f
C549 B.n509 VSUBS 0.021505f
C550 B.n510 VSUBS 0.021505f
C551 B.n511 VSUBS 0.022747f
C552 B.n512 VSUBS 0.008903f
C553 B.n513 VSUBS 0.008903f
C554 B.n514 VSUBS 0.008903f
C555 B.n515 VSUBS 0.008903f
C556 B.n516 VSUBS 0.008903f
C557 B.n517 VSUBS 0.008903f
C558 B.n518 VSUBS 0.008903f
C559 B.n519 VSUBS 0.008903f
C560 B.n520 VSUBS 0.008903f
C561 B.n521 VSUBS 0.008903f
C562 B.n522 VSUBS 0.008903f
C563 B.n523 VSUBS 0.008903f
C564 B.n524 VSUBS 0.008903f
C565 B.n525 VSUBS 0.008903f
C566 B.n526 VSUBS 0.008903f
C567 B.n527 VSUBS 0.008903f
C568 B.n528 VSUBS 0.008903f
C569 B.n529 VSUBS 0.008903f
C570 B.n530 VSUBS 0.008903f
C571 B.n531 VSUBS 0.008903f
C572 B.n532 VSUBS 0.008903f
C573 B.n533 VSUBS 0.008903f
C574 B.n534 VSUBS 0.008903f
C575 B.n535 VSUBS 0.008903f
C576 B.n536 VSUBS 0.008903f
C577 B.n537 VSUBS 0.008903f
C578 B.n538 VSUBS 0.008903f
C579 B.n539 VSUBS 0.008903f
C580 B.n540 VSUBS 0.008903f
C581 B.n541 VSUBS 0.008903f
C582 B.n542 VSUBS 0.008903f
C583 B.n543 VSUBS 0.008903f
C584 B.n544 VSUBS 0.008903f
C585 B.n545 VSUBS 0.008903f
C586 B.n546 VSUBS 0.008903f
C587 B.n547 VSUBS 0.008903f
C588 B.n548 VSUBS 0.008903f
C589 B.n549 VSUBS 0.008903f
C590 B.n550 VSUBS 0.008903f
C591 B.n551 VSUBS 0.008903f
C592 B.n552 VSUBS 0.008903f
C593 B.n553 VSUBS 0.008903f
C594 B.n554 VSUBS 0.008903f
C595 B.n555 VSUBS 0.008903f
C596 B.n556 VSUBS 0.006153f
C597 B.n557 VSUBS 0.020627f
C598 B.n558 VSUBS 0.007201f
C599 B.n559 VSUBS 0.008903f
C600 B.n560 VSUBS 0.008903f
C601 B.n561 VSUBS 0.008903f
C602 B.n562 VSUBS 0.008903f
C603 B.n563 VSUBS 0.008903f
C604 B.n564 VSUBS 0.008903f
C605 B.n565 VSUBS 0.008903f
C606 B.n566 VSUBS 0.008903f
C607 B.n567 VSUBS 0.008903f
C608 B.n568 VSUBS 0.008903f
C609 B.n569 VSUBS 0.008903f
C610 B.n570 VSUBS 0.007201f
C611 B.n571 VSUBS 0.008903f
C612 B.n572 VSUBS 0.008903f
C613 B.n573 VSUBS 0.006153f
C614 B.n574 VSUBS 0.008903f
C615 B.n575 VSUBS 0.008903f
C616 B.n576 VSUBS 0.008903f
C617 B.n577 VSUBS 0.008903f
C618 B.n578 VSUBS 0.008903f
C619 B.n579 VSUBS 0.008903f
C620 B.n580 VSUBS 0.008903f
C621 B.n581 VSUBS 0.008903f
C622 B.n582 VSUBS 0.008903f
C623 B.n583 VSUBS 0.008903f
C624 B.n584 VSUBS 0.008903f
C625 B.n585 VSUBS 0.008903f
C626 B.n586 VSUBS 0.008903f
C627 B.n587 VSUBS 0.008903f
C628 B.n588 VSUBS 0.008903f
C629 B.n589 VSUBS 0.008903f
C630 B.n590 VSUBS 0.008903f
C631 B.n591 VSUBS 0.008903f
C632 B.n592 VSUBS 0.008903f
C633 B.n593 VSUBS 0.008903f
C634 B.n594 VSUBS 0.008903f
C635 B.n595 VSUBS 0.008903f
C636 B.n596 VSUBS 0.008903f
C637 B.n597 VSUBS 0.008903f
C638 B.n598 VSUBS 0.008903f
C639 B.n599 VSUBS 0.008903f
C640 B.n600 VSUBS 0.008903f
C641 B.n601 VSUBS 0.008903f
C642 B.n602 VSUBS 0.008903f
C643 B.n603 VSUBS 0.008903f
C644 B.n604 VSUBS 0.008903f
C645 B.n605 VSUBS 0.008903f
C646 B.n606 VSUBS 0.008903f
C647 B.n607 VSUBS 0.008903f
C648 B.n608 VSUBS 0.008903f
C649 B.n609 VSUBS 0.008903f
C650 B.n610 VSUBS 0.008903f
C651 B.n611 VSUBS 0.008903f
C652 B.n612 VSUBS 0.008903f
C653 B.n613 VSUBS 0.008903f
C654 B.n614 VSUBS 0.008903f
C655 B.n615 VSUBS 0.008903f
C656 B.n616 VSUBS 0.008903f
C657 B.n617 VSUBS 0.022747f
C658 B.n618 VSUBS 0.022747f
C659 B.n619 VSUBS 0.021505f
C660 B.n620 VSUBS 0.008903f
C661 B.n621 VSUBS 0.008903f
C662 B.n622 VSUBS 0.008903f
C663 B.n623 VSUBS 0.008903f
C664 B.n624 VSUBS 0.008903f
C665 B.n625 VSUBS 0.008903f
C666 B.n626 VSUBS 0.008903f
C667 B.n627 VSUBS 0.008903f
C668 B.n628 VSUBS 0.008903f
C669 B.n629 VSUBS 0.008903f
C670 B.n630 VSUBS 0.008903f
C671 B.n631 VSUBS 0.008903f
C672 B.n632 VSUBS 0.008903f
C673 B.n633 VSUBS 0.008903f
C674 B.n634 VSUBS 0.008903f
C675 B.n635 VSUBS 0.008903f
C676 B.n636 VSUBS 0.008903f
C677 B.n637 VSUBS 0.008903f
C678 B.n638 VSUBS 0.008903f
C679 B.n639 VSUBS 0.008903f
C680 B.n640 VSUBS 0.008903f
C681 B.n641 VSUBS 0.008903f
C682 B.n642 VSUBS 0.008903f
C683 B.n643 VSUBS 0.008903f
C684 B.n644 VSUBS 0.008903f
C685 B.n645 VSUBS 0.008903f
C686 B.n646 VSUBS 0.008903f
C687 B.n647 VSUBS 0.008903f
C688 B.n648 VSUBS 0.008903f
C689 B.n649 VSUBS 0.008903f
C690 B.n650 VSUBS 0.008903f
C691 B.n651 VSUBS 0.008903f
C692 B.n652 VSUBS 0.008903f
C693 B.n653 VSUBS 0.008903f
C694 B.n654 VSUBS 0.008903f
C695 B.n655 VSUBS 0.008903f
C696 B.n656 VSUBS 0.008903f
C697 B.n657 VSUBS 0.008903f
C698 B.n658 VSUBS 0.008903f
C699 B.n659 VSUBS 0.008903f
C700 B.n660 VSUBS 0.008903f
C701 B.n661 VSUBS 0.008903f
C702 B.n662 VSUBS 0.008903f
C703 B.n663 VSUBS 0.008903f
C704 B.n664 VSUBS 0.008903f
C705 B.n665 VSUBS 0.008903f
C706 B.n666 VSUBS 0.008903f
C707 B.n667 VSUBS 0.008903f
C708 B.n668 VSUBS 0.008903f
C709 B.n669 VSUBS 0.008903f
C710 B.n670 VSUBS 0.008903f
C711 B.n671 VSUBS 0.008903f
C712 B.n672 VSUBS 0.008903f
C713 B.n673 VSUBS 0.008903f
C714 B.n674 VSUBS 0.008903f
C715 B.n675 VSUBS 0.008903f
C716 B.n676 VSUBS 0.008903f
C717 B.n677 VSUBS 0.008903f
C718 B.n678 VSUBS 0.008903f
C719 B.n679 VSUBS 0.008903f
C720 B.n680 VSUBS 0.008903f
C721 B.n681 VSUBS 0.008903f
C722 B.n682 VSUBS 0.008903f
C723 B.n683 VSUBS 0.008903f
C724 B.n684 VSUBS 0.008903f
C725 B.n685 VSUBS 0.008903f
C726 B.n686 VSUBS 0.008903f
C727 B.n687 VSUBS 0.008903f
C728 B.n688 VSUBS 0.008903f
C729 B.n689 VSUBS 0.008903f
C730 B.n690 VSUBS 0.008903f
C731 B.n691 VSUBS 0.011618f
C732 B.n692 VSUBS 0.012376f
C733 B.n693 VSUBS 0.02461f
C734 VDD2.t0 VSUBS 1.89466f
C735 VDD2.t2 VSUBS 0.194513f
C736 VDD2.t3 VSUBS 0.194513f
C737 VDD2.n0 VSUBS 1.42957f
C738 VDD2.n1 VSUBS 4.00516f
C739 VDD2.t5 VSUBS 1.87471f
C740 VDD2.n2 VSUBS 3.42992f
C741 VDD2.t1 VSUBS 0.194513f
C742 VDD2.t4 VSUBS 0.194513f
C743 VDD2.n3 VSUBS 1.42953f
C744 VN.t2 VSUBS 2.2087f
C745 VN.n0 VSUBS 0.912515f
C746 VN.n1 VSUBS 0.03078f
C747 VN.n2 VSUBS 0.025041f
C748 VN.n3 VSUBS 0.03078f
C749 VN.t3 VSUBS 2.2087f
C750 VN.n4 VSUBS 0.896746f
C751 VN.t5 VSUBS 2.55787f
C752 VN.n5 VSUBS 0.85298f
C753 VN.n6 VSUBS 0.358569f
C754 VN.n7 VSUBS 0.043205f
C755 VN.n8 VSUBS 0.057366f
C756 VN.n9 VSUBS 0.06171f
C757 VN.n10 VSUBS 0.03078f
C758 VN.n11 VSUBS 0.03078f
C759 VN.n12 VSUBS 0.03078f
C760 VN.n13 VSUBS 0.060482f
C761 VN.n14 VSUBS 0.057366f
C762 VN.n15 VSUBS 0.045471f
C763 VN.n16 VSUBS 0.049678f
C764 VN.n17 VSUBS 0.073926f
C765 VN.t0 VSUBS 2.2087f
C766 VN.n18 VSUBS 0.912515f
C767 VN.n19 VSUBS 0.03078f
C768 VN.n20 VSUBS 0.025041f
C769 VN.n21 VSUBS 0.03078f
C770 VN.t4 VSUBS 2.2087f
C771 VN.n22 VSUBS 0.896746f
C772 VN.t1 VSUBS 2.55787f
C773 VN.n23 VSUBS 0.85298f
C774 VN.n24 VSUBS 0.358569f
C775 VN.n25 VSUBS 0.043205f
C776 VN.n26 VSUBS 0.057366f
C777 VN.n27 VSUBS 0.06171f
C778 VN.n28 VSUBS 0.03078f
C779 VN.n29 VSUBS 0.03078f
C780 VN.n30 VSUBS 0.03078f
C781 VN.n31 VSUBS 0.060482f
C782 VN.n32 VSUBS 0.057366f
C783 VN.n33 VSUBS 0.045471f
C784 VN.n34 VSUBS 0.049678f
C785 VN.n35 VSUBS 1.67938f
C786 VTAIL.t3 VSUBS 0.207391f
C787 VTAIL.t1 VSUBS 0.207391f
C788 VTAIL.n0 VSUBS 1.38519f
C789 VTAIL.n1 VSUBS 0.912246f
C790 VTAIL.t7 VSUBS 1.85532f
C791 VTAIL.n2 VSUBS 1.23472f
C792 VTAIL.t9 VSUBS 0.207391f
C793 VTAIL.t8 VSUBS 0.207391f
C794 VTAIL.n3 VSUBS 1.38519f
C795 VTAIL.n4 VSUBS 2.71527f
C796 VTAIL.t4 VSUBS 0.207391f
C797 VTAIL.t2 VSUBS 0.207391f
C798 VTAIL.n5 VSUBS 1.38519f
C799 VTAIL.n6 VSUBS 2.71526f
C800 VTAIL.t0 VSUBS 1.85533f
C801 VTAIL.n7 VSUBS 1.23471f
C802 VTAIL.t6 VSUBS 0.207391f
C803 VTAIL.t11 VSUBS 0.207391f
C804 VTAIL.n8 VSUBS 1.38519f
C805 VTAIL.n9 VSUBS 1.13923f
C806 VTAIL.t10 VSUBS 1.85532f
C807 VTAIL.n10 VSUBS 2.50019f
C808 VTAIL.t5 VSUBS 1.85532f
C809 VTAIL.n11 VSUBS 2.41663f
C810 VDD1.t1 VSUBS 1.67121f
C811 VDD1.t5 VSUBS 1.67009f
C812 VDD1.t0 VSUBS 0.171458f
C813 VDD1.t4 VSUBS 0.171458f
C814 VDD1.n0 VSUBS 1.26013f
C815 VDD1.n1 VSUBS 3.67318f
C816 VDD1.t2 VSUBS 0.171458f
C817 VDD1.t3 VSUBS 0.171458f
C818 VDD1.n2 VSUBS 1.25369f
C819 VDD1.n3 VSUBS 3.02686f
C820 VP.t4 VSUBS 2.47451f
C821 VP.n0 VSUBS 1.02233f
C822 VP.n1 VSUBS 0.034484f
C823 VP.n2 VSUBS 0.028055f
C824 VP.n3 VSUBS 0.034484f
C825 VP.t3 VSUBS 2.47451f
C826 VP.n4 VSUBS 0.891034f
C827 VP.n5 VSUBS 0.034484f
C828 VP.n6 VSUBS 0.028055f
C829 VP.n7 VSUBS 0.034484f
C830 VP.t2 VSUBS 2.47451f
C831 VP.n8 VSUBS 1.02233f
C832 VP.t1 VSUBS 2.47451f
C833 VP.n9 VSUBS 1.02233f
C834 VP.n10 VSUBS 0.034484f
C835 VP.n11 VSUBS 0.028055f
C836 VP.n12 VSUBS 0.034484f
C837 VP.t0 VSUBS 2.47451f
C838 VP.n13 VSUBS 1.00467f
C839 VP.t5 VSUBS 2.8657f
C840 VP.n14 VSUBS 0.955634f
C841 VP.n15 VSUBS 0.401722f
C842 VP.n16 VSUBS 0.048405f
C843 VP.n17 VSUBS 0.06427f
C844 VP.n18 VSUBS 0.069136f
C845 VP.n19 VSUBS 0.034484f
C846 VP.n20 VSUBS 0.034484f
C847 VP.n21 VSUBS 0.034484f
C848 VP.n22 VSUBS 0.067761f
C849 VP.n23 VSUBS 0.06427f
C850 VP.n24 VSUBS 0.050943f
C851 VP.n25 VSUBS 0.055657f
C852 VP.n26 VSUBS 1.8672f
C853 VP.n27 VSUBS 1.89284f
C854 VP.n28 VSUBS 0.055657f
C855 VP.n29 VSUBS 0.050943f
C856 VP.n30 VSUBS 0.06427f
C857 VP.n31 VSUBS 0.067761f
C858 VP.n32 VSUBS 0.034484f
C859 VP.n33 VSUBS 0.034484f
C860 VP.n34 VSUBS 0.034484f
C861 VP.n35 VSUBS 0.069136f
C862 VP.n36 VSUBS 0.06427f
C863 VP.n37 VSUBS 0.048405f
C864 VP.n38 VSUBS 0.034484f
C865 VP.n39 VSUBS 0.034484f
C866 VP.n40 VSUBS 0.048405f
C867 VP.n41 VSUBS 0.06427f
C868 VP.n42 VSUBS 0.069136f
C869 VP.n43 VSUBS 0.034484f
C870 VP.n44 VSUBS 0.034484f
C871 VP.n45 VSUBS 0.034484f
C872 VP.n46 VSUBS 0.067761f
C873 VP.n47 VSUBS 0.06427f
C874 VP.n48 VSUBS 0.050943f
C875 VP.n49 VSUBS 0.055657f
C876 VP.n50 VSUBS 0.082822f
.ends

