* NGSPICE file created from diff_pair_sample_0787.ext - technology: sky130A

.subckt diff_pair_sample_0787 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=3.14
X1 VDD1.t7 VP.t0 VTAIL.t12 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X2 VDD2.t7 VN.t0 VTAIL.t1 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X3 VTAIL.t0 VN.t1 VDD2.t6 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X4 VTAIL.t2 VN.t2 VDD2.t5 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X5 VDD1.t6 VP.t1 VTAIL.t10 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X6 VTAIL.t14 VP.t2 VDD1.t5 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X7 VDD2.t4 VN.t3 VTAIL.t6 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=3.14
X8 VDD2.t3 VN.t4 VTAIL.t15 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=3.14
X9 VTAIL.t13 VP.t3 VDD1.t4 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=3.14
X10 VTAIL.t7 VP.t4 VDD1.t3 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=3.14
X11 B.t8 B.t6 B.t7 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=3.14
X12 VDD1.t2 VP.t5 VTAIL.t8 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=3.14
X13 VTAIL.t3 VN.t5 VDD2.t2 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=3.14
X14 B.t5 B.t3 B.t4 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=3.14
X15 VTAIL.t11 VP.t6 VDD1.t1 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X16 VTAIL.t5 VN.t6 VDD2.t1 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=2.16975 ps=13.48 w=13.15 l=3.14
X17 B.t2 B.t0 B.t1 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=5.1285 pd=27.08 as=0 ps=0 w=13.15 l=3.14
X18 VDD2.t0 VN.t7 VTAIL.t4 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=2.16975 ps=13.48 w=13.15 l=3.14
X19 VDD1.t0 VP.t7 VTAIL.t9 w_n4440_n3598# sky130_fd_pr__pfet_01v8 ad=2.16975 pd=13.48 as=5.1285 ps=27.08 w=13.15 l=3.14
R0 B.n647 B.n646 585
R1 B.n648 B.n85 585
R2 B.n650 B.n649 585
R3 B.n651 B.n84 585
R4 B.n653 B.n652 585
R5 B.n654 B.n83 585
R6 B.n656 B.n655 585
R7 B.n657 B.n82 585
R8 B.n659 B.n658 585
R9 B.n660 B.n81 585
R10 B.n662 B.n661 585
R11 B.n663 B.n80 585
R12 B.n665 B.n664 585
R13 B.n666 B.n79 585
R14 B.n668 B.n667 585
R15 B.n669 B.n78 585
R16 B.n671 B.n670 585
R17 B.n672 B.n77 585
R18 B.n674 B.n673 585
R19 B.n675 B.n76 585
R20 B.n677 B.n676 585
R21 B.n678 B.n75 585
R22 B.n680 B.n679 585
R23 B.n681 B.n74 585
R24 B.n683 B.n682 585
R25 B.n684 B.n73 585
R26 B.n686 B.n685 585
R27 B.n687 B.n72 585
R28 B.n689 B.n688 585
R29 B.n690 B.n71 585
R30 B.n692 B.n691 585
R31 B.n693 B.n70 585
R32 B.n695 B.n694 585
R33 B.n696 B.n69 585
R34 B.n698 B.n697 585
R35 B.n699 B.n68 585
R36 B.n701 B.n700 585
R37 B.n702 B.n67 585
R38 B.n704 B.n703 585
R39 B.n705 B.n66 585
R40 B.n707 B.n706 585
R41 B.n708 B.n65 585
R42 B.n710 B.n709 585
R43 B.n711 B.n64 585
R44 B.n713 B.n712 585
R45 B.n715 B.n61 585
R46 B.n717 B.n716 585
R47 B.n718 B.n60 585
R48 B.n720 B.n719 585
R49 B.n721 B.n59 585
R50 B.n723 B.n722 585
R51 B.n724 B.n58 585
R52 B.n726 B.n725 585
R53 B.n727 B.n57 585
R54 B.n729 B.n728 585
R55 B.n731 B.n730 585
R56 B.n732 B.n53 585
R57 B.n734 B.n733 585
R58 B.n735 B.n52 585
R59 B.n737 B.n736 585
R60 B.n738 B.n51 585
R61 B.n740 B.n739 585
R62 B.n741 B.n50 585
R63 B.n743 B.n742 585
R64 B.n744 B.n49 585
R65 B.n746 B.n745 585
R66 B.n747 B.n48 585
R67 B.n749 B.n748 585
R68 B.n750 B.n47 585
R69 B.n752 B.n751 585
R70 B.n753 B.n46 585
R71 B.n755 B.n754 585
R72 B.n756 B.n45 585
R73 B.n758 B.n757 585
R74 B.n759 B.n44 585
R75 B.n761 B.n760 585
R76 B.n762 B.n43 585
R77 B.n764 B.n763 585
R78 B.n765 B.n42 585
R79 B.n767 B.n766 585
R80 B.n768 B.n41 585
R81 B.n770 B.n769 585
R82 B.n771 B.n40 585
R83 B.n773 B.n772 585
R84 B.n774 B.n39 585
R85 B.n776 B.n775 585
R86 B.n777 B.n38 585
R87 B.n779 B.n778 585
R88 B.n780 B.n37 585
R89 B.n782 B.n781 585
R90 B.n783 B.n36 585
R91 B.n785 B.n784 585
R92 B.n786 B.n35 585
R93 B.n788 B.n787 585
R94 B.n789 B.n34 585
R95 B.n791 B.n790 585
R96 B.n792 B.n33 585
R97 B.n794 B.n793 585
R98 B.n795 B.n32 585
R99 B.n797 B.n796 585
R100 B.n645 B.n86 585
R101 B.n644 B.n643 585
R102 B.n642 B.n87 585
R103 B.n641 B.n640 585
R104 B.n639 B.n88 585
R105 B.n638 B.n637 585
R106 B.n636 B.n89 585
R107 B.n635 B.n634 585
R108 B.n633 B.n90 585
R109 B.n632 B.n631 585
R110 B.n630 B.n91 585
R111 B.n629 B.n628 585
R112 B.n627 B.n92 585
R113 B.n626 B.n625 585
R114 B.n624 B.n93 585
R115 B.n623 B.n622 585
R116 B.n621 B.n94 585
R117 B.n620 B.n619 585
R118 B.n618 B.n95 585
R119 B.n617 B.n616 585
R120 B.n615 B.n96 585
R121 B.n614 B.n613 585
R122 B.n612 B.n97 585
R123 B.n611 B.n610 585
R124 B.n609 B.n98 585
R125 B.n608 B.n607 585
R126 B.n606 B.n99 585
R127 B.n605 B.n604 585
R128 B.n603 B.n100 585
R129 B.n602 B.n601 585
R130 B.n600 B.n101 585
R131 B.n599 B.n598 585
R132 B.n597 B.n102 585
R133 B.n596 B.n595 585
R134 B.n594 B.n103 585
R135 B.n593 B.n592 585
R136 B.n591 B.n104 585
R137 B.n590 B.n589 585
R138 B.n588 B.n105 585
R139 B.n587 B.n586 585
R140 B.n585 B.n106 585
R141 B.n584 B.n583 585
R142 B.n582 B.n107 585
R143 B.n581 B.n580 585
R144 B.n579 B.n108 585
R145 B.n578 B.n577 585
R146 B.n576 B.n109 585
R147 B.n575 B.n574 585
R148 B.n573 B.n110 585
R149 B.n572 B.n571 585
R150 B.n570 B.n111 585
R151 B.n569 B.n568 585
R152 B.n567 B.n112 585
R153 B.n566 B.n565 585
R154 B.n564 B.n113 585
R155 B.n563 B.n562 585
R156 B.n561 B.n114 585
R157 B.n560 B.n559 585
R158 B.n558 B.n115 585
R159 B.n557 B.n556 585
R160 B.n555 B.n116 585
R161 B.n554 B.n553 585
R162 B.n552 B.n117 585
R163 B.n551 B.n550 585
R164 B.n549 B.n118 585
R165 B.n548 B.n547 585
R166 B.n546 B.n119 585
R167 B.n545 B.n544 585
R168 B.n543 B.n120 585
R169 B.n542 B.n541 585
R170 B.n540 B.n121 585
R171 B.n539 B.n538 585
R172 B.n537 B.n122 585
R173 B.n536 B.n535 585
R174 B.n534 B.n123 585
R175 B.n533 B.n532 585
R176 B.n531 B.n124 585
R177 B.n530 B.n529 585
R178 B.n528 B.n125 585
R179 B.n527 B.n526 585
R180 B.n525 B.n126 585
R181 B.n524 B.n523 585
R182 B.n522 B.n127 585
R183 B.n521 B.n520 585
R184 B.n519 B.n128 585
R185 B.n518 B.n517 585
R186 B.n516 B.n129 585
R187 B.n515 B.n514 585
R188 B.n513 B.n130 585
R189 B.n512 B.n511 585
R190 B.n510 B.n131 585
R191 B.n509 B.n508 585
R192 B.n507 B.n132 585
R193 B.n506 B.n505 585
R194 B.n504 B.n133 585
R195 B.n503 B.n502 585
R196 B.n501 B.n134 585
R197 B.n500 B.n499 585
R198 B.n498 B.n135 585
R199 B.n497 B.n496 585
R200 B.n495 B.n136 585
R201 B.n494 B.n493 585
R202 B.n492 B.n137 585
R203 B.n491 B.n490 585
R204 B.n489 B.n138 585
R205 B.n488 B.n487 585
R206 B.n486 B.n139 585
R207 B.n485 B.n484 585
R208 B.n483 B.n140 585
R209 B.n482 B.n481 585
R210 B.n480 B.n141 585
R211 B.n479 B.n478 585
R212 B.n477 B.n142 585
R213 B.n476 B.n475 585
R214 B.n474 B.n143 585
R215 B.n473 B.n472 585
R216 B.n471 B.n144 585
R217 B.n470 B.n469 585
R218 B.n468 B.n145 585
R219 B.n317 B.n316 585
R220 B.n318 B.n199 585
R221 B.n320 B.n319 585
R222 B.n321 B.n198 585
R223 B.n323 B.n322 585
R224 B.n324 B.n197 585
R225 B.n326 B.n325 585
R226 B.n327 B.n196 585
R227 B.n329 B.n328 585
R228 B.n330 B.n195 585
R229 B.n332 B.n331 585
R230 B.n333 B.n194 585
R231 B.n335 B.n334 585
R232 B.n336 B.n193 585
R233 B.n338 B.n337 585
R234 B.n339 B.n192 585
R235 B.n341 B.n340 585
R236 B.n342 B.n191 585
R237 B.n344 B.n343 585
R238 B.n345 B.n190 585
R239 B.n347 B.n346 585
R240 B.n348 B.n189 585
R241 B.n350 B.n349 585
R242 B.n351 B.n188 585
R243 B.n353 B.n352 585
R244 B.n354 B.n187 585
R245 B.n356 B.n355 585
R246 B.n357 B.n186 585
R247 B.n359 B.n358 585
R248 B.n360 B.n185 585
R249 B.n362 B.n361 585
R250 B.n363 B.n184 585
R251 B.n365 B.n364 585
R252 B.n366 B.n183 585
R253 B.n368 B.n367 585
R254 B.n369 B.n182 585
R255 B.n371 B.n370 585
R256 B.n372 B.n181 585
R257 B.n374 B.n373 585
R258 B.n375 B.n180 585
R259 B.n377 B.n376 585
R260 B.n378 B.n179 585
R261 B.n380 B.n379 585
R262 B.n381 B.n178 585
R263 B.n383 B.n382 585
R264 B.n385 B.n175 585
R265 B.n387 B.n386 585
R266 B.n388 B.n174 585
R267 B.n390 B.n389 585
R268 B.n391 B.n173 585
R269 B.n393 B.n392 585
R270 B.n394 B.n172 585
R271 B.n396 B.n395 585
R272 B.n397 B.n171 585
R273 B.n399 B.n398 585
R274 B.n401 B.n400 585
R275 B.n402 B.n167 585
R276 B.n404 B.n403 585
R277 B.n405 B.n166 585
R278 B.n407 B.n406 585
R279 B.n408 B.n165 585
R280 B.n410 B.n409 585
R281 B.n411 B.n164 585
R282 B.n413 B.n412 585
R283 B.n414 B.n163 585
R284 B.n416 B.n415 585
R285 B.n417 B.n162 585
R286 B.n419 B.n418 585
R287 B.n420 B.n161 585
R288 B.n422 B.n421 585
R289 B.n423 B.n160 585
R290 B.n425 B.n424 585
R291 B.n426 B.n159 585
R292 B.n428 B.n427 585
R293 B.n429 B.n158 585
R294 B.n431 B.n430 585
R295 B.n432 B.n157 585
R296 B.n434 B.n433 585
R297 B.n435 B.n156 585
R298 B.n437 B.n436 585
R299 B.n438 B.n155 585
R300 B.n440 B.n439 585
R301 B.n441 B.n154 585
R302 B.n443 B.n442 585
R303 B.n444 B.n153 585
R304 B.n446 B.n445 585
R305 B.n447 B.n152 585
R306 B.n449 B.n448 585
R307 B.n450 B.n151 585
R308 B.n452 B.n451 585
R309 B.n453 B.n150 585
R310 B.n455 B.n454 585
R311 B.n456 B.n149 585
R312 B.n458 B.n457 585
R313 B.n459 B.n148 585
R314 B.n461 B.n460 585
R315 B.n462 B.n147 585
R316 B.n464 B.n463 585
R317 B.n465 B.n146 585
R318 B.n467 B.n466 585
R319 B.n315 B.n200 585
R320 B.n314 B.n313 585
R321 B.n312 B.n201 585
R322 B.n311 B.n310 585
R323 B.n309 B.n202 585
R324 B.n308 B.n307 585
R325 B.n306 B.n203 585
R326 B.n305 B.n304 585
R327 B.n303 B.n204 585
R328 B.n302 B.n301 585
R329 B.n300 B.n205 585
R330 B.n299 B.n298 585
R331 B.n297 B.n206 585
R332 B.n296 B.n295 585
R333 B.n294 B.n207 585
R334 B.n293 B.n292 585
R335 B.n291 B.n208 585
R336 B.n290 B.n289 585
R337 B.n288 B.n209 585
R338 B.n287 B.n286 585
R339 B.n285 B.n210 585
R340 B.n284 B.n283 585
R341 B.n282 B.n211 585
R342 B.n281 B.n280 585
R343 B.n279 B.n212 585
R344 B.n278 B.n277 585
R345 B.n276 B.n213 585
R346 B.n275 B.n274 585
R347 B.n273 B.n214 585
R348 B.n272 B.n271 585
R349 B.n270 B.n215 585
R350 B.n269 B.n268 585
R351 B.n267 B.n216 585
R352 B.n266 B.n265 585
R353 B.n264 B.n217 585
R354 B.n263 B.n262 585
R355 B.n261 B.n218 585
R356 B.n260 B.n259 585
R357 B.n258 B.n219 585
R358 B.n257 B.n256 585
R359 B.n255 B.n220 585
R360 B.n254 B.n253 585
R361 B.n252 B.n221 585
R362 B.n251 B.n250 585
R363 B.n249 B.n222 585
R364 B.n248 B.n247 585
R365 B.n246 B.n223 585
R366 B.n245 B.n244 585
R367 B.n243 B.n224 585
R368 B.n242 B.n241 585
R369 B.n240 B.n225 585
R370 B.n239 B.n238 585
R371 B.n237 B.n226 585
R372 B.n236 B.n235 585
R373 B.n234 B.n227 585
R374 B.n233 B.n232 585
R375 B.n231 B.n228 585
R376 B.n230 B.n229 585
R377 B.n2 B.n0 585
R378 B.n885 B.n1 585
R379 B.n884 B.n883 585
R380 B.n882 B.n3 585
R381 B.n881 B.n880 585
R382 B.n879 B.n4 585
R383 B.n878 B.n877 585
R384 B.n876 B.n5 585
R385 B.n875 B.n874 585
R386 B.n873 B.n6 585
R387 B.n872 B.n871 585
R388 B.n870 B.n7 585
R389 B.n869 B.n868 585
R390 B.n867 B.n8 585
R391 B.n866 B.n865 585
R392 B.n864 B.n9 585
R393 B.n863 B.n862 585
R394 B.n861 B.n10 585
R395 B.n860 B.n859 585
R396 B.n858 B.n11 585
R397 B.n857 B.n856 585
R398 B.n855 B.n12 585
R399 B.n854 B.n853 585
R400 B.n852 B.n13 585
R401 B.n851 B.n850 585
R402 B.n849 B.n14 585
R403 B.n848 B.n847 585
R404 B.n846 B.n15 585
R405 B.n845 B.n844 585
R406 B.n843 B.n16 585
R407 B.n842 B.n841 585
R408 B.n840 B.n17 585
R409 B.n839 B.n838 585
R410 B.n837 B.n18 585
R411 B.n836 B.n835 585
R412 B.n834 B.n19 585
R413 B.n833 B.n832 585
R414 B.n831 B.n20 585
R415 B.n830 B.n829 585
R416 B.n828 B.n21 585
R417 B.n827 B.n826 585
R418 B.n825 B.n22 585
R419 B.n824 B.n823 585
R420 B.n822 B.n23 585
R421 B.n821 B.n820 585
R422 B.n819 B.n24 585
R423 B.n818 B.n817 585
R424 B.n816 B.n25 585
R425 B.n815 B.n814 585
R426 B.n813 B.n26 585
R427 B.n812 B.n811 585
R428 B.n810 B.n27 585
R429 B.n809 B.n808 585
R430 B.n807 B.n28 585
R431 B.n806 B.n805 585
R432 B.n804 B.n29 585
R433 B.n803 B.n802 585
R434 B.n801 B.n30 585
R435 B.n800 B.n799 585
R436 B.n798 B.n31 585
R437 B.n887 B.n886 585
R438 B.n316 B.n315 487.695
R439 B.n796 B.n31 487.695
R440 B.n466 B.n145 487.695
R441 B.n646 B.n645 487.695
R442 B.n168 B.t0 309.666
R443 B.n176 B.t9 309.666
R444 B.n54 B.t3 309.666
R445 B.n62 B.t6 309.666
R446 B.n168 B.t2 178.624
R447 B.n62 B.t7 178.624
R448 B.n176 B.t11 178.607
R449 B.n54 B.t4 178.607
R450 B.n315 B.n314 163.367
R451 B.n314 B.n201 163.367
R452 B.n310 B.n201 163.367
R453 B.n310 B.n309 163.367
R454 B.n309 B.n308 163.367
R455 B.n308 B.n203 163.367
R456 B.n304 B.n203 163.367
R457 B.n304 B.n303 163.367
R458 B.n303 B.n302 163.367
R459 B.n302 B.n205 163.367
R460 B.n298 B.n205 163.367
R461 B.n298 B.n297 163.367
R462 B.n297 B.n296 163.367
R463 B.n296 B.n207 163.367
R464 B.n292 B.n207 163.367
R465 B.n292 B.n291 163.367
R466 B.n291 B.n290 163.367
R467 B.n290 B.n209 163.367
R468 B.n286 B.n209 163.367
R469 B.n286 B.n285 163.367
R470 B.n285 B.n284 163.367
R471 B.n284 B.n211 163.367
R472 B.n280 B.n211 163.367
R473 B.n280 B.n279 163.367
R474 B.n279 B.n278 163.367
R475 B.n278 B.n213 163.367
R476 B.n274 B.n213 163.367
R477 B.n274 B.n273 163.367
R478 B.n273 B.n272 163.367
R479 B.n272 B.n215 163.367
R480 B.n268 B.n215 163.367
R481 B.n268 B.n267 163.367
R482 B.n267 B.n266 163.367
R483 B.n266 B.n217 163.367
R484 B.n262 B.n217 163.367
R485 B.n262 B.n261 163.367
R486 B.n261 B.n260 163.367
R487 B.n260 B.n219 163.367
R488 B.n256 B.n219 163.367
R489 B.n256 B.n255 163.367
R490 B.n255 B.n254 163.367
R491 B.n254 B.n221 163.367
R492 B.n250 B.n221 163.367
R493 B.n250 B.n249 163.367
R494 B.n249 B.n248 163.367
R495 B.n248 B.n223 163.367
R496 B.n244 B.n223 163.367
R497 B.n244 B.n243 163.367
R498 B.n243 B.n242 163.367
R499 B.n242 B.n225 163.367
R500 B.n238 B.n225 163.367
R501 B.n238 B.n237 163.367
R502 B.n237 B.n236 163.367
R503 B.n236 B.n227 163.367
R504 B.n232 B.n227 163.367
R505 B.n232 B.n231 163.367
R506 B.n231 B.n230 163.367
R507 B.n230 B.n2 163.367
R508 B.n886 B.n2 163.367
R509 B.n886 B.n885 163.367
R510 B.n885 B.n884 163.367
R511 B.n884 B.n3 163.367
R512 B.n880 B.n3 163.367
R513 B.n880 B.n879 163.367
R514 B.n879 B.n878 163.367
R515 B.n878 B.n5 163.367
R516 B.n874 B.n5 163.367
R517 B.n874 B.n873 163.367
R518 B.n873 B.n872 163.367
R519 B.n872 B.n7 163.367
R520 B.n868 B.n7 163.367
R521 B.n868 B.n867 163.367
R522 B.n867 B.n866 163.367
R523 B.n866 B.n9 163.367
R524 B.n862 B.n9 163.367
R525 B.n862 B.n861 163.367
R526 B.n861 B.n860 163.367
R527 B.n860 B.n11 163.367
R528 B.n856 B.n11 163.367
R529 B.n856 B.n855 163.367
R530 B.n855 B.n854 163.367
R531 B.n854 B.n13 163.367
R532 B.n850 B.n13 163.367
R533 B.n850 B.n849 163.367
R534 B.n849 B.n848 163.367
R535 B.n848 B.n15 163.367
R536 B.n844 B.n15 163.367
R537 B.n844 B.n843 163.367
R538 B.n843 B.n842 163.367
R539 B.n842 B.n17 163.367
R540 B.n838 B.n17 163.367
R541 B.n838 B.n837 163.367
R542 B.n837 B.n836 163.367
R543 B.n836 B.n19 163.367
R544 B.n832 B.n19 163.367
R545 B.n832 B.n831 163.367
R546 B.n831 B.n830 163.367
R547 B.n830 B.n21 163.367
R548 B.n826 B.n21 163.367
R549 B.n826 B.n825 163.367
R550 B.n825 B.n824 163.367
R551 B.n824 B.n23 163.367
R552 B.n820 B.n23 163.367
R553 B.n820 B.n819 163.367
R554 B.n819 B.n818 163.367
R555 B.n818 B.n25 163.367
R556 B.n814 B.n25 163.367
R557 B.n814 B.n813 163.367
R558 B.n813 B.n812 163.367
R559 B.n812 B.n27 163.367
R560 B.n808 B.n27 163.367
R561 B.n808 B.n807 163.367
R562 B.n807 B.n806 163.367
R563 B.n806 B.n29 163.367
R564 B.n802 B.n29 163.367
R565 B.n802 B.n801 163.367
R566 B.n801 B.n800 163.367
R567 B.n800 B.n31 163.367
R568 B.n316 B.n199 163.367
R569 B.n320 B.n199 163.367
R570 B.n321 B.n320 163.367
R571 B.n322 B.n321 163.367
R572 B.n322 B.n197 163.367
R573 B.n326 B.n197 163.367
R574 B.n327 B.n326 163.367
R575 B.n328 B.n327 163.367
R576 B.n328 B.n195 163.367
R577 B.n332 B.n195 163.367
R578 B.n333 B.n332 163.367
R579 B.n334 B.n333 163.367
R580 B.n334 B.n193 163.367
R581 B.n338 B.n193 163.367
R582 B.n339 B.n338 163.367
R583 B.n340 B.n339 163.367
R584 B.n340 B.n191 163.367
R585 B.n344 B.n191 163.367
R586 B.n345 B.n344 163.367
R587 B.n346 B.n345 163.367
R588 B.n346 B.n189 163.367
R589 B.n350 B.n189 163.367
R590 B.n351 B.n350 163.367
R591 B.n352 B.n351 163.367
R592 B.n352 B.n187 163.367
R593 B.n356 B.n187 163.367
R594 B.n357 B.n356 163.367
R595 B.n358 B.n357 163.367
R596 B.n358 B.n185 163.367
R597 B.n362 B.n185 163.367
R598 B.n363 B.n362 163.367
R599 B.n364 B.n363 163.367
R600 B.n364 B.n183 163.367
R601 B.n368 B.n183 163.367
R602 B.n369 B.n368 163.367
R603 B.n370 B.n369 163.367
R604 B.n370 B.n181 163.367
R605 B.n374 B.n181 163.367
R606 B.n375 B.n374 163.367
R607 B.n376 B.n375 163.367
R608 B.n376 B.n179 163.367
R609 B.n380 B.n179 163.367
R610 B.n381 B.n380 163.367
R611 B.n382 B.n381 163.367
R612 B.n382 B.n175 163.367
R613 B.n387 B.n175 163.367
R614 B.n388 B.n387 163.367
R615 B.n389 B.n388 163.367
R616 B.n389 B.n173 163.367
R617 B.n393 B.n173 163.367
R618 B.n394 B.n393 163.367
R619 B.n395 B.n394 163.367
R620 B.n395 B.n171 163.367
R621 B.n399 B.n171 163.367
R622 B.n400 B.n399 163.367
R623 B.n400 B.n167 163.367
R624 B.n404 B.n167 163.367
R625 B.n405 B.n404 163.367
R626 B.n406 B.n405 163.367
R627 B.n406 B.n165 163.367
R628 B.n410 B.n165 163.367
R629 B.n411 B.n410 163.367
R630 B.n412 B.n411 163.367
R631 B.n412 B.n163 163.367
R632 B.n416 B.n163 163.367
R633 B.n417 B.n416 163.367
R634 B.n418 B.n417 163.367
R635 B.n418 B.n161 163.367
R636 B.n422 B.n161 163.367
R637 B.n423 B.n422 163.367
R638 B.n424 B.n423 163.367
R639 B.n424 B.n159 163.367
R640 B.n428 B.n159 163.367
R641 B.n429 B.n428 163.367
R642 B.n430 B.n429 163.367
R643 B.n430 B.n157 163.367
R644 B.n434 B.n157 163.367
R645 B.n435 B.n434 163.367
R646 B.n436 B.n435 163.367
R647 B.n436 B.n155 163.367
R648 B.n440 B.n155 163.367
R649 B.n441 B.n440 163.367
R650 B.n442 B.n441 163.367
R651 B.n442 B.n153 163.367
R652 B.n446 B.n153 163.367
R653 B.n447 B.n446 163.367
R654 B.n448 B.n447 163.367
R655 B.n448 B.n151 163.367
R656 B.n452 B.n151 163.367
R657 B.n453 B.n452 163.367
R658 B.n454 B.n453 163.367
R659 B.n454 B.n149 163.367
R660 B.n458 B.n149 163.367
R661 B.n459 B.n458 163.367
R662 B.n460 B.n459 163.367
R663 B.n460 B.n147 163.367
R664 B.n464 B.n147 163.367
R665 B.n465 B.n464 163.367
R666 B.n466 B.n465 163.367
R667 B.n470 B.n145 163.367
R668 B.n471 B.n470 163.367
R669 B.n472 B.n471 163.367
R670 B.n472 B.n143 163.367
R671 B.n476 B.n143 163.367
R672 B.n477 B.n476 163.367
R673 B.n478 B.n477 163.367
R674 B.n478 B.n141 163.367
R675 B.n482 B.n141 163.367
R676 B.n483 B.n482 163.367
R677 B.n484 B.n483 163.367
R678 B.n484 B.n139 163.367
R679 B.n488 B.n139 163.367
R680 B.n489 B.n488 163.367
R681 B.n490 B.n489 163.367
R682 B.n490 B.n137 163.367
R683 B.n494 B.n137 163.367
R684 B.n495 B.n494 163.367
R685 B.n496 B.n495 163.367
R686 B.n496 B.n135 163.367
R687 B.n500 B.n135 163.367
R688 B.n501 B.n500 163.367
R689 B.n502 B.n501 163.367
R690 B.n502 B.n133 163.367
R691 B.n506 B.n133 163.367
R692 B.n507 B.n506 163.367
R693 B.n508 B.n507 163.367
R694 B.n508 B.n131 163.367
R695 B.n512 B.n131 163.367
R696 B.n513 B.n512 163.367
R697 B.n514 B.n513 163.367
R698 B.n514 B.n129 163.367
R699 B.n518 B.n129 163.367
R700 B.n519 B.n518 163.367
R701 B.n520 B.n519 163.367
R702 B.n520 B.n127 163.367
R703 B.n524 B.n127 163.367
R704 B.n525 B.n524 163.367
R705 B.n526 B.n525 163.367
R706 B.n526 B.n125 163.367
R707 B.n530 B.n125 163.367
R708 B.n531 B.n530 163.367
R709 B.n532 B.n531 163.367
R710 B.n532 B.n123 163.367
R711 B.n536 B.n123 163.367
R712 B.n537 B.n536 163.367
R713 B.n538 B.n537 163.367
R714 B.n538 B.n121 163.367
R715 B.n542 B.n121 163.367
R716 B.n543 B.n542 163.367
R717 B.n544 B.n543 163.367
R718 B.n544 B.n119 163.367
R719 B.n548 B.n119 163.367
R720 B.n549 B.n548 163.367
R721 B.n550 B.n549 163.367
R722 B.n550 B.n117 163.367
R723 B.n554 B.n117 163.367
R724 B.n555 B.n554 163.367
R725 B.n556 B.n555 163.367
R726 B.n556 B.n115 163.367
R727 B.n560 B.n115 163.367
R728 B.n561 B.n560 163.367
R729 B.n562 B.n561 163.367
R730 B.n562 B.n113 163.367
R731 B.n566 B.n113 163.367
R732 B.n567 B.n566 163.367
R733 B.n568 B.n567 163.367
R734 B.n568 B.n111 163.367
R735 B.n572 B.n111 163.367
R736 B.n573 B.n572 163.367
R737 B.n574 B.n573 163.367
R738 B.n574 B.n109 163.367
R739 B.n578 B.n109 163.367
R740 B.n579 B.n578 163.367
R741 B.n580 B.n579 163.367
R742 B.n580 B.n107 163.367
R743 B.n584 B.n107 163.367
R744 B.n585 B.n584 163.367
R745 B.n586 B.n585 163.367
R746 B.n586 B.n105 163.367
R747 B.n590 B.n105 163.367
R748 B.n591 B.n590 163.367
R749 B.n592 B.n591 163.367
R750 B.n592 B.n103 163.367
R751 B.n596 B.n103 163.367
R752 B.n597 B.n596 163.367
R753 B.n598 B.n597 163.367
R754 B.n598 B.n101 163.367
R755 B.n602 B.n101 163.367
R756 B.n603 B.n602 163.367
R757 B.n604 B.n603 163.367
R758 B.n604 B.n99 163.367
R759 B.n608 B.n99 163.367
R760 B.n609 B.n608 163.367
R761 B.n610 B.n609 163.367
R762 B.n610 B.n97 163.367
R763 B.n614 B.n97 163.367
R764 B.n615 B.n614 163.367
R765 B.n616 B.n615 163.367
R766 B.n616 B.n95 163.367
R767 B.n620 B.n95 163.367
R768 B.n621 B.n620 163.367
R769 B.n622 B.n621 163.367
R770 B.n622 B.n93 163.367
R771 B.n626 B.n93 163.367
R772 B.n627 B.n626 163.367
R773 B.n628 B.n627 163.367
R774 B.n628 B.n91 163.367
R775 B.n632 B.n91 163.367
R776 B.n633 B.n632 163.367
R777 B.n634 B.n633 163.367
R778 B.n634 B.n89 163.367
R779 B.n638 B.n89 163.367
R780 B.n639 B.n638 163.367
R781 B.n640 B.n639 163.367
R782 B.n640 B.n87 163.367
R783 B.n644 B.n87 163.367
R784 B.n645 B.n644 163.367
R785 B.n796 B.n795 163.367
R786 B.n795 B.n794 163.367
R787 B.n794 B.n33 163.367
R788 B.n790 B.n33 163.367
R789 B.n790 B.n789 163.367
R790 B.n789 B.n788 163.367
R791 B.n788 B.n35 163.367
R792 B.n784 B.n35 163.367
R793 B.n784 B.n783 163.367
R794 B.n783 B.n782 163.367
R795 B.n782 B.n37 163.367
R796 B.n778 B.n37 163.367
R797 B.n778 B.n777 163.367
R798 B.n777 B.n776 163.367
R799 B.n776 B.n39 163.367
R800 B.n772 B.n39 163.367
R801 B.n772 B.n771 163.367
R802 B.n771 B.n770 163.367
R803 B.n770 B.n41 163.367
R804 B.n766 B.n41 163.367
R805 B.n766 B.n765 163.367
R806 B.n765 B.n764 163.367
R807 B.n764 B.n43 163.367
R808 B.n760 B.n43 163.367
R809 B.n760 B.n759 163.367
R810 B.n759 B.n758 163.367
R811 B.n758 B.n45 163.367
R812 B.n754 B.n45 163.367
R813 B.n754 B.n753 163.367
R814 B.n753 B.n752 163.367
R815 B.n752 B.n47 163.367
R816 B.n748 B.n47 163.367
R817 B.n748 B.n747 163.367
R818 B.n747 B.n746 163.367
R819 B.n746 B.n49 163.367
R820 B.n742 B.n49 163.367
R821 B.n742 B.n741 163.367
R822 B.n741 B.n740 163.367
R823 B.n740 B.n51 163.367
R824 B.n736 B.n51 163.367
R825 B.n736 B.n735 163.367
R826 B.n735 B.n734 163.367
R827 B.n734 B.n53 163.367
R828 B.n730 B.n53 163.367
R829 B.n730 B.n729 163.367
R830 B.n729 B.n57 163.367
R831 B.n725 B.n57 163.367
R832 B.n725 B.n724 163.367
R833 B.n724 B.n723 163.367
R834 B.n723 B.n59 163.367
R835 B.n719 B.n59 163.367
R836 B.n719 B.n718 163.367
R837 B.n718 B.n717 163.367
R838 B.n717 B.n61 163.367
R839 B.n712 B.n61 163.367
R840 B.n712 B.n711 163.367
R841 B.n711 B.n710 163.367
R842 B.n710 B.n65 163.367
R843 B.n706 B.n65 163.367
R844 B.n706 B.n705 163.367
R845 B.n705 B.n704 163.367
R846 B.n704 B.n67 163.367
R847 B.n700 B.n67 163.367
R848 B.n700 B.n699 163.367
R849 B.n699 B.n698 163.367
R850 B.n698 B.n69 163.367
R851 B.n694 B.n69 163.367
R852 B.n694 B.n693 163.367
R853 B.n693 B.n692 163.367
R854 B.n692 B.n71 163.367
R855 B.n688 B.n71 163.367
R856 B.n688 B.n687 163.367
R857 B.n687 B.n686 163.367
R858 B.n686 B.n73 163.367
R859 B.n682 B.n73 163.367
R860 B.n682 B.n681 163.367
R861 B.n681 B.n680 163.367
R862 B.n680 B.n75 163.367
R863 B.n676 B.n75 163.367
R864 B.n676 B.n675 163.367
R865 B.n675 B.n674 163.367
R866 B.n674 B.n77 163.367
R867 B.n670 B.n77 163.367
R868 B.n670 B.n669 163.367
R869 B.n669 B.n668 163.367
R870 B.n668 B.n79 163.367
R871 B.n664 B.n79 163.367
R872 B.n664 B.n663 163.367
R873 B.n663 B.n662 163.367
R874 B.n662 B.n81 163.367
R875 B.n658 B.n81 163.367
R876 B.n658 B.n657 163.367
R877 B.n657 B.n656 163.367
R878 B.n656 B.n83 163.367
R879 B.n652 B.n83 163.367
R880 B.n652 B.n651 163.367
R881 B.n651 B.n650 163.367
R882 B.n650 B.n85 163.367
R883 B.n646 B.n85 163.367
R884 B.n169 B.t1 111.326
R885 B.n63 B.t8 111.326
R886 B.n177 B.t10 111.311
R887 B.n55 B.t5 111.311
R888 B.n169 B.n168 67.2975
R889 B.n177 B.n176 67.2975
R890 B.n55 B.n54 67.2975
R891 B.n63 B.n62 67.2975
R892 B.n170 B.n169 59.5399
R893 B.n384 B.n177 59.5399
R894 B.n56 B.n55 59.5399
R895 B.n714 B.n63 59.5399
R896 B.n798 B.n797 31.6883
R897 B.n647 B.n86 31.6883
R898 B.n468 B.n467 31.6883
R899 B.n317 B.n200 31.6883
R900 B B.n887 18.0485
R901 B.n797 B.n32 10.6151
R902 B.n793 B.n32 10.6151
R903 B.n793 B.n792 10.6151
R904 B.n792 B.n791 10.6151
R905 B.n791 B.n34 10.6151
R906 B.n787 B.n34 10.6151
R907 B.n787 B.n786 10.6151
R908 B.n786 B.n785 10.6151
R909 B.n785 B.n36 10.6151
R910 B.n781 B.n36 10.6151
R911 B.n781 B.n780 10.6151
R912 B.n780 B.n779 10.6151
R913 B.n779 B.n38 10.6151
R914 B.n775 B.n38 10.6151
R915 B.n775 B.n774 10.6151
R916 B.n774 B.n773 10.6151
R917 B.n773 B.n40 10.6151
R918 B.n769 B.n40 10.6151
R919 B.n769 B.n768 10.6151
R920 B.n768 B.n767 10.6151
R921 B.n767 B.n42 10.6151
R922 B.n763 B.n42 10.6151
R923 B.n763 B.n762 10.6151
R924 B.n762 B.n761 10.6151
R925 B.n761 B.n44 10.6151
R926 B.n757 B.n44 10.6151
R927 B.n757 B.n756 10.6151
R928 B.n756 B.n755 10.6151
R929 B.n755 B.n46 10.6151
R930 B.n751 B.n46 10.6151
R931 B.n751 B.n750 10.6151
R932 B.n750 B.n749 10.6151
R933 B.n749 B.n48 10.6151
R934 B.n745 B.n48 10.6151
R935 B.n745 B.n744 10.6151
R936 B.n744 B.n743 10.6151
R937 B.n743 B.n50 10.6151
R938 B.n739 B.n50 10.6151
R939 B.n739 B.n738 10.6151
R940 B.n738 B.n737 10.6151
R941 B.n737 B.n52 10.6151
R942 B.n733 B.n52 10.6151
R943 B.n733 B.n732 10.6151
R944 B.n732 B.n731 10.6151
R945 B.n728 B.n727 10.6151
R946 B.n727 B.n726 10.6151
R947 B.n726 B.n58 10.6151
R948 B.n722 B.n58 10.6151
R949 B.n722 B.n721 10.6151
R950 B.n721 B.n720 10.6151
R951 B.n720 B.n60 10.6151
R952 B.n716 B.n60 10.6151
R953 B.n716 B.n715 10.6151
R954 B.n713 B.n64 10.6151
R955 B.n709 B.n64 10.6151
R956 B.n709 B.n708 10.6151
R957 B.n708 B.n707 10.6151
R958 B.n707 B.n66 10.6151
R959 B.n703 B.n66 10.6151
R960 B.n703 B.n702 10.6151
R961 B.n702 B.n701 10.6151
R962 B.n701 B.n68 10.6151
R963 B.n697 B.n68 10.6151
R964 B.n697 B.n696 10.6151
R965 B.n696 B.n695 10.6151
R966 B.n695 B.n70 10.6151
R967 B.n691 B.n70 10.6151
R968 B.n691 B.n690 10.6151
R969 B.n690 B.n689 10.6151
R970 B.n689 B.n72 10.6151
R971 B.n685 B.n72 10.6151
R972 B.n685 B.n684 10.6151
R973 B.n684 B.n683 10.6151
R974 B.n683 B.n74 10.6151
R975 B.n679 B.n74 10.6151
R976 B.n679 B.n678 10.6151
R977 B.n678 B.n677 10.6151
R978 B.n677 B.n76 10.6151
R979 B.n673 B.n76 10.6151
R980 B.n673 B.n672 10.6151
R981 B.n672 B.n671 10.6151
R982 B.n671 B.n78 10.6151
R983 B.n667 B.n78 10.6151
R984 B.n667 B.n666 10.6151
R985 B.n666 B.n665 10.6151
R986 B.n665 B.n80 10.6151
R987 B.n661 B.n80 10.6151
R988 B.n661 B.n660 10.6151
R989 B.n660 B.n659 10.6151
R990 B.n659 B.n82 10.6151
R991 B.n655 B.n82 10.6151
R992 B.n655 B.n654 10.6151
R993 B.n654 B.n653 10.6151
R994 B.n653 B.n84 10.6151
R995 B.n649 B.n84 10.6151
R996 B.n649 B.n648 10.6151
R997 B.n648 B.n647 10.6151
R998 B.n469 B.n468 10.6151
R999 B.n469 B.n144 10.6151
R1000 B.n473 B.n144 10.6151
R1001 B.n474 B.n473 10.6151
R1002 B.n475 B.n474 10.6151
R1003 B.n475 B.n142 10.6151
R1004 B.n479 B.n142 10.6151
R1005 B.n480 B.n479 10.6151
R1006 B.n481 B.n480 10.6151
R1007 B.n481 B.n140 10.6151
R1008 B.n485 B.n140 10.6151
R1009 B.n486 B.n485 10.6151
R1010 B.n487 B.n486 10.6151
R1011 B.n487 B.n138 10.6151
R1012 B.n491 B.n138 10.6151
R1013 B.n492 B.n491 10.6151
R1014 B.n493 B.n492 10.6151
R1015 B.n493 B.n136 10.6151
R1016 B.n497 B.n136 10.6151
R1017 B.n498 B.n497 10.6151
R1018 B.n499 B.n498 10.6151
R1019 B.n499 B.n134 10.6151
R1020 B.n503 B.n134 10.6151
R1021 B.n504 B.n503 10.6151
R1022 B.n505 B.n504 10.6151
R1023 B.n505 B.n132 10.6151
R1024 B.n509 B.n132 10.6151
R1025 B.n510 B.n509 10.6151
R1026 B.n511 B.n510 10.6151
R1027 B.n511 B.n130 10.6151
R1028 B.n515 B.n130 10.6151
R1029 B.n516 B.n515 10.6151
R1030 B.n517 B.n516 10.6151
R1031 B.n517 B.n128 10.6151
R1032 B.n521 B.n128 10.6151
R1033 B.n522 B.n521 10.6151
R1034 B.n523 B.n522 10.6151
R1035 B.n523 B.n126 10.6151
R1036 B.n527 B.n126 10.6151
R1037 B.n528 B.n527 10.6151
R1038 B.n529 B.n528 10.6151
R1039 B.n529 B.n124 10.6151
R1040 B.n533 B.n124 10.6151
R1041 B.n534 B.n533 10.6151
R1042 B.n535 B.n534 10.6151
R1043 B.n535 B.n122 10.6151
R1044 B.n539 B.n122 10.6151
R1045 B.n540 B.n539 10.6151
R1046 B.n541 B.n540 10.6151
R1047 B.n541 B.n120 10.6151
R1048 B.n545 B.n120 10.6151
R1049 B.n546 B.n545 10.6151
R1050 B.n547 B.n546 10.6151
R1051 B.n547 B.n118 10.6151
R1052 B.n551 B.n118 10.6151
R1053 B.n552 B.n551 10.6151
R1054 B.n553 B.n552 10.6151
R1055 B.n553 B.n116 10.6151
R1056 B.n557 B.n116 10.6151
R1057 B.n558 B.n557 10.6151
R1058 B.n559 B.n558 10.6151
R1059 B.n559 B.n114 10.6151
R1060 B.n563 B.n114 10.6151
R1061 B.n564 B.n563 10.6151
R1062 B.n565 B.n564 10.6151
R1063 B.n565 B.n112 10.6151
R1064 B.n569 B.n112 10.6151
R1065 B.n570 B.n569 10.6151
R1066 B.n571 B.n570 10.6151
R1067 B.n571 B.n110 10.6151
R1068 B.n575 B.n110 10.6151
R1069 B.n576 B.n575 10.6151
R1070 B.n577 B.n576 10.6151
R1071 B.n577 B.n108 10.6151
R1072 B.n581 B.n108 10.6151
R1073 B.n582 B.n581 10.6151
R1074 B.n583 B.n582 10.6151
R1075 B.n583 B.n106 10.6151
R1076 B.n587 B.n106 10.6151
R1077 B.n588 B.n587 10.6151
R1078 B.n589 B.n588 10.6151
R1079 B.n589 B.n104 10.6151
R1080 B.n593 B.n104 10.6151
R1081 B.n594 B.n593 10.6151
R1082 B.n595 B.n594 10.6151
R1083 B.n595 B.n102 10.6151
R1084 B.n599 B.n102 10.6151
R1085 B.n600 B.n599 10.6151
R1086 B.n601 B.n600 10.6151
R1087 B.n601 B.n100 10.6151
R1088 B.n605 B.n100 10.6151
R1089 B.n606 B.n605 10.6151
R1090 B.n607 B.n606 10.6151
R1091 B.n607 B.n98 10.6151
R1092 B.n611 B.n98 10.6151
R1093 B.n612 B.n611 10.6151
R1094 B.n613 B.n612 10.6151
R1095 B.n613 B.n96 10.6151
R1096 B.n617 B.n96 10.6151
R1097 B.n618 B.n617 10.6151
R1098 B.n619 B.n618 10.6151
R1099 B.n619 B.n94 10.6151
R1100 B.n623 B.n94 10.6151
R1101 B.n624 B.n623 10.6151
R1102 B.n625 B.n624 10.6151
R1103 B.n625 B.n92 10.6151
R1104 B.n629 B.n92 10.6151
R1105 B.n630 B.n629 10.6151
R1106 B.n631 B.n630 10.6151
R1107 B.n631 B.n90 10.6151
R1108 B.n635 B.n90 10.6151
R1109 B.n636 B.n635 10.6151
R1110 B.n637 B.n636 10.6151
R1111 B.n637 B.n88 10.6151
R1112 B.n641 B.n88 10.6151
R1113 B.n642 B.n641 10.6151
R1114 B.n643 B.n642 10.6151
R1115 B.n643 B.n86 10.6151
R1116 B.n318 B.n317 10.6151
R1117 B.n319 B.n318 10.6151
R1118 B.n319 B.n198 10.6151
R1119 B.n323 B.n198 10.6151
R1120 B.n324 B.n323 10.6151
R1121 B.n325 B.n324 10.6151
R1122 B.n325 B.n196 10.6151
R1123 B.n329 B.n196 10.6151
R1124 B.n330 B.n329 10.6151
R1125 B.n331 B.n330 10.6151
R1126 B.n331 B.n194 10.6151
R1127 B.n335 B.n194 10.6151
R1128 B.n336 B.n335 10.6151
R1129 B.n337 B.n336 10.6151
R1130 B.n337 B.n192 10.6151
R1131 B.n341 B.n192 10.6151
R1132 B.n342 B.n341 10.6151
R1133 B.n343 B.n342 10.6151
R1134 B.n343 B.n190 10.6151
R1135 B.n347 B.n190 10.6151
R1136 B.n348 B.n347 10.6151
R1137 B.n349 B.n348 10.6151
R1138 B.n349 B.n188 10.6151
R1139 B.n353 B.n188 10.6151
R1140 B.n354 B.n353 10.6151
R1141 B.n355 B.n354 10.6151
R1142 B.n355 B.n186 10.6151
R1143 B.n359 B.n186 10.6151
R1144 B.n360 B.n359 10.6151
R1145 B.n361 B.n360 10.6151
R1146 B.n361 B.n184 10.6151
R1147 B.n365 B.n184 10.6151
R1148 B.n366 B.n365 10.6151
R1149 B.n367 B.n366 10.6151
R1150 B.n367 B.n182 10.6151
R1151 B.n371 B.n182 10.6151
R1152 B.n372 B.n371 10.6151
R1153 B.n373 B.n372 10.6151
R1154 B.n373 B.n180 10.6151
R1155 B.n377 B.n180 10.6151
R1156 B.n378 B.n377 10.6151
R1157 B.n379 B.n378 10.6151
R1158 B.n379 B.n178 10.6151
R1159 B.n383 B.n178 10.6151
R1160 B.n386 B.n385 10.6151
R1161 B.n386 B.n174 10.6151
R1162 B.n390 B.n174 10.6151
R1163 B.n391 B.n390 10.6151
R1164 B.n392 B.n391 10.6151
R1165 B.n392 B.n172 10.6151
R1166 B.n396 B.n172 10.6151
R1167 B.n397 B.n396 10.6151
R1168 B.n398 B.n397 10.6151
R1169 B.n402 B.n401 10.6151
R1170 B.n403 B.n402 10.6151
R1171 B.n403 B.n166 10.6151
R1172 B.n407 B.n166 10.6151
R1173 B.n408 B.n407 10.6151
R1174 B.n409 B.n408 10.6151
R1175 B.n409 B.n164 10.6151
R1176 B.n413 B.n164 10.6151
R1177 B.n414 B.n413 10.6151
R1178 B.n415 B.n414 10.6151
R1179 B.n415 B.n162 10.6151
R1180 B.n419 B.n162 10.6151
R1181 B.n420 B.n419 10.6151
R1182 B.n421 B.n420 10.6151
R1183 B.n421 B.n160 10.6151
R1184 B.n425 B.n160 10.6151
R1185 B.n426 B.n425 10.6151
R1186 B.n427 B.n426 10.6151
R1187 B.n427 B.n158 10.6151
R1188 B.n431 B.n158 10.6151
R1189 B.n432 B.n431 10.6151
R1190 B.n433 B.n432 10.6151
R1191 B.n433 B.n156 10.6151
R1192 B.n437 B.n156 10.6151
R1193 B.n438 B.n437 10.6151
R1194 B.n439 B.n438 10.6151
R1195 B.n439 B.n154 10.6151
R1196 B.n443 B.n154 10.6151
R1197 B.n444 B.n443 10.6151
R1198 B.n445 B.n444 10.6151
R1199 B.n445 B.n152 10.6151
R1200 B.n449 B.n152 10.6151
R1201 B.n450 B.n449 10.6151
R1202 B.n451 B.n450 10.6151
R1203 B.n451 B.n150 10.6151
R1204 B.n455 B.n150 10.6151
R1205 B.n456 B.n455 10.6151
R1206 B.n457 B.n456 10.6151
R1207 B.n457 B.n148 10.6151
R1208 B.n461 B.n148 10.6151
R1209 B.n462 B.n461 10.6151
R1210 B.n463 B.n462 10.6151
R1211 B.n463 B.n146 10.6151
R1212 B.n467 B.n146 10.6151
R1213 B.n313 B.n200 10.6151
R1214 B.n313 B.n312 10.6151
R1215 B.n312 B.n311 10.6151
R1216 B.n311 B.n202 10.6151
R1217 B.n307 B.n202 10.6151
R1218 B.n307 B.n306 10.6151
R1219 B.n306 B.n305 10.6151
R1220 B.n305 B.n204 10.6151
R1221 B.n301 B.n204 10.6151
R1222 B.n301 B.n300 10.6151
R1223 B.n300 B.n299 10.6151
R1224 B.n299 B.n206 10.6151
R1225 B.n295 B.n206 10.6151
R1226 B.n295 B.n294 10.6151
R1227 B.n294 B.n293 10.6151
R1228 B.n293 B.n208 10.6151
R1229 B.n289 B.n208 10.6151
R1230 B.n289 B.n288 10.6151
R1231 B.n288 B.n287 10.6151
R1232 B.n287 B.n210 10.6151
R1233 B.n283 B.n210 10.6151
R1234 B.n283 B.n282 10.6151
R1235 B.n282 B.n281 10.6151
R1236 B.n281 B.n212 10.6151
R1237 B.n277 B.n212 10.6151
R1238 B.n277 B.n276 10.6151
R1239 B.n276 B.n275 10.6151
R1240 B.n275 B.n214 10.6151
R1241 B.n271 B.n214 10.6151
R1242 B.n271 B.n270 10.6151
R1243 B.n270 B.n269 10.6151
R1244 B.n269 B.n216 10.6151
R1245 B.n265 B.n216 10.6151
R1246 B.n265 B.n264 10.6151
R1247 B.n264 B.n263 10.6151
R1248 B.n263 B.n218 10.6151
R1249 B.n259 B.n218 10.6151
R1250 B.n259 B.n258 10.6151
R1251 B.n258 B.n257 10.6151
R1252 B.n257 B.n220 10.6151
R1253 B.n253 B.n220 10.6151
R1254 B.n253 B.n252 10.6151
R1255 B.n252 B.n251 10.6151
R1256 B.n251 B.n222 10.6151
R1257 B.n247 B.n222 10.6151
R1258 B.n247 B.n246 10.6151
R1259 B.n246 B.n245 10.6151
R1260 B.n245 B.n224 10.6151
R1261 B.n241 B.n224 10.6151
R1262 B.n241 B.n240 10.6151
R1263 B.n240 B.n239 10.6151
R1264 B.n239 B.n226 10.6151
R1265 B.n235 B.n226 10.6151
R1266 B.n235 B.n234 10.6151
R1267 B.n234 B.n233 10.6151
R1268 B.n233 B.n228 10.6151
R1269 B.n229 B.n228 10.6151
R1270 B.n229 B.n0 10.6151
R1271 B.n883 B.n1 10.6151
R1272 B.n883 B.n882 10.6151
R1273 B.n882 B.n881 10.6151
R1274 B.n881 B.n4 10.6151
R1275 B.n877 B.n4 10.6151
R1276 B.n877 B.n876 10.6151
R1277 B.n876 B.n875 10.6151
R1278 B.n875 B.n6 10.6151
R1279 B.n871 B.n6 10.6151
R1280 B.n871 B.n870 10.6151
R1281 B.n870 B.n869 10.6151
R1282 B.n869 B.n8 10.6151
R1283 B.n865 B.n8 10.6151
R1284 B.n865 B.n864 10.6151
R1285 B.n864 B.n863 10.6151
R1286 B.n863 B.n10 10.6151
R1287 B.n859 B.n10 10.6151
R1288 B.n859 B.n858 10.6151
R1289 B.n858 B.n857 10.6151
R1290 B.n857 B.n12 10.6151
R1291 B.n853 B.n12 10.6151
R1292 B.n853 B.n852 10.6151
R1293 B.n852 B.n851 10.6151
R1294 B.n851 B.n14 10.6151
R1295 B.n847 B.n14 10.6151
R1296 B.n847 B.n846 10.6151
R1297 B.n846 B.n845 10.6151
R1298 B.n845 B.n16 10.6151
R1299 B.n841 B.n16 10.6151
R1300 B.n841 B.n840 10.6151
R1301 B.n840 B.n839 10.6151
R1302 B.n839 B.n18 10.6151
R1303 B.n835 B.n18 10.6151
R1304 B.n835 B.n834 10.6151
R1305 B.n834 B.n833 10.6151
R1306 B.n833 B.n20 10.6151
R1307 B.n829 B.n20 10.6151
R1308 B.n829 B.n828 10.6151
R1309 B.n828 B.n827 10.6151
R1310 B.n827 B.n22 10.6151
R1311 B.n823 B.n22 10.6151
R1312 B.n823 B.n822 10.6151
R1313 B.n822 B.n821 10.6151
R1314 B.n821 B.n24 10.6151
R1315 B.n817 B.n24 10.6151
R1316 B.n817 B.n816 10.6151
R1317 B.n816 B.n815 10.6151
R1318 B.n815 B.n26 10.6151
R1319 B.n811 B.n26 10.6151
R1320 B.n811 B.n810 10.6151
R1321 B.n810 B.n809 10.6151
R1322 B.n809 B.n28 10.6151
R1323 B.n805 B.n28 10.6151
R1324 B.n805 B.n804 10.6151
R1325 B.n804 B.n803 10.6151
R1326 B.n803 B.n30 10.6151
R1327 B.n799 B.n30 10.6151
R1328 B.n799 B.n798 10.6151
R1329 B.n731 B.n56 9.36635
R1330 B.n714 B.n713 9.36635
R1331 B.n384 B.n383 9.36635
R1332 B.n401 B.n170 9.36635
R1333 B.n887 B.n0 2.81026
R1334 B.n887 B.n1 2.81026
R1335 B.n728 B.n56 1.24928
R1336 B.n715 B.n714 1.24928
R1337 B.n385 B.n384 1.24928
R1338 B.n398 B.n170 1.24928
R1339 VP.n21 VP.n18 161.3
R1340 VP.n23 VP.n22 161.3
R1341 VP.n24 VP.n17 161.3
R1342 VP.n26 VP.n25 161.3
R1343 VP.n27 VP.n16 161.3
R1344 VP.n29 VP.n28 161.3
R1345 VP.n31 VP.n30 161.3
R1346 VP.n32 VP.n14 161.3
R1347 VP.n34 VP.n33 161.3
R1348 VP.n35 VP.n13 161.3
R1349 VP.n37 VP.n36 161.3
R1350 VP.n38 VP.n12 161.3
R1351 VP.n40 VP.n39 161.3
R1352 VP.n75 VP.n74 161.3
R1353 VP.n73 VP.n1 161.3
R1354 VP.n72 VP.n71 161.3
R1355 VP.n70 VP.n2 161.3
R1356 VP.n69 VP.n68 161.3
R1357 VP.n67 VP.n3 161.3
R1358 VP.n66 VP.n65 161.3
R1359 VP.n64 VP.n63 161.3
R1360 VP.n62 VP.n5 161.3
R1361 VP.n61 VP.n60 161.3
R1362 VP.n59 VP.n6 161.3
R1363 VP.n58 VP.n57 161.3
R1364 VP.n56 VP.n7 161.3
R1365 VP.n54 VP.n53 161.3
R1366 VP.n52 VP.n8 161.3
R1367 VP.n51 VP.n50 161.3
R1368 VP.n49 VP.n9 161.3
R1369 VP.n48 VP.n47 161.3
R1370 VP.n46 VP.n10 161.3
R1371 VP.n45 VP.n44 161.3
R1372 VP.n19 VP.t3 134.344
R1373 VP.n43 VP.t4 100.928
R1374 VP.n55 VP.t1 100.928
R1375 VP.n4 VP.t2 100.928
R1376 VP.n0 VP.t7 100.928
R1377 VP.n11 VP.t5 100.928
R1378 VP.n15 VP.t6 100.928
R1379 VP.n20 VP.t0 100.928
R1380 VP.n43 VP.n42 67.8024
R1381 VP.n76 VP.n0 67.8024
R1382 VP.n41 VP.n11 67.8024
R1383 VP.n49 VP.n48 56.5193
R1384 VP.n61 VP.n6 56.5193
R1385 VP.n72 VP.n2 56.5193
R1386 VP.n37 VP.n13 56.5193
R1387 VP.n26 VP.n17 56.5193
R1388 VP.n42 VP.n41 54.4842
R1389 VP.n20 VP.n19 50.2421
R1390 VP.n44 VP.n10 24.4675
R1391 VP.n48 VP.n10 24.4675
R1392 VP.n50 VP.n49 24.4675
R1393 VP.n50 VP.n8 24.4675
R1394 VP.n54 VP.n8 24.4675
R1395 VP.n57 VP.n56 24.4675
R1396 VP.n57 VP.n6 24.4675
R1397 VP.n62 VP.n61 24.4675
R1398 VP.n63 VP.n62 24.4675
R1399 VP.n67 VP.n66 24.4675
R1400 VP.n68 VP.n67 24.4675
R1401 VP.n68 VP.n2 24.4675
R1402 VP.n73 VP.n72 24.4675
R1403 VP.n74 VP.n73 24.4675
R1404 VP.n38 VP.n37 24.4675
R1405 VP.n39 VP.n38 24.4675
R1406 VP.n27 VP.n26 24.4675
R1407 VP.n28 VP.n27 24.4675
R1408 VP.n32 VP.n31 24.4675
R1409 VP.n33 VP.n32 24.4675
R1410 VP.n33 VP.n13 24.4675
R1411 VP.n22 VP.n21 24.4675
R1412 VP.n22 VP.n17 24.4675
R1413 VP.n56 VP.n55 23.7335
R1414 VP.n63 VP.n4 23.7335
R1415 VP.n28 VP.n15 23.7335
R1416 VP.n21 VP.n20 23.7335
R1417 VP.n44 VP.n43 22.2655
R1418 VP.n74 VP.n0 22.2655
R1419 VP.n39 VP.n11 22.2655
R1420 VP.n19 VP.n18 3.80563
R1421 VP.n55 VP.n54 0.73451
R1422 VP.n66 VP.n4 0.73451
R1423 VP.n31 VP.n15 0.73451
R1424 VP.n41 VP.n40 0.354971
R1425 VP.n45 VP.n42 0.354971
R1426 VP.n76 VP.n75 0.354971
R1427 VP VP.n76 0.26696
R1428 VP.n23 VP.n18 0.189894
R1429 VP.n24 VP.n23 0.189894
R1430 VP.n25 VP.n24 0.189894
R1431 VP.n25 VP.n16 0.189894
R1432 VP.n29 VP.n16 0.189894
R1433 VP.n30 VP.n29 0.189894
R1434 VP.n30 VP.n14 0.189894
R1435 VP.n34 VP.n14 0.189894
R1436 VP.n35 VP.n34 0.189894
R1437 VP.n36 VP.n35 0.189894
R1438 VP.n36 VP.n12 0.189894
R1439 VP.n40 VP.n12 0.189894
R1440 VP.n46 VP.n45 0.189894
R1441 VP.n47 VP.n46 0.189894
R1442 VP.n47 VP.n9 0.189894
R1443 VP.n51 VP.n9 0.189894
R1444 VP.n52 VP.n51 0.189894
R1445 VP.n53 VP.n52 0.189894
R1446 VP.n53 VP.n7 0.189894
R1447 VP.n58 VP.n7 0.189894
R1448 VP.n59 VP.n58 0.189894
R1449 VP.n60 VP.n59 0.189894
R1450 VP.n60 VP.n5 0.189894
R1451 VP.n64 VP.n5 0.189894
R1452 VP.n65 VP.n64 0.189894
R1453 VP.n65 VP.n3 0.189894
R1454 VP.n69 VP.n3 0.189894
R1455 VP.n70 VP.n69 0.189894
R1456 VP.n71 VP.n70 0.189894
R1457 VP.n71 VP.n1 0.189894
R1458 VP.n75 VP.n1 0.189894
R1459 VTAIL.n11 VTAIL.t13 57.4581
R1460 VTAIL.n10 VTAIL.t15 57.4581
R1461 VTAIL.n7 VTAIL.t5 57.4581
R1462 VTAIL.n15 VTAIL.t6 57.4578
R1463 VTAIL.n2 VTAIL.t3 57.4578
R1464 VTAIL.n3 VTAIL.t9 57.4578
R1465 VTAIL.n6 VTAIL.t7 57.4578
R1466 VTAIL.n14 VTAIL.t8 57.4578
R1467 VTAIL.n13 VTAIL.n12 54.9862
R1468 VTAIL.n9 VTAIL.n8 54.9862
R1469 VTAIL.n1 VTAIL.n0 54.9861
R1470 VTAIL.n5 VTAIL.n4 54.9861
R1471 VTAIL.n15 VTAIL.n14 26.6945
R1472 VTAIL.n7 VTAIL.n6 26.6945
R1473 VTAIL.n9 VTAIL.n7 2.99188
R1474 VTAIL.n10 VTAIL.n9 2.99188
R1475 VTAIL.n13 VTAIL.n11 2.99188
R1476 VTAIL.n14 VTAIL.n13 2.99188
R1477 VTAIL.n6 VTAIL.n5 2.99188
R1478 VTAIL.n5 VTAIL.n3 2.99188
R1479 VTAIL.n2 VTAIL.n1 2.99188
R1480 VTAIL VTAIL.n15 2.93369
R1481 VTAIL.n0 VTAIL.t4 2.47236
R1482 VTAIL.n0 VTAIL.t0 2.47236
R1483 VTAIL.n4 VTAIL.t10 2.47236
R1484 VTAIL.n4 VTAIL.t14 2.47236
R1485 VTAIL.n12 VTAIL.t12 2.47236
R1486 VTAIL.n12 VTAIL.t11 2.47236
R1487 VTAIL.n8 VTAIL.t1 2.47236
R1488 VTAIL.n8 VTAIL.t2 2.47236
R1489 VTAIL.n11 VTAIL.n10 0.470328
R1490 VTAIL.n3 VTAIL.n2 0.470328
R1491 VTAIL VTAIL.n1 0.0586897
R1492 VDD1 VDD1.n0 73.2189
R1493 VDD1.n3 VDD1.n2 73.1053
R1494 VDD1.n3 VDD1.n1 73.1053
R1495 VDD1.n5 VDD1.n4 71.6648
R1496 VDD1.n5 VDD1.n3 49.0957
R1497 VDD1.n4 VDD1.t1 2.47236
R1498 VDD1.n4 VDD1.t2 2.47236
R1499 VDD1.n0 VDD1.t4 2.47236
R1500 VDD1.n0 VDD1.t7 2.47236
R1501 VDD1.n2 VDD1.t5 2.47236
R1502 VDD1.n2 VDD1.t0 2.47236
R1503 VDD1.n1 VDD1.t3 2.47236
R1504 VDD1.n1 VDD1.t6 2.47236
R1505 VDD1 VDD1.n5 1.438
R1506 VN.n60 VN.n59 161.3
R1507 VN.n58 VN.n32 161.3
R1508 VN.n57 VN.n56 161.3
R1509 VN.n55 VN.n33 161.3
R1510 VN.n54 VN.n53 161.3
R1511 VN.n52 VN.n34 161.3
R1512 VN.n51 VN.n50 161.3
R1513 VN.n49 VN.n48 161.3
R1514 VN.n47 VN.n36 161.3
R1515 VN.n46 VN.n45 161.3
R1516 VN.n44 VN.n37 161.3
R1517 VN.n43 VN.n42 161.3
R1518 VN.n41 VN.n38 161.3
R1519 VN.n29 VN.n28 161.3
R1520 VN.n27 VN.n1 161.3
R1521 VN.n26 VN.n25 161.3
R1522 VN.n24 VN.n2 161.3
R1523 VN.n23 VN.n22 161.3
R1524 VN.n21 VN.n3 161.3
R1525 VN.n20 VN.n19 161.3
R1526 VN.n18 VN.n17 161.3
R1527 VN.n16 VN.n5 161.3
R1528 VN.n15 VN.n14 161.3
R1529 VN.n13 VN.n6 161.3
R1530 VN.n12 VN.n11 161.3
R1531 VN.n10 VN.n7 161.3
R1532 VN.n39 VN.t4 134.344
R1533 VN.n8 VN.t5 134.344
R1534 VN.n9 VN.t7 100.928
R1535 VN.n4 VN.t1 100.928
R1536 VN.n0 VN.t3 100.928
R1537 VN.n40 VN.t2 100.928
R1538 VN.n35 VN.t0 100.928
R1539 VN.n31 VN.t6 100.928
R1540 VN.n30 VN.n0 67.8024
R1541 VN.n61 VN.n31 67.8024
R1542 VN.n15 VN.n6 56.5193
R1543 VN.n26 VN.n2 56.5193
R1544 VN.n46 VN.n37 56.5193
R1545 VN.n57 VN.n33 56.5193
R1546 VN VN.n61 54.6495
R1547 VN.n40 VN.n39 50.2421
R1548 VN.n9 VN.n8 50.2421
R1549 VN.n11 VN.n10 24.4675
R1550 VN.n11 VN.n6 24.4675
R1551 VN.n16 VN.n15 24.4675
R1552 VN.n17 VN.n16 24.4675
R1553 VN.n21 VN.n20 24.4675
R1554 VN.n22 VN.n21 24.4675
R1555 VN.n22 VN.n2 24.4675
R1556 VN.n27 VN.n26 24.4675
R1557 VN.n28 VN.n27 24.4675
R1558 VN.n42 VN.n37 24.4675
R1559 VN.n42 VN.n41 24.4675
R1560 VN.n53 VN.n33 24.4675
R1561 VN.n53 VN.n52 24.4675
R1562 VN.n52 VN.n51 24.4675
R1563 VN.n48 VN.n47 24.4675
R1564 VN.n47 VN.n46 24.4675
R1565 VN.n59 VN.n58 24.4675
R1566 VN.n58 VN.n57 24.4675
R1567 VN.n10 VN.n9 23.7335
R1568 VN.n17 VN.n4 23.7335
R1569 VN.n41 VN.n40 23.7335
R1570 VN.n48 VN.n35 23.7335
R1571 VN.n28 VN.n0 22.2655
R1572 VN.n59 VN.n31 22.2655
R1573 VN.n39 VN.n38 3.80565
R1574 VN.n8 VN.n7 3.80565
R1575 VN.n20 VN.n4 0.73451
R1576 VN.n51 VN.n35 0.73451
R1577 VN.n61 VN.n60 0.354971
R1578 VN.n30 VN.n29 0.354971
R1579 VN VN.n30 0.26696
R1580 VN.n60 VN.n32 0.189894
R1581 VN.n56 VN.n32 0.189894
R1582 VN.n56 VN.n55 0.189894
R1583 VN.n55 VN.n54 0.189894
R1584 VN.n54 VN.n34 0.189894
R1585 VN.n50 VN.n34 0.189894
R1586 VN.n50 VN.n49 0.189894
R1587 VN.n49 VN.n36 0.189894
R1588 VN.n45 VN.n36 0.189894
R1589 VN.n45 VN.n44 0.189894
R1590 VN.n44 VN.n43 0.189894
R1591 VN.n43 VN.n38 0.189894
R1592 VN.n12 VN.n7 0.189894
R1593 VN.n13 VN.n12 0.189894
R1594 VN.n14 VN.n13 0.189894
R1595 VN.n14 VN.n5 0.189894
R1596 VN.n18 VN.n5 0.189894
R1597 VN.n19 VN.n18 0.189894
R1598 VN.n19 VN.n3 0.189894
R1599 VN.n23 VN.n3 0.189894
R1600 VN.n24 VN.n23 0.189894
R1601 VN.n25 VN.n24 0.189894
R1602 VN.n25 VN.n1 0.189894
R1603 VN.n29 VN.n1 0.189894
R1604 VDD2.n2 VDD2.n1 73.1053
R1605 VDD2.n2 VDD2.n0 73.1053
R1606 VDD2 VDD2.n5 73.1023
R1607 VDD2.n4 VDD2.n3 71.665
R1608 VDD2.n4 VDD2.n2 48.5127
R1609 VDD2.n5 VDD2.t5 2.47236
R1610 VDD2.n5 VDD2.t3 2.47236
R1611 VDD2.n3 VDD2.t1 2.47236
R1612 VDD2.n3 VDD2.t7 2.47236
R1613 VDD2.n1 VDD2.t6 2.47236
R1614 VDD2.n1 VDD2.t4 2.47236
R1615 VDD2.n0 VDD2.t2 2.47236
R1616 VDD2.n0 VDD2.t0 2.47236
R1617 VDD2 VDD2.n4 1.55438
C0 VDD1 VDD2 2.05959f
C1 VTAIL VDD2 8.65874f
C2 VDD1 VP 10.23f
C3 VTAIL VP 10.348599f
C4 w_n4440_n3598# VN 9.19862f
C5 w_n4440_n3598# B 11.264799f
C6 B VN 1.36438f
C7 VDD1 w_n4440_n3598# 2.16246f
C8 w_n4440_n3598# VTAIL 4.51422f
C9 VDD1 VN 0.152829f
C10 VTAIL VN 10.3345f
C11 VDD2 VP 0.577257f
C12 VDD1 B 1.84471f
C13 B VTAIL 5.60501f
C14 VDD1 VTAIL 8.6007f
C15 w_n4440_n3598# VDD2 2.29982f
C16 w_n4440_n3598# VP 9.77662f
C17 VDD2 VN 9.807281f
C18 VN VP 8.53445f
C19 B VDD2 1.95773f
C20 B VP 2.33618f
C21 VDD2 VSUBS 2.204078f
C22 VDD1 VSUBS 2.94465f
C23 VTAIL VSUBS 1.482269f
C24 VN VSUBS 7.49895f
C25 VP VSUBS 4.195594f
C26 B VSUBS 5.703357f
C27 w_n4440_n3598# VSUBS 0.196337p
C28 VDD2.t2 VSUBS 0.311077f
C29 VDD2.t0 VSUBS 0.311077f
C30 VDD2.n0 VSUBS 2.47904f
C31 VDD2.t6 VSUBS 0.311077f
C32 VDD2.t4 VSUBS 0.311077f
C33 VDD2.n1 VSUBS 2.47904f
C34 VDD2.n2 VSUBS 5.03816f
C35 VDD2.t1 VSUBS 0.311077f
C36 VDD2.t7 VSUBS 0.311077f
C37 VDD2.n3 VSUBS 2.45901f
C38 VDD2.n4 VSUBS 4.19222f
C39 VDD2.t5 VSUBS 0.311077f
C40 VDD2.t3 VSUBS 0.311077f
C41 VDD2.n5 VSUBS 2.47898f
C42 VN.t3 VSUBS 2.87726f
C43 VN.n0 VSUBS 1.1167f
C44 VN.n1 VSUBS 0.025511f
C45 VN.n2 VSUBS 0.035109f
C46 VN.n3 VSUBS 0.025511f
C47 VN.t1 VSUBS 2.87726f
C48 VN.n4 VSUBS 1.0075f
C49 VN.n5 VSUBS 0.025511f
C50 VN.n6 VSUBS 0.037242f
C51 VN.n7 VSUBS 0.290507f
C52 VN.t7 VSUBS 2.87726f
C53 VN.t5 VSUBS 3.17407f
C54 VN.n8 VSUBS 1.04826f
C55 VN.n9 VSUBS 1.10314f
C56 VN.n10 VSUBS 0.046841f
C57 VN.n11 VSUBS 0.047547f
C58 VN.n12 VSUBS 0.025511f
C59 VN.n13 VSUBS 0.025511f
C60 VN.n14 VSUBS 0.025511f
C61 VN.n15 VSUBS 0.037242f
C62 VN.n16 VSUBS 0.047547f
C63 VN.n17 VSUBS 0.046841f
C64 VN.n18 VSUBS 0.025511f
C65 VN.n19 VSUBS 0.025511f
C66 VN.n20 VSUBS 0.024776f
C67 VN.n21 VSUBS 0.047547f
C68 VN.n22 VSUBS 0.047547f
C69 VN.n23 VSUBS 0.025511f
C70 VN.n24 VSUBS 0.025511f
C71 VN.n25 VSUBS 0.025511f
C72 VN.n26 VSUBS 0.039375f
C73 VN.n27 VSUBS 0.047547f
C74 VN.n28 VSUBS 0.045433f
C75 VN.n29 VSUBS 0.041175f
C76 VN.n30 VSUBS 0.051374f
C77 VN.t6 VSUBS 2.87726f
C78 VN.n31 VSUBS 1.1167f
C79 VN.n32 VSUBS 0.025511f
C80 VN.n33 VSUBS 0.035109f
C81 VN.n34 VSUBS 0.025511f
C82 VN.t0 VSUBS 2.87726f
C83 VN.n35 VSUBS 1.0075f
C84 VN.n36 VSUBS 0.025511f
C85 VN.n37 VSUBS 0.037242f
C86 VN.n38 VSUBS 0.290507f
C87 VN.t2 VSUBS 2.87726f
C88 VN.t4 VSUBS 3.17407f
C89 VN.n39 VSUBS 1.04826f
C90 VN.n40 VSUBS 1.10314f
C91 VN.n41 VSUBS 0.046841f
C92 VN.n42 VSUBS 0.047547f
C93 VN.n43 VSUBS 0.025511f
C94 VN.n44 VSUBS 0.025511f
C95 VN.n45 VSUBS 0.025511f
C96 VN.n46 VSUBS 0.037242f
C97 VN.n47 VSUBS 0.047547f
C98 VN.n48 VSUBS 0.046841f
C99 VN.n49 VSUBS 0.025511f
C100 VN.n50 VSUBS 0.025511f
C101 VN.n51 VSUBS 0.024776f
C102 VN.n52 VSUBS 0.047547f
C103 VN.n53 VSUBS 0.047547f
C104 VN.n54 VSUBS 0.025511f
C105 VN.n55 VSUBS 0.025511f
C106 VN.n56 VSUBS 0.025511f
C107 VN.n57 VSUBS 0.039375f
C108 VN.n58 VSUBS 0.047547f
C109 VN.n59 VSUBS 0.045433f
C110 VN.n60 VSUBS 0.041175f
C111 VN.n61 VSUBS 1.63944f
C112 VDD1.t4 VSUBS 0.312286f
C113 VDD1.t7 VSUBS 0.312286f
C114 VDD1.n0 VSUBS 2.49046f
C115 VDD1.t3 VSUBS 0.312286f
C116 VDD1.t6 VSUBS 0.312286f
C117 VDD1.n1 VSUBS 2.48868f
C118 VDD1.t5 VSUBS 0.312286f
C119 VDD1.t0 VSUBS 0.312286f
C120 VDD1.n2 VSUBS 2.48868f
C121 VDD1.n3 VSUBS 5.11993f
C122 VDD1.t1 VSUBS 0.312286f
C123 VDD1.t2 VSUBS 0.312286f
C124 VDD1.n4 VSUBS 2.46855f
C125 VDD1.n5 VSUBS 4.24606f
C126 VTAIL.t4 VSUBS 0.261164f
C127 VTAIL.t0 VSUBS 0.261164f
C128 VTAIL.n0 VSUBS 1.91894f
C129 VTAIL.n1 VSUBS 0.84283f
C130 VTAIL.t3 VSUBS 2.52924f
C131 VTAIL.n2 VSUBS 0.978131f
C132 VTAIL.t9 VSUBS 2.52924f
C133 VTAIL.n3 VSUBS 0.978131f
C134 VTAIL.t10 VSUBS 0.261164f
C135 VTAIL.t14 VSUBS 0.261164f
C136 VTAIL.n4 VSUBS 1.91894f
C137 VTAIL.n5 VSUBS 1.08037f
C138 VTAIL.t7 VSUBS 2.52924f
C139 VTAIL.n6 VSUBS 2.44176f
C140 VTAIL.t5 VSUBS 2.52925f
C141 VTAIL.n7 VSUBS 2.44175f
C142 VTAIL.t1 VSUBS 0.261164f
C143 VTAIL.t2 VSUBS 0.261164f
C144 VTAIL.n8 VSUBS 1.91894f
C145 VTAIL.n9 VSUBS 1.08036f
C146 VTAIL.t15 VSUBS 2.52925f
C147 VTAIL.n10 VSUBS 0.978123f
C148 VTAIL.t13 VSUBS 2.52925f
C149 VTAIL.n11 VSUBS 0.978123f
C150 VTAIL.t12 VSUBS 0.261164f
C151 VTAIL.t11 VSUBS 0.261164f
C152 VTAIL.n12 VSUBS 1.91894f
C153 VTAIL.n13 VSUBS 1.08036f
C154 VTAIL.t8 VSUBS 2.52924f
C155 VTAIL.n14 VSUBS 2.44176f
C156 VTAIL.t6 VSUBS 2.52924f
C157 VTAIL.n15 VSUBS 2.43705f
C158 VP.t7 VSUBS 3.13142f
C159 VP.n0 VSUBS 1.21534f
C160 VP.n1 VSUBS 0.027765f
C161 VP.n2 VSUBS 0.038211f
C162 VP.n3 VSUBS 0.027765f
C163 VP.t2 VSUBS 3.13142f
C164 VP.n4 VSUBS 1.0965f
C165 VP.n5 VSUBS 0.027765f
C166 VP.n6 VSUBS 0.040532f
C167 VP.n7 VSUBS 0.027765f
C168 VP.t1 VSUBS 3.13142f
C169 VP.n8 VSUBS 0.051747f
C170 VP.n9 VSUBS 0.027765f
C171 VP.n10 VSUBS 0.051747f
C172 VP.t5 VSUBS 3.13142f
C173 VP.n11 VSUBS 1.21534f
C174 VP.n12 VSUBS 0.027765f
C175 VP.n13 VSUBS 0.038211f
C176 VP.n14 VSUBS 0.027765f
C177 VP.t6 VSUBS 3.13142f
C178 VP.n15 VSUBS 1.0965f
C179 VP.n16 VSUBS 0.027765f
C180 VP.n17 VSUBS 0.040532f
C181 VP.n18 VSUBS 0.31617f
C182 VP.t0 VSUBS 3.13142f
C183 VP.t3 VSUBS 3.45444f
C184 VP.n19 VSUBS 1.14086f
C185 VP.n20 VSUBS 1.20058f
C186 VP.n21 VSUBS 0.050979f
C187 VP.n22 VSUBS 0.051747f
C188 VP.n23 VSUBS 0.027765f
C189 VP.n24 VSUBS 0.027765f
C190 VP.n25 VSUBS 0.027765f
C191 VP.n26 VSUBS 0.040532f
C192 VP.n27 VSUBS 0.051747f
C193 VP.n28 VSUBS 0.050979f
C194 VP.n29 VSUBS 0.027765f
C195 VP.n30 VSUBS 0.027765f
C196 VP.n31 VSUBS 0.026964f
C197 VP.n32 VSUBS 0.051747f
C198 VP.n33 VSUBS 0.051747f
C199 VP.n34 VSUBS 0.027765f
C200 VP.n35 VSUBS 0.027765f
C201 VP.n36 VSUBS 0.027765f
C202 VP.n37 VSUBS 0.042853f
C203 VP.n38 VSUBS 0.051747f
C204 VP.n39 VSUBS 0.049446f
C205 VP.n40 VSUBS 0.044812f
C206 VP.n41 VSUBS 1.77323f
C207 VP.n42 VSUBS 1.79155f
C208 VP.t4 VSUBS 3.13142f
C209 VP.n43 VSUBS 1.21534f
C210 VP.n44 VSUBS 0.049446f
C211 VP.n45 VSUBS 0.044812f
C212 VP.n46 VSUBS 0.027765f
C213 VP.n47 VSUBS 0.027765f
C214 VP.n48 VSUBS 0.042853f
C215 VP.n49 VSUBS 0.038211f
C216 VP.n50 VSUBS 0.051747f
C217 VP.n51 VSUBS 0.027765f
C218 VP.n52 VSUBS 0.027765f
C219 VP.n53 VSUBS 0.027765f
C220 VP.n54 VSUBS 0.026964f
C221 VP.n55 VSUBS 1.0965f
C222 VP.n56 VSUBS 0.050979f
C223 VP.n57 VSUBS 0.051747f
C224 VP.n58 VSUBS 0.027765f
C225 VP.n59 VSUBS 0.027765f
C226 VP.n60 VSUBS 0.027765f
C227 VP.n61 VSUBS 0.040532f
C228 VP.n62 VSUBS 0.051747f
C229 VP.n63 VSUBS 0.050979f
C230 VP.n64 VSUBS 0.027765f
C231 VP.n65 VSUBS 0.027765f
C232 VP.n66 VSUBS 0.026964f
C233 VP.n67 VSUBS 0.051747f
C234 VP.n68 VSUBS 0.051747f
C235 VP.n69 VSUBS 0.027765f
C236 VP.n70 VSUBS 0.027765f
C237 VP.n71 VSUBS 0.027765f
C238 VP.n72 VSUBS 0.042853f
C239 VP.n73 VSUBS 0.051747f
C240 VP.n74 VSUBS 0.049446f
C241 VP.n75 VSUBS 0.044812f
C242 VP.n76 VSUBS 0.055912f
C243 B.n0 VSUBS 0.004524f
C244 B.n1 VSUBS 0.004524f
C245 B.n2 VSUBS 0.007155f
C246 B.n3 VSUBS 0.007155f
C247 B.n4 VSUBS 0.007155f
C248 B.n5 VSUBS 0.007155f
C249 B.n6 VSUBS 0.007155f
C250 B.n7 VSUBS 0.007155f
C251 B.n8 VSUBS 0.007155f
C252 B.n9 VSUBS 0.007155f
C253 B.n10 VSUBS 0.007155f
C254 B.n11 VSUBS 0.007155f
C255 B.n12 VSUBS 0.007155f
C256 B.n13 VSUBS 0.007155f
C257 B.n14 VSUBS 0.007155f
C258 B.n15 VSUBS 0.007155f
C259 B.n16 VSUBS 0.007155f
C260 B.n17 VSUBS 0.007155f
C261 B.n18 VSUBS 0.007155f
C262 B.n19 VSUBS 0.007155f
C263 B.n20 VSUBS 0.007155f
C264 B.n21 VSUBS 0.007155f
C265 B.n22 VSUBS 0.007155f
C266 B.n23 VSUBS 0.007155f
C267 B.n24 VSUBS 0.007155f
C268 B.n25 VSUBS 0.007155f
C269 B.n26 VSUBS 0.007155f
C270 B.n27 VSUBS 0.007155f
C271 B.n28 VSUBS 0.007155f
C272 B.n29 VSUBS 0.007155f
C273 B.n30 VSUBS 0.007155f
C274 B.n31 VSUBS 0.015745f
C275 B.n32 VSUBS 0.007155f
C276 B.n33 VSUBS 0.007155f
C277 B.n34 VSUBS 0.007155f
C278 B.n35 VSUBS 0.007155f
C279 B.n36 VSUBS 0.007155f
C280 B.n37 VSUBS 0.007155f
C281 B.n38 VSUBS 0.007155f
C282 B.n39 VSUBS 0.007155f
C283 B.n40 VSUBS 0.007155f
C284 B.n41 VSUBS 0.007155f
C285 B.n42 VSUBS 0.007155f
C286 B.n43 VSUBS 0.007155f
C287 B.n44 VSUBS 0.007155f
C288 B.n45 VSUBS 0.007155f
C289 B.n46 VSUBS 0.007155f
C290 B.n47 VSUBS 0.007155f
C291 B.n48 VSUBS 0.007155f
C292 B.n49 VSUBS 0.007155f
C293 B.n50 VSUBS 0.007155f
C294 B.n51 VSUBS 0.007155f
C295 B.n52 VSUBS 0.007155f
C296 B.n53 VSUBS 0.007155f
C297 B.t5 VSUBS 0.442144f
C298 B.t4 VSUBS 0.466836f
C299 B.t3 VSUBS 1.93571f
C300 B.n54 VSUBS 0.25941f
C301 B.n55 VSUBS 0.075739f
C302 B.n56 VSUBS 0.016577f
C303 B.n57 VSUBS 0.007155f
C304 B.n58 VSUBS 0.007155f
C305 B.n59 VSUBS 0.007155f
C306 B.n60 VSUBS 0.007155f
C307 B.n61 VSUBS 0.007155f
C308 B.t8 VSUBS 0.442134f
C309 B.t7 VSUBS 0.466828f
C310 B.t6 VSUBS 1.93571f
C311 B.n62 VSUBS 0.259418f
C312 B.n63 VSUBS 0.075749f
C313 B.n64 VSUBS 0.007155f
C314 B.n65 VSUBS 0.007155f
C315 B.n66 VSUBS 0.007155f
C316 B.n67 VSUBS 0.007155f
C317 B.n68 VSUBS 0.007155f
C318 B.n69 VSUBS 0.007155f
C319 B.n70 VSUBS 0.007155f
C320 B.n71 VSUBS 0.007155f
C321 B.n72 VSUBS 0.007155f
C322 B.n73 VSUBS 0.007155f
C323 B.n74 VSUBS 0.007155f
C324 B.n75 VSUBS 0.007155f
C325 B.n76 VSUBS 0.007155f
C326 B.n77 VSUBS 0.007155f
C327 B.n78 VSUBS 0.007155f
C328 B.n79 VSUBS 0.007155f
C329 B.n80 VSUBS 0.007155f
C330 B.n81 VSUBS 0.007155f
C331 B.n82 VSUBS 0.007155f
C332 B.n83 VSUBS 0.007155f
C333 B.n84 VSUBS 0.007155f
C334 B.n85 VSUBS 0.007155f
C335 B.n86 VSUBS 0.016616f
C336 B.n87 VSUBS 0.007155f
C337 B.n88 VSUBS 0.007155f
C338 B.n89 VSUBS 0.007155f
C339 B.n90 VSUBS 0.007155f
C340 B.n91 VSUBS 0.007155f
C341 B.n92 VSUBS 0.007155f
C342 B.n93 VSUBS 0.007155f
C343 B.n94 VSUBS 0.007155f
C344 B.n95 VSUBS 0.007155f
C345 B.n96 VSUBS 0.007155f
C346 B.n97 VSUBS 0.007155f
C347 B.n98 VSUBS 0.007155f
C348 B.n99 VSUBS 0.007155f
C349 B.n100 VSUBS 0.007155f
C350 B.n101 VSUBS 0.007155f
C351 B.n102 VSUBS 0.007155f
C352 B.n103 VSUBS 0.007155f
C353 B.n104 VSUBS 0.007155f
C354 B.n105 VSUBS 0.007155f
C355 B.n106 VSUBS 0.007155f
C356 B.n107 VSUBS 0.007155f
C357 B.n108 VSUBS 0.007155f
C358 B.n109 VSUBS 0.007155f
C359 B.n110 VSUBS 0.007155f
C360 B.n111 VSUBS 0.007155f
C361 B.n112 VSUBS 0.007155f
C362 B.n113 VSUBS 0.007155f
C363 B.n114 VSUBS 0.007155f
C364 B.n115 VSUBS 0.007155f
C365 B.n116 VSUBS 0.007155f
C366 B.n117 VSUBS 0.007155f
C367 B.n118 VSUBS 0.007155f
C368 B.n119 VSUBS 0.007155f
C369 B.n120 VSUBS 0.007155f
C370 B.n121 VSUBS 0.007155f
C371 B.n122 VSUBS 0.007155f
C372 B.n123 VSUBS 0.007155f
C373 B.n124 VSUBS 0.007155f
C374 B.n125 VSUBS 0.007155f
C375 B.n126 VSUBS 0.007155f
C376 B.n127 VSUBS 0.007155f
C377 B.n128 VSUBS 0.007155f
C378 B.n129 VSUBS 0.007155f
C379 B.n130 VSUBS 0.007155f
C380 B.n131 VSUBS 0.007155f
C381 B.n132 VSUBS 0.007155f
C382 B.n133 VSUBS 0.007155f
C383 B.n134 VSUBS 0.007155f
C384 B.n135 VSUBS 0.007155f
C385 B.n136 VSUBS 0.007155f
C386 B.n137 VSUBS 0.007155f
C387 B.n138 VSUBS 0.007155f
C388 B.n139 VSUBS 0.007155f
C389 B.n140 VSUBS 0.007155f
C390 B.n141 VSUBS 0.007155f
C391 B.n142 VSUBS 0.007155f
C392 B.n143 VSUBS 0.007155f
C393 B.n144 VSUBS 0.007155f
C394 B.n145 VSUBS 0.015745f
C395 B.n146 VSUBS 0.007155f
C396 B.n147 VSUBS 0.007155f
C397 B.n148 VSUBS 0.007155f
C398 B.n149 VSUBS 0.007155f
C399 B.n150 VSUBS 0.007155f
C400 B.n151 VSUBS 0.007155f
C401 B.n152 VSUBS 0.007155f
C402 B.n153 VSUBS 0.007155f
C403 B.n154 VSUBS 0.007155f
C404 B.n155 VSUBS 0.007155f
C405 B.n156 VSUBS 0.007155f
C406 B.n157 VSUBS 0.007155f
C407 B.n158 VSUBS 0.007155f
C408 B.n159 VSUBS 0.007155f
C409 B.n160 VSUBS 0.007155f
C410 B.n161 VSUBS 0.007155f
C411 B.n162 VSUBS 0.007155f
C412 B.n163 VSUBS 0.007155f
C413 B.n164 VSUBS 0.007155f
C414 B.n165 VSUBS 0.007155f
C415 B.n166 VSUBS 0.007155f
C416 B.n167 VSUBS 0.007155f
C417 B.t1 VSUBS 0.442134f
C418 B.t2 VSUBS 0.466828f
C419 B.t0 VSUBS 1.93571f
C420 B.n168 VSUBS 0.259418f
C421 B.n169 VSUBS 0.075749f
C422 B.n170 VSUBS 0.016577f
C423 B.n171 VSUBS 0.007155f
C424 B.n172 VSUBS 0.007155f
C425 B.n173 VSUBS 0.007155f
C426 B.n174 VSUBS 0.007155f
C427 B.n175 VSUBS 0.007155f
C428 B.t10 VSUBS 0.442144f
C429 B.t11 VSUBS 0.466836f
C430 B.t9 VSUBS 1.93571f
C431 B.n176 VSUBS 0.25941f
C432 B.n177 VSUBS 0.075739f
C433 B.n178 VSUBS 0.007155f
C434 B.n179 VSUBS 0.007155f
C435 B.n180 VSUBS 0.007155f
C436 B.n181 VSUBS 0.007155f
C437 B.n182 VSUBS 0.007155f
C438 B.n183 VSUBS 0.007155f
C439 B.n184 VSUBS 0.007155f
C440 B.n185 VSUBS 0.007155f
C441 B.n186 VSUBS 0.007155f
C442 B.n187 VSUBS 0.007155f
C443 B.n188 VSUBS 0.007155f
C444 B.n189 VSUBS 0.007155f
C445 B.n190 VSUBS 0.007155f
C446 B.n191 VSUBS 0.007155f
C447 B.n192 VSUBS 0.007155f
C448 B.n193 VSUBS 0.007155f
C449 B.n194 VSUBS 0.007155f
C450 B.n195 VSUBS 0.007155f
C451 B.n196 VSUBS 0.007155f
C452 B.n197 VSUBS 0.007155f
C453 B.n198 VSUBS 0.007155f
C454 B.n199 VSUBS 0.007155f
C455 B.n200 VSUBS 0.015745f
C456 B.n201 VSUBS 0.007155f
C457 B.n202 VSUBS 0.007155f
C458 B.n203 VSUBS 0.007155f
C459 B.n204 VSUBS 0.007155f
C460 B.n205 VSUBS 0.007155f
C461 B.n206 VSUBS 0.007155f
C462 B.n207 VSUBS 0.007155f
C463 B.n208 VSUBS 0.007155f
C464 B.n209 VSUBS 0.007155f
C465 B.n210 VSUBS 0.007155f
C466 B.n211 VSUBS 0.007155f
C467 B.n212 VSUBS 0.007155f
C468 B.n213 VSUBS 0.007155f
C469 B.n214 VSUBS 0.007155f
C470 B.n215 VSUBS 0.007155f
C471 B.n216 VSUBS 0.007155f
C472 B.n217 VSUBS 0.007155f
C473 B.n218 VSUBS 0.007155f
C474 B.n219 VSUBS 0.007155f
C475 B.n220 VSUBS 0.007155f
C476 B.n221 VSUBS 0.007155f
C477 B.n222 VSUBS 0.007155f
C478 B.n223 VSUBS 0.007155f
C479 B.n224 VSUBS 0.007155f
C480 B.n225 VSUBS 0.007155f
C481 B.n226 VSUBS 0.007155f
C482 B.n227 VSUBS 0.007155f
C483 B.n228 VSUBS 0.007155f
C484 B.n229 VSUBS 0.007155f
C485 B.n230 VSUBS 0.007155f
C486 B.n231 VSUBS 0.007155f
C487 B.n232 VSUBS 0.007155f
C488 B.n233 VSUBS 0.007155f
C489 B.n234 VSUBS 0.007155f
C490 B.n235 VSUBS 0.007155f
C491 B.n236 VSUBS 0.007155f
C492 B.n237 VSUBS 0.007155f
C493 B.n238 VSUBS 0.007155f
C494 B.n239 VSUBS 0.007155f
C495 B.n240 VSUBS 0.007155f
C496 B.n241 VSUBS 0.007155f
C497 B.n242 VSUBS 0.007155f
C498 B.n243 VSUBS 0.007155f
C499 B.n244 VSUBS 0.007155f
C500 B.n245 VSUBS 0.007155f
C501 B.n246 VSUBS 0.007155f
C502 B.n247 VSUBS 0.007155f
C503 B.n248 VSUBS 0.007155f
C504 B.n249 VSUBS 0.007155f
C505 B.n250 VSUBS 0.007155f
C506 B.n251 VSUBS 0.007155f
C507 B.n252 VSUBS 0.007155f
C508 B.n253 VSUBS 0.007155f
C509 B.n254 VSUBS 0.007155f
C510 B.n255 VSUBS 0.007155f
C511 B.n256 VSUBS 0.007155f
C512 B.n257 VSUBS 0.007155f
C513 B.n258 VSUBS 0.007155f
C514 B.n259 VSUBS 0.007155f
C515 B.n260 VSUBS 0.007155f
C516 B.n261 VSUBS 0.007155f
C517 B.n262 VSUBS 0.007155f
C518 B.n263 VSUBS 0.007155f
C519 B.n264 VSUBS 0.007155f
C520 B.n265 VSUBS 0.007155f
C521 B.n266 VSUBS 0.007155f
C522 B.n267 VSUBS 0.007155f
C523 B.n268 VSUBS 0.007155f
C524 B.n269 VSUBS 0.007155f
C525 B.n270 VSUBS 0.007155f
C526 B.n271 VSUBS 0.007155f
C527 B.n272 VSUBS 0.007155f
C528 B.n273 VSUBS 0.007155f
C529 B.n274 VSUBS 0.007155f
C530 B.n275 VSUBS 0.007155f
C531 B.n276 VSUBS 0.007155f
C532 B.n277 VSUBS 0.007155f
C533 B.n278 VSUBS 0.007155f
C534 B.n279 VSUBS 0.007155f
C535 B.n280 VSUBS 0.007155f
C536 B.n281 VSUBS 0.007155f
C537 B.n282 VSUBS 0.007155f
C538 B.n283 VSUBS 0.007155f
C539 B.n284 VSUBS 0.007155f
C540 B.n285 VSUBS 0.007155f
C541 B.n286 VSUBS 0.007155f
C542 B.n287 VSUBS 0.007155f
C543 B.n288 VSUBS 0.007155f
C544 B.n289 VSUBS 0.007155f
C545 B.n290 VSUBS 0.007155f
C546 B.n291 VSUBS 0.007155f
C547 B.n292 VSUBS 0.007155f
C548 B.n293 VSUBS 0.007155f
C549 B.n294 VSUBS 0.007155f
C550 B.n295 VSUBS 0.007155f
C551 B.n296 VSUBS 0.007155f
C552 B.n297 VSUBS 0.007155f
C553 B.n298 VSUBS 0.007155f
C554 B.n299 VSUBS 0.007155f
C555 B.n300 VSUBS 0.007155f
C556 B.n301 VSUBS 0.007155f
C557 B.n302 VSUBS 0.007155f
C558 B.n303 VSUBS 0.007155f
C559 B.n304 VSUBS 0.007155f
C560 B.n305 VSUBS 0.007155f
C561 B.n306 VSUBS 0.007155f
C562 B.n307 VSUBS 0.007155f
C563 B.n308 VSUBS 0.007155f
C564 B.n309 VSUBS 0.007155f
C565 B.n310 VSUBS 0.007155f
C566 B.n311 VSUBS 0.007155f
C567 B.n312 VSUBS 0.007155f
C568 B.n313 VSUBS 0.007155f
C569 B.n314 VSUBS 0.007155f
C570 B.n315 VSUBS 0.015745f
C571 B.n316 VSUBS 0.017083f
C572 B.n317 VSUBS 0.017083f
C573 B.n318 VSUBS 0.007155f
C574 B.n319 VSUBS 0.007155f
C575 B.n320 VSUBS 0.007155f
C576 B.n321 VSUBS 0.007155f
C577 B.n322 VSUBS 0.007155f
C578 B.n323 VSUBS 0.007155f
C579 B.n324 VSUBS 0.007155f
C580 B.n325 VSUBS 0.007155f
C581 B.n326 VSUBS 0.007155f
C582 B.n327 VSUBS 0.007155f
C583 B.n328 VSUBS 0.007155f
C584 B.n329 VSUBS 0.007155f
C585 B.n330 VSUBS 0.007155f
C586 B.n331 VSUBS 0.007155f
C587 B.n332 VSUBS 0.007155f
C588 B.n333 VSUBS 0.007155f
C589 B.n334 VSUBS 0.007155f
C590 B.n335 VSUBS 0.007155f
C591 B.n336 VSUBS 0.007155f
C592 B.n337 VSUBS 0.007155f
C593 B.n338 VSUBS 0.007155f
C594 B.n339 VSUBS 0.007155f
C595 B.n340 VSUBS 0.007155f
C596 B.n341 VSUBS 0.007155f
C597 B.n342 VSUBS 0.007155f
C598 B.n343 VSUBS 0.007155f
C599 B.n344 VSUBS 0.007155f
C600 B.n345 VSUBS 0.007155f
C601 B.n346 VSUBS 0.007155f
C602 B.n347 VSUBS 0.007155f
C603 B.n348 VSUBS 0.007155f
C604 B.n349 VSUBS 0.007155f
C605 B.n350 VSUBS 0.007155f
C606 B.n351 VSUBS 0.007155f
C607 B.n352 VSUBS 0.007155f
C608 B.n353 VSUBS 0.007155f
C609 B.n354 VSUBS 0.007155f
C610 B.n355 VSUBS 0.007155f
C611 B.n356 VSUBS 0.007155f
C612 B.n357 VSUBS 0.007155f
C613 B.n358 VSUBS 0.007155f
C614 B.n359 VSUBS 0.007155f
C615 B.n360 VSUBS 0.007155f
C616 B.n361 VSUBS 0.007155f
C617 B.n362 VSUBS 0.007155f
C618 B.n363 VSUBS 0.007155f
C619 B.n364 VSUBS 0.007155f
C620 B.n365 VSUBS 0.007155f
C621 B.n366 VSUBS 0.007155f
C622 B.n367 VSUBS 0.007155f
C623 B.n368 VSUBS 0.007155f
C624 B.n369 VSUBS 0.007155f
C625 B.n370 VSUBS 0.007155f
C626 B.n371 VSUBS 0.007155f
C627 B.n372 VSUBS 0.007155f
C628 B.n373 VSUBS 0.007155f
C629 B.n374 VSUBS 0.007155f
C630 B.n375 VSUBS 0.007155f
C631 B.n376 VSUBS 0.007155f
C632 B.n377 VSUBS 0.007155f
C633 B.n378 VSUBS 0.007155f
C634 B.n379 VSUBS 0.007155f
C635 B.n380 VSUBS 0.007155f
C636 B.n381 VSUBS 0.007155f
C637 B.n382 VSUBS 0.007155f
C638 B.n383 VSUBS 0.006734f
C639 B.n384 VSUBS 0.016577f
C640 B.n385 VSUBS 0.003998f
C641 B.n386 VSUBS 0.007155f
C642 B.n387 VSUBS 0.007155f
C643 B.n388 VSUBS 0.007155f
C644 B.n389 VSUBS 0.007155f
C645 B.n390 VSUBS 0.007155f
C646 B.n391 VSUBS 0.007155f
C647 B.n392 VSUBS 0.007155f
C648 B.n393 VSUBS 0.007155f
C649 B.n394 VSUBS 0.007155f
C650 B.n395 VSUBS 0.007155f
C651 B.n396 VSUBS 0.007155f
C652 B.n397 VSUBS 0.007155f
C653 B.n398 VSUBS 0.003998f
C654 B.n399 VSUBS 0.007155f
C655 B.n400 VSUBS 0.007155f
C656 B.n401 VSUBS 0.006734f
C657 B.n402 VSUBS 0.007155f
C658 B.n403 VSUBS 0.007155f
C659 B.n404 VSUBS 0.007155f
C660 B.n405 VSUBS 0.007155f
C661 B.n406 VSUBS 0.007155f
C662 B.n407 VSUBS 0.007155f
C663 B.n408 VSUBS 0.007155f
C664 B.n409 VSUBS 0.007155f
C665 B.n410 VSUBS 0.007155f
C666 B.n411 VSUBS 0.007155f
C667 B.n412 VSUBS 0.007155f
C668 B.n413 VSUBS 0.007155f
C669 B.n414 VSUBS 0.007155f
C670 B.n415 VSUBS 0.007155f
C671 B.n416 VSUBS 0.007155f
C672 B.n417 VSUBS 0.007155f
C673 B.n418 VSUBS 0.007155f
C674 B.n419 VSUBS 0.007155f
C675 B.n420 VSUBS 0.007155f
C676 B.n421 VSUBS 0.007155f
C677 B.n422 VSUBS 0.007155f
C678 B.n423 VSUBS 0.007155f
C679 B.n424 VSUBS 0.007155f
C680 B.n425 VSUBS 0.007155f
C681 B.n426 VSUBS 0.007155f
C682 B.n427 VSUBS 0.007155f
C683 B.n428 VSUBS 0.007155f
C684 B.n429 VSUBS 0.007155f
C685 B.n430 VSUBS 0.007155f
C686 B.n431 VSUBS 0.007155f
C687 B.n432 VSUBS 0.007155f
C688 B.n433 VSUBS 0.007155f
C689 B.n434 VSUBS 0.007155f
C690 B.n435 VSUBS 0.007155f
C691 B.n436 VSUBS 0.007155f
C692 B.n437 VSUBS 0.007155f
C693 B.n438 VSUBS 0.007155f
C694 B.n439 VSUBS 0.007155f
C695 B.n440 VSUBS 0.007155f
C696 B.n441 VSUBS 0.007155f
C697 B.n442 VSUBS 0.007155f
C698 B.n443 VSUBS 0.007155f
C699 B.n444 VSUBS 0.007155f
C700 B.n445 VSUBS 0.007155f
C701 B.n446 VSUBS 0.007155f
C702 B.n447 VSUBS 0.007155f
C703 B.n448 VSUBS 0.007155f
C704 B.n449 VSUBS 0.007155f
C705 B.n450 VSUBS 0.007155f
C706 B.n451 VSUBS 0.007155f
C707 B.n452 VSUBS 0.007155f
C708 B.n453 VSUBS 0.007155f
C709 B.n454 VSUBS 0.007155f
C710 B.n455 VSUBS 0.007155f
C711 B.n456 VSUBS 0.007155f
C712 B.n457 VSUBS 0.007155f
C713 B.n458 VSUBS 0.007155f
C714 B.n459 VSUBS 0.007155f
C715 B.n460 VSUBS 0.007155f
C716 B.n461 VSUBS 0.007155f
C717 B.n462 VSUBS 0.007155f
C718 B.n463 VSUBS 0.007155f
C719 B.n464 VSUBS 0.007155f
C720 B.n465 VSUBS 0.007155f
C721 B.n466 VSUBS 0.017083f
C722 B.n467 VSUBS 0.017083f
C723 B.n468 VSUBS 0.015745f
C724 B.n469 VSUBS 0.007155f
C725 B.n470 VSUBS 0.007155f
C726 B.n471 VSUBS 0.007155f
C727 B.n472 VSUBS 0.007155f
C728 B.n473 VSUBS 0.007155f
C729 B.n474 VSUBS 0.007155f
C730 B.n475 VSUBS 0.007155f
C731 B.n476 VSUBS 0.007155f
C732 B.n477 VSUBS 0.007155f
C733 B.n478 VSUBS 0.007155f
C734 B.n479 VSUBS 0.007155f
C735 B.n480 VSUBS 0.007155f
C736 B.n481 VSUBS 0.007155f
C737 B.n482 VSUBS 0.007155f
C738 B.n483 VSUBS 0.007155f
C739 B.n484 VSUBS 0.007155f
C740 B.n485 VSUBS 0.007155f
C741 B.n486 VSUBS 0.007155f
C742 B.n487 VSUBS 0.007155f
C743 B.n488 VSUBS 0.007155f
C744 B.n489 VSUBS 0.007155f
C745 B.n490 VSUBS 0.007155f
C746 B.n491 VSUBS 0.007155f
C747 B.n492 VSUBS 0.007155f
C748 B.n493 VSUBS 0.007155f
C749 B.n494 VSUBS 0.007155f
C750 B.n495 VSUBS 0.007155f
C751 B.n496 VSUBS 0.007155f
C752 B.n497 VSUBS 0.007155f
C753 B.n498 VSUBS 0.007155f
C754 B.n499 VSUBS 0.007155f
C755 B.n500 VSUBS 0.007155f
C756 B.n501 VSUBS 0.007155f
C757 B.n502 VSUBS 0.007155f
C758 B.n503 VSUBS 0.007155f
C759 B.n504 VSUBS 0.007155f
C760 B.n505 VSUBS 0.007155f
C761 B.n506 VSUBS 0.007155f
C762 B.n507 VSUBS 0.007155f
C763 B.n508 VSUBS 0.007155f
C764 B.n509 VSUBS 0.007155f
C765 B.n510 VSUBS 0.007155f
C766 B.n511 VSUBS 0.007155f
C767 B.n512 VSUBS 0.007155f
C768 B.n513 VSUBS 0.007155f
C769 B.n514 VSUBS 0.007155f
C770 B.n515 VSUBS 0.007155f
C771 B.n516 VSUBS 0.007155f
C772 B.n517 VSUBS 0.007155f
C773 B.n518 VSUBS 0.007155f
C774 B.n519 VSUBS 0.007155f
C775 B.n520 VSUBS 0.007155f
C776 B.n521 VSUBS 0.007155f
C777 B.n522 VSUBS 0.007155f
C778 B.n523 VSUBS 0.007155f
C779 B.n524 VSUBS 0.007155f
C780 B.n525 VSUBS 0.007155f
C781 B.n526 VSUBS 0.007155f
C782 B.n527 VSUBS 0.007155f
C783 B.n528 VSUBS 0.007155f
C784 B.n529 VSUBS 0.007155f
C785 B.n530 VSUBS 0.007155f
C786 B.n531 VSUBS 0.007155f
C787 B.n532 VSUBS 0.007155f
C788 B.n533 VSUBS 0.007155f
C789 B.n534 VSUBS 0.007155f
C790 B.n535 VSUBS 0.007155f
C791 B.n536 VSUBS 0.007155f
C792 B.n537 VSUBS 0.007155f
C793 B.n538 VSUBS 0.007155f
C794 B.n539 VSUBS 0.007155f
C795 B.n540 VSUBS 0.007155f
C796 B.n541 VSUBS 0.007155f
C797 B.n542 VSUBS 0.007155f
C798 B.n543 VSUBS 0.007155f
C799 B.n544 VSUBS 0.007155f
C800 B.n545 VSUBS 0.007155f
C801 B.n546 VSUBS 0.007155f
C802 B.n547 VSUBS 0.007155f
C803 B.n548 VSUBS 0.007155f
C804 B.n549 VSUBS 0.007155f
C805 B.n550 VSUBS 0.007155f
C806 B.n551 VSUBS 0.007155f
C807 B.n552 VSUBS 0.007155f
C808 B.n553 VSUBS 0.007155f
C809 B.n554 VSUBS 0.007155f
C810 B.n555 VSUBS 0.007155f
C811 B.n556 VSUBS 0.007155f
C812 B.n557 VSUBS 0.007155f
C813 B.n558 VSUBS 0.007155f
C814 B.n559 VSUBS 0.007155f
C815 B.n560 VSUBS 0.007155f
C816 B.n561 VSUBS 0.007155f
C817 B.n562 VSUBS 0.007155f
C818 B.n563 VSUBS 0.007155f
C819 B.n564 VSUBS 0.007155f
C820 B.n565 VSUBS 0.007155f
C821 B.n566 VSUBS 0.007155f
C822 B.n567 VSUBS 0.007155f
C823 B.n568 VSUBS 0.007155f
C824 B.n569 VSUBS 0.007155f
C825 B.n570 VSUBS 0.007155f
C826 B.n571 VSUBS 0.007155f
C827 B.n572 VSUBS 0.007155f
C828 B.n573 VSUBS 0.007155f
C829 B.n574 VSUBS 0.007155f
C830 B.n575 VSUBS 0.007155f
C831 B.n576 VSUBS 0.007155f
C832 B.n577 VSUBS 0.007155f
C833 B.n578 VSUBS 0.007155f
C834 B.n579 VSUBS 0.007155f
C835 B.n580 VSUBS 0.007155f
C836 B.n581 VSUBS 0.007155f
C837 B.n582 VSUBS 0.007155f
C838 B.n583 VSUBS 0.007155f
C839 B.n584 VSUBS 0.007155f
C840 B.n585 VSUBS 0.007155f
C841 B.n586 VSUBS 0.007155f
C842 B.n587 VSUBS 0.007155f
C843 B.n588 VSUBS 0.007155f
C844 B.n589 VSUBS 0.007155f
C845 B.n590 VSUBS 0.007155f
C846 B.n591 VSUBS 0.007155f
C847 B.n592 VSUBS 0.007155f
C848 B.n593 VSUBS 0.007155f
C849 B.n594 VSUBS 0.007155f
C850 B.n595 VSUBS 0.007155f
C851 B.n596 VSUBS 0.007155f
C852 B.n597 VSUBS 0.007155f
C853 B.n598 VSUBS 0.007155f
C854 B.n599 VSUBS 0.007155f
C855 B.n600 VSUBS 0.007155f
C856 B.n601 VSUBS 0.007155f
C857 B.n602 VSUBS 0.007155f
C858 B.n603 VSUBS 0.007155f
C859 B.n604 VSUBS 0.007155f
C860 B.n605 VSUBS 0.007155f
C861 B.n606 VSUBS 0.007155f
C862 B.n607 VSUBS 0.007155f
C863 B.n608 VSUBS 0.007155f
C864 B.n609 VSUBS 0.007155f
C865 B.n610 VSUBS 0.007155f
C866 B.n611 VSUBS 0.007155f
C867 B.n612 VSUBS 0.007155f
C868 B.n613 VSUBS 0.007155f
C869 B.n614 VSUBS 0.007155f
C870 B.n615 VSUBS 0.007155f
C871 B.n616 VSUBS 0.007155f
C872 B.n617 VSUBS 0.007155f
C873 B.n618 VSUBS 0.007155f
C874 B.n619 VSUBS 0.007155f
C875 B.n620 VSUBS 0.007155f
C876 B.n621 VSUBS 0.007155f
C877 B.n622 VSUBS 0.007155f
C878 B.n623 VSUBS 0.007155f
C879 B.n624 VSUBS 0.007155f
C880 B.n625 VSUBS 0.007155f
C881 B.n626 VSUBS 0.007155f
C882 B.n627 VSUBS 0.007155f
C883 B.n628 VSUBS 0.007155f
C884 B.n629 VSUBS 0.007155f
C885 B.n630 VSUBS 0.007155f
C886 B.n631 VSUBS 0.007155f
C887 B.n632 VSUBS 0.007155f
C888 B.n633 VSUBS 0.007155f
C889 B.n634 VSUBS 0.007155f
C890 B.n635 VSUBS 0.007155f
C891 B.n636 VSUBS 0.007155f
C892 B.n637 VSUBS 0.007155f
C893 B.n638 VSUBS 0.007155f
C894 B.n639 VSUBS 0.007155f
C895 B.n640 VSUBS 0.007155f
C896 B.n641 VSUBS 0.007155f
C897 B.n642 VSUBS 0.007155f
C898 B.n643 VSUBS 0.007155f
C899 B.n644 VSUBS 0.007155f
C900 B.n645 VSUBS 0.015745f
C901 B.n646 VSUBS 0.017083f
C902 B.n647 VSUBS 0.016212f
C903 B.n648 VSUBS 0.007155f
C904 B.n649 VSUBS 0.007155f
C905 B.n650 VSUBS 0.007155f
C906 B.n651 VSUBS 0.007155f
C907 B.n652 VSUBS 0.007155f
C908 B.n653 VSUBS 0.007155f
C909 B.n654 VSUBS 0.007155f
C910 B.n655 VSUBS 0.007155f
C911 B.n656 VSUBS 0.007155f
C912 B.n657 VSUBS 0.007155f
C913 B.n658 VSUBS 0.007155f
C914 B.n659 VSUBS 0.007155f
C915 B.n660 VSUBS 0.007155f
C916 B.n661 VSUBS 0.007155f
C917 B.n662 VSUBS 0.007155f
C918 B.n663 VSUBS 0.007155f
C919 B.n664 VSUBS 0.007155f
C920 B.n665 VSUBS 0.007155f
C921 B.n666 VSUBS 0.007155f
C922 B.n667 VSUBS 0.007155f
C923 B.n668 VSUBS 0.007155f
C924 B.n669 VSUBS 0.007155f
C925 B.n670 VSUBS 0.007155f
C926 B.n671 VSUBS 0.007155f
C927 B.n672 VSUBS 0.007155f
C928 B.n673 VSUBS 0.007155f
C929 B.n674 VSUBS 0.007155f
C930 B.n675 VSUBS 0.007155f
C931 B.n676 VSUBS 0.007155f
C932 B.n677 VSUBS 0.007155f
C933 B.n678 VSUBS 0.007155f
C934 B.n679 VSUBS 0.007155f
C935 B.n680 VSUBS 0.007155f
C936 B.n681 VSUBS 0.007155f
C937 B.n682 VSUBS 0.007155f
C938 B.n683 VSUBS 0.007155f
C939 B.n684 VSUBS 0.007155f
C940 B.n685 VSUBS 0.007155f
C941 B.n686 VSUBS 0.007155f
C942 B.n687 VSUBS 0.007155f
C943 B.n688 VSUBS 0.007155f
C944 B.n689 VSUBS 0.007155f
C945 B.n690 VSUBS 0.007155f
C946 B.n691 VSUBS 0.007155f
C947 B.n692 VSUBS 0.007155f
C948 B.n693 VSUBS 0.007155f
C949 B.n694 VSUBS 0.007155f
C950 B.n695 VSUBS 0.007155f
C951 B.n696 VSUBS 0.007155f
C952 B.n697 VSUBS 0.007155f
C953 B.n698 VSUBS 0.007155f
C954 B.n699 VSUBS 0.007155f
C955 B.n700 VSUBS 0.007155f
C956 B.n701 VSUBS 0.007155f
C957 B.n702 VSUBS 0.007155f
C958 B.n703 VSUBS 0.007155f
C959 B.n704 VSUBS 0.007155f
C960 B.n705 VSUBS 0.007155f
C961 B.n706 VSUBS 0.007155f
C962 B.n707 VSUBS 0.007155f
C963 B.n708 VSUBS 0.007155f
C964 B.n709 VSUBS 0.007155f
C965 B.n710 VSUBS 0.007155f
C966 B.n711 VSUBS 0.007155f
C967 B.n712 VSUBS 0.007155f
C968 B.n713 VSUBS 0.006734f
C969 B.n714 VSUBS 0.016577f
C970 B.n715 VSUBS 0.003998f
C971 B.n716 VSUBS 0.007155f
C972 B.n717 VSUBS 0.007155f
C973 B.n718 VSUBS 0.007155f
C974 B.n719 VSUBS 0.007155f
C975 B.n720 VSUBS 0.007155f
C976 B.n721 VSUBS 0.007155f
C977 B.n722 VSUBS 0.007155f
C978 B.n723 VSUBS 0.007155f
C979 B.n724 VSUBS 0.007155f
C980 B.n725 VSUBS 0.007155f
C981 B.n726 VSUBS 0.007155f
C982 B.n727 VSUBS 0.007155f
C983 B.n728 VSUBS 0.003998f
C984 B.n729 VSUBS 0.007155f
C985 B.n730 VSUBS 0.007155f
C986 B.n731 VSUBS 0.006734f
C987 B.n732 VSUBS 0.007155f
C988 B.n733 VSUBS 0.007155f
C989 B.n734 VSUBS 0.007155f
C990 B.n735 VSUBS 0.007155f
C991 B.n736 VSUBS 0.007155f
C992 B.n737 VSUBS 0.007155f
C993 B.n738 VSUBS 0.007155f
C994 B.n739 VSUBS 0.007155f
C995 B.n740 VSUBS 0.007155f
C996 B.n741 VSUBS 0.007155f
C997 B.n742 VSUBS 0.007155f
C998 B.n743 VSUBS 0.007155f
C999 B.n744 VSUBS 0.007155f
C1000 B.n745 VSUBS 0.007155f
C1001 B.n746 VSUBS 0.007155f
C1002 B.n747 VSUBS 0.007155f
C1003 B.n748 VSUBS 0.007155f
C1004 B.n749 VSUBS 0.007155f
C1005 B.n750 VSUBS 0.007155f
C1006 B.n751 VSUBS 0.007155f
C1007 B.n752 VSUBS 0.007155f
C1008 B.n753 VSUBS 0.007155f
C1009 B.n754 VSUBS 0.007155f
C1010 B.n755 VSUBS 0.007155f
C1011 B.n756 VSUBS 0.007155f
C1012 B.n757 VSUBS 0.007155f
C1013 B.n758 VSUBS 0.007155f
C1014 B.n759 VSUBS 0.007155f
C1015 B.n760 VSUBS 0.007155f
C1016 B.n761 VSUBS 0.007155f
C1017 B.n762 VSUBS 0.007155f
C1018 B.n763 VSUBS 0.007155f
C1019 B.n764 VSUBS 0.007155f
C1020 B.n765 VSUBS 0.007155f
C1021 B.n766 VSUBS 0.007155f
C1022 B.n767 VSUBS 0.007155f
C1023 B.n768 VSUBS 0.007155f
C1024 B.n769 VSUBS 0.007155f
C1025 B.n770 VSUBS 0.007155f
C1026 B.n771 VSUBS 0.007155f
C1027 B.n772 VSUBS 0.007155f
C1028 B.n773 VSUBS 0.007155f
C1029 B.n774 VSUBS 0.007155f
C1030 B.n775 VSUBS 0.007155f
C1031 B.n776 VSUBS 0.007155f
C1032 B.n777 VSUBS 0.007155f
C1033 B.n778 VSUBS 0.007155f
C1034 B.n779 VSUBS 0.007155f
C1035 B.n780 VSUBS 0.007155f
C1036 B.n781 VSUBS 0.007155f
C1037 B.n782 VSUBS 0.007155f
C1038 B.n783 VSUBS 0.007155f
C1039 B.n784 VSUBS 0.007155f
C1040 B.n785 VSUBS 0.007155f
C1041 B.n786 VSUBS 0.007155f
C1042 B.n787 VSUBS 0.007155f
C1043 B.n788 VSUBS 0.007155f
C1044 B.n789 VSUBS 0.007155f
C1045 B.n790 VSUBS 0.007155f
C1046 B.n791 VSUBS 0.007155f
C1047 B.n792 VSUBS 0.007155f
C1048 B.n793 VSUBS 0.007155f
C1049 B.n794 VSUBS 0.007155f
C1050 B.n795 VSUBS 0.007155f
C1051 B.n796 VSUBS 0.017083f
C1052 B.n797 VSUBS 0.017083f
C1053 B.n798 VSUBS 0.015745f
C1054 B.n799 VSUBS 0.007155f
C1055 B.n800 VSUBS 0.007155f
C1056 B.n801 VSUBS 0.007155f
C1057 B.n802 VSUBS 0.007155f
C1058 B.n803 VSUBS 0.007155f
C1059 B.n804 VSUBS 0.007155f
C1060 B.n805 VSUBS 0.007155f
C1061 B.n806 VSUBS 0.007155f
C1062 B.n807 VSUBS 0.007155f
C1063 B.n808 VSUBS 0.007155f
C1064 B.n809 VSUBS 0.007155f
C1065 B.n810 VSUBS 0.007155f
C1066 B.n811 VSUBS 0.007155f
C1067 B.n812 VSUBS 0.007155f
C1068 B.n813 VSUBS 0.007155f
C1069 B.n814 VSUBS 0.007155f
C1070 B.n815 VSUBS 0.007155f
C1071 B.n816 VSUBS 0.007155f
C1072 B.n817 VSUBS 0.007155f
C1073 B.n818 VSUBS 0.007155f
C1074 B.n819 VSUBS 0.007155f
C1075 B.n820 VSUBS 0.007155f
C1076 B.n821 VSUBS 0.007155f
C1077 B.n822 VSUBS 0.007155f
C1078 B.n823 VSUBS 0.007155f
C1079 B.n824 VSUBS 0.007155f
C1080 B.n825 VSUBS 0.007155f
C1081 B.n826 VSUBS 0.007155f
C1082 B.n827 VSUBS 0.007155f
C1083 B.n828 VSUBS 0.007155f
C1084 B.n829 VSUBS 0.007155f
C1085 B.n830 VSUBS 0.007155f
C1086 B.n831 VSUBS 0.007155f
C1087 B.n832 VSUBS 0.007155f
C1088 B.n833 VSUBS 0.007155f
C1089 B.n834 VSUBS 0.007155f
C1090 B.n835 VSUBS 0.007155f
C1091 B.n836 VSUBS 0.007155f
C1092 B.n837 VSUBS 0.007155f
C1093 B.n838 VSUBS 0.007155f
C1094 B.n839 VSUBS 0.007155f
C1095 B.n840 VSUBS 0.007155f
C1096 B.n841 VSUBS 0.007155f
C1097 B.n842 VSUBS 0.007155f
C1098 B.n843 VSUBS 0.007155f
C1099 B.n844 VSUBS 0.007155f
C1100 B.n845 VSUBS 0.007155f
C1101 B.n846 VSUBS 0.007155f
C1102 B.n847 VSUBS 0.007155f
C1103 B.n848 VSUBS 0.007155f
C1104 B.n849 VSUBS 0.007155f
C1105 B.n850 VSUBS 0.007155f
C1106 B.n851 VSUBS 0.007155f
C1107 B.n852 VSUBS 0.007155f
C1108 B.n853 VSUBS 0.007155f
C1109 B.n854 VSUBS 0.007155f
C1110 B.n855 VSUBS 0.007155f
C1111 B.n856 VSUBS 0.007155f
C1112 B.n857 VSUBS 0.007155f
C1113 B.n858 VSUBS 0.007155f
C1114 B.n859 VSUBS 0.007155f
C1115 B.n860 VSUBS 0.007155f
C1116 B.n861 VSUBS 0.007155f
C1117 B.n862 VSUBS 0.007155f
C1118 B.n863 VSUBS 0.007155f
C1119 B.n864 VSUBS 0.007155f
C1120 B.n865 VSUBS 0.007155f
C1121 B.n866 VSUBS 0.007155f
C1122 B.n867 VSUBS 0.007155f
C1123 B.n868 VSUBS 0.007155f
C1124 B.n869 VSUBS 0.007155f
C1125 B.n870 VSUBS 0.007155f
C1126 B.n871 VSUBS 0.007155f
C1127 B.n872 VSUBS 0.007155f
C1128 B.n873 VSUBS 0.007155f
C1129 B.n874 VSUBS 0.007155f
C1130 B.n875 VSUBS 0.007155f
C1131 B.n876 VSUBS 0.007155f
C1132 B.n877 VSUBS 0.007155f
C1133 B.n878 VSUBS 0.007155f
C1134 B.n879 VSUBS 0.007155f
C1135 B.n880 VSUBS 0.007155f
C1136 B.n881 VSUBS 0.007155f
C1137 B.n882 VSUBS 0.007155f
C1138 B.n883 VSUBS 0.007155f
C1139 B.n884 VSUBS 0.007155f
C1140 B.n885 VSUBS 0.007155f
C1141 B.n886 VSUBS 0.007155f
C1142 B.n887 VSUBS 0.016201f
.ends

