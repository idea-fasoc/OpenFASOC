* NGSPICE file created from diff_pair_sample_0942.ext - technology: sky130A

.subckt diff_pair_sample_0942 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2704 pd=14.09 as=5.3664 ps=28.3 w=13.76 l=2.98
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=0 ps=0 w=13.76 l=2.98
X2 VTAIL.t5 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=2.2704 ps=14.09 w=13.76 l=2.98
X3 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=2.2704 ps=14.09 w=13.76 l=2.98
X4 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2704 pd=14.09 as=5.3664 ps=28.3 w=13.76 l=2.98
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=0 ps=0 w=13.76 l=2.98
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=0 ps=0 w=13.76 l=2.98
X7 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2704 pd=14.09 as=5.3664 ps=28.3 w=13.76 l=2.98
X8 VTAIL.t7 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=2.2704 ps=14.09 w=13.76 l=2.98
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=0 ps=0 w=13.76 l=2.98
X10 VDD1.t0 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2704 pd=14.09 as=5.3664 ps=28.3 w=13.76 l=2.98
X11 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3664 pd=28.3 as=2.2704 ps=14.09 w=13.76 l=2.98
R0 VP.n15 VP.n14 161.3
R1 VP.n13 VP.n1 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n7 VP.n3 161.3
R6 VP.n4 VP.t1 145.775
R7 VP.n4 VP.t0 144.788
R8 VP.n6 VP.t2 111.281
R9 VP.n0 VP.t3 111.281
R10 VP.n6 VP.n5 70.3262
R11 VP.n16 VP.n0 70.3262
R12 VP.n12 VP.n2 56.5617
R13 VP.n5 VP.n4 51.8729
R14 VP.n8 VP.n7 24.5923
R15 VP.n8 VP.n2 24.5923
R16 VP.n13 VP.n12 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n6 19.9199
R19 VP.n14 VP.n0 19.9199
R20 VP.n5 VP.n3 0.354861
R21 VP.n16 VP.n15 0.354861
R22 VP VP.n16 0.267071
R23 VP.n9 VP.n3 0.189894
R24 VP.n10 VP.n9 0.189894
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n1 0.189894
R27 VP.n15 VP.n1 0.189894
R28 VTAIL.n5 VTAIL.t5 49.7061
R29 VTAIL.n4 VTAIL.t1 49.7061
R30 VTAIL.n3 VTAIL.t0 49.7061
R31 VTAIL.n7 VTAIL.t2 49.7059
R32 VTAIL.n0 VTAIL.t3 49.7059
R33 VTAIL.n1 VTAIL.t4 49.7059
R34 VTAIL.n2 VTAIL.t7 49.7059
R35 VTAIL.n6 VTAIL.t6 49.7059
R36 VTAIL.n7 VTAIL.n6 27.0824
R37 VTAIL.n3 VTAIL.n2 27.0824
R38 VTAIL.n4 VTAIL.n3 2.85395
R39 VTAIL.n6 VTAIL.n5 2.85395
R40 VTAIL.n2 VTAIL.n1 2.85395
R41 VTAIL VTAIL.n0 1.48541
R42 VTAIL VTAIL.n7 1.36903
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 109.608
R46 VDD1 VDD1.n0 65.0039
R47 VDD1.n0 VDD1.t2 1.43945
R48 VDD1.n0 VDD1.t3 1.43945
R49 VDD1.n1 VDD1.t1 1.43945
R50 VDD1.n1 VDD1.t0 1.43945
R51 B.n828 B.n827 585
R52 B.n829 B.n828 585
R53 B.n331 B.n122 585
R54 B.n330 B.n329 585
R55 B.n328 B.n327 585
R56 B.n326 B.n325 585
R57 B.n324 B.n323 585
R58 B.n322 B.n321 585
R59 B.n320 B.n319 585
R60 B.n318 B.n317 585
R61 B.n316 B.n315 585
R62 B.n314 B.n313 585
R63 B.n312 B.n311 585
R64 B.n310 B.n309 585
R65 B.n308 B.n307 585
R66 B.n306 B.n305 585
R67 B.n304 B.n303 585
R68 B.n302 B.n301 585
R69 B.n300 B.n299 585
R70 B.n298 B.n297 585
R71 B.n296 B.n295 585
R72 B.n294 B.n293 585
R73 B.n292 B.n291 585
R74 B.n290 B.n289 585
R75 B.n288 B.n287 585
R76 B.n286 B.n285 585
R77 B.n284 B.n283 585
R78 B.n282 B.n281 585
R79 B.n280 B.n279 585
R80 B.n278 B.n277 585
R81 B.n276 B.n275 585
R82 B.n274 B.n273 585
R83 B.n272 B.n271 585
R84 B.n270 B.n269 585
R85 B.n268 B.n267 585
R86 B.n266 B.n265 585
R87 B.n264 B.n263 585
R88 B.n262 B.n261 585
R89 B.n260 B.n259 585
R90 B.n258 B.n257 585
R91 B.n256 B.n255 585
R92 B.n254 B.n253 585
R93 B.n252 B.n251 585
R94 B.n250 B.n249 585
R95 B.n248 B.n247 585
R96 B.n246 B.n245 585
R97 B.n244 B.n243 585
R98 B.n242 B.n241 585
R99 B.n240 B.n239 585
R100 B.n238 B.n237 585
R101 B.n236 B.n235 585
R102 B.n234 B.n233 585
R103 B.n232 B.n231 585
R104 B.n230 B.n229 585
R105 B.n228 B.n227 585
R106 B.n226 B.n225 585
R107 B.n224 B.n223 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n179 B.n178 585
R130 B.n177 B.n176 585
R131 B.n175 B.n174 585
R132 B.n173 B.n172 585
R133 B.n171 B.n170 585
R134 B.n169 B.n168 585
R135 B.n167 B.n166 585
R136 B.n165 B.n164 585
R137 B.n163 B.n162 585
R138 B.n161 B.n160 585
R139 B.n159 B.n158 585
R140 B.n157 B.n156 585
R141 B.n155 B.n154 585
R142 B.n153 B.n152 585
R143 B.n151 B.n150 585
R144 B.n149 B.n148 585
R145 B.n147 B.n146 585
R146 B.n145 B.n144 585
R147 B.n143 B.n142 585
R148 B.n141 B.n140 585
R149 B.n139 B.n138 585
R150 B.n137 B.n136 585
R151 B.n135 B.n134 585
R152 B.n133 B.n132 585
R153 B.n131 B.n130 585
R154 B.n129 B.n128 585
R155 B.n826 B.n70 585
R156 B.n830 B.n70 585
R157 B.n825 B.n69 585
R158 B.n831 B.n69 585
R159 B.n824 B.n823 585
R160 B.n823 B.n65 585
R161 B.n822 B.n64 585
R162 B.n837 B.n64 585
R163 B.n821 B.n63 585
R164 B.n838 B.n63 585
R165 B.n820 B.n62 585
R166 B.n839 B.n62 585
R167 B.n819 B.n818 585
R168 B.n818 B.n58 585
R169 B.n817 B.n57 585
R170 B.n845 B.n57 585
R171 B.n816 B.n56 585
R172 B.n846 B.n56 585
R173 B.n815 B.n55 585
R174 B.n847 B.n55 585
R175 B.n814 B.n813 585
R176 B.n813 B.n51 585
R177 B.n812 B.n50 585
R178 B.n853 B.n50 585
R179 B.n811 B.n49 585
R180 B.n854 B.n49 585
R181 B.n810 B.n48 585
R182 B.n855 B.n48 585
R183 B.n809 B.n808 585
R184 B.n808 B.n44 585
R185 B.n807 B.n43 585
R186 B.n861 B.n43 585
R187 B.n806 B.n42 585
R188 B.n862 B.n42 585
R189 B.n805 B.n41 585
R190 B.n863 B.n41 585
R191 B.n804 B.n803 585
R192 B.n803 B.n37 585
R193 B.n802 B.n36 585
R194 B.n869 B.n36 585
R195 B.n801 B.n35 585
R196 B.n870 B.n35 585
R197 B.n800 B.n34 585
R198 B.n871 B.n34 585
R199 B.n799 B.n798 585
R200 B.n798 B.n30 585
R201 B.n797 B.n29 585
R202 B.n877 B.n29 585
R203 B.n796 B.n28 585
R204 B.n878 B.n28 585
R205 B.n795 B.n27 585
R206 B.n879 B.n27 585
R207 B.n794 B.n793 585
R208 B.n793 B.n23 585
R209 B.n792 B.n22 585
R210 B.n885 B.n22 585
R211 B.n791 B.n21 585
R212 B.n886 B.n21 585
R213 B.n790 B.n20 585
R214 B.n887 B.n20 585
R215 B.n789 B.n788 585
R216 B.n788 B.n16 585
R217 B.n787 B.n15 585
R218 B.n893 B.n15 585
R219 B.n786 B.n14 585
R220 B.n894 B.n14 585
R221 B.n785 B.n13 585
R222 B.n895 B.n13 585
R223 B.n784 B.n783 585
R224 B.n783 B.n12 585
R225 B.n782 B.n781 585
R226 B.n782 B.n8 585
R227 B.n780 B.n7 585
R228 B.n902 B.n7 585
R229 B.n779 B.n6 585
R230 B.n903 B.n6 585
R231 B.n778 B.n5 585
R232 B.n904 B.n5 585
R233 B.n777 B.n776 585
R234 B.n776 B.n4 585
R235 B.n775 B.n332 585
R236 B.n775 B.n774 585
R237 B.n765 B.n333 585
R238 B.n334 B.n333 585
R239 B.n767 B.n766 585
R240 B.n768 B.n767 585
R241 B.n764 B.n339 585
R242 B.n339 B.n338 585
R243 B.n763 B.n762 585
R244 B.n762 B.n761 585
R245 B.n341 B.n340 585
R246 B.n342 B.n341 585
R247 B.n754 B.n753 585
R248 B.n755 B.n754 585
R249 B.n752 B.n347 585
R250 B.n347 B.n346 585
R251 B.n751 B.n750 585
R252 B.n750 B.n749 585
R253 B.n349 B.n348 585
R254 B.n350 B.n349 585
R255 B.n742 B.n741 585
R256 B.n743 B.n742 585
R257 B.n740 B.n355 585
R258 B.n355 B.n354 585
R259 B.n739 B.n738 585
R260 B.n738 B.n737 585
R261 B.n357 B.n356 585
R262 B.n358 B.n357 585
R263 B.n730 B.n729 585
R264 B.n731 B.n730 585
R265 B.n728 B.n363 585
R266 B.n363 B.n362 585
R267 B.n727 B.n726 585
R268 B.n726 B.n725 585
R269 B.n365 B.n364 585
R270 B.n366 B.n365 585
R271 B.n718 B.n717 585
R272 B.n719 B.n718 585
R273 B.n716 B.n371 585
R274 B.n371 B.n370 585
R275 B.n715 B.n714 585
R276 B.n714 B.n713 585
R277 B.n373 B.n372 585
R278 B.n374 B.n373 585
R279 B.n706 B.n705 585
R280 B.n707 B.n706 585
R281 B.n704 B.n379 585
R282 B.n379 B.n378 585
R283 B.n703 B.n702 585
R284 B.n702 B.n701 585
R285 B.n381 B.n380 585
R286 B.n382 B.n381 585
R287 B.n694 B.n693 585
R288 B.n695 B.n694 585
R289 B.n692 B.n386 585
R290 B.n390 B.n386 585
R291 B.n691 B.n690 585
R292 B.n690 B.n689 585
R293 B.n388 B.n387 585
R294 B.n389 B.n388 585
R295 B.n682 B.n681 585
R296 B.n683 B.n682 585
R297 B.n680 B.n395 585
R298 B.n395 B.n394 585
R299 B.n679 B.n678 585
R300 B.n678 B.n677 585
R301 B.n397 B.n396 585
R302 B.n398 B.n397 585
R303 B.n670 B.n669 585
R304 B.n671 B.n670 585
R305 B.n668 B.n403 585
R306 B.n403 B.n402 585
R307 B.n662 B.n661 585
R308 B.n660 B.n456 585
R309 B.n659 B.n455 585
R310 B.n664 B.n455 585
R311 B.n658 B.n657 585
R312 B.n656 B.n655 585
R313 B.n654 B.n653 585
R314 B.n652 B.n651 585
R315 B.n650 B.n649 585
R316 B.n648 B.n647 585
R317 B.n646 B.n645 585
R318 B.n644 B.n643 585
R319 B.n642 B.n641 585
R320 B.n640 B.n639 585
R321 B.n638 B.n637 585
R322 B.n636 B.n635 585
R323 B.n634 B.n633 585
R324 B.n632 B.n631 585
R325 B.n630 B.n629 585
R326 B.n628 B.n627 585
R327 B.n626 B.n625 585
R328 B.n624 B.n623 585
R329 B.n622 B.n621 585
R330 B.n620 B.n619 585
R331 B.n618 B.n617 585
R332 B.n616 B.n615 585
R333 B.n614 B.n613 585
R334 B.n612 B.n611 585
R335 B.n610 B.n609 585
R336 B.n608 B.n607 585
R337 B.n606 B.n605 585
R338 B.n604 B.n603 585
R339 B.n602 B.n601 585
R340 B.n600 B.n599 585
R341 B.n598 B.n597 585
R342 B.n596 B.n595 585
R343 B.n594 B.n593 585
R344 B.n592 B.n591 585
R345 B.n590 B.n589 585
R346 B.n588 B.n587 585
R347 B.n586 B.n585 585
R348 B.n584 B.n583 585
R349 B.n582 B.n581 585
R350 B.n580 B.n579 585
R351 B.n578 B.n577 585
R352 B.n576 B.n575 585
R353 B.n574 B.n573 585
R354 B.n572 B.n571 585
R355 B.n570 B.n569 585
R356 B.n568 B.n567 585
R357 B.n566 B.n565 585
R358 B.n564 B.n563 585
R359 B.n562 B.n561 585
R360 B.n560 B.n559 585
R361 B.n558 B.n557 585
R362 B.n556 B.n555 585
R363 B.n554 B.n553 585
R364 B.n551 B.n550 585
R365 B.n549 B.n548 585
R366 B.n547 B.n546 585
R367 B.n545 B.n544 585
R368 B.n543 B.n542 585
R369 B.n541 B.n540 585
R370 B.n539 B.n538 585
R371 B.n537 B.n536 585
R372 B.n535 B.n534 585
R373 B.n533 B.n532 585
R374 B.n531 B.n530 585
R375 B.n529 B.n528 585
R376 B.n527 B.n526 585
R377 B.n525 B.n524 585
R378 B.n523 B.n522 585
R379 B.n521 B.n520 585
R380 B.n519 B.n518 585
R381 B.n517 B.n516 585
R382 B.n515 B.n514 585
R383 B.n513 B.n512 585
R384 B.n511 B.n510 585
R385 B.n509 B.n508 585
R386 B.n507 B.n506 585
R387 B.n505 B.n504 585
R388 B.n503 B.n502 585
R389 B.n501 B.n500 585
R390 B.n499 B.n498 585
R391 B.n497 B.n496 585
R392 B.n495 B.n494 585
R393 B.n493 B.n492 585
R394 B.n491 B.n490 585
R395 B.n489 B.n488 585
R396 B.n487 B.n486 585
R397 B.n485 B.n484 585
R398 B.n483 B.n482 585
R399 B.n481 B.n480 585
R400 B.n479 B.n478 585
R401 B.n477 B.n476 585
R402 B.n475 B.n474 585
R403 B.n473 B.n472 585
R404 B.n471 B.n470 585
R405 B.n469 B.n468 585
R406 B.n467 B.n466 585
R407 B.n465 B.n464 585
R408 B.n463 B.n462 585
R409 B.n405 B.n404 585
R410 B.n667 B.n666 585
R411 B.n401 B.n400 585
R412 B.n402 B.n401 585
R413 B.n673 B.n672 585
R414 B.n672 B.n671 585
R415 B.n674 B.n399 585
R416 B.n399 B.n398 585
R417 B.n676 B.n675 585
R418 B.n677 B.n676 585
R419 B.n393 B.n392 585
R420 B.n394 B.n393 585
R421 B.n685 B.n684 585
R422 B.n684 B.n683 585
R423 B.n686 B.n391 585
R424 B.n391 B.n389 585
R425 B.n688 B.n687 585
R426 B.n689 B.n688 585
R427 B.n385 B.n384 585
R428 B.n390 B.n385 585
R429 B.n697 B.n696 585
R430 B.n696 B.n695 585
R431 B.n698 B.n383 585
R432 B.n383 B.n382 585
R433 B.n700 B.n699 585
R434 B.n701 B.n700 585
R435 B.n377 B.n376 585
R436 B.n378 B.n377 585
R437 B.n709 B.n708 585
R438 B.n708 B.n707 585
R439 B.n710 B.n375 585
R440 B.n375 B.n374 585
R441 B.n712 B.n711 585
R442 B.n713 B.n712 585
R443 B.n369 B.n368 585
R444 B.n370 B.n369 585
R445 B.n721 B.n720 585
R446 B.n720 B.n719 585
R447 B.n722 B.n367 585
R448 B.n367 B.n366 585
R449 B.n724 B.n723 585
R450 B.n725 B.n724 585
R451 B.n361 B.n360 585
R452 B.n362 B.n361 585
R453 B.n733 B.n732 585
R454 B.n732 B.n731 585
R455 B.n734 B.n359 585
R456 B.n359 B.n358 585
R457 B.n736 B.n735 585
R458 B.n737 B.n736 585
R459 B.n353 B.n352 585
R460 B.n354 B.n353 585
R461 B.n745 B.n744 585
R462 B.n744 B.n743 585
R463 B.n746 B.n351 585
R464 B.n351 B.n350 585
R465 B.n748 B.n747 585
R466 B.n749 B.n748 585
R467 B.n345 B.n344 585
R468 B.n346 B.n345 585
R469 B.n757 B.n756 585
R470 B.n756 B.n755 585
R471 B.n758 B.n343 585
R472 B.n343 B.n342 585
R473 B.n760 B.n759 585
R474 B.n761 B.n760 585
R475 B.n337 B.n336 585
R476 B.n338 B.n337 585
R477 B.n770 B.n769 585
R478 B.n769 B.n768 585
R479 B.n771 B.n335 585
R480 B.n335 B.n334 585
R481 B.n773 B.n772 585
R482 B.n774 B.n773 585
R483 B.n3 B.n0 585
R484 B.n4 B.n3 585
R485 B.n901 B.n1 585
R486 B.n902 B.n901 585
R487 B.n900 B.n899 585
R488 B.n900 B.n8 585
R489 B.n898 B.n9 585
R490 B.n12 B.n9 585
R491 B.n897 B.n896 585
R492 B.n896 B.n895 585
R493 B.n11 B.n10 585
R494 B.n894 B.n11 585
R495 B.n892 B.n891 585
R496 B.n893 B.n892 585
R497 B.n890 B.n17 585
R498 B.n17 B.n16 585
R499 B.n889 B.n888 585
R500 B.n888 B.n887 585
R501 B.n19 B.n18 585
R502 B.n886 B.n19 585
R503 B.n884 B.n883 585
R504 B.n885 B.n884 585
R505 B.n882 B.n24 585
R506 B.n24 B.n23 585
R507 B.n881 B.n880 585
R508 B.n880 B.n879 585
R509 B.n26 B.n25 585
R510 B.n878 B.n26 585
R511 B.n876 B.n875 585
R512 B.n877 B.n876 585
R513 B.n874 B.n31 585
R514 B.n31 B.n30 585
R515 B.n873 B.n872 585
R516 B.n872 B.n871 585
R517 B.n33 B.n32 585
R518 B.n870 B.n33 585
R519 B.n868 B.n867 585
R520 B.n869 B.n868 585
R521 B.n866 B.n38 585
R522 B.n38 B.n37 585
R523 B.n865 B.n864 585
R524 B.n864 B.n863 585
R525 B.n40 B.n39 585
R526 B.n862 B.n40 585
R527 B.n860 B.n859 585
R528 B.n861 B.n860 585
R529 B.n858 B.n45 585
R530 B.n45 B.n44 585
R531 B.n857 B.n856 585
R532 B.n856 B.n855 585
R533 B.n47 B.n46 585
R534 B.n854 B.n47 585
R535 B.n852 B.n851 585
R536 B.n853 B.n852 585
R537 B.n850 B.n52 585
R538 B.n52 B.n51 585
R539 B.n849 B.n848 585
R540 B.n848 B.n847 585
R541 B.n54 B.n53 585
R542 B.n846 B.n54 585
R543 B.n844 B.n843 585
R544 B.n845 B.n844 585
R545 B.n842 B.n59 585
R546 B.n59 B.n58 585
R547 B.n841 B.n840 585
R548 B.n840 B.n839 585
R549 B.n61 B.n60 585
R550 B.n838 B.n61 585
R551 B.n836 B.n835 585
R552 B.n837 B.n836 585
R553 B.n834 B.n66 585
R554 B.n66 B.n65 585
R555 B.n833 B.n832 585
R556 B.n832 B.n831 585
R557 B.n68 B.n67 585
R558 B.n830 B.n68 585
R559 B.n905 B.n904 585
R560 B.n903 B.n2 585
R561 B.n128 B.n68 482.89
R562 B.n828 B.n70 482.89
R563 B.n666 B.n403 482.89
R564 B.n662 B.n401 482.89
R565 B.n126 B.t8 319.837
R566 B.n123 B.t15 319.837
R567 B.n460 B.t4 319.837
R568 B.n457 B.t12 319.837
R569 B.n829 B.n121 256.663
R570 B.n829 B.n120 256.663
R571 B.n829 B.n119 256.663
R572 B.n829 B.n118 256.663
R573 B.n829 B.n117 256.663
R574 B.n829 B.n116 256.663
R575 B.n829 B.n115 256.663
R576 B.n829 B.n114 256.663
R577 B.n829 B.n113 256.663
R578 B.n829 B.n112 256.663
R579 B.n829 B.n111 256.663
R580 B.n829 B.n110 256.663
R581 B.n829 B.n109 256.663
R582 B.n829 B.n108 256.663
R583 B.n829 B.n107 256.663
R584 B.n829 B.n106 256.663
R585 B.n829 B.n105 256.663
R586 B.n829 B.n104 256.663
R587 B.n829 B.n103 256.663
R588 B.n829 B.n102 256.663
R589 B.n829 B.n101 256.663
R590 B.n829 B.n100 256.663
R591 B.n829 B.n99 256.663
R592 B.n829 B.n98 256.663
R593 B.n829 B.n97 256.663
R594 B.n829 B.n96 256.663
R595 B.n829 B.n95 256.663
R596 B.n829 B.n94 256.663
R597 B.n829 B.n93 256.663
R598 B.n829 B.n92 256.663
R599 B.n829 B.n91 256.663
R600 B.n829 B.n90 256.663
R601 B.n829 B.n89 256.663
R602 B.n829 B.n88 256.663
R603 B.n829 B.n87 256.663
R604 B.n829 B.n86 256.663
R605 B.n829 B.n85 256.663
R606 B.n829 B.n84 256.663
R607 B.n829 B.n83 256.663
R608 B.n829 B.n82 256.663
R609 B.n829 B.n81 256.663
R610 B.n829 B.n80 256.663
R611 B.n829 B.n79 256.663
R612 B.n829 B.n78 256.663
R613 B.n829 B.n77 256.663
R614 B.n829 B.n76 256.663
R615 B.n829 B.n75 256.663
R616 B.n829 B.n74 256.663
R617 B.n829 B.n73 256.663
R618 B.n829 B.n72 256.663
R619 B.n829 B.n71 256.663
R620 B.n664 B.n663 256.663
R621 B.n664 B.n406 256.663
R622 B.n664 B.n407 256.663
R623 B.n664 B.n408 256.663
R624 B.n664 B.n409 256.663
R625 B.n664 B.n410 256.663
R626 B.n664 B.n411 256.663
R627 B.n664 B.n412 256.663
R628 B.n664 B.n413 256.663
R629 B.n664 B.n414 256.663
R630 B.n664 B.n415 256.663
R631 B.n664 B.n416 256.663
R632 B.n664 B.n417 256.663
R633 B.n664 B.n418 256.663
R634 B.n664 B.n419 256.663
R635 B.n664 B.n420 256.663
R636 B.n664 B.n421 256.663
R637 B.n664 B.n422 256.663
R638 B.n664 B.n423 256.663
R639 B.n664 B.n424 256.663
R640 B.n664 B.n425 256.663
R641 B.n664 B.n426 256.663
R642 B.n664 B.n427 256.663
R643 B.n664 B.n428 256.663
R644 B.n664 B.n429 256.663
R645 B.n664 B.n430 256.663
R646 B.n664 B.n431 256.663
R647 B.n664 B.n432 256.663
R648 B.n664 B.n433 256.663
R649 B.n664 B.n434 256.663
R650 B.n664 B.n435 256.663
R651 B.n664 B.n436 256.663
R652 B.n664 B.n437 256.663
R653 B.n664 B.n438 256.663
R654 B.n664 B.n439 256.663
R655 B.n664 B.n440 256.663
R656 B.n664 B.n441 256.663
R657 B.n664 B.n442 256.663
R658 B.n664 B.n443 256.663
R659 B.n664 B.n444 256.663
R660 B.n664 B.n445 256.663
R661 B.n664 B.n446 256.663
R662 B.n664 B.n447 256.663
R663 B.n664 B.n448 256.663
R664 B.n664 B.n449 256.663
R665 B.n664 B.n450 256.663
R666 B.n664 B.n451 256.663
R667 B.n664 B.n452 256.663
R668 B.n664 B.n453 256.663
R669 B.n664 B.n454 256.663
R670 B.n665 B.n664 256.663
R671 B.n907 B.n906 256.663
R672 B.n132 B.n131 163.367
R673 B.n136 B.n135 163.367
R674 B.n140 B.n139 163.367
R675 B.n144 B.n143 163.367
R676 B.n148 B.n147 163.367
R677 B.n152 B.n151 163.367
R678 B.n156 B.n155 163.367
R679 B.n160 B.n159 163.367
R680 B.n164 B.n163 163.367
R681 B.n168 B.n167 163.367
R682 B.n172 B.n171 163.367
R683 B.n176 B.n175 163.367
R684 B.n180 B.n179 163.367
R685 B.n184 B.n183 163.367
R686 B.n188 B.n187 163.367
R687 B.n192 B.n191 163.367
R688 B.n196 B.n195 163.367
R689 B.n200 B.n199 163.367
R690 B.n204 B.n203 163.367
R691 B.n208 B.n207 163.367
R692 B.n212 B.n211 163.367
R693 B.n216 B.n215 163.367
R694 B.n220 B.n219 163.367
R695 B.n225 B.n224 163.367
R696 B.n229 B.n228 163.367
R697 B.n233 B.n232 163.367
R698 B.n237 B.n236 163.367
R699 B.n241 B.n240 163.367
R700 B.n245 B.n244 163.367
R701 B.n249 B.n248 163.367
R702 B.n253 B.n252 163.367
R703 B.n257 B.n256 163.367
R704 B.n261 B.n260 163.367
R705 B.n265 B.n264 163.367
R706 B.n269 B.n268 163.367
R707 B.n273 B.n272 163.367
R708 B.n277 B.n276 163.367
R709 B.n281 B.n280 163.367
R710 B.n285 B.n284 163.367
R711 B.n289 B.n288 163.367
R712 B.n293 B.n292 163.367
R713 B.n297 B.n296 163.367
R714 B.n301 B.n300 163.367
R715 B.n305 B.n304 163.367
R716 B.n309 B.n308 163.367
R717 B.n313 B.n312 163.367
R718 B.n317 B.n316 163.367
R719 B.n321 B.n320 163.367
R720 B.n325 B.n324 163.367
R721 B.n329 B.n328 163.367
R722 B.n828 B.n122 163.367
R723 B.n670 B.n403 163.367
R724 B.n670 B.n397 163.367
R725 B.n678 B.n397 163.367
R726 B.n678 B.n395 163.367
R727 B.n682 B.n395 163.367
R728 B.n682 B.n388 163.367
R729 B.n690 B.n388 163.367
R730 B.n690 B.n386 163.367
R731 B.n694 B.n386 163.367
R732 B.n694 B.n381 163.367
R733 B.n702 B.n381 163.367
R734 B.n702 B.n379 163.367
R735 B.n706 B.n379 163.367
R736 B.n706 B.n373 163.367
R737 B.n714 B.n373 163.367
R738 B.n714 B.n371 163.367
R739 B.n718 B.n371 163.367
R740 B.n718 B.n365 163.367
R741 B.n726 B.n365 163.367
R742 B.n726 B.n363 163.367
R743 B.n730 B.n363 163.367
R744 B.n730 B.n357 163.367
R745 B.n738 B.n357 163.367
R746 B.n738 B.n355 163.367
R747 B.n742 B.n355 163.367
R748 B.n742 B.n349 163.367
R749 B.n750 B.n349 163.367
R750 B.n750 B.n347 163.367
R751 B.n754 B.n347 163.367
R752 B.n754 B.n341 163.367
R753 B.n762 B.n341 163.367
R754 B.n762 B.n339 163.367
R755 B.n767 B.n339 163.367
R756 B.n767 B.n333 163.367
R757 B.n775 B.n333 163.367
R758 B.n776 B.n775 163.367
R759 B.n776 B.n5 163.367
R760 B.n6 B.n5 163.367
R761 B.n7 B.n6 163.367
R762 B.n782 B.n7 163.367
R763 B.n783 B.n782 163.367
R764 B.n783 B.n13 163.367
R765 B.n14 B.n13 163.367
R766 B.n15 B.n14 163.367
R767 B.n788 B.n15 163.367
R768 B.n788 B.n20 163.367
R769 B.n21 B.n20 163.367
R770 B.n22 B.n21 163.367
R771 B.n793 B.n22 163.367
R772 B.n793 B.n27 163.367
R773 B.n28 B.n27 163.367
R774 B.n29 B.n28 163.367
R775 B.n798 B.n29 163.367
R776 B.n798 B.n34 163.367
R777 B.n35 B.n34 163.367
R778 B.n36 B.n35 163.367
R779 B.n803 B.n36 163.367
R780 B.n803 B.n41 163.367
R781 B.n42 B.n41 163.367
R782 B.n43 B.n42 163.367
R783 B.n808 B.n43 163.367
R784 B.n808 B.n48 163.367
R785 B.n49 B.n48 163.367
R786 B.n50 B.n49 163.367
R787 B.n813 B.n50 163.367
R788 B.n813 B.n55 163.367
R789 B.n56 B.n55 163.367
R790 B.n57 B.n56 163.367
R791 B.n818 B.n57 163.367
R792 B.n818 B.n62 163.367
R793 B.n63 B.n62 163.367
R794 B.n64 B.n63 163.367
R795 B.n823 B.n64 163.367
R796 B.n823 B.n69 163.367
R797 B.n70 B.n69 163.367
R798 B.n456 B.n455 163.367
R799 B.n657 B.n455 163.367
R800 B.n655 B.n654 163.367
R801 B.n651 B.n650 163.367
R802 B.n647 B.n646 163.367
R803 B.n643 B.n642 163.367
R804 B.n639 B.n638 163.367
R805 B.n635 B.n634 163.367
R806 B.n631 B.n630 163.367
R807 B.n627 B.n626 163.367
R808 B.n623 B.n622 163.367
R809 B.n619 B.n618 163.367
R810 B.n615 B.n614 163.367
R811 B.n611 B.n610 163.367
R812 B.n607 B.n606 163.367
R813 B.n603 B.n602 163.367
R814 B.n599 B.n598 163.367
R815 B.n595 B.n594 163.367
R816 B.n591 B.n590 163.367
R817 B.n587 B.n586 163.367
R818 B.n583 B.n582 163.367
R819 B.n579 B.n578 163.367
R820 B.n575 B.n574 163.367
R821 B.n571 B.n570 163.367
R822 B.n567 B.n566 163.367
R823 B.n563 B.n562 163.367
R824 B.n559 B.n558 163.367
R825 B.n555 B.n554 163.367
R826 B.n550 B.n549 163.367
R827 B.n546 B.n545 163.367
R828 B.n542 B.n541 163.367
R829 B.n538 B.n537 163.367
R830 B.n534 B.n533 163.367
R831 B.n530 B.n529 163.367
R832 B.n526 B.n525 163.367
R833 B.n522 B.n521 163.367
R834 B.n518 B.n517 163.367
R835 B.n514 B.n513 163.367
R836 B.n510 B.n509 163.367
R837 B.n506 B.n505 163.367
R838 B.n502 B.n501 163.367
R839 B.n498 B.n497 163.367
R840 B.n494 B.n493 163.367
R841 B.n490 B.n489 163.367
R842 B.n486 B.n485 163.367
R843 B.n482 B.n481 163.367
R844 B.n478 B.n477 163.367
R845 B.n474 B.n473 163.367
R846 B.n470 B.n469 163.367
R847 B.n466 B.n465 163.367
R848 B.n462 B.n405 163.367
R849 B.n672 B.n401 163.367
R850 B.n672 B.n399 163.367
R851 B.n676 B.n399 163.367
R852 B.n676 B.n393 163.367
R853 B.n684 B.n393 163.367
R854 B.n684 B.n391 163.367
R855 B.n688 B.n391 163.367
R856 B.n688 B.n385 163.367
R857 B.n696 B.n385 163.367
R858 B.n696 B.n383 163.367
R859 B.n700 B.n383 163.367
R860 B.n700 B.n377 163.367
R861 B.n708 B.n377 163.367
R862 B.n708 B.n375 163.367
R863 B.n712 B.n375 163.367
R864 B.n712 B.n369 163.367
R865 B.n720 B.n369 163.367
R866 B.n720 B.n367 163.367
R867 B.n724 B.n367 163.367
R868 B.n724 B.n361 163.367
R869 B.n732 B.n361 163.367
R870 B.n732 B.n359 163.367
R871 B.n736 B.n359 163.367
R872 B.n736 B.n353 163.367
R873 B.n744 B.n353 163.367
R874 B.n744 B.n351 163.367
R875 B.n748 B.n351 163.367
R876 B.n748 B.n345 163.367
R877 B.n756 B.n345 163.367
R878 B.n756 B.n343 163.367
R879 B.n760 B.n343 163.367
R880 B.n760 B.n337 163.367
R881 B.n769 B.n337 163.367
R882 B.n769 B.n335 163.367
R883 B.n773 B.n335 163.367
R884 B.n773 B.n3 163.367
R885 B.n905 B.n3 163.367
R886 B.n901 B.n2 163.367
R887 B.n901 B.n900 163.367
R888 B.n900 B.n9 163.367
R889 B.n896 B.n9 163.367
R890 B.n896 B.n11 163.367
R891 B.n892 B.n11 163.367
R892 B.n892 B.n17 163.367
R893 B.n888 B.n17 163.367
R894 B.n888 B.n19 163.367
R895 B.n884 B.n19 163.367
R896 B.n884 B.n24 163.367
R897 B.n880 B.n24 163.367
R898 B.n880 B.n26 163.367
R899 B.n876 B.n26 163.367
R900 B.n876 B.n31 163.367
R901 B.n872 B.n31 163.367
R902 B.n872 B.n33 163.367
R903 B.n868 B.n33 163.367
R904 B.n868 B.n38 163.367
R905 B.n864 B.n38 163.367
R906 B.n864 B.n40 163.367
R907 B.n860 B.n40 163.367
R908 B.n860 B.n45 163.367
R909 B.n856 B.n45 163.367
R910 B.n856 B.n47 163.367
R911 B.n852 B.n47 163.367
R912 B.n852 B.n52 163.367
R913 B.n848 B.n52 163.367
R914 B.n848 B.n54 163.367
R915 B.n844 B.n54 163.367
R916 B.n844 B.n59 163.367
R917 B.n840 B.n59 163.367
R918 B.n840 B.n61 163.367
R919 B.n836 B.n61 163.367
R920 B.n836 B.n66 163.367
R921 B.n832 B.n66 163.367
R922 B.n832 B.n68 163.367
R923 B.n123 B.t16 134.879
R924 B.n460 B.t7 134.879
R925 B.n126 B.t10 134.861
R926 B.n457 B.t14 134.861
R927 B.n128 B.n71 71.676
R928 B.n132 B.n72 71.676
R929 B.n136 B.n73 71.676
R930 B.n140 B.n74 71.676
R931 B.n144 B.n75 71.676
R932 B.n148 B.n76 71.676
R933 B.n152 B.n77 71.676
R934 B.n156 B.n78 71.676
R935 B.n160 B.n79 71.676
R936 B.n164 B.n80 71.676
R937 B.n168 B.n81 71.676
R938 B.n172 B.n82 71.676
R939 B.n176 B.n83 71.676
R940 B.n180 B.n84 71.676
R941 B.n184 B.n85 71.676
R942 B.n188 B.n86 71.676
R943 B.n192 B.n87 71.676
R944 B.n196 B.n88 71.676
R945 B.n200 B.n89 71.676
R946 B.n204 B.n90 71.676
R947 B.n208 B.n91 71.676
R948 B.n212 B.n92 71.676
R949 B.n216 B.n93 71.676
R950 B.n220 B.n94 71.676
R951 B.n225 B.n95 71.676
R952 B.n229 B.n96 71.676
R953 B.n233 B.n97 71.676
R954 B.n237 B.n98 71.676
R955 B.n241 B.n99 71.676
R956 B.n245 B.n100 71.676
R957 B.n249 B.n101 71.676
R958 B.n253 B.n102 71.676
R959 B.n257 B.n103 71.676
R960 B.n261 B.n104 71.676
R961 B.n265 B.n105 71.676
R962 B.n269 B.n106 71.676
R963 B.n273 B.n107 71.676
R964 B.n277 B.n108 71.676
R965 B.n281 B.n109 71.676
R966 B.n285 B.n110 71.676
R967 B.n289 B.n111 71.676
R968 B.n293 B.n112 71.676
R969 B.n297 B.n113 71.676
R970 B.n301 B.n114 71.676
R971 B.n305 B.n115 71.676
R972 B.n309 B.n116 71.676
R973 B.n313 B.n117 71.676
R974 B.n317 B.n118 71.676
R975 B.n321 B.n119 71.676
R976 B.n325 B.n120 71.676
R977 B.n329 B.n121 71.676
R978 B.n122 B.n121 71.676
R979 B.n328 B.n120 71.676
R980 B.n324 B.n119 71.676
R981 B.n320 B.n118 71.676
R982 B.n316 B.n117 71.676
R983 B.n312 B.n116 71.676
R984 B.n308 B.n115 71.676
R985 B.n304 B.n114 71.676
R986 B.n300 B.n113 71.676
R987 B.n296 B.n112 71.676
R988 B.n292 B.n111 71.676
R989 B.n288 B.n110 71.676
R990 B.n284 B.n109 71.676
R991 B.n280 B.n108 71.676
R992 B.n276 B.n107 71.676
R993 B.n272 B.n106 71.676
R994 B.n268 B.n105 71.676
R995 B.n264 B.n104 71.676
R996 B.n260 B.n103 71.676
R997 B.n256 B.n102 71.676
R998 B.n252 B.n101 71.676
R999 B.n248 B.n100 71.676
R1000 B.n244 B.n99 71.676
R1001 B.n240 B.n98 71.676
R1002 B.n236 B.n97 71.676
R1003 B.n232 B.n96 71.676
R1004 B.n228 B.n95 71.676
R1005 B.n224 B.n94 71.676
R1006 B.n219 B.n93 71.676
R1007 B.n215 B.n92 71.676
R1008 B.n211 B.n91 71.676
R1009 B.n207 B.n90 71.676
R1010 B.n203 B.n89 71.676
R1011 B.n199 B.n88 71.676
R1012 B.n195 B.n87 71.676
R1013 B.n191 B.n86 71.676
R1014 B.n187 B.n85 71.676
R1015 B.n183 B.n84 71.676
R1016 B.n179 B.n83 71.676
R1017 B.n175 B.n82 71.676
R1018 B.n171 B.n81 71.676
R1019 B.n167 B.n80 71.676
R1020 B.n163 B.n79 71.676
R1021 B.n159 B.n78 71.676
R1022 B.n155 B.n77 71.676
R1023 B.n151 B.n76 71.676
R1024 B.n147 B.n75 71.676
R1025 B.n143 B.n74 71.676
R1026 B.n139 B.n73 71.676
R1027 B.n135 B.n72 71.676
R1028 B.n131 B.n71 71.676
R1029 B.n663 B.n662 71.676
R1030 B.n657 B.n406 71.676
R1031 B.n654 B.n407 71.676
R1032 B.n650 B.n408 71.676
R1033 B.n646 B.n409 71.676
R1034 B.n642 B.n410 71.676
R1035 B.n638 B.n411 71.676
R1036 B.n634 B.n412 71.676
R1037 B.n630 B.n413 71.676
R1038 B.n626 B.n414 71.676
R1039 B.n622 B.n415 71.676
R1040 B.n618 B.n416 71.676
R1041 B.n614 B.n417 71.676
R1042 B.n610 B.n418 71.676
R1043 B.n606 B.n419 71.676
R1044 B.n602 B.n420 71.676
R1045 B.n598 B.n421 71.676
R1046 B.n594 B.n422 71.676
R1047 B.n590 B.n423 71.676
R1048 B.n586 B.n424 71.676
R1049 B.n582 B.n425 71.676
R1050 B.n578 B.n426 71.676
R1051 B.n574 B.n427 71.676
R1052 B.n570 B.n428 71.676
R1053 B.n566 B.n429 71.676
R1054 B.n562 B.n430 71.676
R1055 B.n558 B.n431 71.676
R1056 B.n554 B.n432 71.676
R1057 B.n549 B.n433 71.676
R1058 B.n545 B.n434 71.676
R1059 B.n541 B.n435 71.676
R1060 B.n537 B.n436 71.676
R1061 B.n533 B.n437 71.676
R1062 B.n529 B.n438 71.676
R1063 B.n525 B.n439 71.676
R1064 B.n521 B.n440 71.676
R1065 B.n517 B.n441 71.676
R1066 B.n513 B.n442 71.676
R1067 B.n509 B.n443 71.676
R1068 B.n505 B.n444 71.676
R1069 B.n501 B.n445 71.676
R1070 B.n497 B.n446 71.676
R1071 B.n493 B.n447 71.676
R1072 B.n489 B.n448 71.676
R1073 B.n485 B.n449 71.676
R1074 B.n481 B.n450 71.676
R1075 B.n477 B.n451 71.676
R1076 B.n473 B.n452 71.676
R1077 B.n469 B.n453 71.676
R1078 B.n465 B.n454 71.676
R1079 B.n665 B.n405 71.676
R1080 B.n663 B.n456 71.676
R1081 B.n655 B.n406 71.676
R1082 B.n651 B.n407 71.676
R1083 B.n647 B.n408 71.676
R1084 B.n643 B.n409 71.676
R1085 B.n639 B.n410 71.676
R1086 B.n635 B.n411 71.676
R1087 B.n631 B.n412 71.676
R1088 B.n627 B.n413 71.676
R1089 B.n623 B.n414 71.676
R1090 B.n619 B.n415 71.676
R1091 B.n615 B.n416 71.676
R1092 B.n611 B.n417 71.676
R1093 B.n607 B.n418 71.676
R1094 B.n603 B.n419 71.676
R1095 B.n599 B.n420 71.676
R1096 B.n595 B.n421 71.676
R1097 B.n591 B.n422 71.676
R1098 B.n587 B.n423 71.676
R1099 B.n583 B.n424 71.676
R1100 B.n579 B.n425 71.676
R1101 B.n575 B.n426 71.676
R1102 B.n571 B.n427 71.676
R1103 B.n567 B.n428 71.676
R1104 B.n563 B.n429 71.676
R1105 B.n559 B.n430 71.676
R1106 B.n555 B.n431 71.676
R1107 B.n550 B.n432 71.676
R1108 B.n546 B.n433 71.676
R1109 B.n542 B.n434 71.676
R1110 B.n538 B.n435 71.676
R1111 B.n534 B.n436 71.676
R1112 B.n530 B.n437 71.676
R1113 B.n526 B.n438 71.676
R1114 B.n522 B.n439 71.676
R1115 B.n518 B.n440 71.676
R1116 B.n514 B.n441 71.676
R1117 B.n510 B.n442 71.676
R1118 B.n506 B.n443 71.676
R1119 B.n502 B.n444 71.676
R1120 B.n498 B.n445 71.676
R1121 B.n494 B.n446 71.676
R1122 B.n490 B.n447 71.676
R1123 B.n486 B.n448 71.676
R1124 B.n482 B.n449 71.676
R1125 B.n478 B.n450 71.676
R1126 B.n474 B.n451 71.676
R1127 B.n470 B.n452 71.676
R1128 B.n466 B.n453 71.676
R1129 B.n462 B.n454 71.676
R1130 B.n666 B.n665 71.676
R1131 B.n906 B.n905 71.676
R1132 B.n906 B.n2 71.676
R1133 B.n124 B.t17 70.6844
R1134 B.n461 B.t6 70.6844
R1135 B.n127 B.t11 70.6666
R1136 B.n458 B.t13 70.6666
R1137 B.n127 B.n126 64.1944
R1138 B.n124 B.n123 64.1944
R1139 B.n461 B.n460 64.1944
R1140 B.n458 B.n457 64.1944
R1141 B.n664 B.n402 64.1455
R1142 B.n830 B.n829 64.1455
R1143 B.n222 B.n127 59.5399
R1144 B.n125 B.n124 59.5399
R1145 B.n552 B.n461 59.5399
R1146 B.n459 B.n458 59.5399
R1147 B.n671 B.n402 39.2965
R1148 B.n671 B.n398 39.2965
R1149 B.n677 B.n398 39.2965
R1150 B.n677 B.n394 39.2965
R1151 B.n683 B.n394 39.2965
R1152 B.n683 B.n389 39.2965
R1153 B.n689 B.n389 39.2965
R1154 B.n689 B.n390 39.2965
R1155 B.n695 B.n382 39.2965
R1156 B.n701 B.n382 39.2965
R1157 B.n701 B.n378 39.2965
R1158 B.n707 B.n378 39.2965
R1159 B.n707 B.n374 39.2965
R1160 B.n713 B.n374 39.2965
R1161 B.n713 B.n370 39.2965
R1162 B.n719 B.n370 39.2965
R1163 B.n719 B.n366 39.2965
R1164 B.n725 B.n366 39.2965
R1165 B.n725 B.n362 39.2965
R1166 B.n731 B.n362 39.2965
R1167 B.n737 B.n358 39.2965
R1168 B.n737 B.n354 39.2965
R1169 B.n743 B.n354 39.2965
R1170 B.n743 B.n350 39.2965
R1171 B.n749 B.n350 39.2965
R1172 B.n749 B.n346 39.2965
R1173 B.n755 B.n346 39.2965
R1174 B.n755 B.n342 39.2965
R1175 B.n761 B.n342 39.2965
R1176 B.n768 B.n338 39.2965
R1177 B.n768 B.n334 39.2965
R1178 B.n774 B.n334 39.2965
R1179 B.n774 B.n4 39.2965
R1180 B.n904 B.n4 39.2965
R1181 B.n904 B.n903 39.2965
R1182 B.n903 B.n902 39.2965
R1183 B.n902 B.n8 39.2965
R1184 B.n12 B.n8 39.2965
R1185 B.n895 B.n12 39.2965
R1186 B.n895 B.n894 39.2965
R1187 B.n893 B.n16 39.2965
R1188 B.n887 B.n16 39.2965
R1189 B.n887 B.n886 39.2965
R1190 B.n886 B.n885 39.2965
R1191 B.n885 B.n23 39.2965
R1192 B.n879 B.n23 39.2965
R1193 B.n879 B.n878 39.2965
R1194 B.n878 B.n877 39.2965
R1195 B.n877 B.n30 39.2965
R1196 B.n871 B.n870 39.2965
R1197 B.n870 B.n869 39.2965
R1198 B.n869 B.n37 39.2965
R1199 B.n863 B.n37 39.2965
R1200 B.n863 B.n862 39.2965
R1201 B.n862 B.n861 39.2965
R1202 B.n861 B.n44 39.2965
R1203 B.n855 B.n44 39.2965
R1204 B.n855 B.n854 39.2965
R1205 B.n854 B.n853 39.2965
R1206 B.n853 B.n51 39.2965
R1207 B.n847 B.n51 39.2965
R1208 B.n846 B.n845 39.2965
R1209 B.n845 B.n58 39.2965
R1210 B.n839 B.n58 39.2965
R1211 B.n839 B.n838 39.2965
R1212 B.n838 B.n837 39.2965
R1213 B.n837 B.n65 39.2965
R1214 B.n831 B.n65 39.2965
R1215 B.n831 B.n830 39.2965
R1216 B.t1 B.n338 38.1408
R1217 B.n894 B.t3 38.1408
R1218 B.n661 B.n400 31.3761
R1219 B.n668 B.n667 31.3761
R1220 B.n827 B.n826 31.3761
R1221 B.n129 B.n67 31.3761
R1222 B.t0 B.n358 27.7389
R1223 B.t2 B.n30 27.7389
R1224 B.n695 B.t5 25.4273
R1225 B.n847 B.t9 25.4273
R1226 B B.n907 18.0485
R1227 B.n390 B.t5 13.8697
R1228 B.t9 B.n846 13.8697
R1229 B.n731 B.t0 11.5582
R1230 B.n871 B.t2 11.5582
R1231 B.n673 B.n400 10.6151
R1232 B.n674 B.n673 10.6151
R1233 B.n675 B.n674 10.6151
R1234 B.n675 B.n392 10.6151
R1235 B.n685 B.n392 10.6151
R1236 B.n686 B.n685 10.6151
R1237 B.n687 B.n686 10.6151
R1238 B.n687 B.n384 10.6151
R1239 B.n697 B.n384 10.6151
R1240 B.n698 B.n697 10.6151
R1241 B.n699 B.n698 10.6151
R1242 B.n699 B.n376 10.6151
R1243 B.n709 B.n376 10.6151
R1244 B.n710 B.n709 10.6151
R1245 B.n711 B.n710 10.6151
R1246 B.n711 B.n368 10.6151
R1247 B.n721 B.n368 10.6151
R1248 B.n722 B.n721 10.6151
R1249 B.n723 B.n722 10.6151
R1250 B.n723 B.n360 10.6151
R1251 B.n733 B.n360 10.6151
R1252 B.n734 B.n733 10.6151
R1253 B.n735 B.n734 10.6151
R1254 B.n735 B.n352 10.6151
R1255 B.n745 B.n352 10.6151
R1256 B.n746 B.n745 10.6151
R1257 B.n747 B.n746 10.6151
R1258 B.n747 B.n344 10.6151
R1259 B.n757 B.n344 10.6151
R1260 B.n758 B.n757 10.6151
R1261 B.n759 B.n758 10.6151
R1262 B.n759 B.n336 10.6151
R1263 B.n770 B.n336 10.6151
R1264 B.n771 B.n770 10.6151
R1265 B.n772 B.n771 10.6151
R1266 B.n772 B.n0 10.6151
R1267 B.n661 B.n660 10.6151
R1268 B.n660 B.n659 10.6151
R1269 B.n659 B.n658 10.6151
R1270 B.n658 B.n656 10.6151
R1271 B.n656 B.n653 10.6151
R1272 B.n653 B.n652 10.6151
R1273 B.n652 B.n649 10.6151
R1274 B.n649 B.n648 10.6151
R1275 B.n648 B.n645 10.6151
R1276 B.n645 B.n644 10.6151
R1277 B.n644 B.n641 10.6151
R1278 B.n641 B.n640 10.6151
R1279 B.n640 B.n637 10.6151
R1280 B.n637 B.n636 10.6151
R1281 B.n636 B.n633 10.6151
R1282 B.n633 B.n632 10.6151
R1283 B.n632 B.n629 10.6151
R1284 B.n629 B.n628 10.6151
R1285 B.n628 B.n625 10.6151
R1286 B.n625 B.n624 10.6151
R1287 B.n624 B.n621 10.6151
R1288 B.n621 B.n620 10.6151
R1289 B.n620 B.n617 10.6151
R1290 B.n617 B.n616 10.6151
R1291 B.n616 B.n613 10.6151
R1292 B.n613 B.n612 10.6151
R1293 B.n612 B.n609 10.6151
R1294 B.n609 B.n608 10.6151
R1295 B.n608 B.n605 10.6151
R1296 B.n605 B.n604 10.6151
R1297 B.n604 B.n601 10.6151
R1298 B.n601 B.n600 10.6151
R1299 B.n600 B.n597 10.6151
R1300 B.n597 B.n596 10.6151
R1301 B.n596 B.n593 10.6151
R1302 B.n593 B.n592 10.6151
R1303 B.n592 B.n589 10.6151
R1304 B.n589 B.n588 10.6151
R1305 B.n588 B.n585 10.6151
R1306 B.n585 B.n584 10.6151
R1307 B.n584 B.n581 10.6151
R1308 B.n581 B.n580 10.6151
R1309 B.n580 B.n577 10.6151
R1310 B.n577 B.n576 10.6151
R1311 B.n576 B.n573 10.6151
R1312 B.n573 B.n572 10.6151
R1313 B.n569 B.n568 10.6151
R1314 B.n568 B.n565 10.6151
R1315 B.n565 B.n564 10.6151
R1316 B.n564 B.n561 10.6151
R1317 B.n561 B.n560 10.6151
R1318 B.n560 B.n557 10.6151
R1319 B.n557 B.n556 10.6151
R1320 B.n556 B.n553 10.6151
R1321 B.n551 B.n548 10.6151
R1322 B.n548 B.n547 10.6151
R1323 B.n547 B.n544 10.6151
R1324 B.n544 B.n543 10.6151
R1325 B.n543 B.n540 10.6151
R1326 B.n540 B.n539 10.6151
R1327 B.n539 B.n536 10.6151
R1328 B.n536 B.n535 10.6151
R1329 B.n535 B.n532 10.6151
R1330 B.n532 B.n531 10.6151
R1331 B.n531 B.n528 10.6151
R1332 B.n528 B.n527 10.6151
R1333 B.n527 B.n524 10.6151
R1334 B.n524 B.n523 10.6151
R1335 B.n523 B.n520 10.6151
R1336 B.n520 B.n519 10.6151
R1337 B.n519 B.n516 10.6151
R1338 B.n516 B.n515 10.6151
R1339 B.n515 B.n512 10.6151
R1340 B.n512 B.n511 10.6151
R1341 B.n511 B.n508 10.6151
R1342 B.n508 B.n507 10.6151
R1343 B.n507 B.n504 10.6151
R1344 B.n504 B.n503 10.6151
R1345 B.n503 B.n500 10.6151
R1346 B.n500 B.n499 10.6151
R1347 B.n499 B.n496 10.6151
R1348 B.n496 B.n495 10.6151
R1349 B.n495 B.n492 10.6151
R1350 B.n492 B.n491 10.6151
R1351 B.n491 B.n488 10.6151
R1352 B.n488 B.n487 10.6151
R1353 B.n487 B.n484 10.6151
R1354 B.n484 B.n483 10.6151
R1355 B.n483 B.n480 10.6151
R1356 B.n480 B.n479 10.6151
R1357 B.n479 B.n476 10.6151
R1358 B.n476 B.n475 10.6151
R1359 B.n475 B.n472 10.6151
R1360 B.n472 B.n471 10.6151
R1361 B.n471 B.n468 10.6151
R1362 B.n468 B.n467 10.6151
R1363 B.n467 B.n464 10.6151
R1364 B.n464 B.n463 10.6151
R1365 B.n463 B.n404 10.6151
R1366 B.n667 B.n404 10.6151
R1367 B.n669 B.n668 10.6151
R1368 B.n669 B.n396 10.6151
R1369 B.n679 B.n396 10.6151
R1370 B.n680 B.n679 10.6151
R1371 B.n681 B.n680 10.6151
R1372 B.n681 B.n387 10.6151
R1373 B.n691 B.n387 10.6151
R1374 B.n692 B.n691 10.6151
R1375 B.n693 B.n692 10.6151
R1376 B.n693 B.n380 10.6151
R1377 B.n703 B.n380 10.6151
R1378 B.n704 B.n703 10.6151
R1379 B.n705 B.n704 10.6151
R1380 B.n705 B.n372 10.6151
R1381 B.n715 B.n372 10.6151
R1382 B.n716 B.n715 10.6151
R1383 B.n717 B.n716 10.6151
R1384 B.n717 B.n364 10.6151
R1385 B.n727 B.n364 10.6151
R1386 B.n728 B.n727 10.6151
R1387 B.n729 B.n728 10.6151
R1388 B.n729 B.n356 10.6151
R1389 B.n739 B.n356 10.6151
R1390 B.n740 B.n739 10.6151
R1391 B.n741 B.n740 10.6151
R1392 B.n741 B.n348 10.6151
R1393 B.n751 B.n348 10.6151
R1394 B.n752 B.n751 10.6151
R1395 B.n753 B.n752 10.6151
R1396 B.n753 B.n340 10.6151
R1397 B.n763 B.n340 10.6151
R1398 B.n764 B.n763 10.6151
R1399 B.n766 B.n764 10.6151
R1400 B.n766 B.n765 10.6151
R1401 B.n765 B.n332 10.6151
R1402 B.n777 B.n332 10.6151
R1403 B.n778 B.n777 10.6151
R1404 B.n779 B.n778 10.6151
R1405 B.n780 B.n779 10.6151
R1406 B.n781 B.n780 10.6151
R1407 B.n784 B.n781 10.6151
R1408 B.n785 B.n784 10.6151
R1409 B.n786 B.n785 10.6151
R1410 B.n787 B.n786 10.6151
R1411 B.n789 B.n787 10.6151
R1412 B.n790 B.n789 10.6151
R1413 B.n791 B.n790 10.6151
R1414 B.n792 B.n791 10.6151
R1415 B.n794 B.n792 10.6151
R1416 B.n795 B.n794 10.6151
R1417 B.n796 B.n795 10.6151
R1418 B.n797 B.n796 10.6151
R1419 B.n799 B.n797 10.6151
R1420 B.n800 B.n799 10.6151
R1421 B.n801 B.n800 10.6151
R1422 B.n802 B.n801 10.6151
R1423 B.n804 B.n802 10.6151
R1424 B.n805 B.n804 10.6151
R1425 B.n806 B.n805 10.6151
R1426 B.n807 B.n806 10.6151
R1427 B.n809 B.n807 10.6151
R1428 B.n810 B.n809 10.6151
R1429 B.n811 B.n810 10.6151
R1430 B.n812 B.n811 10.6151
R1431 B.n814 B.n812 10.6151
R1432 B.n815 B.n814 10.6151
R1433 B.n816 B.n815 10.6151
R1434 B.n817 B.n816 10.6151
R1435 B.n819 B.n817 10.6151
R1436 B.n820 B.n819 10.6151
R1437 B.n821 B.n820 10.6151
R1438 B.n822 B.n821 10.6151
R1439 B.n824 B.n822 10.6151
R1440 B.n825 B.n824 10.6151
R1441 B.n826 B.n825 10.6151
R1442 B.n899 B.n1 10.6151
R1443 B.n899 B.n898 10.6151
R1444 B.n898 B.n897 10.6151
R1445 B.n897 B.n10 10.6151
R1446 B.n891 B.n10 10.6151
R1447 B.n891 B.n890 10.6151
R1448 B.n890 B.n889 10.6151
R1449 B.n889 B.n18 10.6151
R1450 B.n883 B.n18 10.6151
R1451 B.n883 B.n882 10.6151
R1452 B.n882 B.n881 10.6151
R1453 B.n881 B.n25 10.6151
R1454 B.n875 B.n25 10.6151
R1455 B.n875 B.n874 10.6151
R1456 B.n874 B.n873 10.6151
R1457 B.n873 B.n32 10.6151
R1458 B.n867 B.n32 10.6151
R1459 B.n867 B.n866 10.6151
R1460 B.n866 B.n865 10.6151
R1461 B.n865 B.n39 10.6151
R1462 B.n859 B.n39 10.6151
R1463 B.n859 B.n858 10.6151
R1464 B.n858 B.n857 10.6151
R1465 B.n857 B.n46 10.6151
R1466 B.n851 B.n46 10.6151
R1467 B.n851 B.n850 10.6151
R1468 B.n850 B.n849 10.6151
R1469 B.n849 B.n53 10.6151
R1470 B.n843 B.n53 10.6151
R1471 B.n843 B.n842 10.6151
R1472 B.n842 B.n841 10.6151
R1473 B.n841 B.n60 10.6151
R1474 B.n835 B.n60 10.6151
R1475 B.n835 B.n834 10.6151
R1476 B.n834 B.n833 10.6151
R1477 B.n833 B.n67 10.6151
R1478 B.n130 B.n129 10.6151
R1479 B.n133 B.n130 10.6151
R1480 B.n134 B.n133 10.6151
R1481 B.n137 B.n134 10.6151
R1482 B.n138 B.n137 10.6151
R1483 B.n141 B.n138 10.6151
R1484 B.n142 B.n141 10.6151
R1485 B.n145 B.n142 10.6151
R1486 B.n146 B.n145 10.6151
R1487 B.n149 B.n146 10.6151
R1488 B.n150 B.n149 10.6151
R1489 B.n153 B.n150 10.6151
R1490 B.n154 B.n153 10.6151
R1491 B.n157 B.n154 10.6151
R1492 B.n158 B.n157 10.6151
R1493 B.n161 B.n158 10.6151
R1494 B.n162 B.n161 10.6151
R1495 B.n165 B.n162 10.6151
R1496 B.n166 B.n165 10.6151
R1497 B.n169 B.n166 10.6151
R1498 B.n170 B.n169 10.6151
R1499 B.n173 B.n170 10.6151
R1500 B.n174 B.n173 10.6151
R1501 B.n177 B.n174 10.6151
R1502 B.n178 B.n177 10.6151
R1503 B.n181 B.n178 10.6151
R1504 B.n182 B.n181 10.6151
R1505 B.n185 B.n182 10.6151
R1506 B.n186 B.n185 10.6151
R1507 B.n189 B.n186 10.6151
R1508 B.n190 B.n189 10.6151
R1509 B.n193 B.n190 10.6151
R1510 B.n194 B.n193 10.6151
R1511 B.n197 B.n194 10.6151
R1512 B.n198 B.n197 10.6151
R1513 B.n201 B.n198 10.6151
R1514 B.n202 B.n201 10.6151
R1515 B.n205 B.n202 10.6151
R1516 B.n206 B.n205 10.6151
R1517 B.n209 B.n206 10.6151
R1518 B.n210 B.n209 10.6151
R1519 B.n213 B.n210 10.6151
R1520 B.n214 B.n213 10.6151
R1521 B.n217 B.n214 10.6151
R1522 B.n218 B.n217 10.6151
R1523 B.n221 B.n218 10.6151
R1524 B.n226 B.n223 10.6151
R1525 B.n227 B.n226 10.6151
R1526 B.n230 B.n227 10.6151
R1527 B.n231 B.n230 10.6151
R1528 B.n234 B.n231 10.6151
R1529 B.n235 B.n234 10.6151
R1530 B.n238 B.n235 10.6151
R1531 B.n239 B.n238 10.6151
R1532 B.n243 B.n242 10.6151
R1533 B.n246 B.n243 10.6151
R1534 B.n247 B.n246 10.6151
R1535 B.n250 B.n247 10.6151
R1536 B.n251 B.n250 10.6151
R1537 B.n254 B.n251 10.6151
R1538 B.n255 B.n254 10.6151
R1539 B.n258 B.n255 10.6151
R1540 B.n259 B.n258 10.6151
R1541 B.n262 B.n259 10.6151
R1542 B.n263 B.n262 10.6151
R1543 B.n266 B.n263 10.6151
R1544 B.n267 B.n266 10.6151
R1545 B.n270 B.n267 10.6151
R1546 B.n271 B.n270 10.6151
R1547 B.n274 B.n271 10.6151
R1548 B.n275 B.n274 10.6151
R1549 B.n278 B.n275 10.6151
R1550 B.n279 B.n278 10.6151
R1551 B.n282 B.n279 10.6151
R1552 B.n283 B.n282 10.6151
R1553 B.n286 B.n283 10.6151
R1554 B.n287 B.n286 10.6151
R1555 B.n290 B.n287 10.6151
R1556 B.n291 B.n290 10.6151
R1557 B.n294 B.n291 10.6151
R1558 B.n295 B.n294 10.6151
R1559 B.n298 B.n295 10.6151
R1560 B.n299 B.n298 10.6151
R1561 B.n302 B.n299 10.6151
R1562 B.n303 B.n302 10.6151
R1563 B.n306 B.n303 10.6151
R1564 B.n307 B.n306 10.6151
R1565 B.n310 B.n307 10.6151
R1566 B.n311 B.n310 10.6151
R1567 B.n314 B.n311 10.6151
R1568 B.n315 B.n314 10.6151
R1569 B.n318 B.n315 10.6151
R1570 B.n319 B.n318 10.6151
R1571 B.n322 B.n319 10.6151
R1572 B.n323 B.n322 10.6151
R1573 B.n326 B.n323 10.6151
R1574 B.n327 B.n326 10.6151
R1575 B.n330 B.n327 10.6151
R1576 B.n331 B.n330 10.6151
R1577 B.n827 B.n331 10.6151
R1578 B.n907 B.n0 8.11757
R1579 B.n907 B.n1 8.11757
R1580 B.n569 B.n459 6.5566
R1581 B.n553 B.n552 6.5566
R1582 B.n223 B.n222 6.5566
R1583 B.n239 B.n125 6.5566
R1584 B.n572 B.n459 4.05904
R1585 B.n552 B.n551 4.05904
R1586 B.n222 B.n221 4.05904
R1587 B.n242 B.n125 4.05904
R1588 B.n761 B.t1 1.15627
R1589 B.t3 B.n893 1.15627
R1590 VN.n1 VN.t2 145.775
R1591 VN.n0 VN.t0 145.775
R1592 VN.n1 VN.t3 144.788
R1593 VN.n0 VN.t1 144.788
R1594 VN VN.n1 52.0381
R1595 VN VN.n0 3.03434
R1596 VDD2.n2 VDD2.n0 109.082
R1597 VDD2.n2 VDD2.n1 64.9457
R1598 VDD2.n1 VDD2.t0 1.43945
R1599 VDD2.n1 VDD2.t1 1.43945
R1600 VDD2.n0 VDD2.t3 1.43945
R1601 VDD2.n0 VDD2.t2 1.43945
R1602 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 5.41641f
C1 VP VDD1 5.79237f
C2 VDD1 VDD2 1.1182f
C3 VP VDD2 0.41896f
C4 VN VDD1 0.149818f
C5 VN VP 6.78888f
C6 VN VDD2 5.52406f
C7 VTAIL VDD1 5.88206f
C8 VP VTAIL 5.43051f
C9 VTAIL VDD2 5.93882f
C10 VDD2 B 4.121726f
C11 VDD1 B 8.59868f
C12 VTAIL B 11.350632f
C13 VN B 11.557321f
C14 VP B 9.875049f
C15 VDD2.t3 B 0.289904f
C16 VDD2.t2 B 0.289904f
C17 VDD2.n0 B 3.34145f
C18 VDD2.t0 B 0.289904f
C19 VDD2.t1 B 0.289904f
C20 VDD2.n1 B 2.61374f
C21 VDD2.n2 B 4.03432f
C22 VN.t1 B 2.80156f
C23 VN.t0 B 2.80853f
C24 VN.n0 B 1.75357f
C25 VN.t2 B 2.80853f
C26 VN.t3 B 2.80156f
C27 VN.n1 B 3.14535f
C28 VDD1.t2 B 0.294986f
C29 VDD1.t3 B 0.294986f
C30 VDD1.n0 B 2.65998f
C31 VDD1.t1 B 0.294986f
C32 VDD1.t0 B 0.294986f
C33 VDD1.n1 B 3.42707f
C34 VTAIL.t3 B 1.96727f
C35 VTAIL.n0 B 0.305632f
C36 VTAIL.t4 B 1.96727f
C37 VTAIL.n1 B 0.376917f
C38 VTAIL.t7 B 1.96727f
C39 VTAIL.n2 B 1.33854f
C40 VTAIL.t0 B 1.96727f
C41 VTAIL.n3 B 1.33854f
C42 VTAIL.t1 B 1.96727f
C43 VTAIL.n4 B 0.376915f
C44 VTAIL.t5 B 1.96727f
C45 VTAIL.n5 B 0.376915f
C46 VTAIL.t6 B 1.96727f
C47 VTAIL.n6 B 1.33854f
C48 VTAIL.t2 B 1.96727f
C49 VTAIL.n7 B 1.2612f
C50 VP.t3 B 2.6068f
C51 VP.n0 B 1.00223f
C52 VP.n1 B 0.023248f
C53 VP.n2 B 0.033794f
C54 VP.n3 B 0.037516f
C55 VP.t2 B 2.6068f
C56 VP.t1 B 2.86131f
C57 VP.t0 B 2.85422f
C58 VP.n4 B 3.19516f
C59 VP.n5 B 1.37766f
C60 VP.n6 B 1.00223f
C61 VP.n7 B 0.039067f
C62 VP.n8 B 0.043111f
C63 VP.n9 B 0.023248f
C64 VP.n10 B 0.023248f
C65 VP.n11 B 0.023248f
C66 VP.n12 B 0.033794f
C67 VP.n13 B 0.043111f
C68 VP.n14 B 0.039067f
C69 VP.n15 B 0.037516f
C70 VP.n16 B 0.048384f
.ends

