* NGSPICE file created from diff_pair_sample_0118.ext - technology: sky130A

.subckt diff_pair_sample_0118 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t15 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.72
X1 B.t11 B.t9 B.t10 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.72
X2 VDD1.t9 VP.t0 VTAIL.t2 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.72
X3 B.t8 B.t6 B.t7 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.72
X4 VDD1.t8 VP.t1 VTAIL.t18 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X5 VDD2.t8 VN.t1 VTAIL.t9 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X6 VTAIL.t5 VP.t2 VDD1.t7 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X7 VDD2.t7 VN.t2 VTAIL.t13 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.72
X8 VTAIL.t0 VP.t3 VDD1.t6 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X9 VTAIL.t14 VN.t3 VDD2.t6 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X10 VDD1.t5 VP.t4 VTAIL.t19 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.72
X11 VDD2.t5 VN.t4 VTAIL.t16 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.72
X12 VTAIL.t12 VN.t5 VDD2.t4 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X13 VTAIL.t1 VP.t5 VDD1.t4 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X14 VDD1.t3 VP.t6 VTAIL.t4 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.72
X15 VDD2.t3 VN.t6 VTAIL.t10 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X16 B.t5 B.t3 B.t4 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.72
X17 VDD1.t2 VP.t7 VTAIL.t7 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.72
X18 VTAIL.t6 VP.t8 VDD1.t1 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X19 VTAIL.t11 VN.t7 VDD2.t2 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X20 VDD2.t1 VN.t8 VTAIL.t17 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.72
X21 VTAIL.t8 VN.t9 VDD2.t0 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
X22 B.t2 B.t0 B.t1 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.72
X23 VDD1.t0 VP.t9 VTAIL.t3 w_n2230_n4576# sky130_fd_pr__pfet_01v8 ad=2.9766 pd=18.37 as=2.9766 ps=18.37 w=18.04 l=0.72
R0 VN.n3 VN.t8 682.245
R1 VN.n17 VN.t2 682.245
R2 VN.n4 VN.t3 658.399
R3 VN.n6 VN.t1 658.399
R4 VN.n10 VN.t9 658.399
R5 VN.n12 VN.t4 658.399
R6 VN.n18 VN.t5 658.399
R7 VN.n20 VN.t6 658.399
R8 VN.n24 VN.t7 658.399
R9 VN.n26 VN.t0 658.399
R10 VN.n13 VN.n12 161.3
R11 VN.n27 VN.n26 161.3
R12 VN.n25 VN.n14 161.3
R13 VN.n24 VN.n23 161.3
R14 VN.n22 VN.n15 161.3
R15 VN.n21 VN.n20 161.3
R16 VN.n19 VN.n16 161.3
R17 VN.n11 VN.n0 161.3
R18 VN.n10 VN.n9 161.3
R19 VN.n8 VN.n1 161.3
R20 VN.n7 VN.n6 161.3
R21 VN.n5 VN.n2 161.3
R22 VN VN.n27 47.885
R23 VN.n17 VN.n16 44.9119
R24 VN.n3 VN.n2 44.9119
R25 VN.n12 VN.n11 35.055
R26 VN.n26 VN.n25 35.055
R27 VN.n5 VN.n4 27.752
R28 VN.n10 VN.n1 27.752
R29 VN.n19 VN.n18 27.752
R30 VN.n24 VN.n15 27.752
R31 VN.n6 VN.n5 20.449
R32 VN.n6 VN.n1 20.449
R33 VN.n20 VN.n19 20.449
R34 VN.n20 VN.n15 20.449
R35 VN.n4 VN.n3 17.739
R36 VN.n18 VN.n17 17.739
R37 VN.n11 VN.n10 13.146
R38 VN.n25 VN.n24 13.146
R39 VN.n27 VN.n14 0.189894
R40 VN.n23 VN.n14 0.189894
R41 VN.n23 VN.n22 0.189894
R42 VN.n22 VN.n21 0.189894
R43 VN.n21 VN.n16 0.189894
R44 VN.n7 VN.n2 0.189894
R45 VN.n8 VN.n7 0.189894
R46 VN.n9 VN.n8 0.189894
R47 VN.n9 VN.n0 0.189894
R48 VN.n13 VN.n0 0.189894
R49 VN VN.n13 0.0516364
R50 VTAIL.n412 VTAIL.n411 756.745
R51 VTAIL.n100 VTAIL.n99 756.745
R52 VTAIL.n312 VTAIL.n311 756.745
R53 VTAIL.n208 VTAIL.n207 756.745
R54 VTAIL.n347 VTAIL.n346 585
R55 VTAIL.n344 VTAIL.n343 585
R56 VTAIL.n353 VTAIL.n352 585
R57 VTAIL.n355 VTAIL.n354 585
R58 VTAIL.n340 VTAIL.n339 585
R59 VTAIL.n361 VTAIL.n360 585
R60 VTAIL.n364 VTAIL.n363 585
R61 VTAIL.n362 VTAIL.n336 585
R62 VTAIL.n369 VTAIL.n335 585
R63 VTAIL.n371 VTAIL.n370 585
R64 VTAIL.n373 VTAIL.n372 585
R65 VTAIL.n332 VTAIL.n331 585
R66 VTAIL.n379 VTAIL.n378 585
R67 VTAIL.n381 VTAIL.n380 585
R68 VTAIL.n328 VTAIL.n327 585
R69 VTAIL.n387 VTAIL.n386 585
R70 VTAIL.n389 VTAIL.n388 585
R71 VTAIL.n324 VTAIL.n323 585
R72 VTAIL.n395 VTAIL.n394 585
R73 VTAIL.n397 VTAIL.n396 585
R74 VTAIL.n320 VTAIL.n319 585
R75 VTAIL.n403 VTAIL.n402 585
R76 VTAIL.n405 VTAIL.n404 585
R77 VTAIL.n316 VTAIL.n315 585
R78 VTAIL.n411 VTAIL.n410 585
R79 VTAIL.n35 VTAIL.n34 585
R80 VTAIL.n32 VTAIL.n31 585
R81 VTAIL.n41 VTAIL.n40 585
R82 VTAIL.n43 VTAIL.n42 585
R83 VTAIL.n28 VTAIL.n27 585
R84 VTAIL.n49 VTAIL.n48 585
R85 VTAIL.n52 VTAIL.n51 585
R86 VTAIL.n50 VTAIL.n24 585
R87 VTAIL.n57 VTAIL.n23 585
R88 VTAIL.n59 VTAIL.n58 585
R89 VTAIL.n61 VTAIL.n60 585
R90 VTAIL.n20 VTAIL.n19 585
R91 VTAIL.n67 VTAIL.n66 585
R92 VTAIL.n69 VTAIL.n68 585
R93 VTAIL.n16 VTAIL.n15 585
R94 VTAIL.n75 VTAIL.n74 585
R95 VTAIL.n77 VTAIL.n76 585
R96 VTAIL.n12 VTAIL.n11 585
R97 VTAIL.n83 VTAIL.n82 585
R98 VTAIL.n85 VTAIL.n84 585
R99 VTAIL.n8 VTAIL.n7 585
R100 VTAIL.n91 VTAIL.n90 585
R101 VTAIL.n93 VTAIL.n92 585
R102 VTAIL.n4 VTAIL.n3 585
R103 VTAIL.n99 VTAIL.n98 585
R104 VTAIL.n311 VTAIL.n310 585
R105 VTAIL.n216 VTAIL.n215 585
R106 VTAIL.n305 VTAIL.n304 585
R107 VTAIL.n303 VTAIL.n302 585
R108 VTAIL.n220 VTAIL.n219 585
R109 VTAIL.n297 VTAIL.n296 585
R110 VTAIL.n295 VTAIL.n294 585
R111 VTAIL.n224 VTAIL.n223 585
R112 VTAIL.n289 VTAIL.n288 585
R113 VTAIL.n287 VTAIL.n286 585
R114 VTAIL.n228 VTAIL.n227 585
R115 VTAIL.n281 VTAIL.n280 585
R116 VTAIL.n279 VTAIL.n278 585
R117 VTAIL.n232 VTAIL.n231 585
R118 VTAIL.n273 VTAIL.n272 585
R119 VTAIL.n271 VTAIL.n270 585
R120 VTAIL.n269 VTAIL.n235 585
R121 VTAIL.n239 VTAIL.n236 585
R122 VTAIL.n264 VTAIL.n263 585
R123 VTAIL.n262 VTAIL.n261 585
R124 VTAIL.n241 VTAIL.n240 585
R125 VTAIL.n256 VTAIL.n255 585
R126 VTAIL.n254 VTAIL.n253 585
R127 VTAIL.n245 VTAIL.n244 585
R128 VTAIL.n248 VTAIL.n247 585
R129 VTAIL.n207 VTAIL.n206 585
R130 VTAIL.n112 VTAIL.n111 585
R131 VTAIL.n201 VTAIL.n200 585
R132 VTAIL.n199 VTAIL.n198 585
R133 VTAIL.n116 VTAIL.n115 585
R134 VTAIL.n193 VTAIL.n192 585
R135 VTAIL.n191 VTAIL.n190 585
R136 VTAIL.n120 VTAIL.n119 585
R137 VTAIL.n185 VTAIL.n184 585
R138 VTAIL.n183 VTAIL.n182 585
R139 VTAIL.n124 VTAIL.n123 585
R140 VTAIL.n177 VTAIL.n176 585
R141 VTAIL.n175 VTAIL.n174 585
R142 VTAIL.n128 VTAIL.n127 585
R143 VTAIL.n169 VTAIL.n168 585
R144 VTAIL.n167 VTAIL.n166 585
R145 VTAIL.n165 VTAIL.n131 585
R146 VTAIL.n135 VTAIL.n132 585
R147 VTAIL.n160 VTAIL.n159 585
R148 VTAIL.n158 VTAIL.n157 585
R149 VTAIL.n137 VTAIL.n136 585
R150 VTAIL.n152 VTAIL.n151 585
R151 VTAIL.n150 VTAIL.n149 585
R152 VTAIL.n141 VTAIL.n140 585
R153 VTAIL.n144 VTAIL.n143 585
R154 VTAIL.t16 VTAIL.n345 329.036
R155 VTAIL.t7 VTAIL.n33 329.036
R156 VTAIL.t13 VTAIL.n142 329.036
R157 VTAIL.t19 VTAIL.n246 329.036
R158 VTAIL.n346 VTAIL.n343 171.744
R159 VTAIL.n353 VTAIL.n343 171.744
R160 VTAIL.n354 VTAIL.n353 171.744
R161 VTAIL.n354 VTAIL.n339 171.744
R162 VTAIL.n361 VTAIL.n339 171.744
R163 VTAIL.n363 VTAIL.n361 171.744
R164 VTAIL.n363 VTAIL.n362 171.744
R165 VTAIL.n362 VTAIL.n335 171.744
R166 VTAIL.n371 VTAIL.n335 171.744
R167 VTAIL.n372 VTAIL.n371 171.744
R168 VTAIL.n372 VTAIL.n331 171.744
R169 VTAIL.n379 VTAIL.n331 171.744
R170 VTAIL.n380 VTAIL.n379 171.744
R171 VTAIL.n380 VTAIL.n327 171.744
R172 VTAIL.n387 VTAIL.n327 171.744
R173 VTAIL.n388 VTAIL.n387 171.744
R174 VTAIL.n388 VTAIL.n323 171.744
R175 VTAIL.n395 VTAIL.n323 171.744
R176 VTAIL.n396 VTAIL.n395 171.744
R177 VTAIL.n396 VTAIL.n319 171.744
R178 VTAIL.n403 VTAIL.n319 171.744
R179 VTAIL.n404 VTAIL.n403 171.744
R180 VTAIL.n404 VTAIL.n315 171.744
R181 VTAIL.n411 VTAIL.n315 171.744
R182 VTAIL.n34 VTAIL.n31 171.744
R183 VTAIL.n41 VTAIL.n31 171.744
R184 VTAIL.n42 VTAIL.n41 171.744
R185 VTAIL.n42 VTAIL.n27 171.744
R186 VTAIL.n49 VTAIL.n27 171.744
R187 VTAIL.n51 VTAIL.n49 171.744
R188 VTAIL.n51 VTAIL.n50 171.744
R189 VTAIL.n50 VTAIL.n23 171.744
R190 VTAIL.n59 VTAIL.n23 171.744
R191 VTAIL.n60 VTAIL.n59 171.744
R192 VTAIL.n60 VTAIL.n19 171.744
R193 VTAIL.n67 VTAIL.n19 171.744
R194 VTAIL.n68 VTAIL.n67 171.744
R195 VTAIL.n68 VTAIL.n15 171.744
R196 VTAIL.n75 VTAIL.n15 171.744
R197 VTAIL.n76 VTAIL.n75 171.744
R198 VTAIL.n76 VTAIL.n11 171.744
R199 VTAIL.n83 VTAIL.n11 171.744
R200 VTAIL.n84 VTAIL.n83 171.744
R201 VTAIL.n84 VTAIL.n7 171.744
R202 VTAIL.n91 VTAIL.n7 171.744
R203 VTAIL.n92 VTAIL.n91 171.744
R204 VTAIL.n92 VTAIL.n3 171.744
R205 VTAIL.n99 VTAIL.n3 171.744
R206 VTAIL.n311 VTAIL.n215 171.744
R207 VTAIL.n304 VTAIL.n215 171.744
R208 VTAIL.n304 VTAIL.n303 171.744
R209 VTAIL.n303 VTAIL.n219 171.744
R210 VTAIL.n296 VTAIL.n219 171.744
R211 VTAIL.n296 VTAIL.n295 171.744
R212 VTAIL.n295 VTAIL.n223 171.744
R213 VTAIL.n288 VTAIL.n223 171.744
R214 VTAIL.n288 VTAIL.n287 171.744
R215 VTAIL.n287 VTAIL.n227 171.744
R216 VTAIL.n280 VTAIL.n227 171.744
R217 VTAIL.n280 VTAIL.n279 171.744
R218 VTAIL.n279 VTAIL.n231 171.744
R219 VTAIL.n272 VTAIL.n231 171.744
R220 VTAIL.n272 VTAIL.n271 171.744
R221 VTAIL.n271 VTAIL.n235 171.744
R222 VTAIL.n239 VTAIL.n235 171.744
R223 VTAIL.n263 VTAIL.n239 171.744
R224 VTAIL.n263 VTAIL.n262 171.744
R225 VTAIL.n262 VTAIL.n240 171.744
R226 VTAIL.n255 VTAIL.n240 171.744
R227 VTAIL.n255 VTAIL.n254 171.744
R228 VTAIL.n254 VTAIL.n244 171.744
R229 VTAIL.n247 VTAIL.n244 171.744
R230 VTAIL.n207 VTAIL.n111 171.744
R231 VTAIL.n200 VTAIL.n111 171.744
R232 VTAIL.n200 VTAIL.n199 171.744
R233 VTAIL.n199 VTAIL.n115 171.744
R234 VTAIL.n192 VTAIL.n115 171.744
R235 VTAIL.n192 VTAIL.n191 171.744
R236 VTAIL.n191 VTAIL.n119 171.744
R237 VTAIL.n184 VTAIL.n119 171.744
R238 VTAIL.n184 VTAIL.n183 171.744
R239 VTAIL.n183 VTAIL.n123 171.744
R240 VTAIL.n176 VTAIL.n123 171.744
R241 VTAIL.n176 VTAIL.n175 171.744
R242 VTAIL.n175 VTAIL.n127 171.744
R243 VTAIL.n168 VTAIL.n127 171.744
R244 VTAIL.n168 VTAIL.n167 171.744
R245 VTAIL.n167 VTAIL.n131 171.744
R246 VTAIL.n135 VTAIL.n131 171.744
R247 VTAIL.n159 VTAIL.n135 171.744
R248 VTAIL.n159 VTAIL.n158 171.744
R249 VTAIL.n158 VTAIL.n136 171.744
R250 VTAIL.n151 VTAIL.n136 171.744
R251 VTAIL.n151 VTAIL.n150 171.744
R252 VTAIL.n150 VTAIL.n140 171.744
R253 VTAIL.n143 VTAIL.n140 171.744
R254 VTAIL.n346 VTAIL.t16 85.8723
R255 VTAIL.n34 VTAIL.t7 85.8723
R256 VTAIL.n247 VTAIL.t19 85.8723
R257 VTAIL.n143 VTAIL.t13 85.8723
R258 VTAIL.n213 VTAIL.n212 54.763
R259 VTAIL.n211 VTAIL.n210 54.763
R260 VTAIL.n109 VTAIL.n108 54.763
R261 VTAIL.n107 VTAIL.n106 54.763
R262 VTAIL.n415 VTAIL.n414 54.7629
R263 VTAIL.n1 VTAIL.n0 54.7629
R264 VTAIL.n103 VTAIL.n102 54.7629
R265 VTAIL.n105 VTAIL.n104 54.7629
R266 VTAIL.n413 VTAIL.n412 34.1247
R267 VTAIL.n101 VTAIL.n100 34.1247
R268 VTAIL.n313 VTAIL.n312 34.1247
R269 VTAIL.n209 VTAIL.n208 34.1247
R270 VTAIL.n107 VTAIL.n105 29.7289
R271 VTAIL.n413 VTAIL.n313 28.8238
R272 VTAIL.n370 VTAIL.n369 13.1884
R273 VTAIL.n58 VTAIL.n57 13.1884
R274 VTAIL.n270 VTAIL.n269 13.1884
R275 VTAIL.n166 VTAIL.n165 13.1884
R276 VTAIL.n368 VTAIL.n336 12.8005
R277 VTAIL.n373 VTAIL.n334 12.8005
R278 VTAIL.n56 VTAIL.n24 12.8005
R279 VTAIL.n61 VTAIL.n22 12.8005
R280 VTAIL.n273 VTAIL.n234 12.8005
R281 VTAIL.n268 VTAIL.n236 12.8005
R282 VTAIL.n169 VTAIL.n130 12.8005
R283 VTAIL.n164 VTAIL.n132 12.8005
R284 VTAIL.n365 VTAIL.n364 12.0247
R285 VTAIL.n374 VTAIL.n332 12.0247
R286 VTAIL.n410 VTAIL.n314 12.0247
R287 VTAIL.n53 VTAIL.n52 12.0247
R288 VTAIL.n62 VTAIL.n20 12.0247
R289 VTAIL.n98 VTAIL.n2 12.0247
R290 VTAIL.n310 VTAIL.n214 12.0247
R291 VTAIL.n274 VTAIL.n232 12.0247
R292 VTAIL.n265 VTAIL.n264 12.0247
R293 VTAIL.n206 VTAIL.n110 12.0247
R294 VTAIL.n170 VTAIL.n128 12.0247
R295 VTAIL.n161 VTAIL.n160 12.0247
R296 VTAIL.n360 VTAIL.n338 11.249
R297 VTAIL.n378 VTAIL.n377 11.249
R298 VTAIL.n409 VTAIL.n316 11.249
R299 VTAIL.n48 VTAIL.n26 11.249
R300 VTAIL.n66 VTAIL.n65 11.249
R301 VTAIL.n97 VTAIL.n4 11.249
R302 VTAIL.n309 VTAIL.n216 11.249
R303 VTAIL.n278 VTAIL.n277 11.249
R304 VTAIL.n261 VTAIL.n238 11.249
R305 VTAIL.n205 VTAIL.n112 11.249
R306 VTAIL.n174 VTAIL.n173 11.249
R307 VTAIL.n157 VTAIL.n134 11.249
R308 VTAIL.n347 VTAIL.n345 10.7239
R309 VTAIL.n35 VTAIL.n33 10.7239
R310 VTAIL.n248 VTAIL.n246 10.7239
R311 VTAIL.n144 VTAIL.n142 10.7239
R312 VTAIL.n359 VTAIL.n340 10.4732
R313 VTAIL.n381 VTAIL.n330 10.4732
R314 VTAIL.n406 VTAIL.n405 10.4732
R315 VTAIL.n47 VTAIL.n28 10.4732
R316 VTAIL.n69 VTAIL.n18 10.4732
R317 VTAIL.n94 VTAIL.n93 10.4732
R318 VTAIL.n306 VTAIL.n305 10.4732
R319 VTAIL.n281 VTAIL.n230 10.4732
R320 VTAIL.n260 VTAIL.n241 10.4732
R321 VTAIL.n202 VTAIL.n201 10.4732
R322 VTAIL.n177 VTAIL.n126 10.4732
R323 VTAIL.n156 VTAIL.n137 10.4732
R324 VTAIL.n356 VTAIL.n355 9.69747
R325 VTAIL.n382 VTAIL.n328 9.69747
R326 VTAIL.n402 VTAIL.n318 9.69747
R327 VTAIL.n44 VTAIL.n43 9.69747
R328 VTAIL.n70 VTAIL.n16 9.69747
R329 VTAIL.n90 VTAIL.n6 9.69747
R330 VTAIL.n302 VTAIL.n218 9.69747
R331 VTAIL.n282 VTAIL.n228 9.69747
R332 VTAIL.n257 VTAIL.n256 9.69747
R333 VTAIL.n198 VTAIL.n114 9.69747
R334 VTAIL.n178 VTAIL.n124 9.69747
R335 VTAIL.n153 VTAIL.n152 9.69747
R336 VTAIL.n408 VTAIL.n314 9.45567
R337 VTAIL.n96 VTAIL.n2 9.45567
R338 VTAIL.n308 VTAIL.n214 9.45567
R339 VTAIL.n204 VTAIL.n110 9.45567
R340 VTAIL.n393 VTAIL.n392 9.3005
R341 VTAIL.n322 VTAIL.n321 9.3005
R342 VTAIL.n399 VTAIL.n398 9.3005
R343 VTAIL.n401 VTAIL.n400 9.3005
R344 VTAIL.n318 VTAIL.n317 9.3005
R345 VTAIL.n407 VTAIL.n406 9.3005
R346 VTAIL.n409 VTAIL.n408 9.3005
R347 VTAIL.n326 VTAIL.n325 9.3005
R348 VTAIL.n385 VTAIL.n384 9.3005
R349 VTAIL.n383 VTAIL.n382 9.3005
R350 VTAIL.n330 VTAIL.n329 9.3005
R351 VTAIL.n377 VTAIL.n376 9.3005
R352 VTAIL.n375 VTAIL.n374 9.3005
R353 VTAIL.n334 VTAIL.n333 9.3005
R354 VTAIL.n349 VTAIL.n348 9.3005
R355 VTAIL.n351 VTAIL.n350 9.3005
R356 VTAIL.n342 VTAIL.n341 9.3005
R357 VTAIL.n357 VTAIL.n356 9.3005
R358 VTAIL.n359 VTAIL.n358 9.3005
R359 VTAIL.n338 VTAIL.n337 9.3005
R360 VTAIL.n366 VTAIL.n365 9.3005
R361 VTAIL.n368 VTAIL.n367 9.3005
R362 VTAIL.n391 VTAIL.n390 9.3005
R363 VTAIL.n81 VTAIL.n80 9.3005
R364 VTAIL.n10 VTAIL.n9 9.3005
R365 VTAIL.n87 VTAIL.n86 9.3005
R366 VTAIL.n89 VTAIL.n88 9.3005
R367 VTAIL.n6 VTAIL.n5 9.3005
R368 VTAIL.n95 VTAIL.n94 9.3005
R369 VTAIL.n97 VTAIL.n96 9.3005
R370 VTAIL.n14 VTAIL.n13 9.3005
R371 VTAIL.n73 VTAIL.n72 9.3005
R372 VTAIL.n71 VTAIL.n70 9.3005
R373 VTAIL.n18 VTAIL.n17 9.3005
R374 VTAIL.n65 VTAIL.n64 9.3005
R375 VTAIL.n63 VTAIL.n62 9.3005
R376 VTAIL.n22 VTAIL.n21 9.3005
R377 VTAIL.n37 VTAIL.n36 9.3005
R378 VTAIL.n39 VTAIL.n38 9.3005
R379 VTAIL.n30 VTAIL.n29 9.3005
R380 VTAIL.n45 VTAIL.n44 9.3005
R381 VTAIL.n47 VTAIL.n46 9.3005
R382 VTAIL.n26 VTAIL.n25 9.3005
R383 VTAIL.n54 VTAIL.n53 9.3005
R384 VTAIL.n56 VTAIL.n55 9.3005
R385 VTAIL.n79 VTAIL.n78 9.3005
R386 VTAIL.n309 VTAIL.n308 9.3005
R387 VTAIL.n307 VTAIL.n306 9.3005
R388 VTAIL.n218 VTAIL.n217 9.3005
R389 VTAIL.n301 VTAIL.n300 9.3005
R390 VTAIL.n299 VTAIL.n298 9.3005
R391 VTAIL.n222 VTAIL.n221 9.3005
R392 VTAIL.n293 VTAIL.n292 9.3005
R393 VTAIL.n291 VTAIL.n290 9.3005
R394 VTAIL.n226 VTAIL.n225 9.3005
R395 VTAIL.n285 VTAIL.n284 9.3005
R396 VTAIL.n283 VTAIL.n282 9.3005
R397 VTAIL.n230 VTAIL.n229 9.3005
R398 VTAIL.n277 VTAIL.n276 9.3005
R399 VTAIL.n275 VTAIL.n274 9.3005
R400 VTAIL.n234 VTAIL.n233 9.3005
R401 VTAIL.n268 VTAIL.n267 9.3005
R402 VTAIL.n266 VTAIL.n265 9.3005
R403 VTAIL.n238 VTAIL.n237 9.3005
R404 VTAIL.n260 VTAIL.n259 9.3005
R405 VTAIL.n258 VTAIL.n257 9.3005
R406 VTAIL.n243 VTAIL.n242 9.3005
R407 VTAIL.n252 VTAIL.n251 9.3005
R408 VTAIL.n250 VTAIL.n249 9.3005
R409 VTAIL.n146 VTAIL.n145 9.3005
R410 VTAIL.n148 VTAIL.n147 9.3005
R411 VTAIL.n139 VTAIL.n138 9.3005
R412 VTAIL.n154 VTAIL.n153 9.3005
R413 VTAIL.n156 VTAIL.n155 9.3005
R414 VTAIL.n134 VTAIL.n133 9.3005
R415 VTAIL.n162 VTAIL.n161 9.3005
R416 VTAIL.n164 VTAIL.n163 9.3005
R417 VTAIL.n118 VTAIL.n117 9.3005
R418 VTAIL.n195 VTAIL.n194 9.3005
R419 VTAIL.n197 VTAIL.n196 9.3005
R420 VTAIL.n114 VTAIL.n113 9.3005
R421 VTAIL.n203 VTAIL.n202 9.3005
R422 VTAIL.n205 VTAIL.n204 9.3005
R423 VTAIL.n189 VTAIL.n188 9.3005
R424 VTAIL.n187 VTAIL.n186 9.3005
R425 VTAIL.n122 VTAIL.n121 9.3005
R426 VTAIL.n181 VTAIL.n180 9.3005
R427 VTAIL.n179 VTAIL.n178 9.3005
R428 VTAIL.n126 VTAIL.n125 9.3005
R429 VTAIL.n173 VTAIL.n172 9.3005
R430 VTAIL.n171 VTAIL.n170 9.3005
R431 VTAIL.n130 VTAIL.n129 9.3005
R432 VTAIL.n352 VTAIL.n342 8.92171
R433 VTAIL.n386 VTAIL.n385 8.92171
R434 VTAIL.n401 VTAIL.n320 8.92171
R435 VTAIL.n40 VTAIL.n30 8.92171
R436 VTAIL.n74 VTAIL.n73 8.92171
R437 VTAIL.n89 VTAIL.n8 8.92171
R438 VTAIL.n301 VTAIL.n220 8.92171
R439 VTAIL.n286 VTAIL.n285 8.92171
R440 VTAIL.n253 VTAIL.n243 8.92171
R441 VTAIL.n197 VTAIL.n116 8.92171
R442 VTAIL.n182 VTAIL.n181 8.92171
R443 VTAIL.n149 VTAIL.n139 8.92171
R444 VTAIL.n351 VTAIL.n344 8.14595
R445 VTAIL.n389 VTAIL.n326 8.14595
R446 VTAIL.n398 VTAIL.n397 8.14595
R447 VTAIL.n39 VTAIL.n32 8.14595
R448 VTAIL.n77 VTAIL.n14 8.14595
R449 VTAIL.n86 VTAIL.n85 8.14595
R450 VTAIL.n298 VTAIL.n297 8.14595
R451 VTAIL.n289 VTAIL.n226 8.14595
R452 VTAIL.n252 VTAIL.n245 8.14595
R453 VTAIL.n194 VTAIL.n193 8.14595
R454 VTAIL.n185 VTAIL.n122 8.14595
R455 VTAIL.n148 VTAIL.n141 8.14595
R456 VTAIL.n348 VTAIL.n347 7.3702
R457 VTAIL.n390 VTAIL.n324 7.3702
R458 VTAIL.n394 VTAIL.n322 7.3702
R459 VTAIL.n36 VTAIL.n35 7.3702
R460 VTAIL.n78 VTAIL.n12 7.3702
R461 VTAIL.n82 VTAIL.n10 7.3702
R462 VTAIL.n294 VTAIL.n222 7.3702
R463 VTAIL.n290 VTAIL.n224 7.3702
R464 VTAIL.n249 VTAIL.n248 7.3702
R465 VTAIL.n190 VTAIL.n118 7.3702
R466 VTAIL.n186 VTAIL.n120 7.3702
R467 VTAIL.n145 VTAIL.n144 7.3702
R468 VTAIL.n393 VTAIL.n324 6.59444
R469 VTAIL.n394 VTAIL.n393 6.59444
R470 VTAIL.n81 VTAIL.n12 6.59444
R471 VTAIL.n82 VTAIL.n81 6.59444
R472 VTAIL.n294 VTAIL.n293 6.59444
R473 VTAIL.n293 VTAIL.n224 6.59444
R474 VTAIL.n190 VTAIL.n189 6.59444
R475 VTAIL.n189 VTAIL.n120 6.59444
R476 VTAIL.n348 VTAIL.n344 5.81868
R477 VTAIL.n390 VTAIL.n389 5.81868
R478 VTAIL.n397 VTAIL.n322 5.81868
R479 VTAIL.n36 VTAIL.n32 5.81868
R480 VTAIL.n78 VTAIL.n77 5.81868
R481 VTAIL.n85 VTAIL.n10 5.81868
R482 VTAIL.n297 VTAIL.n222 5.81868
R483 VTAIL.n290 VTAIL.n289 5.81868
R484 VTAIL.n249 VTAIL.n245 5.81868
R485 VTAIL.n193 VTAIL.n118 5.81868
R486 VTAIL.n186 VTAIL.n185 5.81868
R487 VTAIL.n145 VTAIL.n141 5.81868
R488 VTAIL.n352 VTAIL.n351 5.04292
R489 VTAIL.n386 VTAIL.n326 5.04292
R490 VTAIL.n398 VTAIL.n320 5.04292
R491 VTAIL.n40 VTAIL.n39 5.04292
R492 VTAIL.n74 VTAIL.n14 5.04292
R493 VTAIL.n86 VTAIL.n8 5.04292
R494 VTAIL.n298 VTAIL.n220 5.04292
R495 VTAIL.n286 VTAIL.n226 5.04292
R496 VTAIL.n253 VTAIL.n252 5.04292
R497 VTAIL.n194 VTAIL.n116 5.04292
R498 VTAIL.n182 VTAIL.n122 5.04292
R499 VTAIL.n149 VTAIL.n148 5.04292
R500 VTAIL.n355 VTAIL.n342 4.26717
R501 VTAIL.n385 VTAIL.n328 4.26717
R502 VTAIL.n402 VTAIL.n401 4.26717
R503 VTAIL.n43 VTAIL.n30 4.26717
R504 VTAIL.n73 VTAIL.n16 4.26717
R505 VTAIL.n90 VTAIL.n89 4.26717
R506 VTAIL.n302 VTAIL.n301 4.26717
R507 VTAIL.n285 VTAIL.n228 4.26717
R508 VTAIL.n256 VTAIL.n243 4.26717
R509 VTAIL.n198 VTAIL.n197 4.26717
R510 VTAIL.n181 VTAIL.n124 4.26717
R511 VTAIL.n152 VTAIL.n139 4.26717
R512 VTAIL.n356 VTAIL.n340 3.49141
R513 VTAIL.n382 VTAIL.n381 3.49141
R514 VTAIL.n405 VTAIL.n318 3.49141
R515 VTAIL.n44 VTAIL.n28 3.49141
R516 VTAIL.n70 VTAIL.n69 3.49141
R517 VTAIL.n93 VTAIL.n6 3.49141
R518 VTAIL.n305 VTAIL.n218 3.49141
R519 VTAIL.n282 VTAIL.n281 3.49141
R520 VTAIL.n257 VTAIL.n241 3.49141
R521 VTAIL.n201 VTAIL.n114 3.49141
R522 VTAIL.n178 VTAIL.n177 3.49141
R523 VTAIL.n153 VTAIL.n137 3.49141
R524 VTAIL.n360 VTAIL.n359 2.71565
R525 VTAIL.n378 VTAIL.n330 2.71565
R526 VTAIL.n406 VTAIL.n316 2.71565
R527 VTAIL.n48 VTAIL.n47 2.71565
R528 VTAIL.n66 VTAIL.n18 2.71565
R529 VTAIL.n94 VTAIL.n4 2.71565
R530 VTAIL.n306 VTAIL.n216 2.71565
R531 VTAIL.n278 VTAIL.n230 2.71565
R532 VTAIL.n261 VTAIL.n260 2.71565
R533 VTAIL.n202 VTAIL.n112 2.71565
R534 VTAIL.n174 VTAIL.n126 2.71565
R535 VTAIL.n157 VTAIL.n156 2.71565
R536 VTAIL.n349 VTAIL.n345 2.41282
R537 VTAIL.n37 VTAIL.n33 2.41282
R538 VTAIL.n250 VTAIL.n246 2.41282
R539 VTAIL.n146 VTAIL.n142 2.41282
R540 VTAIL.n364 VTAIL.n338 1.93989
R541 VTAIL.n377 VTAIL.n332 1.93989
R542 VTAIL.n410 VTAIL.n409 1.93989
R543 VTAIL.n52 VTAIL.n26 1.93989
R544 VTAIL.n65 VTAIL.n20 1.93989
R545 VTAIL.n98 VTAIL.n97 1.93989
R546 VTAIL.n310 VTAIL.n309 1.93989
R547 VTAIL.n277 VTAIL.n232 1.93989
R548 VTAIL.n264 VTAIL.n238 1.93989
R549 VTAIL.n206 VTAIL.n205 1.93989
R550 VTAIL.n173 VTAIL.n128 1.93989
R551 VTAIL.n160 VTAIL.n134 1.93989
R552 VTAIL.n414 VTAIL.t9 1.80233
R553 VTAIL.n414 VTAIL.t8 1.80233
R554 VTAIL.n0 VTAIL.t17 1.80233
R555 VTAIL.n0 VTAIL.t14 1.80233
R556 VTAIL.n102 VTAIL.t3 1.80233
R557 VTAIL.n102 VTAIL.t0 1.80233
R558 VTAIL.n104 VTAIL.t2 1.80233
R559 VTAIL.n104 VTAIL.t1 1.80233
R560 VTAIL.n212 VTAIL.t18 1.80233
R561 VTAIL.n212 VTAIL.t5 1.80233
R562 VTAIL.n210 VTAIL.t4 1.80233
R563 VTAIL.n210 VTAIL.t6 1.80233
R564 VTAIL.n108 VTAIL.t10 1.80233
R565 VTAIL.n108 VTAIL.t12 1.80233
R566 VTAIL.n106 VTAIL.t15 1.80233
R567 VTAIL.n106 VTAIL.t11 1.80233
R568 VTAIL.n365 VTAIL.n336 1.16414
R569 VTAIL.n374 VTAIL.n373 1.16414
R570 VTAIL.n412 VTAIL.n314 1.16414
R571 VTAIL.n53 VTAIL.n24 1.16414
R572 VTAIL.n62 VTAIL.n61 1.16414
R573 VTAIL.n100 VTAIL.n2 1.16414
R574 VTAIL.n312 VTAIL.n214 1.16414
R575 VTAIL.n274 VTAIL.n273 1.16414
R576 VTAIL.n265 VTAIL.n236 1.16414
R577 VTAIL.n208 VTAIL.n110 1.16414
R578 VTAIL.n170 VTAIL.n169 1.16414
R579 VTAIL.n161 VTAIL.n132 1.16414
R580 VTAIL.n211 VTAIL.n209 0.922914
R581 VTAIL.n101 VTAIL.n1 0.922914
R582 VTAIL.n109 VTAIL.n107 0.905672
R583 VTAIL.n209 VTAIL.n109 0.905672
R584 VTAIL.n213 VTAIL.n211 0.905672
R585 VTAIL.n313 VTAIL.n213 0.905672
R586 VTAIL.n105 VTAIL.n103 0.905672
R587 VTAIL.n103 VTAIL.n101 0.905672
R588 VTAIL.n415 VTAIL.n413 0.905672
R589 VTAIL VTAIL.n1 0.737569
R590 VTAIL.n369 VTAIL.n368 0.388379
R591 VTAIL.n370 VTAIL.n334 0.388379
R592 VTAIL.n57 VTAIL.n56 0.388379
R593 VTAIL.n58 VTAIL.n22 0.388379
R594 VTAIL.n270 VTAIL.n234 0.388379
R595 VTAIL.n269 VTAIL.n268 0.388379
R596 VTAIL.n166 VTAIL.n130 0.388379
R597 VTAIL.n165 VTAIL.n164 0.388379
R598 VTAIL VTAIL.n415 0.168603
R599 VTAIL.n350 VTAIL.n349 0.155672
R600 VTAIL.n350 VTAIL.n341 0.155672
R601 VTAIL.n357 VTAIL.n341 0.155672
R602 VTAIL.n358 VTAIL.n357 0.155672
R603 VTAIL.n358 VTAIL.n337 0.155672
R604 VTAIL.n366 VTAIL.n337 0.155672
R605 VTAIL.n367 VTAIL.n366 0.155672
R606 VTAIL.n367 VTAIL.n333 0.155672
R607 VTAIL.n375 VTAIL.n333 0.155672
R608 VTAIL.n376 VTAIL.n375 0.155672
R609 VTAIL.n376 VTAIL.n329 0.155672
R610 VTAIL.n383 VTAIL.n329 0.155672
R611 VTAIL.n384 VTAIL.n383 0.155672
R612 VTAIL.n384 VTAIL.n325 0.155672
R613 VTAIL.n391 VTAIL.n325 0.155672
R614 VTAIL.n392 VTAIL.n391 0.155672
R615 VTAIL.n392 VTAIL.n321 0.155672
R616 VTAIL.n399 VTAIL.n321 0.155672
R617 VTAIL.n400 VTAIL.n399 0.155672
R618 VTAIL.n400 VTAIL.n317 0.155672
R619 VTAIL.n407 VTAIL.n317 0.155672
R620 VTAIL.n408 VTAIL.n407 0.155672
R621 VTAIL.n38 VTAIL.n37 0.155672
R622 VTAIL.n38 VTAIL.n29 0.155672
R623 VTAIL.n45 VTAIL.n29 0.155672
R624 VTAIL.n46 VTAIL.n45 0.155672
R625 VTAIL.n46 VTAIL.n25 0.155672
R626 VTAIL.n54 VTAIL.n25 0.155672
R627 VTAIL.n55 VTAIL.n54 0.155672
R628 VTAIL.n55 VTAIL.n21 0.155672
R629 VTAIL.n63 VTAIL.n21 0.155672
R630 VTAIL.n64 VTAIL.n63 0.155672
R631 VTAIL.n64 VTAIL.n17 0.155672
R632 VTAIL.n71 VTAIL.n17 0.155672
R633 VTAIL.n72 VTAIL.n71 0.155672
R634 VTAIL.n72 VTAIL.n13 0.155672
R635 VTAIL.n79 VTAIL.n13 0.155672
R636 VTAIL.n80 VTAIL.n79 0.155672
R637 VTAIL.n80 VTAIL.n9 0.155672
R638 VTAIL.n87 VTAIL.n9 0.155672
R639 VTAIL.n88 VTAIL.n87 0.155672
R640 VTAIL.n88 VTAIL.n5 0.155672
R641 VTAIL.n95 VTAIL.n5 0.155672
R642 VTAIL.n96 VTAIL.n95 0.155672
R643 VTAIL.n308 VTAIL.n307 0.155672
R644 VTAIL.n307 VTAIL.n217 0.155672
R645 VTAIL.n300 VTAIL.n217 0.155672
R646 VTAIL.n300 VTAIL.n299 0.155672
R647 VTAIL.n299 VTAIL.n221 0.155672
R648 VTAIL.n292 VTAIL.n221 0.155672
R649 VTAIL.n292 VTAIL.n291 0.155672
R650 VTAIL.n291 VTAIL.n225 0.155672
R651 VTAIL.n284 VTAIL.n225 0.155672
R652 VTAIL.n284 VTAIL.n283 0.155672
R653 VTAIL.n283 VTAIL.n229 0.155672
R654 VTAIL.n276 VTAIL.n229 0.155672
R655 VTAIL.n276 VTAIL.n275 0.155672
R656 VTAIL.n275 VTAIL.n233 0.155672
R657 VTAIL.n267 VTAIL.n233 0.155672
R658 VTAIL.n267 VTAIL.n266 0.155672
R659 VTAIL.n266 VTAIL.n237 0.155672
R660 VTAIL.n259 VTAIL.n237 0.155672
R661 VTAIL.n259 VTAIL.n258 0.155672
R662 VTAIL.n258 VTAIL.n242 0.155672
R663 VTAIL.n251 VTAIL.n242 0.155672
R664 VTAIL.n251 VTAIL.n250 0.155672
R665 VTAIL.n204 VTAIL.n203 0.155672
R666 VTAIL.n203 VTAIL.n113 0.155672
R667 VTAIL.n196 VTAIL.n113 0.155672
R668 VTAIL.n196 VTAIL.n195 0.155672
R669 VTAIL.n195 VTAIL.n117 0.155672
R670 VTAIL.n188 VTAIL.n117 0.155672
R671 VTAIL.n188 VTAIL.n187 0.155672
R672 VTAIL.n187 VTAIL.n121 0.155672
R673 VTAIL.n180 VTAIL.n121 0.155672
R674 VTAIL.n180 VTAIL.n179 0.155672
R675 VTAIL.n179 VTAIL.n125 0.155672
R676 VTAIL.n172 VTAIL.n125 0.155672
R677 VTAIL.n172 VTAIL.n171 0.155672
R678 VTAIL.n171 VTAIL.n129 0.155672
R679 VTAIL.n163 VTAIL.n129 0.155672
R680 VTAIL.n163 VTAIL.n162 0.155672
R681 VTAIL.n162 VTAIL.n133 0.155672
R682 VTAIL.n155 VTAIL.n133 0.155672
R683 VTAIL.n155 VTAIL.n154 0.155672
R684 VTAIL.n154 VTAIL.n138 0.155672
R685 VTAIL.n147 VTAIL.n138 0.155672
R686 VTAIL.n147 VTAIL.n146 0.155672
R687 VDD2.n201 VDD2.n200 756.745
R688 VDD2.n98 VDD2.n97 756.745
R689 VDD2.n200 VDD2.n199 585
R690 VDD2.n105 VDD2.n104 585
R691 VDD2.n194 VDD2.n193 585
R692 VDD2.n192 VDD2.n191 585
R693 VDD2.n109 VDD2.n108 585
R694 VDD2.n186 VDD2.n185 585
R695 VDD2.n184 VDD2.n183 585
R696 VDD2.n113 VDD2.n112 585
R697 VDD2.n178 VDD2.n177 585
R698 VDD2.n176 VDD2.n175 585
R699 VDD2.n117 VDD2.n116 585
R700 VDD2.n170 VDD2.n169 585
R701 VDD2.n168 VDD2.n167 585
R702 VDD2.n121 VDD2.n120 585
R703 VDD2.n162 VDD2.n161 585
R704 VDD2.n160 VDD2.n159 585
R705 VDD2.n158 VDD2.n124 585
R706 VDD2.n128 VDD2.n125 585
R707 VDD2.n153 VDD2.n152 585
R708 VDD2.n151 VDD2.n150 585
R709 VDD2.n130 VDD2.n129 585
R710 VDD2.n145 VDD2.n144 585
R711 VDD2.n143 VDD2.n142 585
R712 VDD2.n134 VDD2.n133 585
R713 VDD2.n137 VDD2.n136 585
R714 VDD2.n33 VDD2.n32 585
R715 VDD2.n30 VDD2.n29 585
R716 VDD2.n39 VDD2.n38 585
R717 VDD2.n41 VDD2.n40 585
R718 VDD2.n26 VDD2.n25 585
R719 VDD2.n47 VDD2.n46 585
R720 VDD2.n50 VDD2.n49 585
R721 VDD2.n48 VDD2.n22 585
R722 VDD2.n55 VDD2.n21 585
R723 VDD2.n57 VDD2.n56 585
R724 VDD2.n59 VDD2.n58 585
R725 VDD2.n18 VDD2.n17 585
R726 VDD2.n65 VDD2.n64 585
R727 VDD2.n67 VDD2.n66 585
R728 VDD2.n14 VDD2.n13 585
R729 VDD2.n73 VDD2.n72 585
R730 VDD2.n75 VDD2.n74 585
R731 VDD2.n10 VDD2.n9 585
R732 VDD2.n81 VDD2.n80 585
R733 VDD2.n83 VDD2.n82 585
R734 VDD2.n6 VDD2.n5 585
R735 VDD2.n89 VDD2.n88 585
R736 VDD2.n91 VDD2.n90 585
R737 VDD2.n2 VDD2.n1 585
R738 VDD2.n97 VDD2.n96 585
R739 VDD2.t9 VDD2.n135 329.036
R740 VDD2.t1 VDD2.n31 329.036
R741 VDD2.n200 VDD2.n104 171.744
R742 VDD2.n193 VDD2.n104 171.744
R743 VDD2.n193 VDD2.n192 171.744
R744 VDD2.n192 VDD2.n108 171.744
R745 VDD2.n185 VDD2.n108 171.744
R746 VDD2.n185 VDD2.n184 171.744
R747 VDD2.n184 VDD2.n112 171.744
R748 VDD2.n177 VDD2.n112 171.744
R749 VDD2.n177 VDD2.n176 171.744
R750 VDD2.n176 VDD2.n116 171.744
R751 VDD2.n169 VDD2.n116 171.744
R752 VDD2.n169 VDD2.n168 171.744
R753 VDD2.n168 VDD2.n120 171.744
R754 VDD2.n161 VDD2.n120 171.744
R755 VDD2.n161 VDD2.n160 171.744
R756 VDD2.n160 VDD2.n124 171.744
R757 VDD2.n128 VDD2.n124 171.744
R758 VDD2.n152 VDD2.n128 171.744
R759 VDD2.n152 VDD2.n151 171.744
R760 VDD2.n151 VDD2.n129 171.744
R761 VDD2.n144 VDD2.n129 171.744
R762 VDD2.n144 VDD2.n143 171.744
R763 VDD2.n143 VDD2.n133 171.744
R764 VDD2.n136 VDD2.n133 171.744
R765 VDD2.n32 VDD2.n29 171.744
R766 VDD2.n39 VDD2.n29 171.744
R767 VDD2.n40 VDD2.n39 171.744
R768 VDD2.n40 VDD2.n25 171.744
R769 VDD2.n47 VDD2.n25 171.744
R770 VDD2.n49 VDD2.n47 171.744
R771 VDD2.n49 VDD2.n48 171.744
R772 VDD2.n48 VDD2.n21 171.744
R773 VDD2.n57 VDD2.n21 171.744
R774 VDD2.n58 VDD2.n57 171.744
R775 VDD2.n58 VDD2.n17 171.744
R776 VDD2.n65 VDD2.n17 171.744
R777 VDD2.n66 VDD2.n65 171.744
R778 VDD2.n66 VDD2.n13 171.744
R779 VDD2.n73 VDD2.n13 171.744
R780 VDD2.n74 VDD2.n73 171.744
R781 VDD2.n74 VDD2.n9 171.744
R782 VDD2.n81 VDD2.n9 171.744
R783 VDD2.n82 VDD2.n81 171.744
R784 VDD2.n82 VDD2.n5 171.744
R785 VDD2.n89 VDD2.n5 171.744
R786 VDD2.n90 VDD2.n89 171.744
R787 VDD2.n90 VDD2.n1 171.744
R788 VDD2.n97 VDD2.n1 171.744
R789 VDD2.n136 VDD2.t9 85.8723
R790 VDD2.n32 VDD2.t1 85.8723
R791 VDD2.n102 VDD2.n101 72.0652
R792 VDD2 VDD2.n205 72.0613
R793 VDD2.n204 VDD2.n203 71.4418
R794 VDD2.n100 VDD2.n99 71.4416
R795 VDD2.n100 VDD2.n98 51.7087
R796 VDD2.n202 VDD2.n201 50.8035
R797 VDD2.n202 VDD2.n102 43.5666
R798 VDD2.n159 VDD2.n158 13.1884
R799 VDD2.n56 VDD2.n55 13.1884
R800 VDD2.n162 VDD2.n123 12.8005
R801 VDD2.n157 VDD2.n125 12.8005
R802 VDD2.n54 VDD2.n22 12.8005
R803 VDD2.n59 VDD2.n20 12.8005
R804 VDD2.n199 VDD2.n103 12.0247
R805 VDD2.n163 VDD2.n121 12.0247
R806 VDD2.n154 VDD2.n153 12.0247
R807 VDD2.n51 VDD2.n50 12.0247
R808 VDD2.n60 VDD2.n18 12.0247
R809 VDD2.n96 VDD2.n0 12.0247
R810 VDD2.n198 VDD2.n105 11.249
R811 VDD2.n167 VDD2.n166 11.249
R812 VDD2.n150 VDD2.n127 11.249
R813 VDD2.n46 VDD2.n24 11.249
R814 VDD2.n64 VDD2.n63 11.249
R815 VDD2.n95 VDD2.n2 11.249
R816 VDD2.n137 VDD2.n135 10.7239
R817 VDD2.n33 VDD2.n31 10.7239
R818 VDD2.n195 VDD2.n194 10.4732
R819 VDD2.n170 VDD2.n119 10.4732
R820 VDD2.n149 VDD2.n130 10.4732
R821 VDD2.n45 VDD2.n26 10.4732
R822 VDD2.n67 VDD2.n16 10.4732
R823 VDD2.n92 VDD2.n91 10.4732
R824 VDD2.n191 VDD2.n107 9.69747
R825 VDD2.n171 VDD2.n117 9.69747
R826 VDD2.n146 VDD2.n145 9.69747
R827 VDD2.n42 VDD2.n41 9.69747
R828 VDD2.n68 VDD2.n14 9.69747
R829 VDD2.n88 VDD2.n4 9.69747
R830 VDD2.n197 VDD2.n103 9.45567
R831 VDD2.n94 VDD2.n0 9.45567
R832 VDD2.n139 VDD2.n138 9.3005
R833 VDD2.n141 VDD2.n140 9.3005
R834 VDD2.n132 VDD2.n131 9.3005
R835 VDD2.n147 VDD2.n146 9.3005
R836 VDD2.n149 VDD2.n148 9.3005
R837 VDD2.n127 VDD2.n126 9.3005
R838 VDD2.n155 VDD2.n154 9.3005
R839 VDD2.n157 VDD2.n156 9.3005
R840 VDD2.n111 VDD2.n110 9.3005
R841 VDD2.n188 VDD2.n187 9.3005
R842 VDD2.n190 VDD2.n189 9.3005
R843 VDD2.n107 VDD2.n106 9.3005
R844 VDD2.n196 VDD2.n195 9.3005
R845 VDD2.n198 VDD2.n197 9.3005
R846 VDD2.n182 VDD2.n181 9.3005
R847 VDD2.n180 VDD2.n179 9.3005
R848 VDD2.n115 VDD2.n114 9.3005
R849 VDD2.n174 VDD2.n173 9.3005
R850 VDD2.n172 VDD2.n171 9.3005
R851 VDD2.n119 VDD2.n118 9.3005
R852 VDD2.n166 VDD2.n165 9.3005
R853 VDD2.n164 VDD2.n163 9.3005
R854 VDD2.n123 VDD2.n122 9.3005
R855 VDD2.n79 VDD2.n78 9.3005
R856 VDD2.n8 VDD2.n7 9.3005
R857 VDD2.n85 VDD2.n84 9.3005
R858 VDD2.n87 VDD2.n86 9.3005
R859 VDD2.n4 VDD2.n3 9.3005
R860 VDD2.n93 VDD2.n92 9.3005
R861 VDD2.n95 VDD2.n94 9.3005
R862 VDD2.n12 VDD2.n11 9.3005
R863 VDD2.n71 VDD2.n70 9.3005
R864 VDD2.n69 VDD2.n68 9.3005
R865 VDD2.n16 VDD2.n15 9.3005
R866 VDD2.n63 VDD2.n62 9.3005
R867 VDD2.n61 VDD2.n60 9.3005
R868 VDD2.n20 VDD2.n19 9.3005
R869 VDD2.n35 VDD2.n34 9.3005
R870 VDD2.n37 VDD2.n36 9.3005
R871 VDD2.n28 VDD2.n27 9.3005
R872 VDD2.n43 VDD2.n42 9.3005
R873 VDD2.n45 VDD2.n44 9.3005
R874 VDD2.n24 VDD2.n23 9.3005
R875 VDD2.n52 VDD2.n51 9.3005
R876 VDD2.n54 VDD2.n53 9.3005
R877 VDD2.n77 VDD2.n76 9.3005
R878 VDD2.n190 VDD2.n109 8.92171
R879 VDD2.n175 VDD2.n174 8.92171
R880 VDD2.n142 VDD2.n132 8.92171
R881 VDD2.n38 VDD2.n28 8.92171
R882 VDD2.n72 VDD2.n71 8.92171
R883 VDD2.n87 VDD2.n6 8.92171
R884 VDD2.n187 VDD2.n186 8.14595
R885 VDD2.n178 VDD2.n115 8.14595
R886 VDD2.n141 VDD2.n134 8.14595
R887 VDD2.n37 VDD2.n30 8.14595
R888 VDD2.n75 VDD2.n12 8.14595
R889 VDD2.n84 VDD2.n83 8.14595
R890 VDD2.n183 VDD2.n111 7.3702
R891 VDD2.n179 VDD2.n113 7.3702
R892 VDD2.n138 VDD2.n137 7.3702
R893 VDD2.n34 VDD2.n33 7.3702
R894 VDD2.n76 VDD2.n10 7.3702
R895 VDD2.n80 VDD2.n8 7.3702
R896 VDD2.n183 VDD2.n182 6.59444
R897 VDD2.n182 VDD2.n113 6.59444
R898 VDD2.n79 VDD2.n10 6.59444
R899 VDD2.n80 VDD2.n79 6.59444
R900 VDD2.n186 VDD2.n111 5.81868
R901 VDD2.n179 VDD2.n178 5.81868
R902 VDD2.n138 VDD2.n134 5.81868
R903 VDD2.n34 VDD2.n30 5.81868
R904 VDD2.n76 VDD2.n75 5.81868
R905 VDD2.n83 VDD2.n8 5.81868
R906 VDD2.n187 VDD2.n109 5.04292
R907 VDD2.n175 VDD2.n115 5.04292
R908 VDD2.n142 VDD2.n141 5.04292
R909 VDD2.n38 VDD2.n37 5.04292
R910 VDD2.n72 VDD2.n12 5.04292
R911 VDD2.n84 VDD2.n6 5.04292
R912 VDD2.n191 VDD2.n190 4.26717
R913 VDD2.n174 VDD2.n117 4.26717
R914 VDD2.n145 VDD2.n132 4.26717
R915 VDD2.n41 VDD2.n28 4.26717
R916 VDD2.n71 VDD2.n14 4.26717
R917 VDD2.n88 VDD2.n87 4.26717
R918 VDD2.n194 VDD2.n107 3.49141
R919 VDD2.n171 VDD2.n170 3.49141
R920 VDD2.n146 VDD2.n130 3.49141
R921 VDD2.n42 VDD2.n26 3.49141
R922 VDD2.n68 VDD2.n67 3.49141
R923 VDD2.n91 VDD2.n4 3.49141
R924 VDD2.n195 VDD2.n105 2.71565
R925 VDD2.n167 VDD2.n119 2.71565
R926 VDD2.n150 VDD2.n149 2.71565
R927 VDD2.n46 VDD2.n45 2.71565
R928 VDD2.n64 VDD2.n16 2.71565
R929 VDD2.n92 VDD2.n2 2.71565
R930 VDD2.n139 VDD2.n135 2.41282
R931 VDD2.n35 VDD2.n31 2.41282
R932 VDD2.n199 VDD2.n198 1.93989
R933 VDD2.n166 VDD2.n121 1.93989
R934 VDD2.n153 VDD2.n127 1.93989
R935 VDD2.n50 VDD2.n24 1.93989
R936 VDD2.n63 VDD2.n18 1.93989
R937 VDD2.n96 VDD2.n95 1.93989
R938 VDD2.n205 VDD2.t4 1.80233
R939 VDD2.n205 VDD2.t7 1.80233
R940 VDD2.n203 VDD2.t2 1.80233
R941 VDD2.n203 VDD2.t3 1.80233
R942 VDD2.n101 VDD2.t0 1.80233
R943 VDD2.n101 VDD2.t5 1.80233
R944 VDD2.n99 VDD2.t6 1.80233
R945 VDD2.n99 VDD2.t8 1.80233
R946 VDD2.n201 VDD2.n103 1.16414
R947 VDD2.n163 VDD2.n162 1.16414
R948 VDD2.n154 VDD2.n125 1.16414
R949 VDD2.n51 VDD2.n22 1.16414
R950 VDD2.n60 VDD2.n59 1.16414
R951 VDD2.n98 VDD2.n0 1.16414
R952 VDD2.n204 VDD2.n202 0.905672
R953 VDD2.n159 VDD2.n123 0.388379
R954 VDD2.n158 VDD2.n157 0.388379
R955 VDD2.n55 VDD2.n54 0.388379
R956 VDD2.n56 VDD2.n20 0.388379
R957 VDD2 VDD2.n204 0.284983
R958 VDD2.n102 VDD2.n100 0.171447
R959 VDD2.n197 VDD2.n196 0.155672
R960 VDD2.n196 VDD2.n106 0.155672
R961 VDD2.n189 VDD2.n106 0.155672
R962 VDD2.n189 VDD2.n188 0.155672
R963 VDD2.n188 VDD2.n110 0.155672
R964 VDD2.n181 VDD2.n110 0.155672
R965 VDD2.n181 VDD2.n180 0.155672
R966 VDD2.n180 VDD2.n114 0.155672
R967 VDD2.n173 VDD2.n114 0.155672
R968 VDD2.n173 VDD2.n172 0.155672
R969 VDD2.n172 VDD2.n118 0.155672
R970 VDD2.n165 VDD2.n118 0.155672
R971 VDD2.n165 VDD2.n164 0.155672
R972 VDD2.n164 VDD2.n122 0.155672
R973 VDD2.n156 VDD2.n122 0.155672
R974 VDD2.n156 VDD2.n155 0.155672
R975 VDD2.n155 VDD2.n126 0.155672
R976 VDD2.n148 VDD2.n126 0.155672
R977 VDD2.n148 VDD2.n147 0.155672
R978 VDD2.n147 VDD2.n131 0.155672
R979 VDD2.n140 VDD2.n131 0.155672
R980 VDD2.n140 VDD2.n139 0.155672
R981 VDD2.n36 VDD2.n35 0.155672
R982 VDD2.n36 VDD2.n27 0.155672
R983 VDD2.n43 VDD2.n27 0.155672
R984 VDD2.n44 VDD2.n43 0.155672
R985 VDD2.n44 VDD2.n23 0.155672
R986 VDD2.n52 VDD2.n23 0.155672
R987 VDD2.n53 VDD2.n52 0.155672
R988 VDD2.n53 VDD2.n19 0.155672
R989 VDD2.n61 VDD2.n19 0.155672
R990 VDD2.n62 VDD2.n61 0.155672
R991 VDD2.n62 VDD2.n15 0.155672
R992 VDD2.n69 VDD2.n15 0.155672
R993 VDD2.n70 VDD2.n69 0.155672
R994 VDD2.n70 VDD2.n11 0.155672
R995 VDD2.n77 VDD2.n11 0.155672
R996 VDD2.n78 VDD2.n77 0.155672
R997 VDD2.n78 VDD2.n7 0.155672
R998 VDD2.n85 VDD2.n7 0.155672
R999 VDD2.n86 VDD2.n85 0.155672
R1000 VDD2.n86 VDD2.n3 0.155672
R1001 VDD2.n93 VDD2.n3 0.155672
R1002 VDD2.n94 VDD2.n93 0.155672
R1003 B.n314 B.t6 806.566
R1004 B.n141 B.t0 806.566
R1005 B.n53 B.t3 806.566
R1006 B.n46 B.t9 806.566
R1007 B.n422 B.n111 585
R1008 B.n421 B.n420 585
R1009 B.n419 B.n112 585
R1010 B.n418 B.n417 585
R1011 B.n416 B.n113 585
R1012 B.n415 B.n414 585
R1013 B.n413 B.n114 585
R1014 B.n412 B.n411 585
R1015 B.n410 B.n115 585
R1016 B.n409 B.n408 585
R1017 B.n407 B.n116 585
R1018 B.n406 B.n405 585
R1019 B.n404 B.n117 585
R1020 B.n403 B.n402 585
R1021 B.n401 B.n118 585
R1022 B.n400 B.n399 585
R1023 B.n398 B.n119 585
R1024 B.n397 B.n396 585
R1025 B.n395 B.n120 585
R1026 B.n394 B.n393 585
R1027 B.n392 B.n121 585
R1028 B.n391 B.n390 585
R1029 B.n389 B.n122 585
R1030 B.n388 B.n387 585
R1031 B.n386 B.n123 585
R1032 B.n385 B.n384 585
R1033 B.n383 B.n124 585
R1034 B.n382 B.n381 585
R1035 B.n380 B.n125 585
R1036 B.n379 B.n378 585
R1037 B.n377 B.n126 585
R1038 B.n376 B.n375 585
R1039 B.n374 B.n127 585
R1040 B.n373 B.n372 585
R1041 B.n371 B.n128 585
R1042 B.n370 B.n369 585
R1043 B.n368 B.n129 585
R1044 B.n367 B.n366 585
R1045 B.n365 B.n130 585
R1046 B.n364 B.n363 585
R1047 B.n362 B.n131 585
R1048 B.n361 B.n360 585
R1049 B.n359 B.n132 585
R1050 B.n358 B.n357 585
R1051 B.n356 B.n133 585
R1052 B.n355 B.n354 585
R1053 B.n353 B.n134 585
R1054 B.n352 B.n351 585
R1055 B.n350 B.n135 585
R1056 B.n349 B.n348 585
R1057 B.n347 B.n136 585
R1058 B.n346 B.n345 585
R1059 B.n344 B.n137 585
R1060 B.n343 B.n342 585
R1061 B.n341 B.n138 585
R1062 B.n340 B.n339 585
R1063 B.n338 B.n139 585
R1064 B.n337 B.n336 585
R1065 B.n335 B.n140 585
R1066 B.n333 B.n332 585
R1067 B.n331 B.n143 585
R1068 B.n330 B.n329 585
R1069 B.n328 B.n144 585
R1070 B.n327 B.n326 585
R1071 B.n325 B.n145 585
R1072 B.n324 B.n323 585
R1073 B.n322 B.n146 585
R1074 B.n321 B.n320 585
R1075 B.n319 B.n147 585
R1076 B.n318 B.n317 585
R1077 B.n313 B.n148 585
R1078 B.n312 B.n311 585
R1079 B.n310 B.n149 585
R1080 B.n309 B.n308 585
R1081 B.n307 B.n150 585
R1082 B.n306 B.n305 585
R1083 B.n304 B.n151 585
R1084 B.n303 B.n302 585
R1085 B.n301 B.n152 585
R1086 B.n300 B.n299 585
R1087 B.n298 B.n153 585
R1088 B.n297 B.n296 585
R1089 B.n295 B.n154 585
R1090 B.n294 B.n293 585
R1091 B.n292 B.n155 585
R1092 B.n291 B.n290 585
R1093 B.n289 B.n156 585
R1094 B.n288 B.n287 585
R1095 B.n286 B.n157 585
R1096 B.n285 B.n284 585
R1097 B.n283 B.n158 585
R1098 B.n282 B.n281 585
R1099 B.n280 B.n159 585
R1100 B.n279 B.n278 585
R1101 B.n277 B.n160 585
R1102 B.n276 B.n275 585
R1103 B.n274 B.n161 585
R1104 B.n273 B.n272 585
R1105 B.n271 B.n162 585
R1106 B.n270 B.n269 585
R1107 B.n268 B.n163 585
R1108 B.n267 B.n266 585
R1109 B.n265 B.n164 585
R1110 B.n264 B.n263 585
R1111 B.n262 B.n165 585
R1112 B.n261 B.n260 585
R1113 B.n259 B.n166 585
R1114 B.n258 B.n257 585
R1115 B.n256 B.n167 585
R1116 B.n255 B.n254 585
R1117 B.n253 B.n168 585
R1118 B.n252 B.n251 585
R1119 B.n250 B.n169 585
R1120 B.n249 B.n248 585
R1121 B.n247 B.n170 585
R1122 B.n246 B.n245 585
R1123 B.n244 B.n171 585
R1124 B.n243 B.n242 585
R1125 B.n241 B.n172 585
R1126 B.n240 B.n239 585
R1127 B.n238 B.n173 585
R1128 B.n237 B.n236 585
R1129 B.n235 B.n174 585
R1130 B.n234 B.n233 585
R1131 B.n232 B.n175 585
R1132 B.n231 B.n230 585
R1133 B.n229 B.n176 585
R1134 B.n228 B.n227 585
R1135 B.n424 B.n423 585
R1136 B.n425 B.n110 585
R1137 B.n427 B.n426 585
R1138 B.n428 B.n109 585
R1139 B.n430 B.n429 585
R1140 B.n431 B.n108 585
R1141 B.n433 B.n432 585
R1142 B.n434 B.n107 585
R1143 B.n436 B.n435 585
R1144 B.n437 B.n106 585
R1145 B.n439 B.n438 585
R1146 B.n440 B.n105 585
R1147 B.n442 B.n441 585
R1148 B.n443 B.n104 585
R1149 B.n445 B.n444 585
R1150 B.n446 B.n103 585
R1151 B.n448 B.n447 585
R1152 B.n449 B.n102 585
R1153 B.n451 B.n450 585
R1154 B.n452 B.n101 585
R1155 B.n454 B.n453 585
R1156 B.n455 B.n100 585
R1157 B.n457 B.n456 585
R1158 B.n458 B.n99 585
R1159 B.n460 B.n459 585
R1160 B.n461 B.n98 585
R1161 B.n463 B.n462 585
R1162 B.n464 B.n97 585
R1163 B.n466 B.n465 585
R1164 B.n467 B.n96 585
R1165 B.n469 B.n468 585
R1166 B.n470 B.n95 585
R1167 B.n472 B.n471 585
R1168 B.n473 B.n94 585
R1169 B.n475 B.n474 585
R1170 B.n476 B.n93 585
R1171 B.n478 B.n477 585
R1172 B.n479 B.n92 585
R1173 B.n481 B.n480 585
R1174 B.n482 B.n91 585
R1175 B.n484 B.n483 585
R1176 B.n485 B.n90 585
R1177 B.n487 B.n486 585
R1178 B.n488 B.n89 585
R1179 B.n490 B.n489 585
R1180 B.n491 B.n88 585
R1181 B.n493 B.n492 585
R1182 B.n494 B.n87 585
R1183 B.n496 B.n495 585
R1184 B.n497 B.n86 585
R1185 B.n499 B.n498 585
R1186 B.n500 B.n85 585
R1187 B.n502 B.n501 585
R1188 B.n503 B.n84 585
R1189 B.n696 B.n15 585
R1190 B.n695 B.n694 585
R1191 B.n693 B.n16 585
R1192 B.n692 B.n691 585
R1193 B.n690 B.n17 585
R1194 B.n689 B.n688 585
R1195 B.n687 B.n18 585
R1196 B.n686 B.n685 585
R1197 B.n684 B.n19 585
R1198 B.n683 B.n682 585
R1199 B.n681 B.n20 585
R1200 B.n680 B.n679 585
R1201 B.n678 B.n21 585
R1202 B.n677 B.n676 585
R1203 B.n675 B.n22 585
R1204 B.n674 B.n673 585
R1205 B.n672 B.n23 585
R1206 B.n671 B.n670 585
R1207 B.n669 B.n24 585
R1208 B.n668 B.n667 585
R1209 B.n666 B.n25 585
R1210 B.n665 B.n664 585
R1211 B.n663 B.n26 585
R1212 B.n662 B.n661 585
R1213 B.n660 B.n27 585
R1214 B.n659 B.n658 585
R1215 B.n657 B.n28 585
R1216 B.n656 B.n655 585
R1217 B.n654 B.n29 585
R1218 B.n653 B.n652 585
R1219 B.n651 B.n30 585
R1220 B.n650 B.n649 585
R1221 B.n648 B.n31 585
R1222 B.n647 B.n646 585
R1223 B.n645 B.n32 585
R1224 B.n644 B.n643 585
R1225 B.n642 B.n33 585
R1226 B.n641 B.n640 585
R1227 B.n639 B.n34 585
R1228 B.n638 B.n637 585
R1229 B.n636 B.n35 585
R1230 B.n635 B.n634 585
R1231 B.n633 B.n36 585
R1232 B.n632 B.n631 585
R1233 B.n630 B.n37 585
R1234 B.n629 B.n628 585
R1235 B.n627 B.n38 585
R1236 B.n626 B.n625 585
R1237 B.n624 B.n39 585
R1238 B.n623 B.n622 585
R1239 B.n621 B.n40 585
R1240 B.n620 B.n619 585
R1241 B.n618 B.n41 585
R1242 B.n617 B.n616 585
R1243 B.n615 B.n42 585
R1244 B.n614 B.n613 585
R1245 B.n612 B.n43 585
R1246 B.n611 B.n610 585
R1247 B.n609 B.n44 585
R1248 B.n608 B.n607 585
R1249 B.n606 B.n45 585
R1250 B.n605 B.n604 585
R1251 B.n603 B.n49 585
R1252 B.n602 B.n601 585
R1253 B.n600 B.n50 585
R1254 B.n599 B.n598 585
R1255 B.n597 B.n51 585
R1256 B.n596 B.n595 585
R1257 B.n594 B.n52 585
R1258 B.n592 B.n591 585
R1259 B.n590 B.n55 585
R1260 B.n589 B.n588 585
R1261 B.n587 B.n56 585
R1262 B.n586 B.n585 585
R1263 B.n584 B.n57 585
R1264 B.n583 B.n582 585
R1265 B.n581 B.n58 585
R1266 B.n580 B.n579 585
R1267 B.n578 B.n59 585
R1268 B.n577 B.n576 585
R1269 B.n575 B.n60 585
R1270 B.n574 B.n573 585
R1271 B.n572 B.n61 585
R1272 B.n571 B.n570 585
R1273 B.n569 B.n62 585
R1274 B.n568 B.n567 585
R1275 B.n566 B.n63 585
R1276 B.n565 B.n564 585
R1277 B.n563 B.n64 585
R1278 B.n562 B.n561 585
R1279 B.n560 B.n65 585
R1280 B.n559 B.n558 585
R1281 B.n557 B.n66 585
R1282 B.n556 B.n555 585
R1283 B.n554 B.n67 585
R1284 B.n553 B.n552 585
R1285 B.n551 B.n68 585
R1286 B.n550 B.n549 585
R1287 B.n548 B.n69 585
R1288 B.n547 B.n546 585
R1289 B.n545 B.n70 585
R1290 B.n544 B.n543 585
R1291 B.n542 B.n71 585
R1292 B.n541 B.n540 585
R1293 B.n539 B.n72 585
R1294 B.n538 B.n537 585
R1295 B.n536 B.n73 585
R1296 B.n535 B.n534 585
R1297 B.n533 B.n74 585
R1298 B.n532 B.n531 585
R1299 B.n530 B.n75 585
R1300 B.n529 B.n528 585
R1301 B.n527 B.n76 585
R1302 B.n526 B.n525 585
R1303 B.n524 B.n77 585
R1304 B.n523 B.n522 585
R1305 B.n521 B.n78 585
R1306 B.n520 B.n519 585
R1307 B.n518 B.n79 585
R1308 B.n517 B.n516 585
R1309 B.n515 B.n80 585
R1310 B.n514 B.n513 585
R1311 B.n512 B.n81 585
R1312 B.n511 B.n510 585
R1313 B.n509 B.n82 585
R1314 B.n508 B.n507 585
R1315 B.n506 B.n83 585
R1316 B.n505 B.n504 585
R1317 B.n698 B.n697 585
R1318 B.n699 B.n14 585
R1319 B.n701 B.n700 585
R1320 B.n702 B.n13 585
R1321 B.n704 B.n703 585
R1322 B.n705 B.n12 585
R1323 B.n707 B.n706 585
R1324 B.n708 B.n11 585
R1325 B.n710 B.n709 585
R1326 B.n711 B.n10 585
R1327 B.n713 B.n712 585
R1328 B.n714 B.n9 585
R1329 B.n716 B.n715 585
R1330 B.n717 B.n8 585
R1331 B.n719 B.n718 585
R1332 B.n720 B.n7 585
R1333 B.n722 B.n721 585
R1334 B.n723 B.n6 585
R1335 B.n725 B.n724 585
R1336 B.n726 B.n5 585
R1337 B.n728 B.n727 585
R1338 B.n729 B.n4 585
R1339 B.n731 B.n730 585
R1340 B.n732 B.n3 585
R1341 B.n734 B.n733 585
R1342 B.n735 B.n0 585
R1343 B.n2 B.n1 585
R1344 B.n190 B.n189 585
R1345 B.n192 B.n191 585
R1346 B.n193 B.n188 585
R1347 B.n195 B.n194 585
R1348 B.n196 B.n187 585
R1349 B.n198 B.n197 585
R1350 B.n199 B.n186 585
R1351 B.n201 B.n200 585
R1352 B.n202 B.n185 585
R1353 B.n204 B.n203 585
R1354 B.n205 B.n184 585
R1355 B.n207 B.n206 585
R1356 B.n208 B.n183 585
R1357 B.n210 B.n209 585
R1358 B.n211 B.n182 585
R1359 B.n213 B.n212 585
R1360 B.n214 B.n181 585
R1361 B.n216 B.n215 585
R1362 B.n217 B.n180 585
R1363 B.n219 B.n218 585
R1364 B.n220 B.n179 585
R1365 B.n222 B.n221 585
R1366 B.n223 B.n178 585
R1367 B.n225 B.n224 585
R1368 B.n226 B.n177 585
R1369 B.n227 B.n226 550.159
R1370 B.n423 B.n422 550.159
R1371 B.n505 B.n84 550.159
R1372 B.n698 B.n15 550.159
R1373 B.n141 B.t1 504.574
R1374 B.n53 B.t5 504.574
R1375 B.n314 B.t7 504.574
R1376 B.n46 B.t11 504.574
R1377 B.n142 B.t2 484.211
R1378 B.n54 B.t4 484.211
R1379 B.n315 B.t8 484.211
R1380 B.n47 B.t10 484.211
R1381 B.n737 B.n736 256.663
R1382 B.n736 B.n735 235.042
R1383 B.n736 B.n2 235.042
R1384 B.n227 B.n176 163.367
R1385 B.n231 B.n176 163.367
R1386 B.n232 B.n231 163.367
R1387 B.n233 B.n232 163.367
R1388 B.n233 B.n174 163.367
R1389 B.n237 B.n174 163.367
R1390 B.n238 B.n237 163.367
R1391 B.n239 B.n238 163.367
R1392 B.n239 B.n172 163.367
R1393 B.n243 B.n172 163.367
R1394 B.n244 B.n243 163.367
R1395 B.n245 B.n244 163.367
R1396 B.n245 B.n170 163.367
R1397 B.n249 B.n170 163.367
R1398 B.n250 B.n249 163.367
R1399 B.n251 B.n250 163.367
R1400 B.n251 B.n168 163.367
R1401 B.n255 B.n168 163.367
R1402 B.n256 B.n255 163.367
R1403 B.n257 B.n256 163.367
R1404 B.n257 B.n166 163.367
R1405 B.n261 B.n166 163.367
R1406 B.n262 B.n261 163.367
R1407 B.n263 B.n262 163.367
R1408 B.n263 B.n164 163.367
R1409 B.n267 B.n164 163.367
R1410 B.n268 B.n267 163.367
R1411 B.n269 B.n268 163.367
R1412 B.n269 B.n162 163.367
R1413 B.n273 B.n162 163.367
R1414 B.n274 B.n273 163.367
R1415 B.n275 B.n274 163.367
R1416 B.n275 B.n160 163.367
R1417 B.n279 B.n160 163.367
R1418 B.n280 B.n279 163.367
R1419 B.n281 B.n280 163.367
R1420 B.n281 B.n158 163.367
R1421 B.n285 B.n158 163.367
R1422 B.n286 B.n285 163.367
R1423 B.n287 B.n286 163.367
R1424 B.n287 B.n156 163.367
R1425 B.n291 B.n156 163.367
R1426 B.n292 B.n291 163.367
R1427 B.n293 B.n292 163.367
R1428 B.n293 B.n154 163.367
R1429 B.n297 B.n154 163.367
R1430 B.n298 B.n297 163.367
R1431 B.n299 B.n298 163.367
R1432 B.n299 B.n152 163.367
R1433 B.n303 B.n152 163.367
R1434 B.n304 B.n303 163.367
R1435 B.n305 B.n304 163.367
R1436 B.n305 B.n150 163.367
R1437 B.n309 B.n150 163.367
R1438 B.n310 B.n309 163.367
R1439 B.n311 B.n310 163.367
R1440 B.n311 B.n148 163.367
R1441 B.n318 B.n148 163.367
R1442 B.n319 B.n318 163.367
R1443 B.n320 B.n319 163.367
R1444 B.n320 B.n146 163.367
R1445 B.n324 B.n146 163.367
R1446 B.n325 B.n324 163.367
R1447 B.n326 B.n325 163.367
R1448 B.n326 B.n144 163.367
R1449 B.n330 B.n144 163.367
R1450 B.n331 B.n330 163.367
R1451 B.n332 B.n331 163.367
R1452 B.n332 B.n140 163.367
R1453 B.n337 B.n140 163.367
R1454 B.n338 B.n337 163.367
R1455 B.n339 B.n338 163.367
R1456 B.n339 B.n138 163.367
R1457 B.n343 B.n138 163.367
R1458 B.n344 B.n343 163.367
R1459 B.n345 B.n344 163.367
R1460 B.n345 B.n136 163.367
R1461 B.n349 B.n136 163.367
R1462 B.n350 B.n349 163.367
R1463 B.n351 B.n350 163.367
R1464 B.n351 B.n134 163.367
R1465 B.n355 B.n134 163.367
R1466 B.n356 B.n355 163.367
R1467 B.n357 B.n356 163.367
R1468 B.n357 B.n132 163.367
R1469 B.n361 B.n132 163.367
R1470 B.n362 B.n361 163.367
R1471 B.n363 B.n362 163.367
R1472 B.n363 B.n130 163.367
R1473 B.n367 B.n130 163.367
R1474 B.n368 B.n367 163.367
R1475 B.n369 B.n368 163.367
R1476 B.n369 B.n128 163.367
R1477 B.n373 B.n128 163.367
R1478 B.n374 B.n373 163.367
R1479 B.n375 B.n374 163.367
R1480 B.n375 B.n126 163.367
R1481 B.n379 B.n126 163.367
R1482 B.n380 B.n379 163.367
R1483 B.n381 B.n380 163.367
R1484 B.n381 B.n124 163.367
R1485 B.n385 B.n124 163.367
R1486 B.n386 B.n385 163.367
R1487 B.n387 B.n386 163.367
R1488 B.n387 B.n122 163.367
R1489 B.n391 B.n122 163.367
R1490 B.n392 B.n391 163.367
R1491 B.n393 B.n392 163.367
R1492 B.n393 B.n120 163.367
R1493 B.n397 B.n120 163.367
R1494 B.n398 B.n397 163.367
R1495 B.n399 B.n398 163.367
R1496 B.n399 B.n118 163.367
R1497 B.n403 B.n118 163.367
R1498 B.n404 B.n403 163.367
R1499 B.n405 B.n404 163.367
R1500 B.n405 B.n116 163.367
R1501 B.n409 B.n116 163.367
R1502 B.n410 B.n409 163.367
R1503 B.n411 B.n410 163.367
R1504 B.n411 B.n114 163.367
R1505 B.n415 B.n114 163.367
R1506 B.n416 B.n415 163.367
R1507 B.n417 B.n416 163.367
R1508 B.n417 B.n112 163.367
R1509 B.n421 B.n112 163.367
R1510 B.n422 B.n421 163.367
R1511 B.n501 B.n84 163.367
R1512 B.n501 B.n500 163.367
R1513 B.n500 B.n499 163.367
R1514 B.n499 B.n86 163.367
R1515 B.n495 B.n86 163.367
R1516 B.n495 B.n494 163.367
R1517 B.n494 B.n493 163.367
R1518 B.n493 B.n88 163.367
R1519 B.n489 B.n88 163.367
R1520 B.n489 B.n488 163.367
R1521 B.n488 B.n487 163.367
R1522 B.n487 B.n90 163.367
R1523 B.n483 B.n90 163.367
R1524 B.n483 B.n482 163.367
R1525 B.n482 B.n481 163.367
R1526 B.n481 B.n92 163.367
R1527 B.n477 B.n92 163.367
R1528 B.n477 B.n476 163.367
R1529 B.n476 B.n475 163.367
R1530 B.n475 B.n94 163.367
R1531 B.n471 B.n94 163.367
R1532 B.n471 B.n470 163.367
R1533 B.n470 B.n469 163.367
R1534 B.n469 B.n96 163.367
R1535 B.n465 B.n96 163.367
R1536 B.n465 B.n464 163.367
R1537 B.n464 B.n463 163.367
R1538 B.n463 B.n98 163.367
R1539 B.n459 B.n98 163.367
R1540 B.n459 B.n458 163.367
R1541 B.n458 B.n457 163.367
R1542 B.n457 B.n100 163.367
R1543 B.n453 B.n100 163.367
R1544 B.n453 B.n452 163.367
R1545 B.n452 B.n451 163.367
R1546 B.n451 B.n102 163.367
R1547 B.n447 B.n102 163.367
R1548 B.n447 B.n446 163.367
R1549 B.n446 B.n445 163.367
R1550 B.n445 B.n104 163.367
R1551 B.n441 B.n104 163.367
R1552 B.n441 B.n440 163.367
R1553 B.n440 B.n439 163.367
R1554 B.n439 B.n106 163.367
R1555 B.n435 B.n106 163.367
R1556 B.n435 B.n434 163.367
R1557 B.n434 B.n433 163.367
R1558 B.n433 B.n108 163.367
R1559 B.n429 B.n108 163.367
R1560 B.n429 B.n428 163.367
R1561 B.n428 B.n427 163.367
R1562 B.n427 B.n110 163.367
R1563 B.n423 B.n110 163.367
R1564 B.n694 B.n15 163.367
R1565 B.n694 B.n693 163.367
R1566 B.n693 B.n692 163.367
R1567 B.n692 B.n17 163.367
R1568 B.n688 B.n17 163.367
R1569 B.n688 B.n687 163.367
R1570 B.n687 B.n686 163.367
R1571 B.n686 B.n19 163.367
R1572 B.n682 B.n19 163.367
R1573 B.n682 B.n681 163.367
R1574 B.n681 B.n680 163.367
R1575 B.n680 B.n21 163.367
R1576 B.n676 B.n21 163.367
R1577 B.n676 B.n675 163.367
R1578 B.n675 B.n674 163.367
R1579 B.n674 B.n23 163.367
R1580 B.n670 B.n23 163.367
R1581 B.n670 B.n669 163.367
R1582 B.n669 B.n668 163.367
R1583 B.n668 B.n25 163.367
R1584 B.n664 B.n25 163.367
R1585 B.n664 B.n663 163.367
R1586 B.n663 B.n662 163.367
R1587 B.n662 B.n27 163.367
R1588 B.n658 B.n27 163.367
R1589 B.n658 B.n657 163.367
R1590 B.n657 B.n656 163.367
R1591 B.n656 B.n29 163.367
R1592 B.n652 B.n29 163.367
R1593 B.n652 B.n651 163.367
R1594 B.n651 B.n650 163.367
R1595 B.n650 B.n31 163.367
R1596 B.n646 B.n31 163.367
R1597 B.n646 B.n645 163.367
R1598 B.n645 B.n644 163.367
R1599 B.n644 B.n33 163.367
R1600 B.n640 B.n33 163.367
R1601 B.n640 B.n639 163.367
R1602 B.n639 B.n638 163.367
R1603 B.n638 B.n35 163.367
R1604 B.n634 B.n35 163.367
R1605 B.n634 B.n633 163.367
R1606 B.n633 B.n632 163.367
R1607 B.n632 B.n37 163.367
R1608 B.n628 B.n37 163.367
R1609 B.n628 B.n627 163.367
R1610 B.n627 B.n626 163.367
R1611 B.n626 B.n39 163.367
R1612 B.n622 B.n39 163.367
R1613 B.n622 B.n621 163.367
R1614 B.n621 B.n620 163.367
R1615 B.n620 B.n41 163.367
R1616 B.n616 B.n41 163.367
R1617 B.n616 B.n615 163.367
R1618 B.n615 B.n614 163.367
R1619 B.n614 B.n43 163.367
R1620 B.n610 B.n43 163.367
R1621 B.n610 B.n609 163.367
R1622 B.n609 B.n608 163.367
R1623 B.n608 B.n45 163.367
R1624 B.n604 B.n45 163.367
R1625 B.n604 B.n603 163.367
R1626 B.n603 B.n602 163.367
R1627 B.n602 B.n50 163.367
R1628 B.n598 B.n50 163.367
R1629 B.n598 B.n597 163.367
R1630 B.n597 B.n596 163.367
R1631 B.n596 B.n52 163.367
R1632 B.n591 B.n52 163.367
R1633 B.n591 B.n590 163.367
R1634 B.n590 B.n589 163.367
R1635 B.n589 B.n56 163.367
R1636 B.n585 B.n56 163.367
R1637 B.n585 B.n584 163.367
R1638 B.n584 B.n583 163.367
R1639 B.n583 B.n58 163.367
R1640 B.n579 B.n58 163.367
R1641 B.n579 B.n578 163.367
R1642 B.n578 B.n577 163.367
R1643 B.n577 B.n60 163.367
R1644 B.n573 B.n60 163.367
R1645 B.n573 B.n572 163.367
R1646 B.n572 B.n571 163.367
R1647 B.n571 B.n62 163.367
R1648 B.n567 B.n62 163.367
R1649 B.n567 B.n566 163.367
R1650 B.n566 B.n565 163.367
R1651 B.n565 B.n64 163.367
R1652 B.n561 B.n64 163.367
R1653 B.n561 B.n560 163.367
R1654 B.n560 B.n559 163.367
R1655 B.n559 B.n66 163.367
R1656 B.n555 B.n66 163.367
R1657 B.n555 B.n554 163.367
R1658 B.n554 B.n553 163.367
R1659 B.n553 B.n68 163.367
R1660 B.n549 B.n68 163.367
R1661 B.n549 B.n548 163.367
R1662 B.n548 B.n547 163.367
R1663 B.n547 B.n70 163.367
R1664 B.n543 B.n70 163.367
R1665 B.n543 B.n542 163.367
R1666 B.n542 B.n541 163.367
R1667 B.n541 B.n72 163.367
R1668 B.n537 B.n72 163.367
R1669 B.n537 B.n536 163.367
R1670 B.n536 B.n535 163.367
R1671 B.n535 B.n74 163.367
R1672 B.n531 B.n74 163.367
R1673 B.n531 B.n530 163.367
R1674 B.n530 B.n529 163.367
R1675 B.n529 B.n76 163.367
R1676 B.n525 B.n76 163.367
R1677 B.n525 B.n524 163.367
R1678 B.n524 B.n523 163.367
R1679 B.n523 B.n78 163.367
R1680 B.n519 B.n78 163.367
R1681 B.n519 B.n518 163.367
R1682 B.n518 B.n517 163.367
R1683 B.n517 B.n80 163.367
R1684 B.n513 B.n80 163.367
R1685 B.n513 B.n512 163.367
R1686 B.n512 B.n511 163.367
R1687 B.n511 B.n82 163.367
R1688 B.n507 B.n82 163.367
R1689 B.n507 B.n506 163.367
R1690 B.n506 B.n505 163.367
R1691 B.n699 B.n698 163.367
R1692 B.n700 B.n699 163.367
R1693 B.n700 B.n13 163.367
R1694 B.n704 B.n13 163.367
R1695 B.n705 B.n704 163.367
R1696 B.n706 B.n705 163.367
R1697 B.n706 B.n11 163.367
R1698 B.n710 B.n11 163.367
R1699 B.n711 B.n710 163.367
R1700 B.n712 B.n711 163.367
R1701 B.n712 B.n9 163.367
R1702 B.n716 B.n9 163.367
R1703 B.n717 B.n716 163.367
R1704 B.n718 B.n717 163.367
R1705 B.n718 B.n7 163.367
R1706 B.n722 B.n7 163.367
R1707 B.n723 B.n722 163.367
R1708 B.n724 B.n723 163.367
R1709 B.n724 B.n5 163.367
R1710 B.n728 B.n5 163.367
R1711 B.n729 B.n728 163.367
R1712 B.n730 B.n729 163.367
R1713 B.n730 B.n3 163.367
R1714 B.n734 B.n3 163.367
R1715 B.n735 B.n734 163.367
R1716 B.n190 B.n2 163.367
R1717 B.n191 B.n190 163.367
R1718 B.n191 B.n188 163.367
R1719 B.n195 B.n188 163.367
R1720 B.n196 B.n195 163.367
R1721 B.n197 B.n196 163.367
R1722 B.n197 B.n186 163.367
R1723 B.n201 B.n186 163.367
R1724 B.n202 B.n201 163.367
R1725 B.n203 B.n202 163.367
R1726 B.n203 B.n184 163.367
R1727 B.n207 B.n184 163.367
R1728 B.n208 B.n207 163.367
R1729 B.n209 B.n208 163.367
R1730 B.n209 B.n182 163.367
R1731 B.n213 B.n182 163.367
R1732 B.n214 B.n213 163.367
R1733 B.n215 B.n214 163.367
R1734 B.n215 B.n180 163.367
R1735 B.n219 B.n180 163.367
R1736 B.n220 B.n219 163.367
R1737 B.n221 B.n220 163.367
R1738 B.n221 B.n178 163.367
R1739 B.n225 B.n178 163.367
R1740 B.n226 B.n225 163.367
R1741 B.n316 B.n315 59.5399
R1742 B.n334 B.n142 59.5399
R1743 B.n593 B.n54 59.5399
R1744 B.n48 B.n47 59.5399
R1745 B.n697 B.n696 35.7468
R1746 B.n504 B.n503 35.7468
R1747 B.n228 B.n177 35.7468
R1748 B.n424 B.n111 35.7468
R1749 B.n315 B.n314 20.3641
R1750 B.n142 B.n141 20.3641
R1751 B.n54 B.n53 20.3641
R1752 B.n47 B.n46 20.3641
R1753 B B.n737 18.0485
R1754 B.n697 B.n14 10.6151
R1755 B.n701 B.n14 10.6151
R1756 B.n702 B.n701 10.6151
R1757 B.n703 B.n702 10.6151
R1758 B.n703 B.n12 10.6151
R1759 B.n707 B.n12 10.6151
R1760 B.n708 B.n707 10.6151
R1761 B.n709 B.n708 10.6151
R1762 B.n709 B.n10 10.6151
R1763 B.n713 B.n10 10.6151
R1764 B.n714 B.n713 10.6151
R1765 B.n715 B.n714 10.6151
R1766 B.n715 B.n8 10.6151
R1767 B.n719 B.n8 10.6151
R1768 B.n720 B.n719 10.6151
R1769 B.n721 B.n720 10.6151
R1770 B.n721 B.n6 10.6151
R1771 B.n725 B.n6 10.6151
R1772 B.n726 B.n725 10.6151
R1773 B.n727 B.n726 10.6151
R1774 B.n727 B.n4 10.6151
R1775 B.n731 B.n4 10.6151
R1776 B.n732 B.n731 10.6151
R1777 B.n733 B.n732 10.6151
R1778 B.n733 B.n0 10.6151
R1779 B.n696 B.n695 10.6151
R1780 B.n695 B.n16 10.6151
R1781 B.n691 B.n16 10.6151
R1782 B.n691 B.n690 10.6151
R1783 B.n690 B.n689 10.6151
R1784 B.n689 B.n18 10.6151
R1785 B.n685 B.n18 10.6151
R1786 B.n685 B.n684 10.6151
R1787 B.n684 B.n683 10.6151
R1788 B.n683 B.n20 10.6151
R1789 B.n679 B.n20 10.6151
R1790 B.n679 B.n678 10.6151
R1791 B.n678 B.n677 10.6151
R1792 B.n677 B.n22 10.6151
R1793 B.n673 B.n22 10.6151
R1794 B.n673 B.n672 10.6151
R1795 B.n672 B.n671 10.6151
R1796 B.n671 B.n24 10.6151
R1797 B.n667 B.n24 10.6151
R1798 B.n667 B.n666 10.6151
R1799 B.n666 B.n665 10.6151
R1800 B.n665 B.n26 10.6151
R1801 B.n661 B.n26 10.6151
R1802 B.n661 B.n660 10.6151
R1803 B.n660 B.n659 10.6151
R1804 B.n659 B.n28 10.6151
R1805 B.n655 B.n28 10.6151
R1806 B.n655 B.n654 10.6151
R1807 B.n654 B.n653 10.6151
R1808 B.n653 B.n30 10.6151
R1809 B.n649 B.n30 10.6151
R1810 B.n649 B.n648 10.6151
R1811 B.n648 B.n647 10.6151
R1812 B.n647 B.n32 10.6151
R1813 B.n643 B.n32 10.6151
R1814 B.n643 B.n642 10.6151
R1815 B.n642 B.n641 10.6151
R1816 B.n641 B.n34 10.6151
R1817 B.n637 B.n34 10.6151
R1818 B.n637 B.n636 10.6151
R1819 B.n636 B.n635 10.6151
R1820 B.n635 B.n36 10.6151
R1821 B.n631 B.n36 10.6151
R1822 B.n631 B.n630 10.6151
R1823 B.n630 B.n629 10.6151
R1824 B.n629 B.n38 10.6151
R1825 B.n625 B.n38 10.6151
R1826 B.n625 B.n624 10.6151
R1827 B.n624 B.n623 10.6151
R1828 B.n623 B.n40 10.6151
R1829 B.n619 B.n40 10.6151
R1830 B.n619 B.n618 10.6151
R1831 B.n618 B.n617 10.6151
R1832 B.n617 B.n42 10.6151
R1833 B.n613 B.n42 10.6151
R1834 B.n613 B.n612 10.6151
R1835 B.n612 B.n611 10.6151
R1836 B.n611 B.n44 10.6151
R1837 B.n607 B.n606 10.6151
R1838 B.n606 B.n605 10.6151
R1839 B.n605 B.n49 10.6151
R1840 B.n601 B.n49 10.6151
R1841 B.n601 B.n600 10.6151
R1842 B.n600 B.n599 10.6151
R1843 B.n599 B.n51 10.6151
R1844 B.n595 B.n51 10.6151
R1845 B.n595 B.n594 10.6151
R1846 B.n592 B.n55 10.6151
R1847 B.n588 B.n55 10.6151
R1848 B.n588 B.n587 10.6151
R1849 B.n587 B.n586 10.6151
R1850 B.n586 B.n57 10.6151
R1851 B.n582 B.n57 10.6151
R1852 B.n582 B.n581 10.6151
R1853 B.n581 B.n580 10.6151
R1854 B.n580 B.n59 10.6151
R1855 B.n576 B.n59 10.6151
R1856 B.n576 B.n575 10.6151
R1857 B.n575 B.n574 10.6151
R1858 B.n574 B.n61 10.6151
R1859 B.n570 B.n61 10.6151
R1860 B.n570 B.n569 10.6151
R1861 B.n569 B.n568 10.6151
R1862 B.n568 B.n63 10.6151
R1863 B.n564 B.n63 10.6151
R1864 B.n564 B.n563 10.6151
R1865 B.n563 B.n562 10.6151
R1866 B.n562 B.n65 10.6151
R1867 B.n558 B.n65 10.6151
R1868 B.n558 B.n557 10.6151
R1869 B.n557 B.n556 10.6151
R1870 B.n556 B.n67 10.6151
R1871 B.n552 B.n67 10.6151
R1872 B.n552 B.n551 10.6151
R1873 B.n551 B.n550 10.6151
R1874 B.n550 B.n69 10.6151
R1875 B.n546 B.n69 10.6151
R1876 B.n546 B.n545 10.6151
R1877 B.n545 B.n544 10.6151
R1878 B.n544 B.n71 10.6151
R1879 B.n540 B.n71 10.6151
R1880 B.n540 B.n539 10.6151
R1881 B.n539 B.n538 10.6151
R1882 B.n538 B.n73 10.6151
R1883 B.n534 B.n73 10.6151
R1884 B.n534 B.n533 10.6151
R1885 B.n533 B.n532 10.6151
R1886 B.n532 B.n75 10.6151
R1887 B.n528 B.n75 10.6151
R1888 B.n528 B.n527 10.6151
R1889 B.n527 B.n526 10.6151
R1890 B.n526 B.n77 10.6151
R1891 B.n522 B.n77 10.6151
R1892 B.n522 B.n521 10.6151
R1893 B.n521 B.n520 10.6151
R1894 B.n520 B.n79 10.6151
R1895 B.n516 B.n79 10.6151
R1896 B.n516 B.n515 10.6151
R1897 B.n515 B.n514 10.6151
R1898 B.n514 B.n81 10.6151
R1899 B.n510 B.n81 10.6151
R1900 B.n510 B.n509 10.6151
R1901 B.n509 B.n508 10.6151
R1902 B.n508 B.n83 10.6151
R1903 B.n504 B.n83 10.6151
R1904 B.n503 B.n502 10.6151
R1905 B.n502 B.n85 10.6151
R1906 B.n498 B.n85 10.6151
R1907 B.n498 B.n497 10.6151
R1908 B.n497 B.n496 10.6151
R1909 B.n496 B.n87 10.6151
R1910 B.n492 B.n87 10.6151
R1911 B.n492 B.n491 10.6151
R1912 B.n491 B.n490 10.6151
R1913 B.n490 B.n89 10.6151
R1914 B.n486 B.n89 10.6151
R1915 B.n486 B.n485 10.6151
R1916 B.n485 B.n484 10.6151
R1917 B.n484 B.n91 10.6151
R1918 B.n480 B.n91 10.6151
R1919 B.n480 B.n479 10.6151
R1920 B.n479 B.n478 10.6151
R1921 B.n478 B.n93 10.6151
R1922 B.n474 B.n93 10.6151
R1923 B.n474 B.n473 10.6151
R1924 B.n473 B.n472 10.6151
R1925 B.n472 B.n95 10.6151
R1926 B.n468 B.n95 10.6151
R1927 B.n468 B.n467 10.6151
R1928 B.n467 B.n466 10.6151
R1929 B.n466 B.n97 10.6151
R1930 B.n462 B.n97 10.6151
R1931 B.n462 B.n461 10.6151
R1932 B.n461 B.n460 10.6151
R1933 B.n460 B.n99 10.6151
R1934 B.n456 B.n99 10.6151
R1935 B.n456 B.n455 10.6151
R1936 B.n455 B.n454 10.6151
R1937 B.n454 B.n101 10.6151
R1938 B.n450 B.n101 10.6151
R1939 B.n450 B.n449 10.6151
R1940 B.n449 B.n448 10.6151
R1941 B.n448 B.n103 10.6151
R1942 B.n444 B.n103 10.6151
R1943 B.n444 B.n443 10.6151
R1944 B.n443 B.n442 10.6151
R1945 B.n442 B.n105 10.6151
R1946 B.n438 B.n105 10.6151
R1947 B.n438 B.n437 10.6151
R1948 B.n437 B.n436 10.6151
R1949 B.n436 B.n107 10.6151
R1950 B.n432 B.n107 10.6151
R1951 B.n432 B.n431 10.6151
R1952 B.n431 B.n430 10.6151
R1953 B.n430 B.n109 10.6151
R1954 B.n426 B.n109 10.6151
R1955 B.n426 B.n425 10.6151
R1956 B.n425 B.n424 10.6151
R1957 B.n189 B.n1 10.6151
R1958 B.n192 B.n189 10.6151
R1959 B.n193 B.n192 10.6151
R1960 B.n194 B.n193 10.6151
R1961 B.n194 B.n187 10.6151
R1962 B.n198 B.n187 10.6151
R1963 B.n199 B.n198 10.6151
R1964 B.n200 B.n199 10.6151
R1965 B.n200 B.n185 10.6151
R1966 B.n204 B.n185 10.6151
R1967 B.n205 B.n204 10.6151
R1968 B.n206 B.n205 10.6151
R1969 B.n206 B.n183 10.6151
R1970 B.n210 B.n183 10.6151
R1971 B.n211 B.n210 10.6151
R1972 B.n212 B.n211 10.6151
R1973 B.n212 B.n181 10.6151
R1974 B.n216 B.n181 10.6151
R1975 B.n217 B.n216 10.6151
R1976 B.n218 B.n217 10.6151
R1977 B.n218 B.n179 10.6151
R1978 B.n222 B.n179 10.6151
R1979 B.n223 B.n222 10.6151
R1980 B.n224 B.n223 10.6151
R1981 B.n224 B.n177 10.6151
R1982 B.n229 B.n228 10.6151
R1983 B.n230 B.n229 10.6151
R1984 B.n230 B.n175 10.6151
R1985 B.n234 B.n175 10.6151
R1986 B.n235 B.n234 10.6151
R1987 B.n236 B.n235 10.6151
R1988 B.n236 B.n173 10.6151
R1989 B.n240 B.n173 10.6151
R1990 B.n241 B.n240 10.6151
R1991 B.n242 B.n241 10.6151
R1992 B.n242 B.n171 10.6151
R1993 B.n246 B.n171 10.6151
R1994 B.n247 B.n246 10.6151
R1995 B.n248 B.n247 10.6151
R1996 B.n248 B.n169 10.6151
R1997 B.n252 B.n169 10.6151
R1998 B.n253 B.n252 10.6151
R1999 B.n254 B.n253 10.6151
R2000 B.n254 B.n167 10.6151
R2001 B.n258 B.n167 10.6151
R2002 B.n259 B.n258 10.6151
R2003 B.n260 B.n259 10.6151
R2004 B.n260 B.n165 10.6151
R2005 B.n264 B.n165 10.6151
R2006 B.n265 B.n264 10.6151
R2007 B.n266 B.n265 10.6151
R2008 B.n266 B.n163 10.6151
R2009 B.n270 B.n163 10.6151
R2010 B.n271 B.n270 10.6151
R2011 B.n272 B.n271 10.6151
R2012 B.n272 B.n161 10.6151
R2013 B.n276 B.n161 10.6151
R2014 B.n277 B.n276 10.6151
R2015 B.n278 B.n277 10.6151
R2016 B.n278 B.n159 10.6151
R2017 B.n282 B.n159 10.6151
R2018 B.n283 B.n282 10.6151
R2019 B.n284 B.n283 10.6151
R2020 B.n284 B.n157 10.6151
R2021 B.n288 B.n157 10.6151
R2022 B.n289 B.n288 10.6151
R2023 B.n290 B.n289 10.6151
R2024 B.n290 B.n155 10.6151
R2025 B.n294 B.n155 10.6151
R2026 B.n295 B.n294 10.6151
R2027 B.n296 B.n295 10.6151
R2028 B.n296 B.n153 10.6151
R2029 B.n300 B.n153 10.6151
R2030 B.n301 B.n300 10.6151
R2031 B.n302 B.n301 10.6151
R2032 B.n302 B.n151 10.6151
R2033 B.n306 B.n151 10.6151
R2034 B.n307 B.n306 10.6151
R2035 B.n308 B.n307 10.6151
R2036 B.n308 B.n149 10.6151
R2037 B.n312 B.n149 10.6151
R2038 B.n313 B.n312 10.6151
R2039 B.n317 B.n313 10.6151
R2040 B.n321 B.n147 10.6151
R2041 B.n322 B.n321 10.6151
R2042 B.n323 B.n322 10.6151
R2043 B.n323 B.n145 10.6151
R2044 B.n327 B.n145 10.6151
R2045 B.n328 B.n327 10.6151
R2046 B.n329 B.n328 10.6151
R2047 B.n329 B.n143 10.6151
R2048 B.n333 B.n143 10.6151
R2049 B.n336 B.n335 10.6151
R2050 B.n336 B.n139 10.6151
R2051 B.n340 B.n139 10.6151
R2052 B.n341 B.n340 10.6151
R2053 B.n342 B.n341 10.6151
R2054 B.n342 B.n137 10.6151
R2055 B.n346 B.n137 10.6151
R2056 B.n347 B.n346 10.6151
R2057 B.n348 B.n347 10.6151
R2058 B.n348 B.n135 10.6151
R2059 B.n352 B.n135 10.6151
R2060 B.n353 B.n352 10.6151
R2061 B.n354 B.n353 10.6151
R2062 B.n354 B.n133 10.6151
R2063 B.n358 B.n133 10.6151
R2064 B.n359 B.n358 10.6151
R2065 B.n360 B.n359 10.6151
R2066 B.n360 B.n131 10.6151
R2067 B.n364 B.n131 10.6151
R2068 B.n365 B.n364 10.6151
R2069 B.n366 B.n365 10.6151
R2070 B.n366 B.n129 10.6151
R2071 B.n370 B.n129 10.6151
R2072 B.n371 B.n370 10.6151
R2073 B.n372 B.n371 10.6151
R2074 B.n372 B.n127 10.6151
R2075 B.n376 B.n127 10.6151
R2076 B.n377 B.n376 10.6151
R2077 B.n378 B.n377 10.6151
R2078 B.n378 B.n125 10.6151
R2079 B.n382 B.n125 10.6151
R2080 B.n383 B.n382 10.6151
R2081 B.n384 B.n383 10.6151
R2082 B.n384 B.n123 10.6151
R2083 B.n388 B.n123 10.6151
R2084 B.n389 B.n388 10.6151
R2085 B.n390 B.n389 10.6151
R2086 B.n390 B.n121 10.6151
R2087 B.n394 B.n121 10.6151
R2088 B.n395 B.n394 10.6151
R2089 B.n396 B.n395 10.6151
R2090 B.n396 B.n119 10.6151
R2091 B.n400 B.n119 10.6151
R2092 B.n401 B.n400 10.6151
R2093 B.n402 B.n401 10.6151
R2094 B.n402 B.n117 10.6151
R2095 B.n406 B.n117 10.6151
R2096 B.n407 B.n406 10.6151
R2097 B.n408 B.n407 10.6151
R2098 B.n408 B.n115 10.6151
R2099 B.n412 B.n115 10.6151
R2100 B.n413 B.n412 10.6151
R2101 B.n414 B.n413 10.6151
R2102 B.n414 B.n113 10.6151
R2103 B.n418 B.n113 10.6151
R2104 B.n419 B.n418 10.6151
R2105 B.n420 B.n419 10.6151
R2106 B.n420 B.n111 10.6151
R2107 B.n48 B.n44 9.36635
R2108 B.n593 B.n592 9.36635
R2109 B.n317 B.n316 9.36635
R2110 B.n335 B.n334 9.36635
R2111 B.n737 B.n0 8.11757
R2112 B.n737 B.n1 8.11757
R2113 B.n607 B.n48 1.24928
R2114 B.n594 B.n593 1.24928
R2115 B.n316 B.n147 1.24928
R2116 B.n334 B.n333 1.24928
R2117 VP.n7 VP.t6 682.245
R2118 VP.n18 VP.t0 658.399
R2119 VP.n22 VP.t5 658.399
R2120 VP.n24 VP.t9 658.399
R2121 VP.n28 VP.t3 658.399
R2122 VP.n30 VP.t7 658.399
R2123 VP.n16 VP.t4 658.399
R2124 VP.n14 VP.t2 658.399
R2125 VP.n6 VP.t1 658.399
R2126 VP.n8 VP.t8 658.399
R2127 VP.n31 VP.n30 161.3
R2128 VP.n10 VP.n9 161.3
R2129 VP.n11 VP.n6 161.3
R2130 VP.n13 VP.n12 161.3
R2131 VP.n14 VP.n5 161.3
R2132 VP.n15 VP.n4 161.3
R2133 VP.n17 VP.n16 161.3
R2134 VP.n29 VP.n0 161.3
R2135 VP.n28 VP.n27 161.3
R2136 VP.n26 VP.n1 161.3
R2137 VP.n25 VP.n24 161.3
R2138 VP.n23 VP.n2 161.3
R2139 VP.n22 VP.n21 161.3
R2140 VP.n20 VP.n3 161.3
R2141 VP.n19 VP.n18 161.3
R2142 VP.n19 VP.n17 47.5043
R2143 VP.n10 VP.n7 44.9119
R2144 VP.n18 VP.n3 35.055
R2145 VP.n30 VP.n29 35.055
R2146 VP.n16 VP.n15 35.055
R2147 VP.n23 VP.n22 27.752
R2148 VP.n28 VP.n1 27.752
R2149 VP.n14 VP.n13 27.752
R2150 VP.n9 VP.n8 27.752
R2151 VP.n24 VP.n23 20.449
R2152 VP.n24 VP.n1 20.449
R2153 VP.n13 VP.n6 20.449
R2154 VP.n9 VP.n6 20.449
R2155 VP.n8 VP.n7 17.739
R2156 VP.n22 VP.n3 13.146
R2157 VP.n29 VP.n28 13.146
R2158 VP.n15 VP.n14 13.146
R2159 VP.n11 VP.n10 0.189894
R2160 VP.n12 VP.n11 0.189894
R2161 VP.n12 VP.n5 0.189894
R2162 VP.n5 VP.n4 0.189894
R2163 VP.n17 VP.n4 0.189894
R2164 VP.n20 VP.n19 0.189894
R2165 VP.n21 VP.n20 0.189894
R2166 VP.n21 VP.n2 0.189894
R2167 VP.n25 VP.n2 0.189894
R2168 VP.n26 VP.n25 0.189894
R2169 VP.n27 VP.n26 0.189894
R2170 VP.n27 VP.n0 0.189894
R2171 VP.n31 VP.n0 0.189894
R2172 VP VP.n31 0.0516364
R2173 VDD1.n98 VDD1.n97 756.745
R2174 VDD1.n199 VDD1.n198 756.745
R2175 VDD1.n97 VDD1.n96 585
R2176 VDD1.n2 VDD1.n1 585
R2177 VDD1.n91 VDD1.n90 585
R2178 VDD1.n89 VDD1.n88 585
R2179 VDD1.n6 VDD1.n5 585
R2180 VDD1.n83 VDD1.n82 585
R2181 VDD1.n81 VDD1.n80 585
R2182 VDD1.n10 VDD1.n9 585
R2183 VDD1.n75 VDD1.n74 585
R2184 VDD1.n73 VDD1.n72 585
R2185 VDD1.n14 VDD1.n13 585
R2186 VDD1.n67 VDD1.n66 585
R2187 VDD1.n65 VDD1.n64 585
R2188 VDD1.n18 VDD1.n17 585
R2189 VDD1.n59 VDD1.n58 585
R2190 VDD1.n57 VDD1.n56 585
R2191 VDD1.n55 VDD1.n21 585
R2192 VDD1.n25 VDD1.n22 585
R2193 VDD1.n50 VDD1.n49 585
R2194 VDD1.n48 VDD1.n47 585
R2195 VDD1.n27 VDD1.n26 585
R2196 VDD1.n42 VDD1.n41 585
R2197 VDD1.n40 VDD1.n39 585
R2198 VDD1.n31 VDD1.n30 585
R2199 VDD1.n34 VDD1.n33 585
R2200 VDD1.n134 VDD1.n133 585
R2201 VDD1.n131 VDD1.n130 585
R2202 VDD1.n140 VDD1.n139 585
R2203 VDD1.n142 VDD1.n141 585
R2204 VDD1.n127 VDD1.n126 585
R2205 VDD1.n148 VDD1.n147 585
R2206 VDD1.n151 VDD1.n150 585
R2207 VDD1.n149 VDD1.n123 585
R2208 VDD1.n156 VDD1.n122 585
R2209 VDD1.n158 VDD1.n157 585
R2210 VDD1.n160 VDD1.n159 585
R2211 VDD1.n119 VDD1.n118 585
R2212 VDD1.n166 VDD1.n165 585
R2213 VDD1.n168 VDD1.n167 585
R2214 VDD1.n115 VDD1.n114 585
R2215 VDD1.n174 VDD1.n173 585
R2216 VDD1.n176 VDD1.n175 585
R2217 VDD1.n111 VDD1.n110 585
R2218 VDD1.n182 VDD1.n181 585
R2219 VDD1.n184 VDD1.n183 585
R2220 VDD1.n107 VDD1.n106 585
R2221 VDD1.n190 VDD1.n189 585
R2222 VDD1.n192 VDD1.n191 585
R2223 VDD1.n103 VDD1.n102 585
R2224 VDD1.n198 VDD1.n197 585
R2225 VDD1.t3 VDD1.n32 329.036
R2226 VDD1.t9 VDD1.n132 329.036
R2227 VDD1.n97 VDD1.n1 171.744
R2228 VDD1.n90 VDD1.n1 171.744
R2229 VDD1.n90 VDD1.n89 171.744
R2230 VDD1.n89 VDD1.n5 171.744
R2231 VDD1.n82 VDD1.n5 171.744
R2232 VDD1.n82 VDD1.n81 171.744
R2233 VDD1.n81 VDD1.n9 171.744
R2234 VDD1.n74 VDD1.n9 171.744
R2235 VDD1.n74 VDD1.n73 171.744
R2236 VDD1.n73 VDD1.n13 171.744
R2237 VDD1.n66 VDD1.n13 171.744
R2238 VDD1.n66 VDD1.n65 171.744
R2239 VDD1.n65 VDD1.n17 171.744
R2240 VDD1.n58 VDD1.n17 171.744
R2241 VDD1.n58 VDD1.n57 171.744
R2242 VDD1.n57 VDD1.n21 171.744
R2243 VDD1.n25 VDD1.n21 171.744
R2244 VDD1.n49 VDD1.n25 171.744
R2245 VDD1.n49 VDD1.n48 171.744
R2246 VDD1.n48 VDD1.n26 171.744
R2247 VDD1.n41 VDD1.n26 171.744
R2248 VDD1.n41 VDD1.n40 171.744
R2249 VDD1.n40 VDD1.n30 171.744
R2250 VDD1.n33 VDD1.n30 171.744
R2251 VDD1.n133 VDD1.n130 171.744
R2252 VDD1.n140 VDD1.n130 171.744
R2253 VDD1.n141 VDD1.n140 171.744
R2254 VDD1.n141 VDD1.n126 171.744
R2255 VDD1.n148 VDD1.n126 171.744
R2256 VDD1.n150 VDD1.n148 171.744
R2257 VDD1.n150 VDD1.n149 171.744
R2258 VDD1.n149 VDD1.n122 171.744
R2259 VDD1.n158 VDD1.n122 171.744
R2260 VDD1.n159 VDD1.n158 171.744
R2261 VDD1.n159 VDD1.n118 171.744
R2262 VDD1.n166 VDD1.n118 171.744
R2263 VDD1.n167 VDD1.n166 171.744
R2264 VDD1.n167 VDD1.n114 171.744
R2265 VDD1.n174 VDD1.n114 171.744
R2266 VDD1.n175 VDD1.n174 171.744
R2267 VDD1.n175 VDD1.n110 171.744
R2268 VDD1.n182 VDD1.n110 171.744
R2269 VDD1.n183 VDD1.n182 171.744
R2270 VDD1.n183 VDD1.n106 171.744
R2271 VDD1.n190 VDD1.n106 171.744
R2272 VDD1.n191 VDD1.n190 171.744
R2273 VDD1.n191 VDD1.n102 171.744
R2274 VDD1.n198 VDD1.n102 171.744
R2275 VDD1.n33 VDD1.t3 85.8723
R2276 VDD1.n133 VDD1.t9 85.8723
R2277 VDD1.n203 VDD1.n202 72.0652
R2278 VDD1.n100 VDD1.n99 71.4418
R2279 VDD1.n201 VDD1.n200 71.4416
R2280 VDD1.n205 VDD1.n204 71.4406
R2281 VDD1.n100 VDD1.n98 51.7087
R2282 VDD1.n201 VDD1.n199 51.7087
R2283 VDD1.n205 VDD1.n203 44.6022
R2284 VDD1.n56 VDD1.n55 13.1884
R2285 VDD1.n157 VDD1.n156 13.1884
R2286 VDD1.n59 VDD1.n20 12.8005
R2287 VDD1.n54 VDD1.n22 12.8005
R2288 VDD1.n155 VDD1.n123 12.8005
R2289 VDD1.n160 VDD1.n121 12.8005
R2290 VDD1.n96 VDD1.n0 12.0247
R2291 VDD1.n60 VDD1.n18 12.0247
R2292 VDD1.n51 VDD1.n50 12.0247
R2293 VDD1.n152 VDD1.n151 12.0247
R2294 VDD1.n161 VDD1.n119 12.0247
R2295 VDD1.n197 VDD1.n101 12.0247
R2296 VDD1.n95 VDD1.n2 11.249
R2297 VDD1.n64 VDD1.n63 11.249
R2298 VDD1.n47 VDD1.n24 11.249
R2299 VDD1.n147 VDD1.n125 11.249
R2300 VDD1.n165 VDD1.n164 11.249
R2301 VDD1.n196 VDD1.n103 11.249
R2302 VDD1.n34 VDD1.n32 10.7239
R2303 VDD1.n134 VDD1.n132 10.7239
R2304 VDD1.n92 VDD1.n91 10.4732
R2305 VDD1.n67 VDD1.n16 10.4732
R2306 VDD1.n46 VDD1.n27 10.4732
R2307 VDD1.n146 VDD1.n127 10.4732
R2308 VDD1.n168 VDD1.n117 10.4732
R2309 VDD1.n193 VDD1.n192 10.4732
R2310 VDD1.n88 VDD1.n4 9.69747
R2311 VDD1.n68 VDD1.n14 9.69747
R2312 VDD1.n43 VDD1.n42 9.69747
R2313 VDD1.n143 VDD1.n142 9.69747
R2314 VDD1.n169 VDD1.n115 9.69747
R2315 VDD1.n189 VDD1.n105 9.69747
R2316 VDD1.n94 VDD1.n0 9.45567
R2317 VDD1.n195 VDD1.n101 9.45567
R2318 VDD1.n36 VDD1.n35 9.3005
R2319 VDD1.n38 VDD1.n37 9.3005
R2320 VDD1.n29 VDD1.n28 9.3005
R2321 VDD1.n44 VDD1.n43 9.3005
R2322 VDD1.n46 VDD1.n45 9.3005
R2323 VDD1.n24 VDD1.n23 9.3005
R2324 VDD1.n52 VDD1.n51 9.3005
R2325 VDD1.n54 VDD1.n53 9.3005
R2326 VDD1.n8 VDD1.n7 9.3005
R2327 VDD1.n85 VDD1.n84 9.3005
R2328 VDD1.n87 VDD1.n86 9.3005
R2329 VDD1.n4 VDD1.n3 9.3005
R2330 VDD1.n93 VDD1.n92 9.3005
R2331 VDD1.n95 VDD1.n94 9.3005
R2332 VDD1.n79 VDD1.n78 9.3005
R2333 VDD1.n77 VDD1.n76 9.3005
R2334 VDD1.n12 VDD1.n11 9.3005
R2335 VDD1.n71 VDD1.n70 9.3005
R2336 VDD1.n69 VDD1.n68 9.3005
R2337 VDD1.n16 VDD1.n15 9.3005
R2338 VDD1.n63 VDD1.n62 9.3005
R2339 VDD1.n61 VDD1.n60 9.3005
R2340 VDD1.n20 VDD1.n19 9.3005
R2341 VDD1.n180 VDD1.n179 9.3005
R2342 VDD1.n109 VDD1.n108 9.3005
R2343 VDD1.n186 VDD1.n185 9.3005
R2344 VDD1.n188 VDD1.n187 9.3005
R2345 VDD1.n105 VDD1.n104 9.3005
R2346 VDD1.n194 VDD1.n193 9.3005
R2347 VDD1.n196 VDD1.n195 9.3005
R2348 VDD1.n113 VDD1.n112 9.3005
R2349 VDD1.n172 VDD1.n171 9.3005
R2350 VDD1.n170 VDD1.n169 9.3005
R2351 VDD1.n117 VDD1.n116 9.3005
R2352 VDD1.n164 VDD1.n163 9.3005
R2353 VDD1.n162 VDD1.n161 9.3005
R2354 VDD1.n121 VDD1.n120 9.3005
R2355 VDD1.n136 VDD1.n135 9.3005
R2356 VDD1.n138 VDD1.n137 9.3005
R2357 VDD1.n129 VDD1.n128 9.3005
R2358 VDD1.n144 VDD1.n143 9.3005
R2359 VDD1.n146 VDD1.n145 9.3005
R2360 VDD1.n125 VDD1.n124 9.3005
R2361 VDD1.n153 VDD1.n152 9.3005
R2362 VDD1.n155 VDD1.n154 9.3005
R2363 VDD1.n178 VDD1.n177 9.3005
R2364 VDD1.n87 VDD1.n6 8.92171
R2365 VDD1.n72 VDD1.n71 8.92171
R2366 VDD1.n39 VDD1.n29 8.92171
R2367 VDD1.n139 VDD1.n129 8.92171
R2368 VDD1.n173 VDD1.n172 8.92171
R2369 VDD1.n188 VDD1.n107 8.92171
R2370 VDD1.n84 VDD1.n83 8.14595
R2371 VDD1.n75 VDD1.n12 8.14595
R2372 VDD1.n38 VDD1.n31 8.14595
R2373 VDD1.n138 VDD1.n131 8.14595
R2374 VDD1.n176 VDD1.n113 8.14595
R2375 VDD1.n185 VDD1.n184 8.14595
R2376 VDD1.n80 VDD1.n8 7.3702
R2377 VDD1.n76 VDD1.n10 7.3702
R2378 VDD1.n35 VDD1.n34 7.3702
R2379 VDD1.n135 VDD1.n134 7.3702
R2380 VDD1.n177 VDD1.n111 7.3702
R2381 VDD1.n181 VDD1.n109 7.3702
R2382 VDD1.n80 VDD1.n79 6.59444
R2383 VDD1.n79 VDD1.n10 6.59444
R2384 VDD1.n180 VDD1.n111 6.59444
R2385 VDD1.n181 VDD1.n180 6.59444
R2386 VDD1.n83 VDD1.n8 5.81868
R2387 VDD1.n76 VDD1.n75 5.81868
R2388 VDD1.n35 VDD1.n31 5.81868
R2389 VDD1.n135 VDD1.n131 5.81868
R2390 VDD1.n177 VDD1.n176 5.81868
R2391 VDD1.n184 VDD1.n109 5.81868
R2392 VDD1.n84 VDD1.n6 5.04292
R2393 VDD1.n72 VDD1.n12 5.04292
R2394 VDD1.n39 VDD1.n38 5.04292
R2395 VDD1.n139 VDD1.n138 5.04292
R2396 VDD1.n173 VDD1.n113 5.04292
R2397 VDD1.n185 VDD1.n107 5.04292
R2398 VDD1.n88 VDD1.n87 4.26717
R2399 VDD1.n71 VDD1.n14 4.26717
R2400 VDD1.n42 VDD1.n29 4.26717
R2401 VDD1.n142 VDD1.n129 4.26717
R2402 VDD1.n172 VDD1.n115 4.26717
R2403 VDD1.n189 VDD1.n188 4.26717
R2404 VDD1.n91 VDD1.n4 3.49141
R2405 VDD1.n68 VDD1.n67 3.49141
R2406 VDD1.n43 VDD1.n27 3.49141
R2407 VDD1.n143 VDD1.n127 3.49141
R2408 VDD1.n169 VDD1.n168 3.49141
R2409 VDD1.n192 VDD1.n105 3.49141
R2410 VDD1.n92 VDD1.n2 2.71565
R2411 VDD1.n64 VDD1.n16 2.71565
R2412 VDD1.n47 VDD1.n46 2.71565
R2413 VDD1.n147 VDD1.n146 2.71565
R2414 VDD1.n165 VDD1.n117 2.71565
R2415 VDD1.n193 VDD1.n103 2.71565
R2416 VDD1.n36 VDD1.n32 2.41282
R2417 VDD1.n136 VDD1.n132 2.41282
R2418 VDD1.n96 VDD1.n95 1.93989
R2419 VDD1.n63 VDD1.n18 1.93989
R2420 VDD1.n50 VDD1.n24 1.93989
R2421 VDD1.n151 VDD1.n125 1.93989
R2422 VDD1.n164 VDD1.n119 1.93989
R2423 VDD1.n197 VDD1.n196 1.93989
R2424 VDD1.n204 VDD1.t7 1.80233
R2425 VDD1.n204 VDD1.t5 1.80233
R2426 VDD1.n99 VDD1.t1 1.80233
R2427 VDD1.n99 VDD1.t8 1.80233
R2428 VDD1.n202 VDD1.t6 1.80233
R2429 VDD1.n202 VDD1.t2 1.80233
R2430 VDD1.n200 VDD1.t4 1.80233
R2431 VDD1.n200 VDD1.t0 1.80233
R2432 VDD1.n98 VDD1.n0 1.16414
R2433 VDD1.n60 VDD1.n59 1.16414
R2434 VDD1.n51 VDD1.n22 1.16414
R2435 VDD1.n152 VDD1.n123 1.16414
R2436 VDD1.n161 VDD1.n160 1.16414
R2437 VDD1.n199 VDD1.n101 1.16414
R2438 VDD1 VDD1.n205 0.62119
R2439 VDD1.n56 VDD1.n20 0.388379
R2440 VDD1.n55 VDD1.n54 0.388379
R2441 VDD1.n156 VDD1.n155 0.388379
R2442 VDD1.n157 VDD1.n121 0.388379
R2443 VDD1 VDD1.n100 0.284983
R2444 VDD1.n203 VDD1.n201 0.171447
R2445 VDD1.n94 VDD1.n93 0.155672
R2446 VDD1.n93 VDD1.n3 0.155672
R2447 VDD1.n86 VDD1.n3 0.155672
R2448 VDD1.n86 VDD1.n85 0.155672
R2449 VDD1.n85 VDD1.n7 0.155672
R2450 VDD1.n78 VDD1.n7 0.155672
R2451 VDD1.n78 VDD1.n77 0.155672
R2452 VDD1.n77 VDD1.n11 0.155672
R2453 VDD1.n70 VDD1.n11 0.155672
R2454 VDD1.n70 VDD1.n69 0.155672
R2455 VDD1.n69 VDD1.n15 0.155672
R2456 VDD1.n62 VDD1.n15 0.155672
R2457 VDD1.n62 VDD1.n61 0.155672
R2458 VDD1.n61 VDD1.n19 0.155672
R2459 VDD1.n53 VDD1.n19 0.155672
R2460 VDD1.n53 VDD1.n52 0.155672
R2461 VDD1.n52 VDD1.n23 0.155672
R2462 VDD1.n45 VDD1.n23 0.155672
R2463 VDD1.n45 VDD1.n44 0.155672
R2464 VDD1.n44 VDD1.n28 0.155672
R2465 VDD1.n37 VDD1.n28 0.155672
R2466 VDD1.n37 VDD1.n36 0.155672
R2467 VDD1.n137 VDD1.n136 0.155672
R2468 VDD1.n137 VDD1.n128 0.155672
R2469 VDD1.n144 VDD1.n128 0.155672
R2470 VDD1.n145 VDD1.n144 0.155672
R2471 VDD1.n145 VDD1.n124 0.155672
R2472 VDD1.n153 VDD1.n124 0.155672
R2473 VDD1.n154 VDD1.n153 0.155672
R2474 VDD1.n154 VDD1.n120 0.155672
R2475 VDD1.n162 VDD1.n120 0.155672
R2476 VDD1.n163 VDD1.n162 0.155672
R2477 VDD1.n163 VDD1.n116 0.155672
R2478 VDD1.n170 VDD1.n116 0.155672
R2479 VDD1.n171 VDD1.n170 0.155672
R2480 VDD1.n171 VDD1.n112 0.155672
R2481 VDD1.n178 VDD1.n112 0.155672
R2482 VDD1.n179 VDD1.n178 0.155672
R2483 VDD1.n179 VDD1.n108 0.155672
R2484 VDD1.n186 VDD1.n108 0.155672
R2485 VDD1.n187 VDD1.n186 0.155672
R2486 VDD1.n187 VDD1.n104 0.155672
R2487 VDD1.n194 VDD1.n104 0.155672
R2488 VDD1.n195 VDD1.n194 0.155672
C0 B VP 1.34482f
C1 VDD2 B 2.19734f
C2 VP VDD1 10.1839f
C3 B VTAIL 3.8262f
C4 VDD2 VDD1 0.984587f
C5 VTAIL VDD1 19.827f
C6 w_n2230_n4576# VN 4.30872f
C7 B VDD1 2.1523f
C8 w_n2230_n4576# VP 4.59325f
C9 VDD2 w_n2230_n4576# 2.53582f
C10 w_n2230_n4576# VTAIL 3.93475f
C11 VP VN 6.74094f
C12 VDD2 VN 9.99471f
C13 VN VTAIL 9.61297f
C14 w_n2230_n4576# B 9.081111f
C15 w_n2230_n4576# VDD1 2.49019f
C16 B VN 0.876729f
C17 VDD2 VP 0.345068f
C18 VN VDD1 0.1491f
C19 VP VTAIL 9.62781f
C20 VDD2 VTAIL 19.858099f
C21 VDD2 VSUBS 1.696726f
C22 VDD1 VSUBS 1.364362f
C23 VTAIL VSUBS 0.953737f
C24 VN VSUBS 5.40922f
C25 VP VSUBS 2.070095f
C26 B VSUBS 3.548458f
C27 w_n2230_n4576# VSUBS 0.124782p
C28 VDD1.n0 VSUBS 0.015872f
C29 VDD1.n1 VSUBS 0.035814f
C30 VDD1.n2 VSUBS 0.016043f
C31 VDD1.n3 VSUBS 0.028197f
C32 VDD1.n4 VSUBS 0.015152f
C33 VDD1.n5 VSUBS 0.035814f
C34 VDD1.n6 VSUBS 0.016043f
C35 VDD1.n7 VSUBS 0.028197f
C36 VDD1.n8 VSUBS 0.015152f
C37 VDD1.n9 VSUBS 0.035814f
C38 VDD1.n10 VSUBS 0.016043f
C39 VDD1.n11 VSUBS 0.028197f
C40 VDD1.n12 VSUBS 0.015152f
C41 VDD1.n13 VSUBS 0.035814f
C42 VDD1.n14 VSUBS 0.016043f
C43 VDD1.n15 VSUBS 0.028197f
C44 VDD1.n16 VSUBS 0.015152f
C45 VDD1.n17 VSUBS 0.035814f
C46 VDD1.n18 VSUBS 0.016043f
C47 VDD1.n19 VSUBS 0.028197f
C48 VDD1.n20 VSUBS 0.015152f
C49 VDD1.n21 VSUBS 0.035814f
C50 VDD1.n22 VSUBS 0.016043f
C51 VDD1.n23 VSUBS 0.028197f
C52 VDD1.n24 VSUBS 0.015152f
C53 VDD1.n25 VSUBS 0.035814f
C54 VDD1.n26 VSUBS 0.035814f
C55 VDD1.n27 VSUBS 0.016043f
C56 VDD1.n28 VSUBS 0.028197f
C57 VDD1.n29 VSUBS 0.015152f
C58 VDD1.n30 VSUBS 0.035814f
C59 VDD1.n31 VSUBS 0.016043f
C60 VDD1.n32 VSUBS 0.299076f
C61 VDD1.t3 VSUBS 0.077749f
C62 VDD1.n33 VSUBS 0.02686f
C63 VDD1.n34 VSUBS 0.026941f
C64 VDD1.n35 VSUBS 0.015152f
C65 VDD1.n36 VSUBS 2.13167f
C66 VDD1.n37 VSUBS 0.028197f
C67 VDD1.n38 VSUBS 0.015152f
C68 VDD1.n39 VSUBS 0.016043f
C69 VDD1.n40 VSUBS 0.035814f
C70 VDD1.n41 VSUBS 0.035814f
C71 VDD1.n42 VSUBS 0.016043f
C72 VDD1.n43 VSUBS 0.015152f
C73 VDD1.n44 VSUBS 0.028197f
C74 VDD1.n45 VSUBS 0.028197f
C75 VDD1.n46 VSUBS 0.015152f
C76 VDD1.n47 VSUBS 0.016043f
C77 VDD1.n48 VSUBS 0.035814f
C78 VDD1.n49 VSUBS 0.035814f
C79 VDD1.n50 VSUBS 0.016043f
C80 VDD1.n51 VSUBS 0.015152f
C81 VDD1.n52 VSUBS 0.028197f
C82 VDD1.n53 VSUBS 0.028197f
C83 VDD1.n54 VSUBS 0.015152f
C84 VDD1.n55 VSUBS 0.015598f
C85 VDD1.n56 VSUBS 0.015598f
C86 VDD1.n57 VSUBS 0.035814f
C87 VDD1.n58 VSUBS 0.035814f
C88 VDD1.n59 VSUBS 0.016043f
C89 VDD1.n60 VSUBS 0.015152f
C90 VDD1.n61 VSUBS 0.028197f
C91 VDD1.n62 VSUBS 0.028197f
C92 VDD1.n63 VSUBS 0.015152f
C93 VDD1.n64 VSUBS 0.016043f
C94 VDD1.n65 VSUBS 0.035814f
C95 VDD1.n66 VSUBS 0.035814f
C96 VDD1.n67 VSUBS 0.016043f
C97 VDD1.n68 VSUBS 0.015152f
C98 VDD1.n69 VSUBS 0.028197f
C99 VDD1.n70 VSUBS 0.028197f
C100 VDD1.n71 VSUBS 0.015152f
C101 VDD1.n72 VSUBS 0.016043f
C102 VDD1.n73 VSUBS 0.035814f
C103 VDD1.n74 VSUBS 0.035814f
C104 VDD1.n75 VSUBS 0.016043f
C105 VDD1.n76 VSUBS 0.015152f
C106 VDD1.n77 VSUBS 0.028197f
C107 VDD1.n78 VSUBS 0.028197f
C108 VDD1.n79 VSUBS 0.015152f
C109 VDD1.n80 VSUBS 0.016043f
C110 VDD1.n81 VSUBS 0.035814f
C111 VDD1.n82 VSUBS 0.035814f
C112 VDD1.n83 VSUBS 0.016043f
C113 VDD1.n84 VSUBS 0.015152f
C114 VDD1.n85 VSUBS 0.028197f
C115 VDD1.n86 VSUBS 0.028197f
C116 VDD1.n87 VSUBS 0.015152f
C117 VDD1.n88 VSUBS 0.016043f
C118 VDD1.n89 VSUBS 0.035814f
C119 VDD1.n90 VSUBS 0.035814f
C120 VDD1.n91 VSUBS 0.016043f
C121 VDD1.n92 VSUBS 0.015152f
C122 VDD1.n93 VSUBS 0.028197f
C123 VDD1.n94 VSUBS 0.07134f
C124 VDD1.n95 VSUBS 0.015152f
C125 VDD1.n96 VSUBS 0.016043f
C126 VDD1.n97 VSUBS 0.078157f
C127 VDD1.n98 VSUBS 0.073997f
C128 VDD1.t1 VSUBS 0.401973f
C129 VDD1.t8 VSUBS 0.401973f
C130 VDD1.n99 VSUBS 3.3646f
C131 VDD1.n100 VSUBS 0.776386f
C132 VDD1.n101 VSUBS 0.015872f
C133 VDD1.n102 VSUBS 0.035814f
C134 VDD1.n103 VSUBS 0.016043f
C135 VDD1.n104 VSUBS 0.028197f
C136 VDD1.n105 VSUBS 0.015152f
C137 VDD1.n106 VSUBS 0.035814f
C138 VDD1.n107 VSUBS 0.016043f
C139 VDD1.n108 VSUBS 0.028197f
C140 VDD1.n109 VSUBS 0.015152f
C141 VDD1.n110 VSUBS 0.035814f
C142 VDD1.n111 VSUBS 0.016043f
C143 VDD1.n112 VSUBS 0.028197f
C144 VDD1.n113 VSUBS 0.015152f
C145 VDD1.n114 VSUBS 0.035814f
C146 VDD1.n115 VSUBS 0.016043f
C147 VDD1.n116 VSUBS 0.028197f
C148 VDD1.n117 VSUBS 0.015152f
C149 VDD1.n118 VSUBS 0.035814f
C150 VDD1.n119 VSUBS 0.016043f
C151 VDD1.n120 VSUBS 0.028197f
C152 VDD1.n121 VSUBS 0.015152f
C153 VDD1.n122 VSUBS 0.035814f
C154 VDD1.n123 VSUBS 0.016043f
C155 VDD1.n124 VSUBS 0.028197f
C156 VDD1.n125 VSUBS 0.015152f
C157 VDD1.n126 VSUBS 0.035814f
C158 VDD1.n127 VSUBS 0.016043f
C159 VDD1.n128 VSUBS 0.028197f
C160 VDD1.n129 VSUBS 0.015152f
C161 VDD1.n130 VSUBS 0.035814f
C162 VDD1.n131 VSUBS 0.016043f
C163 VDD1.n132 VSUBS 0.299076f
C164 VDD1.t9 VSUBS 0.077749f
C165 VDD1.n133 VSUBS 0.02686f
C166 VDD1.n134 VSUBS 0.026941f
C167 VDD1.n135 VSUBS 0.015152f
C168 VDD1.n136 VSUBS 2.13167f
C169 VDD1.n137 VSUBS 0.028197f
C170 VDD1.n138 VSUBS 0.015152f
C171 VDD1.n139 VSUBS 0.016043f
C172 VDD1.n140 VSUBS 0.035814f
C173 VDD1.n141 VSUBS 0.035814f
C174 VDD1.n142 VSUBS 0.016043f
C175 VDD1.n143 VSUBS 0.015152f
C176 VDD1.n144 VSUBS 0.028197f
C177 VDD1.n145 VSUBS 0.028197f
C178 VDD1.n146 VSUBS 0.015152f
C179 VDD1.n147 VSUBS 0.016043f
C180 VDD1.n148 VSUBS 0.035814f
C181 VDD1.n149 VSUBS 0.035814f
C182 VDD1.n150 VSUBS 0.035814f
C183 VDD1.n151 VSUBS 0.016043f
C184 VDD1.n152 VSUBS 0.015152f
C185 VDD1.n153 VSUBS 0.028197f
C186 VDD1.n154 VSUBS 0.028197f
C187 VDD1.n155 VSUBS 0.015152f
C188 VDD1.n156 VSUBS 0.015598f
C189 VDD1.n157 VSUBS 0.015598f
C190 VDD1.n158 VSUBS 0.035814f
C191 VDD1.n159 VSUBS 0.035814f
C192 VDD1.n160 VSUBS 0.016043f
C193 VDD1.n161 VSUBS 0.015152f
C194 VDD1.n162 VSUBS 0.028197f
C195 VDD1.n163 VSUBS 0.028197f
C196 VDD1.n164 VSUBS 0.015152f
C197 VDD1.n165 VSUBS 0.016043f
C198 VDD1.n166 VSUBS 0.035814f
C199 VDD1.n167 VSUBS 0.035814f
C200 VDD1.n168 VSUBS 0.016043f
C201 VDD1.n169 VSUBS 0.015152f
C202 VDD1.n170 VSUBS 0.028197f
C203 VDD1.n171 VSUBS 0.028197f
C204 VDD1.n172 VSUBS 0.015152f
C205 VDD1.n173 VSUBS 0.016043f
C206 VDD1.n174 VSUBS 0.035814f
C207 VDD1.n175 VSUBS 0.035814f
C208 VDD1.n176 VSUBS 0.016043f
C209 VDD1.n177 VSUBS 0.015152f
C210 VDD1.n178 VSUBS 0.028197f
C211 VDD1.n179 VSUBS 0.028197f
C212 VDD1.n180 VSUBS 0.015152f
C213 VDD1.n181 VSUBS 0.016043f
C214 VDD1.n182 VSUBS 0.035814f
C215 VDD1.n183 VSUBS 0.035814f
C216 VDD1.n184 VSUBS 0.016043f
C217 VDD1.n185 VSUBS 0.015152f
C218 VDD1.n186 VSUBS 0.028197f
C219 VDD1.n187 VSUBS 0.028197f
C220 VDD1.n188 VSUBS 0.015152f
C221 VDD1.n189 VSUBS 0.016043f
C222 VDD1.n190 VSUBS 0.035814f
C223 VDD1.n191 VSUBS 0.035814f
C224 VDD1.n192 VSUBS 0.016043f
C225 VDD1.n193 VSUBS 0.015152f
C226 VDD1.n194 VSUBS 0.028197f
C227 VDD1.n195 VSUBS 0.07134f
C228 VDD1.n196 VSUBS 0.015152f
C229 VDD1.n197 VSUBS 0.016043f
C230 VDD1.n198 VSUBS 0.078157f
C231 VDD1.n199 VSUBS 0.073997f
C232 VDD1.t4 VSUBS 0.401973f
C233 VDD1.t0 VSUBS 0.401973f
C234 VDD1.n200 VSUBS 3.36459f
C235 VDD1.n201 VSUBS 0.769904f
C236 VDD1.t6 VSUBS 0.401973f
C237 VDD1.t2 VSUBS 0.401973f
C238 VDD1.n202 VSUBS 3.3705f
C239 VDD1.n203 VSUBS 2.96718f
C240 VDD1.t7 VSUBS 0.401973f
C241 VDD1.t5 VSUBS 0.401973f
C242 VDD1.n204 VSUBS 3.36459f
C243 VDD1.n205 VSUBS 3.52389f
C244 VP.n0 VSUBS 0.04964f
C245 VP.n1 VSUBS 0.011264f
C246 VP.n2 VSUBS 0.04964f
C247 VP.n3 VSUBS 0.011264f
C248 VP.n4 VSUBS 0.04964f
C249 VP.t4 VSUBS 1.82798f
C250 VP.t2 VSUBS 1.82798f
C251 VP.n5 VSUBS 0.04964f
C252 VP.t1 VSUBS 1.82798f
C253 VP.n6 VSUBS 0.688507f
C254 VP.t6 VSUBS 1.85207f
C255 VP.n7 VSUBS 0.669354f
C256 VP.t8 VSUBS 1.82798f
C257 VP.n8 VSUBS 0.694656f
C258 VP.n9 VSUBS 0.011264f
C259 VP.n10 VSUBS 0.210371f
C260 VP.n11 VSUBS 0.04964f
C261 VP.n12 VSUBS 0.04964f
C262 VP.n13 VSUBS 0.011264f
C263 VP.n14 VSUBS 0.688507f
C264 VP.n15 VSUBS 0.011264f
C265 VP.n16 VSUBS 0.687283f
C266 VP.n17 VSUBS 2.49615f
C267 VP.t0 VSUBS 1.82798f
C268 VP.n18 VSUBS 0.687283f
C269 VP.n19 VSUBS 2.53382f
C270 VP.n20 VSUBS 0.04964f
C271 VP.n21 VSUBS 0.04964f
C272 VP.t5 VSUBS 1.82798f
C273 VP.n22 VSUBS 0.688507f
C274 VP.n23 VSUBS 0.011264f
C275 VP.t9 VSUBS 1.82798f
C276 VP.n24 VSUBS 0.688507f
C277 VP.n25 VSUBS 0.04964f
C278 VP.n26 VSUBS 0.04964f
C279 VP.n27 VSUBS 0.04964f
C280 VP.t3 VSUBS 1.82798f
C281 VP.n28 VSUBS 0.688507f
C282 VP.n29 VSUBS 0.011264f
C283 VP.t7 VSUBS 1.82798f
C284 VP.n30 VSUBS 0.687283f
C285 VP.n31 VSUBS 0.038469f
C286 B.n0 VSUBS 0.008011f
C287 B.n1 VSUBS 0.008011f
C288 B.n2 VSUBS 0.011847f
C289 B.n3 VSUBS 0.009079f
C290 B.n4 VSUBS 0.009079f
C291 B.n5 VSUBS 0.009079f
C292 B.n6 VSUBS 0.009079f
C293 B.n7 VSUBS 0.009079f
C294 B.n8 VSUBS 0.009079f
C295 B.n9 VSUBS 0.009079f
C296 B.n10 VSUBS 0.009079f
C297 B.n11 VSUBS 0.009079f
C298 B.n12 VSUBS 0.009079f
C299 B.n13 VSUBS 0.009079f
C300 B.n14 VSUBS 0.009079f
C301 B.n15 VSUBS 0.023005f
C302 B.n16 VSUBS 0.009079f
C303 B.n17 VSUBS 0.009079f
C304 B.n18 VSUBS 0.009079f
C305 B.n19 VSUBS 0.009079f
C306 B.n20 VSUBS 0.009079f
C307 B.n21 VSUBS 0.009079f
C308 B.n22 VSUBS 0.009079f
C309 B.n23 VSUBS 0.009079f
C310 B.n24 VSUBS 0.009079f
C311 B.n25 VSUBS 0.009079f
C312 B.n26 VSUBS 0.009079f
C313 B.n27 VSUBS 0.009079f
C314 B.n28 VSUBS 0.009079f
C315 B.n29 VSUBS 0.009079f
C316 B.n30 VSUBS 0.009079f
C317 B.n31 VSUBS 0.009079f
C318 B.n32 VSUBS 0.009079f
C319 B.n33 VSUBS 0.009079f
C320 B.n34 VSUBS 0.009079f
C321 B.n35 VSUBS 0.009079f
C322 B.n36 VSUBS 0.009079f
C323 B.n37 VSUBS 0.009079f
C324 B.n38 VSUBS 0.009079f
C325 B.n39 VSUBS 0.009079f
C326 B.n40 VSUBS 0.009079f
C327 B.n41 VSUBS 0.009079f
C328 B.n42 VSUBS 0.009079f
C329 B.n43 VSUBS 0.009079f
C330 B.n44 VSUBS 0.008545f
C331 B.n45 VSUBS 0.009079f
C332 B.t10 VSUBS 0.456295f
C333 B.t11 VSUBS 0.472607f
C334 B.t9 VSUBS 0.680081f
C335 B.n46 VSUBS 0.572074f
C336 B.n47 VSUBS 0.417129f
C337 B.n48 VSUBS 0.021034f
C338 B.n49 VSUBS 0.009079f
C339 B.n50 VSUBS 0.009079f
C340 B.n51 VSUBS 0.009079f
C341 B.n52 VSUBS 0.009079f
C342 B.t4 VSUBS 0.4563f
C343 B.t5 VSUBS 0.472612f
C344 B.t3 VSUBS 0.680081f
C345 B.n53 VSUBS 0.57207f
C346 B.n54 VSUBS 0.417124f
C347 B.n55 VSUBS 0.009079f
C348 B.n56 VSUBS 0.009079f
C349 B.n57 VSUBS 0.009079f
C350 B.n58 VSUBS 0.009079f
C351 B.n59 VSUBS 0.009079f
C352 B.n60 VSUBS 0.009079f
C353 B.n61 VSUBS 0.009079f
C354 B.n62 VSUBS 0.009079f
C355 B.n63 VSUBS 0.009079f
C356 B.n64 VSUBS 0.009079f
C357 B.n65 VSUBS 0.009079f
C358 B.n66 VSUBS 0.009079f
C359 B.n67 VSUBS 0.009079f
C360 B.n68 VSUBS 0.009079f
C361 B.n69 VSUBS 0.009079f
C362 B.n70 VSUBS 0.009079f
C363 B.n71 VSUBS 0.009079f
C364 B.n72 VSUBS 0.009079f
C365 B.n73 VSUBS 0.009079f
C366 B.n74 VSUBS 0.009079f
C367 B.n75 VSUBS 0.009079f
C368 B.n76 VSUBS 0.009079f
C369 B.n77 VSUBS 0.009079f
C370 B.n78 VSUBS 0.009079f
C371 B.n79 VSUBS 0.009079f
C372 B.n80 VSUBS 0.009079f
C373 B.n81 VSUBS 0.009079f
C374 B.n82 VSUBS 0.009079f
C375 B.n83 VSUBS 0.009079f
C376 B.n84 VSUBS 0.022121f
C377 B.n85 VSUBS 0.009079f
C378 B.n86 VSUBS 0.009079f
C379 B.n87 VSUBS 0.009079f
C380 B.n88 VSUBS 0.009079f
C381 B.n89 VSUBS 0.009079f
C382 B.n90 VSUBS 0.009079f
C383 B.n91 VSUBS 0.009079f
C384 B.n92 VSUBS 0.009079f
C385 B.n93 VSUBS 0.009079f
C386 B.n94 VSUBS 0.009079f
C387 B.n95 VSUBS 0.009079f
C388 B.n96 VSUBS 0.009079f
C389 B.n97 VSUBS 0.009079f
C390 B.n98 VSUBS 0.009079f
C391 B.n99 VSUBS 0.009079f
C392 B.n100 VSUBS 0.009079f
C393 B.n101 VSUBS 0.009079f
C394 B.n102 VSUBS 0.009079f
C395 B.n103 VSUBS 0.009079f
C396 B.n104 VSUBS 0.009079f
C397 B.n105 VSUBS 0.009079f
C398 B.n106 VSUBS 0.009079f
C399 B.n107 VSUBS 0.009079f
C400 B.n108 VSUBS 0.009079f
C401 B.n109 VSUBS 0.009079f
C402 B.n110 VSUBS 0.009079f
C403 B.n111 VSUBS 0.022025f
C404 B.n112 VSUBS 0.009079f
C405 B.n113 VSUBS 0.009079f
C406 B.n114 VSUBS 0.009079f
C407 B.n115 VSUBS 0.009079f
C408 B.n116 VSUBS 0.009079f
C409 B.n117 VSUBS 0.009079f
C410 B.n118 VSUBS 0.009079f
C411 B.n119 VSUBS 0.009079f
C412 B.n120 VSUBS 0.009079f
C413 B.n121 VSUBS 0.009079f
C414 B.n122 VSUBS 0.009079f
C415 B.n123 VSUBS 0.009079f
C416 B.n124 VSUBS 0.009079f
C417 B.n125 VSUBS 0.009079f
C418 B.n126 VSUBS 0.009079f
C419 B.n127 VSUBS 0.009079f
C420 B.n128 VSUBS 0.009079f
C421 B.n129 VSUBS 0.009079f
C422 B.n130 VSUBS 0.009079f
C423 B.n131 VSUBS 0.009079f
C424 B.n132 VSUBS 0.009079f
C425 B.n133 VSUBS 0.009079f
C426 B.n134 VSUBS 0.009079f
C427 B.n135 VSUBS 0.009079f
C428 B.n136 VSUBS 0.009079f
C429 B.n137 VSUBS 0.009079f
C430 B.n138 VSUBS 0.009079f
C431 B.n139 VSUBS 0.009079f
C432 B.n140 VSUBS 0.009079f
C433 B.t2 VSUBS 0.4563f
C434 B.t1 VSUBS 0.472612f
C435 B.t0 VSUBS 0.680081f
C436 B.n141 VSUBS 0.57207f
C437 B.n142 VSUBS 0.417124f
C438 B.n143 VSUBS 0.009079f
C439 B.n144 VSUBS 0.009079f
C440 B.n145 VSUBS 0.009079f
C441 B.n146 VSUBS 0.009079f
C442 B.n147 VSUBS 0.005073f
C443 B.n148 VSUBS 0.009079f
C444 B.n149 VSUBS 0.009079f
C445 B.n150 VSUBS 0.009079f
C446 B.n151 VSUBS 0.009079f
C447 B.n152 VSUBS 0.009079f
C448 B.n153 VSUBS 0.009079f
C449 B.n154 VSUBS 0.009079f
C450 B.n155 VSUBS 0.009079f
C451 B.n156 VSUBS 0.009079f
C452 B.n157 VSUBS 0.009079f
C453 B.n158 VSUBS 0.009079f
C454 B.n159 VSUBS 0.009079f
C455 B.n160 VSUBS 0.009079f
C456 B.n161 VSUBS 0.009079f
C457 B.n162 VSUBS 0.009079f
C458 B.n163 VSUBS 0.009079f
C459 B.n164 VSUBS 0.009079f
C460 B.n165 VSUBS 0.009079f
C461 B.n166 VSUBS 0.009079f
C462 B.n167 VSUBS 0.009079f
C463 B.n168 VSUBS 0.009079f
C464 B.n169 VSUBS 0.009079f
C465 B.n170 VSUBS 0.009079f
C466 B.n171 VSUBS 0.009079f
C467 B.n172 VSUBS 0.009079f
C468 B.n173 VSUBS 0.009079f
C469 B.n174 VSUBS 0.009079f
C470 B.n175 VSUBS 0.009079f
C471 B.n176 VSUBS 0.009079f
C472 B.n177 VSUBS 0.022121f
C473 B.n178 VSUBS 0.009079f
C474 B.n179 VSUBS 0.009079f
C475 B.n180 VSUBS 0.009079f
C476 B.n181 VSUBS 0.009079f
C477 B.n182 VSUBS 0.009079f
C478 B.n183 VSUBS 0.009079f
C479 B.n184 VSUBS 0.009079f
C480 B.n185 VSUBS 0.009079f
C481 B.n186 VSUBS 0.009079f
C482 B.n187 VSUBS 0.009079f
C483 B.n188 VSUBS 0.009079f
C484 B.n189 VSUBS 0.009079f
C485 B.n190 VSUBS 0.009079f
C486 B.n191 VSUBS 0.009079f
C487 B.n192 VSUBS 0.009079f
C488 B.n193 VSUBS 0.009079f
C489 B.n194 VSUBS 0.009079f
C490 B.n195 VSUBS 0.009079f
C491 B.n196 VSUBS 0.009079f
C492 B.n197 VSUBS 0.009079f
C493 B.n198 VSUBS 0.009079f
C494 B.n199 VSUBS 0.009079f
C495 B.n200 VSUBS 0.009079f
C496 B.n201 VSUBS 0.009079f
C497 B.n202 VSUBS 0.009079f
C498 B.n203 VSUBS 0.009079f
C499 B.n204 VSUBS 0.009079f
C500 B.n205 VSUBS 0.009079f
C501 B.n206 VSUBS 0.009079f
C502 B.n207 VSUBS 0.009079f
C503 B.n208 VSUBS 0.009079f
C504 B.n209 VSUBS 0.009079f
C505 B.n210 VSUBS 0.009079f
C506 B.n211 VSUBS 0.009079f
C507 B.n212 VSUBS 0.009079f
C508 B.n213 VSUBS 0.009079f
C509 B.n214 VSUBS 0.009079f
C510 B.n215 VSUBS 0.009079f
C511 B.n216 VSUBS 0.009079f
C512 B.n217 VSUBS 0.009079f
C513 B.n218 VSUBS 0.009079f
C514 B.n219 VSUBS 0.009079f
C515 B.n220 VSUBS 0.009079f
C516 B.n221 VSUBS 0.009079f
C517 B.n222 VSUBS 0.009079f
C518 B.n223 VSUBS 0.009079f
C519 B.n224 VSUBS 0.009079f
C520 B.n225 VSUBS 0.009079f
C521 B.n226 VSUBS 0.022121f
C522 B.n227 VSUBS 0.023005f
C523 B.n228 VSUBS 0.023005f
C524 B.n229 VSUBS 0.009079f
C525 B.n230 VSUBS 0.009079f
C526 B.n231 VSUBS 0.009079f
C527 B.n232 VSUBS 0.009079f
C528 B.n233 VSUBS 0.009079f
C529 B.n234 VSUBS 0.009079f
C530 B.n235 VSUBS 0.009079f
C531 B.n236 VSUBS 0.009079f
C532 B.n237 VSUBS 0.009079f
C533 B.n238 VSUBS 0.009079f
C534 B.n239 VSUBS 0.009079f
C535 B.n240 VSUBS 0.009079f
C536 B.n241 VSUBS 0.009079f
C537 B.n242 VSUBS 0.009079f
C538 B.n243 VSUBS 0.009079f
C539 B.n244 VSUBS 0.009079f
C540 B.n245 VSUBS 0.009079f
C541 B.n246 VSUBS 0.009079f
C542 B.n247 VSUBS 0.009079f
C543 B.n248 VSUBS 0.009079f
C544 B.n249 VSUBS 0.009079f
C545 B.n250 VSUBS 0.009079f
C546 B.n251 VSUBS 0.009079f
C547 B.n252 VSUBS 0.009079f
C548 B.n253 VSUBS 0.009079f
C549 B.n254 VSUBS 0.009079f
C550 B.n255 VSUBS 0.009079f
C551 B.n256 VSUBS 0.009079f
C552 B.n257 VSUBS 0.009079f
C553 B.n258 VSUBS 0.009079f
C554 B.n259 VSUBS 0.009079f
C555 B.n260 VSUBS 0.009079f
C556 B.n261 VSUBS 0.009079f
C557 B.n262 VSUBS 0.009079f
C558 B.n263 VSUBS 0.009079f
C559 B.n264 VSUBS 0.009079f
C560 B.n265 VSUBS 0.009079f
C561 B.n266 VSUBS 0.009079f
C562 B.n267 VSUBS 0.009079f
C563 B.n268 VSUBS 0.009079f
C564 B.n269 VSUBS 0.009079f
C565 B.n270 VSUBS 0.009079f
C566 B.n271 VSUBS 0.009079f
C567 B.n272 VSUBS 0.009079f
C568 B.n273 VSUBS 0.009079f
C569 B.n274 VSUBS 0.009079f
C570 B.n275 VSUBS 0.009079f
C571 B.n276 VSUBS 0.009079f
C572 B.n277 VSUBS 0.009079f
C573 B.n278 VSUBS 0.009079f
C574 B.n279 VSUBS 0.009079f
C575 B.n280 VSUBS 0.009079f
C576 B.n281 VSUBS 0.009079f
C577 B.n282 VSUBS 0.009079f
C578 B.n283 VSUBS 0.009079f
C579 B.n284 VSUBS 0.009079f
C580 B.n285 VSUBS 0.009079f
C581 B.n286 VSUBS 0.009079f
C582 B.n287 VSUBS 0.009079f
C583 B.n288 VSUBS 0.009079f
C584 B.n289 VSUBS 0.009079f
C585 B.n290 VSUBS 0.009079f
C586 B.n291 VSUBS 0.009079f
C587 B.n292 VSUBS 0.009079f
C588 B.n293 VSUBS 0.009079f
C589 B.n294 VSUBS 0.009079f
C590 B.n295 VSUBS 0.009079f
C591 B.n296 VSUBS 0.009079f
C592 B.n297 VSUBS 0.009079f
C593 B.n298 VSUBS 0.009079f
C594 B.n299 VSUBS 0.009079f
C595 B.n300 VSUBS 0.009079f
C596 B.n301 VSUBS 0.009079f
C597 B.n302 VSUBS 0.009079f
C598 B.n303 VSUBS 0.009079f
C599 B.n304 VSUBS 0.009079f
C600 B.n305 VSUBS 0.009079f
C601 B.n306 VSUBS 0.009079f
C602 B.n307 VSUBS 0.009079f
C603 B.n308 VSUBS 0.009079f
C604 B.n309 VSUBS 0.009079f
C605 B.n310 VSUBS 0.009079f
C606 B.n311 VSUBS 0.009079f
C607 B.n312 VSUBS 0.009079f
C608 B.n313 VSUBS 0.009079f
C609 B.t8 VSUBS 0.456295f
C610 B.t7 VSUBS 0.472607f
C611 B.t6 VSUBS 0.680081f
C612 B.n314 VSUBS 0.572074f
C613 B.n315 VSUBS 0.417129f
C614 B.n316 VSUBS 0.021034f
C615 B.n317 VSUBS 0.008545f
C616 B.n318 VSUBS 0.009079f
C617 B.n319 VSUBS 0.009079f
C618 B.n320 VSUBS 0.009079f
C619 B.n321 VSUBS 0.009079f
C620 B.n322 VSUBS 0.009079f
C621 B.n323 VSUBS 0.009079f
C622 B.n324 VSUBS 0.009079f
C623 B.n325 VSUBS 0.009079f
C624 B.n326 VSUBS 0.009079f
C625 B.n327 VSUBS 0.009079f
C626 B.n328 VSUBS 0.009079f
C627 B.n329 VSUBS 0.009079f
C628 B.n330 VSUBS 0.009079f
C629 B.n331 VSUBS 0.009079f
C630 B.n332 VSUBS 0.009079f
C631 B.n333 VSUBS 0.005073f
C632 B.n334 VSUBS 0.021034f
C633 B.n335 VSUBS 0.008545f
C634 B.n336 VSUBS 0.009079f
C635 B.n337 VSUBS 0.009079f
C636 B.n338 VSUBS 0.009079f
C637 B.n339 VSUBS 0.009079f
C638 B.n340 VSUBS 0.009079f
C639 B.n341 VSUBS 0.009079f
C640 B.n342 VSUBS 0.009079f
C641 B.n343 VSUBS 0.009079f
C642 B.n344 VSUBS 0.009079f
C643 B.n345 VSUBS 0.009079f
C644 B.n346 VSUBS 0.009079f
C645 B.n347 VSUBS 0.009079f
C646 B.n348 VSUBS 0.009079f
C647 B.n349 VSUBS 0.009079f
C648 B.n350 VSUBS 0.009079f
C649 B.n351 VSUBS 0.009079f
C650 B.n352 VSUBS 0.009079f
C651 B.n353 VSUBS 0.009079f
C652 B.n354 VSUBS 0.009079f
C653 B.n355 VSUBS 0.009079f
C654 B.n356 VSUBS 0.009079f
C655 B.n357 VSUBS 0.009079f
C656 B.n358 VSUBS 0.009079f
C657 B.n359 VSUBS 0.009079f
C658 B.n360 VSUBS 0.009079f
C659 B.n361 VSUBS 0.009079f
C660 B.n362 VSUBS 0.009079f
C661 B.n363 VSUBS 0.009079f
C662 B.n364 VSUBS 0.009079f
C663 B.n365 VSUBS 0.009079f
C664 B.n366 VSUBS 0.009079f
C665 B.n367 VSUBS 0.009079f
C666 B.n368 VSUBS 0.009079f
C667 B.n369 VSUBS 0.009079f
C668 B.n370 VSUBS 0.009079f
C669 B.n371 VSUBS 0.009079f
C670 B.n372 VSUBS 0.009079f
C671 B.n373 VSUBS 0.009079f
C672 B.n374 VSUBS 0.009079f
C673 B.n375 VSUBS 0.009079f
C674 B.n376 VSUBS 0.009079f
C675 B.n377 VSUBS 0.009079f
C676 B.n378 VSUBS 0.009079f
C677 B.n379 VSUBS 0.009079f
C678 B.n380 VSUBS 0.009079f
C679 B.n381 VSUBS 0.009079f
C680 B.n382 VSUBS 0.009079f
C681 B.n383 VSUBS 0.009079f
C682 B.n384 VSUBS 0.009079f
C683 B.n385 VSUBS 0.009079f
C684 B.n386 VSUBS 0.009079f
C685 B.n387 VSUBS 0.009079f
C686 B.n388 VSUBS 0.009079f
C687 B.n389 VSUBS 0.009079f
C688 B.n390 VSUBS 0.009079f
C689 B.n391 VSUBS 0.009079f
C690 B.n392 VSUBS 0.009079f
C691 B.n393 VSUBS 0.009079f
C692 B.n394 VSUBS 0.009079f
C693 B.n395 VSUBS 0.009079f
C694 B.n396 VSUBS 0.009079f
C695 B.n397 VSUBS 0.009079f
C696 B.n398 VSUBS 0.009079f
C697 B.n399 VSUBS 0.009079f
C698 B.n400 VSUBS 0.009079f
C699 B.n401 VSUBS 0.009079f
C700 B.n402 VSUBS 0.009079f
C701 B.n403 VSUBS 0.009079f
C702 B.n404 VSUBS 0.009079f
C703 B.n405 VSUBS 0.009079f
C704 B.n406 VSUBS 0.009079f
C705 B.n407 VSUBS 0.009079f
C706 B.n408 VSUBS 0.009079f
C707 B.n409 VSUBS 0.009079f
C708 B.n410 VSUBS 0.009079f
C709 B.n411 VSUBS 0.009079f
C710 B.n412 VSUBS 0.009079f
C711 B.n413 VSUBS 0.009079f
C712 B.n414 VSUBS 0.009079f
C713 B.n415 VSUBS 0.009079f
C714 B.n416 VSUBS 0.009079f
C715 B.n417 VSUBS 0.009079f
C716 B.n418 VSUBS 0.009079f
C717 B.n419 VSUBS 0.009079f
C718 B.n420 VSUBS 0.009079f
C719 B.n421 VSUBS 0.009079f
C720 B.n422 VSUBS 0.023005f
C721 B.n423 VSUBS 0.022121f
C722 B.n424 VSUBS 0.023101f
C723 B.n425 VSUBS 0.009079f
C724 B.n426 VSUBS 0.009079f
C725 B.n427 VSUBS 0.009079f
C726 B.n428 VSUBS 0.009079f
C727 B.n429 VSUBS 0.009079f
C728 B.n430 VSUBS 0.009079f
C729 B.n431 VSUBS 0.009079f
C730 B.n432 VSUBS 0.009079f
C731 B.n433 VSUBS 0.009079f
C732 B.n434 VSUBS 0.009079f
C733 B.n435 VSUBS 0.009079f
C734 B.n436 VSUBS 0.009079f
C735 B.n437 VSUBS 0.009079f
C736 B.n438 VSUBS 0.009079f
C737 B.n439 VSUBS 0.009079f
C738 B.n440 VSUBS 0.009079f
C739 B.n441 VSUBS 0.009079f
C740 B.n442 VSUBS 0.009079f
C741 B.n443 VSUBS 0.009079f
C742 B.n444 VSUBS 0.009079f
C743 B.n445 VSUBS 0.009079f
C744 B.n446 VSUBS 0.009079f
C745 B.n447 VSUBS 0.009079f
C746 B.n448 VSUBS 0.009079f
C747 B.n449 VSUBS 0.009079f
C748 B.n450 VSUBS 0.009079f
C749 B.n451 VSUBS 0.009079f
C750 B.n452 VSUBS 0.009079f
C751 B.n453 VSUBS 0.009079f
C752 B.n454 VSUBS 0.009079f
C753 B.n455 VSUBS 0.009079f
C754 B.n456 VSUBS 0.009079f
C755 B.n457 VSUBS 0.009079f
C756 B.n458 VSUBS 0.009079f
C757 B.n459 VSUBS 0.009079f
C758 B.n460 VSUBS 0.009079f
C759 B.n461 VSUBS 0.009079f
C760 B.n462 VSUBS 0.009079f
C761 B.n463 VSUBS 0.009079f
C762 B.n464 VSUBS 0.009079f
C763 B.n465 VSUBS 0.009079f
C764 B.n466 VSUBS 0.009079f
C765 B.n467 VSUBS 0.009079f
C766 B.n468 VSUBS 0.009079f
C767 B.n469 VSUBS 0.009079f
C768 B.n470 VSUBS 0.009079f
C769 B.n471 VSUBS 0.009079f
C770 B.n472 VSUBS 0.009079f
C771 B.n473 VSUBS 0.009079f
C772 B.n474 VSUBS 0.009079f
C773 B.n475 VSUBS 0.009079f
C774 B.n476 VSUBS 0.009079f
C775 B.n477 VSUBS 0.009079f
C776 B.n478 VSUBS 0.009079f
C777 B.n479 VSUBS 0.009079f
C778 B.n480 VSUBS 0.009079f
C779 B.n481 VSUBS 0.009079f
C780 B.n482 VSUBS 0.009079f
C781 B.n483 VSUBS 0.009079f
C782 B.n484 VSUBS 0.009079f
C783 B.n485 VSUBS 0.009079f
C784 B.n486 VSUBS 0.009079f
C785 B.n487 VSUBS 0.009079f
C786 B.n488 VSUBS 0.009079f
C787 B.n489 VSUBS 0.009079f
C788 B.n490 VSUBS 0.009079f
C789 B.n491 VSUBS 0.009079f
C790 B.n492 VSUBS 0.009079f
C791 B.n493 VSUBS 0.009079f
C792 B.n494 VSUBS 0.009079f
C793 B.n495 VSUBS 0.009079f
C794 B.n496 VSUBS 0.009079f
C795 B.n497 VSUBS 0.009079f
C796 B.n498 VSUBS 0.009079f
C797 B.n499 VSUBS 0.009079f
C798 B.n500 VSUBS 0.009079f
C799 B.n501 VSUBS 0.009079f
C800 B.n502 VSUBS 0.009079f
C801 B.n503 VSUBS 0.022121f
C802 B.n504 VSUBS 0.023005f
C803 B.n505 VSUBS 0.023005f
C804 B.n506 VSUBS 0.009079f
C805 B.n507 VSUBS 0.009079f
C806 B.n508 VSUBS 0.009079f
C807 B.n509 VSUBS 0.009079f
C808 B.n510 VSUBS 0.009079f
C809 B.n511 VSUBS 0.009079f
C810 B.n512 VSUBS 0.009079f
C811 B.n513 VSUBS 0.009079f
C812 B.n514 VSUBS 0.009079f
C813 B.n515 VSUBS 0.009079f
C814 B.n516 VSUBS 0.009079f
C815 B.n517 VSUBS 0.009079f
C816 B.n518 VSUBS 0.009079f
C817 B.n519 VSUBS 0.009079f
C818 B.n520 VSUBS 0.009079f
C819 B.n521 VSUBS 0.009079f
C820 B.n522 VSUBS 0.009079f
C821 B.n523 VSUBS 0.009079f
C822 B.n524 VSUBS 0.009079f
C823 B.n525 VSUBS 0.009079f
C824 B.n526 VSUBS 0.009079f
C825 B.n527 VSUBS 0.009079f
C826 B.n528 VSUBS 0.009079f
C827 B.n529 VSUBS 0.009079f
C828 B.n530 VSUBS 0.009079f
C829 B.n531 VSUBS 0.009079f
C830 B.n532 VSUBS 0.009079f
C831 B.n533 VSUBS 0.009079f
C832 B.n534 VSUBS 0.009079f
C833 B.n535 VSUBS 0.009079f
C834 B.n536 VSUBS 0.009079f
C835 B.n537 VSUBS 0.009079f
C836 B.n538 VSUBS 0.009079f
C837 B.n539 VSUBS 0.009079f
C838 B.n540 VSUBS 0.009079f
C839 B.n541 VSUBS 0.009079f
C840 B.n542 VSUBS 0.009079f
C841 B.n543 VSUBS 0.009079f
C842 B.n544 VSUBS 0.009079f
C843 B.n545 VSUBS 0.009079f
C844 B.n546 VSUBS 0.009079f
C845 B.n547 VSUBS 0.009079f
C846 B.n548 VSUBS 0.009079f
C847 B.n549 VSUBS 0.009079f
C848 B.n550 VSUBS 0.009079f
C849 B.n551 VSUBS 0.009079f
C850 B.n552 VSUBS 0.009079f
C851 B.n553 VSUBS 0.009079f
C852 B.n554 VSUBS 0.009079f
C853 B.n555 VSUBS 0.009079f
C854 B.n556 VSUBS 0.009079f
C855 B.n557 VSUBS 0.009079f
C856 B.n558 VSUBS 0.009079f
C857 B.n559 VSUBS 0.009079f
C858 B.n560 VSUBS 0.009079f
C859 B.n561 VSUBS 0.009079f
C860 B.n562 VSUBS 0.009079f
C861 B.n563 VSUBS 0.009079f
C862 B.n564 VSUBS 0.009079f
C863 B.n565 VSUBS 0.009079f
C864 B.n566 VSUBS 0.009079f
C865 B.n567 VSUBS 0.009079f
C866 B.n568 VSUBS 0.009079f
C867 B.n569 VSUBS 0.009079f
C868 B.n570 VSUBS 0.009079f
C869 B.n571 VSUBS 0.009079f
C870 B.n572 VSUBS 0.009079f
C871 B.n573 VSUBS 0.009079f
C872 B.n574 VSUBS 0.009079f
C873 B.n575 VSUBS 0.009079f
C874 B.n576 VSUBS 0.009079f
C875 B.n577 VSUBS 0.009079f
C876 B.n578 VSUBS 0.009079f
C877 B.n579 VSUBS 0.009079f
C878 B.n580 VSUBS 0.009079f
C879 B.n581 VSUBS 0.009079f
C880 B.n582 VSUBS 0.009079f
C881 B.n583 VSUBS 0.009079f
C882 B.n584 VSUBS 0.009079f
C883 B.n585 VSUBS 0.009079f
C884 B.n586 VSUBS 0.009079f
C885 B.n587 VSUBS 0.009079f
C886 B.n588 VSUBS 0.009079f
C887 B.n589 VSUBS 0.009079f
C888 B.n590 VSUBS 0.009079f
C889 B.n591 VSUBS 0.009079f
C890 B.n592 VSUBS 0.008545f
C891 B.n593 VSUBS 0.021034f
C892 B.n594 VSUBS 0.005073f
C893 B.n595 VSUBS 0.009079f
C894 B.n596 VSUBS 0.009079f
C895 B.n597 VSUBS 0.009079f
C896 B.n598 VSUBS 0.009079f
C897 B.n599 VSUBS 0.009079f
C898 B.n600 VSUBS 0.009079f
C899 B.n601 VSUBS 0.009079f
C900 B.n602 VSUBS 0.009079f
C901 B.n603 VSUBS 0.009079f
C902 B.n604 VSUBS 0.009079f
C903 B.n605 VSUBS 0.009079f
C904 B.n606 VSUBS 0.009079f
C905 B.n607 VSUBS 0.005073f
C906 B.n608 VSUBS 0.009079f
C907 B.n609 VSUBS 0.009079f
C908 B.n610 VSUBS 0.009079f
C909 B.n611 VSUBS 0.009079f
C910 B.n612 VSUBS 0.009079f
C911 B.n613 VSUBS 0.009079f
C912 B.n614 VSUBS 0.009079f
C913 B.n615 VSUBS 0.009079f
C914 B.n616 VSUBS 0.009079f
C915 B.n617 VSUBS 0.009079f
C916 B.n618 VSUBS 0.009079f
C917 B.n619 VSUBS 0.009079f
C918 B.n620 VSUBS 0.009079f
C919 B.n621 VSUBS 0.009079f
C920 B.n622 VSUBS 0.009079f
C921 B.n623 VSUBS 0.009079f
C922 B.n624 VSUBS 0.009079f
C923 B.n625 VSUBS 0.009079f
C924 B.n626 VSUBS 0.009079f
C925 B.n627 VSUBS 0.009079f
C926 B.n628 VSUBS 0.009079f
C927 B.n629 VSUBS 0.009079f
C928 B.n630 VSUBS 0.009079f
C929 B.n631 VSUBS 0.009079f
C930 B.n632 VSUBS 0.009079f
C931 B.n633 VSUBS 0.009079f
C932 B.n634 VSUBS 0.009079f
C933 B.n635 VSUBS 0.009079f
C934 B.n636 VSUBS 0.009079f
C935 B.n637 VSUBS 0.009079f
C936 B.n638 VSUBS 0.009079f
C937 B.n639 VSUBS 0.009079f
C938 B.n640 VSUBS 0.009079f
C939 B.n641 VSUBS 0.009079f
C940 B.n642 VSUBS 0.009079f
C941 B.n643 VSUBS 0.009079f
C942 B.n644 VSUBS 0.009079f
C943 B.n645 VSUBS 0.009079f
C944 B.n646 VSUBS 0.009079f
C945 B.n647 VSUBS 0.009079f
C946 B.n648 VSUBS 0.009079f
C947 B.n649 VSUBS 0.009079f
C948 B.n650 VSUBS 0.009079f
C949 B.n651 VSUBS 0.009079f
C950 B.n652 VSUBS 0.009079f
C951 B.n653 VSUBS 0.009079f
C952 B.n654 VSUBS 0.009079f
C953 B.n655 VSUBS 0.009079f
C954 B.n656 VSUBS 0.009079f
C955 B.n657 VSUBS 0.009079f
C956 B.n658 VSUBS 0.009079f
C957 B.n659 VSUBS 0.009079f
C958 B.n660 VSUBS 0.009079f
C959 B.n661 VSUBS 0.009079f
C960 B.n662 VSUBS 0.009079f
C961 B.n663 VSUBS 0.009079f
C962 B.n664 VSUBS 0.009079f
C963 B.n665 VSUBS 0.009079f
C964 B.n666 VSUBS 0.009079f
C965 B.n667 VSUBS 0.009079f
C966 B.n668 VSUBS 0.009079f
C967 B.n669 VSUBS 0.009079f
C968 B.n670 VSUBS 0.009079f
C969 B.n671 VSUBS 0.009079f
C970 B.n672 VSUBS 0.009079f
C971 B.n673 VSUBS 0.009079f
C972 B.n674 VSUBS 0.009079f
C973 B.n675 VSUBS 0.009079f
C974 B.n676 VSUBS 0.009079f
C975 B.n677 VSUBS 0.009079f
C976 B.n678 VSUBS 0.009079f
C977 B.n679 VSUBS 0.009079f
C978 B.n680 VSUBS 0.009079f
C979 B.n681 VSUBS 0.009079f
C980 B.n682 VSUBS 0.009079f
C981 B.n683 VSUBS 0.009079f
C982 B.n684 VSUBS 0.009079f
C983 B.n685 VSUBS 0.009079f
C984 B.n686 VSUBS 0.009079f
C985 B.n687 VSUBS 0.009079f
C986 B.n688 VSUBS 0.009079f
C987 B.n689 VSUBS 0.009079f
C988 B.n690 VSUBS 0.009079f
C989 B.n691 VSUBS 0.009079f
C990 B.n692 VSUBS 0.009079f
C991 B.n693 VSUBS 0.009079f
C992 B.n694 VSUBS 0.009079f
C993 B.n695 VSUBS 0.009079f
C994 B.n696 VSUBS 0.023005f
C995 B.n697 VSUBS 0.022121f
C996 B.n698 VSUBS 0.022121f
C997 B.n699 VSUBS 0.009079f
C998 B.n700 VSUBS 0.009079f
C999 B.n701 VSUBS 0.009079f
C1000 B.n702 VSUBS 0.009079f
C1001 B.n703 VSUBS 0.009079f
C1002 B.n704 VSUBS 0.009079f
C1003 B.n705 VSUBS 0.009079f
C1004 B.n706 VSUBS 0.009079f
C1005 B.n707 VSUBS 0.009079f
C1006 B.n708 VSUBS 0.009079f
C1007 B.n709 VSUBS 0.009079f
C1008 B.n710 VSUBS 0.009079f
C1009 B.n711 VSUBS 0.009079f
C1010 B.n712 VSUBS 0.009079f
C1011 B.n713 VSUBS 0.009079f
C1012 B.n714 VSUBS 0.009079f
C1013 B.n715 VSUBS 0.009079f
C1014 B.n716 VSUBS 0.009079f
C1015 B.n717 VSUBS 0.009079f
C1016 B.n718 VSUBS 0.009079f
C1017 B.n719 VSUBS 0.009079f
C1018 B.n720 VSUBS 0.009079f
C1019 B.n721 VSUBS 0.009079f
C1020 B.n722 VSUBS 0.009079f
C1021 B.n723 VSUBS 0.009079f
C1022 B.n724 VSUBS 0.009079f
C1023 B.n725 VSUBS 0.009079f
C1024 B.n726 VSUBS 0.009079f
C1025 B.n727 VSUBS 0.009079f
C1026 B.n728 VSUBS 0.009079f
C1027 B.n729 VSUBS 0.009079f
C1028 B.n730 VSUBS 0.009079f
C1029 B.n731 VSUBS 0.009079f
C1030 B.n732 VSUBS 0.009079f
C1031 B.n733 VSUBS 0.009079f
C1032 B.n734 VSUBS 0.009079f
C1033 B.n735 VSUBS 0.011847f
C1034 B.n736 VSUBS 0.01262f
C1035 B.n737 VSUBS 0.025097f
C1036 VDD2.n0 VSUBS 0.015874f
C1037 VDD2.n1 VSUBS 0.035818f
C1038 VDD2.n2 VSUBS 0.016045f
C1039 VDD2.n3 VSUBS 0.028201f
C1040 VDD2.n4 VSUBS 0.015154f
C1041 VDD2.n5 VSUBS 0.035818f
C1042 VDD2.n6 VSUBS 0.016045f
C1043 VDD2.n7 VSUBS 0.028201f
C1044 VDD2.n8 VSUBS 0.015154f
C1045 VDD2.n9 VSUBS 0.035818f
C1046 VDD2.n10 VSUBS 0.016045f
C1047 VDD2.n11 VSUBS 0.028201f
C1048 VDD2.n12 VSUBS 0.015154f
C1049 VDD2.n13 VSUBS 0.035818f
C1050 VDD2.n14 VSUBS 0.016045f
C1051 VDD2.n15 VSUBS 0.028201f
C1052 VDD2.n16 VSUBS 0.015154f
C1053 VDD2.n17 VSUBS 0.035818f
C1054 VDD2.n18 VSUBS 0.016045f
C1055 VDD2.n19 VSUBS 0.028201f
C1056 VDD2.n20 VSUBS 0.015154f
C1057 VDD2.n21 VSUBS 0.035818f
C1058 VDD2.n22 VSUBS 0.016045f
C1059 VDD2.n23 VSUBS 0.028201f
C1060 VDD2.n24 VSUBS 0.015154f
C1061 VDD2.n25 VSUBS 0.035818f
C1062 VDD2.n26 VSUBS 0.016045f
C1063 VDD2.n27 VSUBS 0.028201f
C1064 VDD2.n28 VSUBS 0.015154f
C1065 VDD2.n29 VSUBS 0.035818f
C1066 VDD2.n30 VSUBS 0.016045f
C1067 VDD2.n31 VSUBS 0.299112f
C1068 VDD2.t1 VSUBS 0.077758f
C1069 VDD2.n32 VSUBS 0.026864f
C1070 VDD2.n33 VSUBS 0.026944f
C1071 VDD2.n34 VSUBS 0.015154f
C1072 VDD2.n35 VSUBS 2.13192f
C1073 VDD2.n36 VSUBS 0.028201f
C1074 VDD2.n37 VSUBS 0.015154f
C1075 VDD2.n38 VSUBS 0.016045f
C1076 VDD2.n39 VSUBS 0.035818f
C1077 VDD2.n40 VSUBS 0.035818f
C1078 VDD2.n41 VSUBS 0.016045f
C1079 VDD2.n42 VSUBS 0.015154f
C1080 VDD2.n43 VSUBS 0.028201f
C1081 VDD2.n44 VSUBS 0.028201f
C1082 VDD2.n45 VSUBS 0.015154f
C1083 VDD2.n46 VSUBS 0.016045f
C1084 VDD2.n47 VSUBS 0.035818f
C1085 VDD2.n48 VSUBS 0.035818f
C1086 VDD2.n49 VSUBS 0.035818f
C1087 VDD2.n50 VSUBS 0.016045f
C1088 VDD2.n51 VSUBS 0.015154f
C1089 VDD2.n52 VSUBS 0.028201f
C1090 VDD2.n53 VSUBS 0.028201f
C1091 VDD2.n54 VSUBS 0.015154f
C1092 VDD2.n55 VSUBS 0.015599f
C1093 VDD2.n56 VSUBS 0.015599f
C1094 VDD2.n57 VSUBS 0.035818f
C1095 VDD2.n58 VSUBS 0.035818f
C1096 VDD2.n59 VSUBS 0.016045f
C1097 VDD2.n60 VSUBS 0.015154f
C1098 VDD2.n61 VSUBS 0.028201f
C1099 VDD2.n62 VSUBS 0.028201f
C1100 VDD2.n63 VSUBS 0.015154f
C1101 VDD2.n64 VSUBS 0.016045f
C1102 VDD2.n65 VSUBS 0.035818f
C1103 VDD2.n66 VSUBS 0.035818f
C1104 VDD2.n67 VSUBS 0.016045f
C1105 VDD2.n68 VSUBS 0.015154f
C1106 VDD2.n69 VSUBS 0.028201f
C1107 VDD2.n70 VSUBS 0.028201f
C1108 VDD2.n71 VSUBS 0.015154f
C1109 VDD2.n72 VSUBS 0.016045f
C1110 VDD2.n73 VSUBS 0.035818f
C1111 VDD2.n74 VSUBS 0.035818f
C1112 VDD2.n75 VSUBS 0.016045f
C1113 VDD2.n76 VSUBS 0.015154f
C1114 VDD2.n77 VSUBS 0.028201f
C1115 VDD2.n78 VSUBS 0.028201f
C1116 VDD2.n79 VSUBS 0.015154f
C1117 VDD2.n80 VSUBS 0.016045f
C1118 VDD2.n81 VSUBS 0.035818f
C1119 VDD2.n82 VSUBS 0.035818f
C1120 VDD2.n83 VSUBS 0.016045f
C1121 VDD2.n84 VSUBS 0.015154f
C1122 VDD2.n85 VSUBS 0.028201f
C1123 VDD2.n86 VSUBS 0.028201f
C1124 VDD2.n87 VSUBS 0.015154f
C1125 VDD2.n88 VSUBS 0.016045f
C1126 VDD2.n89 VSUBS 0.035818f
C1127 VDD2.n90 VSUBS 0.035818f
C1128 VDD2.n91 VSUBS 0.016045f
C1129 VDD2.n92 VSUBS 0.015154f
C1130 VDD2.n93 VSUBS 0.028201f
C1131 VDD2.n94 VSUBS 0.071348f
C1132 VDD2.n95 VSUBS 0.015154f
C1133 VDD2.n96 VSUBS 0.016045f
C1134 VDD2.n97 VSUBS 0.078166f
C1135 VDD2.n98 VSUBS 0.074006f
C1136 VDD2.t6 VSUBS 0.402021f
C1137 VDD2.t8 VSUBS 0.402021f
C1138 VDD2.n99 VSUBS 3.365f
C1139 VDD2.n100 VSUBS 0.769996f
C1140 VDD2.t0 VSUBS 0.402021f
C1141 VDD2.t5 VSUBS 0.402021f
C1142 VDD2.n101 VSUBS 3.37091f
C1143 VDD2.n102 VSUBS 2.87838f
C1144 VDD2.n103 VSUBS 0.015874f
C1145 VDD2.n104 VSUBS 0.035818f
C1146 VDD2.n105 VSUBS 0.016045f
C1147 VDD2.n106 VSUBS 0.028201f
C1148 VDD2.n107 VSUBS 0.015154f
C1149 VDD2.n108 VSUBS 0.035818f
C1150 VDD2.n109 VSUBS 0.016045f
C1151 VDD2.n110 VSUBS 0.028201f
C1152 VDD2.n111 VSUBS 0.015154f
C1153 VDD2.n112 VSUBS 0.035818f
C1154 VDD2.n113 VSUBS 0.016045f
C1155 VDD2.n114 VSUBS 0.028201f
C1156 VDD2.n115 VSUBS 0.015154f
C1157 VDD2.n116 VSUBS 0.035818f
C1158 VDD2.n117 VSUBS 0.016045f
C1159 VDD2.n118 VSUBS 0.028201f
C1160 VDD2.n119 VSUBS 0.015154f
C1161 VDD2.n120 VSUBS 0.035818f
C1162 VDD2.n121 VSUBS 0.016045f
C1163 VDD2.n122 VSUBS 0.028201f
C1164 VDD2.n123 VSUBS 0.015154f
C1165 VDD2.n124 VSUBS 0.035818f
C1166 VDD2.n125 VSUBS 0.016045f
C1167 VDD2.n126 VSUBS 0.028201f
C1168 VDD2.n127 VSUBS 0.015154f
C1169 VDD2.n128 VSUBS 0.035818f
C1170 VDD2.n129 VSUBS 0.035818f
C1171 VDD2.n130 VSUBS 0.016045f
C1172 VDD2.n131 VSUBS 0.028201f
C1173 VDD2.n132 VSUBS 0.015154f
C1174 VDD2.n133 VSUBS 0.035818f
C1175 VDD2.n134 VSUBS 0.016045f
C1176 VDD2.n135 VSUBS 0.299112f
C1177 VDD2.t9 VSUBS 0.077758f
C1178 VDD2.n136 VSUBS 0.026864f
C1179 VDD2.n137 VSUBS 0.026944f
C1180 VDD2.n138 VSUBS 0.015154f
C1181 VDD2.n139 VSUBS 2.13192f
C1182 VDD2.n140 VSUBS 0.028201f
C1183 VDD2.n141 VSUBS 0.015154f
C1184 VDD2.n142 VSUBS 0.016045f
C1185 VDD2.n143 VSUBS 0.035818f
C1186 VDD2.n144 VSUBS 0.035818f
C1187 VDD2.n145 VSUBS 0.016045f
C1188 VDD2.n146 VSUBS 0.015154f
C1189 VDD2.n147 VSUBS 0.028201f
C1190 VDD2.n148 VSUBS 0.028201f
C1191 VDD2.n149 VSUBS 0.015154f
C1192 VDD2.n150 VSUBS 0.016045f
C1193 VDD2.n151 VSUBS 0.035818f
C1194 VDD2.n152 VSUBS 0.035818f
C1195 VDD2.n153 VSUBS 0.016045f
C1196 VDD2.n154 VSUBS 0.015154f
C1197 VDD2.n155 VSUBS 0.028201f
C1198 VDD2.n156 VSUBS 0.028201f
C1199 VDD2.n157 VSUBS 0.015154f
C1200 VDD2.n158 VSUBS 0.015599f
C1201 VDD2.n159 VSUBS 0.015599f
C1202 VDD2.n160 VSUBS 0.035818f
C1203 VDD2.n161 VSUBS 0.035818f
C1204 VDD2.n162 VSUBS 0.016045f
C1205 VDD2.n163 VSUBS 0.015154f
C1206 VDD2.n164 VSUBS 0.028201f
C1207 VDD2.n165 VSUBS 0.028201f
C1208 VDD2.n166 VSUBS 0.015154f
C1209 VDD2.n167 VSUBS 0.016045f
C1210 VDD2.n168 VSUBS 0.035818f
C1211 VDD2.n169 VSUBS 0.035818f
C1212 VDD2.n170 VSUBS 0.016045f
C1213 VDD2.n171 VSUBS 0.015154f
C1214 VDD2.n172 VSUBS 0.028201f
C1215 VDD2.n173 VSUBS 0.028201f
C1216 VDD2.n174 VSUBS 0.015154f
C1217 VDD2.n175 VSUBS 0.016045f
C1218 VDD2.n176 VSUBS 0.035818f
C1219 VDD2.n177 VSUBS 0.035818f
C1220 VDD2.n178 VSUBS 0.016045f
C1221 VDD2.n179 VSUBS 0.015154f
C1222 VDD2.n180 VSUBS 0.028201f
C1223 VDD2.n181 VSUBS 0.028201f
C1224 VDD2.n182 VSUBS 0.015154f
C1225 VDD2.n183 VSUBS 0.016045f
C1226 VDD2.n184 VSUBS 0.035818f
C1227 VDD2.n185 VSUBS 0.035818f
C1228 VDD2.n186 VSUBS 0.016045f
C1229 VDD2.n187 VSUBS 0.015154f
C1230 VDD2.n188 VSUBS 0.028201f
C1231 VDD2.n189 VSUBS 0.028201f
C1232 VDD2.n190 VSUBS 0.015154f
C1233 VDD2.n191 VSUBS 0.016045f
C1234 VDD2.n192 VSUBS 0.035818f
C1235 VDD2.n193 VSUBS 0.035818f
C1236 VDD2.n194 VSUBS 0.016045f
C1237 VDD2.n195 VSUBS 0.015154f
C1238 VDD2.n196 VSUBS 0.028201f
C1239 VDD2.n197 VSUBS 0.071348f
C1240 VDD2.n198 VSUBS 0.015154f
C1241 VDD2.n199 VSUBS 0.016045f
C1242 VDD2.n200 VSUBS 0.078166f
C1243 VDD2.n201 VSUBS 0.071577f
C1244 VDD2.n202 VSUBS 2.966f
C1245 VDD2.t2 VSUBS 0.402021f
C1246 VDD2.t3 VSUBS 0.402021f
C1247 VDD2.n203 VSUBS 3.36501f
C1248 VDD2.n204 VSUBS 0.640148f
C1249 VDD2.t4 VSUBS 0.402021f
C1250 VDD2.t7 VSUBS 0.402021f
C1251 VDD2.n205 VSUBS 3.37087f
C1252 VTAIL.t17 VSUBS 0.402914f
C1253 VTAIL.t14 VSUBS 0.402914f
C1254 VTAIL.n0 VSUBS 3.2117f
C1255 VTAIL.n1 VSUBS 0.806718f
C1256 VTAIL.n2 VSUBS 0.015909f
C1257 VTAIL.n3 VSUBS 0.035898f
C1258 VTAIL.n4 VSUBS 0.016081f
C1259 VTAIL.n5 VSUBS 0.028263f
C1260 VTAIL.n6 VSUBS 0.015187f
C1261 VTAIL.n7 VSUBS 0.035898f
C1262 VTAIL.n8 VSUBS 0.016081f
C1263 VTAIL.n9 VSUBS 0.028263f
C1264 VTAIL.n10 VSUBS 0.015187f
C1265 VTAIL.n11 VSUBS 0.035898f
C1266 VTAIL.n12 VSUBS 0.016081f
C1267 VTAIL.n13 VSUBS 0.028263f
C1268 VTAIL.n14 VSUBS 0.015187f
C1269 VTAIL.n15 VSUBS 0.035898f
C1270 VTAIL.n16 VSUBS 0.016081f
C1271 VTAIL.n17 VSUBS 0.028263f
C1272 VTAIL.n18 VSUBS 0.015187f
C1273 VTAIL.n19 VSUBS 0.035898f
C1274 VTAIL.n20 VSUBS 0.016081f
C1275 VTAIL.n21 VSUBS 0.028263f
C1276 VTAIL.n22 VSUBS 0.015187f
C1277 VTAIL.n23 VSUBS 0.035898f
C1278 VTAIL.n24 VSUBS 0.016081f
C1279 VTAIL.n25 VSUBS 0.028263f
C1280 VTAIL.n26 VSUBS 0.015187f
C1281 VTAIL.n27 VSUBS 0.035898f
C1282 VTAIL.n28 VSUBS 0.016081f
C1283 VTAIL.n29 VSUBS 0.028263f
C1284 VTAIL.n30 VSUBS 0.015187f
C1285 VTAIL.n31 VSUBS 0.035898f
C1286 VTAIL.n32 VSUBS 0.016081f
C1287 VTAIL.n33 VSUBS 0.299776f
C1288 VTAIL.t7 VSUBS 0.077931f
C1289 VTAIL.n34 VSUBS 0.026923f
C1290 VTAIL.n35 VSUBS 0.027004f
C1291 VTAIL.n36 VSUBS 0.015187f
C1292 VTAIL.n37 VSUBS 2.13666f
C1293 VTAIL.n38 VSUBS 0.028263f
C1294 VTAIL.n39 VSUBS 0.015187f
C1295 VTAIL.n40 VSUBS 0.016081f
C1296 VTAIL.n41 VSUBS 0.035898f
C1297 VTAIL.n42 VSUBS 0.035898f
C1298 VTAIL.n43 VSUBS 0.016081f
C1299 VTAIL.n44 VSUBS 0.015187f
C1300 VTAIL.n45 VSUBS 0.028263f
C1301 VTAIL.n46 VSUBS 0.028263f
C1302 VTAIL.n47 VSUBS 0.015187f
C1303 VTAIL.n48 VSUBS 0.016081f
C1304 VTAIL.n49 VSUBS 0.035898f
C1305 VTAIL.n50 VSUBS 0.035898f
C1306 VTAIL.n51 VSUBS 0.035898f
C1307 VTAIL.n52 VSUBS 0.016081f
C1308 VTAIL.n53 VSUBS 0.015187f
C1309 VTAIL.n54 VSUBS 0.028263f
C1310 VTAIL.n55 VSUBS 0.028263f
C1311 VTAIL.n56 VSUBS 0.015187f
C1312 VTAIL.n57 VSUBS 0.015634f
C1313 VTAIL.n58 VSUBS 0.015634f
C1314 VTAIL.n59 VSUBS 0.035898f
C1315 VTAIL.n60 VSUBS 0.035898f
C1316 VTAIL.n61 VSUBS 0.016081f
C1317 VTAIL.n62 VSUBS 0.015187f
C1318 VTAIL.n63 VSUBS 0.028263f
C1319 VTAIL.n64 VSUBS 0.028263f
C1320 VTAIL.n65 VSUBS 0.015187f
C1321 VTAIL.n66 VSUBS 0.016081f
C1322 VTAIL.n67 VSUBS 0.035898f
C1323 VTAIL.n68 VSUBS 0.035898f
C1324 VTAIL.n69 VSUBS 0.016081f
C1325 VTAIL.n70 VSUBS 0.015187f
C1326 VTAIL.n71 VSUBS 0.028263f
C1327 VTAIL.n72 VSUBS 0.028263f
C1328 VTAIL.n73 VSUBS 0.015187f
C1329 VTAIL.n74 VSUBS 0.016081f
C1330 VTAIL.n75 VSUBS 0.035898f
C1331 VTAIL.n76 VSUBS 0.035898f
C1332 VTAIL.n77 VSUBS 0.016081f
C1333 VTAIL.n78 VSUBS 0.015187f
C1334 VTAIL.n79 VSUBS 0.028263f
C1335 VTAIL.n80 VSUBS 0.028263f
C1336 VTAIL.n81 VSUBS 0.015187f
C1337 VTAIL.n82 VSUBS 0.016081f
C1338 VTAIL.n83 VSUBS 0.035898f
C1339 VTAIL.n84 VSUBS 0.035898f
C1340 VTAIL.n85 VSUBS 0.016081f
C1341 VTAIL.n86 VSUBS 0.015187f
C1342 VTAIL.n87 VSUBS 0.028263f
C1343 VTAIL.n88 VSUBS 0.028263f
C1344 VTAIL.n89 VSUBS 0.015187f
C1345 VTAIL.n90 VSUBS 0.016081f
C1346 VTAIL.n91 VSUBS 0.035898f
C1347 VTAIL.n92 VSUBS 0.035898f
C1348 VTAIL.n93 VSUBS 0.016081f
C1349 VTAIL.n94 VSUBS 0.015187f
C1350 VTAIL.n95 VSUBS 0.028263f
C1351 VTAIL.n96 VSUBS 0.071507f
C1352 VTAIL.n97 VSUBS 0.015187f
C1353 VTAIL.n98 VSUBS 0.016081f
C1354 VTAIL.n99 VSUBS 0.07834f
C1355 VTAIL.n100 VSUBS 0.052249f
C1356 VTAIL.n101 VSUBS 0.19276f
C1357 VTAIL.t3 VSUBS 0.402914f
C1358 VTAIL.t0 VSUBS 0.402914f
C1359 VTAIL.n102 VSUBS 3.2117f
C1360 VTAIL.n103 VSUBS 0.820457f
C1361 VTAIL.t2 VSUBS 0.402914f
C1362 VTAIL.t1 VSUBS 0.402914f
C1363 VTAIL.n104 VSUBS 3.2117f
C1364 VTAIL.n105 VSUBS 2.70312f
C1365 VTAIL.t15 VSUBS 0.402914f
C1366 VTAIL.t11 VSUBS 0.402914f
C1367 VTAIL.n106 VSUBS 3.21172f
C1368 VTAIL.n107 VSUBS 2.7031f
C1369 VTAIL.t10 VSUBS 0.402914f
C1370 VTAIL.t12 VSUBS 0.402914f
C1371 VTAIL.n108 VSUBS 3.21172f
C1372 VTAIL.n109 VSUBS 0.820444f
C1373 VTAIL.n110 VSUBS 0.015909f
C1374 VTAIL.n111 VSUBS 0.035898f
C1375 VTAIL.n112 VSUBS 0.016081f
C1376 VTAIL.n113 VSUBS 0.028263f
C1377 VTAIL.n114 VSUBS 0.015187f
C1378 VTAIL.n115 VSUBS 0.035898f
C1379 VTAIL.n116 VSUBS 0.016081f
C1380 VTAIL.n117 VSUBS 0.028263f
C1381 VTAIL.n118 VSUBS 0.015187f
C1382 VTAIL.n119 VSUBS 0.035898f
C1383 VTAIL.n120 VSUBS 0.016081f
C1384 VTAIL.n121 VSUBS 0.028263f
C1385 VTAIL.n122 VSUBS 0.015187f
C1386 VTAIL.n123 VSUBS 0.035898f
C1387 VTAIL.n124 VSUBS 0.016081f
C1388 VTAIL.n125 VSUBS 0.028263f
C1389 VTAIL.n126 VSUBS 0.015187f
C1390 VTAIL.n127 VSUBS 0.035898f
C1391 VTAIL.n128 VSUBS 0.016081f
C1392 VTAIL.n129 VSUBS 0.028263f
C1393 VTAIL.n130 VSUBS 0.015187f
C1394 VTAIL.n131 VSUBS 0.035898f
C1395 VTAIL.n132 VSUBS 0.016081f
C1396 VTAIL.n133 VSUBS 0.028263f
C1397 VTAIL.n134 VSUBS 0.015187f
C1398 VTAIL.n135 VSUBS 0.035898f
C1399 VTAIL.n136 VSUBS 0.035898f
C1400 VTAIL.n137 VSUBS 0.016081f
C1401 VTAIL.n138 VSUBS 0.028263f
C1402 VTAIL.n139 VSUBS 0.015187f
C1403 VTAIL.n140 VSUBS 0.035898f
C1404 VTAIL.n141 VSUBS 0.016081f
C1405 VTAIL.n142 VSUBS 0.299776f
C1406 VTAIL.t13 VSUBS 0.077931f
C1407 VTAIL.n143 VSUBS 0.026923f
C1408 VTAIL.n144 VSUBS 0.027004f
C1409 VTAIL.n145 VSUBS 0.015187f
C1410 VTAIL.n146 VSUBS 2.13666f
C1411 VTAIL.n147 VSUBS 0.028263f
C1412 VTAIL.n148 VSUBS 0.015187f
C1413 VTAIL.n149 VSUBS 0.016081f
C1414 VTAIL.n150 VSUBS 0.035898f
C1415 VTAIL.n151 VSUBS 0.035898f
C1416 VTAIL.n152 VSUBS 0.016081f
C1417 VTAIL.n153 VSUBS 0.015187f
C1418 VTAIL.n154 VSUBS 0.028263f
C1419 VTAIL.n155 VSUBS 0.028263f
C1420 VTAIL.n156 VSUBS 0.015187f
C1421 VTAIL.n157 VSUBS 0.016081f
C1422 VTAIL.n158 VSUBS 0.035898f
C1423 VTAIL.n159 VSUBS 0.035898f
C1424 VTAIL.n160 VSUBS 0.016081f
C1425 VTAIL.n161 VSUBS 0.015187f
C1426 VTAIL.n162 VSUBS 0.028263f
C1427 VTAIL.n163 VSUBS 0.028263f
C1428 VTAIL.n164 VSUBS 0.015187f
C1429 VTAIL.n165 VSUBS 0.015634f
C1430 VTAIL.n166 VSUBS 0.015634f
C1431 VTAIL.n167 VSUBS 0.035898f
C1432 VTAIL.n168 VSUBS 0.035898f
C1433 VTAIL.n169 VSUBS 0.016081f
C1434 VTAIL.n170 VSUBS 0.015187f
C1435 VTAIL.n171 VSUBS 0.028263f
C1436 VTAIL.n172 VSUBS 0.028263f
C1437 VTAIL.n173 VSUBS 0.015187f
C1438 VTAIL.n174 VSUBS 0.016081f
C1439 VTAIL.n175 VSUBS 0.035898f
C1440 VTAIL.n176 VSUBS 0.035898f
C1441 VTAIL.n177 VSUBS 0.016081f
C1442 VTAIL.n178 VSUBS 0.015187f
C1443 VTAIL.n179 VSUBS 0.028263f
C1444 VTAIL.n180 VSUBS 0.028263f
C1445 VTAIL.n181 VSUBS 0.015187f
C1446 VTAIL.n182 VSUBS 0.016081f
C1447 VTAIL.n183 VSUBS 0.035898f
C1448 VTAIL.n184 VSUBS 0.035898f
C1449 VTAIL.n185 VSUBS 0.016081f
C1450 VTAIL.n186 VSUBS 0.015187f
C1451 VTAIL.n187 VSUBS 0.028263f
C1452 VTAIL.n188 VSUBS 0.028263f
C1453 VTAIL.n189 VSUBS 0.015187f
C1454 VTAIL.n190 VSUBS 0.016081f
C1455 VTAIL.n191 VSUBS 0.035898f
C1456 VTAIL.n192 VSUBS 0.035898f
C1457 VTAIL.n193 VSUBS 0.016081f
C1458 VTAIL.n194 VSUBS 0.015187f
C1459 VTAIL.n195 VSUBS 0.028263f
C1460 VTAIL.n196 VSUBS 0.028263f
C1461 VTAIL.n197 VSUBS 0.015187f
C1462 VTAIL.n198 VSUBS 0.016081f
C1463 VTAIL.n199 VSUBS 0.035898f
C1464 VTAIL.n200 VSUBS 0.035898f
C1465 VTAIL.n201 VSUBS 0.016081f
C1466 VTAIL.n202 VSUBS 0.015187f
C1467 VTAIL.n203 VSUBS 0.028263f
C1468 VTAIL.n204 VSUBS 0.071507f
C1469 VTAIL.n205 VSUBS 0.015187f
C1470 VTAIL.n206 VSUBS 0.016081f
C1471 VTAIL.n207 VSUBS 0.07834f
C1472 VTAIL.n208 VSUBS 0.052249f
C1473 VTAIL.n209 VSUBS 0.19276f
C1474 VTAIL.t4 VSUBS 0.402914f
C1475 VTAIL.t6 VSUBS 0.402914f
C1476 VTAIL.n210 VSUBS 3.21172f
C1477 VTAIL.n211 VSUBS 0.822014f
C1478 VTAIL.t18 VSUBS 0.402914f
C1479 VTAIL.t5 VSUBS 0.402914f
C1480 VTAIL.n212 VSUBS 3.21172f
C1481 VTAIL.n213 VSUBS 0.820444f
C1482 VTAIL.n214 VSUBS 0.015909f
C1483 VTAIL.n215 VSUBS 0.035898f
C1484 VTAIL.n216 VSUBS 0.016081f
C1485 VTAIL.n217 VSUBS 0.028263f
C1486 VTAIL.n218 VSUBS 0.015187f
C1487 VTAIL.n219 VSUBS 0.035898f
C1488 VTAIL.n220 VSUBS 0.016081f
C1489 VTAIL.n221 VSUBS 0.028263f
C1490 VTAIL.n222 VSUBS 0.015187f
C1491 VTAIL.n223 VSUBS 0.035898f
C1492 VTAIL.n224 VSUBS 0.016081f
C1493 VTAIL.n225 VSUBS 0.028263f
C1494 VTAIL.n226 VSUBS 0.015187f
C1495 VTAIL.n227 VSUBS 0.035898f
C1496 VTAIL.n228 VSUBS 0.016081f
C1497 VTAIL.n229 VSUBS 0.028263f
C1498 VTAIL.n230 VSUBS 0.015187f
C1499 VTAIL.n231 VSUBS 0.035898f
C1500 VTAIL.n232 VSUBS 0.016081f
C1501 VTAIL.n233 VSUBS 0.028263f
C1502 VTAIL.n234 VSUBS 0.015187f
C1503 VTAIL.n235 VSUBS 0.035898f
C1504 VTAIL.n236 VSUBS 0.016081f
C1505 VTAIL.n237 VSUBS 0.028263f
C1506 VTAIL.n238 VSUBS 0.015187f
C1507 VTAIL.n239 VSUBS 0.035898f
C1508 VTAIL.n240 VSUBS 0.035898f
C1509 VTAIL.n241 VSUBS 0.016081f
C1510 VTAIL.n242 VSUBS 0.028263f
C1511 VTAIL.n243 VSUBS 0.015187f
C1512 VTAIL.n244 VSUBS 0.035898f
C1513 VTAIL.n245 VSUBS 0.016081f
C1514 VTAIL.n246 VSUBS 0.299776f
C1515 VTAIL.t19 VSUBS 0.077931f
C1516 VTAIL.n247 VSUBS 0.026923f
C1517 VTAIL.n248 VSUBS 0.027004f
C1518 VTAIL.n249 VSUBS 0.015187f
C1519 VTAIL.n250 VSUBS 2.13666f
C1520 VTAIL.n251 VSUBS 0.028263f
C1521 VTAIL.n252 VSUBS 0.015187f
C1522 VTAIL.n253 VSUBS 0.016081f
C1523 VTAIL.n254 VSUBS 0.035898f
C1524 VTAIL.n255 VSUBS 0.035898f
C1525 VTAIL.n256 VSUBS 0.016081f
C1526 VTAIL.n257 VSUBS 0.015187f
C1527 VTAIL.n258 VSUBS 0.028263f
C1528 VTAIL.n259 VSUBS 0.028263f
C1529 VTAIL.n260 VSUBS 0.015187f
C1530 VTAIL.n261 VSUBS 0.016081f
C1531 VTAIL.n262 VSUBS 0.035898f
C1532 VTAIL.n263 VSUBS 0.035898f
C1533 VTAIL.n264 VSUBS 0.016081f
C1534 VTAIL.n265 VSUBS 0.015187f
C1535 VTAIL.n266 VSUBS 0.028263f
C1536 VTAIL.n267 VSUBS 0.028263f
C1537 VTAIL.n268 VSUBS 0.015187f
C1538 VTAIL.n269 VSUBS 0.015634f
C1539 VTAIL.n270 VSUBS 0.015634f
C1540 VTAIL.n271 VSUBS 0.035898f
C1541 VTAIL.n272 VSUBS 0.035898f
C1542 VTAIL.n273 VSUBS 0.016081f
C1543 VTAIL.n274 VSUBS 0.015187f
C1544 VTAIL.n275 VSUBS 0.028263f
C1545 VTAIL.n276 VSUBS 0.028263f
C1546 VTAIL.n277 VSUBS 0.015187f
C1547 VTAIL.n278 VSUBS 0.016081f
C1548 VTAIL.n279 VSUBS 0.035898f
C1549 VTAIL.n280 VSUBS 0.035898f
C1550 VTAIL.n281 VSUBS 0.016081f
C1551 VTAIL.n282 VSUBS 0.015187f
C1552 VTAIL.n283 VSUBS 0.028263f
C1553 VTAIL.n284 VSUBS 0.028263f
C1554 VTAIL.n285 VSUBS 0.015187f
C1555 VTAIL.n286 VSUBS 0.016081f
C1556 VTAIL.n287 VSUBS 0.035898f
C1557 VTAIL.n288 VSUBS 0.035898f
C1558 VTAIL.n289 VSUBS 0.016081f
C1559 VTAIL.n290 VSUBS 0.015187f
C1560 VTAIL.n291 VSUBS 0.028263f
C1561 VTAIL.n292 VSUBS 0.028263f
C1562 VTAIL.n293 VSUBS 0.015187f
C1563 VTAIL.n294 VSUBS 0.016081f
C1564 VTAIL.n295 VSUBS 0.035898f
C1565 VTAIL.n296 VSUBS 0.035898f
C1566 VTAIL.n297 VSUBS 0.016081f
C1567 VTAIL.n298 VSUBS 0.015187f
C1568 VTAIL.n299 VSUBS 0.028263f
C1569 VTAIL.n300 VSUBS 0.028263f
C1570 VTAIL.n301 VSUBS 0.015187f
C1571 VTAIL.n302 VSUBS 0.016081f
C1572 VTAIL.n303 VSUBS 0.035898f
C1573 VTAIL.n304 VSUBS 0.035898f
C1574 VTAIL.n305 VSUBS 0.016081f
C1575 VTAIL.n306 VSUBS 0.015187f
C1576 VTAIL.n307 VSUBS 0.028263f
C1577 VTAIL.n308 VSUBS 0.071507f
C1578 VTAIL.n309 VSUBS 0.015187f
C1579 VTAIL.n310 VSUBS 0.016081f
C1580 VTAIL.n311 VSUBS 0.07834f
C1581 VTAIL.n312 VSUBS 0.052249f
C1582 VTAIL.n313 VSUBS 1.99142f
C1583 VTAIL.n314 VSUBS 0.015909f
C1584 VTAIL.n315 VSUBS 0.035898f
C1585 VTAIL.n316 VSUBS 0.016081f
C1586 VTAIL.n317 VSUBS 0.028263f
C1587 VTAIL.n318 VSUBS 0.015187f
C1588 VTAIL.n319 VSUBS 0.035898f
C1589 VTAIL.n320 VSUBS 0.016081f
C1590 VTAIL.n321 VSUBS 0.028263f
C1591 VTAIL.n322 VSUBS 0.015187f
C1592 VTAIL.n323 VSUBS 0.035898f
C1593 VTAIL.n324 VSUBS 0.016081f
C1594 VTAIL.n325 VSUBS 0.028263f
C1595 VTAIL.n326 VSUBS 0.015187f
C1596 VTAIL.n327 VSUBS 0.035898f
C1597 VTAIL.n328 VSUBS 0.016081f
C1598 VTAIL.n329 VSUBS 0.028263f
C1599 VTAIL.n330 VSUBS 0.015187f
C1600 VTAIL.n331 VSUBS 0.035898f
C1601 VTAIL.n332 VSUBS 0.016081f
C1602 VTAIL.n333 VSUBS 0.028263f
C1603 VTAIL.n334 VSUBS 0.015187f
C1604 VTAIL.n335 VSUBS 0.035898f
C1605 VTAIL.n336 VSUBS 0.016081f
C1606 VTAIL.n337 VSUBS 0.028263f
C1607 VTAIL.n338 VSUBS 0.015187f
C1608 VTAIL.n339 VSUBS 0.035898f
C1609 VTAIL.n340 VSUBS 0.016081f
C1610 VTAIL.n341 VSUBS 0.028263f
C1611 VTAIL.n342 VSUBS 0.015187f
C1612 VTAIL.n343 VSUBS 0.035898f
C1613 VTAIL.n344 VSUBS 0.016081f
C1614 VTAIL.n345 VSUBS 0.299776f
C1615 VTAIL.t16 VSUBS 0.077931f
C1616 VTAIL.n346 VSUBS 0.026923f
C1617 VTAIL.n347 VSUBS 0.027004f
C1618 VTAIL.n348 VSUBS 0.015187f
C1619 VTAIL.n349 VSUBS 2.13666f
C1620 VTAIL.n350 VSUBS 0.028263f
C1621 VTAIL.n351 VSUBS 0.015187f
C1622 VTAIL.n352 VSUBS 0.016081f
C1623 VTAIL.n353 VSUBS 0.035898f
C1624 VTAIL.n354 VSUBS 0.035898f
C1625 VTAIL.n355 VSUBS 0.016081f
C1626 VTAIL.n356 VSUBS 0.015187f
C1627 VTAIL.n357 VSUBS 0.028263f
C1628 VTAIL.n358 VSUBS 0.028263f
C1629 VTAIL.n359 VSUBS 0.015187f
C1630 VTAIL.n360 VSUBS 0.016081f
C1631 VTAIL.n361 VSUBS 0.035898f
C1632 VTAIL.n362 VSUBS 0.035898f
C1633 VTAIL.n363 VSUBS 0.035898f
C1634 VTAIL.n364 VSUBS 0.016081f
C1635 VTAIL.n365 VSUBS 0.015187f
C1636 VTAIL.n366 VSUBS 0.028263f
C1637 VTAIL.n367 VSUBS 0.028263f
C1638 VTAIL.n368 VSUBS 0.015187f
C1639 VTAIL.n369 VSUBS 0.015634f
C1640 VTAIL.n370 VSUBS 0.015634f
C1641 VTAIL.n371 VSUBS 0.035898f
C1642 VTAIL.n372 VSUBS 0.035898f
C1643 VTAIL.n373 VSUBS 0.016081f
C1644 VTAIL.n374 VSUBS 0.015187f
C1645 VTAIL.n375 VSUBS 0.028263f
C1646 VTAIL.n376 VSUBS 0.028263f
C1647 VTAIL.n377 VSUBS 0.015187f
C1648 VTAIL.n378 VSUBS 0.016081f
C1649 VTAIL.n379 VSUBS 0.035898f
C1650 VTAIL.n380 VSUBS 0.035898f
C1651 VTAIL.n381 VSUBS 0.016081f
C1652 VTAIL.n382 VSUBS 0.015187f
C1653 VTAIL.n383 VSUBS 0.028263f
C1654 VTAIL.n384 VSUBS 0.028263f
C1655 VTAIL.n385 VSUBS 0.015187f
C1656 VTAIL.n386 VSUBS 0.016081f
C1657 VTAIL.n387 VSUBS 0.035898f
C1658 VTAIL.n388 VSUBS 0.035898f
C1659 VTAIL.n389 VSUBS 0.016081f
C1660 VTAIL.n390 VSUBS 0.015187f
C1661 VTAIL.n391 VSUBS 0.028263f
C1662 VTAIL.n392 VSUBS 0.028263f
C1663 VTAIL.n393 VSUBS 0.015187f
C1664 VTAIL.n394 VSUBS 0.016081f
C1665 VTAIL.n395 VSUBS 0.035898f
C1666 VTAIL.n396 VSUBS 0.035898f
C1667 VTAIL.n397 VSUBS 0.016081f
C1668 VTAIL.n398 VSUBS 0.015187f
C1669 VTAIL.n399 VSUBS 0.028263f
C1670 VTAIL.n400 VSUBS 0.028263f
C1671 VTAIL.n401 VSUBS 0.015187f
C1672 VTAIL.n402 VSUBS 0.016081f
C1673 VTAIL.n403 VSUBS 0.035898f
C1674 VTAIL.n404 VSUBS 0.035898f
C1675 VTAIL.n405 VSUBS 0.016081f
C1676 VTAIL.n406 VSUBS 0.015187f
C1677 VTAIL.n407 VSUBS 0.028263f
C1678 VTAIL.n408 VSUBS 0.071507f
C1679 VTAIL.n409 VSUBS 0.015187f
C1680 VTAIL.n410 VSUBS 0.016081f
C1681 VTAIL.n411 VSUBS 0.07834f
C1682 VTAIL.n412 VSUBS 0.052249f
C1683 VTAIL.n413 VSUBS 1.99142f
C1684 VTAIL.t9 VSUBS 0.402914f
C1685 VTAIL.t8 VSUBS 0.402914f
C1686 VTAIL.n414 VSUBS 3.2117f
C1687 VTAIL.n415 VSUBS 0.753332f
C1688 VN.n0 VSUBS 0.048733f
C1689 VN.n1 VSUBS 0.011059f
C1690 VN.n2 VSUBS 0.206525f
C1691 VN.t8 VSUBS 1.81821f
C1692 VN.n3 VSUBS 0.657119f
C1693 VN.t3 VSUBS 1.79456f
C1694 VN.n4 VSUBS 0.681958f
C1695 VN.n5 VSUBS 0.011059f
C1696 VN.t1 VSUBS 1.79456f
C1697 VN.n6 VSUBS 0.675921f
C1698 VN.n7 VSUBS 0.048733f
C1699 VN.n8 VSUBS 0.048733f
C1700 VN.n9 VSUBS 0.048733f
C1701 VN.t9 VSUBS 1.79456f
C1702 VN.n10 VSUBS 0.675921f
C1703 VN.n11 VSUBS 0.011059f
C1704 VN.t4 VSUBS 1.79456f
C1705 VN.n12 VSUBS 0.674719f
C1706 VN.n13 VSUBS 0.037766f
C1707 VN.n14 VSUBS 0.048733f
C1708 VN.n15 VSUBS 0.011059f
C1709 VN.t7 VSUBS 1.79456f
C1710 VN.n16 VSUBS 0.206525f
C1711 VN.t2 VSUBS 1.81821f
C1712 VN.n17 VSUBS 0.657119f
C1713 VN.t5 VSUBS 1.79456f
C1714 VN.n18 VSUBS 0.681958f
C1715 VN.n19 VSUBS 0.011059f
C1716 VN.t6 VSUBS 1.79456f
C1717 VN.n20 VSUBS 0.675921f
C1718 VN.n21 VSUBS 0.048733f
C1719 VN.n22 VSUBS 0.048733f
C1720 VN.n23 VSUBS 0.048733f
C1721 VN.n24 VSUBS 0.675921f
C1722 VN.n25 VSUBS 0.011059f
C1723 VN.t0 VSUBS 1.79456f
C1724 VN.n26 VSUBS 0.674719f
C1725 VN.n27 VSUBS 2.48228f
.ends

