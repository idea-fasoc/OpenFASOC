* NGSPICE file created from diff_pair_sample_1434.ext - technology: sky130A

.subckt diff_pair_sample_1434 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=0 ps=0 w=18.43 l=2.85
X1 VTAIL.t7 VN.t0 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=3.04095 ps=18.76 w=18.43 l=2.85
X2 VDD2.t1 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.04095 pd=18.76 as=7.1877 ps=37.64 w=18.43 l=2.85
X3 VTAIL.t5 VN.t2 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=3.04095 ps=18.76 w=18.43 l=2.85
X4 VTAIL.t0 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=3.04095 ps=18.76 w=18.43 l=2.85
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=0 ps=0 w=18.43 l=2.85
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=0 ps=0 w=18.43 l=2.85
X7 VDD2.t3 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.04095 pd=18.76 as=7.1877 ps=37.64 w=18.43 l=2.85
X8 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=3.04095 ps=18.76 w=18.43 l=2.85
X9 VDD1.t1 VP.t2 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.04095 pd=18.76 as=7.1877 ps=37.64 w=18.43 l=2.85
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1877 pd=37.64 as=0 ps=0 w=18.43 l=2.85
X11 VDD1.t0 VP.t3 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.04095 pd=18.76 as=7.1877 ps=37.64 w=18.43 l=2.85
R0 B.n956 B.n955 585
R1 B.n957 B.n956 585
R2 B.n397 B.n134 585
R3 B.n396 B.n395 585
R4 B.n394 B.n393 585
R5 B.n392 B.n391 585
R6 B.n390 B.n389 585
R7 B.n388 B.n387 585
R8 B.n386 B.n385 585
R9 B.n384 B.n383 585
R10 B.n382 B.n381 585
R11 B.n380 B.n379 585
R12 B.n378 B.n377 585
R13 B.n376 B.n375 585
R14 B.n374 B.n373 585
R15 B.n372 B.n371 585
R16 B.n370 B.n369 585
R17 B.n368 B.n367 585
R18 B.n366 B.n365 585
R19 B.n364 B.n363 585
R20 B.n362 B.n361 585
R21 B.n360 B.n359 585
R22 B.n358 B.n357 585
R23 B.n356 B.n355 585
R24 B.n354 B.n353 585
R25 B.n352 B.n351 585
R26 B.n350 B.n349 585
R27 B.n348 B.n347 585
R28 B.n346 B.n345 585
R29 B.n344 B.n343 585
R30 B.n342 B.n341 585
R31 B.n340 B.n339 585
R32 B.n338 B.n337 585
R33 B.n336 B.n335 585
R34 B.n334 B.n333 585
R35 B.n332 B.n331 585
R36 B.n330 B.n329 585
R37 B.n328 B.n327 585
R38 B.n326 B.n325 585
R39 B.n324 B.n323 585
R40 B.n322 B.n321 585
R41 B.n320 B.n319 585
R42 B.n318 B.n317 585
R43 B.n316 B.n315 585
R44 B.n314 B.n313 585
R45 B.n312 B.n311 585
R46 B.n310 B.n309 585
R47 B.n308 B.n307 585
R48 B.n306 B.n305 585
R49 B.n304 B.n303 585
R50 B.n302 B.n301 585
R51 B.n300 B.n299 585
R52 B.n298 B.n297 585
R53 B.n296 B.n295 585
R54 B.n294 B.n293 585
R55 B.n292 B.n291 585
R56 B.n290 B.n289 585
R57 B.n288 B.n287 585
R58 B.n286 B.n285 585
R59 B.n284 B.n283 585
R60 B.n282 B.n281 585
R61 B.n280 B.n279 585
R62 B.n278 B.n277 585
R63 B.n276 B.n275 585
R64 B.n274 B.n273 585
R65 B.n272 B.n271 585
R66 B.n270 B.n269 585
R67 B.n268 B.n267 585
R68 B.n266 B.n265 585
R69 B.n264 B.n263 585
R70 B.n262 B.n261 585
R71 B.n259 B.n258 585
R72 B.n257 B.n256 585
R73 B.n255 B.n254 585
R74 B.n253 B.n252 585
R75 B.n251 B.n250 585
R76 B.n249 B.n248 585
R77 B.n247 B.n246 585
R78 B.n245 B.n244 585
R79 B.n243 B.n242 585
R80 B.n241 B.n240 585
R81 B.n239 B.n238 585
R82 B.n237 B.n236 585
R83 B.n235 B.n234 585
R84 B.n233 B.n232 585
R85 B.n231 B.n230 585
R86 B.n229 B.n228 585
R87 B.n227 B.n226 585
R88 B.n225 B.n224 585
R89 B.n223 B.n222 585
R90 B.n221 B.n220 585
R91 B.n219 B.n218 585
R92 B.n217 B.n216 585
R93 B.n215 B.n214 585
R94 B.n213 B.n212 585
R95 B.n211 B.n210 585
R96 B.n209 B.n208 585
R97 B.n207 B.n206 585
R98 B.n205 B.n204 585
R99 B.n203 B.n202 585
R100 B.n201 B.n200 585
R101 B.n199 B.n198 585
R102 B.n197 B.n196 585
R103 B.n195 B.n194 585
R104 B.n193 B.n192 585
R105 B.n191 B.n190 585
R106 B.n189 B.n188 585
R107 B.n187 B.n186 585
R108 B.n185 B.n184 585
R109 B.n183 B.n182 585
R110 B.n181 B.n180 585
R111 B.n179 B.n178 585
R112 B.n177 B.n176 585
R113 B.n175 B.n174 585
R114 B.n173 B.n172 585
R115 B.n171 B.n170 585
R116 B.n169 B.n168 585
R117 B.n167 B.n166 585
R118 B.n165 B.n164 585
R119 B.n163 B.n162 585
R120 B.n161 B.n160 585
R121 B.n159 B.n158 585
R122 B.n157 B.n156 585
R123 B.n155 B.n154 585
R124 B.n153 B.n152 585
R125 B.n151 B.n150 585
R126 B.n149 B.n148 585
R127 B.n147 B.n146 585
R128 B.n145 B.n144 585
R129 B.n143 B.n142 585
R130 B.n141 B.n140 585
R131 B.n67 B.n66 585
R132 B.n954 B.n68 585
R133 B.n958 B.n68 585
R134 B.n953 B.n952 585
R135 B.n952 B.n64 585
R136 B.n951 B.n63 585
R137 B.n964 B.n63 585
R138 B.n950 B.n62 585
R139 B.n965 B.n62 585
R140 B.n949 B.n61 585
R141 B.n966 B.n61 585
R142 B.n948 B.n947 585
R143 B.n947 B.n57 585
R144 B.n946 B.n56 585
R145 B.n972 B.n56 585
R146 B.n945 B.n55 585
R147 B.n973 B.n55 585
R148 B.n944 B.n54 585
R149 B.n974 B.n54 585
R150 B.n943 B.n942 585
R151 B.n942 B.n50 585
R152 B.n941 B.n49 585
R153 B.n980 B.n49 585
R154 B.n940 B.n48 585
R155 B.n981 B.n48 585
R156 B.n939 B.n47 585
R157 B.n982 B.n47 585
R158 B.n938 B.n937 585
R159 B.n937 B.n43 585
R160 B.n936 B.n42 585
R161 B.n988 B.n42 585
R162 B.n935 B.n41 585
R163 B.n989 B.n41 585
R164 B.n934 B.n40 585
R165 B.n990 B.n40 585
R166 B.n933 B.n932 585
R167 B.n932 B.n36 585
R168 B.n931 B.n35 585
R169 B.n996 B.n35 585
R170 B.n930 B.n34 585
R171 B.n997 B.n34 585
R172 B.n929 B.n33 585
R173 B.n998 B.n33 585
R174 B.n928 B.n927 585
R175 B.n927 B.n29 585
R176 B.n926 B.n28 585
R177 B.n1004 B.n28 585
R178 B.n925 B.n27 585
R179 B.n1005 B.n27 585
R180 B.n924 B.n26 585
R181 B.n1006 B.n26 585
R182 B.n923 B.n922 585
R183 B.n922 B.n22 585
R184 B.n921 B.n21 585
R185 B.n1012 B.n21 585
R186 B.n920 B.n20 585
R187 B.n1013 B.n20 585
R188 B.n919 B.n19 585
R189 B.n1014 B.n19 585
R190 B.n918 B.n917 585
R191 B.n917 B.n18 585
R192 B.n916 B.n14 585
R193 B.n1020 B.n14 585
R194 B.n915 B.n13 585
R195 B.n1021 B.n13 585
R196 B.n914 B.n12 585
R197 B.n1022 B.n12 585
R198 B.n913 B.n912 585
R199 B.n912 B.n8 585
R200 B.n911 B.n7 585
R201 B.n1028 B.n7 585
R202 B.n910 B.n6 585
R203 B.n1029 B.n6 585
R204 B.n909 B.n5 585
R205 B.n1030 B.n5 585
R206 B.n908 B.n907 585
R207 B.n907 B.n4 585
R208 B.n906 B.n398 585
R209 B.n906 B.n905 585
R210 B.n896 B.n399 585
R211 B.n400 B.n399 585
R212 B.n898 B.n897 585
R213 B.n899 B.n898 585
R214 B.n895 B.n405 585
R215 B.n405 B.n404 585
R216 B.n894 B.n893 585
R217 B.n893 B.n892 585
R218 B.n407 B.n406 585
R219 B.n885 B.n407 585
R220 B.n884 B.n883 585
R221 B.n886 B.n884 585
R222 B.n882 B.n412 585
R223 B.n412 B.n411 585
R224 B.n881 B.n880 585
R225 B.n880 B.n879 585
R226 B.n414 B.n413 585
R227 B.n415 B.n414 585
R228 B.n872 B.n871 585
R229 B.n873 B.n872 585
R230 B.n870 B.n420 585
R231 B.n420 B.n419 585
R232 B.n869 B.n868 585
R233 B.n868 B.n867 585
R234 B.n422 B.n421 585
R235 B.n423 B.n422 585
R236 B.n860 B.n859 585
R237 B.n861 B.n860 585
R238 B.n858 B.n428 585
R239 B.n428 B.n427 585
R240 B.n857 B.n856 585
R241 B.n856 B.n855 585
R242 B.n430 B.n429 585
R243 B.n431 B.n430 585
R244 B.n848 B.n847 585
R245 B.n849 B.n848 585
R246 B.n846 B.n436 585
R247 B.n436 B.n435 585
R248 B.n845 B.n844 585
R249 B.n844 B.n843 585
R250 B.n438 B.n437 585
R251 B.n439 B.n438 585
R252 B.n836 B.n835 585
R253 B.n837 B.n836 585
R254 B.n834 B.n444 585
R255 B.n444 B.n443 585
R256 B.n833 B.n832 585
R257 B.n832 B.n831 585
R258 B.n446 B.n445 585
R259 B.n447 B.n446 585
R260 B.n824 B.n823 585
R261 B.n825 B.n824 585
R262 B.n822 B.n451 585
R263 B.n455 B.n451 585
R264 B.n821 B.n820 585
R265 B.n820 B.n819 585
R266 B.n453 B.n452 585
R267 B.n454 B.n453 585
R268 B.n812 B.n811 585
R269 B.n813 B.n812 585
R270 B.n810 B.n460 585
R271 B.n460 B.n459 585
R272 B.n809 B.n808 585
R273 B.n808 B.n807 585
R274 B.n462 B.n461 585
R275 B.n463 B.n462 585
R276 B.n800 B.n799 585
R277 B.n801 B.n800 585
R278 B.n466 B.n465 585
R279 B.n540 B.n539 585
R280 B.n541 B.n537 585
R281 B.n537 B.n467 585
R282 B.n543 B.n542 585
R283 B.n545 B.n536 585
R284 B.n548 B.n547 585
R285 B.n549 B.n535 585
R286 B.n551 B.n550 585
R287 B.n553 B.n534 585
R288 B.n556 B.n555 585
R289 B.n557 B.n533 585
R290 B.n559 B.n558 585
R291 B.n561 B.n532 585
R292 B.n564 B.n563 585
R293 B.n565 B.n531 585
R294 B.n567 B.n566 585
R295 B.n569 B.n530 585
R296 B.n572 B.n571 585
R297 B.n573 B.n529 585
R298 B.n575 B.n574 585
R299 B.n577 B.n528 585
R300 B.n580 B.n579 585
R301 B.n581 B.n527 585
R302 B.n583 B.n582 585
R303 B.n585 B.n526 585
R304 B.n588 B.n587 585
R305 B.n589 B.n525 585
R306 B.n591 B.n590 585
R307 B.n593 B.n524 585
R308 B.n596 B.n595 585
R309 B.n597 B.n523 585
R310 B.n599 B.n598 585
R311 B.n601 B.n522 585
R312 B.n604 B.n603 585
R313 B.n605 B.n521 585
R314 B.n607 B.n606 585
R315 B.n609 B.n520 585
R316 B.n612 B.n611 585
R317 B.n613 B.n519 585
R318 B.n615 B.n614 585
R319 B.n617 B.n518 585
R320 B.n620 B.n619 585
R321 B.n621 B.n517 585
R322 B.n623 B.n622 585
R323 B.n625 B.n516 585
R324 B.n628 B.n627 585
R325 B.n629 B.n515 585
R326 B.n631 B.n630 585
R327 B.n633 B.n514 585
R328 B.n636 B.n635 585
R329 B.n637 B.n513 585
R330 B.n639 B.n638 585
R331 B.n641 B.n512 585
R332 B.n644 B.n643 585
R333 B.n645 B.n511 585
R334 B.n647 B.n646 585
R335 B.n649 B.n510 585
R336 B.n652 B.n651 585
R337 B.n653 B.n509 585
R338 B.n655 B.n654 585
R339 B.n657 B.n508 585
R340 B.n660 B.n659 585
R341 B.n661 B.n504 585
R342 B.n663 B.n662 585
R343 B.n665 B.n503 585
R344 B.n668 B.n667 585
R345 B.n669 B.n502 585
R346 B.n671 B.n670 585
R347 B.n673 B.n501 585
R348 B.n676 B.n675 585
R349 B.n678 B.n498 585
R350 B.n680 B.n679 585
R351 B.n682 B.n497 585
R352 B.n685 B.n684 585
R353 B.n686 B.n496 585
R354 B.n688 B.n687 585
R355 B.n690 B.n495 585
R356 B.n693 B.n692 585
R357 B.n694 B.n494 585
R358 B.n696 B.n695 585
R359 B.n698 B.n493 585
R360 B.n701 B.n700 585
R361 B.n702 B.n492 585
R362 B.n704 B.n703 585
R363 B.n706 B.n491 585
R364 B.n709 B.n708 585
R365 B.n710 B.n490 585
R366 B.n712 B.n711 585
R367 B.n714 B.n489 585
R368 B.n717 B.n716 585
R369 B.n718 B.n488 585
R370 B.n720 B.n719 585
R371 B.n722 B.n487 585
R372 B.n725 B.n724 585
R373 B.n726 B.n486 585
R374 B.n728 B.n727 585
R375 B.n730 B.n485 585
R376 B.n733 B.n732 585
R377 B.n734 B.n484 585
R378 B.n736 B.n735 585
R379 B.n738 B.n483 585
R380 B.n741 B.n740 585
R381 B.n742 B.n482 585
R382 B.n744 B.n743 585
R383 B.n746 B.n481 585
R384 B.n749 B.n748 585
R385 B.n750 B.n480 585
R386 B.n752 B.n751 585
R387 B.n754 B.n479 585
R388 B.n757 B.n756 585
R389 B.n758 B.n478 585
R390 B.n760 B.n759 585
R391 B.n762 B.n477 585
R392 B.n765 B.n764 585
R393 B.n766 B.n476 585
R394 B.n768 B.n767 585
R395 B.n770 B.n475 585
R396 B.n773 B.n772 585
R397 B.n774 B.n474 585
R398 B.n776 B.n775 585
R399 B.n778 B.n473 585
R400 B.n781 B.n780 585
R401 B.n782 B.n472 585
R402 B.n784 B.n783 585
R403 B.n786 B.n471 585
R404 B.n789 B.n788 585
R405 B.n790 B.n470 585
R406 B.n792 B.n791 585
R407 B.n794 B.n469 585
R408 B.n797 B.n796 585
R409 B.n798 B.n468 585
R410 B.n803 B.n802 585
R411 B.n802 B.n801 585
R412 B.n804 B.n464 585
R413 B.n464 B.n463 585
R414 B.n806 B.n805 585
R415 B.n807 B.n806 585
R416 B.n458 B.n457 585
R417 B.n459 B.n458 585
R418 B.n815 B.n814 585
R419 B.n814 B.n813 585
R420 B.n816 B.n456 585
R421 B.n456 B.n454 585
R422 B.n818 B.n817 585
R423 B.n819 B.n818 585
R424 B.n450 B.n449 585
R425 B.n455 B.n450 585
R426 B.n827 B.n826 585
R427 B.n826 B.n825 585
R428 B.n828 B.n448 585
R429 B.n448 B.n447 585
R430 B.n830 B.n829 585
R431 B.n831 B.n830 585
R432 B.n442 B.n441 585
R433 B.n443 B.n442 585
R434 B.n839 B.n838 585
R435 B.n838 B.n837 585
R436 B.n840 B.n440 585
R437 B.n440 B.n439 585
R438 B.n842 B.n841 585
R439 B.n843 B.n842 585
R440 B.n434 B.n433 585
R441 B.n435 B.n434 585
R442 B.n851 B.n850 585
R443 B.n850 B.n849 585
R444 B.n852 B.n432 585
R445 B.n432 B.n431 585
R446 B.n854 B.n853 585
R447 B.n855 B.n854 585
R448 B.n426 B.n425 585
R449 B.n427 B.n426 585
R450 B.n863 B.n862 585
R451 B.n862 B.n861 585
R452 B.n864 B.n424 585
R453 B.n424 B.n423 585
R454 B.n866 B.n865 585
R455 B.n867 B.n866 585
R456 B.n418 B.n417 585
R457 B.n419 B.n418 585
R458 B.n875 B.n874 585
R459 B.n874 B.n873 585
R460 B.n876 B.n416 585
R461 B.n416 B.n415 585
R462 B.n878 B.n877 585
R463 B.n879 B.n878 585
R464 B.n410 B.n409 585
R465 B.n411 B.n410 585
R466 B.n888 B.n887 585
R467 B.n887 B.n886 585
R468 B.n889 B.n408 585
R469 B.n885 B.n408 585
R470 B.n891 B.n890 585
R471 B.n892 B.n891 585
R472 B.n403 B.n402 585
R473 B.n404 B.n403 585
R474 B.n901 B.n900 585
R475 B.n900 B.n899 585
R476 B.n902 B.n401 585
R477 B.n401 B.n400 585
R478 B.n904 B.n903 585
R479 B.n905 B.n904 585
R480 B.n2 B.n0 585
R481 B.n4 B.n2 585
R482 B.n3 B.n1 585
R483 B.n1029 B.n3 585
R484 B.n1027 B.n1026 585
R485 B.n1028 B.n1027 585
R486 B.n1025 B.n9 585
R487 B.n9 B.n8 585
R488 B.n1024 B.n1023 585
R489 B.n1023 B.n1022 585
R490 B.n11 B.n10 585
R491 B.n1021 B.n11 585
R492 B.n1019 B.n1018 585
R493 B.n1020 B.n1019 585
R494 B.n1017 B.n15 585
R495 B.n18 B.n15 585
R496 B.n1016 B.n1015 585
R497 B.n1015 B.n1014 585
R498 B.n17 B.n16 585
R499 B.n1013 B.n17 585
R500 B.n1011 B.n1010 585
R501 B.n1012 B.n1011 585
R502 B.n1009 B.n23 585
R503 B.n23 B.n22 585
R504 B.n1008 B.n1007 585
R505 B.n1007 B.n1006 585
R506 B.n25 B.n24 585
R507 B.n1005 B.n25 585
R508 B.n1003 B.n1002 585
R509 B.n1004 B.n1003 585
R510 B.n1001 B.n30 585
R511 B.n30 B.n29 585
R512 B.n1000 B.n999 585
R513 B.n999 B.n998 585
R514 B.n32 B.n31 585
R515 B.n997 B.n32 585
R516 B.n995 B.n994 585
R517 B.n996 B.n995 585
R518 B.n993 B.n37 585
R519 B.n37 B.n36 585
R520 B.n992 B.n991 585
R521 B.n991 B.n990 585
R522 B.n39 B.n38 585
R523 B.n989 B.n39 585
R524 B.n987 B.n986 585
R525 B.n988 B.n987 585
R526 B.n985 B.n44 585
R527 B.n44 B.n43 585
R528 B.n984 B.n983 585
R529 B.n983 B.n982 585
R530 B.n46 B.n45 585
R531 B.n981 B.n46 585
R532 B.n979 B.n978 585
R533 B.n980 B.n979 585
R534 B.n977 B.n51 585
R535 B.n51 B.n50 585
R536 B.n976 B.n975 585
R537 B.n975 B.n974 585
R538 B.n53 B.n52 585
R539 B.n973 B.n53 585
R540 B.n971 B.n970 585
R541 B.n972 B.n971 585
R542 B.n969 B.n58 585
R543 B.n58 B.n57 585
R544 B.n968 B.n967 585
R545 B.n967 B.n966 585
R546 B.n60 B.n59 585
R547 B.n965 B.n60 585
R548 B.n963 B.n962 585
R549 B.n964 B.n963 585
R550 B.n961 B.n65 585
R551 B.n65 B.n64 585
R552 B.n960 B.n959 585
R553 B.n959 B.n958 585
R554 B.n1032 B.n1031 585
R555 B.n1031 B.n1030 585
R556 B.n802 B.n466 497.305
R557 B.n959 B.n67 497.305
R558 B.n800 B.n468 497.305
R559 B.n956 B.n68 497.305
R560 B.n499 B.t8 364.243
R561 B.n505 B.t12 364.243
R562 B.n138 B.t4 364.243
R563 B.n135 B.t15 364.243
R564 B.n957 B.n133 256.663
R565 B.n957 B.n132 256.663
R566 B.n957 B.n131 256.663
R567 B.n957 B.n130 256.663
R568 B.n957 B.n129 256.663
R569 B.n957 B.n128 256.663
R570 B.n957 B.n127 256.663
R571 B.n957 B.n126 256.663
R572 B.n957 B.n125 256.663
R573 B.n957 B.n124 256.663
R574 B.n957 B.n123 256.663
R575 B.n957 B.n122 256.663
R576 B.n957 B.n121 256.663
R577 B.n957 B.n120 256.663
R578 B.n957 B.n119 256.663
R579 B.n957 B.n118 256.663
R580 B.n957 B.n117 256.663
R581 B.n957 B.n116 256.663
R582 B.n957 B.n115 256.663
R583 B.n957 B.n114 256.663
R584 B.n957 B.n113 256.663
R585 B.n957 B.n112 256.663
R586 B.n957 B.n111 256.663
R587 B.n957 B.n110 256.663
R588 B.n957 B.n109 256.663
R589 B.n957 B.n108 256.663
R590 B.n957 B.n107 256.663
R591 B.n957 B.n106 256.663
R592 B.n957 B.n105 256.663
R593 B.n957 B.n104 256.663
R594 B.n957 B.n103 256.663
R595 B.n957 B.n102 256.663
R596 B.n957 B.n101 256.663
R597 B.n957 B.n100 256.663
R598 B.n957 B.n99 256.663
R599 B.n957 B.n98 256.663
R600 B.n957 B.n97 256.663
R601 B.n957 B.n96 256.663
R602 B.n957 B.n95 256.663
R603 B.n957 B.n94 256.663
R604 B.n957 B.n93 256.663
R605 B.n957 B.n92 256.663
R606 B.n957 B.n91 256.663
R607 B.n957 B.n90 256.663
R608 B.n957 B.n89 256.663
R609 B.n957 B.n88 256.663
R610 B.n957 B.n87 256.663
R611 B.n957 B.n86 256.663
R612 B.n957 B.n85 256.663
R613 B.n957 B.n84 256.663
R614 B.n957 B.n83 256.663
R615 B.n957 B.n82 256.663
R616 B.n957 B.n81 256.663
R617 B.n957 B.n80 256.663
R618 B.n957 B.n79 256.663
R619 B.n957 B.n78 256.663
R620 B.n957 B.n77 256.663
R621 B.n957 B.n76 256.663
R622 B.n957 B.n75 256.663
R623 B.n957 B.n74 256.663
R624 B.n957 B.n73 256.663
R625 B.n957 B.n72 256.663
R626 B.n957 B.n71 256.663
R627 B.n957 B.n70 256.663
R628 B.n957 B.n69 256.663
R629 B.n538 B.n467 256.663
R630 B.n544 B.n467 256.663
R631 B.n546 B.n467 256.663
R632 B.n552 B.n467 256.663
R633 B.n554 B.n467 256.663
R634 B.n560 B.n467 256.663
R635 B.n562 B.n467 256.663
R636 B.n568 B.n467 256.663
R637 B.n570 B.n467 256.663
R638 B.n576 B.n467 256.663
R639 B.n578 B.n467 256.663
R640 B.n584 B.n467 256.663
R641 B.n586 B.n467 256.663
R642 B.n592 B.n467 256.663
R643 B.n594 B.n467 256.663
R644 B.n600 B.n467 256.663
R645 B.n602 B.n467 256.663
R646 B.n608 B.n467 256.663
R647 B.n610 B.n467 256.663
R648 B.n616 B.n467 256.663
R649 B.n618 B.n467 256.663
R650 B.n624 B.n467 256.663
R651 B.n626 B.n467 256.663
R652 B.n632 B.n467 256.663
R653 B.n634 B.n467 256.663
R654 B.n640 B.n467 256.663
R655 B.n642 B.n467 256.663
R656 B.n648 B.n467 256.663
R657 B.n650 B.n467 256.663
R658 B.n656 B.n467 256.663
R659 B.n658 B.n467 256.663
R660 B.n664 B.n467 256.663
R661 B.n666 B.n467 256.663
R662 B.n672 B.n467 256.663
R663 B.n674 B.n467 256.663
R664 B.n681 B.n467 256.663
R665 B.n683 B.n467 256.663
R666 B.n689 B.n467 256.663
R667 B.n691 B.n467 256.663
R668 B.n697 B.n467 256.663
R669 B.n699 B.n467 256.663
R670 B.n705 B.n467 256.663
R671 B.n707 B.n467 256.663
R672 B.n713 B.n467 256.663
R673 B.n715 B.n467 256.663
R674 B.n721 B.n467 256.663
R675 B.n723 B.n467 256.663
R676 B.n729 B.n467 256.663
R677 B.n731 B.n467 256.663
R678 B.n737 B.n467 256.663
R679 B.n739 B.n467 256.663
R680 B.n745 B.n467 256.663
R681 B.n747 B.n467 256.663
R682 B.n753 B.n467 256.663
R683 B.n755 B.n467 256.663
R684 B.n761 B.n467 256.663
R685 B.n763 B.n467 256.663
R686 B.n769 B.n467 256.663
R687 B.n771 B.n467 256.663
R688 B.n777 B.n467 256.663
R689 B.n779 B.n467 256.663
R690 B.n785 B.n467 256.663
R691 B.n787 B.n467 256.663
R692 B.n793 B.n467 256.663
R693 B.n795 B.n467 256.663
R694 B.n802 B.n464 163.367
R695 B.n806 B.n464 163.367
R696 B.n806 B.n458 163.367
R697 B.n814 B.n458 163.367
R698 B.n814 B.n456 163.367
R699 B.n818 B.n456 163.367
R700 B.n818 B.n450 163.367
R701 B.n826 B.n450 163.367
R702 B.n826 B.n448 163.367
R703 B.n830 B.n448 163.367
R704 B.n830 B.n442 163.367
R705 B.n838 B.n442 163.367
R706 B.n838 B.n440 163.367
R707 B.n842 B.n440 163.367
R708 B.n842 B.n434 163.367
R709 B.n850 B.n434 163.367
R710 B.n850 B.n432 163.367
R711 B.n854 B.n432 163.367
R712 B.n854 B.n426 163.367
R713 B.n862 B.n426 163.367
R714 B.n862 B.n424 163.367
R715 B.n866 B.n424 163.367
R716 B.n866 B.n418 163.367
R717 B.n874 B.n418 163.367
R718 B.n874 B.n416 163.367
R719 B.n878 B.n416 163.367
R720 B.n878 B.n410 163.367
R721 B.n887 B.n410 163.367
R722 B.n887 B.n408 163.367
R723 B.n891 B.n408 163.367
R724 B.n891 B.n403 163.367
R725 B.n900 B.n403 163.367
R726 B.n900 B.n401 163.367
R727 B.n904 B.n401 163.367
R728 B.n904 B.n2 163.367
R729 B.n1031 B.n2 163.367
R730 B.n1031 B.n3 163.367
R731 B.n1027 B.n3 163.367
R732 B.n1027 B.n9 163.367
R733 B.n1023 B.n9 163.367
R734 B.n1023 B.n11 163.367
R735 B.n1019 B.n11 163.367
R736 B.n1019 B.n15 163.367
R737 B.n1015 B.n15 163.367
R738 B.n1015 B.n17 163.367
R739 B.n1011 B.n17 163.367
R740 B.n1011 B.n23 163.367
R741 B.n1007 B.n23 163.367
R742 B.n1007 B.n25 163.367
R743 B.n1003 B.n25 163.367
R744 B.n1003 B.n30 163.367
R745 B.n999 B.n30 163.367
R746 B.n999 B.n32 163.367
R747 B.n995 B.n32 163.367
R748 B.n995 B.n37 163.367
R749 B.n991 B.n37 163.367
R750 B.n991 B.n39 163.367
R751 B.n987 B.n39 163.367
R752 B.n987 B.n44 163.367
R753 B.n983 B.n44 163.367
R754 B.n983 B.n46 163.367
R755 B.n979 B.n46 163.367
R756 B.n979 B.n51 163.367
R757 B.n975 B.n51 163.367
R758 B.n975 B.n53 163.367
R759 B.n971 B.n53 163.367
R760 B.n971 B.n58 163.367
R761 B.n967 B.n58 163.367
R762 B.n967 B.n60 163.367
R763 B.n963 B.n60 163.367
R764 B.n963 B.n65 163.367
R765 B.n959 B.n65 163.367
R766 B.n539 B.n537 163.367
R767 B.n543 B.n537 163.367
R768 B.n547 B.n545 163.367
R769 B.n551 B.n535 163.367
R770 B.n555 B.n553 163.367
R771 B.n559 B.n533 163.367
R772 B.n563 B.n561 163.367
R773 B.n567 B.n531 163.367
R774 B.n571 B.n569 163.367
R775 B.n575 B.n529 163.367
R776 B.n579 B.n577 163.367
R777 B.n583 B.n527 163.367
R778 B.n587 B.n585 163.367
R779 B.n591 B.n525 163.367
R780 B.n595 B.n593 163.367
R781 B.n599 B.n523 163.367
R782 B.n603 B.n601 163.367
R783 B.n607 B.n521 163.367
R784 B.n611 B.n609 163.367
R785 B.n615 B.n519 163.367
R786 B.n619 B.n617 163.367
R787 B.n623 B.n517 163.367
R788 B.n627 B.n625 163.367
R789 B.n631 B.n515 163.367
R790 B.n635 B.n633 163.367
R791 B.n639 B.n513 163.367
R792 B.n643 B.n641 163.367
R793 B.n647 B.n511 163.367
R794 B.n651 B.n649 163.367
R795 B.n655 B.n509 163.367
R796 B.n659 B.n657 163.367
R797 B.n663 B.n504 163.367
R798 B.n667 B.n665 163.367
R799 B.n671 B.n502 163.367
R800 B.n675 B.n673 163.367
R801 B.n680 B.n498 163.367
R802 B.n684 B.n682 163.367
R803 B.n688 B.n496 163.367
R804 B.n692 B.n690 163.367
R805 B.n696 B.n494 163.367
R806 B.n700 B.n698 163.367
R807 B.n704 B.n492 163.367
R808 B.n708 B.n706 163.367
R809 B.n712 B.n490 163.367
R810 B.n716 B.n714 163.367
R811 B.n720 B.n488 163.367
R812 B.n724 B.n722 163.367
R813 B.n728 B.n486 163.367
R814 B.n732 B.n730 163.367
R815 B.n736 B.n484 163.367
R816 B.n740 B.n738 163.367
R817 B.n744 B.n482 163.367
R818 B.n748 B.n746 163.367
R819 B.n752 B.n480 163.367
R820 B.n756 B.n754 163.367
R821 B.n760 B.n478 163.367
R822 B.n764 B.n762 163.367
R823 B.n768 B.n476 163.367
R824 B.n772 B.n770 163.367
R825 B.n776 B.n474 163.367
R826 B.n780 B.n778 163.367
R827 B.n784 B.n472 163.367
R828 B.n788 B.n786 163.367
R829 B.n792 B.n470 163.367
R830 B.n796 B.n794 163.367
R831 B.n800 B.n462 163.367
R832 B.n808 B.n462 163.367
R833 B.n808 B.n460 163.367
R834 B.n812 B.n460 163.367
R835 B.n812 B.n453 163.367
R836 B.n820 B.n453 163.367
R837 B.n820 B.n451 163.367
R838 B.n824 B.n451 163.367
R839 B.n824 B.n446 163.367
R840 B.n832 B.n446 163.367
R841 B.n832 B.n444 163.367
R842 B.n836 B.n444 163.367
R843 B.n836 B.n438 163.367
R844 B.n844 B.n438 163.367
R845 B.n844 B.n436 163.367
R846 B.n848 B.n436 163.367
R847 B.n848 B.n430 163.367
R848 B.n856 B.n430 163.367
R849 B.n856 B.n428 163.367
R850 B.n860 B.n428 163.367
R851 B.n860 B.n422 163.367
R852 B.n868 B.n422 163.367
R853 B.n868 B.n420 163.367
R854 B.n872 B.n420 163.367
R855 B.n872 B.n414 163.367
R856 B.n880 B.n414 163.367
R857 B.n880 B.n412 163.367
R858 B.n884 B.n412 163.367
R859 B.n884 B.n407 163.367
R860 B.n893 B.n407 163.367
R861 B.n893 B.n405 163.367
R862 B.n898 B.n405 163.367
R863 B.n898 B.n399 163.367
R864 B.n906 B.n399 163.367
R865 B.n907 B.n906 163.367
R866 B.n907 B.n5 163.367
R867 B.n6 B.n5 163.367
R868 B.n7 B.n6 163.367
R869 B.n912 B.n7 163.367
R870 B.n912 B.n12 163.367
R871 B.n13 B.n12 163.367
R872 B.n14 B.n13 163.367
R873 B.n917 B.n14 163.367
R874 B.n917 B.n19 163.367
R875 B.n20 B.n19 163.367
R876 B.n21 B.n20 163.367
R877 B.n922 B.n21 163.367
R878 B.n922 B.n26 163.367
R879 B.n27 B.n26 163.367
R880 B.n28 B.n27 163.367
R881 B.n927 B.n28 163.367
R882 B.n927 B.n33 163.367
R883 B.n34 B.n33 163.367
R884 B.n35 B.n34 163.367
R885 B.n932 B.n35 163.367
R886 B.n932 B.n40 163.367
R887 B.n41 B.n40 163.367
R888 B.n42 B.n41 163.367
R889 B.n937 B.n42 163.367
R890 B.n937 B.n47 163.367
R891 B.n48 B.n47 163.367
R892 B.n49 B.n48 163.367
R893 B.n942 B.n49 163.367
R894 B.n942 B.n54 163.367
R895 B.n55 B.n54 163.367
R896 B.n56 B.n55 163.367
R897 B.n947 B.n56 163.367
R898 B.n947 B.n61 163.367
R899 B.n62 B.n61 163.367
R900 B.n63 B.n62 163.367
R901 B.n952 B.n63 163.367
R902 B.n952 B.n68 163.367
R903 B.n142 B.n141 163.367
R904 B.n146 B.n145 163.367
R905 B.n150 B.n149 163.367
R906 B.n154 B.n153 163.367
R907 B.n158 B.n157 163.367
R908 B.n162 B.n161 163.367
R909 B.n166 B.n165 163.367
R910 B.n170 B.n169 163.367
R911 B.n174 B.n173 163.367
R912 B.n178 B.n177 163.367
R913 B.n182 B.n181 163.367
R914 B.n186 B.n185 163.367
R915 B.n190 B.n189 163.367
R916 B.n194 B.n193 163.367
R917 B.n198 B.n197 163.367
R918 B.n202 B.n201 163.367
R919 B.n206 B.n205 163.367
R920 B.n210 B.n209 163.367
R921 B.n214 B.n213 163.367
R922 B.n218 B.n217 163.367
R923 B.n222 B.n221 163.367
R924 B.n226 B.n225 163.367
R925 B.n230 B.n229 163.367
R926 B.n234 B.n233 163.367
R927 B.n238 B.n237 163.367
R928 B.n242 B.n241 163.367
R929 B.n246 B.n245 163.367
R930 B.n250 B.n249 163.367
R931 B.n254 B.n253 163.367
R932 B.n258 B.n257 163.367
R933 B.n263 B.n262 163.367
R934 B.n267 B.n266 163.367
R935 B.n271 B.n270 163.367
R936 B.n275 B.n274 163.367
R937 B.n279 B.n278 163.367
R938 B.n283 B.n282 163.367
R939 B.n287 B.n286 163.367
R940 B.n291 B.n290 163.367
R941 B.n295 B.n294 163.367
R942 B.n299 B.n298 163.367
R943 B.n303 B.n302 163.367
R944 B.n307 B.n306 163.367
R945 B.n311 B.n310 163.367
R946 B.n315 B.n314 163.367
R947 B.n319 B.n318 163.367
R948 B.n323 B.n322 163.367
R949 B.n327 B.n326 163.367
R950 B.n331 B.n330 163.367
R951 B.n335 B.n334 163.367
R952 B.n339 B.n338 163.367
R953 B.n343 B.n342 163.367
R954 B.n347 B.n346 163.367
R955 B.n351 B.n350 163.367
R956 B.n355 B.n354 163.367
R957 B.n359 B.n358 163.367
R958 B.n363 B.n362 163.367
R959 B.n367 B.n366 163.367
R960 B.n371 B.n370 163.367
R961 B.n375 B.n374 163.367
R962 B.n379 B.n378 163.367
R963 B.n383 B.n382 163.367
R964 B.n387 B.n386 163.367
R965 B.n391 B.n390 163.367
R966 B.n395 B.n394 163.367
R967 B.n956 B.n134 163.367
R968 B.n499 B.t11 130.255
R969 B.n135 B.t16 130.255
R970 B.n505 B.t14 130.23
R971 B.n138 B.t6 130.23
R972 B.n538 B.n466 71.676
R973 B.n544 B.n543 71.676
R974 B.n547 B.n546 71.676
R975 B.n552 B.n551 71.676
R976 B.n555 B.n554 71.676
R977 B.n560 B.n559 71.676
R978 B.n563 B.n562 71.676
R979 B.n568 B.n567 71.676
R980 B.n571 B.n570 71.676
R981 B.n576 B.n575 71.676
R982 B.n579 B.n578 71.676
R983 B.n584 B.n583 71.676
R984 B.n587 B.n586 71.676
R985 B.n592 B.n591 71.676
R986 B.n595 B.n594 71.676
R987 B.n600 B.n599 71.676
R988 B.n603 B.n602 71.676
R989 B.n608 B.n607 71.676
R990 B.n611 B.n610 71.676
R991 B.n616 B.n615 71.676
R992 B.n619 B.n618 71.676
R993 B.n624 B.n623 71.676
R994 B.n627 B.n626 71.676
R995 B.n632 B.n631 71.676
R996 B.n635 B.n634 71.676
R997 B.n640 B.n639 71.676
R998 B.n643 B.n642 71.676
R999 B.n648 B.n647 71.676
R1000 B.n651 B.n650 71.676
R1001 B.n656 B.n655 71.676
R1002 B.n659 B.n658 71.676
R1003 B.n664 B.n663 71.676
R1004 B.n667 B.n666 71.676
R1005 B.n672 B.n671 71.676
R1006 B.n675 B.n674 71.676
R1007 B.n681 B.n680 71.676
R1008 B.n684 B.n683 71.676
R1009 B.n689 B.n688 71.676
R1010 B.n692 B.n691 71.676
R1011 B.n697 B.n696 71.676
R1012 B.n700 B.n699 71.676
R1013 B.n705 B.n704 71.676
R1014 B.n708 B.n707 71.676
R1015 B.n713 B.n712 71.676
R1016 B.n716 B.n715 71.676
R1017 B.n721 B.n720 71.676
R1018 B.n724 B.n723 71.676
R1019 B.n729 B.n728 71.676
R1020 B.n732 B.n731 71.676
R1021 B.n737 B.n736 71.676
R1022 B.n740 B.n739 71.676
R1023 B.n745 B.n744 71.676
R1024 B.n748 B.n747 71.676
R1025 B.n753 B.n752 71.676
R1026 B.n756 B.n755 71.676
R1027 B.n761 B.n760 71.676
R1028 B.n764 B.n763 71.676
R1029 B.n769 B.n768 71.676
R1030 B.n772 B.n771 71.676
R1031 B.n777 B.n776 71.676
R1032 B.n780 B.n779 71.676
R1033 B.n785 B.n784 71.676
R1034 B.n788 B.n787 71.676
R1035 B.n793 B.n792 71.676
R1036 B.n796 B.n795 71.676
R1037 B.n69 B.n67 71.676
R1038 B.n142 B.n70 71.676
R1039 B.n146 B.n71 71.676
R1040 B.n150 B.n72 71.676
R1041 B.n154 B.n73 71.676
R1042 B.n158 B.n74 71.676
R1043 B.n162 B.n75 71.676
R1044 B.n166 B.n76 71.676
R1045 B.n170 B.n77 71.676
R1046 B.n174 B.n78 71.676
R1047 B.n178 B.n79 71.676
R1048 B.n182 B.n80 71.676
R1049 B.n186 B.n81 71.676
R1050 B.n190 B.n82 71.676
R1051 B.n194 B.n83 71.676
R1052 B.n198 B.n84 71.676
R1053 B.n202 B.n85 71.676
R1054 B.n206 B.n86 71.676
R1055 B.n210 B.n87 71.676
R1056 B.n214 B.n88 71.676
R1057 B.n218 B.n89 71.676
R1058 B.n222 B.n90 71.676
R1059 B.n226 B.n91 71.676
R1060 B.n230 B.n92 71.676
R1061 B.n234 B.n93 71.676
R1062 B.n238 B.n94 71.676
R1063 B.n242 B.n95 71.676
R1064 B.n246 B.n96 71.676
R1065 B.n250 B.n97 71.676
R1066 B.n254 B.n98 71.676
R1067 B.n258 B.n99 71.676
R1068 B.n263 B.n100 71.676
R1069 B.n267 B.n101 71.676
R1070 B.n271 B.n102 71.676
R1071 B.n275 B.n103 71.676
R1072 B.n279 B.n104 71.676
R1073 B.n283 B.n105 71.676
R1074 B.n287 B.n106 71.676
R1075 B.n291 B.n107 71.676
R1076 B.n295 B.n108 71.676
R1077 B.n299 B.n109 71.676
R1078 B.n303 B.n110 71.676
R1079 B.n307 B.n111 71.676
R1080 B.n311 B.n112 71.676
R1081 B.n315 B.n113 71.676
R1082 B.n319 B.n114 71.676
R1083 B.n323 B.n115 71.676
R1084 B.n327 B.n116 71.676
R1085 B.n331 B.n117 71.676
R1086 B.n335 B.n118 71.676
R1087 B.n339 B.n119 71.676
R1088 B.n343 B.n120 71.676
R1089 B.n347 B.n121 71.676
R1090 B.n351 B.n122 71.676
R1091 B.n355 B.n123 71.676
R1092 B.n359 B.n124 71.676
R1093 B.n363 B.n125 71.676
R1094 B.n367 B.n126 71.676
R1095 B.n371 B.n127 71.676
R1096 B.n375 B.n128 71.676
R1097 B.n379 B.n129 71.676
R1098 B.n383 B.n130 71.676
R1099 B.n387 B.n131 71.676
R1100 B.n391 B.n132 71.676
R1101 B.n395 B.n133 71.676
R1102 B.n134 B.n133 71.676
R1103 B.n394 B.n132 71.676
R1104 B.n390 B.n131 71.676
R1105 B.n386 B.n130 71.676
R1106 B.n382 B.n129 71.676
R1107 B.n378 B.n128 71.676
R1108 B.n374 B.n127 71.676
R1109 B.n370 B.n126 71.676
R1110 B.n366 B.n125 71.676
R1111 B.n362 B.n124 71.676
R1112 B.n358 B.n123 71.676
R1113 B.n354 B.n122 71.676
R1114 B.n350 B.n121 71.676
R1115 B.n346 B.n120 71.676
R1116 B.n342 B.n119 71.676
R1117 B.n338 B.n118 71.676
R1118 B.n334 B.n117 71.676
R1119 B.n330 B.n116 71.676
R1120 B.n326 B.n115 71.676
R1121 B.n322 B.n114 71.676
R1122 B.n318 B.n113 71.676
R1123 B.n314 B.n112 71.676
R1124 B.n310 B.n111 71.676
R1125 B.n306 B.n110 71.676
R1126 B.n302 B.n109 71.676
R1127 B.n298 B.n108 71.676
R1128 B.n294 B.n107 71.676
R1129 B.n290 B.n106 71.676
R1130 B.n286 B.n105 71.676
R1131 B.n282 B.n104 71.676
R1132 B.n278 B.n103 71.676
R1133 B.n274 B.n102 71.676
R1134 B.n270 B.n101 71.676
R1135 B.n266 B.n100 71.676
R1136 B.n262 B.n99 71.676
R1137 B.n257 B.n98 71.676
R1138 B.n253 B.n97 71.676
R1139 B.n249 B.n96 71.676
R1140 B.n245 B.n95 71.676
R1141 B.n241 B.n94 71.676
R1142 B.n237 B.n93 71.676
R1143 B.n233 B.n92 71.676
R1144 B.n229 B.n91 71.676
R1145 B.n225 B.n90 71.676
R1146 B.n221 B.n89 71.676
R1147 B.n217 B.n88 71.676
R1148 B.n213 B.n87 71.676
R1149 B.n209 B.n86 71.676
R1150 B.n205 B.n85 71.676
R1151 B.n201 B.n84 71.676
R1152 B.n197 B.n83 71.676
R1153 B.n193 B.n82 71.676
R1154 B.n189 B.n81 71.676
R1155 B.n185 B.n80 71.676
R1156 B.n181 B.n79 71.676
R1157 B.n177 B.n78 71.676
R1158 B.n173 B.n77 71.676
R1159 B.n169 B.n76 71.676
R1160 B.n165 B.n75 71.676
R1161 B.n161 B.n74 71.676
R1162 B.n157 B.n73 71.676
R1163 B.n153 B.n72 71.676
R1164 B.n149 B.n71 71.676
R1165 B.n145 B.n70 71.676
R1166 B.n141 B.n69 71.676
R1167 B.n539 B.n538 71.676
R1168 B.n545 B.n544 71.676
R1169 B.n546 B.n535 71.676
R1170 B.n553 B.n552 71.676
R1171 B.n554 B.n533 71.676
R1172 B.n561 B.n560 71.676
R1173 B.n562 B.n531 71.676
R1174 B.n569 B.n568 71.676
R1175 B.n570 B.n529 71.676
R1176 B.n577 B.n576 71.676
R1177 B.n578 B.n527 71.676
R1178 B.n585 B.n584 71.676
R1179 B.n586 B.n525 71.676
R1180 B.n593 B.n592 71.676
R1181 B.n594 B.n523 71.676
R1182 B.n601 B.n600 71.676
R1183 B.n602 B.n521 71.676
R1184 B.n609 B.n608 71.676
R1185 B.n610 B.n519 71.676
R1186 B.n617 B.n616 71.676
R1187 B.n618 B.n517 71.676
R1188 B.n625 B.n624 71.676
R1189 B.n626 B.n515 71.676
R1190 B.n633 B.n632 71.676
R1191 B.n634 B.n513 71.676
R1192 B.n641 B.n640 71.676
R1193 B.n642 B.n511 71.676
R1194 B.n649 B.n648 71.676
R1195 B.n650 B.n509 71.676
R1196 B.n657 B.n656 71.676
R1197 B.n658 B.n504 71.676
R1198 B.n665 B.n664 71.676
R1199 B.n666 B.n502 71.676
R1200 B.n673 B.n672 71.676
R1201 B.n674 B.n498 71.676
R1202 B.n682 B.n681 71.676
R1203 B.n683 B.n496 71.676
R1204 B.n690 B.n689 71.676
R1205 B.n691 B.n494 71.676
R1206 B.n698 B.n697 71.676
R1207 B.n699 B.n492 71.676
R1208 B.n706 B.n705 71.676
R1209 B.n707 B.n490 71.676
R1210 B.n714 B.n713 71.676
R1211 B.n715 B.n488 71.676
R1212 B.n722 B.n721 71.676
R1213 B.n723 B.n486 71.676
R1214 B.n730 B.n729 71.676
R1215 B.n731 B.n484 71.676
R1216 B.n738 B.n737 71.676
R1217 B.n739 B.n482 71.676
R1218 B.n746 B.n745 71.676
R1219 B.n747 B.n480 71.676
R1220 B.n754 B.n753 71.676
R1221 B.n755 B.n478 71.676
R1222 B.n762 B.n761 71.676
R1223 B.n763 B.n476 71.676
R1224 B.n770 B.n769 71.676
R1225 B.n771 B.n474 71.676
R1226 B.n778 B.n777 71.676
R1227 B.n779 B.n472 71.676
R1228 B.n786 B.n785 71.676
R1229 B.n787 B.n470 71.676
R1230 B.n794 B.n793 71.676
R1231 B.n795 B.n468 71.676
R1232 B.n500 B.t10 68.5813
R1233 B.n136 B.t17 68.5813
R1234 B.n506 B.t13 68.5566
R1235 B.n139 B.t7 68.5566
R1236 B.n801 B.n467 62.6455
R1237 B.n958 B.n957 62.6455
R1238 B.n500 B.n499 61.6732
R1239 B.n506 B.n505 61.6732
R1240 B.n139 B.n138 61.6732
R1241 B.n136 B.n135 61.6732
R1242 B.n677 B.n500 59.5399
R1243 B.n507 B.n506 59.5399
R1244 B.n260 B.n139 59.5399
R1245 B.n137 B.n136 59.5399
R1246 B.n960 B.n66 32.3127
R1247 B.n955 B.n954 32.3127
R1248 B.n799 B.n798 32.3127
R1249 B.n803 B.n465 32.3127
R1250 B.n801 B.n463 31.555
R1251 B.n807 B.n463 31.555
R1252 B.n807 B.n459 31.555
R1253 B.n813 B.n459 31.555
R1254 B.n813 B.n454 31.555
R1255 B.n819 B.n454 31.555
R1256 B.n819 B.n455 31.555
R1257 B.n825 B.n447 31.555
R1258 B.n831 B.n447 31.555
R1259 B.n831 B.n443 31.555
R1260 B.n837 B.n443 31.555
R1261 B.n837 B.n439 31.555
R1262 B.n843 B.n439 31.555
R1263 B.n843 B.n435 31.555
R1264 B.n849 B.n435 31.555
R1265 B.n849 B.n431 31.555
R1266 B.n855 B.n431 31.555
R1267 B.n855 B.n427 31.555
R1268 B.n861 B.n427 31.555
R1269 B.n867 B.n423 31.555
R1270 B.n867 B.n419 31.555
R1271 B.n873 B.n419 31.555
R1272 B.n873 B.n415 31.555
R1273 B.n879 B.n415 31.555
R1274 B.n879 B.n411 31.555
R1275 B.n886 B.n411 31.555
R1276 B.n886 B.n885 31.555
R1277 B.n892 B.n404 31.555
R1278 B.n899 B.n404 31.555
R1279 B.n899 B.n400 31.555
R1280 B.n905 B.n400 31.555
R1281 B.n905 B.n4 31.555
R1282 B.n1030 B.n4 31.555
R1283 B.n1030 B.n1029 31.555
R1284 B.n1029 B.n1028 31.555
R1285 B.n1028 B.n8 31.555
R1286 B.n1022 B.n8 31.555
R1287 B.n1022 B.n1021 31.555
R1288 B.n1021 B.n1020 31.555
R1289 B.n1014 B.n18 31.555
R1290 B.n1014 B.n1013 31.555
R1291 B.n1013 B.n1012 31.555
R1292 B.n1012 B.n22 31.555
R1293 B.n1006 B.n22 31.555
R1294 B.n1006 B.n1005 31.555
R1295 B.n1005 B.n1004 31.555
R1296 B.n1004 B.n29 31.555
R1297 B.n998 B.n997 31.555
R1298 B.n997 B.n996 31.555
R1299 B.n996 B.n36 31.555
R1300 B.n990 B.n36 31.555
R1301 B.n990 B.n989 31.555
R1302 B.n989 B.n988 31.555
R1303 B.n988 B.n43 31.555
R1304 B.n982 B.n43 31.555
R1305 B.n982 B.n981 31.555
R1306 B.n981 B.n980 31.555
R1307 B.n980 B.n50 31.555
R1308 B.n974 B.n50 31.555
R1309 B.n973 B.n972 31.555
R1310 B.n972 B.n57 31.555
R1311 B.n966 B.n57 31.555
R1312 B.n966 B.n965 31.555
R1313 B.n965 B.n964 31.555
R1314 B.n964 B.n64 31.555
R1315 B.n958 B.n64 31.555
R1316 B.n455 B.t9 25.5225
R1317 B.t5 B.n973 25.5225
R1318 B.n885 B.t2 22.7383
R1319 B.n18 B.t1 22.7383
R1320 B.t3 B.n423 19.9541
R1321 B.t0 B.n29 19.9541
R1322 B B.n1032 18.0485
R1323 B.n861 B.t3 11.6014
R1324 B.n998 B.t0 11.6014
R1325 B.n140 B.n66 10.6151
R1326 B.n143 B.n140 10.6151
R1327 B.n144 B.n143 10.6151
R1328 B.n147 B.n144 10.6151
R1329 B.n148 B.n147 10.6151
R1330 B.n151 B.n148 10.6151
R1331 B.n152 B.n151 10.6151
R1332 B.n155 B.n152 10.6151
R1333 B.n156 B.n155 10.6151
R1334 B.n159 B.n156 10.6151
R1335 B.n160 B.n159 10.6151
R1336 B.n163 B.n160 10.6151
R1337 B.n164 B.n163 10.6151
R1338 B.n167 B.n164 10.6151
R1339 B.n168 B.n167 10.6151
R1340 B.n171 B.n168 10.6151
R1341 B.n172 B.n171 10.6151
R1342 B.n175 B.n172 10.6151
R1343 B.n176 B.n175 10.6151
R1344 B.n179 B.n176 10.6151
R1345 B.n180 B.n179 10.6151
R1346 B.n183 B.n180 10.6151
R1347 B.n184 B.n183 10.6151
R1348 B.n187 B.n184 10.6151
R1349 B.n188 B.n187 10.6151
R1350 B.n191 B.n188 10.6151
R1351 B.n192 B.n191 10.6151
R1352 B.n195 B.n192 10.6151
R1353 B.n196 B.n195 10.6151
R1354 B.n199 B.n196 10.6151
R1355 B.n200 B.n199 10.6151
R1356 B.n203 B.n200 10.6151
R1357 B.n204 B.n203 10.6151
R1358 B.n207 B.n204 10.6151
R1359 B.n208 B.n207 10.6151
R1360 B.n211 B.n208 10.6151
R1361 B.n212 B.n211 10.6151
R1362 B.n215 B.n212 10.6151
R1363 B.n216 B.n215 10.6151
R1364 B.n219 B.n216 10.6151
R1365 B.n220 B.n219 10.6151
R1366 B.n223 B.n220 10.6151
R1367 B.n224 B.n223 10.6151
R1368 B.n227 B.n224 10.6151
R1369 B.n228 B.n227 10.6151
R1370 B.n231 B.n228 10.6151
R1371 B.n232 B.n231 10.6151
R1372 B.n235 B.n232 10.6151
R1373 B.n236 B.n235 10.6151
R1374 B.n239 B.n236 10.6151
R1375 B.n240 B.n239 10.6151
R1376 B.n243 B.n240 10.6151
R1377 B.n244 B.n243 10.6151
R1378 B.n247 B.n244 10.6151
R1379 B.n248 B.n247 10.6151
R1380 B.n251 B.n248 10.6151
R1381 B.n252 B.n251 10.6151
R1382 B.n255 B.n252 10.6151
R1383 B.n256 B.n255 10.6151
R1384 B.n259 B.n256 10.6151
R1385 B.n264 B.n261 10.6151
R1386 B.n265 B.n264 10.6151
R1387 B.n268 B.n265 10.6151
R1388 B.n269 B.n268 10.6151
R1389 B.n272 B.n269 10.6151
R1390 B.n273 B.n272 10.6151
R1391 B.n276 B.n273 10.6151
R1392 B.n277 B.n276 10.6151
R1393 B.n281 B.n280 10.6151
R1394 B.n284 B.n281 10.6151
R1395 B.n285 B.n284 10.6151
R1396 B.n288 B.n285 10.6151
R1397 B.n289 B.n288 10.6151
R1398 B.n292 B.n289 10.6151
R1399 B.n293 B.n292 10.6151
R1400 B.n296 B.n293 10.6151
R1401 B.n297 B.n296 10.6151
R1402 B.n300 B.n297 10.6151
R1403 B.n301 B.n300 10.6151
R1404 B.n304 B.n301 10.6151
R1405 B.n305 B.n304 10.6151
R1406 B.n308 B.n305 10.6151
R1407 B.n309 B.n308 10.6151
R1408 B.n312 B.n309 10.6151
R1409 B.n313 B.n312 10.6151
R1410 B.n316 B.n313 10.6151
R1411 B.n317 B.n316 10.6151
R1412 B.n320 B.n317 10.6151
R1413 B.n321 B.n320 10.6151
R1414 B.n324 B.n321 10.6151
R1415 B.n325 B.n324 10.6151
R1416 B.n328 B.n325 10.6151
R1417 B.n329 B.n328 10.6151
R1418 B.n332 B.n329 10.6151
R1419 B.n333 B.n332 10.6151
R1420 B.n336 B.n333 10.6151
R1421 B.n337 B.n336 10.6151
R1422 B.n340 B.n337 10.6151
R1423 B.n341 B.n340 10.6151
R1424 B.n344 B.n341 10.6151
R1425 B.n345 B.n344 10.6151
R1426 B.n348 B.n345 10.6151
R1427 B.n349 B.n348 10.6151
R1428 B.n352 B.n349 10.6151
R1429 B.n353 B.n352 10.6151
R1430 B.n356 B.n353 10.6151
R1431 B.n357 B.n356 10.6151
R1432 B.n360 B.n357 10.6151
R1433 B.n361 B.n360 10.6151
R1434 B.n364 B.n361 10.6151
R1435 B.n365 B.n364 10.6151
R1436 B.n368 B.n365 10.6151
R1437 B.n369 B.n368 10.6151
R1438 B.n372 B.n369 10.6151
R1439 B.n373 B.n372 10.6151
R1440 B.n376 B.n373 10.6151
R1441 B.n377 B.n376 10.6151
R1442 B.n380 B.n377 10.6151
R1443 B.n381 B.n380 10.6151
R1444 B.n384 B.n381 10.6151
R1445 B.n385 B.n384 10.6151
R1446 B.n388 B.n385 10.6151
R1447 B.n389 B.n388 10.6151
R1448 B.n392 B.n389 10.6151
R1449 B.n393 B.n392 10.6151
R1450 B.n396 B.n393 10.6151
R1451 B.n397 B.n396 10.6151
R1452 B.n955 B.n397 10.6151
R1453 B.n799 B.n461 10.6151
R1454 B.n809 B.n461 10.6151
R1455 B.n810 B.n809 10.6151
R1456 B.n811 B.n810 10.6151
R1457 B.n811 B.n452 10.6151
R1458 B.n821 B.n452 10.6151
R1459 B.n822 B.n821 10.6151
R1460 B.n823 B.n822 10.6151
R1461 B.n823 B.n445 10.6151
R1462 B.n833 B.n445 10.6151
R1463 B.n834 B.n833 10.6151
R1464 B.n835 B.n834 10.6151
R1465 B.n835 B.n437 10.6151
R1466 B.n845 B.n437 10.6151
R1467 B.n846 B.n845 10.6151
R1468 B.n847 B.n846 10.6151
R1469 B.n847 B.n429 10.6151
R1470 B.n857 B.n429 10.6151
R1471 B.n858 B.n857 10.6151
R1472 B.n859 B.n858 10.6151
R1473 B.n859 B.n421 10.6151
R1474 B.n869 B.n421 10.6151
R1475 B.n870 B.n869 10.6151
R1476 B.n871 B.n870 10.6151
R1477 B.n871 B.n413 10.6151
R1478 B.n881 B.n413 10.6151
R1479 B.n882 B.n881 10.6151
R1480 B.n883 B.n882 10.6151
R1481 B.n883 B.n406 10.6151
R1482 B.n894 B.n406 10.6151
R1483 B.n895 B.n894 10.6151
R1484 B.n897 B.n895 10.6151
R1485 B.n897 B.n896 10.6151
R1486 B.n896 B.n398 10.6151
R1487 B.n908 B.n398 10.6151
R1488 B.n909 B.n908 10.6151
R1489 B.n910 B.n909 10.6151
R1490 B.n911 B.n910 10.6151
R1491 B.n913 B.n911 10.6151
R1492 B.n914 B.n913 10.6151
R1493 B.n915 B.n914 10.6151
R1494 B.n916 B.n915 10.6151
R1495 B.n918 B.n916 10.6151
R1496 B.n919 B.n918 10.6151
R1497 B.n920 B.n919 10.6151
R1498 B.n921 B.n920 10.6151
R1499 B.n923 B.n921 10.6151
R1500 B.n924 B.n923 10.6151
R1501 B.n925 B.n924 10.6151
R1502 B.n926 B.n925 10.6151
R1503 B.n928 B.n926 10.6151
R1504 B.n929 B.n928 10.6151
R1505 B.n930 B.n929 10.6151
R1506 B.n931 B.n930 10.6151
R1507 B.n933 B.n931 10.6151
R1508 B.n934 B.n933 10.6151
R1509 B.n935 B.n934 10.6151
R1510 B.n936 B.n935 10.6151
R1511 B.n938 B.n936 10.6151
R1512 B.n939 B.n938 10.6151
R1513 B.n940 B.n939 10.6151
R1514 B.n941 B.n940 10.6151
R1515 B.n943 B.n941 10.6151
R1516 B.n944 B.n943 10.6151
R1517 B.n945 B.n944 10.6151
R1518 B.n946 B.n945 10.6151
R1519 B.n948 B.n946 10.6151
R1520 B.n949 B.n948 10.6151
R1521 B.n950 B.n949 10.6151
R1522 B.n951 B.n950 10.6151
R1523 B.n953 B.n951 10.6151
R1524 B.n954 B.n953 10.6151
R1525 B.n540 B.n465 10.6151
R1526 B.n541 B.n540 10.6151
R1527 B.n542 B.n541 10.6151
R1528 B.n542 B.n536 10.6151
R1529 B.n548 B.n536 10.6151
R1530 B.n549 B.n548 10.6151
R1531 B.n550 B.n549 10.6151
R1532 B.n550 B.n534 10.6151
R1533 B.n556 B.n534 10.6151
R1534 B.n557 B.n556 10.6151
R1535 B.n558 B.n557 10.6151
R1536 B.n558 B.n532 10.6151
R1537 B.n564 B.n532 10.6151
R1538 B.n565 B.n564 10.6151
R1539 B.n566 B.n565 10.6151
R1540 B.n566 B.n530 10.6151
R1541 B.n572 B.n530 10.6151
R1542 B.n573 B.n572 10.6151
R1543 B.n574 B.n573 10.6151
R1544 B.n574 B.n528 10.6151
R1545 B.n580 B.n528 10.6151
R1546 B.n581 B.n580 10.6151
R1547 B.n582 B.n581 10.6151
R1548 B.n582 B.n526 10.6151
R1549 B.n588 B.n526 10.6151
R1550 B.n589 B.n588 10.6151
R1551 B.n590 B.n589 10.6151
R1552 B.n590 B.n524 10.6151
R1553 B.n596 B.n524 10.6151
R1554 B.n597 B.n596 10.6151
R1555 B.n598 B.n597 10.6151
R1556 B.n598 B.n522 10.6151
R1557 B.n604 B.n522 10.6151
R1558 B.n605 B.n604 10.6151
R1559 B.n606 B.n605 10.6151
R1560 B.n606 B.n520 10.6151
R1561 B.n612 B.n520 10.6151
R1562 B.n613 B.n612 10.6151
R1563 B.n614 B.n613 10.6151
R1564 B.n614 B.n518 10.6151
R1565 B.n620 B.n518 10.6151
R1566 B.n621 B.n620 10.6151
R1567 B.n622 B.n621 10.6151
R1568 B.n622 B.n516 10.6151
R1569 B.n628 B.n516 10.6151
R1570 B.n629 B.n628 10.6151
R1571 B.n630 B.n629 10.6151
R1572 B.n630 B.n514 10.6151
R1573 B.n636 B.n514 10.6151
R1574 B.n637 B.n636 10.6151
R1575 B.n638 B.n637 10.6151
R1576 B.n638 B.n512 10.6151
R1577 B.n644 B.n512 10.6151
R1578 B.n645 B.n644 10.6151
R1579 B.n646 B.n645 10.6151
R1580 B.n646 B.n510 10.6151
R1581 B.n652 B.n510 10.6151
R1582 B.n653 B.n652 10.6151
R1583 B.n654 B.n653 10.6151
R1584 B.n654 B.n508 10.6151
R1585 B.n661 B.n660 10.6151
R1586 B.n662 B.n661 10.6151
R1587 B.n662 B.n503 10.6151
R1588 B.n668 B.n503 10.6151
R1589 B.n669 B.n668 10.6151
R1590 B.n670 B.n669 10.6151
R1591 B.n670 B.n501 10.6151
R1592 B.n676 B.n501 10.6151
R1593 B.n679 B.n678 10.6151
R1594 B.n679 B.n497 10.6151
R1595 B.n685 B.n497 10.6151
R1596 B.n686 B.n685 10.6151
R1597 B.n687 B.n686 10.6151
R1598 B.n687 B.n495 10.6151
R1599 B.n693 B.n495 10.6151
R1600 B.n694 B.n693 10.6151
R1601 B.n695 B.n694 10.6151
R1602 B.n695 B.n493 10.6151
R1603 B.n701 B.n493 10.6151
R1604 B.n702 B.n701 10.6151
R1605 B.n703 B.n702 10.6151
R1606 B.n703 B.n491 10.6151
R1607 B.n709 B.n491 10.6151
R1608 B.n710 B.n709 10.6151
R1609 B.n711 B.n710 10.6151
R1610 B.n711 B.n489 10.6151
R1611 B.n717 B.n489 10.6151
R1612 B.n718 B.n717 10.6151
R1613 B.n719 B.n718 10.6151
R1614 B.n719 B.n487 10.6151
R1615 B.n725 B.n487 10.6151
R1616 B.n726 B.n725 10.6151
R1617 B.n727 B.n726 10.6151
R1618 B.n727 B.n485 10.6151
R1619 B.n733 B.n485 10.6151
R1620 B.n734 B.n733 10.6151
R1621 B.n735 B.n734 10.6151
R1622 B.n735 B.n483 10.6151
R1623 B.n741 B.n483 10.6151
R1624 B.n742 B.n741 10.6151
R1625 B.n743 B.n742 10.6151
R1626 B.n743 B.n481 10.6151
R1627 B.n749 B.n481 10.6151
R1628 B.n750 B.n749 10.6151
R1629 B.n751 B.n750 10.6151
R1630 B.n751 B.n479 10.6151
R1631 B.n757 B.n479 10.6151
R1632 B.n758 B.n757 10.6151
R1633 B.n759 B.n758 10.6151
R1634 B.n759 B.n477 10.6151
R1635 B.n765 B.n477 10.6151
R1636 B.n766 B.n765 10.6151
R1637 B.n767 B.n766 10.6151
R1638 B.n767 B.n475 10.6151
R1639 B.n773 B.n475 10.6151
R1640 B.n774 B.n773 10.6151
R1641 B.n775 B.n774 10.6151
R1642 B.n775 B.n473 10.6151
R1643 B.n781 B.n473 10.6151
R1644 B.n782 B.n781 10.6151
R1645 B.n783 B.n782 10.6151
R1646 B.n783 B.n471 10.6151
R1647 B.n789 B.n471 10.6151
R1648 B.n790 B.n789 10.6151
R1649 B.n791 B.n790 10.6151
R1650 B.n791 B.n469 10.6151
R1651 B.n797 B.n469 10.6151
R1652 B.n798 B.n797 10.6151
R1653 B.n804 B.n803 10.6151
R1654 B.n805 B.n804 10.6151
R1655 B.n805 B.n457 10.6151
R1656 B.n815 B.n457 10.6151
R1657 B.n816 B.n815 10.6151
R1658 B.n817 B.n816 10.6151
R1659 B.n817 B.n449 10.6151
R1660 B.n827 B.n449 10.6151
R1661 B.n828 B.n827 10.6151
R1662 B.n829 B.n828 10.6151
R1663 B.n829 B.n441 10.6151
R1664 B.n839 B.n441 10.6151
R1665 B.n840 B.n839 10.6151
R1666 B.n841 B.n840 10.6151
R1667 B.n841 B.n433 10.6151
R1668 B.n851 B.n433 10.6151
R1669 B.n852 B.n851 10.6151
R1670 B.n853 B.n852 10.6151
R1671 B.n853 B.n425 10.6151
R1672 B.n863 B.n425 10.6151
R1673 B.n864 B.n863 10.6151
R1674 B.n865 B.n864 10.6151
R1675 B.n865 B.n417 10.6151
R1676 B.n875 B.n417 10.6151
R1677 B.n876 B.n875 10.6151
R1678 B.n877 B.n876 10.6151
R1679 B.n877 B.n409 10.6151
R1680 B.n888 B.n409 10.6151
R1681 B.n889 B.n888 10.6151
R1682 B.n890 B.n889 10.6151
R1683 B.n890 B.n402 10.6151
R1684 B.n901 B.n402 10.6151
R1685 B.n902 B.n901 10.6151
R1686 B.n903 B.n902 10.6151
R1687 B.n903 B.n0 10.6151
R1688 B.n1026 B.n1 10.6151
R1689 B.n1026 B.n1025 10.6151
R1690 B.n1025 B.n1024 10.6151
R1691 B.n1024 B.n10 10.6151
R1692 B.n1018 B.n10 10.6151
R1693 B.n1018 B.n1017 10.6151
R1694 B.n1017 B.n1016 10.6151
R1695 B.n1016 B.n16 10.6151
R1696 B.n1010 B.n16 10.6151
R1697 B.n1010 B.n1009 10.6151
R1698 B.n1009 B.n1008 10.6151
R1699 B.n1008 B.n24 10.6151
R1700 B.n1002 B.n24 10.6151
R1701 B.n1002 B.n1001 10.6151
R1702 B.n1001 B.n1000 10.6151
R1703 B.n1000 B.n31 10.6151
R1704 B.n994 B.n31 10.6151
R1705 B.n994 B.n993 10.6151
R1706 B.n993 B.n992 10.6151
R1707 B.n992 B.n38 10.6151
R1708 B.n986 B.n38 10.6151
R1709 B.n986 B.n985 10.6151
R1710 B.n985 B.n984 10.6151
R1711 B.n984 B.n45 10.6151
R1712 B.n978 B.n45 10.6151
R1713 B.n978 B.n977 10.6151
R1714 B.n977 B.n976 10.6151
R1715 B.n976 B.n52 10.6151
R1716 B.n970 B.n52 10.6151
R1717 B.n970 B.n969 10.6151
R1718 B.n969 B.n968 10.6151
R1719 B.n968 B.n59 10.6151
R1720 B.n962 B.n59 10.6151
R1721 B.n962 B.n961 10.6151
R1722 B.n961 B.n960 10.6151
R1723 B.n892 B.t2 8.8172
R1724 B.n1020 B.t1 8.8172
R1725 B.n261 B.n260 6.5566
R1726 B.n277 B.n137 6.5566
R1727 B.n660 B.n507 6.5566
R1728 B.n677 B.n676 6.5566
R1729 B.n825 B.t9 6.03298
R1730 B.n974 B.t5 6.03298
R1731 B.n260 B.n259 4.05904
R1732 B.n280 B.n137 4.05904
R1733 B.n508 B.n507 4.05904
R1734 B.n678 B.n677 4.05904
R1735 B.n1032 B.n0 2.81026
R1736 B.n1032 B.n1 2.81026
R1737 VN.n0 VN.t2 191.249
R1738 VN.n1 VN.t3 191.249
R1739 VN.n0 VN.t1 190.351
R1740 VN.n1 VN.t0 190.351
R1741 VN VN.n1 55.6753
R1742 VN VN.n0 3.43665
R1743 VDD2.n2 VDD2.n0 111.65
R1744 VDD2.n2 VDD2.n1 63.8216
R1745 VDD2.n1 VDD2.t2 1.07484
R1746 VDD2.n1 VDD2.t3 1.07484
R1747 VDD2.n0 VDD2.t0 1.07484
R1748 VDD2.n0 VDD2.t1 1.07484
R1749 VDD2 VDD2.n2 0.0586897
R1750 VTAIL.n5 VTAIL.t0 48.2182
R1751 VTAIL.n4 VTAIL.t4 48.2182
R1752 VTAIL.n3 VTAIL.t7 48.2182
R1753 VTAIL.n7 VTAIL.t6 48.2172
R1754 VTAIL.n0 VTAIL.t5 48.2172
R1755 VTAIL.n1 VTAIL.t1 48.2172
R1756 VTAIL.n2 VTAIL.t3 48.2172
R1757 VTAIL.n6 VTAIL.t2 48.2171
R1758 VTAIL.n7 VTAIL.n6 30.9962
R1759 VTAIL.n3 VTAIL.n2 30.9962
R1760 VTAIL.n4 VTAIL.n3 2.74188
R1761 VTAIL.n6 VTAIL.n5 2.74188
R1762 VTAIL.n2 VTAIL.n1 2.74188
R1763 VTAIL VTAIL.n0 1.42938
R1764 VTAIL VTAIL.n7 1.313
R1765 VTAIL.n5 VTAIL.n4 0.470328
R1766 VTAIL.n1 VTAIL.n0 0.470328
R1767 VP.n4 VP.t0 191.249
R1768 VP.n4 VP.t3 190.351
R1769 VP.n16 VP.n0 161.3
R1770 VP.n15 VP.n14 161.3
R1771 VP.n13 VP.n1 161.3
R1772 VP.n12 VP.n11 161.3
R1773 VP.n10 VP.n2 161.3
R1774 VP.n9 VP.n8 161.3
R1775 VP.n7 VP.n3 161.3
R1776 VP.n5 VP.t1 155.847
R1777 VP.n17 VP.t2 155.847
R1778 VP.n6 VP.n5 106.353
R1779 VP.n18 VP.n17 106.353
R1780 VP.n6 VP.n4 55.3964
R1781 VP.n11 VP.n10 40.4934
R1782 VP.n11 VP.n1 40.4934
R1783 VP.n9 VP.n3 24.4675
R1784 VP.n10 VP.n9 24.4675
R1785 VP.n15 VP.n1 24.4675
R1786 VP.n16 VP.n15 24.4675
R1787 VP.n5 VP.n3 4.40456
R1788 VP.n17 VP.n16 4.40456
R1789 VP.n7 VP.n6 0.278367
R1790 VP.n18 VP.n0 0.278367
R1791 VP.n8 VP.n7 0.189894
R1792 VP.n8 VP.n2 0.189894
R1793 VP.n12 VP.n2 0.189894
R1794 VP.n13 VP.n12 0.189894
R1795 VP.n14 VP.n13 0.189894
R1796 VP.n14 VP.n0 0.189894
R1797 VP VP.n18 0.153454
R1798 VDD1 VDD1.n1 112.174
R1799 VDD1 VDD1.n0 63.8798
R1800 VDD1.n0 VDD1.t3 1.07484
R1801 VDD1.n0 VDD1.t0 1.07484
R1802 VDD1.n1 VDD1.t2 1.07484
R1803 VDD1.n1 VDD1.t1 1.07484
C0 VDD1 VN 0.149065f
C1 VTAIL VP 6.91513f
C2 VDD1 VDD2 1.0826f
C3 VTAIL VN 6.90102f
C4 VN VP 7.56029f
C5 VTAIL VDD2 6.986629f
C6 VP VDD2 0.410052f
C7 VTAIL VDD1 6.93074f
C8 VN VDD2 7.24651f
C9 VDD1 VP 7.5067f
C10 VDD2 B 4.409372f
C11 VDD1 B 9.27781f
C12 VTAIL B 14.094606f
C13 VN B 11.69158f
C14 VP B 9.89332f
C15 VDD1.t3 B 0.388079f
C16 VDD1.t0 B 0.388079f
C17 VDD1.n0 B 3.54931f
C18 VDD1.t2 B 0.388079f
C19 VDD1.t1 B 0.388079f
C20 VDD1.n1 B 4.47846f
C21 VP.n0 B 0.030402f
C22 VP.t2 B 3.33306f
C23 VP.n1 B 0.045832f
C24 VP.n2 B 0.02306f
C25 VP.n3 B 0.025579f
C26 VP.t3 B 3.57035f
C27 VP.t0 B 3.57634f
C28 VP.n4 B 3.75103f
C29 VP.t1 B 3.33306f
C30 VP.n5 B 1.2306f
C31 VP.n6 B 1.47839f
C32 VP.n7 B 0.030402f
C33 VP.n8 B 0.02306f
C34 VP.n9 B 0.042978f
C35 VP.n10 B 0.045832f
C36 VP.n11 B 0.018642f
C37 VP.n12 B 0.02306f
C38 VP.n13 B 0.02306f
C39 VP.n14 B 0.02306f
C40 VP.n15 B 0.042978f
C41 VP.n16 B 0.025579f
C42 VP.n17 B 1.2306f
C43 VP.n18 B 0.042686f
C44 VTAIL.t5 B 2.55528f
C45 VTAIL.n0 B 0.2898f
C46 VTAIL.t1 B 2.55528f
C47 VTAIL.n1 B 0.354629f
C48 VTAIL.t3 B 2.55528f
C49 VTAIL.n2 B 1.45981f
C50 VTAIL.t7 B 2.55527f
C51 VTAIL.n3 B 1.45982f
C52 VTAIL.t4 B 2.55527f
C53 VTAIL.n4 B 0.354636f
C54 VTAIL.t0 B 2.55527f
C55 VTAIL.n5 B 0.354636f
C56 VTAIL.t2 B 2.55527f
C57 VTAIL.n6 B 1.45982f
C58 VTAIL.t6 B 2.55528f
C59 VTAIL.n7 B 1.38924f
C60 VDD2.t0 B 0.385323f
C61 VDD2.t1 B 0.385323f
C62 VDD2.n0 B 4.41871f
C63 VDD2.t2 B 0.385323f
C64 VDD2.t3 B 0.385323f
C65 VDD2.n1 B 3.52368f
C66 VDD2.n2 B 4.47692f
C67 VN.t2 B 3.52238f
C68 VN.t1 B 3.51648f
C69 VN.n0 B 2.23148f
C70 VN.t3 B 3.52238f
C71 VN.t0 B 3.51648f
C72 VN.n1 B 3.70631f
.ends

