* NGSPICE file created from diff_pair_sample_1058.ext - technology: sky130A

.subckt diff_pair_sample_1058 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t3 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=2.1186 ps=13.17 w=12.84 l=2.05
X1 VDD1.t4 VP.t1 VTAIL.t9 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=5.0076 ps=26.46 w=12.84 l=2.05
X2 VDD2.t5 VN.t0 VTAIL.t0 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=5.0076 ps=26.46 w=12.84 l=2.05
X3 VTAIL.t4 VN.t1 VDD2.t4 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=2.1186 ps=13.17 w=12.84 l=2.05
X4 VDD1.t1 VP.t2 VTAIL.t8 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=5.0076 ps=26.46 w=12.84 l=2.05
X5 VDD1.t2 VP.t3 VTAIL.t7 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=2.1186 ps=13.17 w=12.84 l=2.05
X6 B.t11 B.t9 B.t10 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=0 ps=0 w=12.84 l=2.05
X7 VDD2.t3 VN.t2 VTAIL.t11 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=5.0076 ps=26.46 w=12.84 l=2.05
X8 VTAIL.t1 VN.t3 VDD2.t2 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=2.1186 ps=13.17 w=12.84 l=2.05
X9 B.t8 B.t6 B.t7 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=0 ps=0 w=12.84 l=2.05
X10 VTAIL.t6 VP.t4 VDD1.t0 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=2.1186 pd=13.17 as=2.1186 ps=13.17 w=12.84 l=2.05
X11 B.t5 B.t3 B.t4 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=0 ps=0 w=12.84 l=2.05
X12 VDD1.t5 VP.t5 VTAIL.t5 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=2.1186 ps=13.17 w=12.84 l=2.05
X13 VDD2.t1 VN.t4 VTAIL.t3 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=2.1186 ps=13.17 w=12.84 l=2.05
X14 B.t2 B.t0 B.t1 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=0 ps=0 w=12.84 l=2.05
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n2874_n3536# sky130_fd_pr__pfet_01v8 ad=5.0076 pd=26.46 as=2.1186 ps=13.17 w=12.84 l=2.05
R0 VP.n7 VP.t5 184.941
R1 VP.n10 VP.n9 161.3
R2 VP.n11 VP.n6 161.3
R3 VP.n13 VP.n12 161.3
R4 VP.n14 VP.n5 161.3
R5 VP.n31 VP.n0 161.3
R6 VP.n30 VP.n29 161.3
R7 VP.n28 VP.n1 161.3
R8 VP.n27 VP.n26 161.3
R9 VP.n25 VP.n2 161.3
R10 VP.n24 VP.n23 161.3
R11 VP.n22 VP.n3 161.3
R12 VP.n21 VP.n20 161.3
R13 VP.n19 VP.n4 161.3
R14 VP.n25 VP.t4 150.948
R15 VP.n18 VP.t3 150.948
R16 VP.n32 VP.t1 150.948
R17 VP.n8 VP.t0 150.948
R18 VP.n15 VP.t2 150.948
R19 VP.n18 VP.n17 92.2184
R20 VP.n33 VP.n32 92.2184
R21 VP.n16 VP.n15 92.2184
R22 VP.n20 VP.n3 56.5617
R23 VP.n30 VP.n1 56.5617
R24 VP.n13 VP.n6 56.5617
R25 VP.n17 VP.n16 47.1739
R26 VP.n8 VP.n7 46.044
R27 VP.n20 VP.n19 24.5923
R28 VP.n24 VP.n3 24.5923
R29 VP.n25 VP.n24 24.5923
R30 VP.n26 VP.n25 24.5923
R31 VP.n26 VP.n1 24.5923
R32 VP.n31 VP.n30 24.5923
R33 VP.n14 VP.n13 24.5923
R34 VP.n9 VP.n8 24.5923
R35 VP.n9 VP.n6 24.5923
R36 VP.n19 VP.n18 18.6903
R37 VP.n32 VP.n31 18.6903
R38 VP.n15 VP.n14 18.6903
R39 VP.n10 VP.n7 9.07974
R40 VP.n16 VP.n5 0.278335
R41 VP.n17 VP.n4 0.278335
R42 VP.n33 VP.n0 0.278335
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153485
R55 VDD1.n64 VDD1.n0 756.745
R56 VDD1.n133 VDD1.n69 756.745
R57 VDD1.n65 VDD1.n64 585
R58 VDD1.n63 VDD1.n62 585
R59 VDD1.n4 VDD1.n3 585
R60 VDD1.n57 VDD1.n56 585
R61 VDD1.n55 VDD1.n54 585
R62 VDD1.n8 VDD1.n7 585
R63 VDD1.n49 VDD1.n48 585
R64 VDD1.n47 VDD1.n46 585
R65 VDD1.n45 VDD1.n11 585
R66 VDD1.n15 VDD1.n12 585
R67 VDD1.n40 VDD1.n39 585
R68 VDD1.n38 VDD1.n37 585
R69 VDD1.n17 VDD1.n16 585
R70 VDD1.n32 VDD1.n31 585
R71 VDD1.n30 VDD1.n29 585
R72 VDD1.n21 VDD1.n20 585
R73 VDD1.n24 VDD1.n23 585
R74 VDD1.n92 VDD1.n91 585
R75 VDD1.n89 VDD1.n88 585
R76 VDD1.n98 VDD1.n97 585
R77 VDD1.n100 VDD1.n99 585
R78 VDD1.n85 VDD1.n84 585
R79 VDD1.n106 VDD1.n105 585
R80 VDD1.n109 VDD1.n108 585
R81 VDD1.n107 VDD1.n81 585
R82 VDD1.n114 VDD1.n80 585
R83 VDD1.n116 VDD1.n115 585
R84 VDD1.n118 VDD1.n117 585
R85 VDD1.n77 VDD1.n76 585
R86 VDD1.n124 VDD1.n123 585
R87 VDD1.n126 VDD1.n125 585
R88 VDD1.n73 VDD1.n72 585
R89 VDD1.n132 VDD1.n131 585
R90 VDD1.n134 VDD1.n133 585
R91 VDD1.t2 VDD1.n90 329.036
R92 VDD1.t5 VDD1.n22 329.036
R93 VDD1.n64 VDD1.n63 171.744
R94 VDD1.n63 VDD1.n3 171.744
R95 VDD1.n56 VDD1.n3 171.744
R96 VDD1.n56 VDD1.n55 171.744
R97 VDD1.n55 VDD1.n7 171.744
R98 VDD1.n48 VDD1.n7 171.744
R99 VDD1.n48 VDD1.n47 171.744
R100 VDD1.n47 VDD1.n11 171.744
R101 VDD1.n15 VDD1.n11 171.744
R102 VDD1.n39 VDD1.n15 171.744
R103 VDD1.n39 VDD1.n38 171.744
R104 VDD1.n38 VDD1.n16 171.744
R105 VDD1.n31 VDD1.n16 171.744
R106 VDD1.n31 VDD1.n30 171.744
R107 VDD1.n30 VDD1.n20 171.744
R108 VDD1.n23 VDD1.n20 171.744
R109 VDD1.n91 VDD1.n88 171.744
R110 VDD1.n98 VDD1.n88 171.744
R111 VDD1.n99 VDD1.n98 171.744
R112 VDD1.n99 VDD1.n84 171.744
R113 VDD1.n106 VDD1.n84 171.744
R114 VDD1.n108 VDD1.n106 171.744
R115 VDD1.n108 VDD1.n107 171.744
R116 VDD1.n107 VDD1.n80 171.744
R117 VDD1.n116 VDD1.n80 171.744
R118 VDD1.n117 VDD1.n116 171.744
R119 VDD1.n117 VDD1.n76 171.744
R120 VDD1.n124 VDD1.n76 171.744
R121 VDD1.n125 VDD1.n124 171.744
R122 VDD1.n125 VDD1.n72 171.744
R123 VDD1.n132 VDD1.n72 171.744
R124 VDD1.n133 VDD1.n132 171.744
R125 VDD1.n23 VDD1.t5 85.8723
R126 VDD1.n91 VDD1.t2 85.8723
R127 VDD1.n139 VDD1.n138 73.469
R128 VDD1.n141 VDD1.n140 73.0112
R129 VDD1 VDD1.n68 50.4611
R130 VDD1.n139 VDD1.n137 50.3476
R131 VDD1.n141 VDD1.n139 43.0612
R132 VDD1.n46 VDD1.n45 13.1884
R133 VDD1.n115 VDD1.n114 13.1884
R134 VDD1.n49 VDD1.n10 12.8005
R135 VDD1.n44 VDD1.n12 12.8005
R136 VDD1.n113 VDD1.n81 12.8005
R137 VDD1.n118 VDD1.n79 12.8005
R138 VDD1.n50 VDD1.n8 12.0247
R139 VDD1.n41 VDD1.n40 12.0247
R140 VDD1.n110 VDD1.n109 12.0247
R141 VDD1.n119 VDD1.n77 12.0247
R142 VDD1.n54 VDD1.n53 11.249
R143 VDD1.n37 VDD1.n14 11.249
R144 VDD1.n105 VDD1.n83 11.249
R145 VDD1.n123 VDD1.n122 11.249
R146 VDD1.n24 VDD1.n22 10.7239
R147 VDD1.n92 VDD1.n90 10.7239
R148 VDD1.n57 VDD1.n6 10.4732
R149 VDD1.n36 VDD1.n17 10.4732
R150 VDD1.n104 VDD1.n85 10.4732
R151 VDD1.n126 VDD1.n75 10.4732
R152 VDD1.n58 VDD1.n4 9.69747
R153 VDD1.n33 VDD1.n32 9.69747
R154 VDD1.n101 VDD1.n100 9.69747
R155 VDD1.n127 VDD1.n73 9.69747
R156 VDD1.n68 VDD1.n67 9.45567
R157 VDD1.n137 VDD1.n136 9.45567
R158 VDD1.n26 VDD1.n25 9.3005
R159 VDD1.n28 VDD1.n27 9.3005
R160 VDD1.n19 VDD1.n18 9.3005
R161 VDD1.n34 VDD1.n33 9.3005
R162 VDD1.n36 VDD1.n35 9.3005
R163 VDD1.n14 VDD1.n13 9.3005
R164 VDD1.n42 VDD1.n41 9.3005
R165 VDD1.n44 VDD1.n43 9.3005
R166 VDD1.n67 VDD1.n66 9.3005
R167 VDD1.n2 VDD1.n1 9.3005
R168 VDD1.n61 VDD1.n60 9.3005
R169 VDD1.n59 VDD1.n58 9.3005
R170 VDD1.n6 VDD1.n5 9.3005
R171 VDD1.n53 VDD1.n52 9.3005
R172 VDD1.n51 VDD1.n50 9.3005
R173 VDD1.n10 VDD1.n9 9.3005
R174 VDD1.n71 VDD1.n70 9.3005
R175 VDD1.n130 VDD1.n129 9.3005
R176 VDD1.n128 VDD1.n127 9.3005
R177 VDD1.n75 VDD1.n74 9.3005
R178 VDD1.n122 VDD1.n121 9.3005
R179 VDD1.n120 VDD1.n119 9.3005
R180 VDD1.n79 VDD1.n78 9.3005
R181 VDD1.n94 VDD1.n93 9.3005
R182 VDD1.n96 VDD1.n95 9.3005
R183 VDD1.n87 VDD1.n86 9.3005
R184 VDD1.n102 VDD1.n101 9.3005
R185 VDD1.n104 VDD1.n103 9.3005
R186 VDD1.n83 VDD1.n82 9.3005
R187 VDD1.n111 VDD1.n110 9.3005
R188 VDD1.n113 VDD1.n112 9.3005
R189 VDD1.n136 VDD1.n135 9.3005
R190 VDD1.n62 VDD1.n61 8.92171
R191 VDD1.n29 VDD1.n19 8.92171
R192 VDD1.n97 VDD1.n87 8.92171
R193 VDD1.n131 VDD1.n130 8.92171
R194 VDD1.n65 VDD1.n2 8.14595
R195 VDD1.n28 VDD1.n21 8.14595
R196 VDD1.n96 VDD1.n89 8.14595
R197 VDD1.n134 VDD1.n71 8.14595
R198 VDD1.n66 VDD1.n0 7.3702
R199 VDD1.n25 VDD1.n24 7.3702
R200 VDD1.n93 VDD1.n92 7.3702
R201 VDD1.n135 VDD1.n69 7.3702
R202 VDD1.n68 VDD1.n0 6.59444
R203 VDD1.n137 VDD1.n69 6.59444
R204 VDD1.n66 VDD1.n65 5.81868
R205 VDD1.n25 VDD1.n21 5.81868
R206 VDD1.n93 VDD1.n89 5.81868
R207 VDD1.n135 VDD1.n134 5.81868
R208 VDD1.n62 VDD1.n2 5.04292
R209 VDD1.n29 VDD1.n28 5.04292
R210 VDD1.n97 VDD1.n96 5.04292
R211 VDD1.n131 VDD1.n71 5.04292
R212 VDD1.n61 VDD1.n4 4.26717
R213 VDD1.n32 VDD1.n19 4.26717
R214 VDD1.n100 VDD1.n87 4.26717
R215 VDD1.n130 VDD1.n73 4.26717
R216 VDD1.n58 VDD1.n57 3.49141
R217 VDD1.n33 VDD1.n17 3.49141
R218 VDD1.n101 VDD1.n85 3.49141
R219 VDD1.n127 VDD1.n126 3.49141
R220 VDD1.n54 VDD1.n6 2.71565
R221 VDD1.n37 VDD1.n36 2.71565
R222 VDD1.n105 VDD1.n104 2.71565
R223 VDD1.n123 VDD1.n75 2.71565
R224 VDD1.n140 VDD1.t3 2.53204
R225 VDD1.n140 VDD1.t1 2.53204
R226 VDD1.n138 VDD1.t0 2.53204
R227 VDD1.n138 VDD1.t4 2.53204
R228 VDD1.n26 VDD1.n22 2.41282
R229 VDD1.n94 VDD1.n90 2.41282
R230 VDD1.n53 VDD1.n8 1.93989
R231 VDD1.n40 VDD1.n14 1.93989
R232 VDD1.n109 VDD1.n83 1.93989
R233 VDD1.n122 VDD1.n77 1.93989
R234 VDD1.n50 VDD1.n49 1.16414
R235 VDD1.n41 VDD1.n12 1.16414
R236 VDD1.n110 VDD1.n81 1.16414
R237 VDD1.n119 VDD1.n118 1.16414
R238 VDD1 VDD1.n141 0.455241
R239 VDD1.n46 VDD1.n10 0.388379
R240 VDD1.n45 VDD1.n44 0.388379
R241 VDD1.n114 VDD1.n113 0.388379
R242 VDD1.n115 VDD1.n79 0.388379
R243 VDD1.n67 VDD1.n1 0.155672
R244 VDD1.n60 VDD1.n1 0.155672
R245 VDD1.n60 VDD1.n59 0.155672
R246 VDD1.n59 VDD1.n5 0.155672
R247 VDD1.n52 VDD1.n5 0.155672
R248 VDD1.n52 VDD1.n51 0.155672
R249 VDD1.n51 VDD1.n9 0.155672
R250 VDD1.n43 VDD1.n9 0.155672
R251 VDD1.n43 VDD1.n42 0.155672
R252 VDD1.n42 VDD1.n13 0.155672
R253 VDD1.n35 VDD1.n13 0.155672
R254 VDD1.n35 VDD1.n34 0.155672
R255 VDD1.n34 VDD1.n18 0.155672
R256 VDD1.n27 VDD1.n18 0.155672
R257 VDD1.n27 VDD1.n26 0.155672
R258 VDD1.n95 VDD1.n94 0.155672
R259 VDD1.n95 VDD1.n86 0.155672
R260 VDD1.n102 VDD1.n86 0.155672
R261 VDD1.n103 VDD1.n102 0.155672
R262 VDD1.n103 VDD1.n82 0.155672
R263 VDD1.n111 VDD1.n82 0.155672
R264 VDD1.n112 VDD1.n111 0.155672
R265 VDD1.n112 VDD1.n78 0.155672
R266 VDD1.n120 VDD1.n78 0.155672
R267 VDD1.n121 VDD1.n120 0.155672
R268 VDD1.n121 VDD1.n74 0.155672
R269 VDD1.n128 VDD1.n74 0.155672
R270 VDD1.n129 VDD1.n128 0.155672
R271 VDD1.n129 VDD1.n70 0.155672
R272 VDD1.n136 VDD1.n70 0.155672
R273 VTAIL.n282 VTAIL.n218 756.745
R274 VTAIL.n66 VTAIL.n2 756.745
R275 VTAIL.n212 VTAIL.n148 756.745
R276 VTAIL.n140 VTAIL.n76 756.745
R277 VTAIL.n241 VTAIL.n240 585
R278 VTAIL.n238 VTAIL.n237 585
R279 VTAIL.n247 VTAIL.n246 585
R280 VTAIL.n249 VTAIL.n248 585
R281 VTAIL.n234 VTAIL.n233 585
R282 VTAIL.n255 VTAIL.n254 585
R283 VTAIL.n258 VTAIL.n257 585
R284 VTAIL.n256 VTAIL.n230 585
R285 VTAIL.n263 VTAIL.n229 585
R286 VTAIL.n265 VTAIL.n264 585
R287 VTAIL.n267 VTAIL.n266 585
R288 VTAIL.n226 VTAIL.n225 585
R289 VTAIL.n273 VTAIL.n272 585
R290 VTAIL.n275 VTAIL.n274 585
R291 VTAIL.n222 VTAIL.n221 585
R292 VTAIL.n281 VTAIL.n280 585
R293 VTAIL.n283 VTAIL.n282 585
R294 VTAIL.n25 VTAIL.n24 585
R295 VTAIL.n22 VTAIL.n21 585
R296 VTAIL.n31 VTAIL.n30 585
R297 VTAIL.n33 VTAIL.n32 585
R298 VTAIL.n18 VTAIL.n17 585
R299 VTAIL.n39 VTAIL.n38 585
R300 VTAIL.n42 VTAIL.n41 585
R301 VTAIL.n40 VTAIL.n14 585
R302 VTAIL.n47 VTAIL.n13 585
R303 VTAIL.n49 VTAIL.n48 585
R304 VTAIL.n51 VTAIL.n50 585
R305 VTAIL.n10 VTAIL.n9 585
R306 VTAIL.n57 VTAIL.n56 585
R307 VTAIL.n59 VTAIL.n58 585
R308 VTAIL.n6 VTAIL.n5 585
R309 VTAIL.n65 VTAIL.n64 585
R310 VTAIL.n67 VTAIL.n66 585
R311 VTAIL.n213 VTAIL.n212 585
R312 VTAIL.n211 VTAIL.n210 585
R313 VTAIL.n152 VTAIL.n151 585
R314 VTAIL.n205 VTAIL.n204 585
R315 VTAIL.n203 VTAIL.n202 585
R316 VTAIL.n156 VTAIL.n155 585
R317 VTAIL.n197 VTAIL.n196 585
R318 VTAIL.n195 VTAIL.n194 585
R319 VTAIL.n193 VTAIL.n159 585
R320 VTAIL.n163 VTAIL.n160 585
R321 VTAIL.n188 VTAIL.n187 585
R322 VTAIL.n186 VTAIL.n185 585
R323 VTAIL.n165 VTAIL.n164 585
R324 VTAIL.n180 VTAIL.n179 585
R325 VTAIL.n178 VTAIL.n177 585
R326 VTAIL.n169 VTAIL.n168 585
R327 VTAIL.n172 VTAIL.n171 585
R328 VTAIL.n141 VTAIL.n140 585
R329 VTAIL.n139 VTAIL.n138 585
R330 VTAIL.n80 VTAIL.n79 585
R331 VTAIL.n133 VTAIL.n132 585
R332 VTAIL.n131 VTAIL.n130 585
R333 VTAIL.n84 VTAIL.n83 585
R334 VTAIL.n125 VTAIL.n124 585
R335 VTAIL.n123 VTAIL.n122 585
R336 VTAIL.n121 VTAIL.n87 585
R337 VTAIL.n91 VTAIL.n88 585
R338 VTAIL.n116 VTAIL.n115 585
R339 VTAIL.n114 VTAIL.n113 585
R340 VTAIL.n93 VTAIL.n92 585
R341 VTAIL.n108 VTAIL.n107 585
R342 VTAIL.n106 VTAIL.n105 585
R343 VTAIL.n97 VTAIL.n96 585
R344 VTAIL.n100 VTAIL.n99 585
R345 VTAIL.t11 VTAIL.n239 329.036
R346 VTAIL.t9 VTAIL.n23 329.036
R347 VTAIL.t8 VTAIL.n170 329.036
R348 VTAIL.t0 VTAIL.n98 329.036
R349 VTAIL.n240 VTAIL.n237 171.744
R350 VTAIL.n247 VTAIL.n237 171.744
R351 VTAIL.n248 VTAIL.n247 171.744
R352 VTAIL.n248 VTAIL.n233 171.744
R353 VTAIL.n255 VTAIL.n233 171.744
R354 VTAIL.n257 VTAIL.n255 171.744
R355 VTAIL.n257 VTAIL.n256 171.744
R356 VTAIL.n256 VTAIL.n229 171.744
R357 VTAIL.n265 VTAIL.n229 171.744
R358 VTAIL.n266 VTAIL.n265 171.744
R359 VTAIL.n266 VTAIL.n225 171.744
R360 VTAIL.n273 VTAIL.n225 171.744
R361 VTAIL.n274 VTAIL.n273 171.744
R362 VTAIL.n274 VTAIL.n221 171.744
R363 VTAIL.n281 VTAIL.n221 171.744
R364 VTAIL.n282 VTAIL.n281 171.744
R365 VTAIL.n24 VTAIL.n21 171.744
R366 VTAIL.n31 VTAIL.n21 171.744
R367 VTAIL.n32 VTAIL.n31 171.744
R368 VTAIL.n32 VTAIL.n17 171.744
R369 VTAIL.n39 VTAIL.n17 171.744
R370 VTAIL.n41 VTAIL.n39 171.744
R371 VTAIL.n41 VTAIL.n40 171.744
R372 VTAIL.n40 VTAIL.n13 171.744
R373 VTAIL.n49 VTAIL.n13 171.744
R374 VTAIL.n50 VTAIL.n49 171.744
R375 VTAIL.n50 VTAIL.n9 171.744
R376 VTAIL.n57 VTAIL.n9 171.744
R377 VTAIL.n58 VTAIL.n57 171.744
R378 VTAIL.n58 VTAIL.n5 171.744
R379 VTAIL.n65 VTAIL.n5 171.744
R380 VTAIL.n66 VTAIL.n65 171.744
R381 VTAIL.n212 VTAIL.n211 171.744
R382 VTAIL.n211 VTAIL.n151 171.744
R383 VTAIL.n204 VTAIL.n151 171.744
R384 VTAIL.n204 VTAIL.n203 171.744
R385 VTAIL.n203 VTAIL.n155 171.744
R386 VTAIL.n196 VTAIL.n155 171.744
R387 VTAIL.n196 VTAIL.n195 171.744
R388 VTAIL.n195 VTAIL.n159 171.744
R389 VTAIL.n163 VTAIL.n159 171.744
R390 VTAIL.n187 VTAIL.n163 171.744
R391 VTAIL.n187 VTAIL.n186 171.744
R392 VTAIL.n186 VTAIL.n164 171.744
R393 VTAIL.n179 VTAIL.n164 171.744
R394 VTAIL.n179 VTAIL.n178 171.744
R395 VTAIL.n178 VTAIL.n168 171.744
R396 VTAIL.n171 VTAIL.n168 171.744
R397 VTAIL.n140 VTAIL.n139 171.744
R398 VTAIL.n139 VTAIL.n79 171.744
R399 VTAIL.n132 VTAIL.n79 171.744
R400 VTAIL.n132 VTAIL.n131 171.744
R401 VTAIL.n131 VTAIL.n83 171.744
R402 VTAIL.n124 VTAIL.n83 171.744
R403 VTAIL.n124 VTAIL.n123 171.744
R404 VTAIL.n123 VTAIL.n87 171.744
R405 VTAIL.n91 VTAIL.n87 171.744
R406 VTAIL.n115 VTAIL.n91 171.744
R407 VTAIL.n115 VTAIL.n114 171.744
R408 VTAIL.n114 VTAIL.n92 171.744
R409 VTAIL.n107 VTAIL.n92 171.744
R410 VTAIL.n107 VTAIL.n106 171.744
R411 VTAIL.n106 VTAIL.n96 171.744
R412 VTAIL.n99 VTAIL.n96 171.744
R413 VTAIL.n240 VTAIL.t11 85.8723
R414 VTAIL.n24 VTAIL.t9 85.8723
R415 VTAIL.n171 VTAIL.t8 85.8723
R416 VTAIL.n99 VTAIL.t0 85.8723
R417 VTAIL.n1 VTAIL.n0 56.3326
R418 VTAIL.n73 VTAIL.n72 56.3326
R419 VTAIL.n147 VTAIL.n146 56.3326
R420 VTAIL.n75 VTAIL.n74 56.3326
R421 VTAIL.n287 VTAIL.n286 32.1853
R422 VTAIL.n71 VTAIL.n70 32.1853
R423 VTAIL.n217 VTAIL.n216 32.1853
R424 VTAIL.n145 VTAIL.n144 32.1853
R425 VTAIL.n75 VTAIL.n73 27.5393
R426 VTAIL.n287 VTAIL.n217 25.4876
R427 VTAIL.n264 VTAIL.n263 13.1884
R428 VTAIL.n48 VTAIL.n47 13.1884
R429 VTAIL.n194 VTAIL.n193 13.1884
R430 VTAIL.n122 VTAIL.n121 13.1884
R431 VTAIL.n262 VTAIL.n230 12.8005
R432 VTAIL.n267 VTAIL.n228 12.8005
R433 VTAIL.n46 VTAIL.n14 12.8005
R434 VTAIL.n51 VTAIL.n12 12.8005
R435 VTAIL.n197 VTAIL.n158 12.8005
R436 VTAIL.n192 VTAIL.n160 12.8005
R437 VTAIL.n125 VTAIL.n86 12.8005
R438 VTAIL.n120 VTAIL.n88 12.8005
R439 VTAIL.n259 VTAIL.n258 12.0247
R440 VTAIL.n268 VTAIL.n226 12.0247
R441 VTAIL.n43 VTAIL.n42 12.0247
R442 VTAIL.n52 VTAIL.n10 12.0247
R443 VTAIL.n198 VTAIL.n156 12.0247
R444 VTAIL.n189 VTAIL.n188 12.0247
R445 VTAIL.n126 VTAIL.n84 12.0247
R446 VTAIL.n117 VTAIL.n116 12.0247
R447 VTAIL.n254 VTAIL.n232 11.249
R448 VTAIL.n272 VTAIL.n271 11.249
R449 VTAIL.n38 VTAIL.n16 11.249
R450 VTAIL.n56 VTAIL.n55 11.249
R451 VTAIL.n202 VTAIL.n201 11.249
R452 VTAIL.n185 VTAIL.n162 11.249
R453 VTAIL.n130 VTAIL.n129 11.249
R454 VTAIL.n113 VTAIL.n90 11.249
R455 VTAIL.n241 VTAIL.n239 10.7239
R456 VTAIL.n25 VTAIL.n23 10.7239
R457 VTAIL.n172 VTAIL.n170 10.7239
R458 VTAIL.n100 VTAIL.n98 10.7239
R459 VTAIL.n253 VTAIL.n234 10.4732
R460 VTAIL.n275 VTAIL.n224 10.4732
R461 VTAIL.n37 VTAIL.n18 10.4732
R462 VTAIL.n59 VTAIL.n8 10.4732
R463 VTAIL.n205 VTAIL.n154 10.4732
R464 VTAIL.n184 VTAIL.n165 10.4732
R465 VTAIL.n133 VTAIL.n82 10.4732
R466 VTAIL.n112 VTAIL.n93 10.4732
R467 VTAIL.n250 VTAIL.n249 9.69747
R468 VTAIL.n276 VTAIL.n222 9.69747
R469 VTAIL.n34 VTAIL.n33 9.69747
R470 VTAIL.n60 VTAIL.n6 9.69747
R471 VTAIL.n206 VTAIL.n152 9.69747
R472 VTAIL.n181 VTAIL.n180 9.69747
R473 VTAIL.n134 VTAIL.n80 9.69747
R474 VTAIL.n109 VTAIL.n108 9.69747
R475 VTAIL.n286 VTAIL.n285 9.45567
R476 VTAIL.n70 VTAIL.n69 9.45567
R477 VTAIL.n216 VTAIL.n215 9.45567
R478 VTAIL.n144 VTAIL.n143 9.45567
R479 VTAIL.n220 VTAIL.n219 9.3005
R480 VTAIL.n279 VTAIL.n278 9.3005
R481 VTAIL.n277 VTAIL.n276 9.3005
R482 VTAIL.n224 VTAIL.n223 9.3005
R483 VTAIL.n271 VTAIL.n270 9.3005
R484 VTAIL.n269 VTAIL.n268 9.3005
R485 VTAIL.n228 VTAIL.n227 9.3005
R486 VTAIL.n243 VTAIL.n242 9.3005
R487 VTAIL.n245 VTAIL.n244 9.3005
R488 VTAIL.n236 VTAIL.n235 9.3005
R489 VTAIL.n251 VTAIL.n250 9.3005
R490 VTAIL.n253 VTAIL.n252 9.3005
R491 VTAIL.n232 VTAIL.n231 9.3005
R492 VTAIL.n260 VTAIL.n259 9.3005
R493 VTAIL.n262 VTAIL.n261 9.3005
R494 VTAIL.n285 VTAIL.n284 9.3005
R495 VTAIL.n4 VTAIL.n3 9.3005
R496 VTAIL.n63 VTAIL.n62 9.3005
R497 VTAIL.n61 VTAIL.n60 9.3005
R498 VTAIL.n8 VTAIL.n7 9.3005
R499 VTAIL.n55 VTAIL.n54 9.3005
R500 VTAIL.n53 VTAIL.n52 9.3005
R501 VTAIL.n12 VTAIL.n11 9.3005
R502 VTAIL.n27 VTAIL.n26 9.3005
R503 VTAIL.n29 VTAIL.n28 9.3005
R504 VTAIL.n20 VTAIL.n19 9.3005
R505 VTAIL.n35 VTAIL.n34 9.3005
R506 VTAIL.n37 VTAIL.n36 9.3005
R507 VTAIL.n16 VTAIL.n15 9.3005
R508 VTAIL.n44 VTAIL.n43 9.3005
R509 VTAIL.n46 VTAIL.n45 9.3005
R510 VTAIL.n69 VTAIL.n68 9.3005
R511 VTAIL.n174 VTAIL.n173 9.3005
R512 VTAIL.n176 VTAIL.n175 9.3005
R513 VTAIL.n167 VTAIL.n166 9.3005
R514 VTAIL.n182 VTAIL.n181 9.3005
R515 VTAIL.n184 VTAIL.n183 9.3005
R516 VTAIL.n162 VTAIL.n161 9.3005
R517 VTAIL.n190 VTAIL.n189 9.3005
R518 VTAIL.n192 VTAIL.n191 9.3005
R519 VTAIL.n215 VTAIL.n214 9.3005
R520 VTAIL.n150 VTAIL.n149 9.3005
R521 VTAIL.n209 VTAIL.n208 9.3005
R522 VTAIL.n207 VTAIL.n206 9.3005
R523 VTAIL.n154 VTAIL.n153 9.3005
R524 VTAIL.n201 VTAIL.n200 9.3005
R525 VTAIL.n199 VTAIL.n198 9.3005
R526 VTAIL.n158 VTAIL.n157 9.3005
R527 VTAIL.n102 VTAIL.n101 9.3005
R528 VTAIL.n104 VTAIL.n103 9.3005
R529 VTAIL.n95 VTAIL.n94 9.3005
R530 VTAIL.n110 VTAIL.n109 9.3005
R531 VTAIL.n112 VTAIL.n111 9.3005
R532 VTAIL.n90 VTAIL.n89 9.3005
R533 VTAIL.n118 VTAIL.n117 9.3005
R534 VTAIL.n120 VTAIL.n119 9.3005
R535 VTAIL.n143 VTAIL.n142 9.3005
R536 VTAIL.n78 VTAIL.n77 9.3005
R537 VTAIL.n137 VTAIL.n136 9.3005
R538 VTAIL.n135 VTAIL.n134 9.3005
R539 VTAIL.n82 VTAIL.n81 9.3005
R540 VTAIL.n129 VTAIL.n128 9.3005
R541 VTAIL.n127 VTAIL.n126 9.3005
R542 VTAIL.n86 VTAIL.n85 9.3005
R543 VTAIL.n246 VTAIL.n236 8.92171
R544 VTAIL.n280 VTAIL.n279 8.92171
R545 VTAIL.n30 VTAIL.n20 8.92171
R546 VTAIL.n64 VTAIL.n63 8.92171
R547 VTAIL.n210 VTAIL.n209 8.92171
R548 VTAIL.n177 VTAIL.n167 8.92171
R549 VTAIL.n138 VTAIL.n137 8.92171
R550 VTAIL.n105 VTAIL.n95 8.92171
R551 VTAIL.n245 VTAIL.n238 8.14595
R552 VTAIL.n283 VTAIL.n220 8.14595
R553 VTAIL.n29 VTAIL.n22 8.14595
R554 VTAIL.n67 VTAIL.n4 8.14595
R555 VTAIL.n213 VTAIL.n150 8.14595
R556 VTAIL.n176 VTAIL.n169 8.14595
R557 VTAIL.n141 VTAIL.n78 8.14595
R558 VTAIL.n104 VTAIL.n97 8.14595
R559 VTAIL.n242 VTAIL.n241 7.3702
R560 VTAIL.n284 VTAIL.n218 7.3702
R561 VTAIL.n26 VTAIL.n25 7.3702
R562 VTAIL.n68 VTAIL.n2 7.3702
R563 VTAIL.n214 VTAIL.n148 7.3702
R564 VTAIL.n173 VTAIL.n172 7.3702
R565 VTAIL.n142 VTAIL.n76 7.3702
R566 VTAIL.n101 VTAIL.n100 7.3702
R567 VTAIL.n286 VTAIL.n218 6.59444
R568 VTAIL.n70 VTAIL.n2 6.59444
R569 VTAIL.n216 VTAIL.n148 6.59444
R570 VTAIL.n144 VTAIL.n76 6.59444
R571 VTAIL.n242 VTAIL.n238 5.81868
R572 VTAIL.n284 VTAIL.n283 5.81868
R573 VTAIL.n26 VTAIL.n22 5.81868
R574 VTAIL.n68 VTAIL.n67 5.81868
R575 VTAIL.n214 VTAIL.n213 5.81868
R576 VTAIL.n173 VTAIL.n169 5.81868
R577 VTAIL.n142 VTAIL.n141 5.81868
R578 VTAIL.n101 VTAIL.n97 5.81868
R579 VTAIL.n246 VTAIL.n245 5.04292
R580 VTAIL.n280 VTAIL.n220 5.04292
R581 VTAIL.n30 VTAIL.n29 5.04292
R582 VTAIL.n64 VTAIL.n4 5.04292
R583 VTAIL.n210 VTAIL.n150 5.04292
R584 VTAIL.n177 VTAIL.n176 5.04292
R585 VTAIL.n138 VTAIL.n78 5.04292
R586 VTAIL.n105 VTAIL.n104 5.04292
R587 VTAIL.n249 VTAIL.n236 4.26717
R588 VTAIL.n279 VTAIL.n222 4.26717
R589 VTAIL.n33 VTAIL.n20 4.26717
R590 VTAIL.n63 VTAIL.n6 4.26717
R591 VTAIL.n209 VTAIL.n152 4.26717
R592 VTAIL.n180 VTAIL.n167 4.26717
R593 VTAIL.n137 VTAIL.n80 4.26717
R594 VTAIL.n108 VTAIL.n95 4.26717
R595 VTAIL.n250 VTAIL.n234 3.49141
R596 VTAIL.n276 VTAIL.n275 3.49141
R597 VTAIL.n34 VTAIL.n18 3.49141
R598 VTAIL.n60 VTAIL.n59 3.49141
R599 VTAIL.n206 VTAIL.n205 3.49141
R600 VTAIL.n181 VTAIL.n165 3.49141
R601 VTAIL.n134 VTAIL.n133 3.49141
R602 VTAIL.n109 VTAIL.n93 3.49141
R603 VTAIL.n254 VTAIL.n253 2.71565
R604 VTAIL.n272 VTAIL.n224 2.71565
R605 VTAIL.n38 VTAIL.n37 2.71565
R606 VTAIL.n56 VTAIL.n8 2.71565
R607 VTAIL.n202 VTAIL.n154 2.71565
R608 VTAIL.n185 VTAIL.n184 2.71565
R609 VTAIL.n130 VTAIL.n82 2.71565
R610 VTAIL.n113 VTAIL.n112 2.71565
R611 VTAIL.n0 VTAIL.t2 2.53204
R612 VTAIL.n0 VTAIL.t4 2.53204
R613 VTAIL.n72 VTAIL.t7 2.53204
R614 VTAIL.n72 VTAIL.t6 2.53204
R615 VTAIL.n146 VTAIL.t5 2.53204
R616 VTAIL.n146 VTAIL.t10 2.53204
R617 VTAIL.n74 VTAIL.t3 2.53204
R618 VTAIL.n74 VTAIL.t1 2.53204
R619 VTAIL.n243 VTAIL.n239 2.41282
R620 VTAIL.n27 VTAIL.n23 2.41282
R621 VTAIL.n174 VTAIL.n170 2.41282
R622 VTAIL.n102 VTAIL.n98 2.41282
R623 VTAIL.n145 VTAIL.n75 2.05222
R624 VTAIL.n217 VTAIL.n147 2.05222
R625 VTAIL.n73 VTAIL.n71 2.05222
R626 VTAIL.n258 VTAIL.n232 1.93989
R627 VTAIL.n271 VTAIL.n226 1.93989
R628 VTAIL.n42 VTAIL.n16 1.93989
R629 VTAIL.n55 VTAIL.n10 1.93989
R630 VTAIL.n201 VTAIL.n156 1.93989
R631 VTAIL.n188 VTAIL.n162 1.93989
R632 VTAIL.n129 VTAIL.n84 1.93989
R633 VTAIL.n116 VTAIL.n90 1.93989
R634 VTAIL.n147 VTAIL.n145 1.49619
R635 VTAIL.n71 VTAIL.n1 1.49619
R636 VTAIL VTAIL.n287 1.4811
R637 VTAIL.n259 VTAIL.n230 1.16414
R638 VTAIL.n268 VTAIL.n267 1.16414
R639 VTAIL.n43 VTAIL.n14 1.16414
R640 VTAIL.n52 VTAIL.n51 1.16414
R641 VTAIL.n198 VTAIL.n197 1.16414
R642 VTAIL.n189 VTAIL.n160 1.16414
R643 VTAIL.n126 VTAIL.n125 1.16414
R644 VTAIL.n117 VTAIL.n88 1.16414
R645 VTAIL VTAIL.n1 0.571621
R646 VTAIL.n263 VTAIL.n262 0.388379
R647 VTAIL.n264 VTAIL.n228 0.388379
R648 VTAIL.n47 VTAIL.n46 0.388379
R649 VTAIL.n48 VTAIL.n12 0.388379
R650 VTAIL.n194 VTAIL.n158 0.388379
R651 VTAIL.n193 VTAIL.n192 0.388379
R652 VTAIL.n122 VTAIL.n86 0.388379
R653 VTAIL.n121 VTAIL.n120 0.388379
R654 VTAIL.n244 VTAIL.n243 0.155672
R655 VTAIL.n244 VTAIL.n235 0.155672
R656 VTAIL.n251 VTAIL.n235 0.155672
R657 VTAIL.n252 VTAIL.n251 0.155672
R658 VTAIL.n252 VTAIL.n231 0.155672
R659 VTAIL.n260 VTAIL.n231 0.155672
R660 VTAIL.n261 VTAIL.n260 0.155672
R661 VTAIL.n261 VTAIL.n227 0.155672
R662 VTAIL.n269 VTAIL.n227 0.155672
R663 VTAIL.n270 VTAIL.n269 0.155672
R664 VTAIL.n270 VTAIL.n223 0.155672
R665 VTAIL.n277 VTAIL.n223 0.155672
R666 VTAIL.n278 VTAIL.n277 0.155672
R667 VTAIL.n278 VTAIL.n219 0.155672
R668 VTAIL.n285 VTAIL.n219 0.155672
R669 VTAIL.n28 VTAIL.n27 0.155672
R670 VTAIL.n28 VTAIL.n19 0.155672
R671 VTAIL.n35 VTAIL.n19 0.155672
R672 VTAIL.n36 VTAIL.n35 0.155672
R673 VTAIL.n36 VTAIL.n15 0.155672
R674 VTAIL.n44 VTAIL.n15 0.155672
R675 VTAIL.n45 VTAIL.n44 0.155672
R676 VTAIL.n45 VTAIL.n11 0.155672
R677 VTAIL.n53 VTAIL.n11 0.155672
R678 VTAIL.n54 VTAIL.n53 0.155672
R679 VTAIL.n54 VTAIL.n7 0.155672
R680 VTAIL.n61 VTAIL.n7 0.155672
R681 VTAIL.n62 VTAIL.n61 0.155672
R682 VTAIL.n62 VTAIL.n3 0.155672
R683 VTAIL.n69 VTAIL.n3 0.155672
R684 VTAIL.n215 VTAIL.n149 0.155672
R685 VTAIL.n208 VTAIL.n149 0.155672
R686 VTAIL.n208 VTAIL.n207 0.155672
R687 VTAIL.n207 VTAIL.n153 0.155672
R688 VTAIL.n200 VTAIL.n153 0.155672
R689 VTAIL.n200 VTAIL.n199 0.155672
R690 VTAIL.n199 VTAIL.n157 0.155672
R691 VTAIL.n191 VTAIL.n157 0.155672
R692 VTAIL.n191 VTAIL.n190 0.155672
R693 VTAIL.n190 VTAIL.n161 0.155672
R694 VTAIL.n183 VTAIL.n161 0.155672
R695 VTAIL.n183 VTAIL.n182 0.155672
R696 VTAIL.n182 VTAIL.n166 0.155672
R697 VTAIL.n175 VTAIL.n166 0.155672
R698 VTAIL.n175 VTAIL.n174 0.155672
R699 VTAIL.n143 VTAIL.n77 0.155672
R700 VTAIL.n136 VTAIL.n77 0.155672
R701 VTAIL.n136 VTAIL.n135 0.155672
R702 VTAIL.n135 VTAIL.n81 0.155672
R703 VTAIL.n128 VTAIL.n81 0.155672
R704 VTAIL.n128 VTAIL.n127 0.155672
R705 VTAIL.n127 VTAIL.n85 0.155672
R706 VTAIL.n119 VTAIL.n85 0.155672
R707 VTAIL.n119 VTAIL.n118 0.155672
R708 VTAIL.n118 VTAIL.n89 0.155672
R709 VTAIL.n111 VTAIL.n89 0.155672
R710 VTAIL.n111 VTAIL.n110 0.155672
R711 VTAIL.n110 VTAIL.n94 0.155672
R712 VTAIL.n103 VTAIL.n94 0.155672
R713 VTAIL.n103 VTAIL.n102 0.155672
R714 VN.n2 VN.t5 184.941
R715 VN.n14 VN.t0 184.941
R716 VN.n21 VN.n12 161.3
R717 VN.n20 VN.n19 161.3
R718 VN.n18 VN.n13 161.3
R719 VN.n17 VN.n16 161.3
R720 VN.n9 VN.n0 161.3
R721 VN.n8 VN.n7 161.3
R722 VN.n6 VN.n1 161.3
R723 VN.n5 VN.n4 161.3
R724 VN.n3 VN.t1 150.948
R725 VN.n10 VN.t2 150.948
R726 VN.n15 VN.t3 150.948
R727 VN.n22 VN.t4 150.948
R728 VN.n11 VN.n10 92.2184
R729 VN.n23 VN.n22 92.2184
R730 VN.n8 VN.n1 56.5617
R731 VN.n20 VN.n13 56.5617
R732 VN VN.n23 47.4527
R733 VN.n15 VN.n14 46.044
R734 VN.n3 VN.n2 46.044
R735 VN.n4 VN.n3 24.5923
R736 VN.n4 VN.n1 24.5923
R737 VN.n9 VN.n8 24.5923
R738 VN.n16 VN.n13 24.5923
R739 VN.n16 VN.n15 24.5923
R740 VN.n21 VN.n20 24.5923
R741 VN.n10 VN.n9 18.6903
R742 VN.n22 VN.n21 18.6903
R743 VN.n17 VN.n14 9.07974
R744 VN.n5 VN.n2 9.07974
R745 VN.n23 VN.n12 0.278335
R746 VN.n11 VN.n0 0.278335
R747 VN.n19 VN.n12 0.189894
R748 VN.n19 VN.n18 0.189894
R749 VN.n18 VN.n17 0.189894
R750 VN.n6 VN.n5 0.189894
R751 VN.n7 VN.n6 0.189894
R752 VN.n7 VN.n0 0.189894
R753 VN VN.n11 0.153485
R754 VDD2.n135 VDD2.n71 756.745
R755 VDD2.n64 VDD2.n0 756.745
R756 VDD2.n136 VDD2.n135 585
R757 VDD2.n134 VDD2.n133 585
R758 VDD2.n75 VDD2.n74 585
R759 VDD2.n128 VDD2.n127 585
R760 VDD2.n126 VDD2.n125 585
R761 VDD2.n79 VDD2.n78 585
R762 VDD2.n120 VDD2.n119 585
R763 VDD2.n118 VDD2.n117 585
R764 VDD2.n116 VDD2.n82 585
R765 VDD2.n86 VDD2.n83 585
R766 VDD2.n111 VDD2.n110 585
R767 VDD2.n109 VDD2.n108 585
R768 VDD2.n88 VDD2.n87 585
R769 VDD2.n103 VDD2.n102 585
R770 VDD2.n101 VDD2.n100 585
R771 VDD2.n92 VDD2.n91 585
R772 VDD2.n95 VDD2.n94 585
R773 VDD2.n23 VDD2.n22 585
R774 VDD2.n20 VDD2.n19 585
R775 VDD2.n29 VDD2.n28 585
R776 VDD2.n31 VDD2.n30 585
R777 VDD2.n16 VDD2.n15 585
R778 VDD2.n37 VDD2.n36 585
R779 VDD2.n40 VDD2.n39 585
R780 VDD2.n38 VDD2.n12 585
R781 VDD2.n45 VDD2.n11 585
R782 VDD2.n47 VDD2.n46 585
R783 VDD2.n49 VDD2.n48 585
R784 VDD2.n8 VDD2.n7 585
R785 VDD2.n55 VDD2.n54 585
R786 VDD2.n57 VDD2.n56 585
R787 VDD2.n4 VDD2.n3 585
R788 VDD2.n63 VDD2.n62 585
R789 VDD2.n65 VDD2.n64 585
R790 VDD2.t0 VDD2.n21 329.036
R791 VDD2.t1 VDD2.n93 329.036
R792 VDD2.n135 VDD2.n134 171.744
R793 VDD2.n134 VDD2.n74 171.744
R794 VDD2.n127 VDD2.n74 171.744
R795 VDD2.n127 VDD2.n126 171.744
R796 VDD2.n126 VDD2.n78 171.744
R797 VDD2.n119 VDD2.n78 171.744
R798 VDD2.n119 VDD2.n118 171.744
R799 VDD2.n118 VDD2.n82 171.744
R800 VDD2.n86 VDD2.n82 171.744
R801 VDD2.n110 VDD2.n86 171.744
R802 VDD2.n110 VDD2.n109 171.744
R803 VDD2.n109 VDD2.n87 171.744
R804 VDD2.n102 VDD2.n87 171.744
R805 VDD2.n102 VDD2.n101 171.744
R806 VDD2.n101 VDD2.n91 171.744
R807 VDD2.n94 VDD2.n91 171.744
R808 VDD2.n22 VDD2.n19 171.744
R809 VDD2.n29 VDD2.n19 171.744
R810 VDD2.n30 VDD2.n29 171.744
R811 VDD2.n30 VDD2.n15 171.744
R812 VDD2.n37 VDD2.n15 171.744
R813 VDD2.n39 VDD2.n37 171.744
R814 VDD2.n39 VDD2.n38 171.744
R815 VDD2.n38 VDD2.n11 171.744
R816 VDD2.n47 VDD2.n11 171.744
R817 VDD2.n48 VDD2.n47 171.744
R818 VDD2.n48 VDD2.n7 171.744
R819 VDD2.n55 VDD2.n7 171.744
R820 VDD2.n56 VDD2.n55 171.744
R821 VDD2.n56 VDD2.n3 171.744
R822 VDD2.n63 VDD2.n3 171.744
R823 VDD2.n64 VDD2.n63 171.744
R824 VDD2.n94 VDD2.t1 85.8723
R825 VDD2.n22 VDD2.t0 85.8723
R826 VDD2.n70 VDD2.n69 73.469
R827 VDD2 VDD2.n141 73.4659
R828 VDD2.n70 VDD2.n68 50.3476
R829 VDD2.n140 VDD2.n139 48.8641
R830 VDD2.n140 VDD2.n70 41.4524
R831 VDD2.n117 VDD2.n116 13.1884
R832 VDD2.n46 VDD2.n45 13.1884
R833 VDD2.n120 VDD2.n81 12.8005
R834 VDD2.n115 VDD2.n83 12.8005
R835 VDD2.n44 VDD2.n12 12.8005
R836 VDD2.n49 VDD2.n10 12.8005
R837 VDD2.n121 VDD2.n79 12.0247
R838 VDD2.n112 VDD2.n111 12.0247
R839 VDD2.n41 VDD2.n40 12.0247
R840 VDD2.n50 VDD2.n8 12.0247
R841 VDD2.n125 VDD2.n124 11.249
R842 VDD2.n108 VDD2.n85 11.249
R843 VDD2.n36 VDD2.n14 11.249
R844 VDD2.n54 VDD2.n53 11.249
R845 VDD2.n95 VDD2.n93 10.7239
R846 VDD2.n23 VDD2.n21 10.7239
R847 VDD2.n128 VDD2.n77 10.4732
R848 VDD2.n107 VDD2.n88 10.4732
R849 VDD2.n35 VDD2.n16 10.4732
R850 VDD2.n57 VDD2.n6 10.4732
R851 VDD2.n129 VDD2.n75 9.69747
R852 VDD2.n104 VDD2.n103 9.69747
R853 VDD2.n32 VDD2.n31 9.69747
R854 VDD2.n58 VDD2.n4 9.69747
R855 VDD2.n139 VDD2.n138 9.45567
R856 VDD2.n68 VDD2.n67 9.45567
R857 VDD2.n97 VDD2.n96 9.3005
R858 VDD2.n99 VDD2.n98 9.3005
R859 VDD2.n90 VDD2.n89 9.3005
R860 VDD2.n105 VDD2.n104 9.3005
R861 VDD2.n107 VDD2.n106 9.3005
R862 VDD2.n85 VDD2.n84 9.3005
R863 VDD2.n113 VDD2.n112 9.3005
R864 VDD2.n115 VDD2.n114 9.3005
R865 VDD2.n138 VDD2.n137 9.3005
R866 VDD2.n73 VDD2.n72 9.3005
R867 VDD2.n132 VDD2.n131 9.3005
R868 VDD2.n130 VDD2.n129 9.3005
R869 VDD2.n77 VDD2.n76 9.3005
R870 VDD2.n124 VDD2.n123 9.3005
R871 VDD2.n122 VDD2.n121 9.3005
R872 VDD2.n81 VDD2.n80 9.3005
R873 VDD2.n2 VDD2.n1 9.3005
R874 VDD2.n61 VDD2.n60 9.3005
R875 VDD2.n59 VDD2.n58 9.3005
R876 VDD2.n6 VDD2.n5 9.3005
R877 VDD2.n53 VDD2.n52 9.3005
R878 VDD2.n51 VDD2.n50 9.3005
R879 VDD2.n10 VDD2.n9 9.3005
R880 VDD2.n25 VDD2.n24 9.3005
R881 VDD2.n27 VDD2.n26 9.3005
R882 VDD2.n18 VDD2.n17 9.3005
R883 VDD2.n33 VDD2.n32 9.3005
R884 VDD2.n35 VDD2.n34 9.3005
R885 VDD2.n14 VDD2.n13 9.3005
R886 VDD2.n42 VDD2.n41 9.3005
R887 VDD2.n44 VDD2.n43 9.3005
R888 VDD2.n67 VDD2.n66 9.3005
R889 VDD2.n133 VDD2.n132 8.92171
R890 VDD2.n100 VDD2.n90 8.92171
R891 VDD2.n28 VDD2.n18 8.92171
R892 VDD2.n62 VDD2.n61 8.92171
R893 VDD2.n136 VDD2.n73 8.14595
R894 VDD2.n99 VDD2.n92 8.14595
R895 VDD2.n27 VDD2.n20 8.14595
R896 VDD2.n65 VDD2.n2 8.14595
R897 VDD2.n137 VDD2.n71 7.3702
R898 VDD2.n96 VDD2.n95 7.3702
R899 VDD2.n24 VDD2.n23 7.3702
R900 VDD2.n66 VDD2.n0 7.3702
R901 VDD2.n139 VDD2.n71 6.59444
R902 VDD2.n68 VDD2.n0 6.59444
R903 VDD2.n137 VDD2.n136 5.81868
R904 VDD2.n96 VDD2.n92 5.81868
R905 VDD2.n24 VDD2.n20 5.81868
R906 VDD2.n66 VDD2.n65 5.81868
R907 VDD2.n133 VDD2.n73 5.04292
R908 VDD2.n100 VDD2.n99 5.04292
R909 VDD2.n28 VDD2.n27 5.04292
R910 VDD2.n62 VDD2.n2 5.04292
R911 VDD2.n132 VDD2.n75 4.26717
R912 VDD2.n103 VDD2.n90 4.26717
R913 VDD2.n31 VDD2.n18 4.26717
R914 VDD2.n61 VDD2.n4 4.26717
R915 VDD2.n129 VDD2.n128 3.49141
R916 VDD2.n104 VDD2.n88 3.49141
R917 VDD2.n32 VDD2.n16 3.49141
R918 VDD2.n58 VDD2.n57 3.49141
R919 VDD2.n125 VDD2.n77 2.71565
R920 VDD2.n108 VDD2.n107 2.71565
R921 VDD2.n36 VDD2.n35 2.71565
R922 VDD2.n54 VDD2.n6 2.71565
R923 VDD2.n141 VDD2.t2 2.53204
R924 VDD2.n141 VDD2.t5 2.53204
R925 VDD2.n69 VDD2.t4 2.53204
R926 VDD2.n69 VDD2.t3 2.53204
R927 VDD2.n97 VDD2.n93 2.41282
R928 VDD2.n25 VDD2.n21 2.41282
R929 VDD2.n124 VDD2.n79 1.93989
R930 VDD2.n111 VDD2.n85 1.93989
R931 VDD2.n40 VDD2.n14 1.93989
R932 VDD2.n53 VDD2.n8 1.93989
R933 VDD2 VDD2.n140 1.59748
R934 VDD2.n121 VDD2.n120 1.16414
R935 VDD2.n112 VDD2.n83 1.16414
R936 VDD2.n41 VDD2.n12 1.16414
R937 VDD2.n50 VDD2.n49 1.16414
R938 VDD2.n117 VDD2.n81 0.388379
R939 VDD2.n116 VDD2.n115 0.388379
R940 VDD2.n45 VDD2.n44 0.388379
R941 VDD2.n46 VDD2.n10 0.388379
R942 VDD2.n138 VDD2.n72 0.155672
R943 VDD2.n131 VDD2.n72 0.155672
R944 VDD2.n131 VDD2.n130 0.155672
R945 VDD2.n130 VDD2.n76 0.155672
R946 VDD2.n123 VDD2.n76 0.155672
R947 VDD2.n123 VDD2.n122 0.155672
R948 VDD2.n122 VDD2.n80 0.155672
R949 VDD2.n114 VDD2.n80 0.155672
R950 VDD2.n114 VDD2.n113 0.155672
R951 VDD2.n113 VDD2.n84 0.155672
R952 VDD2.n106 VDD2.n84 0.155672
R953 VDD2.n106 VDD2.n105 0.155672
R954 VDD2.n105 VDD2.n89 0.155672
R955 VDD2.n98 VDD2.n89 0.155672
R956 VDD2.n98 VDD2.n97 0.155672
R957 VDD2.n26 VDD2.n25 0.155672
R958 VDD2.n26 VDD2.n17 0.155672
R959 VDD2.n33 VDD2.n17 0.155672
R960 VDD2.n34 VDD2.n33 0.155672
R961 VDD2.n34 VDD2.n13 0.155672
R962 VDD2.n42 VDD2.n13 0.155672
R963 VDD2.n43 VDD2.n42 0.155672
R964 VDD2.n43 VDD2.n9 0.155672
R965 VDD2.n51 VDD2.n9 0.155672
R966 VDD2.n52 VDD2.n51 0.155672
R967 VDD2.n52 VDD2.n5 0.155672
R968 VDD2.n59 VDD2.n5 0.155672
R969 VDD2.n60 VDD2.n59 0.155672
R970 VDD2.n60 VDD2.n1 0.155672
R971 VDD2.n67 VDD2.n1 0.155672
R972 B.n492 B.n73 585
R973 B.n494 B.n493 585
R974 B.n495 B.n72 585
R975 B.n497 B.n496 585
R976 B.n498 B.n71 585
R977 B.n500 B.n499 585
R978 B.n501 B.n70 585
R979 B.n503 B.n502 585
R980 B.n504 B.n69 585
R981 B.n506 B.n505 585
R982 B.n507 B.n68 585
R983 B.n509 B.n508 585
R984 B.n510 B.n67 585
R985 B.n512 B.n511 585
R986 B.n513 B.n66 585
R987 B.n515 B.n514 585
R988 B.n516 B.n65 585
R989 B.n518 B.n517 585
R990 B.n519 B.n64 585
R991 B.n521 B.n520 585
R992 B.n522 B.n63 585
R993 B.n524 B.n523 585
R994 B.n525 B.n62 585
R995 B.n527 B.n526 585
R996 B.n528 B.n61 585
R997 B.n530 B.n529 585
R998 B.n531 B.n60 585
R999 B.n533 B.n532 585
R1000 B.n534 B.n59 585
R1001 B.n536 B.n535 585
R1002 B.n537 B.n58 585
R1003 B.n539 B.n538 585
R1004 B.n540 B.n57 585
R1005 B.n542 B.n541 585
R1006 B.n543 B.n56 585
R1007 B.n545 B.n544 585
R1008 B.n546 B.n55 585
R1009 B.n548 B.n547 585
R1010 B.n549 B.n54 585
R1011 B.n551 B.n550 585
R1012 B.n552 B.n53 585
R1013 B.n554 B.n553 585
R1014 B.n555 B.n52 585
R1015 B.n557 B.n556 585
R1016 B.n559 B.n49 585
R1017 B.n561 B.n560 585
R1018 B.n562 B.n48 585
R1019 B.n564 B.n563 585
R1020 B.n565 B.n47 585
R1021 B.n567 B.n566 585
R1022 B.n568 B.n46 585
R1023 B.n570 B.n569 585
R1024 B.n571 B.n45 585
R1025 B.n573 B.n572 585
R1026 B.n575 B.n574 585
R1027 B.n576 B.n41 585
R1028 B.n578 B.n577 585
R1029 B.n579 B.n40 585
R1030 B.n581 B.n580 585
R1031 B.n582 B.n39 585
R1032 B.n584 B.n583 585
R1033 B.n585 B.n38 585
R1034 B.n587 B.n586 585
R1035 B.n588 B.n37 585
R1036 B.n590 B.n589 585
R1037 B.n591 B.n36 585
R1038 B.n593 B.n592 585
R1039 B.n594 B.n35 585
R1040 B.n596 B.n595 585
R1041 B.n597 B.n34 585
R1042 B.n599 B.n598 585
R1043 B.n600 B.n33 585
R1044 B.n602 B.n601 585
R1045 B.n603 B.n32 585
R1046 B.n605 B.n604 585
R1047 B.n606 B.n31 585
R1048 B.n608 B.n607 585
R1049 B.n609 B.n30 585
R1050 B.n611 B.n610 585
R1051 B.n612 B.n29 585
R1052 B.n614 B.n613 585
R1053 B.n615 B.n28 585
R1054 B.n617 B.n616 585
R1055 B.n618 B.n27 585
R1056 B.n620 B.n619 585
R1057 B.n621 B.n26 585
R1058 B.n623 B.n622 585
R1059 B.n624 B.n25 585
R1060 B.n626 B.n625 585
R1061 B.n627 B.n24 585
R1062 B.n629 B.n628 585
R1063 B.n630 B.n23 585
R1064 B.n632 B.n631 585
R1065 B.n633 B.n22 585
R1066 B.n635 B.n634 585
R1067 B.n636 B.n21 585
R1068 B.n638 B.n637 585
R1069 B.n639 B.n20 585
R1070 B.n491 B.n490 585
R1071 B.n489 B.n74 585
R1072 B.n488 B.n487 585
R1073 B.n486 B.n75 585
R1074 B.n485 B.n484 585
R1075 B.n483 B.n76 585
R1076 B.n482 B.n481 585
R1077 B.n480 B.n77 585
R1078 B.n479 B.n478 585
R1079 B.n477 B.n78 585
R1080 B.n476 B.n475 585
R1081 B.n474 B.n79 585
R1082 B.n473 B.n472 585
R1083 B.n471 B.n80 585
R1084 B.n470 B.n469 585
R1085 B.n468 B.n81 585
R1086 B.n467 B.n466 585
R1087 B.n465 B.n82 585
R1088 B.n464 B.n463 585
R1089 B.n462 B.n83 585
R1090 B.n461 B.n460 585
R1091 B.n459 B.n84 585
R1092 B.n458 B.n457 585
R1093 B.n456 B.n85 585
R1094 B.n455 B.n454 585
R1095 B.n453 B.n86 585
R1096 B.n452 B.n451 585
R1097 B.n450 B.n87 585
R1098 B.n449 B.n448 585
R1099 B.n447 B.n88 585
R1100 B.n446 B.n445 585
R1101 B.n444 B.n89 585
R1102 B.n443 B.n442 585
R1103 B.n441 B.n90 585
R1104 B.n440 B.n439 585
R1105 B.n438 B.n91 585
R1106 B.n437 B.n436 585
R1107 B.n435 B.n92 585
R1108 B.n434 B.n433 585
R1109 B.n432 B.n93 585
R1110 B.n431 B.n430 585
R1111 B.n429 B.n94 585
R1112 B.n428 B.n427 585
R1113 B.n426 B.n95 585
R1114 B.n425 B.n424 585
R1115 B.n423 B.n96 585
R1116 B.n422 B.n421 585
R1117 B.n420 B.n97 585
R1118 B.n419 B.n418 585
R1119 B.n417 B.n98 585
R1120 B.n416 B.n415 585
R1121 B.n414 B.n99 585
R1122 B.n413 B.n412 585
R1123 B.n411 B.n100 585
R1124 B.n410 B.n409 585
R1125 B.n408 B.n101 585
R1126 B.n407 B.n406 585
R1127 B.n405 B.n102 585
R1128 B.n404 B.n403 585
R1129 B.n402 B.n103 585
R1130 B.n401 B.n400 585
R1131 B.n399 B.n104 585
R1132 B.n398 B.n397 585
R1133 B.n396 B.n105 585
R1134 B.n395 B.n394 585
R1135 B.n393 B.n106 585
R1136 B.n392 B.n391 585
R1137 B.n390 B.n107 585
R1138 B.n389 B.n388 585
R1139 B.n387 B.n108 585
R1140 B.n386 B.n385 585
R1141 B.n384 B.n109 585
R1142 B.n383 B.n382 585
R1143 B.n234 B.n163 585
R1144 B.n236 B.n235 585
R1145 B.n237 B.n162 585
R1146 B.n239 B.n238 585
R1147 B.n240 B.n161 585
R1148 B.n242 B.n241 585
R1149 B.n243 B.n160 585
R1150 B.n245 B.n244 585
R1151 B.n246 B.n159 585
R1152 B.n248 B.n247 585
R1153 B.n249 B.n158 585
R1154 B.n251 B.n250 585
R1155 B.n252 B.n157 585
R1156 B.n254 B.n253 585
R1157 B.n255 B.n156 585
R1158 B.n257 B.n256 585
R1159 B.n258 B.n155 585
R1160 B.n260 B.n259 585
R1161 B.n261 B.n154 585
R1162 B.n263 B.n262 585
R1163 B.n264 B.n153 585
R1164 B.n266 B.n265 585
R1165 B.n267 B.n152 585
R1166 B.n269 B.n268 585
R1167 B.n270 B.n151 585
R1168 B.n272 B.n271 585
R1169 B.n273 B.n150 585
R1170 B.n275 B.n274 585
R1171 B.n276 B.n149 585
R1172 B.n278 B.n277 585
R1173 B.n279 B.n148 585
R1174 B.n281 B.n280 585
R1175 B.n282 B.n147 585
R1176 B.n284 B.n283 585
R1177 B.n285 B.n146 585
R1178 B.n287 B.n286 585
R1179 B.n288 B.n145 585
R1180 B.n290 B.n289 585
R1181 B.n291 B.n144 585
R1182 B.n293 B.n292 585
R1183 B.n294 B.n143 585
R1184 B.n296 B.n295 585
R1185 B.n297 B.n142 585
R1186 B.n299 B.n298 585
R1187 B.n301 B.n139 585
R1188 B.n303 B.n302 585
R1189 B.n304 B.n138 585
R1190 B.n306 B.n305 585
R1191 B.n307 B.n137 585
R1192 B.n309 B.n308 585
R1193 B.n310 B.n136 585
R1194 B.n312 B.n311 585
R1195 B.n313 B.n135 585
R1196 B.n315 B.n314 585
R1197 B.n317 B.n316 585
R1198 B.n318 B.n131 585
R1199 B.n320 B.n319 585
R1200 B.n321 B.n130 585
R1201 B.n323 B.n322 585
R1202 B.n324 B.n129 585
R1203 B.n326 B.n325 585
R1204 B.n327 B.n128 585
R1205 B.n329 B.n328 585
R1206 B.n330 B.n127 585
R1207 B.n332 B.n331 585
R1208 B.n333 B.n126 585
R1209 B.n335 B.n334 585
R1210 B.n336 B.n125 585
R1211 B.n338 B.n337 585
R1212 B.n339 B.n124 585
R1213 B.n341 B.n340 585
R1214 B.n342 B.n123 585
R1215 B.n344 B.n343 585
R1216 B.n345 B.n122 585
R1217 B.n347 B.n346 585
R1218 B.n348 B.n121 585
R1219 B.n350 B.n349 585
R1220 B.n351 B.n120 585
R1221 B.n353 B.n352 585
R1222 B.n354 B.n119 585
R1223 B.n356 B.n355 585
R1224 B.n357 B.n118 585
R1225 B.n359 B.n358 585
R1226 B.n360 B.n117 585
R1227 B.n362 B.n361 585
R1228 B.n363 B.n116 585
R1229 B.n365 B.n364 585
R1230 B.n366 B.n115 585
R1231 B.n368 B.n367 585
R1232 B.n369 B.n114 585
R1233 B.n371 B.n370 585
R1234 B.n372 B.n113 585
R1235 B.n374 B.n373 585
R1236 B.n375 B.n112 585
R1237 B.n377 B.n376 585
R1238 B.n378 B.n111 585
R1239 B.n380 B.n379 585
R1240 B.n381 B.n110 585
R1241 B.n233 B.n232 585
R1242 B.n231 B.n164 585
R1243 B.n230 B.n229 585
R1244 B.n228 B.n165 585
R1245 B.n227 B.n226 585
R1246 B.n225 B.n166 585
R1247 B.n224 B.n223 585
R1248 B.n222 B.n167 585
R1249 B.n221 B.n220 585
R1250 B.n219 B.n168 585
R1251 B.n218 B.n217 585
R1252 B.n216 B.n169 585
R1253 B.n215 B.n214 585
R1254 B.n213 B.n170 585
R1255 B.n212 B.n211 585
R1256 B.n210 B.n171 585
R1257 B.n209 B.n208 585
R1258 B.n207 B.n172 585
R1259 B.n206 B.n205 585
R1260 B.n204 B.n173 585
R1261 B.n203 B.n202 585
R1262 B.n201 B.n174 585
R1263 B.n200 B.n199 585
R1264 B.n198 B.n175 585
R1265 B.n197 B.n196 585
R1266 B.n195 B.n176 585
R1267 B.n194 B.n193 585
R1268 B.n192 B.n177 585
R1269 B.n191 B.n190 585
R1270 B.n189 B.n178 585
R1271 B.n188 B.n187 585
R1272 B.n186 B.n179 585
R1273 B.n185 B.n184 585
R1274 B.n183 B.n180 585
R1275 B.n182 B.n181 585
R1276 B.n2 B.n0 585
R1277 B.n693 B.n1 585
R1278 B.n692 B.n691 585
R1279 B.n690 B.n3 585
R1280 B.n689 B.n688 585
R1281 B.n687 B.n4 585
R1282 B.n686 B.n685 585
R1283 B.n684 B.n5 585
R1284 B.n683 B.n682 585
R1285 B.n681 B.n6 585
R1286 B.n680 B.n679 585
R1287 B.n678 B.n7 585
R1288 B.n677 B.n676 585
R1289 B.n675 B.n8 585
R1290 B.n674 B.n673 585
R1291 B.n672 B.n9 585
R1292 B.n671 B.n670 585
R1293 B.n669 B.n10 585
R1294 B.n668 B.n667 585
R1295 B.n666 B.n11 585
R1296 B.n665 B.n664 585
R1297 B.n663 B.n12 585
R1298 B.n662 B.n661 585
R1299 B.n660 B.n13 585
R1300 B.n659 B.n658 585
R1301 B.n657 B.n14 585
R1302 B.n656 B.n655 585
R1303 B.n654 B.n15 585
R1304 B.n653 B.n652 585
R1305 B.n651 B.n16 585
R1306 B.n650 B.n649 585
R1307 B.n648 B.n17 585
R1308 B.n647 B.n646 585
R1309 B.n645 B.n18 585
R1310 B.n644 B.n643 585
R1311 B.n642 B.n19 585
R1312 B.n641 B.n640 585
R1313 B.n695 B.n694 585
R1314 B.n232 B.n163 497.305
R1315 B.n640 B.n639 497.305
R1316 B.n382 B.n381 497.305
R1317 B.n490 B.n73 497.305
R1318 B.n132 B.t2 437.038
R1319 B.n50 B.t10 437.038
R1320 B.n140 B.t8 437.038
R1321 B.n42 B.t4 437.038
R1322 B.n133 B.t1 390.88
R1323 B.n51 B.t11 390.88
R1324 B.n141 B.t7 390.88
R1325 B.n43 B.t5 390.88
R1326 B.n132 B.t0 357.981
R1327 B.n140 B.t6 357.981
R1328 B.n42 B.t3 357.981
R1329 B.n50 B.t9 357.981
R1330 B.n232 B.n231 163.367
R1331 B.n231 B.n230 163.367
R1332 B.n230 B.n165 163.367
R1333 B.n226 B.n165 163.367
R1334 B.n226 B.n225 163.367
R1335 B.n225 B.n224 163.367
R1336 B.n224 B.n167 163.367
R1337 B.n220 B.n167 163.367
R1338 B.n220 B.n219 163.367
R1339 B.n219 B.n218 163.367
R1340 B.n218 B.n169 163.367
R1341 B.n214 B.n169 163.367
R1342 B.n214 B.n213 163.367
R1343 B.n213 B.n212 163.367
R1344 B.n212 B.n171 163.367
R1345 B.n208 B.n171 163.367
R1346 B.n208 B.n207 163.367
R1347 B.n207 B.n206 163.367
R1348 B.n206 B.n173 163.367
R1349 B.n202 B.n173 163.367
R1350 B.n202 B.n201 163.367
R1351 B.n201 B.n200 163.367
R1352 B.n200 B.n175 163.367
R1353 B.n196 B.n175 163.367
R1354 B.n196 B.n195 163.367
R1355 B.n195 B.n194 163.367
R1356 B.n194 B.n177 163.367
R1357 B.n190 B.n177 163.367
R1358 B.n190 B.n189 163.367
R1359 B.n189 B.n188 163.367
R1360 B.n188 B.n179 163.367
R1361 B.n184 B.n179 163.367
R1362 B.n184 B.n183 163.367
R1363 B.n183 B.n182 163.367
R1364 B.n182 B.n2 163.367
R1365 B.n694 B.n2 163.367
R1366 B.n694 B.n693 163.367
R1367 B.n693 B.n692 163.367
R1368 B.n692 B.n3 163.367
R1369 B.n688 B.n3 163.367
R1370 B.n688 B.n687 163.367
R1371 B.n687 B.n686 163.367
R1372 B.n686 B.n5 163.367
R1373 B.n682 B.n5 163.367
R1374 B.n682 B.n681 163.367
R1375 B.n681 B.n680 163.367
R1376 B.n680 B.n7 163.367
R1377 B.n676 B.n7 163.367
R1378 B.n676 B.n675 163.367
R1379 B.n675 B.n674 163.367
R1380 B.n674 B.n9 163.367
R1381 B.n670 B.n9 163.367
R1382 B.n670 B.n669 163.367
R1383 B.n669 B.n668 163.367
R1384 B.n668 B.n11 163.367
R1385 B.n664 B.n11 163.367
R1386 B.n664 B.n663 163.367
R1387 B.n663 B.n662 163.367
R1388 B.n662 B.n13 163.367
R1389 B.n658 B.n13 163.367
R1390 B.n658 B.n657 163.367
R1391 B.n657 B.n656 163.367
R1392 B.n656 B.n15 163.367
R1393 B.n652 B.n15 163.367
R1394 B.n652 B.n651 163.367
R1395 B.n651 B.n650 163.367
R1396 B.n650 B.n17 163.367
R1397 B.n646 B.n17 163.367
R1398 B.n646 B.n645 163.367
R1399 B.n645 B.n644 163.367
R1400 B.n644 B.n19 163.367
R1401 B.n640 B.n19 163.367
R1402 B.n236 B.n163 163.367
R1403 B.n237 B.n236 163.367
R1404 B.n238 B.n237 163.367
R1405 B.n238 B.n161 163.367
R1406 B.n242 B.n161 163.367
R1407 B.n243 B.n242 163.367
R1408 B.n244 B.n243 163.367
R1409 B.n244 B.n159 163.367
R1410 B.n248 B.n159 163.367
R1411 B.n249 B.n248 163.367
R1412 B.n250 B.n249 163.367
R1413 B.n250 B.n157 163.367
R1414 B.n254 B.n157 163.367
R1415 B.n255 B.n254 163.367
R1416 B.n256 B.n255 163.367
R1417 B.n256 B.n155 163.367
R1418 B.n260 B.n155 163.367
R1419 B.n261 B.n260 163.367
R1420 B.n262 B.n261 163.367
R1421 B.n262 B.n153 163.367
R1422 B.n266 B.n153 163.367
R1423 B.n267 B.n266 163.367
R1424 B.n268 B.n267 163.367
R1425 B.n268 B.n151 163.367
R1426 B.n272 B.n151 163.367
R1427 B.n273 B.n272 163.367
R1428 B.n274 B.n273 163.367
R1429 B.n274 B.n149 163.367
R1430 B.n278 B.n149 163.367
R1431 B.n279 B.n278 163.367
R1432 B.n280 B.n279 163.367
R1433 B.n280 B.n147 163.367
R1434 B.n284 B.n147 163.367
R1435 B.n285 B.n284 163.367
R1436 B.n286 B.n285 163.367
R1437 B.n286 B.n145 163.367
R1438 B.n290 B.n145 163.367
R1439 B.n291 B.n290 163.367
R1440 B.n292 B.n291 163.367
R1441 B.n292 B.n143 163.367
R1442 B.n296 B.n143 163.367
R1443 B.n297 B.n296 163.367
R1444 B.n298 B.n297 163.367
R1445 B.n298 B.n139 163.367
R1446 B.n303 B.n139 163.367
R1447 B.n304 B.n303 163.367
R1448 B.n305 B.n304 163.367
R1449 B.n305 B.n137 163.367
R1450 B.n309 B.n137 163.367
R1451 B.n310 B.n309 163.367
R1452 B.n311 B.n310 163.367
R1453 B.n311 B.n135 163.367
R1454 B.n315 B.n135 163.367
R1455 B.n316 B.n315 163.367
R1456 B.n316 B.n131 163.367
R1457 B.n320 B.n131 163.367
R1458 B.n321 B.n320 163.367
R1459 B.n322 B.n321 163.367
R1460 B.n322 B.n129 163.367
R1461 B.n326 B.n129 163.367
R1462 B.n327 B.n326 163.367
R1463 B.n328 B.n327 163.367
R1464 B.n328 B.n127 163.367
R1465 B.n332 B.n127 163.367
R1466 B.n333 B.n332 163.367
R1467 B.n334 B.n333 163.367
R1468 B.n334 B.n125 163.367
R1469 B.n338 B.n125 163.367
R1470 B.n339 B.n338 163.367
R1471 B.n340 B.n339 163.367
R1472 B.n340 B.n123 163.367
R1473 B.n344 B.n123 163.367
R1474 B.n345 B.n344 163.367
R1475 B.n346 B.n345 163.367
R1476 B.n346 B.n121 163.367
R1477 B.n350 B.n121 163.367
R1478 B.n351 B.n350 163.367
R1479 B.n352 B.n351 163.367
R1480 B.n352 B.n119 163.367
R1481 B.n356 B.n119 163.367
R1482 B.n357 B.n356 163.367
R1483 B.n358 B.n357 163.367
R1484 B.n358 B.n117 163.367
R1485 B.n362 B.n117 163.367
R1486 B.n363 B.n362 163.367
R1487 B.n364 B.n363 163.367
R1488 B.n364 B.n115 163.367
R1489 B.n368 B.n115 163.367
R1490 B.n369 B.n368 163.367
R1491 B.n370 B.n369 163.367
R1492 B.n370 B.n113 163.367
R1493 B.n374 B.n113 163.367
R1494 B.n375 B.n374 163.367
R1495 B.n376 B.n375 163.367
R1496 B.n376 B.n111 163.367
R1497 B.n380 B.n111 163.367
R1498 B.n381 B.n380 163.367
R1499 B.n382 B.n109 163.367
R1500 B.n386 B.n109 163.367
R1501 B.n387 B.n386 163.367
R1502 B.n388 B.n387 163.367
R1503 B.n388 B.n107 163.367
R1504 B.n392 B.n107 163.367
R1505 B.n393 B.n392 163.367
R1506 B.n394 B.n393 163.367
R1507 B.n394 B.n105 163.367
R1508 B.n398 B.n105 163.367
R1509 B.n399 B.n398 163.367
R1510 B.n400 B.n399 163.367
R1511 B.n400 B.n103 163.367
R1512 B.n404 B.n103 163.367
R1513 B.n405 B.n404 163.367
R1514 B.n406 B.n405 163.367
R1515 B.n406 B.n101 163.367
R1516 B.n410 B.n101 163.367
R1517 B.n411 B.n410 163.367
R1518 B.n412 B.n411 163.367
R1519 B.n412 B.n99 163.367
R1520 B.n416 B.n99 163.367
R1521 B.n417 B.n416 163.367
R1522 B.n418 B.n417 163.367
R1523 B.n418 B.n97 163.367
R1524 B.n422 B.n97 163.367
R1525 B.n423 B.n422 163.367
R1526 B.n424 B.n423 163.367
R1527 B.n424 B.n95 163.367
R1528 B.n428 B.n95 163.367
R1529 B.n429 B.n428 163.367
R1530 B.n430 B.n429 163.367
R1531 B.n430 B.n93 163.367
R1532 B.n434 B.n93 163.367
R1533 B.n435 B.n434 163.367
R1534 B.n436 B.n435 163.367
R1535 B.n436 B.n91 163.367
R1536 B.n440 B.n91 163.367
R1537 B.n441 B.n440 163.367
R1538 B.n442 B.n441 163.367
R1539 B.n442 B.n89 163.367
R1540 B.n446 B.n89 163.367
R1541 B.n447 B.n446 163.367
R1542 B.n448 B.n447 163.367
R1543 B.n448 B.n87 163.367
R1544 B.n452 B.n87 163.367
R1545 B.n453 B.n452 163.367
R1546 B.n454 B.n453 163.367
R1547 B.n454 B.n85 163.367
R1548 B.n458 B.n85 163.367
R1549 B.n459 B.n458 163.367
R1550 B.n460 B.n459 163.367
R1551 B.n460 B.n83 163.367
R1552 B.n464 B.n83 163.367
R1553 B.n465 B.n464 163.367
R1554 B.n466 B.n465 163.367
R1555 B.n466 B.n81 163.367
R1556 B.n470 B.n81 163.367
R1557 B.n471 B.n470 163.367
R1558 B.n472 B.n471 163.367
R1559 B.n472 B.n79 163.367
R1560 B.n476 B.n79 163.367
R1561 B.n477 B.n476 163.367
R1562 B.n478 B.n477 163.367
R1563 B.n478 B.n77 163.367
R1564 B.n482 B.n77 163.367
R1565 B.n483 B.n482 163.367
R1566 B.n484 B.n483 163.367
R1567 B.n484 B.n75 163.367
R1568 B.n488 B.n75 163.367
R1569 B.n489 B.n488 163.367
R1570 B.n490 B.n489 163.367
R1571 B.n639 B.n638 163.367
R1572 B.n638 B.n21 163.367
R1573 B.n634 B.n21 163.367
R1574 B.n634 B.n633 163.367
R1575 B.n633 B.n632 163.367
R1576 B.n632 B.n23 163.367
R1577 B.n628 B.n23 163.367
R1578 B.n628 B.n627 163.367
R1579 B.n627 B.n626 163.367
R1580 B.n626 B.n25 163.367
R1581 B.n622 B.n25 163.367
R1582 B.n622 B.n621 163.367
R1583 B.n621 B.n620 163.367
R1584 B.n620 B.n27 163.367
R1585 B.n616 B.n27 163.367
R1586 B.n616 B.n615 163.367
R1587 B.n615 B.n614 163.367
R1588 B.n614 B.n29 163.367
R1589 B.n610 B.n29 163.367
R1590 B.n610 B.n609 163.367
R1591 B.n609 B.n608 163.367
R1592 B.n608 B.n31 163.367
R1593 B.n604 B.n31 163.367
R1594 B.n604 B.n603 163.367
R1595 B.n603 B.n602 163.367
R1596 B.n602 B.n33 163.367
R1597 B.n598 B.n33 163.367
R1598 B.n598 B.n597 163.367
R1599 B.n597 B.n596 163.367
R1600 B.n596 B.n35 163.367
R1601 B.n592 B.n35 163.367
R1602 B.n592 B.n591 163.367
R1603 B.n591 B.n590 163.367
R1604 B.n590 B.n37 163.367
R1605 B.n586 B.n37 163.367
R1606 B.n586 B.n585 163.367
R1607 B.n585 B.n584 163.367
R1608 B.n584 B.n39 163.367
R1609 B.n580 B.n39 163.367
R1610 B.n580 B.n579 163.367
R1611 B.n579 B.n578 163.367
R1612 B.n578 B.n41 163.367
R1613 B.n574 B.n41 163.367
R1614 B.n574 B.n573 163.367
R1615 B.n573 B.n45 163.367
R1616 B.n569 B.n45 163.367
R1617 B.n569 B.n568 163.367
R1618 B.n568 B.n567 163.367
R1619 B.n567 B.n47 163.367
R1620 B.n563 B.n47 163.367
R1621 B.n563 B.n562 163.367
R1622 B.n562 B.n561 163.367
R1623 B.n561 B.n49 163.367
R1624 B.n556 B.n49 163.367
R1625 B.n556 B.n555 163.367
R1626 B.n555 B.n554 163.367
R1627 B.n554 B.n53 163.367
R1628 B.n550 B.n53 163.367
R1629 B.n550 B.n549 163.367
R1630 B.n549 B.n548 163.367
R1631 B.n548 B.n55 163.367
R1632 B.n544 B.n55 163.367
R1633 B.n544 B.n543 163.367
R1634 B.n543 B.n542 163.367
R1635 B.n542 B.n57 163.367
R1636 B.n538 B.n57 163.367
R1637 B.n538 B.n537 163.367
R1638 B.n537 B.n536 163.367
R1639 B.n536 B.n59 163.367
R1640 B.n532 B.n59 163.367
R1641 B.n532 B.n531 163.367
R1642 B.n531 B.n530 163.367
R1643 B.n530 B.n61 163.367
R1644 B.n526 B.n61 163.367
R1645 B.n526 B.n525 163.367
R1646 B.n525 B.n524 163.367
R1647 B.n524 B.n63 163.367
R1648 B.n520 B.n63 163.367
R1649 B.n520 B.n519 163.367
R1650 B.n519 B.n518 163.367
R1651 B.n518 B.n65 163.367
R1652 B.n514 B.n65 163.367
R1653 B.n514 B.n513 163.367
R1654 B.n513 B.n512 163.367
R1655 B.n512 B.n67 163.367
R1656 B.n508 B.n67 163.367
R1657 B.n508 B.n507 163.367
R1658 B.n507 B.n506 163.367
R1659 B.n506 B.n69 163.367
R1660 B.n502 B.n69 163.367
R1661 B.n502 B.n501 163.367
R1662 B.n501 B.n500 163.367
R1663 B.n500 B.n71 163.367
R1664 B.n496 B.n71 163.367
R1665 B.n496 B.n495 163.367
R1666 B.n495 B.n494 163.367
R1667 B.n494 B.n73 163.367
R1668 B.n134 B.n133 59.5399
R1669 B.n300 B.n141 59.5399
R1670 B.n44 B.n43 59.5399
R1671 B.n558 B.n51 59.5399
R1672 B.n133 B.n132 46.1581
R1673 B.n141 B.n140 46.1581
R1674 B.n43 B.n42 46.1581
R1675 B.n51 B.n50 46.1581
R1676 B.n641 B.n20 32.3127
R1677 B.n492 B.n491 32.3127
R1678 B.n383 B.n110 32.3127
R1679 B.n234 B.n233 32.3127
R1680 B B.n695 18.0485
R1681 B.n637 B.n20 10.6151
R1682 B.n637 B.n636 10.6151
R1683 B.n636 B.n635 10.6151
R1684 B.n635 B.n22 10.6151
R1685 B.n631 B.n22 10.6151
R1686 B.n631 B.n630 10.6151
R1687 B.n630 B.n629 10.6151
R1688 B.n629 B.n24 10.6151
R1689 B.n625 B.n24 10.6151
R1690 B.n625 B.n624 10.6151
R1691 B.n624 B.n623 10.6151
R1692 B.n623 B.n26 10.6151
R1693 B.n619 B.n26 10.6151
R1694 B.n619 B.n618 10.6151
R1695 B.n618 B.n617 10.6151
R1696 B.n617 B.n28 10.6151
R1697 B.n613 B.n28 10.6151
R1698 B.n613 B.n612 10.6151
R1699 B.n612 B.n611 10.6151
R1700 B.n611 B.n30 10.6151
R1701 B.n607 B.n30 10.6151
R1702 B.n607 B.n606 10.6151
R1703 B.n606 B.n605 10.6151
R1704 B.n605 B.n32 10.6151
R1705 B.n601 B.n32 10.6151
R1706 B.n601 B.n600 10.6151
R1707 B.n600 B.n599 10.6151
R1708 B.n599 B.n34 10.6151
R1709 B.n595 B.n34 10.6151
R1710 B.n595 B.n594 10.6151
R1711 B.n594 B.n593 10.6151
R1712 B.n593 B.n36 10.6151
R1713 B.n589 B.n36 10.6151
R1714 B.n589 B.n588 10.6151
R1715 B.n588 B.n587 10.6151
R1716 B.n587 B.n38 10.6151
R1717 B.n583 B.n38 10.6151
R1718 B.n583 B.n582 10.6151
R1719 B.n582 B.n581 10.6151
R1720 B.n581 B.n40 10.6151
R1721 B.n577 B.n40 10.6151
R1722 B.n577 B.n576 10.6151
R1723 B.n576 B.n575 10.6151
R1724 B.n572 B.n571 10.6151
R1725 B.n571 B.n570 10.6151
R1726 B.n570 B.n46 10.6151
R1727 B.n566 B.n46 10.6151
R1728 B.n566 B.n565 10.6151
R1729 B.n565 B.n564 10.6151
R1730 B.n564 B.n48 10.6151
R1731 B.n560 B.n48 10.6151
R1732 B.n560 B.n559 10.6151
R1733 B.n557 B.n52 10.6151
R1734 B.n553 B.n52 10.6151
R1735 B.n553 B.n552 10.6151
R1736 B.n552 B.n551 10.6151
R1737 B.n551 B.n54 10.6151
R1738 B.n547 B.n54 10.6151
R1739 B.n547 B.n546 10.6151
R1740 B.n546 B.n545 10.6151
R1741 B.n545 B.n56 10.6151
R1742 B.n541 B.n56 10.6151
R1743 B.n541 B.n540 10.6151
R1744 B.n540 B.n539 10.6151
R1745 B.n539 B.n58 10.6151
R1746 B.n535 B.n58 10.6151
R1747 B.n535 B.n534 10.6151
R1748 B.n534 B.n533 10.6151
R1749 B.n533 B.n60 10.6151
R1750 B.n529 B.n60 10.6151
R1751 B.n529 B.n528 10.6151
R1752 B.n528 B.n527 10.6151
R1753 B.n527 B.n62 10.6151
R1754 B.n523 B.n62 10.6151
R1755 B.n523 B.n522 10.6151
R1756 B.n522 B.n521 10.6151
R1757 B.n521 B.n64 10.6151
R1758 B.n517 B.n64 10.6151
R1759 B.n517 B.n516 10.6151
R1760 B.n516 B.n515 10.6151
R1761 B.n515 B.n66 10.6151
R1762 B.n511 B.n66 10.6151
R1763 B.n511 B.n510 10.6151
R1764 B.n510 B.n509 10.6151
R1765 B.n509 B.n68 10.6151
R1766 B.n505 B.n68 10.6151
R1767 B.n505 B.n504 10.6151
R1768 B.n504 B.n503 10.6151
R1769 B.n503 B.n70 10.6151
R1770 B.n499 B.n70 10.6151
R1771 B.n499 B.n498 10.6151
R1772 B.n498 B.n497 10.6151
R1773 B.n497 B.n72 10.6151
R1774 B.n493 B.n72 10.6151
R1775 B.n493 B.n492 10.6151
R1776 B.n384 B.n383 10.6151
R1777 B.n385 B.n384 10.6151
R1778 B.n385 B.n108 10.6151
R1779 B.n389 B.n108 10.6151
R1780 B.n390 B.n389 10.6151
R1781 B.n391 B.n390 10.6151
R1782 B.n391 B.n106 10.6151
R1783 B.n395 B.n106 10.6151
R1784 B.n396 B.n395 10.6151
R1785 B.n397 B.n396 10.6151
R1786 B.n397 B.n104 10.6151
R1787 B.n401 B.n104 10.6151
R1788 B.n402 B.n401 10.6151
R1789 B.n403 B.n402 10.6151
R1790 B.n403 B.n102 10.6151
R1791 B.n407 B.n102 10.6151
R1792 B.n408 B.n407 10.6151
R1793 B.n409 B.n408 10.6151
R1794 B.n409 B.n100 10.6151
R1795 B.n413 B.n100 10.6151
R1796 B.n414 B.n413 10.6151
R1797 B.n415 B.n414 10.6151
R1798 B.n415 B.n98 10.6151
R1799 B.n419 B.n98 10.6151
R1800 B.n420 B.n419 10.6151
R1801 B.n421 B.n420 10.6151
R1802 B.n421 B.n96 10.6151
R1803 B.n425 B.n96 10.6151
R1804 B.n426 B.n425 10.6151
R1805 B.n427 B.n426 10.6151
R1806 B.n427 B.n94 10.6151
R1807 B.n431 B.n94 10.6151
R1808 B.n432 B.n431 10.6151
R1809 B.n433 B.n432 10.6151
R1810 B.n433 B.n92 10.6151
R1811 B.n437 B.n92 10.6151
R1812 B.n438 B.n437 10.6151
R1813 B.n439 B.n438 10.6151
R1814 B.n439 B.n90 10.6151
R1815 B.n443 B.n90 10.6151
R1816 B.n444 B.n443 10.6151
R1817 B.n445 B.n444 10.6151
R1818 B.n445 B.n88 10.6151
R1819 B.n449 B.n88 10.6151
R1820 B.n450 B.n449 10.6151
R1821 B.n451 B.n450 10.6151
R1822 B.n451 B.n86 10.6151
R1823 B.n455 B.n86 10.6151
R1824 B.n456 B.n455 10.6151
R1825 B.n457 B.n456 10.6151
R1826 B.n457 B.n84 10.6151
R1827 B.n461 B.n84 10.6151
R1828 B.n462 B.n461 10.6151
R1829 B.n463 B.n462 10.6151
R1830 B.n463 B.n82 10.6151
R1831 B.n467 B.n82 10.6151
R1832 B.n468 B.n467 10.6151
R1833 B.n469 B.n468 10.6151
R1834 B.n469 B.n80 10.6151
R1835 B.n473 B.n80 10.6151
R1836 B.n474 B.n473 10.6151
R1837 B.n475 B.n474 10.6151
R1838 B.n475 B.n78 10.6151
R1839 B.n479 B.n78 10.6151
R1840 B.n480 B.n479 10.6151
R1841 B.n481 B.n480 10.6151
R1842 B.n481 B.n76 10.6151
R1843 B.n485 B.n76 10.6151
R1844 B.n486 B.n485 10.6151
R1845 B.n487 B.n486 10.6151
R1846 B.n487 B.n74 10.6151
R1847 B.n491 B.n74 10.6151
R1848 B.n235 B.n234 10.6151
R1849 B.n235 B.n162 10.6151
R1850 B.n239 B.n162 10.6151
R1851 B.n240 B.n239 10.6151
R1852 B.n241 B.n240 10.6151
R1853 B.n241 B.n160 10.6151
R1854 B.n245 B.n160 10.6151
R1855 B.n246 B.n245 10.6151
R1856 B.n247 B.n246 10.6151
R1857 B.n247 B.n158 10.6151
R1858 B.n251 B.n158 10.6151
R1859 B.n252 B.n251 10.6151
R1860 B.n253 B.n252 10.6151
R1861 B.n253 B.n156 10.6151
R1862 B.n257 B.n156 10.6151
R1863 B.n258 B.n257 10.6151
R1864 B.n259 B.n258 10.6151
R1865 B.n259 B.n154 10.6151
R1866 B.n263 B.n154 10.6151
R1867 B.n264 B.n263 10.6151
R1868 B.n265 B.n264 10.6151
R1869 B.n265 B.n152 10.6151
R1870 B.n269 B.n152 10.6151
R1871 B.n270 B.n269 10.6151
R1872 B.n271 B.n270 10.6151
R1873 B.n271 B.n150 10.6151
R1874 B.n275 B.n150 10.6151
R1875 B.n276 B.n275 10.6151
R1876 B.n277 B.n276 10.6151
R1877 B.n277 B.n148 10.6151
R1878 B.n281 B.n148 10.6151
R1879 B.n282 B.n281 10.6151
R1880 B.n283 B.n282 10.6151
R1881 B.n283 B.n146 10.6151
R1882 B.n287 B.n146 10.6151
R1883 B.n288 B.n287 10.6151
R1884 B.n289 B.n288 10.6151
R1885 B.n289 B.n144 10.6151
R1886 B.n293 B.n144 10.6151
R1887 B.n294 B.n293 10.6151
R1888 B.n295 B.n294 10.6151
R1889 B.n295 B.n142 10.6151
R1890 B.n299 B.n142 10.6151
R1891 B.n302 B.n301 10.6151
R1892 B.n302 B.n138 10.6151
R1893 B.n306 B.n138 10.6151
R1894 B.n307 B.n306 10.6151
R1895 B.n308 B.n307 10.6151
R1896 B.n308 B.n136 10.6151
R1897 B.n312 B.n136 10.6151
R1898 B.n313 B.n312 10.6151
R1899 B.n314 B.n313 10.6151
R1900 B.n318 B.n317 10.6151
R1901 B.n319 B.n318 10.6151
R1902 B.n319 B.n130 10.6151
R1903 B.n323 B.n130 10.6151
R1904 B.n324 B.n323 10.6151
R1905 B.n325 B.n324 10.6151
R1906 B.n325 B.n128 10.6151
R1907 B.n329 B.n128 10.6151
R1908 B.n330 B.n329 10.6151
R1909 B.n331 B.n330 10.6151
R1910 B.n331 B.n126 10.6151
R1911 B.n335 B.n126 10.6151
R1912 B.n336 B.n335 10.6151
R1913 B.n337 B.n336 10.6151
R1914 B.n337 B.n124 10.6151
R1915 B.n341 B.n124 10.6151
R1916 B.n342 B.n341 10.6151
R1917 B.n343 B.n342 10.6151
R1918 B.n343 B.n122 10.6151
R1919 B.n347 B.n122 10.6151
R1920 B.n348 B.n347 10.6151
R1921 B.n349 B.n348 10.6151
R1922 B.n349 B.n120 10.6151
R1923 B.n353 B.n120 10.6151
R1924 B.n354 B.n353 10.6151
R1925 B.n355 B.n354 10.6151
R1926 B.n355 B.n118 10.6151
R1927 B.n359 B.n118 10.6151
R1928 B.n360 B.n359 10.6151
R1929 B.n361 B.n360 10.6151
R1930 B.n361 B.n116 10.6151
R1931 B.n365 B.n116 10.6151
R1932 B.n366 B.n365 10.6151
R1933 B.n367 B.n366 10.6151
R1934 B.n367 B.n114 10.6151
R1935 B.n371 B.n114 10.6151
R1936 B.n372 B.n371 10.6151
R1937 B.n373 B.n372 10.6151
R1938 B.n373 B.n112 10.6151
R1939 B.n377 B.n112 10.6151
R1940 B.n378 B.n377 10.6151
R1941 B.n379 B.n378 10.6151
R1942 B.n379 B.n110 10.6151
R1943 B.n233 B.n164 10.6151
R1944 B.n229 B.n164 10.6151
R1945 B.n229 B.n228 10.6151
R1946 B.n228 B.n227 10.6151
R1947 B.n227 B.n166 10.6151
R1948 B.n223 B.n166 10.6151
R1949 B.n223 B.n222 10.6151
R1950 B.n222 B.n221 10.6151
R1951 B.n221 B.n168 10.6151
R1952 B.n217 B.n168 10.6151
R1953 B.n217 B.n216 10.6151
R1954 B.n216 B.n215 10.6151
R1955 B.n215 B.n170 10.6151
R1956 B.n211 B.n170 10.6151
R1957 B.n211 B.n210 10.6151
R1958 B.n210 B.n209 10.6151
R1959 B.n209 B.n172 10.6151
R1960 B.n205 B.n172 10.6151
R1961 B.n205 B.n204 10.6151
R1962 B.n204 B.n203 10.6151
R1963 B.n203 B.n174 10.6151
R1964 B.n199 B.n174 10.6151
R1965 B.n199 B.n198 10.6151
R1966 B.n198 B.n197 10.6151
R1967 B.n197 B.n176 10.6151
R1968 B.n193 B.n176 10.6151
R1969 B.n193 B.n192 10.6151
R1970 B.n192 B.n191 10.6151
R1971 B.n191 B.n178 10.6151
R1972 B.n187 B.n178 10.6151
R1973 B.n187 B.n186 10.6151
R1974 B.n186 B.n185 10.6151
R1975 B.n185 B.n180 10.6151
R1976 B.n181 B.n180 10.6151
R1977 B.n181 B.n0 10.6151
R1978 B.n691 B.n1 10.6151
R1979 B.n691 B.n690 10.6151
R1980 B.n690 B.n689 10.6151
R1981 B.n689 B.n4 10.6151
R1982 B.n685 B.n4 10.6151
R1983 B.n685 B.n684 10.6151
R1984 B.n684 B.n683 10.6151
R1985 B.n683 B.n6 10.6151
R1986 B.n679 B.n6 10.6151
R1987 B.n679 B.n678 10.6151
R1988 B.n678 B.n677 10.6151
R1989 B.n677 B.n8 10.6151
R1990 B.n673 B.n8 10.6151
R1991 B.n673 B.n672 10.6151
R1992 B.n672 B.n671 10.6151
R1993 B.n671 B.n10 10.6151
R1994 B.n667 B.n10 10.6151
R1995 B.n667 B.n666 10.6151
R1996 B.n666 B.n665 10.6151
R1997 B.n665 B.n12 10.6151
R1998 B.n661 B.n12 10.6151
R1999 B.n661 B.n660 10.6151
R2000 B.n660 B.n659 10.6151
R2001 B.n659 B.n14 10.6151
R2002 B.n655 B.n14 10.6151
R2003 B.n655 B.n654 10.6151
R2004 B.n654 B.n653 10.6151
R2005 B.n653 B.n16 10.6151
R2006 B.n649 B.n16 10.6151
R2007 B.n649 B.n648 10.6151
R2008 B.n648 B.n647 10.6151
R2009 B.n647 B.n18 10.6151
R2010 B.n643 B.n18 10.6151
R2011 B.n643 B.n642 10.6151
R2012 B.n642 B.n641 10.6151
R2013 B.n575 B.n44 9.36635
R2014 B.n558 B.n557 9.36635
R2015 B.n300 B.n299 9.36635
R2016 B.n317 B.n134 9.36635
R2017 B.n695 B.n0 2.81026
R2018 B.n695 B.n1 2.81026
R2019 B.n572 B.n44 1.24928
R2020 B.n559 B.n558 1.24928
R2021 B.n301 B.n300 1.24928
R2022 B.n314 B.n134 1.24928
C0 VDD2 VDD1 1.20223f
C1 VTAIL VDD2 8.10218f
C2 VDD2 w_n2874_n3536# 2.28614f
C3 VTAIL VDD1 8.05597f
C4 w_n2874_n3536# VDD1 2.21859f
C5 VTAIL w_n2874_n3536# 3.05802f
C6 VDD2 VP 0.412212f
C7 VN B 1.06424f
C8 VP VDD1 7.07084f
C9 VTAIL VP 6.8227f
C10 w_n2874_n3536# VP 5.69266f
C11 B VDD2 2.07307f
C12 B VDD1 2.01217f
C13 VTAIL B 3.63639f
C14 B w_n2874_n3536# 9.151421f
C15 VN VDD2 6.81258f
C16 B VP 1.67928f
C17 VN VDD1 0.150394f
C18 VTAIL VN 6.80835f
C19 VN w_n2874_n3536# 5.32262f
C20 VN VP 6.54518f
C21 VDD2 VSUBS 1.795007f
C22 VDD1 VSUBS 1.658889f
C23 VTAIL VSUBS 1.117785f
C24 VN VSUBS 5.3591f
C25 VP VSUBS 2.545576f
C26 B VSUBS 4.164638f
C27 w_n2874_n3536# VSUBS 0.12495p
C28 B.n0 VSUBS 0.00524f
C29 B.n1 VSUBS 0.00524f
C30 B.n2 VSUBS 0.008287f
C31 B.n3 VSUBS 0.008287f
C32 B.n4 VSUBS 0.008287f
C33 B.n5 VSUBS 0.008287f
C34 B.n6 VSUBS 0.008287f
C35 B.n7 VSUBS 0.008287f
C36 B.n8 VSUBS 0.008287f
C37 B.n9 VSUBS 0.008287f
C38 B.n10 VSUBS 0.008287f
C39 B.n11 VSUBS 0.008287f
C40 B.n12 VSUBS 0.008287f
C41 B.n13 VSUBS 0.008287f
C42 B.n14 VSUBS 0.008287f
C43 B.n15 VSUBS 0.008287f
C44 B.n16 VSUBS 0.008287f
C45 B.n17 VSUBS 0.008287f
C46 B.n18 VSUBS 0.008287f
C47 B.n19 VSUBS 0.008287f
C48 B.n20 VSUBS 0.019919f
C49 B.n21 VSUBS 0.008287f
C50 B.n22 VSUBS 0.008287f
C51 B.n23 VSUBS 0.008287f
C52 B.n24 VSUBS 0.008287f
C53 B.n25 VSUBS 0.008287f
C54 B.n26 VSUBS 0.008287f
C55 B.n27 VSUBS 0.008287f
C56 B.n28 VSUBS 0.008287f
C57 B.n29 VSUBS 0.008287f
C58 B.n30 VSUBS 0.008287f
C59 B.n31 VSUBS 0.008287f
C60 B.n32 VSUBS 0.008287f
C61 B.n33 VSUBS 0.008287f
C62 B.n34 VSUBS 0.008287f
C63 B.n35 VSUBS 0.008287f
C64 B.n36 VSUBS 0.008287f
C65 B.n37 VSUBS 0.008287f
C66 B.n38 VSUBS 0.008287f
C67 B.n39 VSUBS 0.008287f
C68 B.n40 VSUBS 0.008287f
C69 B.n41 VSUBS 0.008287f
C70 B.t5 VSUBS 0.272306f
C71 B.t4 VSUBS 0.303684f
C72 B.t3 VSUBS 1.38944f
C73 B.n42 VSUBS 0.470905f
C74 B.n43 VSUBS 0.308918f
C75 B.n44 VSUBS 0.0192f
C76 B.n45 VSUBS 0.008287f
C77 B.n46 VSUBS 0.008287f
C78 B.n47 VSUBS 0.008287f
C79 B.n48 VSUBS 0.008287f
C80 B.n49 VSUBS 0.008287f
C81 B.t11 VSUBS 0.27231f
C82 B.t10 VSUBS 0.303687f
C83 B.t9 VSUBS 1.38944f
C84 B.n50 VSUBS 0.470901f
C85 B.n51 VSUBS 0.308915f
C86 B.n52 VSUBS 0.008287f
C87 B.n53 VSUBS 0.008287f
C88 B.n54 VSUBS 0.008287f
C89 B.n55 VSUBS 0.008287f
C90 B.n56 VSUBS 0.008287f
C91 B.n57 VSUBS 0.008287f
C92 B.n58 VSUBS 0.008287f
C93 B.n59 VSUBS 0.008287f
C94 B.n60 VSUBS 0.008287f
C95 B.n61 VSUBS 0.008287f
C96 B.n62 VSUBS 0.008287f
C97 B.n63 VSUBS 0.008287f
C98 B.n64 VSUBS 0.008287f
C99 B.n65 VSUBS 0.008287f
C100 B.n66 VSUBS 0.008287f
C101 B.n67 VSUBS 0.008287f
C102 B.n68 VSUBS 0.008287f
C103 B.n69 VSUBS 0.008287f
C104 B.n70 VSUBS 0.008287f
C105 B.n71 VSUBS 0.008287f
C106 B.n72 VSUBS 0.008287f
C107 B.n73 VSUBS 0.019919f
C108 B.n74 VSUBS 0.008287f
C109 B.n75 VSUBS 0.008287f
C110 B.n76 VSUBS 0.008287f
C111 B.n77 VSUBS 0.008287f
C112 B.n78 VSUBS 0.008287f
C113 B.n79 VSUBS 0.008287f
C114 B.n80 VSUBS 0.008287f
C115 B.n81 VSUBS 0.008287f
C116 B.n82 VSUBS 0.008287f
C117 B.n83 VSUBS 0.008287f
C118 B.n84 VSUBS 0.008287f
C119 B.n85 VSUBS 0.008287f
C120 B.n86 VSUBS 0.008287f
C121 B.n87 VSUBS 0.008287f
C122 B.n88 VSUBS 0.008287f
C123 B.n89 VSUBS 0.008287f
C124 B.n90 VSUBS 0.008287f
C125 B.n91 VSUBS 0.008287f
C126 B.n92 VSUBS 0.008287f
C127 B.n93 VSUBS 0.008287f
C128 B.n94 VSUBS 0.008287f
C129 B.n95 VSUBS 0.008287f
C130 B.n96 VSUBS 0.008287f
C131 B.n97 VSUBS 0.008287f
C132 B.n98 VSUBS 0.008287f
C133 B.n99 VSUBS 0.008287f
C134 B.n100 VSUBS 0.008287f
C135 B.n101 VSUBS 0.008287f
C136 B.n102 VSUBS 0.008287f
C137 B.n103 VSUBS 0.008287f
C138 B.n104 VSUBS 0.008287f
C139 B.n105 VSUBS 0.008287f
C140 B.n106 VSUBS 0.008287f
C141 B.n107 VSUBS 0.008287f
C142 B.n108 VSUBS 0.008287f
C143 B.n109 VSUBS 0.008287f
C144 B.n110 VSUBS 0.019919f
C145 B.n111 VSUBS 0.008287f
C146 B.n112 VSUBS 0.008287f
C147 B.n113 VSUBS 0.008287f
C148 B.n114 VSUBS 0.008287f
C149 B.n115 VSUBS 0.008287f
C150 B.n116 VSUBS 0.008287f
C151 B.n117 VSUBS 0.008287f
C152 B.n118 VSUBS 0.008287f
C153 B.n119 VSUBS 0.008287f
C154 B.n120 VSUBS 0.008287f
C155 B.n121 VSUBS 0.008287f
C156 B.n122 VSUBS 0.008287f
C157 B.n123 VSUBS 0.008287f
C158 B.n124 VSUBS 0.008287f
C159 B.n125 VSUBS 0.008287f
C160 B.n126 VSUBS 0.008287f
C161 B.n127 VSUBS 0.008287f
C162 B.n128 VSUBS 0.008287f
C163 B.n129 VSUBS 0.008287f
C164 B.n130 VSUBS 0.008287f
C165 B.n131 VSUBS 0.008287f
C166 B.t1 VSUBS 0.27231f
C167 B.t2 VSUBS 0.303687f
C168 B.t0 VSUBS 1.38944f
C169 B.n132 VSUBS 0.470901f
C170 B.n133 VSUBS 0.308915f
C171 B.n134 VSUBS 0.0192f
C172 B.n135 VSUBS 0.008287f
C173 B.n136 VSUBS 0.008287f
C174 B.n137 VSUBS 0.008287f
C175 B.n138 VSUBS 0.008287f
C176 B.n139 VSUBS 0.008287f
C177 B.t7 VSUBS 0.272306f
C178 B.t8 VSUBS 0.303684f
C179 B.t6 VSUBS 1.38944f
C180 B.n140 VSUBS 0.470905f
C181 B.n141 VSUBS 0.308918f
C182 B.n142 VSUBS 0.008287f
C183 B.n143 VSUBS 0.008287f
C184 B.n144 VSUBS 0.008287f
C185 B.n145 VSUBS 0.008287f
C186 B.n146 VSUBS 0.008287f
C187 B.n147 VSUBS 0.008287f
C188 B.n148 VSUBS 0.008287f
C189 B.n149 VSUBS 0.008287f
C190 B.n150 VSUBS 0.008287f
C191 B.n151 VSUBS 0.008287f
C192 B.n152 VSUBS 0.008287f
C193 B.n153 VSUBS 0.008287f
C194 B.n154 VSUBS 0.008287f
C195 B.n155 VSUBS 0.008287f
C196 B.n156 VSUBS 0.008287f
C197 B.n157 VSUBS 0.008287f
C198 B.n158 VSUBS 0.008287f
C199 B.n159 VSUBS 0.008287f
C200 B.n160 VSUBS 0.008287f
C201 B.n161 VSUBS 0.008287f
C202 B.n162 VSUBS 0.008287f
C203 B.n163 VSUBS 0.019919f
C204 B.n164 VSUBS 0.008287f
C205 B.n165 VSUBS 0.008287f
C206 B.n166 VSUBS 0.008287f
C207 B.n167 VSUBS 0.008287f
C208 B.n168 VSUBS 0.008287f
C209 B.n169 VSUBS 0.008287f
C210 B.n170 VSUBS 0.008287f
C211 B.n171 VSUBS 0.008287f
C212 B.n172 VSUBS 0.008287f
C213 B.n173 VSUBS 0.008287f
C214 B.n174 VSUBS 0.008287f
C215 B.n175 VSUBS 0.008287f
C216 B.n176 VSUBS 0.008287f
C217 B.n177 VSUBS 0.008287f
C218 B.n178 VSUBS 0.008287f
C219 B.n179 VSUBS 0.008287f
C220 B.n180 VSUBS 0.008287f
C221 B.n181 VSUBS 0.008287f
C222 B.n182 VSUBS 0.008287f
C223 B.n183 VSUBS 0.008287f
C224 B.n184 VSUBS 0.008287f
C225 B.n185 VSUBS 0.008287f
C226 B.n186 VSUBS 0.008287f
C227 B.n187 VSUBS 0.008287f
C228 B.n188 VSUBS 0.008287f
C229 B.n189 VSUBS 0.008287f
C230 B.n190 VSUBS 0.008287f
C231 B.n191 VSUBS 0.008287f
C232 B.n192 VSUBS 0.008287f
C233 B.n193 VSUBS 0.008287f
C234 B.n194 VSUBS 0.008287f
C235 B.n195 VSUBS 0.008287f
C236 B.n196 VSUBS 0.008287f
C237 B.n197 VSUBS 0.008287f
C238 B.n198 VSUBS 0.008287f
C239 B.n199 VSUBS 0.008287f
C240 B.n200 VSUBS 0.008287f
C241 B.n201 VSUBS 0.008287f
C242 B.n202 VSUBS 0.008287f
C243 B.n203 VSUBS 0.008287f
C244 B.n204 VSUBS 0.008287f
C245 B.n205 VSUBS 0.008287f
C246 B.n206 VSUBS 0.008287f
C247 B.n207 VSUBS 0.008287f
C248 B.n208 VSUBS 0.008287f
C249 B.n209 VSUBS 0.008287f
C250 B.n210 VSUBS 0.008287f
C251 B.n211 VSUBS 0.008287f
C252 B.n212 VSUBS 0.008287f
C253 B.n213 VSUBS 0.008287f
C254 B.n214 VSUBS 0.008287f
C255 B.n215 VSUBS 0.008287f
C256 B.n216 VSUBS 0.008287f
C257 B.n217 VSUBS 0.008287f
C258 B.n218 VSUBS 0.008287f
C259 B.n219 VSUBS 0.008287f
C260 B.n220 VSUBS 0.008287f
C261 B.n221 VSUBS 0.008287f
C262 B.n222 VSUBS 0.008287f
C263 B.n223 VSUBS 0.008287f
C264 B.n224 VSUBS 0.008287f
C265 B.n225 VSUBS 0.008287f
C266 B.n226 VSUBS 0.008287f
C267 B.n227 VSUBS 0.008287f
C268 B.n228 VSUBS 0.008287f
C269 B.n229 VSUBS 0.008287f
C270 B.n230 VSUBS 0.008287f
C271 B.n231 VSUBS 0.008287f
C272 B.n232 VSUBS 0.018592f
C273 B.n233 VSUBS 0.018592f
C274 B.n234 VSUBS 0.019919f
C275 B.n235 VSUBS 0.008287f
C276 B.n236 VSUBS 0.008287f
C277 B.n237 VSUBS 0.008287f
C278 B.n238 VSUBS 0.008287f
C279 B.n239 VSUBS 0.008287f
C280 B.n240 VSUBS 0.008287f
C281 B.n241 VSUBS 0.008287f
C282 B.n242 VSUBS 0.008287f
C283 B.n243 VSUBS 0.008287f
C284 B.n244 VSUBS 0.008287f
C285 B.n245 VSUBS 0.008287f
C286 B.n246 VSUBS 0.008287f
C287 B.n247 VSUBS 0.008287f
C288 B.n248 VSUBS 0.008287f
C289 B.n249 VSUBS 0.008287f
C290 B.n250 VSUBS 0.008287f
C291 B.n251 VSUBS 0.008287f
C292 B.n252 VSUBS 0.008287f
C293 B.n253 VSUBS 0.008287f
C294 B.n254 VSUBS 0.008287f
C295 B.n255 VSUBS 0.008287f
C296 B.n256 VSUBS 0.008287f
C297 B.n257 VSUBS 0.008287f
C298 B.n258 VSUBS 0.008287f
C299 B.n259 VSUBS 0.008287f
C300 B.n260 VSUBS 0.008287f
C301 B.n261 VSUBS 0.008287f
C302 B.n262 VSUBS 0.008287f
C303 B.n263 VSUBS 0.008287f
C304 B.n264 VSUBS 0.008287f
C305 B.n265 VSUBS 0.008287f
C306 B.n266 VSUBS 0.008287f
C307 B.n267 VSUBS 0.008287f
C308 B.n268 VSUBS 0.008287f
C309 B.n269 VSUBS 0.008287f
C310 B.n270 VSUBS 0.008287f
C311 B.n271 VSUBS 0.008287f
C312 B.n272 VSUBS 0.008287f
C313 B.n273 VSUBS 0.008287f
C314 B.n274 VSUBS 0.008287f
C315 B.n275 VSUBS 0.008287f
C316 B.n276 VSUBS 0.008287f
C317 B.n277 VSUBS 0.008287f
C318 B.n278 VSUBS 0.008287f
C319 B.n279 VSUBS 0.008287f
C320 B.n280 VSUBS 0.008287f
C321 B.n281 VSUBS 0.008287f
C322 B.n282 VSUBS 0.008287f
C323 B.n283 VSUBS 0.008287f
C324 B.n284 VSUBS 0.008287f
C325 B.n285 VSUBS 0.008287f
C326 B.n286 VSUBS 0.008287f
C327 B.n287 VSUBS 0.008287f
C328 B.n288 VSUBS 0.008287f
C329 B.n289 VSUBS 0.008287f
C330 B.n290 VSUBS 0.008287f
C331 B.n291 VSUBS 0.008287f
C332 B.n292 VSUBS 0.008287f
C333 B.n293 VSUBS 0.008287f
C334 B.n294 VSUBS 0.008287f
C335 B.n295 VSUBS 0.008287f
C336 B.n296 VSUBS 0.008287f
C337 B.n297 VSUBS 0.008287f
C338 B.n298 VSUBS 0.008287f
C339 B.n299 VSUBS 0.0078f
C340 B.n300 VSUBS 0.0192f
C341 B.n301 VSUBS 0.004631f
C342 B.n302 VSUBS 0.008287f
C343 B.n303 VSUBS 0.008287f
C344 B.n304 VSUBS 0.008287f
C345 B.n305 VSUBS 0.008287f
C346 B.n306 VSUBS 0.008287f
C347 B.n307 VSUBS 0.008287f
C348 B.n308 VSUBS 0.008287f
C349 B.n309 VSUBS 0.008287f
C350 B.n310 VSUBS 0.008287f
C351 B.n311 VSUBS 0.008287f
C352 B.n312 VSUBS 0.008287f
C353 B.n313 VSUBS 0.008287f
C354 B.n314 VSUBS 0.004631f
C355 B.n315 VSUBS 0.008287f
C356 B.n316 VSUBS 0.008287f
C357 B.n317 VSUBS 0.0078f
C358 B.n318 VSUBS 0.008287f
C359 B.n319 VSUBS 0.008287f
C360 B.n320 VSUBS 0.008287f
C361 B.n321 VSUBS 0.008287f
C362 B.n322 VSUBS 0.008287f
C363 B.n323 VSUBS 0.008287f
C364 B.n324 VSUBS 0.008287f
C365 B.n325 VSUBS 0.008287f
C366 B.n326 VSUBS 0.008287f
C367 B.n327 VSUBS 0.008287f
C368 B.n328 VSUBS 0.008287f
C369 B.n329 VSUBS 0.008287f
C370 B.n330 VSUBS 0.008287f
C371 B.n331 VSUBS 0.008287f
C372 B.n332 VSUBS 0.008287f
C373 B.n333 VSUBS 0.008287f
C374 B.n334 VSUBS 0.008287f
C375 B.n335 VSUBS 0.008287f
C376 B.n336 VSUBS 0.008287f
C377 B.n337 VSUBS 0.008287f
C378 B.n338 VSUBS 0.008287f
C379 B.n339 VSUBS 0.008287f
C380 B.n340 VSUBS 0.008287f
C381 B.n341 VSUBS 0.008287f
C382 B.n342 VSUBS 0.008287f
C383 B.n343 VSUBS 0.008287f
C384 B.n344 VSUBS 0.008287f
C385 B.n345 VSUBS 0.008287f
C386 B.n346 VSUBS 0.008287f
C387 B.n347 VSUBS 0.008287f
C388 B.n348 VSUBS 0.008287f
C389 B.n349 VSUBS 0.008287f
C390 B.n350 VSUBS 0.008287f
C391 B.n351 VSUBS 0.008287f
C392 B.n352 VSUBS 0.008287f
C393 B.n353 VSUBS 0.008287f
C394 B.n354 VSUBS 0.008287f
C395 B.n355 VSUBS 0.008287f
C396 B.n356 VSUBS 0.008287f
C397 B.n357 VSUBS 0.008287f
C398 B.n358 VSUBS 0.008287f
C399 B.n359 VSUBS 0.008287f
C400 B.n360 VSUBS 0.008287f
C401 B.n361 VSUBS 0.008287f
C402 B.n362 VSUBS 0.008287f
C403 B.n363 VSUBS 0.008287f
C404 B.n364 VSUBS 0.008287f
C405 B.n365 VSUBS 0.008287f
C406 B.n366 VSUBS 0.008287f
C407 B.n367 VSUBS 0.008287f
C408 B.n368 VSUBS 0.008287f
C409 B.n369 VSUBS 0.008287f
C410 B.n370 VSUBS 0.008287f
C411 B.n371 VSUBS 0.008287f
C412 B.n372 VSUBS 0.008287f
C413 B.n373 VSUBS 0.008287f
C414 B.n374 VSUBS 0.008287f
C415 B.n375 VSUBS 0.008287f
C416 B.n376 VSUBS 0.008287f
C417 B.n377 VSUBS 0.008287f
C418 B.n378 VSUBS 0.008287f
C419 B.n379 VSUBS 0.008287f
C420 B.n380 VSUBS 0.008287f
C421 B.n381 VSUBS 0.019919f
C422 B.n382 VSUBS 0.018592f
C423 B.n383 VSUBS 0.018592f
C424 B.n384 VSUBS 0.008287f
C425 B.n385 VSUBS 0.008287f
C426 B.n386 VSUBS 0.008287f
C427 B.n387 VSUBS 0.008287f
C428 B.n388 VSUBS 0.008287f
C429 B.n389 VSUBS 0.008287f
C430 B.n390 VSUBS 0.008287f
C431 B.n391 VSUBS 0.008287f
C432 B.n392 VSUBS 0.008287f
C433 B.n393 VSUBS 0.008287f
C434 B.n394 VSUBS 0.008287f
C435 B.n395 VSUBS 0.008287f
C436 B.n396 VSUBS 0.008287f
C437 B.n397 VSUBS 0.008287f
C438 B.n398 VSUBS 0.008287f
C439 B.n399 VSUBS 0.008287f
C440 B.n400 VSUBS 0.008287f
C441 B.n401 VSUBS 0.008287f
C442 B.n402 VSUBS 0.008287f
C443 B.n403 VSUBS 0.008287f
C444 B.n404 VSUBS 0.008287f
C445 B.n405 VSUBS 0.008287f
C446 B.n406 VSUBS 0.008287f
C447 B.n407 VSUBS 0.008287f
C448 B.n408 VSUBS 0.008287f
C449 B.n409 VSUBS 0.008287f
C450 B.n410 VSUBS 0.008287f
C451 B.n411 VSUBS 0.008287f
C452 B.n412 VSUBS 0.008287f
C453 B.n413 VSUBS 0.008287f
C454 B.n414 VSUBS 0.008287f
C455 B.n415 VSUBS 0.008287f
C456 B.n416 VSUBS 0.008287f
C457 B.n417 VSUBS 0.008287f
C458 B.n418 VSUBS 0.008287f
C459 B.n419 VSUBS 0.008287f
C460 B.n420 VSUBS 0.008287f
C461 B.n421 VSUBS 0.008287f
C462 B.n422 VSUBS 0.008287f
C463 B.n423 VSUBS 0.008287f
C464 B.n424 VSUBS 0.008287f
C465 B.n425 VSUBS 0.008287f
C466 B.n426 VSUBS 0.008287f
C467 B.n427 VSUBS 0.008287f
C468 B.n428 VSUBS 0.008287f
C469 B.n429 VSUBS 0.008287f
C470 B.n430 VSUBS 0.008287f
C471 B.n431 VSUBS 0.008287f
C472 B.n432 VSUBS 0.008287f
C473 B.n433 VSUBS 0.008287f
C474 B.n434 VSUBS 0.008287f
C475 B.n435 VSUBS 0.008287f
C476 B.n436 VSUBS 0.008287f
C477 B.n437 VSUBS 0.008287f
C478 B.n438 VSUBS 0.008287f
C479 B.n439 VSUBS 0.008287f
C480 B.n440 VSUBS 0.008287f
C481 B.n441 VSUBS 0.008287f
C482 B.n442 VSUBS 0.008287f
C483 B.n443 VSUBS 0.008287f
C484 B.n444 VSUBS 0.008287f
C485 B.n445 VSUBS 0.008287f
C486 B.n446 VSUBS 0.008287f
C487 B.n447 VSUBS 0.008287f
C488 B.n448 VSUBS 0.008287f
C489 B.n449 VSUBS 0.008287f
C490 B.n450 VSUBS 0.008287f
C491 B.n451 VSUBS 0.008287f
C492 B.n452 VSUBS 0.008287f
C493 B.n453 VSUBS 0.008287f
C494 B.n454 VSUBS 0.008287f
C495 B.n455 VSUBS 0.008287f
C496 B.n456 VSUBS 0.008287f
C497 B.n457 VSUBS 0.008287f
C498 B.n458 VSUBS 0.008287f
C499 B.n459 VSUBS 0.008287f
C500 B.n460 VSUBS 0.008287f
C501 B.n461 VSUBS 0.008287f
C502 B.n462 VSUBS 0.008287f
C503 B.n463 VSUBS 0.008287f
C504 B.n464 VSUBS 0.008287f
C505 B.n465 VSUBS 0.008287f
C506 B.n466 VSUBS 0.008287f
C507 B.n467 VSUBS 0.008287f
C508 B.n468 VSUBS 0.008287f
C509 B.n469 VSUBS 0.008287f
C510 B.n470 VSUBS 0.008287f
C511 B.n471 VSUBS 0.008287f
C512 B.n472 VSUBS 0.008287f
C513 B.n473 VSUBS 0.008287f
C514 B.n474 VSUBS 0.008287f
C515 B.n475 VSUBS 0.008287f
C516 B.n476 VSUBS 0.008287f
C517 B.n477 VSUBS 0.008287f
C518 B.n478 VSUBS 0.008287f
C519 B.n479 VSUBS 0.008287f
C520 B.n480 VSUBS 0.008287f
C521 B.n481 VSUBS 0.008287f
C522 B.n482 VSUBS 0.008287f
C523 B.n483 VSUBS 0.008287f
C524 B.n484 VSUBS 0.008287f
C525 B.n485 VSUBS 0.008287f
C526 B.n486 VSUBS 0.008287f
C527 B.n487 VSUBS 0.008287f
C528 B.n488 VSUBS 0.008287f
C529 B.n489 VSUBS 0.008287f
C530 B.n490 VSUBS 0.018592f
C531 B.n491 VSUBS 0.019581f
C532 B.n492 VSUBS 0.01893f
C533 B.n493 VSUBS 0.008287f
C534 B.n494 VSUBS 0.008287f
C535 B.n495 VSUBS 0.008287f
C536 B.n496 VSUBS 0.008287f
C537 B.n497 VSUBS 0.008287f
C538 B.n498 VSUBS 0.008287f
C539 B.n499 VSUBS 0.008287f
C540 B.n500 VSUBS 0.008287f
C541 B.n501 VSUBS 0.008287f
C542 B.n502 VSUBS 0.008287f
C543 B.n503 VSUBS 0.008287f
C544 B.n504 VSUBS 0.008287f
C545 B.n505 VSUBS 0.008287f
C546 B.n506 VSUBS 0.008287f
C547 B.n507 VSUBS 0.008287f
C548 B.n508 VSUBS 0.008287f
C549 B.n509 VSUBS 0.008287f
C550 B.n510 VSUBS 0.008287f
C551 B.n511 VSUBS 0.008287f
C552 B.n512 VSUBS 0.008287f
C553 B.n513 VSUBS 0.008287f
C554 B.n514 VSUBS 0.008287f
C555 B.n515 VSUBS 0.008287f
C556 B.n516 VSUBS 0.008287f
C557 B.n517 VSUBS 0.008287f
C558 B.n518 VSUBS 0.008287f
C559 B.n519 VSUBS 0.008287f
C560 B.n520 VSUBS 0.008287f
C561 B.n521 VSUBS 0.008287f
C562 B.n522 VSUBS 0.008287f
C563 B.n523 VSUBS 0.008287f
C564 B.n524 VSUBS 0.008287f
C565 B.n525 VSUBS 0.008287f
C566 B.n526 VSUBS 0.008287f
C567 B.n527 VSUBS 0.008287f
C568 B.n528 VSUBS 0.008287f
C569 B.n529 VSUBS 0.008287f
C570 B.n530 VSUBS 0.008287f
C571 B.n531 VSUBS 0.008287f
C572 B.n532 VSUBS 0.008287f
C573 B.n533 VSUBS 0.008287f
C574 B.n534 VSUBS 0.008287f
C575 B.n535 VSUBS 0.008287f
C576 B.n536 VSUBS 0.008287f
C577 B.n537 VSUBS 0.008287f
C578 B.n538 VSUBS 0.008287f
C579 B.n539 VSUBS 0.008287f
C580 B.n540 VSUBS 0.008287f
C581 B.n541 VSUBS 0.008287f
C582 B.n542 VSUBS 0.008287f
C583 B.n543 VSUBS 0.008287f
C584 B.n544 VSUBS 0.008287f
C585 B.n545 VSUBS 0.008287f
C586 B.n546 VSUBS 0.008287f
C587 B.n547 VSUBS 0.008287f
C588 B.n548 VSUBS 0.008287f
C589 B.n549 VSUBS 0.008287f
C590 B.n550 VSUBS 0.008287f
C591 B.n551 VSUBS 0.008287f
C592 B.n552 VSUBS 0.008287f
C593 B.n553 VSUBS 0.008287f
C594 B.n554 VSUBS 0.008287f
C595 B.n555 VSUBS 0.008287f
C596 B.n556 VSUBS 0.008287f
C597 B.n557 VSUBS 0.0078f
C598 B.n558 VSUBS 0.0192f
C599 B.n559 VSUBS 0.004631f
C600 B.n560 VSUBS 0.008287f
C601 B.n561 VSUBS 0.008287f
C602 B.n562 VSUBS 0.008287f
C603 B.n563 VSUBS 0.008287f
C604 B.n564 VSUBS 0.008287f
C605 B.n565 VSUBS 0.008287f
C606 B.n566 VSUBS 0.008287f
C607 B.n567 VSUBS 0.008287f
C608 B.n568 VSUBS 0.008287f
C609 B.n569 VSUBS 0.008287f
C610 B.n570 VSUBS 0.008287f
C611 B.n571 VSUBS 0.008287f
C612 B.n572 VSUBS 0.004631f
C613 B.n573 VSUBS 0.008287f
C614 B.n574 VSUBS 0.008287f
C615 B.n575 VSUBS 0.0078f
C616 B.n576 VSUBS 0.008287f
C617 B.n577 VSUBS 0.008287f
C618 B.n578 VSUBS 0.008287f
C619 B.n579 VSUBS 0.008287f
C620 B.n580 VSUBS 0.008287f
C621 B.n581 VSUBS 0.008287f
C622 B.n582 VSUBS 0.008287f
C623 B.n583 VSUBS 0.008287f
C624 B.n584 VSUBS 0.008287f
C625 B.n585 VSUBS 0.008287f
C626 B.n586 VSUBS 0.008287f
C627 B.n587 VSUBS 0.008287f
C628 B.n588 VSUBS 0.008287f
C629 B.n589 VSUBS 0.008287f
C630 B.n590 VSUBS 0.008287f
C631 B.n591 VSUBS 0.008287f
C632 B.n592 VSUBS 0.008287f
C633 B.n593 VSUBS 0.008287f
C634 B.n594 VSUBS 0.008287f
C635 B.n595 VSUBS 0.008287f
C636 B.n596 VSUBS 0.008287f
C637 B.n597 VSUBS 0.008287f
C638 B.n598 VSUBS 0.008287f
C639 B.n599 VSUBS 0.008287f
C640 B.n600 VSUBS 0.008287f
C641 B.n601 VSUBS 0.008287f
C642 B.n602 VSUBS 0.008287f
C643 B.n603 VSUBS 0.008287f
C644 B.n604 VSUBS 0.008287f
C645 B.n605 VSUBS 0.008287f
C646 B.n606 VSUBS 0.008287f
C647 B.n607 VSUBS 0.008287f
C648 B.n608 VSUBS 0.008287f
C649 B.n609 VSUBS 0.008287f
C650 B.n610 VSUBS 0.008287f
C651 B.n611 VSUBS 0.008287f
C652 B.n612 VSUBS 0.008287f
C653 B.n613 VSUBS 0.008287f
C654 B.n614 VSUBS 0.008287f
C655 B.n615 VSUBS 0.008287f
C656 B.n616 VSUBS 0.008287f
C657 B.n617 VSUBS 0.008287f
C658 B.n618 VSUBS 0.008287f
C659 B.n619 VSUBS 0.008287f
C660 B.n620 VSUBS 0.008287f
C661 B.n621 VSUBS 0.008287f
C662 B.n622 VSUBS 0.008287f
C663 B.n623 VSUBS 0.008287f
C664 B.n624 VSUBS 0.008287f
C665 B.n625 VSUBS 0.008287f
C666 B.n626 VSUBS 0.008287f
C667 B.n627 VSUBS 0.008287f
C668 B.n628 VSUBS 0.008287f
C669 B.n629 VSUBS 0.008287f
C670 B.n630 VSUBS 0.008287f
C671 B.n631 VSUBS 0.008287f
C672 B.n632 VSUBS 0.008287f
C673 B.n633 VSUBS 0.008287f
C674 B.n634 VSUBS 0.008287f
C675 B.n635 VSUBS 0.008287f
C676 B.n636 VSUBS 0.008287f
C677 B.n637 VSUBS 0.008287f
C678 B.n638 VSUBS 0.008287f
C679 B.n639 VSUBS 0.019919f
C680 B.n640 VSUBS 0.018592f
C681 B.n641 VSUBS 0.018592f
C682 B.n642 VSUBS 0.008287f
C683 B.n643 VSUBS 0.008287f
C684 B.n644 VSUBS 0.008287f
C685 B.n645 VSUBS 0.008287f
C686 B.n646 VSUBS 0.008287f
C687 B.n647 VSUBS 0.008287f
C688 B.n648 VSUBS 0.008287f
C689 B.n649 VSUBS 0.008287f
C690 B.n650 VSUBS 0.008287f
C691 B.n651 VSUBS 0.008287f
C692 B.n652 VSUBS 0.008287f
C693 B.n653 VSUBS 0.008287f
C694 B.n654 VSUBS 0.008287f
C695 B.n655 VSUBS 0.008287f
C696 B.n656 VSUBS 0.008287f
C697 B.n657 VSUBS 0.008287f
C698 B.n658 VSUBS 0.008287f
C699 B.n659 VSUBS 0.008287f
C700 B.n660 VSUBS 0.008287f
C701 B.n661 VSUBS 0.008287f
C702 B.n662 VSUBS 0.008287f
C703 B.n663 VSUBS 0.008287f
C704 B.n664 VSUBS 0.008287f
C705 B.n665 VSUBS 0.008287f
C706 B.n666 VSUBS 0.008287f
C707 B.n667 VSUBS 0.008287f
C708 B.n668 VSUBS 0.008287f
C709 B.n669 VSUBS 0.008287f
C710 B.n670 VSUBS 0.008287f
C711 B.n671 VSUBS 0.008287f
C712 B.n672 VSUBS 0.008287f
C713 B.n673 VSUBS 0.008287f
C714 B.n674 VSUBS 0.008287f
C715 B.n675 VSUBS 0.008287f
C716 B.n676 VSUBS 0.008287f
C717 B.n677 VSUBS 0.008287f
C718 B.n678 VSUBS 0.008287f
C719 B.n679 VSUBS 0.008287f
C720 B.n680 VSUBS 0.008287f
C721 B.n681 VSUBS 0.008287f
C722 B.n682 VSUBS 0.008287f
C723 B.n683 VSUBS 0.008287f
C724 B.n684 VSUBS 0.008287f
C725 B.n685 VSUBS 0.008287f
C726 B.n686 VSUBS 0.008287f
C727 B.n687 VSUBS 0.008287f
C728 B.n688 VSUBS 0.008287f
C729 B.n689 VSUBS 0.008287f
C730 B.n690 VSUBS 0.008287f
C731 B.n691 VSUBS 0.008287f
C732 B.n692 VSUBS 0.008287f
C733 B.n693 VSUBS 0.008287f
C734 B.n694 VSUBS 0.008287f
C735 B.n695 VSUBS 0.018765f
C736 VDD2.n0 VSUBS 0.030861f
C737 VDD2.n1 VSUBS 0.027764f
C738 VDD2.n2 VSUBS 0.014919f
C739 VDD2.n3 VSUBS 0.035264f
C740 VDD2.n4 VSUBS 0.015797f
C741 VDD2.n5 VSUBS 0.027764f
C742 VDD2.n6 VSUBS 0.014919f
C743 VDD2.n7 VSUBS 0.035264f
C744 VDD2.n8 VSUBS 0.015797f
C745 VDD2.n9 VSUBS 0.027764f
C746 VDD2.n10 VSUBS 0.014919f
C747 VDD2.n11 VSUBS 0.035264f
C748 VDD2.n12 VSUBS 0.015797f
C749 VDD2.n13 VSUBS 0.027764f
C750 VDD2.n14 VSUBS 0.014919f
C751 VDD2.n15 VSUBS 0.035264f
C752 VDD2.n16 VSUBS 0.015797f
C753 VDD2.n17 VSUBS 0.027764f
C754 VDD2.n18 VSUBS 0.014919f
C755 VDD2.n19 VSUBS 0.035264f
C756 VDD2.n20 VSUBS 0.015797f
C757 VDD2.n21 VSUBS 0.229201f
C758 VDD2.t0 VSUBS 0.076066f
C759 VDD2.n22 VSUBS 0.026448f
C760 VDD2.n23 VSUBS 0.026527f
C761 VDD2.n24 VSUBS 0.014919f
C762 VDD2.n25 VSUBS 1.46632f
C763 VDD2.n26 VSUBS 0.027764f
C764 VDD2.n27 VSUBS 0.014919f
C765 VDD2.n28 VSUBS 0.015797f
C766 VDD2.n29 VSUBS 0.035264f
C767 VDD2.n30 VSUBS 0.035264f
C768 VDD2.n31 VSUBS 0.015797f
C769 VDD2.n32 VSUBS 0.014919f
C770 VDD2.n33 VSUBS 0.027764f
C771 VDD2.n34 VSUBS 0.027764f
C772 VDD2.n35 VSUBS 0.014919f
C773 VDD2.n36 VSUBS 0.015797f
C774 VDD2.n37 VSUBS 0.035264f
C775 VDD2.n38 VSUBS 0.035264f
C776 VDD2.n39 VSUBS 0.035264f
C777 VDD2.n40 VSUBS 0.015797f
C778 VDD2.n41 VSUBS 0.014919f
C779 VDD2.n42 VSUBS 0.027764f
C780 VDD2.n43 VSUBS 0.027764f
C781 VDD2.n44 VSUBS 0.014919f
C782 VDD2.n45 VSUBS 0.015358f
C783 VDD2.n46 VSUBS 0.015358f
C784 VDD2.n47 VSUBS 0.035264f
C785 VDD2.n48 VSUBS 0.035264f
C786 VDD2.n49 VSUBS 0.015797f
C787 VDD2.n50 VSUBS 0.014919f
C788 VDD2.n51 VSUBS 0.027764f
C789 VDD2.n52 VSUBS 0.027764f
C790 VDD2.n53 VSUBS 0.014919f
C791 VDD2.n54 VSUBS 0.015797f
C792 VDD2.n55 VSUBS 0.035264f
C793 VDD2.n56 VSUBS 0.035264f
C794 VDD2.n57 VSUBS 0.015797f
C795 VDD2.n58 VSUBS 0.014919f
C796 VDD2.n59 VSUBS 0.027764f
C797 VDD2.n60 VSUBS 0.027764f
C798 VDD2.n61 VSUBS 0.014919f
C799 VDD2.n62 VSUBS 0.015797f
C800 VDD2.n63 VSUBS 0.035264f
C801 VDD2.n64 VSUBS 0.086577f
C802 VDD2.n65 VSUBS 0.015797f
C803 VDD2.n66 VSUBS 0.014919f
C804 VDD2.n67 VSUBS 0.064175f
C805 VDD2.n68 VSUBS 0.068261f
C806 VDD2.t4 VSUBS 0.281709f
C807 VDD2.t3 VSUBS 0.281709f
C808 VDD2.n69 VSUBS 2.22721f
C809 VDD2.n70 VSUBS 3.0659f
C810 VDD2.n71 VSUBS 0.030861f
C811 VDD2.n72 VSUBS 0.027764f
C812 VDD2.n73 VSUBS 0.014919f
C813 VDD2.n74 VSUBS 0.035264f
C814 VDD2.n75 VSUBS 0.015797f
C815 VDD2.n76 VSUBS 0.027764f
C816 VDD2.n77 VSUBS 0.014919f
C817 VDD2.n78 VSUBS 0.035264f
C818 VDD2.n79 VSUBS 0.015797f
C819 VDD2.n80 VSUBS 0.027764f
C820 VDD2.n81 VSUBS 0.014919f
C821 VDD2.n82 VSUBS 0.035264f
C822 VDD2.n83 VSUBS 0.015797f
C823 VDD2.n84 VSUBS 0.027764f
C824 VDD2.n85 VSUBS 0.014919f
C825 VDD2.n86 VSUBS 0.035264f
C826 VDD2.n87 VSUBS 0.035264f
C827 VDD2.n88 VSUBS 0.015797f
C828 VDD2.n89 VSUBS 0.027764f
C829 VDD2.n90 VSUBS 0.014919f
C830 VDD2.n91 VSUBS 0.035264f
C831 VDD2.n92 VSUBS 0.015797f
C832 VDD2.n93 VSUBS 0.229201f
C833 VDD2.t1 VSUBS 0.076066f
C834 VDD2.n94 VSUBS 0.026448f
C835 VDD2.n95 VSUBS 0.026527f
C836 VDD2.n96 VSUBS 0.014919f
C837 VDD2.n97 VSUBS 1.46632f
C838 VDD2.n98 VSUBS 0.027764f
C839 VDD2.n99 VSUBS 0.014919f
C840 VDD2.n100 VSUBS 0.015797f
C841 VDD2.n101 VSUBS 0.035264f
C842 VDD2.n102 VSUBS 0.035264f
C843 VDD2.n103 VSUBS 0.015797f
C844 VDD2.n104 VSUBS 0.014919f
C845 VDD2.n105 VSUBS 0.027764f
C846 VDD2.n106 VSUBS 0.027764f
C847 VDD2.n107 VSUBS 0.014919f
C848 VDD2.n108 VSUBS 0.015797f
C849 VDD2.n109 VSUBS 0.035264f
C850 VDD2.n110 VSUBS 0.035264f
C851 VDD2.n111 VSUBS 0.015797f
C852 VDD2.n112 VSUBS 0.014919f
C853 VDD2.n113 VSUBS 0.027764f
C854 VDD2.n114 VSUBS 0.027764f
C855 VDD2.n115 VSUBS 0.014919f
C856 VDD2.n116 VSUBS 0.015358f
C857 VDD2.n117 VSUBS 0.015358f
C858 VDD2.n118 VSUBS 0.035264f
C859 VDD2.n119 VSUBS 0.035264f
C860 VDD2.n120 VSUBS 0.015797f
C861 VDD2.n121 VSUBS 0.014919f
C862 VDD2.n122 VSUBS 0.027764f
C863 VDD2.n123 VSUBS 0.027764f
C864 VDD2.n124 VSUBS 0.014919f
C865 VDD2.n125 VSUBS 0.015797f
C866 VDD2.n126 VSUBS 0.035264f
C867 VDD2.n127 VSUBS 0.035264f
C868 VDD2.n128 VSUBS 0.015797f
C869 VDD2.n129 VSUBS 0.014919f
C870 VDD2.n130 VSUBS 0.027764f
C871 VDD2.n131 VSUBS 0.027764f
C872 VDD2.n132 VSUBS 0.014919f
C873 VDD2.n133 VSUBS 0.015797f
C874 VDD2.n134 VSUBS 0.035264f
C875 VDD2.n135 VSUBS 0.086577f
C876 VDD2.n136 VSUBS 0.015797f
C877 VDD2.n137 VSUBS 0.014919f
C878 VDD2.n138 VSUBS 0.064175f
C879 VDD2.n139 VSUBS 0.062763f
C880 VDD2.n140 VSUBS 2.7501f
C881 VDD2.t2 VSUBS 0.281709f
C882 VDD2.t5 VSUBS 0.281709f
C883 VDD2.n141 VSUBS 2.22717f
C884 VN.n0 VSUBS 0.04457f
C885 VN.t2 VSUBS 2.42917f
C886 VN.n1 VSUBS 0.043533f
C887 VN.t5 VSUBS 2.62011f
C888 VN.n2 VSUBS 0.93466f
C889 VN.t1 VSUBS 2.42917f
C890 VN.n3 VSUBS 0.961794f
C891 VN.n4 VSUBS 0.062694f
C892 VN.n5 VSUBS 0.283087f
C893 VN.n6 VSUBS 0.033808f
C894 VN.n7 VSUBS 0.033808f
C895 VN.n8 VSUBS 0.054758f
C896 VN.n9 VSUBS 0.055266f
C897 VN.n10 VSUBS 0.965422f
C898 VN.n11 VSUBS 0.042479f
C899 VN.n12 VSUBS 0.04457f
C900 VN.t4 VSUBS 2.42917f
C901 VN.n13 VSUBS 0.043533f
C902 VN.t0 VSUBS 2.62011f
C903 VN.n14 VSUBS 0.93466f
C904 VN.t3 VSUBS 2.42917f
C905 VN.n15 VSUBS 0.961794f
C906 VN.n16 VSUBS 0.062694f
C907 VN.n17 VSUBS 0.283087f
C908 VN.n18 VSUBS 0.033808f
C909 VN.n19 VSUBS 0.033808f
C910 VN.n20 VSUBS 0.054758f
C911 VN.n21 VSUBS 0.055266f
C912 VN.n22 VSUBS 0.965422f
C913 VN.n23 VSUBS 1.72982f
C914 VTAIL.t2 VSUBS 0.28876f
C915 VTAIL.t4 VSUBS 0.28876f
C916 VTAIL.n0 VSUBS 2.11922f
C917 VTAIL.n1 VSUBS 0.851639f
C918 VTAIL.n2 VSUBS 0.031634f
C919 VTAIL.n3 VSUBS 0.028459f
C920 VTAIL.n4 VSUBS 0.015293f
C921 VTAIL.n5 VSUBS 0.036146f
C922 VTAIL.n6 VSUBS 0.016192f
C923 VTAIL.n7 VSUBS 0.028459f
C924 VTAIL.n8 VSUBS 0.015293f
C925 VTAIL.n9 VSUBS 0.036146f
C926 VTAIL.n10 VSUBS 0.016192f
C927 VTAIL.n11 VSUBS 0.028459f
C928 VTAIL.n12 VSUBS 0.015293f
C929 VTAIL.n13 VSUBS 0.036146f
C930 VTAIL.n14 VSUBS 0.016192f
C931 VTAIL.n15 VSUBS 0.028459f
C932 VTAIL.n16 VSUBS 0.015293f
C933 VTAIL.n17 VSUBS 0.036146f
C934 VTAIL.n18 VSUBS 0.016192f
C935 VTAIL.n19 VSUBS 0.028459f
C936 VTAIL.n20 VSUBS 0.015293f
C937 VTAIL.n21 VSUBS 0.036146f
C938 VTAIL.n22 VSUBS 0.016192f
C939 VTAIL.n23 VSUBS 0.234939f
C940 VTAIL.t9 VSUBS 0.07797f
C941 VTAIL.n24 VSUBS 0.02711f
C942 VTAIL.n25 VSUBS 0.027191f
C943 VTAIL.n26 VSUBS 0.015293f
C944 VTAIL.n27 VSUBS 1.50303f
C945 VTAIL.n28 VSUBS 0.028459f
C946 VTAIL.n29 VSUBS 0.015293f
C947 VTAIL.n30 VSUBS 0.016192f
C948 VTAIL.n31 VSUBS 0.036146f
C949 VTAIL.n32 VSUBS 0.036146f
C950 VTAIL.n33 VSUBS 0.016192f
C951 VTAIL.n34 VSUBS 0.015293f
C952 VTAIL.n35 VSUBS 0.028459f
C953 VTAIL.n36 VSUBS 0.028459f
C954 VTAIL.n37 VSUBS 0.015293f
C955 VTAIL.n38 VSUBS 0.016192f
C956 VTAIL.n39 VSUBS 0.036146f
C957 VTAIL.n40 VSUBS 0.036146f
C958 VTAIL.n41 VSUBS 0.036146f
C959 VTAIL.n42 VSUBS 0.016192f
C960 VTAIL.n43 VSUBS 0.015293f
C961 VTAIL.n44 VSUBS 0.028459f
C962 VTAIL.n45 VSUBS 0.028459f
C963 VTAIL.n46 VSUBS 0.015293f
C964 VTAIL.n47 VSUBS 0.015742f
C965 VTAIL.n48 VSUBS 0.015742f
C966 VTAIL.n49 VSUBS 0.036146f
C967 VTAIL.n50 VSUBS 0.036146f
C968 VTAIL.n51 VSUBS 0.016192f
C969 VTAIL.n52 VSUBS 0.015293f
C970 VTAIL.n53 VSUBS 0.028459f
C971 VTAIL.n54 VSUBS 0.028459f
C972 VTAIL.n55 VSUBS 0.015293f
C973 VTAIL.n56 VSUBS 0.016192f
C974 VTAIL.n57 VSUBS 0.036146f
C975 VTAIL.n58 VSUBS 0.036146f
C976 VTAIL.n59 VSUBS 0.016192f
C977 VTAIL.n60 VSUBS 0.015293f
C978 VTAIL.n61 VSUBS 0.028459f
C979 VTAIL.n62 VSUBS 0.028459f
C980 VTAIL.n63 VSUBS 0.015293f
C981 VTAIL.n64 VSUBS 0.016192f
C982 VTAIL.n65 VSUBS 0.036146f
C983 VTAIL.n66 VSUBS 0.088744f
C984 VTAIL.n67 VSUBS 0.016192f
C985 VTAIL.n68 VSUBS 0.015293f
C986 VTAIL.n69 VSUBS 0.065781f
C987 VTAIL.n70 VSUBS 0.044684f
C988 VTAIL.n71 VSUBS 0.349608f
C989 VTAIL.t7 VSUBS 0.28876f
C990 VTAIL.t6 VSUBS 0.28876f
C991 VTAIL.n72 VSUBS 2.11922f
C992 VTAIL.n73 VSUBS 2.62817f
C993 VTAIL.t3 VSUBS 0.28876f
C994 VTAIL.t1 VSUBS 0.28876f
C995 VTAIL.n74 VSUBS 2.11923f
C996 VTAIL.n75 VSUBS 2.62816f
C997 VTAIL.n76 VSUBS 0.031634f
C998 VTAIL.n77 VSUBS 0.028459f
C999 VTAIL.n78 VSUBS 0.015293f
C1000 VTAIL.n79 VSUBS 0.036146f
C1001 VTAIL.n80 VSUBS 0.016192f
C1002 VTAIL.n81 VSUBS 0.028459f
C1003 VTAIL.n82 VSUBS 0.015293f
C1004 VTAIL.n83 VSUBS 0.036146f
C1005 VTAIL.n84 VSUBS 0.016192f
C1006 VTAIL.n85 VSUBS 0.028459f
C1007 VTAIL.n86 VSUBS 0.015293f
C1008 VTAIL.n87 VSUBS 0.036146f
C1009 VTAIL.n88 VSUBS 0.016192f
C1010 VTAIL.n89 VSUBS 0.028459f
C1011 VTAIL.n90 VSUBS 0.015293f
C1012 VTAIL.n91 VSUBS 0.036146f
C1013 VTAIL.n92 VSUBS 0.036146f
C1014 VTAIL.n93 VSUBS 0.016192f
C1015 VTAIL.n94 VSUBS 0.028459f
C1016 VTAIL.n95 VSUBS 0.015293f
C1017 VTAIL.n96 VSUBS 0.036146f
C1018 VTAIL.n97 VSUBS 0.016192f
C1019 VTAIL.n98 VSUBS 0.234939f
C1020 VTAIL.t0 VSUBS 0.07797f
C1021 VTAIL.n99 VSUBS 0.02711f
C1022 VTAIL.n100 VSUBS 0.027191f
C1023 VTAIL.n101 VSUBS 0.015293f
C1024 VTAIL.n102 VSUBS 1.50303f
C1025 VTAIL.n103 VSUBS 0.028459f
C1026 VTAIL.n104 VSUBS 0.015293f
C1027 VTAIL.n105 VSUBS 0.016192f
C1028 VTAIL.n106 VSUBS 0.036146f
C1029 VTAIL.n107 VSUBS 0.036146f
C1030 VTAIL.n108 VSUBS 0.016192f
C1031 VTAIL.n109 VSUBS 0.015293f
C1032 VTAIL.n110 VSUBS 0.028459f
C1033 VTAIL.n111 VSUBS 0.028459f
C1034 VTAIL.n112 VSUBS 0.015293f
C1035 VTAIL.n113 VSUBS 0.016192f
C1036 VTAIL.n114 VSUBS 0.036146f
C1037 VTAIL.n115 VSUBS 0.036146f
C1038 VTAIL.n116 VSUBS 0.016192f
C1039 VTAIL.n117 VSUBS 0.015293f
C1040 VTAIL.n118 VSUBS 0.028459f
C1041 VTAIL.n119 VSUBS 0.028459f
C1042 VTAIL.n120 VSUBS 0.015293f
C1043 VTAIL.n121 VSUBS 0.015742f
C1044 VTAIL.n122 VSUBS 0.015742f
C1045 VTAIL.n123 VSUBS 0.036146f
C1046 VTAIL.n124 VSUBS 0.036146f
C1047 VTAIL.n125 VSUBS 0.016192f
C1048 VTAIL.n126 VSUBS 0.015293f
C1049 VTAIL.n127 VSUBS 0.028459f
C1050 VTAIL.n128 VSUBS 0.028459f
C1051 VTAIL.n129 VSUBS 0.015293f
C1052 VTAIL.n130 VSUBS 0.016192f
C1053 VTAIL.n131 VSUBS 0.036146f
C1054 VTAIL.n132 VSUBS 0.036146f
C1055 VTAIL.n133 VSUBS 0.016192f
C1056 VTAIL.n134 VSUBS 0.015293f
C1057 VTAIL.n135 VSUBS 0.028459f
C1058 VTAIL.n136 VSUBS 0.028459f
C1059 VTAIL.n137 VSUBS 0.015293f
C1060 VTAIL.n138 VSUBS 0.016192f
C1061 VTAIL.n139 VSUBS 0.036146f
C1062 VTAIL.n140 VSUBS 0.088744f
C1063 VTAIL.n141 VSUBS 0.016192f
C1064 VTAIL.n142 VSUBS 0.015293f
C1065 VTAIL.n143 VSUBS 0.065781f
C1066 VTAIL.n144 VSUBS 0.044684f
C1067 VTAIL.n145 VSUBS 0.349608f
C1068 VTAIL.t5 VSUBS 0.28876f
C1069 VTAIL.t10 VSUBS 0.28876f
C1070 VTAIL.n146 VSUBS 2.11923f
C1071 VTAIL.n147 VSUBS 0.987403f
C1072 VTAIL.n148 VSUBS 0.031634f
C1073 VTAIL.n149 VSUBS 0.028459f
C1074 VTAIL.n150 VSUBS 0.015293f
C1075 VTAIL.n151 VSUBS 0.036146f
C1076 VTAIL.n152 VSUBS 0.016192f
C1077 VTAIL.n153 VSUBS 0.028459f
C1078 VTAIL.n154 VSUBS 0.015293f
C1079 VTAIL.n155 VSUBS 0.036146f
C1080 VTAIL.n156 VSUBS 0.016192f
C1081 VTAIL.n157 VSUBS 0.028459f
C1082 VTAIL.n158 VSUBS 0.015293f
C1083 VTAIL.n159 VSUBS 0.036146f
C1084 VTAIL.n160 VSUBS 0.016192f
C1085 VTAIL.n161 VSUBS 0.028459f
C1086 VTAIL.n162 VSUBS 0.015293f
C1087 VTAIL.n163 VSUBS 0.036146f
C1088 VTAIL.n164 VSUBS 0.036146f
C1089 VTAIL.n165 VSUBS 0.016192f
C1090 VTAIL.n166 VSUBS 0.028459f
C1091 VTAIL.n167 VSUBS 0.015293f
C1092 VTAIL.n168 VSUBS 0.036146f
C1093 VTAIL.n169 VSUBS 0.016192f
C1094 VTAIL.n170 VSUBS 0.234939f
C1095 VTAIL.t8 VSUBS 0.07797f
C1096 VTAIL.n171 VSUBS 0.02711f
C1097 VTAIL.n172 VSUBS 0.027191f
C1098 VTAIL.n173 VSUBS 0.015293f
C1099 VTAIL.n174 VSUBS 1.50303f
C1100 VTAIL.n175 VSUBS 0.028459f
C1101 VTAIL.n176 VSUBS 0.015293f
C1102 VTAIL.n177 VSUBS 0.016192f
C1103 VTAIL.n178 VSUBS 0.036146f
C1104 VTAIL.n179 VSUBS 0.036146f
C1105 VTAIL.n180 VSUBS 0.016192f
C1106 VTAIL.n181 VSUBS 0.015293f
C1107 VTAIL.n182 VSUBS 0.028459f
C1108 VTAIL.n183 VSUBS 0.028459f
C1109 VTAIL.n184 VSUBS 0.015293f
C1110 VTAIL.n185 VSUBS 0.016192f
C1111 VTAIL.n186 VSUBS 0.036146f
C1112 VTAIL.n187 VSUBS 0.036146f
C1113 VTAIL.n188 VSUBS 0.016192f
C1114 VTAIL.n189 VSUBS 0.015293f
C1115 VTAIL.n190 VSUBS 0.028459f
C1116 VTAIL.n191 VSUBS 0.028459f
C1117 VTAIL.n192 VSUBS 0.015293f
C1118 VTAIL.n193 VSUBS 0.015742f
C1119 VTAIL.n194 VSUBS 0.015742f
C1120 VTAIL.n195 VSUBS 0.036146f
C1121 VTAIL.n196 VSUBS 0.036146f
C1122 VTAIL.n197 VSUBS 0.016192f
C1123 VTAIL.n198 VSUBS 0.015293f
C1124 VTAIL.n199 VSUBS 0.028459f
C1125 VTAIL.n200 VSUBS 0.028459f
C1126 VTAIL.n201 VSUBS 0.015293f
C1127 VTAIL.n202 VSUBS 0.016192f
C1128 VTAIL.n203 VSUBS 0.036146f
C1129 VTAIL.n204 VSUBS 0.036146f
C1130 VTAIL.n205 VSUBS 0.016192f
C1131 VTAIL.n206 VSUBS 0.015293f
C1132 VTAIL.n207 VSUBS 0.028459f
C1133 VTAIL.n208 VSUBS 0.028459f
C1134 VTAIL.n209 VSUBS 0.015293f
C1135 VTAIL.n210 VSUBS 0.016192f
C1136 VTAIL.n211 VSUBS 0.036146f
C1137 VTAIL.n212 VSUBS 0.088744f
C1138 VTAIL.n213 VSUBS 0.016192f
C1139 VTAIL.n214 VSUBS 0.015293f
C1140 VTAIL.n215 VSUBS 0.065781f
C1141 VTAIL.n216 VSUBS 0.044684f
C1142 VTAIL.n217 VSUBS 1.80222f
C1143 VTAIL.n218 VSUBS 0.031634f
C1144 VTAIL.n219 VSUBS 0.028459f
C1145 VTAIL.n220 VSUBS 0.015293f
C1146 VTAIL.n221 VSUBS 0.036146f
C1147 VTAIL.n222 VSUBS 0.016192f
C1148 VTAIL.n223 VSUBS 0.028459f
C1149 VTAIL.n224 VSUBS 0.015293f
C1150 VTAIL.n225 VSUBS 0.036146f
C1151 VTAIL.n226 VSUBS 0.016192f
C1152 VTAIL.n227 VSUBS 0.028459f
C1153 VTAIL.n228 VSUBS 0.015293f
C1154 VTAIL.n229 VSUBS 0.036146f
C1155 VTAIL.n230 VSUBS 0.016192f
C1156 VTAIL.n231 VSUBS 0.028459f
C1157 VTAIL.n232 VSUBS 0.015293f
C1158 VTAIL.n233 VSUBS 0.036146f
C1159 VTAIL.n234 VSUBS 0.016192f
C1160 VTAIL.n235 VSUBS 0.028459f
C1161 VTAIL.n236 VSUBS 0.015293f
C1162 VTAIL.n237 VSUBS 0.036146f
C1163 VTAIL.n238 VSUBS 0.016192f
C1164 VTAIL.n239 VSUBS 0.234939f
C1165 VTAIL.t11 VSUBS 0.07797f
C1166 VTAIL.n240 VSUBS 0.02711f
C1167 VTAIL.n241 VSUBS 0.027191f
C1168 VTAIL.n242 VSUBS 0.015293f
C1169 VTAIL.n243 VSUBS 1.50303f
C1170 VTAIL.n244 VSUBS 0.028459f
C1171 VTAIL.n245 VSUBS 0.015293f
C1172 VTAIL.n246 VSUBS 0.016192f
C1173 VTAIL.n247 VSUBS 0.036146f
C1174 VTAIL.n248 VSUBS 0.036146f
C1175 VTAIL.n249 VSUBS 0.016192f
C1176 VTAIL.n250 VSUBS 0.015293f
C1177 VTAIL.n251 VSUBS 0.028459f
C1178 VTAIL.n252 VSUBS 0.028459f
C1179 VTAIL.n253 VSUBS 0.015293f
C1180 VTAIL.n254 VSUBS 0.016192f
C1181 VTAIL.n255 VSUBS 0.036146f
C1182 VTAIL.n256 VSUBS 0.036146f
C1183 VTAIL.n257 VSUBS 0.036146f
C1184 VTAIL.n258 VSUBS 0.016192f
C1185 VTAIL.n259 VSUBS 0.015293f
C1186 VTAIL.n260 VSUBS 0.028459f
C1187 VTAIL.n261 VSUBS 0.028459f
C1188 VTAIL.n262 VSUBS 0.015293f
C1189 VTAIL.n263 VSUBS 0.015742f
C1190 VTAIL.n264 VSUBS 0.015742f
C1191 VTAIL.n265 VSUBS 0.036146f
C1192 VTAIL.n266 VSUBS 0.036146f
C1193 VTAIL.n267 VSUBS 0.016192f
C1194 VTAIL.n268 VSUBS 0.015293f
C1195 VTAIL.n269 VSUBS 0.028459f
C1196 VTAIL.n270 VSUBS 0.028459f
C1197 VTAIL.n271 VSUBS 0.015293f
C1198 VTAIL.n272 VSUBS 0.016192f
C1199 VTAIL.n273 VSUBS 0.036146f
C1200 VTAIL.n274 VSUBS 0.036146f
C1201 VTAIL.n275 VSUBS 0.016192f
C1202 VTAIL.n276 VSUBS 0.015293f
C1203 VTAIL.n277 VSUBS 0.028459f
C1204 VTAIL.n278 VSUBS 0.028459f
C1205 VTAIL.n279 VSUBS 0.015293f
C1206 VTAIL.n280 VSUBS 0.016192f
C1207 VTAIL.n281 VSUBS 0.036146f
C1208 VTAIL.n282 VSUBS 0.088744f
C1209 VTAIL.n283 VSUBS 0.016192f
C1210 VTAIL.n284 VSUBS 0.015293f
C1211 VTAIL.n285 VSUBS 0.065781f
C1212 VTAIL.n286 VSUBS 0.044684f
C1213 VTAIL.n287 VSUBS 1.74984f
C1214 VDD1.n0 VSUBS 0.030857f
C1215 VDD1.n1 VSUBS 0.02776f
C1216 VDD1.n2 VSUBS 0.014917f
C1217 VDD1.n3 VSUBS 0.035259f
C1218 VDD1.n4 VSUBS 0.015795f
C1219 VDD1.n5 VSUBS 0.02776f
C1220 VDD1.n6 VSUBS 0.014917f
C1221 VDD1.n7 VSUBS 0.035259f
C1222 VDD1.n8 VSUBS 0.015795f
C1223 VDD1.n9 VSUBS 0.02776f
C1224 VDD1.n10 VSUBS 0.014917f
C1225 VDD1.n11 VSUBS 0.035259f
C1226 VDD1.n12 VSUBS 0.015795f
C1227 VDD1.n13 VSUBS 0.02776f
C1228 VDD1.n14 VSUBS 0.014917f
C1229 VDD1.n15 VSUBS 0.035259f
C1230 VDD1.n16 VSUBS 0.035259f
C1231 VDD1.n17 VSUBS 0.015795f
C1232 VDD1.n18 VSUBS 0.02776f
C1233 VDD1.n19 VSUBS 0.014917f
C1234 VDD1.n20 VSUBS 0.035259f
C1235 VDD1.n21 VSUBS 0.015795f
C1236 VDD1.n22 VSUBS 0.229171f
C1237 VDD1.t5 VSUBS 0.076056f
C1238 VDD1.n23 VSUBS 0.026444f
C1239 VDD1.n24 VSUBS 0.026524f
C1240 VDD1.n25 VSUBS 0.014917f
C1241 VDD1.n26 VSUBS 1.46613f
C1242 VDD1.n27 VSUBS 0.02776f
C1243 VDD1.n28 VSUBS 0.014917f
C1244 VDD1.n29 VSUBS 0.015795f
C1245 VDD1.n30 VSUBS 0.035259f
C1246 VDD1.n31 VSUBS 0.035259f
C1247 VDD1.n32 VSUBS 0.015795f
C1248 VDD1.n33 VSUBS 0.014917f
C1249 VDD1.n34 VSUBS 0.02776f
C1250 VDD1.n35 VSUBS 0.02776f
C1251 VDD1.n36 VSUBS 0.014917f
C1252 VDD1.n37 VSUBS 0.015795f
C1253 VDD1.n38 VSUBS 0.035259f
C1254 VDD1.n39 VSUBS 0.035259f
C1255 VDD1.n40 VSUBS 0.015795f
C1256 VDD1.n41 VSUBS 0.014917f
C1257 VDD1.n42 VSUBS 0.02776f
C1258 VDD1.n43 VSUBS 0.02776f
C1259 VDD1.n44 VSUBS 0.014917f
C1260 VDD1.n45 VSUBS 0.015356f
C1261 VDD1.n46 VSUBS 0.015356f
C1262 VDD1.n47 VSUBS 0.035259f
C1263 VDD1.n48 VSUBS 0.035259f
C1264 VDD1.n49 VSUBS 0.015795f
C1265 VDD1.n50 VSUBS 0.014917f
C1266 VDD1.n51 VSUBS 0.02776f
C1267 VDD1.n52 VSUBS 0.02776f
C1268 VDD1.n53 VSUBS 0.014917f
C1269 VDD1.n54 VSUBS 0.015795f
C1270 VDD1.n55 VSUBS 0.035259f
C1271 VDD1.n56 VSUBS 0.035259f
C1272 VDD1.n57 VSUBS 0.015795f
C1273 VDD1.n58 VSUBS 0.014917f
C1274 VDD1.n59 VSUBS 0.02776f
C1275 VDD1.n60 VSUBS 0.02776f
C1276 VDD1.n61 VSUBS 0.014917f
C1277 VDD1.n62 VSUBS 0.015795f
C1278 VDD1.n63 VSUBS 0.035259f
C1279 VDD1.n64 VSUBS 0.086566f
C1280 VDD1.n65 VSUBS 0.015795f
C1281 VDD1.n66 VSUBS 0.014917f
C1282 VDD1.n67 VSUBS 0.064167f
C1283 VDD1.n68 VSUBS 0.068967f
C1284 VDD1.n69 VSUBS 0.030857f
C1285 VDD1.n70 VSUBS 0.02776f
C1286 VDD1.n71 VSUBS 0.014917f
C1287 VDD1.n72 VSUBS 0.035259f
C1288 VDD1.n73 VSUBS 0.015795f
C1289 VDD1.n74 VSUBS 0.02776f
C1290 VDD1.n75 VSUBS 0.014917f
C1291 VDD1.n76 VSUBS 0.035259f
C1292 VDD1.n77 VSUBS 0.015795f
C1293 VDD1.n78 VSUBS 0.02776f
C1294 VDD1.n79 VSUBS 0.014917f
C1295 VDD1.n80 VSUBS 0.035259f
C1296 VDD1.n81 VSUBS 0.015795f
C1297 VDD1.n82 VSUBS 0.02776f
C1298 VDD1.n83 VSUBS 0.014917f
C1299 VDD1.n84 VSUBS 0.035259f
C1300 VDD1.n85 VSUBS 0.015795f
C1301 VDD1.n86 VSUBS 0.02776f
C1302 VDD1.n87 VSUBS 0.014917f
C1303 VDD1.n88 VSUBS 0.035259f
C1304 VDD1.n89 VSUBS 0.015795f
C1305 VDD1.n90 VSUBS 0.229171f
C1306 VDD1.t2 VSUBS 0.076056f
C1307 VDD1.n91 VSUBS 0.026444f
C1308 VDD1.n92 VSUBS 0.026524f
C1309 VDD1.n93 VSUBS 0.014917f
C1310 VDD1.n94 VSUBS 1.46613f
C1311 VDD1.n95 VSUBS 0.02776f
C1312 VDD1.n96 VSUBS 0.014917f
C1313 VDD1.n97 VSUBS 0.015795f
C1314 VDD1.n98 VSUBS 0.035259f
C1315 VDD1.n99 VSUBS 0.035259f
C1316 VDD1.n100 VSUBS 0.015795f
C1317 VDD1.n101 VSUBS 0.014917f
C1318 VDD1.n102 VSUBS 0.02776f
C1319 VDD1.n103 VSUBS 0.02776f
C1320 VDD1.n104 VSUBS 0.014917f
C1321 VDD1.n105 VSUBS 0.015795f
C1322 VDD1.n106 VSUBS 0.035259f
C1323 VDD1.n107 VSUBS 0.035259f
C1324 VDD1.n108 VSUBS 0.035259f
C1325 VDD1.n109 VSUBS 0.015795f
C1326 VDD1.n110 VSUBS 0.014917f
C1327 VDD1.n111 VSUBS 0.02776f
C1328 VDD1.n112 VSUBS 0.02776f
C1329 VDD1.n113 VSUBS 0.014917f
C1330 VDD1.n114 VSUBS 0.015356f
C1331 VDD1.n115 VSUBS 0.015356f
C1332 VDD1.n116 VSUBS 0.035259f
C1333 VDD1.n117 VSUBS 0.035259f
C1334 VDD1.n118 VSUBS 0.015795f
C1335 VDD1.n119 VSUBS 0.014917f
C1336 VDD1.n120 VSUBS 0.02776f
C1337 VDD1.n121 VSUBS 0.02776f
C1338 VDD1.n122 VSUBS 0.014917f
C1339 VDD1.n123 VSUBS 0.015795f
C1340 VDD1.n124 VSUBS 0.035259f
C1341 VDD1.n125 VSUBS 0.035259f
C1342 VDD1.n126 VSUBS 0.015795f
C1343 VDD1.n127 VSUBS 0.014917f
C1344 VDD1.n128 VSUBS 0.02776f
C1345 VDD1.n129 VSUBS 0.02776f
C1346 VDD1.n130 VSUBS 0.014917f
C1347 VDD1.n131 VSUBS 0.015795f
C1348 VDD1.n132 VSUBS 0.035259f
C1349 VDD1.n133 VSUBS 0.086566f
C1350 VDD1.n134 VSUBS 0.015795f
C1351 VDD1.n135 VSUBS 0.014917f
C1352 VDD1.n136 VSUBS 0.064167f
C1353 VDD1.n137 VSUBS 0.068252f
C1354 VDD1.t0 VSUBS 0.281672f
C1355 VDD1.t4 VSUBS 0.281672f
C1356 VDD1.n138 VSUBS 2.22692f
C1357 VDD1.n139 VSUBS 3.18824f
C1358 VDD1.t3 VSUBS 0.281672f
C1359 VDD1.t1 VSUBS 0.281672f
C1360 VDD1.n140 VSUBS 2.22215f
C1361 VDD1.n141 VSUBS 3.29725f
C1362 VP.n0 VSUBS 0.045884f
C1363 VP.t1 VSUBS 2.50079f
C1364 VP.n1 VSUBS 0.044817f
C1365 VP.n2 VSUBS 0.034805f
C1366 VP.t4 VSUBS 2.50079f
C1367 VP.n3 VSUBS 0.044817f
C1368 VP.n4 VSUBS 0.045884f
C1369 VP.t3 VSUBS 2.50079f
C1370 VP.n5 VSUBS 0.045884f
C1371 VP.t2 VSUBS 2.50079f
C1372 VP.n6 VSUBS 0.044817f
C1373 VP.t5 VSUBS 2.69736f
C1374 VP.n7 VSUBS 0.962218f
C1375 VP.t0 VSUBS 2.50079f
C1376 VP.n8 VSUBS 0.990153f
C1377 VP.n9 VSUBS 0.064543f
C1378 VP.n10 VSUBS 0.291434f
C1379 VP.n11 VSUBS 0.034805f
C1380 VP.n12 VSUBS 0.034805f
C1381 VP.n13 VSUBS 0.056372f
C1382 VP.n14 VSUBS 0.056896f
C1383 VP.n15 VSUBS 0.993887f
C1384 VP.n16 VSUBS 1.76194f
C1385 VP.n17 VSUBS 1.78854f
C1386 VP.n18 VSUBS 0.993887f
C1387 VP.n19 VSUBS 0.056896f
C1388 VP.n20 VSUBS 0.056372f
C1389 VP.n21 VSUBS 0.034805f
C1390 VP.n22 VSUBS 0.034805f
C1391 VP.n23 VSUBS 0.034805f
C1392 VP.n24 VSUBS 0.064543f
C1393 VP.n25 VSUBS 0.920357f
C1394 VP.n26 VSUBS 0.064543f
C1395 VP.n27 VSUBS 0.034805f
C1396 VP.n28 VSUBS 0.034805f
C1397 VP.n29 VSUBS 0.034805f
C1398 VP.n30 VSUBS 0.056372f
C1399 VP.n31 VSUBS 0.056896f
C1400 VP.n32 VSUBS 0.993887f
C1401 VP.n33 VSUBS 0.043731f
.ends

