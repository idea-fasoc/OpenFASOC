* NGSPICE file created from diff_pair_sample_1282.ext - technology: sky130A

.subckt diff_pair_sample_1282 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0 ps=0 w=5.9 l=2
X1 VDD2.t5 VN.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0.9735 ps=6.23 w=5.9 l=2
X2 VDD1.t5 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=2.301 ps=12.58 w=5.9 l=2
X3 VDD1.t4 VP.t1 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=2.301 ps=12.58 w=5.9 l=2
X4 VTAIL.t7 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=0.9735 ps=6.23 w=5.9 l=2
X5 VDD1.t3 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0.9735 ps=6.23 w=5.9 l=2
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0 ps=0 w=5.9 l=2
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0 ps=0 w=5.9 l=2
X8 VDD2.t3 VN.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0.9735 ps=6.23 w=5.9 l=2
X9 VDD2.t2 VN.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=2.301 ps=12.58 w=5.9 l=2
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0 ps=0 w=5.9 l=2
X11 VTAIL.t8 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=0.9735 ps=6.23 w=5.9 l=2
X12 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.301 pd=12.58 as=0.9735 ps=6.23 w=5.9 l=2
X13 VTAIL.t0 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=0.9735 ps=6.23 w=5.9 l=2
X14 VTAIL.t3 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=0.9735 ps=6.23 w=5.9 l=2
X15 VDD2.t0 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9735 pd=6.23 as=2.301 ps=12.58 w=5.9 l=2
R0 B.n579 B.n578 585
R1 B.n580 B.n579 585
R2 B.n210 B.n96 585
R3 B.n209 B.n208 585
R4 B.n207 B.n206 585
R5 B.n205 B.n204 585
R6 B.n203 B.n202 585
R7 B.n201 B.n200 585
R8 B.n199 B.n198 585
R9 B.n197 B.n196 585
R10 B.n195 B.n194 585
R11 B.n193 B.n192 585
R12 B.n191 B.n190 585
R13 B.n189 B.n188 585
R14 B.n187 B.n186 585
R15 B.n185 B.n184 585
R16 B.n183 B.n182 585
R17 B.n181 B.n180 585
R18 B.n179 B.n178 585
R19 B.n177 B.n176 585
R20 B.n175 B.n174 585
R21 B.n173 B.n172 585
R22 B.n171 B.n170 585
R23 B.n169 B.n168 585
R24 B.n167 B.n166 585
R25 B.n164 B.n163 585
R26 B.n162 B.n161 585
R27 B.n160 B.n159 585
R28 B.n158 B.n157 585
R29 B.n156 B.n155 585
R30 B.n154 B.n153 585
R31 B.n152 B.n151 585
R32 B.n150 B.n149 585
R33 B.n148 B.n147 585
R34 B.n146 B.n145 585
R35 B.n144 B.n143 585
R36 B.n142 B.n141 585
R37 B.n140 B.n139 585
R38 B.n138 B.n137 585
R39 B.n136 B.n135 585
R40 B.n134 B.n133 585
R41 B.n132 B.n131 585
R42 B.n130 B.n129 585
R43 B.n128 B.n127 585
R44 B.n126 B.n125 585
R45 B.n124 B.n123 585
R46 B.n122 B.n121 585
R47 B.n120 B.n119 585
R48 B.n118 B.n117 585
R49 B.n116 B.n115 585
R50 B.n114 B.n113 585
R51 B.n112 B.n111 585
R52 B.n110 B.n109 585
R53 B.n108 B.n107 585
R54 B.n106 B.n105 585
R55 B.n104 B.n103 585
R56 B.n68 B.n67 585
R57 B.n583 B.n582 585
R58 B.n577 B.n97 585
R59 B.n97 B.n65 585
R60 B.n576 B.n64 585
R61 B.n587 B.n64 585
R62 B.n575 B.n63 585
R63 B.n588 B.n63 585
R64 B.n574 B.n62 585
R65 B.n589 B.n62 585
R66 B.n573 B.n572 585
R67 B.n572 B.n58 585
R68 B.n571 B.n57 585
R69 B.n595 B.n57 585
R70 B.n570 B.n56 585
R71 B.n596 B.n56 585
R72 B.n569 B.n55 585
R73 B.n597 B.n55 585
R74 B.n568 B.n567 585
R75 B.n567 B.n51 585
R76 B.n566 B.n50 585
R77 B.n603 B.n50 585
R78 B.n565 B.n49 585
R79 B.n604 B.n49 585
R80 B.n564 B.n48 585
R81 B.n605 B.n48 585
R82 B.n563 B.n562 585
R83 B.n562 B.n44 585
R84 B.n561 B.n43 585
R85 B.n611 B.n43 585
R86 B.n560 B.n42 585
R87 B.n612 B.n42 585
R88 B.n559 B.n41 585
R89 B.n613 B.n41 585
R90 B.n558 B.n557 585
R91 B.n557 B.n40 585
R92 B.n556 B.n36 585
R93 B.n619 B.n36 585
R94 B.n555 B.n35 585
R95 B.n620 B.n35 585
R96 B.n554 B.n34 585
R97 B.n621 B.n34 585
R98 B.n553 B.n552 585
R99 B.n552 B.n30 585
R100 B.n551 B.n29 585
R101 B.n627 B.n29 585
R102 B.n550 B.n28 585
R103 B.n628 B.n28 585
R104 B.n549 B.n27 585
R105 B.n629 B.n27 585
R106 B.n548 B.n547 585
R107 B.n547 B.n23 585
R108 B.n546 B.n22 585
R109 B.n635 B.n22 585
R110 B.n545 B.n21 585
R111 B.n636 B.n21 585
R112 B.n544 B.n20 585
R113 B.n637 B.n20 585
R114 B.n543 B.n542 585
R115 B.n542 B.n16 585
R116 B.n541 B.n15 585
R117 B.n643 B.n15 585
R118 B.n540 B.n14 585
R119 B.n644 B.n14 585
R120 B.n539 B.n13 585
R121 B.n645 B.n13 585
R122 B.n538 B.n537 585
R123 B.n537 B.n12 585
R124 B.n536 B.n535 585
R125 B.n536 B.n8 585
R126 B.n534 B.n7 585
R127 B.n652 B.n7 585
R128 B.n533 B.n6 585
R129 B.n653 B.n6 585
R130 B.n532 B.n5 585
R131 B.n654 B.n5 585
R132 B.n531 B.n530 585
R133 B.n530 B.n4 585
R134 B.n529 B.n211 585
R135 B.n529 B.n528 585
R136 B.n519 B.n212 585
R137 B.n213 B.n212 585
R138 B.n521 B.n520 585
R139 B.n522 B.n521 585
R140 B.n518 B.n217 585
R141 B.n221 B.n217 585
R142 B.n517 B.n516 585
R143 B.n516 B.n515 585
R144 B.n219 B.n218 585
R145 B.n220 B.n219 585
R146 B.n508 B.n507 585
R147 B.n509 B.n508 585
R148 B.n506 B.n226 585
R149 B.n226 B.n225 585
R150 B.n505 B.n504 585
R151 B.n504 B.n503 585
R152 B.n228 B.n227 585
R153 B.n229 B.n228 585
R154 B.n496 B.n495 585
R155 B.n497 B.n496 585
R156 B.n494 B.n234 585
R157 B.n234 B.n233 585
R158 B.n493 B.n492 585
R159 B.n492 B.n491 585
R160 B.n236 B.n235 585
R161 B.n237 B.n236 585
R162 B.n484 B.n483 585
R163 B.n485 B.n484 585
R164 B.n482 B.n242 585
R165 B.n242 B.n241 585
R166 B.n481 B.n480 585
R167 B.n480 B.n479 585
R168 B.n244 B.n243 585
R169 B.n472 B.n244 585
R170 B.n471 B.n470 585
R171 B.n473 B.n471 585
R172 B.n469 B.n249 585
R173 B.n249 B.n248 585
R174 B.n468 B.n467 585
R175 B.n467 B.n466 585
R176 B.n251 B.n250 585
R177 B.n252 B.n251 585
R178 B.n459 B.n458 585
R179 B.n460 B.n459 585
R180 B.n457 B.n257 585
R181 B.n257 B.n256 585
R182 B.n456 B.n455 585
R183 B.n455 B.n454 585
R184 B.n259 B.n258 585
R185 B.n260 B.n259 585
R186 B.n447 B.n446 585
R187 B.n448 B.n447 585
R188 B.n445 B.n264 585
R189 B.n268 B.n264 585
R190 B.n444 B.n443 585
R191 B.n443 B.n442 585
R192 B.n266 B.n265 585
R193 B.n267 B.n266 585
R194 B.n435 B.n434 585
R195 B.n436 B.n435 585
R196 B.n433 B.n273 585
R197 B.n273 B.n272 585
R198 B.n432 B.n431 585
R199 B.n431 B.n430 585
R200 B.n275 B.n274 585
R201 B.n276 B.n275 585
R202 B.n426 B.n425 585
R203 B.n279 B.n278 585
R204 B.n422 B.n421 585
R205 B.n423 B.n422 585
R206 B.n420 B.n307 585
R207 B.n419 B.n418 585
R208 B.n417 B.n416 585
R209 B.n415 B.n414 585
R210 B.n413 B.n412 585
R211 B.n411 B.n410 585
R212 B.n409 B.n408 585
R213 B.n407 B.n406 585
R214 B.n405 B.n404 585
R215 B.n403 B.n402 585
R216 B.n401 B.n400 585
R217 B.n399 B.n398 585
R218 B.n397 B.n396 585
R219 B.n395 B.n394 585
R220 B.n393 B.n392 585
R221 B.n391 B.n390 585
R222 B.n389 B.n388 585
R223 B.n387 B.n386 585
R224 B.n385 B.n384 585
R225 B.n383 B.n382 585
R226 B.n381 B.n380 585
R227 B.n378 B.n377 585
R228 B.n376 B.n375 585
R229 B.n374 B.n373 585
R230 B.n372 B.n371 585
R231 B.n370 B.n369 585
R232 B.n368 B.n367 585
R233 B.n366 B.n365 585
R234 B.n364 B.n363 585
R235 B.n362 B.n361 585
R236 B.n360 B.n359 585
R237 B.n358 B.n357 585
R238 B.n356 B.n355 585
R239 B.n354 B.n353 585
R240 B.n352 B.n351 585
R241 B.n350 B.n349 585
R242 B.n348 B.n347 585
R243 B.n346 B.n345 585
R244 B.n344 B.n343 585
R245 B.n342 B.n341 585
R246 B.n340 B.n339 585
R247 B.n338 B.n337 585
R248 B.n336 B.n335 585
R249 B.n334 B.n333 585
R250 B.n332 B.n331 585
R251 B.n330 B.n329 585
R252 B.n328 B.n327 585
R253 B.n326 B.n325 585
R254 B.n324 B.n323 585
R255 B.n322 B.n321 585
R256 B.n320 B.n319 585
R257 B.n318 B.n317 585
R258 B.n316 B.n315 585
R259 B.n314 B.n313 585
R260 B.n427 B.n277 585
R261 B.n277 B.n276 585
R262 B.n429 B.n428 585
R263 B.n430 B.n429 585
R264 B.n271 B.n270 585
R265 B.n272 B.n271 585
R266 B.n438 B.n437 585
R267 B.n437 B.n436 585
R268 B.n439 B.n269 585
R269 B.n269 B.n267 585
R270 B.n441 B.n440 585
R271 B.n442 B.n441 585
R272 B.n263 B.n262 585
R273 B.n268 B.n263 585
R274 B.n450 B.n449 585
R275 B.n449 B.n448 585
R276 B.n451 B.n261 585
R277 B.n261 B.n260 585
R278 B.n453 B.n452 585
R279 B.n454 B.n453 585
R280 B.n255 B.n254 585
R281 B.n256 B.n255 585
R282 B.n462 B.n461 585
R283 B.n461 B.n460 585
R284 B.n463 B.n253 585
R285 B.n253 B.n252 585
R286 B.n465 B.n464 585
R287 B.n466 B.n465 585
R288 B.n247 B.n246 585
R289 B.n248 B.n247 585
R290 B.n475 B.n474 585
R291 B.n474 B.n473 585
R292 B.n476 B.n245 585
R293 B.n472 B.n245 585
R294 B.n478 B.n477 585
R295 B.n479 B.n478 585
R296 B.n240 B.n239 585
R297 B.n241 B.n240 585
R298 B.n487 B.n486 585
R299 B.n486 B.n485 585
R300 B.n488 B.n238 585
R301 B.n238 B.n237 585
R302 B.n490 B.n489 585
R303 B.n491 B.n490 585
R304 B.n232 B.n231 585
R305 B.n233 B.n232 585
R306 B.n499 B.n498 585
R307 B.n498 B.n497 585
R308 B.n500 B.n230 585
R309 B.n230 B.n229 585
R310 B.n502 B.n501 585
R311 B.n503 B.n502 585
R312 B.n224 B.n223 585
R313 B.n225 B.n224 585
R314 B.n511 B.n510 585
R315 B.n510 B.n509 585
R316 B.n512 B.n222 585
R317 B.n222 B.n220 585
R318 B.n514 B.n513 585
R319 B.n515 B.n514 585
R320 B.n216 B.n215 585
R321 B.n221 B.n216 585
R322 B.n524 B.n523 585
R323 B.n523 B.n522 585
R324 B.n525 B.n214 585
R325 B.n214 B.n213 585
R326 B.n527 B.n526 585
R327 B.n528 B.n527 585
R328 B.n3 B.n0 585
R329 B.n4 B.n3 585
R330 B.n651 B.n1 585
R331 B.n652 B.n651 585
R332 B.n650 B.n649 585
R333 B.n650 B.n8 585
R334 B.n648 B.n9 585
R335 B.n12 B.n9 585
R336 B.n647 B.n646 585
R337 B.n646 B.n645 585
R338 B.n11 B.n10 585
R339 B.n644 B.n11 585
R340 B.n642 B.n641 585
R341 B.n643 B.n642 585
R342 B.n640 B.n17 585
R343 B.n17 B.n16 585
R344 B.n639 B.n638 585
R345 B.n638 B.n637 585
R346 B.n19 B.n18 585
R347 B.n636 B.n19 585
R348 B.n634 B.n633 585
R349 B.n635 B.n634 585
R350 B.n632 B.n24 585
R351 B.n24 B.n23 585
R352 B.n631 B.n630 585
R353 B.n630 B.n629 585
R354 B.n26 B.n25 585
R355 B.n628 B.n26 585
R356 B.n626 B.n625 585
R357 B.n627 B.n626 585
R358 B.n624 B.n31 585
R359 B.n31 B.n30 585
R360 B.n623 B.n622 585
R361 B.n622 B.n621 585
R362 B.n33 B.n32 585
R363 B.n620 B.n33 585
R364 B.n618 B.n617 585
R365 B.n619 B.n618 585
R366 B.n616 B.n37 585
R367 B.n40 B.n37 585
R368 B.n615 B.n614 585
R369 B.n614 B.n613 585
R370 B.n39 B.n38 585
R371 B.n612 B.n39 585
R372 B.n610 B.n609 585
R373 B.n611 B.n610 585
R374 B.n608 B.n45 585
R375 B.n45 B.n44 585
R376 B.n607 B.n606 585
R377 B.n606 B.n605 585
R378 B.n47 B.n46 585
R379 B.n604 B.n47 585
R380 B.n602 B.n601 585
R381 B.n603 B.n602 585
R382 B.n600 B.n52 585
R383 B.n52 B.n51 585
R384 B.n599 B.n598 585
R385 B.n598 B.n597 585
R386 B.n54 B.n53 585
R387 B.n596 B.n54 585
R388 B.n594 B.n593 585
R389 B.n595 B.n594 585
R390 B.n592 B.n59 585
R391 B.n59 B.n58 585
R392 B.n591 B.n590 585
R393 B.n590 B.n589 585
R394 B.n61 B.n60 585
R395 B.n588 B.n61 585
R396 B.n586 B.n585 585
R397 B.n587 B.n586 585
R398 B.n584 B.n66 585
R399 B.n66 B.n65 585
R400 B.n655 B.n654 585
R401 B.n653 B.n2 585
R402 B.n582 B.n66 497.305
R403 B.n579 B.n97 497.305
R404 B.n313 B.n275 497.305
R405 B.n425 B.n277 497.305
R406 B.n100 B.t17 278.012
R407 B.n98 B.t13 278.012
R408 B.n310 B.t10 278.012
R409 B.n308 B.t6 278.012
R410 B.n580 B.n95 256.663
R411 B.n580 B.n94 256.663
R412 B.n580 B.n93 256.663
R413 B.n580 B.n92 256.663
R414 B.n580 B.n91 256.663
R415 B.n580 B.n90 256.663
R416 B.n580 B.n89 256.663
R417 B.n580 B.n88 256.663
R418 B.n580 B.n87 256.663
R419 B.n580 B.n86 256.663
R420 B.n580 B.n85 256.663
R421 B.n580 B.n84 256.663
R422 B.n580 B.n83 256.663
R423 B.n580 B.n82 256.663
R424 B.n580 B.n81 256.663
R425 B.n580 B.n80 256.663
R426 B.n580 B.n79 256.663
R427 B.n580 B.n78 256.663
R428 B.n580 B.n77 256.663
R429 B.n580 B.n76 256.663
R430 B.n580 B.n75 256.663
R431 B.n580 B.n74 256.663
R432 B.n580 B.n73 256.663
R433 B.n580 B.n72 256.663
R434 B.n580 B.n71 256.663
R435 B.n580 B.n70 256.663
R436 B.n580 B.n69 256.663
R437 B.n581 B.n580 256.663
R438 B.n424 B.n423 256.663
R439 B.n423 B.n280 256.663
R440 B.n423 B.n281 256.663
R441 B.n423 B.n282 256.663
R442 B.n423 B.n283 256.663
R443 B.n423 B.n284 256.663
R444 B.n423 B.n285 256.663
R445 B.n423 B.n286 256.663
R446 B.n423 B.n287 256.663
R447 B.n423 B.n288 256.663
R448 B.n423 B.n289 256.663
R449 B.n423 B.n290 256.663
R450 B.n423 B.n291 256.663
R451 B.n423 B.n292 256.663
R452 B.n423 B.n293 256.663
R453 B.n423 B.n294 256.663
R454 B.n423 B.n295 256.663
R455 B.n423 B.n296 256.663
R456 B.n423 B.n297 256.663
R457 B.n423 B.n298 256.663
R458 B.n423 B.n299 256.663
R459 B.n423 B.n300 256.663
R460 B.n423 B.n301 256.663
R461 B.n423 B.n302 256.663
R462 B.n423 B.n303 256.663
R463 B.n423 B.n304 256.663
R464 B.n423 B.n305 256.663
R465 B.n423 B.n306 256.663
R466 B.n657 B.n656 256.663
R467 B.n98 B.t15 222.236
R468 B.n310 B.t12 222.236
R469 B.n100 B.t18 222.236
R470 B.n308 B.t9 222.236
R471 B.n99 B.t16 177.048
R472 B.n311 B.t11 177.048
R473 B.n101 B.t19 177.048
R474 B.n309 B.t8 177.048
R475 B.n103 B.n68 163.367
R476 B.n107 B.n106 163.367
R477 B.n111 B.n110 163.367
R478 B.n115 B.n114 163.367
R479 B.n119 B.n118 163.367
R480 B.n123 B.n122 163.367
R481 B.n127 B.n126 163.367
R482 B.n131 B.n130 163.367
R483 B.n135 B.n134 163.367
R484 B.n139 B.n138 163.367
R485 B.n143 B.n142 163.367
R486 B.n147 B.n146 163.367
R487 B.n151 B.n150 163.367
R488 B.n155 B.n154 163.367
R489 B.n159 B.n158 163.367
R490 B.n163 B.n162 163.367
R491 B.n168 B.n167 163.367
R492 B.n172 B.n171 163.367
R493 B.n176 B.n175 163.367
R494 B.n180 B.n179 163.367
R495 B.n184 B.n183 163.367
R496 B.n188 B.n187 163.367
R497 B.n192 B.n191 163.367
R498 B.n196 B.n195 163.367
R499 B.n200 B.n199 163.367
R500 B.n204 B.n203 163.367
R501 B.n208 B.n207 163.367
R502 B.n579 B.n96 163.367
R503 B.n431 B.n275 163.367
R504 B.n431 B.n273 163.367
R505 B.n435 B.n273 163.367
R506 B.n435 B.n266 163.367
R507 B.n443 B.n266 163.367
R508 B.n443 B.n264 163.367
R509 B.n447 B.n264 163.367
R510 B.n447 B.n259 163.367
R511 B.n455 B.n259 163.367
R512 B.n455 B.n257 163.367
R513 B.n459 B.n257 163.367
R514 B.n459 B.n251 163.367
R515 B.n467 B.n251 163.367
R516 B.n467 B.n249 163.367
R517 B.n471 B.n249 163.367
R518 B.n471 B.n244 163.367
R519 B.n480 B.n244 163.367
R520 B.n480 B.n242 163.367
R521 B.n484 B.n242 163.367
R522 B.n484 B.n236 163.367
R523 B.n492 B.n236 163.367
R524 B.n492 B.n234 163.367
R525 B.n496 B.n234 163.367
R526 B.n496 B.n228 163.367
R527 B.n504 B.n228 163.367
R528 B.n504 B.n226 163.367
R529 B.n508 B.n226 163.367
R530 B.n508 B.n219 163.367
R531 B.n516 B.n219 163.367
R532 B.n516 B.n217 163.367
R533 B.n521 B.n217 163.367
R534 B.n521 B.n212 163.367
R535 B.n529 B.n212 163.367
R536 B.n530 B.n529 163.367
R537 B.n530 B.n5 163.367
R538 B.n6 B.n5 163.367
R539 B.n7 B.n6 163.367
R540 B.n536 B.n7 163.367
R541 B.n537 B.n536 163.367
R542 B.n537 B.n13 163.367
R543 B.n14 B.n13 163.367
R544 B.n15 B.n14 163.367
R545 B.n542 B.n15 163.367
R546 B.n542 B.n20 163.367
R547 B.n21 B.n20 163.367
R548 B.n22 B.n21 163.367
R549 B.n547 B.n22 163.367
R550 B.n547 B.n27 163.367
R551 B.n28 B.n27 163.367
R552 B.n29 B.n28 163.367
R553 B.n552 B.n29 163.367
R554 B.n552 B.n34 163.367
R555 B.n35 B.n34 163.367
R556 B.n36 B.n35 163.367
R557 B.n557 B.n36 163.367
R558 B.n557 B.n41 163.367
R559 B.n42 B.n41 163.367
R560 B.n43 B.n42 163.367
R561 B.n562 B.n43 163.367
R562 B.n562 B.n48 163.367
R563 B.n49 B.n48 163.367
R564 B.n50 B.n49 163.367
R565 B.n567 B.n50 163.367
R566 B.n567 B.n55 163.367
R567 B.n56 B.n55 163.367
R568 B.n57 B.n56 163.367
R569 B.n572 B.n57 163.367
R570 B.n572 B.n62 163.367
R571 B.n63 B.n62 163.367
R572 B.n64 B.n63 163.367
R573 B.n97 B.n64 163.367
R574 B.n422 B.n279 163.367
R575 B.n422 B.n307 163.367
R576 B.n418 B.n417 163.367
R577 B.n414 B.n413 163.367
R578 B.n410 B.n409 163.367
R579 B.n406 B.n405 163.367
R580 B.n402 B.n401 163.367
R581 B.n398 B.n397 163.367
R582 B.n394 B.n393 163.367
R583 B.n390 B.n389 163.367
R584 B.n386 B.n385 163.367
R585 B.n382 B.n381 163.367
R586 B.n377 B.n376 163.367
R587 B.n373 B.n372 163.367
R588 B.n369 B.n368 163.367
R589 B.n365 B.n364 163.367
R590 B.n361 B.n360 163.367
R591 B.n357 B.n356 163.367
R592 B.n353 B.n352 163.367
R593 B.n349 B.n348 163.367
R594 B.n345 B.n344 163.367
R595 B.n341 B.n340 163.367
R596 B.n337 B.n336 163.367
R597 B.n333 B.n332 163.367
R598 B.n329 B.n328 163.367
R599 B.n325 B.n324 163.367
R600 B.n321 B.n320 163.367
R601 B.n317 B.n316 163.367
R602 B.n429 B.n277 163.367
R603 B.n429 B.n271 163.367
R604 B.n437 B.n271 163.367
R605 B.n437 B.n269 163.367
R606 B.n441 B.n269 163.367
R607 B.n441 B.n263 163.367
R608 B.n449 B.n263 163.367
R609 B.n449 B.n261 163.367
R610 B.n453 B.n261 163.367
R611 B.n453 B.n255 163.367
R612 B.n461 B.n255 163.367
R613 B.n461 B.n253 163.367
R614 B.n465 B.n253 163.367
R615 B.n465 B.n247 163.367
R616 B.n474 B.n247 163.367
R617 B.n474 B.n245 163.367
R618 B.n478 B.n245 163.367
R619 B.n478 B.n240 163.367
R620 B.n486 B.n240 163.367
R621 B.n486 B.n238 163.367
R622 B.n490 B.n238 163.367
R623 B.n490 B.n232 163.367
R624 B.n498 B.n232 163.367
R625 B.n498 B.n230 163.367
R626 B.n502 B.n230 163.367
R627 B.n502 B.n224 163.367
R628 B.n510 B.n224 163.367
R629 B.n510 B.n222 163.367
R630 B.n514 B.n222 163.367
R631 B.n514 B.n216 163.367
R632 B.n523 B.n216 163.367
R633 B.n523 B.n214 163.367
R634 B.n527 B.n214 163.367
R635 B.n527 B.n3 163.367
R636 B.n655 B.n3 163.367
R637 B.n651 B.n2 163.367
R638 B.n651 B.n650 163.367
R639 B.n650 B.n9 163.367
R640 B.n646 B.n9 163.367
R641 B.n646 B.n11 163.367
R642 B.n642 B.n11 163.367
R643 B.n642 B.n17 163.367
R644 B.n638 B.n17 163.367
R645 B.n638 B.n19 163.367
R646 B.n634 B.n19 163.367
R647 B.n634 B.n24 163.367
R648 B.n630 B.n24 163.367
R649 B.n630 B.n26 163.367
R650 B.n626 B.n26 163.367
R651 B.n626 B.n31 163.367
R652 B.n622 B.n31 163.367
R653 B.n622 B.n33 163.367
R654 B.n618 B.n33 163.367
R655 B.n618 B.n37 163.367
R656 B.n614 B.n37 163.367
R657 B.n614 B.n39 163.367
R658 B.n610 B.n39 163.367
R659 B.n610 B.n45 163.367
R660 B.n606 B.n45 163.367
R661 B.n606 B.n47 163.367
R662 B.n602 B.n47 163.367
R663 B.n602 B.n52 163.367
R664 B.n598 B.n52 163.367
R665 B.n598 B.n54 163.367
R666 B.n594 B.n54 163.367
R667 B.n594 B.n59 163.367
R668 B.n590 B.n59 163.367
R669 B.n590 B.n61 163.367
R670 B.n586 B.n61 163.367
R671 B.n586 B.n66 163.367
R672 B.n423 B.n276 123.043
R673 B.n580 B.n65 123.043
R674 B.n582 B.n581 71.676
R675 B.n103 B.n69 71.676
R676 B.n107 B.n70 71.676
R677 B.n111 B.n71 71.676
R678 B.n115 B.n72 71.676
R679 B.n119 B.n73 71.676
R680 B.n123 B.n74 71.676
R681 B.n127 B.n75 71.676
R682 B.n131 B.n76 71.676
R683 B.n135 B.n77 71.676
R684 B.n139 B.n78 71.676
R685 B.n143 B.n79 71.676
R686 B.n147 B.n80 71.676
R687 B.n151 B.n81 71.676
R688 B.n155 B.n82 71.676
R689 B.n159 B.n83 71.676
R690 B.n163 B.n84 71.676
R691 B.n168 B.n85 71.676
R692 B.n172 B.n86 71.676
R693 B.n176 B.n87 71.676
R694 B.n180 B.n88 71.676
R695 B.n184 B.n89 71.676
R696 B.n188 B.n90 71.676
R697 B.n192 B.n91 71.676
R698 B.n196 B.n92 71.676
R699 B.n200 B.n93 71.676
R700 B.n204 B.n94 71.676
R701 B.n208 B.n95 71.676
R702 B.n96 B.n95 71.676
R703 B.n207 B.n94 71.676
R704 B.n203 B.n93 71.676
R705 B.n199 B.n92 71.676
R706 B.n195 B.n91 71.676
R707 B.n191 B.n90 71.676
R708 B.n187 B.n89 71.676
R709 B.n183 B.n88 71.676
R710 B.n179 B.n87 71.676
R711 B.n175 B.n86 71.676
R712 B.n171 B.n85 71.676
R713 B.n167 B.n84 71.676
R714 B.n162 B.n83 71.676
R715 B.n158 B.n82 71.676
R716 B.n154 B.n81 71.676
R717 B.n150 B.n80 71.676
R718 B.n146 B.n79 71.676
R719 B.n142 B.n78 71.676
R720 B.n138 B.n77 71.676
R721 B.n134 B.n76 71.676
R722 B.n130 B.n75 71.676
R723 B.n126 B.n74 71.676
R724 B.n122 B.n73 71.676
R725 B.n118 B.n72 71.676
R726 B.n114 B.n71 71.676
R727 B.n110 B.n70 71.676
R728 B.n106 B.n69 71.676
R729 B.n581 B.n68 71.676
R730 B.n425 B.n424 71.676
R731 B.n307 B.n280 71.676
R732 B.n417 B.n281 71.676
R733 B.n413 B.n282 71.676
R734 B.n409 B.n283 71.676
R735 B.n405 B.n284 71.676
R736 B.n401 B.n285 71.676
R737 B.n397 B.n286 71.676
R738 B.n393 B.n287 71.676
R739 B.n389 B.n288 71.676
R740 B.n385 B.n289 71.676
R741 B.n381 B.n290 71.676
R742 B.n376 B.n291 71.676
R743 B.n372 B.n292 71.676
R744 B.n368 B.n293 71.676
R745 B.n364 B.n294 71.676
R746 B.n360 B.n295 71.676
R747 B.n356 B.n296 71.676
R748 B.n352 B.n297 71.676
R749 B.n348 B.n298 71.676
R750 B.n344 B.n299 71.676
R751 B.n340 B.n300 71.676
R752 B.n336 B.n301 71.676
R753 B.n332 B.n302 71.676
R754 B.n328 B.n303 71.676
R755 B.n324 B.n304 71.676
R756 B.n320 B.n305 71.676
R757 B.n316 B.n306 71.676
R758 B.n424 B.n279 71.676
R759 B.n418 B.n280 71.676
R760 B.n414 B.n281 71.676
R761 B.n410 B.n282 71.676
R762 B.n406 B.n283 71.676
R763 B.n402 B.n284 71.676
R764 B.n398 B.n285 71.676
R765 B.n394 B.n286 71.676
R766 B.n390 B.n287 71.676
R767 B.n386 B.n288 71.676
R768 B.n382 B.n289 71.676
R769 B.n377 B.n290 71.676
R770 B.n373 B.n291 71.676
R771 B.n369 B.n292 71.676
R772 B.n365 B.n293 71.676
R773 B.n361 B.n294 71.676
R774 B.n357 B.n295 71.676
R775 B.n353 B.n296 71.676
R776 B.n349 B.n297 71.676
R777 B.n345 B.n298 71.676
R778 B.n341 B.n299 71.676
R779 B.n337 B.n300 71.676
R780 B.n333 B.n301 71.676
R781 B.n329 B.n302 71.676
R782 B.n325 B.n303 71.676
R783 B.n321 B.n304 71.676
R784 B.n317 B.n305 71.676
R785 B.n313 B.n306 71.676
R786 B.n656 B.n655 71.676
R787 B.n656 B.n2 71.676
R788 B.n430 B.n276 66.9356
R789 B.n430 B.n272 66.9356
R790 B.n436 B.n272 66.9356
R791 B.n436 B.n267 66.9356
R792 B.n442 B.n267 66.9356
R793 B.n442 B.n268 66.9356
R794 B.n448 B.n260 66.9356
R795 B.n454 B.n260 66.9356
R796 B.n454 B.n256 66.9356
R797 B.n460 B.n256 66.9356
R798 B.n460 B.n252 66.9356
R799 B.n466 B.n252 66.9356
R800 B.n466 B.n248 66.9356
R801 B.n473 B.n248 66.9356
R802 B.n473 B.n472 66.9356
R803 B.n479 B.n241 66.9356
R804 B.n485 B.n241 66.9356
R805 B.n485 B.n237 66.9356
R806 B.n491 B.n237 66.9356
R807 B.n491 B.n233 66.9356
R808 B.n497 B.n233 66.9356
R809 B.n503 B.n229 66.9356
R810 B.n503 B.n225 66.9356
R811 B.n509 B.n225 66.9356
R812 B.n509 B.n220 66.9356
R813 B.n515 B.n220 66.9356
R814 B.n515 B.n221 66.9356
R815 B.n522 B.n213 66.9356
R816 B.n528 B.n213 66.9356
R817 B.n528 B.n4 66.9356
R818 B.n654 B.n4 66.9356
R819 B.n654 B.n653 66.9356
R820 B.n653 B.n652 66.9356
R821 B.n652 B.n8 66.9356
R822 B.n12 B.n8 66.9356
R823 B.n645 B.n12 66.9356
R824 B.n644 B.n643 66.9356
R825 B.n643 B.n16 66.9356
R826 B.n637 B.n16 66.9356
R827 B.n637 B.n636 66.9356
R828 B.n636 B.n635 66.9356
R829 B.n635 B.n23 66.9356
R830 B.n629 B.n628 66.9356
R831 B.n628 B.n627 66.9356
R832 B.n627 B.n30 66.9356
R833 B.n621 B.n30 66.9356
R834 B.n621 B.n620 66.9356
R835 B.n620 B.n619 66.9356
R836 B.n613 B.n40 66.9356
R837 B.n613 B.n612 66.9356
R838 B.n612 B.n611 66.9356
R839 B.n611 B.n44 66.9356
R840 B.n605 B.n44 66.9356
R841 B.n605 B.n604 66.9356
R842 B.n604 B.n603 66.9356
R843 B.n603 B.n51 66.9356
R844 B.n597 B.n51 66.9356
R845 B.n596 B.n595 66.9356
R846 B.n595 B.n58 66.9356
R847 B.n589 B.n58 66.9356
R848 B.n589 B.n588 66.9356
R849 B.n588 B.n587 66.9356
R850 B.n587 B.n65 66.9356
R851 B.n102 B.n101 59.5399
R852 B.n165 B.n99 59.5399
R853 B.n312 B.n311 59.5399
R854 B.n379 B.n309 59.5399
R855 B.n472 B.t4 51.1862
R856 B.n40 B.t0 51.1862
R857 B.n268 B.t7 47.2488
R858 B.t14 B.n596 47.2488
R859 B.n101 B.n100 45.1884
R860 B.n99 B.n98 45.1884
R861 B.n311 B.n310 45.1884
R862 B.n309 B.n308 45.1884
R863 B.n497 B.t1 41.3428
R864 B.n629 B.t2 41.3428
R865 B.n522 B.t3 35.4367
R866 B.n645 B.t5 35.4367
R867 B.n427 B.n426 32.3127
R868 B.n314 B.n274 32.3127
R869 B.n578 B.n577 32.3127
R870 B.n584 B.n583 32.3127
R871 B.n221 B.t3 31.4994
R872 B.t5 B.n644 31.4994
R873 B.t1 B.n229 25.5933
R874 B.t2 B.n23 25.5933
R875 B.n448 B.t7 19.6873
R876 B.n597 B.t14 19.6873
R877 B B.n657 18.0485
R878 B.n479 B.t4 15.7499
R879 B.n619 B.t0 15.7499
R880 B.n428 B.n427 10.6151
R881 B.n428 B.n270 10.6151
R882 B.n438 B.n270 10.6151
R883 B.n439 B.n438 10.6151
R884 B.n440 B.n439 10.6151
R885 B.n440 B.n262 10.6151
R886 B.n450 B.n262 10.6151
R887 B.n451 B.n450 10.6151
R888 B.n452 B.n451 10.6151
R889 B.n452 B.n254 10.6151
R890 B.n462 B.n254 10.6151
R891 B.n463 B.n462 10.6151
R892 B.n464 B.n463 10.6151
R893 B.n464 B.n246 10.6151
R894 B.n475 B.n246 10.6151
R895 B.n476 B.n475 10.6151
R896 B.n477 B.n476 10.6151
R897 B.n477 B.n239 10.6151
R898 B.n487 B.n239 10.6151
R899 B.n488 B.n487 10.6151
R900 B.n489 B.n488 10.6151
R901 B.n489 B.n231 10.6151
R902 B.n499 B.n231 10.6151
R903 B.n500 B.n499 10.6151
R904 B.n501 B.n500 10.6151
R905 B.n501 B.n223 10.6151
R906 B.n511 B.n223 10.6151
R907 B.n512 B.n511 10.6151
R908 B.n513 B.n512 10.6151
R909 B.n513 B.n215 10.6151
R910 B.n524 B.n215 10.6151
R911 B.n525 B.n524 10.6151
R912 B.n526 B.n525 10.6151
R913 B.n526 B.n0 10.6151
R914 B.n426 B.n278 10.6151
R915 B.n421 B.n278 10.6151
R916 B.n421 B.n420 10.6151
R917 B.n420 B.n419 10.6151
R918 B.n419 B.n416 10.6151
R919 B.n416 B.n415 10.6151
R920 B.n415 B.n412 10.6151
R921 B.n412 B.n411 10.6151
R922 B.n411 B.n408 10.6151
R923 B.n408 B.n407 10.6151
R924 B.n407 B.n404 10.6151
R925 B.n404 B.n403 10.6151
R926 B.n403 B.n400 10.6151
R927 B.n400 B.n399 10.6151
R928 B.n399 B.n396 10.6151
R929 B.n396 B.n395 10.6151
R930 B.n395 B.n392 10.6151
R931 B.n392 B.n391 10.6151
R932 B.n391 B.n388 10.6151
R933 B.n388 B.n387 10.6151
R934 B.n387 B.n384 10.6151
R935 B.n384 B.n383 10.6151
R936 B.n383 B.n380 10.6151
R937 B.n378 B.n375 10.6151
R938 B.n375 B.n374 10.6151
R939 B.n374 B.n371 10.6151
R940 B.n371 B.n370 10.6151
R941 B.n370 B.n367 10.6151
R942 B.n367 B.n366 10.6151
R943 B.n366 B.n363 10.6151
R944 B.n363 B.n362 10.6151
R945 B.n359 B.n358 10.6151
R946 B.n358 B.n355 10.6151
R947 B.n355 B.n354 10.6151
R948 B.n354 B.n351 10.6151
R949 B.n351 B.n350 10.6151
R950 B.n350 B.n347 10.6151
R951 B.n347 B.n346 10.6151
R952 B.n346 B.n343 10.6151
R953 B.n343 B.n342 10.6151
R954 B.n342 B.n339 10.6151
R955 B.n339 B.n338 10.6151
R956 B.n338 B.n335 10.6151
R957 B.n335 B.n334 10.6151
R958 B.n334 B.n331 10.6151
R959 B.n331 B.n330 10.6151
R960 B.n330 B.n327 10.6151
R961 B.n327 B.n326 10.6151
R962 B.n326 B.n323 10.6151
R963 B.n323 B.n322 10.6151
R964 B.n322 B.n319 10.6151
R965 B.n319 B.n318 10.6151
R966 B.n318 B.n315 10.6151
R967 B.n315 B.n314 10.6151
R968 B.n432 B.n274 10.6151
R969 B.n433 B.n432 10.6151
R970 B.n434 B.n433 10.6151
R971 B.n434 B.n265 10.6151
R972 B.n444 B.n265 10.6151
R973 B.n445 B.n444 10.6151
R974 B.n446 B.n445 10.6151
R975 B.n446 B.n258 10.6151
R976 B.n456 B.n258 10.6151
R977 B.n457 B.n456 10.6151
R978 B.n458 B.n457 10.6151
R979 B.n458 B.n250 10.6151
R980 B.n468 B.n250 10.6151
R981 B.n469 B.n468 10.6151
R982 B.n470 B.n469 10.6151
R983 B.n470 B.n243 10.6151
R984 B.n481 B.n243 10.6151
R985 B.n482 B.n481 10.6151
R986 B.n483 B.n482 10.6151
R987 B.n483 B.n235 10.6151
R988 B.n493 B.n235 10.6151
R989 B.n494 B.n493 10.6151
R990 B.n495 B.n494 10.6151
R991 B.n495 B.n227 10.6151
R992 B.n505 B.n227 10.6151
R993 B.n506 B.n505 10.6151
R994 B.n507 B.n506 10.6151
R995 B.n507 B.n218 10.6151
R996 B.n517 B.n218 10.6151
R997 B.n518 B.n517 10.6151
R998 B.n520 B.n518 10.6151
R999 B.n520 B.n519 10.6151
R1000 B.n519 B.n211 10.6151
R1001 B.n531 B.n211 10.6151
R1002 B.n532 B.n531 10.6151
R1003 B.n533 B.n532 10.6151
R1004 B.n534 B.n533 10.6151
R1005 B.n535 B.n534 10.6151
R1006 B.n538 B.n535 10.6151
R1007 B.n539 B.n538 10.6151
R1008 B.n540 B.n539 10.6151
R1009 B.n541 B.n540 10.6151
R1010 B.n543 B.n541 10.6151
R1011 B.n544 B.n543 10.6151
R1012 B.n545 B.n544 10.6151
R1013 B.n546 B.n545 10.6151
R1014 B.n548 B.n546 10.6151
R1015 B.n549 B.n548 10.6151
R1016 B.n550 B.n549 10.6151
R1017 B.n551 B.n550 10.6151
R1018 B.n553 B.n551 10.6151
R1019 B.n554 B.n553 10.6151
R1020 B.n555 B.n554 10.6151
R1021 B.n556 B.n555 10.6151
R1022 B.n558 B.n556 10.6151
R1023 B.n559 B.n558 10.6151
R1024 B.n560 B.n559 10.6151
R1025 B.n561 B.n560 10.6151
R1026 B.n563 B.n561 10.6151
R1027 B.n564 B.n563 10.6151
R1028 B.n565 B.n564 10.6151
R1029 B.n566 B.n565 10.6151
R1030 B.n568 B.n566 10.6151
R1031 B.n569 B.n568 10.6151
R1032 B.n570 B.n569 10.6151
R1033 B.n571 B.n570 10.6151
R1034 B.n573 B.n571 10.6151
R1035 B.n574 B.n573 10.6151
R1036 B.n575 B.n574 10.6151
R1037 B.n576 B.n575 10.6151
R1038 B.n577 B.n576 10.6151
R1039 B.n649 B.n1 10.6151
R1040 B.n649 B.n648 10.6151
R1041 B.n648 B.n647 10.6151
R1042 B.n647 B.n10 10.6151
R1043 B.n641 B.n10 10.6151
R1044 B.n641 B.n640 10.6151
R1045 B.n640 B.n639 10.6151
R1046 B.n639 B.n18 10.6151
R1047 B.n633 B.n18 10.6151
R1048 B.n633 B.n632 10.6151
R1049 B.n632 B.n631 10.6151
R1050 B.n631 B.n25 10.6151
R1051 B.n625 B.n25 10.6151
R1052 B.n625 B.n624 10.6151
R1053 B.n624 B.n623 10.6151
R1054 B.n623 B.n32 10.6151
R1055 B.n617 B.n32 10.6151
R1056 B.n617 B.n616 10.6151
R1057 B.n616 B.n615 10.6151
R1058 B.n615 B.n38 10.6151
R1059 B.n609 B.n38 10.6151
R1060 B.n609 B.n608 10.6151
R1061 B.n608 B.n607 10.6151
R1062 B.n607 B.n46 10.6151
R1063 B.n601 B.n46 10.6151
R1064 B.n601 B.n600 10.6151
R1065 B.n600 B.n599 10.6151
R1066 B.n599 B.n53 10.6151
R1067 B.n593 B.n53 10.6151
R1068 B.n593 B.n592 10.6151
R1069 B.n592 B.n591 10.6151
R1070 B.n591 B.n60 10.6151
R1071 B.n585 B.n60 10.6151
R1072 B.n585 B.n584 10.6151
R1073 B.n583 B.n67 10.6151
R1074 B.n104 B.n67 10.6151
R1075 B.n105 B.n104 10.6151
R1076 B.n108 B.n105 10.6151
R1077 B.n109 B.n108 10.6151
R1078 B.n112 B.n109 10.6151
R1079 B.n113 B.n112 10.6151
R1080 B.n116 B.n113 10.6151
R1081 B.n117 B.n116 10.6151
R1082 B.n120 B.n117 10.6151
R1083 B.n121 B.n120 10.6151
R1084 B.n124 B.n121 10.6151
R1085 B.n125 B.n124 10.6151
R1086 B.n128 B.n125 10.6151
R1087 B.n129 B.n128 10.6151
R1088 B.n132 B.n129 10.6151
R1089 B.n133 B.n132 10.6151
R1090 B.n136 B.n133 10.6151
R1091 B.n137 B.n136 10.6151
R1092 B.n140 B.n137 10.6151
R1093 B.n141 B.n140 10.6151
R1094 B.n144 B.n141 10.6151
R1095 B.n145 B.n144 10.6151
R1096 B.n149 B.n148 10.6151
R1097 B.n152 B.n149 10.6151
R1098 B.n153 B.n152 10.6151
R1099 B.n156 B.n153 10.6151
R1100 B.n157 B.n156 10.6151
R1101 B.n160 B.n157 10.6151
R1102 B.n161 B.n160 10.6151
R1103 B.n164 B.n161 10.6151
R1104 B.n169 B.n166 10.6151
R1105 B.n170 B.n169 10.6151
R1106 B.n173 B.n170 10.6151
R1107 B.n174 B.n173 10.6151
R1108 B.n177 B.n174 10.6151
R1109 B.n178 B.n177 10.6151
R1110 B.n181 B.n178 10.6151
R1111 B.n182 B.n181 10.6151
R1112 B.n185 B.n182 10.6151
R1113 B.n186 B.n185 10.6151
R1114 B.n189 B.n186 10.6151
R1115 B.n190 B.n189 10.6151
R1116 B.n193 B.n190 10.6151
R1117 B.n194 B.n193 10.6151
R1118 B.n197 B.n194 10.6151
R1119 B.n198 B.n197 10.6151
R1120 B.n201 B.n198 10.6151
R1121 B.n202 B.n201 10.6151
R1122 B.n205 B.n202 10.6151
R1123 B.n206 B.n205 10.6151
R1124 B.n209 B.n206 10.6151
R1125 B.n210 B.n209 10.6151
R1126 B.n578 B.n210 10.6151
R1127 B.n657 B.n0 8.11757
R1128 B.n657 B.n1 8.11757
R1129 B.n379 B.n378 6.5566
R1130 B.n362 B.n312 6.5566
R1131 B.n148 B.n102 6.5566
R1132 B.n165 B.n164 6.5566
R1133 B.n380 B.n379 4.05904
R1134 B.n359 B.n312 4.05904
R1135 B.n145 B.n102 4.05904
R1136 B.n166 B.n165 4.05904
R1137 VN.n21 VN.n12 161.3
R1138 VN.n20 VN.n19 161.3
R1139 VN.n18 VN.n13 161.3
R1140 VN.n17 VN.n16 161.3
R1141 VN.n9 VN.n0 161.3
R1142 VN.n8 VN.n7 161.3
R1143 VN.n6 VN.n1 161.3
R1144 VN.n5 VN.n4 161.3
R1145 VN.n2 VN.t0 104.612
R1146 VN.n14 VN.t3 104.612
R1147 VN.n11 VN.n10 94.6776
R1148 VN.n23 VN.n22 94.6776
R1149 VN.n3 VN.t4 71.0955
R1150 VN.n10 VN.t5 71.0955
R1151 VN.n15 VN.t1 71.0955
R1152 VN.n22 VN.t2 71.0955
R1153 VN.n8 VN.n1 56.5617
R1154 VN.n20 VN.n13 56.5617
R1155 VN.n15 VN.n14 45.8151
R1156 VN.n3 VN.n2 45.8151
R1157 VN VN.n23 41.9489
R1158 VN.n4 VN.n3 24.5923
R1159 VN.n4 VN.n1 24.5923
R1160 VN.n9 VN.n8 24.5923
R1161 VN.n16 VN.n13 24.5923
R1162 VN.n16 VN.n15 24.5923
R1163 VN.n21 VN.n20 24.5923
R1164 VN.n10 VN.n9 16.2311
R1165 VN.n22 VN.n21 16.2311
R1166 VN.n5 VN.n2 9.3086
R1167 VN.n17 VN.n14 9.3086
R1168 VN.n23 VN.n12 0.278335
R1169 VN.n11 VN.n0 0.278335
R1170 VN.n19 VN.n12 0.189894
R1171 VN.n19 VN.n18 0.189894
R1172 VN.n18 VN.n17 0.189894
R1173 VN.n6 VN.n5 0.189894
R1174 VN.n7 VN.n6 0.189894
R1175 VN.n7 VN.n0 0.189894
R1176 VN VN.n11 0.153485
R1177 VTAIL.n130 VTAIL.n104 289.615
R1178 VTAIL.n28 VTAIL.n2 289.615
R1179 VTAIL.n98 VTAIL.n72 289.615
R1180 VTAIL.n64 VTAIL.n38 289.615
R1181 VTAIL.n115 VTAIL.n114 185
R1182 VTAIL.n112 VTAIL.n111 185
R1183 VTAIL.n121 VTAIL.n120 185
R1184 VTAIL.n123 VTAIL.n122 185
R1185 VTAIL.n108 VTAIL.n107 185
R1186 VTAIL.n129 VTAIL.n128 185
R1187 VTAIL.n131 VTAIL.n130 185
R1188 VTAIL.n13 VTAIL.n12 185
R1189 VTAIL.n10 VTAIL.n9 185
R1190 VTAIL.n19 VTAIL.n18 185
R1191 VTAIL.n21 VTAIL.n20 185
R1192 VTAIL.n6 VTAIL.n5 185
R1193 VTAIL.n27 VTAIL.n26 185
R1194 VTAIL.n29 VTAIL.n28 185
R1195 VTAIL.n99 VTAIL.n98 185
R1196 VTAIL.n97 VTAIL.n96 185
R1197 VTAIL.n76 VTAIL.n75 185
R1198 VTAIL.n91 VTAIL.n90 185
R1199 VTAIL.n89 VTAIL.n88 185
R1200 VTAIL.n80 VTAIL.n79 185
R1201 VTAIL.n83 VTAIL.n82 185
R1202 VTAIL.n65 VTAIL.n64 185
R1203 VTAIL.n63 VTAIL.n62 185
R1204 VTAIL.n42 VTAIL.n41 185
R1205 VTAIL.n57 VTAIL.n56 185
R1206 VTAIL.n55 VTAIL.n54 185
R1207 VTAIL.n46 VTAIL.n45 185
R1208 VTAIL.n49 VTAIL.n48 185
R1209 VTAIL.t10 VTAIL.n113 147.661
R1210 VTAIL.t1 VTAIL.n11 147.661
R1211 VTAIL.t2 VTAIL.n81 147.661
R1212 VTAIL.t11 VTAIL.n47 147.661
R1213 VTAIL.n114 VTAIL.n111 104.615
R1214 VTAIL.n121 VTAIL.n111 104.615
R1215 VTAIL.n122 VTAIL.n121 104.615
R1216 VTAIL.n122 VTAIL.n107 104.615
R1217 VTAIL.n129 VTAIL.n107 104.615
R1218 VTAIL.n130 VTAIL.n129 104.615
R1219 VTAIL.n12 VTAIL.n9 104.615
R1220 VTAIL.n19 VTAIL.n9 104.615
R1221 VTAIL.n20 VTAIL.n19 104.615
R1222 VTAIL.n20 VTAIL.n5 104.615
R1223 VTAIL.n27 VTAIL.n5 104.615
R1224 VTAIL.n28 VTAIL.n27 104.615
R1225 VTAIL.n98 VTAIL.n97 104.615
R1226 VTAIL.n97 VTAIL.n75 104.615
R1227 VTAIL.n90 VTAIL.n75 104.615
R1228 VTAIL.n90 VTAIL.n89 104.615
R1229 VTAIL.n89 VTAIL.n79 104.615
R1230 VTAIL.n82 VTAIL.n79 104.615
R1231 VTAIL.n64 VTAIL.n63 104.615
R1232 VTAIL.n63 VTAIL.n41 104.615
R1233 VTAIL.n56 VTAIL.n41 104.615
R1234 VTAIL.n56 VTAIL.n55 104.615
R1235 VTAIL.n55 VTAIL.n45 104.615
R1236 VTAIL.n48 VTAIL.n45 104.615
R1237 VTAIL.n114 VTAIL.t10 52.3082
R1238 VTAIL.n12 VTAIL.t1 52.3082
R1239 VTAIL.n82 VTAIL.t2 52.3082
R1240 VTAIL.n48 VTAIL.t11 52.3082
R1241 VTAIL.n71 VTAIL.n70 48.5726
R1242 VTAIL.n37 VTAIL.n36 48.5726
R1243 VTAIL.n1 VTAIL.n0 48.5725
R1244 VTAIL.n35 VTAIL.n34 48.5725
R1245 VTAIL.n135 VTAIL.n134 30.246
R1246 VTAIL.n33 VTAIL.n32 30.246
R1247 VTAIL.n103 VTAIL.n102 30.246
R1248 VTAIL.n69 VTAIL.n68 30.246
R1249 VTAIL.n37 VTAIL.n35 21.4703
R1250 VTAIL.n135 VTAIL.n103 19.4617
R1251 VTAIL.n115 VTAIL.n113 15.6674
R1252 VTAIL.n13 VTAIL.n11 15.6674
R1253 VTAIL.n83 VTAIL.n81 15.6674
R1254 VTAIL.n49 VTAIL.n47 15.6674
R1255 VTAIL.n116 VTAIL.n112 12.8005
R1256 VTAIL.n14 VTAIL.n10 12.8005
R1257 VTAIL.n84 VTAIL.n80 12.8005
R1258 VTAIL.n50 VTAIL.n46 12.8005
R1259 VTAIL.n120 VTAIL.n119 12.0247
R1260 VTAIL.n18 VTAIL.n17 12.0247
R1261 VTAIL.n88 VTAIL.n87 12.0247
R1262 VTAIL.n54 VTAIL.n53 12.0247
R1263 VTAIL.n123 VTAIL.n110 11.249
R1264 VTAIL.n21 VTAIL.n8 11.249
R1265 VTAIL.n91 VTAIL.n78 11.249
R1266 VTAIL.n57 VTAIL.n44 11.249
R1267 VTAIL.n124 VTAIL.n108 10.4732
R1268 VTAIL.n22 VTAIL.n6 10.4732
R1269 VTAIL.n92 VTAIL.n76 10.4732
R1270 VTAIL.n58 VTAIL.n42 10.4732
R1271 VTAIL.n128 VTAIL.n127 9.69747
R1272 VTAIL.n26 VTAIL.n25 9.69747
R1273 VTAIL.n96 VTAIL.n95 9.69747
R1274 VTAIL.n62 VTAIL.n61 9.69747
R1275 VTAIL.n134 VTAIL.n133 9.45567
R1276 VTAIL.n32 VTAIL.n31 9.45567
R1277 VTAIL.n102 VTAIL.n101 9.45567
R1278 VTAIL.n68 VTAIL.n67 9.45567
R1279 VTAIL.n133 VTAIL.n132 9.3005
R1280 VTAIL.n106 VTAIL.n105 9.3005
R1281 VTAIL.n127 VTAIL.n126 9.3005
R1282 VTAIL.n125 VTAIL.n124 9.3005
R1283 VTAIL.n110 VTAIL.n109 9.3005
R1284 VTAIL.n119 VTAIL.n118 9.3005
R1285 VTAIL.n117 VTAIL.n116 9.3005
R1286 VTAIL.n31 VTAIL.n30 9.3005
R1287 VTAIL.n4 VTAIL.n3 9.3005
R1288 VTAIL.n25 VTAIL.n24 9.3005
R1289 VTAIL.n23 VTAIL.n22 9.3005
R1290 VTAIL.n8 VTAIL.n7 9.3005
R1291 VTAIL.n17 VTAIL.n16 9.3005
R1292 VTAIL.n15 VTAIL.n14 9.3005
R1293 VTAIL.n101 VTAIL.n100 9.3005
R1294 VTAIL.n74 VTAIL.n73 9.3005
R1295 VTAIL.n95 VTAIL.n94 9.3005
R1296 VTAIL.n93 VTAIL.n92 9.3005
R1297 VTAIL.n78 VTAIL.n77 9.3005
R1298 VTAIL.n87 VTAIL.n86 9.3005
R1299 VTAIL.n85 VTAIL.n84 9.3005
R1300 VTAIL.n67 VTAIL.n66 9.3005
R1301 VTAIL.n40 VTAIL.n39 9.3005
R1302 VTAIL.n61 VTAIL.n60 9.3005
R1303 VTAIL.n59 VTAIL.n58 9.3005
R1304 VTAIL.n44 VTAIL.n43 9.3005
R1305 VTAIL.n53 VTAIL.n52 9.3005
R1306 VTAIL.n51 VTAIL.n50 9.3005
R1307 VTAIL.n131 VTAIL.n106 8.92171
R1308 VTAIL.n29 VTAIL.n4 8.92171
R1309 VTAIL.n99 VTAIL.n74 8.92171
R1310 VTAIL.n65 VTAIL.n40 8.92171
R1311 VTAIL.n132 VTAIL.n104 8.14595
R1312 VTAIL.n30 VTAIL.n2 8.14595
R1313 VTAIL.n100 VTAIL.n72 8.14595
R1314 VTAIL.n66 VTAIL.n38 8.14595
R1315 VTAIL.n134 VTAIL.n104 5.81868
R1316 VTAIL.n32 VTAIL.n2 5.81868
R1317 VTAIL.n102 VTAIL.n72 5.81868
R1318 VTAIL.n68 VTAIL.n38 5.81868
R1319 VTAIL.n132 VTAIL.n131 5.04292
R1320 VTAIL.n30 VTAIL.n29 5.04292
R1321 VTAIL.n100 VTAIL.n99 5.04292
R1322 VTAIL.n66 VTAIL.n65 5.04292
R1323 VTAIL.n117 VTAIL.n113 4.38594
R1324 VTAIL.n15 VTAIL.n11 4.38594
R1325 VTAIL.n85 VTAIL.n81 4.38594
R1326 VTAIL.n51 VTAIL.n47 4.38594
R1327 VTAIL.n128 VTAIL.n106 4.26717
R1328 VTAIL.n26 VTAIL.n4 4.26717
R1329 VTAIL.n96 VTAIL.n74 4.26717
R1330 VTAIL.n62 VTAIL.n40 4.26717
R1331 VTAIL.n127 VTAIL.n108 3.49141
R1332 VTAIL.n25 VTAIL.n6 3.49141
R1333 VTAIL.n95 VTAIL.n76 3.49141
R1334 VTAIL.n61 VTAIL.n42 3.49141
R1335 VTAIL.n0 VTAIL.t6 3.35643
R1336 VTAIL.n0 VTAIL.t8 3.35643
R1337 VTAIL.n34 VTAIL.t4 3.35643
R1338 VTAIL.n34 VTAIL.t3 3.35643
R1339 VTAIL.n70 VTAIL.t5 3.35643
R1340 VTAIL.n70 VTAIL.t0 3.35643
R1341 VTAIL.n36 VTAIL.t9 3.35643
R1342 VTAIL.n36 VTAIL.t7 3.35643
R1343 VTAIL.n124 VTAIL.n123 2.71565
R1344 VTAIL.n22 VTAIL.n21 2.71565
R1345 VTAIL.n92 VTAIL.n91 2.71565
R1346 VTAIL.n58 VTAIL.n57 2.71565
R1347 VTAIL.n69 VTAIL.n37 2.00912
R1348 VTAIL.n103 VTAIL.n71 2.00912
R1349 VTAIL.n35 VTAIL.n33 2.00912
R1350 VTAIL.n120 VTAIL.n110 1.93989
R1351 VTAIL.n18 VTAIL.n8 1.93989
R1352 VTAIL.n88 VTAIL.n78 1.93989
R1353 VTAIL.n54 VTAIL.n44 1.93989
R1354 VTAIL.n71 VTAIL.n69 1.47464
R1355 VTAIL.n33 VTAIL.n1 1.47464
R1356 VTAIL VTAIL.n135 1.44878
R1357 VTAIL.n119 VTAIL.n112 1.16414
R1358 VTAIL.n17 VTAIL.n10 1.16414
R1359 VTAIL.n87 VTAIL.n80 1.16414
R1360 VTAIL.n53 VTAIL.n46 1.16414
R1361 VTAIL VTAIL.n1 0.560845
R1362 VTAIL.n116 VTAIL.n115 0.388379
R1363 VTAIL.n14 VTAIL.n13 0.388379
R1364 VTAIL.n84 VTAIL.n83 0.388379
R1365 VTAIL.n50 VTAIL.n49 0.388379
R1366 VTAIL.n118 VTAIL.n117 0.155672
R1367 VTAIL.n118 VTAIL.n109 0.155672
R1368 VTAIL.n125 VTAIL.n109 0.155672
R1369 VTAIL.n126 VTAIL.n125 0.155672
R1370 VTAIL.n126 VTAIL.n105 0.155672
R1371 VTAIL.n133 VTAIL.n105 0.155672
R1372 VTAIL.n16 VTAIL.n15 0.155672
R1373 VTAIL.n16 VTAIL.n7 0.155672
R1374 VTAIL.n23 VTAIL.n7 0.155672
R1375 VTAIL.n24 VTAIL.n23 0.155672
R1376 VTAIL.n24 VTAIL.n3 0.155672
R1377 VTAIL.n31 VTAIL.n3 0.155672
R1378 VTAIL.n101 VTAIL.n73 0.155672
R1379 VTAIL.n94 VTAIL.n73 0.155672
R1380 VTAIL.n94 VTAIL.n93 0.155672
R1381 VTAIL.n93 VTAIL.n77 0.155672
R1382 VTAIL.n86 VTAIL.n77 0.155672
R1383 VTAIL.n86 VTAIL.n85 0.155672
R1384 VTAIL.n67 VTAIL.n39 0.155672
R1385 VTAIL.n60 VTAIL.n39 0.155672
R1386 VTAIL.n60 VTAIL.n59 0.155672
R1387 VTAIL.n59 VTAIL.n43 0.155672
R1388 VTAIL.n52 VTAIL.n43 0.155672
R1389 VTAIL.n52 VTAIL.n51 0.155672
R1390 VDD2.n59 VDD2.n33 289.615
R1391 VDD2.n26 VDD2.n0 289.615
R1392 VDD2.n60 VDD2.n59 185
R1393 VDD2.n58 VDD2.n57 185
R1394 VDD2.n37 VDD2.n36 185
R1395 VDD2.n52 VDD2.n51 185
R1396 VDD2.n50 VDD2.n49 185
R1397 VDD2.n41 VDD2.n40 185
R1398 VDD2.n44 VDD2.n43 185
R1399 VDD2.n11 VDD2.n10 185
R1400 VDD2.n8 VDD2.n7 185
R1401 VDD2.n17 VDD2.n16 185
R1402 VDD2.n19 VDD2.n18 185
R1403 VDD2.n4 VDD2.n3 185
R1404 VDD2.n25 VDD2.n24 185
R1405 VDD2.n27 VDD2.n26 185
R1406 VDD2.t3 VDD2.n42 147.661
R1407 VDD2.t5 VDD2.n9 147.661
R1408 VDD2.n59 VDD2.n58 104.615
R1409 VDD2.n58 VDD2.n36 104.615
R1410 VDD2.n51 VDD2.n36 104.615
R1411 VDD2.n51 VDD2.n50 104.615
R1412 VDD2.n50 VDD2.n40 104.615
R1413 VDD2.n43 VDD2.n40 104.615
R1414 VDD2.n10 VDD2.n7 104.615
R1415 VDD2.n17 VDD2.n7 104.615
R1416 VDD2.n18 VDD2.n17 104.615
R1417 VDD2.n18 VDD2.n3 104.615
R1418 VDD2.n25 VDD2.n3 104.615
R1419 VDD2.n26 VDD2.n25 104.615
R1420 VDD2.n32 VDD2.n31 65.6981
R1421 VDD2 VDD2.n65 65.6952
R1422 VDD2.n43 VDD2.t3 52.3082
R1423 VDD2.n10 VDD2.t5 52.3082
R1424 VDD2.n32 VDD2.n30 48.3759
R1425 VDD2.n64 VDD2.n63 46.9247
R1426 VDD2.n64 VDD2.n32 35.3295
R1427 VDD2.n44 VDD2.n42 15.6674
R1428 VDD2.n11 VDD2.n9 15.6674
R1429 VDD2.n45 VDD2.n41 12.8005
R1430 VDD2.n12 VDD2.n8 12.8005
R1431 VDD2.n49 VDD2.n48 12.0247
R1432 VDD2.n16 VDD2.n15 12.0247
R1433 VDD2.n52 VDD2.n39 11.249
R1434 VDD2.n19 VDD2.n6 11.249
R1435 VDD2.n53 VDD2.n37 10.4732
R1436 VDD2.n20 VDD2.n4 10.4732
R1437 VDD2.n57 VDD2.n56 9.69747
R1438 VDD2.n24 VDD2.n23 9.69747
R1439 VDD2.n63 VDD2.n62 9.45567
R1440 VDD2.n30 VDD2.n29 9.45567
R1441 VDD2.n62 VDD2.n61 9.3005
R1442 VDD2.n35 VDD2.n34 9.3005
R1443 VDD2.n56 VDD2.n55 9.3005
R1444 VDD2.n54 VDD2.n53 9.3005
R1445 VDD2.n39 VDD2.n38 9.3005
R1446 VDD2.n48 VDD2.n47 9.3005
R1447 VDD2.n46 VDD2.n45 9.3005
R1448 VDD2.n29 VDD2.n28 9.3005
R1449 VDD2.n2 VDD2.n1 9.3005
R1450 VDD2.n23 VDD2.n22 9.3005
R1451 VDD2.n21 VDD2.n20 9.3005
R1452 VDD2.n6 VDD2.n5 9.3005
R1453 VDD2.n15 VDD2.n14 9.3005
R1454 VDD2.n13 VDD2.n12 9.3005
R1455 VDD2.n60 VDD2.n35 8.92171
R1456 VDD2.n27 VDD2.n2 8.92171
R1457 VDD2.n61 VDD2.n33 8.14595
R1458 VDD2.n28 VDD2.n0 8.14595
R1459 VDD2.n63 VDD2.n33 5.81868
R1460 VDD2.n30 VDD2.n0 5.81868
R1461 VDD2.n61 VDD2.n60 5.04292
R1462 VDD2.n28 VDD2.n27 5.04292
R1463 VDD2.n46 VDD2.n42 4.38594
R1464 VDD2.n13 VDD2.n9 4.38594
R1465 VDD2.n57 VDD2.n35 4.26717
R1466 VDD2.n24 VDD2.n2 4.26717
R1467 VDD2.n56 VDD2.n37 3.49141
R1468 VDD2.n23 VDD2.n4 3.49141
R1469 VDD2.n65 VDD2.t4 3.35643
R1470 VDD2.n65 VDD2.t2 3.35643
R1471 VDD2.n31 VDD2.t1 3.35643
R1472 VDD2.n31 VDD2.t0 3.35643
R1473 VDD2.n53 VDD2.n52 2.71565
R1474 VDD2.n20 VDD2.n19 2.71565
R1475 VDD2.n49 VDD2.n39 1.93989
R1476 VDD2.n16 VDD2.n6 1.93989
R1477 VDD2 VDD2.n64 1.56516
R1478 VDD2.n48 VDD2.n41 1.16414
R1479 VDD2.n15 VDD2.n8 1.16414
R1480 VDD2.n45 VDD2.n44 0.388379
R1481 VDD2.n12 VDD2.n11 0.388379
R1482 VDD2.n62 VDD2.n34 0.155672
R1483 VDD2.n55 VDD2.n34 0.155672
R1484 VDD2.n55 VDD2.n54 0.155672
R1485 VDD2.n54 VDD2.n38 0.155672
R1486 VDD2.n47 VDD2.n38 0.155672
R1487 VDD2.n47 VDD2.n46 0.155672
R1488 VDD2.n14 VDD2.n13 0.155672
R1489 VDD2.n14 VDD2.n5 0.155672
R1490 VDD2.n21 VDD2.n5 0.155672
R1491 VDD2.n22 VDD2.n21 0.155672
R1492 VDD2.n22 VDD2.n1 0.155672
R1493 VDD2.n29 VDD2.n1 0.155672
R1494 VP.n10 VP.n9 161.3
R1495 VP.n11 VP.n6 161.3
R1496 VP.n13 VP.n12 161.3
R1497 VP.n14 VP.n5 161.3
R1498 VP.n31 VP.n0 161.3
R1499 VP.n30 VP.n29 161.3
R1500 VP.n28 VP.n1 161.3
R1501 VP.n27 VP.n26 161.3
R1502 VP.n25 VP.n2 161.3
R1503 VP.n24 VP.n23 161.3
R1504 VP.n22 VP.n3 161.3
R1505 VP.n21 VP.n20 161.3
R1506 VP.n19 VP.n4 161.3
R1507 VP.n7 VP.t2 104.612
R1508 VP.n18 VP.n17 94.6776
R1509 VP.n33 VP.n32 94.6776
R1510 VP.n16 VP.n15 94.6776
R1511 VP.n25 VP.t5 71.0955
R1512 VP.n18 VP.t3 71.0955
R1513 VP.n32 VP.t1 71.0955
R1514 VP.n15 VP.t0 71.0955
R1515 VP.n8 VP.t4 71.0955
R1516 VP.n20 VP.n3 56.5617
R1517 VP.n30 VP.n1 56.5617
R1518 VP.n13 VP.n6 56.5617
R1519 VP.n8 VP.n7 45.8151
R1520 VP.n17 VP.n16 41.6701
R1521 VP.n20 VP.n19 24.5923
R1522 VP.n24 VP.n3 24.5923
R1523 VP.n25 VP.n24 24.5923
R1524 VP.n26 VP.n25 24.5923
R1525 VP.n26 VP.n1 24.5923
R1526 VP.n31 VP.n30 24.5923
R1527 VP.n14 VP.n13 24.5923
R1528 VP.n9 VP.n8 24.5923
R1529 VP.n9 VP.n6 24.5923
R1530 VP.n19 VP.n18 16.2311
R1531 VP.n32 VP.n31 16.2311
R1532 VP.n15 VP.n14 16.2311
R1533 VP.n10 VP.n7 9.3086
R1534 VP.n16 VP.n5 0.278335
R1535 VP.n17 VP.n4 0.278335
R1536 VP.n33 VP.n0 0.278335
R1537 VP.n11 VP.n10 0.189894
R1538 VP.n12 VP.n11 0.189894
R1539 VP.n12 VP.n5 0.189894
R1540 VP.n21 VP.n4 0.189894
R1541 VP.n22 VP.n21 0.189894
R1542 VP.n23 VP.n22 0.189894
R1543 VP.n23 VP.n2 0.189894
R1544 VP.n27 VP.n2 0.189894
R1545 VP.n28 VP.n27 0.189894
R1546 VP.n29 VP.n28 0.189894
R1547 VP.n29 VP.n0 0.189894
R1548 VP VP.n33 0.153485
R1549 VDD1.n26 VDD1.n0 289.615
R1550 VDD1.n57 VDD1.n31 289.615
R1551 VDD1.n27 VDD1.n26 185
R1552 VDD1.n25 VDD1.n24 185
R1553 VDD1.n4 VDD1.n3 185
R1554 VDD1.n19 VDD1.n18 185
R1555 VDD1.n17 VDD1.n16 185
R1556 VDD1.n8 VDD1.n7 185
R1557 VDD1.n11 VDD1.n10 185
R1558 VDD1.n42 VDD1.n41 185
R1559 VDD1.n39 VDD1.n38 185
R1560 VDD1.n48 VDD1.n47 185
R1561 VDD1.n50 VDD1.n49 185
R1562 VDD1.n35 VDD1.n34 185
R1563 VDD1.n56 VDD1.n55 185
R1564 VDD1.n58 VDD1.n57 185
R1565 VDD1.t3 VDD1.n9 147.661
R1566 VDD1.t2 VDD1.n40 147.661
R1567 VDD1.n26 VDD1.n25 104.615
R1568 VDD1.n25 VDD1.n3 104.615
R1569 VDD1.n18 VDD1.n3 104.615
R1570 VDD1.n18 VDD1.n17 104.615
R1571 VDD1.n17 VDD1.n7 104.615
R1572 VDD1.n10 VDD1.n7 104.615
R1573 VDD1.n41 VDD1.n38 104.615
R1574 VDD1.n48 VDD1.n38 104.615
R1575 VDD1.n49 VDD1.n48 104.615
R1576 VDD1.n49 VDD1.n34 104.615
R1577 VDD1.n56 VDD1.n34 104.615
R1578 VDD1.n57 VDD1.n56 104.615
R1579 VDD1.n63 VDD1.n62 65.6981
R1580 VDD1.n65 VDD1.n64 65.2513
R1581 VDD1.n10 VDD1.t3 52.3082
R1582 VDD1.n41 VDD1.t2 52.3082
R1583 VDD1 VDD1.n30 48.4894
R1584 VDD1.n63 VDD1.n61 48.3759
R1585 VDD1.n65 VDD1.n63 36.9168
R1586 VDD1.n11 VDD1.n9 15.6674
R1587 VDD1.n42 VDD1.n40 15.6674
R1588 VDD1.n12 VDD1.n8 12.8005
R1589 VDD1.n43 VDD1.n39 12.8005
R1590 VDD1.n16 VDD1.n15 12.0247
R1591 VDD1.n47 VDD1.n46 12.0247
R1592 VDD1.n19 VDD1.n6 11.249
R1593 VDD1.n50 VDD1.n37 11.249
R1594 VDD1.n20 VDD1.n4 10.4732
R1595 VDD1.n51 VDD1.n35 10.4732
R1596 VDD1.n24 VDD1.n23 9.69747
R1597 VDD1.n55 VDD1.n54 9.69747
R1598 VDD1.n30 VDD1.n29 9.45567
R1599 VDD1.n61 VDD1.n60 9.45567
R1600 VDD1.n29 VDD1.n28 9.3005
R1601 VDD1.n2 VDD1.n1 9.3005
R1602 VDD1.n23 VDD1.n22 9.3005
R1603 VDD1.n21 VDD1.n20 9.3005
R1604 VDD1.n6 VDD1.n5 9.3005
R1605 VDD1.n15 VDD1.n14 9.3005
R1606 VDD1.n13 VDD1.n12 9.3005
R1607 VDD1.n60 VDD1.n59 9.3005
R1608 VDD1.n33 VDD1.n32 9.3005
R1609 VDD1.n54 VDD1.n53 9.3005
R1610 VDD1.n52 VDD1.n51 9.3005
R1611 VDD1.n37 VDD1.n36 9.3005
R1612 VDD1.n46 VDD1.n45 9.3005
R1613 VDD1.n44 VDD1.n43 9.3005
R1614 VDD1.n27 VDD1.n2 8.92171
R1615 VDD1.n58 VDD1.n33 8.92171
R1616 VDD1.n28 VDD1.n0 8.14595
R1617 VDD1.n59 VDD1.n31 8.14595
R1618 VDD1.n30 VDD1.n0 5.81868
R1619 VDD1.n61 VDD1.n31 5.81868
R1620 VDD1.n28 VDD1.n27 5.04292
R1621 VDD1.n59 VDD1.n58 5.04292
R1622 VDD1.n13 VDD1.n9 4.38594
R1623 VDD1.n44 VDD1.n40 4.38594
R1624 VDD1.n24 VDD1.n2 4.26717
R1625 VDD1.n55 VDD1.n33 4.26717
R1626 VDD1.n23 VDD1.n4 3.49141
R1627 VDD1.n54 VDD1.n35 3.49141
R1628 VDD1.n64 VDD1.t1 3.35643
R1629 VDD1.n64 VDD1.t5 3.35643
R1630 VDD1.n62 VDD1.t0 3.35643
R1631 VDD1.n62 VDD1.t4 3.35643
R1632 VDD1.n20 VDD1.n19 2.71565
R1633 VDD1.n51 VDD1.n50 2.71565
R1634 VDD1.n16 VDD1.n6 1.93989
R1635 VDD1.n47 VDD1.n37 1.93989
R1636 VDD1.n15 VDD1.n8 1.16414
R1637 VDD1.n46 VDD1.n39 1.16414
R1638 VDD1 VDD1.n65 0.444466
R1639 VDD1.n12 VDD1.n11 0.388379
R1640 VDD1.n43 VDD1.n42 0.388379
R1641 VDD1.n29 VDD1.n1 0.155672
R1642 VDD1.n22 VDD1.n1 0.155672
R1643 VDD1.n22 VDD1.n21 0.155672
R1644 VDD1.n21 VDD1.n5 0.155672
R1645 VDD1.n14 VDD1.n5 0.155672
R1646 VDD1.n14 VDD1.n13 0.155672
R1647 VDD1.n45 VDD1.n44 0.155672
R1648 VDD1.n45 VDD1.n36 0.155672
R1649 VDD1.n52 VDD1.n36 0.155672
R1650 VDD1.n53 VDD1.n52 0.155672
R1651 VDD1.n53 VDD1.n32 0.155672
R1652 VDD1.n60 VDD1.n32 0.155672
C0 VTAIL VDD1 5.27321f
C1 VDD2 VP 0.407306f
C2 VP VN 5.21386f
C3 VP VTAIL 3.72395f
C4 VP VDD1 3.56942f
C5 VDD2 VN 3.31455f
C6 VDD2 VTAIL 5.32105f
C7 VN VTAIL 3.70972f
C8 VDD2 VDD1 1.18445f
C9 VN VDD1 0.150316f
C10 VDD2 B 4.42688f
C11 VDD1 B 4.524248f
C12 VTAIL B 4.754739f
C13 VN B 10.534949f
C14 VP B 9.162529f
C15 VDD1.n0 B 0.029926f
C16 VDD1.n1 B 0.022364f
C17 VDD1.n2 B 0.012017f
C18 VDD1.n3 B 0.028405f
C19 VDD1.n4 B 0.012724f
C20 VDD1.n5 B 0.022364f
C21 VDD1.n6 B 0.012017f
C22 VDD1.n7 B 0.028405f
C23 VDD1.n8 B 0.012724f
C24 VDD1.n9 B 0.095081f
C25 VDD1.t3 B 0.04626f
C26 VDD1.n10 B 0.021303f
C27 VDD1.n11 B 0.016778f
C28 VDD1.n12 B 0.012017f
C29 VDD1.n13 B 0.521964f
C30 VDD1.n14 B 0.022364f
C31 VDD1.n15 B 0.012017f
C32 VDD1.n16 B 0.012724f
C33 VDD1.n17 B 0.028405f
C34 VDD1.n18 B 0.028405f
C35 VDD1.n19 B 0.012724f
C36 VDD1.n20 B 0.012017f
C37 VDD1.n21 B 0.022364f
C38 VDD1.n22 B 0.022364f
C39 VDD1.n23 B 0.012017f
C40 VDD1.n24 B 0.012724f
C41 VDD1.n25 B 0.028405f
C42 VDD1.n26 B 0.058823f
C43 VDD1.n27 B 0.012724f
C44 VDD1.n28 B 0.012017f
C45 VDD1.n29 B 0.048638f
C46 VDD1.n30 B 0.052982f
C47 VDD1.n31 B 0.029926f
C48 VDD1.n32 B 0.022364f
C49 VDD1.n33 B 0.012017f
C50 VDD1.n34 B 0.028405f
C51 VDD1.n35 B 0.012724f
C52 VDD1.n36 B 0.022364f
C53 VDD1.n37 B 0.012017f
C54 VDD1.n38 B 0.028405f
C55 VDD1.n39 B 0.012724f
C56 VDD1.n40 B 0.095081f
C57 VDD1.t2 B 0.04626f
C58 VDD1.n41 B 0.021303f
C59 VDD1.n42 B 0.016778f
C60 VDD1.n43 B 0.012017f
C61 VDD1.n44 B 0.521964f
C62 VDD1.n45 B 0.022364f
C63 VDD1.n46 B 0.012017f
C64 VDD1.n47 B 0.012724f
C65 VDD1.n48 B 0.028405f
C66 VDD1.n49 B 0.028405f
C67 VDD1.n50 B 0.012724f
C68 VDD1.n51 B 0.012017f
C69 VDD1.n52 B 0.022364f
C70 VDD1.n53 B 0.022364f
C71 VDD1.n54 B 0.012017f
C72 VDD1.n55 B 0.012724f
C73 VDD1.n56 B 0.028405f
C74 VDD1.n57 B 0.058823f
C75 VDD1.n58 B 0.012724f
C76 VDD1.n59 B 0.012017f
C77 VDD1.n60 B 0.048638f
C78 VDD1.n61 B 0.052398f
C79 VDD1.t0 B 0.104268f
C80 VDD1.t4 B 0.104268f
C81 VDD1.n62 B 0.869643f
C82 VDD1.n63 B 1.92375f
C83 VDD1.t1 B 0.104268f
C84 VDD1.t5 B 0.104268f
C85 VDD1.n64 B 0.867134f
C86 VDD1.n65 B 1.91702f
C87 VP.n0 B 0.040649f
C88 VP.t1 B 0.962053f
C89 VP.n1 B 0.037571f
C90 VP.n2 B 0.030834f
C91 VP.t5 B 0.962053f
C92 VP.n3 B 0.037571f
C93 VP.n4 B 0.040649f
C94 VP.t3 B 0.962053f
C95 VP.n5 B 0.040649f
C96 VP.t0 B 0.962053f
C97 VP.n6 B 0.037571f
C98 VP.t2 B 1.1299f
C99 VP.n7 B 0.432106f
C100 VP.t4 B 0.962053f
C101 VP.n8 B 0.457484f
C102 VP.n9 B 0.057179f
C103 VP.n10 B 0.256624f
C104 VP.n11 B 0.030834f
C105 VP.n12 B 0.030834f
C106 VP.n13 B 0.052074f
C107 VP.n14 B 0.047582f
C108 VP.n15 B 0.455638f
C109 VP.n16 B 1.28408f
C110 VP.n17 B 1.31075f
C111 VP.n18 B 0.455638f
C112 VP.n19 B 0.047582f
C113 VP.n20 B 0.052074f
C114 VP.n21 B 0.030834f
C115 VP.n22 B 0.030834f
C116 VP.n23 B 0.030834f
C117 VP.n24 B 0.057179f
C118 VP.n25 B 0.397066f
C119 VP.n26 B 0.057179f
C120 VP.n27 B 0.030834f
C121 VP.n28 B 0.030834f
C122 VP.n29 B 0.030834f
C123 VP.n30 B 0.052074f
C124 VP.n31 B 0.047582f
C125 VP.n32 B 0.455638f
C126 VP.n33 B 0.040412f
C127 VDD2.n0 B 0.029188f
C128 VDD2.n1 B 0.021812f
C129 VDD2.n2 B 0.011721f
C130 VDD2.n3 B 0.027704f
C131 VDD2.n4 B 0.01241f
C132 VDD2.n5 B 0.021812f
C133 VDD2.n6 B 0.011721f
C134 VDD2.n7 B 0.027704f
C135 VDD2.n8 B 0.01241f
C136 VDD2.n9 B 0.092737f
C137 VDD2.t5 B 0.045119f
C138 VDD2.n10 B 0.020778f
C139 VDD2.n11 B 0.016365f
C140 VDD2.n12 B 0.011721f
C141 VDD2.n13 B 0.509095f
C142 VDD2.n14 B 0.021812f
C143 VDD2.n15 B 0.011721f
C144 VDD2.n16 B 0.01241f
C145 VDD2.n17 B 0.027704f
C146 VDD2.n18 B 0.027704f
C147 VDD2.n19 B 0.01241f
C148 VDD2.n20 B 0.011721f
C149 VDD2.n21 B 0.021812f
C150 VDD2.n22 B 0.021812f
C151 VDD2.n23 B 0.011721f
C152 VDD2.n24 B 0.01241f
C153 VDD2.n25 B 0.027704f
C154 VDD2.n26 B 0.057373f
C155 VDD2.n27 B 0.01241f
C156 VDD2.n28 B 0.011721f
C157 VDD2.n29 B 0.047439f
C158 VDD2.n30 B 0.051106f
C159 VDD2.t1 B 0.101697f
C160 VDD2.t0 B 0.101697f
C161 VDD2.n31 B 0.848202f
C162 VDD2.n32 B 1.78576f
C163 VDD2.n33 B 0.029188f
C164 VDD2.n34 B 0.021812f
C165 VDD2.n35 B 0.011721f
C166 VDD2.n36 B 0.027704f
C167 VDD2.n37 B 0.01241f
C168 VDD2.n38 B 0.021812f
C169 VDD2.n39 B 0.011721f
C170 VDD2.n40 B 0.027704f
C171 VDD2.n41 B 0.01241f
C172 VDD2.n42 B 0.092737f
C173 VDD2.t3 B 0.045119f
C174 VDD2.n43 B 0.020778f
C175 VDD2.n44 B 0.016365f
C176 VDD2.n45 B 0.011721f
C177 VDD2.n46 B 0.509095f
C178 VDD2.n47 B 0.021812f
C179 VDD2.n48 B 0.011721f
C180 VDD2.n49 B 0.01241f
C181 VDD2.n50 B 0.027704f
C182 VDD2.n51 B 0.027704f
C183 VDD2.n52 B 0.01241f
C184 VDD2.n53 B 0.011721f
C185 VDD2.n54 B 0.021812f
C186 VDD2.n55 B 0.021812f
C187 VDD2.n56 B 0.011721f
C188 VDD2.n57 B 0.01241f
C189 VDD2.n58 B 0.027704f
C190 VDD2.n59 B 0.057373f
C191 VDD2.n60 B 0.01241f
C192 VDD2.n61 B 0.011721f
C193 VDD2.n62 B 0.047439f
C194 VDD2.n63 B 0.046827f
C195 VDD2.n64 B 1.67143f
C196 VDD2.t4 B 0.101697f
C197 VDD2.t2 B 0.101697f
C198 VDD2.n65 B 0.848177f
C199 VTAIL.t6 B 0.123044f
C200 VTAIL.t8 B 0.123044f
C201 VTAIL.n0 B 0.951301f
C202 VTAIL.n1 B 0.423775f
C203 VTAIL.n2 B 0.035314f
C204 VTAIL.n3 B 0.026391f
C205 VTAIL.n4 B 0.014181f
C206 VTAIL.n5 B 0.03352f
C207 VTAIL.n6 B 0.015016f
C208 VTAIL.n7 B 0.026391f
C209 VTAIL.n8 B 0.014181f
C210 VTAIL.n9 B 0.03352f
C211 VTAIL.n10 B 0.015016f
C212 VTAIL.n11 B 0.112203f
C213 VTAIL.t1 B 0.05459f
C214 VTAIL.n12 B 0.02514f
C215 VTAIL.n13 B 0.0198f
C216 VTAIL.n14 B 0.014181f
C217 VTAIL.n15 B 0.615958f
C218 VTAIL.n16 B 0.026391f
C219 VTAIL.n17 B 0.014181f
C220 VTAIL.n18 B 0.015016f
C221 VTAIL.n19 B 0.03352f
C222 VTAIL.n20 B 0.03352f
C223 VTAIL.n21 B 0.015016f
C224 VTAIL.n22 B 0.014181f
C225 VTAIL.n23 B 0.026391f
C226 VTAIL.n24 B 0.026391f
C227 VTAIL.n25 B 0.014181f
C228 VTAIL.n26 B 0.015016f
C229 VTAIL.n27 B 0.03352f
C230 VTAIL.n28 B 0.069416f
C231 VTAIL.n29 B 0.015016f
C232 VTAIL.n30 B 0.014181f
C233 VTAIL.n31 B 0.057396f
C234 VTAIL.n32 B 0.038403f
C235 VTAIL.n33 B 0.316674f
C236 VTAIL.t4 B 0.123044f
C237 VTAIL.t3 B 0.123044f
C238 VTAIL.n34 B 0.951301f
C239 VTAIL.n35 B 1.5542f
C240 VTAIL.t9 B 0.123044f
C241 VTAIL.t7 B 0.123044f
C242 VTAIL.n36 B 0.951308f
C243 VTAIL.n37 B 1.5542f
C244 VTAIL.n38 B 0.035314f
C245 VTAIL.n39 B 0.026391f
C246 VTAIL.n40 B 0.014181f
C247 VTAIL.n41 B 0.03352f
C248 VTAIL.n42 B 0.015016f
C249 VTAIL.n43 B 0.026391f
C250 VTAIL.n44 B 0.014181f
C251 VTAIL.n45 B 0.03352f
C252 VTAIL.n46 B 0.015016f
C253 VTAIL.n47 B 0.112203f
C254 VTAIL.t11 B 0.05459f
C255 VTAIL.n48 B 0.02514f
C256 VTAIL.n49 B 0.0198f
C257 VTAIL.n50 B 0.014181f
C258 VTAIL.n51 B 0.615958f
C259 VTAIL.n52 B 0.026391f
C260 VTAIL.n53 B 0.014181f
C261 VTAIL.n54 B 0.015016f
C262 VTAIL.n55 B 0.03352f
C263 VTAIL.n56 B 0.03352f
C264 VTAIL.n57 B 0.015016f
C265 VTAIL.n58 B 0.014181f
C266 VTAIL.n59 B 0.026391f
C267 VTAIL.n60 B 0.026391f
C268 VTAIL.n61 B 0.014181f
C269 VTAIL.n62 B 0.015016f
C270 VTAIL.n63 B 0.03352f
C271 VTAIL.n64 B 0.069416f
C272 VTAIL.n65 B 0.015016f
C273 VTAIL.n66 B 0.014181f
C274 VTAIL.n67 B 0.057396f
C275 VTAIL.n68 B 0.038403f
C276 VTAIL.n69 B 0.316674f
C277 VTAIL.t5 B 0.123044f
C278 VTAIL.t0 B 0.123044f
C279 VTAIL.n70 B 0.951308f
C280 VTAIL.n71 B 0.546926f
C281 VTAIL.n72 B 0.035314f
C282 VTAIL.n73 B 0.026391f
C283 VTAIL.n74 B 0.014181f
C284 VTAIL.n75 B 0.03352f
C285 VTAIL.n76 B 0.015016f
C286 VTAIL.n77 B 0.026391f
C287 VTAIL.n78 B 0.014181f
C288 VTAIL.n79 B 0.03352f
C289 VTAIL.n80 B 0.015016f
C290 VTAIL.n81 B 0.112203f
C291 VTAIL.t2 B 0.05459f
C292 VTAIL.n82 B 0.02514f
C293 VTAIL.n83 B 0.0198f
C294 VTAIL.n84 B 0.014181f
C295 VTAIL.n85 B 0.615958f
C296 VTAIL.n86 B 0.026391f
C297 VTAIL.n87 B 0.014181f
C298 VTAIL.n88 B 0.015016f
C299 VTAIL.n89 B 0.03352f
C300 VTAIL.n90 B 0.03352f
C301 VTAIL.n91 B 0.015016f
C302 VTAIL.n92 B 0.014181f
C303 VTAIL.n93 B 0.026391f
C304 VTAIL.n94 B 0.026391f
C305 VTAIL.n95 B 0.014181f
C306 VTAIL.n96 B 0.015016f
C307 VTAIL.n97 B 0.03352f
C308 VTAIL.n98 B 0.069416f
C309 VTAIL.n99 B 0.015016f
C310 VTAIL.n100 B 0.014181f
C311 VTAIL.n101 B 0.057396f
C312 VTAIL.n102 B 0.038403f
C313 VTAIL.n103 B 1.15314f
C314 VTAIL.n104 B 0.035314f
C315 VTAIL.n105 B 0.026391f
C316 VTAIL.n106 B 0.014181f
C317 VTAIL.n107 B 0.03352f
C318 VTAIL.n108 B 0.015016f
C319 VTAIL.n109 B 0.026391f
C320 VTAIL.n110 B 0.014181f
C321 VTAIL.n111 B 0.03352f
C322 VTAIL.n112 B 0.015016f
C323 VTAIL.n113 B 0.112203f
C324 VTAIL.t10 B 0.05459f
C325 VTAIL.n114 B 0.02514f
C326 VTAIL.n115 B 0.0198f
C327 VTAIL.n116 B 0.014181f
C328 VTAIL.n117 B 0.615958f
C329 VTAIL.n118 B 0.026391f
C330 VTAIL.n119 B 0.014181f
C331 VTAIL.n120 B 0.015016f
C332 VTAIL.n121 B 0.03352f
C333 VTAIL.n122 B 0.03352f
C334 VTAIL.n123 B 0.015016f
C335 VTAIL.n124 B 0.014181f
C336 VTAIL.n125 B 0.026391f
C337 VTAIL.n126 B 0.026391f
C338 VTAIL.n127 B 0.014181f
C339 VTAIL.n128 B 0.015016f
C340 VTAIL.n129 B 0.03352f
C341 VTAIL.n130 B 0.069416f
C342 VTAIL.n131 B 0.015016f
C343 VTAIL.n132 B 0.014181f
C344 VTAIL.n133 B 0.057396f
C345 VTAIL.n134 B 0.038403f
C346 VTAIL.n135 B 1.10549f
C347 VN.n0 B 0.039537f
C348 VN.t5 B 0.935719f
C349 VN.n1 B 0.036543f
C350 VN.t0 B 1.09897f
C351 VN.n2 B 0.420278f
C352 VN.t4 B 0.935719f
C353 VN.n3 B 0.444961f
C354 VN.n4 B 0.055614f
C355 VN.n5 B 0.249599f
C356 VN.n6 B 0.02999f
C357 VN.n7 B 0.02999f
C358 VN.n8 B 0.050648f
C359 VN.n9 B 0.046279f
C360 VN.n10 B 0.443167f
C361 VN.n11 B 0.039306f
C362 VN.n12 B 0.039537f
C363 VN.t2 B 0.935719f
C364 VN.n13 B 0.036543f
C365 VN.t3 B 1.09897f
C366 VN.n14 B 0.420278f
C367 VN.t1 B 0.935719f
C368 VN.n15 B 0.444961f
C369 VN.n16 B 0.055614f
C370 VN.n17 B 0.249599f
C371 VN.n18 B 0.02999f
C372 VN.n19 B 0.02999f
C373 VN.n20 B 0.050648f
C374 VN.n21 B 0.046279f
C375 VN.n22 B 0.443167f
C376 VN.n23 B 1.26556f
.ends

