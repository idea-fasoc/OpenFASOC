* NGSPICE file created from diff_pair_sample_0182.ext - technology: sky130A

.subckt diff_pair_sample_0182 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=0 ps=0 w=17.53 l=2.75
X1 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=6.8367 ps=35.84 w=17.53 l=2.75
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=0 ps=0 w=17.53 l=2.75
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=6.8367 ps=35.84 w=17.53 l=2.75
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=6.8367 ps=35.84 w=17.53 l=2.75
X5 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=6.8367 ps=35.84 w=17.53 l=2.75
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=0 ps=0 w=17.53 l=2.75
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8367 pd=35.84 as=0 ps=0 w=17.53 l=2.75
R0 B.n598 B.n597 585
R1 B.n598 B.n50 585
R2 B.n601 B.n600 585
R3 B.n602 B.n117 585
R4 B.n604 B.n603 585
R5 B.n606 B.n116 585
R6 B.n609 B.n608 585
R7 B.n610 B.n115 585
R8 B.n612 B.n611 585
R9 B.n614 B.n114 585
R10 B.n617 B.n616 585
R11 B.n618 B.n113 585
R12 B.n620 B.n619 585
R13 B.n622 B.n112 585
R14 B.n625 B.n624 585
R15 B.n626 B.n111 585
R16 B.n628 B.n627 585
R17 B.n630 B.n110 585
R18 B.n633 B.n632 585
R19 B.n634 B.n109 585
R20 B.n636 B.n635 585
R21 B.n638 B.n108 585
R22 B.n641 B.n640 585
R23 B.n642 B.n107 585
R24 B.n644 B.n643 585
R25 B.n646 B.n106 585
R26 B.n649 B.n648 585
R27 B.n650 B.n105 585
R28 B.n652 B.n651 585
R29 B.n654 B.n104 585
R30 B.n657 B.n656 585
R31 B.n658 B.n103 585
R32 B.n660 B.n659 585
R33 B.n662 B.n102 585
R34 B.n665 B.n664 585
R35 B.n666 B.n101 585
R36 B.n668 B.n667 585
R37 B.n670 B.n100 585
R38 B.n673 B.n672 585
R39 B.n674 B.n99 585
R40 B.n676 B.n675 585
R41 B.n678 B.n98 585
R42 B.n681 B.n680 585
R43 B.n682 B.n97 585
R44 B.n684 B.n683 585
R45 B.n686 B.n96 585
R46 B.n689 B.n688 585
R47 B.n690 B.n95 585
R48 B.n692 B.n691 585
R49 B.n694 B.n94 585
R50 B.n697 B.n696 585
R51 B.n698 B.n93 585
R52 B.n700 B.n699 585
R53 B.n702 B.n92 585
R54 B.n705 B.n704 585
R55 B.n706 B.n91 585
R56 B.n708 B.n707 585
R57 B.n710 B.n90 585
R58 B.n713 B.n712 585
R59 B.n715 B.n87 585
R60 B.n717 B.n716 585
R61 B.n719 B.n86 585
R62 B.n722 B.n721 585
R63 B.n723 B.n85 585
R64 B.n725 B.n724 585
R65 B.n727 B.n84 585
R66 B.n729 B.n728 585
R67 B.n731 B.n730 585
R68 B.n734 B.n733 585
R69 B.n735 B.n79 585
R70 B.n737 B.n736 585
R71 B.n739 B.n78 585
R72 B.n742 B.n741 585
R73 B.n743 B.n77 585
R74 B.n745 B.n744 585
R75 B.n747 B.n76 585
R76 B.n750 B.n749 585
R77 B.n751 B.n75 585
R78 B.n753 B.n752 585
R79 B.n755 B.n74 585
R80 B.n758 B.n757 585
R81 B.n759 B.n73 585
R82 B.n761 B.n760 585
R83 B.n763 B.n72 585
R84 B.n766 B.n765 585
R85 B.n767 B.n71 585
R86 B.n769 B.n768 585
R87 B.n771 B.n70 585
R88 B.n774 B.n773 585
R89 B.n775 B.n69 585
R90 B.n777 B.n776 585
R91 B.n779 B.n68 585
R92 B.n782 B.n781 585
R93 B.n783 B.n67 585
R94 B.n785 B.n784 585
R95 B.n787 B.n66 585
R96 B.n790 B.n789 585
R97 B.n791 B.n65 585
R98 B.n793 B.n792 585
R99 B.n795 B.n64 585
R100 B.n798 B.n797 585
R101 B.n799 B.n63 585
R102 B.n801 B.n800 585
R103 B.n803 B.n62 585
R104 B.n806 B.n805 585
R105 B.n807 B.n61 585
R106 B.n809 B.n808 585
R107 B.n811 B.n60 585
R108 B.n814 B.n813 585
R109 B.n815 B.n59 585
R110 B.n817 B.n816 585
R111 B.n819 B.n58 585
R112 B.n822 B.n821 585
R113 B.n823 B.n57 585
R114 B.n825 B.n824 585
R115 B.n827 B.n56 585
R116 B.n830 B.n829 585
R117 B.n831 B.n55 585
R118 B.n833 B.n832 585
R119 B.n835 B.n54 585
R120 B.n838 B.n837 585
R121 B.n839 B.n53 585
R122 B.n841 B.n840 585
R123 B.n843 B.n52 585
R124 B.n846 B.n845 585
R125 B.n847 B.n51 585
R126 B.n596 B.n49 585
R127 B.n850 B.n49 585
R128 B.n595 B.n48 585
R129 B.n851 B.n48 585
R130 B.n594 B.n47 585
R131 B.n852 B.n47 585
R132 B.n593 B.n592 585
R133 B.n592 B.n43 585
R134 B.n591 B.n42 585
R135 B.n858 B.n42 585
R136 B.n590 B.n41 585
R137 B.n859 B.n41 585
R138 B.n589 B.n40 585
R139 B.n860 B.n40 585
R140 B.n588 B.n587 585
R141 B.n587 B.n39 585
R142 B.n586 B.n35 585
R143 B.n866 B.n35 585
R144 B.n585 B.n34 585
R145 B.n867 B.n34 585
R146 B.n584 B.n33 585
R147 B.n868 B.n33 585
R148 B.n583 B.n582 585
R149 B.n582 B.n29 585
R150 B.n581 B.n28 585
R151 B.n874 B.n28 585
R152 B.n580 B.n27 585
R153 B.n875 B.n27 585
R154 B.n579 B.n26 585
R155 B.n876 B.n26 585
R156 B.n578 B.n577 585
R157 B.n577 B.n22 585
R158 B.n576 B.n21 585
R159 B.n882 B.n21 585
R160 B.n575 B.n20 585
R161 B.n883 B.n20 585
R162 B.n574 B.n19 585
R163 B.n884 B.n19 585
R164 B.n573 B.n572 585
R165 B.n572 B.n18 585
R166 B.n571 B.n14 585
R167 B.n890 B.n14 585
R168 B.n570 B.n13 585
R169 B.n891 B.n13 585
R170 B.n569 B.n12 585
R171 B.n892 B.n12 585
R172 B.n568 B.n567 585
R173 B.n567 B.n8 585
R174 B.n566 B.n7 585
R175 B.n898 B.n7 585
R176 B.n565 B.n6 585
R177 B.n899 B.n6 585
R178 B.n564 B.n5 585
R179 B.n900 B.n5 585
R180 B.n563 B.n562 585
R181 B.n562 B.n4 585
R182 B.n561 B.n118 585
R183 B.n561 B.n560 585
R184 B.n551 B.n119 585
R185 B.n120 B.n119 585
R186 B.n553 B.n552 585
R187 B.n554 B.n553 585
R188 B.n550 B.n125 585
R189 B.n125 B.n124 585
R190 B.n549 B.n548 585
R191 B.n548 B.n547 585
R192 B.n127 B.n126 585
R193 B.n540 B.n127 585
R194 B.n539 B.n538 585
R195 B.n541 B.n539 585
R196 B.n537 B.n132 585
R197 B.n132 B.n131 585
R198 B.n536 B.n535 585
R199 B.n535 B.n534 585
R200 B.n134 B.n133 585
R201 B.n135 B.n134 585
R202 B.n527 B.n526 585
R203 B.n528 B.n527 585
R204 B.n525 B.n140 585
R205 B.n140 B.n139 585
R206 B.n524 B.n523 585
R207 B.n523 B.n522 585
R208 B.n142 B.n141 585
R209 B.n143 B.n142 585
R210 B.n515 B.n514 585
R211 B.n516 B.n515 585
R212 B.n513 B.n148 585
R213 B.n148 B.n147 585
R214 B.n512 B.n511 585
R215 B.n511 B.n510 585
R216 B.n150 B.n149 585
R217 B.n503 B.n150 585
R218 B.n502 B.n501 585
R219 B.n504 B.n502 585
R220 B.n500 B.n155 585
R221 B.n155 B.n154 585
R222 B.n499 B.n498 585
R223 B.n498 B.n497 585
R224 B.n157 B.n156 585
R225 B.n158 B.n157 585
R226 B.n490 B.n489 585
R227 B.n491 B.n490 585
R228 B.n488 B.n163 585
R229 B.n163 B.n162 585
R230 B.n487 B.n486 585
R231 B.n486 B.n485 585
R232 B.n482 B.n167 585
R233 B.n481 B.n480 585
R234 B.n478 B.n168 585
R235 B.n478 B.n166 585
R236 B.n477 B.n476 585
R237 B.n475 B.n474 585
R238 B.n473 B.n170 585
R239 B.n471 B.n470 585
R240 B.n469 B.n171 585
R241 B.n468 B.n467 585
R242 B.n465 B.n172 585
R243 B.n463 B.n462 585
R244 B.n461 B.n173 585
R245 B.n460 B.n459 585
R246 B.n457 B.n174 585
R247 B.n455 B.n454 585
R248 B.n453 B.n175 585
R249 B.n452 B.n451 585
R250 B.n449 B.n176 585
R251 B.n447 B.n446 585
R252 B.n445 B.n177 585
R253 B.n444 B.n443 585
R254 B.n441 B.n178 585
R255 B.n439 B.n438 585
R256 B.n437 B.n179 585
R257 B.n436 B.n435 585
R258 B.n433 B.n180 585
R259 B.n431 B.n430 585
R260 B.n429 B.n181 585
R261 B.n428 B.n427 585
R262 B.n425 B.n182 585
R263 B.n423 B.n422 585
R264 B.n421 B.n183 585
R265 B.n420 B.n419 585
R266 B.n417 B.n184 585
R267 B.n415 B.n414 585
R268 B.n413 B.n185 585
R269 B.n412 B.n411 585
R270 B.n409 B.n186 585
R271 B.n407 B.n406 585
R272 B.n405 B.n187 585
R273 B.n404 B.n403 585
R274 B.n401 B.n188 585
R275 B.n399 B.n398 585
R276 B.n397 B.n189 585
R277 B.n396 B.n395 585
R278 B.n393 B.n190 585
R279 B.n391 B.n390 585
R280 B.n389 B.n191 585
R281 B.n388 B.n387 585
R282 B.n385 B.n192 585
R283 B.n383 B.n382 585
R284 B.n381 B.n193 585
R285 B.n380 B.n379 585
R286 B.n377 B.n194 585
R287 B.n375 B.n374 585
R288 B.n373 B.n195 585
R289 B.n372 B.n371 585
R290 B.n369 B.n196 585
R291 B.n367 B.n366 585
R292 B.n365 B.n197 585
R293 B.n364 B.n363 585
R294 B.n361 B.n201 585
R295 B.n359 B.n358 585
R296 B.n357 B.n202 585
R297 B.n356 B.n355 585
R298 B.n353 B.n203 585
R299 B.n351 B.n350 585
R300 B.n348 B.n204 585
R301 B.n347 B.n346 585
R302 B.n344 B.n207 585
R303 B.n342 B.n341 585
R304 B.n340 B.n208 585
R305 B.n339 B.n338 585
R306 B.n336 B.n209 585
R307 B.n334 B.n333 585
R308 B.n332 B.n210 585
R309 B.n331 B.n330 585
R310 B.n328 B.n211 585
R311 B.n326 B.n325 585
R312 B.n324 B.n212 585
R313 B.n323 B.n322 585
R314 B.n320 B.n213 585
R315 B.n318 B.n317 585
R316 B.n316 B.n214 585
R317 B.n315 B.n314 585
R318 B.n312 B.n215 585
R319 B.n310 B.n309 585
R320 B.n308 B.n216 585
R321 B.n307 B.n306 585
R322 B.n304 B.n217 585
R323 B.n302 B.n301 585
R324 B.n300 B.n218 585
R325 B.n299 B.n298 585
R326 B.n296 B.n219 585
R327 B.n294 B.n293 585
R328 B.n292 B.n220 585
R329 B.n291 B.n290 585
R330 B.n288 B.n221 585
R331 B.n286 B.n285 585
R332 B.n284 B.n222 585
R333 B.n283 B.n282 585
R334 B.n280 B.n223 585
R335 B.n278 B.n277 585
R336 B.n276 B.n224 585
R337 B.n275 B.n274 585
R338 B.n272 B.n225 585
R339 B.n270 B.n269 585
R340 B.n268 B.n226 585
R341 B.n267 B.n266 585
R342 B.n264 B.n227 585
R343 B.n262 B.n261 585
R344 B.n260 B.n228 585
R345 B.n259 B.n258 585
R346 B.n256 B.n229 585
R347 B.n254 B.n253 585
R348 B.n252 B.n230 585
R349 B.n251 B.n250 585
R350 B.n248 B.n231 585
R351 B.n246 B.n245 585
R352 B.n244 B.n232 585
R353 B.n243 B.n242 585
R354 B.n240 B.n233 585
R355 B.n238 B.n237 585
R356 B.n236 B.n235 585
R357 B.n165 B.n164 585
R358 B.n484 B.n483 585
R359 B.n485 B.n484 585
R360 B.n161 B.n160 585
R361 B.n162 B.n161 585
R362 B.n493 B.n492 585
R363 B.n492 B.n491 585
R364 B.n494 B.n159 585
R365 B.n159 B.n158 585
R366 B.n496 B.n495 585
R367 B.n497 B.n496 585
R368 B.n153 B.n152 585
R369 B.n154 B.n153 585
R370 B.n506 B.n505 585
R371 B.n505 B.n504 585
R372 B.n507 B.n151 585
R373 B.n503 B.n151 585
R374 B.n509 B.n508 585
R375 B.n510 B.n509 585
R376 B.n146 B.n145 585
R377 B.n147 B.n146 585
R378 B.n518 B.n517 585
R379 B.n517 B.n516 585
R380 B.n519 B.n144 585
R381 B.n144 B.n143 585
R382 B.n521 B.n520 585
R383 B.n522 B.n521 585
R384 B.n138 B.n137 585
R385 B.n139 B.n138 585
R386 B.n530 B.n529 585
R387 B.n529 B.n528 585
R388 B.n531 B.n136 585
R389 B.n136 B.n135 585
R390 B.n533 B.n532 585
R391 B.n534 B.n533 585
R392 B.n130 B.n129 585
R393 B.n131 B.n130 585
R394 B.n543 B.n542 585
R395 B.n542 B.n541 585
R396 B.n544 B.n128 585
R397 B.n540 B.n128 585
R398 B.n546 B.n545 585
R399 B.n547 B.n546 585
R400 B.n123 B.n122 585
R401 B.n124 B.n123 585
R402 B.n556 B.n555 585
R403 B.n555 B.n554 585
R404 B.n557 B.n121 585
R405 B.n121 B.n120 585
R406 B.n559 B.n558 585
R407 B.n560 B.n559 585
R408 B.n2 B.n0 585
R409 B.n4 B.n2 585
R410 B.n3 B.n1 585
R411 B.n899 B.n3 585
R412 B.n897 B.n896 585
R413 B.n898 B.n897 585
R414 B.n895 B.n9 585
R415 B.n9 B.n8 585
R416 B.n894 B.n893 585
R417 B.n893 B.n892 585
R418 B.n11 B.n10 585
R419 B.n891 B.n11 585
R420 B.n889 B.n888 585
R421 B.n890 B.n889 585
R422 B.n887 B.n15 585
R423 B.n18 B.n15 585
R424 B.n886 B.n885 585
R425 B.n885 B.n884 585
R426 B.n17 B.n16 585
R427 B.n883 B.n17 585
R428 B.n881 B.n880 585
R429 B.n882 B.n881 585
R430 B.n879 B.n23 585
R431 B.n23 B.n22 585
R432 B.n878 B.n877 585
R433 B.n877 B.n876 585
R434 B.n25 B.n24 585
R435 B.n875 B.n25 585
R436 B.n873 B.n872 585
R437 B.n874 B.n873 585
R438 B.n871 B.n30 585
R439 B.n30 B.n29 585
R440 B.n870 B.n869 585
R441 B.n869 B.n868 585
R442 B.n32 B.n31 585
R443 B.n867 B.n32 585
R444 B.n865 B.n864 585
R445 B.n866 B.n865 585
R446 B.n863 B.n36 585
R447 B.n39 B.n36 585
R448 B.n862 B.n861 585
R449 B.n861 B.n860 585
R450 B.n38 B.n37 585
R451 B.n859 B.n38 585
R452 B.n857 B.n856 585
R453 B.n858 B.n857 585
R454 B.n855 B.n44 585
R455 B.n44 B.n43 585
R456 B.n854 B.n853 585
R457 B.n853 B.n852 585
R458 B.n46 B.n45 585
R459 B.n851 B.n46 585
R460 B.n849 B.n848 585
R461 B.n850 B.n849 585
R462 B.n902 B.n901 585
R463 B.n901 B.n900 585
R464 B.n484 B.n167 564.573
R465 B.n849 B.n51 564.573
R466 B.n486 B.n165 564.573
R467 B.n598 B.n49 564.573
R468 B.n205 B.t5 437.187
R469 B.n88 B.t8 437.187
R470 B.n198 B.t15 437.187
R471 B.n80 B.t11 437.187
R472 B.n206 B.t4 377.452
R473 B.n89 B.t9 377.452
R474 B.n199 B.t14 377.452
R475 B.n81 B.t12 377.452
R476 B.n205 B.t2 361.889
R477 B.n198 B.t13 361.889
R478 B.n80 B.t10 361.889
R479 B.n88 B.t6 361.889
R480 B.n599 B.n50 256.663
R481 B.n605 B.n50 256.663
R482 B.n607 B.n50 256.663
R483 B.n613 B.n50 256.663
R484 B.n615 B.n50 256.663
R485 B.n621 B.n50 256.663
R486 B.n623 B.n50 256.663
R487 B.n629 B.n50 256.663
R488 B.n631 B.n50 256.663
R489 B.n637 B.n50 256.663
R490 B.n639 B.n50 256.663
R491 B.n645 B.n50 256.663
R492 B.n647 B.n50 256.663
R493 B.n653 B.n50 256.663
R494 B.n655 B.n50 256.663
R495 B.n661 B.n50 256.663
R496 B.n663 B.n50 256.663
R497 B.n669 B.n50 256.663
R498 B.n671 B.n50 256.663
R499 B.n677 B.n50 256.663
R500 B.n679 B.n50 256.663
R501 B.n685 B.n50 256.663
R502 B.n687 B.n50 256.663
R503 B.n693 B.n50 256.663
R504 B.n695 B.n50 256.663
R505 B.n701 B.n50 256.663
R506 B.n703 B.n50 256.663
R507 B.n709 B.n50 256.663
R508 B.n711 B.n50 256.663
R509 B.n718 B.n50 256.663
R510 B.n720 B.n50 256.663
R511 B.n726 B.n50 256.663
R512 B.n83 B.n50 256.663
R513 B.n732 B.n50 256.663
R514 B.n738 B.n50 256.663
R515 B.n740 B.n50 256.663
R516 B.n746 B.n50 256.663
R517 B.n748 B.n50 256.663
R518 B.n754 B.n50 256.663
R519 B.n756 B.n50 256.663
R520 B.n762 B.n50 256.663
R521 B.n764 B.n50 256.663
R522 B.n770 B.n50 256.663
R523 B.n772 B.n50 256.663
R524 B.n778 B.n50 256.663
R525 B.n780 B.n50 256.663
R526 B.n786 B.n50 256.663
R527 B.n788 B.n50 256.663
R528 B.n794 B.n50 256.663
R529 B.n796 B.n50 256.663
R530 B.n802 B.n50 256.663
R531 B.n804 B.n50 256.663
R532 B.n810 B.n50 256.663
R533 B.n812 B.n50 256.663
R534 B.n818 B.n50 256.663
R535 B.n820 B.n50 256.663
R536 B.n826 B.n50 256.663
R537 B.n828 B.n50 256.663
R538 B.n834 B.n50 256.663
R539 B.n836 B.n50 256.663
R540 B.n842 B.n50 256.663
R541 B.n844 B.n50 256.663
R542 B.n479 B.n166 256.663
R543 B.n169 B.n166 256.663
R544 B.n472 B.n166 256.663
R545 B.n466 B.n166 256.663
R546 B.n464 B.n166 256.663
R547 B.n458 B.n166 256.663
R548 B.n456 B.n166 256.663
R549 B.n450 B.n166 256.663
R550 B.n448 B.n166 256.663
R551 B.n442 B.n166 256.663
R552 B.n440 B.n166 256.663
R553 B.n434 B.n166 256.663
R554 B.n432 B.n166 256.663
R555 B.n426 B.n166 256.663
R556 B.n424 B.n166 256.663
R557 B.n418 B.n166 256.663
R558 B.n416 B.n166 256.663
R559 B.n410 B.n166 256.663
R560 B.n408 B.n166 256.663
R561 B.n402 B.n166 256.663
R562 B.n400 B.n166 256.663
R563 B.n394 B.n166 256.663
R564 B.n392 B.n166 256.663
R565 B.n386 B.n166 256.663
R566 B.n384 B.n166 256.663
R567 B.n378 B.n166 256.663
R568 B.n376 B.n166 256.663
R569 B.n370 B.n166 256.663
R570 B.n368 B.n166 256.663
R571 B.n362 B.n166 256.663
R572 B.n360 B.n166 256.663
R573 B.n354 B.n166 256.663
R574 B.n352 B.n166 256.663
R575 B.n345 B.n166 256.663
R576 B.n343 B.n166 256.663
R577 B.n337 B.n166 256.663
R578 B.n335 B.n166 256.663
R579 B.n329 B.n166 256.663
R580 B.n327 B.n166 256.663
R581 B.n321 B.n166 256.663
R582 B.n319 B.n166 256.663
R583 B.n313 B.n166 256.663
R584 B.n311 B.n166 256.663
R585 B.n305 B.n166 256.663
R586 B.n303 B.n166 256.663
R587 B.n297 B.n166 256.663
R588 B.n295 B.n166 256.663
R589 B.n289 B.n166 256.663
R590 B.n287 B.n166 256.663
R591 B.n281 B.n166 256.663
R592 B.n279 B.n166 256.663
R593 B.n273 B.n166 256.663
R594 B.n271 B.n166 256.663
R595 B.n265 B.n166 256.663
R596 B.n263 B.n166 256.663
R597 B.n257 B.n166 256.663
R598 B.n255 B.n166 256.663
R599 B.n249 B.n166 256.663
R600 B.n247 B.n166 256.663
R601 B.n241 B.n166 256.663
R602 B.n239 B.n166 256.663
R603 B.n234 B.n166 256.663
R604 B.n484 B.n161 163.367
R605 B.n492 B.n161 163.367
R606 B.n492 B.n159 163.367
R607 B.n496 B.n159 163.367
R608 B.n496 B.n153 163.367
R609 B.n505 B.n153 163.367
R610 B.n505 B.n151 163.367
R611 B.n509 B.n151 163.367
R612 B.n509 B.n146 163.367
R613 B.n517 B.n146 163.367
R614 B.n517 B.n144 163.367
R615 B.n521 B.n144 163.367
R616 B.n521 B.n138 163.367
R617 B.n529 B.n138 163.367
R618 B.n529 B.n136 163.367
R619 B.n533 B.n136 163.367
R620 B.n533 B.n130 163.367
R621 B.n542 B.n130 163.367
R622 B.n542 B.n128 163.367
R623 B.n546 B.n128 163.367
R624 B.n546 B.n123 163.367
R625 B.n555 B.n123 163.367
R626 B.n555 B.n121 163.367
R627 B.n559 B.n121 163.367
R628 B.n559 B.n2 163.367
R629 B.n901 B.n2 163.367
R630 B.n901 B.n3 163.367
R631 B.n897 B.n3 163.367
R632 B.n897 B.n9 163.367
R633 B.n893 B.n9 163.367
R634 B.n893 B.n11 163.367
R635 B.n889 B.n11 163.367
R636 B.n889 B.n15 163.367
R637 B.n885 B.n15 163.367
R638 B.n885 B.n17 163.367
R639 B.n881 B.n17 163.367
R640 B.n881 B.n23 163.367
R641 B.n877 B.n23 163.367
R642 B.n877 B.n25 163.367
R643 B.n873 B.n25 163.367
R644 B.n873 B.n30 163.367
R645 B.n869 B.n30 163.367
R646 B.n869 B.n32 163.367
R647 B.n865 B.n32 163.367
R648 B.n865 B.n36 163.367
R649 B.n861 B.n36 163.367
R650 B.n861 B.n38 163.367
R651 B.n857 B.n38 163.367
R652 B.n857 B.n44 163.367
R653 B.n853 B.n44 163.367
R654 B.n853 B.n46 163.367
R655 B.n849 B.n46 163.367
R656 B.n480 B.n478 163.367
R657 B.n478 B.n477 163.367
R658 B.n474 B.n473 163.367
R659 B.n471 B.n171 163.367
R660 B.n467 B.n465 163.367
R661 B.n463 B.n173 163.367
R662 B.n459 B.n457 163.367
R663 B.n455 B.n175 163.367
R664 B.n451 B.n449 163.367
R665 B.n447 B.n177 163.367
R666 B.n443 B.n441 163.367
R667 B.n439 B.n179 163.367
R668 B.n435 B.n433 163.367
R669 B.n431 B.n181 163.367
R670 B.n427 B.n425 163.367
R671 B.n423 B.n183 163.367
R672 B.n419 B.n417 163.367
R673 B.n415 B.n185 163.367
R674 B.n411 B.n409 163.367
R675 B.n407 B.n187 163.367
R676 B.n403 B.n401 163.367
R677 B.n399 B.n189 163.367
R678 B.n395 B.n393 163.367
R679 B.n391 B.n191 163.367
R680 B.n387 B.n385 163.367
R681 B.n383 B.n193 163.367
R682 B.n379 B.n377 163.367
R683 B.n375 B.n195 163.367
R684 B.n371 B.n369 163.367
R685 B.n367 B.n197 163.367
R686 B.n363 B.n361 163.367
R687 B.n359 B.n202 163.367
R688 B.n355 B.n353 163.367
R689 B.n351 B.n204 163.367
R690 B.n346 B.n344 163.367
R691 B.n342 B.n208 163.367
R692 B.n338 B.n336 163.367
R693 B.n334 B.n210 163.367
R694 B.n330 B.n328 163.367
R695 B.n326 B.n212 163.367
R696 B.n322 B.n320 163.367
R697 B.n318 B.n214 163.367
R698 B.n314 B.n312 163.367
R699 B.n310 B.n216 163.367
R700 B.n306 B.n304 163.367
R701 B.n302 B.n218 163.367
R702 B.n298 B.n296 163.367
R703 B.n294 B.n220 163.367
R704 B.n290 B.n288 163.367
R705 B.n286 B.n222 163.367
R706 B.n282 B.n280 163.367
R707 B.n278 B.n224 163.367
R708 B.n274 B.n272 163.367
R709 B.n270 B.n226 163.367
R710 B.n266 B.n264 163.367
R711 B.n262 B.n228 163.367
R712 B.n258 B.n256 163.367
R713 B.n254 B.n230 163.367
R714 B.n250 B.n248 163.367
R715 B.n246 B.n232 163.367
R716 B.n242 B.n240 163.367
R717 B.n238 B.n235 163.367
R718 B.n486 B.n163 163.367
R719 B.n490 B.n163 163.367
R720 B.n490 B.n157 163.367
R721 B.n498 B.n157 163.367
R722 B.n498 B.n155 163.367
R723 B.n502 B.n155 163.367
R724 B.n502 B.n150 163.367
R725 B.n511 B.n150 163.367
R726 B.n511 B.n148 163.367
R727 B.n515 B.n148 163.367
R728 B.n515 B.n142 163.367
R729 B.n523 B.n142 163.367
R730 B.n523 B.n140 163.367
R731 B.n527 B.n140 163.367
R732 B.n527 B.n134 163.367
R733 B.n535 B.n134 163.367
R734 B.n535 B.n132 163.367
R735 B.n539 B.n132 163.367
R736 B.n539 B.n127 163.367
R737 B.n548 B.n127 163.367
R738 B.n548 B.n125 163.367
R739 B.n553 B.n125 163.367
R740 B.n553 B.n119 163.367
R741 B.n561 B.n119 163.367
R742 B.n562 B.n561 163.367
R743 B.n562 B.n5 163.367
R744 B.n6 B.n5 163.367
R745 B.n7 B.n6 163.367
R746 B.n567 B.n7 163.367
R747 B.n567 B.n12 163.367
R748 B.n13 B.n12 163.367
R749 B.n14 B.n13 163.367
R750 B.n572 B.n14 163.367
R751 B.n572 B.n19 163.367
R752 B.n20 B.n19 163.367
R753 B.n21 B.n20 163.367
R754 B.n577 B.n21 163.367
R755 B.n577 B.n26 163.367
R756 B.n27 B.n26 163.367
R757 B.n28 B.n27 163.367
R758 B.n582 B.n28 163.367
R759 B.n582 B.n33 163.367
R760 B.n34 B.n33 163.367
R761 B.n35 B.n34 163.367
R762 B.n587 B.n35 163.367
R763 B.n587 B.n40 163.367
R764 B.n41 B.n40 163.367
R765 B.n42 B.n41 163.367
R766 B.n592 B.n42 163.367
R767 B.n592 B.n47 163.367
R768 B.n48 B.n47 163.367
R769 B.n49 B.n48 163.367
R770 B.n845 B.n843 163.367
R771 B.n841 B.n53 163.367
R772 B.n837 B.n835 163.367
R773 B.n833 B.n55 163.367
R774 B.n829 B.n827 163.367
R775 B.n825 B.n57 163.367
R776 B.n821 B.n819 163.367
R777 B.n817 B.n59 163.367
R778 B.n813 B.n811 163.367
R779 B.n809 B.n61 163.367
R780 B.n805 B.n803 163.367
R781 B.n801 B.n63 163.367
R782 B.n797 B.n795 163.367
R783 B.n793 B.n65 163.367
R784 B.n789 B.n787 163.367
R785 B.n785 B.n67 163.367
R786 B.n781 B.n779 163.367
R787 B.n777 B.n69 163.367
R788 B.n773 B.n771 163.367
R789 B.n769 B.n71 163.367
R790 B.n765 B.n763 163.367
R791 B.n761 B.n73 163.367
R792 B.n757 B.n755 163.367
R793 B.n753 B.n75 163.367
R794 B.n749 B.n747 163.367
R795 B.n745 B.n77 163.367
R796 B.n741 B.n739 163.367
R797 B.n737 B.n79 163.367
R798 B.n733 B.n731 163.367
R799 B.n728 B.n727 163.367
R800 B.n725 B.n85 163.367
R801 B.n721 B.n719 163.367
R802 B.n717 B.n87 163.367
R803 B.n712 B.n710 163.367
R804 B.n708 B.n91 163.367
R805 B.n704 B.n702 163.367
R806 B.n700 B.n93 163.367
R807 B.n696 B.n694 163.367
R808 B.n692 B.n95 163.367
R809 B.n688 B.n686 163.367
R810 B.n684 B.n97 163.367
R811 B.n680 B.n678 163.367
R812 B.n676 B.n99 163.367
R813 B.n672 B.n670 163.367
R814 B.n668 B.n101 163.367
R815 B.n664 B.n662 163.367
R816 B.n660 B.n103 163.367
R817 B.n656 B.n654 163.367
R818 B.n652 B.n105 163.367
R819 B.n648 B.n646 163.367
R820 B.n644 B.n107 163.367
R821 B.n640 B.n638 163.367
R822 B.n636 B.n109 163.367
R823 B.n632 B.n630 163.367
R824 B.n628 B.n111 163.367
R825 B.n624 B.n622 163.367
R826 B.n620 B.n113 163.367
R827 B.n616 B.n614 163.367
R828 B.n612 B.n115 163.367
R829 B.n608 B.n606 163.367
R830 B.n604 B.n117 163.367
R831 B.n600 B.n598 163.367
R832 B.n479 B.n167 71.676
R833 B.n477 B.n169 71.676
R834 B.n473 B.n472 71.676
R835 B.n466 B.n171 71.676
R836 B.n465 B.n464 71.676
R837 B.n458 B.n173 71.676
R838 B.n457 B.n456 71.676
R839 B.n450 B.n175 71.676
R840 B.n449 B.n448 71.676
R841 B.n442 B.n177 71.676
R842 B.n441 B.n440 71.676
R843 B.n434 B.n179 71.676
R844 B.n433 B.n432 71.676
R845 B.n426 B.n181 71.676
R846 B.n425 B.n424 71.676
R847 B.n418 B.n183 71.676
R848 B.n417 B.n416 71.676
R849 B.n410 B.n185 71.676
R850 B.n409 B.n408 71.676
R851 B.n402 B.n187 71.676
R852 B.n401 B.n400 71.676
R853 B.n394 B.n189 71.676
R854 B.n393 B.n392 71.676
R855 B.n386 B.n191 71.676
R856 B.n385 B.n384 71.676
R857 B.n378 B.n193 71.676
R858 B.n377 B.n376 71.676
R859 B.n370 B.n195 71.676
R860 B.n369 B.n368 71.676
R861 B.n362 B.n197 71.676
R862 B.n361 B.n360 71.676
R863 B.n354 B.n202 71.676
R864 B.n353 B.n352 71.676
R865 B.n345 B.n204 71.676
R866 B.n344 B.n343 71.676
R867 B.n337 B.n208 71.676
R868 B.n336 B.n335 71.676
R869 B.n329 B.n210 71.676
R870 B.n328 B.n327 71.676
R871 B.n321 B.n212 71.676
R872 B.n320 B.n319 71.676
R873 B.n313 B.n214 71.676
R874 B.n312 B.n311 71.676
R875 B.n305 B.n216 71.676
R876 B.n304 B.n303 71.676
R877 B.n297 B.n218 71.676
R878 B.n296 B.n295 71.676
R879 B.n289 B.n220 71.676
R880 B.n288 B.n287 71.676
R881 B.n281 B.n222 71.676
R882 B.n280 B.n279 71.676
R883 B.n273 B.n224 71.676
R884 B.n272 B.n271 71.676
R885 B.n265 B.n226 71.676
R886 B.n264 B.n263 71.676
R887 B.n257 B.n228 71.676
R888 B.n256 B.n255 71.676
R889 B.n249 B.n230 71.676
R890 B.n248 B.n247 71.676
R891 B.n241 B.n232 71.676
R892 B.n240 B.n239 71.676
R893 B.n235 B.n234 71.676
R894 B.n844 B.n51 71.676
R895 B.n843 B.n842 71.676
R896 B.n836 B.n53 71.676
R897 B.n835 B.n834 71.676
R898 B.n828 B.n55 71.676
R899 B.n827 B.n826 71.676
R900 B.n820 B.n57 71.676
R901 B.n819 B.n818 71.676
R902 B.n812 B.n59 71.676
R903 B.n811 B.n810 71.676
R904 B.n804 B.n61 71.676
R905 B.n803 B.n802 71.676
R906 B.n796 B.n63 71.676
R907 B.n795 B.n794 71.676
R908 B.n788 B.n65 71.676
R909 B.n787 B.n786 71.676
R910 B.n780 B.n67 71.676
R911 B.n779 B.n778 71.676
R912 B.n772 B.n69 71.676
R913 B.n771 B.n770 71.676
R914 B.n764 B.n71 71.676
R915 B.n763 B.n762 71.676
R916 B.n756 B.n73 71.676
R917 B.n755 B.n754 71.676
R918 B.n748 B.n75 71.676
R919 B.n747 B.n746 71.676
R920 B.n740 B.n77 71.676
R921 B.n739 B.n738 71.676
R922 B.n732 B.n79 71.676
R923 B.n731 B.n83 71.676
R924 B.n727 B.n726 71.676
R925 B.n720 B.n85 71.676
R926 B.n719 B.n718 71.676
R927 B.n711 B.n87 71.676
R928 B.n710 B.n709 71.676
R929 B.n703 B.n91 71.676
R930 B.n702 B.n701 71.676
R931 B.n695 B.n93 71.676
R932 B.n694 B.n693 71.676
R933 B.n687 B.n95 71.676
R934 B.n686 B.n685 71.676
R935 B.n679 B.n97 71.676
R936 B.n678 B.n677 71.676
R937 B.n671 B.n99 71.676
R938 B.n670 B.n669 71.676
R939 B.n663 B.n101 71.676
R940 B.n662 B.n661 71.676
R941 B.n655 B.n103 71.676
R942 B.n654 B.n653 71.676
R943 B.n647 B.n105 71.676
R944 B.n646 B.n645 71.676
R945 B.n639 B.n107 71.676
R946 B.n638 B.n637 71.676
R947 B.n631 B.n109 71.676
R948 B.n630 B.n629 71.676
R949 B.n623 B.n111 71.676
R950 B.n622 B.n621 71.676
R951 B.n615 B.n113 71.676
R952 B.n614 B.n613 71.676
R953 B.n607 B.n115 71.676
R954 B.n606 B.n605 71.676
R955 B.n599 B.n117 71.676
R956 B.n600 B.n599 71.676
R957 B.n605 B.n604 71.676
R958 B.n608 B.n607 71.676
R959 B.n613 B.n612 71.676
R960 B.n616 B.n615 71.676
R961 B.n621 B.n620 71.676
R962 B.n624 B.n623 71.676
R963 B.n629 B.n628 71.676
R964 B.n632 B.n631 71.676
R965 B.n637 B.n636 71.676
R966 B.n640 B.n639 71.676
R967 B.n645 B.n644 71.676
R968 B.n648 B.n647 71.676
R969 B.n653 B.n652 71.676
R970 B.n656 B.n655 71.676
R971 B.n661 B.n660 71.676
R972 B.n664 B.n663 71.676
R973 B.n669 B.n668 71.676
R974 B.n672 B.n671 71.676
R975 B.n677 B.n676 71.676
R976 B.n680 B.n679 71.676
R977 B.n685 B.n684 71.676
R978 B.n688 B.n687 71.676
R979 B.n693 B.n692 71.676
R980 B.n696 B.n695 71.676
R981 B.n701 B.n700 71.676
R982 B.n704 B.n703 71.676
R983 B.n709 B.n708 71.676
R984 B.n712 B.n711 71.676
R985 B.n718 B.n717 71.676
R986 B.n721 B.n720 71.676
R987 B.n726 B.n725 71.676
R988 B.n728 B.n83 71.676
R989 B.n733 B.n732 71.676
R990 B.n738 B.n737 71.676
R991 B.n741 B.n740 71.676
R992 B.n746 B.n745 71.676
R993 B.n749 B.n748 71.676
R994 B.n754 B.n753 71.676
R995 B.n757 B.n756 71.676
R996 B.n762 B.n761 71.676
R997 B.n765 B.n764 71.676
R998 B.n770 B.n769 71.676
R999 B.n773 B.n772 71.676
R1000 B.n778 B.n777 71.676
R1001 B.n781 B.n780 71.676
R1002 B.n786 B.n785 71.676
R1003 B.n789 B.n788 71.676
R1004 B.n794 B.n793 71.676
R1005 B.n797 B.n796 71.676
R1006 B.n802 B.n801 71.676
R1007 B.n805 B.n804 71.676
R1008 B.n810 B.n809 71.676
R1009 B.n813 B.n812 71.676
R1010 B.n818 B.n817 71.676
R1011 B.n821 B.n820 71.676
R1012 B.n826 B.n825 71.676
R1013 B.n829 B.n828 71.676
R1014 B.n834 B.n833 71.676
R1015 B.n837 B.n836 71.676
R1016 B.n842 B.n841 71.676
R1017 B.n845 B.n844 71.676
R1018 B.n480 B.n479 71.676
R1019 B.n474 B.n169 71.676
R1020 B.n472 B.n471 71.676
R1021 B.n467 B.n466 71.676
R1022 B.n464 B.n463 71.676
R1023 B.n459 B.n458 71.676
R1024 B.n456 B.n455 71.676
R1025 B.n451 B.n450 71.676
R1026 B.n448 B.n447 71.676
R1027 B.n443 B.n442 71.676
R1028 B.n440 B.n439 71.676
R1029 B.n435 B.n434 71.676
R1030 B.n432 B.n431 71.676
R1031 B.n427 B.n426 71.676
R1032 B.n424 B.n423 71.676
R1033 B.n419 B.n418 71.676
R1034 B.n416 B.n415 71.676
R1035 B.n411 B.n410 71.676
R1036 B.n408 B.n407 71.676
R1037 B.n403 B.n402 71.676
R1038 B.n400 B.n399 71.676
R1039 B.n395 B.n394 71.676
R1040 B.n392 B.n391 71.676
R1041 B.n387 B.n386 71.676
R1042 B.n384 B.n383 71.676
R1043 B.n379 B.n378 71.676
R1044 B.n376 B.n375 71.676
R1045 B.n371 B.n370 71.676
R1046 B.n368 B.n367 71.676
R1047 B.n363 B.n362 71.676
R1048 B.n360 B.n359 71.676
R1049 B.n355 B.n354 71.676
R1050 B.n352 B.n351 71.676
R1051 B.n346 B.n345 71.676
R1052 B.n343 B.n342 71.676
R1053 B.n338 B.n337 71.676
R1054 B.n335 B.n334 71.676
R1055 B.n330 B.n329 71.676
R1056 B.n327 B.n326 71.676
R1057 B.n322 B.n321 71.676
R1058 B.n319 B.n318 71.676
R1059 B.n314 B.n313 71.676
R1060 B.n311 B.n310 71.676
R1061 B.n306 B.n305 71.676
R1062 B.n303 B.n302 71.676
R1063 B.n298 B.n297 71.676
R1064 B.n295 B.n294 71.676
R1065 B.n290 B.n289 71.676
R1066 B.n287 B.n286 71.676
R1067 B.n282 B.n281 71.676
R1068 B.n279 B.n278 71.676
R1069 B.n274 B.n273 71.676
R1070 B.n271 B.n270 71.676
R1071 B.n266 B.n265 71.676
R1072 B.n263 B.n262 71.676
R1073 B.n258 B.n257 71.676
R1074 B.n255 B.n254 71.676
R1075 B.n250 B.n249 71.676
R1076 B.n247 B.n246 71.676
R1077 B.n242 B.n241 71.676
R1078 B.n239 B.n238 71.676
R1079 B.n234 B.n165 71.676
R1080 B.n485 B.n166 67.0472
R1081 B.n850 B.n50 67.0472
R1082 B.n206 B.n205 59.7338
R1083 B.n199 B.n198 59.7338
R1084 B.n81 B.n80 59.7338
R1085 B.n89 B.n88 59.7338
R1086 B.n349 B.n206 59.5399
R1087 B.n200 B.n199 59.5399
R1088 B.n82 B.n81 59.5399
R1089 B.n714 B.n89 59.5399
R1090 B.n848 B.n847 36.6834
R1091 B.n597 B.n596 36.6834
R1092 B.n487 B.n164 36.6834
R1093 B.n483 B.n482 36.6834
R1094 B.n485 B.n162 32.8003
R1095 B.n491 B.n162 32.8003
R1096 B.n491 B.n158 32.8003
R1097 B.n497 B.n158 32.8003
R1098 B.n497 B.n154 32.8003
R1099 B.n504 B.n154 32.8003
R1100 B.n504 B.n503 32.8003
R1101 B.n510 B.n147 32.8003
R1102 B.n516 B.n147 32.8003
R1103 B.n516 B.n143 32.8003
R1104 B.n522 B.n143 32.8003
R1105 B.n522 B.n139 32.8003
R1106 B.n528 B.n139 32.8003
R1107 B.n528 B.n135 32.8003
R1108 B.n534 B.n135 32.8003
R1109 B.n534 B.n131 32.8003
R1110 B.n541 B.n131 32.8003
R1111 B.n541 B.n540 32.8003
R1112 B.n547 B.n124 32.8003
R1113 B.n554 B.n124 32.8003
R1114 B.n554 B.n120 32.8003
R1115 B.n560 B.n120 32.8003
R1116 B.n560 B.n4 32.8003
R1117 B.n900 B.n4 32.8003
R1118 B.n900 B.n899 32.8003
R1119 B.n899 B.n898 32.8003
R1120 B.n898 B.n8 32.8003
R1121 B.n892 B.n8 32.8003
R1122 B.n892 B.n891 32.8003
R1123 B.n891 B.n890 32.8003
R1124 B.n884 B.n18 32.8003
R1125 B.n884 B.n883 32.8003
R1126 B.n883 B.n882 32.8003
R1127 B.n882 B.n22 32.8003
R1128 B.n876 B.n22 32.8003
R1129 B.n876 B.n875 32.8003
R1130 B.n875 B.n874 32.8003
R1131 B.n874 B.n29 32.8003
R1132 B.n868 B.n29 32.8003
R1133 B.n868 B.n867 32.8003
R1134 B.n867 B.n866 32.8003
R1135 B.n860 B.n39 32.8003
R1136 B.n860 B.n859 32.8003
R1137 B.n859 B.n858 32.8003
R1138 B.n858 B.n43 32.8003
R1139 B.n852 B.n43 32.8003
R1140 B.n852 B.n851 32.8003
R1141 B.n851 B.n850 32.8003
R1142 B.n540 B.t1 28.4592
R1143 B.n18 B.t0 28.4592
R1144 B.n503 B.t3 19.7769
R1145 B.n39 B.t7 19.7769
R1146 B B.n902 18.0485
R1147 B.n510 B.t3 13.024
R1148 B.n866 B.t7 13.024
R1149 B.n847 B.n846 10.6151
R1150 B.n846 B.n52 10.6151
R1151 B.n840 B.n52 10.6151
R1152 B.n840 B.n839 10.6151
R1153 B.n839 B.n838 10.6151
R1154 B.n838 B.n54 10.6151
R1155 B.n832 B.n54 10.6151
R1156 B.n832 B.n831 10.6151
R1157 B.n831 B.n830 10.6151
R1158 B.n830 B.n56 10.6151
R1159 B.n824 B.n56 10.6151
R1160 B.n824 B.n823 10.6151
R1161 B.n823 B.n822 10.6151
R1162 B.n822 B.n58 10.6151
R1163 B.n816 B.n58 10.6151
R1164 B.n816 B.n815 10.6151
R1165 B.n815 B.n814 10.6151
R1166 B.n814 B.n60 10.6151
R1167 B.n808 B.n60 10.6151
R1168 B.n808 B.n807 10.6151
R1169 B.n807 B.n806 10.6151
R1170 B.n806 B.n62 10.6151
R1171 B.n800 B.n62 10.6151
R1172 B.n800 B.n799 10.6151
R1173 B.n799 B.n798 10.6151
R1174 B.n798 B.n64 10.6151
R1175 B.n792 B.n64 10.6151
R1176 B.n792 B.n791 10.6151
R1177 B.n791 B.n790 10.6151
R1178 B.n790 B.n66 10.6151
R1179 B.n784 B.n66 10.6151
R1180 B.n784 B.n783 10.6151
R1181 B.n783 B.n782 10.6151
R1182 B.n782 B.n68 10.6151
R1183 B.n776 B.n68 10.6151
R1184 B.n776 B.n775 10.6151
R1185 B.n775 B.n774 10.6151
R1186 B.n774 B.n70 10.6151
R1187 B.n768 B.n70 10.6151
R1188 B.n768 B.n767 10.6151
R1189 B.n767 B.n766 10.6151
R1190 B.n766 B.n72 10.6151
R1191 B.n760 B.n72 10.6151
R1192 B.n760 B.n759 10.6151
R1193 B.n759 B.n758 10.6151
R1194 B.n758 B.n74 10.6151
R1195 B.n752 B.n74 10.6151
R1196 B.n752 B.n751 10.6151
R1197 B.n751 B.n750 10.6151
R1198 B.n750 B.n76 10.6151
R1199 B.n744 B.n76 10.6151
R1200 B.n744 B.n743 10.6151
R1201 B.n743 B.n742 10.6151
R1202 B.n742 B.n78 10.6151
R1203 B.n736 B.n78 10.6151
R1204 B.n736 B.n735 10.6151
R1205 B.n735 B.n734 10.6151
R1206 B.n730 B.n729 10.6151
R1207 B.n729 B.n84 10.6151
R1208 B.n724 B.n84 10.6151
R1209 B.n724 B.n723 10.6151
R1210 B.n723 B.n722 10.6151
R1211 B.n722 B.n86 10.6151
R1212 B.n716 B.n86 10.6151
R1213 B.n716 B.n715 10.6151
R1214 B.n713 B.n90 10.6151
R1215 B.n707 B.n90 10.6151
R1216 B.n707 B.n706 10.6151
R1217 B.n706 B.n705 10.6151
R1218 B.n705 B.n92 10.6151
R1219 B.n699 B.n92 10.6151
R1220 B.n699 B.n698 10.6151
R1221 B.n698 B.n697 10.6151
R1222 B.n697 B.n94 10.6151
R1223 B.n691 B.n94 10.6151
R1224 B.n691 B.n690 10.6151
R1225 B.n690 B.n689 10.6151
R1226 B.n689 B.n96 10.6151
R1227 B.n683 B.n96 10.6151
R1228 B.n683 B.n682 10.6151
R1229 B.n682 B.n681 10.6151
R1230 B.n681 B.n98 10.6151
R1231 B.n675 B.n98 10.6151
R1232 B.n675 B.n674 10.6151
R1233 B.n674 B.n673 10.6151
R1234 B.n673 B.n100 10.6151
R1235 B.n667 B.n100 10.6151
R1236 B.n667 B.n666 10.6151
R1237 B.n666 B.n665 10.6151
R1238 B.n665 B.n102 10.6151
R1239 B.n659 B.n102 10.6151
R1240 B.n659 B.n658 10.6151
R1241 B.n658 B.n657 10.6151
R1242 B.n657 B.n104 10.6151
R1243 B.n651 B.n104 10.6151
R1244 B.n651 B.n650 10.6151
R1245 B.n650 B.n649 10.6151
R1246 B.n649 B.n106 10.6151
R1247 B.n643 B.n106 10.6151
R1248 B.n643 B.n642 10.6151
R1249 B.n642 B.n641 10.6151
R1250 B.n641 B.n108 10.6151
R1251 B.n635 B.n108 10.6151
R1252 B.n635 B.n634 10.6151
R1253 B.n634 B.n633 10.6151
R1254 B.n633 B.n110 10.6151
R1255 B.n627 B.n110 10.6151
R1256 B.n627 B.n626 10.6151
R1257 B.n626 B.n625 10.6151
R1258 B.n625 B.n112 10.6151
R1259 B.n619 B.n112 10.6151
R1260 B.n619 B.n618 10.6151
R1261 B.n618 B.n617 10.6151
R1262 B.n617 B.n114 10.6151
R1263 B.n611 B.n114 10.6151
R1264 B.n611 B.n610 10.6151
R1265 B.n610 B.n609 10.6151
R1266 B.n609 B.n116 10.6151
R1267 B.n603 B.n116 10.6151
R1268 B.n603 B.n602 10.6151
R1269 B.n602 B.n601 10.6151
R1270 B.n601 B.n597 10.6151
R1271 B.n488 B.n487 10.6151
R1272 B.n489 B.n488 10.6151
R1273 B.n489 B.n156 10.6151
R1274 B.n499 B.n156 10.6151
R1275 B.n500 B.n499 10.6151
R1276 B.n501 B.n500 10.6151
R1277 B.n501 B.n149 10.6151
R1278 B.n512 B.n149 10.6151
R1279 B.n513 B.n512 10.6151
R1280 B.n514 B.n513 10.6151
R1281 B.n514 B.n141 10.6151
R1282 B.n524 B.n141 10.6151
R1283 B.n525 B.n524 10.6151
R1284 B.n526 B.n525 10.6151
R1285 B.n526 B.n133 10.6151
R1286 B.n536 B.n133 10.6151
R1287 B.n537 B.n536 10.6151
R1288 B.n538 B.n537 10.6151
R1289 B.n538 B.n126 10.6151
R1290 B.n549 B.n126 10.6151
R1291 B.n550 B.n549 10.6151
R1292 B.n552 B.n550 10.6151
R1293 B.n552 B.n551 10.6151
R1294 B.n551 B.n118 10.6151
R1295 B.n563 B.n118 10.6151
R1296 B.n564 B.n563 10.6151
R1297 B.n565 B.n564 10.6151
R1298 B.n566 B.n565 10.6151
R1299 B.n568 B.n566 10.6151
R1300 B.n569 B.n568 10.6151
R1301 B.n570 B.n569 10.6151
R1302 B.n571 B.n570 10.6151
R1303 B.n573 B.n571 10.6151
R1304 B.n574 B.n573 10.6151
R1305 B.n575 B.n574 10.6151
R1306 B.n576 B.n575 10.6151
R1307 B.n578 B.n576 10.6151
R1308 B.n579 B.n578 10.6151
R1309 B.n580 B.n579 10.6151
R1310 B.n581 B.n580 10.6151
R1311 B.n583 B.n581 10.6151
R1312 B.n584 B.n583 10.6151
R1313 B.n585 B.n584 10.6151
R1314 B.n586 B.n585 10.6151
R1315 B.n588 B.n586 10.6151
R1316 B.n589 B.n588 10.6151
R1317 B.n590 B.n589 10.6151
R1318 B.n591 B.n590 10.6151
R1319 B.n593 B.n591 10.6151
R1320 B.n594 B.n593 10.6151
R1321 B.n595 B.n594 10.6151
R1322 B.n596 B.n595 10.6151
R1323 B.n482 B.n481 10.6151
R1324 B.n481 B.n168 10.6151
R1325 B.n476 B.n168 10.6151
R1326 B.n476 B.n475 10.6151
R1327 B.n475 B.n170 10.6151
R1328 B.n470 B.n170 10.6151
R1329 B.n470 B.n469 10.6151
R1330 B.n469 B.n468 10.6151
R1331 B.n468 B.n172 10.6151
R1332 B.n462 B.n172 10.6151
R1333 B.n462 B.n461 10.6151
R1334 B.n461 B.n460 10.6151
R1335 B.n460 B.n174 10.6151
R1336 B.n454 B.n174 10.6151
R1337 B.n454 B.n453 10.6151
R1338 B.n453 B.n452 10.6151
R1339 B.n452 B.n176 10.6151
R1340 B.n446 B.n176 10.6151
R1341 B.n446 B.n445 10.6151
R1342 B.n445 B.n444 10.6151
R1343 B.n444 B.n178 10.6151
R1344 B.n438 B.n178 10.6151
R1345 B.n438 B.n437 10.6151
R1346 B.n437 B.n436 10.6151
R1347 B.n436 B.n180 10.6151
R1348 B.n430 B.n180 10.6151
R1349 B.n430 B.n429 10.6151
R1350 B.n429 B.n428 10.6151
R1351 B.n428 B.n182 10.6151
R1352 B.n422 B.n182 10.6151
R1353 B.n422 B.n421 10.6151
R1354 B.n421 B.n420 10.6151
R1355 B.n420 B.n184 10.6151
R1356 B.n414 B.n184 10.6151
R1357 B.n414 B.n413 10.6151
R1358 B.n413 B.n412 10.6151
R1359 B.n412 B.n186 10.6151
R1360 B.n406 B.n186 10.6151
R1361 B.n406 B.n405 10.6151
R1362 B.n405 B.n404 10.6151
R1363 B.n404 B.n188 10.6151
R1364 B.n398 B.n188 10.6151
R1365 B.n398 B.n397 10.6151
R1366 B.n397 B.n396 10.6151
R1367 B.n396 B.n190 10.6151
R1368 B.n390 B.n190 10.6151
R1369 B.n390 B.n389 10.6151
R1370 B.n389 B.n388 10.6151
R1371 B.n388 B.n192 10.6151
R1372 B.n382 B.n192 10.6151
R1373 B.n382 B.n381 10.6151
R1374 B.n381 B.n380 10.6151
R1375 B.n380 B.n194 10.6151
R1376 B.n374 B.n194 10.6151
R1377 B.n374 B.n373 10.6151
R1378 B.n373 B.n372 10.6151
R1379 B.n372 B.n196 10.6151
R1380 B.n366 B.n365 10.6151
R1381 B.n365 B.n364 10.6151
R1382 B.n364 B.n201 10.6151
R1383 B.n358 B.n201 10.6151
R1384 B.n358 B.n357 10.6151
R1385 B.n357 B.n356 10.6151
R1386 B.n356 B.n203 10.6151
R1387 B.n350 B.n203 10.6151
R1388 B.n348 B.n347 10.6151
R1389 B.n347 B.n207 10.6151
R1390 B.n341 B.n207 10.6151
R1391 B.n341 B.n340 10.6151
R1392 B.n340 B.n339 10.6151
R1393 B.n339 B.n209 10.6151
R1394 B.n333 B.n209 10.6151
R1395 B.n333 B.n332 10.6151
R1396 B.n332 B.n331 10.6151
R1397 B.n331 B.n211 10.6151
R1398 B.n325 B.n211 10.6151
R1399 B.n325 B.n324 10.6151
R1400 B.n324 B.n323 10.6151
R1401 B.n323 B.n213 10.6151
R1402 B.n317 B.n213 10.6151
R1403 B.n317 B.n316 10.6151
R1404 B.n316 B.n315 10.6151
R1405 B.n315 B.n215 10.6151
R1406 B.n309 B.n215 10.6151
R1407 B.n309 B.n308 10.6151
R1408 B.n308 B.n307 10.6151
R1409 B.n307 B.n217 10.6151
R1410 B.n301 B.n217 10.6151
R1411 B.n301 B.n300 10.6151
R1412 B.n300 B.n299 10.6151
R1413 B.n299 B.n219 10.6151
R1414 B.n293 B.n219 10.6151
R1415 B.n293 B.n292 10.6151
R1416 B.n292 B.n291 10.6151
R1417 B.n291 B.n221 10.6151
R1418 B.n285 B.n221 10.6151
R1419 B.n285 B.n284 10.6151
R1420 B.n284 B.n283 10.6151
R1421 B.n283 B.n223 10.6151
R1422 B.n277 B.n223 10.6151
R1423 B.n277 B.n276 10.6151
R1424 B.n276 B.n275 10.6151
R1425 B.n275 B.n225 10.6151
R1426 B.n269 B.n225 10.6151
R1427 B.n269 B.n268 10.6151
R1428 B.n268 B.n267 10.6151
R1429 B.n267 B.n227 10.6151
R1430 B.n261 B.n227 10.6151
R1431 B.n261 B.n260 10.6151
R1432 B.n260 B.n259 10.6151
R1433 B.n259 B.n229 10.6151
R1434 B.n253 B.n229 10.6151
R1435 B.n253 B.n252 10.6151
R1436 B.n252 B.n251 10.6151
R1437 B.n251 B.n231 10.6151
R1438 B.n245 B.n231 10.6151
R1439 B.n245 B.n244 10.6151
R1440 B.n244 B.n243 10.6151
R1441 B.n243 B.n233 10.6151
R1442 B.n237 B.n233 10.6151
R1443 B.n237 B.n236 10.6151
R1444 B.n236 B.n164 10.6151
R1445 B.n483 B.n160 10.6151
R1446 B.n493 B.n160 10.6151
R1447 B.n494 B.n493 10.6151
R1448 B.n495 B.n494 10.6151
R1449 B.n495 B.n152 10.6151
R1450 B.n506 B.n152 10.6151
R1451 B.n507 B.n506 10.6151
R1452 B.n508 B.n507 10.6151
R1453 B.n508 B.n145 10.6151
R1454 B.n518 B.n145 10.6151
R1455 B.n519 B.n518 10.6151
R1456 B.n520 B.n519 10.6151
R1457 B.n520 B.n137 10.6151
R1458 B.n530 B.n137 10.6151
R1459 B.n531 B.n530 10.6151
R1460 B.n532 B.n531 10.6151
R1461 B.n532 B.n129 10.6151
R1462 B.n543 B.n129 10.6151
R1463 B.n544 B.n543 10.6151
R1464 B.n545 B.n544 10.6151
R1465 B.n545 B.n122 10.6151
R1466 B.n556 B.n122 10.6151
R1467 B.n557 B.n556 10.6151
R1468 B.n558 B.n557 10.6151
R1469 B.n558 B.n0 10.6151
R1470 B.n896 B.n1 10.6151
R1471 B.n896 B.n895 10.6151
R1472 B.n895 B.n894 10.6151
R1473 B.n894 B.n10 10.6151
R1474 B.n888 B.n10 10.6151
R1475 B.n888 B.n887 10.6151
R1476 B.n887 B.n886 10.6151
R1477 B.n886 B.n16 10.6151
R1478 B.n880 B.n16 10.6151
R1479 B.n880 B.n879 10.6151
R1480 B.n879 B.n878 10.6151
R1481 B.n878 B.n24 10.6151
R1482 B.n872 B.n24 10.6151
R1483 B.n872 B.n871 10.6151
R1484 B.n871 B.n870 10.6151
R1485 B.n870 B.n31 10.6151
R1486 B.n864 B.n31 10.6151
R1487 B.n864 B.n863 10.6151
R1488 B.n863 B.n862 10.6151
R1489 B.n862 B.n37 10.6151
R1490 B.n856 B.n37 10.6151
R1491 B.n856 B.n855 10.6151
R1492 B.n855 B.n854 10.6151
R1493 B.n854 B.n45 10.6151
R1494 B.n848 B.n45 10.6151
R1495 B.n730 B.n82 6.5566
R1496 B.n715 B.n714 6.5566
R1497 B.n366 B.n200 6.5566
R1498 B.n350 B.n349 6.5566
R1499 B.n547 B.t1 4.34165
R1500 B.n890 B.t0 4.34165
R1501 B.n734 B.n82 4.05904
R1502 B.n714 B.n713 4.05904
R1503 B.n200 B.n196 4.05904
R1504 B.n349 B.n348 4.05904
R1505 B.n902 B.n0 2.81026
R1506 B.n902 B.n1 2.81026
R1507 VN VN.t1 243.969
R1508 VN VN.t0 195.155
R1509 VTAIL.n386 VTAIL.n294 289.615
R1510 VTAIL.n92 VTAIL.n0 289.615
R1511 VTAIL.n288 VTAIL.n196 289.615
R1512 VTAIL.n190 VTAIL.n98 289.615
R1513 VTAIL.n327 VTAIL.n326 185
R1514 VTAIL.n329 VTAIL.n328 185
R1515 VTAIL.n322 VTAIL.n321 185
R1516 VTAIL.n335 VTAIL.n334 185
R1517 VTAIL.n337 VTAIL.n336 185
R1518 VTAIL.n318 VTAIL.n317 185
R1519 VTAIL.n343 VTAIL.n342 185
R1520 VTAIL.n345 VTAIL.n344 185
R1521 VTAIL.n314 VTAIL.n313 185
R1522 VTAIL.n351 VTAIL.n350 185
R1523 VTAIL.n353 VTAIL.n352 185
R1524 VTAIL.n310 VTAIL.n309 185
R1525 VTAIL.n359 VTAIL.n358 185
R1526 VTAIL.n361 VTAIL.n360 185
R1527 VTAIL.n306 VTAIL.n305 185
R1528 VTAIL.n368 VTAIL.n367 185
R1529 VTAIL.n369 VTAIL.n304 185
R1530 VTAIL.n371 VTAIL.n370 185
R1531 VTAIL.n302 VTAIL.n301 185
R1532 VTAIL.n377 VTAIL.n376 185
R1533 VTAIL.n379 VTAIL.n378 185
R1534 VTAIL.n298 VTAIL.n297 185
R1535 VTAIL.n385 VTAIL.n384 185
R1536 VTAIL.n387 VTAIL.n386 185
R1537 VTAIL.n33 VTAIL.n32 185
R1538 VTAIL.n35 VTAIL.n34 185
R1539 VTAIL.n28 VTAIL.n27 185
R1540 VTAIL.n41 VTAIL.n40 185
R1541 VTAIL.n43 VTAIL.n42 185
R1542 VTAIL.n24 VTAIL.n23 185
R1543 VTAIL.n49 VTAIL.n48 185
R1544 VTAIL.n51 VTAIL.n50 185
R1545 VTAIL.n20 VTAIL.n19 185
R1546 VTAIL.n57 VTAIL.n56 185
R1547 VTAIL.n59 VTAIL.n58 185
R1548 VTAIL.n16 VTAIL.n15 185
R1549 VTAIL.n65 VTAIL.n64 185
R1550 VTAIL.n67 VTAIL.n66 185
R1551 VTAIL.n12 VTAIL.n11 185
R1552 VTAIL.n74 VTAIL.n73 185
R1553 VTAIL.n75 VTAIL.n10 185
R1554 VTAIL.n77 VTAIL.n76 185
R1555 VTAIL.n8 VTAIL.n7 185
R1556 VTAIL.n83 VTAIL.n82 185
R1557 VTAIL.n85 VTAIL.n84 185
R1558 VTAIL.n4 VTAIL.n3 185
R1559 VTAIL.n91 VTAIL.n90 185
R1560 VTAIL.n93 VTAIL.n92 185
R1561 VTAIL.n289 VTAIL.n288 185
R1562 VTAIL.n287 VTAIL.n286 185
R1563 VTAIL.n200 VTAIL.n199 185
R1564 VTAIL.n281 VTAIL.n280 185
R1565 VTAIL.n279 VTAIL.n278 185
R1566 VTAIL.n204 VTAIL.n203 185
R1567 VTAIL.n208 VTAIL.n206 185
R1568 VTAIL.n273 VTAIL.n272 185
R1569 VTAIL.n271 VTAIL.n270 185
R1570 VTAIL.n210 VTAIL.n209 185
R1571 VTAIL.n265 VTAIL.n264 185
R1572 VTAIL.n263 VTAIL.n262 185
R1573 VTAIL.n214 VTAIL.n213 185
R1574 VTAIL.n257 VTAIL.n256 185
R1575 VTAIL.n255 VTAIL.n254 185
R1576 VTAIL.n218 VTAIL.n217 185
R1577 VTAIL.n249 VTAIL.n248 185
R1578 VTAIL.n247 VTAIL.n246 185
R1579 VTAIL.n222 VTAIL.n221 185
R1580 VTAIL.n241 VTAIL.n240 185
R1581 VTAIL.n239 VTAIL.n238 185
R1582 VTAIL.n226 VTAIL.n225 185
R1583 VTAIL.n233 VTAIL.n232 185
R1584 VTAIL.n231 VTAIL.n230 185
R1585 VTAIL.n191 VTAIL.n190 185
R1586 VTAIL.n189 VTAIL.n188 185
R1587 VTAIL.n102 VTAIL.n101 185
R1588 VTAIL.n183 VTAIL.n182 185
R1589 VTAIL.n181 VTAIL.n180 185
R1590 VTAIL.n106 VTAIL.n105 185
R1591 VTAIL.n110 VTAIL.n108 185
R1592 VTAIL.n175 VTAIL.n174 185
R1593 VTAIL.n173 VTAIL.n172 185
R1594 VTAIL.n112 VTAIL.n111 185
R1595 VTAIL.n167 VTAIL.n166 185
R1596 VTAIL.n165 VTAIL.n164 185
R1597 VTAIL.n116 VTAIL.n115 185
R1598 VTAIL.n159 VTAIL.n158 185
R1599 VTAIL.n157 VTAIL.n156 185
R1600 VTAIL.n120 VTAIL.n119 185
R1601 VTAIL.n151 VTAIL.n150 185
R1602 VTAIL.n149 VTAIL.n148 185
R1603 VTAIL.n124 VTAIL.n123 185
R1604 VTAIL.n143 VTAIL.n142 185
R1605 VTAIL.n141 VTAIL.n140 185
R1606 VTAIL.n128 VTAIL.n127 185
R1607 VTAIL.n135 VTAIL.n134 185
R1608 VTAIL.n133 VTAIL.n132 185
R1609 VTAIL.n325 VTAIL.t0 147.659
R1610 VTAIL.n31 VTAIL.t3 147.659
R1611 VTAIL.n229 VTAIL.t2 147.659
R1612 VTAIL.n131 VTAIL.t1 147.659
R1613 VTAIL.n328 VTAIL.n327 104.615
R1614 VTAIL.n328 VTAIL.n321 104.615
R1615 VTAIL.n335 VTAIL.n321 104.615
R1616 VTAIL.n336 VTAIL.n335 104.615
R1617 VTAIL.n336 VTAIL.n317 104.615
R1618 VTAIL.n343 VTAIL.n317 104.615
R1619 VTAIL.n344 VTAIL.n343 104.615
R1620 VTAIL.n344 VTAIL.n313 104.615
R1621 VTAIL.n351 VTAIL.n313 104.615
R1622 VTAIL.n352 VTAIL.n351 104.615
R1623 VTAIL.n352 VTAIL.n309 104.615
R1624 VTAIL.n359 VTAIL.n309 104.615
R1625 VTAIL.n360 VTAIL.n359 104.615
R1626 VTAIL.n360 VTAIL.n305 104.615
R1627 VTAIL.n368 VTAIL.n305 104.615
R1628 VTAIL.n369 VTAIL.n368 104.615
R1629 VTAIL.n370 VTAIL.n369 104.615
R1630 VTAIL.n370 VTAIL.n301 104.615
R1631 VTAIL.n377 VTAIL.n301 104.615
R1632 VTAIL.n378 VTAIL.n377 104.615
R1633 VTAIL.n378 VTAIL.n297 104.615
R1634 VTAIL.n385 VTAIL.n297 104.615
R1635 VTAIL.n386 VTAIL.n385 104.615
R1636 VTAIL.n34 VTAIL.n33 104.615
R1637 VTAIL.n34 VTAIL.n27 104.615
R1638 VTAIL.n41 VTAIL.n27 104.615
R1639 VTAIL.n42 VTAIL.n41 104.615
R1640 VTAIL.n42 VTAIL.n23 104.615
R1641 VTAIL.n49 VTAIL.n23 104.615
R1642 VTAIL.n50 VTAIL.n49 104.615
R1643 VTAIL.n50 VTAIL.n19 104.615
R1644 VTAIL.n57 VTAIL.n19 104.615
R1645 VTAIL.n58 VTAIL.n57 104.615
R1646 VTAIL.n58 VTAIL.n15 104.615
R1647 VTAIL.n65 VTAIL.n15 104.615
R1648 VTAIL.n66 VTAIL.n65 104.615
R1649 VTAIL.n66 VTAIL.n11 104.615
R1650 VTAIL.n74 VTAIL.n11 104.615
R1651 VTAIL.n75 VTAIL.n74 104.615
R1652 VTAIL.n76 VTAIL.n75 104.615
R1653 VTAIL.n76 VTAIL.n7 104.615
R1654 VTAIL.n83 VTAIL.n7 104.615
R1655 VTAIL.n84 VTAIL.n83 104.615
R1656 VTAIL.n84 VTAIL.n3 104.615
R1657 VTAIL.n91 VTAIL.n3 104.615
R1658 VTAIL.n92 VTAIL.n91 104.615
R1659 VTAIL.n288 VTAIL.n287 104.615
R1660 VTAIL.n287 VTAIL.n199 104.615
R1661 VTAIL.n280 VTAIL.n199 104.615
R1662 VTAIL.n280 VTAIL.n279 104.615
R1663 VTAIL.n279 VTAIL.n203 104.615
R1664 VTAIL.n208 VTAIL.n203 104.615
R1665 VTAIL.n272 VTAIL.n208 104.615
R1666 VTAIL.n272 VTAIL.n271 104.615
R1667 VTAIL.n271 VTAIL.n209 104.615
R1668 VTAIL.n264 VTAIL.n209 104.615
R1669 VTAIL.n264 VTAIL.n263 104.615
R1670 VTAIL.n263 VTAIL.n213 104.615
R1671 VTAIL.n256 VTAIL.n213 104.615
R1672 VTAIL.n256 VTAIL.n255 104.615
R1673 VTAIL.n255 VTAIL.n217 104.615
R1674 VTAIL.n248 VTAIL.n217 104.615
R1675 VTAIL.n248 VTAIL.n247 104.615
R1676 VTAIL.n247 VTAIL.n221 104.615
R1677 VTAIL.n240 VTAIL.n221 104.615
R1678 VTAIL.n240 VTAIL.n239 104.615
R1679 VTAIL.n239 VTAIL.n225 104.615
R1680 VTAIL.n232 VTAIL.n225 104.615
R1681 VTAIL.n232 VTAIL.n231 104.615
R1682 VTAIL.n190 VTAIL.n189 104.615
R1683 VTAIL.n189 VTAIL.n101 104.615
R1684 VTAIL.n182 VTAIL.n101 104.615
R1685 VTAIL.n182 VTAIL.n181 104.615
R1686 VTAIL.n181 VTAIL.n105 104.615
R1687 VTAIL.n110 VTAIL.n105 104.615
R1688 VTAIL.n174 VTAIL.n110 104.615
R1689 VTAIL.n174 VTAIL.n173 104.615
R1690 VTAIL.n173 VTAIL.n111 104.615
R1691 VTAIL.n166 VTAIL.n111 104.615
R1692 VTAIL.n166 VTAIL.n165 104.615
R1693 VTAIL.n165 VTAIL.n115 104.615
R1694 VTAIL.n158 VTAIL.n115 104.615
R1695 VTAIL.n158 VTAIL.n157 104.615
R1696 VTAIL.n157 VTAIL.n119 104.615
R1697 VTAIL.n150 VTAIL.n119 104.615
R1698 VTAIL.n150 VTAIL.n149 104.615
R1699 VTAIL.n149 VTAIL.n123 104.615
R1700 VTAIL.n142 VTAIL.n123 104.615
R1701 VTAIL.n142 VTAIL.n141 104.615
R1702 VTAIL.n141 VTAIL.n127 104.615
R1703 VTAIL.n134 VTAIL.n127 104.615
R1704 VTAIL.n134 VTAIL.n133 104.615
R1705 VTAIL.n327 VTAIL.t0 52.3082
R1706 VTAIL.n33 VTAIL.t3 52.3082
R1707 VTAIL.n231 VTAIL.t2 52.3082
R1708 VTAIL.n133 VTAIL.t1 52.3082
R1709 VTAIL.n195 VTAIL.n97 32.7893
R1710 VTAIL.n391 VTAIL.n390 32.3793
R1711 VTAIL.n97 VTAIL.n96 32.3793
R1712 VTAIL.n293 VTAIL.n292 32.3793
R1713 VTAIL.n195 VTAIL.n194 32.3793
R1714 VTAIL.n391 VTAIL.n293 30.1341
R1715 VTAIL.n326 VTAIL.n325 15.6677
R1716 VTAIL.n32 VTAIL.n31 15.6677
R1717 VTAIL.n230 VTAIL.n229 15.6677
R1718 VTAIL.n132 VTAIL.n131 15.6677
R1719 VTAIL.n371 VTAIL.n302 13.1884
R1720 VTAIL.n77 VTAIL.n8 13.1884
R1721 VTAIL.n206 VTAIL.n204 13.1884
R1722 VTAIL.n108 VTAIL.n106 13.1884
R1723 VTAIL.n329 VTAIL.n324 12.8005
R1724 VTAIL.n372 VTAIL.n304 12.8005
R1725 VTAIL.n376 VTAIL.n375 12.8005
R1726 VTAIL.n35 VTAIL.n30 12.8005
R1727 VTAIL.n78 VTAIL.n10 12.8005
R1728 VTAIL.n82 VTAIL.n81 12.8005
R1729 VTAIL.n278 VTAIL.n277 12.8005
R1730 VTAIL.n274 VTAIL.n273 12.8005
R1731 VTAIL.n233 VTAIL.n228 12.8005
R1732 VTAIL.n180 VTAIL.n179 12.8005
R1733 VTAIL.n176 VTAIL.n175 12.8005
R1734 VTAIL.n135 VTAIL.n130 12.8005
R1735 VTAIL.n330 VTAIL.n322 12.0247
R1736 VTAIL.n367 VTAIL.n366 12.0247
R1737 VTAIL.n379 VTAIL.n300 12.0247
R1738 VTAIL.n36 VTAIL.n28 12.0247
R1739 VTAIL.n73 VTAIL.n72 12.0247
R1740 VTAIL.n85 VTAIL.n6 12.0247
R1741 VTAIL.n281 VTAIL.n202 12.0247
R1742 VTAIL.n270 VTAIL.n207 12.0247
R1743 VTAIL.n234 VTAIL.n226 12.0247
R1744 VTAIL.n183 VTAIL.n104 12.0247
R1745 VTAIL.n172 VTAIL.n109 12.0247
R1746 VTAIL.n136 VTAIL.n128 12.0247
R1747 VTAIL.n334 VTAIL.n333 11.249
R1748 VTAIL.n365 VTAIL.n306 11.249
R1749 VTAIL.n380 VTAIL.n298 11.249
R1750 VTAIL.n40 VTAIL.n39 11.249
R1751 VTAIL.n71 VTAIL.n12 11.249
R1752 VTAIL.n86 VTAIL.n4 11.249
R1753 VTAIL.n282 VTAIL.n200 11.249
R1754 VTAIL.n269 VTAIL.n210 11.249
R1755 VTAIL.n238 VTAIL.n237 11.249
R1756 VTAIL.n184 VTAIL.n102 11.249
R1757 VTAIL.n171 VTAIL.n112 11.249
R1758 VTAIL.n140 VTAIL.n139 11.249
R1759 VTAIL.n337 VTAIL.n320 10.4732
R1760 VTAIL.n362 VTAIL.n361 10.4732
R1761 VTAIL.n384 VTAIL.n383 10.4732
R1762 VTAIL.n43 VTAIL.n26 10.4732
R1763 VTAIL.n68 VTAIL.n67 10.4732
R1764 VTAIL.n90 VTAIL.n89 10.4732
R1765 VTAIL.n286 VTAIL.n285 10.4732
R1766 VTAIL.n266 VTAIL.n265 10.4732
R1767 VTAIL.n241 VTAIL.n224 10.4732
R1768 VTAIL.n188 VTAIL.n187 10.4732
R1769 VTAIL.n168 VTAIL.n167 10.4732
R1770 VTAIL.n143 VTAIL.n126 10.4732
R1771 VTAIL.n338 VTAIL.n318 9.69747
R1772 VTAIL.n358 VTAIL.n308 9.69747
R1773 VTAIL.n387 VTAIL.n296 9.69747
R1774 VTAIL.n44 VTAIL.n24 9.69747
R1775 VTAIL.n64 VTAIL.n14 9.69747
R1776 VTAIL.n93 VTAIL.n2 9.69747
R1777 VTAIL.n289 VTAIL.n198 9.69747
R1778 VTAIL.n262 VTAIL.n212 9.69747
R1779 VTAIL.n242 VTAIL.n222 9.69747
R1780 VTAIL.n191 VTAIL.n100 9.69747
R1781 VTAIL.n164 VTAIL.n114 9.69747
R1782 VTAIL.n144 VTAIL.n124 9.69747
R1783 VTAIL.n390 VTAIL.n389 9.45567
R1784 VTAIL.n96 VTAIL.n95 9.45567
R1785 VTAIL.n292 VTAIL.n291 9.45567
R1786 VTAIL.n194 VTAIL.n193 9.45567
R1787 VTAIL.n389 VTAIL.n388 9.3005
R1788 VTAIL.n296 VTAIL.n295 9.3005
R1789 VTAIL.n383 VTAIL.n382 9.3005
R1790 VTAIL.n381 VTAIL.n380 9.3005
R1791 VTAIL.n300 VTAIL.n299 9.3005
R1792 VTAIL.n375 VTAIL.n374 9.3005
R1793 VTAIL.n347 VTAIL.n346 9.3005
R1794 VTAIL.n316 VTAIL.n315 9.3005
R1795 VTAIL.n341 VTAIL.n340 9.3005
R1796 VTAIL.n339 VTAIL.n338 9.3005
R1797 VTAIL.n320 VTAIL.n319 9.3005
R1798 VTAIL.n333 VTAIL.n332 9.3005
R1799 VTAIL.n331 VTAIL.n330 9.3005
R1800 VTAIL.n324 VTAIL.n323 9.3005
R1801 VTAIL.n349 VTAIL.n348 9.3005
R1802 VTAIL.n312 VTAIL.n311 9.3005
R1803 VTAIL.n355 VTAIL.n354 9.3005
R1804 VTAIL.n357 VTAIL.n356 9.3005
R1805 VTAIL.n308 VTAIL.n307 9.3005
R1806 VTAIL.n363 VTAIL.n362 9.3005
R1807 VTAIL.n365 VTAIL.n364 9.3005
R1808 VTAIL.n366 VTAIL.n303 9.3005
R1809 VTAIL.n373 VTAIL.n372 9.3005
R1810 VTAIL.n95 VTAIL.n94 9.3005
R1811 VTAIL.n2 VTAIL.n1 9.3005
R1812 VTAIL.n89 VTAIL.n88 9.3005
R1813 VTAIL.n87 VTAIL.n86 9.3005
R1814 VTAIL.n6 VTAIL.n5 9.3005
R1815 VTAIL.n81 VTAIL.n80 9.3005
R1816 VTAIL.n53 VTAIL.n52 9.3005
R1817 VTAIL.n22 VTAIL.n21 9.3005
R1818 VTAIL.n47 VTAIL.n46 9.3005
R1819 VTAIL.n45 VTAIL.n44 9.3005
R1820 VTAIL.n26 VTAIL.n25 9.3005
R1821 VTAIL.n39 VTAIL.n38 9.3005
R1822 VTAIL.n37 VTAIL.n36 9.3005
R1823 VTAIL.n30 VTAIL.n29 9.3005
R1824 VTAIL.n55 VTAIL.n54 9.3005
R1825 VTAIL.n18 VTAIL.n17 9.3005
R1826 VTAIL.n61 VTAIL.n60 9.3005
R1827 VTAIL.n63 VTAIL.n62 9.3005
R1828 VTAIL.n14 VTAIL.n13 9.3005
R1829 VTAIL.n69 VTAIL.n68 9.3005
R1830 VTAIL.n71 VTAIL.n70 9.3005
R1831 VTAIL.n72 VTAIL.n9 9.3005
R1832 VTAIL.n79 VTAIL.n78 9.3005
R1833 VTAIL.n216 VTAIL.n215 9.3005
R1834 VTAIL.n259 VTAIL.n258 9.3005
R1835 VTAIL.n261 VTAIL.n260 9.3005
R1836 VTAIL.n212 VTAIL.n211 9.3005
R1837 VTAIL.n267 VTAIL.n266 9.3005
R1838 VTAIL.n269 VTAIL.n268 9.3005
R1839 VTAIL.n207 VTAIL.n205 9.3005
R1840 VTAIL.n275 VTAIL.n274 9.3005
R1841 VTAIL.n291 VTAIL.n290 9.3005
R1842 VTAIL.n198 VTAIL.n197 9.3005
R1843 VTAIL.n285 VTAIL.n284 9.3005
R1844 VTAIL.n283 VTAIL.n282 9.3005
R1845 VTAIL.n202 VTAIL.n201 9.3005
R1846 VTAIL.n277 VTAIL.n276 9.3005
R1847 VTAIL.n253 VTAIL.n252 9.3005
R1848 VTAIL.n251 VTAIL.n250 9.3005
R1849 VTAIL.n220 VTAIL.n219 9.3005
R1850 VTAIL.n245 VTAIL.n244 9.3005
R1851 VTAIL.n243 VTAIL.n242 9.3005
R1852 VTAIL.n224 VTAIL.n223 9.3005
R1853 VTAIL.n237 VTAIL.n236 9.3005
R1854 VTAIL.n235 VTAIL.n234 9.3005
R1855 VTAIL.n228 VTAIL.n227 9.3005
R1856 VTAIL.n118 VTAIL.n117 9.3005
R1857 VTAIL.n161 VTAIL.n160 9.3005
R1858 VTAIL.n163 VTAIL.n162 9.3005
R1859 VTAIL.n114 VTAIL.n113 9.3005
R1860 VTAIL.n169 VTAIL.n168 9.3005
R1861 VTAIL.n171 VTAIL.n170 9.3005
R1862 VTAIL.n109 VTAIL.n107 9.3005
R1863 VTAIL.n177 VTAIL.n176 9.3005
R1864 VTAIL.n193 VTAIL.n192 9.3005
R1865 VTAIL.n100 VTAIL.n99 9.3005
R1866 VTAIL.n187 VTAIL.n186 9.3005
R1867 VTAIL.n185 VTAIL.n184 9.3005
R1868 VTAIL.n104 VTAIL.n103 9.3005
R1869 VTAIL.n179 VTAIL.n178 9.3005
R1870 VTAIL.n155 VTAIL.n154 9.3005
R1871 VTAIL.n153 VTAIL.n152 9.3005
R1872 VTAIL.n122 VTAIL.n121 9.3005
R1873 VTAIL.n147 VTAIL.n146 9.3005
R1874 VTAIL.n145 VTAIL.n144 9.3005
R1875 VTAIL.n126 VTAIL.n125 9.3005
R1876 VTAIL.n139 VTAIL.n138 9.3005
R1877 VTAIL.n137 VTAIL.n136 9.3005
R1878 VTAIL.n130 VTAIL.n129 9.3005
R1879 VTAIL.n342 VTAIL.n341 8.92171
R1880 VTAIL.n357 VTAIL.n310 8.92171
R1881 VTAIL.n388 VTAIL.n294 8.92171
R1882 VTAIL.n48 VTAIL.n47 8.92171
R1883 VTAIL.n63 VTAIL.n16 8.92171
R1884 VTAIL.n94 VTAIL.n0 8.92171
R1885 VTAIL.n290 VTAIL.n196 8.92171
R1886 VTAIL.n261 VTAIL.n214 8.92171
R1887 VTAIL.n246 VTAIL.n245 8.92171
R1888 VTAIL.n192 VTAIL.n98 8.92171
R1889 VTAIL.n163 VTAIL.n116 8.92171
R1890 VTAIL.n148 VTAIL.n147 8.92171
R1891 VTAIL.n345 VTAIL.n316 8.14595
R1892 VTAIL.n354 VTAIL.n353 8.14595
R1893 VTAIL.n51 VTAIL.n22 8.14595
R1894 VTAIL.n60 VTAIL.n59 8.14595
R1895 VTAIL.n258 VTAIL.n257 8.14595
R1896 VTAIL.n249 VTAIL.n220 8.14595
R1897 VTAIL.n160 VTAIL.n159 8.14595
R1898 VTAIL.n151 VTAIL.n122 8.14595
R1899 VTAIL.n346 VTAIL.n314 7.3702
R1900 VTAIL.n350 VTAIL.n312 7.3702
R1901 VTAIL.n52 VTAIL.n20 7.3702
R1902 VTAIL.n56 VTAIL.n18 7.3702
R1903 VTAIL.n254 VTAIL.n216 7.3702
R1904 VTAIL.n250 VTAIL.n218 7.3702
R1905 VTAIL.n156 VTAIL.n118 7.3702
R1906 VTAIL.n152 VTAIL.n120 7.3702
R1907 VTAIL.n349 VTAIL.n314 6.59444
R1908 VTAIL.n350 VTAIL.n349 6.59444
R1909 VTAIL.n55 VTAIL.n20 6.59444
R1910 VTAIL.n56 VTAIL.n55 6.59444
R1911 VTAIL.n254 VTAIL.n253 6.59444
R1912 VTAIL.n253 VTAIL.n218 6.59444
R1913 VTAIL.n156 VTAIL.n155 6.59444
R1914 VTAIL.n155 VTAIL.n120 6.59444
R1915 VTAIL.n346 VTAIL.n345 5.81868
R1916 VTAIL.n353 VTAIL.n312 5.81868
R1917 VTAIL.n52 VTAIL.n51 5.81868
R1918 VTAIL.n59 VTAIL.n18 5.81868
R1919 VTAIL.n257 VTAIL.n216 5.81868
R1920 VTAIL.n250 VTAIL.n249 5.81868
R1921 VTAIL.n159 VTAIL.n118 5.81868
R1922 VTAIL.n152 VTAIL.n151 5.81868
R1923 VTAIL.n342 VTAIL.n316 5.04292
R1924 VTAIL.n354 VTAIL.n310 5.04292
R1925 VTAIL.n390 VTAIL.n294 5.04292
R1926 VTAIL.n48 VTAIL.n22 5.04292
R1927 VTAIL.n60 VTAIL.n16 5.04292
R1928 VTAIL.n96 VTAIL.n0 5.04292
R1929 VTAIL.n292 VTAIL.n196 5.04292
R1930 VTAIL.n258 VTAIL.n214 5.04292
R1931 VTAIL.n246 VTAIL.n220 5.04292
R1932 VTAIL.n194 VTAIL.n98 5.04292
R1933 VTAIL.n160 VTAIL.n116 5.04292
R1934 VTAIL.n148 VTAIL.n122 5.04292
R1935 VTAIL.n325 VTAIL.n323 4.38563
R1936 VTAIL.n31 VTAIL.n29 4.38563
R1937 VTAIL.n229 VTAIL.n227 4.38563
R1938 VTAIL.n131 VTAIL.n129 4.38563
R1939 VTAIL.n341 VTAIL.n318 4.26717
R1940 VTAIL.n358 VTAIL.n357 4.26717
R1941 VTAIL.n388 VTAIL.n387 4.26717
R1942 VTAIL.n47 VTAIL.n24 4.26717
R1943 VTAIL.n64 VTAIL.n63 4.26717
R1944 VTAIL.n94 VTAIL.n93 4.26717
R1945 VTAIL.n290 VTAIL.n289 4.26717
R1946 VTAIL.n262 VTAIL.n261 4.26717
R1947 VTAIL.n245 VTAIL.n222 4.26717
R1948 VTAIL.n192 VTAIL.n191 4.26717
R1949 VTAIL.n164 VTAIL.n163 4.26717
R1950 VTAIL.n147 VTAIL.n124 4.26717
R1951 VTAIL.n338 VTAIL.n337 3.49141
R1952 VTAIL.n361 VTAIL.n308 3.49141
R1953 VTAIL.n384 VTAIL.n296 3.49141
R1954 VTAIL.n44 VTAIL.n43 3.49141
R1955 VTAIL.n67 VTAIL.n14 3.49141
R1956 VTAIL.n90 VTAIL.n2 3.49141
R1957 VTAIL.n286 VTAIL.n198 3.49141
R1958 VTAIL.n265 VTAIL.n212 3.49141
R1959 VTAIL.n242 VTAIL.n241 3.49141
R1960 VTAIL.n188 VTAIL.n100 3.49141
R1961 VTAIL.n167 VTAIL.n114 3.49141
R1962 VTAIL.n144 VTAIL.n143 3.49141
R1963 VTAIL.n334 VTAIL.n320 2.71565
R1964 VTAIL.n362 VTAIL.n306 2.71565
R1965 VTAIL.n383 VTAIL.n298 2.71565
R1966 VTAIL.n40 VTAIL.n26 2.71565
R1967 VTAIL.n68 VTAIL.n12 2.71565
R1968 VTAIL.n89 VTAIL.n4 2.71565
R1969 VTAIL.n285 VTAIL.n200 2.71565
R1970 VTAIL.n266 VTAIL.n210 2.71565
R1971 VTAIL.n238 VTAIL.n224 2.71565
R1972 VTAIL.n187 VTAIL.n102 2.71565
R1973 VTAIL.n168 VTAIL.n112 2.71565
R1974 VTAIL.n140 VTAIL.n126 2.71565
R1975 VTAIL.n333 VTAIL.n322 1.93989
R1976 VTAIL.n367 VTAIL.n365 1.93989
R1977 VTAIL.n380 VTAIL.n379 1.93989
R1978 VTAIL.n39 VTAIL.n28 1.93989
R1979 VTAIL.n73 VTAIL.n71 1.93989
R1980 VTAIL.n86 VTAIL.n85 1.93989
R1981 VTAIL.n282 VTAIL.n281 1.93989
R1982 VTAIL.n270 VTAIL.n269 1.93989
R1983 VTAIL.n237 VTAIL.n226 1.93989
R1984 VTAIL.n184 VTAIL.n183 1.93989
R1985 VTAIL.n172 VTAIL.n171 1.93989
R1986 VTAIL.n139 VTAIL.n128 1.93989
R1987 VTAIL.n293 VTAIL.n195 1.79791
R1988 VTAIL VTAIL.n97 1.19231
R1989 VTAIL.n330 VTAIL.n329 1.16414
R1990 VTAIL.n366 VTAIL.n304 1.16414
R1991 VTAIL.n376 VTAIL.n300 1.16414
R1992 VTAIL.n36 VTAIL.n35 1.16414
R1993 VTAIL.n72 VTAIL.n10 1.16414
R1994 VTAIL.n82 VTAIL.n6 1.16414
R1995 VTAIL.n278 VTAIL.n202 1.16414
R1996 VTAIL.n273 VTAIL.n207 1.16414
R1997 VTAIL.n234 VTAIL.n233 1.16414
R1998 VTAIL.n180 VTAIL.n104 1.16414
R1999 VTAIL.n175 VTAIL.n109 1.16414
R2000 VTAIL.n136 VTAIL.n135 1.16414
R2001 VTAIL VTAIL.n391 0.606103
R2002 VTAIL.n326 VTAIL.n324 0.388379
R2003 VTAIL.n372 VTAIL.n371 0.388379
R2004 VTAIL.n375 VTAIL.n302 0.388379
R2005 VTAIL.n32 VTAIL.n30 0.388379
R2006 VTAIL.n78 VTAIL.n77 0.388379
R2007 VTAIL.n81 VTAIL.n8 0.388379
R2008 VTAIL.n277 VTAIL.n204 0.388379
R2009 VTAIL.n274 VTAIL.n206 0.388379
R2010 VTAIL.n230 VTAIL.n228 0.388379
R2011 VTAIL.n179 VTAIL.n106 0.388379
R2012 VTAIL.n176 VTAIL.n108 0.388379
R2013 VTAIL.n132 VTAIL.n130 0.388379
R2014 VTAIL.n331 VTAIL.n323 0.155672
R2015 VTAIL.n332 VTAIL.n331 0.155672
R2016 VTAIL.n332 VTAIL.n319 0.155672
R2017 VTAIL.n339 VTAIL.n319 0.155672
R2018 VTAIL.n340 VTAIL.n339 0.155672
R2019 VTAIL.n340 VTAIL.n315 0.155672
R2020 VTAIL.n347 VTAIL.n315 0.155672
R2021 VTAIL.n348 VTAIL.n347 0.155672
R2022 VTAIL.n348 VTAIL.n311 0.155672
R2023 VTAIL.n355 VTAIL.n311 0.155672
R2024 VTAIL.n356 VTAIL.n355 0.155672
R2025 VTAIL.n356 VTAIL.n307 0.155672
R2026 VTAIL.n363 VTAIL.n307 0.155672
R2027 VTAIL.n364 VTAIL.n363 0.155672
R2028 VTAIL.n364 VTAIL.n303 0.155672
R2029 VTAIL.n373 VTAIL.n303 0.155672
R2030 VTAIL.n374 VTAIL.n373 0.155672
R2031 VTAIL.n374 VTAIL.n299 0.155672
R2032 VTAIL.n381 VTAIL.n299 0.155672
R2033 VTAIL.n382 VTAIL.n381 0.155672
R2034 VTAIL.n382 VTAIL.n295 0.155672
R2035 VTAIL.n389 VTAIL.n295 0.155672
R2036 VTAIL.n37 VTAIL.n29 0.155672
R2037 VTAIL.n38 VTAIL.n37 0.155672
R2038 VTAIL.n38 VTAIL.n25 0.155672
R2039 VTAIL.n45 VTAIL.n25 0.155672
R2040 VTAIL.n46 VTAIL.n45 0.155672
R2041 VTAIL.n46 VTAIL.n21 0.155672
R2042 VTAIL.n53 VTAIL.n21 0.155672
R2043 VTAIL.n54 VTAIL.n53 0.155672
R2044 VTAIL.n54 VTAIL.n17 0.155672
R2045 VTAIL.n61 VTAIL.n17 0.155672
R2046 VTAIL.n62 VTAIL.n61 0.155672
R2047 VTAIL.n62 VTAIL.n13 0.155672
R2048 VTAIL.n69 VTAIL.n13 0.155672
R2049 VTAIL.n70 VTAIL.n69 0.155672
R2050 VTAIL.n70 VTAIL.n9 0.155672
R2051 VTAIL.n79 VTAIL.n9 0.155672
R2052 VTAIL.n80 VTAIL.n79 0.155672
R2053 VTAIL.n80 VTAIL.n5 0.155672
R2054 VTAIL.n87 VTAIL.n5 0.155672
R2055 VTAIL.n88 VTAIL.n87 0.155672
R2056 VTAIL.n88 VTAIL.n1 0.155672
R2057 VTAIL.n95 VTAIL.n1 0.155672
R2058 VTAIL.n291 VTAIL.n197 0.155672
R2059 VTAIL.n284 VTAIL.n197 0.155672
R2060 VTAIL.n284 VTAIL.n283 0.155672
R2061 VTAIL.n283 VTAIL.n201 0.155672
R2062 VTAIL.n276 VTAIL.n201 0.155672
R2063 VTAIL.n276 VTAIL.n275 0.155672
R2064 VTAIL.n275 VTAIL.n205 0.155672
R2065 VTAIL.n268 VTAIL.n205 0.155672
R2066 VTAIL.n268 VTAIL.n267 0.155672
R2067 VTAIL.n267 VTAIL.n211 0.155672
R2068 VTAIL.n260 VTAIL.n211 0.155672
R2069 VTAIL.n260 VTAIL.n259 0.155672
R2070 VTAIL.n259 VTAIL.n215 0.155672
R2071 VTAIL.n252 VTAIL.n215 0.155672
R2072 VTAIL.n252 VTAIL.n251 0.155672
R2073 VTAIL.n251 VTAIL.n219 0.155672
R2074 VTAIL.n244 VTAIL.n219 0.155672
R2075 VTAIL.n244 VTAIL.n243 0.155672
R2076 VTAIL.n243 VTAIL.n223 0.155672
R2077 VTAIL.n236 VTAIL.n223 0.155672
R2078 VTAIL.n236 VTAIL.n235 0.155672
R2079 VTAIL.n235 VTAIL.n227 0.155672
R2080 VTAIL.n193 VTAIL.n99 0.155672
R2081 VTAIL.n186 VTAIL.n99 0.155672
R2082 VTAIL.n186 VTAIL.n185 0.155672
R2083 VTAIL.n185 VTAIL.n103 0.155672
R2084 VTAIL.n178 VTAIL.n103 0.155672
R2085 VTAIL.n178 VTAIL.n177 0.155672
R2086 VTAIL.n177 VTAIL.n107 0.155672
R2087 VTAIL.n170 VTAIL.n107 0.155672
R2088 VTAIL.n170 VTAIL.n169 0.155672
R2089 VTAIL.n169 VTAIL.n113 0.155672
R2090 VTAIL.n162 VTAIL.n113 0.155672
R2091 VTAIL.n162 VTAIL.n161 0.155672
R2092 VTAIL.n161 VTAIL.n117 0.155672
R2093 VTAIL.n154 VTAIL.n117 0.155672
R2094 VTAIL.n154 VTAIL.n153 0.155672
R2095 VTAIL.n153 VTAIL.n121 0.155672
R2096 VTAIL.n146 VTAIL.n121 0.155672
R2097 VTAIL.n146 VTAIL.n145 0.155672
R2098 VTAIL.n145 VTAIL.n125 0.155672
R2099 VTAIL.n138 VTAIL.n125 0.155672
R2100 VTAIL.n138 VTAIL.n137 0.155672
R2101 VTAIL.n137 VTAIL.n129 0.155672
R2102 VDD2.n189 VDD2.n97 289.615
R2103 VDD2.n92 VDD2.n0 289.615
R2104 VDD2.n190 VDD2.n189 185
R2105 VDD2.n188 VDD2.n187 185
R2106 VDD2.n101 VDD2.n100 185
R2107 VDD2.n182 VDD2.n181 185
R2108 VDD2.n180 VDD2.n179 185
R2109 VDD2.n105 VDD2.n104 185
R2110 VDD2.n109 VDD2.n107 185
R2111 VDD2.n174 VDD2.n173 185
R2112 VDD2.n172 VDD2.n171 185
R2113 VDD2.n111 VDD2.n110 185
R2114 VDD2.n166 VDD2.n165 185
R2115 VDD2.n164 VDD2.n163 185
R2116 VDD2.n115 VDD2.n114 185
R2117 VDD2.n158 VDD2.n157 185
R2118 VDD2.n156 VDD2.n155 185
R2119 VDD2.n119 VDD2.n118 185
R2120 VDD2.n150 VDD2.n149 185
R2121 VDD2.n148 VDD2.n147 185
R2122 VDD2.n123 VDD2.n122 185
R2123 VDD2.n142 VDD2.n141 185
R2124 VDD2.n140 VDD2.n139 185
R2125 VDD2.n127 VDD2.n126 185
R2126 VDD2.n134 VDD2.n133 185
R2127 VDD2.n132 VDD2.n131 185
R2128 VDD2.n33 VDD2.n32 185
R2129 VDD2.n35 VDD2.n34 185
R2130 VDD2.n28 VDD2.n27 185
R2131 VDD2.n41 VDD2.n40 185
R2132 VDD2.n43 VDD2.n42 185
R2133 VDD2.n24 VDD2.n23 185
R2134 VDD2.n49 VDD2.n48 185
R2135 VDD2.n51 VDD2.n50 185
R2136 VDD2.n20 VDD2.n19 185
R2137 VDD2.n57 VDD2.n56 185
R2138 VDD2.n59 VDD2.n58 185
R2139 VDD2.n16 VDD2.n15 185
R2140 VDD2.n65 VDD2.n64 185
R2141 VDD2.n67 VDD2.n66 185
R2142 VDD2.n12 VDD2.n11 185
R2143 VDD2.n74 VDD2.n73 185
R2144 VDD2.n75 VDD2.n10 185
R2145 VDD2.n77 VDD2.n76 185
R2146 VDD2.n8 VDD2.n7 185
R2147 VDD2.n83 VDD2.n82 185
R2148 VDD2.n85 VDD2.n84 185
R2149 VDD2.n4 VDD2.n3 185
R2150 VDD2.n91 VDD2.n90 185
R2151 VDD2.n93 VDD2.n92 185
R2152 VDD2.n130 VDD2.t0 147.659
R2153 VDD2.n31 VDD2.t1 147.659
R2154 VDD2.n189 VDD2.n188 104.615
R2155 VDD2.n188 VDD2.n100 104.615
R2156 VDD2.n181 VDD2.n100 104.615
R2157 VDD2.n181 VDD2.n180 104.615
R2158 VDD2.n180 VDD2.n104 104.615
R2159 VDD2.n109 VDD2.n104 104.615
R2160 VDD2.n173 VDD2.n109 104.615
R2161 VDD2.n173 VDD2.n172 104.615
R2162 VDD2.n172 VDD2.n110 104.615
R2163 VDD2.n165 VDD2.n110 104.615
R2164 VDD2.n165 VDD2.n164 104.615
R2165 VDD2.n164 VDD2.n114 104.615
R2166 VDD2.n157 VDD2.n114 104.615
R2167 VDD2.n157 VDD2.n156 104.615
R2168 VDD2.n156 VDD2.n118 104.615
R2169 VDD2.n149 VDD2.n118 104.615
R2170 VDD2.n149 VDD2.n148 104.615
R2171 VDD2.n148 VDD2.n122 104.615
R2172 VDD2.n141 VDD2.n122 104.615
R2173 VDD2.n141 VDD2.n140 104.615
R2174 VDD2.n140 VDD2.n126 104.615
R2175 VDD2.n133 VDD2.n126 104.615
R2176 VDD2.n133 VDD2.n132 104.615
R2177 VDD2.n34 VDD2.n33 104.615
R2178 VDD2.n34 VDD2.n27 104.615
R2179 VDD2.n41 VDD2.n27 104.615
R2180 VDD2.n42 VDD2.n41 104.615
R2181 VDD2.n42 VDD2.n23 104.615
R2182 VDD2.n49 VDD2.n23 104.615
R2183 VDD2.n50 VDD2.n49 104.615
R2184 VDD2.n50 VDD2.n19 104.615
R2185 VDD2.n57 VDD2.n19 104.615
R2186 VDD2.n58 VDD2.n57 104.615
R2187 VDD2.n58 VDD2.n15 104.615
R2188 VDD2.n65 VDD2.n15 104.615
R2189 VDD2.n66 VDD2.n65 104.615
R2190 VDD2.n66 VDD2.n11 104.615
R2191 VDD2.n74 VDD2.n11 104.615
R2192 VDD2.n75 VDD2.n74 104.615
R2193 VDD2.n76 VDD2.n75 104.615
R2194 VDD2.n76 VDD2.n7 104.615
R2195 VDD2.n83 VDD2.n7 104.615
R2196 VDD2.n84 VDD2.n83 104.615
R2197 VDD2.n84 VDD2.n3 104.615
R2198 VDD2.n91 VDD2.n3 104.615
R2199 VDD2.n92 VDD2.n91 104.615
R2200 VDD2.n194 VDD2.n96 93.1399
R2201 VDD2.n132 VDD2.t0 52.3082
R2202 VDD2.n33 VDD2.t1 52.3082
R2203 VDD2.n194 VDD2.n193 49.0581
R2204 VDD2.n131 VDD2.n130 15.6677
R2205 VDD2.n32 VDD2.n31 15.6677
R2206 VDD2.n107 VDD2.n105 13.1884
R2207 VDD2.n77 VDD2.n8 13.1884
R2208 VDD2.n179 VDD2.n178 12.8005
R2209 VDD2.n175 VDD2.n174 12.8005
R2210 VDD2.n134 VDD2.n129 12.8005
R2211 VDD2.n35 VDD2.n30 12.8005
R2212 VDD2.n78 VDD2.n10 12.8005
R2213 VDD2.n82 VDD2.n81 12.8005
R2214 VDD2.n182 VDD2.n103 12.0247
R2215 VDD2.n171 VDD2.n108 12.0247
R2216 VDD2.n135 VDD2.n127 12.0247
R2217 VDD2.n36 VDD2.n28 12.0247
R2218 VDD2.n73 VDD2.n72 12.0247
R2219 VDD2.n85 VDD2.n6 12.0247
R2220 VDD2.n183 VDD2.n101 11.249
R2221 VDD2.n170 VDD2.n111 11.249
R2222 VDD2.n139 VDD2.n138 11.249
R2223 VDD2.n40 VDD2.n39 11.249
R2224 VDD2.n71 VDD2.n12 11.249
R2225 VDD2.n86 VDD2.n4 11.249
R2226 VDD2.n187 VDD2.n186 10.4732
R2227 VDD2.n167 VDD2.n166 10.4732
R2228 VDD2.n142 VDD2.n125 10.4732
R2229 VDD2.n43 VDD2.n26 10.4732
R2230 VDD2.n68 VDD2.n67 10.4732
R2231 VDD2.n90 VDD2.n89 10.4732
R2232 VDD2.n190 VDD2.n99 9.69747
R2233 VDD2.n163 VDD2.n113 9.69747
R2234 VDD2.n143 VDD2.n123 9.69747
R2235 VDD2.n44 VDD2.n24 9.69747
R2236 VDD2.n64 VDD2.n14 9.69747
R2237 VDD2.n93 VDD2.n2 9.69747
R2238 VDD2.n193 VDD2.n192 9.45567
R2239 VDD2.n96 VDD2.n95 9.45567
R2240 VDD2.n117 VDD2.n116 9.3005
R2241 VDD2.n160 VDD2.n159 9.3005
R2242 VDD2.n162 VDD2.n161 9.3005
R2243 VDD2.n113 VDD2.n112 9.3005
R2244 VDD2.n168 VDD2.n167 9.3005
R2245 VDD2.n170 VDD2.n169 9.3005
R2246 VDD2.n108 VDD2.n106 9.3005
R2247 VDD2.n176 VDD2.n175 9.3005
R2248 VDD2.n192 VDD2.n191 9.3005
R2249 VDD2.n99 VDD2.n98 9.3005
R2250 VDD2.n186 VDD2.n185 9.3005
R2251 VDD2.n184 VDD2.n183 9.3005
R2252 VDD2.n103 VDD2.n102 9.3005
R2253 VDD2.n178 VDD2.n177 9.3005
R2254 VDD2.n154 VDD2.n153 9.3005
R2255 VDD2.n152 VDD2.n151 9.3005
R2256 VDD2.n121 VDD2.n120 9.3005
R2257 VDD2.n146 VDD2.n145 9.3005
R2258 VDD2.n144 VDD2.n143 9.3005
R2259 VDD2.n125 VDD2.n124 9.3005
R2260 VDD2.n138 VDD2.n137 9.3005
R2261 VDD2.n136 VDD2.n135 9.3005
R2262 VDD2.n129 VDD2.n128 9.3005
R2263 VDD2.n95 VDD2.n94 9.3005
R2264 VDD2.n2 VDD2.n1 9.3005
R2265 VDD2.n89 VDD2.n88 9.3005
R2266 VDD2.n87 VDD2.n86 9.3005
R2267 VDD2.n6 VDD2.n5 9.3005
R2268 VDD2.n81 VDD2.n80 9.3005
R2269 VDD2.n53 VDD2.n52 9.3005
R2270 VDD2.n22 VDD2.n21 9.3005
R2271 VDD2.n47 VDD2.n46 9.3005
R2272 VDD2.n45 VDD2.n44 9.3005
R2273 VDD2.n26 VDD2.n25 9.3005
R2274 VDD2.n39 VDD2.n38 9.3005
R2275 VDD2.n37 VDD2.n36 9.3005
R2276 VDD2.n30 VDD2.n29 9.3005
R2277 VDD2.n55 VDD2.n54 9.3005
R2278 VDD2.n18 VDD2.n17 9.3005
R2279 VDD2.n61 VDD2.n60 9.3005
R2280 VDD2.n63 VDD2.n62 9.3005
R2281 VDD2.n14 VDD2.n13 9.3005
R2282 VDD2.n69 VDD2.n68 9.3005
R2283 VDD2.n71 VDD2.n70 9.3005
R2284 VDD2.n72 VDD2.n9 9.3005
R2285 VDD2.n79 VDD2.n78 9.3005
R2286 VDD2.n191 VDD2.n97 8.92171
R2287 VDD2.n162 VDD2.n115 8.92171
R2288 VDD2.n147 VDD2.n146 8.92171
R2289 VDD2.n48 VDD2.n47 8.92171
R2290 VDD2.n63 VDD2.n16 8.92171
R2291 VDD2.n94 VDD2.n0 8.92171
R2292 VDD2.n159 VDD2.n158 8.14595
R2293 VDD2.n150 VDD2.n121 8.14595
R2294 VDD2.n51 VDD2.n22 8.14595
R2295 VDD2.n60 VDD2.n59 8.14595
R2296 VDD2.n155 VDD2.n117 7.3702
R2297 VDD2.n151 VDD2.n119 7.3702
R2298 VDD2.n52 VDD2.n20 7.3702
R2299 VDD2.n56 VDD2.n18 7.3702
R2300 VDD2.n155 VDD2.n154 6.59444
R2301 VDD2.n154 VDD2.n119 6.59444
R2302 VDD2.n55 VDD2.n20 6.59444
R2303 VDD2.n56 VDD2.n55 6.59444
R2304 VDD2.n158 VDD2.n117 5.81868
R2305 VDD2.n151 VDD2.n150 5.81868
R2306 VDD2.n52 VDD2.n51 5.81868
R2307 VDD2.n59 VDD2.n18 5.81868
R2308 VDD2.n193 VDD2.n97 5.04292
R2309 VDD2.n159 VDD2.n115 5.04292
R2310 VDD2.n147 VDD2.n121 5.04292
R2311 VDD2.n48 VDD2.n22 5.04292
R2312 VDD2.n60 VDD2.n16 5.04292
R2313 VDD2.n96 VDD2.n0 5.04292
R2314 VDD2.n130 VDD2.n128 4.38563
R2315 VDD2.n31 VDD2.n29 4.38563
R2316 VDD2.n191 VDD2.n190 4.26717
R2317 VDD2.n163 VDD2.n162 4.26717
R2318 VDD2.n146 VDD2.n123 4.26717
R2319 VDD2.n47 VDD2.n24 4.26717
R2320 VDD2.n64 VDD2.n63 4.26717
R2321 VDD2.n94 VDD2.n93 4.26717
R2322 VDD2.n187 VDD2.n99 3.49141
R2323 VDD2.n166 VDD2.n113 3.49141
R2324 VDD2.n143 VDD2.n142 3.49141
R2325 VDD2.n44 VDD2.n43 3.49141
R2326 VDD2.n67 VDD2.n14 3.49141
R2327 VDD2.n90 VDD2.n2 3.49141
R2328 VDD2.n186 VDD2.n101 2.71565
R2329 VDD2.n167 VDD2.n111 2.71565
R2330 VDD2.n139 VDD2.n125 2.71565
R2331 VDD2.n40 VDD2.n26 2.71565
R2332 VDD2.n68 VDD2.n12 2.71565
R2333 VDD2.n89 VDD2.n4 2.71565
R2334 VDD2.n183 VDD2.n182 1.93989
R2335 VDD2.n171 VDD2.n170 1.93989
R2336 VDD2.n138 VDD2.n127 1.93989
R2337 VDD2.n39 VDD2.n28 1.93989
R2338 VDD2.n73 VDD2.n71 1.93989
R2339 VDD2.n86 VDD2.n85 1.93989
R2340 VDD2.n179 VDD2.n103 1.16414
R2341 VDD2.n174 VDD2.n108 1.16414
R2342 VDD2.n135 VDD2.n134 1.16414
R2343 VDD2.n36 VDD2.n35 1.16414
R2344 VDD2.n72 VDD2.n10 1.16414
R2345 VDD2.n82 VDD2.n6 1.16414
R2346 VDD2 VDD2.n194 0.722483
R2347 VDD2.n178 VDD2.n105 0.388379
R2348 VDD2.n175 VDD2.n107 0.388379
R2349 VDD2.n131 VDD2.n129 0.388379
R2350 VDD2.n32 VDD2.n30 0.388379
R2351 VDD2.n78 VDD2.n77 0.388379
R2352 VDD2.n81 VDD2.n8 0.388379
R2353 VDD2.n192 VDD2.n98 0.155672
R2354 VDD2.n185 VDD2.n98 0.155672
R2355 VDD2.n185 VDD2.n184 0.155672
R2356 VDD2.n184 VDD2.n102 0.155672
R2357 VDD2.n177 VDD2.n102 0.155672
R2358 VDD2.n177 VDD2.n176 0.155672
R2359 VDD2.n176 VDD2.n106 0.155672
R2360 VDD2.n169 VDD2.n106 0.155672
R2361 VDD2.n169 VDD2.n168 0.155672
R2362 VDD2.n168 VDD2.n112 0.155672
R2363 VDD2.n161 VDD2.n112 0.155672
R2364 VDD2.n161 VDD2.n160 0.155672
R2365 VDD2.n160 VDD2.n116 0.155672
R2366 VDD2.n153 VDD2.n116 0.155672
R2367 VDD2.n153 VDD2.n152 0.155672
R2368 VDD2.n152 VDD2.n120 0.155672
R2369 VDD2.n145 VDD2.n120 0.155672
R2370 VDD2.n145 VDD2.n144 0.155672
R2371 VDD2.n144 VDD2.n124 0.155672
R2372 VDD2.n137 VDD2.n124 0.155672
R2373 VDD2.n137 VDD2.n136 0.155672
R2374 VDD2.n136 VDD2.n128 0.155672
R2375 VDD2.n37 VDD2.n29 0.155672
R2376 VDD2.n38 VDD2.n37 0.155672
R2377 VDD2.n38 VDD2.n25 0.155672
R2378 VDD2.n45 VDD2.n25 0.155672
R2379 VDD2.n46 VDD2.n45 0.155672
R2380 VDD2.n46 VDD2.n21 0.155672
R2381 VDD2.n53 VDD2.n21 0.155672
R2382 VDD2.n54 VDD2.n53 0.155672
R2383 VDD2.n54 VDD2.n17 0.155672
R2384 VDD2.n61 VDD2.n17 0.155672
R2385 VDD2.n62 VDD2.n61 0.155672
R2386 VDD2.n62 VDD2.n13 0.155672
R2387 VDD2.n69 VDD2.n13 0.155672
R2388 VDD2.n70 VDD2.n69 0.155672
R2389 VDD2.n70 VDD2.n9 0.155672
R2390 VDD2.n79 VDD2.n9 0.155672
R2391 VDD2.n80 VDD2.n79 0.155672
R2392 VDD2.n80 VDD2.n5 0.155672
R2393 VDD2.n87 VDD2.n5 0.155672
R2394 VDD2.n88 VDD2.n87 0.155672
R2395 VDD2.n88 VDD2.n1 0.155672
R2396 VDD2.n95 VDD2.n1 0.155672
R2397 VP.n0 VP.t1 243.966
R2398 VP.n0 VP.t0 194.722
R2399 VP VP.n0 0.431811
R2400 VDD1.n92 VDD1.n0 289.615
R2401 VDD1.n189 VDD1.n97 289.615
R2402 VDD1.n93 VDD1.n92 185
R2403 VDD1.n91 VDD1.n90 185
R2404 VDD1.n4 VDD1.n3 185
R2405 VDD1.n85 VDD1.n84 185
R2406 VDD1.n83 VDD1.n82 185
R2407 VDD1.n8 VDD1.n7 185
R2408 VDD1.n12 VDD1.n10 185
R2409 VDD1.n77 VDD1.n76 185
R2410 VDD1.n75 VDD1.n74 185
R2411 VDD1.n14 VDD1.n13 185
R2412 VDD1.n69 VDD1.n68 185
R2413 VDD1.n67 VDD1.n66 185
R2414 VDD1.n18 VDD1.n17 185
R2415 VDD1.n61 VDD1.n60 185
R2416 VDD1.n59 VDD1.n58 185
R2417 VDD1.n22 VDD1.n21 185
R2418 VDD1.n53 VDD1.n52 185
R2419 VDD1.n51 VDD1.n50 185
R2420 VDD1.n26 VDD1.n25 185
R2421 VDD1.n45 VDD1.n44 185
R2422 VDD1.n43 VDD1.n42 185
R2423 VDD1.n30 VDD1.n29 185
R2424 VDD1.n37 VDD1.n36 185
R2425 VDD1.n35 VDD1.n34 185
R2426 VDD1.n130 VDD1.n129 185
R2427 VDD1.n132 VDD1.n131 185
R2428 VDD1.n125 VDD1.n124 185
R2429 VDD1.n138 VDD1.n137 185
R2430 VDD1.n140 VDD1.n139 185
R2431 VDD1.n121 VDD1.n120 185
R2432 VDD1.n146 VDD1.n145 185
R2433 VDD1.n148 VDD1.n147 185
R2434 VDD1.n117 VDD1.n116 185
R2435 VDD1.n154 VDD1.n153 185
R2436 VDD1.n156 VDD1.n155 185
R2437 VDD1.n113 VDD1.n112 185
R2438 VDD1.n162 VDD1.n161 185
R2439 VDD1.n164 VDD1.n163 185
R2440 VDD1.n109 VDD1.n108 185
R2441 VDD1.n171 VDD1.n170 185
R2442 VDD1.n172 VDD1.n107 185
R2443 VDD1.n174 VDD1.n173 185
R2444 VDD1.n105 VDD1.n104 185
R2445 VDD1.n180 VDD1.n179 185
R2446 VDD1.n182 VDD1.n181 185
R2447 VDD1.n101 VDD1.n100 185
R2448 VDD1.n188 VDD1.n187 185
R2449 VDD1.n190 VDD1.n189 185
R2450 VDD1.n33 VDD1.t0 147.659
R2451 VDD1.n128 VDD1.t1 147.659
R2452 VDD1.n92 VDD1.n91 104.615
R2453 VDD1.n91 VDD1.n3 104.615
R2454 VDD1.n84 VDD1.n3 104.615
R2455 VDD1.n84 VDD1.n83 104.615
R2456 VDD1.n83 VDD1.n7 104.615
R2457 VDD1.n12 VDD1.n7 104.615
R2458 VDD1.n76 VDD1.n12 104.615
R2459 VDD1.n76 VDD1.n75 104.615
R2460 VDD1.n75 VDD1.n13 104.615
R2461 VDD1.n68 VDD1.n13 104.615
R2462 VDD1.n68 VDD1.n67 104.615
R2463 VDD1.n67 VDD1.n17 104.615
R2464 VDD1.n60 VDD1.n17 104.615
R2465 VDD1.n60 VDD1.n59 104.615
R2466 VDD1.n59 VDD1.n21 104.615
R2467 VDD1.n52 VDD1.n21 104.615
R2468 VDD1.n52 VDD1.n51 104.615
R2469 VDD1.n51 VDD1.n25 104.615
R2470 VDD1.n44 VDD1.n25 104.615
R2471 VDD1.n44 VDD1.n43 104.615
R2472 VDD1.n43 VDD1.n29 104.615
R2473 VDD1.n36 VDD1.n29 104.615
R2474 VDD1.n36 VDD1.n35 104.615
R2475 VDD1.n131 VDD1.n130 104.615
R2476 VDD1.n131 VDD1.n124 104.615
R2477 VDD1.n138 VDD1.n124 104.615
R2478 VDD1.n139 VDD1.n138 104.615
R2479 VDD1.n139 VDD1.n120 104.615
R2480 VDD1.n146 VDD1.n120 104.615
R2481 VDD1.n147 VDD1.n146 104.615
R2482 VDD1.n147 VDD1.n116 104.615
R2483 VDD1.n154 VDD1.n116 104.615
R2484 VDD1.n155 VDD1.n154 104.615
R2485 VDD1.n155 VDD1.n112 104.615
R2486 VDD1.n162 VDD1.n112 104.615
R2487 VDD1.n163 VDD1.n162 104.615
R2488 VDD1.n163 VDD1.n108 104.615
R2489 VDD1.n171 VDD1.n108 104.615
R2490 VDD1.n172 VDD1.n171 104.615
R2491 VDD1.n173 VDD1.n172 104.615
R2492 VDD1.n173 VDD1.n104 104.615
R2493 VDD1.n180 VDD1.n104 104.615
R2494 VDD1.n181 VDD1.n180 104.615
R2495 VDD1.n181 VDD1.n100 104.615
R2496 VDD1.n188 VDD1.n100 104.615
R2497 VDD1.n189 VDD1.n188 104.615
R2498 VDD1 VDD1.n193 94.3286
R2499 VDD1.n35 VDD1.t0 52.3082
R2500 VDD1.n130 VDD1.t1 52.3082
R2501 VDD1 VDD1.n96 49.7801
R2502 VDD1.n34 VDD1.n33 15.6677
R2503 VDD1.n129 VDD1.n128 15.6677
R2504 VDD1.n10 VDD1.n8 13.1884
R2505 VDD1.n174 VDD1.n105 13.1884
R2506 VDD1.n82 VDD1.n81 12.8005
R2507 VDD1.n78 VDD1.n77 12.8005
R2508 VDD1.n37 VDD1.n32 12.8005
R2509 VDD1.n132 VDD1.n127 12.8005
R2510 VDD1.n175 VDD1.n107 12.8005
R2511 VDD1.n179 VDD1.n178 12.8005
R2512 VDD1.n85 VDD1.n6 12.0247
R2513 VDD1.n74 VDD1.n11 12.0247
R2514 VDD1.n38 VDD1.n30 12.0247
R2515 VDD1.n133 VDD1.n125 12.0247
R2516 VDD1.n170 VDD1.n169 12.0247
R2517 VDD1.n182 VDD1.n103 12.0247
R2518 VDD1.n86 VDD1.n4 11.249
R2519 VDD1.n73 VDD1.n14 11.249
R2520 VDD1.n42 VDD1.n41 11.249
R2521 VDD1.n137 VDD1.n136 11.249
R2522 VDD1.n168 VDD1.n109 11.249
R2523 VDD1.n183 VDD1.n101 11.249
R2524 VDD1.n90 VDD1.n89 10.4732
R2525 VDD1.n70 VDD1.n69 10.4732
R2526 VDD1.n45 VDD1.n28 10.4732
R2527 VDD1.n140 VDD1.n123 10.4732
R2528 VDD1.n165 VDD1.n164 10.4732
R2529 VDD1.n187 VDD1.n186 10.4732
R2530 VDD1.n93 VDD1.n2 9.69747
R2531 VDD1.n66 VDD1.n16 9.69747
R2532 VDD1.n46 VDD1.n26 9.69747
R2533 VDD1.n141 VDD1.n121 9.69747
R2534 VDD1.n161 VDD1.n111 9.69747
R2535 VDD1.n190 VDD1.n99 9.69747
R2536 VDD1.n96 VDD1.n95 9.45567
R2537 VDD1.n193 VDD1.n192 9.45567
R2538 VDD1.n20 VDD1.n19 9.3005
R2539 VDD1.n63 VDD1.n62 9.3005
R2540 VDD1.n65 VDD1.n64 9.3005
R2541 VDD1.n16 VDD1.n15 9.3005
R2542 VDD1.n71 VDD1.n70 9.3005
R2543 VDD1.n73 VDD1.n72 9.3005
R2544 VDD1.n11 VDD1.n9 9.3005
R2545 VDD1.n79 VDD1.n78 9.3005
R2546 VDD1.n95 VDD1.n94 9.3005
R2547 VDD1.n2 VDD1.n1 9.3005
R2548 VDD1.n89 VDD1.n88 9.3005
R2549 VDD1.n87 VDD1.n86 9.3005
R2550 VDD1.n6 VDD1.n5 9.3005
R2551 VDD1.n81 VDD1.n80 9.3005
R2552 VDD1.n57 VDD1.n56 9.3005
R2553 VDD1.n55 VDD1.n54 9.3005
R2554 VDD1.n24 VDD1.n23 9.3005
R2555 VDD1.n49 VDD1.n48 9.3005
R2556 VDD1.n47 VDD1.n46 9.3005
R2557 VDD1.n28 VDD1.n27 9.3005
R2558 VDD1.n41 VDD1.n40 9.3005
R2559 VDD1.n39 VDD1.n38 9.3005
R2560 VDD1.n32 VDD1.n31 9.3005
R2561 VDD1.n192 VDD1.n191 9.3005
R2562 VDD1.n99 VDD1.n98 9.3005
R2563 VDD1.n186 VDD1.n185 9.3005
R2564 VDD1.n184 VDD1.n183 9.3005
R2565 VDD1.n103 VDD1.n102 9.3005
R2566 VDD1.n178 VDD1.n177 9.3005
R2567 VDD1.n150 VDD1.n149 9.3005
R2568 VDD1.n119 VDD1.n118 9.3005
R2569 VDD1.n144 VDD1.n143 9.3005
R2570 VDD1.n142 VDD1.n141 9.3005
R2571 VDD1.n123 VDD1.n122 9.3005
R2572 VDD1.n136 VDD1.n135 9.3005
R2573 VDD1.n134 VDD1.n133 9.3005
R2574 VDD1.n127 VDD1.n126 9.3005
R2575 VDD1.n152 VDD1.n151 9.3005
R2576 VDD1.n115 VDD1.n114 9.3005
R2577 VDD1.n158 VDD1.n157 9.3005
R2578 VDD1.n160 VDD1.n159 9.3005
R2579 VDD1.n111 VDD1.n110 9.3005
R2580 VDD1.n166 VDD1.n165 9.3005
R2581 VDD1.n168 VDD1.n167 9.3005
R2582 VDD1.n169 VDD1.n106 9.3005
R2583 VDD1.n176 VDD1.n175 9.3005
R2584 VDD1.n94 VDD1.n0 8.92171
R2585 VDD1.n65 VDD1.n18 8.92171
R2586 VDD1.n50 VDD1.n49 8.92171
R2587 VDD1.n145 VDD1.n144 8.92171
R2588 VDD1.n160 VDD1.n113 8.92171
R2589 VDD1.n191 VDD1.n97 8.92171
R2590 VDD1.n62 VDD1.n61 8.14595
R2591 VDD1.n53 VDD1.n24 8.14595
R2592 VDD1.n148 VDD1.n119 8.14595
R2593 VDD1.n157 VDD1.n156 8.14595
R2594 VDD1.n58 VDD1.n20 7.3702
R2595 VDD1.n54 VDD1.n22 7.3702
R2596 VDD1.n149 VDD1.n117 7.3702
R2597 VDD1.n153 VDD1.n115 7.3702
R2598 VDD1.n58 VDD1.n57 6.59444
R2599 VDD1.n57 VDD1.n22 6.59444
R2600 VDD1.n152 VDD1.n117 6.59444
R2601 VDD1.n153 VDD1.n152 6.59444
R2602 VDD1.n61 VDD1.n20 5.81868
R2603 VDD1.n54 VDD1.n53 5.81868
R2604 VDD1.n149 VDD1.n148 5.81868
R2605 VDD1.n156 VDD1.n115 5.81868
R2606 VDD1.n96 VDD1.n0 5.04292
R2607 VDD1.n62 VDD1.n18 5.04292
R2608 VDD1.n50 VDD1.n24 5.04292
R2609 VDD1.n145 VDD1.n119 5.04292
R2610 VDD1.n157 VDD1.n113 5.04292
R2611 VDD1.n193 VDD1.n97 5.04292
R2612 VDD1.n33 VDD1.n31 4.38563
R2613 VDD1.n128 VDD1.n126 4.38563
R2614 VDD1.n94 VDD1.n93 4.26717
R2615 VDD1.n66 VDD1.n65 4.26717
R2616 VDD1.n49 VDD1.n26 4.26717
R2617 VDD1.n144 VDD1.n121 4.26717
R2618 VDD1.n161 VDD1.n160 4.26717
R2619 VDD1.n191 VDD1.n190 4.26717
R2620 VDD1.n90 VDD1.n2 3.49141
R2621 VDD1.n69 VDD1.n16 3.49141
R2622 VDD1.n46 VDD1.n45 3.49141
R2623 VDD1.n141 VDD1.n140 3.49141
R2624 VDD1.n164 VDD1.n111 3.49141
R2625 VDD1.n187 VDD1.n99 3.49141
R2626 VDD1.n89 VDD1.n4 2.71565
R2627 VDD1.n70 VDD1.n14 2.71565
R2628 VDD1.n42 VDD1.n28 2.71565
R2629 VDD1.n137 VDD1.n123 2.71565
R2630 VDD1.n165 VDD1.n109 2.71565
R2631 VDD1.n186 VDD1.n101 2.71565
R2632 VDD1.n86 VDD1.n85 1.93989
R2633 VDD1.n74 VDD1.n73 1.93989
R2634 VDD1.n41 VDD1.n30 1.93989
R2635 VDD1.n136 VDD1.n125 1.93989
R2636 VDD1.n170 VDD1.n168 1.93989
R2637 VDD1.n183 VDD1.n182 1.93989
R2638 VDD1.n82 VDD1.n6 1.16414
R2639 VDD1.n77 VDD1.n11 1.16414
R2640 VDD1.n38 VDD1.n37 1.16414
R2641 VDD1.n133 VDD1.n132 1.16414
R2642 VDD1.n169 VDD1.n107 1.16414
R2643 VDD1.n179 VDD1.n103 1.16414
R2644 VDD1.n81 VDD1.n8 0.388379
R2645 VDD1.n78 VDD1.n10 0.388379
R2646 VDD1.n34 VDD1.n32 0.388379
R2647 VDD1.n129 VDD1.n127 0.388379
R2648 VDD1.n175 VDD1.n174 0.388379
R2649 VDD1.n178 VDD1.n105 0.388379
R2650 VDD1.n95 VDD1.n1 0.155672
R2651 VDD1.n88 VDD1.n1 0.155672
R2652 VDD1.n88 VDD1.n87 0.155672
R2653 VDD1.n87 VDD1.n5 0.155672
R2654 VDD1.n80 VDD1.n5 0.155672
R2655 VDD1.n80 VDD1.n79 0.155672
R2656 VDD1.n79 VDD1.n9 0.155672
R2657 VDD1.n72 VDD1.n9 0.155672
R2658 VDD1.n72 VDD1.n71 0.155672
R2659 VDD1.n71 VDD1.n15 0.155672
R2660 VDD1.n64 VDD1.n15 0.155672
R2661 VDD1.n64 VDD1.n63 0.155672
R2662 VDD1.n63 VDD1.n19 0.155672
R2663 VDD1.n56 VDD1.n19 0.155672
R2664 VDD1.n56 VDD1.n55 0.155672
R2665 VDD1.n55 VDD1.n23 0.155672
R2666 VDD1.n48 VDD1.n23 0.155672
R2667 VDD1.n48 VDD1.n47 0.155672
R2668 VDD1.n47 VDD1.n27 0.155672
R2669 VDD1.n40 VDD1.n27 0.155672
R2670 VDD1.n40 VDD1.n39 0.155672
R2671 VDD1.n39 VDD1.n31 0.155672
R2672 VDD1.n134 VDD1.n126 0.155672
R2673 VDD1.n135 VDD1.n134 0.155672
R2674 VDD1.n135 VDD1.n122 0.155672
R2675 VDD1.n142 VDD1.n122 0.155672
R2676 VDD1.n143 VDD1.n142 0.155672
R2677 VDD1.n143 VDD1.n118 0.155672
R2678 VDD1.n150 VDD1.n118 0.155672
R2679 VDD1.n151 VDD1.n150 0.155672
R2680 VDD1.n151 VDD1.n114 0.155672
R2681 VDD1.n158 VDD1.n114 0.155672
R2682 VDD1.n159 VDD1.n158 0.155672
R2683 VDD1.n159 VDD1.n110 0.155672
R2684 VDD1.n166 VDD1.n110 0.155672
R2685 VDD1.n167 VDD1.n166 0.155672
R2686 VDD1.n167 VDD1.n106 0.155672
R2687 VDD1.n176 VDD1.n106 0.155672
R2688 VDD1.n177 VDD1.n176 0.155672
R2689 VDD1.n177 VDD1.n102 0.155672
R2690 VDD1.n184 VDD1.n102 0.155672
R2691 VDD1.n185 VDD1.n184 0.155672
R2692 VDD1.n185 VDD1.n98 0.155672
R2693 VDD1.n192 VDD1.n98 0.155672
C0 VDD1 VTAIL 6.53565f
C1 VP VDD2 0.339786f
C2 VDD2 VN 3.98049f
C3 VDD1 VDD2 0.693334f
C4 VDD2 VTAIL 6.58621f
C5 VP VN 6.55257f
C6 VP VDD1 4.16871f
C7 VDD1 VN 0.148191f
C8 VP VTAIL 3.42431f
C9 VN VTAIL 3.40996f
C10 VDD2 B 5.475072f
C11 VDD1 B 8.63856f
C12 VTAIL B 9.661626f
C13 VN B 12.2124f
C14 VP B 6.965181f
C15 VDD1.n0 B 0.027805f
C16 VDD1.n1 B 0.02007f
C17 VDD1.n2 B 0.010785f
C18 VDD1.n3 B 0.025492f
C19 VDD1.n4 B 0.011419f
C20 VDD1.n5 B 0.02007f
C21 VDD1.n6 B 0.010785f
C22 VDD1.n7 B 0.025492f
C23 VDD1.n8 B 0.011102f
C24 VDD1.n9 B 0.02007f
C25 VDD1.n10 B 0.011102f
C26 VDD1.n11 B 0.010785f
C27 VDD1.n12 B 0.025492f
C28 VDD1.n13 B 0.025492f
C29 VDD1.n14 B 0.011419f
C30 VDD1.n15 B 0.02007f
C31 VDD1.n16 B 0.010785f
C32 VDD1.n17 B 0.025492f
C33 VDD1.n18 B 0.011419f
C34 VDD1.n19 B 0.02007f
C35 VDD1.n20 B 0.010785f
C36 VDD1.n21 B 0.025492f
C37 VDD1.n22 B 0.011419f
C38 VDD1.n23 B 0.02007f
C39 VDD1.n24 B 0.010785f
C40 VDD1.n25 B 0.025492f
C41 VDD1.n26 B 0.011419f
C42 VDD1.n27 B 0.02007f
C43 VDD1.n28 B 0.010785f
C44 VDD1.n29 B 0.025492f
C45 VDD1.n30 B 0.011419f
C46 VDD1.n31 B 1.53853f
C47 VDD1.n32 B 0.010785f
C48 VDD1.t0 B 0.042207f
C49 VDD1.n33 B 0.143635f
C50 VDD1.n34 B 0.015059f
C51 VDD1.n35 B 0.019119f
C52 VDD1.n36 B 0.025492f
C53 VDD1.n37 B 0.011419f
C54 VDD1.n38 B 0.010785f
C55 VDD1.n39 B 0.02007f
C56 VDD1.n40 B 0.02007f
C57 VDD1.n41 B 0.010785f
C58 VDD1.n42 B 0.011419f
C59 VDD1.n43 B 0.025492f
C60 VDD1.n44 B 0.025492f
C61 VDD1.n45 B 0.011419f
C62 VDD1.n46 B 0.010785f
C63 VDD1.n47 B 0.02007f
C64 VDD1.n48 B 0.02007f
C65 VDD1.n49 B 0.010785f
C66 VDD1.n50 B 0.011419f
C67 VDD1.n51 B 0.025492f
C68 VDD1.n52 B 0.025492f
C69 VDD1.n53 B 0.011419f
C70 VDD1.n54 B 0.010785f
C71 VDD1.n55 B 0.02007f
C72 VDD1.n56 B 0.02007f
C73 VDD1.n57 B 0.010785f
C74 VDD1.n58 B 0.011419f
C75 VDD1.n59 B 0.025492f
C76 VDD1.n60 B 0.025492f
C77 VDD1.n61 B 0.011419f
C78 VDD1.n62 B 0.010785f
C79 VDD1.n63 B 0.02007f
C80 VDD1.n64 B 0.02007f
C81 VDD1.n65 B 0.010785f
C82 VDD1.n66 B 0.011419f
C83 VDD1.n67 B 0.025492f
C84 VDD1.n68 B 0.025492f
C85 VDD1.n69 B 0.011419f
C86 VDD1.n70 B 0.010785f
C87 VDD1.n71 B 0.02007f
C88 VDD1.n72 B 0.02007f
C89 VDD1.n73 B 0.010785f
C90 VDD1.n74 B 0.011419f
C91 VDD1.n75 B 0.025492f
C92 VDD1.n76 B 0.025492f
C93 VDD1.n77 B 0.011419f
C94 VDD1.n78 B 0.010785f
C95 VDD1.n79 B 0.02007f
C96 VDD1.n80 B 0.02007f
C97 VDD1.n81 B 0.010785f
C98 VDD1.n82 B 0.011419f
C99 VDD1.n83 B 0.025492f
C100 VDD1.n84 B 0.025492f
C101 VDD1.n85 B 0.011419f
C102 VDD1.n86 B 0.010785f
C103 VDD1.n87 B 0.02007f
C104 VDD1.n88 B 0.02007f
C105 VDD1.n89 B 0.010785f
C106 VDD1.n90 B 0.011419f
C107 VDD1.n91 B 0.025492f
C108 VDD1.n92 B 0.054467f
C109 VDD1.n93 B 0.011419f
C110 VDD1.n94 B 0.010785f
C111 VDD1.n95 B 0.046666f
C112 VDD1.n96 B 0.045507f
C113 VDD1.n97 B 0.027805f
C114 VDD1.n98 B 0.02007f
C115 VDD1.n99 B 0.010785f
C116 VDD1.n100 B 0.025492f
C117 VDD1.n101 B 0.011419f
C118 VDD1.n102 B 0.02007f
C119 VDD1.n103 B 0.010785f
C120 VDD1.n104 B 0.025492f
C121 VDD1.n105 B 0.011102f
C122 VDD1.n106 B 0.02007f
C123 VDD1.n107 B 0.011419f
C124 VDD1.n108 B 0.025492f
C125 VDD1.n109 B 0.011419f
C126 VDD1.n110 B 0.02007f
C127 VDD1.n111 B 0.010785f
C128 VDD1.n112 B 0.025492f
C129 VDD1.n113 B 0.011419f
C130 VDD1.n114 B 0.02007f
C131 VDD1.n115 B 0.010785f
C132 VDD1.n116 B 0.025492f
C133 VDD1.n117 B 0.011419f
C134 VDD1.n118 B 0.02007f
C135 VDD1.n119 B 0.010785f
C136 VDD1.n120 B 0.025492f
C137 VDD1.n121 B 0.011419f
C138 VDD1.n122 B 0.02007f
C139 VDD1.n123 B 0.010785f
C140 VDD1.n124 B 0.025492f
C141 VDD1.n125 B 0.011419f
C142 VDD1.n126 B 1.53853f
C143 VDD1.n127 B 0.010785f
C144 VDD1.t1 B 0.042207f
C145 VDD1.n128 B 0.143635f
C146 VDD1.n129 B 0.015059f
C147 VDD1.n130 B 0.019119f
C148 VDD1.n131 B 0.025492f
C149 VDD1.n132 B 0.011419f
C150 VDD1.n133 B 0.010785f
C151 VDD1.n134 B 0.02007f
C152 VDD1.n135 B 0.02007f
C153 VDD1.n136 B 0.010785f
C154 VDD1.n137 B 0.011419f
C155 VDD1.n138 B 0.025492f
C156 VDD1.n139 B 0.025492f
C157 VDD1.n140 B 0.011419f
C158 VDD1.n141 B 0.010785f
C159 VDD1.n142 B 0.02007f
C160 VDD1.n143 B 0.02007f
C161 VDD1.n144 B 0.010785f
C162 VDD1.n145 B 0.011419f
C163 VDD1.n146 B 0.025492f
C164 VDD1.n147 B 0.025492f
C165 VDD1.n148 B 0.011419f
C166 VDD1.n149 B 0.010785f
C167 VDD1.n150 B 0.02007f
C168 VDD1.n151 B 0.02007f
C169 VDD1.n152 B 0.010785f
C170 VDD1.n153 B 0.011419f
C171 VDD1.n154 B 0.025492f
C172 VDD1.n155 B 0.025492f
C173 VDD1.n156 B 0.011419f
C174 VDD1.n157 B 0.010785f
C175 VDD1.n158 B 0.02007f
C176 VDD1.n159 B 0.02007f
C177 VDD1.n160 B 0.010785f
C178 VDD1.n161 B 0.011419f
C179 VDD1.n162 B 0.025492f
C180 VDD1.n163 B 0.025492f
C181 VDD1.n164 B 0.011419f
C182 VDD1.n165 B 0.010785f
C183 VDD1.n166 B 0.02007f
C184 VDD1.n167 B 0.02007f
C185 VDD1.n168 B 0.010785f
C186 VDD1.n169 B 0.010785f
C187 VDD1.n170 B 0.011419f
C188 VDD1.n171 B 0.025492f
C189 VDD1.n172 B 0.025492f
C190 VDD1.n173 B 0.025492f
C191 VDD1.n174 B 0.011102f
C192 VDD1.n175 B 0.010785f
C193 VDD1.n176 B 0.02007f
C194 VDD1.n177 B 0.02007f
C195 VDD1.n178 B 0.010785f
C196 VDD1.n179 B 0.011419f
C197 VDD1.n180 B 0.025492f
C198 VDD1.n181 B 0.025492f
C199 VDD1.n182 B 0.011419f
C200 VDD1.n183 B 0.010785f
C201 VDD1.n184 B 0.02007f
C202 VDD1.n185 B 0.02007f
C203 VDD1.n186 B 0.010785f
C204 VDD1.n187 B 0.011419f
C205 VDD1.n188 B 0.025492f
C206 VDD1.n189 B 0.054467f
C207 VDD1.n190 B 0.011419f
C208 VDD1.n191 B 0.010785f
C209 VDD1.n192 B 0.046666f
C210 VDD1.n193 B 0.805883f
C211 VP.t0 B 4.17784f
C212 VP.t1 B 4.76553f
C213 VP.n0 B 5.17761f
C214 VDD2.n0 B 0.027737f
C215 VDD2.n1 B 0.020022f
C216 VDD2.n2 B 0.010759f
C217 VDD2.n3 B 0.02543f
C218 VDD2.n4 B 0.011392f
C219 VDD2.n5 B 0.020022f
C220 VDD2.n6 B 0.010759f
C221 VDD2.n7 B 0.02543f
C222 VDD2.n8 B 0.011075f
C223 VDD2.n9 B 0.020022f
C224 VDD2.n10 B 0.011392f
C225 VDD2.n11 B 0.02543f
C226 VDD2.n12 B 0.011392f
C227 VDD2.n13 B 0.020022f
C228 VDD2.n14 B 0.010759f
C229 VDD2.n15 B 0.02543f
C230 VDD2.n16 B 0.011392f
C231 VDD2.n17 B 0.020022f
C232 VDD2.n18 B 0.010759f
C233 VDD2.n19 B 0.02543f
C234 VDD2.n20 B 0.011392f
C235 VDD2.n21 B 0.020022f
C236 VDD2.n22 B 0.010759f
C237 VDD2.n23 B 0.02543f
C238 VDD2.n24 B 0.011392f
C239 VDD2.n25 B 0.020022f
C240 VDD2.n26 B 0.010759f
C241 VDD2.n27 B 0.02543f
C242 VDD2.n28 B 0.011392f
C243 VDD2.n29 B 1.53478f
C244 VDD2.n30 B 0.010759f
C245 VDD2.t1 B 0.042104f
C246 VDD2.n31 B 0.143285f
C247 VDD2.n32 B 0.015022f
C248 VDD2.n33 B 0.019072f
C249 VDD2.n34 B 0.02543f
C250 VDD2.n35 B 0.011392f
C251 VDD2.n36 B 0.010759f
C252 VDD2.n37 B 0.020022f
C253 VDD2.n38 B 0.020022f
C254 VDD2.n39 B 0.010759f
C255 VDD2.n40 B 0.011392f
C256 VDD2.n41 B 0.02543f
C257 VDD2.n42 B 0.02543f
C258 VDD2.n43 B 0.011392f
C259 VDD2.n44 B 0.010759f
C260 VDD2.n45 B 0.020022f
C261 VDD2.n46 B 0.020022f
C262 VDD2.n47 B 0.010759f
C263 VDD2.n48 B 0.011392f
C264 VDD2.n49 B 0.02543f
C265 VDD2.n50 B 0.02543f
C266 VDD2.n51 B 0.011392f
C267 VDD2.n52 B 0.010759f
C268 VDD2.n53 B 0.020022f
C269 VDD2.n54 B 0.020022f
C270 VDD2.n55 B 0.010759f
C271 VDD2.n56 B 0.011392f
C272 VDD2.n57 B 0.02543f
C273 VDD2.n58 B 0.02543f
C274 VDD2.n59 B 0.011392f
C275 VDD2.n60 B 0.010759f
C276 VDD2.n61 B 0.020022f
C277 VDD2.n62 B 0.020022f
C278 VDD2.n63 B 0.010759f
C279 VDD2.n64 B 0.011392f
C280 VDD2.n65 B 0.02543f
C281 VDD2.n66 B 0.02543f
C282 VDD2.n67 B 0.011392f
C283 VDD2.n68 B 0.010759f
C284 VDD2.n69 B 0.020022f
C285 VDD2.n70 B 0.020022f
C286 VDD2.n71 B 0.010759f
C287 VDD2.n72 B 0.010759f
C288 VDD2.n73 B 0.011392f
C289 VDD2.n74 B 0.02543f
C290 VDD2.n75 B 0.02543f
C291 VDD2.n76 B 0.02543f
C292 VDD2.n77 B 0.011075f
C293 VDD2.n78 B 0.010759f
C294 VDD2.n79 B 0.020022f
C295 VDD2.n80 B 0.020022f
C296 VDD2.n81 B 0.010759f
C297 VDD2.n82 B 0.011392f
C298 VDD2.n83 B 0.02543f
C299 VDD2.n84 B 0.02543f
C300 VDD2.n85 B 0.011392f
C301 VDD2.n86 B 0.010759f
C302 VDD2.n87 B 0.020022f
C303 VDD2.n88 B 0.020022f
C304 VDD2.n89 B 0.010759f
C305 VDD2.n90 B 0.011392f
C306 VDD2.n91 B 0.02543f
C307 VDD2.n92 B 0.054334f
C308 VDD2.n93 B 0.011392f
C309 VDD2.n94 B 0.010759f
C310 VDD2.n95 B 0.046553f
C311 VDD2.n96 B 0.760067f
C312 VDD2.n97 B 0.027737f
C313 VDD2.n98 B 0.020022f
C314 VDD2.n99 B 0.010759f
C315 VDD2.n100 B 0.02543f
C316 VDD2.n101 B 0.011392f
C317 VDD2.n102 B 0.020022f
C318 VDD2.n103 B 0.010759f
C319 VDD2.n104 B 0.02543f
C320 VDD2.n105 B 0.011075f
C321 VDD2.n106 B 0.020022f
C322 VDD2.n107 B 0.011075f
C323 VDD2.n108 B 0.010759f
C324 VDD2.n109 B 0.02543f
C325 VDD2.n110 B 0.02543f
C326 VDD2.n111 B 0.011392f
C327 VDD2.n112 B 0.020022f
C328 VDD2.n113 B 0.010759f
C329 VDD2.n114 B 0.02543f
C330 VDD2.n115 B 0.011392f
C331 VDD2.n116 B 0.020022f
C332 VDD2.n117 B 0.010759f
C333 VDD2.n118 B 0.02543f
C334 VDD2.n119 B 0.011392f
C335 VDD2.n120 B 0.020022f
C336 VDD2.n121 B 0.010759f
C337 VDD2.n122 B 0.02543f
C338 VDD2.n123 B 0.011392f
C339 VDD2.n124 B 0.020022f
C340 VDD2.n125 B 0.010759f
C341 VDD2.n126 B 0.02543f
C342 VDD2.n127 B 0.011392f
C343 VDD2.n128 B 1.53478f
C344 VDD2.n129 B 0.010759f
C345 VDD2.t0 B 0.042104f
C346 VDD2.n130 B 0.143285f
C347 VDD2.n131 B 0.015022f
C348 VDD2.n132 B 0.019072f
C349 VDD2.n133 B 0.02543f
C350 VDD2.n134 B 0.011392f
C351 VDD2.n135 B 0.010759f
C352 VDD2.n136 B 0.020022f
C353 VDD2.n137 B 0.020022f
C354 VDD2.n138 B 0.010759f
C355 VDD2.n139 B 0.011392f
C356 VDD2.n140 B 0.02543f
C357 VDD2.n141 B 0.02543f
C358 VDD2.n142 B 0.011392f
C359 VDD2.n143 B 0.010759f
C360 VDD2.n144 B 0.020022f
C361 VDD2.n145 B 0.020022f
C362 VDD2.n146 B 0.010759f
C363 VDD2.n147 B 0.011392f
C364 VDD2.n148 B 0.02543f
C365 VDD2.n149 B 0.02543f
C366 VDD2.n150 B 0.011392f
C367 VDD2.n151 B 0.010759f
C368 VDD2.n152 B 0.020022f
C369 VDD2.n153 B 0.020022f
C370 VDD2.n154 B 0.010759f
C371 VDD2.n155 B 0.011392f
C372 VDD2.n156 B 0.02543f
C373 VDD2.n157 B 0.02543f
C374 VDD2.n158 B 0.011392f
C375 VDD2.n159 B 0.010759f
C376 VDD2.n160 B 0.020022f
C377 VDD2.n161 B 0.020022f
C378 VDD2.n162 B 0.010759f
C379 VDD2.n163 B 0.011392f
C380 VDD2.n164 B 0.02543f
C381 VDD2.n165 B 0.02543f
C382 VDD2.n166 B 0.011392f
C383 VDD2.n167 B 0.010759f
C384 VDD2.n168 B 0.020022f
C385 VDD2.n169 B 0.020022f
C386 VDD2.n170 B 0.010759f
C387 VDD2.n171 B 0.011392f
C388 VDD2.n172 B 0.02543f
C389 VDD2.n173 B 0.02543f
C390 VDD2.n174 B 0.011392f
C391 VDD2.n175 B 0.010759f
C392 VDD2.n176 B 0.020022f
C393 VDD2.n177 B 0.020022f
C394 VDD2.n178 B 0.010759f
C395 VDD2.n179 B 0.011392f
C396 VDD2.n180 B 0.02543f
C397 VDD2.n181 B 0.02543f
C398 VDD2.n182 B 0.011392f
C399 VDD2.n183 B 0.010759f
C400 VDD2.n184 B 0.020022f
C401 VDD2.n185 B 0.020022f
C402 VDD2.n186 B 0.010759f
C403 VDD2.n187 B 0.011392f
C404 VDD2.n188 B 0.02543f
C405 VDD2.n189 B 0.054334f
C406 VDD2.n190 B 0.011392f
C407 VDD2.n191 B 0.010759f
C408 VDD2.n192 B 0.046553f
C409 VDD2.n193 B 0.044159f
C410 VDD2.n194 B 2.91974f
C411 VTAIL.n0 B 0.027384f
C412 VTAIL.n1 B 0.019767f
C413 VTAIL.n2 B 0.010622f
C414 VTAIL.n3 B 0.025107f
C415 VTAIL.n4 B 0.011247f
C416 VTAIL.n5 B 0.019767f
C417 VTAIL.n6 B 0.010622f
C418 VTAIL.n7 B 0.025107f
C419 VTAIL.n8 B 0.010934f
C420 VTAIL.n9 B 0.019767f
C421 VTAIL.n10 B 0.011247f
C422 VTAIL.n11 B 0.025107f
C423 VTAIL.n12 B 0.011247f
C424 VTAIL.n13 B 0.019767f
C425 VTAIL.n14 B 0.010622f
C426 VTAIL.n15 B 0.025107f
C427 VTAIL.n16 B 0.011247f
C428 VTAIL.n17 B 0.019767f
C429 VTAIL.n18 B 0.010622f
C430 VTAIL.n19 B 0.025107f
C431 VTAIL.n20 B 0.011247f
C432 VTAIL.n21 B 0.019767f
C433 VTAIL.n22 B 0.010622f
C434 VTAIL.n23 B 0.025107f
C435 VTAIL.n24 B 0.011247f
C436 VTAIL.n25 B 0.019767f
C437 VTAIL.n26 B 0.010622f
C438 VTAIL.n27 B 0.025107f
C439 VTAIL.n28 B 0.011247f
C440 VTAIL.n29 B 1.51528f
C441 VTAIL.n30 B 0.010622f
C442 VTAIL.t3 B 0.041569f
C443 VTAIL.n31 B 0.141465f
C444 VTAIL.n32 B 0.014831f
C445 VTAIL.n33 B 0.01883f
C446 VTAIL.n34 B 0.025107f
C447 VTAIL.n35 B 0.011247f
C448 VTAIL.n36 B 0.010622f
C449 VTAIL.n37 B 0.019767f
C450 VTAIL.n38 B 0.019767f
C451 VTAIL.n39 B 0.010622f
C452 VTAIL.n40 B 0.011247f
C453 VTAIL.n41 B 0.025107f
C454 VTAIL.n42 B 0.025107f
C455 VTAIL.n43 B 0.011247f
C456 VTAIL.n44 B 0.010622f
C457 VTAIL.n45 B 0.019767f
C458 VTAIL.n46 B 0.019767f
C459 VTAIL.n47 B 0.010622f
C460 VTAIL.n48 B 0.011247f
C461 VTAIL.n49 B 0.025107f
C462 VTAIL.n50 B 0.025107f
C463 VTAIL.n51 B 0.011247f
C464 VTAIL.n52 B 0.010622f
C465 VTAIL.n53 B 0.019767f
C466 VTAIL.n54 B 0.019767f
C467 VTAIL.n55 B 0.010622f
C468 VTAIL.n56 B 0.011247f
C469 VTAIL.n57 B 0.025107f
C470 VTAIL.n58 B 0.025107f
C471 VTAIL.n59 B 0.011247f
C472 VTAIL.n60 B 0.010622f
C473 VTAIL.n61 B 0.019767f
C474 VTAIL.n62 B 0.019767f
C475 VTAIL.n63 B 0.010622f
C476 VTAIL.n64 B 0.011247f
C477 VTAIL.n65 B 0.025107f
C478 VTAIL.n66 B 0.025107f
C479 VTAIL.n67 B 0.011247f
C480 VTAIL.n68 B 0.010622f
C481 VTAIL.n69 B 0.019767f
C482 VTAIL.n70 B 0.019767f
C483 VTAIL.n71 B 0.010622f
C484 VTAIL.n72 B 0.010622f
C485 VTAIL.n73 B 0.011247f
C486 VTAIL.n74 B 0.025107f
C487 VTAIL.n75 B 0.025107f
C488 VTAIL.n76 B 0.025107f
C489 VTAIL.n77 B 0.010934f
C490 VTAIL.n78 B 0.010622f
C491 VTAIL.n79 B 0.019767f
C492 VTAIL.n80 B 0.019767f
C493 VTAIL.n81 B 0.010622f
C494 VTAIL.n82 B 0.011247f
C495 VTAIL.n83 B 0.025107f
C496 VTAIL.n84 B 0.025107f
C497 VTAIL.n85 B 0.011247f
C498 VTAIL.n86 B 0.010622f
C499 VTAIL.n87 B 0.019767f
C500 VTAIL.n88 B 0.019767f
C501 VTAIL.n89 B 0.010622f
C502 VTAIL.n90 B 0.011247f
C503 VTAIL.n91 B 0.025107f
C504 VTAIL.n92 B 0.053644f
C505 VTAIL.n93 B 0.011247f
C506 VTAIL.n94 B 0.010622f
C507 VTAIL.n95 B 0.045961f
C508 VTAIL.n96 B 0.029951f
C509 VTAIL.n97 B 1.66225f
C510 VTAIL.n98 B 0.027384f
C511 VTAIL.n99 B 0.019767f
C512 VTAIL.n100 B 0.010622f
C513 VTAIL.n101 B 0.025107f
C514 VTAIL.n102 B 0.011247f
C515 VTAIL.n103 B 0.019767f
C516 VTAIL.n104 B 0.010622f
C517 VTAIL.n105 B 0.025107f
C518 VTAIL.n106 B 0.010934f
C519 VTAIL.n107 B 0.019767f
C520 VTAIL.n108 B 0.010934f
C521 VTAIL.n109 B 0.010622f
C522 VTAIL.n110 B 0.025107f
C523 VTAIL.n111 B 0.025107f
C524 VTAIL.n112 B 0.011247f
C525 VTAIL.n113 B 0.019767f
C526 VTAIL.n114 B 0.010622f
C527 VTAIL.n115 B 0.025107f
C528 VTAIL.n116 B 0.011247f
C529 VTAIL.n117 B 0.019767f
C530 VTAIL.n118 B 0.010622f
C531 VTAIL.n119 B 0.025107f
C532 VTAIL.n120 B 0.011247f
C533 VTAIL.n121 B 0.019767f
C534 VTAIL.n122 B 0.010622f
C535 VTAIL.n123 B 0.025107f
C536 VTAIL.n124 B 0.011247f
C537 VTAIL.n125 B 0.019767f
C538 VTAIL.n126 B 0.010622f
C539 VTAIL.n127 B 0.025107f
C540 VTAIL.n128 B 0.011247f
C541 VTAIL.n129 B 1.51528f
C542 VTAIL.n130 B 0.010622f
C543 VTAIL.t1 B 0.041569f
C544 VTAIL.n131 B 0.141465f
C545 VTAIL.n132 B 0.014831f
C546 VTAIL.n133 B 0.01883f
C547 VTAIL.n134 B 0.025107f
C548 VTAIL.n135 B 0.011247f
C549 VTAIL.n136 B 0.010622f
C550 VTAIL.n137 B 0.019767f
C551 VTAIL.n138 B 0.019767f
C552 VTAIL.n139 B 0.010622f
C553 VTAIL.n140 B 0.011247f
C554 VTAIL.n141 B 0.025107f
C555 VTAIL.n142 B 0.025107f
C556 VTAIL.n143 B 0.011247f
C557 VTAIL.n144 B 0.010622f
C558 VTAIL.n145 B 0.019767f
C559 VTAIL.n146 B 0.019767f
C560 VTAIL.n147 B 0.010622f
C561 VTAIL.n148 B 0.011247f
C562 VTAIL.n149 B 0.025107f
C563 VTAIL.n150 B 0.025107f
C564 VTAIL.n151 B 0.011247f
C565 VTAIL.n152 B 0.010622f
C566 VTAIL.n153 B 0.019767f
C567 VTAIL.n154 B 0.019767f
C568 VTAIL.n155 B 0.010622f
C569 VTAIL.n156 B 0.011247f
C570 VTAIL.n157 B 0.025107f
C571 VTAIL.n158 B 0.025107f
C572 VTAIL.n159 B 0.011247f
C573 VTAIL.n160 B 0.010622f
C574 VTAIL.n161 B 0.019767f
C575 VTAIL.n162 B 0.019767f
C576 VTAIL.n163 B 0.010622f
C577 VTAIL.n164 B 0.011247f
C578 VTAIL.n165 B 0.025107f
C579 VTAIL.n166 B 0.025107f
C580 VTAIL.n167 B 0.011247f
C581 VTAIL.n168 B 0.010622f
C582 VTAIL.n169 B 0.019767f
C583 VTAIL.n170 B 0.019767f
C584 VTAIL.n171 B 0.010622f
C585 VTAIL.n172 B 0.011247f
C586 VTAIL.n173 B 0.025107f
C587 VTAIL.n174 B 0.025107f
C588 VTAIL.n175 B 0.011247f
C589 VTAIL.n176 B 0.010622f
C590 VTAIL.n177 B 0.019767f
C591 VTAIL.n178 B 0.019767f
C592 VTAIL.n179 B 0.010622f
C593 VTAIL.n180 B 0.011247f
C594 VTAIL.n181 B 0.025107f
C595 VTAIL.n182 B 0.025107f
C596 VTAIL.n183 B 0.011247f
C597 VTAIL.n184 B 0.010622f
C598 VTAIL.n185 B 0.019767f
C599 VTAIL.n186 B 0.019767f
C600 VTAIL.n187 B 0.010622f
C601 VTAIL.n188 B 0.011247f
C602 VTAIL.n189 B 0.025107f
C603 VTAIL.n190 B 0.053644f
C604 VTAIL.n191 B 0.011247f
C605 VTAIL.n192 B 0.010622f
C606 VTAIL.n193 B 0.045961f
C607 VTAIL.n194 B 0.029951f
C608 VTAIL.n195 B 1.70083f
C609 VTAIL.n196 B 0.027384f
C610 VTAIL.n197 B 0.019767f
C611 VTAIL.n198 B 0.010622f
C612 VTAIL.n199 B 0.025107f
C613 VTAIL.n200 B 0.011247f
C614 VTAIL.n201 B 0.019767f
C615 VTAIL.n202 B 0.010622f
C616 VTAIL.n203 B 0.025107f
C617 VTAIL.n204 B 0.010934f
C618 VTAIL.n205 B 0.019767f
C619 VTAIL.n206 B 0.010934f
C620 VTAIL.n207 B 0.010622f
C621 VTAIL.n208 B 0.025107f
C622 VTAIL.n209 B 0.025107f
C623 VTAIL.n210 B 0.011247f
C624 VTAIL.n211 B 0.019767f
C625 VTAIL.n212 B 0.010622f
C626 VTAIL.n213 B 0.025107f
C627 VTAIL.n214 B 0.011247f
C628 VTAIL.n215 B 0.019767f
C629 VTAIL.n216 B 0.010622f
C630 VTAIL.n217 B 0.025107f
C631 VTAIL.n218 B 0.011247f
C632 VTAIL.n219 B 0.019767f
C633 VTAIL.n220 B 0.010622f
C634 VTAIL.n221 B 0.025107f
C635 VTAIL.n222 B 0.011247f
C636 VTAIL.n223 B 0.019767f
C637 VTAIL.n224 B 0.010622f
C638 VTAIL.n225 B 0.025107f
C639 VTAIL.n226 B 0.011247f
C640 VTAIL.n227 B 1.51528f
C641 VTAIL.n228 B 0.010622f
C642 VTAIL.t2 B 0.041569f
C643 VTAIL.n229 B 0.141465f
C644 VTAIL.n230 B 0.014831f
C645 VTAIL.n231 B 0.01883f
C646 VTAIL.n232 B 0.025107f
C647 VTAIL.n233 B 0.011247f
C648 VTAIL.n234 B 0.010622f
C649 VTAIL.n235 B 0.019767f
C650 VTAIL.n236 B 0.019767f
C651 VTAIL.n237 B 0.010622f
C652 VTAIL.n238 B 0.011247f
C653 VTAIL.n239 B 0.025107f
C654 VTAIL.n240 B 0.025107f
C655 VTAIL.n241 B 0.011247f
C656 VTAIL.n242 B 0.010622f
C657 VTAIL.n243 B 0.019767f
C658 VTAIL.n244 B 0.019767f
C659 VTAIL.n245 B 0.010622f
C660 VTAIL.n246 B 0.011247f
C661 VTAIL.n247 B 0.025107f
C662 VTAIL.n248 B 0.025107f
C663 VTAIL.n249 B 0.011247f
C664 VTAIL.n250 B 0.010622f
C665 VTAIL.n251 B 0.019767f
C666 VTAIL.n252 B 0.019767f
C667 VTAIL.n253 B 0.010622f
C668 VTAIL.n254 B 0.011247f
C669 VTAIL.n255 B 0.025107f
C670 VTAIL.n256 B 0.025107f
C671 VTAIL.n257 B 0.011247f
C672 VTAIL.n258 B 0.010622f
C673 VTAIL.n259 B 0.019767f
C674 VTAIL.n260 B 0.019767f
C675 VTAIL.n261 B 0.010622f
C676 VTAIL.n262 B 0.011247f
C677 VTAIL.n263 B 0.025107f
C678 VTAIL.n264 B 0.025107f
C679 VTAIL.n265 B 0.011247f
C680 VTAIL.n266 B 0.010622f
C681 VTAIL.n267 B 0.019767f
C682 VTAIL.n268 B 0.019767f
C683 VTAIL.n269 B 0.010622f
C684 VTAIL.n270 B 0.011247f
C685 VTAIL.n271 B 0.025107f
C686 VTAIL.n272 B 0.025107f
C687 VTAIL.n273 B 0.011247f
C688 VTAIL.n274 B 0.010622f
C689 VTAIL.n275 B 0.019767f
C690 VTAIL.n276 B 0.019767f
C691 VTAIL.n277 B 0.010622f
C692 VTAIL.n278 B 0.011247f
C693 VTAIL.n279 B 0.025107f
C694 VTAIL.n280 B 0.025107f
C695 VTAIL.n281 B 0.011247f
C696 VTAIL.n282 B 0.010622f
C697 VTAIL.n283 B 0.019767f
C698 VTAIL.n284 B 0.019767f
C699 VTAIL.n285 B 0.010622f
C700 VTAIL.n286 B 0.011247f
C701 VTAIL.n287 B 0.025107f
C702 VTAIL.n288 B 0.053644f
C703 VTAIL.n289 B 0.011247f
C704 VTAIL.n290 B 0.010622f
C705 VTAIL.n291 B 0.045961f
C706 VTAIL.n292 B 0.029951f
C707 VTAIL.n293 B 1.53171f
C708 VTAIL.n294 B 0.027384f
C709 VTAIL.n295 B 0.019767f
C710 VTAIL.n296 B 0.010622f
C711 VTAIL.n297 B 0.025107f
C712 VTAIL.n298 B 0.011247f
C713 VTAIL.n299 B 0.019767f
C714 VTAIL.n300 B 0.010622f
C715 VTAIL.n301 B 0.025107f
C716 VTAIL.n302 B 0.010934f
C717 VTAIL.n303 B 0.019767f
C718 VTAIL.n304 B 0.011247f
C719 VTAIL.n305 B 0.025107f
C720 VTAIL.n306 B 0.011247f
C721 VTAIL.n307 B 0.019767f
C722 VTAIL.n308 B 0.010622f
C723 VTAIL.n309 B 0.025107f
C724 VTAIL.n310 B 0.011247f
C725 VTAIL.n311 B 0.019767f
C726 VTAIL.n312 B 0.010622f
C727 VTAIL.n313 B 0.025107f
C728 VTAIL.n314 B 0.011247f
C729 VTAIL.n315 B 0.019767f
C730 VTAIL.n316 B 0.010622f
C731 VTAIL.n317 B 0.025107f
C732 VTAIL.n318 B 0.011247f
C733 VTAIL.n319 B 0.019767f
C734 VTAIL.n320 B 0.010622f
C735 VTAIL.n321 B 0.025107f
C736 VTAIL.n322 B 0.011247f
C737 VTAIL.n323 B 1.51528f
C738 VTAIL.n324 B 0.010622f
C739 VTAIL.t0 B 0.041569f
C740 VTAIL.n325 B 0.141465f
C741 VTAIL.n326 B 0.014831f
C742 VTAIL.n327 B 0.01883f
C743 VTAIL.n328 B 0.025107f
C744 VTAIL.n329 B 0.011247f
C745 VTAIL.n330 B 0.010622f
C746 VTAIL.n331 B 0.019767f
C747 VTAIL.n332 B 0.019767f
C748 VTAIL.n333 B 0.010622f
C749 VTAIL.n334 B 0.011247f
C750 VTAIL.n335 B 0.025107f
C751 VTAIL.n336 B 0.025107f
C752 VTAIL.n337 B 0.011247f
C753 VTAIL.n338 B 0.010622f
C754 VTAIL.n339 B 0.019767f
C755 VTAIL.n340 B 0.019767f
C756 VTAIL.n341 B 0.010622f
C757 VTAIL.n342 B 0.011247f
C758 VTAIL.n343 B 0.025107f
C759 VTAIL.n344 B 0.025107f
C760 VTAIL.n345 B 0.011247f
C761 VTAIL.n346 B 0.010622f
C762 VTAIL.n347 B 0.019767f
C763 VTAIL.n348 B 0.019767f
C764 VTAIL.n349 B 0.010622f
C765 VTAIL.n350 B 0.011247f
C766 VTAIL.n351 B 0.025107f
C767 VTAIL.n352 B 0.025107f
C768 VTAIL.n353 B 0.011247f
C769 VTAIL.n354 B 0.010622f
C770 VTAIL.n355 B 0.019767f
C771 VTAIL.n356 B 0.019767f
C772 VTAIL.n357 B 0.010622f
C773 VTAIL.n358 B 0.011247f
C774 VTAIL.n359 B 0.025107f
C775 VTAIL.n360 B 0.025107f
C776 VTAIL.n361 B 0.011247f
C777 VTAIL.n362 B 0.010622f
C778 VTAIL.n363 B 0.019767f
C779 VTAIL.n364 B 0.019767f
C780 VTAIL.n365 B 0.010622f
C781 VTAIL.n366 B 0.010622f
C782 VTAIL.n367 B 0.011247f
C783 VTAIL.n368 B 0.025107f
C784 VTAIL.n369 B 0.025107f
C785 VTAIL.n370 B 0.025107f
C786 VTAIL.n371 B 0.010934f
C787 VTAIL.n372 B 0.010622f
C788 VTAIL.n373 B 0.019767f
C789 VTAIL.n374 B 0.019767f
C790 VTAIL.n375 B 0.010622f
C791 VTAIL.n376 B 0.011247f
C792 VTAIL.n377 B 0.025107f
C793 VTAIL.n378 B 0.025107f
C794 VTAIL.n379 B 0.011247f
C795 VTAIL.n380 B 0.010622f
C796 VTAIL.n381 B 0.019767f
C797 VTAIL.n382 B 0.019767f
C798 VTAIL.n383 B 0.010622f
C799 VTAIL.n384 B 0.011247f
C800 VTAIL.n385 B 0.025107f
C801 VTAIL.n386 B 0.053644f
C802 VTAIL.n387 B 0.011247f
C803 VTAIL.n388 B 0.010622f
C804 VTAIL.n389 B 0.045961f
C805 VTAIL.n390 B 0.029951f
C806 VTAIL.n391 B 1.45579f
C807 VN.t0 B 4.11013f
C808 VN.t1 B 4.68624f
.ends

