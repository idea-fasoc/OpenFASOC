* NGSPICE file created from diff_pair_sample_1677.ext - technology: sky130A

.subckt diff_pair_sample_1677 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=0 ps=0 w=13.97 l=1.73
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=0 ps=0 w=13.97 l=1.73
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=0 ps=0 w=13.97 l=1.73
X3 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=5.4483 ps=28.72 w=13.97 l=1.73
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=5.4483 ps=28.72 w=13.97 l=1.73
X5 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=5.4483 ps=28.72 w=13.97 l=1.73
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=5.4483 ps=28.72 w=13.97 l=1.73
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4483 pd=28.72 as=0 ps=0 w=13.97 l=1.73
R0 B.n692 B.n691 585
R1 B.n301 B.n92 585
R2 B.n300 B.n299 585
R3 B.n298 B.n297 585
R4 B.n296 B.n295 585
R5 B.n294 B.n293 585
R6 B.n292 B.n291 585
R7 B.n290 B.n289 585
R8 B.n288 B.n287 585
R9 B.n286 B.n285 585
R10 B.n284 B.n283 585
R11 B.n282 B.n281 585
R12 B.n280 B.n279 585
R13 B.n278 B.n277 585
R14 B.n276 B.n275 585
R15 B.n274 B.n273 585
R16 B.n272 B.n271 585
R17 B.n270 B.n269 585
R18 B.n268 B.n267 585
R19 B.n266 B.n265 585
R20 B.n264 B.n263 585
R21 B.n262 B.n261 585
R22 B.n260 B.n259 585
R23 B.n258 B.n257 585
R24 B.n256 B.n255 585
R25 B.n254 B.n253 585
R26 B.n252 B.n251 585
R27 B.n250 B.n249 585
R28 B.n248 B.n247 585
R29 B.n246 B.n245 585
R30 B.n244 B.n243 585
R31 B.n242 B.n241 585
R32 B.n240 B.n239 585
R33 B.n238 B.n237 585
R34 B.n236 B.n235 585
R35 B.n234 B.n233 585
R36 B.n232 B.n231 585
R37 B.n230 B.n229 585
R38 B.n228 B.n227 585
R39 B.n226 B.n225 585
R40 B.n224 B.n223 585
R41 B.n222 B.n221 585
R42 B.n220 B.n219 585
R43 B.n218 B.n217 585
R44 B.n216 B.n215 585
R45 B.n214 B.n213 585
R46 B.n212 B.n211 585
R47 B.n209 B.n208 585
R48 B.n207 B.n206 585
R49 B.n205 B.n204 585
R50 B.n203 B.n202 585
R51 B.n201 B.n200 585
R52 B.n199 B.n198 585
R53 B.n197 B.n196 585
R54 B.n195 B.n194 585
R55 B.n193 B.n192 585
R56 B.n191 B.n190 585
R57 B.n188 B.n187 585
R58 B.n186 B.n185 585
R59 B.n184 B.n183 585
R60 B.n182 B.n181 585
R61 B.n180 B.n179 585
R62 B.n178 B.n177 585
R63 B.n176 B.n175 585
R64 B.n174 B.n173 585
R65 B.n172 B.n171 585
R66 B.n170 B.n169 585
R67 B.n168 B.n167 585
R68 B.n166 B.n165 585
R69 B.n164 B.n163 585
R70 B.n162 B.n161 585
R71 B.n160 B.n159 585
R72 B.n158 B.n157 585
R73 B.n156 B.n155 585
R74 B.n154 B.n153 585
R75 B.n152 B.n151 585
R76 B.n150 B.n149 585
R77 B.n148 B.n147 585
R78 B.n146 B.n145 585
R79 B.n144 B.n143 585
R80 B.n142 B.n141 585
R81 B.n140 B.n139 585
R82 B.n138 B.n137 585
R83 B.n136 B.n135 585
R84 B.n134 B.n133 585
R85 B.n132 B.n131 585
R86 B.n130 B.n129 585
R87 B.n128 B.n127 585
R88 B.n126 B.n125 585
R89 B.n124 B.n123 585
R90 B.n122 B.n121 585
R91 B.n120 B.n119 585
R92 B.n118 B.n117 585
R93 B.n116 B.n115 585
R94 B.n114 B.n113 585
R95 B.n112 B.n111 585
R96 B.n110 B.n109 585
R97 B.n108 B.n107 585
R98 B.n106 B.n105 585
R99 B.n104 B.n103 585
R100 B.n102 B.n101 585
R101 B.n100 B.n99 585
R102 B.n98 B.n97 585
R103 B.n39 B.n38 585
R104 B.n690 B.n40 585
R105 B.n695 B.n40 585
R106 B.n689 B.n688 585
R107 B.n688 B.n36 585
R108 B.n687 B.n35 585
R109 B.n701 B.n35 585
R110 B.n686 B.n34 585
R111 B.n702 B.n34 585
R112 B.n685 B.n33 585
R113 B.n703 B.n33 585
R114 B.n684 B.n683 585
R115 B.n683 B.n29 585
R116 B.n682 B.n28 585
R117 B.n709 B.n28 585
R118 B.n681 B.n27 585
R119 B.n710 B.n27 585
R120 B.n680 B.n26 585
R121 B.n711 B.n26 585
R122 B.n679 B.n678 585
R123 B.n678 B.n22 585
R124 B.n677 B.n21 585
R125 B.n717 B.n21 585
R126 B.n676 B.n20 585
R127 B.n718 B.n20 585
R128 B.n675 B.n19 585
R129 B.n719 B.n19 585
R130 B.n674 B.n673 585
R131 B.n673 B.n15 585
R132 B.n672 B.n14 585
R133 B.n725 B.n14 585
R134 B.n671 B.n13 585
R135 B.n726 B.n13 585
R136 B.n670 B.n12 585
R137 B.n727 B.n12 585
R138 B.n669 B.n668 585
R139 B.n668 B.n8 585
R140 B.n667 B.n7 585
R141 B.n733 B.n7 585
R142 B.n666 B.n6 585
R143 B.n734 B.n6 585
R144 B.n665 B.n5 585
R145 B.n735 B.n5 585
R146 B.n664 B.n663 585
R147 B.n663 B.n4 585
R148 B.n662 B.n302 585
R149 B.n662 B.n661 585
R150 B.n652 B.n303 585
R151 B.n304 B.n303 585
R152 B.n654 B.n653 585
R153 B.n655 B.n654 585
R154 B.n651 B.n308 585
R155 B.n312 B.n308 585
R156 B.n650 B.n649 585
R157 B.n649 B.n648 585
R158 B.n310 B.n309 585
R159 B.n311 B.n310 585
R160 B.n641 B.n640 585
R161 B.n642 B.n641 585
R162 B.n639 B.n317 585
R163 B.n317 B.n316 585
R164 B.n638 B.n637 585
R165 B.n637 B.n636 585
R166 B.n319 B.n318 585
R167 B.n320 B.n319 585
R168 B.n629 B.n628 585
R169 B.n630 B.n629 585
R170 B.n627 B.n325 585
R171 B.n325 B.n324 585
R172 B.n626 B.n625 585
R173 B.n625 B.n624 585
R174 B.n327 B.n326 585
R175 B.n328 B.n327 585
R176 B.n617 B.n616 585
R177 B.n618 B.n617 585
R178 B.n615 B.n333 585
R179 B.n333 B.n332 585
R180 B.n614 B.n613 585
R181 B.n613 B.n612 585
R182 B.n335 B.n334 585
R183 B.n336 B.n335 585
R184 B.n605 B.n604 585
R185 B.n606 B.n605 585
R186 B.n339 B.n338 585
R187 B.n400 B.n399 585
R188 B.n401 B.n397 585
R189 B.n397 B.n340 585
R190 B.n403 B.n402 585
R191 B.n405 B.n396 585
R192 B.n408 B.n407 585
R193 B.n409 B.n395 585
R194 B.n411 B.n410 585
R195 B.n413 B.n394 585
R196 B.n416 B.n415 585
R197 B.n417 B.n393 585
R198 B.n419 B.n418 585
R199 B.n421 B.n392 585
R200 B.n424 B.n423 585
R201 B.n425 B.n391 585
R202 B.n427 B.n426 585
R203 B.n429 B.n390 585
R204 B.n432 B.n431 585
R205 B.n433 B.n389 585
R206 B.n435 B.n434 585
R207 B.n437 B.n388 585
R208 B.n440 B.n439 585
R209 B.n441 B.n387 585
R210 B.n443 B.n442 585
R211 B.n445 B.n386 585
R212 B.n448 B.n447 585
R213 B.n449 B.n385 585
R214 B.n451 B.n450 585
R215 B.n453 B.n384 585
R216 B.n456 B.n455 585
R217 B.n457 B.n383 585
R218 B.n459 B.n458 585
R219 B.n461 B.n382 585
R220 B.n464 B.n463 585
R221 B.n465 B.n381 585
R222 B.n467 B.n466 585
R223 B.n469 B.n380 585
R224 B.n472 B.n471 585
R225 B.n473 B.n379 585
R226 B.n475 B.n474 585
R227 B.n477 B.n378 585
R228 B.n480 B.n479 585
R229 B.n481 B.n377 585
R230 B.n483 B.n482 585
R231 B.n485 B.n376 585
R232 B.n488 B.n487 585
R233 B.n489 B.n373 585
R234 B.n492 B.n491 585
R235 B.n494 B.n372 585
R236 B.n497 B.n496 585
R237 B.n498 B.n371 585
R238 B.n500 B.n499 585
R239 B.n502 B.n370 585
R240 B.n505 B.n504 585
R241 B.n506 B.n369 585
R242 B.n508 B.n507 585
R243 B.n510 B.n368 585
R244 B.n513 B.n512 585
R245 B.n514 B.n364 585
R246 B.n516 B.n515 585
R247 B.n518 B.n363 585
R248 B.n521 B.n520 585
R249 B.n522 B.n362 585
R250 B.n524 B.n523 585
R251 B.n526 B.n361 585
R252 B.n529 B.n528 585
R253 B.n530 B.n360 585
R254 B.n532 B.n531 585
R255 B.n534 B.n359 585
R256 B.n537 B.n536 585
R257 B.n538 B.n358 585
R258 B.n540 B.n539 585
R259 B.n542 B.n357 585
R260 B.n545 B.n544 585
R261 B.n546 B.n356 585
R262 B.n548 B.n547 585
R263 B.n550 B.n355 585
R264 B.n553 B.n552 585
R265 B.n554 B.n354 585
R266 B.n556 B.n555 585
R267 B.n558 B.n353 585
R268 B.n561 B.n560 585
R269 B.n562 B.n352 585
R270 B.n564 B.n563 585
R271 B.n566 B.n351 585
R272 B.n569 B.n568 585
R273 B.n570 B.n350 585
R274 B.n572 B.n571 585
R275 B.n574 B.n349 585
R276 B.n577 B.n576 585
R277 B.n578 B.n348 585
R278 B.n580 B.n579 585
R279 B.n582 B.n347 585
R280 B.n585 B.n584 585
R281 B.n586 B.n346 585
R282 B.n588 B.n587 585
R283 B.n590 B.n345 585
R284 B.n593 B.n592 585
R285 B.n594 B.n344 585
R286 B.n596 B.n595 585
R287 B.n598 B.n343 585
R288 B.n599 B.n342 585
R289 B.n602 B.n601 585
R290 B.n603 B.n341 585
R291 B.n341 B.n340 585
R292 B.n608 B.n607 585
R293 B.n607 B.n606 585
R294 B.n609 B.n337 585
R295 B.n337 B.n336 585
R296 B.n611 B.n610 585
R297 B.n612 B.n611 585
R298 B.n331 B.n330 585
R299 B.n332 B.n331 585
R300 B.n620 B.n619 585
R301 B.n619 B.n618 585
R302 B.n621 B.n329 585
R303 B.n329 B.n328 585
R304 B.n623 B.n622 585
R305 B.n624 B.n623 585
R306 B.n323 B.n322 585
R307 B.n324 B.n323 585
R308 B.n632 B.n631 585
R309 B.n631 B.n630 585
R310 B.n633 B.n321 585
R311 B.n321 B.n320 585
R312 B.n635 B.n634 585
R313 B.n636 B.n635 585
R314 B.n315 B.n314 585
R315 B.n316 B.n315 585
R316 B.n644 B.n643 585
R317 B.n643 B.n642 585
R318 B.n645 B.n313 585
R319 B.n313 B.n311 585
R320 B.n647 B.n646 585
R321 B.n648 B.n647 585
R322 B.n307 B.n306 585
R323 B.n312 B.n307 585
R324 B.n657 B.n656 585
R325 B.n656 B.n655 585
R326 B.n658 B.n305 585
R327 B.n305 B.n304 585
R328 B.n660 B.n659 585
R329 B.n661 B.n660 585
R330 B.n2 B.n0 585
R331 B.n4 B.n2 585
R332 B.n3 B.n1 585
R333 B.n734 B.n3 585
R334 B.n732 B.n731 585
R335 B.n733 B.n732 585
R336 B.n730 B.n9 585
R337 B.n9 B.n8 585
R338 B.n729 B.n728 585
R339 B.n728 B.n727 585
R340 B.n11 B.n10 585
R341 B.n726 B.n11 585
R342 B.n724 B.n723 585
R343 B.n725 B.n724 585
R344 B.n722 B.n16 585
R345 B.n16 B.n15 585
R346 B.n721 B.n720 585
R347 B.n720 B.n719 585
R348 B.n18 B.n17 585
R349 B.n718 B.n18 585
R350 B.n716 B.n715 585
R351 B.n717 B.n716 585
R352 B.n714 B.n23 585
R353 B.n23 B.n22 585
R354 B.n713 B.n712 585
R355 B.n712 B.n711 585
R356 B.n25 B.n24 585
R357 B.n710 B.n25 585
R358 B.n708 B.n707 585
R359 B.n709 B.n708 585
R360 B.n706 B.n30 585
R361 B.n30 B.n29 585
R362 B.n705 B.n704 585
R363 B.n704 B.n703 585
R364 B.n32 B.n31 585
R365 B.n702 B.n32 585
R366 B.n700 B.n699 585
R367 B.n701 B.n700 585
R368 B.n698 B.n37 585
R369 B.n37 B.n36 585
R370 B.n697 B.n696 585
R371 B.n696 B.n695 585
R372 B.n737 B.n736 585
R373 B.n736 B.n735 585
R374 B.n607 B.n339 569.379
R375 B.n696 B.n39 569.379
R376 B.n605 B.n341 569.379
R377 B.n692 B.n40 569.379
R378 B.n365 B.t6 400.815
R379 B.n374 B.t13 400.815
R380 B.n95 B.t10 400.815
R381 B.n93 B.t2 400.815
R382 B.n365 B.t9 355.74
R383 B.n93 B.t4 355.74
R384 B.n374 B.t15 355.74
R385 B.n95 B.t11 355.74
R386 B.n366 B.t8 315.788
R387 B.n94 B.t5 315.788
R388 B.n375 B.t14 315.788
R389 B.n96 B.t12 315.788
R390 B.n694 B.n693 256.663
R391 B.n694 B.n91 256.663
R392 B.n694 B.n90 256.663
R393 B.n694 B.n89 256.663
R394 B.n694 B.n88 256.663
R395 B.n694 B.n87 256.663
R396 B.n694 B.n86 256.663
R397 B.n694 B.n85 256.663
R398 B.n694 B.n84 256.663
R399 B.n694 B.n83 256.663
R400 B.n694 B.n82 256.663
R401 B.n694 B.n81 256.663
R402 B.n694 B.n80 256.663
R403 B.n694 B.n79 256.663
R404 B.n694 B.n78 256.663
R405 B.n694 B.n77 256.663
R406 B.n694 B.n76 256.663
R407 B.n694 B.n75 256.663
R408 B.n694 B.n74 256.663
R409 B.n694 B.n73 256.663
R410 B.n694 B.n72 256.663
R411 B.n694 B.n71 256.663
R412 B.n694 B.n70 256.663
R413 B.n694 B.n69 256.663
R414 B.n694 B.n68 256.663
R415 B.n694 B.n67 256.663
R416 B.n694 B.n66 256.663
R417 B.n694 B.n65 256.663
R418 B.n694 B.n64 256.663
R419 B.n694 B.n63 256.663
R420 B.n694 B.n62 256.663
R421 B.n694 B.n61 256.663
R422 B.n694 B.n60 256.663
R423 B.n694 B.n59 256.663
R424 B.n694 B.n58 256.663
R425 B.n694 B.n57 256.663
R426 B.n694 B.n56 256.663
R427 B.n694 B.n55 256.663
R428 B.n694 B.n54 256.663
R429 B.n694 B.n53 256.663
R430 B.n694 B.n52 256.663
R431 B.n694 B.n51 256.663
R432 B.n694 B.n50 256.663
R433 B.n694 B.n49 256.663
R434 B.n694 B.n48 256.663
R435 B.n694 B.n47 256.663
R436 B.n694 B.n46 256.663
R437 B.n694 B.n45 256.663
R438 B.n694 B.n44 256.663
R439 B.n694 B.n43 256.663
R440 B.n694 B.n42 256.663
R441 B.n694 B.n41 256.663
R442 B.n398 B.n340 256.663
R443 B.n404 B.n340 256.663
R444 B.n406 B.n340 256.663
R445 B.n412 B.n340 256.663
R446 B.n414 B.n340 256.663
R447 B.n420 B.n340 256.663
R448 B.n422 B.n340 256.663
R449 B.n428 B.n340 256.663
R450 B.n430 B.n340 256.663
R451 B.n436 B.n340 256.663
R452 B.n438 B.n340 256.663
R453 B.n444 B.n340 256.663
R454 B.n446 B.n340 256.663
R455 B.n452 B.n340 256.663
R456 B.n454 B.n340 256.663
R457 B.n460 B.n340 256.663
R458 B.n462 B.n340 256.663
R459 B.n468 B.n340 256.663
R460 B.n470 B.n340 256.663
R461 B.n476 B.n340 256.663
R462 B.n478 B.n340 256.663
R463 B.n484 B.n340 256.663
R464 B.n486 B.n340 256.663
R465 B.n493 B.n340 256.663
R466 B.n495 B.n340 256.663
R467 B.n501 B.n340 256.663
R468 B.n503 B.n340 256.663
R469 B.n509 B.n340 256.663
R470 B.n511 B.n340 256.663
R471 B.n517 B.n340 256.663
R472 B.n519 B.n340 256.663
R473 B.n525 B.n340 256.663
R474 B.n527 B.n340 256.663
R475 B.n533 B.n340 256.663
R476 B.n535 B.n340 256.663
R477 B.n541 B.n340 256.663
R478 B.n543 B.n340 256.663
R479 B.n549 B.n340 256.663
R480 B.n551 B.n340 256.663
R481 B.n557 B.n340 256.663
R482 B.n559 B.n340 256.663
R483 B.n565 B.n340 256.663
R484 B.n567 B.n340 256.663
R485 B.n573 B.n340 256.663
R486 B.n575 B.n340 256.663
R487 B.n581 B.n340 256.663
R488 B.n583 B.n340 256.663
R489 B.n589 B.n340 256.663
R490 B.n591 B.n340 256.663
R491 B.n597 B.n340 256.663
R492 B.n600 B.n340 256.663
R493 B.n607 B.n337 163.367
R494 B.n611 B.n337 163.367
R495 B.n611 B.n331 163.367
R496 B.n619 B.n331 163.367
R497 B.n619 B.n329 163.367
R498 B.n623 B.n329 163.367
R499 B.n623 B.n323 163.367
R500 B.n631 B.n323 163.367
R501 B.n631 B.n321 163.367
R502 B.n635 B.n321 163.367
R503 B.n635 B.n315 163.367
R504 B.n643 B.n315 163.367
R505 B.n643 B.n313 163.367
R506 B.n647 B.n313 163.367
R507 B.n647 B.n307 163.367
R508 B.n656 B.n307 163.367
R509 B.n656 B.n305 163.367
R510 B.n660 B.n305 163.367
R511 B.n660 B.n2 163.367
R512 B.n736 B.n2 163.367
R513 B.n736 B.n3 163.367
R514 B.n732 B.n3 163.367
R515 B.n732 B.n9 163.367
R516 B.n728 B.n9 163.367
R517 B.n728 B.n11 163.367
R518 B.n724 B.n11 163.367
R519 B.n724 B.n16 163.367
R520 B.n720 B.n16 163.367
R521 B.n720 B.n18 163.367
R522 B.n716 B.n18 163.367
R523 B.n716 B.n23 163.367
R524 B.n712 B.n23 163.367
R525 B.n712 B.n25 163.367
R526 B.n708 B.n25 163.367
R527 B.n708 B.n30 163.367
R528 B.n704 B.n30 163.367
R529 B.n704 B.n32 163.367
R530 B.n700 B.n32 163.367
R531 B.n700 B.n37 163.367
R532 B.n696 B.n37 163.367
R533 B.n399 B.n397 163.367
R534 B.n403 B.n397 163.367
R535 B.n407 B.n405 163.367
R536 B.n411 B.n395 163.367
R537 B.n415 B.n413 163.367
R538 B.n419 B.n393 163.367
R539 B.n423 B.n421 163.367
R540 B.n427 B.n391 163.367
R541 B.n431 B.n429 163.367
R542 B.n435 B.n389 163.367
R543 B.n439 B.n437 163.367
R544 B.n443 B.n387 163.367
R545 B.n447 B.n445 163.367
R546 B.n451 B.n385 163.367
R547 B.n455 B.n453 163.367
R548 B.n459 B.n383 163.367
R549 B.n463 B.n461 163.367
R550 B.n467 B.n381 163.367
R551 B.n471 B.n469 163.367
R552 B.n475 B.n379 163.367
R553 B.n479 B.n477 163.367
R554 B.n483 B.n377 163.367
R555 B.n487 B.n485 163.367
R556 B.n492 B.n373 163.367
R557 B.n496 B.n494 163.367
R558 B.n500 B.n371 163.367
R559 B.n504 B.n502 163.367
R560 B.n508 B.n369 163.367
R561 B.n512 B.n510 163.367
R562 B.n516 B.n364 163.367
R563 B.n520 B.n518 163.367
R564 B.n524 B.n362 163.367
R565 B.n528 B.n526 163.367
R566 B.n532 B.n360 163.367
R567 B.n536 B.n534 163.367
R568 B.n540 B.n358 163.367
R569 B.n544 B.n542 163.367
R570 B.n548 B.n356 163.367
R571 B.n552 B.n550 163.367
R572 B.n556 B.n354 163.367
R573 B.n560 B.n558 163.367
R574 B.n564 B.n352 163.367
R575 B.n568 B.n566 163.367
R576 B.n572 B.n350 163.367
R577 B.n576 B.n574 163.367
R578 B.n580 B.n348 163.367
R579 B.n584 B.n582 163.367
R580 B.n588 B.n346 163.367
R581 B.n592 B.n590 163.367
R582 B.n596 B.n344 163.367
R583 B.n599 B.n598 163.367
R584 B.n601 B.n341 163.367
R585 B.n605 B.n335 163.367
R586 B.n613 B.n335 163.367
R587 B.n613 B.n333 163.367
R588 B.n617 B.n333 163.367
R589 B.n617 B.n327 163.367
R590 B.n625 B.n327 163.367
R591 B.n625 B.n325 163.367
R592 B.n629 B.n325 163.367
R593 B.n629 B.n319 163.367
R594 B.n637 B.n319 163.367
R595 B.n637 B.n317 163.367
R596 B.n641 B.n317 163.367
R597 B.n641 B.n310 163.367
R598 B.n649 B.n310 163.367
R599 B.n649 B.n308 163.367
R600 B.n654 B.n308 163.367
R601 B.n654 B.n303 163.367
R602 B.n662 B.n303 163.367
R603 B.n663 B.n662 163.367
R604 B.n663 B.n5 163.367
R605 B.n6 B.n5 163.367
R606 B.n7 B.n6 163.367
R607 B.n668 B.n7 163.367
R608 B.n668 B.n12 163.367
R609 B.n13 B.n12 163.367
R610 B.n14 B.n13 163.367
R611 B.n673 B.n14 163.367
R612 B.n673 B.n19 163.367
R613 B.n20 B.n19 163.367
R614 B.n21 B.n20 163.367
R615 B.n678 B.n21 163.367
R616 B.n678 B.n26 163.367
R617 B.n27 B.n26 163.367
R618 B.n28 B.n27 163.367
R619 B.n683 B.n28 163.367
R620 B.n683 B.n33 163.367
R621 B.n34 B.n33 163.367
R622 B.n35 B.n34 163.367
R623 B.n688 B.n35 163.367
R624 B.n688 B.n40 163.367
R625 B.n99 B.n98 163.367
R626 B.n103 B.n102 163.367
R627 B.n107 B.n106 163.367
R628 B.n111 B.n110 163.367
R629 B.n115 B.n114 163.367
R630 B.n119 B.n118 163.367
R631 B.n123 B.n122 163.367
R632 B.n127 B.n126 163.367
R633 B.n131 B.n130 163.367
R634 B.n135 B.n134 163.367
R635 B.n139 B.n138 163.367
R636 B.n143 B.n142 163.367
R637 B.n147 B.n146 163.367
R638 B.n151 B.n150 163.367
R639 B.n155 B.n154 163.367
R640 B.n159 B.n158 163.367
R641 B.n163 B.n162 163.367
R642 B.n167 B.n166 163.367
R643 B.n171 B.n170 163.367
R644 B.n175 B.n174 163.367
R645 B.n179 B.n178 163.367
R646 B.n183 B.n182 163.367
R647 B.n187 B.n186 163.367
R648 B.n192 B.n191 163.367
R649 B.n196 B.n195 163.367
R650 B.n200 B.n199 163.367
R651 B.n204 B.n203 163.367
R652 B.n208 B.n207 163.367
R653 B.n213 B.n212 163.367
R654 B.n217 B.n216 163.367
R655 B.n221 B.n220 163.367
R656 B.n225 B.n224 163.367
R657 B.n229 B.n228 163.367
R658 B.n233 B.n232 163.367
R659 B.n237 B.n236 163.367
R660 B.n241 B.n240 163.367
R661 B.n245 B.n244 163.367
R662 B.n249 B.n248 163.367
R663 B.n253 B.n252 163.367
R664 B.n257 B.n256 163.367
R665 B.n261 B.n260 163.367
R666 B.n265 B.n264 163.367
R667 B.n269 B.n268 163.367
R668 B.n273 B.n272 163.367
R669 B.n277 B.n276 163.367
R670 B.n281 B.n280 163.367
R671 B.n285 B.n284 163.367
R672 B.n289 B.n288 163.367
R673 B.n293 B.n292 163.367
R674 B.n297 B.n296 163.367
R675 B.n299 B.n92 163.367
R676 B.n606 B.n340 79.4497
R677 B.n695 B.n694 79.4497
R678 B.n398 B.n339 71.676
R679 B.n404 B.n403 71.676
R680 B.n407 B.n406 71.676
R681 B.n412 B.n411 71.676
R682 B.n415 B.n414 71.676
R683 B.n420 B.n419 71.676
R684 B.n423 B.n422 71.676
R685 B.n428 B.n427 71.676
R686 B.n431 B.n430 71.676
R687 B.n436 B.n435 71.676
R688 B.n439 B.n438 71.676
R689 B.n444 B.n443 71.676
R690 B.n447 B.n446 71.676
R691 B.n452 B.n451 71.676
R692 B.n455 B.n454 71.676
R693 B.n460 B.n459 71.676
R694 B.n463 B.n462 71.676
R695 B.n468 B.n467 71.676
R696 B.n471 B.n470 71.676
R697 B.n476 B.n475 71.676
R698 B.n479 B.n478 71.676
R699 B.n484 B.n483 71.676
R700 B.n487 B.n486 71.676
R701 B.n493 B.n492 71.676
R702 B.n496 B.n495 71.676
R703 B.n501 B.n500 71.676
R704 B.n504 B.n503 71.676
R705 B.n509 B.n508 71.676
R706 B.n512 B.n511 71.676
R707 B.n517 B.n516 71.676
R708 B.n520 B.n519 71.676
R709 B.n525 B.n524 71.676
R710 B.n528 B.n527 71.676
R711 B.n533 B.n532 71.676
R712 B.n536 B.n535 71.676
R713 B.n541 B.n540 71.676
R714 B.n544 B.n543 71.676
R715 B.n549 B.n548 71.676
R716 B.n552 B.n551 71.676
R717 B.n557 B.n556 71.676
R718 B.n560 B.n559 71.676
R719 B.n565 B.n564 71.676
R720 B.n568 B.n567 71.676
R721 B.n573 B.n572 71.676
R722 B.n576 B.n575 71.676
R723 B.n581 B.n580 71.676
R724 B.n584 B.n583 71.676
R725 B.n589 B.n588 71.676
R726 B.n592 B.n591 71.676
R727 B.n597 B.n596 71.676
R728 B.n600 B.n599 71.676
R729 B.n41 B.n39 71.676
R730 B.n99 B.n42 71.676
R731 B.n103 B.n43 71.676
R732 B.n107 B.n44 71.676
R733 B.n111 B.n45 71.676
R734 B.n115 B.n46 71.676
R735 B.n119 B.n47 71.676
R736 B.n123 B.n48 71.676
R737 B.n127 B.n49 71.676
R738 B.n131 B.n50 71.676
R739 B.n135 B.n51 71.676
R740 B.n139 B.n52 71.676
R741 B.n143 B.n53 71.676
R742 B.n147 B.n54 71.676
R743 B.n151 B.n55 71.676
R744 B.n155 B.n56 71.676
R745 B.n159 B.n57 71.676
R746 B.n163 B.n58 71.676
R747 B.n167 B.n59 71.676
R748 B.n171 B.n60 71.676
R749 B.n175 B.n61 71.676
R750 B.n179 B.n62 71.676
R751 B.n183 B.n63 71.676
R752 B.n187 B.n64 71.676
R753 B.n192 B.n65 71.676
R754 B.n196 B.n66 71.676
R755 B.n200 B.n67 71.676
R756 B.n204 B.n68 71.676
R757 B.n208 B.n69 71.676
R758 B.n213 B.n70 71.676
R759 B.n217 B.n71 71.676
R760 B.n221 B.n72 71.676
R761 B.n225 B.n73 71.676
R762 B.n229 B.n74 71.676
R763 B.n233 B.n75 71.676
R764 B.n237 B.n76 71.676
R765 B.n241 B.n77 71.676
R766 B.n245 B.n78 71.676
R767 B.n249 B.n79 71.676
R768 B.n253 B.n80 71.676
R769 B.n257 B.n81 71.676
R770 B.n261 B.n82 71.676
R771 B.n265 B.n83 71.676
R772 B.n269 B.n84 71.676
R773 B.n273 B.n85 71.676
R774 B.n277 B.n86 71.676
R775 B.n281 B.n87 71.676
R776 B.n285 B.n88 71.676
R777 B.n289 B.n89 71.676
R778 B.n293 B.n90 71.676
R779 B.n297 B.n91 71.676
R780 B.n693 B.n92 71.676
R781 B.n693 B.n692 71.676
R782 B.n299 B.n91 71.676
R783 B.n296 B.n90 71.676
R784 B.n292 B.n89 71.676
R785 B.n288 B.n88 71.676
R786 B.n284 B.n87 71.676
R787 B.n280 B.n86 71.676
R788 B.n276 B.n85 71.676
R789 B.n272 B.n84 71.676
R790 B.n268 B.n83 71.676
R791 B.n264 B.n82 71.676
R792 B.n260 B.n81 71.676
R793 B.n256 B.n80 71.676
R794 B.n252 B.n79 71.676
R795 B.n248 B.n78 71.676
R796 B.n244 B.n77 71.676
R797 B.n240 B.n76 71.676
R798 B.n236 B.n75 71.676
R799 B.n232 B.n74 71.676
R800 B.n228 B.n73 71.676
R801 B.n224 B.n72 71.676
R802 B.n220 B.n71 71.676
R803 B.n216 B.n70 71.676
R804 B.n212 B.n69 71.676
R805 B.n207 B.n68 71.676
R806 B.n203 B.n67 71.676
R807 B.n199 B.n66 71.676
R808 B.n195 B.n65 71.676
R809 B.n191 B.n64 71.676
R810 B.n186 B.n63 71.676
R811 B.n182 B.n62 71.676
R812 B.n178 B.n61 71.676
R813 B.n174 B.n60 71.676
R814 B.n170 B.n59 71.676
R815 B.n166 B.n58 71.676
R816 B.n162 B.n57 71.676
R817 B.n158 B.n56 71.676
R818 B.n154 B.n55 71.676
R819 B.n150 B.n54 71.676
R820 B.n146 B.n53 71.676
R821 B.n142 B.n52 71.676
R822 B.n138 B.n51 71.676
R823 B.n134 B.n50 71.676
R824 B.n130 B.n49 71.676
R825 B.n126 B.n48 71.676
R826 B.n122 B.n47 71.676
R827 B.n118 B.n46 71.676
R828 B.n114 B.n45 71.676
R829 B.n110 B.n44 71.676
R830 B.n106 B.n43 71.676
R831 B.n102 B.n42 71.676
R832 B.n98 B.n41 71.676
R833 B.n399 B.n398 71.676
R834 B.n405 B.n404 71.676
R835 B.n406 B.n395 71.676
R836 B.n413 B.n412 71.676
R837 B.n414 B.n393 71.676
R838 B.n421 B.n420 71.676
R839 B.n422 B.n391 71.676
R840 B.n429 B.n428 71.676
R841 B.n430 B.n389 71.676
R842 B.n437 B.n436 71.676
R843 B.n438 B.n387 71.676
R844 B.n445 B.n444 71.676
R845 B.n446 B.n385 71.676
R846 B.n453 B.n452 71.676
R847 B.n454 B.n383 71.676
R848 B.n461 B.n460 71.676
R849 B.n462 B.n381 71.676
R850 B.n469 B.n468 71.676
R851 B.n470 B.n379 71.676
R852 B.n477 B.n476 71.676
R853 B.n478 B.n377 71.676
R854 B.n485 B.n484 71.676
R855 B.n486 B.n373 71.676
R856 B.n494 B.n493 71.676
R857 B.n495 B.n371 71.676
R858 B.n502 B.n501 71.676
R859 B.n503 B.n369 71.676
R860 B.n510 B.n509 71.676
R861 B.n511 B.n364 71.676
R862 B.n518 B.n517 71.676
R863 B.n519 B.n362 71.676
R864 B.n526 B.n525 71.676
R865 B.n527 B.n360 71.676
R866 B.n534 B.n533 71.676
R867 B.n535 B.n358 71.676
R868 B.n542 B.n541 71.676
R869 B.n543 B.n356 71.676
R870 B.n550 B.n549 71.676
R871 B.n551 B.n354 71.676
R872 B.n558 B.n557 71.676
R873 B.n559 B.n352 71.676
R874 B.n566 B.n565 71.676
R875 B.n567 B.n350 71.676
R876 B.n574 B.n573 71.676
R877 B.n575 B.n348 71.676
R878 B.n582 B.n581 71.676
R879 B.n583 B.n346 71.676
R880 B.n590 B.n589 71.676
R881 B.n591 B.n344 71.676
R882 B.n598 B.n597 71.676
R883 B.n601 B.n600 71.676
R884 B.n367 B.n366 59.5399
R885 B.n490 B.n375 59.5399
R886 B.n189 B.n96 59.5399
R887 B.n210 B.n94 59.5399
R888 B.n366 B.n365 39.952
R889 B.n375 B.n374 39.952
R890 B.n96 B.n95 39.952
R891 B.n94 B.n93 39.952
R892 B.n606 B.n336 38.8677
R893 B.n612 B.n336 38.8677
R894 B.n612 B.n332 38.8677
R895 B.n618 B.n332 38.8677
R896 B.n618 B.n328 38.8677
R897 B.n624 B.n328 38.8677
R898 B.n630 B.n324 38.8677
R899 B.n630 B.n320 38.8677
R900 B.n636 B.n320 38.8677
R901 B.n636 B.n316 38.8677
R902 B.n642 B.n316 38.8677
R903 B.n642 B.n311 38.8677
R904 B.n648 B.n311 38.8677
R905 B.n648 B.n312 38.8677
R906 B.n655 B.n304 38.8677
R907 B.n661 B.n304 38.8677
R908 B.n661 B.n4 38.8677
R909 B.n735 B.n4 38.8677
R910 B.n735 B.n734 38.8677
R911 B.n734 B.n733 38.8677
R912 B.n733 B.n8 38.8677
R913 B.n727 B.n8 38.8677
R914 B.n726 B.n725 38.8677
R915 B.n725 B.n15 38.8677
R916 B.n719 B.n15 38.8677
R917 B.n719 B.n718 38.8677
R918 B.n718 B.n717 38.8677
R919 B.n717 B.n22 38.8677
R920 B.n711 B.n22 38.8677
R921 B.n711 B.n710 38.8677
R922 B.n709 B.n29 38.8677
R923 B.n703 B.n29 38.8677
R924 B.n703 B.n702 38.8677
R925 B.n702 B.n701 38.8677
R926 B.n701 B.n36 38.8677
R927 B.n695 B.n36 38.8677
R928 B.n697 B.n38 36.9956
R929 B.n691 B.n690 36.9956
R930 B.n604 B.n603 36.9956
R931 B.n608 B.n338 36.9956
R932 B.t7 B.n324 34.8667
R933 B.n710 B.t3 34.8667
R934 B.n655 B.t0 24.5783
R935 B.n727 B.t1 24.5783
R936 B B.n737 18.0485
R937 B.n312 B.t0 14.2899
R938 B.t1 B.n726 14.2899
R939 B.n97 B.n38 10.6151
R940 B.n100 B.n97 10.6151
R941 B.n101 B.n100 10.6151
R942 B.n104 B.n101 10.6151
R943 B.n105 B.n104 10.6151
R944 B.n108 B.n105 10.6151
R945 B.n109 B.n108 10.6151
R946 B.n112 B.n109 10.6151
R947 B.n113 B.n112 10.6151
R948 B.n116 B.n113 10.6151
R949 B.n117 B.n116 10.6151
R950 B.n120 B.n117 10.6151
R951 B.n121 B.n120 10.6151
R952 B.n124 B.n121 10.6151
R953 B.n125 B.n124 10.6151
R954 B.n128 B.n125 10.6151
R955 B.n129 B.n128 10.6151
R956 B.n132 B.n129 10.6151
R957 B.n133 B.n132 10.6151
R958 B.n136 B.n133 10.6151
R959 B.n137 B.n136 10.6151
R960 B.n140 B.n137 10.6151
R961 B.n141 B.n140 10.6151
R962 B.n144 B.n141 10.6151
R963 B.n145 B.n144 10.6151
R964 B.n148 B.n145 10.6151
R965 B.n149 B.n148 10.6151
R966 B.n152 B.n149 10.6151
R967 B.n153 B.n152 10.6151
R968 B.n156 B.n153 10.6151
R969 B.n157 B.n156 10.6151
R970 B.n160 B.n157 10.6151
R971 B.n161 B.n160 10.6151
R972 B.n164 B.n161 10.6151
R973 B.n165 B.n164 10.6151
R974 B.n168 B.n165 10.6151
R975 B.n169 B.n168 10.6151
R976 B.n172 B.n169 10.6151
R977 B.n173 B.n172 10.6151
R978 B.n176 B.n173 10.6151
R979 B.n177 B.n176 10.6151
R980 B.n180 B.n177 10.6151
R981 B.n181 B.n180 10.6151
R982 B.n184 B.n181 10.6151
R983 B.n185 B.n184 10.6151
R984 B.n188 B.n185 10.6151
R985 B.n193 B.n190 10.6151
R986 B.n194 B.n193 10.6151
R987 B.n197 B.n194 10.6151
R988 B.n198 B.n197 10.6151
R989 B.n201 B.n198 10.6151
R990 B.n202 B.n201 10.6151
R991 B.n205 B.n202 10.6151
R992 B.n206 B.n205 10.6151
R993 B.n209 B.n206 10.6151
R994 B.n214 B.n211 10.6151
R995 B.n215 B.n214 10.6151
R996 B.n218 B.n215 10.6151
R997 B.n219 B.n218 10.6151
R998 B.n222 B.n219 10.6151
R999 B.n223 B.n222 10.6151
R1000 B.n226 B.n223 10.6151
R1001 B.n227 B.n226 10.6151
R1002 B.n230 B.n227 10.6151
R1003 B.n231 B.n230 10.6151
R1004 B.n234 B.n231 10.6151
R1005 B.n235 B.n234 10.6151
R1006 B.n238 B.n235 10.6151
R1007 B.n239 B.n238 10.6151
R1008 B.n242 B.n239 10.6151
R1009 B.n243 B.n242 10.6151
R1010 B.n246 B.n243 10.6151
R1011 B.n247 B.n246 10.6151
R1012 B.n250 B.n247 10.6151
R1013 B.n251 B.n250 10.6151
R1014 B.n254 B.n251 10.6151
R1015 B.n255 B.n254 10.6151
R1016 B.n258 B.n255 10.6151
R1017 B.n259 B.n258 10.6151
R1018 B.n262 B.n259 10.6151
R1019 B.n263 B.n262 10.6151
R1020 B.n266 B.n263 10.6151
R1021 B.n267 B.n266 10.6151
R1022 B.n270 B.n267 10.6151
R1023 B.n271 B.n270 10.6151
R1024 B.n274 B.n271 10.6151
R1025 B.n275 B.n274 10.6151
R1026 B.n278 B.n275 10.6151
R1027 B.n279 B.n278 10.6151
R1028 B.n282 B.n279 10.6151
R1029 B.n283 B.n282 10.6151
R1030 B.n286 B.n283 10.6151
R1031 B.n287 B.n286 10.6151
R1032 B.n290 B.n287 10.6151
R1033 B.n291 B.n290 10.6151
R1034 B.n294 B.n291 10.6151
R1035 B.n295 B.n294 10.6151
R1036 B.n298 B.n295 10.6151
R1037 B.n300 B.n298 10.6151
R1038 B.n301 B.n300 10.6151
R1039 B.n691 B.n301 10.6151
R1040 B.n604 B.n334 10.6151
R1041 B.n614 B.n334 10.6151
R1042 B.n615 B.n614 10.6151
R1043 B.n616 B.n615 10.6151
R1044 B.n616 B.n326 10.6151
R1045 B.n626 B.n326 10.6151
R1046 B.n627 B.n626 10.6151
R1047 B.n628 B.n627 10.6151
R1048 B.n628 B.n318 10.6151
R1049 B.n638 B.n318 10.6151
R1050 B.n639 B.n638 10.6151
R1051 B.n640 B.n639 10.6151
R1052 B.n640 B.n309 10.6151
R1053 B.n650 B.n309 10.6151
R1054 B.n651 B.n650 10.6151
R1055 B.n653 B.n651 10.6151
R1056 B.n653 B.n652 10.6151
R1057 B.n652 B.n302 10.6151
R1058 B.n664 B.n302 10.6151
R1059 B.n665 B.n664 10.6151
R1060 B.n666 B.n665 10.6151
R1061 B.n667 B.n666 10.6151
R1062 B.n669 B.n667 10.6151
R1063 B.n670 B.n669 10.6151
R1064 B.n671 B.n670 10.6151
R1065 B.n672 B.n671 10.6151
R1066 B.n674 B.n672 10.6151
R1067 B.n675 B.n674 10.6151
R1068 B.n676 B.n675 10.6151
R1069 B.n677 B.n676 10.6151
R1070 B.n679 B.n677 10.6151
R1071 B.n680 B.n679 10.6151
R1072 B.n681 B.n680 10.6151
R1073 B.n682 B.n681 10.6151
R1074 B.n684 B.n682 10.6151
R1075 B.n685 B.n684 10.6151
R1076 B.n686 B.n685 10.6151
R1077 B.n687 B.n686 10.6151
R1078 B.n689 B.n687 10.6151
R1079 B.n690 B.n689 10.6151
R1080 B.n400 B.n338 10.6151
R1081 B.n401 B.n400 10.6151
R1082 B.n402 B.n401 10.6151
R1083 B.n402 B.n396 10.6151
R1084 B.n408 B.n396 10.6151
R1085 B.n409 B.n408 10.6151
R1086 B.n410 B.n409 10.6151
R1087 B.n410 B.n394 10.6151
R1088 B.n416 B.n394 10.6151
R1089 B.n417 B.n416 10.6151
R1090 B.n418 B.n417 10.6151
R1091 B.n418 B.n392 10.6151
R1092 B.n424 B.n392 10.6151
R1093 B.n425 B.n424 10.6151
R1094 B.n426 B.n425 10.6151
R1095 B.n426 B.n390 10.6151
R1096 B.n432 B.n390 10.6151
R1097 B.n433 B.n432 10.6151
R1098 B.n434 B.n433 10.6151
R1099 B.n434 B.n388 10.6151
R1100 B.n440 B.n388 10.6151
R1101 B.n441 B.n440 10.6151
R1102 B.n442 B.n441 10.6151
R1103 B.n442 B.n386 10.6151
R1104 B.n448 B.n386 10.6151
R1105 B.n449 B.n448 10.6151
R1106 B.n450 B.n449 10.6151
R1107 B.n450 B.n384 10.6151
R1108 B.n456 B.n384 10.6151
R1109 B.n457 B.n456 10.6151
R1110 B.n458 B.n457 10.6151
R1111 B.n458 B.n382 10.6151
R1112 B.n464 B.n382 10.6151
R1113 B.n465 B.n464 10.6151
R1114 B.n466 B.n465 10.6151
R1115 B.n466 B.n380 10.6151
R1116 B.n472 B.n380 10.6151
R1117 B.n473 B.n472 10.6151
R1118 B.n474 B.n473 10.6151
R1119 B.n474 B.n378 10.6151
R1120 B.n480 B.n378 10.6151
R1121 B.n481 B.n480 10.6151
R1122 B.n482 B.n481 10.6151
R1123 B.n482 B.n376 10.6151
R1124 B.n488 B.n376 10.6151
R1125 B.n489 B.n488 10.6151
R1126 B.n491 B.n372 10.6151
R1127 B.n497 B.n372 10.6151
R1128 B.n498 B.n497 10.6151
R1129 B.n499 B.n498 10.6151
R1130 B.n499 B.n370 10.6151
R1131 B.n505 B.n370 10.6151
R1132 B.n506 B.n505 10.6151
R1133 B.n507 B.n506 10.6151
R1134 B.n507 B.n368 10.6151
R1135 B.n514 B.n513 10.6151
R1136 B.n515 B.n514 10.6151
R1137 B.n515 B.n363 10.6151
R1138 B.n521 B.n363 10.6151
R1139 B.n522 B.n521 10.6151
R1140 B.n523 B.n522 10.6151
R1141 B.n523 B.n361 10.6151
R1142 B.n529 B.n361 10.6151
R1143 B.n530 B.n529 10.6151
R1144 B.n531 B.n530 10.6151
R1145 B.n531 B.n359 10.6151
R1146 B.n537 B.n359 10.6151
R1147 B.n538 B.n537 10.6151
R1148 B.n539 B.n538 10.6151
R1149 B.n539 B.n357 10.6151
R1150 B.n545 B.n357 10.6151
R1151 B.n546 B.n545 10.6151
R1152 B.n547 B.n546 10.6151
R1153 B.n547 B.n355 10.6151
R1154 B.n553 B.n355 10.6151
R1155 B.n554 B.n553 10.6151
R1156 B.n555 B.n554 10.6151
R1157 B.n555 B.n353 10.6151
R1158 B.n561 B.n353 10.6151
R1159 B.n562 B.n561 10.6151
R1160 B.n563 B.n562 10.6151
R1161 B.n563 B.n351 10.6151
R1162 B.n569 B.n351 10.6151
R1163 B.n570 B.n569 10.6151
R1164 B.n571 B.n570 10.6151
R1165 B.n571 B.n349 10.6151
R1166 B.n577 B.n349 10.6151
R1167 B.n578 B.n577 10.6151
R1168 B.n579 B.n578 10.6151
R1169 B.n579 B.n347 10.6151
R1170 B.n585 B.n347 10.6151
R1171 B.n586 B.n585 10.6151
R1172 B.n587 B.n586 10.6151
R1173 B.n587 B.n345 10.6151
R1174 B.n593 B.n345 10.6151
R1175 B.n594 B.n593 10.6151
R1176 B.n595 B.n594 10.6151
R1177 B.n595 B.n343 10.6151
R1178 B.n343 B.n342 10.6151
R1179 B.n602 B.n342 10.6151
R1180 B.n603 B.n602 10.6151
R1181 B.n609 B.n608 10.6151
R1182 B.n610 B.n609 10.6151
R1183 B.n610 B.n330 10.6151
R1184 B.n620 B.n330 10.6151
R1185 B.n621 B.n620 10.6151
R1186 B.n622 B.n621 10.6151
R1187 B.n622 B.n322 10.6151
R1188 B.n632 B.n322 10.6151
R1189 B.n633 B.n632 10.6151
R1190 B.n634 B.n633 10.6151
R1191 B.n634 B.n314 10.6151
R1192 B.n644 B.n314 10.6151
R1193 B.n645 B.n644 10.6151
R1194 B.n646 B.n645 10.6151
R1195 B.n646 B.n306 10.6151
R1196 B.n657 B.n306 10.6151
R1197 B.n658 B.n657 10.6151
R1198 B.n659 B.n658 10.6151
R1199 B.n659 B.n0 10.6151
R1200 B.n731 B.n1 10.6151
R1201 B.n731 B.n730 10.6151
R1202 B.n730 B.n729 10.6151
R1203 B.n729 B.n10 10.6151
R1204 B.n723 B.n10 10.6151
R1205 B.n723 B.n722 10.6151
R1206 B.n722 B.n721 10.6151
R1207 B.n721 B.n17 10.6151
R1208 B.n715 B.n17 10.6151
R1209 B.n715 B.n714 10.6151
R1210 B.n714 B.n713 10.6151
R1211 B.n713 B.n24 10.6151
R1212 B.n707 B.n24 10.6151
R1213 B.n707 B.n706 10.6151
R1214 B.n706 B.n705 10.6151
R1215 B.n705 B.n31 10.6151
R1216 B.n699 B.n31 10.6151
R1217 B.n699 B.n698 10.6151
R1218 B.n698 B.n697 10.6151
R1219 B.n189 B.n188 9.36635
R1220 B.n211 B.n210 9.36635
R1221 B.n490 B.n489 9.36635
R1222 B.n513 B.n367 9.36635
R1223 B.n624 B.t7 4.00154
R1224 B.t3 B.n709 4.00154
R1225 B.n737 B.n0 2.81026
R1226 B.n737 B.n1 2.81026
R1227 B.n190 B.n189 1.24928
R1228 B.n210 B.n209 1.24928
R1229 B.n491 B.n490 1.24928
R1230 B.n368 B.n367 1.24928
R1231 VN VN.t0 297.505
R1232 VN VN.t1 253.714
R1233 VTAIL.n306 VTAIL.n234 289.615
R1234 VTAIL.n72 VTAIL.n0 289.615
R1235 VTAIL.n228 VTAIL.n156 289.615
R1236 VTAIL.n150 VTAIL.n78 289.615
R1237 VTAIL.n258 VTAIL.n257 185
R1238 VTAIL.n263 VTAIL.n262 185
R1239 VTAIL.n265 VTAIL.n264 185
R1240 VTAIL.n254 VTAIL.n253 185
R1241 VTAIL.n271 VTAIL.n270 185
R1242 VTAIL.n273 VTAIL.n272 185
R1243 VTAIL.n250 VTAIL.n249 185
R1244 VTAIL.n279 VTAIL.n278 185
R1245 VTAIL.n281 VTAIL.n280 185
R1246 VTAIL.n246 VTAIL.n245 185
R1247 VTAIL.n287 VTAIL.n286 185
R1248 VTAIL.n289 VTAIL.n288 185
R1249 VTAIL.n242 VTAIL.n241 185
R1250 VTAIL.n295 VTAIL.n294 185
R1251 VTAIL.n297 VTAIL.n296 185
R1252 VTAIL.n238 VTAIL.n237 185
R1253 VTAIL.n304 VTAIL.n303 185
R1254 VTAIL.n305 VTAIL.n236 185
R1255 VTAIL.n307 VTAIL.n306 185
R1256 VTAIL.n24 VTAIL.n23 185
R1257 VTAIL.n29 VTAIL.n28 185
R1258 VTAIL.n31 VTAIL.n30 185
R1259 VTAIL.n20 VTAIL.n19 185
R1260 VTAIL.n37 VTAIL.n36 185
R1261 VTAIL.n39 VTAIL.n38 185
R1262 VTAIL.n16 VTAIL.n15 185
R1263 VTAIL.n45 VTAIL.n44 185
R1264 VTAIL.n47 VTAIL.n46 185
R1265 VTAIL.n12 VTAIL.n11 185
R1266 VTAIL.n53 VTAIL.n52 185
R1267 VTAIL.n55 VTAIL.n54 185
R1268 VTAIL.n8 VTAIL.n7 185
R1269 VTAIL.n61 VTAIL.n60 185
R1270 VTAIL.n63 VTAIL.n62 185
R1271 VTAIL.n4 VTAIL.n3 185
R1272 VTAIL.n70 VTAIL.n69 185
R1273 VTAIL.n71 VTAIL.n2 185
R1274 VTAIL.n73 VTAIL.n72 185
R1275 VTAIL.n229 VTAIL.n228 185
R1276 VTAIL.n227 VTAIL.n158 185
R1277 VTAIL.n226 VTAIL.n225 185
R1278 VTAIL.n161 VTAIL.n159 185
R1279 VTAIL.n220 VTAIL.n219 185
R1280 VTAIL.n218 VTAIL.n217 185
R1281 VTAIL.n165 VTAIL.n164 185
R1282 VTAIL.n212 VTAIL.n211 185
R1283 VTAIL.n210 VTAIL.n209 185
R1284 VTAIL.n169 VTAIL.n168 185
R1285 VTAIL.n204 VTAIL.n203 185
R1286 VTAIL.n202 VTAIL.n201 185
R1287 VTAIL.n173 VTAIL.n172 185
R1288 VTAIL.n196 VTAIL.n195 185
R1289 VTAIL.n194 VTAIL.n193 185
R1290 VTAIL.n177 VTAIL.n176 185
R1291 VTAIL.n188 VTAIL.n187 185
R1292 VTAIL.n186 VTAIL.n185 185
R1293 VTAIL.n181 VTAIL.n180 185
R1294 VTAIL.n151 VTAIL.n150 185
R1295 VTAIL.n149 VTAIL.n80 185
R1296 VTAIL.n148 VTAIL.n147 185
R1297 VTAIL.n83 VTAIL.n81 185
R1298 VTAIL.n142 VTAIL.n141 185
R1299 VTAIL.n140 VTAIL.n139 185
R1300 VTAIL.n87 VTAIL.n86 185
R1301 VTAIL.n134 VTAIL.n133 185
R1302 VTAIL.n132 VTAIL.n131 185
R1303 VTAIL.n91 VTAIL.n90 185
R1304 VTAIL.n126 VTAIL.n125 185
R1305 VTAIL.n124 VTAIL.n123 185
R1306 VTAIL.n95 VTAIL.n94 185
R1307 VTAIL.n118 VTAIL.n117 185
R1308 VTAIL.n116 VTAIL.n115 185
R1309 VTAIL.n99 VTAIL.n98 185
R1310 VTAIL.n110 VTAIL.n109 185
R1311 VTAIL.n108 VTAIL.n107 185
R1312 VTAIL.n103 VTAIL.n102 185
R1313 VTAIL.n259 VTAIL.t2 147.659
R1314 VTAIL.n25 VTAIL.t0 147.659
R1315 VTAIL.n182 VTAIL.t1 147.659
R1316 VTAIL.n104 VTAIL.t3 147.659
R1317 VTAIL.n263 VTAIL.n257 104.615
R1318 VTAIL.n264 VTAIL.n263 104.615
R1319 VTAIL.n264 VTAIL.n253 104.615
R1320 VTAIL.n271 VTAIL.n253 104.615
R1321 VTAIL.n272 VTAIL.n271 104.615
R1322 VTAIL.n272 VTAIL.n249 104.615
R1323 VTAIL.n279 VTAIL.n249 104.615
R1324 VTAIL.n280 VTAIL.n279 104.615
R1325 VTAIL.n280 VTAIL.n245 104.615
R1326 VTAIL.n287 VTAIL.n245 104.615
R1327 VTAIL.n288 VTAIL.n287 104.615
R1328 VTAIL.n288 VTAIL.n241 104.615
R1329 VTAIL.n295 VTAIL.n241 104.615
R1330 VTAIL.n296 VTAIL.n295 104.615
R1331 VTAIL.n296 VTAIL.n237 104.615
R1332 VTAIL.n304 VTAIL.n237 104.615
R1333 VTAIL.n305 VTAIL.n304 104.615
R1334 VTAIL.n306 VTAIL.n305 104.615
R1335 VTAIL.n29 VTAIL.n23 104.615
R1336 VTAIL.n30 VTAIL.n29 104.615
R1337 VTAIL.n30 VTAIL.n19 104.615
R1338 VTAIL.n37 VTAIL.n19 104.615
R1339 VTAIL.n38 VTAIL.n37 104.615
R1340 VTAIL.n38 VTAIL.n15 104.615
R1341 VTAIL.n45 VTAIL.n15 104.615
R1342 VTAIL.n46 VTAIL.n45 104.615
R1343 VTAIL.n46 VTAIL.n11 104.615
R1344 VTAIL.n53 VTAIL.n11 104.615
R1345 VTAIL.n54 VTAIL.n53 104.615
R1346 VTAIL.n54 VTAIL.n7 104.615
R1347 VTAIL.n61 VTAIL.n7 104.615
R1348 VTAIL.n62 VTAIL.n61 104.615
R1349 VTAIL.n62 VTAIL.n3 104.615
R1350 VTAIL.n70 VTAIL.n3 104.615
R1351 VTAIL.n71 VTAIL.n70 104.615
R1352 VTAIL.n72 VTAIL.n71 104.615
R1353 VTAIL.n228 VTAIL.n227 104.615
R1354 VTAIL.n227 VTAIL.n226 104.615
R1355 VTAIL.n226 VTAIL.n159 104.615
R1356 VTAIL.n219 VTAIL.n159 104.615
R1357 VTAIL.n219 VTAIL.n218 104.615
R1358 VTAIL.n218 VTAIL.n164 104.615
R1359 VTAIL.n211 VTAIL.n164 104.615
R1360 VTAIL.n211 VTAIL.n210 104.615
R1361 VTAIL.n210 VTAIL.n168 104.615
R1362 VTAIL.n203 VTAIL.n168 104.615
R1363 VTAIL.n203 VTAIL.n202 104.615
R1364 VTAIL.n202 VTAIL.n172 104.615
R1365 VTAIL.n195 VTAIL.n172 104.615
R1366 VTAIL.n195 VTAIL.n194 104.615
R1367 VTAIL.n194 VTAIL.n176 104.615
R1368 VTAIL.n187 VTAIL.n176 104.615
R1369 VTAIL.n187 VTAIL.n186 104.615
R1370 VTAIL.n186 VTAIL.n180 104.615
R1371 VTAIL.n150 VTAIL.n149 104.615
R1372 VTAIL.n149 VTAIL.n148 104.615
R1373 VTAIL.n148 VTAIL.n81 104.615
R1374 VTAIL.n141 VTAIL.n81 104.615
R1375 VTAIL.n141 VTAIL.n140 104.615
R1376 VTAIL.n140 VTAIL.n86 104.615
R1377 VTAIL.n133 VTAIL.n86 104.615
R1378 VTAIL.n133 VTAIL.n132 104.615
R1379 VTAIL.n132 VTAIL.n90 104.615
R1380 VTAIL.n125 VTAIL.n90 104.615
R1381 VTAIL.n125 VTAIL.n124 104.615
R1382 VTAIL.n124 VTAIL.n94 104.615
R1383 VTAIL.n117 VTAIL.n94 104.615
R1384 VTAIL.n117 VTAIL.n116 104.615
R1385 VTAIL.n116 VTAIL.n98 104.615
R1386 VTAIL.n109 VTAIL.n98 104.615
R1387 VTAIL.n109 VTAIL.n108 104.615
R1388 VTAIL.n108 VTAIL.n102 104.615
R1389 VTAIL.t2 VTAIL.n257 52.3082
R1390 VTAIL.t0 VTAIL.n23 52.3082
R1391 VTAIL.t1 VTAIL.n180 52.3082
R1392 VTAIL.t3 VTAIL.n102 52.3082
R1393 VTAIL.n311 VTAIL.n310 33.155
R1394 VTAIL.n77 VTAIL.n76 33.155
R1395 VTAIL.n233 VTAIL.n232 33.155
R1396 VTAIL.n155 VTAIL.n154 33.155
R1397 VTAIL.n155 VTAIL.n77 27.9617
R1398 VTAIL.n311 VTAIL.n233 26.1858
R1399 VTAIL.n259 VTAIL.n258 15.6677
R1400 VTAIL.n25 VTAIL.n24 15.6677
R1401 VTAIL.n182 VTAIL.n181 15.6677
R1402 VTAIL.n104 VTAIL.n103 15.6677
R1403 VTAIL.n307 VTAIL.n236 13.1884
R1404 VTAIL.n73 VTAIL.n2 13.1884
R1405 VTAIL.n229 VTAIL.n158 13.1884
R1406 VTAIL.n151 VTAIL.n80 13.1884
R1407 VTAIL.n262 VTAIL.n261 12.8005
R1408 VTAIL.n303 VTAIL.n302 12.8005
R1409 VTAIL.n308 VTAIL.n234 12.8005
R1410 VTAIL.n28 VTAIL.n27 12.8005
R1411 VTAIL.n69 VTAIL.n68 12.8005
R1412 VTAIL.n74 VTAIL.n0 12.8005
R1413 VTAIL.n230 VTAIL.n156 12.8005
R1414 VTAIL.n225 VTAIL.n160 12.8005
R1415 VTAIL.n185 VTAIL.n184 12.8005
R1416 VTAIL.n152 VTAIL.n78 12.8005
R1417 VTAIL.n147 VTAIL.n82 12.8005
R1418 VTAIL.n107 VTAIL.n106 12.8005
R1419 VTAIL.n265 VTAIL.n256 12.0247
R1420 VTAIL.n301 VTAIL.n238 12.0247
R1421 VTAIL.n31 VTAIL.n22 12.0247
R1422 VTAIL.n67 VTAIL.n4 12.0247
R1423 VTAIL.n224 VTAIL.n161 12.0247
R1424 VTAIL.n188 VTAIL.n179 12.0247
R1425 VTAIL.n146 VTAIL.n83 12.0247
R1426 VTAIL.n110 VTAIL.n101 12.0247
R1427 VTAIL.n266 VTAIL.n254 11.249
R1428 VTAIL.n298 VTAIL.n297 11.249
R1429 VTAIL.n32 VTAIL.n20 11.249
R1430 VTAIL.n64 VTAIL.n63 11.249
R1431 VTAIL.n221 VTAIL.n220 11.249
R1432 VTAIL.n189 VTAIL.n177 11.249
R1433 VTAIL.n143 VTAIL.n142 11.249
R1434 VTAIL.n111 VTAIL.n99 11.249
R1435 VTAIL.n270 VTAIL.n269 10.4732
R1436 VTAIL.n294 VTAIL.n240 10.4732
R1437 VTAIL.n36 VTAIL.n35 10.4732
R1438 VTAIL.n60 VTAIL.n6 10.4732
R1439 VTAIL.n217 VTAIL.n163 10.4732
R1440 VTAIL.n193 VTAIL.n192 10.4732
R1441 VTAIL.n139 VTAIL.n85 10.4732
R1442 VTAIL.n115 VTAIL.n114 10.4732
R1443 VTAIL.n273 VTAIL.n252 9.69747
R1444 VTAIL.n293 VTAIL.n242 9.69747
R1445 VTAIL.n39 VTAIL.n18 9.69747
R1446 VTAIL.n59 VTAIL.n8 9.69747
R1447 VTAIL.n216 VTAIL.n165 9.69747
R1448 VTAIL.n196 VTAIL.n175 9.69747
R1449 VTAIL.n138 VTAIL.n87 9.69747
R1450 VTAIL.n118 VTAIL.n97 9.69747
R1451 VTAIL.n310 VTAIL.n309 9.45567
R1452 VTAIL.n76 VTAIL.n75 9.45567
R1453 VTAIL.n232 VTAIL.n231 9.45567
R1454 VTAIL.n154 VTAIL.n153 9.45567
R1455 VTAIL.n309 VTAIL.n308 9.3005
R1456 VTAIL.n248 VTAIL.n247 9.3005
R1457 VTAIL.n277 VTAIL.n276 9.3005
R1458 VTAIL.n275 VTAIL.n274 9.3005
R1459 VTAIL.n252 VTAIL.n251 9.3005
R1460 VTAIL.n269 VTAIL.n268 9.3005
R1461 VTAIL.n267 VTAIL.n266 9.3005
R1462 VTAIL.n256 VTAIL.n255 9.3005
R1463 VTAIL.n261 VTAIL.n260 9.3005
R1464 VTAIL.n283 VTAIL.n282 9.3005
R1465 VTAIL.n285 VTAIL.n284 9.3005
R1466 VTAIL.n244 VTAIL.n243 9.3005
R1467 VTAIL.n291 VTAIL.n290 9.3005
R1468 VTAIL.n293 VTAIL.n292 9.3005
R1469 VTAIL.n240 VTAIL.n239 9.3005
R1470 VTAIL.n299 VTAIL.n298 9.3005
R1471 VTAIL.n301 VTAIL.n300 9.3005
R1472 VTAIL.n302 VTAIL.n235 9.3005
R1473 VTAIL.n75 VTAIL.n74 9.3005
R1474 VTAIL.n14 VTAIL.n13 9.3005
R1475 VTAIL.n43 VTAIL.n42 9.3005
R1476 VTAIL.n41 VTAIL.n40 9.3005
R1477 VTAIL.n18 VTAIL.n17 9.3005
R1478 VTAIL.n35 VTAIL.n34 9.3005
R1479 VTAIL.n33 VTAIL.n32 9.3005
R1480 VTAIL.n22 VTAIL.n21 9.3005
R1481 VTAIL.n27 VTAIL.n26 9.3005
R1482 VTAIL.n49 VTAIL.n48 9.3005
R1483 VTAIL.n51 VTAIL.n50 9.3005
R1484 VTAIL.n10 VTAIL.n9 9.3005
R1485 VTAIL.n57 VTAIL.n56 9.3005
R1486 VTAIL.n59 VTAIL.n58 9.3005
R1487 VTAIL.n6 VTAIL.n5 9.3005
R1488 VTAIL.n65 VTAIL.n64 9.3005
R1489 VTAIL.n67 VTAIL.n66 9.3005
R1490 VTAIL.n68 VTAIL.n1 9.3005
R1491 VTAIL.n208 VTAIL.n207 9.3005
R1492 VTAIL.n167 VTAIL.n166 9.3005
R1493 VTAIL.n214 VTAIL.n213 9.3005
R1494 VTAIL.n216 VTAIL.n215 9.3005
R1495 VTAIL.n163 VTAIL.n162 9.3005
R1496 VTAIL.n222 VTAIL.n221 9.3005
R1497 VTAIL.n224 VTAIL.n223 9.3005
R1498 VTAIL.n160 VTAIL.n157 9.3005
R1499 VTAIL.n231 VTAIL.n230 9.3005
R1500 VTAIL.n206 VTAIL.n205 9.3005
R1501 VTAIL.n171 VTAIL.n170 9.3005
R1502 VTAIL.n200 VTAIL.n199 9.3005
R1503 VTAIL.n198 VTAIL.n197 9.3005
R1504 VTAIL.n175 VTAIL.n174 9.3005
R1505 VTAIL.n192 VTAIL.n191 9.3005
R1506 VTAIL.n190 VTAIL.n189 9.3005
R1507 VTAIL.n179 VTAIL.n178 9.3005
R1508 VTAIL.n184 VTAIL.n183 9.3005
R1509 VTAIL.n130 VTAIL.n129 9.3005
R1510 VTAIL.n89 VTAIL.n88 9.3005
R1511 VTAIL.n136 VTAIL.n135 9.3005
R1512 VTAIL.n138 VTAIL.n137 9.3005
R1513 VTAIL.n85 VTAIL.n84 9.3005
R1514 VTAIL.n144 VTAIL.n143 9.3005
R1515 VTAIL.n146 VTAIL.n145 9.3005
R1516 VTAIL.n82 VTAIL.n79 9.3005
R1517 VTAIL.n153 VTAIL.n152 9.3005
R1518 VTAIL.n128 VTAIL.n127 9.3005
R1519 VTAIL.n93 VTAIL.n92 9.3005
R1520 VTAIL.n122 VTAIL.n121 9.3005
R1521 VTAIL.n120 VTAIL.n119 9.3005
R1522 VTAIL.n97 VTAIL.n96 9.3005
R1523 VTAIL.n114 VTAIL.n113 9.3005
R1524 VTAIL.n112 VTAIL.n111 9.3005
R1525 VTAIL.n101 VTAIL.n100 9.3005
R1526 VTAIL.n106 VTAIL.n105 9.3005
R1527 VTAIL.n274 VTAIL.n250 8.92171
R1528 VTAIL.n290 VTAIL.n289 8.92171
R1529 VTAIL.n40 VTAIL.n16 8.92171
R1530 VTAIL.n56 VTAIL.n55 8.92171
R1531 VTAIL.n213 VTAIL.n212 8.92171
R1532 VTAIL.n197 VTAIL.n173 8.92171
R1533 VTAIL.n135 VTAIL.n134 8.92171
R1534 VTAIL.n119 VTAIL.n95 8.92171
R1535 VTAIL.n278 VTAIL.n277 8.14595
R1536 VTAIL.n286 VTAIL.n244 8.14595
R1537 VTAIL.n44 VTAIL.n43 8.14595
R1538 VTAIL.n52 VTAIL.n10 8.14595
R1539 VTAIL.n209 VTAIL.n167 8.14595
R1540 VTAIL.n201 VTAIL.n200 8.14595
R1541 VTAIL.n131 VTAIL.n89 8.14595
R1542 VTAIL.n123 VTAIL.n122 8.14595
R1543 VTAIL.n281 VTAIL.n248 7.3702
R1544 VTAIL.n285 VTAIL.n246 7.3702
R1545 VTAIL.n47 VTAIL.n14 7.3702
R1546 VTAIL.n51 VTAIL.n12 7.3702
R1547 VTAIL.n208 VTAIL.n169 7.3702
R1548 VTAIL.n204 VTAIL.n171 7.3702
R1549 VTAIL.n130 VTAIL.n91 7.3702
R1550 VTAIL.n126 VTAIL.n93 7.3702
R1551 VTAIL.n282 VTAIL.n281 6.59444
R1552 VTAIL.n282 VTAIL.n246 6.59444
R1553 VTAIL.n48 VTAIL.n47 6.59444
R1554 VTAIL.n48 VTAIL.n12 6.59444
R1555 VTAIL.n205 VTAIL.n169 6.59444
R1556 VTAIL.n205 VTAIL.n204 6.59444
R1557 VTAIL.n127 VTAIL.n91 6.59444
R1558 VTAIL.n127 VTAIL.n126 6.59444
R1559 VTAIL.n278 VTAIL.n248 5.81868
R1560 VTAIL.n286 VTAIL.n285 5.81868
R1561 VTAIL.n44 VTAIL.n14 5.81868
R1562 VTAIL.n52 VTAIL.n51 5.81868
R1563 VTAIL.n209 VTAIL.n208 5.81868
R1564 VTAIL.n201 VTAIL.n171 5.81868
R1565 VTAIL.n131 VTAIL.n130 5.81868
R1566 VTAIL.n123 VTAIL.n93 5.81868
R1567 VTAIL.n277 VTAIL.n250 5.04292
R1568 VTAIL.n289 VTAIL.n244 5.04292
R1569 VTAIL.n43 VTAIL.n16 5.04292
R1570 VTAIL.n55 VTAIL.n10 5.04292
R1571 VTAIL.n212 VTAIL.n167 5.04292
R1572 VTAIL.n200 VTAIL.n173 5.04292
R1573 VTAIL.n134 VTAIL.n89 5.04292
R1574 VTAIL.n122 VTAIL.n95 5.04292
R1575 VTAIL.n260 VTAIL.n259 4.38563
R1576 VTAIL.n26 VTAIL.n25 4.38563
R1577 VTAIL.n183 VTAIL.n182 4.38563
R1578 VTAIL.n105 VTAIL.n104 4.38563
R1579 VTAIL.n274 VTAIL.n273 4.26717
R1580 VTAIL.n290 VTAIL.n242 4.26717
R1581 VTAIL.n40 VTAIL.n39 4.26717
R1582 VTAIL.n56 VTAIL.n8 4.26717
R1583 VTAIL.n213 VTAIL.n165 4.26717
R1584 VTAIL.n197 VTAIL.n196 4.26717
R1585 VTAIL.n135 VTAIL.n87 4.26717
R1586 VTAIL.n119 VTAIL.n118 4.26717
R1587 VTAIL.n270 VTAIL.n252 3.49141
R1588 VTAIL.n294 VTAIL.n293 3.49141
R1589 VTAIL.n36 VTAIL.n18 3.49141
R1590 VTAIL.n60 VTAIL.n59 3.49141
R1591 VTAIL.n217 VTAIL.n216 3.49141
R1592 VTAIL.n193 VTAIL.n175 3.49141
R1593 VTAIL.n139 VTAIL.n138 3.49141
R1594 VTAIL.n115 VTAIL.n97 3.49141
R1595 VTAIL.n269 VTAIL.n254 2.71565
R1596 VTAIL.n297 VTAIL.n240 2.71565
R1597 VTAIL.n35 VTAIL.n20 2.71565
R1598 VTAIL.n63 VTAIL.n6 2.71565
R1599 VTAIL.n220 VTAIL.n163 2.71565
R1600 VTAIL.n192 VTAIL.n177 2.71565
R1601 VTAIL.n142 VTAIL.n85 2.71565
R1602 VTAIL.n114 VTAIL.n99 2.71565
R1603 VTAIL.n266 VTAIL.n265 1.93989
R1604 VTAIL.n298 VTAIL.n238 1.93989
R1605 VTAIL.n32 VTAIL.n31 1.93989
R1606 VTAIL.n64 VTAIL.n4 1.93989
R1607 VTAIL.n221 VTAIL.n161 1.93989
R1608 VTAIL.n189 VTAIL.n188 1.93989
R1609 VTAIL.n143 VTAIL.n83 1.93989
R1610 VTAIL.n111 VTAIL.n110 1.93989
R1611 VTAIL.n233 VTAIL.n155 1.35826
R1612 VTAIL.n262 VTAIL.n256 1.16414
R1613 VTAIL.n303 VTAIL.n301 1.16414
R1614 VTAIL.n310 VTAIL.n234 1.16414
R1615 VTAIL.n28 VTAIL.n22 1.16414
R1616 VTAIL.n69 VTAIL.n67 1.16414
R1617 VTAIL.n76 VTAIL.n0 1.16414
R1618 VTAIL.n232 VTAIL.n156 1.16414
R1619 VTAIL.n225 VTAIL.n224 1.16414
R1620 VTAIL.n185 VTAIL.n179 1.16414
R1621 VTAIL.n154 VTAIL.n78 1.16414
R1622 VTAIL.n147 VTAIL.n146 1.16414
R1623 VTAIL.n107 VTAIL.n101 1.16414
R1624 VTAIL VTAIL.n77 0.972483
R1625 VTAIL.n261 VTAIL.n258 0.388379
R1626 VTAIL.n302 VTAIL.n236 0.388379
R1627 VTAIL.n308 VTAIL.n307 0.388379
R1628 VTAIL.n27 VTAIL.n24 0.388379
R1629 VTAIL.n68 VTAIL.n2 0.388379
R1630 VTAIL.n74 VTAIL.n73 0.388379
R1631 VTAIL.n230 VTAIL.n229 0.388379
R1632 VTAIL.n160 VTAIL.n158 0.388379
R1633 VTAIL.n184 VTAIL.n181 0.388379
R1634 VTAIL.n152 VTAIL.n151 0.388379
R1635 VTAIL.n82 VTAIL.n80 0.388379
R1636 VTAIL.n106 VTAIL.n103 0.388379
R1637 VTAIL VTAIL.n311 0.386276
R1638 VTAIL.n260 VTAIL.n255 0.155672
R1639 VTAIL.n267 VTAIL.n255 0.155672
R1640 VTAIL.n268 VTAIL.n267 0.155672
R1641 VTAIL.n268 VTAIL.n251 0.155672
R1642 VTAIL.n275 VTAIL.n251 0.155672
R1643 VTAIL.n276 VTAIL.n275 0.155672
R1644 VTAIL.n276 VTAIL.n247 0.155672
R1645 VTAIL.n283 VTAIL.n247 0.155672
R1646 VTAIL.n284 VTAIL.n283 0.155672
R1647 VTAIL.n284 VTAIL.n243 0.155672
R1648 VTAIL.n291 VTAIL.n243 0.155672
R1649 VTAIL.n292 VTAIL.n291 0.155672
R1650 VTAIL.n292 VTAIL.n239 0.155672
R1651 VTAIL.n299 VTAIL.n239 0.155672
R1652 VTAIL.n300 VTAIL.n299 0.155672
R1653 VTAIL.n300 VTAIL.n235 0.155672
R1654 VTAIL.n309 VTAIL.n235 0.155672
R1655 VTAIL.n26 VTAIL.n21 0.155672
R1656 VTAIL.n33 VTAIL.n21 0.155672
R1657 VTAIL.n34 VTAIL.n33 0.155672
R1658 VTAIL.n34 VTAIL.n17 0.155672
R1659 VTAIL.n41 VTAIL.n17 0.155672
R1660 VTAIL.n42 VTAIL.n41 0.155672
R1661 VTAIL.n42 VTAIL.n13 0.155672
R1662 VTAIL.n49 VTAIL.n13 0.155672
R1663 VTAIL.n50 VTAIL.n49 0.155672
R1664 VTAIL.n50 VTAIL.n9 0.155672
R1665 VTAIL.n57 VTAIL.n9 0.155672
R1666 VTAIL.n58 VTAIL.n57 0.155672
R1667 VTAIL.n58 VTAIL.n5 0.155672
R1668 VTAIL.n65 VTAIL.n5 0.155672
R1669 VTAIL.n66 VTAIL.n65 0.155672
R1670 VTAIL.n66 VTAIL.n1 0.155672
R1671 VTAIL.n75 VTAIL.n1 0.155672
R1672 VTAIL.n231 VTAIL.n157 0.155672
R1673 VTAIL.n223 VTAIL.n157 0.155672
R1674 VTAIL.n223 VTAIL.n222 0.155672
R1675 VTAIL.n222 VTAIL.n162 0.155672
R1676 VTAIL.n215 VTAIL.n162 0.155672
R1677 VTAIL.n215 VTAIL.n214 0.155672
R1678 VTAIL.n214 VTAIL.n166 0.155672
R1679 VTAIL.n207 VTAIL.n166 0.155672
R1680 VTAIL.n207 VTAIL.n206 0.155672
R1681 VTAIL.n206 VTAIL.n170 0.155672
R1682 VTAIL.n199 VTAIL.n170 0.155672
R1683 VTAIL.n199 VTAIL.n198 0.155672
R1684 VTAIL.n198 VTAIL.n174 0.155672
R1685 VTAIL.n191 VTAIL.n174 0.155672
R1686 VTAIL.n191 VTAIL.n190 0.155672
R1687 VTAIL.n190 VTAIL.n178 0.155672
R1688 VTAIL.n183 VTAIL.n178 0.155672
R1689 VTAIL.n153 VTAIL.n79 0.155672
R1690 VTAIL.n145 VTAIL.n79 0.155672
R1691 VTAIL.n145 VTAIL.n144 0.155672
R1692 VTAIL.n144 VTAIL.n84 0.155672
R1693 VTAIL.n137 VTAIL.n84 0.155672
R1694 VTAIL.n137 VTAIL.n136 0.155672
R1695 VTAIL.n136 VTAIL.n88 0.155672
R1696 VTAIL.n129 VTAIL.n88 0.155672
R1697 VTAIL.n129 VTAIL.n128 0.155672
R1698 VTAIL.n128 VTAIL.n92 0.155672
R1699 VTAIL.n121 VTAIL.n92 0.155672
R1700 VTAIL.n121 VTAIL.n120 0.155672
R1701 VTAIL.n120 VTAIL.n96 0.155672
R1702 VTAIL.n113 VTAIL.n96 0.155672
R1703 VTAIL.n113 VTAIL.n112 0.155672
R1704 VTAIL.n112 VTAIL.n100 0.155672
R1705 VTAIL.n105 VTAIL.n100 0.155672
R1706 VDD2.n149 VDD2.n77 289.615
R1707 VDD2.n72 VDD2.n0 289.615
R1708 VDD2.n150 VDD2.n149 185
R1709 VDD2.n148 VDD2.n79 185
R1710 VDD2.n147 VDD2.n146 185
R1711 VDD2.n82 VDD2.n80 185
R1712 VDD2.n141 VDD2.n140 185
R1713 VDD2.n139 VDD2.n138 185
R1714 VDD2.n86 VDD2.n85 185
R1715 VDD2.n133 VDD2.n132 185
R1716 VDD2.n131 VDD2.n130 185
R1717 VDD2.n90 VDD2.n89 185
R1718 VDD2.n125 VDD2.n124 185
R1719 VDD2.n123 VDD2.n122 185
R1720 VDD2.n94 VDD2.n93 185
R1721 VDD2.n117 VDD2.n116 185
R1722 VDD2.n115 VDD2.n114 185
R1723 VDD2.n98 VDD2.n97 185
R1724 VDD2.n109 VDD2.n108 185
R1725 VDD2.n107 VDD2.n106 185
R1726 VDD2.n102 VDD2.n101 185
R1727 VDD2.n24 VDD2.n23 185
R1728 VDD2.n29 VDD2.n28 185
R1729 VDD2.n31 VDD2.n30 185
R1730 VDD2.n20 VDD2.n19 185
R1731 VDD2.n37 VDD2.n36 185
R1732 VDD2.n39 VDD2.n38 185
R1733 VDD2.n16 VDD2.n15 185
R1734 VDD2.n45 VDD2.n44 185
R1735 VDD2.n47 VDD2.n46 185
R1736 VDD2.n12 VDD2.n11 185
R1737 VDD2.n53 VDD2.n52 185
R1738 VDD2.n55 VDD2.n54 185
R1739 VDD2.n8 VDD2.n7 185
R1740 VDD2.n61 VDD2.n60 185
R1741 VDD2.n63 VDD2.n62 185
R1742 VDD2.n4 VDD2.n3 185
R1743 VDD2.n70 VDD2.n69 185
R1744 VDD2.n71 VDD2.n2 185
R1745 VDD2.n73 VDD2.n72 185
R1746 VDD2.n103 VDD2.t1 147.659
R1747 VDD2.n25 VDD2.t0 147.659
R1748 VDD2.n149 VDD2.n148 104.615
R1749 VDD2.n148 VDD2.n147 104.615
R1750 VDD2.n147 VDD2.n80 104.615
R1751 VDD2.n140 VDD2.n80 104.615
R1752 VDD2.n140 VDD2.n139 104.615
R1753 VDD2.n139 VDD2.n85 104.615
R1754 VDD2.n132 VDD2.n85 104.615
R1755 VDD2.n132 VDD2.n131 104.615
R1756 VDD2.n131 VDD2.n89 104.615
R1757 VDD2.n124 VDD2.n89 104.615
R1758 VDD2.n124 VDD2.n123 104.615
R1759 VDD2.n123 VDD2.n93 104.615
R1760 VDD2.n116 VDD2.n93 104.615
R1761 VDD2.n116 VDD2.n115 104.615
R1762 VDD2.n115 VDD2.n97 104.615
R1763 VDD2.n108 VDD2.n97 104.615
R1764 VDD2.n108 VDD2.n107 104.615
R1765 VDD2.n107 VDD2.n101 104.615
R1766 VDD2.n29 VDD2.n23 104.615
R1767 VDD2.n30 VDD2.n29 104.615
R1768 VDD2.n30 VDD2.n19 104.615
R1769 VDD2.n37 VDD2.n19 104.615
R1770 VDD2.n38 VDD2.n37 104.615
R1771 VDD2.n38 VDD2.n15 104.615
R1772 VDD2.n45 VDD2.n15 104.615
R1773 VDD2.n46 VDD2.n45 104.615
R1774 VDD2.n46 VDD2.n11 104.615
R1775 VDD2.n53 VDD2.n11 104.615
R1776 VDD2.n54 VDD2.n53 104.615
R1777 VDD2.n54 VDD2.n7 104.615
R1778 VDD2.n61 VDD2.n7 104.615
R1779 VDD2.n62 VDD2.n61 104.615
R1780 VDD2.n62 VDD2.n3 104.615
R1781 VDD2.n70 VDD2.n3 104.615
R1782 VDD2.n71 VDD2.n70 104.615
R1783 VDD2.n72 VDD2.n71 104.615
R1784 VDD2.n154 VDD2.n76 89.0881
R1785 VDD2.t1 VDD2.n101 52.3082
R1786 VDD2.t0 VDD2.n23 52.3082
R1787 VDD2.n154 VDD2.n153 49.8338
R1788 VDD2.n103 VDD2.n102 15.6677
R1789 VDD2.n25 VDD2.n24 15.6677
R1790 VDD2.n150 VDD2.n79 13.1884
R1791 VDD2.n73 VDD2.n2 13.1884
R1792 VDD2.n151 VDD2.n77 12.8005
R1793 VDD2.n146 VDD2.n81 12.8005
R1794 VDD2.n106 VDD2.n105 12.8005
R1795 VDD2.n28 VDD2.n27 12.8005
R1796 VDD2.n69 VDD2.n68 12.8005
R1797 VDD2.n74 VDD2.n0 12.8005
R1798 VDD2.n145 VDD2.n82 12.0247
R1799 VDD2.n109 VDD2.n100 12.0247
R1800 VDD2.n31 VDD2.n22 12.0247
R1801 VDD2.n67 VDD2.n4 12.0247
R1802 VDD2.n142 VDD2.n141 11.249
R1803 VDD2.n110 VDD2.n98 11.249
R1804 VDD2.n32 VDD2.n20 11.249
R1805 VDD2.n64 VDD2.n63 11.249
R1806 VDD2.n138 VDD2.n84 10.4732
R1807 VDD2.n114 VDD2.n113 10.4732
R1808 VDD2.n36 VDD2.n35 10.4732
R1809 VDD2.n60 VDD2.n6 10.4732
R1810 VDD2.n137 VDD2.n86 9.69747
R1811 VDD2.n117 VDD2.n96 9.69747
R1812 VDD2.n39 VDD2.n18 9.69747
R1813 VDD2.n59 VDD2.n8 9.69747
R1814 VDD2.n153 VDD2.n152 9.45567
R1815 VDD2.n76 VDD2.n75 9.45567
R1816 VDD2.n129 VDD2.n128 9.3005
R1817 VDD2.n88 VDD2.n87 9.3005
R1818 VDD2.n135 VDD2.n134 9.3005
R1819 VDD2.n137 VDD2.n136 9.3005
R1820 VDD2.n84 VDD2.n83 9.3005
R1821 VDD2.n143 VDD2.n142 9.3005
R1822 VDD2.n145 VDD2.n144 9.3005
R1823 VDD2.n81 VDD2.n78 9.3005
R1824 VDD2.n152 VDD2.n151 9.3005
R1825 VDD2.n127 VDD2.n126 9.3005
R1826 VDD2.n92 VDD2.n91 9.3005
R1827 VDD2.n121 VDD2.n120 9.3005
R1828 VDD2.n119 VDD2.n118 9.3005
R1829 VDD2.n96 VDD2.n95 9.3005
R1830 VDD2.n113 VDD2.n112 9.3005
R1831 VDD2.n111 VDD2.n110 9.3005
R1832 VDD2.n100 VDD2.n99 9.3005
R1833 VDD2.n105 VDD2.n104 9.3005
R1834 VDD2.n75 VDD2.n74 9.3005
R1835 VDD2.n14 VDD2.n13 9.3005
R1836 VDD2.n43 VDD2.n42 9.3005
R1837 VDD2.n41 VDD2.n40 9.3005
R1838 VDD2.n18 VDD2.n17 9.3005
R1839 VDD2.n35 VDD2.n34 9.3005
R1840 VDD2.n33 VDD2.n32 9.3005
R1841 VDD2.n22 VDD2.n21 9.3005
R1842 VDD2.n27 VDD2.n26 9.3005
R1843 VDD2.n49 VDD2.n48 9.3005
R1844 VDD2.n51 VDD2.n50 9.3005
R1845 VDD2.n10 VDD2.n9 9.3005
R1846 VDD2.n57 VDD2.n56 9.3005
R1847 VDD2.n59 VDD2.n58 9.3005
R1848 VDD2.n6 VDD2.n5 9.3005
R1849 VDD2.n65 VDD2.n64 9.3005
R1850 VDD2.n67 VDD2.n66 9.3005
R1851 VDD2.n68 VDD2.n1 9.3005
R1852 VDD2.n134 VDD2.n133 8.92171
R1853 VDD2.n118 VDD2.n94 8.92171
R1854 VDD2.n40 VDD2.n16 8.92171
R1855 VDD2.n56 VDD2.n55 8.92171
R1856 VDD2.n130 VDD2.n88 8.14595
R1857 VDD2.n122 VDD2.n121 8.14595
R1858 VDD2.n44 VDD2.n43 8.14595
R1859 VDD2.n52 VDD2.n10 8.14595
R1860 VDD2.n129 VDD2.n90 7.3702
R1861 VDD2.n125 VDD2.n92 7.3702
R1862 VDD2.n47 VDD2.n14 7.3702
R1863 VDD2.n51 VDD2.n12 7.3702
R1864 VDD2.n126 VDD2.n90 6.59444
R1865 VDD2.n126 VDD2.n125 6.59444
R1866 VDD2.n48 VDD2.n47 6.59444
R1867 VDD2.n48 VDD2.n12 6.59444
R1868 VDD2.n130 VDD2.n129 5.81868
R1869 VDD2.n122 VDD2.n92 5.81868
R1870 VDD2.n44 VDD2.n14 5.81868
R1871 VDD2.n52 VDD2.n51 5.81868
R1872 VDD2.n133 VDD2.n88 5.04292
R1873 VDD2.n121 VDD2.n94 5.04292
R1874 VDD2.n43 VDD2.n16 5.04292
R1875 VDD2.n55 VDD2.n10 5.04292
R1876 VDD2.n104 VDD2.n103 4.38563
R1877 VDD2.n26 VDD2.n25 4.38563
R1878 VDD2.n134 VDD2.n86 4.26717
R1879 VDD2.n118 VDD2.n117 4.26717
R1880 VDD2.n40 VDD2.n39 4.26717
R1881 VDD2.n56 VDD2.n8 4.26717
R1882 VDD2.n138 VDD2.n137 3.49141
R1883 VDD2.n114 VDD2.n96 3.49141
R1884 VDD2.n36 VDD2.n18 3.49141
R1885 VDD2.n60 VDD2.n59 3.49141
R1886 VDD2.n141 VDD2.n84 2.71565
R1887 VDD2.n113 VDD2.n98 2.71565
R1888 VDD2.n35 VDD2.n20 2.71565
R1889 VDD2.n63 VDD2.n6 2.71565
R1890 VDD2.n142 VDD2.n82 1.93989
R1891 VDD2.n110 VDD2.n109 1.93989
R1892 VDD2.n32 VDD2.n31 1.93989
R1893 VDD2.n64 VDD2.n4 1.93989
R1894 VDD2.n153 VDD2.n77 1.16414
R1895 VDD2.n146 VDD2.n145 1.16414
R1896 VDD2.n106 VDD2.n100 1.16414
R1897 VDD2.n28 VDD2.n22 1.16414
R1898 VDD2.n69 VDD2.n67 1.16414
R1899 VDD2.n76 VDD2.n0 1.16414
R1900 VDD2 VDD2.n154 0.502655
R1901 VDD2.n151 VDD2.n150 0.388379
R1902 VDD2.n81 VDD2.n79 0.388379
R1903 VDD2.n105 VDD2.n102 0.388379
R1904 VDD2.n27 VDD2.n24 0.388379
R1905 VDD2.n68 VDD2.n2 0.388379
R1906 VDD2.n74 VDD2.n73 0.388379
R1907 VDD2.n152 VDD2.n78 0.155672
R1908 VDD2.n144 VDD2.n78 0.155672
R1909 VDD2.n144 VDD2.n143 0.155672
R1910 VDD2.n143 VDD2.n83 0.155672
R1911 VDD2.n136 VDD2.n83 0.155672
R1912 VDD2.n136 VDD2.n135 0.155672
R1913 VDD2.n135 VDD2.n87 0.155672
R1914 VDD2.n128 VDD2.n87 0.155672
R1915 VDD2.n128 VDD2.n127 0.155672
R1916 VDD2.n127 VDD2.n91 0.155672
R1917 VDD2.n120 VDD2.n91 0.155672
R1918 VDD2.n120 VDD2.n119 0.155672
R1919 VDD2.n119 VDD2.n95 0.155672
R1920 VDD2.n112 VDD2.n95 0.155672
R1921 VDD2.n112 VDD2.n111 0.155672
R1922 VDD2.n111 VDD2.n99 0.155672
R1923 VDD2.n104 VDD2.n99 0.155672
R1924 VDD2.n26 VDD2.n21 0.155672
R1925 VDD2.n33 VDD2.n21 0.155672
R1926 VDD2.n34 VDD2.n33 0.155672
R1927 VDD2.n34 VDD2.n17 0.155672
R1928 VDD2.n41 VDD2.n17 0.155672
R1929 VDD2.n42 VDD2.n41 0.155672
R1930 VDD2.n42 VDD2.n13 0.155672
R1931 VDD2.n49 VDD2.n13 0.155672
R1932 VDD2.n50 VDD2.n49 0.155672
R1933 VDD2.n50 VDD2.n9 0.155672
R1934 VDD2.n57 VDD2.n9 0.155672
R1935 VDD2.n58 VDD2.n57 0.155672
R1936 VDD2.n58 VDD2.n5 0.155672
R1937 VDD2.n65 VDD2.n5 0.155672
R1938 VDD2.n66 VDD2.n65 0.155672
R1939 VDD2.n66 VDD2.n1 0.155672
R1940 VDD2.n75 VDD2.n1 0.155672
R1941 VP.n0 VP.t1 297.313
R1942 VP.n0 VP.t0 253.472
R1943 VP VP.n0 0.241678
R1944 VDD1.n72 VDD1.n0 289.615
R1945 VDD1.n149 VDD1.n77 289.615
R1946 VDD1.n73 VDD1.n72 185
R1947 VDD1.n71 VDD1.n2 185
R1948 VDD1.n70 VDD1.n69 185
R1949 VDD1.n5 VDD1.n3 185
R1950 VDD1.n64 VDD1.n63 185
R1951 VDD1.n62 VDD1.n61 185
R1952 VDD1.n9 VDD1.n8 185
R1953 VDD1.n56 VDD1.n55 185
R1954 VDD1.n54 VDD1.n53 185
R1955 VDD1.n13 VDD1.n12 185
R1956 VDD1.n48 VDD1.n47 185
R1957 VDD1.n46 VDD1.n45 185
R1958 VDD1.n17 VDD1.n16 185
R1959 VDD1.n40 VDD1.n39 185
R1960 VDD1.n38 VDD1.n37 185
R1961 VDD1.n21 VDD1.n20 185
R1962 VDD1.n32 VDD1.n31 185
R1963 VDD1.n30 VDD1.n29 185
R1964 VDD1.n25 VDD1.n24 185
R1965 VDD1.n101 VDD1.n100 185
R1966 VDD1.n106 VDD1.n105 185
R1967 VDD1.n108 VDD1.n107 185
R1968 VDD1.n97 VDD1.n96 185
R1969 VDD1.n114 VDD1.n113 185
R1970 VDD1.n116 VDD1.n115 185
R1971 VDD1.n93 VDD1.n92 185
R1972 VDD1.n122 VDD1.n121 185
R1973 VDD1.n124 VDD1.n123 185
R1974 VDD1.n89 VDD1.n88 185
R1975 VDD1.n130 VDD1.n129 185
R1976 VDD1.n132 VDD1.n131 185
R1977 VDD1.n85 VDD1.n84 185
R1978 VDD1.n138 VDD1.n137 185
R1979 VDD1.n140 VDD1.n139 185
R1980 VDD1.n81 VDD1.n80 185
R1981 VDD1.n147 VDD1.n146 185
R1982 VDD1.n148 VDD1.n79 185
R1983 VDD1.n150 VDD1.n149 185
R1984 VDD1.n26 VDD1.t0 147.659
R1985 VDD1.n102 VDD1.t1 147.659
R1986 VDD1.n72 VDD1.n71 104.615
R1987 VDD1.n71 VDD1.n70 104.615
R1988 VDD1.n70 VDD1.n3 104.615
R1989 VDD1.n63 VDD1.n3 104.615
R1990 VDD1.n63 VDD1.n62 104.615
R1991 VDD1.n62 VDD1.n8 104.615
R1992 VDD1.n55 VDD1.n8 104.615
R1993 VDD1.n55 VDD1.n54 104.615
R1994 VDD1.n54 VDD1.n12 104.615
R1995 VDD1.n47 VDD1.n12 104.615
R1996 VDD1.n47 VDD1.n46 104.615
R1997 VDD1.n46 VDD1.n16 104.615
R1998 VDD1.n39 VDD1.n16 104.615
R1999 VDD1.n39 VDD1.n38 104.615
R2000 VDD1.n38 VDD1.n20 104.615
R2001 VDD1.n31 VDD1.n20 104.615
R2002 VDD1.n31 VDD1.n30 104.615
R2003 VDD1.n30 VDD1.n24 104.615
R2004 VDD1.n106 VDD1.n100 104.615
R2005 VDD1.n107 VDD1.n106 104.615
R2006 VDD1.n107 VDD1.n96 104.615
R2007 VDD1.n114 VDD1.n96 104.615
R2008 VDD1.n115 VDD1.n114 104.615
R2009 VDD1.n115 VDD1.n92 104.615
R2010 VDD1.n122 VDD1.n92 104.615
R2011 VDD1.n123 VDD1.n122 104.615
R2012 VDD1.n123 VDD1.n88 104.615
R2013 VDD1.n130 VDD1.n88 104.615
R2014 VDD1.n131 VDD1.n130 104.615
R2015 VDD1.n131 VDD1.n84 104.615
R2016 VDD1.n138 VDD1.n84 104.615
R2017 VDD1.n139 VDD1.n138 104.615
R2018 VDD1.n139 VDD1.n80 104.615
R2019 VDD1.n147 VDD1.n80 104.615
R2020 VDD1.n148 VDD1.n147 104.615
R2021 VDD1.n149 VDD1.n148 104.615
R2022 VDD1 VDD1.n153 90.0569
R2023 VDD1.t0 VDD1.n24 52.3082
R2024 VDD1.t1 VDD1.n100 52.3082
R2025 VDD1 VDD1.n76 50.336
R2026 VDD1.n26 VDD1.n25 15.6677
R2027 VDD1.n102 VDD1.n101 15.6677
R2028 VDD1.n73 VDD1.n2 13.1884
R2029 VDD1.n150 VDD1.n79 13.1884
R2030 VDD1.n74 VDD1.n0 12.8005
R2031 VDD1.n69 VDD1.n4 12.8005
R2032 VDD1.n29 VDD1.n28 12.8005
R2033 VDD1.n105 VDD1.n104 12.8005
R2034 VDD1.n146 VDD1.n145 12.8005
R2035 VDD1.n151 VDD1.n77 12.8005
R2036 VDD1.n68 VDD1.n5 12.0247
R2037 VDD1.n32 VDD1.n23 12.0247
R2038 VDD1.n108 VDD1.n99 12.0247
R2039 VDD1.n144 VDD1.n81 12.0247
R2040 VDD1.n65 VDD1.n64 11.249
R2041 VDD1.n33 VDD1.n21 11.249
R2042 VDD1.n109 VDD1.n97 11.249
R2043 VDD1.n141 VDD1.n140 11.249
R2044 VDD1.n61 VDD1.n7 10.4732
R2045 VDD1.n37 VDD1.n36 10.4732
R2046 VDD1.n113 VDD1.n112 10.4732
R2047 VDD1.n137 VDD1.n83 10.4732
R2048 VDD1.n60 VDD1.n9 9.69747
R2049 VDD1.n40 VDD1.n19 9.69747
R2050 VDD1.n116 VDD1.n95 9.69747
R2051 VDD1.n136 VDD1.n85 9.69747
R2052 VDD1.n76 VDD1.n75 9.45567
R2053 VDD1.n153 VDD1.n152 9.45567
R2054 VDD1.n52 VDD1.n51 9.3005
R2055 VDD1.n11 VDD1.n10 9.3005
R2056 VDD1.n58 VDD1.n57 9.3005
R2057 VDD1.n60 VDD1.n59 9.3005
R2058 VDD1.n7 VDD1.n6 9.3005
R2059 VDD1.n66 VDD1.n65 9.3005
R2060 VDD1.n68 VDD1.n67 9.3005
R2061 VDD1.n4 VDD1.n1 9.3005
R2062 VDD1.n75 VDD1.n74 9.3005
R2063 VDD1.n50 VDD1.n49 9.3005
R2064 VDD1.n15 VDD1.n14 9.3005
R2065 VDD1.n44 VDD1.n43 9.3005
R2066 VDD1.n42 VDD1.n41 9.3005
R2067 VDD1.n19 VDD1.n18 9.3005
R2068 VDD1.n36 VDD1.n35 9.3005
R2069 VDD1.n34 VDD1.n33 9.3005
R2070 VDD1.n23 VDD1.n22 9.3005
R2071 VDD1.n28 VDD1.n27 9.3005
R2072 VDD1.n152 VDD1.n151 9.3005
R2073 VDD1.n91 VDD1.n90 9.3005
R2074 VDD1.n120 VDD1.n119 9.3005
R2075 VDD1.n118 VDD1.n117 9.3005
R2076 VDD1.n95 VDD1.n94 9.3005
R2077 VDD1.n112 VDD1.n111 9.3005
R2078 VDD1.n110 VDD1.n109 9.3005
R2079 VDD1.n99 VDD1.n98 9.3005
R2080 VDD1.n104 VDD1.n103 9.3005
R2081 VDD1.n126 VDD1.n125 9.3005
R2082 VDD1.n128 VDD1.n127 9.3005
R2083 VDD1.n87 VDD1.n86 9.3005
R2084 VDD1.n134 VDD1.n133 9.3005
R2085 VDD1.n136 VDD1.n135 9.3005
R2086 VDD1.n83 VDD1.n82 9.3005
R2087 VDD1.n142 VDD1.n141 9.3005
R2088 VDD1.n144 VDD1.n143 9.3005
R2089 VDD1.n145 VDD1.n78 9.3005
R2090 VDD1.n57 VDD1.n56 8.92171
R2091 VDD1.n41 VDD1.n17 8.92171
R2092 VDD1.n117 VDD1.n93 8.92171
R2093 VDD1.n133 VDD1.n132 8.92171
R2094 VDD1.n53 VDD1.n11 8.14595
R2095 VDD1.n45 VDD1.n44 8.14595
R2096 VDD1.n121 VDD1.n120 8.14595
R2097 VDD1.n129 VDD1.n87 8.14595
R2098 VDD1.n52 VDD1.n13 7.3702
R2099 VDD1.n48 VDD1.n15 7.3702
R2100 VDD1.n124 VDD1.n91 7.3702
R2101 VDD1.n128 VDD1.n89 7.3702
R2102 VDD1.n49 VDD1.n13 6.59444
R2103 VDD1.n49 VDD1.n48 6.59444
R2104 VDD1.n125 VDD1.n124 6.59444
R2105 VDD1.n125 VDD1.n89 6.59444
R2106 VDD1.n53 VDD1.n52 5.81868
R2107 VDD1.n45 VDD1.n15 5.81868
R2108 VDD1.n121 VDD1.n91 5.81868
R2109 VDD1.n129 VDD1.n128 5.81868
R2110 VDD1.n56 VDD1.n11 5.04292
R2111 VDD1.n44 VDD1.n17 5.04292
R2112 VDD1.n120 VDD1.n93 5.04292
R2113 VDD1.n132 VDD1.n87 5.04292
R2114 VDD1.n27 VDD1.n26 4.38563
R2115 VDD1.n103 VDD1.n102 4.38563
R2116 VDD1.n57 VDD1.n9 4.26717
R2117 VDD1.n41 VDD1.n40 4.26717
R2118 VDD1.n117 VDD1.n116 4.26717
R2119 VDD1.n133 VDD1.n85 4.26717
R2120 VDD1.n61 VDD1.n60 3.49141
R2121 VDD1.n37 VDD1.n19 3.49141
R2122 VDD1.n113 VDD1.n95 3.49141
R2123 VDD1.n137 VDD1.n136 3.49141
R2124 VDD1.n64 VDD1.n7 2.71565
R2125 VDD1.n36 VDD1.n21 2.71565
R2126 VDD1.n112 VDD1.n97 2.71565
R2127 VDD1.n140 VDD1.n83 2.71565
R2128 VDD1.n65 VDD1.n5 1.93989
R2129 VDD1.n33 VDD1.n32 1.93989
R2130 VDD1.n109 VDD1.n108 1.93989
R2131 VDD1.n141 VDD1.n81 1.93989
R2132 VDD1.n76 VDD1.n0 1.16414
R2133 VDD1.n69 VDD1.n68 1.16414
R2134 VDD1.n29 VDD1.n23 1.16414
R2135 VDD1.n105 VDD1.n99 1.16414
R2136 VDD1.n146 VDD1.n144 1.16414
R2137 VDD1.n153 VDD1.n77 1.16414
R2138 VDD1.n74 VDD1.n73 0.388379
R2139 VDD1.n4 VDD1.n2 0.388379
R2140 VDD1.n28 VDD1.n25 0.388379
R2141 VDD1.n104 VDD1.n101 0.388379
R2142 VDD1.n145 VDD1.n79 0.388379
R2143 VDD1.n151 VDD1.n150 0.388379
R2144 VDD1.n75 VDD1.n1 0.155672
R2145 VDD1.n67 VDD1.n1 0.155672
R2146 VDD1.n67 VDD1.n66 0.155672
R2147 VDD1.n66 VDD1.n6 0.155672
R2148 VDD1.n59 VDD1.n6 0.155672
R2149 VDD1.n59 VDD1.n58 0.155672
R2150 VDD1.n58 VDD1.n10 0.155672
R2151 VDD1.n51 VDD1.n10 0.155672
R2152 VDD1.n51 VDD1.n50 0.155672
R2153 VDD1.n50 VDD1.n14 0.155672
R2154 VDD1.n43 VDD1.n14 0.155672
R2155 VDD1.n43 VDD1.n42 0.155672
R2156 VDD1.n42 VDD1.n18 0.155672
R2157 VDD1.n35 VDD1.n18 0.155672
R2158 VDD1.n35 VDD1.n34 0.155672
R2159 VDD1.n34 VDD1.n22 0.155672
R2160 VDD1.n27 VDD1.n22 0.155672
R2161 VDD1.n103 VDD1.n98 0.155672
R2162 VDD1.n110 VDD1.n98 0.155672
R2163 VDD1.n111 VDD1.n110 0.155672
R2164 VDD1.n111 VDD1.n94 0.155672
R2165 VDD1.n118 VDD1.n94 0.155672
R2166 VDD1.n119 VDD1.n118 0.155672
R2167 VDD1.n119 VDD1.n90 0.155672
R2168 VDD1.n126 VDD1.n90 0.155672
R2169 VDD1.n127 VDD1.n126 0.155672
R2170 VDD1.n127 VDD1.n86 0.155672
R2171 VDD1.n134 VDD1.n86 0.155672
R2172 VDD1.n135 VDD1.n134 0.155672
R2173 VDD1.n135 VDD1.n82 0.155672
R2174 VDD1.n142 VDD1.n82 0.155672
R2175 VDD1.n143 VDD1.n142 0.155672
R2176 VDD1.n143 VDD1.n78 0.155672
R2177 VDD1.n152 VDD1.n78 0.155672
C0 VDD1 VP 3.10969f
C1 VP VDD2 0.296812f
C2 VN VP 5.41431f
C3 VDD1 VTAIL 5.59491f
C4 VTAIL VDD2 5.63781f
C5 VTAIL VN 2.48417f
C6 VTAIL VP 2.49859f
C7 VDD1 VDD2 0.572513f
C8 VDD1 VN 0.147723f
C9 VN VDD2 2.96417f
C10 VDD2 B 4.479456f
C11 VDD1 B 7.19328f
C12 VTAIL B 7.700065f
C13 VN B 10.440551f
C14 VP B 5.457789f
C15 VDD1.n0 B 0.025743f
C16 VDD1.n1 B 0.020152f
C17 VDD1.n2 B 0.011148f
C18 VDD1.n3 B 0.025596f
C19 VDD1.n4 B 0.010829f
C20 VDD1.n5 B 0.011466f
C21 VDD1.n6 B 0.020152f
C22 VDD1.n7 B 0.010829f
C23 VDD1.n8 B 0.025596f
C24 VDD1.n9 B 0.011466f
C25 VDD1.n10 B 0.020152f
C26 VDD1.n11 B 0.010829f
C27 VDD1.n12 B 0.025596f
C28 VDD1.n13 B 0.011466f
C29 VDD1.n14 B 0.020152f
C30 VDD1.n15 B 0.010829f
C31 VDD1.n16 B 0.025596f
C32 VDD1.n17 B 0.011466f
C33 VDD1.n18 B 0.020152f
C34 VDD1.n19 B 0.010829f
C35 VDD1.n20 B 0.025596f
C36 VDD1.n21 B 0.011466f
C37 VDD1.n22 B 0.020152f
C38 VDD1.n23 B 0.010829f
C39 VDD1.n24 B 0.019197f
C40 VDD1.n25 B 0.01512f
C41 VDD1.t0 B 0.042133f
C42 VDD1.n26 B 0.126233f
C43 VDD1.n27 B 1.21601f
C44 VDD1.n28 B 0.010829f
C45 VDD1.n29 B 0.011466f
C46 VDD1.n30 B 0.025596f
C47 VDD1.n31 B 0.025596f
C48 VDD1.n32 B 0.011466f
C49 VDD1.n33 B 0.010829f
C50 VDD1.n34 B 0.020152f
C51 VDD1.n35 B 0.020152f
C52 VDD1.n36 B 0.010829f
C53 VDD1.n37 B 0.011466f
C54 VDD1.n38 B 0.025596f
C55 VDD1.n39 B 0.025596f
C56 VDD1.n40 B 0.011466f
C57 VDD1.n41 B 0.010829f
C58 VDD1.n42 B 0.020152f
C59 VDD1.n43 B 0.020152f
C60 VDD1.n44 B 0.010829f
C61 VDD1.n45 B 0.011466f
C62 VDD1.n46 B 0.025596f
C63 VDD1.n47 B 0.025596f
C64 VDD1.n48 B 0.011466f
C65 VDD1.n49 B 0.010829f
C66 VDD1.n50 B 0.020152f
C67 VDD1.n51 B 0.020152f
C68 VDD1.n52 B 0.010829f
C69 VDD1.n53 B 0.011466f
C70 VDD1.n54 B 0.025596f
C71 VDD1.n55 B 0.025596f
C72 VDD1.n56 B 0.011466f
C73 VDD1.n57 B 0.010829f
C74 VDD1.n58 B 0.020152f
C75 VDD1.n59 B 0.020152f
C76 VDD1.n60 B 0.010829f
C77 VDD1.n61 B 0.011466f
C78 VDD1.n62 B 0.025596f
C79 VDD1.n63 B 0.025596f
C80 VDD1.n64 B 0.011466f
C81 VDD1.n65 B 0.010829f
C82 VDD1.n66 B 0.020152f
C83 VDD1.n67 B 0.020152f
C84 VDD1.n68 B 0.010829f
C85 VDD1.n69 B 0.011466f
C86 VDD1.n70 B 0.025596f
C87 VDD1.n71 B 0.025596f
C88 VDD1.n72 B 0.050842f
C89 VDD1.n73 B 0.011148f
C90 VDD1.n74 B 0.010829f
C91 VDD1.n75 B 0.047957f
C92 VDD1.n76 B 0.042645f
C93 VDD1.n77 B 0.025743f
C94 VDD1.n78 B 0.020152f
C95 VDD1.n79 B 0.011148f
C96 VDD1.n80 B 0.025596f
C97 VDD1.n81 B 0.011466f
C98 VDD1.n82 B 0.020152f
C99 VDD1.n83 B 0.010829f
C100 VDD1.n84 B 0.025596f
C101 VDD1.n85 B 0.011466f
C102 VDD1.n86 B 0.020152f
C103 VDD1.n87 B 0.010829f
C104 VDD1.n88 B 0.025596f
C105 VDD1.n89 B 0.011466f
C106 VDD1.n90 B 0.020152f
C107 VDD1.n91 B 0.010829f
C108 VDD1.n92 B 0.025596f
C109 VDD1.n93 B 0.011466f
C110 VDD1.n94 B 0.020152f
C111 VDD1.n95 B 0.010829f
C112 VDD1.n96 B 0.025596f
C113 VDD1.n97 B 0.011466f
C114 VDD1.n98 B 0.020152f
C115 VDD1.n99 B 0.010829f
C116 VDD1.n100 B 0.019197f
C117 VDD1.n101 B 0.01512f
C118 VDD1.t1 B 0.042133f
C119 VDD1.n102 B 0.126233f
C120 VDD1.n103 B 1.21601f
C121 VDD1.n104 B 0.010829f
C122 VDD1.n105 B 0.011466f
C123 VDD1.n106 B 0.025596f
C124 VDD1.n107 B 0.025596f
C125 VDD1.n108 B 0.011466f
C126 VDD1.n109 B 0.010829f
C127 VDD1.n110 B 0.020152f
C128 VDD1.n111 B 0.020152f
C129 VDD1.n112 B 0.010829f
C130 VDD1.n113 B 0.011466f
C131 VDD1.n114 B 0.025596f
C132 VDD1.n115 B 0.025596f
C133 VDD1.n116 B 0.011466f
C134 VDD1.n117 B 0.010829f
C135 VDD1.n118 B 0.020152f
C136 VDD1.n119 B 0.020152f
C137 VDD1.n120 B 0.010829f
C138 VDD1.n121 B 0.011466f
C139 VDD1.n122 B 0.025596f
C140 VDD1.n123 B 0.025596f
C141 VDD1.n124 B 0.011466f
C142 VDD1.n125 B 0.010829f
C143 VDD1.n126 B 0.020152f
C144 VDD1.n127 B 0.020152f
C145 VDD1.n128 B 0.010829f
C146 VDD1.n129 B 0.011466f
C147 VDD1.n130 B 0.025596f
C148 VDD1.n131 B 0.025596f
C149 VDD1.n132 B 0.011466f
C150 VDD1.n133 B 0.010829f
C151 VDD1.n134 B 0.020152f
C152 VDD1.n135 B 0.020152f
C153 VDD1.n136 B 0.010829f
C154 VDD1.n137 B 0.011466f
C155 VDD1.n138 B 0.025596f
C156 VDD1.n139 B 0.025596f
C157 VDD1.n140 B 0.011466f
C158 VDD1.n141 B 0.010829f
C159 VDD1.n142 B 0.020152f
C160 VDD1.n143 B 0.020152f
C161 VDD1.n144 B 0.010829f
C162 VDD1.n145 B 0.010829f
C163 VDD1.n146 B 0.011466f
C164 VDD1.n147 B 0.025596f
C165 VDD1.n148 B 0.025596f
C166 VDD1.n149 B 0.050842f
C167 VDD1.n150 B 0.011148f
C168 VDD1.n151 B 0.010829f
C169 VDD1.n152 B 0.047957f
C170 VDD1.n153 B 0.62859f
C171 VP.t1 B 3.22064f
C172 VP.t0 B 2.82914f
C173 VP.n0 B 4.89319f
C174 VDD2.n0 B 0.025666f
C175 VDD2.n1 B 0.020093f
C176 VDD2.n2 B 0.011114f
C177 VDD2.n3 B 0.02552f
C178 VDD2.n4 B 0.011432f
C179 VDD2.n5 B 0.020093f
C180 VDD2.n6 B 0.010797f
C181 VDD2.n7 B 0.02552f
C182 VDD2.n8 B 0.011432f
C183 VDD2.n9 B 0.020093f
C184 VDD2.n10 B 0.010797f
C185 VDD2.n11 B 0.02552f
C186 VDD2.n12 B 0.011432f
C187 VDD2.n13 B 0.020093f
C188 VDD2.n14 B 0.010797f
C189 VDD2.n15 B 0.02552f
C190 VDD2.n16 B 0.011432f
C191 VDD2.n17 B 0.020093f
C192 VDD2.n18 B 0.010797f
C193 VDD2.n19 B 0.02552f
C194 VDD2.n20 B 0.011432f
C195 VDD2.n21 B 0.020093f
C196 VDD2.n22 B 0.010797f
C197 VDD2.n23 B 0.01914f
C198 VDD2.n24 B 0.015075f
C199 VDD2.t0 B 0.042008f
C200 VDD2.n25 B 0.125859f
C201 VDD2.n26 B 1.2124f
C202 VDD2.n27 B 0.010797f
C203 VDD2.n28 B 0.011432f
C204 VDD2.n29 B 0.02552f
C205 VDD2.n30 B 0.02552f
C206 VDD2.n31 B 0.011432f
C207 VDD2.n32 B 0.010797f
C208 VDD2.n33 B 0.020093f
C209 VDD2.n34 B 0.020093f
C210 VDD2.n35 B 0.010797f
C211 VDD2.n36 B 0.011432f
C212 VDD2.n37 B 0.02552f
C213 VDD2.n38 B 0.02552f
C214 VDD2.n39 B 0.011432f
C215 VDD2.n40 B 0.010797f
C216 VDD2.n41 B 0.020093f
C217 VDD2.n42 B 0.020093f
C218 VDD2.n43 B 0.010797f
C219 VDD2.n44 B 0.011432f
C220 VDD2.n45 B 0.02552f
C221 VDD2.n46 B 0.02552f
C222 VDD2.n47 B 0.011432f
C223 VDD2.n48 B 0.010797f
C224 VDD2.n49 B 0.020093f
C225 VDD2.n50 B 0.020093f
C226 VDD2.n51 B 0.010797f
C227 VDD2.n52 B 0.011432f
C228 VDD2.n53 B 0.02552f
C229 VDD2.n54 B 0.02552f
C230 VDD2.n55 B 0.011432f
C231 VDD2.n56 B 0.010797f
C232 VDD2.n57 B 0.020093f
C233 VDD2.n58 B 0.020093f
C234 VDD2.n59 B 0.010797f
C235 VDD2.n60 B 0.011432f
C236 VDD2.n61 B 0.02552f
C237 VDD2.n62 B 0.02552f
C238 VDD2.n63 B 0.011432f
C239 VDD2.n64 B 0.010797f
C240 VDD2.n65 B 0.020093f
C241 VDD2.n66 B 0.020093f
C242 VDD2.n67 B 0.010797f
C243 VDD2.n68 B 0.010797f
C244 VDD2.n69 B 0.011432f
C245 VDD2.n70 B 0.02552f
C246 VDD2.n71 B 0.02552f
C247 VDD2.n72 B 0.050691f
C248 VDD2.n73 B 0.011114f
C249 VDD2.n74 B 0.010797f
C250 VDD2.n75 B 0.047815f
C251 VDD2.n76 B 0.592472f
C252 VDD2.n77 B 0.025666f
C253 VDD2.n78 B 0.020093f
C254 VDD2.n79 B 0.011114f
C255 VDD2.n80 B 0.02552f
C256 VDD2.n81 B 0.010797f
C257 VDD2.n82 B 0.011432f
C258 VDD2.n83 B 0.020093f
C259 VDD2.n84 B 0.010797f
C260 VDD2.n85 B 0.02552f
C261 VDD2.n86 B 0.011432f
C262 VDD2.n87 B 0.020093f
C263 VDD2.n88 B 0.010797f
C264 VDD2.n89 B 0.02552f
C265 VDD2.n90 B 0.011432f
C266 VDD2.n91 B 0.020093f
C267 VDD2.n92 B 0.010797f
C268 VDD2.n93 B 0.02552f
C269 VDD2.n94 B 0.011432f
C270 VDD2.n95 B 0.020093f
C271 VDD2.n96 B 0.010797f
C272 VDD2.n97 B 0.02552f
C273 VDD2.n98 B 0.011432f
C274 VDD2.n99 B 0.020093f
C275 VDD2.n100 B 0.010797f
C276 VDD2.n101 B 0.01914f
C277 VDD2.n102 B 0.015075f
C278 VDD2.t1 B 0.042008f
C279 VDD2.n103 B 0.125859f
C280 VDD2.n104 B 1.2124f
C281 VDD2.n105 B 0.010797f
C282 VDD2.n106 B 0.011432f
C283 VDD2.n107 B 0.02552f
C284 VDD2.n108 B 0.02552f
C285 VDD2.n109 B 0.011432f
C286 VDD2.n110 B 0.010797f
C287 VDD2.n111 B 0.020093f
C288 VDD2.n112 B 0.020093f
C289 VDD2.n113 B 0.010797f
C290 VDD2.n114 B 0.011432f
C291 VDD2.n115 B 0.02552f
C292 VDD2.n116 B 0.02552f
C293 VDD2.n117 B 0.011432f
C294 VDD2.n118 B 0.010797f
C295 VDD2.n119 B 0.020093f
C296 VDD2.n120 B 0.020093f
C297 VDD2.n121 B 0.010797f
C298 VDD2.n122 B 0.011432f
C299 VDD2.n123 B 0.02552f
C300 VDD2.n124 B 0.02552f
C301 VDD2.n125 B 0.011432f
C302 VDD2.n126 B 0.010797f
C303 VDD2.n127 B 0.020093f
C304 VDD2.n128 B 0.020093f
C305 VDD2.n129 B 0.010797f
C306 VDD2.n130 B 0.011432f
C307 VDD2.n131 B 0.02552f
C308 VDD2.n132 B 0.02552f
C309 VDD2.n133 B 0.011432f
C310 VDD2.n134 B 0.010797f
C311 VDD2.n135 B 0.020093f
C312 VDD2.n136 B 0.020093f
C313 VDD2.n137 B 0.010797f
C314 VDD2.n138 B 0.011432f
C315 VDD2.n139 B 0.02552f
C316 VDD2.n140 B 0.02552f
C317 VDD2.n141 B 0.011432f
C318 VDD2.n142 B 0.010797f
C319 VDD2.n143 B 0.020093f
C320 VDD2.n144 B 0.020093f
C321 VDD2.n145 B 0.010797f
C322 VDD2.n146 B 0.011432f
C323 VDD2.n147 B 0.02552f
C324 VDD2.n148 B 0.02552f
C325 VDD2.n149 B 0.050691f
C326 VDD2.n150 B 0.011114f
C327 VDD2.n151 B 0.010797f
C328 VDD2.n152 B 0.047815f
C329 VDD2.n153 B 0.0418f
C330 VDD2.n154 B 2.48825f
C331 VTAIL.n0 B 0.025651f
C332 VTAIL.n1 B 0.020081f
C333 VTAIL.n2 B 0.011108f
C334 VTAIL.n3 B 0.025505f
C335 VTAIL.n4 B 0.011425f
C336 VTAIL.n5 B 0.020081f
C337 VTAIL.n6 B 0.010791f
C338 VTAIL.n7 B 0.025505f
C339 VTAIL.n8 B 0.011425f
C340 VTAIL.n9 B 0.020081f
C341 VTAIL.n10 B 0.010791f
C342 VTAIL.n11 B 0.025505f
C343 VTAIL.n12 B 0.011425f
C344 VTAIL.n13 B 0.020081f
C345 VTAIL.n14 B 0.010791f
C346 VTAIL.n15 B 0.025505f
C347 VTAIL.n16 B 0.011425f
C348 VTAIL.n17 B 0.020081f
C349 VTAIL.n18 B 0.010791f
C350 VTAIL.n19 B 0.025505f
C351 VTAIL.n20 B 0.011425f
C352 VTAIL.n21 B 0.020081f
C353 VTAIL.n22 B 0.010791f
C354 VTAIL.n23 B 0.019129f
C355 VTAIL.n24 B 0.015067f
C356 VTAIL.t0 B 0.041984f
C357 VTAIL.n25 B 0.125787f
C358 VTAIL.n26 B 1.2117f
C359 VTAIL.n27 B 0.010791f
C360 VTAIL.n28 B 0.011425f
C361 VTAIL.n29 B 0.025505f
C362 VTAIL.n30 B 0.025505f
C363 VTAIL.n31 B 0.011425f
C364 VTAIL.n32 B 0.010791f
C365 VTAIL.n33 B 0.020081f
C366 VTAIL.n34 B 0.020081f
C367 VTAIL.n35 B 0.010791f
C368 VTAIL.n36 B 0.011425f
C369 VTAIL.n37 B 0.025505f
C370 VTAIL.n38 B 0.025505f
C371 VTAIL.n39 B 0.011425f
C372 VTAIL.n40 B 0.010791f
C373 VTAIL.n41 B 0.020081f
C374 VTAIL.n42 B 0.020081f
C375 VTAIL.n43 B 0.010791f
C376 VTAIL.n44 B 0.011425f
C377 VTAIL.n45 B 0.025505f
C378 VTAIL.n46 B 0.025505f
C379 VTAIL.n47 B 0.011425f
C380 VTAIL.n48 B 0.010791f
C381 VTAIL.n49 B 0.020081f
C382 VTAIL.n50 B 0.020081f
C383 VTAIL.n51 B 0.010791f
C384 VTAIL.n52 B 0.011425f
C385 VTAIL.n53 B 0.025505f
C386 VTAIL.n54 B 0.025505f
C387 VTAIL.n55 B 0.011425f
C388 VTAIL.n56 B 0.010791f
C389 VTAIL.n57 B 0.020081f
C390 VTAIL.n58 B 0.020081f
C391 VTAIL.n59 B 0.010791f
C392 VTAIL.n60 B 0.011425f
C393 VTAIL.n61 B 0.025505f
C394 VTAIL.n62 B 0.025505f
C395 VTAIL.n63 B 0.011425f
C396 VTAIL.n64 B 0.010791f
C397 VTAIL.n65 B 0.020081f
C398 VTAIL.n66 B 0.020081f
C399 VTAIL.n67 B 0.010791f
C400 VTAIL.n68 B 0.010791f
C401 VTAIL.n69 B 0.011425f
C402 VTAIL.n70 B 0.025505f
C403 VTAIL.n71 B 0.025505f
C404 VTAIL.n72 B 0.050662f
C405 VTAIL.n73 B 0.011108f
C406 VTAIL.n74 B 0.010791f
C407 VTAIL.n75 B 0.047788f
C408 VTAIL.n76 B 0.027921f
C409 VTAIL.n77 B 1.36266f
C410 VTAIL.n78 B 0.025651f
C411 VTAIL.n79 B 0.020081f
C412 VTAIL.n80 B 0.011108f
C413 VTAIL.n81 B 0.025505f
C414 VTAIL.n82 B 0.010791f
C415 VTAIL.n83 B 0.011425f
C416 VTAIL.n84 B 0.020081f
C417 VTAIL.n85 B 0.010791f
C418 VTAIL.n86 B 0.025505f
C419 VTAIL.n87 B 0.011425f
C420 VTAIL.n88 B 0.020081f
C421 VTAIL.n89 B 0.010791f
C422 VTAIL.n90 B 0.025505f
C423 VTAIL.n91 B 0.011425f
C424 VTAIL.n92 B 0.020081f
C425 VTAIL.n93 B 0.010791f
C426 VTAIL.n94 B 0.025505f
C427 VTAIL.n95 B 0.011425f
C428 VTAIL.n96 B 0.020081f
C429 VTAIL.n97 B 0.010791f
C430 VTAIL.n98 B 0.025505f
C431 VTAIL.n99 B 0.011425f
C432 VTAIL.n100 B 0.020081f
C433 VTAIL.n101 B 0.010791f
C434 VTAIL.n102 B 0.019129f
C435 VTAIL.n103 B 0.015067f
C436 VTAIL.t3 B 0.041984f
C437 VTAIL.n104 B 0.125787f
C438 VTAIL.n105 B 1.2117f
C439 VTAIL.n106 B 0.010791f
C440 VTAIL.n107 B 0.011425f
C441 VTAIL.n108 B 0.025505f
C442 VTAIL.n109 B 0.025505f
C443 VTAIL.n110 B 0.011425f
C444 VTAIL.n111 B 0.010791f
C445 VTAIL.n112 B 0.020081f
C446 VTAIL.n113 B 0.020081f
C447 VTAIL.n114 B 0.010791f
C448 VTAIL.n115 B 0.011425f
C449 VTAIL.n116 B 0.025505f
C450 VTAIL.n117 B 0.025505f
C451 VTAIL.n118 B 0.011425f
C452 VTAIL.n119 B 0.010791f
C453 VTAIL.n120 B 0.020081f
C454 VTAIL.n121 B 0.020081f
C455 VTAIL.n122 B 0.010791f
C456 VTAIL.n123 B 0.011425f
C457 VTAIL.n124 B 0.025505f
C458 VTAIL.n125 B 0.025505f
C459 VTAIL.n126 B 0.011425f
C460 VTAIL.n127 B 0.010791f
C461 VTAIL.n128 B 0.020081f
C462 VTAIL.n129 B 0.020081f
C463 VTAIL.n130 B 0.010791f
C464 VTAIL.n131 B 0.011425f
C465 VTAIL.n132 B 0.025505f
C466 VTAIL.n133 B 0.025505f
C467 VTAIL.n134 B 0.011425f
C468 VTAIL.n135 B 0.010791f
C469 VTAIL.n136 B 0.020081f
C470 VTAIL.n137 B 0.020081f
C471 VTAIL.n138 B 0.010791f
C472 VTAIL.n139 B 0.011425f
C473 VTAIL.n140 B 0.025505f
C474 VTAIL.n141 B 0.025505f
C475 VTAIL.n142 B 0.011425f
C476 VTAIL.n143 B 0.010791f
C477 VTAIL.n144 B 0.020081f
C478 VTAIL.n145 B 0.020081f
C479 VTAIL.n146 B 0.010791f
C480 VTAIL.n147 B 0.011425f
C481 VTAIL.n148 B 0.025505f
C482 VTAIL.n149 B 0.025505f
C483 VTAIL.n150 B 0.050662f
C484 VTAIL.n151 B 0.011108f
C485 VTAIL.n152 B 0.010791f
C486 VTAIL.n153 B 0.047788f
C487 VTAIL.n154 B 0.027921f
C488 VTAIL.n155 B 1.38762f
C489 VTAIL.n156 B 0.025651f
C490 VTAIL.n157 B 0.020081f
C491 VTAIL.n158 B 0.011108f
C492 VTAIL.n159 B 0.025505f
C493 VTAIL.n160 B 0.010791f
C494 VTAIL.n161 B 0.011425f
C495 VTAIL.n162 B 0.020081f
C496 VTAIL.n163 B 0.010791f
C497 VTAIL.n164 B 0.025505f
C498 VTAIL.n165 B 0.011425f
C499 VTAIL.n166 B 0.020081f
C500 VTAIL.n167 B 0.010791f
C501 VTAIL.n168 B 0.025505f
C502 VTAIL.n169 B 0.011425f
C503 VTAIL.n170 B 0.020081f
C504 VTAIL.n171 B 0.010791f
C505 VTAIL.n172 B 0.025505f
C506 VTAIL.n173 B 0.011425f
C507 VTAIL.n174 B 0.020081f
C508 VTAIL.n175 B 0.010791f
C509 VTAIL.n176 B 0.025505f
C510 VTAIL.n177 B 0.011425f
C511 VTAIL.n178 B 0.020081f
C512 VTAIL.n179 B 0.010791f
C513 VTAIL.n180 B 0.019129f
C514 VTAIL.n181 B 0.015067f
C515 VTAIL.t1 B 0.041984f
C516 VTAIL.n182 B 0.125787f
C517 VTAIL.n183 B 1.2117f
C518 VTAIL.n184 B 0.010791f
C519 VTAIL.n185 B 0.011425f
C520 VTAIL.n186 B 0.025505f
C521 VTAIL.n187 B 0.025505f
C522 VTAIL.n188 B 0.011425f
C523 VTAIL.n189 B 0.010791f
C524 VTAIL.n190 B 0.020081f
C525 VTAIL.n191 B 0.020081f
C526 VTAIL.n192 B 0.010791f
C527 VTAIL.n193 B 0.011425f
C528 VTAIL.n194 B 0.025505f
C529 VTAIL.n195 B 0.025505f
C530 VTAIL.n196 B 0.011425f
C531 VTAIL.n197 B 0.010791f
C532 VTAIL.n198 B 0.020081f
C533 VTAIL.n199 B 0.020081f
C534 VTAIL.n200 B 0.010791f
C535 VTAIL.n201 B 0.011425f
C536 VTAIL.n202 B 0.025505f
C537 VTAIL.n203 B 0.025505f
C538 VTAIL.n204 B 0.011425f
C539 VTAIL.n205 B 0.010791f
C540 VTAIL.n206 B 0.020081f
C541 VTAIL.n207 B 0.020081f
C542 VTAIL.n208 B 0.010791f
C543 VTAIL.n209 B 0.011425f
C544 VTAIL.n210 B 0.025505f
C545 VTAIL.n211 B 0.025505f
C546 VTAIL.n212 B 0.011425f
C547 VTAIL.n213 B 0.010791f
C548 VTAIL.n214 B 0.020081f
C549 VTAIL.n215 B 0.020081f
C550 VTAIL.n216 B 0.010791f
C551 VTAIL.n217 B 0.011425f
C552 VTAIL.n218 B 0.025505f
C553 VTAIL.n219 B 0.025505f
C554 VTAIL.n220 B 0.011425f
C555 VTAIL.n221 B 0.010791f
C556 VTAIL.n222 B 0.020081f
C557 VTAIL.n223 B 0.020081f
C558 VTAIL.n224 B 0.010791f
C559 VTAIL.n225 B 0.011425f
C560 VTAIL.n226 B 0.025505f
C561 VTAIL.n227 B 0.025505f
C562 VTAIL.n228 B 0.050662f
C563 VTAIL.n229 B 0.011108f
C564 VTAIL.n230 B 0.010791f
C565 VTAIL.n231 B 0.047788f
C566 VTAIL.n232 B 0.027921f
C567 VTAIL.n233 B 1.27272f
C568 VTAIL.n234 B 0.025651f
C569 VTAIL.n235 B 0.020081f
C570 VTAIL.n236 B 0.011108f
C571 VTAIL.n237 B 0.025505f
C572 VTAIL.n238 B 0.011425f
C573 VTAIL.n239 B 0.020081f
C574 VTAIL.n240 B 0.010791f
C575 VTAIL.n241 B 0.025505f
C576 VTAIL.n242 B 0.011425f
C577 VTAIL.n243 B 0.020081f
C578 VTAIL.n244 B 0.010791f
C579 VTAIL.n245 B 0.025505f
C580 VTAIL.n246 B 0.011425f
C581 VTAIL.n247 B 0.020081f
C582 VTAIL.n248 B 0.010791f
C583 VTAIL.n249 B 0.025505f
C584 VTAIL.n250 B 0.011425f
C585 VTAIL.n251 B 0.020081f
C586 VTAIL.n252 B 0.010791f
C587 VTAIL.n253 B 0.025505f
C588 VTAIL.n254 B 0.011425f
C589 VTAIL.n255 B 0.020081f
C590 VTAIL.n256 B 0.010791f
C591 VTAIL.n257 B 0.019129f
C592 VTAIL.n258 B 0.015067f
C593 VTAIL.t2 B 0.041984f
C594 VTAIL.n259 B 0.125787f
C595 VTAIL.n260 B 1.2117f
C596 VTAIL.n261 B 0.010791f
C597 VTAIL.n262 B 0.011425f
C598 VTAIL.n263 B 0.025505f
C599 VTAIL.n264 B 0.025505f
C600 VTAIL.n265 B 0.011425f
C601 VTAIL.n266 B 0.010791f
C602 VTAIL.n267 B 0.020081f
C603 VTAIL.n268 B 0.020081f
C604 VTAIL.n269 B 0.010791f
C605 VTAIL.n270 B 0.011425f
C606 VTAIL.n271 B 0.025505f
C607 VTAIL.n272 B 0.025505f
C608 VTAIL.n273 B 0.011425f
C609 VTAIL.n274 B 0.010791f
C610 VTAIL.n275 B 0.020081f
C611 VTAIL.n276 B 0.020081f
C612 VTAIL.n277 B 0.010791f
C613 VTAIL.n278 B 0.011425f
C614 VTAIL.n279 B 0.025505f
C615 VTAIL.n280 B 0.025505f
C616 VTAIL.n281 B 0.011425f
C617 VTAIL.n282 B 0.010791f
C618 VTAIL.n283 B 0.020081f
C619 VTAIL.n284 B 0.020081f
C620 VTAIL.n285 B 0.010791f
C621 VTAIL.n286 B 0.011425f
C622 VTAIL.n287 B 0.025505f
C623 VTAIL.n288 B 0.025505f
C624 VTAIL.n289 B 0.011425f
C625 VTAIL.n290 B 0.010791f
C626 VTAIL.n291 B 0.020081f
C627 VTAIL.n292 B 0.020081f
C628 VTAIL.n293 B 0.010791f
C629 VTAIL.n294 B 0.011425f
C630 VTAIL.n295 B 0.025505f
C631 VTAIL.n296 B 0.025505f
C632 VTAIL.n297 B 0.011425f
C633 VTAIL.n298 B 0.010791f
C634 VTAIL.n299 B 0.020081f
C635 VTAIL.n300 B 0.020081f
C636 VTAIL.n301 B 0.010791f
C637 VTAIL.n302 B 0.010791f
C638 VTAIL.n303 B 0.011425f
C639 VTAIL.n304 B 0.025505f
C640 VTAIL.n305 B 0.025505f
C641 VTAIL.n306 B 0.050662f
C642 VTAIL.n307 B 0.011108f
C643 VTAIL.n308 B 0.010791f
C644 VTAIL.n309 B 0.047788f
C645 VTAIL.n310 B 0.027921f
C646 VTAIL.n311 B 1.20982f
C647 VN.t1 B 2.79043f
C648 VN.t0 B 3.1796f
.ends

