* NGSPICE file created from diff_pair_sample_0806.ext - technology: sky130A

.subckt diff_pair_sample_0806 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=3.3696 ps=18.06 w=8.64 l=3.37
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.37
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=3.3696 ps=18.06 w=8.64 l=3.37
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.37
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=3.3696 ps=18.06 w=8.64 l=3.37
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.37
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.37
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=3.3696 ps=18.06 w=8.64 l=3.37
R0 VP.n0 VP.t1 144.672
R1 VP.n0 VP.t0 100.519
R2 VP VP.n0 0.526368
R3 VTAIL.n178 VTAIL.n138 289.615
R4 VTAIL.n40 VTAIL.n0 289.615
R5 VTAIL.n132 VTAIL.n92 289.615
R6 VTAIL.n86 VTAIL.n46 289.615
R7 VTAIL.n153 VTAIL.n152 185
R8 VTAIL.n150 VTAIL.n149 185
R9 VTAIL.n159 VTAIL.n158 185
R10 VTAIL.n161 VTAIL.n160 185
R11 VTAIL.n146 VTAIL.n145 185
R12 VTAIL.n167 VTAIL.n166 185
R13 VTAIL.n170 VTAIL.n169 185
R14 VTAIL.n168 VTAIL.n142 185
R15 VTAIL.n175 VTAIL.n141 185
R16 VTAIL.n177 VTAIL.n176 185
R17 VTAIL.n179 VTAIL.n178 185
R18 VTAIL.n15 VTAIL.n14 185
R19 VTAIL.n12 VTAIL.n11 185
R20 VTAIL.n21 VTAIL.n20 185
R21 VTAIL.n23 VTAIL.n22 185
R22 VTAIL.n8 VTAIL.n7 185
R23 VTAIL.n29 VTAIL.n28 185
R24 VTAIL.n32 VTAIL.n31 185
R25 VTAIL.n30 VTAIL.n4 185
R26 VTAIL.n37 VTAIL.n3 185
R27 VTAIL.n39 VTAIL.n38 185
R28 VTAIL.n41 VTAIL.n40 185
R29 VTAIL.n133 VTAIL.n132 185
R30 VTAIL.n131 VTAIL.n130 185
R31 VTAIL.n129 VTAIL.n95 185
R32 VTAIL.n99 VTAIL.n96 185
R33 VTAIL.n124 VTAIL.n123 185
R34 VTAIL.n122 VTAIL.n121 185
R35 VTAIL.n101 VTAIL.n100 185
R36 VTAIL.n116 VTAIL.n115 185
R37 VTAIL.n114 VTAIL.n113 185
R38 VTAIL.n105 VTAIL.n104 185
R39 VTAIL.n108 VTAIL.n107 185
R40 VTAIL.n87 VTAIL.n86 185
R41 VTAIL.n85 VTAIL.n84 185
R42 VTAIL.n83 VTAIL.n49 185
R43 VTAIL.n53 VTAIL.n50 185
R44 VTAIL.n78 VTAIL.n77 185
R45 VTAIL.n76 VTAIL.n75 185
R46 VTAIL.n55 VTAIL.n54 185
R47 VTAIL.n70 VTAIL.n69 185
R48 VTAIL.n68 VTAIL.n67 185
R49 VTAIL.n59 VTAIL.n58 185
R50 VTAIL.n62 VTAIL.n61 185
R51 VTAIL.t0 VTAIL.n151 149.524
R52 VTAIL.t2 VTAIL.n13 149.524
R53 VTAIL.t3 VTAIL.n106 149.524
R54 VTAIL.t1 VTAIL.n60 149.524
R55 VTAIL.n152 VTAIL.n149 104.615
R56 VTAIL.n159 VTAIL.n149 104.615
R57 VTAIL.n160 VTAIL.n159 104.615
R58 VTAIL.n160 VTAIL.n145 104.615
R59 VTAIL.n167 VTAIL.n145 104.615
R60 VTAIL.n169 VTAIL.n167 104.615
R61 VTAIL.n169 VTAIL.n168 104.615
R62 VTAIL.n168 VTAIL.n141 104.615
R63 VTAIL.n177 VTAIL.n141 104.615
R64 VTAIL.n178 VTAIL.n177 104.615
R65 VTAIL.n14 VTAIL.n11 104.615
R66 VTAIL.n21 VTAIL.n11 104.615
R67 VTAIL.n22 VTAIL.n21 104.615
R68 VTAIL.n22 VTAIL.n7 104.615
R69 VTAIL.n29 VTAIL.n7 104.615
R70 VTAIL.n31 VTAIL.n29 104.615
R71 VTAIL.n31 VTAIL.n30 104.615
R72 VTAIL.n30 VTAIL.n3 104.615
R73 VTAIL.n39 VTAIL.n3 104.615
R74 VTAIL.n40 VTAIL.n39 104.615
R75 VTAIL.n132 VTAIL.n131 104.615
R76 VTAIL.n131 VTAIL.n95 104.615
R77 VTAIL.n99 VTAIL.n95 104.615
R78 VTAIL.n123 VTAIL.n99 104.615
R79 VTAIL.n123 VTAIL.n122 104.615
R80 VTAIL.n122 VTAIL.n100 104.615
R81 VTAIL.n115 VTAIL.n100 104.615
R82 VTAIL.n115 VTAIL.n114 104.615
R83 VTAIL.n114 VTAIL.n104 104.615
R84 VTAIL.n107 VTAIL.n104 104.615
R85 VTAIL.n86 VTAIL.n85 104.615
R86 VTAIL.n85 VTAIL.n49 104.615
R87 VTAIL.n53 VTAIL.n49 104.615
R88 VTAIL.n77 VTAIL.n53 104.615
R89 VTAIL.n77 VTAIL.n76 104.615
R90 VTAIL.n76 VTAIL.n54 104.615
R91 VTAIL.n69 VTAIL.n54 104.615
R92 VTAIL.n69 VTAIL.n68 104.615
R93 VTAIL.n68 VTAIL.n58 104.615
R94 VTAIL.n61 VTAIL.n58 104.615
R95 VTAIL.n152 VTAIL.t0 52.3082
R96 VTAIL.n14 VTAIL.t2 52.3082
R97 VTAIL.n107 VTAIL.t3 52.3082
R98 VTAIL.n61 VTAIL.t1 52.3082
R99 VTAIL.n183 VTAIL.n182 34.5126
R100 VTAIL.n45 VTAIL.n44 34.5126
R101 VTAIL.n137 VTAIL.n136 34.5126
R102 VTAIL.n91 VTAIL.n90 34.5126
R103 VTAIL.n91 VTAIL.n45 26.1945
R104 VTAIL.n183 VTAIL.n137 23.0048
R105 VTAIL.n176 VTAIL.n175 13.1884
R106 VTAIL.n38 VTAIL.n37 13.1884
R107 VTAIL.n130 VTAIL.n129 13.1884
R108 VTAIL.n84 VTAIL.n83 13.1884
R109 VTAIL.n174 VTAIL.n142 12.8005
R110 VTAIL.n179 VTAIL.n140 12.8005
R111 VTAIL.n36 VTAIL.n4 12.8005
R112 VTAIL.n41 VTAIL.n2 12.8005
R113 VTAIL.n133 VTAIL.n94 12.8005
R114 VTAIL.n128 VTAIL.n96 12.8005
R115 VTAIL.n87 VTAIL.n48 12.8005
R116 VTAIL.n82 VTAIL.n50 12.8005
R117 VTAIL.n171 VTAIL.n170 12.0247
R118 VTAIL.n180 VTAIL.n138 12.0247
R119 VTAIL.n33 VTAIL.n32 12.0247
R120 VTAIL.n42 VTAIL.n0 12.0247
R121 VTAIL.n134 VTAIL.n92 12.0247
R122 VTAIL.n125 VTAIL.n124 12.0247
R123 VTAIL.n88 VTAIL.n46 12.0247
R124 VTAIL.n79 VTAIL.n78 12.0247
R125 VTAIL.n166 VTAIL.n144 11.249
R126 VTAIL.n28 VTAIL.n6 11.249
R127 VTAIL.n121 VTAIL.n98 11.249
R128 VTAIL.n75 VTAIL.n52 11.249
R129 VTAIL.n165 VTAIL.n146 10.4732
R130 VTAIL.n27 VTAIL.n8 10.4732
R131 VTAIL.n120 VTAIL.n101 10.4732
R132 VTAIL.n74 VTAIL.n55 10.4732
R133 VTAIL.n153 VTAIL.n151 10.2747
R134 VTAIL.n15 VTAIL.n13 10.2747
R135 VTAIL.n108 VTAIL.n106 10.2747
R136 VTAIL.n62 VTAIL.n60 10.2747
R137 VTAIL.n162 VTAIL.n161 9.69747
R138 VTAIL.n24 VTAIL.n23 9.69747
R139 VTAIL.n117 VTAIL.n116 9.69747
R140 VTAIL.n71 VTAIL.n70 9.69747
R141 VTAIL.n182 VTAIL.n181 9.45567
R142 VTAIL.n44 VTAIL.n43 9.45567
R143 VTAIL.n136 VTAIL.n135 9.45567
R144 VTAIL.n90 VTAIL.n89 9.45567
R145 VTAIL.n181 VTAIL.n180 9.3005
R146 VTAIL.n140 VTAIL.n139 9.3005
R147 VTAIL.n155 VTAIL.n154 9.3005
R148 VTAIL.n157 VTAIL.n156 9.3005
R149 VTAIL.n148 VTAIL.n147 9.3005
R150 VTAIL.n163 VTAIL.n162 9.3005
R151 VTAIL.n165 VTAIL.n164 9.3005
R152 VTAIL.n144 VTAIL.n143 9.3005
R153 VTAIL.n172 VTAIL.n171 9.3005
R154 VTAIL.n174 VTAIL.n173 9.3005
R155 VTAIL.n43 VTAIL.n42 9.3005
R156 VTAIL.n2 VTAIL.n1 9.3005
R157 VTAIL.n17 VTAIL.n16 9.3005
R158 VTAIL.n19 VTAIL.n18 9.3005
R159 VTAIL.n10 VTAIL.n9 9.3005
R160 VTAIL.n25 VTAIL.n24 9.3005
R161 VTAIL.n27 VTAIL.n26 9.3005
R162 VTAIL.n6 VTAIL.n5 9.3005
R163 VTAIL.n34 VTAIL.n33 9.3005
R164 VTAIL.n36 VTAIL.n35 9.3005
R165 VTAIL.n110 VTAIL.n109 9.3005
R166 VTAIL.n112 VTAIL.n111 9.3005
R167 VTAIL.n103 VTAIL.n102 9.3005
R168 VTAIL.n118 VTAIL.n117 9.3005
R169 VTAIL.n120 VTAIL.n119 9.3005
R170 VTAIL.n98 VTAIL.n97 9.3005
R171 VTAIL.n126 VTAIL.n125 9.3005
R172 VTAIL.n128 VTAIL.n127 9.3005
R173 VTAIL.n135 VTAIL.n134 9.3005
R174 VTAIL.n94 VTAIL.n93 9.3005
R175 VTAIL.n64 VTAIL.n63 9.3005
R176 VTAIL.n66 VTAIL.n65 9.3005
R177 VTAIL.n57 VTAIL.n56 9.3005
R178 VTAIL.n72 VTAIL.n71 9.3005
R179 VTAIL.n74 VTAIL.n73 9.3005
R180 VTAIL.n52 VTAIL.n51 9.3005
R181 VTAIL.n80 VTAIL.n79 9.3005
R182 VTAIL.n82 VTAIL.n81 9.3005
R183 VTAIL.n89 VTAIL.n88 9.3005
R184 VTAIL.n48 VTAIL.n47 9.3005
R185 VTAIL.n158 VTAIL.n148 8.92171
R186 VTAIL.n20 VTAIL.n10 8.92171
R187 VTAIL.n113 VTAIL.n103 8.92171
R188 VTAIL.n67 VTAIL.n57 8.92171
R189 VTAIL.n157 VTAIL.n150 8.14595
R190 VTAIL.n19 VTAIL.n12 8.14595
R191 VTAIL.n112 VTAIL.n105 8.14595
R192 VTAIL.n66 VTAIL.n59 8.14595
R193 VTAIL.n154 VTAIL.n153 7.3702
R194 VTAIL.n16 VTAIL.n15 7.3702
R195 VTAIL.n109 VTAIL.n108 7.3702
R196 VTAIL.n63 VTAIL.n62 7.3702
R197 VTAIL.n154 VTAIL.n150 5.81868
R198 VTAIL.n16 VTAIL.n12 5.81868
R199 VTAIL.n109 VTAIL.n105 5.81868
R200 VTAIL.n63 VTAIL.n59 5.81868
R201 VTAIL.n158 VTAIL.n157 5.04292
R202 VTAIL.n20 VTAIL.n19 5.04292
R203 VTAIL.n113 VTAIL.n112 5.04292
R204 VTAIL.n67 VTAIL.n66 5.04292
R205 VTAIL.n161 VTAIL.n148 4.26717
R206 VTAIL.n23 VTAIL.n10 4.26717
R207 VTAIL.n116 VTAIL.n103 4.26717
R208 VTAIL.n70 VTAIL.n57 4.26717
R209 VTAIL.n162 VTAIL.n146 3.49141
R210 VTAIL.n24 VTAIL.n8 3.49141
R211 VTAIL.n117 VTAIL.n101 3.49141
R212 VTAIL.n71 VTAIL.n55 3.49141
R213 VTAIL.n155 VTAIL.n151 2.84303
R214 VTAIL.n17 VTAIL.n13 2.84303
R215 VTAIL.n110 VTAIL.n106 2.84303
R216 VTAIL.n64 VTAIL.n60 2.84303
R217 VTAIL.n166 VTAIL.n165 2.71565
R218 VTAIL.n28 VTAIL.n27 2.71565
R219 VTAIL.n121 VTAIL.n120 2.71565
R220 VTAIL.n75 VTAIL.n74 2.71565
R221 VTAIL.n137 VTAIL.n91 2.06516
R222 VTAIL.n170 VTAIL.n144 1.93989
R223 VTAIL.n182 VTAIL.n138 1.93989
R224 VTAIL.n32 VTAIL.n6 1.93989
R225 VTAIL.n44 VTAIL.n0 1.93989
R226 VTAIL.n136 VTAIL.n92 1.93989
R227 VTAIL.n124 VTAIL.n98 1.93989
R228 VTAIL.n90 VTAIL.n46 1.93989
R229 VTAIL.n78 VTAIL.n52 1.93989
R230 VTAIL VTAIL.n45 1.32593
R231 VTAIL.n171 VTAIL.n142 1.16414
R232 VTAIL.n180 VTAIL.n179 1.16414
R233 VTAIL.n33 VTAIL.n4 1.16414
R234 VTAIL.n42 VTAIL.n41 1.16414
R235 VTAIL.n134 VTAIL.n133 1.16414
R236 VTAIL.n125 VTAIL.n96 1.16414
R237 VTAIL.n88 VTAIL.n87 1.16414
R238 VTAIL.n79 VTAIL.n50 1.16414
R239 VTAIL VTAIL.n183 0.739724
R240 VTAIL.n175 VTAIL.n174 0.388379
R241 VTAIL.n176 VTAIL.n140 0.388379
R242 VTAIL.n37 VTAIL.n36 0.388379
R243 VTAIL.n38 VTAIL.n2 0.388379
R244 VTAIL.n130 VTAIL.n94 0.388379
R245 VTAIL.n129 VTAIL.n128 0.388379
R246 VTAIL.n84 VTAIL.n48 0.388379
R247 VTAIL.n83 VTAIL.n82 0.388379
R248 VTAIL.n156 VTAIL.n155 0.155672
R249 VTAIL.n156 VTAIL.n147 0.155672
R250 VTAIL.n163 VTAIL.n147 0.155672
R251 VTAIL.n164 VTAIL.n163 0.155672
R252 VTAIL.n164 VTAIL.n143 0.155672
R253 VTAIL.n172 VTAIL.n143 0.155672
R254 VTAIL.n173 VTAIL.n172 0.155672
R255 VTAIL.n173 VTAIL.n139 0.155672
R256 VTAIL.n181 VTAIL.n139 0.155672
R257 VTAIL.n18 VTAIL.n17 0.155672
R258 VTAIL.n18 VTAIL.n9 0.155672
R259 VTAIL.n25 VTAIL.n9 0.155672
R260 VTAIL.n26 VTAIL.n25 0.155672
R261 VTAIL.n26 VTAIL.n5 0.155672
R262 VTAIL.n34 VTAIL.n5 0.155672
R263 VTAIL.n35 VTAIL.n34 0.155672
R264 VTAIL.n35 VTAIL.n1 0.155672
R265 VTAIL.n43 VTAIL.n1 0.155672
R266 VTAIL.n135 VTAIL.n93 0.155672
R267 VTAIL.n127 VTAIL.n93 0.155672
R268 VTAIL.n127 VTAIL.n126 0.155672
R269 VTAIL.n126 VTAIL.n97 0.155672
R270 VTAIL.n119 VTAIL.n97 0.155672
R271 VTAIL.n119 VTAIL.n118 0.155672
R272 VTAIL.n118 VTAIL.n102 0.155672
R273 VTAIL.n111 VTAIL.n102 0.155672
R274 VTAIL.n111 VTAIL.n110 0.155672
R275 VTAIL.n89 VTAIL.n47 0.155672
R276 VTAIL.n81 VTAIL.n47 0.155672
R277 VTAIL.n81 VTAIL.n80 0.155672
R278 VTAIL.n80 VTAIL.n51 0.155672
R279 VTAIL.n73 VTAIL.n51 0.155672
R280 VTAIL.n73 VTAIL.n72 0.155672
R281 VTAIL.n72 VTAIL.n56 0.155672
R282 VTAIL.n65 VTAIL.n56 0.155672
R283 VTAIL.n65 VTAIL.n64 0.155672
R284 VDD1.n40 VDD1.n0 289.615
R285 VDD1.n85 VDD1.n45 289.615
R286 VDD1.n41 VDD1.n40 185
R287 VDD1.n39 VDD1.n38 185
R288 VDD1.n37 VDD1.n3 185
R289 VDD1.n7 VDD1.n4 185
R290 VDD1.n32 VDD1.n31 185
R291 VDD1.n30 VDD1.n29 185
R292 VDD1.n9 VDD1.n8 185
R293 VDD1.n24 VDD1.n23 185
R294 VDD1.n22 VDD1.n21 185
R295 VDD1.n13 VDD1.n12 185
R296 VDD1.n16 VDD1.n15 185
R297 VDD1.n60 VDD1.n59 185
R298 VDD1.n57 VDD1.n56 185
R299 VDD1.n66 VDD1.n65 185
R300 VDD1.n68 VDD1.n67 185
R301 VDD1.n53 VDD1.n52 185
R302 VDD1.n74 VDD1.n73 185
R303 VDD1.n77 VDD1.n76 185
R304 VDD1.n75 VDD1.n49 185
R305 VDD1.n82 VDD1.n48 185
R306 VDD1.n84 VDD1.n83 185
R307 VDD1.n86 VDD1.n85 185
R308 VDD1.t0 VDD1.n14 149.524
R309 VDD1.t1 VDD1.n58 149.524
R310 VDD1.n40 VDD1.n39 104.615
R311 VDD1.n39 VDD1.n3 104.615
R312 VDD1.n7 VDD1.n3 104.615
R313 VDD1.n31 VDD1.n7 104.615
R314 VDD1.n31 VDD1.n30 104.615
R315 VDD1.n30 VDD1.n8 104.615
R316 VDD1.n23 VDD1.n8 104.615
R317 VDD1.n23 VDD1.n22 104.615
R318 VDD1.n22 VDD1.n12 104.615
R319 VDD1.n15 VDD1.n12 104.615
R320 VDD1.n59 VDD1.n56 104.615
R321 VDD1.n66 VDD1.n56 104.615
R322 VDD1.n67 VDD1.n66 104.615
R323 VDD1.n67 VDD1.n52 104.615
R324 VDD1.n74 VDD1.n52 104.615
R325 VDD1.n76 VDD1.n74 104.615
R326 VDD1.n76 VDD1.n75 104.615
R327 VDD1.n75 VDD1.n48 104.615
R328 VDD1.n84 VDD1.n48 104.615
R329 VDD1.n85 VDD1.n84 104.615
R330 VDD1 VDD1.n89 90.0007
R331 VDD1.n15 VDD1.t0 52.3082
R332 VDD1.n59 VDD1.t1 52.3082
R333 VDD1 VDD1.n44 52.047
R334 VDD1.n38 VDD1.n37 13.1884
R335 VDD1.n83 VDD1.n82 13.1884
R336 VDD1.n41 VDD1.n2 12.8005
R337 VDD1.n36 VDD1.n4 12.8005
R338 VDD1.n81 VDD1.n49 12.8005
R339 VDD1.n86 VDD1.n47 12.8005
R340 VDD1.n42 VDD1.n0 12.0247
R341 VDD1.n33 VDD1.n32 12.0247
R342 VDD1.n78 VDD1.n77 12.0247
R343 VDD1.n87 VDD1.n45 12.0247
R344 VDD1.n29 VDD1.n6 11.249
R345 VDD1.n73 VDD1.n51 11.249
R346 VDD1.n28 VDD1.n9 10.4732
R347 VDD1.n72 VDD1.n53 10.4732
R348 VDD1.n16 VDD1.n14 10.2747
R349 VDD1.n60 VDD1.n58 10.2747
R350 VDD1.n25 VDD1.n24 9.69747
R351 VDD1.n69 VDD1.n68 9.69747
R352 VDD1.n44 VDD1.n43 9.45567
R353 VDD1.n89 VDD1.n88 9.45567
R354 VDD1.n18 VDD1.n17 9.3005
R355 VDD1.n20 VDD1.n19 9.3005
R356 VDD1.n11 VDD1.n10 9.3005
R357 VDD1.n26 VDD1.n25 9.3005
R358 VDD1.n28 VDD1.n27 9.3005
R359 VDD1.n6 VDD1.n5 9.3005
R360 VDD1.n34 VDD1.n33 9.3005
R361 VDD1.n36 VDD1.n35 9.3005
R362 VDD1.n43 VDD1.n42 9.3005
R363 VDD1.n2 VDD1.n1 9.3005
R364 VDD1.n88 VDD1.n87 9.3005
R365 VDD1.n47 VDD1.n46 9.3005
R366 VDD1.n62 VDD1.n61 9.3005
R367 VDD1.n64 VDD1.n63 9.3005
R368 VDD1.n55 VDD1.n54 9.3005
R369 VDD1.n70 VDD1.n69 9.3005
R370 VDD1.n72 VDD1.n71 9.3005
R371 VDD1.n51 VDD1.n50 9.3005
R372 VDD1.n79 VDD1.n78 9.3005
R373 VDD1.n81 VDD1.n80 9.3005
R374 VDD1.n21 VDD1.n11 8.92171
R375 VDD1.n65 VDD1.n55 8.92171
R376 VDD1.n20 VDD1.n13 8.14595
R377 VDD1.n64 VDD1.n57 8.14595
R378 VDD1.n17 VDD1.n16 7.3702
R379 VDD1.n61 VDD1.n60 7.3702
R380 VDD1.n17 VDD1.n13 5.81868
R381 VDD1.n61 VDD1.n57 5.81868
R382 VDD1.n21 VDD1.n20 5.04292
R383 VDD1.n65 VDD1.n64 5.04292
R384 VDD1.n24 VDD1.n11 4.26717
R385 VDD1.n68 VDD1.n55 4.26717
R386 VDD1.n25 VDD1.n9 3.49141
R387 VDD1.n69 VDD1.n53 3.49141
R388 VDD1.n62 VDD1.n58 2.84303
R389 VDD1.n18 VDD1.n14 2.84303
R390 VDD1.n29 VDD1.n28 2.71565
R391 VDD1.n73 VDD1.n72 2.71565
R392 VDD1.n44 VDD1.n0 1.93989
R393 VDD1.n32 VDD1.n6 1.93989
R394 VDD1.n77 VDD1.n51 1.93989
R395 VDD1.n89 VDD1.n45 1.93989
R396 VDD1.n42 VDD1.n41 1.16414
R397 VDD1.n33 VDD1.n4 1.16414
R398 VDD1.n78 VDD1.n49 1.16414
R399 VDD1.n87 VDD1.n86 1.16414
R400 VDD1.n38 VDD1.n2 0.388379
R401 VDD1.n37 VDD1.n36 0.388379
R402 VDD1.n82 VDD1.n81 0.388379
R403 VDD1.n83 VDD1.n47 0.388379
R404 VDD1.n43 VDD1.n1 0.155672
R405 VDD1.n35 VDD1.n1 0.155672
R406 VDD1.n35 VDD1.n34 0.155672
R407 VDD1.n34 VDD1.n5 0.155672
R408 VDD1.n27 VDD1.n5 0.155672
R409 VDD1.n27 VDD1.n26 0.155672
R410 VDD1.n26 VDD1.n10 0.155672
R411 VDD1.n19 VDD1.n10 0.155672
R412 VDD1.n19 VDD1.n18 0.155672
R413 VDD1.n63 VDD1.n62 0.155672
R414 VDD1.n63 VDD1.n54 0.155672
R415 VDD1.n70 VDD1.n54 0.155672
R416 VDD1.n71 VDD1.n70 0.155672
R417 VDD1.n71 VDD1.n50 0.155672
R418 VDD1.n79 VDD1.n50 0.155672
R419 VDD1.n80 VDD1.n79 0.155672
R420 VDD1.n80 VDD1.n46 0.155672
R421 VDD1.n88 VDD1.n46 0.155672
R422 B.n473 B.n98 585
R423 B.n98 B.n57 585
R424 B.n475 B.n474 585
R425 B.n477 B.n97 585
R426 B.n480 B.n479 585
R427 B.n481 B.n96 585
R428 B.n483 B.n482 585
R429 B.n485 B.n95 585
R430 B.n488 B.n487 585
R431 B.n489 B.n94 585
R432 B.n491 B.n490 585
R433 B.n493 B.n93 585
R434 B.n496 B.n495 585
R435 B.n497 B.n92 585
R436 B.n499 B.n498 585
R437 B.n501 B.n91 585
R438 B.n504 B.n503 585
R439 B.n505 B.n90 585
R440 B.n507 B.n506 585
R441 B.n509 B.n89 585
R442 B.n512 B.n511 585
R443 B.n513 B.n88 585
R444 B.n515 B.n514 585
R445 B.n517 B.n87 585
R446 B.n520 B.n519 585
R447 B.n521 B.n86 585
R448 B.n523 B.n522 585
R449 B.n525 B.n85 585
R450 B.n528 B.n527 585
R451 B.n529 B.n84 585
R452 B.n531 B.n530 585
R453 B.n533 B.n83 585
R454 B.n536 B.n535 585
R455 B.n538 B.n80 585
R456 B.n540 B.n539 585
R457 B.n542 B.n79 585
R458 B.n545 B.n544 585
R459 B.n546 B.n78 585
R460 B.n548 B.n547 585
R461 B.n550 B.n77 585
R462 B.n553 B.n552 585
R463 B.n554 B.n74 585
R464 B.n557 B.n556 585
R465 B.n559 B.n73 585
R466 B.n562 B.n561 585
R467 B.n563 B.n72 585
R468 B.n565 B.n564 585
R469 B.n567 B.n71 585
R470 B.n570 B.n569 585
R471 B.n571 B.n70 585
R472 B.n573 B.n572 585
R473 B.n575 B.n69 585
R474 B.n578 B.n577 585
R475 B.n579 B.n68 585
R476 B.n581 B.n580 585
R477 B.n583 B.n67 585
R478 B.n586 B.n585 585
R479 B.n587 B.n66 585
R480 B.n589 B.n588 585
R481 B.n591 B.n65 585
R482 B.n594 B.n593 585
R483 B.n595 B.n64 585
R484 B.n597 B.n596 585
R485 B.n599 B.n63 585
R486 B.n602 B.n601 585
R487 B.n603 B.n62 585
R488 B.n605 B.n604 585
R489 B.n607 B.n61 585
R490 B.n610 B.n609 585
R491 B.n611 B.n60 585
R492 B.n613 B.n612 585
R493 B.n615 B.n59 585
R494 B.n618 B.n617 585
R495 B.n619 B.n58 585
R496 B.n472 B.n56 585
R497 B.n622 B.n56 585
R498 B.n471 B.n55 585
R499 B.n623 B.n55 585
R500 B.n470 B.n54 585
R501 B.n624 B.n54 585
R502 B.n469 B.n468 585
R503 B.n468 B.n50 585
R504 B.n467 B.n49 585
R505 B.n630 B.n49 585
R506 B.n466 B.n48 585
R507 B.n631 B.n48 585
R508 B.n465 B.n47 585
R509 B.n632 B.n47 585
R510 B.n464 B.n463 585
R511 B.n463 B.n43 585
R512 B.n462 B.n42 585
R513 B.n638 B.n42 585
R514 B.n461 B.n41 585
R515 B.n639 B.n41 585
R516 B.n460 B.n40 585
R517 B.n640 B.n40 585
R518 B.n459 B.n458 585
R519 B.n458 B.n36 585
R520 B.n457 B.n35 585
R521 B.n646 B.n35 585
R522 B.n456 B.n34 585
R523 B.n647 B.n34 585
R524 B.n455 B.n33 585
R525 B.n648 B.n33 585
R526 B.n454 B.n453 585
R527 B.n453 B.n29 585
R528 B.n452 B.n28 585
R529 B.n654 B.n28 585
R530 B.n451 B.n27 585
R531 B.n655 B.n27 585
R532 B.n450 B.n26 585
R533 B.n656 B.n26 585
R534 B.n449 B.n448 585
R535 B.n448 B.n22 585
R536 B.n447 B.n21 585
R537 B.n662 B.n21 585
R538 B.n446 B.n20 585
R539 B.n663 B.n20 585
R540 B.n445 B.n19 585
R541 B.n664 B.n19 585
R542 B.n444 B.n443 585
R543 B.n443 B.n15 585
R544 B.n442 B.n14 585
R545 B.n670 B.n14 585
R546 B.n441 B.n13 585
R547 B.n671 B.n13 585
R548 B.n440 B.n12 585
R549 B.n672 B.n12 585
R550 B.n439 B.n438 585
R551 B.n438 B.n8 585
R552 B.n437 B.n7 585
R553 B.n678 B.n7 585
R554 B.n436 B.n6 585
R555 B.n679 B.n6 585
R556 B.n435 B.n5 585
R557 B.n680 B.n5 585
R558 B.n434 B.n433 585
R559 B.n433 B.n4 585
R560 B.n432 B.n99 585
R561 B.n432 B.n431 585
R562 B.n422 B.n100 585
R563 B.n101 B.n100 585
R564 B.n424 B.n423 585
R565 B.n425 B.n424 585
R566 B.n421 B.n106 585
R567 B.n106 B.n105 585
R568 B.n420 B.n419 585
R569 B.n419 B.n418 585
R570 B.n108 B.n107 585
R571 B.n109 B.n108 585
R572 B.n411 B.n410 585
R573 B.n412 B.n411 585
R574 B.n409 B.n114 585
R575 B.n114 B.n113 585
R576 B.n408 B.n407 585
R577 B.n407 B.n406 585
R578 B.n116 B.n115 585
R579 B.n117 B.n116 585
R580 B.n399 B.n398 585
R581 B.n400 B.n399 585
R582 B.n397 B.n122 585
R583 B.n122 B.n121 585
R584 B.n396 B.n395 585
R585 B.n395 B.n394 585
R586 B.n124 B.n123 585
R587 B.n125 B.n124 585
R588 B.n387 B.n386 585
R589 B.n388 B.n387 585
R590 B.n385 B.n130 585
R591 B.n130 B.n129 585
R592 B.n384 B.n383 585
R593 B.n383 B.n382 585
R594 B.n132 B.n131 585
R595 B.n133 B.n132 585
R596 B.n375 B.n374 585
R597 B.n376 B.n375 585
R598 B.n373 B.n138 585
R599 B.n138 B.n137 585
R600 B.n372 B.n371 585
R601 B.n371 B.n370 585
R602 B.n140 B.n139 585
R603 B.n141 B.n140 585
R604 B.n363 B.n362 585
R605 B.n364 B.n363 585
R606 B.n361 B.n146 585
R607 B.n146 B.n145 585
R608 B.n360 B.n359 585
R609 B.n359 B.n358 585
R610 B.n148 B.n147 585
R611 B.n149 B.n148 585
R612 B.n351 B.n350 585
R613 B.n352 B.n351 585
R614 B.n349 B.n154 585
R615 B.n154 B.n153 585
R616 B.n348 B.n347 585
R617 B.n347 B.n346 585
R618 B.n343 B.n158 585
R619 B.n342 B.n341 585
R620 B.n339 B.n159 585
R621 B.n339 B.n157 585
R622 B.n338 B.n337 585
R623 B.n336 B.n335 585
R624 B.n334 B.n161 585
R625 B.n332 B.n331 585
R626 B.n330 B.n162 585
R627 B.n329 B.n328 585
R628 B.n326 B.n163 585
R629 B.n324 B.n323 585
R630 B.n322 B.n164 585
R631 B.n321 B.n320 585
R632 B.n318 B.n165 585
R633 B.n316 B.n315 585
R634 B.n314 B.n166 585
R635 B.n313 B.n312 585
R636 B.n310 B.n167 585
R637 B.n308 B.n307 585
R638 B.n306 B.n168 585
R639 B.n305 B.n304 585
R640 B.n302 B.n169 585
R641 B.n300 B.n299 585
R642 B.n298 B.n170 585
R643 B.n297 B.n296 585
R644 B.n294 B.n171 585
R645 B.n292 B.n291 585
R646 B.n290 B.n172 585
R647 B.n289 B.n288 585
R648 B.n286 B.n173 585
R649 B.n284 B.n283 585
R650 B.n282 B.n174 585
R651 B.n280 B.n279 585
R652 B.n277 B.n177 585
R653 B.n275 B.n274 585
R654 B.n273 B.n178 585
R655 B.n272 B.n271 585
R656 B.n269 B.n179 585
R657 B.n267 B.n266 585
R658 B.n265 B.n180 585
R659 B.n264 B.n263 585
R660 B.n261 B.n260 585
R661 B.n259 B.n258 585
R662 B.n257 B.n185 585
R663 B.n255 B.n254 585
R664 B.n253 B.n186 585
R665 B.n252 B.n251 585
R666 B.n249 B.n187 585
R667 B.n247 B.n246 585
R668 B.n245 B.n188 585
R669 B.n244 B.n243 585
R670 B.n241 B.n189 585
R671 B.n239 B.n238 585
R672 B.n237 B.n190 585
R673 B.n236 B.n235 585
R674 B.n233 B.n191 585
R675 B.n231 B.n230 585
R676 B.n229 B.n192 585
R677 B.n228 B.n227 585
R678 B.n225 B.n193 585
R679 B.n223 B.n222 585
R680 B.n221 B.n194 585
R681 B.n220 B.n219 585
R682 B.n217 B.n195 585
R683 B.n215 B.n214 585
R684 B.n213 B.n196 585
R685 B.n212 B.n211 585
R686 B.n209 B.n197 585
R687 B.n207 B.n206 585
R688 B.n205 B.n198 585
R689 B.n204 B.n203 585
R690 B.n201 B.n199 585
R691 B.n156 B.n155 585
R692 B.n345 B.n344 585
R693 B.n346 B.n345 585
R694 B.n152 B.n151 585
R695 B.n153 B.n152 585
R696 B.n354 B.n353 585
R697 B.n353 B.n352 585
R698 B.n355 B.n150 585
R699 B.n150 B.n149 585
R700 B.n357 B.n356 585
R701 B.n358 B.n357 585
R702 B.n144 B.n143 585
R703 B.n145 B.n144 585
R704 B.n366 B.n365 585
R705 B.n365 B.n364 585
R706 B.n367 B.n142 585
R707 B.n142 B.n141 585
R708 B.n369 B.n368 585
R709 B.n370 B.n369 585
R710 B.n136 B.n135 585
R711 B.n137 B.n136 585
R712 B.n378 B.n377 585
R713 B.n377 B.n376 585
R714 B.n379 B.n134 585
R715 B.n134 B.n133 585
R716 B.n381 B.n380 585
R717 B.n382 B.n381 585
R718 B.n128 B.n127 585
R719 B.n129 B.n128 585
R720 B.n390 B.n389 585
R721 B.n389 B.n388 585
R722 B.n391 B.n126 585
R723 B.n126 B.n125 585
R724 B.n393 B.n392 585
R725 B.n394 B.n393 585
R726 B.n120 B.n119 585
R727 B.n121 B.n120 585
R728 B.n402 B.n401 585
R729 B.n401 B.n400 585
R730 B.n403 B.n118 585
R731 B.n118 B.n117 585
R732 B.n405 B.n404 585
R733 B.n406 B.n405 585
R734 B.n112 B.n111 585
R735 B.n113 B.n112 585
R736 B.n414 B.n413 585
R737 B.n413 B.n412 585
R738 B.n415 B.n110 585
R739 B.n110 B.n109 585
R740 B.n417 B.n416 585
R741 B.n418 B.n417 585
R742 B.n104 B.n103 585
R743 B.n105 B.n104 585
R744 B.n427 B.n426 585
R745 B.n426 B.n425 585
R746 B.n428 B.n102 585
R747 B.n102 B.n101 585
R748 B.n430 B.n429 585
R749 B.n431 B.n430 585
R750 B.n2 B.n0 585
R751 B.n4 B.n2 585
R752 B.n3 B.n1 585
R753 B.n679 B.n3 585
R754 B.n677 B.n676 585
R755 B.n678 B.n677 585
R756 B.n675 B.n9 585
R757 B.n9 B.n8 585
R758 B.n674 B.n673 585
R759 B.n673 B.n672 585
R760 B.n11 B.n10 585
R761 B.n671 B.n11 585
R762 B.n669 B.n668 585
R763 B.n670 B.n669 585
R764 B.n667 B.n16 585
R765 B.n16 B.n15 585
R766 B.n666 B.n665 585
R767 B.n665 B.n664 585
R768 B.n18 B.n17 585
R769 B.n663 B.n18 585
R770 B.n661 B.n660 585
R771 B.n662 B.n661 585
R772 B.n659 B.n23 585
R773 B.n23 B.n22 585
R774 B.n658 B.n657 585
R775 B.n657 B.n656 585
R776 B.n25 B.n24 585
R777 B.n655 B.n25 585
R778 B.n653 B.n652 585
R779 B.n654 B.n653 585
R780 B.n651 B.n30 585
R781 B.n30 B.n29 585
R782 B.n650 B.n649 585
R783 B.n649 B.n648 585
R784 B.n32 B.n31 585
R785 B.n647 B.n32 585
R786 B.n645 B.n644 585
R787 B.n646 B.n645 585
R788 B.n643 B.n37 585
R789 B.n37 B.n36 585
R790 B.n642 B.n641 585
R791 B.n641 B.n640 585
R792 B.n39 B.n38 585
R793 B.n639 B.n39 585
R794 B.n637 B.n636 585
R795 B.n638 B.n637 585
R796 B.n635 B.n44 585
R797 B.n44 B.n43 585
R798 B.n634 B.n633 585
R799 B.n633 B.n632 585
R800 B.n46 B.n45 585
R801 B.n631 B.n46 585
R802 B.n629 B.n628 585
R803 B.n630 B.n629 585
R804 B.n627 B.n51 585
R805 B.n51 B.n50 585
R806 B.n626 B.n625 585
R807 B.n625 B.n624 585
R808 B.n53 B.n52 585
R809 B.n623 B.n53 585
R810 B.n621 B.n620 585
R811 B.n622 B.n621 585
R812 B.n682 B.n681 585
R813 B.n681 B.n680 585
R814 B.n345 B.n158 482.89
R815 B.n621 B.n58 482.89
R816 B.n347 B.n156 482.89
R817 B.n98 B.n56 482.89
R818 B.n181 B.t5 295.983
R819 B.n81 B.t8 295.983
R820 B.n175 B.t12 295.983
R821 B.n75 B.t14 295.983
R822 B.n181 B.t2 270.76
R823 B.n175 B.t10 270.76
R824 B.n75 B.t13 270.76
R825 B.n81 B.t6 270.76
R826 B.n476 B.n57 256.663
R827 B.n478 B.n57 256.663
R828 B.n484 B.n57 256.663
R829 B.n486 B.n57 256.663
R830 B.n492 B.n57 256.663
R831 B.n494 B.n57 256.663
R832 B.n500 B.n57 256.663
R833 B.n502 B.n57 256.663
R834 B.n508 B.n57 256.663
R835 B.n510 B.n57 256.663
R836 B.n516 B.n57 256.663
R837 B.n518 B.n57 256.663
R838 B.n524 B.n57 256.663
R839 B.n526 B.n57 256.663
R840 B.n532 B.n57 256.663
R841 B.n534 B.n57 256.663
R842 B.n541 B.n57 256.663
R843 B.n543 B.n57 256.663
R844 B.n549 B.n57 256.663
R845 B.n551 B.n57 256.663
R846 B.n558 B.n57 256.663
R847 B.n560 B.n57 256.663
R848 B.n566 B.n57 256.663
R849 B.n568 B.n57 256.663
R850 B.n574 B.n57 256.663
R851 B.n576 B.n57 256.663
R852 B.n582 B.n57 256.663
R853 B.n584 B.n57 256.663
R854 B.n590 B.n57 256.663
R855 B.n592 B.n57 256.663
R856 B.n598 B.n57 256.663
R857 B.n600 B.n57 256.663
R858 B.n606 B.n57 256.663
R859 B.n608 B.n57 256.663
R860 B.n614 B.n57 256.663
R861 B.n616 B.n57 256.663
R862 B.n340 B.n157 256.663
R863 B.n160 B.n157 256.663
R864 B.n333 B.n157 256.663
R865 B.n327 B.n157 256.663
R866 B.n325 B.n157 256.663
R867 B.n319 B.n157 256.663
R868 B.n317 B.n157 256.663
R869 B.n311 B.n157 256.663
R870 B.n309 B.n157 256.663
R871 B.n303 B.n157 256.663
R872 B.n301 B.n157 256.663
R873 B.n295 B.n157 256.663
R874 B.n293 B.n157 256.663
R875 B.n287 B.n157 256.663
R876 B.n285 B.n157 256.663
R877 B.n278 B.n157 256.663
R878 B.n276 B.n157 256.663
R879 B.n270 B.n157 256.663
R880 B.n268 B.n157 256.663
R881 B.n262 B.n157 256.663
R882 B.n184 B.n157 256.663
R883 B.n256 B.n157 256.663
R884 B.n250 B.n157 256.663
R885 B.n248 B.n157 256.663
R886 B.n242 B.n157 256.663
R887 B.n240 B.n157 256.663
R888 B.n234 B.n157 256.663
R889 B.n232 B.n157 256.663
R890 B.n226 B.n157 256.663
R891 B.n224 B.n157 256.663
R892 B.n218 B.n157 256.663
R893 B.n216 B.n157 256.663
R894 B.n210 B.n157 256.663
R895 B.n208 B.n157 256.663
R896 B.n202 B.n157 256.663
R897 B.n200 B.n157 256.663
R898 B.n182 B.t4 224.225
R899 B.n82 B.t9 224.225
R900 B.n176 B.t11 224.225
R901 B.n76 B.t15 224.225
R902 B.n345 B.n152 163.367
R903 B.n353 B.n152 163.367
R904 B.n353 B.n150 163.367
R905 B.n357 B.n150 163.367
R906 B.n357 B.n144 163.367
R907 B.n365 B.n144 163.367
R908 B.n365 B.n142 163.367
R909 B.n369 B.n142 163.367
R910 B.n369 B.n136 163.367
R911 B.n377 B.n136 163.367
R912 B.n377 B.n134 163.367
R913 B.n381 B.n134 163.367
R914 B.n381 B.n128 163.367
R915 B.n389 B.n128 163.367
R916 B.n389 B.n126 163.367
R917 B.n393 B.n126 163.367
R918 B.n393 B.n120 163.367
R919 B.n401 B.n120 163.367
R920 B.n401 B.n118 163.367
R921 B.n405 B.n118 163.367
R922 B.n405 B.n112 163.367
R923 B.n413 B.n112 163.367
R924 B.n413 B.n110 163.367
R925 B.n417 B.n110 163.367
R926 B.n417 B.n104 163.367
R927 B.n426 B.n104 163.367
R928 B.n426 B.n102 163.367
R929 B.n430 B.n102 163.367
R930 B.n430 B.n2 163.367
R931 B.n681 B.n2 163.367
R932 B.n681 B.n3 163.367
R933 B.n677 B.n3 163.367
R934 B.n677 B.n9 163.367
R935 B.n673 B.n9 163.367
R936 B.n673 B.n11 163.367
R937 B.n669 B.n11 163.367
R938 B.n669 B.n16 163.367
R939 B.n665 B.n16 163.367
R940 B.n665 B.n18 163.367
R941 B.n661 B.n18 163.367
R942 B.n661 B.n23 163.367
R943 B.n657 B.n23 163.367
R944 B.n657 B.n25 163.367
R945 B.n653 B.n25 163.367
R946 B.n653 B.n30 163.367
R947 B.n649 B.n30 163.367
R948 B.n649 B.n32 163.367
R949 B.n645 B.n32 163.367
R950 B.n645 B.n37 163.367
R951 B.n641 B.n37 163.367
R952 B.n641 B.n39 163.367
R953 B.n637 B.n39 163.367
R954 B.n637 B.n44 163.367
R955 B.n633 B.n44 163.367
R956 B.n633 B.n46 163.367
R957 B.n629 B.n46 163.367
R958 B.n629 B.n51 163.367
R959 B.n625 B.n51 163.367
R960 B.n625 B.n53 163.367
R961 B.n621 B.n53 163.367
R962 B.n341 B.n339 163.367
R963 B.n339 B.n338 163.367
R964 B.n335 B.n334 163.367
R965 B.n332 B.n162 163.367
R966 B.n328 B.n326 163.367
R967 B.n324 B.n164 163.367
R968 B.n320 B.n318 163.367
R969 B.n316 B.n166 163.367
R970 B.n312 B.n310 163.367
R971 B.n308 B.n168 163.367
R972 B.n304 B.n302 163.367
R973 B.n300 B.n170 163.367
R974 B.n296 B.n294 163.367
R975 B.n292 B.n172 163.367
R976 B.n288 B.n286 163.367
R977 B.n284 B.n174 163.367
R978 B.n279 B.n277 163.367
R979 B.n275 B.n178 163.367
R980 B.n271 B.n269 163.367
R981 B.n267 B.n180 163.367
R982 B.n263 B.n261 163.367
R983 B.n258 B.n257 163.367
R984 B.n255 B.n186 163.367
R985 B.n251 B.n249 163.367
R986 B.n247 B.n188 163.367
R987 B.n243 B.n241 163.367
R988 B.n239 B.n190 163.367
R989 B.n235 B.n233 163.367
R990 B.n231 B.n192 163.367
R991 B.n227 B.n225 163.367
R992 B.n223 B.n194 163.367
R993 B.n219 B.n217 163.367
R994 B.n215 B.n196 163.367
R995 B.n211 B.n209 163.367
R996 B.n207 B.n198 163.367
R997 B.n203 B.n201 163.367
R998 B.n347 B.n154 163.367
R999 B.n351 B.n154 163.367
R1000 B.n351 B.n148 163.367
R1001 B.n359 B.n148 163.367
R1002 B.n359 B.n146 163.367
R1003 B.n363 B.n146 163.367
R1004 B.n363 B.n140 163.367
R1005 B.n371 B.n140 163.367
R1006 B.n371 B.n138 163.367
R1007 B.n375 B.n138 163.367
R1008 B.n375 B.n132 163.367
R1009 B.n383 B.n132 163.367
R1010 B.n383 B.n130 163.367
R1011 B.n387 B.n130 163.367
R1012 B.n387 B.n124 163.367
R1013 B.n395 B.n124 163.367
R1014 B.n395 B.n122 163.367
R1015 B.n399 B.n122 163.367
R1016 B.n399 B.n116 163.367
R1017 B.n407 B.n116 163.367
R1018 B.n407 B.n114 163.367
R1019 B.n411 B.n114 163.367
R1020 B.n411 B.n108 163.367
R1021 B.n419 B.n108 163.367
R1022 B.n419 B.n106 163.367
R1023 B.n424 B.n106 163.367
R1024 B.n424 B.n100 163.367
R1025 B.n432 B.n100 163.367
R1026 B.n433 B.n432 163.367
R1027 B.n433 B.n5 163.367
R1028 B.n6 B.n5 163.367
R1029 B.n7 B.n6 163.367
R1030 B.n438 B.n7 163.367
R1031 B.n438 B.n12 163.367
R1032 B.n13 B.n12 163.367
R1033 B.n14 B.n13 163.367
R1034 B.n443 B.n14 163.367
R1035 B.n443 B.n19 163.367
R1036 B.n20 B.n19 163.367
R1037 B.n21 B.n20 163.367
R1038 B.n448 B.n21 163.367
R1039 B.n448 B.n26 163.367
R1040 B.n27 B.n26 163.367
R1041 B.n28 B.n27 163.367
R1042 B.n453 B.n28 163.367
R1043 B.n453 B.n33 163.367
R1044 B.n34 B.n33 163.367
R1045 B.n35 B.n34 163.367
R1046 B.n458 B.n35 163.367
R1047 B.n458 B.n40 163.367
R1048 B.n41 B.n40 163.367
R1049 B.n42 B.n41 163.367
R1050 B.n463 B.n42 163.367
R1051 B.n463 B.n47 163.367
R1052 B.n48 B.n47 163.367
R1053 B.n49 B.n48 163.367
R1054 B.n468 B.n49 163.367
R1055 B.n468 B.n54 163.367
R1056 B.n55 B.n54 163.367
R1057 B.n56 B.n55 163.367
R1058 B.n617 B.n615 163.367
R1059 B.n613 B.n60 163.367
R1060 B.n609 B.n607 163.367
R1061 B.n605 B.n62 163.367
R1062 B.n601 B.n599 163.367
R1063 B.n597 B.n64 163.367
R1064 B.n593 B.n591 163.367
R1065 B.n589 B.n66 163.367
R1066 B.n585 B.n583 163.367
R1067 B.n581 B.n68 163.367
R1068 B.n577 B.n575 163.367
R1069 B.n573 B.n70 163.367
R1070 B.n569 B.n567 163.367
R1071 B.n565 B.n72 163.367
R1072 B.n561 B.n559 163.367
R1073 B.n557 B.n74 163.367
R1074 B.n552 B.n550 163.367
R1075 B.n548 B.n78 163.367
R1076 B.n544 B.n542 163.367
R1077 B.n540 B.n80 163.367
R1078 B.n535 B.n533 163.367
R1079 B.n531 B.n84 163.367
R1080 B.n527 B.n525 163.367
R1081 B.n523 B.n86 163.367
R1082 B.n519 B.n517 163.367
R1083 B.n515 B.n88 163.367
R1084 B.n511 B.n509 163.367
R1085 B.n507 B.n90 163.367
R1086 B.n503 B.n501 163.367
R1087 B.n499 B.n92 163.367
R1088 B.n495 B.n493 163.367
R1089 B.n491 B.n94 163.367
R1090 B.n487 B.n485 163.367
R1091 B.n483 B.n96 163.367
R1092 B.n479 B.n477 163.367
R1093 B.n475 B.n98 163.367
R1094 B.n346 B.n157 90.9096
R1095 B.n622 B.n57 90.9096
R1096 B.n182 B.n181 71.7581
R1097 B.n176 B.n175 71.7581
R1098 B.n76 B.n75 71.7581
R1099 B.n82 B.n81 71.7581
R1100 B.n340 B.n158 71.676
R1101 B.n338 B.n160 71.676
R1102 B.n334 B.n333 71.676
R1103 B.n327 B.n162 71.676
R1104 B.n326 B.n325 71.676
R1105 B.n319 B.n164 71.676
R1106 B.n318 B.n317 71.676
R1107 B.n311 B.n166 71.676
R1108 B.n310 B.n309 71.676
R1109 B.n303 B.n168 71.676
R1110 B.n302 B.n301 71.676
R1111 B.n295 B.n170 71.676
R1112 B.n294 B.n293 71.676
R1113 B.n287 B.n172 71.676
R1114 B.n286 B.n285 71.676
R1115 B.n278 B.n174 71.676
R1116 B.n277 B.n276 71.676
R1117 B.n270 B.n178 71.676
R1118 B.n269 B.n268 71.676
R1119 B.n262 B.n180 71.676
R1120 B.n261 B.n184 71.676
R1121 B.n257 B.n256 71.676
R1122 B.n250 B.n186 71.676
R1123 B.n249 B.n248 71.676
R1124 B.n242 B.n188 71.676
R1125 B.n241 B.n240 71.676
R1126 B.n234 B.n190 71.676
R1127 B.n233 B.n232 71.676
R1128 B.n226 B.n192 71.676
R1129 B.n225 B.n224 71.676
R1130 B.n218 B.n194 71.676
R1131 B.n217 B.n216 71.676
R1132 B.n210 B.n196 71.676
R1133 B.n209 B.n208 71.676
R1134 B.n202 B.n198 71.676
R1135 B.n201 B.n200 71.676
R1136 B.n616 B.n58 71.676
R1137 B.n615 B.n614 71.676
R1138 B.n608 B.n60 71.676
R1139 B.n607 B.n606 71.676
R1140 B.n600 B.n62 71.676
R1141 B.n599 B.n598 71.676
R1142 B.n592 B.n64 71.676
R1143 B.n591 B.n590 71.676
R1144 B.n584 B.n66 71.676
R1145 B.n583 B.n582 71.676
R1146 B.n576 B.n68 71.676
R1147 B.n575 B.n574 71.676
R1148 B.n568 B.n70 71.676
R1149 B.n567 B.n566 71.676
R1150 B.n560 B.n72 71.676
R1151 B.n559 B.n558 71.676
R1152 B.n551 B.n74 71.676
R1153 B.n550 B.n549 71.676
R1154 B.n543 B.n78 71.676
R1155 B.n542 B.n541 71.676
R1156 B.n534 B.n80 71.676
R1157 B.n533 B.n532 71.676
R1158 B.n526 B.n84 71.676
R1159 B.n525 B.n524 71.676
R1160 B.n518 B.n86 71.676
R1161 B.n517 B.n516 71.676
R1162 B.n510 B.n88 71.676
R1163 B.n509 B.n508 71.676
R1164 B.n502 B.n90 71.676
R1165 B.n501 B.n500 71.676
R1166 B.n494 B.n92 71.676
R1167 B.n493 B.n492 71.676
R1168 B.n486 B.n94 71.676
R1169 B.n485 B.n484 71.676
R1170 B.n478 B.n96 71.676
R1171 B.n477 B.n476 71.676
R1172 B.n476 B.n475 71.676
R1173 B.n479 B.n478 71.676
R1174 B.n484 B.n483 71.676
R1175 B.n487 B.n486 71.676
R1176 B.n492 B.n491 71.676
R1177 B.n495 B.n494 71.676
R1178 B.n500 B.n499 71.676
R1179 B.n503 B.n502 71.676
R1180 B.n508 B.n507 71.676
R1181 B.n511 B.n510 71.676
R1182 B.n516 B.n515 71.676
R1183 B.n519 B.n518 71.676
R1184 B.n524 B.n523 71.676
R1185 B.n527 B.n526 71.676
R1186 B.n532 B.n531 71.676
R1187 B.n535 B.n534 71.676
R1188 B.n541 B.n540 71.676
R1189 B.n544 B.n543 71.676
R1190 B.n549 B.n548 71.676
R1191 B.n552 B.n551 71.676
R1192 B.n558 B.n557 71.676
R1193 B.n561 B.n560 71.676
R1194 B.n566 B.n565 71.676
R1195 B.n569 B.n568 71.676
R1196 B.n574 B.n573 71.676
R1197 B.n577 B.n576 71.676
R1198 B.n582 B.n581 71.676
R1199 B.n585 B.n584 71.676
R1200 B.n590 B.n589 71.676
R1201 B.n593 B.n592 71.676
R1202 B.n598 B.n597 71.676
R1203 B.n601 B.n600 71.676
R1204 B.n606 B.n605 71.676
R1205 B.n609 B.n608 71.676
R1206 B.n614 B.n613 71.676
R1207 B.n617 B.n616 71.676
R1208 B.n341 B.n340 71.676
R1209 B.n335 B.n160 71.676
R1210 B.n333 B.n332 71.676
R1211 B.n328 B.n327 71.676
R1212 B.n325 B.n324 71.676
R1213 B.n320 B.n319 71.676
R1214 B.n317 B.n316 71.676
R1215 B.n312 B.n311 71.676
R1216 B.n309 B.n308 71.676
R1217 B.n304 B.n303 71.676
R1218 B.n301 B.n300 71.676
R1219 B.n296 B.n295 71.676
R1220 B.n293 B.n292 71.676
R1221 B.n288 B.n287 71.676
R1222 B.n285 B.n284 71.676
R1223 B.n279 B.n278 71.676
R1224 B.n276 B.n275 71.676
R1225 B.n271 B.n270 71.676
R1226 B.n268 B.n267 71.676
R1227 B.n263 B.n262 71.676
R1228 B.n258 B.n184 71.676
R1229 B.n256 B.n255 71.676
R1230 B.n251 B.n250 71.676
R1231 B.n248 B.n247 71.676
R1232 B.n243 B.n242 71.676
R1233 B.n240 B.n239 71.676
R1234 B.n235 B.n234 71.676
R1235 B.n232 B.n231 71.676
R1236 B.n227 B.n226 71.676
R1237 B.n224 B.n223 71.676
R1238 B.n219 B.n218 71.676
R1239 B.n216 B.n215 71.676
R1240 B.n211 B.n210 71.676
R1241 B.n208 B.n207 71.676
R1242 B.n203 B.n202 71.676
R1243 B.n200 B.n156 71.676
R1244 B.n183 B.n182 59.5399
R1245 B.n281 B.n176 59.5399
R1246 B.n555 B.n76 59.5399
R1247 B.n537 B.n82 59.5399
R1248 B.n346 B.n153 53.7554
R1249 B.n352 B.n153 53.7554
R1250 B.n352 B.n149 53.7554
R1251 B.n358 B.n149 53.7554
R1252 B.n358 B.n145 53.7554
R1253 B.n364 B.n145 53.7554
R1254 B.n364 B.n141 53.7554
R1255 B.n370 B.n141 53.7554
R1256 B.n376 B.n137 53.7554
R1257 B.n376 B.n133 53.7554
R1258 B.n382 B.n133 53.7554
R1259 B.n382 B.n129 53.7554
R1260 B.n388 B.n129 53.7554
R1261 B.n388 B.n125 53.7554
R1262 B.n394 B.n125 53.7554
R1263 B.n394 B.n121 53.7554
R1264 B.n400 B.n121 53.7554
R1265 B.n400 B.n117 53.7554
R1266 B.n406 B.n117 53.7554
R1267 B.n406 B.n113 53.7554
R1268 B.n412 B.n113 53.7554
R1269 B.n418 B.n109 53.7554
R1270 B.n418 B.n105 53.7554
R1271 B.n425 B.n105 53.7554
R1272 B.n425 B.n101 53.7554
R1273 B.n431 B.n101 53.7554
R1274 B.n431 B.n4 53.7554
R1275 B.n680 B.n4 53.7554
R1276 B.n680 B.n679 53.7554
R1277 B.n679 B.n678 53.7554
R1278 B.n678 B.n8 53.7554
R1279 B.n672 B.n8 53.7554
R1280 B.n672 B.n671 53.7554
R1281 B.n671 B.n670 53.7554
R1282 B.n670 B.n15 53.7554
R1283 B.n664 B.n663 53.7554
R1284 B.n663 B.n662 53.7554
R1285 B.n662 B.n22 53.7554
R1286 B.n656 B.n22 53.7554
R1287 B.n656 B.n655 53.7554
R1288 B.n655 B.n654 53.7554
R1289 B.n654 B.n29 53.7554
R1290 B.n648 B.n29 53.7554
R1291 B.n648 B.n647 53.7554
R1292 B.n647 B.n646 53.7554
R1293 B.n646 B.n36 53.7554
R1294 B.n640 B.n36 53.7554
R1295 B.n640 B.n639 53.7554
R1296 B.n638 B.n43 53.7554
R1297 B.n632 B.n43 53.7554
R1298 B.n632 B.n631 53.7554
R1299 B.n631 B.n630 53.7554
R1300 B.n630 B.n50 53.7554
R1301 B.n624 B.n50 53.7554
R1302 B.n624 B.n623 53.7554
R1303 B.n623 B.n622 53.7554
R1304 B.n412 B.t1 51.3839
R1305 B.n664 B.t0 51.3839
R1306 B.n370 B.t3 46.6408
R1307 B.t7 B.n638 46.6408
R1308 B.n620 B.n619 31.3761
R1309 B.n473 B.n472 31.3761
R1310 B.n348 B.n155 31.3761
R1311 B.n344 B.n343 31.3761
R1312 B B.n682 18.0485
R1313 B.n619 B.n618 10.6151
R1314 B.n618 B.n59 10.6151
R1315 B.n612 B.n59 10.6151
R1316 B.n612 B.n611 10.6151
R1317 B.n611 B.n610 10.6151
R1318 B.n610 B.n61 10.6151
R1319 B.n604 B.n61 10.6151
R1320 B.n604 B.n603 10.6151
R1321 B.n603 B.n602 10.6151
R1322 B.n602 B.n63 10.6151
R1323 B.n596 B.n63 10.6151
R1324 B.n596 B.n595 10.6151
R1325 B.n595 B.n594 10.6151
R1326 B.n594 B.n65 10.6151
R1327 B.n588 B.n65 10.6151
R1328 B.n588 B.n587 10.6151
R1329 B.n587 B.n586 10.6151
R1330 B.n586 B.n67 10.6151
R1331 B.n580 B.n67 10.6151
R1332 B.n580 B.n579 10.6151
R1333 B.n579 B.n578 10.6151
R1334 B.n578 B.n69 10.6151
R1335 B.n572 B.n69 10.6151
R1336 B.n572 B.n571 10.6151
R1337 B.n571 B.n570 10.6151
R1338 B.n570 B.n71 10.6151
R1339 B.n564 B.n71 10.6151
R1340 B.n564 B.n563 10.6151
R1341 B.n563 B.n562 10.6151
R1342 B.n562 B.n73 10.6151
R1343 B.n556 B.n73 10.6151
R1344 B.n554 B.n553 10.6151
R1345 B.n553 B.n77 10.6151
R1346 B.n547 B.n77 10.6151
R1347 B.n547 B.n546 10.6151
R1348 B.n546 B.n545 10.6151
R1349 B.n545 B.n79 10.6151
R1350 B.n539 B.n79 10.6151
R1351 B.n539 B.n538 10.6151
R1352 B.n536 B.n83 10.6151
R1353 B.n530 B.n83 10.6151
R1354 B.n530 B.n529 10.6151
R1355 B.n529 B.n528 10.6151
R1356 B.n528 B.n85 10.6151
R1357 B.n522 B.n85 10.6151
R1358 B.n522 B.n521 10.6151
R1359 B.n521 B.n520 10.6151
R1360 B.n520 B.n87 10.6151
R1361 B.n514 B.n87 10.6151
R1362 B.n514 B.n513 10.6151
R1363 B.n513 B.n512 10.6151
R1364 B.n512 B.n89 10.6151
R1365 B.n506 B.n89 10.6151
R1366 B.n506 B.n505 10.6151
R1367 B.n505 B.n504 10.6151
R1368 B.n504 B.n91 10.6151
R1369 B.n498 B.n91 10.6151
R1370 B.n498 B.n497 10.6151
R1371 B.n497 B.n496 10.6151
R1372 B.n496 B.n93 10.6151
R1373 B.n490 B.n93 10.6151
R1374 B.n490 B.n489 10.6151
R1375 B.n489 B.n488 10.6151
R1376 B.n488 B.n95 10.6151
R1377 B.n482 B.n95 10.6151
R1378 B.n482 B.n481 10.6151
R1379 B.n481 B.n480 10.6151
R1380 B.n480 B.n97 10.6151
R1381 B.n474 B.n97 10.6151
R1382 B.n474 B.n473 10.6151
R1383 B.n349 B.n348 10.6151
R1384 B.n350 B.n349 10.6151
R1385 B.n350 B.n147 10.6151
R1386 B.n360 B.n147 10.6151
R1387 B.n361 B.n360 10.6151
R1388 B.n362 B.n361 10.6151
R1389 B.n362 B.n139 10.6151
R1390 B.n372 B.n139 10.6151
R1391 B.n373 B.n372 10.6151
R1392 B.n374 B.n373 10.6151
R1393 B.n374 B.n131 10.6151
R1394 B.n384 B.n131 10.6151
R1395 B.n385 B.n384 10.6151
R1396 B.n386 B.n385 10.6151
R1397 B.n386 B.n123 10.6151
R1398 B.n396 B.n123 10.6151
R1399 B.n397 B.n396 10.6151
R1400 B.n398 B.n397 10.6151
R1401 B.n398 B.n115 10.6151
R1402 B.n408 B.n115 10.6151
R1403 B.n409 B.n408 10.6151
R1404 B.n410 B.n409 10.6151
R1405 B.n410 B.n107 10.6151
R1406 B.n420 B.n107 10.6151
R1407 B.n421 B.n420 10.6151
R1408 B.n423 B.n421 10.6151
R1409 B.n423 B.n422 10.6151
R1410 B.n422 B.n99 10.6151
R1411 B.n434 B.n99 10.6151
R1412 B.n435 B.n434 10.6151
R1413 B.n436 B.n435 10.6151
R1414 B.n437 B.n436 10.6151
R1415 B.n439 B.n437 10.6151
R1416 B.n440 B.n439 10.6151
R1417 B.n441 B.n440 10.6151
R1418 B.n442 B.n441 10.6151
R1419 B.n444 B.n442 10.6151
R1420 B.n445 B.n444 10.6151
R1421 B.n446 B.n445 10.6151
R1422 B.n447 B.n446 10.6151
R1423 B.n449 B.n447 10.6151
R1424 B.n450 B.n449 10.6151
R1425 B.n451 B.n450 10.6151
R1426 B.n452 B.n451 10.6151
R1427 B.n454 B.n452 10.6151
R1428 B.n455 B.n454 10.6151
R1429 B.n456 B.n455 10.6151
R1430 B.n457 B.n456 10.6151
R1431 B.n459 B.n457 10.6151
R1432 B.n460 B.n459 10.6151
R1433 B.n461 B.n460 10.6151
R1434 B.n462 B.n461 10.6151
R1435 B.n464 B.n462 10.6151
R1436 B.n465 B.n464 10.6151
R1437 B.n466 B.n465 10.6151
R1438 B.n467 B.n466 10.6151
R1439 B.n469 B.n467 10.6151
R1440 B.n470 B.n469 10.6151
R1441 B.n471 B.n470 10.6151
R1442 B.n472 B.n471 10.6151
R1443 B.n343 B.n342 10.6151
R1444 B.n342 B.n159 10.6151
R1445 B.n337 B.n159 10.6151
R1446 B.n337 B.n336 10.6151
R1447 B.n336 B.n161 10.6151
R1448 B.n331 B.n161 10.6151
R1449 B.n331 B.n330 10.6151
R1450 B.n330 B.n329 10.6151
R1451 B.n329 B.n163 10.6151
R1452 B.n323 B.n163 10.6151
R1453 B.n323 B.n322 10.6151
R1454 B.n322 B.n321 10.6151
R1455 B.n321 B.n165 10.6151
R1456 B.n315 B.n165 10.6151
R1457 B.n315 B.n314 10.6151
R1458 B.n314 B.n313 10.6151
R1459 B.n313 B.n167 10.6151
R1460 B.n307 B.n167 10.6151
R1461 B.n307 B.n306 10.6151
R1462 B.n306 B.n305 10.6151
R1463 B.n305 B.n169 10.6151
R1464 B.n299 B.n169 10.6151
R1465 B.n299 B.n298 10.6151
R1466 B.n298 B.n297 10.6151
R1467 B.n297 B.n171 10.6151
R1468 B.n291 B.n171 10.6151
R1469 B.n291 B.n290 10.6151
R1470 B.n290 B.n289 10.6151
R1471 B.n289 B.n173 10.6151
R1472 B.n283 B.n173 10.6151
R1473 B.n283 B.n282 10.6151
R1474 B.n280 B.n177 10.6151
R1475 B.n274 B.n177 10.6151
R1476 B.n274 B.n273 10.6151
R1477 B.n273 B.n272 10.6151
R1478 B.n272 B.n179 10.6151
R1479 B.n266 B.n179 10.6151
R1480 B.n266 B.n265 10.6151
R1481 B.n265 B.n264 10.6151
R1482 B.n260 B.n259 10.6151
R1483 B.n259 B.n185 10.6151
R1484 B.n254 B.n185 10.6151
R1485 B.n254 B.n253 10.6151
R1486 B.n253 B.n252 10.6151
R1487 B.n252 B.n187 10.6151
R1488 B.n246 B.n187 10.6151
R1489 B.n246 B.n245 10.6151
R1490 B.n245 B.n244 10.6151
R1491 B.n244 B.n189 10.6151
R1492 B.n238 B.n189 10.6151
R1493 B.n238 B.n237 10.6151
R1494 B.n237 B.n236 10.6151
R1495 B.n236 B.n191 10.6151
R1496 B.n230 B.n191 10.6151
R1497 B.n230 B.n229 10.6151
R1498 B.n229 B.n228 10.6151
R1499 B.n228 B.n193 10.6151
R1500 B.n222 B.n193 10.6151
R1501 B.n222 B.n221 10.6151
R1502 B.n221 B.n220 10.6151
R1503 B.n220 B.n195 10.6151
R1504 B.n214 B.n195 10.6151
R1505 B.n214 B.n213 10.6151
R1506 B.n213 B.n212 10.6151
R1507 B.n212 B.n197 10.6151
R1508 B.n206 B.n197 10.6151
R1509 B.n206 B.n205 10.6151
R1510 B.n205 B.n204 10.6151
R1511 B.n204 B.n199 10.6151
R1512 B.n199 B.n155 10.6151
R1513 B.n344 B.n151 10.6151
R1514 B.n354 B.n151 10.6151
R1515 B.n355 B.n354 10.6151
R1516 B.n356 B.n355 10.6151
R1517 B.n356 B.n143 10.6151
R1518 B.n366 B.n143 10.6151
R1519 B.n367 B.n366 10.6151
R1520 B.n368 B.n367 10.6151
R1521 B.n368 B.n135 10.6151
R1522 B.n378 B.n135 10.6151
R1523 B.n379 B.n378 10.6151
R1524 B.n380 B.n379 10.6151
R1525 B.n380 B.n127 10.6151
R1526 B.n390 B.n127 10.6151
R1527 B.n391 B.n390 10.6151
R1528 B.n392 B.n391 10.6151
R1529 B.n392 B.n119 10.6151
R1530 B.n402 B.n119 10.6151
R1531 B.n403 B.n402 10.6151
R1532 B.n404 B.n403 10.6151
R1533 B.n404 B.n111 10.6151
R1534 B.n414 B.n111 10.6151
R1535 B.n415 B.n414 10.6151
R1536 B.n416 B.n415 10.6151
R1537 B.n416 B.n103 10.6151
R1538 B.n427 B.n103 10.6151
R1539 B.n428 B.n427 10.6151
R1540 B.n429 B.n428 10.6151
R1541 B.n429 B.n0 10.6151
R1542 B.n676 B.n1 10.6151
R1543 B.n676 B.n675 10.6151
R1544 B.n675 B.n674 10.6151
R1545 B.n674 B.n10 10.6151
R1546 B.n668 B.n10 10.6151
R1547 B.n668 B.n667 10.6151
R1548 B.n667 B.n666 10.6151
R1549 B.n666 B.n17 10.6151
R1550 B.n660 B.n17 10.6151
R1551 B.n660 B.n659 10.6151
R1552 B.n659 B.n658 10.6151
R1553 B.n658 B.n24 10.6151
R1554 B.n652 B.n24 10.6151
R1555 B.n652 B.n651 10.6151
R1556 B.n651 B.n650 10.6151
R1557 B.n650 B.n31 10.6151
R1558 B.n644 B.n31 10.6151
R1559 B.n644 B.n643 10.6151
R1560 B.n643 B.n642 10.6151
R1561 B.n642 B.n38 10.6151
R1562 B.n636 B.n38 10.6151
R1563 B.n636 B.n635 10.6151
R1564 B.n635 B.n634 10.6151
R1565 B.n634 B.n45 10.6151
R1566 B.n628 B.n45 10.6151
R1567 B.n628 B.n627 10.6151
R1568 B.n627 B.n626 10.6151
R1569 B.n626 B.n52 10.6151
R1570 B.n620 B.n52 10.6151
R1571 B.t3 B.n137 7.11512
R1572 B.n639 B.t7 7.11512
R1573 B.n555 B.n554 6.5566
R1574 B.n538 B.n537 6.5566
R1575 B.n281 B.n280 6.5566
R1576 B.n264 B.n183 6.5566
R1577 B.n556 B.n555 4.05904
R1578 B.n537 B.n536 4.05904
R1579 B.n282 B.n281 4.05904
R1580 B.n260 B.n183 4.05904
R1581 B.n682 B.n0 2.81026
R1582 B.n682 B.n1 2.81026
R1583 B.t1 B.n109 2.37204
R1584 B.t0 B.n15 2.37204
R1585 VN VN.t1 144.578
R1586 VN VN.t0 101.044
R1587 VDD2.n85 VDD2.n45 289.615
R1588 VDD2.n40 VDD2.n0 289.615
R1589 VDD2.n86 VDD2.n85 185
R1590 VDD2.n84 VDD2.n83 185
R1591 VDD2.n82 VDD2.n48 185
R1592 VDD2.n52 VDD2.n49 185
R1593 VDD2.n77 VDD2.n76 185
R1594 VDD2.n75 VDD2.n74 185
R1595 VDD2.n54 VDD2.n53 185
R1596 VDD2.n69 VDD2.n68 185
R1597 VDD2.n67 VDD2.n66 185
R1598 VDD2.n58 VDD2.n57 185
R1599 VDD2.n61 VDD2.n60 185
R1600 VDD2.n15 VDD2.n14 185
R1601 VDD2.n12 VDD2.n11 185
R1602 VDD2.n21 VDD2.n20 185
R1603 VDD2.n23 VDD2.n22 185
R1604 VDD2.n8 VDD2.n7 185
R1605 VDD2.n29 VDD2.n28 185
R1606 VDD2.n32 VDD2.n31 185
R1607 VDD2.n30 VDD2.n4 185
R1608 VDD2.n37 VDD2.n3 185
R1609 VDD2.n39 VDD2.n38 185
R1610 VDD2.n41 VDD2.n40 185
R1611 VDD2.t0 VDD2.n59 149.524
R1612 VDD2.t1 VDD2.n13 149.524
R1613 VDD2.n85 VDD2.n84 104.615
R1614 VDD2.n84 VDD2.n48 104.615
R1615 VDD2.n52 VDD2.n48 104.615
R1616 VDD2.n76 VDD2.n52 104.615
R1617 VDD2.n76 VDD2.n75 104.615
R1618 VDD2.n75 VDD2.n53 104.615
R1619 VDD2.n68 VDD2.n53 104.615
R1620 VDD2.n68 VDD2.n67 104.615
R1621 VDD2.n67 VDD2.n57 104.615
R1622 VDD2.n60 VDD2.n57 104.615
R1623 VDD2.n14 VDD2.n11 104.615
R1624 VDD2.n21 VDD2.n11 104.615
R1625 VDD2.n22 VDD2.n21 104.615
R1626 VDD2.n22 VDD2.n7 104.615
R1627 VDD2.n29 VDD2.n7 104.615
R1628 VDD2.n31 VDD2.n29 104.615
R1629 VDD2.n31 VDD2.n30 104.615
R1630 VDD2.n30 VDD2.n3 104.615
R1631 VDD2.n39 VDD2.n3 104.615
R1632 VDD2.n40 VDD2.n39 104.615
R1633 VDD2.n90 VDD2.n44 88.6784
R1634 VDD2.n60 VDD2.t0 52.3082
R1635 VDD2.n14 VDD2.t1 52.3082
R1636 VDD2.n90 VDD2.n89 51.1914
R1637 VDD2.n83 VDD2.n82 13.1884
R1638 VDD2.n38 VDD2.n37 13.1884
R1639 VDD2.n86 VDD2.n47 12.8005
R1640 VDD2.n81 VDD2.n49 12.8005
R1641 VDD2.n36 VDD2.n4 12.8005
R1642 VDD2.n41 VDD2.n2 12.8005
R1643 VDD2.n87 VDD2.n45 12.0247
R1644 VDD2.n78 VDD2.n77 12.0247
R1645 VDD2.n33 VDD2.n32 12.0247
R1646 VDD2.n42 VDD2.n0 12.0247
R1647 VDD2.n74 VDD2.n51 11.249
R1648 VDD2.n28 VDD2.n6 11.249
R1649 VDD2.n73 VDD2.n54 10.4732
R1650 VDD2.n27 VDD2.n8 10.4732
R1651 VDD2.n61 VDD2.n59 10.2747
R1652 VDD2.n15 VDD2.n13 10.2747
R1653 VDD2.n70 VDD2.n69 9.69747
R1654 VDD2.n24 VDD2.n23 9.69747
R1655 VDD2.n89 VDD2.n88 9.45567
R1656 VDD2.n44 VDD2.n43 9.45567
R1657 VDD2.n63 VDD2.n62 9.3005
R1658 VDD2.n65 VDD2.n64 9.3005
R1659 VDD2.n56 VDD2.n55 9.3005
R1660 VDD2.n71 VDD2.n70 9.3005
R1661 VDD2.n73 VDD2.n72 9.3005
R1662 VDD2.n51 VDD2.n50 9.3005
R1663 VDD2.n79 VDD2.n78 9.3005
R1664 VDD2.n81 VDD2.n80 9.3005
R1665 VDD2.n88 VDD2.n87 9.3005
R1666 VDD2.n47 VDD2.n46 9.3005
R1667 VDD2.n43 VDD2.n42 9.3005
R1668 VDD2.n2 VDD2.n1 9.3005
R1669 VDD2.n17 VDD2.n16 9.3005
R1670 VDD2.n19 VDD2.n18 9.3005
R1671 VDD2.n10 VDD2.n9 9.3005
R1672 VDD2.n25 VDD2.n24 9.3005
R1673 VDD2.n27 VDD2.n26 9.3005
R1674 VDD2.n6 VDD2.n5 9.3005
R1675 VDD2.n34 VDD2.n33 9.3005
R1676 VDD2.n36 VDD2.n35 9.3005
R1677 VDD2.n66 VDD2.n56 8.92171
R1678 VDD2.n20 VDD2.n10 8.92171
R1679 VDD2.n65 VDD2.n58 8.14595
R1680 VDD2.n19 VDD2.n12 8.14595
R1681 VDD2.n62 VDD2.n61 7.3702
R1682 VDD2.n16 VDD2.n15 7.3702
R1683 VDD2.n62 VDD2.n58 5.81868
R1684 VDD2.n16 VDD2.n12 5.81868
R1685 VDD2.n66 VDD2.n65 5.04292
R1686 VDD2.n20 VDD2.n19 5.04292
R1687 VDD2.n69 VDD2.n56 4.26717
R1688 VDD2.n23 VDD2.n10 4.26717
R1689 VDD2.n70 VDD2.n54 3.49141
R1690 VDD2.n24 VDD2.n8 3.49141
R1691 VDD2.n17 VDD2.n13 2.84303
R1692 VDD2.n63 VDD2.n59 2.84303
R1693 VDD2.n74 VDD2.n73 2.71565
R1694 VDD2.n28 VDD2.n27 2.71565
R1695 VDD2.n89 VDD2.n45 1.93989
R1696 VDD2.n77 VDD2.n51 1.93989
R1697 VDD2.n32 VDD2.n6 1.93989
R1698 VDD2.n44 VDD2.n0 1.93989
R1699 VDD2.n87 VDD2.n86 1.16414
R1700 VDD2.n78 VDD2.n49 1.16414
R1701 VDD2.n33 VDD2.n4 1.16414
R1702 VDD2.n42 VDD2.n41 1.16414
R1703 VDD2 VDD2.n90 0.856103
R1704 VDD2.n83 VDD2.n47 0.388379
R1705 VDD2.n82 VDD2.n81 0.388379
R1706 VDD2.n37 VDD2.n36 0.388379
R1707 VDD2.n38 VDD2.n2 0.388379
R1708 VDD2.n88 VDD2.n46 0.155672
R1709 VDD2.n80 VDD2.n46 0.155672
R1710 VDD2.n80 VDD2.n79 0.155672
R1711 VDD2.n79 VDD2.n50 0.155672
R1712 VDD2.n72 VDD2.n50 0.155672
R1713 VDD2.n72 VDD2.n71 0.155672
R1714 VDD2.n71 VDD2.n55 0.155672
R1715 VDD2.n64 VDD2.n55 0.155672
R1716 VDD2.n64 VDD2.n63 0.155672
R1717 VDD2.n18 VDD2.n17 0.155672
R1718 VDD2.n18 VDD2.n9 0.155672
R1719 VDD2.n25 VDD2.n9 0.155672
R1720 VDD2.n26 VDD2.n25 0.155672
R1721 VDD2.n26 VDD2.n5 0.155672
R1722 VDD2.n34 VDD2.n5 0.155672
R1723 VDD2.n35 VDD2.n34 0.155672
R1724 VDD2.n35 VDD2.n1 0.155672
R1725 VDD2.n43 VDD2.n1 0.155672
C0 VDD2 VTAIL 4.4165f
C1 VDD2 VDD1 0.768261f
C2 VTAIL VN 2.01804f
C3 VDD2 VP 0.364865f
C4 VDD1 VN 0.148141f
C5 VTAIL VDD1 4.35945f
C6 VP VN 5.1991f
C7 VTAIL VP 2.03224f
C8 VP VDD1 2.35976f
C9 VDD2 VN 2.14478f
C10 VDD2 B 4.097579f
C11 VDD1 B 6.80754f
C12 VTAIL B 6.356205f
C13 VN B 10.7161f
C14 VP B 7.135497f
C15 VDD2.n0 B 0.027822f
C16 VDD2.n1 B 0.020584f
C17 VDD2.n2 B 0.011061f
C18 VDD2.n3 B 0.026144f
C19 VDD2.n4 B 0.011712f
C20 VDD2.n5 B 0.020584f
C21 VDD2.n6 B 0.011061f
C22 VDD2.n7 B 0.026144f
C23 VDD2.n8 B 0.011712f
C24 VDD2.n9 B 0.020584f
C25 VDD2.n10 B 0.011061f
C26 VDD2.n11 B 0.026144f
C27 VDD2.n12 B 0.011712f
C28 VDD2.n13 B 0.121868f
C29 VDD2.t1 B 0.04379f
C30 VDD2.n14 B 0.019608f
C31 VDD2.n15 B 0.018482f
C32 VDD2.n16 B 0.011061f
C33 VDD2.n17 B 0.730782f
C34 VDD2.n18 B 0.020584f
C35 VDD2.n19 B 0.011061f
C36 VDD2.n20 B 0.011712f
C37 VDD2.n21 B 0.026144f
C38 VDD2.n22 B 0.026144f
C39 VDD2.n23 B 0.011712f
C40 VDD2.n24 B 0.011061f
C41 VDD2.n25 B 0.020584f
C42 VDD2.n26 B 0.020584f
C43 VDD2.n27 B 0.011061f
C44 VDD2.n28 B 0.011712f
C45 VDD2.n29 B 0.026144f
C46 VDD2.n30 B 0.026144f
C47 VDD2.n31 B 0.026144f
C48 VDD2.n32 B 0.011712f
C49 VDD2.n33 B 0.011061f
C50 VDD2.n34 B 0.020584f
C51 VDD2.n35 B 0.020584f
C52 VDD2.n36 B 0.011061f
C53 VDD2.n37 B 0.011386f
C54 VDD2.n38 B 0.011386f
C55 VDD2.n39 B 0.026144f
C56 VDD2.n40 B 0.054633f
C57 VDD2.n41 B 0.011712f
C58 VDD2.n42 B 0.011061f
C59 VDD2.n43 B 0.050953f
C60 VDD2.n44 B 0.536352f
C61 VDD2.n45 B 0.027822f
C62 VDD2.n46 B 0.020584f
C63 VDD2.n47 B 0.011061f
C64 VDD2.n48 B 0.026144f
C65 VDD2.n49 B 0.011712f
C66 VDD2.n50 B 0.020584f
C67 VDD2.n51 B 0.011061f
C68 VDD2.n52 B 0.026144f
C69 VDD2.n53 B 0.026144f
C70 VDD2.n54 B 0.011712f
C71 VDD2.n55 B 0.020584f
C72 VDD2.n56 B 0.011061f
C73 VDD2.n57 B 0.026144f
C74 VDD2.n58 B 0.011712f
C75 VDD2.n59 B 0.121868f
C76 VDD2.t0 B 0.04379f
C77 VDD2.n60 B 0.019608f
C78 VDD2.n61 B 0.018482f
C79 VDD2.n62 B 0.011061f
C80 VDD2.n63 B 0.730782f
C81 VDD2.n64 B 0.020584f
C82 VDD2.n65 B 0.011061f
C83 VDD2.n66 B 0.011712f
C84 VDD2.n67 B 0.026144f
C85 VDD2.n68 B 0.026144f
C86 VDD2.n69 B 0.011712f
C87 VDD2.n70 B 0.011061f
C88 VDD2.n71 B 0.020584f
C89 VDD2.n72 B 0.020584f
C90 VDD2.n73 B 0.011061f
C91 VDD2.n74 B 0.011712f
C92 VDD2.n75 B 0.026144f
C93 VDD2.n76 B 0.026144f
C94 VDD2.n77 B 0.011712f
C95 VDD2.n78 B 0.011061f
C96 VDD2.n79 B 0.020584f
C97 VDD2.n80 B 0.020584f
C98 VDD2.n81 B 0.011061f
C99 VDD2.n82 B 0.011386f
C100 VDD2.n83 B 0.011386f
C101 VDD2.n84 B 0.026144f
C102 VDD2.n85 B 0.054633f
C103 VDD2.n86 B 0.011712f
C104 VDD2.n87 B 0.011061f
C105 VDD2.n88 B 0.050953f
C106 VDD2.n89 B 0.044656f
C107 VDD2.n90 B 2.36593f
C108 VN.t0 B 2.56055f
C109 VN.t1 B 3.18627f
C110 VDD1.n0 B 0.028769f
C111 VDD1.n1 B 0.021285f
C112 VDD1.n2 B 0.011438f
C113 VDD1.n3 B 0.027035f
C114 VDD1.n4 B 0.012111f
C115 VDD1.n5 B 0.021285f
C116 VDD1.n6 B 0.011438f
C117 VDD1.n7 B 0.027035f
C118 VDD1.n8 B 0.027035f
C119 VDD1.n9 B 0.012111f
C120 VDD1.n10 B 0.021285f
C121 VDD1.n11 B 0.011438f
C122 VDD1.n12 B 0.027035f
C123 VDD1.n13 B 0.012111f
C124 VDD1.n14 B 0.126019f
C125 VDD1.t0 B 0.045282f
C126 VDD1.n15 B 0.020276f
C127 VDD1.n16 B 0.019111f
C128 VDD1.n17 B 0.011438f
C129 VDD1.n18 B 0.755672f
C130 VDD1.n19 B 0.021285f
C131 VDD1.n20 B 0.011438f
C132 VDD1.n21 B 0.012111f
C133 VDD1.n22 B 0.027035f
C134 VDD1.n23 B 0.027035f
C135 VDD1.n24 B 0.012111f
C136 VDD1.n25 B 0.011438f
C137 VDD1.n26 B 0.021285f
C138 VDD1.n27 B 0.021285f
C139 VDD1.n28 B 0.011438f
C140 VDD1.n29 B 0.012111f
C141 VDD1.n30 B 0.027035f
C142 VDD1.n31 B 0.027035f
C143 VDD1.n32 B 0.012111f
C144 VDD1.n33 B 0.011438f
C145 VDD1.n34 B 0.021285f
C146 VDD1.n35 B 0.021285f
C147 VDD1.n36 B 0.011438f
C148 VDD1.n37 B 0.011774f
C149 VDD1.n38 B 0.011774f
C150 VDD1.n39 B 0.027035f
C151 VDD1.n40 B 0.056493f
C152 VDD1.n41 B 0.012111f
C153 VDD1.n42 B 0.011438f
C154 VDD1.n43 B 0.052689f
C155 VDD1.n44 B 0.047848f
C156 VDD1.n45 B 0.028769f
C157 VDD1.n46 B 0.021285f
C158 VDD1.n47 B 0.011438f
C159 VDD1.n48 B 0.027035f
C160 VDD1.n49 B 0.012111f
C161 VDD1.n50 B 0.021285f
C162 VDD1.n51 B 0.011438f
C163 VDD1.n52 B 0.027035f
C164 VDD1.n53 B 0.012111f
C165 VDD1.n54 B 0.021285f
C166 VDD1.n55 B 0.011438f
C167 VDD1.n56 B 0.027035f
C168 VDD1.n57 B 0.012111f
C169 VDD1.n58 B 0.126019f
C170 VDD1.t1 B 0.045282f
C171 VDD1.n59 B 0.020276f
C172 VDD1.n60 B 0.019111f
C173 VDD1.n61 B 0.011438f
C174 VDD1.n62 B 0.755672f
C175 VDD1.n63 B 0.021285f
C176 VDD1.n64 B 0.011438f
C177 VDD1.n65 B 0.012111f
C178 VDD1.n66 B 0.027035f
C179 VDD1.n67 B 0.027035f
C180 VDD1.n68 B 0.012111f
C181 VDD1.n69 B 0.011438f
C182 VDD1.n70 B 0.021285f
C183 VDD1.n71 B 0.021285f
C184 VDD1.n72 B 0.011438f
C185 VDD1.n73 B 0.012111f
C186 VDD1.n74 B 0.027035f
C187 VDD1.n75 B 0.027035f
C188 VDD1.n76 B 0.027035f
C189 VDD1.n77 B 0.012111f
C190 VDD1.n78 B 0.011438f
C191 VDD1.n79 B 0.021285f
C192 VDD1.n80 B 0.021285f
C193 VDD1.n81 B 0.011438f
C194 VDD1.n82 B 0.011774f
C195 VDD1.n83 B 0.011774f
C196 VDD1.n84 B 0.027035f
C197 VDD1.n85 B 0.056493f
C198 VDD1.n86 B 0.012111f
C199 VDD1.n87 B 0.011438f
C200 VDD1.n88 B 0.052689f
C201 VDD1.n89 B 0.598503f
C202 VTAIL.n0 B 0.029948f
C203 VTAIL.n1 B 0.022157f
C204 VTAIL.n2 B 0.011906f
C205 VTAIL.n3 B 0.028142f
C206 VTAIL.n4 B 0.012606f
C207 VTAIL.n5 B 0.022157f
C208 VTAIL.n6 B 0.011906f
C209 VTAIL.n7 B 0.028142f
C210 VTAIL.n8 B 0.012606f
C211 VTAIL.n9 B 0.022157f
C212 VTAIL.n10 B 0.011906f
C213 VTAIL.n11 B 0.028142f
C214 VTAIL.n12 B 0.012606f
C215 VTAIL.n13 B 0.13118f
C216 VTAIL.t2 B 0.047136f
C217 VTAIL.n14 B 0.021106f
C218 VTAIL.n15 B 0.019894f
C219 VTAIL.n16 B 0.011906f
C220 VTAIL.n17 B 0.786623f
C221 VTAIL.n18 B 0.022157f
C222 VTAIL.n19 B 0.011906f
C223 VTAIL.n20 B 0.012606f
C224 VTAIL.n21 B 0.028142f
C225 VTAIL.n22 B 0.028142f
C226 VTAIL.n23 B 0.012606f
C227 VTAIL.n24 B 0.011906f
C228 VTAIL.n25 B 0.022157f
C229 VTAIL.n26 B 0.022157f
C230 VTAIL.n27 B 0.011906f
C231 VTAIL.n28 B 0.012606f
C232 VTAIL.n29 B 0.028142f
C233 VTAIL.n30 B 0.028142f
C234 VTAIL.n31 B 0.028142f
C235 VTAIL.n32 B 0.012606f
C236 VTAIL.n33 B 0.011906f
C237 VTAIL.n34 B 0.022157f
C238 VTAIL.n35 B 0.022157f
C239 VTAIL.n36 B 0.011906f
C240 VTAIL.n37 B 0.012256f
C241 VTAIL.n38 B 0.012256f
C242 VTAIL.n39 B 0.028142f
C243 VTAIL.n40 B 0.058807f
C244 VTAIL.n41 B 0.012606f
C245 VTAIL.n42 B 0.011906f
C246 VTAIL.n43 B 0.054847f
C247 VTAIL.n44 B 0.032796f
C248 VTAIL.n45 B 1.40379f
C249 VTAIL.n46 B 0.029948f
C250 VTAIL.n47 B 0.022157f
C251 VTAIL.n48 B 0.011906f
C252 VTAIL.n49 B 0.028142f
C253 VTAIL.n50 B 0.012606f
C254 VTAIL.n51 B 0.022157f
C255 VTAIL.n52 B 0.011906f
C256 VTAIL.n53 B 0.028142f
C257 VTAIL.n54 B 0.028142f
C258 VTAIL.n55 B 0.012606f
C259 VTAIL.n56 B 0.022157f
C260 VTAIL.n57 B 0.011906f
C261 VTAIL.n58 B 0.028142f
C262 VTAIL.n59 B 0.012606f
C263 VTAIL.n60 B 0.13118f
C264 VTAIL.t1 B 0.047136f
C265 VTAIL.n61 B 0.021106f
C266 VTAIL.n62 B 0.019894f
C267 VTAIL.n63 B 0.011906f
C268 VTAIL.n64 B 0.786623f
C269 VTAIL.n65 B 0.022157f
C270 VTAIL.n66 B 0.011906f
C271 VTAIL.n67 B 0.012606f
C272 VTAIL.n68 B 0.028142f
C273 VTAIL.n69 B 0.028142f
C274 VTAIL.n70 B 0.012606f
C275 VTAIL.n71 B 0.011906f
C276 VTAIL.n72 B 0.022157f
C277 VTAIL.n73 B 0.022157f
C278 VTAIL.n74 B 0.011906f
C279 VTAIL.n75 B 0.012606f
C280 VTAIL.n76 B 0.028142f
C281 VTAIL.n77 B 0.028142f
C282 VTAIL.n78 B 0.012606f
C283 VTAIL.n79 B 0.011906f
C284 VTAIL.n80 B 0.022157f
C285 VTAIL.n81 B 0.022157f
C286 VTAIL.n82 B 0.011906f
C287 VTAIL.n83 B 0.012256f
C288 VTAIL.n84 B 0.012256f
C289 VTAIL.n85 B 0.028142f
C290 VTAIL.n86 B 0.058807f
C291 VTAIL.n87 B 0.012606f
C292 VTAIL.n88 B 0.011906f
C293 VTAIL.n89 B 0.054847f
C294 VTAIL.n90 B 0.032796f
C295 VTAIL.n91 B 1.45657f
C296 VTAIL.n92 B 0.029948f
C297 VTAIL.n93 B 0.022157f
C298 VTAIL.n94 B 0.011906f
C299 VTAIL.n95 B 0.028142f
C300 VTAIL.n96 B 0.012606f
C301 VTAIL.n97 B 0.022157f
C302 VTAIL.n98 B 0.011906f
C303 VTAIL.n99 B 0.028142f
C304 VTAIL.n100 B 0.028142f
C305 VTAIL.n101 B 0.012606f
C306 VTAIL.n102 B 0.022157f
C307 VTAIL.n103 B 0.011906f
C308 VTAIL.n104 B 0.028142f
C309 VTAIL.n105 B 0.012606f
C310 VTAIL.n106 B 0.13118f
C311 VTAIL.t3 B 0.047136f
C312 VTAIL.n107 B 0.021106f
C313 VTAIL.n108 B 0.019894f
C314 VTAIL.n109 B 0.011906f
C315 VTAIL.n110 B 0.786623f
C316 VTAIL.n111 B 0.022157f
C317 VTAIL.n112 B 0.011906f
C318 VTAIL.n113 B 0.012606f
C319 VTAIL.n114 B 0.028142f
C320 VTAIL.n115 B 0.028142f
C321 VTAIL.n116 B 0.012606f
C322 VTAIL.n117 B 0.011906f
C323 VTAIL.n118 B 0.022157f
C324 VTAIL.n119 B 0.022157f
C325 VTAIL.n120 B 0.011906f
C326 VTAIL.n121 B 0.012606f
C327 VTAIL.n122 B 0.028142f
C328 VTAIL.n123 B 0.028142f
C329 VTAIL.n124 B 0.012606f
C330 VTAIL.n125 B 0.011906f
C331 VTAIL.n126 B 0.022157f
C332 VTAIL.n127 B 0.022157f
C333 VTAIL.n128 B 0.011906f
C334 VTAIL.n129 B 0.012256f
C335 VTAIL.n130 B 0.012256f
C336 VTAIL.n131 B 0.028142f
C337 VTAIL.n132 B 0.058807f
C338 VTAIL.n133 B 0.012606f
C339 VTAIL.n134 B 0.011906f
C340 VTAIL.n135 B 0.054847f
C341 VTAIL.n136 B 0.032796f
C342 VTAIL.n137 B 1.22884f
C343 VTAIL.n138 B 0.029948f
C344 VTAIL.n139 B 0.022157f
C345 VTAIL.n140 B 0.011906f
C346 VTAIL.n141 B 0.028142f
C347 VTAIL.n142 B 0.012606f
C348 VTAIL.n143 B 0.022157f
C349 VTAIL.n144 B 0.011906f
C350 VTAIL.n145 B 0.028142f
C351 VTAIL.n146 B 0.012606f
C352 VTAIL.n147 B 0.022157f
C353 VTAIL.n148 B 0.011906f
C354 VTAIL.n149 B 0.028142f
C355 VTAIL.n150 B 0.012606f
C356 VTAIL.n151 B 0.13118f
C357 VTAIL.t0 B 0.047136f
C358 VTAIL.n152 B 0.021106f
C359 VTAIL.n153 B 0.019894f
C360 VTAIL.n154 B 0.011906f
C361 VTAIL.n155 B 0.786623f
C362 VTAIL.n156 B 0.022157f
C363 VTAIL.n157 B 0.011906f
C364 VTAIL.n158 B 0.012606f
C365 VTAIL.n159 B 0.028142f
C366 VTAIL.n160 B 0.028142f
C367 VTAIL.n161 B 0.012606f
C368 VTAIL.n162 B 0.011906f
C369 VTAIL.n163 B 0.022157f
C370 VTAIL.n164 B 0.022157f
C371 VTAIL.n165 B 0.011906f
C372 VTAIL.n166 B 0.012606f
C373 VTAIL.n167 B 0.028142f
C374 VTAIL.n168 B 0.028142f
C375 VTAIL.n169 B 0.028142f
C376 VTAIL.n170 B 0.012606f
C377 VTAIL.n171 B 0.011906f
C378 VTAIL.n172 B 0.022157f
C379 VTAIL.n173 B 0.022157f
C380 VTAIL.n174 B 0.011906f
C381 VTAIL.n175 B 0.012256f
C382 VTAIL.n176 B 0.012256f
C383 VTAIL.n177 B 0.028142f
C384 VTAIL.n178 B 0.058807f
C385 VTAIL.n179 B 0.012606f
C386 VTAIL.n180 B 0.011906f
C387 VTAIL.n181 B 0.054847f
C388 VTAIL.n182 B 0.032796f
C389 VTAIL.n183 B 1.13422f
C390 VP.t1 B 3.30258f
C391 VP.t0 B 2.64995f
C392 VP.n0 B 3.54453f
.ends

