* NGSPICE file created from diff_pair_sample_0125.ext - technology: sky130A

.subckt diff_pair_sample_0125 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t2 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X1 VDD1.t9 VP.t0 VTAIL.t7 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=4.1925 ps=22.28 w=10.75 l=3.09
X2 VTAIL.t17 VN.t1 VDD2.t8 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X3 VTAIL.t16 VN.t2 VDD2.t9 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X4 VDD2.t1 VN.t3 VTAIL.t15 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=4.1925 ps=22.28 w=10.75 l=3.09
X5 VDD2.t0 VN.t4 VTAIL.t14 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=4.1925 ps=22.28 w=10.75 l=3.09
X6 VDD2.t3 VN.t5 VTAIL.t13 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=1.77375 ps=11.08 w=10.75 l=3.09
X7 VTAIL.t2 VP.t1 VDD1.t8 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X8 VDD1.t7 VP.t2 VTAIL.t4 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=1.77375 ps=11.08 w=10.75 l=3.09
X9 VTAIL.t12 VN.t6 VDD2.t6 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X10 VDD1.t6 VP.t3 VTAIL.t0 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X11 VTAIL.t8 VP.t4 VDD1.t5 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X12 VTAIL.t5 VP.t5 VDD1.t4 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X13 VDD1.t3 VP.t6 VTAIL.t3 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=1.77375 ps=11.08 w=10.75 l=3.09
X14 VDD1.t2 VP.t7 VTAIL.t6 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X15 B.t11 B.t9 B.t10 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=0 ps=0 w=10.75 l=3.09
X16 VDD2.t4 VN.t7 VTAIL.t11 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X17 B.t8 B.t6 B.t7 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=0 ps=0 w=10.75 l=3.09
X18 VDD1.t1 VP.t8 VTAIL.t19 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=4.1925 ps=22.28 w=10.75 l=3.09
X19 B.t5 B.t3 B.t4 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=0 ps=0 w=10.75 l=3.09
X20 VDD2.t7 VN.t8 VTAIL.t10 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X21 VTAIL.t1 VP.t9 VDD1.t0 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=1.77375 pd=11.08 as=1.77375 ps=11.08 w=10.75 l=3.09
X22 B.t2 B.t0 B.t1 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=0 ps=0 w=10.75 l=3.09
X23 VDD2.t5 VN.t9 VTAIL.t9 w_n5074_n3118# sky130_fd_pr__pfet_01v8 ad=4.1925 pd=22.28 as=1.77375 ps=11.08 w=10.75 l=3.09
R0 VN.n88 VN.n87 161.3
R1 VN.n86 VN.n46 161.3
R2 VN.n85 VN.n84 161.3
R3 VN.n83 VN.n47 161.3
R4 VN.n82 VN.n81 161.3
R5 VN.n80 VN.n48 161.3
R6 VN.n79 VN.n78 161.3
R7 VN.n77 VN.n76 161.3
R8 VN.n75 VN.n50 161.3
R9 VN.n74 VN.n73 161.3
R10 VN.n72 VN.n51 161.3
R11 VN.n71 VN.n70 161.3
R12 VN.n69 VN.n52 161.3
R13 VN.n68 VN.n67 161.3
R14 VN.n66 VN.n53 161.3
R15 VN.n65 VN.n64 161.3
R16 VN.n63 VN.n54 161.3
R17 VN.n62 VN.n61 161.3
R18 VN.n60 VN.n55 161.3
R19 VN.n59 VN.n58 161.3
R20 VN.n43 VN.n42 161.3
R21 VN.n41 VN.n1 161.3
R22 VN.n40 VN.n39 161.3
R23 VN.n38 VN.n2 161.3
R24 VN.n37 VN.n36 161.3
R25 VN.n35 VN.n3 161.3
R26 VN.n34 VN.n33 161.3
R27 VN.n32 VN.n31 161.3
R28 VN.n30 VN.n5 161.3
R29 VN.n29 VN.n28 161.3
R30 VN.n27 VN.n6 161.3
R31 VN.n26 VN.n25 161.3
R32 VN.n24 VN.n7 161.3
R33 VN.n23 VN.n22 161.3
R34 VN.n21 VN.n8 161.3
R35 VN.n20 VN.n19 161.3
R36 VN.n18 VN.n9 161.3
R37 VN.n17 VN.n16 161.3
R38 VN.n15 VN.n10 161.3
R39 VN.n14 VN.n13 161.3
R40 VN.n56 VN.t3 117.066
R41 VN.n11 VN.t9 117.066
R42 VN.n23 VN.t8 83.8435
R43 VN.n12 VN.t1 83.8435
R44 VN.n4 VN.t0 83.8435
R45 VN.n0 VN.t4 83.8435
R46 VN.n68 VN.t7 83.8435
R47 VN.n57 VN.t6 83.8435
R48 VN.n49 VN.t2 83.8435
R49 VN.n45 VN.t5 83.8435
R50 VN.n44 VN.n0 73.4298
R51 VN.n89 VN.n45 73.4298
R52 VN.n18 VN.n17 56.5193
R53 VN.n29 VN.n6 56.5193
R54 VN.n63 VN.n62 56.5193
R55 VN.n74 VN.n51 56.5193
R56 VN VN.n89 55.0889
R57 VN.n12 VN.n11 53.3325
R58 VN.n57 VN.n56 53.3325
R59 VN.n40 VN.n2 53.1199
R60 VN.n85 VN.n47 53.1199
R61 VN.n36 VN.n2 27.8669
R62 VN.n81 VN.n47 27.8669
R63 VN.n13 VN.n10 24.4675
R64 VN.n17 VN.n10 24.4675
R65 VN.n19 VN.n18 24.4675
R66 VN.n19 VN.n8 24.4675
R67 VN.n23 VN.n8 24.4675
R68 VN.n24 VN.n23 24.4675
R69 VN.n25 VN.n24 24.4675
R70 VN.n25 VN.n6 24.4675
R71 VN.n30 VN.n29 24.4675
R72 VN.n31 VN.n30 24.4675
R73 VN.n35 VN.n34 24.4675
R74 VN.n36 VN.n35 24.4675
R75 VN.n41 VN.n40 24.4675
R76 VN.n42 VN.n41 24.4675
R77 VN.n62 VN.n55 24.4675
R78 VN.n58 VN.n55 24.4675
R79 VN.n70 VN.n51 24.4675
R80 VN.n70 VN.n69 24.4675
R81 VN.n69 VN.n68 24.4675
R82 VN.n68 VN.n53 24.4675
R83 VN.n64 VN.n53 24.4675
R84 VN.n64 VN.n63 24.4675
R85 VN.n81 VN.n80 24.4675
R86 VN.n80 VN.n79 24.4675
R87 VN.n76 VN.n75 24.4675
R88 VN.n75 VN.n74 24.4675
R89 VN.n87 VN.n86 24.4675
R90 VN.n86 VN.n85 24.4675
R91 VN.n13 VN.n12 20.5528
R92 VN.n31 VN.n4 20.5528
R93 VN.n58 VN.n57 20.5528
R94 VN.n76 VN.n49 20.5528
R95 VN.n42 VN.n0 16.6381
R96 VN.n87 VN.n45 16.6381
R97 VN.n59 VN.n56 4.07053
R98 VN.n14 VN.n11 4.07053
R99 VN.n34 VN.n4 3.91522
R100 VN.n79 VN.n49 3.91522
R101 VN.n89 VN.n88 0.354971
R102 VN.n44 VN.n43 0.354971
R103 VN VN.n44 0.26696
R104 VN.n88 VN.n46 0.189894
R105 VN.n84 VN.n46 0.189894
R106 VN.n84 VN.n83 0.189894
R107 VN.n83 VN.n82 0.189894
R108 VN.n82 VN.n48 0.189894
R109 VN.n78 VN.n48 0.189894
R110 VN.n78 VN.n77 0.189894
R111 VN.n77 VN.n50 0.189894
R112 VN.n73 VN.n50 0.189894
R113 VN.n73 VN.n72 0.189894
R114 VN.n72 VN.n71 0.189894
R115 VN.n71 VN.n52 0.189894
R116 VN.n67 VN.n52 0.189894
R117 VN.n67 VN.n66 0.189894
R118 VN.n66 VN.n65 0.189894
R119 VN.n65 VN.n54 0.189894
R120 VN.n61 VN.n54 0.189894
R121 VN.n61 VN.n60 0.189894
R122 VN.n60 VN.n59 0.189894
R123 VN.n15 VN.n14 0.189894
R124 VN.n16 VN.n15 0.189894
R125 VN.n16 VN.n9 0.189894
R126 VN.n20 VN.n9 0.189894
R127 VN.n21 VN.n20 0.189894
R128 VN.n22 VN.n21 0.189894
R129 VN.n22 VN.n7 0.189894
R130 VN.n26 VN.n7 0.189894
R131 VN.n27 VN.n26 0.189894
R132 VN.n28 VN.n27 0.189894
R133 VN.n28 VN.n5 0.189894
R134 VN.n32 VN.n5 0.189894
R135 VN.n33 VN.n32 0.189894
R136 VN.n33 VN.n3 0.189894
R137 VN.n37 VN.n3 0.189894
R138 VN.n38 VN.n37 0.189894
R139 VN.n39 VN.n38 0.189894
R140 VN.n39 VN.n1 0.189894
R141 VN.n43 VN.n1 0.189894
R142 VDD2.n113 VDD2.n61 756.745
R143 VDD2.n52 VDD2.n0 756.745
R144 VDD2.n114 VDD2.n113 585
R145 VDD2.n112 VDD2.n111 585
R146 VDD2.n65 VDD2.n64 585
R147 VDD2.n106 VDD2.n105 585
R148 VDD2.n104 VDD2.n103 585
R149 VDD2.n102 VDD2.n68 585
R150 VDD2.n72 VDD2.n69 585
R151 VDD2.n97 VDD2.n96 585
R152 VDD2.n95 VDD2.n94 585
R153 VDD2.n74 VDD2.n73 585
R154 VDD2.n89 VDD2.n88 585
R155 VDD2.n87 VDD2.n86 585
R156 VDD2.n78 VDD2.n77 585
R157 VDD2.n81 VDD2.n80 585
R158 VDD2.n19 VDD2.n18 585
R159 VDD2.n16 VDD2.n15 585
R160 VDD2.n25 VDD2.n24 585
R161 VDD2.n27 VDD2.n26 585
R162 VDD2.n12 VDD2.n11 585
R163 VDD2.n33 VDD2.n32 585
R164 VDD2.n36 VDD2.n35 585
R165 VDD2.n34 VDD2.n8 585
R166 VDD2.n41 VDD2.n7 585
R167 VDD2.n43 VDD2.n42 585
R168 VDD2.n45 VDD2.n44 585
R169 VDD2.n4 VDD2.n3 585
R170 VDD2.n51 VDD2.n50 585
R171 VDD2.n53 VDD2.n52 585
R172 VDD2.t3 VDD2.n79 329.038
R173 VDD2.t5 VDD2.n17 329.038
R174 VDD2.n113 VDD2.n112 171.744
R175 VDD2.n112 VDD2.n64 171.744
R176 VDD2.n105 VDD2.n64 171.744
R177 VDD2.n105 VDD2.n104 171.744
R178 VDD2.n104 VDD2.n68 171.744
R179 VDD2.n72 VDD2.n68 171.744
R180 VDD2.n96 VDD2.n72 171.744
R181 VDD2.n96 VDD2.n95 171.744
R182 VDD2.n95 VDD2.n73 171.744
R183 VDD2.n88 VDD2.n73 171.744
R184 VDD2.n88 VDD2.n87 171.744
R185 VDD2.n87 VDD2.n77 171.744
R186 VDD2.n80 VDD2.n77 171.744
R187 VDD2.n18 VDD2.n15 171.744
R188 VDD2.n25 VDD2.n15 171.744
R189 VDD2.n26 VDD2.n25 171.744
R190 VDD2.n26 VDD2.n11 171.744
R191 VDD2.n33 VDD2.n11 171.744
R192 VDD2.n35 VDD2.n33 171.744
R193 VDD2.n35 VDD2.n34 171.744
R194 VDD2.n34 VDD2.n7 171.744
R195 VDD2.n43 VDD2.n7 171.744
R196 VDD2.n44 VDD2.n43 171.744
R197 VDD2.n44 VDD2.n3 171.744
R198 VDD2.n51 VDD2.n3 171.744
R199 VDD2.n52 VDD2.n51 171.744
R200 VDD2.n80 VDD2.t3 85.8723
R201 VDD2.n18 VDD2.t5 85.8723
R202 VDD2.n60 VDD2.n59 79.3794
R203 VDD2 VDD2.n121 79.3766
R204 VDD2.n120 VDD2.n119 77.2237
R205 VDD2.n58 VDD2.n57 77.2235
R206 VDD2.n58 VDD2.n56 53.17
R207 VDD2.n118 VDD2.n117 50.2217
R208 VDD2.n118 VDD2.n60 46.9868
R209 VDD2.n103 VDD2.n102 13.1884
R210 VDD2.n42 VDD2.n41 13.1884
R211 VDD2.n106 VDD2.n67 12.8005
R212 VDD2.n101 VDD2.n69 12.8005
R213 VDD2.n40 VDD2.n8 12.8005
R214 VDD2.n45 VDD2.n6 12.8005
R215 VDD2.n107 VDD2.n65 12.0247
R216 VDD2.n98 VDD2.n97 12.0247
R217 VDD2.n37 VDD2.n36 12.0247
R218 VDD2.n46 VDD2.n4 12.0247
R219 VDD2.n111 VDD2.n110 11.249
R220 VDD2.n94 VDD2.n71 11.249
R221 VDD2.n32 VDD2.n10 11.249
R222 VDD2.n50 VDD2.n49 11.249
R223 VDD2.n81 VDD2.n79 10.7239
R224 VDD2.n19 VDD2.n17 10.7239
R225 VDD2.n114 VDD2.n63 10.4732
R226 VDD2.n93 VDD2.n74 10.4732
R227 VDD2.n31 VDD2.n12 10.4732
R228 VDD2.n53 VDD2.n2 10.4732
R229 VDD2.n115 VDD2.n61 9.69747
R230 VDD2.n90 VDD2.n89 9.69747
R231 VDD2.n28 VDD2.n27 9.69747
R232 VDD2.n54 VDD2.n0 9.69747
R233 VDD2.n117 VDD2.n116 9.45567
R234 VDD2.n56 VDD2.n55 9.45567
R235 VDD2.n83 VDD2.n82 9.3005
R236 VDD2.n85 VDD2.n84 9.3005
R237 VDD2.n76 VDD2.n75 9.3005
R238 VDD2.n91 VDD2.n90 9.3005
R239 VDD2.n93 VDD2.n92 9.3005
R240 VDD2.n71 VDD2.n70 9.3005
R241 VDD2.n99 VDD2.n98 9.3005
R242 VDD2.n101 VDD2.n100 9.3005
R243 VDD2.n116 VDD2.n115 9.3005
R244 VDD2.n63 VDD2.n62 9.3005
R245 VDD2.n110 VDD2.n109 9.3005
R246 VDD2.n108 VDD2.n107 9.3005
R247 VDD2.n67 VDD2.n66 9.3005
R248 VDD2.n55 VDD2.n54 9.3005
R249 VDD2.n2 VDD2.n1 9.3005
R250 VDD2.n49 VDD2.n48 9.3005
R251 VDD2.n47 VDD2.n46 9.3005
R252 VDD2.n6 VDD2.n5 9.3005
R253 VDD2.n21 VDD2.n20 9.3005
R254 VDD2.n23 VDD2.n22 9.3005
R255 VDD2.n14 VDD2.n13 9.3005
R256 VDD2.n29 VDD2.n28 9.3005
R257 VDD2.n31 VDD2.n30 9.3005
R258 VDD2.n10 VDD2.n9 9.3005
R259 VDD2.n38 VDD2.n37 9.3005
R260 VDD2.n40 VDD2.n39 9.3005
R261 VDD2.n86 VDD2.n76 8.92171
R262 VDD2.n24 VDD2.n14 8.92171
R263 VDD2.n85 VDD2.n78 8.14595
R264 VDD2.n23 VDD2.n16 8.14595
R265 VDD2.n82 VDD2.n81 7.3702
R266 VDD2.n20 VDD2.n19 7.3702
R267 VDD2.n82 VDD2.n78 5.81868
R268 VDD2.n20 VDD2.n16 5.81868
R269 VDD2.n86 VDD2.n85 5.04292
R270 VDD2.n24 VDD2.n23 5.04292
R271 VDD2.n117 VDD2.n61 4.26717
R272 VDD2.n89 VDD2.n76 4.26717
R273 VDD2.n27 VDD2.n14 4.26717
R274 VDD2.n56 VDD2.n0 4.26717
R275 VDD2.n115 VDD2.n114 3.49141
R276 VDD2.n90 VDD2.n74 3.49141
R277 VDD2.n28 VDD2.n12 3.49141
R278 VDD2.n54 VDD2.n53 3.49141
R279 VDD2.n121 VDD2.t6 3.02422
R280 VDD2.n121 VDD2.t1 3.02422
R281 VDD2.n119 VDD2.t9 3.02422
R282 VDD2.n119 VDD2.t4 3.02422
R283 VDD2.n59 VDD2.t2 3.02422
R284 VDD2.n59 VDD2.t0 3.02422
R285 VDD2.n57 VDD2.t8 3.02422
R286 VDD2.n57 VDD2.t7 3.02422
R287 VDD2.n120 VDD2.n118 2.94878
R288 VDD2.n111 VDD2.n63 2.71565
R289 VDD2.n94 VDD2.n93 2.71565
R290 VDD2.n32 VDD2.n31 2.71565
R291 VDD2.n50 VDD2.n2 2.71565
R292 VDD2.n83 VDD2.n79 2.41282
R293 VDD2.n21 VDD2.n17 2.41282
R294 VDD2.n110 VDD2.n65 1.93989
R295 VDD2.n97 VDD2.n71 1.93989
R296 VDD2.n36 VDD2.n10 1.93989
R297 VDD2.n49 VDD2.n4 1.93989
R298 VDD2.n107 VDD2.n106 1.16414
R299 VDD2.n98 VDD2.n69 1.16414
R300 VDD2.n37 VDD2.n8 1.16414
R301 VDD2.n46 VDD2.n45 1.16414
R302 VDD2 VDD2.n120 0.795759
R303 VDD2.n60 VDD2.n58 0.682223
R304 VDD2.n103 VDD2.n67 0.388379
R305 VDD2.n102 VDD2.n101 0.388379
R306 VDD2.n41 VDD2.n40 0.388379
R307 VDD2.n42 VDD2.n6 0.388379
R308 VDD2.n116 VDD2.n62 0.155672
R309 VDD2.n109 VDD2.n62 0.155672
R310 VDD2.n109 VDD2.n108 0.155672
R311 VDD2.n108 VDD2.n66 0.155672
R312 VDD2.n100 VDD2.n66 0.155672
R313 VDD2.n100 VDD2.n99 0.155672
R314 VDD2.n99 VDD2.n70 0.155672
R315 VDD2.n92 VDD2.n70 0.155672
R316 VDD2.n92 VDD2.n91 0.155672
R317 VDD2.n91 VDD2.n75 0.155672
R318 VDD2.n84 VDD2.n75 0.155672
R319 VDD2.n84 VDD2.n83 0.155672
R320 VDD2.n22 VDD2.n21 0.155672
R321 VDD2.n22 VDD2.n13 0.155672
R322 VDD2.n29 VDD2.n13 0.155672
R323 VDD2.n30 VDD2.n29 0.155672
R324 VDD2.n30 VDD2.n9 0.155672
R325 VDD2.n38 VDD2.n9 0.155672
R326 VDD2.n39 VDD2.n38 0.155672
R327 VDD2.n39 VDD2.n5 0.155672
R328 VDD2.n47 VDD2.n5 0.155672
R329 VDD2.n48 VDD2.n47 0.155672
R330 VDD2.n48 VDD2.n1 0.155672
R331 VDD2.n55 VDD2.n1 0.155672
R332 VTAIL.n240 VTAIL.n188 756.745
R333 VTAIL.n54 VTAIL.n2 756.745
R334 VTAIL.n182 VTAIL.n130 756.745
R335 VTAIL.n120 VTAIL.n68 756.745
R336 VTAIL.n207 VTAIL.n206 585
R337 VTAIL.n204 VTAIL.n203 585
R338 VTAIL.n213 VTAIL.n212 585
R339 VTAIL.n215 VTAIL.n214 585
R340 VTAIL.n200 VTAIL.n199 585
R341 VTAIL.n221 VTAIL.n220 585
R342 VTAIL.n224 VTAIL.n223 585
R343 VTAIL.n222 VTAIL.n196 585
R344 VTAIL.n229 VTAIL.n195 585
R345 VTAIL.n231 VTAIL.n230 585
R346 VTAIL.n233 VTAIL.n232 585
R347 VTAIL.n192 VTAIL.n191 585
R348 VTAIL.n239 VTAIL.n238 585
R349 VTAIL.n241 VTAIL.n240 585
R350 VTAIL.n21 VTAIL.n20 585
R351 VTAIL.n18 VTAIL.n17 585
R352 VTAIL.n27 VTAIL.n26 585
R353 VTAIL.n29 VTAIL.n28 585
R354 VTAIL.n14 VTAIL.n13 585
R355 VTAIL.n35 VTAIL.n34 585
R356 VTAIL.n38 VTAIL.n37 585
R357 VTAIL.n36 VTAIL.n10 585
R358 VTAIL.n43 VTAIL.n9 585
R359 VTAIL.n45 VTAIL.n44 585
R360 VTAIL.n47 VTAIL.n46 585
R361 VTAIL.n6 VTAIL.n5 585
R362 VTAIL.n53 VTAIL.n52 585
R363 VTAIL.n55 VTAIL.n54 585
R364 VTAIL.n183 VTAIL.n182 585
R365 VTAIL.n181 VTAIL.n180 585
R366 VTAIL.n134 VTAIL.n133 585
R367 VTAIL.n175 VTAIL.n174 585
R368 VTAIL.n173 VTAIL.n172 585
R369 VTAIL.n171 VTAIL.n137 585
R370 VTAIL.n141 VTAIL.n138 585
R371 VTAIL.n166 VTAIL.n165 585
R372 VTAIL.n164 VTAIL.n163 585
R373 VTAIL.n143 VTAIL.n142 585
R374 VTAIL.n158 VTAIL.n157 585
R375 VTAIL.n156 VTAIL.n155 585
R376 VTAIL.n147 VTAIL.n146 585
R377 VTAIL.n150 VTAIL.n149 585
R378 VTAIL.n121 VTAIL.n120 585
R379 VTAIL.n119 VTAIL.n118 585
R380 VTAIL.n72 VTAIL.n71 585
R381 VTAIL.n113 VTAIL.n112 585
R382 VTAIL.n111 VTAIL.n110 585
R383 VTAIL.n109 VTAIL.n75 585
R384 VTAIL.n79 VTAIL.n76 585
R385 VTAIL.n104 VTAIL.n103 585
R386 VTAIL.n102 VTAIL.n101 585
R387 VTAIL.n81 VTAIL.n80 585
R388 VTAIL.n96 VTAIL.n95 585
R389 VTAIL.n94 VTAIL.n93 585
R390 VTAIL.n85 VTAIL.n84 585
R391 VTAIL.n88 VTAIL.n87 585
R392 VTAIL.t7 VTAIL.n148 329.038
R393 VTAIL.t15 VTAIL.n86 329.038
R394 VTAIL.t14 VTAIL.n205 329.038
R395 VTAIL.t19 VTAIL.n19 329.038
R396 VTAIL.n206 VTAIL.n203 171.744
R397 VTAIL.n213 VTAIL.n203 171.744
R398 VTAIL.n214 VTAIL.n213 171.744
R399 VTAIL.n214 VTAIL.n199 171.744
R400 VTAIL.n221 VTAIL.n199 171.744
R401 VTAIL.n223 VTAIL.n221 171.744
R402 VTAIL.n223 VTAIL.n222 171.744
R403 VTAIL.n222 VTAIL.n195 171.744
R404 VTAIL.n231 VTAIL.n195 171.744
R405 VTAIL.n232 VTAIL.n231 171.744
R406 VTAIL.n232 VTAIL.n191 171.744
R407 VTAIL.n239 VTAIL.n191 171.744
R408 VTAIL.n240 VTAIL.n239 171.744
R409 VTAIL.n20 VTAIL.n17 171.744
R410 VTAIL.n27 VTAIL.n17 171.744
R411 VTAIL.n28 VTAIL.n27 171.744
R412 VTAIL.n28 VTAIL.n13 171.744
R413 VTAIL.n35 VTAIL.n13 171.744
R414 VTAIL.n37 VTAIL.n35 171.744
R415 VTAIL.n37 VTAIL.n36 171.744
R416 VTAIL.n36 VTAIL.n9 171.744
R417 VTAIL.n45 VTAIL.n9 171.744
R418 VTAIL.n46 VTAIL.n45 171.744
R419 VTAIL.n46 VTAIL.n5 171.744
R420 VTAIL.n53 VTAIL.n5 171.744
R421 VTAIL.n54 VTAIL.n53 171.744
R422 VTAIL.n182 VTAIL.n181 171.744
R423 VTAIL.n181 VTAIL.n133 171.744
R424 VTAIL.n174 VTAIL.n133 171.744
R425 VTAIL.n174 VTAIL.n173 171.744
R426 VTAIL.n173 VTAIL.n137 171.744
R427 VTAIL.n141 VTAIL.n137 171.744
R428 VTAIL.n165 VTAIL.n141 171.744
R429 VTAIL.n165 VTAIL.n164 171.744
R430 VTAIL.n164 VTAIL.n142 171.744
R431 VTAIL.n157 VTAIL.n142 171.744
R432 VTAIL.n157 VTAIL.n156 171.744
R433 VTAIL.n156 VTAIL.n146 171.744
R434 VTAIL.n149 VTAIL.n146 171.744
R435 VTAIL.n120 VTAIL.n119 171.744
R436 VTAIL.n119 VTAIL.n71 171.744
R437 VTAIL.n112 VTAIL.n71 171.744
R438 VTAIL.n112 VTAIL.n111 171.744
R439 VTAIL.n111 VTAIL.n75 171.744
R440 VTAIL.n79 VTAIL.n75 171.744
R441 VTAIL.n103 VTAIL.n79 171.744
R442 VTAIL.n103 VTAIL.n102 171.744
R443 VTAIL.n102 VTAIL.n80 171.744
R444 VTAIL.n95 VTAIL.n80 171.744
R445 VTAIL.n95 VTAIL.n94 171.744
R446 VTAIL.n94 VTAIL.n84 171.744
R447 VTAIL.n87 VTAIL.n84 171.744
R448 VTAIL.n206 VTAIL.t14 85.8723
R449 VTAIL.n20 VTAIL.t19 85.8723
R450 VTAIL.n149 VTAIL.t7 85.8723
R451 VTAIL.n87 VTAIL.t15 85.8723
R452 VTAIL.n129 VTAIL.n128 60.5449
R453 VTAIL.n127 VTAIL.n126 60.5449
R454 VTAIL.n67 VTAIL.n66 60.5449
R455 VTAIL.n65 VTAIL.n64 60.5449
R456 VTAIL.n247 VTAIL.n246 60.5448
R457 VTAIL.n1 VTAIL.n0 60.5448
R458 VTAIL.n61 VTAIL.n60 60.5448
R459 VTAIL.n63 VTAIL.n62 60.5448
R460 VTAIL.n245 VTAIL.n244 33.5429
R461 VTAIL.n59 VTAIL.n58 33.5429
R462 VTAIL.n187 VTAIL.n186 33.5429
R463 VTAIL.n125 VTAIL.n124 33.5429
R464 VTAIL.n65 VTAIL.n63 27.5307
R465 VTAIL.n245 VTAIL.n187 24.5824
R466 VTAIL.n230 VTAIL.n229 13.1884
R467 VTAIL.n44 VTAIL.n43 13.1884
R468 VTAIL.n172 VTAIL.n171 13.1884
R469 VTAIL.n110 VTAIL.n109 13.1884
R470 VTAIL.n228 VTAIL.n196 12.8005
R471 VTAIL.n233 VTAIL.n194 12.8005
R472 VTAIL.n42 VTAIL.n10 12.8005
R473 VTAIL.n47 VTAIL.n8 12.8005
R474 VTAIL.n175 VTAIL.n136 12.8005
R475 VTAIL.n170 VTAIL.n138 12.8005
R476 VTAIL.n113 VTAIL.n74 12.8005
R477 VTAIL.n108 VTAIL.n76 12.8005
R478 VTAIL.n225 VTAIL.n224 12.0247
R479 VTAIL.n234 VTAIL.n192 12.0247
R480 VTAIL.n39 VTAIL.n38 12.0247
R481 VTAIL.n48 VTAIL.n6 12.0247
R482 VTAIL.n176 VTAIL.n134 12.0247
R483 VTAIL.n167 VTAIL.n166 12.0247
R484 VTAIL.n114 VTAIL.n72 12.0247
R485 VTAIL.n105 VTAIL.n104 12.0247
R486 VTAIL.n220 VTAIL.n198 11.249
R487 VTAIL.n238 VTAIL.n237 11.249
R488 VTAIL.n34 VTAIL.n12 11.249
R489 VTAIL.n52 VTAIL.n51 11.249
R490 VTAIL.n180 VTAIL.n179 11.249
R491 VTAIL.n163 VTAIL.n140 11.249
R492 VTAIL.n118 VTAIL.n117 11.249
R493 VTAIL.n101 VTAIL.n78 11.249
R494 VTAIL.n207 VTAIL.n205 10.7239
R495 VTAIL.n21 VTAIL.n19 10.7239
R496 VTAIL.n150 VTAIL.n148 10.7239
R497 VTAIL.n88 VTAIL.n86 10.7239
R498 VTAIL.n219 VTAIL.n200 10.4732
R499 VTAIL.n241 VTAIL.n190 10.4732
R500 VTAIL.n33 VTAIL.n14 10.4732
R501 VTAIL.n55 VTAIL.n4 10.4732
R502 VTAIL.n183 VTAIL.n132 10.4732
R503 VTAIL.n162 VTAIL.n143 10.4732
R504 VTAIL.n121 VTAIL.n70 10.4732
R505 VTAIL.n100 VTAIL.n81 10.4732
R506 VTAIL.n216 VTAIL.n215 9.69747
R507 VTAIL.n242 VTAIL.n188 9.69747
R508 VTAIL.n30 VTAIL.n29 9.69747
R509 VTAIL.n56 VTAIL.n2 9.69747
R510 VTAIL.n184 VTAIL.n130 9.69747
R511 VTAIL.n159 VTAIL.n158 9.69747
R512 VTAIL.n122 VTAIL.n68 9.69747
R513 VTAIL.n97 VTAIL.n96 9.69747
R514 VTAIL.n244 VTAIL.n243 9.45567
R515 VTAIL.n58 VTAIL.n57 9.45567
R516 VTAIL.n186 VTAIL.n185 9.45567
R517 VTAIL.n124 VTAIL.n123 9.45567
R518 VTAIL.n243 VTAIL.n242 9.3005
R519 VTAIL.n190 VTAIL.n189 9.3005
R520 VTAIL.n237 VTAIL.n236 9.3005
R521 VTAIL.n235 VTAIL.n234 9.3005
R522 VTAIL.n194 VTAIL.n193 9.3005
R523 VTAIL.n209 VTAIL.n208 9.3005
R524 VTAIL.n211 VTAIL.n210 9.3005
R525 VTAIL.n202 VTAIL.n201 9.3005
R526 VTAIL.n217 VTAIL.n216 9.3005
R527 VTAIL.n219 VTAIL.n218 9.3005
R528 VTAIL.n198 VTAIL.n197 9.3005
R529 VTAIL.n226 VTAIL.n225 9.3005
R530 VTAIL.n228 VTAIL.n227 9.3005
R531 VTAIL.n57 VTAIL.n56 9.3005
R532 VTAIL.n4 VTAIL.n3 9.3005
R533 VTAIL.n51 VTAIL.n50 9.3005
R534 VTAIL.n49 VTAIL.n48 9.3005
R535 VTAIL.n8 VTAIL.n7 9.3005
R536 VTAIL.n23 VTAIL.n22 9.3005
R537 VTAIL.n25 VTAIL.n24 9.3005
R538 VTAIL.n16 VTAIL.n15 9.3005
R539 VTAIL.n31 VTAIL.n30 9.3005
R540 VTAIL.n33 VTAIL.n32 9.3005
R541 VTAIL.n12 VTAIL.n11 9.3005
R542 VTAIL.n40 VTAIL.n39 9.3005
R543 VTAIL.n42 VTAIL.n41 9.3005
R544 VTAIL.n152 VTAIL.n151 9.3005
R545 VTAIL.n154 VTAIL.n153 9.3005
R546 VTAIL.n145 VTAIL.n144 9.3005
R547 VTAIL.n160 VTAIL.n159 9.3005
R548 VTAIL.n162 VTAIL.n161 9.3005
R549 VTAIL.n140 VTAIL.n139 9.3005
R550 VTAIL.n168 VTAIL.n167 9.3005
R551 VTAIL.n170 VTAIL.n169 9.3005
R552 VTAIL.n185 VTAIL.n184 9.3005
R553 VTAIL.n132 VTAIL.n131 9.3005
R554 VTAIL.n179 VTAIL.n178 9.3005
R555 VTAIL.n177 VTAIL.n176 9.3005
R556 VTAIL.n136 VTAIL.n135 9.3005
R557 VTAIL.n90 VTAIL.n89 9.3005
R558 VTAIL.n92 VTAIL.n91 9.3005
R559 VTAIL.n83 VTAIL.n82 9.3005
R560 VTAIL.n98 VTAIL.n97 9.3005
R561 VTAIL.n100 VTAIL.n99 9.3005
R562 VTAIL.n78 VTAIL.n77 9.3005
R563 VTAIL.n106 VTAIL.n105 9.3005
R564 VTAIL.n108 VTAIL.n107 9.3005
R565 VTAIL.n123 VTAIL.n122 9.3005
R566 VTAIL.n70 VTAIL.n69 9.3005
R567 VTAIL.n117 VTAIL.n116 9.3005
R568 VTAIL.n115 VTAIL.n114 9.3005
R569 VTAIL.n74 VTAIL.n73 9.3005
R570 VTAIL.n212 VTAIL.n202 8.92171
R571 VTAIL.n26 VTAIL.n16 8.92171
R572 VTAIL.n155 VTAIL.n145 8.92171
R573 VTAIL.n93 VTAIL.n83 8.92171
R574 VTAIL.n211 VTAIL.n204 8.14595
R575 VTAIL.n25 VTAIL.n18 8.14595
R576 VTAIL.n154 VTAIL.n147 8.14595
R577 VTAIL.n92 VTAIL.n85 8.14595
R578 VTAIL.n208 VTAIL.n207 7.3702
R579 VTAIL.n22 VTAIL.n21 7.3702
R580 VTAIL.n151 VTAIL.n150 7.3702
R581 VTAIL.n89 VTAIL.n88 7.3702
R582 VTAIL.n208 VTAIL.n204 5.81868
R583 VTAIL.n22 VTAIL.n18 5.81868
R584 VTAIL.n151 VTAIL.n147 5.81868
R585 VTAIL.n89 VTAIL.n85 5.81868
R586 VTAIL.n212 VTAIL.n211 5.04292
R587 VTAIL.n26 VTAIL.n25 5.04292
R588 VTAIL.n155 VTAIL.n154 5.04292
R589 VTAIL.n93 VTAIL.n92 5.04292
R590 VTAIL.n215 VTAIL.n202 4.26717
R591 VTAIL.n244 VTAIL.n188 4.26717
R592 VTAIL.n29 VTAIL.n16 4.26717
R593 VTAIL.n58 VTAIL.n2 4.26717
R594 VTAIL.n186 VTAIL.n130 4.26717
R595 VTAIL.n158 VTAIL.n145 4.26717
R596 VTAIL.n124 VTAIL.n68 4.26717
R597 VTAIL.n96 VTAIL.n83 4.26717
R598 VTAIL.n216 VTAIL.n200 3.49141
R599 VTAIL.n242 VTAIL.n241 3.49141
R600 VTAIL.n30 VTAIL.n14 3.49141
R601 VTAIL.n56 VTAIL.n55 3.49141
R602 VTAIL.n184 VTAIL.n183 3.49141
R603 VTAIL.n159 VTAIL.n143 3.49141
R604 VTAIL.n122 VTAIL.n121 3.49141
R605 VTAIL.n97 VTAIL.n81 3.49141
R606 VTAIL.n246 VTAIL.t10 3.02422
R607 VTAIL.n246 VTAIL.t18 3.02422
R608 VTAIL.n0 VTAIL.t9 3.02422
R609 VTAIL.n0 VTAIL.t17 3.02422
R610 VTAIL.n60 VTAIL.t6 3.02422
R611 VTAIL.n60 VTAIL.t2 3.02422
R612 VTAIL.n62 VTAIL.t4 3.02422
R613 VTAIL.n62 VTAIL.t1 3.02422
R614 VTAIL.n128 VTAIL.t0 3.02422
R615 VTAIL.n128 VTAIL.t8 3.02422
R616 VTAIL.n126 VTAIL.t3 3.02422
R617 VTAIL.n126 VTAIL.t5 3.02422
R618 VTAIL.n66 VTAIL.t11 3.02422
R619 VTAIL.n66 VTAIL.t12 3.02422
R620 VTAIL.n64 VTAIL.t13 3.02422
R621 VTAIL.n64 VTAIL.t16 3.02422
R622 VTAIL.n67 VTAIL.n65 2.94878
R623 VTAIL.n125 VTAIL.n67 2.94878
R624 VTAIL.n129 VTAIL.n127 2.94878
R625 VTAIL.n187 VTAIL.n129 2.94878
R626 VTAIL.n63 VTAIL.n61 2.94878
R627 VTAIL.n61 VTAIL.n59 2.94878
R628 VTAIL.n247 VTAIL.n245 2.94878
R629 VTAIL.n220 VTAIL.n219 2.71565
R630 VTAIL.n238 VTAIL.n190 2.71565
R631 VTAIL.n34 VTAIL.n33 2.71565
R632 VTAIL.n52 VTAIL.n4 2.71565
R633 VTAIL.n180 VTAIL.n132 2.71565
R634 VTAIL.n163 VTAIL.n162 2.71565
R635 VTAIL.n118 VTAIL.n70 2.71565
R636 VTAIL.n101 VTAIL.n100 2.71565
R637 VTAIL.n209 VTAIL.n205 2.41282
R638 VTAIL.n23 VTAIL.n19 2.41282
R639 VTAIL.n152 VTAIL.n148 2.41282
R640 VTAIL.n90 VTAIL.n86 2.41282
R641 VTAIL VTAIL.n1 2.2699
R642 VTAIL.n127 VTAIL.n125 1.94447
R643 VTAIL.n59 VTAIL.n1 1.94447
R644 VTAIL.n224 VTAIL.n198 1.93989
R645 VTAIL.n237 VTAIL.n192 1.93989
R646 VTAIL.n38 VTAIL.n12 1.93989
R647 VTAIL.n51 VTAIL.n6 1.93989
R648 VTAIL.n179 VTAIL.n134 1.93989
R649 VTAIL.n166 VTAIL.n140 1.93989
R650 VTAIL.n117 VTAIL.n72 1.93989
R651 VTAIL.n104 VTAIL.n78 1.93989
R652 VTAIL.n225 VTAIL.n196 1.16414
R653 VTAIL.n234 VTAIL.n233 1.16414
R654 VTAIL.n39 VTAIL.n10 1.16414
R655 VTAIL.n48 VTAIL.n47 1.16414
R656 VTAIL.n176 VTAIL.n175 1.16414
R657 VTAIL.n167 VTAIL.n138 1.16414
R658 VTAIL.n114 VTAIL.n113 1.16414
R659 VTAIL.n105 VTAIL.n76 1.16414
R660 VTAIL VTAIL.n247 0.679379
R661 VTAIL.n229 VTAIL.n228 0.388379
R662 VTAIL.n230 VTAIL.n194 0.388379
R663 VTAIL.n43 VTAIL.n42 0.388379
R664 VTAIL.n44 VTAIL.n8 0.388379
R665 VTAIL.n172 VTAIL.n136 0.388379
R666 VTAIL.n171 VTAIL.n170 0.388379
R667 VTAIL.n110 VTAIL.n74 0.388379
R668 VTAIL.n109 VTAIL.n108 0.388379
R669 VTAIL.n210 VTAIL.n209 0.155672
R670 VTAIL.n210 VTAIL.n201 0.155672
R671 VTAIL.n217 VTAIL.n201 0.155672
R672 VTAIL.n218 VTAIL.n217 0.155672
R673 VTAIL.n218 VTAIL.n197 0.155672
R674 VTAIL.n226 VTAIL.n197 0.155672
R675 VTAIL.n227 VTAIL.n226 0.155672
R676 VTAIL.n227 VTAIL.n193 0.155672
R677 VTAIL.n235 VTAIL.n193 0.155672
R678 VTAIL.n236 VTAIL.n235 0.155672
R679 VTAIL.n236 VTAIL.n189 0.155672
R680 VTAIL.n243 VTAIL.n189 0.155672
R681 VTAIL.n24 VTAIL.n23 0.155672
R682 VTAIL.n24 VTAIL.n15 0.155672
R683 VTAIL.n31 VTAIL.n15 0.155672
R684 VTAIL.n32 VTAIL.n31 0.155672
R685 VTAIL.n32 VTAIL.n11 0.155672
R686 VTAIL.n40 VTAIL.n11 0.155672
R687 VTAIL.n41 VTAIL.n40 0.155672
R688 VTAIL.n41 VTAIL.n7 0.155672
R689 VTAIL.n49 VTAIL.n7 0.155672
R690 VTAIL.n50 VTAIL.n49 0.155672
R691 VTAIL.n50 VTAIL.n3 0.155672
R692 VTAIL.n57 VTAIL.n3 0.155672
R693 VTAIL.n185 VTAIL.n131 0.155672
R694 VTAIL.n178 VTAIL.n131 0.155672
R695 VTAIL.n178 VTAIL.n177 0.155672
R696 VTAIL.n177 VTAIL.n135 0.155672
R697 VTAIL.n169 VTAIL.n135 0.155672
R698 VTAIL.n169 VTAIL.n168 0.155672
R699 VTAIL.n168 VTAIL.n139 0.155672
R700 VTAIL.n161 VTAIL.n139 0.155672
R701 VTAIL.n161 VTAIL.n160 0.155672
R702 VTAIL.n160 VTAIL.n144 0.155672
R703 VTAIL.n153 VTAIL.n144 0.155672
R704 VTAIL.n153 VTAIL.n152 0.155672
R705 VTAIL.n123 VTAIL.n69 0.155672
R706 VTAIL.n116 VTAIL.n69 0.155672
R707 VTAIL.n116 VTAIL.n115 0.155672
R708 VTAIL.n115 VTAIL.n73 0.155672
R709 VTAIL.n107 VTAIL.n73 0.155672
R710 VTAIL.n107 VTAIL.n106 0.155672
R711 VTAIL.n106 VTAIL.n77 0.155672
R712 VTAIL.n99 VTAIL.n77 0.155672
R713 VTAIL.n99 VTAIL.n98 0.155672
R714 VTAIL.n98 VTAIL.n82 0.155672
R715 VTAIL.n91 VTAIL.n82 0.155672
R716 VTAIL.n91 VTAIL.n90 0.155672
R717 VP.n29 VP.n28 161.3
R718 VP.n30 VP.n25 161.3
R719 VP.n32 VP.n31 161.3
R720 VP.n33 VP.n24 161.3
R721 VP.n35 VP.n34 161.3
R722 VP.n36 VP.n23 161.3
R723 VP.n38 VP.n37 161.3
R724 VP.n39 VP.n22 161.3
R725 VP.n41 VP.n40 161.3
R726 VP.n42 VP.n21 161.3
R727 VP.n44 VP.n43 161.3
R728 VP.n45 VP.n20 161.3
R729 VP.n47 VP.n46 161.3
R730 VP.n49 VP.n48 161.3
R731 VP.n50 VP.n18 161.3
R732 VP.n52 VP.n51 161.3
R733 VP.n53 VP.n17 161.3
R734 VP.n55 VP.n54 161.3
R735 VP.n56 VP.n16 161.3
R736 VP.n58 VP.n57 161.3
R737 VP.n103 VP.n102 161.3
R738 VP.n101 VP.n1 161.3
R739 VP.n100 VP.n99 161.3
R740 VP.n98 VP.n2 161.3
R741 VP.n97 VP.n96 161.3
R742 VP.n95 VP.n3 161.3
R743 VP.n94 VP.n93 161.3
R744 VP.n92 VP.n91 161.3
R745 VP.n90 VP.n5 161.3
R746 VP.n89 VP.n88 161.3
R747 VP.n87 VP.n6 161.3
R748 VP.n86 VP.n85 161.3
R749 VP.n84 VP.n7 161.3
R750 VP.n83 VP.n82 161.3
R751 VP.n81 VP.n8 161.3
R752 VP.n80 VP.n79 161.3
R753 VP.n78 VP.n9 161.3
R754 VP.n77 VP.n76 161.3
R755 VP.n75 VP.n10 161.3
R756 VP.n74 VP.n73 161.3
R757 VP.n71 VP.n11 161.3
R758 VP.n70 VP.n69 161.3
R759 VP.n68 VP.n12 161.3
R760 VP.n67 VP.n66 161.3
R761 VP.n65 VP.n13 161.3
R762 VP.n64 VP.n63 161.3
R763 VP.n62 VP.n14 161.3
R764 VP.n26 VP.t6 117.064
R765 VP.n83 VP.t7 83.8435
R766 VP.n60 VP.t2 83.8435
R767 VP.n72 VP.t9 83.8435
R768 VP.n4 VP.t1 83.8435
R769 VP.n0 VP.t8 83.8435
R770 VP.n38 VP.t3 83.8435
R771 VP.n15 VP.t0 83.8435
R772 VP.n19 VP.t4 83.8435
R773 VP.n27 VP.t5 83.8435
R774 VP.n61 VP.n60 73.4298
R775 VP.n104 VP.n0 73.4298
R776 VP.n59 VP.n15 73.4298
R777 VP.n78 VP.n77 56.5193
R778 VP.n89 VP.n6 56.5193
R779 VP.n44 VP.n21 56.5193
R780 VP.n33 VP.n32 56.5193
R781 VP.n61 VP.n59 54.9236
R782 VP.n27 VP.n26 53.3325
R783 VP.n66 VP.n65 53.1199
R784 VP.n100 VP.n2 53.1199
R785 VP.n55 VP.n17 53.1199
R786 VP.n66 VP.n12 27.8669
R787 VP.n96 VP.n2 27.8669
R788 VP.n51 VP.n17 27.8669
R789 VP.n64 VP.n14 24.4675
R790 VP.n65 VP.n64 24.4675
R791 VP.n70 VP.n12 24.4675
R792 VP.n71 VP.n70 24.4675
R793 VP.n73 VP.n10 24.4675
R794 VP.n77 VP.n10 24.4675
R795 VP.n79 VP.n78 24.4675
R796 VP.n79 VP.n8 24.4675
R797 VP.n83 VP.n8 24.4675
R798 VP.n84 VP.n83 24.4675
R799 VP.n85 VP.n84 24.4675
R800 VP.n85 VP.n6 24.4675
R801 VP.n90 VP.n89 24.4675
R802 VP.n91 VP.n90 24.4675
R803 VP.n95 VP.n94 24.4675
R804 VP.n96 VP.n95 24.4675
R805 VP.n101 VP.n100 24.4675
R806 VP.n102 VP.n101 24.4675
R807 VP.n56 VP.n55 24.4675
R808 VP.n57 VP.n56 24.4675
R809 VP.n45 VP.n44 24.4675
R810 VP.n46 VP.n45 24.4675
R811 VP.n50 VP.n49 24.4675
R812 VP.n51 VP.n50 24.4675
R813 VP.n34 VP.n33 24.4675
R814 VP.n34 VP.n23 24.4675
R815 VP.n38 VP.n23 24.4675
R816 VP.n39 VP.n38 24.4675
R817 VP.n40 VP.n39 24.4675
R818 VP.n40 VP.n21 24.4675
R819 VP.n28 VP.n25 24.4675
R820 VP.n32 VP.n25 24.4675
R821 VP.n73 VP.n72 20.5528
R822 VP.n91 VP.n4 20.5528
R823 VP.n46 VP.n19 20.5528
R824 VP.n28 VP.n27 20.5528
R825 VP.n60 VP.n14 16.6381
R826 VP.n102 VP.n0 16.6381
R827 VP.n57 VP.n15 16.6381
R828 VP.n29 VP.n26 4.0705
R829 VP.n72 VP.n71 3.91522
R830 VP.n94 VP.n4 3.91522
R831 VP.n49 VP.n19 3.91522
R832 VP.n59 VP.n58 0.354971
R833 VP.n62 VP.n61 0.354971
R834 VP.n104 VP.n103 0.354971
R835 VP VP.n104 0.26696
R836 VP.n30 VP.n29 0.189894
R837 VP.n31 VP.n30 0.189894
R838 VP.n31 VP.n24 0.189894
R839 VP.n35 VP.n24 0.189894
R840 VP.n36 VP.n35 0.189894
R841 VP.n37 VP.n36 0.189894
R842 VP.n37 VP.n22 0.189894
R843 VP.n41 VP.n22 0.189894
R844 VP.n42 VP.n41 0.189894
R845 VP.n43 VP.n42 0.189894
R846 VP.n43 VP.n20 0.189894
R847 VP.n47 VP.n20 0.189894
R848 VP.n48 VP.n47 0.189894
R849 VP.n48 VP.n18 0.189894
R850 VP.n52 VP.n18 0.189894
R851 VP.n53 VP.n52 0.189894
R852 VP.n54 VP.n53 0.189894
R853 VP.n54 VP.n16 0.189894
R854 VP.n58 VP.n16 0.189894
R855 VP.n63 VP.n62 0.189894
R856 VP.n63 VP.n13 0.189894
R857 VP.n67 VP.n13 0.189894
R858 VP.n68 VP.n67 0.189894
R859 VP.n69 VP.n68 0.189894
R860 VP.n69 VP.n11 0.189894
R861 VP.n74 VP.n11 0.189894
R862 VP.n75 VP.n74 0.189894
R863 VP.n76 VP.n75 0.189894
R864 VP.n76 VP.n9 0.189894
R865 VP.n80 VP.n9 0.189894
R866 VP.n81 VP.n80 0.189894
R867 VP.n82 VP.n81 0.189894
R868 VP.n82 VP.n7 0.189894
R869 VP.n86 VP.n7 0.189894
R870 VP.n87 VP.n86 0.189894
R871 VP.n88 VP.n87 0.189894
R872 VP.n88 VP.n5 0.189894
R873 VP.n92 VP.n5 0.189894
R874 VP.n93 VP.n92 0.189894
R875 VP.n93 VP.n3 0.189894
R876 VP.n97 VP.n3 0.189894
R877 VP.n98 VP.n97 0.189894
R878 VP.n99 VP.n98 0.189894
R879 VP.n99 VP.n1 0.189894
R880 VP.n103 VP.n1 0.189894
R881 VDD1.n52 VDD1.n0 756.745
R882 VDD1.n111 VDD1.n59 756.745
R883 VDD1.n53 VDD1.n52 585
R884 VDD1.n51 VDD1.n50 585
R885 VDD1.n4 VDD1.n3 585
R886 VDD1.n45 VDD1.n44 585
R887 VDD1.n43 VDD1.n42 585
R888 VDD1.n41 VDD1.n7 585
R889 VDD1.n11 VDD1.n8 585
R890 VDD1.n36 VDD1.n35 585
R891 VDD1.n34 VDD1.n33 585
R892 VDD1.n13 VDD1.n12 585
R893 VDD1.n28 VDD1.n27 585
R894 VDD1.n26 VDD1.n25 585
R895 VDD1.n17 VDD1.n16 585
R896 VDD1.n20 VDD1.n19 585
R897 VDD1.n78 VDD1.n77 585
R898 VDD1.n75 VDD1.n74 585
R899 VDD1.n84 VDD1.n83 585
R900 VDD1.n86 VDD1.n85 585
R901 VDD1.n71 VDD1.n70 585
R902 VDD1.n92 VDD1.n91 585
R903 VDD1.n95 VDD1.n94 585
R904 VDD1.n93 VDD1.n67 585
R905 VDD1.n100 VDD1.n66 585
R906 VDD1.n102 VDD1.n101 585
R907 VDD1.n104 VDD1.n103 585
R908 VDD1.n63 VDD1.n62 585
R909 VDD1.n110 VDD1.n109 585
R910 VDD1.n112 VDD1.n111 585
R911 VDD1.t3 VDD1.n18 329.038
R912 VDD1.t7 VDD1.n76 329.038
R913 VDD1.n52 VDD1.n51 171.744
R914 VDD1.n51 VDD1.n3 171.744
R915 VDD1.n44 VDD1.n3 171.744
R916 VDD1.n44 VDD1.n43 171.744
R917 VDD1.n43 VDD1.n7 171.744
R918 VDD1.n11 VDD1.n7 171.744
R919 VDD1.n35 VDD1.n11 171.744
R920 VDD1.n35 VDD1.n34 171.744
R921 VDD1.n34 VDD1.n12 171.744
R922 VDD1.n27 VDD1.n12 171.744
R923 VDD1.n27 VDD1.n26 171.744
R924 VDD1.n26 VDD1.n16 171.744
R925 VDD1.n19 VDD1.n16 171.744
R926 VDD1.n77 VDD1.n74 171.744
R927 VDD1.n84 VDD1.n74 171.744
R928 VDD1.n85 VDD1.n84 171.744
R929 VDD1.n85 VDD1.n70 171.744
R930 VDD1.n92 VDD1.n70 171.744
R931 VDD1.n94 VDD1.n92 171.744
R932 VDD1.n94 VDD1.n93 171.744
R933 VDD1.n93 VDD1.n66 171.744
R934 VDD1.n102 VDD1.n66 171.744
R935 VDD1.n103 VDD1.n102 171.744
R936 VDD1.n103 VDD1.n62 171.744
R937 VDD1.n110 VDD1.n62 171.744
R938 VDD1.n111 VDD1.n110 171.744
R939 VDD1.n19 VDD1.t3 85.8723
R940 VDD1.n77 VDD1.t7 85.8723
R941 VDD1.n119 VDD1.n118 79.3794
R942 VDD1.n58 VDD1.n57 77.2237
R943 VDD1.n121 VDD1.n120 77.2235
R944 VDD1.n117 VDD1.n116 77.2235
R945 VDD1.n58 VDD1.n56 53.17
R946 VDD1.n117 VDD1.n115 53.17
R947 VDD1.n121 VDD1.n119 49.044
R948 VDD1.n42 VDD1.n41 13.1884
R949 VDD1.n101 VDD1.n100 13.1884
R950 VDD1.n45 VDD1.n6 12.8005
R951 VDD1.n40 VDD1.n8 12.8005
R952 VDD1.n99 VDD1.n67 12.8005
R953 VDD1.n104 VDD1.n65 12.8005
R954 VDD1.n46 VDD1.n4 12.0247
R955 VDD1.n37 VDD1.n36 12.0247
R956 VDD1.n96 VDD1.n95 12.0247
R957 VDD1.n105 VDD1.n63 12.0247
R958 VDD1.n50 VDD1.n49 11.249
R959 VDD1.n33 VDD1.n10 11.249
R960 VDD1.n91 VDD1.n69 11.249
R961 VDD1.n109 VDD1.n108 11.249
R962 VDD1.n20 VDD1.n18 10.7239
R963 VDD1.n78 VDD1.n76 10.7239
R964 VDD1.n53 VDD1.n2 10.4732
R965 VDD1.n32 VDD1.n13 10.4732
R966 VDD1.n90 VDD1.n71 10.4732
R967 VDD1.n112 VDD1.n61 10.4732
R968 VDD1.n54 VDD1.n0 9.69747
R969 VDD1.n29 VDD1.n28 9.69747
R970 VDD1.n87 VDD1.n86 9.69747
R971 VDD1.n113 VDD1.n59 9.69747
R972 VDD1.n56 VDD1.n55 9.45567
R973 VDD1.n115 VDD1.n114 9.45567
R974 VDD1.n22 VDD1.n21 9.3005
R975 VDD1.n24 VDD1.n23 9.3005
R976 VDD1.n15 VDD1.n14 9.3005
R977 VDD1.n30 VDD1.n29 9.3005
R978 VDD1.n32 VDD1.n31 9.3005
R979 VDD1.n10 VDD1.n9 9.3005
R980 VDD1.n38 VDD1.n37 9.3005
R981 VDD1.n40 VDD1.n39 9.3005
R982 VDD1.n55 VDD1.n54 9.3005
R983 VDD1.n2 VDD1.n1 9.3005
R984 VDD1.n49 VDD1.n48 9.3005
R985 VDD1.n47 VDD1.n46 9.3005
R986 VDD1.n6 VDD1.n5 9.3005
R987 VDD1.n114 VDD1.n113 9.3005
R988 VDD1.n61 VDD1.n60 9.3005
R989 VDD1.n108 VDD1.n107 9.3005
R990 VDD1.n106 VDD1.n105 9.3005
R991 VDD1.n65 VDD1.n64 9.3005
R992 VDD1.n80 VDD1.n79 9.3005
R993 VDD1.n82 VDD1.n81 9.3005
R994 VDD1.n73 VDD1.n72 9.3005
R995 VDD1.n88 VDD1.n87 9.3005
R996 VDD1.n90 VDD1.n89 9.3005
R997 VDD1.n69 VDD1.n68 9.3005
R998 VDD1.n97 VDD1.n96 9.3005
R999 VDD1.n99 VDD1.n98 9.3005
R1000 VDD1.n25 VDD1.n15 8.92171
R1001 VDD1.n83 VDD1.n73 8.92171
R1002 VDD1.n24 VDD1.n17 8.14595
R1003 VDD1.n82 VDD1.n75 8.14595
R1004 VDD1.n21 VDD1.n20 7.3702
R1005 VDD1.n79 VDD1.n78 7.3702
R1006 VDD1.n21 VDD1.n17 5.81868
R1007 VDD1.n79 VDD1.n75 5.81868
R1008 VDD1.n25 VDD1.n24 5.04292
R1009 VDD1.n83 VDD1.n82 5.04292
R1010 VDD1.n56 VDD1.n0 4.26717
R1011 VDD1.n28 VDD1.n15 4.26717
R1012 VDD1.n86 VDD1.n73 4.26717
R1013 VDD1.n115 VDD1.n59 4.26717
R1014 VDD1.n54 VDD1.n53 3.49141
R1015 VDD1.n29 VDD1.n13 3.49141
R1016 VDD1.n87 VDD1.n71 3.49141
R1017 VDD1.n113 VDD1.n112 3.49141
R1018 VDD1.n120 VDD1.t5 3.02422
R1019 VDD1.n120 VDD1.t9 3.02422
R1020 VDD1.n57 VDD1.t4 3.02422
R1021 VDD1.n57 VDD1.t6 3.02422
R1022 VDD1.n118 VDD1.t8 3.02422
R1023 VDD1.n118 VDD1.t1 3.02422
R1024 VDD1.n116 VDD1.t0 3.02422
R1025 VDD1.n116 VDD1.t2 3.02422
R1026 VDD1.n50 VDD1.n2 2.71565
R1027 VDD1.n33 VDD1.n32 2.71565
R1028 VDD1.n91 VDD1.n90 2.71565
R1029 VDD1.n109 VDD1.n61 2.71565
R1030 VDD1.n22 VDD1.n18 2.41282
R1031 VDD1.n80 VDD1.n76 2.41282
R1032 VDD1 VDD1.n121 2.15352
R1033 VDD1.n49 VDD1.n4 1.93989
R1034 VDD1.n36 VDD1.n10 1.93989
R1035 VDD1.n95 VDD1.n69 1.93989
R1036 VDD1.n108 VDD1.n63 1.93989
R1037 VDD1.n46 VDD1.n45 1.16414
R1038 VDD1.n37 VDD1.n8 1.16414
R1039 VDD1.n96 VDD1.n67 1.16414
R1040 VDD1.n105 VDD1.n104 1.16414
R1041 VDD1 VDD1.n58 0.795759
R1042 VDD1.n119 VDD1.n117 0.682223
R1043 VDD1.n42 VDD1.n6 0.388379
R1044 VDD1.n41 VDD1.n40 0.388379
R1045 VDD1.n100 VDD1.n99 0.388379
R1046 VDD1.n101 VDD1.n65 0.388379
R1047 VDD1.n55 VDD1.n1 0.155672
R1048 VDD1.n48 VDD1.n1 0.155672
R1049 VDD1.n48 VDD1.n47 0.155672
R1050 VDD1.n47 VDD1.n5 0.155672
R1051 VDD1.n39 VDD1.n5 0.155672
R1052 VDD1.n39 VDD1.n38 0.155672
R1053 VDD1.n38 VDD1.n9 0.155672
R1054 VDD1.n31 VDD1.n9 0.155672
R1055 VDD1.n31 VDD1.n30 0.155672
R1056 VDD1.n30 VDD1.n14 0.155672
R1057 VDD1.n23 VDD1.n14 0.155672
R1058 VDD1.n23 VDD1.n22 0.155672
R1059 VDD1.n81 VDD1.n80 0.155672
R1060 VDD1.n81 VDD1.n72 0.155672
R1061 VDD1.n88 VDD1.n72 0.155672
R1062 VDD1.n89 VDD1.n88 0.155672
R1063 VDD1.n89 VDD1.n68 0.155672
R1064 VDD1.n97 VDD1.n68 0.155672
R1065 VDD1.n98 VDD1.n97 0.155672
R1066 VDD1.n98 VDD1.n64 0.155672
R1067 VDD1.n106 VDD1.n64 0.155672
R1068 VDD1.n107 VDD1.n106 0.155672
R1069 VDD1.n107 VDD1.n60 0.155672
R1070 VDD1.n114 VDD1.n60 0.155672
R1071 B.n461 B.n460 585
R1072 B.n459 B.n152 585
R1073 B.n458 B.n457 585
R1074 B.n456 B.n153 585
R1075 B.n455 B.n454 585
R1076 B.n453 B.n154 585
R1077 B.n452 B.n451 585
R1078 B.n450 B.n155 585
R1079 B.n449 B.n448 585
R1080 B.n447 B.n156 585
R1081 B.n446 B.n445 585
R1082 B.n444 B.n157 585
R1083 B.n443 B.n442 585
R1084 B.n441 B.n158 585
R1085 B.n440 B.n439 585
R1086 B.n438 B.n159 585
R1087 B.n437 B.n436 585
R1088 B.n435 B.n160 585
R1089 B.n434 B.n433 585
R1090 B.n432 B.n161 585
R1091 B.n431 B.n430 585
R1092 B.n429 B.n162 585
R1093 B.n428 B.n427 585
R1094 B.n426 B.n163 585
R1095 B.n425 B.n424 585
R1096 B.n423 B.n164 585
R1097 B.n422 B.n421 585
R1098 B.n420 B.n165 585
R1099 B.n419 B.n418 585
R1100 B.n417 B.n166 585
R1101 B.n416 B.n415 585
R1102 B.n414 B.n167 585
R1103 B.n413 B.n412 585
R1104 B.n411 B.n168 585
R1105 B.n410 B.n409 585
R1106 B.n408 B.n169 585
R1107 B.n407 B.n406 585
R1108 B.n405 B.n170 585
R1109 B.n404 B.n403 585
R1110 B.n399 B.n171 585
R1111 B.n398 B.n397 585
R1112 B.n396 B.n172 585
R1113 B.n395 B.n394 585
R1114 B.n393 B.n173 585
R1115 B.n392 B.n391 585
R1116 B.n390 B.n174 585
R1117 B.n389 B.n388 585
R1118 B.n386 B.n175 585
R1119 B.n385 B.n384 585
R1120 B.n383 B.n178 585
R1121 B.n382 B.n381 585
R1122 B.n380 B.n179 585
R1123 B.n379 B.n378 585
R1124 B.n377 B.n180 585
R1125 B.n376 B.n375 585
R1126 B.n374 B.n181 585
R1127 B.n373 B.n372 585
R1128 B.n371 B.n182 585
R1129 B.n370 B.n369 585
R1130 B.n368 B.n183 585
R1131 B.n367 B.n366 585
R1132 B.n365 B.n184 585
R1133 B.n364 B.n363 585
R1134 B.n362 B.n185 585
R1135 B.n361 B.n360 585
R1136 B.n359 B.n186 585
R1137 B.n358 B.n357 585
R1138 B.n356 B.n187 585
R1139 B.n355 B.n354 585
R1140 B.n353 B.n188 585
R1141 B.n352 B.n351 585
R1142 B.n350 B.n189 585
R1143 B.n349 B.n348 585
R1144 B.n347 B.n190 585
R1145 B.n346 B.n345 585
R1146 B.n344 B.n191 585
R1147 B.n343 B.n342 585
R1148 B.n341 B.n192 585
R1149 B.n340 B.n339 585
R1150 B.n338 B.n193 585
R1151 B.n337 B.n336 585
R1152 B.n335 B.n194 585
R1153 B.n334 B.n333 585
R1154 B.n332 B.n195 585
R1155 B.n331 B.n330 585
R1156 B.n462 B.n151 585
R1157 B.n464 B.n463 585
R1158 B.n465 B.n150 585
R1159 B.n467 B.n466 585
R1160 B.n468 B.n149 585
R1161 B.n470 B.n469 585
R1162 B.n471 B.n148 585
R1163 B.n473 B.n472 585
R1164 B.n474 B.n147 585
R1165 B.n476 B.n475 585
R1166 B.n477 B.n146 585
R1167 B.n479 B.n478 585
R1168 B.n480 B.n145 585
R1169 B.n482 B.n481 585
R1170 B.n483 B.n144 585
R1171 B.n485 B.n484 585
R1172 B.n486 B.n143 585
R1173 B.n488 B.n487 585
R1174 B.n489 B.n142 585
R1175 B.n491 B.n490 585
R1176 B.n492 B.n141 585
R1177 B.n494 B.n493 585
R1178 B.n495 B.n140 585
R1179 B.n497 B.n496 585
R1180 B.n498 B.n139 585
R1181 B.n500 B.n499 585
R1182 B.n501 B.n138 585
R1183 B.n503 B.n502 585
R1184 B.n504 B.n137 585
R1185 B.n506 B.n505 585
R1186 B.n507 B.n136 585
R1187 B.n509 B.n508 585
R1188 B.n510 B.n135 585
R1189 B.n512 B.n511 585
R1190 B.n513 B.n134 585
R1191 B.n515 B.n514 585
R1192 B.n516 B.n133 585
R1193 B.n518 B.n517 585
R1194 B.n519 B.n132 585
R1195 B.n521 B.n520 585
R1196 B.n522 B.n131 585
R1197 B.n524 B.n523 585
R1198 B.n525 B.n130 585
R1199 B.n527 B.n526 585
R1200 B.n528 B.n129 585
R1201 B.n530 B.n529 585
R1202 B.n531 B.n128 585
R1203 B.n533 B.n532 585
R1204 B.n534 B.n127 585
R1205 B.n536 B.n535 585
R1206 B.n537 B.n126 585
R1207 B.n539 B.n538 585
R1208 B.n540 B.n125 585
R1209 B.n542 B.n541 585
R1210 B.n543 B.n124 585
R1211 B.n545 B.n544 585
R1212 B.n546 B.n123 585
R1213 B.n548 B.n547 585
R1214 B.n549 B.n122 585
R1215 B.n551 B.n550 585
R1216 B.n552 B.n121 585
R1217 B.n554 B.n553 585
R1218 B.n555 B.n120 585
R1219 B.n557 B.n556 585
R1220 B.n558 B.n119 585
R1221 B.n560 B.n559 585
R1222 B.n561 B.n118 585
R1223 B.n563 B.n562 585
R1224 B.n564 B.n117 585
R1225 B.n566 B.n565 585
R1226 B.n567 B.n116 585
R1227 B.n569 B.n568 585
R1228 B.n570 B.n115 585
R1229 B.n572 B.n571 585
R1230 B.n573 B.n114 585
R1231 B.n575 B.n574 585
R1232 B.n576 B.n113 585
R1233 B.n578 B.n577 585
R1234 B.n579 B.n112 585
R1235 B.n581 B.n580 585
R1236 B.n582 B.n111 585
R1237 B.n584 B.n583 585
R1238 B.n585 B.n110 585
R1239 B.n587 B.n586 585
R1240 B.n588 B.n109 585
R1241 B.n590 B.n589 585
R1242 B.n591 B.n108 585
R1243 B.n593 B.n592 585
R1244 B.n594 B.n107 585
R1245 B.n596 B.n595 585
R1246 B.n597 B.n106 585
R1247 B.n599 B.n598 585
R1248 B.n600 B.n105 585
R1249 B.n602 B.n601 585
R1250 B.n603 B.n104 585
R1251 B.n605 B.n604 585
R1252 B.n606 B.n103 585
R1253 B.n608 B.n607 585
R1254 B.n609 B.n102 585
R1255 B.n611 B.n610 585
R1256 B.n612 B.n101 585
R1257 B.n614 B.n613 585
R1258 B.n615 B.n100 585
R1259 B.n617 B.n616 585
R1260 B.n618 B.n99 585
R1261 B.n620 B.n619 585
R1262 B.n621 B.n98 585
R1263 B.n623 B.n622 585
R1264 B.n624 B.n97 585
R1265 B.n626 B.n625 585
R1266 B.n627 B.n96 585
R1267 B.n629 B.n628 585
R1268 B.n630 B.n95 585
R1269 B.n632 B.n631 585
R1270 B.n633 B.n94 585
R1271 B.n635 B.n634 585
R1272 B.n636 B.n93 585
R1273 B.n638 B.n637 585
R1274 B.n639 B.n92 585
R1275 B.n641 B.n640 585
R1276 B.n642 B.n91 585
R1277 B.n644 B.n643 585
R1278 B.n645 B.n90 585
R1279 B.n647 B.n646 585
R1280 B.n648 B.n89 585
R1281 B.n650 B.n649 585
R1282 B.n651 B.n88 585
R1283 B.n653 B.n652 585
R1284 B.n654 B.n87 585
R1285 B.n656 B.n655 585
R1286 B.n657 B.n86 585
R1287 B.n659 B.n658 585
R1288 B.n660 B.n85 585
R1289 B.n662 B.n661 585
R1290 B.n663 B.n84 585
R1291 B.n665 B.n664 585
R1292 B.n666 B.n83 585
R1293 B.n668 B.n667 585
R1294 B.n797 B.n36 585
R1295 B.n796 B.n795 585
R1296 B.n794 B.n37 585
R1297 B.n793 B.n792 585
R1298 B.n791 B.n38 585
R1299 B.n790 B.n789 585
R1300 B.n788 B.n39 585
R1301 B.n787 B.n786 585
R1302 B.n785 B.n40 585
R1303 B.n784 B.n783 585
R1304 B.n782 B.n41 585
R1305 B.n781 B.n780 585
R1306 B.n779 B.n42 585
R1307 B.n778 B.n777 585
R1308 B.n776 B.n43 585
R1309 B.n775 B.n774 585
R1310 B.n773 B.n44 585
R1311 B.n772 B.n771 585
R1312 B.n770 B.n45 585
R1313 B.n769 B.n768 585
R1314 B.n767 B.n46 585
R1315 B.n766 B.n765 585
R1316 B.n764 B.n47 585
R1317 B.n763 B.n762 585
R1318 B.n761 B.n48 585
R1319 B.n760 B.n759 585
R1320 B.n758 B.n49 585
R1321 B.n757 B.n756 585
R1322 B.n755 B.n50 585
R1323 B.n754 B.n753 585
R1324 B.n752 B.n51 585
R1325 B.n751 B.n750 585
R1326 B.n749 B.n52 585
R1327 B.n748 B.n747 585
R1328 B.n746 B.n53 585
R1329 B.n745 B.n744 585
R1330 B.n743 B.n54 585
R1331 B.n742 B.n741 585
R1332 B.n739 B.n55 585
R1333 B.n738 B.n737 585
R1334 B.n736 B.n58 585
R1335 B.n735 B.n734 585
R1336 B.n733 B.n59 585
R1337 B.n732 B.n731 585
R1338 B.n730 B.n60 585
R1339 B.n729 B.n728 585
R1340 B.n727 B.n61 585
R1341 B.n725 B.n724 585
R1342 B.n723 B.n64 585
R1343 B.n722 B.n721 585
R1344 B.n720 B.n65 585
R1345 B.n719 B.n718 585
R1346 B.n717 B.n66 585
R1347 B.n716 B.n715 585
R1348 B.n714 B.n67 585
R1349 B.n713 B.n712 585
R1350 B.n711 B.n68 585
R1351 B.n710 B.n709 585
R1352 B.n708 B.n69 585
R1353 B.n707 B.n706 585
R1354 B.n705 B.n70 585
R1355 B.n704 B.n703 585
R1356 B.n702 B.n71 585
R1357 B.n701 B.n700 585
R1358 B.n699 B.n72 585
R1359 B.n698 B.n697 585
R1360 B.n696 B.n73 585
R1361 B.n695 B.n694 585
R1362 B.n693 B.n74 585
R1363 B.n692 B.n691 585
R1364 B.n690 B.n75 585
R1365 B.n689 B.n688 585
R1366 B.n687 B.n76 585
R1367 B.n686 B.n685 585
R1368 B.n684 B.n77 585
R1369 B.n683 B.n682 585
R1370 B.n681 B.n78 585
R1371 B.n680 B.n679 585
R1372 B.n678 B.n79 585
R1373 B.n677 B.n676 585
R1374 B.n675 B.n80 585
R1375 B.n674 B.n673 585
R1376 B.n672 B.n81 585
R1377 B.n671 B.n670 585
R1378 B.n669 B.n82 585
R1379 B.n799 B.n798 585
R1380 B.n800 B.n35 585
R1381 B.n802 B.n801 585
R1382 B.n803 B.n34 585
R1383 B.n805 B.n804 585
R1384 B.n806 B.n33 585
R1385 B.n808 B.n807 585
R1386 B.n809 B.n32 585
R1387 B.n811 B.n810 585
R1388 B.n812 B.n31 585
R1389 B.n814 B.n813 585
R1390 B.n815 B.n30 585
R1391 B.n817 B.n816 585
R1392 B.n818 B.n29 585
R1393 B.n820 B.n819 585
R1394 B.n821 B.n28 585
R1395 B.n823 B.n822 585
R1396 B.n824 B.n27 585
R1397 B.n826 B.n825 585
R1398 B.n827 B.n26 585
R1399 B.n829 B.n828 585
R1400 B.n830 B.n25 585
R1401 B.n832 B.n831 585
R1402 B.n833 B.n24 585
R1403 B.n835 B.n834 585
R1404 B.n836 B.n23 585
R1405 B.n838 B.n837 585
R1406 B.n839 B.n22 585
R1407 B.n841 B.n840 585
R1408 B.n842 B.n21 585
R1409 B.n844 B.n843 585
R1410 B.n845 B.n20 585
R1411 B.n847 B.n846 585
R1412 B.n848 B.n19 585
R1413 B.n850 B.n849 585
R1414 B.n851 B.n18 585
R1415 B.n853 B.n852 585
R1416 B.n854 B.n17 585
R1417 B.n856 B.n855 585
R1418 B.n857 B.n16 585
R1419 B.n859 B.n858 585
R1420 B.n860 B.n15 585
R1421 B.n862 B.n861 585
R1422 B.n863 B.n14 585
R1423 B.n865 B.n864 585
R1424 B.n866 B.n13 585
R1425 B.n868 B.n867 585
R1426 B.n869 B.n12 585
R1427 B.n871 B.n870 585
R1428 B.n872 B.n11 585
R1429 B.n874 B.n873 585
R1430 B.n875 B.n10 585
R1431 B.n877 B.n876 585
R1432 B.n878 B.n9 585
R1433 B.n880 B.n879 585
R1434 B.n881 B.n8 585
R1435 B.n883 B.n882 585
R1436 B.n884 B.n7 585
R1437 B.n886 B.n885 585
R1438 B.n887 B.n6 585
R1439 B.n889 B.n888 585
R1440 B.n890 B.n5 585
R1441 B.n892 B.n891 585
R1442 B.n893 B.n4 585
R1443 B.n895 B.n894 585
R1444 B.n896 B.n3 585
R1445 B.n898 B.n897 585
R1446 B.n899 B.n0 585
R1447 B.n2 B.n1 585
R1448 B.n230 B.n229 585
R1449 B.n232 B.n231 585
R1450 B.n233 B.n228 585
R1451 B.n235 B.n234 585
R1452 B.n236 B.n227 585
R1453 B.n238 B.n237 585
R1454 B.n239 B.n226 585
R1455 B.n241 B.n240 585
R1456 B.n242 B.n225 585
R1457 B.n244 B.n243 585
R1458 B.n245 B.n224 585
R1459 B.n247 B.n246 585
R1460 B.n248 B.n223 585
R1461 B.n250 B.n249 585
R1462 B.n251 B.n222 585
R1463 B.n253 B.n252 585
R1464 B.n254 B.n221 585
R1465 B.n256 B.n255 585
R1466 B.n257 B.n220 585
R1467 B.n259 B.n258 585
R1468 B.n260 B.n219 585
R1469 B.n262 B.n261 585
R1470 B.n263 B.n218 585
R1471 B.n265 B.n264 585
R1472 B.n266 B.n217 585
R1473 B.n268 B.n267 585
R1474 B.n269 B.n216 585
R1475 B.n271 B.n270 585
R1476 B.n272 B.n215 585
R1477 B.n274 B.n273 585
R1478 B.n275 B.n214 585
R1479 B.n277 B.n276 585
R1480 B.n278 B.n213 585
R1481 B.n280 B.n279 585
R1482 B.n281 B.n212 585
R1483 B.n283 B.n282 585
R1484 B.n284 B.n211 585
R1485 B.n286 B.n285 585
R1486 B.n287 B.n210 585
R1487 B.n289 B.n288 585
R1488 B.n290 B.n209 585
R1489 B.n292 B.n291 585
R1490 B.n293 B.n208 585
R1491 B.n295 B.n294 585
R1492 B.n296 B.n207 585
R1493 B.n298 B.n297 585
R1494 B.n299 B.n206 585
R1495 B.n301 B.n300 585
R1496 B.n302 B.n205 585
R1497 B.n304 B.n303 585
R1498 B.n305 B.n204 585
R1499 B.n307 B.n306 585
R1500 B.n308 B.n203 585
R1501 B.n310 B.n309 585
R1502 B.n311 B.n202 585
R1503 B.n313 B.n312 585
R1504 B.n314 B.n201 585
R1505 B.n316 B.n315 585
R1506 B.n317 B.n200 585
R1507 B.n319 B.n318 585
R1508 B.n320 B.n199 585
R1509 B.n322 B.n321 585
R1510 B.n323 B.n198 585
R1511 B.n325 B.n324 585
R1512 B.n326 B.n197 585
R1513 B.n328 B.n327 585
R1514 B.n329 B.n196 585
R1515 B.n330 B.n329 530.939
R1516 B.n460 B.n151 530.939
R1517 B.n669 B.n668 530.939
R1518 B.n798 B.n797 530.939
R1519 B.n400 B.t1 419.502
R1520 B.n62 B.t8 419.502
R1521 B.n176 B.t10 419.502
R1522 B.n56 B.t5 419.502
R1523 B.n401 B.t2 353.175
R1524 B.n63 B.t7 353.175
R1525 B.n177 B.t11 353.173
R1526 B.n57 B.t4 353.173
R1527 B.n176 B.t9 292.526
R1528 B.n400 B.t0 292.526
R1529 B.n62 B.t6 292.526
R1530 B.n56 B.t3 292.526
R1531 B.n901 B.n900 256.663
R1532 B.n900 B.n899 235.042
R1533 B.n900 B.n2 235.042
R1534 B.n330 B.n195 163.367
R1535 B.n334 B.n195 163.367
R1536 B.n335 B.n334 163.367
R1537 B.n336 B.n335 163.367
R1538 B.n336 B.n193 163.367
R1539 B.n340 B.n193 163.367
R1540 B.n341 B.n340 163.367
R1541 B.n342 B.n341 163.367
R1542 B.n342 B.n191 163.367
R1543 B.n346 B.n191 163.367
R1544 B.n347 B.n346 163.367
R1545 B.n348 B.n347 163.367
R1546 B.n348 B.n189 163.367
R1547 B.n352 B.n189 163.367
R1548 B.n353 B.n352 163.367
R1549 B.n354 B.n353 163.367
R1550 B.n354 B.n187 163.367
R1551 B.n358 B.n187 163.367
R1552 B.n359 B.n358 163.367
R1553 B.n360 B.n359 163.367
R1554 B.n360 B.n185 163.367
R1555 B.n364 B.n185 163.367
R1556 B.n365 B.n364 163.367
R1557 B.n366 B.n365 163.367
R1558 B.n366 B.n183 163.367
R1559 B.n370 B.n183 163.367
R1560 B.n371 B.n370 163.367
R1561 B.n372 B.n371 163.367
R1562 B.n372 B.n181 163.367
R1563 B.n376 B.n181 163.367
R1564 B.n377 B.n376 163.367
R1565 B.n378 B.n377 163.367
R1566 B.n378 B.n179 163.367
R1567 B.n382 B.n179 163.367
R1568 B.n383 B.n382 163.367
R1569 B.n384 B.n383 163.367
R1570 B.n384 B.n175 163.367
R1571 B.n389 B.n175 163.367
R1572 B.n390 B.n389 163.367
R1573 B.n391 B.n390 163.367
R1574 B.n391 B.n173 163.367
R1575 B.n395 B.n173 163.367
R1576 B.n396 B.n395 163.367
R1577 B.n397 B.n396 163.367
R1578 B.n397 B.n171 163.367
R1579 B.n404 B.n171 163.367
R1580 B.n405 B.n404 163.367
R1581 B.n406 B.n405 163.367
R1582 B.n406 B.n169 163.367
R1583 B.n410 B.n169 163.367
R1584 B.n411 B.n410 163.367
R1585 B.n412 B.n411 163.367
R1586 B.n412 B.n167 163.367
R1587 B.n416 B.n167 163.367
R1588 B.n417 B.n416 163.367
R1589 B.n418 B.n417 163.367
R1590 B.n418 B.n165 163.367
R1591 B.n422 B.n165 163.367
R1592 B.n423 B.n422 163.367
R1593 B.n424 B.n423 163.367
R1594 B.n424 B.n163 163.367
R1595 B.n428 B.n163 163.367
R1596 B.n429 B.n428 163.367
R1597 B.n430 B.n429 163.367
R1598 B.n430 B.n161 163.367
R1599 B.n434 B.n161 163.367
R1600 B.n435 B.n434 163.367
R1601 B.n436 B.n435 163.367
R1602 B.n436 B.n159 163.367
R1603 B.n440 B.n159 163.367
R1604 B.n441 B.n440 163.367
R1605 B.n442 B.n441 163.367
R1606 B.n442 B.n157 163.367
R1607 B.n446 B.n157 163.367
R1608 B.n447 B.n446 163.367
R1609 B.n448 B.n447 163.367
R1610 B.n448 B.n155 163.367
R1611 B.n452 B.n155 163.367
R1612 B.n453 B.n452 163.367
R1613 B.n454 B.n453 163.367
R1614 B.n454 B.n153 163.367
R1615 B.n458 B.n153 163.367
R1616 B.n459 B.n458 163.367
R1617 B.n460 B.n459 163.367
R1618 B.n668 B.n83 163.367
R1619 B.n664 B.n83 163.367
R1620 B.n664 B.n663 163.367
R1621 B.n663 B.n662 163.367
R1622 B.n662 B.n85 163.367
R1623 B.n658 B.n85 163.367
R1624 B.n658 B.n657 163.367
R1625 B.n657 B.n656 163.367
R1626 B.n656 B.n87 163.367
R1627 B.n652 B.n87 163.367
R1628 B.n652 B.n651 163.367
R1629 B.n651 B.n650 163.367
R1630 B.n650 B.n89 163.367
R1631 B.n646 B.n89 163.367
R1632 B.n646 B.n645 163.367
R1633 B.n645 B.n644 163.367
R1634 B.n644 B.n91 163.367
R1635 B.n640 B.n91 163.367
R1636 B.n640 B.n639 163.367
R1637 B.n639 B.n638 163.367
R1638 B.n638 B.n93 163.367
R1639 B.n634 B.n93 163.367
R1640 B.n634 B.n633 163.367
R1641 B.n633 B.n632 163.367
R1642 B.n632 B.n95 163.367
R1643 B.n628 B.n95 163.367
R1644 B.n628 B.n627 163.367
R1645 B.n627 B.n626 163.367
R1646 B.n626 B.n97 163.367
R1647 B.n622 B.n97 163.367
R1648 B.n622 B.n621 163.367
R1649 B.n621 B.n620 163.367
R1650 B.n620 B.n99 163.367
R1651 B.n616 B.n99 163.367
R1652 B.n616 B.n615 163.367
R1653 B.n615 B.n614 163.367
R1654 B.n614 B.n101 163.367
R1655 B.n610 B.n101 163.367
R1656 B.n610 B.n609 163.367
R1657 B.n609 B.n608 163.367
R1658 B.n608 B.n103 163.367
R1659 B.n604 B.n103 163.367
R1660 B.n604 B.n603 163.367
R1661 B.n603 B.n602 163.367
R1662 B.n602 B.n105 163.367
R1663 B.n598 B.n105 163.367
R1664 B.n598 B.n597 163.367
R1665 B.n597 B.n596 163.367
R1666 B.n596 B.n107 163.367
R1667 B.n592 B.n107 163.367
R1668 B.n592 B.n591 163.367
R1669 B.n591 B.n590 163.367
R1670 B.n590 B.n109 163.367
R1671 B.n586 B.n109 163.367
R1672 B.n586 B.n585 163.367
R1673 B.n585 B.n584 163.367
R1674 B.n584 B.n111 163.367
R1675 B.n580 B.n111 163.367
R1676 B.n580 B.n579 163.367
R1677 B.n579 B.n578 163.367
R1678 B.n578 B.n113 163.367
R1679 B.n574 B.n113 163.367
R1680 B.n574 B.n573 163.367
R1681 B.n573 B.n572 163.367
R1682 B.n572 B.n115 163.367
R1683 B.n568 B.n115 163.367
R1684 B.n568 B.n567 163.367
R1685 B.n567 B.n566 163.367
R1686 B.n566 B.n117 163.367
R1687 B.n562 B.n117 163.367
R1688 B.n562 B.n561 163.367
R1689 B.n561 B.n560 163.367
R1690 B.n560 B.n119 163.367
R1691 B.n556 B.n119 163.367
R1692 B.n556 B.n555 163.367
R1693 B.n555 B.n554 163.367
R1694 B.n554 B.n121 163.367
R1695 B.n550 B.n121 163.367
R1696 B.n550 B.n549 163.367
R1697 B.n549 B.n548 163.367
R1698 B.n548 B.n123 163.367
R1699 B.n544 B.n123 163.367
R1700 B.n544 B.n543 163.367
R1701 B.n543 B.n542 163.367
R1702 B.n542 B.n125 163.367
R1703 B.n538 B.n125 163.367
R1704 B.n538 B.n537 163.367
R1705 B.n537 B.n536 163.367
R1706 B.n536 B.n127 163.367
R1707 B.n532 B.n127 163.367
R1708 B.n532 B.n531 163.367
R1709 B.n531 B.n530 163.367
R1710 B.n530 B.n129 163.367
R1711 B.n526 B.n129 163.367
R1712 B.n526 B.n525 163.367
R1713 B.n525 B.n524 163.367
R1714 B.n524 B.n131 163.367
R1715 B.n520 B.n131 163.367
R1716 B.n520 B.n519 163.367
R1717 B.n519 B.n518 163.367
R1718 B.n518 B.n133 163.367
R1719 B.n514 B.n133 163.367
R1720 B.n514 B.n513 163.367
R1721 B.n513 B.n512 163.367
R1722 B.n512 B.n135 163.367
R1723 B.n508 B.n135 163.367
R1724 B.n508 B.n507 163.367
R1725 B.n507 B.n506 163.367
R1726 B.n506 B.n137 163.367
R1727 B.n502 B.n137 163.367
R1728 B.n502 B.n501 163.367
R1729 B.n501 B.n500 163.367
R1730 B.n500 B.n139 163.367
R1731 B.n496 B.n139 163.367
R1732 B.n496 B.n495 163.367
R1733 B.n495 B.n494 163.367
R1734 B.n494 B.n141 163.367
R1735 B.n490 B.n141 163.367
R1736 B.n490 B.n489 163.367
R1737 B.n489 B.n488 163.367
R1738 B.n488 B.n143 163.367
R1739 B.n484 B.n143 163.367
R1740 B.n484 B.n483 163.367
R1741 B.n483 B.n482 163.367
R1742 B.n482 B.n145 163.367
R1743 B.n478 B.n145 163.367
R1744 B.n478 B.n477 163.367
R1745 B.n477 B.n476 163.367
R1746 B.n476 B.n147 163.367
R1747 B.n472 B.n147 163.367
R1748 B.n472 B.n471 163.367
R1749 B.n471 B.n470 163.367
R1750 B.n470 B.n149 163.367
R1751 B.n466 B.n149 163.367
R1752 B.n466 B.n465 163.367
R1753 B.n465 B.n464 163.367
R1754 B.n464 B.n151 163.367
R1755 B.n797 B.n796 163.367
R1756 B.n796 B.n37 163.367
R1757 B.n792 B.n37 163.367
R1758 B.n792 B.n791 163.367
R1759 B.n791 B.n790 163.367
R1760 B.n790 B.n39 163.367
R1761 B.n786 B.n39 163.367
R1762 B.n786 B.n785 163.367
R1763 B.n785 B.n784 163.367
R1764 B.n784 B.n41 163.367
R1765 B.n780 B.n41 163.367
R1766 B.n780 B.n779 163.367
R1767 B.n779 B.n778 163.367
R1768 B.n778 B.n43 163.367
R1769 B.n774 B.n43 163.367
R1770 B.n774 B.n773 163.367
R1771 B.n773 B.n772 163.367
R1772 B.n772 B.n45 163.367
R1773 B.n768 B.n45 163.367
R1774 B.n768 B.n767 163.367
R1775 B.n767 B.n766 163.367
R1776 B.n766 B.n47 163.367
R1777 B.n762 B.n47 163.367
R1778 B.n762 B.n761 163.367
R1779 B.n761 B.n760 163.367
R1780 B.n760 B.n49 163.367
R1781 B.n756 B.n49 163.367
R1782 B.n756 B.n755 163.367
R1783 B.n755 B.n754 163.367
R1784 B.n754 B.n51 163.367
R1785 B.n750 B.n51 163.367
R1786 B.n750 B.n749 163.367
R1787 B.n749 B.n748 163.367
R1788 B.n748 B.n53 163.367
R1789 B.n744 B.n53 163.367
R1790 B.n744 B.n743 163.367
R1791 B.n743 B.n742 163.367
R1792 B.n742 B.n55 163.367
R1793 B.n737 B.n55 163.367
R1794 B.n737 B.n736 163.367
R1795 B.n736 B.n735 163.367
R1796 B.n735 B.n59 163.367
R1797 B.n731 B.n59 163.367
R1798 B.n731 B.n730 163.367
R1799 B.n730 B.n729 163.367
R1800 B.n729 B.n61 163.367
R1801 B.n724 B.n61 163.367
R1802 B.n724 B.n723 163.367
R1803 B.n723 B.n722 163.367
R1804 B.n722 B.n65 163.367
R1805 B.n718 B.n65 163.367
R1806 B.n718 B.n717 163.367
R1807 B.n717 B.n716 163.367
R1808 B.n716 B.n67 163.367
R1809 B.n712 B.n67 163.367
R1810 B.n712 B.n711 163.367
R1811 B.n711 B.n710 163.367
R1812 B.n710 B.n69 163.367
R1813 B.n706 B.n69 163.367
R1814 B.n706 B.n705 163.367
R1815 B.n705 B.n704 163.367
R1816 B.n704 B.n71 163.367
R1817 B.n700 B.n71 163.367
R1818 B.n700 B.n699 163.367
R1819 B.n699 B.n698 163.367
R1820 B.n698 B.n73 163.367
R1821 B.n694 B.n73 163.367
R1822 B.n694 B.n693 163.367
R1823 B.n693 B.n692 163.367
R1824 B.n692 B.n75 163.367
R1825 B.n688 B.n75 163.367
R1826 B.n688 B.n687 163.367
R1827 B.n687 B.n686 163.367
R1828 B.n686 B.n77 163.367
R1829 B.n682 B.n77 163.367
R1830 B.n682 B.n681 163.367
R1831 B.n681 B.n680 163.367
R1832 B.n680 B.n79 163.367
R1833 B.n676 B.n79 163.367
R1834 B.n676 B.n675 163.367
R1835 B.n675 B.n674 163.367
R1836 B.n674 B.n81 163.367
R1837 B.n670 B.n81 163.367
R1838 B.n670 B.n669 163.367
R1839 B.n798 B.n35 163.367
R1840 B.n802 B.n35 163.367
R1841 B.n803 B.n802 163.367
R1842 B.n804 B.n803 163.367
R1843 B.n804 B.n33 163.367
R1844 B.n808 B.n33 163.367
R1845 B.n809 B.n808 163.367
R1846 B.n810 B.n809 163.367
R1847 B.n810 B.n31 163.367
R1848 B.n814 B.n31 163.367
R1849 B.n815 B.n814 163.367
R1850 B.n816 B.n815 163.367
R1851 B.n816 B.n29 163.367
R1852 B.n820 B.n29 163.367
R1853 B.n821 B.n820 163.367
R1854 B.n822 B.n821 163.367
R1855 B.n822 B.n27 163.367
R1856 B.n826 B.n27 163.367
R1857 B.n827 B.n826 163.367
R1858 B.n828 B.n827 163.367
R1859 B.n828 B.n25 163.367
R1860 B.n832 B.n25 163.367
R1861 B.n833 B.n832 163.367
R1862 B.n834 B.n833 163.367
R1863 B.n834 B.n23 163.367
R1864 B.n838 B.n23 163.367
R1865 B.n839 B.n838 163.367
R1866 B.n840 B.n839 163.367
R1867 B.n840 B.n21 163.367
R1868 B.n844 B.n21 163.367
R1869 B.n845 B.n844 163.367
R1870 B.n846 B.n845 163.367
R1871 B.n846 B.n19 163.367
R1872 B.n850 B.n19 163.367
R1873 B.n851 B.n850 163.367
R1874 B.n852 B.n851 163.367
R1875 B.n852 B.n17 163.367
R1876 B.n856 B.n17 163.367
R1877 B.n857 B.n856 163.367
R1878 B.n858 B.n857 163.367
R1879 B.n858 B.n15 163.367
R1880 B.n862 B.n15 163.367
R1881 B.n863 B.n862 163.367
R1882 B.n864 B.n863 163.367
R1883 B.n864 B.n13 163.367
R1884 B.n868 B.n13 163.367
R1885 B.n869 B.n868 163.367
R1886 B.n870 B.n869 163.367
R1887 B.n870 B.n11 163.367
R1888 B.n874 B.n11 163.367
R1889 B.n875 B.n874 163.367
R1890 B.n876 B.n875 163.367
R1891 B.n876 B.n9 163.367
R1892 B.n880 B.n9 163.367
R1893 B.n881 B.n880 163.367
R1894 B.n882 B.n881 163.367
R1895 B.n882 B.n7 163.367
R1896 B.n886 B.n7 163.367
R1897 B.n887 B.n886 163.367
R1898 B.n888 B.n887 163.367
R1899 B.n888 B.n5 163.367
R1900 B.n892 B.n5 163.367
R1901 B.n893 B.n892 163.367
R1902 B.n894 B.n893 163.367
R1903 B.n894 B.n3 163.367
R1904 B.n898 B.n3 163.367
R1905 B.n899 B.n898 163.367
R1906 B.n229 B.n2 163.367
R1907 B.n232 B.n229 163.367
R1908 B.n233 B.n232 163.367
R1909 B.n234 B.n233 163.367
R1910 B.n234 B.n227 163.367
R1911 B.n238 B.n227 163.367
R1912 B.n239 B.n238 163.367
R1913 B.n240 B.n239 163.367
R1914 B.n240 B.n225 163.367
R1915 B.n244 B.n225 163.367
R1916 B.n245 B.n244 163.367
R1917 B.n246 B.n245 163.367
R1918 B.n246 B.n223 163.367
R1919 B.n250 B.n223 163.367
R1920 B.n251 B.n250 163.367
R1921 B.n252 B.n251 163.367
R1922 B.n252 B.n221 163.367
R1923 B.n256 B.n221 163.367
R1924 B.n257 B.n256 163.367
R1925 B.n258 B.n257 163.367
R1926 B.n258 B.n219 163.367
R1927 B.n262 B.n219 163.367
R1928 B.n263 B.n262 163.367
R1929 B.n264 B.n263 163.367
R1930 B.n264 B.n217 163.367
R1931 B.n268 B.n217 163.367
R1932 B.n269 B.n268 163.367
R1933 B.n270 B.n269 163.367
R1934 B.n270 B.n215 163.367
R1935 B.n274 B.n215 163.367
R1936 B.n275 B.n274 163.367
R1937 B.n276 B.n275 163.367
R1938 B.n276 B.n213 163.367
R1939 B.n280 B.n213 163.367
R1940 B.n281 B.n280 163.367
R1941 B.n282 B.n281 163.367
R1942 B.n282 B.n211 163.367
R1943 B.n286 B.n211 163.367
R1944 B.n287 B.n286 163.367
R1945 B.n288 B.n287 163.367
R1946 B.n288 B.n209 163.367
R1947 B.n292 B.n209 163.367
R1948 B.n293 B.n292 163.367
R1949 B.n294 B.n293 163.367
R1950 B.n294 B.n207 163.367
R1951 B.n298 B.n207 163.367
R1952 B.n299 B.n298 163.367
R1953 B.n300 B.n299 163.367
R1954 B.n300 B.n205 163.367
R1955 B.n304 B.n205 163.367
R1956 B.n305 B.n304 163.367
R1957 B.n306 B.n305 163.367
R1958 B.n306 B.n203 163.367
R1959 B.n310 B.n203 163.367
R1960 B.n311 B.n310 163.367
R1961 B.n312 B.n311 163.367
R1962 B.n312 B.n201 163.367
R1963 B.n316 B.n201 163.367
R1964 B.n317 B.n316 163.367
R1965 B.n318 B.n317 163.367
R1966 B.n318 B.n199 163.367
R1967 B.n322 B.n199 163.367
R1968 B.n323 B.n322 163.367
R1969 B.n324 B.n323 163.367
R1970 B.n324 B.n197 163.367
R1971 B.n328 B.n197 163.367
R1972 B.n329 B.n328 163.367
R1973 B.n177 B.n176 66.3278
R1974 B.n401 B.n400 66.3278
R1975 B.n63 B.n62 66.3278
R1976 B.n57 B.n56 66.3278
R1977 B.n387 B.n177 59.5399
R1978 B.n402 B.n401 59.5399
R1979 B.n726 B.n63 59.5399
R1980 B.n740 B.n57 59.5399
R1981 B.n799 B.n36 34.4981
R1982 B.n667 B.n82 34.4981
R1983 B.n462 B.n461 34.4981
R1984 B.n331 B.n196 34.4981
R1985 B B.n901 18.0485
R1986 B.n800 B.n799 10.6151
R1987 B.n801 B.n800 10.6151
R1988 B.n801 B.n34 10.6151
R1989 B.n805 B.n34 10.6151
R1990 B.n806 B.n805 10.6151
R1991 B.n807 B.n806 10.6151
R1992 B.n807 B.n32 10.6151
R1993 B.n811 B.n32 10.6151
R1994 B.n812 B.n811 10.6151
R1995 B.n813 B.n812 10.6151
R1996 B.n813 B.n30 10.6151
R1997 B.n817 B.n30 10.6151
R1998 B.n818 B.n817 10.6151
R1999 B.n819 B.n818 10.6151
R2000 B.n819 B.n28 10.6151
R2001 B.n823 B.n28 10.6151
R2002 B.n824 B.n823 10.6151
R2003 B.n825 B.n824 10.6151
R2004 B.n825 B.n26 10.6151
R2005 B.n829 B.n26 10.6151
R2006 B.n830 B.n829 10.6151
R2007 B.n831 B.n830 10.6151
R2008 B.n831 B.n24 10.6151
R2009 B.n835 B.n24 10.6151
R2010 B.n836 B.n835 10.6151
R2011 B.n837 B.n836 10.6151
R2012 B.n837 B.n22 10.6151
R2013 B.n841 B.n22 10.6151
R2014 B.n842 B.n841 10.6151
R2015 B.n843 B.n842 10.6151
R2016 B.n843 B.n20 10.6151
R2017 B.n847 B.n20 10.6151
R2018 B.n848 B.n847 10.6151
R2019 B.n849 B.n848 10.6151
R2020 B.n849 B.n18 10.6151
R2021 B.n853 B.n18 10.6151
R2022 B.n854 B.n853 10.6151
R2023 B.n855 B.n854 10.6151
R2024 B.n855 B.n16 10.6151
R2025 B.n859 B.n16 10.6151
R2026 B.n860 B.n859 10.6151
R2027 B.n861 B.n860 10.6151
R2028 B.n861 B.n14 10.6151
R2029 B.n865 B.n14 10.6151
R2030 B.n866 B.n865 10.6151
R2031 B.n867 B.n866 10.6151
R2032 B.n867 B.n12 10.6151
R2033 B.n871 B.n12 10.6151
R2034 B.n872 B.n871 10.6151
R2035 B.n873 B.n872 10.6151
R2036 B.n873 B.n10 10.6151
R2037 B.n877 B.n10 10.6151
R2038 B.n878 B.n877 10.6151
R2039 B.n879 B.n878 10.6151
R2040 B.n879 B.n8 10.6151
R2041 B.n883 B.n8 10.6151
R2042 B.n884 B.n883 10.6151
R2043 B.n885 B.n884 10.6151
R2044 B.n885 B.n6 10.6151
R2045 B.n889 B.n6 10.6151
R2046 B.n890 B.n889 10.6151
R2047 B.n891 B.n890 10.6151
R2048 B.n891 B.n4 10.6151
R2049 B.n895 B.n4 10.6151
R2050 B.n896 B.n895 10.6151
R2051 B.n897 B.n896 10.6151
R2052 B.n897 B.n0 10.6151
R2053 B.n795 B.n36 10.6151
R2054 B.n795 B.n794 10.6151
R2055 B.n794 B.n793 10.6151
R2056 B.n793 B.n38 10.6151
R2057 B.n789 B.n38 10.6151
R2058 B.n789 B.n788 10.6151
R2059 B.n788 B.n787 10.6151
R2060 B.n787 B.n40 10.6151
R2061 B.n783 B.n40 10.6151
R2062 B.n783 B.n782 10.6151
R2063 B.n782 B.n781 10.6151
R2064 B.n781 B.n42 10.6151
R2065 B.n777 B.n42 10.6151
R2066 B.n777 B.n776 10.6151
R2067 B.n776 B.n775 10.6151
R2068 B.n775 B.n44 10.6151
R2069 B.n771 B.n44 10.6151
R2070 B.n771 B.n770 10.6151
R2071 B.n770 B.n769 10.6151
R2072 B.n769 B.n46 10.6151
R2073 B.n765 B.n46 10.6151
R2074 B.n765 B.n764 10.6151
R2075 B.n764 B.n763 10.6151
R2076 B.n763 B.n48 10.6151
R2077 B.n759 B.n48 10.6151
R2078 B.n759 B.n758 10.6151
R2079 B.n758 B.n757 10.6151
R2080 B.n757 B.n50 10.6151
R2081 B.n753 B.n50 10.6151
R2082 B.n753 B.n752 10.6151
R2083 B.n752 B.n751 10.6151
R2084 B.n751 B.n52 10.6151
R2085 B.n747 B.n52 10.6151
R2086 B.n747 B.n746 10.6151
R2087 B.n746 B.n745 10.6151
R2088 B.n745 B.n54 10.6151
R2089 B.n741 B.n54 10.6151
R2090 B.n739 B.n738 10.6151
R2091 B.n738 B.n58 10.6151
R2092 B.n734 B.n58 10.6151
R2093 B.n734 B.n733 10.6151
R2094 B.n733 B.n732 10.6151
R2095 B.n732 B.n60 10.6151
R2096 B.n728 B.n60 10.6151
R2097 B.n728 B.n727 10.6151
R2098 B.n725 B.n64 10.6151
R2099 B.n721 B.n64 10.6151
R2100 B.n721 B.n720 10.6151
R2101 B.n720 B.n719 10.6151
R2102 B.n719 B.n66 10.6151
R2103 B.n715 B.n66 10.6151
R2104 B.n715 B.n714 10.6151
R2105 B.n714 B.n713 10.6151
R2106 B.n713 B.n68 10.6151
R2107 B.n709 B.n68 10.6151
R2108 B.n709 B.n708 10.6151
R2109 B.n708 B.n707 10.6151
R2110 B.n707 B.n70 10.6151
R2111 B.n703 B.n70 10.6151
R2112 B.n703 B.n702 10.6151
R2113 B.n702 B.n701 10.6151
R2114 B.n701 B.n72 10.6151
R2115 B.n697 B.n72 10.6151
R2116 B.n697 B.n696 10.6151
R2117 B.n696 B.n695 10.6151
R2118 B.n695 B.n74 10.6151
R2119 B.n691 B.n74 10.6151
R2120 B.n691 B.n690 10.6151
R2121 B.n690 B.n689 10.6151
R2122 B.n689 B.n76 10.6151
R2123 B.n685 B.n76 10.6151
R2124 B.n685 B.n684 10.6151
R2125 B.n684 B.n683 10.6151
R2126 B.n683 B.n78 10.6151
R2127 B.n679 B.n78 10.6151
R2128 B.n679 B.n678 10.6151
R2129 B.n678 B.n677 10.6151
R2130 B.n677 B.n80 10.6151
R2131 B.n673 B.n80 10.6151
R2132 B.n673 B.n672 10.6151
R2133 B.n672 B.n671 10.6151
R2134 B.n671 B.n82 10.6151
R2135 B.n667 B.n666 10.6151
R2136 B.n666 B.n665 10.6151
R2137 B.n665 B.n84 10.6151
R2138 B.n661 B.n84 10.6151
R2139 B.n661 B.n660 10.6151
R2140 B.n660 B.n659 10.6151
R2141 B.n659 B.n86 10.6151
R2142 B.n655 B.n86 10.6151
R2143 B.n655 B.n654 10.6151
R2144 B.n654 B.n653 10.6151
R2145 B.n653 B.n88 10.6151
R2146 B.n649 B.n88 10.6151
R2147 B.n649 B.n648 10.6151
R2148 B.n648 B.n647 10.6151
R2149 B.n647 B.n90 10.6151
R2150 B.n643 B.n90 10.6151
R2151 B.n643 B.n642 10.6151
R2152 B.n642 B.n641 10.6151
R2153 B.n641 B.n92 10.6151
R2154 B.n637 B.n92 10.6151
R2155 B.n637 B.n636 10.6151
R2156 B.n636 B.n635 10.6151
R2157 B.n635 B.n94 10.6151
R2158 B.n631 B.n94 10.6151
R2159 B.n631 B.n630 10.6151
R2160 B.n630 B.n629 10.6151
R2161 B.n629 B.n96 10.6151
R2162 B.n625 B.n96 10.6151
R2163 B.n625 B.n624 10.6151
R2164 B.n624 B.n623 10.6151
R2165 B.n623 B.n98 10.6151
R2166 B.n619 B.n98 10.6151
R2167 B.n619 B.n618 10.6151
R2168 B.n618 B.n617 10.6151
R2169 B.n617 B.n100 10.6151
R2170 B.n613 B.n100 10.6151
R2171 B.n613 B.n612 10.6151
R2172 B.n612 B.n611 10.6151
R2173 B.n611 B.n102 10.6151
R2174 B.n607 B.n102 10.6151
R2175 B.n607 B.n606 10.6151
R2176 B.n606 B.n605 10.6151
R2177 B.n605 B.n104 10.6151
R2178 B.n601 B.n104 10.6151
R2179 B.n601 B.n600 10.6151
R2180 B.n600 B.n599 10.6151
R2181 B.n599 B.n106 10.6151
R2182 B.n595 B.n106 10.6151
R2183 B.n595 B.n594 10.6151
R2184 B.n594 B.n593 10.6151
R2185 B.n593 B.n108 10.6151
R2186 B.n589 B.n108 10.6151
R2187 B.n589 B.n588 10.6151
R2188 B.n588 B.n587 10.6151
R2189 B.n587 B.n110 10.6151
R2190 B.n583 B.n110 10.6151
R2191 B.n583 B.n582 10.6151
R2192 B.n582 B.n581 10.6151
R2193 B.n581 B.n112 10.6151
R2194 B.n577 B.n112 10.6151
R2195 B.n577 B.n576 10.6151
R2196 B.n576 B.n575 10.6151
R2197 B.n575 B.n114 10.6151
R2198 B.n571 B.n114 10.6151
R2199 B.n571 B.n570 10.6151
R2200 B.n570 B.n569 10.6151
R2201 B.n569 B.n116 10.6151
R2202 B.n565 B.n116 10.6151
R2203 B.n565 B.n564 10.6151
R2204 B.n564 B.n563 10.6151
R2205 B.n563 B.n118 10.6151
R2206 B.n559 B.n118 10.6151
R2207 B.n559 B.n558 10.6151
R2208 B.n558 B.n557 10.6151
R2209 B.n557 B.n120 10.6151
R2210 B.n553 B.n120 10.6151
R2211 B.n553 B.n552 10.6151
R2212 B.n552 B.n551 10.6151
R2213 B.n551 B.n122 10.6151
R2214 B.n547 B.n122 10.6151
R2215 B.n547 B.n546 10.6151
R2216 B.n546 B.n545 10.6151
R2217 B.n545 B.n124 10.6151
R2218 B.n541 B.n124 10.6151
R2219 B.n541 B.n540 10.6151
R2220 B.n540 B.n539 10.6151
R2221 B.n539 B.n126 10.6151
R2222 B.n535 B.n126 10.6151
R2223 B.n535 B.n534 10.6151
R2224 B.n534 B.n533 10.6151
R2225 B.n533 B.n128 10.6151
R2226 B.n529 B.n128 10.6151
R2227 B.n529 B.n528 10.6151
R2228 B.n528 B.n527 10.6151
R2229 B.n527 B.n130 10.6151
R2230 B.n523 B.n130 10.6151
R2231 B.n523 B.n522 10.6151
R2232 B.n522 B.n521 10.6151
R2233 B.n521 B.n132 10.6151
R2234 B.n517 B.n132 10.6151
R2235 B.n517 B.n516 10.6151
R2236 B.n516 B.n515 10.6151
R2237 B.n515 B.n134 10.6151
R2238 B.n511 B.n134 10.6151
R2239 B.n511 B.n510 10.6151
R2240 B.n510 B.n509 10.6151
R2241 B.n509 B.n136 10.6151
R2242 B.n505 B.n136 10.6151
R2243 B.n505 B.n504 10.6151
R2244 B.n504 B.n503 10.6151
R2245 B.n503 B.n138 10.6151
R2246 B.n499 B.n138 10.6151
R2247 B.n499 B.n498 10.6151
R2248 B.n498 B.n497 10.6151
R2249 B.n497 B.n140 10.6151
R2250 B.n493 B.n140 10.6151
R2251 B.n493 B.n492 10.6151
R2252 B.n492 B.n491 10.6151
R2253 B.n491 B.n142 10.6151
R2254 B.n487 B.n142 10.6151
R2255 B.n487 B.n486 10.6151
R2256 B.n486 B.n485 10.6151
R2257 B.n485 B.n144 10.6151
R2258 B.n481 B.n144 10.6151
R2259 B.n481 B.n480 10.6151
R2260 B.n480 B.n479 10.6151
R2261 B.n479 B.n146 10.6151
R2262 B.n475 B.n146 10.6151
R2263 B.n475 B.n474 10.6151
R2264 B.n474 B.n473 10.6151
R2265 B.n473 B.n148 10.6151
R2266 B.n469 B.n148 10.6151
R2267 B.n469 B.n468 10.6151
R2268 B.n468 B.n467 10.6151
R2269 B.n467 B.n150 10.6151
R2270 B.n463 B.n150 10.6151
R2271 B.n463 B.n462 10.6151
R2272 B.n230 B.n1 10.6151
R2273 B.n231 B.n230 10.6151
R2274 B.n231 B.n228 10.6151
R2275 B.n235 B.n228 10.6151
R2276 B.n236 B.n235 10.6151
R2277 B.n237 B.n236 10.6151
R2278 B.n237 B.n226 10.6151
R2279 B.n241 B.n226 10.6151
R2280 B.n242 B.n241 10.6151
R2281 B.n243 B.n242 10.6151
R2282 B.n243 B.n224 10.6151
R2283 B.n247 B.n224 10.6151
R2284 B.n248 B.n247 10.6151
R2285 B.n249 B.n248 10.6151
R2286 B.n249 B.n222 10.6151
R2287 B.n253 B.n222 10.6151
R2288 B.n254 B.n253 10.6151
R2289 B.n255 B.n254 10.6151
R2290 B.n255 B.n220 10.6151
R2291 B.n259 B.n220 10.6151
R2292 B.n260 B.n259 10.6151
R2293 B.n261 B.n260 10.6151
R2294 B.n261 B.n218 10.6151
R2295 B.n265 B.n218 10.6151
R2296 B.n266 B.n265 10.6151
R2297 B.n267 B.n266 10.6151
R2298 B.n267 B.n216 10.6151
R2299 B.n271 B.n216 10.6151
R2300 B.n272 B.n271 10.6151
R2301 B.n273 B.n272 10.6151
R2302 B.n273 B.n214 10.6151
R2303 B.n277 B.n214 10.6151
R2304 B.n278 B.n277 10.6151
R2305 B.n279 B.n278 10.6151
R2306 B.n279 B.n212 10.6151
R2307 B.n283 B.n212 10.6151
R2308 B.n284 B.n283 10.6151
R2309 B.n285 B.n284 10.6151
R2310 B.n285 B.n210 10.6151
R2311 B.n289 B.n210 10.6151
R2312 B.n290 B.n289 10.6151
R2313 B.n291 B.n290 10.6151
R2314 B.n291 B.n208 10.6151
R2315 B.n295 B.n208 10.6151
R2316 B.n296 B.n295 10.6151
R2317 B.n297 B.n296 10.6151
R2318 B.n297 B.n206 10.6151
R2319 B.n301 B.n206 10.6151
R2320 B.n302 B.n301 10.6151
R2321 B.n303 B.n302 10.6151
R2322 B.n303 B.n204 10.6151
R2323 B.n307 B.n204 10.6151
R2324 B.n308 B.n307 10.6151
R2325 B.n309 B.n308 10.6151
R2326 B.n309 B.n202 10.6151
R2327 B.n313 B.n202 10.6151
R2328 B.n314 B.n313 10.6151
R2329 B.n315 B.n314 10.6151
R2330 B.n315 B.n200 10.6151
R2331 B.n319 B.n200 10.6151
R2332 B.n320 B.n319 10.6151
R2333 B.n321 B.n320 10.6151
R2334 B.n321 B.n198 10.6151
R2335 B.n325 B.n198 10.6151
R2336 B.n326 B.n325 10.6151
R2337 B.n327 B.n326 10.6151
R2338 B.n327 B.n196 10.6151
R2339 B.n332 B.n331 10.6151
R2340 B.n333 B.n332 10.6151
R2341 B.n333 B.n194 10.6151
R2342 B.n337 B.n194 10.6151
R2343 B.n338 B.n337 10.6151
R2344 B.n339 B.n338 10.6151
R2345 B.n339 B.n192 10.6151
R2346 B.n343 B.n192 10.6151
R2347 B.n344 B.n343 10.6151
R2348 B.n345 B.n344 10.6151
R2349 B.n345 B.n190 10.6151
R2350 B.n349 B.n190 10.6151
R2351 B.n350 B.n349 10.6151
R2352 B.n351 B.n350 10.6151
R2353 B.n351 B.n188 10.6151
R2354 B.n355 B.n188 10.6151
R2355 B.n356 B.n355 10.6151
R2356 B.n357 B.n356 10.6151
R2357 B.n357 B.n186 10.6151
R2358 B.n361 B.n186 10.6151
R2359 B.n362 B.n361 10.6151
R2360 B.n363 B.n362 10.6151
R2361 B.n363 B.n184 10.6151
R2362 B.n367 B.n184 10.6151
R2363 B.n368 B.n367 10.6151
R2364 B.n369 B.n368 10.6151
R2365 B.n369 B.n182 10.6151
R2366 B.n373 B.n182 10.6151
R2367 B.n374 B.n373 10.6151
R2368 B.n375 B.n374 10.6151
R2369 B.n375 B.n180 10.6151
R2370 B.n379 B.n180 10.6151
R2371 B.n380 B.n379 10.6151
R2372 B.n381 B.n380 10.6151
R2373 B.n381 B.n178 10.6151
R2374 B.n385 B.n178 10.6151
R2375 B.n386 B.n385 10.6151
R2376 B.n388 B.n174 10.6151
R2377 B.n392 B.n174 10.6151
R2378 B.n393 B.n392 10.6151
R2379 B.n394 B.n393 10.6151
R2380 B.n394 B.n172 10.6151
R2381 B.n398 B.n172 10.6151
R2382 B.n399 B.n398 10.6151
R2383 B.n403 B.n399 10.6151
R2384 B.n407 B.n170 10.6151
R2385 B.n408 B.n407 10.6151
R2386 B.n409 B.n408 10.6151
R2387 B.n409 B.n168 10.6151
R2388 B.n413 B.n168 10.6151
R2389 B.n414 B.n413 10.6151
R2390 B.n415 B.n414 10.6151
R2391 B.n415 B.n166 10.6151
R2392 B.n419 B.n166 10.6151
R2393 B.n420 B.n419 10.6151
R2394 B.n421 B.n420 10.6151
R2395 B.n421 B.n164 10.6151
R2396 B.n425 B.n164 10.6151
R2397 B.n426 B.n425 10.6151
R2398 B.n427 B.n426 10.6151
R2399 B.n427 B.n162 10.6151
R2400 B.n431 B.n162 10.6151
R2401 B.n432 B.n431 10.6151
R2402 B.n433 B.n432 10.6151
R2403 B.n433 B.n160 10.6151
R2404 B.n437 B.n160 10.6151
R2405 B.n438 B.n437 10.6151
R2406 B.n439 B.n438 10.6151
R2407 B.n439 B.n158 10.6151
R2408 B.n443 B.n158 10.6151
R2409 B.n444 B.n443 10.6151
R2410 B.n445 B.n444 10.6151
R2411 B.n445 B.n156 10.6151
R2412 B.n449 B.n156 10.6151
R2413 B.n450 B.n449 10.6151
R2414 B.n451 B.n450 10.6151
R2415 B.n451 B.n154 10.6151
R2416 B.n455 B.n154 10.6151
R2417 B.n456 B.n455 10.6151
R2418 B.n457 B.n456 10.6151
R2419 B.n457 B.n152 10.6151
R2420 B.n461 B.n152 10.6151
R2421 B.n901 B.n0 8.11757
R2422 B.n901 B.n1 8.11757
R2423 B.n740 B.n739 6.5566
R2424 B.n727 B.n726 6.5566
R2425 B.n388 B.n387 6.5566
R2426 B.n403 B.n402 6.5566
R2427 B.n741 B.n740 4.05904
R2428 B.n726 B.n725 4.05904
R2429 B.n387 B.n386 4.05904
R2430 B.n402 B.n170 4.05904
C0 VDD2 B 2.70891f
C1 VP w_n5074_n3118# 11.6439f
C2 VN w_n5074_n3118# 10.9818f
C3 VDD1 w_n5074_n3118# 2.89069f
C4 VP VN 8.892469f
C5 VP VDD1 10.406099f
C6 VTAIL w_n5074_n3118# 3.11171f
C7 VN VDD1 0.154577f
C8 VP VTAIL 10.843401f
C9 VN VTAIL 10.8292f
C10 VTAIL VDD1 10.036f
C11 VDD2 w_n5074_n3118# 3.05971f
C12 VP VDD2 0.646101f
C13 w_n5074_n3118# B 11.0205f
C14 VP B 2.50937f
C15 VN VDD2 9.918231f
C16 VDD1 VDD2 2.49408f
C17 VN B 1.39327f
C18 VDD1 B 2.57191f
C19 VTAIL VDD2 10.0909f
C20 VTAIL B 3.63694f
C21 VDD2 VSUBS 2.33155f
C22 VDD1 VSUBS 2.131503f
C23 VTAIL VSUBS 1.381538f
C24 VN VSUBS 8.47552f
C25 VP VSUBS 4.826609f
C26 B VSUBS 5.869558f
C27 w_n5074_n3118# VSUBS 0.195146p
C28 B.n0 VSUBS 0.008338f
C29 B.n1 VSUBS 0.008338f
C30 B.n2 VSUBS 0.012332f
C31 B.n3 VSUBS 0.00945f
C32 B.n4 VSUBS 0.00945f
C33 B.n5 VSUBS 0.00945f
C34 B.n6 VSUBS 0.00945f
C35 B.n7 VSUBS 0.00945f
C36 B.n8 VSUBS 0.00945f
C37 B.n9 VSUBS 0.00945f
C38 B.n10 VSUBS 0.00945f
C39 B.n11 VSUBS 0.00945f
C40 B.n12 VSUBS 0.00945f
C41 B.n13 VSUBS 0.00945f
C42 B.n14 VSUBS 0.00945f
C43 B.n15 VSUBS 0.00945f
C44 B.n16 VSUBS 0.00945f
C45 B.n17 VSUBS 0.00945f
C46 B.n18 VSUBS 0.00945f
C47 B.n19 VSUBS 0.00945f
C48 B.n20 VSUBS 0.00945f
C49 B.n21 VSUBS 0.00945f
C50 B.n22 VSUBS 0.00945f
C51 B.n23 VSUBS 0.00945f
C52 B.n24 VSUBS 0.00945f
C53 B.n25 VSUBS 0.00945f
C54 B.n26 VSUBS 0.00945f
C55 B.n27 VSUBS 0.00945f
C56 B.n28 VSUBS 0.00945f
C57 B.n29 VSUBS 0.00945f
C58 B.n30 VSUBS 0.00945f
C59 B.n31 VSUBS 0.00945f
C60 B.n32 VSUBS 0.00945f
C61 B.n33 VSUBS 0.00945f
C62 B.n34 VSUBS 0.00945f
C63 B.n35 VSUBS 0.00945f
C64 B.n36 VSUBS 0.023201f
C65 B.n37 VSUBS 0.00945f
C66 B.n38 VSUBS 0.00945f
C67 B.n39 VSUBS 0.00945f
C68 B.n40 VSUBS 0.00945f
C69 B.n41 VSUBS 0.00945f
C70 B.n42 VSUBS 0.00945f
C71 B.n43 VSUBS 0.00945f
C72 B.n44 VSUBS 0.00945f
C73 B.n45 VSUBS 0.00945f
C74 B.n46 VSUBS 0.00945f
C75 B.n47 VSUBS 0.00945f
C76 B.n48 VSUBS 0.00945f
C77 B.n49 VSUBS 0.00945f
C78 B.n50 VSUBS 0.00945f
C79 B.n51 VSUBS 0.00945f
C80 B.n52 VSUBS 0.00945f
C81 B.n53 VSUBS 0.00945f
C82 B.n54 VSUBS 0.00945f
C83 B.n55 VSUBS 0.00945f
C84 B.t4 VSUBS 0.247933f
C85 B.t5 VSUBS 0.296187f
C86 B.t3 VSUBS 2.07865f
C87 B.n56 VSUBS 0.475821f
C88 B.n57 VSUBS 0.318671f
C89 B.n58 VSUBS 0.00945f
C90 B.n59 VSUBS 0.00945f
C91 B.n60 VSUBS 0.00945f
C92 B.n61 VSUBS 0.00945f
C93 B.t7 VSUBS 0.247937f
C94 B.t8 VSUBS 0.29619f
C95 B.t6 VSUBS 2.07865f
C96 B.n62 VSUBS 0.475818f
C97 B.n63 VSUBS 0.318667f
C98 B.n64 VSUBS 0.00945f
C99 B.n65 VSUBS 0.00945f
C100 B.n66 VSUBS 0.00945f
C101 B.n67 VSUBS 0.00945f
C102 B.n68 VSUBS 0.00945f
C103 B.n69 VSUBS 0.00945f
C104 B.n70 VSUBS 0.00945f
C105 B.n71 VSUBS 0.00945f
C106 B.n72 VSUBS 0.00945f
C107 B.n73 VSUBS 0.00945f
C108 B.n74 VSUBS 0.00945f
C109 B.n75 VSUBS 0.00945f
C110 B.n76 VSUBS 0.00945f
C111 B.n77 VSUBS 0.00945f
C112 B.n78 VSUBS 0.00945f
C113 B.n79 VSUBS 0.00945f
C114 B.n80 VSUBS 0.00945f
C115 B.n81 VSUBS 0.00945f
C116 B.n82 VSUBS 0.023201f
C117 B.n83 VSUBS 0.00945f
C118 B.n84 VSUBS 0.00945f
C119 B.n85 VSUBS 0.00945f
C120 B.n86 VSUBS 0.00945f
C121 B.n87 VSUBS 0.00945f
C122 B.n88 VSUBS 0.00945f
C123 B.n89 VSUBS 0.00945f
C124 B.n90 VSUBS 0.00945f
C125 B.n91 VSUBS 0.00945f
C126 B.n92 VSUBS 0.00945f
C127 B.n93 VSUBS 0.00945f
C128 B.n94 VSUBS 0.00945f
C129 B.n95 VSUBS 0.00945f
C130 B.n96 VSUBS 0.00945f
C131 B.n97 VSUBS 0.00945f
C132 B.n98 VSUBS 0.00945f
C133 B.n99 VSUBS 0.00945f
C134 B.n100 VSUBS 0.00945f
C135 B.n101 VSUBS 0.00945f
C136 B.n102 VSUBS 0.00945f
C137 B.n103 VSUBS 0.00945f
C138 B.n104 VSUBS 0.00945f
C139 B.n105 VSUBS 0.00945f
C140 B.n106 VSUBS 0.00945f
C141 B.n107 VSUBS 0.00945f
C142 B.n108 VSUBS 0.00945f
C143 B.n109 VSUBS 0.00945f
C144 B.n110 VSUBS 0.00945f
C145 B.n111 VSUBS 0.00945f
C146 B.n112 VSUBS 0.00945f
C147 B.n113 VSUBS 0.00945f
C148 B.n114 VSUBS 0.00945f
C149 B.n115 VSUBS 0.00945f
C150 B.n116 VSUBS 0.00945f
C151 B.n117 VSUBS 0.00945f
C152 B.n118 VSUBS 0.00945f
C153 B.n119 VSUBS 0.00945f
C154 B.n120 VSUBS 0.00945f
C155 B.n121 VSUBS 0.00945f
C156 B.n122 VSUBS 0.00945f
C157 B.n123 VSUBS 0.00945f
C158 B.n124 VSUBS 0.00945f
C159 B.n125 VSUBS 0.00945f
C160 B.n126 VSUBS 0.00945f
C161 B.n127 VSUBS 0.00945f
C162 B.n128 VSUBS 0.00945f
C163 B.n129 VSUBS 0.00945f
C164 B.n130 VSUBS 0.00945f
C165 B.n131 VSUBS 0.00945f
C166 B.n132 VSUBS 0.00945f
C167 B.n133 VSUBS 0.00945f
C168 B.n134 VSUBS 0.00945f
C169 B.n135 VSUBS 0.00945f
C170 B.n136 VSUBS 0.00945f
C171 B.n137 VSUBS 0.00945f
C172 B.n138 VSUBS 0.00945f
C173 B.n139 VSUBS 0.00945f
C174 B.n140 VSUBS 0.00945f
C175 B.n141 VSUBS 0.00945f
C176 B.n142 VSUBS 0.00945f
C177 B.n143 VSUBS 0.00945f
C178 B.n144 VSUBS 0.00945f
C179 B.n145 VSUBS 0.00945f
C180 B.n146 VSUBS 0.00945f
C181 B.n147 VSUBS 0.00945f
C182 B.n148 VSUBS 0.00945f
C183 B.n149 VSUBS 0.00945f
C184 B.n150 VSUBS 0.00945f
C185 B.n151 VSUBS 0.02266f
C186 B.n152 VSUBS 0.00945f
C187 B.n153 VSUBS 0.00945f
C188 B.n154 VSUBS 0.00945f
C189 B.n155 VSUBS 0.00945f
C190 B.n156 VSUBS 0.00945f
C191 B.n157 VSUBS 0.00945f
C192 B.n158 VSUBS 0.00945f
C193 B.n159 VSUBS 0.00945f
C194 B.n160 VSUBS 0.00945f
C195 B.n161 VSUBS 0.00945f
C196 B.n162 VSUBS 0.00945f
C197 B.n163 VSUBS 0.00945f
C198 B.n164 VSUBS 0.00945f
C199 B.n165 VSUBS 0.00945f
C200 B.n166 VSUBS 0.00945f
C201 B.n167 VSUBS 0.00945f
C202 B.n168 VSUBS 0.00945f
C203 B.n169 VSUBS 0.00945f
C204 B.n170 VSUBS 0.006532f
C205 B.n171 VSUBS 0.00945f
C206 B.n172 VSUBS 0.00945f
C207 B.n173 VSUBS 0.00945f
C208 B.n174 VSUBS 0.00945f
C209 B.n175 VSUBS 0.00945f
C210 B.t11 VSUBS 0.247933f
C211 B.t10 VSUBS 0.296187f
C212 B.t9 VSUBS 2.07865f
C213 B.n176 VSUBS 0.475821f
C214 B.n177 VSUBS 0.318671f
C215 B.n178 VSUBS 0.00945f
C216 B.n179 VSUBS 0.00945f
C217 B.n180 VSUBS 0.00945f
C218 B.n181 VSUBS 0.00945f
C219 B.n182 VSUBS 0.00945f
C220 B.n183 VSUBS 0.00945f
C221 B.n184 VSUBS 0.00945f
C222 B.n185 VSUBS 0.00945f
C223 B.n186 VSUBS 0.00945f
C224 B.n187 VSUBS 0.00945f
C225 B.n188 VSUBS 0.00945f
C226 B.n189 VSUBS 0.00945f
C227 B.n190 VSUBS 0.00945f
C228 B.n191 VSUBS 0.00945f
C229 B.n192 VSUBS 0.00945f
C230 B.n193 VSUBS 0.00945f
C231 B.n194 VSUBS 0.00945f
C232 B.n195 VSUBS 0.00945f
C233 B.n196 VSUBS 0.02266f
C234 B.n197 VSUBS 0.00945f
C235 B.n198 VSUBS 0.00945f
C236 B.n199 VSUBS 0.00945f
C237 B.n200 VSUBS 0.00945f
C238 B.n201 VSUBS 0.00945f
C239 B.n202 VSUBS 0.00945f
C240 B.n203 VSUBS 0.00945f
C241 B.n204 VSUBS 0.00945f
C242 B.n205 VSUBS 0.00945f
C243 B.n206 VSUBS 0.00945f
C244 B.n207 VSUBS 0.00945f
C245 B.n208 VSUBS 0.00945f
C246 B.n209 VSUBS 0.00945f
C247 B.n210 VSUBS 0.00945f
C248 B.n211 VSUBS 0.00945f
C249 B.n212 VSUBS 0.00945f
C250 B.n213 VSUBS 0.00945f
C251 B.n214 VSUBS 0.00945f
C252 B.n215 VSUBS 0.00945f
C253 B.n216 VSUBS 0.00945f
C254 B.n217 VSUBS 0.00945f
C255 B.n218 VSUBS 0.00945f
C256 B.n219 VSUBS 0.00945f
C257 B.n220 VSUBS 0.00945f
C258 B.n221 VSUBS 0.00945f
C259 B.n222 VSUBS 0.00945f
C260 B.n223 VSUBS 0.00945f
C261 B.n224 VSUBS 0.00945f
C262 B.n225 VSUBS 0.00945f
C263 B.n226 VSUBS 0.00945f
C264 B.n227 VSUBS 0.00945f
C265 B.n228 VSUBS 0.00945f
C266 B.n229 VSUBS 0.00945f
C267 B.n230 VSUBS 0.00945f
C268 B.n231 VSUBS 0.00945f
C269 B.n232 VSUBS 0.00945f
C270 B.n233 VSUBS 0.00945f
C271 B.n234 VSUBS 0.00945f
C272 B.n235 VSUBS 0.00945f
C273 B.n236 VSUBS 0.00945f
C274 B.n237 VSUBS 0.00945f
C275 B.n238 VSUBS 0.00945f
C276 B.n239 VSUBS 0.00945f
C277 B.n240 VSUBS 0.00945f
C278 B.n241 VSUBS 0.00945f
C279 B.n242 VSUBS 0.00945f
C280 B.n243 VSUBS 0.00945f
C281 B.n244 VSUBS 0.00945f
C282 B.n245 VSUBS 0.00945f
C283 B.n246 VSUBS 0.00945f
C284 B.n247 VSUBS 0.00945f
C285 B.n248 VSUBS 0.00945f
C286 B.n249 VSUBS 0.00945f
C287 B.n250 VSUBS 0.00945f
C288 B.n251 VSUBS 0.00945f
C289 B.n252 VSUBS 0.00945f
C290 B.n253 VSUBS 0.00945f
C291 B.n254 VSUBS 0.00945f
C292 B.n255 VSUBS 0.00945f
C293 B.n256 VSUBS 0.00945f
C294 B.n257 VSUBS 0.00945f
C295 B.n258 VSUBS 0.00945f
C296 B.n259 VSUBS 0.00945f
C297 B.n260 VSUBS 0.00945f
C298 B.n261 VSUBS 0.00945f
C299 B.n262 VSUBS 0.00945f
C300 B.n263 VSUBS 0.00945f
C301 B.n264 VSUBS 0.00945f
C302 B.n265 VSUBS 0.00945f
C303 B.n266 VSUBS 0.00945f
C304 B.n267 VSUBS 0.00945f
C305 B.n268 VSUBS 0.00945f
C306 B.n269 VSUBS 0.00945f
C307 B.n270 VSUBS 0.00945f
C308 B.n271 VSUBS 0.00945f
C309 B.n272 VSUBS 0.00945f
C310 B.n273 VSUBS 0.00945f
C311 B.n274 VSUBS 0.00945f
C312 B.n275 VSUBS 0.00945f
C313 B.n276 VSUBS 0.00945f
C314 B.n277 VSUBS 0.00945f
C315 B.n278 VSUBS 0.00945f
C316 B.n279 VSUBS 0.00945f
C317 B.n280 VSUBS 0.00945f
C318 B.n281 VSUBS 0.00945f
C319 B.n282 VSUBS 0.00945f
C320 B.n283 VSUBS 0.00945f
C321 B.n284 VSUBS 0.00945f
C322 B.n285 VSUBS 0.00945f
C323 B.n286 VSUBS 0.00945f
C324 B.n287 VSUBS 0.00945f
C325 B.n288 VSUBS 0.00945f
C326 B.n289 VSUBS 0.00945f
C327 B.n290 VSUBS 0.00945f
C328 B.n291 VSUBS 0.00945f
C329 B.n292 VSUBS 0.00945f
C330 B.n293 VSUBS 0.00945f
C331 B.n294 VSUBS 0.00945f
C332 B.n295 VSUBS 0.00945f
C333 B.n296 VSUBS 0.00945f
C334 B.n297 VSUBS 0.00945f
C335 B.n298 VSUBS 0.00945f
C336 B.n299 VSUBS 0.00945f
C337 B.n300 VSUBS 0.00945f
C338 B.n301 VSUBS 0.00945f
C339 B.n302 VSUBS 0.00945f
C340 B.n303 VSUBS 0.00945f
C341 B.n304 VSUBS 0.00945f
C342 B.n305 VSUBS 0.00945f
C343 B.n306 VSUBS 0.00945f
C344 B.n307 VSUBS 0.00945f
C345 B.n308 VSUBS 0.00945f
C346 B.n309 VSUBS 0.00945f
C347 B.n310 VSUBS 0.00945f
C348 B.n311 VSUBS 0.00945f
C349 B.n312 VSUBS 0.00945f
C350 B.n313 VSUBS 0.00945f
C351 B.n314 VSUBS 0.00945f
C352 B.n315 VSUBS 0.00945f
C353 B.n316 VSUBS 0.00945f
C354 B.n317 VSUBS 0.00945f
C355 B.n318 VSUBS 0.00945f
C356 B.n319 VSUBS 0.00945f
C357 B.n320 VSUBS 0.00945f
C358 B.n321 VSUBS 0.00945f
C359 B.n322 VSUBS 0.00945f
C360 B.n323 VSUBS 0.00945f
C361 B.n324 VSUBS 0.00945f
C362 B.n325 VSUBS 0.00945f
C363 B.n326 VSUBS 0.00945f
C364 B.n327 VSUBS 0.00945f
C365 B.n328 VSUBS 0.00945f
C366 B.n329 VSUBS 0.02266f
C367 B.n330 VSUBS 0.023201f
C368 B.n331 VSUBS 0.023201f
C369 B.n332 VSUBS 0.00945f
C370 B.n333 VSUBS 0.00945f
C371 B.n334 VSUBS 0.00945f
C372 B.n335 VSUBS 0.00945f
C373 B.n336 VSUBS 0.00945f
C374 B.n337 VSUBS 0.00945f
C375 B.n338 VSUBS 0.00945f
C376 B.n339 VSUBS 0.00945f
C377 B.n340 VSUBS 0.00945f
C378 B.n341 VSUBS 0.00945f
C379 B.n342 VSUBS 0.00945f
C380 B.n343 VSUBS 0.00945f
C381 B.n344 VSUBS 0.00945f
C382 B.n345 VSUBS 0.00945f
C383 B.n346 VSUBS 0.00945f
C384 B.n347 VSUBS 0.00945f
C385 B.n348 VSUBS 0.00945f
C386 B.n349 VSUBS 0.00945f
C387 B.n350 VSUBS 0.00945f
C388 B.n351 VSUBS 0.00945f
C389 B.n352 VSUBS 0.00945f
C390 B.n353 VSUBS 0.00945f
C391 B.n354 VSUBS 0.00945f
C392 B.n355 VSUBS 0.00945f
C393 B.n356 VSUBS 0.00945f
C394 B.n357 VSUBS 0.00945f
C395 B.n358 VSUBS 0.00945f
C396 B.n359 VSUBS 0.00945f
C397 B.n360 VSUBS 0.00945f
C398 B.n361 VSUBS 0.00945f
C399 B.n362 VSUBS 0.00945f
C400 B.n363 VSUBS 0.00945f
C401 B.n364 VSUBS 0.00945f
C402 B.n365 VSUBS 0.00945f
C403 B.n366 VSUBS 0.00945f
C404 B.n367 VSUBS 0.00945f
C405 B.n368 VSUBS 0.00945f
C406 B.n369 VSUBS 0.00945f
C407 B.n370 VSUBS 0.00945f
C408 B.n371 VSUBS 0.00945f
C409 B.n372 VSUBS 0.00945f
C410 B.n373 VSUBS 0.00945f
C411 B.n374 VSUBS 0.00945f
C412 B.n375 VSUBS 0.00945f
C413 B.n376 VSUBS 0.00945f
C414 B.n377 VSUBS 0.00945f
C415 B.n378 VSUBS 0.00945f
C416 B.n379 VSUBS 0.00945f
C417 B.n380 VSUBS 0.00945f
C418 B.n381 VSUBS 0.00945f
C419 B.n382 VSUBS 0.00945f
C420 B.n383 VSUBS 0.00945f
C421 B.n384 VSUBS 0.00945f
C422 B.n385 VSUBS 0.00945f
C423 B.n386 VSUBS 0.006532f
C424 B.n387 VSUBS 0.021895f
C425 B.n388 VSUBS 0.007644f
C426 B.n389 VSUBS 0.00945f
C427 B.n390 VSUBS 0.00945f
C428 B.n391 VSUBS 0.00945f
C429 B.n392 VSUBS 0.00945f
C430 B.n393 VSUBS 0.00945f
C431 B.n394 VSUBS 0.00945f
C432 B.n395 VSUBS 0.00945f
C433 B.n396 VSUBS 0.00945f
C434 B.n397 VSUBS 0.00945f
C435 B.n398 VSUBS 0.00945f
C436 B.n399 VSUBS 0.00945f
C437 B.t2 VSUBS 0.247937f
C438 B.t1 VSUBS 0.29619f
C439 B.t0 VSUBS 2.07865f
C440 B.n400 VSUBS 0.475818f
C441 B.n401 VSUBS 0.318667f
C442 B.n402 VSUBS 0.021895f
C443 B.n403 VSUBS 0.007644f
C444 B.n404 VSUBS 0.00945f
C445 B.n405 VSUBS 0.00945f
C446 B.n406 VSUBS 0.00945f
C447 B.n407 VSUBS 0.00945f
C448 B.n408 VSUBS 0.00945f
C449 B.n409 VSUBS 0.00945f
C450 B.n410 VSUBS 0.00945f
C451 B.n411 VSUBS 0.00945f
C452 B.n412 VSUBS 0.00945f
C453 B.n413 VSUBS 0.00945f
C454 B.n414 VSUBS 0.00945f
C455 B.n415 VSUBS 0.00945f
C456 B.n416 VSUBS 0.00945f
C457 B.n417 VSUBS 0.00945f
C458 B.n418 VSUBS 0.00945f
C459 B.n419 VSUBS 0.00945f
C460 B.n420 VSUBS 0.00945f
C461 B.n421 VSUBS 0.00945f
C462 B.n422 VSUBS 0.00945f
C463 B.n423 VSUBS 0.00945f
C464 B.n424 VSUBS 0.00945f
C465 B.n425 VSUBS 0.00945f
C466 B.n426 VSUBS 0.00945f
C467 B.n427 VSUBS 0.00945f
C468 B.n428 VSUBS 0.00945f
C469 B.n429 VSUBS 0.00945f
C470 B.n430 VSUBS 0.00945f
C471 B.n431 VSUBS 0.00945f
C472 B.n432 VSUBS 0.00945f
C473 B.n433 VSUBS 0.00945f
C474 B.n434 VSUBS 0.00945f
C475 B.n435 VSUBS 0.00945f
C476 B.n436 VSUBS 0.00945f
C477 B.n437 VSUBS 0.00945f
C478 B.n438 VSUBS 0.00945f
C479 B.n439 VSUBS 0.00945f
C480 B.n440 VSUBS 0.00945f
C481 B.n441 VSUBS 0.00945f
C482 B.n442 VSUBS 0.00945f
C483 B.n443 VSUBS 0.00945f
C484 B.n444 VSUBS 0.00945f
C485 B.n445 VSUBS 0.00945f
C486 B.n446 VSUBS 0.00945f
C487 B.n447 VSUBS 0.00945f
C488 B.n448 VSUBS 0.00945f
C489 B.n449 VSUBS 0.00945f
C490 B.n450 VSUBS 0.00945f
C491 B.n451 VSUBS 0.00945f
C492 B.n452 VSUBS 0.00945f
C493 B.n453 VSUBS 0.00945f
C494 B.n454 VSUBS 0.00945f
C495 B.n455 VSUBS 0.00945f
C496 B.n456 VSUBS 0.00945f
C497 B.n457 VSUBS 0.00945f
C498 B.n458 VSUBS 0.00945f
C499 B.n459 VSUBS 0.00945f
C500 B.n460 VSUBS 0.023201f
C501 B.n461 VSUBS 0.022144f
C502 B.n462 VSUBS 0.023717f
C503 B.n463 VSUBS 0.00945f
C504 B.n464 VSUBS 0.00945f
C505 B.n465 VSUBS 0.00945f
C506 B.n466 VSUBS 0.00945f
C507 B.n467 VSUBS 0.00945f
C508 B.n468 VSUBS 0.00945f
C509 B.n469 VSUBS 0.00945f
C510 B.n470 VSUBS 0.00945f
C511 B.n471 VSUBS 0.00945f
C512 B.n472 VSUBS 0.00945f
C513 B.n473 VSUBS 0.00945f
C514 B.n474 VSUBS 0.00945f
C515 B.n475 VSUBS 0.00945f
C516 B.n476 VSUBS 0.00945f
C517 B.n477 VSUBS 0.00945f
C518 B.n478 VSUBS 0.00945f
C519 B.n479 VSUBS 0.00945f
C520 B.n480 VSUBS 0.00945f
C521 B.n481 VSUBS 0.00945f
C522 B.n482 VSUBS 0.00945f
C523 B.n483 VSUBS 0.00945f
C524 B.n484 VSUBS 0.00945f
C525 B.n485 VSUBS 0.00945f
C526 B.n486 VSUBS 0.00945f
C527 B.n487 VSUBS 0.00945f
C528 B.n488 VSUBS 0.00945f
C529 B.n489 VSUBS 0.00945f
C530 B.n490 VSUBS 0.00945f
C531 B.n491 VSUBS 0.00945f
C532 B.n492 VSUBS 0.00945f
C533 B.n493 VSUBS 0.00945f
C534 B.n494 VSUBS 0.00945f
C535 B.n495 VSUBS 0.00945f
C536 B.n496 VSUBS 0.00945f
C537 B.n497 VSUBS 0.00945f
C538 B.n498 VSUBS 0.00945f
C539 B.n499 VSUBS 0.00945f
C540 B.n500 VSUBS 0.00945f
C541 B.n501 VSUBS 0.00945f
C542 B.n502 VSUBS 0.00945f
C543 B.n503 VSUBS 0.00945f
C544 B.n504 VSUBS 0.00945f
C545 B.n505 VSUBS 0.00945f
C546 B.n506 VSUBS 0.00945f
C547 B.n507 VSUBS 0.00945f
C548 B.n508 VSUBS 0.00945f
C549 B.n509 VSUBS 0.00945f
C550 B.n510 VSUBS 0.00945f
C551 B.n511 VSUBS 0.00945f
C552 B.n512 VSUBS 0.00945f
C553 B.n513 VSUBS 0.00945f
C554 B.n514 VSUBS 0.00945f
C555 B.n515 VSUBS 0.00945f
C556 B.n516 VSUBS 0.00945f
C557 B.n517 VSUBS 0.00945f
C558 B.n518 VSUBS 0.00945f
C559 B.n519 VSUBS 0.00945f
C560 B.n520 VSUBS 0.00945f
C561 B.n521 VSUBS 0.00945f
C562 B.n522 VSUBS 0.00945f
C563 B.n523 VSUBS 0.00945f
C564 B.n524 VSUBS 0.00945f
C565 B.n525 VSUBS 0.00945f
C566 B.n526 VSUBS 0.00945f
C567 B.n527 VSUBS 0.00945f
C568 B.n528 VSUBS 0.00945f
C569 B.n529 VSUBS 0.00945f
C570 B.n530 VSUBS 0.00945f
C571 B.n531 VSUBS 0.00945f
C572 B.n532 VSUBS 0.00945f
C573 B.n533 VSUBS 0.00945f
C574 B.n534 VSUBS 0.00945f
C575 B.n535 VSUBS 0.00945f
C576 B.n536 VSUBS 0.00945f
C577 B.n537 VSUBS 0.00945f
C578 B.n538 VSUBS 0.00945f
C579 B.n539 VSUBS 0.00945f
C580 B.n540 VSUBS 0.00945f
C581 B.n541 VSUBS 0.00945f
C582 B.n542 VSUBS 0.00945f
C583 B.n543 VSUBS 0.00945f
C584 B.n544 VSUBS 0.00945f
C585 B.n545 VSUBS 0.00945f
C586 B.n546 VSUBS 0.00945f
C587 B.n547 VSUBS 0.00945f
C588 B.n548 VSUBS 0.00945f
C589 B.n549 VSUBS 0.00945f
C590 B.n550 VSUBS 0.00945f
C591 B.n551 VSUBS 0.00945f
C592 B.n552 VSUBS 0.00945f
C593 B.n553 VSUBS 0.00945f
C594 B.n554 VSUBS 0.00945f
C595 B.n555 VSUBS 0.00945f
C596 B.n556 VSUBS 0.00945f
C597 B.n557 VSUBS 0.00945f
C598 B.n558 VSUBS 0.00945f
C599 B.n559 VSUBS 0.00945f
C600 B.n560 VSUBS 0.00945f
C601 B.n561 VSUBS 0.00945f
C602 B.n562 VSUBS 0.00945f
C603 B.n563 VSUBS 0.00945f
C604 B.n564 VSUBS 0.00945f
C605 B.n565 VSUBS 0.00945f
C606 B.n566 VSUBS 0.00945f
C607 B.n567 VSUBS 0.00945f
C608 B.n568 VSUBS 0.00945f
C609 B.n569 VSUBS 0.00945f
C610 B.n570 VSUBS 0.00945f
C611 B.n571 VSUBS 0.00945f
C612 B.n572 VSUBS 0.00945f
C613 B.n573 VSUBS 0.00945f
C614 B.n574 VSUBS 0.00945f
C615 B.n575 VSUBS 0.00945f
C616 B.n576 VSUBS 0.00945f
C617 B.n577 VSUBS 0.00945f
C618 B.n578 VSUBS 0.00945f
C619 B.n579 VSUBS 0.00945f
C620 B.n580 VSUBS 0.00945f
C621 B.n581 VSUBS 0.00945f
C622 B.n582 VSUBS 0.00945f
C623 B.n583 VSUBS 0.00945f
C624 B.n584 VSUBS 0.00945f
C625 B.n585 VSUBS 0.00945f
C626 B.n586 VSUBS 0.00945f
C627 B.n587 VSUBS 0.00945f
C628 B.n588 VSUBS 0.00945f
C629 B.n589 VSUBS 0.00945f
C630 B.n590 VSUBS 0.00945f
C631 B.n591 VSUBS 0.00945f
C632 B.n592 VSUBS 0.00945f
C633 B.n593 VSUBS 0.00945f
C634 B.n594 VSUBS 0.00945f
C635 B.n595 VSUBS 0.00945f
C636 B.n596 VSUBS 0.00945f
C637 B.n597 VSUBS 0.00945f
C638 B.n598 VSUBS 0.00945f
C639 B.n599 VSUBS 0.00945f
C640 B.n600 VSUBS 0.00945f
C641 B.n601 VSUBS 0.00945f
C642 B.n602 VSUBS 0.00945f
C643 B.n603 VSUBS 0.00945f
C644 B.n604 VSUBS 0.00945f
C645 B.n605 VSUBS 0.00945f
C646 B.n606 VSUBS 0.00945f
C647 B.n607 VSUBS 0.00945f
C648 B.n608 VSUBS 0.00945f
C649 B.n609 VSUBS 0.00945f
C650 B.n610 VSUBS 0.00945f
C651 B.n611 VSUBS 0.00945f
C652 B.n612 VSUBS 0.00945f
C653 B.n613 VSUBS 0.00945f
C654 B.n614 VSUBS 0.00945f
C655 B.n615 VSUBS 0.00945f
C656 B.n616 VSUBS 0.00945f
C657 B.n617 VSUBS 0.00945f
C658 B.n618 VSUBS 0.00945f
C659 B.n619 VSUBS 0.00945f
C660 B.n620 VSUBS 0.00945f
C661 B.n621 VSUBS 0.00945f
C662 B.n622 VSUBS 0.00945f
C663 B.n623 VSUBS 0.00945f
C664 B.n624 VSUBS 0.00945f
C665 B.n625 VSUBS 0.00945f
C666 B.n626 VSUBS 0.00945f
C667 B.n627 VSUBS 0.00945f
C668 B.n628 VSUBS 0.00945f
C669 B.n629 VSUBS 0.00945f
C670 B.n630 VSUBS 0.00945f
C671 B.n631 VSUBS 0.00945f
C672 B.n632 VSUBS 0.00945f
C673 B.n633 VSUBS 0.00945f
C674 B.n634 VSUBS 0.00945f
C675 B.n635 VSUBS 0.00945f
C676 B.n636 VSUBS 0.00945f
C677 B.n637 VSUBS 0.00945f
C678 B.n638 VSUBS 0.00945f
C679 B.n639 VSUBS 0.00945f
C680 B.n640 VSUBS 0.00945f
C681 B.n641 VSUBS 0.00945f
C682 B.n642 VSUBS 0.00945f
C683 B.n643 VSUBS 0.00945f
C684 B.n644 VSUBS 0.00945f
C685 B.n645 VSUBS 0.00945f
C686 B.n646 VSUBS 0.00945f
C687 B.n647 VSUBS 0.00945f
C688 B.n648 VSUBS 0.00945f
C689 B.n649 VSUBS 0.00945f
C690 B.n650 VSUBS 0.00945f
C691 B.n651 VSUBS 0.00945f
C692 B.n652 VSUBS 0.00945f
C693 B.n653 VSUBS 0.00945f
C694 B.n654 VSUBS 0.00945f
C695 B.n655 VSUBS 0.00945f
C696 B.n656 VSUBS 0.00945f
C697 B.n657 VSUBS 0.00945f
C698 B.n658 VSUBS 0.00945f
C699 B.n659 VSUBS 0.00945f
C700 B.n660 VSUBS 0.00945f
C701 B.n661 VSUBS 0.00945f
C702 B.n662 VSUBS 0.00945f
C703 B.n663 VSUBS 0.00945f
C704 B.n664 VSUBS 0.00945f
C705 B.n665 VSUBS 0.00945f
C706 B.n666 VSUBS 0.00945f
C707 B.n667 VSUBS 0.02266f
C708 B.n668 VSUBS 0.02266f
C709 B.n669 VSUBS 0.023201f
C710 B.n670 VSUBS 0.00945f
C711 B.n671 VSUBS 0.00945f
C712 B.n672 VSUBS 0.00945f
C713 B.n673 VSUBS 0.00945f
C714 B.n674 VSUBS 0.00945f
C715 B.n675 VSUBS 0.00945f
C716 B.n676 VSUBS 0.00945f
C717 B.n677 VSUBS 0.00945f
C718 B.n678 VSUBS 0.00945f
C719 B.n679 VSUBS 0.00945f
C720 B.n680 VSUBS 0.00945f
C721 B.n681 VSUBS 0.00945f
C722 B.n682 VSUBS 0.00945f
C723 B.n683 VSUBS 0.00945f
C724 B.n684 VSUBS 0.00945f
C725 B.n685 VSUBS 0.00945f
C726 B.n686 VSUBS 0.00945f
C727 B.n687 VSUBS 0.00945f
C728 B.n688 VSUBS 0.00945f
C729 B.n689 VSUBS 0.00945f
C730 B.n690 VSUBS 0.00945f
C731 B.n691 VSUBS 0.00945f
C732 B.n692 VSUBS 0.00945f
C733 B.n693 VSUBS 0.00945f
C734 B.n694 VSUBS 0.00945f
C735 B.n695 VSUBS 0.00945f
C736 B.n696 VSUBS 0.00945f
C737 B.n697 VSUBS 0.00945f
C738 B.n698 VSUBS 0.00945f
C739 B.n699 VSUBS 0.00945f
C740 B.n700 VSUBS 0.00945f
C741 B.n701 VSUBS 0.00945f
C742 B.n702 VSUBS 0.00945f
C743 B.n703 VSUBS 0.00945f
C744 B.n704 VSUBS 0.00945f
C745 B.n705 VSUBS 0.00945f
C746 B.n706 VSUBS 0.00945f
C747 B.n707 VSUBS 0.00945f
C748 B.n708 VSUBS 0.00945f
C749 B.n709 VSUBS 0.00945f
C750 B.n710 VSUBS 0.00945f
C751 B.n711 VSUBS 0.00945f
C752 B.n712 VSUBS 0.00945f
C753 B.n713 VSUBS 0.00945f
C754 B.n714 VSUBS 0.00945f
C755 B.n715 VSUBS 0.00945f
C756 B.n716 VSUBS 0.00945f
C757 B.n717 VSUBS 0.00945f
C758 B.n718 VSUBS 0.00945f
C759 B.n719 VSUBS 0.00945f
C760 B.n720 VSUBS 0.00945f
C761 B.n721 VSUBS 0.00945f
C762 B.n722 VSUBS 0.00945f
C763 B.n723 VSUBS 0.00945f
C764 B.n724 VSUBS 0.00945f
C765 B.n725 VSUBS 0.006532f
C766 B.n726 VSUBS 0.021895f
C767 B.n727 VSUBS 0.007644f
C768 B.n728 VSUBS 0.00945f
C769 B.n729 VSUBS 0.00945f
C770 B.n730 VSUBS 0.00945f
C771 B.n731 VSUBS 0.00945f
C772 B.n732 VSUBS 0.00945f
C773 B.n733 VSUBS 0.00945f
C774 B.n734 VSUBS 0.00945f
C775 B.n735 VSUBS 0.00945f
C776 B.n736 VSUBS 0.00945f
C777 B.n737 VSUBS 0.00945f
C778 B.n738 VSUBS 0.00945f
C779 B.n739 VSUBS 0.007644f
C780 B.n740 VSUBS 0.021895f
C781 B.n741 VSUBS 0.006532f
C782 B.n742 VSUBS 0.00945f
C783 B.n743 VSUBS 0.00945f
C784 B.n744 VSUBS 0.00945f
C785 B.n745 VSUBS 0.00945f
C786 B.n746 VSUBS 0.00945f
C787 B.n747 VSUBS 0.00945f
C788 B.n748 VSUBS 0.00945f
C789 B.n749 VSUBS 0.00945f
C790 B.n750 VSUBS 0.00945f
C791 B.n751 VSUBS 0.00945f
C792 B.n752 VSUBS 0.00945f
C793 B.n753 VSUBS 0.00945f
C794 B.n754 VSUBS 0.00945f
C795 B.n755 VSUBS 0.00945f
C796 B.n756 VSUBS 0.00945f
C797 B.n757 VSUBS 0.00945f
C798 B.n758 VSUBS 0.00945f
C799 B.n759 VSUBS 0.00945f
C800 B.n760 VSUBS 0.00945f
C801 B.n761 VSUBS 0.00945f
C802 B.n762 VSUBS 0.00945f
C803 B.n763 VSUBS 0.00945f
C804 B.n764 VSUBS 0.00945f
C805 B.n765 VSUBS 0.00945f
C806 B.n766 VSUBS 0.00945f
C807 B.n767 VSUBS 0.00945f
C808 B.n768 VSUBS 0.00945f
C809 B.n769 VSUBS 0.00945f
C810 B.n770 VSUBS 0.00945f
C811 B.n771 VSUBS 0.00945f
C812 B.n772 VSUBS 0.00945f
C813 B.n773 VSUBS 0.00945f
C814 B.n774 VSUBS 0.00945f
C815 B.n775 VSUBS 0.00945f
C816 B.n776 VSUBS 0.00945f
C817 B.n777 VSUBS 0.00945f
C818 B.n778 VSUBS 0.00945f
C819 B.n779 VSUBS 0.00945f
C820 B.n780 VSUBS 0.00945f
C821 B.n781 VSUBS 0.00945f
C822 B.n782 VSUBS 0.00945f
C823 B.n783 VSUBS 0.00945f
C824 B.n784 VSUBS 0.00945f
C825 B.n785 VSUBS 0.00945f
C826 B.n786 VSUBS 0.00945f
C827 B.n787 VSUBS 0.00945f
C828 B.n788 VSUBS 0.00945f
C829 B.n789 VSUBS 0.00945f
C830 B.n790 VSUBS 0.00945f
C831 B.n791 VSUBS 0.00945f
C832 B.n792 VSUBS 0.00945f
C833 B.n793 VSUBS 0.00945f
C834 B.n794 VSUBS 0.00945f
C835 B.n795 VSUBS 0.00945f
C836 B.n796 VSUBS 0.00945f
C837 B.n797 VSUBS 0.023201f
C838 B.n798 VSUBS 0.02266f
C839 B.n799 VSUBS 0.02266f
C840 B.n800 VSUBS 0.00945f
C841 B.n801 VSUBS 0.00945f
C842 B.n802 VSUBS 0.00945f
C843 B.n803 VSUBS 0.00945f
C844 B.n804 VSUBS 0.00945f
C845 B.n805 VSUBS 0.00945f
C846 B.n806 VSUBS 0.00945f
C847 B.n807 VSUBS 0.00945f
C848 B.n808 VSUBS 0.00945f
C849 B.n809 VSUBS 0.00945f
C850 B.n810 VSUBS 0.00945f
C851 B.n811 VSUBS 0.00945f
C852 B.n812 VSUBS 0.00945f
C853 B.n813 VSUBS 0.00945f
C854 B.n814 VSUBS 0.00945f
C855 B.n815 VSUBS 0.00945f
C856 B.n816 VSUBS 0.00945f
C857 B.n817 VSUBS 0.00945f
C858 B.n818 VSUBS 0.00945f
C859 B.n819 VSUBS 0.00945f
C860 B.n820 VSUBS 0.00945f
C861 B.n821 VSUBS 0.00945f
C862 B.n822 VSUBS 0.00945f
C863 B.n823 VSUBS 0.00945f
C864 B.n824 VSUBS 0.00945f
C865 B.n825 VSUBS 0.00945f
C866 B.n826 VSUBS 0.00945f
C867 B.n827 VSUBS 0.00945f
C868 B.n828 VSUBS 0.00945f
C869 B.n829 VSUBS 0.00945f
C870 B.n830 VSUBS 0.00945f
C871 B.n831 VSUBS 0.00945f
C872 B.n832 VSUBS 0.00945f
C873 B.n833 VSUBS 0.00945f
C874 B.n834 VSUBS 0.00945f
C875 B.n835 VSUBS 0.00945f
C876 B.n836 VSUBS 0.00945f
C877 B.n837 VSUBS 0.00945f
C878 B.n838 VSUBS 0.00945f
C879 B.n839 VSUBS 0.00945f
C880 B.n840 VSUBS 0.00945f
C881 B.n841 VSUBS 0.00945f
C882 B.n842 VSUBS 0.00945f
C883 B.n843 VSUBS 0.00945f
C884 B.n844 VSUBS 0.00945f
C885 B.n845 VSUBS 0.00945f
C886 B.n846 VSUBS 0.00945f
C887 B.n847 VSUBS 0.00945f
C888 B.n848 VSUBS 0.00945f
C889 B.n849 VSUBS 0.00945f
C890 B.n850 VSUBS 0.00945f
C891 B.n851 VSUBS 0.00945f
C892 B.n852 VSUBS 0.00945f
C893 B.n853 VSUBS 0.00945f
C894 B.n854 VSUBS 0.00945f
C895 B.n855 VSUBS 0.00945f
C896 B.n856 VSUBS 0.00945f
C897 B.n857 VSUBS 0.00945f
C898 B.n858 VSUBS 0.00945f
C899 B.n859 VSUBS 0.00945f
C900 B.n860 VSUBS 0.00945f
C901 B.n861 VSUBS 0.00945f
C902 B.n862 VSUBS 0.00945f
C903 B.n863 VSUBS 0.00945f
C904 B.n864 VSUBS 0.00945f
C905 B.n865 VSUBS 0.00945f
C906 B.n866 VSUBS 0.00945f
C907 B.n867 VSUBS 0.00945f
C908 B.n868 VSUBS 0.00945f
C909 B.n869 VSUBS 0.00945f
C910 B.n870 VSUBS 0.00945f
C911 B.n871 VSUBS 0.00945f
C912 B.n872 VSUBS 0.00945f
C913 B.n873 VSUBS 0.00945f
C914 B.n874 VSUBS 0.00945f
C915 B.n875 VSUBS 0.00945f
C916 B.n876 VSUBS 0.00945f
C917 B.n877 VSUBS 0.00945f
C918 B.n878 VSUBS 0.00945f
C919 B.n879 VSUBS 0.00945f
C920 B.n880 VSUBS 0.00945f
C921 B.n881 VSUBS 0.00945f
C922 B.n882 VSUBS 0.00945f
C923 B.n883 VSUBS 0.00945f
C924 B.n884 VSUBS 0.00945f
C925 B.n885 VSUBS 0.00945f
C926 B.n886 VSUBS 0.00945f
C927 B.n887 VSUBS 0.00945f
C928 B.n888 VSUBS 0.00945f
C929 B.n889 VSUBS 0.00945f
C930 B.n890 VSUBS 0.00945f
C931 B.n891 VSUBS 0.00945f
C932 B.n892 VSUBS 0.00945f
C933 B.n893 VSUBS 0.00945f
C934 B.n894 VSUBS 0.00945f
C935 B.n895 VSUBS 0.00945f
C936 B.n896 VSUBS 0.00945f
C937 B.n897 VSUBS 0.00945f
C938 B.n898 VSUBS 0.00945f
C939 B.n899 VSUBS 0.012332f
C940 B.n900 VSUBS 0.013137f
C941 B.n901 VSUBS 0.026124f
C942 VDD1.n0 VSUBS 0.033951f
C943 VDD1.n1 VSUBS 0.031137f
C944 VDD1.n2 VSUBS 0.016732f
C945 VDD1.n3 VSUBS 0.039548f
C946 VDD1.n4 VSUBS 0.017716f
C947 VDD1.n5 VSUBS 0.031137f
C948 VDD1.n6 VSUBS 0.016732f
C949 VDD1.n7 VSUBS 0.039548f
C950 VDD1.n8 VSUBS 0.017716f
C951 VDD1.n9 VSUBS 0.031137f
C952 VDD1.n10 VSUBS 0.016732f
C953 VDD1.n11 VSUBS 0.039548f
C954 VDD1.n12 VSUBS 0.039548f
C955 VDD1.n13 VSUBS 0.017716f
C956 VDD1.n14 VSUBS 0.031137f
C957 VDD1.n15 VSUBS 0.016732f
C958 VDD1.n16 VSUBS 0.039548f
C959 VDD1.n17 VSUBS 0.017716f
C960 VDD1.n18 VSUBS 0.227636f
C961 VDD1.t3 VSUBS 0.085103f
C962 VDD1.n19 VSUBS 0.029661f
C963 VDD1.n20 VSUBS 0.02975f
C964 VDD1.n21 VSUBS 0.016732f
C965 VDD1.n22 VSUBS 1.3593f
C966 VDD1.n23 VSUBS 0.031137f
C967 VDD1.n24 VSUBS 0.016732f
C968 VDD1.n25 VSUBS 0.017716f
C969 VDD1.n26 VSUBS 0.039548f
C970 VDD1.n27 VSUBS 0.039548f
C971 VDD1.n28 VSUBS 0.017716f
C972 VDD1.n29 VSUBS 0.016732f
C973 VDD1.n30 VSUBS 0.031137f
C974 VDD1.n31 VSUBS 0.031137f
C975 VDD1.n32 VSUBS 0.016732f
C976 VDD1.n33 VSUBS 0.017716f
C977 VDD1.n34 VSUBS 0.039548f
C978 VDD1.n35 VSUBS 0.039548f
C979 VDD1.n36 VSUBS 0.017716f
C980 VDD1.n37 VSUBS 0.016732f
C981 VDD1.n38 VSUBS 0.031137f
C982 VDD1.n39 VSUBS 0.031137f
C983 VDD1.n40 VSUBS 0.016732f
C984 VDD1.n41 VSUBS 0.017224f
C985 VDD1.n42 VSUBS 0.017224f
C986 VDD1.n43 VSUBS 0.039548f
C987 VDD1.n44 VSUBS 0.039548f
C988 VDD1.n45 VSUBS 0.017716f
C989 VDD1.n46 VSUBS 0.016732f
C990 VDD1.n47 VSUBS 0.031137f
C991 VDD1.n48 VSUBS 0.031137f
C992 VDD1.n49 VSUBS 0.016732f
C993 VDD1.n50 VSUBS 0.017716f
C994 VDD1.n51 VSUBS 0.039548f
C995 VDD1.n52 VSUBS 0.094848f
C996 VDD1.n53 VSUBS 0.017716f
C997 VDD1.n54 VSUBS 0.016732f
C998 VDD1.n55 VSUBS 0.074949f
C999 VDD1.n56 VSUBS 0.089047f
C1000 VDD1.t4 VSUBS 0.264509f
C1001 VDD1.t6 VSUBS 0.264509f
C1002 VDD1.n57 VSUBS 2.02937f
C1003 VDD1.n58 VSUBS 1.27994f
C1004 VDD1.n59 VSUBS 0.033951f
C1005 VDD1.n60 VSUBS 0.031137f
C1006 VDD1.n61 VSUBS 0.016732f
C1007 VDD1.n62 VSUBS 0.039548f
C1008 VDD1.n63 VSUBS 0.017716f
C1009 VDD1.n64 VSUBS 0.031137f
C1010 VDD1.n65 VSUBS 0.016732f
C1011 VDD1.n66 VSUBS 0.039548f
C1012 VDD1.n67 VSUBS 0.017716f
C1013 VDD1.n68 VSUBS 0.031137f
C1014 VDD1.n69 VSUBS 0.016732f
C1015 VDD1.n70 VSUBS 0.039548f
C1016 VDD1.n71 VSUBS 0.017716f
C1017 VDD1.n72 VSUBS 0.031137f
C1018 VDD1.n73 VSUBS 0.016732f
C1019 VDD1.n74 VSUBS 0.039548f
C1020 VDD1.n75 VSUBS 0.017716f
C1021 VDD1.n76 VSUBS 0.227636f
C1022 VDD1.t7 VSUBS 0.085103f
C1023 VDD1.n77 VSUBS 0.029661f
C1024 VDD1.n78 VSUBS 0.02975f
C1025 VDD1.n79 VSUBS 0.016732f
C1026 VDD1.n80 VSUBS 1.3593f
C1027 VDD1.n81 VSUBS 0.031137f
C1028 VDD1.n82 VSUBS 0.016732f
C1029 VDD1.n83 VSUBS 0.017716f
C1030 VDD1.n84 VSUBS 0.039548f
C1031 VDD1.n85 VSUBS 0.039548f
C1032 VDD1.n86 VSUBS 0.017716f
C1033 VDD1.n87 VSUBS 0.016732f
C1034 VDD1.n88 VSUBS 0.031137f
C1035 VDD1.n89 VSUBS 0.031137f
C1036 VDD1.n90 VSUBS 0.016732f
C1037 VDD1.n91 VSUBS 0.017716f
C1038 VDD1.n92 VSUBS 0.039548f
C1039 VDD1.n93 VSUBS 0.039548f
C1040 VDD1.n94 VSUBS 0.039548f
C1041 VDD1.n95 VSUBS 0.017716f
C1042 VDD1.n96 VSUBS 0.016732f
C1043 VDD1.n97 VSUBS 0.031137f
C1044 VDD1.n98 VSUBS 0.031137f
C1045 VDD1.n99 VSUBS 0.016732f
C1046 VDD1.n100 VSUBS 0.017224f
C1047 VDD1.n101 VSUBS 0.017224f
C1048 VDD1.n102 VSUBS 0.039548f
C1049 VDD1.n103 VSUBS 0.039548f
C1050 VDD1.n104 VSUBS 0.017716f
C1051 VDD1.n105 VSUBS 0.016732f
C1052 VDD1.n106 VSUBS 0.031137f
C1053 VDD1.n107 VSUBS 0.031137f
C1054 VDD1.n108 VSUBS 0.016732f
C1055 VDD1.n109 VSUBS 0.017716f
C1056 VDD1.n110 VSUBS 0.039548f
C1057 VDD1.n111 VSUBS 0.094848f
C1058 VDD1.n112 VSUBS 0.017716f
C1059 VDD1.n113 VSUBS 0.016732f
C1060 VDD1.n114 VSUBS 0.074949f
C1061 VDD1.n115 VSUBS 0.089047f
C1062 VDD1.t0 VSUBS 0.264509f
C1063 VDD1.t2 VSUBS 0.264509f
C1064 VDD1.n116 VSUBS 2.02936f
C1065 VDD1.n117 VSUBS 1.26962f
C1066 VDD1.t8 VSUBS 0.264509f
C1067 VDD1.t1 VSUBS 0.264509f
C1068 VDD1.n118 VSUBS 2.05901f
C1069 VDD1.n119 VSUBS 4.31828f
C1070 VDD1.t5 VSUBS 0.264509f
C1071 VDD1.t9 VSUBS 0.264509f
C1072 VDD1.n120 VSUBS 2.02936f
C1073 VDD1.n121 VSUBS 4.39686f
C1074 VP.t8 VSUBS 2.62427f
C1075 VP.n0 VSUBS 1.04094f
C1076 VP.n1 VSUBS 0.029093f
C1077 VP.n2 VSUBS 0.030513f
C1078 VP.n3 VSUBS 0.029093f
C1079 VP.t1 VSUBS 2.62427f
C1080 VP.n4 VSUBS 0.929519f
C1081 VP.n5 VSUBS 0.029093f
C1082 VP.n6 VSUBS 0.039227f
C1083 VP.n7 VSUBS 0.029093f
C1084 VP.t7 VSUBS 2.62427f
C1085 VP.n8 VSUBS 0.054221f
C1086 VP.n9 VSUBS 0.029093f
C1087 VP.n10 VSUBS 0.054221f
C1088 VP.n11 VSUBS 0.029093f
C1089 VP.t9 VSUBS 2.62427f
C1090 VP.n12 VSUBS 0.057028f
C1091 VP.n13 VSUBS 0.029093f
C1092 VP.n14 VSUBS 0.045655f
C1093 VP.t0 VSUBS 2.62427f
C1094 VP.n15 VSUBS 1.04094f
C1095 VP.n16 VSUBS 0.029093f
C1096 VP.n17 VSUBS 0.030513f
C1097 VP.n18 VSUBS 0.029093f
C1098 VP.t4 VSUBS 2.62427f
C1099 VP.n19 VSUBS 0.929519f
C1100 VP.n20 VSUBS 0.029093f
C1101 VP.n21 VSUBS 0.039227f
C1102 VP.n22 VSUBS 0.029093f
C1103 VP.t3 VSUBS 2.62427f
C1104 VP.n23 VSUBS 0.054221f
C1105 VP.n24 VSUBS 0.029093f
C1106 VP.n25 VSUBS 0.054221f
C1107 VP.t6 VSUBS 2.94551f
C1108 VP.n26 VSUBS 0.979989f
C1109 VP.t5 VSUBS 2.62427f
C1110 VP.n27 VSUBS 1.03313f
C1111 VP.n28 VSUBS 0.049938f
C1112 VP.n29 VSUBS 0.333455f
C1113 VP.n30 VSUBS 0.029093f
C1114 VP.n31 VSUBS 0.029093f
C1115 VP.n32 VSUBS 0.045713f
C1116 VP.n33 VSUBS 0.039227f
C1117 VP.n34 VSUBS 0.054221f
C1118 VP.n35 VSUBS 0.029093f
C1119 VP.n36 VSUBS 0.029093f
C1120 VP.n37 VSUBS 0.029093f
C1121 VP.n38 VSUBS 0.956971f
C1122 VP.n39 VSUBS 0.054221f
C1123 VP.n40 VSUBS 0.054221f
C1124 VP.n41 VSUBS 0.029093f
C1125 VP.n42 VSUBS 0.029093f
C1126 VP.n43 VSUBS 0.029093f
C1127 VP.n44 VSUBS 0.045713f
C1128 VP.n45 VSUBS 0.054221f
C1129 VP.n46 VSUBS 0.049938f
C1130 VP.n47 VSUBS 0.029093f
C1131 VP.n48 VSUBS 0.029093f
C1132 VP.n49 VSUBS 0.031735f
C1133 VP.n50 VSUBS 0.054221f
C1134 VP.n51 VSUBS 0.057028f
C1135 VP.n52 VSUBS 0.029093f
C1136 VP.n53 VSUBS 0.029093f
C1137 VP.n54 VSUBS 0.029093f
C1138 VP.n55 VSUBS 0.05162f
C1139 VP.n56 VSUBS 0.054221f
C1140 VP.n57 VSUBS 0.045655f
C1141 VP.n58 VSUBS 0.046955f
C1142 VP.n59 VSUBS 1.88317f
C1143 VP.t2 VSUBS 2.62427f
C1144 VP.n60 VSUBS 1.04094f
C1145 VP.n61 VSUBS 1.90222f
C1146 VP.n62 VSUBS 0.046955f
C1147 VP.n63 VSUBS 0.029093f
C1148 VP.n64 VSUBS 0.054221f
C1149 VP.n65 VSUBS 0.05162f
C1150 VP.n66 VSUBS 0.030513f
C1151 VP.n67 VSUBS 0.029093f
C1152 VP.n68 VSUBS 0.029093f
C1153 VP.n69 VSUBS 0.029093f
C1154 VP.n70 VSUBS 0.054221f
C1155 VP.n71 VSUBS 0.031735f
C1156 VP.n72 VSUBS 0.929519f
C1157 VP.n73 VSUBS 0.049938f
C1158 VP.n74 VSUBS 0.029093f
C1159 VP.n75 VSUBS 0.029093f
C1160 VP.n76 VSUBS 0.029093f
C1161 VP.n77 VSUBS 0.045713f
C1162 VP.n78 VSUBS 0.039227f
C1163 VP.n79 VSUBS 0.054221f
C1164 VP.n80 VSUBS 0.029093f
C1165 VP.n81 VSUBS 0.029093f
C1166 VP.n82 VSUBS 0.029093f
C1167 VP.n83 VSUBS 0.956971f
C1168 VP.n84 VSUBS 0.054221f
C1169 VP.n85 VSUBS 0.054221f
C1170 VP.n86 VSUBS 0.029093f
C1171 VP.n87 VSUBS 0.029093f
C1172 VP.n88 VSUBS 0.029093f
C1173 VP.n89 VSUBS 0.045713f
C1174 VP.n90 VSUBS 0.054221f
C1175 VP.n91 VSUBS 0.049938f
C1176 VP.n92 VSUBS 0.029093f
C1177 VP.n93 VSUBS 0.029093f
C1178 VP.n94 VSUBS 0.031735f
C1179 VP.n95 VSUBS 0.054221f
C1180 VP.n96 VSUBS 0.057028f
C1181 VP.n97 VSUBS 0.029093f
C1182 VP.n98 VSUBS 0.029093f
C1183 VP.n99 VSUBS 0.029093f
C1184 VP.n100 VSUBS 0.05162f
C1185 VP.n101 VSUBS 0.054221f
C1186 VP.n102 VSUBS 0.045655f
C1187 VP.n103 VSUBS 0.046955f
C1188 VP.n104 VSUBS 0.065674f
C1189 VTAIL.t9 VSUBS 0.253703f
C1190 VTAIL.t17 VSUBS 0.253703f
C1191 VTAIL.n0 VSUBS 1.79828f
C1192 VTAIL.n1 VSUBS 1.0566f
C1193 VTAIL.n2 VSUBS 0.032564f
C1194 VTAIL.n3 VSUBS 0.029865f
C1195 VTAIL.n4 VSUBS 0.016048f
C1196 VTAIL.n5 VSUBS 0.037932f
C1197 VTAIL.n6 VSUBS 0.016992f
C1198 VTAIL.n7 VSUBS 0.029865f
C1199 VTAIL.n8 VSUBS 0.016048f
C1200 VTAIL.n9 VSUBS 0.037932f
C1201 VTAIL.n10 VSUBS 0.016992f
C1202 VTAIL.n11 VSUBS 0.029865f
C1203 VTAIL.n12 VSUBS 0.016048f
C1204 VTAIL.n13 VSUBS 0.037932f
C1205 VTAIL.n14 VSUBS 0.016992f
C1206 VTAIL.n15 VSUBS 0.029865f
C1207 VTAIL.n16 VSUBS 0.016048f
C1208 VTAIL.n17 VSUBS 0.037932f
C1209 VTAIL.n18 VSUBS 0.016992f
C1210 VTAIL.n19 VSUBS 0.218336f
C1211 VTAIL.t19 VSUBS 0.081626f
C1212 VTAIL.n20 VSUBS 0.028449f
C1213 VTAIL.n21 VSUBS 0.028534f
C1214 VTAIL.n22 VSUBS 0.016048f
C1215 VTAIL.n23 VSUBS 1.30377f
C1216 VTAIL.n24 VSUBS 0.029865f
C1217 VTAIL.n25 VSUBS 0.016048f
C1218 VTAIL.n26 VSUBS 0.016992f
C1219 VTAIL.n27 VSUBS 0.037932f
C1220 VTAIL.n28 VSUBS 0.037932f
C1221 VTAIL.n29 VSUBS 0.016992f
C1222 VTAIL.n30 VSUBS 0.016048f
C1223 VTAIL.n31 VSUBS 0.029865f
C1224 VTAIL.n32 VSUBS 0.029865f
C1225 VTAIL.n33 VSUBS 0.016048f
C1226 VTAIL.n34 VSUBS 0.016992f
C1227 VTAIL.n35 VSUBS 0.037932f
C1228 VTAIL.n36 VSUBS 0.037932f
C1229 VTAIL.n37 VSUBS 0.037932f
C1230 VTAIL.n38 VSUBS 0.016992f
C1231 VTAIL.n39 VSUBS 0.016048f
C1232 VTAIL.n40 VSUBS 0.029865f
C1233 VTAIL.n41 VSUBS 0.029865f
C1234 VTAIL.n42 VSUBS 0.016048f
C1235 VTAIL.n43 VSUBS 0.01652f
C1236 VTAIL.n44 VSUBS 0.01652f
C1237 VTAIL.n45 VSUBS 0.037932f
C1238 VTAIL.n46 VSUBS 0.037932f
C1239 VTAIL.n47 VSUBS 0.016992f
C1240 VTAIL.n48 VSUBS 0.016048f
C1241 VTAIL.n49 VSUBS 0.029865f
C1242 VTAIL.n50 VSUBS 0.029865f
C1243 VTAIL.n51 VSUBS 0.016048f
C1244 VTAIL.n52 VSUBS 0.016992f
C1245 VTAIL.n53 VSUBS 0.037932f
C1246 VTAIL.n54 VSUBS 0.090973f
C1247 VTAIL.n55 VSUBS 0.016992f
C1248 VTAIL.n56 VSUBS 0.016048f
C1249 VTAIL.n57 VSUBS 0.071887f
C1250 VTAIL.n58 VSUBS 0.045798f
C1251 VTAIL.n59 VSUBS 0.49791f
C1252 VTAIL.t6 VSUBS 0.253703f
C1253 VTAIL.t2 VSUBS 0.253703f
C1254 VTAIL.n60 VSUBS 1.79828f
C1255 VTAIL.n61 VSUBS 1.21858f
C1256 VTAIL.t4 VSUBS 0.253703f
C1257 VTAIL.t1 VSUBS 0.253703f
C1258 VTAIL.n62 VSUBS 1.79828f
C1259 VTAIL.n63 VSUBS 2.79978f
C1260 VTAIL.t13 VSUBS 0.253703f
C1261 VTAIL.t16 VSUBS 0.253703f
C1262 VTAIL.n64 VSUBS 1.79829f
C1263 VTAIL.n65 VSUBS 2.79977f
C1264 VTAIL.t11 VSUBS 0.253703f
C1265 VTAIL.t12 VSUBS 0.253703f
C1266 VTAIL.n66 VSUBS 1.79829f
C1267 VTAIL.n67 VSUBS 1.21857f
C1268 VTAIL.n68 VSUBS 0.032564f
C1269 VTAIL.n69 VSUBS 0.029865f
C1270 VTAIL.n70 VSUBS 0.016048f
C1271 VTAIL.n71 VSUBS 0.037932f
C1272 VTAIL.n72 VSUBS 0.016992f
C1273 VTAIL.n73 VSUBS 0.029865f
C1274 VTAIL.n74 VSUBS 0.016048f
C1275 VTAIL.n75 VSUBS 0.037932f
C1276 VTAIL.n76 VSUBS 0.016992f
C1277 VTAIL.n77 VSUBS 0.029865f
C1278 VTAIL.n78 VSUBS 0.016048f
C1279 VTAIL.n79 VSUBS 0.037932f
C1280 VTAIL.n80 VSUBS 0.037932f
C1281 VTAIL.n81 VSUBS 0.016992f
C1282 VTAIL.n82 VSUBS 0.029865f
C1283 VTAIL.n83 VSUBS 0.016048f
C1284 VTAIL.n84 VSUBS 0.037932f
C1285 VTAIL.n85 VSUBS 0.016992f
C1286 VTAIL.n86 VSUBS 0.218336f
C1287 VTAIL.t15 VSUBS 0.081626f
C1288 VTAIL.n87 VSUBS 0.028449f
C1289 VTAIL.n88 VSUBS 0.028534f
C1290 VTAIL.n89 VSUBS 0.016048f
C1291 VTAIL.n90 VSUBS 1.30377f
C1292 VTAIL.n91 VSUBS 0.029865f
C1293 VTAIL.n92 VSUBS 0.016048f
C1294 VTAIL.n93 VSUBS 0.016992f
C1295 VTAIL.n94 VSUBS 0.037932f
C1296 VTAIL.n95 VSUBS 0.037932f
C1297 VTAIL.n96 VSUBS 0.016992f
C1298 VTAIL.n97 VSUBS 0.016048f
C1299 VTAIL.n98 VSUBS 0.029865f
C1300 VTAIL.n99 VSUBS 0.029865f
C1301 VTAIL.n100 VSUBS 0.016048f
C1302 VTAIL.n101 VSUBS 0.016992f
C1303 VTAIL.n102 VSUBS 0.037932f
C1304 VTAIL.n103 VSUBS 0.037932f
C1305 VTAIL.n104 VSUBS 0.016992f
C1306 VTAIL.n105 VSUBS 0.016048f
C1307 VTAIL.n106 VSUBS 0.029865f
C1308 VTAIL.n107 VSUBS 0.029865f
C1309 VTAIL.n108 VSUBS 0.016048f
C1310 VTAIL.n109 VSUBS 0.01652f
C1311 VTAIL.n110 VSUBS 0.01652f
C1312 VTAIL.n111 VSUBS 0.037932f
C1313 VTAIL.n112 VSUBS 0.037932f
C1314 VTAIL.n113 VSUBS 0.016992f
C1315 VTAIL.n114 VSUBS 0.016048f
C1316 VTAIL.n115 VSUBS 0.029865f
C1317 VTAIL.n116 VSUBS 0.029865f
C1318 VTAIL.n117 VSUBS 0.016048f
C1319 VTAIL.n118 VSUBS 0.016992f
C1320 VTAIL.n119 VSUBS 0.037932f
C1321 VTAIL.n120 VSUBS 0.090973f
C1322 VTAIL.n121 VSUBS 0.016992f
C1323 VTAIL.n122 VSUBS 0.016048f
C1324 VTAIL.n123 VSUBS 0.071887f
C1325 VTAIL.n124 VSUBS 0.045798f
C1326 VTAIL.n125 VSUBS 0.49791f
C1327 VTAIL.t3 VSUBS 0.253703f
C1328 VTAIL.t5 VSUBS 0.253703f
C1329 VTAIL.n126 VSUBS 1.79829f
C1330 VTAIL.n127 VSUBS 1.12192f
C1331 VTAIL.t0 VSUBS 0.253703f
C1332 VTAIL.t8 VSUBS 0.253703f
C1333 VTAIL.n128 VSUBS 1.79829f
C1334 VTAIL.n129 VSUBS 1.21857f
C1335 VTAIL.n130 VSUBS 0.032564f
C1336 VTAIL.n131 VSUBS 0.029865f
C1337 VTAIL.n132 VSUBS 0.016048f
C1338 VTAIL.n133 VSUBS 0.037932f
C1339 VTAIL.n134 VSUBS 0.016992f
C1340 VTAIL.n135 VSUBS 0.029865f
C1341 VTAIL.n136 VSUBS 0.016048f
C1342 VTAIL.n137 VSUBS 0.037932f
C1343 VTAIL.n138 VSUBS 0.016992f
C1344 VTAIL.n139 VSUBS 0.029865f
C1345 VTAIL.n140 VSUBS 0.016048f
C1346 VTAIL.n141 VSUBS 0.037932f
C1347 VTAIL.n142 VSUBS 0.037932f
C1348 VTAIL.n143 VSUBS 0.016992f
C1349 VTAIL.n144 VSUBS 0.029865f
C1350 VTAIL.n145 VSUBS 0.016048f
C1351 VTAIL.n146 VSUBS 0.037932f
C1352 VTAIL.n147 VSUBS 0.016992f
C1353 VTAIL.n148 VSUBS 0.218336f
C1354 VTAIL.t7 VSUBS 0.081626f
C1355 VTAIL.n149 VSUBS 0.028449f
C1356 VTAIL.n150 VSUBS 0.028534f
C1357 VTAIL.n151 VSUBS 0.016048f
C1358 VTAIL.n152 VSUBS 1.30377f
C1359 VTAIL.n153 VSUBS 0.029865f
C1360 VTAIL.n154 VSUBS 0.016048f
C1361 VTAIL.n155 VSUBS 0.016992f
C1362 VTAIL.n156 VSUBS 0.037932f
C1363 VTAIL.n157 VSUBS 0.037932f
C1364 VTAIL.n158 VSUBS 0.016992f
C1365 VTAIL.n159 VSUBS 0.016048f
C1366 VTAIL.n160 VSUBS 0.029865f
C1367 VTAIL.n161 VSUBS 0.029865f
C1368 VTAIL.n162 VSUBS 0.016048f
C1369 VTAIL.n163 VSUBS 0.016992f
C1370 VTAIL.n164 VSUBS 0.037932f
C1371 VTAIL.n165 VSUBS 0.037932f
C1372 VTAIL.n166 VSUBS 0.016992f
C1373 VTAIL.n167 VSUBS 0.016048f
C1374 VTAIL.n168 VSUBS 0.029865f
C1375 VTAIL.n169 VSUBS 0.029865f
C1376 VTAIL.n170 VSUBS 0.016048f
C1377 VTAIL.n171 VSUBS 0.01652f
C1378 VTAIL.n172 VSUBS 0.01652f
C1379 VTAIL.n173 VSUBS 0.037932f
C1380 VTAIL.n174 VSUBS 0.037932f
C1381 VTAIL.n175 VSUBS 0.016992f
C1382 VTAIL.n176 VSUBS 0.016048f
C1383 VTAIL.n177 VSUBS 0.029865f
C1384 VTAIL.n178 VSUBS 0.029865f
C1385 VTAIL.n179 VSUBS 0.016048f
C1386 VTAIL.n180 VSUBS 0.016992f
C1387 VTAIL.n181 VSUBS 0.037932f
C1388 VTAIL.n182 VSUBS 0.090973f
C1389 VTAIL.n183 VSUBS 0.016992f
C1390 VTAIL.n184 VSUBS 0.016048f
C1391 VTAIL.n185 VSUBS 0.071887f
C1392 VTAIL.n186 VSUBS 0.045798f
C1393 VTAIL.n187 VSUBS 1.89204f
C1394 VTAIL.n188 VSUBS 0.032564f
C1395 VTAIL.n189 VSUBS 0.029865f
C1396 VTAIL.n190 VSUBS 0.016048f
C1397 VTAIL.n191 VSUBS 0.037932f
C1398 VTAIL.n192 VSUBS 0.016992f
C1399 VTAIL.n193 VSUBS 0.029865f
C1400 VTAIL.n194 VSUBS 0.016048f
C1401 VTAIL.n195 VSUBS 0.037932f
C1402 VTAIL.n196 VSUBS 0.016992f
C1403 VTAIL.n197 VSUBS 0.029865f
C1404 VTAIL.n198 VSUBS 0.016048f
C1405 VTAIL.n199 VSUBS 0.037932f
C1406 VTAIL.n200 VSUBS 0.016992f
C1407 VTAIL.n201 VSUBS 0.029865f
C1408 VTAIL.n202 VSUBS 0.016048f
C1409 VTAIL.n203 VSUBS 0.037932f
C1410 VTAIL.n204 VSUBS 0.016992f
C1411 VTAIL.n205 VSUBS 0.218336f
C1412 VTAIL.t14 VSUBS 0.081626f
C1413 VTAIL.n206 VSUBS 0.028449f
C1414 VTAIL.n207 VSUBS 0.028534f
C1415 VTAIL.n208 VSUBS 0.016048f
C1416 VTAIL.n209 VSUBS 1.30377f
C1417 VTAIL.n210 VSUBS 0.029865f
C1418 VTAIL.n211 VSUBS 0.016048f
C1419 VTAIL.n212 VSUBS 0.016992f
C1420 VTAIL.n213 VSUBS 0.037932f
C1421 VTAIL.n214 VSUBS 0.037932f
C1422 VTAIL.n215 VSUBS 0.016992f
C1423 VTAIL.n216 VSUBS 0.016048f
C1424 VTAIL.n217 VSUBS 0.029865f
C1425 VTAIL.n218 VSUBS 0.029865f
C1426 VTAIL.n219 VSUBS 0.016048f
C1427 VTAIL.n220 VSUBS 0.016992f
C1428 VTAIL.n221 VSUBS 0.037932f
C1429 VTAIL.n222 VSUBS 0.037932f
C1430 VTAIL.n223 VSUBS 0.037932f
C1431 VTAIL.n224 VSUBS 0.016992f
C1432 VTAIL.n225 VSUBS 0.016048f
C1433 VTAIL.n226 VSUBS 0.029865f
C1434 VTAIL.n227 VSUBS 0.029865f
C1435 VTAIL.n228 VSUBS 0.016048f
C1436 VTAIL.n229 VSUBS 0.01652f
C1437 VTAIL.n230 VSUBS 0.01652f
C1438 VTAIL.n231 VSUBS 0.037932f
C1439 VTAIL.n232 VSUBS 0.037932f
C1440 VTAIL.n233 VSUBS 0.016992f
C1441 VTAIL.n234 VSUBS 0.016048f
C1442 VTAIL.n235 VSUBS 0.029865f
C1443 VTAIL.n236 VSUBS 0.029865f
C1444 VTAIL.n237 VSUBS 0.016048f
C1445 VTAIL.n238 VSUBS 0.016992f
C1446 VTAIL.n239 VSUBS 0.037932f
C1447 VTAIL.n240 VSUBS 0.090973f
C1448 VTAIL.n241 VSUBS 0.016992f
C1449 VTAIL.n242 VSUBS 0.016048f
C1450 VTAIL.n243 VSUBS 0.071887f
C1451 VTAIL.n244 VSUBS 0.045798f
C1452 VTAIL.n245 VSUBS 1.89204f
C1453 VTAIL.t10 VSUBS 0.253703f
C1454 VTAIL.t18 VSUBS 0.253703f
C1455 VTAIL.n246 VSUBS 1.79828f
C1456 VTAIL.n247 VSUBS 1.00019f
C1457 VDD2.n0 VSUBS 0.033969f
C1458 VDD2.n1 VSUBS 0.031154f
C1459 VDD2.n2 VSUBS 0.016741f
C1460 VDD2.n3 VSUBS 0.039569f
C1461 VDD2.n4 VSUBS 0.017725f
C1462 VDD2.n5 VSUBS 0.031154f
C1463 VDD2.n6 VSUBS 0.016741f
C1464 VDD2.n7 VSUBS 0.039569f
C1465 VDD2.n8 VSUBS 0.017725f
C1466 VDD2.n9 VSUBS 0.031154f
C1467 VDD2.n10 VSUBS 0.016741f
C1468 VDD2.n11 VSUBS 0.039569f
C1469 VDD2.n12 VSUBS 0.017725f
C1470 VDD2.n13 VSUBS 0.031154f
C1471 VDD2.n14 VSUBS 0.016741f
C1472 VDD2.n15 VSUBS 0.039569f
C1473 VDD2.n16 VSUBS 0.017725f
C1474 VDD2.n17 VSUBS 0.227757f
C1475 VDD2.t5 VSUBS 0.085148f
C1476 VDD2.n18 VSUBS 0.029677f
C1477 VDD2.n19 VSUBS 0.029766f
C1478 VDD2.n20 VSUBS 0.016741f
C1479 VDD2.n21 VSUBS 1.36002f
C1480 VDD2.n22 VSUBS 0.031154f
C1481 VDD2.n23 VSUBS 0.016741f
C1482 VDD2.n24 VSUBS 0.017725f
C1483 VDD2.n25 VSUBS 0.039569f
C1484 VDD2.n26 VSUBS 0.039569f
C1485 VDD2.n27 VSUBS 0.017725f
C1486 VDD2.n28 VSUBS 0.016741f
C1487 VDD2.n29 VSUBS 0.031154f
C1488 VDD2.n30 VSUBS 0.031154f
C1489 VDD2.n31 VSUBS 0.016741f
C1490 VDD2.n32 VSUBS 0.017725f
C1491 VDD2.n33 VSUBS 0.039569f
C1492 VDD2.n34 VSUBS 0.039569f
C1493 VDD2.n35 VSUBS 0.039569f
C1494 VDD2.n36 VSUBS 0.017725f
C1495 VDD2.n37 VSUBS 0.016741f
C1496 VDD2.n38 VSUBS 0.031154f
C1497 VDD2.n39 VSUBS 0.031154f
C1498 VDD2.n40 VSUBS 0.016741f
C1499 VDD2.n41 VSUBS 0.017233f
C1500 VDD2.n42 VSUBS 0.017233f
C1501 VDD2.n43 VSUBS 0.039569f
C1502 VDD2.n44 VSUBS 0.039569f
C1503 VDD2.n45 VSUBS 0.017725f
C1504 VDD2.n46 VSUBS 0.016741f
C1505 VDD2.n47 VSUBS 0.031154f
C1506 VDD2.n48 VSUBS 0.031154f
C1507 VDD2.n49 VSUBS 0.016741f
C1508 VDD2.n50 VSUBS 0.017725f
C1509 VDD2.n51 VSUBS 0.039569f
C1510 VDD2.n52 VSUBS 0.094898f
C1511 VDD2.n53 VSUBS 0.017725f
C1512 VDD2.n54 VSUBS 0.016741f
C1513 VDD2.n55 VSUBS 0.074989f
C1514 VDD2.n56 VSUBS 0.089094f
C1515 VDD2.t8 VSUBS 0.264649f
C1516 VDD2.t7 VSUBS 0.264649f
C1517 VDD2.n57 VSUBS 2.03044f
C1518 VDD2.n58 VSUBS 1.27029f
C1519 VDD2.t2 VSUBS 0.264649f
C1520 VDD2.t0 VSUBS 0.264649f
C1521 VDD2.n59 VSUBS 2.0601f
C1522 VDD2.n60 VSUBS 4.14931f
C1523 VDD2.n61 VSUBS 0.033969f
C1524 VDD2.n62 VSUBS 0.031154f
C1525 VDD2.n63 VSUBS 0.016741f
C1526 VDD2.n64 VSUBS 0.039569f
C1527 VDD2.n65 VSUBS 0.017725f
C1528 VDD2.n66 VSUBS 0.031154f
C1529 VDD2.n67 VSUBS 0.016741f
C1530 VDD2.n68 VSUBS 0.039569f
C1531 VDD2.n69 VSUBS 0.017725f
C1532 VDD2.n70 VSUBS 0.031154f
C1533 VDD2.n71 VSUBS 0.016741f
C1534 VDD2.n72 VSUBS 0.039569f
C1535 VDD2.n73 VSUBS 0.039569f
C1536 VDD2.n74 VSUBS 0.017725f
C1537 VDD2.n75 VSUBS 0.031154f
C1538 VDD2.n76 VSUBS 0.016741f
C1539 VDD2.n77 VSUBS 0.039569f
C1540 VDD2.n78 VSUBS 0.017725f
C1541 VDD2.n79 VSUBS 0.227757f
C1542 VDD2.t3 VSUBS 0.085148f
C1543 VDD2.n80 VSUBS 0.029677f
C1544 VDD2.n81 VSUBS 0.029766f
C1545 VDD2.n82 VSUBS 0.016741f
C1546 VDD2.n83 VSUBS 1.36002f
C1547 VDD2.n84 VSUBS 0.031154f
C1548 VDD2.n85 VSUBS 0.016741f
C1549 VDD2.n86 VSUBS 0.017725f
C1550 VDD2.n87 VSUBS 0.039569f
C1551 VDD2.n88 VSUBS 0.039569f
C1552 VDD2.n89 VSUBS 0.017725f
C1553 VDD2.n90 VSUBS 0.016741f
C1554 VDD2.n91 VSUBS 0.031154f
C1555 VDD2.n92 VSUBS 0.031154f
C1556 VDD2.n93 VSUBS 0.016741f
C1557 VDD2.n94 VSUBS 0.017725f
C1558 VDD2.n95 VSUBS 0.039569f
C1559 VDD2.n96 VSUBS 0.039569f
C1560 VDD2.n97 VSUBS 0.017725f
C1561 VDD2.n98 VSUBS 0.016741f
C1562 VDD2.n99 VSUBS 0.031154f
C1563 VDD2.n100 VSUBS 0.031154f
C1564 VDD2.n101 VSUBS 0.016741f
C1565 VDD2.n102 VSUBS 0.017233f
C1566 VDD2.n103 VSUBS 0.017233f
C1567 VDD2.n104 VSUBS 0.039569f
C1568 VDD2.n105 VSUBS 0.039569f
C1569 VDD2.n106 VSUBS 0.017725f
C1570 VDD2.n107 VSUBS 0.016741f
C1571 VDD2.n108 VSUBS 0.031154f
C1572 VDD2.n109 VSUBS 0.031154f
C1573 VDD2.n110 VSUBS 0.016741f
C1574 VDD2.n111 VSUBS 0.017725f
C1575 VDD2.n112 VSUBS 0.039569f
C1576 VDD2.n113 VSUBS 0.094898f
C1577 VDD2.n114 VSUBS 0.017725f
C1578 VDD2.n115 VSUBS 0.016741f
C1579 VDD2.n116 VSUBS 0.074989f
C1580 VDD2.n117 VSUBS 0.069262f
C1581 VDD2.n118 VSUBS 3.72139f
C1582 VDD2.t9 VSUBS 0.264649f
C1583 VDD2.t4 VSUBS 0.264649f
C1584 VDD2.n119 VSUBS 2.03045f
C1585 VDD2.n120 VSUBS 0.942796f
C1586 VDD2.t6 VSUBS 0.264649f
C1587 VDD2.t1 VSUBS 0.264649f
C1588 VDD2.n121 VSUBS 2.06005f
C1589 VN.t4 VSUBS 2.4083f
C1590 VN.n0 VSUBS 0.955274f
C1591 VN.n1 VSUBS 0.026698f
C1592 VN.n2 VSUBS 0.028002f
C1593 VN.n3 VSUBS 0.026698f
C1594 VN.t0 VSUBS 2.4083f
C1595 VN.n4 VSUBS 0.853023f
C1596 VN.n5 VSUBS 0.026698f
C1597 VN.n6 VSUBS 0.035999f
C1598 VN.n7 VSUBS 0.026698f
C1599 VN.t8 VSUBS 2.4083f
C1600 VN.n8 VSUBS 0.049759f
C1601 VN.n9 VSUBS 0.026698f
C1602 VN.n10 VSUBS 0.049759f
C1603 VN.t9 VSUBS 2.70311f
C1604 VN.n11 VSUBS 0.899337f
C1605 VN.t1 VSUBS 2.4083f
C1606 VN.n12 VSUBS 0.948104f
C1607 VN.n13 VSUBS 0.045828f
C1608 VN.n14 VSUBS 0.306012f
C1609 VN.n15 VSUBS 0.026698f
C1610 VN.n16 VSUBS 0.026698f
C1611 VN.n17 VSUBS 0.041951f
C1612 VN.n18 VSUBS 0.035999f
C1613 VN.n19 VSUBS 0.049759f
C1614 VN.n20 VSUBS 0.026698f
C1615 VN.n21 VSUBS 0.026698f
C1616 VN.n22 VSUBS 0.026698f
C1617 VN.n23 VSUBS 0.878215f
C1618 VN.n24 VSUBS 0.049759f
C1619 VN.n25 VSUBS 0.049759f
C1620 VN.n26 VSUBS 0.026698f
C1621 VN.n27 VSUBS 0.026698f
C1622 VN.n28 VSUBS 0.026698f
C1623 VN.n29 VSUBS 0.041951f
C1624 VN.n30 VSUBS 0.049759f
C1625 VN.n31 VSUBS 0.045828f
C1626 VN.n32 VSUBS 0.026698f
C1627 VN.n33 VSUBS 0.026698f
C1628 VN.n34 VSUBS 0.029123f
C1629 VN.n35 VSUBS 0.049759f
C1630 VN.n36 VSUBS 0.052335f
C1631 VN.n37 VSUBS 0.026698f
C1632 VN.n38 VSUBS 0.026698f
C1633 VN.n39 VSUBS 0.026698f
C1634 VN.n40 VSUBS 0.047371f
C1635 VN.n41 VSUBS 0.049759f
C1636 VN.n42 VSUBS 0.041898f
C1637 VN.n43 VSUBS 0.04309f
C1638 VN.n44 VSUBS 0.060269f
C1639 VN.t5 VSUBS 2.4083f
C1640 VN.n45 VSUBS 0.955274f
C1641 VN.n46 VSUBS 0.026698f
C1642 VN.n47 VSUBS 0.028002f
C1643 VN.n48 VSUBS 0.026698f
C1644 VN.t2 VSUBS 2.4083f
C1645 VN.n49 VSUBS 0.853023f
C1646 VN.n50 VSUBS 0.026698f
C1647 VN.n51 VSUBS 0.035999f
C1648 VN.n52 VSUBS 0.026698f
C1649 VN.t7 VSUBS 2.4083f
C1650 VN.n53 VSUBS 0.049759f
C1651 VN.n54 VSUBS 0.026698f
C1652 VN.n55 VSUBS 0.049759f
C1653 VN.t3 VSUBS 2.70311f
C1654 VN.n56 VSUBS 0.899337f
C1655 VN.t6 VSUBS 2.4083f
C1656 VN.n57 VSUBS 0.948104f
C1657 VN.n58 VSUBS 0.045828f
C1658 VN.n59 VSUBS 0.306012f
C1659 VN.n60 VSUBS 0.026698f
C1660 VN.n61 VSUBS 0.026698f
C1661 VN.n62 VSUBS 0.041951f
C1662 VN.n63 VSUBS 0.035999f
C1663 VN.n64 VSUBS 0.049759f
C1664 VN.n65 VSUBS 0.026698f
C1665 VN.n66 VSUBS 0.026698f
C1666 VN.n67 VSUBS 0.026698f
C1667 VN.n68 VSUBS 0.878215f
C1668 VN.n69 VSUBS 0.049759f
C1669 VN.n70 VSUBS 0.049759f
C1670 VN.n71 VSUBS 0.026698f
C1671 VN.n72 VSUBS 0.026698f
C1672 VN.n73 VSUBS 0.026698f
C1673 VN.n74 VSUBS 0.041951f
C1674 VN.n75 VSUBS 0.049759f
C1675 VN.n76 VSUBS 0.045828f
C1676 VN.n77 VSUBS 0.026698f
C1677 VN.n78 VSUBS 0.026698f
C1678 VN.n79 VSUBS 0.029123f
C1679 VN.n80 VSUBS 0.049759f
C1680 VN.n81 VSUBS 0.052335f
C1681 VN.n82 VSUBS 0.026698f
C1682 VN.n83 VSUBS 0.026698f
C1683 VN.n84 VSUBS 0.026698f
C1684 VN.n85 VSUBS 0.047371f
C1685 VN.n86 VSUBS 0.049759f
C1686 VN.n87 VSUBS 0.041898f
C1687 VN.n88 VSUBS 0.04309f
C1688 VN.n89 VSUBS 1.73879f
.ends

