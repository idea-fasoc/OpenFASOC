* NGSPICE file created from diff_pair_sample_0893.ext - technology: sky130A

.subckt diff_pair_sample_0893 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=2.66
X1 VDD2.t5 VN.t0 VTAIL.t1 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=2.66
X2 VTAIL.t5 VN.t1 VDD2.t4 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=2.66
X3 B.t11 B.t9 B.t10 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=2.66
X4 VTAIL.t7 VP.t1 VDD1.t4 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=2.66
X5 VDD2.t3 VN.t2 VTAIL.t2 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=2.66
X6 VTAIL.t3 VN.t3 VDD2.t2 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=2.66
X7 B.t8 B.t6 B.t7 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=2.66
X8 B.t5 B.t3 B.t4 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=2.66
X9 VDD1.t3 VP.t2 VTAIL.t6 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=2.66
X10 VDD2.t1 VN.t4 VTAIL.t4 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=2.66
X11 VDD2.t0 VN.t5 VTAIL.t0 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=2.66
X12 VDD1.t2 VP.t3 VTAIL.t9 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=5.148 ps=27.18 w=13.2 l=2.66
X13 B.t2 B.t0 B.t1 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=0 ps=0 w=13.2 l=2.66
X14 VTAIL.t11 VP.t4 VDD1.t1 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=2.178 pd=13.53 as=2.178 ps=13.53 w=13.2 l=2.66
X15 VDD1.t0 VP.t5 VTAIL.t10 w_n3362_n3608# sky130_fd_pr__pfet_01v8 ad=5.148 pd=27.18 as=2.178 ps=13.53 w=13.2 l=2.66
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n38 VP.n37 161.3
R6 VP.n36 VP.n1 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n33 VP.n2 161.3
R9 VP.n32 VP.n31 161.3
R10 VP.n30 VP.n3 161.3
R11 VP.n29 VP.n28 161.3
R12 VP.n27 VP.n4 161.3
R13 VP.n26 VP.n25 161.3
R14 VP.n24 VP.n5 161.3
R15 VP.n23 VP.n22 161.3
R16 VP.n10 VP.t2 151.821
R17 VP.n30 VP.t4 119.594
R18 VP.n6 VP.t5 119.594
R19 VP.n0 VP.t3 119.594
R20 VP.n11 VP.t1 119.594
R21 VP.n7 VP.t0 119.594
R22 VP.n21 VP.n6 66.1456
R23 VP.n39 VP.n0 66.1456
R24 VP.n20 VP.n7 66.1456
R25 VP.n21 VP.n20 49.92
R26 VP.n11 VP.n10 49.0206
R27 VP.n25 VP.n4 41.0614
R28 VP.n35 VP.n2 41.0614
R29 VP.n16 VP.n9 41.0614
R30 VP.n25 VP.n24 40.0926
R31 VP.n36 VP.n35 40.0926
R32 VP.n17 VP.n16 40.0926
R33 VP.n24 VP.n23 24.5923
R34 VP.n29 VP.n4 24.5923
R35 VP.n30 VP.n29 24.5923
R36 VP.n31 VP.n30 24.5923
R37 VP.n31 VP.n2 24.5923
R38 VP.n37 VP.n36 24.5923
R39 VP.n18 VP.n17 24.5923
R40 VP.n12 VP.n11 24.5923
R41 VP.n12 VP.n9 24.5923
R42 VP.n23 VP.n6 24.1005
R43 VP.n37 VP.n0 24.1005
R44 VP.n18 VP.n7 24.1005
R45 VP.n13 VP.n10 5.20743
R46 VP.n20 VP.n19 0.354861
R47 VP.n22 VP.n21 0.354861
R48 VP.n39 VP.n38 0.354861
R49 VP VP.n39 0.267071
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n8 0.189894
R53 VP.n19 VP.n8 0.189894
R54 VP.n22 VP.n5 0.189894
R55 VP.n26 VP.n5 0.189894
R56 VP.n27 VP.n26 0.189894
R57 VP.n28 VP.n27 0.189894
R58 VP.n28 VP.n3 0.189894
R59 VP.n32 VP.n3 0.189894
R60 VP.n33 VP.n32 0.189894
R61 VP.n34 VP.n33 0.189894
R62 VP.n34 VP.n1 0.189894
R63 VP.n38 VP.n1 0.189894
R64 VTAIL.n7 VTAIL.t4 58.4184
R65 VTAIL.n11 VTAIL.t0 58.4181
R66 VTAIL.n2 VTAIL.t9 58.4181
R67 VTAIL.n10 VTAIL.t8 58.4181
R68 VTAIL.n9 VTAIL.n8 55.9559
R69 VTAIL.n6 VTAIL.n5 55.9559
R70 VTAIL.n1 VTAIL.n0 55.9558
R71 VTAIL.n4 VTAIL.n3 55.9558
R72 VTAIL.n6 VTAIL.n4 28.9014
R73 VTAIL.n11 VTAIL.n10 26.3238
R74 VTAIL.n7 VTAIL.n6 2.57809
R75 VTAIL.n10 VTAIL.n9 2.57809
R76 VTAIL.n4 VTAIL.n2 2.57809
R77 VTAIL.n0 VTAIL.t1 2.463
R78 VTAIL.n0 VTAIL.t5 2.463
R79 VTAIL.n3 VTAIL.t10 2.463
R80 VTAIL.n3 VTAIL.t11 2.463
R81 VTAIL.n8 VTAIL.t6 2.463
R82 VTAIL.n8 VTAIL.t7 2.463
R83 VTAIL.n5 VTAIL.t2 2.463
R84 VTAIL.n5 VTAIL.t3 2.463
R85 VTAIL VTAIL.n11 1.8755
R86 VTAIL.n9 VTAIL.n7 1.75912
R87 VTAIL.n2 VTAIL.n1 1.75912
R88 VTAIL VTAIL.n1 0.703086
R89 VDD1 VDD1.t3 77.0886
R90 VDD1.n1 VDD1.t0 76.9748
R91 VDD1.n1 VDD1.n0 73.2237
R92 VDD1.n3 VDD1.n2 72.6345
R93 VDD1.n3 VDD1.n1 45.3436
R94 VDD1.n2 VDD1.t4 2.463
R95 VDD1.n2 VDD1.t5 2.463
R96 VDD1.n0 VDD1.t1 2.463
R97 VDD1.n0 VDD1.t2 2.463
R98 VDD1 VDD1.n3 0.586707
R99 VN.n26 VN.n25 161.3
R100 VN.n24 VN.n15 161.3
R101 VN.n23 VN.n22 161.3
R102 VN.n21 VN.n16 161.3
R103 VN.n20 VN.n19 161.3
R104 VN.n12 VN.n11 161.3
R105 VN.n10 VN.n1 161.3
R106 VN.n9 VN.n8 161.3
R107 VN.n7 VN.n2 161.3
R108 VN.n6 VN.n5 161.3
R109 VN.n17 VN.t4 151.821
R110 VN.n3 VN.t0 151.821
R111 VN.n4 VN.t1 119.594
R112 VN.n0 VN.t5 119.594
R113 VN.n18 VN.t3 119.594
R114 VN.n14 VN.t2 119.594
R115 VN.n13 VN.n0 66.1456
R116 VN.n27 VN.n14 66.1456
R117 VN VN.n27 50.0853
R118 VN.n4 VN.n3 49.0206
R119 VN.n18 VN.n17 49.0206
R120 VN.n9 VN.n2 41.0614
R121 VN.n23 VN.n16 41.0614
R122 VN.n10 VN.n9 40.0926
R123 VN.n24 VN.n23 40.0926
R124 VN.n5 VN.n4 24.5923
R125 VN.n5 VN.n2 24.5923
R126 VN.n11 VN.n10 24.5923
R127 VN.n19 VN.n16 24.5923
R128 VN.n19 VN.n18 24.5923
R129 VN.n25 VN.n24 24.5923
R130 VN.n11 VN.n0 24.1005
R131 VN.n25 VN.n14 24.1005
R132 VN.n20 VN.n17 5.20746
R133 VN.n6 VN.n3 5.20746
R134 VN.n27 VN.n26 0.354861
R135 VN.n13 VN.n12 0.354861
R136 VN VN.n13 0.267071
R137 VN.n26 VN.n15 0.189894
R138 VN.n22 VN.n15 0.189894
R139 VN.n22 VN.n21 0.189894
R140 VN.n21 VN.n20 0.189894
R141 VN.n7 VN.n6 0.189894
R142 VN.n8 VN.n7 0.189894
R143 VN.n8 VN.n1 0.189894
R144 VN.n12 VN.n1 0.189894
R145 VDD2.n1 VDD2.t5 76.9748
R146 VDD2.n2 VDD2.t3 75.0972
R147 VDD2.n1 VDD2.n0 73.2237
R148 VDD2 VDD2.n3 73.2207
R149 VDD2.n2 VDD2.n1 43.4718
R150 VDD2.n3 VDD2.t2 2.463
R151 VDD2.n3 VDD2.t1 2.463
R152 VDD2.n0 VDD2.t4 2.463
R153 VDD2.n0 VDD2.t0 2.463
R154 VDD2 VDD2.n2 1.99188
R155 B.n411 B.n122 585
R156 B.n410 B.n409 585
R157 B.n408 B.n123 585
R158 B.n407 B.n406 585
R159 B.n405 B.n124 585
R160 B.n404 B.n403 585
R161 B.n402 B.n125 585
R162 B.n401 B.n400 585
R163 B.n399 B.n126 585
R164 B.n398 B.n397 585
R165 B.n396 B.n127 585
R166 B.n395 B.n394 585
R167 B.n393 B.n128 585
R168 B.n392 B.n391 585
R169 B.n390 B.n129 585
R170 B.n389 B.n388 585
R171 B.n387 B.n130 585
R172 B.n386 B.n385 585
R173 B.n384 B.n131 585
R174 B.n383 B.n382 585
R175 B.n381 B.n132 585
R176 B.n380 B.n379 585
R177 B.n378 B.n133 585
R178 B.n377 B.n376 585
R179 B.n375 B.n134 585
R180 B.n374 B.n373 585
R181 B.n372 B.n135 585
R182 B.n371 B.n370 585
R183 B.n369 B.n136 585
R184 B.n368 B.n367 585
R185 B.n366 B.n137 585
R186 B.n365 B.n364 585
R187 B.n363 B.n138 585
R188 B.n362 B.n361 585
R189 B.n360 B.n139 585
R190 B.n359 B.n358 585
R191 B.n357 B.n140 585
R192 B.n356 B.n355 585
R193 B.n354 B.n141 585
R194 B.n353 B.n352 585
R195 B.n351 B.n142 585
R196 B.n350 B.n349 585
R197 B.n348 B.n143 585
R198 B.n347 B.n346 585
R199 B.n345 B.n144 585
R200 B.n344 B.n343 585
R201 B.n339 B.n145 585
R202 B.n338 B.n337 585
R203 B.n336 B.n146 585
R204 B.n335 B.n334 585
R205 B.n333 B.n147 585
R206 B.n332 B.n331 585
R207 B.n330 B.n148 585
R208 B.n329 B.n328 585
R209 B.n327 B.n149 585
R210 B.n325 B.n324 585
R211 B.n323 B.n152 585
R212 B.n322 B.n321 585
R213 B.n320 B.n153 585
R214 B.n319 B.n318 585
R215 B.n317 B.n154 585
R216 B.n316 B.n315 585
R217 B.n314 B.n155 585
R218 B.n313 B.n312 585
R219 B.n311 B.n156 585
R220 B.n310 B.n309 585
R221 B.n308 B.n157 585
R222 B.n307 B.n306 585
R223 B.n305 B.n158 585
R224 B.n304 B.n303 585
R225 B.n302 B.n159 585
R226 B.n301 B.n300 585
R227 B.n299 B.n160 585
R228 B.n298 B.n297 585
R229 B.n296 B.n161 585
R230 B.n295 B.n294 585
R231 B.n293 B.n162 585
R232 B.n292 B.n291 585
R233 B.n290 B.n163 585
R234 B.n289 B.n288 585
R235 B.n287 B.n164 585
R236 B.n286 B.n285 585
R237 B.n284 B.n165 585
R238 B.n283 B.n282 585
R239 B.n281 B.n166 585
R240 B.n280 B.n279 585
R241 B.n278 B.n167 585
R242 B.n277 B.n276 585
R243 B.n275 B.n168 585
R244 B.n274 B.n273 585
R245 B.n272 B.n169 585
R246 B.n271 B.n270 585
R247 B.n269 B.n170 585
R248 B.n268 B.n267 585
R249 B.n266 B.n171 585
R250 B.n265 B.n264 585
R251 B.n263 B.n172 585
R252 B.n262 B.n261 585
R253 B.n260 B.n173 585
R254 B.n259 B.n258 585
R255 B.n413 B.n412 585
R256 B.n414 B.n121 585
R257 B.n416 B.n415 585
R258 B.n417 B.n120 585
R259 B.n419 B.n418 585
R260 B.n420 B.n119 585
R261 B.n422 B.n421 585
R262 B.n423 B.n118 585
R263 B.n425 B.n424 585
R264 B.n426 B.n117 585
R265 B.n428 B.n427 585
R266 B.n429 B.n116 585
R267 B.n431 B.n430 585
R268 B.n432 B.n115 585
R269 B.n434 B.n433 585
R270 B.n435 B.n114 585
R271 B.n437 B.n436 585
R272 B.n438 B.n113 585
R273 B.n440 B.n439 585
R274 B.n441 B.n112 585
R275 B.n443 B.n442 585
R276 B.n444 B.n111 585
R277 B.n446 B.n445 585
R278 B.n447 B.n110 585
R279 B.n449 B.n448 585
R280 B.n450 B.n109 585
R281 B.n452 B.n451 585
R282 B.n453 B.n108 585
R283 B.n455 B.n454 585
R284 B.n456 B.n107 585
R285 B.n458 B.n457 585
R286 B.n459 B.n106 585
R287 B.n461 B.n460 585
R288 B.n462 B.n105 585
R289 B.n464 B.n463 585
R290 B.n465 B.n104 585
R291 B.n467 B.n466 585
R292 B.n468 B.n103 585
R293 B.n470 B.n469 585
R294 B.n471 B.n102 585
R295 B.n473 B.n472 585
R296 B.n474 B.n101 585
R297 B.n476 B.n475 585
R298 B.n477 B.n100 585
R299 B.n479 B.n478 585
R300 B.n480 B.n99 585
R301 B.n482 B.n481 585
R302 B.n483 B.n98 585
R303 B.n485 B.n484 585
R304 B.n486 B.n97 585
R305 B.n488 B.n487 585
R306 B.n489 B.n96 585
R307 B.n491 B.n490 585
R308 B.n492 B.n95 585
R309 B.n494 B.n493 585
R310 B.n495 B.n94 585
R311 B.n497 B.n496 585
R312 B.n498 B.n93 585
R313 B.n500 B.n499 585
R314 B.n501 B.n92 585
R315 B.n503 B.n502 585
R316 B.n504 B.n91 585
R317 B.n506 B.n505 585
R318 B.n507 B.n90 585
R319 B.n509 B.n508 585
R320 B.n510 B.n89 585
R321 B.n512 B.n511 585
R322 B.n513 B.n88 585
R323 B.n515 B.n514 585
R324 B.n516 B.n87 585
R325 B.n518 B.n517 585
R326 B.n519 B.n86 585
R327 B.n521 B.n520 585
R328 B.n522 B.n85 585
R329 B.n524 B.n523 585
R330 B.n525 B.n84 585
R331 B.n527 B.n526 585
R332 B.n528 B.n83 585
R333 B.n530 B.n529 585
R334 B.n531 B.n82 585
R335 B.n533 B.n532 585
R336 B.n534 B.n81 585
R337 B.n536 B.n535 585
R338 B.n537 B.n80 585
R339 B.n539 B.n538 585
R340 B.n540 B.n79 585
R341 B.n542 B.n541 585
R342 B.n543 B.n78 585
R343 B.n695 B.n694 585
R344 B.n693 B.n24 585
R345 B.n692 B.n691 585
R346 B.n690 B.n25 585
R347 B.n689 B.n688 585
R348 B.n687 B.n26 585
R349 B.n686 B.n685 585
R350 B.n684 B.n27 585
R351 B.n683 B.n682 585
R352 B.n681 B.n28 585
R353 B.n680 B.n679 585
R354 B.n678 B.n29 585
R355 B.n677 B.n676 585
R356 B.n675 B.n30 585
R357 B.n674 B.n673 585
R358 B.n672 B.n31 585
R359 B.n671 B.n670 585
R360 B.n669 B.n32 585
R361 B.n668 B.n667 585
R362 B.n666 B.n33 585
R363 B.n665 B.n664 585
R364 B.n663 B.n34 585
R365 B.n662 B.n661 585
R366 B.n660 B.n35 585
R367 B.n659 B.n658 585
R368 B.n657 B.n36 585
R369 B.n656 B.n655 585
R370 B.n654 B.n37 585
R371 B.n653 B.n652 585
R372 B.n651 B.n38 585
R373 B.n650 B.n649 585
R374 B.n648 B.n39 585
R375 B.n647 B.n646 585
R376 B.n645 B.n40 585
R377 B.n644 B.n643 585
R378 B.n642 B.n41 585
R379 B.n641 B.n640 585
R380 B.n639 B.n42 585
R381 B.n638 B.n637 585
R382 B.n636 B.n43 585
R383 B.n635 B.n634 585
R384 B.n633 B.n44 585
R385 B.n632 B.n631 585
R386 B.n630 B.n45 585
R387 B.n629 B.n628 585
R388 B.n627 B.n626 585
R389 B.n625 B.n49 585
R390 B.n624 B.n623 585
R391 B.n622 B.n50 585
R392 B.n621 B.n620 585
R393 B.n619 B.n51 585
R394 B.n618 B.n617 585
R395 B.n616 B.n52 585
R396 B.n615 B.n614 585
R397 B.n613 B.n53 585
R398 B.n611 B.n610 585
R399 B.n609 B.n56 585
R400 B.n608 B.n607 585
R401 B.n606 B.n57 585
R402 B.n605 B.n604 585
R403 B.n603 B.n58 585
R404 B.n602 B.n601 585
R405 B.n600 B.n59 585
R406 B.n599 B.n598 585
R407 B.n597 B.n60 585
R408 B.n596 B.n595 585
R409 B.n594 B.n61 585
R410 B.n593 B.n592 585
R411 B.n591 B.n62 585
R412 B.n590 B.n589 585
R413 B.n588 B.n63 585
R414 B.n587 B.n586 585
R415 B.n585 B.n64 585
R416 B.n584 B.n583 585
R417 B.n582 B.n65 585
R418 B.n581 B.n580 585
R419 B.n579 B.n66 585
R420 B.n578 B.n577 585
R421 B.n576 B.n67 585
R422 B.n575 B.n574 585
R423 B.n573 B.n68 585
R424 B.n572 B.n571 585
R425 B.n570 B.n69 585
R426 B.n569 B.n568 585
R427 B.n567 B.n70 585
R428 B.n566 B.n565 585
R429 B.n564 B.n71 585
R430 B.n563 B.n562 585
R431 B.n561 B.n72 585
R432 B.n560 B.n559 585
R433 B.n558 B.n73 585
R434 B.n557 B.n556 585
R435 B.n555 B.n74 585
R436 B.n554 B.n553 585
R437 B.n552 B.n75 585
R438 B.n551 B.n550 585
R439 B.n549 B.n76 585
R440 B.n548 B.n547 585
R441 B.n546 B.n77 585
R442 B.n545 B.n544 585
R443 B.n696 B.n23 585
R444 B.n698 B.n697 585
R445 B.n699 B.n22 585
R446 B.n701 B.n700 585
R447 B.n702 B.n21 585
R448 B.n704 B.n703 585
R449 B.n705 B.n20 585
R450 B.n707 B.n706 585
R451 B.n708 B.n19 585
R452 B.n710 B.n709 585
R453 B.n711 B.n18 585
R454 B.n713 B.n712 585
R455 B.n714 B.n17 585
R456 B.n716 B.n715 585
R457 B.n717 B.n16 585
R458 B.n719 B.n718 585
R459 B.n720 B.n15 585
R460 B.n722 B.n721 585
R461 B.n723 B.n14 585
R462 B.n725 B.n724 585
R463 B.n726 B.n13 585
R464 B.n728 B.n727 585
R465 B.n729 B.n12 585
R466 B.n731 B.n730 585
R467 B.n732 B.n11 585
R468 B.n734 B.n733 585
R469 B.n735 B.n10 585
R470 B.n737 B.n736 585
R471 B.n738 B.n9 585
R472 B.n740 B.n739 585
R473 B.n741 B.n8 585
R474 B.n743 B.n742 585
R475 B.n744 B.n7 585
R476 B.n746 B.n745 585
R477 B.n747 B.n6 585
R478 B.n749 B.n748 585
R479 B.n750 B.n5 585
R480 B.n752 B.n751 585
R481 B.n753 B.n4 585
R482 B.n755 B.n754 585
R483 B.n756 B.n3 585
R484 B.n758 B.n757 585
R485 B.n759 B.n0 585
R486 B.n2 B.n1 585
R487 B.n196 B.n195 585
R488 B.n197 B.n194 585
R489 B.n199 B.n198 585
R490 B.n200 B.n193 585
R491 B.n202 B.n201 585
R492 B.n203 B.n192 585
R493 B.n205 B.n204 585
R494 B.n206 B.n191 585
R495 B.n208 B.n207 585
R496 B.n209 B.n190 585
R497 B.n211 B.n210 585
R498 B.n212 B.n189 585
R499 B.n214 B.n213 585
R500 B.n215 B.n188 585
R501 B.n217 B.n216 585
R502 B.n218 B.n187 585
R503 B.n220 B.n219 585
R504 B.n221 B.n186 585
R505 B.n223 B.n222 585
R506 B.n224 B.n185 585
R507 B.n226 B.n225 585
R508 B.n227 B.n184 585
R509 B.n229 B.n228 585
R510 B.n230 B.n183 585
R511 B.n232 B.n231 585
R512 B.n233 B.n182 585
R513 B.n235 B.n234 585
R514 B.n236 B.n181 585
R515 B.n238 B.n237 585
R516 B.n239 B.n180 585
R517 B.n241 B.n240 585
R518 B.n242 B.n179 585
R519 B.n244 B.n243 585
R520 B.n245 B.n178 585
R521 B.n247 B.n246 585
R522 B.n248 B.n177 585
R523 B.n250 B.n249 585
R524 B.n251 B.n176 585
R525 B.n253 B.n252 585
R526 B.n254 B.n175 585
R527 B.n256 B.n255 585
R528 B.n257 B.n174 585
R529 B.n258 B.n257 454.062
R530 B.n412 B.n411 454.062
R531 B.n544 B.n543 454.062
R532 B.n694 B.n23 454.062
R533 B.n150 B.t9 327.729
R534 B.n340 B.t6 327.729
R535 B.n54 B.t0 327.729
R536 B.n46 B.t3 327.729
R537 B.n761 B.n760 256.663
R538 B.n760 B.n759 235.042
R539 B.n760 B.n2 235.042
R540 B.n340 B.t7 170.274
R541 B.n54 B.t2 170.274
R542 B.n150 B.t10 170.258
R543 B.n46 B.t5 170.258
R544 B.n258 B.n173 163.367
R545 B.n262 B.n173 163.367
R546 B.n263 B.n262 163.367
R547 B.n264 B.n263 163.367
R548 B.n264 B.n171 163.367
R549 B.n268 B.n171 163.367
R550 B.n269 B.n268 163.367
R551 B.n270 B.n269 163.367
R552 B.n270 B.n169 163.367
R553 B.n274 B.n169 163.367
R554 B.n275 B.n274 163.367
R555 B.n276 B.n275 163.367
R556 B.n276 B.n167 163.367
R557 B.n280 B.n167 163.367
R558 B.n281 B.n280 163.367
R559 B.n282 B.n281 163.367
R560 B.n282 B.n165 163.367
R561 B.n286 B.n165 163.367
R562 B.n287 B.n286 163.367
R563 B.n288 B.n287 163.367
R564 B.n288 B.n163 163.367
R565 B.n292 B.n163 163.367
R566 B.n293 B.n292 163.367
R567 B.n294 B.n293 163.367
R568 B.n294 B.n161 163.367
R569 B.n298 B.n161 163.367
R570 B.n299 B.n298 163.367
R571 B.n300 B.n299 163.367
R572 B.n300 B.n159 163.367
R573 B.n304 B.n159 163.367
R574 B.n305 B.n304 163.367
R575 B.n306 B.n305 163.367
R576 B.n306 B.n157 163.367
R577 B.n310 B.n157 163.367
R578 B.n311 B.n310 163.367
R579 B.n312 B.n311 163.367
R580 B.n312 B.n155 163.367
R581 B.n316 B.n155 163.367
R582 B.n317 B.n316 163.367
R583 B.n318 B.n317 163.367
R584 B.n318 B.n153 163.367
R585 B.n322 B.n153 163.367
R586 B.n323 B.n322 163.367
R587 B.n324 B.n323 163.367
R588 B.n324 B.n149 163.367
R589 B.n329 B.n149 163.367
R590 B.n330 B.n329 163.367
R591 B.n331 B.n330 163.367
R592 B.n331 B.n147 163.367
R593 B.n335 B.n147 163.367
R594 B.n336 B.n335 163.367
R595 B.n337 B.n336 163.367
R596 B.n337 B.n145 163.367
R597 B.n344 B.n145 163.367
R598 B.n345 B.n344 163.367
R599 B.n346 B.n345 163.367
R600 B.n346 B.n143 163.367
R601 B.n350 B.n143 163.367
R602 B.n351 B.n350 163.367
R603 B.n352 B.n351 163.367
R604 B.n352 B.n141 163.367
R605 B.n356 B.n141 163.367
R606 B.n357 B.n356 163.367
R607 B.n358 B.n357 163.367
R608 B.n358 B.n139 163.367
R609 B.n362 B.n139 163.367
R610 B.n363 B.n362 163.367
R611 B.n364 B.n363 163.367
R612 B.n364 B.n137 163.367
R613 B.n368 B.n137 163.367
R614 B.n369 B.n368 163.367
R615 B.n370 B.n369 163.367
R616 B.n370 B.n135 163.367
R617 B.n374 B.n135 163.367
R618 B.n375 B.n374 163.367
R619 B.n376 B.n375 163.367
R620 B.n376 B.n133 163.367
R621 B.n380 B.n133 163.367
R622 B.n381 B.n380 163.367
R623 B.n382 B.n381 163.367
R624 B.n382 B.n131 163.367
R625 B.n386 B.n131 163.367
R626 B.n387 B.n386 163.367
R627 B.n388 B.n387 163.367
R628 B.n388 B.n129 163.367
R629 B.n392 B.n129 163.367
R630 B.n393 B.n392 163.367
R631 B.n394 B.n393 163.367
R632 B.n394 B.n127 163.367
R633 B.n398 B.n127 163.367
R634 B.n399 B.n398 163.367
R635 B.n400 B.n399 163.367
R636 B.n400 B.n125 163.367
R637 B.n404 B.n125 163.367
R638 B.n405 B.n404 163.367
R639 B.n406 B.n405 163.367
R640 B.n406 B.n123 163.367
R641 B.n410 B.n123 163.367
R642 B.n411 B.n410 163.367
R643 B.n543 B.n542 163.367
R644 B.n542 B.n79 163.367
R645 B.n538 B.n79 163.367
R646 B.n538 B.n537 163.367
R647 B.n537 B.n536 163.367
R648 B.n536 B.n81 163.367
R649 B.n532 B.n81 163.367
R650 B.n532 B.n531 163.367
R651 B.n531 B.n530 163.367
R652 B.n530 B.n83 163.367
R653 B.n526 B.n83 163.367
R654 B.n526 B.n525 163.367
R655 B.n525 B.n524 163.367
R656 B.n524 B.n85 163.367
R657 B.n520 B.n85 163.367
R658 B.n520 B.n519 163.367
R659 B.n519 B.n518 163.367
R660 B.n518 B.n87 163.367
R661 B.n514 B.n87 163.367
R662 B.n514 B.n513 163.367
R663 B.n513 B.n512 163.367
R664 B.n512 B.n89 163.367
R665 B.n508 B.n89 163.367
R666 B.n508 B.n507 163.367
R667 B.n507 B.n506 163.367
R668 B.n506 B.n91 163.367
R669 B.n502 B.n91 163.367
R670 B.n502 B.n501 163.367
R671 B.n501 B.n500 163.367
R672 B.n500 B.n93 163.367
R673 B.n496 B.n93 163.367
R674 B.n496 B.n495 163.367
R675 B.n495 B.n494 163.367
R676 B.n494 B.n95 163.367
R677 B.n490 B.n95 163.367
R678 B.n490 B.n489 163.367
R679 B.n489 B.n488 163.367
R680 B.n488 B.n97 163.367
R681 B.n484 B.n97 163.367
R682 B.n484 B.n483 163.367
R683 B.n483 B.n482 163.367
R684 B.n482 B.n99 163.367
R685 B.n478 B.n99 163.367
R686 B.n478 B.n477 163.367
R687 B.n477 B.n476 163.367
R688 B.n476 B.n101 163.367
R689 B.n472 B.n101 163.367
R690 B.n472 B.n471 163.367
R691 B.n471 B.n470 163.367
R692 B.n470 B.n103 163.367
R693 B.n466 B.n103 163.367
R694 B.n466 B.n465 163.367
R695 B.n465 B.n464 163.367
R696 B.n464 B.n105 163.367
R697 B.n460 B.n105 163.367
R698 B.n460 B.n459 163.367
R699 B.n459 B.n458 163.367
R700 B.n458 B.n107 163.367
R701 B.n454 B.n107 163.367
R702 B.n454 B.n453 163.367
R703 B.n453 B.n452 163.367
R704 B.n452 B.n109 163.367
R705 B.n448 B.n109 163.367
R706 B.n448 B.n447 163.367
R707 B.n447 B.n446 163.367
R708 B.n446 B.n111 163.367
R709 B.n442 B.n111 163.367
R710 B.n442 B.n441 163.367
R711 B.n441 B.n440 163.367
R712 B.n440 B.n113 163.367
R713 B.n436 B.n113 163.367
R714 B.n436 B.n435 163.367
R715 B.n435 B.n434 163.367
R716 B.n434 B.n115 163.367
R717 B.n430 B.n115 163.367
R718 B.n430 B.n429 163.367
R719 B.n429 B.n428 163.367
R720 B.n428 B.n117 163.367
R721 B.n424 B.n117 163.367
R722 B.n424 B.n423 163.367
R723 B.n423 B.n422 163.367
R724 B.n422 B.n119 163.367
R725 B.n418 B.n119 163.367
R726 B.n418 B.n417 163.367
R727 B.n417 B.n416 163.367
R728 B.n416 B.n121 163.367
R729 B.n412 B.n121 163.367
R730 B.n694 B.n693 163.367
R731 B.n693 B.n692 163.367
R732 B.n692 B.n25 163.367
R733 B.n688 B.n25 163.367
R734 B.n688 B.n687 163.367
R735 B.n687 B.n686 163.367
R736 B.n686 B.n27 163.367
R737 B.n682 B.n27 163.367
R738 B.n682 B.n681 163.367
R739 B.n681 B.n680 163.367
R740 B.n680 B.n29 163.367
R741 B.n676 B.n29 163.367
R742 B.n676 B.n675 163.367
R743 B.n675 B.n674 163.367
R744 B.n674 B.n31 163.367
R745 B.n670 B.n31 163.367
R746 B.n670 B.n669 163.367
R747 B.n669 B.n668 163.367
R748 B.n668 B.n33 163.367
R749 B.n664 B.n33 163.367
R750 B.n664 B.n663 163.367
R751 B.n663 B.n662 163.367
R752 B.n662 B.n35 163.367
R753 B.n658 B.n35 163.367
R754 B.n658 B.n657 163.367
R755 B.n657 B.n656 163.367
R756 B.n656 B.n37 163.367
R757 B.n652 B.n37 163.367
R758 B.n652 B.n651 163.367
R759 B.n651 B.n650 163.367
R760 B.n650 B.n39 163.367
R761 B.n646 B.n39 163.367
R762 B.n646 B.n645 163.367
R763 B.n645 B.n644 163.367
R764 B.n644 B.n41 163.367
R765 B.n640 B.n41 163.367
R766 B.n640 B.n639 163.367
R767 B.n639 B.n638 163.367
R768 B.n638 B.n43 163.367
R769 B.n634 B.n43 163.367
R770 B.n634 B.n633 163.367
R771 B.n633 B.n632 163.367
R772 B.n632 B.n45 163.367
R773 B.n628 B.n45 163.367
R774 B.n628 B.n627 163.367
R775 B.n627 B.n49 163.367
R776 B.n623 B.n49 163.367
R777 B.n623 B.n622 163.367
R778 B.n622 B.n621 163.367
R779 B.n621 B.n51 163.367
R780 B.n617 B.n51 163.367
R781 B.n617 B.n616 163.367
R782 B.n616 B.n615 163.367
R783 B.n615 B.n53 163.367
R784 B.n610 B.n53 163.367
R785 B.n610 B.n609 163.367
R786 B.n609 B.n608 163.367
R787 B.n608 B.n57 163.367
R788 B.n604 B.n57 163.367
R789 B.n604 B.n603 163.367
R790 B.n603 B.n602 163.367
R791 B.n602 B.n59 163.367
R792 B.n598 B.n59 163.367
R793 B.n598 B.n597 163.367
R794 B.n597 B.n596 163.367
R795 B.n596 B.n61 163.367
R796 B.n592 B.n61 163.367
R797 B.n592 B.n591 163.367
R798 B.n591 B.n590 163.367
R799 B.n590 B.n63 163.367
R800 B.n586 B.n63 163.367
R801 B.n586 B.n585 163.367
R802 B.n585 B.n584 163.367
R803 B.n584 B.n65 163.367
R804 B.n580 B.n65 163.367
R805 B.n580 B.n579 163.367
R806 B.n579 B.n578 163.367
R807 B.n578 B.n67 163.367
R808 B.n574 B.n67 163.367
R809 B.n574 B.n573 163.367
R810 B.n573 B.n572 163.367
R811 B.n572 B.n69 163.367
R812 B.n568 B.n69 163.367
R813 B.n568 B.n567 163.367
R814 B.n567 B.n566 163.367
R815 B.n566 B.n71 163.367
R816 B.n562 B.n71 163.367
R817 B.n562 B.n561 163.367
R818 B.n561 B.n560 163.367
R819 B.n560 B.n73 163.367
R820 B.n556 B.n73 163.367
R821 B.n556 B.n555 163.367
R822 B.n555 B.n554 163.367
R823 B.n554 B.n75 163.367
R824 B.n550 B.n75 163.367
R825 B.n550 B.n549 163.367
R826 B.n549 B.n548 163.367
R827 B.n548 B.n77 163.367
R828 B.n544 B.n77 163.367
R829 B.n698 B.n23 163.367
R830 B.n699 B.n698 163.367
R831 B.n700 B.n699 163.367
R832 B.n700 B.n21 163.367
R833 B.n704 B.n21 163.367
R834 B.n705 B.n704 163.367
R835 B.n706 B.n705 163.367
R836 B.n706 B.n19 163.367
R837 B.n710 B.n19 163.367
R838 B.n711 B.n710 163.367
R839 B.n712 B.n711 163.367
R840 B.n712 B.n17 163.367
R841 B.n716 B.n17 163.367
R842 B.n717 B.n716 163.367
R843 B.n718 B.n717 163.367
R844 B.n718 B.n15 163.367
R845 B.n722 B.n15 163.367
R846 B.n723 B.n722 163.367
R847 B.n724 B.n723 163.367
R848 B.n724 B.n13 163.367
R849 B.n728 B.n13 163.367
R850 B.n729 B.n728 163.367
R851 B.n730 B.n729 163.367
R852 B.n730 B.n11 163.367
R853 B.n734 B.n11 163.367
R854 B.n735 B.n734 163.367
R855 B.n736 B.n735 163.367
R856 B.n736 B.n9 163.367
R857 B.n740 B.n9 163.367
R858 B.n741 B.n740 163.367
R859 B.n742 B.n741 163.367
R860 B.n742 B.n7 163.367
R861 B.n746 B.n7 163.367
R862 B.n747 B.n746 163.367
R863 B.n748 B.n747 163.367
R864 B.n748 B.n5 163.367
R865 B.n752 B.n5 163.367
R866 B.n753 B.n752 163.367
R867 B.n754 B.n753 163.367
R868 B.n754 B.n3 163.367
R869 B.n758 B.n3 163.367
R870 B.n759 B.n758 163.367
R871 B.n196 B.n2 163.367
R872 B.n197 B.n196 163.367
R873 B.n198 B.n197 163.367
R874 B.n198 B.n193 163.367
R875 B.n202 B.n193 163.367
R876 B.n203 B.n202 163.367
R877 B.n204 B.n203 163.367
R878 B.n204 B.n191 163.367
R879 B.n208 B.n191 163.367
R880 B.n209 B.n208 163.367
R881 B.n210 B.n209 163.367
R882 B.n210 B.n189 163.367
R883 B.n214 B.n189 163.367
R884 B.n215 B.n214 163.367
R885 B.n216 B.n215 163.367
R886 B.n216 B.n187 163.367
R887 B.n220 B.n187 163.367
R888 B.n221 B.n220 163.367
R889 B.n222 B.n221 163.367
R890 B.n222 B.n185 163.367
R891 B.n226 B.n185 163.367
R892 B.n227 B.n226 163.367
R893 B.n228 B.n227 163.367
R894 B.n228 B.n183 163.367
R895 B.n232 B.n183 163.367
R896 B.n233 B.n232 163.367
R897 B.n234 B.n233 163.367
R898 B.n234 B.n181 163.367
R899 B.n238 B.n181 163.367
R900 B.n239 B.n238 163.367
R901 B.n240 B.n239 163.367
R902 B.n240 B.n179 163.367
R903 B.n244 B.n179 163.367
R904 B.n245 B.n244 163.367
R905 B.n246 B.n245 163.367
R906 B.n246 B.n177 163.367
R907 B.n250 B.n177 163.367
R908 B.n251 B.n250 163.367
R909 B.n252 B.n251 163.367
R910 B.n252 B.n175 163.367
R911 B.n256 B.n175 163.367
R912 B.n257 B.n256 163.367
R913 B.n341 B.t8 112.287
R914 B.n55 B.t1 112.287
R915 B.n151 B.t11 112.27
R916 B.n47 B.t4 112.27
R917 B.n326 B.n151 59.5399
R918 B.n342 B.n341 59.5399
R919 B.n612 B.n55 59.5399
R920 B.n48 B.n47 59.5399
R921 B.n151 B.n150 57.9884
R922 B.n341 B.n340 57.9884
R923 B.n55 B.n54 57.9884
R924 B.n47 B.n46 57.9884
R925 B.n696 B.n695 29.5029
R926 B.n545 B.n78 29.5029
R927 B.n259 B.n174 29.5029
R928 B.n413 B.n122 29.5029
R929 B B.n761 18.0485
R930 B.n697 B.n696 10.6151
R931 B.n697 B.n22 10.6151
R932 B.n701 B.n22 10.6151
R933 B.n702 B.n701 10.6151
R934 B.n703 B.n702 10.6151
R935 B.n703 B.n20 10.6151
R936 B.n707 B.n20 10.6151
R937 B.n708 B.n707 10.6151
R938 B.n709 B.n708 10.6151
R939 B.n709 B.n18 10.6151
R940 B.n713 B.n18 10.6151
R941 B.n714 B.n713 10.6151
R942 B.n715 B.n714 10.6151
R943 B.n715 B.n16 10.6151
R944 B.n719 B.n16 10.6151
R945 B.n720 B.n719 10.6151
R946 B.n721 B.n720 10.6151
R947 B.n721 B.n14 10.6151
R948 B.n725 B.n14 10.6151
R949 B.n726 B.n725 10.6151
R950 B.n727 B.n726 10.6151
R951 B.n727 B.n12 10.6151
R952 B.n731 B.n12 10.6151
R953 B.n732 B.n731 10.6151
R954 B.n733 B.n732 10.6151
R955 B.n733 B.n10 10.6151
R956 B.n737 B.n10 10.6151
R957 B.n738 B.n737 10.6151
R958 B.n739 B.n738 10.6151
R959 B.n739 B.n8 10.6151
R960 B.n743 B.n8 10.6151
R961 B.n744 B.n743 10.6151
R962 B.n745 B.n744 10.6151
R963 B.n745 B.n6 10.6151
R964 B.n749 B.n6 10.6151
R965 B.n750 B.n749 10.6151
R966 B.n751 B.n750 10.6151
R967 B.n751 B.n4 10.6151
R968 B.n755 B.n4 10.6151
R969 B.n756 B.n755 10.6151
R970 B.n757 B.n756 10.6151
R971 B.n757 B.n0 10.6151
R972 B.n695 B.n24 10.6151
R973 B.n691 B.n24 10.6151
R974 B.n691 B.n690 10.6151
R975 B.n690 B.n689 10.6151
R976 B.n689 B.n26 10.6151
R977 B.n685 B.n26 10.6151
R978 B.n685 B.n684 10.6151
R979 B.n684 B.n683 10.6151
R980 B.n683 B.n28 10.6151
R981 B.n679 B.n28 10.6151
R982 B.n679 B.n678 10.6151
R983 B.n678 B.n677 10.6151
R984 B.n677 B.n30 10.6151
R985 B.n673 B.n30 10.6151
R986 B.n673 B.n672 10.6151
R987 B.n672 B.n671 10.6151
R988 B.n671 B.n32 10.6151
R989 B.n667 B.n32 10.6151
R990 B.n667 B.n666 10.6151
R991 B.n666 B.n665 10.6151
R992 B.n665 B.n34 10.6151
R993 B.n661 B.n34 10.6151
R994 B.n661 B.n660 10.6151
R995 B.n660 B.n659 10.6151
R996 B.n659 B.n36 10.6151
R997 B.n655 B.n36 10.6151
R998 B.n655 B.n654 10.6151
R999 B.n654 B.n653 10.6151
R1000 B.n653 B.n38 10.6151
R1001 B.n649 B.n38 10.6151
R1002 B.n649 B.n648 10.6151
R1003 B.n648 B.n647 10.6151
R1004 B.n647 B.n40 10.6151
R1005 B.n643 B.n40 10.6151
R1006 B.n643 B.n642 10.6151
R1007 B.n642 B.n641 10.6151
R1008 B.n641 B.n42 10.6151
R1009 B.n637 B.n42 10.6151
R1010 B.n637 B.n636 10.6151
R1011 B.n636 B.n635 10.6151
R1012 B.n635 B.n44 10.6151
R1013 B.n631 B.n44 10.6151
R1014 B.n631 B.n630 10.6151
R1015 B.n630 B.n629 10.6151
R1016 B.n626 B.n625 10.6151
R1017 B.n625 B.n624 10.6151
R1018 B.n624 B.n50 10.6151
R1019 B.n620 B.n50 10.6151
R1020 B.n620 B.n619 10.6151
R1021 B.n619 B.n618 10.6151
R1022 B.n618 B.n52 10.6151
R1023 B.n614 B.n52 10.6151
R1024 B.n614 B.n613 10.6151
R1025 B.n611 B.n56 10.6151
R1026 B.n607 B.n56 10.6151
R1027 B.n607 B.n606 10.6151
R1028 B.n606 B.n605 10.6151
R1029 B.n605 B.n58 10.6151
R1030 B.n601 B.n58 10.6151
R1031 B.n601 B.n600 10.6151
R1032 B.n600 B.n599 10.6151
R1033 B.n599 B.n60 10.6151
R1034 B.n595 B.n60 10.6151
R1035 B.n595 B.n594 10.6151
R1036 B.n594 B.n593 10.6151
R1037 B.n593 B.n62 10.6151
R1038 B.n589 B.n62 10.6151
R1039 B.n589 B.n588 10.6151
R1040 B.n588 B.n587 10.6151
R1041 B.n587 B.n64 10.6151
R1042 B.n583 B.n64 10.6151
R1043 B.n583 B.n582 10.6151
R1044 B.n582 B.n581 10.6151
R1045 B.n581 B.n66 10.6151
R1046 B.n577 B.n66 10.6151
R1047 B.n577 B.n576 10.6151
R1048 B.n576 B.n575 10.6151
R1049 B.n575 B.n68 10.6151
R1050 B.n571 B.n68 10.6151
R1051 B.n571 B.n570 10.6151
R1052 B.n570 B.n569 10.6151
R1053 B.n569 B.n70 10.6151
R1054 B.n565 B.n70 10.6151
R1055 B.n565 B.n564 10.6151
R1056 B.n564 B.n563 10.6151
R1057 B.n563 B.n72 10.6151
R1058 B.n559 B.n72 10.6151
R1059 B.n559 B.n558 10.6151
R1060 B.n558 B.n557 10.6151
R1061 B.n557 B.n74 10.6151
R1062 B.n553 B.n74 10.6151
R1063 B.n553 B.n552 10.6151
R1064 B.n552 B.n551 10.6151
R1065 B.n551 B.n76 10.6151
R1066 B.n547 B.n76 10.6151
R1067 B.n547 B.n546 10.6151
R1068 B.n546 B.n545 10.6151
R1069 B.n541 B.n78 10.6151
R1070 B.n541 B.n540 10.6151
R1071 B.n540 B.n539 10.6151
R1072 B.n539 B.n80 10.6151
R1073 B.n535 B.n80 10.6151
R1074 B.n535 B.n534 10.6151
R1075 B.n534 B.n533 10.6151
R1076 B.n533 B.n82 10.6151
R1077 B.n529 B.n82 10.6151
R1078 B.n529 B.n528 10.6151
R1079 B.n528 B.n527 10.6151
R1080 B.n527 B.n84 10.6151
R1081 B.n523 B.n84 10.6151
R1082 B.n523 B.n522 10.6151
R1083 B.n522 B.n521 10.6151
R1084 B.n521 B.n86 10.6151
R1085 B.n517 B.n86 10.6151
R1086 B.n517 B.n516 10.6151
R1087 B.n516 B.n515 10.6151
R1088 B.n515 B.n88 10.6151
R1089 B.n511 B.n88 10.6151
R1090 B.n511 B.n510 10.6151
R1091 B.n510 B.n509 10.6151
R1092 B.n509 B.n90 10.6151
R1093 B.n505 B.n90 10.6151
R1094 B.n505 B.n504 10.6151
R1095 B.n504 B.n503 10.6151
R1096 B.n503 B.n92 10.6151
R1097 B.n499 B.n92 10.6151
R1098 B.n499 B.n498 10.6151
R1099 B.n498 B.n497 10.6151
R1100 B.n497 B.n94 10.6151
R1101 B.n493 B.n94 10.6151
R1102 B.n493 B.n492 10.6151
R1103 B.n492 B.n491 10.6151
R1104 B.n491 B.n96 10.6151
R1105 B.n487 B.n96 10.6151
R1106 B.n487 B.n486 10.6151
R1107 B.n486 B.n485 10.6151
R1108 B.n485 B.n98 10.6151
R1109 B.n481 B.n98 10.6151
R1110 B.n481 B.n480 10.6151
R1111 B.n480 B.n479 10.6151
R1112 B.n479 B.n100 10.6151
R1113 B.n475 B.n100 10.6151
R1114 B.n475 B.n474 10.6151
R1115 B.n474 B.n473 10.6151
R1116 B.n473 B.n102 10.6151
R1117 B.n469 B.n102 10.6151
R1118 B.n469 B.n468 10.6151
R1119 B.n468 B.n467 10.6151
R1120 B.n467 B.n104 10.6151
R1121 B.n463 B.n104 10.6151
R1122 B.n463 B.n462 10.6151
R1123 B.n462 B.n461 10.6151
R1124 B.n461 B.n106 10.6151
R1125 B.n457 B.n106 10.6151
R1126 B.n457 B.n456 10.6151
R1127 B.n456 B.n455 10.6151
R1128 B.n455 B.n108 10.6151
R1129 B.n451 B.n108 10.6151
R1130 B.n451 B.n450 10.6151
R1131 B.n450 B.n449 10.6151
R1132 B.n449 B.n110 10.6151
R1133 B.n445 B.n110 10.6151
R1134 B.n445 B.n444 10.6151
R1135 B.n444 B.n443 10.6151
R1136 B.n443 B.n112 10.6151
R1137 B.n439 B.n112 10.6151
R1138 B.n439 B.n438 10.6151
R1139 B.n438 B.n437 10.6151
R1140 B.n437 B.n114 10.6151
R1141 B.n433 B.n114 10.6151
R1142 B.n433 B.n432 10.6151
R1143 B.n432 B.n431 10.6151
R1144 B.n431 B.n116 10.6151
R1145 B.n427 B.n116 10.6151
R1146 B.n427 B.n426 10.6151
R1147 B.n426 B.n425 10.6151
R1148 B.n425 B.n118 10.6151
R1149 B.n421 B.n118 10.6151
R1150 B.n421 B.n420 10.6151
R1151 B.n420 B.n419 10.6151
R1152 B.n419 B.n120 10.6151
R1153 B.n415 B.n120 10.6151
R1154 B.n415 B.n414 10.6151
R1155 B.n414 B.n413 10.6151
R1156 B.n195 B.n1 10.6151
R1157 B.n195 B.n194 10.6151
R1158 B.n199 B.n194 10.6151
R1159 B.n200 B.n199 10.6151
R1160 B.n201 B.n200 10.6151
R1161 B.n201 B.n192 10.6151
R1162 B.n205 B.n192 10.6151
R1163 B.n206 B.n205 10.6151
R1164 B.n207 B.n206 10.6151
R1165 B.n207 B.n190 10.6151
R1166 B.n211 B.n190 10.6151
R1167 B.n212 B.n211 10.6151
R1168 B.n213 B.n212 10.6151
R1169 B.n213 B.n188 10.6151
R1170 B.n217 B.n188 10.6151
R1171 B.n218 B.n217 10.6151
R1172 B.n219 B.n218 10.6151
R1173 B.n219 B.n186 10.6151
R1174 B.n223 B.n186 10.6151
R1175 B.n224 B.n223 10.6151
R1176 B.n225 B.n224 10.6151
R1177 B.n225 B.n184 10.6151
R1178 B.n229 B.n184 10.6151
R1179 B.n230 B.n229 10.6151
R1180 B.n231 B.n230 10.6151
R1181 B.n231 B.n182 10.6151
R1182 B.n235 B.n182 10.6151
R1183 B.n236 B.n235 10.6151
R1184 B.n237 B.n236 10.6151
R1185 B.n237 B.n180 10.6151
R1186 B.n241 B.n180 10.6151
R1187 B.n242 B.n241 10.6151
R1188 B.n243 B.n242 10.6151
R1189 B.n243 B.n178 10.6151
R1190 B.n247 B.n178 10.6151
R1191 B.n248 B.n247 10.6151
R1192 B.n249 B.n248 10.6151
R1193 B.n249 B.n176 10.6151
R1194 B.n253 B.n176 10.6151
R1195 B.n254 B.n253 10.6151
R1196 B.n255 B.n254 10.6151
R1197 B.n255 B.n174 10.6151
R1198 B.n260 B.n259 10.6151
R1199 B.n261 B.n260 10.6151
R1200 B.n261 B.n172 10.6151
R1201 B.n265 B.n172 10.6151
R1202 B.n266 B.n265 10.6151
R1203 B.n267 B.n266 10.6151
R1204 B.n267 B.n170 10.6151
R1205 B.n271 B.n170 10.6151
R1206 B.n272 B.n271 10.6151
R1207 B.n273 B.n272 10.6151
R1208 B.n273 B.n168 10.6151
R1209 B.n277 B.n168 10.6151
R1210 B.n278 B.n277 10.6151
R1211 B.n279 B.n278 10.6151
R1212 B.n279 B.n166 10.6151
R1213 B.n283 B.n166 10.6151
R1214 B.n284 B.n283 10.6151
R1215 B.n285 B.n284 10.6151
R1216 B.n285 B.n164 10.6151
R1217 B.n289 B.n164 10.6151
R1218 B.n290 B.n289 10.6151
R1219 B.n291 B.n290 10.6151
R1220 B.n291 B.n162 10.6151
R1221 B.n295 B.n162 10.6151
R1222 B.n296 B.n295 10.6151
R1223 B.n297 B.n296 10.6151
R1224 B.n297 B.n160 10.6151
R1225 B.n301 B.n160 10.6151
R1226 B.n302 B.n301 10.6151
R1227 B.n303 B.n302 10.6151
R1228 B.n303 B.n158 10.6151
R1229 B.n307 B.n158 10.6151
R1230 B.n308 B.n307 10.6151
R1231 B.n309 B.n308 10.6151
R1232 B.n309 B.n156 10.6151
R1233 B.n313 B.n156 10.6151
R1234 B.n314 B.n313 10.6151
R1235 B.n315 B.n314 10.6151
R1236 B.n315 B.n154 10.6151
R1237 B.n319 B.n154 10.6151
R1238 B.n320 B.n319 10.6151
R1239 B.n321 B.n320 10.6151
R1240 B.n321 B.n152 10.6151
R1241 B.n325 B.n152 10.6151
R1242 B.n328 B.n327 10.6151
R1243 B.n328 B.n148 10.6151
R1244 B.n332 B.n148 10.6151
R1245 B.n333 B.n332 10.6151
R1246 B.n334 B.n333 10.6151
R1247 B.n334 B.n146 10.6151
R1248 B.n338 B.n146 10.6151
R1249 B.n339 B.n338 10.6151
R1250 B.n343 B.n339 10.6151
R1251 B.n347 B.n144 10.6151
R1252 B.n348 B.n347 10.6151
R1253 B.n349 B.n348 10.6151
R1254 B.n349 B.n142 10.6151
R1255 B.n353 B.n142 10.6151
R1256 B.n354 B.n353 10.6151
R1257 B.n355 B.n354 10.6151
R1258 B.n355 B.n140 10.6151
R1259 B.n359 B.n140 10.6151
R1260 B.n360 B.n359 10.6151
R1261 B.n361 B.n360 10.6151
R1262 B.n361 B.n138 10.6151
R1263 B.n365 B.n138 10.6151
R1264 B.n366 B.n365 10.6151
R1265 B.n367 B.n366 10.6151
R1266 B.n367 B.n136 10.6151
R1267 B.n371 B.n136 10.6151
R1268 B.n372 B.n371 10.6151
R1269 B.n373 B.n372 10.6151
R1270 B.n373 B.n134 10.6151
R1271 B.n377 B.n134 10.6151
R1272 B.n378 B.n377 10.6151
R1273 B.n379 B.n378 10.6151
R1274 B.n379 B.n132 10.6151
R1275 B.n383 B.n132 10.6151
R1276 B.n384 B.n383 10.6151
R1277 B.n385 B.n384 10.6151
R1278 B.n385 B.n130 10.6151
R1279 B.n389 B.n130 10.6151
R1280 B.n390 B.n389 10.6151
R1281 B.n391 B.n390 10.6151
R1282 B.n391 B.n128 10.6151
R1283 B.n395 B.n128 10.6151
R1284 B.n396 B.n395 10.6151
R1285 B.n397 B.n396 10.6151
R1286 B.n397 B.n126 10.6151
R1287 B.n401 B.n126 10.6151
R1288 B.n402 B.n401 10.6151
R1289 B.n403 B.n402 10.6151
R1290 B.n403 B.n124 10.6151
R1291 B.n407 B.n124 10.6151
R1292 B.n408 B.n407 10.6151
R1293 B.n409 B.n408 10.6151
R1294 B.n409 B.n122 10.6151
R1295 B.n629 B.n48 9.36635
R1296 B.n612 B.n611 9.36635
R1297 B.n326 B.n325 9.36635
R1298 B.n342 B.n144 9.36635
R1299 B.n761 B.n0 8.11757
R1300 B.n761 B.n1 8.11757
R1301 B.n626 B.n48 1.24928
R1302 B.n613 B.n612 1.24928
R1303 B.n327 B.n326 1.24928
R1304 B.n343 B.n342 1.24928
C0 VP VN 7.20708f
C1 VDD1 VDD2 1.42904f
C2 VDD1 w_n3362_n3608# 2.38567f
C3 VDD2 VTAIL 8.22317f
C4 w_n3362_n3608# VTAIL 3.13964f
C5 VP VDD2 0.463625f
C6 w_n3362_n3608# VP 6.85032f
C7 VDD2 VN 7.39496f
C8 w_n3362_n3608# VN 6.4155f
C9 VDD1 B 2.20355f
C10 B VTAIL 3.98861f
C11 w_n3362_n3608# VDD2 2.47262f
C12 VP B 1.92399f
C13 B VN 1.1977f
C14 VDD1 VTAIL 8.17214f
C15 VDD1 VP 7.70426f
C16 VP VTAIL 7.52573f
C17 VDD1 VN 0.150946f
C18 B VDD2 2.27908f
C19 w_n3362_n3608# B 10.0955f
C20 VN VTAIL 7.511431f
C21 VDD2 VSUBS 1.969963f
C22 VDD1 VSUBS 2.45717f
C23 VTAIL VSUBS 1.239996f
C24 VN VSUBS 5.93997f
C25 VP VSUBS 3.036598f
C26 B VSUBS 4.799499f
C27 w_n3362_n3608# VSUBS 0.149071p
C28 B.n0 VSUBS 0.006901f
C29 B.n1 VSUBS 0.006901f
C30 B.n2 VSUBS 0.010207f
C31 B.n3 VSUBS 0.007821f
C32 B.n4 VSUBS 0.007821f
C33 B.n5 VSUBS 0.007821f
C34 B.n6 VSUBS 0.007821f
C35 B.n7 VSUBS 0.007821f
C36 B.n8 VSUBS 0.007821f
C37 B.n9 VSUBS 0.007821f
C38 B.n10 VSUBS 0.007821f
C39 B.n11 VSUBS 0.007821f
C40 B.n12 VSUBS 0.007821f
C41 B.n13 VSUBS 0.007821f
C42 B.n14 VSUBS 0.007821f
C43 B.n15 VSUBS 0.007821f
C44 B.n16 VSUBS 0.007821f
C45 B.n17 VSUBS 0.007821f
C46 B.n18 VSUBS 0.007821f
C47 B.n19 VSUBS 0.007821f
C48 B.n20 VSUBS 0.007821f
C49 B.n21 VSUBS 0.007821f
C50 B.n22 VSUBS 0.007821f
C51 B.n23 VSUBS 0.016777f
C52 B.n24 VSUBS 0.007821f
C53 B.n25 VSUBS 0.007821f
C54 B.n26 VSUBS 0.007821f
C55 B.n27 VSUBS 0.007821f
C56 B.n28 VSUBS 0.007821f
C57 B.n29 VSUBS 0.007821f
C58 B.n30 VSUBS 0.007821f
C59 B.n31 VSUBS 0.007821f
C60 B.n32 VSUBS 0.007821f
C61 B.n33 VSUBS 0.007821f
C62 B.n34 VSUBS 0.007821f
C63 B.n35 VSUBS 0.007821f
C64 B.n36 VSUBS 0.007821f
C65 B.n37 VSUBS 0.007821f
C66 B.n38 VSUBS 0.007821f
C67 B.n39 VSUBS 0.007821f
C68 B.n40 VSUBS 0.007821f
C69 B.n41 VSUBS 0.007821f
C70 B.n42 VSUBS 0.007821f
C71 B.n43 VSUBS 0.007821f
C72 B.n44 VSUBS 0.007821f
C73 B.n45 VSUBS 0.007821f
C74 B.t4 VSUBS 0.485355f
C75 B.t5 VSUBS 0.509f
C76 B.t3 VSUBS 1.77912f
C77 B.n46 VSUBS 0.270521f
C78 B.n47 VSUBS 0.080578f
C79 B.n48 VSUBS 0.018122f
C80 B.n49 VSUBS 0.007821f
C81 B.n50 VSUBS 0.007821f
C82 B.n51 VSUBS 0.007821f
C83 B.n52 VSUBS 0.007821f
C84 B.n53 VSUBS 0.007821f
C85 B.t1 VSUBS 0.485345f
C86 B.t2 VSUBS 0.50899f
C87 B.t0 VSUBS 1.77912f
C88 B.n54 VSUBS 0.27053f
C89 B.n55 VSUBS 0.080588f
C90 B.n56 VSUBS 0.007821f
C91 B.n57 VSUBS 0.007821f
C92 B.n58 VSUBS 0.007821f
C93 B.n59 VSUBS 0.007821f
C94 B.n60 VSUBS 0.007821f
C95 B.n61 VSUBS 0.007821f
C96 B.n62 VSUBS 0.007821f
C97 B.n63 VSUBS 0.007821f
C98 B.n64 VSUBS 0.007821f
C99 B.n65 VSUBS 0.007821f
C100 B.n66 VSUBS 0.007821f
C101 B.n67 VSUBS 0.007821f
C102 B.n68 VSUBS 0.007821f
C103 B.n69 VSUBS 0.007821f
C104 B.n70 VSUBS 0.007821f
C105 B.n71 VSUBS 0.007821f
C106 B.n72 VSUBS 0.007821f
C107 B.n73 VSUBS 0.007821f
C108 B.n74 VSUBS 0.007821f
C109 B.n75 VSUBS 0.007821f
C110 B.n76 VSUBS 0.007821f
C111 B.n77 VSUBS 0.007821f
C112 B.n78 VSUBS 0.016777f
C113 B.n79 VSUBS 0.007821f
C114 B.n80 VSUBS 0.007821f
C115 B.n81 VSUBS 0.007821f
C116 B.n82 VSUBS 0.007821f
C117 B.n83 VSUBS 0.007821f
C118 B.n84 VSUBS 0.007821f
C119 B.n85 VSUBS 0.007821f
C120 B.n86 VSUBS 0.007821f
C121 B.n87 VSUBS 0.007821f
C122 B.n88 VSUBS 0.007821f
C123 B.n89 VSUBS 0.007821f
C124 B.n90 VSUBS 0.007821f
C125 B.n91 VSUBS 0.007821f
C126 B.n92 VSUBS 0.007821f
C127 B.n93 VSUBS 0.007821f
C128 B.n94 VSUBS 0.007821f
C129 B.n95 VSUBS 0.007821f
C130 B.n96 VSUBS 0.007821f
C131 B.n97 VSUBS 0.007821f
C132 B.n98 VSUBS 0.007821f
C133 B.n99 VSUBS 0.007821f
C134 B.n100 VSUBS 0.007821f
C135 B.n101 VSUBS 0.007821f
C136 B.n102 VSUBS 0.007821f
C137 B.n103 VSUBS 0.007821f
C138 B.n104 VSUBS 0.007821f
C139 B.n105 VSUBS 0.007821f
C140 B.n106 VSUBS 0.007821f
C141 B.n107 VSUBS 0.007821f
C142 B.n108 VSUBS 0.007821f
C143 B.n109 VSUBS 0.007821f
C144 B.n110 VSUBS 0.007821f
C145 B.n111 VSUBS 0.007821f
C146 B.n112 VSUBS 0.007821f
C147 B.n113 VSUBS 0.007821f
C148 B.n114 VSUBS 0.007821f
C149 B.n115 VSUBS 0.007821f
C150 B.n116 VSUBS 0.007821f
C151 B.n117 VSUBS 0.007821f
C152 B.n118 VSUBS 0.007821f
C153 B.n119 VSUBS 0.007821f
C154 B.n120 VSUBS 0.007821f
C155 B.n121 VSUBS 0.007821f
C156 B.n122 VSUBS 0.016477f
C157 B.n123 VSUBS 0.007821f
C158 B.n124 VSUBS 0.007821f
C159 B.n125 VSUBS 0.007821f
C160 B.n126 VSUBS 0.007821f
C161 B.n127 VSUBS 0.007821f
C162 B.n128 VSUBS 0.007821f
C163 B.n129 VSUBS 0.007821f
C164 B.n130 VSUBS 0.007821f
C165 B.n131 VSUBS 0.007821f
C166 B.n132 VSUBS 0.007821f
C167 B.n133 VSUBS 0.007821f
C168 B.n134 VSUBS 0.007821f
C169 B.n135 VSUBS 0.007821f
C170 B.n136 VSUBS 0.007821f
C171 B.n137 VSUBS 0.007821f
C172 B.n138 VSUBS 0.007821f
C173 B.n139 VSUBS 0.007821f
C174 B.n140 VSUBS 0.007821f
C175 B.n141 VSUBS 0.007821f
C176 B.n142 VSUBS 0.007821f
C177 B.n143 VSUBS 0.007821f
C178 B.n144 VSUBS 0.007361f
C179 B.n145 VSUBS 0.007821f
C180 B.n146 VSUBS 0.007821f
C181 B.n147 VSUBS 0.007821f
C182 B.n148 VSUBS 0.007821f
C183 B.n149 VSUBS 0.007821f
C184 B.t11 VSUBS 0.485355f
C185 B.t10 VSUBS 0.509f
C186 B.t9 VSUBS 1.77912f
C187 B.n150 VSUBS 0.270521f
C188 B.n151 VSUBS 0.080578f
C189 B.n152 VSUBS 0.007821f
C190 B.n153 VSUBS 0.007821f
C191 B.n154 VSUBS 0.007821f
C192 B.n155 VSUBS 0.007821f
C193 B.n156 VSUBS 0.007821f
C194 B.n157 VSUBS 0.007821f
C195 B.n158 VSUBS 0.007821f
C196 B.n159 VSUBS 0.007821f
C197 B.n160 VSUBS 0.007821f
C198 B.n161 VSUBS 0.007821f
C199 B.n162 VSUBS 0.007821f
C200 B.n163 VSUBS 0.007821f
C201 B.n164 VSUBS 0.007821f
C202 B.n165 VSUBS 0.007821f
C203 B.n166 VSUBS 0.007821f
C204 B.n167 VSUBS 0.007821f
C205 B.n168 VSUBS 0.007821f
C206 B.n169 VSUBS 0.007821f
C207 B.n170 VSUBS 0.007821f
C208 B.n171 VSUBS 0.007821f
C209 B.n172 VSUBS 0.007821f
C210 B.n173 VSUBS 0.007821f
C211 B.n174 VSUBS 0.016777f
C212 B.n175 VSUBS 0.007821f
C213 B.n176 VSUBS 0.007821f
C214 B.n177 VSUBS 0.007821f
C215 B.n178 VSUBS 0.007821f
C216 B.n179 VSUBS 0.007821f
C217 B.n180 VSUBS 0.007821f
C218 B.n181 VSUBS 0.007821f
C219 B.n182 VSUBS 0.007821f
C220 B.n183 VSUBS 0.007821f
C221 B.n184 VSUBS 0.007821f
C222 B.n185 VSUBS 0.007821f
C223 B.n186 VSUBS 0.007821f
C224 B.n187 VSUBS 0.007821f
C225 B.n188 VSUBS 0.007821f
C226 B.n189 VSUBS 0.007821f
C227 B.n190 VSUBS 0.007821f
C228 B.n191 VSUBS 0.007821f
C229 B.n192 VSUBS 0.007821f
C230 B.n193 VSUBS 0.007821f
C231 B.n194 VSUBS 0.007821f
C232 B.n195 VSUBS 0.007821f
C233 B.n196 VSUBS 0.007821f
C234 B.n197 VSUBS 0.007821f
C235 B.n198 VSUBS 0.007821f
C236 B.n199 VSUBS 0.007821f
C237 B.n200 VSUBS 0.007821f
C238 B.n201 VSUBS 0.007821f
C239 B.n202 VSUBS 0.007821f
C240 B.n203 VSUBS 0.007821f
C241 B.n204 VSUBS 0.007821f
C242 B.n205 VSUBS 0.007821f
C243 B.n206 VSUBS 0.007821f
C244 B.n207 VSUBS 0.007821f
C245 B.n208 VSUBS 0.007821f
C246 B.n209 VSUBS 0.007821f
C247 B.n210 VSUBS 0.007821f
C248 B.n211 VSUBS 0.007821f
C249 B.n212 VSUBS 0.007821f
C250 B.n213 VSUBS 0.007821f
C251 B.n214 VSUBS 0.007821f
C252 B.n215 VSUBS 0.007821f
C253 B.n216 VSUBS 0.007821f
C254 B.n217 VSUBS 0.007821f
C255 B.n218 VSUBS 0.007821f
C256 B.n219 VSUBS 0.007821f
C257 B.n220 VSUBS 0.007821f
C258 B.n221 VSUBS 0.007821f
C259 B.n222 VSUBS 0.007821f
C260 B.n223 VSUBS 0.007821f
C261 B.n224 VSUBS 0.007821f
C262 B.n225 VSUBS 0.007821f
C263 B.n226 VSUBS 0.007821f
C264 B.n227 VSUBS 0.007821f
C265 B.n228 VSUBS 0.007821f
C266 B.n229 VSUBS 0.007821f
C267 B.n230 VSUBS 0.007821f
C268 B.n231 VSUBS 0.007821f
C269 B.n232 VSUBS 0.007821f
C270 B.n233 VSUBS 0.007821f
C271 B.n234 VSUBS 0.007821f
C272 B.n235 VSUBS 0.007821f
C273 B.n236 VSUBS 0.007821f
C274 B.n237 VSUBS 0.007821f
C275 B.n238 VSUBS 0.007821f
C276 B.n239 VSUBS 0.007821f
C277 B.n240 VSUBS 0.007821f
C278 B.n241 VSUBS 0.007821f
C279 B.n242 VSUBS 0.007821f
C280 B.n243 VSUBS 0.007821f
C281 B.n244 VSUBS 0.007821f
C282 B.n245 VSUBS 0.007821f
C283 B.n246 VSUBS 0.007821f
C284 B.n247 VSUBS 0.007821f
C285 B.n248 VSUBS 0.007821f
C286 B.n249 VSUBS 0.007821f
C287 B.n250 VSUBS 0.007821f
C288 B.n251 VSUBS 0.007821f
C289 B.n252 VSUBS 0.007821f
C290 B.n253 VSUBS 0.007821f
C291 B.n254 VSUBS 0.007821f
C292 B.n255 VSUBS 0.007821f
C293 B.n256 VSUBS 0.007821f
C294 B.n257 VSUBS 0.016777f
C295 B.n258 VSUBS 0.0175f
C296 B.n259 VSUBS 0.0175f
C297 B.n260 VSUBS 0.007821f
C298 B.n261 VSUBS 0.007821f
C299 B.n262 VSUBS 0.007821f
C300 B.n263 VSUBS 0.007821f
C301 B.n264 VSUBS 0.007821f
C302 B.n265 VSUBS 0.007821f
C303 B.n266 VSUBS 0.007821f
C304 B.n267 VSUBS 0.007821f
C305 B.n268 VSUBS 0.007821f
C306 B.n269 VSUBS 0.007821f
C307 B.n270 VSUBS 0.007821f
C308 B.n271 VSUBS 0.007821f
C309 B.n272 VSUBS 0.007821f
C310 B.n273 VSUBS 0.007821f
C311 B.n274 VSUBS 0.007821f
C312 B.n275 VSUBS 0.007821f
C313 B.n276 VSUBS 0.007821f
C314 B.n277 VSUBS 0.007821f
C315 B.n278 VSUBS 0.007821f
C316 B.n279 VSUBS 0.007821f
C317 B.n280 VSUBS 0.007821f
C318 B.n281 VSUBS 0.007821f
C319 B.n282 VSUBS 0.007821f
C320 B.n283 VSUBS 0.007821f
C321 B.n284 VSUBS 0.007821f
C322 B.n285 VSUBS 0.007821f
C323 B.n286 VSUBS 0.007821f
C324 B.n287 VSUBS 0.007821f
C325 B.n288 VSUBS 0.007821f
C326 B.n289 VSUBS 0.007821f
C327 B.n290 VSUBS 0.007821f
C328 B.n291 VSUBS 0.007821f
C329 B.n292 VSUBS 0.007821f
C330 B.n293 VSUBS 0.007821f
C331 B.n294 VSUBS 0.007821f
C332 B.n295 VSUBS 0.007821f
C333 B.n296 VSUBS 0.007821f
C334 B.n297 VSUBS 0.007821f
C335 B.n298 VSUBS 0.007821f
C336 B.n299 VSUBS 0.007821f
C337 B.n300 VSUBS 0.007821f
C338 B.n301 VSUBS 0.007821f
C339 B.n302 VSUBS 0.007821f
C340 B.n303 VSUBS 0.007821f
C341 B.n304 VSUBS 0.007821f
C342 B.n305 VSUBS 0.007821f
C343 B.n306 VSUBS 0.007821f
C344 B.n307 VSUBS 0.007821f
C345 B.n308 VSUBS 0.007821f
C346 B.n309 VSUBS 0.007821f
C347 B.n310 VSUBS 0.007821f
C348 B.n311 VSUBS 0.007821f
C349 B.n312 VSUBS 0.007821f
C350 B.n313 VSUBS 0.007821f
C351 B.n314 VSUBS 0.007821f
C352 B.n315 VSUBS 0.007821f
C353 B.n316 VSUBS 0.007821f
C354 B.n317 VSUBS 0.007821f
C355 B.n318 VSUBS 0.007821f
C356 B.n319 VSUBS 0.007821f
C357 B.n320 VSUBS 0.007821f
C358 B.n321 VSUBS 0.007821f
C359 B.n322 VSUBS 0.007821f
C360 B.n323 VSUBS 0.007821f
C361 B.n324 VSUBS 0.007821f
C362 B.n325 VSUBS 0.007361f
C363 B.n326 VSUBS 0.018122f
C364 B.n327 VSUBS 0.004371f
C365 B.n328 VSUBS 0.007821f
C366 B.n329 VSUBS 0.007821f
C367 B.n330 VSUBS 0.007821f
C368 B.n331 VSUBS 0.007821f
C369 B.n332 VSUBS 0.007821f
C370 B.n333 VSUBS 0.007821f
C371 B.n334 VSUBS 0.007821f
C372 B.n335 VSUBS 0.007821f
C373 B.n336 VSUBS 0.007821f
C374 B.n337 VSUBS 0.007821f
C375 B.n338 VSUBS 0.007821f
C376 B.n339 VSUBS 0.007821f
C377 B.t8 VSUBS 0.485345f
C378 B.t7 VSUBS 0.50899f
C379 B.t6 VSUBS 1.77912f
C380 B.n340 VSUBS 0.27053f
C381 B.n341 VSUBS 0.080588f
C382 B.n342 VSUBS 0.018122f
C383 B.n343 VSUBS 0.004371f
C384 B.n344 VSUBS 0.007821f
C385 B.n345 VSUBS 0.007821f
C386 B.n346 VSUBS 0.007821f
C387 B.n347 VSUBS 0.007821f
C388 B.n348 VSUBS 0.007821f
C389 B.n349 VSUBS 0.007821f
C390 B.n350 VSUBS 0.007821f
C391 B.n351 VSUBS 0.007821f
C392 B.n352 VSUBS 0.007821f
C393 B.n353 VSUBS 0.007821f
C394 B.n354 VSUBS 0.007821f
C395 B.n355 VSUBS 0.007821f
C396 B.n356 VSUBS 0.007821f
C397 B.n357 VSUBS 0.007821f
C398 B.n358 VSUBS 0.007821f
C399 B.n359 VSUBS 0.007821f
C400 B.n360 VSUBS 0.007821f
C401 B.n361 VSUBS 0.007821f
C402 B.n362 VSUBS 0.007821f
C403 B.n363 VSUBS 0.007821f
C404 B.n364 VSUBS 0.007821f
C405 B.n365 VSUBS 0.007821f
C406 B.n366 VSUBS 0.007821f
C407 B.n367 VSUBS 0.007821f
C408 B.n368 VSUBS 0.007821f
C409 B.n369 VSUBS 0.007821f
C410 B.n370 VSUBS 0.007821f
C411 B.n371 VSUBS 0.007821f
C412 B.n372 VSUBS 0.007821f
C413 B.n373 VSUBS 0.007821f
C414 B.n374 VSUBS 0.007821f
C415 B.n375 VSUBS 0.007821f
C416 B.n376 VSUBS 0.007821f
C417 B.n377 VSUBS 0.007821f
C418 B.n378 VSUBS 0.007821f
C419 B.n379 VSUBS 0.007821f
C420 B.n380 VSUBS 0.007821f
C421 B.n381 VSUBS 0.007821f
C422 B.n382 VSUBS 0.007821f
C423 B.n383 VSUBS 0.007821f
C424 B.n384 VSUBS 0.007821f
C425 B.n385 VSUBS 0.007821f
C426 B.n386 VSUBS 0.007821f
C427 B.n387 VSUBS 0.007821f
C428 B.n388 VSUBS 0.007821f
C429 B.n389 VSUBS 0.007821f
C430 B.n390 VSUBS 0.007821f
C431 B.n391 VSUBS 0.007821f
C432 B.n392 VSUBS 0.007821f
C433 B.n393 VSUBS 0.007821f
C434 B.n394 VSUBS 0.007821f
C435 B.n395 VSUBS 0.007821f
C436 B.n396 VSUBS 0.007821f
C437 B.n397 VSUBS 0.007821f
C438 B.n398 VSUBS 0.007821f
C439 B.n399 VSUBS 0.007821f
C440 B.n400 VSUBS 0.007821f
C441 B.n401 VSUBS 0.007821f
C442 B.n402 VSUBS 0.007821f
C443 B.n403 VSUBS 0.007821f
C444 B.n404 VSUBS 0.007821f
C445 B.n405 VSUBS 0.007821f
C446 B.n406 VSUBS 0.007821f
C447 B.n407 VSUBS 0.007821f
C448 B.n408 VSUBS 0.007821f
C449 B.n409 VSUBS 0.007821f
C450 B.n410 VSUBS 0.007821f
C451 B.n411 VSUBS 0.0175f
C452 B.n412 VSUBS 0.016777f
C453 B.n413 VSUBS 0.017799f
C454 B.n414 VSUBS 0.007821f
C455 B.n415 VSUBS 0.007821f
C456 B.n416 VSUBS 0.007821f
C457 B.n417 VSUBS 0.007821f
C458 B.n418 VSUBS 0.007821f
C459 B.n419 VSUBS 0.007821f
C460 B.n420 VSUBS 0.007821f
C461 B.n421 VSUBS 0.007821f
C462 B.n422 VSUBS 0.007821f
C463 B.n423 VSUBS 0.007821f
C464 B.n424 VSUBS 0.007821f
C465 B.n425 VSUBS 0.007821f
C466 B.n426 VSUBS 0.007821f
C467 B.n427 VSUBS 0.007821f
C468 B.n428 VSUBS 0.007821f
C469 B.n429 VSUBS 0.007821f
C470 B.n430 VSUBS 0.007821f
C471 B.n431 VSUBS 0.007821f
C472 B.n432 VSUBS 0.007821f
C473 B.n433 VSUBS 0.007821f
C474 B.n434 VSUBS 0.007821f
C475 B.n435 VSUBS 0.007821f
C476 B.n436 VSUBS 0.007821f
C477 B.n437 VSUBS 0.007821f
C478 B.n438 VSUBS 0.007821f
C479 B.n439 VSUBS 0.007821f
C480 B.n440 VSUBS 0.007821f
C481 B.n441 VSUBS 0.007821f
C482 B.n442 VSUBS 0.007821f
C483 B.n443 VSUBS 0.007821f
C484 B.n444 VSUBS 0.007821f
C485 B.n445 VSUBS 0.007821f
C486 B.n446 VSUBS 0.007821f
C487 B.n447 VSUBS 0.007821f
C488 B.n448 VSUBS 0.007821f
C489 B.n449 VSUBS 0.007821f
C490 B.n450 VSUBS 0.007821f
C491 B.n451 VSUBS 0.007821f
C492 B.n452 VSUBS 0.007821f
C493 B.n453 VSUBS 0.007821f
C494 B.n454 VSUBS 0.007821f
C495 B.n455 VSUBS 0.007821f
C496 B.n456 VSUBS 0.007821f
C497 B.n457 VSUBS 0.007821f
C498 B.n458 VSUBS 0.007821f
C499 B.n459 VSUBS 0.007821f
C500 B.n460 VSUBS 0.007821f
C501 B.n461 VSUBS 0.007821f
C502 B.n462 VSUBS 0.007821f
C503 B.n463 VSUBS 0.007821f
C504 B.n464 VSUBS 0.007821f
C505 B.n465 VSUBS 0.007821f
C506 B.n466 VSUBS 0.007821f
C507 B.n467 VSUBS 0.007821f
C508 B.n468 VSUBS 0.007821f
C509 B.n469 VSUBS 0.007821f
C510 B.n470 VSUBS 0.007821f
C511 B.n471 VSUBS 0.007821f
C512 B.n472 VSUBS 0.007821f
C513 B.n473 VSUBS 0.007821f
C514 B.n474 VSUBS 0.007821f
C515 B.n475 VSUBS 0.007821f
C516 B.n476 VSUBS 0.007821f
C517 B.n477 VSUBS 0.007821f
C518 B.n478 VSUBS 0.007821f
C519 B.n479 VSUBS 0.007821f
C520 B.n480 VSUBS 0.007821f
C521 B.n481 VSUBS 0.007821f
C522 B.n482 VSUBS 0.007821f
C523 B.n483 VSUBS 0.007821f
C524 B.n484 VSUBS 0.007821f
C525 B.n485 VSUBS 0.007821f
C526 B.n486 VSUBS 0.007821f
C527 B.n487 VSUBS 0.007821f
C528 B.n488 VSUBS 0.007821f
C529 B.n489 VSUBS 0.007821f
C530 B.n490 VSUBS 0.007821f
C531 B.n491 VSUBS 0.007821f
C532 B.n492 VSUBS 0.007821f
C533 B.n493 VSUBS 0.007821f
C534 B.n494 VSUBS 0.007821f
C535 B.n495 VSUBS 0.007821f
C536 B.n496 VSUBS 0.007821f
C537 B.n497 VSUBS 0.007821f
C538 B.n498 VSUBS 0.007821f
C539 B.n499 VSUBS 0.007821f
C540 B.n500 VSUBS 0.007821f
C541 B.n501 VSUBS 0.007821f
C542 B.n502 VSUBS 0.007821f
C543 B.n503 VSUBS 0.007821f
C544 B.n504 VSUBS 0.007821f
C545 B.n505 VSUBS 0.007821f
C546 B.n506 VSUBS 0.007821f
C547 B.n507 VSUBS 0.007821f
C548 B.n508 VSUBS 0.007821f
C549 B.n509 VSUBS 0.007821f
C550 B.n510 VSUBS 0.007821f
C551 B.n511 VSUBS 0.007821f
C552 B.n512 VSUBS 0.007821f
C553 B.n513 VSUBS 0.007821f
C554 B.n514 VSUBS 0.007821f
C555 B.n515 VSUBS 0.007821f
C556 B.n516 VSUBS 0.007821f
C557 B.n517 VSUBS 0.007821f
C558 B.n518 VSUBS 0.007821f
C559 B.n519 VSUBS 0.007821f
C560 B.n520 VSUBS 0.007821f
C561 B.n521 VSUBS 0.007821f
C562 B.n522 VSUBS 0.007821f
C563 B.n523 VSUBS 0.007821f
C564 B.n524 VSUBS 0.007821f
C565 B.n525 VSUBS 0.007821f
C566 B.n526 VSUBS 0.007821f
C567 B.n527 VSUBS 0.007821f
C568 B.n528 VSUBS 0.007821f
C569 B.n529 VSUBS 0.007821f
C570 B.n530 VSUBS 0.007821f
C571 B.n531 VSUBS 0.007821f
C572 B.n532 VSUBS 0.007821f
C573 B.n533 VSUBS 0.007821f
C574 B.n534 VSUBS 0.007821f
C575 B.n535 VSUBS 0.007821f
C576 B.n536 VSUBS 0.007821f
C577 B.n537 VSUBS 0.007821f
C578 B.n538 VSUBS 0.007821f
C579 B.n539 VSUBS 0.007821f
C580 B.n540 VSUBS 0.007821f
C581 B.n541 VSUBS 0.007821f
C582 B.n542 VSUBS 0.007821f
C583 B.n543 VSUBS 0.016777f
C584 B.n544 VSUBS 0.0175f
C585 B.n545 VSUBS 0.0175f
C586 B.n546 VSUBS 0.007821f
C587 B.n547 VSUBS 0.007821f
C588 B.n548 VSUBS 0.007821f
C589 B.n549 VSUBS 0.007821f
C590 B.n550 VSUBS 0.007821f
C591 B.n551 VSUBS 0.007821f
C592 B.n552 VSUBS 0.007821f
C593 B.n553 VSUBS 0.007821f
C594 B.n554 VSUBS 0.007821f
C595 B.n555 VSUBS 0.007821f
C596 B.n556 VSUBS 0.007821f
C597 B.n557 VSUBS 0.007821f
C598 B.n558 VSUBS 0.007821f
C599 B.n559 VSUBS 0.007821f
C600 B.n560 VSUBS 0.007821f
C601 B.n561 VSUBS 0.007821f
C602 B.n562 VSUBS 0.007821f
C603 B.n563 VSUBS 0.007821f
C604 B.n564 VSUBS 0.007821f
C605 B.n565 VSUBS 0.007821f
C606 B.n566 VSUBS 0.007821f
C607 B.n567 VSUBS 0.007821f
C608 B.n568 VSUBS 0.007821f
C609 B.n569 VSUBS 0.007821f
C610 B.n570 VSUBS 0.007821f
C611 B.n571 VSUBS 0.007821f
C612 B.n572 VSUBS 0.007821f
C613 B.n573 VSUBS 0.007821f
C614 B.n574 VSUBS 0.007821f
C615 B.n575 VSUBS 0.007821f
C616 B.n576 VSUBS 0.007821f
C617 B.n577 VSUBS 0.007821f
C618 B.n578 VSUBS 0.007821f
C619 B.n579 VSUBS 0.007821f
C620 B.n580 VSUBS 0.007821f
C621 B.n581 VSUBS 0.007821f
C622 B.n582 VSUBS 0.007821f
C623 B.n583 VSUBS 0.007821f
C624 B.n584 VSUBS 0.007821f
C625 B.n585 VSUBS 0.007821f
C626 B.n586 VSUBS 0.007821f
C627 B.n587 VSUBS 0.007821f
C628 B.n588 VSUBS 0.007821f
C629 B.n589 VSUBS 0.007821f
C630 B.n590 VSUBS 0.007821f
C631 B.n591 VSUBS 0.007821f
C632 B.n592 VSUBS 0.007821f
C633 B.n593 VSUBS 0.007821f
C634 B.n594 VSUBS 0.007821f
C635 B.n595 VSUBS 0.007821f
C636 B.n596 VSUBS 0.007821f
C637 B.n597 VSUBS 0.007821f
C638 B.n598 VSUBS 0.007821f
C639 B.n599 VSUBS 0.007821f
C640 B.n600 VSUBS 0.007821f
C641 B.n601 VSUBS 0.007821f
C642 B.n602 VSUBS 0.007821f
C643 B.n603 VSUBS 0.007821f
C644 B.n604 VSUBS 0.007821f
C645 B.n605 VSUBS 0.007821f
C646 B.n606 VSUBS 0.007821f
C647 B.n607 VSUBS 0.007821f
C648 B.n608 VSUBS 0.007821f
C649 B.n609 VSUBS 0.007821f
C650 B.n610 VSUBS 0.007821f
C651 B.n611 VSUBS 0.007361f
C652 B.n612 VSUBS 0.018122f
C653 B.n613 VSUBS 0.004371f
C654 B.n614 VSUBS 0.007821f
C655 B.n615 VSUBS 0.007821f
C656 B.n616 VSUBS 0.007821f
C657 B.n617 VSUBS 0.007821f
C658 B.n618 VSUBS 0.007821f
C659 B.n619 VSUBS 0.007821f
C660 B.n620 VSUBS 0.007821f
C661 B.n621 VSUBS 0.007821f
C662 B.n622 VSUBS 0.007821f
C663 B.n623 VSUBS 0.007821f
C664 B.n624 VSUBS 0.007821f
C665 B.n625 VSUBS 0.007821f
C666 B.n626 VSUBS 0.004371f
C667 B.n627 VSUBS 0.007821f
C668 B.n628 VSUBS 0.007821f
C669 B.n629 VSUBS 0.007361f
C670 B.n630 VSUBS 0.007821f
C671 B.n631 VSUBS 0.007821f
C672 B.n632 VSUBS 0.007821f
C673 B.n633 VSUBS 0.007821f
C674 B.n634 VSUBS 0.007821f
C675 B.n635 VSUBS 0.007821f
C676 B.n636 VSUBS 0.007821f
C677 B.n637 VSUBS 0.007821f
C678 B.n638 VSUBS 0.007821f
C679 B.n639 VSUBS 0.007821f
C680 B.n640 VSUBS 0.007821f
C681 B.n641 VSUBS 0.007821f
C682 B.n642 VSUBS 0.007821f
C683 B.n643 VSUBS 0.007821f
C684 B.n644 VSUBS 0.007821f
C685 B.n645 VSUBS 0.007821f
C686 B.n646 VSUBS 0.007821f
C687 B.n647 VSUBS 0.007821f
C688 B.n648 VSUBS 0.007821f
C689 B.n649 VSUBS 0.007821f
C690 B.n650 VSUBS 0.007821f
C691 B.n651 VSUBS 0.007821f
C692 B.n652 VSUBS 0.007821f
C693 B.n653 VSUBS 0.007821f
C694 B.n654 VSUBS 0.007821f
C695 B.n655 VSUBS 0.007821f
C696 B.n656 VSUBS 0.007821f
C697 B.n657 VSUBS 0.007821f
C698 B.n658 VSUBS 0.007821f
C699 B.n659 VSUBS 0.007821f
C700 B.n660 VSUBS 0.007821f
C701 B.n661 VSUBS 0.007821f
C702 B.n662 VSUBS 0.007821f
C703 B.n663 VSUBS 0.007821f
C704 B.n664 VSUBS 0.007821f
C705 B.n665 VSUBS 0.007821f
C706 B.n666 VSUBS 0.007821f
C707 B.n667 VSUBS 0.007821f
C708 B.n668 VSUBS 0.007821f
C709 B.n669 VSUBS 0.007821f
C710 B.n670 VSUBS 0.007821f
C711 B.n671 VSUBS 0.007821f
C712 B.n672 VSUBS 0.007821f
C713 B.n673 VSUBS 0.007821f
C714 B.n674 VSUBS 0.007821f
C715 B.n675 VSUBS 0.007821f
C716 B.n676 VSUBS 0.007821f
C717 B.n677 VSUBS 0.007821f
C718 B.n678 VSUBS 0.007821f
C719 B.n679 VSUBS 0.007821f
C720 B.n680 VSUBS 0.007821f
C721 B.n681 VSUBS 0.007821f
C722 B.n682 VSUBS 0.007821f
C723 B.n683 VSUBS 0.007821f
C724 B.n684 VSUBS 0.007821f
C725 B.n685 VSUBS 0.007821f
C726 B.n686 VSUBS 0.007821f
C727 B.n687 VSUBS 0.007821f
C728 B.n688 VSUBS 0.007821f
C729 B.n689 VSUBS 0.007821f
C730 B.n690 VSUBS 0.007821f
C731 B.n691 VSUBS 0.007821f
C732 B.n692 VSUBS 0.007821f
C733 B.n693 VSUBS 0.007821f
C734 B.n694 VSUBS 0.0175f
C735 B.n695 VSUBS 0.0175f
C736 B.n696 VSUBS 0.016777f
C737 B.n697 VSUBS 0.007821f
C738 B.n698 VSUBS 0.007821f
C739 B.n699 VSUBS 0.007821f
C740 B.n700 VSUBS 0.007821f
C741 B.n701 VSUBS 0.007821f
C742 B.n702 VSUBS 0.007821f
C743 B.n703 VSUBS 0.007821f
C744 B.n704 VSUBS 0.007821f
C745 B.n705 VSUBS 0.007821f
C746 B.n706 VSUBS 0.007821f
C747 B.n707 VSUBS 0.007821f
C748 B.n708 VSUBS 0.007821f
C749 B.n709 VSUBS 0.007821f
C750 B.n710 VSUBS 0.007821f
C751 B.n711 VSUBS 0.007821f
C752 B.n712 VSUBS 0.007821f
C753 B.n713 VSUBS 0.007821f
C754 B.n714 VSUBS 0.007821f
C755 B.n715 VSUBS 0.007821f
C756 B.n716 VSUBS 0.007821f
C757 B.n717 VSUBS 0.007821f
C758 B.n718 VSUBS 0.007821f
C759 B.n719 VSUBS 0.007821f
C760 B.n720 VSUBS 0.007821f
C761 B.n721 VSUBS 0.007821f
C762 B.n722 VSUBS 0.007821f
C763 B.n723 VSUBS 0.007821f
C764 B.n724 VSUBS 0.007821f
C765 B.n725 VSUBS 0.007821f
C766 B.n726 VSUBS 0.007821f
C767 B.n727 VSUBS 0.007821f
C768 B.n728 VSUBS 0.007821f
C769 B.n729 VSUBS 0.007821f
C770 B.n730 VSUBS 0.007821f
C771 B.n731 VSUBS 0.007821f
C772 B.n732 VSUBS 0.007821f
C773 B.n733 VSUBS 0.007821f
C774 B.n734 VSUBS 0.007821f
C775 B.n735 VSUBS 0.007821f
C776 B.n736 VSUBS 0.007821f
C777 B.n737 VSUBS 0.007821f
C778 B.n738 VSUBS 0.007821f
C779 B.n739 VSUBS 0.007821f
C780 B.n740 VSUBS 0.007821f
C781 B.n741 VSUBS 0.007821f
C782 B.n742 VSUBS 0.007821f
C783 B.n743 VSUBS 0.007821f
C784 B.n744 VSUBS 0.007821f
C785 B.n745 VSUBS 0.007821f
C786 B.n746 VSUBS 0.007821f
C787 B.n747 VSUBS 0.007821f
C788 B.n748 VSUBS 0.007821f
C789 B.n749 VSUBS 0.007821f
C790 B.n750 VSUBS 0.007821f
C791 B.n751 VSUBS 0.007821f
C792 B.n752 VSUBS 0.007821f
C793 B.n753 VSUBS 0.007821f
C794 B.n754 VSUBS 0.007821f
C795 B.n755 VSUBS 0.007821f
C796 B.n756 VSUBS 0.007821f
C797 B.n757 VSUBS 0.007821f
C798 B.n758 VSUBS 0.007821f
C799 B.n759 VSUBS 0.010207f
C800 B.n760 VSUBS 0.010873f
C801 B.n761 VSUBS 0.021621f
C802 VDD2.t5 VSUBS 3.02467f
C803 VDD2.t4 VSUBS 0.290764f
C804 VDD2.t0 VSUBS 0.290764f
C805 VDD2.n0 VSUBS 2.31072f
C806 VDD2.n1 VSUBS 3.97164f
C807 VDD2.t3 VSUBS 3.00502f
C808 VDD2.n2 VSUBS 3.56039f
C809 VDD2.t2 VSUBS 0.290764f
C810 VDD2.t1 VSUBS 0.290764f
C811 VDD2.n3 VSUBS 2.31067f
C812 VN.t5 VSUBS 2.80503f
C813 VN.n0 VSUBS 1.09706f
C814 VN.n1 VSUBS 0.029245f
C815 VN.n2 VSUBS 0.057668f
C816 VN.t0 VSUBS 3.05387f
C817 VN.n3 VSUBS 1.0463f
C818 VN.t1 VSUBS 2.80503f
C819 VN.n4 VSUBS 1.08799f
C820 VN.n5 VSUBS 0.054232f
C821 VN.n6 VSUBS 0.302455f
C822 VN.n7 VSUBS 0.029245f
C823 VN.n8 VSUBS 0.029245f
C824 VN.n9 VSUBS 0.023629f
C825 VN.n10 VSUBS 0.057958f
C826 VN.n11 VSUBS 0.053696f
C827 VN.n12 VSUBS 0.047193f
C828 VN.n13 VSUBS 0.05251f
C829 VN.t2 VSUBS 2.80503f
C830 VN.n14 VSUBS 1.09706f
C831 VN.n15 VSUBS 0.029245f
C832 VN.n16 VSUBS 0.057668f
C833 VN.t4 VSUBS 3.05387f
C834 VN.n17 VSUBS 1.0463f
C835 VN.t3 VSUBS 2.80503f
C836 VN.n18 VSUBS 1.08799f
C837 VN.n19 VSUBS 0.054232f
C838 VN.n20 VSUBS 0.302455f
C839 VN.n21 VSUBS 0.029245f
C840 VN.n22 VSUBS 0.029245f
C841 VN.n23 VSUBS 0.023629f
C842 VN.n24 VSUBS 0.057958f
C843 VN.n25 VSUBS 0.053696f
C844 VN.n26 VSUBS 0.047193f
C845 VN.n27 VSUBS 1.65101f
C846 VDD1.t3 VSUBS 3.02565f
C847 VDD1.t0 VSUBS 3.02424f
C848 VDD1.t1 VSUBS 0.290722f
C849 VDD1.t2 VSUBS 0.290722f
C850 VDD1.n0 VSUBS 2.31039f
C851 VDD1.n1 VSUBS 4.11221f
C852 VDD1.t4 VSUBS 0.290722f
C853 VDD1.t5 VSUBS 0.290722f
C854 VDD1.n2 VSUBS 2.30371f
C855 VDD1.n3 VSUBS 3.53497f
C856 VTAIL.t1 VSUBS 0.299543f
C857 VTAIL.t5 VSUBS 0.299543f
C858 VTAIL.n0 VSUBS 2.2114f
C859 VTAIL.n1 VSUBS 0.900565f
C860 VTAIL.t9 VSUBS 2.91331f
C861 VTAIL.n2 VSUBS 1.18909f
C862 VTAIL.t10 VSUBS 0.299543f
C863 VTAIL.t11 VSUBS 0.299543f
C864 VTAIL.n3 VSUBS 2.2114f
C865 VTAIL.n4 VSUBS 2.83136f
C866 VTAIL.t2 VSUBS 0.299543f
C867 VTAIL.t3 VSUBS 0.299543f
C868 VTAIL.n5 VSUBS 2.21141f
C869 VTAIL.n6 VSUBS 2.83136f
C870 VTAIL.t4 VSUBS 2.91332f
C871 VTAIL.n7 VSUBS 1.18908f
C872 VTAIL.t6 VSUBS 0.299543f
C873 VTAIL.t7 VSUBS 0.299543f
C874 VTAIL.n8 VSUBS 2.21141f
C875 VTAIL.n9 VSUBS 1.07406f
C876 VTAIL.t8 VSUBS 2.91331f
C877 VTAIL.n10 VSUBS 2.70789f
C878 VTAIL.t0 VSUBS 2.91331f
C879 VTAIL.n11 VSUBS 2.64288f
C880 VP.t3 VSUBS 2.88794f
C881 VP.n0 VSUBS 1.12949f
C882 VP.n1 VSUBS 0.030109f
C883 VP.n2 VSUBS 0.059373f
C884 VP.n3 VSUBS 0.030109f
C885 VP.t4 VSUBS 2.88794f
C886 VP.n4 VSUBS 0.059373f
C887 VP.n5 VSUBS 0.030109f
C888 VP.t5 VSUBS 2.88794f
C889 VP.n6 VSUBS 1.12949f
C890 VP.t0 VSUBS 2.88794f
C891 VP.n7 VSUBS 1.12949f
C892 VP.n8 VSUBS 0.030109f
C893 VP.n9 VSUBS 0.059373f
C894 VP.t2 VSUBS 3.14413f
C895 VP.n10 VSUBS 1.07722f
C896 VP.t1 VSUBS 2.88794f
C897 VP.n11 VSUBS 1.12015f
C898 VP.n12 VSUBS 0.055835f
C899 VP.n13 VSUBS 0.311395f
C900 VP.n14 VSUBS 0.030109f
C901 VP.n15 VSUBS 0.030109f
C902 VP.n16 VSUBS 0.024328f
C903 VP.n17 VSUBS 0.059671f
C904 VP.n18 VSUBS 0.055283f
C905 VP.n19 VSUBS 0.048588f
C906 VP.n20 VSUBS 1.68747f
C907 VP.n21 VSUBS 1.70921f
C908 VP.n22 VSUBS 0.048588f
C909 VP.n23 VSUBS 0.055283f
C910 VP.n24 VSUBS 0.059671f
C911 VP.n25 VSUBS 0.024328f
C912 VP.n26 VSUBS 0.030109f
C913 VP.n27 VSUBS 0.030109f
C914 VP.n28 VSUBS 0.030109f
C915 VP.n29 VSUBS 0.055835f
C916 VP.n30 VSUBS 1.04342f
C917 VP.n31 VSUBS 0.055835f
C918 VP.n32 VSUBS 0.030109f
C919 VP.n33 VSUBS 0.030109f
C920 VP.n34 VSUBS 0.030109f
C921 VP.n35 VSUBS 0.024328f
C922 VP.n36 VSUBS 0.059671f
C923 VP.n37 VSUBS 0.055283f
C924 VP.n38 VSUBS 0.048588f
C925 VP.n39 VSUBS 0.054062f
.ends

