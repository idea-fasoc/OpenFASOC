* NGSPICE file created from diff_pair_sample_0972.ext - technology: sky130A

.subckt diff_pair_sample_0972 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VN.t0 VDD2.t0 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=1.22265 ps=7.74 w=7.41 l=0.17
X1 VTAIL.t11 VN.t1 VDD2.t4 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X2 VTAIL.t2 VP.t0 VDD1.t7 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=1.22265 ps=7.74 w=7.41 l=0.17
X3 B.t11 B.t9 B.t10 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=0 ps=0 w=7.41 l=0.17
X4 VDD1.t6 VP.t1 VTAIL.t4 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=2.8899 ps=15.6 w=7.41 l=0.17
X5 VDD2.t1 VN.t2 VTAIL.t10 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=2.8899 ps=15.6 w=7.41 l=0.17
X6 VTAIL.t1 VP.t2 VDD1.t5 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=1.22265 ps=7.74 w=7.41 l=0.17
X7 VDD1.t4 VP.t3 VTAIL.t13 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X8 VTAIL.t9 VN.t3 VDD2.t6 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=1.22265 ps=7.74 w=7.41 l=0.17
X9 B.t8 B.t6 B.t7 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=0 ps=0 w=7.41 l=0.17
X10 B.t5 B.t3 B.t4 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=0 ps=0 w=7.41 l=0.17
X11 VTAIL.t14 VP.t4 VDD1.t3 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X12 VTAIL.t15 VP.t5 VDD1.t2 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X13 VDD1.t1 VP.t6 VTAIL.t0 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=2.8899 ps=15.6 w=7.41 l=0.17
X14 B.t2 B.t0 B.t1 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=2.8899 pd=15.6 as=0 ps=0 w=7.41 l=0.17
X15 VDD2.t5 VN.t4 VTAIL.t8 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=2.8899 ps=15.6 w=7.41 l=0.17
X16 VDD2.t7 VN.t5 VTAIL.t7 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X17 VTAIL.t6 VN.t6 VDD2.t2 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X18 VDD2.t3 VN.t7 VTAIL.t5 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
X19 VDD1.t0 VP.t7 VTAIL.t3 w_n1470_n2450# sky130_fd_pr__pfet_01v8 ad=1.22265 pd=7.74 as=1.22265 ps=7.74 w=7.41 l=0.17
R0 VN.n5 VN.t4 1272.7
R1 VN.n1 VN.t0 1272.7
R2 VN.n12 VN.t3 1272.7
R3 VN.n8 VN.t2 1272.7
R4 VN.n4 VN.t6 1236.19
R5 VN.n2 VN.t7 1236.19
R6 VN.n11 VN.t5 1236.19
R7 VN.n9 VN.t1 1236.19
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN.n2 VN.n1 36.5157
R15 VN.n3 VN.n2 36.5157
R16 VN.n4 VN.n3 36.5157
R17 VN.n5 VN.n4 36.5157
R18 VN.n12 VN.n11 36.5157
R19 VN.n11 VN.n10 36.5157
R20 VN.n10 VN.n9 36.5157
R21 VN.n9 VN.n8 36.5157
R22 VN VN.n13 36.4418
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VDD2.n2 VDD2.n1 84.8807
R27 VDD2.n2 VDD2.n0 84.8807
R28 VDD2 VDD2.n5 84.8779
R29 VDD2.n4 VDD2.n3 84.7207
R30 VDD2.n4 VDD2.n2 32.0429
R31 VDD2.n5 VDD2.t4 4.38714
R32 VDD2.n5 VDD2.t1 4.38714
R33 VDD2.n3 VDD2.t6 4.38714
R34 VDD2.n3 VDD2.t7 4.38714
R35 VDD2.n1 VDD2.t2 4.38714
R36 VDD2.n1 VDD2.t5 4.38714
R37 VDD2.n0 VDD2.t0 4.38714
R38 VDD2.n0 VDD2.t3 4.38714
R39 VDD2 VDD2.n4 0.274207
R40 VTAIL.n322 VTAIL.n288 756.745
R41 VTAIL.n36 VTAIL.n2 756.745
R42 VTAIL.n76 VTAIL.n42 756.745
R43 VTAIL.n118 VTAIL.n84 756.745
R44 VTAIL.n282 VTAIL.n248 756.745
R45 VTAIL.n240 VTAIL.n206 756.745
R46 VTAIL.n200 VTAIL.n166 756.745
R47 VTAIL.n158 VTAIL.n124 756.745
R48 VTAIL.n300 VTAIL.n299 585
R49 VTAIL.n305 VTAIL.n304 585
R50 VTAIL.n307 VTAIL.n306 585
R51 VTAIL.n296 VTAIL.n295 585
R52 VTAIL.n313 VTAIL.n312 585
R53 VTAIL.n315 VTAIL.n314 585
R54 VTAIL.n292 VTAIL.n291 585
R55 VTAIL.n321 VTAIL.n320 585
R56 VTAIL.n323 VTAIL.n322 585
R57 VTAIL.n14 VTAIL.n13 585
R58 VTAIL.n19 VTAIL.n18 585
R59 VTAIL.n21 VTAIL.n20 585
R60 VTAIL.n10 VTAIL.n9 585
R61 VTAIL.n27 VTAIL.n26 585
R62 VTAIL.n29 VTAIL.n28 585
R63 VTAIL.n6 VTAIL.n5 585
R64 VTAIL.n35 VTAIL.n34 585
R65 VTAIL.n37 VTAIL.n36 585
R66 VTAIL.n54 VTAIL.n53 585
R67 VTAIL.n59 VTAIL.n58 585
R68 VTAIL.n61 VTAIL.n60 585
R69 VTAIL.n50 VTAIL.n49 585
R70 VTAIL.n67 VTAIL.n66 585
R71 VTAIL.n69 VTAIL.n68 585
R72 VTAIL.n46 VTAIL.n45 585
R73 VTAIL.n75 VTAIL.n74 585
R74 VTAIL.n77 VTAIL.n76 585
R75 VTAIL.n96 VTAIL.n95 585
R76 VTAIL.n101 VTAIL.n100 585
R77 VTAIL.n103 VTAIL.n102 585
R78 VTAIL.n92 VTAIL.n91 585
R79 VTAIL.n109 VTAIL.n108 585
R80 VTAIL.n111 VTAIL.n110 585
R81 VTAIL.n88 VTAIL.n87 585
R82 VTAIL.n117 VTAIL.n116 585
R83 VTAIL.n119 VTAIL.n118 585
R84 VTAIL.n283 VTAIL.n282 585
R85 VTAIL.n281 VTAIL.n280 585
R86 VTAIL.n252 VTAIL.n251 585
R87 VTAIL.n275 VTAIL.n274 585
R88 VTAIL.n273 VTAIL.n272 585
R89 VTAIL.n256 VTAIL.n255 585
R90 VTAIL.n267 VTAIL.n266 585
R91 VTAIL.n265 VTAIL.n264 585
R92 VTAIL.n260 VTAIL.n259 585
R93 VTAIL.n241 VTAIL.n240 585
R94 VTAIL.n239 VTAIL.n238 585
R95 VTAIL.n210 VTAIL.n209 585
R96 VTAIL.n233 VTAIL.n232 585
R97 VTAIL.n231 VTAIL.n230 585
R98 VTAIL.n214 VTAIL.n213 585
R99 VTAIL.n225 VTAIL.n224 585
R100 VTAIL.n223 VTAIL.n222 585
R101 VTAIL.n218 VTAIL.n217 585
R102 VTAIL.n201 VTAIL.n200 585
R103 VTAIL.n199 VTAIL.n198 585
R104 VTAIL.n170 VTAIL.n169 585
R105 VTAIL.n193 VTAIL.n192 585
R106 VTAIL.n191 VTAIL.n190 585
R107 VTAIL.n174 VTAIL.n173 585
R108 VTAIL.n185 VTAIL.n184 585
R109 VTAIL.n183 VTAIL.n182 585
R110 VTAIL.n178 VTAIL.n177 585
R111 VTAIL.n159 VTAIL.n158 585
R112 VTAIL.n157 VTAIL.n156 585
R113 VTAIL.n128 VTAIL.n127 585
R114 VTAIL.n151 VTAIL.n150 585
R115 VTAIL.n149 VTAIL.n148 585
R116 VTAIL.n132 VTAIL.n131 585
R117 VTAIL.n143 VTAIL.n142 585
R118 VTAIL.n141 VTAIL.n140 585
R119 VTAIL.n136 VTAIL.n135 585
R120 VTAIL.n301 VTAIL.t8 327.483
R121 VTAIL.n15 VTAIL.t12 327.483
R122 VTAIL.n55 VTAIL.t0 327.483
R123 VTAIL.n97 VTAIL.t1 327.483
R124 VTAIL.n261 VTAIL.t4 327.483
R125 VTAIL.n219 VTAIL.t2 327.483
R126 VTAIL.n179 VTAIL.t10 327.483
R127 VTAIL.n137 VTAIL.t9 327.483
R128 VTAIL.n305 VTAIL.n299 171.744
R129 VTAIL.n306 VTAIL.n305 171.744
R130 VTAIL.n306 VTAIL.n295 171.744
R131 VTAIL.n313 VTAIL.n295 171.744
R132 VTAIL.n314 VTAIL.n313 171.744
R133 VTAIL.n314 VTAIL.n291 171.744
R134 VTAIL.n321 VTAIL.n291 171.744
R135 VTAIL.n322 VTAIL.n321 171.744
R136 VTAIL.n19 VTAIL.n13 171.744
R137 VTAIL.n20 VTAIL.n19 171.744
R138 VTAIL.n20 VTAIL.n9 171.744
R139 VTAIL.n27 VTAIL.n9 171.744
R140 VTAIL.n28 VTAIL.n27 171.744
R141 VTAIL.n28 VTAIL.n5 171.744
R142 VTAIL.n35 VTAIL.n5 171.744
R143 VTAIL.n36 VTAIL.n35 171.744
R144 VTAIL.n59 VTAIL.n53 171.744
R145 VTAIL.n60 VTAIL.n59 171.744
R146 VTAIL.n60 VTAIL.n49 171.744
R147 VTAIL.n67 VTAIL.n49 171.744
R148 VTAIL.n68 VTAIL.n67 171.744
R149 VTAIL.n68 VTAIL.n45 171.744
R150 VTAIL.n75 VTAIL.n45 171.744
R151 VTAIL.n76 VTAIL.n75 171.744
R152 VTAIL.n101 VTAIL.n95 171.744
R153 VTAIL.n102 VTAIL.n101 171.744
R154 VTAIL.n102 VTAIL.n91 171.744
R155 VTAIL.n109 VTAIL.n91 171.744
R156 VTAIL.n110 VTAIL.n109 171.744
R157 VTAIL.n110 VTAIL.n87 171.744
R158 VTAIL.n117 VTAIL.n87 171.744
R159 VTAIL.n118 VTAIL.n117 171.744
R160 VTAIL.n282 VTAIL.n281 171.744
R161 VTAIL.n281 VTAIL.n251 171.744
R162 VTAIL.n274 VTAIL.n251 171.744
R163 VTAIL.n274 VTAIL.n273 171.744
R164 VTAIL.n273 VTAIL.n255 171.744
R165 VTAIL.n266 VTAIL.n255 171.744
R166 VTAIL.n266 VTAIL.n265 171.744
R167 VTAIL.n265 VTAIL.n259 171.744
R168 VTAIL.n240 VTAIL.n239 171.744
R169 VTAIL.n239 VTAIL.n209 171.744
R170 VTAIL.n232 VTAIL.n209 171.744
R171 VTAIL.n232 VTAIL.n231 171.744
R172 VTAIL.n231 VTAIL.n213 171.744
R173 VTAIL.n224 VTAIL.n213 171.744
R174 VTAIL.n224 VTAIL.n223 171.744
R175 VTAIL.n223 VTAIL.n217 171.744
R176 VTAIL.n200 VTAIL.n199 171.744
R177 VTAIL.n199 VTAIL.n169 171.744
R178 VTAIL.n192 VTAIL.n169 171.744
R179 VTAIL.n192 VTAIL.n191 171.744
R180 VTAIL.n191 VTAIL.n173 171.744
R181 VTAIL.n184 VTAIL.n173 171.744
R182 VTAIL.n184 VTAIL.n183 171.744
R183 VTAIL.n183 VTAIL.n177 171.744
R184 VTAIL.n158 VTAIL.n157 171.744
R185 VTAIL.n157 VTAIL.n127 171.744
R186 VTAIL.n150 VTAIL.n127 171.744
R187 VTAIL.n150 VTAIL.n149 171.744
R188 VTAIL.n149 VTAIL.n131 171.744
R189 VTAIL.n142 VTAIL.n131 171.744
R190 VTAIL.n142 VTAIL.n141 171.744
R191 VTAIL.n141 VTAIL.n135 171.744
R192 VTAIL.t8 VTAIL.n299 85.8723
R193 VTAIL.t12 VTAIL.n13 85.8723
R194 VTAIL.t0 VTAIL.n53 85.8723
R195 VTAIL.t1 VTAIL.n95 85.8723
R196 VTAIL.t4 VTAIL.n259 85.8723
R197 VTAIL.t2 VTAIL.n217 85.8723
R198 VTAIL.t10 VTAIL.n177 85.8723
R199 VTAIL.t9 VTAIL.n135 85.8723
R200 VTAIL.n247 VTAIL.n246 68.0419
R201 VTAIL.n165 VTAIL.n164 68.0419
R202 VTAIL.n1 VTAIL.n0 68.0418
R203 VTAIL.n83 VTAIL.n82 68.0418
R204 VTAIL.n327 VTAIL.n326 31.6035
R205 VTAIL.n41 VTAIL.n40 31.6035
R206 VTAIL.n81 VTAIL.n80 31.6035
R207 VTAIL.n123 VTAIL.n122 31.6035
R208 VTAIL.n287 VTAIL.n286 31.6035
R209 VTAIL.n245 VTAIL.n244 31.6035
R210 VTAIL.n205 VTAIL.n204 31.6035
R211 VTAIL.n163 VTAIL.n162 31.6035
R212 VTAIL.n327 VTAIL.n287 19.1858
R213 VTAIL.n163 VTAIL.n123 19.1858
R214 VTAIL.n301 VTAIL.n300 16.3891
R215 VTAIL.n15 VTAIL.n14 16.3891
R216 VTAIL.n55 VTAIL.n54 16.3891
R217 VTAIL.n97 VTAIL.n96 16.3891
R218 VTAIL.n261 VTAIL.n260 16.3891
R219 VTAIL.n219 VTAIL.n218 16.3891
R220 VTAIL.n179 VTAIL.n178 16.3891
R221 VTAIL.n137 VTAIL.n136 16.3891
R222 VTAIL.n304 VTAIL.n303 12.8005
R223 VTAIL.n18 VTAIL.n17 12.8005
R224 VTAIL.n58 VTAIL.n57 12.8005
R225 VTAIL.n100 VTAIL.n99 12.8005
R226 VTAIL.n264 VTAIL.n263 12.8005
R227 VTAIL.n222 VTAIL.n221 12.8005
R228 VTAIL.n182 VTAIL.n181 12.8005
R229 VTAIL.n140 VTAIL.n139 12.8005
R230 VTAIL.n307 VTAIL.n298 12.0247
R231 VTAIL.n21 VTAIL.n12 12.0247
R232 VTAIL.n61 VTAIL.n52 12.0247
R233 VTAIL.n103 VTAIL.n94 12.0247
R234 VTAIL.n267 VTAIL.n258 12.0247
R235 VTAIL.n225 VTAIL.n216 12.0247
R236 VTAIL.n185 VTAIL.n176 12.0247
R237 VTAIL.n143 VTAIL.n134 12.0247
R238 VTAIL.n308 VTAIL.n296 11.249
R239 VTAIL.n22 VTAIL.n10 11.249
R240 VTAIL.n62 VTAIL.n50 11.249
R241 VTAIL.n104 VTAIL.n92 11.249
R242 VTAIL.n268 VTAIL.n256 11.249
R243 VTAIL.n226 VTAIL.n214 11.249
R244 VTAIL.n186 VTAIL.n174 11.249
R245 VTAIL.n144 VTAIL.n132 11.249
R246 VTAIL.n312 VTAIL.n311 10.4732
R247 VTAIL.n26 VTAIL.n25 10.4732
R248 VTAIL.n66 VTAIL.n65 10.4732
R249 VTAIL.n108 VTAIL.n107 10.4732
R250 VTAIL.n272 VTAIL.n271 10.4732
R251 VTAIL.n230 VTAIL.n229 10.4732
R252 VTAIL.n190 VTAIL.n189 10.4732
R253 VTAIL.n148 VTAIL.n147 10.4732
R254 VTAIL.n315 VTAIL.n294 9.69747
R255 VTAIL.n29 VTAIL.n8 9.69747
R256 VTAIL.n69 VTAIL.n48 9.69747
R257 VTAIL.n111 VTAIL.n90 9.69747
R258 VTAIL.n275 VTAIL.n254 9.69747
R259 VTAIL.n233 VTAIL.n212 9.69747
R260 VTAIL.n193 VTAIL.n172 9.69747
R261 VTAIL.n151 VTAIL.n130 9.69747
R262 VTAIL.n326 VTAIL.n325 9.45567
R263 VTAIL.n40 VTAIL.n39 9.45567
R264 VTAIL.n80 VTAIL.n79 9.45567
R265 VTAIL.n122 VTAIL.n121 9.45567
R266 VTAIL.n286 VTAIL.n285 9.45567
R267 VTAIL.n244 VTAIL.n243 9.45567
R268 VTAIL.n204 VTAIL.n203 9.45567
R269 VTAIL.n162 VTAIL.n161 9.45567
R270 VTAIL.n325 VTAIL.n324 9.3005
R271 VTAIL.n319 VTAIL.n318 9.3005
R272 VTAIL.n317 VTAIL.n316 9.3005
R273 VTAIL.n294 VTAIL.n293 9.3005
R274 VTAIL.n311 VTAIL.n310 9.3005
R275 VTAIL.n309 VTAIL.n308 9.3005
R276 VTAIL.n298 VTAIL.n297 9.3005
R277 VTAIL.n303 VTAIL.n302 9.3005
R278 VTAIL.n290 VTAIL.n289 9.3005
R279 VTAIL.n39 VTAIL.n38 9.3005
R280 VTAIL.n33 VTAIL.n32 9.3005
R281 VTAIL.n31 VTAIL.n30 9.3005
R282 VTAIL.n8 VTAIL.n7 9.3005
R283 VTAIL.n25 VTAIL.n24 9.3005
R284 VTAIL.n23 VTAIL.n22 9.3005
R285 VTAIL.n12 VTAIL.n11 9.3005
R286 VTAIL.n17 VTAIL.n16 9.3005
R287 VTAIL.n4 VTAIL.n3 9.3005
R288 VTAIL.n79 VTAIL.n78 9.3005
R289 VTAIL.n73 VTAIL.n72 9.3005
R290 VTAIL.n71 VTAIL.n70 9.3005
R291 VTAIL.n48 VTAIL.n47 9.3005
R292 VTAIL.n65 VTAIL.n64 9.3005
R293 VTAIL.n63 VTAIL.n62 9.3005
R294 VTAIL.n52 VTAIL.n51 9.3005
R295 VTAIL.n57 VTAIL.n56 9.3005
R296 VTAIL.n44 VTAIL.n43 9.3005
R297 VTAIL.n121 VTAIL.n120 9.3005
R298 VTAIL.n115 VTAIL.n114 9.3005
R299 VTAIL.n113 VTAIL.n112 9.3005
R300 VTAIL.n90 VTAIL.n89 9.3005
R301 VTAIL.n107 VTAIL.n106 9.3005
R302 VTAIL.n105 VTAIL.n104 9.3005
R303 VTAIL.n94 VTAIL.n93 9.3005
R304 VTAIL.n99 VTAIL.n98 9.3005
R305 VTAIL.n86 VTAIL.n85 9.3005
R306 VTAIL.n285 VTAIL.n284 9.3005
R307 VTAIL.n250 VTAIL.n249 9.3005
R308 VTAIL.n279 VTAIL.n278 9.3005
R309 VTAIL.n277 VTAIL.n276 9.3005
R310 VTAIL.n254 VTAIL.n253 9.3005
R311 VTAIL.n271 VTAIL.n270 9.3005
R312 VTAIL.n269 VTAIL.n268 9.3005
R313 VTAIL.n258 VTAIL.n257 9.3005
R314 VTAIL.n263 VTAIL.n262 9.3005
R315 VTAIL.n243 VTAIL.n242 9.3005
R316 VTAIL.n208 VTAIL.n207 9.3005
R317 VTAIL.n237 VTAIL.n236 9.3005
R318 VTAIL.n235 VTAIL.n234 9.3005
R319 VTAIL.n212 VTAIL.n211 9.3005
R320 VTAIL.n229 VTAIL.n228 9.3005
R321 VTAIL.n227 VTAIL.n226 9.3005
R322 VTAIL.n216 VTAIL.n215 9.3005
R323 VTAIL.n221 VTAIL.n220 9.3005
R324 VTAIL.n203 VTAIL.n202 9.3005
R325 VTAIL.n168 VTAIL.n167 9.3005
R326 VTAIL.n197 VTAIL.n196 9.3005
R327 VTAIL.n195 VTAIL.n194 9.3005
R328 VTAIL.n172 VTAIL.n171 9.3005
R329 VTAIL.n189 VTAIL.n188 9.3005
R330 VTAIL.n187 VTAIL.n186 9.3005
R331 VTAIL.n176 VTAIL.n175 9.3005
R332 VTAIL.n181 VTAIL.n180 9.3005
R333 VTAIL.n161 VTAIL.n160 9.3005
R334 VTAIL.n126 VTAIL.n125 9.3005
R335 VTAIL.n155 VTAIL.n154 9.3005
R336 VTAIL.n153 VTAIL.n152 9.3005
R337 VTAIL.n130 VTAIL.n129 9.3005
R338 VTAIL.n147 VTAIL.n146 9.3005
R339 VTAIL.n145 VTAIL.n144 9.3005
R340 VTAIL.n134 VTAIL.n133 9.3005
R341 VTAIL.n139 VTAIL.n138 9.3005
R342 VTAIL.n316 VTAIL.n292 8.92171
R343 VTAIL.n30 VTAIL.n6 8.92171
R344 VTAIL.n70 VTAIL.n46 8.92171
R345 VTAIL.n112 VTAIL.n88 8.92171
R346 VTAIL.n276 VTAIL.n252 8.92171
R347 VTAIL.n234 VTAIL.n210 8.92171
R348 VTAIL.n194 VTAIL.n170 8.92171
R349 VTAIL.n152 VTAIL.n128 8.92171
R350 VTAIL.n320 VTAIL.n319 8.14595
R351 VTAIL.n34 VTAIL.n33 8.14595
R352 VTAIL.n74 VTAIL.n73 8.14595
R353 VTAIL.n116 VTAIL.n115 8.14595
R354 VTAIL.n280 VTAIL.n279 8.14595
R355 VTAIL.n238 VTAIL.n237 8.14595
R356 VTAIL.n198 VTAIL.n197 8.14595
R357 VTAIL.n156 VTAIL.n155 8.14595
R358 VTAIL.n323 VTAIL.n290 7.3702
R359 VTAIL.n326 VTAIL.n288 7.3702
R360 VTAIL.n37 VTAIL.n4 7.3702
R361 VTAIL.n40 VTAIL.n2 7.3702
R362 VTAIL.n77 VTAIL.n44 7.3702
R363 VTAIL.n80 VTAIL.n42 7.3702
R364 VTAIL.n119 VTAIL.n86 7.3702
R365 VTAIL.n122 VTAIL.n84 7.3702
R366 VTAIL.n286 VTAIL.n248 7.3702
R367 VTAIL.n283 VTAIL.n250 7.3702
R368 VTAIL.n244 VTAIL.n206 7.3702
R369 VTAIL.n241 VTAIL.n208 7.3702
R370 VTAIL.n204 VTAIL.n166 7.3702
R371 VTAIL.n201 VTAIL.n168 7.3702
R372 VTAIL.n162 VTAIL.n124 7.3702
R373 VTAIL.n159 VTAIL.n126 7.3702
R374 VTAIL.n324 VTAIL.n323 6.59444
R375 VTAIL.n324 VTAIL.n288 6.59444
R376 VTAIL.n38 VTAIL.n37 6.59444
R377 VTAIL.n38 VTAIL.n2 6.59444
R378 VTAIL.n78 VTAIL.n77 6.59444
R379 VTAIL.n78 VTAIL.n42 6.59444
R380 VTAIL.n120 VTAIL.n119 6.59444
R381 VTAIL.n120 VTAIL.n84 6.59444
R382 VTAIL.n284 VTAIL.n248 6.59444
R383 VTAIL.n284 VTAIL.n283 6.59444
R384 VTAIL.n242 VTAIL.n206 6.59444
R385 VTAIL.n242 VTAIL.n241 6.59444
R386 VTAIL.n202 VTAIL.n166 6.59444
R387 VTAIL.n202 VTAIL.n201 6.59444
R388 VTAIL.n160 VTAIL.n124 6.59444
R389 VTAIL.n160 VTAIL.n159 6.59444
R390 VTAIL.n320 VTAIL.n290 5.81868
R391 VTAIL.n34 VTAIL.n4 5.81868
R392 VTAIL.n74 VTAIL.n44 5.81868
R393 VTAIL.n116 VTAIL.n86 5.81868
R394 VTAIL.n280 VTAIL.n250 5.81868
R395 VTAIL.n238 VTAIL.n208 5.81868
R396 VTAIL.n198 VTAIL.n168 5.81868
R397 VTAIL.n156 VTAIL.n126 5.81868
R398 VTAIL.n319 VTAIL.n292 5.04292
R399 VTAIL.n33 VTAIL.n6 5.04292
R400 VTAIL.n73 VTAIL.n46 5.04292
R401 VTAIL.n115 VTAIL.n88 5.04292
R402 VTAIL.n279 VTAIL.n252 5.04292
R403 VTAIL.n237 VTAIL.n210 5.04292
R404 VTAIL.n197 VTAIL.n170 5.04292
R405 VTAIL.n155 VTAIL.n128 5.04292
R406 VTAIL.n0 VTAIL.t5 4.38714
R407 VTAIL.n0 VTAIL.t6 4.38714
R408 VTAIL.n82 VTAIL.t13 4.38714
R409 VTAIL.n82 VTAIL.t14 4.38714
R410 VTAIL.n246 VTAIL.t3 4.38714
R411 VTAIL.n246 VTAIL.t15 4.38714
R412 VTAIL.n164 VTAIL.t7 4.38714
R413 VTAIL.n164 VTAIL.t11 4.38714
R414 VTAIL.n316 VTAIL.n315 4.26717
R415 VTAIL.n30 VTAIL.n29 4.26717
R416 VTAIL.n70 VTAIL.n69 4.26717
R417 VTAIL.n112 VTAIL.n111 4.26717
R418 VTAIL.n276 VTAIL.n275 4.26717
R419 VTAIL.n234 VTAIL.n233 4.26717
R420 VTAIL.n194 VTAIL.n193 4.26717
R421 VTAIL.n152 VTAIL.n151 4.26717
R422 VTAIL.n302 VTAIL.n301 3.71019
R423 VTAIL.n16 VTAIL.n15 3.71019
R424 VTAIL.n56 VTAIL.n55 3.71019
R425 VTAIL.n98 VTAIL.n97 3.71019
R426 VTAIL.n262 VTAIL.n261 3.71019
R427 VTAIL.n220 VTAIL.n219 3.71019
R428 VTAIL.n180 VTAIL.n179 3.71019
R429 VTAIL.n138 VTAIL.n137 3.71019
R430 VTAIL.n312 VTAIL.n294 3.49141
R431 VTAIL.n26 VTAIL.n8 3.49141
R432 VTAIL.n66 VTAIL.n48 3.49141
R433 VTAIL.n108 VTAIL.n90 3.49141
R434 VTAIL.n272 VTAIL.n254 3.49141
R435 VTAIL.n230 VTAIL.n212 3.49141
R436 VTAIL.n190 VTAIL.n172 3.49141
R437 VTAIL.n148 VTAIL.n130 3.49141
R438 VTAIL.n311 VTAIL.n296 2.71565
R439 VTAIL.n25 VTAIL.n10 2.71565
R440 VTAIL.n65 VTAIL.n50 2.71565
R441 VTAIL.n107 VTAIL.n92 2.71565
R442 VTAIL.n271 VTAIL.n256 2.71565
R443 VTAIL.n229 VTAIL.n214 2.71565
R444 VTAIL.n189 VTAIL.n174 2.71565
R445 VTAIL.n147 VTAIL.n132 2.71565
R446 VTAIL.n308 VTAIL.n307 1.93989
R447 VTAIL.n22 VTAIL.n21 1.93989
R448 VTAIL.n62 VTAIL.n61 1.93989
R449 VTAIL.n104 VTAIL.n103 1.93989
R450 VTAIL.n268 VTAIL.n267 1.93989
R451 VTAIL.n226 VTAIL.n225 1.93989
R452 VTAIL.n186 VTAIL.n185 1.93989
R453 VTAIL.n144 VTAIL.n143 1.93989
R454 VTAIL.n304 VTAIL.n298 1.16414
R455 VTAIL.n18 VTAIL.n12 1.16414
R456 VTAIL.n58 VTAIL.n52 1.16414
R457 VTAIL.n100 VTAIL.n94 1.16414
R458 VTAIL.n264 VTAIL.n258 1.16414
R459 VTAIL.n222 VTAIL.n216 1.16414
R460 VTAIL.n182 VTAIL.n176 1.16414
R461 VTAIL.n140 VTAIL.n134 1.16414
R462 VTAIL.n245 VTAIL.n205 0.470328
R463 VTAIL.n81 VTAIL.n41 0.470328
R464 VTAIL.n165 VTAIL.n163 0.431534
R465 VTAIL.n205 VTAIL.n165 0.431534
R466 VTAIL.n247 VTAIL.n245 0.431534
R467 VTAIL.n287 VTAIL.n247 0.431534
R468 VTAIL.n123 VTAIL.n83 0.431534
R469 VTAIL.n83 VTAIL.n81 0.431534
R470 VTAIL.n41 VTAIL.n1 0.431534
R471 VTAIL.n303 VTAIL.n300 0.388379
R472 VTAIL.n17 VTAIL.n14 0.388379
R473 VTAIL.n57 VTAIL.n54 0.388379
R474 VTAIL.n99 VTAIL.n96 0.388379
R475 VTAIL.n263 VTAIL.n260 0.388379
R476 VTAIL.n221 VTAIL.n218 0.388379
R477 VTAIL.n181 VTAIL.n178 0.388379
R478 VTAIL.n139 VTAIL.n136 0.388379
R479 VTAIL VTAIL.n327 0.373345
R480 VTAIL.n302 VTAIL.n297 0.155672
R481 VTAIL.n309 VTAIL.n297 0.155672
R482 VTAIL.n310 VTAIL.n309 0.155672
R483 VTAIL.n310 VTAIL.n293 0.155672
R484 VTAIL.n317 VTAIL.n293 0.155672
R485 VTAIL.n318 VTAIL.n317 0.155672
R486 VTAIL.n318 VTAIL.n289 0.155672
R487 VTAIL.n325 VTAIL.n289 0.155672
R488 VTAIL.n16 VTAIL.n11 0.155672
R489 VTAIL.n23 VTAIL.n11 0.155672
R490 VTAIL.n24 VTAIL.n23 0.155672
R491 VTAIL.n24 VTAIL.n7 0.155672
R492 VTAIL.n31 VTAIL.n7 0.155672
R493 VTAIL.n32 VTAIL.n31 0.155672
R494 VTAIL.n32 VTAIL.n3 0.155672
R495 VTAIL.n39 VTAIL.n3 0.155672
R496 VTAIL.n56 VTAIL.n51 0.155672
R497 VTAIL.n63 VTAIL.n51 0.155672
R498 VTAIL.n64 VTAIL.n63 0.155672
R499 VTAIL.n64 VTAIL.n47 0.155672
R500 VTAIL.n71 VTAIL.n47 0.155672
R501 VTAIL.n72 VTAIL.n71 0.155672
R502 VTAIL.n72 VTAIL.n43 0.155672
R503 VTAIL.n79 VTAIL.n43 0.155672
R504 VTAIL.n98 VTAIL.n93 0.155672
R505 VTAIL.n105 VTAIL.n93 0.155672
R506 VTAIL.n106 VTAIL.n105 0.155672
R507 VTAIL.n106 VTAIL.n89 0.155672
R508 VTAIL.n113 VTAIL.n89 0.155672
R509 VTAIL.n114 VTAIL.n113 0.155672
R510 VTAIL.n114 VTAIL.n85 0.155672
R511 VTAIL.n121 VTAIL.n85 0.155672
R512 VTAIL.n285 VTAIL.n249 0.155672
R513 VTAIL.n278 VTAIL.n249 0.155672
R514 VTAIL.n278 VTAIL.n277 0.155672
R515 VTAIL.n277 VTAIL.n253 0.155672
R516 VTAIL.n270 VTAIL.n253 0.155672
R517 VTAIL.n270 VTAIL.n269 0.155672
R518 VTAIL.n269 VTAIL.n257 0.155672
R519 VTAIL.n262 VTAIL.n257 0.155672
R520 VTAIL.n243 VTAIL.n207 0.155672
R521 VTAIL.n236 VTAIL.n207 0.155672
R522 VTAIL.n236 VTAIL.n235 0.155672
R523 VTAIL.n235 VTAIL.n211 0.155672
R524 VTAIL.n228 VTAIL.n211 0.155672
R525 VTAIL.n228 VTAIL.n227 0.155672
R526 VTAIL.n227 VTAIL.n215 0.155672
R527 VTAIL.n220 VTAIL.n215 0.155672
R528 VTAIL.n203 VTAIL.n167 0.155672
R529 VTAIL.n196 VTAIL.n167 0.155672
R530 VTAIL.n196 VTAIL.n195 0.155672
R531 VTAIL.n195 VTAIL.n171 0.155672
R532 VTAIL.n188 VTAIL.n171 0.155672
R533 VTAIL.n188 VTAIL.n187 0.155672
R534 VTAIL.n187 VTAIL.n175 0.155672
R535 VTAIL.n180 VTAIL.n175 0.155672
R536 VTAIL.n161 VTAIL.n125 0.155672
R537 VTAIL.n154 VTAIL.n125 0.155672
R538 VTAIL.n154 VTAIL.n153 0.155672
R539 VTAIL.n153 VTAIL.n129 0.155672
R540 VTAIL.n146 VTAIL.n129 0.155672
R541 VTAIL.n146 VTAIL.n145 0.155672
R542 VTAIL.n145 VTAIL.n133 0.155672
R543 VTAIL.n138 VTAIL.n133 0.155672
R544 VTAIL VTAIL.n1 0.0586897
R545 VP.n13 VP.t6 1272.7
R546 VP.n9 VP.t2 1272.7
R547 VP.n2 VP.t0 1272.7
R548 VP.n6 VP.t1 1272.7
R549 VP.n12 VP.t4 1236.19
R550 VP.n10 VP.t3 1236.19
R551 VP.n3 VP.t7 1236.19
R552 VP.n5 VP.t5 1236.19
R553 VP.n2 VP.n1 161.489
R554 VP.n14 VP.n13 161.3
R555 VP.n4 VP.n1 161.3
R556 VP.n7 VP.n6 161.3
R557 VP.n11 VP.n0 161.3
R558 VP.n9 VP.n8 161.3
R559 VP.n10 VP.n9 36.5157
R560 VP.n11 VP.n10 36.5157
R561 VP.n12 VP.n11 36.5157
R562 VP.n13 VP.n12 36.5157
R563 VP.n3 VP.n2 36.5157
R564 VP.n4 VP.n3 36.5157
R565 VP.n5 VP.n4 36.5157
R566 VP.n6 VP.n5 36.5157
R567 VP.n8 VP.n7 36.0611
R568 VP.n7 VP.n1 0.189894
R569 VP.n8 VP.n0 0.189894
R570 VP.n14 VP.n0 0.189894
R571 VP VP.n14 0.0516364
R572 VDD1 VDD1.n0 84.9944
R573 VDD1.n3 VDD1.n2 84.8807
R574 VDD1.n3 VDD1.n1 84.8807
R575 VDD1.n5 VDD1.n4 84.7205
R576 VDD1.n5 VDD1.n3 32.6259
R577 VDD1.n4 VDD1.t2 4.38714
R578 VDD1.n4 VDD1.t6 4.38714
R579 VDD1.n0 VDD1.t7 4.38714
R580 VDD1.n0 VDD1.t0 4.38714
R581 VDD1.n2 VDD1.t3 4.38714
R582 VDD1.n2 VDD1.t1 4.38714
R583 VDD1.n1 VDD1.t5 4.38714
R584 VDD1.n1 VDD1.t4 4.38714
R585 VDD1 VDD1.n5 0.157828
R586 B.n83 B.t6 1297.46
R587 B.n183 B.t3 1297.46
R588 B.n32 B.t9 1297.46
R589 B.n24 B.t0 1297.46
R590 B.n229 B.n228 585
R591 B.n227 B.n64 585
R592 B.n226 B.n225 585
R593 B.n224 B.n65 585
R594 B.n223 B.n222 585
R595 B.n221 B.n66 585
R596 B.n220 B.n219 585
R597 B.n218 B.n67 585
R598 B.n217 B.n216 585
R599 B.n215 B.n68 585
R600 B.n214 B.n213 585
R601 B.n212 B.n69 585
R602 B.n211 B.n210 585
R603 B.n209 B.n70 585
R604 B.n208 B.n207 585
R605 B.n206 B.n71 585
R606 B.n205 B.n204 585
R607 B.n203 B.n72 585
R608 B.n202 B.n201 585
R609 B.n200 B.n73 585
R610 B.n199 B.n198 585
R611 B.n197 B.n74 585
R612 B.n196 B.n195 585
R613 B.n194 B.n75 585
R614 B.n193 B.n192 585
R615 B.n191 B.n76 585
R616 B.n190 B.n189 585
R617 B.n188 B.n77 585
R618 B.n187 B.n186 585
R619 B.n182 B.n78 585
R620 B.n181 B.n180 585
R621 B.n179 B.n79 585
R622 B.n178 B.n177 585
R623 B.n176 B.n80 585
R624 B.n175 B.n174 585
R625 B.n173 B.n81 585
R626 B.n172 B.n171 585
R627 B.n170 B.n82 585
R628 B.n168 B.n167 585
R629 B.n166 B.n85 585
R630 B.n165 B.n164 585
R631 B.n163 B.n86 585
R632 B.n162 B.n161 585
R633 B.n160 B.n87 585
R634 B.n159 B.n158 585
R635 B.n157 B.n88 585
R636 B.n156 B.n155 585
R637 B.n154 B.n89 585
R638 B.n153 B.n152 585
R639 B.n151 B.n90 585
R640 B.n150 B.n149 585
R641 B.n148 B.n91 585
R642 B.n147 B.n146 585
R643 B.n145 B.n92 585
R644 B.n144 B.n143 585
R645 B.n142 B.n93 585
R646 B.n141 B.n140 585
R647 B.n139 B.n94 585
R648 B.n138 B.n137 585
R649 B.n136 B.n95 585
R650 B.n135 B.n134 585
R651 B.n133 B.n96 585
R652 B.n132 B.n131 585
R653 B.n130 B.n97 585
R654 B.n129 B.n128 585
R655 B.n127 B.n98 585
R656 B.n230 B.n63 585
R657 B.n232 B.n231 585
R658 B.n233 B.n62 585
R659 B.n235 B.n234 585
R660 B.n236 B.n61 585
R661 B.n238 B.n237 585
R662 B.n239 B.n60 585
R663 B.n241 B.n240 585
R664 B.n242 B.n59 585
R665 B.n244 B.n243 585
R666 B.n245 B.n58 585
R667 B.n247 B.n246 585
R668 B.n248 B.n57 585
R669 B.n250 B.n249 585
R670 B.n251 B.n56 585
R671 B.n253 B.n252 585
R672 B.n254 B.n55 585
R673 B.n256 B.n255 585
R674 B.n257 B.n54 585
R675 B.n259 B.n258 585
R676 B.n260 B.n53 585
R677 B.n262 B.n261 585
R678 B.n263 B.n52 585
R679 B.n265 B.n264 585
R680 B.n266 B.n51 585
R681 B.n268 B.n267 585
R682 B.n269 B.n50 585
R683 B.n271 B.n270 585
R684 B.n272 B.n49 585
R685 B.n274 B.n273 585
R686 B.n275 B.n48 585
R687 B.n277 B.n276 585
R688 B.n377 B.n376 585
R689 B.n375 B.n10 585
R690 B.n374 B.n373 585
R691 B.n372 B.n11 585
R692 B.n371 B.n370 585
R693 B.n369 B.n12 585
R694 B.n368 B.n367 585
R695 B.n366 B.n13 585
R696 B.n365 B.n364 585
R697 B.n363 B.n14 585
R698 B.n362 B.n361 585
R699 B.n360 B.n15 585
R700 B.n359 B.n358 585
R701 B.n357 B.n16 585
R702 B.n356 B.n355 585
R703 B.n354 B.n17 585
R704 B.n353 B.n352 585
R705 B.n351 B.n18 585
R706 B.n350 B.n349 585
R707 B.n348 B.n19 585
R708 B.n347 B.n346 585
R709 B.n345 B.n20 585
R710 B.n344 B.n343 585
R711 B.n342 B.n21 585
R712 B.n341 B.n340 585
R713 B.n339 B.n22 585
R714 B.n338 B.n337 585
R715 B.n336 B.n23 585
R716 B.n334 B.n333 585
R717 B.n332 B.n26 585
R718 B.n331 B.n330 585
R719 B.n329 B.n27 585
R720 B.n328 B.n327 585
R721 B.n326 B.n28 585
R722 B.n325 B.n324 585
R723 B.n323 B.n29 585
R724 B.n322 B.n321 585
R725 B.n320 B.n30 585
R726 B.n319 B.n318 585
R727 B.n317 B.n31 585
R728 B.n316 B.n315 585
R729 B.n314 B.n35 585
R730 B.n313 B.n312 585
R731 B.n311 B.n36 585
R732 B.n310 B.n309 585
R733 B.n308 B.n37 585
R734 B.n307 B.n306 585
R735 B.n305 B.n38 585
R736 B.n304 B.n303 585
R737 B.n302 B.n39 585
R738 B.n301 B.n300 585
R739 B.n299 B.n40 585
R740 B.n298 B.n297 585
R741 B.n296 B.n41 585
R742 B.n295 B.n294 585
R743 B.n293 B.n42 585
R744 B.n292 B.n291 585
R745 B.n290 B.n43 585
R746 B.n289 B.n288 585
R747 B.n287 B.n44 585
R748 B.n286 B.n285 585
R749 B.n284 B.n45 585
R750 B.n283 B.n282 585
R751 B.n281 B.n46 585
R752 B.n280 B.n279 585
R753 B.n278 B.n47 585
R754 B.n378 B.n9 585
R755 B.n380 B.n379 585
R756 B.n381 B.n8 585
R757 B.n383 B.n382 585
R758 B.n384 B.n7 585
R759 B.n386 B.n385 585
R760 B.n387 B.n6 585
R761 B.n389 B.n388 585
R762 B.n390 B.n5 585
R763 B.n392 B.n391 585
R764 B.n393 B.n4 585
R765 B.n395 B.n394 585
R766 B.n396 B.n3 585
R767 B.n398 B.n397 585
R768 B.n399 B.n0 585
R769 B.n2 B.n1 585
R770 B.n106 B.n105 585
R771 B.n108 B.n107 585
R772 B.n109 B.n104 585
R773 B.n111 B.n110 585
R774 B.n112 B.n103 585
R775 B.n114 B.n113 585
R776 B.n115 B.n102 585
R777 B.n117 B.n116 585
R778 B.n118 B.n101 585
R779 B.n120 B.n119 585
R780 B.n121 B.n100 585
R781 B.n123 B.n122 585
R782 B.n124 B.n99 585
R783 B.n126 B.n125 585
R784 B.n125 B.n98 478.086
R785 B.n230 B.n229 478.086
R786 B.n278 B.n277 478.086
R787 B.n376 B.n9 478.086
R788 B.n183 B.t4 302.962
R789 B.n32 B.t11 302.962
R790 B.n83 B.t7 302.962
R791 B.n24 B.t2 302.962
R792 B.n184 B.t5 293.265
R793 B.n33 B.t10 293.265
R794 B.n84 B.t8 293.265
R795 B.n25 B.t1 293.265
R796 B.n401 B.n400 256.663
R797 B.n400 B.n399 235.042
R798 B.n400 B.n2 235.042
R799 B.n129 B.n98 163.367
R800 B.n130 B.n129 163.367
R801 B.n131 B.n130 163.367
R802 B.n131 B.n96 163.367
R803 B.n135 B.n96 163.367
R804 B.n136 B.n135 163.367
R805 B.n137 B.n136 163.367
R806 B.n137 B.n94 163.367
R807 B.n141 B.n94 163.367
R808 B.n142 B.n141 163.367
R809 B.n143 B.n142 163.367
R810 B.n143 B.n92 163.367
R811 B.n147 B.n92 163.367
R812 B.n148 B.n147 163.367
R813 B.n149 B.n148 163.367
R814 B.n149 B.n90 163.367
R815 B.n153 B.n90 163.367
R816 B.n154 B.n153 163.367
R817 B.n155 B.n154 163.367
R818 B.n155 B.n88 163.367
R819 B.n159 B.n88 163.367
R820 B.n160 B.n159 163.367
R821 B.n161 B.n160 163.367
R822 B.n161 B.n86 163.367
R823 B.n165 B.n86 163.367
R824 B.n166 B.n165 163.367
R825 B.n167 B.n166 163.367
R826 B.n167 B.n82 163.367
R827 B.n172 B.n82 163.367
R828 B.n173 B.n172 163.367
R829 B.n174 B.n173 163.367
R830 B.n174 B.n80 163.367
R831 B.n178 B.n80 163.367
R832 B.n179 B.n178 163.367
R833 B.n180 B.n179 163.367
R834 B.n180 B.n78 163.367
R835 B.n187 B.n78 163.367
R836 B.n188 B.n187 163.367
R837 B.n189 B.n188 163.367
R838 B.n189 B.n76 163.367
R839 B.n193 B.n76 163.367
R840 B.n194 B.n193 163.367
R841 B.n195 B.n194 163.367
R842 B.n195 B.n74 163.367
R843 B.n199 B.n74 163.367
R844 B.n200 B.n199 163.367
R845 B.n201 B.n200 163.367
R846 B.n201 B.n72 163.367
R847 B.n205 B.n72 163.367
R848 B.n206 B.n205 163.367
R849 B.n207 B.n206 163.367
R850 B.n207 B.n70 163.367
R851 B.n211 B.n70 163.367
R852 B.n212 B.n211 163.367
R853 B.n213 B.n212 163.367
R854 B.n213 B.n68 163.367
R855 B.n217 B.n68 163.367
R856 B.n218 B.n217 163.367
R857 B.n219 B.n218 163.367
R858 B.n219 B.n66 163.367
R859 B.n223 B.n66 163.367
R860 B.n224 B.n223 163.367
R861 B.n225 B.n224 163.367
R862 B.n225 B.n64 163.367
R863 B.n229 B.n64 163.367
R864 B.n277 B.n48 163.367
R865 B.n273 B.n48 163.367
R866 B.n273 B.n272 163.367
R867 B.n272 B.n271 163.367
R868 B.n271 B.n50 163.367
R869 B.n267 B.n50 163.367
R870 B.n267 B.n266 163.367
R871 B.n266 B.n265 163.367
R872 B.n265 B.n52 163.367
R873 B.n261 B.n52 163.367
R874 B.n261 B.n260 163.367
R875 B.n260 B.n259 163.367
R876 B.n259 B.n54 163.367
R877 B.n255 B.n54 163.367
R878 B.n255 B.n254 163.367
R879 B.n254 B.n253 163.367
R880 B.n253 B.n56 163.367
R881 B.n249 B.n56 163.367
R882 B.n249 B.n248 163.367
R883 B.n248 B.n247 163.367
R884 B.n247 B.n58 163.367
R885 B.n243 B.n58 163.367
R886 B.n243 B.n242 163.367
R887 B.n242 B.n241 163.367
R888 B.n241 B.n60 163.367
R889 B.n237 B.n60 163.367
R890 B.n237 B.n236 163.367
R891 B.n236 B.n235 163.367
R892 B.n235 B.n62 163.367
R893 B.n231 B.n62 163.367
R894 B.n231 B.n230 163.367
R895 B.n376 B.n375 163.367
R896 B.n375 B.n374 163.367
R897 B.n374 B.n11 163.367
R898 B.n370 B.n11 163.367
R899 B.n370 B.n369 163.367
R900 B.n369 B.n368 163.367
R901 B.n368 B.n13 163.367
R902 B.n364 B.n13 163.367
R903 B.n364 B.n363 163.367
R904 B.n363 B.n362 163.367
R905 B.n362 B.n15 163.367
R906 B.n358 B.n15 163.367
R907 B.n358 B.n357 163.367
R908 B.n357 B.n356 163.367
R909 B.n356 B.n17 163.367
R910 B.n352 B.n17 163.367
R911 B.n352 B.n351 163.367
R912 B.n351 B.n350 163.367
R913 B.n350 B.n19 163.367
R914 B.n346 B.n19 163.367
R915 B.n346 B.n345 163.367
R916 B.n345 B.n344 163.367
R917 B.n344 B.n21 163.367
R918 B.n340 B.n21 163.367
R919 B.n340 B.n339 163.367
R920 B.n339 B.n338 163.367
R921 B.n338 B.n23 163.367
R922 B.n333 B.n23 163.367
R923 B.n333 B.n332 163.367
R924 B.n332 B.n331 163.367
R925 B.n331 B.n27 163.367
R926 B.n327 B.n27 163.367
R927 B.n327 B.n326 163.367
R928 B.n326 B.n325 163.367
R929 B.n325 B.n29 163.367
R930 B.n321 B.n29 163.367
R931 B.n321 B.n320 163.367
R932 B.n320 B.n319 163.367
R933 B.n319 B.n31 163.367
R934 B.n315 B.n31 163.367
R935 B.n315 B.n314 163.367
R936 B.n314 B.n313 163.367
R937 B.n313 B.n36 163.367
R938 B.n309 B.n36 163.367
R939 B.n309 B.n308 163.367
R940 B.n308 B.n307 163.367
R941 B.n307 B.n38 163.367
R942 B.n303 B.n38 163.367
R943 B.n303 B.n302 163.367
R944 B.n302 B.n301 163.367
R945 B.n301 B.n40 163.367
R946 B.n297 B.n40 163.367
R947 B.n297 B.n296 163.367
R948 B.n296 B.n295 163.367
R949 B.n295 B.n42 163.367
R950 B.n291 B.n42 163.367
R951 B.n291 B.n290 163.367
R952 B.n290 B.n289 163.367
R953 B.n289 B.n44 163.367
R954 B.n285 B.n44 163.367
R955 B.n285 B.n284 163.367
R956 B.n284 B.n283 163.367
R957 B.n283 B.n46 163.367
R958 B.n279 B.n46 163.367
R959 B.n279 B.n278 163.367
R960 B.n380 B.n9 163.367
R961 B.n381 B.n380 163.367
R962 B.n382 B.n381 163.367
R963 B.n382 B.n7 163.367
R964 B.n386 B.n7 163.367
R965 B.n387 B.n386 163.367
R966 B.n388 B.n387 163.367
R967 B.n388 B.n5 163.367
R968 B.n392 B.n5 163.367
R969 B.n393 B.n392 163.367
R970 B.n394 B.n393 163.367
R971 B.n394 B.n3 163.367
R972 B.n398 B.n3 163.367
R973 B.n399 B.n398 163.367
R974 B.n106 B.n2 163.367
R975 B.n107 B.n106 163.367
R976 B.n107 B.n104 163.367
R977 B.n111 B.n104 163.367
R978 B.n112 B.n111 163.367
R979 B.n113 B.n112 163.367
R980 B.n113 B.n102 163.367
R981 B.n117 B.n102 163.367
R982 B.n118 B.n117 163.367
R983 B.n119 B.n118 163.367
R984 B.n119 B.n100 163.367
R985 B.n123 B.n100 163.367
R986 B.n124 B.n123 163.367
R987 B.n125 B.n124 163.367
R988 B.n169 B.n84 59.5399
R989 B.n185 B.n184 59.5399
R990 B.n34 B.n33 59.5399
R991 B.n335 B.n25 59.5399
R992 B.n378 B.n377 31.0639
R993 B.n276 B.n47 31.0639
R994 B.n228 B.n63 31.0639
R995 B.n127 B.n126 31.0639
R996 B B.n401 18.0485
R997 B.n379 B.n378 10.6151
R998 B.n379 B.n8 10.6151
R999 B.n383 B.n8 10.6151
R1000 B.n384 B.n383 10.6151
R1001 B.n385 B.n384 10.6151
R1002 B.n385 B.n6 10.6151
R1003 B.n389 B.n6 10.6151
R1004 B.n390 B.n389 10.6151
R1005 B.n391 B.n390 10.6151
R1006 B.n391 B.n4 10.6151
R1007 B.n395 B.n4 10.6151
R1008 B.n396 B.n395 10.6151
R1009 B.n397 B.n396 10.6151
R1010 B.n397 B.n0 10.6151
R1011 B.n377 B.n10 10.6151
R1012 B.n373 B.n10 10.6151
R1013 B.n373 B.n372 10.6151
R1014 B.n372 B.n371 10.6151
R1015 B.n371 B.n12 10.6151
R1016 B.n367 B.n12 10.6151
R1017 B.n367 B.n366 10.6151
R1018 B.n366 B.n365 10.6151
R1019 B.n365 B.n14 10.6151
R1020 B.n361 B.n14 10.6151
R1021 B.n361 B.n360 10.6151
R1022 B.n360 B.n359 10.6151
R1023 B.n359 B.n16 10.6151
R1024 B.n355 B.n16 10.6151
R1025 B.n355 B.n354 10.6151
R1026 B.n354 B.n353 10.6151
R1027 B.n353 B.n18 10.6151
R1028 B.n349 B.n18 10.6151
R1029 B.n349 B.n348 10.6151
R1030 B.n348 B.n347 10.6151
R1031 B.n347 B.n20 10.6151
R1032 B.n343 B.n20 10.6151
R1033 B.n343 B.n342 10.6151
R1034 B.n342 B.n341 10.6151
R1035 B.n341 B.n22 10.6151
R1036 B.n337 B.n22 10.6151
R1037 B.n337 B.n336 10.6151
R1038 B.n334 B.n26 10.6151
R1039 B.n330 B.n26 10.6151
R1040 B.n330 B.n329 10.6151
R1041 B.n329 B.n328 10.6151
R1042 B.n328 B.n28 10.6151
R1043 B.n324 B.n28 10.6151
R1044 B.n324 B.n323 10.6151
R1045 B.n323 B.n322 10.6151
R1046 B.n322 B.n30 10.6151
R1047 B.n318 B.n317 10.6151
R1048 B.n317 B.n316 10.6151
R1049 B.n316 B.n35 10.6151
R1050 B.n312 B.n35 10.6151
R1051 B.n312 B.n311 10.6151
R1052 B.n311 B.n310 10.6151
R1053 B.n310 B.n37 10.6151
R1054 B.n306 B.n37 10.6151
R1055 B.n306 B.n305 10.6151
R1056 B.n305 B.n304 10.6151
R1057 B.n304 B.n39 10.6151
R1058 B.n300 B.n39 10.6151
R1059 B.n300 B.n299 10.6151
R1060 B.n299 B.n298 10.6151
R1061 B.n298 B.n41 10.6151
R1062 B.n294 B.n41 10.6151
R1063 B.n294 B.n293 10.6151
R1064 B.n293 B.n292 10.6151
R1065 B.n292 B.n43 10.6151
R1066 B.n288 B.n43 10.6151
R1067 B.n288 B.n287 10.6151
R1068 B.n287 B.n286 10.6151
R1069 B.n286 B.n45 10.6151
R1070 B.n282 B.n45 10.6151
R1071 B.n282 B.n281 10.6151
R1072 B.n281 B.n280 10.6151
R1073 B.n280 B.n47 10.6151
R1074 B.n276 B.n275 10.6151
R1075 B.n275 B.n274 10.6151
R1076 B.n274 B.n49 10.6151
R1077 B.n270 B.n49 10.6151
R1078 B.n270 B.n269 10.6151
R1079 B.n269 B.n268 10.6151
R1080 B.n268 B.n51 10.6151
R1081 B.n264 B.n51 10.6151
R1082 B.n264 B.n263 10.6151
R1083 B.n263 B.n262 10.6151
R1084 B.n262 B.n53 10.6151
R1085 B.n258 B.n53 10.6151
R1086 B.n258 B.n257 10.6151
R1087 B.n257 B.n256 10.6151
R1088 B.n256 B.n55 10.6151
R1089 B.n252 B.n55 10.6151
R1090 B.n252 B.n251 10.6151
R1091 B.n251 B.n250 10.6151
R1092 B.n250 B.n57 10.6151
R1093 B.n246 B.n57 10.6151
R1094 B.n246 B.n245 10.6151
R1095 B.n245 B.n244 10.6151
R1096 B.n244 B.n59 10.6151
R1097 B.n240 B.n59 10.6151
R1098 B.n240 B.n239 10.6151
R1099 B.n239 B.n238 10.6151
R1100 B.n238 B.n61 10.6151
R1101 B.n234 B.n61 10.6151
R1102 B.n234 B.n233 10.6151
R1103 B.n233 B.n232 10.6151
R1104 B.n232 B.n63 10.6151
R1105 B.n105 B.n1 10.6151
R1106 B.n108 B.n105 10.6151
R1107 B.n109 B.n108 10.6151
R1108 B.n110 B.n109 10.6151
R1109 B.n110 B.n103 10.6151
R1110 B.n114 B.n103 10.6151
R1111 B.n115 B.n114 10.6151
R1112 B.n116 B.n115 10.6151
R1113 B.n116 B.n101 10.6151
R1114 B.n120 B.n101 10.6151
R1115 B.n121 B.n120 10.6151
R1116 B.n122 B.n121 10.6151
R1117 B.n122 B.n99 10.6151
R1118 B.n126 B.n99 10.6151
R1119 B.n128 B.n127 10.6151
R1120 B.n128 B.n97 10.6151
R1121 B.n132 B.n97 10.6151
R1122 B.n133 B.n132 10.6151
R1123 B.n134 B.n133 10.6151
R1124 B.n134 B.n95 10.6151
R1125 B.n138 B.n95 10.6151
R1126 B.n139 B.n138 10.6151
R1127 B.n140 B.n139 10.6151
R1128 B.n140 B.n93 10.6151
R1129 B.n144 B.n93 10.6151
R1130 B.n145 B.n144 10.6151
R1131 B.n146 B.n145 10.6151
R1132 B.n146 B.n91 10.6151
R1133 B.n150 B.n91 10.6151
R1134 B.n151 B.n150 10.6151
R1135 B.n152 B.n151 10.6151
R1136 B.n152 B.n89 10.6151
R1137 B.n156 B.n89 10.6151
R1138 B.n157 B.n156 10.6151
R1139 B.n158 B.n157 10.6151
R1140 B.n158 B.n87 10.6151
R1141 B.n162 B.n87 10.6151
R1142 B.n163 B.n162 10.6151
R1143 B.n164 B.n163 10.6151
R1144 B.n164 B.n85 10.6151
R1145 B.n168 B.n85 10.6151
R1146 B.n171 B.n170 10.6151
R1147 B.n171 B.n81 10.6151
R1148 B.n175 B.n81 10.6151
R1149 B.n176 B.n175 10.6151
R1150 B.n177 B.n176 10.6151
R1151 B.n177 B.n79 10.6151
R1152 B.n181 B.n79 10.6151
R1153 B.n182 B.n181 10.6151
R1154 B.n186 B.n182 10.6151
R1155 B.n190 B.n77 10.6151
R1156 B.n191 B.n190 10.6151
R1157 B.n192 B.n191 10.6151
R1158 B.n192 B.n75 10.6151
R1159 B.n196 B.n75 10.6151
R1160 B.n197 B.n196 10.6151
R1161 B.n198 B.n197 10.6151
R1162 B.n198 B.n73 10.6151
R1163 B.n202 B.n73 10.6151
R1164 B.n203 B.n202 10.6151
R1165 B.n204 B.n203 10.6151
R1166 B.n204 B.n71 10.6151
R1167 B.n208 B.n71 10.6151
R1168 B.n209 B.n208 10.6151
R1169 B.n210 B.n209 10.6151
R1170 B.n210 B.n69 10.6151
R1171 B.n214 B.n69 10.6151
R1172 B.n215 B.n214 10.6151
R1173 B.n216 B.n215 10.6151
R1174 B.n216 B.n67 10.6151
R1175 B.n220 B.n67 10.6151
R1176 B.n221 B.n220 10.6151
R1177 B.n222 B.n221 10.6151
R1178 B.n222 B.n65 10.6151
R1179 B.n226 B.n65 10.6151
R1180 B.n227 B.n226 10.6151
R1181 B.n228 B.n227 10.6151
R1182 B.n84 B.n83 9.69747
R1183 B.n184 B.n183 9.69747
R1184 B.n33 B.n32 9.69747
R1185 B.n25 B.n24 9.69747
R1186 B.n336 B.n335 9.36635
R1187 B.n318 B.n34 9.36635
R1188 B.n169 B.n168 9.36635
R1189 B.n185 B.n77 9.36635
R1190 B.n401 B.n0 8.11757
R1191 B.n401 B.n1 8.11757
R1192 B.n335 B.n334 1.24928
R1193 B.n34 B.n30 1.24928
R1194 B.n170 B.n169 1.24928
R1195 B.n186 B.n185 1.24928
C0 w_n1470_n2450# VP 2.42501f
C1 w_n1470_n2450# B 5.18306f
C2 B VP 0.895012f
C3 VN VTAIL 1.28004f
C4 VN VDD1 0.14676f
C5 VDD2 VN 1.59498f
C6 w_n1470_n2450# VN 2.24133f
C7 VDD1 VTAIL 13.476099f
C8 VP VN 3.84348f
C9 B VN 0.600067f
C10 VDD2 VTAIL 13.5142f
C11 VDD2 VDD1 0.568086f
C12 w_n1470_n2450# VTAIL 3.0942f
C13 w_n1470_n2450# VDD1 0.946116f
C14 VP VTAIL 1.29415f
C15 VP VDD1 1.70857f
C16 B VTAIL 2.25892f
C17 B VDD1 0.784231f
C18 w_n1470_n2450# VDD2 0.959572f
C19 VDD2 VP 0.260519f
C20 VDD2 B 0.805126f
C21 VDD2 VSUBS 1.19451f
C22 VDD1 VSUBS 1.3872f
C23 VTAIL VSUBS 0.498117f
C24 VN VSUBS 3.20516f
C25 VP VSUBS 0.929143f
C26 B VSUBS 1.893959f
C27 w_n1470_n2450# VSUBS 44.752697f
C28 B.n0 VSUBS 0.00843f
C29 B.n1 VSUBS 0.00843f
C30 B.n2 VSUBS 0.012467f
C31 B.n3 VSUBS 0.009554f
C32 B.n4 VSUBS 0.009554f
C33 B.n5 VSUBS 0.009554f
C34 B.n6 VSUBS 0.009554f
C35 B.n7 VSUBS 0.009554f
C36 B.n8 VSUBS 0.009554f
C37 B.n9 VSUBS 0.021014f
C38 B.n10 VSUBS 0.009554f
C39 B.n11 VSUBS 0.009554f
C40 B.n12 VSUBS 0.009554f
C41 B.n13 VSUBS 0.009554f
C42 B.n14 VSUBS 0.009554f
C43 B.n15 VSUBS 0.009554f
C44 B.n16 VSUBS 0.009554f
C45 B.n17 VSUBS 0.009554f
C46 B.n18 VSUBS 0.009554f
C47 B.n19 VSUBS 0.009554f
C48 B.n20 VSUBS 0.009554f
C49 B.n21 VSUBS 0.009554f
C50 B.n22 VSUBS 0.009554f
C51 B.n23 VSUBS 0.009554f
C52 B.t1 VSUBS 0.157469f
C53 B.t2 VSUBS 0.164522f
C54 B.t0 VSUBS 0.067328f
C55 B.n24 VSUBS 0.245451f
C56 B.n25 VSUBS 0.23401f
C57 B.n26 VSUBS 0.009554f
C58 B.n27 VSUBS 0.009554f
C59 B.n28 VSUBS 0.009554f
C60 B.n29 VSUBS 0.009554f
C61 B.n30 VSUBS 0.005339f
C62 B.n31 VSUBS 0.009554f
C63 B.t10 VSUBS 0.157472f
C64 B.t11 VSUBS 0.164525f
C65 B.t9 VSUBS 0.067328f
C66 B.n32 VSUBS 0.245448f
C67 B.n33 VSUBS 0.234007f
C68 B.n34 VSUBS 0.022135f
C69 B.n35 VSUBS 0.009554f
C70 B.n36 VSUBS 0.009554f
C71 B.n37 VSUBS 0.009554f
C72 B.n38 VSUBS 0.009554f
C73 B.n39 VSUBS 0.009554f
C74 B.n40 VSUBS 0.009554f
C75 B.n41 VSUBS 0.009554f
C76 B.n42 VSUBS 0.009554f
C77 B.n43 VSUBS 0.009554f
C78 B.n44 VSUBS 0.009554f
C79 B.n45 VSUBS 0.009554f
C80 B.n46 VSUBS 0.009554f
C81 B.n47 VSUBS 0.022258f
C82 B.n48 VSUBS 0.009554f
C83 B.n49 VSUBS 0.009554f
C84 B.n50 VSUBS 0.009554f
C85 B.n51 VSUBS 0.009554f
C86 B.n52 VSUBS 0.009554f
C87 B.n53 VSUBS 0.009554f
C88 B.n54 VSUBS 0.009554f
C89 B.n55 VSUBS 0.009554f
C90 B.n56 VSUBS 0.009554f
C91 B.n57 VSUBS 0.009554f
C92 B.n58 VSUBS 0.009554f
C93 B.n59 VSUBS 0.009554f
C94 B.n60 VSUBS 0.009554f
C95 B.n61 VSUBS 0.009554f
C96 B.n62 VSUBS 0.009554f
C97 B.n63 VSUBS 0.022201f
C98 B.n64 VSUBS 0.009554f
C99 B.n65 VSUBS 0.009554f
C100 B.n66 VSUBS 0.009554f
C101 B.n67 VSUBS 0.009554f
C102 B.n68 VSUBS 0.009554f
C103 B.n69 VSUBS 0.009554f
C104 B.n70 VSUBS 0.009554f
C105 B.n71 VSUBS 0.009554f
C106 B.n72 VSUBS 0.009554f
C107 B.n73 VSUBS 0.009554f
C108 B.n74 VSUBS 0.009554f
C109 B.n75 VSUBS 0.009554f
C110 B.n76 VSUBS 0.009554f
C111 B.n77 VSUBS 0.008992f
C112 B.n78 VSUBS 0.009554f
C113 B.n79 VSUBS 0.009554f
C114 B.n80 VSUBS 0.009554f
C115 B.n81 VSUBS 0.009554f
C116 B.n82 VSUBS 0.009554f
C117 B.t8 VSUBS 0.157469f
C118 B.t7 VSUBS 0.164522f
C119 B.t6 VSUBS 0.067328f
C120 B.n83 VSUBS 0.245451f
C121 B.n84 VSUBS 0.23401f
C122 B.n85 VSUBS 0.009554f
C123 B.n86 VSUBS 0.009554f
C124 B.n87 VSUBS 0.009554f
C125 B.n88 VSUBS 0.009554f
C126 B.n89 VSUBS 0.009554f
C127 B.n90 VSUBS 0.009554f
C128 B.n91 VSUBS 0.009554f
C129 B.n92 VSUBS 0.009554f
C130 B.n93 VSUBS 0.009554f
C131 B.n94 VSUBS 0.009554f
C132 B.n95 VSUBS 0.009554f
C133 B.n96 VSUBS 0.009554f
C134 B.n97 VSUBS 0.009554f
C135 B.n98 VSUBS 0.022258f
C136 B.n99 VSUBS 0.009554f
C137 B.n100 VSUBS 0.009554f
C138 B.n101 VSUBS 0.009554f
C139 B.n102 VSUBS 0.009554f
C140 B.n103 VSUBS 0.009554f
C141 B.n104 VSUBS 0.009554f
C142 B.n105 VSUBS 0.009554f
C143 B.n106 VSUBS 0.009554f
C144 B.n107 VSUBS 0.009554f
C145 B.n108 VSUBS 0.009554f
C146 B.n109 VSUBS 0.009554f
C147 B.n110 VSUBS 0.009554f
C148 B.n111 VSUBS 0.009554f
C149 B.n112 VSUBS 0.009554f
C150 B.n113 VSUBS 0.009554f
C151 B.n114 VSUBS 0.009554f
C152 B.n115 VSUBS 0.009554f
C153 B.n116 VSUBS 0.009554f
C154 B.n117 VSUBS 0.009554f
C155 B.n118 VSUBS 0.009554f
C156 B.n119 VSUBS 0.009554f
C157 B.n120 VSUBS 0.009554f
C158 B.n121 VSUBS 0.009554f
C159 B.n122 VSUBS 0.009554f
C160 B.n123 VSUBS 0.009554f
C161 B.n124 VSUBS 0.009554f
C162 B.n125 VSUBS 0.021014f
C163 B.n126 VSUBS 0.021014f
C164 B.n127 VSUBS 0.022258f
C165 B.n128 VSUBS 0.009554f
C166 B.n129 VSUBS 0.009554f
C167 B.n130 VSUBS 0.009554f
C168 B.n131 VSUBS 0.009554f
C169 B.n132 VSUBS 0.009554f
C170 B.n133 VSUBS 0.009554f
C171 B.n134 VSUBS 0.009554f
C172 B.n135 VSUBS 0.009554f
C173 B.n136 VSUBS 0.009554f
C174 B.n137 VSUBS 0.009554f
C175 B.n138 VSUBS 0.009554f
C176 B.n139 VSUBS 0.009554f
C177 B.n140 VSUBS 0.009554f
C178 B.n141 VSUBS 0.009554f
C179 B.n142 VSUBS 0.009554f
C180 B.n143 VSUBS 0.009554f
C181 B.n144 VSUBS 0.009554f
C182 B.n145 VSUBS 0.009554f
C183 B.n146 VSUBS 0.009554f
C184 B.n147 VSUBS 0.009554f
C185 B.n148 VSUBS 0.009554f
C186 B.n149 VSUBS 0.009554f
C187 B.n150 VSUBS 0.009554f
C188 B.n151 VSUBS 0.009554f
C189 B.n152 VSUBS 0.009554f
C190 B.n153 VSUBS 0.009554f
C191 B.n154 VSUBS 0.009554f
C192 B.n155 VSUBS 0.009554f
C193 B.n156 VSUBS 0.009554f
C194 B.n157 VSUBS 0.009554f
C195 B.n158 VSUBS 0.009554f
C196 B.n159 VSUBS 0.009554f
C197 B.n160 VSUBS 0.009554f
C198 B.n161 VSUBS 0.009554f
C199 B.n162 VSUBS 0.009554f
C200 B.n163 VSUBS 0.009554f
C201 B.n164 VSUBS 0.009554f
C202 B.n165 VSUBS 0.009554f
C203 B.n166 VSUBS 0.009554f
C204 B.n167 VSUBS 0.009554f
C205 B.n168 VSUBS 0.008992f
C206 B.n169 VSUBS 0.022135f
C207 B.n170 VSUBS 0.005339f
C208 B.n171 VSUBS 0.009554f
C209 B.n172 VSUBS 0.009554f
C210 B.n173 VSUBS 0.009554f
C211 B.n174 VSUBS 0.009554f
C212 B.n175 VSUBS 0.009554f
C213 B.n176 VSUBS 0.009554f
C214 B.n177 VSUBS 0.009554f
C215 B.n178 VSUBS 0.009554f
C216 B.n179 VSUBS 0.009554f
C217 B.n180 VSUBS 0.009554f
C218 B.n181 VSUBS 0.009554f
C219 B.n182 VSUBS 0.009554f
C220 B.t5 VSUBS 0.157472f
C221 B.t4 VSUBS 0.164525f
C222 B.t3 VSUBS 0.067328f
C223 B.n183 VSUBS 0.245448f
C224 B.n184 VSUBS 0.234007f
C225 B.n185 VSUBS 0.022135f
C226 B.n186 VSUBS 0.005339f
C227 B.n187 VSUBS 0.009554f
C228 B.n188 VSUBS 0.009554f
C229 B.n189 VSUBS 0.009554f
C230 B.n190 VSUBS 0.009554f
C231 B.n191 VSUBS 0.009554f
C232 B.n192 VSUBS 0.009554f
C233 B.n193 VSUBS 0.009554f
C234 B.n194 VSUBS 0.009554f
C235 B.n195 VSUBS 0.009554f
C236 B.n196 VSUBS 0.009554f
C237 B.n197 VSUBS 0.009554f
C238 B.n198 VSUBS 0.009554f
C239 B.n199 VSUBS 0.009554f
C240 B.n200 VSUBS 0.009554f
C241 B.n201 VSUBS 0.009554f
C242 B.n202 VSUBS 0.009554f
C243 B.n203 VSUBS 0.009554f
C244 B.n204 VSUBS 0.009554f
C245 B.n205 VSUBS 0.009554f
C246 B.n206 VSUBS 0.009554f
C247 B.n207 VSUBS 0.009554f
C248 B.n208 VSUBS 0.009554f
C249 B.n209 VSUBS 0.009554f
C250 B.n210 VSUBS 0.009554f
C251 B.n211 VSUBS 0.009554f
C252 B.n212 VSUBS 0.009554f
C253 B.n213 VSUBS 0.009554f
C254 B.n214 VSUBS 0.009554f
C255 B.n215 VSUBS 0.009554f
C256 B.n216 VSUBS 0.009554f
C257 B.n217 VSUBS 0.009554f
C258 B.n218 VSUBS 0.009554f
C259 B.n219 VSUBS 0.009554f
C260 B.n220 VSUBS 0.009554f
C261 B.n221 VSUBS 0.009554f
C262 B.n222 VSUBS 0.009554f
C263 B.n223 VSUBS 0.009554f
C264 B.n224 VSUBS 0.009554f
C265 B.n225 VSUBS 0.009554f
C266 B.n226 VSUBS 0.009554f
C267 B.n227 VSUBS 0.009554f
C268 B.n228 VSUBS 0.021072f
C269 B.n229 VSUBS 0.022258f
C270 B.n230 VSUBS 0.021014f
C271 B.n231 VSUBS 0.009554f
C272 B.n232 VSUBS 0.009554f
C273 B.n233 VSUBS 0.009554f
C274 B.n234 VSUBS 0.009554f
C275 B.n235 VSUBS 0.009554f
C276 B.n236 VSUBS 0.009554f
C277 B.n237 VSUBS 0.009554f
C278 B.n238 VSUBS 0.009554f
C279 B.n239 VSUBS 0.009554f
C280 B.n240 VSUBS 0.009554f
C281 B.n241 VSUBS 0.009554f
C282 B.n242 VSUBS 0.009554f
C283 B.n243 VSUBS 0.009554f
C284 B.n244 VSUBS 0.009554f
C285 B.n245 VSUBS 0.009554f
C286 B.n246 VSUBS 0.009554f
C287 B.n247 VSUBS 0.009554f
C288 B.n248 VSUBS 0.009554f
C289 B.n249 VSUBS 0.009554f
C290 B.n250 VSUBS 0.009554f
C291 B.n251 VSUBS 0.009554f
C292 B.n252 VSUBS 0.009554f
C293 B.n253 VSUBS 0.009554f
C294 B.n254 VSUBS 0.009554f
C295 B.n255 VSUBS 0.009554f
C296 B.n256 VSUBS 0.009554f
C297 B.n257 VSUBS 0.009554f
C298 B.n258 VSUBS 0.009554f
C299 B.n259 VSUBS 0.009554f
C300 B.n260 VSUBS 0.009554f
C301 B.n261 VSUBS 0.009554f
C302 B.n262 VSUBS 0.009554f
C303 B.n263 VSUBS 0.009554f
C304 B.n264 VSUBS 0.009554f
C305 B.n265 VSUBS 0.009554f
C306 B.n266 VSUBS 0.009554f
C307 B.n267 VSUBS 0.009554f
C308 B.n268 VSUBS 0.009554f
C309 B.n269 VSUBS 0.009554f
C310 B.n270 VSUBS 0.009554f
C311 B.n271 VSUBS 0.009554f
C312 B.n272 VSUBS 0.009554f
C313 B.n273 VSUBS 0.009554f
C314 B.n274 VSUBS 0.009554f
C315 B.n275 VSUBS 0.009554f
C316 B.n276 VSUBS 0.021014f
C317 B.n277 VSUBS 0.021014f
C318 B.n278 VSUBS 0.022258f
C319 B.n279 VSUBS 0.009554f
C320 B.n280 VSUBS 0.009554f
C321 B.n281 VSUBS 0.009554f
C322 B.n282 VSUBS 0.009554f
C323 B.n283 VSUBS 0.009554f
C324 B.n284 VSUBS 0.009554f
C325 B.n285 VSUBS 0.009554f
C326 B.n286 VSUBS 0.009554f
C327 B.n287 VSUBS 0.009554f
C328 B.n288 VSUBS 0.009554f
C329 B.n289 VSUBS 0.009554f
C330 B.n290 VSUBS 0.009554f
C331 B.n291 VSUBS 0.009554f
C332 B.n292 VSUBS 0.009554f
C333 B.n293 VSUBS 0.009554f
C334 B.n294 VSUBS 0.009554f
C335 B.n295 VSUBS 0.009554f
C336 B.n296 VSUBS 0.009554f
C337 B.n297 VSUBS 0.009554f
C338 B.n298 VSUBS 0.009554f
C339 B.n299 VSUBS 0.009554f
C340 B.n300 VSUBS 0.009554f
C341 B.n301 VSUBS 0.009554f
C342 B.n302 VSUBS 0.009554f
C343 B.n303 VSUBS 0.009554f
C344 B.n304 VSUBS 0.009554f
C345 B.n305 VSUBS 0.009554f
C346 B.n306 VSUBS 0.009554f
C347 B.n307 VSUBS 0.009554f
C348 B.n308 VSUBS 0.009554f
C349 B.n309 VSUBS 0.009554f
C350 B.n310 VSUBS 0.009554f
C351 B.n311 VSUBS 0.009554f
C352 B.n312 VSUBS 0.009554f
C353 B.n313 VSUBS 0.009554f
C354 B.n314 VSUBS 0.009554f
C355 B.n315 VSUBS 0.009554f
C356 B.n316 VSUBS 0.009554f
C357 B.n317 VSUBS 0.009554f
C358 B.n318 VSUBS 0.008992f
C359 B.n319 VSUBS 0.009554f
C360 B.n320 VSUBS 0.009554f
C361 B.n321 VSUBS 0.009554f
C362 B.n322 VSUBS 0.009554f
C363 B.n323 VSUBS 0.009554f
C364 B.n324 VSUBS 0.009554f
C365 B.n325 VSUBS 0.009554f
C366 B.n326 VSUBS 0.009554f
C367 B.n327 VSUBS 0.009554f
C368 B.n328 VSUBS 0.009554f
C369 B.n329 VSUBS 0.009554f
C370 B.n330 VSUBS 0.009554f
C371 B.n331 VSUBS 0.009554f
C372 B.n332 VSUBS 0.009554f
C373 B.n333 VSUBS 0.009554f
C374 B.n334 VSUBS 0.005339f
C375 B.n335 VSUBS 0.022135f
C376 B.n336 VSUBS 0.008992f
C377 B.n337 VSUBS 0.009554f
C378 B.n338 VSUBS 0.009554f
C379 B.n339 VSUBS 0.009554f
C380 B.n340 VSUBS 0.009554f
C381 B.n341 VSUBS 0.009554f
C382 B.n342 VSUBS 0.009554f
C383 B.n343 VSUBS 0.009554f
C384 B.n344 VSUBS 0.009554f
C385 B.n345 VSUBS 0.009554f
C386 B.n346 VSUBS 0.009554f
C387 B.n347 VSUBS 0.009554f
C388 B.n348 VSUBS 0.009554f
C389 B.n349 VSUBS 0.009554f
C390 B.n350 VSUBS 0.009554f
C391 B.n351 VSUBS 0.009554f
C392 B.n352 VSUBS 0.009554f
C393 B.n353 VSUBS 0.009554f
C394 B.n354 VSUBS 0.009554f
C395 B.n355 VSUBS 0.009554f
C396 B.n356 VSUBS 0.009554f
C397 B.n357 VSUBS 0.009554f
C398 B.n358 VSUBS 0.009554f
C399 B.n359 VSUBS 0.009554f
C400 B.n360 VSUBS 0.009554f
C401 B.n361 VSUBS 0.009554f
C402 B.n362 VSUBS 0.009554f
C403 B.n363 VSUBS 0.009554f
C404 B.n364 VSUBS 0.009554f
C405 B.n365 VSUBS 0.009554f
C406 B.n366 VSUBS 0.009554f
C407 B.n367 VSUBS 0.009554f
C408 B.n368 VSUBS 0.009554f
C409 B.n369 VSUBS 0.009554f
C410 B.n370 VSUBS 0.009554f
C411 B.n371 VSUBS 0.009554f
C412 B.n372 VSUBS 0.009554f
C413 B.n373 VSUBS 0.009554f
C414 B.n374 VSUBS 0.009554f
C415 B.n375 VSUBS 0.009554f
C416 B.n376 VSUBS 0.022258f
C417 B.n377 VSUBS 0.022258f
C418 B.n378 VSUBS 0.021014f
C419 B.n379 VSUBS 0.009554f
C420 B.n380 VSUBS 0.009554f
C421 B.n381 VSUBS 0.009554f
C422 B.n382 VSUBS 0.009554f
C423 B.n383 VSUBS 0.009554f
C424 B.n384 VSUBS 0.009554f
C425 B.n385 VSUBS 0.009554f
C426 B.n386 VSUBS 0.009554f
C427 B.n387 VSUBS 0.009554f
C428 B.n388 VSUBS 0.009554f
C429 B.n389 VSUBS 0.009554f
C430 B.n390 VSUBS 0.009554f
C431 B.n391 VSUBS 0.009554f
C432 B.n392 VSUBS 0.009554f
C433 B.n393 VSUBS 0.009554f
C434 B.n394 VSUBS 0.009554f
C435 B.n395 VSUBS 0.009554f
C436 B.n396 VSUBS 0.009554f
C437 B.n397 VSUBS 0.009554f
C438 B.n398 VSUBS 0.009554f
C439 B.n399 VSUBS 0.012467f
C440 B.n400 VSUBS 0.01328f
C441 B.n401 VSUBS 0.026409f
C442 VDD1.t7 VSUBS 0.199697f
C443 VDD1.t0 VSUBS 0.199697f
C444 VDD1.n0 VSUBS 1.39867f
C445 VDD1.t5 VSUBS 0.199697f
C446 VDD1.t4 VSUBS 0.199697f
C447 VDD1.n1 VSUBS 1.39774f
C448 VDD1.t3 VSUBS 0.199697f
C449 VDD1.t1 VSUBS 0.199697f
C450 VDD1.n2 VSUBS 1.39774f
C451 VDD1.n3 VSUBS 2.85884f
C452 VDD1.t2 VSUBS 0.199697f
C453 VDD1.t6 VSUBS 0.199697f
C454 VDD1.n4 VSUBS 1.39647f
C455 VDD1.n5 VSUBS 2.72615f
C456 VP.n0 VSUBS 0.055229f
C457 VP.t4 VSUBS 0.197692f
C458 VP.t3 VSUBS 0.197692f
C459 VP.t2 VSUBS 0.200297f
C460 VP.n1 VSUBS 0.116175f
C461 VP.t5 VSUBS 0.197692f
C462 VP.t7 VSUBS 0.197692f
C463 VP.t0 VSUBS 0.200297f
C464 VP.n2 VSUBS 0.10657f
C465 VP.n3 VSUBS 0.093506f
C466 VP.n4 VSUBS 0.018321f
C467 VP.n5 VSUBS 0.093506f
C468 VP.t1 VSUBS 0.200297f
C469 VP.n6 VSUBS 0.106499f
C470 VP.n7 VSUBS 1.74192f
C471 VP.n8 VSUBS 1.79697f
C472 VP.n9 VSUBS 0.106499f
C473 VP.n10 VSUBS 0.093506f
C474 VP.n11 VSUBS 0.018321f
C475 VP.n12 VSUBS 0.093506f
C476 VP.t6 VSUBS 0.200297f
C477 VP.n13 VSUBS 0.106499f
C478 VP.n14 VSUBS 0.0428f
C479 VTAIL.t5 VSUBS 0.184566f
C480 VTAIL.t6 VSUBS 0.184566f
C481 VTAIL.n0 VSUBS 1.15836f
C482 VTAIL.n1 VSUBS 0.684862f
C483 VTAIL.n2 VSUBS 0.03517f
C484 VTAIL.n3 VSUBS 0.03152f
C485 VTAIL.n4 VSUBS 0.016937f
C486 VTAIL.n5 VSUBS 0.040034f
C487 VTAIL.n6 VSUBS 0.017934f
C488 VTAIL.n7 VSUBS 0.03152f
C489 VTAIL.n8 VSUBS 0.016937f
C490 VTAIL.n9 VSUBS 0.040034f
C491 VTAIL.n10 VSUBS 0.017934f
C492 VTAIL.n11 VSUBS 0.03152f
C493 VTAIL.n12 VSUBS 0.016937f
C494 VTAIL.n13 VSUBS 0.030025f
C495 VTAIL.n14 VSUBS 0.025466f
C496 VTAIL.t12 VSUBS 0.085458f
C497 VTAIL.n15 VSUBS 0.151964f
C498 VTAIL.n16 VSUBS 0.925844f
C499 VTAIL.n17 VSUBS 0.016937f
C500 VTAIL.n18 VSUBS 0.017934f
C501 VTAIL.n19 VSUBS 0.040034f
C502 VTAIL.n20 VSUBS 0.040034f
C503 VTAIL.n21 VSUBS 0.017934f
C504 VTAIL.n22 VSUBS 0.016937f
C505 VTAIL.n23 VSUBS 0.03152f
C506 VTAIL.n24 VSUBS 0.03152f
C507 VTAIL.n25 VSUBS 0.016937f
C508 VTAIL.n26 VSUBS 0.017934f
C509 VTAIL.n27 VSUBS 0.040034f
C510 VTAIL.n28 VSUBS 0.040034f
C511 VTAIL.n29 VSUBS 0.017934f
C512 VTAIL.n30 VSUBS 0.016937f
C513 VTAIL.n31 VSUBS 0.03152f
C514 VTAIL.n32 VSUBS 0.03152f
C515 VTAIL.n33 VSUBS 0.016937f
C516 VTAIL.n34 VSUBS 0.017934f
C517 VTAIL.n35 VSUBS 0.040034f
C518 VTAIL.n36 VSUBS 0.098743f
C519 VTAIL.n37 VSUBS 0.017934f
C520 VTAIL.n38 VSUBS 0.016937f
C521 VTAIL.n39 VSUBS 0.071564f
C522 VTAIL.n40 VSUBS 0.049698f
C523 VTAIL.n41 VSUBS 0.117685f
C524 VTAIL.n42 VSUBS 0.03517f
C525 VTAIL.n43 VSUBS 0.03152f
C526 VTAIL.n44 VSUBS 0.016937f
C527 VTAIL.n45 VSUBS 0.040034f
C528 VTAIL.n46 VSUBS 0.017934f
C529 VTAIL.n47 VSUBS 0.03152f
C530 VTAIL.n48 VSUBS 0.016937f
C531 VTAIL.n49 VSUBS 0.040034f
C532 VTAIL.n50 VSUBS 0.017934f
C533 VTAIL.n51 VSUBS 0.03152f
C534 VTAIL.n52 VSUBS 0.016937f
C535 VTAIL.n53 VSUBS 0.030025f
C536 VTAIL.n54 VSUBS 0.025466f
C537 VTAIL.t0 VSUBS 0.085458f
C538 VTAIL.n55 VSUBS 0.151964f
C539 VTAIL.n56 VSUBS 0.925844f
C540 VTAIL.n57 VSUBS 0.016937f
C541 VTAIL.n58 VSUBS 0.017934f
C542 VTAIL.n59 VSUBS 0.040034f
C543 VTAIL.n60 VSUBS 0.040034f
C544 VTAIL.n61 VSUBS 0.017934f
C545 VTAIL.n62 VSUBS 0.016937f
C546 VTAIL.n63 VSUBS 0.03152f
C547 VTAIL.n64 VSUBS 0.03152f
C548 VTAIL.n65 VSUBS 0.016937f
C549 VTAIL.n66 VSUBS 0.017934f
C550 VTAIL.n67 VSUBS 0.040034f
C551 VTAIL.n68 VSUBS 0.040034f
C552 VTAIL.n69 VSUBS 0.017934f
C553 VTAIL.n70 VSUBS 0.016937f
C554 VTAIL.n71 VSUBS 0.03152f
C555 VTAIL.n72 VSUBS 0.03152f
C556 VTAIL.n73 VSUBS 0.016937f
C557 VTAIL.n74 VSUBS 0.017934f
C558 VTAIL.n75 VSUBS 0.040034f
C559 VTAIL.n76 VSUBS 0.098743f
C560 VTAIL.n77 VSUBS 0.017934f
C561 VTAIL.n78 VSUBS 0.016937f
C562 VTAIL.n79 VSUBS 0.071564f
C563 VTAIL.n80 VSUBS 0.049698f
C564 VTAIL.n81 VSUBS 0.117685f
C565 VTAIL.t13 VSUBS 0.184566f
C566 VTAIL.t14 VSUBS 0.184566f
C567 VTAIL.n82 VSUBS 1.15836f
C568 VTAIL.n83 VSUBS 0.72273f
C569 VTAIL.n84 VSUBS 0.03517f
C570 VTAIL.n85 VSUBS 0.03152f
C571 VTAIL.n86 VSUBS 0.016937f
C572 VTAIL.n87 VSUBS 0.040034f
C573 VTAIL.n88 VSUBS 0.017934f
C574 VTAIL.n89 VSUBS 0.03152f
C575 VTAIL.n90 VSUBS 0.016937f
C576 VTAIL.n91 VSUBS 0.040034f
C577 VTAIL.n92 VSUBS 0.017934f
C578 VTAIL.n93 VSUBS 0.03152f
C579 VTAIL.n94 VSUBS 0.016937f
C580 VTAIL.n95 VSUBS 0.030025f
C581 VTAIL.n96 VSUBS 0.025466f
C582 VTAIL.t1 VSUBS 0.085458f
C583 VTAIL.n97 VSUBS 0.151964f
C584 VTAIL.n98 VSUBS 0.925844f
C585 VTAIL.n99 VSUBS 0.016937f
C586 VTAIL.n100 VSUBS 0.017934f
C587 VTAIL.n101 VSUBS 0.040034f
C588 VTAIL.n102 VSUBS 0.040034f
C589 VTAIL.n103 VSUBS 0.017934f
C590 VTAIL.n104 VSUBS 0.016937f
C591 VTAIL.n105 VSUBS 0.03152f
C592 VTAIL.n106 VSUBS 0.03152f
C593 VTAIL.n107 VSUBS 0.016937f
C594 VTAIL.n108 VSUBS 0.017934f
C595 VTAIL.n109 VSUBS 0.040034f
C596 VTAIL.n110 VSUBS 0.040034f
C597 VTAIL.n111 VSUBS 0.017934f
C598 VTAIL.n112 VSUBS 0.016937f
C599 VTAIL.n113 VSUBS 0.03152f
C600 VTAIL.n114 VSUBS 0.03152f
C601 VTAIL.n115 VSUBS 0.016937f
C602 VTAIL.n116 VSUBS 0.017934f
C603 VTAIL.n117 VSUBS 0.040034f
C604 VTAIL.n118 VSUBS 0.098743f
C605 VTAIL.n119 VSUBS 0.017934f
C606 VTAIL.n120 VSUBS 0.016937f
C607 VTAIL.n121 VSUBS 0.071564f
C608 VTAIL.n122 VSUBS 0.049698f
C609 VTAIL.n123 VSUBS 1.19068f
C610 VTAIL.n124 VSUBS 0.03517f
C611 VTAIL.n125 VSUBS 0.03152f
C612 VTAIL.n126 VSUBS 0.016937f
C613 VTAIL.n127 VSUBS 0.040034f
C614 VTAIL.n128 VSUBS 0.017934f
C615 VTAIL.n129 VSUBS 0.03152f
C616 VTAIL.n130 VSUBS 0.016937f
C617 VTAIL.n131 VSUBS 0.040034f
C618 VTAIL.n132 VSUBS 0.017934f
C619 VTAIL.n133 VSUBS 0.03152f
C620 VTAIL.n134 VSUBS 0.016937f
C621 VTAIL.n135 VSUBS 0.030025f
C622 VTAIL.n136 VSUBS 0.025466f
C623 VTAIL.t9 VSUBS 0.085458f
C624 VTAIL.n137 VSUBS 0.151964f
C625 VTAIL.n138 VSUBS 0.925844f
C626 VTAIL.n139 VSUBS 0.016937f
C627 VTAIL.n140 VSUBS 0.017934f
C628 VTAIL.n141 VSUBS 0.040034f
C629 VTAIL.n142 VSUBS 0.040034f
C630 VTAIL.n143 VSUBS 0.017934f
C631 VTAIL.n144 VSUBS 0.016937f
C632 VTAIL.n145 VSUBS 0.03152f
C633 VTAIL.n146 VSUBS 0.03152f
C634 VTAIL.n147 VSUBS 0.016937f
C635 VTAIL.n148 VSUBS 0.017934f
C636 VTAIL.n149 VSUBS 0.040034f
C637 VTAIL.n150 VSUBS 0.040034f
C638 VTAIL.n151 VSUBS 0.017934f
C639 VTAIL.n152 VSUBS 0.016937f
C640 VTAIL.n153 VSUBS 0.03152f
C641 VTAIL.n154 VSUBS 0.03152f
C642 VTAIL.n155 VSUBS 0.016937f
C643 VTAIL.n156 VSUBS 0.017934f
C644 VTAIL.n157 VSUBS 0.040034f
C645 VTAIL.n158 VSUBS 0.098743f
C646 VTAIL.n159 VSUBS 0.017934f
C647 VTAIL.n160 VSUBS 0.016937f
C648 VTAIL.n161 VSUBS 0.071564f
C649 VTAIL.n162 VSUBS 0.049698f
C650 VTAIL.n163 VSUBS 1.19068f
C651 VTAIL.t7 VSUBS 0.184566f
C652 VTAIL.t11 VSUBS 0.184566f
C653 VTAIL.n164 VSUBS 1.15837f
C654 VTAIL.n165 VSUBS 0.722721f
C655 VTAIL.n166 VSUBS 0.03517f
C656 VTAIL.n167 VSUBS 0.03152f
C657 VTAIL.n168 VSUBS 0.016937f
C658 VTAIL.n169 VSUBS 0.040034f
C659 VTAIL.n170 VSUBS 0.017934f
C660 VTAIL.n171 VSUBS 0.03152f
C661 VTAIL.n172 VSUBS 0.016937f
C662 VTAIL.n173 VSUBS 0.040034f
C663 VTAIL.n174 VSUBS 0.017934f
C664 VTAIL.n175 VSUBS 0.03152f
C665 VTAIL.n176 VSUBS 0.016937f
C666 VTAIL.n177 VSUBS 0.030025f
C667 VTAIL.n178 VSUBS 0.025466f
C668 VTAIL.t10 VSUBS 0.085458f
C669 VTAIL.n179 VSUBS 0.151964f
C670 VTAIL.n180 VSUBS 0.925844f
C671 VTAIL.n181 VSUBS 0.016937f
C672 VTAIL.n182 VSUBS 0.017934f
C673 VTAIL.n183 VSUBS 0.040034f
C674 VTAIL.n184 VSUBS 0.040034f
C675 VTAIL.n185 VSUBS 0.017934f
C676 VTAIL.n186 VSUBS 0.016937f
C677 VTAIL.n187 VSUBS 0.03152f
C678 VTAIL.n188 VSUBS 0.03152f
C679 VTAIL.n189 VSUBS 0.016937f
C680 VTAIL.n190 VSUBS 0.017934f
C681 VTAIL.n191 VSUBS 0.040034f
C682 VTAIL.n192 VSUBS 0.040034f
C683 VTAIL.n193 VSUBS 0.017934f
C684 VTAIL.n194 VSUBS 0.016937f
C685 VTAIL.n195 VSUBS 0.03152f
C686 VTAIL.n196 VSUBS 0.03152f
C687 VTAIL.n197 VSUBS 0.016937f
C688 VTAIL.n198 VSUBS 0.017934f
C689 VTAIL.n199 VSUBS 0.040034f
C690 VTAIL.n200 VSUBS 0.098743f
C691 VTAIL.n201 VSUBS 0.017934f
C692 VTAIL.n202 VSUBS 0.016937f
C693 VTAIL.n203 VSUBS 0.071564f
C694 VTAIL.n204 VSUBS 0.049698f
C695 VTAIL.n205 VSUBS 0.117685f
C696 VTAIL.n206 VSUBS 0.03517f
C697 VTAIL.n207 VSUBS 0.03152f
C698 VTAIL.n208 VSUBS 0.016937f
C699 VTAIL.n209 VSUBS 0.040034f
C700 VTAIL.n210 VSUBS 0.017934f
C701 VTAIL.n211 VSUBS 0.03152f
C702 VTAIL.n212 VSUBS 0.016937f
C703 VTAIL.n213 VSUBS 0.040034f
C704 VTAIL.n214 VSUBS 0.017934f
C705 VTAIL.n215 VSUBS 0.03152f
C706 VTAIL.n216 VSUBS 0.016937f
C707 VTAIL.n217 VSUBS 0.030025f
C708 VTAIL.n218 VSUBS 0.025466f
C709 VTAIL.t2 VSUBS 0.085458f
C710 VTAIL.n219 VSUBS 0.151964f
C711 VTAIL.n220 VSUBS 0.925844f
C712 VTAIL.n221 VSUBS 0.016937f
C713 VTAIL.n222 VSUBS 0.017934f
C714 VTAIL.n223 VSUBS 0.040034f
C715 VTAIL.n224 VSUBS 0.040034f
C716 VTAIL.n225 VSUBS 0.017934f
C717 VTAIL.n226 VSUBS 0.016937f
C718 VTAIL.n227 VSUBS 0.03152f
C719 VTAIL.n228 VSUBS 0.03152f
C720 VTAIL.n229 VSUBS 0.016937f
C721 VTAIL.n230 VSUBS 0.017934f
C722 VTAIL.n231 VSUBS 0.040034f
C723 VTAIL.n232 VSUBS 0.040034f
C724 VTAIL.n233 VSUBS 0.017934f
C725 VTAIL.n234 VSUBS 0.016937f
C726 VTAIL.n235 VSUBS 0.03152f
C727 VTAIL.n236 VSUBS 0.03152f
C728 VTAIL.n237 VSUBS 0.016937f
C729 VTAIL.n238 VSUBS 0.017934f
C730 VTAIL.n239 VSUBS 0.040034f
C731 VTAIL.n240 VSUBS 0.098743f
C732 VTAIL.n241 VSUBS 0.017934f
C733 VTAIL.n242 VSUBS 0.016937f
C734 VTAIL.n243 VSUBS 0.071564f
C735 VTAIL.n244 VSUBS 0.049698f
C736 VTAIL.n245 VSUBS 0.117685f
C737 VTAIL.t3 VSUBS 0.184566f
C738 VTAIL.t15 VSUBS 0.184566f
C739 VTAIL.n246 VSUBS 1.15837f
C740 VTAIL.n247 VSUBS 0.722721f
C741 VTAIL.n248 VSUBS 0.03517f
C742 VTAIL.n249 VSUBS 0.03152f
C743 VTAIL.n250 VSUBS 0.016937f
C744 VTAIL.n251 VSUBS 0.040034f
C745 VTAIL.n252 VSUBS 0.017934f
C746 VTAIL.n253 VSUBS 0.03152f
C747 VTAIL.n254 VSUBS 0.016937f
C748 VTAIL.n255 VSUBS 0.040034f
C749 VTAIL.n256 VSUBS 0.017934f
C750 VTAIL.n257 VSUBS 0.03152f
C751 VTAIL.n258 VSUBS 0.016937f
C752 VTAIL.n259 VSUBS 0.030025f
C753 VTAIL.n260 VSUBS 0.025466f
C754 VTAIL.t4 VSUBS 0.085458f
C755 VTAIL.n261 VSUBS 0.151964f
C756 VTAIL.n262 VSUBS 0.925844f
C757 VTAIL.n263 VSUBS 0.016937f
C758 VTAIL.n264 VSUBS 0.017934f
C759 VTAIL.n265 VSUBS 0.040034f
C760 VTAIL.n266 VSUBS 0.040034f
C761 VTAIL.n267 VSUBS 0.017934f
C762 VTAIL.n268 VSUBS 0.016937f
C763 VTAIL.n269 VSUBS 0.03152f
C764 VTAIL.n270 VSUBS 0.03152f
C765 VTAIL.n271 VSUBS 0.016937f
C766 VTAIL.n272 VSUBS 0.017934f
C767 VTAIL.n273 VSUBS 0.040034f
C768 VTAIL.n274 VSUBS 0.040034f
C769 VTAIL.n275 VSUBS 0.017934f
C770 VTAIL.n276 VSUBS 0.016937f
C771 VTAIL.n277 VSUBS 0.03152f
C772 VTAIL.n278 VSUBS 0.03152f
C773 VTAIL.n279 VSUBS 0.016937f
C774 VTAIL.n280 VSUBS 0.017934f
C775 VTAIL.n281 VSUBS 0.040034f
C776 VTAIL.n282 VSUBS 0.098743f
C777 VTAIL.n283 VSUBS 0.017934f
C778 VTAIL.n284 VSUBS 0.016937f
C779 VTAIL.n285 VSUBS 0.071564f
C780 VTAIL.n286 VSUBS 0.049698f
C781 VTAIL.n287 VSUBS 1.19068f
C782 VTAIL.n288 VSUBS 0.03517f
C783 VTAIL.n289 VSUBS 0.03152f
C784 VTAIL.n290 VSUBS 0.016937f
C785 VTAIL.n291 VSUBS 0.040034f
C786 VTAIL.n292 VSUBS 0.017934f
C787 VTAIL.n293 VSUBS 0.03152f
C788 VTAIL.n294 VSUBS 0.016937f
C789 VTAIL.n295 VSUBS 0.040034f
C790 VTAIL.n296 VSUBS 0.017934f
C791 VTAIL.n297 VSUBS 0.03152f
C792 VTAIL.n298 VSUBS 0.016937f
C793 VTAIL.n299 VSUBS 0.030025f
C794 VTAIL.n300 VSUBS 0.025466f
C795 VTAIL.t8 VSUBS 0.085458f
C796 VTAIL.n301 VSUBS 0.151964f
C797 VTAIL.n302 VSUBS 0.925844f
C798 VTAIL.n303 VSUBS 0.016937f
C799 VTAIL.n304 VSUBS 0.017934f
C800 VTAIL.n305 VSUBS 0.040034f
C801 VTAIL.n306 VSUBS 0.040034f
C802 VTAIL.n307 VSUBS 0.017934f
C803 VTAIL.n308 VSUBS 0.016937f
C804 VTAIL.n309 VSUBS 0.03152f
C805 VTAIL.n310 VSUBS 0.03152f
C806 VTAIL.n311 VSUBS 0.016937f
C807 VTAIL.n312 VSUBS 0.017934f
C808 VTAIL.n313 VSUBS 0.040034f
C809 VTAIL.n314 VSUBS 0.040034f
C810 VTAIL.n315 VSUBS 0.017934f
C811 VTAIL.n316 VSUBS 0.016937f
C812 VTAIL.n317 VSUBS 0.03152f
C813 VTAIL.n318 VSUBS 0.03152f
C814 VTAIL.n319 VSUBS 0.016937f
C815 VTAIL.n320 VSUBS 0.017934f
C816 VTAIL.n321 VSUBS 0.040034f
C817 VTAIL.n322 VSUBS 0.098743f
C818 VTAIL.n323 VSUBS 0.017934f
C819 VTAIL.n324 VSUBS 0.016937f
C820 VTAIL.n325 VSUBS 0.071564f
C821 VTAIL.n326 VSUBS 0.049698f
C822 VTAIL.n327 VSUBS 1.18477f
C823 VDD2.t0 VSUBS 0.201578f
C824 VDD2.t3 VSUBS 0.201578f
C825 VDD2.n0 VSUBS 1.41091f
C826 VDD2.t2 VSUBS 0.201578f
C827 VDD2.t5 VSUBS 0.201578f
C828 VDD2.n1 VSUBS 1.41091f
C829 VDD2.n2 VSUBS 2.81139f
C830 VDD2.t6 VSUBS 0.201578f
C831 VDD2.t7 VSUBS 0.201578f
C832 VDD2.n3 VSUBS 1.40963f
C833 VDD2.n4 VSUBS 2.71196f
C834 VDD2.t4 VSUBS 0.201578f
C835 VDD2.t1 VSUBS 0.201578f
C836 VDD2.n5 VSUBS 1.41087f
C837 VN.n0 VSUBS 0.111037f
C838 VN.t6 VSUBS 0.188949f
C839 VN.t7 VSUBS 0.188949f
C840 VN.t0 VSUBS 0.191439f
C841 VN.n1 VSUBS 0.101857f
C842 VN.n2 VSUBS 0.089371f
C843 VN.n3 VSUBS 0.017511f
C844 VN.n4 VSUBS 0.089371f
C845 VN.t4 VSUBS 0.191439f
C846 VN.n5 VSUBS 0.101789f
C847 VN.n6 VSUBS 0.040908f
C848 VN.n7 VSUBS 0.111037f
C849 VN.t3 VSUBS 0.191439f
C850 VN.t5 VSUBS 0.188949f
C851 VN.t1 VSUBS 0.188949f
C852 VN.t2 VSUBS 0.191439f
C853 VN.n8 VSUBS 0.101857f
C854 VN.n9 VSUBS 0.089371f
C855 VN.n10 VSUBS 0.017511f
C856 VN.n11 VSUBS 0.089371f
C857 VN.n12 VSUBS 0.101789f
C858 VN.n13 VSUBS 1.69989f
.ends

