* NGSPICE file created from diff_pair_sample_0525.ext - technology: sky130A

.subckt diff_pair_sample_0525 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=1.52295 ps=9.56 w=9.23 l=0.73
X1 B.t11 B.t9 B.t10 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=0 ps=0 w=9.23 l=0.73
X2 B.t8 B.t6 B.t7 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=0 ps=0 w=9.23 l=0.73
X3 VDD1.t4 VP.t1 VTAIL.t10 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=3.5997 ps=19.24 w=9.23 l=0.73
X4 VTAIL.t9 VP.t2 VDD1.t3 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=1.52295 ps=9.56 w=9.23 l=0.73
X5 VDD1.t2 VP.t3 VTAIL.t8 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=1.52295 ps=9.56 w=9.23 l=0.73
X6 VDD1.t1 VP.t4 VTAIL.t11 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=3.5997 ps=19.24 w=9.23 l=0.73
X7 VDD2.t5 VN.t0 VTAIL.t1 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=3.5997 ps=19.24 w=9.23 l=0.73
X8 VDD2.t4 VN.t1 VTAIL.t0 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=1.52295 ps=9.56 w=9.23 l=0.73
X9 B.t5 B.t3 B.t4 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=0 ps=0 w=9.23 l=0.73
X10 VTAIL.t7 VP.t5 VDD1.t0 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=1.52295 ps=9.56 w=9.23 l=0.73
X11 B.t2 B.t0 B.t1 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=0 ps=0 w=9.23 l=0.73
X12 VTAIL.t5 VN.t2 VDD2.t3 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=1.52295 ps=9.56 w=9.23 l=0.73
X13 VDD2.t2 VN.t3 VTAIL.t4 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=3.5997 pd=19.24 as=1.52295 ps=9.56 w=9.23 l=0.73
X14 VDD2.t1 VN.t4 VTAIL.t3 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=3.5997 ps=19.24 w=9.23 l=0.73
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n1818_n2814# sky130_fd_pr__pfet_01v8 ad=1.52295 pd=9.56 as=1.52295 ps=9.56 w=9.23 l=0.73
R0 VP.n3 VP.t0 381.038
R1 VP.n8 VP.t3 358.86
R2 VP.n12 VP.t2 358.86
R3 VP.n14 VP.t4 358.86
R4 VP.n6 VP.t1 358.86
R5 VP.n4 VP.t5 358.86
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.862
R14 VP.n9 VP.n7 39.2505
R15 VP.n8 VP.n1 28.4823
R16 VP.n14 VP.n13 28.4823
R17 VP.n6 VP.n5 28.4823
R18 VP.n12 VP.n1 19.7187
R19 VP.n13 VP.n12 19.7187
R20 VP.n5 VP.n4 19.7187
R21 VP.n4 VP.n3 19.7081
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VTAIL.n202 VTAIL.n158 756.745
R29 VTAIL.n46 VTAIL.n2 756.745
R30 VTAIL.n152 VTAIL.n108 756.745
R31 VTAIL.n100 VTAIL.n56 756.745
R32 VTAIL.n175 VTAIL.n174 585
R33 VTAIL.n177 VTAIL.n176 585
R34 VTAIL.n170 VTAIL.n169 585
R35 VTAIL.n183 VTAIL.n182 585
R36 VTAIL.n185 VTAIL.n184 585
R37 VTAIL.n166 VTAIL.n165 585
R38 VTAIL.n192 VTAIL.n191 585
R39 VTAIL.n193 VTAIL.n164 585
R40 VTAIL.n195 VTAIL.n194 585
R41 VTAIL.n162 VTAIL.n161 585
R42 VTAIL.n201 VTAIL.n200 585
R43 VTAIL.n203 VTAIL.n202 585
R44 VTAIL.n19 VTAIL.n18 585
R45 VTAIL.n21 VTAIL.n20 585
R46 VTAIL.n14 VTAIL.n13 585
R47 VTAIL.n27 VTAIL.n26 585
R48 VTAIL.n29 VTAIL.n28 585
R49 VTAIL.n10 VTAIL.n9 585
R50 VTAIL.n36 VTAIL.n35 585
R51 VTAIL.n37 VTAIL.n8 585
R52 VTAIL.n39 VTAIL.n38 585
R53 VTAIL.n6 VTAIL.n5 585
R54 VTAIL.n45 VTAIL.n44 585
R55 VTAIL.n47 VTAIL.n46 585
R56 VTAIL.n153 VTAIL.n152 585
R57 VTAIL.n151 VTAIL.n150 585
R58 VTAIL.n112 VTAIL.n111 585
R59 VTAIL.n116 VTAIL.n114 585
R60 VTAIL.n145 VTAIL.n144 585
R61 VTAIL.n143 VTAIL.n142 585
R62 VTAIL.n118 VTAIL.n117 585
R63 VTAIL.n137 VTAIL.n136 585
R64 VTAIL.n135 VTAIL.n134 585
R65 VTAIL.n122 VTAIL.n121 585
R66 VTAIL.n129 VTAIL.n128 585
R67 VTAIL.n127 VTAIL.n126 585
R68 VTAIL.n101 VTAIL.n100 585
R69 VTAIL.n99 VTAIL.n98 585
R70 VTAIL.n60 VTAIL.n59 585
R71 VTAIL.n64 VTAIL.n62 585
R72 VTAIL.n93 VTAIL.n92 585
R73 VTAIL.n91 VTAIL.n90 585
R74 VTAIL.n66 VTAIL.n65 585
R75 VTAIL.n85 VTAIL.n84 585
R76 VTAIL.n83 VTAIL.n82 585
R77 VTAIL.n70 VTAIL.n69 585
R78 VTAIL.n77 VTAIL.n76 585
R79 VTAIL.n75 VTAIL.n74 585
R80 VTAIL.n173 VTAIL.t3 329.038
R81 VTAIL.n17 VTAIL.t11 329.038
R82 VTAIL.n125 VTAIL.t10 329.038
R83 VTAIL.n73 VTAIL.t1 329.038
R84 VTAIL.n176 VTAIL.n175 171.744
R85 VTAIL.n176 VTAIL.n169 171.744
R86 VTAIL.n183 VTAIL.n169 171.744
R87 VTAIL.n184 VTAIL.n183 171.744
R88 VTAIL.n184 VTAIL.n165 171.744
R89 VTAIL.n192 VTAIL.n165 171.744
R90 VTAIL.n193 VTAIL.n192 171.744
R91 VTAIL.n194 VTAIL.n193 171.744
R92 VTAIL.n194 VTAIL.n161 171.744
R93 VTAIL.n201 VTAIL.n161 171.744
R94 VTAIL.n202 VTAIL.n201 171.744
R95 VTAIL.n20 VTAIL.n19 171.744
R96 VTAIL.n20 VTAIL.n13 171.744
R97 VTAIL.n27 VTAIL.n13 171.744
R98 VTAIL.n28 VTAIL.n27 171.744
R99 VTAIL.n28 VTAIL.n9 171.744
R100 VTAIL.n36 VTAIL.n9 171.744
R101 VTAIL.n37 VTAIL.n36 171.744
R102 VTAIL.n38 VTAIL.n37 171.744
R103 VTAIL.n38 VTAIL.n5 171.744
R104 VTAIL.n45 VTAIL.n5 171.744
R105 VTAIL.n46 VTAIL.n45 171.744
R106 VTAIL.n152 VTAIL.n151 171.744
R107 VTAIL.n151 VTAIL.n111 171.744
R108 VTAIL.n116 VTAIL.n111 171.744
R109 VTAIL.n144 VTAIL.n116 171.744
R110 VTAIL.n144 VTAIL.n143 171.744
R111 VTAIL.n143 VTAIL.n117 171.744
R112 VTAIL.n136 VTAIL.n117 171.744
R113 VTAIL.n136 VTAIL.n135 171.744
R114 VTAIL.n135 VTAIL.n121 171.744
R115 VTAIL.n128 VTAIL.n121 171.744
R116 VTAIL.n128 VTAIL.n127 171.744
R117 VTAIL.n100 VTAIL.n99 171.744
R118 VTAIL.n99 VTAIL.n59 171.744
R119 VTAIL.n64 VTAIL.n59 171.744
R120 VTAIL.n92 VTAIL.n64 171.744
R121 VTAIL.n92 VTAIL.n91 171.744
R122 VTAIL.n91 VTAIL.n65 171.744
R123 VTAIL.n84 VTAIL.n65 171.744
R124 VTAIL.n84 VTAIL.n83 171.744
R125 VTAIL.n83 VTAIL.n69 171.744
R126 VTAIL.n76 VTAIL.n69 171.744
R127 VTAIL.n76 VTAIL.n75 171.744
R128 VTAIL.n175 VTAIL.t3 85.8723
R129 VTAIL.n19 VTAIL.t11 85.8723
R130 VTAIL.n127 VTAIL.t10 85.8723
R131 VTAIL.n75 VTAIL.t1 85.8723
R132 VTAIL.n107 VTAIL.n106 61.7082
R133 VTAIL.n55 VTAIL.n54 61.7082
R134 VTAIL.n1 VTAIL.n0 61.708
R135 VTAIL.n53 VTAIL.n52 61.708
R136 VTAIL.n207 VTAIL.n206 31.9914
R137 VTAIL.n51 VTAIL.n50 31.9914
R138 VTAIL.n157 VTAIL.n156 31.9914
R139 VTAIL.n105 VTAIL.n104 31.9914
R140 VTAIL.n55 VTAIL.n53 22.1514
R141 VTAIL.n207 VTAIL.n157 21.2376
R142 VTAIL.n195 VTAIL.n162 13.1884
R143 VTAIL.n39 VTAIL.n6 13.1884
R144 VTAIL.n114 VTAIL.n112 13.1884
R145 VTAIL.n62 VTAIL.n60 13.1884
R146 VTAIL.n196 VTAIL.n164 12.8005
R147 VTAIL.n200 VTAIL.n199 12.8005
R148 VTAIL.n40 VTAIL.n8 12.8005
R149 VTAIL.n44 VTAIL.n43 12.8005
R150 VTAIL.n150 VTAIL.n149 12.8005
R151 VTAIL.n146 VTAIL.n145 12.8005
R152 VTAIL.n98 VTAIL.n97 12.8005
R153 VTAIL.n94 VTAIL.n93 12.8005
R154 VTAIL.n191 VTAIL.n190 12.0247
R155 VTAIL.n203 VTAIL.n160 12.0247
R156 VTAIL.n35 VTAIL.n34 12.0247
R157 VTAIL.n47 VTAIL.n4 12.0247
R158 VTAIL.n153 VTAIL.n110 12.0247
R159 VTAIL.n142 VTAIL.n115 12.0247
R160 VTAIL.n101 VTAIL.n58 12.0247
R161 VTAIL.n90 VTAIL.n63 12.0247
R162 VTAIL.n189 VTAIL.n166 11.249
R163 VTAIL.n204 VTAIL.n158 11.249
R164 VTAIL.n33 VTAIL.n10 11.249
R165 VTAIL.n48 VTAIL.n2 11.249
R166 VTAIL.n154 VTAIL.n108 11.249
R167 VTAIL.n141 VTAIL.n118 11.249
R168 VTAIL.n102 VTAIL.n56 11.249
R169 VTAIL.n89 VTAIL.n66 11.249
R170 VTAIL.n174 VTAIL.n173 10.7239
R171 VTAIL.n18 VTAIL.n17 10.7239
R172 VTAIL.n126 VTAIL.n125 10.7239
R173 VTAIL.n74 VTAIL.n73 10.7239
R174 VTAIL.n186 VTAIL.n185 10.4732
R175 VTAIL.n30 VTAIL.n29 10.4732
R176 VTAIL.n138 VTAIL.n137 10.4732
R177 VTAIL.n86 VTAIL.n85 10.4732
R178 VTAIL.n182 VTAIL.n168 9.69747
R179 VTAIL.n26 VTAIL.n12 9.69747
R180 VTAIL.n134 VTAIL.n120 9.69747
R181 VTAIL.n82 VTAIL.n68 9.69747
R182 VTAIL.n206 VTAIL.n205 9.45567
R183 VTAIL.n50 VTAIL.n49 9.45567
R184 VTAIL.n156 VTAIL.n155 9.45567
R185 VTAIL.n104 VTAIL.n103 9.45567
R186 VTAIL.n205 VTAIL.n204 9.3005
R187 VTAIL.n160 VTAIL.n159 9.3005
R188 VTAIL.n199 VTAIL.n198 9.3005
R189 VTAIL.n172 VTAIL.n171 9.3005
R190 VTAIL.n179 VTAIL.n178 9.3005
R191 VTAIL.n181 VTAIL.n180 9.3005
R192 VTAIL.n168 VTAIL.n167 9.3005
R193 VTAIL.n187 VTAIL.n186 9.3005
R194 VTAIL.n189 VTAIL.n188 9.3005
R195 VTAIL.n190 VTAIL.n163 9.3005
R196 VTAIL.n197 VTAIL.n196 9.3005
R197 VTAIL.n49 VTAIL.n48 9.3005
R198 VTAIL.n4 VTAIL.n3 9.3005
R199 VTAIL.n43 VTAIL.n42 9.3005
R200 VTAIL.n16 VTAIL.n15 9.3005
R201 VTAIL.n23 VTAIL.n22 9.3005
R202 VTAIL.n25 VTAIL.n24 9.3005
R203 VTAIL.n12 VTAIL.n11 9.3005
R204 VTAIL.n31 VTAIL.n30 9.3005
R205 VTAIL.n33 VTAIL.n32 9.3005
R206 VTAIL.n34 VTAIL.n7 9.3005
R207 VTAIL.n41 VTAIL.n40 9.3005
R208 VTAIL.n124 VTAIL.n123 9.3005
R209 VTAIL.n131 VTAIL.n130 9.3005
R210 VTAIL.n133 VTAIL.n132 9.3005
R211 VTAIL.n120 VTAIL.n119 9.3005
R212 VTAIL.n139 VTAIL.n138 9.3005
R213 VTAIL.n141 VTAIL.n140 9.3005
R214 VTAIL.n115 VTAIL.n113 9.3005
R215 VTAIL.n147 VTAIL.n146 9.3005
R216 VTAIL.n155 VTAIL.n154 9.3005
R217 VTAIL.n110 VTAIL.n109 9.3005
R218 VTAIL.n149 VTAIL.n148 9.3005
R219 VTAIL.n72 VTAIL.n71 9.3005
R220 VTAIL.n79 VTAIL.n78 9.3005
R221 VTAIL.n81 VTAIL.n80 9.3005
R222 VTAIL.n68 VTAIL.n67 9.3005
R223 VTAIL.n87 VTAIL.n86 9.3005
R224 VTAIL.n89 VTAIL.n88 9.3005
R225 VTAIL.n63 VTAIL.n61 9.3005
R226 VTAIL.n95 VTAIL.n94 9.3005
R227 VTAIL.n103 VTAIL.n102 9.3005
R228 VTAIL.n58 VTAIL.n57 9.3005
R229 VTAIL.n97 VTAIL.n96 9.3005
R230 VTAIL.n181 VTAIL.n170 8.92171
R231 VTAIL.n25 VTAIL.n14 8.92171
R232 VTAIL.n133 VTAIL.n122 8.92171
R233 VTAIL.n81 VTAIL.n70 8.92171
R234 VTAIL.n178 VTAIL.n177 8.14595
R235 VTAIL.n22 VTAIL.n21 8.14595
R236 VTAIL.n130 VTAIL.n129 8.14595
R237 VTAIL.n78 VTAIL.n77 8.14595
R238 VTAIL.n174 VTAIL.n172 7.3702
R239 VTAIL.n18 VTAIL.n16 7.3702
R240 VTAIL.n126 VTAIL.n124 7.3702
R241 VTAIL.n74 VTAIL.n72 7.3702
R242 VTAIL.n177 VTAIL.n172 5.81868
R243 VTAIL.n21 VTAIL.n16 5.81868
R244 VTAIL.n129 VTAIL.n124 5.81868
R245 VTAIL.n77 VTAIL.n72 5.81868
R246 VTAIL.n178 VTAIL.n170 5.04292
R247 VTAIL.n22 VTAIL.n14 5.04292
R248 VTAIL.n130 VTAIL.n122 5.04292
R249 VTAIL.n78 VTAIL.n70 5.04292
R250 VTAIL.n182 VTAIL.n181 4.26717
R251 VTAIL.n26 VTAIL.n25 4.26717
R252 VTAIL.n134 VTAIL.n133 4.26717
R253 VTAIL.n82 VTAIL.n81 4.26717
R254 VTAIL.n0 VTAIL.t4 3.52217
R255 VTAIL.n0 VTAIL.t5 3.52217
R256 VTAIL.n52 VTAIL.t8 3.52217
R257 VTAIL.n52 VTAIL.t9 3.52217
R258 VTAIL.n106 VTAIL.t6 3.52217
R259 VTAIL.n106 VTAIL.t7 3.52217
R260 VTAIL.n54 VTAIL.t0 3.52217
R261 VTAIL.n54 VTAIL.t2 3.52217
R262 VTAIL.n185 VTAIL.n168 3.49141
R263 VTAIL.n29 VTAIL.n12 3.49141
R264 VTAIL.n137 VTAIL.n120 3.49141
R265 VTAIL.n85 VTAIL.n68 3.49141
R266 VTAIL.n186 VTAIL.n166 2.71565
R267 VTAIL.n206 VTAIL.n158 2.71565
R268 VTAIL.n30 VTAIL.n10 2.71565
R269 VTAIL.n50 VTAIL.n2 2.71565
R270 VTAIL.n156 VTAIL.n108 2.71565
R271 VTAIL.n138 VTAIL.n118 2.71565
R272 VTAIL.n104 VTAIL.n56 2.71565
R273 VTAIL.n86 VTAIL.n66 2.71565
R274 VTAIL.n173 VTAIL.n171 2.41283
R275 VTAIL.n17 VTAIL.n15 2.41283
R276 VTAIL.n125 VTAIL.n123 2.41283
R277 VTAIL.n73 VTAIL.n71 2.41283
R278 VTAIL.n191 VTAIL.n189 1.93989
R279 VTAIL.n204 VTAIL.n203 1.93989
R280 VTAIL.n35 VTAIL.n33 1.93989
R281 VTAIL.n48 VTAIL.n47 1.93989
R282 VTAIL.n154 VTAIL.n153 1.93989
R283 VTAIL.n142 VTAIL.n141 1.93989
R284 VTAIL.n102 VTAIL.n101 1.93989
R285 VTAIL.n90 VTAIL.n89 1.93989
R286 VTAIL.n190 VTAIL.n164 1.16414
R287 VTAIL.n200 VTAIL.n160 1.16414
R288 VTAIL.n34 VTAIL.n8 1.16414
R289 VTAIL.n44 VTAIL.n4 1.16414
R290 VTAIL.n150 VTAIL.n110 1.16414
R291 VTAIL.n145 VTAIL.n115 1.16414
R292 VTAIL.n98 VTAIL.n58 1.16414
R293 VTAIL.n93 VTAIL.n63 1.16414
R294 VTAIL.n107 VTAIL.n105 0.927224
R295 VTAIL.n51 VTAIL.n1 0.927224
R296 VTAIL.n105 VTAIL.n55 0.914293
R297 VTAIL.n157 VTAIL.n107 0.914293
R298 VTAIL.n53 VTAIL.n51 0.914293
R299 VTAIL VTAIL.n207 0.627655
R300 VTAIL.n196 VTAIL.n195 0.388379
R301 VTAIL.n199 VTAIL.n162 0.388379
R302 VTAIL.n40 VTAIL.n39 0.388379
R303 VTAIL.n43 VTAIL.n6 0.388379
R304 VTAIL.n149 VTAIL.n112 0.388379
R305 VTAIL.n146 VTAIL.n114 0.388379
R306 VTAIL.n97 VTAIL.n60 0.388379
R307 VTAIL.n94 VTAIL.n62 0.388379
R308 VTAIL VTAIL.n1 0.287138
R309 VTAIL.n179 VTAIL.n171 0.155672
R310 VTAIL.n180 VTAIL.n179 0.155672
R311 VTAIL.n180 VTAIL.n167 0.155672
R312 VTAIL.n187 VTAIL.n167 0.155672
R313 VTAIL.n188 VTAIL.n187 0.155672
R314 VTAIL.n188 VTAIL.n163 0.155672
R315 VTAIL.n197 VTAIL.n163 0.155672
R316 VTAIL.n198 VTAIL.n197 0.155672
R317 VTAIL.n198 VTAIL.n159 0.155672
R318 VTAIL.n205 VTAIL.n159 0.155672
R319 VTAIL.n23 VTAIL.n15 0.155672
R320 VTAIL.n24 VTAIL.n23 0.155672
R321 VTAIL.n24 VTAIL.n11 0.155672
R322 VTAIL.n31 VTAIL.n11 0.155672
R323 VTAIL.n32 VTAIL.n31 0.155672
R324 VTAIL.n32 VTAIL.n7 0.155672
R325 VTAIL.n41 VTAIL.n7 0.155672
R326 VTAIL.n42 VTAIL.n41 0.155672
R327 VTAIL.n42 VTAIL.n3 0.155672
R328 VTAIL.n49 VTAIL.n3 0.155672
R329 VTAIL.n155 VTAIL.n109 0.155672
R330 VTAIL.n148 VTAIL.n109 0.155672
R331 VTAIL.n148 VTAIL.n147 0.155672
R332 VTAIL.n147 VTAIL.n113 0.155672
R333 VTAIL.n140 VTAIL.n113 0.155672
R334 VTAIL.n140 VTAIL.n139 0.155672
R335 VTAIL.n139 VTAIL.n119 0.155672
R336 VTAIL.n132 VTAIL.n119 0.155672
R337 VTAIL.n132 VTAIL.n131 0.155672
R338 VTAIL.n131 VTAIL.n123 0.155672
R339 VTAIL.n103 VTAIL.n57 0.155672
R340 VTAIL.n96 VTAIL.n57 0.155672
R341 VTAIL.n96 VTAIL.n95 0.155672
R342 VTAIL.n95 VTAIL.n61 0.155672
R343 VTAIL.n88 VTAIL.n61 0.155672
R344 VTAIL.n88 VTAIL.n87 0.155672
R345 VTAIL.n87 VTAIL.n67 0.155672
R346 VTAIL.n80 VTAIL.n67 0.155672
R347 VTAIL.n80 VTAIL.n79 0.155672
R348 VTAIL.n79 VTAIL.n71 0.155672
R349 VDD1.n44 VDD1.n0 756.745
R350 VDD1.n93 VDD1.n49 756.745
R351 VDD1.n45 VDD1.n44 585
R352 VDD1.n43 VDD1.n42 585
R353 VDD1.n4 VDD1.n3 585
R354 VDD1.n8 VDD1.n6 585
R355 VDD1.n37 VDD1.n36 585
R356 VDD1.n35 VDD1.n34 585
R357 VDD1.n10 VDD1.n9 585
R358 VDD1.n29 VDD1.n28 585
R359 VDD1.n27 VDD1.n26 585
R360 VDD1.n14 VDD1.n13 585
R361 VDD1.n21 VDD1.n20 585
R362 VDD1.n19 VDD1.n18 585
R363 VDD1.n66 VDD1.n65 585
R364 VDD1.n68 VDD1.n67 585
R365 VDD1.n61 VDD1.n60 585
R366 VDD1.n74 VDD1.n73 585
R367 VDD1.n76 VDD1.n75 585
R368 VDD1.n57 VDD1.n56 585
R369 VDD1.n83 VDD1.n82 585
R370 VDD1.n84 VDD1.n55 585
R371 VDD1.n86 VDD1.n85 585
R372 VDD1.n53 VDD1.n52 585
R373 VDD1.n92 VDD1.n91 585
R374 VDD1.n94 VDD1.n93 585
R375 VDD1.n17 VDD1.t5 329.038
R376 VDD1.n64 VDD1.t2 329.038
R377 VDD1.n44 VDD1.n43 171.744
R378 VDD1.n43 VDD1.n3 171.744
R379 VDD1.n8 VDD1.n3 171.744
R380 VDD1.n36 VDD1.n8 171.744
R381 VDD1.n36 VDD1.n35 171.744
R382 VDD1.n35 VDD1.n9 171.744
R383 VDD1.n28 VDD1.n9 171.744
R384 VDD1.n28 VDD1.n27 171.744
R385 VDD1.n27 VDD1.n13 171.744
R386 VDD1.n20 VDD1.n13 171.744
R387 VDD1.n20 VDD1.n19 171.744
R388 VDD1.n67 VDD1.n66 171.744
R389 VDD1.n67 VDD1.n60 171.744
R390 VDD1.n74 VDD1.n60 171.744
R391 VDD1.n75 VDD1.n74 171.744
R392 VDD1.n75 VDD1.n56 171.744
R393 VDD1.n83 VDD1.n56 171.744
R394 VDD1.n84 VDD1.n83 171.744
R395 VDD1.n85 VDD1.n84 171.744
R396 VDD1.n85 VDD1.n52 171.744
R397 VDD1.n92 VDD1.n52 171.744
R398 VDD1.n93 VDD1.n92 171.744
R399 VDD1.n19 VDD1.t5 85.8723
R400 VDD1.n66 VDD1.t2 85.8723
R401 VDD1.n99 VDD1.n98 78.5599
R402 VDD1.n101 VDD1.n100 78.3868
R403 VDD1 VDD1.n48 49.4137
R404 VDD1.n99 VDD1.n97 49.3002
R405 VDD1.n101 VDD1.n99 35.6819
R406 VDD1.n6 VDD1.n4 13.1884
R407 VDD1.n86 VDD1.n53 13.1884
R408 VDD1.n42 VDD1.n41 12.8005
R409 VDD1.n38 VDD1.n37 12.8005
R410 VDD1.n87 VDD1.n55 12.8005
R411 VDD1.n91 VDD1.n90 12.8005
R412 VDD1.n45 VDD1.n2 12.0247
R413 VDD1.n34 VDD1.n7 12.0247
R414 VDD1.n82 VDD1.n81 12.0247
R415 VDD1.n94 VDD1.n51 12.0247
R416 VDD1.n46 VDD1.n0 11.249
R417 VDD1.n33 VDD1.n10 11.249
R418 VDD1.n80 VDD1.n57 11.249
R419 VDD1.n95 VDD1.n49 11.249
R420 VDD1.n18 VDD1.n17 10.7239
R421 VDD1.n65 VDD1.n64 10.7239
R422 VDD1.n30 VDD1.n29 10.4732
R423 VDD1.n77 VDD1.n76 10.4732
R424 VDD1.n26 VDD1.n12 9.69747
R425 VDD1.n73 VDD1.n59 9.69747
R426 VDD1.n48 VDD1.n47 9.45567
R427 VDD1.n97 VDD1.n96 9.45567
R428 VDD1.n16 VDD1.n15 9.3005
R429 VDD1.n23 VDD1.n22 9.3005
R430 VDD1.n25 VDD1.n24 9.3005
R431 VDD1.n12 VDD1.n11 9.3005
R432 VDD1.n31 VDD1.n30 9.3005
R433 VDD1.n33 VDD1.n32 9.3005
R434 VDD1.n7 VDD1.n5 9.3005
R435 VDD1.n39 VDD1.n38 9.3005
R436 VDD1.n47 VDD1.n46 9.3005
R437 VDD1.n2 VDD1.n1 9.3005
R438 VDD1.n41 VDD1.n40 9.3005
R439 VDD1.n96 VDD1.n95 9.3005
R440 VDD1.n51 VDD1.n50 9.3005
R441 VDD1.n90 VDD1.n89 9.3005
R442 VDD1.n63 VDD1.n62 9.3005
R443 VDD1.n70 VDD1.n69 9.3005
R444 VDD1.n72 VDD1.n71 9.3005
R445 VDD1.n59 VDD1.n58 9.3005
R446 VDD1.n78 VDD1.n77 9.3005
R447 VDD1.n80 VDD1.n79 9.3005
R448 VDD1.n81 VDD1.n54 9.3005
R449 VDD1.n88 VDD1.n87 9.3005
R450 VDD1.n25 VDD1.n14 8.92171
R451 VDD1.n72 VDD1.n61 8.92171
R452 VDD1.n22 VDD1.n21 8.14595
R453 VDD1.n69 VDD1.n68 8.14595
R454 VDD1.n18 VDD1.n16 7.3702
R455 VDD1.n65 VDD1.n63 7.3702
R456 VDD1.n21 VDD1.n16 5.81868
R457 VDD1.n68 VDD1.n63 5.81868
R458 VDD1.n22 VDD1.n14 5.04292
R459 VDD1.n69 VDD1.n61 5.04292
R460 VDD1.n26 VDD1.n25 4.26717
R461 VDD1.n73 VDD1.n72 4.26717
R462 VDD1.n100 VDD1.t0 3.52217
R463 VDD1.n100 VDD1.t4 3.52217
R464 VDD1.n98 VDD1.t3 3.52217
R465 VDD1.n98 VDD1.t1 3.52217
R466 VDD1.n29 VDD1.n12 3.49141
R467 VDD1.n76 VDD1.n59 3.49141
R468 VDD1.n48 VDD1.n0 2.71565
R469 VDD1.n30 VDD1.n10 2.71565
R470 VDD1.n77 VDD1.n57 2.71565
R471 VDD1.n97 VDD1.n49 2.71565
R472 VDD1.n17 VDD1.n15 2.41283
R473 VDD1.n64 VDD1.n62 2.41283
R474 VDD1.n46 VDD1.n45 1.93989
R475 VDD1.n34 VDD1.n33 1.93989
R476 VDD1.n82 VDD1.n80 1.93989
R477 VDD1.n95 VDD1.n94 1.93989
R478 VDD1.n42 VDD1.n2 1.16414
R479 VDD1.n37 VDD1.n7 1.16414
R480 VDD1.n81 VDD1.n55 1.16414
R481 VDD1.n91 VDD1.n51 1.16414
R482 VDD1.n41 VDD1.n4 0.388379
R483 VDD1.n38 VDD1.n6 0.388379
R484 VDD1.n87 VDD1.n86 0.388379
R485 VDD1.n90 VDD1.n53 0.388379
R486 VDD1 VDD1.n101 0.170759
R487 VDD1.n47 VDD1.n1 0.155672
R488 VDD1.n40 VDD1.n1 0.155672
R489 VDD1.n40 VDD1.n39 0.155672
R490 VDD1.n39 VDD1.n5 0.155672
R491 VDD1.n32 VDD1.n5 0.155672
R492 VDD1.n32 VDD1.n31 0.155672
R493 VDD1.n31 VDD1.n11 0.155672
R494 VDD1.n24 VDD1.n11 0.155672
R495 VDD1.n24 VDD1.n23 0.155672
R496 VDD1.n23 VDD1.n15 0.155672
R497 VDD1.n70 VDD1.n62 0.155672
R498 VDD1.n71 VDD1.n70 0.155672
R499 VDD1.n71 VDD1.n58 0.155672
R500 VDD1.n78 VDD1.n58 0.155672
R501 VDD1.n79 VDD1.n78 0.155672
R502 VDD1.n79 VDD1.n54 0.155672
R503 VDD1.n88 VDD1.n54 0.155672
R504 VDD1.n89 VDD1.n88 0.155672
R505 VDD1.n89 VDD1.n50 0.155672
R506 VDD1.n96 VDD1.n50 0.155672
R507 B.n273 B.n272 585
R508 B.n271 B.n76 585
R509 B.n270 B.n269 585
R510 B.n268 B.n77 585
R511 B.n267 B.n266 585
R512 B.n265 B.n78 585
R513 B.n264 B.n263 585
R514 B.n262 B.n79 585
R515 B.n261 B.n260 585
R516 B.n259 B.n80 585
R517 B.n258 B.n257 585
R518 B.n256 B.n81 585
R519 B.n255 B.n254 585
R520 B.n253 B.n82 585
R521 B.n252 B.n251 585
R522 B.n250 B.n83 585
R523 B.n249 B.n248 585
R524 B.n247 B.n84 585
R525 B.n246 B.n245 585
R526 B.n244 B.n85 585
R527 B.n243 B.n242 585
R528 B.n241 B.n86 585
R529 B.n240 B.n239 585
R530 B.n238 B.n87 585
R531 B.n237 B.n236 585
R532 B.n235 B.n88 585
R533 B.n234 B.n233 585
R534 B.n232 B.n89 585
R535 B.n231 B.n230 585
R536 B.n229 B.n90 585
R537 B.n228 B.n227 585
R538 B.n226 B.n91 585
R539 B.n225 B.n224 585
R540 B.n223 B.n92 585
R541 B.n222 B.n221 585
R542 B.n217 B.n93 585
R543 B.n216 B.n215 585
R544 B.n214 B.n94 585
R545 B.n213 B.n212 585
R546 B.n211 B.n95 585
R547 B.n210 B.n209 585
R548 B.n208 B.n96 585
R549 B.n207 B.n206 585
R550 B.n204 B.n97 585
R551 B.n203 B.n202 585
R552 B.n201 B.n100 585
R553 B.n200 B.n199 585
R554 B.n198 B.n101 585
R555 B.n197 B.n196 585
R556 B.n195 B.n102 585
R557 B.n194 B.n193 585
R558 B.n192 B.n103 585
R559 B.n191 B.n190 585
R560 B.n189 B.n104 585
R561 B.n188 B.n187 585
R562 B.n186 B.n105 585
R563 B.n185 B.n184 585
R564 B.n183 B.n106 585
R565 B.n182 B.n181 585
R566 B.n180 B.n107 585
R567 B.n179 B.n178 585
R568 B.n177 B.n108 585
R569 B.n176 B.n175 585
R570 B.n174 B.n109 585
R571 B.n173 B.n172 585
R572 B.n171 B.n110 585
R573 B.n170 B.n169 585
R574 B.n168 B.n111 585
R575 B.n167 B.n166 585
R576 B.n165 B.n112 585
R577 B.n164 B.n163 585
R578 B.n162 B.n113 585
R579 B.n161 B.n160 585
R580 B.n159 B.n114 585
R581 B.n158 B.n157 585
R582 B.n156 B.n115 585
R583 B.n155 B.n154 585
R584 B.n274 B.n75 585
R585 B.n276 B.n275 585
R586 B.n277 B.n74 585
R587 B.n279 B.n278 585
R588 B.n280 B.n73 585
R589 B.n282 B.n281 585
R590 B.n283 B.n72 585
R591 B.n285 B.n284 585
R592 B.n286 B.n71 585
R593 B.n288 B.n287 585
R594 B.n289 B.n70 585
R595 B.n291 B.n290 585
R596 B.n292 B.n69 585
R597 B.n294 B.n293 585
R598 B.n295 B.n68 585
R599 B.n297 B.n296 585
R600 B.n298 B.n67 585
R601 B.n300 B.n299 585
R602 B.n301 B.n66 585
R603 B.n303 B.n302 585
R604 B.n304 B.n65 585
R605 B.n306 B.n305 585
R606 B.n307 B.n64 585
R607 B.n309 B.n308 585
R608 B.n310 B.n63 585
R609 B.n312 B.n311 585
R610 B.n313 B.n62 585
R611 B.n315 B.n314 585
R612 B.n316 B.n61 585
R613 B.n318 B.n317 585
R614 B.n319 B.n60 585
R615 B.n321 B.n320 585
R616 B.n322 B.n59 585
R617 B.n324 B.n323 585
R618 B.n325 B.n58 585
R619 B.n327 B.n326 585
R620 B.n328 B.n57 585
R621 B.n330 B.n329 585
R622 B.n331 B.n56 585
R623 B.n333 B.n332 585
R624 B.n334 B.n55 585
R625 B.n336 B.n335 585
R626 B.n453 B.n12 585
R627 B.n452 B.n451 585
R628 B.n450 B.n13 585
R629 B.n449 B.n448 585
R630 B.n447 B.n14 585
R631 B.n446 B.n445 585
R632 B.n444 B.n15 585
R633 B.n443 B.n442 585
R634 B.n441 B.n16 585
R635 B.n440 B.n439 585
R636 B.n438 B.n17 585
R637 B.n437 B.n436 585
R638 B.n435 B.n18 585
R639 B.n434 B.n433 585
R640 B.n432 B.n19 585
R641 B.n431 B.n430 585
R642 B.n429 B.n20 585
R643 B.n428 B.n427 585
R644 B.n426 B.n21 585
R645 B.n425 B.n424 585
R646 B.n423 B.n22 585
R647 B.n422 B.n421 585
R648 B.n420 B.n23 585
R649 B.n419 B.n418 585
R650 B.n417 B.n24 585
R651 B.n416 B.n415 585
R652 B.n414 B.n25 585
R653 B.n413 B.n412 585
R654 B.n411 B.n26 585
R655 B.n410 B.n409 585
R656 B.n408 B.n27 585
R657 B.n407 B.n406 585
R658 B.n405 B.n28 585
R659 B.n404 B.n403 585
R660 B.n401 B.n29 585
R661 B.n400 B.n399 585
R662 B.n398 B.n32 585
R663 B.n397 B.n396 585
R664 B.n395 B.n33 585
R665 B.n394 B.n393 585
R666 B.n392 B.n34 585
R667 B.n391 B.n390 585
R668 B.n389 B.n35 585
R669 B.n387 B.n386 585
R670 B.n385 B.n38 585
R671 B.n384 B.n383 585
R672 B.n382 B.n39 585
R673 B.n381 B.n380 585
R674 B.n379 B.n40 585
R675 B.n378 B.n377 585
R676 B.n376 B.n41 585
R677 B.n375 B.n374 585
R678 B.n373 B.n42 585
R679 B.n372 B.n371 585
R680 B.n370 B.n43 585
R681 B.n369 B.n368 585
R682 B.n367 B.n44 585
R683 B.n366 B.n365 585
R684 B.n364 B.n45 585
R685 B.n363 B.n362 585
R686 B.n361 B.n46 585
R687 B.n360 B.n359 585
R688 B.n358 B.n47 585
R689 B.n357 B.n356 585
R690 B.n355 B.n48 585
R691 B.n354 B.n353 585
R692 B.n352 B.n49 585
R693 B.n351 B.n350 585
R694 B.n349 B.n50 585
R695 B.n348 B.n347 585
R696 B.n346 B.n51 585
R697 B.n345 B.n344 585
R698 B.n343 B.n52 585
R699 B.n342 B.n341 585
R700 B.n340 B.n53 585
R701 B.n339 B.n338 585
R702 B.n337 B.n54 585
R703 B.n455 B.n454 585
R704 B.n456 B.n11 585
R705 B.n458 B.n457 585
R706 B.n459 B.n10 585
R707 B.n461 B.n460 585
R708 B.n462 B.n9 585
R709 B.n464 B.n463 585
R710 B.n465 B.n8 585
R711 B.n467 B.n466 585
R712 B.n468 B.n7 585
R713 B.n470 B.n469 585
R714 B.n471 B.n6 585
R715 B.n473 B.n472 585
R716 B.n474 B.n5 585
R717 B.n476 B.n475 585
R718 B.n477 B.n4 585
R719 B.n479 B.n478 585
R720 B.n480 B.n3 585
R721 B.n482 B.n481 585
R722 B.n483 B.n0 585
R723 B.n2 B.n1 585
R724 B.n126 B.n125 585
R725 B.n128 B.n127 585
R726 B.n129 B.n124 585
R727 B.n131 B.n130 585
R728 B.n132 B.n123 585
R729 B.n134 B.n133 585
R730 B.n135 B.n122 585
R731 B.n137 B.n136 585
R732 B.n138 B.n121 585
R733 B.n140 B.n139 585
R734 B.n141 B.n120 585
R735 B.n143 B.n142 585
R736 B.n144 B.n119 585
R737 B.n146 B.n145 585
R738 B.n147 B.n118 585
R739 B.n149 B.n148 585
R740 B.n150 B.n117 585
R741 B.n152 B.n151 585
R742 B.n153 B.n116 585
R743 B.n98 B.t9 507.327
R744 B.n218 B.t0 507.327
R745 B.n36 B.t6 507.327
R746 B.n30 B.t3 507.327
R747 B.n154 B.n153 473.281
R748 B.n272 B.n75 473.281
R749 B.n337 B.n336 473.281
R750 B.n454 B.n453 473.281
R751 B.n218 B.t1 346.154
R752 B.n36 B.t8 346.154
R753 B.n98 B.t10 346.154
R754 B.n30 B.t5 346.154
R755 B.n219 B.t2 325.596
R756 B.n37 B.t7 325.596
R757 B.n99 B.t11 325.596
R758 B.n31 B.t4 325.596
R759 B.n485 B.n484 256.663
R760 B.n484 B.n483 235.042
R761 B.n484 B.n2 235.042
R762 B.n154 B.n115 163.367
R763 B.n158 B.n115 163.367
R764 B.n159 B.n158 163.367
R765 B.n160 B.n159 163.367
R766 B.n160 B.n113 163.367
R767 B.n164 B.n113 163.367
R768 B.n165 B.n164 163.367
R769 B.n166 B.n165 163.367
R770 B.n166 B.n111 163.367
R771 B.n170 B.n111 163.367
R772 B.n171 B.n170 163.367
R773 B.n172 B.n171 163.367
R774 B.n172 B.n109 163.367
R775 B.n176 B.n109 163.367
R776 B.n177 B.n176 163.367
R777 B.n178 B.n177 163.367
R778 B.n178 B.n107 163.367
R779 B.n182 B.n107 163.367
R780 B.n183 B.n182 163.367
R781 B.n184 B.n183 163.367
R782 B.n184 B.n105 163.367
R783 B.n188 B.n105 163.367
R784 B.n189 B.n188 163.367
R785 B.n190 B.n189 163.367
R786 B.n190 B.n103 163.367
R787 B.n194 B.n103 163.367
R788 B.n195 B.n194 163.367
R789 B.n196 B.n195 163.367
R790 B.n196 B.n101 163.367
R791 B.n200 B.n101 163.367
R792 B.n201 B.n200 163.367
R793 B.n202 B.n201 163.367
R794 B.n202 B.n97 163.367
R795 B.n207 B.n97 163.367
R796 B.n208 B.n207 163.367
R797 B.n209 B.n208 163.367
R798 B.n209 B.n95 163.367
R799 B.n213 B.n95 163.367
R800 B.n214 B.n213 163.367
R801 B.n215 B.n214 163.367
R802 B.n215 B.n93 163.367
R803 B.n222 B.n93 163.367
R804 B.n223 B.n222 163.367
R805 B.n224 B.n223 163.367
R806 B.n224 B.n91 163.367
R807 B.n228 B.n91 163.367
R808 B.n229 B.n228 163.367
R809 B.n230 B.n229 163.367
R810 B.n230 B.n89 163.367
R811 B.n234 B.n89 163.367
R812 B.n235 B.n234 163.367
R813 B.n236 B.n235 163.367
R814 B.n236 B.n87 163.367
R815 B.n240 B.n87 163.367
R816 B.n241 B.n240 163.367
R817 B.n242 B.n241 163.367
R818 B.n242 B.n85 163.367
R819 B.n246 B.n85 163.367
R820 B.n247 B.n246 163.367
R821 B.n248 B.n247 163.367
R822 B.n248 B.n83 163.367
R823 B.n252 B.n83 163.367
R824 B.n253 B.n252 163.367
R825 B.n254 B.n253 163.367
R826 B.n254 B.n81 163.367
R827 B.n258 B.n81 163.367
R828 B.n259 B.n258 163.367
R829 B.n260 B.n259 163.367
R830 B.n260 B.n79 163.367
R831 B.n264 B.n79 163.367
R832 B.n265 B.n264 163.367
R833 B.n266 B.n265 163.367
R834 B.n266 B.n77 163.367
R835 B.n270 B.n77 163.367
R836 B.n271 B.n270 163.367
R837 B.n272 B.n271 163.367
R838 B.n336 B.n55 163.367
R839 B.n332 B.n55 163.367
R840 B.n332 B.n331 163.367
R841 B.n331 B.n330 163.367
R842 B.n330 B.n57 163.367
R843 B.n326 B.n57 163.367
R844 B.n326 B.n325 163.367
R845 B.n325 B.n324 163.367
R846 B.n324 B.n59 163.367
R847 B.n320 B.n59 163.367
R848 B.n320 B.n319 163.367
R849 B.n319 B.n318 163.367
R850 B.n318 B.n61 163.367
R851 B.n314 B.n61 163.367
R852 B.n314 B.n313 163.367
R853 B.n313 B.n312 163.367
R854 B.n312 B.n63 163.367
R855 B.n308 B.n63 163.367
R856 B.n308 B.n307 163.367
R857 B.n307 B.n306 163.367
R858 B.n306 B.n65 163.367
R859 B.n302 B.n65 163.367
R860 B.n302 B.n301 163.367
R861 B.n301 B.n300 163.367
R862 B.n300 B.n67 163.367
R863 B.n296 B.n67 163.367
R864 B.n296 B.n295 163.367
R865 B.n295 B.n294 163.367
R866 B.n294 B.n69 163.367
R867 B.n290 B.n69 163.367
R868 B.n290 B.n289 163.367
R869 B.n289 B.n288 163.367
R870 B.n288 B.n71 163.367
R871 B.n284 B.n71 163.367
R872 B.n284 B.n283 163.367
R873 B.n283 B.n282 163.367
R874 B.n282 B.n73 163.367
R875 B.n278 B.n73 163.367
R876 B.n278 B.n277 163.367
R877 B.n277 B.n276 163.367
R878 B.n276 B.n75 163.367
R879 B.n453 B.n452 163.367
R880 B.n452 B.n13 163.367
R881 B.n448 B.n13 163.367
R882 B.n448 B.n447 163.367
R883 B.n447 B.n446 163.367
R884 B.n446 B.n15 163.367
R885 B.n442 B.n15 163.367
R886 B.n442 B.n441 163.367
R887 B.n441 B.n440 163.367
R888 B.n440 B.n17 163.367
R889 B.n436 B.n17 163.367
R890 B.n436 B.n435 163.367
R891 B.n435 B.n434 163.367
R892 B.n434 B.n19 163.367
R893 B.n430 B.n19 163.367
R894 B.n430 B.n429 163.367
R895 B.n429 B.n428 163.367
R896 B.n428 B.n21 163.367
R897 B.n424 B.n21 163.367
R898 B.n424 B.n423 163.367
R899 B.n423 B.n422 163.367
R900 B.n422 B.n23 163.367
R901 B.n418 B.n23 163.367
R902 B.n418 B.n417 163.367
R903 B.n417 B.n416 163.367
R904 B.n416 B.n25 163.367
R905 B.n412 B.n25 163.367
R906 B.n412 B.n411 163.367
R907 B.n411 B.n410 163.367
R908 B.n410 B.n27 163.367
R909 B.n406 B.n27 163.367
R910 B.n406 B.n405 163.367
R911 B.n405 B.n404 163.367
R912 B.n404 B.n29 163.367
R913 B.n399 B.n29 163.367
R914 B.n399 B.n398 163.367
R915 B.n398 B.n397 163.367
R916 B.n397 B.n33 163.367
R917 B.n393 B.n33 163.367
R918 B.n393 B.n392 163.367
R919 B.n392 B.n391 163.367
R920 B.n391 B.n35 163.367
R921 B.n386 B.n35 163.367
R922 B.n386 B.n385 163.367
R923 B.n385 B.n384 163.367
R924 B.n384 B.n39 163.367
R925 B.n380 B.n39 163.367
R926 B.n380 B.n379 163.367
R927 B.n379 B.n378 163.367
R928 B.n378 B.n41 163.367
R929 B.n374 B.n41 163.367
R930 B.n374 B.n373 163.367
R931 B.n373 B.n372 163.367
R932 B.n372 B.n43 163.367
R933 B.n368 B.n43 163.367
R934 B.n368 B.n367 163.367
R935 B.n367 B.n366 163.367
R936 B.n366 B.n45 163.367
R937 B.n362 B.n45 163.367
R938 B.n362 B.n361 163.367
R939 B.n361 B.n360 163.367
R940 B.n360 B.n47 163.367
R941 B.n356 B.n47 163.367
R942 B.n356 B.n355 163.367
R943 B.n355 B.n354 163.367
R944 B.n354 B.n49 163.367
R945 B.n350 B.n49 163.367
R946 B.n350 B.n349 163.367
R947 B.n349 B.n348 163.367
R948 B.n348 B.n51 163.367
R949 B.n344 B.n51 163.367
R950 B.n344 B.n343 163.367
R951 B.n343 B.n342 163.367
R952 B.n342 B.n53 163.367
R953 B.n338 B.n53 163.367
R954 B.n338 B.n337 163.367
R955 B.n454 B.n11 163.367
R956 B.n458 B.n11 163.367
R957 B.n459 B.n458 163.367
R958 B.n460 B.n459 163.367
R959 B.n460 B.n9 163.367
R960 B.n464 B.n9 163.367
R961 B.n465 B.n464 163.367
R962 B.n466 B.n465 163.367
R963 B.n466 B.n7 163.367
R964 B.n470 B.n7 163.367
R965 B.n471 B.n470 163.367
R966 B.n472 B.n471 163.367
R967 B.n472 B.n5 163.367
R968 B.n476 B.n5 163.367
R969 B.n477 B.n476 163.367
R970 B.n478 B.n477 163.367
R971 B.n478 B.n3 163.367
R972 B.n482 B.n3 163.367
R973 B.n483 B.n482 163.367
R974 B.n125 B.n2 163.367
R975 B.n128 B.n125 163.367
R976 B.n129 B.n128 163.367
R977 B.n130 B.n129 163.367
R978 B.n130 B.n123 163.367
R979 B.n134 B.n123 163.367
R980 B.n135 B.n134 163.367
R981 B.n136 B.n135 163.367
R982 B.n136 B.n121 163.367
R983 B.n140 B.n121 163.367
R984 B.n141 B.n140 163.367
R985 B.n142 B.n141 163.367
R986 B.n142 B.n119 163.367
R987 B.n146 B.n119 163.367
R988 B.n147 B.n146 163.367
R989 B.n148 B.n147 163.367
R990 B.n148 B.n117 163.367
R991 B.n152 B.n117 163.367
R992 B.n153 B.n152 163.367
R993 B.n205 B.n99 59.5399
R994 B.n220 B.n219 59.5399
R995 B.n388 B.n37 59.5399
R996 B.n402 B.n31 59.5399
R997 B.n455 B.n12 30.7517
R998 B.n335 B.n54 30.7517
R999 B.n274 B.n273 30.7517
R1000 B.n155 B.n116 30.7517
R1001 B.n99 B.n98 20.5581
R1002 B.n219 B.n218 20.5581
R1003 B.n37 B.n36 20.5581
R1004 B.n31 B.n30 20.5581
R1005 B B.n485 18.0485
R1006 B.n456 B.n455 10.6151
R1007 B.n457 B.n456 10.6151
R1008 B.n457 B.n10 10.6151
R1009 B.n461 B.n10 10.6151
R1010 B.n462 B.n461 10.6151
R1011 B.n463 B.n462 10.6151
R1012 B.n463 B.n8 10.6151
R1013 B.n467 B.n8 10.6151
R1014 B.n468 B.n467 10.6151
R1015 B.n469 B.n468 10.6151
R1016 B.n469 B.n6 10.6151
R1017 B.n473 B.n6 10.6151
R1018 B.n474 B.n473 10.6151
R1019 B.n475 B.n474 10.6151
R1020 B.n475 B.n4 10.6151
R1021 B.n479 B.n4 10.6151
R1022 B.n480 B.n479 10.6151
R1023 B.n481 B.n480 10.6151
R1024 B.n481 B.n0 10.6151
R1025 B.n451 B.n12 10.6151
R1026 B.n451 B.n450 10.6151
R1027 B.n450 B.n449 10.6151
R1028 B.n449 B.n14 10.6151
R1029 B.n445 B.n14 10.6151
R1030 B.n445 B.n444 10.6151
R1031 B.n444 B.n443 10.6151
R1032 B.n443 B.n16 10.6151
R1033 B.n439 B.n16 10.6151
R1034 B.n439 B.n438 10.6151
R1035 B.n438 B.n437 10.6151
R1036 B.n437 B.n18 10.6151
R1037 B.n433 B.n18 10.6151
R1038 B.n433 B.n432 10.6151
R1039 B.n432 B.n431 10.6151
R1040 B.n431 B.n20 10.6151
R1041 B.n427 B.n20 10.6151
R1042 B.n427 B.n426 10.6151
R1043 B.n426 B.n425 10.6151
R1044 B.n425 B.n22 10.6151
R1045 B.n421 B.n22 10.6151
R1046 B.n421 B.n420 10.6151
R1047 B.n420 B.n419 10.6151
R1048 B.n419 B.n24 10.6151
R1049 B.n415 B.n24 10.6151
R1050 B.n415 B.n414 10.6151
R1051 B.n414 B.n413 10.6151
R1052 B.n413 B.n26 10.6151
R1053 B.n409 B.n26 10.6151
R1054 B.n409 B.n408 10.6151
R1055 B.n408 B.n407 10.6151
R1056 B.n407 B.n28 10.6151
R1057 B.n403 B.n28 10.6151
R1058 B.n401 B.n400 10.6151
R1059 B.n400 B.n32 10.6151
R1060 B.n396 B.n32 10.6151
R1061 B.n396 B.n395 10.6151
R1062 B.n395 B.n394 10.6151
R1063 B.n394 B.n34 10.6151
R1064 B.n390 B.n34 10.6151
R1065 B.n390 B.n389 10.6151
R1066 B.n387 B.n38 10.6151
R1067 B.n383 B.n38 10.6151
R1068 B.n383 B.n382 10.6151
R1069 B.n382 B.n381 10.6151
R1070 B.n381 B.n40 10.6151
R1071 B.n377 B.n40 10.6151
R1072 B.n377 B.n376 10.6151
R1073 B.n376 B.n375 10.6151
R1074 B.n375 B.n42 10.6151
R1075 B.n371 B.n42 10.6151
R1076 B.n371 B.n370 10.6151
R1077 B.n370 B.n369 10.6151
R1078 B.n369 B.n44 10.6151
R1079 B.n365 B.n44 10.6151
R1080 B.n365 B.n364 10.6151
R1081 B.n364 B.n363 10.6151
R1082 B.n363 B.n46 10.6151
R1083 B.n359 B.n46 10.6151
R1084 B.n359 B.n358 10.6151
R1085 B.n358 B.n357 10.6151
R1086 B.n357 B.n48 10.6151
R1087 B.n353 B.n48 10.6151
R1088 B.n353 B.n352 10.6151
R1089 B.n352 B.n351 10.6151
R1090 B.n351 B.n50 10.6151
R1091 B.n347 B.n50 10.6151
R1092 B.n347 B.n346 10.6151
R1093 B.n346 B.n345 10.6151
R1094 B.n345 B.n52 10.6151
R1095 B.n341 B.n52 10.6151
R1096 B.n341 B.n340 10.6151
R1097 B.n340 B.n339 10.6151
R1098 B.n339 B.n54 10.6151
R1099 B.n335 B.n334 10.6151
R1100 B.n334 B.n333 10.6151
R1101 B.n333 B.n56 10.6151
R1102 B.n329 B.n56 10.6151
R1103 B.n329 B.n328 10.6151
R1104 B.n328 B.n327 10.6151
R1105 B.n327 B.n58 10.6151
R1106 B.n323 B.n58 10.6151
R1107 B.n323 B.n322 10.6151
R1108 B.n322 B.n321 10.6151
R1109 B.n321 B.n60 10.6151
R1110 B.n317 B.n60 10.6151
R1111 B.n317 B.n316 10.6151
R1112 B.n316 B.n315 10.6151
R1113 B.n315 B.n62 10.6151
R1114 B.n311 B.n62 10.6151
R1115 B.n311 B.n310 10.6151
R1116 B.n310 B.n309 10.6151
R1117 B.n309 B.n64 10.6151
R1118 B.n305 B.n64 10.6151
R1119 B.n305 B.n304 10.6151
R1120 B.n304 B.n303 10.6151
R1121 B.n303 B.n66 10.6151
R1122 B.n299 B.n66 10.6151
R1123 B.n299 B.n298 10.6151
R1124 B.n298 B.n297 10.6151
R1125 B.n297 B.n68 10.6151
R1126 B.n293 B.n68 10.6151
R1127 B.n293 B.n292 10.6151
R1128 B.n292 B.n291 10.6151
R1129 B.n291 B.n70 10.6151
R1130 B.n287 B.n70 10.6151
R1131 B.n287 B.n286 10.6151
R1132 B.n286 B.n285 10.6151
R1133 B.n285 B.n72 10.6151
R1134 B.n281 B.n72 10.6151
R1135 B.n281 B.n280 10.6151
R1136 B.n280 B.n279 10.6151
R1137 B.n279 B.n74 10.6151
R1138 B.n275 B.n74 10.6151
R1139 B.n275 B.n274 10.6151
R1140 B.n126 B.n1 10.6151
R1141 B.n127 B.n126 10.6151
R1142 B.n127 B.n124 10.6151
R1143 B.n131 B.n124 10.6151
R1144 B.n132 B.n131 10.6151
R1145 B.n133 B.n132 10.6151
R1146 B.n133 B.n122 10.6151
R1147 B.n137 B.n122 10.6151
R1148 B.n138 B.n137 10.6151
R1149 B.n139 B.n138 10.6151
R1150 B.n139 B.n120 10.6151
R1151 B.n143 B.n120 10.6151
R1152 B.n144 B.n143 10.6151
R1153 B.n145 B.n144 10.6151
R1154 B.n145 B.n118 10.6151
R1155 B.n149 B.n118 10.6151
R1156 B.n150 B.n149 10.6151
R1157 B.n151 B.n150 10.6151
R1158 B.n151 B.n116 10.6151
R1159 B.n156 B.n155 10.6151
R1160 B.n157 B.n156 10.6151
R1161 B.n157 B.n114 10.6151
R1162 B.n161 B.n114 10.6151
R1163 B.n162 B.n161 10.6151
R1164 B.n163 B.n162 10.6151
R1165 B.n163 B.n112 10.6151
R1166 B.n167 B.n112 10.6151
R1167 B.n168 B.n167 10.6151
R1168 B.n169 B.n168 10.6151
R1169 B.n169 B.n110 10.6151
R1170 B.n173 B.n110 10.6151
R1171 B.n174 B.n173 10.6151
R1172 B.n175 B.n174 10.6151
R1173 B.n175 B.n108 10.6151
R1174 B.n179 B.n108 10.6151
R1175 B.n180 B.n179 10.6151
R1176 B.n181 B.n180 10.6151
R1177 B.n181 B.n106 10.6151
R1178 B.n185 B.n106 10.6151
R1179 B.n186 B.n185 10.6151
R1180 B.n187 B.n186 10.6151
R1181 B.n187 B.n104 10.6151
R1182 B.n191 B.n104 10.6151
R1183 B.n192 B.n191 10.6151
R1184 B.n193 B.n192 10.6151
R1185 B.n193 B.n102 10.6151
R1186 B.n197 B.n102 10.6151
R1187 B.n198 B.n197 10.6151
R1188 B.n199 B.n198 10.6151
R1189 B.n199 B.n100 10.6151
R1190 B.n203 B.n100 10.6151
R1191 B.n204 B.n203 10.6151
R1192 B.n206 B.n96 10.6151
R1193 B.n210 B.n96 10.6151
R1194 B.n211 B.n210 10.6151
R1195 B.n212 B.n211 10.6151
R1196 B.n212 B.n94 10.6151
R1197 B.n216 B.n94 10.6151
R1198 B.n217 B.n216 10.6151
R1199 B.n221 B.n217 10.6151
R1200 B.n225 B.n92 10.6151
R1201 B.n226 B.n225 10.6151
R1202 B.n227 B.n226 10.6151
R1203 B.n227 B.n90 10.6151
R1204 B.n231 B.n90 10.6151
R1205 B.n232 B.n231 10.6151
R1206 B.n233 B.n232 10.6151
R1207 B.n233 B.n88 10.6151
R1208 B.n237 B.n88 10.6151
R1209 B.n238 B.n237 10.6151
R1210 B.n239 B.n238 10.6151
R1211 B.n239 B.n86 10.6151
R1212 B.n243 B.n86 10.6151
R1213 B.n244 B.n243 10.6151
R1214 B.n245 B.n244 10.6151
R1215 B.n245 B.n84 10.6151
R1216 B.n249 B.n84 10.6151
R1217 B.n250 B.n249 10.6151
R1218 B.n251 B.n250 10.6151
R1219 B.n251 B.n82 10.6151
R1220 B.n255 B.n82 10.6151
R1221 B.n256 B.n255 10.6151
R1222 B.n257 B.n256 10.6151
R1223 B.n257 B.n80 10.6151
R1224 B.n261 B.n80 10.6151
R1225 B.n262 B.n261 10.6151
R1226 B.n263 B.n262 10.6151
R1227 B.n263 B.n78 10.6151
R1228 B.n267 B.n78 10.6151
R1229 B.n268 B.n267 10.6151
R1230 B.n269 B.n268 10.6151
R1231 B.n269 B.n76 10.6151
R1232 B.n273 B.n76 10.6151
R1233 B.n485 B.n0 8.11757
R1234 B.n485 B.n1 8.11757
R1235 B.n402 B.n401 6.5566
R1236 B.n389 B.n388 6.5566
R1237 B.n206 B.n205 6.5566
R1238 B.n221 B.n220 6.5566
R1239 B.n403 B.n402 4.05904
R1240 B.n388 B.n387 4.05904
R1241 B.n205 B.n204 4.05904
R1242 B.n220 B.n92 4.05904
R1243 VN.n1 VN.t3 381.038
R1244 VN.n7 VN.t0 381.038
R1245 VN.n2 VN.t2 358.86
R1246 VN.n4 VN.t4 358.86
R1247 VN.n8 VN.t5 358.86
R1248 VN.n10 VN.t1 358.86
R1249 VN.n5 VN.n4 161.3
R1250 VN.n11 VN.n10 161.3
R1251 VN.n9 VN.n6 161.3
R1252 VN.n3 VN.n0 161.3
R1253 VN.n7 VN.n6 44.862
R1254 VN.n1 VN.n0 44.862
R1255 VN VN.n11 39.6312
R1256 VN.n4 VN.n3 28.4823
R1257 VN.n10 VN.n9 28.4823
R1258 VN.n3 VN.n2 19.7187
R1259 VN.n9 VN.n8 19.7187
R1260 VN.n2 VN.n1 19.7081
R1261 VN.n8 VN.n7 19.7081
R1262 VN.n11 VN.n6 0.189894
R1263 VN.n5 VN.n0 0.189894
R1264 VN VN.n5 0.0516364
R1265 VDD2.n95 VDD2.n51 756.745
R1266 VDD2.n44 VDD2.n0 756.745
R1267 VDD2.n96 VDD2.n95 585
R1268 VDD2.n94 VDD2.n93 585
R1269 VDD2.n55 VDD2.n54 585
R1270 VDD2.n59 VDD2.n57 585
R1271 VDD2.n88 VDD2.n87 585
R1272 VDD2.n86 VDD2.n85 585
R1273 VDD2.n61 VDD2.n60 585
R1274 VDD2.n80 VDD2.n79 585
R1275 VDD2.n78 VDD2.n77 585
R1276 VDD2.n65 VDD2.n64 585
R1277 VDD2.n72 VDD2.n71 585
R1278 VDD2.n70 VDD2.n69 585
R1279 VDD2.n17 VDD2.n16 585
R1280 VDD2.n19 VDD2.n18 585
R1281 VDD2.n12 VDD2.n11 585
R1282 VDD2.n25 VDD2.n24 585
R1283 VDD2.n27 VDD2.n26 585
R1284 VDD2.n8 VDD2.n7 585
R1285 VDD2.n34 VDD2.n33 585
R1286 VDD2.n35 VDD2.n6 585
R1287 VDD2.n37 VDD2.n36 585
R1288 VDD2.n4 VDD2.n3 585
R1289 VDD2.n43 VDD2.n42 585
R1290 VDD2.n45 VDD2.n44 585
R1291 VDD2.n68 VDD2.t4 329.038
R1292 VDD2.n15 VDD2.t2 329.038
R1293 VDD2.n95 VDD2.n94 171.744
R1294 VDD2.n94 VDD2.n54 171.744
R1295 VDD2.n59 VDD2.n54 171.744
R1296 VDD2.n87 VDD2.n59 171.744
R1297 VDD2.n87 VDD2.n86 171.744
R1298 VDD2.n86 VDD2.n60 171.744
R1299 VDD2.n79 VDD2.n60 171.744
R1300 VDD2.n79 VDD2.n78 171.744
R1301 VDD2.n78 VDD2.n64 171.744
R1302 VDD2.n71 VDD2.n64 171.744
R1303 VDD2.n71 VDD2.n70 171.744
R1304 VDD2.n18 VDD2.n17 171.744
R1305 VDD2.n18 VDD2.n11 171.744
R1306 VDD2.n25 VDD2.n11 171.744
R1307 VDD2.n26 VDD2.n25 171.744
R1308 VDD2.n26 VDD2.n7 171.744
R1309 VDD2.n34 VDD2.n7 171.744
R1310 VDD2.n35 VDD2.n34 171.744
R1311 VDD2.n36 VDD2.n35 171.744
R1312 VDD2.n36 VDD2.n3 171.744
R1313 VDD2.n43 VDD2.n3 171.744
R1314 VDD2.n44 VDD2.n43 171.744
R1315 VDD2.n70 VDD2.t4 85.8723
R1316 VDD2.n17 VDD2.t2 85.8723
R1317 VDD2.n50 VDD2.n49 78.5599
R1318 VDD2 VDD2.n101 78.557
R1319 VDD2.n50 VDD2.n48 49.3002
R1320 VDD2.n100 VDD2.n99 48.6702
R1321 VDD2.n100 VDD2.n50 34.642
R1322 VDD2.n57 VDD2.n55 13.1884
R1323 VDD2.n37 VDD2.n4 13.1884
R1324 VDD2.n93 VDD2.n92 12.8005
R1325 VDD2.n89 VDD2.n88 12.8005
R1326 VDD2.n38 VDD2.n6 12.8005
R1327 VDD2.n42 VDD2.n41 12.8005
R1328 VDD2.n96 VDD2.n53 12.0247
R1329 VDD2.n85 VDD2.n58 12.0247
R1330 VDD2.n33 VDD2.n32 12.0247
R1331 VDD2.n45 VDD2.n2 12.0247
R1332 VDD2.n97 VDD2.n51 11.249
R1333 VDD2.n84 VDD2.n61 11.249
R1334 VDD2.n31 VDD2.n8 11.249
R1335 VDD2.n46 VDD2.n0 11.249
R1336 VDD2.n69 VDD2.n68 10.7239
R1337 VDD2.n16 VDD2.n15 10.7239
R1338 VDD2.n81 VDD2.n80 10.4732
R1339 VDD2.n28 VDD2.n27 10.4732
R1340 VDD2.n77 VDD2.n63 9.69747
R1341 VDD2.n24 VDD2.n10 9.69747
R1342 VDD2.n99 VDD2.n98 9.45567
R1343 VDD2.n48 VDD2.n47 9.45567
R1344 VDD2.n67 VDD2.n66 9.3005
R1345 VDD2.n74 VDD2.n73 9.3005
R1346 VDD2.n76 VDD2.n75 9.3005
R1347 VDD2.n63 VDD2.n62 9.3005
R1348 VDD2.n82 VDD2.n81 9.3005
R1349 VDD2.n84 VDD2.n83 9.3005
R1350 VDD2.n58 VDD2.n56 9.3005
R1351 VDD2.n90 VDD2.n89 9.3005
R1352 VDD2.n98 VDD2.n97 9.3005
R1353 VDD2.n53 VDD2.n52 9.3005
R1354 VDD2.n92 VDD2.n91 9.3005
R1355 VDD2.n47 VDD2.n46 9.3005
R1356 VDD2.n2 VDD2.n1 9.3005
R1357 VDD2.n41 VDD2.n40 9.3005
R1358 VDD2.n14 VDD2.n13 9.3005
R1359 VDD2.n21 VDD2.n20 9.3005
R1360 VDD2.n23 VDD2.n22 9.3005
R1361 VDD2.n10 VDD2.n9 9.3005
R1362 VDD2.n29 VDD2.n28 9.3005
R1363 VDD2.n31 VDD2.n30 9.3005
R1364 VDD2.n32 VDD2.n5 9.3005
R1365 VDD2.n39 VDD2.n38 9.3005
R1366 VDD2.n76 VDD2.n65 8.92171
R1367 VDD2.n23 VDD2.n12 8.92171
R1368 VDD2.n73 VDD2.n72 8.14595
R1369 VDD2.n20 VDD2.n19 8.14595
R1370 VDD2.n69 VDD2.n67 7.3702
R1371 VDD2.n16 VDD2.n14 7.3702
R1372 VDD2.n72 VDD2.n67 5.81868
R1373 VDD2.n19 VDD2.n14 5.81868
R1374 VDD2.n73 VDD2.n65 5.04292
R1375 VDD2.n20 VDD2.n12 5.04292
R1376 VDD2.n77 VDD2.n76 4.26717
R1377 VDD2.n24 VDD2.n23 4.26717
R1378 VDD2.n101 VDD2.t0 3.52217
R1379 VDD2.n101 VDD2.t5 3.52217
R1380 VDD2.n49 VDD2.t3 3.52217
R1381 VDD2.n49 VDD2.t1 3.52217
R1382 VDD2.n80 VDD2.n63 3.49141
R1383 VDD2.n27 VDD2.n10 3.49141
R1384 VDD2.n99 VDD2.n51 2.71565
R1385 VDD2.n81 VDD2.n61 2.71565
R1386 VDD2.n28 VDD2.n8 2.71565
R1387 VDD2.n48 VDD2.n0 2.71565
R1388 VDD2.n68 VDD2.n66 2.41283
R1389 VDD2.n15 VDD2.n13 2.41283
R1390 VDD2.n97 VDD2.n96 1.93989
R1391 VDD2.n85 VDD2.n84 1.93989
R1392 VDD2.n33 VDD2.n31 1.93989
R1393 VDD2.n46 VDD2.n45 1.93989
R1394 VDD2.n93 VDD2.n53 1.16414
R1395 VDD2.n88 VDD2.n58 1.16414
R1396 VDD2.n32 VDD2.n6 1.16414
R1397 VDD2.n42 VDD2.n2 1.16414
R1398 VDD2 VDD2.n100 0.744035
R1399 VDD2.n92 VDD2.n55 0.388379
R1400 VDD2.n89 VDD2.n57 0.388379
R1401 VDD2.n38 VDD2.n37 0.388379
R1402 VDD2.n41 VDD2.n4 0.388379
R1403 VDD2.n98 VDD2.n52 0.155672
R1404 VDD2.n91 VDD2.n52 0.155672
R1405 VDD2.n91 VDD2.n90 0.155672
R1406 VDD2.n90 VDD2.n56 0.155672
R1407 VDD2.n83 VDD2.n56 0.155672
R1408 VDD2.n83 VDD2.n82 0.155672
R1409 VDD2.n82 VDD2.n62 0.155672
R1410 VDD2.n75 VDD2.n62 0.155672
R1411 VDD2.n75 VDD2.n74 0.155672
R1412 VDD2.n74 VDD2.n66 0.155672
R1413 VDD2.n21 VDD2.n13 0.155672
R1414 VDD2.n22 VDD2.n21 0.155672
R1415 VDD2.n22 VDD2.n9 0.155672
R1416 VDD2.n29 VDD2.n9 0.155672
R1417 VDD2.n30 VDD2.n29 0.155672
R1418 VDD2.n30 VDD2.n5 0.155672
R1419 VDD2.n39 VDD2.n5 0.155672
R1420 VDD2.n40 VDD2.n39 0.155672
R1421 VDD2.n40 VDD2.n1 0.155672
R1422 VDD2.n47 VDD2.n1 0.155672
C0 VTAIL w_n1818_n2814# 2.49619f
C1 VDD1 w_n1818_n2814# 1.61226f
C2 w_n1818_n2814# VP 3.17391f
C3 VDD1 VTAIL 7.96148f
C4 VTAIL VP 3.30486f
C5 VDD1 VP 3.63253f
C6 VDD2 VN 3.48451f
C7 B VN 0.738092f
C8 VN w_n1818_n2814# 2.94408f
C9 VDD2 B 1.39652f
C10 VTAIL VN 3.29038f
C11 VDD1 VN 0.147992f
C12 VN VP 4.59675f
C13 VDD2 w_n1818_n2814# 1.6373f
C14 VDD2 VTAIL 7.99738f
C15 VDD2 VDD1 0.719587f
C16 VDD2 VP 0.29955f
C17 B w_n1818_n2814# 6.31796f
C18 VTAIL B 2.23165f
C19 VDD1 B 1.36684f
C20 B VP 1.1124f
C21 VDD2 VSUBS 1.206681f
C22 VDD1 VSUBS 1.059294f
C23 VTAIL VSUBS 0.683978f
C24 VN VSUBS 4.23738f
C25 VP VSUBS 1.387946f
C26 B VSUBS 2.548783f
C27 w_n1818_n2814# VSUBS 63.2882f
C28 VDD2.n0 VSUBS 0.023818f
C29 VDD2.n1 VSUBS 0.023293f
C30 VDD2.n2 VSUBS 0.012517f
C31 VDD2.n3 VSUBS 0.029585f
C32 VDD2.n4 VSUBS 0.012885f
C33 VDD2.n5 VSUBS 0.023293f
C34 VDD2.n6 VSUBS 0.013253f
C35 VDD2.n7 VSUBS 0.029585f
C36 VDD2.n8 VSUBS 0.013253f
C37 VDD2.n9 VSUBS 0.023293f
C38 VDD2.n10 VSUBS 0.012517f
C39 VDD2.n11 VSUBS 0.029585f
C40 VDD2.n12 VSUBS 0.013253f
C41 VDD2.n13 VSUBS 0.861706f
C42 VDD2.n14 VSUBS 0.012517f
C43 VDD2.t2 VSUBS 0.06356f
C44 VDD2.n15 VSUBS 0.154295f
C45 VDD2.n16 VSUBS 0.022255f
C46 VDD2.n17 VSUBS 0.022189f
C47 VDD2.n18 VSUBS 0.029585f
C48 VDD2.n19 VSUBS 0.013253f
C49 VDD2.n20 VSUBS 0.012517f
C50 VDD2.n21 VSUBS 0.023293f
C51 VDD2.n22 VSUBS 0.023293f
C52 VDD2.n23 VSUBS 0.012517f
C53 VDD2.n24 VSUBS 0.013253f
C54 VDD2.n25 VSUBS 0.029585f
C55 VDD2.n26 VSUBS 0.029585f
C56 VDD2.n27 VSUBS 0.013253f
C57 VDD2.n28 VSUBS 0.012517f
C58 VDD2.n29 VSUBS 0.023293f
C59 VDD2.n30 VSUBS 0.023293f
C60 VDD2.n31 VSUBS 0.012517f
C61 VDD2.n32 VSUBS 0.012517f
C62 VDD2.n33 VSUBS 0.013253f
C63 VDD2.n34 VSUBS 0.029585f
C64 VDD2.n35 VSUBS 0.029585f
C65 VDD2.n36 VSUBS 0.029585f
C66 VDD2.n37 VSUBS 0.012885f
C67 VDD2.n38 VSUBS 0.012517f
C68 VDD2.n39 VSUBS 0.023293f
C69 VDD2.n40 VSUBS 0.023293f
C70 VDD2.n41 VSUBS 0.012517f
C71 VDD2.n42 VSUBS 0.013253f
C72 VDD2.n43 VSUBS 0.029585f
C73 VDD2.n44 VSUBS 0.065573f
C74 VDD2.n45 VSUBS 0.013253f
C75 VDD2.n46 VSUBS 0.012517f
C76 VDD2.n47 VSUBS 0.053523f
C77 VDD2.n48 VSUBS 0.049969f
C78 VDD2.t3 VSUBS 0.169896f
C79 VDD2.t1 VSUBS 0.169896f
C80 VDD2.n49 VSUBS 1.26327f
C81 VDD2.n50 VSUBS 1.80418f
C82 VDD2.n51 VSUBS 0.023818f
C83 VDD2.n52 VSUBS 0.023293f
C84 VDD2.n53 VSUBS 0.012517f
C85 VDD2.n54 VSUBS 0.029585f
C86 VDD2.n55 VSUBS 0.012885f
C87 VDD2.n56 VSUBS 0.023293f
C88 VDD2.n57 VSUBS 0.012885f
C89 VDD2.n58 VSUBS 0.012517f
C90 VDD2.n59 VSUBS 0.029585f
C91 VDD2.n60 VSUBS 0.029585f
C92 VDD2.n61 VSUBS 0.013253f
C93 VDD2.n62 VSUBS 0.023293f
C94 VDD2.n63 VSUBS 0.012517f
C95 VDD2.n64 VSUBS 0.029585f
C96 VDD2.n65 VSUBS 0.013253f
C97 VDD2.n66 VSUBS 0.861705f
C98 VDD2.n67 VSUBS 0.012517f
C99 VDD2.t4 VSUBS 0.06356f
C100 VDD2.n68 VSUBS 0.154295f
C101 VDD2.n69 VSUBS 0.022255f
C102 VDD2.n70 VSUBS 0.022189f
C103 VDD2.n71 VSUBS 0.029585f
C104 VDD2.n72 VSUBS 0.013253f
C105 VDD2.n73 VSUBS 0.012517f
C106 VDD2.n74 VSUBS 0.023293f
C107 VDD2.n75 VSUBS 0.023293f
C108 VDD2.n76 VSUBS 0.012517f
C109 VDD2.n77 VSUBS 0.013253f
C110 VDD2.n78 VSUBS 0.029585f
C111 VDD2.n79 VSUBS 0.029585f
C112 VDD2.n80 VSUBS 0.013253f
C113 VDD2.n81 VSUBS 0.012517f
C114 VDD2.n82 VSUBS 0.023293f
C115 VDD2.n83 VSUBS 0.023293f
C116 VDD2.n84 VSUBS 0.012517f
C117 VDD2.n85 VSUBS 0.013253f
C118 VDD2.n86 VSUBS 0.029585f
C119 VDD2.n87 VSUBS 0.029585f
C120 VDD2.n88 VSUBS 0.013253f
C121 VDD2.n89 VSUBS 0.012517f
C122 VDD2.n90 VSUBS 0.023293f
C123 VDD2.n91 VSUBS 0.023293f
C124 VDD2.n92 VSUBS 0.012517f
C125 VDD2.n93 VSUBS 0.013253f
C126 VDD2.n94 VSUBS 0.029585f
C127 VDD2.n95 VSUBS 0.065573f
C128 VDD2.n96 VSUBS 0.013253f
C129 VDD2.n97 VSUBS 0.012517f
C130 VDD2.n98 VSUBS 0.053523f
C131 VDD2.n99 VSUBS 0.048783f
C132 VDD2.n100 VSUBS 1.70874f
C133 VDD2.t0 VSUBS 0.169896f
C134 VDD2.t5 VSUBS 0.169896f
C135 VDD2.n101 VSUBS 1.26325f
C136 VN.n0 VSUBS 0.240686f
C137 VN.t3 VSUBS 1.13532f
C138 VN.n1 VSUBS 0.441418f
C139 VN.t2 VSUBS 1.10838f
C140 VN.n2 VSUBS 0.467188f
C141 VN.n3 VSUBS 0.013019f
C142 VN.t4 VSUBS 1.10838f
C143 VN.n4 VSUBS 0.459343f
C144 VN.n5 VSUBS 0.044461f
C145 VN.n6 VSUBS 0.240686f
C146 VN.t0 VSUBS 1.13532f
C147 VN.n7 VSUBS 0.441418f
C148 VN.t5 VSUBS 1.10838f
C149 VN.n8 VSUBS 0.467188f
C150 VN.n9 VSUBS 0.013019f
C151 VN.t1 VSUBS 1.10838f
C152 VN.n10 VSUBS 0.459343f
C153 VN.n11 VSUBS 2.14749f
C154 B.n0 VSUBS 0.006778f
C155 B.n1 VSUBS 0.006778f
C156 B.n2 VSUBS 0.010024f
C157 B.n3 VSUBS 0.007682f
C158 B.n4 VSUBS 0.007682f
C159 B.n5 VSUBS 0.007682f
C160 B.n6 VSUBS 0.007682f
C161 B.n7 VSUBS 0.007682f
C162 B.n8 VSUBS 0.007682f
C163 B.n9 VSUBS 0.007682f
C164 B.n10 VSUBS 0.007682f
C165 B.n11 VSUBS 0.007682f
C166 B.n12 VSUBS 0.018001f
C167 B.n13 VSUBS 0.007682f
C168 B.n14 VSUBS 0.007682f
C169 B.n15 VSUBS 0.007682f
C170 B.n16 VSUBS 0.007682f
C171 B.n17 VSUBS 0.007682f
C172 B.n18 VSUBS 0.007682f
C173 B.n19 VSUBS 0.007682f
C174 B.n20 VSUBS 0.007682f
C175 B.n21 VSUBS 0.007682f
C176 B.n22 VSUBS 0.007682f
C177 B.n23 VSUBS 0.007682f
C178 B.n24 VSUBS 0.007682f
C179 B.n25 VSUBS 0.007682f
C180 B.n26 VSUBS 0.007682f
C181 B.n27 VSUBS 0.007682f
C182 B.n28 VSUBS 0.007682f
C183 B.n29 VSUBS 0.007682f
C184 B.t4 VSUBS 0.165966f
C185 B.t5 VSUBS 0.178593f
C186 B.t3 VSUBS 0.311212f
C187 B.n30 VSUBS 0.275715f
C188 B.n31 VSUBS 0.22357f
C189 B.n32 VSUBS 0.007682f
C190 B.n33 VSUBS 0.007682f
C191 B.n34 VSUBS 0.007682f
C192 B.n35 VSUBS 0.007682f
C193 B.t7 VSUBS 0.165969f
C194 B.t8 VSUBS 0.178595f
C195 B.t6 VSUBS 0.311212f
C196 B.n36 VSUBS 0.275712f
C197 B.n37 VSUBS 0.223567f
C198 B.n38 VSUBS 0.007682f
C199 B.n39 VSUBS 0.007682f
C200 B.n40 VSUBS 0.007682f
C201 B.n41 VSUBS 0.007682f
C202 B.n42 VSUBS 0.007682f
C203 B.n43 VSUBS 0.007682f
C204 B.n44 VSUBS 0.007682f
C205 B.n45 VSUBS 0.007682f
C206 B.n46 VSUBS 0.007682f
C207 B.n47 VSUBS 0.007682f
C208 B.n48 VSUBS 0.007682f
C209 B.n49 VSUBS 0.007682f
C210 B.n50 VSUBS 0.007682f
C211 B.n51 VSUBS 0.007682f
C212 B.n52 VSUBS 0.007682f
C213 B.n53 VSUBS 0.007682f
C214 B.n54 VSUBS 0.018001f
C215 B.n55 VSUBS 0.007682f
C216 B.n56 VSUBS 0.007682f
C217 B.n57 VSUBS 0.007682f
C218 B.n58 VSUBS 0.007682f
C219 B.n59 VSUBS 0.007682f
C220 B.n60 VSUBS 0.007682f
C221 B.n61 VSUBS 0.007682f
C222 B.n62 VSUBS 0.007682f
C223 B.n63 VSUBS 0.007682f
C224 B.n64 VSUBS 0.007682f
C225 B.n65 VSUBS 0.007682f
C226 B.n66 VSUBS 0.007682f
C227 B.n67 VSUBS 0.007682f
C228 B.n68 VSUBS 0.007682f
C229 B.n69 VSUBS 0.007682f
C230 B.n70 VSUBS 0.007682f
C231 B.n71 VSUBS 0.007682f
C232 B.n72 VSUBS 0.007682f
C233 B.n73 VSUBS 0.007682f
C234 B.n74 VSUBS 0.007682f
C235 B.n75 VSUBS 0.016567f
C236 B.n76 VSUBS 0.007682f
C237 B.n77 VSUBS 0.007682f
C238 B.n78 VSUBS 0.007682f
C239 B.n79 VSUBS 0.007682f
C240 B.n80 VSUBS 0.007682f
C241 B.n81 VSUBS 0.007682f
C242 B.n82 VSUBS 0.007682f
C243 B.n83 VSUBS 0.007682f
C244 B.n84 VSUBS 0.007682f
C245 B.n85 VSUBS 0.007682f
C246 B.n86 VSUBS 0.007682f
C247 B.n87 VSUBS 0.007682f
C248 B.n88 VSUBS 0.007682f
C249 B.n89 VSUBS 0.007682f
C250 B.n90 VSUBS 0.007682f
C251 B.n91 VSUBS 0.007682f
C252 B.n92 VSUBS 0.005309f
C253 B.n93 VSUBS 0.007682f
C254 B.n94 VSUBS 0.007682f
C255 B.n95 VSUBS 0.007682f
C256 B.n96 VSUBS 0.007682f
C257 B.n97 VSUBS 0.007682f
C258 B.t11 VSUBS 0.165966f
C259 B.t10 VSUBS 0.178593f
C260 B.t9 VSUBS 0.311212f
C261 B.n98 VSUBS 0.275715f
C262 B.n99 VSUBS 0.22357f
C263 B.n100 VSUBS 0.007682f
C264 B.n101 VSUBS 0.007682f
C265 B.n102 VSUBS 0.007682f
C266 B.n103 VSUBS 0.007682f
C267 B.n104 VSUBS 0.007682f
C268 B.n105 VSUBS 0.007682f
C269 B.n106 VSUBS 0.007682f
C270 B.n107 VSUBS 0.007682f
C271 B.n108 VSUBS 0.007682f
C272 B.n109 VSUBS 0.007682f
C273 B.n110 VSUBS 0.007682f
C274 B.n111 VSUBS 0.007682f
C275 B.n112 VSUBS 0.007682f
C276 B.n113 VSUBS 0.007682f
C277 B.n114 VSUBS 0.007682f
C278 B.n115 VSUBS 0.007682f
C279 B.n116 VSUBS 0.016567f
C280 B.n117 VSUBS 0.007682f
C281 B.n118 VSUBS 0.007682f
C282 B.n119 VSUBS 0.007682f
C283 B.n120 VSUBS 0.007682f
C284 B.n121 VSUBS 0.007682f
C285 B.n122 VSUBS 0.007682f
C286 B.n123 VSUBS 0.007682f
C287 B.n124 VSUBS 0.007682f
C288 B.n125 VSUBS 0.007682f
C289 B.n126 VSUBS 0.007682f
C290 B.n127 VSUBS 0.007682f
C291 B.n128 VSUBS 0.007682f
C292 B.n129 VSUBS 0.007682f
C293 B.n130 VSUBS 0.007682f
C294 B.n131 VSUBS 0.007682f
C295 B.n132 VSUBS 0.007682f
C296 B.n133 VSUBS 0.007682f
C297 B.n134 VSUBS 0.007682f
C298 B.n135 VSUBS 0.007682f
C299 B.n136 VSUBS 0.007682f
C300 B.n137 VSUBS 0.007682f
C301 B.n138 VSUBS 0.007682f
C302 B.n139 VSUBS 0.007682f
C303 B.n140 VSUBS 0.007682f
C304 B.n141 VSUBS 0.007682f
C305 B.n142 VSUBS 0.007682f
C306 B.n143 VSUBS 0.007682f
C307 B.n144 VSUBS 0.007682f
C308 B.n145 VSUBS 0.007682f
C309 B.n146 VSUBS 0.007682f
C310 B.n147 VSUBS 0.007682f
C311 B.n148 VSUBS 0.007682f
C312 B.n149 VSUBS 0.007682f
C313 B.n150 VSUBS 0.007682f
C314 B.n151 VSUBS 0.007682f
C315 B.n152 VSUBS 0.007682f
C316 B.n153 VSUBS 0.016567f
C317 B.n154 VSUBS 0.018001f
C318 B.n155 VSUBS 0.018001f
C319 B.n156 VSUBS 0.007682f
C320 B.n157 VSUBS 0.007682f
C321 B.n158 VSUBS 0.007682f
C322 B.n159 VSUBS 0.007682f
C323 B.n160 VSUBS 0.007682f
C324 B.n161 VSUBS 0.007682f
C325 B.n162 VSUBS 0.007682f
C326 B.n163 VSUBS 0.007682f
C327 B.n164 VSUBS 0.007682f
C328 B.n165 VSUBS 0.007682f
C329 B.n166 VSUBS 0.007682f
C330 B.n167 VSUBS 0.007682f
C331 B.n168 VSUBS 0.007682f
C332 B.n169 VSUBS 0.007682f
C333 B.n170 VSUBS 0.007682f
C334 B.n171 VSUBS 0.007682f
C335 B.n172 VSUBS 0.007682f
C336 B.n173 VSUBS 0.007682f
C337 B.n174 VSUBS 0.007682f
C338 B.n175 VSUBS 0.007682f
C339 B.n176 VSUBS 0.007682f
C340 B.n177 VSUBS 0.007682f
C341 B.n178 VSUBS 0.007682f
C342 B.n179 VSUBS 0.007682f
C343 B.n180 VSUBS 0.007682f
C344 B.n181 VSUBS 0.007682f
C345 B.n182 VSUBS 0.007682f
C346 B.n183 VSUBS 0.007682f
C347 B.n184 VSUBS 0.007682f
C348 B.n185 VSUBS 0.007682f
C349 B.n186 VSUBS 0.007682f
C350 B.n187 VSUBS 0.007682f
C351 B.n188 VSUBS 0.007682f
C352 B.n189 VSUBS 0.007682f
C353 B.n190 VSUBS 0.007682f
C354 B.n191 VSUBS 0.007682f
C355 B.n192 VSUBS 0.007682f
C356 B.n193 VSUBS 0.007682f
C357 B.n194 VSUBS 0.007682f
C358 B.n195 VSUBS 0.007682f
C359 B.n196 VSUBS 0.007682f
C360 B.n197 VSUBS 0.007682f
C361 B.n198 VSUBS 0.007682f
C362 B.n199 VSUBS 0.007682f
C363 B.n200 VSUBS 0.007682f
C364 B.n201 VSUBS 0.007682f
C365 B.n202 VSUBS 0.007682f
C366 B.n203 VSUBS 0.007682f
C367 B.n204 VSUBS 0.005309f
C368 B.n205 VSUBS 0.017798f
C369 B.n206 VSUBS 0.006213f
C370 B.n207 VSUBS 0.007682f
C371 B.n208 VSUBS 0.007682f
C372 B.n209 VSUBS 0.007682f
C373 B.n210 VSUBS 0.007682f
C374 B.n211 VSUBS 0.007682f
C375 B.n212 VSUBS 0.007682f
C376 B.n213 VSUBS 0.007682f
C377 B.n214 VSUBS 0.007682f
C378 B.n215 VSUBS 0.007682f
C379 B.n216 VSUBS 0.007682f
C380 B.n217 VSUBS 0.007682f
C381 B.t2 VSUBS 0.165969f
C382 B.t1 VSUBS 0.178595f
C383 B.t0 VSUBS 0.311212f
C384 B.n218 VSUBS 0.275712f
C385 B.n219 VSUBS 0.223567f
C386 B.n220 VSUBS 0.017798f
C387 B.n221 VSUBS 0.006213f
C388 B.n222 VSUBS 0.007682f
C389 B.n223 VSUBS 0.007682f
C390 B.n224 VSUBS 0.007682f
C391 B.n225 VSUBS 0.007682f
C392 B.n226 VSUBS 0.007682f
C393 B.n227 VSUBS 0.007682f
C394 B.n228 VSUBS 0.007682f
C395 B.n229 VSUBS 0.007682f
C396 B.n230 VSUBS 0.007682f
C397 B.n231 VSUBS 0.007682f
C398 B.n232 VSUBS 0.007682f
C399 B.n233 VSUBS 0.007682f
C400 B.n234 VSUBS 0.007682f
C401 B.n235 VSUBS 0.007682f
C402 B.n236 VSUBS 0.007682f
C403 B.n237 VSUBS 0.007682f
C404 B.n238 VSUBS 0.007682f
C405 B.n239 VSUBS 0.007682f
C406 B.n240 VSUBS 0.007682f
C407 B.n241 VSUBS 0.007682f
C408 B.n242 VSUBS 0.007682f
C409 B.n243 VSUBS 0.007682f
C410 B.n244 VSUBS 0.007682f
C411 B.n245 VSUBS 0.007682f
C412 B.n246 VSUBS 0.007682f
C413 B.n247 VSUBS 0.007682f
C414 B.n248 VSUBS 0.007682f
C415 B.n249 VSUBS 0.007682f
C416 B.n250 VSUBS 0.007682f
C417 B.n251 VSUBS 0.007682f
C418 B.n252 VSUBS 0.007682f
C419 B.n253 VSUBS 0.007682f
C420 B.n254 VSUBS 0.007682f
C421 B.n255 VSUBS 0.007682f
C422 B.n256 VSUBS 0.007682f
C423 B.n257 VSUBS 0.007682f
C424 B.n258 VSUBS 0.007682f
C425 B.n259 VSUBS 0.007682f
C426 B.n260 VSUBS 0.007682f
C427 B.n261 VSUBS 0.007682f
C428 B.n262 VSUBS 0.007682f
C429 B.n263 VSUBS 0.007682f
C430 B.n264 VSUBS 0.007682f
C431 B.n265 VSUBS 0.007682f
C432 B.n266 VSUBS 0.007682f
C433 B.n267 VSUBS 0.007682f
C434 B.n268 VSUBS 0.007682f
C435 B.n269 VSUBS 0.007682f
C436 B.n270 VSUBS 0.007682f
C437 B.n271 VSUBS 0.007682f
C438 B.n272 VSUBS 0.018001f
C439 B.n273 VSUBS 0.017037f
C440 B.n274 VSUBS 0.017531f
C441 B.n275 VSUBS 0.007682f
C442 B.n276 VSUBS 0.007682f
C443 B.n277 VSUBS 0.007682f
C444 B.n278 VSUBS 0.007682f
C445 B.n279 VSUBS 0.007682f
C446 B.n280 VSUBS 0.007682f
C447 B.n281 VSUBS 0.007682f
C448 B.n282 VSUBS 0.007682f
C449 B.n283 VSUBS 0.007682f
C450 B.n284 VSUBS 0.007682f
C451 B.n285 VSUBS 0.007682f
C452 B.n286 VSUBS 0.007682f
C453 B.n287 VSUBS 0.007682f
C454 B.n288 VSUBS 0.007682f
C455 B.n289 VSUBS 0.007682f
C456 B.n290 VSUBS 0.007682f
C457 B.n291 VSUBS 0.007682f
C458 B.n292 VSUBS 0.007682f
C459 B.n293 VSUBS 0.007682f
C460 B.n294 VSUBS 0.007682f
C461 B.n295 VSUBS 0.007682f
C462 B.n296 VSUBS 0.007682f
C463 B.n297 VSUBS 0.007682f
C464 B.n298 VSUBS 0.007682f
C465 B.n299 VSUBS 0.007682f
C466 B.n300 VSUBS 0.007682f
C467 B.n301 VSUBS 0.007682f
C468 B.n302 VSUBS 0.007682f
C469 B.n303 VSUBS 0.007682f
C470 B.n304 VSUBS 0.007682f
C471 B.n305 VSUBS 0.007682f
C472 B.n306 VSUBS 0.007682f
C473 B.n307 VSUBS 0.007682f
C474 B.n308 VSUBS 0.007682f
C475 B.n309 VSUBS 0.007682f
C476 B.n310 VSUBS 0.007682f
C477 B.n311 VSUBS 0.007682f
C478 B.n312 VSUBS 0.007682f
C479 B.n313 VSUBS 0.007682f
C480 B.n314 VSUBS 0.007682f
C481 B.n315 VSUBS 0.007682f
C482 B.n316 VSUBS 0.007682f
C483 B.n317 VSUBS 0.007682f
C484 B.n318 VSUBS 0.007682f
C485 B.n319 VSUBS 0.007682f
C486 B.n320 VSUBS 0.007682f
C487 B.n321 VSUBS 0.007682f
C488 B.n322 VSUBS 0.007682f
C489 B.n323 VSUBS 0.007682f
C490 B.n324 VSUBS 0.007682f
C491 B.n325 VSUBS 0.007682f
C492 B.n326 VSUBS 0.007682f
C493 B.n327 VSUBS 0.007682f
C494 B.n328 VSUBS 0.007682f
C495 B.n329 VSUBS 0.007682f
C496 B.n330 VSUBS 0.007682f
C497 B.n331 VSUBS 0.007682f
C498 B.n332 VSUBS 0.007682f
C499 B.n333 VSUBS 0.007682f
C500 B.n334 VSUBS 0.007682f
C501 B.n335 VSUBS 0.016567f
C502 B.n336 VSUBS 0.016567f
C503 B.n337 VSUBS 0.018001f
C504 B.n338 VSUBS 0.007682f
C505 B.n339 VSUBS 0.007682f
C506 B.n340 VSUBS 0.007682f
C507 B.n341 VSUBS 0.007682f
C508 B.n342 VSUBS 0.007682f
C509 B.n343 VSUBS 0.007682f
C510 B.n344 VSUBS 0.007682f
C511 B.n345 VSUBS 0.007682f
C512 B.n346 VSUBS 0.007682f
C513 B.n347 VSUBS 0.007682f
C514 B.n348 VSUBS 0.007682f
C515 B.n349 VSUBS 0.007682f
C516 B.n350 VSUBS 0.007682f
C517 B.n351 VSUBS 0.007682f
C518 B.n352 VSUBS 0.007682f
C519 B.n353 VSUBS 0.007682f
C520 B.n354 VSUBS 0.007682f
C521 B.n355 VSUBS 0.007682f
C522 B.n356 VSUBS 0.007682f
C523 B.n357 VSUBS 0.007682f
C524 B.n358 VSUBS 0.007682f
C525 B.n359 VSUBS 0.007682f
C526 B.n360 VSUBS 0.007682f
C527 B.n361 VSUBS 0.007682f
C528 B.n362 VSUBS 0.007682f
C529 B.n363 VSUBS 0.007682f
C530 B.n364 VSUBS 0.007682f
C531 B.n365 VSUBS 0.007682f
C532 B.n366 VSUBS 0.007682f
C533 B.n367 VSUBS 0.007682f
C534 B.n368 VSUBS 0.007682f
C535 B.n369 VSUBS 0.007682f
C536 B.n370 VSUBS 0.007682f
C537 B.n371 VSUBS 0.007682f
C538 B.n372 VSUBS 0.007682f
C539 B.n373 VSUBS 0.007682f
C540 B.n374 VSUBS 0.007682f
C541 B.n375 VSUBS 0.007682f
C542 B.n376 VSUBS 0.007682f
C543 B.n377 VSUBS 0.007682f
C544 B.n378 VSUBS 0.007682f
C545 B.n379 VSUBS 0.007682f
C546 B.n380 VSUBS 0.007682f
C547 B.n381 VSUBS 0.007682f
C548 B.n382 VSUBS 0.007682f
C549 B.n383 VSUBS 0.007682f
C550 B.n384 VSUBS 0.007682f
C551 B.n385 VSUBS 0.007682f
C552 B.n386 VSUBS 0.007682f
C553 B.n387 VSUBS 0.005309f
C554 B.n388 VSUBS 0.017798f
C555 B.n389 VSUBS 0.006213f
C556 B.n390 VSUBS 0.007682f
C557 B.n391 VSUBS 0.007682f
C558 B.n392 VSUBS 0.007682f
C559 B.n393 VSUBS 0.007682f
C560 B.n394 VSUBS 0.007682f
C561 B.n395 VSUBS 0.007682f
C562 B.n396 VSUBS 0.007682f
C563 B.n397 VSUBS 0.007682f
C564 B.n398 VSUBS 0.007682f
C565 B.n399 VSUBS 0.007682f
C566 B.n400 VSUBS 0.007682f
C567 B.n401 VSUBS 0.006213f
C568 B.n402 VSUBS 0.017798f
C569 B.n403 VSUBS 0.005309f
C570 B.n404 VSUBS 0.007682f
C571 B.n405 VSUBS 0.007682f
C572 B.n406 VSUBS 0.007682f
C573 B.n407 VSUBS 0.007682f
C574 B.n408 VSUBS 0.007682f
C575 B.n409 VSUBS 0.007682f
C576 B.n410 VSUBS 0.007682f
C577 B.n411 VSUBS 0.007682f
C578 B.n412 VSUBS 0.007682f
C579 B.n413 VSUBS 0.007682f
C580 B.n414 VSUBS 0.007682f
C581 B.n415 VSUBS 0.007682f
C582 B.n416 VSUBS 0.007682f
C583 B.n417 VSUBS 0.007682f
C584 B.n418 VSUBS 0.007682f
C585 B.n419 VSUBS 0.007682f
C586 B.n420 VSUBS 0.007682f
C587 B.n421 VSUBS 0.007682f
C588 B.n422 VSUBS 0.007682f
C589 B.n423 VSUBS 0.007682f
C590 B.n424 VSUBS 0.007682f
C591 B.n425 VSUBS 0.007682f
C592 B.n426 VSUBS 0.007682f
C593 B.n427 VSUBS 0.007682f
C594 B.n428 VSUBS 0.007682f
C595 B.n429 VSUBS 0.007682f
C596 B.n430 VSUBS 0.007682f
C597 B.n431 VSUBS 0.007682f
C598 B.n432 VSUBS 0.007682f
C599 B.n433 VSUBS 0.007682f
C600 B.n434 VSUBS 0.007682f
C601 B.n435 VSUBS 0.007682f
C602 B.n436 VSUBS 0.007682f
C603 B.n437 VSUBS 0.007682f
C604 B.n438 VSUBS 0.007682f
C605 B.n439 VSUBS 0.007682f
C606 B.n440 VSUBS 0.007682f
C607 B.n441 VSUBS 0.007682f
C608 B.n442 VSUBS 0.007682f
C609 B.n443 VSUBS 0.007682f
C610 B.n444 VSUBS 0.007682f
C611 B.n445 VSUBS 0.007682f
C612 B.n446 VSUBS 0.007682f
C613 B.n447 VSUBS 0.007682f
C614 B.n448 VSUBS 0.007682f
C615 B.n449 VSUBS 0.007682f
C616 B.n450 VSUBS 0.007682f
C617 B.n451 VSUBS 0.007682f
C618 B.n452 VSUBS 0.007682f
C619 B.n453 VSUBS 0.018001f
C620 B.n454 VSUBS 0.016567f
C621 B.n455 VSUBS 0.016567f
C622 B.n456 VSUBS 0.007682f
C623 B.n457 VSUBS 0.007682f
C624 B.n458 VSUBS 0.007682f
C625 B.n459 VSUBS 0.007682f
C626 B.n460 VSUBS 0.007682f
C627 B.n461 VSUBS 0.007682f
C628 B.n462 VSUBS 0.007682f
C629 B.n463 VSUBS 0.007682f
C630 B.n464 VSUBS 0.007682f
C631 B.n465 VSUBS 0.007682f
C632 B.n466 VSUBS 0.007682f
C633 B.n467 VSUBS 0.007682f
C634 B.n468 VSUBS 0.007682f
C635 B.n469 VSUBS 0.007682f
C636 B.n470 VSUBS 0.007682f
C637 B.n471 VSUBS 0.007682f
C638 B.n472 VSUBS 0.007682f
C639 B.n473 VSUBS 0.007682f
C640 B.n474 VSUBS 0.007682f
C641 B.n475 VSUBS 0.007682f
C642 B.n476 VSUBS 0.007682f
C643 B.n477 VSUBS 0.007682f
C644 B.n478 VSUBS 0.007682f
C645 B.n479 VSUBS 0.007682f
C646 B.n480 VSUBS 0.007682f
C647 B.n481 VSUBS 0.007682f
C648 B.n482 VSUBS 0.007682f
C649 B.n483 VSUBS 0.010024f
C650 B.n484 VSUBS 0.010679f
C651 B.n485 VSUBS 0.021235f
C652 VDD1.n0 VSUBS 0.023847f
C653 VDD1.n1 VSUBS 0.023321f
C654 VDD1.n2 VSUBS 0.012532f
C655 VDD1.n3 VSUBS 0.029621f
C656 VDD1.n4 VSUBS 0.0129f
C657 VDD1.n5 VSUBS 0.023321f
C658 VDD1.n6 VSUBS 0.0129f
C659 VDD1.n7 VSUBS 0.012532f
C660 VDD1.n8 VSUBS 0.029621f
C661 VDD1.n9 VSUBS 0.029621f
C662 VDD1.n10 VSUBS 0.013269f
C663 VDD1.n11 VSUBS 0.023321f
C664 VDD1.n12 VSUBS 0.012532f
C665 VDD1.n13 VSUBS 0.029621f
C666 VDD1.n14 VSUBS 0.013269f
C667 VDD1.n15 VSUBS 0.862744f
C668 VDD1.n16 VSUBS 0.012532f
C669 VDD1.t5 VSUBS 0.063637f
C670 VDD1.n17 VSUBS 0.154481f
C671 VDD1.n18 VSUBS 0.022282f
C672 VDD1.n19 VSUBS 0.022216f
C673 VDD1.n20 VSUBS 0.029621f
C674 VDD1.n21 VSUBS 0.013269f
C675 VDD1.n22 VSUBS 0.012532f
C676 VDD1.n23 VSUBS 0.023321f
C677 VDD1.n24 VSUBS 0.023321f
C678 VDD1.n25 VSUBS 0.012532f
C679 VDD1.n26 VSUBS 0.013269f
C680 VDD1.n27 VSUBS 0.029621f
C681 VDD1.n28 VSUBS 0.029621f
C682 VDD1.n29 VSUBS 0.013269f
C683 VDD1.n30 VSUBS 0.012532f
C684 VDD1.n31 VSUBS 0.023321f
C685 VDD1.n32 VSUBS 0.023321f
C686 VDD1.n33 VSUBS 0.012532f
C687 VDD1.n34 VSUBS 0.013269f
C688 VDD1.n35 VSUBS 0.029621f
C689 VDD1.n36 VSUBS 0.029621f
C690 VDD1.n37 VSUBS 0.013269f
C691 VDD1.n38 VSUBS 0.012532f
C692 VDD1.n39 VSUBS 0.023321f
C693 VDD1.n40 VSUBS 0.023321f
C694 VDD1.n41 VSUBS 0.012532f
C695 VDD1.n42 VSUBS 0.013269f
C696 VDD1.n43 VSUBS 0.029621f
C697 VDD1.n44 VSUBS 0.065652f
C698 VDD1.n45 VSUBS 0.013269f
C699 VDD1.n46 VSUBS 0.012532f
C700 VDD1.n47 VSUBS 0.053587f
C701 VDD1.n48 VSUBS 0.050356f
C702 VDD1.n49 VSUBS 0.023847f
C703 VDD1.n50 VSUBS 0.023321f
C704 VDD1.n51 VSUBS 0.012532f
C705 VDD1.n52 VSUBS 0.029621f
C706 VDD1.n53 VSUBS 0.0129f
C707 VDD1.n54 VSUBS 0.023321f
C708 VDD1.n55 VSUBS 0.013269f
C709 VDD1.n56 VSUBS 0.029621f
C710 VDD1.n57 VSUBS 0.013269f
C711 VDD1.n58 VSUBS 0.023321f
C712 VDD1.n59 VSUBS 0.012532f
C713 VDD1.n60 VSUBS 0.029621f
C714 VDD1.n61 VSUBS 0.013269f
C715 VDD1.n62 VSUBS 0.862744f
C716 VDD1.n63 VSUBS 0.012532f
C717 VDD1.t2 VSUBS 0.063637f
C718 VDD1.n64 VSUBS 0.154481f
C719 VDD1.n65 VSUBS 0.022282f
C720 VDD1.n66 VSUBS 0.022216f
C721 VDD1.n67 VSUBS 0.029621f
C722 VDD1.n68 VSUBS 0.013269f
C723 VDD1.n69 VSUBS 0.012532f
C724 VDD1.n70 VSUBS 0.023321f
C725 VDD1.n71 VSUBS 0.023321f
C726 VDD1.n72 VSUBS 0.012532f
C727 VDD1.n73 VSUBS 0.013269f
C728 VDD1.n74 VSUBS 0.029621f
C729 VDD1.n75 VSUBS 0.029621f
C730 VDD1.n76 VSUBS 0.013269f
C731 VDD1.n77 VSUBS 0.012532f
C732 VDD1.n78 VSUBS 0.023321f
C733 VDD1.n79 VSUBS 0.023321f
C734 VDD1.n80 VSUBS 0.012532f
C735 VDD1.n81 VSUBS 0.012532f
C736 VDD1.n82 VSUBS 0.013269f
C737 VDD1.n83 VSUBS 0.029621f
C738 VDD1.n84 VSUBS 0.029621f
C739 VDD1.n85 VSUBS 0.029621f
C740 VDD1.n86 VSUBS 0.0129f
C741 VDD1.n87 VSUBS 0.012532f
C742 VDD1.n88 VSUBS 0.023321f
C743 VDD1.n89 VSUBS 0.023321f
C744 VDD1.n90 VSUBS 0.012532f
C745 VDD1.n91 VSUBS 0.013269f
C746 VDD1.n92 VSUBS 0.029621f
C747 VDD1.n93 VSUBS 0.065652f
C748 VDD1.n94 VSUBS 0.013269f
C749 VDD1.n95 VSUBS 0.012532f
C750 VDD1.n96 VSUBS 0.053587f
C751 VDD1.n97 VSUBS 0.05003f
C752 VDD1.t3 VSUBS 0.170101f
C753 VDD1.t1 VSUBS 0.170101f
C754 VDD1.n98 VSUBS 1.2648f
C755 VDD1.n99 VSUBS 1.87798f
C756 VDD1.t0 VSUBS 0.170101f
C757 VDD1.t4 VSUBS 0.170101f
C758 VDD1.n100 VSUBS 1.26368f
C759 VDD1.n101 VSUBS 2.12978f
C760 VTAIL.t4 VSUBS 0.218173f
C761 VTAIL.t5 VSUBS 0.218173f
C762 VTAIL.n0 VSUBS 1.47876f
C763 VTAIL.n1 VSUBS 0.749601f
C764 VTAIL.n2 VSUBS 0.030586f
C765 VTAIL.n3 VSUBS 0.029912f
C766 VTAIL.n4 VSUBS 0.016073f
C767 VTAIL.n5 VSUBS 0.037992f
C768 VTAIL.n6 VSUBS 0.016546f
C769 VTAIL.n7 VSUBS 0.029912f
C770 VTAIL.n8 VSUBS 0.017019f
C771 VTAIL.n9 VSUBS 0.037992f
C772 VTAIL.n10 VSUBS 0.017019f
C773 VTAIL.n11 VSUBS 0.029912f
C774 VTAIL.n12 VSUBS 0.016073f
C775 VTAIL.n13 VSUBS 0.037992f
C776 VTAIL.n14 VSUBS 0.017019f
C777 VTAIL.n15 VSUBS 1.10657f
C778 VTAIL.n16 VSUBS 0.016073f
C779 VTAIL.t11 VSUBS 0.081622f
C780 VTAIL.n17 VSUBS 0.198139f
C781 VTAIL.n18 VSUBS 0.028579f
C782 VTAIL.n19 VSUBS 0.028494f
C783 VTAIL.n20 VSUBS 0.037992f
C784 VTAIL.n21 VSUBS 0.017019f
C785 VTAIL.n22 VSUBS 0.016073f
C786 VTAIL.n23 VSUBS 0.029912f
C787 VTAIL.n24 VSUBS 0.029912f
C788 VTAIL.n25 VSUBS 0.016073f
C789 VTAIL.n26 VSUBS 0.017019f
C790 VTAIL.n27 VSUBS 0.037992f
C791 VTAIL.n28 VSUBS 0.037992f
C792 VTAIL.n29 VSUBS 0.017019f
C793 VTAIL.n30 VSUBS 0.016073f
C794 VTAIL.n31 VSUBS 0.029912f
C795 VTAIL.n32 VSUBS 0.029912f
C796 VTAIL.n33 VSUBS 0.016073f
C797 VTAIL.n34 VSUBS 0.016073f
C798 VTAIL.n35 VSUBS 0.017019f
C799 VTAIL.n36 VSUBS 0.037992f
C800 VTAIL.n37 VSUBS 0.037992f
C801 VTAIL.n38 VSUBS 0.037992f
C802 VTAIL.n39 VSUBS 0.016546f
C803 VTAIL.n40 VSUBS 0.016073f
C804 VTAIL.n41 VSUBS 0.029912f
C805 VTAIL.n42 VSUBS 0.029912f
C806 VTAIL.n43 VSUBS 0.016073f
C807 VTAIL.n44 VSUBS 0.017019f
C808 VTAIL.n45 VSUBS 0.037992f
C809 VTAIL.n46 VSUBS 0.084206f
C810 VTAIL.n47 VSUBS 0.017019f
C811 VTAIL.n48 VSUBS 0.016073f
C812 VTAIL.n49 VSUBS 0.068732f
C813 VTAIL.n50 VSUBS 0.041989f
C814 VTAIL.n51 VSUBS 0.202712f
C815 VTAIL.t8 VSUBS 0.218173f
C816 VTAIL.t9 VSUBS 0.218173f
C817 VTAIL.n52 VSUBS 1.47876f
C818 VTAIL.n53 VSUBS 2.07011f
C819 VTAIL.t0 VSUBS 0.218173f
C820 VTAIL.t2 VSUBS 0.218173f
C821 VTAIL.n54 VSUBS 1.47877f
C822 VTAIL.n55 VSUBS 2.0701f
C823 VTAIL.n56 VSUBS 0.030586f
C824 VTAIL.n57 VSUBS 0.029912f
C825 VTAIL.n58 VSUBS 0.016073f
C826 VTAIL.n59 VSUBS 0.037992f
C827 VTAIL.n60 VSUBS 0.016546f
C828 VTAIL.n61 VSUBS 0.029912f
C829 VTAIL.n62 VSUBS 0.016546f
C830 VTAIL.n63 VSUBS 0.016073f
C831 VTAIL.n64 VSUBS 0.037992f
C832 VTAIL.n65 VSUBS 0.037992f
C833 VTAIL.n66 VSUBS 0.017019f
C834 VTAIL.n67 VSUBS 0.029912f
C835 VTAIL.n68 VSUBS 0.016073f
C836 VTAIL.n69 VSUBS 0.037992f
C837 VTAIL.n70 VSUBS 0.017019f
C838 VTAIL.n71 VSUBS 1.10657f
C839 VTAIL.n72 VSUBS 0.016073f
C840 VTAIL.t1 VSUBS 0.081622f
C841 VTAIL.n73 VSUBS 0.198139f
C842 VTAIL.n74 VSUBS 0.028579f
C843 VTAIL.n75 VSUBS 0.028494f
C844 VTAIL.n76 VSUBS 0.037992f
C845 VTAIL.n77 VSUBS 0.017019f
C846 VTAIL.n78 VSUBS 0.016073f
C847 VTAIL.n79 VSUBS 0.029912f
C848 VTAIL.n80 VSUBS 0.029912f
C849 VTAIL.n81 VSUBS 0.016073f
C850 VTAIL.n82 VSUBS 0.017019f
C851 VTAIL.n83 VSUBS 0.037992f
C852 VTAIL.n84 VSUBS 0.037992f
C853 VTAIL.n85 VSUBS 0.017019f
C854 VTAIL.n86 VSUBS 0.016073f
C855 VTAIL.n87 VSUBS 0.029912f
C856 VTAIL.n88 VSUBS 0.029912f
C857 VTAIL.n89 VSUBS 0.016073f
C858 VTAIL.n90 VSUBS 0.017019f
C859 VTAIL.n91 VSUBS 0.037992f
C860 VTAIL.n92 VSUBS 0.037992f
C861 VTAIL.n93 VSUBS 0.017019f
C862 VTAIL.n94 VSUBS 0.016073f
C863 VTAIL.n95 VSUBS 0.029912f
C864 VTAIL.n96 VSUBS 0.029912f
C865 VTAIL.n97 VSUBS 0.016073f
C866 VTAIL.n98 VSUBS 0.017019f
C867 VTAIL.n99 VSUBS 0.037992f
C868 VTAIL.n100 VSUBS 0.084206f
C869 VTAIL.n101 VSUBS 0.017019f
C870 VTAIL.n102 VSUBS 0.016073f
C871 VTAIL.n103 VSUBS 0.068732f
C872 VTAIL.n104 VSUBS 0.041989f
C873 VTAIL.n105 VSUBS 0.202712f
C874 VTAIL.t6 VSUBS 0.218173f
C875 VTAIL.t7 VSUBS 0.218173f
C876 VTAIL.n106 VSUBS 1.47877f
C877 VTAIL.n107 VSUBS 0.810038f
C878 VTAIL.n108 VSUBS 0.030586f
C879 VTAIL.n109 VSUBS 0.029912f
C880 VTAIL.n110 VSUBS 0.016073f
C881 VTAIL.n111 VSUBS 0.037992f
C882 VTAIL.n112 VSUBS 0.016546f
C883 VTAIL.n113 VSUBS 0.029912f
C884 VTAIL.n114 VSUBS 0.016546f
C885 VTAIL.n115 VSUBS 0.016073f
C886 VTAIL.n116 VSUBS 0.037992f
C887 VTAIL.n117 VSUBS 0.037992f
C888 VTAIL.n118 VSUBS 0.017019f
C889 VTAIL.n119 VSUBS 0.029912f
C890 VTAIL.n120 VSUBS 0.016073f
C891 VTAIL.n121 VSUBS 0.037992f
C892 VTAIL.n122 VSUBS 0.017019f
C893 VTAIL.n123 VSUBS 1.10657f
C894 VTAIL.n124 VSUBS 0.016073f
C895 VTAIL.t10 VSUBS 0.081622f
C896 VTAIL.n125 VSUBS 0.198139f
C897 VTAIL.n126 VSUBS 0.028579f
C898 VTAIL.n127 VSUBS 0.028494f
C899 VTAIL.n128 VSUBS 0.037992f
C900 VTAIL.n129 VSUBS 0.017019f
C901 VTAIL.n130 VSUBS 0.016073f
C902 VTAIL.n131 VSUBS 0.029912f
C903 VTAIL.n132 VSUBS 0.029912f
C904 VTAIL.n133 VSUBS 0.016073f
C905 VTAIL.n134 VSUBS 0.017019f
C906 VTAIL.n135 VSUBS 0.037992f
C907 VTAIL.n136 VSUBS 0.037992f
C908 VTAIL.n137 VSUBS 0.017019f
C909 VTAIL.n138 VSUBS 0.016073f
C910 VTAIL.n139 VSUBS 0.029912f
C911 VTAIL.n140 VSUBS 0.029912f
C912 VTAIL.n141 VSUBS 0.016073f
C913 VTAIL.n142 VSUBS 0.017019f
C914 VTAIL.n143 VSUBS 0.037992f
C915 VTAIL.n144 VSUBS 0.037992f
C916 VTAIL.n145 VSUBS 0.017019f
C917 VTAIL.n146 VSUBS 0.016073f
C918 VTAIL.n147 VSUBS 0.029912f
C919 VTAIL.n148 VSUBS 0.029912f
C920 VTAIL.n149 VSUBS 0.016073f
C921 VTAIL.n150 VSUBS 0.017019f
C922 VTAIL.n151 VSUBS 0.037992f
C923 VTAIL.n152 VSUBS 0.084206f
C924 VTAIL.n153 VSUBS 0.017019f
C925 VTAIL.n154 VSUBS 0.016073f
C926 VTAIL.n155 VSUBS 0.068732f
C927 VTAIL.n156 VSUBS 0.041989f
C928 VTAIL.n157 VSUBS 1.3747f
C929 VTAIL.n158 VSUBS 0.030586f
C930 VTAIL.n159 VSUBS 0.029912f
C931 VTAIL.n160 VSUBS 0.016073f
C932 VTAIL.n161 VSUBS 0.037992f
C933 VTAIL.n162 VSUBS 0.016546f
C934 VTAIL.n163 VSUBS 0.029912f
C935 VTAIL.n164 VSUBS 0.017019f
C936 VTAIL.n165 VSUBS 0.037992f
C937 VTAIL.n166 VSUBS 0.017019f
C938 VTAIL.n167 VSUBS 0.029912f
C939 VTAIL.n168 VSUBS 0.016073f
C940 VTAIL.n169 VSUBS 0.037992f
C941 VTAIL.n170 VSUBS 0.017019f
C942 VTAIL.n171 VSUBS 1.10657f
C943 VTAIL.n172 VSUBS 0.016073f
C944 VTAIL.t3 VSUBS 0.081622f
C945 VTAIL.n173 VSUBS 0.198139f
C946 VTAIL.n174 VSUBS 0.028579f
C947 VTAIL.n175 VSUBS 0.028494f
C948 VTAIL.n176 VSUBS 0.037992f
C949 VTAIL.n177 VSUBS 0.017019f
C950 VTAIL.n178 VSUBS 0.016073f
C951 VTAIL.n179 VSUBS 0.029912f
C952 VTAIL.n180 VSUBS 0.029912f
C953 VTAIL.n181 VSUBS 0.016073f
C954 VTAIL.n182 VSUBS 0.017019f
C955 VTAIL.n183 VSUBS 0.037992f
C956 VTAIL.n184 VSUBS 0.037992f
C957 VTAIL.n185 VSUBS 0.017019f
C958 VTAIL.n186 VSUBS 0.016073f
C959 VTAIL.n187 VSUBS 0.029912f
C960 VTAIL.n188 VSUBS 0.029912f
C961 VTAIL.n189 VSUBS 0.016073f
C962 VTAIL.n190 VSUBS 0.016073f
C963 VTAIL.n191 VSUBS 0.017019f
C964 VTAIL.n192 VSUBS 0.037992f
C965 VTAIL.n193 VSUBS 0.037992f
C966 VTAIL.n194 VSUBS 0.037992f
C967 VTAIL.n195 VSUBS 0.016546f
C968 VTAIL.n196 VSUBS 0.016073f
C969 VTAIL.n197 VSUBS 0.029912f
C970 VTAIL.n198 VSUBS 0.029912f
C971 VTAIL.n199 VSUBS 0.016073f
C972 VTAIL.n200 VSUBS 0.017019f
C973 VTAIL.n201 VSUBS 0.037992f
C974 VTAIL.n202 VSUBS 0.084206f
C975 VTAIL.n203 VSUBS 0.017019f
C976 VTAIL.n204 VSUBS 0.016073f
C977 VTAIL.n205 VSUBS 0.068732f
C978 VTAIL.n206 VSUBS 0.041989f
C979 VTAIL.n207 VSUBS 1.34707f
C980 VP.n0 VSUBS 0.059311f
C981 VP.n1 VSUBS 0.013459f
C982 VP.n2 VSUBS 0.248822f
C983 VP.t1 VSUBS 1.14585f
C984 VP.t5 VSUBS 1.14585f
C985 VP.t0 VSUBS 1.17369f
C986 VP.n3 VSUBS 0.456339f
C987 VP.n4 VSUBS 0.48298f
C988 VP.n5 VSUBS 0.013459f
C989 VP.n6 VSUBS 0.47487f
C990 VP.n7 VSUBS 2.18098f
C991 VP.t3 VSUBS 1.14585f
C992 VP.n8 VSUBS 0.47487f
C993 VP.n9 VSUBS 2.2353f
C994 VP.n10 VSUBS 0.059311f
C995 VP.n11 VSUBS 0.059311f
C996 VP.t2 VSUBS 1.14585f
C997 VP.n12 VSUBS 0.477613f
C998 VP.n13 VSUBS 0.013459f
C999 VP.t4 VSUBS 1.14585f
C1000 VP.n14 VSUBS 0.47487f
C1001 VP.n15 VSUBS 0.045964f
.ends

