* NGSPICE file created from diff_pair_sample_0500.ext - technology: sky130A

.subckt diff_pair_sample_0500 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=1.68
X1 VTAIL.t15 VP.t0 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=1.68
X2 VDD1.t6 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X3 VTAIL.t13 VP.t2 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X4 VDD1.t2 VP.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=1.68
X5 VTAIL.t11 VP.t4 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X6 VTAIL.t5 VN.t0 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=1.68
X7 VDD1.t4 VP.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X8 VDD1.t3 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=1.68
X9 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X10 VDD2.t5 VN.t2 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=1.68
X11 VTAIL.t4 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=1.68
X12 VDD2.t3 VN.t4 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=1.68
X13 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=1.68
X14 VDD2.t2 VN.t5 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X15 VTAIL.t6 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=1.68
X17 VTAIL.t8 VP.t7 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=1.68
X18 VDD2.t0 VN.t7 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=1.68
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=1.68
R0 B.n638 B.n637 585
R1 B.n639 B.n638 585
R2 B.n236 B.n103 585
R3 B.n235 B.n234 585
R4 B.n233 B.n232 585
R5 B.n231 B.n230 585
R6 B.n229 B.n228 585
R7 B.n227 B.n226 585
R8 B.n225 B.n224 585
R9 B.n223 B.n222 585
R10 B.n221 B.n220 585
R11 B.n219 B.n218 585
R12 B.n217 B.n216 585
R13 B.n215 B.n214 585
R14 B.n213 B.n212 585
R15 B.n211 B.n210 585
R16 B.n209 B.n208 585
R17 B.n207 B.n206 585
R18 B.n205 B.n204 585
R19 B.n203 B.n202 585
R20 B.n201 B.n200 585
R21 B.n199 B.n198 585
R22 B.n197 B.n196 585
R23 B.n195 B.n194 585
R24 B.n193 B.n192 585
R25 B.n191 B.n190 585
R26 B.n189 B.n188 585
R27 B.n187 B.n186 585
R28 B.n185 B.n184 585
R29 B.n182 B.n181 585
R30 B.n180 B.n179 585
R31 B.n178 B.n177 585
R32 B.n176 B.n175 585
R33 B.n174 B.n173 585
R34 B.n172 B.n171 585
R35 B.n170 B.n169 585
R36 B.n168 B.n167 585
R37 B.n166 B.n165 585
R38 B.n164 B.n163 585
R39 B.n162 B.n161 585
R40 B.n160 B.n159 585
R41 B.n158 B.n157 585
R42 B.n156 B.n155 585
R43 B.n154 B.n153 585
R44 B.n152 B.n151 585
R45 B.n150 B.n149 585
R46 B.n148 B.n147 585
R47 B.n146 B.n145 585
R48 B.n144 B.n143 585
R49 B.n142 B.n141 585
R50 B.n140 B.n139 585
R51 B.n138 B.n137 585
R52 B.n136 B.n135 585
R53 B.n134 B.n133 585
R54 B.n132 B.n131 585
R55 B.n130 B.n129 585
R56 B.n128 B.n127 585
R57 B.n126 B.n125 585
R58 B.n124 B.n123 585
R59 B.n122 B.n121 585
R60 B.n120 B.n119 585
R61 B.n118 B.n117 585
R62 B.n116 B.n115 585
R63 B.n114 B.n113 585
R64 B.n112 B.n111 585
R65 B.n110 B.n109 585
R66 B.n636 B.n70 585
R67 B.n640 B.n70 585
R68 B.n635 B.n69 585
R69 B.n641 B.n69 585
R70 B.n634 B.n633 585
R71 B.n633 B.n65 585
R72 B.n632 B.n64 585
R73 B.n647 B.n64 585
R74 B.n631 B.n63 585
R75 B.n648 B.n63 585
R76 B.n630 B.n62 585
R77 B.n649 B.n62 585
R78 B.n629 B.n628 585
R79 B.n628 B.n61 585
R80 B.n627 B.n57 585
R81 B.n655 B.n57 585
R82 B.n626 B.n56 585
R83 B.n656 B.n56 585
R84 B.n625 B.n55 585
R85 B.n657 B.n55 585
R86 B.n624 B.n623 585
R87 B.n623 B.n51 585
R88 B.n622 B.n50 585
R89 B.n663 B.n50 585
R90 B.n621 B.n49 585
R91 B.n664 B.n49 585
R92 B.n620 B.n48 585
R93 B.n665 B.n48 585
R94 B.n619 B.n618 585
R95 B.n618 B.n44 585
R96 B.n617 B.n43 585
R97 B.n671 B.n43 585
R98 B.n616 B.n42 585
R99 B.n672 B.n42 585
R100 B.n615 B.n41 585
R101 B.n673 B.n41 585
R102 B.n614 B.n613 585
R103 B.n613 B.n37 585
R104 B.n612 B.n36 585
R105 B.n679 B.n36 585
R106 B.n611 B.n35 585
R107 B.n680 B.n35 585
R108 B.n610 B.n34 585
R109 B.n681 B.n34 585
R110 B.n609 B.n608 585
R111 B.n608 B.n30 585
R112 B.n607 B.n29 585
R113 B.n687 B.n29 585
R114 B.n606 B.n28 585
R115 B.n688 B.n28 585
R116 B.n605 B.n27 585
R117 B.n689 B.n27 585
R118 B.n604 B.n603 585
R119 B.n603 B.n23 585
R120 B.n602 B.n22 585
R121 B.n695 B.n22 585
R122 B.n601 B.n21 585
R123 B.n696 B.n21 585
R124 B.n600 B.n20 585
R125 B.n697 B.n20 585
R126 B.n599 B.n598 585
R127 B.n598 B.n16 585
R128 B.n597 B.n15 585
R129 B.n703 B.n15 585
R130 B.n596 B.n14 585
R131 B.n704 B.n14 585
R132 B.n595 B.n13 585
R133 B.n705 B.n13 585
R134 B.n594 B.n593 585
R135 B.n593 B.n12 585
R136 B.n592 B.n591 585
R137 B.n592 B.n8 585
R138 B.n590 B.n7 585
R139 B.n712 B.n7 585
R140 B.n589 B.n6 585
R141 B.n713 B.n6 585
R142 B.n588 B.n5 585
R143 B.n714 B.n5 585
R144 B.n587 B.n586 585
R145 B.n586 B.n4 585
R146 B.n585 B.n237 585
R147 B.n585 B.n584 585
R148 B.n575 B.n238 585
R149 B.n239 B.n238 585
R150 B.n577 B.n576 585
R151 B.n578 B.n577 585
R152 B.n574 B.n243 585
R153 B.n247 B.n243 585
R154 B.n573 B.n572 585
R155 B.n572 B.n571 585
R156 B.n245 B.n244 585
R157 B.n246 B.n245 585
R158 B.n564 B.n563 585
R159 B.n565 B.n564 585
R160 B.n562 B.n252 585
R161 B.n252 B.n251 585
R162 B.n561 B.n560 585
R163 B.n560 B.n559 585
R164 B.n254 B.n253 585
R165 B.n255 B.n254 585
R166 B.n552 B.n551 585
R167 B.n553 B.n552 585
R168 B.n550 B.n260 585
R169 B.n260 B.n259 585
R170 B.n549 B.n548 585
R171 B.n548 B.n547 585
R172 B.n262 B.n261 585
R173 B.n263 B.n262 585
R174 B.n540 B.n539 585
R175 B.n541 B.n540 585
R176 B.n538 B.n268 585
R177 B.n268 B.n267 585
R178 B.n537 B.n536 585
R179 B.n536 B.n535 585
R180 B.n270 B.n269 585
R181 B.n271 B.n270 585
R182 B.n528 B.n527 585
R183 B.n529 B.n528 585
R184 B.n526 B.n276 585
R185 B.n276 B.n275 585
R186 B.n525 B.n524 585
R187 B.n524 B.n523 585
R188 B.n278 B.n277 585
R189 B.n279 B.n278 585
R190 B.n516 B.n515 585
R191 B.n517 B.n516 585
R192 B.n514 B.n284 585
R193 B.n284 B.n283 585
R194 B.n513 B.n512 585
R195 B.n512 B.n511 585
R196 B.n286 B.n285 585
R197 B.n287 B.n286 585
R198 B.n504 B.n503 585
R199 B.n505 B.n504 585
R200 B.n502 B.n292 585
R201 B.n292 B.n291 585
R202 B.n501 B.n500 585
R203 B.n500 B.n499 585
R204 B.n294 B.n293 585
R205 B.n492 B.n294 585
R206 B.n491 B.n490 585
R207 B.n493 B.n491 585
R208 B.n489 B.n299 585
R209 B.n299 B.n298 585
R210 B.n488 B.n487 585
R211 B.n487 B.n486 585
R212 B.n301 B.n300 585
R213 B.n302 B.n301 585
R214 B.n479 B.n478 585
R215 B.n480 B.n479 585
R216 B.n477 B.n307 585
R217 B.n307 B.n306 585
R218 B.n471 B.n470 585
R219 B.n469 B.n341 585
R220 B.n468 B.n340 585
R221 B.n473 B.n340 585
R222 B.n467 B.n466 585
R223 B.n465 B.n464 585
R224 B.n463 B.n462 585
R225 B.n461 B.n460 585
R226 B.n459 B.n458 585
R227 B.n457 B.n456 585
R228 B.n455 B.n454 585
R229 B.n453 B.n452 585
R230 B.n451 B.n450 585
R231 B.n449 B.n448 585
R232 B.n447 B.n446 585
R233 B.n445 B.n444 585
R234 B.n443 B.n442 585
R235 B.n441 B.n440 585
R236 B.n439 B.n438 585
R237 B.n437 B.n436 585
R238 B.n435 B.n434 585
R239 B.n433 B.n432 585
R240 B.n431 B.n430 585
R241 B.n429 B.n428 585
R242 B.n427 B.n426 585
R243 B.n425 B.n424 585
R244 B.n423 B.n422 585
R245 B.n421 B.n420 585
R246 B.n419 B.n418 585
R247 B.n416 B.n415 585
R248 B.n414 B.n413 585
R249 B.n412 B.n411 585
R250 B.n410 B.n409 585
R251 B.n408 B.n407 585
R252 B.n406 B.n405 585
R253 B.n404 B.n403 585
R254 B.n402 B.n401 585
R255 B.n400 B.n399 585
R256 B.n398 B.n397 585
R257 B.n396 B.n395 585
R258 B.n394 B.n393 585
R259 B.n392 B.n391 585
R260 B.n390 B.n389 585
R261 B.n388 B.n387 585
R262 B.n386 B.n385 585
R263 B.n384 B.n383 585
R264 B.n382 B.n381 585
R265 B.n380 B.n379 585
R266 B.n378 B.n377 585
R267 B.n376 B.n375 585
R268 B.n374 B.n373 585
R269 B.n372 B.n371 585
R270 B.n370 B.n369 585
R271 B.n368 B.n367 585
R272 B.n366 B.n365 585
R273 B.n364 B.n363 585
R274 B.n362 B.n361 585
R275 B.n360 B.n359 585
R276 B.n358 B.n357 585
R277 B.n356 B.n355 585
R278 B.n354 B.n353 585
R279 B.n352 B.n351 585
R280 B.n350 B.n349 585
R281 B.n348 B.n347 585
R282 B.n309 B.n308 585
R283 B.n476 B.n475 585
R284 B.n305 B.n304 585
R285 B.n306 B.n305 585
R286 B.n482 B.n481 585
R287 B.n481 B.n480 585
R288 B.n483 B.n303 585
R289 B.n303 B.n302 585
R290 B.n485 B.n484 585
R291 B.n486 B.n485 585
R292 B.n297 B.n296 585
R293 B.n298 B.n297 585
R294 B.n495 B.n494 585
R295 B.n494 B.n493 585
R296 B.n496 B.n295 585
R297 B.n492 B.n295 585
R298 B.n498 B.n497 585
R299 B.n499 B.n498 585
R300 B.n290 B.n289 585
R301 B.n291 B.n290 585
R302 B.n507 B.n506 585
R303 B.n506 B.n505 585
R304 B.n508 B.n288 585
R305 B.n288 B.n287 585
R306 B.n510 B.n509 585
R307 B.n511 B.n510 585
R308 B.n282 B.n281 585
R309 B.n283 B.n282 585
R310 B.n519 B.n518 585
R311 B.n518 B.n517 585
R312 B.n520 B.n280 585
R313 B.n280 B.n279 585
R314 B.n522 B.n521 585
R315 B.n523 B.n522 585
R316 B.n274 B.n273 585
R317 B.n275 B.n274 585
R318 B.n531 B.n530 585
R319 B.n530 B.n529 585
R320 B.n532 B.n272 585
R321 B.n272 B.n271 585
R322 B.n534 B.n533 585
R323 B.n535 B.n534 585
R324 B.n266 B.n265 585
R325 B.n267 B.n266 585
R326 B.n543 B.n542 585
R327 B.n542 B.n541 585
R328 B.n544 B.n264 585
R329 B.n264 B.n263 585
R330 B.n546 B.n545 585
R331 B.n547 B.n546 585
R332 B.n258 B.n257 585
R333 B.n259 B.n258 585
R334 B.n555 B.n554 585
R335 B.n554 B.n553 585
R336 B.n556 B.n256 585
R337 B.n256 B.n255 585
R338 B.n558 B.n557 585
R339 B.n559 B.n558 585
R340 B.n250 B.n249 585
R341 B.n251 B.n250 585
R342 B.n567 B.n566 585
R343 B.n566 B.n565 585
R344 B.n568 B.n248 585
R345 B.n248 B.n246 585
R346 B.n570 B.n569 585
R347 B.n571 B.n570 585
R348 B.n242 B.n241 585
R349 B.n247 B.n242 585
R350 B.n580 B.n579 585
R351 B.n579 B.n578 585
R352 B.n581 B.n240 585
R353 B.n240 B.n239 585
R354 B.n583 B.n582 585
R355 B.n584 B.n583 585
R356 B.n3 B.n0 585
R357 B.n4 B.n3 585
R358 B.n711 B.n1 585
R359 B.n712 B.n711 585
R360 B.n710 B.n709 585
R361 B.n710 B.n8 585
R362 B.n708 B.n9 585
R363 B.n12 B.n9 585
R364 B.n707 B.n706 585
R365 B.n706 B.n705 585
R366 B.n11 B.n10 585
R367 B.n704 B.n11 585
R368 B.n702 B.n701 585
R369 B.n703 B.n702 585
R370 B.n700 B.n17 585
R371 B.n17 B.n16 585
R372 B.n699 B.n698 585
R373 B.n698 B.n697 585
R374 B.n19 B.n18 585
R375 B.n696 B.n19 585
R376 B.n694 B.n693 585
R377 B.n695 B.n694 585
R378 B.n692 B.n24 585
R379 B.n24 B.n23 585
R380 B.n691 B.n690 585
R381 B.n690 B.n689 585
R382 B.n26 B.n25 585
R383 B.n688 B.n26 585
R384 B.n686 B.n685 585
R385 B.n687 B.n686 585
R386 B.n684 B.n31 585
R387 B.n31 B.n30 585
R388 B.n683 B.n682 585
R389 B.n682 B.n681 585
R390 B.n33 B.n32 585
R391 B.n680 B.n33 585
R392 B.n678 B.n677 585
R393 B.n679 B.n678 585
R394 B.n676 B.n38 585
R395 B.n38 B.n37 585
R396 B.n675 B.n674 585
R397 B.n674 B.n673 585
R398 B.n40 B.n39 585
R399 B.n672 B.n40 585
R400 B.n670 B.n669 585
R401 B.n671 B.n670 585
R402 B.n668 B.n45 585
R403 B.n45 B.n44 585
R404 B.n667 B.n666 585
R405 B.n666 B.n665 585
R406 B.n47 B.n46 585
R407 B.n664 B.n47 585
R408 B.n662 B.n661 585
R409 B.n663 B.n662 585
R410 B.n660 B.n52 585
R411 B.n52 B.n51 585
R412 B.n659 B.n658 585
R413 B.n658 B.n657 585
R414 B.n54 B.n53 585
R415 B.n656 B.n54 585
R416 B.n654 B.n653 585
R417 B.n655 B.n654 585
R418 B.n652 B.n58 585
R419 B.n61 B.n58 585
R420 B.n651 B.n650 585
R421 B.n650 B.n649 585
R422 B.n60 B.n59 585
R423 B.n648 B.n60 585
R424 B.n646 B.n645 585
R425 B.n647 B.n646 585
R426 B.n644 B.n66 585
R427 B.n66 B.n65 585
R428 B.n643 B.n642 585
R429 B.n642 B.n641 585
R430 B.n68 B.n67 585
R431 B.n640 B.n68 585
R432 B.n715 B.n714 585
R433 B.n713 B.n2 585
R434 B.n109 B.n68 516.524
R435 B.n638 B.n70 516.524
R436 B.n475 B.n307 516.524
R437 B.n471 B.n305 516.524
R438 B.n106 B.t8 310.055
R439 B.n104 B.t16 310.055
R440 B.n344 B.t19 310.055
R441 B.n342 B.t12 310.055
R442 B.n639 B.n102 256.663
R443 B.n639 B.n101 256.663
R444 B.n639 B.n100 256.663
R445 B.n639 B.n99 256.663
R446 B.n639 B.n98 256.663
R447 B.n639 B.n97 256.663
R448 B.n639 B.n96 256.663
R449 B.n639 B.n95 256.663
R450 B.n639 B.n94 256.663
R451 B.n639 B.n93 256.663
R452 B.n639 B.n92 256.663
R453 B.n639 B.n91 256.663
R454 B.n639 B.n90 256.663
R455 B.n639 B.n89 256.663
R456 B.n639 B.n88 256.663
R457 B.n639 B.n87 256.663
R458 B.n639 B.n86 256.663
R459 B.n639 B.n85 256.663
R460 B.n639 B.n84 256.663
R461 B.n639 B.n83 256.663
R462 B.n639 B.n82 256.663
R463 B.n639 B.n81 256.663
R464 B.n639 B.n80 256.663
R465 B.n639 B.n79 256.663
R466 B.n639 B.n78 256.663
R467 B.n639 B.n77 256.663
R468 B.n639 B.n76 256.663
R469 B.n639 B.n75 256.663
R470 B.n639 B.n74 256.663
R471 B.n639 B.n73 256.663
R472 B.n639 B.n72 256.663
R473 B.n639 B.n71 256.663
R474 B.n473 B.n472 256.663
R475 B.n473 B.n310 256.663
R476 B.n473 B.n311 256.663
R477 B.n473 B.n312 256.663
R478 B.n473 B.n313 256.663
R479 B.n473 B.n314 256.663
R480 B.n473 B.n315 256.663
R481 B.n473 B.n316 256.663
R482 B.n473 B.n317 256.663
R483 B.n473 B.n318 256.663
R484 B.n473 B.n319 256.663
R485 B.n473 B.n320 256.663
R486 B.n473 B.n321 256.663
R487 B.n473 B.n322 256.663
R488 B.n473 B.n323 256.663
R489 B.n473 B.n324 256.663
R490 B.n473 B.n325 256.663
R491 B.n473 B.n326 256.663
R492 B.n473 B.n327 256.663
R493 B.n473 B.n328 256.663
R494 B.n473 B.n329 256.663
R495 B.n473 B.n330 256.663
R496 B.n473 B.n331 256.663
R497 B.n473 B.n332 256.663
R498 B.n473 B.n333 256.663
R499 B.n473 B.n334 256.663
R500 B.n473 B.n335 256.663
R501 B.n473 B.n336 256.663
R502 B.n473 B.n337 256.663
R503 B.n473 B.n338 256.663
R504 B.n473 B.n339 256.663
R505 B.n474 B.n473 256.663
R506 B.n717 B.n716 256.663
R507 B.n104 B.t17 239.21
R508 B.n344 B.t21 239.21
R509 B.n106 B.t10 239.21
R510 B.n342 B.t15 239.21
R511 B.n105 B.t18 200.228
R512 B.n345 B.t20 200.228
R513 B.n107 B.t11 200.228
R514 B.n343 B.t14 200.228
R515 B.n113 B.n112 163.367
R516 B.n117 B.n116 163.367
R517 B.n121 B.n120 163.367
R518 B.n125 B.n124 163.367
R519 B.n129 B.n128 163.367
R520 B.n133 B.n132 163.367
R521 B.n137 B.n136 163.367
R522 B.n141 B.n140 163.367
R523 B.n145 B.n144 163.367
R524 B.n149 B.n148 163.367
R525 B.n153 B.n152 163.367
R526 B.n157 B.n156 163.367
R527 B.n161 B.n160 163.367
R528 B.n165 B.n164 163.367
R529 B.n169 B.n168 163.367
R530 B.n173 B.n172 163.367
R531 B.n177 B.n176 163.367
R532 B.n181 B.n180 163.367
R533 B.n186 B.n185 163.367
R534 B.n190 B.n189 163.367
R535 B.n194 B.n193 163.367
R536 B.n198 B.n197 163.367
R537 B.n202 B.n201 163.367
R538 B.n206 B.n205 163.367
R539 B.n210 B.n209 163.367
R540 B.n214 B.n213 163.367
R541 B.n218 B.n217 163.367
R542 B.n222 B.n221 163.367
R543 B.n226 B.n225 163.367
R544 B.n230 B.n229 163.367
R545 B.n234 B.n233 163.367
R546 B.n638 B.n103 163.367
R547 B.n479 B.n307 163.367
R548 B.n479 B.n301 163.367
R549 B.n487 B.n301 163.367
R550 B.n487 B.n299 163.367
R551 B.n491 B.n299 163.367
R552 B.n491 B.n294 163.367
R553 B.n500 B.n294 163.367
R554 B.n500 B.n292 163.367
R555 B.n504 B.n292 163.367
R556 B.n504 B.n286 163.367
R557 B.n512 B.n286 163.367
R558 B.n512 B.n284 163.367
R559 B.n516 B.n284 163.367
R560 B.n516 B.n278 163.367
R561 B.n524 B.n278 163.367
R562 B.n524 B.n276 163.367
R563 B.n528 B.n276 163.367
R564 B.n528 B.n270 163.367
R565 B.n536 B.n270 163.367
R566 B.n536 B.n268 163.367
R567 B.n540 B.n268 163.367
R568 B.n540 B.n262 163.367
R569 B.n548 B.n262 163.367
R570 B.n548 B.n260 163.367
R571 B.n552 B.n260 163.367
R572 B.n552 B.n254 163.367
R573 B.n560 B.n254 163.367
R574 B.n560 B.n252 163.367
R575 B.n564 B.n252 163.367
R576 B.n564 B.n245 163.367
R577 B.n572 B.n245 163.367
R578 B.n572 B.n243 163.367
R579 B.n577 B.n243 163.367
R580 B.n577 B.n238 163.367
R581 B.n585 B.n238 163.367
R582 B.n586 B.n585 163.367
R583 B.n586 B.n5 163.367
R584 B.n6 B.n5 163.367
R585 B.n7 B.n6 163.367
R586 B.n592 B.n7 163.367
R587 B.n593 B.n592 163.367
R588 B.n593 B.n13 163.367
R589 B.n14 B.n13 163.367
R590 B.n15 B.n14 163.367
R591 B.n598 B.n15 163.367
R592 B.n598 B.n20 163.367
R593 B.n21 B.n20 163.367
R594 B.n22 B.n21 163.367
R595 B.n603 B.n22 163.367
R596 B.n603 B.n27 163.367
R597 B.n28 B.n27 163.367
R598 B.n29 B.n28 163.367
R599 B.n608 B.n29 163.367
R600 B.n608 B.n34 163.367
R601 B.n35 B.n34 163.367
R602 B.n36 B.n35 163.367
R603 B.n613 B.n36 163.367
R604 B.n613 B.n41 163.367
R605 B.n42 B.n41 163.367
R606 B.n43 B.n42 163.367
R607 B.n618 B.n43 163.367
R608 B.n618 B.n48 163.367
R609 B.n49 B.n48 163.367
R610 B.n50 B.n49 163.367
R611 B.n623 B.n50 163.367
R612 B.n623 B.n55 163.367
R613 B.n56 B.n55 163.367
R614 B.n57 B.n56 163.367
R615 B.n628 B.n57 163.367
R616 B.n628 B.n62 163.367
R617 B.n63 B.n62 163.367
R618 B.n64 B.n63 163.367
R619 B.n633 B.n64 163.367
R620 B.n633 B.n69 163.367
R621 B.n70 B.n69 163.367
R622 B.n341 B.n340 163.367
R623 B.n466 B.n340 163.367
R624 B.n464 B.n463 163.367
R625 B.n460 B.n459 163.367
R626 B.n456 B.n455 163.367
R627 B.n452 B.n451 163.367
R628 B.n448 B.n447 163.367
R629 B.n444 B.n443 163.367
R630 B.n440 B.n439 163.367
R631 B.n436 B.n435 163.367
R632 B.n432 B.n431 163.367
R633 B.n428 B.n427 163.367
R634 B.n424 B.n423 163.367
R635 B.n420 B.n419 163.367
R636 B.n415 B.n414 163.367
R637 B.n411 B.n410 163.367
R638 B.n407 B.n406 163.367
R639 B.n403 B.n402 163.367
R640 B.n399 B.n398 163.367
R641 B.n395 B.n394 163.367
R642 B.n391 B.n390 163.367
R643 B.n387 B.n386 163.367
R644 B.n383 B.n382 163.367
R645 B.n379 B.n378 163.367
R646 B.n375 B.n374 163.367
R647 B.n371 B.n370 163.367
R648 B.n367 B.n366 163.367
R649 B.n363 B.n362 163.367
R650 B.n359 B.n358 163.367
R651 B.n355 B.n354 163.367
R652 B.n351 B.n350 163.367
R653 B.n347 B.n309 163.367
R654 B.n481 B.n305 163.367
R655 B.n481 B.n303 163.367
R656 B.n485 B.n303 163.367
R657 B.n485 B.n297 163.367
R658 B.n494 B.n297 163.367
R659 B.n494 B.n295 163.367
R660 B.n498 B.n295 163.367
R661 B.n498 B.n290 163.367
R662 B.n506 B.n290 163.367
R663 B.n506 B.n288 163.367
R664 B.n510 B.n288 163.367
R665 B.n510 B.n282 163.367
R666 B.n518 B.n282 163.367
R667 B.n518 B.n280 163.367
R668 B.n522 B.n280 163.367
R669 B.n522 B.n274 163.367
R670 B.n530 B.n274 163.367
R671 B.n530 B.n272 163.367
R672 B.n534 B.n272 163.367
R673 B.n534 B.n266 163.367
R674 B.n542 B.n266 163.367
R675 B.n542 B.n264 163.367
R676 B.n546 B.n264 163.367
R677 B.n546 B.n258 163.367
R678 B.n554 B.n258 163.367
R679 B.n554 B.n256 163.367
R680 B.n558 B.n256 163.367
R681 B.n558 B.n250 163.367
R682 B.n566 B.n250 163.367
R683 B.n566 B.n248 163.367
R684 B.n570 B.n248 163.367
R685 B.n570 B.n242 163.367
R686 B.n579 B.n242 163.367
R687 B.n579 B.n240 163.367
R688 B.n583 B.n240 163.367
R689 B.n583 B.n3 163.367
R690 B.n715 B.n3 163.367
R691 B.n711 B.n2 163.367
R692 B.n711 B.n710 163.367
R693 B.n710 B.n9 163.367
R694 B.n706 B.n9 163.367
R695 B.n706 B.n11 163.367
R696 B.n702 B.n11 163.367
R697 B.n702 B.n17 163.367
R698 B.n698 B.n17 163.367
R699 B.n698 B.n19 163.367
R700 B.n694 B.n19 163.367
R701 B.n694 B.n24 163.367
R702 B.n690 B.n24 163.367
R703 B.n690 B.n26 163.367
R704 B.n686 B.n26 163.367
R705 B.n686 B.n31 163.367
R706 B.n682 B.n31 163.367
R707 B.n682 B.n33 163.367
R708 B.n678 B.n33 163.367
R709 B.n678 B.n38 163.367
R710 B.n674 B.n38 163.367
R711 B.n674 B.n40 163.367
R712 B.n670 B.n40 163.367
R713 B.n670 B.n45 163.367
R714 B.n666 B.n45 163.367
R715 B.n666 B.n47 163.367
R716 B.n662 B.n47 163.367
R717 B.n662 B.n52 163.367
R718 B.n658 B.n52 163.367
R719 B.n658 B.n54 163.367
R720 B.n654 B.n54 163.367
R721 B.n654 B.n58 163.367
R722 B.n650 B.n58 163.367
R723 B.n650 B.n60 163.367
R724 B.n646 B.n60 163.367
R725 B.n646 B.n66 163.367
R726 B.n642 B.n66 163.367
R727 B.n642 B.n68 163.367
R728 B.n473 B.n306 118.564
R729 B.n640 B.n639 118.564
R730 B.n109 B.n71 71.676
R731 B.n113 B.n72 71.676
R732 B.n117 B.n73 71.676
R733 B.n121 B.n74 71.676
R734 B.n125 B.n75 71.676
R735 B.n129 B.n76 71.676
R736 B.n133 B.n77 71.676
R737 B.n137 B.n78 71.676
R738 B.n141 B.n79 71.676
R739 B.n145 B.n80 71.676
R740 B.n149 B.n81 71.676
R741 B.n153 B.n82 71.676
R742 B.n157 B.n83 71.676
R743 B.n161 B.n84 71.676
R744 B.n165 B.n85 71.676
R745 B.n169 B.n86 71.676
R746 B.n173 B.n87 71.676
R747 B.n177 B.n88 71.676
R748 B.n181 B.n89 71.676
R749 B.n186 B.n90 71.676
R750 B.n190 B.n91 71.676
R751 B.n194 B.n92 71.676
R752 B.n198 B.n93 71.676
R753 B.n202 B.n94 71.676
R754 B.n206 B.n95 71.676
R755 B.n210 B.n96 71.676
R756 B.n214 B.n97 71.676
R757 B.n218 B.n98 71.676
R758 B.n222 B.n99 71.676
R759 B.n226 B.n100 71.676
R760 B.n230 B.n101 71.676
R761 B.n234 B.n102 71.676
R762 B.n103 B.n102 71.676
R763 B.n233 B.n101 71.676
R764 B.n229 B.n100 71.676
R765 B.n225 B.n99 71.676
R766 B.n221 B.n98 71.676
R767 B.n217 B.n97 71.676
R768 B.n213 B.n96 71.676
R769 B.n209 B.n95 71.676
R770 B.n205 B.n94 71.676
R771 B.n201 B.n93 71.676
R772 B.n197 B.n92 71.676
R773 B.n193 B.n91 71.676
R774 B.n189 B.n90 71.676
R775 B.n185 B.n89 71.676
R776 B.n180 B.n88 71.676
R777 B.n176 B.n87 71.676
R778 B.n172 B.n86 71.676
R779 B.n168 B.n85 71.676
R780 B.n164 B.n84 71.676
R781 B.n160 B.n83 71.676
R782 B.n156 B.n82 71.676
R783 B.n152 B.n81 71.676
R784 B.n148 B.n80 71.676
R785 B.n144 B.n79 71.676
R786 B.n140 B.n78 71.676
R787 B.n136 B.n77 71.676
R788 B.n132 B.n76 71.676
R789 B.n128 B.n75 71.676
R790 B.n124 B.n74 71.676
R791 B.n120 B.n73 71.676
R792 B.n116 B.n72 71.676
R793 B.n112 B.n71 71.676
R794 B.n472 B.n471 71.676
R795 B.n466 B.n310 71.676
R796 B.n463 B.n311 71.676
R797 B.n459 B.n312 71.676
R798 B.n455 B.n313 71.676
R799 B.n451 B.n314 71.676
R800 B.n447 B.n315 71.676
R801 B.n443 B.n316 71.676
R802 B.n439 B.n317 71.676
R803 B.n435 B.n318 71.676
R804 B.n431 B.n319 71.676
R805 B.n427 B.n320 71.676
R806 B.n423 B.n321 71.676
R807 B.n419 B.n322 71.676
R808 B.n414 B.n323 71.676
R809 B.n410 B.n324 71.676
R810 B.n406 B.n325 71.676
R811 B.n402 B.n326 71.676
R812 B.n398 B.n327 71.676
R813 B.n394 B.n328 71.676
R814 B.n390 B.n329 71.676
R815 B.n386 B.n330 71.676
R816 B.n382 B.n331 71.676
R817 B.n378 B.n332 71.676
R818 B.n374 B.n333 71.676
R819 B.n370 B.n334 71.676
R820 B.n366 B.n335 71.676
R821 B.n362 B.n336 71.676
R822 B.n358 B.n337 71.676
R823 B.n354 B.n338 71.676
R824 B.n350 B.n339 71.676
R825 B.n474 B.n309 71.676
R826 B.n472 B.n341 71.676
R827 B.n464 B.n310 71.676
R828 B.n460 B.n311 71.676
R829 B.n456 B.n312 71.676
R830 B.n452 B.n313 71.676
R831 B.n448 B.n314 71.676
R832 B.n444 B.n315 71.676
R833 B.n440 B.n316 71.676
R834 B.n436 B.n317 71.676
R835 B.n432 B.n318 71.676
R836 B.n428 B.n319 71.676
R837 B.n424 B.n320 71.676
R838 B.n420 B.n321 71.676
R839 B.n415 B.n322 71.676
R840 B.n411 B.n323 71.676
R841 B.n407 B.n324 71.676
R842 B.n403 B.n325 71.676
R843 B.n399 B.n326 71.676
R844 B.n395 B.n327 71.676
R845 B.n391 B.n328 71.676
R846 B.n387 B.n329 71.676
R847 B.n383 B.n330 71.676
R848 B.n379 B.n331 71.676
R849 B.n375 B.n332 71.676
R850 B.n371 B.n333 71.676
R851 B.n367 B.n334 71.676
R852 B.n363 B.n335 71.676
R853 B.n359 B.n336 71.676
R854 B.n355 B.n337 71.676
R855 B.n351 B.n338 71.676
R856 B.n347 B.n339 71.676
R857 B.n475 B.n474 71.676
R858 B.n716 B.n715 71.676
R859 B.n716 B.n2 71.676
R860 B.n480 B.n306 59.7211
R861 B.n480 B.n302 59.7211
R862 B.n486 B.n302 59.7211
R863 B.n486 B.n298 59.7211
R864 B.n493 B.n298 59.7211
R865 B.n493 B.n492 59.7211
R866 B.n499 B.n291 59.7211
R867 B.n505 B.n291 59.7211
R868 B.n505 B.n287 59.7211
R869 B.n511 B.n287 59.7211
R870 B.n511 B.n283 59.7211
R871 B.n517 B.n283 59.7211
R872 B.n517 B.n279 59.7211
R873 B.n523 B.n279 59.7211
R874 B.n529 B.n275 59.7211
R875 B.n529 B.n271 59.7211
R876 B.n535 B.n271 59.7211
R877 B.n535 B.n267 59.7211
R878 B.n541 B.n267 59.7211
R879 B.n547 B.n263 59.7211
R880 B.n547 B.n259 59.7211
R881 B.n553 B.n259 59.7211
R882 B.n553 B.n255 59.7211
R883 B.n559 B.n255 59.7211
R884 B.n565 B.n251 59.7211
R885 B.n565 B.n246 59.7211
R886 B.n571 B.n246 59.7211
R887 B.n571 B.n247 59.7211
R888 B.n578 B.n239 59.7211
R889 B.n584 B.n239 59.7211
R890 B.n584 B.n4 59.7211
R891 B.n714 B.n4 59.7211
R892 B.n714 B.n713 59.7211
R893 B.n713 B.n712 59.7211
R894 B.n712 B.n8 59.7211
R895 B.n12 B.n8 59.7211
R896 B.n705 B.n12 59.7211
R897 B.n704 B.n703 59.7211
R898 B.n703 B.n16 59.7211
R899 B.n697 B.n16 59.7211
R900 B.n697 B.n696 59.7211
R901 B.n695 B.n23 59.7211
R902 B.n689 B.n23 59.7211
R903 B.n689 B.n688 59.7211
R904 B.n688 B.n687 59.7211
R905 B.n687 B.n30 59.7211
R906 B.n681 B.n680 59.7211
R907 B.n680 B.n679 59.7211
R908 B.n679 B.n37 59.7211
R909 B.n673 B.n37 59.7211
R910 B.n673 B.n672 59.7211
R911 B.n671 B.n44 59.7211
R912 B.n665 B.n44 59.7211
R913 B.n665 B.n664 59.7211
R914 B.n664 B.n663 59.7211
R915 B.n663 B.n51 59.7211
R916 B.n657 B.n51 59.7211
R917 B.n657 B.n656 59.7211
R918 B.n656 B.n655 59.7211
R919 B.n649 B.n61 59.7211
R920 B.n649 B.n648 59.7211
R921 B.n648 B.n647 59.7211
R922 B.n647 B.n65 59.7211
R923 B.n641 B.n65 59.7211
R924 B.n641 B.n640 59.7211
R925 B.n108 B.n107 59.5399
R926 B.n183 B.n105 59.5399
R927 B.n346 B.n345 59.5399
R928 B.n417 B.n343 59.5399
R929 B.t6 B.n251 57.9646
R930 B.n696 B.t1 57.9646
R931 B.n247 B.t3 56.2081
R932 B.t7 B.n704 56.2081
R933 B.n499 B.t13 54.4516
R934 B.n655 B.t9 54.4516
R935 B.t2 B.n263 52.6951
R936 B.t0 B.n30 52.6951
R937 B.t4 B.n275 47.4256
R938 B.n672 B.t5 47.4256
R939 B.n107 B.n106 38.9823
R940 B.n105 B.n104 38.9823
R941 B.n345 B.n344 38.9823
R942 B.n343 B.n342 38.9823
R943 B.n470 B.n304 33.5615
R944 B.n477 B.n476 33.5615
R945 B.n637 B.n636 33.5615
R946 B.n110 B.n67 33.5615
R947 B B.n717 18.0485
R948 B.n523 B.t4 12.2959
R949 B.t5 B.n671 12.2959
R950 B.n482 B.n304 10.6151
R951 B.n483 B.n482 10.6151
R952 B.n484 B.n483 10.6151
R953 B.n484 B.n296 10.6151
R954 B.n495 B.n296 10.6151
R955 B.n496 B.n495 10.6151
R956 B.n497 B.n496 10.6151
R957 B.n497 B.n289 10.6151
R958 B.n507 B.n289 10.6151
R959 B.n508 B.n507 10.6151
R960 B.n509 B.n508 10.6151
R961 B.n509 B.n281 10.6151
R962 B.n519 B.n281 10.6151
R963 B.n520 B.n519 10.6151
R964 B.n521 B.n520 10.6151
R965 B.n521 B.n273 10.6151
R966 B.n531 B.n273 10.6151
R967 B.n532 B.n531 10.6151
R968 B.n533 B.n532 10.6151
R969 B.n533 B.n265 10.6151
R970 B.n543 B.n265 10.6151
R971 B.n544 B.n543 10.6151
R972 B.n545 B.n544 10.6151
R973 B.n545 B.n257 10.6151
R974 B.n555 B.n257 10.6151
R975 B.n556 B.n555 10.6151
R976 B.n557 B.n556 10.6151
R977 B.n557 B.n249 10.6151
R978 B.n567 B.n249 10.6151
R979 B.n568 B.n567 10.6151
R980 B.n569 B.n568 10.6151
R981 B.n569 B.n241 10.6151
R982 B.n580 B.n241 10.6151
R983 B.n581 B.n580 10.6151
R984 B.n582 B.n581 10.6151
R985 B.n582 B.n0 10.6151
R986 B.n470 B.n469 10.6151
R987 B.n469 B.n468 10.6151
R988 B.n468 B.n467 10.6151
R989 B.n467 B.n465 10.6151
R990 B.n465 B.n462 10.6151
R991 B.n462 B.n461 10.6151
R992 B.n461 B.n458 10.6151
R993 B.n458 B.n457 10.6151
R994 B.n457 B.n454 10.6151
R995 B.n454 B.n453 10.6151
R996 B.n453 B.n450 10.6151
R997 B.n450 B.n449 10.6151
R998 B.n449 B.n446 10.6151
R999 B.n446 B.n445 10.6151
R1000 B.n445 B.n442 10.6151
R1001 B.n442 B.n441 10.6151
R1002 B.n441 B.n438 10.6151
R1003 B.n438 B.n437 10.6151
R1004 B.n437 B.n434 10.6151
R1005 B.n434 B.n433 10.6151
R1006 B.n433 B.n430 10.6151
R1007 B.n430 B.n429 10.6151
R1008 B.n429 B.n426 10.6151
R1009 B.n426 B.n425 10.6151
R1010 B.n425 B.n422 10.6151
R1011 B.n422 B.n421 10.6151
R1012 B.n421 B.n418 10.6151
R1013 B.n416 B.n413 10.6151
R1014 B.n413 B.n412 10.6151
R1015 B.n412 B.n409 10.6151
R1016 B.n409 B.n408 10.6151
R1017 B.n408 B.n405 10.6151
R1018 B.n405 B.n404 10.6151
R1019 B.n404 B.n401 10.6151
R1020 B.n401 B.n400 10.6151
R1021 B.n397 B.n396 10.6151
R1022 B.n396 B.n393 10.6151
R1023 B.n393 B.n392 10.6151
R1024 B.n392 B.n389 10.6151
R1025 B.n389 B.n388 10.6151
R1026 B.n388 B.n385 10.6151
R1027 B.n385 B.n384 10.6151
R1028 B.n384 B.n381 10.6151
R1029 B.n381 B.n380 10.6151
R1030 B.n380 B.n377 10.6151
R1031 B.n377 B.n376 10.6151
R1032 B.n376 B.n373 10.6151
R1033 B.n373 B.n372 10.6151
R1034 B.n372 B.n369 10.6151
R1035 B.n369 B.n368 10.6151
R1036 B.n368 B.n365 10.6151
R1037 B.n365 B.n364 10.6151
R1038 B.n364 B.n361 10.6151
R1039 B.n361 B.n360 10.6151
R1040 B.n360 B.n357 10.6151
R1041 B.n357 B.n356 10.6151
R1042 B.n356 B.n353 10.6151
R1043 B.n353 B.n352 10.6151
R1044 B.n352 B.n349 10.6151
R1045 B.n349 B.n348 10.6151
R1046 B.n348 B.n308 10.6151
R1047 B.n476 B.n308 10.6151
R1048 B.n478 B.n477 10.6151
R1049 B.n478 B.n300 10.6151
R1050 B.n488 B.n300 10.6151
R1051 B.n489 B.n488 10.6151
R1052 B.n490 B.n489 10.6151
R1053 B.n490 B.n293 10.6151
R1054 B.n501 B.n293 10.6151
R1055 B.n502 B.n501 10.6151
R1056 B.n503 B.n502 10.6151
R1057 B.n503 B.n285 10.6151
R1058 B.n513 B.n285 10.6151
R1059 B.n514 B.n513 10.6151
R1060 B.n515 B.n514 10.6151
R1061 B.n515 B.n277 10.6151
R1062 B.n525 B.n277 10.6151
R1063 B.n526 B.n525 10.6151
R1064 B.n527 B.n526 10.6151
R1065 B.n527 B.n269 10.6151
R1066 B.n537 B.n269 10.6151
R1067 B.n538 B.n537 10.6151
R1068 B.n539 B.n538 10.6151
R1069 B.n539 B.n261 10.6151
R1070 B.n549 B.n261 10.6151
R1071 B.n550 B.n549 10.6151
R1072 B.n551 B.n550 10.6151
R1073 B.n551 B.n253 10.6151
R1074 B.n561 B.n253 10.6151
R1075 B.n562 B.n561 10.6151
R1076 B.n563 B.n562 10.6151
R1077 B.n563 B.n244 10.6151
R1078 B.n573 B.n244 10.6151
R1079 B.n574 B.n573 10.6151
R1080 B.n576 B.n574 10.6151
R1081 B.n576 B.n575 10.6151
R1082 B.n575 B.n237 10.6151
R1083 B.n587 B.n237 10.6151
R1084 B.n588 B.n587 10.6151
R1085 B.n589 B.n588 10.6151
R1086 B.n590 B.n589 10.6151
R1087 B.n591 B.n590 10.6151
R1088 B.n594 B.n591 10.6151
R1089 B.n595 B.n594 10.6151
R1090 B.n596 B.n595 10.6151
R1091 B.n597 B.n596 10.6151
R1092 B.n599 B.n597 10.6151
R1093 B.n600 B.n599 10.6151
R1094 B.n601 B.n600 10.6151
R1095 B.n602 B.n601 10.6151
R1096 B.n604 B.n602 10.6151
R1097 B.n605 B.n604 10.6151
R1098 B.n606 B.n605 10.6151
R1099 B.n607 B.n606 10.6151
R1100 B.n609 B.n607 10.6151
R1101 B.n610 B.n609 10.6151
R1102 B.n611 B.n610 10.6151
R1103 B.n612 B.n611 10.6151
R1104 B.n614 B.n612 10.6151
R1105 B.n615 B.n614 10.6151
R1106 B.n616 B.n615 10.6151
R1107 B.n617 B.n616 10.6151
R1108 B.n619 B.n617 10.6151
R1109 B.n620 B.n619 10.6151
R1110 B.n621 B.n620 10.6151
R1111 B.n622 B.n621 10.6151
R1112 B.n624 B.n622 10.6151
R1113 B.n625 B.n624 10.6151
R1114 B.n626 B.n625 10.6151
R1115 B.n627 B.n626 10.6151
R1116 B.n629 B.n627 10.6151
R1117 B.n630 B.n629 10.6151
R1118 B.n631 B.n630 10.6151
R1119 B.n632 B.n631 10.6151
R1120 B.n634 B.n632 10.6151
R1121 B.n635 B.n634 10.6151
R1122 B.n636 B.n635 10.6151
R1123 B.n709 B.n1 10.6151
R1124 B.n709 B.n708 10.6151
R1125 B.n708 B.n707 10.6151
R1126 B.n707 B.n10 10.6151
R1127 B.n701 B.n10 10.6151
R1128 B.n701 B.n700 10.6151
R1129 B.n700 B.n699 10.6151
R1130 B.n699 B.n18 10.6151
R1131 B.n693 B.n18 10.6151
R1132 B.n693 B.n692 10.6151
R1133 B.n692 B.n691 10.6151
R1134 B.n691 B.n25 10.6151
R1135 B.n685 B.n25 10.6151
R1136 B.n685 B.n684 10.6151
R1137 B.n684 B.n683 10.6151
R1138 B.n683 B.n32 10.6151
R1139 B.n677 B.n32 10.6151
R1140 B.n677 B.n676 10.6151
R1141 B.n676 B.n675 10.6151
R1142 B.n675 B.n39 10.6151
R1143 B.n669 B.n39 10.6151
R1144 B.n669 B.n668 10.6151
R1145 B.n668 B.n667 10.6151
R1146 B.n667 B.n46 10.6151
R1147 B.n661 B.n46 10.6151
R1148 B.n661 B.n660 10.6151
R1149 B.n660 B.n659 10.6151
R1150 B.n659 B.n53 10.6151
R1151 B.n653 B.n53 10.6151
R1152 B.n653 B.n652 10.6151
R1153 B.n652 B.n651 10.6151
R1154 B.n651 B.n59 10.6151
R1155 B.n645 B.n59 10.6151
R1156 B.n645 B.n644 10.6151
R1157 B.n644 B.n643 10.6151
R1158 B.n643 B.n67 10.6151
R1159 B.n111 B.n110 10.6151
R1160 B.n114 B.n111 10.6151
R1161 B.n115 B.n114 10.6151
R1162 B.n118 B.n115 10.6151
R1163 B.n119 B.n118 10.6151
R1164 B.n122 B.n119 10.6151
R1165 B.n123 B.n122 10.6151
R1166 B.n126 B.n123 10.6151
R1167 B.n127 B.n126 10.6151
R1168 B.n130 B.n127 10.6151
R1169 B.n131 B.n130 10.6151
R1170 B.n134 B.n131 10.6151
R1171 B.n135 B.n134 10.6151
R1172 B.n138 B.n135 10.6151
R1173 B.n139 B.n138 10.6151
R1174 B.n142 B.n139 10.6151
R1175 B.n143 B.n142 10.6151
R1176 B.n146 B.n143 10.6151
R1177 B.n147 B.n146 10.6151
R1178 B.n150 B.n147 10.6151
R1179 B.n151 B.n150 10.6151
R1180 B.n154 B.n151 10.6151
R1181 B.n155 B.n154 10.6151
R1182 B.n158 B.n155 10.6151
R1183 B.n159 B.n158 10.6151
R1184 B.n162 B.n159 10.6151
R1185 B.n163 B.n162 10.6151
R1186 B.n167 B.n166 10.6151
R1187 B.n170 B.n167 10.6151
R1188 B.n171 B.n170 10.6151
R1189 B.n174 B.n171 10.6151
R1190 B.n175 B.n174 10.6151
R1191 B.n178 B.n175 10.6151
R1192 B.n179 B.n178 10.6151
R1193 B.n182 B.n179 10.6151
R1194 B.n187 B.n184 10.6151
R1195 B.n188 B.n187 10.6151
R1196 B.n191 B.n188 10.6151
R1197 B.n192 B.n191 10.6151
R1198 B.n195 B.n192 10.6151
R1199 B.n196 B.n195 10.6151
R1200 B.n199 B.n196 10.6151
R1201 B.n200 B.n199 10.6151
R1202 B.n203 B.n200 10.6151
R1203 B.n204 B.n203 10.6151
R1204 B.n207 B.n204 10.6151
R1205 B.n208 B.n207 10.6151
R1206 B.n211 B.n208 10.6151
R1207 B.n212 B.n211 10.6151
R1208 B.n215 B.n212 10.6151
R1209 B.n216 B.n215 10.6151
R1210 B.n219 B.n216 10.6151
R1211 B.n220 B.n219 10.6151
R1212 B.n223 B.n220 10.6151
R1213 B.n224 B.n223 10.6151
R1214 B.n227 B.n224 10.6151
R1215 B.n228 B.n227 10.6151
R1216 B.n231 B.n228 10.6151
R1217 B.n232 B.n231 10.6151
R1218 B.n235 B.n232 10.6151
R1219 B.n236 B.n235 10.6151
R1220 B.n637 B.n236 10.6151
R1221 B.n717 B.n0 8.11757
R1222 B.n717 B.n1 8.11757
R1223 B.n541 B.t2 7.02645
R1224 B.n681 B.t0 7.02645
R1225 B.n417 B.n416 6.5566
R1226 B.n400 B.n346 6.5566
R1227 B.n166 B.n108 6.5566
R1228 B.n183 B.n182 6.5566
R1229 B.n492 B.t13 5.26996
R1230 B.n61 B.t9 5.26996
R1231 B.n418 B.n417 4.05904
R1232 B.n397 B.n346 4.05904
R1233 B.n163 B.n108 4.05904
R1234 B.n184 B.n183 4.05904
R1235 B.n578 B.t3 3.51347
R1236 B.n705 B.t7 3.51347
R1237 B.n559 B.t6 1.75699
R1238 B.t1 B.n695 1.75699
R1239 VP.n31 VP.n30 185.034
R1240 VP.n54 VP.n53 185.034
R1241 VP.n29 VP.n28 185.034
R1242 VP.n14 VP.n11 161.3
R1243 VP.n16 VP.n15 161.3
R1244 VP.n17 VP.n10 161.3
R1245 VP.n19 VP.n18 161.3
R1246 VP.n20 VP.n9 161.3
R1247 VP.n23 VP.n22 161.3
R1248 VP.n24 VP.n8 161.3
R1249 VP.n26 VP.n25 161.3
R1250 VP.n27 VP.n7 161.3
R1251 VP.n52 VP.n0 161.3
R1252 VP.n51 VP.n50 161.3
R1253 VP.n49 VP.n1 161.3
R1254 VP.n48 VP.n47 161.3
R1255 VP.n45 VP.n2 161.3
R1256 VP.n44 VP.n43 161.3
R1257 VP.n42 VP.n3 161.3
R1258 VP.n41 VP.n40 161.3
R1259 VP.n39 VP.n4 161.3
R1260 VP.n37 VP.n36 161.3
R1261 VP.n35 VP.n5 161.3
R1262 VP.n34 VP.n33 161.3
R1263 VP.n32 VP.n6 161.3
R1264 VP.n12 VP.t7 131.504
R1265 VP.n31 VP.t0 104.004
R1266 VP.n38 VP.t5 104.004
R1267 VP.n46 VP.t4 104.004
R1268 VP.n53 VP.t3 104.004
R1269 VP.n28 VP.t6 104.004
R1270 VP.n21 VP.t2 104.004
R1271 VP.n13 VP.t1 104.004
R1272 VP.n13 VP.n12 68.7155
R1273 VP.n30 VP.n29 42.8187
R1274 VP.n33 VP.n5 41.4647
R1275 VP.n51 VP.n1 41.4647
R1276 VP.n26 VP.n8 41.4647
R1277 VP.n40 VP.n3 40.4934
R1278 VP.n44 VP.n3 40.4934
R1279 VP.n19 VP.n10 40.4934
R1280 VP.n15 VP.n10 40.4934
R1281 VP.n37 VP.n5 39.5221
R1282 VP.n47 VP.n1 39.5221
R1283 VP.n22 VP.n8 39.5221
R1284 VP.n33 VP.n32 24.4675
R1285 VP.n40 VP.n39 24.4675
R1286 VP.n45 VP.n44 24.4675
R1287 VP.n52 VP.n51 24.4675
R1288 VP.n27 VP.n26 24.4675
R1289 VP.n20 VP.n19 24.4675
R1290 VP.n15 VP.n14 24.4675
R1291 VP.n38 VP.n37 24.2228
R1292 VP.n47 VP.n46 24.2228
R1293 VP.n22 VP.n21 24.2228
R1294 VP.n12 VP.n11 18.9997
R1295 VP.n32 VP.n31 0.73451
R1296 VP.n53 VP.n52 0.73451
R1297 VP.n28 VP.n27 0.73451
R1298 VP.n39 VP.n38 0.24517
R1299 VP.n46 VP.n45 0.24517
R1300 VP.n21 VP.n20 0.24517
R1301 VP.n14 VP.n13 0.24517
R1302 VP.n16 VP.n11 0.189894
R1303 VP.n17 VP.n16 0.189894
R1304 VP.n18 VP.n17 0.189894
R1305 VP.n18 VP.n9 0.189894
R1306 VP.n23 VP.n9 0.189894
R1307 VP.n24 VP.n23 0.189894
R1308 VP.n25 VP.n24 0.189894
R1309 VP.n25 VP.n7 0.189894
R1310 VP.n29 VP.n7 0.189894
R1311 VP.n30 VP.n6 0.189894
R1312 VP.n34 VP.n6 0.189894
R1313 VP.n35 VP.n34 0.189894
R1314 VP.n36 VP.n35 0.189894
R1315 VP.n36 VP.n4 0.189894
R1316 VP.n41 VP.n4 0.189894
R1317 VP.n42 VP.n41 0.189894
R1318 VP.n43 VP.n42 0.189894
R1319 VP.n43 VP.n2 0.189894
R1320 VP.n48 VP.n2 0.189894
R1321 VP.n49 VP.n48 0.189894
R1322 VP.n50 VP.n49 0.189894
R1323 VP.n50 VP.n0 0.189894
R1324 VP.n54 VP.n0 0.189894
R1325 VP VP.n54 0.0516364
R1326 VDD1 VDD1.n0 68.8564
R1327 VDD1.n3 VDD1.n2 68.7428
R1328 VDD1.n3 VDD1.n1 68.7428
R1329 VDD1.n5 VDD1.n4 67.9318
R1330 VDD1.n5 VDD1.n3 38.3457
R1331 VDD1.n4 VDD1.t0 2.73153
R1332 VDD1.n4 VDD1.t3 2.73153
R1333 VDD1.n0 VDD1.t5 2.73153
R1334 VDD1.n0 VDD1.t6 2.73153
R1335 VDD1.n2 VDD1.t7 2.73153
R1336 VDD1.n2 VDD1.t2 2.73153
R1337 VDD1.n1 VDD1.t1 2.73153
R1338 VDD1.n1 VDD1.t4 2.73153
R1339 VDD1 VDD1.n5 0.80869
R1340 VTAIL.n290 VTAIL.n260 214.453
R1341 VTAIL.n32 VTAIL.n2 214.453
R1342 VTAIL.n68 VTAIL.n38 214.453
R1343 VTAIL.n106 VTAIL.n76 214.453
R1344 VTAIL.n254 VTAIL.n224 214.453
R1345 VTAIL.n216 VTAIL.n186 214.453
R1346 VTAIL.n180 VTAIL.n150 214.453
R1347 VTAIL.n142 VTAIL.n112 214.453
R1348 VTAIL.n273 VTAIL.n272 185
R1349 VTAIL.n275 VTAIL.n274 185
R1350 VTAIL.n268 VTAIL.n267 185
R1351 VTAIL.n281 VTAIL.n280 185
R1352 VTAIL.n283 VTAIL.n282 185
R1353 VTAIL.n264 VTAIL.n263 185
R1354 VTAIL.n289 VTAIL.n288 185
R1355 VTAIL.n291 VTAIL.n290 185
R1356 VTAIL.n15 VTAIL.n14 185
R1357 VTAIL.n17 VTAIL.n16 185
R1358 VTAIL.n10 VTAIL.n9 185
R1359 VTAIL.n23 VTAIL.n22 185
R1360 VTAIL.n25 VTAIL.n24 185
R1361 VTAIL.n6 VTAIL.n5 185
R1362 VTAIL.n31 VTAIL.n30 185
R1363 VTAIL.n33 VTAIL.n32 185
R1364 VTAIL.n51 VTAIL.n50 185
R1365 VTAIL.n53 VTAIL.n52 185
R1366 VTAIL.n46 VTAIL.n45 185
R1367 VTAIL.n59 VTAIL.n58 185
R1368 VTAIL.n61 VTAIL.n60 185
R1369 VTAIL.n42 VTAIL.n41 185
R1370 VTAIL.n67 VTAIL.n66 185
R1371 VTAIL.n69 VTAIL.n68 185
R1372 VTAIL.n89 VTAIL.n88 185
R1373 VTAIL.n91 VTAIL.n90 185
R1374 VTAIL.n84 VTAIL.n83 185
R1375 VTAIL.n97 VTAIL.n96 185
R1376 VTAIL.n99 VTAIL.n98 185
R1377 VTAIL.n80 VTAIL.n79 185
R1378 VTAIL.n105 VTAIL.n104 185
R1379 VTAIL.n107 VTAIL.n106 185
R1380 VTAIL.n255 VTAIL.n254 185
R1381 VTAIL.n253 VTAIL.n252 185
R1382 VTAIL.n228 VTAIL.n227 185
R1383 VTAIL.n247 VTAIL.n246 185
R1384 VTAIL.n245 VTAIL.n244 185
R1385 VTAIL.n232 VTAIL.n231 185
R1386 VTAIL.n239 VTAIL.n238 185
R1387 VTAIL.n237 VTAIL.n236 185
R1388 VTAIL.n217 VTAIL.n216 185
R1389 VTAIL.n215 VTAIL.n214 185
R1390 VTAIL.n190 VTAIL.n189 185
R1391 VTAIL.n209 VTAIL.n208 185
R1392 VTAIL.n207 VTAIL.n206 185
R1393 VTAIL.n194 VTAIL.n193 185
R1394 VTAIL.n201 VTAIL.n200 185
R1395 VTAIL.n199 VTAIL.n198 185
R1396 VTAIL.n181 VTAIL.n180 185
R1397 VTAIL.n179 VTAIL.n178 185
R1398 VTAIL.n154 VTAIL.n153 185
R1399 VTAIL.n173 VTAIL.n172 185
R1400 VTAIL.n171 VTAIL.n170 185
R1401 VTAIL.n158 VTAIL.n157 185
R1402 VTAIL.n165 VTAIL.n164 185
R1403 VTAIL.n163 VTAIL.n162 185
R1404 VTAIL.n143 VTAIL.n142 185
R1405 VTAIL.n141 VTAIL.n140 185
R1406 VTAIL.n116 VTAIL.n115 185
R1407 VTAIL.n135 VTAIL.n134 185
R1408 VTAIL.n133 VTAIL.n132 185
R1409 VTAIL.n120 VTAIL.n119 185
R1410 VTAIL.n127 VTAIL.n126 185
R1411 VTAIL.n125 VTAIL.n124 185
R1412 VTAIL.n271 VTAIL.t7 149.524
R1413 VTAIL.n13 VTAIL.t4 149.524
R1414 VTAIL.n49 VTAIL.t12 149.524
R1415 VTAIL.n87 VTAIL.t15 149.524
R1416 VTAIL.n235 VTAIL.t9 149.524
R1417 VTAIL.n197 VTAIL.t8 149.524
R1418 VTAIL.n161 VTAIL.t2 149.524
R1419 VTAIL.n123 VTAIL.t5 149.524
R1420 VTAIL.n274 VTAIL.n273 104.615
R1421 VTAIL.n274 VTAIL.n267 104.615
R1422 VTAIL.n281 VTAIL.n267 104.615
R1423 VTAIL.n282 VTAIL.n281 104.615
R1424 VTAIL.n282 VTAIL.n263 104.615
R1425 VTAIL.n289 VTAIL.n263 104.615
R1426 VTAIL.n290 VTAIL.n289 104.615
R1427 VTAIL.n16 VTAIL.n15 104.615
R1428 VTAIL.n16 VTAIL.n9 104.615
R1429 VTAIL.n23 VTAIL.n9 104.615
R1430 VTAIL.n24 VTAIL.n23 104.615
R1431 VTAIL.n24 VTAIL.n5 104.615
R1432 VTAIL.n31 VTAIL.n5 104.615
R1433 VTAIL.n32 VTAIL.n31 104.615
R1434 VTAIL.n52 VTAIL.n51 104.615
R1435 VTAIL.n52 VTAIL.n45 104.615
R1436 VTAIL.n59 VTAIL.n45 104.615
R1437 VTAIL.n60 VTAIL.n59 104.615
R1438 VTAIL.n60 VTAIL.n41 104.615
R1439 VTAIL.n67 VTAIL.n41 104.615
R1440 VTAIL.n68 VTAIL.n67 104.615
R1441 VTAIL.n90 VTAIL.n89 104.615
R1442 VTAIL.n90 VTAIL.n83 104.615
R1443 VTAIL.n97 VTAIL.n83 104.615
R1444 VTAIL.n98 VTAIL.n97 104.615
R1445 VTAIL.n98 VTAIL.n79 104.615
R1446 VTAIL.n105 VTAIL.n79 104.615
R1447 VTAIL.n106 VTAIL.n105 104.615
R1448 VTAIL.n254 VTAIL.n253 104.615
R1449 VTAIL.n253 VTAIL.n227 104.615
R1450 VTAIL.n246 VTAIL.n227 104.615
R1451 VTAIL.n246 VTAIL.n245 104.615
R1452 VTAIL.n245 VTAIL.n231 104.615
R1453 VTAIL.n238 VTAIL.n231 104.615
R1454 VTAIL.n238 VTAIL.n237 104.615
R1455 VTAIL.n216 VTAIL.n215 104.615
R1456 VTAIL.n215 VTAIL.n189 104.615
R1457 VTAIL.n208 VTAIL.n189 104.615
R1458 VTAIL.n208 VTAIL.n207 104.615
R1459 VTAIL.n207 VTAIL.n193 104.615
R1460 VTAIL.n200 VTAIL.n193 104.615
R1461 VTAIL.n200 VTAIL.n199 104.615
R1462 VTAIL.n180 VTAIL.n179 104.615
R1463 VTAIL.n179 VTAIL.n153 104.615
R1464 VTAIL.n172 VTAIL.n153 104.615
R1465 VTAIL.n172 VTAIL.n171 104.615
R1466 VTAIL.n171 VTAIL.n157 104.615
R1467 VTAIL.n164 VTAIL.n157 104.615
R1468 VTAIL.n164 VTAIL.n163 104.615
R1469 VTAIL.n142 VTAIL.n141 104.615
R1470 VTAIL.n141 VTAIL.n115 104.615
R1471 VTAIL.n134 VTAIL.n115 104.615
R1472 VTAIL.n134 VTAIL.n133 104.615
R1473 VTAIL.n133 VTAIL.n119 104.615
R1474 VTAIL.n126 VTAIL.n119 104.615
R1475 VTAIL.n126 VTAIL.n125 104.615
R1476 VTAIL.n273 VTAIL.t7 52.3082
R1477 VTAIL.n15 VTAIL.t4 52.3082
R1478 VTAIL.n51 VTAIL.t12 52.3082
R1479 VTAIL.n89 VTAIL.t15 52.3082
R1480 VTAIL.n237 VTAIL.t9 52.3082
R1481 VTAIL.n199 VTAIL.t8 52.3082
R1482 VTAIL.n163 VTAIL.t2 52.3082
R1483 VTAIL.n125 VTAIL.t5 52.3082
R1484 VTAIL.n223 VTAIL.n222 51.2531
R1485 VTAIL.n149 VTAIL.n148 51.2531
R1486 VTAIL.n1 VTAIL.n0 51.253
R1487 VTAIL.n75 VTAIL.n74 51.253
R1488 VTAIL.n295 VTAIL.n294 35.4823
R1489 VTAIL.n37 VTAIL.n36 35.4823
R1490 VTAIL.n73 VTAIL.n72 35.4823
R1491 VTAIL.n111 VTAIL.n110 35.4823
R1492 VTAIL.n259 VTAIL.n258 35.4823
R1493 VTAIL.n221 VTAIL.n220 35.4823
R1494 VTAIL.n185 VTAIL.n184 35.4823
R1495 VTAIL.n147 VTAIL.n146 35.4823
R1496 VTAIL.n295 VTAIL.n259 20.3496
R1497 VTAIL.n147 VTAIL.n111 20.3496
R1498 VTAIL.n292 VTAIL.n291 12.8005
R1499 VTAIL.n34 VTAIL.n33 12.8005
R1500 VTAIL.n70 VTAIL.n69 12.8005
R1501 VTAIL.n108 VTAIL.n107 12.8005
R1502 VTAIL.n256 VTAIL.n255 12.8005
R1503 VTAIL.n218 VTAIL.n217 12.8005
R1504 VTAIL.n182 VTAIL.n181 12.8005
R1505 VTAIL.n144 VTAIL.n143 12.8005
R1506 VTAIL.n288 VTAIL.n262 12.0247
R1507 VTAIL.n30 VTAIL.n4 12.0247
R1508 VTAIL.n66 VTAIL.n40 12.0247
R1509 VTAIL.n104 VTAIL.n78 12.0247
R1510 VTAIL.n252 VTAIL.n226 12.0247
R1511 VTAIL.n214 VTAIL.n188 12.0247
R1512 VTAIL.n178 VTAIL.n152 12.0247
R1513 VTAIL.n140 VTAIL.n114 12.0247
R1514 VTAIL.n287 VTAIL.n264 11.249
R1515 VTAIL.n29 VTAIL.n6 11.249
R1516 VTAIL.n65 VTAIL.n42 11.249
R1517 VTAIL.n103 VTAIL.n80 11.249
R1518 VTAIL.n251 VTAIL.n228 11.249
R1519 VTAIL.n213 VTAIL.n190 11.249
R1520 VTAIL.n177 VTAIL.n154 11.249
R1521 VTAIL.n139 VTAIL.n116 11.249
R1522 VTAIL.n284 VTAIL.n283 10.4732
R1523 VTAIL.n26 VTAIL.n25 10.4732
R1524 VTAIL.n62 VTAIL.n61 10.4732
R1525 VTAIL.n100 VTAIL.n99 10.4732
R1526 VTAIL.n248 VTAIL.n247 10.4732
R1527 VTAIL.n210 VTAIL.n209 10.4732
R1528 VTAIL.n174 VTAIL.n173 10.4732
R1529 VTAIL.n136 VTAIL.n135 10.4732
R1530 VTAIL.n272 VTAIL.n271 10.2747
R1531 VTAIL.n14 VTAIL.n13 10.2747
R1532 VTAIL.n50 VTAIL.n49 10.2747
R1533 VTAIL.n88 VTAIL.n87 10.2747
R1534 VTAIL.n236 VTAIL.n235 10.2747
R1535 VTAIL.n198 VTAIL.n197 10.2747
R1536 VTAIL.n162 VTAIL.n161 10.2747
R1537 VTAIL.n124 VTAIL.n123 10.2747
R1538 VTAIL.n280 VTAIL.n266 9.69747
R1539 VTAIL.n22 VTAIL.n8 9.69747
R1540 VTAIL.n58 VTAIL.n44 9.69747
R1541 VTAIL.n96 VTAIL.n82 9.69747
R1542 VTAIL.n244 VTAIL.n230 9.69747
R1543 VTAIL.n206 VTAIL.n192 9.69747
R1544 VTAIL.n170 VTAIL.n156 9.69747
R1545 VTAIL.n132 VTAIL.n118 9.69747
R1546 VTAIL.n294 VTAIL.n293 9.45567
R1547 VTAIL.n36 VTAIL.n35 9.45567
R1548 VTAIL.n72 VTAIL.n71 9.45567
R1549 VTAIL.n110 VTAIL.n109 9.45567
R1550 VTAIL.n258 VTAIL.n257 9.45567
R1551 VTAIL.n220 VTAIL.n219 9.45567
R1552 VTAIL.n184 VTAIL.n183 9.45567
R1553 VTAIL.n146 VTAIL.n145 9.45567
R1554 VTAIL.n270 VTAIL.n269 9.3005
R1555 VTAIL.n277 VTAIL.n276 9.3005
R1556 VTAIL.n279 VTAIL.n278 9.3005
R1557 VTAIL.n266 VTAIL.n265 9.3005
R1558 VTAIL.n285 VTAIL.n284 9.3005
R1559 VTAIL.n287 VTAIL.n286 9.3005
R1560 VTAIL.n262 VTAIL.n261 9.3005
R1561 VTAIL.n293 VTAIL.n292 9.3005
R1562 VTAIL.n12 VTAIL.n11 9.3005
R1563 VTAIL.n19 VTAIL.n18 9.3005
R1564 VTAIL.n21 VTAIL.n20 9.3005
R1565 VTAIL.n8 VTAIL.n7 9.3005
R1566 VTAIL.n27 VTAIL.n26 9.3005
R1567 VTAIL.n29 VTAIL.n28 9.3005
R1568 VTAIL.n4 VTAIL.n3 9.3005
R1569 VTAIL.n35 VTAIL.n34 9.3005
R1570 VTAIL.n48 VTAIL.n47 9.3005
R1571 VTAIL.n55 VTAIL.n54 9.3005
R1572 VTAIL.n57 VTAIL.n56 9.3005
R1573 VTAIL.n44 VTAIL.n43 9.3005
R1574 VTAIL.n63 VTAIL.n62 9.3005
R1575 VTAIL.n65 VTAIL.n64 9.3005
R1576 VTAIL.n40 VTAIL.n39 9.3005
R1577 VTAIL.n71 VTAIL.n70 9.3005
R1578 VTAIL.n86 VTAIL.n85 9.3005
R1579 VTAIL.n93 VTAIL.n92 9.3005
R1580 VTAIL.n95 VTAIL.n94 9.3005
R1581 VTAIL.n82 VTAIL.n81 9.3005
R1582 VTAIL.n101 VTAIL.n100 9.3005
R1583 VTAIL.n103 VTAIL.n102 9.3005
R1584 VTAIL.n78 VTAIL.n77 9.3005
R1585 VTAIL.n109 VTAIL.n108 9.3005
R1586 VTAIL.n234 VTAIL.n233 9.3005
R1587 VTAIL.n241 VTAIL.n240 9.3005
R1588 VTAIL.n243 VTAIL.n242 9.3005
R1589 VTAIL.n230 VTAIL.n229 9.3005
R1590 VTAIL.n249 VTAIL.n248 9.3005
R1591 VTAIL.n251 VTAIL.n250 9.3005
R1592 VTAIL.n226 VTAIL.n225 9.3005
R1593 VTAIL.n257 VTAIL.n256 9.3005
R1594 VTAIL.n196 VTAIL.n195 9.3005
R1595 VTAIL.n203 VTAIL.n202 9.3005
R1596 VTAIL.n205 VTAIL.n204 9.3005
R1597 VTAIL.n192 VTAIL.n191 9.3005
R1598 VTAIL.n211 VTAIL.n210 9.3005
R1599 VTAIL.n213 VTAIL.n212 9.3005
R1600 VTAIL.n188 VTAIL.n187 9.3005
R1601 VTAIL.n219 VTAIL.n218 9.3005
R1602 VTAIL.n160 VTAIL.n159 9.3005
R1603 VTAIL.n167 VTAIL.n166 9.3005
R1604 VTAIL.n169 VTAIL.n168 9.3005
R1605 VTAIL.n156 VTAIL.n155 9.3005
R1606 VTAIL.n175 VTAIL.n174 9.3005
R1607 VTAIL.n177 VTAIL.n176 9.3005
R1608 VTAIL.n152 VTAIL.n151 9.3005
R1609 VTAIL.n183 VTAIL.n182 9.3005
R1610 VTAIL.n122 VTAIL.n121 9.3005
R1611 VTAIL.n129 VTAIL.n128 9.3005
R1612 VTAIL.n131 VTAIL.n130 9.3005
R1613 VTAIL.n118 VTAIL.n117 9.3005
R1614 VTAIL.n137 VTAIL.n136 9.3005
R1615 VTAIL.n139 VTAIL.n138 9.3005
R1616 VTAIL.n114 VTAIL.n113 9.3005
R1617 VTAIL.n145 VTAIL.n144 9.3005
R1618 VTAIL.n279 VTAIL.n268 8.92171
R1619 VTAIL.n21 VTAIL.n10 8.92171
R1620 VTAIL.n57 VTAIL.n46 8.92171
R1621 VTAIL.n95 VTAIL.n84 8.92171
R1622 VTAIL.n243 VTAIL.n232 8.92171
R1623 VTAIL.n205 VTAIL.n194 8.92171
R1624 VTAIL.n169 VTAIL.n158 8.92171
R1625 VTAIL.n131 VTAIL.n120 8.92171
R1626 VTAIL.n294 VTAIL.n260 8.2187
R1627 VTAIL.n36 VTAIL.n2 8.2187
R1628 VTAIL.n72 VTAIL.n38 8.2187
R1629 VTAIL.n110 VTAIL.n76 8.2187
R1630 VTAIL.n258 VTAIL.n224 8.2187
R1631 VTAIL.n220 VTAIL.n186 8.2187
R1632 VTAIL.n184 VTAIL.n150 8.2187
R1633 VTAIL.n146 VTAIL.n112 8.2187
R1634 VTAIL.n276 VTAIL.n275 8.14595
R1635 VTAIL.n18 VTAIL.n17 8.14595
R1636 VTAIL.n54 VTAIL.n53 8.14595
R1637 VTAIL.n92 VTAIL.n91 8.14595
R1638 VTAIL.n240 VTAIL.n239 8.14595
R1639 VTAIL.n202 VTAIL.n201 8.14595
R1640 VTAIL.n166 VTAIL.n165 8.14595
R1641 VTAIL.n128 VTAIL.n127 8.14595
R1642 VTAIL.n272 VTAIL.n270 7.3702
R1643 VTAIL.n14 VTAIL.n12 7.3702
R1644 VTAIL.n50 VTAIL.n48 7.3702
R1645 VTAIL.n88 VTAIL.n86 7.3702
R1646 VTAIL.n236 VTAIL.n234 7.3702
R1647 VTAIL.n198 VTAIL.n196 7.3702
R1648 VTAIL.n162 VTAIL.n160 7.3702
R1649 VTAIL.n124 VTAIL.n122 7.3702
R1650 VTAIL.n275 VTAIL.n270 5.81868
R1651 VTAIL.n17 VTAIL.n12 5.81868
R1652 VTAIL.n53 VTAIL.n48 5.81868
R1653 VTAIL.n91 VTAIL.n86 5.81868
R1654 VTAIL.n239 VTAIL.n234 5.81868
R1655 VTAIL.n201 VTAIL.n196 5.81868
R1656 VTAIL.n165 VTAIL.n160 5.81868
R1657 VTAIL.n127 VTAIL.n122 5.81868
R1658 VTAIL.n292 VTAIL.n260 5.3904
R1659 VTAIL.n34 VTAIL.n2 5.3904
R1660 VTAIL.n70 VTAIL.n38 5.3904
R1661 VTAIL.n108 VTAIL.n76 5.3904
R1662 VTAIL.n256 VTAIL.n224 5.3904
R1663 VTAIL.n218 VTAIL.n186 5.3904
R1664 VTAIL.n182 VTAIL.n150 5.3904
R1665 VTAIL.n144 VTAIL.n112 5.3904
R1666 VTAIL.n276 VTAIL.n268 5.04292
R1667 VTAIL.n18 VTAIL.n10 5.04292
R1668 VTAIL.n54 VTAIL.n46 5.04292
R1669 VTAIL.n92 VTAIL.n84 5.04292
R1670 VTAIL.n240 VTAIL.n232 5.04292
R1671 VTAIL.n202 VTAIL.n194 5.04292
R1672 VTAIL.n166 VTAIL.n158 5.04292
R1673 VTAIL.n128 VTAIL.n120 5.04292
R1674 VTAIL.n280 VTAIL.n279 4.26717
R1675 VTAIL.n22 VTAIL.n21 4.26717
R1676 VTAIL.n58 VTAIL.n57 4.26717
R1677 VTAIL.n96 VTAIL.n95 4.26717
R1678 VTAIL.n244 VTAIL.n243 4.26717
R1679 VTAIL.n206 VTAIL.n205 4.26717
R1680 VTAIL.n170 VTAIL.n169 4.26717
R1681 VTAIL.n132 VTAIL.n131 4.26717
R1682 VTAIL.n283 VTAIL.n266 3.49141
R1683 VTAIL.n25 VTAIL.n8 3.49141
R1684 VTAIL.n61 VTAIL.n44 3.49141
R1685 VTAIL.n99 VTAIL.n82 3.49141
R1686 VTAIL.n247 VTAIL.n230 3.49141
R1687 VTAIL.n209 VTAIL.n192 3.49141
R1688 VTAIL.n173 VTAIL.n156 3.49141
R1689 VTAIL.n135 VTAIL.n118 3.49141
R1690 VTAIL.n271 VTAIL.n269 2.84305
R1691 VTAIL.n13 VTAIL.n11 2.84305
R1692 VTAIL.n49 VTAIL.n47 2.84305
R1693 VTAIL.n87 VTAIL.n85 2.84305
R1694 VTAIL.n235 VTAIL.n233 2.84305
R1695 VTAIL.n197 VTAIL.n195 2.84305
R1696 VTAIL.n161 VTAIL.n159 2.84305
R1697 VTAIL.n123 VTAIL.n121 2.84305
R1698 VTAIL.n0 VTAIL.t3 2.73153
R1699 VTAIL.n0 VTAIL.t0 2.73153
R1700 VTAIL.n74 VTAIL.t10 2.73153
R1701 VTAIL.n74 VTAIL.t11 2.73153
R1702 VTAIL.n222 VTAIL.t14 2.73153
R1703 VTAIL.n222 VTAIL.t13 2.73153
R1704 VTAIL.n148 VTAIL.t1 2.73153
R1705 VTAIL.n148 VTAIL.t6 2.73153
R1706 VTAIL.n284 VTAIL.n264 2.71565
R1707 VTAIL.n26 VTAIL.n6 2.71565
R1708 VTAIL.n62 VTAIL.n42 2.71565
R1709 VTAIL.n100 VTAIL.n80 2.71565
R1710 VTAIL.n248 VTAIL.n228 2.71565
R1711 VTAIL.n210 VTAIL.n190 2.71565
R1712 VTAIL.n174 VTAIL.n154 2.71565
R1713 VTAIL.n136 VTAIL.n116 2.71565
R1714 VTAIL.n288 VTAIL.n287 1.93989
R1715 VTAIL.n30 VTAIL.n29 1.93989
R1716 VTAIL.n66 VTAIL.n65 1.93989
R1717 VTAIL.n104 VTAIL.n103 1.93989
R1718 VTAIL.n252 VTAIL.n251 1.93989
R1719 VTAIL.n214 VTAIL.n213 1.93989
R1720 VTAIL.n178 VTAIL.n177 1.93989
R1721 VTAIL.n140 VTAIL.n139 1.93989
R1722 VTAIL.n149 VTAIL.n147 1.73326
R1723 VTAIL.n185 VTAIL.n149 1.73326
R1724 VTAIL.n223 VTAIL.n221 1.73326
R1725 VTAIL.n259 VTAIL.n223 1.73326
R1726 VTAIL.n111 VTAIL.n75 1.73326
R1727 VTAIL.n75 VTAIL.n73 1.73326
R1728 VTAIL.n37 VTAIL.n1 1.73326
R1729 VTAIL VTAIL.n295 1.67507
R1730 VTAIL.n291 VTAIL.n262 1.16414
R1731 VTAIL.n33 VTAIL.n4 1.16414
R1732 VTAIL.n69 VTAIL.n40 1.16414
R1733 VTAIL.n107 VTAIL.n78 1.16414
R1734 VTAIL.n255 VTAIL.n226 1.16414
R1735 VTAIL.n217 VTAIL.n188 1.16414
R1736 VTAIL.n181 VTAIL.n152 1.16414
R1737 VTAIL.n143 VTAIL.n114 1.16414
R1738 VTAIL.n221 VTAIL.n185 0.470328
R1739 VTAIL.n73 VTAIL.n37 0.470328
R1740 VTAIL.n277 VTAIL.n269 0.155672
R1741 VTAIL.n278 VTAIL.n277 0.155672
R1742 VTAIL.n278 VTAIL.n265 0.155672
R1743 VTAIL.n285 VTAIL.n265 0.155672
R1744 VTAIL.n286 VTAIL.n285 0.155672
R1745 VTAIL.n286 VTAIL.n261 0.155672
R1746 VTAIL.n293 VTAIL.n261 0.155672
R1747 VTAIL.n19 VTAIL.n11 0.155672
R1748 VTAIL.n20 VTAIL.n19 0.155672
R1749 VTAIL.n20 VTAIL.n7 0.155672
R1750 VTAIL.n27 VTAIL.n7 0.155672
R1751 VTAIL.n28 VTAIL.n27 0.155672
R1752 VTAIL.n28 VTAIL.n3 0.155672
R1753 VTAIL.n35 VTAIL.n3 0.155672
R1754 VTAIL.n55 VTAIL.n47 0.155672
R1755 VTAIL.n56 VTAIL.n55 0.155672
R1756 VTAIL.n56 VTAIL.n43 0.155672
R1757 VTAIL.n63 VTAIL.n43 0.155672
R1758 VTAIL.n64 VTAIL.n63 0.155672
R1759 VTAIL.n64 VTAIL.n39 0.155672
R1760 VTAIL.n71 VTAIL.n39 0.155672
R1761 VTAIL.n93 VTAIL.n85 0.155672
R1762 VTAIL.n94 VTAIL.n93 0.155672
R1763 VTAIL.n94 VTAIL.n81 0.155672
R1764 VTAIL.n101 VTAIL.n81 0.155672
R1765 VTAIL.n102 VTAIL.n101 0.155672
R1766 VTAIL.n102 VTAIL.n77 0.155672
R1767 VTAIL.n109 VTAIL.n77 0.155672
R1768 VTAIL.n257 VTAIL.n225 0.155672
R1769 VTAIL.n250 VTAIL.n225 0.155672
R1770 VTAIL.n250 VTAIL.n249 0.155672
R1771 VTAIL.n249 VTAIL.n229 0.155672
R1772 VTAIL.n242 VTAIL.n229 0.155672
R1773 VTAIL.n242 VTAIL.n241 0.155672
R1774 VTAIL.n241 VTAIL.n233 0.155672
R1775 VTAIL.n219 VTAIL.n187 0.155672
R1776 VTAIL.n212 VTAIL.n187 0.155672
R1777 VTAIL.n212 VTAIL.n211 0.155672
R1778 VTAIL.n211 VTAIL.n191 0.155672
R1779 VTAIL.n204 VTAIL.n191 0.155672
R1780 VTAIL.n204 VTAIL.n203 0.155672
R1781 VTAIL.n203 VTAIL.n195 0.155672
R1782 VTAIL.n183 VTAIL.n151 0.155672
R1783 VTAIL.n176 VTAIL.n151 0.155672
R1784 VTAIL.n176 VTAIL.n175 0.155672
R1785 VTAIL.n175 VTAIL.n155 0.155672
R1786 VTAIL.n168 VTAIL.n155 0.155672
R1787 VTAIL.n168 VTAIL.n167 0.155672
R1788 VTAIL.n167 VTAIL.n159 0.155672
R1789 VTAIL.n145 VTAIL.n113 0.155672
R1790 VTAIL.n138 VTAIL.n113 0.155672
R1791 VTAIL.n138 VTAIL.n137 0.155672
R1792 VTAIL.n137 VTAIL.n117 0.155672
R1793 VTAIL.n130 VTAIL.n117 0.155672
R1794 VTAIL.n130 VTAIL.n129 0.155672
R1795 VTAIL.n129 VTAIL.n121 0.155672
R1796 VTAIL VTAIL.n1 0.0586897
R1797 VN.n22 VN.n21 185.034
R1798 VN.n45 VN.n44 185.034
R1799 VN.n43 VN.n23 161.3
R1800 VN.n42 VN.n41 161.3
R1801 VN.n40 VN.n24 161.3
R1802 VN.n39 VN.n38 161.3
R1803 VN.n36 VN.n25 161.3
R1804 VN.n35 VN.n34 161.3
R1805 VN.n33 VN.n26 161.3
R1806 VN.n32 VN.n31 161.3
R1807 VN.n30 VN.n27 161.3
R1808 VN.n20 VN.n0 161.3
R1809 VN.n19 VN.n18 161.3
R1810 VN.n17 VN.n1 161.3
R1811 VN.n16 VN.n15 161.3
R1812 VN.n13 VN.n2 161.3
R1813 VN.n12 VN.n11 161.3
R1814 VN.n10 VN.n3 161.3
R1815 VN.n9 VN.n8 161.3
R1816 VN.n7 VN.n4 161.3
R1817 VN.n5 VN.t3 131.504
R1818 VN.n28 VN.t4 131.504
R1819 VN.n6 VN.t5 104.004
R1820 VN.n14 VN.t1 104.004
R1821 VN.n21 VN.t2 104.004
R1822 VN.n29 VN.t6 104.004
R1823 VN.n37 VN.t7 104.004
R1824 VN.n44 VN.t0 104.004
R1825 VN.n6 VN.n5 68.7155
R1826 VN.n29 VN.n28 68.7155
R1827 VN VN.n45 43.1994
R1828 VN.n19 VN.n1 41.4647
R1829 VN.n42 VN.n24 41.4647
R1830 VN.n8 VN.n3 40.4934
R1831 VN.n12 VN.n3 40.4934
R1832 VN.n31 VN.n26 40.4934
R1833 VN.n35 VN.n26 40.4934
R1834 VN.n15 VN.n1 39.5221
R1835 VN.n38 VN.n24 39.5221
R1836 VN.n8 VN.n7 24.4675
R1837 VN.n13 VN.n12 24.4675
R1838 VN.n20 VN.n19 24.4675
R1839 VN.n31 VN.n30 24.4675
R1840 VN.n36 VN.n35 24.4675
R1841 VN.n43 VN.n42 24.4675
R1842 VN.n15 VN.n14 24.2228
R1843 VN.n38 VN.n37 24.2228
R1844 VN.n28 VN.n27 18.9997
R1845 VN.n5 VN.n4 18.9997
R1846 VN.n21 VN.n20 0.73451
R1847 VN.n44 VN.n43 0.73451
R1848 VN.n7 VN.n6 0.24517
R1849 VN.n14 VN.n13 0.24517
R1850 VN.n30 VN.n29 0.24517
R1851 VN.n37 VN.n36 0.24517
R1852 VN.n45 VN.n23 0.189894
R1853 VN.n41 VN.n23 0.189894
R1854 VN.n41 VN.n40 0.189894
R1855 VN.n40 VN.n39 0.189894
R1856 VN.n39 VN.n25 0.189894
R1857 VN.n34 VN.n25 0.189894
R1858 VN.n34 VN.n33 0.189894
R1859 VN.n33 VN.n32 0.189894
R1860 VN.n32 VN.n27 0.189894
R1861 VN.n9 VN.n4 0.189894
R1862 VN.n10 VN.n9 0.189894
R1863 VN.n11 VN.n10 0.189894
R1864 VN.n11 VN.n2 0.189894
R1865 VN.n16 VN.n2 0.189894
R1866 VN.n17 VN.n16 0.189894
R1867 VN.n18 VN.n17 0.189894
R1868 VN.n18 VN.n0 0.189894
R1869 VN.n22 VN.n0 0.189894
R1870 VN VN.n22 0.0516364
R1871 VDD2.n2 VDD2.n1 68.7428
R1872 VDD2.n2 VDD2.n0 68.7428
R1873 VDD2 VDD2.n5 68.74
R1874 VDD2.n4 VDD2.n3 67.9319
R1875 VDD2.n4 VDD2.n2 37.7627
R1876 VDD2.n5 VDD2.t1 2.73153
R1877 VDD2.n5 VDD2.t3 2.73153
R1878 VDD2.n3 VDD2.t7 2.73153
R1879 VDD2.n3 VDD2.t0 2.73153
R1880 VDD2.n1 VDD2.t6 2.73153
R1881 VDD2.n1 VDD2.t5 2.73153
R1882 VDD2.n0 VDD2.t4 2.73153
R1883 VDD2.n0 VDD2.t2 2.73153
R1884 VDD2 VDD2.n4 0.925069
C0 VTAIL VP 5.20967f
C1 VTAIL VN 5.19556f
C2 VDD1 VP 5.17538f
C3 VDD1 VN 0.149573f
C4 VDD2 VTAIL 6.28099f
C5 VDD2 VDD1 1.29537f
C6 VN VP 5.66091f
C7 VTAIL VDD1 6.23275f
C8 VDD2 VP 0.421282f
C9 VDD2 VN 4.9046f
C10 VDD2 B 4.083084f
C11 VDD1 B 4.42217f
C12 VTAIL B 6.996604f
C13 VN B 11.60905f
C14 VP B 10.152308f
C15 VDD2.t4 B 0.141787f
C16 VDD2.t2 B 0.141787f
C17 VDD2.n0 B 1.22282f
C18 VDD2.t6 B 0.141787f
C19 VDD2.t5 B 0.141787f
C20 VDD2.n1 B 1.22282f
C21 VDD2.n2 B 2.41044f
C22 VDD2.t7 B 0.141787f
C23 VDD2.t0 B 0.141787f
C24 VDD2.n3 B 1.21802f
C25 VDD2.n4 B 2.22874f
C26 VDD2.t1 B 0.141787f
C27 VDD2.t3 B 0.141787f
C28 VDD2.n5 B 1.22279f
C29 VN.n0 B 0.030391f
C30 VN.t2 B 0.989673f
C31 VN.n1 B 0.024607f
C32 VN.n2 B 0.030391f
C33 VN.t1 B 0.989673f
C34 VN.n3 B 0.024568f
C35 VN.n4 B 0.191913f
C36 VN.t5 B 0.989673f
C37 VN.t3 B 1.09425f
C38 VN.n5 B 0.454524f
C39 VN.n6 B 0.424915f
C40 VN.n7 B 0.028955f
C41 VN.n8 B 0.060402f
C42 VN.n9 B 0.030391f
C43 VN.n10 B 0.030391f
C44 VN.n11 B 0.030391f
C45 VN.n12 B 0.060402f
C46 VN.n13 B 0.028955f
C47 VN.n14 B 0.373751f
C48 VN.n15 B 0.060406f
C49 VN.n16 B 0.030391f
C50 VN.n17 B 0.030391f
C51 VN.n18 B 0.030391f
C52 VN.n19 B 0.060078f
C53 VN.n20 B 0.029515f
C54 VN.n21 B 0.432633f
C55 VN.n22 B 0.032215f
C56 VN.n23 B 0.030391f
C57 VN.t0 B 0.989673f
C58 VN.n24 B 0.024607f
C59 VN.n25 B 0.030391f
C60 VN.t7 B 0.989673f
C61 VN.n26 B 0.024568f
C62 VN.n27 B 0.191913f
C63 VN.t6 B 0.989673f
C64 VN.t4 B 1.09425f
C65 VN.n28 B 0.454524f
C66 VN.n29 B 0.424915f
C67 VN.n30 B 0.028955f
C68 VN.n31 B 0.060402f
C69 VN.n32 B 0.030391f
C70 VN.n33 B 0.030391f
C71 VN.n34 B 0.030391f
C72 VN.n35 B 0.060402f
C73 VN.n36 B 0.028955f
C74 VN.n37 B 0.373751f
C75 VN.n38 B 0.060406f
C76 VN.n39 B 0.030391f
C77 VN.n40 B 0.030391f
C78 VN.n41 B 0.030391f
C79 VN.n42 B 0.060078f
C80 VN.n43 B 0.029515f
C81 VN.n44 B 0.432633f
C82 VN.n45 B 1.32378f
C83 VTAIL.t3 B 0.120163f
C84 VTAIL.t0 B 0.120163f
C85 VTAIL.n0 B 0.980023f
C86 VTAIL.n1 B 0.309239f
C87 VTAIL.n2 B 0.028927f
C88 VTAIL.n3 B 0.020974f
C89 VTAIL.n4 B 0.01127f
C90 VTAIL.n5 B 0.026639f
C91 VTAIL.n6 B 0.011933f
C92 VTAIL.n7 B 0.020974f
C93 VTAIL.n8 B 0.01127f
C94 VTAIL.n9 B 0.026639f
C95 VTAIL.n10 B 0.011933f
C96 VTAIL.n11 B 0.61489f
C97 VTAIL.n12 B 0.01127f
C98 VTAIL.t4 B 0.044485f
C99 VTAIL.n13 B 0.113023f
C100 VTAIL.n14 B 0.018832f
C101 VTAIL.n15 B 0.019979f
C102 VTAIL.n16 B 0.026639f
C103 VTAIL.n17 B 0.011933f
C104 VTAIL.n18 B 0.01127f
C105 VTAIL.n19 B 0.020974f
C106 VTAIL.n20 B 0.020974f
C107 VTAIL.n21 B 0.01127f
C108 VTAIL.n22 B 0.011933f
C109 VTAIL.n23 B 0.026639f
C110 VTAIL.n24 B 0.026639f
C111 VTAIL.n25 B 0.011933f
C112 VTAIL.n26 B 0.01127f
C113 VTAIL.n27 B 0.020974f
C114 VTAIL.n28 B 0.020974f
C115 VTAIL.n29 B 0.01127f
C116 VTAIL.n30 B 0.011933f
C117 VTAIL.n31 B 0.026639f
C118 VTAIL.n32 B 0.054766f
C119 VTAIL.n33 B 0.011933f
C120 VTAIL.n34 B 0.022037f
C121 VTAIL.n35 B 0.053351f
C122 VTAIL.n36 B 0.056879f
C123 VTAIL.n37 B 0.169525f
C124 VTAIL.n38 B 0.028927f
C125 VTAIL.n39 B 0.020974f
C126 VTAIL.n40 B 0.01127f
C127 VTAIL.n41 B 0.026639f
C128 VTAIL.n42 B 0.011933f
C129 VTAIL.n43 B 0.020974f
C130 VTAIL.n44 B 0.01127f
C131 VTAIL.n45 B 0.026639f
C132 VTAIL.n46 B 0.011933f
C133 VTAIL.n47 B 0.61489f
C134 VTAIL.n48 B 0.01127f
C135 VTAIL.t12 B 0.044485f
C136 VTAIL.n49 B 0.113023f
C137 VTAIL.n50 B 0.018832f
C138 VTAIL.n51 B 0.019979f
C139 VTAIL.n52 B 0.026639f
C140 VTAIL.n53 B 0.011933f
C141 VTAIL.n54 B 0.01127f
C142 VTAIL.n55 B 0.020974f
C143 VTAIL.n56 B 0.020974f
C144 VTAIL.n57 B 0.01127f
C145 VTAIL.n58 B 0.011933f
C146 VTAIL.n59 B 0.026639f
C147 VTAIL.n60 B 0.026639f
C148 VTAIL.n61 B 0.011933f
C149 VTAIL.n62 B 0.01127f
C150 VTAIL.n63 B 0.020974f
C151 VTAIL.n64 B 0.020974f
C152 VTAIL.n65 B 0.01127f
C153 VTAIL.n66 B 0.011933f
C154 VTAIL.n67 B 0.026639f
C155 VTAIL.n68 B 0.054766f
C156 VTAIL.n69 B 0.011933f
C157 VTAIL.n70 B 0.022037f
C158 VTAIL.n71 B 0.053351f
C159 VTAIL.n72 B 0.056879f
C160 VTAIL.n73 B 0.169525f
C161 VTAIL.t10 B 0.120163f
C162 VTAIL.t11 B 0.120163f
C163 VTAIL.n74 B 0.980023f
C164 VTAIL.n75 B 0.42241f
C165 VTAIL.n76 B 0.028927f
C166 VTAIL.n77 B 0.020974f
C167 VTAIL.n78 B 0.01127f
C168 VTAIL.n79 B 0.026639f
C169 VTAIL.n80 B 0.011933f
C170 VTAIL.n81 B 0.020974f
C171 VTAIL.n82 B 0.01127f
C172 VTAIL.n83 B 0.026639f
C173 VTAIL.n84 B 0.011933f
C174 VTAIL.n85 B 0.61489f
C175 VTAIL.n86 B 0.01127f
C176 VTAIL.t15 B 0.044485f
C177 VTAIL.n87 B 0.113023f
C178 VTAIL.n88 B 0.018832f
C179 VTAIL.n89 B 0.019979f
C180 VTAIL.n90 B 0.026639f
C181 VTAIL.n91 B 0.011933f
C182 VTAIL.n92 B 0.01127f
C183 VTAIL.n93 B 0.020974f
C184 VTAIL.n94 B 0.020974f
C185 VTAIL.n95 B 0.01127f
C186 VTAIL.n96 B 0.011933f
C187 VTAIL.n97 B 0.026639f
C188 VTAIL.n98 B 0.026639f
C189 VTAIL.n99 B 0.011933f
C190 VTAIL.n100 B 0.01127f
C191 VTAIL.n101 B 0.020974f
C192 VTAIL.n102 B 0.020974f
C193 VTAIL.n103 B 0.01127f
C194 VTAIL.n104 B 0.011933f
C195 VTAIL.n105 B 0.026639f
C196 VTAIL.n106 B 0.054766f
C197 VTAIL.n107 B 0.011933f
C198 VTAIL.n108 B 0.022037f
C199 VTAIL.n109 B 0.053351f
C200 VTAIL.n110 B 0.056879f
C201 VTAIL.n111 B 0.962171f
C202 VTAIL.n112 B 0.028927f
C203 VTAIL.n113 B 0.020974f
C204 VTAIL.n114 B 0.01127f
C205 VTAIL.n115 B 0.026639f
C206 VTAIL.n116 B 0.011933f
C207 VTAIL.n117 B 0.020974f
C208 VTAIL.n118 B 0.01127f
C209 VTAIL.n119 B 0.026639f
C210 VTAIL.n120 B 0.011933f
C211 VTAIL.n121 B 0.61489f
C212 VTAIL.n122 B 0.01127f
C213 VTAIL.t5 B 0.044485f
C214 VTAIL.n123 B 0.113023f
C215 VTAIL.n124 B 0.018832f
C216 VTAIL.n125 B 0.019979f
C217 VTAIL.n126 B 0.026639f
C218 VTAIL.n127 B 0.011933f
C219 VTAIL.n128 B 0.01127f
C220 VTAIL.n129 B 0.020974f
C221 VTAIL.n130 B 0.020974f
C222 VTAIL.n131 B 0.01127f
C223 VTAIL.n132 B 0.011933f
C224 VTAIL.n133 B 0.026639f
C225 VTAIL.n134 B 0.026639f
C226 VTAIL.n135 B 0.011933f
C227 VTAIL.n136 B 0.01127f
C228 VTAIL.n137 B 0.020974f
C229 VTAIL.n138 B 0.020974f
C230 VTAIL.n139 B 0.01127f
C231 VTAIL.n140 B 0.011933f
C232 VTAIL.n141 B 0.026639f
C233 VTAIL.n142 B 0.054766f
C234 VTAIL.n143 B 0.011933f
C235 VTAIL.n144 B 0.022037f
C236 VTAIL.n145 B 0.053351f
C237 VTAIL.n146 B 0.056879f
C238 VTAIL.n147 B 0.962171f
C239 VTAIL.t1 B 0.120163f
C240 VTAIL.t6 B 0.120163f
C241 VTAIL.n148 B 0.98003f
C242 VTAIL.n149 B 0.422404f
C243 VTAIL.n150 B 0.028927f
C244 VTAIL.n151 B 0.020974f
C245 VTAIL.n152 B 0.01127f
C246 VTAIL.n153 B 0.026639f
C247 VTAIL.n154 B 0.011933f
C248 VTAIL.n155 B 0.020974f
C249 VTAIL.n156 B 0.01127f
C250 VTAIL.n157 B 0.026639f
C251 VTAIL.n158 B 0.011933f
C252 VTAIL.n159 B 0.61489f
C253 VTAIL.n160 B 0.01127f
C254 VTAIL.t2 B 0.044485f
C255 VTAIL.n161 B 0.113023f
C256 VTAIL.n162 B 0.018832f
C257 VTAIL.n163 B 0.019979f
C258 VTAIL.n164 B 0.026639f
C259 VTAIL.n165 B 0.011933f
C260 VTAIL.n166 B 0.01127f
C261 VTAIL.n167 B 0.020974f
C262 VTAIL.n168 B 0.020974f
C263 VTAIL.n169 B 0.01127f
C264 VTAIL.n170 B 0.011933f
C265 VTAIL.n171 B 0.026639f
C266 VTAIL.n172 B 0.026639f
C267 VTAIL.n173 B 0.011933f
C268 VTAIL.n174 B 0.01127f
C269 VTAIL.n175 B 0.020974f
C270 VTAIL.n176 B 0.020974f
C271 VTAIL.n177 B 0.01127f
C272 VTAIL.n178 B 0.011933f
C273 VTAIL.n179 B 0.026639f
C274 VTAIL.n180 B 0.054766f
C275 VTAIL.n181 B 0.011933f
C276 VTAIL.n182 B 0.022037f
C277 VTAIL.n183 B 0.053351f
C278 VTAIL.n184 B 0.056879f
C279 VTAIL.n185 B 0.169525f
C280 VTAIL.n186 B 0.028927f
C281 VTAIL.n187 B 0.020974f
C282 VTAIL.n188 B 0.01127f
C283 VTAIL.n189 B 0.026639f
C284 VTAIL.n190 B 0.011933f
C285 VTAIL.n191 B 0.020974f
C286 VTAIL.n192 B 0.01127f
C287 VTAIL.n193 B 0.026639f
C288 VTAIL.n194 B 0.011933f
C289 VTAIL.n195 B 0.61489f
C290 VTAIL.n196 B 0.01127f
C291 VTAIL.t8 B 0.044485f
C292 VTAIL.n197 B 0.113023f
C293 VTAIL.n198 B 0.018832f
C294 VTAIL.n199 B 0.019979f
C295 VTAIL.n200 B 0.026639f
C296 VTAIL.n201 B 0.011933f
C297 VTAIL.n202 B 0.01127f
C298 VTAIL.n203 B 0.020974f
C299 VTAIL.n204 B 0.020974f
C300 VTAIL.n205 B 0.01127f
C301 VTAIL.n206 B 0.011933f
C302 VTAIL.n207 B 0.026639f
C303 VTAIL.n208 B 0.026639f
C304 VTAIL.n209 B 0.011933f
C305 VTAIL.n210 B 0.01127f
C306 VTAIL.n211 B 0.020974f
C307 VTAIL.n212 B 0.020974f
C308 VTAIL.n213 B 0.01127f
C309 VTAIL.n214 B 0.011933f
C310 VTAIL.n215 B 0.026639f
C311 VTAIL.n216 B 0.054766f
C312 VTAIL.n217 B 0.011933f
C313 VTAIL.n218 B 0.022037f
C314 VTAIL.n219 B 0.053351f
C315 VTAIL.n220 B 0.056879f
C316 VTAIL.n221 B 0.169525f
C317 VTAIL.t14 B 0.120163f
C318 VTAIL.t13 B 0.120163f
C319 VTAIL.n222 B 0.98003f
C320 VTAIL.n223 B 0.422404f
C321 VTAIL.n224 B 0.028927f
C322 VTAIL.n225 B 0.020974f
C323 VTAIL.n226 B 0.01127f
C324 VTAIL.n227 B 0.026639f
C325 VTAIL.n228 B 0.011933f
C326 VTAIL.n229 B 0.020974f
C327 VTAIL.n230 B 0.01127f
C328 VTAIL.n231 B 0.026639f
C329 VTAIL.n232 B 0.011933f
C330 VTAIL.n233 B 0.61489f
C331 VTAIL.n234 B 0.01127f
C332 VTAIL.t9 B 0.044485f
C333 VTAIL.n235 B 0.113023f
C334 VTAIL.n236 B 0.018832f
C335 VTAIL.n237 B 0.019979f
C336 VTAIL.n238 B 0.026639f
C337 VTAIL.n239 B 0.011933f
C338 VTAIL.n240 B 0.01127f
C339 VTAIL.n241 B 0.020974f
C340 VTAIL.n242 B 0.020974f
C341 VTAIL.n243 B 0.01127f
C342 VTAIL.n244 B 0.011933f
C343 VTAIL.n245 B 0.026639f
C344 VTAIL.n246 B 0.026639f
C345 VTAIL.n247 B 0.011933f
C346 VTAIL.n248 B 0.01127f
C347 VTAIL.n249 B 0.020974f
C348 VTAIL.n250 B 0.020974f
C349 VTAIL.n251 B 0.01127f
C350 VTAIL.n252 B 0.011933f
C351 VTAIL.n253 B 0.026639f
C352 VTAIL.n254 B 0.054766f
C353 VTAIL.n255 B 0.011933f
C354 VTAIL.n256 B 0.022037f
C355 VTAIL.n257 B 0.053351f
C356 VTAIL.n258 B 0.056879f
C357 VTAIL.n259 B 0.96217f
C358 VTAIL.n260 B 0.028927f
C359 VTAIL.n261 B 0.020974f
C360 VTAIL.n262 B 0.01127f
C361 VTAIL.n263 B 0.026639f
C362 VTAIL.n264 B 0.011933f
C363 VTAIL.n265 B 0.020974f
C364 VTAIL.n266 B 0.01127f
C365 VTAIL.n267 B 0.026639f
C366 VTAIL.n268 B 0.011933f
C367 VTAIL.n269 B 0.61489f
C368 VTAIL.n270 B 0.01127f
C369 VTAIL.t7 B 0.044485f
C370 VTAIL.n271 B 0.113023f
C371 VTAIL.n272 B 0.018832f
C372 VTAIL.n273 B 0.019979f
C373 VTAIL.n274 B 0.026639f
C374 VTAIL.n275 B 0.011933f
C375 VTAIL.n276 B 0.01127f
C376 VTAIL.n277 B 0.020974f
C377 VTAIL.n278 B 0.020974f
C378 VTAIL.n279 B 0.01127f
C379 VTAIL.n280 B 0.011933f
C380 VTAIL.n281 B 0.026639f
C381 VTAIL.n282 B 0.026639f
C382 VTAIL.n283 B 0.011933f
C383 VTAIL.n284 B 0.01127f
C384 VTAIL.n285 B 0.020974f
C385 VTAIL.n286 B 0.020974f
C386 VTAIL.n287 B 0.01127f
C387 VTAIL.n288 B 0.011933f
C388 VTAIL.n289 B 0.026639f
C389 VTAIL.n290 B 0.054766f
C390 VTAIL.n291 B 0.011933f
C391 VTAIL.n292 B 0.022037f
C392 VTAIL.n293 B 0.053351f
C393 VTAIL.n294 B 0.056879f
C394 VTAIL.n295 B 0.958238f
C395 VDD1.t5 B 0.14315f
C396 VDD1.t6 B 0.14315f
C397 VDD1.n0 B 1.23537f
C398 VDD1.t1 B 0.14315f
C399 VDD1.t4 B 0.14315f
C400 VDD1.n1 B 1.23458f
C401 VDD1.t7 B 0.14315f
C402 VDD1.t2 B 0.14315f
C403 VDD1.n2 B 1.23458f
C404 VDD1.n3 B 2.4864f
C405 VDD1.t0 B 0.14315f
C406 VDD1.t3 B 0.14315f
C407 VDD1.n4 B 1.22973f
C408 VDD1.n5 B 2.28031f
C409 VP.n0 B 0.031052f
C410 VP.t3 B 1.0112f
C411 VP.n1 B 0.025143f
C412 VP.n2 B 0.031052f
C413 VP.t4 B 1.0112f
C414 VP.n3 B 0.025103f
C415 VP.n4 B 0.031052f
C416 VP.t5 B 1.0112f
C417 VP.n5 B 0.025143f
C418 VP.n6 B 0.031052f
C419 VP.t0 B 1.0112f
C420 VP.n7 B 0.031052f
C421 VP.t6 B 1.0112f
C422 VP.n8 B 0.025143f
C423 VP.n9 B 0.031052f
C424 VP.t2 B 1.0112f
C425 VP.n10 B 0.025103f
C426 VP.n11 B 0.196087f
C427 VP.t1 B 1.0112f
C428 VP.t7 B 1.11805f
C429 VP.n12 B 0.46441f
C430 VP.n13 B 0.434156f
C431 VP.n14 B 0.029585f
C432 VP.n15 B 0.061716f
C433 VP.n16 B 0.031052f
C434 VP.n17 B 0.031052f
C435 VP.n18 B 0.031052f
C436 VP.n19 B 0.061716f
C437 VP.n20 B 0.029585f
C438 VP.n21 B 0.38188f
C439 VP.n22 B 0.061719f
C440 VP.n23 B 0.031052f
C441 VP.n24 B 0.031052f
C442 VP.n25 B 0.031052f
C443 VP.n26 B 0.061384f
C444 VP.n27 B 0.030157f
C445 VP.n28 B 0.442043f
C446 VP.n29 B 1.33222f
C447 VP.n30 B 1.35828f
C448 VP.n31 B 0.442043f
C449 VP.n32 B 0.030157f
C450 VP.n33 B 0.061384f
C451 VP.n34 B 0.031052f
C452 VP.n35 B 0.031052f
C453 VP.n36 B 0.031052f
C454 VP.n37 B 0.061719f
C455 VP.n38 B 0.38188f
C456 VP.n39 B 0.029585f
C457 VP.n40 B 0.061716f
C458 VP.n41 B 0.031052f
C459 VP.n42 B 0.031052f
C460 VP.n43 B 0.031052f
C461 VP.n44 B 0.061716f
C462 VP.n45 B 0.029585f
C463 VP.n46 B 0.38188f
C464 VP.n47 B 0.061719f
C465 VP.n48 B 0.031052f
C466 VP.n49 B 0.031052f
C467 VP.n50 B 0.031052f
C468 VP.n51 B 0.061384f
C469 VP.n52 B 0.030157f
C470 VP.n53 B 0.442043f
C471 VP.n54 B 0.032916f
.ends

