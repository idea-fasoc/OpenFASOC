* NGSPICE file created from diff_pair_sample_0356.ext - technology: sky130A

.subckt diff_pair_sample_0356 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=0.51
X1 VTAIL.t16 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X2 VDD2.t9 VN.t0 VTAIL.t19 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=0.51
X4 VDD1.t4 VP.t1 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X5 VTAIL.t14 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=0.51
X7 VDD1.t1 VP.t3 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=3.0954 ps=19.09 w=18.76 l=0.51
X8 VTAIL.t12 VP.t4 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X9 VTAIL.t3 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X10 VDD2.t7 VN.t2 VTAIL.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=3.0954 ps=19.09 w=18.76 l=0.51
X11 VDD1.t0 VP.t5 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=3.0954 ps=19.09 w=18.76 l=0.51
X12 VDD1.t9 VP.t6 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=7.3164 ps=38.3 w=18.76 l=0.51
X13 VTAIL.t5 VN.t3 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X14 VDD2.t5 VN.t4 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=7.3164 ps=38.3 w=18.76 l=0.51
X15 VDD2.t4 VN.t5 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=3.0954 ps=19.09 w=18.76 l=0.51
X16 VDD2.t3 VN.t6 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X17 VTAIL.t9 VP.t7 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X18 VTAIL.t17 VN.t7 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X19 VTAIL.t6 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
X20 VDD1.t8 VP.t8 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=7.3164 ps=38.3 w=18.76 l=0.51
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=0.51
X22 VDD2.t0 VN.t9 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=7.3164 ps=38.3 w=18.76 l=0.51
X23 VDD1.t5 VP.t9 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0954 pd=19.09 as=3.0954 ps=19.09 w=18.76 l=0.51
R0 B.n490 B.t14 1092.67
R1 B.n488 B.t18 1092.67
R2 B.n116 B.t10 1092.67
R3 B.n114 B.t21 1092.67
R4 B.n860 B.n859 585
R5 B.n861 B.n860 585
R6 B.n378 B.n112 585
R7 B.n377 B.n376 585
R8 B.n375 B.n374 585
R9 B.n373 B.n372 585
R10 B.n371 B.n370 585
R11 B.n369 B.n368 585
R12 B.n367 B.n366 585
R13 B.n365 B.n364 585
R14 B.n363 B.n362 585
R15 B.n361 B.n360 585
R16 B.n359 B.n358 585
R17 B.n357 B.n356 585
R18 B.n355 B.n354 585
R19 B.n353 B.n352 585
R20 B.n351 B.n350 585
R21 B.n349 B.n348 585
R22 B.n347 B.n346 585
R23 B.n345 B.n344 585
R24 B.n343 B.n342 585
R25 B.n341 B.n340 585
R26 B.n339 B.n338 585
R27 B.n337 B.n336 585
R28 B.n335 B.n334 585
R29 B.n333 B.n332 585
R30 B.n331 B.n330 585
R31 B.n329 B.n328 585
R32 B.n327 B.n326 585
R33 B.n325 B.n324 585
R34 B.n323 B.n322 585
R35 B.n321 B.n320 585
R36 B.n319 B.n318 585
R37 B.n317 B.n316 585
R38 B.n315 B.n314 585
R39 B.n313 B.n312 585
R40 B.n311 B.n310 585
R41 B.n309 B.n308 585
R42 B.n307 B.n306 585
R43 B.n305 B.n304 585
R44 B.n303 B.n302 585
R45 B.n301 B.n300 585
R46 B.n299 B.n298 585
R47 B.n297 B.n296 585
R48 B.n295 B.n294 585
R49 B.n293 B.n292 585
R50 B.n291 B.n290 585
R51 B.n289 B.n288 585
R52 B.n287 B.n286 585
R53 B.n285 B.n284 585
R54 B.n283 B.n282 585
R55 B.n281 B.n280 585
R56 B.n279 B.n278 585
R57 B.n277 B.n276 585
R58 B.n275 B.n274 585
R59 B.n273 B.n272 585
R60 B.n271 B.n270 585
R61 B.n269 B.n268 585
R62 B.n267 B.n266 585
R63 B.n265 B.n264 585
R64 B.n263 B.n262 585
R65 B.n261 B.n260 585
R66 B.n259 B.n258 585
R67 B.n256 B.n255 585
R68 B.n254 B.n253 585
R69 B.n252 B.n251 585
R70 B.n250 B.n249 585
R71 B.n248 B.n247 585
R72 B.n246 B.n245 585
R73 B.n244 B.n243 585
R74 B.n242 B.n241 585
R75 B.n240 B.n239 585
R76 B.n238 B.n237 585
R77 B.n236 B.n235 585
R78 B.n234 B.n233 585
R79 B.n232 B.n231 585
R80 B.n230 B.n229 585
R81 B.n228 B.n227 585
R82 B.n226 B.n225 585
R83 B.n224 B.n223 585
R84 B.n222 B.n221 585
R85 B.n220 B.n219 585
R86 B.n218 B.n217 585
R87 B.n216 B.n215 585
R88 B.n214 B.n213 585
R89 B.n212 B.n211 585
R90 B.n210 B.n209 585
R91 B.n208 B.n207 585
R92 B.n206 B.n205 585
R93 B.n204 B.n203 585
R94 B.n202 B.n201 585
R95 B.n200 B.n199 585
R96 B.n198 B.n197 585
R97 B.n196 B.n195 585
R98 B.n194 B.n193 585
R99 B.n192 B.n191 585
R100 B.n190 B.n189 585
R101 B.n188 B.n187 585
R102 B.n186 B.n185 585
R103 B.n184 B.n183 585
R104 B.n182 B.n181 585
R105 B.n180 B.n179 585
R106 B.n178 B.n177 585
R107 B.n176 B.n175 585
R108 B.n174 B.n173 585
R109 B.n172 B.n171 585
R110 B.n170 B.n169 585
R111 B.n168 B.n167 585
R112 B.n166 B.n165 585
R113 B.n164 B.n163 585
R114 B.n162 B.n161 585
R115 B.n160 B.n159 585
R116 B.n158 B.n157 585
R117 B.n156 B.n155 585
R118 B.n154 B.n153 585
R119 B.n152 B.n151 585
R120 B.n150 B.n149 585
R121 B.n148 B.n147 585
R122 B.n146 B.n145 585
R123 B.n144 B.n143 585
R124 B.n142 B.n141 585
R125 B.n140 B.n139 585
R126 B.n138 B.n137 585
R127 B.n136 B.n135 585
R128 B.n134 B.n133 585
R129 B.n132 B.n131 585
R130 B.n130 B.n129 585
R131 B.n128 B.n127 585
R132 B.n126 B.n125 585
R133 B.n124 B.n123 585
R134 B.n122 B.n121 585
R135 B.n120 B.n119 585
R136 B.n46 B.n45 585
R137 B.n864 B.n863 585
R138 B.n858 B.n113 585
R139 B.n113 B.n43 585
R140 B.n857 B.n42 585
R141 B.n868 B.n42 585
R142 B.n856 B.n41 585
R143 B.n869 B.n41 585
R144 B.n855 B.n40 585
R145 B.n870 B.n40 585
R146 B.n854 B.n853 585
R147 B.n853 B.n39 585
R148 B.n852 B.n35 585
R149 B.n876 B.n35 585
R150 B.n851 B.n34 585
R151 B.n877 B.n34 585
R152 B.n850 B.n33 585
R153 B.n878 B.n33 585
R154 B.n849 B.n848 585
R155 B.n848 B.n29 585
R156 B.n847 B.n28 585
R157 B.n884 B.n28 585
R158 B.n846 B.n27 585
R159 B.n885 B.n27 585
R160 B.n845 B.n26 585
R161 B.n886 B.n26 585
R162 B.n844 B.n843 585
R163 B.n843 B.n25 585
R164 B.n842 B.n21 585
R165 B.n892 B.n21 585
R166 B.n841 B.n20 585
R167 B.n893 B.n20 585
R168 B.n840 B.n19 585
R169 B.n894 B.n19 585
R170 B.n839 B.n838 585
R171 B.n838 B.n15 585
R172 B.n837 B.n14 585
R173 B.n900 B.n14 585
R174 B.n836 B.n13 585
R175 B.n901 B.n13 585
R176 B.n835 B.n12 585
R177 B.n902 B.n12 585
R178 B.n834 B.n833 585
R179 B.n833 B.n11 585
R180 B.n832 B.n7 585
R181 B.n908 B.n7 585
R182 B.n831 B.n6 585
R183 B.n909 B.n6 585
R184 B.n830 B.n5 585
R185 B.n910 B.n5 585
R186 B.n829 B.n828 585
R187 B.n828 B.n4 585
R188 B.n827 B.n379 585
R189 B.n827 B.n826 585
R190 B.n816 B.n380 585
R191 B.n819 B.n380 585
R192 B.n818 B.n817 585
R193 B.n820 B.n818 585
R194 B.n815 B.n385 585
R195 B.n385 B.n384 585
R196 B.n814 B.n813 585
R197 B.n813 B.n812 585
R198 B.n387 B.n386 585
R199 B.n388 B.n387 585
R200 B.n805 B.n804 585
R201 B.n806 B.n805 585
R202 B.n803 B.n393 585
R203 B.n393 B.n392 585
R204 B.n802 B.n801 585
R205 B.n801 B.n800 585
R206 B.n395 B.n394 585
R207 B.n793 B.n395 585
R208 B.n792 B.n791 585
R209 B.n794 B.n792 585
R210 B.n790 B.n399 585
R211 B.n403 B.n399 585
R212 B.n789 B.n788 585
R213 B.n788 B.n787 585
R214 B.n401 B.n400 585
R215 B.n402 B.n401 585
R216 B.n780 B.n779 585
R217 B.n781 B.n780 585
R218 B.n778 B.n408 585
R219 B.n408 B.n407 585
R220 B.n777 B.n776 585
R221 B.n776 B.n775 585
R222 B.n410 B.n409 585
R223 B.n768 B.n410 585
R224 B.n767 B.n766 585
R225 B.n769 B.n767 585
R226 B.n765 B.n415 585
R227 B.n415 B.n414 585
R228 B.n764 B.n763 585
R229 B.n763 B.n762 585
R230 B.n417 B.n416 585
R231 B.n418 B.n417 585
R232 B.n758 B.n757 585
R233 B.n421 B.n420 585
R234 B.n754 B.n753 585
R235 B.n755 B.n754 585
R236 B.n752 B.n487 585
R237 B.n751 B.n750 585
R238 B.n749 B.n748 585
R239 B.n747 B.n746 585
R240 B.n745 B.n744 585
R241 B.n743 B.n742 585
R242 B.n741 B.n740 585
R243 B.n739 B.n738 585
R244 B.n737 B.n736 585
R245 B.n735 B.n734 585
R246 B.n733 B.n732 585
R247 B.n731 B.n730 585
R248 B.n729 B.n728 585
R249 B.n727 B.n726 585
R250 B.n725 B.n724 585
R251 B.n723 B.n722 585
R252 B.n721 B.n720 585
R253 B.n719 B.n718 585
R254 B.n717 B.n716 585
R255 B.n715 B.n714 585
R256 B.n713 B.n712 585
R257 B.n711 B.n710 585
R258 B.n709 B.n708 585
R259 B.n707 B.n706 585
R260 B.n705 B.n704 585
R261 B.n703 B.n702 585
R262 B.n701 B.n700 585
R263 B.n699 B.n698 585
R264 B.n697 B.n696 585
R265 B.n695 B.n694 585
R266 B.n693 B.n692 585
R267 B.n691 B.n690 585
R268 B.n689 B.n688 585
R269 B.n687 B.n686 585
R270 B.n685 B.n684 585
R271 B.n683 B.n682 585
R272 B.n681 B.n680 585
R273 B.n679 B.n678 585
R274 B.n677 B.n676 585
R275 B.n675 B.n674 585
R276 B.n673 B.n672 585
R277 B.n671 B.n670 585
R278 B.n669 B.n668 585
R279 B.n667 B.n666 585
R280 B.n665 B.n664 585
R281 B.n663 B.n662 585
R282 B.n661 B.n660 585
R283 B.n659 B.n658 585
R284 B.n657 B.n656 585
R285 B.n655 B.n654 585
R286 B.n653 B.n652 585
R287 B.n651 B.n650 585
R288 B.n649 B.n648 585
R289 B.n647 B.n646 585
R290 B.n645 B.n644 585
R291 B.n643 B.n642 585
R292 B.n641 B.n640 585
R293 B.n639 B.n638 585
R294 B.n637 B.n636 585
R295 B.n634 B.n633 585
R296 B.n632 B.n631 585
R297 B.n630 B.n629 585
R298 B.n628 B.n627 585
R299 B.n626 B.n625 585
R300 B.n624 B.n623 585
R301 B.n622 B.n621 585
R302 B.n620 B.n619 585
R303 B.n618 B.n617 585
R304 B.n616 B.n615 585
R305 B.n614 B.n613 585
R306 B.n612 B.n611 585
R307 B.n610 B.n609 585
R308 B.n608 B.n607 585
R309 B.n606 B.n605 585
R310 B.n604 B.n603 585
R311 B.n602 B.n601 585
R312 B.n600 B.n599 585
R313 B.n598 B.n597 585
R314 B.n596 B.n595 585
R315 B.n594 B.n593 585
R316 B.n592 B.n591 585
R317 B.n590 B.n589 585
R318 B.n588 B.n587 585
R319 B.n586 B.n585 585
R320 B.n584 B.n583 585
R321 B.n582 B.n581 585
R322 B.n580 B.n579 585
R323 B.n578 B.n577 585
R324 B.n576 B.n575 585
R325 B.n574 B.n573 585
R326 B.n572 B.n571 585
R327 B.n570 B.n569 585
R328 B.n568 B.n567 585
R329 B.n566 B.n565 585
R330 B.n564 B.n563 585
R331 B.n562 B.n561 585
R332 B.n560 B.n559 585
R333 B.n558 B.n557 585
R334 B.n556 B.n555 585
R335 B.n554 B.n553 585
R336 B.n552 B.n551 585
R337 B.n550 B.n549 585
R338 B.n548 B.n547 585
R339 B.n546 B.n545 585
R340 B.n544 B.n543 585
R341 B.n542 B.n541 585
R342 B.n540 B.n539 585
R343 B.n538 B.n537 585
R344 B.n536 B.n535 585
R345 B.n534 B.n533 585
R346 B.n532 B.n531 585
R347 B.n530 B.n529 585
R348 B.n528 B.n527 585
R349 B.n526 B.n525 585
R350 B.n524 B.n523 585
R351 B.n522 B.n521 585
R352 B.n520 B.n519 585
R353 B.n518 B.n517 585
R354 B.n516 B.n515 585
R355 B.n514 B.n513 585
R356 B.n512 B.n511 585
R357 B.n510 B.n509 585
R358 B.n508 B.n507 585
R359 B.n506 B.n505 585
R360 B.n504 B.n503 585
R361 B.n502 B.n501 585
R362 B.n500 B.n499 585
R363 B.n498 B.n497 585
R364 B.n496 B.n495 585
R365 B.n494 B.n493 585
R366 B.n759 B.n419 585
R367 B.n419 B.n418 585
R368 B.n761 B.n760 585
R369 B.n762 B.n761 585
R370 B.n413 B.n412 585
R371 B.n414 B.n413 585
R372 B.n771 B.n770 585
R373 B.n770 B.n769 585
R374 B.n772 B.n411 585
R375 B.n768 B.n411 585
R376 B.n774 B.n773 585
R377 B.n775 B.n774 585
R378 B.n406 B.n405 585
R379 B.n407 B.n406 585
R380 B.n783 B.n782 585
R381 B.n782 B.n781 585
R382 B.n784 B.n404 585
R383 B.n404 B.n402 585
R384 B.n786 B.n785 585
R385 B.n787 B.n786 585
R386 B.n398 B.n397 585
R387 B.n403 B.n398 585
R388 B.n796 B.n795 585
R389 B.n795 B.n794 585
R390 B.n797 B.n396 585
R391 B.n793 B.n396 585
R392 B.n799 B.n798 585
R393 B.n800 B.n799 585
R394 B.n391 B.n390 585
R395 B.n392 B.n391 585
R396 B.n808 B.n807 585
R397 B.n807 B.n806 585
R398 B.n809 B.n389 585
R399 B.n389 B.n388 585
R400 B.n811 B.n810 585
R401 B.n812 B.n811 585
R402 B.n383 B.n382 585
R403 B.n384 B.n383 585
R404 B.n822 B.n821 585
R405 B.n821 B.n820 585
R406 B.n823 B.n381 585
R407 B.n819 B.n381 585
R408 B.n825 B.n824 585
R409 B.n826 B.n825 585
R410 B.n2 B.n0 585
R411 B.n4 B.n2 585
R412 B.n3 B.n1 585
R413 B.n909 B.n3 585
R414 B.n907 B.n906 585
R415 B.n908 B.n907 585
R416 B.n905 B.n8 585
R417 B.n11 B.n8 585
R418 B.n904 B.n903 585
R419 B.n903 B.n902 585
R420 B.n10 B.n9 585
R421 B.n901 B.n10 585
R422 B.n899 B.n898 585
R423 B.n900 B.n899 585
R424 B.n897 B.n16 585
R425 B.n16 B.n15 585
R426 B.n896 B.n895 585
R427 B.n895 B.n894 585
R428 B.n18 B.n17 585
R429 B.n893 B.n18 585
R430 B.n891 B.n890 585
R431 B.n892 B.n891 585
R432 B.n889 B.n22 585
R433 B.n25 B.n22 585
R434 B.n888 B.n887 585
R435 B.n887 B.n886 585
R436 B.n24 B.n23 585
R437 B.n885 B.n24 585
R438 B.n883 B.n882 585
R439 B.n884 B.n883 585
R440 B.n881 B.n30 585
R441 B.n30 B.n29 585
R442 B.n880 B.n879 585
R443 B.n879 B.n878 585
R444 B.n32 B.n31 585
R445 B.n877 B.n32 585
R446 B.n875 B.n874 585
R447 B.n876 B.n875 585
R448 B.n873 B.n36 585
R449 B.n39 B.n36 585
R450 B.n872 B.n871 585
R451 B.n871 B.n870 585
R452 B.n38 B.n37 585
R453 B.n869 B.n38 585
R454 B.n867 B.n866 585
R455 B.n868 B.n867 585
R456 B.n865 B.n44 585
R457 B.n44 B.n43 585
R458 B.n912 B.n911 585
R459 B.n911 B.n910 585
R460 B.n757 B.n419 454.062
R461 B.n863 B.n44 454.062
R462 B.n493 B.n417 454.062
R463 B.n860 B.n113 454.062
R464 B.n490 B.t17 414.647
R465 B.n114 B.t22 414.647
R466 B.n488 B.t20 414.647
R467 B.n116 B.t12 414.647
R468 B.n491 B.t16 398.356
R469 B.n115 B.t23 398.356
R470 B.n489 B.t19 398.356
R471 B.n117 B.t13 398.356
R472 B.n861 B.n111 256.663
R473 B.n861 B.n110 256.663
R474 B.n861 B.n109 256.663
R475 B.n861 B.n108 256.663
R476 B.n861 B.n107 256.663
R477 B.n861 B.n106 256.663
R478 B.n861 B.n105 256.663
R479 B.n861 B.n104 256.663
R480 B.n861 B.n103 256.663
R481 B.n861 B.n102 256.663
R482 B.n861 B.n101 256.663
R483 B.n861 B.n100 256.663
R484 B.n861 B.n99 256.663
R485 B.n861 B.n98 256.663
R486 B.n861 B.n97 256.663
R487 B.n861 B.n96 256.663
R488 B.n861 B.n95 256.663
R489 B.n861 B.n94 256.663
R490 B.n861 B.n93 256.663
R491 B.n861 B.n92 256.663
R492 B.n861 B.n91 256.663
R493 B.n861 B.n90 256.663
R494 B.n861 B.n89 256.663
R495 B.n861 B.n88 256.663
R496 B.n861 B.n87 256.663
R497 B.n861 B.n86 256.663
R498 B.n861 B.n85 256.663
R499 B.n861 B.n84 256.663
R500 B.n861 B.n83 256.663
R501 B.n861 B.n82 256.663
R502 B.n861 B.n81 256.663
R503 B.n861 B.n80 256.663
R504 B.n861 B.n79 256.663
R505 B.n861 B.n78 256.663
R506 B.n861 B.n77 256.663
R507 B.n861 B.n76 256.663
R508 B.n861 B.n75 256.663
R509 B.n861 B.n74 256.663
R510 B.n861 B.n73 256.663
R511 B.n861 B.n72 256.663
R512 B.n861 B.n71 256.663
R513 B.n861 B.n70 256.663
R514 B.n861 B.n69 256.663
R515 B.n861 B.n68 256.663
R516 B.n861 B.n67 256.663
R517 B.n861 B.n66 256.663
R518 B.n861 B.n65 256.663
R519 B.n861 B.n64 256.663
R520 B.n861 B.n63 256.663
R521 B.n861 B.n62 256.663
R522 B.n861 B.n61 256.663
R523 B.n861 B.n60 256.663
R524 B.n861 B.n59 256.663
R525 B.n861 B.n58 256.663
R526 B.n861 B.n57 256.663
R527 B.n861 B.n56 256.663
R528 B.n861 B.n55 256.663
R529 B.n861 B.n54 256.663
R530 B.n861 B.n53 256.663
R531 B.n861 B.n52 256.663
R532 B.n861 B.n51 256.663
R533 B.n861 B.n50 256.663
R534 B.n861 B.n49 256.663
R535 B.n861 B.n48 256.663
R536 B.n861 B.n47 256.663
R537 B.n862 B.n861 256.663
R538 B.n756 B.n755 256.663
R539 B.n755 B.n422 256.663
R540 B.n755 B.n423 256.663
R541 B.n755 B.n424 256.663
R542 B.n755 B.n425 256.663
R543 B.n755 B.n426 256.663
R544 B.n755 B.n427 256.663
R545 B.n755 B.n428 256.663
R546 B.n755 B.n429 256.663
R547 B.n755 B.n430 256.663
R548 B.n755 B.n431 256.663
R549 B.n755 B.n432 256.663
R550 B.n755 B.n433 256.663
R551 B.n755 B.n434 256.663
R552 B.n755 B.n435 256.663
R553 B.n755 B.n436 256.663
R554 B.n755 B.n437 256.663
R555 B.n755 B.n438 256.663
R556 B.n755 B.n439 256.663
R557 B.n755 B.n440 256.663
R558 B.n755 B.n441 256.663
R559 B.n755 B.n442 256.663
R560 B.n755 B.n443 256.663
R561 B.n755 B.n444 256.663
R562 B.n755 B.n445 256.663
R563 B.n755 B.n446 256.663
R564 B.n755 B.n447 256.663
R565 B.n755 B.n448 256.663
R566 B.n755 B.n449 256.663
R567 B.n755 B.n450 256.663
R568 B.n755 B.n451 256.663
R569 B.n755 B.n452 256.663
R570 B.n755 B.n453 256.663
R571 B.n755 B.n454 256.663
R572 B.n755 B.n455 256.663
R573 B.n755 B.n456 256.663
R574 B.n755 B.n457 256.663
R575 B.n755 B.n458 256.663
R576 B.n755 B.n459 256.663
R577 B.n755 B.n460 256.663
R578 B.n755 B.n461 256.663
R579 B.n755 B.n462 256.663
R580 B.n755 B.n463 256.663
R581 B.n755 B.n464 256.663
R582 B.n755 B.n465 256.663
R583 B.n755 B.n466 256.663
R584 B.n755 B.n467 256.663
R585 B.n755 B.n468 256.663
R586 B.n755 B.n469 256.663
R587 B.n755 B.n470 256.663
R588 B.n755 B.n471 256.663
R589 B.n755 B.n472 256.663
R590 B.n755 B.n473 256.663
R591 B.n755 B.n474 256.663
R592 B.n755 B.n475 256.663
R593 B.n755 B.n476 256.663
R594 B.n755 B.n477 256.663
R595 B.n755 B.n478 256.663
R596 B.n755 B.n479 256.663
R597 B.n755 B.n480 256.663
R598 B.n755 B.n481 256.663
R599 B.n755 B.n482 256.663
R600 B.n755 B.n483 256.663
R601 B.n755 B.n484 256.663
R602 B.n755 B.n485 256.663
R603 B.n755 B.n486 256.663
R604 B.n761 B.n419 163.367
R605 B.n761 B.n413 163.367
R606 B.n770 B.n413 163.367
R607 B.n770 B.n411 163.367
R608 B.n774 B.n411 163.367
R609 B.n774 B.n406 163.367
R610 B.n782 B.n406 163.367
R611 B.n782 B.n404 163.367
R612 B.n786 B.n404 163.367
R613 B.n786 B.n398 163.367
R614 B.n795 B.n398 163.367
R615 B.n795 B.n396 163.367
R616 B.n799 B.n396 163.367
R617 B.n799 B.n391 163.367
R618 B.n807 B.n391 163.367
R619 B.n807 B.n389 163.367
R620 B.n811 B.n389 163.367
R621 B.n811 B.n383 163.367
R622 B.n821 B.n383 163.367
R623 B.n821 B.n381 163.367
R624 B.n825 B.n381 163.367
R625 B.n825 B.n2 163.367
R626 B.n911 B.n2 163.367
R627 B.n911 B.n3 163.367
R628 B.n907 B.n3 163.367
R629 B.n907 B.n8 163.367
R630 B.n903 B.n8 163.367
R631 B.n903 B.n10 163.367
R632 B.n899 B.n10 163.367
R633 B.n899 B.n16 163.367
R634 B.n895 B.n16 163.367
R635 B.n895 B.n18 163.367
R636 B.n891 B.n18 163.367
R637 B.n891 B.n22 163.367
R638 B.n887 B.n22 163.367
R639 B.n887 B.n24 163.367
R640 B.n883 B.n24 163.367
R641 B.n883 B.n30 163.367
R642 B.n879 B.n30 163.367
R643 B.n879 B.n32 163.367
R644 B.n875 B.n32 163.367
R645 B.n875 B.n36 163.367
R646 B.n871 B.n36 163.367
R647 B.n871 B.n38 163.367
R648 B.n867 B.n38 163.367
R649 B.n867 B.n44 163.367
R650 B.n754 B.n421 163.367
R651 B.n754 B.n487 163.367
R652 B.n750 B.n749 163.367
R653 B.n746 B.n745 163.367
R654 B.n742 B.n741 163.367
R655 B.n738 B.n737 163.367
R656 B.n734 B.n733 163.367
R657 B.n730 B.n729 163.367
R658 B.n726 B.n725 163.367
R659 B.n722 B.n721 163.367
R660 B.n718 B.n717 163.367
R661 B.n714 B.n713 163.367
R662 B.n710 B.n709 163.367
R663 B.n706 B.n705 163.367
R664 B.n702 B.n701 163.367
R665 B.n698 B.n697 163.367
R666 B.n694 B.n693 163.367
R667 B.n690 B.n689 163.367
R668 B.n686 B.n685 163.367
R669 B.n682 B.n681 163.367
R670 B.n678 B.n677 163.367
R671 B.n674 B.n673 163.367
R672 B.n670 B.n669 163.367
R673 B.n666 B.n665 163.367
R674 B.n662 B.n661 163.367
R675 B.n658 B.n657 163.367
R676 B.n654 B.n653 163.367
R677 B.n650 B.n649 163.367
R678 B.n646 B.n645 163.367
R679 B.n642 B.n641 163.367
R680 B.n638 B.n637 163.367
R681 B.n633 B.n632 163.367
R682 B.n629 B.n628 163.367
R683 B.n625 B.n624 163.367
R684 B.n621 B.n620 163.367
R685 B.n617 B.n616 163.367
R686 B.n613 B.n612 163.367
R687 B.n609 B.n608 163.367
R688 B.n605 B.n604 163.367
R689 B.n601 B.n600 163.367
R690 B.n597 B.n596 163.367
R691 B.n593 B.n592 163.367
R692 B.n589 B.n588 163.367
R693 B.n585 B.n584 163.367
R694 B.n581 B.n580 163.367
R695 B.n577 B.n576 163.367
R696 B.n573 B.n572 163.367
R697 B.n569 B.n568 163.367
R698 B.n565 B.n564 163.367
R699 B.n561 B.n560 163.367
R700 B.n557 B.n556 163.367
R701 B.n553 B.n552 163.367
R702 B.n549 B.n548 163.367
R703 B.n545 B.n544 163.367
R704 B.n541 B.n540 163.367
R705 B.n537 B.n536 163.367
R706 B.n533 B.n532 163.367
R707 B.n529 B.n528 163.367
R708 B.n525 B.n524 163.367
R709 B.n521 B.n520 163.367
R710 B.n517 B.n516 163.367
R711 B.n513 B.n512 163.367
R712 B.n509 B.n508 163.367
R713 B.n505 B.n504 163.367
R714 B.n501 B.n500 163.367
R715 B.n497 B.n496 163.367
R716 B.n763 B.n417 163.367
R717 B.n763 B.n415 163.367
R718 B.n767 B.n415 163.367
R719 B.n767 B.n410 163.367
R720 B.n776 B.n410 163.367
R721 B.n776 B.n408 163.367
R722 B.n780 B.n408 163.367
R723 B.n780 B.n401 163.367
R724 B.n788 B.n401 163.367
R725 B.n788 B.n399 163.367
R726 B.n792 B.n399 163.367
R727 B.n792 B.n395 163.367
R728 B.n801 B.n395 163.367
R729 B.n801 B.n393 163.367
R730 B.n805 B.n393 163.367
R731 B.n805 B.n387 163.367
R732 B.n813 B.n387 163.367
R733 B.n813 B.n385 163.367
R734 B.n818 B.n385 163.367
R735 B.n818 B.n380 163.367
R736 B.n827 B.n380 163.367
R737 B.n828 B.n827 163.367
R738 B.n828 B.n5 163.367
R739 B.n6 B.n5 163.367
R740 B.n7 B.n6 163.367
R741 B.n833 B.n7 163.367
R742 B.n833 B.n12 163.367
R743 B.n13 B.n12 163.367
R744 B.n14 B.n13 163.367
R745 B.n838 B.n14 163.367
R746 B.n838 B.n19 163.367
R747 B.n20 B.n19 163.367
R748 B.n21 B.n20 163.367
R749 B.n843 B.n21 163.367
R750 B.n843 B.n26 163.367
R751 B.n27 B.n26 163.367
R752 B.n28 B.n27 163.367
R753 B.n848 B.n28 163.367
R754 B.n848 B.n33 163.367
R755 B.n34 B.n33 163.367
R756 B.n35 B.n34 163.367
R757 B.n853 B.n35 163.367
R758 B.n853 B.n40 163.367
R759 B.n41 B.n40 163.367
R760 B.n42 B.n41 163.367
R761 B.n113 B.n42 163.367
R762 B.n119 B.n46 163.367
R763 B.n123 B.n122 163.367
R764 B.n127 B.n126 163.367
R765 B.n131 B.n130 163.367
R766 B.n135 B.n134 163.367
R767 B.n139 B.n138 163.367
R768 B.n143 B.n142 163.367
R769 B.n147 B.n146 163.367
R770 B.n151 B.n150 163.367
R771 B.n155 B.n154 163.367
R772 B.n159 B.n158 163.367
R773 B.n163 B.n162 163.367
R774 B.n167 B.n166 163.367
R775 B.n171 B.n170 163.367
R776 B.n175 B.n174 163.367
R777 B.n179 B.n178 163.367
R778 B.n183 B.n182 163.367
R779 B.n187 B.n186 163.367
R780 B.n191 B.n190 163.367
R781 B.n195 B.n194 163.367
R782 B.n199 B.n198 163.367
R783 B.n203 B.n202 163.367
R784 B.n207 B.n206 163.367
R785 B.n211 B.n210 163.367
R786 B.n215 B.n214 163.367
R787 B.n219 B.n218 163.367
R788 B.n223 B.n222 163.367
R789 B.n227 B.n226 163.367
R790 B.n231 B.n230 163.367
R791 B.n235 B.n234 163.367
R792 B.n239 B.n238 163.367
R793 B.n243 B.n242 163.367
R794 B.n247 B.n246 163.367
R795 B.n251 B.n250 163.367
R796 B.n255 B.n254 163.367
R797 B.n260 B.n259 163.367
R798 B.n264 B.n263 163.367
R799 B.n268 B.n267 163.367
R800 B.n272 B.n271 163.367
R801 B.n276 B.n275 163.367
R802 B.n280 B.n279 163.367
R803 B.n284 B.n283 163.367
R804 B.n288 B.n287 163.367
R805 B.n292 B.n291 163.367
R806 B.n296 B.n295 163.367
R807 B.n300 B.n299 163.367
R808 B.n304 B.n303 163.367
R809 B.n308 B.n307 163.367
R810 B.n312 B.n311 163.367
R811 B.n316 B.n315 163.367
R812 B.n320 B.n319 163.367
R813 B.n324 B.n323 163.367
R814 B.n328 B.n327 163.367
R815 B.n332 B.n331 163.367
R816 B.n336 B.n335 163.367
R817 B.n340 B.n339 163.367
R818 B.n344 B.n343 163.367
R819 B.n348 B.n347 163.367
R820 B.n352 B.n351 163.367
R821 B.n356 B.n355 163.367
R822 B.n360 B.n359 163.367
R823 B.n364 B.n363 163.367
R824 B.n368 B.n367 163.367
R825 B.n372 B.n371 163.367
R826 B.n376 B.n375 163.367
R827 B.n860 B.n112 163.367
R828 B.n757 B.n756 71.676
R829 B.n487 B.n422 71.676
R830 B.n749 B.n423 71.676
R831 B.n745 B.n424 71.676
R832 B.n741 B.n425 71.676
R833 B.n737 B.n426 71.676
R834 B.n733 B.n427 71.676
R835 B.n729 B.n428 71.676
R836 B.n725 B.n429 71.676
R837 B.n721 B.n430 71.676
R838 B.n717 B.n431 71.676
R839 B.n713 B.n432 71.676
R840 B.n709 B.n433 71.676
R841 B.n705 B.n434 71.676
R842 B.n701 B.n435 71.676
R843 B.n697 B.n436 71.676
R844 B.n693 B.n437 71.676
R845 B.n689 B.n438 71.676
R846 B.n685 B.n439 71.676
R847 B.n681 B.n440 71.676
R848 B.n677 B.n441 71.676
R849 B.n673 B.n442 71.676
R850 B.n669 B.n443 71.676
R851 B.n665 B.n444 71.676
R852 B.n661 B.n445 71.676
R853 B.n657 B.n446 71.676
R854 B.n653 B.n447 71.676
R855 B.n649 B.n448 71.676
R856 B.n645 B.n449 71.676
R857 B.n641 B.n450 71.676
R858 B.n637 B.n451 71.676
R859 B.n632 B.n452 71.676
R860 B.n628 B.n453 71.676
R861 B.n624 B.n454 71.676
R862 B.n620 B.n455 71.676
R863 B.n616 B.n456 71.676
R864 B.n612 B.n457 71.676
R865 B.n608 B.n458 71.676
R866 B.n604 B.n459 71.676
R867 B.n600 B.n460 71.676
R868 B.n596 B.n461 71.676
R869 B.n592 B.n462 71.676
R870 B.n588 B.n463 71.676
R871 B.n584 B.n464 71.676
R872 B.n580 B.n465 71.676
R873 B.n576 B.n466 71.676
R874 B.n572 B.n467 71.676
R875 B.n568 B.n468 71.676
R876 B.n564 B.n469 71.676
R877 B.n560 B.n470 71.676
R878 B.n556 B.n471 71.676
R879 B.n552 B.n472 71.676
R880 B.n548 B.n473 71.676
R881 B.n544 B.n474 71.676
R882 B.n540 B.n475 71.676
R883 B.n536 B.n476 71.676
R884 B.n532 B.n477 71.676
R885 B.n528 B.n478 71.676
R886 B.n524 B.n479 71.676
R887 B.n520 B.n480 71.676
R888 B.n516 B.n481 71.676
R889 B.n512 B.n482 71.676
R890 B.n508 B.n483 71.676
R891 B.n504 B.n484 71.676
R892 B.n500 B.n485 71.676
R893 B.n496 B.n486 71.676
R894 B.n863 B.n862 71.676
R895 B.n119 B.n47 71.676
R896 B.n123 B.n48 71.676
R897 B.n127 B.n49 71.676
R898 B.n131 B.n50 71.676
R899 B.n135 B.n51 71.676
R900 B.n139 B.n52 71.676
R901 B.n143 B.n53 71.676
R902 B.n147 B.n54 71.676
R903 B.n151 B.n55 71.676
R904 B.n155 B.n56 71.676
R905 B.n159 B.n57 71.676
R906 B.n163 B.n58 71.676
R907 B.n167 B.n59 71.676
R908 B.n171 B.n60 71.676
R909 B.n175 B.n61 71.676
R910 B.n179 B.n62 71.676
R911 B.n183 B.n63 71.676
R912 B.n187 B.n64 71.676
R913 B.n191 B.n65 71.676
R914 B.n195 B.n66 71.676
R915 B.n199 B.n67 71.676
R916 B.n203 B.n68 71.676
R917 B.n207 B.n69 71.676
R918 B.n211 B.n70 71.676
R919 B.n215 B.n71 71.676
R920 B.n219 B.n72 71.676
R921 B.n223 B.n73 71.676
R922 B.n227 B.n74 71.676
R923 B.n231 B.n75 71.676
R924 B.n235 B.n76 71.676
R925 B.n239 B.n77 71.676
R926 B.n243 B.n78 71.676
R927 B.n247 B.n79 71.676
R928 B.n251 B.n80 71.676
R929 B.n255 B.n81 71.676
R930 B.n260 B.n82 71.676
R931 B.n264 B.n83 71.676
R932 B.n268 B.n84 71.676
R933 B.n272 B.n85 71.676
R934 B.n276 B.n86 71.676
R935 B.n280 B.n87 71.676
R936 B.n284 B.n88 71.676
R937 B.n288 B.n89 71.676
R938 B.n292 B.n90 71.676
R939 B.n296 B.n91 71.676
R940 B.n300 B.n92 71.676
R941 B.n304 B.n93 71.676
R942 B.n308 B.n94 71.676
R943 B.n312 B.n95 71.676
R944 B.n316 B.n96 71.676
R945 B.n320 B.n97 71.676
R946 B.n324 B.n98 71.676
R947 B.n328 B.n99 71.676
R948 B.n332 B.n100 71.676
R949 B.n336 B.n101 71.676
R950 B.n340 B.n102 71.676
R951 B.n344 B.n103 71.676
R952 B.n348 B.n104 71.676
R953 B.n352 B.n105 71.676
R954 B.n356 B.n106 71.676
R955 B.n360 B.n107 71.676
R956 B.n364 B.n108 71.676
R957 B.n368 B.n109 71.676
R958 B.n372 B.n110 71.676
R959 B.n376 B.n111 71.676
R960 B.n112 B.n111 71.676
R961 B.n375 B.n110 71.676
R962 B.n371 B.n109 71.676
R963 B.n367 B.n108 71.676
R964 B.n363 B.n107 71.676
R965 B.n359 B.n106 71.676
R966 B.n355 B.n105 71.676
R967 B.n351 B.n104 71.676
R968 B.n347 B.n103 71.676
R969 B.n343 B.n102 71.676
R970 B.n339 B.n101 71.676
R971 B.n335 B.n100 71.676
R972 B.n331 B.n99 71.676
R973 B.n327 B.n98 71.676
R974 B.n323 B.n97 71.676
R975 B.n319 B.n96 71.676
R976 B.n315 B.n95 71.676
R977 B.n311 B.n94 71.676
R978 B.n307 B.n93 71.676
R979 B.n303 B.n92 71.676
R980 B.n299 B.n91 71.676
R981 B.n295 B.n90 71.676
R982 B.n291 B.n89 71.676
R983 B.n287 B.n88 71.676
R984 B.n283 B.n87 71.676
R985 B.n279 B.n86 71.676
R986 B.n275 B.n85 71.676
R987 B.n271 B.n84 71.676
R988 B.n267 B.n83 71.676
R989 B.n263 B.n82 71.676
R990 B.n259 B.n81 71.676
R991 B.n254 B.n80 71.676
R992 B.n250 B.n79 71.676
R993 B.n246 B.n78 71.676
R994 B.n242 B.n77 71.676
R995 B.n238 B.n76 71.676
R996 B.n234 B.n75 71.676
R997 B.n230 B.n74 71.676
R998 B.n226 B.n73 71.676
R999 B.n222 B.n72 71.676
R1000 B.n218 B.n71 71.676
R1001 B.n214 B.n70 71.676
R1002 B.n210 B.n69 71.676
R1003 B.n206 B.n68 71.676
R1004 B.n202 B.n67 71.676
R1005 B.n198 B.n66 71.676
R1006 B.n194 B.n65 71.676
R1007 B.n190 B.n64 71.676
R1008 B.n186 B.n63 71.676
R1009 B.n182 B.n62 71.676
R1010 B.n178 B.n61 71.676
R1011 B.n174 B.n60 71.676
R1012 B.n170 B.n59 71.676
R1013 B.n166 B.n58 71.676
R1014 B.n162 B.n57 71.676
R1015 B.n158 B.n56 71.676
R1016 B.n154 B.n55 71.676
R1017 B.n150 B.n54 71.676
R1018 B.n146 B.n53 71.676
R1019 B.n142 B.n52 71.676
R1020 B.n138 B.n51 71.676
R1021 B.n134 B.n50 71.676
R1022 B.n130 B.n49 71.676
R1023 B.n126 B.n48 71.676
R1024 B.n122 B.n47 71.676
R1025 B.n862 B.n46 71.676
R1026 B.n756 B.n421 71.676
R1027 B.n750 B.n422 71.676
R1028 B.n746 B.n423 71.676
R1029 B.n742 B.n424 71.676
R1030 B.n738 B.n425 71.676
R1031 B.n734 B.n426 71.676
R1032 B.n730 B.n427 71.676
R1033 B.n726 B.n428 71.676
R1034 B.n722 B.n429 71.676
R1035 B.n718 B.n430 71.676
R1036 B.n714 B.n431 71.676
R1037 B.n710 B.n432 71.676
R1038 B.n706 B.n433 71.676
R1039 B.n702 B.n434 71.676
R1040 B.n698 B.n435 71.676
R1041 B.n694 B.n436 71.676
R1042 B.n690 B.n437 71.676
R1043 B.n686 B.n438 71.676
R1044 B.n682 B.n439 71.676
R1045 B.n678 B.n440 71.676
R1046 B.n674 B.n441 71.676
R1047 B.n670 B.n442 71.676
R1048 B.n666 B.n443 71.676
R1049 B.n662 B.n444 71.676
R1050 B.n658 B.n445 71.676
R1051 B.n654 B.n446 71.676
R1052 B.n650 B.n447 71.676
R1053 B.n646 B.n448 71.676
R1054 B.n642 B.n449 71.676
R1055 B.n638 B.n450 71.676
R1056 B.n633 B.n451 71.676
R1057 B.n629 B.n452 71.676
R1058 B.n625 B.n453 71.676
R1059 B.n621 B.n454 71.676
R1060 B.n617 B.n455 71.676
R1061 B.n613 B.n456 71.676
R1062 B.n609 B.n457 71.676
R1063 B.n605 B.n458 71.676
R1064 B.n601 B.n459 71.676
R1065 B.n597 B.n460 71.676
R1066 B.n593 B.n461 71.676
R1067 B.n589 B.n462 71.676
R1068 B.n585 B.n463 71.676
R1069 B.n581 B.n464 71.676
R1070 B.n577 B.n465 71.676
R1071 B.n573 B.n466 71.676
R1072 B.n569 B.n467 71.676
R1073 B.n565 B.n468 71.676
R1074 B.n561 B.n469 71.676
R1075 B.n557 B.n470 71.676
R1076 B.n553 B.n471 71.676
R1077 B.n549 B.n472 71.676
R1078 B.n545 B.n473 71.676
R1079 B.n541 B.n474 71.676
R1080 B.n537 B.n475 71.676
R1081 B.n533 B.n476 71.676
R1082 B.n529 B.n477 71.676
R1083 B.n525 B.n478 71.676
R1084 B.n521 B.n479 71.676
R1085 B.n517 B.n480 71.676
R1086 B.n513 B.n481 71.676
R1087 B.n509 B.n482 71.676
R1088 B.n505 B.n483 71.676
R1089 B.n501 B.n484 71.676
R1090 B.n497 B.n485 71.676
R1091 B.n493 B.n486 71.676
R1092 B.n492 B.n491 59.5399
R1093 B.n635 B.n489 59.5399
R1094 B.n118 B.n117 59.5399
R1095 B.n257 B.n115 59.5399
R1096 B.n755 B.n418 54.4627
R1097 B.n861 B.n43 54.4627
R1098 B.n762 B.n418 31.1218
R1099 B.n762 B.n414 31.1218
R1100 B.n769 B.n414 31.1218
R1101 B.n769 B.n768 31.1218
R1102 B.n775 B.n407 31.1218
R1103 B.n781 B.n407 31.1218
R1104 B.n781 B.n402 31.1218
R1105 B.n787 B.n402 31.1218
R1106 B.n787 B.n403 31.1218
R1107 B.n794 B.n793 31.1218
R1108 B.n800 B.n392 31.1218
R1109 B.n806 B.n392 31.1218
R1110 B.n812 B.n388 31.1218
R1111 B.n820 B.n384 31.1218
R1112 B.n820 B.n819 31.1218
R1113 B.n826 B.n4 31.1218
R1114 B.n910 B.n4 31.1218
R1115 B.n910 B.n909 31.1218
R1116 B.n909 B.n908 31.1218
R1117 B.n902 B.n11 31.1218
R1118 B.n902 B.n901 31.1218
R1119 B.n900 B.n15 31.1218
R1120 B.n894 B.n893 31.1218
R1121 B.n893 B.n892 31.1218
R1122 B.n886 B.n25 31.1218
R1123 B.n885 B.n884 31.1218
R1124 B.n884 B.n29 31.1218
R1125 B.n878 B.n29 31.1218
R1126 B.n878 B.n877 31.1218
R1127 B.n877 B.n876 31.1218
R1128 B.n870 B.n39 31.1218
R1129 B.n870 B.n869 31.1218
R1130 B.n869 B.n868 31.1218
R1131 B.n868 B.n43 31.1218
R1132 B.n859 B.n858 29.5029
R1133 B.n865 B.n864 29.5029
R1134 B.n494 B.n416 29.5029
R1135 B.n759 B.n758 29.5029
R1136 B.n826 B.t3 26.0875
R1137 B.n908 B.t7 26.0875
R1138 B.t0 B.n388 24.2568
R1139 B.t8 B.n15 24.2568
R1140 B.n793 B.t1 23.3415
R1141 B.n25 B.t9 23.3415
R1142 B.n794 B.t5 22.4261
R1143 B.n886 B.t2 22.4261
R1144 B.n812 B.t4 21.5108
R1145 B.t6 B.n900 21.5108
R1146 B.n768 B.t15 18.7648
R1147 B.n39 B.t11 18.7648
R1148 B B.n912 18.0485
R1149 B.n491 B.n490 16.2914
R1150 B.n489 B.n488 16.2914
R1151 B.n117 B.n116 16.2914
R1152 B.n115 B.n114 16.2914
R1153 B.n775 B.t15 12.3575
R1154 B.n876 B.t11 12.3575
R1155 B.n864 B.n45 10.6151
R1156 B.n120 B.n45 10.6151
R1157 B.n121 B.n120 10.6151
R1158 B.n124 B.n121 10.6151
R1159 B.n125 B.n124 10.6151
R1160 B.n128 B.n125 10.6151
R1161 B.n129 B.n128 10.6151
R1162 B.n132 B.n129 10.6151
R1163 B.n133 B.n132 10.6151
R1164 B.n136 B.n133 10.6151
R1165 B.n137 B.n136 10.6151
R1166 B.n140 B.n137 10.6151
R1167 B.n141 B.n140 10.6151
R1168 B.n144 B.n141 10.6151
R1169 B.n145 B.n144 10.6151
R1170 B.n148 B.n145 10.6151
R1171 B.n149 B.n148 10.6151
R1172 B.n152 B.n149 10.6151
R1173 B.n153 B.n152 10.6151
R1174 B.n156 B.n153 10.6151
R1175 B.n157 B.n156 10.6151
R1176 B.n160 B.n157 10.6151
R1177 B.n161 B.n160 10.6151
R1178 B.n164 B.n161 10.6151
R1179 B.n165 B.n164 10.6151
R1180 B.n168 B.n165 10.6151
R1181 B.n169 B.n168 10.6151
R1182 B.n172 B.n169 10.6151
R1183 B.n173 B.n172 10.6151
R1184 B.n176 B.n173 10.6151
R1185 B.n177 B.n176 10.6151
R1186 B.n180 B.n177 10.6151
R1187 B.n181 B.n180 10.6151
R1188 B.n184 B.n181 10.6151
R1189 B.n185 B.n184 10.6151
R1190 B.n188 B.n185 10.6151
R1191 B.n189 B.n188 10.6151
R1192 B.n192 B.n189 10.6151
R1193 B.n193 B.n192 10.6151
R1194 B.n196 B.n193 10.6151
R1195 B.n197 B.n196 10.6151
R1196 B.n200 B.n197 10.6151
R1197 B.n201 B.n200 10.6151
R1198 B.n204 B.n201 10.6151
R1199 B.n205 B.n204 10.6151
R1200 B.n208 B.n205 10.6151
R1201 B.n209 B.n208 10.6151
R1202 B.n212 B.n209 10.6151
R1203 B.n213 B.n212 10.6151
R1204 B.n216 B.n213 10.6151
R1205 B.n217 B.n216 10.6151
R1206 B.n220 B.n217 10.6151
R1207 B.n221 B.n220 10.6151
R1208 B.n224 B.n221 10.6151
R1209 B.n225 B.n224 10.6151
R1210 B.n228 B.n225 10.6151
R1211 B.n229 B.n228 10.6151
R1212 B.n232 B.n229 10.6151
R1213 B.n233 B.n232 10.6151
R1214 B.n236 B.n233 10.6151
R1215 B.n237 B.n236 10.6151
R1216 B.n241 B.n240 10.6151
R1217 B.n244 B.n241 10.6151
R1218 B.n245 B.n244 10.6151
R1219 B.n248 B.n245 10.6151
R1220 B.n249 B.n248 10.6151
R1221 B.n252 B.n249 10.6151
R1222 B.n253 B.n252 10.6151
R1223 B.n256 B.n253 10.6151
R1224 B.n261 B.n258 10.6151
R1225 B.n262 B.n261 10.6151
R1226 B.n265 B.n262 10.6151
R1227 B.n266 B.n265 10.6151
R1228 B.n269 B.n266 10.6151
R1229 B.n270 B.n269 10.6151
R1230 B.n273 B.n270 10.6151
R1231 B.n274 B.n273 10.6151
R1232 B.n277 B.n274 10.6151
R1233 B.n278 B.n277 10.6151
R1234 B.n281 B.n278 10.6151
R1235 B.n282 B.n281 10.6151
R1236 B.n285 B.n282 10.6151
R1237 B.n286 B.n285 10.6151
R1238 B.n289 B.n286 10.6151
R1239 B.n290 B.n289 10.6151
R1240 B.n293 B.n290 10.6151
R1241 B.n294 B.n293 10.6151
R1242 B.n297 B.n294 10.6151
R1243 B.n298 B.n297 10.6151
R1244 B.n301 B.n298 10.6151
R1245 B.n302 B.n301 10.6151
R1246 B.n305 B.n302 10.6151
R1247 B.n306 B.n305 10.6151
R1248 B.n309 B.n306 10.6151
R1249 B.n310 B.n309 10.6151
R1250 B.n313 B.n310 10.6151
R1251 B.n314 B.n313 10.6151
R1252 B.n317 B.n314 10.6151
R1253 B.n318 B.n317 10.6151
R1254 B.n321 B.n318 10.6151
R1255 B.n322 B.n321 10.6151
R1256 B.n325 B.n322 10.6151
R1257 B.n326 B.n325 10.6151
R1258 B.n329 B.n326 10.6151
R1259 B.n330 B.n329 10.6151
R1260 B.n333 B.n330 10.6151
R1261 B.n334 B.n333 10.6151
R1262 B.n337 B.n334 10.6151
R1263 B.n338 B.n337 10.6151
R1264 B.n341 B.n338 10.6151
R1265 B.n342 B.n341 10.6151
R1266 B.n345 B.n342 10.6151
R1267 B.n346 B.n345 10.6151
R1268 B.n349 B.n346 10.6151
R1269 B.n350 B.n349 10.6151
R1270 B.n353 B.n350 10.6151
R1271 B.n354 B.n353 10.6151
R1272 B.n357 B.n354 10.6151
R1273 B.n358 B.n357 10.6151
R1274 B.n361 B.n358 10.6151
R1275 B.n362 B.n361 10.6151
R1276 B.n365 B.n362 10.6151
R1277 B.n366 B.n365 10.6151
R1278 B.n369 B.n366 10.6151
R1279 B.n370 B.n369 10.6151
R1280 B.n373 B.n370 10.6151
R1281 B.n374 B.n373 10.6151
R1282 B.n377 B.n374 10.6151
R1283 B.n378 B.n377 10.6151
R1284 B.n859 B.n378 10.6151
R1285 B.n764 B.n416 10.6151
R1286 B.n765 B.n764 10.6151
R1287 B.n766 B.n765 10.6151
R1288 B.n766 B.n409 10.6151
R1289 B.n777 B.n409 10.6151
R1290 B.n778 B.n777 10.6151
R1291 B.n779 B.n778 10.6151
R1292 B.n779 B.n400 10.6151
R1293 B.n789 B.n400 10.6151
R1294 B.n790 B.n789 10.6151
R1295 B.n791 B.n790 10.6151
R1296 B.n791 B.n394 10.6151
R1297 B.n802 B.n394 10.6151
R1298 B.n803 B.n802 10.6151
R1299 B.n804 B.n803 10.6151
R1300 B.n804 B.n386 10.6151
R1301 B.n814 B.n386 10.6151
R1302 B.n815 B.n814 10.6151
R1303 B.n817 B.n815 10.6151
R1304 B.n817 B.n816 10.6151
R1305 B.n816 B.n379 10.6151
R1306 B.n829 B.n379 10.6151
R1307 B.n830 B.n829 10.6151
R1308 B.n831 B.n830 10.6151
R1309 B.n832 B.n831 10.6151
R1310 B.n834 B.n832 10.6151
R1311 B.n835 B.n834 10.6151
R1312 B.n836 B.n835 10.6151
R1313 B.n837 B.n836 10.6151
R1314 B.n839 B.n837 10.6151
R1315 B.n840 B.n839 10.6151
R1316 B.n841 B.n840 10.6151
R1317 B.n842 B.n841 10.6151
R1318 B.n844 B.n842 10.6151
R1319 B.n845 B.n844 10.6151
R1320 B.n846 B.n845 10.6151
R1321 B.n847 B.n846 10.6151
R1322 B.n849 B.n847 10.6151
R1323 B.n850 B.n849 10.6151
R1324 B.n851 B.n850 10.6151
R1325 B.n852 B.n851 10.6151
R1326 B.n854 B.n852 10.6151
R1327 B.n855 B.n854 10.6151
R1328 B.n856 B.n855 10.6151
R1329 B.n857 B.n856 10.6151
R1330 B.n858 B.n857 10.6151
R1331 B.n758 B.n420 10.6151
R1332 B.n753 B.n420 10.6151
R1333 B.n753 B.n752 10.6151
R1334 B.n752 B.n751 10.6151
R1335 B.n751 B.n748 10.6151
R1336 B.n748 B.n747 10.6151
R1337 B.n747 B.n744 10.6151
R1338 B.n744 B.n743 10.6151
R1339 B.n743 B.n740 10.6151
R1340 B.n740 B.n739 10.6151
R1341 B.n739 B.n736 10.6151
R1342 B.n736 B.n735 10.6151
R1343 B.n735 B.n732 10.6151
R1344 B.n732 B.n731 10.6151
R1345 B.n731 B.n728 10.6151
R1346 B.n728 B.n727 10.6151
R1347 B.n727 B.n724 10.6151
R1348 B.n724 B.n723 10.6151
R1349 B.n723 B.n720 10.6151
R1350 B.n720 B.n719 10.6151
R1351 B.n719 B.n716 10.6151
R1352 B.n716 B.n715 10.6151
R1353 B.n715 B.n712 10.6151
R1354 B.n712 B.n711 10.6151
R1355 B.n711 B.n708 10.6151
R1356 B.n708 B.n707 10.6151
R1357 B.n707 B.n704 10.6151
R1358 B.n704 B.n703 10.6151
R1359 B.n703 B.n700 10.6151
R1360 B.n700 B.n699 10.6151
R1361 B.n699 B.n696 10.6151
R1362 B.n696 B.n695 10.6151
R1363 B.n695 B.n692 10.6151
R1364 B.n692 B.n691 10.6151
R1365 B.n691 B.n688 10.6151
R1366 B.n688 B.n687 10.6151
R1367 B.n687 B.n684 10.6151
R1368 B.n684 B.n683 10.6151
R1369 B.n683 B.n680 10.6151
R1370 B.n680 B.n679 10.6151
R1371 B.n679 B.n676 10.6151
R1372 B.n676 B.n675 10.6151
R1373 B.n675 B.n672 10.6151
R1374 B.n672 B.n671 10.6151
R1375 B.n671 B.n668 10.6151
R1376 B.n668 B.n667 10.6151
R1377 B.n667 B.n664 10.6151
R1378 B.n664 B.n663 10.6151
R1379 B.n663 B.n660 10.6151
R1380 B.n660 B.n659 10.6151
R1381 B.n659 B.n656 10.6151
R1382 B.n656 B.n655 10.6151
R1383 B.n655 B.n652 10.6151
R1384 B.n652 B.n651 10.6151
R1385 B.n651 B.n648 10.6151
R1386 B.n648 B.n647 10.6151
R1387 B.n647 B.n644 10.6151
R1388 B.n644 B.n643 10.6151
R1389 B.n643 B.n640 10.6151
R1390 B.n640 B.n639 10.6151
R1391 B.n639 B.n636 10.6151
R1392 B.n634 B.n631 10.6151
R1393 B.n631 B.n630 10.6151
R1394 B.n630 B.n627 10.6151
R1395 B.n627 B.n626 10.6151
R1396 B.n626 B.n623 10.6151
R1397 B.n623 B.n622 10.6151
R1398 B.n622 B.n619 10.6151
R1399 B.n619 B.n618 10.6151
R1400 B.n615 B.n614 10.6151
R1401 B.n614 B.n611 10.6151
R1402 B.n611 B.n610 10.6151
R1403 B.n610 B.n607 10.6151
R1404 B.n607 B.n606 10.6151
R1405 B.n606 B.n603 10.6151
R1406 B.n603 B.n602 10.6151
R1407 B.n602 B.n599 10.6151
R1408 B.n599 B.n598 10.6151
R1409 B.n598 B.n595 10.6151
R1410 B.n595 B.n594 10.6151
R1411 B.n594 B.n591 10.6151
R1412 B.n591 B.n590 10.6151
R1413 B.n590 B.n587 10.6151
R1414 B.n587 B.n586 10.6151
R1415 B.n586 B.n583 10.6151
R1416 B.n583 B.n582 10.6151
R1417 B.n582 B.n579 10.6151
R1418 B.n579 B.n578 10.6151
R1419 B.n578 B.n575 10.6151
R1420 B.n575 B.n574 10.6151
R1421 B.n574 B.n571 10.6151
R1422 B.n571 B.n570 10.6151
R1423 B.n570 B.n567 10.6151
R1424 B.n567 B.n566 10.6151
R1425 B.n566 B.n563 10.6151
R1426 B.n563 B.n562 10.6151
R1427 B.n562 B.n559 10.6151
R1428 B.n559 B.n558 10.6151
R1429 B.n558 B.n555 10.6151
R1430 B.n555 B.n554 10.6151
R1431 B.n554 B.n551 10.6151
R1432 B.n551 B.n550 10.6151
R1433 B.n550 B.n547 10.6151
R1434 B.n547 B.n546 10.6151
R1435 B.n546 B.n543 10.6151
R1436 B.n543 B.n542 10.6151
R1437 B.n542 B.n539 10.6151
R1438 B.n539 B.n538 10.6151
R1439 B.n538 B.n535 10.6151
R1440 B.n535 B.n534 10.6151
R1441 B.n534 B.n531 10.6151
R1442 B.n531 B.n530 10.6151
R1443 B.n530 B.n527 10.6151
R1444 B.n527 B.n526 10.6151
R1445 B.n526 B.n523 10.6151
R1446 B.n523 B.n522 10.6151
R1447 B.n522 B.n519 10.6151
R1448 B.n519 B.n518 10.6151
R1449 B.n518 B.n515 10.6151
R1450 B.n515 B.n514 10.6151
R1451 B.n514 B.n511 10.6151
R1452 B.n511 B.n510 10.6151
R1453 B.n510 B.n507 10.6151
R1454 B.n507 B.n506 10.6151
R1455 B.n506 B.n503 10.6151
R1456 B.n503 B.n502 10.6151
R1457 B.n502 B.n499 10.6151
R1458 B.n499 B.n498 10.6151
R1459 B.n498 B.n495 10.6151
R1460 B.n495 B.n494 10.6151
R1461 B.n760 B.n759 10.6151
R1462 B.n760 B.n412 10.6151
R1463 B.n771 B.n412 10.6151
R1464 B.n772 B.n771 10.6151
R1465 B.n773 B.n772 10.6151
R1466 B.n773 B.n405 10.6151
R1467 B.n783 B.n405 10.6151
R1468 B.n784 B.n783 10.6151
R1469 B.n785 B.n784 10.6151
R1470 B.n785 B.n397 10.6151
R1471 B.n796 B.n397 10.6151
R1472 B.n797 B.n796 10.6151
R1473 B.n798 B.n797 10.6151
R1474 B.n798 B.n390 10.6151
R1475 B.n808 B.n390 10.6151
R1476 B.n809 B.n808 10.6151
R1477 B.n810 B.n809 10.6151
R1478 B.n810 B.n382 10.6151
R1479 B.n822 B.n382 10.6151
R1480 B.n823 B.n822 10.6151
R1481 B.n824 B.n823 10.6151
R1482 B.n824 B.n0 10.6151
R1483 B.n906 B.n1 10.6151
R1484 B.n906 B.n905 10.6151
R1485 B.n905 B.n904 10.6151
R1486 B.n904 B.n9 10.6151
R1487 B.n898 B.n9 10.6151
R1488 B.n898 B.n897 10.6151
R1489 B.n897 B.n896 10.6151
R1490 B.n896 B.n17 10.6151
R1491 B.n890 B.n17 10.6151
R1492 B.n890 B.n889 10.6151
R1493 B.n889 B.n888 10.6151
R1494 B.n888 B.n23 10.6151
R1495 B.n882 B.n23 10.6151
R1496 B.n882 B.n881 10.6151
R1497 B.n881 B.n880 10.6151
R1498 B.n880 B.n31 10.6151
R1499 B.n874 B.n31 10.6151
R1500 B.n874 B.n873 10.6151
R1501 B.n873 B.n872 10.6151
R1502 B.n872 B.n37 10.6151
R1503 B.n866 B.n37 10.6151
R1504 B.n866 B.n865 10.6151
R1505 B.t4 B.n384 9.61148
R1506 B.n901 B.t6 9.61148
R1507 B.n403 B.t5 8.69615
R1508 B.t2 B.n885 8.69615
R1509 B.n800 B.t1 7.78082
R1510 B.n892 B.t9 7.78082
R1511 B.n806 B.t0 6.86549
R1512 B.n894 B.t8 6.86549
R1513 B.n240 B.n118 6.5566
R1514 B.n257 B.n256 6.5566
R1515 B.n635 B.n634 6.5566
R1516 B.n618 B.n492 6.5566
R1517 B.n819 B.t3 5.03482
R1518 B.n11 B.t7 5.03482
R1519 B.n237 B.n118 4.05904
R1520 B.n258 B.n257 4.05904
R1521 B.n636 B.n635 4.05904
R1522 B.n615 B.n492 4.05904
R1523 B.n912 B.n0 2.81026
R1524 B.n912 B.n1 2.81026
R1525 VP.n5 VP.t5 985.455
R1526 VP.n16 VP.t3 964.472
R1527 VP.n17 VP.t2 964.472
R1528 VP.n1 VP.t1 964.472
R1529 VP.n23 VP.t0 964.472
R1530 VP.n24 VP.t8 964.472
R1531 VP.n13 VP.t6 964.472
R1532 VP.n12 VP.t7 964.472
R1533 VP.n4 VP.t9 964.472
R1534 VP.n6 VP.t4 964.472
R1535 VP.n25 VP.n24 161.3
R1536 VP.n8 VP.n7 161.3
R1537 VP.n9 VP.n4 161.3
R1538 VP.n11 VP.n10 161.3
R1539 VP.n12 VP.n3 161.3
R1540 VP.n14 VP.n13 161.3
R1541 VP.n23 VP.n0 161.3
R1542 VP.n22 VP.n21 161.3
R1543 VP.n20 VP.n1 161.3
R1544 VP.n19 VP.n18 161.3
R1545 VP.n17 VP.n2 161.3
R1546 VP.n16 VP.n15 161.3
R1547 VP.n8 VP.n5 70.4033
R1548 VP.n17 VP.n16 48.2005
R1549 VP.n24 VP.n23 48.2005
R1550 VP.n13 VP.n12 48.2005
R1551 VP.n15 VP.n14 46.9172
R1552 VP.n18 VP.n1 35.7853
R1553 VP.n22 VP.n1 35.7853
R1554 VP.n11 VP.n4 35.7853
R1555 VP.n7 VP.n4 35.7853
R1556 VP.n6 VP.n5 20.9576
R1557 VP.n18 VP.n17 12.4157
R1558 VP.n23 VP.n22 12.4157
R1559 VP.n12 VP.n11 12.4157
R1560 VP.n7 VP.n6 12.4157
R1561 VP.n9 VP.n8 0.189894
R1562 VP.n10 VP.n9 0.189894
R1563 VP.n10 VP.n3 0.189894
R1564 VP.n14 VP.n3 0.189894
R1565 VP.n15 VP.n2 0.189894
R1566 VP.n19 VP.n2 0.189894
R1567 VP.n20 VP.n19 0.189894
R1568 VP.n21 VP.n20 0.189894
R1569 VP.n21 VP.n0 0.189894
R1570 VP.n25 VP.n0 0.189894
R1571 VP VP.n25 0.0516364
R1572 VDD1.n102 VDD1.n101 289.615
R1573 VDD1.n207 VDD1.n206 289.615
R1574 VDD1.n101 VDD1.n100 185
R1575 VDD1.n2 VDD1.n1 185
R1576 VDD1.n95 VDD1.n94 185
R1577 VDD1.n93 VDD1.n92 185
R1578 VDD1.n6 VDD1.n5 185
R1579 VDD1.n87 VDD1.n86 185
R1580 VDD1.n85 VDD1.n84 185
R1581 VDD1.n10 VDD1.n9 185
R1582 VDD1.n79 VDD1.n78 185
R1583 VDD1.n77 VDD1.n76 185
R1584 VDD1.n14 VDD1.n13 185
R1585 VDD1.n71 VDD1.n70 185
R1586 VDD1.n69 VDD1.n68 185
R1587 VDD1.n18 VDD1.n17 185
R1588 VDD1.n63 VDD1.n62 185
R1589 VDD1.n61 VDD1.n60 185
R1590 VDD1.n22 VDD1.n21 185
R1591 VDD1.n26 VDD1.n24 185
R1592 VDD1.n55 VDD1.n54 185
R1593 VDD1.n53 VDD1.n52 185
R1594 VDD1.n28 VDD1.n27 185
R1595 VDD1.n47 VDD1.n46 185
R1596 VDD1.n45 VDD1.n44 185
R1597 VDD1.n32 VDD1.n31 185
R1598 VDD1.n39 VDD1.n38 185
R1599 VDD1.n37 VDD1.n36 185
R1600 VDD1.n140 VDD1.n139 185
R1601 VDD1.n142 VDD1.n141 185
R1602 VDD1.n135 VDD1.n134 185
R1603 VDD1.n148 VDD1.n147 185
R1604 VDD1.n150 VDD1.n149 185
R1605 VDD1.n131 VDD1.n130 185
R1606 VDD1.n157 VDD1.n156 185
R1607 VDD1.n158 VDD1.n129 185
R1608 VDD1.n160 VDD1.n159 185
R1609 VDD1.n127 VDD1.n126 185
R1610 VDD1.n166 VDD1.n165 185
R1611 VDD1.n168 VDD1.n167 185
R1612 VDD1.n123 VDD1.n122 185
R1613 VDD1.n174 VDD1.n173 185
R1614 VDD1.n176 VDD1.n175 185
R1615 VDD1.n119 VDD1.n118 185
R1616 VDD1.n182 VDD1.n181 185
R1617 VDD1.n184 VDD1.n183 185
R1618 VDD1.n115 VDD1.n114 185
R1619 VDD1.n190 VDD1.n189 185
R1620 VDD1.n192 VDD1.n191 185
R1621 VDD1.n111 VDD1.n110 185
R1622 VDD1.n198 VDD1.n197 185
R1623 VDD1.n200 VDD1.n199 185
R1624 VDD1.n107 VDD1.n106 185
R1625 VDD1.n206 VDD1.n205 185
R1626 VDD1.n35 VDD1.t0 149.524
R1627 VDD1.n138 VDD1.t1 149.524
R1628 VDD1.n101 VDD1.n1 104.615
R1629 VDD1.n94 VDD1.n1 104.615
R1630 VDD1.n94 VDD1.n93 104.615
R1631 VDD1.n93 VDD1.n5 104.615
R1632 VDD1.n86 VDD1.n5 104.615
R1633 VDD1.n86 VDD1.n85 104.615
R1634 VDD1.n85 VDD1.n9 104.615
R1635 VDD1.n78 VDD1.n9 104.615
R1636 VDD1.n78 VDD1.n77 104.615
R1637 VDD1.n77 VDD1.n13 104.615
R1638 VDD1.n70 VDD1.n13 104.615
R1639 VDD1.n70 VDD1.n69 104.615
R1640 VDD1.n69 VDD1.n17 104.615
R1641 VDD1.n62 VDD1.n17 104.615
R1642 VDD1.n62 VDD1.n61 104.615
R1643 VDD1.n61 VDD1.n21 104.615
R1644 VDD1.n26 VDD1.n21 104.615
R1645 VDD1.n54 VDD1.n26 104.615
R1646 VDD1.n54 VDD1.n53 104.615
R1647 VDD1.n53 VDD1.n27 104.615
R1648 VDD1.n46 VDD1.n27 104.615
R1649 VDD1.n46 VDD1.n45 104.615
R1650 VDD1.n45 VDD1.n31 104.615
R1651 VDD1.n38 VDD1.n31 104.615
R1652 VDD1.n38 VDD1.n37 104.615
R1653 VDD1.n141 VDD1.n140 104.615
R1654 VDD1.n141 VDD1.n134 104.615
R1655 VDD1.n148 VDD1.n134 104.615
R1656 VDD1.n149 VDD1.n148 104.615
R1657 VDD1.n149 VDD1.n130 104.615
R1658 VDD1.n157 VDD1.n130 104.615
R1659 VDD1.n158 VDD1.n157 104.615
R1660 VDD1.n159 VDD1.n158 104.615
R1661 VDD1.n159 VDD1.n126 104.615
R1662 VDD1.n166 VDD1.n126 104.615
R1663 VDD1.n167 VDD1.n166 104.615
R1664 VDD1.n167 VDD1.n122 104.615
R1665 VDD1.n174 VDD1.n122 104.615
R1666 VDD1.n175 VDD1.n174 104.615
R1667 VDD1.n175 VDD1.n118 104.615
R1668 VDD1.n182 VDD1.n118 104.615
R1669 VDD1.n183 VDD1.n182 104.615
R1670 VDD1.n183 VDD1.n114 104.615
R1671 VDD1.n190 VDD1.n114 104.615
R1672 VDD1.n191 VDD1.n190 104.615
R1673 VDD1.n191 VDD1.n110 104.615
R1674 VDD1.n198 VDD1.n110 104.615
R1675 VDD1.n199 VDD1.n198 104.615
R1676 VDD1.n199 VDD1.n106 104.615
R1677 VDD1.n206 VDD1.n106 104.615
R1678 VDD1.n211 VDD1.n210 63.7589
R1679 VDD1.n104 VDD1.n103 63.2721
R1680 VDD1.n209 VDD1.n208 63.2711
R1681 VDD1.n213 VDD1.n212 63.271
R1682 VDD1.n37 VDD1.t0 52.3082
R1683 VDD1.n140 VDD1.t1 52.3082
R1684 VDD1.n104 VDD1.n102 52.3034
R1685 VDD1.n209 VDD1.n207 52.3034
R1686 VDD1.n213 VDD1.n211 44.2724
R1687 VDD1.n24 VDD1.n22 13.1884
R1688 VDD1.n160 VDD1.n127 13.1884
R1689 VDD1.n100 VDD1.n0 12.8005
R1690 VDD1.n60 VDD1.n59 12.8005
R1691 VDD1.n56 VDD1.n55 12.8005
R1692 VDD1.n161 VDD1.n129 12.8005
R1693 VDD1.n165 VDD1.n164 12.8005
R1694 VDD1.n205 VDD1.n105 12.8005
R1695 VDD1.n99 VDD1.n2 12.0247
R1696 VDD1.n63 VDD1.n20 12.0247
R1697 VDD1.n52 VDD1.n25 12.0247
R1698 VDD1.n156 VDD1.n155 12.0247
R1699 VDD1.n168 VDD1.n125 12.0247
R1700 VDD1.n204 VDD1.n107 12.0247
R1701 VDD1.n96 VDD1.n95 11.249
R1702 VDD1.n64 VDD1.n18 11.249
R1703 VDD1.n51 VDD1.n28 11.249
R1704 VDD1.n154 VDD1.n131 11.249
R1705 VDD1.n169 VDD1.n123 11.249
R1706 VDD1.n201 VDD1.n200 11.249
R1707 VDD1.n92 VDD1.n4 10.4732
R1708 VDD1.n68 VDD1.n67 10.4732
R1709 VDD1.n48 VDD1.n47 10.4732
R1710 VDD1.n151 VDD1.n150 10.4732
R1711 VDD1.n173 VDD1.n172 10.4732
R1712 VDD1.n197 VDD1.n109 10.4732
R1713 VDD1.n36 VDD1.n35 10.2747
R1714 VDD1.n139 VDD1.n138 10.2747
R1715 VDD1.n91 VDD1.n6 9.69747
R1716 VDD1.n71 VDD1.n16 9.69747
R1717 VDD1.n44 VDD1.n30 9.69747
R1718 VDD1.n147 VDD1.n133 9.69747
R1719 VDD1.n176 VDD1.n121 9.69747
R1720 VDD1.n196 VDD1.n111 9.69747
R1721 VDD1.n98 VDD1.n0 9.45567
R1722 VDD1.n203 VDD1.n105 9.45567
R1723 VDD1.n34 VDD1.n33 9.3005
R1724 VDD1.n41 VDD1.n40 9.3005
R1725 VDD1.n43 VDD1.n42 9.3005
R1726 VDD1.n30 VDD1.n29 9.3005
R1727 VDD1.n49 VDD1.n48 9.3005
R1728 VDD1.n51 VDD1.n50 9.3005
R1729 VDD1.n25 VDD1.n23 9.3005
R1730 VDD1.n57 VDD1.n56 9.3005
R1731 VDD1.n83 VDD1.n82 9.3005
R1732 VDD1.n8 VDD1.n7 9.3005
R1733 VDD1.n89 VDD1.n88 9.3005
R1734 VDD1.n91 VDD1.n90 9.3005
R1735 VDD1.n4 VDD1.n3 9.3005
R1736 VDD1.n97 VDD1.n96 9.3005
R1737 VDD1.n99 VDD1.n98 9.3005
R1738 VDD1.n81 VDD1.n80 9.3005
R1739 VDD1.n12 VDD1.n11 9.3005
R1740 VDD1.n75 VDD1.n74 9.3005
R1741 VDD1.n73 VDD1.n72 9.3005
R1742 VDD1.n16 VDD1.n15 9.3005
R1743 VDD1.n67 VDD1.n66 9.3005
R1744 VDD1.n65 VDD1.n64 9.3005
R1745 VDD1.n20 VDD1.n19 9.3005
R1746 VDD1.n59 VDD1.n58 9.3005
R1747 VDD1.n186 VDD1.n185 9.3005
R1748 VDD1.n188 VDD1.n187 9.3005
R1749 VDD1.n113 VDD1.n112 9.3005
R1750 VDD1.n194 VDD1.n193 9.3005
R1751 VDD1.n196 VDD1.n195 9.3005
R1752 VDD1.n109 VDD1.n108 9.3005
R1753 VDD1.n202 VDD1.n201 9.3005
R1754 VDD1.n204 VDD1.n203 9.3005
R1755 VDD1.n180 VDD1.n179 9.3005
R1756 VDD1.n178 VDD1.n177 9.3005
R1757 VDD1.n121 VDD1.n120 9.3005
R1758 VDD1.n172 VDD1.n171 9.3005
R1759 VDD1.n170 VDD1.n169 9.3005
R1760 VDD1.n125 VDD1.n124 9.3005
R1761 VDD1.n164 VDD1.n163 9.3005
R1762 VDD1.n137 VDD1.n136 9.3005
R1763 VDD1.n144 VDD1.n143 9.3005
R1764 VDD1.n146 VDD1.n145 9.3005
R1765 VDD1.n133 VDD1.n132 9.3005
R1766 VDD1.n152 VDD1.n151 9.3005
R1767 VDD1.n154 VDD1.n153 9.3005
R1768 VDD1.n155 VDD1.n128 9.3005
R1769 VDD1.n162 VDD1.n161 9.3005
R1770 VDD1.n117 VDD1.n116 9.3005
R1771 VDD1.n88 VDD1.n87 8.92171
R1772 VDD1.n72 VDD1.n14 8.92171
R1773 VDD1.n43 VDD1.n32 8.92171
R1774 VDD1.n146 VDD1.n135 8.92171
R1775 VDD1.n177 VDD1.n119 8.92171
R1776 VDD1.n193 VDD1.n192 8.92171
R1777 VDD1.n84 VDD1.n8 8.14595
R1778 VDD1.n76 VDD1.n75 8.14595
R1779 VDD1.n40 VDD1.n39 8.14595
R1780 VDD1.n143 VDD1.n142 8.14595
R1781 VDD1.n181 VDD1.n180 8.14595
R1782 VDD1.n189 VDD1.n113 8.14595
R1783 VDD1.n83 VDD1.n10 7.3702
R1784 VDD1.n79 VDD1.n12 7.3702
R1785 VDD1.n36 VDD1.n34 7.3702
R1786 VDD1.n139 VDD1.n137 7.3702
R1787 VDD1.n184 VDD1.n117 7.3702
R1788 VDD1.n188 VDD1.n115 7.3702
R1789 VDD1.n80 VDD1.n10 6.59444
R1790 VDD1.n80 VDD1.n79 6.59444
R1791 VDD1.n185 VDD1.n184 6.59444
R1792 VDD1.n185 VDD1.n115 6.59444
R1793 VDD1.n84 VDD1.n83 5.81868
R1794 VDD1.n76 VDD1.n12 5.81868
R1795 VDD1.n39 VDD1.n34 5.81868
R1796 VDD1.n142 VDD1.n137 5.81868
R1797 VDD1.n181 VDD1.n117 5.81868
R1798 VDD1.n189 VDD1.n188 5.81868
R1799 VDD1.n87 VDD1.n8 5.04292
R1800 VDD1.n75 VDD1.n14 5.04292
R1801 VDD1.n40 VDD1.n32 5.04292
R1802 VDD1.n143 VDD1.n135 5.04292
R1803 VDD1.n180 VDD1.n119 5.04292
R1804 VDD1.n192 VDD1.n113 5.04292
R1805 VDD1.n88 VDD1.n6 4.26717
R1806 VDD1.n72 VDD1.n71 4.26717
R1807 VDD1.n44 VDD1.n43 4.26717
R1808 VDD1.n147 VDD1.n146 4.26717
R1809 VDD1.n177 VDD1.n176 4.26717
R1810 VDD1.n193 VDD1.n111 4.26717
R1811 VDD1.n92 VDD1.n91 3.49141
R1812 VDD1.n68 VDD1.n16 3.49141
R1813 VDD1.n47 VDD1.n30 3.49141
R1814 VDD1.n150 VDD1.n133 3.49141
R1815 VDD1.n173 VDD1.n121 3.49141
R1816 VDD1.n197 VDD1.n196 3.49141
R1817 VDD1.n138 VDD1.n136 2.84303
R1818 VDD1.n35 VDD1.n33 2.84303
R1819 VDD1.n95 VDD1.n4 2.71565
R1820 VDD1.n67 VDD1.n18 2.71565
R1821 VDD1.n48 VDD1.n28 2.71565
R1822 VDD1.n151 VDD1.n131 2.71565
R1823 VDD1.n172 VDD1.n123 2.71565
R1824 VDD1.n200 VDD1.n109 2.71565
R1825 VDD1.n96 VDD1.n2 1.93989
R1826 VDD1.n64 VDD1.n63 1.93989
R1827 VDD1.n52 VDD1.n51 1.93989
R1828 VDD1.n156 VDD1.n154 1.93989
R1829 VDD1.n169 VDD1.n168 1.93989
R1830 VDD1.n201 VDD1.n107 1.93989
R1831 VDD1.n100 VDD1.n99 1.16414
R1832 VDD1.n60 VDD1.n20 1.16414
R1833 VDD1.n55 VDD1.n25 1.16414
R1834 VDD1.n155 VDD1.n129 1.16414
R1835 VDD1.n165 VDD1.n125 1.16414
R1836 VDD1.n205 VDD1.n204 1.16414
R1837 VDD1.n212 VDD1.t6 1.05594
R1838 VDD1.n212 VDD1.t9 1.05594
R1839 VDD1.n103 VDD1.t2 1.05594
R1840 VDD1.n103 VDD1.t5 1.05594
R1841 VDD1.n210 VDD1.t7 1.05594
R1842 VDD1.n210 VDD1.t8 1.05594
R1843 VDD1.n208 VDD1.t3 1.05594
R1844 VDD1.n208 VDD1.t4 1.05594
R1845 VDD1 VDD1.n213 0.485414
R1846 VDD1.n102 VDD1.n0 0.388379
R1847 VDD1.n59 VDD1.n22 0.388379
R1848 VDD1.n56 VDD1.n24 0.388379
R1849 VDD1.n161 VDD1.n160 0.388379
R1850 VDD1.n164 VDD1.n127 0.388379
R1851 VDD1.n207 VDD1.n105 0.388379
R1852 VDD1 VDD1.n104 0.239724
R1853 VDD1.n98 VDD1.n97 0.155672
R1854 VDD1.n97 VDD1.n3 0.155672
R1855 VDD1.n90 VDD1.n3 0.155672
R1856 VDD1.n90 VDD1.n89 0.155672
R1857 VDD1.n89 VDD1.n7 0.155672
R1858 VDD1.n82 VDD1.n7 0.155672
R1859 VDD1.n82 VDD1.n81 0.155672
R1860 VDD1.n81 VDD1.n11 0.155672
R1861 VDD1.n74 VDD1.n11 0.155672
R1862 VDD1.n74 VDD1.n73 0.155672
R1863 VDD1.n73 VDD1.n15 0.155672
R1864 VDD1.n66 VDD1.n15 0.155672
R1865 VDD1.n66 VDD1.n65 0.155672
R1866 VDD1.n65 VDD1.n19 0.155672
R1867 VDD1.n58 VDD1.n19 0.155672
R1868 VDD1.n58 VDD1.n57 0.155672
R1869 VDD1.n57 VDD1.n23 0.155672
R1870 VDD1.n50 VDD1.n23 0.155672
R1871 VDD1.n50 VDD1.n49 0.155672
R1872 VDD1.n49 VDD1.n29 0.155672
R1873 VDD1.n42 VDD1.n29 0.155672
R1874 VDD1.n42 VDD1.n41 0.155672
R1875 VDD1.n41 VDD1.n33 0.155672
R1876 VDD1.n144 VDD1.n136 0.155672
R1877 VDD1.n145 VDD1.n144 0.155672
R1878 VDD1.n145 VDD1.n132 0.155672
R1879 VDD1.n152 VDD1.n132 0.155672
R1880 VDD1.n153 VDD1.n152 0.155672
R1881 VDD1.n153 VDD1.n128 0.155672
R1882 VDD1.n162 VDD1.n128 0.155672
R1883 VDD1.n163 VDD1.n162 0.155672
R1884 VDD1.n163 VDD1.n124 0.155672
R1885 VDD1.n170 VDD1.n124 0.155672
R1886 VDD1.n171 VDD1.n170 0.155672
R1887 VDD1.n171 VDD1.n120 0.155672
R1888 VDD1.n178 VDD1.n120 0.155672
R1889 VDD1.n179 VDD1.n178 0.155672
R1890 VDD1.n179 VDD1.n116 0.155672
R1891 VDD1.n186 VDD1.n116 0.155672
R1892 VDD1.n187 VDD1.n186 0.155672
R1893 VDD1.n187 VDD1.n112 0.155672
R1894 VDD1.n194 VDD1.n112 0.155672
R1895 VDD1.n195 VDD1.n194 0.155672
R1896 VDD1.n195 VDD1.n108 0.155672
R1897 VDD1.n202 VDD1.n108 0.155672
R1898 VDD1.n203 VDD1.n202 0.155672
R1899 VDD1.n211 VDD1.n209 0.126188
R1900 VTAIL.n428 VTAIL.n427 289.615
R1901 VTAIL.n104 VTAIL.n103 289.615
R1902 VTAIL.n324 VTAIL.n323 289.615
R1903 VTAIL.n216 VTAIL.n215 289.615
R1904 VTAIL.n361 VTAIL.n360 185
R1905 VTAIL.n363 VTAIL.n362 185
R1906 VTAIL.n356 VTAIL.n355 185
R1907 VTAIL.n369 VTAIL.n368 185
R1908 VTAIL.n371 VTAIL.n370 185
R1909 VTAIL.n352 VTAIL.n351 185
R1910 VTAIL.n378 VTAIL.n377 185
R1911 VTAIL.n379 VTAIL.n350 185
R1912 VTAIL.n381 VTAIL.n380 185
R1913 VTAIL.n348 VTAIL.n347 185
R1914 VTAIL.n387 VTAIL.n386 185
R1915 VTAIL.n389 VTAIL.n388 185
R1916 VTAIL.n344 VTAIL.n343 185
R1917 VTAIL.n395 VTAIL.n394 185
R1918 VTAIL.n397 VTAIL.n396 185
R1919 VTAIL.n340 VTAIL.n339 185
R1920 VTAIL.n403 VTAIL.n402 185
R1921 VTAIL.n405 VTAIL.n404 185
R1922 VTAIL.n336 VTAIL.n335 185
R1923 VTAIL.n411 VTAIL.n410 185
R1924 VTAIL.n413 VTAIL.n412 185
R1925 VTAIL.n332 VTAIL.n331 185
R1926 VTAIL.n419 VTAIL.n418 185
R1927 VTAIL.n421 VTAIL.n420 185
R1928 VTAIL.n328 VTAIL.n327 185
R1929 VTAIL.n427 VTAIL.n426 185
R1930 VTAIL.n37 VTAIL.n36 185
R1931 VTAIL.n39 VTAIL.n38 185
R1932 VTAIL.n32 VTAIL.n31 185
R1933 VTAIL.n45 VTAIL.n44 185
R1934 VTAIL.n47 VTAIL.n46 185
R1935 VTAIL.n28 VTAIL.n27 185
R1936 VTAIL.n54 VTAIL.n53 185
R1937 VTAIL.n55 VTAIL.n26 185
R1938 VTAIL.n57 VTAIL.n56 185
R1939 VTAIL.n24 VTAIL.n23 185
R1940 VTAIL.n63 VTAIL.n62 185
R1941 VTAIL.n65 VTAIL.n64 185
R1942 VTAIL.n20 VTAIL.n19 185
R1943 VTAIL.n71 VTAIL.n70 185
R1944 VTAIL.n73 VTAIL.n72 185
R1945 VTAIL.n16 VTAIL.n15 185
R1946 VTAIL.n79 VTAIL.n78 185
R1947 VTAIL.n81 VTAIL.n80 185
R1948 VTAIL.n12 VTAIL.n11 185
R1949 VTAIL.n87 VTAIL.n86 185
R1950 VTAIL.n89 VTAIL.n88 185
R1951 VTAIL.n8 VTAIL.n7 185
R1952 VTAIL.n95 VTAIL.n94 185
R1953 VTAIL.n97 VTAIL.n96 185
R1954 VTAIL.n4 VTAIL.n3 185
R1955 VTAIL.n103 VTAIL.n102 185
R1956 VTAIL.n323 VTAIL.n322 185
R1957 VTAIL.n224 VTAIL.n223 185
R1958 VTAIL.n317 VTAIL.n316 185
R1959 VTAIL.n315 VTAIL.n314 185
R1960 VTAIL.n228 VTAIL.n227 185
R1961 VTAIL.n309 VTAIL.n308 185
R1962 VTAIL.n307 VTAIL.n306 185
R1963 VTAIL.n232 VTAIL.n231 185
R1964 VTAIL.n301 VTAIL.n300 185
R1965 VTAIL.n299 VTAIL.n298 185
R1966 VTAIL.n236 VTAIL.n235 185
R1967 VTAIL.n293 VTAIL.n292 185
R1968 VTAIL.n291 VTAIL.n290 185
R1969 VTAIL.n240 VTAIL.n239 185
R1970 VTAIL.n285 VTAIL.n284 185
R1971 VTAIL.n283 VTAIL.n282 185
R1972 VTAIL.n244 VTAIL.n243 185
R1973 VTAIL.n248 VTAIL.n246 185
R1974 VTAIL.n277 VTAIL.n276 185
R1975 VTAIL.n275 VTAIL.n274 185
R1976 VTAIL.n250 VTAIL.n249 185
R1977 VTAIL.n269 VTAIL.n268 185
R1978 VTAIL.n267 VTAIL.n266 185
R1979 VTAIL.n254 VTAIL.n253 185
R1980 VTAIL.n261 VTAIL.n260 185
R1981 VTAIL.n259 VTAIL.n258 185
R1982 VTAIL.n215 VTAIL.n214 185
R1983 VTAIL.n116 VTAIL.n115 185
R1984 VTAIL.n209 VTAIL.n208 185
R1985 VTAIL.n207 VTAIL.n206 185
R1986 VTAIL.n120 VTAIL.n119 185
R1987 VTAIL.n201 VTAIL.n200 185
R1988 VTAIL.n199 VTAIL.n198 185
R1989 VTAIL.n124 VTAIL.n123 185
R1990 VTAIL.n193 VTAIL.n192 185
R1991 VTAIL.n191 VTAIL.n190 185
R1992 VTAIL.n128 VTAIL.n127 185
R1993 VTAIL.n185 VTAIL.n184 185
R1994 VTAIL.n183 VTAIL.n182 185
R1995 VTAIL.n132 VTAIL.n131 185
R1996 VTAIL.n177 VTAIL.n176 185
R1997 VTAIL.n175 VTAIL.n174 185
R1998 VTAIL.n136 VTAIL.n135 185
R1999 VTAIL.n140 VTAIL.n138 185
R2000 VTAIL.n169 VTAIL.n168 185
R2001 VTAIL.n167 VTAIL.n166 185
R2002 VTAIL.n142 VTAIL.n141 185
R2003 VTAIL.n161 VTAIL.n160 185
R2004 VTAIL.n159 VTAIL.n158 185
R2005 VTAIL.n146 VTAIL.n145 185
R2006 VTAIL.n153 VTAIL.n152 185
R2007 VTAIL.n151 VTAIL.n150 185
R2008 VTAIL.n359 VTAIL.t0 149.524
R2009 VTAIL.n35 VTAIL.t8 149.524
R2010 VTAIL.n257 VTAIL.t10 149.524
R2011 VTAIL.n149 VTAIL.t1 149.524
R2012 VTAIL.n362 VTAIL.n361 104.615
R2013 VTAIL.n362 VTAIL.n355 104.615
R2014 VTAIL.n369 VTAIL.n355 104.615
R2015 VTAIL.n370 VTAIL.n369 104.615
R2016 VTAIL.n370 VTAIL.n351 104.615
R2017 VTAIL.n378 VTAIL.n351 104.615
R2018 VTAIL.n379 VTAIL.n378 104.615
R2019 VTAIL.n380 VTAIL.n379 104.615
R2020 VTAIL.n380 VTAIL.n347 104.615
R2021 VTAIL.n387 VTAIL.n347 104.615
R2022 VTAIL.n388 VTAIL.n387 104.615
R2023 VTAIL.n388 VTAIL.n343 104.615
R2024 VTAIL.n395 VTAIL.n343 104.615
R2025 VTAIL.n396 VTAIL.n395 104.615
R2026 VTAIL.n396 VTAIL.n339 104.615
R2027 VTAIL.n403 VTAIL.n339 104.615
R2028 VTAIL.n404 VTAIL.n403 104.615
R2029 VTAIL.n404 VTAIL.n335 104.615
R2030 VTAIL.n411 VTAIL.n335 104.615
R2031 VTAIL.n412 VTAIL.n411 104.615
R2032 VTAIL.n412 VTAIL.n331 104.615
R2033 VTAIL.n419 VTAIL.n331 104.615
R2034 VTAIL.n420 VTAIL.n419 104.615
R2035 VTAIL.n420 VTAIL.n327 104.615
R2036 VTAIL.n427 VTAIL.n327 104.615
R2037 VTAIL.n38 VTAIL.n37 104.615
R2038 VTAIL.n38 VTAIL.n31 104.615
R2039 VTAIL.n45 VTAIL.n31 104.615
R2040 VTAIL.n46 VTAIL.n45 104.615
R2041 VTAIL.n46 VTAIL.n27 104.615
R2042 VTAIL.n54 VTAIL.n27 104.615
R2043 VTAIL.n55 VTAIL.n54 104.615
R2044 VTAIL.n56 VTAIL.n55 104.615
R2045 VTAIL.n56 VTAIL.n23 104.615
R2046 VTAIL.n63 VTAIL.n23 104.615
R2047 VTAIL.n64 VTAIL.n63 104.615
R2048 VTAIL.n64 VTAIL.n19 104.615
R2049 VTAIL.n71 VTAIL.n19 104.615
R2050 VTAIL.n72 VTAIL.n71 104.615
R2051 VTAIL.n72 VTAIL.n15 104.615
R2052 VTAIL.n79 VTAIL.n15 104.615
R2053 VTAIL.n80 VTAIL.n79 104.615
R2054 VTAIL.n80 VTAIL.n11 104.615
R2055 VTAIL.n87 VTAIL.n11 104.615
R2056 VTAIL.n88 VTAIL.n87 104.615
R2057 VTAIL.n88 VTAIL.n7 104.615
R2058 VTAIL.n95 VTAIL.n7 104.615
R2059 VTAIL.n96 VTAIL.n95 104.615
R2060 VTAIL.n96 VTAIL.n3 104.615
R2061 VTAIL.n103 VTAIL.n3 104.615
R2062 VTAIL.n323 VTAIL.n223 104.615
R2063 VTAIL.n316 VTAIL.n223 104.615
R2064 VTAIL.n316 VTAIL.n315 104.615
R2065 VTAIL.n315 VTAIL.n227 104.615
R2066 VTAIL.n308 VTAIL.n227 104.615
R2067 VTAIL.n308 VTAIL.n307 104.615
R2068 VTAIL.n307 VTAIL.n231 104.615
R2069 VTAIL.n300 VTAIL.n231 104.615
R2070 VTAIL.n300 VTAIL.n299 104.615
R2071 VTAIL.n299 VTAIL.n235 104.615
R2072 VTAIL.n292 VTAIL.n235 104.615
R2073 VTAIL.n292 VTAIL.n291 104.615
R2074 VTAIL.n291 VTAIL.n239 104.615
R2075 VTAIL.n284 VTAIL.n239 104.615
R2076 VTAIL.n284 VTAIL.n283 104.615
R2077 VTAIL.n283 VTAIL.n243 104.615
R2078 VTAIL.n248 VTAIL.n243 104.615
R2079 VTAIL.n276 VTAIL.n248 104.615
R2080 VTAIL.n276 VTAIL.n275 104.615
R2081 VTAIL.n275 VTAIL.n249 104.615
R2082 VTAIL.n268 VTAIL.n249 104.615
R2083 VTAIL.n268 VTAIL.n267 104.615
R2084 VTAIL.n267 VTAIL.n253 104.615
R2085 VTAIL.n260 VTAIL.n253 104.615
R2086 VTAIL.n260 VTAIL.n259 104.615
R2087 VTAIL.n215 VTAIL.n115 104.615
R2088 VTAIL.n208 VTAIL.n115 104.615
R2089 VTAIL.n208 VTAIL.n207 104.615
R2090 VTAIL.n207 VTAIL.n119 104.615
R2091 VTAIL.n200 VTAIL.n119 104.615
R2092 VTAIL.n200 VTAIL.n199 104.615
R2093 VTAIL.n199 VTAIL.n123 104.615
R2094 VTAIL.n192 VTAIL.n123 104.615
R2095 VTAIL.n192 VTAIL.n191 104.615
R2096 VTAIL.n191 VTAIL.n127 104.615
R2097 VTAIL.n184 VTAIL.n127 104.615
R2098 VTAIL.n184 VTAIL.n183 104.615
R2099 VTAIL.n183 VTAIL.n131 104.615
R2100 VTAIL.n176 VTAIL.n131 104.615
R2101 VTAIL.n176 VTAIL.n175 104.615
R2102 VTAIL.n175 VTAIL.n135 104.615
R2103 VTAIL.n140 VTAIL.n135 104.615
R2104 VTAIL.n168 VTAIL.n140 104.615
R2105 VTAIL.n168 VTAIL.n167 104.615
R2106 VTAIL.n167 VTAIL.n141 104.615
R2107 VTAIL.n160 VTAIL.n141 104.615
R2108 VTAIL.n160 VTAIL.n159 104.615
R2109 VTAIL.n159 VTAIL.n145 104.615
R2110 VTAIL.n152 VTAIL.n145 104.615
R2111 VTAIL.n152 VTAIL.n151 104.615
R2112 VTAIL.n361 VTAIL.t0 52.3082
R2113 VTAIL.n37 VTAIL.t8 52.3082
R2114 VTAIL.n259 VTAIL.t10 52.3082
R2115 VTAIL.n151 VTAIL.t1 52.3082
R2116 VTAIL.n221 VTAIL.n220 46.5933
R2117 VTAIL.n219 VTAIL.n218 46.5933
R2118 VTAIL.n113 VTAIL.n112 46.5933
R2119 VTAIL.n111 VTAIL.n110 46.5933
R2120 VTAIL.n431 VTAIL.n430 46.5923
R2121 VTAIL.n1 VTAIL.n0 46.5923
R2122 VTAIL.n107 VTAIL.n106 46.5923
R2123 VTAIL.n109 VTAIL.n108 46.5923
R2124 VTAIL.n429 VTAIL.n428 34.9005
R2125 VTAIL.n105 VTAIL.n104 34.9005
R2126 VTAIL.n325 VTAIL.n324 34.9005
R2127 VTAIL.n217 VTAIL.n216 34.9005
R2128 VTAIL.n111 VTAIL.n109 29.9876
R2129 VTAIL.n429 VTAIL.n325 29.2634
R2130 VTAIL.n381 VTAIL.n348 13.1884
R2131 VTAIL.n57 VTAIL.n24 13.1884
R2132 VTAIL.n246 VTAIL.n244 13.1884
R2133 VTAIL.n138 VTAIL.n136 13.1884
R2134 VTAIL.n382 VTAIL.n350 12.8005
R2135 VTAIL.n386 VTAIL.n385 12.8005
R2136 VTAIL.n426 VTAIL.n326 12.8005
R2137 VTAIL.n58 VTAIL.n26 12.8005
R2138 VTAIL.n62 VTAIL.n61 12.8005
R2139 VTAIL.n102 VTAIL.n2 12.8005
R2140 VTAIL.n322 VTAIL.n222 12.8005
R2141 VTAIL.n282 VTAIL.n281 12.8005
R2142 VTAIL.n278 VTAIL.n277 12.8005
R2143 VTAIL.n214 VTAIL.n114 12.8005
R2144 VTAIL.n174 VTAIL.n173 12.8005
R2145 VTAIL.n170 VTAIL.n169 12.8005
R2146 VTAIL.n377 VTAIL.n376 12.0247
R2147 VTAIL.n389 VTAIL.n346 12.0247
R2148 VTAIL.n425 VTAIL.n328 12.0247
R2149 VTAIL.n53 VTAIL.n52 12.0247
R2150 VTAIL.n65 VTAIL.n22 12.0247
R2151 VTAIL.n101 VTAIL.n4 12.0247
R2152 VTAIL.n321 VTAIL.n224 12.0247
R2153 VTAIL.n285 VTAIL.n242 12.0247
R2154 VTAIL.n274 VTAIL.n247 12.0247
R2155 VTAIL.n213 VTAIL.n116 12.0247
R2156 VTAIL.n177 VTAIL.n134 12.0247
R2157 VTAIL.n166 VTAIL.n139 12.0247
R2158 VTAIL.n375 VTAIL.n352 11.249
R2159 VTAIL.n390 VTAIL.n344 11.249
R2160 VTAIL.n422 VTAIL.n421 11.249
R2161 VTAIL.n51 VTAIL.n28 11.249
R2162 VTAIL.n66 VTAIL.n20 11.249
R2163 VTAIL.n98 VTAIL.n97 11.249
R2164 VTAIL.n318 VTAIL.n317 11.249
R2165 VTAIL.n286 VTAIL.n240 11.249
R2166 VTAIL.n273 VTAIL.n250 11.249
R2167 VTAIL.n210 VTAIL.n209 11.249
R2168 VTAIL.n178 VTAIL.n132 11.249
R2169 VTAIL.n165 VTAIL.n142 11.249
R2170 VTAIL.n372 VTAIL.n371 10.4732
R2171 VTAIL.n394 VTAIL.n393 10.4732
R2172 VTAIL.n418 VTAIL.n330 10.4732
R2173 VTAIL.n48 VTAIL.n47 10.4732
R2174 VTAIL.n70 VTAIL.n69 10.4732
R2175 VTAIL.n94 VTAIL.n6 10.4732
R2176 VTAIL.n314 VTAIL.n226 10.4732
R2177 VTAIL.n290 VTAIL.n289 10.4732
R2178 VTAIL.n270 VTAIL.n269 10.4732
R2179 VTAIL.n206 VTAIL.n118 10.4732
R2180 VTAIL.n182 VTAIL.n181 10.4732
R2181 VTAIL.n162 VTAIL.n161 10.4732
R2182 VTAIL.n360 VTAIL.n359 10.2747
R2183 VTAIL.n36 VTAIL.n35 10.2747
R2184 VTAIL.n258 VTAIL.n257 10.2747
R2185 VTAIL.n150 VTAIL.n149 10.2747
R2186 VTAIL.n368 VTAIL.n354 9.69747
R2187 VTAIL.n397 VTAIL.n342 9.69747
R2188 VTAIL.n417 VTAIL.n332 9.69747
R2189 VTAIL.n44 VTAIL.n30 9.69747
R2190 VTAIL.n73 VTAIL.n18 9.69747
R2191 VTAIL.n93 VTAIL.n8 9.69747
R2192 VTAIL.n313 VTAIL.n228 9.69747
R2193 VTAIL.n293 VTAIL.n238 9.69747
R2194 VTAIL.n266 VTAIL.n252 9.69747
R2195 VTAIL.n205 VTAIL.n120 9.69747
R2196 VTAIL.n185 VTAIL.n130 9.69747
R2197 VTAIL.n158 VTAIL.n144 9.69747
R2198 VTAIL.n424 VTAIL.n326 9.45567
R2199 VTAIL.n100 VTAIL.n2 9.45567
R2200 VTAIL.n320 VTAIL.n222 9.45567
R2201 VTAIL.n212 VTAIL.n114 9.45567
R2202 VTAIL.n407 VTAIL.n406 9.3005
R2203 VTAIL.n409 VTAIL.n408 9.3005
R2204 VTAIL.n334 VTAIL.n333 9.3005
R2205 VTAIL.n415 VTAIL.n414 9.3005
R2206 VTAIL.n417 VTAIL.n416 9.3005
R2207 VTAIL.n330 VTAIL.n329 9.3005
R2208 VTAIL.n423 VTAIL.n422 9.3005
R2209 VTAIL.n425 VTAIL.n424 9.3005
R2210 VTAIL.n401 VTAIL.n400 9.3005
R2211 VTAIL.n399 VTAIL.n398 9.3005
R2212 VTAIL.n342 VTAIL.n341 9.3005
R2213 VTAIL.n393 VTAIL.n392 9.3005
R2214 VTAIL.n391 VTAIL.n390 9.3005
R2215 VTAIL.n346 VTAIL.n345 9.3005
R2216 VTAIL.n385 VTAIL.n384 9.3005
R2217 VTAIL.n358 VTAIL.n357 9.3005
R2218 VTAIL.n365 VTAIL.n364 9.3005
R2219 VTAIL.n367 VTAIL.n366 9.3005
R2220 VTAIL.n354 VTAIL.n353 9.3005
R2221 VTAIL.n373 VTAIL.n372 9.3005
R2222 VTAIL.n375 VTAIL.n374 9.3005
R2223 VTAIL.n376 VTAIL.n349 9.3005
R2224 VTAIL.n383 VTAIL.n382 9.3005
R2225 VTAIL.n338 VTAIL.n337 9.3005
R2226 VTAIL.n83 VTAIL.n82 9.3005
R2227 VTAIL.n85 VTAIL.n84 9.3005
R2228 VTAIL.n10 VTAIL.n9 9.3005
R2229 VTAIL.n91 VTAIL.n90 9.3005
R2230 VTAIL.n93 VTAIL.n92 9.3005
R2231 VTAIL.n6 VTAIL.n5 9.3005
R2232 VTAIL.n99 VTAIL.n98 9.3005
R2233 VTAIL.n101 VTAIL.n100 9.3005
R2234 VTAIL.n77 VTAIL.n76 9.3005
R2235 VTAIL.n75 VTAIL.n74 9.3005
R2236 VTAIL.n18 VTAIL.n17 9.3005
R2237 VTAIL.n69 VTAIL.n68 9.3005
R2238 VTAIL.n67 VTAIL.n66 9.3005
R2239 VTAIL.n22 VTAIL.n21 9.3005
R2240 VTAIL.n61 VTAIL.n60 9.3005
R2241 VTAIL.n34 VTAIL.n33 9.3005
R2242 VTAIL.n41 VTAIL.n40 9.3005
R2243 VTAIL.n43 VTAIL.n42 9.3005
R2244 VTAIL.n30 VTAIL.n29 9.3005
R2245 VTAIL.n49 VTAIL.n48 9.3005
R2246 VTAIL.n51 VTAIL.n50 9.3005
R2247 VTAIL.n52 VTAIL.n25 9.3005
R2248 VTAIL.n59 VTAIL.n58 9.3005
R2249 VTAIL.n14 VTAIL.n13 9.3005
R2250 VTAIL.n321 VTAIL.n320 9.3005
R2251 VTAIL.n319 VTAIL.n318 9.3005
R2252 VTAIL.n226 VTAIL.n225 9.3005
R2253 VTAIL.n313 VTAIL.n312 9.3005
R2254 VTAIL.n311 VTAIL.n310 9.3005
R2255 VTAIL.n230 VTAIL.n229 9.3005
R2256 VTAIL.n305 VTAIL.n304 9.3005
R2257 VTAIL.n303 VTAIL.n302 9.3005
R2258 VTAIL.n234 VTAIL.n233 9.3005
R2259 VTAIL.n297 VTAIL.n296 9.3005
R2260 VTAIL.n295 VTAIL.n294 9.3005
R2261 VTAIL.n238 VTAIL.n237 9.3005
R2262 VTAIL.n289 VTAIL.n288 9.3005
R2263 VTAIL.n287 VTAIL.n286 9.3005
R2264 VTAIL.n242 VTAIL.n241 9.3005
R2265 VTAIL.n281 VTAIL.n280 9.3005
R2266 VTAIL.n279 VTAIL.n278 9.3005
R2267 VTAIL.n247 VTAIL.n245 9.3005
R2268 VTAIL.n273 VTAIL.n272 9.3005
R2269 VTAIL.n271 VTAIL.n270 9.3005
R2270 VTAIL.n252 VTAIL.n251 9.3005
R2271 VTAIL.n265 VTAIL.n264 9.3005
R2272 VTAIL.n263 VTAIL.n262 9.3005
R2273 VTAIL.n256 VTAIL.n255 9.3005
R2274 VTAIL.n148 VTAIL.n147 9.3005
R2275 VTAIL.n155 VTAIL.n154 9.3005
R2276 VTAIL.n157 VTAIL.n156 9.3005
R2277 VTAIL.n144 VTAIL.n143 9.3005
R2278 VTAIL.n163 VTAIL.n162 9.3005
R2279 VTAIL.n165 VTAIL.n164 9.3005
R2280 VTAIL.n139 VTAIL.n137 9.3005
R2281 VTAIL.n171 VTAIL.n170 9.3005
R2282 VTAIL.n197 VTAIL.n196 9.3005
R2283 VTAIL.n122 VTAIL.n121 9.3005
R2284 VTAIL.n203 VTAIL.n202 9.3005
R2285 VTAIL.n205 VTAIL.n204 9.3005
R2286 VTAIL.n118 VTAIL.n117 9.3005
R2287 VTAIL.n211 VTAIL.n210 9.3005
R2288 VTAIL.n213 VTAIL.n212 9.3005
R2289 VTAIL.n195 VTAIL.n194 9.3005
R2290 VTAIL.n126 VTAIL.n125 9.3005
R2291 VTAIL.n189 VTAIL.n188 9.3005
R2292 VTAIL.n187 VTAIL.n186 9.3005
R2293 VTAIL.n130 VTAIL.n129 9.3005
R2294 VTAIL.n181 VTAIL.n180 9.3005
R2295 VTAIL.n179 VTAIL.n178 9.3005
R2296 VTAIL.n134 VTAIL.n133 9.3005
R2297 VTAIL.n173 VTAIL.n172 9.3005
R2298 VTAIL.n367 VTAIL.n356 8.92171
R2299 VTAIL.n398 VTAIL.n340 8.92171
R2300 VTAIL.n414 VTAIL.n413 8.92171
R2301 VTAIL.n43 VTAIL.n32 8.92171
R2302 VTAIL.n74 VTAIL.n16 8.92171
R2303 VTAIL.n90 VTAIL.n89 8.92171
R2304 VTAIL.n310 VTAIL.n309 8.92171
R2305 VTAIL.n294 VTAIL.n236 8.92171
R2306 VTAIL.n265 VTAIL.n254 8.92171
R2307 VTAIL.n202 VTAIL.n201 8.92171
R2308 VTAIL.n186 VTAIL.n128 8.92171
R2309 VTAIL.n157 VTAIL.n146 8.92171
R2310 VTAIL.n364 VTAIL.n363 8.14595
R2311 VTAIL.n402 VTAIL.n401 8.14595
R2312 VTAIL.n410 VTAIL.n334 8.14595
R2313 VTAIL.n40 VTAIL.n39 8.14595
R2314 VTAIL.n78 VTAIL.n77 8.14595
R2315 VTAIL.n86 VTAIL.n10 8.14595
R2316 VTAIL.n306 VTAIL.n230 8.14595
R2317 VTAIL.n298 VTAIL.n297 8.14595
R2318 VTAIL.n262 VTAIL.n261 8.14595
R2319 VTAIL.n198 VTAIL.n122 8.14595
R2320 VTAIL.n190 VTAIL.n189 8.14595
R2321 VTAIL.n154 VTAIL.n153 8.14595
R2322 VTAIL.n360 VTAIL.n358 7.3702
R2323 VTAIL.n405 VTAIL.n338 7.3702
R2324 VTAIL.n409 VTAIL.n336 7.3702
R2325 VTAIL.n36 VTAIL.n34 7.3702
R2326 VTAIL.n81 VTAIL.n14 7.3702
R2327 VTAIL.n85 VTAIL.n12 7.3702
R2328 VTAIL.n305 VTAIL.n232 7.3702
R2329 VTAIL.n301 VTAIL.n234 7.3702
R2330 VTAIL.n258 VTAIL.n256 7.3702
R2331 VTAIL.n197 VTAIL.n124 7.3702
R2332 VTAIL.n193 VTAIL.n126 7.3702
R2333 VTAIL.n150 VTAIL.n148 7.3702
R2334 VTAIL.n406 VTAIL.n405 6.59444
R2335 VTAIL.n406 VTAIL.n336 6.59444
R2336 VTAIL.n82 VTAIL.n81 6.59444
R2337 VTAIL.n82 VTAIL.n12 6.59444
R2338 VTAIL.n302 VTAIL.n232 6.59444
R2339 VTAIL.n302 VTAIL.n301 6.59444
R2340 VTAIL.n194 VTAIL.n124 6.59444
R2341 VTAIL.n194 VTAIL.n193 6.59444
R2342 VTAIL.n363 VTAIL.n358 5.81868
R2343 VTAIL.n402 VTAIL.n338 5.81868
R2344 VTAIL.n410 VTAIL.n409 5.81868
R2345 VTAIL.n39 VTAIL.n34 5.81868
R2346 VTAIL.n78 VTAIL.n14 5.81868
R2347 VTAIL.n86 VTAIL.n85 5.81868
R2348 VTAIL.n306 VTAIL.n305 5.81868
R2349 VTAIL.n298 VTAIL.n234 5.81868
R2350 VTAIL.n261 VTAIL.n256 5.81868
R2351 VTAIL.n198 VTAIL.n197 5.81868
R2352 VTAIL.n190 VTAIL.n126 5.81868
R2353 VTAIL.n153 VTAIL.n148 5.81868
R2354 VTAIL.n364 VTAIL.n356 5.04292
R2355 VTAIL.n401 VTAIL.n340 5.04292
R2356 VTAIL.n413 VTAIL.n334 5.04292
R2357 VTAIL.n40 VTAIL.n32 5.04292
R2358 VTAIL.n77 VTAIL.n16 5.04292
R2359 VTAIL.n89 VTAIL.n10 5.04292
R2360 VTAIL.n309 VTAIL.n230 5.04292
R2361 VTAIL.n297 VTAIL.n236 5.04292
R2362 VTAIL.n262 VTAIL.n254 5.04292
R2363 VTAIL.n201 VTAIL.n122 5.04292
R2364 VTAIL.n189 VTAIL.n128 5.04292
R2365 VTAIL.n154 VTAIL.n146 5.04292
R2366 VTAIL.n368 VTAIL.n367 4.26717
R2367 VTAIL.n398 VTAIL.n397 4.26717
R2368 VTAIL.n414 VTAIL.n332 4.26717
R2369 VTAIL.n44 VTAIL.n43 4.26717
R2370 VTAIL.n74 VTAIL.n73 4.26717
R2371 VTAIL.n90 VTAIL.n8 4.26717
R2372 VTAIL.n310 VTAIL.n228 4.26717
R2373 VTAIL.n294 VTAIL.n293 4.26717
R2374 VTAIL.n266 VTAIL.n265 4.26717
R2375 VTAIL.n202 VTAIL.n120 4.26717
R2376 VTAIL.n186 VTAIL.n185 4.26717
R2377 VTAIL.n158 VTAIL.n157 4.26717
R2378 VTAIL.n371 VTAIL.n354 3.49141
R2379 VTAIL.n394 VTAIL.n342 3.49141
R2380 VTAIL.n418 VTAIL.n417 3.49141
R2381 VTAIL.n47 VTAIL.n30 3.49141
R2382 VTAIL.n70 VTAIL.n18 3.49141
R2383 VTAIL.n94 VTAIL.n93 3.49141
R2384 VTAIL.n314 VTAIL.n313 3.49141
R2385 VTAIL.n290 VTAIL.n238 3.49141
R2386 VTAIL.n269 VTAIL.n252 3.49141
R2387 VTAIL.n206 VTAIL.n205 3.49141
R2388 VTAIL.n182 VTAIL.n130 3.49141
R2389 VTAIL.n161 VTAIL.n144 3.49141
R2390 VTAIL.n359 VTAIL.n357 2.84303
R2391 VTAIL.n35 VTAIL.n33 2.84303
R2392 VTAIL.n257 VTAIL.n255 2.84303
R2393 VTAIL.n149 VTAIL.n147 2.84303
R2394 VTAIL.n372 VTAIL.n352 2.71565
R2395 VTAIL.n393 VTAIL.n344 2.71565
R2396 VTAIL.n421 VTAIL.n330 2.71565
R2397 VTAIL.n48 VTAIL.n28 2.71565
R2398 VTAIL.n69 VTAIL.n20 2.71565
R2399 VTAIL.n97 VTAIL.n6 2.71565
R2400 VTAIL.n317 VTAIL.n226 2.71565
R2401 VTAIL.n289 VTAIL.n240 2.71565
R2402 VTAIL.n270 VTAIL.n250 2.71565
R2403 VTAIL.n209 VTAIL.n118 2.71565
R2404 VTAIL.n181 VTAIL.n132 2.71565
R2405 VTAIL.n162 VTAIL.n142 2.71565
R2406 VTAIL.n377 VTAIL.n375 1.93989
R2407 VTAIL.n390 VTAIL.n389 1.93989
R2408 VTAIL.n422 VTAIL.n328 1.93989
R2409 VTAIL.n53 VTAIL.n51 1.93989
R2410 VTAIL.n66 VTAIL.n65 1.93989
R2411 VTAIL.n98 VTAIL.n4 1.93989
R2412 VTAIL.n318 VTAIL.n224 1.93989
R2413 VTAIL.n286 VTAIL.n285 1.93989
R2414 VTAIL.n274 VTAIL.n273 1.93989
R2415 VTAIL.n210 VTAIL.n116 1.93989
R2416 VTAIL.n178 VTAIL.n177 1.93989
R2417 VTAIL.n166 VTAIL.n165 1.93989
R2418 VTAIL.n376 VTAIL.n350 1.16414
R2419 VTAIL.n386 VTAIL.n346 1.16414
R2420 VTAIL.n426 VTAIL.n425 1.16414
R2421 VTAIL.n52 VTAIL.n26 1.16414
R2422 VTAIL.n62 VTAIL.n22 1.16414
R2423 VTAIL.n102 VTAIL.n101 1.16414
R2424 VTAIL.n322 VTAIL.n321 1.16414
R2425 VTAIL.n282 VTAIL.n242 1.16414
R2426 VTAIL.n277 VTAIL.n247 1.16414
R2427 VTAIL.n214 VTAIL.n213 1.16414
R2428 VTAIL.n174 VTAIL.n134 1.16414
R2429 VTAIL.n169 VTAIL.n139 1.16414
R2430 VTAIL.n430 VTAIL.t18 1.05594
R2431 VTAIL.n430 VTAIL.t17 1.05594
R2432 VTAIL.n0 VTAIL.t2 1.05594
R2433 VTAIL.n0 VTAIL.t5 1.05594
R2434 VTAIL.n106 VTAIL.t15 1.05594
R2435 VTAIL.n106 VTAIL.t16 1.05594
R2436 VTAIL.n108 VTAIL.t13 1.05594
R2437 VTAIL.n108 VTAIL.t14 1.05594
R2438 VTAIL.n220 VTAIL.t7 1.05594
R2439 VTAIL.n220 VTAIL.t9 1.05594
R2440 VTAIL.n218 VTAIL.t11 1.05594
R2441 VTAIL.n218 VTAIL.t12 1.05594
R2442 VTAIL.n112 VTAIL.t19 1.05594
R2443 VTAIL.n112 VTAIL.t3 1.05594
R2444 VTAIL.n110 VTAIL.t4 1.05594
R2445 VTAIL.n110 VTAIL.t6 1.05594
R2446 VTAIL.n219 VTAIL.n217 0.832397
R2447 VTAIL.n105 VTAIL.n1 0.832397
R2448 VTAIL.n113 VTAIL.n111 0.724638
R2449 VTAIL.n217 VTAIL.n113 0.724638
R2450 VTAIL.n221 VTAIL.n219 0.724638
R2451 VTAIL.n325 VTAIL.n221 0.724638
R2452 VTAIL.n109 VTAIL.n107 0.724638
R2453 VTAIL.n107 VTAIL.n105 0.724638
R2454 VTAIL.n431 VTAIL.n429 0.724638
R2455 VTAIL VTAIL.n1 0.601793
R2456 VTAIL.n382 VTAIL.n381 0.388379
R2457 VTAIL.n385 VTAIL.n348 0.388379
R2458 VTAIL.n428 VTAIL.n326 0.388379
R2459 VTAIL.n58 VTAIL.n57 0.388379
R2460 VTAIL.n61 VTAIL.n24 0.388379
R2461 VTAIL.n104 VTAIL.n2 0.388379
R2462 VTAIL.n324 VTAIL.n222 0.388379
R2463 VTAIL.n281 VTAIL.n244 0.388379
R2464 VTAIL.n278 VTAIL.n246 0.388379
R2465 VTAIL.n216 VTAIL.n114 0.388379
R2466 VTAIL.n173 VTAIL.n136 0.388379
R2467 VTAIL.n170 VTAIL.n138 0.388379
R2468 VTAIL.n365 VTAIL.n357 0.155672
R2469 VTAIL.n366 VTAIL.n365 0.155672
R2470 VTAIL.n366 VTAIL.n353 0.155672
R2471 VTAIL.n373 VTAIL.n353 0.155672
R2472 VTAIL.n374 VTAIL.n373 0.155672
R2473 VTAIL.n374 VTAIL.n349 0.155672
R2474 VTAIL.n383 VTAIL.n349 0.155672
R2475 VTAIL.n384 VTAIL.n383 0.155672
R2476 VTAIL.n384 VTAIL.n345 0.155672
R2477 VTAIL.n391 VTAIL.n345 0.155672
R2478 VTAIL.n392 VTAIL.n391 0.155672
R2479 VTAIL.n392 VTAIL.n341 0.155672
R2480 VTAIL.n399 VTAIL.n341 0.155672
R2481 VTAIL.n400 VTAIL.n399 0.155672
R2482 VTAIL.n400 VTAIL.n337 0.155672
R2483 VTAIL.n407 VTAIL.n337 0.155672
R2484 VTAIL.n408 VTAIL.n407 0.155672
R2485 VTAIL.n408 VTAIL.n333 0.155672
R2486 VTAIL.n415 VTAIL.n333 0.155672
R2487 VTAIL.n416 VTAIL.n415 0.155672
R2488 VTAIL.n416 VTAIL.n329 0.155672
R2489 VTAIL.n423 VTAIL.n329 0.155672
R2490 VTAIL.n424 VTAIL.n423 0.155672
R2491 VTAIL.n41 VTAIL.n33 0.155672
R2492 VTAIL.n42 VTAIL.n41 0.155672
R2493 VTAIL.n42 VTAIL.n29 0.155672
R2494 VTAIL.n49 VTAIL.n29 0.155672
R2495 VTAIL.n50 VTAIL.n49 0.155672
R2496 VTAIL.n50 VTAIL.n25 0.155672
R2497 VTAIL.n59 VTAIL.n25 0.155672
R2498 VTAIL.n60 VTAIL.n59 0.155672
R2499 VTAIL.n60 VTAIL.n21 0.155672
R2500 VTAIL.n67 VTAIL.n21 0.155672
R2501 VTAIL.n68 VTAIL.n67 0.155672
R2502 VTAIL.n68 VTAIL.n17 0.155672
R2503 VTAIL.n75 VTAIL.n17 0.155672
R2504 VTAIL.n76 VTAIL.n75 0.155672
R2505 VTAIL.n76 VTAIL.n13 0.155672
R2506 VTAIL.n83 VTAIL.n13 0.155672
R2507 VTAIL.n84 VTAIL.n83 0.155672
R2508 VTAIL.n84 VTAIL.n9 0.155672
R2509 VTAIL.n91 VTAIL.n9 0.155672
R2510 VTAIL.n92 VTAIL.n91 0.155672
R2511 VTAIL.n92 VTAIL.n5 0.155672
R2512 VTAIL.n99 VTAIL.n5 0.155672
R2513 VTAIL.n100 VTAIL.n99 0.155672
R2514 VTAIL.n320 VTAIL.n319 0.155672
R2515 VTAIL.n319 VTAIL.n225 0.155672
R2516 VTAIL.n312 VTAIL.n225 0.155672
R2517 VTAIL.n312 VTAIL.n311 0.155672
R2518 VTAIL.n311 VTAIL.n229 0.155672
R2519 VTAIL.n304 VTAIL.n229 0.155672
R2520 VTAIL.n304 VTAIL.n303 0.155672
R2521 VTAIL.n303 VTAIL.n233 0.155672
R2522 VTAIL.n296 VTAIL.n233 0.155672
R2523 VTAIL.n296 VTAIL.n295 0.155672
R2524 VTAIL.n295 VTAIL.n237 0.155672
R2525 VTAIL.n288 VTAIL.n237 0.155672
R2526 VTAIL.n288 VTAIL.n287 0.155672
R2527 VTAIL.n287 VTAIL.n241 0.155672
R2528 VTAIL.n280 VTAIL.n241 0.155672
R2529 VTAIL.n280 VTAIL.n279 0.155672
R2530 VTAIL.n279 VTAIL.n245 0.155672
R2531 VTAIL.n272 VTAIL.n245 0.155672
R2532 VTAIL.n272 VTAIL.n271 0.155672
R2533 VTAIL.n271 VTAIL.n251 0.155672
R2534 VTAIL.n264 VTAIL.n251 0.155672
R2535 VTAIL.n264 VTAIL.n263 0.155672
R2536 VTAIL.n263 VTAIL.n255 0.155672
R2537 VTAIL.n212 VTAIL.n211 0.155672
R2538 VTAIL.n211 VTAIL.n117 0.155672
R2539 VTAIL.n204 VTAIL.n117 0.155672
R2540 VTAIL.n204 VTAIL.n203 0.155672
R2541 VTAIL.n203 VTAIL.n121 0.155672
R2542 VTAIL.n196 VTAIL.n121 0.155672
R2543 VTAIL.n196 VTAIL.n195 0.155672
R2544 VTAIL.n195 VTAIL.n125 0.155672
R2545 VTAIL.n188 VTAIL.n125 0.155672
R2546 VTAIL.n188 VTAIL.n187 0.155672
R2547 VTAIL.n187 VTAIL.n129 0.155672
R2548 VTAIL.n180 VTAIL.n129 0.155672
R2549 VTAIL.n180 VTAIL.n179 0.155672
R2550 VTAIL.n179 VTAIL.n133 0.155672
R2551 VTAIL.n172 VTAIL.n133 0.155672
R2552 VTAIL.n172 VTAIL.n171 0.155672
R2553 VTAIL.n171 VTAIL.n137 0.155672
R2554 VTAIL.n164 VTAIL.n137 0.155672
R2555 VTAIL.n164 VTAIL.n163 0.155672
R2556 VTAIL.n163 VTAIL.n143 0.155672
R2557 VTAIL.n156 VTAIL.n143 0.155672
R2558 VTAIL.n156 VTAIL.n155 0.155672
R2559 VTAIL.n155 VTAIL.n147 0.155672
R2560 VTAIL VTAIL.n431 0.123345
R2561 VN.n2 VN.t2 985.455
R2562 VN.n14 VN.t4 985.455
R2563 VN.n3 VN.t3 964.472
R2564 VN.n1 VN.t6 964.472
R2565 VN.n9 VN.t7 964.472
R2566 VN.n10 VN.t9 964.472
R2567 VN.n15 VN.t1 964.472
R2568 VN.n13 VN.t0 964.472
R2569 VN.n21 VN.t8 964.472
R2570 VN.n22 VN.t5 964.472
R2571 VN.n11 VN.n10 161.3
R2572 VN.n23 VN.n22 161.3
R2573 VN.n21 VN.n12 161.3
R2574 VN.n20 VN.n19 161.3
R2575 VN.n18 VN.n13 161.3
R2576 VN.n17 VN.n16 161.3
R2577 VN.n9 VN.n0 161.3
R2578 VN.n8 VN.n7 161.3
R2579 VN.n6 VN.n1 161.3
R2580 VN.n5 VN.n4 161.3
R2581 VN.n17 VN.n14 70.4033
R2582 VN.n5 VN.n2 70.4033
R2583 VN.n10 VN.n9 48.2005
R2584 VN.n22 VN.n21 48.2005
R2585 VN VN.n23 47.2978
R2586 VN.n4 VN.n1 35.7853
R2587 VN.n8 VN.n1 35.7853
R2588 VN.n16 VN.n13 35.7853
R2589 VN.n20 VN.n13 35.7853
R2590 VN.n15 VN.n14 20.9576
R2591 VN.n3 VN.n2 20.9576
R2592 VN.n4 VN.n3 12.4157
R2593 VN.n9 VN.n8 12.4157
R2594 VN.n16 VN.n15 12.4157
R2595 VN.n21 VN.n20 12.4157
R2596 VN.n23 VN.n12 0.189894
R2597 VN.n19 VN.n12 0.189894
R2598 VN.n19 VN.n18 0.189894
R2599 VN.n18 VN.n17 0.189894
R2600 VN.n6 VN.n5 0.189894
R2601 VN.n7 VN.n6 0.189894
R2602 VN.n7 VN.n0 0.189894
R2603 VN.n11 VN.n0 0.189894
R2604 VN VN.n11 0.0516364
R2605 VDD2.n209 VDD2.n208 289.615
R2606 VDD2.n102 VDD2.n101 289.615
R2607 VDD2.n208 VDD2.n207 185
R2608 VDD2.n109 VDD2.n108 185
R2609 VDD2.n202 VDD2.n201 185
R2610 VDD2.n200 VDD2.n199 185
R2611 VDD2.n113 VDD2.n112 185
R2612 VDD2.n194 VDD2.n193 185
R2613 VDD2.n192 VDD2.n191 185
R2614 VDD2.n117 VDD2.n116 185
R2615 VDD2.n186 VDD2.n185 185
R2616 VDD2.n184 VDD2.n183 185
R2617 VDD2.n121 VDD2.n120 185
R2618 VDD2.n178 VDD2.n177 185
R2619 VDD2.n176 VDD2.n175 185
R2620 VDD2.n125 VDD2.n124 185
R2621 VDD2.n170 VDD2.n169 185
R2622 VDD2.n168 VDD2.n167 185
R2623 VDD2.n129 VDD2.n128 185
R2624 VDD2.n133 VDD2.n131 185
R2625 VDD2.n162 VDD2.n161 185
R2626 VDD2.n160 VDD2.n159 185
R2627 VDD2.n135 VDD2.n134 185
R2628 VDD2.n154 VDD2.n153 185
R2629 VDD2.n152 VDD2.n151 185
R2630 VDD2.n139 VDD2.n138 185
R2631 VDD2.n146 VDD2.n145 185
R2632 VDD2.n144 VDD2.n143 185
R2633 VDD2.n35 VDD2.n34 185
R2634 VDD2.n37 VDD2.n36 185
R2635 VDD2.n30 VDD2.n29 185
R2636 VDD2.n43 VDD2.n42 185
R2637 VDD2.n45 VDD2.n44 185
R2638 VDD2.n26 VDD2.n25 185
R2639 VDD2.n52 VDD2.n51 185
R2640 VDD2.n53 VDD2.n24 185
R2641 VDD2.n55 VDD2.n54 185
R2642 VDD2.n22 VDD2.n21 185
R2643 VDD2.n61 VDD2.n60 185
R2644 VDD2.n63 VDD2.n62 185
R2645 VDD2.n18 VDD2.n17 185
R2646 VDD2.n69 VDD2.n68 185
R2647 VDD2.n71 VDD2.n70 185
R2648 VDD2.n14 VDD2.n13 185
R2649 VDD2.n77 VDD2.n76 185
R2650 VDD2.n79 VDD2.n78 185
R2651 VDD2.n10 VDD2.n9 185
R2652 VDD2.n85 VDD2.n84 185
R2653 VDD2.n87 VDD2.n86 185
R2654 VDD2.n6 VDD2.n5 185
R2655 VDD2.n93 VDD2.n92 185
R2656 VDD2.n95 VDD2.n94 185
R2657 VDD2.n2 VDD2.n1 185
R2658 VDD2.n101 VDD2.n100 185
R2659 VDD2.n142 VDD2.t4 149.524
R2660 VDD2.n33 VDD2.t7 149.524
R2661 VDD2.n208 VDD2.n108 104.615
R2662 VDD2.n201 VDD2.n108 104.615
R2663 VDD2.n201 VDD2.n200 104.615
R2664 VDD2.n200 VDD2.n112 104.615
R2665 VDD2.n193 VDD2.n112 104.615
R2666 VDD2.n193 VDD2.n192 104.615
R2667 VDD2.n192 VDD2.n116 104.615
R2668 VDD2.n185 VDD2.n116 104.615
R2669 VDD2.n185 VDD2.n184 104.615
R2670 VDD2.n184 VDD2.n120 104.615
R2671 VDD2.n177 VDD2.n120 104.615
R2672 VDD2.n177 VDD2.n176 104.615
R2673 VDD2.n176 VDD2.n124 104.615
R2674 VDD2.n169 VDD2.n124 104.615
R2675 VDD2.n169 VDD2.n168 104.615
R2676 VDD2.n168 VDD2.n128 104.615
R2677 VDD2.n133 VDD2.n128 104.615
R2678 VDD2.n161 VDD2.n133 104.615
R2679 VDD2.n161 VDD2.n160 104.615
R2680 VDD2.n160 VDD2.n134 104.615
R2681 VDD2.n153 VDD2.n134 104.615
R2682 VDD2.n153 VDD2.n152 104.615
R2683 VDD2.n152 VDD2.n138 104.615
R2684 VDD2.n145 VDD2.n138 104.615
R2685 VDD2.n145 VDD2.n144 104.615
R2686 VDD2.n36 VDD2.n35 104.615
R2687 VDD2.n36 VDD2.n29 104.615
R2688 VDD2.n43 VDD2.n29 104.615
R2689 VDD2.n44 VDD2.n43 104.615
R2690 VDD2.n44 VDD2.n25 104.615
R2691 VDD2.n52 VDD2.n25 104.615
R2692 VDD2.n53 VDD2.n52 104.615
R2693 VDD2.n54 VDD2.n53 104.615
R2694 VDD2.n54 VDD2.n21 104.615
R2695 VDD2.n61 VDD2.n21 104.615
R2696 VDD2.n62 VDD2.n61 104.615
R2697 VDD2.n62 VDD2.n17 104.615
R2698 VDD2.n69 VDD2.n17 104.615
R2699 VDD2.n70 VDD2.n69 104.615
R2700 VDD2.n70 VDD2.n13 104.615
R2701 VDD2.n77 VDD2.n13 104.615
R2702 VDD2.n78 VDD2.n77 104.615
R2703 VDD2.n78 VDD2.n9 104.615
R2704 VDD2.n85 VDD2.n9 104.615
R2705 VDD2.n86 VDD2.n85 104.615
R2706 VDD2.n86 VDD2.n5 104.615
R2707 VDD2.n93 VDD2.n5 104.615
R2708 VDD2.n94 VDD2.n93 104.615
R2709 VDD2.n94 VDD2.n1 104.615
R2710 VDD2.n101 VDD2.n1 104.615
R2711 VDD2.n106 VDD2.n105 63.7589
R2712 VDD2 VDD2.n213 63.7559
R2713 VDD2.n212 VDD2.n211 63.2721
R2714 VDD2.n104 VDD2.n103 63.2711
R2715 VDD2.n144 VDD2.t4 52.3082
R2716 VDD2.n35 VDD2.t7 52.3082
R2717 VDD2.n104 VDD2.n102 52.3034
R2718 VDD2.n210 VDD2.n209 51.5793
R2719 VDD2.n210 VDD2.n106 43.3274
R2720 VDD2.n131 VDD2.n129 13.1884
R2721 VDD2.n55 VDD2.n22 13.1884
R2722 VDD2.n207 VDD2.n107 12.8005
R2723 VDD2.n167 VDD2.n166 12.8005
R2724 VDD2.n163 VDD2.n162 12.8005
R2725 VDD2.n56 VDD2.n24 12.8005
R2726 VDD2.n60 VDD2.n59 12.8005
R2727 VDD2.n100 VDD2.n0 12.8005
R2728 VDD2.n206 VDD2.n109 12.0247
R2729 VDD2.n170 VDD2.n127 12.0247
R2730 VDD2.n159 VDD2.n132 12.0247
R2731 VDD2.n51 VDD2.n50 12.0247
R2732 VDD2.n63 VDD2.n20 12.0247
R2733 VDD2.n99 VDD2.n2 12.0247
R2734 VDD2.n203 VDD2.n202 11.249
R2735 VDD2.n171 VDD2.n125 11.249
R2736 VDD2.n158 VDD2.n135 11.249
R2737 VDD2.n49 VDD2.n26 11.249
R2738 VDD2.n64 VDD2.n18 11.249
R2739 VDD2.n96 VDD2.n95 11.249
R2740 VDD2.n199 VDD2.n111 10.4732
R2741 VDD2.n175 VDD2.n174 10.4732
R2742 VDD2.n155 VDD2.n154 10.4732
R2743 VDD2.n46 VDD2.n45 10.4732
R2744 VDD2.n68 VDD2.n67 10.4732
R2745 VDD2.n92 VDD2.n4 10.4732
R2746 VDD2.n143 VDD2.n142 10.2747
R2747 VDD2.n34 VDD2.n33 10.2747
R2748 VDD2.n198 VDD2.n113 9.69747
R2749 VDD2.n178 VDD2.n123 9.69747
R2750 VDD2.n151 VDD2.n137 9.69747
R2751 VDD2.n42 VDD2.n28 9.69747
R2752 VDD2.n71 VDD2.n16 9.69747
R2753 VDD2.n91 VDD2.n6 9.69747
R2754 VDD2.n205 VDD2.n107 9.45567
R2755 VDD2.n98 VDD2.n0 9.45567
R2756 VDD2.n141 VDD2.n140 9.3005
R2757 VDD2.n148 VDD2.n147 9.3005
R2758 VDD2.n150 VDD2.n149 9.3005
R2759 VDD2.n137 VDD2.n136 9.3005
R2760 VDD2.n156 VDD2.n155 9.3005
R2761 VDD2.n158 VDD2.n157 9.3005
R2762 VDD2.n132 VDD2.n130 9.3005
R2763 VDD2.n164 VDD2.n163 9.3005
R2764 VDD2.n190 VDD2.n189 9.3005
R2765 VDD2.n115 VDD2.n114 9.3005
R2766 VDD2.n196 VDD2.n195 9.3005
R2767 VDD2.n198 VDD2.n197 9.3005
R2768 VDD2.n111 VDD2.n110 9.3005
R2769 VDD2.n204 VDD2.n203 9.3005
R2770 VDD2.n206 VDD2.n205 9.3005
R2771 VDD2.n188 VDD2.n187 9.3005
R2772 VDD2.n119 VDD2.n118 9.3005
R2773 VDD2.n182 VDD2.n181 9.3005
R2774 VDD2.n180 VDD2.n179 9.3005
R2775 VDD2.n123 VDD2.n122 9.3005
R2776 VDD2.n174 VDD2.n173 9.3005
R2777 VDD2.n172 VDD2.n171 9.3005
R2778 VDD2.n127 VDD2.n126 9.3005
R2779 VDD2.n166 VDD2.n165 9.3005
R2780 VDD2.n81 VDD2.n80 9.3005
R2781 VDD2.n83 VDD2.n82 9.3005
R2782 VDD2.n8 VDD2.n7 9.3005
R2783 VDD2.n89 VDD2.n88 9.3005
R2784 VDD2.n91 VDD2.n90 9.3005
R2785 VDD2.n4 VDD2.n3 9.3005
R2786 VDD2.n97 VDD2.n96 9.3005
R2787 VDD2.n99 VDD2.n98 9.3005
R2788 VDD2.n75 VDD2.n74 9.3005
R2789 VDD2.n73 VDD2.n72 9.3005
R2790 VDD2.n16 VDD2.n15 9.3005
R2791 VDD2.n67 VDD2.n66 9.3005
R2792 VDD2.n65 VDD2.n64 9.3005
R2793 VDD2.n20 VDD2.n19 9.3005
R2794 VDD2.n59 VDD2.n58 9.3005
R2795 VDD2.n32 VDD2.n31 9.3005
R2796 VDD2.n39 VDD2.n38 9.3005
R2797 VDD2.n41 VDD2.n40 9.3005
R2798 VDD2.n28 VDD2.n27 9.3005
R2799 VDD2.n47 VDD2.n46 9.3005
R2800 VDD2.n49 VDD2.n48 9.3005
R2801 VDD2.n50 VDD2.n23 9.3005
R2802 VDD2.n57 VDD2.n56 9.3005
R2803 VDD2.n12 VDD2.n11 9.3005
R2804 VDD2.n195 VDD2.n194 8.92171
R2805 VDD2.n179 VDD2.n121 8.92171
R2806 VDD2.n150 VDD2.n139 8.92171
R2807 VDD2.n41 VDD2.n30 8.92171
R2808 VDD2.n72 VDD2.n14 8.92171
R2809 VDD2.n88 VDD2.n87 8.92171
R2810 VDD2.n191 VDD2.n115 8.14595
R2811 VDD2.n183 VDD2.n182 8.14595
R2812 VDD2.n147 VDD2.n146 8.14595
R2813 VDD2.n38 VDD2.n37 8.14595
R2814 VDD2.n76 VDD2.n75 8.14595
R2815 VDD2.n84 VDD2.n8 8.14595
R2816 VDD2.n190 VDD2.n117 7.3702
R2817 VDD2.n186 VDD2.n119 7.3702
R2818 VDD2.n143 VDD2.n141 7.3702
R2819 VDD2.n34 VDD2.n32 7.3702
R2820 VDD2.n79 VDD2.n12 7.3702
R2821 VDD2.n83 VDD2.n10 7.3702
R2822 VDD2.n187 VDD2.n117 6.59444
R2823 VDD2.n187 VDD2.n186 6.59444
R2824 VDD2.n80 VDD2.n79 6.59444
R2825 VDD2.n80 VDD2.n10 6.59444
R2826 VDD2.n191 VDD2.n190 5.81868
R2827 VDD2.n183 VDD2.n119 5.81868
R2828 VDD2.n146 VDD2.n141 5.81868
R2829 VDD2.n37 VDD2.n32 5.81868
R2830 VDD2.n76 VDD2.n12 5.81868
R2831 VDD2.n84 VDD2.n83 5.81868
R2832 VDD2.n194 VDD2.n115 5.04292
R2833 VDD2.n182 VDD2.n121 5.04292
R2834 VDD2.n147 VDD2.n139 5.04292
R2835 VDD2.n38 VDD2.n30 5.04292
R2836 VDD2.n75 VDD2.n14 5.04292
R2837 VDD2.n87 VDD2.n8 5.04292
R2838 VDD2.n195 VDD2.n113 4.26717
R2839 VDD2.n179 VDD2.n178 4.26717
R2840 VDD2.n151 VDD2.n150 4.26717
R2841 VDD2.n42 VDD2.n41 4.26717
R2842 VDD2.n72 VDD2.n71 4.26717
R2843 VDD2.n88 VDD2.n6 4.26717
R2844 VDD2.n199 VDD2.n198 3.49141
R2845 VDD2.n175 VDD2.n123 3.49141
R2846 VDD2.n154 VDD2.n137 3.49141
R2847 VDD2.n45 VDD2.n28 3.49141
R2848 VDD2.n68 VDD2.n16 3.49141
R2849 VDD2.n92 VDD2.n91 3.49141
R2850 VDD2.n33 VDD2.n31 2.84303
R2851 VDD2.n142 VDD2.n140 2.84303
R2852 VDD2.n202 VDD2.n111 2.71565
R2853 VDD2.n174 VDD2.n125 2.71565
R2854 VDD2.n155 VDD2.n135 2.71565
R2855 VDD2.n46 VDD2.n26 2.71565
R2856 VDD2.n67 VDD2.n18 2.71565
R2857 VDD2.n95 VDD2.n4 2.71565
R2858 VDD2.n203 VDD2.n109 1.93989
R2859 VDD2.n171 VDD2.n170 1.93989
R2860 VDD2.n159 VDD2.n158 1.93989
R2861 VDD2.n51 VDD2.n49 1.93989
R2862 VDD2.n64 VDD2.n63 1.93989
R2863 VDD2.n96 VDD2.n2 1.93989
R2864 VDD2.n207 VDD2.n206 1.16414
R2865 VDD2.n167 VDD2.n127 1.16414
R2866 VDD2.n162 VDD2.n132 1.16414
R2867 VDD2.n50 VDD2.n24 1.16414
R2868 VDD2.n60 VDD2.n20 1.16414
R2869 VDD2.n100 VDD2.n99 1.16414
R2870 VDD2.n213 VDD2.t8 1.05594
R2871 VDD2.n213 VDD2.t5 1.05594
R2872 VDD2.n211 VDD2.t1 1.05594
R2873 VDD2.n211 VDD2.t9 1.05594
R2874 VDD2.n105 VDD2.t2 1.05594
R2875 VDD2.n105 VDD2.t0 1.05594
R2876 VDD2.n103 VDD2.t6 1.05594
R2877 VDD2.n103 VDD2.t3 1.05594
R2878 VDD2.n212 VDD2.n210 0.724638
R2879 VDD2.n209 VDD2.n107 0.388379
R2880 VDD2.n166 VDD2.n129 0.388379
R2881 VDD2.n163 VDD2.n131 0.388379
R2882 VDD2.n56 VDD2.n55 0.388379
R2883 VDD2.n59 VDD2.n22 0.388379
R2884 VDD2.n102 VDD2.n0 0.388379
R2885 VDD2 VDD2.n212 0.239724
R2886 VDD2.n205 VDD2.n204 0.155672
R2887 VDD2.n204 VDD2.n110 0.155672
R2888 VDD2.n197 VDD2.n110 0.155672
R2889 VDD2.n197 VDD2.n196 0.155672
R2890 VDD2.n196 VDD2.n114 0.155672
R2891 VDD2.n189 VDD2.n114 0.155672
R2892 VDD2.n189 VDD2.n188 0.155672
R2893 VDD2.n188 VDD2.n118 0.155672
R2894 VDD2.n181 VDD2.n118 0.155672
R2895 VDD2.n181 VDD2.n180 0.155672
R2896 VDD2.n180 VDD2.n122 0.155672
R2897 VDD2.n173 VDD2.n122 0.155672
R2898 VDD2.n173 VDD2.n172 0.155672
R2899 VDD2.n172 VDD2.n126 0.155672
R2900 VDD2.n165 VDD2.n126 0.155672
R2901 VDD2.n165 VDD2.n164 0.155672
R2902 VDD2.n164 VDD2.n130 0.155672
R2903 VDD2.n157 VDD2.n130 0.155672
R2904 VDD2.n157 VDD2.n156 0.155672
R2905 VDD2.n156 VDD2.n136 0.155672
R2906 VDD2.n149 VDD2.n136 0.155672
R2907 VDD2.n149 VDD2.n148 0.155672
R2908 VDD2.n148 VDD2.n140 0.155672
R2909 VDD2.n39 VDD2.n31 0.155672
R2910 VDD2.n40 VDD2.n39 0.155672
R2911 VDD2.n40 VDD2.n27 0.155672
R2912 VDD2.n47 VDD2.n27 0.155672
R2913 VDD2.n48 VDD2.n47 0.155672
R2914 VDD2.n48 VDD2.n23 0.155672
R2915 VDD2.n57 VDD2.n23 0.155672
R2916 VDD2.n58 VDD2.n57 0.155672
R2917 VDD2.n58 VDD2.n19 0.155672
R2918 VDD2.n65 VDD2.n19 0.155672
R2919 VDD2.n66 VDD2.n65 0.155672
R2920 VDD2.n66 VDD2.n15 0.155672
R2921 VDD2.n73 VDD2.n15 0.155672
R2922 VDD2.n74 VDD2.n73 0.155672
R2923 VDD2.n74 VDD2.n11 0.155672
R2924 VDD2.n81 VDD2.n11 0.155672
R2925 VDD2.n82 VDD2.n81 0.155672
R2926 VDD2.n82 VDD2.n7 0.155672
R2927 VDD2.n89 VDD2.n7 0.155672
R2928 VDD2.n90 VDD2.n89 0.155672
R2929 VDD2.n90 VDD2.n3 0.155672
R2930 VDD2.n97 VDD2.n3 0.155672
R2931 VDD2.n98 VDD2.n97 0.155672
R2932 VDD2.n106 VDD2.n104 0.126188
C0 VN VTAIL 7.96114f
C1 VDD1 VN 0.148217f
C2 VDD1 VTAIL 24.331f
C3 VDD2 VN 8.50316f
C4 VDD2 VTAIL 24.3588f
C5 VN VP 6.57199f
C6 VTAIL VP 7.97613f
C7 VDD1 VDD2 0.856267f
C8 VDD1 VP 8.66564f
C9 VDD2 VP 0.318183f
C10 VDD2 B 5.959951f
C11 VDD1 B 5.867868f
C12 VTAIL B 8.722138f
C13 VN B 9.50574f
C14 VP B 7.043589f
C15 VDD2.n0 B 0.014701f
C16 VDD2.n1 B 0.033172f
C17 VDD2.n2 B 0.01486f
C18 VDD2.n3 B 0.026118f
C19 VDD2.n4 B 0.014035f
C20 VDD2.n5 B 0.033172f
C21 VDD2.n6 B 0.01486f
C22 VDD2.n7 B 0.026118f
C23 VDD2.n8 B 0.014035f
C24 VDD2.n9 B 0.033172f
C25 VDD2.n10 B 0.01486f
C26 VDD2.n11 B 0.026118f
C27 VDD2.n12 B 0.014035f
C28 VDD2.n13 B 0.033172f
C29 VDD2.n14 B 0.01486f
C30 VDD2.n15 B 0.026118f
C31 VDD2.n16 B 0.014035f
C32 VDD2.n17 B 0.033172f
C33 VDD2.n18 B 0.01486f
C34 VDD2.n19 B 0.026118f
C35 VDD2.n20 B 0.014035f
C36 VDD2.n21 B 0.033172f
C37 VDD2.n22 B 0.014447f
C38 VDD2.n23 B 0.026118f
C39 VDD2.n24 B 0.01486f
C40 VDD2.n25 B 0.033172f
C41 VDD2.n26 B 0.01486f
C42 VDD2.n27 B 0.026118f
C43 VDD2.n28 B 0.014035f
C44 VDD2.n29 B 0.033172f
C45 VDD2.n30 B 0.01486f
C46 VDD2.n31 B 2.10288f
C47 VDD2.n32 B 0.014035f
C48 VDD2.t7 B 0.056977f
C49 VDD2.n33 B 0.256088f
C50 VDD2.n34 B 0.02345f
C51 VDD2.n35 B 0.024879f
C52 VDD2.n36 B 0.033172f
C53 VDD2.n37 B 0.01486f
C54 VDD2.n38 B 0.014035f
C55 VDD2.n39 B 0.026118f
C56 VDD2.n40 B 0.026118f
C57 VDD2.n41 B 0.014035f
C58 VDD2.n42 B 0.01486f
C59 VDD2.n43 B 0.033172f
C60 VDD2.n44 B 0.033172f
C61 VDD2.n45 B 0.01486f
C62 VDD2.n46 B 0.014035f
C63 VDD2.n47 B 0.026118f
C64 VDD2.n48 B 0.026118f
C65 VDD2.n49 B 0.014035f
C66 VDD2.n50 B 0.014035f
C67 VDD2.n51 B 0.01486f
C68 VDD2.n52 B 0.033172f
C69 VDD2.n53 B 0.033172f
C70 VDD2.n54 B 0.033172f
C71 VDD2.n55 B 0.014447f
C72 VDD2.n56 B 0.014035f
C73 VDD2.n57 B 0.026118f
C74 VDD2.n58 B 0.026118f
C75 VDD2.n59 B 0.014035f
C76 VDD2.n60 B 0.01486f
C77 VDD2.n61 B 0.033172f
C78 VDD2.n62 B 0.033172f
C79 VDD2.n63 B 0.01486f
C80 VDD2.n64 B 0.014035f
C81 VDD2.n65 B 0.026118f
C82 VDD2.n66 B 0.026118f
C83 VDD2.n67 B 0.014035f
C84 VDD2.n68 B 0.01486f
C85 VDD2.n69 B 0.033172f
C86 VDD2.n70 B 0.033172f
C87 VDD2.n71 B 0.01486f
C88 VDD2.n72 B 0.014035f
C89 VDD2.n73 B 0.026118f
C90 VDD2.n74 B 0.026118f
C91 VDD2.n75 B 0.014035f
C92 VDD2.n76 B 0.01486f
C93 VDD2.n77 B 0.033172f
C94 VDD2.n78 B 0.033172f
C95 VDD2.n79 B 0.01486f
C96 VDD2.n80 B 0.014035f
C97 VDD2.n81 B 0.026118f
C98 VDD2.n82 B 0.026118f
C99 VDD2.n83 B 0.014035f
C100 VDD2.n84 B 0.01486f
C101 VDD2.n85 B 0.033172f
C102 VDD2.n86 B 0.033172f
C103 VDD2.n87 B 0.01486f
C104 VDD2.n88 B 0.014035f
C105 VDD2.n89 B 0.026118f
C106 VDD2.n90 B 0.026118f
C107 VDD2.n91 B 0.014035f
C108 VDD2.n92 B 0.01486f
C109 VDD2.n93 B 0.033172f
C110 VDD2.n94 B 0.033172f
C111 VDD2.n95 B 0.01486f
C112 VDD2.n96 B 0.014035f
C113 VDD2.n97 B 0.026118f
C114 VDD2.n98 B 0.066078f
C115 VDD2.n99 B 0.014035f
C116 VDD2.n100 B 0.01486f
C117 VDD2.n101 B 0.066827f
C118 VDD2.n102 B 0.075394f
C119 VDD2.t6 B 0.387187f
C120 VDD2.t3 B 0.387187f
C121 VDD2.n103 B 3.54213f
C122 VDD2.n104 B 0.397318f
C123 VDD2.t2 B 0.387187f
C124 VDD2.t0 B 0.387187f
C125 VDD2.n105 B 3.54459f
C126 VDD2.n106 B 2.31238f
C127 VDD2.n107 B 0.014701f
C128 VDD2.n108 B 0.033172f
C129 VDD2.n109 B 0.01486f
C130 VDD2.n110 B 0.026118f
C131 VDD2.n111 B 0.014035f
C132 VDD2.n112 B 0.033172f
C133 VDD2.n113 B 0.01486f
C134 VDD2.n114 B 0.026118f
C135 VDD2.n115 B 0.014035f
C136 VDD2.n116 B 0.033172f
C137 VDD2.n117 B 0.01486f
C138 VDD2.n118 B 0.026118f
C139 VDD2.n119 B 0.014035f
C140 VDD2.n120 B 0.033172f
C141 VDD2.n121 B 0.01486f
C142 VDD2.n122 B 0.026118f
C143 VDD2.n123 B 0.014035f
C144 VDD2.n124 B 0.033172f
C145 VDD2.n125 B 0.01486f
C146 VDD2.n126 B 0.026118f
C147 VDD2.n127 B 0.014035f
C148 VDD2.n128 B 0.033172f
C149 VDD2.n129 B 0.014447f
C150 VDD2.n130 B 0.026118f
C151 VDD2.n131 B 0.014447f
C152 VDD2.n132 B 0.014035f
C153 VDD2.n133 B 0.033172f
C154 VDD2.n134 B 0.033172f
C155 VDD2.n135 B 0.01486f
C156 VDD2.n136 B 0.026118f
C157 VDD2.n137 B 0.014035f
C158 VDD2.n138 B 0.033172f
C159 VDD2.n139 B 0.01486f
C160 VDD2.n140 B 2.10288f
C161 VDD2.n141 B 0.014035f
C162 VDD2.t4 B 0.056977f
C163 VDD2.n142 B 0.256088f
C164 VDD2.n143 B 0.02345f
C165 VDD2.n144 B 0.024879f
C166 VDD2.n145 B 0.033172f
C167 VDD2.n146 B 0.01486f
C168 VDD2.n147 B 0.014035f
C169 VDD2.n148 B 0.026118f
C170 VDD2.n149 B 0.026118f
C171 VDD2.n150 B 0.014035f
C172 VDD2.n151 B 0.01486f
C173 VDD2.n152 B 0.033172f
C174 VDD2.n153 B 0.033172f
C175 VDD2.n154 B 0.01486f
C176 VDD2.n155 B 0.014035f
C177 VDD2.n156 B 0.026118f
C178 VDD2.n157 B 0.026118f
C179 VDD2.n158 B 0.014035f
C180 VDD2.n159 B 0.01486f
C181 VDD2.n160 B 0.033172f
C182 VDD2.n161 B 0.033172f
C183 VDD2.n162 B 0.01486f
C184 VDD2.n163 B 0.014035f
C185 VDD2.n164 B 0.026118f
C186 VDD2.n165 B 0.026118f
C187 VDD2.n166 B 0.014035f
C188 VDD2.n167 B 0.01486f
C189 VDD2.n168 B 0.033172f
C190 VDD2.n169 B 0.033172f
C191 VDD2.n170 B 0.01486f
C192 VDD2.n171 B 0.014035f
C193 VDD2.n172 B 0.026118f
C194 VDD2.n173 B 0.026118f
C195 VDD2.n174 B 0.014035f
C196 VDD2.n175 B 0.01486f
C197 VDD2.n176 B 0.033172f
C198 VDD2.n177 B 0.033172f
C199 VDD2.n178 B 0.01486f
C200 VDD2.n179 B 0.014035f
C201 VDD2.n180 B 0.026118f
C202 VDD2.n181 B 0.026118f
C203 VDD2.n182 B 0.014035f
C204 VDD2.n183 B 0.01486f
C205 VDD2.n184 B 0.033172f
C206 VDD2.n185 B 0.033172f
C207 VDD2.n186 B 0.01486f
C208 VDD2.n187 B 0.014035f
C209 VDD2.n188 B 0.026118f
C210 VDD2.n189 B 0.026118f
C211 VDD2.n190 B 0.014035f
C212 VDD2.n191 B 0.01486f
C213 VDD2.n192 B 0.033172f
C214 VDD2.n193 B 0.033172f
C215 VDD2.n194 B 0.01486f
C216 VDD2.n195 B 0.014035f
C217 VDD2.n196 B 0.026118f
C218 VDD2.n197 B 0.026118f
C219 VDD2.n198 B 0.014035f
C220 VDD2.n199 B 0.01486f
C221 VDD2.n200 B 0.033172f
C222 VDD2.n201 B 0.033172f
C223 VDD2.n202 B 0.01486f
C224 VDD2.n203 B 0.014035f
C225 VDD2.n204 B 0.026118f
C226 VDD2.n205 B 0.066078f
C227 VDD2.n206 B 0.014035f
C228 VDD2.n207 B 0.01486f
C229 VDD2.n208 B 0.066827f
C230 VDD2.n209 B 0.073815f
C231 VDD2.n210 B 2.72118f
C232 VDD2.t1 B 0.387187f
C233 VDD2.t9 B 0.387187f
C234 VDD2.n211 B 3.54212f
C235 VDD2.n212 B 0.289549f
C236 VDD2.t8 B 0.387187f
C237 VDD2.t5 B 0.387187f
C238 VDD2.n213 B 3.54456f
C239 VN.n0 B 0.047291f
C240 VN.t6 B 1.28264f
C241 VN.n1 B 0.490106f
C242 VN.t2 B 1.29298f
C243 VN.n2 B 0.475455f
C244 VN.t3 B 1.28264f
C245 VN.n3 B 0.48792f
C246 VN.n4 B 0.010731f
C247 VN.n5 B 0.152308f
C248 VN.n6 B 0.047291f
C249 VN.n7 B 0.047291f
C250 VN.n8 B 0.010731f
C251 VN.t7 B 1.28264f
C252 VN.n9 B 0.48792f
C253 VN.t9 B 1.28264f
C254 VN.n10 B 0.485441f
C255 VN.n11 B 0.036648f
C256 VN.n12 B 0.047291f
C257 VN.t0 B 1.28264f
C258 VN.n13 B 0.490106f
C259 VN.t4 B 1.29298f
C260 VN.n14 B 0.475455f
C261 VN.t1 B 1.28264f
C262 VN.n15 B 0.48792f
C263 VN.n16 B 0.010731f
C264 VN.n17 B 0.152308f
C265 VN.n18 B 0.047291f
C266 VN.n19 B 0.047291f
C267 VN.n20 B 0.010731f
C268 VN.t8 B 1.28264f
C269 VN.n21 B 0.48792f
C270 VN.t5 B 1.28264f
C271 VN.n22 B 0.485441f
C272 VN.n23 B 2.36352f
C273 VTAIL.t2 B 0.394603f
C274 VTAIL.t5 B 0.394603f
C275 VTAIL.n0 B 3.53574f
C276 VTAIL.n1 B 0.373448f
C277 VTAIL.n2 B 0.014983f
C278 VTAIL.n3 B 0.033808f
C279 VTAIL.n4 B 0.015145f
C280 VTAIL.n5 B 0.026618f
C281 VTAIL.n6 B 0.014303f
C282 VTAIL.n7 B 0.033808f
C283 VTAIL.n8 B 0.015145f
C284 VTAIL.n9 B 0.026618f
C285 VTAIL.n10 B 0.014303f
C286 VTAIL.n11 B 0.033808f
C287 VTAIL.n12 B 0.015145f
C288 VTAIL.n13 B 0.026618f
C289 VTAIL.n14 B 0.014303f
C290 VTAIL.n15 B 0.033808f
C291 VTAIL.n16 B 0.015145f
C292 VTAIL.n17 B 0.026618f
C293 VTAIL.n18 B 0.014303f
C294 VTAIL.n19 B 0.033808f
C295 VTAIL.n20 B 0.015145f
C296 VTAIL.n21 B 0.026618f
C297 VTAIL.n22 B 0.014303f
C298 VTAIL.n23 B 0.033808f
C299 VTAIL.n24 B 0.014724f
C300 VTAIL.n25 B 0.026618f
C301 VTAIL.n26 B 0.015145f
C302 VTAIL.n27 B 0.033808f
C303 VTAIL.n28 B 0.015145f
C304 VTAIL.n29 B 0.026618f
C305 VTAIL.n30 B 0.014303f
C306 VTAIL.n31 B 0.033808f
C307 VTAIL.n32 B 0.015145f
C308 VTAIL.n33 B 2.14316f
C309 VTAIL.n34 B 0.014303f
C310 VTAIL.t8 B 0.058068f
C311 VTAIL.n35 B 0.260993f
C312 VTAIL.n36 B 0.023899f
C313 VTAIL.n37 B 0.025356f
C314 VTAIL.n38 B 0.033808f
C315 VTAIL.n39 B 0.015145f
C316 VTAIL.n40 B 0.014303f
C317 VTAIL.n41 B 0.026618f
C318 VTAIL.n42 B 0.026618f
C319 VTAIL.n43 B 0.014303f
C320 VTAIL.n44 B 0.015145f
C321 VTAIL.n45 B 0.033808f
C322 VTAIL.n46 B 0.033808f
C323 VTAIL.n47 B 0.015145f
C324 VTAIL.n48 B 0.014303f
C325 VTAIL.n49 B 0.026618f
C326 VTAIL.n50 B 0.026618f
C327 VTAIL.n51 B 0.014303f
C328 VTAIL.n52 B 0.014303f
C329 VTAIL.n53 B 0.015145f
C330 VTAIL.n54 B 0.033808f
C331 VTAIL.n55 B 0.033808f
C332 VTAIL.n56 B 0.033808f
C333 VTAIL.n57 B 0.014724f
C334 VTAIL.n58 B 0.014303f
C335 VTAIL.n59 B 0.026618f
C336 VTAIL.n60 B 0.026618f
C337 VTAIL.n61 B 0.014303f
C338 VTAIL.n62 B 0.015145f
C339 VTAIL.n63 B 0.033808f
C340 VTAIL.n64 B 0.033808f
C341 VTAIL.n65 B 0.015145f
C342 VTAIL.n66 B 0.014303f
C343 VTAIL.n67 B 0.026618f
C344 VTAIL.n68 B 0.026618f
C345 VTAIL.n69 B 0.014303f
C346 VTAIL.n70 B 0.015145f
C347 VTAIL.n71 B 0.033808f
C348 VTAIL.n72 B 0.033808f
C349 VTAIL.n73 B 0.015145f
C350 VTAIL.n74 B 0.014303f
C351 VTAIL.n75 B 0.026618f
C352 VTAIL.n76 B 0.026618f
C353 VTAIL.n77 B 0.014303f
C354 VTAIL.n78 B 0.015145f
C355 VTAIL.n79 B 0.033808f
C356 VTAIL.n80 B 0.033808f
C357 VTAIL.n81 B 0.015145f
C358 VTAIL.n82 B 0.014303f
C359 VTAIL.n83 B 0.026618f
C360 VTAIL.n84 B 0.026618f
C361 VTAIL.n85 B 0.014303f
C362 VTAIL.n86 B 0.015145f
C363 VTAIL.n87 B 0.033808f
C364 VTAIL.n88 B 0.033808f
C365 VTAIL.n89 B 0.015145f
C366 VTAIL.n90 B 0.014303f
C367 VTAIL.n91 B 0.026618f
C368 VTAIL.n92 B 0.026618f
C369 VTAIL.n93 B 0.014303f
C370 VTAIL.n94 B 0.015145f
C371 VTAIL.n95 B 0.033808f
C372 VTAIL.n96 B 0.033808f
C373 VTAIL.n97 B 0.015145f
C374 VTAIL.n98 B 0.014303f
C375 VTAIL.n99 B 0.026618f
C376 VTAIL.n100 B 0.067344f
C377 VTAIL.n101 B 0.014303f
C378 VTAIL.n102 B 0.015145f
C379 VTAIL.n103 B 0.068107f
C380 VTAIL.n104 B 0.056886f
C381 VTAIL.n105 B 0.159072f
C382 VTAIL.t15 B 0.394603f
C383 VTAIL.t16 B 0.394603f
C384 VTAIL.n106 B 3.53574f
C385 VTAIL.n107 B 0.374742f
C386 VTAIL.t13 B 0.394603f
C387 VTAIL.t14 B 0.394603f
C388 VTAIL.n108 B 3.53574f
C389 VTAIL.n109 B 2.18551f
C390 VTAIL.t4 B 0.394603f
C391 VTAIL.t6 B 0.394603f
C392 VTAIL.n110 B 3.53573f
C393 VTAIL.n111 B 2.18552f
C394 VTAIL.t19 B 0.394603f
C395 VTAIL.t3 B 0.394603f
C396 VTAIL.n112 B 3.53573f
C397 VTAIL.n113 B 0.374751f
C398 VTAIL.n114 B 0.014983f
C399 VTAIL.n115 B 0.033808f
C400 VTAIL.n116 B 0.015145f
C401 VTAIL.n117 B 0.026618f
C402 VTAIL.n118 B 0.014303f
C403 VTAIL.n119 B 0.033808f
C404 VTAIL.n120 B 0.015145f
C405 VTAIL.n121 B 0.026618f
C406 VTAIL.n122 B 0.014303f
C407 VTAIL.n123 B 0.033808f
C408 VTAIL.n124 B 0.015145f
C409 VTAIL.n125 B 0.026618f
C410 VTAIL.n126 B 0.014303f
C411 VTAIL.n127 B 0.033808f
C412 VTAIL.n128 B 0.015145f
C413 VTAIL.n129 B 0.026618f
C414 VTAIL.n130 B 0.014303f
C415 VTAIL.n131 B 0.033808f
C416 VTAIL.n132 B 0.015145f
C417 VTAIL.n133 B 0.026618f
C418 VTAIL.n134 B 0.014303f
C419 VTAIL.n135 B 0.033808f
C420 VTAIL.n136 B 0.014724f
C421 VTAIL.n137 B 0.026618f
C422 VTAIL.n138 B 0.014724f
C423 VTAIL.n139 B 0.014303f
C424 VTAIL.n140 B 0.033808f
C425 VTAIL.n141 B 0.033808f
C426 VTAIL.n142 B 0.015145f
C427 VTAIL.n143 B 0.026618f
C428 VTAIL.n144 B 0.014303f
C429 VTAIL.n145 B 0.033808f
C430 VTAIL.n146 B 0.015145f
C431 VTAIL.n147 B 2.14316f
C432 VTAIL.n148 B 0.014303f
C433 VTAIL.t1 B 0.058068f
C434 VTAIL.n149 B 0.260993f
C435 VTAIL.n150 B 0.023899f
C436 VTAIL.n151 B 0.025356f
C437 VTAIL.n152 B 0.033808f
C438 VTAIL.n153 B 0.015145f
C439 VTAIL.n154 B 0.014303f
C440 VTAIL.n155 B 0.026618f
C441 VTAIL.n156 B 0.026618f
C442 VTAIL.n157 B 0.014303f
C443 VTAIL.n158 B 0.015145f
C444 VTAIL.n159 B 0.033808f
C445 VTAIL.n160 B 0.033808f
C446 VTAIL.n161 B 0.015145f
C447 VTAIL.n162 B 0.014303f
C448 VTAIL.n163 B 0.026618f
C449 VTAIL.n164 B 0.026618f
C450 VTAIL.n165 B 0.014303f
C451 VTAIL.n166 B 0.015145f
C452 VTAIL.n167 B 0.033808f
C453 VTAIL.n168 B 0.033808f
C454 VTAIL.n169 B 0.015145f
C455 VTAIL.n170 B 0.014303f
C456 VTAIL.n171 B 0.026618f
C457 VTAIL.n172 B 0.026618f
C458 VTAIL.n173 B 0.014303f
C459 VTAIL.n174 B 0.015145f
C460 VTAIL.n175 B 0.033808f
C461 VTAIL.n176 B 0.033808f
C462 VTAIL.n177 B 0.015145f
C463 VTAIL.n178 B 0.014303f
C464 VTAIL.n179 B 0.026618f
C465 VTAIL.n180 B 0.026618f
C466 VTAIL.n181 B 0.014303f
C467 VTAIL.n182 B 0.015145f
C468 VTAIL.n183 B 0.033808f
C469 VTAIL.n184 B 0.033808f
C470 VTAIL.n185 B 0.015145f
C471 VTAIL.n186 B 0.014303f
C472 VTAIL.n187 B 0.026618f
C473 VTAIL.n188 B 0.026618f
C474 VTAIL.n189 B 0.014303f
C475 VTAIL.n190 B 0.015145f
C476 VTAIL.n191 B 0.033808f
C477 VTAIL.n192 B 0.033808f
C478 VTAIL.n193 B 0.015145f
C479 VTAIL.n194 B 0.014303f
C480 VTAIL.n195 B 0.026618f
C481 VTAIL.n196 B 0.026618f
C482 VTAIL.n197 B 0.014303f
C483 VTAIL.n198 B 0.015145f
C484 VTAIL.n199 B 0.033808f
C485 VTAIL.n200 B 0.033808f
C486 VTAIL.n201 B 0.015145f
C487 VTAIL.n202 B 0.014303f
C488 VTAIL.n203 B 0.026618f
C489 VTAIL.n204 B 0.026618f
C490 VTAIL.n205 B 0.014303f
C491 VTAIL.n206 B 0.015145f
C492 VTAIL.n207 B 0.033808f
C493 VTAIL.n208 B 0.033808f
C494 VTAIL.n209 B 0.015145f
C495 VTAIL.n210 B 0.014303f
C496 VTAIL.n211 B 0.026618f
C497 VTAIL.n212 B 0.067344f
C498 VTAIL.n213 B 0.014303f
C499 VTAIL.n214 B 0.015145f
C500 VTAIL.n215 B 0.068107f
C501 VTAIL.n216 B 0.056886f
C502 VTAIL.n217 B 0.159072f
C503 VTAIL.t11 B 0.394603f
C504 VTAIL.t12 B 0.394603f
C505 VTAIL.n218 B 3.53573f
C506 VTAIL.n219 B 0.383993f
C507 VTAIL.t7 B 0.394603f
C508 VTAIL.t9 B 0.394603f
C509 VTAIL.n220 B 3.53573f
C510 VTAIL.n221 B 0.374751f
C511 VTAIL.n222 B 0.014983f
C512 VTAIL.n223 B 0.033808f
C513 VTAIL.n224 B 0.015145f
C514 VTAIL.n225 B 0.026618f
C515 VTAIL.n226 B 0.014303f
C516 VTAIL.n227 B 0.033808f
C517 VTAIL.n228 B 0.015145f
C518 VTAIL.n229 B 0.026618f
C519 VTAIL.n230 B 0.014303f
C520 VTAIL.n231 B 0.033808f
C521 VTAIL.n232 B 0.015145f
C522 VTAIL.n233 B 0.026618f
C523 VTAIL.n234 B 0.014303f
C524 VTAIL.n235 B 0.033808f
C525 VTAIL.n236 B 0.015145f
C526 VTAIL.n237 B 0.026618f
C527 VTAIL.n238 B 0.014303f
C528 VTAIL.n239 B 0.033808f
C529 VTAIL.n240 B 0.015145f
C530 VTAIL.n241 B 0.026618f
C531 VTAIL.n242 B 0.014303f
C532 VTAIL.n243 B 0.033808f
C533 VTAIL.n244 B 0.014724f
C534 VTAIL.n245 B 0.026618f
C535 VTAIL.n246 B 0.014724f
C536 VTAIL.n247 B 0.014303f
C537 VTAIL.n248 B 0.033808f
C538 VTAIL.n249 B 0.033808f
C539 VTAIL.n250 B 0.015145f
C540 VTAIL.n251 B 0.026618f
C541 VTAIL.n252 B 0.014303f
C542 VTAIL.n253 B 0.033808f
C543 VTAIL.n254 B 0.015145f
C544 VTAIL.n255 B 2.14316f
C545 VTAIL.n256 B 0.014303f
C546 VTAIL.t10 B 0.058068f
C547 VTAIL.n257 B 0.260993f
C548 VTAIL.n258 B 0.023899f
C549 VTAIL.n259 B 0.025356f
C550 VTAIL.n260 B 0.033808f
C551 VTAIL.n261 B 0.015145f
C552 VTAIL.n262 B 0.014303f
C553 VTAIL.n263 B 0.026618f
C554 VTAIL.n264 B 0.026618f
C555 VTAIL.n265 B 0.014303f
C556 VTAIL.n266 B 0.015145f
C557 VTAIL.n267 B 0.033808f
C558 VTAIL.n268 B 0.033808f
C559 VTAIL.n269 B 0.015145f
C560 VTAIL.n270 B 0.014303f
C561 VTAIL.n271 B 0.026618f
C562 VTAIL.n272 B 0.026618f
C563 VTAIL.n273 B 0.014303f
C564 VTAIL.n274 B 0.015145f
C565 VTAIL.n275 B 0.033808f
C566 VTAIL.n276 B 0.033808f
C567 VTAIL.n277 B 0.015145f
C568 VTAIL.n278 B 0.014303f
C569 VTAIL.n279 B 0.026618f
C570 VTAIL.n280 B 0.026618f
C571 VTAIL.n281 B 0.014303f
C572 VTAIL.n282 B 0.015145f
C573 VTAIL.n283 B 0.033808f
C574 VTAIL.n284 B 0.033808f
C575 VTAIL.n285 B 0.015145f
C576 VTAIL.n286 B 0.014303f
C577 VTAIL.n287 B 0.026618f
C578 VTAIL.n288 B 0.026618f
C579 VTAIL.n289 B 0.014303f
C580 VTAIL.n290 B 0.015145f
C581 VTAIL.n291 B 0.033808f
C582 VTAIL.n292 B 0.033808f
C583 VTAIL.n293 B 0.015145f
C584 VTAIL.n294 B 0.014303f
C585 VTAIL.n295 B 0.026618f
C586 VTAIL.n296 B 0.026618f
C587 VTAIL.n297 B 0.014303f
C588 VTAIL.n298 B 0.015145f
C589 VTAIL.n299 B 0.033808f
C590 VTAIL.n300 B 0.033808f
C591 VTAIL.n301 B 0.015145f
C592 VTAIL.n302 B 0.014303f
C593 VTAIL.n303 B 0.026618f
C594 VTAIL.n304 B 0.026618f
C595 VTAIL.n305 B 0.014303f
C596 VTAIL.n306 B 0.015145f
C597 VTAIL.n307 B 0.033808f
C598 VTAIL.n308 B 0.033808f
C599 VTAIL.n309 B 0.015145f
C600 VTAIL.n310 B 0.014303f
C601 VTAIL.n311 B 0.026618f
C602 VTAIL.n312 B 0.026618f
C603 VTAIL.n313 B 0.014303f
C604 VTAIL.n314 B 0.015145f
C605 VTAIL.n315 B 0.033808f
C606 VTAIL.n316 B 0.033808f
C607 VTAIL.n317 B 0.015145f
C608 VTAIL.n318 B 0.014303f
C609 VTAIL.n319 B 0.026618f
C610 VTAIL.n320 B 0.067344f
C611 VTAIL.n321 B 0.014303f
C612 VTAIL.n322 B 0.015145f
C613 VTAIL.n323 B 0.068107f
C614 VTAIL.n324 B 0.056886f
C615 VTAIL.n325 B 1.89849f
C616 VTAIL.n326 B 0.014983f
C617 VTAIL.n327 B 0.033808f
C618 VTAIL.n328 B 0.015145f
C619 VTAIL.n329 B 0.026618f
C620 VTAIL.n330 B 0.014303f
C621 VTAIL.n331 B 0.033808f
C622 VTAIL.n332 B 0.015145f
C623 VTAIL.n333 B 0.026618f
C624 VTAIL.n334 B 0.014303f
C625 VTAIL.n335 B 0.033808f
C626 VTAIL.n336 B 0.015145f
C627 VTAIL.n337 B 0.026618f
C628 VTAIL.n338 B 0.014303f
C629 VTAIL.n339 B 0.033808f
C630 VTAIL.n340 B 0.015145f
C631 VTAIL.n341 B 0.026618f
C632 VTAIL.n342 B 0.014303f
C633 VTAIL.n343 B 0.033808f
C634 VTAIL.n344 B 0.015145f
C635 VTAIL.n345 B 0.026618f
C636 VTAIL.n346 B 0.014303f
C637 VTAIL.n347 B 0.033808f
C638 VTAIL.n348 B 0.014724f
C639 VTAIL.n349 B 0.026618f
C640 VTAIL.n350 B 0.015145f
C641 VTAIL.n351 B 0.033808f
C642 VTAIL.n352 B 0.015145f
C643 VTAIL.n353 B 0.026618f
C644 VTAIL.n354 B 0.014303f
C645 VTAIL.n355 B 0.033808f
C646 VTAIL.n356 B 0.015145f
C647 VTAIL.n357 B 2.14316f
C648 VTAIL.n358 B 0.014303f
C649 VTAIL.t0 B 0.058068f
C650 VTAIL.n359 B 0.260993f
C651 VTAIL.n360 B 0.023899f
C652 VTAIL.n361 B 0.025356f
C653 VTAIL.n362 B 0.033808f
C654 VTAIL.n363 B 0.015145f
C655 VTAIL.n364 B 0.014303f
C656 VTAIL.n365 B 0.026618f
C657 VTAIL.n366 B 0.026618f
C658 VTAIL.n367 B 0.014303f
C659 VTAIL.n368 B 0.015145f
C660 VTAIL.n369 B 0.033808f
C661 VTAIL.n370 B 0.033808f
C662 VTAIL.n371 B 0.015145f
C663 VTAIL.n372 B 0.014303f
C664 VTAIL.n373 B 0.026618f
C665 VTAIL.n374 B 0.026618f
C666 VTAIL.n375 B 0.014303f
C667 VTAIL.n376 B 0.014303f
C668 VTAIL.n377 B 0.015145f
C669 VTAIL.n378 B 0.033808f
C670 VTAIL.n379 B 0.033808f
C671 VTAIL.n380 B 0.033808f
C672 VTAIL.n381 B 0.014724f
C673 VTAIL.n382 B 0.014303f
C674 VTAIL.n383 B 0.026618f
C675 VTAIL.n384 B 0.026618f
C676 VTAIL.n385 B 0.014303f
C677 VTAIL.n386 B 0.015145f
C678 VTAIL.n387 B 0.033808f
C679 VTAIL.n388 B 0.033808f
C680 VTAIL.n389 B 0.015145f
C681 VTAIL.n390 B 0.014303f
C682 VTAIL.n391 B 0.026618f
C683 VTAIL.n392 B 0.026618f
C684 VTAIL.n393 B 0.014303f
C685 VTAIL.n394 B 0.015145f
C686 VTAIL.n395 B 0.033808f
C687 VTAIL.n396 B 0.033808f
C688 VTAIL.n397 B 0.015145f
C689 VTAIL.n398 B 0.014303f
C690 VTAIL.n399 B 0.026618f
C691 VTAIL.n400 B 0.026618f
C692 VTAIL.n401 B 0.014303f
C693 VTAIL.n402 B 0.015145f
C694 VTAIL.n403 B 0.033808f
C695 VTAIL.n404 B 0.033808f
C696 VTAIL.n405 B 0.015145f
C697 VTAIL.n406 B 0.014303f
C698 VTAIL.n407 B 0.026618f
C699 VTAIL.n408 B 0.026618f
C700 VTAIL.n409 B 0.014303f
C701 VTAIL.n410 B 0.015145f
C702 VTAIL.n411 B 0.033808f
C703 VTAIL.n412 B 0.033808f
C704 VTAIL.n413 B 0.015145f
C705 VTAIL.n414 B 0.014303f
C706 VTAIL.n415 B 0.026618f
C707 VTAIL.n416 B 0.026618f
C708 VTAIL.n417 B 0.014303f
C709 VTAIL.n418 B 0.015145f
C710 VTAIL.n419 B 0.033808f
C711 VTAIL.n420 B 0.033808f
C712 VTAIL.n421 B 0.015145f
C713 VTAIL.n422 B 0.014303f
C714 VTAIL.n423 B 0.026618f
C715 VTAIL.n424 B 0.067344f
C716 VTAIL.n425 B 0.014303f
C717 VTAIL.n426 B 0.015145f
C718 VTAIL.n427 B 0.068107f
C719 VTAIL.n428 B 0.056886f
C720 VTAIL.n429 B 1.89849f
C721 VTAIL.t18 B 0.394603f
C722 VTAIL.t17 B 0.394603f
C723 VTAIL.n430 B 3.53574f
C724 VTAIL.n431 B 0.323169f
C725 VDD1.n0 B 0.014703f
C726 VDD1.n1 B 0.033176f
C727 VDD1.n2 B 0.014862f
C728 VDD1.n3 B 0.02612f
C729 VDD1.n4 B 0.014036f
C730 VDD1.n5 B 0.033176f
C731 VDD1.n6 B 0.014862f
C732 VDD1.n7 B 0.02612f
C733 VDD1.n8 B 0.014036f
C734 VDD1.n9 B 0.033176f
C735 VDD1.n10 B 0.014862f
C736 VDD1.n11 B 0.02612f
C737 VDD1.n12 B 0.014036f
C738 VDD1.n13 B 0.033176f
C739 VDD1.n14 B 0.014862f
C740 VDD1.n15 B 0.02612f
C741 VDD1.n16 B 0.014036f
C742 VDD1.n17 B 0.033176f
C743 VDD1.n18 B 0.014862f
C744 VDD1.n19 B 0.02612f
C745 VDD1.n20 B 0.014036f
C746 VDD1.n21 B 0.033176f
C747 VDD1.n22 B 0.014449f
C748 VDD1.n23 B 0.02612f
C749 VDD1.n24 B 0.014449f
C750 VDD1.n25 B 0.014036f
C751 VDD1.n26 B 0.033176f
C752 VDD1.n27 B 0.033176f
C753 VDD1.n28 B 0.014862f
C754 VDD1.n29 B 0.02612f
C755 VDD1.n30 B 0.014036f
C756 VDD1.n31 B 0.033176f
C757 VDD1.n32 B 0.014862f
C758 VDD1.n33 B 2.10311f
C759 VDD1.n34 B 0.014036f
C760 VDD1.t0 B 0.056983f
C761 VDD1.n35 B 0.256115f
C762 VDD1.n36 B 0.023453f
C763 VDD1.n37 B 0.024882f
C764 VDD1.n38 B 0.033176f
C765 VDD1.n39 B 0.014862f
C766 VDD1.n40 B 0.014036f
C767 VDD1.n41 B 0.02612f
C768 VDD1.n42 B 0.02612f
C769 VDD1.n43 B 0.014036f
C770 VDD1.n44 B 0.014862f
C771 VDD1.n45 B 0.033176f
C772 VDD1.n46 B 0.033176f
C773 VDD1.n47 B 0.014862f
C774 VDD1.n48 B 0.014036f
C775 VDD1.n49 B 0.02612f
C776 VDD1.n50 B 0.02612f
C777 VDD1.n51 B 0.014036f
C778 VDD1.n52 B 0.014862f
C779 VDD1.n53 B 0.033176f
C780 VDD1.n54 B 0.033176f
C781 VDD1.n55 B 0.014862f
C782 VDD1.n56 B 0.014036f
C783 VDD1.n57 B 0.02612f
C784 VDD1.n58 B 0.02612f
C785 VDD1.n59 B 0.014036f
C786 VDD1.n60 B 0.014862f
C787 VDD1.n61 B 0.033176f
C788 VDD1.n62 B 0.033176f
C789 VDD1.n63 B 0.014862f
C790 VDD1.n64 B 0.014036f
C791 VDD1.n65 B 0.02612f
C792 VDD1.n66 B 0.02612f
C793 VDD1.n67 B 0.014036f
C794 VDD1.n68 B 0.014862f
C795 VDD1.n69 B 0.033176f
C796 VDD1.n70 B 0.033176f
C797 VDD1.n71 B 0.014862f
C798 VDD1.n72 B 0.014036f
C799 VDD1.n73 B 0.02612f
C800 VDD1.n74 B 0.02612f
C801 VDD1.n75 B 0.014036f
C802 VDD1.n76 B 0.014862f
C803 VDD1.n77 B 0.033176f
C804 VDD1.n78 B 0.033176f
C805 VDD1.n79 B 0.014862f
C806 VDD1.n80 B 0.014036f
C807 VDD1.n81 B 0.02612f
C808 VDD1.n82 B 0.02612f
C809 VDD1.n83 B 0.014036f
C810 VDD1.n84 B 0.014862f
C811 VDD1.n85 B 0.033176f
C812 VDD1.n86 B 0.033176f
C813 VDD1.n87 B 0.014862f
C814 VDD1.n88 B 0.014036f
C815 VDD1.n89 B 0.02612f
C816 VDD1.n90 B 0.02612f
C817 VDD1.n91 B 0.014036f
C818 VDD1.n92 B 0.014862f
C819 VDD1.n93 B 0.033176f
C820 VDD1.n94 B 0.033176f
C821 VDD1.n95 B 0.014862f
C822 VDD1.n96 B 0.014036f
C823 VDD1.n97 B 0.02612f
C824 VDD1.n98 B 0.066085f
C825 VDD1.n99 B 0.014036f
C826 VDD1.n100 B 0.014862f
C827 VDD1.n101 B 0.066834f
C828 VDD1.n102 B 0.075402f
C829 VDD1.t2 B 0.387228f
C830 VDD1.t5 B 0.387228f
C831 VDD1.n103 B 3.5425f
C832 VDD1.n104 B 0.402106f
C833 VDD1.n105 B 0.014703f
C834 VDD1.n106 B 0.033176f
C835 VDD1.n107 B 0.014862f
C836 VDD1.n108 B 0.02612f
C837 VDD1.n109 B 0.014036f
C838 VDD1.n110 B 0.033176f
C839 VDD1.n111 B 0.014862f
C840 VDD1.n112 B 0.02612f
C841 VDD1.n113 B 0.014036f
C842 VDD1.n114 B 0.033176f
C843 VDD1.n115 B 0.014862f
C844 VDD1.n116 B 0.02612f
C845 VDD1.n117 B 0.014036f
C846 VDD1.n118 B 0.033176f
C847 VDD1.n119 B 0.014862f
C848 VDD1.n120 B 0.02612f
C849 VDD1.n121 B 0.014036f
C850 VDD1.n122 B 0.033176f
C851 VDD1.n123 B 0.014862f
C852 VDD1.n124 B 0.02612f
C853 VDD1.n125 B 0.014036f
C854 VDD1.n126 B 0.033176f
C855 VDD1.n127 B 0.014449f
C856 VDD1.n128 B 0.02612f
C857 VDD1.n129 B 0.014862f
C858 VDD1.n130 B 0.033176f
C859 VDD1.n131 B 0.014862f
C860 VDD1.n132 B 0.02612f
C861 VDD1.n133 B 0.014036f
C862 VDD1.n134 B 0.033176f
C863 VDD1.n135 B 0.014862f
C864 VDD1.n136 B 2.10311f
C865 VDD1.n137 B 0.014036f
C866 VDD1.t1 B 0.056983f
C867 VDD1.n138 B 0.256115f
C868 VDD1.n139 B 0.023453f
C869 VDD1.n140 B 0.024882f
C870 VDD1.n141 B 0.033176f
C871 VDD1.n142 B 0.014862f
C872 VDD1.n143 B 0.014036f
C873 VDD1.n144 B 0.02612f
C874 VDD1.n145 B 0.02612f
C875 VDD1.n146 B 0.014036f
C876 VDD1.n147 B 0.014862f
C877 VDD1.n148 B 0.033176f
C878 VDD1.n149 B 0.033176f
C879 VDD1.n150 B 0.014862f
C880 VDD1.n151 B 0.014036f
C881 VDD1.n152 B 0.02612f
C882 VDD1.n153 B 0.02612f
C883 VDD1.n154 B 0.014036f
C884 VDD1.n155 B 0.014036f
C885 VDD1.n156 B 0.014862f
C886 VDD1.n157 B 0.033176f
C887 VDD1.n158 B 0.033176f
C888 VDD1.n159 B 0.033176f
C889 VDD1.n160 B 0.014449f
C890 VDD1.n161 B 0.014036f
C891 VDD1.n162 B 0.02612f
C892 VDD1.n163 B 0.02612f
C893 VDD1.n164 B 0.014036f
C894 VDD1.n165 B 0.014862f
C895 VDD1.n166 B 0.033176f
C896 VDD1.n167 B 0.033176f
C897 VDD1.n168 B 0.014862f
C898 VDD1.n169 B 0.014036f
C899 VDD1.n170 B 0.02612f
C900 VDD1.n171 B 0.02612f
C901 VDD1.n172 B 0.014036f
C902 VDD1.n173 B 0.014862f
C903 VDD1.n174 B 0.033176f
C904 VDD1.n175 B 0.033176f
C905 VDD1.n176 B 0.014862f
C906 VDD1.n177 B 0.014036f
C907 VDD1.n178 B 0.02612f
C908 VDD1.n179 B 0.02612f
C909 VDD1.n180 B 0.014036f
C910 VDD1.n181 B 0.014862f
C911 VDD1.n182 B 0.033176f
C912 VDD1.n183 B 0.033176f
C913 VDD1.n184 B 0.014862f
C914 VDD1.n185 B 0.014036f
C915 VDD1.n186 B 0.02612f
C916 VDD1.n187 B 0.02612f
C917 VDD1.n188 B 0.014036f
C918 VDD1.n189 B 0.014862f
C919 VDD1.n190 B 0.033176f
C920 VDD1.n191 B 0.033176f
C921 VDD1.n192 B 0.014862f
C922 VDD1.n193 B 0.014036f
C923 VDD1.n194 B 0.02612f
C924 VDD1.n195 B 0.02612f
C925 VDD1.n196 B 0.014036f
C926 VDD1.n197 B 0.014862f
C927 VDD1.n198 B 0.033176f
C928 VDD1.n199 B 0.033176f
C929 VDD1.n200 B 0.014862f
C930 VDD1.n201 B 0.014036f
C931 VDD1.n202 B 0.02612f
C932 VDD1.n203 B 0.066085f
C933 VDD1.n204 B 0.014036f
C934 VDD1.n205 B 0.014862f
C935 VDD1.n206 B 0.066834f
C936 VDD1.n207 B 0.075402f
C937 VDD1.t3 B 0.387228f
C938 VDD1.t4 B 0.387228f
C939 VDD1.n208 B 3.54251f
C940 VDD1.n209 B 0.39736f
C941 VDD1.t7 B 0.387228f
C942 VDD1.t8 B 0.387228f
C943 VDD1.n210 B 3.54497f
C944 VDD1.n211 B 2.38988f
C945 VDD1.t6 B 0.387228f
C946 VDD1.t9 B 0.387228f
C947 VDD1.n212 B 3.5425f
C948 VDD1.n213 B 2.94737f
C949 VP.n0 B 0.047838f
C950 VP.t1 B 1.29748f
C951 VP.n1 B 0.495776f
C952 VP.n2 B 0.047838f
C953 VP.n3 B 0.047838f
C954 VP.t6 B 1.29748f
C955 VP.t7 B 1.29748f
C956 VP.t9 B 1.29748f
C957 VP.n4 B 0.495776f
C958 VP.t5 B 1.30794f
C959 VP.n5 B 0.480956f
C960 VP.t4 B 1.29748f
C961 VP.n6 B 0.493564f
C962 VP.n7 B 0.010855f
C963 VP.n8 B 0.15407f
C964 VP.n9 B 0.047838f
C965 VP.n10 B 0.047838f
C966 VP.n11 B 0.010855f
C967 VP.n12 B 0.493564f
C968 VP.n13 B 0.491057f
C969 VP.n14 B 2.35966f
C970 VP.n15 B 2.39621f
C971 VP.t3 B 1.29748f
C972 VP.n16 B 0.491057f
C973 VP.t2 B 1.29748f
C974 VP.n17 B 0.493564f
C975 VP.n18 B 0.010855f
C976 VP.n19 B 0.047838f
C977 VP.n20 B 0.047838f
C978 VP.n21 B 0.047838f
C979 VP.n22 B 0.010855f
C980 VP.t0 B 1.29748f
C981 VP.n23 B 0.493564f
C982 VP.t8 B 1.29748f
C983 VP.n24 B 0.491057f
C984 VP.n25 B 0.037072f
.ends

