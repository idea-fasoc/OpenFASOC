* NGSPICE file created from diff_pair_sample_1395.ext - technology: sky130A

.subckt diff_pair_sample_1395 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X1 B.t11 B.t9 B.t10 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=0 ps=0 w=6.32 l=0.54
X2 B.t8 B.t6 B.t7 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=0 ps=0 w=6.32 l=0.54
X3 VTAIL.t13 VP.t1 VDD1.t6 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X4 VDD1.t5 VP.t2 VTAIL.t12 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X5 B.t5 B.t3 B.t4 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=0 ps=0 w=6.32 l=0.54
X6 VTAIL.t3 VN.t0 VDD2.t7 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X7 VTAIL.t11 VP.t3 VDD1.t4 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=1.0428 ps=6.65 w=6.32 l=0.54
X8 VDD2.t6 VN.t1 VTAIL.t4 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=2.4648 ps=13.42 w=6.32 l=0.54
X9 VTAIL.t15 VP.t4 VDD1.t3 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=1.0428 ps=6.65 w=6.32 l=0.54
X10 B.t2 B.t0 B.t1 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=0 ps=0 w=6.32 l=0.54
X11 VTAIL.t5 VN.t2 VDD2.t5 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=1.0428 ps=6.65 w=6.32 l=0.54
X12 VDD1.t2 VP.t5 VTAIL.t10 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=2.4648 ps=13.42 w=6.32 l=0.54
X13 VTAIL.t2 VN.t3 VDD2.t4 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=2.4648 pd=13.42 as=1.0428 ps=6.65 w=6.32 l=0.54
X14 VDD2.t3 VN.t4 VTAIL.t1 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X15 VTAIL.t0 VN.t5 VDD2.t2 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X16 VDD2.t1 VN.t6 VTAIL.t7 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X17 VDD1.t1 VP.t6 VTAIL.t14 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=2.4648 ps=13.42 w=6.32 l=0.54
X18 VTAIL.t9 VP.t7 VDD1.t0 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=1.0428 ps=6.65 w=6.32 l=0.54
X19 VDD2.t0 VN.t7 VTAIL.t6 w_n1840_n2232# sky130_fd_pr__pfet_01v8 ad=1.0428 pd=6.65 as=2.4648 ps=13.42 w=6.32 l=0.54
R0 VP.n4 VP.t4 380.2
R1 VP.n11 VP.t3 354.807
R2 VP.n1 VP.t0 354.807
R3 VP.n16 VP.t1 354.807
R4 VP.n18 VP.t6 354.807
R5 VP.n8 VP.t5 354.807
R6 VP.n6 VP.t7 354.807
R7 VP.n5 VP.t2 354.807
R8 VP.n19 VP.n18 161.3
R9 VP.n6 VP.n3 161.3
R10 VP.n7 VP.n2 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n17 VP.n0 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n14 VP.n1 161.3
R15 VP.n13 VP.n12 161.3
R16 VP.n11 VP.n10 161.3
R17 VP.n16 VP.n1 48.2005
R18 VP.n6 VP.n5 48.2005
R19 VP.n4 VP.n3 45.0031
R20 VP.n12 VP.n11 41.6278
R21 VP.n18 VP.n17 41.6278
R22 VP.n8 VP.n7 41.6278
R23 VP.n10 VP.n9 36.9096
R24 VP.n5 VP.n4 15.6319
R25 VP.n12 VP.n1 6.57323
R26 VP.n17 VP.n16 6.57323
R27 VP.n7 VP.n6 6.57323
R28 VP.n3 VP.n2 0.189894
R29 VP.n9 VP.n2 0.189894
R30 VP.n13 VP.n10 0.189894
R31 VP.n14 VP.n13 0.189894
R32 VP.n15 VP.n14 0.189894
R33 VP.n15 VP.n0 0.189894
R34 VP.n19 VP.n0 0.189894
R35 VP VP.n19 0.0516364
R36 VTAIL.n11 VTAIL.t15 77.917
R37 VTAIL.n10 VTAIL.t4 77.917
R38 VTAIL.n7 VTAIL.t2 77.917
R39 VTAIL.n15 VTAIL.t6 77.9169
R40 VTAIL.n2 VTAIL.t5 77.9169
R41 VTAIL.n3 VTAIL.t14 77.9169
R42 VTAIL.n6 VTAIL.t11 77.9169
R43 VTAIL.n14 VTAIL.t10 77.9169
R44 VTAIL.n13 VTAIL.n12 72.7739
R45 VTAIL.n9 VTAIL.n8 72.7739
R46 VTAIL.n1 VTAIL.n0 72.7737
R47 VTAIL.n5 VTAIL.n4 72.7737
R48 VTAIL.n15 VTAIL.n14 18.5652
R49 VTAIL.n7 VTAIL.n6 18.5652
R50 VTAIL.n0 VTAIL.t1 5.1437
R51 VTAIL.n0 VTAIL.t0 5.1437
R52 VTAIL.n4 VTAIL.t8 5.1437
R53 VTAIL.n4 VTAIL.t13 5.1437
R54 VTAIL.n12 VTAIL.t12 5.1437
R55 VTAIL.n12 VTAIL.t9 5.1437
R56 VTAIL.n8 VTAIL.t7 5.1437
R57 VTAIL.n8 VTAIL.t3 5.1437
R58 VTAIL.n9 VTAIL.n7 0.7505
R59 VTAIL.n10 VTAIL.n9 0.7505
R60 VTAIL.n13 VTAIL.n11 0.7505
R61 VTAIL.n14 VTAIL.n13 0.7505
R62 VTAIL.n6 VTAIL.n5 0.7505
R63 VTAIL.n5 VTAIL.n3 0.7505
R64 VTAIL.n2 VTAIL.n1 0.7505
R65 VTAIL VTAIL.n15 0.69231
R66 VTAIL.n11 VTAIL.n10 0.470328
R67 VTAIL.n3 VTAIL.n2 0.470328
R68 VTAIL VTAIL.n1 0.0586897
R69 VDD1 VDD1.n0 89.8859
R70 VDD1.n3 VDD1.n2 89.7721
R71 VDD1.n3 VDD1.n1 89.7721
R72 VDD1.n5 VDD1.n4 89.4525
R73 VDD1.n5 VDD1.n3 33.1216
R74 VDD1.n4 VDD1.t0 5.1437
R75 VDD1.n4 VDD1.t2 5.1437
R76 VDD1.n0 VDD1.t3 5.1437
R77 VDD1.n0 VDD1.t5 5.1437
R78 VDD1.n2 VDD1.t6 5.1437
R79 VDD1.n2 VDD1.t1 5.1437
R80 VDD1.n1 VDD1.t4 5.1437
R81 VDD1.n1 VDD1.t7 5.1437
R82 VDD1 VDD1.n5 0.31731
R83 B.n297 B.n296 585
R84 B.n298 B.n45 585
R85 B.n300 B.n299 585
R86 B.n301 B.n44 585
R87 B.n303 B.n302 585
R88 B.n304 B.n43 585
R89 B.n306 B.n305 585
R90 B.n307 B.n42 585
R91 B.n309 B.n308 585
R92 B.n310 B.n41 585
R93 B.n312 B.n311 585
R94 B.n313 B.n40 585
R95 B.n315 B.n314 585
R96 B.n316 B.n39 585
R97 B.n318 B.n317 585
R98 B.n319 B.n38 585
R99 B.n321 B.n320 585
R100 B.n322 B.n37 585
R101 B.n324 B.n323 585
R102 B.n325 B.n36 585
R103 B.n327 B.n326 585
R104 B.n328 B.n35 585
R105 B.n330 B.n329 585
R106 B.n331 B.n34 585
R107 B.n333 B.n332 585
R108 B.n335 B.n31 585
R109 B.n337 B.n336 585
R110 B.n338 B.n30 585
R111 B.n340 B.n339 585
R112 B.n341 B.n29 585
R113 B.n343 B.n342 585
R114 B.n344 B.n28 585
R115 B.n346 B.n345 585
R116 B.n347 B.n25 585
R117 B.n350 B.n349 585
R118 B.n351 B.n24 585
R119 B.n353 B.n352 585
R120 B.n354 B.n23 585
R121 B.n356 B.n355 585
R122 B.n357 B.n22 585
R123 B.n359 B.n358 585
R124 B.n360 B.n21 585
R125 B.n362 B.n361 585
R126 B.n363 B.n20 585
R127 B.n365 B.n364 585
R128 B.n366 B.n19 585
R129 B.n368 B.n367 585
R130 B.n369 B.n18 585
R131 B.n371 B.n370 585
R132 B.n372 B.n17 585
R133 B.n374 B.n373 585
R134 B.n375 B.n16 585
R135 B.n377 B.n376 585
R136 B.n378 B.n15 585
R137 B.n380 B.n379 585
R138 B.n381 B.n14 585
R139 B.n383 B.n382 585
R140 B.n384 B.n13 585
R141 B.n386 B.n385 585
R142 B.n295 B.n46 585
R143 B.n294 B.n293 585
R144 B.n292 B.n47 585
R145 B.n291 B.n290 585
R146 B.n289 B.n48 585
R147 B.n288 B.n287 585
R148 B.n286 B.n49 585
R149 B.n285 B.n284 585
R150 B.n283 B.n50 585
R151 B.n282 B.n281 585
R152 B.n280 B.n51 585
R153 B.n279 B.n278 585
R154 B.n277 B.n52 585
R155 B.n276 B.n275 585
R156 B.n274 B.n53 585
R157 B.n273 B.n272 585
R158 B.n271 B.n54 585
R159 B.n270 B.n269 585
R160 B.n268 B.n55 585
R161 B.n267 B.n266 585
R162 B.n265 B.n56 585
R163 B.n264 B.n263 585
R164 B.n262 B.n57 585
R165 B.n261 B.n260 585
R166 B.n259 B.n58 585
R167 B.n258 B.n257 585
R168 B.n256 B.n59 585
R169 B.n255 B.n254 585
R170 B.n253 B.n60 585
R171 B.n252 B.n251 585
R172 B.n250 B.n61 585
R173 B.n249 B.n248 585
R174 B.n247 B.n62 585
R175 B.n246 B.n245 585
R176 B.n244 B.n63 585
R177 B.n243 B.n242 585
R178 B.n241 B.n64 585
R179 B.n240 B.n239 585
R180 B.n238 B.n65 585
R181 B.n237 B.n236 585
R182 B.n235 B.n66 585
R183 B.n234 B.n233 585
R184 B.n232 B.n67 585
R185 B.n142 B.n101 585
R186 B.n144 B.n143 585
R187 B.n145 B.n100 585
R188 B.n147 B.n146 585
R189 B.n148 B.n99 585
R190 B.n150 B.n149 585
R191 B.n151 B.n98 585
R192 B.n153 B.n152 585
R193 B.n154 B.n97 585
R194 B.n156 B.n155 585
R195 B.n157 B.n96 585
R196 B.n159 B.n158 585
R197 B.n160 B.n95 585
R198 B.n162 B.n161 585
R199 B.n163 B.n94 585
R200 B.n165 B.n164 585
R201 B.n166 B.n93 585
R202 B.n168 B.n167 585
R203 B.n169 B.n92 585
R204 B.n171 B.n170 585
R205 B.n172 B.n91 585
R206 B.n174 B.n173 585
R207 B.n175 B.n90 585
R208 B.n177 B.n176 585
R209 B.n178 B.n87 585
R210 B.n181 B.n180 585
R211 B.n182 B.n86 585
R212 B.n184 B.n183 585
R213 B.n185 B.n85 585
R214 B.n187 B.n186 585
R215 B.n188 B.n84 585
R216 B.n190 B.n189 585
R217 B.n191 B.n83 585
R218 B.n193 B.n192 585
R219 B.n195 B.n194 585
R220 B.n196 B.n79 585
R221 B.n198 B.n197 585
R222 B.n199 B.n78 585
R223 B.n201 B.n200 585
R224 B.n202 B.n77 585
R225 B.n204 B.n203 585
R226 B.n205 B.n76 585
R227 B.n207 B.n206 585
R228 B.n208 B.n75 585
R229 B.n210 B.n209 585
R230 B.n211 B.n74 585
R231 B.n213 B.n212 585
R232 B.n214 B.n73 585
R233 B.n216 B.n215 585
R234 B.n217 B.n72 585
R235 B.n219 B.n218 585
R236 B.n220 B.n71 585
R237 B.n222 B.n221 585
R238 B.n223 B.n70 585
R239 B.n225 B.n224 585
R240 B.n226 B.n69 585
R241 B.n228 B.n227 585
R242 B.n229 B.n68 585
R243 B.n231 B.n230 585
R244 B.n141 B.n140 585
R245 B.n139 B.n102 585
R246 B.n138 B.n137 585
R247 B.n136 B.n103 585
R248 B.n135 B.n134 585
R249 B.n133 B.n104 585
R250 B.n132 B.n131 585
R251 B.n130 B.n105 585
R252 B.n129 B.n128 585
R253 B.n127 B.n106 585
R254 B.n126 B.n125 585
R255 B.n124 B.n107 585
R256 B.n123 B.n122 585
R257 B.n121 B.n108 585
R258 B.n120 B.n119 585
R259 B.n118 B.n109 585
R260 B.n117 B.n116 585
R261 B.n115 B.n110 585
R262 B.n114 B.n113 585
R263 B.n112 B.n111 585
R264 B.n2 B.n0 585
R265 B.n417 B.n1 585
R266 B.n416 B.n415 585
R267 B.n414 B.n3 585
R268 B.n413 B.n412 585
R269 B.n411 B.n4 585
R270 B.n410 B.n409 585
R271 B.n408 B.n5 585
R272 B.n407 B.n406 585
R273 B.n405 B.n6 585
R274 B.n404 B.n403 585
R275 B.n402 B.n7 585
R276 B.n401 B.n400 585
R277 B.n399 B.n8 585
R278 B.n398 B.n397 585
R279 B.n396 B.n9 585
R280 B.n395 B.n394 585
R281 B.n393 B.n10 585
R282 B.n392 B.n391 585
R283 B.n390 B.n11 585
R284 B.n389 B.n388 585
R285 B.n387 B.n12 585
R286 B.n419 B.n418 585
R287 B.n140 B.n101 516.524
R288 B.n387 B.n386 516.524
R289 B.n230 B.n67 516.524
R290 B.n296 B.n295 516.524
R291 B.n80 B.t0 487.575
R292 B.n88 B.t3 487.575
R293 B.n26 B.t9 487.575
R294 B.n32 B.t6 487.575
R295 B.n140 B.n139 163.367
R296 B.n139 B.n138 163.367
R297 B.n138 B.n103 163.367
R298 B.n134 B.n103 163.367
R299 B.n134 B.n133 163.367
R300 B.n133 B.n132 163.367
R301 B.n132 B.n105 163.367
R302 B.n128 B.n105 163.367
R303 B.n128 B.n127 163.367
R304 B.n127 B.n126 163.367
R305 B.n126 B.n107 163.367
R306 B.n122 B.n107 163.367
R307 B.n122 B.n121 163.367
R308 B.n121 B.n120 163.367
R309 B.n120 B.n109 163.367
R310 B.n116 B.n109 163.367
R311 B.n116 B.n115 163.367
R312 B.n115 B.n114 163.367
R313 B.n114 B.n111 163.367
R314 B.n111 B.n2 163.367
R315 B.n418 B.n2 163.367
R316 B.n418 B.n417 163.367
R317 B.n417 B.n416 163.367
R318 B.n416 B.n3 163.367
R319 B.n412 B.n3 163.367
R320 B.n412 B.n411 163.367
R321 B.n411 B.n410 163.367
R322 B.n410 B.n5 163.367
R323 B.n406 B.n5 163.367
R324 B.n406 B.n405 163.367
R325 B.n405 B.n404 163.367
R326 B.n404 B.n7 163.367
R327 B.n400 B.n7 163.367
R328 B.n400 B.n399 163.367
R329 B.n399 B.n398 163.367
R330 B.n398 B.n9 163.367
R331 B.n394 B.n9 163.367
R332 B.n394 B.n393 163.367
R333 B.n393 B.n392 163.367
R334 B.n392 B.n11 163.367
R335 B.n388 B.n11 163.367
R336 B.n388 B.n387 163.367
R337 B.n144 B.n101 163.367
R338 B.n145 B.n144 163.367
R339 B.n146 B.n145 163.367
R340 B.n146 B.n99 163.367
R341 B.n150 B.n99 163.367
R342 B.n151 B.n150 163.367
R343 B.n152 B.n151 163.367
R344 B.n152 B.n97 163.367
R345 B.n156 B.n97 163.367
R346 B.n157 B.n156 163.367
R347 B.n158 B.n157 163.367
R348 B.n158 B.n95 163.367
R349 B.n162 B.n95 163.367
R350 B.n163 B.n162 163.367
R351 B.n164 B.n163 163.367
R352 B.n164 B.n93 163.367
R353 B.n168 B.n93 163.367
R354 B.n169 B.n168 163.367
R355 B.n170 B.n169 163.367
R356 B.n170 B.n91 163.367
R357 B.n174 B.n91 163.367
R358 B.n175 B.n174 163.367
R359 B.n176 B.n175 163.367
R360 B.n176 B.n87 163.367
R361 B.n181 B.n87 163.367
R362 B.n182 B.n181 163.367
R363 B.n183 B.n182 163.367
R364 B.n183 B.n85 163.367
R365 B.n187 B.n85 163.367
R366 B.n188 B.n187 163.367
R367 B.n189 B.n188 163.367
R368 B.n189 B.n83 163.367
R369 B.n193 B.n83 163.367
R370 B.n194 B.n193 163.367
R371 B.n194 B.n79 163.367
R372 B.n198 B.n79 163.367
R373 B.n199 B.n198 163.367
R374 B.n200 B.n199 163.367
R375 B.n200 B.n77 163.367
R376 B.n204 B.n77 163.367
R377 B.n205 B.n204 163.367
R378 B.n206 B.n205 163.367
R379 B.n206 B.n75 163.367
R380 B.n210 B.n75 163.367
R381 B.n211 B.n210 163.367
R382 B.n212 B.n211 163.367
R383 B.n212 B.n73 163.367
R384 B.n216 B.n73 163.367
R385 B.n217 B.n216 163.367
R386 B.n218 B.n217 163.367
R387 B.n218 B.n71 163.367
R388 B.n222 B.n71 163.367
R389 B.n223 B.n222 163.367
R390 B.n224 B.n223 163.367
R391 B.n224 B.n69 163.367
R392 B.n228 B.n69 163.367
R393 B.n229 B.n228 163.367
R394 B.n230 B.n229 163.367
R395 B.n234 B.n67 163.367
R396 B.n235 B.n234 163.367
R397 B.n236 B.n235 163.367
R398 B.n236 B.n65 163.367
R399 B.n240 B.n65 163.367
R400 B.n241 B.n240 163.367
R401 B.n242 B.n241 163.367
R402 B.n242 B.n63 163.367
R403 B.n246 B.n63 163.367
R404 B.n247 B.n246 163.367
R405 B.n248 B.n247 163.367
R406 B.n248 B.n61 163.367
R407 B.n252 B.n61 163.367
R408 B.n253 B.n252 163.367
R409 B.n254 B.n253 163.367
R410 B.n254 B.n59 163.367
R411 B.n258 B.n59 163.367
R412 B.n259 B.n258 163.367
R413 B.n260 B.n259 163.367
R414 B.n260 B.n57 163.367
R415 B.n264 B.n57 163.367
R416 B.n265 B.n264 163.367
R417 B.n266 B.n265 163.367
R418 B.n266 B.n55 163.367
R419 B.n270 B.n55 163.367
R420 B.n271 B.n270 163.367
R421 B.n272 B.n271 163.367
R422 B.n272 B.n53 163.367
R423 B.n276 B.n53 163.367
R424 B.n277 B.n276 163.367
R425 B.n278 B.n277 163.367
R426 B.n278 B.n51 163.367
R427 B.n282 B.n51 163.367
R428 B.n283 B.n282 163.367
R429 B.n284 B.n283 163.367
R430 B.n284 B.n49 163.367
R431 B.n288 B.n49 163.367
R432 B.n289 B.n288 163.367
R433 B.n290 B.n289 163.367
R434 B.n290 B.n47 163.367
R435 B.n294 B.n47 163.367
R436 B.n295 B.n294 163.367
R437 B.n386 B.n13 163.367
R438 B.n382 B.n13 163.367
R439 B.n382 B.n381 163.367
R440 B.n381 B.n380 163.367
R441 B.n380 B.n15 163.367
R442 B.n376 B.n15 163.367
R443 B.n376 B.n375 163.367
R444 B.n375 B.n374 163.367
R445 B.n374 B.n17 163.367
R446 B.n370 B.n17 163.367
R447 B.n370 B.n369 163.367
R448 B.n369 B.n368 163.367
R449 B.n368 B.n19 163.367
R450 B.n364 B.n19 163.367
R451 B.n364 B.n363 163.367
R452 B.n363 B.n362 163.367
R453 B.n362 B.n21 163.367
R454 B.n358 B.n21 163.367
R455 B.n358 B.n357 163.367
R456 B.n357 B.n356 163.367
R457 B.n356 B.n23 163.367
R458 B.n352 B.n23 163.367
R459 B.n352 B.n351 163.367
R460 B.n351 B.n350 163.367
R461 B.n350 B.n25 163.367
R462 B.n345 B.n25 163.367
R463 B.n345 B.n344 163.367
R464 B.n344 B.n343 163.367
R465 B.n343 B.n29 163.367
R466 B.n339 B.n29 163.367
R467 B.n339 B.n338 163.367
R468 B.n338 B.n337 163.367
R469 B.n337 B.n31 163.367
R470 B.n332 B.n31 163.367
R471 B.n332 B.n331 163.367
R472 B.n331 B.n330 163.367
R473 B.n330 B.n35 163.367
R474 B.n326 B.n35 163.367
R475 B.n326 B.n325 163.367
R476 B.n325 B.n324 163.367
R477 B.n324 B.n37 163.367
R478 B.n320 B.n37 163.367
R479 B.n320 B.n319 163.367
R480 B.n319 B.n318 163.367
R481 B.n318 B.n39 163.367
R482 B.n314 B.n39 163.367
R483 B.n314 B.n313 163.367
R484 B.n313 B.n312 163.367
R485 B.n312 B.n41 163.367
R486 B.n308 B.n41 163.367
R487 B.n308 B.n307 163.367
R488 B.n307 B.n306 163.367
R489 B.n306 B.n43 163.367
R490 B.n302 B.n43 163.367
R491 B.n302 B.n301 163.367
R492 B.n301 B.n300 163.367
R493 B.n300 B.n45 163.367
R494 B.n296 B.n45 163.367
R495 B.n80 B.t2 131.357
R496 B.n32 B.t7 131.357
R497 B.n88 B.t5 131.351
R498 B.n26 B.t10 131.351
R499 B.n81 B.t1 114.484
R500 B.n33 B.t8 114.484
R501 B.n89 B.t4 114.478
R502 B.n27 B.t11 114.478
R503 B.n82 B.n81 59.5399
R504 B.n179 B.n89 59.5399
R505 B.n348 B.n27 59.5399
R506 B.n334 B.n33 59.5399
R507 B.n385 B.n12 33.5615
R508 B.n297 B.n46 33.5615
R509 B.n232 B.n231 33.5615
R510 B.n142 B.n141 33.5615
R511 B B.n419 18.0485
R512 B.n81 B.n80 16.8732
R513 B.n89 B.n88 16.8732
R514 B.n27 B.n26 16.8732
R515 B.n33 B.n32 16.8732
R516 B.n385 B.n384 10.6151
R517 B.n384 B.n383 10.6151
R518 B.n383 B.n14 10.6151
R519 B.n379 B.n14 10.6151
R520 B.n379 B.n378 10.6151
R521 B.n378 B.n377 10.6151
R522 B.n377 B.n16 10.6151
R523 B.n373 B.n16 10.6151
R524 B.n373 B.n372 10.6151
R525 B.n372 B.n371 10.6151
R526 B.n371 B.n18 10.6151
R527 B.n367 B.n18 10.6151
R528 B.n367 B.n366 10.6151
R529 B.n366 B.n365 10.6151
R530 B.n365 B.n20 10.6151
R531 B.n361 B.n20 10.6151
R532 B.n361 B.n360 10.6151
R533 B.n360 B.n359 10.6151
R534 B.n359 B.n22 10.6151
R535 B.n355 B.n22 10.6151
R536 B.n355 B.n354 10.6151
R537 B.n354 B.n353 10.6151
R538 B.n353 B.n24 10.6151
R539 B.n349 B.n24 10.6151
R540 B.n347 B.n346 10.6151
R541 B.n346 B.n28 10.6151
R542 B.n342 B.n28 10.6151
R543 B.n342 B.n341 10.6151
R544 B.n341 B.n340 10.6151
R545 B.n340 B.n30 10.6151
R546 B.n336 B.n30 10.6151
R547 B.n336 B.n335 10.6151
R548 B.n333 B.n34 10.6151
R549 B.n329 B.n34 10.6151
R550 B.n329 B.n328 10.6151
R551 B.n328 B.n327 10.6151
R552 B.n327 B.n36 10.6151
R553 B.n323 B.n36 10.6151
R554 B.n323 B.n322 10.6151
R555 B.n322 B.n321 10.6151
R556 B.n321 B.n38 10.6151
R557 B.n317 B.n38 10.6151
R558 B.n317 B.n316 10.6151
R559 B.n316 B.n315 10.6151
R560 B.n315 B.n40 10.6151
R561 B.n311 B.n40 10.6151
R562 B.n311 B.n310 10.6151
R563 B.n310 B.n309 10.6151
R564 B.n309 B.n42 10.6151
R565 B.n305 B.n42 10.6151
R566 B.n305 B.n304 10.6151
R567 B.n304 B.n303 10.6151
R568 B.n303 B.n44 10.6151
R569 B.n299 B.n44 10.6151
R570 B.n299 B.n298 10.6151
R571 B.n298 B.n297 10.6151
R572 B.n233 B.n232 10.6151
R573 B.n233 B.n66 10.6151
R574 B.n237 B.n66 10.6151
R575 B.n238 B.n237 10.6151
R576 B.n239 B.n238 10.6151
R577 B.n239 B.n64 10.6151
R578 B.n243 B.n64 10.6151
R579 B.n244 B.n243 10.6151
R580 B.n245 B.n244 10.6151
R581 B.n245 B.n62 10.6151
R582 B.n249 B.n62 10.6151
R583 B.n250 B.n249 10.6151
R584 B.n251 B.n250 10.6151
R585 B.n251 B.n60 10.6151
R586 B.n255 B.n60 10.6151
R587 B.n256 B.n255 10.6151
R588 B.n257 B.n256 10.6151
R589 B.n257 B.n58 10.6151
R590 B.n261 B.n58 10.6151
R591 B.n262 B.n261 10.6151
R592 B.n263 B.n262 10.6151
R593 B.n263 B.n56 10.6151
R594 B.n267 B.n56 10.6151
R595 B.n268 B.n267 10.6151
R596 B.n269 B.n268 10.6151
R597 B.n269 B.n54 10.6151
R598 B.n273 B.n54 10.6151
R599 B.n274 B.n273 10.6151
R600 B.n275 B.n274 10.6151
R601 B.n275 B.n52 10.6151
R602 B.n279 B.n52 10.6151
R603 B.n280 B.n279 10.6151
R604 B.n281 B.n280 10.6151
R605 B.n281 B.n50 10.6151
R606 B.n285 B.n50 10.6151
R607 B.n286 B.n285 10.6151
R608 B.n287 B.n286 10.6151
R609 B.n287 B.n48 10.6151
R610 B.n291 B.n48 10.6151
R611 B.n292 B.n291 10.6151
R612 B.n293 B.n292 10.6151
R613 B.n293 B.n46 10.6151
R614 B.n143 B.n142 10.6151
R615 B.n143 B.n100 10.6151
R616 B.n147 B.n100 10.6151
R617 B.n148 B.n147 10.6151
R618 B.n149 B.n148 10.6151
R619 B.n149 B.n98 10.6151
R620 B.n153 B.n98 10.6151
R621 B.n154 B.n153 10.6151
R622 B.n155 B.n154 10.6151
R623 B.n155 B.n96 10.6151
R624 B.n159 B.n96 10.6151
R625 B.n160 B.n159 10.6151
R626 B.n161 B.n160 10.6151
R627 B.n161 B.n94 10.6151
R628 B.n165 B.n94 10.6151
R629 B.n166 B.n165 10.6151
R630 B.n167 B.n166 10.6151
R631 B.n167 B.n92 10.6151
R632 B.n171 B.n92 10.6151
R633 B.n172 B.n171 10.6151
R634 B.n173 B.n172 10.6151
R635 B.n173 B.n90 10.6151
R636 B.n177 B.n90 10.6151
R637 B.n178 B.n177 10.6151
R638 B.n180 B.n86 10.6151
R639 B.n184 B.n86 10.6151
R640 B.n185 B.n184 10.6151
R641 B.n186 B.n185 10.6151
R642 B.n186 B.n84 10.6151
R643 B.n190 B.n84 10.6151
R644 B.n191 B.n190 10.6151
R645 B.n192 B.n191 10.6151
R646 B.n196 B.n195 10.6151
R647 B.n197 B.n196 10.6151
R648 B.n197 B.n78 10.6151
R649 B.n201 B.n78 10.6151
R650 B.n202 B.n201 10.6151
R651 B.n203 B.n202 10.6151
R652 B.n203 B.n76 10.6151
R653 B.n207 B.n76 10.6151
R654 B.n208 B.n207 10.6151
R655 B.n209 B.n208 10.6151
R656 B.n209 B.n74 10.6151
R657 B.n213 B.n74 10.6151
R658 B.n214 B.n213 10.6151
R659 B.n215 B.n214 10.6151
R660 B.n215 B.n72 10.6151
R661 B.n219 B.n72 10.6151
R662 B.n220 B.n219 10.6151
R663 B.n221 B.n220 10.6151
R664 B.n221 B.n70 10.6151
R665 B.n225 B.n70 10.6151
R666 B.n226 B.n225 10.6151
R667 B.n227 B.n226 10.6151
R668 B.n227 B.n68 10.6151
R669 B.n231 B.n68 10.6151
R670 B.n141 B.n102 10.6151
R671 B.n137 B.n102 10.6151
R672 B.n137 B.n136 10.6151
R673 B.n136 B.n135 10.6151
R674 B.n135 B.n104 10.6151
R675 B.n131 B.n104 10.6151
R676 B.n131 B.n130 10.6151
R677 B.n130 B.n129 10.6151
R678 B.n129 B.n106 10.6151
R679 B.n125 B.n106 10.6151
R680 B.n125 B.n124 10.6151
R681 B.n124 B.n123 10.6151
R682 B.n123 B.n108 10.6151
R683 B.n119 B.n108 10.6151
R684 B.n119 B.n118 10.6151
R685 B.n118 B.n117 10.6151
R686 B.n117 B.n110 10.6151
R687 B.n113 B.n110 10.6151
R688 B.n113 B.n112 10.6151
R689 B.n112 B.n0 10.6151
R690 B.n415 B.n1 10.6151
R691 B.n415 B.n414 10.6151
R692 B.n414 B.n413 10.6151
R693 B.n413 B.n4 10.6151
R694 B.n409 B.n4 10.6151
R695 B.n409 B.n408 10.6151
R696 B.n408 B.n407 10.6151
R697 B.n407 B.n6 10.6151
R698 B.n403 B.n6 10.6151
R699 B.n403 B.n402 10.6151
R700 B.n402 B.n401 10.6151
R701 B.n401 B.n8 10.6151
R702 B.n397 B.n8 10.6151
R703 B.n397 B.n396 10.6151
R704 B.n396 B.n395 10.6151
R705 B.n395 B.n10 10.6151
R706 B.n391 B.n10 10.6151
R707 B.n391 B.n390 10.6151
R708 B.n390 B.n389 10.6151
R709 B.n389 B.n12 10.6151
R710 B.n348 B.n347 6.5566
R711 B.n335 B.n334 6.5566
R712 B.n180 B.n179 6.5566
R713 B.n192 B.n82 6.5566
R714 B.n349 B.n348 4.05904
R715 B.n334 B.n333 4.05904
R716 B.n179 B.n178 4.05904
R717 B.n195 B.n82 4.05904
R718 B.n419 B.n0 2.81026
R719 B.n419 B.n1 2.81026
R720 VN.n2 VN.t2 380.2
R721 VN.n10 VN.t1 380.2
R722 VN.n1 VN.t4 354.807
R723 VN.n4 VN.t5 354.807
R724 VN.n6 VN.t7 354.807
R725 VN.n9 VN.t0 354.807
R726 VN.n12 VN.t6 354.807
R727 VN.n14 VN.t3 354.807
R728 VN.n7 VN.n6 161.3
R729 VN.n15 VN.n14 161.3
R730 VN.n13 VN.n8 161.3
R731 VN.n12 VN.n11 161.3
R732 VN.n5 VN.n0 161.3
R733 VN.n4 VN.n3 161.3
R734 VN.n4 VN.n1 48.2005
R735 VN.n12 VN.n9 48.2005
R736 VN.n11 VN.n10 45.0031
R737 VN.n3 VN.n2 45.0031
R738 VN.n6 VN.n5 41.6278
R739 VN.n14 VN.n13 41.6278
R740 VN VN.n15 37.2903
R741 VN.n2 VN.n1 15.6319
R742 VN.n10 VN.n9 15.6319
R743 VN.n5 VN.n4 6.57323
R744 VN.n13 VN.n12 6.57323
R745 VN.n15 VN.n8 0.189894
R746 VN.n11 VN.n8 0.189894
R747 VN.n3 VN.n0 0.189894
R748 VN.n7 VN.n0 0.189894
R749 VN VN.n7 0.0516364
R750 VDD2.n2 VDD2.n1 89.7721
R751 VDD2.n2 VDD2.n0 89.7721
R752 VDD2 VDD2.n5 89.7693
R753 VDD2.n4 VDD2.n3 89.4527
R754 VDD2.n4 VDD2.n2 32.5386
R755 VDD2.n5 VDD2.t7 5.1437
R756 VDD2.n5 VDD2.t6 5.1437
R757 VDD2.n3 VDD2.t4 5.1437
R758 VDD2.n3 VDD2.t1 5.1437
R759 VDD2.n1 VDD2.t2 5.1437
R760 VDD2.n1 VDD2.t0 5.1437
R761 VDD2.n0 VDD2.t5 5.1437
R762 VDD2.n0 VDD2.t3 5.1437
R763 VDD2 VDD2.n4 0.43369
C0 VDD2 B 0.899927f
C1 w_n1840_n2232# VN 3.06558f
C2 VTAIL VP 2.67764f
C3 w_n1840_n2232# VDD1 1.08257f
C4 VDD1 VN 0.148197f
C5 VDD2 VP 0.300659f
C6 w_n1840_n2232# B 5.37348f
C7 VN B 0.677526f
C8 VDD2 VTAIL 7.54592f
C9 VDD1 B 0.868205f
C10 w_n1840_n2232# VP 3.29838f
C11 VN VP 4.09178f
C12 w_n1840_n2232# VTAIL 2.78188f
C13 VTAIL VN 2.66353f
C14 VDD1 VP 2.84869f
C15 VP B 1.05679f
C16 w_n1840_n2232# VDD2 1.11079f
C17 VDD2 VN 2.69658f
C18 VDD1 VTAIL 7.50532f
C19 VTAIL B 2.21599f
C20 VDD2 VDD1 0.746651f
C21 VDD2 VSUBS 1.115922f
C22 VDD1 VSUBS 1.39338f
C23 VTAIL VSUBS 0.496435f
C24 VN VSUBS 4.09491f
C25 VP VSUBS 1.202993f
C26 B VSUBS 2.221283f
C27 w_n1840_n2232# VSUBS 51.203503f
C28 VDD2.t5 VSUBS 0.140383f
C29 VDD2.t3 VSUBS 0.140383f
C30 VDD2.n0 VSUBS 0.943937f
C31 VDD2.t2 VSUBS 0.140383f
C32 VDD2.t0 VSUBS 0.140383f
C33 VDD2.n1 VSUBS 0.943937f
C34 VDD2.n2 VSUBS 2.42259f
C35 VDD2.t4 VSUBS 0.140383f
C36 VDD2.t1 VSUBS 0.140383f
C37 VDD2.n3 VSUBS 0.941891f
C38 VDD2.n4 VSUBS 2.24141f
C39 VDD2.t7 VSUBS 0.140383f
C40 VDD2.t6 VSUBS 0.140383f
C41 VDD2.n5 VSUBS 0.94391f
C42 VN.n0 VSUBS 0.06463f
C43 VN.t4 VSUBS 0.638681f
C44 VN.n1 VSUBS 0.307976f
C45 VN.t2 VSUBS 0.658371f
C46 VN.n2 VSUBS 0.279024f
C47 VN.n3 VSUBS 0.263219f
C48 VN.t5 VSUBS 0.638681f
C49 VN.n4 VSUBS 0.297166f
C50 VN.n5 VSUBS 0.014666f
C51 VN.t7 VSUBS 0.638681f
C52 VN.n6 VSUBS 0.293579f
C53 VN.n7 VSUBS 0.050086f
C54 VN.n8 VSUBS 0.06463f
C55 VN.t0 VSUBS 0.638681f
C56 VN.n9 VSUBS 0.307976f
C57 VN.t6 VSUBS 0.638681f
C58 VN.t1 VSUBS 0.658371f
C59 VN.n10 VSUBS 0.279024f
C60 VN.n11 VSUBS 0.263219f
C61 VN.n12 VSUBS 0.297166f
C62 VN.n13 VSUBS 0.014666f
C63 VN.t3 VSUBS 0.638681f
C64 VN.n14 VSUBS 0.293579f
C65 VN.n15 VSUBS 2.17113f
C66 B.n0 VSUBS 0.005838f
C67 B.n1 VSUBS 0.005838f
C68 B.n2 VSUBS 0.009233f
C69 B.n3 VSUBS 0.009233f
C70 B.n4 VSUBS 0.009233f
C71 B.n5 VSUBS 0.009233f
C72 B.n6 VSUBS 0.009233f
C73 B.n7 VSUBS 0.009233f
C74 B.n8 VSUBS 0.009233f
C75 B.n9 VSUBS 0.009233f
C76 B.n10 VSUBS 0.009233f
C77 B.n11 VSUBS 0.009233f
C78 B.n12 VSUBS 0.021749f
C79 B.n13 VSUBS 0.009233f
C80 B.n14 VSUBS 0.009233f
C81 B.n15 VSUBS 0.009233f
C82 B.n16 VSUBS 0.009233f
C83 B.n17 VSUBS 0.009233f
C84 B.n18 VSUBS 0.009233f
C85 B.n19 VSUBS 0.009233f
C86 B.n20 VSUBS 0.009233f
C87 B.n21 VSUBS 0.009233f
C88 B.n22 VSUBS 0.009233f
C89 B.n23 VSUBS 0.009233f
C90 B.n24 VSUBS 0.009233f
C91 B.n25 VSUBS 0.009233f
C92 B.t11 VSUBS 0.245957f
C93 B.t10 VSUBS 0.254852f
C94 B.t9 VSUBS 0.190301f
C95 B.n26 VSUBS 0.112795f
C96 B.n27 VSUBS 0.08241f
C97 B.n28 VSUBS 0.009233f
C98 B.n29 VSUBS 0.009233f
C99 B.n30 VSUBS 0.009233f
C100 B.n31 VSUBS 0.009233f
C101 B.t8 VSUBS 0.245957f
C102 B.t7 VSUBS 0.254851f
C103 B.t6 VSUBS 0.190301f
C104 B.n32 VSUBS 0.112796f
C105 B.n33 VSUBS 0.082411f
C106 B.n34 VSUBS 0.009233f
C107 B.n35 VSUBS 0.009233f
C108 B.n36 VSUBS 0.009233f
C109 B.n37 VSUBS 0.009233f
C110 B.n38 VSUBS 0.009233f
C111 B.n39 VSUBS 0.009233f
C112 B.n40 VSUBS 0.009233f
C113 B.n41 VSUBS 0.009233f
C114 B.n42 VSUBS 0.009233f
C115 B.n43 VSUBS 0.009233f
C116 B.n44 VSUBS 0.009233f
C117 B.n45 VSUBS 0.009233f
C118 B.n46 VSUBS 0.022811f
C119 B.n47 VSUBS 0.009233f
C120 B.n48 VSUBS 0.009233f
C121 B.n49 VSUBS 0.009233f
C122 B.n50 VSUBS 0.009233f
C123 B.n51 VSUBS 0.009233f
C124 B.n52 VSUBS 0.009233f
C125 B.n53 VSUBS 0.009233f
C126 B.n54 VSUBS 0.009233f
C127 B.n55 VSUBS 0.009233f
C128 B.n56 VSUBS 0.009233f
C129 B.n57 VSUBS 0.009233f
C130 B.n58 VSUBS 0.009233f
C131 B.n59 VSUBS 0.009233f
C132 B.n60 VSUBS 0.009233f
C133 B.n61 VSUBS 0.009233f
C134 B.n62 VSUBS 0.009233f
C135 B.n63 VSUBS 0.009233f
C136 B.n64 VSUBS 0.009233f
C137 B.n65 VSUBS 0.009233f
C138 B.n66 VSUBS 0.009233f
C139 B.n67 VSUBS 0.021749f
C140 B.n68 VSUBS 0.009233f
C141 B.n69 VSUBS 0.009233f
C142 B.n70 VSUBS 0.009233f
C143 B.n71 VSUBS 0.009233f
C144 B.n72 VSUBS 0.009233f
C145 B.n73 VSUBS 0.009233f
C146 B.n74 VSUBS 0.009233f
C147 B.n75 VSUBS 0.009233f
C148 B.n76 VSUBS 0.009233f
C149 B.n77 VSUBS 0.009233f
C150 B.n78 VSUBS 0.009233f
C151 B.n79 VSUBS 0.009233f
C152 B.t1 VSUBS 0.245957f
C153 B.t2 VSUBS 0.254851f
C154 B.t0 VSUBS 0.190301f
C155 B.n80 VSUBS 0.112796f
C156 B.n81 VSUBS 0.082411f
C157 B.n82 VSUBS 0.021391f
C158 B.n83 VSUBS 0.009233f
C159 B.n84 VSUBS 0.009233f
C160 B.n85 VSUBS 0.009233f
C161 B.n86 VSUBS 0.009233f
C162 B.n87 VSUBS 0.009233f
C163 B.t4 VSUBS 0.245957f
C164 B.t5 VSUBS 0.254852f
C165 B.t3 VSUBS 0.190301f
C166 B.n88 VSUBS 0.112795f
C167 B.n89 VSUBS 0.08241f
C168 B.n90 VSUBS 0.009233f
C169 B.n91 VSUBS 0.009233f
C170 B.n92 VSUBS 0.009233f
C171 B.n93 VSUBS 0.009233f
C172 B.n94 VSUBS 0.009233f
C173 B.n95 VSUBS 0.009233f
C174 B.n96 VSUBS 0.009233f
C175 B.n97 VSUBS 0.009233f
C176 B.n98 VSUBS 0.009233f
C177 B.n99 VSUBS 0.009233f
C178 B.n100 VSUBS 0.009233f
C179 B.n101 VSUBS 0.022241f
C180 B.n102 VSUBS 0.009233f
C181 B.n103 VSUBS 0.009233f
C182 B.n104 VSUBS 0.009233f
C183 B.n105 VSUBS 0.009233f
C184 B.n106 VSUBS 0.009233f
C185 B.n107 VSUBS 0.009233f
C186 B.n108 VSUBS 0.009233f
C187 B.n109 VSUBS 0.009233f
C188 B.n110 VSUBS 0.009233f
C189 B.n111 VSUBS 0.009233f
C190 B.n112 VSUBS 0.009233f
C191 B.n113 VSUBS 0.009233f
C192 B.n114 VSUBS 0.009233f
C193 B.n115 VSUBS 0.009233f
C194 B.n116 VSUBS 0.009233f
C195 B.n117 VSUBS 0.009233f
C196 B.n118 VSUBS 0.009233f
C197 B.n119 VSUBS 0.009233f
C198 B.n120 VSUBS 0.009233f
C199 B.n121 VSUBS 0.009233f
C200 B.n122 VSUBS 0.009233f
C201 B.n123 VSUBS 0.009233f
C202 B.n124 VSUBS 0.009233f
C203 B.n125 VSUBS 0.009233f
C204 B.n126 VSUBS 0.009233f
C205 B.n127 VSUBS 0.009233f
C206 B.n128 VSUBS 0.009233f
C207 B.n129 VSUBS 0.009233f
C208 B.n130 VSUBS 0.009233f
C209 B.n131 VSUBS 0.009233f
C210 B.n132 VSUBS 0.009233f
C211 B.n133 VSUBS 0.009233f
C212 B.n134 VSUBS 0.009233f
C213 B.n135 VSUBS 0.009233f
C214 B.n136 VSUBS 0.009233f
C215 B.n137 VSUBS 0.009233f
C216 B.n138 VSUBS 0.009233f
C217 B.n139 VSUBS 0.009233f
C218 B.n140 VSUBS 0.021749f
C219 B.n141 VSUBS 0.021749f
C220 B.n142 VSUBS 0.022241f
C221 B.n143 VSUBS 0.009233f
C222 B.n144 VSUBS 0.009233f
C223 B.n145 VSUBS 0.009233f
C224 B.n146 VSUBS 0.009233f
C225 B.n147 VSUBS 0.009233f
C226 B.n148 VSUBS 0.009233f
C227 B.n149 VSUBS 0.009233f
C228 B.n150 VSUBS 0.009233f
C229 B.n151 VSUBS 0.009233f
C230 B.n152 VSUBS 0.009233f
C231 B.n153 VSUBS 0.009233f
C232 B.n154 VSUBS 0.009233f
C233 B.n155 VSUBS 0.009233f
C234 B.n156 VSUBS 0.009233f
C235 B.n157 VSUBS 0.009233f
C236 B.n158 VSUBS 0.009233f
C237 B.n159 VSUBS 0.009233f
C238 B.n160 VSUBS 0.009233f
C239 B.n161 VSUBS 0.009233f
C240 B.n162 VSUBS 0.009233f
C241 B.n163 VSUBS 0.009233f
C242 B.n164 VSUBS 0.009233f
C243 B.n165 VSUBS 0.009233f
C244 B.n166 VSUBS 0.009233f
C245 B.n167 VSUBS 0.009233f
C246 B.n168 VSUBS 0.009233f
C247 B.n169 VSUBS 0.009233f
C248 B.n170 VSUBS 0.009233f
C249 B.n171 VSUBS 0.009233f
C250 B.n172 VSUBS 0.009233f
C251 B.n173 VSUBS 0.009233f
C252 B.n174 VSUBS 0.009233f
C253 B.n175 VSUBS 0.009233f
C254 B.n176 VSUBS 0.009233f
C255 B.n177 VSUBS 0.009233f
C256 B.n178 VSUBS 0.006381f
C257 B.n179 VSUBS 0.021391f
C258 B.n180 VSUBS 0.007468f
C259 B.n181 VSUBS 0.009233f
C260 B.n182 VSUBS 0.009233f
C261 B.n183 VSUBS 0.009233f
C262 B.n184 VSUBS 0.009233f
C263 B.n185 VSUBS 0.009233f
C264 B.n186 VSUBS 0.009233f
C265 B.n187 VSUBS 0.009233f
C266 B.n188 VSUBS 0.009233f
C267 B.n189 VSUBS 0.009233f
C268 B.n190 VSUBS 0.009233f
C269 B.n191 VSUBS 0.009233f
C270 B.n192 VSUBS 0.007468f
C271 B.n193 VSUBS 0.009233f
C272 B.n194 VSUBS 0.009233f
C273 B.n195 VSUBS 0.006381f
C274 B.n196 VSUBS 0.009233f
C275 B.n197 VSUBS 0.009233f
C276 B.n198 VSUBS 0.009233f
C277 B.n199 VSUBS 0.009233f
C278 B.n200 VSUBS 0.009233f
C279 B.n201 VSUBS 0.009233f
C280 B.n202 VSUBS 0.009233f
C281 B.n203 VSUBS 0.009233f
C282 B.n204 VSUBS 0.009233f
C283 B.n205 VSUBS 0.009233f
C284 B.n206 VSUBS 0.009233f
C285 B.n207 VSUBS 0.009233f
C286 B.n208 VSUBS 0.009233f
C287 B.n209 VSUBS 0.009233f
C288 B.n210 VSUBS 0.009233f
C289 B.n211 VSUBS 0.009233f
C290 B.n212 VSUBS 0.009233f
C291 B.n213 VSUBS 0.009233f
C292 B.n214 VSUBS 0.009233f
C293 B.n215 VSUBS 0.009233f
C294 B.n216 VSUBS 0.009233f
C295 B.n217 VSUBS 0.009233f
C296 B.n218 VSUBS 0.009233f
C297 B.n219 VSUBS 0.009233f
C298 B.n220 VSUBS 0.009233f
C299 B.n221 VSUBS 0.009233f
C300 B.n222 VSUBS 0.009233f
C301 B.n223 VSUBS 0.009233f
C302 B.n224 VSUBS 0.009233f
C303 B.n225 VSUBS 0.009233f
C304 B.n226 VSUBS 0.009233f
C305 B.n227 VSUBS 0.009233f
C306 B.n228 VSUBS 0.009233f
C307 B.n229 VSUBS 0.009233f
C308 B.n230 VSUBS 0.022241f
C309 B.n231 VSUBS 0.022241f
C310 B.n232 VSUBS 0.021749f
C311 B.n233 VSUBS 0.009233f
C312 B.n234 VSUBS 0.009233f
C313 B.n235 VSUBS 0.009233f
C314 B.n236 VSUBS 0.009233f
C315 B.n237 VSUBS 0.009233f
C316 B.n238 VSUBS 0.009233f
C317 B.n239 VSUBS 0.009233f
C318 B.n240 VSUBS 0.009233f
C319 B.n241 VSUBS 0.009233f
C320 B.n242 VSUBS 0.009233f
C321 B.n243 VSUBS 0.009233f
C322 B.n244 VSUBS 0.009233f
C323 B.n245 VSUBS 0.009233f
C324 B.n246 VSUBS 0.009233f
C325 B.n247 VSUBS 0.009233f
C326 B.n248 VSUBS 0.009233f
C327 B.n249 VSUBS 0.009233f
C328 B.n250 VSUBS 0.009233f
C329 B.n251 VSUBS 0.009233f
C330 B.n252 VSUBS 0.009233f
C331 B.n253 VSUBS 0.009233f
C332 B.n254 VSUBS 0.009233f
C333 B.n255 VSUBS 0.009233f
C334 B.n256 VSUBS 0.009233f
C335 B.n257 VSUBS 0.009233f
C336 B.n258 VSUBS 0.009233f
C337 B.n259 VSUBS 0.009233f
C338 B.n260 VSUBS 0.009233f
C339 B.n261 VSUBS 0.009233f
C340 B.n262 VSUBS 0.009233f
C341 B.n263 VSUBS 0.009233f
C342 B.n264 VSUBS 0.009233f
C343 B.n265 VSUBS 0.009233f
C344 B.n266 VSUBS 0.009233f
C345 B.n267 VSUBS 0.009233f
C346 B.n268 VSUBS 0.009233f
C347 B.n269 VSUBS 0.009233f
C348 B.n270 VSUBS 0.009233f
C349 B.n271 VSUBS 0.009233f
C350 B.n272 VSUBS 0.009233f
C351 B.n273 VSUBS 0.009233f
C352 B.n274 VSUBS 0.009233f
C353 B.n275 VSUBS 0.009233f
C354 B.n276 VSUBS 0.009233f
C355 B.n277 VSUBS 0.009233f
C356 B.n278 VSUBS 0.009233f
C357 B.n279 VSUBS 0.009233f
C358 B.n280 VSUBS 0.009233f
C359 B.n281 VSUBS 0.009233f
C360 B.n282 VSUBS 0.009233f
C361 B.n283 VSUBS 0.009233f
C362 B.n284 VSUBS 0.009233f
C363 B.n285 VSUBS 0.009233f
C364 B.n286 VSUBS 0.009233f
C365 B.n287 VSUBS 0.009233f
C366 B.n288 VSUBS 0.009233f
C367 B.n289 VSUBS 0.009233f
C368 B.n290 VSUBS 0.009233f
C369 B.n291 VSUBS 0.009233f
C370 B.n292 VSUBS 0.009233f
C371 B.n293 VSUBS 0.009233f
C372 B.n294 VSUBS 0.009233f
C373 B.n295 VSUBS 0.021749f
C374 B.n296 VSUBS 0.022241f
C375 B.n297 VSUBS 0.02118f
C376 B.n298 VSUBS 0.009233f
C377 B.n299 VSUBS 0.009233f
C378 B.n300 VSUBS 0.009233f
C379 B.n301 VSUBS 0.009233f
C380 B.n302 VSUBS 0.009233f
C381 B.n303 VSUBS 0.009233f
C382 B.n304 VSUBS 0.009233f
C383 B.n305 VSUBS 0.009233f
C384 B.n306 VSUBS 0.009233f
C385 B.n307 VSUBS 0.009233f
C386 B.n308 VSUBS 0.009233f
C387 B.n309 VSUBS 0.009233f
C388 B.n310 VSUBS 0.009233f
C389 B.n311 VSUBS 0.009233f
C390 B.n312 VSUBS 0.009233f
C391 B.n313 VSUBS 0.009233f
C392 B.n314 VSUBS 0.009233f
C393 B.n315 VSUBS 0.009233f
C394 B.n316 VSUBS 0.009233f
C395 B.n317 VSUBS 0.009233f
C396 B.n318 VSUBS 0.009233f
C397 B.n319 VSUBS 0.009233f
C398 B.n320 VSUBS 0.009233f
C399 B.n321 VSUBS 0.009233f
C400 B.n322 VSUBS 0.009233f
C401 B.n323 VSUBS 0.009233f
C402 B.n324 VSUBS 0.009233f
C403 B.n325 VSUBS 0.009233f
C404 B.n326 VSUBS 0.009233f
C405 B.n327 VSUBS 0.009233f
C406 B.n328 VSUBS 0.009233f
C407 B.n329 VSUBS 0.009233f
C408 B.n330 VSUBS 0.009233f
C409 B.n331 VSUBS 0.009233f
C410 B.n332 VSUBS 0.009233f
C411 B.n333 VSUBS 0.006381f
C412 B.n334 VSUBS 0.021391f
C413 B.n335 VSUBS 0.007468f
C414 B.n336 VSUBS 0.009233f
C415 B.n337 VSUBS 0.009233f
C416 B.n338 VSUBS 0.009233f
C417 B.n339 VSUBS 0.009233f
C418 B.n340 VSUBS 0.009233f
C419 B.n341 VSUBS 0.009233f
C420 B.n342 VSUBS 0.009233f
C421 B.n343 VSUBS 0.009233f
C422 B.n344 VSUBS 0.009233f
C423 B.n345 VSUBS 0.009233f
C424 B.n346 VSUBS 0.009233f
C425 B.n347 VSUBS 0.007468f
C426 B.n348 VSUBS 0.021391f
C427 B.n349 VSUBS 0.006381f
C428 B.n350 VSUBS 0.009233f
C429 B.n351 VSUBS 0.009233f
C430 B.n352 VSUBS 0.009233f
C431 B.n353 VSUBS 0.009233f
C432 B.n354 VSUBS 0.009233f
C433 B.n355 VSUBS 0.009233f
C434 B.n356 VSUBS 0.009233f
C435 B.n357 VSUBS 0.009233f
C436 B.n358 VSUBS 0.009233f
C437 B.n359 VSUBS 0.009233f
C438 B.n360 VSUBS 0.009233f
C439 B.n361 VSUBS 0.009233f
C440 B.n362 VSUBS 0.009233f
C441 B.n363 VSUBS 0.009233f
C442 B.n364 VSUBS 0.009233f
C443 B.n365 VSUBS 0.009233f
C444 B.n366 VSUBS 0.009233f
C445 B.n367 VSUBS 0.009233f
C446 B.n368 VSUBS 0.009233f
C447 B.n369 VSUBS 0.009233f
C448 B.n370 VSUBS 0.009233f
C449 B.n371 VSUBS 0.009233f
C450 B.n372 VSUBS 0.009233f
C451 B.n373 VSUBS 0.009233f
C452 B.n374 VSUBS 0.009233f
C453 B.n375 VSUBS 0.009233f
C454 B.n376 VSUBS 0.009233f
C455 B.n377 VSUBS 0.009233f
C456 B.n378 VSUBS 0.009233f
C457 B.n379 VSUBS 0.009233f
C458 B.n380 VSUBS 0.009233f
C459 B.n381 VSUBS 0.009233f
C460 B.n382 VSUBS 0.009233f
C461 B.n383 VSUBS 0.009233f
C462 B.n384 VSUBS 0.009233f
C463 B.n385 VSUBS 0.022241f
C464 B.n386 VSUBS 0.022241f
C465 B.n387 VSUBS 0.021749f
C466 B.n388 VSUBS 0.009233f
C467 B.n389 VSUBS 0.009233f
C468 B.n390 VSUBS 0.009233f
C469 B.n391 VSUBS 0.009233f
C470 B.n392 VSUBS 0.009233f
C471 B.n393 VSUBS 0.009233f
C472 B.n394 VSUBS 0.009233f
C473 B.n395 VSUBS 0.009233f
C474 B.n396 VSUBS 0.009233f
C475 B.n397 VSUBS 0.009233f
C476 B.n398 VSUBS 0.009233f
C477 B.n399 VSUBS 0.009233f
C478 B.n400 VSUBS 0.009233f
C479 B.n401 VSUBS 0.009233f
C480 B.n402 VSUBS 0.009233f
C481 B.n403 VSUBS 0.009233f
C482 B.n404 VSUBS 0.009233f
C483 B.n405 VSUBS 0.009233f
C484 B.n406 VSUBS 0.009233f
C485 B.n407 VSUBS 0.009233f
C486 B.n408 VSUBS 0.009233f
C487 B.n409 VSUBS 0.009233f
C488 B.n410 VSUBS 0.009233f
C489 B.n411 VSUBS 0.009233f
C490 B.n412 VSUBS 0.009233f
C491 B.n413 VSUBS 0.009233f
C492 B.n414 VSUBS 0.009233f
C493 B.n415 VSUBS 0.009233f
C494 B.n416 VSUBS 0.009233f
C495 B.n417 VSUBS 0.009233f
C496 B.n418 VSUBS 0.009233f
C497 B.n419 VSUBS 0.020906f
C498 VDD1.t3 VSUBS 0.140331f
C499 VDD1.t5 VSUBS 0.140331f
C500 VDD1.n0 VSUBS 0.944355f
C501 VDD1.t4 VSUBS 0.140331f
C502 VDD1.t7 VSUBS 0.140331f
C503 VDD1.n1 VSUBS 0.943587f
C504 VDD1.t6 VSUBS 0.140331f
C505 VDD1.t1 VSUBS 0.140331f
C506 VDD1.n2 VSUBS 0.943587f
C507 VDD1.n3 VSUBS 2.48206f
C508 VDD1.t0 VSUBS 0.140331f
C509 VDD1.t2 VSUBS 0.140331f
C510 VDD1.n4 VSUBS 0.941537f
C511 VDD1.n5 VSUBS 2.27346f
C512 VTAIL.t1 VSUBS 0.139042f
C513 VTAIL.t0 VSUBS 0.139042f
C514 VTAIL.n0 VSUBS 0.828457f
C515 VTAIL.n1 VSUBS 0.600051f
C516 VTAIL.t5 VSUBS 1.13712f
C517 VTAIL.n2 VSUBS 0.707518f
C518 VTAIL.t14 VSUBS 1.13712f
C519 VTAIL.n3 VSUBS 0.707518f
C520 VTAIL.t8 VSUBS 0.139042f
C521 VTAIL.t13 VSUBS 0.139042f
C522 VTAIL.n4 VSUBS 0.828457f
C523 VTAIL.n5 VSUBS 0.662112f
C524 VTAIL.t11 VSUBS 1.13712f
C525 VTAIL.n6 VSUBS 1.59958f
C526 VTAIL.t2 VSUBS 1.13713f
C527 VTAIL.n7 VSUBS 1.59958f
C528 VTAIL.t7 VSUBS 0.139042f
C529 VTAIL.t3 VSUBS 0.139042f
C530 VTAIL.n8 VSUBS 0.828462f
C531 VTAIL.n9 VSUBS 0.662107f
C532 VTAIL.t4 VSUBS 1.13713f
C533 VTAIL.n10 VSUBS 0.707511f
C534 VTAIL.t15 VSUBS 1.13713f
C535 VTAIL.n11 VSUBS 0.707511f
C536 VTAIL.t12 VSUBS 0.139042f
C537 VTAIL.t9 VSUBS 0.139042f
C538 VTAIL.n12 VSUBS 0.828462f
C539 VTAIL.n13 VSUBS 0.662107f
C540 VTAIL.t10 VSUBS 1.13712f
C541 VTAIL.n14 VSUBS 1.59958f
C542 VTAIL.t6 VSUBS 1.13712f
C543 VTAIL.n15 VSUBS 1.59436f
C544 VP.n0 VSUBS 0.06665f
C545 VP.t0 VSUBS 0.658636f
C546 VP.n1 VSUBS 0.306451f
C547 VP.n2 VSUBS 0.06665f
C548 VP.t5 VSUBS 0.658636f
C549 VP.t7 VSUBS 0.658636f
C550 VP.n3 VSUBS 0.271443f
C551 VP.t2 VSUBS 0.658636f
C552 VP.t4 VSUBS 0.678942f
C553 VP.n4 VSUBS 0.287742f
C554 VP.n5 VSUBS 0.317598f
C555 VP.n6 VSUBS 0.306451f
C556 VP.n7 VSUBS 0.015124f
C557 VP.n8 VSUBS 0.302752f
C558 VP.n9 VSUBS 2.19484f
C559 VP.n10 VSUBS 2.25994f
C560 VP.t3 VSUBS 0.658636f
C561 VP.n11 VSUBS 0.302752f
C562 VP.n12 VSUBS 0.015124f
C563 VP.n13 VSUBS 0.06665f
C564 VP.n14 VSUBS 0.06665f
C565 VP.n15 VSUBS 0.06665f
C566 VP.t1 VSUBS 0.658636f
C567 VP.n16 VSUBS 0.306451f
C568 VP.n17 VSUBS 0.015124f
C569 VP.t6 VSUBS 0.658636f
C570 VP.n18 VSUBS 0.302752f
C571 VP.n19 VSUBS 0.051651f
.ends

