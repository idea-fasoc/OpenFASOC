* NGSPICE file created from diff_pair_sample_0987.ext - technology: sky130A

.subckt diff_pair_sample_0987 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0 ps=0 w=0.66 l=3.2
X1 VTAIL.t7 VP.t0 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0.1089 ps=0.99 w=0.66 l=3.2
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0 ps=0 w=0.66 l=3.2
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0 ps=0 w=0.66 l=3.2
X4 VDD1.t3 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1089 pd=0.99 as=0.2574 ps=2.1 w=0.66 l=3.2
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0 ps=0 w=0.66 l=3.2
X6 VDD1.t2 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1089 pd=0.99 as=0.2574 ps=2.1 w=0.66 l=3.2
X7 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0.1089 ps=0.99 w=0.66 l=3.2
X8 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1089 pd=0.99 as=0.2574 ps=2.1 w=0.66 l=3.2
X9 VTAIL.t4 VP.t3 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0.1089 ps=0.99 w=0.66 l=3.2
X10 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1089 pd=0.99 as=0.2574 ps=2.1 w=0.66 l=3.2
X11 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2574 pd=2.1 as=0.1089 ps=0.99 w=0.66 l=3.2
R0 B.n452 B.n451 585
R1 B.n138 B.n86 585
R2 B.n137 B.n136 585
R3 B.n135 B.n134 585
R4 B.n133 B.n132 585
R5 B.n131 B.n130 585
R6 B.n129 B.n128 585
R7 B.n127 B.n126 585
R8 B.n125 B.n124 585
R9 B.n123 B.n122 585
R10 B.n121 B.n120 585
R11 B.n119 B.n118 585
R12 B.n117 B.n116 585
R13 B.n115 B.n114 585
R14 B.n113 B.n112 585
R15 B.n111 B.n110 585
R16 B.n109 B.n108 585
R17 B.n107 B.n106 585
R18 B.n105 B.n104 585
R19 B.n103 B.n102 585
R20 B.n101 B.n100 585
R21 B.n99 B.n98 585
R22 B.n97 B.n96 585
R23 B.n95 B.n94 585
R24 B.n74 B.n73 585
R25 B.n457 B.n456 585
R26 B.n450 B.n87 585
R27 B.n87 B.n71 585
R28 B.n449 B.n70 585
R29 B.n461 B.n70 585
R30 B.n448 B.n69 585
R31 B.n462 B.n69 585
R32 B.n447 B.n68 585
R33 B.n463 B.n68 585
R34 B.n446 B.n445 585
R35 B.n445 B.n64 585
R36 B.n444 B.n63 585
R37 B.n469 B.n63 585
R38 B.n443 B.n62 585
R39 B.n470 B.n62 585
R40 B.n442 B.n61 585
R41 B.n471 B.n61 585
R42 B.n441 B.n440 585
R43 B.n440 B.n60 585
R44 B.n439 B.n56 585
R45 B.n477 B.n56 585
R46 B.n438 B.n55 585
R47 B.n478 B.n55 585
R48 B.n437 B.n54 585
R49 B.n479 B.n54 585
R50 B.n436 B.n435 585
R51 B.n435 B.n50 585
R52 B.n434 B.n49 585
R53 B.n485 B.n49 585
R54 B.n433 B.n48 585
R55 B.n486 B.n48 585
R56 B.n432 B.n47 585
R57 B.n487 B.n47 585
R58 B.n431 B.n430 585
R59 B.n430 B.n43 585
R60 B.n429 B.n42 585
R61 B.n493 B.n42 585
R62 B.n428 B.n41 585
R63 B.n494 B.n41 585
R64 B.n427 B.n40 585
R65 B.n495 B.n40 585
R66 B.n426 B.n425 585
R67 B.n425 B.n36 585
R68 B.n424 B.n35 585
R69 B.n501 B.n35 585
R70 B.n423 B.n34 585
R71 B.n502 B.n34 585
R72 B.n422 B.n33 585
R73 B.n503 B.n33 585
R74 B.n421 B.n420 585
R75 B.n420 B.n29 585
R76 B.n419 B.n28 585
R77 B.n509 B.n28 585
R78 B.n418 B.n27 585
R79 B.n510 B.n27 585
R80 B.n417 B.n26 585
R81 B.n511 B.n26 585
R82 B.n416 B.n415 585
R83 B.n415 B.n22 585
R84 B.n414 B.n21 585
R85 B.n517 B.n21 585
R86 B.n413 B.n20 585
R87 B.n518 B.n20 585
R88 B.n412 B.n19 585
R89 B.n519 B.n19 585
R90 B.n411 B.n410 585
R91 B.n410 B.n18 585
R92 B.n409 B.n14 585
R93 B.n525 B.n14 585
R94 B.n408 B.n13 585
R95 B.n526 B.n13 585
R96 B.n407 B.n12 585
R97 B.n527 B.n12 585
R98 B.n406 B.n405 585
R99 B.n405 B.n8 585
R100 B.n404 B.n7 585
R101 B.n533 B.n7 585
R102 B.n403 B.n6 585
R103 B.n534 B.n6 585
R104 B.n402 B.n5 585
R105 B.n535 B.n5 585
R106 B.n401 B.n400 585
R107 B.n400 B.n4 585
R108 B.n399 B.n139 585
R109 B.n399 B.n398 585
R110 B.n389 B.n140 585
R111 B.n141 B.n140 585
R112 B.n391 B.n390 585
R113 B.n392 B.n391 585
R114 B.n388 B.n146 585
R115 B.n146 B.n145 585
R116 B.n387 B.n386 585
R117 B.n386 B.n385 585
R118 B.n148 B.n147 585
R119 B.n378 B.n148 585
R120 B.n377 B.n376 585
R121 B.n379 B.n377 585
R122 B.n375 B.n153 585
R123 B.n153 B.n152 585
R124 B.n374 B.n373 585
R125 B.n373 B.n372 585
R126 B.n155 B.n154 585
R127 B.n156 B.n155 585
R128 B.n365 B.n364 585
R129 B.n366 B.n365 585
R130 B.n363 B.n161 585
R131 B.n161 B.n160 585
R132 B.n362 B.n361 585
R133 B.n361 B.n360 585
R134 B.n163 B.n162 585
R135 B.n164 B.n163 585
R136 B.n353 B.n352 585
R137 B.n354 B.n353 585
R138 B.n351 B.n169 585
R139 B.n169 B.n168 585
R140 B.n350 B.n349 585
R141 B.n349 B.n348 585
R142 B.n171 B.n170 585
R143 B.n172 B.n171 585
R144 B.n341 B.n340 585
R145 B.n342 B.n341 585
R146 B.n339 B.n177 585
R147 B.n177 B.n176 585
R148 B.n338 B.n337 585
R149 B.n337 B.n336 585
R150 B.n179 B.n178 585
R151 B.n180 B.n179 585
R152 B.n329 B.n328 585
R153 B.n330 B.n329 585
R154 B.n327 B.n185 585
R155 B.n185 B.n184 585
R156 B.n326 B.n325 585
R157 B.n325 B.n324 585
R158 B.n187 B.n186 585
R159 B.n188 B.n187 585
R160 B.n317 B.n316 585
R161 B.n318 B.n317 585
R162 B.n315 B.n193 585
R163 B.n193 B.n192 585
R164 B.n314 B.n313 585
R165 B.n313 B.n312 585
R166 B.n195 B.n194 585
R167 B.n305 B.n195 585
R168 B.n304 B.n303 585
R169 B.n306 B.n304 585
R170 B.n302 B.n200 585
R171 B.n200 B.n199 585
R172 B.n301 B.n300 585
R173 B.n300 B.n299 585
R174 B.n202 B.n201 585
R175 B.n203 B.n202 585
R176 B.n292 B.n291 585
R177 B.n293 B.n292 585
R178 B.n290 B.n208 585
R179 B.n208 B.n207 585
R180 B.n289 B.n288 585
R181 B.n288 B.n287 585
R182 B.n210 B.n209 585
R183 B.n211 B.n210 585
R184 B.n283 B.n282 585
R185 B.n214 B.n213 585
R186 B.n279 B.n278 585
R187 B.n280 B.n279 585
R188 B.n277 B.n227 585
R189 B.n276 B.n275 585
R190 B.n274 B.n273 585
R191 B.n272 B.n271 585
R192 B.n270 B.n269 585
R193 B.n267 B.n266 585
R194 B.n265 B.n264 585
R195 B.n263 B.n262 585
R196 B.n261 B.n260 585
R197 B.n259 B.n258 585
R198 B.n257 B.n256 585
R199 B.n255 B.n254 585
R200 B.n253 B.n252 585
R201 B.n251 B.n250 585
R202 B.n249 B.n248 585
R203 B.n246 B.n245 585
R204 B.n244 B.n243 585
R205 B.n242 B.n241 585
R206 B.n240 B.n239 585
R207 B.n238 B.n237 585
R208 B.n236 B.n235 585
R209 B.n234 B.n233 585
R210 B.n232 B.n226 585
R211 B.n280 B.n226 585
R212 B.n284 B.n212 585
R213 B.n212 B.n211 585
R214 B.n286 B.n285 585
R215 B.n287 B.n286 585
R216 B.n206 B.n205 585
R217 B.n207 B.n206 585
R218 B.n295 B.n294 585
R219 B.n294 B.n293 585
R220 B.n296 B.n204 585
R221 B.n204 B.n203 585
R222 B.n298 B.n297 585
R223 B.n299 B.n298 585
R224 B.n198 B.n197 585
R225 B.n199 B.n198 585
R226 B.n308 B.n307 585
R227 B.n307 B.n306 585
R228 B.n309 B.n196 585
R229 B.n305 B.n196 585
R230 B.n311 B.n310 585
R231 B.n312 B.n311 585
R232 B.n191 B.n190 585
R233 B.n192 B.n191 585
R234 B.n320 B.n319 585
R235 B.n319 B.n318 585
R236 B.n321 B.n189 585
R237 B.n189 B.n188 585
R238 B.n323 B.n322 585
R239 B.n324 B.n323 585
R240 B.n183 B.n182 585
R241 B.n184 B.n183 585
R242 B.n332 B.n331 585
R243 B.n331 B.n330 585
R244 B.n333 B.n181 585
R245 B.n181 B.n180 585
R246 B.n335 B.n334 585
R247 B.n336 B.n335 585
R248 B.n175 B.n174 585
R249 B.n176 B.n175 585
R250 B.n344 B.n343 585
R251 B.n343 B.n342 585
R252 B.n345 B.n173 585
R253 B.n173 B.n172 585
R254 B.n347 B.n346 585
R255 B.n348 B.n347 585
R256 B.n167 B.n166 585
R257 B.n168 B.n167 585
R258 B.n356 B.n355 585
R259 B.n355 B.n354 585
R260 B.n357 B.n165 585
R261 B.n165 B.n164 585
R262 B.n359 B.n358 585
R263 B.n360 B.n359 585
R264 B.n159 B.n158 585
R265 B.n160 B.n159 585
R266 B.n368 B.n367 585
R267 B.n367 B.n366 585
R268 B.n369 B.n157 585
R269 B.n157 B.n156 585
R270 B.n371 B.n370 585
R271 B.n372 B.n371 585
R272 B.n151 B.n150 585
R273 B.n152 B.n151 585
R274 B.n381 B.n380 585
R275 B.n380 B.n379 585
R276 B.n382 B.n149 585
R277 B.n378 B.n149 585
R278 B.n384 B.n383 585
R279 B.n385 B.n384 585
R280 B.n144 B.n143 585
R281 B.n145 B.n144 585
R282 B.n394 B.n393 585
R283 B.n393 B.n392 585
R284 B.n395 B.n142 585
R285 B.n142 B.n141 585
R286 B.n397 B.n396 585
R287 B.n398 B.n397 585
R288 B.n2 B.n0 585
R289 B.n4 B.n2 585
R290 B.n3 B.n1 585
R291 B.n534 B.n3 585
R292 B.n532 B.n531 585
R293 B.n533 B.n532 585
R294 B.n530 B.n9 585
R295 B.n9 B.n8 585
R296 B.n529 B.n528 585
R297 B.n528 B.n527 585
R298 B.n11 B.n10 585
R299 B.n526 B.n11 585
R300 B.n524 B.n523 585
R301 B.n525 B.n524 585
R302 B.n522 B.n15 585
R303 B.n18 B.n15 585
R304 B.n521 B.n520 585
R305 B.n520 B.n519 585
R306 B.n17 B.n16 585
R307 B.n518 B.n17 585
R308 B.n516 B.n515 585
R309 B.n517 B.n516 585
R310 B.n514 B.n23 585
R311 B.n23 B.n22 585
R312 B.n513 B.n512 585
R313 B.n512 B.n511 585
R314 B.n25 B.n24 585
R315 B.n510 B.n25 585
R316 B.n508 B.n507 585
R317 B.n509 B.n508 585
R318 B.n506 B.n30 585
R319 B.n30 B.n29 585
R320 B.n505 B.n504 585
R321 B.n504 B.n503 585
R322 B.n32 B.n31 585
R323 B.n502 B.n32 585
R324 B.n500 B.n499 585
R325 B.n501 B.n500 585
R326 B.n498 B.n37 585
R327 B.n37 B.n36 585
R328 B.n497 B.n496 585
R329 B.n496 B.n495 585
R330 B.n39 B.n38 585
R331 B.n494 B.n39 585
R332 B.n492 B.n491 585
R333 B.n493 B.n492 585
R334 B.n490 B.n44 585
R335 B.n44 B.n43 585
R336 B.n489 B.n488 585
R337 B.n488 B.n487 585
R338 B.n46 B.n45 585
R339 B.n486 B.n46 585
R340 B.n484 B.n483 585
R341 B.n485 B.n484 585
R342 B.n482 B.n51 585
R343 B.n51 B.n50 585
R344 B.n481 B.n480 585
R345 B.n480 B.n479 585
R346 B.n53 B.n52 585
R347 B.n478 B.n53 585
R348 B.n476 B.n475 585
R349 B.n477 B.n476 585
R350 B.n474 B.n57 585
R351 B.n60 B.n57 585
R352 B.n473 B.n472 585
R353 B.n472 B.n471 585
R354 B.n59 B.n58 585
R355 B.n470 B.n59 585
R356 B.n468 B.n467 585
R357 B.n469 B.n468 585
R358 B.n466 B.n65 585
R359 B.n65 B.n64 585
R360 B.n465 B.n464 585
R361 B.n464 B.n463 585
R362 B.n67 B.n66 585
R363 B.n462 B.n67 585
R364 B.n460 B.n459 585
R365 B.n461 B.n460 585
R366 B.n458 B.n72 585
R367 B.n72 B.n71 585
R368 B.n537 B.n536 585
R369 B.n536 B.n535 585
R370 B.n282 B.n212 550.159
R371 B.n456 B.n72 550.159
R372 B.n226 B.n210 550.159
R373 B.n452 B.n87 550.159
R374 B.n230 B.t7 306.151
R375 B.n228 B.t14 306.151
R376 B.n91 B.t16 306.151
R377 B.n88 B.t10 306.151
R378 B.n280 B.n211 261.332
R379 B.n454 B.n71 261.332
R380 B.n454 B.n453 256.663
R381 B.n454 B.n85 256.663
R382 B.n454 B.n84 256.663
R383 B.n454 B.n83 256.663
R384 B.n454 B.n82 256.663
R385 B.n454 B.n81 256.663
R386 B.n454 B.n80 256.663
R387 B.n454 B.n79 256.663
R388 B.n454 B.n78 256.663
R389 B.n454 B.n77 256.663
R390 B.n454 B.n76 256.663
R391 B.n454 B.n75 256.663
R392 B.n455 B.n454 256.663
R393 B.n281 B.n280 256.663
R394 B.n280 B.n215 256.663
R395 B.n280 B.n216 256.663
R396 B.n280 B.n217 256.663
R397 B.n280 B.n218 256.663
R398 B.n280 B.n219 256.663
R399 B.n280 B.n220 256.663
R400 B.n280 B.n221 256.663
R401 B.n280 B.n222 256.663
R402 B.n280 B.n223 256.663
R403 B.n280 B.n224 256.663
R404 B.n280 B.n225 256.663
R405 B.n231 B.t6 237.691
R406 B.n229 B.t13 237.691
R407 B.n92 B.t17 237.691
R408 B.n89 B.t11 237.691
R409 B.n230 B.t4 210.529
R410 B.n88 B.t8 210.529
R411 B.n228 B.t12 210.316
R412 B.n91 B.t15 210.316
R413 B.n286 B.n212 163.367
R414 B.n286 B.n206 163.367
R415 B.n294 B.n206 163.367
R416 B.n294 B.n204 163.367
R417 B.n298 B.n204 163.367
R418 B.n298 B.n198 163.367
R419 B.n307 B.n198 163.367
R420 B.n307 B.n196 163.367
R421 B.n311 B.n196 163.367
R422 B.n311 B.n191 163.367
R423 B.n319 B.n191 163.367
R424 B.n319 B.n189 163.367
R425 B.n323 B.n189 163.367
R426 B.n323 B.n183 163.367
R427 B.n331 B.n183 163.367
R428 B.n331 B.n181 163.367
R429 B.n335 B.n181 163.367
R430 B.n335 B.n175 163.367
R431 B.n343 B.n175 163.367
R432 B.n343 B.n173 163.367
R433 B.n347 B.n173 163.367
R434 B.n347 B.n167 163.367
R435 B.n355 B.n167 163.367
R436 B.n355 B.n165 163.367
R437 B.n359 B.n165 163.367
R438 B.n359 B.n159 163.367
R439 B.n367 B.n159 163.367
R440 B.n367 B.n157 163.367
R441 B.n371 B.n157 163.367
R442 B.n371 B.n151 163.367
R443 B.n380 B.n151 163.367
R444 B.n380 B.n149 163.367
R445 B.n384 B.n149 163.367
R446 B.n384 B.n144 163.367
R447 B.n393 B.n144 163.367
R448 B.n393 B.n142 163.367
R449 B.n397 B.n142 163.367
R450 B.n397 B.n2 163.367
R451 B.n536 B.n2 163.367
R452 B.n536 B.n3 163.367
R453 B.n532 B.n3 163.367
R454 B.n532 B.n9 163.367
R455 B.n528 B.n9 163.367
R456 B.n528 B.n11 163.367
R457 B.n524 B.n11 163.367
R458 B.n524 B.n15 163.367
R459 B.n520 B.n15 163.367
R460 B.n520 B.n17 163.367
R461 B.n516 B.n17 163.367
R462 B.n516 B.n23 163.367
R463 B.n512 B.n23 163.367
R464 B.n512 B.n25 163.367
R465 B.n508 B.n25 163.367
R466 B.n508 B.n30 163.367
R467 B.n504 B.n30 163.367
R468 B.n504 B.n32 163.367
R469 B.n500 B.n32 163.367
R470 B.n500 B.n37 163.367
R471 B.n496 B.n37 163.367
R472 B.n496 B.n39 163.367
R473 B.n492 B.n39 163.367
R474 B.n492 B.n44 163.367
R475 B.n488 B.n44 163.367
R476 B.n488 B.n46 163.367
R477 B.n484 B.n46 163.367
R478 B.n484 B.n51 163.367
R479 B.n480 B.n51 163.367
R480 B.n480 B.n53 163.367
R481 B.n476 B.n53 163.367
R482 B.n476 B.n57 163.367
R483 B.n472 B.n57 163.367
R484 B.n472 B.n59 163.367
R485 B.n468 B.n59 163.367
R486 B.n468 B.n65 163.367
R487 B.n464 B.n65 163.367
R488 B.n464 B.n67 163.367
R489 B.n460 B.n67 163.367
R490 B.n460 B.n72 163.367
R491 B.n279 B.n214 163.367
R492 B.n279 B.n227 163.367
R493 B.n275 B.n274 163.367
R494 B.n271 B.n270 163.367
R495 B.n266 B.n265 163.367
R496 B.n262 B.n261 163.367
R497 B.n258 B.n257 163.367
R498 B.n254 B.n253 163.367
R499 B.n250 B.n249 163.367
R500 B.n245 B.n244 163.367
R501 B.n241 B.n240 163.367
R502 B.n237 B.n236 163.367
R503 B.n233 B.n226 163.367
R504 B.n288 B.n210 163.367
R505 B.n288 B.n208 163.367
R506 B.n292 B.n208 163.367
R507 B.n292 B.n202 163.367
R508 B.n300 B.n202 163.367
R509 B.n300 B.n200 163.367
R510 B.n304 B.n200 163.367
R511 B.n304 B.n195 163.367
R512 B.n313 B.n195 163.367
R513 B.n313 B.n193 163.367
R514 B.n317 B.n193 163.367
R515 B.n317 B.n187 163.367
R516 B.n325 B.n187 163.367
R517 B.n325 B.n185 163.367
R518 B.n329 B.n185 163.367
R519 B.n329 B.n179 163.367
R520 B.n337 B.n179 163.367
R521 B.n337 B.n177 163.367
R522 B.n341 B.n177 163.367
R523 B.n341 B.n171 163.367
R524 B.n349 B.n171 163.367
R525 B.n349 B.n169 163.367
R526 B.n353 B.n169 163.367
R527 B.n353 B.n163 163.367
R528 B.n361 B.n163 163.367
R529 B.n361 B.n161 163.367
R530 B.n365 B.n161 163.367
R531 B.n365 B.n155 163.367
R532 B.n373 B.n155 163.367
R533 B.n373 B.n153 163.367
R534 B.n377 B.n153 163.367
R535 B.n377 B.n148 163.367
R536 B.n386 B.n148 163.367
R537 B.n386 B.n146 163.367
R538 B.n391 B.n146 163.367
R539 B.n391 B.n140 163.367
R540 B.n399 B.n140 163.367
R541 B.n400 B.n399 163.367
R542 B.n400 B.n5 163.367
R543 B.n6 B.n5 163.367
R544 B.n7 B.n6 163.367
R545 B.n405 B.n7 163.367
R546 B.n405 B.n12 163.367
R547 B.n13 B.n12 163.367
R548 B.n14 B.n13 163.367
R549 B.n410 B.n14 163.367
R550 B.n410 B.n19 163.367
R551 B.n20 B.n19 163.367
R552 B.n21 B.n20 163.367
R553 B.n415 B.n21 163.367
R554 B.n415 B.n26 163.367
R555 B.n27 B.n26 163.367
R556 B.n28 B.n27 163.367
R557 B.n420 B.n28 163.367
R558 B.n420 B.n33 163.367
R559 B.n34 B.n33 163.367
R560 B.n35 B.n34 163.367
R561 B.n425 B.n35 163.367
R562 B.n425 B.n40 163.367
R563 B.n41 B.n40 163.367
R564 B.n42 B.n41 163.367
R565 B.n430 B.n42 163.367
R566 B.n430 B.n47 163.367
R567 B.n48 B.n47 163.367
R568 B.n49 B.n48 163.367
R569 B.n435 B.n49 163.367
R570 B.n435 B.n54 163.367
R571 B.n55 B.n54 163.367
R572 B.n56 B.n55 163.367
R573 B.n440 B.n56 163.367
R574 B.n440 B.n61 163.367
R575 B.n62 B.n61 163.367
R576 B.n63 B.n62 163.367
R577 B.n445 B.n63 163.367
R578 B.n445 B.n68 163.367
R579 B.n69 B.n68 163.367
R580 B.n70 B.n69 163.367
R581 B.n87 B.n70 163.367
R582 B.n94 B.n74 163.367
R583 B.n98 B.n97 163.367
R584 B.n102 B.n101 163.367
R585 B.n106 B.n105 163.367
R586 B.n110 B.n109 163.367
R587 B.n114 B.n113 163.367
R588 B.n118 B.n117 163.367
R589 B.n122 B.n121 163.367
R590 B.n126 B.n125 163.367
R591 B.n130 B.n129 163.367
R592 B.n134 B.n133 163.367
R593 B.n136 B.n86 163.367
R594 B.n287 B.n211 126.032
R595 B.n287 B.n207 126.032
R596 B.n293 B.n207 126.032
R597 B.n293 B.n203 126.032
R598 B.n299 B.n203 126.032
R599 B.n299 B.n199 126.032
R600 B.n306 B.n199 126.032
R601 B.n306 B.n305 126.032
R602 B.n312 B.n192 126.032
R603 B.n318 B.n192 126.032
R604 B.n318 B.n188 126.032
R605 B.n324 B.n188 126.032
R606 B.n324 B.n184 126.032
R607 B.n330 B.n184 126.032
R608 B.n330 B.n180 126.032
R609 B.n336 B.n180 126.032
R610 B.n336 B.n176 126.032
R611 B.n342 B.n176 126.032
R612 B.n342 B.n172 126.032
R613 B.n348 B.n172 126.032
R614 B.n354 B.n168 126.032
R615 B.n354 B.n164 126.032
R616 B.n360 B.n164 126.032
R617 B.n360 B.n160 126.032
R618 B.n366 B.n160 126.032
R619 B.n366 B.n156 126.032
R620 B.n372 B.n156 126.032
R621 B.n372 B.n152 126.032
R622 B.n379 B.n152 126.032
R623 B.n379 B.n378 126.032
R624 B.n385 B.n145 126.032
R625 B.n392 B.n145 126.032
R626 B.n392 B.n141 126.032
R627 B.n398 B.n141 126.032
R628 B.n398 B.n4 126.032
R629 B.n535 B.n4 126.032
R630 B.n535 B.n534 126.032
R631 B.n534 B.n533 126.032
R632 B.n533 B.n8 126.032
R633 B.n527 B.n8 126.032
R634 B.n527 B.n526 126.032
R635 B.n526 B.n525 126.032
R636 B.n519 B.n18 126.032
R637 B.n519 B.n518 126.032
R638 B.n518 B.n517 126.032
R639 B.n517 B.n22 126.032
R640 B.n511 B.n22 126.032
R641 B.n511 B.n510 126.032
R642 B.n510 B.n509 126.032
R643 B.n509 B.n29 126.032
R644 B.n503 B.n29 126.032
R645 B.n503 B.n502 126.032
R646 B.n501 B.n36 126.032
R647 B.n495 B.n36 126.032
R648 B.n495 B.n494 126.032
R649 B.n494 B.n493 126.032
R650 B.n493 B.n43 126.032
R651 B.n487 B.n43 126.032
R652 B.n487 B.n486 126.032
R653 B.n486 B.n485 126.032
R654 B.n485 B.n50 126.032
R655 B.n479 B.n50 126.032
R656 B.n479 B.n478 126.032
R657 B.n478 B.n477 126.032
R658 B.n471 B.n60 126.032
R659 B.n471 B.n470 126.032
R660 B.n470 B.n469 126.032
R661 B.n469 B.n64 126.032
R662 B.n463 B.n64 126.032
R663 B.n463 B.n462 126.032
R664 B.n462 B.n461 126.032
R665 B.n461 B.n71 126.032
R666 B.n348 B.t1 103.791
R667 B.t3 B.n501 103.791
R668 B.n385 B.t2 100.085
R669 B.n525 B.t0 100.085
R670 B.n312 B.t5 96.3779
R671 B.n477 B.t9 96.3779
R672 B.n282 B.n281 71.676
R673 B.n227 B.n215 71.676
R674 B.n274 B.n216 71.676
R675 B.n270 B.n217 71.676
R676 B.n265 B.n218 71.676
R677 B.n261 B.n219 71.676
R678 B.n257 B.n220 71.676
R679 B.n253 B.n221 71.676
R680 B.n249 B.n222 71.676
R681 B.n244 B.n223 71.676
R682 B.n240 B.n224 71.676
R683 B.n236 B.n225 71.676
R684 B.n456 B.n455 71.676
R685 B.n94 B.n75 71.676
R686 B.n98 B.n76 71.676
R687 B.n102 B.n77 71.676
R688 B.n106 B.n78 71.676
R689 B.n110 B.n79 71.676
R690 B.n114 B.n80 71.676
R691 B.n118 B.n81 71.676
R692 B.n122 B.n82 71.676
R693 B.n126 B.n83 71.676
R694 B.n130 B.n84 71.676
R695 B.n134 B.n85 71.676
R696 B.n453 B.n86 71.676
R697 B.n453 B.n452 71.676
R698 B.n136 B.n85 71.676
R699 B.n133 B.n84 71.676
R700 B.n129 B.n83 71.676
R701 B.n125 B.n82 71.676
R702 B.n121 B.n81 71.676
R703 B.n117 B.n80 71.676
R704 B.n113 B.n79 71.676
R705 B.n109 B.n78 71.676
R706 B.n105 B.n77 71.676
R707 B.n101 B.n76 71.676
R708 B.n97 B.n75 71.676
R709 B.n455 B.n74 71.676
R710 B.n281 B.n214 71.676
R711 B.n275 B.n215 71.676
R712 B.n271 B.n216 71.676
R713 B.n266 B.n217 71.676
R714 B.n262 B.n218 71.676
R715 B.n258 B.n219 71.676
R716 B.n254 B.n220 71.676
R717 B.n250 B.n221 71.676
R718 B.n245 B.n222 71.676
R719 B.n241 B.n223 71.676
R720 B.n237 B.n224 71.676
R721 B.n233 B.n225 71.676
R722 B.n231 B.n230 68.4611
R723 B.n229 B.n228 68.4611
R724 B.n92 B.n91 68.4611
R725 B.n89 B.n88 68.4611
R726 B.n247 B.n231 59.5399
R727 B.n268 B.n229 59.5399
R728 B.n93 B.n92 59.5399
R729 B.n90 B.n89 59.5399
R730 B.n451 B.n450 35.7468
R731 B.n458 B.n457 35.7468
R732 B.n232 B.n209 35.7468
R733 B.n284 B.n283 35.7468
R734 B.n305 B.t5 29.6551
R735 B.n60 B.t9 29.6551
R736 B.n378 B.t2 25.9483
R737 B.n18 B.t0 25.9483
R738 B.t1 B.n168 22.2414
R739 B.n502 B.t3 22.2414
R740 B B.n537 18.0485
R741 B.n457 B.n73 10.6151
R742 B.n95 B.n73 10.6151
R743 B.n96 B.n95 10.6151
R744 B.n99 B.n96 10.6151
R745 B.n100 B.n99 10.6151
R746 B.n103 B.n100 10.6151
R747 B.n104 B.n103 10.6151
R748 B.n108 B.n107 10.6151
R749 B.n111 B.n108 10.6151
R750 B.n112 B.n111 10.6151
R751 B.n115 B.n112 10.6151
R752 B.n116 B.n115 10.6151
R753 B.n119 B.n116 10.6151
R754 B.n120 B.n119 10.6151
R755 B.n123 B.n120 10.6151
R756 B.n124 B.n123 10.6151
R757 B.n128 B.n127 10.6151
R758 B.n131 B.n128 10.6151
R759 B.n132 B.n131 10.6151
R760 B.n135 B.n132 10.6151
R761 B.n137 B.n135 10.6151
R762 B.n138 B.n137 10.6151
R763 B.n451 B.n138 10.6151
R764 B.n289 B.n209 10.6151
R765 B.n290 B.n289 10.6151
R766 B.n291 B.n290 10.6151
R767 B.n291 B.n201 10.6151
R768 B.n301 B.n201 10.6151
R769 B.n302 B.n301 10.6151
R770 B.n303 B.n302 10.6151
R771 B.n303 B.n194 10.6151
R772 B.n314 B.n194 10.6151
R773 B.n315 B.n314 10.6151
R774 B.n316 B.n315 10.6151
R775 B.n316 B.n186 10.6151
R776 B.n326 B.n186 10.6151
R777 B.n327 B.n326 10.6151
R778 B.n328 B.n327 10.6151
R779 B.n328 B.n178 10.6151
R780 B.n338 B.n178 10.6151
R781 B.n339 B.n338 10.6151
R782 B.n340 B.n339 10.6151
R783 B.n340 B.n170 10.6151
R784 B.n350 B.n170 10.6151
R785 B.n351 B.n350 10.6151
R786 B.n352 B.n351 10.6151
R787 B.n352 B.n162 10.6151
R788 B.n362 B.n162 10.6151
R789 B.n363 B.n362 10.6151
R790 B.n364 B.n363 10.6151
R791 B.n364 B.n154 10.6151
R792 B.n374 B.n154 10.6151
R793 B.n375 B.n374 10.6151
R794 B.n376 B.n375 10.6151
R795 B.n376 B.n147 10.6151
R796 B.n387 B.n147 10.6151
R797 B.n388 B.n387 10.6151
R798 B.n390 B.n388 10.6151
R799 B.n390 B.n389 10.6151
R800 B.n389 B.n139 10.6151
R801 B.n401 B.n139 10.6151
R802 B.n402 B.n401 10.6151
R803 B.n403 B.n402 10.6151
R804 B.n404 B.n403 10.6151
R805 B.n406 B.n404 10.6151
R806 B.n407 B.n406 10.6151
R807 B.n408 B.n407 10.6151
R808 B.n409 B.n408 10.6151
R809 B.n411 B.n409 10.6151
R810 B.n412 B.n411 10.6151
R811 B.n413 B.n412 10.6151
R812 B.n414 B.n413 10.6151
R813 B.n416 B.n414 10.6151
R814 B.n417 B.n416 10.6151
R815 B.n418 B.n417 10.6151
R816 B.n419 B.n418 10.6151
R817 B.n421 B.n419 10.6151
R818 B.n422 B.n421 10.6151
R819 B.n423 B.n422 10.6151
R820 B.n424 B.n423 10.6151
R821 B.n426 B.n424 10.6151
R822 B.n427 B.n426 10.6151
R823 B.n428 B.n427 10.6151
R824 B.n429 B.n428 10.6151
R825 B.n431 B.n429 10.6151
R826 B.n432 B.n431 10.6151
R827 B.n433 B.n432 10.6151
R828 B.n434 B.n433 10.6151
R829 B.n436 B.n434 10.6151
R830 B.n437 B.n436 10.6151
R831 B.n438 B.n437 10.6151
R832 B.n439 B.n438 10.6151
R833 B.n441 B.n439 10.6151
R834 B.n442 B.n441 10.6151
R835 B.n443 B.n442 10.6151
R836 B.n444 B.n443 10.6151
R837 B.n446 B.n444 10.6151
R838 B.n447 B.n446 10.6151
R839 B.n448 B.n447 10.6151
R840 B.n449 B.n448 10.6151
R841 B.n450 B.n449 10.6151
R842 B.n283 B.n213 10.6151
R843 B.n278 B.n213 10.6151
R844 B.n278 B.n277 10.6151
R845 B.n277 B.n276 10.6151
R846 B.n276 B.n273 10.6151
R847 B.n273 B.n272 10.6151
R848 B.n272 B.n269 10.6151
R849 B.n267 B.n264 10.6151
R850 B.n264 B.n263 10.6151
R851 B.n263 B.n260 10.6151
R852 B.n260 B.n259 10.6151
R853 B.n259 B.n256 10.6151
R854 B.n256 B.n255 10.6151
R855 B.n255 B.n252 10.6151
R856 B.n252 B.n251 10.6151
R857 B.n251 B.n248 10.6151
R858 B.n246 B.n243 10.6151
R859 B.n243 B.n242 10.6151
R860 B.n242 B.n239 10.6151
R861 B.n239 B.n238 10.6151
R862 B.n238 B.n235 10.6151
R863 B.n235 B.n234 10.6151
R864 B.n234 B.n232 10.6151
R865 B.n285 B.n284 10.6151
R866 B.n285 B.n205 10.6151
R867 B.n295 B.n205 10.6151
R868 B.n296 B.n295 10.6151
R869 B.n297 B.n296 10.6151
R870 B.n297 B.n197 10.6151
R871 B.n308 B.n197 10.6151
R872 B.n309 B.n308 10.6151
R873 B.n310 B.n309 10.6151
R874 B.n310 B.n190 10.6151
R875 B.n320 B.n190 10.6151
R876 B.n321 B.n320 10.6151
R877 B.n322 B.n321 10.6151
R878 B.n322 B.n182 10.6151
R879 B.n332 B.n182 10.6151
R880 B.n333 B.n332 10.6151
R881 B.n334 B.n333 10.6151
R882 B.n334 B.n174 10.6151
R883 B.n344 B.n174 10.6151
R884 B.n345 B.n344 10.6151
R885 B.n346 B.n345 10.6151
R886 B.n346 B.n166 10.6151
R887 B.n356 B.n166 10.6151
R888 B.n357 B.n356 10.6151
R889 B.n358 B.n357 10.6151
R890 B.n358 B.n158 10.6151
R891 B.n368 B.n158 10.6151
R892 B.n369 B.n368 10.6151
R893 B.n370 B.n369 10.6151
R894 B.n370 B.n150 10.6151
R895 B.n381 B.n150 10.6151
R896 B.n382 B.n381 10.6151
R897 B.n383 B.n382 10.6151
R898 B.n383 B.n143 10.6151
R899 B.n394 B.n143 10.6151
R900 B.n395 B.n394 10.6151
R901 B.n396 B.n395 10.6151
R902 B.n396 B.n0 10.6151
R903 B.n531 B.n1 10.6151
R904 B.n531 B.n530 10.6151
R905 B.n530 B.n529 10.6151
R906 B.n529 B.n10 10.6151
R907 B.n523 B.n10 10.6151
R908 B.n523 B.n522 10.6151
R909 B.n522 B.n521 10.6151
R910 B.n521 B.n16 10.6151
R911 B.n515 B.n16 10.6151
R912 B.n515 B.n514 10.6151
R913 B.n514 B.n513 10.6151
R914 B.n513 B.n24 10.6151
R915 B.n507 B.n24 10.6151
R916 B.n507 B.n506 10.6151
R917 B.n506 B.n505 10.6151
R918 B.n505 B.n31 10.6151
R919 B.n499 B.n31 10.6151
R920 B.n499 B.n498 10.6151
R921 B.n498 B.n497 10.6151
R922 B.n497 B.n38 10.6151
R923 B.n491 B.n38 10.6151
R924 B.n491 B.n490 10.6151
R925 B.n490 B.n489 10.6151
R926 B.n489 B.n45 10.6151
R927 B.n483 B.n45 10.6151
R928 B.n483 B.n482 10.6151
R929 B.n482 B.n481 10.6151
R930 B.n481 B.n52 10.6151
R931 B.n475 B.n52 10.6151
R932 B.n475 B.n474 10.6151
R933 B.n474 B.n473 10.6151
R934 B.n473 B.n58 10.6151
R935 B.n467 B.n58 10.6151
R936 B.n467 B.n466 10.6151
R937 B.n466 B.n465 10.6151
R938 B.n465 B.n66 10.6151
R939 B.n459 B.n66 10.6151
R940 B.n459 B.n458 10.6151
R941 B.n104 B.n93 9.52245
R942 B.n127 B.n90 9.52245
R943 B.n269 B.n268 9.52245
R944 B.n247 B.n246 9.52245
R945 B.n537 B.n0 2.81026
R946 B.n537 B.n1 2.81026
R947 B.n107 B.n93 1.09318
R948 B.n124 B.n90 1.09318
R949 B.n268 B.n267 1.09318
R950 B.n248 B.n247 1.09318
R951 VP.n17 VP.n16 161.3
R952 VP.n15 VP.n1 161.3
R953 VP.n14 VP.n13 161.3
R954 VP.n12 VP.n2 161.3
R955 VP.n11 VP.n10 161.3
R956 VP.n9 VP.n3 161.3
R957 VP.n8 VP.n7 161.3
R958 VP.n6 VP.n4 76.989
R959 VP.n18 VP.n0 76.989
R960 VP.n6 VP.n5 42.1887
R961 VP.n10 VP.n2 40.4106
R962 VP.n14 VP.n2 40.4106
R963 VP.n5 VP.t3 39.5417
R964 VP.n5 VP.t2 38.4474
R965 VP.n9 VP.n8 24.3439
R966 VP.n10 VP.n9 24.3439
R967 VP.n15 VP.n14 24.3439
R968 VP.n16 VP.n15 24.3439
R969 VP.n8 VP.n4 12.9025
R970 VP.n16 VP.n0 12.9025
R971 VP.n4 VP.t0 4.97112
R972 VP.n0 VP.t1 4.97112
R973 VP.n7 VP.n6 0.355081
R974 VP.n18 VP.n17 0.355081
R975 VP VP.n18 0.26685
R976 VP.n7 VP.n3 0.189894
R977 VP.n11 VP.n3 0.189894
R978 VP.n12 VP.n11 0.189894
R979 VP.n13 VP.n12 0.189894
R980 VP.n13 VP.n1 0.189894
R981 VP.n17 VP.n1 0.189894
R982 VDD1 VDD1.n1 268.966
R983 VDD1 VDD1.n0 235.085
R984 VDD1.n0 VDD1.t1 30.0005
R985 VDD1.n0 VDD1.t2 30.0005
R986 VDD1.n1 VDD1.t0 30.0005
R987 VDD1.n1 VDD1.t3 30.0005
R988 VTAIL.n7 VTAIL.t3 248.349
R989 VTAIL.n0 VTAIL.t0 248.349
R990 VTAIL.n1 VTAIL.t6 248.349
R991 VTAIL.n2 VTAIL.t7 248.349
R992 VTAIL.n6 VTAIL.t5 248.349
R993 VTAIL.n5 VTAIL.t4 248.349
R994 VTAIL.n4 VTAIL.t2 248.349
R995 VTAIL.n3 VTAIL.t1 248.349
R996 VTAIL.n7 VTAIL.n6 15.9789
R997 VTAIL.n3 VTAIL.n2 15.9789
R998 VTAIL.n4 VTAIL.n3 3.0436
R999 VTAIL.n6 VTAIL.n5 3.0436
R1000 VTAIL.n2 VTAIL.n1 3.0436
R1001 VTAIL VTAIL.n0 1.58024
R1002 VTAIL VTAIL.n7 1.46386
R1003 VTAIL.n5 VTAIL.n4 0.470328
R1004 VTAIL.n1 VTAIL.n0 0.470328
R1005 VN VN.n1 42.3542
R1006 VN.n1 VN.t1 39.5418
R1007 VN.n0 VN.t3 39.5418
R1008 VN.n1 VN.t0 38.4474
R1009 VN.n0 VN.t2 38.4474
R1010 VN VN.n0 2.63069
R1011 VDD2.n2 VDD2.n0 268.44
R1012 VDD2.n2 VDD2.n1 235.028
R1013 VDD2.n1 VDD2.t3 30.0005
R1014 VDD2.n1 VDD2.t2 30.0005
R1015 VDD2.n0 VDD2.t0 30.0005
R1016 VDD2.n0 VDD2.t1 30.0005
R1017 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 1.51828f
C1 VP VTAIL 1.53238f
C2 VDD2 VTAIL 3.10391f
C3 VN VDD1 0.156638f
C4 VP VDD1 0.877654f
C5 VDD2 VDD1 1.17328f
C6 VP VN 4.54124f
C7 VDD2 VP 0.441415f
C8 VDD2 VN 0.595918f
C9 VTAIL VDD1 3.04568f
C10 VDD2 B 3.212089f
C11 VDD1 B 6.01608f
C12 VTAIL B 3.007083f
C13 VN B 10.73898f
C14 VP B 9.165438f
C15 VDD2.t0 B 0.01442f
C16 VDD2.t1 B 0.01442f
C17 VDD2.n0 B 0.141209f
C18 VDD2.t3 B 0.01442f
C19 VDD2.t2 B 0.01442f
C20 VDD2.n1 B 0.036066f
C21 VDD2.n2 B 2.58797f
C22 VN.t2 B 0.307108f
C23 VN.t3 B 0.316047f
C24 VN.n0 B 0.271124f
C25 VN.t0 B 0.307108f
C26 VN.t1 B 0.316047f
C27 VN.n1 B 1.53137f
C28 VTAIL.t0 B 0.06485f
C29 VTAIL.n0 B 0.231051f
C30 VTAIL.t6 B 0.06485f
C31 VTAIL.n1 B 0.363832f
C32 VTAIL.t7 B 0.06485f
C33 VTAIL.n2 B 1.03147f
C34 VTAIL.t1 B 0.06485f
C35 VTAIL.n3 B 1.03147f
C36 VTAIL.t2 B 0.06485f
C37 VTAIL.n4 B 0.363832f
C38 VTAIL.t4 B 0.06485f
C39 VTAIL.n5 B 0.363832f
C40 VTAIL.t5 B 0.06485f
C41 VTAIL.n6 B 1.03147f
C42 VTAIL.t3 B 0.06485f
C43 VTAIL.n7 B 0.888127f
C44 VDD1.t1 B 0.01351f
C45 VDD1.t2 B 0.01351f
C46 VDD1.n0 B 0.033873f
C47 VDD1.t0 B 0.01351f
C48 VDD1.t3 B 0.01351f
C49 VDD1.n1 B 0.140248f
C50 VP.t1 B 0.077163f
C51 VP.n0 B 0.178676f
C52 VP.n1 B 0.026889f
C53 VP.n2 B 0.021759f
C54 VP.n3 B 0.026889f
C55 VP.t0 B 0.077163f
C56 VP.n4 B 0.178675f
C57 VP.t3 B 0.318701f
C58 VP.t2 B 0.309687f
C59 VP.n5 B 1.53262f
C60 VP.n6 B 1.1822f
C61 VP.n7 B 0.043405f
C62 VP.n8 B 0.038678f
C63 VP.n9 B 0.050365f
C64 VP.n10 B 0.053727f
C65 VP.n11 B 0.026889f
C66 VP.n12 B 0.026889f
C67 VP.n13 B 0.026889f
C68 VP.n14 B 0.053727f
C69 VP.n15 B 0.050365f
C70 VP.n16 B 0.038678f
C71 VP.n17 B 0.043405f
C72 VP.n18 B 0.065752f
.ends

