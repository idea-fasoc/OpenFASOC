* NGSPICE file created from diff_pair_sample_1035.ext - technology: sky130A

.subckt diff_pair_sample_1035 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X1 VDD2.t9 VN.t0 VTAIL.t2 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=1.88595 ps=11.76 w=11.43 l=2.81
X2 VTAIL.t1 VN.t1 VDD2.t8 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X3 VTAIL.t10 VP.t1 VDD1.t8 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X4 VTAIL.t14 VP.t2 VDD1.t7 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X5 B.t11 B.t9 B.t10 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=0 ps=0 w=11.43 l=2.81
X6 VTAIL.t16 VN.t2 VDD2.t7 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X7 VDD2.t6 VN.t3 VTAIL.t15 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=4.4577 ps=23.64 w=11.43 l=2.81
X8 VTAIL.t3 VN.t4 VDD2.t5 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X9 B.t8 B.t6 B.t7 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=0 ps=0 w=11.43 l=2.81
X10 VDD1.t6 VP.t3 VTAIL.t9 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=1.88595 ps=11.76 w=11.43 l=2.81
X11 VDD1.t5 VP.t4 VTAIL.t5 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X12 VDD2.t4 VN.t5 VTAIL.t4 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=4.4577 ps=23.64 w=11.43 l=2.81
X13 VDD2.t3 VN.t6 VTAIL.t0 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X14 VTAIL.t18 VN.t7 VDD2.t2 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X15 B.t5 B.t3 B.t4 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=0 ps=0 w=11.43 l=2.81
X16 VTAIL.t6 VP.t5 VDD1.t4 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X17 VDD2.t1 VN.t8 VTAIL.t19 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=1.88595 ps=11.76 w=11.43 l=2.81
X18 VTAIL.t8 VP.t6 VDD1.t3 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X19 VDD1.t2 VP.t7 VTAIL.t13 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=1.88595 ps=11.76 w=11.43 l=2.81
X20 VDD2.t0 VN.t9 VTAIL.t17 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=1.88595 ps=11.76 w=11.43 l=2.81
X21 VDD1.t1 VP.t8 VTAIL.t7 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=4.4577 ps=23.64 w=11.43 l=2.81
X22 VDD1.t0 VP.t9 VTAIL.t12 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=1.88595 pd=11.76 as=4.4577 ps=23.64 w=11.43 l=2.81
X23 B.t2 B.t0 B.t1 w_n4738_n3254# sky130_fd_pr__pfet_01v8 ad=4.4577 pd=23.64 as=0 ps=0 w=11.43 l=2.81
R0 VP.n26 VP.n23 161.3
R1 VP.n28 VP.n27 161.3
R2 VP.n29 VP.n22 161.3
R3 VP.n31 VP.n30 161.3
R4 VP.n32 VP.n21 161.3
R5 VP.n34 VP.n33 161.3
R6 VP.n36 VP.n20 161.3
R7 VP.n38 VP.n37 161.3
R8 VP.n39 VP.n19 161.3
R9 VP.n41 VP.n40 161.3
R10 VP.n42 VP.n18 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n17 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n49 VP.n16 161.3
R15 VP.n51 VP.n50 161.3
R16 VP.n52 VP.n15 161.3
R17 VP.n54 VP.n53 161.3
R18 VP.n55 VP.n14 161.3
R19 VP.n100 VP.n0 161.3
R20 VP.n99 VP.n98 161.3
R21 VP.n97 VP.n1 161.3
R22 VP.n96 VP.n95 161.3
R23 VP.n94 VP.n2 161.3
R24 VP.n93 VP.n92 161.3
R25 VP.n91 VP.n3 161.3
R26 VP.n90 VP.n89 161.3
R27 VP.n87 VP.n4 161.3
R28 VP.n86 VP.n85 161.3
R29 VP.n84 VP.n5 161.3
R30 VP.n83 VP.n82 161.3
R31 VP.n81 VP.n6 161.3
R32 VP.n79 VP.n78 161.3
R33 VP.n77 VP.n7 161.3
R34 VP.n76 VP.n75 161.3
R35 VP.n74 VP.n8 161.3
R36 VP.n73 VP.n72 161.3
R37 VP.n71 VP.n9 161.3
R38 VP.n70 VP.n69 161.3
R39 VP.n67 VP.n10 161.3
R40 VP.n66 VP.n65 161.3
R41 VP.n64 VP.n11 161.3
R42 VP.n63 VP.n62 161.3
R43 VP.n61 VP.n12 161.3
R44 VP.n60 VP.n59 161.3
R45 VP.n25 VP.t7 130.656
R46 VP.n58 VP.n13 109.288
R47 VP.n102 VP.n101 109.288
R48 VP.n57 VP.n56 109.288
R49 VP.n13 VP.t3 98.03
R50 VP.n68 VP.t1 98.03
R51 VP.n80 VP.t4 98.03
R52 VP.n88 VP.t2 98.03
R53 VP.n101 VP.t8 98.03
R54 VP.n56 VP.t9 98.03
R55 VP.n43 VP.t5 98.03
R56 VP.n35 VP.t0 98.03
R57 VP.n24 VP.t6 98.03
R58 VP.n75 VP.n74 56.5193
R59 VP.n41 VP.n19 56.5193
R60 VP.n86 VP.n5 56.5193
R61 VP.n30 VP.n29 56.5193
R62 VP.n25 VP.n24 54.5315
R63 VP.n58 VP.n57 53.7647
R64 VP.n66 VP.n11 44.3785
R65 VP.n95 VP.n94 44.3785
R66 VP.n50 VP.n49 44.3785
R67 VP.n62 VP.n11 36.6083
R68 VP.n95 VP.n1 36.6083
R69 VP.n50 VP.n15 36.6083
R70 VP.n61 VP.n60 24.4675
R71 VP.n62 VP.n61 24.4675
R72 VP.n67 VP.n66 24.4675
R73 VP.n69 VP.n67 24.4675
R74 VP.n73 VP.n9 24.4675
R75 VP.n74 VP.n73 24.4675
R76 VP.n75 VP.n7 24.4675
R77 VP.n79 VP.n7 24.4675
R78 VP.n82 VP.n81 24.4675
R79 VP.n82 VP.n5 24.4675
R80 VP.n87 VP.n86 24.4675
R81 VP.n89 VP.n87 24.4675
R82 VP.n93 VP.n3 24.4675
R83 VP.n94 VP.n93 24.4675
R84 VP.n99 VP.n1 24.4675
R85 VP.n100 VP.n99 24.4675
R86 VP.n54 VP.n15 24.4675
R87 VP.n55 VP.n54 24.4675
R88 VP.n42 VP.n41 24.4675
R89 VP.n44 VP.n42 24.4675
R90 VP.n48 VP.n17 24.4675
R91 VP.n49 VP.n48 24.4675
R92 VP.n30 VP.n21 24.4675
R93 VP.n34 VP.n21 24.4675
R94 VP.n37 VP.n36 24.4675
R95 VP.n37 VP.n19 24.4675
R96 VP.n28 VP.n23 24.4675
R97 VP.n29 VP.n28 24.4675
R98 VP.n68 VP.n9 19.0848
R99 VP.n89 VP.n88 19.0848
R100 VP.n44 VP.n43 19.0848
R101 VP.n24 VP.n23 19.0848
R102 VP.n80 VP.n79 12.234
R103 VP.n81 VP.n80 12.234
R104 VP.n35 VP.n34 12.234
R105 VP.n36 VP.n35 12.234
R106 VP.n69 VP.n68 5.38324
R107 VP.n88 VP.n3 5.38324
R108 VP.n43 VP.n17 5.38324
R109 VP.n26 VP.n25 5.13245
R110 VP.n60 VP.n13 1.46852
R111 VP.n101 VP.n100 1.46852
R112 VP.n56 VP.n55 1.46852
R113 VP.n57 VP.n14 0.278367
R114 VP.n59 VP.n58 0.278367
R115 VP.n102 VP.n0 0.278367
R116 VP.n27 VP.n26 0.189894
R117 VP.n27 VP.n22 0.189894
R118 VP.n31 VP.n22 0.189894
R119 VP.n32 VP.n31 0.189894
R120 VP.n33 VP.n32 0.189894
R121 VP.n33 VP.n20 0.189894
R122 VP.n38 VP.n20 0.189894
R123 VP.n39 VP.n38 0.189894
R124 VP.n40 VP.n39 0.189894
R125 VP.n40 VP.n18 0.189894
R126 VP.n45 VP.n18 0.189894
R127 VP.n46 VP.n45 0.189894
R128 VP.n47 VP.n46 0.189894
R129 VP.n47 VP.n16 0.189894
R130 VP.n51 VP.n16 0.189894
R131 VP.n52 VP.n51 0.189894
R132 VP.n53 VP.n52 0.189894
R133 VP.n53 VP.n14 0.189894
R134 VP.n59 VP.n12 0.189894
R135 VP.n63 VP.n12 0.189894
R136 VP.n64 VP.n63 0.189894
R137 VP.n65 VP.n64 0.189894
R138 VP.n65 VP.n10 0.189894
R139 VP.n70 VP.n10 0.189894
R140 VP.n71 VP.n70 0.189894
R141 VP.n72 VP.n71 0.189894
R142 VP.n72 VP.n8 0.189894
R143 VP.n76 VP.n8 0.189894
R144 VP.n77 VP.n76 0.189894
R145 VP.n78 VP.n77 0.189894
R146 VP.n78 VP.n6 0.189894
R147 VP.n83 VP.n6 0.189894
R148 VP.n84 VP.n83 0.189894
R149 VP.n85 VP.n84 0.189894
R150 VP.n85 VP.n4 0.189894
R151 VP.n90 VP.n4 0.189894
R152 VP.n91 VP.n90 0.189894
R153 VP.n92 VP.n91 0.189894
R154 VP.n92 VP.n2 0.189894
R155 VP.n96 VP.n2 0.189894
R156 VP.n97 VP.n96 0.189894
R157 VP.n98 VP.n97 0.189894
R158 VP.n98 VP.n0 0.189894
R159 VP VP.n102 0.153454
R160 VTAIL.n256 VTAIL.n200 756.745
R161 VTAIL.n58 VTAIL.n2 756.745
R162 VTAIL.n194 VTAIL.n138 756.745
R163 VTAIL.n128 VTAIL.n72 756.745
R164 VTAIL.n221 VTAIL.n220 585
R165 VTAIL.n223 VTAIL.n222 585
R166 VTAIL.n216 VTAIL.n215 585
R167 VTAIL.n229 VTAIL.n228 585
R168 VTAIL.n231 VTAIL.n230 585
R169 VTAIL.n212 VTAIL.n211 585
R170 VTAIL.n238 VTAIL.n237 585
R171 VTAIL.n239 VTAIL.n210 585
R172 VTAIL.n241 VTAIL.n240 585
R173 VTAIL.n208 VTAIL.n207 585
R174 VTAIL.n247 VTAIL.n246 585
R175 VTAIL.n249 VTAIL.n248 585
R176 VTAIL.n204 VTAIL.n203 585
R177 VTAIL.n255 VTAIL.n254 585
R178 VTAIL.n257 VTAIL.n256 585
R179 VTAIL.n23 VTAIL.n22 585
R180 VTAIL.n25 VTAIL.n24 585
R181 VTAIL.n18 VTAIL.n17 585
R182 VTAIL.n31 VTAIL.n30 585
R183 VTAIL.n33 VTAIL.n32 585
R184 VTAIL.n14 VTAIL.n13 585
R185 VTAIL.n40 VTAIL.n39 585
R186 VTAIL.n41 VTAIL.n12 585
R187 VTAIL.n43 VTAIL.n42 585
R188 VTAIL.n10 VTAIL.n9 585
R189 VTAIL.n49 VTAIL.n48 585
R190 VTAIL.n51 VTAIL.n50 585
R191 VTAIL.n6 VTAIL.n5 585
R192 VTAIL.n57 VTAIL.n56 585
R193 VTAIL.n59 VTAIL.n58 585
R194 VTAIL.n195 VTAIL.n194 585
R195 VTAIL.n193 VTAIL.n192 585
R196 VTAIL.n142 VTAIL.n141 585
R197 VTAIL.n187 VTAIL.n186 585
R198 VTAIL.n185 VTAIL.n184 585
R199 VTAIL.n146 VTAIL.n145 585
R200 VTAIL.n150 VTAIL.n148 585
R201 VTAIL.n179 VTAIL.n178 585
R202 VTAIL.n177 VTAIL.n176 585
R203 VTAIL.n152 VTAIL.n151 585
R204 VTAIL.n171 VTAIL.n170 585
R205 VTAIL.n169 VTAIL.n168 585
R206 VTAIL.n156 VTAIL.n155 585
R207 VTAIL.n163 VTAIL.n162 585
R208 VTAIL.n161 VTAIL.n160 585
R209 VTAIL.n129 VTAIL.n128 585
R210 VTAIL.n127 VTAIL.n126 585
R211 VTAIL.n76 VTAIL.n75 585
R212 VTAIL.n121 VTAIL.n120 585
R213 VTAIL.n119 VTAIL.n118 585
R214 VTAIL.n80 VTAIL.n79 585
R215 VTAIL.n84 VTAIL.n82 585
R216 VTAIL.n113 VTAIL.n112 585
R217 VTAIL.n111 VTAIL.n110 585
R218 VTAIL.n86 VTAIL.n85 585
R219 VTAIL.n105 VTAIL.n104 585
R220 VTAIL.n103 VTAIL.n102 585
R221 VTAIL.n90 VTAIL.n89 585
R222 VTAIL.n97 VTAIL.n96 585
R223 VTAIL.n95 VTAIL.n94 585
R224 VTAIL.n219 VTAIL.t4 329.036
R225 VTAIL.n21 VTAIL.t7 329.036
R226 VTAIL.n159 VTAIL.t12 329.036
R227 VTAIL.n93 VTAIL.t15 329.036
R228 VTAIL.n222 VTAIL.n221 171.744
R229 VTAIL.n222 VTAIL.n215 171.744
R230 VTAIL.n229 VTAIL.n215 171.744
R231 VTAIL.n230 VTAIL.n229 171.744
R232 VTAIL.n230 VTAIL.n211 171.744
R233 VTAIL.n238 VTAIL.n211 171.744
R234 VTAIL.n239 VTAIL.n238 171.744
R235 VTAIL.n240 VTAIL.n239 171.744
R236 VTAIL.n240 VTAIL.n207 171.744
R237 VTAIL.n247 VTAIL.n207 171.744
R238 VTAIL.n248 VTAIL.n247 171.744
R239 VTAIL.n248 VTAIL.n203 171.744
R240 VTAIL.n255 VTAIL.n203 171.744
R241 VTAIL.n256 VTAIL.n255 171.744
R242 VTAIL.n24 VTAIL.n23 171.744
R243 VTAIL.n24 VTAIL.n17 171.744
R244 VTAIL.n31 VTAIL.n17 171.744
R245 VTAIL.n32 VTAIL.n31 171.744
R246 VTAIL.n32 VTAIL.n13 171.744
R247 VTAIL.n40 VTAIL.n13 171.744
R248 VTAIL.n41 VTAIL.n40 171.744
R249 VTAIL.n42 VTAIL.n41 171.744
R250 VTAIL.n42 VTAIL.n9 171.744
R251 VTAIL.n49 VTAIL.n9 171.744
R252 VTAIL.n50 VTAIL.n49 171.744
R253 VTAIL.n50 VTAIL.n5 171.744
R254 VTAIL.n57 VTAIL.n5 171.744
R255 VTAIL.n58 VTAIL.n57 171.744
R256 VTAIL.n194 VTAIL.n193 171.744
R257 VTAIL.n193 VTAIL.n141 171.744
R258 VTAIL.n186 VTAIL.n141 171.744
R259 VTAIL.n186 VTAIL.n185 171.744
R260 VTAIL.n185 VTAIL.n145 171.744
R261 VTAIL.n150 VTAIL.n145 171.744
R262 VTAIL.n178 VTAIL.n150 171.744
R263 VTAIL.n178 VTAIL.n177 171.744
R264 VTAIL.n177 VTAIL.n151 171.744
R265 VTAIL.n170 VTAIL.n151 171.744
R266 VTAIL.n170 VTAIL.n169 171.744
R267 VTAIL.n169 VTAIL.n155 171.744
R268 VTAIL.n162 VTAIL.n155 171.744
R269 VTAIL.n162 VTAIL.n161 171.744
R270 VTAIL.n128 VTAIL.n127 171.744
R271 VTAIL.n127 VTAIL.n75 171.744
R272 VTAIL.n120 VTAIL.n75 171.744
R273 VTAIL.n120 VTAIL.n119 171.744
R274 VTAIL.n119 VTAIL.n79 171.744
R275 VTAIL.n84 VTAIL.n79 171.744
R276 VTAIL.n112 VTAIL.n84 171.744
R277 VTAIL.n112 VTAIL.n111 171.744
R278 VTAIL.n111 VTAIL.n85 171.744
R279 VTAIL.n104 VTAIL.n85 171.744
R280 VTAIL.n104 VTAIL.n103 171.744
R281 VTAIL.n103 VTAIL.n89 171.744
R282 VTAIL.n96 VTAIL.n89 171.744
R283 VTAIL.n96 VTAIL.n95 171.744
R284 VTAIL.n221 VTAIL.t4 85.8723
R285 VTAIL.n23 VTAIL.t7 85.8723
R286 VTAIL.n161 VTAIL.t12 85.8723
R287 VTAIL.n95 VTAIL.t15 85.8723
R288 VTAIL.n137 VTAIL.n136 58.686
R289 VTAIL.n135 VTAIL.n134 58.686
R290 VTAIL.n71 VTAIL.n70 58.686
R291 VTAIL.n69 VTAIL.n68 58.686
R292 VTAIL.n263 VTAIL.n262 58.6858
R293 VTAIL.n1 VTAIL.n0 58.6858
R294 VTAIL.n65 VTAIL.n64 58.6858
R295 VTAIL.n67 VTAIL.n66 58.6858
R296 VTAIL.n261 VTAIL.n260 32.7672
R297 VTAIL.n63 VTAIL.n62 32.7672
R298 VTAIL.n199 VTAIL.n198 32.7672
R299 VTAIL.n133 VTAIL.n132 32.7672
R300 VTAIL.n69 VTAIL.n67 27.6341
R301 VTAIL.n261 VTAIL.n199 24.9272
R302 VTAIL.n241 VTAIL.n208 13.1884
R303 VTAIL.n43 VTAIL.n10 13.1884
R304 VTAIL.n148 VTAIL.n146 13.1884
R305 VTAIL.n82 VTAIL.n80 13.1884
R306 VTAIL.n242 VTAIL.n210 12.8005
R307 VTAIL.n246 VTAIL.n245 12.8005
R308 VTAIL.n44 VTAIL.n12 12.8005
R309 VTAIL.n48 VTAIL.n47 12.8005
R310 VTAIL.n184 VTAIL.n183 12.8005
R311 VTAIL.n180 VTAIL.n179 12.8005
R312 VTAIL.n118 VTAIL.n117 12.8005
R313 VTAIL.n114 VTAIL.n113 12.8005
R314 VTAIL.n237 VTAIL.n236 12.0247
R315 VTAIL.n249 VTAIL.n206 12.0247
R316 VTAIL.n39 VTAIL.n38 12.0247
R317 VTAIL.n51 VTAIL.n8 12.0247
R318 VTAIL.n187 VTAIL.n144 12.0247
R319 VTAIL.n176 VTAIL.n149 12.0247
R320 VTAIL.n121 VTAIL.n78 12.0247
R321 VTAIL.n110 VTAIL.n83 12.0247
R322 VTAIL.n235 VTAIL.n212 11.249
R323 VTAIL.n250 VTAIL.n204 11.249
R324 VTAIL.n37 VTAIL.n14 11.249
R325 VTAIL.n52 VTAIL.n6 11.249
R326 VTAIL.n188 VTAIL.n142 11.249
R327 VTAIL.n175 VTAIL.n152 11.249
R328 VTAIL.n122 VTAIL.n76 11.249
R329 VTAIL.n109 VTAIL.n86 11.249
R330 VTAIL.n220 VTAIL.n219 10.7239
R331 VTAIL.n22 VTAIL.n21 10.7239
R332 VTAIL.n160 VTAIL.n159 10.7239
R333 VTAIL.n94 VTAIL.n93 10.7239
R334 VTAIL.n232 VTAIL.n231 10.4732
R335 VTAIL.n254 VTAIL.n253 10.4732
R336 VTAIL.n34 VTAIL.n33 10.4732
R337 VTAIL.n56 VTAIL.n55 10.4732
R338 VTAIL.n192 VTAIL.n191 10.4732
R339 VTAIL.n172 VTAIL.n171 10.4732
R340 VTAIL.n126 VTAIL.n125 10.4732
R341 VTAIL.n106 VTAIL.n105 10.4732
R342 VTAIL.n228 VTAIL.n214 9.69747
R343 VTAIL.n257 VTAIL.n202 9.69747
R344 VTAIL.n30 VTAIL.n16 9.69747
R345 VTAIL.n59 VTAIL.n4 9.69747
R346 VTAIL.n195 VTAIL.n140 9.69747
R347 VTAIL.n168 VTAIL.n154 9.69747
R348 VTAIL.n129 VTAIL.n74 9.69747
R349 VTAIL.n102 VTAIL.n88 9.69747
R350 VTAIL.n260 VTAIL.n259 9.45567
R351 VTAIL.n62 VTAIL.n61 9.45567
R352 VTAIL.n198 VTAIL.n197 9.45567
R353 VTAIL.n132 VTAIL.n131 9.45567
R354 VTAIL.n259 VTAIL.n258 9.3005
R355 VTAIL.n202 VTAIL.n201 9.3005
R356 VTAIL.n253 VTAIL.n252 9.3005
R357 VTAIL.n251 VTAIL.n250 9.3005
R358 VTAIL.n206 VTAIL.n205 9.3005
R359 VTAIL.n245 VTAIL.n244 9.3005
R360 VTAIL.n218 VTAIL.n217 9.3005
R361 VTAIL.n225 VTAIL.n224 9.3005
R362 VTAIL.n227 VTAIL.n226 9.3005
R363 VTAIL.n214 VTAIL.n213 9.3005
R364 VTAIL.n233 VTAIL.n232 9.3005
R365 VTAIL.n235 VTAIL.n234 9.3005
R366 VTAIL.n236 VTAIL.n209 9.3005
R367 VTAIL.n243 VTAIL.n242 9.3005
R368 VTAIL.n61 VTAIL.n60 9.3005
R369 VTAIL.n4 VTAIL.n3 9.3005
R370 VTAIL.n55 VTAIL.n54 9.3005
R371 VTAIL.n53 VTAIL.n52 9.3005
R372 VTAIL.n8 VTAIL.n7 9.3005
R373 VTAIL.n47 VTAIL.n46 9.3005
R374 VTAIL.n20 VTAIL.n19 9.3005
R375 VTAIL.n27 VTAIL.n26 9.3005
R376 VTAIL.n29 VTAIL.n28 9.3005
R377 VTAIL.n16 VTAIL.n15 9.3005
R378 VTAIL.n35 VTAIL.n34 9.3005
R379 VTAIL.n37 VTAIL.n36 9.3005
R380 VTAIL.n38 VTAIL.n11 9.3005
R381 VTAIL.n45 VTAIL.n44 9.3005
R382 VTAIL.n158 VTAIL.n157 9.3005
R383 VTAIL.n165 VTAIL.n164 9.3005
R384 VTAIL.n167 VTAIL.n166 9.3005
R385 VTAIL.n154 VTAIL.n153 9.3005
R386 VTAIL.n173 VTAIL.n172 9.3005
R387 VTAIL.n175 VTAIL.n174 9.3005
R388 VTAIL.n149 VTAIL.n147 9.3005
R389 VTAIL.n181 VTAIL.n180 9.3005
R390 VTAIL.n197 VTAIL.n196 9.3005
R391 VTAIL.n140 VTAIL.n139 9.3005
R392 VTAIL.n191 VTAIL.n190 9.3005
R393 VTAIL.n189 VTAIL.n188 9.3005
R394 VTAIL.n144 VTAIL.n143 9.3005
R395 VTAIL.n183 VTAIL.n182 9.3005
R396 VTAIL.n92 VTAIL.n91 9.3005
R397 VTAIL.n99 VTAIL.n98 9.3005
R398 VTAIL.n101 VTAIL.n100 9.3005
R399 VTAIL.n88 VTAIL.n87 9.3005
R400 VTAIL.n107 VTAIL.n106 9.3005
R401 VTAIL.n109 VTAIL.n108 9.3005
R402 VTAIL.n83 VTAIL.n81 9.3005
R403 VTAIL.n115 VTAIL.n114 9.3005
R404 VTAIL.n131 VTAIL.n130 9.3005
R405 VTAIL.n74 VTAIL.n73 9.3005
R406 VTAIL.n125 VTAIL.n124 9.3005
R407 VTAIL.n123 VTAIL.n122 9.3005
R408 VTAIL.n78 VTAIL.n77 9.3005
R409 VTAIL.n117 VTAIL.n116 9.3005
R410 VTAIL.n227 VTAIL.n216 8.92171
R411 VTAIL.n258 VTAIL.n200 8.92171
R412 VTAIL.n29 VTAIL.n18 8.92171
R413 VTAIL.n60 VTAIL.n2 8.92171
R414 VTAIL.n196 VTAIL.n138 8.92171
R415 VTAIL.n167 VTAIL.n156 8.92171
R416 VTAIL.n130 VTAIL.n72 8.92171
R417 VTAIL.n101 VTAIL.n90 8.92171
R418 VTAIL.n224 VTAIL.n223 8.14595
R419 VTAIL.n26 VTAIL.n25 8.14595
R420 VTAIL.n164 VTAIL.n163 8.14595
R421 VTAIL.n98 VTAIL.n97 8.14595
R422 VTAIL.n220 VTAIL.n218 7.3702
R423 VTAIL.n22 VTAIL.n20 7.3702
R424 VTAIL.n160 VTAIL.n158 7.3702
R425 VTAIL.n94 VTAIL.n92 7.3702
R426 VTAIL.n223 VTAIL.n218 5.81868
R427 VTAIL.n25 VTAIL.n20 5.81868
R428 VTAIL.n163 VTAIL.n158 5.81868
R429 VTAIL.n97 VTAIL.n92 5.81868
R430 VTAIL.n224 VTAIL.n216 5.04292
R431 VTAIL.n260 VTAIL.n200 5.04292
R432 VTAIL.n26 VTAIL.n18 5.04292
R433 VTAIL.n62 VTAIL.n2 5.04292
R434 VTAIL.n198 VTAIL.n138 5.04292
R435 VTAIL.n164 VTAIL.n156 5.04292
R436 VTAIL.n132 VTAIL.n72 5.04292
R437 VTAIL.n98 VTAIL.n90 5.04292
R438 VTAIL.n228 VTAIL.n227 4.26717
R439 VTAIL.n258 VTAIL.n257 4.26717
R440 VTAIL.n30 VTAIL.n29 4.26717
R441 VTAIL.n60 VTAIL.n59 4.26717
R442 VTAIL.n196 VTAIL.n195 4.26717
R443 VTAIL.n168 VTAIL.n167 4.26717
R444 VTAIL.n130 VTAIL.n129 4.26717
R445 VTAIL.n102 VTAIL.n101 4.26717
R446 VTAIL.n231 VTAIL.n214 3.49141
R447 VTAIL.n254 VTAIL.n202 3.49141
R448 VTAIL.n33 VTAIL.n16 3.49141
R449 VTAIL.n56 VTAIL.n4 3.49141
R450 VTAIL.n192 VTAIL.n140 3.49141
R451 VTAIL.n171 VTAIL.n154 3.49141
R452 VTAIL.n126 VTAIL.n74 3.49141
R453 VTAIL.n105 VTAIL.n88 3.49141
R454 VTAIL.n262 VTAIL.t17 2.84433
R455 VTAIL.n262 VTAIL.t1 2.84433
R456 VTAIL.n0 VTAIL.t2 2.84433
R457 VTAIL.n0 VTAIL.t16 2.84433
R458 VTAIL.n64 VTAIL.t5 2.84433
R459 VTAIL.n64 VTAIL.t14 2.84433
R460 VTAIL.n66 VTAIL.t9 2.84433
R461 VTAIL.n66 VTAIL.t10 2.84433
R462 VTAIL.n136 VTAIL.t11 2.84433
R463 VTAIL.n136 VTAIL.t6 2.84433
R464 VTAIL.n134 VTAIL.t13 2.84433
R465 VTAIL.n134 VTAIL.t8 2.84433
R466 VTAIL.n70 VTAIL.t0 2.84433
R467 VTAIL.n70 VTAIL.t3 2.84433
R468 VTAIL.n68 VTAIL.t19 2.84433
R469 VTAIL.n68 VTAIL.t18 2.84433
R470 VTAIL.n232 VTAIL.n212 2.71565
R471 VTAIL.n253 VTAIL.n204 2.71565
R472 VTAIL.n34 VTAIL.n14 2.71565
R473 VTAIL.n55 VTAIL.n6 2.71565
R474 VTAIL.n191 VTAIL.n142 2.71565
R475 VTAIL.n172 VTAIL.n152 2.71565
R476 VTAIL.n125 VTAIL.n76 2.71565
R477 VTAIL.n106 VTAIL.n86 2.71565
R478 VTAIL.n71 VTAIL.n69 2.7074
R479 VTAIL.n133 VTAIL.n71 2.7074
R480 VTAIL.n137 VTAIL.n135 2.7074
R481 VTAIL.n199 VTAIL.n137 2.7074
R482 VTAIL.n67 VTAIL.n65 2.7074
R483 VTAIL.n65 VTAIL.n63 2.7074
R484 VTAIL.n263 VTAIL.n261 2.7074
R485 VTAIL.n219 VTAIL.n217 2.41282
R486 VTAIL.n21 VTAIL.n19 2.41282
R487 VTAIL.n159 VTAIL.n157 2.41282
R488 VTAIL.n93 VTAIL.n91 2.41282
R489 VTAIL VTAIL.n1 2.08886
R490 VTAIL.n237 VTAIL.n235 1.93989
R491 VTAIL.n250 VTAIL.n249 1.93989
R492 VTAIL.n39 VTAIL.n37 1.93989
R493 VTAIL.n52 VTAIL.n51 1.93989
R494 VTAIL.n188 VTAIL.n187 1.93989
R495 VTAIL.n176 VTAIL.n175 1.93989
R496 VTAIL.n122 VTAIL.n121 1.93989
R497 VTAIL.n110 VTAIL.n109 1.93989
R498 VTAIL.n135 VTAIL.n133 1.82378
R499 VTAIL.n63 VTAIL.n1 1.82378
R500 VTAIL.n236 VTAIL.n210 1.16414
R501 VTAIL.n246 VTAIL.n206 1.16414
R502 VTAIL.n38 VTAIL.n12 1.16414
R503 VTAIL.n48 VTAIL.n8 1.16414
R504 VTAIL.n184 VTAIL.n144 1.16414
R505 VTAIL.n179 VTAIL.n149 1.16414
R506 VTAIL.n118 VTAIL.n78 1.16414
R507 VTAIL.n113 VTAIL.n83 1.16414
R508 VTAIL VTAIL.n263 0.619035
R509 VTAIL.n242 VTAIL.n241 0.388379
R510 VTAIL.n245 VTAIL.n208 0.388379
R511 VTAIL.n44 VTAIL.n43 0.388379
R512 VTAIL.n47 VTAIL.n10 0.388379
R513 VTAIL.n183 VTAIL.n146 0.388379
R514 VTAIL.n180 VTAIL.n148 0.388379
R515 VTAIL.n117 VTAIL.n80 0.388379
R516 VTAIL.n114 VTAIL.n82 0.388379
R517 VTAIL.n225 VTAIL.n217 0.155672
R518 VTAIL.n226 VTAIL.n225 0.155672
R519 VTAIL.n226 VTAIL.n213 0.155672
R520 VTAIL.n233 VTAIL.n213 0.155672
R521 VTAIL.n234 VTAIL.n233 0.155672
R522 VTAIL.n234 VTAIL.n209 0.155672
R523 VTAIL.n243 VTAIL.n209 0.155672
R524 VTAIL.n244 VTAIL.n243 0.155672
R525 VTAIL.n244 VTAIL.n205 0.155672
R526 VTAIL.n251 VTAIL.n205 0.155672
R527 VTAIL.n252 VTAIL.n251 0.155672
R528 VTAIL.n252 VTAIL.n201 0.155672
R529 VTAIL.n259 VTAIL.n201 0.155672
R530 VTAIL.n27 VTAIL.n19 0.155672
R531 VTAIL.n28 VTAIL.n27 0.155672
R532 VTAIL.n28 VTAIL.n15 0.155672
R533 VTAIL.n35 VTAIL.n15 0.155672
R534 VTAIL.n36 VTAIL.n35 0.155672
R535 VTAIL.n36 VTAIL.n11 0.155672
R536 VTAIL.n45 VTAIL.n11 0.155672
R537 VTAIL.n46 VTAIL.n45 0.155672
R538 VTAIL.n46 VTAIL.n7 0.155672
R539 VTAIL.n53 VTAIL.n7 0.155672
R540 VTAIL.n54 VTAIL.n53 0.155672
R541 VTAIL.n54 VTAIL.n3 0.155672
R542 VTAIL.n61 VTAIL.n3 0.155672
R543 VTAIL.n197 VTAIL.n139 0.155672
R544 VTAIL.n190 VTAIL.n139 0.155672
R545 VTAIL.n190 VTAIL.n189 0.155672
R546 VTAIL.n189 VTAIL.n143 0.155672
R547 VTAIL.n182 VTAIL.n143 0.155672
R548 VTAIL.n182 VTAIL.n181 0.155672
R549 VTAIL.n181 VTAIL.n147 0.155672
R550 VTAIL.n174 VTAIL.n147 0.155672
R551 VTAIL.n174 VTAIL.n173 0.155672
R552 VTAIL.n173 VTAIL.n153 0.155672
R553 VTAIL.n166 VTAIL.n153 0.155672
R554 VTAIL.n166 VTAIL.n165 0.155672
R555 VTAIL.n165 VTAIL.n157 0.155672
R556 VTAIL.n131 VTAIL.n73 0.155672
R557 VTAIL.n124 VTAIL.n73 0.155672
R558 VTAIL.n124 VTAIL.n123 0.155672
R559 VTAIL.n123 VTAIL.n77 0.155672
R560 VTAIL.n116 VTAIL.n77 0.155672
R561 VTAIL.n116 VTAIL.n115 0.155672
R562 VTAIL.n115 VTAIL.n81 0.155672
R563 VTAIL.n108 VTAIL.n81 0.155672
R564 VTAIL.n108 VTAIL.n107 0.155672
R565 VTAIL.n107 VTAIL.n87 0.155672
R566 VTAIL.n100 VTAIL.n87 0.155672
R567 VTAIL.n100 VTAIL.n99 0.155672
R568 VTAIL.n99 VTAIL.n91 0.155672
R569 VDD1.n56 VDD1.n0 756.745
R570 VDD1.n119 VDD1.n63 756.745
R571 VDD1.n57 VDD1.n56 585
R572 VDD1.n55 VDD1.n54 585
R573 VDD1.n4 VDD1.n3 585
R574 VDD1.n49 VDD1.n48 585
R575 VDD1.n47 VDD1.n46 585
R576 VDD1.n8 VDD1.n7 585
R577 VDD1.n12 VDD1.n10 585
R578 VDD1.n41 VDD1.n40 585
R579 VDD1.n39 VDD1.n38 585
R580 VDD1.n14 VDD1.n13 585
R581 VDD1.n33 VDD1.n32 585
R582 VDD1.n31 VDD1.n30 585
R583 VDD1.n18 VDD1.n17 585
R584 VDD1.n25 VDD1.n24 585
R585 VDD1.n23 VDD1.n22 585
R586 VDD1.n84 VDD1.n83 585
R587 VDD1.n86 VDD1.n85 585
R588 VDD1.n79 VDD1.n78 585
R589 VDD1.n92 VDD1.n91 585
R590 VDD1.n94 VDD1.n93 585
R591 VDD1.n75 VDD1.n74 585
R592 VDD1.n101 VDD1.n100 585
R593 VDD1.n102 VDD1.n73 585
R594 VDD1.n104 VDD1.n103 585
R595 VDD1.n71 VDD1.n70 585
R596 VDD1.n110 VDD1.n109 585
R597 VDD1.n112 VDD1.n111 585
R598 VDD1.n67 VDD1.n66 585
R599 VDD1.n118 VDD1.n117 585
R600 VDD1.n120 VDD1.n119 585
R601 VDD1.n21 VDD1.t2 329.036
R602 VDD1.n82 VDD1.t6 329.036
R603 VDD1.n56 VDD1.n55 171.744
R604 VDD1.n55 VDD1.n3 171.744
R605 VDD1.n48 VDD1.n3 171.744
R606 VDD1.n48 VDD1.n47 171.744
R607 VDD1.n47 VDD1.n7 171.744
R608 VDD1.n12 VDD1.n7 171.744
R609 VDD1.n40 VDD1.n12 171.744
R610 VDD1.n40 VDD1.n39 171.744
R611 VDD1.n39 VDD1.n13 171.744
R612 VDD1.n32 VDD1.n13 171.744
R613 VDD1.n32 VDD1.n31 171.744
R614 VDD1.n31 VDD1.n17 171.744
R615 VDD1.n24 VDD1.n17 171.744
R616 VDD1.n24 VDD1.n23 171.744
R617 VDD1.n85 VDD1.n84 171.744
R618 VDD1.n85 VDD1.n78 171.744
R619 VDD1.n92 VDD1.n78 171.744
R620 VDD1.n93 VDD1.n92 171.744
R621 VDD1.n93 VDD1.n74 171.744
R622 VDD1.n101 VDD1.n74 171.744
R623 VDD1.n102 VDD1.n101 171.744
R624 VDD1.n103 VDD1.n102 171.744
R625 VDD1.n103 VDD1.n70 171.744
R626 VDD1.n110 VDD1.n70 171.744
R627 VDD1.n111 VDD1.n110 171.744
R628 VDD1.n111 VDD1.n66 171.744
R629 VDD1.n118 VDD1.n66 171.744
R630 VDD1.n119 VDD1.n118 171.744
R631 VDD1.n23 VDD1.t2 85.8723
R632 VDD1.n84 VDD1.t6 85.8723
R633 VDD1.n127 VDD1.n126 77.3394
R634 VDD1.n62 VDD1.n61 75.3648
R635 VDD1.n129 VDD1.n128 75.3646
R636 VDD1.n125 VDD1.n124 75.3646
R637 VDD1.n62 VDD1.n60 52.1529
R638 VDD1.n125 VDD1.n123 52.1529
R639 VDD1.n129 VDD1.n127 48.363
R640 VDD1.n10 VDD1.n8 13.1884
R641 VDD1.n104 VDD1.n71 13.1884
R642 VDD1.n46 VDD1.n45 12.8005
R643 VDD1.n42 VDD1.n41 12.8005
R644 VDD1.n105 VDD1.n73 12.8005
R645 VDD1.n109 VDD1.n108 12.8005
R646 VDD1.n49 VDD1.n6 12.0247
R647 VDD1.n38 VDD1.n11 12.0247
R648 VDD1.n100 VDD1.n99 12.0247
R649 VDD1.n112 VDD1.n69 12.0247
R650 VDD1.n50 VDD1.n4 11.249
R651 VDD1.n37 VDD1.n14 11.249
R652 VDD1.n98 VDD1.n75 11.249
R653 VDD1.n113 VDD1.n67 11.249
R654 VDD1.n22 VDD1.n21 10.7239
R655 VDD1.n83 VDD1.n82 10.7239
R656 VDD1.n54 VDD1.n53 10.4732
R657 VDD1.n34 VDD1.n33 10.4732
R658 VDD1.n95 VDD1.n94 10.4732
R659 VDD1.n117 VDD1.n116 10.4732
R660 VDD1.n57 VDD1.n2 9.69747
R661 VDD1.n30 VDD1.n16 9.69747
R662 VDD1.n91 VDD1.n77 9.69747
R663 VDD1.n120 VDD1.n65 9.69747
R664 VDD1.n60 VDD1.n59 9.45567
R665 VDD1.n123 VDD1.n122 9.45567
R666 VDD1.n20 VDD1.n19 9.3005
R667 VDD1.n27 VDD1.n26 9.3005
R668 VDD1.n29 VDD1.n28 9.3005
R669 VDD1.n16 VDD1.n15 9.3005
R670 VDD1.n35 VDD1.n34 9.3005
R671 VDD1.n37 VDD1.n36 9.3005
R672 VDD1.n11 VDD1.n9 9.3005
R673 VDD1.n43 VDD1.n42 9.3005
R674 VDD1.n59 VDD1.n58 9.3005
R675 VDD1.n2 VDD1.n1 9.3005
R676 VDD1.n53 VDD1.n52 9.3005
R677 VDD1.n51 VDD1.n50 9.3005
R678 VDD1.n6 VDD1.n5 9.3005
R679 VDD1.n45 VDD1.n44 9.3005
R680 VDD1.n122 VDD1.n121 9.3005
R681 VDD1.n65 VDD1.n64 9.3005
R682 VDD1.n116 VDD1.n115 9.3005
R683 VDD1.n114 VDD1.n113 9.3005
R684 VDD1.n69 VDD1.n68 9.3005
R685 VDD1.n108 VDD1.n107 9.3005
R686 VDD1.n81 VDD1.n80 9.3005
R687 VDD1.n88 VDD1.n87 9.3005
R688 VDD1.n90 VDD1.n89 9.3005
R689 VDD1.n77 VDD1.n76 9.3005
R690 VDD1.n96 VDD1.n95 9.3005
R691 VDD1.n98 VDD1.n97 9.3005
R692 VDD1.n99 VDD1.n72 9.3005
R693 VDD1.n106 VDD1.n105 9.3005
R694 VDD1.n58 VDD1.n0 8.92171
R695 VDD1.n29 VDD1.n18 8.92171
R696 VDD1.n90 VDD1.n79 8.92171
R697 VDD1.n121 VDD1.n63 8.92171
R698 VDD1.n26 VDD1.n25 8.14595
R699 VDD1.n87 VDD1.n86 8.14595
R700 VDD1.n22 VDD1.n20 7.3702
R701 VDD1.n83 VDD1.n81 7.3702
R702 VDD1.n25 VDD1.n20 5.81868
R703 VDD1.n86 VDD1.n81 5.81868
R704 VDD1.n60 VDD1.n0 5.04292
R705 VDD1.n26 VDD1.n18 5.04292
R706 VDD1.n87 VDD1.n79 5.04292
R707 VDD1.n123 VDD1.n63 5.04292
R708 VDD1.n58 VDD1.n57 4.26717
R709 VDD1.n30 VDD1.n29 4.26717
R710 VDD1.n91 VDD1.n90 4.26717
R711 VDD1.n121 VDD1.n120 4.26717
R712 VDD1.n54 VDD1.n2 3.49141
R713 VDD1.n33 VDD1.n16 3.49141
R714 VDD1.n94 VDD1.n77 3.49141
R715 VDD1.n117 VDD1.n65 3.49141
R716 VDD1.n128 VDD1.t4 2.84433
R717 VDD1.n128 VDD1.t0 2.84433
R718 VDD1.n61 VDD1.t3 2.84433
R719 VDD1.n61 VDD1.t9 2.84433
R720 VDD1.n126 VDD1.t7 2.84433
R721 VDD1.n126 VDD1.t1 2.84433
R722 VDD1.n124 VDD1.t8 2.84433
R723 VDD1.n124 VDD1.t5 2.84433
R724 VDD1.n53 VDD1.n4 2.71565
R725 VDD1.n34 VDD1.n14 2.71565
R726 VDD1.n95 VDD1.n75 2.71565
R727 VDD1.n116 VDD1.n67 2.71565
R728 VDD1.n21 VDD1.n19 2.41282
R729 VDD1.n82 VDD1.n80 2.41282
R730 VDD1 VDD1.n129 1.97248
R731 VDD1.n50 VDD1.n49 1.93989
R732 VDD1.n38 VDD1.n37 1.93989
R733 VDD1.n100 VDD1.n98 1.93989
R734 VDD1.n113 VDD1.n112 1.93989
R735 VDD1.n46 VDD1.n6 1.16414
R736 VDD1.n41 VDD1.n11 1.16414
R737 VDD1.n99 VDD1.n73 1.16414
R738 VDD1.n109 VDD1.n69 1.16414
R739 VDD1 VDD1.n62 0.735414
R740 VDD1.n127 VDD1.n125 0.621878
R741 VDD1.n45 VDD1.n8 0.388379
R742 VDD1.n42 VDD1.n10 0.388379
R743 VDD1.n105 VDD1.n104 0.388379
R744 VDD1.n108 VDD1.n71 0.388379
R745 VDD1.n59 VDD1.n1 0.155672
R746 VDD1.n52 VDD1.n1 0.155672
R747 VDD1.n52 VDD1.n51 0.155672
R748 VDD1.n51 VDD1.n5 0.155672
R749 VDD1.n44 VDD1.n5 0.155672
R750 VDD1.n44 VDD1.n43 0.155672
R751 VDD1.n43 VDD1.n9 0.155672
R752 VDD1.n36 VDD1.n9 0.155672
R753 VDD1.n36 VDD1.n35 0.155672
R754 VDD1.n35 VDD1.n15 0.155672
R755 VDD1.n28 VDD1.n15 0.155672
R756 VDD1.n28 VDD1.n27 0.155672
R757 VDD1.n27 VDD1.n19 0.155672
R758 VDD1.n88 VDD1.n80 0.155672
R759 VDD1.n89 VDD1.n88 0.155672
R760 VDD1.n89 VDD1.n76 0.155672
R761 VDD1.n96 VDD1.n76 0.155672
R762 VDD1.n97 VDD1.n96 0.155672
R763 VDD1.n97 VDD1.n72 0.155672
R764 VDD1.n106 VDD1.n72 0.155672
R765 VDD1.n107 VDD1.n106 0.155672
R766 VDD1.n107 VDD1.n68 0.155672
R767 VDD1.n114 VDD1.n68 0.155672
R768 VDD1.n115 VDD1.n114 0.155672
R769 VDD1.n115 VDD1.n64 0.155672
R770 VDD1.n122 VDD1.n64 0.155672
R771 VN.n85 VN.n44 161.3
R772 VN.n84 VN.n83 161.3
R773 VN.n82 VN.n45 161.3
R774 VN.n81 VN.n80 161.3
R775 VN.n79 VN.n46 161.3
R776 VN.n78 VN.n77 161.3
R777 VN.n76 VN.n47 161.3
R778 VN.n75 VN.n74 161.3
R779 VN.n73 VN.n48 161.3
R780 VN.n72 VN.n71 161.3
R781 VN.n70 VN.n50 161.3
R782 VN.n69 VN.n68 161.3
R783 VN.n67 VN.n51 161.3
R784 VN.n65 VN.n64 161.3
R785 VN.n63 VN.n52 161.3
R786 VN.n62 VN.n61 161.3
R787 VN.n60 VN.n53 161.3
R788 VN.n59 VN.n58 161.3
R789 VN.n57 VN.n54 161.3
R790 VN.n41 VN.n0 161.3
R791 VN.n40 VN.n39 161.3
R792 VN.n38 VN.n1 161.3
R793 VN.n37 VN.n36 161.3
R794 VN.n35 VN.n2 161.3
R795 VN.n34 VN.n33 161.3
R796 VN.n32 VN.n3 161.3
R797 VN.n31 VN.n30 161.3
R798 VN.n28 VN.n4 161.3
R799 VN.n27 VN.n26 161.3
R800 VN.n25 VN.n5 161.3
R801 VN.n24 VN.n23 161.3
R802 VN.n22 VN.n6 161.3
R803 VN.n20 VN.n19 161.3
R804 VN.n18 VN.n7 161.3
R805 VN.n17 VN.n16 161.3
R806 VN.n15 VN.n8 161.3
R807 VN.n14 VN.n13 161.3
R808 VN.n12 VN.n9 161.3
R809 VN.n11 VN.t0 130.656
R810 VN.n56 VN.t3 130.656
R811 VN.n43 VN.n42 109.288
R812 VN.n87 VN.n86 109.288
R813 VN.n10 VN.t2 98.03
R814 VN.n21 VN.t9 98.03
R815 VN.n29 VN.t1 98.03
R816 VN.n42 VN.t5 98.03
R817 VN.n55 VN.t4 98.03
R818 VN.n66 VN.t6 98.03
R819 VN.n49 VN.t7 98.03
R820 VN.n86 VN.t8 98.03
R821 VN.n16 VN.n15 56.5193
R822 VN.n61 VN.n60 56.5193
R823 VN.n27 VN.n5 56.5193
R824 VN.n72 VN.n50 56.5193
R825 VN.n11 VN.n10 54.5315
R826 VN.n56 VN.n55 54.5315
R827 VN VN.n87 54.0436
R828 VN.n36 VN.n35 44.3785
R829 VN.n80 VN.n79 44.3785
R830 VN.n36 VN.n1 36.6083
R831 VN.n80 VN.n45 36.6083
R832 VN.n14 VN.n9 24.4675
R833 VN.n15 VN.n14 24.4675
R834 VN.n16 VN.n7 24.4675
R835 VN.n20 VN.n7 24.4675
R836 VN.n23 VN.n22 24.4675
R837 VN.n23 VN.n5 24.4675
R838 VN.n28 VN.n27 24.4675
R839 VN.n30 VN.n28 24.4675
R840 VN.n34 VN.n3 24.4675
R841 VN.n35 VN.n34 24.4675
R842 VN.n40 VN.n1 24.4675
R843 VN.n41 VN.n40 24.4675
R844 VN.n60 VN.n59 24.4675
R845 VN.n59 VN.n54 24.4675
R846 VN.n68 VN.n50 24.4675
R847 VN.n68 VN.n67 24.4675
R848 VN.n65 VN.n52 24.4675
R849 VN.n61 VN.n52 24.4675
R850 VN.n79 VN.n78 24.4675
R851 VN.n78 VN.n47 24.4675
R852 VN.n74 VN.n73 24.4675
R853 VN.n73 VN.n72 24.4675
R854 VN.n85 VN.n84 24.4675
R855 VN.n84 VN.n45 24.4675
R856 VN.n10 VN.n9 19.0848
R857 VN.n30 VN.n29 19.0848
R858 VN.n55 VN.n54 19.0848
R859 VN.n74 VN.n49 19.0848
R860 VN.n21 VN.n20 12.234
R861 VN.n22 VN.n21 12.234
R862 VN.n67 VN.n66 12.234
R863 VN.n66 VN.n65 12.234
R864 VN.n29 VN.n3 5.38324
R865 VN.n49 VN.n47 5.38324
R866 VN.n57 VN.n56 5.13245
R867 VN.n12 VN.n11 5.13245
R868 VN.n42 VN.n41 1.46852
R869 VN.n86 VN.n85 1.46852
R870 VN.n87 VN.n44 0.278367
R871 VN.n43 VN.n0 0.278367
R872 VN.n83 VN.n44 0.189894
R873 VN.n83 VN.n82 0.189894
R874 VN.n82 VN.n81 0.189894
R875 VN.n81 VN.n46 0.189894
R876 VN.n77 VN.n46 0.189894
R877 VN.n77 VN.n76 0.189894
R878 VN.n76 VN.n75 0.189894
R879 VN.n75 VN.n48 0.189894
R880 VN.n71 VN.n48 0.189894
R881 VN.n71 VN.n70 0.189894
R882 VN.n70 VN.n69 0.189894
R883 VN.n69 VN.n51 0.189894
R884 VN.n64 VN.n51 0.189894
R885 VN.n64 VN.n63 0.189894
R886 VN.n63 VN.n62 0.189894
R887 VN.n62 VN.n53 0.189894
R888 VN.n58 VN.n53 0.189894
R889 VN.n58 VN.n57 0.189894
R890 VN.n13 VN.n12 0.189894
R891 VN.n13 VN.n8 0.189894
R892 VN.n17 VN.n8 0.189894
R893 VN.n18 VN.n17 0.189894
R894 VN.n19 VN.n18 0.189894
R895 VN.n19 VN.n6 0.189894
R896 VN.n24 VN.n6 0.189894
R897 VN.n25 VN.n24 0.189894
R898 VN.n26 VN.n25 0.189894
R899 VN.n26 VN.n4 0.189894
R900 VN.n31 VN.n4 0.189894
R901 VN.n32 VN.n31 0.189894
R902 VN.n33 VN.n32 0.189894
R903 VN.n33 VN.n2 0.189894
R904 VN.n37 VN.n2 0.189894
R905 VN.n38 VN.n37 0.189894
R906 VN.n39 VN.n38 0.189894
R907 VN.n39 VN.n0 0.189894
R908 VN VN.n43 0.153454
R909 VDD2.n121 VDD2.n65 756.745
R910 VDD2.n56 VDD2.n0 756.745
R911 VDD2.n122 VDD2.n121 585
R912 VDD2.n120 VDD2.n119 585
R913 VDD2.n69 VDD2.n68 585
R914 VDD2.n114 VDD2.n113 585
R915 VDD2.n112 VDD2.n111 585
R916 VDD2.n73 VDD2.n72 585
R917 VDD2.n77 VDD2.n75 585
R918 VDD2.n106 VDD2.n105 585
R919 VDD2.n104 VDD2.n103 585
R920 VDD2.n79 VDD2.n78 585
R921 VDD2.n98 VDD2.n97 585
R922 VDD2.n96 VDD2.n95 585
R923 VDD2.n83 VDD2.n82 585
R924 VDD2.n90 VDD2.n89 585
R925 VDD2.n88 VDD2.n87 585
R926 VDD2.n21 VDD2.n20 585
R927 VDD2.n23 VDD2.n22 585
R928 VDD2.n16 VDD2.n15 585
R929 VDD2.n29 VDD2.n28 585
R930 VDD2.n31 VDD2.n30 585
R931 VDD2.n12 VDD2.n11 585
R932 VDD2.n38 VDD2.n37 585
R933 VDD2.n39 VDD2.n10 585
R934 VDD2.n41 VDD2.n40 585
R935 VDD2.n8 VDD2.n7 585
R936 VDD2.n47 VDD2.n46 585
R937 VDD2.n49 VDD2.n48 585
R938 VDD2.n4 VDD2.n3 585
R939 VDD2.n55 VDD2.n54 585
R940 VDD2.n57 VDD2.n56 585
R941 VDD2.n86 VDD2.t1 329.036
R942 VDD2.n19 VDD2.t9 329.036
R943 VDD2.n121 VDD2.n120 171.744
R944 VDD2.n120 VDD2.n68 171.744
R945 VDD2.n113 VDD2.n68 171.744
R946 VDD2.n113 VDD2.n112 171.744
R947 VDD2.n112 VDD2.n72 171.744
R948 VDD2.n77 VDD2.n72 171.744
R949 VDD2.n105 VDD2.n77 171.744
R950 VDD2.n105 VDD2.n104 171.744
R951 VDD2.n104 VDD2.n78 171.744
R952 VDD2.n97 VDD2.n78 171.744
R953 VDD2.n97 VDD2.n96 171.744
R954 VDD2.n96 VDD2.n82 171.744
R955 VDD2.n89 VDD2.n82 171.744
R956 VDD2.n89 VDD2.n88 171.744
R957 VDD2.n22 VDD2.n21 171.744
R958 VDD2.n22 VDD2.n15 171.744
R959 VDD2.n29 VDD2.n15 171.744
R960 VDD2.n30 VDD2.n29 171.744
R961 VDD2.n30 VDD2.n11 171.744
R962 VDD2.n38 VDD2.n11 171.744
R963 VDD2.n39 VDD2.n38 171.744
R964 VDD2.n40 VDD2.n39 171.744
R965 VDD2.n40 VDD2.n7 171.744
R966 VDD2.n47 VDD2.n7 171.744
R967 VDD2.n48 VDD2.n47 171.744
R968 VDD2.n48 VDD2.n3 171.744
R969 VDD2.n55 VDD2.n3 171.744
R970 VDD2.n56 VDD2.n55 171.744
R971 VDD2.n88 VDD2.t1 85.8723
R972 VDD2.n21 VDD2.t9 85.8723
R973 VDD2.n64 VDD2.n63 77.3394
R974 VDD2 VDD2.n129 77.3366
R975 VDD2.n128 VDD2.n127 75.3648
R976 VDD2.n62 VDD2.n61 75.3646
R977 VDD2.n62 VDD2.n60 52.1529
R978 VDD2.n126 VDD2.n125 49.446
R979 VDD2.n126 VDD2.n64 46.4265
R980 VDD2.n75 VDD2.n73 13.1884
R981 VDD2.n41 VDD2.n8 13.1884
R982 VDD2.n111 VDD2.n110 12.8005
R983 VDD2.n107 VDD2.n106 12.8005
R984 VDD2.n42 VDD2.n10 12.8005
R985 VDD2.n46 VDD2.n45 12.8005
R986 VDD2.n114 VDD2.n71 12.0247
R987 VDD2.n103 VDD2.n76 12.0247
R988 VDD2.n37 VDD2.n36 12.0247
R989 VDD2.n49 VDD2.n6 12.0247
R990 VDD2.n115 VDD2.n69 11.249
R991 VDD2.n102 VDD2.n79 11.249
R992 VDD2.n35 VDD2.n12 11.249
R993 VDD2.n50 VDD2.n4 11.249
R994 VDD2.n87 VDD2.n86 10.7239
R995 VDD2.n20 VDD2.n19 10.7239
R996 VDD2.n119 VDD2.n118 10.4732
R997 VDD2.n99 VDD2.n98 10.4732
R998 VDD2.n32 VDD2.n31 10.4732
R999 VDD2.n54 VDD2.n53 10.4732
R1000 VDD2.n122 VDD2.n67 9.69747
R1001 VDD2.n95 VDD2.n81 9.69747
R1002 VDD2.n28 VDD2.n14 9.69747
R1003 VDD2.n57 VDD2.n2 9.69747
R1004 VDD2.n125 VDD2.n124 9.45567
R1005 VDD2.n60 VDD2.n59 9.45567
R1006 VDD2.n85 VDD2.n84 9.3005
R1007 VDD2.n92 VDD2.n91 9.3005
R1008 VDD2.n94 VDD2.n93 9.3005
R1009 VDD2.n81 VDD2.n80 9.3005
R1010 VDD2.n100 VDD2.n99 9.3005
R1011 VDD2.n102 VDD2.n101 9.3005
R1012 VDD2.n76 VDD2.n74 9.3005
R1013 VDD2.n108 VDD2.n107 9.3005
R1014 VDD2.n124 VDD2.n123 9.3005
R1015 VDD2.n67 VDD2.n66 9.3005
R1016 VDD2.n118 VDD2.n117 9.3005
R1017 VDD2.n116 VDD2.n115 9.3005
R1018 VDD2.n71 VDD2.n70 9.3005
R1019 VDD2.n110 VDD2.n109 9.3005
R1020 VDD2.n59 VDD2.n58 9.3005
R1021 VDD2.n2 VDD2.n1 9.3005
R1022 VDD2.n53 VDD2.n52 9.3005
R1023 VDD2.n51 VDD2.n50 9.3005
R1024 VDD2.n6 VDD2.n5 9.3005
R1025 VDD2.n45 VDD2.n44 9.3005
R1026 VDD2.n18 VDD2.n17 9.3005
R1027 VDD2.n25 VDD2.n24 9.3005
R1028 VDD2.n27 VDD2.n26 9.3005
R1029 VDD2.n14 VDD2.n13 9.3005
R1030 VDD2.n33 VDD2.n32 9.3005
R1031 VDD2.n35 VDD2.n34 9.3005
R1032 VDD2.n36 VDD2.n9 9.3005
R1033 VDD2.n43 VDD2.n42 9.3005
R1034 VDD2.n123 VDD2.n65 8.92171
R1035 VDD2.n94 VDD2.n83 8.92171
R1036 VDD2.n27 VDD2.n16 8.92171
R1037 VDD2.n58 VDD2.n0 8.92171
R1038 VDD2.n91 VDD2.n90 8.14595
R1039 VDD2.n24 VDD2.n23 8.14595
R1040 VDD2.n87 VDD2.n85 7.3702
R1041 VDD2.n20 VDD2.n18 7.3702
R1042 VDD2.n90 VDD2.n85 5.81868
R1043 VDD2.n23 VDD2.n18 5.81868
R1044 VDD2.n125 VDD2.n65 5.04292
R1045 VDD2.n91 VDD2.n83 5.04292
R1046 VDD2.n24 VDD2.n16 5.04292
R1047 VDD2.n60 VDD2.n0 5.04292
R1048 VDD2.n123 VDD2.n122 4.26717
R1049 VDD2.n95 VDD2.n94 4.26717
R1050 VDD2.n28 VDD2.n27 4.26717
R1051 VDD2.n58 VDD2.n57 4.26717
R1052 VDD2.n119 VDD2.n67 3.49141
R1053 VDD2.n98 VDD2.n81 3.49141
R1054 VDD2.n31 VDD2.n14 3.49141
R1055 VDD2.n54 VDD2.n2 3.49141
R1056 VDD2.n129 VDD2.t5 2.84433
R1057 VDD2.n129 VDD2.t6 2.84433
R1058 VDD2.n127 VDD2.t2 2.84433
R1059 VDD2.n127 VDD2.t3 2.84433
R1060 VDD2.n63 VDD2.t8 2.84433
R1061 VDD2.n63 VDD2.t4 2.84433
R1062 VDD2.n61 VDD2.t7 2.84433
R1063 VDD2.n61 VDD2.t0 2.84433
R1064 VDD2.n118 VDD2.n69 2.71565
R1065 VDD2.n99 VDD2.n79 2.71565
R1066 VDD2.n32 VDD2.n12 2.71565
R1067 VDD2.n53 VDD2.n4 2.71565
R1068 VDD2.n128 VDD2.n126 2.7074
R1069 VDD2.n86 VDD2.n84 2.41282
R1070 VDD2.n19 VDD2.n17 2.41282
R1071 VDD2.n115 VDD2.n114 1.93989
R1072 VDD2.n103 VDD2.n102 1.93989
R1073 VDD2.n37 VDD2.n35 1.93989
R1074 VDD2.n50 VDD2.n49 1.93989
R1075 VDD2.n111 VDD2.n71 1.16414
R1076 VDD2.n106 VDD2.n76 1.16414
R1077 VDD2.n36 VDD2.n10 1.16414
R1078 VDD2.n46 VDD2.n6 1.16414
R1079 VDD2 VDD2.n128 0.735414
R1080 VDD2.n64 VDD2.n62 0.621878
R1081 VDD2.n110 VDD2.n73 0.388379
R1082 VDD2.n107 VDD2.n75 0.388379
R1083 VDD2.n42 VDD2.n41 0.388379
R1084 VDD2.n45 VDD2.n8 0.388379
R1085 VDD2.n124 VDD2.n66 0.155672
R1086 VDD2.n117 VDD2.n66 0.155672
R1087 VDD2.n117 VDD2.n116 0.155672
R1088 VDD2.n116 VDD2.n70 0.155672
R1089 VDD2.n109 VDD2.n70 0.155672
R1090 VDD2.n109 VDD2.n108 0.155672
R1091 VDD2.n108 VDD2.n74 0.155672
R1092 VDD2.n101 VDD2.n74 0.155672
R1093 VDD2.n101 VDD2.n100 0.155672
R1094 VDD2.n100 VDD2.n80 0.155672
R1095 VDD2.n93 VDD2.n80 0.155672
R1096 VDD2.n93 VDD2.n92 0.155672
R1097 VDD2.n92 VDD2.n84 0.155672
R1098 VDD2.n25 VDD2.n17 0.155672
R1099 VDD2.n26 VDD2.n25 0.155672
R1100 VDD2.n26 VDD2.n13 0.155672
R1101 VDD2.n33 VDD2.n13 0.155672
R1102 VDD2.n34 VDD2.n33 0.155672
R1103 VDD2.n34 VDD2.n9 0.155672
R1104 VDD2.n43 VDD2.n9 0.155672
R1105 VDD2.n44 VDD2.n43 0.155672
R1106 VDD2.n44 VDD2.n5 0.155672
R1107 VDD2.n51 VDD2.n5 0.155672
R1108 VDD2.n52 VDD2.n51 0.155672
R1109 VDD2.n52 VDD2.n1 0.155672
R1110 VDD2.n59 VDD2.n1 0.155672
R1111 B.n454 B.n453 585
R1112 B.n452 B.n147 585
R1113 B.n451 B.n450 585
R1114 B.n449 B.n148 585
R1115 B.n448 B.n447 585
R1116 B.n446 B.n149 585
R1117 B.n445 B.n444 585
R1118 B.n443 B.n150 585
R1119 B.n442 B.n441 585
R1120 B.n440 B.n151 585
R1121 B.n439 B.n438 585
R1122 B.n437 B.n152 585
R1123 B.n436 B.n435 585
R1124 B.n434 B.n153 585
R1125 B.n433 B.n432 585
R1126 B.n431 B.n154 585
R1127 B.n430 B.n429 585
R1128 B.n428 B.n155 585
R1129 B.n427 B.n426 585
R1130 B.n425 B.n156 585
R1131 B.n424 B.n423 585
R1132 B.n422 B.n157 585
R1133 B.n421 B.n420 585
R1134 B.n419 B.n158 585
R1135 B.n418 B.n417 585
R1136 B.n416 B.n159 585
R1137 B.n415 B.n414 585
R1138 B.n413 B.n160 585
R1139 B.n412 B.n411 585
R1140 B.n410 B.n161 585
R1141 B.n409 B.n408 585
R1142 B.n407 B.n162 585
R1143 B.n406 B.n405 585
R1144 B.n404 B.n163 585
R1145 B.n403 B.n402 585
R1146 B.n401 B.n164 585
R1147 B.n400 B.n399 585
R1148 B.n398 B.n165 585
R1149 B.n397 B.n396 585
R1150 B.n395 B.n166 585
R1151 B.n394 B.n393 585
R1152 B.n389 B.n167 585
R1153 B.n388 B.n387 585
R1154 B.n386 B.n168 585
R1155 B.n385 B.n384 585
R1156 B.n383 B.n169 585
R1157 B.n382 B.n381 585
R1158 B.n380 B.n170 585
R1159 B.n379 B.n378 585
R1160 B.n376 B.n171 585
R1161 B.n375 B.n374 585
R1162 B.n373 B.n174 585
R1163 B.n372 B.n371 585
R1164 B.n370 B.n175 585
R1165 B.n369 B.n368 585
R1166 B.n367 B.n176 585
R1167 B.n366 B.n365 585
R1168 B.n364 B.n177 585
R1169 B.n363 B.n362 585
R1170 B.n361 B.n178 585
R1171 B.n360 B.n359 585
R1172 B.n358 B.n179 585
R1173 B.n357 B.n356 585
R1174 B.n355 B.n180 585
R1175 B.n354 B.n353 585
R1176 B.n352 B.n181 585
R1177 B.n351 B.n350 585
R1178 B.n349 B.n182 585
R1179 B.n348 B.n347 585
R1180 B.n346 B.n183 585
R1181 B.n345 B.n344 585
R1182 B.n343 B.n184 585
R1183 B.n342 B.n341 585
R1184 B.n340 B.n185 585
R1185 B.n339 B.n338 585
R1186 B.n337 B.n186 585
R1187 B.n336 B.n335 585
R1188 B.n334 B.n187 585
R1189 B.n333 B.n332 585
R1190 B.n331 B.n188 585
R1191 B.n330 B.n329 585
R1192 B.n328 B.n189 585
R1193 B.n327 B.n326 585
R1194 B.n325 B.n190 585
R1195 B.n324 B.n323 585
R1196 B.n322 B.n191 585
R1197 B.n321 B.n320 585
R1198 B.n319 B.n192 585
R1199 B.n318 B.n317 585
R1200 B.n455 B.n146 585
R1201 B.n457 B.n456 585
R1202 B.n458 B.n145 585
R1203 B.n460 B.n459 585
R1204 B.n461 B.n144 585
R1205 B.n463 B.n462 585
R1206 B.n464 B.n143 585
R1207 B.n466 B.n465 585
R1208 B.n467 B.n142 585
R1209 B.n469 B.n468 585
R1210 B.n470 B.n141 585
R1211 B.n472 B.n471 585
R1212 B.n473 B.n140 585
R1213 B.n475 B.n474 585
R1214 B.n476 B.n139 585
R1215 B.n478 B.n477 585
R1216 B.n479 B.n138 585
R1217 B.n481 B.n480 585
R1218 B.n482 B.n137 585
R1219 B.n484 B.n483 585
R1220 B.n485 B.n136 585
R1221 B.n487 B.n486 585
R1222 B.n488 B.n135 585
R1223 B.n490 B.n489 585
R1224 B.n491 B.n134 585
R1225 B.n493 B.n492 585
R1226 B.n494 B.n133 585
R1227 B.n496 B.n495 585
R1228 B.n497 B.n132 585
R1229 B.n499 B.n498 585
R1230 B.n500 B.n131 585
R1231 B.n502 B.n501 585
R1232 B.n503 B.n130 585
R1233 B.n505 B.n504 585
R1234 B.n506 B.n129 585
R1235 B.n508 B.n507 585
R1236 B.n509 B.n128 585
R1237 B.n511 B.n510 585
R1238 B.n512 B.n127 585
R1239 B.n514 B.n513 585
R1240 B.n515 B.n126 585
R1241 B.n517 B.n516 585
R1242 B.n518 B.n125 585
R1243 B.n520 B.n519 585
R1244 B.n521 B.n124 585
R1245 B.n523 B.n522 585
R1246 B.n524 B.n123 585
R1247 B.n526 B.n525 585
R1248 B.n527 B.n122 585
R1249 B.n529 B.n528 585
R1250 B.n530 B.n121 585
R1251 B.n532 B.n531 585
R1252 B.n533 B.n120 585
R1253 B.n535 B.n534 585
R1254 B.n536 B.n119 585
R1255 B.n538 B.n537 585
R1256 B.n539 B.n118 585
R1257 B.n541 B.n540 585
R1258 B.n542 B.n117 585
R1259 B.n544 B.n543 585
R1260 B.n545 B.n116 585
R1261 B.n547 B.n546 585
R1262 B.n548 B.n115 585
R1263 B.n550 B.n549 585
R1264 B.n551 B.n114 585
R1265 B.n553 B.n552 585
R1266 B.n554 B.n113 585
R1267 B.n556 B.n555 585
R1268 B.n557 B.n112 585
R1269 B.n559 B.n558 585
R1270 B.n560 B.n111 585
R1271 B.n562 B.n561 585
R1272 B.n563 B.n110 585
R1273 B.n565 B.n564 585
R1274 B.n566 B.n109 585
R1275 B.n568 B.n567 585
R1276 B.n569 B.n108 585
R1277 B.n571 B.n570 585
R1278 B.n572 B.n107 585
R1279 B.n574 B.n573 585
R1280 B.n575 B.n106 585
R1281 B.n577 B.n576 585
R1282 B.n578 B.n105 585
R1283 B.n580 B.n579 585
R1284 B.n581 B.n104 585
R1285 B.n583 B.n582 585
R1286 B.n584 B.n103 585
R1287 B.n586 B.n585 585
R1288 B.n587 B.n102 585
R1289 B.n589 B.n588 585
R1290 B.n590 B.n101 585
R1291 B.n592 B.n591 585
R1292 B.n593 B.n100 585
R1293 B.n595 B.n594 585
R1294 B.n596 B.n99 585
R1295 B.n598 B.n597 585
R1296 B.n599 B.n98 585
R1297 B.n601 B.n600 585
R1298 B.n602 B.n97 585
R1299 B.n604 B.n603 585
R1300 B.n605 B.n96 585
R1301 B.n607 B.n606 585
R1302 B.n608 B.n95 585
R1303 B.n610 B.n609 585
R1304 B.n611 B.n94 585
R1305 B.n613 B.n612 585
R1306 B.n614 B.n93 585
R1307 B.n616 B.n615 585
R1308 B.n617 B.n92 585
R1309 B.n619 B.n618 585
R1310 B.n620 B.n91 585
R1311 B.n622 B.n621 585
R1312 B.n623 B.n90 585
R1313 B.n625 B.n624 585
R1314 B.n626 B.n89 585
R1315 B.n628 B.n627 585
R1316 B.n629 B.n88 585
R1317 B.n631 B.n630 585
R1318 B.n632 B.n87 585
R1319 B.n634 B.n633 585
R1320 B.n635 B.n86 585
R1321 B.n637 B.n636 585
R1322 B.n638 B.n85 585
R1323 B.n640 B.n639 585
R1324 B.n641 B.n84 585
R1325 B.n643 B.n642 585
R1326 B.n644 B.n83 585
R1327 B.n646 B.n645 585
R1328 B.n781 B.n780 585
R1329 B.n779 B.n34 585
R1330 B.n778 B.n777 585
R1331 B.n776 B.n35 585
R1332 B.n775 B.n774 585
R1333 B.n773 B.n36 585
R1334 B.n772 B.n771 585
R1335 B.n770 B.n37 585
R1336 B.n769 B.n768 585
R1337 B.n767 B.n38 585
R1338 B.n766 B.n765 585
R1339 B.n764 B.n39 585
R1340 B.n763 B.n762 585
R1341 B.n761 B.n40 585
R1342 B.n760 B.n759 585
R1343 B.n758 B.n41 585
R1344 B.n757 B.n756 585
R1345 B.n755 B.n42 585
R1346 B.n754 B.n753 585
R1347 B.n752 B.n43 585
R1348 B.n751 B.n750 585
R1349 B.n749 B.n44 585
R1350 B.n748 B.n747 585
R1351 B.n746 B.n45 585
R1352 B.n745 B.n744 585
R1353 B.n743 B.n46 585
R1354 B.n742 B.n741 585
R1355 B.n740 B.n47 585
R1356 B.n739 B.n738 585
R1357 B.n737 B.n48 585
R1358 B.n736 B.n735 585
R1359 B.n734 B.n49 585
R1360 B.n733 B.n732 585
R1361 B.n731 B.n50 585
R1362 B.n730 B.n729 585
R1363 B.n728 B.n51 585
R1364 B.n727 B.n726 585
R1365 B.n725 B.n52 585
R1366 B.n724 B.n723 585
R1367 B.n722 B.n53 585
R1368 B.n720 B.n719 585
R1369 B.n718 B.n56 585
R1370 B.n717 B.n716 585
R1371 B.n715 B.n57 585
R1372 B.n714 B.n713 585
R1373 B.n712 B.n58 585
R1374 B.n711 B.n710 585
R1375 B.n709 B.n59 585
R1376 B.n708 B.n707 585
R1377 B.n706 B.n705 585
R1378 B.n704 B.n63 585
R1379 B.n703 B.n702 585
R1380 B.n701 B.n64 585
R1381 B.n700 B.n699 585
R1382 B.n698 B.n65 585
R1383 B.n697 B.n696 585
R1384 B.n695 B.n66 585
R1385 B.n694 B.n693 585
R1386 B.n692 B.n67 585
R1387 B.n691 B.n690 585
R1388 B.n689 B.n68 585
R1389 B.n688 B.n687 585
R1390 B.n686 B.n69 585
R1391 B.n685 B.n684 585
R1392 B.n683 B.n70 585
R1393 B.n682 B.n681 585
R1394 B.n680 B.n71 585
R1395 B.n679 B.n678 585
R1396 B.n677 B.n72 585
R1397 B.n676 B.n675 585
R1398 B.n674 B.n73 585
R1399 B.n673 B.n672 585
R1400 B.n671 B.n74 585
R1401 B.n670 B.n669 585
R1402 B.n668 B.n75 585
R1403 B.n667 B.n666 585
R1404 B.n665 B.n76 585
R1405 B.n664 B.n663 585
R1406 B.n662 B.n77 585
R1407 B.n661 B.n660 585
R1408 B.n659 B.n78 585
R1409 B.n658 B.n657 585
R1410 B.n656 B.n79 585
R1411 B.n655 B.n654 585
R1412 B.n653 B.n80 585
R1413 B.n652 B.n651 585
R1414 B.n650 B.n81 585
R1415 B.n649 B.n648 585
R1416 B.n647 B.n82 585
R1417 B.n782 B.n33 585
R1418 B.n784 B.n783 585
R1419 B.n785 B.n32 585
R1420 B.n787 B.n786 585
R1421 B.n788 B.n31 585
R1422 B.n790 B.n789 585
R1423 B.n791 B.n30 585
R1424 B.n793 B.n792 585
R1425 B.n794 B.n29 585
R1426 B.n796 B.n795 585
R1427 B.n797 B.n28 585
R1428 B.n799 B.n798 585
R1429 B.n800 B.n27 585
R1430 B.n802 B.n801 585
R1431 B.n803 B.n26 585
R1432 B.n805 B.n804 585
R1433 B.n806 B.n25 585
R1434 B.n808 B.n807 585
R1435 B.n809 B.n24 585
R1436 B.n811 B.n810 585
R1437 B.n812 B.n23 585
R1438 B.n814 B.n813 585
R1439 B.n815 B.n22 585
R1440 B.n817 B.n816 585
R1441 B.n818 B.n21 585
R1442 B.n820 B.n819 585
R1443 B.n821 B.n20 585
R1444 B.n823 B.n822 585
R1445 B.n824 B.n19 585
R1446 B.n826 B.n825 585
R1447 B.n827 B.n18 585
R1448 B.n829 B.n828 585
R1449 B.n830 B.n17 585
R1450 B.n832 B.n831 585
R1451 B.n833 B.n16 585
R1452 B.n835 B.n834 585
R1453 B.n836 B.n15 585
R1454 B.n838 B.n837 585
R1455 B.n839 B.n14 585
R1456 B.n841 B.n840 585
R1457 B.n842 B.n13 585
R1458 B.n844 B.n843 585
R1459 B.n845 B.n12 585
R1460 B.n847 B.n846 585
R1461 B.n848 B.n11 585
R1462 B.n850 B.n849 585
R1463 B.n851 B.n10 585
R1464 B.n853 B.n852 585
R1465 B.n854 B.n9 585
R1466 B.n856 B.n855 585
R1467 B.n857 B.n8 585
R1468 B.n859 B.n858 585
R1469 B.n860 B.n7 585
R1470 B.n862 B.n861 585
R1471 B.n863 B.n6 585
R1472 B.n865 B.n864 585
R1473 B.n866 B.n5 585
R1474 B.n868 B.n867 585
R1475 B.n869 B.n4 585
R1476 B.n871 B.n870 585
R1477 B.n872 B.n3 585
R1478 B.n874 B.n873 585
R1479 B.n875 B.n0 585
R1480 B.n2 B.n1 585
R1481 B.n225 B.n224 585
R1482 B.n226 B.n223 585
R1483 B.n228 B.n227 585
R1484 B.n229 B.n222 585
R1485 B.n231 B.n230 585
R1486 B.n232 B.n221 585
R1487 B.n234 B.n233 585
R1488 B.n235 B.n220 585
R1489 B.n237 B.n236 585
R1490 B.n238 B.n219 585
R1491 B.n240 B.n239 585
R1492 B.n241 B.n218 585
R1493 B.n243 B.n242 585
R1494 B.n244 B.n217 585
R1495 B.n246 B.n245 585
R1496 B.n247 B.n216 585
R1497 B.n249 B.n248 585
R1498 B.n250 B.n215 585
R1499 B.n252 B.n251 585
R1500 B.n253 B.n214 585
R1501 B.n255 B.n254 585
R1502 B.n256 B.n213 585
R1503 B.n258 B.n257 585
R1504 B.n259 B.n212 585
R1505 B.n261 B.n260 585
R1506 B.n262 B.n211 585
R1507 B.n264 B.n263 585
R1508 B.n265 B.n210 585
R1509 B.n267 B.n266 585
R1510 B.n268 B.n209 585
R1511 B.n270 B.n269 585
R1512 B.n271 B.n208 585
R1513 B.n273 B.n272 585
R1514 B.n274 B.n207 585
R1515 B.n276 B.n275 585
R1516 B.n277 B.n206 585
R1517 B.n279 B.n278 585
R1518 B.n280 B.n205 585
R1519 B.n282 B.n281 585
R1520 B.n283 B.n204 585
R1521 B.n285 B.n284 585
R1522 B.n286 B.n203 585
R1523 B.n288 B.n287 585
R1524 B.n289 B.n202 585
R1525 B.n291 B.n290 585
R1526 B.n292 B.n201 585
R1527 B.n294 B.n293 585
R1528 B.n295 B.n200 585
R1529 B.n297 B.n296 585
R1530 B.n298 B.n199 585
R1531 B.n300 B.n299 585
R1532 B.n301 B.n198 585
R1533 B.n303 B.n302 585
R1534 B.n304 B.n197 585
R1535 B.n306 B.n305 585
R1536 B.n307 B.n196 585
R1537 B.n309 B.n308 585
R1538 B.n310 B.n195 585
R1539 B.n312 B.n311 585
R1540 B.n313 B.n194 585
R1541 B.n315 B.n314 585
R1542 B.n316 B.n193 585
R1543 B.n318 B.n193 540.549
R1544 B.n455 B.n454 540.549
R1545 B.n647 B.n646 540.549
R1546 B.n780 B.n33 540.549
R1547 B.n390 B.t4 426.315
R1548 B.n60 B.t2 426.315
R1549 B.n172 B.t10 426.315
R1550 B.n54 B.t8 426.315
R1551 B.n391 B.t5 365.418
R1552 B.n61 B.t1 365.418
R1553 B.n173 B.t11 365.418
R1554 B.n55 B.t7 365.418
R1555 B.n172 B.t9 306.373
R1556 B.n390 B.t3 306.373
R1557 B.n60 B.t0 306.373
R1558 B.n54 B.t6 306.373
R1559 B.n877 B.n876 256.663
R1560 B.n876 B.n875 235.042
R1561 B.n876 B.n2 235.042
R1562 B.n319 B.n318 163.367
R1563 B.n320 B.n319 163.367
R1564 B.n320 B.n191 163.367
R1565 B.n324 B.n191 163.367
R1566 B.n325 B.n324 163.367
R1567 B.n326 B.n325 163.367
R1568 B.n326 B.n189 163.367
R1569 B.n330 B.n189 163.367
R1570 B.n331 B.n330 163.367
R1571 B.n332 B.n331 163.367
R1572 B.n332 B.n187 163.367
R1573 B.n336 B.n187 163.367
R1574 B.n337 B.n336 163.367
R1575 B.n338 B.n337 163.367
R1576 B.n338 B.n185 163.367
R1577 B.n342 B.n185 163.367
R1578 B.n343 B.n342 163.367
R1579 B.n344 B.n343 163.367
R1580 B.n344 B.n183 163.367
R1581 B.n348 B.n183 163.367
R1582 B.n349 B.n348 163.367
R1583 B.n350 B.n349 163.367
R1584 B.n350 B.n181 163.367
R1585 B.n354 B.n181 163.367
R1586 B.n355 B.n354 163.367
R1587 B.n356 B.n355 163.367
R1588 B.n356 B.n179 163.367
R1589 B.n360 B.n179 163.367
R1590 B.n361 B.n360 163.367
R1591 B.n362 B.n361 163.367
R1592 B.n362 B.n177 163.367
R1593 B.n366 B.n177 163.367
R1594 B.n367 B.n366 163.367
R1595 B.n368 B.n367 163.367
R1596 B.n368 B.n175 163.367
R1597 B.n372 B.n175 163.367
R1598 B.n373 B.n372 163.367
R1599 B.n374 B.n373 163.367
R1600 B.n374 B.n171 163.367
R1601 B.n379 B.n171 163.367
R1602 B.n380 B.n379 163.367
R1603 B.n381 B.n380 163.367
R1604 B.n381 B.n169 163.367
R1605 B.n385 B.n169 163.367
R1606 B.n386 B.n385 163.367
R1607 B.n387 B.n386 163.367
R1608 B.n387 B.n167 163.367
R1609 B.n394 B.n167 163.367
R1610 B.n395 B.n394 163.367
R1611 B.n396 B.n395 163.367
R1612 B.n396 B.n165 163.367
R1613 B.n400 B.n165 163.367
R1614 B.n401 B.n400 163.367
R1615 B.n402 B.n401 163.367
R1616 B.n402 B.n163 163.367
R1617 B.n406 B.n163 163.367
R1618 B.n407 B.n406 163.367
R1619 B.n408 B.n407 163.367
R1620 B.n408 B.n161 163.367
R1621 B.n412 B.n161 163.367
R1622 B.n413 B.n412 163.367
R1623 B.n414 B.n413 163.367
R1624 B.n414 B.n159 163.367
R1625 B.n418 B.n159 163.367
R1626 B.n419 B.n418 163.367
R1627 B.n420 B.n419 163.367
R1628 B.n420 B.n157 163.367
R1629 B.n424 B.n157 163.367
R1630 B.n425 B.n424 163.367
R1631 B.n426 B.n425 163.367
R1632 B.n426 B.n155 163.367
R1633 B.n430 B.n155 163.367
R1634 B.n431 B.n430 163.367
R1635 B.n432 B.n431 163.367
R1636 B.n432 B.n153 163.367
R1637 B.n436 B.n153 163.367
R1638 B.n437 B.n436 163.367
R1639 B.n438 B.n437 163.367
R1640 B.n438 B.n151 163.367
R1641 B.n442 B.n151 163.367
R1642 B.n443 B.n442 163.367
R1643 B.n444 B.n443 163.367
R1644 B.n444 B.n149 163.367
R1645 B.n448 B.n149 163.367
R1646 B.n449 B.n448 163.367
R1647 B.n450 B.n449 163.367
R1648 B.n450 B.n147 163.367
R1649 B.n454 B.n147 163.367
R1650 B.n646 B.n83 163.367
R1651 B.n642 B.n83 163.367
R1652 B.n642 B.n641 163.367
R1653 B.n641 B.n640 163.367
R1654 B.n640 B.n85 163.367
R1655 B.n636 B.n85 163.367
R1656 B.n636 B.n635 163.367
R1657 B.n635 B.n634 163.367
R1658 B.n634 B.n87 163.367
R1659 B.n630 B.n87 163.367
R1660 B.n630 B.n629 163.367
R1661 B.n629 B.n628 163.367
R1662 B.n628 B.n89 163.367
R1663 B.n624 B.n89 163.367
R1664 B.n624 B.n623 163.367
R1665 B.n623 B.n622 163.367
R1666 B.n622 B.n91 163.367
R1667 B.n618 B.n91 163.367
R1668 B.n618 B.n617 163.367
R1669 B.n617 B.n616 163.367
R1670 B.n616 B.n93 163.367
R1671 B.n612 B.n93 163.367
R1672 B.n612 B.n611 163.367
R1673 B.n611 B.n610 163.367
R1674 B.n610 B.n95 163.367
R1675 B.n606 B.n95 163.367
R1676 B.n606 B.n605 163.367
R1677 B.n605 B.n604 163.367
R1678 B.n604 B.n97 163.367
R1679 B.n600 B.n97 163.367
R1680 B.n600 B.n599 163.367
R1681 B.n599 B.n598 163.367
R1682 B.n598 B.n99 163.367
R1683 B.n594 B.n99 163.367
R1684 B.n594 B.n593 163.367
R1685 B.n593 B.n592 163.367
R1686 B.n592 B.n101 163.367
R1687 B.n588 B.n101 163.367
R1688 B.n588 B.n587 163.367
R1689 B.n587 B.n586 163.367
R1690 B.n586 B.n103 163.367
R1691 B.n582 B.n103 163.367
R1692 B.n582 B.n581 163.367
R1693 B.n581 B.n580 163.367
R1694 B.n580 B.n105 163.367
R1695 B.n576 B.n105 163.367
R1696 B.n576 B.n575 163.367
R1697 B.n575 B.n574 163.367
R1698 B.n574 B.n107 163.367
R1699 B.n570 B.n107 163.367
R1700 B.n570 B.n569 163.367
R1701 B.n569 B.n568 163.367
R1702 B.n568 B.n109 163.367
R1703 B.n564 B.n109 163.367
R1704 B.n564 B.n563 163.367
R1705 B.n563 B.n562 163.367
R1706 B.n562 B.n111 163.367
R1707 B.n558 B.n111 163.367
R1708 B.n558 B.n557 163.367
R1709 B.n557 B.n556 163.367
R1710 B.n556 B.n113 163.367
R1711 B.n552 B.n113 163.367
R1712 B.n552 B.n551 163.367
R1713 B.n551 B.n550 163.367
R1714 B.n550 B.n115 163.367
R1715 B.n546 B.n115 163.367
R1716 B.n546 B.n545 163.367
R1717 B.n545 B.n544 163.367
R1718 B.n544 B.n117 163.367
R1719 B.n540 B.n117 163.367
R1720 B.n540 B.n539 163.367
R1721 B.n539 B.n538 163.367
R1722 B.n538 B.n119 163.367
R1723 B.n534 B.n119 163.367
R1724 B.n534 B.n533 163.367
R1725 B.n533 B.n532 163.367
R1726 B.n532 B.n121 163.367
R1727 B.n528 B.n121 163.367
R1728 B.n528 B.n527 163.367
R1729 B.n527 B.n526 163.367
R1730 B.n526 B.n123 163.367
R1731 B.n522 B.n123 163.367
R1732 B.n522 B.n521 163.367
R1733 B.n521 B.n520 163.367
R1734 B.n520 B.n125 163.367
R1735 B.n516 B.n125 163.367
R1736 B.n516 B.n515 163.367
R1737 B.n515 B.n514 163.367
R1738 B.n514 B.n127 163.367
R1739 B.n510 B.n127 163.367
R1740 B.n510 B.n509 163.367
R1741 B.n509 B.n508 163.367
R1742 B.n508 B.n129 163.367
R1743 B.n504 B.n129 163.367
R1744 B.n504 B.n503 163.367
R1745 B.n503 B.n502 163.367
R1746 B.n502 B.n131 163.367
R1747 B.n498 B.n131 163.367
R1748 B.n498 B.n497 163.367
R1749 B.n497 B.n496 163.367
R1750 B.n496 B.n133 163.367
R1751 B.n492 B.n133 163.367
R1752 B.n492 B.n491 163.367
R1753 B.n491 B.n490 163.367
R1754 B.n490 B.n135 163.367
R1755 B.n486 B.n135 163.367
R1756 B.n486 B.n485 163.367
R1757 B.n485 B.n484 163.367
R1758 B.n484 B.n137 163.367
R1759 B.n480 B.n137 163.367
R1760 B.n480 B.n479 163.367
R1761 B.n479 B.n478 163.367
R1762 B.n478 B.n139 163.367
R1763 B.n474 B.n139 163.367
R1764 B.n474 B.n473 163.367
R1765 B.n473 B.n472 163.367
R1766 B.n472 B.n141 163.367
R1767 B.n468 B.n141 163.367
R1768 B.n468 B.n467 163.367
R1769 B.n467 B.n466 163.367
R1770 B.n466 B.n143 163.367
R1771 B.n462 B.n143 163.367
R1772 B.n462 B.n461 163.367
R1773 B.n461 B.n460 163.367
R1774 B.n460 B.n145 163.367
R1775 B.n456 B.n145 163.367
R1776 B.n456 B.n455 163.367
R1777 B.n780 B.n779 163.367
R1778 B.n779 B.n778 163.367
R1779 B.n778 B.n35 163.367
R1780 B.n774 B.n35 163.367
R1781 B.n774 B.n773 163.367
R1782 B.n773 B.n772 163.367
R1783 B.n772 B.n37 163.367
R1784 B.n768 B.n37 163.367
R1785 B.n768 B.n767 163.367
R1786 B.n767 B.n766 163.367
R1787 B.n766 B.n39 163.367
R1788 B.n762 B.n39 163.367
R1789 B.n762 B.n761 163.367
R1790 B.n761 B.n760 163.367
R1791 B.n760 B.n41 163.367
R1792 B.n756 B.n41 163.367
R1793 B.n756 B.n755 163.367
R1794 B.n755 B.n754 163.367
R1795 B.n754 B.n43 163.367
R1796 B.n750 B.n43 163.367
R1797 B.n750 B.n749 163.367
R1798 B.n749 B.n748 163.367
R1799 B.n748 B.n45 163.367
R1800 B.n744 B.n45 163.367
R1801 B.n744 B.n743 163.367
R1802 B.n743 B.n742 163.367
R1803 B.n742 B.n47 163.367
R1804 B.n738 B.n47 163.367
R1805 B.n738 B.n737 163.367
R1806 B.n737 B.n736 163.367
R1807 B.n736 B.n49 163.367
R1808 B.n732 B.n49 163.367
R1809 B.n732 B.n731 163.367
R1810 B.n731 B.n730 163.367
R1811 B.n730 B.n51 163.367
R1812 B.n726 B.n51 163.367
R1813 B.n726 B.n725 163.367
R1814 B.n725 B.n724 163.367
R1815 B.n724 B.n53 163.367
R1816 B.n719 B.n53 163.367
R1817 B.n719 B.n718 163.367
R1818 B.n718 B.n717 163.367
R1819 B.n717 B.n57 163.367
R1820 B.n713 B.n57 163.367
R1821 B.n713 B.n712 163.367
R1822 B.n712 B.n711 163.367
R1823 B.n711 B.n59 163.367
R1824 B.n707 B.n59 163.367
R1825 B.n707 B.n706 163.367
R1826 B.n706 B.n63 163.367
R1827 B.n702 B.n63 163.367
R1828 B.n702 B.n701 163.367
R1829 B.n701 B.n700 163.367
R1830 B.n700 B.n65 163.367
R1831 B.n696 B.n65 163.367
R1832 B.n696 B.n695 163.367
R1833 B.n695 B.n694 163.367
R1834 B.n694 B.n67 163.367
R1835 B.n690 B.n67 163.367
R1836 B.n690 B.n689 163.367
R1837 B.n689 B.n688 163.367
R1838 B.n688 B.n69 163.367
R1839 B.n684 B.n69 163.367
R1840 B.n684 B.n683 163.367
R1841 B.n683 B.n682 163.367
R1842 B.n682 B.n71 163.367
R1843 B.n678 B.n71 163.367
R1844 B.n678 B.n677 163.367
R1845 B.n677 B.n676 163.367
R1846 B.n676 B.n73 163.367
R1847 B.n672 B.n73 163.367
R1848 B.n672 B.n671 163.367
R1849 B.n671 B.n670 163.367
R1850 B.n670 B.n75 163.367
R1851 B.n666 B.n75 163.367
R1852 B.n666 B.n665 163.367
R1853 B.n665 B.n664 163.367
R1854 B.n664 B.n77 163.367
R1855 B.n660 B.n77 163.367
R1856 B.n660 B.n659 163.367
R1857 B.n659 B.n658 163.367
R1858 B.n658 B.n79 163.367
R1859 B.n654 B.n79 163.367
R1860 B.n654 B.n653 163.367
R1861 B.n653 B.n652 163.367
R1862 B.n652 B.n81 163.367
R1863 B.n648 B.n81 163.367
R1864 B.n648 B.n647 163.367
R1865 B.n784 B.n33 163.367
R1866 B.n785 B.n784 163.367
R1867 B.n786 B.n785 163.367
R1868 B.n786 B.n31 163.367
R1869 B.n790 B.n31 163.367
R1870 B.n791 B.n790 163.367
R1871 B.n792 B.n791 163.367
R1872 B.n792 B.n29 163.367
R1873 B.n796 B.n29 163.367
R1874 B.n797 B.n796 163.367
R1875 B.n798 B.n797 163.367
R1876 B.n798 B.n27 163.367
R1877 B.n802 B.n27 163.367
R1878 B.n803 B.n802 163.367
R1879 B.n804 B.n803 163.367
R1880 B.n804 B.n25 163.367
R1881 B.n808 B.n25 163.367
R1882 B.n809 B.n808 163.367
R1883 B.n810 B.n809 163.367
R1884 B.n810 B.n23 163.367
R1885 B.n814 B.n23 163.367
R1886 B.n815 B.n814 163.367
R1887 B.n816 B.n815 163.367
R1888 B.n816 B.n21 163.367
R1889 B.n820 B.n21 163.367
R1890 B.n821 B.n820 163.367
R1891 B.n822 B.n821 163.367
R1892 B.n822 B.n19 163.367
R1893 B.n826 B.n19 163.367
R1894 B.n827 B.n826 163.367
R1895 B.n828 B.n827 163.367
R1896 B.n828 B.n17 163.367
R1897 B.n832 B.n17 163.367
R1898 B.n833 B.n832 163.367
R1899 B.n834 B.n833 163.367
R1900 B.n834 B.n15 163.367
R1901 B.n838 B.n15 163.367
R1902 B.n839 B.n838 163.367
R1903 B.n840 B.n839 163.367
R1904 B.n840 B.n13 163.367
R1905 B.n844 B.n13 163.367
R1906 B.n845 B.n844 163.367
R1907 B.n846 B.n845 163.367
R1908 B.n846 B.n11 163.367
R1909 B.n850 B.n11 163.367
R1910 B.n851 B.n850 163.367
R1911 B.n852 B.n851 163.367
R1912 B.n852 B.n9 163.367
R1913 B.n856 B.n9 163.367
R1914 B.n857 B.n856 163.367
R1915 B.n858 B.n857 163.367
R1916 B.n858 B.n7 163.367
R1917 B.n862 B.n7 163.367
R1918 B.n863 B.n862 163.367
R1919 B.n864 B.n863 163.367
R1920 B.n864 B.n5 163.367
R1921 B.n868 B.n5 163.367
R1922 B.n869 B.n868 163.367
R1923 B.n870 B.n869 163.367
R1924 B.n870 B.n3 163.367
R1925 B.n874 B.n3 163.367
R1926 B.n875 B.n874 163.367
R1927 B.n224 B.n2 163.367
R1928 B.n224 B.n223 163.367
R1929 B.n228 B.n223 163.367
R1930 B.n229 B.n228 163.367
R1931 B.n230 B.n229 163.367
R1932 B.n230 B.n221 163.367
R1933 B.n234 B.n221 163.367
R1934 B.n235 B.n234 163.367
R1935 B.n236 B.n235 163.367
R1936 B.n236 B.n219 163.367
R1937 B.n240 B.n219 163.367
R1938 B.n241 B.n240 163.367
R1939 B.n242 B.n241 163.367
R1940 B.n242 B.n217 163.367
R1941 B.n246 B.n217 163.367
R1942 B.n247 B.n246 163.367
R1943 B.n248 B.n247 163.367
R1944 B.n248 B.n215 163.367
R1945 B.n252 B.n215 163.367
R1946 B.n253 B.n252 163.367
R1947 B.n254 B.n253 163.367
R1948 B.n254 B.n213 163.367
R1949 B.n258 B.n213 163.367
R1950 B.n259 B.n258 163.367
R1951 B.n260 B.n259 163.367
R1952 B.n260 B.n211 163.367
R1953 B.n264 B.n211 163.367
R1954 B.n265 B.n264 163.367
R1955 B.n266 B.n265 163.367
R1956 B.n266 B.n209 163.367
R1957 B.n270 B.n209 163.367
R1958 B.n271 B.n270 163.367
R1959 B.n272 B.n271 163.367
R1960 B.n272 B.n207 163.367
R1961 B.n276 B.n207 163.367
R1962 B.n277 B.n276 163.367
R1963 B.n278 B.n277 163.367
R1964 B.n278 B.n205 163.367
R1965 B.n282 B.n205 163.367
R1966 B.n283 B.n282 163.367
R1967 B.n284 B.n283 163.367
R1968 B.n284 B.n203 163.367
R1969 B.n288 B.n203 163.367
R1970 B.n289 B.n288 163.367
R1971 B.n290 B.n289 163.367
R1972 B.n290 B.n201 163.367
R1973 B.n294 B.n201 163.367
R1974 B.n295 B.n294 163.367
R1975 B.n296 B.n295 163.367
R1976 B.n296 B.n199 163.367
R1977 B.n300 B.n199 163.367
R1978 B.n301 B.n300 163.367
R1979 B.n302 B.n301 163.367
R1980 B.n302 B.n197 163.367
R1981 B.n306 B.n197 163.367
R1982 B.n307 B.n306 163.367
R1983 B.n308 B.n307 163.367
R1984 B.n308 B.n195 163.367
R1985 B.n312 B.n195 163.367
R1986 B.n313 B.n312 163.367
R1987 B.n314 B.n313 163.367
R1988 B.n314 B.n193 163.367
R1989 B.n173 B.n172 60.8975
R1990 B.n391 B.n390 60.8975
R1991 B.n61 B.n60 60.8975
R1992 B.n55 B.n54 60.8975
R1993 B.n377 B.n173 59.5399
R1994 B.n392 B.n391 59.5399
R1995 B.n62 B.n61 59.5399
R1996 B.n721 B.n55 59.5399
R1997 B.n782 B.n781 35.1225
R1998 B.n645 B.n82 35.1225
R1999 B.n453 B.n146 35.1225
R2000 B.n317 B.n316 35.1225
R2001 B B.n877 18.0485
R2002 B.n783 B.n782 10.6151
R2003 B.n783 B.n32 10.6151
R2004 B.n787 B.n32 10.6151
R2005 B.n788 B.n787 10.6151
R2006 B.n789 B.n788 10.6151
R2007 B.n789 B.n30 10.6151
R2008 B.n793 B.n30 10.6151
R2009 B.n794 B.n793 10.6151
R2010 B.n795 B.n794 10.6151
R2011 B.n795 B.n28 10.6151
R2012 B.n799 B.n28 10.6151
R2013 B.n800 B.n799 10.6151
R2014 B.n801 B.n800 10.6151
R2015 B.n801 B.n26 10.6151
R2016 B.n805 B.n26 10.6151
R2017 B.n806 B.n805 10.6151
R2018 B.n807 B.n806 10.6151
R2019 B.n807 B.n24 10.6151
R2020 B.n811 B.n24 10.6151
R2021 B.n812 B.n811 10.6151
R2022 B.n813 B.n812 10.6151
R2023 B.n813 B.n22 10.6151
R2024 B.n817 B.n22 10.6151
R2025 B.n818 B.n817 10.6151
R2026 B.n819 B.n818 10.6151
R2027 B.n819 B.n20 10.6151
R2028 B.n823 B.n20 10.6151
R2029 B.n824 B.n823 10.6151
R2030 B.n825 B.n824 10.6151
R2031 B.n825 B.n18 10.6151
R2032 B.n829 B.n18 10.6151
R2033 B.n830 B.n829 10.6151
R2034 B.n831 B.n830 10.6151
R2035 B.n831 B.n16 10.6151
R2036 B.n835 B.n16 10.6151
R2037 B.n836 B.n835 10.6151
R2038 B.n837 B.n836 10.6151
R2039 B.n837 B.n14 10.6151
R2040 B.n841 B.n14 10.6151
R2041 B.n842 B.n841 10.6151
R2042 B.n843 B.n842 10.6151
R2043 B.n843 B.n12 10.6151
R2044 B.n847 B.n12 10.6151
R2045 B.n848 B.n847 10.6151
R2046 B.n849 B.n848 10.6151
R2047 B.n849 B.n10 10.6151
R2048 B.n853 B.n10 10.6151
R2049 B.n854 B.n853 10.6151
R2050 B.n855 B.n854 10.6151
R2051 B.n855 B.n8 10.6151
R2052 B.n859 B.n8 10.6151
R2053 B.n860 B.n859 10.6151
R2054 B.n861 B.n860 10.6151
R2055 B.n861 B.n6 10.6151
R2056 B.n865 B.n6 10.6151
R2057 B.n866 B.n865 10.6151
R2058 B.n867 B.n866 10.6151
R2059 B.n867 B.n4 10.6151
R2060 B.n871 B.n4 10.6151
R2061 B.n872 B.n871 10.6151
R2062 B.n873 B.n872 10.6151
R2063 B.n873 B.n0 10.6151
R2064 B.n781 B.n34 10.6151
R2065 B.n777 B.n34 10.6151
R2066 B.n777 B.n776 10.6151
R2067 B.n776 B.n775 10.6151
R2068 B.n775 B.n36 10.6151
R2069 B.n771 B.n36 10.6151
R2070 B.n771 B.n770 10.6151
R2071 B.n770 B.n769 10.6151
R2072 B.n769 B.n38 10.6151
R2073 B.n765 B.n38 10.6151
R2074 B.n765 B.n764 10.6151
R2075 B.n764 B.n763 10.6151
R2076 B.n763 B.n40 10.6151
R2077 B.n759 B.n40 10.6151
R2078 B.n759 B.n758 10.6151
R2079 B.n758 B.n757 10.6151
R2080 B.n757 B.n42 10.6151
R2081 B.n753 B.n42 10.6151
R2082 B.n753 B.n752 10.6151
R2083 B.n752 B.n751 10.6151
R2084 B.n751 B.n44 10.6151
R2085 B.n747 B.n44 10.6151
R2086 B.n747 B.n746 10.6151
R2087 B.n746 B.n745 10.6151
R2088 B.n745 B.n46 10.6151
R2089 B.n741 B.n46 10.6151
R2090 B.n741 B.n740 10.6151
R2091 B.n740 B.n739 10.6151
R2092 B.n739 B.n48 10.6151
R2093 B.n735 B.n48 10.6151
R2094 B.n735 B.n734 10.6151
R2095 B.n734 B.n733 10.6151
R2096 B.n733 B.n50 10.6151
R2097 B.n729 B.n50 10.6151
R2098 B.n729 B.n728 10.6151
R2099 B.n728 B.n727 10.6151
R2100 B.n727 B.n52 10.6151
R2101 B.n723 B.n52 10.6151
R2102 B.n723 B.n722 10.6151
R2103 B.n720 B.n56 10.6151
R2104 B.n716 B.n56 10.6151
R2105 B.n716 B.n715 10.6151
R2106 B.n715 B.n714 10.6151
R2107 B.n714 B.n58 10.6151
R2108 B.n710 B.n58 10.6151
R2109 B.n710 B.n709 10.6151
R2110 B.n709 B.n708 10.6151
R2111 B.n705 B.n704 10.6151
R2112 B.n704 B.n703 10.6151
R2113 B.n703 B.n64 10.6151
R2114 B.n699 B.n64 10.6151
R2115 B.n699 B.n698 10.6151
R2116 B.n698 B.n697 10.6151
R2117 B.n697 B.n66 10.6151
R2118 B.n693 B.n66 10.6151
R2119 B.n693 B.n692 10.6151
R2120 B.n692 B.n691 10.6151
R2121 B.n691 B.n68 10.6151
R2122 B.n687 B.n68 10.6151
R2123 B.n687 B.n686 10.6151
R2124 B.n686 B.n685 10.6151
R2125 B.n685 B.n70 10.6151
R2126 B.n681 B.n70 10.6151
R2127 B.n681 B.n680 10.6151
R2128 B.n680 B.n679 10.6151
R2129 B.n679 B.n72 10.6151
R2130 B.n675 B.n72 10.6151
R2131 B.n675 B.n674 10.6151
R2132 B.n674 B.n673 10.6151
R2133 B.n673 B.n74 10.6151
R2134 B.n669 B.n74 10.6151
R2135 B.n669 B.n668 10.6151
R2136 B.n668 B.n667 10.6151
R2137 B.n667 B.n76 10.6151
R2138 B.n663 B.n76 10.6151
R2139 B.n663 B.n662 10.6151
R2140 B.n662 B.n661 10.6151
R2141 B.n661 B.n78 10.6151
R2142 B.n657 B.n78 10.6151
R2143 B.n657 B.n656 10.6151
R2144 B.n656 B.n655 10.6151
R2145 B.n655 B.n80 10.6151
R2146 B.n651 B.n80 10.6151
R2147 B.n651 B.n650 10.6151
R2148 B.n650 B.n649 10.6151
R2149 B.n649 B.n82 10.6151
R2150 B.n645 B.n644 10.6151
R2151 B.n644 B.n643 10.6151
R2152 B.n643 B.n84 10.6151
R2153 B.n639 B.n84 10.6151
R2154 B.n639 B.n638 10.6151
R2155 B.n638 B.n637 10.6151
R2156 B.n637 B.n86 10.6151
R2157 B.n633 B.n86 10.6151
R2158 B.n633 B.n632 10.6151
R2159 B.n632 B.n631 10.6151
R2160 B.n631 B.n88 10.6151
R2161 B.n627 B.n88 10.6151
R2162 B.n627 B.n626 10.6151
R2163 B.n626 B.n625 10.6151
R2164 B.n625 B.n90 10.6151
R2165 B.n621 B.n90 10.6151
R2166 B.n621 B.n620 10.6151
R2167 B.n620 B.n619 10.6151
R2168 B.n619 B.n92 10.6151
R2169 B.n615 B.n92 10.6151
R2170 B.n615 B.n614 10.6151
R2171 B.n614 B.n613 10.6151
R2172 B.n613 B.n94 10.6151
R2173 B.n609 B.n94 10.6151
R2174 B.n609 B.n608 10.6151
R2175 B.n608 B.n607 10.6151
R2176 B.n607 B.n96 10.6151
R2177 B.n603 B.n96 10.6151
R2178 B.n603 B.n602 10.6151
R2179 B.n602 B.n601 10.6151
R2180 B.n601 B.n98 10.6151
R2181 B.n597 B.n98 10.6151
R2182 B.n597 B.n596 10.6151
R2183 B.n596 B.n595 10.6151
R2184 B.n595 B.n100 10.6151
R2185 B.n591 B.n100 10.6151
R2186 B.n591 B.n590 10.6151
R2187 B.n590 B.n589 10.6151
R2188 B.n589 B.n102 10.6151
R2189 B.n585 B.n102 10.6151
R2190 B.n585 B.n584 10.6151
R2191 B.n584 B.n583 10.6151
R2192 B.n583 B.n104 10.6151
R2193 B.n579 B.n104 10.6151
R2194 B.n579 B.n578 10.6151
R2195 B.n578 B.n577 10.6151
R2196 B.n577 B.n106 10.6151
R2197 B.n573 B.n106 10.6151
R2198 B.n573 B.n572 10.6151
R2199 B.n572 B.n571 10.6151
R2200 B.n571 B.n108 10.6151
R2201 B.n567 B.n108 10.6151
R2202 B.n567 B.n566 10.6151
R2203 B.n566 B.n565 10.6151
R2204 B.n565 B.n110 10.6151
R2205 B.n561 B.n110 10.6151
R2206 B.n561 B.n560 10.6151
R2207 B.n560 B.n559 10.6151
R2208 B.n559 B.n112 10.6151
R2209 B.n555 B.n112 10.6151
R2210 B.n555 B.n554 10.6151
R2211 B.n554 B.n553 10.6151
R2212 B.n553 B.n114 10.6151
R2213 B.n549 B.n114 10.6151
R2214 B.n549 B.n548 10.6151
R2215 B.n548 B.n547 10.6151
R2216 B.n547 B.n116 10.6151
R2217 B.n543 B.n116 10.6151
R2218 B.n543 B.n542 10.6151
R2219 B.n542 B.n541 10.6151
R2220 B.n541 B.n118 10.6151
R2221 B.n537 B.n118 10.6151
R2222 B.n537 B.n536 10.6151
R2223 B.n536 B.n535 10.6151
R2224 B.n535 B.n120 10.6151
R2225 B.n531 B.n120 10.6151
R2226 B.n531 B.n530 10.6151
R2227 B.n530 B.n529 10.6151
R2228 B.n529 B.n122 10.6151
R2229 B.n525 B.n122 10.6151
R2230 B.n525 B.n524 10.6151
R2231 B.n524 B.n523 10.6151
R2232 B.n523 B.n124 10.6151
R2233 B.n519 B.n124 10.6151
R2234 B.n519 B.n518 10.6151
R2235 B.n518 B.n517 10.6151
R2236 B.n517 B.n126 10.6151
R2237 B.n513 B.n126 10.6151
R2238 B.n513 B.n512 10.6151
R2239 B.n512 B.n511 10.6151
R2240 B.n511 B.n128 10.6151
R2241 B.n507 B.n128 10.6151
R2242 B.n507 B.n506 10.6151
R2243 B.n506 B.n505 10.6151
R2244 B.n505 B.n130 10.6151
R2245 B.n501 B.n130 10.6151
R2246 B.n501 B.n500 10.6151
R2247 B.n500 B.n499 10.6151
R2248 B.n499 B.n132 10.6151
R2249 B.n495 B.n132 10.6151
R2250 B.n495 B.n494 10.6151
R2251 B.n494 B.n493 10.6151
R2252 B.n493 B.n134 10.6151
R2253 B.n489 B.n134 10.6151
R2254 B.n489 B.n488 10.6151
R2255 B.n488 B.n487 10.6151
R2256 B.n487 B.n136 10.6151
R2257 B.n483 B.n136 10.6151
R2258 B.n483 B.n482 10.6151
R2259 B.n482 B.n481 10.6151
R2260 B.n481 B.n138 10.6151
R2261 B.n477 B.n138 10.6151
R2262 B.n477 B.n476 10.6151
R2263 B.n476 B.n475 10.6151
R2264 B.n475 B.n140 10.6151
R2265 B.n471 B.n140 10.6151
R2266 B.n471 B.n470 10.6151
R2267 B.n470 B.n469 10.6151
R2268 B.n469 B.n142 10.6151
R2269 B.n465 B.n142 10.6151
R2270 B.n465 B.n464 10.6151
R2271 B.n464 B.n463 10.6151
R2272 B.n463 B.n144 10.6151
R2273 B.n459 B.n144 10.6151
R2274 B.n459 B.n458 10.6151
R2275 B.n458 B.n457 10.6151
R2276 B.n457 B.n146 10.6151
R2277 B.n225 B.n1 10.6151
R2278 B.n226 B.n225 10.6151
R2279 B.n227 B.n226 10.6151
R2280 B.n227 B.n222 10.6151
R2281 B.n231 B.n222 10.6151
R2282 B.n232 B.n231 10.6151
R2283 B.n233 B.n232 10.6151
R2284 B.n233 B.n220 10.6151
R2285 B.n237 B.n220 10.6151
R2286 B.n238 B.n237 10.6151
R2287 B.n239 B.n238 10.6151
R2288 B.n239 B.n218 10.6151
R2289 B.n243 B.n218 10.6151
R2290 B.n244 B.n243 10.6151
R2291 B.n245 B.n244 10.6151
R2292 B.n245 B.n216 10.6151
R2293 B.n249 B.n216 10.6151
R2294 B.n250 B.n249 10.6151
R2295 B.n251 B.n250 10.6151
R2296 B.n251 B.n214 10.6151
R2297 B.n255 B.n214 10.6151
R2298 B.n256 B.n255 10.6151
R2299 B.n257 B.n256 10.6151
R2300 B.n257 B.n212 10.6151
R2301 B.n261 B.n212 10.6151
R2302 B.n262 B.n261 10.6151
R2303 B.n263 B.n262 10.6151
R2304 B.n263 B.n210 10.6151
R2305 B.n267 B.n210 10.6151
R2306 B.n268 B.n267 10.6151
R2307 B.n269 B.n268 10.6151
R2308 B.n269 B.n208 10.6151
R2309 B.n273 B.n208 10.6151
R2310 B.n274 B.n273 10.6151
R2311 B.n275 B.n274 10.6151
R2312 B.n275 B.n206 10.6151
R2313 B.n279 B.n206 10.6151
R2314 B.n280 B.n279 10.6151
R2315 B.n281 B.n280 10.6151
R2316 B.n281 B.n204 10.6151
R2317 B.n285 B.n204 10.6151
R2318 B.n286 B.n285 10.6151
R2319 B.n287 B.n286 10.6151
R2320 B.n287 B.n202 10.6151
R2321 B.n291 B.n202 10.6151
R2322 B.n292 B.n291 10.6151
R2323 B.n293 B.n292 10.6151
R2324 B.n293 B.n200 10.6151
R2325 B.n297 B.n200 10.6151
R2326 B.n298 B.n297 10.6151
R2327 B.n299 B.n298 10.6151
R2328 B.n299 B.n198 10.6151
R2329 B.n303 B.n198 10.6151
R2330 B.n304 B.n303 10.6151
R2331 B.n305 B.n304 10.6151
R2332 B.n305 B.n196 10.6151
R2333 B.n309 B.n196 10.6151
R2334 B.n310 B.n309 10.6151
R2335 B.n311 B.n310 10.6151
R2336 B.n311 B.n194 10.6151
R2337 B.n315 B.n194 10.6151
R2338 B.n316 B.n315 10.6151
R2339 B.n317 B.n192 10.6151
R2340 B.n321 B.n192 10.6151
R2341 B.n322 B.n321 10.6151
R2342 B.n323 B.n322 10.6151
R2343 B.n323 B.n190 10.6151
R2344 B.n327 B.n190 10.6151
R2345 B.n328 B.n327 10.6151
R2346 B.n329 B.n328 10.6151
R2347 B.n329 B.n188 10.6151
R2348 B.n333 B.n188 10.6151
R2349 B.n334 B.n333 10.6151
R2350 B.n335 B.n334 10.6151
R2351 B.n335 B.n186 10.6151
R2352 B.n339 B.n186 10.6151
R2353 B.n340 B.n339 10.6151
R2354 B.n341 B.n340 10.6151
R2355 B.n341 B.n184 10.6151
R2356 B.n345 B.n184 10.6151
R2357 B.n346 B.n345 10.6151
R2358 B.n347 B.n346 10.6151
R2359 B.n347 B.n182 10.6151
R2360 B.n351 B.n182 10.6151
R2361 B.n352 B.n351 10.6151
R2362 B.n353 B.n352 10.6151
R2363 B.n353 B.n180 10.6151
R2364 B.n357 B.n180 10.6151
R2365 B.n358 B.n357 10.6151
R2366 B.n359 B.n358 10.6151
R2367 B.n359 B.n178 10.6151
R2368 B.n363 B.n178 10.6151
R2369 B.n364 B.n363 10.6151
R2370 B.n365 B.n364 10.6151
R2371 B.n365 B.n176 10.6151
R2372 B.n369 B.n176 10.6151
R2373 B.n370 B.n369 10.6151
R2374 B.n371 B.n370 10.6151
R2375 B.n371 B.n174 10.6151
R2376 B.n375 B.n174 10.6151
R2377 B.n376 B.n375 10.6151
R2378 B.n378 B.n170 10.6151
R2379 B.n382 B.n170 10.6151
R2380 B.n383 B.n382 10.6151
R2381 B.n384 B.n383 10.6151
R2382 B.n384 B.n168 10.6151
R2383 B.n388 B.n168 10.6151
R2384 B.n389 B.n388 10.6151
R2385 B.n393 B.n389 10.6151
R2386 B.n397 B.n166 10.6151
R2387 B.n398 B.n397 10.6151
R2388 B.n399 B.n398 10.6151
R2389 B.n399 B.n164 10.6151
R2390 B.n403 B.n164 10.6151
R2391 B.n404 B.n403 10.6151
R2392 B.n405 B.n404 10.6151
R2393 B.n405 B.n162 10.6151
R2394 B.n409 B.n162 10.6151
R2395 B.n410 B.n409 10.6151
R2396 B.n411 B.n410 10.6151
R2397 B.n411 B.n160 10.6151
R2398 B.n415 B.n160 10.6151
R2399 B.n416 B.n415 10.6151
R2400 B.n417 B.n416 10.6151
R2401 B.n417 B.n158 10.6151
R2402 B.n421 B.n158 10.6151
R2403 B.n422 B.n421 10.6151
R2404 B.n423 B.n422 10.6151
R2405 B.n423 B.n156 10.6151
R2406 B.n427 B.n156 10.6151
R2407 B.n428 B.n427 10.6151
R2408 B.n429 B.n428 10.6151
R2409 B.n429 B.n154 10.6151
R2410 B.n433 B.n154 10.6151
R2411 B.n434 B.n433 10.6151
R2412 B.n435 B.n434 10.6151
R2413 B.n435 B.n152 10.6151
R2414 B.n439 B.n152 10.6151
R2415 B.n440 B.n439 10.6151
R2416 B.n441 B.n440 10.6151
R2417 B.n441 B.n150 10.6151
R2418 B.n445 B.n150 10.6151
R2419 B.n446 B.n445 10.6151
R2420 B.n447 B.n446 10.6151
R2421 B.n447 B.n148 10.6151
R2422 B.n451 B.n148 10.6151
R2423 B.n452 B.n451 10.6151
R2424 B.n453 B.n452 10.6151
R2425 B.n877 B.n0 8.11757
R2426 B.n877 B.n1 8.11757
R2427 B.n721 B.n720 6.5566
R2428 B.n708 B.n62 6.5566
R2429 B.n378 B.n377 6.5566
R2430 B.n393 B.n392 6.5566
R2431 B.n722 B.n721 4.05904
R2432 B.n705 B.n62 4.05904
R2433 B.n377 B.n376 4.05904
R2434 B.n392 B.n166 4.05904
C0 VDD2 B 2.64341f
C1 VDD1 VDD2 2.31061f
C2 VDD1 B 2.51732f
C3 VP VDD2 0.610257f
C4 VP B 2.36959f
C5 VP VDD1 10.7927f
C6 VTAIL VDD2 10.2494f
C7 VN VDD2 10.34f
C8 VTAIL B 3.68708f
C9 VN B 1.33005f
C10 VTAIL VDD1 10.1967f
C11 VN VDD1 0.153773f
C12 VP VTAIL 11.1118f
C13 VP VN 8.603769f
C14 VN VTAIL 11.097501f
C15 VDD2 w_n4738_n3254# 2.98286f
C16 w_n4738_n3254# B 10.7404f
C17 VDD1 w_n4738_n3254# 2.8284f
C18 VP w_n4738_n3254# 10.8079f
C19 VTAIL w_n4738_n3254# 3.1591f
C20 VN w_n4738_n3254# 10.1904f
C21 VDD2 VSUBS 2.23674f
C22 VDD1 VSUBS 2.03164f
C23 VTAIL VSUBS 1.332692f
C24 VN VSUBS 7.996409f
C25 VP VSUBS 4.475866f
C26 B VSUBS 5.58033f
C27 w_n4738_n3254# VSUBS 0.189956p
C28 B.n0 VSUBS 0.008256f
C29 B.n1 VSUBS 0.008256f
C30 B.n2 VSUBS 0.012209f
C31 B.n3 VSUBS 0.009356f
C32 B.n4 VSUBS 0.009356f
C33 B.n5 VSUBS 0.009356f
C34 B.n6 VSUBS 0.009356f
C35 B.n7 VSUBS 0.009356f
C36 B.n8 VSUBS 0.009356f
C37 B.n9 VSUBS 0.009356f
C38 B.n10 VSUBS 0.009356f
C39 B.n11 VSUBS 0.009356f
C40 B.n12 VSUBS 0.009356f
C41 B.n13 VSUBS 0.009356f
C42 B.n14 VSUBS 0.009356f
C43 B.n15 VSUBS 0.009356f
C44 B.n16 VSUBS 0.009356f
C45 B.n17 VSUBS 0.009356f
C46 B.n18 VSUBS 0.009356f
C47 B.n19 VSUBS 0.009356f
C48 B.n20 VSUBS 0.009356f
C49 B.n21 VSUBS 0.009356f
C50 B.n22 VSUBS 0.009356f
C51 B.n23 VSUBS 0.009356f
C52 B.n24 VSUBS 0.009356f
C53 B.n25 VSUBS 0.009356f
C54 B.n26 VSUBS 0.009356f
C55 B.n27 VSUBS 0.009356f
C56 B.n28 VSUBS 0.009356f
C57 B.n29 VSUBS 0.009356f
C58 B.n30 VSUBS 0.009356f
C59 B.n31 VSUBS 0.009356f
C60 B.n32 VSUBS 0.009356f
C61 B.n33 VSUBS 0.022664f
C62 B.n34 VSUBS 0.009356f
C63 B.n35 VSUBS 0.009356f
C64 B.n36 VSUBS 0.009356f
C65 B.n37 VSUBS 0.009356f
C66 B.n38 VSUBS 0.009356f
C67 B.n39 VSUBS 0.009356f
C68 B.n40 VSUBS 0.009356f
C69 B.n41 VSUBS 0.009356f
C70 B.n42 VSUBS 0.009356f
C71 B.n43 VSUBS 0.009356f
C72 B.n44 VSUBS 0.009356f
C73 B.n45 VSUBS 0.009356f
C74 B.n46 VSUBS 0.009356f
C75 B.n47 VSUBS 0.009356f
C76 B.n48 VSUBS 0.009356f
C77 B.n49 VSUBS 0.009356f
C78 B.n50 VSUBS 0.009356f
C79 B.n51 VSUBS 0.009356f
C80 B.n52 VSUBS 0.009356f
C81 B.n53 VSUBS 0.009356f
C82 B.t7 VSUBS 0.26528f
C83 B.t8 VSUBS 0.310084f
C84 B.t6 VSUBS 1.97121f
C85 B.n54 VSUBS 0.495437f
C86 B.n55 VSUBS 0.326998f
C87 B.n56 VSUBS 0.009356f
C88 B.n57 VSUBS 0.009356f
C89 B.n58 VSUBS 0.009356f
C90 B.n59 VSUBS 0.009356f
C91 B.t1 VSUBS 0.265284f
C92 B.t2 VSUBS 0.310087f
C93 B.t0 VSUBS 1.97121f
C94 B.n60 VSUBS 0.495433f
C95 B.n61 VSUBS 0.326994f
C96 B.n62 VSUBS 0.021677f
C97 B.n63 VSUBS 0.009356f
C98 B.n64 VSUBS 0.009356f
C99 B.n65 VSUBS 0.009356f
C100 B.n66 VSUBS 0.009356f
C101 B.n67 VSUBS 0.009356f
C102 B.n68 VSUBS 0.009356f
C103 B.n69 VSUBS 0.009356f
C104 B.n70 VSUBS 0.009356f
C105 B.n71 VSUBS 0.009356f
C106 B.n72 VSUBS 0.009356f
C107 B.n73 VSUBS 0.009356f
C108 B.n74 VSUBS 0.009356f
C109 B.n75 VSUBS 0.009356f
C110 B.n76 VSUBS 0.009356f
C111 B.n77 VSUBS 0.009356f
C112 B.n78 VSUBS 0.009356f
C113 B.n79 VSUBS 0.009356f
C114 B.n80 VSUBS 0.009356f
C115 B.n81 VSUBS 0.009356f
C116 B.n82 VSUBS 0.023291f
C117 B.n83 VSUBS 0.009356f
C118 B.n84 VSUBS 0.009356f
C119 B.n85 VSUBS 0.009356f
C120 B.n86 VSUBS 0.009356f
C121 B.n87 VSUBS 0.009356f
C122 B.n88 VSUBS 0.009356f
C123 B.n89 VSUBS 0.009356f
C124 B.n90 VSUBS 0.009356f
C125 B.n91 VSUBS 0.009356f
C126 B.n92 VSUBS 0.009356f
C127 B.n93 VSUBS 0.009356f
C128 B.n94 VSUBS 0.009356f
C129 B.n95 VSUBS 0.009356f
C130 B.n96 VSUBS 0.009356f
C131 B.n97 VSUBS 0.009356f
C132 B.n98 VSUBS 0.009356f
C133 B.n99 VSUBS 0.009356f
C134 B.n100 VSUBS 0.009356f
C135 B.n101 VSUBS 0.009356f
C136 B.n102 VSUBS 0.009356f
C137 B.n103 VSUBS 0.009356f
C138 B.n104 VSUBS 0.009356f
C139 B.n105 VSUBS 0.009356f
C140 B.n106 VSUBS 0.009356f
C141 B.n107 VSUBS 0.009356f
C142 B.n108 VSUBS 0.009356f
C143 B.n109 VSUBS 0.009356f
C144 B.n110 VSUBS 0.009356f
C145 B.n111 VSUBS 0.009356f
C146 B.n112 VSUBS 0.009356f
C147 B.n113 VSUBS 0.009356f
C148 B.n114 VSUBS 0.009356f
C149 B.n115 VSUBS 0.009356f
C150 B.n116 VSUBS 0.009356f
C151 B.n117 VSUBS 0.009356f
C152 B.n118 VSUBS 0.009356f
C153 B.n119 VSUBS 0.009356f
C154 B.n120 VSUBS 0.009356f
C155 B.n121 VSUBS 0.009356f
C156 B.n122 VSUBS 0.009356f
C157 B.n123 VSUBS 0.009356f
C158 B.n124 VSUBS 0.009356f
C159 B.n125 VSUBS 0.009356f
C160 B.n126 VSUBS 0.009356f
C161 B.n127 VSUBS 0.009356f
C162 B.n128 VSUBS 0.009356f
C163 B.n129 VSUBS 0.009356f
C164 B.n130 VSUBS 0.009356f
C165 B.n131 VSUBS 0.009356f
C166 B.n132 VSUBS 0.009356f
C167 B.n133 VSUBS 0.009356f
C168 B.n134 VSUBS 0.009356f
C169 B.n135 VSUBS 0.009356f
C170 B.n136 VSUBS 0.009356f
C171 B.n137 VSUBS 0.009356f
C172 B.n138 VSUBS 0.009356f
C173 B.n139 VSUBS 0.009356f
C174 B.n140 VSUBS 0.009356f
C175 B.n141 VSUBS 0.009356f
C176 B.n142 VSUBS 0.009356f
C177 B.n143 VSUBS 0.009356f
C178 B.n144 VSUBS 0.009356f
C179 B.n145 VSUBS 0.009356f
C180 B.n146 VSUBS 0.023692f
C181 B.n147 VSUBS 0.009356f
C182 B.n148 VSUBS 0.009356f
C183 B.n149 VSUBS 0.009356f
C184 B.n150 VSUBS 0.009356f
C185 B.n151 VSUBS 0.009356f
C186 B.n152 VSUBS 0.009356f
C187 B.n153 VSUBS 0.009356f
C188 B.n154 VSUBS 0.009356f
C189 B.n155 VSUBS 0.009356f
C190 B.n156 VSUBS 0.009356f
C191 B.n157 VSUBS 0.009356f
C192 B.n158 VSUBS 0.009356f
C193 B.n159 VSUBS 0.009356f
C194 B.n160 VSUBS 0.009356f
C195 B.n161 VSUBS 0.009356f
C196 B.n162 VSUBS 0.009356f
C197 B.n163 VSUBS 0.009356f
C198 B.n164 VSUBS 0.009356f
C199 B.n165 VSUBS 0.009356f
C200 B.n166 VSUBS 0.006467f
C201 B.n167 VSUBS 0.009356f
C202 B.n168 VSUBS 0.009356f
C203 B.n169 VSUBS 0.009356f
C204 B.n170 VSUBS 0.009356f
C205 B.n171 VSUBS 0.009356f
C206 B.t11 VSUBS 0.26528f
C207 B.t10 VSUBS 0.310084f
C208 B.t9 VSUBS 1.97121f
C209 B.n172 VSUBS 0.495437f
C210 B.n173 VSUBS 0.326998f
C211 B.n174 VSUBS 0.009356f
C212 B.n175 VSUBS 0.009356f
C213 B.n176 VSUBS 0.009356f
C214 B.n177 VSUBS 0.009356f
C215 B.n178 VSUBS 0.009356f
C216 B.n179 VSUBS 0.009356f
C217 B.n180 VSUBS 0.009356f
C218 B.n181 VSUBS 0.009356f
C219 B.n182 VSUBS 0.009356f
C220 B.n183 VSUBS 0.009356f
C221 B.n184 VSUBS 0.009356f
C222 B.n185 VSUBS 0.009356f
C223 B.n186 VSUBS 0.009356f
C224 B.n187 VSUBS 0.009356f
C225 B.n188 VSUBS 0.009356f
C226 B.n189 VSUBS 0.009356f
C227 B.n190 VSUBS 0.009356f
C228 B.n191 VSUBS 0.009356f
C229 B.n192 VSUBS 0.009356f
C230 B.n193 VSUBS 0.022664f
C231 B.n194 VSUBS 0.009356f
C232 B.n195 VSUBS 0.009356f
C233 B.n196 VSUBS 0.009356f
C234 B.n197 VSUBS 0.009356f
C235 B.n198 VSUBS 0.009356f
C236 B.n199 VSUBS 0.009356f
C237 B.n200 VSUBS 0.009356f
C238 B.n201 VSUBS 0.009356f
C239 B.n202 VSUBS 0.009356f
C240 B.n203 VSUBS 0.009356f
C241 B.n204 VSUBS 0.009356f
C242 B.n205 VSUBS 0.009356f
C243 B.n206 VSUBS 0.009356f
C244 B.n207 VSUBS 0.009356f
C245 B.n208 VSUBS 0.009356f
C246 B.n209 VSUBS 0.009356f
C247 B.n210 VSUBS 0.009356f
C248 B.n211 VSUBS 0.009356f
C249 B.n212 VSUBS 0.009356f
C250 B.n213 VSUBS 0.009356f
C251 B.n214 VSUBS 0.009356f
C252 B.n215 VSUBS 0.009356f
C253 B.n216 VSUBS 0.009356f
C254 B.n217 VSUBS 0.009356f
C255 B.n218 VSUBS 0.009356f
C256 B.n219 VSUBS 0.009356f
C257 B.n220 VSUBS 0.009356f
C258 B.n221 VSUBS 0.009356f
C259 B.n222 VSUBS 0.009356f
C260 B.n223 VSUBS 0.009356f
C261 B.n224 VSUBS 0.009356f
C262 B.n225 VSUBS 0.009356f
C263 B.n226 VSUBS 0.009356f
C264 B.n227 VSUBS 0.009356f
C265 B.n228 VSUBS 0.009356f
C266 B.n229 VSUBS 0.009356f
C267 B.n230 VSUBS 0.009356f
C268 B.n231 VSUBS 0.009356f
C269 B.n232 VSUBS 0.009356f
C270 B.n233 VSUBS 0.009356f
C271 B.n234 VSUBS 0.009356f
C272 B.n235 VSUBS 0.009356f
C273 B.n236 VSUBS 0.009356f
C274 B.n237 VSUBS 0.009356f
C275 B.n238 VSUBS 0.009356f
C276 B.n239 VSUBS 0.009356f
C277 B.n240 VSUBS 0.009356f
C278 B.n241 VSUBS 0.009356f
C279 B.n242 VSUBS 0.009356f
C280 B.n243 VSUBS 0.009356f
C281 B.n244 VSUBS 0.009356f
C282 B.n245 VSUBS 0.009356f
C283 B.n246 VSUBS 0.009356f
C284 B.n247 VSUBS 0.009356f
C285 B.n248 VSUBS 0.009356f
C286 B.n249 VSUBS 0.009356f
C287 B.n250 VSUBS 0.009356f
C288 B.n251 VSUBS 0.009356f
C289 B.n252 VSUBS 0.009356f
C290 B.n253 VSUBS 0.009356f
C291 B.n254 VSUBS 0.009356f
C292 B.n255 VSUBS 0.009356f
C293 B.n256 VSUBS 0.009356f
C294 B.n257 VSUBS 0.009356f
C295 B.n258 VSUBS 0.009356f
C296 B.n259 VSUBS 0.009356f
C297 B.n260 VSUBS 0.009356f
C298 B.n261 VSUBS 0.009356f
C299 B.n262 VSUBS 0.009356f
C300 B.n263 VSUBS 0.009356f
C301 B.n264 VSUBS 0.009356f
C302 B.n265 VSUBS 0.009356f
C303 B.n266 VSUBS 0.009356f
C304 B.n267 VSUBS 0.009356f
C305 B.n268 VSUBS 0.009356f
C306 B.n269 VSUBS 0.009356f
C307 B.n270 VSUBS 0.009356f
C308 B.n271 VSUBS 0.009356f
C309 B.n272 VSUBS 0.009356f
C310 B.n273 VSUBS 0.009356f
C311 B.n274 VSUBS 0.009356f
C312 B.n275 VSUBS 0.009356f
C313 B.n276 VSUBS 0.009356f
C314 B.n277 VSUBS 0.009356f
C315 B.n278 VSUBS 0.009356f
C316 B.n279 VSUBS 0.009356f
C317 B.n280 VSUBS 0.009356f
C318 B.n281 VSUBS 0.009356f
C319 B.n282 VSUBS 0.009356f
C320 B.n283 VSUBS 0.009356f
C321 B.n284 VSUBS 0.009356f
C322 B.n285 VSUBS 0.009356f
C323 B.n286 VSUBS 0.009356f
C324 B.n287 VSUBS 0.009356f
C325 B.n288 VSUBS 0.009356f
C326 B.n289 VSUBS 0.009356f
C327 B.n290 VSUBS 0.009356f
C328 B.n291 VSUBS 0.009356f
C329 B.n292 VSUBS 0.009356f
C330 B.n293 VSUBS 0.009356f
C331 B.n294 VSUBS 0.009356f
C332 B.n295 VSUBS 0.009356f
C333 B.n296 VSUBS 0.009356f
C334 B.n297 VSUBS 0.009356f
C335 B.n298 VSUBS 0.009356f
C336 B.n299 VSUBS 0.009356f
C337 B.n300 VSUBS 0.009356f
C338 B.n301 VSUBS 0.009356f
C339 B.n302 VSUBS 0.009356f
C340 B.n303 VSUBS 0.009356f
C341 B.n304 VSUBS 0.009356f
C342 B.n305 VSUBS 0.009356f
C343 B.n306 VSUBS 0.009356f
C344 B.n307 VSUBS 0.009356f
C345 B.n308 VSUBS 0.009356f
C346 B.n309 VSUBS 0.009356f
C347 B.n310 VSUBS 0.009356f
C348 B.n311 VSUBS 0.009356f
C349 B.n312 VSUBS 0.009356f
C350 B.n313 VSUBS 0.009356f
C351 B.n314 VSUBS 0.009356f
C352 B.n315 VSUBS 0.009356f
C353 B.n316 VSUBS 0.022664f
C354 B.n317 VSUBS 0.023291f
C355 B.n318 VSUBS 0.023291f
C356 B.n319 VSUBS 0.009356f
C357 B.n320 VSUBS 0.009356f
C358 B.n321 VSUBS 0.009356f
C359 B.n322 VSUBS 0.009356f
C360 B.n323 VSUBS 0.009356f
C361 B.n324 VSUBS 0.009356f
C362 B.n325 VSUBS 0.009356f
C363 B.n326 VSUBS 0.009356f
C364 B.n327 VSUBS 0.009356f
C365 B.n328 VSUBS 0.009356f
C366 B.n329 VSUBS 0.009356f
C367 B.n330 VSUBS 0.009356f
C368 B.n331 VSUBS 0.009356f
C369 B.n332 VSUBS 0.009356f
C370 B.n333 VSUBS 0.009356f
C371 B.n334 VSUBS 0.009356f
C372 B.n335 VSUBS 0.009356f
C373 B.n336 VSUBS 0.009356f
C374 B.n337 VSUBS 0.009356f
C375 B.n338 VSUBS 0.009356f
C376 B.n339 VSUBS 0.009356f
C377 B.n340 VSUBS 0.009356f
C378 B.n341 VSUBS 0.009356f
C379 B.n342 VSUBS 0.009356f
C380 B.n343 VSUBS 0.009356f
C381 B.n344 VSUBS 0.009356f
C382 B.n345 VSUBS 0.009356f
C383 B.n346 VSUBS 0.009356f
C384 B.n347 VSUBS 0.009356f
C385 B.n348 VSUBS 0.009356f
C386 B.n349 VSUBS 0.009356f
C387 B.n350 VSUBS 0.009356f
C388 B.n351 VSUBS 0.009356f
C389 B.n352 VSUBS 0.009356f
C390 B.n353 VSUBS 0.009356f
C391 B.n354 VSUBS 0.009356f
C392 B.n355 VSUBS 0.009356f
C393 B.n356 VSUBS 0.009356f
C394 B.n357 VSUBS 0.009356f
C395 B.n358 VSUBS 0.009356f
C396 B.n359 VSUBS 0.009356f
C397 B.n360 VSUBS 0.009356f
C398 B.n361 VSUBS 0.009356f
C399 B.n362 VSUBS 0.009356f
C400 B.n363 VSUBS 0.009356f
C401 B.n364 VSUBS 0.009356f
C402 B.n365 VSUBS 0.009356f
C403 B.n366 VSUBS 0.009356f
C404 B.n367 VSUBS 0.009356f
C405 B.n368 VSUBS 0.009356f
C406 B.n369 VSUBS 0.009356f
C407 B.n370 VSUBS 0.009356f
C408 B.n371 VSUBS 0.009356f
C409 B.n372 VSUBS 0.009356f
C410 B.n373 VSUBS 0.009356f
C411 B.n374 VSUBS 0.009356f
C412 B.n375 VSUBS 0.009356f
C413 B.n376 VSUBS 0.006467f
C414 B.n377 VSUBS 0.021677f
C415 B.n378 VSUBS 0.007568f
C416 B.n379 VSUBS 0.009356f
C417 B.n380 VSUBS 0.009356f
C418 B.n381 VSUBS 0.009356f
C419 B.n382 VSUBS 0.009356f
C420 B.n383 VSUBS 0.009356f
C421 B.n384 VSUBS 0.009356f
C422 B.n385 VSUBS 0.009356f
C423 B.n386 VSUBS 0.009356f
C424 B.n387 VSUBS 0.009356f
C425 B.n388 VSUBS 0.009356f
C426 B.n389 VSUBS 0.009356f
C427 B.t5 VSUBS 0.265284f
C428 B.t4 VSUBS 0.310087f
C429 B.t3 VSUBS 1.97121f
C430 B.n390 VSUBS 0.495433f
C431 B.n391 VSUBS 0.326994f
C432 B.n392 VSUBS 0.021677f
C433 B.n393 VSUBS 0.007568f
C434 B.n394 VSUBS 0.009356f
C435 B.n395 VSUBS 0.009356f
C436 B.n396 VSUBS 0.009356f
C437 B.n397 VSUBS 0.009356f
C438 B.n398 VSUBS 0.009356f
C439 B.n399 VSUBS 0.009356f
C440 B.n400 VSUBS 0.009356f
C441 B.n401 VSUBS 0.009356f
C442 B.n402 VSUBS 0.009356f
C443 B.n403 VSUBS 0.009356f
C444 B.n404 VSUBS 0.009356f
C445 B.n405 VSUBS 0.009356f
C446 B.n406 VSUBS 0.009356f
C447 B.n407 VSUBS 0.009356f
C448 B.n408 VSUBS 0.009356f
C449 B.n409 VSUBS 0.009356f
C450 B.n410 VSUBS 0.009356f
C451 B.n411 VSUBS 0.009356f
C452 B.n412 VSUBS 0.009356f
C453 B.n413 VSUBS 0.009356f
C454 B.n414 VSUBS 0.009356f
C455 B.n415 VSUBS 0.009356f
C456 B.n416 VSUBS 0.009356f
C457 B.n417 VSUBS 0.009356f
C458 B.n418 VSUBS 0.009356f
C459 B.n419 VSUBS 0.009356f
C460 B.n420 VSUBS 0.009356f
C461 B.n421 VSUBS 0.009356f
C462 B.n422 VSUBS 0.009356f
C463 B.n423 VSUBS 0.009356f
C464 B.n424 VSUBS 0.009356f
C465 B.n425 VSUBS 0.009356f
C466 B.n426 VSUBS 0.009356f
C467 B.n427 VSUBS 0.009356f
C468 B.n428 VSUBS 0.009356f
C469 B.n429 VSUBS 0.009356f
C470 B.n430 VSUBS 0.009356f
C471 B.n431 VSUBS 0.009356f
C472 B.n432 VSUBS 0.009356f
C473 B.n433 VSUBS 0.009356f
C474 B.n434 VSUBS 0.009356f
C475 B.n435 VSUBS 0.009356f
C476 B.n436 VSUBS 0.009356f
C477 B.n437 VSUBS 0.009356f
C478 B.n438 VSUBS 0.009356f
C479 B.n439 VSUBS 0.009356f
C480 B.n440 VSUBS 0.009356f
C481 B.n441 VSUBS 0.009356f
C482 B.n442 VSUBS 0.009356f
C483 B.n443 VSUBS 0.009356f
C484 B.n444 VSUBS 0.009356f
C485 B.n445 VSUBS 0.009356f
C486 B.n446 VSUBS 0.009356f
C487 B.n447 VSUBS 0.009356f
C488 B.n448 VSUBS 0.009356f
C489 B.n449 VSUBS 0.009356f
C490 B.n450 VSUBS 0.009356f
C491 B.n451 VSUBS 0.009356f
C492 B.n452 VSUBS 0.009356f
C493 B.n453 VSUBS 0.022263f
C494 B.n454 VSUBS 0.023291f
C495 B.n455 VSUBS 0.022664f
C496 B.n456 VSUBS 0.009356f
C497 B.n457 VSUBS 0.009356f
C498 B.n458 VSUBS 0.009356f
C499 B.n459 VSUBS 0.009356f
C500 B.n460 VSUBS 0.009356f
C501 B.n461 VSUBS 0.009356f
C502 B.n462 VSUBS 0.009356f
C503 B.n463 VSUBS 0.009356f
C504 B.n464 VSUBS 0.009356f
C505 B.n465 VSUBS 0.009356f
C506 B.n466 VSUBS 0.009356f
C507 B.n467 VSUBS 0.009356f
C508 B.n468 VSUBS 0.009356f
C509 B.n469 VSUBS 0.009356f
C510 B.n470 VSUBS 0.009356f
C511 B.n471 VSUBS 0.009356f
C512 B.n472 VSUBS 0.009356f
C513 B.n473 VSUBS 0.009356f
C514 B.n474 VSUBS 0.009356f
C515 B.n475 VSUBS 0.009356f
C516 B.n476 VSUBS 0.009356f
C517 B.n477 VSUBS 0.009356f
C518 B.n478 VSUBS 0.009356f
C519 B.n479 VSUBS 0.009356f
C520 B.n480 VSUBS 0.009356f
C521 B.n481 VSUBS 0.009356f
C522 B.n482 VSUBS 0.009356f
C523 B.n483 VSUBS 0.009356f
C524 B.n484 VSUBS 0.009356f
C525 B.n485 VSUBS 0.009356f
C526 B.n486 VSUBS 0.009356f
C527 B.n487 VSUBS 0.009356f
C528 B.n488 VSUBS 0.009356f
C529 B.n489 VSUBS 0.009356f
C530 B.n490 VSUBS 0.009356f
C531 B.n491 VSUBS 0.009356f
C532 B.n492 VSUBS 0.009356f
C533 B.n493 VSUBS 0.009356f
C534 B.n494 VSUBS 0.009356f
C535 B.n495 VSUBS 0.009356f
C536 B.n496 VSUBS 0.009356f
C537 B.n497 VSUBS 0.009356f
C538 B.n498 VSUBS 0.009356f
C539 B.n499 VSUBS 0.009356f
C540 B.n500 VSUBS 0.009356f
C541 B.n501 VSUBS 0.009356f
C542 B.n502 VSUBS 0.009356f
C543 B.n503 VSUBS 0.009356f
C544 B.n504 VSUBS 0.009356f
C545 B.n505 VSUBS 0.009356f
C546 B.n506 VSUBS 0.009356f
C547 B.n507 VSUBS 0.009356f
C548 B.n508 VSUBS 0.009356f
C549 B.n509 VSUBS 0.009356f
C550 B.n510 VSUBS 0.009356f
C551 B.n511 VSUBS 0.009356f
C552 B.n512 VSUBS 0.009356f
C553 B.n513 VSUBS 0.009356f
C554 B.n514 VSUBS 0.009356f
C555 B.n515 VSUBS 0.009356f
C556 B.n516 VSUBS 0.009356f
C557 B.n517 VSUBS 0.009356f
C558 B.n518 VSUBS 0.009356f
C559 B.n519 VSUBS 0.009356f
C560 B.n520 VSUBS 0.009356f
C561 B.n521 VSUBS 0.009356f
C562 B.n522 VSUBS 0.009356f
C563 B.n523 VSUBS 0.009356f
C564 B.n524 VSUBS 0.009356f
C565 B.n525 VSUBS 0.009356f
C566 B.n526 VSUBS 0.009356f
C567 B.n527 VSUBS 0.009356f
C568 B.n528 VSUBS 0.009356f
C569 B.n529 VSUBS 0.009356f
C570 B.n530 VSUBS 0.009356f
C571 B.n531 VSUBS 0.009356f
C572 B.n532 VSUBS 0.009356f
C573 B.n533 VSUBS 0.009356f
C574 B.n534 VSUBS 0.009356f
C575 B.n535 VSUBS 0.009356f
C576 B.n536 VSUBS 0.009356f
C577 B.n537 VSUBS 0.009356f
C578 B.n538 VSUBS 0.009356f
C579 B.n539 VSUBS 0.009356f
C580 B.n540 VSUBS 0.009356f
C581 B.n541 VSUBS 0.009356f
C582 B.n542 VSUBS 0.009356f
C583 B.n543 VSUBS 0.009356f
C584 B.n544 VSUBS 0.009356f
C585 B.n545 VSUBS 0.009356f
C586 B.n546 VSUBS 0.009356f
C587 B.n547 VSUBS 0.009356f
C588 B.n548 VSUBS 0.009356f
C589 B.n549 VSUBS 0.009356f
C590 B.n550 VSUBS 0.009356f
C591 B.n551 VSUBS 0.009356f
C592 B.n552 VSUBS 0.009356f
C593 B.n553 VSUBS 0.009356f
C594 B.n554 VSUBS 0.009356f
C595 B.n555 VSUBS 0.009356f
C596 B.n556 VSUBS 0.009356f
C597 B.n557 VSUBS 0.009356f
C598 B.n558 VSUBS 0.009356f
C599 B.n559 VSUBS 0.009356f
C600 B.n560 VSUBS 0.009356f
C601 B.n561 VSUBS 0.009356f
C602 B.n562 VSUBS 0.009356f
C603 B.n563 VSUBS 0.009356f
C604 B.n564 VSUBS 0.009356f
C605 B.n565 VSUBS 0.009356f
C606 B.n566 VSUBS 0.009356f
C607 B.n567 VSUBS 0.009356f
C608 B.n568 VSUBS 0.009356f
C609 B.n569 VSUBS 0.009356f
C610 B.n570 VSUBS 0.009356f
C611 B.n571 VSUBS 0.009356f
C612 B.n572 VSUBS 0.009356f
C613 B.n573 VSUBS 0.009356f
C614 B.n574 VSUBS 0.009356f
C615 B.n575 VSUBS 0.009356f
C616 B.n576 VSUBS 0.009356f
C617 B.n577 VSUBS 0.009356f
C618 B.n578 VSUBS 0.009356f
C619 B.n579 VSUBS 0.009356f
C620 B.n580 VSUBS 0.009356f
C621 B.n581 VSUBS 0.009356f
C622 B.n582 VSUBS 0.009356f
C623 B.n583 VSUBS 0.009356f
C624 B.n584 VSUBS 0.009356f
C625 B.n585 VSUBS 0.009356f
C626 B.n586 VSUBS 0.009356f
C627 B.n587 VSUBS 0.009356f
C628 B.n588 VSUBS 0.009356f
C629 B.n589 VSUBS 0.009356f
C630 B.n590 VSUBS 0.009356f
C631 B.n591 VSUBS 0.009356f
C632 B.n592 VSUBS 0.009356f
C633 B.n593 VSUBS 0.009356f
C634 B.n594 VSUBS 0.009356f
C635 B.n595 VSUBS 0.009356f
C636 B.n596 VSUBS 0.009356f
C637 B.n597 VSUBS 0.009356f
C638 B.n598 VSUBS 0.009356f
C639 B.n599 VSUBS 0.009356f
C640 B.n600 VSUBS 0.009356f
C641 B.n601 VSUBS 0.009356f
C642 B.n602 VSUBS 0.009356f
C643 B.n603 VSUBS 0.009356f
C644 B.n604 VSUBS 0.009356f
C645 B.n605 VSUBS 0.009356f
C646 B.n606 VSUBS 0.009356f
C647 B.n607 VSUBS 0.009356f
C648 B.n608 VSUBS 0.009356f
C649 B.n609 VSUBS 0.009356f
C650 B.n610 VSUBS 0.009356f
C651 B.n611 VSUBS 0.009356f
C652 B.n612 VSUBS 0.009356f
C653 B.n613 VSUBS 0.009356f
C654 B.n614 VSUBS 0.009356f
C655 B.n615 VSUBS 0.009356f
C656 B.n616 VSUBS 0.009356f
C657 B.n617 VSUBS 0.009356f
C658 B.n618 VSUBS 0.009356f
C659 B.n619 VSUBS 0.009356f
C660 B.n620 VSUBS 0.009356f
C661 B.n621 VSUBS 0.009356f
C662 B.n622 VSUBS 0.009356f
C663 B.n623 VSUBS 0.009356f
C664 B.n624 VSUBS 0.009356f
C665 B.n625 VSUBS 0.009356f
C666 B.n626 VSUBS 0.009356f
C667 B.n627 VSUBS 0.009356f
C668 B.n628 VSUBS 0.009356f
C669 B.n629 VSUBS 0.009356f
C670 B.n630 VSUBS 0.009356f
C671 B.n631 VSUBS 0.009356f
C672 B.n632 VSUBS 0.009356f
C673 B.n633 VSUBS 0.009356f
C674 B.n634 VSUBS 0.009356f
C675 B.n635 VSUBS 0.009356f
C676 B.n636 VSUBS 0.009356f
C677 B.n637 VSUBS 0.009356f
C678 B.n638 VSUBS 0.009356f
C679 B.n639 VSUBS 0.009356f
C680 B.n640 VSUBS 0.009356f
C681 B.n641 VSUBS 0.009356f
C682 B.n642 VSUBS 0.009356f
C683 B.n643 VSUBS 0.009356f
C684 B.n644 VSUBS 0.009356f
C685 B.n645 VSUBS 0.022664f
C686 B.n646 VSUBS 0.022664f
C687 B.n647 VSUBS 0.023291f
C688 B.n648 VSUBS 0.009356f
C689 B.n649 VSUBS 0.009356f
C690 B.n650 VSUBS 0.009356f
C691 B.n651 VSUBS 0.009356f
C692 B.n652 VSUBS 0.009356f
C693 B.n653 VSUBS 0.009356f
C694 B.n654 VSUBS 0.009356f
C695 B.n655 VSUBS 0.009356f
C696 B.n656 VSUBS 0.009356f
C697 B.n657 VSUBS 0.009356f
C698 B.n658 VSUBS 0.009356f
C699 B.n659 VSUBS 0.009356f
C700 B.n660 VSUBS 0.009356f
C701 B.n661 VSUBS 0.009356f
C702 B.n662 VSUBS 0.009356f
C703 B.n663 VSUBS 0.009356f
C704 B.n664 VSUBS 0.009356f
C705 B.n665 VSUBS 0.009356f
C706 B.n666 VSUBS 0.009356f
C707 B.n667 VSUBS 0.009356f
C708 B.n668 VSUBS 0.009356f
C709 B.n669 VSUBS 0.009356f
C710 B.n670 VSUBS 0.009356f
C711 B.n671 VSUBS 0.009356f
C712 B.n672 VSUBS 0.009356f
C713 B.n673 VSUBS 0.009356f
C714 B.n674 VSUBS 0.009356f
C715 B.n675 VSUBS 0.009356f
C716 B.n676 VSUBS 0.009356f
C717 B.n677 VSUBS 0.009356f
C718 B.n678 VSUBS 0.009356f
C719 B.n679 VSUBS 0.009356f
C720 B.n680 VSUBS 0.009356f
C721 B.n681 VSUBS 0.009356f
C722 B.n682 VSUBS 0.009356f
C723 B.n683 VSUBS 0.009356f
C724 B.n684 VSUBS 0.009356f
C725 B.n685 VSUBS 0.009356f
C726 B.n686 VSUBS 0.009356f
C727 B.n687 VSUBS 0.009356f
C728 B.n688 VSUBS 0.009356f
C729 B.n689 VSUBS 0.009356f
C730 B.n690 VSUBS 0.009356f
C731 B.n691 VSUBS 0.009356f
C732 B.n692 VSUBS 0.009356f
C733 B.n693 VSUBS 0.009356f
C734 B.n694 VSUBS 0.009356f
C735 B.n695 VSUBS 0.009356f
C736 B.n696 VSUBS 0.009356f
C737 B.n697 VSUBS 0.009356f
C738 B.n698 VSUBS 0.009356f
C739 B.n699 VSUBS 0.009356f
C740 B.n700 VSUBS 0.009356f
C741 B.n701 VSUBS 0.009356f
C742 B.n702 VSUBS 0.009356f
C743 B.n703 VSUBS 0.009356f
C744 B.n704 VSUBS 0.009356f
C745 B.n705 VSUBS 0.006467f
C746 B.n706 VSUBS 0.009356f
C747 B.n707 VSUBS 0.009356f
C748 B.n708 VSUBS 0.007568f
C749 B.n709 VSUBS 0.009356f
C750 B.n710 VSUBS 0.009356f
C751 B.n711 VSUBS 0.009356f
C752 B.n712 VSUBS 0.009356f
C753 B.n713 VSUBS 0.009356f
C754 B.n714 VSUBS 0.009356f
C755 B.n715 VSUBS 0.009356f
C756 B.n716 VSUBS 0.009356f
C757 B.n717 VSUBS 0.009356f
C758 B.n718 VSUBS 0.009356f
C759 B.n719 VSUBS 0.009356f
C760 B.n720 VSUBS 0.007568f
C761 B.n721 VSUBS 0.021677f
C762 B.n722 VSUBS 0.006467f
C763 B.n723 VSUBS 0.009356f
C764 B.n724 VSUBS 0.009356f
C765 B.n725 VSUBS 0.009356f
C766 B.n726 VSUBS 0.009356f
C767 B.n727 VSUBS 0.009356f
C768 B.n728 VSUBS 0.009356f
C769 B.n729 VSUBS 0.009356f
C770 B.n730 VSUBS 0.009356f
C771 B.n731 VSUBS 0.009356f
C772 B.n732 VSUBS 0.009356f
C773 B.n733 VSUBS 0.009356f
C774 B.n734 VSUBS 0.009356f
C775 B.n735 VSUBS 0.009356f
C776 B.n736 VSUBS 0.009356f
C777 B.n737 VSUBS 0.009356f
C778 B.n738 VSUBS 0.009356f
C779 B.n739 VSUBS 0.009356f
C780 B.n740 VSUBS 0.009356f
C781 B.n741 VSUBS 0.009356f
C782 B.n742 VSUBS 0.009356f
C783 B.n743 VSUBS 0.009356f
C784 B.n744 VSUBS 0.009356f
C785 B.n745 VSUBS 0.009356f
C786 B.n746 VSUBS 0.009356f
C787 B.n747 VSUBS 0.009356f
C788 B.n748 VSUBS 0.009356f
C789 B.n749 VSUBS 0.009356f
C790 B.n750 VSUBS 0.009356f
C791 B.n751 VSUBS 0.009356f
C792 B.n752 VSUBS 0.009356f
C793 B.n753 VSUBS 0.009356f
C794 B.n754 VSUBS 0.009356f
C795 B.n755 VSUBS 0.009356f
C796 B.n756 VSUBS 0.009356f
C797 B.n757 VSUBS 0.009356f
C798 B.n758 VSUBS 0.009356f
C799 B.n759 VSUBS 0.009356f
C800 B.n760 VSUBS 0.009356f
C801 B.n761 VSUBS 0.009356f
C802 B.n762 VSUBS 0.009356f
C803 B.n763 VSUBS 0.009356f
C804 B.n764 VSUBS 0.009356f
C805 B.n765 VSUBS 0.009356f
C806 B.n766 VSUBS 0.009356f
C807 B.n767 VSUBS 0.009356f
C808 B.n768 VSUBS 0.009356f
C809 B.n769 VSUBS 0.009356f
C810 B.n770 VSUBS 0.009356f
C811 B.n771 VSUBS 0.009356f
C812 B.n772 VSUBS 0.009356f
C813 B.n773 VSUBS 0.009356f
C814 B.n774 VSUBS 0.009356f
C815 B.n775 VSUBS 0.009356f
C816 B.n776 VSUBS 0.009356f
C817 B.n777 VSUBS 0.009356f
C818 B.n778 VSUBS 0.009356f
C819 B.n779 VSUBS 0.009356f
C820 B.n780 VSUBS 0.023291f
C821 B.n781 VSUBS 0.023291f
C822 B.n782 VSUBS 0.022664f
C823 B.n783 VSUBS 0.009356f
C824 B.n784 VSUBS 0.009356f
C825 B.n785 VSUBS 0.009356f
C826 B.n786 VSUBS 0.009356f
C827 B.n787 VSUBS 0.009356f
C828 B.n788 VSUBS 0.009356f
C829 B.n789 VSUBS 0.009356f
C830 B.n790 VSUBS 0.009356f
C831 B.n791 VSUBS 0.009356f
C832 B.n792 VSUBS 0.009356f
C833 B.n793 VSUBS 0.009356f
C834 B.n794 VSUBS 0.009356f
C835 B.n795 VSUBS 0.009356f
C836 B.n796 VSUBS 0.009356f
C837 B.n797 VSUBS 0.009356f
C838 B.n798 VSUBS 0.009356f
C839 B.n799 VSUBS 0.009356f
C840 B.n800 VSUBS 0.009356f
C841 B.n801 VSUBS 0.009356f
C842 B.n802 VSUBS 0.009356f
C843 B.n803 VSUBS 0.009356f
C844 B.n804 VSUBS 0.009356f
C845 B.n805 VSUBS 0.009356f
C846 B.n806 VSUBS 0.009356f
C847 B.n807 VSUBS 0.009356f
C848 B.n808 VSUBS 0.009356f
C849 B.n809 VSUBS 0.009356f
C850 B.n810 VSUBS 0.009356f
C851 B.n811 VSUBS 0.009356f
C852 B.n812 VSUBS 0.009356f
C853 B.n813 VSUBS 0.009356f
C854 B.n814 VSUBS 0.009356f
C855 B.n815 VSUBS 0.009356f
C856 B.n816 VSUBS 0.009356f
C857 B.n817 VSUBS 0.009356f
C858 B.n818 VSUBS 0.009356f
C859 B.n819 VSUBS 0.009356f
C860 B.n820 VSUBS 0.009356f
C861 B.n821 VSUBS 0.009356f
C862 B.n822 VSUBS 0.009356f
C863 B.n823 VSUBS 0.009356f
C864 B.n824 VSUBS 0.009356f
C865 B.n825 VSUBS 0.009356f
C866 B.n826 VSUBS 0.009356f
C867 B.n827 VSUBS 0.009356f
C868 B.n828 VSUBS 0.009356f
C869 B.n829 VSUBS 0.009356f
C870 B.n830 VSUBS 0.009356f
C871 B.n831 VSUBS 0.009356f
C872 B.n832 VSUBS 0.009356f
C873 B.n833 VSUBS 0.009356f
C874 B.n834 VSUBS 0.009356f
C875 B.n835 VSUBS 0.009356f
C876 B.n836 VSUBS 0.009356f
C877 B.n837 VSUBS 0.009356f
C878 B.n838 VSUBS 0.009356f
C879 B.n839 VSUBS 0.009356f
C880 B.n840 VSUBS 0.009356f
C881 B.n841 VSUBS 0.009356f
C882 B.n842 VSUBS 0.009356f
C883 B.n843 VSUBS 0.009356f
C884 B.n844 VSUBS 0.009356f
C885 B.n845 VSUBS 0.009356f
C886 B.n846 VSUBS 0.009356f
C887 B.n847 VSUBS 0.009356f
C888 B.n848 VSUBS 0.009356f
C889 B.n849 VSUBS 0.009356f
C890 B.n850 VSUBS 0.009356f
C891 B.n851 VSUBS 0.009356f
C892 B.n852 VSUBS 0.009356f
C893 B.n853 VSUBS 0.009356f
C894 B.n854 VSUBS 0.009356f
C895 B.n855 VSUBS 0.009356f
C896 B.n856 VSUBS 0.009356f
C897 B.n857 VSUBS 0.009356f
C898 B.n858 VSUBS 0.009356f
C899 B.n859 VSUBS 0.009356f
C900 B.n860 VSUBS 0.009356f
C901 B.n861 VSUBS 0.009356f
C902 B.n862 VSUBS 0.009356f
C903 B.n863 VSUBS 0.009356f
C904 B.n864 VSUBS 0.009356f
C905 B.n865 VSUBS 0.009356f
C906 B.n866 VSUBS 0.009356f
C907 B.n867 VSUBS 0.009356f
C908 B.n868 VSUBS 0.009356f
C909 B.n869 VSUBS 0.009356f
C910 B.n870 VSUBS 0.009356f
C911 B.n871 VSUBS 0.009356f
C912 B.n872 VSUBS 0.009356f
C913 B.n873 VSUBS 0.009356f
C914 B.n874 VSUBS 0.009356f
C915 B.n875 VSUBS 0.012209f
C916 B.n876 VSUBS 0.013006f
C917 B.n877 VSUBS 0.025864f
C918 VDD2.n0 VSUBS 0.033122f
C919 VDD2.n1 VSUBS 0.030377f
C920 VDD2.n2 VSUBS 0.016323f
C921 VDD2.n3 VSUBS 0.038582f
C922 VDD2.n4 VSUBS 0.017283f
C923 VDD2.n5 VSUBS 0.030377f
C924 VDD2.n6 VSUBS 0.016323f
C925 VDD2.n7 VSUBS 0.038582f
C926 VDD2.n8 VSUBS 0.016803f
C927 VDD2.n9 VSUBS 0.030377f
C928 VDD2.n10 VSUBS 0.017283f
C929 VDD2.n11 VSUBS 0.038582f
C930 VDD2.n12 VSUBS 0.017283f
C931 VDD2.n13 VSUBS 0.030377f
C932 VDD2.n14 VSUBS 0.016323f
C933 VDD2.n15 VSUBS 0.038582f
C934 VDD2.n16 VSUBS 0.017283f
C935 VDD2.n17 VSUBS 1.41664f
C936 VDD2.n18 VSUBS 0.016323f
C937 VDD2.t9 VSUBS 0.083087f
C938 VDD2.n19 VSUBS 0.231411f
C939 VDD2.n20 VSUBS 0.029024f
C940 VDD2.n21 VSUBS 0.028937f
C941 VDD2.n22 VSUBS 0.038582f
C942 VDD2.n23 VSUBS 0.017283f
C943 VDD2.n24 VSUBS 0.016323f
C944 VDD2.n25 VSUBS 0.030377f
C945 VDD2.n26 VSUBS 0.030377f
C946 VDD2.n27 VSUBS 0.016323f
C947 VDD2.n28 VSUBS 0.017283f
C948 VDD2.n29 VSUBS 0.038582f
C949 VDD2.n30 VSUBS 0.038582f
C950 VDD2.n31 VSUBS 0.017283f
C951 VDD2.n32 VSUBS 0.016323f
C952 VDD2.n33 VSUBS 0.030377f
C953 VDD2.n34 VSUBS 0.030377f
C954 VDD2.n35 VSUBS 0.016323f
C955 VDD2.n36 VSUBS 0.016323f
C956 VDD2.n37 VSUBS 0.017283f
C957 VDD2.n38 VSUBS 0.038582f
C958 VDD2.n39 VSUBS 0.038582f
C959 VDD2.n40 VSUBS 0.038582f
C960 VDD2.n41 VSUBS 0.016803f
C961 VDD2.n42 VSUBS 0.016323f
C962 VDD2.n43 VSUBS 0.030377f
C963 VDD2.n44 VSUBS 0.030377f
C964 VDD2.n45 VSUBS 0.016323f
C965 VDD2.n46 VSUBS 0.017283f
C966 VDD2.n47 VSUBS 0.038582f
C967 VDD2.n48 VSUBS 0.038582f
C968 VDD2.n49 VSUBS 0.017283f
C969 VDD2.n50 VSUBS 0.016323f
C970 VDD2.n51 VSUBS 0.030377f
C971 VDD2.n52 VSUBS 0.030377f
C972 VDD2.n53 VSUBS 0.016323f
C973 VDD2.n54 VSUBS 0.017283f
C974 VDD2.n55 VSUBS 0.038582f
C975 VDD2.n56 VSUBS 0.092532f
C976 VDD2.n57 VSUBS 0.017283f
C977 VDD2.n58 VSUBS 0.016323f
C978 VDD2.n59 VSUBS 0.07146f
C979 VDD2.n60 VSUBS 0.084323f
C980 VDD2.t7 VSUBS 0.274375f
C981 VDD2.t0 VSUBS 0.274375f
C982 VDD2.n61 VSUBS 2.12505f
C983 VDD2.n62 VSUBS 1.19721f
C984 VDD2.t8 VSUBS 0.274375f
C985 VDD2.t4 VSUBS 0.274375f
C986 VDD2.n63 VSUBS 2.15145f
C987 VDD2.n64 VSUBS 3.92914f
C988 VDD2.n65 VSUBS 0.033122f
C989 VDD2.n66 VSUBS 0.030377f
C990 VDD2.n67 VSUBS 0.016323f
C991 VDD2.n68 VSUBS 0.038582f
C992 VDD2.n69 VSUBS 0.017283f
C993 VDD2.n70 VSUBS 0.030377f
C994 VDD2.n71 VSUBS 0.016323f
C995 VDD2.n72 VSUBS 0.038582f
C996 VDD2.n73 VSUBS 0.016803f
C997 VDD2.n74 VSUBS 0.030377f
C998 VDD2.n75 VSUBS 0.016803f
C999 VDD2.n76 VSUBS 0.016323f
C1000 VDD2.n77 VSUBS 0.038582f
C1001 VDD2.n78 VSUBS 0.038582f
C1002 VDD2.n79 VSUBS 0.017283f
C1003 VDD2.n80 VSUBS 0.030377f
C1004 VDD2.n81 VSUBS 0.016323f
C1005 VDD2.n82 VSUBS 0.038582f
C1006 VDD2.n83 VSUBS 0.017283f
C1007 VDD2.n84 VSUBS 1.41664f
C1008 VDD2.n85 VSUBS 0.016323f
C1009 VDD2.t1 VSUBS 0.083087f
C1010 VDD2.n86 VSUBS 0.231411f
C1011 VDD2.n87 VSUBS 0.029024f
C1012 VDD2.n88 VSUBS 0.028937f
C1013 VDD2.n89 VSUBS 0.038582f
C1014 VDD2.n90 VSUBS 0.017283f
C1015 VDD2.n91 VSUBS 0.016323f
C1016 VDD2.n92 VSUBS 0.030377f
C1017 VDD2.n93 VSUBS 0.030377f
C1018 VDD2.n94 VSUBS 0.016323f
C1019 VDD2.n95 VSUBS 0.017283f
C1020 VDD2.n96 VSUBS 0.038582f
C1021 VDD2.n97 VSUBS 0.038582f
C1022 VDD2.n98 VSUBS 0.017283f
C1023 VDD2.n99 VSUBS 0.016323f
C1024 VDD2.n100 VSUBS 0.030377f
C1025 VDD2.n101 VSUBS 0.030377f
C1026 VDD2.n102 VSUBS 0.016323f
C1027 VDD2.n103 VSUBS 0.017283f
C1028 VDD2.n104 VSUBS 0.038582f
C1029 VDD2.n105 VSUBS 0.038582f
C1030 VDD2.n106 VSUBS 0.017283f
C1031 VDD2.n107 VSUBS 0.016323f
C1032 VDD2.n108 VSUBS 0.030377f
C1033 VDD2.n109 VSUBS 0.030377f
C1034 VDD2.n110 VSUBS 0.016323f
C1035 VDD2.n111 VSUBS 0.017283f
C1036 VDD2.n112 VSUBS 0.038582f
C1037 VDD2.n113 VSUBS 0.038582f
C1038 VDD2.n114 VSUBS 0.017283f
C1039 VDD2.n115 VSUBS 0.016323f
C1040 VDD2.n116 VSUBS 0.030377f
C1041 VDD2.n117 VSUBS 0.030377f
C1042 VDD2.n118 VSUBS 0.016323f
C1043 VDD2.n119 VSUBS 0.017283f
C1044 VDD2.n120 VSUBS 0.038582f
C1045 VDD2.n121 VSUBS 0.092532f
C1046 VDD2.n122 VSUBS 0.017283f
C1047 VDD2.n123 VSUBS 0.016323f
C1048 VDD2.n124 VSUBS 0.07146f
C1049 VDD2.n125 VSUBS 0.067498f
C1050 VDD2.n126 VSUBS 3.55859f
C1051 VDD2.t2 VSUBS 0.274375f
C1052 VDD2.t3 VSUBS 0.274375f
C1053 VDD2.n127 VSUBS 2.12506f
C1054 VDD2.n128 VSUBS 0.89984f
C1055 VDD2.t5 VSUBS 0.274375f
C1056 VDD2.t6 VSUBS 0.274375f
C1057 VDD2.n129 VSUBS 2.15139f
C1058 VN.n0 VSUBS 0.03623f
C1059 VN.t5 VSUBS 2.40135f
C1060 VN.n1 VSUBS 0.055407f
C1061 VN.n2 VSUBS 0.02748f
C1062 VN.n3 VSUBS 0.031493f
C1063 VN.n4 VSUBS 0.02748f
C1064 VN.n5 VSUBS 0.045476f
C1065 VN.n6 VSUBS 0.02748f
C1066 VN.t9 VSUBS 2.40135f
C1067 VN.n7 VSUBS 0.051216f
C1068 VN.n8 VSUBS 0.02748f
C1069 VN.n9 VSUBS 0.045653f
C1070 VN.t0 VSUBS 2.6593f
C1071 VN.t2 VSUBS 2.40135f
C1072 VN.n10 VSUBS 0.941646f
C1073 VN.n11 VSUBS 0.904731f
C1074 VN.n12 VSUBS 0.28875f
C1075 VN.n13 VSUBS 0.02748f
C1076 VN.n14 VSUBS 0.051216f
C1077 VN.n15 VSUBS 0.034756f
C1078 VN.n16 VSUBS 0.045476f
C1079 VN.n17 VSUBS 0.02748f
C1080 VN.n18 VSUBS 0.02748f
C1081 VN.n19 VSUBS 0.02748f
C1082 VN.n20 VSUBS 0.038573f
C1083 VN.n21 VSUBS 0.849781f
C1084 VN.n22 VSUBS 0.038573f
C1085 VN.n23 VSUBS 0.051216f
C1086 VN.n24 VSUBS 0.02748f
C1087 VN.n25 VSUBS 0.02748f
C1088 VN.n26 VSUBS 0.02748f
C1089 VN.n27 VSUBS 0.034756f
C1090 VN.n28 VSUBS 0.051216f
C1091 VN.t1 VSUBS 2.40135f
C1092 VN.n29 VSUBS 0.849781f
C1093 VN.n30 VSUBS 0.045653f
C1094 VN.n31 VSUBS 0.02748f
C1095 VN.n32 VSUBS 0.02748f
C1096 VN.n33 VSUBS 0.02748f
C1097 VN.n34 VSUBS 0.051216f
C1098 VN.n35 VSUBS 0.053256f
C1099 VN.n36 VSUBS 0.022785f
C1100 VN.n37 VSUBS 0.02748f
C1101 VN.n38 VSUBS 0.02748f
C1102 VN.n39 VSUBS 0.02748f
C1103 VN.n40 VSUBS 0.051216f
C1104 VN.n41 VSUBS 0.027447f
C1105 VN.n42 VSUBS 0.936961f
C1106 VN.n43 VSUBS 0.052166f
C1107 VN.n44 VSUBS 0.03623f
C1108 VN.t8 VSUBS 2.40135f
C1109 VN.n45 VSUBS 0.055407f
C1110 VN.n46 VSUBS 0.02748f
C1111 VN.n47 VSUBS 0.031493f
C1112 VN.n48 VSUBS 0.02748f
C1113 VN.t7 VSUBS 2.40135f
C1114 VN.n49 VSUBS 0.849781f
C1115 VN.n50 VSUBS 0.045476f
C1116 VN.n51 VSUBS 0.02748f
C1117 VN.t6 VSUBS 2.40135f
C1118 VN.n52 VSUBS 0.051216f
C1119 VN.n53 VSUBS 0.02748f
C1120 VN.n54 VSUBS 0.045653f
C1121 VN.t3 VSUBS 2.6593f
C1122 VN.t4 VSUBS 2.40135f
C1123 VN.n55 VSUBS 0.941646f
C1124 VN.n56 VSUBS 0.904731f
C1125 VN.n57 VSUBS 0.28875f
C1126 VN.n58 VSUBS 0.02748f
C1127 VN.n59 VSUBS 0.051216f
C1128 VN.n60 VSUBS 0.034756f
C1129 VN.n61 VSUBS 0.045476f
C1130 VN.n62 VSUBS 0.02748f
C1131 VN.n63 VSUBS 0.02748f
C1132 VN.n64 VSUBS 0.02748f
C1133 VN.n65 VSUBS 0.038573f
C1134 VN.n66 VSUBS 0.849781f
C1135 VN.n67 VSUBS 0.038573f
C1136 VN.n68 VSUBS 0.051216f
C1137 VN.n69 VSUBS 0.02748f
C1138 VN.n70 VSUBS 0.02748f
C1139 VN.n71 VSUBS 0.02748f
C1140 VN.n72 VSUBS 0.034756f
C1141 VN.n73 VSUBS 0.051216f
C1142 VN.n74 VSUBS 0.045653f
C1143 VN.n75 VSUBS 0.02748f
C1144 VN.n76 VSUBS 0.02748f
C1145 VN.n77 VSUBS 0.02748f
C1146 VN.n78 VSUBS 0.051216f
C1147 VN.n79 VSUBS 0.053256f
C1148 VN.n80 VSUBS 0.022785f
C1149 VN.n81 VSUBS 0.02748f
C1150 VN.n82 VSUBS 0.02748f
C1151 VN.n83 VSUBS 0.02748f
C1152 VN.n84 VSUBS 0.051216f
C1153 VN.n85 VSUBS 0.027447f
C1154 VN.n86 VSUBS 0.936961f
C1155 VN.n87 VSUBS 1.71975f
C1156 VDD1.n0 VSUBS 0.033224f
C1157 VDD1.n1 VSUBS 0.030471f
C1158 VDD1.n2 VSUBS 0.016374f
C1159 VDD1.n3 VSUBS 0.038701f
C1160 VDD1.n4 VSUBS 0.017337f
C1161 VDD1.n5 VSUBS 0.030471f
C1162 VDD1.n6 VSUBS 0.016374f
C1163 VDD1.n7 VSUBS 0.038701f
C1164 VDD1.n8 VSUBS 0.016855f
C1165 VDD1.n9 VSUBS 0.030471f
C1166 VDD1.n10 VSUBS 0.016855f
C1167 VDD1.n11 VSUBS 0.016374f
C1168 VDD1.n12 VSUBS 0.038701f
C1169 VDD1.n13 VSUBS 0.038701f
C1170 VDD1.n14 VSUBS 0.017337f
C1171 VDD1.n15 VSUBS 0.030471f
C1172 VDD1.n16 VSUBS 0.016374f
C1173 VDD1.n17 VSUBS 0.038701f
C1174 VDD1.n18 VSUBS 0.017337f
C1175 VDD1.n19 VSUBS 1.421f
C1176 VDD1.n20 VSUBS 0.016374f
C1177 VDD1.t2 VSUBS 0.083343f
C1178 VDD1.n21 VSUBS 0.232124f
C1179 VDD1.n22 VSUBS 0.029113f
C1180 VDD1.n23 VSUBS 0.029026f
C1181 VDD1.n24 VSUBS 0.038701f
C1182 VDD1.n25 VSUBS 0.017337f
C1183 VDD1.n26 VSUBS 0.016374f
C1184 VDD1.n27 VSUBS 0.030471f
C1185 VDD1.n28 VSUBS 0.030471f
C1186 VDD1.n29 VSUBS 0.016374f
C1187 VDD1.n30 VSUBS 0.017337f
C1188 VDD1.n31 VSUBS 0.038701f
C1189 VDD1.n32 VSUBS 0.038701f
C1190 VDD1.n33 VSUBS 0.017337f
C1191 VDD1.n34 VSUBS 0.016374f
C1192 VDD1.n35 VSUBS 0.030471f
C1193 VDD1.n36 VSUBS 0.030471f
C1194 VDD1.n37 VSUBS 0.016374f
C1195 VDD1.n38 VSUBS 0.017337f
C1196 VDD1.n39 VSUBS 0.038701f
C1197 VDD1.n40 VSUBS 0.038701f
C1198 VDD1.n41 VSUBS 0.017337f
C1199 VDD1.n42 VSUBS 0.016374f
C1200 VDD1.n43 VSUBS 0.030471f
C1201 VDD1.n44 VSUBS 0.030471f
C1202 VDD1.n45 VSUBS 0.016374f
C1203 VDD1.n46 VSUBS 0.017337f
C1204 VDD1.n47 VSUBS 0.038701f
C1205 VDD1.n48 VSUBS 0.038701f
C1206 VDD1.n49 VSUBS 0.017337f
C1207 VDD1.n50 VSUBS 0.016374f
C1208 VDD1.n51 VSUBS 0.030471f
C1209 VDD1.n52 VSUBS 0.030471f
C1210 VDD1.n53 VSUBS 0.016374f
C1211 VDD1.n54 VSUBS 0.017337f
C1212 VDD1.n55 VSUBS 0.038701f
C1213 VDD1.n56 VSUBS 0.092817f
C1214 VDD1.n57 VSUBS 0.017337f
C1215 VDD1.n58 VSUBS 0.016374f
C1216 VDD1.n59 VSUBS 0.07168f
C1217 VDD1.n60 VSUBS 0.084582f
C1218 VDD1.t3 VSUBS 0.275219f
C1219 VDD1.t9 VSUBS 0.275219f
C1220 VDD1.n61 VSUBS 2.1316f
C1221 VDD1.n62 VSUBS 1.21089f
C1222 VDD1.n63 VSUBS 0.033224f
C1223 VDD1.n64 VSUBS 0.030471f
C1224 VDD1.n65 VSUBS 0.016374f
C1225 VDD1.n66 VSUBS 0.038701f
C1226 VDD1.n67 VSUBS 0.017337f
C1227 VDD1.n68 VSUBS 0.030471f
C1228 VDD1.n69 VSUBS 0.016374f
C1229 VDD1.n70 VSUBS 0.038701f
C1230 VDD1.n71 VSUBS 0.016855f
C1231 VDD1.n72 VSUBS 0.030471f
C1232 VDD1.n73 VSUBS 0.017337f
C1233 VDD1.n74 VSUBS 0.038701f
C1234 VDD1.n75 VSUBS 0.017337f
C1235 VDD1.n76 VSUBS 0.030471f
C1236 VDD1.n77 VSUBS 0.016374f
C1237 VDD1.n78 VSUBS 0.038701f
C1238 VDD1.n79 VSUBS 0.017337f
C1239 VDD1.n80 VSUBS 1.421f
C1240 VDD1.n81 VSUBS 0.016374f
C1241 VDD1.t6 VSUBS 0.083343f
C1242 VDD1.n82 VSUBS 0.232124f
C1243 VDD1.n83 VSUBS 0.029113f
C1244 VDD1.n84 VSUBS 0.029026f
C1245 VDD1.n85 VSUBS 0.038701f
C1246 VDD1.n86 VSUBS 0.017337f
C1247 VDD1.n87 VSUBS 0.016374f
C1248 VDD1.n88 VSUBS 0.030471f
C1249 VDD1.n89 VSUBS 0.030471f
C1250 VDD1.n90 VSUBS 0.016374f
C1251 VDD1.n91 VSUBS 0.017337f
C1252 VDD1.n92 VSUBS 0.038701f
C1253 VDD1.n93 VSUBS 0.038701f
C1254 VDD1.n94 VSUBS 0.017337f
C1255 VDD1.n95 VSUBS 0.016374f
C1256 VDD1.n96 VSUBS 0.030471f
C1257 VDD1.n97 VSUBS 0.030471f
C1258 VDD1.n98 VSUBS 0.016374f
C1259 VDD1.n99 VSUBS 0.016374f
C1260 VDD1.n100 VSUBS 0.017337f
C1261 VDD1.n101 VSUBS 0.038701f
C1262 VDD1.n102 VSUBS 0.038701f
C1263 VDD1.n103 VSUBS 0.038701f
C1264 VDD1.n104 VSUBS 0.016855f
C1265 VDD1.n105 VSUBS 0.016374f
C1266 VDD1.n106 VSUBS 0.030471f
C1267 VDD1.n107 VSUBS 0.030471f
C1268 VDD1.n108 VSUBS 0.016374f
C1269 VDD1.n109 VSUBS 0.017337f
C1270 VDD1.n110 VSUBS 0.038701f
C1271 VDD1.n111 VSUBS 0.038701f
C1272 VDD1.n112 VSUBS 0.017337f
C1273 VDD1.n113 VSUBS 0.016374f
C1274 VDD1.n114 VSUBS 0.030471f
C1275 VDD1.n115 VSUBS 0.030471f
C1276 VDD1.n116 VSUBS 0.016374f
C1277 VDD1.n117 VSUBS 0.017337f
C1278 VDD1.n118 VSUBS 0.038701f
C1279 VDD1.n119 VSUBS 0.092817f
C1280 VDD1.n120 VSUBS 0.017337f
C1281 VDD1.n121 VSUBS 0.016374f
C1282 VDD1.n122 VSUBS 0.07168f
C1283 VDD1.n123 VSUBS 0.084582f
C1284 VDD1.t8 VSUBS 0.275219f
C1285 VDD1.t5 VSUBS 0.275219f
C1286 VDD1.n124 VSUBS 2.13159f
C1287 VDD1.n125 VSUBS 1.20089f
C1288 VDD1.t7 VSUBS 0.275219f
C1289 VDD1.t1 VSUBS 0.275219f
C1290 VDD1.n126 VSUBS 2.15807f
C1291 VDD1.n127 VSUBS 4.10009f
C1292 VDD1.t4 VSUBS 0.275219f
C1293 VDD1.t0 VSUBS 0.275219f
C1294 VDD1.n128 VSUBS 2.13159f
C1295 VDD1.n129 VSUBS 4.23444f
C1296 VTAIL.t2 VSUBS 0.26529f
C1297 VTAIL.t16 VSUBS 0.26529f
C1298 VTAIL.n0 VSUBS 1.90158f
C1299 VTAIL.n1 VSUBS 1.02771f
C1300 VTAIL.n2 VSUBS 0.032025f
C1301 VTAIL.n3 VSUBS 0.029371f
C1302 VTAIL.n4 VSUBS 0.015783f
C1303 VTAIL.n5 VSUBS 0.037305f
C1304 VTAIL.n6 VSUBS 0.016711f
C1305 VTAIL.n7 VSUBS 0.029371f
C1306 VTAIL.n8 VSUBS 0.015783f
C1307 VTAIL.n9 VSUBS 0.037305f
C1308 VTAIL.n10 VSUBS 0.016247f
C1309 VTAIL.n11 VSUBS 0.029371f
C1310 VTAIL.n12 VSUBS 0.016711f
C1311 VTAIL.n13 VSUBS 0.037305f
C1312 VTAIL.n14 VSUBS 0.016711f
C1313 VTAIL.n15 VSUBS 0.029371f
C1314 VTAIL.n16 VSUBS 0.015783f
C1315 VTAIL.n17 VSUBS 0.037305f
C1316 VTAIL.n18 VSUBS 0.016711f
C1317 VTAIL.n19 VSUBS 1.36973f
C1318 VTAIL.n20 VSUBS 0.015783f
C1319 VTAIL.t7 VSUBS 0.080336f
C1320 VTAIL.n21 VSUBS 0.223749f
C1321 VTAIL.n22 VSUBS 0.028063f
C1322 VTAIL.n23 VSUBS 0.027979f
C1323 VTAIL.n24 VSUBS 0.037305f
C1324 VTAIL.n25 VSUBS 0.016711f
C1325 VTAIL.n26 VSUBS 0.015783f
C1326 VTAIL.n27 VSUBS 0.029371f
C1327 VTAIL.n28 VSUBS 0.029371f
C1328 VTAIL.n29 VSUBS 0.015783f
C1329 VTAIL.n30 VSUBS 0.016711f
C1330 VTAIL.n31 VSUBS 0.037305f
C1331 VTAIL.n32 VSUBS 0.037305f
C1332 VTAIL.n33 VSUBS 0.016711f
C1333 VTAIL.n34 VSUBS 0.015783f
C1334 VTAIL.n35 VSUBS 0.029371f
C1335 VTAIL.n36 VSUBS 0.029371f
C1336 VTAIL.n37 VSUBS 0.015783f
C1337 VTAIL.n38 VSUBS 0.015783f
C1338 VTAIL.n39 VSUBS 0.016711f
C1339 VTAIL.n40 VSUBS 0.037305f
C1340 VTAIL.n41 VSUBS 0.037305f
C1341 VTAIL.n42 VSUBS 0.037305f
C1342 VTAIL.n43 VSUBS 0.016247f
C1343 VTAIL.n44 VSUBS 0.015783f
C1344 VTAIL.n45 VSUBS 0.029371f
C1345 VTAIL.n46 VSUBS 0.029371f
C1346 VTAIL.n47 VSUBS 0.015783f
C1347 VTAIL.n48 VSUBS 0.016711f
C1348 VTAIL.n49 VSUBS 0.037305f
C1349 VTAIL.n50 VSUBS 0.037305f
C1350 VTAIL.n51 VSUBS 0.016711f
C1351 VTAIL.n52 VSUBS 0.015783f
C1352 VTAIL.n53 VSUBS 0.029371f
C1353 VTAIL.n54 VSUBS 0.029371f
C1354 VTAIL.n55 VSUBS 0.015783f
C1355 VTAIL.n56 VSUBS 0.016711f
C1356 VTAIL.n57 VSUBS 0.037305f
C1357 VTAIL.n58 VSUBS 0.089468f
C1358 VTAIL.n59 VSUBS 0.016711f
C1359 VTAIL.n60 VSUBS 0.015783f
C1360 VTAIL.n61 VSUBS 0.069094f
C1361 VTAIL.n62 VSUBS 0.044992f
C1362 VTAIL.n63 VSUBS 0.454502f
C1363 VTAIL.t5 VSUBS 0.26529f
C1364 VTAIL.t14 VSUBS 0.26529f
C1365 VTAIL.n64 VSUBS 1.90158f
C1366 VTAIL.n65 VSUBS 1.16987f
C1367 VTAIL.t9 VSUBS 0.26529f
C1368 VTAIL.t10 VSUBS 0.26529f
C1369 VTAIL.n66 VSUBS 1.90158f
C1370 VTAIL.n67 VSUBS 2.75756f
C1371 VTAIL.t19 VSUBS 0.26529f
C1372 VTAIL.t18 VSUBS 0.26529f
C1373 VTAIL.n68 VSUBS 1.90159f
C1374 VTAIL.n69 VSUBS 2.75755f
C1375 VTAIL.t0 VSUBS 0.26529f
C1376 VTAIL.t3 VSUBS 0.26529f
C1377 VTAIL.n70 VSUBS 1.90159f
C1378 VTAIL.n71 VSUBS 1.16986f
C1379 VTAIL.n72 VSUBS 0.032025f
C1380 VTAIL.n73 VSUBS 0.029371f
C1381 VTAIL.n74 VSUBS 0.015783f
C1382 VTAIL.n75 VSUBS 0.037305f
C1383 VTAIL.n76 VSUBS 0.016711f
C1384 VTAIL.n77 VSUBS 0.029371f
C1385 VTAIL.n78 VSUBS 0.015783f
C1386 VTAIL.n79 VSUBS 0.037305f
C1387 VTAIL.n80 VSUBS 0.016247f
C1388 VTAIL.n81 VSUBS 0.029371f
C1389 VTAIL.n82 VSUBS 0.016247f
C1390 VTAIL.n83 VSUBS 0.015783f
C1391 VTAIL.n84 VSUBS 0.037305f
C1392 VTAIL.n85 VSUBS 0.037305f
C1393 VTAIL.n86 VSUBS 0.016711f
C1394 VTAIL.n87 VSUBS 0.029371f
C1395 VTAIL.n88 VSUBS 0.015783f
C1396 VTAIL.n89 VSUBS 0.037305f
C1397 VTAIL.n90 VSUBS 0.016711f
C1398 VTAIL.n91 VSUBS 1.36973f
C1399 VTAIL.n92 VSUBS 0.015783f
C1400 VTAIL.t15 VSUBS 0.080336f
C1401 VTAIL.n93 VSUBS 0.223749f
C1402 VTAIL.n94 VSUBS 0.028063f
C1403 VTAIL.n95 VSUBS 0.027979f
C1404 VTAIL.n96 VSUBS 0.037305f
C1405 VTAIL.n97 VSUBS 0.016711f
C1406 VTAIL.n98 VSUBS 0.015783f
C1407 VTAIL.n99 VSUBS 0.029371f
C1408 VTAIL.n100 VSUBS 0.029371f
C1409 VTAIL.n101 VSUBS 0.015783f
C1410 VTAIL.n102 VSUBS 0.016711f
C1411 VTAIL.n103 VSUBS 0.037305f
C1412 VTAIL.n104 VSUBS 0.037305f
C1413 VTAIL.n105 VSUBS 0.016711f
C1414 VTAIL.n106 VSUBS 0.015783f
C1415 VTAIL.n107 VSUBS 0.029371f
C1416 VTAIL.n108 VSUBS 0.029371f
C1417 VTAIL.n109 VSUBS 0.015783f
C1418 VTAIL.n110 VSUBS 0.016711f
C1419 VTAIL.n111 VSUBS 0.037305f
C1420 VTAIL.n112 VSUBS 0.037305f
C1421 VTAIL.n113 VSUBS 0.016711f
C1422 VTAIL.n114 VSUBS 0.015783f
C1423 VTAIL.n115 VSUBS 0.029371f
C1424 VTAIL.n116 VSUBS 0.029371f
C1425 VTAIL.n117 VSUBS 0.015783f
C1426 VTAIL.n118 VSUBS 0.016711f
C1427 VTAIL.n119 VSUBS 0.037305f
C1428 VTAIL.n120 VSUBS 0.037305f
C1429 VTAIL.n121 VSUBS 0.016711f
C1430 VTAIL.n122 VSUBS 0.015783f
C1431 VTAIL.n123 VSUBS 0.029371f
C1432 VTAIL.n124 VSUBS 0.029371f
C1433 VTAIL.n125 VSUBS 0.015783f
C1434 VTAIL.n126 VSUBS 0.016711f
C1435 VTAIL.n127 VSUBS 0.037305f
C1436 VTAIL.n128 VSUBS 0.089468f
C1437 VTAIL.n129 VSUBS 0.016711f
C1438 VTAIL.n130 VSUBS 0.015783f
C1439 VTAIL.n131 VSUBS 0.069094f
C1440 VTAIL.n132 VSUBS 0.044992f
C1441 VTAIL.n133 VSUBS 0.454502f
C1442 VTAIL.t13 VSUBS 0.26529f
C1443 VTAIL.t8 VSUBS 0.26529f
C1444 VTAIL.n134 VSUBS 1.90159f
C1445 VTAIL.n135 VSUBS 1.08623f
C1446 VTAIL.t11 VSUBS 0.26529f
C1447 VTAIL.t6 VSUBS 0.26529f
C1448 VTAIL.n136 VSUBS 1.90159f
C1449 VTAIL.n137 VSUBS 1.16986f
C1450 VTAIL.n138 VSUBS 0.032025f
C1451 VTAIL.n139 VSUBS 0.029371f
C1452 VTAIL.n140 VSUBS 0.015783f
C1453 VTAIL.n141 VSUBS 0.037305f
C1454 VTAIL.n142 VSUBS 0.016711f
C1455 VTAIL.n143 VSUBS 0.029371f
C1456 VTAIL.n144 VSUBS 0.015783f
C1457 VTAIL.n145 VSUBS 0.037305f
C1458 VTAIL.n146 VSUBS 0.016247f
C1459 VTAIL.n147 VSUBS 0.029371f
C1460 VTAIL.n148 VSUBS 0.016247f
C1461 VTAIL.n149 VSUBS 0.015783f
C1462 VTAIL.n150 VSUBS 0.037305f
C1463 VTAIL.n151 VSUBS 0.037305f
C1464 VTAIL.n152 VSUBS 0.016711f
C1465 VTAIL.n153 VSUBS 0.029371f
C1466 VTAIL.n154 VSUBS 0.015783f
C1467 VTAIL.n155 VSUBS 0.037305f
C1468 VTAIL.n156 VSUBS 0.016711f
C1469 VTAIL.n157 VSUBS 1.36973f
C1470 VTAIL.n158 VSUBS 0.015783f
C1471 VTAIL.t12 VSUBS 0.080336f
C1472 VTAIL.n159 VSUBS 0.223749f
C1473 VTAIL.n160 VSUBS 0.028063f
C1474 VTAIL.n161 VSUBS 0.027979f
C1475 VTAIL.n162 VSUBS 0.037305f
C1476 VTAIL.n163 VSUBS 0.016711f
C1477 VTAIL.n164 VSUBS 0.015783f
C1478 VTAIL.n165 VSUBS 0.029371f
C1479 VTAIL.n166 VSUBS 0.029371f
C1480 VTAIL.n167 VSUBS 0.015783f
C1481 VTAIL.n168 VSUBS 0.016711f
C1482 VTAIL.n169 VSUBS 0.037305f
C1483 VTAIL.n170 VSUBS 0.037305f
C1484 VTAIL.n171 VSUBS 0.016711f
C1485 VTAIL.n172 VSUBS 0.015783f
C1486 VTAIL.n173 VSUBS 0.029371f
C1487 VTAIL.n174 VSUBS 0.029371f
C1488 VTAIL.n175 VSUBS 0.015783f
C1489 VTAIL.n176 VSUBS 0.016711f
C1490 VTAIL.n177 VSUBS 0.037305f
C1491 VTAIL.n178 VSUBS 0.037305f
C1492 VTAIL.n179 VSUBS 0.016711f
C1493 VTAIL.n180 VSUBS 0.015783f
C1494 VTAIL.n181 VSUBS 0.029371f
C1495 VTAIL.n182 VSUBS 0.029371f
C1496 VTAIL.n183 VSUBS 0.015783f
C1497 VTAIL.n184 VSUBS 0.016711f
C1498 VTAIL.n185 VSUBS 0.037305f
C1499 VTAIL.n186 VSUBS 0.037305f
C1500 VTAIL.n187 VSUBS 0.016711f
C1501 VTAIL.n188 VSUBS 0.015783f
C1502 VTAIL.n189 VSUBS 0.029371f
C1503 VTAIL.n190 VSUBS 0.029371f
C1504 VTAIL.n191 VSUBS 0.015783f
C1505 VTAIL.n192 VSUBS 0.016711f
C1506 VTAIL.n193 VSUBS 0.037305f
C1507 VTAIL.n194 VSUBS 0.089468f
C1508 VTAIL.n195 VSUBS 0.016711f
C1509 VTAIL.n196 VSUBS 0.015783f
C1510 VTAIL.n197 VSUBS 0.069094f
C1511 VTAIL.n198 VSUBS 0.044992f
C1512 VTAIL.n199 VSUBS 1.86963f
C1513 VTAIL.n200 VSUBS 0.032025f
C1514 VTAIL.n201 VSUBS 0.029371f
C1515 VTAIL.n202 VSUBS 0.015783f
C1516 VTAIL.n203 VSUBS 0.037305f
C1517 VTAIL.n204 VSUBS 0.016711f
C1518 VTAIL.n205 VSUBS 0.029371f
C1519 VTAIL.n206 VSUBS 0.015783f
C1520 VTAIL.n207 VSUBS 0.037305f
C1521 VTAIL.n208 VSUBS 0.016247f
C1522 VTAIL.n209 VSUBS 0.029371f
C1523 VTAIL.n210 VSUBS 0.016711f
C1524 VTAIL.n211 VSUBS 0.037305f
C1525 VTAIL.n212 VSUBS 0.016711f
C1526 VTAIL.n213 VSUBS 0.029371f
C1527 VTAIL.n214 VSUBS 0.015783f
C1528 VTAIL.n215 VSUBS 0.037305f
C1529 VTAIL.n216 VSUBS 0.016711f
C1530 VTAIL.n217 VSUBS 1.36973f
C1531 VTAIL.n218 VSUBS 0.015783f
C1532 VTAIL.t4 VSUBS 0.080336f
C1533 VTAIL.n219 VSUBS 0.223749f
C1534 VTAIL.n220 VSUBS 0.028063f
C1535 VTAIL.n221 VSUBS 0.027979f
C1536 VTAIL.n222 VSUBS 0.037305f
C1537 VTAIL.n223 VSUBS 0.016711f
C1538 VTAIL.n224 VSUBS 0.015783f
C1539 VTAIL.n225 VSUBS 0.029371f
C1540 VTAIL.n226 VSUBS 0.029371f
C1541 VTAIL.n227 VSUBS 0.015783f
C1542 VTAIL.n228 VSUBS 0.016711f
C1543 VTAIL.n229 VSUBS 0.037305f
C1544 VTAIL.n230 VSUBS 0.037305f
C1545 VTAIL.n231 VSUBS 0.016711f
C1546 VTAIL.n232 VSUBS 0.015783f
C1547 VTAIL.n233 VSUBS 0.029371f
C1548 VTAIL.n234 VSUBS 0.029371f
C1549 VTAIL.n235 VSUBS 0.015783f
C1550 VTAIL.n236 VSUBS 0.015783f
C1551 VTAIL.n237 VSUBS 0.016711f
C1552 VTAIL.n238 VSUBS 0.037305f
C1553 VTAIL.n239 VSUBS 0.037305f
C1554 VTAIL.n240 VSUBS 0.037305f
C1555 VTAIL.n241 VSUBS 0.016247f
C1556 VTAIL.n242 VSUBS 0.015783f
C1557 VTAIL.n243 VSUBS 0.029371f
C1558 VTAIL.n244 VSUBS 0.029371f
C1559 VTAIL.n245 VSUBS 0.015783f
C1560 VTAIL.n246 VSUBS 0.016711f
C1561 VTAIL.n247 VSUBS 0.037305f
C1562 VTAIL.n248 VSUBS 0.037305f
C1563 VTAIL.n249 VSUBS 0.016711f
C1564 VTAIL.n250 VSUBS 0.015783f
C1565 VTAIL.n251 VSUBS 0.029371f
C1566 VTAIL.n252 VSUBS 0.029371f
C1567 VTAIL.n253 VSUBS 0.015783f
C1568 VTAIL.n254 VSUBS 0.016711f
C1569 VTAIL.n255 VSUBS 0.037305f
C1570 VTAIL.n256 VSUBS 0.089468f
C1571 VTAIL.n257 VSUBS 0.016711f
C1572 VTAIL.n258 VSUBS 0.015783f
C1573 VTAIL.n259 VSUBS 0.069094f
C1574 VTAIL.n260 VSUBS 0.044992f
C1575 VTAIL.n261 VSUBS 1.86963f
C1576 VTAIL.t17 VSUBS 0.26529f
C1577 VTAIL.t1 VSUBS 0.26529f
C1578 VTAIL.n262 VSUBS 1.90158f
C1579 VTAIL.n263 VSUBS 0.972231f
C1580 VP.n0 VSUBS 0.039422f
C1581 VP.t8 VSUBS 2.61294f
C1582 VP.n1 VSUBS 0.060289f
C1583 VP.n2 VSUBS 0.029901f
C1584 VP.n3 VSUBS 0.034268f
C1585 VP.n4 VSUBS 0.029901f
C1586 VP.n5 VSUBS 0.049483f
C1587 VP.n6 VSUBS 0.029901f
C1588 VP.t4 VSUBS 2.61294f
C1589 VP.n7 VSUBS 0.055728f
C1590 VP.n8 VSUBS 0.029901f
C1591 VP.n9 VSUBS 0.049675f
C1592 VP.n10 VSUBS 0.029901f
C1593 VP.n11 VSUBS 0.024792f
C1594 VP.n12 VSUBS 0.029901f
C1595 VP.t3 VSUBS 2.61294f
C1596 VP.n13 VSUBS 1.01952f
C1597 VP.n14 VSUBS 0.039422f
C1598 VP.t9 VSUBS 2.61294f
C1599 VP.n15 VSUBS 0.060289f
C1600 VP.n16 VSUBS 0.029901f
C1601 VP.n17 VSUBS 0.034268f
C1602 VP.n18 VSUBS 0.029901f
C1603 VP.n19 VSUBS 0.049483f
C1604 VP.n20 VSUBS 0.029901f
C1605 VP.t0 VSUBS 2.61294f
C1606 VP.n21 VSUBS 0.055728f
C1607 VP.n22 VSUBS 0.029901f
C1608 VP.n23 VSUBS 0.049675f
C1609 VP.t7 VSUBS 2.89361f
C1610 VP.t6 VSUBS 2.61294f
C1611 VP.n24 VSUBS 1.02461f
C1612 VP.n25 VSUBS 0.984447f
C1613 VP.n26 VSUBS 0.314192f
C1614 VP.n27 VSUBS 0.029901f
C1615 VP.n28 VSUBS 0.055728f
C1616 VP.n29 VSUBS 0.037818f
C1617 VP.n30 VSUBS 0.049483f
C1618 VP.n31 VSUBS 0.029901f
C1619 VP.n32 VSUBS 0.029901f
C1620 VP.n33 VSUBS 0.029901f
C1621 VP.n34 VSUBS 0.041972f
C1622 VP.n35 VSUBS 0.924656f
C1623 VP.n36 VSUBS 0.041972f
C1624 VP.n37 VSUBS 0.055728f
C1625 VP.n38 VSUBS 0.029901f
C1626 VP.n39 VSUBS 0.029901f
C1627 VP.n40 VSUBS 0.029901f
C1628 VP.n41 VSUBS 0.037818f
C1629 VP.n42 VSUBS 0.055728f
C1630 VP.t5 VSUBS 2.61294f
C1631 VP.n43 VSUBS 0.924656f
C1632 VP.n44 VSUBS 0.049675f
C1633 VP.n45 VSUBS 0.029901f
C1634 VP.n46 VSUBS 0.029901f
C1635 VP.n47 VSUBS 0.029901f
C1636 VP.n48 VSUBS 0.055728f
C1637 VP.n49 VSUBS 0.057948f
C1638 VP.n50 VSUBS 0.024792f
C1639 VP.n51 VSUBS 0.029901f
C1640 VP.n52 VSUBS 0.029901f
C1641 VP.n53 VSUBS 0.029901f
C1642 VP.n54 VSUBS 0.055728f
C1643 VP.n55 VSUBS 0.029866f
C1644 VP.n56 VSUBS 1.01952f
C1645 VP.n57 VSUBS 1.85539f
C1646 VP.n58 VSUBS 1.87538f
C1647 VP.n59 VSUBS 0.039422f
C1648 VP.n60 VSUBS 0.029866f
C1649 VP.n61 VSUBS 0.055728f
C1650 VP.n62 VSUBS 0.060289f
C1651 VP.n63 VSUBS 0.029901f
C1652 VP.n64 VSUBS 0.029901f
C1653 VP.n65 VSUBS 0.029901f
C1654 VP.n66 VSUBS 0.057948f
C1655 VP.n67 VSUBS 0.055728f
C1656 VP.t1 VSUBS 2.61294f
C1657 VP.n68 VSUBS 0.924656f
C1658 VP.n69 VSUBS 0.034268f
C1659 VP.n70 VSUBS 0.029901f
C1660 VP.n71 VSUBS 0.029901f
C1661 VP.n72 VSUBS 0.029901f
C1662 VP.n73 VSUBS 0.055728f
C1663 VP.n74 VSUBS 0.037818f
C1664 VP.n75 VSUBS 0.049483f
C1665 VP.n76 VSUBS 0.029901f
C1666 VP.n77 VSUBS 0.029901f
C1667 VP.n78 VSUBS 0.029901f
C1668 VP.n79 VSUBS 0.041972f
C1669 VP.n80 VSUBS 0.924656f
C1670 VP.n81 VSUBS 0.041972f
C1671 VP.n82 VSUBS 0.055728f
C1672 VP.n83 VSUBS 0.029901f
C1673 VP.n84 VSUBS 0.029901f
C1674 VP.n85 VSUBS 0.029901f
C1675 VP.n86 VSUBS 0.037818f
C1676 VP.n87 VSUBS 0.055728f
C1677 VP.t2 VSUBS 2.61294f
C1678 VP.n88 VSUBS 0.924656f
C1679 VP.n89 VSUBS 0.049675f
C1680 VP.n90 VSUBS 0.029901f
C1681 VP.n91 VSUBS 0.029901f
C1682 VP.n92 VSUBS 0.029901f
C1683 VP.n93 VSUBS 0.055728f
C1684 VP.n94 VSUBS 0.057948f
C1685 VP.n95 VSUBS 0.024792f
C1686 VP.n96 VSUBS 0.029901f
C1687 VP.n97 VSUBS 0.029901f
C1688 VP.n98 VSUBS 0.029901f
C1689 VP.n99 VSUBS 0.055728f
C1690 VP.n100 VSUBS 0.029866f
C1691 VP.n101 VSUBS 1.01952f
C1692 VP.n102 VSUBS 0.056762f
.ends

