* NGSPICE file created from diff_pair_sample_0996.ext - technology: sky130A

.subckt diff_pair_sample_0996 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8084 pd=11.29 as=4.2744 ps=22.7 w=10.96 l=0.2
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=0 ps=0 w=10.96 l=0.2
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=0 ps=0 w=10.96 l=0.2
X3 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8084 pd=11.29 as=4.2744 ps=22.7 w=10.96 l=0.2
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=0 ps=0 w=10.96 l=0.2
X5 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=1.8084 ps=11.29 w=10.96 l=0.2
X6 VTAIL.t4 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=1.8084 ps=11.29 w=10.96 l=0.2
X7 VDD2.t1 VN.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8084 pd=11.29 as=4.2744 ps=22.7 w=10.96 l=0.2
X8 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8084 pd=11.29 as=4.2744 ps=22.7 w=10.96 l=0.2
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=0 ps=0 w=10.96 l=0.2
X10 VTAIL.t6 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=1.8084 ps=11.29 w=10.96 l=0.2
X11 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=4.2744 pd=22.7 as=1.8084 ps=11.29 w=10.96 l=0.2
R0 VN.n0 VN.t2 1518.45
R1 VN.n0 VN.t1 1518.45
R2 VN.n1 VN.t3 1518.45
R3 VN.n1 VN.t0 1518.45
R4 VN VN.n1 199.803
R5 VN VN.n0 161.351
R6 VTAIL.n5 VTAIL.t2 45.7853
R7 VTAIL.n4 VTAIL.t5 45.7853
R8 VTAIL.n3 VTAIL.t6 45.7853
R9 VTAIL.n7 VTAIL.t7 45.7852
R10 VTAIL.n0 VTAIL.t4 45.7852
R11 VTAIL.n1 VTAIL.t0 45.7852
R12 VTAIL.n2 VTAIL.t3 45.7852
R13 VTAIL.n6 VTAIL.t1 45.7852
R14 VTAIL.n7 VTAIL.n6 22.2893
R15 VTAIL.n3 VTAIL.n2 22.2893
R16 VTAIL.n5 VTAIL.n4 0.470328
R17 VTAIL.n1 VTAIL.n0 0.470328
R18 VTAIL.n4 VTAIL.n3 0.457397
R19 VTAIL.n6 VTAIL.n5 0.457397
R20 VTAIL.n2 VTAIL.n1 0.457397
R21 VTAIL VTAIL.n0 0.287138
R22 VTAIL VTAIL.n7 0.170759
R23 VDD2.n2 VDD2.n0 95.2084
R24 VDD2.n2 VDD2.n1 60.6575
R25 VDD2.n1 VDD2.t0 1.80707
R26 VDD2.n1 VDD2.t3 1.80707
R27 VDD2.n0 VDD2.t2 1.80707
R28 VDD2.n0 VDD2.t1 1.80707
R29 VDD2 VDD2.n2 0.0586897
R30 B.n50 B.t8 1557.03
R31 B.n57 B.t4 1557.03
R32 B.n238 B.t15 1557.03
R33 B.n125 B.t11 1557.03
R34 B.n375 B.n374 585
R35 B.n375 B.n28 585
R36 B.n378 B.n377 585
R37 B.n379 B.n76 585
R38 B.n381 B.n380 585
R39 B.n383 B.n75 585
R40 B.n386 B.n385 585
R41 B.n387 B.n74 585
R42 B.n389 B.n388 585
R43 B.n391 B.n73 585
R44 B.n394 B.n393 585
R45 B.n395 B.n72 585
R46 B.n397 B.n396 585
R47 B.n399 B.n71 585
R48 B.n402 B.n401 585
R49 B.n403 B.n70 585
R50 B.n405 B.n404 585
R51 B.n407 B.n69 585
R52 B.n410 B.n409 585
R53 B.n411 B.n68 585
R54 B.n413 B.n412 585
R55 B.n415 B.n67 585
R56 B.n418 B.n417 585
R57 B.n419 B.n66 585
R58 B.n421 B.n420 585
R59 B.n423 B.n65 585
R60 B.n426 B.n425 585
R61 B.n427 B.n64 585
R62 B.n429 B.n428 585
R63 B.n431 B.n63 585
R64 B.n434 B.n433 585
R65 B.n435 B.n62 585
R66 B.n437 B.n436 585
R67 B.n439 B.n61 585
R68 B.n442 B.n441 585
R69 B.n443 B.n60 585
R70 B.n445 B.n444 585
R71 B.n447 B.n59 585
R72 B.n450 B.n449 585
R73 B.n451 B.n56 585
R74 B.n454 B.n453 585
R75 B.n456 B.n55 585
R76 B.n459 B.n458 585
R77 B.n460 B.n54 585
R78 B.n462 B.n461 585
R79 B.n464 B.n53 585
R80 B.n467 B.n466 585
R81 B.n468 B.n49 585
R82 B.n470 B.n469 585
R83 B.n472 B.n48 585
R84 B.n475 B.n474 585
R85 B.n476 B.n47 585
R86 B.n478 B.n477 585
R87 B.n480 B.n46 585
R88 B.n483 B.n482 585
R89 B.n484 B.n45 585
R90 B.n486 B.n485 585
R91 B.n488 B.n44 585
R92 B.n491 B.n490 585
R93 B.n492 B.n43 585
R94 B.n494 B.n493 585
R95 B.n496 B.n42 585
R96 B.n499 B.n498 585
R97 B.n500 B.n41 585
R98 B.n502 B.n501 585
R99 B.n504 B.n40 585
R100 B.n507 B.n506 585
R101 B.n508 B.n39 585
R102 B.n510 B.n509 585
R103 B.n512 B.n38 585
R104 B.n515 B.n514 585
R105 B.n516 B.n37 585
R106 B.n518 B.n517 585
R107 B.n520 B.n36 585
R108 B.n523 B.n522 585
R109 B.n524 B.n35 585
R110 B.n526 B.n525 585
R111 B.n528 B.n34 585
R112 B.n531 B.n530 585
R113 B.n532 B.n33 585
R114 B.n534 B.n533 585
R115 B.n536 B.n32 585
R116 B.n539 B.n538 585
R117 B.n540 B.n31 585
R118 B.n542 B.n541 585
R119 B.n544 B.n30 585
R120 B.n547 B.n546 585
R121 B.n548 B.n29 585
R122 B.n373 B.n27 585
R123 B.n551 B.n27 585
R124 B.n372 B.n26 585
R125 B.n552 B.n26 585
R126 B.n371 B.n25 585
R127 B.n553 B.n25 585
R128 B.n370 B.n369 585
R129 B.n369 B.n24 585
R130 B.n368 B.n20 585
R131 B.n559 B.n20 585
R132 B.n367 B.n19 585
R133 B.n560 B.n19 585
R134 B.n366 B.n18 585
R135 B.n561 B.n18 585
R136 B.n365 B.n364 585
R137 B.n364 B.n13 585
R138 B.n363 B.n12 585
R139 B.n567 B.n12 585
R140 B.n362 B.n11 585
R141 B.n568 B.n11 585
R142 B.n361 B.n10 585
R143 B.n569 B.n10 585
R144 B.n360 B.n7 585
R145 B.n572 B.n7 585
R146 B.n359 B.n6 585
R147 B.n573 B.n6 585
R148 B.n358 B.n5 585
R149 B.n574 B.n5 585
R150 B.n357 B.n356 585
R151 B.n356 B.n4 585
R152 B.n355 B.n77 585
R153 B.n355 B.n354 585
R154 B.n345 B.n78 585
R155 B.n79 B.n78 585
R156 B.n347 B.n346 585
R157 B.n348 B.n347 585
R158 B.n344 B.n84 585
R159 B.n84 B.n83 585
R160 B.n343 B.n342 585
R161 B.n342 B.n341 585
R162 B.n86 B.n85 585
R163 B.n87 B.n86 585
R164 B.n334 B.n333 585
R165 B.n335 B.n334 585
R166 B.n332 B.n91 585
R167 B.n95 B.n91 585
R168 B.n331 B.n330 585
R169 B.n330 B.n329 585
R170 B.n93 B.n92 585
R171 B.n94 B.n93 585
R172 B.n322 B.n321 585
R173 B.n323 B.n322 585
R174 B.n98 B.n97 585
R175 B.n147 B.n146 585
R176 B.n148 B.n144 585
R177 B.n144 B.n99 585
R178 B.n150 B.n149 585
R179 B.n152 B.n143 585
R180 B.n155 B.n154 585
R181 B.n156 B.n142 585
R182 B.n158 B.n157 585
R183 B.n160 B.n141 585
R184 B.n163 B.n162 585
R185 B.n164 B.n140 585
R186 B.n166 B.n165 585
R187 B.n168 B.n139 585
R188 B.n171 B.n170 585
R189 B.n172 B.n138 585
R190 B.n174 B.n173 585
R191 B.n176 B.n137 585
R192 B.n179 B.n178 585
R193 B.n180 B.n136 585
R194 B.n182 B.n181 585
R195 B.n184 B.n135 585
R196 B.n187 B.n186 585
R197 B.n188 B.n134 585
R198 B.n190 B.n189 585
R199 B.n192 B.n133 585
R200 B.n195 B.n194 585
R201 B.n196 B.n132 585
R202 B.n198 B.n197 585
R203 B.n200 B.n131 585
R204 B.n203 B.n202 585
R205 B.n204 B.n130 585
R206 B.n206 B.n205 585
R207 B.n208 B.n129 585
R208 B.n211 B.n210 585
R209 B.n212 B.n128 585
R210 B.n214 B.n213 585
R211 B.n216 B.n127 585
R212 B.n219 B.n218 585
R213 B.n220 B.n124 585
R214 B.n223 B.n222 585
R215 B.n225 B.n123 585
R216 B.n228 B.n227 585
R217 B.n229 B.n122 585
R218 B.n231 B.n230 585
R219 B.n233 B.n121 585
R220 B.n236 B.n235 585
R221 B.n237 B.n120 585
R222 B.n242 B.n241 585
R223 B.n244 B.n119 585
R224 B.n247 B.n246 585
R225 B.n248 B.n118 585
R226 B.n250 B.n249 585
R227 B.n252 B.n117 585
R228 B.n255 B.n254 585
R229 B.n256 B.n116 585
R230 B.n258 B.n257 585
R231 B.n260 B.n115 585
R232 B.n263 B.n262 585
R233 B.n264 B.n114 585
R234 B.n266 B.n265 585
R235 B.n268 B.n113 585
R236 B.n271 B.n270 585
R237 B.n272 B.n112 585
R238 B.n274 B.n273 585
R239 B.n276 B.n111 585
R240 B.n279 B.n278 585
R241 B.n280 B.n110 585
R242 B.n282 B.n281 585
R243 B.n284 B.n109 585
R244 B.n287 B.n286 585
R245 B.n288 B.n108 585
R246 B.n290 B.n289 585
R247 B.n292 B.n107 585
R248 B.n295 B.n294 585
R249 B.n296 B.n106 585
R250 B.n298 B.n297 585
R251 B.n300 B.n105 585
R252 B.n303 B.n302 585
R253 B.n304 B.n104 585
R254 B.n306 B.n305 585
R255 B.n308 B.n103 585
R256 B.n311 B.n310 585
R257 B.n312 B.n102 585
R258 B.n314 B.n313 585
R259 B.n316 B.n101 585
R260 B.n319 B.n318 585
R261 B.n320 B.n100 585
R262 B.n325 B.n324 585
R263 B.n324 B.n323 585
R264 B.n326 B.n96 585
R265 B.n96 B.n94 585
R266 B.n328 B.n327 585
R267 B.n329 B.n328 585
R268 B.n90 B.n89 585
R269 B.n95 B.n90 585
R270 B.n337 B.n336 585
R271 B.n336 B.n335 585
R272 B.n338 B.n88 585
R273 B.n88 B.n87 585
R274 B.n340 B.n339 585
R275 B.n341 B.n340 585
R276 B.n82 B.n81 585
R277 B.n83 B.n82 585
R278 B.n350 B.n349 585
R279 B.n349 B.n348 585
R280 B.n351 B.n80 585
R281 B.n80 B.n79 585
R282 B.n353 B.n352 585
R283 B.n354 B.n353 585
R284 B.n3 B.n0 585
R285 B.n4 B.n3 585
R286 B.n571 B.n1 585
R287 B.n572 B.n571 585
R288 B.n570 B.n9 585
R289 B.n570 B.n569 585
R290 B.n15 B.n8 585
R291 B.n568 B.n8 585
R292 B.n566 B.n565 585
R293 B.n567 B.n566 585
R294 B.n564 B.n14 585
R295 B.n14 B.n13 585
R296 B.n563 B.n562 585
R297 B.n562 B.n561 585
R298 B.n17 B.n16 585
R299 B.n560 B.n17 585
R300 B.n558 B.n557 585
R301 B.n559 B.n558 585
R302 B.n556 B.n21 585
R303 B.n24 B.n21 585
R304 B.n555 B.n554 585
R305 B.n554 B.n553 585
R306 B.n23 B.n22 585
R307 B.n552 B.n23 585
R308 B.n550 B.n549 585
R309 B.n551 B.n550 585
R310 B.n575 B.n574 585
R311 B.n573 B.n2 585
R312 B.n550 B.n29 530.939
R313 B.n375 B.n27 530.939
R314 B.n322 B.n100 530.939
R315 B.n324 B.n98 530.939
R316 B.n376 B.n28 256.663
R317 B.n382 B.n28 256.663
R318 B.n384 B.n28 256.663
R319 B.n390 B.n28 256.663
R320 B.n392 B.n28 256.663
R321 B.n398 B.n28 256.663
R322 B.n400 B.n28 256.663
R323 B.n406 B.n28 256.663
R324 B.n408 B.n28 256.663
R325 B.n414 B.n28 256.663
R326 B.n416 B.n28 256.663
R327 B.n422 B.n28 256.663
R328 B.n424 B.n28 256.663
R329 B.n430 B.n28 256.663
R330 B.n432 B.n28 256.663
R331 B.n438 B.n28 256.663
R332 B.n440 B.n28 256.663
R333 B.n446 B.n28 256.663
R334 B.n448 B.n28 256.663
R335 B.n455 B.n28 256.663
R336 B.n457 B.n28 256.663
R337 B.n463 B.n28 256.663
R338 B.n465 B.n28 256.663
R339 B.n471 B.n28 256.663
R340 B.n473 B.n28 256.663
R341 B.n479 B.n28 256.663
R342 B.n481 B.n28 256.663
R343 B.n487 B.n28 256.663
R344 B.n489 B.n28 256.663
R345 B.n495 B.n28 256.663
R346 B.n497 B.n28 256.663
R347 B.n503 B.n28 256.663
R348 B.n505 B.n28 256.663
R349 B.n511 B.n28 256.663
R350 B.n513 B.n28 256.663
R351 B.n519 B.n28 256.663
R352 B.n521 B.n28 256.663
R353 B.n527 B.n28 256.663
R354 B.n529 B.n28 256.663
R355 B.n535 B.n28 256.663
R356 B.n537 B.n28 256.663
R357 B.n543 B.n28 256.663
R358 B.n545 B.n28 256.663
R359 B.n145 B.n99 256.663
R360 B.n151 B.n99 256.663
R361 B.n153 B.n99 256.663
R362 B.n159 B.n99 256.663
R363 B.n161 B.n99 256.663
R364 B.n167 B.n99 256.663
R365 B.n169 B.n99 256.663
R366 B.n175 B.n99 256.663
R367 B.n177 B.n99 256.663
R368 B.n183 B.n99 256.663
R369 B.n185 B.n99 256.663
R370 B.n191 B.n99 256.663
R371 B.n193 B.n99 256.663
R372 B.n199 B.n99 256.663
R373 B.n201 B.n99 256.663
R374 B.n207 B.n99 256.663
R375 B.n209 B.n99 256.663
R376 B.n215 B.n99 256.663
R377 B.n217 B.n99 256.663
R378 B.n224 B.n99 256.663
R379 B.n226 B.n99 256.663
R380 B.n232 B.n99 256.663
R381 B.n234 B.n99 256.663
R382 B.n243 B.n99 256.663
R383 B.n245 B.n99 256.663
R384 B.n251 B.n99 256.663
R385 B.n253 B.n99 256.663
R386 B.n259 B.n99 256.663
R387 B.n261 B.n99 256.663
R388 B.n267 B.n99 256.663
R389 B.n269 B.n99 256.663
R390 B.n275 B.n99 256.663
R391 B.n277 B.n99 256.663
R392 B.n283 B.n99 256.663
R393 B.n285 B.n99 256.663
R394 B.n291 B.n99 256.663
R395 B.n293 B.n99 256.663
R396 B.n299 B.n99 256.663
R397 B.n301 B.n99 256.663
R398 B.n307 B.n99 256.663
R399 B.n309 B.n99 256.663
R400 B.n315 B.n99 256.663
R401 B.n317 B.n99 256.663
R402 B.n577 B.n576 256.663
R403 B.n546 B.n544 163.367
R404 B.n542 B.n31 163.367
R405 B.n538 B.n536 163.367
R406 B.n534 B.n33 163.367
R407 B.n530 B.n528 163.367
R408 B.n526 B.n35 163.367
R409 B.n522 B.n520 163.367
R410 B.n518 B.n37 163.367
R411 B.n514 B.n512 163.367
R412 B.n510 B.n39 163.367
R413 B.n506 B.n504 163.367
R414 B.n502 B.n41 163.367
R415 B.n498 B.n496 163.367
R416 B.n494 B.n43 163.367
R417 B.n490 B.n488 163.367
R418 B.n486 B.n45 163.367
R419 B.n482 B.n480 163.367
R420 B.n478 B.n47 163.367
R421 B.n474 B.n472 163.367
R422 B.n470 B.n49 163.367
R423 B.n466 B.n464 163.367
R424 B.n462 B.n54 163.367
R425 B.n458 B.n456 163.367
R426 B.n454 B.n56 163.367
R427 B.n449 B.n447 163.367
R428 B.n445 B.n60 163.367
R429 B.n441 B.n439 163.367
R430 B.n437 B.n62 163.367
R431 B.n433 B.n431 163.367
R432 B.n429 B.n64 163.367
R433 B.n425 B.n423 163.367
R434 B.n421 B.n66 163.367
R435 B.n417 B.n415 163.367
R436 B.n413 B.n68 163.367
R437 B.n409 B.n407 163.367
R438 B.n405 B.n70 163.367
R439 B.n401 B.n399 163.367
R440 B.n397 B.n72 163.367
R441 B.n393 B.n391 163.367
R442 B.n389 B.n74 163.367
R443 B.n385 B.n383 163.367
R444 B.n381 B.n76 163.367
R445 B.n377 B.n375 163.367
R446 B.n322 B.n93 163.367
R447 B.n330 B.n93 163.367
R448 B.n330 B.n91 163.367
R449 B.n334 B.n91 163.367
R450 B.n334 B.n86 163.367
R451 B.n342 B.n86 163.367
R452 B.n342 B.n84 163.367
R453 B.n347 B.n84 163.367
R454 B.n347 B.n78 163.367
R455 B.n355 B.n78 163.367
R456 B.n356 B.n355 163.367
R457 B.n356 B.n5 163.367
R458 B.n6 B.n5 163.367
R459 B.n7 B.n6 163.367
R460 B.n10 B.n7 163.367
R461 B.n11 B.n10 163.367
R462 B.n12 B.n11 163.367
R463 B.n364 B.n12 163.367
R464 B.n364 B.n18 163.367
R465 B.n19 B.n18 163.367
R466 B.n20 B.n19 163.367
R467 B.n369 B.n20 163.367
R468 B.n369 B.n25 163.367
R469 B.n26 B.n25 163.367
R470 B.n27 B.n26 163.367
R471 B.n146 B.n144 163.367
R472 B.n150 B.n144 163.367
R473 B.n154 B.n152 163.367
R474 B.n158 B.n142 163.367
R475 B.n162 B.n160 163.367
R476 B.n166 B.n140 163.367
R477 B.n170 B.n168 163.367
R478 B.n174 B.n138 163.367
R479 B.n178 B.n176 163.367
R480 B.n182 B.n136 163.367
R481 B.n186 B.n184 163.367
R482 B.n190 B.n134 163.367
R483 B.n194 B.n192 163.367
R484 B.n198 B.n132 163.367
R485 B.n202 B.n200 163.367
R486 B.n206 B.n130 163.367
R487 B.n210 B.n208 163.367
R488 B.n214 B.n128 163.367
R489 B.n218 B.n216 163.367
R490 B.n223 B.n124 163.367
R491 B.n227 B.n225 163.367
R492 B.n231 B.n122 163.367
R493 B.n235 B.n233 163.367
R494 B.n242 B.n120 163.367
R495 B.n246 B.n244 163.367
R496 B.n250 B.n118 163.367
R497 B.n254 B.n252 163.367
R498 B.n258 B.n116 163.367
R499 B.n262 B.n260 163.367
R500 B.n266 B.n114 163.367
R501 B.n270 B.n268 163.367
R502 B.n274 B.n112 163.367
R503 B.n278 B.n276 163.367
R504 B.n282 B.n110 163.367
R505 B.n286 B.n284 163.367
R506 B.n290 B.n108 163.367
R507 B.n294 B.n292 163.367
R508 B.n298 B.n106 163.367
R509 B.n302 B.n300 163.367
R510 B.n306 B.n104 163.367
R511 B.n310 B.n308 163.367
R512 B.n314 B.n102 163.367
R513 B.n318 B.n316 163.367
R514 B.n324 B.n96 163.367
R515 B.n328 B.n96 163.367
R516 B.n328 B.n90 163.367
R517 B.n336 B.n90 163.367
R518 B.n336 B.n88 163.367
R519 B.n340 B.n88 163.367
R520 B.n340 B.n82 163.367
R521 B.n349 B.n82 163.367
R522 B.n349 B.n80 163.367
R523 B.n353 B.n80 163.367
R524 B.n353 B.n3 163.367
R525 B.n575 B.n3 163.367
R526 B.n571 B.n2 163.367
R527 B.n571 B.n570 163.367
R528 B.n570 B.n8 163.367
R529 B.n566 B.n8 163.367
R530 B.n566 B.n14 163.367
R531 B.n562 B.n14 163.367
R532 B.n562 B.n17 163.367
R533 B.n558 B.n17 163.367
R534 B.n558 B.n21 163.367
R535 B.n554 B.n21 163.367
R536 B.n554 B.n23 163.367
R537 B.n550 B.n23 163.367
R538 B.n323 B.n99 96.7707
R539 B.n551 B.n28 96.7707
R540 B.n57 B.t6 79.7753
R541 B.n238 B.t17 79.7753
R542 B.n50 B.t9 79.7615
R543 B.n125 B.t14 79.7615
R544 B.n545 B.n29 71.676
R545 B.n544 B.n543 71.676
R546 B.n537 B.n31 71.676
R547 B.n536 B.n535 71.676
R548 B.n529 B.n33 71.676
R549 B.n528 B.n527 71.676
R550 B.n521 B.n35 71.676
R551 B.n520 B.n519 71.676
R552 B.n513 B.n37 71.676
R553 B.n512 B.n511 71.676
R554 B.n505 B.n39 71.676
R555 B.n504 B.n503 71.676
R556 B.n497 B.n41 71.676
R557 B.n496 B.n495 71.676
R558 B.n489 B.n43 71.676
R559 B.n488 B.n487 71.676
R560 B.n481 B.n45 71.676
R561 B.n480 B.n479 71.676
R562 B.n473 B.n47 71.676
R563 B.n472 B.n471 71.676
R564 B.n465 B.n49 71.676
R565 B.n464 B.n463 71.676
R566 B.n457 B.n54 71.676
R567 B.n456 B.n455 71.676
R568 B.n448 B.n56 71.676
R569 B.n447 B.n446 71.676
R570 B.n440 B.n60 71.676
R571 B.n439 B.n438 71.676
R572 B.n432 B.n62 71.676
R573 B.n431 B.n430 71.676
R574 B.n424 B.n64 71.676
R575 B.n423 B.n422 71.676
R576 B.n416 B.n66 71.676
R577 B.n415 B.n414 71.676
R578 B.n408 B.n68 71.676
R579 B.n407 B.n406 71.676
R580 B.n400 B.n70 71.676
R581 B.n399 B.n398 71.676
R582 B.n392 B.n72 71.676
R583 B.n391 B.n390 71.676
R584 B.n384 B.n74 71.676
R585 B.n383 B.n382 71.676
R586 B.n376 B.n76 71.676
R587 B.n377 B.n376 71.676
R588 B.n382 B.n381 71.676
R589 B.n385 B.n384 71.676
R590 B.n390 B.n389 71.676
R591 B.n393 B.n392 71.676
R592 B.n398 B.n397 71.676
R593 B.n401 B.n400 71.676
R594 B.n406 B.n405 71.676
R595 B.n409 B.n408 71.676
R596 B.n414 B.n413 71.676
R597 B.n417 B.n416 71.676
R598 B.n422 B.n421 71.676
R599 B.n425 B.n424 71.676
R600 B.n430 B.n429 71.676
R601 B.n433 B.n432 71.676
R602 B.n438 B.n437 71.676
R603 B.n441 B.n440 71.676
R604 B.n446 B.n445 71.676
R605 B.n449 B.n448 71.676
R606 B.n455 B.n454 71.676
R607 B.n458 B.n457 71.676
R608 B.n463 B.n462 71.676
R609 B.n466 B.n465 71.676
R610 B.n471 B.n470 71.676
R611 B.n474 B.n473 71.676
R612 B.n479 B.n478 71.676
R613 B.n482 B.n481 71.676
R614 B.n487 B.n486 71.676
R615 B.n490 B.n489 71.676
R616 B.n495 B.n494 71.676
R617 B.n498 B.n497 71.676
R618 B.n503 B.n502 71.676
R619 B.n506 B.n505 71.676
R620 B.n511 B.n510 71.676
R621 B.n514 B.n513 71.676
R622 B.n519 B.n518 71.676
R623 B.n522 B.n521 71.676
R624 B.n527 B.n526 71.676
R625 B.n530 B.n529 71.676
R626 B.n535 B.n534 71.676
R627 B.n538 B.n537 71.676
R628 B.n543 B.n542 71.676
R629 B.n546 B.n545 71.676
R630 B.n145 B.n98 71.676
R631 B.n151 B.n150 71.676
R632 B.n154 B.n153 71.676
R633 B.n159 B.n158 71.676
R634 B.n162 B.n161 71.676
R635 B.n167 B.n166 71.676
R636 B.n170 B.n169 71.676
R637 B.n175 B.n174 71.676
R638 B.n178 B.n177 71.676
R639 B.n183 B.n182 71.676
R640 B.n186 B.n185 71.676
R641 B.n191 B.n190 71.676
R642 B.n194 B.n193 71.676
R643 B.n199 B.n198 71.676
R644 B.n202 B.n201 71.676
R645 B.n207 B.n206 71.676
R646 B.n210 B.n209 71.676
R647 B.n215 B.n214 71.676
R648 B.n218 B.n217 71.676
R649 B.n224 B.n223 71.676
R650 B.n227 B.n226 71.676
R651 B.n232 B.n231 71.676
R652 B.n235 B.n234 71.676
R653 B.n243 B.n242 71.676
R654 B.n246 B.n245 71.676
R655 B.n251 B.n250 71.676
R656 B.n254 B.n253 71.676
R657 B.n259 B.n258 71.676
R658 B.n262 B.n261 71.676
R659 B.n267 B.n266 71.676
R660 B.n270 B.n269 71.676
R661 B.n275 B.n274 71.676
R662 B.n278 B.n277 71.676
R663 B.n283 B.n282 71.676
R664 B.n286 B.n285 71.676
R665 B.n291 B.n290 71.676
R666 B.n294 B.n293 71.676
R667 B.n299 B.n298 71.676
R668 B.n302 B.n301 71.676
R669 B.n307 B.n306 71.676
R670 B.n310 B.n309 71.676
R671 B.n315 B.n314 71.676
R672 B.n318 B.n317 71.676
R673 B.n146 B.n145 71.676
R674 B.n152 B.n151 71.676
R675 B.n153 B.n142 71.676
R676 B.n160 B.n159 71.676
R677 B.n161 B.n140 71.676
R678 B.n168 B.n167 71.676
R679 B.n169 B.n138 71.676
R680 B.n176 B.n175 71.676
R681 B.n177 B.n136 71.676
R682 B.n184 B.n183 71.676
R683 B.n185 B.n134 71.676
R684 B.n192 B.n191 71.676
R685 B.n193 B.n132 71.676
R686 B.n200 B.n199 71.676
R687 B.n201 B.n130 71.676
R688 B.n208 B.n207 71.676
R689 B.n209 B.n128 71.676
R690 B.n216 B.n215 71.676
R691 B.n217 B.n124 71.676
R692 B.n225 B.n224 71.676
R693 B.n226 B.n122 71.676
R694 B.n233 B.n232 71.676
R695 B.n234 B.n120 71.676
R696 B.n244 B.n243 71.676
R697 B.n245 B.n118 71.676
R698 B.n252 B.n251 71.676
R699 B.n253 B.n116 71.676
R700 B.n260 B.n259 71.676
R701 B.n261 B.n114 71.676
R702 B.n268 B.n267 71.676
R703 B.n269 B.n112 71.676
R704 B.n276 B.n275 71.676
R705 B.n277 B.n110 71.676
R706 B.n284 B.n283 71.676
R707 B.n285 B.n108 71.676
R708 B.n292 B.n291 71.676
R709 B.n293 B.n106 71.676
R710 B.n300 B.n299 71.676
R711 B.n301 B.n104 71.676
R712 B.n308 B.n307 71.676
R713 B.n309 B.n102 71.676
R714 B.n316 B.n315 71.676
R715 B.n317 B.n100 71.676
R716 B.n576 B.n575 71.676
R717 B.n576 B.n2 71.676
R718 B.n58 B.t7 69.4965
R719 B.n239 B.t16 69.4965
R720 B.n51 B.t10 69.4827
R721 B.n126 B.t13 69.4827
R722 B.n52 B.n51 59.5399
R723 B.n452 B.n58 59.5399
R724 B.n240 B.n239 59.5399
R725 B.n221 B.n126 59.5399
R726 B.n323 B.n94 46.0171
R727 B.n329 B.n94 46.0171
R728 B.n329 B.n95 46.0171
R729 B.n335 B.n87 46.0171
R730 B.n341 B.n87 46.0171
R731 B.n341 B.n83 46.0171
R732 B.n348 B.n83 46.0171
R733 B.n354 B.n79 46.0171
R734 B.n574 B.n4 46.0171
R735 B.n574 B.n573 46.0171
R736 B.n573 B.n572 46.0171
R737 B.n569 B.n568 46.0171
R738 B.n567 B.n13 46.0171
R739 B.n561 B.n13 46.0171
R740 B.n561 B.n560 46.0171
R741 B.n560 B.n559 46.0171
R742 B.n553 B.n24 46.0171
R743 B.n553 B.n552 46.0171
R744 B.n552 B.n551 46.0171
R745 B.t0 B.n4 40.6034
R746 B.n572 B.t2 40.6034
R747 B.n95 B.t12 36.5431
R748 B.n24 B.t5 36.5431
R749 B.n325 B.n97 34.4981
R750 B.n321 B.n320 34.4981
R751 B.n374 B.n373 34.4981
R752 B.n549 B.n548 34.4981
R753 B.n348 B.t3 25.7157
R754 B.t1 B.n567 25.7157
R755 B.t3 B.n79 20.3019
R756 B.n568 B.t1 20.3019
R757 B B.n577 18.0485
R758 B.n326 B.n325 10.6151
R759 B.n327 B.n326 10.6151
R760 B.n327 B.n89 10.6151
R761 B.n337 B.n89 10.6151
R762 B.n338 B.n337 10.6151
R763 B.n339 B.n338 10.6151
R764 B.n339 B.n81 10.6151
R765 B.n350 B.n81 10.6151
R766 B.n351 B.n350 10.6151
R767 B.n352 B.n351 10.6151
R768 B.n352 B.n0 10.6151
R769 B.n147 B.n97 10.6151
R770 B.n148 B.n147 10.6151
R771 B.n149 B.n148 10.6151
R772 B.n149 B.n143 10.6151
R773 B.n155 B.n143 10.6151
R774 B.n156 B.n155 10.6151
R775 B.n157 B.n156 10.6151
R776 B.n157 B.n141 10.6151
R777 B.n163 B.n141 10.6151
R778 B.n164 B.n163 10.6151
R779 B.n165 B.n164 10.6151
R780 B.n165 B.n139 10.6151
R781 B.n171 B.n139 10.6151
R782 B.n172 B.n171 10.6151
R783 B.n173 B.n172 10.6151
R784 B.n173 B.n137 10.6151
R785 B.n179 B.n137 10.6151
R786 B.n180 B.n179 10.6151
R787 B.n181 B.n180 10.6151
R788 B.n181 B.n135 10.6151
R789 B.n187 B.n135 10.6151
R790 B.n188 B.n187 10.6151
R791 B.n189 B.n188 10.6151
R792 B.n189 B.n133 10.6151
R793 B.n195 B.n133 10.6151
R794 B.n196 B.n195 10.6151
R795 B.n197 B.n196 10.6151
R796 B.n197 B.n131 10.6151
R797 B.n203 B.n131 10.6151
R798 B.n204 B.n203 10.6151
R799 B.n205 B.n204 10.6151
R800 B.n205 B.n129 10.6151
R801 B.n211 B.n129 10.6151
R802 B.n212 B.n211 10.6151
R803 B.n213 B.n212 10.6151
R804 B.n213 B.n127 10.6151
R805 B.n219 B.n127 10.6151
R806 B.n220 B.n219 10.6151
R807 B.n222 B.n123 10.6151
R808 B.n228 B.n123 10.6151
R809 B.n229 B.n228 10.6151
R810 B.n230 B.n229 10.6151
R811 B.n230 B.n121 10.6151
R812 B.n236 B.n121 10.6151
R813 B.n237 B.n236 10.6151
R814 B.n241 B.n237 10.6151
R815 B.n247 B.n119 10.6151
R816 B.n248 B.n247 10.6151
R817 B.n249 B.n248 10.6151
R818 B.n249 B.n117 10.6151
R819 B.n255 B.n117 10.6151
R820 B.n256 B.n255 10.6151
R821 B.n257 B.n256 10.6151
R822 B.n257 B.n115 10.6151
R823 B.n263 B.n115 10.6151
R824 B.n264 B.n263 10.6151
R825 B.n265 B.n264 10.6151
R826 B.n265 B.n113 10.6151
R827 B.n271 B.n113 10.6151
R828 B.n272 B.n271 10.6151
R829 B.n273 B.n272 10.6151
R830 B.n273 B.n111 10.6151
R831 B.n279 B.n111 10.6151
R832 B.n280 B.n279 10.6151
R833 B.n281 B.n280 10.6151
R834 B.n281 B.n109 10.6151
R835 B.n287 B.n109 10.6151
R836 B.n288 B.n287 10.6151
R837 B.n289 B.n288 10.6151
R838 B.n289 B.n107 10.6151
R839 B.n295 B.n107 10.6151
R840 B.n296 B.n295 10.6151
R841 B.n297 B.n296 10.6151
R842 B.n297 B.n105 10.6151
R843 B.n303 B.n105 10.6151
R844 B.n304 B.n303 10.6151
R845 B.n305 B.n304 10.6151
R846 B.n305 B.n103 10.6151
R847 B.n311 B.n103 10.6151
R848 B.n312 B.n311 10.6151
R849 B.n313 B.n312 10.6151
R850 B.n313 B.n101 10.6151
R851 B.n319 B.n101 10.6151
R852 B.n320 B.n319 10.6151
R853 B.n321 B.n92 10.6151
R854 B.n331 B.n92 10.6151
R855 B.n332 B.n331 10.6151
R856 B.n333 B.n332 10.6151
R857 B.n333 B.n85 10.6151
R858 B.n343 B.n85 10.6151
R859 B.n344 B.n343 10.6151
R860 B.n346 B.n344 10.6151
R861 B.n346 B.n345 10.6151
R862 B.n345 B.n77 10.6151
R863 B.n357 B.n77 10.6151
R864 B.n358 B.n357 10.6151
R865 B.n359 B.n358 10.6151
R866 B.n360 B.n359 10.6151
R867 B.n361 B.n360 10.6151
R868 B.n362 B.n361 10.6151
R869 B.n363 B.n362 10.6151
R870 B.n365 B.n363 10.6151
R871 B.n366 B.n365 10.6151
R872 B.n367 B.n366 10.6151
R873 B.n368 B.n367 10.6151
R874 B.n370 B.n368 10.6151
R875 B.n371 B.n370 10.6151
R876 B.n372 B.n371 10.6151
R877 B.n373 B.n372 10.6151
R878 B.n9 B.n1 10.6151
R879 B.n15 B.n9 10.6151
R880 B.n565 B.n15 10.6151
R881 B.n565 B.n564 10.6151
R882 B.n564 B.n563 10.6151
R883 B.n563 B.n16 10.6151
R884 B.n557 B.n16 10.6151
R885 B.n557 B.n556 10.6151
R886 B.n556 B.n555 10.6151
R887 B.n555 B.n22 10.6151
R888 B.n549 B.n22 10.6151
R889 B.n548 B.n547 10.6151
R890 B.n547 B.n30 10.6151
R891 B.n541 B.n30 10.6151
R892 B.n541 B.n540 10.6151
R893 B.n540 B.n539 10.6151
R894 B.n539 B.n32 10.6151
R895 B.n533 B.n32 10.6151
R896 B.n533 B.n532 10.6151
R897 B.n532 B.n531 10.6151
R898 B.n531 B.n34 10.6151
R899 B.n525 B.n34 10.6151
R900 B.n525 B.n524 10.6151
R901 B.n524 B.n523 10.6151
R902 B.n523 B.n36 10.6151
R903 B.n517 B.n36 10.6151
R904 B.n517 B.n516 10.6151
R905 B.n516 B.n515 10.6151
R906 B.n515 B.n38 10.6151
R907 B.n509 B.n38 10.6151
R908 B.n509 B.n508 10.6151
R909 B.n508 B.n507 10.6151
R910 B.n507 B.n40 10.6151
R911 B.n501 B.n40 10.6151
R912 B.n501 B.n500 10.6151
R913 B.n500 B.n499 10.6151
R914 B.n499 B.n42 10.6151
R915 B.n493 B.n42 10.6151
R916 B.n493 B.n492 10.6151
R917 B.n492 B.n491 10.6151
R918 B.n491 B.n44 10.6151
R919 B.n485 B.n44 10.6151
R920 B.n485 B.n484 10.6151
R921 B.n484 B.n483 10.6151
R922 B.n483 B.n46 10.6151
R923 B.n477 B.n46 10.6151
R924 B.n477 B.n476 10.6151
R925 B.n476 B.n475 10.6151
R926 B.n475 B.n48 10.6151
R927 B.n469 B.n468 10.6151
R928 B.n468 B.n467 10.6151
R929 B.n467 B.n53 10.6151
R930 B.n461 B.n53 10.6151
R931 B.n461 B.n460 10.6151
R932 B.n460 B.n459 10.6151
R933 B.n459 B.n55 10.6151
R934 B.n453 B.n55 10.6151
R935 B.n451 B.n450 10.6151
R936 B.n450 B.n59 10.6151
R937 B.n444 B.n59 10.6151
R938 B.n444 B.n443 10.6151
R939 B.n443 B.n442 10.6151
R940 B.n442 B.n61 10.6151
R941 B.n436 B.n61 10.6151
R942 B.n436 B.n435 10.6151
R943 B.n435 B.n434 10.6151
R944 B.n434 B.n63 10.6151
R945 B.n428 B.n63 10.6151
R946 B.n428 B.n427 10.6151
R947 B.n427 B.n426 10.6151
R948 B.n426 B.n65 10.6151
R949 B.n420 B.n65 10.6151
R950 B.n420 B.n419 10.6151
R951 B.n419 B.n418 10.6151
R952 B.n418 B.n67 10.6151
R953 B.n412 B.n67 10.6151
R954 B.n412 B.n411 10.6151
R955 B.n411 B.n410 10.6151
R956 B.n410 B.n69 10.6151
R957 B.n404 B.n69 10.6151
R958 B.n404 B.n403 10.6151
R959 B.n403 B.n402 10.6151
R960 B.n402 B.n71 10.6151
R961 B.n396 B.n71 10.6151
R962 B.n396 B.n395 10.6151
R963 B.n395 B.n394 10.6151
R964 B.n394 B.n73 10.6151
R965 B.n388 B.n73 10.6151
R966 B.n388 B.n387 10.6151
R967 B.n387 B.n386 10.6151
R968 B.n386 B.n75 10.6151
R969 B.n380 B.n75 10.6151
R970 B.n380 B.n379 10.6151
R971 B.n379 B.n378 10.6151
R972 B.n378 B.n374 10.6151
R973 B.n51 B.n50 10.2793
R974 B.n58 B.n57 10.2793
R975 B.n239 B.n238 10.2793
R976 B.n126 B.n125 10.2793
R977 B.n335 B.t12 9.47451
R978 B.n559 B.t5 9.47451
R979 B.n577 B.n0 8.11757
R980 B.n577 B.n1 8.11757
R981 B.n222 B.n221 7.18099
R982 B.n241 B.n240 7.18099
R983 B.n469 B.n52 7.18099
R984 B.n453 B.n452 7.18099
R985 B.n354 B.t0 5.41422
R986 B.n569 B.t2 5.41422
R987 B.n221 B.n220 3.43465
R988 B.n240 B.n119 3.43465
R989 B.n52 B.n48 3.43465
R990 B.n452 B.n451 3.43465
R991 VP.n1 VP.t0 1518.45
R992 VP.n1 VP.t1 1518.45
R993 VP.n0 VP.t3 1518.45
R994 VP.n0 VP.t2 1518.45
R995 VP.n2 VP.n0 199.422
R996 VP.n2 VP.n1 161.3
R997 VP VP.n2 0.0516364
R998 VDD1 VDD1.n1 95.7332
R999 VDD1 VDD1.n0 60.7156
R1000 VDD1.n0 VDD1.t0 1.80707
R1001 VDD1.n0 VDD1.t1 1.80707
R1002 VDD1.n1 VDD1.t2 1.80707
R1003 VDD1.n1 VDD1.t3 1.80707
C0 VDD1 VP 1.67779f
C1 VDD1 VN 0.147636f
C2 VDD2 VDD1 0.458222f
C3 VN VP 4.26893f
C4 VDD2 VP 0.242395f
C5 VDD2 VN 1.58317f
C6 VDD1 VTAIL 10.1305f
C7 VTAIL VP 1.07617f
C8 VN VTAIL 1.06206f
C9 VDD2 VTAIL 10.1687f
C10 VDD2 B 2.33246f
C11 VDD1 B 6.05143f
C12 VTAIL B 7.415233f
C13 VN B 6.44759f
C14 VP B 3.764326f
C15 VDD1.t0 B 0.268112f
C16 VDD1.t1 B 0.268112f
C17 VDD1.n0 B 2.37366f
C18 VDD1.t2 B 0.268112f
C19 VDD1.t3 B 0.268112f
C20 VDD1.n1 B 3.01017f
C21 VP.t3 B 0.252142f
C22 VP.t2 B 0.252142f
C23 VP.n0 B 0.485991f
C24 VP.t1 B 0.252142f
C25 VP.t0 B 0.252142f
C26 VP.n1 B 0.216425f
C27 VP.n2 B 2.57426f
C28 VDD2.t2 B 0.273867f
C29 VDD2.t1 B 0.273867f
C30 VDD2.n0 B 3.04512f
C31 VDD2.t0 B 0.273867f
C32 VDD2.t3 B 0.273867f
C33 VDD2.n1 B 2.4243f
C34 VDD2.n2 B 3.58176f
C35 VTAIL.t4 B 1.79865f
C36 VTAIL.n0 B 0.305719f
C37 VTAIL.t0 B 1.79865f
C38 VTAIL.n1 B 0.316248f
C39 VTAIL.t3 B 1.79865f
C40 VTAIL.n2 B 1.16146f
C41 VTAIL.t6 B 1.79866f
C42 VTAIL.n3 B 1.16145f
C43 VTAIL.t5 B 1.79866f
C44 VTAIL.n4 B 0.316235f
C45 VTAIL.t2 B 1.79866f
C46 VTAIL.n5 B 0.316235f
C47 VTAIL.t1 B 1.79865f
C48 VTAIL.n6 B 1.16146f
C49 VTAIL.t7 B 1.79865f
C50 VTAIL.n7 B 1.14374f
C51 VN.t1 B 0.24887f
C52 VN.t2 B 0.24887f
C53 VN.n0 B 0.213627f
C54 VN.t3 B 0.24887f
C55 VN.t0 B 0.24887f
C56 VN.n1 B 0.486882f
.ends

