* NGSPICE file created from diff_pair_sample_1598.ext - technology: sky130A

.subckt diff_pair_sample_1598 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=1.28
X1 VDD1.t9 VP.t0 VTAIL.t14 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=1.28
X2 B.t8 B.t6 B.t7 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=1.28
X3 VTAIL.t11 VP.t1 VDD1.t8 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X4 VDD2.t9 VN.t0 VTAIL.t6 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=1.28
X5 VDD2.t8 VN.t1 VTAIL.t0 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X6 VTAIL.t4 VN.t2 VDD2.t7 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X7 VDD2.t6 VN.t3 VTAIL.t1 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=1.28
X8 VDD1.t7 VP.t2 VTAIL.t15 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=1.28
X9 VTAIL.t19 VP.t3 VDD1.t6 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X10 VDD1.t5 VP.t4 VTAIL.t18 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=1.28
X11 VDD2.t5 VN.t4 VTAIL.t5 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=1.28
X12 VDD1.t4 VP.t5 VTAIL.t17 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X13 VDD1.t3 VP.t6 VTAIL.t12 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=5.8539 ps=30.8 w=15.01 l=1.28
X14 B.t5 B.t3 B.t4 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=1.28
X15 VTAIL.t8 VN.t5 VDD2.t4 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X16 VTAIL.t3 VN.t6 VDD2.t3 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X17 VTAIL.t7 VN.t7 VDD2.t2 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X18 VDD2.t1 VN.t8 VTAIL.t2 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=2.47665 ps=15.34 w=15.01 l=1.28
X19 VTAIL.t16 VP.t7 VDD1.t2 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X20 VTAIL.t13 VP.t8 VDD1.t1 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X21 VDD1.t0 VP.t9 VTAIL.t10 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
X22 B.t2 B.t0 B.t1 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=5.8539 pd=30.8 as=0 ps=0 w=15.01 l=1.28
X23 VDD2.t0 VN.t9 VTAIL.t9 w_n2902_n3970# sky130_fd_pr__pfet_01v8 ad=2.47665 pd=15.34 as=2.47665 ps=15.34 w=15.01 l=1.28
R0 B.n412 B.n411 585
R1 B.n410 B.n117 585
R2 B.n409 B.n408 585
R3 B.n407 B.n118 585
R4 B.n406 B.n405 585
R5 B.n404 B.n119 585
R6 B.n403 B.n402 585
R7 B.n401 B.n120 585
R8 B.n400 B.n399 585
R9 B.n398 B.n121 585
R10 B.n397 B.n396 585
R11 B.n395 B.n122 585
R12 B.n394 B.n393 585
R13 B.n392 B.n123 585
R14 B.n391 B.n390 585
R15 B.n389 B.n124 585
R16 B.n388 B.n387 585
R17 B.n386 B.n125 585
R18 B.n385 B.n384 585
R19 B.n383 B.n126 585
R20 B.n382 B.n381 585
R21 B.n380 B.n127 585
R22 B.n379 B.n378 585
R23 B.n377 B.n128 585
R24 B.n376 B.n375 585
R25 B.n374 B.n129 585
R26 B.n373 B.n372 585
R27 B.n371 B.n130 585
R28 B.n370 B.n369 585
R29 B.n368 B.n131 585
R30 B.n367 B.n366 585
R31 B.n365 B.n132 585
R32 B.n364 B.n363 585
R33 B.n362 B.n133 585
R34 B.n361 B.n360 585
R35 B.n359 B.n134 585
R36 B.n358 B.n357 585
R37 B.n356 B.n135 585
R38 B.n355 B.n354 585
R39 B.n353 B.n136 585
R40 B.n352 B.n351 585
R41 B.n350 B.n137 585
R42 B.n349 B.n348 585
R43 B.n347 B.n138 585
R44 B.n346 B.n345 585
R45 B.n344 B.n139 585
R46 B.n343 B.n342 585
R47 B.n341 B.n140 585
R48 B.n340 B.n339 585
R49 B.n338 B.n141 585
R50 B.n336 B.n335 585
R51 B.n334 B.n144 585
R52 B.n333 B.n332 585
R53 B.n331 B.n145 585
R54 B.n330 B.n329 585
R55 B.n328 B.n146 585
R56 B.n327 B.n326 585
R57 B.n325 B.n147 585
R58 B.n324 B.n323 585
R59 B.n322 B.n148 585
R60 B.n321 B.n320 585
R61 B.n316 B.n149 585
R62 B.n315 B.n314 585
R63 B.n313 B.n150 585
R64 B.n312 B.n311 585
R65 B.n310 B.n151 585
R66 B.n309 B.n308 585
R67 B.n307 B.n152 585
R68 B.n306 B.n305 585
R69 B.n304 B.n153 585
R70 B.n303 B.n302 585
R71 B.n301 B.n154 585
R72 B.n300 B.n299 585
R73 B.n298 B.n155 585
R74 B.n297 B.n296 585
R75 B.n295 B.n156 585
R76 B.n294 B.n293 585
R77 B.n292 B.n157 585
R78 B.n291 B.n290 585
R79 B.n289 B.n158 585
R80 B.n288 B.n287 585
R81 B.n286 B.n159 585
R82 B.n285 B.n284 585
R83 B.n283 B.n160 585
R84 B.n282 B.n281 585
R85 B.n280 B.n161 585
R86 B.n279 B.n278 585
R87 B.n277 B.n162 585
R88 B.n276 B.n275 585
R89 B.n274 B.n163 585
R90 B.n273 B.n272 585
R91 B.n271 B.n164 585
R92 B.n270 B.n269 585
R93 B.n268 B.n165 585
R94 B.n267 B.n266 585
R95 B.n265 B.n166 585
R96 B.n264 B.n263 585
R97 B.n262 B.n167 585
R98 B.n261 B.n260 585
R99 B.n259 B.n168 585
R100 B.n258 B.n257 585
R101 B.n256 B.n169 585
R102 B.n255 B.n254 585
R103 B.n253 B.n170 585
R104 B.n252 B.n251 585
R105 B.n250 B.n171 585
R106 B.n249 B.n248 585
R107 B.n247 B.n172 585
R108 B.n246 B.n245 585
R109 B.n244 B.n173 585
R110 B.n413 B.n116 585
R111 B.n415 B.n414 585
R112 B.n416 B.n115 585
R113 B.n418 B.n417 585
R114 B.n419 B.n114 585
R115 B.n421 B.n420 585
R116 B.n422 B.n113 585
R117 B.n424 B.n423 585
R118 B.n425 B.n112 585
R119 B.n427 B.n426 585
R120 B.n428 B.n111 585
R121 B.n430 B.n429 585
R122 B.n431 B.n110 585
R123 B.n433 B.n432 585
R124 B.n434 B.n109 585
R125 B.n436 B.n435 585
R126 B.n437 B.n108 585
R127 B.n439 B.n438 585
R128 B.n440 B.n107 585
R129 B.n442 B.n441 585
R130 B.n443 B.n106 585
R131 B.n445 B.n444 585
R132 B.n446 B.n105 585
R133 B.n448 B.n447 585
R134 B.n449 B.n104 585
R135 B.n451 B.n450 585
R136 B.n452 B.n103 585
R137 B.n454 B.n453 585
R138 B.n455 B.n102 585
R139 B.n457 B.n456 585
R140 B.n458 B.n101 585
R141 B.n460 B.n459 585
R142 B.n461 B.n100 585
R143 B.n463 B.n462 585
R144 B.n464 B.n99 585
R145 B.n466 B.n465 585
R146 B.n467 B.n98 585
R147 B.n469 B.n468 585
R148 B.n470 B.n97 585
R149 B.n472 B.n471 585
R150 B.n473 B.n96 585
R151 B.n475 B.n474 585
R152 B.n476 B.n95 585
R153 B.n478 B.n477 585
R154 B.n479 B.n94 585
R155 B.n481 B.n480 585
R156 B.n482 B.n93 585
R157 B.n484 B.n483 585
R158 B.n485 B.n92 585
R159 B.n487 B.n486 585
R160 B.n488 B.n91 585
R161 B.n490 B.n489 585
R162 B.n491 B.n90 585
R163 B.n493 B.n492 585
R164 B.n494 B.n89 585
R165 B.n496 B.n495 585
R166 B.n497 B.n88 585
R167 B.n499 B.n498 585
R168 B.n500 B.n87 585
R169 B.n502 B.n501 585
R170 B.n503 B.n86 585
R171 B.n505 B.n504 585
R172 B.n506 B.n85 585
R173 B.n508 B.n507 585
R174 B.n509 B.n84 585
R175 B.n511 B.n510 585
R176 B.n512 B.n83 585
R177 B.n514 B.n513 585
R178 B.n515 B.n82 585
R179 B.n517 B.n516 585
R180 B.n518 B.n81 585
R181 B.n520 B.n519 585
R182 B.n521 B.n80 585
R183 B.n523 B.n522 585
R184 B.n689 B.n20 585
R185 B.n688 B.n687 585
R186 B.n686 B.n21 585
R187 B.n685 B.n684 585
R188 B.n683 B.n22 585
R189 B.n682 B.n681 585
R190 B.n680 B.n23 585
R191 B.n679 B.n678 585
R192 B.n677 B.n24 585
R193 B.n676 B.n675 585
R194 B.n674 B.n25 585
R195 B.n673 B.n672 585
R196 B.n671 B.n26 585
R197 B.n670 B.n669 585
R198 B.n668 B.n27 585
R199 B.n667 B.n666 585
R200 B.n665 B.n28 585
R201 B.n664 B.n663 585
R202 B.n662 B.n29 585
R203 B.n661 B.n660 585
R204 B.n659 B.n30 585
R205 B.n658 B.n657 585
R206 B.n656 B.n31 585
R207 B.n655 B.n654 585
R208 B.n653 B.n32 585
R209 B.n652 B.n651 585
R210 B.n650 B.n33 585
R211 B.n649 B.n648 585
R212 B.n647 B.n34 585
R213 B.n646 B.n645 585
R214 B.n644 B.n35 585
R215 B.n643 B.n642 585
R216 B.n641 B.n36 585
R217 B.n640 B.n639 585
R218 B.n638 B.n37 585
R219 B.n637 B.n636 585
R220 B.n635 B.n38 585
R221 B.n634 B.n633 585
R222 B.n632 B.n39 585
R223 B.n631 B.n630 585
R224 B.n629 B.n40 585
R225 B.n628 B.n627 585
R226 B.n626 B.n41 585
R227 B.n625 B.n624 585
R228 B.n623 B.n42 585
R229 B.n622 B.n621 585
R230 B.n620 B.n43 585
R231 B.n619 B.n618 585
R232 B.n617 B.n44 585
R233 B.n616 B.n615 585
R234 B.n613 B.n45 585
R235 B.n612 B.n611 585
R236 B.n610 B.n48 585
R237 B.n609 B.n608 585
R238 B.n607 B.n49 585
R239 B.n606 B.n605 585
R240 B.n604 B.n50 585
R241 B.n603 B.n602 585
R242 B.n601 B.n51 585
R243 B.n600 B.n599 585
R244 B.n598 B.n597 585
R245 B.n596 B.n55 585
R246 B.n595 B.n594 585
R247 B.n593 B.n56 585
R248 B.n592 B.n591 585
R249 B.n590 B.n57 585
R250 B.n589 B.n588 585
R251 B.n587 B.n58 585
R252 B.n586 B.n585 585
R253 B.n584 B.n59 585
R254 B.n583 B.n582 585
R255 B.n581 B.n60 585
R256 B.n580 B.n579 585
R257 B.n578 B.n61 585
R258 B.n577 B.n576 585
R259 B.n575 B.n62 585
R260 B.n574 B.n573 585
R261 B.n572 B.n63 585
R262 B.n571 B.n570 585
R263 B.n569 B.n64 585
R264 B.n568 B.n567 585
R265 B.n566 B.n65 585
R266 B.n565 B.n564 585
R267 B.n563 B.n66 585
R268 B.n562 B.n561 585
R269 B.n560 B.n67 585
R270 B.n559 B.n558 585
R271 B.n557 B.n68 585
R272 B.n556 B.n555 585
R273 B.n554 B.n69 585
R274 B.n553 B.n552 585
R275 B.n551 B.n70 585
R276 B.n550 B.n549 585
R277 B.n548 B.n71 585
R278 B.n547 B.n546 585
R279 B.n545 B.n72 585
R280 B.n544 B.n543 585
R281 B.n542 B.n73 585
R282 B.n541 B.n540 585
R283 B.n539 B.n74 585
R284 B.n538 B.n537 585
R285 B.n536 B.n75 585
R286 B.n535 B.n534 585
R287 B.n533 B.n76 585
R288 B.n532 B.n531 585
R289 B.n530 B.n77 585
R290 B.n529 B.n528 585
R291 B.n527 B.n78 585
R292 B.n526 B.n525 585
R293 B.n524 B.n79 585
R294 B.n691 B.n690 585
R295 B.n692 B.n19 585
R296 B.n694 B.n693 585
R297 B.n695 B.n18 585
R298 B.n697 B.n696 585
R299 B.n698 B.n17 585
R300 B.n700 B.n699 585
R301 B.n701 B.n16 585
R302 B.n703 B.n702 585
R303 B.n704 B.n15 585
R304 B.n706 B.n705 585
R305 B.n707 B.n14 585
R306 B.n709 B.n708 585
R307 B.n710 B.n13 585
R308 B.n712 B.n711 585
R309 B.n713 B.n12 585
R310 B.n715 B.n714 585
R311 B.n716 B.n11 585
R312 B.n718 B.n717 585
R313 B.n719 B.n10 585
R314 B.n721 B.n720 585
R315 B.n722 B.n9 585
R316 B.n724 B.n723 585
R317 B.n725 B.n8 585
R318 B.n727 B.n726 585
R319 B.n728 B.n7 585
R320 B.n730 B.n729 585
R321 B.n731 B.n6 585
R322 B.n733 B.n732 585
R323 B.n734 B.n5 585
R324 B.n736 B.n735 585
R325 B.n737 B.n4 585
R326 B.n739 B.n738 585
R327 B.n740 B.n3 585
R328 B.n742 B.n741 585
R329 B.n743 B.n0 585
R330 B.n2 B.n1 585
R331 B.n192 B.n191 585
R332 B.n193 B.n190 585
R333 B.n195 B.n194 585
R334 B.n196 B.n189 585
R335 B.n198 B.n197 585
R336 B.n199 B.n188 585
R337 B.n201 B.n200 585
R338 B.n202 B.n187 585
R339 B.n204 B.n203 585
R340 B.n205 B.n186 585
R341 B.n207 B.n206 585
R342 B.n208 B.n185 585
R343 B.n210 B.n209 585
R344 B.n211 B.n184 585
R345 B.n213 B.n212 585
R346 B.n214 B.n183 585
R347 B.n216 B.n215 585
R348 B.n217 B.n182 585
R349 B.n219 B.n218 585
R350 B.n220 B.n181 585
R351 B.n222 B.n221 585
R352 B.n223 B.n180 585
R353 B.n225 B.n224 585
R354 B.n226 B.n179 585
R355 B.n228 B.n227 585
R356 B.n229 B.n178 585
R357 B.n231 B.n230 585
R358 B.n232 B.n177 585
R359 B.n234 B.n233 585
R360 B.n235 B.n176 585
R361 B.n237 B.n236 585
R362 B.n238 B.n175 585
R363 B.n240 B.n239 585
R364 B.n241 B.n174 585
R365 B.n243 B.n242 585
R366 B.n242 B.n173 545.355
R367 B.n413 B.n412 545.355
R368 B.n522 B.n79 545.355
R369 B.n690 B.n689 545.355
R370 B.n317 B.t0 487.125
R371 B.n142 B.t6 487.125
R372 B.n52 B.t3 487.125
R373 B.n46 B.t9 487.125
R374 B.n745 B.n744 256.663
R375 B.n744 B.n743 235.042
R376 B.n744 B.n2 235.042
R377 B.n246 B.n173 163.367
R378 B.n247 B.n246 163.367
R379 B.n248 B.n247 163.367
R380 B.n248 B.n171 163.367
R381 B.n252 B.n171 163.367
R382 B.n253 B.n252 163.367
R383 B.n254 B.n253 163.367
R384 B.n254 B.n169 163.367
R385 B.n258 B.n169 163.367
R386 B.n259 B.n258 163.367
R387 B.n260 B.n259 163.367
R388 B.n260 B.n167 163.367
R389 B.n264 B.n167 163.367
R390 B.n265 B.n264 163.367
R391 B.n266 B.n265 163.367
R392 B.n266 B.n165 163.367
R393 B.n270 B.n165 163.367
R394 B.n271 B.n270 163.367
R395 B.n272 B.n271 163.367
R396 B.n272 B.n163 163.367
R397 B.n276 B.n163 163.367
R398 B.n277 B.n276 163.367
R399 B.n278 B.n277 163.367
R400 B.n278 B.n161 163.367
R401 B.n282 B.n161 163.367
R402 B.n283 B.n282 163.367
R403 B.n284 B.n283 163.367
R404 B.n284 B.n159 163.367
R405 B.n288 B.n159 163.367
R406 B.n289 B.n288 163.367
R407 B.n290 B.n289 163.367
R408 B.n290 B.n157 163.367
R409 B.n294 B.n157 163.367
R410 B.n295 B.n294 163.367
R411 B.n296 B.n295 163.367
R412 B.n296 B.n155 163.367
R413 B.n300 B.n155 163.367
R414 B.n301 B.n300 163.367
R415 B.n302 B.n301 163.367
R416 B.n302 B.n153 163.367
R417 B.n306 B.n153 163.367
R418 B.n307 B.n306 163.367
R419 B.n308 B.n307 163.367
R420 B.n308 B.n151 163.367
R421 B.n312 B.n151 163.367
R422 B.n313 B.n312 163.367
R423 B.n314 B.n313 163.367
R424 B.n314 B.n149 163.367
R425 B.n321 B.n149 163.367
R426 B.n322 B.n321 163.367
R427 B.n323 B.n322 163.367
R428 B.n323 B.n147 163.367
R429 B.n327 B.n147 163.367
R430 B.n328 B.n327 163.367
R431 B.n329 B.n328 163.367
R432 B.n329 B.n145 163.367
R433 B.n333 B.n145 163.367
R434 B.n334 B.n333 163.367
R435 B.n335 B.n334 163.367
R436 B.n335 B.n141 163.367
R437 B.n340 B.n141 163.367
R438 B.n341 B.n340 163.367
R439 B.n342 B.n341 163.367
R440 B.n342 B.n139 163.367
R441 B.n346 B.n139 163.367
R442 B.n347 B.n346 163.367
R443 B.n348 B.n347 163.367
R444 B.n348 B.n137 163.367
R445 B.n352 B.n137 163.367
R446 B.n353 B.n352 163.367
R447 B.n354 B.n353 163.367
R448 B.n354 B.n135 163.367
R449 B.n358 B.n135 163.367
R450 B.n359 B.n358 163.367
R451 B.n360 B.n359 163.367
R452 B.n360 B.n133 163.367
R453 B.n364 B.n133 163.367
R454 B.n365 B.n364 163.367
R455 B.n366 B.n365 163.367
R456 B.n366 B.n131 163.367
R457 B.n370 B.n131 163.367
R458 B.n371 B.n370 163.367
R459 B.n372 B.n371 163.367
R460 B.n372 B.n129 163.367
R461 B.n376 B.n129 163.367
R462 B.n377 B.n376 163.367
R463 B.n378 B.n377 163.367
R464 B.n378 B.n127 163.367
R465 B.n382 B.n127 163.367
R466 B.n383 B.n382 163.367
R467 B.n384 B.n383 163.367
R468 B.n384 B.n125 163.367
R469 B.n388 B.n125 163.367
R470 B.n389 B.n388 163.367
R471 B.n390 B.n389 163.367
R472 B.n390 B.n123 163.367
R473 B.n394 B.n123 163.367
R474 B.n395 B.n394 163.367
R475 B.n396 B.n395 163.367
R476 B.n396 B.n121 163.367
R477 B.n400 B.n121 163.367
R478 B.n401 B.n400 163.367
R479 B.n402 B.n401 163.367
R480 B.n402 B.n119 163.367
R481 B.n406 B.n119 163.367
R482 B.n407 B.n406 163.367
R483 B.n408 B.n407 163.367
R484 B.n408 B.n117 163.367
R485 B.n412 B.n117 163.367
R486 B.n522 B.n521 163.367
R487 B.n521 B.n520 163.367
R488 B.n520 B.n81 163.367
R489 B.n516 B.n81 163.367
R490 B.n516 B.n515 163.367
R491 B.n515 B.n514 163.367
R492 B.n514 B.n83 163.367
R493 B.n510 B.n83 163.367
R494 B.n510 B.n509 163.367
R495 B.n509 B.n508 163.367
R496 B.n508 B.n85 163.367
R497 B.n504 B.n85 163.367
R498 B.n504 B.n503 163.367
R499 B.n503 B.n502 163.367
R500 B.n502 B.n87 163.367
R501 B.n498 B.n87 163.367
R502 B.n498 B.n497 163.367
R503 B.n497 B.n496 163.367
R504 B.n496 B.n89 163.367
R505 B.n492 B.n89 163.367
R506 B.n492 B.n491 163.367
R507 B.n491 B.n490 163.367
R508 B.n490 B.n91 163.367
R509 B.n486 B.n91 163.367
R510 B.n486 B.n485 163.367
R511 B.n485 B.n484 163.367
R512 B.n484 B.n93 163.367
R513 B.n480 B.n93 163.367
R514 B.n480 B.n479 163.367
R515 B.n479 B.n478 163.367
R516 B.n478 B.n95 163.367
R517 B.n474 B.n95 163.367
R518 B.n474 B.n473 163.367
R519 B.n473 B.n472 163.367
R520 B.n472 B.n97 163.367
R521 B.n468 B.n97 163.367
R522 B.n468 B.n467 163.367
R523 B.n467 B.n466 163.367
R524 B.n466 B.n99 163.367
R525 B.n462 B.n99 163.367
R526 B.n462 B.n461 163.367
R527 B.n461 B.n460 163.367
R528 B.n460 B.n101 163.367
R529 B.n456 B.n101 163.367
R530 B.n456 B.n455 163.367
R531 B.n455 B.n454 163.367
R532 B.n454 B.n103 163.367
R533 B.n450 B.n103 163.367
R534 B.n450 B.n449 163.367
R535 B.n449 B.n448 163.367
R536 B.n448 B.n105 163.367
R537 B.n444 B.n105 163.367
R538 B.n444 B.n443 163.367
R539 B.n443 B.n442 163.367
R540 B.n442 B.n107 163.367
R541 B.n438 B.n107 163.367
R542 B.n438 B.n437 163.367
R543 B.n437 B.n436 163.367
R544 B.n436 B.n109 163.367
R545 B.n432 B.n109 163.367
R546 B.n432 B.n431 163.367
R547 B.n431 B.n430 163.367
R548 B.n430 B.n111 163.367
R549 B.n426 B.n111 163.367
R550 B.n426 B.n425 163.367
R551 B.n425 B.n424 163.367
R552 B.n424 B.n113 163.367
R553 B.n420 B.n113 163.367
R554 B.n420 B.n419 163.367
R555 B.n419 B.n418 163.367
R556 B.n418 B.n115 163.367
R557 B.n414 B.n115 163.367
R558 B.n414 B.n413 163.367
R559 B.n689 B.n688 163.367
R560 B.n688 B.n21 163.367
R561 B.n684 B.n21 163.367
R562 B.n684 B.n683 163.367
R563 B.n683 B.n682 163.367
R564 B.n682 B.n23 163.367
R565 B.n678 B.n23 163.367
R566 B.n678 B.n677 163.367
R567 B.n677 B.n676 163.367
R568 B.n676 B.n25 163.367
R569 B.n672 B.n25 163.367
R570 B.n672 B.n671 163.367
R571 B.n671 B.n670 163.367
R572 B.n670 B.n27 163.367
R573 B.n666 B.n27 163.367
R574 B.n666 B.n665 163.367
R575 B.n665 B.n664 163.367
R576 B.n664 B.n29 163.367
R577 B.n660 B.n29 163.367
R578 B.n660 B.n659 163.367
R579 B.n659 B.n658 163.367
R580 B.n658 B.n31 163.367
R581 B.n654 B.n31 163.367
R582 B.n654 B.n653 163.367
R583 B.n653 B.n652 163.367
R584 B.n652 B.n33 163.367
R585 B.n648 B.n33 163.367
R586 B.n648 B.n647 163.367
R587 B.n647 B.n646 163.367
R588 B.n646 B.n35 163.367
R589 B.n642 B.n35 163.367
R590 B.n642 B.n641 163.367
R591 B.n641 B.n640 163.367
R592 B.n640 B.n37 163.367
R593 B.n636 B.n37 163.367
R594 B.n636 B.n635 163.367
R595 B.n635 B.n634 163.367
R596 B.n634 B.n39 163.367
R597 B.n630 B.n39 163.367
R598 B.n630 B.n629 163.367
R599 B.n629 B.n628 163.367
R600 B.n628 B.n41 163.367
R601 B.n624 B.n41 163.367
R602 B.n624 B.n623 163.367
R603 B.n623 B.n622 163.367
R604 B.n622 B.n43 163.367
R605 B.n618 B.n43 163.367
R606 B.n618 B.n617 163.367
R607 B.n617 B.n616 163.367
R608 B.n616 B.n45 163.367
R609 B.n611 B.n45 163.367
R610 B.n611 B.n610 163.367
R611 B.n610 B.n609 163.367
R612 B.n609 B.n49 163.367
R613 B.n605 B.n49 163.367
R614 B.n605 B.n604 163.367
R615 B.n604 B.n603 163.367
R616 B.n603 B.n51 163.367
R617 B.n599 B.n51 163.367
R618 B.n599 B.n598 163.367
R619 B.n598 B.n55 163.367
R620 B.n594 B.n55 163.367
R621 B.n594 B.n593 163.367
R622 B.n593 B.n592 163.367
R623 B.n592 B.n57 163.367
R624 B.n588 B.n57 163.367
R625 B.n588 B.n587 163.367
R626 B.n587 B.n586 163.367
R627 B.n586 B.n59 163.367
R628 B.n582 B.n59 163.367
R629 B.n582 B.n581 163.367
R630 B.n581 B.n580 163.367
R631 B.n580 B.n61 163.367
R632 B.n576 B.n61 163.367
R633 B.n576 B.n575 163.367
R634 B.n575 B.n574 163.367
R635 B.n574 B.n63 163.367
R636 B.n570 B.n63 163.367
R637 B.n570 B.n569 163.367
R638 B.n569 B.n568 163.367
R639 B.n568 B.n65 163.367
R640 B.n564 B.n65 163.367
R641 B.n564 B.n563 163.367
R642 B.n563 B.n562 163.367
R643 B.n562 B.n67 163.367
R644 B.n558 B.n67 163.367
R645 B.n558 B.n557 163.367
R646 B.n557 B.n556 163.367
R647 B.n556 B.n69 163.367
R648 B.n552 B.n69 163.367
R649 B.n552 B.n551 163.367
R650 B.n551 B.n550 163.367
R651 B.n550 B.n71 163.367
R652 B.n546 B.n71 163.367
R653 B.n546 B.n545 163.367
R654 B.n545 B.n544 163.367
R655 B.n544 B.n73 163.367
R656 B.n540 B.n73 163.367
R657 B.n540 B.n539 163.367
R658 B.n539 B.n538 163.367
R659 B.n538 B.n75 163.367
R660 B.n534 B.n75 163.367
R661 B.n534 B.n533 163.367
R662 B.n533 B.n532 163.367
R663 B.n532 B.n77 163.367
R664 B.n528 B.n77 163.367
R665 B.n528 B.n527 163.367
R666 B.n527 B.n526 163.367
R667 B.n526 B.n79 163.367
R668 B.n690 B.n19 163.367
R669 B.n694 B.n19 163.367
R670 B.n695 B.n694 163.367
R671 B.n696 B.n695 163.367
R672 B.n696 B.n17 163.367
R673 B.n700 B.n17 163.367
R674 B.n701 B.n700 163.367
R675 B.n702 B.n701 163.367
R676 B.n702 B.n15 163.367
R677 B.n706 B.n15 163.367
R678 B.n707 B.n706 163.367
R679 B.n708 B.n707 163.367
R680 B.n708 B.n13 163.367
R681 B.n712 B.n13 163.367
R682 B.n713 B.n712 163.367
R683 B.n714 B.n713 163.367
R684 B.n714 B.n11 163.367
R685 B.n718 B.n11 163.367
R686 B.n719 B.n718 163.367
R687 B.n720 B.n719 163.367
R688 B.n720 B.n9 163.367
R689 B.n724 B.n9 163.367
R690 B.n725 B.n724 163.367
R691 B.n726 B.n725 163.367
R692 B.n726 B.n7 163.367
R693 B.n730 B.n7 163.367
R694 B.n731 B.n730 163.367
R695 B.n732 B.n731 163.367
R696 B.n732 B.n5 163.367
R697 B.n736 B.n5 163.367
R698 B.n737 B.n736 163.367
R699 B.n738 B.n737 163.367
R700 B.n738 B.n3 163.367
R701 B.n742 B.n3 163.367
R702 B.n743 B.n742 163.367
R703 B.n192 B.n2 163.367
R704 B.n193 B.n192 163.367
R705 B.n194 B.n193 163.367
R706 B.n194 B.n189 163.367
R707 B.n198 B.n189 163.367
R708 B.n199 B.n198 163.367
R709 B.n200 B.n199 163.367
R710 B.n200 B.n187 163.367
R711 B.n204 B.n187 163.367
R712 B.n205 B.n204 163.367
R713 B.n206 B.n205 163.367
R714 B.n206 B.n185 163.367
R715 B.n210 B.n185 163.367
R716 B.n211 B.n210 163.367
R717 B.n212 B.n211 163.367
R718 B.n212 B.n183 163.367
R719 B.n216 B.n183 163.367
R720 B.n217 B.n216 163.367
R721 B.n218 B.n217 163.367
R722 B.n218 B.n181 163.367
R723 B.n222 B.n181 163.367
R724 B.n223 B.n222 163.367
R725 B.n224 B.n223 163.367
R726 B.n224 B.n179 163.367
R727 B.n228 B.n179 163.367
R728 B.n229 B.n228 163.367
R729 B.n230 B.n229 163.367
R730 B.n230 B.n177 163.367
R731 B.n234 B.n177 163.367
R732 B.n235 B.n234 163.367
R733 B.n236 B.n235 163.367
R734 B.n236 B.n175 163.367
R735 B.n240 B.n175 163.367
R736 B.n241 B.n240 163.367
R737 B.n242 B.n241 163.367
R738 B.n142 B.t7 138.754
R739 B.n52 B.t5 138.754
R740 B.n317 B.t1 138.734
R741 B.n46 B.t11 138.734
R742 B.n143 B.t8 107.529
R743 B.n53 B.t4 107.529
R744 B.n318 B.t2 107.51
R745 B.n47 B.t10 107.51
R746 B.n319 B.n318 59.5399
R747 B.n337 B.n143 59.5399
R748 B.n54 B.n53 59.5399
R749 B.n614 B.n47 59.5399
R750 B.n691 B.n20 35.4346
R751 B.n524 B.n523 35.4346
R752 B.n411 B.n116 35.4346
R753 B.n244 B.n243 35.4346
R754 B.n318 B.n317 31.2247
R755 B.n143 B.n142 31.2247
R756 B.n53 B.n52 31.2247
R757 B.n47 B.n46 31.2247
R758 B B.n745 18.0485
R759 B.n692 B.n691 10.6151
R760 B.n693 B.n692 10.6151
R761 B.n693 B.n18 10.6151
R762 B.n697 B.n18 10.6151
R763 B.n698 B.n697 10.6151
R764 B.n699 B.n698 10.6151
R765 B.n699 B.n16 10.6151
R766 B.n703 B.n16 10.6151
R767 B.n704 B.n703 10.6151
R768 B.n705 B.n704 10.6151
R769 B.n705 B.n14 10.6151
R770 B.n709 B.n14 10.6151
R771 B.n710 B.n709 10.6151
R772 B.n711 B.n710 10.6151
R773 B.n711 B.n12 10.6151
R774 B.n715 B.n12 10.6151
R775 B.n716 B.n715 10.6151
R776 B.n717 B.n716 10.6151
R777 B.n717 B.n10 10.6151
R778 B.n721 B.n10 10.6151
R779 B.n722 B.n721 10.6151
R780 B.n723 B.n722 10.6151
R781 B.n723 B.n8 10.6151
R782 B.n727 B.n8 10.6151
R783 B.n728 B.n727 10.6151
R784 B.n729 B.n728 10.6151
R785 B.n729 B.n6 10.6151
R786 B.n733 B.n6 10.6151
R787 B.n734 B.n733 10.6151
R788 B.n735 B.n734 10.6151
R789 B.n735 B.n4 10.6151
R790 B.n739 B.n4 10.6151
R791 B.n740 B.n739 10.6151
R792 B.n741 B.n740 10.6151
R793 B.n741 B.n0 10.6151
R794 B.n687 B.n20 10.6151
R795 B.n687 B.n686 10.6151
R796 B.n686 B.n685 10.6151
R797 B.n685 B.n22 10.6151
R798 B.n681 B.n22 10.6151
R799 B.n681 B.n680 10.6151
R800 B.n680 B.n679 10.6151
R801 B.n679 B.n24 10.6151
R802 B.n675 B.n24 10.6151
R803 B.n675 B.n674 10.6151
R804 B.n674 B.n673 10.6151
R805 B.n673 B.n26 10.6151
R806 B.n669 B.n26 10.6151
R807 B.n669 B.n668 10.6151
R808 B.n668 B.n667 10.6151
R809 B.n667 B.n28 10.6151
R810 B.n663 B.n28 10.6151
R811 B.n663 B.n662 10.6151
R812 B.n662 B.n661 10.6151
R813 B.n661 B.n30 10.6151
R814 B.n657 B.n30 10.6151
R815 B.n657 B.n656 10.6151
R816 B.n656 B.n655 10.6151
R817 B.n655 B.n32 10.6151
R818 B.n651 B.n32 10.6151
R819 B.n651 B.n650 10.6151
R820 B.n650 B.n649 10.6151
R821 B.n649 B.n34 10.6151
R822 B.n645 B.n34 10.6151
R823 B.n645 B.n644 10.6151
R824 B.n644 B.n643 10.6151
R825 B.n643 B.n36 10.6151
R826 B.n639 B.n36 10.6151
R827 B.n639 B.n638 10.6151
R828 B.n638 B.n637 10.6151
R829 B.n637 B.n38 10.6151
R830 B.n633 B.n38 10.6151
R831 B.n633 B.n632 10.6151
R832 B.n632 B.n631 10.6151
R833 B.n631 B.n40 10.6151
R834 B.n627 B.n40 10.6151
R835 B.n627 B.n626 10.6151
R836 B.n626 B.n625 10.6151
R837 B.n625 B.n42 10.6151
R838 B.n621 B.n42 10.6151
R839 B.n621 B.n620 10.6151
R840 B.n620 B.n619 10.6151
R841 B.n619 B.n44 10.6151
R842 B.n615 B.n44 10.6151
R843 B.n613 B.n612 10.6151
R844 B.n612 B.n48 10.6151
R845 B.n608 B.n48 10.6151
R846 B.n608 B.n607 10.6151
R847 B.n607 B.n606 10.6151
R848 B.n606 B.n50 10.6151
R849 B.n602 B.n50 10.6151
R850 B.n602 B.n601 10.6151
R851 B.n601 B.n600 10.6151
R852 B.n597 B.n596 10.6151
R853 B.n596 B.n595 10.6151
R854 B.n595 B.n56 10.6151
R855 B.n591 B.n56 10.6151
R856 B.n591 B.n590 10.6151
R857 B.n590 B.n589 10.6151
R858 B.n589 B.n58 10.6151
R859 B.n585 B.n58 10.6151
R860 B.n585 B.n584 10.6151
R861 B.n584 B.n583 10.6151
R862 B.n583 B.n60 10.6151
R863 B.n579 B.n60 10.6151
R864 B.n579 B.n578 10.6151
R865 B.n578 B.n577 10.6151
R866 B.n577 B.n62 10.6151
R867 B.n573 B.n62 10.6151
R868 B.n573 B.n572 10.6151
R869 B.n572 B.n571 10.6151
R870 B.n571 B.n64 10.6151
R871 B.n567 B.n64 10.6151
R872 B.n567 B.n566 10.6151
R873 B.n566 B.n565 10.6151
R874 B.n565 B.n66 10.6151
R875 B.n561 B.n66 10.6151
R876 B.n561 B.n560 10.6151
R877 B.n560 B.n559 10.6151
R878 B.n559 B.n68 10.6151
R879 B.n555 B.n68 10.6151
R880 B.n555 B.n554 10.6151
R881 B.n554 B.n553 10.6151
R882 B.n553 B.n70 10.6151
R883 B.n549 B.n70 10.6151
R884 B.n549 B.n548 10.6151
R885 B.n548 B.n547 10.6151
R886 B.n547 B.n72 10.6151
R887 B.n543 B.n72 10.6151
R888 B.n543 B.n542 10.6151
R889 B.n542 B.n541 10.6151
R890 B.n541 B.n74 10.6151
R891 B.n537 B.n74 10.6151
R892 B.n537 B.n536 10.6151
R893 B.n536 B.n535 10.6151
R894 B.n535 B.n76 10.6151
R895 B.n531 B.n76 10.6151
R896 B.n531 B.n530 10.6151
R897 B.n530 B.n529 10.6151
R898 B.n529 B.n78 10.6151
R899 B.n525 B.n78 10.6151
R900 B.n525 B.n524 10.6151
R901 B.n523 B.n80 10.6151
R902 B.n519 B.n80 10.6151
R903 B.n519 B.n518 10.6151
R904 B.n518 B.n517 10.6151
R905 B.n517 B.n82 10.6151
R906 B.n513 B.n82 10.6151
R907 B.n513 B.n512 10.6151
R908 B.n512 B.n511 10.6151
R909 B.n511 B.n84 10.6151
R910 B.n507 B.n84 10.6151
R911 B.n507 B.n506 10.6151
R912 B.n506 B.n505 10.6151
R913 B.n505 B.n86 10.6151
R914 B.n501 B.n86 10.6151
R915 B.n501 B.n500 10.6151
R916 B.n500 B.n499 10.6151
R917 B.n499 B.n88 10.6151
R918 B.n495 B.n88 10.6151
R919 B.n495 B.n494 10.6151
R920 B.n494 B.n493 10.6151
R921 B.n493 B.n90 10.6151
R922 B.n489 B.n90 10.6151
R923 B.n489 B.n488 10.6151
R924 B.n488 B.n487 10.6151
R925 B.n487 B.n92 10.6151
R926 B.n483 B.n92 10.6151
R927 B.n483 B.n482 10.6151
R928 B.n482 B.n481 10.6151
R929 B.n481 B.n94 10.6151
R930 B.n477 B.n94 10.6151
R931 B.n477 B.n476 10.6151
R932 B.n476 B.n475 10.6151
R933 B.n475 B.n96 10.6151
R934 B.n471 B.n96 10.6151
R935 B.n471 B.n470 10.6151
R936 B.n470 B.n469 10.6151
R937 B.n469 B.n98 10.6151
R938 B.n465 B.n98 10.6151
R939 B.n465 B.n464 10.6151
R940 B.n464 B.n463 10.6151
R941 B.n463 B.n100 10.6151
R942 B.n459 B.n100 10.6151
R943 B.n459 B.n458 10.6151
R944 B.n458 B.n457 10.6151
R945 B.n457 B.n102 10.6151
R946 B.n453 B.n102 10.6151
R947 B.n453 B.n452 10.6151
R948 B.n452 B.n451 10.6151
R949 B.n451 B.n104 10.6151
R950 B.n447 B.n104 10.6151
R951 B.n447 B.n446 10.6151
R952 B.n446 B.n445 10.6151
R953 B.n445 B.n106 10.6151
R954 B.n441 B.n106 10.6151
R955 B.n441 B.n440 10.6151
R956 B.n440 B.n439 10.6151
R957 B.n439 B.n108 10.6151
R958 B.n435 B.n108 10.6151
R959 B.n435 B.n434 10.6151
R960 B.n434 B.n433 10.6151
R961 B.n433 B.n110 10.6151
R962 B.n429 B.n110 10.6151
R963 B.n429 B.n428 10.6151
R964 B.n428 B.n427 10.6151
R965 B.n427 B.n112 10.6151
R966 B.n423 B.n112 10.6151
R967 B.n423 B.n422 10.6151
R968 B.n422 B.n421 10.6151
R969 B.n421 B.n114 10.6151
R970 B.n417 B.n114 10.6151
R971 B.n417 B.n416 10.6151
R972 B.n416 B.n415 10.6151
R973 B.n415 B.n116 10.6151
R974 B.n191 B.n1 10.6151
R975 B.n191 B.n190 10.6151
R976 B.n195 B.n190 10.6151
R977 B.n196 B.n195 10.6151
R978 B.n197 B.n196 10.6151
R979 B.n197 B.n188 10.6151
R980 B.n201 B.n188 10.6151
R981 B.n202 B.n201 10.6151
R982 B.n203 B.n202 10.6151
R983 B.n203 B.n186 10.6151
R984 B.n207 B.n186 10.6151
R985 B.n208 B.n207 10.6151
R986 B.n209 B.n208 10.6151
R987 B.n209 B.n184 10.6151
R988 B.n213 B.n184 10.6151
R989 B.n214 B.n213 10.6151
R990 B.n215 B.n214 10.6151
R991 B.n215 B.n182 10.6151
R992 B.n219 B.n182 10.6151
R993 B.n220 B.n219 10.6151
R994 B.n221 B.n220 10.6151
R995 B.n221 B.n180 10.6151
R996 B.n225 B.n180 10.6151
R997 B.n226 B.n225 10.6151
R998 B.n227 B.n226 10.6151
R999 B.n227 B.n178 10.6151
R1000 B.n231 B.n178 10.6151
R1001 B.n232 B.n231 10.6151
R1002 B.n233 B.n232 10.6151
R1003 B.n233 B.n176 10.6151
R1004 B.n237 B.n176 10.6151
R1005 B.n238 B.n237 10.6151
R1006 B.n239 B.n238 10.6151
R1007 B.n239 B.n174 10.6151
R1008 B.n243 B.n174 10.6151
R1009 B.n245 B.n244 10.6151
R1010 B.n245 B.n172 10.6151
R1011 B.n249 B.n172 10.6151
R1012 B.n250 B.n249 10.6151
R1013 B.n251 B.n250 10.6151
R1014 B.n251 B.n170 10.6151
R1015 B.n255 B.n170 10.6151
R1016 B.n256 B.n255 10.6151
R1017 B.n257 B.n256 10.6151
R1018 B.n257 B.n168 10.6151
R1019 B.n261 B.n168 10.6151
R1020 B.n262 B.n261 10.6151
R1021 B.n263 B.n262 10.6151
R1022 B.n263 B.n166 10.6151
R1023 B.n267 B.n166 10.6151
R1024 B.n268 B.n267 10.6151
R1025 B.n269 B.n268 10.6151
R1026 B.n269 B.n164 10.6151
R1027 B.n273 B.n164 10.6151
R1028 B.n274 B.n273 10.6151
R1029 B.n275 B.n274 10.6151
R1030 B.n275 B.n162 10.6151
R1031 B.n279 B.n162 10.6151
R1032 B.n280 B.n279 10.6151
R1033 B.n281 B.n280 10.6151
R1034 B.n281 B.n160 10.6151
R1035 B.n285 B.n160 10.6151
R1036 B.n286 B.n285 10.6151
R1037 B.n287 B.n286 10.6151
R1038 B.n287 B.n158 10.6151
R1039 B.n291 B.n158 10.6151
R1040 B.n292 B.n291 10.6151
R1041 B.n293 B.n292 10.6151
R1042 B.n293 B.n156 10.6151
R1043 B.n297 B.n156 10.6151
R1044 B.n298 B.n297 10.6151
R1045 B.n299 B.n298 10.6151
R1046 B.n299 B.n154 10.6151
R1047 B.n303 B.n154 10.6151
R1048 B.n304 B.n303 10.6151
R1049 B.n305 B.n304 10.6151
R1050 B.n305 B.n152 10.6151
R1051 B.n309 B.n152 10.6151
R1052 B.n310 B.n309 10.6151
R1053 B.n311 B.n310 10.6151
R1054 B.n311 B.n150 10.6151
R1055 B.n315 B.n150 10.6151
R1056 B.n316 B.n315 10.6151
R1057 B.n320 B.n316 10.6151
R1058 B.n324 B.n148 10.6151
R1059 B.n325 B.n324 10.6151
R1060 B.n326 B.n325 10.6151
R1061 B.n326 B.n146 10.6151
R1062 B.n330 B.n146 10.6151
R1063 B.n331 B.n330 10.6151
R1064 B.n332 B.n331 10.6151
R1065 B.n332 B.n144 10.6151
R1066 B.n336 B.n144 10.6151
R1067 B.n339 B.n338 10.6151
R1068 B.n339 B.n140 10.6151
R1069 B.n343 B.n140 10.6151
R1070 B.n344 B.n343 10.6151
R1071 B.n345 B.n344 10.6151
R1072 B.n345 B.n138 10.6151
R1073 B.n349 B.n138 10.6151
R1074 B.n350 B.n349 10.6151
R1075 B.n351 B.n350 10.6151
R1076 B.n351 B.n136 10.6151
R1077 B.n355 B.n136 10.6151
R1078 B.n356 B.n355 10.6151
R1079 B.n357 B.n356 10.6151
R1080 B.n357 B.n134 10.6151
R1081 B.n361 B.n134 10.6151
R1082 B.n362 B.n361 10.6151
R1083 B.n363 B.n362 10.6151
R1084 B.n363 B.n132 10.6151
R1085 B.n367 B.n132 10.6151
R1086 B.n368 B.n367 10.6151
R1087 B.n369 B.n368 10.6151
R1088 B.n369 B.n130 10.6151
R1089 B.n373 B.n130 10.6151
R1090 B.n374 B.n373 10.6151
R1091 B.n375 B.n374 10.6151
R1092 B.n375 B.n128 10.6151
R1093 B.n379 B.n128 10.6151
R1094 B.n380 B.n379 10.6151
R1095 B.n381 B.n380 10.6151
R1096 B.n381 B.n126 10.6151
R1097 B.n385 B.n126 10.6151
R1098 B.n386 B.n385 10.6151
R1099 B.n387 B.n386 10.6151
R1100 B.n387 B.n124 10.6151
R1101 B.n391 B.n124 10.6151
R1102 B.n392 B.n391 10.6151
R1103 B.n393 B.n392 10.6151
R1104 B.n393 B.n122 10.6151
R1105 B.n397 B.n122 10.6151
R1106 B.n398 B.n397 10.6151
R1107 B.n399 B.n398 10.6151
R1108 B.n399 B.n120 10.6151
R1109 B.n403 B.n120 10.6151
R1110 B.n404 B.n403 10.6151
R1111 B.n405 B.n404 10.6151
R1112 B.n405 B.n118 10.6151
R1113 B.n409 B.n118 10.6151
R1114 B.n410 B.n409 10.6151
R1115 B.n411 B.n410 10.6151
R1116 B.n615 B.n614 9.36635
R1117 B.n597 B.n54 9.36635
R1118 B.n320 B.n319 9.36635
R1119 B.n338 B.n337 9.36635
R1120 B.n745 B.n0 8.11757
R1121 B.n745 B.n1 8.11757
R1122 B.n614 B.n613 1.24928
R1123 B.n600 B.n54 1.24928
R1124 B.n319 B.n148 1.24928
R1125 B.n337 B.n336 1.24928
R1126 VP.n14 VP.t4 310.767
R1127 VP.n3 VP.t9 282.611
R1128 VP.n7 VP.t0 282.611
R1129 VP.n5 VP.t7 282.611
R1130 VP.n48 VP.t1 282.611
R1131 VP.n55 VP.t6 282.611
R1132 VP.n11 VP.t5 282.611
R1133 VP.n31 VP.t2 282.611
R1134 VP.n24 VP.t3 282.611
R1135 VP.n13 VP.t8 282.611
R1136 VP.n33 VP.n7 175.002
R1137 VP.n56 VP.n55 175.002
R1138 VP.n32 VP.n31 175.002
R1139 VP.n16 VP.n15 161.3
R1140 VP.n17 VP.n12 161.3
R1141 VP.n19 VP.n18 161.3
R1142 VP.n20 VP.n11 161.3
R1143 VP.n22 VP.n21 161.3
R1144 VP.n23 VP.n10 161.3
R1145 VP.n26 VP.n25 161.3
R1146 VP.n27 VP.n9 161.3
R1147 VP.n29 VP.n28 161.3
R1148 VP.n30 VP.n8 161.3
R1149 VP.n54 VP.n0 161.3
R1150 VP.n53 VP.n52 161.3
R1151 VP.n51 VP.n1 161.3
R1152 VP.n50 VP.n49 161.3
R1153 VP.n47 VP.n2 161.3
R1154 VP.n46 VP.n45 161.3
R1155 VP.n44 VP.n3 161.3
R1156 VP.n43 VP.n42 161.3
R1157 VP.n41 VP.n4 161.3
R1158 VP.n40 VP.n39 161.3
R1159 VP.n38 VP.n37 161.3
R1160 VP.n36 VP.n6 161.3
R1161 VP.n35 VP.n34 161.3
R1162 VP.n14 VP.n13 59.7169
R1163 VP.n42 VP.n41 56.5193
R1164 VP.n47 VP.n46 56.5193
R1165 VP.n23 VP.n22 56.5193
R1166 VP.n18 VP.n17 56.5193
R1167 VP.n37 VP.n36 48.7492
R1168 VP.n53 VP.n1 48.7492
R1169 VP.n29 VP.n9 48.7492
R1170 VP.n33 VP.n32 48.1028
R1171 VP.n36 VP.n35 32.2376
R1172 VP.n54 VP.n53 32.2376
R1173 VP.n30 VP.n29 32.2376
R1174 VP.n15 VP.n14 27.4893
R1175 VP.n41 VP.n40 24.4675
R1176 VP.n42 VP.n3 24.4675
R1177 VP.n46 VP.n3 24.4675
R1178 VP.n49 VP.n47 24.4675
R1179 VP.n25 VP.n23 24.4675
R1180 VP.n18 VP.n11 24.4675
R1181 VP.n22 VP.n11 24.4675
R1182 VP.n17 VP.n16 24.4675
R1183 VP.n37 VP.n5 19.0848
R1184 VP.n48 VP.n1 19.0848
R1185 VP.n24 VP.n9 19.0848
R1186 VP.n35 VP.n7 10.766
R1187 VP.n55 VP.n54 10.766
R1188 VP.n31 VP.n30 10.766
R1189 VP.n40 VP.n5 5.38324
R1190 VP.n49 VP.n48 5.38324
R1191 VP.n25 VP.n24 5.38324
R1192 VP.n16 VP.n13 5.38324
R1193 VP.n15 VP.n12 0.189894
R1194 VP.n19 VP.n12 0.189894
R1195 VP.n20 VP.n19 0.189894
R1196 VP.n21 VP.n20 0.189894
R1197 VP.n21 VP.n10 0.189894
R1198 VP.n26 VP.n10 0.189894
R1199 VP.n27 VP.n26 0.189894
R1200 VP.n28 VP.n27 0.189894
R1201 VP.n28 VP.n8 0.189894
R1202 VP.n32 VP.n8 0.189894
R1203 VP.n34 VP.n33 0.189894
R1204 VP.n34 VP.n6 0.189894
R1205 VP.n38 VP.n6 0.189894
R1206 VP.n39 VP.n38 0.189894
R1207 VP.n39 VP.n4 0.189894
R1208 VP.n43 VP.n4 0.189894
R1209 VP.n44 VP.n43 0.189894
R1210 VP.n45 VP.n44 0.189894
R1211 VP.n45 VP.n2 0.189894
R1212 VP.n50 VP.n2 0.189894
R1213 VP.n51 VP.n50 0.189894
R1214 VP.n52 VP.n51 0.189894
R1215 VP.n52 VP.n0 0.189894
R1216 VP.n56 VP.n0 0.189894
R1217 VP VP.n56 0.0516364
R1218 VTAIL.n11 VTAIL.t1 56.1859
R1219 VTAIL.n17 VTAIL.t6 56.1856
R1220 VTAIL.n2 VTAIL.t12 56.1856
R1221 VTAIL.n16 VTAIL.t15 56.1856
R1222 VTAIL.n15 VTAIL.n14 54.0203
R1223 VTAIL.n13 VTAIL.n12 54.0203
R1224 VTAIL.n10 VTAIL.n9 54.0203
R1225 VTAIL.n8 VTAIL.n7 54.0203
R1226 VTAIL.n19 VTAIL.n18 54.0201
R1227 VTAIL.n1 VTAIL.n0 54.0201
R1228 VTAIL.n4 VTAIL.n3 54.0201
R1229 VTAIL.n6 VTAIL.n5 54.0201
R1230 VTAIL.n8 VTAIL.n6 28.0824
R1231 VTAIL.n17 VTAIL.n16 26.6945
R1232 VTAIL.n18 VTAIL.t9 2.16606
R1233 VTAIL.n18 VTAIL.t3 2.16606
R1234 VTAIL.n0 VTAIL.t2 2.16606
R1235 VTAIL.n0 VTAIL.t7 2.16606
R1236 VTAIL.n3 VTAIL.t10 2.16606
R1237 VTAIL.n3 VTAIL.t11 2.16606
R1238 VTAIL.n5 VTAIL.t14 2.16606
R1239 VTAIL.n5 VTAIL.t16 2.16606
R1240 VTAIL.n14 VTAIL.t17 2.16606
R1241 VTAIL.n14 VTAIL.t19 2.16606
R1242 VTAIL.n12 VTAIL.t18 2.16606
R1243 VTAIL.n12 VTAIL.t13 2.16606
R1244 VTAIL.n9 VTAIL.t0 2.16606
R1245 VTAIL.n9 VTAIL.t4 2.16606
R1246 VTAIL.n7 VTAIL.t5 2.16606
R1247 VTAIL.n7 VTAIL.t8 2.16606
R1248 VTAIL.n10 VTAIL.n8 1.38843
R1249 VTAIL.n11 VTAIL.n10 1.38843
R1250 VTAIL.n15 VTAIL.n13 1.38843
R1251 VTAIL.n16 VTAIL.n15 1.38843
R1252 VTAIL.n6 VTAIL.n4 1.38843
R1253 VTAIL.n4 VTAIL.n2 1.38843
R1254 VTAIL.n19 VTAIL.n17 1.38843
R1255 VTAIL.n13 VTAIL.n11 1.16429
R1256 VTAIL.n2 VTAIL.n1 1.16429
R1257 VTAIL VTAIL.n1 1.09964
R1258 VTAIL VTAIL.n19 0.289293
R1259 VDD1.n1 VDD1.t5 74.2526
R1260 VDD1.n3 VDD1.t9 74.2523
R1261 VDD1.n5 VDD1.n4 71.6844
R1262 VDD1.n1 VDD1.n0 70.6991
R1263 VDD1.n7 VDD1.n6 70.6989
R1264 VDD1.n3 VDD1.n2 70.6988
R1265 VDD1.n7 VDD1.n5 44.5246
R1266 VDD1.n6 VDD1.t6 2.16606
R1267 VDD1.n6 VDD1.t7 2.16606
R1268 VDD1.n0 VDD1.t1 2.16606
R1269 VDD1.n0 VDD1.t4 2.16606
R1270 VDD1.n4 VDD1.t8 2.16606
R1271 VDD1.n4 VDD1.t3 2.16606
R1272 VDD1.n2 VDD1.t2 2.16606
R1273 VDD1.n2 VDD1.t0 2.16606
R1274 VDD1 VDD1.n7 0.983259
R1275 VDD1 VDD1.n1 0.405672
R1276 VDD1.n5 VDD1.n3 0.292137
R1277 VN.n6 VN.t8 310.767
R1278 VN.n32 VN.t3 310.767
R1279 VN.n3 VN.t9 282.611
R1280 VN.n5 VN.t7 282.611
R1281 VN.n16 VN.t6 282.611
R1282 VN.n23 VN.t0 282.611
R1283 VN.n29 VN.t1 282.611
R1284 VN.n31 VN.t2 282.611
R1285 VN.n28 VN.t5 282.611
R1286 VN.n48 VN.t4 282.611
R1287 VN.n24 VN.n23 175.002
R1288 VN.n49 VN.n48 175.002
R1289 VN.n47 VN.n25 161.3
R1290 VN.n46 VN.n45 161.3
R1291 VN.n44 VN.n26 161.3
R1292 VN.n43 VN.n42 161.3
R1293 VN.n41 VN.n27 161.3
R1294 VN.n40 VN.n39 161.3
R1295 VN.n38 VN.n29 161.3
R1296 VN.n37 VN.n36 161.3
R1297 VN.n35 VN.n30 161.3
R1298 VN.n34 VN.n33 161.3
R1299 VN.n22 VN.n0 161.3
R1300 VN.n21 VN.n20 161.3
R1301 VN.n19 VN.n1 161.3
R1302 VN.n18 VN.n17 161.3
R1303 VN.n15 VN.n2 161.3
R1304 VN.n14 VN.n13 161.3
R1305 VN.n12 VN.n3 161.3
R1306 VN.n11 VN.n10 161.3
R1307 VN.n9 VN.n4 161.3
R1308 VN.n8 VN.n7 161.3
R1309 VN.n6 VN.n5 59.7169
R1310 VN.n32 VN.n31 59.7169
R1311 VN.n10 VN.n9 56.5193
R1312 VN.n15 VN.n14 56.5193
R1313 VN.n36 VN.n35 56.5193
R1314 VN.n41 VN.n40 56.5193
R1315 VN.n21 VN.n1 48.7492
R1316 VN.n46 VN.n26 48.7492
R1317 VN VN.n49 48.4835
R1318 VN.n22 VN.n21 32.2376
R1319 VN.n47 VN.n46 32.2376
R1320 VN.n33 VN.n32 27.4893
R1321 VN.n7 VN.n6 27.4893
R1322 VN.n9 VN.n8 24.4675
R1323 VN.n10 VN.n3 24.4675
R1324 VN.n14 VN.n3 24.4675
R1325 VN.n17 VN.n15 24.4675
R1326 VN.n35 VN.n34 24.4675
R1327 VN.n40 VN.n29 24.4675
R1328 VN.n36 VN.n29 24.4675
R1329 VN.n42 VN.n41 24.4675
R1330 VN.n16 VN.n1 19.0848
R1331 VN.n28 VN.n26 19.0848
R1332 VN.n23 VN.n22 10.766
R1333 VN.n48 VN.n47 10.766
R1334 VN.n8 VN.n5 5.38324
R1335 VN.n17 VN.n16 5.38324
R1336 VN.n34 VN.n31 5.38324
R1337 VN.n42 VN.n28 5.38324
R1338 VN.n49 VN.n25 0.189894
R1339 VN.n45 VN.n25 0.189894
R1340 VN.n45 VN.n44 0.189894
R1341 VN.n44 VN.n43 0.189894
R1342 VN.n43 VN.n27 0.189894
R1343 VN.n39 VN.n27 0.189894
R1344 VN.n39 VN.n38 0.189894
R1345 VN.n38 VN.n37 0.189894
R1346 VN.n37 VN.n30 0.189894
R1347 VN.n33 VN.n30 0.189894
R1348 VN.n7 VN.n4 0.189894
R1349 VN.n11 VN.n4 0.189894
R1350 VN.n12 VN.n11 0.189894
R1351 VN.n13 VN.n12 0.189894
R1352 VN.n13 VN.n2 0.189894
R1353 VN.n18 VN.n2 0.189894
R1354 VN.n19 VN.n18 0.189894
R1355 VN.n20 VN.n19 0.189894
R1356 VN.n20 VN.n0 0.189894
R1357 VN.n24 VN.n0 0.189894
R1358 VN VN.n24 0.0516364
R1359 VDD2.n1 VDD2.t1 74.2523
R1360 VDD2.n4 VDD2.t5 72.8647
R1361 VDD2.n3 VDD2.n2 71.6844
R1362 VDD2 VDD2.n7 71.6817
R1363 VDD2.n6 VDD2.n5 70.6991
R1364 VDD2.n1 VDD2.n0 70.6988
R1365 VDD2.n4 VDD2.n3 43.2476
R1366 VDD2.n7 VDD2.t7 2.16606
R1367 VDD2.n7 VDD2.t6 2.16606
R1368 VDD2.n5 VDD2.t4 2.16606
R1369 VDD2.n5 VDD2.t8 2.16606
R1370 VDD2.n2 VDD2.t3 2.16606
R1371 VDD2.n2 VDD2.t9 2.16606
R1372 VDD2.n0 VDD2.t2 2.16606
R1373 VDD2.n0 VDD2.t0 2.16606
R1374 VDD2.n6 VDD2.n4 1.38843
R1375 VDD2 VDD2.n6 0.405672
R1376 VDD2.n3 VDD2.n1 0.292137
C0 VTAIL B 3.684f
C1 VN VDD1 0.150329f
C2 B VDD1 2.17743f
C3 w_n2902_n3970# VP 6.2412f
C4 VDD2 VP 0.415711f
C5 w_n2902_n3970# VDD2 2.57397f
C6 VTAIL VP 10.8372f
C7 w_n2902_n3970# VTAIL 3.50361f
C8 VTAIL VDD2 13.451799f
C9 B VN 0.98264f
C10 VP VDD1 11.1073f
C11 w_n2902_n3970# VDD1 2.49898f
C12 VDD2 VDD1 1.3319f
C13 VTAIL VDD1 13.413099f
C14 VN VP 7.01256f
C15 w_n2902_n3970# VN 5.86744f
C16 VDD2 VN 10.846901f
C17 VTAIL VN 10.822599f
C18 B VP 1.60384f
C19 w_n2902_n3970# B 9.17074f
C20 B VDD2 2.24395f
C21 VDD2 VSUBS 1.753283f
C22 VDD1 VSUBS 1.491155f
C23 VTAIL VSUBS 1.072642f
C24 VN VSUBS 5.79945f
C25 VP VSUBS 2.657897f
C26 B VSUBS 3.984792f
C27 w_n2902_n3970# VSUBS 0.141281p
C28 VDD2.t1 VSUBS 3.41239f
C29 VDD2.t2 VSUBS 0.32213f
C30 VDD2.t0 VSUBS 0.32213f
C31 VDD2.n0 VSUBS 2.61412f
C32 VDD2.n1 VSUBS 1.402f
C33 VDD2.t3 VSUBS 0.32213f
C34 VDD2.t9 VSUBS 0.32213f
C35 VDD2.n2 VSUBS 2.62429f
C36 VDD2.n3 VSUBS 2.89754f
C37 VDD2.t5 VSUBS 3.39843f
C38 VDD2.n4 VSUBS 3.40896f
C39 VDD2.t4 VSUBS 0.32213f
C40 VDD2.t8 VSUBS 0.32213f
C41 VDD2.n5 VSUBS 2.61413f
C42 VDD2.n6 VSUBS 0.67701f
C43 VDD2.t7 VSUBS 0.32213f
C44 VDD2.t6 VSUBS 0.32213f
C45 VDD2.n7 VSUBS 2.62424f
C46 VN.n0 VSUBS 0.038765f
C47 VN.t0 VSUBS 2.04088f
C48 VN.n1 VSUBS 0.064401f
C49 VN.n2 VSUBS 0.038765f
C50 VN.t9 VSUBS 2.04088f
C51 VN.n3 VSUBS 0.767994f
C52 VN.n4 VSUBS 0.038765f
C53 VN.t7 VSUBS 2.04088f
C54 VN.n5 VSUBS 0.784152f
C55 VN.t8 VSUBS 2.11804f
C56 VN.n6 VSUBS 0.827632f
C57 VN.n7 VSUBS 0.202833f
C58 VN.n8 VSUBS 0.044426f
C59 VN.n9 VSUBS 0.050653f
C60 VN.n10 VSUBS 0.062535f
C61 VN.n11 VSUBS 0.038765f
C62 VN.n12 VSUBS 0.038765f
C63 VN.n13 VSUBS 0.038765f
C64 VN.n14 VSUBS 0.062535f
C65 VN.n15 VSUBS 0.050653f
C66 VN.t6 VSUBS 2.04088f
C67 VN.n16 VSUBS 0.731415f
C68 VN.n17 VSUBS 0.044426f
C69 VN.n18 VSUBS 0.038765f
C70 VN.n19 VSUBS 0.038765f
C71 VN.n20 VSUBS 0.038765f
C72 VN.n21 VSUBS 0.035093f
C73 VN.n22 VSUBS 0.05812f
C74 VN.n23 VSUBS 0.798007f
C75 VN.n24 VSUBS 0.035698f
C76 VN.n25 VSUBS 0.038765f
C77 VN.t4 VSUBS 2.04088f
C78 VN.n26 VSUBS 0.064401f
C79 VN.n27 VSUBS 0.038765f
C80 VN.t5 VSUBS 2.04088f
C81 VN.n28 VSUBS 0.731415f
C82 VN.t1 VSUBS 2.04088f
C83 VN.n29 VSUBS 0.767994f
C84 VN.n30 VSUBS 0.038765f
C85 VN.t2 VSUBS 2.04088f
C86 VN.n31 VSUBS 0.784152f
C87 VN.t3 VSUBS 2.11804f
C88 VN.n32 VSUBS 0.827632f
C89 VN.n33 VSUBS 0.202833f
C90 VN.n34 VSUBS 0.044426f
C91 VN.n35 VSUBS 0.050653f
C92 VN.n36 VSUBS 0.062535f
C93 VN.n37 VSUBS 0.038765f
C94 VN.n38 VSUBS 0.038765f
C95 VN.n39 VSUBS 0.038765f
C96 VN.n40 VSUBS 0.062535f
C97 VN.n41 VSUBS 0.050653f
C98 VN.n42 VSUBS 0.044426f
C99 VN.n43 VSUBS 0.038765f
C100 VN.n44 VSUBS 0.038765f
C101 VN.n45 VSUBS 0.038765f
C102 VN.n46 VSUBS 0.035093f
C103 VN.n47 VSUBS 0.05812f
C104 VN.n48 VSUBS 0.798007f
C105 VN.n49 VSUBS 2.01818f
C106 VDD1.t5 VSUBS 3.41236f
C107 VDD1.t1 VSUBS 0.322127f
C108 VDD1.t4 VSUBS 0.322127f
C109 VDD1.n0 VSUBS 2.6141f
C110 VDD1.n1 VSUBS 1.40976f
C111 VDD1.t9 VSUBS 3.41235f
C112 VDD1.t2 VSUBS 0.322127f
C113 VDD1.t0 VSUBS 0.322127f
C114 VDD1.n2 VSUBS 2.6141f
C115 VDD1.n3 VSUBS 1.40199f
C116 VDD1.t8 VSUBS 0.322127f
C117 VDD1.t3 VSUBS 0.322127f
C118 VDD1.n4 VSUBS 2.62426f
C119 VDD1.n5 VSUBS 2.9977f
C120 VDD1.t6 VSUBS 0.322127f
C121 VDD1.t7 VSUBS 0.322127f
C122 VDD1.n6 VSUBS 2.61409f
C123 VDD1.n7 VSUBS 3.40082f
C124 VTAIL.t2 VSUBS 0.326703f
C125 VTAIL.t7 VSUBS 0.326703f
C126 VTAIL.n0 VSUBS 2.48999f
C127 VTAIL.n1 VSUBS 0.852128f
C128 VTAIL.t12 VSUBS 3.26328f
C129 VTAIL.n2 VSUBS 0.995481f
C130 VTAIL.t10 VSUBS 0.326703f
C131 VTAIL.t11 VSUBS 0.326703f
C132 VTAIL.n3 VSUBS 2.48999f
C133 VTAIL.n4 VSUBS 0.897652f
C134 VTAIL.t14 VSUBS 0.326703f
C135 VTAIL.t16 VSUBS 0.326703f
C136 VTAIL.n5 VSUBS 2.48999f
C137 VTAIL.n6 VSUBS 2.54339f
C138 VTAIL.t5 VSUBS 0.326703f
C139 VTAIL.t8 VSUBS 0.326703f
C140 VTAIL.n7 VSUBS 2.48999f
C141 VTAIL.n8 VSUBS 2.54338f
C142 VTAIL.t0 VSUBS 0.326703f
C143 VTAIL.t4 VSUBS 0.326703f
C144 VTAIL.n9 VSUBS 2.48999f
C145 VTAIL.n10 VSUBS 0.897646f
C146 VTAIL.t1 VSUBS 3.26328f
C147 VTAIL.n11 VSUBS 0.995476f
C148 VTAIL.t18 VSUBS 0.326703f
C149 VTAIL.t13 VSUBS 0.326703f
C150 VTAIL.n12 VSUBS 2.48999f
C151 VTAIL.n13 VSUBS 0.877754f
C152 VTAIL.t17 VSUBS 0.326703f
C153 VTAIL.t19 VSUBS 0.326703f
C154 VTAIL.n14 VSUBS 2.48999f
C155 VTAIL.n15 VSUBS 0.897646f
C156 VTAIL.t15 VSUBS 3.26328f
C157 VTAIL.n16 VSUBS 2.53793f
C158 VTAIL.t6 VSUBS 3.26328f
C159 VTAIL.n17 VSUBS 2.53793f
C160 VTAIL.t9 VSUBS 0.326703f
C161 VTAIL.t3 VSUBS 0.326703f
C162 VTAIL.n18 VSUBS 2.48999f
C163 VTAIL.n19 VSUBS 0.800102f
C164 VP.n0 VSUBS 0.039502f
C165 VP.t6 VSUBS 2.07966f
C166 VP.n1 VSUBS 0.065625f
C167 VP.n2 VSUBS 0.039502f
C168 VP.t9 VSUBS 2.07966f
C169 VP.n3 VSUBS 0.782587f
C170 VP.n4 VSUBS 0.039502f
C171 VP.t7 VSUBS 2.07966f
C172 VP.n5 VSUBS 0.745313f
C173 VP.n6 VSUBS 0.039502f
C174 VP.t0 VSUBS 2.07966f
C175 VP.n7 VSUBS 0.81317f
C176 VP.n8 VSUBS 0.039502f
C177 VP.t2 VSUBS 2.07966f
C178 VP.n9 VSUBS 0.065625f
C179 VP.n10 VSUBS 0.039502f
C180 VP.t5 VSUBS 2.07966f
C181 VP.n11 VSUBS 0.782587f
C182 VP.n12 VSUBS 0.039502f
C183 VP.t8 VSUBS 2.07966f
C184 VP.n13 VSUBS 0.799052f
C185 VP.t4 VSUBS 2.15829f
C186 VP.n14 VSUBS 0.843358f
C187 VP.n15 VSUBS 0.206687f
C188 VP.n16 VSUBS 0.04527f
C189 VP.n17 VSUBS 0.051615f
C190 VP.n18 VSUBS 0.063723f
C191 VP.n19 VSUBS 0.039502f
C192 VP.n20 VSUBS 0.039502f
C193 VP.n21 VSUBS 0.039502f
C194 VP.n22 VSUBS 0.063723f
C195 VP.n23 VSUBS 0.051615f
C196 VP.t3 VSUBS 2.07966f
C197 VP.n24 VSUBS 0.745313f
C198 VP.n25 VSUBS 0.04527f
C199 VP.n26 VSUBS 0.039502f
C200 VP.n27 VSUBS 0.039502f
C201 VP.n28 VSUBS 0.039502f
C202 VP.n29 VSUBS 0.035759f
C203 VP.n30 VSUBS 0.059224f
C204 VP.n31 VSUBS 0.81317f
C205 VP.n32 VSUBS 2.0308f
C206 VP.n33 VSUBS 2.06032f
C207 VP.n34 VSUBS 0.039502f
C208 VP.n35 VSUBS 0.059224f
C209 VP.n36 VSUBS 0.035759f
C210 VP.n37 VSUBS 0.065625f
C211 VP.n38 VSUBS 0.039502f
C212 VP.n39 VSUBS 0.039502f
C213 VP.n40 VSUBS 0.04527f
C214 VP.n41 VSUBS 0.051615f
C215 VP.n42 VSUBS 0.063723f
C216 VP.n43 VSUBS 0.039502f
C217 VP.n44 VSUBS 0.039502f
C218 VP.n45 VSUBS 0.039502f
C219 VP.n46 VSUBS 0.063723f
C220 VP.n47 VSUBS 0.051615f
C221 VP.t1 VSUBS 2.07966f
C222 VP.n48 VSUBS 0.745313f
C223 VP.n49 VSUBS 0.04527f
C224 VP.n50 VSUBS 0.039502f
C225 VP.n51 VSUBS 0.039502f
C226 VP.n52 VSUBS 0.039502f
C227 VP.n53 VSUBS 0.035759f
C228 VP.n54 VSUBS 0.059224f
C229 VP.n55 VSUBS 0.81317f
C230 VP.n56 VSUBS 0.036376f
C231 B.n0 VSUBS 0.007741f
C232 B.n1 VSUBS 0.007741f
C233 B.n2 VSUBS 0.011448f
C234 B.n3 VSUBS 0.008773f
C235 B.n4 VSUBS 0.008773f
C236 B.n5 VSUBS 0.008773f
C237 B.n6 VSUBS 0.008773f
C238 B.n7 VSUBS 0.008773f
C239 B.n8 VSUBS 0.008773f
C240 B.n9 VSUBS 0.008773f
C241 B.n10 VSUBS 0.008773f
C242 B.n11 VSUBS 0.008773f
C243 B.n12 VSUBS 0.008773f
C244 B.n13 VSUBS 0.008773f
C245 B.n14 VSUBS 0.008773f
C246 B.n15 VSUBS 0.008773f
C247 B.n16 VSUBS 0.008773f
C248 B.n17 VSUBS 0.008773f
C249 B.n18 VSUBS 0.008773f
C250 B.n19 VSUBS 0.008773f
C251 B.n20 VSUBS 0.021942f
C252 B.n21 VSUBS 0.008773f
C253 B.n22 VSUBS 0.008773f
C254 B.n23 VSUBS 0.008773f
C255 B.n24 VSUBS 0.008773f
C256 B.n25 VSUBS 0.008773f
C257 B.n26 VSUBS 0.008773f
C258 B.n27 VSUBS 0.008773f
C259 B.n28 VSUBS 0.008773f
C260 B.n29 VSUBS 0.008773f
C261 B.n30 VSUBS 0.008773f
C262 B.n31 VSUBS 0.008773f
C263 B.n32 VSUBS 0.008773f
C264 B.n33 VSUBS 0.008773f
C265 B.n34 VSUBS 0.008773f
C266 B.n35 VSUBS 0.008773f
C267 B.n36 VSUBS 0.008773f
C268 B.n37 VSUBS 0.008773f
C269 B.n38 VSUBS 0.008773f
C270 B.n39 VSUBS 0.008773f
C271 B.n40 VSUBS 0.008773f
C272 B.n41 VSUBS 0.008773f
C273 B.n42 VSUBS 0.008773f
C274 B.n43 VSUBS 0.008773f
C275 B.n44 VSUBS 0.008773f
C276 B.n45 VSUBS 0.008773f
C277 B.t10 VSUBS 0.626218f
C278 B.t11 VSUBS 0.642169f
C279 B.t9 VSUBS 1.02406f
C280 B.n46 VSUBS 0.263527f
C281 B.n47 VSUBS 0.083385f
C282 B.n48 VSUBS 0.008773f
C283 B.n49 VSUBS 0.008773f
C284 B.n50 VSUBS 0.008773f
C285 B.n51 VSUBS 0.008773f
C286 B.t4 VSUBS 0.6262f
C287 B.t5 VSUBS 0.642153f
C288 B.t3 VSUBS 1.02406f
C289 B.n52 VSUBS 0.263543f
C290 B.n53 VSUBS 0.083403f
C291 B.n54 VSUBS 0.020325f
C292 B.n55 VSUBS 0.008773f
C293 B.n56 VSUBS 0.008773f
C294 B.n57 VSUBS 0.008773f
C295 B.n58 VSUBS 0.008773f
C296 B.n59 VSUBS 0.008773f
C297 B.n60 VSUBS 0.008773f
C298 B.n61 VSUBS 0.008773f
C299 B.n62 VSUBS 0.008773f
C300 B.n63 VSUBS 0.008773f
C301 B.n64 VSUBS 0.008773f
C302 B.n65 VSUBS 0.008773f
C303 B.n66 VSUBS 0.008773f
C304 B.n67 VSUBS 0.008773f
C305 B.n68 VSUBS 0.008773f
C306 B.n69 VSUBS 0.008773f
C307 B.n70 VSUBS 0.008773f
C308 B.n71 VSUBS 0.008773f
C309 B.n72 VSUBS 0.008773f
C310 B.n73 VSUBS 0.008773f
C311 B.n74 VSUBS 0.008773f
C312 B.n75 VSUBS 0.008773f
C313 B.n76 VSUBS 0.008773f
C314 B.n77 VSUBS 0.008773f
C315 B.n78 VSUBS 0.008773f
C316 B.n79 VSUBS 0.021942f
C317 B.n80 VSUBS 0.008773f
C318 B.n81 VSUBS 0.008773f
C319 B.n82 VSUBS 0.008773f
C320 B.n83 VSUBS 0.008773f
C321 B.n84 VSUBS 0.008773f
C322 B.n85 VSUBS 0.008773f
C323 B.n86 VSUBS 0.008773f
C324 B.n87 VSUBS 0.008773f
C325 B.n88 VSUBS 0.008773f
C326 B.n89 VSUBS 0.008773f
C327 B.n90 VSUBS 0.008773f
C328 B.n91 VSUBS 0.008773f
C329 B.n92 VSUBS 0.008773f
C330 B.n93 VSUBS 0.008773f
C331 B.n94 VSUBS 0.008773f
C332 B.n95 VSUBS 0.008773f
C333 B.n96 VSUBS 0.008773f
C334 B.n97 VSUBS 0.008773f
C335 B.n98 VSUBS 0.008773f
C336 B.n99 VSUBS 0.008773f
C337 B.n100 VSUBS 0.008773f
C338 B.n101 VSUBS 0.008773f
C339 B.n102 VSUBS 0.008773f
C340 B.n103 VSUBS 0.008773f
C341 B.n104 VSUBS 0.008773f
C342 B.n105 VSUBS 0.008773f
C343 B.n106 VSUBS 0.008773f
C344 B.n107 VSUBS 0.008773f
C345 B.n108 VSUBS 0.008773f
C346 B.n109 VSUBS 0.008773f
C347 B.n110 VSUBS 0.008773f
C348 B.n111 VSUBS 0.008773f
C349 B.n112 VSUBS 0.008773f
C350 B.n113 VSUBS 0.008773f
C351 B.n114 VSUBS 0.008773f
C352 B.n115 VSUBS 0.008773f
C353 B.n116 VSUBS 0.022361f
C354 B.n117 VSUBS 0.008773f
C355 B.n118 VSUBS 0.008773f
C356 B.n119 VSUBS 0.008773f
C357 B.n120 VSUBS 0.008773f
C358 B.n121 VSUBS 0.008773f
C359 B.n122 VSUBS 0.008773f
C360 B.n123 VSUBS 0.008773f
C361 B.n124 VSUBS 0.008773f
C362 B.n125 VSUBS 0.008773f
C363 B.n126 VSUBS 0.008773f
C364 B.n127 VSUBS 0.008773f
C365 B.n128 VSUBS 0.008773f
C366 B.n129 VSUBS 0.008773f
C367 B.n130 VSUBS 0.008773f
C368 B.n131 VSUBS 0.008773f
C369 B.n132 VSUBS 0.008773f
C370 B.n133 VSUBS 0.008773f
C371 B.n134 VSUBS 0.008773f
C372 B.n135 VSUBS 0.008773f
C373 B.n136 VSUBS 0.008773f
C374 B.n137 VSUBS 0.008773f
C375 B.n138 VSUBS 0.008773f
C376 B.n139 VSUBS 0.008773f
C377 B.n140 VSUBS 0.008773f
C378 B.n141 VSUBS 0.008773f
C379 B.t8 VSUBS 0.6262f
C380 B.t7 VSUBS 0.642153f
C381 B.t6 VSUBS 1.02406f
C382 B.n142 VSUBS 0.263543f
C383 B.n143 VSUBS 0.083403f
C384 B.n144 VSUBS 0.008773f
C385 B.n145 VSUBS 0.008773f
C386 B.n146 VSUBS 0.008773f
C387 B.n147 VSUBS 0.008773f
C388 B.n148 VSUBS 0.004902f
C389 B.n149 VSUBS 0.008773f
C390 B.n150 VSUBS 0.008773f
C391 B.n151 VSUBS 0.008773f
C392 B.n152 VSUBS 0.008773f
C393 B.n153 VSUBS 0.008773f
C394 B.n154 VSUBS 0.008773f
C395 B.n155 VSUBS 0.008773f
C396 B.n156 VSUBS 0.008773f
C397 B.n157 VSUBS 0.008773f
C398 B.n158 VSUBS 0.008773f
C399 B.n159 VSUBS 0.008773f
C400 B.n160 VSUBS 0.008773f
C401 B.n161 VSUBS 0.008773f
C402 B.n162 VSUBS 0.008773f
C403 B.n163 VSUBS 0.008773f
C404 B.n164 VSUBS 0.008773f
C405 B.n165 VSUBS 0.008773f
C406 B.n166 VSUBS 0.008773f
C407 B.n167 VSUBS 0.008773f
C408 B.n168 VSUBS 0.008773f
C409 B.n169 VSUBS 0.008773f
C410 B.n170 VSUBS 0.008773f
C411 B.n171 VSUBS 0.008773f
C412 B.n172 VSUBS 0.008773f
C413 B.n173 VSUBS 0.021942f
C414 B.n174 VSUBS 0.008773f
C415 B.n175 VSUBS 0.008773f
C416 B.n176 VSUBS 0.008773f
C417 B.n177 VSUBS 0.008773f
C418 B.n178 VSUBS 0.008773f
C419 B.n179 VSUBS 0.008773f
C420 B.n180 VSUBS 0.008773f
C421 B.n181 VSUBS 0.008773f
C422 B.n182 VSUBS 0.008773f
C423 B.n183 VSUBS 0.008773f
C424 B.n184 VSUBS 0.008773f
C425 B.n185 VSUBS 0.008773f
C426 B.n186 VSUBS 0.008773f
C427 B.n187 VSUBS 0.008773f
C428 B.n188 VSUBS 0.008773f
C429 B.n189 VSUBS 0.008773f
C430 B.n190 VSUBS 0.008773f
C431 B.n191 VSUBS 0.008773f
C432 B.n192 VSUBS 0.008773f
C433 B.n193 VSUBS 0.008773f
C434 B.n194 VSUBS 0.008773f
C435 B.n195 VSUBS 0.008773f
C436 B.n196 VSUBS 0.008773f
C437 B.n197 VSUBS 0.008773f
C438 B.n198 VSUBS 0.008773f
C439 B.n199 VSUBS 0.008773f
C440 B.n200 VSUBS 0.008773f
C441 B.n201 VSUBS 0.008773f
C442 B.n202 VSUBS 0.008773f
C443 B.n203 VSUBS 0.008773f
C444 B.n204 VSUBS 0.008773f
C445 B.n205 VSUBS 0.008773f
C446 B.n206 VSUBS 0.008773f
C447 B.n207 VSUBS 0.008773f
C448 B.n208 VSUBS 0.008773f
C449 B.n209 VSUBS 0.008773f
C450 B.n210 VSUBS 0.008773f
C451 B.n211 VSUBS 0.008773f
C452 B.n212 VSUBS 0.008773f
C453 B.n213 VSUBS 0.008773f
C454 B.n214 VSUBS 0.008773f
C455 B.n215 VSUBS 0.008773f
C456 B.n216 VSUBS 0.008773f
C457 B.n217 VSUBS 0.008773f
C458 B.n218 VSUBS 0.008773f
C459 B.n219 VSUBS 0.008773f
C460 B.n220 VSUBS 0.008773f
C461 B.n221 VSUBS 0.008773f
C462 B.n222 VSUBS 0.008773f
C463 B.n223 VSUBS 0.008773f
C464 B.n224 VSUBS 0.008773f
C465 B.n225 VSUBS 0.008773f
C466 B.n226 VSUBS 0.008773f
C467 B.n227 VSUBS 0.008773f
C468 B.n228 VSUBS 0.008773f
C469 B.n229 VSUBS 0.008773f
C470 B.n230 VSUBS 0.008773f
C471 B.n231 VSUBS 0.008773f
C472 B.n232 VSUBS 0.008773f
C473 B.n233 VSUBS 0.008773f
C474 B.n234 VSUBS 0.008773f
C475 B.n235 VSUBS 0.008773f
C476 B.n236 VSUBS 0.008773f
C477 B.n237 VSUBS 0.008773f
C478 B.n238 VSUBS 0.008773f
C479 B.n239 VSUBS 0.008773f
C480 B.n240 VSUBS 0.008773f
C481 B.n241 VSUBS 0.008773f
C482 B.n242 VSUBS 0.021406f
C483 B.n243 VSUBS 0.021406f
C484 B.n244 VSUBS 0.021942f
C485 B.n245 VSUBS 0.008773f
C486 B.n246 VSUBS 0.008773f
C487 B.n247 VSUBS 0.008773f
C488 B.n248 VSUBS 0.008773f
C489 B.n249 VSUBS 0.008773f
C490 B.n250 VSUBS 0.008773f
C491 B.n251 VSUBS 0.008773f
C492 B.n252 VSUBS 0.008773f
C493 B.n253 VSUBS 0.008773f
C494 B.n254 VSUBS 0.008773f
C495 B.n255 VSUBS 0.008773f
C496 B.n256 VSUBS 0.008773f
C497 B.n257 VSUBS 0.008773f
C498 B.n258 VSUBS 0.008773f
C499 B.n259 VSUBS 0.008773f
C500 B.n260 VSUBS 0.008773f
C501 B.n261 VSUBS 0.008773f
C502 B.n262 VSUBS 0.008773f
C503 B.n263 VSUBS 0.008773f
C504 B.n264 VSUBS 0.008773f
C505 B.n265 VSUBS 0.008773f
C506 B.n266 VSUBS 0.008773f
C507 B.n267 VSUBS 0.008773f
C508 B.n268 VSUBS 0.008773f
C509 B.n269 VSUBS 0.008773f
C510 B.n270 VSUBS 0.008773f
C511 B.n271 VSUBS 0.008773f
C512 B.n272 VSUBS 0.008773f
C513 B.n273 VSUBS 0.008773f
C514 B.n274 VSUBS 0.008773f
C515 B.n275 VSUBS 0.008773f
C516 B.n276 VSUBS 0.008773f
C517 B.n277 VSUBS 0.008773f
C518 B.n278 VSUBS 0.008773f
C519 B.n279 VSUBS 0.008773f
C520 B.n280 VSUBS 0.008773f
C521 B.n281 VSUBS 0.008773f
C522 B.n282 VSUBS 0.008773f
C523 B.n283 VSUBS 0.008773f
C524 B.n284 VSUBS 0.008773f
C525 B.n285 VSUBS 0.008773f
C526 B.n286 VSUBS 0.008773f
C527 B.n287 VSUBS 0.008773f
C528 B.n288 VSUBS 0.008773f
C529 B.n289 VSUBS 0.008773f
C530 B.n290 VSUBS 0.008773f
C531 B.n291 VSUBS 0.008773f
C532 B.n292 VSUBS 0.008773f
C533 B.n293 VSUBS 0.008773f
C534 B.n294 VSUBS 0.008773f
C535 B.n295 VSUBS 0.008773f
C536 B.n296 VSUBS 0.008773f
C537 B.n297 VSUBS 0.008773f
C538 B.n298 VSUBS 0.008773f
C539 B.n299 VSUBS 0.008773f
C540 B.n300 VSUBS 0.008773f
C541 B.n301 VSUBS 0.008773f
C542 B.n302 VSUBS 0.008773f
C543 B.n303 VSUBS 0.008773f
C544 B.n304 VSUBS 0.008773f
C545 B.n305 VSUBS 0.008773f
C546 B.n306 VSUBS 0.008773f
C547 B.n307 VSUBS 0.008773f
C548 B.n308 VSUBS 0.008773f
C549 B.n309 VSUBS 0.008773f
C550 B.n310 VSUBS 0.008773f
C551 B.n311 VSUBS 0.008773f
C552 B.n312 VSUBS 0.008773f
C553 B.n313 VSUBS 0.008773f
C554 B.n314 VSUBS 0.008773f
C555 B.n315 VSUBS 0.008773f
C556 B.n316 VSUBS 0.008773f
C557 B.t2 VSUBS 0.626218f
C558 B.t1 VSUBS 0.642169f
C559 B.t0 VSUBS 1.02406f
C560 B.n317 VSUBS 0.263527f
C561 B.n318 VSUBS 0.083385f
C562 B.n319 VSUBS 0.020325f
C563 B.n320 VSUBS 0.008257f
C564 B.n321 VSUBS 0.008773f
C565 B.n322 VSUBS 0.008773f
C566 B.n323 VSUBS 0.008773f
C567 B.n324 VSUBS 0.008773f
C568 B.n325 VSUBS 0.008773f
C569 B.n326 VSUBS 0.008773f
C570 B.n327 VSUBS 0.008773f
C571 B.n328 VSUBS 0.008773f
C572 B.n329 VSUBS 0.008773f
C573 B.n330 VSUBS 0.008773f
C574 B.n331 VSUBS 0.008773f
C575 B.n332 VSUBS 0.008773f
C576 B.n333 VSUBS 0.008773f
C577 B.n334 VSUBS 0.008773f
C578 B.n335 VSUBS 0.008773f
C579 B.n336 VSUBS 0.004902f
C580 B.n337 VSUBS 0.020325f
C581 B.n338 VSUBS 0.008257f
C582 B.n339 VSUBS 0.008773f
C583 B.n340 VSUBS 0.008773f
C584 B.n341 VSUBS 0.008773f
C585 B.n342 VSUBS 0.008773f
C586 B.n343 VSUBS 0.008773f
C587 B.n344 VSUBS 0.008773f
C588 B.n345 VSUBS 0.008773f
C589 B.n346 VSUBS 0.008773f
C590 B.n347 VSUBS 0.008773f
C591 B.n348 VSUBS 0.008773f
C592 B.n349 VSUBS 0.008773f
C593 B.n350 VSUBS 0.008773f
C594 B.n351 VSUBS 0.008773f
C595 B.n352 VSUBS 0.008773f
C596 B.n353 VSUBS 0.008773f
C597 B.n354 VSUBS 0.008773f
C598 B.n355 VSUBS 0.008773f
C599 B.n356 VSUBS 0.008773f
C600 B.n357 VSUBS 0.008773f
C601 B.n358 VSUBS 0.008773f
C602 B.n359 VSUBS 0.008773f
C603 B.n360 VSUBS 0.008773f
C604 B.n361 VSUBS 0.008773f
C605 B.n362 VSUBS 0.008773f
C606 B.n363 VSUBS 0.008773f
C607 B.n364 VSUBS 0.008773f
C608 B.n365 VSUBS 0.008773f
C609 B.n366 VSUBS 0.008773f
C610 B.n367 VSUBS 0.008773f
C611 B.n368 VSUBS 0.008773f
C612 B.n369 VSUBS 0.008773f
C613 B.n370 VSUBS 0.008773f
C614 B.n371 VSUBS 0.008773f
C615 B.n372 VSUBS 0.008773f
C616 B.n373 VSUBS 0.008773f
C617 B.n374 VSUBS 0.008773f
C618 B.n375 VSUBS 0.008773f
C619 B.n376 VSUBS 0.008773f
C620 B.n377 VSUBS 0.008773f
C621 B.n378 VSUBS 0.008773f
C622 B.n379 VSUBS 0.008773f
C623 B.n380 VSUBS 0.008773f
C624 B.n381 VSUBS 0.008773f
C625 B.n382 VSUBS 0.008773f
C626 B.n383 VSUBS 0.008773f
C627 B.n384 VSUBS 0.008773f
C628 B.n385 VSUBS 0.008773f
C629 B.n386 VSUBS 0.008773f
C630 B.n387 VSUBS 0.008773f
C631 B.n388 VSUBS 0.008773f
C632 B.n389 VSUBS 0.008773f
C633 B.n390 VSUBS 0.008773f
C634 B.n391 VSUBS 0.008773f
C635 B.n392 VSUBS 0.008773f
C636 B.n393 VSUBS 0.008773f
C637 B.n394 VSUBS 0.008773f
C638 B.n395 VSUBS 0.008773f
C639 B.n396 VSUBS 0.008773f
C640 B.n397 VSUBS 0.008773f
C641 B.n398 VSUBS 0.008773f
C642 B.n399 VSUBS 0.008773f
C643 B.n400 VSUBS 0.008773f
C644 B.n401 VSUBS 0.008773f
C645 B.n402 VSUBS 0.008773f
C646 B.n403 VSUBS 0.008773f
C647 B.n404 VSUBS 0.008773f
C648 B.n405 VSUBS 0.008773f
C649 B.n406 VSUBS 0.008773f
C650 B.n407 VSUBS 0.008773f
C651 B.n408 VSUBS 0.008773f
C652 B.n409 VSUBS 0.008773f
C653 B.n410 VSUBS 0.008773f
C654 B.n411 VSUBS 0.020986f
C655 B.n412 VSUBS 0.021942f
C656 B.n413 VSUBS 0.021406f
C657 B.n414 VSUBS 0.008773f
C658 B.n415 VSUBS 0.008773f
C659 B.n416 VSUBS 0.008773f
C660 B.n417 VSUBS 0.008773f
C661 B.n418 VSUBS 0.008773f
C662 B.n419 VSUBS 0.008773f
C663 B.n420 VSUBS 0.008773f
C664 B.n421 VSUBS 0.008773f
C665 B.n422 VSUBS 0.008773f
C666 B.n423 VSUBS 0.008773f
C667 B.n424 VSUBS 0.008773f
C668 B.n425 VSUBS 0.008773f
C669 B.n426 VSUBS 0.008773f
C670 B.n427 VSUBS 0.008773f
C671 B.n428 VSUBS 0.008773f
C672 B.n429 VSUBS 0.008773f
C673 B.n430 VSUBS 0.008773f
C674 B.n431 VSUBS 0.008773f
C675 B.n432 VSUBS 0.008773f
C676 B.n433 VSUBS 0.008773f
C677 B.n434 VSUBS 0.008773f
C678 B.n435 VSUBS 0.008773f
C679 B.n436 VSUBS 0.008773f
C680 B.n437 VSUBS 0.008773f
C681 B.n438 VSUBS 0.008773f
C682 B.n439 VSUBS 0.008773f
C683 B.n440 VSUBS 0.008773f
C684 B.n441 VSUBS 0.008773f
C685 B.n442 VSUBS 0.008773f
C686 B.n443 VSUBS 0.008773f
C687 B.n444 VSUBS 0.008773f
C688 B.n445 VSUBS 0.008773f
C689 B.n446 VSUBS 0.008773f
C690 B.n447 VSUBS 0.008773f
C691 B.n448 VSUBS 0.008773f
C692 B.n449 VSUBS 0.008773f
C693 B.n450 VSUBS 0.008773f
C694 B.n451 VSUBS 0.008773f
C695 B.n452 VSUBS 0.008773f
C696 B.n453 VSUBS 0.008773f
C697 B.n454 VSUBS 0.008773f
C698 B.n455 VSUBS 0.008773f
C699 B.n456 VSUBS 0.008773f
C700 B.n457 VSUBS 0.008773f
C701 B.n458 VSUBS 0.008773f
C702 B.n459 VSUBS 0.008773f
C703 B.n460 VSUBS 0.008773f
C704 B.n461 VSUBS 0.008773f
C705 B.n462 VSUBS 0.008773f
C706 B.n463 VSUBS 0.008773f
C707 B.n464 VSUBS 0.008773f
C708 B.n465 VSUBS 0.008773f
C709 B.n466 VSUBS 0.008773f
C710 B.n467 VSUBS 0.008773f
C711 B.n468 VSUBS 0.008773f
C712 B.n469 VSUBS 0.008773f
C713 B.n470 VSUBS 0.008773f
C714 B.n471 VSUBS 0.008773f
C715 B.n472 VSUBS 0.008773f
C716 B.n473 VSUBS 0.008773f
C717 B.n474 VSUBS 0.008773f
C718 B.n475 VSUBS 0.008773f
C719 B.n476 VSUBS 0.008773f
C720 B.n477 VSUBS 0.008773f
C721 B.n478 VSUBS 0.008773f
C722 B.n479 VSUBS 0.008773f
C723 B.n480 VSUBS 0.008773f
C724 B.n481 VSUBS 0.008773f
C725 B.n482 VSUBS 0.008773f
C726 B.n483 VSUBS 0.008773f
C727 B.n484 VSUBS 0.008773f
C728 B.n485 VSUBS 0.008773f
C729 B.n486 VSUBS 0.008773f
C730 B.n487 VSUBS 0.008773f
C731 B.n488 VSUBS 0.008773f
C732 B.n489 VSUBS 0.008773f
C733 B.n490 VSUBS 0.008773f
C734 B.n491 VSUBS 0.008773f
C735 B.n492 VSUBS 0.008773f
C736 B.n493 VSUBS 0.008773f
C737 B.n494 VSUBS 0.008773f
C738 B.n495 VSUBS 0.008773f
C739 B.n496 VSUBS 0.008773f
C740 B.n497 VSUBS 0.008773f
C741 B.n498 VSUBS 0.008773f
C742 B.n499 VSUBS 0.008773f
C743 B.n500 VSUBS 0.008773f
C744 B.n501 VSUBS 0.008773f
C745 B.n502 VSUBS 0.008773f
C746 B.n503 VSUBS 0.008773f
C747 B.n504 VSUBS 0.008773f
C748 B.n505 VSUBS 0.008773f
C749 B.n506 VSUBS 0.008773f
C750 B.n507 VSUBS 0.008773f
C751 B.n508 VSUBS 0.008773f
C752 B.n509 VSUBS 0.008773f
C753 B.n510 VSUBS 0.008773f
C754 B.n511 VSUBS 0.008773f
C755 B.n512 VSUBS 0.008773f
C756 B.n513 VSUBS 0.008773f
C757 B.n514 VSUBS 0.008773f
C758 B.n515 VSUBS 0.008773f
C759 B.n516 VSUBS 0.008773f
C760 B.n517 VSUBS 0.008773f
C761 B.n518 VSUBS 0.008773f
C762 B.n519 VSUBS 0.008773f
C763 B.n520 VSUBS 0.008773f
C764 B.n521 VSUBS 0.008773f
C765 B.n522 VSUBS 0.021406f
C766 B.n523 VSUBS 0.021406f
C767 B.n524 VSUBS 0.021942f
C768 B.n525 VSUBS 0.008773f
C769 B.n526 VSUBS 0.008773f
C770 B.n527 VSUBS 0.008773f
C771 B.n528 VSUBS 0.008773f
C772 B.n529 VSUBS 0.008773f
C773 B.n530 VSUBS 0.008773f
C774 B.n531 VSUBS 0.008773f
C775 B.n532 VSUBS 0.008773f
C776 B.n533 VSUBS 0.008773f
C777 B.n534 VSUBS 0.008773f
C778 B.n535 VSUBS 0.008773f
C779 B.n536 VSUBS 0.008773f
C780 B.n537 VSUBS 0.008773f
C781 B.n538 VSUBS 0.008773f
C782 B.n539 VSUBS 0.008773f
C783 B.n540 VSUBS 0.008773f
C784 B.n541 VSUBS 0.008773f
C785 B.n542 VSUBS 0.008773f
C786 B.n543 VSUBS 0.008773f
C787 B.n544 VSUBS 0.008773f
C788 B.n545 VSUBS 0.008773f
C789 B.n546 VSUBS 0.008773f
C790 B.n547 VSUBS 0.008773f
C791 B.n548 VSUBS 0.008773f
C792 B.n549 VSUBS 0.008773f
C793 B.n550 VSUBS 0.008773f
C794 B.n551 VSUBS 0.008773f
C795 B.n552 VSUBS 0.008773f
C796 B.n553 VSUBS 0.008773f
C797 B.n554 VSUBS 0.008773f
C798 B.n555 VSUBS 0.008773f
C799 B.n556 VSUBS 0.008773f
C800 B.n557 VSUBS 0.008773f
C801 B.n558 VSUBS 0.008773f
C802 B.n559 VSUBS 0.008773f
C803 B.n560 VSUBS 0.008773f
C804 B.n561 VSUBS 0.008773f
C805 B.n562 VSUBS 0.008773f
C806 B.n563 VSUBS 0.008773f
C807 B.n564 VSUBS 0.008773f
C808 B.n565 VSUBS 0.008773f
C809 B.n566 VSUBS 0.008773f
C810 B.n567 VSUBS 0.008773f
C811 B.n568 VSUBS 0.008773f
C812 B.n569 VSUBS 0.008773f
C813 B.n570 VSUBS 0.008773f
C814 B.n571 VSUBS 0.008773f
C815 B.n572 VSUBS 0.008773f
C816 B.n573 VSUBS 0.008773f
C817 B.n574 VSUBS 0.008773f
C818 B.n575 VSUBS 0.008773f
C819 B.n576 VSUBS 0.008773f
C820 B.n577 VSUBS 0.008773f
C821 B.n578 VSUBS 0.008773f
C822 B.n579 VSUBS 0.008773f
C823 B.n580 VSUBS 0.008773f
C824 B.n581 VSUBS 0.008773f
C825 B.n582 VSUBS 0.008773f
C826 B.n583 VSUBS 0.008773f
C827 B.n584 VSUBS 0.008773f
C828 B.n585 VSUBS 0.008773f
C829 B.n586 VSUBS 0.008773f
C830 B.n587 VSUBS 0.008773f
C831 B.n588 VSUBS 0.008773f
C832 B.n589 VSUBS 0.008773f
C833 B.n590 VSUBS 0.008773f
C834 B.n591 VSUBS 0.008773f
C835 B.n592 VSUBS 0.008773f
C836 B.n593 VSUBS 0.008773f
C837 B.n594 VSUBS 0.008773f
C838 B.n595 VSUBS 0.008773f
C839 B.n596 VSUBS 0.008773f
C840 B.n597 VSUBS 0.008257f
C841 B.n598 VSUBS 0.008773f
C842 B.n599 VSUBS 0.008773f
C843 B.n600 VSUBS 0.004902f
C844 B.n601 VSUBS 0.008773f
C845 B.n602 VSUBS 0.008773f
C846 B.n603 VSUBS 0.008773f
C847 B.n604 VSUBS 0.008773f
C848 B.n605 VSUBS 0.008773f
C849 B.n606 VSUBS 0.008773f
C850 B.n607 VSUBS 0.008773f
C851 B.n608 VSUBS 0.008773f
C852 B.n609 VSUBS 0.008773f
C853 B.n610 VSUBS 0.008773f
C854 B.n611 VSUBS 0.008773f
C855 B.n612 VSUBS 0.008773f
C856 B.n613 VSUBS 0.004902f
C857 B.n614 VSUBS 0.020325f
C858 B.n615 VSUBS 0.008257f
C859 B.n616 VSUBS 0.008773f
C860 B.n617 VSUBS 0.008773f
C861 B.n618 VSUBS 0.008773f
C862 B.n619 VSUBS 0.008773f
C863 B.n620 VSUBS 0.008773f
C864 B.n621 VSUBS 0.008773f
C865 B.n622 VSUBS 0.008773f
C866 B.n623 VSUBS 0.008773f
C867 B.n624 VSUBS 0.008773f
C868 B.n625 VSUBS 0.008773f
C869 B.n626 VSUBS 0.008773f
C870 B.n627 VSUBS 0.008773f
C871 B.n628 VSUBS 0.008773f
C872 B.n629 VSUBS 0.008773f
C873 B.n630 VSUBS 0.008773f
C874 B.n631 VSUBS 0.008773f
C875 B.n632 VSUBS 0.008773f
C876 B.n633 VSUBS 0.008773f
C877 B.n634 VSUBS 0.008773f
C878 B.n635 VSUBS 0.008773f
C879 B.n636 VSUBS 0.008773f
C880 B.n637 VSUBS 0.008773f
C881 B.n638 VSUBS 0.008773f
C882 B.n639 VSUBS 0.008773f
C883 B.n640 VSUBS 0.008773f
C884 B.n641 VSUBS 0.008773f
C885 B.n642 VSUBS 0.008773f
C886 B.n643 VSUBS 0.008773f
C887 B.n644 VSUBS 0.008773f
C888 B.n645 VSUBS 0.008773f
C889 B.n646 VSUBS 0.008773f
C890 B.n647 VSUBS 0.008773f
C891 B.n648 VSUBS 0.008773f
C892 B.n649 VSUBS 0.008773f
C893 B.n650 VSUBS 0.008773f
C894 B.n651 VSUBS 0.008773f
C895 B.n652 VSUBS 0.008773f
C896 B.n653 VSUBS 0.008773f
C897 B.n654 VSUBS 0.008773f
C898 B.n655 VSUBS 0.008773f
C899 B.n656 VSUBS 0.008773f
C900 B.n657 VSUBS 0.008773f
C901 B.n658 VSUBS 0.008773f
C902 B.n659 VSUBS 0.008773f
C903 B.n660 VSUBS 0.008773f
C904 B.n661 VSUBS 0.008773f
C905 B.n662 VSUBS 0.008773f
C906 B.n663 VSUBS 0.008773f
C907 B.n664 VSUBS 0.008773f
C908 B.n665 VSUBS 0.008773f
C909 B.n666 VSUBS 0.008773f
C910 B.n667 VSUBS 0.008773f
C911 B.n668 VSUBS 0.008773f
C912 B.n669 VSUBS 0.008773f
C913 B.n670 VSUBS 0.008773f
C914 B.n671 VSUBS 0.008773f
C915 B.n672 VSUBS 0.008773f
C916 B.n673 VSUBS 0.008773f
C917 B.n674 VSUBS 0.008773f
C918 B.n675 VSUBS 0.008773f
C919 B.n676 VSUBS 0.008773f
C920 B.n677 VSUBS 0.008773f
C921 B.n678 VSUBS 0.008773f
C922 B.n679 VSUBS 0.008773f
C923 B.n680 VSUBS 0.008773f
C924 B.n681 VSUBS 0.008773f
C925 B.n682 VSUBS 0.008773f
C926 B.n683 VSUBS 0.008773f
C927 B.n684 VSUBS 0.008773f
C928 B.n685 VSUBS 0.008773f
C929 B.n686 VSUBS 0.008773f
C930 B.n687 VSUBS 0.008773f
C931 B.n688 VSUBS 0.008773f
C932 B.n689 VSUBS 0.021942f
C933 B.n690 VSUBS 0.021406f
C934 B.n691 VSUBS 0.021406f
C935 B.n692 VSUBS 0.008773f
C936 B.n693 VSUBS 0.008773f
C937 B.n694 VSUBS 0.008773f
C938 B.n695 VSUBS 0.008773f
C939 B.n696 VSUBS 0.008773f
C940 B.n697 VSUBS 0.008773f
C941 B.n698 VSUBS 0.008773f
C942 B.n699 VSUBS 0.008773f
C943 B.n700 VSUBS 0.008773f
C944 B.n701 VSUBS 0.008773f
C945 B.n702 VSUBS 0.008773f
C946 B.n703 VSUBS 0.008773f
C947 B.n704 VSUBS 0.008773f
C948 B.n705 VSUBS 0.008773f
C949 B.n706 VSUBS 0.008773f
C950 B.n707 VSUBS 0.008773f
C951 B.n708 VSUBS 0.008773f
C952 B.n709 VSUBS 0.008773f
C953 B.n710 VSUBS 0.008773f
C954 B.n711 VSUBS 0.008773f
C955 B.n712 VSUBS 0.008773f
C956 B.n713 VSUBS 0.008773f
C957 B.n714 VSUBS 0.008773f
C958 B.n715 VSUBS 0.008773f
C959 B.n716 VSUBS 0.008773f
C960 B.n717 VSUBS 0.008773f
C961 B.n718 VSUBS 0.008773f
C962 B.n719 VSUBS 0.008773f
C963 B.n720 VSUBS 0.008773f
C964 B.n721 VSUBS 0.008773f
C965 B.n722 VSUBS 0.008773f
C966 B.n723 VSUBS 0.008773f
C967 B.n724 VSUBS 0.008773f
C968 B.n725 VSUBS 0.008773f
C969 B.n726 VSUBS 0.008773f
C970 B.n727 VSUBS 0.008773f
C971 B.n728 VSUBS 0.008773f
C972 B.n729 VSUBS 0.008773f
C973 B.n730 VSUBS 0.008773f
C974 B.n731 VSUBS 0.008773f
C975 B.n732 VSUBS 0.008773f
C976 B.n733 VSUBS 0.008773f
C977 B.n734 VSUBS 0.008773f
C978 B.n735 VSUBS 0.008773f
C979 B.n736 VSUBS 0.008773f
C980 B.n737 VSUBS 0.008773f
C981 B.n738 VSUBS 0.008773f
C982 B.n739 VSUBS 0.008773f
C983 B.n740 VSUBS 0.008773f
C984 B.n741 VSUBS 0.008773f
C985 B.n742 VSUBS 0.008773f
C986 B.n743 VSUBS 0.011448f
C987 B.n744 VSUBS 0.012195f
C988 B.n745 VSUBS 0.024251f
.ends

