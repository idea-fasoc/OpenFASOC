* NGSPICE file created from diff_pair_sample_1605.ext - technology: sky130A

.subckt diff_pair_sample_1605 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=2
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=2
X2 VDD1.t5 VP.t0 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=2
X3 VDD1.t4 VP.t1 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=2
X4 VTAIL.t6 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=2
X5 VDD1.t3 VP.t2 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=2
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=2
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=2
X8 VDD2.t3 VN.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=2
X9 VDD2.t2 VN.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=2
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=0 ps=0 w=7.25 l=2
X11 VTAIL.t9 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=2
X12 VDD1.t2 VP.t3 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8275 pd=15.28 as=1.19625 ps=7.58 w=7.25 l=2
X13 VTAIL.t2 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=2
X14 VTAIL.t5 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=1.19625 ps=7.58 w=7.25 l=2
X15 VDD2.t0 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.19625 pd=7.58 as=2.8275 ps=15.28 w=7.25 l=2
R0 B.n619 B.n618 585
R1 B.n620 B.n619 585
R2 B.n230 B.n100 585
R3 B.n229 B.n228 585
R4 B.n227 B.n226 585
R5 B.n225 B.n224 585
R6 B.n223 B.n222 585
R7 B.n221 B.n220 585
R8 B.n219 B.n218 585
R9 B.n217 B.n216 585
R10 B.n215 B.n214 585
R11 B.n213 B.n212 585
R12 B.n211 B.n210 585
R13 B.n209 B.n208 585
R14 B.n207 B.n206 585
R15 B.n205 B.n204 585
R16 B.n203 B.n202 585
R17 B.n201 B.n200 585
R18 B.n199 B.n198 585
R19 B.n197 B.n196 585
R20 B.n195 B.n194 585
R21 B.n193 B.n192 585
R22 B.n191 B.n190 585
R23 B.n189 B.n188 585
R24 B.n187 B.n186 585
R25 B.n185 B.n184 585
R26 B.n183 B.n182 585
R27 B.n181 B.n180 585
R28 B.n179 B.n178 585
R29 B.n176 B.n175 585
R30 B.n174 B.n173 585
R31 B.n172 B.n171 585
R32 B.n170 B.n169 585
R33 B.n168 B.n167 585
R34 B.n166 B.n165 585
R35 B.n164 B.n163 585
R36 B.n162 B.n161 585
R37 B.n160 B.n159 585
R38 B.n158 B.n157 585
R39 B.n156 B.n155 585
R40 B.n154 B.n153 585
R41 B.n152 B.n151 585
R42 B.n150 B.n149 585
R43 B.n148 B.n147 585
R44 B.n146 B.n145 585
R45 B.n144 B.n143 585
R46 B.n142 B.n141 585
R47 B.n140 B.n139 585
R48 B.n138 B.n137 585
R49 B.n136 B.n135 585
R50 B.n134 B.n133 585
R51 B.n132 B.n131 585
R52 B.n130 B.n129 585
R53 B.n128 B.n127 585
R54 B.n126 B.n125 585
R55 B.n124 B.n123 585
R56 B.n122 B.n121 585
R57 B.n120 B.n119 585
R58 B.n118 B.n117 585
R59 B.n116 B.n115 585
R60 B.n114 B.n113 585
R61 B.n112 B.n111 585
R62 B.n110 B.n109 585
R63 B.n108 B.n107 585
R64 B.n68 B.n67 585
R65 B.n623 B.n622 585
R66 B.n617 B.n101 585
R67 B.n101 B.n65 585
R68 B.n616 B.n64 585
R69 B.n627 B.n64 585
R70 B.n615 B.n63 585
R71 B.n628 B.n63 585
R72 B.n614 B.n62 585
R73 B.n629 B.n62 585
R74 B.n613 B.n612 585
R75 B.n612 B.n58 585
R76 B.n611 B.n57 585
R77 B.n635 B.n57 585
R78 B.n610 B.n56 585
R79 B.n636 B.n56 585
R80 B.n609 B.n55 585
R81 B.n637 B.n55 585
R82 B.n608 B.n607 585
R83 B.n607 B.n51 585
R84 B.n606 B.n50 585
R85 B.n643 B.n50 585
R86 B.n605 B.n49 585
R87 B.n644 B.n49 585
R88 B.n604 B.n48 585
R89 B.n645 B.n48 585
R90 B.n603 B.n602 585
R91 B.n602 B.n44 585
R92 B.n601 B.n43 585
R93 B.n651 B.n43 585
R94 B.n600 B.n42 585
R95 B.n652 B.n42 585
R96 B.n599 B.n41 585
R97 B.n653 B.n41 585
R98 B.n598 B.n597 585
R99 B.n597 B.n40 585
R100 B.n596 B.n36 585
R101 B.n659 B.n36 585
R102 B.n595 B.n35 585
R103 B.n660 B.n35 585
R104 B.n594 B.n34 585
R105 B.n661 B.n34 585
R106 B.n593 B.n592 585
R107 B.n592 B.n30 585
R108 B.n591 B.n29 585
R109 B.n667 B.n29 585
R110 B.n590 B.n28 585
R111 B.n668 B.n28 585
R112 B.n589 B.n27 585
R113 B.n669 B.n27 585
R114 B.n588 B.n587 585
R115 B.n587 B.n23 585
R116 B.n586 B.n22 585
R117 B.n675 B.n22 585
R118 B.n585 B.n21 585
R119 B.n676 B.n21 585
R120 B.n584 B.n20 585
R121 B.n677 B.n20 585
R122 B.n583 B.n582 585
R123 B.n582 B.n16 585
R124 B.n581 B.n15 585
R125 B.n683 B.n15 585
R126 B.n580 B.n14 585
R127 B.n684 B.n14 585
R128 B.n579 B.n13 585
R129 B.n685 B.n13 585
R130 B.n578 B.n577 585
R131 B.n577 B.n12 585
R132 B.n576 B.n575 585
R133 B.n576 B.n8 585
R134 B.n574 B.n7 585
R135 B.n692 B.n7 585
R136 B.n573 B.n6 585
R137 B.n693 B.n6 585
R138 B.n572 B.n5 585
R139 B.n694 B.n5 585
R140 B.n571 B.n570 585
R141 B.n570 B.n4 585
R142 B.n569 B.n231 585
R143 B.n569 B.n568 585
R144 B.n559 B.n232 585
R145 B.n233 B.n232 585
R146 B.n561 B.n560 585
R147 B.n562 B.n561 585
R148 B.n558 B.n237 585
R149 B.n241 B.n237 585
R150 B.n557 B.n556 585
R151 B.n556 B.n555 585
R152 B.n239 B.n238 585
R153 B.n240 B.n239 585
R154 B.n548 B.n547 585
R155 B.n549 B.n548 585
R156 B.n546 B.n246 585
R157 B.n246 B.n245 585
R158 B.n545 B.n544 585
R159 B.n544 B.n543 585
R160 B.n248 B.n247 585
R161 B.n249 B.n248 585
R162 B.n536 B.n535 585
R163 B.n537 B.n536 585
R164 B.n534 B.n254 585
R165 B.n254 B.n253 585
R166 B.n533 B.n532 585
R167 B.n532 B.n531 585
R168 B.n256 B.n255 585
R169 B.n257 B.n256 585
R170 B.n524 B.n523 585
R171 B.n525 B.n524 585
R172 B.n522 B.n262 585
R173 B.n262 B.n261 585
R174 B.n521 B.n520 585
R175 B.n520 B.n519 585
R176 B.n264 B.n263 585
R177 B.n512 B.n264 585
R178 B.n511 B.n510 585
R179 B.n513 B.n511 585
R180 B.n509 B.n269 585
R181 B.n269 B.n268 585
R182 B.n508 B.n507 585
R183 B.n507 B.n506 585
R184 B.n271 B.n270 585
R185 B.n272 B.n271 585
R186 B.n499 B.n498 585
R187 B.n500 B.n499 585
R188 B.n497 B.n277 585
R189 B.n277 B.n276 585
R190 B.n496 B.n495 585
R191 B.n495 B.n494 585
R192 B.n279 B.n278 585
R193 B.n280 B.n279 585
R194 B.n487 B.n486 585
R195 B.n488 B.n487 585
R196 B.n485 B.n284 585
R197 B.n288 B.n284 585
R198 B.n484 B.n483 585
R199 B.n483 B.n482 585
R200 B.n286 B.n285 585
R201 B.n287 B.n286 585
R202 B.n475 B.n474 585
R203 B.n476 B.n475 585
R204 B.n473 B.n293 585
R205 B.n293 B.n292 585
R206 B.n472 B.n471 585
R207 B.n471 B.n470 585
R208 B.n295 B.n294 585
R209 B.n296 B.n295 585
R210 B.n466 B.n465 585
R211 B.n299 B.n298 585
R212 B.n462 B.n461 585
R213 B.n463 B.n462 585
R214 B.n460 B.n331 585
R215 B.n459 B.n458 585
R216 B.n457 B.n456 585
R217 B.n455 B.n454 585
R218 B.n453 B.n452 585
R219 B.n451 B.n450 585
R220 B.n449 B.n448 585
R221 B.n447 B.n446 585
R222 B.n445 B.n444 585
R223 B.n443 B.n442 585
R224 B.n441 B.n440 585
R225 B.n439 B.n438 585
R226 B.n437 B.n436 585
R227 B.n435 B.n434 585
R228 B.n433 B.n432 585
R229 B.n431 B.n430 585
R230 B.n429 B.n428 585
R231 B.n427 B.n426 585
R232 B.n425 B.n424 585
R233 B.n423 B.n422 585
R234 B.n421 B.n420 585
R235 B.n419 B.n418 585
R236 B.n417 B.n416 585
R237 B.n415 B.n414 585
R238 B.n413 B.n412 585
R239 B.n410 B.n409 585
R240 B.n408 B.n407 585
R241 B.n406 B.n405 585
R242 B.n404 B.n403 585
R243 B.n402 B.n401 585
R244 B.n400 B.n399 585
R245 B.n398 B.n397 585
R246 B.n396 B.n395 585
R247 B.n394 B.n393 585
R248 B.n392 B.n391 585
R249 B.n390 B.n389 585
R250 B.n388 B.n387 585
R251 B.n386 B.n385 585
R252 B.n384 B.n383 585
R253 B.n382 B.n381 585
R254 B.n380 B.n379 585
R255 B.n378 B.n377 585
R256 B.n376 B.n375 585
R257 B.n374 B.n373 585
R258 B.n372 B.n371 585
R259 B.n370 B.n369 585
R260 B.n368 B.n367 585
R261 B.n366 B.n365 585
R262 B.n364 B.n363 585
R263 B.n362 B.n361 585
R264 B.n360 B.n359 585
R265 B.n358 B.n357 585
R266 B.n356 B.n355 585
R267 B.n354 B.n353 585
R268 B.n352 B.n351 585
R269 B.n350 B.n349 585
R270 B.n348 B.n347 585
R271 B.n346 B.n345 585
R272 B.n344 B.n343 585
R273 B.n342 B.n341 585
R274 B.n340 B.n339 585
R275 B.n338 B.n337 585
R276 B.n467 B.n297 585
R277 B.n297 B.n296 585
R278 B.n469 B.n468 585
R279 B.n470 B.n469 585
R280 B.n291 B.n290 585
R281 B.n292 B.n291 585
R282 B.n478 B.n477 585
R283 B.n477 B.n476 585
R284 B.n479 B.n289 585
R285 B.n289 B.n287 585
R286 B.n481 B.n480 585
R287 B.n482 B.n481 585
R288 B.n283 B.n282 585
R289 B.n288 B.n283 585
R290 B.n490 B.n489 585
R291 B.n489 B.n488 585
R292 B.n491 B.n281 585
R293 B.n281 B.n280 585
R294 B.n493 B.n492 585
R295 B.n494 B.n493 585
R296 B.n275 B.n274 585
R297 B.n276 B.n275 585
R298 B.n502 B.n501 585
R299 B.n501 B.n500 585
R300 B.n503 B.n273 585
R301 B.n273 B.n272 585
R302 B.n505 B.n504 585
R303 B.n506 B.n505 585
R304 B.n267 B.n266 585
R305 B.n268 B.n267 585
R306 B.n515 B.n514 585
R307 B.n514 B.n513 585
R308 B.n516 B.n265 585
R309 B.n512 B.n265 585
R310 B.n518 B.n517 585
R311 B.n519 B.n518 585
R312 B.n260 B.n259 585
R313 B.n261 B.n260 585
R314 B.n527 B.n526 585
R315 B.n526 B.n525 585
R316 B.n528 B.n258 585
R317 B.n258 B.n257 585
R318 B.n530 B.n529 585
R319 B.n531 B.n530 585
R320 B.n252 B.n251 585
R321 B.n253 B.n252 585
R322 B.n539 B.n538 585
R323 B.n538 B.n537 585
R324 B.n540 B.n250 585
R325 B.n250 B.n249 585
R326 B.n542 B.n541 585
R327 B.n543 B.n542 585
R328 B.n244 B.n243 585
R329 B.n245 B.n244 585
R330 B.n551 B.n550 585
R331 B.n550 B.n549 585
R332 B.n552 B.n242 585
R333 B.n242 B.n240 585
R334 B.n554 B.n553 585
R335 B.n555 B.n554 585
R336 B.n236 B.n235 585
R337 B.n241 B.n236 585
R338 B.n564 B.n563 585
R339 B.n563 B.n562 585
R340 B.n565 B.n234 585
R341 B.n234 B.n233 585
R342 B.n567 B.n566 585
R343 B.n568 B.n567 585
R344 B.n3 B.n0 585
R345 B.n4 B.n3 585
R346 B.n691 B.n1 585
R347 B.n692 B.n691 585
R348 B.n690 B.n689 585
R349 B.n690 B.n8 585
R350 B.n688 B.n9 585
R351 B.n12 B.n9 585
R352 B.n687 B.n686 585
R353 B.n686 B.n685 585
R354 B.n11 B.n10 585
R355 B.n684 B.n11 585
R356 B.n682 B.n681 585
R357 B.n683 B.n682 585
R358 B.n680 B.n17 585
R359 B.n17 B.n16 585
R360 B.n679 B.n678 585
R361 B.n678 B.n677 585
R362 B.n19 B.n18 585
R363 B.n676 B.n19 585
R364 B.n674 B.n673 585
R365 B.n675 B.n674 585
R366 B.n672 B.n24 585
R367 B.n24 B.n23 585
R368 B.n671 B.n670 585
R369 B.n670 B.n669 585
R370 B.n26 B.n25 585
R371 B.n668 B.n26 585
R372 B.n666 B.n665 585
R373 B.n667 B.n666 585
R374 B.n664 B.n31 585
R375 B.n31 B.n30 585
R376 B.n663 B.n662 585
R377 B.n662 B.n661 585
R378 B.n33 B.n32 585
R379 B.n660 B.n33 585
R380 B.n658 B.n657 585
R381 B.n659 B.n658 585
R382 B.n656 B.n37 585
R383 B.n40 B.n37 585
R384 B.n655 B.n654 585
R385 B.n654 B.n653 585
R386 B.n39 B.n38 585
R387 B.n652 B.n39 585
R388 B.n650 B.n649 585
R389 B.n651 B.n650 585
R390 B.n648 B.n45 585
R391 B.n45 B.n44 585
R392 B.n647 B.n646 585
R393 B.n646 B.n645 585
R394 B.n47 B.n46 585
R395 B.n644 B.n47 585
R396 B.n642 B.n641 585
R397 B.n643 B.n642 585
R398 B.n640 B.n52 585
R399 B.n52 B.n51 585
R400 B.n639 B.n638 585
R401 B.n638 B.n637 585
R402 B.n54 B.n53 585
R403 B.n636 B.n54 585
R404 B.n634 B.n633 585
R405 B.n635 B.n634 585
R406 B.n632 B.n59 585
R407 B.n59 B.n58 585
R408 B.n631 B.n630 585
R409 B.n630 B.n629 585
R410 B.n61 B.n60 585
R411 B.n628 B.n61 585
R412 B.n626 B.n625 585
R413 B.n627 B.n626 585
R414 B.n624 B.n66 585
R415 B.n66 B.n65 585
R416 B.n695 B.n694 585
R417 B.n693 B.n2 585
R418 B.n622 B.n66 492.5
R419 B.n619 B.n101 492.5
R420 B.n337 B.n295 492.5
R421 B.n465 B.n297 492.5
R422 B.n104 B.t17 294.281
R423 B.n102 B.t13 294.281
R424 B.n334 B.t10 294.281
R425 B.n332 B.t6 294.281
R426 B.n620 B.n99 256.663
R427 B.n620 B.n98 256.663
R428 B.n620 B.n97 256.663
R429 B.n620 B.n96 256.663
R430 B.n620 B.n95 256.663
R431 B.n620 B.n94 256.663
R432 B.n620 B.n93 256.663
R433 B.n620 B.n92 256.663
R434 B.n620 B.n91 256.663
R435 B.n620 B.n90 256.663
R436 B.n620 B.n89 256.663
R437 B.n620 B.n88 256.663
R438 B.n620 B.n87 256.663
R439 B.n620 B.n86 256.663
R440 B.n620 B.n85 256.663
R441 B.n620 B.n84 256.663
R442 B.n620 B.n83 256.663
R443 B.n620 B.n82 256.663
R444 B.n620 B.n81 256.663
R445 B.n620 B.n80 256.663
R446 B.n620 B.n79 256.663
R447 B.n620 B.n78 256.663
R448 B.n620 B.n77 256.663
R449 B.n620 B.n76 256.663
R450 B.n620 B.n75 256.663
R451 B.n620 B.n74 256.663
R452 B.n620 B.n73 256.663
R453 B.n620 B.n72 256.663
R454 B.n620 B.n71 256.663
R455 B.n620 B.n70 256.663
R456 B.n620 B.n69 256.663
R457 B.n621 B.n620 256.663
R458 B.n464 B.n463 256.663
R459 B.n463 B.n300 256.663
R460 B.n463 B.n301 256.663
R461 B.n463 B.n302 256.663
R462 B.n463 B.n303 256.663
R463 B.n463 B.n304 256.663
R464 B.n463 B.n305 256.663
R465 B.n463 B.n306 256.663
R466 B.n463 B.n307 256.663
R467 B.n463 B.n308 256.663
R468 B.n463 B.n309 256.663
R469 B.n463 B.n310 256.663
R470 B.n463 B.n311 256.663
R471 B.n463 B.n312 256.663
R472 B.n463 B.n313 256.663
R473 B.n463 B.n314 256.663
R474 B.n463 B.n315 256.663
R475 B.n463 B.n316 256.663
R476 B.n463 B.n317 256.663
R477 B.n463 B.n318 256.663
R478 B.n463 B.n319 256.663
R479 B.n463 B.n320 256.663
R480 B.n463 B.n321 256.663
R481 B.n463 B.n322 256.663
R482 B.n463 B.n323 256.663
R483 B.n463 B.n324 256.663
R484 B.n463 B.n325 256.663
R485 B.n463 B.n326 256.663
R486 B.n463 B.n327 256.663
R487 B.n463 B.n328 256.663
R488 B.n463 B.n329 256.663
R489 B.n463 B.n330 256.663
R490 B.n697 B.n696 256.663
R491 B.n102 B.t15 245.417
R492 B.n334 B.t12 245.417
R493 B.n104 B.t18 245.417
R494 B.n332 B.t9 245.417
R495 B.n103 B.t16 200.228
R496 B.n335 B.t11 200.228
R497 B.n105 B.t19 200.228
R498 B.n333 B.t8 200.228
R499 B.n107 B.n68 163.367
R500 B.n111 B.n110 163.367
R501 B.n115 B.n114 163.367
R502 B.n119 B.n118 163.367
R503 B.n123 B.n122 163.367
R504 B.n127 B.n126 163.367
R505 B.n131 B.n130 163.367
R506 B.n135 B.n134 163.367
R507 B.n139 B.n138 163.367
R508 B.n143 B.n142 163.367
R509 B.n147 B.n146 163.367
R510 B.n151 B.n150 163.367
R511 B.n155 B.n154 163.367
R512 B.n159 B.n158 163.367
R513 B.n163 B.n162 163.367
R514 B.n167 B.n166 163.367
R515 B.n171 B.n170 163.367
R516 B.n175 B.n174 163.367
R517 B.n180 B.n179 163.367
R518 B.n184 B.n183 163.367
R519 B.n188 B.n187 163.367
R520 B.n192 B.n191 163.367
R521 B.n196 B.n195 163.367
R522 B.n200 B.n199 163.367
R523 B.n204 B.n203 163.367
R524 B.n208 B.n207 163.367
R525 B.n212 B.n211 163.367
R526 B.n216 B.n215 163.367
R527 B.n220 B.n219 163.367
R528 B.n224 B.n223 163.367
R529 B.n228 B.n227 163.367
R530 B.n619 B.n100 163.367
R531 B.n471 B.n295 163.367
R532 B.n471 B.n293 163.367
R533 B.n475 B.n293 163.367
R534 B.n475 B.n286 163.367
R535 B.n483 B.n286 163.367
R536 B.n483 B.n284 163.367
R537 B.n487 B.n284 163.367
R538 B.n487 B.n279 163.367
R539 B.n495 B.n279 163.367
R540 B.n495 B.n277 163.367
R541 B.n499 B.n277 163.367
R542 B.n499 B.n271 163.367
R543 B.n507 B.n271 163.367
R544 B.n507 B.n269 163.367
R545 B.n511 B.n269 163.367
R546 B.n511 B.n264 163.367
R547 B.n520 B.n264 163.367
R548 B.n520 B.n262 163.367
R549 B.n524 B.n262 163.367
R550 B.n524 B.n256 163.367
R551 B.n532 B.n256 163.367
R552 B.n532 B.n254 163.367
R553 B.n536 B.n254 163.367
R554 B.n536 B.n248 163.367
R555 B.n544 B.n248 163.367
R556 B.n544 B.n246 163.367
R557 B.n548 B.n246 163.367
R558 B.n548 B.n239 163.367
R559 B.n556 B.n239 163.367
R560 B.n556 B.n237 163.367
R561 B.n561 B.n237 163.367
R562 B.n561 B.n232 163.367
R563 B.n569 B.n232 163.367
R564 B.n570 B.n569 163.367
R565 B.n570 B.n5 163.367
R566 B.n6 B.n5 163.367
R567 B.n7 B.n6 163.367
R568 B.n576 B.n7 163.367
R569 B.n577 B.n576 163.367
R570 B.n577 B.n13 163.367
R571 B.n14 B.n13 163.367
R572 B.n15 B.n14 163.367
R573 B.n582 B.n15 163.367
R574 B.n582 B.n20 163.367
R575 B.n21 B.n20 163.367
R576 B.n22 B.n21 163.367
R577 B.n587 B.n22 163.367
R578 B.n587 B.n27 163.367
R579 B.n28 B.n27 163.367
R580 B.n29 B.n28 163.367
R581 B.n592 B.n29 163.367
R582 B.n592 B.n34 163.367
R583 B.n35 B.n34 163.367
R584 B.n36 B.n35 163.367
R585 B.n597 B.n36 163.367
R586 B.n597 B.n41 163.367
R587 B.n42 B.n41 163.367
R588 B.n43 B.n42 163.367
R589 B.n602 B.n43 163.367
R590 B.n602 B.n48 163.367
R591 B.n49 B.n48 163.367
R592 B.n50 B.n49 163.367
R593 B.n607 B.n50 163.367
R594 B.n607 B.n55 163.367
R595 B.n56 B.n55 163.367
R596 B.n57 B.n56 163.367
R597 B.n612 B.n57 163.367
R598 B.n612 B.n62 163.367
R599 B.n63 B.n62 163.367
R600 B.n64 B.n63 163.367
R601 B.n101 B.n64 163.367
R602 B.n462 B.n299 163.367
R603 B.n462 B.n331 163.367
R604 B.n458 B.n457 163.367
R605 B.n454 B.n453 163.367
R606 B.n450 B.n449 163.367
R607 B.n446 B.n445 163.367
R608 B.n442 B.n441 163.367
R609 B.n438 B.n437 163.367
R610 B.n434 B.n433 163.367
R611 B.n430 B.n429 163.367
R612 B.n426 B.n425 163.367
R613 B.n422 B.n421 163.367
R614 B.n418 B.n417 163.367
R615 B.n414 B.n413 163.367
R616 B.n409 B.n408 163.367
R617 B.n405 B.n404 163.367
R618 B.n401 B.n400 163.367
R619 B.n397 B.n396 163.367
R620 B.n393 B.n392 163.367
R621 B.n389 B.n388 163.367
R622 B.n385 B.n384 163.367
R623 B.n381 B.n380 163.367
R624 B.n377 B.n376 163.367
R625 B.n373 B.n372 163.367
R626 B.n369 B.n368 163.367
R627 B.n365 B.n364 163.367
R628 B.n361 B.n360 163.367
R629 B.n357 B.n356 163.367
R630 B.n353 B.n352 163.367
R631 B.n349 B.n348 163.367
R632 B.n345 B.n344 163.367
R633 B.n341 B.n340 163.367
R634 B.n469 B.n297 163.367
R635 B.n469 B.n291 163.367
R636 B.n477 B.n291 163.367
R637 B.n477 B.n289 163.367
R638 B.n481 B.n289 163.367
R639 B.n481 B.n283 163.367
R640 B.n489 B.n283 163.367
R641 B.n489 B.n281 163.367
R642 B.n493 B.n281 163.367
R643 B.n493 B.n275 163.367
R644 B.n501 B.n275 163.367
R645 B.n501 B.n273 163.367
R646 B.n505 B.n273 163.367
R647 B.n505 B.n267 163.367
R648 B.n514 B.n267 163.367
R649 B.n514 B.n265 163.367
R650 B.n518 B.n265 163.367
R651 B.n518 B.n260 163.367
R652 B.n526 B.n260 163.367
R653 B.n526 B.n258 163.367
R654 B.n530 B.n258 163.367
R655 B.n530 B.n252 163.367
R656 B.n538 B.n252 163.367
R657 B.n538 B.n250 163.367
R658 B.n542 B.n250 163.367
R659 B.n542 B.n244 163.367
R660 B.n550 B.n244 163.367
R661 B.n550 B.n242 163.367
R662 B.n554 B.n242 163.367
R663 B.n554 B.n236 163.367
R664 B.n563 B.n236 163.367
R665 B.n563 B.n234 163.367
R666 B.n567 B.n234 163.367
R667 B.n567 B.n3 163.367
R668 B.n695 B.n3 163.367
R669 B.n691 B.n2 163.367
R670 B.n691 B.n690 163.367
R671 B.n690 B.n9 163.367
R672 B.n686 B.n9 163.367
R673 B.n686 B.n11 163.367
R674 B.n682 B.n11 163.367
R675 B.n682 B.n17 163.367
R676 B.n678 B.n17 163.367
R677 B.n678 B.n19 163.367
R678 B.n674 B.n19 163.367
R679 B.n674 B.n24 163.367
R680 B.n670 B.n24 163.367
R681 B.n670 B.n26 163.367
R682 B.n666 B.n26 163.367
R683 B.n666 B.n31 163.367
R684 B.n662 B.n31 163.367
R685 B.n662 B.n33 163.367
R686 B.n658 B.n33 163.367
R687 B.n658 B.n37 163.367
R688 B.n654 B.n37 163.367
R689 B.n654 B.n39 163.367
R690 B.n650 B.n39 163.367
R691 B.n650 B.n45 163.367
R692 B.n646 B.n45 163.367
R693 B.n646 B.n47 163.367
R694 B.n642 B.n47 163.367
R695 B.n642 B.n52 163.367
R696 B.n638 B.n52 163.367
R697 B.n638 B.n54 163.367
R698 B.n634 B.n54 163.367
R699 B.n634 B.n59 163.367
R700 B.n630 B.n59 163.367
R701 B.n630 B.n61 163.367
R702 B.n626 B.n61 163.367
R703 B.n626 B.n66 163.367
R704 B.n463 B.n296 109.781
R705 B.n620 B.n65 109.781
R706 B.n622 B.n621 71.676
R707 B.n107 B.n69 71.676
R708 B.n111 B.n70 71.676
R709 B.n115 B.n71 71.676
R710 B.n119 B.n72 71.676
R711 B.n123 B.n73 71.676
R712 B.n127 B.n74 71.676
R713 B.n131 B.n75 71.676
R714 B.n135 B.n76 71.676
R715 B.n139 B.n77 71.676
R716 B.n143 B.n78 71.676
R717 B.n147 B.n79 71.676
R718 B.n151 B.n80 71.676
R719 B.n155 B.n81 71.676
R720 B.n159 B.n82 71.676
R721 B.n163 B.n83 71.676
R722 B.n167 B.n84 71.676
R723 B.n171 B.n85 71.676
R724 B.n175 B.n86 71.676
R725 B.n180 B.n87 71.676
R726 B.n184 B.n88 71.676
R727 B.n188 B.n89 71.676
R728 B.n192 B.n90 71.676
R729 B.n196 B.n91 71.676
R730 B.n200 B.n92 71.676
R731 B.n204 B.n93 71.676
R732 B.n208 B.n94 71.676
R733 B.n212 B.n95 71.676
R734 B.n216 B.n96 71.676
R735 B.n220 B.n97 71.676
R736 B.n224 B.n98 71.676
R737 B.n228 B.n99 71.676
R738 B.n100 B.n99 71.676
R739 B.n227 B.n98 71.676
R740 B.n223 B.n97 71.676
R741 B.n219 B.n96 71.676
R742 B.n215 B.n95 71.676
R743 B.n211 B.n94 71.676
R744 B.n207 B.n93 71.676
R745 B.n203 B.n92 71.676
R746 B.n199 B.n91 71.676
R747 B.n195 B.n90 71.676
R748 B.n191 B.n89 71.676
R749 B.n187 B.n88 71.676
R750 B.n183 B.n87 71.676
R751 B.n179 B.n86 71.676
R752 B.n174 B.n85 71.676
R753 B.n170 B.n84 71.676
R754 B.n166 B.n83 71.676
R755 B.n162 B.n82 71.676
R756 B.n158 B.n81 71.676
R757 B.n154 B.n80 71.676
R758 B.n150 B.n79 71.676
R759 B.n146 B.n78 71.676
R760 B.n142 B.n77 71.676
R761 B.n138 B.n76 71.676
R762 B.n134 B.n75 71.676
R763 B.n130 B.n74 71.676
R764 B.n126 B.n73 71.676
R765 B.n122 B.n72 71.676
R766 B.n118 B.n71 71.676
R767 B.n114 B.n70 71.676
R768 B.n110 B.n69 71.676
R769 B.n621 B.n68 71.676
R770 B.n465 B.n464 71.676
R771 B.n331 B.n300 71.676
R772 B.n457 B.n301 71.676
R773 B.n453 B.n302 71.676
R774 B.n449 B.n303 71.676
R775 B.n445 B.n304 71.676
R776 B.n441 B.n305 71.676
R777 B.n437 B.n306 71.676
R778 B.n433 B.n307 71.676
R779 B.n429 B.n308 71.676
R780 B.n425 B.n309 71.676
R781 B.n421 B.n310 71.676
R782 B.n417 B.n311 71.676
R783 B.n413 B.n312 71.676
R784 B.n408 B.n313 71.676
R785 B.n404 B.n314 71.676
R786 B.n400 B.n315 71.676
R787 B.n396 B.n316 71.676
R788 B.n392 B.n317 71.676
R789 B.n388 B.n318 71.676
R790 B.n384 B.n319 71.676
R791 B.n380 B.n320 71.676
R792 B.n376 B.n321 71.676
R793 B.n372 B.n322 71.676
R794 B.n368 B.n323 71.676
R795 B.n364 B.n324 71.676
R796 B.n360 B.n325 71.676
R797 B.n356 B.n326 71.676
R798 B.n352 B.n327 71.676
R799 B.n348 B.n328 71.676
R800 B.n344 B.n329 71.676
R801 B.n340 B.n330 71.676
R802 B.n464 B.n299 71.676
R803 B.n458 B.n300 71.676
R804 B.n454 B.n301 71.676
R805 B.n450 B.n302 71.676
R806 B.n446 B.n303 71.676
R807 B.n442 B.n304 71.676
R808 B.n438 B.n305 71.676
R809 B.n434 B.n306 71.676
R810 B.n430 B.n307 71.676
R811 B.n426 B.n308 71.676
R812 B.n422 B.n309 71.676
R813 B.n418 B.n310 71.676
R814 B.n414 B.n311 71.676
R815 B.n409 B.n312 71.676
R816 B.n405 B.n313 71.676
R817 B.n401 B.n314 71.676
R818 B.n397 B.n315 71.676
R819 B.n393 B.n316 71.676
R820 B.n389 B.n317 71.676
R821 B.n385 B.n318 71.676
R822 B.n381 B.n319 71.676
R823 B.n377 B.n320 71.676
R824 B.n373 B.n321 71.676
R825 B.n369 B.n322 71.676
R826 B.n365 B.n323 71.676
R827 B.n361 B.n324 71.676
R828 B.n357 B.n325 71.676
R829 B.n353 B.n326 71.676
R830 B.n349 B.n327 71.676
R831 B.n345 B.n328 71.676
R832 B.n341 B.n329 71.676
R833 B.n337 B.n330 71.676
R834 B.n696 B.n695 71.676
R835 B.n696 B.n2 71.676
R836 B.n470 B.n296 59.7211
R837 B.n470 B.n292 59.7211
R838 B.n476 B.n292 59.7211
R839 B.n476 B.n287 59.7211
R840 B.n482 B.n287 59.7211
R841 B.n482 B.n288 59.7211
R842 B.n488 B.n280 59.7211
R843 B.n494 B.n280 59.7211
R844 B.n494 B.n276 59.7211
R845 B.n500 B.n276 59.7211
R846 B.n500 B.n272 59.7211
R847 B.n506 B.n272 59.7211
R848 B.n506 B.n268 59.7211
R849 B.n513 B.n268 59.7211
R850 B.n513 B.n512 59.7211
R851 B.n519 B.n261 59.7211
R852 B.n525 B.n261 59.7211
R853 B.n525 B.n257 59.7211
R854 B.n531 B.n257 59.7211
R855 B.n531 B.n253 59.7211
R856 B.n537 B.n253 59.7211
R857 B.n543 B.n249 59.7211
R858 B.n543 B.n245 59.7211
R859 B.n549 B.n245 59.7211
R860 B.n549 B.n240 59.7211
R861 B.n555 B.n240 59.7211
R862 B.n555 B.n241 59.7211
R863 B.n562 B.n233 59.7211
R864 B.n568 B.n233 59.7211
R865 B.n568 B.n4 59.7211
R866 B.n694 B.n4 59.7211
R867 B.n694 B.n693 59.7211
R868 B.n693 B.n692 59.7211
R869 B.n692 B.n8 59.7211
R870 B.n12 B.n8 59.7211
R871 B.n685 B.n12 59.7211
R872 B.n684 B.n683 59.7211
R873 B.n683 B.n16 59.7211
R874 B.n677 B.n16 59.7211
R875 B.n677 B.n676 59.7211
R876 B.n676 B.n675 59.7211
R877 B.n675 B.n23 59.7211
R878 B.n669 B.n668 59.7211
R879 B.n668 B.n667 59.7211
R880 B.n667 B.n30 59.7211
R881 B.n661 B.n30 59.7211
R882 B.n661 B.n660 59.7211
R883 B.n660 B.n659 59.7211
R884 B.n653 B.n40 59.7211
R885 B.n653 B.n652 59.7211
R886 B.n652 B.n651 59.7211
R887 B.n651 B.n44 59.7211
R888 B.n645 B.n44 59.7211
R889 B.n645 B.n644 59.7211
R890 B.n644 B.n643 59.7211
R891 B.n643 B.n51 59.7211
R892 B.n637 B.n51 59.7211
R893 B.n636 B.n635 59.7211
R894 B.n635 B.n58 59.7211
R895 B.n629 B.n58 59.7211
R896 B.n629 B.n628 59.7211
R897 B.n628 B.n627 59.7211
R898 B.n627 B.n65 59.7211
R899 B.n106 B.n105 59.5399
R900 B.n177 B.n103 59.5399
R901 B.n336 B.n335 59.5399
R902 B.n411 B.n333 59.5399
R903 B.n512 B.t2 45.6692
R904 B.n40 B.t5 45.6692
R905 B.n105 B.n104 45.1884
R906 B.n103 B.n102 45.1884
R907 B.n335 B.n334 45.1884
R908 B.n333 B.n332 45.1884
R909 B.n288 B.t7 42.1562
R910 B.t14 B.n636 42.1562
R911 B.n537 B.t1 36.8867
R912 B.n669 B.t4 36.8867
R913 B.n467 B.n466 32.0005
R914 B.n338 B.n294 32.0005
R915 B.n618 B.n617 32.0005
R916 B.n624 B.n623 32.0005
R917 B.n562 B.t0 31.6173
R918 B.n685 B.t3 31.6173
R919 B.n241 B.t0 28.1043
R920 B.t3 B.n684 28.1043
R921 B.t1 B.n249 22.8348
R922 B.t4 B.n23 22.8348
R923 B B.n697 18.0485
R924 B.n488 B.t7 17.5654
R925 B.n637 B.t14 17.5654
R926 B.n519 B.t2 14.0524
R927 B.n659 B.t5 14.0524
R928 B.n468 B.n467 10.6151
R929 B.n468 B.n290 10.6151
R930 B.n478 B.n290 10.6151
R931 B.n479 B.n478 10.6151
R932 B.n480 B.n479 10.6151
R933 B.n480 B.n282 10.6151
R934 B.n490 B.n282 10.6151
R935 B.n491 B.n490 10.6151
R936 B.n492 B.n491 10.6151
R937 B.n492 B.n274 10.6151
R938 B.n502 B.n274 10.6151
R939 B.n503 B.n502 10.6151
R940 B.n504 B.n503 10.6151
R941 B.n504 B.n266 10.6151
R942 B.n515 B.n266 10.6151
R943 B.n516 B.n515 10.6151
R944 B.n517 B.n516 10.6151
R945 B.n517 B.n259 10.6151
R946 B.n527 B.n259 10.6151
R947 B.n528 B.n527 10.6151
R948 B.n529 B.n528 10.6151
R949 B.n529 B.n251 10.6151
R950 B.n539 B.n251 10.6151
R951 B.n540 B.n539 10.6151
R952 B.n541 B.n540 10.6151
R953 B.n541 B.n243 10.6151
R954 B.n551 B.n243 10.6151
R955 B.n552 B.n551 10.6151
R956 B.n553 B.n552 10.6151
R957 B.n553 B.n235 10.6151
R958 B.n564 B.n235 10.6151
R959 B.n565 B.n564 10.6151
R960 B.n566 B.n565 10.6151
R961 B.n566 B.n0 10.6151
R962 B.n466 B.n298 10.6151
R963 B.n461 B.n298 10.6151
R964 B.n461 B.n460 10.6151
R965 B.n460 B.n459 10.6151
R966 B.n459 B.n456 10.6151
R967 B.n456 B.n455 10.6151
R968 B.n455 B.n452 10.6151
R969 B.n452 B.n451 10.6151
R970 B.n451 B.n448 10.6151
R971 B.n448 B.n447 10.6151
R972 B.n447 B.n444 10.6151
R973 B.n444 B.n443 10.6151
R974 B.n443 B.n440 10.6151
R975 B.n440 B.n439 10.6151
R976 B.n439 B.n436 10.6151
R977 B.n436 B.n435 10.6151
R978 B.n435 B.n432 10.6151
R979 B.n432 B.n431 10.6151
R980 B.n431 B.n428 10.6151
R981 B.n428 B.n427 10.6151
R982 B.n427 B.n424 10.6151
R983 B.n424 B.n423 10.6151
R984 B.n423 B.n420 10.6151
R985 B.n420 B.n419 10.6151
R986 B.n419 B.n416 10.6151
R987 B.n416 B.n415 10.6151
R988 B.n415 B.n412 10.6151
R989 B.n410 B.n407 10.6151
R990 B.n407 B.n406 10.6151
R991 B.n406 B.n403 10.6151
R992 B.n403 B.n402 10.6151
R993 B.n402 B.n399 10.6151
R994 B.n399 B.n398 10.6151
R995 B.n398 B.n395 10.6151
R996 B.n395 B.n394 10.6151
R997 B.n391 B.n390 10.6151
R998 B.n390 B.n387 10.6151
R999 B.n387 B.n386 10.6151
R1000 B.n386 B.n383 10.6151
R1001 B.n383 B.n382 10.6151
R1002 B.n382 B.n379 10.6151
R1003 B.n379 B.n378 10.6151
R1004 B.n378 B.n375 10.6151
R1005 B.n375 B.n374 10.6151
R1006 B.n374 B.n371 10.6151
R1007 B.n371 B.n370 10.6151
R1008 B.n370 B.n367 10.6151
R1009 B.n367 B.n366 10.6151
R1010 B.n366 B.n363 10.6151
R1011 B.n363 B.n362 10.6151
R1012 B.n362 B.n359 10.6151
R1013 B.n359 B.n358 10.6151
R1014 B.n358 B.n355 10.6151
R1015 B.n355 B.n354 10.6151
R1016 B.n354 B.n351 10.6151
R1017 B.n351 B.n350 10.6151
R1018 B.n350 B.n347 10.6151
R1019 B.n347 B.n346 10.6151
R1020 B.n346 B.n343 10.6151
R1021 B.n343 B.n342 10.6151
R1022 B.n342 B.n339 10.6151
R1023 B.n339 B.n338 10.6151
R1024 B.n472 B.n294 10.6151
R1025 B.n473 B.n472 10.6151
R1026 B.n474 B.n473 10.6151
R1027 B.n474 B.n285 10.6151
R1028 B.n484 B.n285 10.6151
R1029 B.n485 B.n484 10.6151
R1030 B.n486 B.n485 10.6151
R1031 B.n486 B.n278 10.6151
R1032 B.n496 B.n278 10.6151
R1033 B.n497 B.n496 10.6151
R1034 B.n498 B.n497 10.6151
R1035 B.n498 B.n270 10.6151
R1036 B.n508 B.n270 10.6151
R1037 B.n509 B.n508 10.6151
R1038 B.n510 B.n509 10.6151
R1039 B.n510 B.n263 10.6151
R1040 B.n521 B.n263 10.6151
R1041 B.n522 B.n521 10.6151
R1042 B.n523 B.n522 10.6151
R1043 B.n523 B.n255 10.6151
R1044 B.n533 B.n255 10.6151
R1045 B.n534 B.n533 10.6151
R1046 B.n535 B.n534 10.6151
R1047 B.n535 B.n247 10.6151
R1048 B.n545 B.n247 10.6151
R1049 B.n546 B.n545 10.6151
R1050 B.n547 B.n546 10.6151
R1051 B.n547 B.n238 10.6151
R1052 B.n557 B.n238 10.6151
R1053 B.n558 B.n557 10.6151
R1054 B.n560 B.n558 10.6151
R1055 B.n560 B.n559 10.6151
R1056 B.n559 B.n231 10.6151
R1057 B.n571 B.n231 10.6151
R1058 B.n572 B.n571 10.6151
R1059 B.n573 B.n572 10.6151
R1060 B.n574 B.n573 10.6151
R1061 B.n575 B.n574 10.6151
R1062 B.n578 B.n575 10.6151
R1063 B.n579 B.n578 10.6151
R1064 B.n580 B.n579 10.6151
R1065 B.n581 B.n580 10.6151
R1066 B.n583 B.n581 10.6151
R1067 B.n584 B.n583 10.6151
R1068 B.n585 B.n584 10.6151
R1069 B.n586 B.n585 10.6151
R1070 B.n588 B.n586 10.6151
R1071 B.n589 B.n588 10.6151
R1072 B.n590 B.n589 10.6151
R1073 B.n591 B.n590 10.6151
R1074 B.n593 B.n591 10.6151
R1075 B.n594 B.n593 10.6151
R1076 B.n595 B.n594 10.6151
R1077 B.n596 B.n595 10.6151
R1078 B.n598 B.n596 10.6151
R1079 B.n599 B.n598 10.6151
R1080 B.n600 B.n599 10.6151
R1081 B.n601 B.n600 10.6151
R1082 B.n603 B.n601 10.6151
R1083 B.n604 B.n603 10.6151
R1084 B.n605 B.n604 10.6151
R1085 B.n606 B.n605 10.6151
R1086 B.n608 B.n606 10.6151
R1087 B.n609 B.n608 10.6151
R1088 B.n610 B.n609 10.6151
R1089 B.n611 B.n610 10.6151
R1090 B.n613 B.n611 10.6151
R1091 B.n614 B.n613 10.6151
R1092 B.n615 B.n614 10.6151
R1093 B.n616 B.n615 10.6151
R1094 B.n617 B.n616 10.6151
R1095 B.n689 B.n1 10.6151
R1096 B.n689 B.n688 10.6151
R1097 B.n688 B.n687 10.6151
R1098 B.n687 B.n10 10.6151
R1099 B.n681 B.n10 10.6151
R1100 B.n681 B.n680 10.6151
R1101 B.n680 B.n679 10.6151
R1102 B.n679 B.n18 10.6151
R1103 B.n673 B.n18 10.6151
R1104 B.n673 B.n672 10.6151
R1105 B.n672 B.n671 10.6151
R1106 B.n671 B.n25 10.6151
R1107 B.n665 B.n25 10.6151
R1108 B.n665 B.n664 10.6151
R1109 B.n664 B.n663 10.6151
R1110 B.n663 B.n32 10.6151
R1111 B.n657 B.n32 10.6151
R1112 B.n657 B.n656 10.6151
R1113 B.n656 B.n655 10.6151
R1114 B.n655 B.n38 10.6151
R1115 B.n649 B.n38 10.6151
R1116 B.n649 B.n648 10.6151
R1117 B.n648 B.n647 10.6151
R1118 B.n647 B.n46 10.6151
R1119 B.n641 B.n46 10.6151
R1120 B.n641 B.n640 10.6151
R1121 B.n640 B.n639 10.6151
R1122 B.n639 B.n53 10.6151
R1123 B.n633 B.n53 10.6151
R1124 B.n633 B.n632 10.6151
R1125 B.n632 B.n631 10.6151
R1126 B.n631 B.n60 10.6151
R1127 B.n625 B.n60 10.6151
R1128 B.n625 B.n624 10.6151
R1129 B.n623 B.n67 10.6151
R1130 B.n108 B.n67 10.6151
R1131 B.n109 B.n108 10.6151
R1132 B.n112 B.n109 10.6151
R1133 B.n113 B.n112 10.6151
R1134 B.n116 B.n113 10.6151
R1135 B.n117 B.n116 10.6151
R1136 B.n120 B.n117 10.6151
R1137 B.n121 B.n120 10.6151
R1138 B.n124 B.n121 10.6151
R1139 B.n125 B.n124 10.6151
R1140 B.n128 B.n125 10.6151
R1141 B.n129 B.n128 10.6151
R1142 B.n132 B.n129 10.6151
R1143 B.n133 B.n132 10.6151
R1144 B.n136 B.n133 10.6151
R1145 B.n137 B.n136 10.6151
R1146 B.n140 B.n137 10.6151
R1147 B.n141 B.n140 10.6151
R1148 B.n144 B.n141 10.6151
R1149 B.n145 B.n144 10.6151
R1150 B.n148 B.n145 10.6151
R1151 B.n149 B.n148 10.6151
R1152 B.n152 B.n149 10.6151
R1153 B.n153 B.n152 10.6151
R1154 B.n156 B.n153 10.6151
R1155 B.n157 B.n156 10.6151
R1156 B.n161 B.n160 10.6151
R1157 B.n164 B.n161 10.6151
R1158 B.n165 B.n164 10.6151
R1159 B.n168 B.n165 10.6151
R1160 B.n169 B.n168 10.6151
R1161 B.n172 B.n169 10.6151
R1162 B.n173 B.n172 10.6151
R1163 B.n176 B.n173 10.6151
R1164 B.n181 B.n178 10.6151
R1165 B.n182 B.n181 10.6151
R1166 B.n185 B.n182 10.6151
R1167 B.n186 B.n185 10.6151
R1168 B.n189 B.n186 10.6151
R1169 B.n190 B.n189 10.6151
R1170 B.n193 B.n190 10.6151
R1171 B.n194 B.n193 10.6151
R1172 B.n197 B.n194 10.6151
R1173 B.n198 B.n197 10.6151
R1174 B.n201 B.n198 10.6151
R1175 B.n202 B.n201 10.6151
R1176 B.n205 B.n202 10.6151
R1177 B.n206 B.n205 10.6151
R1178 B.n209 B.n206 10.6151
R1179 B.n210 B.n209 10.6151
R1180 B.n213 B.n210 10.6151
R1181 B.n214 B.n213 10.6151
R1182 B.n217 B.n214 10.6151
R1183 B.n218 B.n217 10.6151
R1184 B.n221 B.n218 10.6151
R1185 B.n222 B.n221 10.6151
R1186 B.n225 B.n222 10.6151
R1187 B.n226 B.n225 10.6151
R1188 B.n229 B.n226 10.6151
R1189 B.n230 B.n229 10.6151
R1190 B.n618 B.n230 10.6151
R1191 B.n697 B.n0 8.11757
R1192 B.n697 B.n1 8.11757
R1193 B.n411 B.n410 6.5566
R1194 B.n394 B.n336 6.5566
R1195 B.n160 B.n106 6.5566
R1196 B.n177 B.n176 6.5566
R1197 B.n412 B.n411 4.05904
R1198 B.n391 B.n336 4.05904
R1199 B.n157 B.n106 4.05904
R1200 B.n178 B.n177 4.05904
R1201 VN.n21 VN.n12 161.3
R1202 VN.n20 VN.n19 161.3
R1203 VN.n18 VN.n13 161.3
R1204 VN.n17 VN.n16 161.3
R1205 VN.n9 VN.n0 161.3
R1206 VN.n8 VN.n7 161.3
R1207 VN.n6 VN.n1 161.3
R1208 VN.n5 VN.n4 161.3
R1209 VN.n2 VN.t0 120.799
R1210 VN.n14 VN.t3 120.799
R1211 VN.n11 VN.n10 94.6082
R1212 VN.n23 VN.n22 94.6082
R1213 VN.n3 VN.t4 87.363
R1214 VN.n10 VN.t5 87.363
R1215 VN.n15 VN.t1 87.363
R1216 VN.n22 VN.t2 87.363
R1217 VN.n8 VN.n1 56.5193
R1218 VN.n20 VN.n13 56.5193
R1219 VN.n15 VN.n14 45.7103
R1220 VN.n3 VN.n2 45.7103
R1221 VN VN.n23 42.9716
R1222 VN.n4 VN.n3 24.4675
R1223 VN.n4 VN.n1 24.4675
R1224 VN.n9 VN.n8 24.4675
R1225 VN.n16 VN.n13 24.4675
R1226 VN.n16 VN.n15 24.4675
R1227 VN.n21 VN.n20 24.4675
R1228 VN.n10 VN.n9 16.1487
R1229 VN.n22 VN.n21 16.1487
R1230 VN.n17 VN.n14 9.33007
R1231 VN.n5 VN.n2 9.33007
R1232 VN.n23 VN.n12 0.278367
R1233 VN.n11 VN.n0 0.278367
R1234 VN.n19 VN.n12 0.189894
R1235 VN.n19 VN.n18 0.189894
R1236 VN.n18 VN.n17 0.189894
R1237 VN.n6 VN.n5 0.189894
R1238 VN.n7 VN.n6 0.189894
R1239 VN.n7 VN.n0 0.189894
R1240 VN VN.n11 0.153454
R1241 VTAIL.n146 VTAIL.n116 214.453
R1242 VTAIL.n32 VTAIL.n2 214.453
R1243 VTAIL.n110 VTAIL.n80 214.453
R1244 VTAIL.n72 VTAIL.n42 214.453
R1245 VTAIL.n129 VTAIL.n128 185
R1246 VTAIL.n131 VTAIL.n130 185
R1247 VTAIL.n124 VTAIL.n123 185
R1248 VTAIL.n137 VTAIL.n136 185
R1249 VTAIL.n139 VTAIL.n138 185
R1250 VTAIL.n120 VTAIL.n119 185
R1251 VTAIL.n145 VTAIL.n144 185
R1252 VTAIL.n147 VTAIL.n146 185
R1253 VTAIL.n15 VTAIL.n14 185
R1254 VTAIL.n17 VTAIL.n16 185
R1255 VTAIL.n10 VTAIL.n9 185
R1256 VTAIL.n23 VTAIL.n22 185
R1257 VTAIL.n25 VTAIL.n24 185
R1258 VTAIL.n6 VTAIL.n5 185
R1259 VTAIL.n31 VTAIL.n30 185
R1260 VTAIL.n33 VTAIL.n32 185
R1261 VTAIL.n111 VTAIL.n110 185
R1262 VTAIL.n109 VTAIL.n108 185
R1263 VTAIL.n84 VTAIL.n83 185
R1264 VTAIL.n103 VTAIL.n102 185
R1265 VTAIL.n101 VTAIL.n100 185
R1266 VTAIL.n88 VTAIL.n87 185
R1267 VTAIL.n95 VTAIL.n94 185
R1268 VTAIL.n93 VTAIL.n92 185
R1269 VTAIL.n73 VTAIL.n72 185
R1270 VTAIL.n71 VTAIL.n70 185
R1271 VTAIL.n46 VTAIL.n45 185
R1272 VTAIL.n65 VTAIL.n64 185
R1273 VTAIL.n63 VTAIL.n62 185
R1274 VTAIL.n50 VTAIL.n49 185
R1275 VTAIL.n57 VTAIL.n56 185
R1276 VTAIL.n55 VTAIL.n54 185
R1277 VTAIL.n127 VTAIL.t10 149.524
R1278 VTAIL.n13 VTAIL.t4 149.524
R1279 VTAIL.n91 VTAIL.t3 149.524
R1280 VTAIL.n53 VTAIL.t8 149.524
R1281 VTAIL.n130 VTAIL.n129 104.615
R1282 VTAIL.n130 VTAIL.n123 104.615
R1283 VTAIL.n137 VTAIL.n123 104.615
R1284 VTAIL.n138 VTAIL.n137 104.615
R1285 VTAIL.n138 VTAIL.n119 104.615
R1286 VTAIL.n145 VTAIL.n119 104.615
R1287 VTAIL.n146 VTAIL.n145 104.615
R1288 VTAIL.n16 VTAIL.n15 104.615
R1289 VTAIL.n16 VTAIL.n9 104.615
R1290 VTAIL.n23 VTAIL.n9 104.615
R1291 VTAIL.n24 VTAIL.n23 104.615
R1292 VTAIL.n24 VTAIL.n5 104.615
R1293 VTAIL.n31 VTAIL.n5 104.615
R1294 VTAIL.n32 VTAIL.n31 104.615
R1295 VTAIL.n110 VTAIL.n109 104.615
R1296 VTAIL.n109 VTAIL.n83 104.615
R1297 VTAIL.n102 VTAIL.n83 104.615
R1298 VTAIL.n102 VTAIL.n101 104.615
R1299 VTAIL.n101 VTAIL.n87 104.615
R1300 VTAIL.n94 VTAIL.n87 104.615
R1301 VTAIL.n94 VTAIL.n93 104.615
R1302 VTAIL.n72 VTAIL.n71 104.615
R1303 VTAIL.n71 VTAIL.n45 104.615
R1304 VTAIL.n64 VTAIL.n45 104.615
R1305 VTAIL.n64 VTAIL.n63 104.615
R1306 VTAIL.n63 VTAIL.n49 104.615
R1307 VTAIL.n56 VTAIL.n49 104.615
R1308 VTAIL.n56 VTAIL.n55 104.615
R1309 VTAIL.n129 VTAIL.t10 52.3082
R1310 VTAIL.n15 VTAIL.t4 52.3082
R1311 VTAIL.n93 VTAIL.t3 52.3082
R1312 VTAIL.n55 VTAIL.t8 52.3082
R1313 VTAIL.n79 VTAIL.n78 51.2531
R1314 VTAIL.n41 VTAIL.n40 51.2531
R1315 VTAIL.n1 VTAIL.n0 51.253
R1316 VTAIL.n39 VTAIL.n38 51.253
R1317 VTAIL.n151 VTAIL.n150 35.4823
R1318 VTAIL.n37 VTAIL.n36 35.4823
R1319 VTAIL.n115 VTAIL.n114 35.4823
R1320 VTAIL.n77 VTAIL.n76 35.4823
R1321 VTAIL.n41 VTAIL.n39 22.6341
R1322 VTAIL.n151 VTAIL.n115 20.6255
R1323 VTAIL.n148 VTAIL.n147 12.8005
R1324 VTAIL.n34 VTAIL.n33 12.8005
R1325 VTAIL.n112 VTAIL.n111 12.8005
R1326 VTAIL.n74 VTAIL.n73 12.8005
R1327 VTAIL.n144 VTAIL.n118 12.0247
R1328 VTAIL.n30 VTAIL.n4 12.0247
R1329 VTAIL.n108 VTAIL.n82 12.0247
R1330 VTAIL.n70 VTAIL.n44 12.0247
R1331 VTAIL.n143 VTAIL.n120 11.249
R1332 VTAIL.n29 VTAIL.n6 11.249
R1333 VTAIL.n107 VTAIL.n84 11.249
R1334 VTAIL.n69 VTAIL.n46 11.249
R1335 VTAIL.n140 VTAIL.n139 10.4732
R1336 VTAIL.n26 VTAIL.n25 10.4732
R1337 VTAIL.n104 VTAIL.n103 10.4732
R1338 VTAIL.n66 VTAIL.n65 10.4732
R1339 VTAIL.n128 VTAIL.n127 10.2747
R1340 VTAIL.n14 VTAIL.n13 10.2747
R1341 VTAIL.n92 VTAIL.n91 10.2747
R1342 VTAIL.n54 VTAIL.n53 10.2747
R1343 VTAIL.n136 VTAIL.n122 9.69747
R1344 VTAIL.n22 VTAIL.n8 9.69747
R1345 VTAIL.n100 VTAIL.n86 9.69747
R1346 VTAIL.n62 VTAIL.n48 9.69747
R1347 VTAIL.n150 VTAIL.n149 9.45567
R1348 VTAIL.n36 VTAIL.n35 9.45567
R1349 VTAIL.n114 VTAIL.n113 9.45567
R1350 VTAIL.n76 VTAIL.n75 9.45567
R1351 VTAIL.n126 VTAIL.n125 9.3005
R1352 VTAIL.n133 VTAIL.n132 9.3005
R1353 VTAIL.n135 VTAIL.n134 9.3005
R1354 VTAIL.n122 VTAIL.n121 9.3005
R1355 VTAIL.n141 VTAIL.n140 9.3005
R1356 VTAIL.n143 VTAIL.n142 9.3005
R1357 VTAIL.n118 VTAIL.n117 9.3005
R1358 VTAIL.n149 VTAIL.n148 9.3005
R1359 VTAIL.n12 VTAIL.n11 9.3005
R1360 VTAIL.n19 VTAIL.n18 9.3005
R1361 VTAIL.n21 VTAIL.n20 9.3005
R1362 VTAIL.n8 VTAIL.n7 9.3005
R1363 VTAIL.n27 VTAIL.n26 9.3005
R1364 VTAIL.n29 VTAIL.n28 9.3005
R1365 VTAIL.n4 VTAIL.n3 9.3005
R1366 VTAIL.n35 VTAIL.n34 9.3005
R1367 VTAIL.n90 VTAIL.n89 9.3005
R1368 VTAIL.n97 VTAIL.n96 9.3005
R1369 VTAIL.n99 VTAIL.n98 9.3005
R1370 VTAIL.n86 VTAIL.n85 9.3005
R1371 VTAIL.n105 VTAIL.n104 9.3005
R1372 VTAIL.n107 VTAIL.n106 9.3005
R1373 VTAIL.n82 VTAIL.n81 9.3005
R1374 VTAIL.n113 VTAIL.n112 9.3005
R1375 VTAIL.n52 VTAIL.n51 9.3005
R1376 VTAIL.n59 VTAIL.n58 9.3005
R1377 VTAIL.n61 VTAIL.n60 9.3005
R1378 VTAIL.n48 VTAIL.n47 9.3005
R1379 VTAIL.n67 VTAIL.n66 9.3005
R1380 VTAIL.n69 VTAIL.n68 9.3005
R1381 VTAIL.n44 VTAIL.n43 9.3005
R1382 VTAIL.n75 VTAIL.n74 9.3005
R1383 VTAIL.n135 VTAIL.n124 8.92171
R1384 VTAIL.n21 VTAIL.n10 8.92171
R1385 VTAIL.n99 VTAIL.n88 8.92171
R1386 VTAIL.n61 VTAIL.n50 8.92171
R1387 VTAIL.n150 VTAIL.n116 8.2187
R1388 VTAIL.n36 VTAIL.n2 8.2187
R1389 VTAIL.n114 VTAIL.n80 8.2187
R1390 VTAIL.n76 VTAIL.n42 8.2187
R1391 VTAIL.n132 VTAIL.n131 8.14595
R1392 VTAIL.n18 VTAIL.n17 8.14595
R1393 VTAIL.n96 VTAIL.n95 8.14595
R1394 VTAIL.n58 VTAIL.n57 8.14595
R1395 VTAIL.n128 VTAIL.n126 7.3702
R1396 VTAIL.n14 VTAIL.n12 7.3702
R1397 VTAIL.n92 VTAIL.n90 7.3702
R1398 VTAIL.n54 VTAIL.n52 7.3702
R1399 VTAIL.n131 VTAIL.n126 5.81868
R1400 VTAIL.n17 VTAIL.n12 5.81868
R1401 VTAIL.n95 VTAIL.n90 5.81868
R1402 VTAIL.n57 VTAIL.n52 5.81868
R1403 VTAIL.n148 VTAIL.n116 5.3904
R1404 VTAIL.n34 VTAIL.n2 5.3904
R1405 VTAIL.n112 VTAIL.n80 5.3904
R1406 VTAIL.n74 VTAIL.n42 5.3904
R1407 VTAIL.n132 VTAIL.n124 5.04292
R1408 VTAIL.n18 VTAIL.n10 5.04292
R1409 VTAIL.n96 VTAIL.n88 5.04292
R1410 VTAIL.n58 VTAIL.n50 5.04292
R1411 VTAIL.n136 VTAIL.n135 4.26717
R1412 VTAIL.n22 VTAIL.n21 4.26717
R1413 VTAIL.n100 VTAIL.n99 4.26717
R1414 VTAIL.n62 VTAIL.n61 4.26717
R1415 VTAIL.n139 VTAIL.n122 3.49141
R1416 VTAIL.n25 VTAIL.n8 3.49141
R1417 VTAIL.n103 VTAIL.n86 3.49141
R1418 VTAIL.n65 VTAIL.n48 3.49141
R1419 VTAIL.n127 VTAIL.n125 2.84305
R1420 VTAIL.n13 VTAIL.n11 2.84305
R1421 VTAIL.n91 VTAIL.n89 2.84305
R1422 VTAIL.n53 VTAIL.n51 2.84305
R1423 VTAIL.n0 VTAIL.t11 2.73153
R1424 VTAIL.n0 VTAIL.t9 2.73153
R1425 VTAIL.n38 VTAIL.t0 2.73153
R1426 VTAIL.n38 VTAIL.t5 2.73153
R1427 VTAIL.n78 VTAIL.t1 2.73153
R1428 VTAIL.n78 VTAIL.t2 2.73153
R1429 VTAIL.n40 VTAIL.t7 2.73153
R1430 VTAIL.n40 VTAIL.t6 2.73153
R1431 VTAIL.n140 VTAIL.n120 2.71565
R1432 VTAIL.n26 VTAIL.n6 2.71565
R1433 VTAIL.n104 VTAIL.n84 2.71565
R1434 VTAIL.n66 VTAIL.n46 2.71565
R1435 VTAIL.n77 VTAIL.n41 2.00912
R1436 VTAIL.n115 VTAIL.n79 2.00912
R1437 VTAIL.n39 VTAIL.n37 2.00912
R1438 VTAIL.n144 VTAIL.n143 1.93989
R1439 VTAIL.n30 VTAIL.n29 1.93989
R1440 VTAIL.n108 VTAIL.n107 1.93989
R1441 VTAIL.n70 VTAIL.n69 1.93989
R1442 VTAIL.n79 VTAIL.n77 1.47464
R1443 VTAIL.n37 VTAIL.n1 1.47464
R1444 VTAIL VTAIL.n151 1.44878
R1445 VTAIL.n147 VTAIL.n118 1.16414
R1446 VTAIL.n33 VTAIL.n4 1.16414
R1447 VTAIL.n111 VTAIL.n82 1.16414
R1448 VTAIL.n73 VTAIL.n44 1.16414
R1449 VTAIL VTAIL.n1 0.560845
R1450 VTAIL.n133 VTAIL.n125 0.155672
R1451 VTAIL.n134 VTAIL.n133 0.155672
R1452 VTAIL.n134 VTAIL.n121 0.155672
R1453 VTAIL.n141 VTAIL.n121 0.155672
R1454 VTAIL.n142 VTAIL.n141 0.155672
R1455 VTAIL.n142 VTAIL.n117 0.155672
R1456 VTAIL.n149 VTAIL.n117 0.155672
R1457 VTAIL.n19 VTAIL.n11 0.155672
R1458 VTAIL.n20 VTAIL.n19 0.155672
R1459 VTAIL.n20 VTAIL.n7 0.155672
R1460 VTAIL.n27 VTAIL.n7 0.155672
R1461 VTAIL.n28 VTAIL.n27 0.155672
R1462 VTAIL.n28 VTAIL.n3 0.155672
R1463 VTAIL.n35 VTAIL.n3 0.155672
R1464 VTAIL.n113 VTAIL.n81 0.155672
R1465 VTAIL.n106 VTAIL.n81 0.155672
R1466 VTAIL.n106 VTAIL.n105 0.155672
R1467 VTAIL.n105 VTAIL.n85 0.155672
R1468 VTAIL.n98 VTAIL.n85 0.155672
R1469 VTAIL.n98 VTAIL.n97 0.155672
R1470 VTAIL.n97 VTAIL.n89 0.155672
R1471 VTAIL.n75 VTAIL.n43 0.155672
R1472 VTAIL.n68 VTAIL.n43 0.155672
R1473 VTAIL.n68 VTAIL.n67 0.155672
R1474 VTAIL.n67 VTAIL.n47 0.155672
R1475 VTAIL.n60 VTAIL.n47 0.155672
R1476 VTAIL.n60 VTAIL.n59 0.155672
R1477 VTAIL.n59 VTAIL.n51 0.155672
R1478 VDD2.n67 VDD2.n37 214.453
R1479 VDD2.n30 VDD2.n0 214.453
R1480 VDD2.n68 VDD2.n67 185
R1481 VDD2.n66 VDD2.n65 185
R1482 VDD2.n41 VDD2.n40 185
R1483 VDD2.n60 VDD2.n59 185
R1484 VDD2.n58 VDD2.n57 185
R1485 VDD2.n45 VDD2.n44 185
R1486 VDD2.n52 VDD2.n51 185
R1487 VDD2.n50 VDD2.n49 185
R1488 VDD2.n13 VDD2.n12 185
R1489 VDD2.n15 VDD2.n14 185
R1490 VDD2.n8 VDD2.n7 185
R1491 VDD2.n21 VDD2.n20 185
R1492 VDD2.n23 VDD2.n22 185
R1493 VDD2.n4 VDD2.n3 185
R1494 VDD2.n29 VDD2.n28 185
R1495 VDD2.n31 VDD2.n30 185
R1496 VDD2.n11 VDD2.t5 149.524
R1497 VDD2.n48 VDD2.t3 149.524
R1498 VDD2.n67 VDD2.n66 104.615
R1499 VDD2.n66 VDD2.n40 104.615
R1500 VDD2.n59 VDD2.n40 104.615
R1501 VDD2.n59 VDD2.n58 104.615
R1502 VDD2.n58 VDD2.n44 104.615
R1503 VDD2.n51 VDD2.n44 104.615
R1504 VDD2.n51 VDD2.n50 104.615
R1505 VDD2.n14 VDD2.n13 104.615
R1506 VDD2.n14 VDD2.n7 104.615
R1507 VDD2.n21 VDD2.n7 104.615
R1508 VDD2.n22 VDD2.n21 104.615
R1509 VDD2.n22 VDD2.n3 104.615
R1510 VDD2.n29 VDD2.n3 104.615
R1511 VDD2.n30 VDD2.n29 104.615
R1512 VDD2.n36 VDD2.n35 68.3786
R1513 VDD2 VDD2.n73 68.3757
R1514 VDD2.n36 VDD2.n34 53.6122
R1515 VDD2.n50 VDD2.t3 52.3082
R1516 VDD2.n13 VDD2.t5 52.3082
R1517 VDD2.n72 VDD2.n71 52.1611
R1518 VDD2.n72 VDD2.n36 36.4933
R1519 VDD2.n69 VDD2.n68 12.8005
R1520 VDD2.n32 VDD2.n31 12.8005
R1521 VDD2.n65 VDD2.n39 12.0247
R1522 VDD2.n28 VDD2.n2 12.0247
R1523 VDD2.n64 VDD2.n41 11.249
R1524 VDD2.n27 VDD2.n4 11.249
R1525 VDD2.n61 VDD2.n60 10.4732
R1526 VDD2.n24 VDD2.n23 10.4732
R1527 VDD2.n49 VDD2.n48 10.2747
R1528 VDD2.n12 VDD2.n11 10.2747
R1529 VDD2.n57 VDD2.n43 9.69747
R1530 VDD2.n20 VDD2.n6 9.69747
R1531 VDD2.n71 VDD2.n70 9.45567
R1532 VDD2.n34 VDD2.n33 9.45567
R1533 VDD2.n47 VDD2.n46 9.3005
R1534 VDD2.n54 VDD2.n53 9.3005
R1535 VDD2.n56 VDD2.n55 9.3005
R1536 VDD2.n43 VDD2.n42 9.3005
R1537 VDD2.n62 VDD2.n61 9.3005
R1538 VDD2.n64 VDD2.n63 9.3005
R1539 VDD2.n39 VDD2.n38 9.3005
R1540 VDD2.n70 VDD2.n69 9.3005
R1541 VDD2.n10 VDD2.n9 9.3005
R1542 VDD2.n17 VDD2.n16 9.3005
R1543 VDD2.n19 VDD2.n18 9.3005
R1544 VDD2.n6 VDD2.n5 9.3005
R1545 VDD2.n25 VDD2.n24 9.3005
R1546 VDD2.n27 VDD2.n26 9.3005
R1547 VDD2.n2 VDD2.n1 9.3005
R1548 VDD2.n33 VDD2.n32 9.3005
R1549 VDD2.n56 VDD2.n45 8.92171
R1550 VDD2.n19 VDD2.n8 8.92171
R1551 VDD2.n71 VDD2.n37 8.2187
R1552 VDD2.n34 VDD2.n0 8.2187
R1553 VDD2.n53 VDD2.n52 8.14595
R1554 VDD2.n16 VDD2.n15 8.14595
R1555 VDD2.n49 VDD2.n47 7.3702
R1556 VDD2.n12 VDD2.n10 7.3702
R1557 VDD2.n52 VDD2.n47 5.81868
R1558 VDD2.n15 VDD2.n10 5.81868
R1559 VDD2.n69 VDD2.n37 5.3904
R1560 VDD2.n32 VDD2.n0 5.3904
R1561 VDD2.n53 VDD2.n45 5.04292
R1562 VDD2.n16 VDD2.n8 5.04292
R1563 VDD2.n57 VDD2.n56 4.26717
R1564 VDD2.n20 VDD2.n19 4.26717
R1565 VDD2.n60 VDD2.n43 3.49141
R1566 VDD2.n23 VDD2.n6 3.49141
R1567 VDD2.n48 VDD2.n46 2.84305
R1568 VDD2.n11 VDD2.n9 2.84305
R1569 VDD2.n73 VDD2.t4 2.73153
R1570 VDD2.n73 VDD2.t2 2.73153
R1571 VDD2.n35 VDD2.t1 2.73153
R1572 VDD2.n35 VDD2.t0 2.73153
R1573 VDD2.n61 VDD2.n41 2.71565
R1574 VDD2.n24 VDD2.n4 2.71565
R1575 VDD2.n65 VDD2.n64 1.93989
R1576 VDD2.n28 VDD2.n27 1.93989
R1577 VDD2 VDD2.n72 1.56516
R1578 VDD2.n68 VDD2.n39 1.16414
R1579 VDD2.n31 VDD2.n2 1.16414
R1580 VDD2.n70 VDD2.n38 0.155672
R1581 VDD2.n63 VDD2.n38 0.155672
R1582 VDD2.n63 VDD2.n62 0.155672
R1583 VDD2.n62 VDD2.n42 0.155672
R1584 VDD2.n55 VDD2.n42 0.155672
R1585 VDD2.n55 VDD2.n54 0.155672
R1586 VDD2.n54 VDD2.n46 0.155672
R1587 VDD2.n17 VDD2.n9 0.155672
R1588 VDD2.n18 VDD2.n17 0.155672
R1589 VDD2.n18 VDD2.n5 0.155672
R1590 VDD2.n25 VDD2.n5 0.155672
R1591 VDD2.n26 VDD2.n25 0.155672
R1592 VDD2.n26 VDD2.n1 0.155672
R1593 VDD2.n33 VDD2.n1 0.155672
R1594 VP.n10 VP.n9 161.3
R1595 VP.n11 VP.n6 161.3
R1596 VP.n13 VP.n12 161.3
R1597 VP.n14 VP.n5 161.3
R1598 VP.n31 VP.n0 161.3
R1599 VP.n30 VP.n29 161.3
R1600 VP.n28 VP.n1 161.3
R1601 VP.n27 VP.n26 161.3
R1602 VP.n25 VP.n2 161.3
R1603 VP.n24 VP.n23 161.3
R1604 VP.n22 VP.n3 161.3
R1605 VP.n21 VP.n20 161.3
R1606 VP.n19 VP.n4 161.3
R1607 VP.n7 VP.t2 120.799
R1608 VP.n18 VP.n17 94.6082
R1609 VP.n33 VP.n32 94.6082
R1610 VP.n16 VP.n15 94.6082
R1611 VP.n25 VP.t5 87.363
R1612 VP.n18 VP.t3 87.363
R1613 VP.n32 VP.t1 87.363
R1614 VP.n15 VP.t0 87.363
R1615 VP.n8 VP.t4 87.363
R1616 VP.n20 VP.n3 56.5193
R1617 VP.n30 VP.n1 56.5193
R1618 VP.n13 VP.n6 56.5193
R1619 VP.n8 VP.n7 45.7103
R1620 VP.n17 VP.n16 42.6928
R1621 VP.n20 VP.n19 24.4675
R1622 VP.n24 VP.n3 24.4675
R1623 VP.n25 VP.n24 24.4675
R1624 VP.n26 VP.n25 24.4675
R1625 VP.n26 VP.n1 24.4675
R1626 VP.n31 VP.n30 24.4675
R1627 VP.n14 VP.n13 24.4675
R1628 VP.n9 VP.n8 24.4675
R1629 VP.n9 VP.n6 24.4675
R1630 VP.n19 VP.n18 16.1487
R1631 VP.n32 VP.n31 16.1487
R1632 VP.n15 VP.n14 16.1487
R1633 VP.n10 VP.n7 9.33007
R1634 VP.n16 VP.n5 0.278367
R1635 VP.n17 VP.n4 0.278367
R1636 VP.n33 VP.n0 0.278367
R1637 VP.n11 VP.n10 0.189894
R1638 VP.n12 VP.n11 0.189894
R1639 VP.n12 VP.n5 0.189894
R1640 VP.n21 VP.n4 0.189894
R1641 VP.n22 VP.n21 0.189894
R1642 VP.n23 VP.n22 0.189894
R1643 VP.n23 VP.n2 0.189894
R1644 VP.n27 VP.n2 0.189894
R1645 VP.n28 VP.n27 0.189894
R1646 VP.n29 VP.n28 0.189894
R1647 VP.n29 VP.n0 0.189894
R1648 VP VP.n33 0.153454
R1649 VDD1.n30 VDD1.n0 214.453
R1650 VDD1.n65 VDD1.n35 214.453
R1651 VDD1.n31 VDD1.n30 185
R1652 VDD1.n29 VDD1.n28 185
R1653 VDD1.n4 VDD1.n3 185
R1654 VDD1.n23 VDD1.n22 185
R1655 VDD1.n21 VDD1.n20 185
R1656 VDD1.n8 VDD1.n7 185
R1657 VDD1.n15 VDD1.n14 185
R1658 VDD1.n13 VDD1.n12 185
R1659 VDD1.n48 VDD1.n47 185
R1660 VDD1.n50 VDD1.n49 185
R1661 VDD1.n43 VDD1.n42 185
R1662 VDD1.n56 VDD1.n55 185
R1663 VDD1.n58 VDD1.n57 185
R1664 VDD1.n39 VDD1.n38 185
R1665 VDD1.n64 VDD1.n63 185
R1666 VDD1.n66 VDD1.n65 185
R1667 VDD1.n46 VDD1.t2 149.524
R1668 VDD1.n11 VDD1.t3 149.524
R1669 VDD1.n30 VDD1.n29 104.615
R1670 VDD1.n29 VDD1.n3 104.615
R1671 VDD1.n22 VDD1.n3 104.615
R1672 VDD1.n22 VDD1.n21 104.615
R1673 VDD1.n21 VDD1.n7 104.615
R1674 VDD1.n14 VDD1.n7 104.615
R1675 VDD1.n14 VDD1.n13 104.615
R1676 VDD1.n49 VDD1.n48 104.615
R1677 VDD1.n49 VDD1.n42 104.615
R1678 VDD1.n56 VDD1.n42 104.615
R1679 VDD1.n57 VDD1.n56 104.615
R1680 VDD1.n57 VDD1.n38 104.615
R1681 VDD1.n64 VDD1.n38 104.615
R1682 VDD1.n65 VDD1.n64 104.615
R1683 VDD1.n71 VDD1.n70 68.3786
R1684 VDD1.n73 VDD1.n72 67.9318
R1685 VDD1 VDD1.n34 53.7258
R1686 VDD1.n71 VDD1.n69 53.6122
R1687 VDD1.n13 VDD1.t3 52.3082
R1688 VDD1.n48 VDD1.t2 52.3082
R1689 VDD1.n73 VDD1.n71 38.0806
R1690 VDD1.n32 VDD1.n31 12.8005
R1691 VDD1.n67 VDD1.n66 12.8005
R1692 VDD1.n28 VDD1.n2 12.0247
R1693 VDD1.n63 VDD1.n37 12.0247
R1694 VDD1.n27 VDD1.n4 11.249
R1695 VDD1.n62 VDD1.n39 11.249
R1696 VDD1.n24 VDD1.n23 10.4732
R1697 VDD1.n59 VDD1.n58 10.4732
R1698 VDD1.n12 VDD1.n11 10.2747
R1699 VDD1.n47 VDD1.n46 10.2747
R1700 VDD1.n20 VDD1.n6 9.69747
R1701 VDD1.n55 VDD1.n41 9.69747
R1702 VDD1.n34 VDD1.n33 9.45567
R1703 VDD1.n69 VDD1.n68 9.45567
R1704 VDD1.n10 VDD1.n9 9.3005
R1705 VDD1.n17 VDD1.n16 9.3005
R1706 VDD1.n19 VDD1.n18 9.3005
R1707 VDD1.n6 VDD1.n5 9.3005
R1708 VDD1.n25 VDD1.n24 9.3005
R1709 VDD1.n27 VDD1.n26 9.3005
R1710 VDD1.n2 VDD1.n1 9.3005
R1711 VDD1.n33 VDD1.n32 9.3005
R1712 VDD1.n45 VDD1.n44 9.3005
R1713 VDD1.n52 VDD1.n51 9.3005
R1714 VDD1.n54 VDD1.n53 9.3005
R1715 VDD1.n41 VDD1.n40 9.3005
R1716 VDD1.n60 VDD1.n59 9.3005
R1717 VDD1.n62 VDD1.n61 9.3005
R1718 VDD1.n37 VDD1.n36 9.3005
R1719 VDD1.n68 VDD1.n67 9.3005
R1720 VDD1.n19 VDD1.n8 8.92171
R1721 VDD1.n54 VDD1.n43 8.92171
R1722 VDD1.n34 VDD1.n0 8.2187
R1723 VDD1.n69 VDD1.n35 8.2187
R1724 VDD1.n16 VDD1.n15 8.14595
R1725 VDD1.n51 VDD1.n50 8.14595
R1726 VDD1.n12 VDD1.n10 7.3702
R1727 VDD1.n47 VDD1.n45 7.3702
R1728 VDD1.n15 VDD1.n10 5.81868
R1729 VDD1.n50 VDD1.n45 5.81868
R1730 VDD1.n32 VDD1.n0 5.3904
R1731 VDD1.n67 VDD1.n35 5.3904
R1732 VDD1.n16 VDD1.n8 5.04292
R1733 VDD1.n51 VDD1.n43 5.04292
R1734 VDD1.n20 VDD1.n19 4.26717
R1735 VDD1.n55 VDD1.n54 4.26717
R1736 VDD1.n23 VDD1.n6 3.49141
R1737 VDD1.n58 VDD1.n41 3.49141
R1738 VDD1.n11 VDD1.n9 2.84305
R1739 VDD1.n46 VDD1.n44 2.84305
R1740 VDD1.n72 VDD1.t1 2.73153
R1741 VDD1.n72 VDD1.t5 2.73153
R1742 VDD1.n70 VDD1.t0 2.73153
R1743 VDD1.n70 VDD1.t4 2.73153
R1744 VDD1.n24 VDD1.n4 2.71565
R1745 VDD1.n59 VDD1.n39 2.71565
R1746 VDD1.n28 VDD1.n27 1.93989
R1747 VDD1.n63 VDD1.n62 1.93989
R1748 VDD1.n31 VDD1.n2 1.16414
R1749 VDD1.n66 VDD1.n37 1.16414
R1750 VDD1 VDD1.n73 0.444466
R1751 VDD1.n33 VDD1.n1 0.155672
R1752 VDD1.n26 VDD1.n1 0.155672
R1753 VDD1.n26 VDD1.n25 0.155672
R1754 VDD1.n25 VDD1.n5 0.155672
R1755 VDD1.n18 VDD1.n5 0.155672
R1756 VDD1.n18 VDD1.n17 0.155672
R1757 VDD1.n17 VDD1.n9 0.155672
R1758 VDD1.n52 VDD1.n44 0.155672
R1759 VDD1.n53 VDD1.n52 0.155672
R1760 VDD1.n53 VDD1.n40 0.155672
R1761 VDD1.n60 VDD1.n40 0.155672
R1762 VDD1.n61 VDD1.n60 0.155672
R1763 VDD1.n61 VDD1.n36 0.155672
R1764 VDD1.n68 VDD1.n36 0.155672
C0 VDD1 VDD2 1.18465f
C1 VN VTAIL 4.20881f
C2 VTAIL VP 4.22306f
C3 VN VP 5.46816f
C4 VDD1 VTAIL 5.81731f
C5 VDD1 VN 0.149983f
C6 VDD1 VP 4.23827f
C7 VDD2 VTAIL 5.86475f
C8 VDD2 VN 3.98356f
C9 VDD2 VP 0.407102f
C10 VDD2 B 4.668662f
C11 VDD1 B 4.769878f
C12 VTAIL B 5.537355f
C13 VN B 10.76734f
C14 VP B 9.383179f
C15 VDD1.n0 B 0.030235f
C16 VDD1.n1 B 0.021922f
C17 VDD1.n2 B 0.01178f
C18 VDD1.n3 B 0.027844f
C19 VDD1.n4 B 0.012473f
C20 VDD1.n5 B 0.021922f
C21 VDD1.n6 B 0.01178f
C22 VDD1.n7 B 0.027844f
C23 VDD1.n8 B 0.012473f
C24 VDD1.n9 B 0.6427f
C25 VDD1.n10 B 0.01178f
C26 VDD1.t3 B 0.046497f
C27 VDD1.n11 B 0.118135f
C28 VDD1.n12 B 0.019684f
C29 VDD1.n13 B 0.020883f
C30 VDD1.n14 B 0.027844f
C31 VDD1.n15 B 0.012473f
C32 VDD1.n16 B 0.01178f
C33 VDD1.n17 B 0.021922f
C34 VDD1.n18 B 0.021922f
C35 VDD1.n19 B 0.01178f
C36 VDD1.n20 B 0.012473f
C37 VDD1.n21 B 0.027844f
C38 VDD1.n22 B 0.027844f
C39 VDD1.n23 B 0.012473f
C40 VDD1.n24 B 0.01178f
C41 VDD1.n25 B 0.021922f
C42 VDD1.n26 B 0.021922f
C43 VDD1.n27 B 0.01178f
C44 VDD1.n28 B 0.012473f
C45 VDD1.n29 B 0.027844f
C46 VDD1.n30 B 0.057243f
C47 VDD1.n31 B 0.012473f
C48 VDD1.n32 B 0.023034f
C49 VDD1.n33 B 0.055764f
C50 VDD1.n34 B 0.079085f
C51 VDD1.n35 B 0.030235f
C52 VDD1.n36 B 0.021922f
C53 VDD1.n37 B 0.01178f
C54 VDD1.n38 B 0.027844f
C55 VDD1.n39 B 0.012473f
C56 VDD1.n40 B 0.021922f
C57 VDD1.n41 B 0.01178f
C58 VDD1.n42 B 0.027844f
C59 VDD1.n43 B 0.012473f
C60 VDD1.n44 B 0.6427f
C61 VDD1.n45 B 0.01178f
C62 VDD1.t2 B 0.046497f
C63 VDD1.n46 B 0.118135f
C64 VDD1.n47 B 0.019684f
C65 VDD1.n48 B 0.020883f
C66 VDD1.n49 B 0.027844f
C67 VDD1.n50 B 0.012473f
C68 VDD1.n51 B 0.01178f
C69 VDD1.n52 B 0.021922f
C70 VDD1.n53 B 0.021922f
C71 VDD1.n54 B 0.01178f
C72 VDD1.n55 B 0.012473f
C73 VDD1.n56 B 0.027844f
C74 VDD1.n57 B 0.027844f
C75 VDD1.n58 B 0.012473f
C76 VDD1.n59 B 0.01178f
C77 VDD1.n60 B 0.021922f
C78 VDD1.n61 B 0.021922f
C79 VDD1.n62 B 0.01178f
C80 VDD1.n63 B 0.012473f
C81 VDD1.n64 B 0.027844f
C82 VDD1.n65 B 0.057243f
C83 VDD1.n66 B 0.012473f
C84 VDD1.n67 B 0.023034f
C85 VDD1.n68 B 0.055764f
C86 VDD1.n69 B 0.078558f
C87 VDD1.t0 B 0.125597f
C88 VDD1.t4 B 0.125597f
C89 VDD1.n70 B 1.08126f
C90 VDD1.n71 B 1.95559f
C91 VDD1.t1 B 0.125597f
C92 VDD1.t5 B 0.125597f
C93 VDD1.n72 B 1.07894f
C94 VDD1.n73 B 1.96608f
C95 VP.n0 B 0.039034f
C96 VP.t1 B 1.1478f
C97 VP.n1 B 0.036211f
C98 VP.n2 B 0.029607f
C99 VP.t5 B 1.1478f
C100 VP.n3 B 0.036211f
C101 VP.n4 B 0.039034f
C102 VP.t3 B 1.1478f
C103 VP.n5 B 0.039034f
C104 VP.t0 B 1.1478f
C105 VP.n6 B 0.036211f
C106 VP.t2 B 1.30799f
C107 VP.n7 B 0.491713f
C108 VP.t4 B 1.1478f
C109 VP.n8 B 0.514578f
C110 VP.n9 B 0.05518f
C111 VP.n10 B 0.246441f
C112 VP.n11 B 0.029607f
C113 VP.n12 B 0.029607f
C114 VP.n13 B 0.050237f
C115 VP.n14 B 0.045918f
C116 VP.n15 B 0.512813f
C117 VP.n16 B 1.28262f
C118 VP.n17 B 1.30755f
C119 VP.n18 B 0.512813f
C120 VP.n19 B 0.045918f
C121 VP.n20 B 0.050237f
C122 VP.n21 B 0.029607f
C123 VP.n22 B 0.029607f
C124 VP.n23 B 0.029607f
C125 VP.n24 B 0.05518f
C126 VP.n25 B 0.456218f
C127 VP.n26 B 0.05518f
C128 VP.n27 B 0.029607f
C129 VP.n28 B 0.029607f
C130 VP.n29 B 0.029607f
C131 VP.n30 B 0.050237f
C132 VP.n31 B 0.045918f
C133 VP.n32 B 0.512813f
C134 VP.n33 B 0.038814f
C135 VDD2.n0 B 0.030177f
C136 VDD2.n1 B 0.02188f
C137 VDD2.n2 B 0.011758f
C138 VDD2.n3 B 0.027791f
C139 VDD2.n4 B 0.012449f
C140 VDD2.n5 B 0.02188f
C141 VDD2.n6 B 0.011758f
C142 VDD2.n7 B 0.027791f
C143 VDD2.n8 B 0.012449f
C144 VDD2.n9 B 0.641467f
C145 VDD2.n10 B 0.011758f
C146 VDD2.t5 B 0.046408f
C147 VDD2.n11 B 0.117908f
C148 VDD2.n12 B 0.019646f
C149 VDD2.n13 B 0.020843f
C150 VDD2.n14 B 0.027791f
C151 VDD2.n15 B 0.012449f
C152 VDD2.n16 B 0.011758f
C153 VDD2.n17 B 0.02188f
C154 VDD2.n18 B 0.02188f
C155 VDD2.n19 B 0.011758f
C156 VDD2.n20 B 0.012449f
C157 VDD2.n21 B 0.027791f
C158 VDD2.n22 B 0.027791f
C159 VDD2.n23 B 0.012449f
C160 VDD2.n24 B 0.011758f
C161 VDD2.n25 B 0.02188f
C162 VDD2.n26 B 0.02188f
C163 VDD2.n27 B 0.011758f
C164 VDD2.n28 B 0.012449f
C165 VDD2.n29 B 0.027791f
C166 VDD2.n30 B 0.057133f
C167 VDD2.n31 B 0.012449f
C168 VDD2.n32 B 0.02299f
C169 VDD2.n33 B 0.055657f
C170 VDD2.n34 B 0.078407f
C171 VDD2.t1 B 0.125356f
C172 VDD2.t0 B 0.125356f
C173 VDD2.n35 B 1.07918f
C174 VDD2.n36 B 1.85989f
C175 VDD2.n37 B 0.030177f
C176 VDD2.n38 B 0.02188f
C177 VDD2.n39 B 0.011758f
C178 VDD2.n40 B 0.027791f
C179 VDD2.n41 B 0.012449f
C180 VDD2.n42 B 0.02188f
C181 VDD2.n43 B 0.011758f
C182 VDD2.n44 B 0.027791f
C183 VDD2.n45 B 0.012449f
C184 VDD2.n46 B 0.641467f
C185 VDD2.n47 B 0.011758f
C186 VDD2.t3 B 0.046408f
C187 VDD2.n48 B 0.117908f
C188 VDD2.n49 B 0.019646f
C189 VDD2.n50 B 0.020843f
C190 VDD2.n51 B 0.027791f
C191 VDD2.n52 B 0.012449f
C192 VDD2.n53 B 0.011758f
C193 VDD2.n54 B 0.02188f
C194 VDD2.n55 B 0.02188f
C195 VDD2.n56 B 0.011758f
C196 VDD2.n57 B 0.012449f
C197 VDD2.n58 B 0.027791f
C198 VDD2.n59 B 0.027791f
C199 VDD2.n60 B 0.012449f
C200 VDD2.n61 B 0.011758f
C201 VDD2.n62 B 0.02188f
C202 VDD2.n63 B 0.02188f
C203 VDD2.n64 B 0.011758f
C204 VDD2.n65 B 0.012449f
C205 VDD2.n66 B 0.027791f
C206 VDD2.n67 B 0.057133f
C207 VDD2.n68 B 0.012449f
C208 VDD2.n69 B 0.02299f
C209 VDD2.n70 B 0.055657f
C210 VDD2.n71 B 0.074409f
C211 VDD2.n72 B 1.77547f
C212 VDD2.t4 B 0.125356f
C213 VDD2.t2 B 0.125356f
C214 VDD2.n73 B 1.07916f
C215 VTAIL.t11 B 0.144229f
C216 VTAIL.t9 B 0.144229f
C217 VTAIL.n0 B 1.1763f
C218 VTAIL.n1 B 0.390928f
C219 VTAIL.n2 B 0.03472f
C220 VTAIL.n3 B 0.025174f
C221 VTAIL.n4 B 0.013528f
C222 VTAIL.n5 B 0.031974f
C223 VTAIL.n6 B 0.014323f
C224 VTAIL.n7 B 0.025174f
C225 VTAIL.n8 B 0.013528f
C226 VTAIL.n9 B 0.031974f
C227 VTAIL.n10 B 0.014323f
C228 VTAIL.n11 B 0.738039f
C229 VTAIL.n12 B 0.013528f
C230 VTAIL.t4 B 0.053395f
C231 VTAIL.n13 B 0.135659f
C232 VTAIL.n14 B 0.022603f
C233 VTAIL.n15 B 0.023981f
C234 VTAIL.n16 B 0.031974f
C235 VTAIL.n17 B 0.014323f
C236 VTAIL.n18 B 0.013528f
C237 VTAIL.n19 B 0.025174f
C238 VTAIL.n20 B 0.025174f
C239 VTAIL.n21 B 0.013528f
C240 VTAIL.n22 B 0.014323f
C241 VTAIL.n23 B 0.031974f
C242 VTAIL.n24 B 0.031974f
C243 VTAIL.n25 B 0.014323f
C244 VTAIL.n26 B 0.013528f
C245 VTAIL.n27 B 0.025174f
C246 VTAIL.n28 B 0.025174f
C247 VTAIL.n29 B 0.013528f
C248 VTAIL.n30 B 0.014323f
C249 VTAIL.n31 B 0.031974f
C250 VTAIL.n32 B 0.065735f
C251 VTAIL.n33 B 0.014323f
C252 VTAIL.n34 B 0.026451f
C253 VTAIL.n35 B 0.064036f
C254 VTAIL.n36 B 0.06827f
C255 VTAIL.n37 B 0.307321f
C256 VTAIL.t0 B 0.144229f
C257 VTAIL.t5 B 0.144229f
C258 VTAIL.n38 B 1.1763f
C259 VTAIL.n39 B 1.56365f
C260 VTAIL.t7 B 0.144229f
C261 VTAIL.t6 B 0.144229f
C262 VTAIL.n40 B 1.17631f
C263 VTAIL.n41 B 1.56364f
C264 VTAIL.n42 B 0.03472f
C265 VTAIL.n43 B 0.025174f
C266 VTAIL.n44 B 0.013528f
C267 VTAIL.n45 B 0.031974f
C268 VTAIL.n46 B 0.014323f
C269 VTAIL.n47 B 0.025174f
C270 VTAIL.n48 B 0.013528f
C271 VTAIL.n49 B 0.031974f
C272 VTAIL.n50 B 0.014323f
C273 VTAIL.n51 B 0.738039f
C274 VTAIL.n52 B 0.013528f
C275 VTAIL.t8 B 0.053395f
C276 VTAIL.n53 B 0.135659f
C277 VTAIL.n54 B 0.022603f
C278 VTAIL.n55 B 0.023981f
C279 VTAIL.n56 B 0.031974f
C280 VTAIL.n57 B 0.014323f
C281 VTAIL.n58 B 0.013528f
C282 VTAIL.n59 B 0.025174f
C283 VTAIL.n60 B 0.025174f
C284 VTAIL.n61 B 0.013528f
C285 VTAIL.n62 B 0.014323f
C286 VTAIL.n63 B 0.031974f
C287 VTAIL.n64 B 0.031974f
C288 VTAIL.n65 B 0.014323f
C289 VTAIL.n66 B 0.013528f
C290 VTAIL.n67 B 0.025174f
C291 VTAIL.n68 B 0.025174f
C292 VTAIL.n69 B 0.013528f
C293 VTAIL.n70 B 0.014323f
C294 VTAIL.n71 B 0.031974f
C295 VTAIL.n72 B 0.065735f
C296 VTAIL.n73 B 0.014323f
C297 VTAIL.n74 B 0.026451f
C298 VTAIL.n75 B 0.064036f
C299 VTAIL.n76 B 0.06827f
C300 VTAIL.n77 B 0.307321f
C301 VTAIL.t1 B 0.144229f
C302 VTAIL.t2 B 0.144229f
C303 VTAIL.n78 B 1.17631f
C304 VTAIL.n79 B 0.508401f
C305 VTAIL.n80 B 0.03472f
C306 VTAIL.n81 B 0.025174f
C307 VTAIL.n82 B 0.013528f
C308 VTAIL.n83 B 0.031974f
C309 VTAIL.n84 B 0.014323f
C310 VTAIL.n85 B 0.025174f
C311 VTAIL.n86 B 0.013528f
C312 VTAIL.n87 B 0.031974f
C313 VTAIL.n88 B 0.014323f
C314 VTAIL.n89 B 0.738039f
C315 VTAIL.n90 B 0.013528f
C316 VTAIL.t3 B 0.053395f
C317 VTAIL.n91 B 0.135659f
C318 VTAIL.n92 B 0.022603f
C319 VTAIL.n93 B 0.023981f
C320 VTAIL.n94 B 0.031974f
C321 VTAIL.n95 B 0.014323f
C322 VTAIL.n96 B 0.013528f
C323 VTAIL.n97 B 0.025174f
C324 VTAIL.n98 B 0.025174f
C325 VTAIL.n99 B 0.013528f
C326 VTAIL.n100 B 0.014323f
C327 VTAIL.n101 B 0.031974f
C328 VTAIL.n102 B 0.031974f
C329 VTAIL.n103 B 0.014323f
C330 VTAIL.n104 B 0.013528f
C331 VTAIL.n105 B 0.025174f
C332 VTAIL.n106 B 0.025174f
C333 VTAIL.n107 B 0.013528f
C334 VTAIL.n108 B 0.014323f
C335 VTAIL.n109 B 0.031974f
C336 VTAIL.n110 B 0.065735f
C337 VTAIL.n111 B 0.014323f
C338 VTAIL.n112 B 0.026451f
C339 VTAIL.n113 B 0.064036f
C340 VTAIL.n114 B 0.06827f
C341 VTAIL.n115 B 1.19963f
C342 VTAIL.n116 B 0.03472f
C343 VTAIL.n117 B 0.025174f
C344 VTAIL.n118 B 0.013528f
C345 VTAIL.n119 B 0.031974f
C346 VTAIL.n120 B 0.014323f
C347 VTAIL.n121 B 0.025174f
C348 VTAIL.n122 B 0.013528f
C349 VTAIL.n123 B 0.031974f
C350 VTAIL.n124 B 0.014323f
C351 VTAIL.n125 B 0.738039f
C352 VTAIL.n126 B 0.013528f
C353 VTAIL.t10 B 0.053395f
C354 VTAIL.n127 B 0.135659f
C355 VTAIL.n128 B 0.022603f
C356 VTAIL.n129 B 0.023981f
C357 VTAIL.n130 B 0.031974f
C358 VTAIL.n131 B 0.014323f
C359 VTAIL.n132 B 0.013528f
C360 VTAIL.n133 B 0.025174f
C361 VTAIL.n134 B 0.025174f
C362 VTAIL.n135 B 0.013528f
C363 VTAIL.n136 B 0.014323f
C364 VTAIL.n137 B 0.031974f
C365 VTAIL.n138 B 0.031974f
C366 VTAIL.n139 B 0.014323f
C367 VTAIL.n140 B 0.013528f
C368 VTAIL.n141 B 0.025174f
C369 VTAIL.n142 B 0.025174f
C370 VTAIL.n143 B 0.013528f
C371 VTAIL.n144 B 0.014323f
C372 VTAIL.n145 B 0.031974f
C373 VTAIL.n146 B 0.065735f
C374 VTAIL.n147 B 0.014323f
C375 VTAIL.n148 B 0.026451f
C376 VTAIL.n149 B 0.064036f
C377 VTAIL.n150 B 0.06827f
C378 VTAIL.n151 B 1.15417f
C379 VN.n0 B 0.038358f
C380 VN.t5 B 1.1279f
C381 VN.n1 B 0.035584f
C382 VN.t0 B 1.28532f
C383 VN.n2 B 0.483191f
C384 VN.t4 B 1.1279f
C385 VN.n3 B 0.50566f
C386 VN.n4 B 0.054224f
C387 VN.n5 B 0.24217f
C388 VN.n6 B 0.029094f
C389 VN.n7 B 0.029094f
C390 VN.n8 B 0.049366f
C391 VN.n9 B 0.045122f
C392 VN.n10 B 0.503926f
C393 VN.n11 B 0.038142f
C394 VN.n12 B 0.038358f
C395 VN.t2 B 1.1279f
C396 VN.n13 B 0.035584f
C397 VN.t3 B 1.28532f
C398 VN.n14 B 0.483191f
C399 VN.t1 B 1.1279f
C400 VN.n15 B 0.50566f
C401 VN.n16 B 0.054224f
C402 VN.n17 B 0.24217f
C403 VN.n18 B 0.029094f
C404 VN.n19 B 0.029094f
C405 VN.n20 B 0.049366f
C406 VN.n21 B 0.045122f
C407 VN.n22 B 0.503926f
C408 VN.n23 B 1.27645f
.ends

