* NGSPICE file created from diff_pair_sample_1709.ext - technology: sky130A

.subckt diff_pair_sample_1709 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X1 VTAIL.t7 VN.t0 VDD2.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X2 VDD1.t8 VP.t1 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=4.7619 ps=25.2 w=12.21 l=3.3
X3 VTAIL.t3 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X4 VTAIL.t16 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=0 ps=0 w=12.21 l=3.3
X6 VDD2.t7 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=2.01465 ps=12.54 w=12.21 l=3.3
X7 VDD1.t6 VP.t3 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=2.01465 ps=12.54 w=12.21 l=3.3
X8 VTAIL.t19 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X9 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X10 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=0 ps=0 w=12.21 l=3.3
X11 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=0 ps=0 w=12.21 l=3.3
X13 VDD2.t4 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X14 VDD2.t3 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=4.7619 ps=25.2 w=12.21 l=3.3
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=0 ps=0 w=12.21 l=3.3
X16 VDD2.t2 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=4.7619 ps=25.2 w=12.21 l=3.3
X17 VDD2.t1 VN.t8 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=2.01465 ps=12.54 w=12.21 l=3.3
X18 VTAIL.t9 VN.t9 VDD2.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X19 VDD1.t4 VP.t5 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X20 VTAIL.t15 VP.t6 VDD1.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X21 VDD1.t2 VP.t7 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=4.7619 pd=25.2 as=2.01465 ps=12.54 w=12.21 l=3.3
X22 VTAIL.t14 VP.t8 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=2.01465 ps=12.54 w=12.21 l=3.3
X23 VDD1.t0 VP.t9 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=2.01465 pd=12.54 as=4.7619 ps=25.2 w=12.21 l=3.3
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n20 161.3
R17 VP.n58 VP.n57 161.3
R18 VP.n59 VP.n19 161.3
R19 VP.n61 VP.n60 161.3
R20 VP.n62 VP.n18 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n111 VP.n110 161.3
R23 VP.n109 VP.n1 161.3
R24 VP.n108 VP.n107 161.3
R25 VP.n106 VP.n2 161.3
R26 VP.n105 VP.n104 161.3
R27 VP.n103 VP.n3 161.3
R28 VP.n102 VP.n101 161.3
R29 VP.n100 VP.n99 161.3
R30 VP.n98 VP.n5 161.3
R31 VP.n97 VP.n96 161.3
R32 VP.n95 VP.n6 161.3
R33 VP.n94 VP.n93 161.3
R34 VP.n92 VP.n7 161.3
R35 VP.n91 VP.n90 161.3
R36 VP.n89 VP.n8 161.3
R37 VP.n88 VP.n87 161.3
R38 VP.n86 VP.n9 161.3
R39 VP.n85 VP.n84 161.3
R40 VP.n83 VP.n10 161.3
R41 VP.n82 VP.n81 161.3
R42 VP.n80 VP.n11 161.3
R43 VP.n79 VP.n78 161.3
R44 VP.n77 VP.n76 161.3
R45 VP.n75 VP.n13 161.3
R46 VP.n74 VP.n73 161.3
R47 VP.n72 VP.n14 161.3
R48 VP.n71 VP.n70 161.3
R49 VP.n69 VP.n15 161.3
R50 VP.n68 VP.n67 161.3
R51 VP.n30 VP.t3 121.791
R52 VP.n8 VP.t5 89.1705
R53 VP.n16 VP.t7 89.1705
R54 VP.n12 VP.t8 89.1705
R55 VP.n4 VP.t2 89.1705
R56 VP.n0 VP.t1 89.1705
R57 VP.n25 VP.t0 89.1705
R58 VP.n17 VP.t9 89.1705
R59 VP.n21 VP.t4 89.1705
R60 VP.n29 VP.t6 89.1705
R61 VP.n66 VP.n16 77.3446
R62 VP.n112 VP.n0 77.3446
R63 VP.n65 VP.n17 77.3446
R64 VP.n30 VP.n29 68.1433
R65 VP.n66 VP.n65 57.1622
R66 VP.n85 VP.n10 56.5193
R67 VP.n93 VP.n6 56.5193
R68 VP.n46 VP.n23 56.5193
R69 VP.n38 VP.n27 56.5193
R70 VP.n74 VP.n14 45.8354
R71 VP.n104 VP.n2 45.8354
R72 VP.n57 VP.n19 45.8354
R73 VP.n70 VP.n14 35.1514
R74 VP.n108 VP.n2 35.1514
R75 VP.n61 VP.n19 35.1514
R76 VP.n69 VP.n68 24.4675
R77 VP.n70 VP.n69 24.4675
R78 VP.n75 VP.n74 24.4675
R79 VP.n76 VP.n75 24.4675
R80 VP.n80 VP.n79 24.4675
R81 VP.n81 VP.n80 24.4675
R82 VP.n81 VP.n10 24.4675
R83 VP.n86 VP.n85 24.4675
R84 VP.n87 VP.n86 24.4675
R85 VP.n87 VP.n8 24.4675
R86 VP.n91 VP.n8 24.4675
R87 VP.n92 VP.n91 24.4675
R88 VP.n93 VP.n92 24.4675
R89 VP.n97 VP.n6 24.4675
R90 VP.n98 VP.n97 24.4675
R91 VP.n99 VP.n98 24.4675
R92 VP.n103 VP.n102 24.4675
R93 VP.n104 VP.n103 24.4675
R94 VP.n109 VP.n108 24.4675
R95 VP.n110 VP.n109 24.4675
R96 VP.n62 VP.n61 24.4675
R97 VP.n63 VP.n62 24.4675
R98 VP.n50 VP.n23 24.4675
R99 VP.n51 VP.n50 24.4675
R100 VP.n52 VP.n51 24.4675
R101 VP.n56 VP.n55 24.4675
R102 VP.n57 VP.n56 24.4675
R103 VP.n39 VP.n38 24.4675
R104 VP.n40 VP.n39 24.4675
R105 VP.n40 VP.n25 24.4675
R106 VP.n44 VP.n25 24.4675
R107 VP.n45 VP.n44 24.4675
R108 VP.n46 VP.n45 24.4675
R109 VP.n33 VP.n32 24.4675
R110 VP.n34 VP.n33 24.4675
R111 VP.n34 VP.n27 24.4675
R112 VP.n76 VP.n12 18.1061
R113 VP.n102 VP.n4 18.1061
R114 VP.n55 VP.n21 18.1061
R115 VP.n68 VP.n16 12.7233
R116 VP.n110 VP.n0 12.7233
R117 VP.n63 VP.n17 12.7233
R118 VP.n79 VP.n12 6.36192
R119 VP.n99 VP.n4 6.36192
R120 VP.n52 VP.n21 6.36192
R121 VP.n32 VP.n29 6.36192
R122 VP.n31 VP.n30 4.26089
R123 VP.n65 VP.n64 0.354971
R124 VP.n67 VP.n66 0.354971
R125 VP.n112 VP.n111 0.354971
R126 VP VP.n112 0.26696
R127 VP.n31 VP.n28 0.189894
R128 VP.n35 VP.n28 0.189894
R129 VP.n36 VP.n35 0.189894
R130 VP.n37 VP.n36 0.189894
R131 VP.n37 VP.n26 0.189894
R132 VP.n41 VP.n26 0.189894
R133 VP.n42 VP.n41 0.189894
R134 VP.n43 VP.n42 0.189894
R135 VP.n43 VP.n24 0.189894
R136 VP.n47 VP.n24 0.189894
R137 VP.n48 VP.n47 0.189894
R138 VP.n49 VP.n48 0.189894
R139 VP.n49 VP.n22 0.189894
R140 VP.n53 VP.n22 0.189894
R141 VP.n54 VP.n53 0.189894
R142 VP.n54 VP.n20 0.189894
R143 VP.n58 VP.n20 0.189894
R144 VP.n59 VP.n58 0.189894
R145 VP.n60 VP.n59 0.189894
R146 VP.n60 VP.n18 0.189894
R147 VP.n64 VP.n18 0.189894
R148 VP.n67 VP.n15 0.189894
R149 VP.n71 VP.n15 0.189894
R150 VP.n72 VP.n71 0.189894
R151 VP.n73 VP.n72 0.189894
R152 VP.n73 VP.n13 0.189894
R153 VP.n77 VP.n13 0.189894
R154 VP.n78 VP.n77 0.189894
R155 VP.n78 VP.n11 0.189894
R156 VP.n82 VP.n11 0.189894
R157 VP.n83 VP.n82 0.189894
R158 VP.n84 VP.n83 0.189894
R159 VP.n84 VP.n9 0.189894
R160 VP.n88 VP.n9 0.189894
R161 VP.n89 VP.n88 0.189894
R162 VP.n90 VP.n89 0.189894
R163 VP.n90 VP.n7 0.189894
R164 VP.n94 VP.n7 0.189894
R165 VP.n95 VP.n94 0.189894
R166 VP.n96 VP.n95 0.189894
R167 VP.n96 VP.n5 0.189894
R168 VP.n100 VP.n5 0.189894
R169 VP.n101 VP.n100 0.189894
R170 VP.n101 VP.n3 0.189894
R171 VP.n105 VP.n3 0.189894
R172 VP.n106 VP.n105 0.189894
R173 VP.n107 VP.n106 0.189894
R174 VP.n107 VP.n1 0.189894
R175 VP.n111 VP.n1 0.189894
R176 VTAIL.n272 VTAIL.n212 289.615
R177 VTAIL.n62 VTAIL.n2 289.615
R178 VTAIL.n206 VTAIL.n146 289.615
R179 VTAIL.n136 VTAIL.n76 289.615
R180 VTAIL.n232 VTAIL.n231 185
R181 VTAIL.n237 VTAIL.n236 185
R182 VTAIL.n239 VTAIL.n238 185
R183 VTAIL.n228 VTAIL.n227 185
R184 VTAIL.n245 VTAIL.n244 185
R185 VTAIL.n247 VTAIL.n246 185
R186 VTAIL.n224 VTAIL.n223 185
R187 VTAIL.n254 VTAIL.n253 185
R188 VTAIL.n255 VTAIL.n222 185
R189 VTAIL.n257 VTAIL.n256 185
R190 VTAIL.n220 VTAIL.n219 185
R191 VTAIL.n263 VTAIL.n262 185
R192 VTAIL.n265 VTAIL.n264 185
R193 VTAIL.n216 VTAIL.n215 185
R194 VTAIL.n271 VTAIL.n270 185
R195 VTAIL.n273 VTAIL.n272 185
R196 VTAIL.n22 VTAIL.n21 185
R197 VTAIL.n27 VTAIL.n26 185
R198 VTAIL.n29 VTAIL.n28 185
R199 VTAIL.n18 VTAIL.n17 185
R200 VTAIL.n35 VTAIL.n34 185
R201 VTAIL.n37 VTAIL.n36 185
R202 VTAIL.n14 VTAIL.n13 185
R203 VTAIL.n44 VTAIL.n43 185
R204 VTAIL.n45 VTAIL.n12 185
R205 VTAIL.n47 VTAIL.n46 185
R206 VTAIL.n10 VTAIL.n9 185
R207 VTAIL.n53 VTAIL.n52 185
R208 VTAIL.n55 VTAIL.n54 185
R209 VTAIL.n6 VTAIL.n5 185
R210 VTAIL.n61 VTAIL.n60 185
R211 VTAIL.n63 VTAIL.n62 185
R212 VTAIL.n207 VTAIL.n206 185
R213 VTAIL.n205 VTAIL.n204 185
R214 VTAIL.n150 VTAIL.n149 185
R215 VTAIL.n199 VTAIL.n198 185
R216 VTAIL.n197 VTAIL.n196 185
R217 VTAIL.n154 VTAIL.n153 185
R218 VTAIL.n191 VTAIL.n190 185
R219 VTAIL.n189 VTAIL.n156 185
R220 VTAIL.n188 VTAIL.n187 185
R221 VTAIL.n159 VTAIL.n157 185
R222 VTAIL.n182 VTAIL.n181 185
R223 VTAIL.n180 VTAIL.n179 185
R224 VTAIL.n163 VTAIL.n162 185
R225 VTAIL.n174 VTAIL.n173 185
R226 VTAIL.n172 VTAIL.n171 185
R227 VTAIL.n167 VTAIL.n166 185
R228 VTAIL.n137 VTAIL.n136 185
R229 VTAIL.n135 VTAIL.n134 185
R230 VTAIL.n80 VTAIL.n79 185
R231 VTAIL.n129 VTAIL.n128 185
R232 VTAIL.n127 VTAIL.n126 185
R233 VTAIL.n84 VTAIL.n83 185
R234 VTAIL.n121 VTAIL.n120 185
R235 VTAIL.n119 VTAIL.n86 185
R236 VTAIL.n118 VTAIL.n117 185
R237 VTAIL.n89 VTAIL.n87 185
R238 VTAIL.n112 VTAIL.n111 185
R239 VTAIL.n110 VTAIL.n109 185
R240 VTAIL.n93 VTAIL.n92 185
R241 VTAIL.n104 VTAIL.n103 185
R242 VTAIL.n102 VTAIL.n101 185
R243 VTAIL.n97 VTAIL.n96 185
R244 VTAIL.n233 VTAIL.t1 149.524
R245 VTAIL.n23 VTAIL.t12 149.524
R246 VTAIL.n168 VTAIL.t18 149.524
R247 VTAIL.n98 VTAIL.t0 149.524
R248 VTAIL.n237 VTAIL.n231 104.615
R249 VTAIL.n238 VTAIL.n237 104.615
R250 VTAIL.n238 VTAIL.n227 104.615
R251 VTAIL.n245 VTAIL.n227 104.615
R252 VTAIL.n246 VTAIL.n245 104.615
R253 VTAIL.n246 VTAIL.n223 104.615
R254 VTAIL.n254 VTAIL.n223 104.615
R255 VTAIL.n255 VTAIL.n254 104.615
R256 VTAIL.n256 VTAIL.n255 104.615
R257 VTAIL.n256 VTAIL.n219 104.615
R258 VTAIL.n263 VTAIL.n219 104.615
R259 VTAIL.n264 VTAIL.n263 104.615
R260 VTAIL.n264 VTAIL.n215 104.615
R261 VTAIL.n271 VTAIL.n215 104.615
R262 VTAIL.n272 VTAIL.n271 104.615
R263 VTAIL.n27 VTAIL.n21 104.615
R264 VTAIL.n28 VTAIL.n27 104.615
R265 VTAIL.n28 VTAIL.n17 104.615
R266 VTAIL.n35 VTAIL.n17 104.615
R267 VTAIL.n36 VTAIL.n35 104.615
R268 VTAIL.n36 VTAIL.n13 104.615
R269 VTAIL.n44 VTAIL.n13 104.615
R270 VTAIL.n45 VTAIL.n44 104.615
R271 VTAIL.n46 VTAIL.n45 104.615
R272 VTAIL.n46 VTAIL.n9 104.615
R273 VTAIL.n53 VTAIL.n9 104.615
R274 VTAIL.n54 VTAIL.n53 104.615
R275 VTAIL.n54 VTAIL.n5 104.615
R276 VTAIL.n61 VTAIL.n5 104.615
R277 VTAIL.n62 VTAIL.n61 104.615
R278 VTAIL.n206 VTAIL.n205 104.615
R279 VTAIL.n205 VTAIL.n149 104.615
R280 VTAIL.n198 VTAIL.n149 104.615
R281 VTAIL.n198 VTAIL.n197 104.615
R282 VTAIL.n197 VTAIL.n153 104.615
R283 VTAIL.n190 VTAIL.n153 104.615
R284 VTAIL.n190 VTAIL.n189 104.615
R285 VTAIL.n189 VTAIL.n188 104.615
R286 VTAIL.n188 VTAIL.n157 104.615
R287 VTAIL.n181 VTAIL.n157 104.615
R288 VTAIL.n181 VTAIL.n180 104.615
R289 VTAIL.n180 VTAIL.n162 104.615
R290 VTAIL.n173 VTAIL.n162 104.615
R291 VTAIL.n173 VTAIL.n172 104.615
R292 VTAIL.n172 VTAIL.n166 104.615
R293 VTAIL.n136 VTAIL.n135 104.615
R294 VTAIL.n135 VTAIL.n79 104.615
R295 VTAIL.n128 VTAIL.n79 104.615
R296 VTAIL.n128 VTAIL.n127 104.615
R297 VTAIL.n127 VTAIL.n83 104.615
R298 VTAIL.n120 VTAIL.n83 104.615
R299 VTAIL.n120 VTAIL.n119 104.615
R300 VTAIL.n119 VTAIL.n118 104.615
R301 VTAIL.n118 VTAIL.n87 104.615
R302 VTAIL.n111 VTAIL.n87 104.615
R303 VTAIL.n111 VTAIL.n110 104.615
R304 VTAIL.n110 VTAIL.n92 104.615
R305 VTAIL.n103 VTAIL.n92 104.615
R306 VTAIL.n103 VTAIL.n102 104.615
R307 VTAIL.n102 VTAIL.n96 104.615
R308 VTAIL.t1 VTAIL.n231 52.3082
R309 VTAIL.t12 VTAIL.n21 52.3082
R310 VTAIL.t18 VTAIL.n166 52.3082
R311 VTAIL.t0 VTAIL.n96 52.3082
R312 VTAIL.n145 VTAIL.n144 46.9466
R313 VTAIL.n143 VTAIL.n142 46.9466
R314 VTAIL.n75 VTAIL.n74 46.9466
R315 VTAIL.n73 VTAIL.n72 46.9466
R316 VTAIL.n279 VTAIL.n278 46.9464
R317 VTAIL.n1 VTAIL.n0 46.9464
R318 VTAIL.n69 VTAIL.n68 46.9464
R319 VTAIL.n71 VTAIL.n70 46.9464
R320 VTAIL.n277 VTAIL.n276 33.9308
R321 VTAIL.n67 VTAIL.n66 33.9308
R322 VTAIL.n211 VTAIL.n210 33.9308
R323 VTAIL.n141 VTAIL.n140 33.9308
R324 VTAIL.n73 VTAIL.n71 29.1514
R325 VTAIL.n277 VTAIL.n211 26.0221
R326 VTAIL.n257 VTAIL.n222 13.1884
R327 VTAIL.n47 VTAIL.n12 13.1884
R328 VTAIL.n191 VTAIL.n156 13.1884
R329 VTAIL.n121 VTAIL.n86 13.1884
R330 VTAIL.n253 VTAIL.n252 12.8005
R331 VTAIL.n258 VTAIL.n220 12.8005
R332 VTAIL.n43 VTAIL.n42 12.8005
R333 VTAIL.n48 VTAIL.n10 12.8005
R334 VTAIL.n192 VTAIL.n154 12.8005
R335 VTAIL.n187 VTAIL.n158 12.8005
R336 VTAIL.n122 VTAIL.n84 12.8005
R337 VTAIL.n117 VTAIL.n88 12.8005
R338 VTAIL.n251 VTAIL.n224 12.0247
R339 VTAIL.n262 VTAIL.n261 12.0247
R340 VTAIL.n41 VTAIL.n14 12.0247
R341 VTAIL.n52 VTAIL.n51 12.0247
R342 VTAIL.n196 VTAIL.n195 12.0247
R343 VTAIL.n186 VTAIL.n159 12.0247
R344 VTAIL.n126 VTAIL.n125 12.0247
R345 VTAIL.n116 VTAIL.n89 12.0247
R346 VTAIL.n248 VTAIL.n247 11.249
R347 VTAIL.n265 VTAIL.n218 11.249
R348 VTAIL.n38 VTAIL.n37 11.249
R349 VTAIL.n55 VTAIL.n8 11.249
R350 VTAIL.n199 VTAIL.n152 11.249
R351 VTAIL.n183 VTAIL.n182 11.249
R352 VTAIL.n129 VTAIL.n82 11.249
R353 VTAIL.n113 VTAIL.n112 11.249
R354 VTAIL.n244 VTAIL.n226 10.4732
R355 VTAIL.n266 VTAIL.n216 10.4732
R356 VTAIL.n34 VTAIL.n16 10.4732
R357 VTAIL.n56 VTAIL.n6 10.4732
R358 VTAIL.n200 VTAIL.n150 10.4732
R359 VTAIL.n179 VTAIL.n161 10.4732
R360 VTAIL.n130 VTAIL.n80 10.4732
R361 VTAIL.n109 VTAIL.n91 10.4732
R362 VTAIL.n233 VTAIL.n232 10.2747
R363 VTAIL.n23 VTAIL.n22 10.2747
R364 VTAIL.n168 VTAIL.n167 10.2747
R365 VTAIL.n98 VTAIL.n97 10.2747
R366 VTAIL.n243 VTAIL.n228 9.69747
R367 VTAIL.n270 VTAIL.n269 9.69747
R368 VTAIL.n33 VTAIL.n18 9.69747
R369 VTAIL.n60 VTAIL.n59 9.69747
R370 VTAIL.n204 VTAIL.n203 9.69747
R371 VTAIL.n178 VTAIL.n163 9.69747
R372 VTAIL.n134 VTAIL.n133 9.69747
R373 VTAIL.n108 VTAIL.n93 9.69747
R374 VTAIL.n276 VTAIL.n275 9.45567
R375 VTAIL.n66 VTAIL.n65 9.45567
R376 VTAIL.n210 VTAIL.n209 9.45567
R377 VTAIL.n140 VTAIL.n139 9.45567
R378 VTAIL.n275 VTAIL.n274 9.3005
R379 VTAIL.n214 VTAIL.n213 9.3005
R380 VTAIL.n269 VTAIL.n268 9.3005
R381 VTAIL.n267 VTAIL.n266 9.3005
R382 VTAIL.n218 VTAIL.n217 9.3005
R383 VTAIL.n261 VTAIL.n260 9.3005
R384 VTAIL.n259 VTAIL.n258 9.3005
R385 VTAIL.n235 VTAIL.n234 9.3005
R386 VTAIL.n230 VTAIL.n229 9.3005
R387 VTAIL.n241 VTAIL.n240 9.3005
R388 VTAIL.n243 VTAIL.n242 9.3005
R389 VTAIL.n226 VTAIL.n225 9.3005
R390 VTAIL.n249 VTAIL.n248 9.3005
R391 VTAIL.n251 VTAIL.n250 9.3005
R392 VTAIL.n252 VTAIL.n221 9.3005
R393 VTAIL.n65 VTAIL.n64 9.3005
R394 VTAIL.n4 VTAIL.n3 9.3005
R395 VTAIL.n59 VTAIL.n58 9.3005
R396 VTAIL.n57 VTAIL.n56 9.3005
R397 VTAIL.n8 VTAIL.n7 9.3005
R398 VTAIL.n51 VTAIL.n50 9.3005
R399 VTAIL.n49 VTAIL.n48 9.3005
R400 VTAIL.n25 VTAIL.n24 9.3005
R401 VTAIL.n20 VTAIL.n19 9.3005
R402 VTAIL.n31 VTAIL.n30 9.3005
R403 VTAIL.n33 VTAIL.n32 9.3005
R404 VTAIL.n16 VTAIL.n15 9.3005
R405 VTAIL.n39 VTAIL.n38 9.3005
R406 VTAIL.n41 VTAIL.n40 9.3005
R407 VTAIL.n42 VTAIL.n11 9.3005
R408 VTAIL.n170 VTAIL.n169 9.3005
R409 VTAIL.n165 VTAIL.n164 9.3005
R410 VTAIL.n176 VTAIL.n175 9.3005
R411 VTAIL.n178 VTAIL.n177 9.3005
R412 VTAIL.n161 VTAIL.n160 9.3005
R413 VTAIL.n184 VTAIL.n183 9.3005
R414 VTAIL.n186 VTAIL.n185 9.3005
R415 VTAIL.n158 VTAIL.n155 9.3005
R416 VTAIL.n209 VTAIL.n208 9.3005
R417 VTAIL.n148 VTAIL.n147 9.3005
R418 VTAIL.n203 VTAIL.n202 9.3005
R419 VTAIL.n201 VTAIL.n200 9.3005
R420 VTAIL.n152 VTAIL.n151 9.3005
R421 VTAIL.n195 VTAIL.n194 9.3005
R422 VTAIL.n193 VTAIL.n192 9.3005
R423 VTAIL.n100 VTAIL.n99 9.3005
R424 VTAIL.n95 VTAIL.n94 9.3005
R425 VTAIL.n106 VTAIL.n105 9.3005
R426 VTAIL.n108 VTAIL.n107 9.3005
R427 VTAIL.n91 VTAIL.n90 9.3005
R428 VTAIL.n114 VTAIL.n113 9.3005
R429 VTAIL.n116 VTAIL.n115 9.3005
R430 VTAIL.n88 VTAIL.n85 9.3005
R431 VTAIL.n139 VTAIL.n138 9.3005
R432 VTAIL.n78 VTAIL.n77 9.3005
R433 VTAIL.n133 VTAIL.n132 9.3005
R434 VTAIL.n131 VTAIL.n130 9.3005
R435 VTAIL.n82 VTAIL.n81 9.3005
R436 VTAIL.n125 VTAIL.n124 9.3005
R437 VTAIL.n123 VTAIL.n122 9.3005
R438 VTAIL.n240 VTAIL.n239 8.92171
R439 VTAIL.n273 VTAIL.n214 8.92171
R440 VTAIL.n30 VTAIL.n29 8.92171
R441 VTAIL.n63 VTAIL.n4 8.92171
R442 VTAIL.n207 VTAIL.n148 8.92171
R443 VTAIL.n175 VTAIL.n174 8.92171
R444 VTAIL.n137 VTAIL.n78 8.92171
R445 VTAIL.n105 VTAIL.n104 8.92171
R446 VTAIL.n236 VTAIL.n230 8.14595
R447 VTAIL.n274 VTAIL.n212 8.14595
R448 VTAIL.n26 VTAIL.n20 8.14595
R449 VTAIL.n64 VTAIL.n2 8.14595
R450 VTAIL.n208 VTAIL.n146 8.14595
R451 VTAIL.n171 VTAIL.n165 8.14595
R452 VTAIL.n138 VTAIL.n76 8.14595
R453 VTAIL.n101 VTAIL.n95 8.14595
R454 VTAIL.n235 VTAIL.n232 7.3702
R455 VTAIL.n25 VTAIL.n22 7.3702
R456 VTAIL.n170 VTAIL.n167 7.3702
R457 VTAIL.n100 VTAIL.n97 7.3702
R458 VTAIL.n236 VTAIL.n235 5.81868
R459 VTAIL.n276 VTAIL.n212 5.81868
R460 VTAIL.n26 VTAIL.n25 5.81868
R461 VTAIL.n66 VTAIL.n2 5.81868
R462 VTAIL.n210 VTAIL.n146 5.81868
R463 VTAIL.n171 VTAIL.n170 5.81868
R464 VTAIL.n140 VTAIL.n76 5.81868
R465 VTAIL.n101 VTAIL.n100 5.81868
R466 VTAIL.n239 VTAIL.n230 5.04292
R467 VTAIL.n274 VTAIL.n273 5.04292
R468 VTAIL.n29 VTAIL.n20 5.04292
R469 VTAIL.n64 VTAIL.n63 5.04292
R470 VTAIL.n208 VTAIL.n207 5.04292
R471 VTAIL.n174 VTAIL.n165 5.04292
R472 VTAIL.n138 VTAIL.n137 5.04292
R473 VTAIL.n104 VTAIL.n95 5.04292
R474 VTAIL.n240 VTAIL.n228 4.26717
R475 VTAIL.n270 VTAIL.n214 4.26717
R476 VTAIL.n30 VTAIL.n18 4.26717
R477 VTAIL.n60 VTAIL.n4 4.26717
R478 VTAIL.n204 VTAIL.n148 4.26717
R479 VTAIL.n175 VTAIL.n163 4.26717
R480 VTAIL.n134 VTAIL.n78 4.26717
R481 VTAIL.n105 VTAIL.n93 4.26717
R482 VTAIL.n244 VTAIL.n243 3.49141
R483 VTAIL.n269 VTAIL.n216 3.49141
R484 VTAIL.n34 VTAIL.n33 3.49141
R485 VTAIL.n59 VTAIL.n6 3.49141
R486 VTAIL.n203 VTAIL.n150 3.49141
R487 VTAIL.n179 VTAIL.n178 3.49141
R488 VTAIL.n133 VTAIL.n80 3.49141
R489 VTAIL.n109 VTAIL.n108 3.49141
R490 VTAIL.n75 VTAIL.n73 3.12981
R491 VTAIL.n141 VTAIL.n75 3.12981
R492 VTAIL.n145 VTAIL.n143 3.12981
R493 VTAIL.n211 VTAIL.n145 3.12981
R494 VTAIL.n71 VTAIL.n69 3.12981
R495 VTAIL.n69 VTAIL.n67 3.12981
R496 VTAIL.n279 VTAIL.n277 3.12981
R497 VTAIL.n234 VTAIL.n233 2.84303
R498 VTAIL.n24 VTAIL.n23 2.84303
R499 VTAIL.n169 VTAIL.n168 2.84303
R500 VTAIL.n99 VTAIL.n98 2.84303
R501 VTAIL.n247 VTAIL.n226 2.71565
R502 VTAIL.n266 VTAIL.n265 2.71565
R503 VTAIL.n37 VTAIL.n16 2.71565
R504 VTAIL.n56 VTAIL.n55 2.71565
R505 VTAIL.n200 VTAIL.n199 2.71565
R506 VTAIL.n182 VTAIL.n161 2.71565
R507 VTAIL.n130 VTAIL.n129 2.71565
R508 VTAIL.n112 VTAIL.n91 2.71565
R509 VTAIL VTAIL.n1 2.40567
R510 VTAIL.n143 VTAIL.n141 2.03498
R511 VTAIL.n67 VTAIL.n1 2.03498
R512 VTAIL.n248 VTAIL.n224 1.93989
R513 VTAIL.n262 VTAIL.n218 1.93989
R514 VTAIL.n38 VTAIL.n14 1.93989
R515 VTAIL.n52 VTAIL.n8 1.93989
R516 VTAIL.n196 VTAIL.n152 1.93989
R517 VTAIL.n183 VTAIL.n159 1.93989
R518 VTAIL.n126 VTAIL.n82 1.93989
R519 VTAIL.n113 VTAIL.n89 1.93989
R520 VTAIL.n278 VTAIL.t6 1.62212
R521 VTAIL.n278 VTAIL.t4 1.62212
R522 VTAIL.n0 VTAIL.t8 1.62212
R523 VTAIL.n0 VTAIL.t9 1.62212
R524 VTAIL.n68 VTAIL.t13 1.62212
R525 VTAIL.n68 VTAIL.t16 1.62212
R526 VTAIL.n70 VTAIL.t10 1.62212
R527 VTAIL.n70 VTAIL.t14 1.62212
R528 VTAIL.n144 VTAIL.t11 1.62212
R529 VTAIL.n144 VTAIL.t19 1.62212
R530 VTAIL.n142 VTAIL.t17 1.62212
R531 VTAIL.n142 VTAIL.t15 1.62212
R532 VTAIL.n74 VTAIL.t5 1.62212
R533 VTAIL.n74 VTAIL.t3 1.62212
R534 VTAIL.n72 VTAIL.t2 1.62212
R535 VTAIL.n72 VTAIL.t7 1.62212
R536 VTAIL.n253 VTAIL.n251 1.16414
R537 VTAIL.n261 VTAIL.n220 1.16414
R538 VTAIL.n43 VTAIL.n41 1.16414
R539 VTAIL.n51 VTAIL.n10 1.16414
R540 VTAIL.n195 VTAIL.n154 1.16414
R541 VTAIL.n187 VTAIL.n186 1.16414
R542 VTAIL.n125 VTAIL.n84 1.16414
R543 VTAIL.n117 VTAIL.n116 1.16414
R544 VTAIL VTAIL.n279 0.724638
R545 VTAIL.n252 VTAIL.n222 0.388379
R546 VTAIL.n258 VTAIL.n257 0.388379
R547 VTAIL.n42 VTAIL.n12 0.388379
R548 VTAIL.n48 VTAIL.n47 0.388379
R549 VTAIL.n192 VTAIL.n191 0.388379
R550 VTAIL.n158 VTAIL.n156 0.388379
R551 VTAIL.n122 VTAIL.n121 0.388379
R552 VTAIL.n88 VTAIL.n86 0.388379
R553 VTAIL.n234 VTAIL.n229 0.155672
R554 VTAIL.n241 VTAIL.n229 0.155672
R555 VTAIL.n242 VTAIL.n241 0.155672
R556 VTAIL.n242 VTAIL.n225 0.155672
R557 VTAIL.n249 VTAIL.n225 0.155672
R558 VTAIL.n250 VTAIL.n249 0.155672
R559 VTAIL.n250 VTAIL.n221 0.155672
R560 VTAIL.n259 VTAIL.n221 0.155672
R561 VTAIL.n260 VTAIL.n259 0.155672
R562 VTAIL.n260 VTAIL.n217 0.155672
R563 VTAIL.n267 VTAIL.n217 0.155672
R564 VTAIL.n268 VTAIL.n267 0.155672
R565 VTAIL.n268 VTAIL.n213 0.155672
R566 VTAIL.n275 VTAIL.n213 0.155672
R567 VTAIL.n24 VTAIL.n19 0.155672
R568 VTAIL.n31 VTAIL.n19 0.155672
R569 VTAIL.n32 VTAIL.n31 0.155672
R570 VTAIL.n32 VTAIL.n15 0.155672
R571 VTAIL.n39 VTAIL.n15 0.155672
R572 VTAIL.n40 VTAIL.n39 0.155672
R573 VTAIL.n40 VTAIL.n11 0.155672
R574 VTAIL.n49 VTAIL.n11 0.155672
R575 VTAIL.n50 VTAIL.n49 0.155672
R576 VTAIL.n50 VTAIL.n7 0.155672
R577 VTAIL.n57 VTAIL.n7 0.155672
R578 VTAIL.n58 VTAIL.n57 0.155672
R579 VTAIL.n58 VTAIL.n3 0.155672
R580 VTAIL.n65 VTAIL.n3 0.155672
R581 VTAIL.n209 VTAIL.n147 0.155672
R582 VTAIL.n202 VTAIL.n147 0.155672
R583 VTAIL.n202 VTAIL.n201 0.155672
R584 VTAIL.n201 VTAIL.n151 0.155672
R585 VTAIL.n194 VTAIL.n151 0.155672
R586 VTAIL.n194 VTAIL.n193 0.155672
R587 VTAIL.n193 VTAIL.n155 0.155672
R588 VTAIL.n185 VTAIL.n155 0.155672
R589 VTAIL.n185 VTAIL.n184 0.155672
R590 VTAIL.n184 VTAIL.n160 0.155672
R591 VTAIL.n177 VTAIL.n160 0.155672
R592 VTAIL.n177 VTAIL.n176 0.155672
R593 VTAIL.n176 VTAIL.n164 0.155672
R594 VTAIL.n169 VTAIL.n164 0.155672
R595 VTAIL.n139 VTAIL.n77 0.155672
R596 VTAIL.n132 VTAIL.n77 0.155672
R597 VTAIL.n132 VTAIL.n131 0.155672
R598 VTAIL.n131 VTAIL.n81 0.155672
R599 VTAIL.n124 VTAIL.n81 0.155672
R600 VTAIL.n124 VTAIL.n123 0.155672
R601 VTAIL.n123 VTAIL.n85 0.155672
R602 VTAIL.n115 VTAIL.n85 0.155672
R603 VTAIL.n115 VTAIL.n114 0.155672
R604 VTAIL.n114 VTAIL.n90 0.155672
R605 VTAIL.n107 VTAIL.n90 0.155672
R606 VTAIL.n107 VTAIL.n106 0.155672
R607 VTAIL.n106 VTAIL.n94 0.155672
R608 VTAIL.n99 VTAIL.n94 0.155672
R609 VDD1.n60 VDD1.n0 289.615
R610 VDD1.n127 VDD1.n67 289.615
R611 VDD1.n61 VDD1.n60 185
R612 VDD1.n59 VDD1.n58 185
R613 VDD1.n4 VDD1.n3 185
R614 VDD1.n53 VDD1.n52 185
R615 VDD1.n51 VDD1.n50 185
R616 VDD1.n8 VDD1.n7 185
R617 VDD1.n45 VDD1.n44 185
R618 VDD1.n43 VDD1.n10 185
R619 VDD1.n42 VDD1.n41 185
R620 VDD1.n13 VDD1.n11 185
R621 VDD1.n36 VDD1.n35 185
R622 VDD1.n34 VDD1.n33 185
R623 VDD1.n17 VDD1.n16 185
R624 VDD1.n28 VDD1.n27 185
R625 VDD1.n26 VDD1.n25 185
R626 VDD1.n21 VDD1.n20 185
R627 VDD1.n87 VDD1.n86 185
R628 VDD1.n92 VDD1.n91 185
R629 VDD1.n94 VDD1.n93 185
R630 VDD1.n83 VDD1.n82 185
R631 VDD1.n100 VDD1.n99 185
R632 VDD1.n102 VDD1.n101 185
R633 VDD1.n79 VDD1.n78 185
R634 VDD1.n109 VDD1.n108 185
R635 VDD1.n110 VDD1.n77 185
R636 VDD1.n112 VDD1.n111 185
R637 VDD1.n75 VDD1.n74 185
R638 VDD1.n118 VDD1.n117 185
R639 VDD1.n120 VDD1.n119 185
R640 VDD1.n71 VDD1.n70 185
R641 VDD1.n126 VDD1.n125 185
R642 VDD1.n128 VDD1.n127 185
R643 VDD1.n22 VDD1.t6 149.524
R644 VDD1.n88 VDD1.t2 149.524
R645 VDD1.n60 VDD1.n59 104.615
R646 VDD1.n59 VDD1.n3 104.615
R647 VDD1.n52 VDD1.n3 104.615
R648 VDD1.n52 VDD1.n51 104.615
R649 VDD1.n51 VDD1.n7 104.615
R650 VDD1.n44 VDD1.n7 104.615
R651 VDD1.n44 VDD1.n43 104.615
R652 VDD1.n43 VDD1.n42 104.615
R653 VDD1.n42 VDD1.n11 104.615
R654 VDD1.n35 VDD1.n11 104.615
R655 VDD1.n35 VDD1.n34 104.615
R656 VDD1.n34 VDD1.n16 104.615
R657 VDD1.n27 VDD1.n16 104.615
R658 VDD1.n27 VDD1.n26 104.615
R659 VDD1.n26 VDD1.n20 104.615
R660 VDD1.n92 VDD1.n86 104.615
R661 VDD1.n93 VDD1.n92 104.615
R662 VDD1.n93 VDD1.n82 104.615
R663 VDD1.n100 VDD1.n82 104.615
R664 VDD1.n101 VDD1.n100 104.615
R665 VDD1.n101 VDD1.n78 104.615
R666 VDD1.n109 VDD1.n78 104.615
R667 VDD1.n110 VDD1.n109 104.615
R668 VDD1.n111 VDD1.n110 104.615
R669 VDD1.n111 VDD1.n74 104.615
R670 VDD1.n118 VDD1.n74 104.615
R671 VDD1.n119 VDD1.n118 104.615
R672 VDD1.n119 VDD1.n70 104.615
R673 VDD1.n126 VDD1.n70 104.615
R674 VDD1.n127 VDD1.n126 104.615
R675 VDD1.n135 VDD1.n134 65.9169
R676 VDD1.n66 VDD1.n65 63.6254
R677 VDD1.n137 VDD1.n136 63.6252
R678 VDD1.n133 VDD1.n132 63.6252
R679 VDD1.n66 VDD1.n64 53.7389
R680 VDD1.n133 VDD1.n131 53.7389
R681 VDD1.t6 VDD1.n20 52.3082
R682 VDD1.t2 VDD1.n86 52.3082
R683 VDD1.n137 VDD1.n135 51.253
R684 VDD1.n45 VDD1.n10 13.1884
R685 VDD1.n112 VDD1.n77 13.1884
R686 VDD1.n46 VDD1.n8 12.8005
R687 VDD1.n41 VDD1.n12 12.8005
R688 VDD1.n108 VDD1.n107 12.8005
R689 VDD1.n113 VDD1.n75 12.8005
R690 VDD1.n50 VDD1.n49 12.0247
R691 VDD1.n40 VDD1.n13 12.0247
R692 VDD1.n106 VDD1.n79 12.0247
R693 VDD1.n117 VDD1.n116 12.0247
R694 VDD1.n53 VDD1.n6 11.249
R695 VDD1.n37 VDD1.n36 11.249
R696 VDD1.n103 VDD1.n102 11.249
R697 VDD1.n120 VDD1.n73 11.249
R698 VDD1.n54 VDD1.n4 10.4732
R699 VDD1.n33 VDD1.n15 10.4732
R700 VDD1.n99 VDD1.n81 10.4732
R701 VDD1.n121 VDD1.n71 10.4732
R702 VDD1.n22 VDD1.n21 10.2747
R703 VDD1.n88 VDD1.n87 10.2747
R704 VDD1.n58 VDD1.n57 9.69747
R705 VDD1.n32 VDD1.n17 9.69747
R706 VDD1.n98 VDD1.n83 9.69747
R707 VDD1.n125 VDD1.n124 9.69747
R708 VDD1.n64 VDD1.n63 9.45567
R709 VDD1.n131 VDD1.n130 9.45567
R710 VDD1.n24 VDD1.n23 9.3005
R711 VDD1.n19 VDD1.n18 9.3005
R712 VDD1.n30 VDD1.n29 9.3005
R713 VDD1.n32 VDD1.n31 9.3005
R714 VDD1.n15 VDD1.n14 9.3005
R715 VDD1.n38 VDD1.n37 9.3005
R716 VDD1.n40 VDD1.n39 9.3005
R717 VDD1.n12 VDD1.n9 9.3005
R718 VDD1.n63 VDD1.n62 9.3005
R719 VDD1.n2 VDD1.n1 9.3005
R720 VDD1.n57 VDD1.n56 9.3005
R721 VDD1.n55 VDD1.n54 9.3005
R722 VDD1.n6 VDD1.n5 9.3005
R723 VDD1.n49 VDD1.n48 9.3005
R724 VDD1.n47 VDD1.n46 9.3005
R725 VDD1.n130 VDD1.n129 9.3005
R726 VDD1.n69 VDD1.n68 9.3005
R727 VDD1.n124 VDD1.n123 9.3005
R728 VDD1.n122 VDD1.n121 9.3005
R729 VDD1.n73 VDD1.n72 9.3005
R730 VDD1.n116 VDD1.n115 9.3005
R731 VDD1.n114 VDD1.n113 9.3005
R732 VDD1.n90 VDD1.n89 9.3005
R733 VDD1.n85 VDD1.n84 9.3005
R734 VDD1.n96 VDD1.n95 9.3005
R735 VDD1.n98 VDD1.n97 9.3005
R736 VDD1.n81 VDD1.n80 9.3005
R737 VDD1.n104 VDD1.n103 9.3005
R738 VDD1.n106 VDD1.n105 9.3005
R739 VDD1.n107 VDD1.n76 9.3005
R740 VDD1.n61 VDD1.n2 8.92171
R741 VDD1.n29 VDD1.n28 8.92171
R742 VDD1.n95 VDD1.n94 8.92171
R743 VDD1.n128 VDD1.n69 8.92171
R744 VDD1.n62 VDD1.n0 8.14595
R745 VDD1.n25 VDD1.n19 8.14595
R746 VDD1.n91 VDD1.n85 8.14595
R747 VDD1.n129 VDD1.n67 8.14595
R748 VDD1.n24 VDD1.n21 7.3702
R749 VDD1.n90 VDD1.n87 7.3702
R750 VDD1.n64 VDD1.n0 5.81868
R751 VDD1.n25 VDD1.n24 5.81868
R752 VDD1.n91 VDD1.n90 5.81868
R753 VDD1.n131 VDD1.n67 5.81868
R754 VDD1.n62 VDD1.n61 5.04292
R755 VDD1.n28 VDD1.n19 5.04292
R756 VDD1.n94 VDD1.n85 5.04292
R757 VDD1.n129 VDD1.n128 5.04292
R758 VDD1.n58 VDD1.n2 4.26717
R759 VDD1.n29 VDD1.n17 4.26717
R760 VDD1.n95 VDD1.n83 4.26717
R761 VDD1.n125 VDD1.n69 4.26717
R762 VDD1.n57 VDD1.n4 3.49141
R763 VDD1.n33 VDD1.n32 3.49141
R764 VDD1.n99 VDD1.n98 3.49141
R765 VDD1.n124 VDD1.n71 3.49141
R766 VDD1.n23 VDD1.n22 2.84303
R767 VDD1.n89 VDD1.n88 2.84303
R768 VDD1.n54 VDD1.n53 2.71565
R769 VDD1.n36 VDD1.n15 2.71565
R770 VDD1.n102 VDD1.n81 2.71565
R771 VDD1.n121 VDD1.n120 2.71565
R772 VDD1 VDD1.n137 2.28929
R773 VDD1.n50 VDD1.n6 1.93989
R774 VDD1.n37 VDD1.n13 1.93989
R775 VDD1.n103 VDD1.n79 1.93989
R776 VDD1.n117 VDD1.n73 1.93989
R777 VDD1.n136 VDD1.t5 1.62212
R778 VDD1.n136 VDD1.t0 1.62212
R779 VDD1.n65 VDD1.t3 1.62212
R780 VDD1.n65 VDD1.t9 1.62212
R781 VDD1.n134 VDD1.t7 1.62212
R782 VDD1.n134 VDD1.t8 1.62212
R783 VDD1.n132 VDD1.t1 1.62212
R784 VDD1.n132 VDD1.t4 1.62212
R785 VDD1.n49 VDD1.n8 1.16414
R786 VDD1.n41 VDD1.n40 1.16414
R787 VDD1.n108 VDD1.n106 1.16414
R788 VDD1.n116 VDD1.n75 1.16414
R789 VDD1 VDD1.n66 0.841017
R790 VDD1.n135 VDD1.n133 0.727482
R791 VDD1.n46 VDD1.n45 0.388379
R792 VDD1.n12 VDD1.n10 0.388379
R793 VDD1.n107 VDD1.n77 0.388379
R794 VDD1.n113 VDD1.n112 0.388379
R795 VDD1.n63 VDD1.n1 0.155672
R796 VDD1.n56 VDD1.n1 0.155672
R797 VDD1.n56 VDD1.n55 0.155672
R798 VDD1.n55 VDD1.n5 0.155672
R799 VDD1.n48 VDD1.n5 0.155672
R800 VDD1.n48 VDD1.n47 0.155672
R801 VDD1.n47 VDD1.n9 0.155672
R802 VDD1.n39 VDD1.n9 0.155672
R803 VDD1.n39 VDD1.n38 0.155672
R804 VDD1.n38 VDD1.n14 0.155672
R805 VDD1.n31 VDD1.n14 0.155672
R806 VDD1.n31 VDD1.n30 0.155672
R807 VDD1.n30 VDD1.n18 0.155672
R808 VDD1.n23 VDD1.n18 0.155672
R809 VDD1.n89 VDD1.n84 0.155672
R810 VDD1.n96 VDD1.n84 0.155672
R811 VDD1.n97 VDD1.n96 0.155672
R812 VDD1.n97 VDD1.n80 0.155672
R813 VDD1.n104 VDD1.n80 0.155672
R814 VDD1.n105 VDD1.n104 0.155672
R815 VDD1.n105 VDD1.n76 0.155672
R816 VDD1.n114 VDD1.n76 0.155672
R817 VDD1.n115 VDD1.n114 0.155672
R818 VDD1.n115 VDD1.n72 0.155672
R819 VDD1.n122 VDD1.n72 0.155672
R820 VDD1.n123 VDD1.n122 0.155672
R821 VDD1.n123 VDD1.n68 0.155672
R822 VDD1.n130 VDD1.n68 0.155672
R823 B.n1058 B.n1057 585
R824 B.n367 B.n178 585
R825 B.n366 B.n365 585
R826 B.n364 B.n363 585
R827 B.n362 B.n361 585
R828 B.n360 B.n359 585
R829 B.n358 B.n357 585
R830 B.n356 B.n355 585
R831 B.n354 B.n353 585
R832 B.n352 B.n351 585
R833 B.n350 B.n349 585
R834 B.n348 B.n347 585
R835 B.n346 B.n345 585
R836 B.n344 B.n343 585
R837 B.n342 B.n341 585
R838 B.n340 B.n339 585
R839 B.n338 B.n337 585
R840 B.n336 B.n335 585
R841 B.n334 B.n333 585
R842 B.n332 B.n331 585
R843 B.n330 B.n329 585
R844 B.n328 B.n327 585
R845 B.n326 B.n325 585
R846 B.n324 B.n323 585
R847 B.n322 B.n321 585
R848 B.n320 B.n319 585
R849 B.n318 B.n317 585
R850 B.n316 B.n315 585
R851 B.n314 B.n313 585
R852 B.n312 B.n311 585
R853 B.n310 B.n309 585
R854 B.n308 B.n307 585
R855 B.n306 B.n305 585
R856 B.n304 B.n303 585
R857 B.n302 B.n301 585
R858 B.n300 B.n299 585
R859 B.n298 B.n297 585
R860 B.n296 B.n295 585
R861 B.n294 B.n293 585
R862 B.n292 B.n291 585
R863 B.n290 B.n289 585
R864 B.n288 B.n287 585
R865 B.n286 B.n285 585
R866 B.n284 B.n283 585
R867 B.n282 B.n281 585
R868 B.n280 B.n279 585
R869 B.n278 B.n277 585
R870 B.n276 B.n275 585
R871 B.n274 B.n273 585
R872 B.n272 B.n271 585
R873 B.n270 B.n269 585
R874 B.n268 B.n267 585
R875 B.n266 B.n265 585
R876 B.n264 B.n263 585
R877 B.n262 B.n261 585
R878 B.n260 B.n259 585
R879 B.n258 B.n257 585
R880 B.n256 B.n255 585
R881 B.n254 B.n253 585
R882 B.n252 B.n251 585
R883 B.n250 B.n249 585
R884 B.n248 B.n247 585
R885 B.n246 B.n245 585
R886 B.n244 B.n243 585
R887 B.n242 B.n241 585
R888 B.n240 B.n239 585
R889 B.n238 B.n237 585
R890 B.n236 B.n235 585
R891 B.n234 B.n233 585
R892 B.n232 B.n231 585
R893 B.n230 B.n229 585
R894 B.n228 B.n227 585
R895 B.n226 B.n225 585
R896 B.n224 B.n223 585
R897 B.n222 B.n221 585
R898 B.n220 B.n219 585
R899 B.n218 B.n217 585
R900 B.n216 B.n215 585
R901 B.n214 B.n213 585
R902 B.n212 B.n211 585
R903 B.n210 B.n209 585
R904 B.n208 B.n207 585
R905 B.n206 B.n205 585
R906 B.n204 B.n203 585
R907 B.n202 B.n201 585
R908 B.n200 B.n199 585
R909 B.n198 B.n197 585
R910 B.n196 B.n195 585
R911 B.n194 B.n193 585
R912 B.n192 B.n191 585
R913 B.n190 B.n189 585
R914 B.n188 B.n187 585
R915 B.n186 B.n185 585
R916 B.n130 B.n129 585
R917 B.n1056 B.n131 585
R918 B.n1061 B.n131 585
R919 B.n1055 B.n1054 585
R920 B.n1054 B.n127 585
R921 B.n1053 B.n126 585
R922 B.n1067 B.n126 585
R923 B.n1052 B.n125 585
R924 B.n1068 B.n125 585
R925 B.n1051 B.n124 585
R926 B.n1069 B.n124 585
R927 B.n1050 B.n1049 585
R928 B.n1049 B.n120 585
R929 B.n1048 B.n119 585
R930 B.n1075 B.n119 585
R931 B.n1047 B.n118 585
R932 B.n1076 B.n118 585
R933 B.n1046 B.n117 585
R934 B.n1077 B.n117 585
R935 B.n1045 B.n1044 585
R936 B.n1044 B.n113 585
R937 B.n1043 B.n112 585
R938 B.n1083 B.n112 585
R939 B.n1042 B.n111 585
R940 B.n1084 B.n111 585
R941 B.n1041 B.n110 585
R942 B.n1085 B.n110 585
R943 B.n1040 B.n1039 585
R944 B.n1039 B.n106 585
R945 B.n1038 B.n105 585
R946 B.n1091 B.n105 585
R947 B.n1037 B.n104 585
R948 B.n1092 B.n104 585
R949 B.n1036 B.n103 585
R950 B.n1093 B.n103 585
R951 B.n1035 B.n1034 585
R952 B.n1034 B.n99 585
R953 B.n1033 B.n98 585
R954 B.n1099 B.n98 585
R955 B.n1032 B.n97 585
R956 B.n1100 B.n97 585
R957 B.n1031 B.n96 585
R958 B.n1101 B.n96 585
R959 B.n1030 B.n1029 585
R960 B.n1029 B.n92 585
R961 B.n1028 B.n91 585
R962 B.n1107 B.n91 585
R963 B.n1027 B.n90 585
R964 B.n1108 B.n90 585
R965 B.n1026 B.n89 585
R966 B.n1109 B.n89 585
R967 B.n1025 B.n1024 585
R968 B.n1024 B.n85 585
R969 B.n1023 B.n84 585
R970 B.n1115 B.n84 585
R971 B.n1022 B.n83 585
R972 B.n1116 B.n83 585
R973 B.n1021 B.n82 585
R974 B.n1117 B.n82 585
R975 B.n1020 B.n1019 585
R976 B.n1019 B.n78 585
R977 B.n1018 B.n77 585
R978 B.n1123 B.n77 585
R979 B.n1017 B.n76 585
R980 B.n1124 B.n76 585
R981 B.n1016 B.n75 585
R982 B.n1125 B.n75 585
R983 B.n1015 B.n1014 585
R984 B.n1014 B.n74 585
R985 B.n1013 B.n70 585
R986 B.n1131 B.n70 585
R987 B.n1012 B.n69 585
R988 B.n1132 B.n69 585
R989 B.n1011 B.n68 585
R990 B.n1133 B.n68 585
R991 B.n1010 B.n1009 585
R992 B.n1009 B.n64 585
R993 B.n1008 B.n63 585
R994 B.n1139 B.n63 585
R995 B.n1007 B.n62 585
R996 B.n1140 B.n62 585
R997 B.n1006 B.n61 585
R998 B.n1141 B.n61 585
R999 B.n1005 B.n1004 585
R1000 B.n1004 B.n57 585
R1001 B.n1003 B.n56 585
R1002 B.n1147 B.n56 585
R1003 B.n1002 B.n55 585
R1004 B.n1148 B.n55 585
R1005 B.n1001 B.n54 585
R1006 B.n1149 B.n54 585
R1007 B.n1000 B.n999 585
R1008 B.n999 B.n50 585
R1009 B.n998 B.n49 585
R1010 B.n1155 B.n49 585
R1011 B.n997 B.n48 585
R1012 B.n1156 B.n48 585
R1013 B.n996 B.n47 585
R1014 B.n1157 B.n47 585
R1015 B.n995 B.n994 585
R1016 B.n994 B.n43 585
R1017 B.n993 B.n42 585
R1018 B.n1163 B.n42 585
R1019 B.n992 B.n41 585
R1020 B.n1164 B.n41 585
R1021 B.n991 B.n40 585
R1022 B.n1165 B.n40 585
R1023 B.n990 B.n989 585
R1024 B.n989 B.n36 585
R1025 B.n988 B.n35 585
R1026 B.n1171 B.n35 585
R1027 B.n987 B.n34 585
R1028 B.n1172 B.n34 585
R1029 B.n986 B.n33 585
R1030 B.n1173 B.n33 585
R1031 B.n985 B.n984 585
R1032 B.n984 B.n29 585
R1033 B.n983 B.n28 585
R1034 B.n1179 B.n28 585
R1035 B.n982 B.n27 585
R1036 B.n1180 B.n27 585
R1037 B.n981 B.n26 585
R1038 B.n1181 B.n26 585
R1039 B.n980 B.n979 585
R1040 B.n979 B.n22 585
R1041 B.n978 B.n21 585
R1042 B.n1187 B.n21 585
R1043 B.n977 B.n20 585
R1044 B.n1188 B.n20 585
R1045 B.n976 B.n19 585
R1046 B.n1189 B.n19 585
R1047 B.n975 B.n974 585
R1048 B.n974 B.n18 585
R1049 B.n973 B.n14 585
R1050 B.n1195 B.n14 585
R1051 B.n972 B.n13 585
R1052 B.n1196 B.n13 585
R1053 B.n971 B.n12 585
R1054 B.n1197 B.n12 585
R1055 B.n970 B.n969 585
R1056 B.n969 B.n8 585
R1057 B.n968 B.n7 585
R1058 B.n1203 B.n7 585
R1059 B.n967 B.n6 585
R1060 B.n1204 B.n6 585
R1061 B.n966 B.n5 585
R1062 B.n1205 B.n5 585
R1063 B.n965 B.n964 585
R1064 B.n964 B.n4 585
R1065 B.n963 B.n368 585
R1066 B.n963 B.n962 585
R1067 B.n953 B.n369 585
R1068 B.n370 B.n369 585
R1069 B.n955 B.n954 585
R1070 B.n956 B.n955 585
R1071 B.n952 B.n375 585
R1072 B.n375 B.n374 585
R1073 B.n951 B.n950 585
R1074 B.n950 B.n949 585
R1075 B.n377 B.n376 585
R1076 B.n942 B.n377 585
R1077 B.n941 B.n940 585
R1078 B.n943 B.n941 585
R1079 B.n939 B.n382 585
R1080 B.n382 B.n381 585
R1081 B.n938 B.n937 585
R1082 B.n937 B.n936 585
R1083 B.n384 B.n383 585
R1084 B.n385 B.n384 585
R1085 B.n929 B.n928 585
R1086 B.n930 B.n929 585
R1087 B.n927 B.n390 585
R1088 B.n390 B.n389 585
R1089 B.n926 B.n925 585
R1090 B.n925 B.n924 585
R1091 B.n392 B.n391 585
R1092 B.n393 B.n392 585
R1093 B.n917 B.n916 585
R1094 B.n918 B.n917 585
R1095 B.n915 B.n398 585
R1096 B.n398 B.n397 585
R1097 B.n914 B.n913 585
R1098 B.n913 B.n912 585
R1099 B.n400 B.n399 585
R1100 B.n401 B.n400 585
R1101 B.n905 B.n904 585
R1102 B.n906 B.n905 585
R1103 B.n903 B.n406 585
R1104 B.n406 B.n405 585
R1105 B.n902 B.n901 585
R1106 B.n901 B.n900 585
R1107 B.n408 B.n407 585
R1108 B.n409 B.n408 585
R1109 B.n893 B.n892 585
R1110 B.n894 B.n893 585
R1111 B.n891 B.n414 585
R1112 B.n414 B.n413 585
R1113 B.n890 B.n889 585
R1114 B.n889 B.n888 585
R1115 B.n416 B.n415 585
R1116 B.n417 B.n416 585
R1117 B.n881 B.n880 585
R1118 B.n882 B.n881 585
R1119 B.n879 B.n421 585
R1120 B.n425 B.n421 585
R1121 B.n878 B.n877 585
R1122 B.n877 B.n876 585
R1123 B.n423 B.n422 585
R1124 B.n424 B.n423 585
R1125 B.n869 B.n868 585
R1126 B.n870 B.n869 585
R1127 B.n867 B.n430 585
R1128 B.n430 B.n429 585
R1129 B.n866 B.n865 585
R1130 B.n865 B.n864 585
R1131 B.n432 B.n431 585
R1132 B.n433 B.n432 585
R1133 B.n857 B.n856 585
R1134 B.n858 B.n857 585
R1135 B.n855 B.n438 585
R1136 B.n438 B.n437 585
R1137 B.n854 B.n853 585
R1138 B.n853 B.n852 585
R1139 B.n440 B.n439 585
R1140 B.n845 B.n440 585
R1141 B.n844 B.n843 585
R1142 B.n846 B.n844 585
R1143 B.n842 B.n445 585
R1144 B.n445 B.n444 585
R1145 B.n841 B.n840 585
R1146 B.n840 B.n839 585
R1147 B.n447 B.n446 585
R1148 B.n448 B.n447 585
R1149 B.n832 B.n831 585
R1150 B.n833 B.n832 585
R1151 B.n830 B.n453 585
R1152 B.n453 B.n452 585
R1153 B.n829 B.n828 585
R1154 B.n828 B.n827 585
R1155 B.n455 B.n454 585
R1156 B.n456 B.n455 585
R1157 B.n820 B.n819 585
R1158 B.n821 B.n820 585
R1159 B.n818 B.n461 585
R1160 B.n461 B.n460 585
R1161 B.n817 B.n816 585
R1162 B.n816 B.n815 585
R1163 B.n463 B.n462 585
R1164 B.n464 B.n463 585
R1165 B.n808 B.n807 585
R1166 B.n809 B.n808 585
R1167 B.n806 B.n469 585
R1168 B.n469 B.n468 585
R1169 B.n805 B.n804 585
R1170 B.n804 B.n803 585
R1171 B.n471 B.n470 585
R1172 B.n472 B.n471 585
R1173 B.n796 B.n795 585
R1174 B.n797 B.n796 585
R1175 B.n794 B.n477 585
R1176 B.n477 B.n476 585
R1177 B.n793 B.n792 585
R1178 B.n792 B.n791 585
R1179 B.n479 B.n478 585
R1180 B.n480 B.n479 585
R1181 B.n784 B.n783 585
R1182 B.n785 B.n784 585
R1183 B.n782 B.n485 585
R1184 B.n485 B.n484 585
R1185 B.n781 B.n780 585
R1186 B.n780 B.n779 585
R1187 B.n487 B.n486 585
R1188 B.n488 B.n487 585
R1189 B.n772 B.n771 585
R1190 B.n773 B.n772 585
R1191 B.n770 B.n493 585
R1192 B.n493 B.n492 585
R1193 B.n769 B.n768 585
R1194 B.n768 B.n767 585
R1195 B.n495 B.n494 585
R1196 B.n496 B.n495 585
R1197 B.n760 B.n759 585
R1198 B.n761 B.n760 585
R1199 B.n758 B.n501 585
R1200 B.n501 B.n500 585
R1201 B.n757 B.n756 585
R1202 B.n756 B.n755 585
R1203 B.n503 B.n502 585
R1204 B.n504 B.n503 585
R1205 B.n748 B.n747 585
R1206 B.n749 B.n748 585
R1207 B.n507 B.n506 585
R1208 B.n560 B.n558 585
R1209 B.n561 B.n557 585
R1210 B.n561 B.n508 585
R1211 B.n564 B.n563 585
R1212 B.n565 B.n556 585
R1213 B.n567 B.n566 585
R1214 B.n569 B.n555 585
R1215 B.n572 B.n571 585
R1216 B.n573 B.n554 585
R1217 B.n575 B.n574 585
R1218 B.n577 B.n553 585
R1219 B.n580 B.n579 585
R1220 B.n581 B.n552 585
R1221 B.n583 B.n582 585
R1222 B.n585 B.n551 585
R1223 B.n588 B.n587 585
R1224 B.n589 B.n550 585
R1225 B.n591 B.n590 585
R1226 B.n593 B.n549 585
R1227 B.n596 B.n595 585
R1228 B.n597 B.n548 585
R1229 B.n599 B.n598 585
R1230 B.n601 B.n547 585
R1231 B.n604 B.n603 585
R1232 B.n605 B.n546 585
R1233 B.n607 B.n606 585
R1234 B.n609 B.n545 585
R1235 B.n612 B.n611 585
R1236 B.n613 B.n544 585
R1237 B.n615 B.n614 585
R1238 B.n617 B.n543 585
R1239 B.n620 B.n619 585
R1240 B.n621 B.n542 585
R1241 B.n623 B.n622 585
R1242 B.n625 B.n541 585
R1243 B.n628 B.n627 585
R1244 B.n629 B.n540 585
R1245 B.n631 B.n630 585
R1246 B.n633 B.n539 585
R1247 B.n636 B.n635 585
R1248 B.n637 B.n538 585
R1249 B.n642 B.n641 585
R1250 B.n644 B.n537 585
R1251 B.n647 B.n646 585
R1252 B.n648 B.n536 585
R1253 B.n650 B.n649 585
R1254 B.n652 B.n535 585
R1255 B.n655 B.n654 585
R1256 B.n656 B.n534 585
R1257 B.n658 B.n657 585
R1258 B.n660 B.n533 585
R1259 B.n663 B.n662 585
R1260 B.n665 B.n530 585
R1261 B.n667 B.n666 585
R1262 B.n669 B.n529 585
R1263 B.n672 B.n671 585
R1264 B.n673 B.n528 585
R1265 B.n675 B.n674 585
R1266 B.n677 B.n527 585
R1267 B.n680 B.n679 585
R1268 B.n681 B.n526 585
R1269 B.n683 B.n682 585
R1270 B.n685 B.n525 585
R1271 B.n688 B.n687 585
R1272 B.n689 B.n524 585
R1273 B.n691 B.n690 585
R1274 B.n693 B.n523 585
R1275 B.n696 B.n695 585
R1276 B.n697 B.n522 585
R1277 B.n699 B.n698 585
R1278 B.n701 B.n521 585
R1279 B.n704 B.n703 585
R1280 B.n705 B.n520 585
R1281 B.n707 B.n706 585
R1282 B.n709 B.n519 585
R1283 B.n712 B.n711 585
R1284 B.n713 B.n518 585
R1285 B.n715 B.n714 585
R1286 B.n717 B.n517 585
R1287 B.n720 B.n719 585
R1288 B.n721 B.n516 585
R1289 B.n723 B.n722 585
R1290 B.n725 B.n515 585
R1291 B.n728 B.n727 585
R1292 B.n729 B.n514 585
R1293 B.n731 B.n730 585
R1294 B.n733 B.n513 585
R1295 B.n736 B.n735 585
R1296 B.n737 B.n512 585
R1297 B.n739 B.n738 585
R1298 B.n741 B.n511 585
R1299 B.n742 B.n510 585
R1300 B.n745 B.n744 585
R1301 B.n746 B.n509 585
R1302 B.n509 B.n508 585
R1303 B.n751 B.n750 585
R1304 B.n750 B.n749 585
R1305 B.n752 B.n505 585
R1306 B.n505 B.n504 585
R1307 B.n754 B.n753 585
R1308 B.n755 B.n754 585
R1309 B.n499 B.n498 585
R1310 B.n500 B.n499 585
R1311 B.n763 B.n762 585
R1312 B.n762 B.n761 585
R1313 B.n764 B.n497 585
R1314 B.n497 B.n496 585
R1315 B.n766 B.n765 585
R1316 B.n767 B.n766 585
R1317 B.n491 B.n490 585
R1318 B.n492 B.n491 585
R1319 B.n775 B.n774 585
R1320 B.n774 B.n773 585
R1321 B.n776 B.n489 585
R1322 B.n489 B.n488 585
R1323 B.n778 B.n777 585
R1324 B.n779 B.n778 585
R1325 B.n483 B.n482 585
R1326 B.n484 B.n483 585
R1327 B.n787 B.n786 585
R1328 B.n786 B.n785 585
R1329 B.n788 B.n481 585
R1330 B.n481 B.n480 585
R1331 B.n790 B.n789 585
R1332 B.n791 B.n790 585
R1333 B.n475 B.n474 585
R1334 B.n476 B.n475 585
R1335 B.n799 B.n798 585
R1336 B.n798 B.n797 585
R1337 B.n800 B.n473 585
R1338 B.n473 B.n472 585
R1339 B.n802 B.n801 585
R1340 B.n803 B.n802 585
R1341 B.n467 B.n466 585
R1342 B.n468 B.n467 585
R1343 B.n811 B.n810 585
R1344 B.n810 B.n809 585
R1345 B.n812 B.n465 585
R1346 B.n465 B.n464 585
R1347 B.n814 B.n813 585
R1348 B.n815 B.n814 585
R1349 B.n459 B.n458 585
R1350 B.n460 B.n459 585
R1351 B.n823 B.n822 585
R1352 B.n822 B.n821 585
R1353 B.n824 B.n457 585
R1354 B.n457 B.n456 585
R1355 B.n826 B.n825 585
R1356 B.n827 B.n826 585
R1357 B.n451 B.n450 585
R1358 B.n452 B.n451 585
R1359 B.n835 B.n834 585
R1360 B.n834 B.n833 585
R1361 B.n836 B.n449 585
R1362 B.n449 B.n448 585
R1363 B.n838 B.n837 585
R1364 B.n839 B.n838 585
R1365 B.n443 B.n442 585
R1366 B.n444 B.n443 585
R1367 B.n848 B.n847 585
R1368 B.n847 B.n846 585
R1369 B.n849 B.n441 585
R1370 B.n845 B.n441 585
R1371 B.n851 B.n850 585
R1372 B.n852 B.n851 585
R1373 B.n436 B.n435 585
R1374 B.n437 B.n436 585
R1375 B.n860 B.n859 585
R1376 B.n859 B.n858 585
R1377 B.n861 B.n434 585
R1378 B.n434 B.n433 585
R1379 B.n863 B.n862 585
R1380 B.n864 B.n863 585
R1381 B.n428 B.n427 585
R1382 B.n429 B.n428 585
R1383 B.n872 B.n871 585
R1384 B.n871 B.n870 585
R1385 B.n873 B.n426 585
R1386 B.n426 B.n424 585
R1387 B.n875 B.n874 585
R1388 B.n876 B.n875 585
R1389 B.n420 B.n419 585
R1390 B.n425 B.n420 585
R1391 B.n884 B.n883 585
R1392 B.n883 B.n882 585
R1393 B.n885 B.n418 585
R1394 B.n418 B.n417 585
R1395 B.n887 B.n886 585
R1396 B.n888 B.n887 585
R1397 B.n412 B.n411 585
R1398 B.n413 B.n412 585
R1399 B.n896 B.n895 585
R1400 B.n895 B.n894 585
R1401 B.n897 B.n410 585
R1402 B.n410 B.n409 585
R1403 B.n899 B.n898 585
R1404 B.n900 B.n899 585
R1405 B.n404 B.n403 585
R1406 B.n405 B.n404 585
R1407 B.n908 B.n907 585
R1408 B.n907 B.n906 585
R1409 B.n909 B.n402 585
R1410 B.n402 B.n401 585
R1411 B.n911 B.n910 585
R1412 B.n912 B.n911 585
R1413 B.n396 B.n395 585
R1414 B.n397 B.n396 585
R1415 B.n920 B.n919 585
R1416 B.n919 B.n918 585
R1417 B.n921 B.n394 585
R1418 B.n394 B.n393 585
R1419 B.n923 B.n922 585
R1420 B.n924 B.n923 585
R1421 B.n388 B.n387 585
R1422 B.n389 B.n388 585
R1423 B.n932 B.n931 585
R1424 B.n931 B.n930 585
R1425 B.n933 B.n386 585
R1426 B.n386 B.n385 585
R1427 B.n935 B.n934 585
R1428 B.n936 B.n935 585
R1429 B.n380 B.n379 585
R1430 B.n381 B.n380 585
R1431 B.n945 B.n944 585
R1432 B.n944 B.n943 585
R1433 B.n946 B.n378 585
R1434 B.n942 B.n378 585
R1435 B.n948 B.n947 585
R1436 B.n949 B.n948 585
R1437 B.n373 B.n372 585
R1438 B.n374 B.n373 585
R1439 B.n958 B.n957 585
R1440 B.n957 B.n956 585
R1441 B.n959 B.n371 585
R1442 B.n371 B.n370 585
R1443 B.n961 B.n960 585
R1444 B.n962 B.n961 585
R1445 B.n2 B.n0 585
R1446 B.n4 B.n2 585
R1447 B.n3 B.n1 585
R1448 B.n1204 B.n3 585
R1449 B.n1202 B.n1201 585
R1450 B.n1203 B.n1202 585
R1451 B.n1200 B.n9 585
R1452 B.n9 B.n8 585
R1453 B.n1199 B.n1198 585
R1454 B.n1198 B.n1197 585
R1455 B.n11 B.n10 585
R1456 B.n1196 B.n11 585
R1457 B.n1194 B.n1193 585
R1458 B.n1195 B.n1194 585
R1459 B.n1192 B.n15 585
R1460 B.n18 B.n15 585
R1461 B.n1191 B.n1190 585
R1462 B.n1190 B.n1189 585
R1463 B.n17 B.n16 585
R1464 B.n1188 B.n17 585
R1465 B.n1186 B.n1185 585
R1466 B.n1187 B.n1186 585
R1467 B.n1184 B.n23 585
R1468 B.n23 B.n22 585
R1469 B.n1183 B.n1182 585
R1470 B.n1182 B.n1181 585
R1471 B.n25 B.n24 585
R1472 B.n1180 B.n25 585
R1473 B.n1178 B.n1177 585
R1474 B.n1179 B.n1178 585
R1475 B.n1176 B.n30 585
R1476 B.n30 B.n29 585
R1477 B.n1175 B.n1174 585
R1478 B.n1174 B.n1173 585
R1479 B.n32 B.n31 585
R1480 B.n1172 B.n32 585
R1481 B.n1170 B.n1169 585
R1482 B.n1171 B.n1170 585
R1483 B.n1168 B.n37 585
R1484 B.n37 B.n36 585
R1485 B.n1167 B.n1166 585
R1486 B.n1166 B.n1165 585
R1487 B.n39 B.n38 585
R1488 B.n1164 B.n39 585
R1489 B.n1162 B.n1161 585
R1490 B.n1163 B.n1162 585
R1491 B.n1160 B.n44 585
R1492 B.n44 B.n43 585
R1493 B.n1159 B.n1158 585
R1494 B.n1158 B.n1157 585
R1495 B.n46 B.n45 585
R1496 B.n1156 B.n46 585
R1497 B.n1154 B.n1153 585
R1498 B.n1155 B.n1154 585
R1499 B.n1152 B.n51 585
R1500 B.n51 B.n50 585
R1501 B.n1151 B.n1150 585
R1502 B.n1150 B.n1149 585
R1503 B.n53 B.n52 585
R1504 B.n1148 B.n53 585
R1505 B.n1146 B.n1145 585
R1506 B.n1147 B.n1146 585
R1507 B.n1144 B.n58 585
R1508 B.n58 B.n57 585
R1509 B.n1143 B.n1142 585
R1510 B.n1142 B.n1141 585
R1511 B.n60 B.n59 585
R1512 B.n1140 B.n60 585
R1513 B.n1138 B.n1137 585
R1514 B.n1139 B.n1138 585
R1515 B.n1136 B.n65 585
R1516 B.n65 B.n64 585
R1517 B.n1135 B.n1134 585
R1518 B.n1134 B.n1133 585
R1519 B.n67 B.n66 585
R1520 B.n1132 B.n67 585
R1521 B.n1130 B.n1129 585
R1522 B.n1131 B.n1130 585
R1523 B.n1128 B.n71 585
R1524 B.n74 B.n71 585
R1525 B.n1127 B.n1126 585
R1526 B.n1126 B.n1125 585
R1527 B.n73 B.n72 585
R1528 B.n1124 B.n73 585
R1529 B.n1122 B.n1121 585
R1530 B.n1123 B.n1122 585
R1531 B.n1120 B.n79 585
R1532 B.n79 B.n78 585
R1533 B.n1119 B.n1118 585
R1534 B.n1118 B.n1117 585
R1535 B.n81 B.n80 585
R1536 B.n1116 B.n81 585
R1537 B.n1114 B.n1113 585
R1538 B.n1115 B.n1114 585
R1539 B.n1112 B.n86 585
R1540 B.n86 B.n85 585
R1541 B.n1111 B.n1110 585
R1542 B.n1110 B.n1109 585
R1543 B.n88 B.n87 585
R1544 B.n1108 B.n88 585
R1545 B.n1106 B.n1105 585
R1546 B.n1107 B.n1106 585
R1547 B.n1104 B.n93 585
R1548 B.n93 B.n92 585
R1549 B.n1103 B.n1102 585
R1550 B.n1102 B.n1101 585
R1551 B.n95 B.n94 585
R1552 B.n1100 B.n95 585
R1553 B.n1098 B.n1097 585
R1554 B.n1099 B.n1098 585
R1555 B.n1096 B.n100 585
R1556 B.n100 B.n99 585
R1557 B.n1095 B.n1094 585
R1558 B.n1094 B.n1093 585
R1559 B.n102 B.n101 585
R1560 B.n1092 B.n102 585
R1561 B.n1090 B.n1089 585
R1562 B.n1091 B.n1090 585
R1563 B.n1088 B.n107 585
R1564 B.n107 B.n106 585
R1565 B.n1087 B.n1086 585
R1566 B.n1086 B.n1085 585
R1567 B.n109 B.n108 585
R1568 B.n1084 B.n109 585
R1569 B.n1082 B.n1081 585
R1570 B.n1083 B.n1082 585
R1571 B.n1080 B.n114 585
R1572 B.n114 B.n113 585
R1573 B.n1079 B.n1078 585
R1574 B.n1078 B.n1077 585
R1575 B.n116 B.n115 585
R1576 B.n1076 B.n116 585
R1577 B.n1074 B.n1073 585
R1578 B.n1075 B.n1074 585
R1579 B.n1072 B.n121 585
R1580 B.n121 B.n120 585
R1581 B.n1071 B.n1070 585
R1582 B.n1070 B.n1069 585
R1583 B.n123 B.n122 585
R1584 B.n1068 B.n123 585
R1585 B.n1066 B.n1065 585
R1586 B.n1067 B.n1066 585
R1587 B.n1064 B.n128 585
R1588 B.n128 B.n127 585
R1589 B.n1063 B.n1062 585
R1590 B.n1062 B.n1061 585
R1591 B.n1207 B.n1206 585
R1592 B.n1206 B.n1205 585
R1593 B.n750 B.n507 530.939
R1594 B.n1062 B.n130 530.939
R1595 B.n748 B.n509 530.939
R1596 B.n1058 B.n131 530.939
R1597 B.n531 B.t17 356.481
R1598 B.n638 B.t23 356.481
R1599 B.n182 B.t12 356.481
R1600 B.n179 B.t19 356.481
R1601 B.n531 B.t14 298.075
R1602 B.n638 B.t21 298.075
R1603 B.n182 B.t10 298.075
R1604 B.n179 B.t18 298.075
R1605 B.n532 B.t16 286.08
R1606 B.n180 B.t20 286.08
R1607 B.n639 B.t22 286.08
R1608 B.n183 B.t13 286.08
R1609 B.n1060 B.n1059 256.663
R1610 B.n1060 B.n177 256.663
R1611 B.n1060 B.n176 256.663
R1612 B.n1060 B.n175 256.663
R1613 B.n1060 B.n174 256.663
R1614 B.n1060 B.n173 256.663
R1615 B.n1060 B.n172 256.663
R1616 B.n1060 B.n171 256.663
R1617 B.n1060 B.n170 256.663
R1618 B.n1060 B.n169 256.663
R1619 B.n1060 B.n168 256.663
R1620 B.n1060 B.n167 256.663
R1621 B.n1060 B.n166 256.663
R1622 B.n1060 B.n165 256.663
R1623 B.n1060 B.n164 256.663
R1624 B.n1060 B.n163 256.663
R1625 B.n1060 B.n162 256.663
R1626 B.n1060 B.n161 256.663
R1627 B.n1060 B.n160 256.663
R1628 B.n1060 B.n159 256.663
R1629 B.n1060 B.n158 256.663
R1630 B.n1060 B.n157 256.663
R1631 B.n1060 B.n156 256.663
R1632 B.n1060 B.n155 256.663
R1633 B.n1060 B.n154 256.663
R1634 B.n1060 B.n153 256.663
R1635 B.n1060 B.n152 256.663
R1636 B.n1060 B.n151 256.663
R1637 B.n1060 B.n150 256.663
R1638 B.n1060 B.n149 256.663
R1639 B.n1060 B.n148 256.663
R1640 B.n1060 B.n147 256.663
R1641 B.n1060 B.n146 256.663
R1642 B.n1060 B.n145 256.663
R1643 B.n1060 B.n144 256.663
R1644 B.n1060 B.n143 256.663
R1645 B.n1060 B.n142 256.663
R1646 B.n1060 B.n141 256.663
R1647 B.n1060 B.n140 256.663
R1648 B.n1060 B.n139 256.663
R1649 B.n1060 B.n138 256.663
R1650 B.n1060 B.n137 256.663
R1651 B.n1060 B.n136 256.663
R1652 B.n1060 B.n135 256.663
R1653 B.n1060 B.n134 256.663
R1654 B.n1060 B.n133 256.663
R1655 B.n1060 B.n132 256.663
R1656 B.n559 B.n508 256.663
R1657 B.n562 B.n508 256.663
R1658 B.n568 B.n508 256.663
R1659 B.n570 B.n508 256.663
R1660 B.n576 B.n508 256.663
R1661 B.n578 B.n508 256.663
R1662 B.n584 B.n508 256.663
R1663 B.n586 B.n508 256.663
R1664 B.n592 B.n508 256.663
R1665 B.n594 B.n508 256.663
R1666 B.n600 B.n508 256.663
R1667 B.n602 B.n508 256.663
R1668 B.n608 B.n508 256.663
R1669 B.n610 B.n508 256.663
R1670 B.n616 B.n508 256.663
R1671 B.n618 B.n508 256.663
R1672 B.n624 B.n508 256.663
R1673 B.n626 B.n508 256.663
R1674 B.n632 B.n508 256.663
R1675 B.n634 B.n508 256.663
R1676 B.n643 B.n508 256.663
R1677 B.n645 B.n508 256.663
R1678 B.n651 B.n508 256.663
R1679 B.n653 B.n508 256.663
R1680 B.n659 B.n508 256.663
R1681 B.n661 B.n508 256.663
R1682 B.n668 B.n508 256.663
R1683 B.n670 B.n508 256.663
R1684 B.n676 B.n508 256.663
R1685 B.n678 B.n508 256.663
R1686 B.n684 B.n508 256.663
R1687 B.n686 B.n508 256.663
R1688 B.n692 B.n508 256.663
R1689 B.n694 B.n508 256.663
R1690 B.n700 B.n508 256.663
R1691 B.n702 B.n508 256.663
R1692 B.n708 B.n508 256.663
R1693 B.n710 B.n508 256.663
R1694 B.n716 B.n508 256.663
R1695 B.n718 B.n508 256.663
R1696 B.n724 B.n508 256.663
R1697 B.n726 B.n508 256.663
R1698 B.n732 B.n508 256.663
R1699 B.n734 B.n508 256.663
R1700 B.n740 B.n508 256.663
R1701 B.n743 B.n508 256.663
R1702 B.n750 B.n505 163.367
R1703 B.n754 B.n505 163.367
R1704 B.n754 B.n499 163.367
R1705 B.n762 B.n499 163.367
R1706 B.n762 B.n497 163.367
R1707 B.n766 B.n497 163.367
R1708 B.n766 B.n491 163.367
R1709 B.n774 B.n491 163.367
R1710 B.n774 B.n489 163.367
R1711 B.n778 B.n489 163.367
R1712 B.n778 B.n483 163.367
R1713 B.n786 B.n483 163.367
R1714 B.n786 B.n481 163.367
R1715 B.n790 B.n481 163.367
R1716 B.n790 B.n475 163.367
R1717 B.n798 B.n475 163.367
R1718 B.n798 B.n473 163.367
R1719 B.n802 B.n473 163.367
R1720 B.n802 B.n467 163.367
R1721 B.n810 B.n467 163.367
R1722 B.n810 B.n465 163.367
R1723 B.n814 B.n465 163.367
R1724 B.n814 B.n459 163.367
R1725 B.n822 B.n459 163.367
R1726 B.n822 B.n457 163.367
R1727 B.n826 B.n457 163.367
R1728 B.n826 B.n451 163.367
R1729 B.n834 B.n451 163.367
R1730 B.n834 B.n449 163.367
R1731 B.n838 B.n449 163.367
R1732 B.n838 B.n443 163.367
R1733 B.n847 B.n443 163.367
R1734 B.n847 B.n441 163.367
R1735 B.n851 B.n441 163.367
R1736 B.n851 B.n436 163.367
R1737 B.n859 B.n436 163.367
R1738 B.n859 B.n434 163.367
R1739 B.n863 B.n434 163.367
R1740 B.n863 B.n428 163.367
R1741 B.n871 B.n428 163.367
R1742 B.n871 B.n426 163.367
R1743 B.n875 B.n426 163.367
R1744 B.n875 B.n420 163.367
R1745 B.n883 B.n420 163.367
R1746 B.n883 B.n418 163.367
R1747 B.n887 B.n418 163.367
R1748 B.n887 B.n412 163.367
R1749 B.n895 B.n412 163.367
R1750 B.n895 B.n410 163.367
R1751 B.n899 B.n410 163.367
R1752 B.n899 B.n404 163.367
R1753 B.n907 B.n404 163.367
R1754 B.n907 B.n402 163.367
R1755 B.n911 B.n402 163.367
R1756 B.n911 B.n396 163.367
R1757 B.n919 B.n396 163.367
R1758 B.n919 B.n394 163.367
R1759 B.n923 B.n394 163.367
R1760 B.n923 B.n388 163.367
R1761 B.n931 B.n388 163.367
R1762 B.n931 B.n386 163.367
R1763 B.n935 B.n386 163.367
R1764 B.n935 B.n380 163.367
R1765 B.n944 B.n380 163.367
R1766 B.n944 B.n378 163.367
R1767 B.n948 B.n378 163.367
R1768 B.n948 B.n373 163.367
R1769 B.n957 B.n373 163.367
R1770 B.n957 B.n371 163.367
R1771 B.n961 B.n371 163.367
R1772 B.n961 B.n2 163.367
R1773 B.n1206 B.n2 163.367
R1774 B.n1206 B.n3 163.367
R1775 B.n1202 B.n3 163.367
R1776 B.n1202 B.n9 163.367
R1777 B.n1198 B.n9 163.367
R1778 B.n1198 B.n11 163.367
R1779 B.n1194 B.n11 163.367
R1780 B.n1194 B.n15 163.367
R1781 B.n1190 B.n15 163.367
R1782 B.n1190 B.n17 163.367
R1783 B.n1186 B.n17 163.367
R1784 B.n1186 B.n23 163.367
R1785 B.n1182 B.n23 163.367
R1786 B.n1182 B.n25 163.367
R1787 B.n1178 B.n25 163.367
R1788 B.n1178 B.n30 163.367
R1789 B.n1174 B.n30 163.367
R1790 B.n1174 B.n32 163.367
R1791 B.n1170 B.n32 163.367
R1792 B.n1170 B.n37 163.367
R1793 B.n1166 B.n37 163.367
R1794 B.n1166 B.n39 163.367
R1795 B.n1162 B.n39 163.367
R1796 B.n1162 B.n44 163.367
R1797 B.n1158 B.n44 163.367
R1798 B.n1158 B.n46 163.367
R1799 B.n1154 B.n46 163.367
R1800 B.n1154 B.n51 163.367
R1801 B.n1150 B.n51 163.367
R1802 B.n1150 B.n53 163.367
R1803 B.n1146 B.n53 163.367
R1804 B.n1146 B.n58 163.367
R1805 B.n1142 B.n58 163.367
R1806 B.n1142 B.n60 163.367
R1807 B.n1138 B.n60 163.367
R1808 B.n1138 B.n65 163.367
R1809 B.n1134 B.n65 163.367
R1810 B.n1134 B.n67 163.367
R1811 B.n1130 B.n67 163.367
R1812 B.n1130 B.n71 163.367
R1813 B.n1126 B.n71 163.367
R1814 B.n1126 B.n73 163.367
R1815 B.n1122 B.n73 163.367
R1816 B.n1122 B.n79 163.367
R1817 B.n1118 B.n79 163.367
R1818 B.n1118 B.n81 163.367
R1819 B.n1114 B.n81 163.367
R1820 B.n1114 B.n86 163.367
R1821 B.n1110 B.n86 163.367
R1822 B.n1110 B.n88 163.367
R1823 B.n1106 B.n88 163.367
R1824 B.n1106 B.n93 163.367
R1825 B.n1102 B.n93 163.367
R1826 B.n1102 B.n95 163.367
R1827 B.n1098 B.n95 163.367
R1828 B.n1098 B.n100 163.367
R1829 B.n1094 B.n100 163.367
R1830 B.n1094 B.n102 163.367
R1831 B.n1090 B.n102 163.367
R1832 B.n1090 B.n107 163.367
R1833 B.n1086 B.n107 163.367
R1834 B.n1086 B.n109 163.367
R1835 B.n1082 B.n109 163.367
R1836 B.n1082 B.n114 163.367
R1837 B.n1078 B.n114 163.367
R1838 B.n1078 B.n116 163.367
R1839 B.n1074 B.n116 163.367
R1840 B.n1074 B.n121 163.367
R1841 B.n1070 B.n121 163.367
R1842 B.n1070 B.n123 163.367
R1843 B.n1066 B.n123 163.367
R1844 B.n1066 B.n128 163.367
R1845 B.n1062 B.n128 163.367
R1846 B.n561 B.n560 163.367
R1847 B.n563 B.n561 163.367
R1848 B.n567 B.n556 163.367
R1849 B.n571 B.n569 163.367
R1850 B.n575 B.n554 163.367
R1851 B.n579 B.n577 163.367
R1852 B.n583 B.n552 163.367
R1853 B.n587 B.n585 163.367
R1854 B.n591 B.n550 163.367
R1855 B.n595 B.n593 163.367
R1856 B.n599 B.n548 163.367
R1857 B.n603 B.n601 163.367
R1858 B.n607 B.n546 163.367
R1859 B.n611 B.n609 163.367
R1860 B.n615 B.n544 163.367
R1861 B.n619 B.n617 163.367
R1862 B.n623 B.n542 163.367
R1863 B.n627 B.n625 163.367
R1864 B.n631 B.n540 163.367
R1865 B.n635 B.n633 163.367
R1866 B.n642 B.n538 163.367
R1867 B.n646 B.n644 163.367
R1868 B.n650 B.n536 163.367
R1869 B.n654 B.n652 163.367
R1870 B.n658 B.n534 163.367
R1871 B.n662 B.n660 163.367
R1872 B.n667 B.n530 163.367
R1873 B.n671 B.n669 163.367
R1874 B.n675 B.n528 163.367
R1875 B.n679 B.n677 163.367
R1876 B.n683 B.n526 163.367
R1877 B.n687 B.n685 163.367
R1878 B.n691 B.n524 163.367
R1879 B.n695 B.n693 163.367
R1880 B.n699 B.n522 163.367
R1881 B.n703 B.n701 163.367
R1882 B.n707 B.n520 163.367
R1883 B.n711 B.n709 163.367
R1884 B.n715 B.n518 163.367
R1885 B.n719 B.n717 163.367
R1886 B.n723 B.n516 163.367
R1887 B.n727 B.n725 163.367
R1888 B.n731 B.n514 163.367
R1889 B.n735 B.n733 163.367
R1890 B.n739 B.n512 163.367
R1891 B.n742 B.n741 163.367
R1892 B.n744 B.n509 163.367
R1893 B.n748 B.n503 163.367
R1894 B.n756 B.n503 163.367
R1895 B.n756 B.n501 163.367
R1896 B.n760 B.n501 163.367
R1897 B.n760 B.n495 163.367
R1898 B.n768 B.n495 163.367
R1899 B.n768 B.n493 163.367
R1900 B.n772 B.n493 163.367
R1901 B.n772 B.n487 163.367
R1902 B.n780 B.n487 163.367
R1903 B.n780 B.n485 163.367
R1904 B.n784 B.n485 163.367
R1905 B.n784 B.n479 163.367
R1906 B.n792 B.n479 163.367
R1907 B.n792 B.n477 163.367
R1908 B.n796 B.n477 163.367
R1909 B.n796 B.n471 163.367
R1910 B.n804 B.n471 163.367
R1911 B.n804 B.n469 163.367
R1912 B.n808 B.n469 163.367
R1913 B.n808 B.n463 163.367
R1914 B.n816 B.n463 163.367
R1915 B.n816 B.n461 163.367
R1916 B.n820 B.n461 163.367
R1917 B.n820 B.n455 163.367
R1918 B.n828 B.n455 163.367
R1919 B.n828 B.n453 163.367
R1920 B.n832 B.n453 163.367
R1921 B.n832 B.n447 163.367
R1922 B.n840 B.n447 163.367
R1923 B.n840 B.n445 163.367
R1924 B.n844 B.n445 163.367
R1925 B.n844 B.n440 163.367
R1926 B.n853 B.n440 163.367
R1927 B.n853 B.n438 163.367
R1928 B.n857 B.n438 163.367
R1929 B.n857 B.n432 163.367
R1930 B.n865 B.n432 163.367
R1931 B.n865 B.n430 163.367
R1932 B.n869 B.n430 163.367
R1933 B.n869 B.n423 163.367
R1934 B.n877 B.n423 163.367
R1935 B.n877 B.n421 163.367
R1936 B.n881 B.n421 163.367
R1937 B.n881 B.n416 163.367
R1938 B.n889 B.n416 163.367
R1939 B.n889 B.n414 163.367
R1940 B.n893 B.n414 163.367
R1941 B.n893 B.n408 163.367
R1942 B.n901 B.n408 163.367
R1943 B.n901 B.n406 163.367
R1944 B.n905 B.n406 163.367
R1945 B.n905 B.n400 163.367
R1946 B.n913 B.n400 163.367
R1947 B.n913 B.n398 163.367
R1948 B.n917 B.n398 163.367
R1949 B.n917 B.n392 163.367
R1950 B.n925 B.n392 163.367
R1951 B.n925 B.n390 163.367
R1952 B.n929 B.n390 163.367
R1953 B.n929 B.n384 163.367
R1954 B.n937 B.n384 163.367
R1955 B.n937 B.n382 163.367
R1956 B.n941 B.n382 163.367
R1957 B.n941 B.n377 163.367
R1958 B.n950 B.n377 163.367
R1959 B.n950 B.n375 163.367
R1960 B.n955 B.n375 163.367
R1961 B.n955 B.n369 163.367
R1962 B.n963 B.n369 163.367
R1963 B.n964 B.n963 163.367
R1964 B.n964 B.n5 163.367
R1965 B.n6 B.n5 163.367
R1966 B.n7 B.n6 163.367
R1967 B.n969 B.n7 163.367
R1968 B.n969 B.n12 163.367
R1969 B.n13 B.n12 163.367
R1970 B.n14 B.n13 163.367
R1971 B.n974 B.n14 163.367
R1972 B.n974 B.n19 163.367
R1973 B.n20 B.n19 163.367
R1974 B.n21 B.n20 163.367
R1975 B.n979 B.n21 163.367
R1976 B.n979 B.n26 163.367
R1977 B.n27 B.n26 163.367
R1978 B.n28 B.n27 163.367
R1979 B.n984 B.n28 163.367
R1980 B.n984 B.n33 163.367
R1981 B.n34 B.n33 163.367
R1982 B.n35 B.n34 163.367
R1983 B.n989 B.n35 163.367
R1984 B.n989 B.n40 163.367
R1985 B.n41 B.n40 163.367
R1986 B.n42 B.n41 163.367
R1987 B.n994 B.n42 163.367
R1988 B.n994 B.n47 163.367
R1989 B.n48 B.n47 163.367
R1990 B.n49 B.n48 163.367
R1991 B.n999 B.n49 163.367
R1992 B.n999 B.n54 163.367
R1993 B.n55 B.n54 163.367
R1994 B.n56 B.n55 163.367
R1995 B.n1004 B.n56 163.367
R1996 B.n1004 B.n61 163.367
R1997 B.n62 B.n61 163.367
R1998 B.n63 B.n62 163.367
R1999 B.n1009 B.n63 163.367
R2000 B.n1009 B.n68 163.367
R2001 B.n69 B.n68 163.367
R2002 B.n70 B.n69 163.367
R2003 B.n1014 B.n70 163.367
R2004 B.n1014 B.n75 163.367
R2005 B.n76 B.n75 163.367
R2006 B.n77 B.n76 163.367
R2007 B.n1019 B.n77 163.367
R2008 B.n1019 B.n82 163.367
R2009 B.n83 B.n82 163.367
R2010 B.n84 B.n83 163.367
R2011 B.n1024 B.n84 163.367
R2012 B.n1024 B.n89 163.367
R2013 B.n90 B.n89 163.367
R2014 B.n91 B.n90 163.367
R2015 B.n1029 B.n91 163.367
R2016 B.n1029 B.n96 163.367
R2017 B.n97 B.n96 163.367
R2018 B.n98 B.n97 163.367
R2019 B.n1034 B.n98 163.367
R2020 B.n1034 B.n103 163.367
R2021 B.n104 B.n103 163.367
R2022 B.n105 B.n104 163.367
R2023 B.n1039 B.n105 163.367
R2024 B.n1039 B.n110 163.367
R2025 B.n111 B.n110 163.367
R2026 B.n112 B.n111 163.367
R2027 B.n1044 B.n112 163.367
R2028 B.n1044 B.n117 163.367
R2029 B.n118 B.n117 163.367
R2030 B.n119 B.n118 163.367
R2031 B.n1049 B.n119 163.367
R2032 B.n1049 B.n124 163.367
R2033 B.n125 B.n124 163.367
R2034 B.n126 B.n125 163.367
R2035 B.n1054 B.n126 163.367
R2036 B.n1054 B.n131 163.367
R2037 B.n187 B.n186 163.367
R2038 B.n191 B.n190 163.367
R2039 B.n195 B.n194 163.367
R2040 B.n199 B.n198 163.367
R2041 B.n203 B.n202 163.367
R2042 B.n207 B.n206 163.367
R2043 B.n211 B.n210 163.367
R2044 B.n215 B.n214 163.367
R2045 B.n219 B.n218 163.367
R2046 B.n223 B.n222 163.367
R2047 B.n227 B.n226 163.367
R2048 B.n231 B.n230 163.367
R2049 B.n235 B.n234 163.367
R2050 B.n239 B.n238 163.367
R2051 B.n243 B.n242 163.367
R2052 B.n247 B.n246 163.367
R2053 B.n251 B.n250 163.367
R2054 B.n255 B.n254 163.367
R2055 B.n259 B.n258 163.367
R2056 B.n263 B.n262 163.367
R2057 B.n267 B.n266 163.367
R2058 B.n271 B.n270 163.367
R2059 B.n275 B.n274 163.367
R2060 B.n279 B.n278 163.367
R2061 B.n283 B.n282 163.367
R2062 B.n287 B.n286 163.367
R2063 B.n291 B.n290 163.367
R2064 B.n295 B.n294 163.367
R2065 B.n299 B.n298 163.367
R2066 B.n303 B.n302 163.367
R2067 B.n307 B.n306 163.367
R2068 B.n311 B.n310 163.367
R2069 B.n315 B.n314 163.367
R2070 B.n319 B.n318 163.367
R2071 B.n323 B.n322 163.367
R2072 B.n327 B.n326 163.367
R2073 B.n331 B.n330 163.367
R2074 B.n335 B.n334 163.367
R2075 B.n339 B.n338 163.367
R2076 B.n343 B.n342 163.367
R2077 B.n347 B.n346 163.367
R2078 B.n351 B.n350 163.367
R2079 B.n355 B.n354 163.367
R2080 B.n359 B.n358 163.367
R2081 B.n363 B.n362 163.367
R2082 B.n365 B.n178 163.367
R2083 B.n749 B.n508 84.9304
R2084 B.n1061 B.n1060 84.9304
R2085 B.n559 B.n507 71.676
R2086 B.n563 B.n562 71.676
R2087 B.n568 B.n567 71.676
R2088 B.n571 B.n570 71.676
R2089 B.n576 B.n575 71.676
R2090 B.n579 B.n578 71.676
R2091 B.n584 B.n583 71.676
R2092 B.n587 B.n586 71.676
R2093 B.n592 B.n591 71.676
R2094 B.n595 B.n594 71.676
R2095 B.n600 B.n599 71.676
R2096 B.n603 B.n602 71.676
R2097 B.n608 B.n607 71.676
R2098 B.n611 B.n610 71.676
R2099 B.n616 B.n615 71.676
R2100 B.n619 B.n618 71.676
R2101 B.n624 B.n623 71.676
R2102 B.n627 B.n626 71.676
R2103 B.n632 B.n631 71.676
R2104 B.n635 B.n634 71.676
R2105 B.n643 B.n642 71.676
R2106 B.n646 B.n645 71.676
R2107 B.n651 B.n650 71.676
R2108 B.n654 B.n653 71.676
R2109 B.n659 B.n658 71.676
R2110 B.n662 B.n661 71.676
R2111 B.n668 B.n667 71.676
R2112 B.n671 B.n670 71.676
R2113 B.n676 B.n675 71.676
R2114 B.n679 B.n678 71.676
R2115 B.n684 B.n683 71.676
R2116 B.n687 B.n686 71.676
R2117 B.n692 B.n691 71.676
R2118 B.n695 B.n694 71.676
R2119 B.n700 B.n699 71.676
R2120 B.n703 B.n702 71.676
R2121 B.n708 B.n707 71.676
R2122 B.n711 B.n710 71.676
R2123 B.n716 B.n715 71.676
R2124 B.n719 B.n718 71.676
R2125 B.n724 B.n723 71.676
R2126 B.n727 B.n726 71.676
R2127 B.n732 B.n731 71.676
R2128 B.n735 B.n734 71.676
R2129 B.n740 B.n739 71.676
R2130 B.n743 B.n742 71.676
R2131 B.n132 B.n130 71.676
R2132 B.n187 B.n133 71.676
R2133 B.n191 B.n134 71.676
R2134 B.n195 B.n135 71.676
R2135 B.n199 B.n136 71.676
R2136 B.n203 B.n137 71.676
R2137 B.n207 B.n138 71.676
R2138 B.n211 B.n139 71.676
R2139 B.n215 B.n140 71.676
R2140 B.n219 B.n141 71.676
R2141 B.n223 B.n142 71.676
R2142 B.n227 B.n143 71.676
R2143 B.n231 B.n144 71.676
R2144 B.n235 B.n145 71.676
R2145 B.n239 B.n146 71.676
R2146 B.n243 B.n147 71.676
R2147 B.n247 B.n148 71.676
R2148 B.n251 B.n149 71.676
R2149 B.n255 B.n150 71.676
R2150 B.n259 B.n151 71.676
R2151 B.n263 B.n152 71.676
R2152 B.n267 B.n153 71.676
R2153 B.n271 B.n154 71.676
R2154 B.n275 B.n155 71.676
R2155 B.n279 B.n156 71.676
R2156 B.n283 B.n157 71.676
R2157 B.n287 B.n158 71.676
R2158 B.n291 B.n159 71.676
R2159 B.n295 B.n160 71.676
R2160 B.n299 B.n161 71.676
R2161 B.n303 B.n162 71.676
R2162 B.n307 B.n163 71.676
R2163 B.n311 B.n164 71.676
R2164 B.n315 B.n165 71.676
R2165 B.n319 B.n166 71.676
R2166 B.n323 B.n167 71.676
R2167 B.n327 B.n168 71.676
R2168 B.n331 B.n169 71.676
R2169 B.n335 B.n170 71.676
R2170 B.n339 B.n171 71.676
R2171 B.n343 B.n172 71.676
R2172 B.n347 B.n173 71.676
R2173 B.n351 B.n174 71.676
R2174 B.n355 B.n175 71.676
R2175 B.n359 B.n176 71.676
R2176 B.n363 B.n177 71.676
R2177 B.n1059 B.n178 71.676
R2178 B.n1059 B.n1058 71.676
R2179 B.n365 B.n177 71.676
R2180 B.n362 B.n176 71.676
R2181 B.n358 B.n175 71.676
R2182 B.n354 B.n174 71.676
R2183 B.n350 B.n173 71.676
R2184 B.n346 B.n172 71.676
R2185 B.n342 B.n171 71.676
R2186 B.n338 B.n170 71.676
R2187 B.n334 B.n169 71.676
R2188 B.n330 B.n168 71.676
R2189 B.n326 B.n167 71.676
R2190 B.n322 B.n166 71.676
R2191 B.n318 B.n165 71.676
R2192 B.n314 B.n164 71.676
R2193 B.n310 B.n163 71.676
R2194 B.n306 B.n162 71.676
R2195 B.n302 B.n161 71.676
R2196 B.n298 B.n160 71.676
R2197 B.n294 B.n159 71.676
R2198 B.n290 B.n158 71.676
R2199 B.n286 B.n157 71.676
R2200 B.n282 B.n156 71.676
R2201 B.n278 B.n155 71.676
R2202 B.n274 B.n154 71.676
R2203 B.n270 B.n153 71.676
R2204 B.n266 B.n152 71.676
R2205 B.n262 B.n151 71.676
R2206 B.n258 B.n150 71.676
R2207 B.n254 B.n149 71.676
R2208 B.n250 B.n148 71.676
R2209 B.n246 B.n147 71.676
R2210 B.n242 B.n146 71.676
R2211 B.n238 B.n145 71.676
R2212 B.n234 B.n144 71.676
R2213 B.n230 B.n143 71.676
R2214 B.n226 B.n142 71.676
R2215 B.n222 B.n141 71.676
R2216 B.n218 B.n140 71.676
R2217 B.n214 B.n139 71.676
R2218 B.n210 B.n138 71.676
R2219 B.n206 B.n137 71.676
R2220 B.n202 B.n136 71.676
R2221 B.n198 B.n135 71.676
R2222 B.n194 B.n134 71.676
R2223 B.n190 B.n133 71.676
R2224 B.n186 B.n132 71.676
R2225 B.n560 B.n559 71.676
R2226 B.n562 B.n556 71.676
R2227 B.n569 B.n568 71.676
R2228 B.n570 B.n554 71.676
R2229 B.n577 B.n576 71.676
R2230 B.n578 B.n552 71.676
R2231 B.n585 B.n584 71.676
R2232 B.n586 B.n550 71.676
R2233 B.n593 B.n592 71.676
R2234 B.n594 B.n548 71.676
R2235 B.n601 B.n600 71.676
R2236 B.n602 B.n546 71.676
R2237 B.n609 B.n608 71.676
R2238 B.n610 B.n544 71.676
R2239 B.n617 B.n616 71.676
R2240 B.n618 B.n542 71.676
R2241 B.n625 B.n624 71.676
R2242 B.n626 B.n540 71.676
R2243 B.n633 B.n632 71.676
R2244 B.n634 B.n538 71.676
R2245 B.n644 B.n643 71.676
R2246 B.n645 B.n536 71.676
R2247 B.n652 B.n651 71.676
R2248 B.n653 B.n534 71.676
R2249 B.n660 B.n659 71.676
R2250 B.n661 B.n530 71.676
R2251 B.n669 B.n668 71.676
R2252 B.n670 B.n528 71.676
R2253 B.n677 B.n676 71.676
R2254 B.n678 B.n526 71.676
R2255 B.n685 B.n684 71.676
R2256 B.n686 B.n524 71.676
R2257 B.n693 B.n692 71.676
R2258 B.n694 B.n522 71.676
R2259 B.n701 B.n700 71.676
R2260 B.n702 B.n520 71.676
R2261 B.n709 B.n708 71.676
R2262 B.n710 B.n518 71.676
R2263 B.n717 B.n716 71.676
R2264 B.n718 B.n516 71.676
R2265 B.n725 B.n724 71.676
R2266 B.n726 B.n514 71.676
R2267 B.n733 B.n732 71.676
R2268 B.n734 B.n512 71.676
R2269 B.n741 B.n740 71.676
R2270 B.n744 B.n743 71.676
R2271 B.n532 B.n531 70.4005
R2272 B.n639 B.n638 70.4005
R2273 B.n183 B.n182 70.4005
R2274 B.n180 B.n179 70.4005
R2275 B.n664 B.n532 59.5399
R2276 B.n640 B.n639 59.5399
R2277 B.n184 B.n183 59.5399
R2278 B.n181 B.n180 59.5399
R2279 B.n749 B.n504 42.78
R2280 B.n755 B.n504 42.78
R2281 B.n755 B.n500 42.78
R2282 B.n761 B.n500 42.78
R2283 B.n761 B.n496 42.78
R2284 B.n767 B.n496 42.78
R2285 B.n767 B.n492 42.78
R2286 B.n773 B.n492 42.78
R2287 B.n779 B.n488 42.78
R2288 B.n779 B.n484 42.78
R2289 B.n785 B.n484 42.78
R2290 B.n785 B.n480 42.78
R2291 B.n791 B.n480 42.78
R2292 B.n791 B.n476 42.78
R2293 B.n797 B.n476 42.78
R2294 B.n797 B.n472 42.78
R2295 B.n803 B.n472 42.78
R2296 B.n803 B.n468 42.78
R2297 B.n809 B.n468 42.78
R2298 B.n809 B.n464 42.78
R2299 B.n815 B.n464 42.78
R2300 B.n821 B.n460 42.78
R2301 B.n821 B.n456 42.78
R2302 B.n827 B.n456 42.78
R2303 B.n827 B.n452 42.78
R2304 B.n833 B.n452 42.78
R2305 B.n833 B.n448 42.78
R2306 B.n839 B.n448 42.78
R2307 B.n839 B.n444 42.78
R2308 B.n846 B.n444 42.78
R2309 B.n846 B.n845 42.78
R2310 B.n852 B.n437 42.78
R2311 B.n858 B.n437 42.78
R2312 B.n858 B.n433 42.78
R2313 B.n864 B.n433 42.78
R2314 B.n864 B.n429 42.78
R2315 B.n870 B.n429 42.78
R2316 B.n870 B.n424 42.78
R2317 B.n876 B.n424 42.78
R2318 B.n876 B.n425 42.78
R2319 B.n882 B.n417 42.78
R2320 B.n888 B.n417 42.78
R2321 B.n888 B.n413 42.78
R2322 B.n894 B.n413 42.78
R2323 B.n894 B.n409 42.78
R2324 B.n900 B.n409 42.78
R2325 B.n900 B.n405 42.78
R2326 B.n906 B.n405 42.78
R2327 B.n906 B.n401 42.78
R2328 B.n912 B.n401 42.78
R2329 B.n918 B.n397 42.78
R2330 B.n918 B.n393 42.78
R2331 B.n924 B.n393 42.78
R2332 B.n924 B.n389 42.78
R2333 B.n930 B.n389 42.78
R2334 B.n930 B.n385 42.78
R2335 B.n936 B.n385 42.78
R2336 B.n936 B.n381 42.78
R2337 B.n943 B.n381 42.78
R2338 B.n943 B.n942 42.78
R2339 B.n949 B.n374 42.78
R2340 B.n956 B.n374 42.78
R2341 B.n956 B.n370 42.78
R2342 B.n962 B.n370 42.78
R2343 B.n962 B.n4 42.78
R2344 B.n1205 B.n4 42.78
R2345 B.n1205 B.n1204 42.78
R2346 B.n1204 B.n1203 42.78
R2347 B.n1203 B.n8 42.78
R2348 B.n1197 B.n8 42.78
R2349 B.n1197 B.n1196 42.78
R2350 B.n1196 B.n1195 42.78
R2351 B.n1189 B.n18 42.78
R2352 B.n1189 B.n1188 42.78
R2353 B.n1188 B.n1187 42.78
R2354 B.n1187 B.n22 42.78
R2355 B.n1181 B.n22 42.78
R2356 B.n1181 B.n1180 42.78
R2357 B.n1180 B.n1179 42.78
R2358 B.n1179 B.n29 42.78
R2359 B.n1173 B.n29 42.78
R2360 B.n1173 B.n1172 42.78
R2361 B.n1171 B.n36 42.78
R2362 B.n1165 B.n36 42.78
R2363 B.n1165 B.n1164 42.78
R2364 B.n1164 B.n1163 42.78
R2365 B.n1163 B.n43 42.78
R2366 B.n1157 B.n43 42.78
R2367 B.n1157 B.n1156 42.78
R2368 B.n1156 B.n1155 42.78
R2369 B.n1155 B.n50 42.78
R2370 B.n1149 B.n50 42.78
R2371 B.n1148 B.n1147 42.78
R2372 B.n1147 B.n57 42.78
R2373 B.n1141 B.n57 42.78
R2374 B.n1141 B.n1140 42.78
R2375 B.n1140 B.n1139 42.78
R2376 B.n1139 B.n64 42.78
R2377 B.n1133 B.n64 42.78
R2378 B.n1133 B.n1132 42.78
R2379 B.n1132 B.n1131 42.78
R2380 B.n1125 B.n74 42.78
R2381 B.n1125 B.n1124 42.78
R2382 B.n1124 B.n1123 42.78
R2383 B.n1123 B.n78 42.78
R2384 B.n1117 B.n78 42.78
R2385 B.n1117 B.n1116 42.78
R2386 B.n1116 B.n1115 42.78
R2387 B.n1115 B.n85 42.78
R2388 B.n1109 B.n85 42.78
R2389 B.n1109 B.n1108 42.78
R2390 B.n1107 B.n92 42.78
R2391 B.n1101 B.n92 42.78
R2392 B.n1101 B.n1100 42.78
R2393 B.n1100 B.n1099 42.78
R2394 B.n1099 B.n99 42.78
R2395 B.n1093 B.n99 42.78
R2396 B.n1093 B.n1092 42.78
R2397 B.n1092 B.n1091 42.78
R2398 B.n1091 B.n106 42.78
R2399 B.n1085 B.n106 42.78
R2400 B.n1085 B.n1084 42.78
R2401 B.n1084 B.n1083 42.78
R2402 B.n1083 B.n113 42.78
R2403 B.n1077 B.n1076 42.78
R2404 B.n1076 B.n1075 42.78
R2405 B.n1075 B.n120 42.78
R2406 B.n1069 B.n120 42.78
R2407 B.n1069 B.n1068 42.78
R2408 B.n1068 B.n1067 42.78
R2409 B.n1067 B.n127 42.78
R2410 B.n1061 B.n127 42.78
R2411 B.n852 B.t7 41.5218
R2412 B.n1131 B.t4 41.5218
R2413 B.n949 B.t0 40.2636
R2414 B.n1195 B.t8 40.2636
R2415 B.n1063 B.n129 34.4981
R2416 B.n1057 B.n1056 34.4981
R2417 B.n747 B.n746 34.4981
R2418 B.n751 B.n506 34.4981
R2419 B.n425 B.t5 30.1978
R2420 B.t6 B.n1148 30.1978
R2421 B.t2 B.n460 27.6814
R2422 B.n1108 B.t1 27.6814
R2423 B.t3 B.n397 26.4231
R2424 B.n1172 B.t9 26.4231
R2425 B.t15 B.n488 22.6485
R2426 B.t11 B.n113 22.6485
R2427 B.n773 B.t15 20.132
R2428 B.n1077 B.t11 20.132
R2429 B B.n1207 18.0485
R2430 B.n912 B.t3 16.3574
R2431 B.t9 B.n1171 16.3574
R2432 B.n815 B.t2 15.0992
R2433 B.t1 B.n1107 15.0992
R2434 B.n882 B.t5 12.5827
R2435 B.n1149 B.t6 12.5827
R2436 B.n185 B.n129 10.6151
R2437 B.n188 B.n185 10.6151
R2438 B.n189 B.n188 10.6151
R2439 B.n192 B.n189 10.6151
R2440 B.n193 B.n192 10.6151
R2441 B.n196 B.n193 10.6151
R2442 B.n197 B.n196 10.6151
R2443 B.n200 B.n197 10.6151
R2444 B.n201 B.n200 10.6151
R2445 B.n204 B.n201 10.6151
R2446 B.n205 B.n204 10.6151
R2447 B.n208 B.n205 10.6151
R2448 B.n209 B.n208 10.6151
R2449 B.n212 B.n209 10.6151
R2450 B.n213 B.n212 10.6151
R2451 B.n216 B.n213 10.6151
R2452 B.n217 B.n216 10.6151
R2453 B.n220 B.n217 10.6151
R2454 B.n221 B.n220 10.6151
R2455 B.n224 B.n221 10.6151
R2456 B.n225 B.n224 10.6151
R2457 B.n228 B.n225 10.6151
R2458 B.n229 B.n228 10.6151
R2459 B.n232 B.n229 10.6151
R2460 B.n233 B.n232 10.6151
R2461 B.n236 B.n233 10.6151
R2462 B.n237 B.n236 10.6151
R2463 B.n240 B.n237 10.6151
R2464 B.n241 B.n240 10.6151
R2465 B.n244 B.n241 10.6151
R2466 B.n245 B.n244 10.6151
R2467 B.n248 B.n245 10.6151
R2468 B.n249 B.n248 10.6151
R2469 B.n252 B.n249 10.6151
R2470 B.n253 B.n252 10.6151
R2471 B.n256 B.n253 10.6151
R2472 B.n257 B.n256 10.6151
R2473 B.n260 B.n257 10.6151
R2474 B.n261 B.n260 10.6151
R2475 B.n264 B.n261 10.6151
R2476 B.n265 B.n264 10.6151
R2477 B.n269 B.n268 10.6151
R2478 B.n272 B.n269 10.6151
R2479 B.n273 B.n272 10.6151
R2480 B.n276 B.n273 10.6151
R2481 B.n277 B.n276 10.6151
R2482 B.n280 B.n277 10.6151
R2483 B.n281 B.n280 10.6151
R2484 B.n284 B.n281 10.6151
R2485 B.n285 B.n284 10.6151
R2486 B.n289 B.n288 10.6151
R2487 B.n292 B.n289 10.6151
R2488 B.n293 B.n292 10.6151
R2489 B.n296 B.n293 10.6151
R2490 B.n297 B.n296 10.6151
R2491 B.n300 B.n297 10.6151
R2492 B.n301 B.n300 10.6151
R2493 B.n304 B.n301 10.6151
R2494 B.n305 B.n304 10.6151
R2495 B.n308 B.n305 10.6151
R2496 B.n309 B.n308 10.6151
R2497 B.n312 B.n309 10.6151
R2498 B.n313 B.n312 10.6151
R2499 B.n316 B.n313 10.6151
R2500 B.n317 B.n316 10.6151
R2501 B.n320 B.n317 10.6151
R2502 B.n321 B.n320 10.6151
R2503 B.n324 B.n321 10.6151
R2504 B.n325 B.n324 10.6151
R2505 B.n328 B.n325 10.6151
R2506 B.n329 B.n328 10.6151
R2507 B.n332 B.n329 10.6151
R2508 B.n333 B.n332 10.6151
R2509 B.n336 B.n333 10.6151
R2510 B.n337 B.n336 10.6151
R2511 B.n340 B.n337 10.6151
R2512 B.n341 B.n340 10.6151
R2513 B.n344 B.n341 10.6151
R2514 B.n345 B.n344 10.6151
R2515 B.n348 B.n345 10.6151
R2516 B.n349 B.n348 10.6151
R2517 B.n352 B.n349 10.6151
R2518 B.n353 B.n352 10.6151
R2519 B.n356 B.n353 10.6151
R2520 B.n357 B.n356 10.6151
R2521 B.n360 B.n357 10.6151
R2522 B.n361 B.n360 10.6151
R2523 B.n364 B.n361 10.6151
R2524 B.n366 B.n364 10.6151
R2525 B.n367 B.n366 10.6151
R2526 B.n1057 B.n367 10.6151
R2527 B.n747 B.n502 10.6151
R2528 B.n757 B.n502 10.6151
R2529 B.n758 B.n757 10.6151
R2530 B.n759 B.n758 10.6151
R2531 B.n759 B.n494 10.6151
R2532 B.n769 B.n494 10.6151
R2533 B.n770 B.n769 10.6151
R2534 B.n771 B.n770 10.6151
R2535 B.n771 B.n486 10.6151
R2536 B.n781 B.n486 10.6151
R2537 B.n782 B.n781 10.6151
R2538 B.n783 B.n782 10.6151
R2539 B.n783 B.n478 10.6151
R2540 B.n793 B.n478 10.6151
R2541 B.n794 B.n793 10.6151
R2542 B.n795 B.n794 10.6151
R2543 B.n795 B.n470 10.6151
R2544 B.n805 B.n470 10.6151
R2545 B.n806 B.n805 10.6151
R2546 B.n807 B.n806 10.6151
R2547 B.n807 B.n462 10.6151
R2548 B.n817 B.n462 10.6151
R2549 B.n818 B.n817 10.6151
R2550 B.n819 B.n818 10.6151
R2551 B.n819 B.n454 10.6151
R2552 B.n829 B.n454 10.6151
R2553 B.n830 B.n829 10.6151
R2554 B.n831 B.n830 10.6151
R2555 B.n831 B.n446 10.6151
R2556 B.n841 B.n446 10.6151
R2557 B.n842 B.n841 10.6151
R2558 B.n843 B.n842 10.6151
R2559 B.n843 B.n439 10.6151
R2560 B.n854 B.n439 10.6151
R2561 B.n855 B.n854 10.6151
R2562 B.n856 B.n855 10.6151
R2563 B.n856 B.n431 10.6151
R2564 B.n866 B.n431 10.6151
R2565 B.n867 B.n866 10.6151
R2566 B.n868 B.n867 10.6151
R2567 B.n868 B.n422 10.6151
R2568 B.n878 B.n422 10.6151
R2569 B.n879 B.n878 10.6151
R2570 B.n880 B.n879 10.6151
R2571 B.n880 B.n415 10.6151
R2572 B.n890 B.n415 10.6151
R2573 B.n891 B.n890 10.6151
R2574 B.n892 B.n891 10.6151
R2575 B.n892 B.n407 10.6151
R2576 B.n902 B.n407 10.6151
R2577 B.n903 B.n902 10.6151
R2578 B.n904 B.n903 10.6151
R2579 B.n904 B.n399 10.6151
R2580 B.n914 B.n399 10.6151
R2581 B.n915 B.n914 10.6151
R2582 B.n916 B.n915 10.6151
R2583 B.n916 B.n391 10.6151
R2584 B.n926 B.n391 10.6151
R2585 B.n927 B.n926 10.6151
R2586 B.n928 B.n927 10.6151
R2587 B.n928 B.n383 10.6151
R2588 B.n938 B.n383 10.6151
R2589 B.n939 B.n938 10.6151
R2590 B.n940 B.n939 10.6151
R2591 B.n940 B.n376 10.6151
R2592 B.n951 B.n376 10.6151
R2593 B.n952 B.n951 10.6151
R2594 B.n954 B.n952 10.6151
R2595 B.n954 B.n953 10.6151
R2596 B.n953 B.n368 10.6151
R2597 B.n965 B.n368 10.6151
R2598 B.n966 B.n965 10.6151
R2599 B.n967 B.n966 10.6151
R2600 B.n968 B.n967 10.6151
R2601 B.n970 B.n968 10.6151
R2602 B.n971 B.n970 10.6151
R2603 B.n972 B.n971 10.6151
R2604 B.n973 B.n972 10.6151
R2605 B.n975 B.n973 10.6151
R2606 B.n976 B.n975 10.6151
R2607 B.n977 B.n976 10.6151
R2608 B.n978 B.n977 10.6151
R2609 B.n980 B.n978 10.6151
R2610 B.n981 B.n980 10.6151
R2611 B.n982 B.n981 10.6151
R2612 B.n983 B.n982 10.6151
R2613 B.n985 B.n983 10.6151
R2614 B.n986 B.n985 10.6151
R2615 B.n987 B.n986 10.6151
R2616 B.n988 B.n987 10.6151
R2617 B.n990 B.n988 10.6151
R2618 B.n991 B.n990 10.6151
R2619 B.n992 B.n991 10.6151
R2620 B.n993 B.n992 10.6151
R2621 B.n995 B.n993 10.6151
R2622 B.n996 B.n995 10.6151
R2623 B.n997 B.n996 10.6151
R2624 B.n998 B.n997 10.6151
R2625 B.n1000 B.n998 10.6151
R2626 B.n1001 B.n1000 10.6151
R2627 B.n1002 B.n1001 10.6151
R2628 B.n1003 B.n1002 10.6151
R2629 B.n1005 B.n1003 10.6151
R2630 B.n1006 B.n1005 10.6151
R2631 B.n1007 B.n1006 10.6151
R2632 B.n1008 B.n1007 10.6151
R2633 B.n1010 B.n1008 10.6151
R2634 B.n1011 B.n1010 10.6151
R2635 B.n1012 B.n1011 10.6151
R2636 B.n1013 B.n1012 10.6151
R2637 B.n1015 B.n1013 10.6151
R2638 B.n1016 B.n1015 10.6151
R2639 B.n1017 B.n1016 10.6151
R2640 B.n1018 B.n1017 10.6151
R2641 B.n1020 B.n1018 10.6151
R2642 B.n1021 B.n1020 10.6151
R2643 B.n1022 B.n1021 10.6151
R2644 B.n1023 B.n1022 10.6151
R2645 B.n1025 B.n1023 10.6151
R2646 B.n1026 B.n1025 10.6151
R2647 B.n1027 B.n1026 10.6151
R2648 B.n1028 B.n1027 10.6151
R2649 B.n1030 B.n1028 10.6151
R2650 B.n1031 B.n1030 10.6151
R2651 B.n1032 B.n1031 10.6151
R2652 B.n1033 B.n1032 10.6151
R2653 B.n1035 B.n1033 10.6151
R2654 B.n1036 B.n1035 10.6151
R2655 B.n1037 B.n1036 10.6151
R2656 B.n1038 B.n1037 10.6151
R2657 B.n1040 B.n1038 10.6151
R2658 B.n1041 B.n1040 10.6151
R2659 B.n1042 B.n1041 10.6151
R2660 B.n1043 B.n1042 10.6151
R2661 B.n1045 B.n1043 10.6151
R2662 B.n1046 B.n1045 10.6151
R2663 B.n1047 B.n1046 10.6151
R2664 B.n1048 B.n1047 10.6151
R2665 B.n1050 B.n1048 10.6151
R2666 B.n1051 B.n1050 10.6151
R2667 B.n1052 B.n1051 10.6151
R2668 B.n1053 B.n1052 10.6151
R2669 B.n1055 B.n1053 10.6151
R2670 B.n1056 B.n1055 10.6151
R2671 B.n558 B.n506 10.6151
R2672 B.n558 B.n557 10.6151
R2673 B.n564 B.n557 10.6151
R2674 B.n565 B.n564 10.6151
R2675 B.n566 B.n565 10.6151
R2676 B.n566 B.n555 10.6151
R2677 B.n572 B.n555 10.6151
R2678 B.n573 B.n572 10.6151
R2679 B.n574 B.n573 10.6151
R2680 B.n574 B.n553 10.6151
R2681 B.n580 B.n553 10.6151
R2682 B.n581 B.n580 10.6151
R2683 B.n582 B.n581 10.6151
R2684 B.n582 B.n551 10.6151
R2685 B.n588 B.n551 10.6151
R2686 B.n589 B.n588 10.6151
R2687 B.n590 B.n589 10.6151
R2688 B.n590 B.n549 10.6151
R2689 B.n596 B.n549 10.6151
R2690 B.n597 B.n596 10.6151
R2691 B.n598 B.n597 10.6151
R2692 B.n598 B.n547 10.6151
R2693 B.n604 B.n547 10.6151
R2694 B.n605 B.n604 10.6151
R2695 B.n606 B.n605 10.6151
R2696 B.n606 B.n545 10.6151
R2697 B.n612 B.n545 10.6151
R2698 B.n613 B.n612 10.6151
R2699 B.n614 B.n613 10.6151
R2700 B.n614 B.n543 10.6151
R2701 B.n620 B.n543 10.6151
R2702 B.n621 B.n620 10.6151
R2703 B.n622 B.n621 10.6151
R2704 B.n622 B.n541 10.6151
R2705 B.n628 B.n541 10.6151
R2706 B.n629 B.n628 10.6151
R2707 B.n630 B.n629 10.6151
R2708 B.n630 B.n539 10.6151
R2709 B.n636 B.n539 10.6151
R2710 B.n637 B.n636 10.6151
R2711 B.n641 B.n637 10.6151
R2712 B.n647 B.n537 10.6151
R2713 B.n648 B.n647 10.6151
R2714 B.n649 B.n648 10.6151
R2715 B.n649 B.n535 10.6151
R2716 B.n655 B.n535 10.6151
R2717 B.n656 B.n655 10.6151
R2718 B.n657 B.n656 10.6151
R2719 B.n657 B.n533 10.6151
R2720 B.n663 B.n533 10.6151
R2721 B.n666 B.n665 10.6151
R2722 B.n666 B.n529 10.6151
R2723 B.n672 B.n529 10.6151
R2724 B.n673 B.n672 10.6151
R2725 B.n674 B.n673 10.6151
R2726 B.n674 B.n527 10.6151
R2727 B.n680 B.n527 10.6151
R2728 B.n681 B.n680 10.6151
R2729 B.n682 B.n681 10.6151
R2730 B.n682 B.n525 10.6151
R2731 B.n688 B.n525 10.6151
R2732 B.n689 B.n688 10.6151
R2733 B.n690 B.n689 10.6151
R2734 B.n690 B.n523 10.6151
R2735 B.n696 B.n523 10.6151
R2736 B.n697 B.n696 10.6151
R2737 B.n698 B.n697 10.6151
R2738 B.n698 B.n521 10.6151
R2739 B.n704 B.n521 10.6151
R2740 B.n705 B.n704 10.6151
R2741 B.n706 B.n705 10.6151
R2742 B.n706 B.n519 10.6151
R2743 B.n712 B.n519 10.6151
R2744 B.n713 B.n712 10.6151
R2745 B.n714 B.n713 10.6151
R2746 B.n714 B.n517 10.6151
R2747 B.n720 B.n517 10.6151
R2748 B.n721 B.n720 10.6151
R2749 B.n722 B.n721 10.6151
R2750 B.n722 B.n515 10.6151
R2751 B.n728 B.n515 10.6151
R2752 B.n729 B.n728 10.6151
R2753 B.n730 B.n729 10.6151
R2754 B.n730 B.n513 10.6151
R2755 B.n736 B.n513 10.6151
R2756 B.n737 B.n736 10.6151
R2757 B.n738 B.n737 10.6151
R2758 B.n738 B.n511 10.6151
R2759 B.n511 B.n510 10.6151
R2760 B.n745 B.n510 10.6151
R2761 B.n746 B.n745 10.6151
R2762 B.n752 B.n751 10.6151
R2763 B.n753 B.n752 10.6151
R2764 B.n753 B.n498 10.6151
R2765 B.n763 B.n498 10.6151
R2766 B.n764 B.n763 10.6151
R2767 B.n765 B.n764 10.6151
R2768 B.n765 B.n490 10.6151
R2769 B.n775 B.n490 10.6151
R2770 B.n776 B.n775 10.6151
R2771 B.n777 B.n776 10.6151
R2772 B.n777 B.n482 10.6151
R2773 B.n787 B.n482 10.6151
R2774 B.n788 B.n787 10.6151
R2775 B.n789 B.n788 10.6151
R2776 B.n789 B.n474 10.6151
R2777 B.n799 B.n474 10.6151
R2778 B.n800 B.n799 10.6151
R2779 B.n801 B.n800 10.6151
R2780 B.n801 B.n466 10.6151
R2781 B.n811 B.n466 10.6151
R2782 B.n812 B.n811 10.6151
R2783 B.n813 B.n812 10.6151
R2784 B.n813 B.n458 10.6151
R2785 B.n823 B.n458 10.6151
R2786 B.n824 B.n823 10.6151
R2787 B.n825 B.n824 10.6151
R2788 B.n825 B.n450 10.6151
R2789 B.n835 B.n450 10.6151
R2790 B.n836 B.n835 10.6151
R2791 B.n837 B.n836 10.6151
R2792 B.n837 B.n442 10.6151
R2793 B.n848 B.n442 10.6151
R2794 B.n849 B.n848 10.6151
R2795 B.n850 B.n849 10.6151
R2796 B.n850 B.n435 10.6151
R2797 B.n860 B.n435 10.6151
R2798 B.n861 B.n860 10.6151
R2799 B.n862 B.n861 10.6151
R2800 B.n862 B.n427 10.6151
R2801 B.n872 B.n427 10.6151
R2802 B.n873 B.n872 10.6151
R2803 B.n874 B.n873 10.6151
R2804 B.n874 B.n419 10.6151
R2805 B.n884 B.n419 10.6151
R2806 B.n885 B.n884 10.6151
R2807 B.n886 B.n885 10.6151
R2808 B.n886 B.n411 10.6151
R2809 B.n896 B.n411 10.6151
R2810 B.n897 B.n896 10.6151
R2811 B.n898 B.n897 10.6151
R2812 B.n898 B.n403 10.6151
R2813 B.n908 B.n403 10.6151
R2814 B.n909 B.n908 10.6151
R2815 B.n910 B.n909 10.6151
R2816 B.n910 B.n395 10.6151
R2817 B.n920 B.n395 10.6151
R2818 B.n921 B.n920 10.6151
R2819 B.n922 B.n921 10.6151
R2820 B.n922 B.n387 10.6151
R2821 B.n932 B.n387 10.6151
R2822 B.n933 B.n932 10.6151
R2823 B.n934 B.n933 10.6151
R2824 B.n934 B.n379 10.6151
R2825 B.n945 B.n379 10.6151
R2826 B.n946 B.n945 10.6151
R2827 B.n947 B.n946 10.6151
R2828 B.n947 B.n372 10.6151
R2829 B.n958 B.n372 10.6151
R2830 B.n959 B.n958 10.6151
R2831 B.n960 B.n959 10.6151
R2832 B.n960 B.n0 10.6151
R2833 B.n1201 B.n1 10.6151
R2834 B.n1201 B.n1200 10.6151
R2835 B.n1200 B.n1199 10.6151
R2836 B.n1199 B.n10 10.6151
R2837 B.n1193 B.n10 10.6151
R2838 B.n1193 B.n1192 10.6151
R2839 B.n1192 B.n1191 10.6151
R2840 B.n1191 B.n16 10.6151
R2841 B.n1185 B.n16 10.6151
R2842 B.n1185 B.n1184 10.6151
R2843 B.n1184 B.n1183 10.6151
R2844 B.n1183 B.n24 10.6151
R2845 B.n1177 B.n24 10.6151
R2846 B.n1177 B.n1176 10.6151
R2847 B.n1176 B.n1175 10.6151
R2848 B.n1175 B.n31 10.6151
R2849 B.n1169 B.n31 10.6151
R2850 B.n1169 B.n1168 10.6151
R2851 B.n1168 B.n1167 10.6151
R2852 B.n1167 B.n38 10.6151
R2853 B.n1161 B.n38 10.6151
R2854 B.n1161 B.n1160 10.6151
R2855 B.n1160 B.n1159 10.6151
R2856 B.n1159 B.n45 10.6151
R2857 B.n1153 B.n45 10.6151
R2858 B.n1153 B.n1152 10.6151
R2859 B.n1152 B.n1151 10.6151
R2860 B.n1151 B.n52 10.6151
R2861 B.n1145 B.n52 10.6151
R2862 B.n1145 B.n1144 10.6151
R2863 B.n1144 B.n1143 10.6151
R2864 B.n1143 B.n59 10.6151
R2865 B.n1137 B.n59 10.6151
R2866 B.n1137 B.n1136 10.6151
R2867 B.n1136 B.n1135 10.6151
R2868 B.n1135 B.n66 10.6151
R2869 B.n1129 B.n66 10.6151
R2870 B.n1129 B.n1128 10.6151
R2871 B.n1128 B.n1127 10.6151
R2872 B.n1127 B.n72 10.6151
R2873 B.n1121 B.n72 10.6151
R2874 B.n1121 B.n1120 10.6151
R2875 B.n1120 B.n1119 10.6151
R2876 B.n1119 B.n80 10.6151
R2877 B.n1113 B.n80 10.6151
R2878 B.n1113 B.n1112 10.6151
R2879 B.n1112 B.n1111 10.6151
R2880 B.n1111 B.n87 10.6151
R2881 B.n1105 B.n87 10.6151
R2882 B.n1105 B.n1104 10.6151
R2883 B.n1104 B.n1103 10.6151
R2884 B.n1103 B.n94 10.6151
R2885 B.n1097 B.n94 10.6151
R2886 B.n1097 B.n1096 10.6151
R2887 B.n1096 B.n1095 10.6151
R2888 B.n1095 B.n101 10.6151
R2889 B.n1089 B.n101 10.6151
R2890 B.n1089 B.n1088 10.6151
R2891 B.n1088 B.n1087 10.6151
R2892 B.n1087 B.n108 10.6151
R2893 B.n1081 B.n108 10.6151
R2894 B.n1081 B.n1080 10.6151
R2895 B.n1080 B.n1079 10.6151
R2896 B.n1079 B.n115 10.6151
R2897 B.n1073 B.n115 10.6151
R2898 B.n1073 B.n1072 10.6151
R2899 B.n1072 B.n1071 10.6151
R2900 B.n1071 B.n122 10.6151
R2901 B.n1065 B.n122 10.6151
R2902 B.n1065 B.n1064 10.6151
R2903 B.n1064 B.n1063 10.6151
R2904 B.n265 B.n184 9.36635
R2905 B.n288 B.n181 9.36635
R2906 B.n641 B.n640 9.36635
R2907 B.n665 B.n664 9.36635
R2908 B.n1207 B.n0 2.81026
R2909 B.n1207 B.n1 2.81026
R2910 B.n942 B.t0 2.51694
R2911 B.n18 B.t8 2.51694
R2912 B.n845 B.t7 1.25872
R2913 B.n74 B.t4 1.25872
R2914 B.n268 B.n184 1.24928
R2915 B.n285 B.n181 1.24928
R2916 B.n640 B.n537 1.24928
R2917 B.n664 B.n663 1.24928
R2918 VN.n96 VN.n95 161.3
R2919 VN.n94 VN.n50 161.3
R2920 VN.n93 VN.n92 161.3
R2921 VN.n91 VN.n51 161.3
R2922 VN.n90 VN.n89 161.3
R2923 VN.n88 VN.n52 161.3
R2924 VN.n87 VN.n86 161.3
R2925 VN.n85 VN.n84 161.3
R2926 VN.n83 VN.n54 161.3
R2927 VN.n82 VN.n81 161.3
R2928 VN.n80 VN.n55 161.3
R2929 VN.n79 VN.n78 161.3
R2930 VN.n77 VN.n56 161.3
R2931 VN.n76 VN.n75 161.3
R2932 VN.n74 VN.n57 161.3
R2933 VN.n73 VN.n72 161.3
R2934 VN.n71 VN.n58 161.3
R2935 VN.n70 VN.n69 161.3
R2936 VN.n68 VN.n59 161.3
R2937 VN.n67 VN.n66 161.3
R2938 VN.n65 VN.n60 161.3
R2939 VN.n64 VN.n63 161.3
R2940 VN.n47 VN.n46 161.3
R2941 VN.n45 VN.n1 161.3
R2942 VN.n44 VN.n43 161.3
R2943 VN.n42 VN.n2 161.3
R2944 VN.n41 VN.n40 161.3
R2945 VN.n39 VN.n3 161.3
R2946 VN.n38 VN.n37 161.3
R2947 VN.n36 VN.n35 161.3
R2948 VN.n34 VN.n5 161.3
R2949 VN.n33 VN.n32 161.3
R2950 VN.n31 VN.n6 161.3
R2951 VN.n30 VN.n29 161.3
R2952 VN.n28 VN.n7 161.3
R2953 VN.n27 VN.n26 161.3
R2954 VN.n25 VN.n8 161.3
R2955 VN.n24 VN.n23 161.3
R2956 VN.n22 VN.n9 161.3
R2957 VN.n21 VN.n20 161.3
R2958 VN.n19 VN.n10 161.3
R2959 VN.n18 VN.n17 161.3
R2960 VN.n16 VN.n11 161.3
R2961 VN.n15 VN.n14 161.3
R2962 VN.n62 VN.t7 121.793
R2963 VN.n13 VN.t8 121.793
R2964 VN.n8 VN.t3 89.1705
R2965 VN.n12 VN.t9 89.1705
R2966 VN.n4 VN.t4 89.1705
R2967 VN.n0 VN.t6 89.1705
R2968 VN.n57 VN.t5 89.1705
R2969 VN.n61 VN.t1 89.1705
R2970 VN.n53 VN.t0 89.1705
R2971 VN.n49 VN.t2 89.1705
R2972 VN.n48 VN.n0 77.3446
R2973 VN.n97 VN.n49 77.3446
R2974 VN.n62 VN.n61 68.1432
R2975 VN.n13 VN.n12 68.1432
R2976 VN VN.n97 57.3276
R2977 VN.n21 VN.n10 56.5193
R2978 VN.n29 VN.n6 56.5193
R2979 VN.n70 VN.n59 56.5193
R2980 VN.n78 VN.n55 56.5193
R2981 VN.n40 VN.n2 45.8354
R2982 VN.n89 VN.n51 45.8354
R2983 VN.n44 VN.n2 35.1514
R2984 VN.n93 VN.n51 35.1514
R2985 VN.n16 VN.n15 24.4675
R2986 VN.n17 VN.n16 24.4675
R2987 VN.n17 VN.n10 24.4675
R2988 VN.n22 VN.n21 24.4675
R2989 VN.n23 VN.n22 24.4675
R2990 VN.n23 VN.n8 24.4675
R2991 VN.n27 VN.n8 24.4675
R2992 VN.n28 VN.n27 24.4675
R2993 VN.n29 VN.n28 24.4675
R2994 VN.n33 VN.n6 24.4675
R2995 VN.n34 VN.n33 24.4675
R2996 VN.n35 VN.n34 24.4675
R2997 VN.n39 VN.n38 24.4675
R2998 VN.n40 VN.n39 24.4675
R2999 VN.n45 VN.n44 24.4675
R3000 VN.n46 VN.n45 24.4675
R3001 VN.n66 VN.n59 24.4675
R3002 VN.n66 VN.n65 24.4675
R3003 VN.n65 VN.n64 24.4675
R3004 VN.n78 VN.n77 24.4675
R3005 VN.n77 VN.n76 24.4675
R3006 VN.n76 VN.n57 24.4675
R3007 VN.n72 VN.n57 24.4675
R3008 VN.n72 VN.n71 24.4675
R3009 VN.n71 VN.n70 24.4675
R3010 VN.n89 VN.n88 24.4675
R3011 VN.n88 VN.n87 24.4675
R3012 VN.n84 VN.n83 24.4675
R3013 VN.n83 VN.n82 24.4675
R3014 VN.n82 VN.n55 24.4675
R3015 VN.n95 VN.n94 24.4675
R3016 VN.n94 VN.n93 24.4675
R3017 VN.n38 VN.n4 18.1061
R3018 VN.n87 VN.n53 18.1061
R3019 VN.n46 VN.n0 12.7233
R3020 VN.n95 VN.n49 12.7233
R3021 VN.n15 VN.n12 6.36192
R3022 VN.n35 VN.n4 6.36192
R3023 VN.n64 VN.n61 6.36192
R3024 VN.n84 VN.n53 6.36192
R3025 VN.n63 VN.n62 4.26091
R3026 VN.n14 VN.n13 4.26091
R3027 VN.n97 VN.n96 0.354971
R3028 VN.n48 VN.n47 0.354971
R3029 VN VN.n48 0.26696
R3030 VN.n96 VN.n50 0.189894
R3031 VN.n92 VN.n50 0.189894
R3032 VN.n92 VN.n91 0.189894
R3033 VN.n91 VN.n90 0.189894
R3034 VN.n90 VN.n52 0.189894
R3035 VN.n86 VN.n52 0.189894
R3036 VN.n86 VN.n85 0.189894
R3037 VN.n85 VN.n54 0.189894
R3038 VN.n81 VN.n54 0.189894
R3039 VN.n81 VN.n80 0.189894
R3040 VN.n80 VN.n79 0.189894
R3041 VN.n79 VN.n56 0.189894
R3042 VN.n75 VN.n56 0.189894
R3043 VN.n75 VN.n74 0.189894
R3044 VN.n74 VN.n73 0.189894
R3045 VN.n73 VN.n58 0.189894
R3046 VN.n69 VN.n58 0.189894
R3047 VN.n69 VN.n68 0.189894
R3048 VN.n68 VN.n67 0.189894
R3049 VN.n67 VN.n60 0.189894
R3050 VN.n63 VN.n60 0.189894
R3051 VN.n14 VN.n11 0.189894
R3052 VN.n18 VN.n11 0.189894
R3053 VN.n19 VN.n18 0.189894
R3054 VN.n20 VN.n19 0.189894
R3055 VN.n20 VN.n9 0.189894
R3056 VN.n24 VN.n9 0.189894
R3057 VN.n25 VN.n24 0.189894
R3058 VN.n26 VN.n25 0.189894
R3059 VN.n26 VN.n7 0.189894
R3060 VN.n30 VN.n7 0.189894
R3061 VN.n31 VN.n30 0.189894
R3062 VN.n32 VN.n31 0.189894
R3063 VN.n32 VN.n5 0.189894
R3064 VN.n36 VN.n5 0.189894
R3065 VN.n37 VN.n36 0.189894
R3066 VN.n37 VN.n3 0.189894
R3067 VN.n41 VN.n3 0.189894
R3068 VN.n42 VN.n41 0.189894
R3069 VN.n43 VN.n42 0.189894
R3070 VN.n43 VN.n1 0.189894
R3071 VN.n47 VN.n1 0.189894
R3072 VDD2.n129 VDD2.n69 289.615
R3073 VDD2.n60 VDD2.n0 289.615
R3074 VDD2.n130 VDD2.n129 185
R3075 VDD2.n128 VDD2.n127 185
R3076 VDD2.n73 VDD2.n72 185
R3077 VDD2.n122 VDD2.n121 185
R3078 VDD2.n120 VDD2.n119 185
R3079 VDD2.n77 VDD2.n76 185
R3080 VDD2.n114 VDD2.n113 185
R3081 VDD2.n112 VDD2.n79 185
R3082 VDD2.n111 VDD2.n110 185
R3083 VDD2.n82 VDD2.n80 185
R3084 VDD2.n105 VDD2.n104 185
R3085 VDD2.n103 VDD2.n102 185
R3086 VDD2.n86 VDD2.n85 185
R3087 VDD2.n97 VDD2.n96 185
R3088 VDD2.n95 VDD2.n94 185
R3089 VDD2.n90 VDD2.n89 185
R3090 VDD2.n20 VDD2.n19 185
R3091 VDD2.n25 VDD2.n24 185
R3092 VDD2.n27 VDD2.n26 185
R3093 VDD2.n16 VDD2.n15 185
R3094 VDD2.n33 VDD2.n32 185
R3095 VDD2.n35 VDD2.n34 185
R3096 VDD2.n12 VDD2.n11 185
R3097 VDD2.n42 VDD2.n41 185
R3098 VDD2.n43 VDD2.n10 185
R3099 VDD2.n45 VDD2.n44 185
R3100 VDD2.n8 VDD2.n7 185
R3101 VDD2.n51 VDD2.n50 185
R3102 VDD2.n53 VDD2.n52 185
R3103 VDD2.n4 VDD2.n3 185
R3104 VDD2.n59 VDD2.n58 185
R3105 VDD2.n61 VDD2.n60 185
R3106 VDD2.n91 VDD2.t7 149.524
R3107 VDD2.n21 VDD2.t1 149.524
R3108 VDD2.n129 VDD2.n128 104.615
R3109 VDD2.n128 VDD2.n72 104.615
R3110 VDD2.n121 VDD2.n72 104.615
R3111 VDD2.n121 VDD2.n120 104.615
R3112 VDD2.n120 VDD2.n76 104.615
R3113 VDD2.n113 VDD2.n76 104.615
R3114 VDD2.n113 VDD2.n112 104.615
R3115 VDD2.n112 VDD2.n111 104.615
R3116 VDD2.n111 VDD2.n80 104.615
R3117 VDD2.n104 VDD2.n80 104.615
R3118 VDD2.n104 VDD2.n103 104.615
R3119 VDD2.n103 VDD2.n85 104.615
R3120 VDD2.n96 VDD2.n85 104.615
R3121 VDD2.n96 VDD2.n95 104.615
R3122 VDD2.n95 VDD2.n89 104.615
R3123 VDD2.n25 VDD2.n19 104.615
R3124 VDD2.n26 VDD2.n25 104.615
R3125 VDD2.n26 VDD2.n15 104.615
R3126 VDD2.n33 VDD2.n15 104.615
R3127 VDD2.n34 VDD2.n33 104.615
R3128 VDD2.n34 VDD2.n11 104.615
R3129 VDD2.n42 VDD2.n11 104.615
R3130 VDD2.n43 VDD2.n42 104.615
R3131 VDD2.n44 VDD2.n43 104.615
R3132 VDD2.n44 VDD2.n7 104.615
R3133 VDD2.n51 VDD2.n7 104.615
R3134 VDD2.n52 VDD2.n51 104.615
R3135 VDD2.n52 VDD2.n3 104.615
R3136 VDD2.n59 VDD2.n3 104.615
R3137 VDD2.n60 VDD2.n59 104.615
R3138 VDD2.n68 VDD2.n67 65.9169
R3139 VDD2 VDD2.n137 65.914
R3140 VDD2.n136 VDD2.n135 63.6254
R3141 VDD2.n66 VDD2.n65 63.6252
R3142 VDD2.n66 VDD2.n64 53.7389
R3143 VDD2.t7 VDD2.n89 52.3082
R3144 VDD2.t1 VDD2.n19 52.3082
R3145 VDD2.n134 VDD2.n133 50.6096
R3146 VDD2.n134 VDD2.n68 49.1054
R3147 VDD2.n114 VDD2.n79 13.1884
R3148 VDD2.n45 VDD2.n10 13.1884
R3149 VDD2.n115 VDD2.n77 12.8005
R3150 VDD2.n110 VDD2.n81 12.8005
R3151 VDD2.n41 VDD2.n40 12.8005
R3152 VDD2.n46 VDD2.n8 12.8005
R3153 VDD2.n119 VDD2.n118 12.0247
R3154 VDD2.n109 VDD2.n82 12.0247
R3155 VDD2.n39 VDD2.n12 12.0247
R3156 VDD2.n50 VDD2.n49 12.0247
R3157 VDD2.n122 VDD2.n75 11.249
R3158 VDD2.n106 VDD2.n105 11.249
R3159 VDD2.n36 VDD2.n35 11.249
R3160 VDD2.n53 VDD2.n6 11.249
R3161 VDD2.n123 VDD2.n73 10.4732
R3162 VDD2.n102 VDD2.n84 10.4732
R3163 VDD2.n32 VDD2.n14 10.4732
R3164 VDD2.n54 VDD2.n4 10.4732
R3165 VDD2.n91 VDD2.n90 10.2747
R3166 VDD2.n21 VDD2.n20 10.2747
R3167 VDD2.n127 VDD2.n126 9.69747
R3168 VDD2.n101 VDD2.n86 9.69747
R3169 VDD2.n31 VDD2.n16 9.69747
R3170 VDD2.n58 VDD2.n57 9.69747
R3171 VDD2.n133 VDD2.n132 9.45567
R3172 VDD2.n64 VDD2.n63 9.45567
R3173 VDD2.n93 VDD2.n92 9.3005
R3174 VDD2.n88 VDD2.n87 9.3005
R3175 VDD2.n99 VDD2.n98 9.3005
R3176 VDD2.n101 VDD2.n100 9.3005
R3177 VDD2.n84 VDD2.n83 9.3005
R3178 VDD2.n107 VDD2.n106 9.3005
R3179 VDD2.n109 VDD2.n108 9.3005
R3180 VDD2.n81 VDD2.n78 9.3005
R3181 VDD2.n132 VDD2.n131 9.3005
R3182 VDD2.n71 VDD2.n70 9.3005
R3183 VDD2.n126 VDD2.n125 9.3005
R3184 VDD2.n124 VDD2.n123 9.3005
R3185 VDD2.n75 VDD2.n74 9.3005
R3186 VDD2.n118 VDD2.n117 9.3005
R3187 VDD2.n116 VDD2.n115 9.3005
R3188 VDD2.n63 VDD2.n62 9.3005
R3189 VDD2.n2 VDD2.n1 9.3005
R3190 VDD2.n57 VDD2.n56 9.3005
R3191 VDD2.n55 VDD2.n54 9.3005
R3192 VDD2.n6 VDD2.n5 9.3005
R3193 VDD2.n49 VDD2.n48 9.3005
R3194 VDD2.n47 VDD2.n46 9.3005
R3195 VDD2.n23 VDD2.n22 9.3005
R3196 VDD2.n18 VDD2.n17 9.3005
R3197 VDD2.n29 VDD2.n28 9.3005
R3198 VDD2.n31 VDD2.n30 9.3005
R3199 VDD2.n14 VDD2.n13 9.3005
R3200 VDD2.n37 VDD2.n36 9.3005
R3201 VDD2.n39 VDD2.n38 9.3005
R3202 VDD2.n40 VDD2.n9 9.3005
R3203 VDD2.n130 VDD2.n71 8.92171
R3204 VDD2.n98 VDD2.n97 8.92171
R3205 VDD2.n28 VDD2.n27 8.92171
R3206 VDD2.n61 VDD2.n2 8.92171
R3207 VDD2.n131 VDD2.n69 8.14595
R3208 VDD2.n94 VDD2.n88 8.14595
R3209 VDD2.n24 VDD2.n18 8.14595
R3210 VDD2.n62 VDD2.n0 8.14595
R3211 VDD2.n93 VDD2.n90 7.3702
R3212 VDD2.n23 VDD2.n20 7.3702
R3213 VDD2.n133 VDD2.n69 5.81868
R3214 VDD2.n94 VDD2.n93 5.81868
R3215 VDD2.n24 VDD2.n23 5.81868
R3216 VDD2.n64 VDD2.n0 5.81868
R3217 VDD2.n131 VDD2.n130 5.04292
R3218 VDD2.n97 VDD2.n88 5.04292
R3219 VDD2.n27 VDD2.n18 5.04292
R3220 VDD2.n62 VDD2.n61 5.04292
R3221 VDD2.n127 VDD2.n71 4.26717
R3222 VDD2.n98 VDD2.n86 4.26717
R3223 VDD2.n28 VDD2.n16 4.26717
R3224 VDD2.n58 VDD2.n2 4.26717
R3225 VDD2.n126 VDD2.n73 3.49141
R3226 VDD2.n102 VDD2.n101 3.49141
R3227 VDD2.n32 VDD2.n31 3.49141
R3228 VDD2.n57 VDD2.n4 3.49141
R3229 VDD2.n136 VDD2.n134 3.12981
R3230 VDD2.n92 VDD2.n91 2.84303
R3231 VDD2.n22 VDD2.n21 2.84303
R3232 VDD2.n123 VDD2.n122 2.71565
R3233 VDD2.n105 VDD2.n84 2.71565
R3234 VDD2.n35 VDD2.n14 2.71565
R3235 VDD2.n54 VDD2.n53 2.71565
R3236 VDD2.n119 VDD2.n75 1.93989
R3237 VDD2.n106 VDD2.n82 1.93989
R3238 VDD2.n36 VDD2.n12 1.93989
R3239 VDD2.n50 VDD2.n6 1.93989
R3240 VDD2.n137 VDD2.t8 1.62212
R3241 VDD2.n137 VDD2.t2 1.62212
R3242 VDD2.n135 VDD2.t9 1.62212
R3243 VDD2.n135 VDD2.t4 1.62212
R3244 VDD2.n67 VDD2.t5 1.62212
R3245 VDD2.n67 VDD2.t3 1.62212
R3246 VDD2.n65 VDD2.t0 1.62212
R3247 VDD2.n65 VDD2.t6 1.62212
R3248 VDD2.n118 VDD2.n77 1.16414
R3249 VDD2.n110 VDD2.n109 1.16414
R3250 VDD2.n41 VDD2.n39 1.16414
R3251 VDD2.n49 VDD2.n8 1.16414
R3252 VDD2 VDD2.n136 0.841017
R3253 VDD2.n68 VDD2.n66 0.727482
R3254 VDD2.n115 VDD2.n114 0.388379
R3255 VDD2.n81 VDD2.n79 0.388379
R3256 VDD2.n40 VDD2.n10 0.388379
R3257 VDD2.n46 VDD2.n45 0.388379
R3258 VDD2.n132 VDD2.n70 0.155672
R3259 VDD2.n125 VDD2.n70 0.155672
R3260 VDD2.n125 VDD2.n124 0.155672
R3261 VDD2.n124 VDD2.n74 0.155672
R3262 VDD2.n117 VDD2.n74 0.155672
R3263 VDD2.n117 VDD2.n116 0.155672
R3264 VDD2.n116 VDD2.n78 0.155672
R3265 VDD2.n108 VDD2.n78 0.155672
R3266 VDD2.n108 VDD2.n107 0.155672
R3267 VDD2.n107 VDD2.n83 0.155672
R3268 VDD2.n100 VDD2.n83 0.155672
R3269 VDD2.n100 VDD2.n99 0.155672
R3270 VDD2.n99 VDD2.n87 0.155672
R3271 VDD2.n92 VDD2.n87 0.155672
R3272 VDD2.n22 VDD2.n17 0.155672
R3273 VDD2.n29 VDD2.n17 0.155672
R3274 VDD2.n30 VDD2.n29 0.155672
R3275 VDD2.n30 VDD2.n13 0.155672
R3276 VDD2.n37 VDD2.n13 0.155672
R3277 VDD2.n38 VDD2.n37 0.155672
R3278 VDD2.n38 VDD2.n9 0.155672
R3279 VDD2.n47 VDD2.n9 0.155672
R3280 VDD2.n48 VDD2.n47 0.155672
R3281 VDD2.n48 VDD2.n5 0.155672
R3282 VDD2.n55 VDD2.n5 0.155672
R3283 VDD2.n56 VDD2.n55 0.155672
R3284 VDD2.n56 VDD2.n1 0.155672
R3285 VDD2.n63 VDD2.n1 0.155672
C0 VTAIL VDD1 10.765699f
C1 VP VDD1 11.8339f
C2 VN VTAIL 12.2527f
C3 VP VN 9.47175f
C4 VN VDD1 0.154928f
C5 VDD2 VTAIL 10.8219f
C6 VDD2 VP 0.672871f
C7 VDD2 VDD1 2.63015f
C8 VDD2 VN 11.3198f
C9 VP VTAIL 12.266901f
C10 VDD2 B 8.063275f
C11 VDD1 B 8.034097f
C12 VTAIL B 8.829302f
C13 VN B 21.5025f
C14 VP B 20.07196f
C15 VDD2.n0 B 0.035885f
C16 VDD2.n1 B 0.024473f
C17 VDD2.n2 B 0.013151f
C18 VDD2.n3 B 0.031083f
C19 VDD2.n4 B 0.013924f
C20 VDD2.n5 B 0.024473f
C21 VDD2.n6 B 0.013151f
C22 VDD2.n7 B 0.031083f
C23 VDD2.n8 B 0.013924f
C24 VDD2.n9 B 0.024473f
C25 VDD2.n10 B 0.013538f
C26 VDD2.n11 B 0.031083f
C27 VDD2.n12 B 0.013924f
C28 VDD2.n13 B 0.024473f
C29 VDD2.n14 B 0.013151f
C30 VDD2.n15 B 0.031083f
C31 VDD2.n16 B 0.013924f
C32 VDD2.n17 B 0.024473f
C33 VDD2.n18 B 0.013151f
C34 VDD2.n19 B 0.023313f
C35 VDD2.n20 B 0.021974f
C36 VDD2.t1 B 0.052526f
C37 VDD2.n21 B 0.17842f
C38 VDD2.n22 B 1.25748f
C39 VDD2.n23 B 0.013151f
C40 VDD2.n24 B 0.013924f
C41 VDD2.n25 B 0.031083f
C42 VDD2.n26 B 0.031083f
C43 VDD2.n27 B 0.013924f
C44 VDD2.n28 B 0.013151f
C45 VDD2.n29 B 0.024473f
C46 VDD2.n30 B 0.024473f
C47 VDD2.n31 B 0.013151f
C48 VDD2.n32 B 0.013924f
C49 VDD2.n33 B 0.031083f
C50 VDD2.n34 B 0.031083f
C51 VDD2.n35 B 0.013924f
C52 VDD2.n36 B 0.013151f
C53 VDD2.n37 B 0.024473f
C54 VDD2.n38 B 0.024473f
C55 VDD2.n39 B 0.013151f
C56 VDD2.n40 B 0.013151f
C57 VDD2.n41 B 0.013924f
C58 VDD2.n42 B 0.031083f
C59 VDD2.n43 B 0.031083f
C60 VDD2.n44 B 0.031083f
C61 VDD2.n45 B 0.013538f
C62 VDD2.n46 B 0.013151f
C63 VDD2.n47 B 0.024473f
C64 VDD2.n48 B 0.024473f
C65 VDD2.n49 B 0.013151f
C66 VDD2.n50 B 0.013924f
C67 VDD2.n51 B 0.031083f
C68 VDD2.n52 B 0.031083f
C69 VDD2.n53 B 0.013924f
C70 VDD2.n54 B 0.013151f
C71 VDD2.n55 B 0.024473f
C72 VDD2.n56 B 0.024473f
C73 VDD2.n57 B 0.013151f
C74 VDD2.n58 B 0.013924f
C75 VDD2.n59 B 0.031083f
C76 VDD2.n60 B 0.069918f
C77 VDD2.n61 B 0.013924f
C78 VDD2.n62 B 0.013151f
C79 VDD2.n63 B 0.059577f
C80 VDD2.n64 B 0.073572f
C81 VDD2.t0 B 0.236132f
C82 VDD2.t6 B 0.236132f
C83 VDD2.n65 B 2.10783f
C84 VDD2.n66 B 0.784558f
C85 VDD2.t5 B 0.236132f
C86 VDD2.t3 B 0.236132f
C87 VDD2.n67 B 2.13004f
C88 VDD2.n68 B 3.21403f
C89 VDD2.n69 B 0.035885f
C90 VDD2.n70 B 0.024473f
C91 VDD2.n71 B 0.013151f
C92 VDD2.n72 B 0.031083f
C93 VDD2.n73 B 0.013924f
C94 VDD2.n74 B 0.024473f
C95 VDD2.n75 B 0.013151f
C96 VDD2.n76 B 0.031083f
C97 VDD2.n77 B 0.013924f
C98 VDD2.n78 B 0.024473f
C99 VDD2.n79 B 0.013538f
C100 VDD2.n80 B 0.031083f
C101 VDD2.n81 B 0.013151f
C102 VDD2.n82 B 0.013924f
C103 VDD2.n83 B 0.024473f
C104 VDD2.n84 B 0.013151f
C105 VDD2.n85 B 0.031083f
C106 VDD2.n86 B 0.013924f
C107 VDD2.n87 B 0.024473f
C108 VDD2.n88 B 0.013151f
C109 VDD2.n89 B 0.023313f
C110 VDD2.n90 B 0.021974f
C111 VDD2.t7 B 0.052526f
C112 VDD2.n91 B 0.17842f
C113 VDD2.n92 B 1.25748f
C114 VDD2.n93 B 0.013151f
C115 VDD2.n94 B 0.013924f
C116 VDD2.n95 B 0.031083f
C117 VDD2.n96 B 0.031083f
C118 VDD2.n97 B 0.013924f
C119 VDD2.n98 B 0.013151f
C120 VDD2.n99 B 0.024473f
C121 VDD2.n100 B 0.024473f
C122 VDD2.n101 B 0.013151f
C123 VDD2.n102 B 0.013924f
C124 VDD2.n103 B 0.031083f
C125 VDD2.n104 B 0.031083f
C126 VDD2.n105 B 0.013924f
C127 VDD2.n106 B 0.013151f
C128 VDD2.n107 B 0.024473f
C129 VDD2.n108 B 0.024473f
C130 VDD2.n109 B 0.013151f
C131 VDD2.n110 B 0.013924f
C132 VDD2.n111 B 0.031083f
C133 VDD2.n112 B 0.031083f
C134 VDD2.n113 B 0.031083f
C135 VDD2.n114 B 0.013538f
C136 VDD2.n115 B 0.013151f
C137 VDD2.n116 B 0.024473f
C138 VDD2.n117 B 0.024473f
C139 VDD2.n118 B 0.013151f
C140 VDD2.n119 B 0.013924f
C141 VDD2.n120 B 0.031083f
C142 VDD2.n121 B 0.031083f
C143 VDD2.n122 B 0.013924f
C144 VDD2.n123 B 0.013151f
C145 VDD2.n124 B 0.024473f
C146 VDD2.n125 B 0.024473f
C147 VDD2.n126 B 0.013151f
C148 VDD2.n127 B 0.013924f
C149 VDD2.n128 B 0.031083f
C150 VDD2.n129 B 0.069918f
C151 VDD2.n130 B 0.013924f
C152 VDD2.n131 B 0.013151f
C153 VDD2.n132 B 0.059577f
C154 VDD2.n133 B 0.056358f
C155 VDD2.n134 B 3.11389f
C156 VDD2.t9 B 0.236132f
C157 VDD2.t4 B 0.236132f
C158 VDD2.n135 B 2.10784f
C159 VDD2.n136 B 0.514321f
C160 VDD2.t8 B 0.236132f
C161 VDD2.t2 B 0.236132f
C162 VDD2.n137 B 2.13f
C163 VN.t6 B 2.01721f
C164 VN.n0 B 0.778215f
C165 VN.n1 B 0.018365f
C166 VN.n2 B 0.015574f
C167 VN.n3 B 0.018365f
C168 VN.t4 B 2.01721f
C169 VN.n4 B 0.708175f
C170 VN.n5 B 0.018365f
C171 VN.n6 B 0.023486f
C172 VN.n7 B 0.018365f
C173 VN.t3 B 2.01721f
C174 VN.n8 B 0.725505f
C175 VN.n9 B 0.018365f
C176 VN.n10 B 0.023486f
C177 VN.n11 B 0.018365f
C178 VN.t9 B 2.01721f
C179 VN.n12 B 0.765923f
C180 VN.t8 B 2.2417f
C181 VN.n13 B 0.732097f
C182 VN.n14 B 0.216458f
C183 VN.n15 B 0.021723f
C184 VN.n16 B 0.034229f
C185 VN.n17 B 0.034229f
C186 VN.n18 B 0.018365f
C187 VN.n19 B 0.018365f
C188 VN.n20 B 0.018365f
C189 VN.n21 B 0.030139f
C190 VN.n22 B 0.034229f
C191 VN.n23 B 0.034229f
C192 VN.n24 B 0.018365f
C193 VN.n25 B 0.018365f
C194 VN.n26 B 0.018365f
C195 VN.n27 B 0.034229f
C196 VN.n28 B 0.034229f
C197 VN.n29 B 0.030139f
C198 VN.n30 B 0.018365f
C199 VN.n31 B 0.018365f
C200 VN.n32 B 0.018365f
C201 VN.n33 B 0.034229f
C202 VN.n34 B 0.034229f
C203 VN.n35 B 0.021723f
C204 VN.n36 B 0.018365f
C205 VN.n37 B 0.018365f
C206 VN.n38 B 0.029835f
C207 VN.n39 B 0.034229f
C208 VN.n40 B 0.035174f
C209 VN.n41 B 0.018365f
C210 VN.n42 B 0.018365f
C211 VN.n43 B 0.018365f
C212 VN.n44 B 0.037105f
C213 VN.n45 B 0.034229f
C214 VN.n46 B 0.026117f
C215 VN.n47 B 0.029642f
C216 VN.n48 B 0.045832f
C217 VN.t2 B 2.01721f
C218 VN.n49 B 0.778215f
C219 VN.n50 B 0.018365f
C220 VN.n51 B 0.015574f
C221 VN.n52 B 0.018365f
C222 VN.t0 B 2.01721f
C223 VN.n53 B 0.708175f
C224 VN.n54 B 0.018365f
C225 VN.n55 B 0.023486f
C226 VN.n56 B 0.018365f
C227 VN.t5 B 2.01721f
C228 VN.n57 B 0.725505f
C229 VN.n58 B 0.018365f
C230 VN.n59 B 0.023486f
C231 VN.n60 B 0.018365f
C232 VN.t1 B 2.01721f
C233 VN.n61 B 0.765923f
C234 VN.t7 B 2.2417f
C235 VN.n62 B 0.732097f
C236 VN.n63 B 0.216458f
C237 VN.n64 B 0.021723f
C238 VN.n65 B 0.034229f
C239 VN.n66 B 0.034229f
C240 VN.n67 B 0.018365f
C241 VN.n68 B 0.018365f
C242 VN.n69 B 0.018365f
C243 VN.n70 B 0.030139f
C244 VN.n71 B 0.034229f
C245 VN.n72 B 0.034229f
C246 VN.n73 B 0.018365f
C247 VN.n74 B 0.018365f
C248 VN.n75 B 0.018365f
C249 VN.n76 B 0.034229f
C250 VN.n77 B 0.034229f
C251 VN.n78 B 0.030139f
C252 VN.n79 B 0.018365f
C253 VN.n80 B 0.018365f
C254 VN.n81 B 0.018365f
C255 VN.n82 B 0.034229f
C256 VN.n83 B 0.034229f
C257 VN.n84 B 0.021723f
C258 VN.n85 B 0.018365f
C259 VN.n86 B 0.018365f
C260 VN.n87 B 0.029835f
C261 VN.n88 B 0.034229f
C262 VN.n89 B 0.035174f
C263 VN.n90 B 0.018365f
C264 VN.n91 B 0.018365f
C265 VN.n92 B 0.018365f
C266 VN.n93 B 0.037105f
C267 VN.n94 B 0.034229f
C268 VN.n95 B 0.026117f
C269 VN.n96 B 0.029642f
C270 VN.n97 B 1.26785f
C271 VDD1.n0 B 0.036478f
C272 VDD1.n1 B 0.024877f
C273 VDD1.n2 B 0.013368f
C274 VDD1.n3 B 0.031597f
C275 VDD1.n4 B 0.014154f
C276 VDD1.n5 B 0.024877f
C277 VDD1.n6 B 0.013368f
C278 VDD1.n7 B 0.031597f
C279 VDD1.n8 B 0.014154f
C280 VDD1.n9 B 0.024877f
C281 VDD1.n10 B 0.013761f
C282 VDD1.n11 B 0.031597f
C283 VDD1.n12 B 0.013368f
C284 VDD1.n13 B 0.014154f
C285 VDD1.n14 B 0.024877f
C286 VDD1.n15 B 0.013368f
C287 VDD1.n16 B 0.031597f
C288 VDD1.n17 B 0.014154f
C289 VDD1.n18 B 0.024877f
C290 VDD1.n19 B 0.013368f
C291 VDD1.n20 B 0.023698f
C292 VDD1.n21 B 0.022337f
C293 VDD1.t6 B 0.053394f
C294 VDD1.n22 B 0.181368f
C295 VDD1.n23 B 1.27825f
C296 VDD1.n24 B 0.013368f
C297 VDD1.n25 B 0.014154f
C298 VDD1.n26 B 0.031597f
C299 VDD1.n27 B 0.031597f
C300 VDD1.n28 B 0.014154f
C301 VDD1.n29 B 0.013368f
C302 VDD1.n30 B 0.024877f
C303 VDD1.n31 B 0.024877f
C304 VDD1.n32 B 0.013368f
C305 VDD1.n33 B 0.014154f
C306 VDD1.n34 B 0.031597f
C307 VDD1.n35 B 0.031597f
C308 VDD1.n36 B 0.014154f
C309 VDD1.n37 B 0.013368f
C310 VDD1.n38 B 0.024877f
C311 VDD1.n39 B 0.024877f
C312 VDD1.n40 B 0.013368f
C313 VDD1.n41 B 0.014154f
C314 VDD1.n42 B 0.031597f
C315 VDD1.n43 B 0.031597f
C316 VDD1.n44 B 0.031597f
C317 VDD1.n45 B 0.013761f
C318 VDD1.n46 B 0.013368f
C319 VDD1.n47 B 0.024877f
C320 VDD1.n48 B 0.024877f
C321 VDD1.n49 B 0.013368f
C322 VDD1.n50 B 0.014154f
C323 VDD1.n51 B 0.031597f
C324 VDD1.n52 B 0.031597f
C325 VDD1.n53 B 0.014154f
C326 VDD1.n54 B 0.013368f
C327 VDD1.n55 B 0.024877f
C328 VDD1.n56 B 0.024877f
C329 VDD1.n57 B 0.013368f
C330 VDD1.n58 B 0.014154f
C331 VDD1.n59 B 0.031597f
C332 VDD1.n60 B 0.071074f
C333 VDD1.n61 B 0.014154f
C334 VDD1.n62 B 0.013368f
C335 VDD1.n63 B 0.060561f
C336 VDD1.n64 B 0.074788f
C337 VDD1.t3 B 0.240034f
C338 VDD1.t9 B 0.240034f
C339 VDD1.n65 B 2.14266f
C340 VDD1.n66 B 0.805821f
C341 VDD1.n67 B 0.036478f
C342 VDD1.n68 B 0.024877f
C343 VDD1.n69 B 0.013368f
C344 VDD1.n70 B 0.031597f
C345 VDD1.n71 B 0.014154f
C346 VDD1.n72 B 0.024877f
C347 VDD1.n73 B 0.013368f
C348 VDD1.n74 B 0.031597f
C349 VDD1.n75 B 0.014154f
C350 VDD1.n76 B 0.024877f
C351 VDD1.n77 B 0.013761f
C352 VDD1.n78 B 0.031597f
C353 VDD1.n79 B 0.014154f
C354 VDD1.n80 B 0.024877f
C355 VDD1.n81 B 0.013368f
C356 VDD1.n82 B 0.031597f
C357 VDD1.n83 B 0.014154f
C358 VDD1.n84 B 0.024877f
C359 VDD1.n85 B 0.013368f
C360 VDD1.n86 B 0.023698f
C361 VDD1.n87 B 0.022337f
C362 VDD1.t2 B 0.053394f
C363 VDD1.n88 B 0.181368f
C364 VDD1.n89 B 1.27825f
C365 VDD1.n90 B 0.013368f
C366 VDD1.n91 B 0.014154f
C367 VDD1.n92 B 0.031597f
C368 VDD1.n93 B 0.031597f
C369 VDD1.n94 B 0.014154f
C370 VDD1.n95 B 0.013368f
C371 VDD1.n96 B 0.024877f
C372 VDD1.n97 B 0.024877f
C373 VDD1.n98 B 0.013368f
C374 VDD1.n99 B 0.014154f
C375 VDD1.n100 B 0.031597f
C376 VDD1.n101 B 0.031597f
C377 VDD1.n102 B 0.014154f
C378 VDD1.n103 B 0.013368f
C379 VDD1.n104 B 0.024877f
C380 VDD1.n105 B 0.024877f
C381 VDD1.n106 B 0.013368f
C382 VDD1.n107 B 0.013368f
C383 VDD1.n108 B 0.014154f
C384 VDD1.n109 B 0.031597f
C385 VDD1.n110 B 0.031597f
C386 VDD1.n111 B 0.031597f
C387 VDD1.n112 B 0.013761f
C388 VDD1.n113 B 0.013368f
C389 VDD1.n114 B 0.024877f
C390 VDD1.n115 B 0.024877f
C391 VDD1.n116 B 0.013368f
C392 VDD1.n117 B 0.014154f
C393 VDD1.n118 B 0.031597f
C394 VDD1.n119 B 0.031597f
C395 VDD1.n120 B 0.014154f
C396 VDD1.n121 B 0.013368f
C397 VDD1.n122 B 0.024877f
C398 VDD1.n123 B 0.024877f
C399 VDD1.n124 B 0.013368f
C400 VDD1.n125 B 0.014154f
C401 VDD1.n126 B 0.031597f
C402 VDD1.n127 B 0.071074f
C403 VDD1.n128 B 0.014154f
C404 VDD1.n129 B 0.013368f
C405 VDD1.n130 B 0.060561f
C406 VDD1.n131 B 0.074788f
C407 VDD1.t1 B 0.240034f
C408 VDD1.t4 B 0.240034f
C409 VDD1.n132 B 2.14266f
C410 VDD1.n133 B 0.797521f
C411 VDD1.t7 B 0.240034f
C412 VDD1.t8 B 0.240034f
C413 VDD1.n134 B 2.16523f
C414 VDD1.n135 B 3.41078f
C415 VDD1.t5 B 0.240034f
C416 VDD1.t0 B 0.240034f
C417 VDD1.n136 B 2.14266f
C418 VDD1.n137 B 3.46203f
C419 VTAIL.t8 B 0.245789f
C420 VTAIL.t9 B 0.245789f
C421 VTAIL.n0 B 2.12132f
C422 VTAIL.n1 B 0.612015f
C423 VTAIL.n2 B 0.037353f
C424 VTAIL.n3 B 0.025474f
C425 VTAIL.n4 B 0.013689f
C426 VTAIL.n5 B 0.032355f
C427 VTAIL.n6 B 0.014494f
C428 VTAIL.n7 B 0.025474f
C429 VTAIL.n8 B 0.013689f
C430 VTAIL.n9 B 0.032355f
C431 VTAIL.n10 B 0.014494f
C432 VTAIL.n11 B 0.025474f
C433 VTAIL.n12 B 0.014091f
C434 VTAIL.n13 B 0.032355f
C435 VTAIL.n14 B 0.014494f
C436 VTAIL.n15 B 0.025474f
C437 VTAIL.n16 B 0.013689f
C438 VTAIL.n17 B 0.032355f
C439 VTAIL.n18 B 0.014494f
C440 VTAIL.n19 B 0.025474f
C441 VTAIL.n20 B 0.013689f
C442 VTAIL.n21 B 0.024266f
C443 VTAIL.n22 B 0.022872f
C444 VTAIL.t12 B 0.054674f
C445 VTAIL.n23 B 0.185717f
C446 VTAIL.n24 B 1.3089f
C447 VTAIL.n25 B 0.013689f
C448 VTAIL.n26 B 0.014494f
C449 VTAIL.n27 B 0.032355f
C450 VTAIL.n28 B 0.032355f
C451 VTAIL.n29 B 0.014494f
C452 VTAIL.n30 B 0.013689f
C453 VTAIL.n31 B 0.025474f
C454 VTAIL.n32 B 0.025474f
C455 VTAIL.n33 B 0.013689f
C456 VTAIL.n34 B 0.014494f
C457 VTAIL.n35 B 0.032355f
C458 VTAIL.n36 B 0.032355f
C459 VTAIL.n37 B 0.014494f
C460 VTAIL.n38 B 0.013689f
C461 VTAIL.n39 B 0.025474f
C462 VTAIL.n40 B 0.025474f
C463 VTAIL.n41 B 0.013689f
C464 VTAIL.n42 B 0.013689f
C465 VTAIL.n43 B 0.014494f
C466 VTAIL.n44 B 0.032355f
C467 VTAIL.n45 B 0.032355f
C468 VTAIL.n46 B 0.032355f
C469 VTAIL.n47 B 0.014091f
C470 VTAIL.n48 B 0.013689f
C471 VTAIL.n49 B 0.025474f
C472 VTAIL.n50 B 0.025474f
C473 VTAIL.n51 B 0.013689f
C474 VTAIL.n52 B 0.014494f
C475 VTAIL.n53 B 0.032355f
C476 VTAIL.n54 B 0.032355f
C477 VTAIL.n55 B 0.014494f
C478 VTAIL.n56 B 0.013689f
C479 VTAIL.n57 B 0.025474f
C480 VTAIL.n58 B 0.025474f
C481 VTAIL.n59 B 0.013689f
C482 VTAIL.n60 B 0.014494f
C483 VTAIL.n61 B 0.032355f
C484 VTAIL.n62 B 0.072778f
C485 VTAIL.n63 B 0.014494f
C486 VTAIL.n64 B 0.013689f
C487 VTAIL.n65 B 0.062013f
C488 VTAIL.n66 B 0.041097f
C489 VTAIL.n67 B 0.447383f
C490 VTAIL.t13 B 0.245789f
C491 VTAIL.t16 B 0.245789f
C492 VTAIL.n68 B 2.12132f
C493 VTAIL.n69 B 0.76132f
C494 VTAIL.t10 B 0.245789f
C495 VTAIL.t14 B 0.245789f
C496 VTAIL.n70 B 2.12132f
C497 VTAIL.n71 B 2.2282f
C498 VTAIL.t2 B 0.245789f
C499 VTAIL.t7 B 0.245789f
C500 VTAIL.n72 B 2.12133f
C501 VTAIL.n73 B 2.22819f
C502 VTAIL.t5 B 0.245789f
C503 VTAIL.t3 B 0.245789f
C504 VTAIL.n74 B 2.12133f
C505 VTAIL.n75 B 0.761309f
C506 VTAIL.n76 B 0.037353f
C507 VTAIL.n77 B 0.025474f
C508 VTAIL.n78 B 0.013689f
C509 VTAIL.n79 B 0.032355f
C510 VTAIL.n80 B 0.014494f
C511 VTAIL.n81 B 0.025474f
C512 VTAIL.n82 B 0.013689f
C513 VTAIL.n83 B 0.032355f
C514 VTAIL.n84 B 0.014494f
C515 VTAIL.n85 B 0.025474f
C516 VTAIL.n86 B 0.014091f
C517 VTAIL.n87 B 0.032355f
C518 VTAIL.n88 B 0.013689f
C519 VTAIL.n89 B 0.014494f
C520 VTAIL.n90 B 0.025474f
C521 VTAIL.n91 B 0.013689f
C522 VTAIL.n92 B 0.032355f
C523 VTAIL.n93 B 0.014494f
C524 VTAIL.n94 B 0.025474f
C525 VTAIL.n95 B 0.013689f
C526 VTAIL.n96 B 0.024266f
C527 VTAIL.n97 B 0.022872f
C528 VTAIL.t0 B 0.054674f
C529 VTAIL.n98 B 0.185717f
C530 VTAIL.n99 B 1.3089f
C531 VTAIL.n100 B 0.013689f
C532 VTAIL.n101 B 0.014494f
C533 VTAIL.n102 B 0.032355f
C534 VTAIL.n103 B 0.032355f
C535 VTAIL.n104 B 0.014494f
C536 VTAIL.n105 B 0.013689f
C537 VTAIL.n106 B 0.025474f
C538 VTAIL.n107 B 0.025474f
C539 VTAIL.n108 B 0.013689f
C540 VTAIL.n109 B 0.014494f
C541 VTAIL.n110 B 0.032355f
C542 VTAIL.n111 B 0.032355f
C543 VTAIL.n112 B 0.014494f
C544 VTAIL.n113 B 0.013689f
C545 VTAIL.n114 B 0.025474f
C546 VTAIL.n115 B 0.025474f
C547 VTAIL.n116 B 0.013689f
C548 VTAIL.n117 B 0.014494f
C549 VTAIL.n118 B 0.032355f
C550 VTAIL.n119 B 0.032355f
C551 VTAIL.n120 B 0.032355f
C552 VTAIL.n121 B 0.014091f
C553 VTAIL.n122 B 0.013689f
C554 VTAIL.n123 B 0.025474f
C555 VTAIL.n124 B 0.025474f
C556 VTAIL.n125 B 0.013689f
C557 VTAIL.n126 B 0.014494f
C558 VTAIL.n127 B 0.032355f
C559 VTAIL.n128 B 0.032355f
C560 VTAIL.n129 B 0.014494f
C561 VTAIL.n130 B 0.013689f
C562 VTAIL.n131 B 0.025474f
C563 VTAIL.n132 B 0.025474f
C564 VTAIL.n133 B 0.013689f
C565 VTAIL.n134 B 0.014494f
C566 VTAIL.n135 B 0.032355f
C567 VTAIL.n136 B 0.072778f
C568 VTAIL.n137 B 0.014494f
C569 VTAIL.n138 B 0.013689f
C570 VTAIL.n139 B 0.062013f
C571 VTAIL.n140 B 0.041097f
C572 VTAIL.n141 B 0.447383f
C573 VTAIL.t17 B 0.245789f
C574 VTAIL.t15 B 0.245789f
C575 VTAIL.n142 B 2.12133f
C576 VTAIL.n143 B 0.671443f
C577 VTAIL.t11 B 0.245789f
C578 VTAIL.t19 B 0.245789f
C579 VTAIL.n144 B 2.12133f
C580 VTAIL.n145 B 0.761309f
C581 VTAIL.n146 B 0.037353f
C582 VTAIL.n147 B 0.025474f
C583 VTAIL.n148 B 0.013689f
C584 VTAIL.n149 B 0.032355f
C585 VTAIL.n150 B 0.014494f
C586 VTAIL.n151 B 0.025474f
C587 VTAIL.n152 B 0.013689f
C588 VTAIL.n153 B 0.032355f
C589 VTAIL.n154 B 0.014494f
C590 VTAIL.n155 B 0.025474f
C591 VTAIL.n156 B 0.014091f
C592 VTAIL.n157 B 0.032355f
C593 VTAIL.n158 B 0.013689f
C594 VTAIL.n159 B 0.014494f
C595 VTAIL.n160 B 0.025474f
C596 VTAIL.n161 B 0.013689f
C597 VTAIL.n162 B 0.032355f
C598 VTAIL.n163 B 0.014494f
C599 VTAIL.n164 B 0.025474f
C600 VTAIL.n165 B 0.013689f
C601 VTAIL.n166 B 0.024266f
C602 VTAIL.n167 B 0.022872f
C603 VTAIL.t18 B 0.054674f
C604 VTAIL.n168 B 0.185717f
C605 VTAIL.n169 B 1.3089f
C606 VTAIL.n170 B 0.013689f
C607 VTAIL.n171 B 0.014494f
C608 VTAIL.n172 B 0.032355f
C609 VTAIL.n173 B 0.032355f
C610 VTAIL.n174 B 0.014494f
C611 VTAIL.n175 B 0.013689f
C612 VTAIL.n176 B 0.025474f
C613 VTAIL.n177 B 0.025474f
C614 VTAIL.n178 B 0.013689f
C615 VTAIL.n179 B 0.014494f
C616 VTAIL.n180 B 0.032355f
C617 VTAIL.n181 B 0.032355f
C618 VTAIL.n182 B 0.014494f
C619 VTAIL.n183 B 0.013689f
C620 VTAIL.n184 B 0.025474f
C621 VTAIL.n185 B 0.025474f
C622 VTAIL.n186 B 0.013689f
C623 VTAIL.n187 B 0.014494f
C624 VTAIL.n188 B 0.032355f
C625 VTAIL.n189 B 0.032355f
C626 VTAIL.n190 B 0.032355f
C627 VTAIL.n191 B 0.014091f
C628 VTAIL.n192 B 0.013689f
C629 VTAIL.n193 B 0.025474f
C630 VTAIL.n194 B 0.025474f
C631 VTAIL.n195 B 0.013689f
C632 VTAIL.n196 B 0.014494f
C633 VTAIL.n197 B 0.032355f
C634 VTAIL.n198 B 0.032355f
C635 VTAIL.n199 B 0.014494f
C636 VTAIL.n200 B 0.013689f
C637 VTAIL.n201 B 0.025474f
C638 VTAIL.n202 B 0.025474f
C639 VTAIL.n203 B 0.013689f
C640 VTAIL.n204 B 0.014494f
C641 VTAIL.n205 B 0.032355f
C642 VTAIL.n206 B 0.072778f
C643 VTAIL.n207 B 0.014494f
C644 VTAIL.n208 B 0.013689f
C645 VTAIL.n209 B 0.062013f
C646 VTAIL.n210 B 0.041097f
C647 VTAIL.n211 B 1.74727f
C648 VTAIL.n212 B 0.037353f
C649 VTAIL.n213 B 0.025474f
C650 VTAIL.n214 B 0.013689f
C651 VTAIL.n215 B 0.032355f
C652 VTAIL.n216 B 0.014494f
C653 VTAIL.n217 B 0.025474f
C654 VTAIL.n218 B 0.013689f
C655 VTAIL.n219 B 0.032355f
C656 VTAIL.n220 B 0.014494f
C657 VTAIL.n221 B 0.025474f
C658 VTAIL.n222 B 0.014091f
C659 VTAIL.n223 B 0.032355f
C660 VTAIL.n224 B 0.014494f
C661 VTAIL.n225 B 0.025474f
C662 VTAIL.n226 B 0.013689f
C663 VTAIL.n227 B 0.032355f
C664 VTAIL.n228 B 0.014494f
C665 VTAIL.n229 B 0.025474f
C666 VTAIL.n230 B 0.013689f
C667 VTAIL.n231 B 0.024266f
C668 VTAIL.n232 B 0.022872f
C669 VTAIL.t1 B 0.054674f
C670 VTAIL.n233 B 0.185717f
C671 VTAIL.n234 B 1.3089f
C672 VTAIL.n235 B 0.013689f
C673 VTAIL.n236 B 0.014494f
C674 VTAIL.n237 B 0.032355f
C675 VTAIL.n238 B 0.032355f
C676 VTAIL.n239 B 0.014494f
C677 VTAIL.n240 B 0.013689f
C678 VTAIL.n241 B 0.025474f
C679 VTAIL.n242 B 0.025474f
C680 VTAIL.n243 B 0.013689f
C681 VTAIL.n244 B 0.014494f
C682 VTAIL.n245 B 0.032355f
C683 VTAIL.n246 B 0.032355f
C684 VTAIL.n247 B 0.014494f
C685 VTAIL.n248 B 0.013689f
C686 VTAIL.n249 B 0.025474f
C687 VTAIL.n250 B 0.025474f
C688 VTAIL.n251 B 0.013689f
C689 VTAIL.n252 B 0.013689f
C690 VTAIL.n253 B 0.014494f
C691 VTAIL.n254 B 0.032355f
C692 VTAIL.n255 B 0.032355f
C693 VTAIL.n256 B 0.032355f
C694 VTAIL.n257 B 0.014091f
C695 VTAIL.n258 B 0.013689f
C696 VTAIL.n259 B 0.025474f
C697 VTAIL.n260 B 0.025474f
C698 VTAIL.n261 B 0.013689f
C699 VTAIL.n262 B 0.014494f
C700 VTAIL.n263 B 0.032355f
C701 VTAIL.n264 B 0.032355f
C702 VTAIL.n265 B 0.014494f
C703 VTAIL.n266 B 0.013689f
C704 VTAIL.n267 B 0.025474f
C705 VTAIL.n268 B 0.025474f
C706 VTAIL.n269 B 0.013689f
C707 VTAIL.n270 B 0.014494f
C708 VTAIL.n271 B 0.032355f
C709 VTAIL.n272 B 0.072778f
C710 VTAIL.n273 B 0.014494f
C711 VTAIL.n274 B 0.013689f
C712 VTAIL.n275 B 0.062013f
C713 VTAIL.n276 B 0.041097f
C714 VTAIL.n277 B 1.74727f
C715 VTAIL.t6 B 0.245789f
C716 VTAIL.t4 B 0.245789f
C717 VTAIL.n278 B 2.12132f
C718 VTAIL.n279 B 0.563898f
C719 VP.t1 B 2.04928f
C720 VP.n0 B 0.790587f
C721 VP.n1 B 0.018657f
C722 VP.n2 B 0.015821f
C723 VP.n3 B 0.018657f
C724 VP.t2 B 2.04928f
C725 VP.n4 B 0.719433f
C726 VP.n5 B 0.018657f
C727 VP.n6 B 0.023859f
C728 VP.n7 B 0.018657f
C729 VP.t5 B 2.04928f
C730 VP.n8 B 0.737039f
C731 VP.n9 B 0.018657f
C732 VP.n10 B 0.023859f
C733 VP.n11 B 0.018657f
C734 VP.t8 B 2.04928f
C735 VP.n12 B 0.719433f
C736 VP.n13 B 0.018657f
C737 VP.n14 B 0.015821f
C738 VP.n15 B 0.018657f
C739 VP.t7 B 2.04928f
C740 VP.n16 B 0.790587f
C741 VP.t9 B 2.04928f
C742 VP.n17 B 0.790587f
C743 VP.n18 B 0.018657f
C744 VP.n19 B 0.015821f
C745 VP.n20 B 0.018657f
C746 VP.t4 B 2.04928f
C747 VP.n21 B 0.719433f
C748 VP.n22 B 0.018657f
C749 VP.n23 B 0.023859f
C750 VP.n24 B 0.018657f
C751 VP.t0 B 2.04928f
C752 VP.n25 B 0.737039f
C753 VP.n26 B 0.018657f
C754 VP.n27 B 0.023859f
C755 VP.n28 B 0.018657f
C756 VP.t6 B 2.04928f
C757 VP.n29 B 0.7781f
C758 VP.t3 B 2.27734f
C759 VP.n30 B 0.743737f
C760 VP.n31 B 0.2199f
C761 VP.n32 B 0.022069f
C762 VP.n33 B 0.034773f
C763 VP.n34 B 0.034773f
C764 VP.n35 B 0.018657f
C765 VP.n36 B 0.018657f
C766 VP.n37 B 0.018657f
C767 VP.n38 B 0.030618f
C768 VP.n39 B 0.034773f
C769 VP.n40 B 0.034773f
C770 VP.n41 B 0.018657f
C771 VP.n42 B 0.018657f
C772 VP.n43 B 0.018657f
C773 VP.n44 B 0.034773f
C774 VP.n45 B 0.034773f
C775 VP.n46 B 0.030618f
C776 VP.n47 B 0.018657f
C777 VP.n48 B 0.018657f
C778 VP.n49 B 0.018657f
C779 VP.n50 B 0.034773f
C780 VP.n51 B 0.034773f
C781 VP.n52 B 0.022069f
C782 VP.n53 B 0.018657f
C783 VP.n54 B 0.018657f
C784 VP.n55 B 0.030309f
C785 VP.n56 B 0.034773f
C786 VP.n57 B 0.035733f
C787 VP.n58 B 0.018657f
C788 VP.n59 B 0.018657f
C789 VP.n60 B 0.018657f
C790 VP.n61 B 0.037695f
C791 VP.n62 B 0.034773f
C792 VP.n63 B 0.026532f
C793 VP.n64 B 0.030113f
C794 VP.n65 B 1.2807f
C795 VP.n66 B 1.29243f
C796 VP.n67 B 0.030113f
C797 VP.n68 B 0.026532f
C798 VP.n69 B 0.034773f
C799 VP.n70 B 0.037695f
C800 VP.n71 B 0.018657f
C801 VP.n72 B 0.018657f
C802 VP.n73 B 0.018657f
C803 VP.n74 B 0.035733f
C804 VP.n75 B 0.034773f
C805 VP.n76 B 0.030309f
C806 VP.n77 B 0.018657f
C807 VP.n78 B 0.018657f
C808 VP.n79 B 0.022069f
C809 VP.n80 B 0.034773f
C810 VP.n81 B 0.034773f
C811 VP.n82 B 0.018657f
C812 VP.n83 B 0.018657f
C813 VP.n84 B 0.018657f
C814 VP.n85 B 0.030618f
C815 VP.n86 B 0.034773f
C816 VP.n87 B 0.034773f
C817 VP.n88 B 0.018657f
C818 VP.n89 B 0.018657f
C819 VP.n90 B 0.018657f
C820 VP.n91 B 0.034773f
C821 VP.n92 B 0.034773f
C822 VP.n93 B 0.030618f
C823 VP.n94 B 0.018657f
C824 VP.n95 B 0.018657f
C825 VP.n96 B 0.018657f
C826 VP.n97 B 0.034773f
C827 VP.n98 B 0.034773f
C828 VP.n99 B 0.022069f
C829 VP.n100 B 0.018657f
C830 VP.n101 B 0.018657f
C831 VP.n102 B 0.030309f
C832 VP.n103 B 0.034773f
C833 VP.n104 B 0.035733f
C834 VP.n105 B 0.018657f
C835 VP.n106 B 0.018657f
C836 VP.n107 B 0.018657f
C837 VP.n108 B 0.037695f
C838 VP.n109 B 0.034773f
C839 VP.n110 B 0.026532f
C840 VP.n111 B 0.030113f
C841 VP.n112 B 0.04656f
.ends

