* NGSPICE file created from diff_pair_sample_0092.ext - technology: sky130A

.subckt diff_pair_sample_0092 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=2.82645 ps=17.46 w=17.13 l=1.99
X1 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=2.82645 ps=17.46 w=17.13 l=1.99
X2 VDD1.t4 VP.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=6.6807 ps=35.04 w=17.13 l=1.99
X3 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=6.6807 ps=35.04 w=17.13 l=1.99
X4 VTAIL.t6 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=2.82645 ps=17.46 w=17.13 l=1.99
X5 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=2.82645 ps=17.46 w=17.13 l=1.99
X6 VDD1.t2 VP.t3 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=2.82645 ps=17.46 w=17.13 l=1.99
X7 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=0 ps=0 w=17.13 l=1.99
X8 VDD1.t1 VP.t4 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=6.6807 ps=35.04 w=17.13 l=1.99
X9 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=0 ps=0 w=17.13 l=1.99
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=0 ps=0 w=17.13 l=1.99
X11 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=6.6807 ps=35.04 w=17.13 l=1.99
X12 VTAIL.t10 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=2.82645 ps=17.46 w=17.13 l=1.99
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=0 ps=0 w=17.13 l=1.99
X14 VTAIL.t11 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.82645 pd=17.46 as=2.82645 ps=17.46 w=17.13 l=1.99
X15 VDD2.t0 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6807 pd=35.04 as=2.82645 ps=17.46 w=17.13 l=1.99
R0 VP.n7 VP.t0 240.774
R1 VP.n25 VP.t5 207.454
R2 VP.n18 VP.t3 207.454
R3 VP.n32 VP.t4 207.454
R4 VP.n8 VP.t2 207.454
R5 VP.n15 VP.t1 207.454
R6 VP.n10 VP.n9 161.3
R7 VP.n11 VP.n6 161.3
R8 VP.n13 VP.n12 161.3
R9 VP.n14 VP.n5 161.3
R10 VP.n31 VP.n0 161.3
R11 VP.n30 VP.n29 161.3
R12 VP.n28 VP.n1 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n25 VP.n2 161.3
R15 VP.n24 VP.n23 161.3
R16 VP.n22 VP.n3 161.3
R17 VP.n21 VP.n20 161.3
R18 VP.n19 VP.n4 161.3
R19 VP.n18 VP.n17 95.0976
R20 VP.n33 VP.n32 95.0976
R21 VP.n16 VP.n15 95.0976
R22 VP.n20 VP.n3 56.0336
R23 VP.n30 VP.n1 56.0336
R24 VP.n13 VP.n6 56.0336
R25 VP.n17 VP.n16 50.1284
R26 VP.n8 VP.n7 45.7215
R27 VP.n24 VP.n3 24.9531
R28 VP.n26 VP.n1 24.9531
R29 VP.n9 VP.n6 24.9531
R30 VP.n20 VP.n19 24.4675
R31 VP.n25 VP.n24 24.4675
R32 VP.n26 VP.n25 24.4675
R33 VP.n31 VP.n30 24.4675
R34 VP.n14 VP.n13 24.4675
R35 VP.n9 VP.n8 24.4675
R36 VP.n19 VP.n18 15.6594
R37 VP.n32 VP.n31 15.6594
R38 VP.n15 VP.n14 15.6594
R39 VP.n10 VP.n7 9.37527
R40 VP.n16 VP.n5 0.278367
R41 VP.n17 VP.n4 0.278367
R42 VP.n33 VP.n0 0.278367
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153454
R55 VTAIL.n7 VTAIL.t3 44.5973
R56 VTAIL.n11 VTAIL.t2 44.5971
R57 VTAIL.n2 VTAIL.t9 44.5971
R58 VTAIL.n10 VTAIL.t5 44.5971
R59 VTAIL.n9 VTAIL.n8 43.4415
R60 VTAIL.n6 VTAIL.n5 43.4415
R61 VTAIL.n1 VTAIL.n0 43.4412
R62 VTAIL.n4 VTAIL.n3 43.4412
R63 VTAIL.n6 VTAIL.n4 31.1341
R64 VTAIL.n11 VTAIL.n10 29.1341
R65 VTAIL.n7 VTAIL.n6 2.0005
R66 VTAIL.n10 VTAIL.n9 2.0005
R67 VTAIL.n4 VTAIL.n2 2.0005
R68 VTAIL.n9 VTAIL.n7 1.47033
R69 VTAIL.n2 VTAIL.n1 1.47033
R70 VTAIL VTAIL.n11 1.44231
R71 VTAIL.n0 VTAIL.t1 1.15637
R72 VTAIL.n0 VTAIL.t0 1.15637
R73 VTAIL.n3 VTAIL.t7 1.15637
R74 VTAIL.n3 VTAIL.t10 1.15637
R75 VTAIL.n8 VTAIL.t8 1.15637
R76 VTAIL.n8 VTAIL.t6 1.15637
R77 VTAIL.n5 VTAIL.t4 1.15637
R78 VTAIL.n5 VTAIL.t11 1.15637
R79 VTAIL VTAIL.n1 0.55869
R80 VDD1 VDD1.t5 62.8342
R81 VDD1.n1 VDD1.t2 62.7206
R82 VDD1.n1 VDD1.n0 60.5647
R83 VDD1.n3 VDD1.n2 60.1201
R84 VDD1.n3 VDD1.n1 46.5655
R85 VDD1.n2 VDD1.t3 1.15637
R86 VDD1.n2 VDD1.t4 1.15637
R87 VDD1.n0 VDD1.t0 1.15637
R88 VDD1.n0 VDD1.t1 1.15637
R89 VDD1 VDD1.n3 0.44231
R90 B.n909 B.n908 585
R91 B.n910 B.n909 585
R92 B.n375 B.n129 585
R93 B.n374 B.n373 585
R94 B.n372 B.n371 585
R95 B.n370 B.n369 585
R96 B.n368 B.n367 585
R97 B.n366 B.n365 585
R98 B.n364 B.n363 585
R99 B.n362 B.n361 585
R100 B.n360 B.n359 585
R101 B.n358 B.n357 585
R102 B.n356 B.n355 585
R103 B.n354 B.n353 585
R104 B.n352 B.n351 585
R105 B.n350 B.n349 585
R106 B.n348 B.n347 585
R107 B.n346 B.n345 585
R108 B.n344 B.n343 585
R109 B.n342 B.n341 585
R110 B.n340 B.n339 585
R111 B.n338 B.n337 585
R112 B.n336 B.n335 585
R113 B.n334 B.n333 585
R114 B.n332 B.n331 585
R115 B.n330 B.n329 585
R116 B.n328 B.n327 585
R117 B.n326 B.n325 585
R118 B.n324 B.n323 585
R119 B.n322 B.n321 585
R120 B.n320 B.n319 585
R121 B.n318 B.n317 585
R122 B.n316 B.n315 585
R123 B.n314 B.n313 585
R124 B.n312 B.n311 585
R125 B.n310 B.n309 585
R126 B.n308 B.n307 585
R127 B.n306 B.n305 585
R128 B.n304 B.n303 585
R129 B.n302 B.n301 585
R130 B.n300 B.n299 585
R131 B.n298 B.n297 585
R132 B.n296 B.n295 585
R133 B.n294 B.n293 585
R134 B.n292 B.n291 585
R135 B.n290 B.n289 585
R136 B.n288 B.n287 585
R137 B.n286 B.n285 585
R138 B.n284 B.n283 585
R139 B.n282 B.n281 585
R140 B.n280 B.n279 585
R141 B.n278 B.n277 585
R142 B.n276 B.n275 585
R143 B.n274 B.n273 585
R144 B.n272 B.n271 585
R145 B.n270 B.n269 585
R146 B.n268 B.n267 585
R147 B.n266 B.n265 585
R148 B.n264 B.n263 585
R149 B.n262 B.n261 585
R150 B.n260 B.n259 585
R151 B.n258 B.n257 585
R152 B.n256 B.n255 585
R153 B.n254 B.n253 585
R154 B.n252 B.n251 585
R155 B.n250 B.n249 585
R156 B.n248 B.n247 585
R157 B.n245 B.n244 585
R158 B.n243 B.n242 585
R159 B.n241 B.n240 585
R160 B.n239 B.n238 585
R161 B.n237 B.n236 585
R162 B.n235 B.n234 585
R163 B.n233 B.n232 585
R164 B.n231 B.n230 585
R165 B.n229 B.n228 585
R166 B.n227 B.n226 585
R167 B.n225 B.n224 585
R168 B.n223 B.n222 585
R169 B.n221 B.n220 585
R170 B.n219 B.n218 585
R171 B.n217 B.n216 585
R172 B.n215 B.n214 585
R173 B.n213 B.n212 585
R174 B.n211 B.n210 585
R175 B.n209 B.n208 585
R176 B.n207 B.n206 585
R177 B.n205 B.n204 585
R178 B.n203 B.n202 585
R179 B.n201 B.n200 585
R180 B.n199 B.n198 585
R181 B.n197 B.n196 585
R182 B.n195 B.n194 585
R183 B.n193 B.n192 585
R184 B.n191 B.n190 585
R185 B.n189 B.n188 585
R186 B.n187 B.n186 585
R187 B.n185 B.n184 585
R188 B.n183 B.n182 585
R189 B.n181 B.n180 585
R190 B.n179 B.n178 585
R191 B.n177 B.n176 585
R192 B.n175 B.n174 585
R193 B.n173 B.n172 585
R194 B.n171 B.n170 585
R195 B.n169 B.n168 585
R196 B.n167 B.n166 585
R197 B.n165 B.n164 585
R198 B.n163 B.n162 585
R199 B.n161 B.n160 585
R200 B.n159 B.n158 585
R201 B.n157 B.n156 585
R202 B.n155 B.n154 585
R203 B.n153 B.n152 585
R204 B.n151 B.n150 585
R205 B.n149 B.n148 585
R206 B.n147 B.n146 585
R207 B.n145 B.n144 585
R208 B.n143 B.n142 585
R209 B.n141 B.n140 585
R210 B.n139 B.n138 585
R211 B.n137 B.n136 585
R212 B.n68 B.n67 585
R213 B.n913 B.n912 585
R214 B.n907 B.n130 585
R215 B.n130 B.n65 585
R216 B.n906 B.n64 585
R217 B.n917 B.n64 585
R218 B.n905 B.n63 585
R219 B.n918 B.n63 585
R220 B.n904 B.n62 585
R221 B.n919 B.n62 585
R222 B.n903 B.n902 585
R223 B.n902 B.n58 585
R224 B.n901 B.n57 585
R225 B.n925 B.n57 585
R226 B.n900 B.n56 585
R227 B.n926 B.n56 585
R228 B.n899 B.n55 585
R229 B.n927 B.n55 585
R230 B.n898 B.n897 585
R231 B.n897 B.n51 585
R232 B.n896 B.n50 585
R233 B.n933 B.n50 585
R234 B.n895 B.n49 585
R235 B.n934 B.n49 585
R236 B.n894 B.n48 585
R237 B.n935 B.n48 585
R238 B.n893 B.n892 585
R239 B.n892 B.n44 585
R240 B.n891 B.n43 585
R241 B.n941 B.n43 585
R242 B.n890 B.n42 585
R243 B.n942 B.n42 585
R244 B.n889 B.n41 585
R245 B.n943 B.n41 585
R246 B.n888 B.n887 585
R247 B.n887 B.n40 585
R248 B.n886 B.n36 585
R249 B.n949 B.n36 585
R250 B.n885 B.n35 585
R251 B.n950 B.n35 585
R252 B.n884 B.n34 585
R253 B.n951 B.n34 585
R254 B.n883 B.n882 585
R255 B.n882 B.n30 585
R256 B.n881 B.n29 585
R257 B.n957 B.n29 585
R258 B.n880 B.n28 585
R259 B.n958 B.n28 585
R260 B.n879 B.n27 585
R261 B.n959 B.n27 585
R262 B.n878 B.n877 585
R263 B.n877 B.n23 585
R264 B.n876 B.n22 585
R265 B.n965 B.n22 585
R266 B.n875 B.n21 585
R267 B.n966 B.n21 585
R268 B.n874 B.n20 585
R269 B.n967 B.n20 585
R270 B.n873 B.n872 585
R271 B.n872 B.n16 585
R272 B.n871 B.n15 585
R273 B.n973 B.n15 585
R274 B.n870 B.n14 585
R275 B.n974 B.n14 585
R276 B.n869 B.n13 585
R277 B.n975 B.n13 585
R278 B.n868 B.n867 585
R279 B.n867 B.n12 585
R280 B.n866 B.n865 585
R281 B.n866 B.n8 585
R282 B.n864 B.n7 585
R283 B.n982 B.n7 585
R284 B.n863 B.n6 585
R285 B.n983 B.n6 585
R286 B.n862 B.n5 585
R287 B.n984 B.n5 585
R288 B.n861 B.n860 585
R289 B.n860 B.n4 585
R290 B.n859 B.n376 585
R291 B.n859 B.n858 585
R292 B.n849 B.n377 585
R293 B.n378 B.n377 585
R294 B.n851 B.n850 585
R295 B.n852 B.n851 585
R296 B.n848 B.n382 585
R297 B.n386 B.n382 585
R298 B.n847 B.n846 585
R299 B.n846 B.n845 585
R300 B.n384 B.n383 585
R301 B.n385 B.n384 585
R302 B.n838 B.n837 585
R303 B.n839 B.n838 585
R304 B.n836 B.n391 585
R305 B.n391 B.n390 585
R306 B.n835 B.n834 585
R307 B.n834 B.n833 585
R308 B.n393 B.n392 585
R309 B.n394 B.n393 585
R310 B.n826 B.n825 585
R311 B.n827 B.n826 585
R312 B.n824 B.n399 585
R313 B.n399 B.n398 585
R314 B.n823 B.n822 585
R315 B.n822 B.n821 585
R316 B.n401 B.n400 585
R317 B.n402 B.n401 585
R318 B.n814 B.n813 585
R319 B.n815 B.n814 585
R320 B.n812 B.n407 585
R321 B.n407 B.n406 585
R322 B.n811 B.n810 585
R323 B.n810 B.n809 585
R324 B.n409 B.n408 585
R325 B.n802 B.n409 585
R326 B.n801 B.n800 585
R327 B.n803 B.n801 585
R328 B.n799 B.n414 585
R329 B.n414 B.n413 585
R330 B.n798 B.n797 585
R331 B.n797 B.n796 585
R332 B.n416 B.n415 585
R333 B.n417 B.n416 585
R334 B.n789 B.n788 585
R335 B.n790 B.n789 585
R336 B.n787 B.n422 585
R337 B.n422 B.n421 585
R338 B.n786 B.n785 585
R339 B.n785 B.n784 585
R340 B.n424 B.n423 585
R341 B.n425 B.n424 585
R342 B.n777 B.n776 585
R343 B.n778 B.n777 585
R344 B.n775 B.n429 585
R345 B.n433 B.n429 585
R346 B.n774 B.n773 585
R347 B.n773 B.n772 585
R348 B.n431 B.n430 585
R349 B.n432 B.n431 585
R350 B.n765 B.n764 585
R351 B.n766 B.n765 585
R352 B.n763 B.n438 585
R353 B.n438 B.n437 585
R354 B.n762 B.n761 585
R355 B.n761 B.n760 585
R356 B.n440 B.n439 585
R357 B.n441 B.n440 585
R358 B.n756 B.n755 585
R359 B.n444 B.n443 585
R360 B.n752 B.n751 585
R361 B.n753 B.n752 585
R362 B.n750 B.n505 585
R363 B.n749 B.n748 585
R364 B.n747 B.n746 585
R365 B.n745 B.n744 585
R366 B.n743 B.n742 585
R367 B.n741 B.n740 585
R368 B.n739 B.n738 585
R369 B.n737 B.n736 585
R370 B.n735 B.n734 585
R371 B.n733 B.n732 585
R372 B.n731 B.n730 585
R373 B.n729 B.n728 585
R374 B.n727 B.n726 585
R375 B.n725 B.n724 585
R376 B.n723 B.n722 585
R377 B.n721 B.n720 585
R378 B.n719 B.n718 585
R379 B.n717 B.n716 585
R380 B.n715 B.n714 585
R381 B.n713 B.n712 585
R382 B.n711 B.n710 585
R383 B.n709 B.n708 585
R384 B.n707 B.n706 585
R385 B.n705 B.n704 585
R386 B.n703 B.n702 585
R387 B.n701 B.n700 585
R388 B.n699 B.n698 585
R389 B.n697 B.n696 585
R390 B.n695 B.n694 585
R391 B.n693 B.n692 585
R392 B.n691 B.n690 585
R393 B.n689 B.n688 585
R394 B.n687 B.n686 585
R395 B.n685 B.n684 585
R396 B.n683 B.n682 585
R397 B.n681 B.n680 585
R398 B.n679 B.n678 585
R399 B.n677 B.n676 585
R400 B.n675 B.n674 585
R401 B.n673 B.n672 585
R402 B.n671 B.n670 585
R403 B.n669 B.n668 585
R404 B.n667 B.n666 585
R405 B.n665 B.n664 585
R406 B.n663 B.n662 585
R407 B.n661 B.n660 585
R408 B.n659 B.n658 585
R409 B.n657 B.n656 585
R410 B.n655 B.n654 585
R411 B.n653 B.n652 585
R412 B.n651 B.n650 585
R413 B.n649 B.n648 585
R414 B.n647 B.n646 585
R415 B.n645 B.n644 585
R416 B.n643 B.n642 585
R417 B.n641 B.n640 585
R418 B.n639 B.n638 585
R419 B.n637 B.n636 585
R420 B.n635 B.n634 585
R421 B.n633 B.n632 585
R422 B.n631 B.n630 585
R423 B.n629 B.n628 585
R424 B.n627 B.n626 585
R425 B.n624 B.n623 585
R426 B.n622 B.n621 585
R427 B.n620 B.n619 585
R428 B.n618 B.n617 585
R429 B.n616 B.n615 585
R430 B.n614 B.n613 585
R431 B.n612 B.n611 585
R432 B.n610 B.n609 585
R433 B.n608 B.n607 585
R434 B.n606 B.n605 585
R435 B.n604 B.n603 585
R436 B.n602 B.n601 585
R437 B.n600 B.n599 585
R438 B.n598 B.n597 585
R439 B.n596 B.n595 585
R440 B.n594 B.n593 585
R441 B.n592 B.n591 585
R442 B.n590 B.n589 585
R443 B.n588 B.n587 585
R444 B.n586 B.n585 585
R445 B.n584 B.n583 585
R446 B.n582 B.n581 585
R447 B.n580 B.n579 585
R448 B.n578 B.n577 585
R449 B.n576 B.n575 585
R450 B.n574 B.n573 585
R451 B.n572 B.n571 585
R452 B.n570 B.n569 585
R453 B.n568 B.n567 585
R454 B.n566 B.n565 585
R455 B.n564 B.n563 585
R456 B.n562 B.n561 585
R457 B.n560 B.n559 585
R458 B.n558 B.n557 585
R459 B.n556 B.n555 585
R460 B.n554 B.n553 585
R461 B.n552 B.n551 585
R462 B.n550 B.n549 585
R463 B.n548 B.n547 585
R464 B.n546 B.n545 585
R465 B.n544 B.n543 585
R466 B.n542 B.n541 585
R467 B.n540 B.n539 585
R468 B.n538 B.n537 585
R469 B.n536 B.n535 585
R470 B.n534 B.n533 585
R471 B.n532 B.n531 585
R472 B.n530 B.n529 585
R473 B.n528 B.n527 585
R474 B.n526 B.n525 585
R475 B.n524 B.n523 585
R476 B.n522 B.n521 585
R477 B.n520 B.n519 585
R478 B.n518 B.n517 585
R479 B.n516 B.n515 585
R480 B.n514 B.n513 585
R481 B.n512 B.n511 585
R482 B.n757 B.n442 585
R483 B.n442 B.n441 585
R484 B.n759 B.n758 585
R485 B.n760 B.n759 585
R486 B.n436 B.n435 585
R487 B.n437 B.n436 585
R488 B.n768 B.n767 585
R489 B.n767 B.n766 585
R490 B.n769 B.n434 585
R491 B.n434 B.n432 585
R492 B.n771 B.n770 585
R493 B.n772 B.n771 585
R494 B.n428 B.n427 585
R495 B.n433 B.n428 585
R496 B.n780 B.n779 585
R497 B.n779 B.n778 585
R498 B.n781 B.n426 585
R499 B.n426 B.n425 585
R500 B.n783 B.n782 585
R501 B.n784 B.n783 585
R502 B.n420 B.n419 585
R503 B.n421 B.n420 585
R504 B.n792 B.n791 585
R505 B.n791 B.n790 585
R506 B.n793 B.n418 585
R507 B.n418 B.n417 585
R508 B.n795 B.n794 585
R509 B.n796 B.n795 585
R510 B.n412 B.n411 585
R511 B.n413 B.n412 585
R512 B.n805 B.n804 585
R513 B.n804 B.n803 585
R514 B.n806 B.n410 585
R515 B.n802 B.n410 585
R516 B.n808 B.n807 585
R517 B.n809 B.n808 585
R518 B.n405 B.n404 585
R519 B.n406 B.n405 585
R520 B.n817 B.n816 585
R521 B.n816 B.n815 585
R522 B.n818 B.n403 585
R523 B.n403 B.n402 585
R524 B.n820 B.n819 585
R525 B.n821 B.n820 585
R526 B.n397 B.n396 585
R527 B.n398 B.n397 585
R528 B.n829 B.n828 585
R529 B.n828 B.n827 585
R530 B.n830 B.n395 585
R531 B.n395 B.n394 585
R532 B.n832 B.n831 585
R533 B.n833 B.n832 585
R534 B.n389 B.n388 585
R535 B.n390 B.n389 585
R536 B.n841 B.n840 585
R537 B.n840 B.n839 585
R538 B.n842 B.n387 585
R539 B.n387 B.n385 585
R540 B.n844 B.n843 585
R541 B.n845 B.n844 585
R542 B.n381 B.n380 585
R543 B.n386 B.n381 585
R544 B.n854 B.n853 585
R545 B.n853 B.n852 585
R546 B.n855 B.n379 585
R547 B.n379 B.n378 585
R548 B.n857 B.n856 585
R549 B.n858 B.n857 585
R550 B.n3 B.n0 585
R551 B.n4 B.n3 585
R552 B.n981 B.n1 585
R553 B.n982 B.n981 585
R554 B.n980 B.n979 585
R555 B.n980 B.n8 585
R556 B.n978 B.n9 585
R557 B.n12 B.n9 585
R558 B.n977 B.n976 585
R559 B.n976 B.n975 585
R560 B.n11 B.n10 585
R561 B.n974 B.n11 585
R562 B.n972 B.n971 585
R563 B.n973 B.n972 585
R564 B.n970 B.n17 585
R565 B.n17 B.n16 585
R566 B.n969 B.n968 585
R567 B.n968 B.n967 585
R568 B.n19 B.n18 585
R569 B.n966 B.n19 585
R570 B.n964 B.n963 585
R571 B.n965 B.n964 585
R572 B.n962 B.n24 585
R573 B.n24 B.n23 585
R574 B.n961 B.n960 585
R575 B.n960 B.n959 585
R576 B.n26 B.n25 585
R577 B.n958 B.n26 585
R578 B.n956 B.n955 585
R579 B.n957 B.n956 585
R580 B.n954 B.n31 585
R581 B.n31 B.n30 585
R582 B.n953 B.n952 585
R583 B.n952 B.n951 585
R584 B.n33 B.n32 585
R585 B.n950 B.n33 585
R586 B.n948 B.n947 585
R587 B.n949 B.n948 585
R588 B.n946 B.n37 585
R589 B.n40 B.n37 585
R590 B.n945 B.n944 585
R591 B.n944 B.n943 585
R592 B.n39 B.n38 585
R593 B.n942 B.n39 585
R594 B.n940 B.n939 585
R595 B.n941 B.n940 585
R596 B.n938 B.n45 585
R597 B.n45 B.n44 585
R598 B.n937 B.n936 585
R599 B.n936 B.n935 585
R600 B.n47 B.n46 585
R601 B.n934 B.n47 585
R602 B.n932 B.n931 585
R603 B.n933 B.n932 585
R604 B.n930 B.n52 585
R605 B.n52 B.n51 585
R606 B.n929 B.n928 585
R607 B.n928 B.n927 585
R608 B.n54 B.n53 585
R609 B.n926 B.n54 585
R610 B.n924 B.n923 585
R611 B.n925 B.n924 585
R612 B.n922 B.n59 585
R613 B.n59 B.n58 585
R614 B.n921 B.n920 585
R615 B.n920 B.n919 585
R616 B.n61 B.n60 585
R617 B.n918 B.n61 585
R618 B.n916 B.n915 585
R619 B.n917 B.n916 585
R620 B.n914 B.n66 585
R621 B.n66 B.n65 585
R622 B.n985 B.n984 585
R623 B.n983 B.n2 585
R624 B.n912 B.n66 482.89
R625 B.n909 B.n130 482.89
R626 B.n511 B.n440 482.89
R627 B.n755 B.n442 482.89
R628 B.n134 B.t10 414.349
R629 B.n131 B.t17 414.349
R630 B.n509 B.t14 414.349
R631 B.n506 B.t6 414.349
R632 B.n910 B.n128 256.663
R633 B.n910 B.n127 256.663
R634 B.n910 B.n126 256.663
R635 B.n910 B.n125 256.663
R636 B.n910 B.n124 256.663
R637 B.n910 B.n123 256.663
R638 B.n910 B.n122 256.663
R639 B.n910 B.n121 256.663
R640 B.n910 B.n120 256.663
R641 B.n910 B.n119 256.663
R642 B.n910 B.n118 256.663
R643 B.n910 B.n117 256.663
R644 B.n910 B.n116 256.663
R645 B.n910 B.n115 256.663
R646 B.n910 B.n114 256.663
R647 B.n910 B.n113 256.663
R648 B.n910 B.n112 256.663
R649 B.n910 B.n111 256.663
R650 B.n910 B.n110 256.663
R651 B.n910 B.n109 256.663
R652 B.n910 B.n108 256.663
R653 B.n910 B.n107 256.663
R654 B.n910 B.n106 256.663
R655 B.n910 B.n105 256.663
R656 B.n910 B.n104 256.663
R657 B.n910 B.n103 256.663
R658 B.n910 B.n102 256.663
R659 B.n910 B.n101 256.663
R660 B.n910 B.n100 256.663
R661 B.n910 B.n99 256.663
R662 B.n910 B.n98 256.663
R663 B.n910 B.n97 256.663
R664 B.n910 B.n96 256.663
R665 B.n910 B.n95 256.663
R666 B.n910 B.n94 256.663
R667 B.n910 B.n93 256.663
R668 B.n910 B.n92 256.663
R669 B.n910 B.n91 256.663
R670 B.n910 B.n90 256.663
R671 B.n910 B.n89 256.663
R672 B.n910 B.n88 256.663
R673 B.n910 B.n87 256.663
R674 B.n910 B.n86 256.663
R675 B.n910 B.n85 256.663
R676 B.n910 B.n84 256.663
R677 B.n910 B.n83 256.663
R678 B.n910 B.n82 256.663
R679 B.n910 B.n81 256.663
R680 B.n910 B.n80 256.663
R681 B.n910 B.n79 256.663
R682 B.n910 B.n78 256.663
R683 B.n910 B.n77 256.663
R684 B.n910 B.n76 256.663
R685 B.n910 B.n75 256.663
R686 B.n910 B.n74 256.663
R687 B.n910 B.n73 256.663
R688 B.n910 B.n72 256.663
R689 B.n910 B.n71 256.663
R690 B.n910 B.n70 256.663
R691 B.n910 B.n69 256.663
R692 B.n911 B.n910 256.663
R693 B.n754 B.n753 256.663
R694 B.n753 B.n445 256.663
R695 B.n753 B.n446 256.663
R696 B.n753 B.n447 256.663
R697 B.n753 B.n448 256.663
R698 B.n753 B.n449 256.663
R699 B.n753 B.n450 256.663
R700 B.n753 B.n451 256.663
R701 B.n753 B.n452 256.663
R702 B.n753 B.n453 256.663
R703 B.n753 B.n454 256.663
R704 B.n753 B.n455 256.663
R705 B.n753 B.n456 256.663
R706 B.n753 B.n457 256.663
R707 B.n753 B.n458 256.663
R708 B.n753 B.n459 256.663
R709 B.n753 B.n460 256.663
R710 B.n753 B.n461 256.663
R711 B.n753 B.n462 256.663
R712 B.n753 B.n463 256.663
R713 B.n753 B.n464 256.663
R714 B.n753 B.n465 256.663
R715 B.n753 B.n466 256.663
R716 B.n753 B.n467 256.663
R717 B.n753 B.n468 256.663
R718 B.n753 B.n469 256.663
R719 B.n753 B.n470 256.663
R720 B.n753 B.n471 256.663
R721 B.n753 B.n472 256.663
R722 B.n753 B.n473 256.663
R723 B.n753 B.n474 256.663
R724 B.n753 B.n475 256.663
R725 B.n753 B.n476 256.663
R726 B.n753 B.n477 256.663
R727 B.n753 B.n478 256.663
R728 B.n753 B.n479 256.663
R729 B.n753 B.n480 256.663
R730 B.n753 B.n481 256.663
R731 B.n753 B.n482 256.663
R732 B.n753 B.n483 256.663
R733 B.n753 B.n484 256.663
R734 B.n753 B.n485 256.663
R735 B.n753 B.n486 256.663
R736 B.n753 B.n487 256.663
R737 B.n753 B.n488 256.663
R738 B.n753 B.n489 256.663
R739 B.n753 B.n490 256.663
R740 B.n753 B.n491 256.663
R741 B.n753 B.n492 256.663
R742 B.n753 B.n493 256.663
R743 B.n753 B.n494 256.663
R744 B.n753 B.n495 256.663
R745 B.n753 B.n496 256.663
R746 B.n753 B.n497 256.663
R747 B.n753 B.n498 256.663
R748 B.n753 B.n499 256.663
R749 B.n753 B.n500 256.663
R750 B.n753 B.n501 256.663
R751 B.n753 B.n502 256.663
R752 B.n753 B.n503 256.663
R753 B.n753 B.n504 256.663
R754 B.n987 B.n986 256.663
R755 B.n136 B.n68 163.367
R756 B.n140 B.n139 163.367
R757 B.n144 B.n143 163.367
R758 B.n148 B.n147 163.367
R759 B.n152 B.n151 163.367
R760 B.n156 B.n155 163.367
R761 B.n160 B.n159 163.367
R762 B.n164 B.n163 163.367
R763 B.n168 B.n167 163.367
R764 B.n172 B.n171 163.367
R765 B.n176 B.n175 163.367
R766 B.n180 B.n179 163.367
R767 B.n184 B.n183 163.367
R768 B.n188 B.n187 163.367
R769 B.n192 B.n191 163.367
R770 B.n196 B.n195 163.367
R771 B.n200 B.n199 163.367
R772 B.n204 B.n203 163.367
R773 B.n208 B.n207 163.367
R774 B.n212 B.n211 163.367
R775 B.n216 B.n215 163.367
R776 B.n220 B.n219 163.367
R777 B.n224 B.n223 163.367
R778 B.n228 B.n227 163.367
R779 B.n232 B.n231 163.367
R780 B.n236 B.n235 163.367
R781 B.n240 B.n239 163.367
R782 B.n244 B.n243 163.367
R783 B.n249 B.n248 163.367
R784 B.n253 B.n252 163.367
R785 B.n257 B.n256 163.367
R786 B.n261 B.n260 163.367
R787 B.n265 B.n264 163.367
R788 B.n269 B.n268 163.367
R789 B.n273 B.n272 163.367
R790 B.n277 B.n276 163.367
R791 B.n281 B.n280 163.367
R792 B.n285 B.n284 163.367
R793 B.n289 B.n288 163.367
R794 B.n293 B.n292 163.367
R795 B.n297 B.n296 163.367
R796 B.n301 B.n300 163.367
R797 B.n305 B.n304 163.367
R798 B.n309 B.n308 163.367
R799 B.n313 B.n312 163.367
R800 B.n317 B.n316 163.367
R801 B.n321 B.n320 163.367
R802 B.n325 B.n324 163.367
R803 B.n329 B.n328 163.367
R804 B.n333 B.n332 163.367
R805 B.n337 B.n336 163.367
R806 B.n341 B.n340 163.367
R807 B.n345 B.n344 163.367
R808 B.n349 B.n348 163.367
R809 B.n353 B.n352 163.367
R810 B.n357 B.n356 163.367
R811 B.n361 B.n360 163.367
R812 B.n365 B.n364 163.367
R813 B.n369 B.n368 163.367
R814 B.n373 B.n372 163.367
R815 B.n909 B.n129 163.367
R816 B.n761 B.n440 163.367
R817 B.n761 B.n438 163.367
R818 B.n765 B.n438 163.367
R819 B.n765 B.n431 163.367
R820 B.n773 B.n431 163.367
R821 B.n773 B.n429 163.367
R822 B.n777 B.n429 163.367
R823 B.n777 B.n424 163.367
R824 B.n785 B.n424 163.367
R825 B.n785 B.n422 163.367
R826 B.n789 B.n422 163.367
R827 B.n789 B.n416 163.367
R828 B.n797 B.n416 163.367
R829 B.n797 B.n414 163.367
R830 B.n801 B.n414 163.367
R831 B.n801 B.n409 163.367
R832 B.n810 B.n409 163.367
R833 B.n810 B.n407 163.367
R834 B.n814 B.n407 163.367
R835 B.n814 B.n401 163.367
R836 B.n822 B.n401 163.367
R837 B.n822 B.n399 163.367
R838 B.n826 B.n399 163.367
R839 B.n826 B.n393 163.367
R840 B.n834 B.n393 163.367
R841 B.n834 B.n391 163.367
R842 B.n838 B.n391 163.367
R843 B.n838 B.n384 163.367
R844 B.n846 B.n384 163.367
R845 B.n846 B.n382 163.367
R846 B.n851 B.n382 163.367
R847 B.n851 B.n377 163.367
R848 B.n859 B.n377 163.367
R849 B.n860 B.n859 163.367
R850 B.n860 B.n5 163.367
R851 B.n6 B.n5 163.367
R852 B.n7 B.n6 163.367
R853 B.n866 B.n7 163.367
R854 B.n867 B.n866 163.367
R855 B.n867 B.n13 163.367
R856 B.n14 B.n13 163.367
R857 B.n15 B.n14 163.367
R858 B.n872 B.n15 163.367
R859 B.n872 B.n20 163.367
R860 B.n21 B.n20 163.367
R861 B.n22 B.n21 163.367
R862 B.n877 B.n22 163.367
R863 B.n877 B.n27 163.367
R864 B.n28 B.n27 163.367
R865 B.n29 B.n28 163.367
R866 B.n882 B.n29 163.367
R867 B.n882 B.n34 163.367
R868 B.n35 B.n34 163.367
R869 B.n36 B.n35 163.367
R870 B.n887 B.n36 163.367
R871 B.n887 B.n41 163.367
R872 B.n42 B.n41 163.367
R873 B.n43 B.n42 163.367
R874 B.n892 B.n43 163.367
R875 B.n892 B.n48 163.367
R876 B.n49 B.n48 163.367
R877 B.n50 B.n49 163.367
R878 B.n897 B.n50 163.367
R879 B.n897 B.n55 163.367
R880 B.n56 B.n55 163.367
R881 B.n57 B.n56 163.367
R882 B.n902 B.n57 163.367
R883 B.n902 B.n62 163.367
R884 B.n63 B.n62 163.367
R885 B.n64 B.n63 163.367
R886 B.n130 B.n64 163.367
R887 B.n752 B.n444 163.367
R888 B.n752 B.n505 163.367
R889 B.n748 B.n747 163.367
R890 B.n744 B.n743 163.367
R891 B.n740 B.n739 163.367
R892 B.n736 B.n735 163.367
R893 B.n732 B.n731 163.367
R894 B.n728 B.n727 163.367
R895 B.n724 B.n723 163.367
R896 B.n720 B.n719 163.367
R897 B.n716 B.n715 163.367
R898 B.n712 B.n711 163.367
R899 B.n708 B.n707 163.367
R900 B.n704 B.n703 163.367
R901 B.n700 B.n699 163.367
R902 B.n696 B.n695 163.367
R903 B.n692 B.n691 163.367
R904 B.n688 B.n687 163.367
R905 B.n684 B.n683 163.367
R906 B.n680 B.n679 163.367
R907 B.n676 B.n675 163.367
R908 B.n672 B.n671 163.367
R909 B.n668 B.n667 163.367
R910 B.n664 B.n663 163.367
R911 B.n660 B.n659 163.367
R912 B.n656 B.n655 163.367
R913 B.n652 B.n651 163.367
R914 B.n648 B.n647 163.367
R915 B.n644 B.n643 163.367
R916 B.n640 B.n639 163.367
R917 B.n636 B.n635 163.367
R918 B.n632 B.n631 163.367
R919 B.n628 B.n627 163.367
R920 B.n623 B.n622 163.367
R921 B.n619 B.n618 163.367
R922 B.n615 B.n614 163.367
R923 B.n611 B.n610 163.367
R924 B.n607 B.n606 163.367
R925 B.n603 B.n602 163.367
R926 B.n599 B.n598 163.367
R927 B.n595 B.n594 163.367
R928 B.n591 B.n590 163.367
R929 B.n587 B.n586 163.367
R930 B.n583 B.n582 163.367
R931 B.n579 B.n578 163.367
R932 B.n575 B.n574 163.367
R933 B.n571 B.n570 163.367
R934 B.n567 B.n566 163.367
R935 B.n563 B.n562 163.367
R936 B.n559 B.n558 163.367
R937 B.n555 B.n554 163.367
R938 B.n551 B.n550 163.367
R939 B.n547 B.n546 163.367
R940 B.n543 B.n542 163.367
R941 B.n539 B.n538 163.367
R942 B.n535 B.n534 163.367
R943 B.n531 B.n530 163.367
R944 B.n527 B.n526 163.367
R945 B.n523 B.n522 163.367
R946 B.n519 B.n518 163.367
R947 B.n515 B.n514 163.367
R948 B.n759 B.n442 163.367
R949 B.n759 B.n436 163.367
R950 B.n767 B.n436 163.367
R951 B.n767 B.n434 163.367
R952 B.n771 B.n434 163.367
R953 B.n771 B.n428 163.367
R954 B.n779 B.n428 163.367
R955 B.n779 B.n426 163.367
R956 B.n783 B.n426 163.367
R957 B.n783 B.n420 163.367
R958 B.n791 B.n420 163.367
R959 B.n791 B.n418 163.367
R960 B.n795 B.n418 163.367
R961 B.n795 B.n412 163.367
R962 B.n804 B.n412 163.367
R963 B.n804 B.n410 163.367
R964 B.n808 B.n410 163.367
R965 B.n808 B.n405 163.367
R966 B.n816 B.n405 163.367
R967 B.n816 B.n403 163.367
R968 B.n820 B.n403 163.367
R969 B.n820 B.n397 163.367
R970 B.n828 B.n397 163.367
R971 B.n828 B.n395 163.367
R972 B.n832 B.n395 163.367
R973 B.n832 B.n389 163.367
R974 B.n840 B.n389 163.367
R975 B.n840 B.n387 163.367
R976 B.n844 B.n387 163.367
R977 B.n844 B.n381 163.367
R978 B.n853 B.n381 163.367
R979 B.n853 B.n379 163.367
R980 B.n857 B.n379 163.367
R981 B.n857 B.n3 163.367
R982 B.n985 B.n3 163.367
R983 B.n981 B.n2 163.367
R984 B.n981 B.n980 163.367
R985 B.n980 B.n9 163.367
R986 B.n976 B.n9 163.367
R987 B.n976 B.n11 163.367
R988 B.n972 B.n11 163.367
R989 B.n972 B.n17 163.367
R990 B.n968 B.n17 163.367
R991 B.n968 B.n19 163.367
R992 B.n964 B.n19 163.367
R993 B.n964 B.n24 163.367
R994 B.n960 B.n24 163.367
R995 B.n960 B.n26 163.367
R996 B.n956 B.n26 163.367
R997 B.n956 B.n31 163.367
R998 B.n952 B.n31 163.367
R999 B.n952 B.n33 163.367
R1000 B.n948 B.n33 163.367
R1001 B.n948 B.n37 163.367
R1002 B.n944 B.n37 163.367
R1003 B.n944 B.n39 163.367
R1004 B.n940 B.n39 163.367
R1005 B.n940 B.n45 163.367
R1006 B.n936 B.n45 163.367
R1007 B.n936 B.n47 163.367
R1008 B.n932 B.n47 163.367
R1009 B.n932 B.n52 163.367
R1010 B.n928 B.n52 163.367
R1011 B.n928 B.n54 163.367
R1012 B.n924 B.n54 163.367
R1013 B.n924 B.n59 163.367
R1014 B.n920 B.n59 163.367
R1015 B.n920 B.n61 163.367
R1016 B.n916 B.n61 163.367
R1017 B.n916 B.n66 163.367
R1018 B.n131 B.t18 114.819
R1019 B.n509 B.t16 114.819
R1020 B.n134 B.t12 114.796
R1021 B.n506 B.t9 114.796
R1022 B.n912 B.n911 71.676
R1023 B.n136 B.n69 71.676
R1024 B.n140 B.n70 71.676
R1025 B.n144 B.n71 71.676
R1026 B.n148 B.n72 71.676
R1027 B.n152 B.n73 71.676
R1028 B.n156 B.n74 71.676
R1029 B.n160 B.n75 71.676
R1030 B.n164 B.n76 71.676
R1031 B.n168 B.n77 71.676
R1032 B.n172 B.n78 71.676
R1033 B.n176 B.n79 71.676
R1034 B.n180 B.n80 71.676
R1035 B.n184 B.n81 71.676
R1036 B.n188 B.n82 71.676
R1037 B.n192 B.n83 71.676
R1038 B.n196 B.n84 71.676
R1039 B.n200 B.n85 71.676
R1040 B.n204 B.n86 71.676
R1041 B.n208 B.n87 71.676
R1042 B.n212 B.n88 71.676
R1043 B.n216 B.n89 71.676
R1044 B.n220 B.n90 71.676
R1045 B.n224 B.n91 71.676
R1046 B.n228 B.n92 71.676
R1047 B.n232 B.n93 71.676
R1048 B.n236 B.n94 71.676
R1049 B.n240 B.n95 71.676
R1050 B.n244 B.n96 71.676
R1051 B.n249 B.n97 71.676
R1052 B.n253 B.n98 71.676
R1053 B.n257 B.n99 71.676
R1054 B.n261 B.n100 71.676
R1055 B.n265 B.n101 71.676
R1056 B.n269 B.n102 71.676
R1057 B.n273 B.n103 71.676
R1058 B.n277 B.n104 71.676
R1059 B.n281 B.n105 71.676
R1060 B.n285 B.n106 71.676
R1061 B.n289 B.n107 71.676
R1062 B.n293 B.n108 71.676
R1063 B.n297 B.n109 71.676
R1064 B.n301 B.n110 71.676
R1065 B.n305 B.n111 71.676
R1066 B.n309 B.n112 71.676
R1067 B.n313 B.n113 71.676
R1068 B.n317 B.n114 71.676
R1069 B.n321 B.n115 71.676
R1070 B.n325 B.n116 71.676
R1071 B.n329 B.n117 71.676
R1072 B.n333 B.n118 71.676
R1073 B.n337 B.n119 71.676
R1074 B.n341 B.n120 71.676
R1075 B.n345 B.n121 71.676
R1076 B.n349 B.n122 71.676
R1077 B.n353 B.n123 71.676
R1078 B.n357 B.n124 71.676
R1079 B.n361 B.n125 71.676
R1080 B.n365 B.n126 71.676
R1081 B.n369 B.n127 71.676
R1082 B.n373 B.n128 71.676
R1083 B.n129 B.n128 71.676
R1084 B.n372 B.n127 71.676
R1085 B.n368 B.n126 71.676
R1086 B.n364 B.n125 71.676
R1087 B.n360 B.n124 71.676
R1088 B.n356 B.n123 71.676
R1089 B.n352 B.n122 71.676
R1090 B.n348 B.n121 71.676
R1091 B.n344 B.n120 71.676
R1092 B.n340 B.n119 71.676
R1093 B.n336 B.n118 71.676
R1094 B.n332 B.n117 71.676
R1095 B.n328 B.n116 71.676
R1096 B.n324 B.n115 71.676
R1097 B.n320 B.n114 71.676
R1098 B.n316 B.n113 71.676
R1099 B.n312 B.n112 71.676
R1100 B.n308 B.n111 71.676
R1101 B.n304 B.n110 71.676
R1102 B.n300 B.n109 71.676
R1103 B.n296 B.n108 71.676
R1104 B.n292 B.n107 71.676
R1105 B.n288 B.n106 71.676
R1106 B.n284 B.n105 71.676
R1107 B.n280 B.n104 71.676
R1108 B.n276 B.n103 71.676
R1109 B.n272 B.n102 71.676
R1110 B.n268 B.n101 71.676
R1111 B.n264 B.n100 71.676
R1112 B.n260 B.n99 71.676
R1113 B.n256 B.n98 71.676
R1114 B.n252 B.n97 71.676
R1115 B.n248 B.n96 71.676
R1116 B.n243 B.n95 71.676
R1117 B.n239 B.n94 71.676
R1118 B.n235 B.n93 71.676
R1119 B.n231 B.n92 71.676
R1120 B.n227 B.n91 71.676
R1121 B.n223 B.n90 71.676
R1122 B.n219 B.n89 71.676
R1123 B.n215 B.n88 71.676
R1124 B.n211 B.n87 71.676
R1125 B.n207 B.n86 71.676
R1126 B.n203 B.n85 71.676
R1127 B.n199 B.n84 71.676
R1128 B.n195 B.n83 71.676
R1129 B.n191 B.n82 71.676
R1130 B.n187 B.n81 71.676
R1131 B.n183 B.n80 71.676
R1132 B.n179 B.n79 71.676
R1133 B.n175 B.n78 71.676
R1134 B.n171 B.n77 71.676
R1135 B.n167 B.n76 71.676
R1136 B.n163 B.n75 71.676
R1137 B.n159 B.n74 71.676
R1138 B.n155 B.n73 71.676
R1139 B.n151 B.n72 71.676
R1140 B.n147 B.n71 71.676
R1141 B.n143 B.n70 71.676
R1142 B.n139 B.n69 71.676
R1143 B.n911 B.n68 71.676
R1144 B.n755 B.n754 71.676
R1145 B.n505 B.n445 71.676
R1146 B.n747 B.n446 71.676
R1147 B.n743 B.n447 71.676
R1148 B.n739 B.n448 71.676
R1149 B.n735 B.n449 71.676
R1150 B.n731 B.n450 71.676
R1151 B.n727 B.n451 71.676
R1152 B.n723 B.n452 71.676
R1153 B.n719 B.n453 71.676
R1154 B.n715 B.n454 71.676
R1155 B.n711 B.n455 71.676
R1156 B.n707 B.n456 71.676
R1157 B.n703 B.n457 71.676
R1158 B.n699 B.n458 71.676
R1159 B.n695 B.n459 71.676
R1160 B.n691 B.n460 71.676
R1161 B.n687 B.n461 71.676
R1162 B.n683 B.n462 71.676
R1163 B.n679 B.n463 71.676
R1164 B.n675 B.n464 71.676
R1165 B.n671 B.n465 71.676
R1166 B.n667 B.n466 71.676
R1167 B.n663 B.n467 71.676
R1168 B.n659 B.n468 71.676
R1169 B.n655 B.n469 71.676
R1170 B.n651 B.n470 71.676
R1171 B.n647 B.n471 71.676
R1172 B.n643 B.n472 71.676
R1173 B.n639 B.n473 71.676
R1174 B.n635 B.n474 71.676
R1175 B.n631 B.n475 71.676
R1176 B.n627 B.n476 71.676
R1177 B.n622 B.n477 71.676
R1178 B.n618 B.n478 71.676
R1179 B.n614 B.n479 71.676
R1180 B.n610 B.n480 71.676
R1181 B.n606 B.n481 71.676
R1182 B.n602 B.n482 71.676
R1183 B.n598 B.n483 71.676
R1184 B.n594 B.n484 71.676
R1185 B.n590 B.n485 71.676
R1186 B.n586 B.n486 71.676
R1187 B.n582 B.n487 71.676
R1188 B.n578 B.n488 71.676
R1189 B.n574 B.n489 71.676
R1190 B.n570 B.n490 71.676
R1191 B.n566 B.n491 71.676
R1192 B.n562 B.n492 71.676
R1193 B.n558 B.n493 71.676
R1194 B.n554 B.n494 71.676
R1195 B.n550 B.n495 71.676
R1196 B.n546 B.n496 71.676
R1197 B.n542 B.n497 71.676
R1198 B.n538 B.n498 71.676
R1199 B.n534 B.n499 71.676
R1200 B.n530 B.n500 71.676
R1201 B.n526 B.n501 71.676
R1202 B.n522 B.n502 71.676
R1203 B.n518 B.n503 71.676
R1204 B.n514 B.n504 71.676
R1205 B.n754 B.n444 71.676
R1206 B.n748 B.n445 71.676
R1207 B.n744 B.n446 71.676
R1208 B.n740 B.n447 71.676
R1209 B.n736 B.n448 71.676
R1210 B.n732 B.n449 71.676
R1211 B.n728 B.n450 71.676
R1212 B.n724 B.n451 71.676
R1213 B.n720 B.n452 71.676
R1214 B.n716 B.n453 71.676
R1215 B.n712 B.n454 71.676
R1216 B.n708 B.n455 71.676
R1217 B.n704 B.n456 71.676
R1218 B.n700 B.n457 71.676
R1219 B.n696 B.n458 71.676
R1220 B.n692 B.n459 71.676
R1221 B.n688 B.n460 71.676
R1222 B.n684 B.n461 71.676
R1223 B.n680 B.n462 71.676
R1224 B.n676 B.n463 71.676
R1225 B.n672 B.n464 71.676
R1226 B.n668 B.n465 71.676
R1227 B.n664 B.n466 71.676
R1228 B.n660 B.n467 71.676
R1229 B.n656 B.n468 71.676
R1230 B.n652 B.n469 71.676
R1231 B.n648 B.n470 71.676
R1232 B.n644 B.n471 71.676
R1233 B.n640 B.n472 71.676
R1234 B.n636 B.n473 71.676
R1235 B.n632 B.n474 71.676
R1236 B.n628 B.n475 71.676
R1237 B.n623 B.n476 71.676
R1238 B.n619 B.n477 71.676
R1239 B.n615 B.n478 71.676
R1240 B.n611 B.n479 71.676
R1241 B.n607 B.n480 71.676
R1242 B.n603 B.n481 71.676
R1243 B.n599 B.n482 71.676
R1244 B.n595 B.n483 71.676
R1245 B.n591 B.n484 71.676
R1246 B.n587 B.n485 71.676
R1247 B.n583 B.n486 71.676
R1248 B.n579 B.n487 71.676
R1249 B.n575 B.n488 71.676
R1250 B.n571 B.n489 71.676
R1251 B.n567 B.n490 71.676
R1252 B.n563 B.n491 71.676
R1253 B.n559 B.n492 71.676
R1254 B.n555 B.n493 71.676
R1255 B.n551 B.n494 71.676
R1256 B.n547 B.n495 71.676
R1257 B.n543 B.n496 71.676
R1258 B.n539 B.n497 71.676
R1259 B.n535 B.n498 71.676
R1260 B.n531 B.n499 71.676
R1261 B.n527 B.n500 71.676
R1262 B.n523 B.n501 71.676
R1263 B.n519 B.n502 71.676
R1264 B.n515 B.n503 71.676
R1265 B.n511 B.n504 71.676
R1266 B.n986 B.n985 71.676
R1267 B.n986 B.n2 71.676
R1268 B.n132 B.t19 69.8245
R1269 B.n510 B.t15 69.8245
R1270 B.n135 B.t13 69.8017
R1271 B.n507 B.t8 69.8017
R1272 B.n246 B.n135 59.5399
R1273 B.n133 B.n132 59.5399
R1274 B.n625 B.n510 59.5399
R1275 B.n508 B.n507 59.5399
R1276 B.n753 B.n441 57.443
R1277 B.n910 B.n65 57.443
R1278 B.n135 B.n134 44.9944
R1279 B.n132 B.n131 44.9944
R1280 B.n510 B.n509 44.9944
R1281 B.n507 B.n506 44.9944
R1282 B.n760 B.n441 33.3859
R1283 B.n760 B.n437 33.3859
R1284 B.n766 B.n437 33.3859
R1285 B.n766 B.n432 33.3859
R1286 B.n772 B.n432 33.3859
R1287 B.n772 B.n433 33.3859
R1288 B.n778 B.n425 33.3859
R1289 B.n784 B.n425 33.3859
R1290 B.n784 B.n421 33.3859
R1291 B.n790 B.n421 33.3859
R1292 B.n790 B.n417 33.3859
R1293 B.n796 B.n417 33.3859
R1294 B.n796 B.n413 33.3859
R1295 B.n803 B.n413 33.3859
R1296 B.n803 B.n802 33.3859
R1297 B.n809 B.n406 33.3859
R1298 B.n815 B.n406 33.3859
R1299 B.n815 B.n402 33.3859
R1300 B.n821 B.n402 33.3859
R1301 B.n821 B.n398 33.3859
R1302 B.n827 B.n398 33.3859
R1303 B.n833 B.n394 33.3859
R1304 B.n833 B.n390 33.3859
R1305 B.n839 B.n390 33.3859
R1306 B.n839 B.n385 33.3859
R1307 B.n845 B.n385 33.3859
R1308 B.n845 B.n386 33.3859
R1309 B.n852 B.n378 33.3859
R1310 B.n858 B.n378 33.3859
R1311 B.n858 B.n4 33.3859
R1312 B.n984 B.n4 33.3859
R1313 B.n984 B.n983 33.3859
R1314 B.n983 B.n982 33.3859
R1315 B.n982 B.n8 33.3859
R1316 B.n12 B.n8 33.3859
R1317 B.n975 B.n12 33.3859
R1318 B.n974 B.n973 33.3859
R1319 B.n973 B.n16 33.3859
R1320 B.n967 B.n16 33.3859
R1321 B.n967 B.n966 33.3859
R1322 B.n966 B.n965 33.3859
R1323 B.n965 B.n23 33.3859
R1324 B.n959 B.n958 33.3859
R1325 B.n958 B.n957 33.3859
R1326 B.n957 B.n30 33.3859
R1327 B.n951 B.n30 33.3859
R1328 B.n951 B.n950 33.3859
R1329 B.n950 B.n949 33.3859
R1330 B.n943 B.n40 33.3859
R1331 B.n943 B.n942 33.3859
R1332 B.n942 B.n941 33.3859
R1333 B.n941 B.n44 33.3859
R1334 B.n935 B.n44 33.3859
R1335 B.n935 B.n934 33.3859
R1336 B.n934 B.n933 33.3859
R1337 B.n933 B.n51 33.3859
R1338 B.n927 B.n51 33.3859
R1339 B.n926 B.n925 33.3859
R1340 B.n925 B.n58 33.3859
R1341 B.n919 B.n58 33.3859
R1342 B.n919 B.n918 33.3859
R1343 B.n918 B.n917 33.3859
R1344 B.n917 B.n65 33.3859
R1345 B.n757 B.n756 31.3761
R1346 B.n512 B.n439 31.3761
R1347 B.n908 B.n907 31.3761
R1348 B.n914 B.n913 31.3761
R1349 B.n802 B.t4 27.9853
R1350 B.n40 B.t2 27.9853
R1351 B.n433 B.t7 27.0034
R1352 B.t11 B.n926 27.0034
R1353 B.n827 B.t5 22.0938
R1354 B.n959 B.t0 22.0938
R1355 B B.n987 18.0485
R1356 B.n852 B.t3 17.1842
R1357 B.n975 B.t1 17.1842
R1358 B.n386 B.t3 16.2022
R1359 B.t1 B.n974 16.2022
R1360 B.t5 B.n394 11.2926
R1361 B.t0 B.n23 11.2926
R1362 B.n758 B.n757 10.6151
R1363 B.n758 B.n435 10.6151
R1364 B.n768 B.n435 10.6151
R1365 B.n769 B.n768 10.6151
R1366 B.n770 B.n769 10.6151
R1367 B.n770 B.n427 10.6151
R1368 B.n780 B.n427 10.6151
R1369 B.n781 B.n780 10.6151
R1370 B.n782 B.n781 10.6151
R1371 B.n782 B.n419 10.6151
R1372 B.n792 B.n419 10.6151
R1373 B.n793 B.n792 10.6151
R1374 B.n794 B.n793 10.6151
R1375 B.n794 B.n411 10.6151
R1376 B.n805 B.n411 10.6151
R1377 B.n806 B.n805 10.6151
R1378 B.n807 B.n806 10.6151
R1379 B.n807 B.n404 10.6151
R1380 B.n817 B.n404 10.6151
R1381 B.n818 B.n817 10.6151
R1382 B.n819 B.n818 10.6151
R1383 B.n819 B.n396 10.6151
R1384 B.n829 B.n396 10.6151
R1385 B.n830 B.n829 10.6151
R1386 B.n831 B.n830 10.6151
R1387 B.n831 B.n388 10.6151
R1388 B.n841 B.n388 10.6151
R1389 B.n842 B.n841 10.6151
R1390 B.n843 B.n842 10.6151
R1391 B.n843 B.n380 10.6151
R1392 B.n854 B.n380 10.6151
R1393 B.n855 B.n854 10.6151
R1394 B.n856 B.n855 10.6151
R1395 B.n856 B.n0 10.6151
R1396 B.n756 B.n443 10.6151
R1397 B.n751 B.n443 10.6151
R1398 B.n751 B.n750 10.6151
R1399 B.n750 B.n749 10.6151
R1400 B.n749 B.n746 10.6151
R1401 B.n746 B.n745 10.6151
R1402 B.n745 B.n742 10.6151
R1403 B.n742 B.n741 10.6151
R1404 B.n741 B.n738 10.6151
R1405 B.n738 B.n737 10.6151
R1406 B.n737 B.n734 10.6151
R1407 B.n734 B.n733 10.6151
R1408 B.n733 B.n730 10.6151
R1409 B.n730 B.n729 10.6151
R1410 B.n729 B.n726 10.6151
R1411 B.n726 B.n725 10.6151
R1412 B.n725 B.n722 10.6151
R1413 B.n722 B.n721 10.6151
R1414 B.n721 B.n718 10.6151
R1415 B.n718 B.n717 10.6151
R1416 B.n717 B.n714 10.6151
R1417 B.n714 B.n713 10.6151
R1418 B.n713 B.n710 10.6151
R1419 B.n710 B.n709 10.6151
R1420 B.n709 B.n706 10.6151
R1421 B.n706 B.n705 10.6151
R1422 B.n705 B.n702 10.6151
R1423 B.n702 B.n701 10.6151
R1424 B.n701 B.n698 10.6151
R1425 B.n698 B.n697 10.6151
R1426 B.n697 B.n694 10.6151
R1427 B.n694 B.n693 10.6151
R1428 B.n693 B.n690 10.6151
R1429 B.n690 B.n689 10.6151
R1430 B.n689 B.n686 10.6151
R1431 B.n686 B.n685 10.6151
R1432 B.n685 B.n682 10.6151
R1433 B.n682 B.n681 10.6151
R1434 B.n681 B.n678 10.6151
R1435 B.n678 B.n677 10.6151
R1436 B.n677 B.n674 10.6151
R1437 B.n674 B.n673 10.6151
R1438 B.n673 B.n670 10.6151
R1439 B.n670 B.n669 10.6151
R1440 B.n669 B.n666 10.6151
R1441 B.n666 B.n665 10.6151
R1442 B.n665 B.n662 10.6151
R1443 B.n662 B.n661 10.6151
R1444 B.n661 B.n658 10.6151
R1445 B.n658 B.n657 10.6151
R1446 B.n657 B.n654 10.6151
R1447 B.n654 B.n653 10.6151
R1448 B.n653 B.n650 10.6151
R1449 B.n650 B.n649 10.6151
R1450 B.n649 B.n646 10.6151
R1451 B.n646 B.n645 10.6151
R1452 B.n642 B.n641 10.6151
R1453 B.n641 B.n638 10.6151
R1454 B.n638 B.n637 10.6151
R1455 B.n637 B.n634 10.6151
R1456 B.n634 B.n633 10.6151
R1457 B.n633 B.n630 10.6151
R1458 B.n630 B.n629 10.6151
R1459 B.n629 B.n626 10.6151
R1460 B.n624 B.n621 10.6151
R1461 B.n621 B.n620 10.6151
R1462 B.n620 B.n617 10.6151
R1463 B.n617 B.n616 10.6151
R1464 B.n616 B.n613 10.6151
R1465 B.n613 B.n612 10.6151
R1466 B.n612 B.n609 10.6151
R1467 B.n609 B.n608 10.6151
R1468 B.n608 B.n605 10.6151
R1469 B.n605 B.n604 10.6151
R1470 B.n604 B.n601 10.6151
R1471 B.n601 B.n600 10.6151
R1472 B.n600 B.n597 10.6151
R1473 B.n597 B.n596 10.6151
R1474 B.n596 B.n593 10.6151
R1475 B.n593 B.n592 10.6151
R1476 B.n592 B.n589 10.6151
R1477 B.n589 B.n588 10.6151
R1478 B.n588 B.n585 10.6151
R1479 B.n585 B.n584 10.6151
R1480 B.n584 B.n581 10.6151
R1481 B.n581 B.n580 10.6151
R1482 B.n580 B.n577 10.6151
R1483 B.n577 B.n576 10.6151
R1484 B.n576 B.n573 10.6151
R1485 B.n573 B.n572 10.6151
R1486 B.n572 B.n569 10.6151
R1487 B.n569 B.n568 10.6151
R1488 B.n568 B.n565 10.6151
R1489 B.n565 B.n564 10.6151
R1490 B.n564 B.n561 10.6151
R1491 B.n561 B.n560 10.6151
R1492 B.n560 B.n557 10.6151
R1493 B.n557 B.n556 10.6151
R1494 B.n556 B.n553 10.6151
R1495 B.n553 B.n552 10.6151
R1496 B.n552 B.n549 10.6151
R1497 B.n549 B.n548 10.6151
R1498 B.n548 B.n545 10.6151
R1499 B.n545 B.n544 10.6151
R1500 B.n544 B.n541 10.6151
R1501 B.n541 B.n540 10.6151
R1502 B.n540 B.n537 10.6151
R1503 B.n537 B.n536 10.6151
R1504 B.n536 B.n533 10.6151
R1505 B.n533 B.n532 10.6151
R1506 B.n532 B.n529 10.6151
R1507 B.n529 B.n528 10.6151
R1508 B.n528 B.n525 10.6151
R1509 B.n525 B.n524 10.6151
R1510 B.n524 B.n521 10.6151
R1511 B.n521 B.n520 10.6151
R1512 B.n520 B.n517 10.6151
R1513 B.n517 B.n516 10.6151
R1514 B.n516 B.n513 10.6151
R1515 B.n513 B.n512 10.6151
R1516 B.n762 B.n439 10.6151
R1517 B.n763 B.n762 10.6151
R1518 B.n764 B.n763 10.6151
R1519 B.n764 B.n430 10.6151
R1520 B.n774 B.n430 10.6151
R1521 B.n775 B.n774 10.6151
R1522 B.n776 B.n775 10.6151
R1523 B.n776 B.n423 10.6151
R1524 B.n786 B.n423 10.6151
R1525 B.n787 B.n786 10.6151
R1526 B.n788 B.n787 10.6151
R1527 B.n788 B.n415 10.6151
R1528 B.n798 B.n415 10.6151
R1529 B.n799 B.n798 10.6151
R1530 B.n800 B.n799 10.6151
R1531 B.n800 B.n408 10.6151
R1532 B.n811 B.n408 10.6151
R1533 B.n812 B.n811 10.6151
R1534 B.n813 B.n812 10.6151
R1535 B.n813 B.n400 10.6151
R1536 B.n823 B.n400 10.6151
R1537 B.n824 B.n823 10.6151
R1538 B.n825 B.n824 10.6151
R1539 B.n825 B.n392 10.6151
R1540 B.n835 B.n392 10.6151
R1541 B.n836 B.n835 10.6151
R1542 B.n837 B.n836 10.6151
R1543 B.n837 B.n383 10.6151
R1544 B.n847 B.n383 10.6151
R1545 B.n848 B.n847 10.6151
R1546 B.n850 B.n848 10.6151
R1547 B.n850 B.n849 10.6151
R1548 B.n849 B.n376 10.6151
R1549 B.n861 B.n376 10.6151
R1550 B.n862 B.n861 10.6151
R1551 B.n863 B.n862 10.6151
R1552 B.n864 B.n863 10.6151
R1553 B.n865 B.n864 10.6151
R1554 B.n868 B.n865 10.6151
R1555 B.n869 B.n868 10.6151
R1556 B.n870 B.n869 10.6151
R1557 B.n871 B.n870 10.6151
R1558 B.n873 B.n871 10.6151
R1559 B.n874 B.n873 10.6151
R1560 B.n875 B.n874 10.6151
R1561 B.n876 B.n875 10.6151
R1562 B.n878 B.n876 10.6151
R1563 B.n879 B.n878 10.6151
R1564 B.n880 B.n879 10.6151
R1565 B.n881 B.n880 10.6151
R1566 B.n883 B.n881 10.6151
R1567 B.n884 B.n883 10.6151
R1568 B.n885 B.n884 10.6151
R1569 B.n886 B.n885 10.6151
R1570 B.n888 B.n886 10.6151
R1571 B.n889 B.n888 10.6151
R1572 B.n890 B.n889 10.6151
R1573 B.n891 B.n890 10.6151
R1574 B.n893 B.n891 10.6151
R1575 B.n894 B.n893 10.6151
R1576 B.n895 B.n894 10.6151
R1577 B.n896 B.n895 10.6151
R1578 B.n898 B.n896 10.6151
R1579 B.n899 B.n898 10.6151
R1580 B.n900 B.n899 10.6151
R1581 B.n901 B.n900 10.6151
R1582 B.n903 B.n901 10.6151
R1583 B.n904 B.n903 10.6151
R1584 B.n905 B.n904 10.6151
R1585 B.n906 B.n905 10.6151
R1586 B.n907 B.n906 10.6151
R1587 B.n979 B.n1 10.6151
R1588 B.n979 B.n978 10.6151
R1589 B.n978 B.n977 10.6151
R1590 B.n977 B.n10 10.6151
R1591 B.n971 B.n10 10.6151
R1592 B.n971 B.n970 10.6151
R1593 B.n970 B.n969 10.6151
R1594 B.n969 B.n18 10.6151
R1595 B.n963 B.n18 10.6151
R1596 B.n963 B.n962 10.6151
R1597 B.n962 B.n961 10.6151
R1598 B.n961 B.n25 10.6151
R1599 B.n955 B.n25 10.6151
R1600 B.n955 B.n954 10.6151
R1601 B.n954 B.n953 10.6151
R1602 B.n953 B.n32 10.6151
R1603 B.n947 B.n32 10.6151
R1604 B.n947 B.n946 10.6151
R1605 B.n946 B.n945 10.6151
R1606 B.n945 B.n38 10.6151
R1607 B.n939 B.n38 10.6151
R1608 B.n939 B.n938 10.6151
R1609 B.n938 B.n937 10.6151
R1610 B.n937 B.n46 10.6151
R1611 B.n931 B.n46 10.6151
R1612 B.n931 B.n930 10.6151
R1613 B.n930 B.n929 10.6151
R1614 B.n929 B.n53 10.6151
R1615 B.n923 B.n53 10.6151
R1616 B.n923 B.n922 10.6151
R1617 B.n922 B.n921 10.6151
R1618 B.n921 B.n60 10.6151
R1619 B.n915 B.n60 10.6151
R1620 B.n915 B.n914 10.6151
R1621 B.n913 B.n67 10.6151
R1622 B.n137 B.n67 10.6151
R1623 B.n138 B.n137 10.6151
R1624 B.n141 B.n138 10.6151
R1625 B.n142 B.n141 10.6151
R1626 B.n145 B.n142 10.6151
R1627 B.n146 B.n145 10.6151
R1628 B.n149 B.n146 10.6151
R1629 B.n150 B.n149 10.6151
R1630 B.n153 B.n150 10.6151
R1631 B.n154 B.n153 10.6151
R1632 B.n157 B.n154 10.6151
R1633 B.n158 B.n157 10.6151
R1634 B.n161 B.n158 10.6151
R1635 B.n162 B.n161 10.6151
R1636 B.n165 B.n162 10.6151
R1637 B.n166 B.n165 10.6151
R1638 B.n169 B.n166 10.6151
R1639 B.n170 B.n169 10.6151
R1640 B.n173 B.n170 10.6151
R1641 B.n174 B.n173 10.6151
R1642 B.n177 B.n174 10.6151
R1643 B.n178 B.n177 10.6151
R1644 B.n181 B.n178 10.6151
R1645 B.n182 B.n181 10.6151
R1646 B.n185 B.n182 10.6151
R1647 B.n186 B.n185 10.6151
R1648 B.n189 B.n186 10.6151
R1649 B.n190 B.n189 10.6151
R1650 B.n193 B.n190 10.6151
R1651 B.n194 B.n193 10.6151
R1652 B.n197 B.n194 10.6151
R1653 B.n198 B.n197 10.6151
R1654 B.n201 B.n198 10.6151
R1655 B.n202 B.n201 10.6151
R1656 B.n205 B.n202 10.6151
R1657 B.n206 B.n205 10.6151
R1658 B.n209 B.n206 10.6151
R1659 B.n210 B.n209 10.6151
R1660 B.n213 B.n210 10.6151
R1661 B.n214 B.n213 10.6151
R1662 B.n217 B.n214 10.6151
R1663 B.n218 B.n217 10.6151
R1664 B.n221 B.n218 10.6151
R1665 B.n222 B.n221 10.6151
R1666 B.n225 B.n222 10.6151
R1667 B.n226 B.n225 10.6151
R1668 B.n229 B.n226 10.6151
R1669 B.n230 B.n229 10.6151
R1670 B.n233 B.n230 10.6151
R1671 B.n234 B.n233 10.6151
R1672 B.n237 B.n234 10.6151
R1673 B.n238 B.n237 10.6151
R1674 B.n241 B.n238 10.6151
R1675 B.n242 B.n241 10.6151
R1676 B.n245 B.n242 10.6151
R1677 B.n250 B.n247 10.6151
R1678 B.n251 B.n250 10.6151
R1679 B.n254 B.n251 10.6151
R1680 B.n255 B.n254 10.6151
R1681 B.n258 B.n255 10.6151
R1682 B.n259 B.n258 10.6151
R1683 B.n262 B.n259 10.6151
R1684 B.n263 B.n262 10.6151
R1685 B.n267 B.n266 10.6151
R1686 B.n270 B.n267 10.6151
R1687 B.n271 B.n270 10.6151
R1688 B.n274 B.n271 10.6151
R1689 B.n275 B.n274 10.6151
R1690 B.n278 B.n275 10.6151
R1691 B.n279 B.n278 10.6151
R1692 B.n282 B.n279 10.6151
R1693 B.n283 B.n282 10.6151
R1694 B.n286 B.n283 10.6151
R1695 B.n287 B.n286 10.6151
R1696 B.n290 B.n287 10.6151
R1697 B.n291 B.n290 10.6151
R1698 B.n294 B.n291 10.6151
R1699 B.n295 B.n294 10.6151
R1700 B.n298 B.n295 10.6151
R1701 B.n299 B.n298 10.6151
R1702 B.n302 B.n299 10.6151
R1703 B.n303 B.n302 10.6151
R1704 B.n306 B.n303 10.6151
R1705 B.n307 B.n306 10.6151
R1706 B.n310 B.n307 10.6151
R1707 B.n311 B.n310 10.6151
R1708 B.n314 B.n311 10.6151
R1709 B.n315 B.n314 10.6151
R1710 B.n318 B.n315 10.6151
R1711 B.n319 B.n318 10.6151
R1712 B.n322 B.n319 10.6151
R1713 B.n323 B.n322 10.6151
R1714 B.n326 B.n323 10.6151
R1715 B.n327 B.n326 10.6151
R1716 B.n330 B.n327 10.6151
R1717 B.n331 B.n330 10.6151
R1718 B.n334 B.n331 10.6151
R1719 B.n335 B.n334 10.6151
R1720 B.n338 B.n335 10.6151
R1721 B.n339 B.n338 10.6151
R1722 B.n342 B.n339 10.6151
R1723 B.n343 B.n342 10.6151
R1724 B.n346 B.n343 10.6151
R1725 B.n347 B.n346 10.6151
R1726 B.n350 B.n347 10.6151
R1727 B.n351 B.n350 10.6151
R1728 B.n354 B.n351 10.6151
R1729 B.n355 B.n354 10.6151
R1730 B.n358 B.n355 10.6151
R1731 B.n359 B.n358 10.6151
R1732 B.n362 B.n359 10.6151
R1733 B.n363 B.n362 10.6151
R1734 B.n366 B.n363 10.6151
R1735 B.n367 B.n366 10.6151
R1736 B.n370 B.n367 10.6151
R1737 B.n371 B.n370 10.6151
R1738 B.n374 B.n371 10.6151
R1739 B.n375 B.n374 10.6151
R1740 B.n908 B.n375 10.6151
R1741 B.n987 B.n0 8.11757
R1742 B.n987 B.n1 8.11757
R1743 B.n642 B.n508 6.5566
R1744 B.n626 B.n625 6.5566
R1745 B.n247 B.n246 6.5566
R1746 B.n263 B.n133 6.5566
R1747 B.n778 B.t7 6.383
R1748 B.n927 B.t11 6.383
R1749 B.n809 B.t4 5.40108
R1750 B.n949 B.t2 5.40108
R1751 B.n645 B.n508 4.05904
R1752 B.n625 B.n624 4.05904
R1753 B.n246 B.n245 4.05904
R1754 B.n266 B.n133 4.05904
R1755 VN.n2 VN.t0 240.774
R1756 VN.n14 VN.t3 240.774
R1757 VN.n3 VN.t2 207.454
R1758 VN.n10 VN.t1 207.454
R1759 VN.n15 VN.t4 207.454
R1760 VN.n22 VN.t5 207.454
R1761 VN.n21 VN.n12 161.3
R1762 VN.n20 VN.n19 161.3
R1763 VN.n18 VN.n13 161.3
R1764 VN.n17 VN.n16 161.3
R1765 VN.n9 VN.n0 161.3
R1766 VN.n8 VN.n7 161.3
R1767 VN.n6 VN.n1 161.3
R1768 VN.n5 VN.n4 161.3
R1769 VN.n11 VN.n10 95.0976
R1770 VN.n23 VN.n22 95.0976
R1771 VN.n8 VN.n1 56.0336
R1772 VN.n20 VN.n13 56.0336
R1773 VN VN.n23 50.4072
R1774 VN.n15 VN.n14 45.7215
R1775 VN.n3 VN.n2 45.7215
R1776 VN.n4 VN.n1 24.9531
R1777 VN.n16 VN.n13 24.9531
R1778 VN.n4 VN.n3 24.4675
R1779 VN.n9 VN.n8 24.4675
R1780 VN.n16 VN.n15 24.4675
R1781 VN.n21 VN.n20 24.4675
R1782 VN.n10 VN.n9 15.6594
R1783 VN.n22 VN.n21 15.6594
R1784 VN.n17 VN.n14 9.37527
R1785 VN.n5 VN.n2 9.37527
R1786 VN.n23 VN.n12 0.278367
R1787 VN.n11 VN.n0 0.278367
R1788 VN.n19 VN.n12 0.189894
R1789 VN.n19 VN.n18 0.189894
R1790 VN.n18 VN.n17 0.189894
R1791 VN.n6 VN.n5 0.189894
R1792 VN.n7 VN.n6 0.189894
R1793 VN.n7 VN.n0 0.189894
R1794 VN VN.n11 0.153454
R1795 VDD2.n1 VDD2.t5 62.7206
R1796 VDD2.n2 VDD2.t0 61.276
R1797 VDD2.n1 VDD2.n0 60.5647
R1798 VDD2 VDD2.n3 60.5619
R1799 VDD2.n2 VDD2.n1 44.9825
R1800 VDD2 VDD2.n2 1.55869
R1801 VDD2.n3 VDD2.t1 1.15637
R1802 VDD2.n3 VDD2.t2 1.15637
R1803 VDD2.n0 VDD2.t3 1.15637
R1804 VDD2.n0 VDD2.t4 1.15637
C0 VN VTAIL 8.70401f
C1 VN VDD2 8.90251f
C2 VTAIL VDD1 9.804389f
C3 VDD2 VDD1 1.1822f
C4 VTAIL VP 8.71846f
C5 VN VDD1 0.149961f
C6 VP VDD2 0.407194f
C7 VN VP 7.28854f
C8 VP VDD1 9.15524f
C9 VTAIL VDD2 9.84883f
C10 VDD2 B 6.424587f
C11 VDD1 B 6.722343f
C12 VTAIL B 9.423057f
C13 VN B 11.62803f
C14 VP B 10.026037f
C15 VDD2.t5 B 3.35589f
C16 VDD2.t3 B 0.288317f
C17 VDD2.t4 B 0.288317f
C18 VDD2.n0 B 2.62308f
C19 VDD2.n1 B 2.52958f
C20 VDD2.t0 B 3.34798f
C21 VDD2.n2 B 2.5792f
C22 VDD2.t1 B 0.288317f
C23 VDD2.t2 B 0.288317f
C24 VDD2.n3 B 2.62305f
C25 VN.n0 B 0.035146f
C26 VN.t1 B 2.49712f
C27 VN.n1 B 0.031829f
C28 VN.t0 B 2.63662f
C29 VN.n2 B 0.933806f
C30 VN.t2 B 2.49712f
C31 VN.n3 B 0.950925f
C32 VN.n4 B 0.05015f
C33 VN.n5 B 0.221588f
C34 VN.n6 B 0.026658f
C35 VN.n7 B 0.026658f
C36 VN.n8 B 0.045535f
C37 VN.n9 B 0.040853f
C38 VN.n10 B 0.948428f
C39 VN.n11 B 0.035202f
C40 VN.n12 B 0.035146f
C41 VN.t5 B 2.49712f
C42 VN.n13 B 0.031829f
C43 VN.t3 B 2.63662f
C44 VN.n14 B 0.933806f
C45 VN.t4 B 2.49712f
C46 VN.n15 B 0.950925f
C47 VN.n16 B 0.05015f
C48 VN.n17 B 0.221588f
C49 VN.n18 B 0.026658f
C50 VN.n19 B 0.026658f
C51 VN.n20 B 0.045535f
C52 VN.n21 B 0.040853f
C53 VN.n22 B 0.948428f
C54 VN.n23 B 1.49359f
C55 VDD1.t5 B 3.39626f
C56 VDD1.t2 B 3.39544f
C57 VDD1.t0 B 0.291715f
C58 VDD1.t1 B 0.291715f
C59 VDD1.n0 B 2.654f
C60 VDD1.n1 B 2.65541f
C61 VDD1.t3 B 0.291715f
C62 VDD1.t4 B 0.291715f
C63 VDD1.n2 B 2.65136f
C64 VDD1.n3 B 2.59503f
C65 VTAIL.t1 B 0.303602f
C66 VTAIL.t0 B 0.303602f
C67 VTAIL.n0 B 2.68945f
C68 VTAIL.n1 B 0.372525f
C69 VTAIL.t9 B 3.43415f
C70 VTAIL.n2 B 0.560029f
C71 VTAIL.t7 B 0.303602f
C72 VTAIL.t10 B 0.303602f
C73 VTAIL.n3 B 2.68945f
C74 VTAIL.n4 B 2.03144f
C75 VTAIL.t4 B 0.303602f
C76 VTAIL.t11 B 0.303602f
C77 VTAIL.n5 B 2.68945f
C78 VTAIL.n6 B 2.03144f
C79 VTAIL.t3 B 3.43417f
C80 VTAIL.n7 B 0.560007f
C81 VTAIL.t8 B 0.303602f
C82 VTAIL.t6 B 0.303602f
C83 VTAIL.n8 B 2.68945f
C84 VTAIL.n9 B 0.476719f
C85 VTAIL.t5 B 3.43415f
C86 VTAIL.n10 B 1.97021f
C87 VTAIL.t2 B 3.43415f
C88 VTAIL.n11 B 1.92987f
C89 VP.n0 B 0.035623f
C90 VP.t4 B 2.53102f
C91 VP.n1 B 0.032261f
C92 VP.n2 B 0.02702f
C93 VP.t5 B 2.53102f
C94 VP.n3 B 0.032261f
C95 VP.n4 B 0.035623f
C96 VP.t3 B 2.53102f
C97 VP.n5 B 0.035623f
C98 VP.t1 B 2.53102f
C99 VP.n6 B 0.032261f
C100 VP.t0 B 2.6724f
C101 VP.n7 B 0.946481f
C102 VP.t2 B 2.53102f
C103 VP.n8 B 0.963832f
C104 VP.n9 B 0.050831f
C105 VP.n10 B 0.224596f
C106 VP.n11 B 0.02702f
C107 VP.n12 B 0.02702f
C108 VP.n13 B 0.046154f
C109 VP.n14 B 0.041407f
C110 VP.n15 B 0.961302f
C111 VP.n16 B 1.49934f
C112 VP.n17 B 1.51872f
C113 VP.n18 B 0.961302f
C114 VP.n19 B 0.041407f
C115 VP.n20 B 0.046154f
C116 VP.n21 B 0.02702f
C117 VP.n22 B 0.02702f
C118 VP.n23 B 0.02702f
C119 VP.n24 B 0.050831f
C120 VP.n25 B 0.910774f
C121 VP.n26 B 0.050831f
C122 VP.n27 B 0.02702f
C123 VP.n28 B 0.02702f
C124 VP.n29 B 0.02702f
C125 VP.n30 B 0.046154f
C126 VP.n31 B 0.041407f
C127 VP.n32 B 0.961302f
C128 VP.n33 B 0.035679f
.ends

