* NGSPICE file created from diff_pair_sample_1261.ext - technology: sky130A

.subckt diff_pair_sample_1261 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=2.21
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=2.21
X2 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=2.21
X3 VTAIL.t7 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=2.21
X4 VDD1.t1 VP.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=2.21
X5 VTAIL.t3 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=2.21
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=2.21
X7 VTAIL.t4 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=2.21
X8 VDD2.t2 VN.t1 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=2.21
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0 ps=0 w=0.7 l=2.21
X10 VTAIL.t1 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.273 pd=2.18 as=0.1155 ps=1.03 w=0.7 l=2.21
X11 VDD2.t0 VN.t3 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.03 as=0.273 ps=2.18 w=0.7 l=2.21
R0 B.n336 B.n335 585
R1 B.n338 B.n76 585
R2 B.n341 B.n340 585
R3 B.n342 B.n75 585
R4 B.n344 B.n343 585
R5 B.n346 B.n74 585
R6 B.n348 B.n347 585
R7 B.n350 B.n349 585
R8 B.n353 B.n352 585
R9 B.n354 B.n69 585
R10 B.n356 B.n355 585
R11 B.n358 B.n68 585
R12 B.n361 B.n360 585
R13 B.n362 B.n67 585
R14 B.n364 B.n363 585
R15 B.n366 B.n66 585
R16 B.n369 B.n368 585
R17 B.n370 B.n63 585
R18 B.n373 B.n372 585
R19 B.n375 B.n62 585
R20 B.n378 B.n377 585
R21 B.n379 B.n61 585
R22 B.n381 B.n380 585
R23 B.n383 B.n60 585
R24 B.n386 B.n385 585
R25 B.n387 B.n59 585
R26 B.n334 B.n57 585
R27 B.n390 B.n57 585
R28 B.n333 B.n56 585
R29 B.n391 B.n56 585
R30 B.n332 B.n55 585
R31 B.n392 B.n55 585
R32 B.n331 B.n330 585
R33 B.n330 B.n51 585
R34 B.n329 B.n50 585
R35 B.n398 B.n50 585
R36 B.n328 B.n49 585
R37 B.n399 B.n49 585
R38 B.n327 B.n48 585
R39 B.n400 B.n48 585
R40 B.n326 B.n325 585
R41 B.n325 B.n47 585
R42 B.n324 B.n43 585
R43 B.n406 B.n43 585
R44 B.n323 B.n42 585
R45 B.n407 B.n42 585
R46 B.n322 B.n41 585
R47 B.n408 B.n41 585
R48 B.n321 B.n320 585
R49 B.n320 B.n37 585
R50 B.n319 B.n36 585
R51 B.n414 B.n36 585
R52 B.n318 B.n35 585
R53 B.n415 B.n35 585
R54 B.n317 B.n34 585
R55 B.n416 B.n34 585
R56 B.n316 B.n315 585
R57 B.n315 B.n30 585
R58 B.n314 B.n29 585
R59 B.n422 B.n29 585
R60 B.n313 B.n28 585
R61 B.n423 B.n28 585
R62 B.n312 B.n27 585
R63 B.n424 B.n27 585
R64 B.n311 B.n310 585
R65 B.n310 B.n23 585
R66 B.n309 B.n22 585
R67 B.n430 B.n22 585
R68 B.n308 B.n21 585
R69 B.n431 B.n21 585
R70 B.n307 B.n20 585
R71 B.n432 B.n20 585
R72 B.n306 B.n305 585
R73 B.n305 B.n16 585
R74 B.n304 B.n15 585
R75 B.n438 B.n15 585
R76 B.n303 B.n14 585
R77 B.n439 B.n14 585
R78 B.n302 B.n13 585
R79 B.n440 B.n13 585
R80 B.n301 B.n300 585
R81 B.n300 B.n12 585
R82 B.n299 B.n298 585
R83 B.n299 B.n8 585
R84 B.n297 B.n7 585
R85 B.n447 B.n7 585
R86 B.n296 B.n6 585
R87 B.n448 B.n6 585
R88 B.n295 B.n5 585
R89 B.n449 B.n5 585
R90 B.n294 B.n293 585
R91 B.n293 B.n4 585
R92 B.n292 B.n77 585
R93 B.n292 B.n291 585
R94 B.n282 B.n78 585
R95 B.n79 B.n78 585
R96 B.n284 B.n283 585
R97 B.n285 B.n284 585
R98 B.n281 B.n83 585
R99 B.n87 B.n83 585
R100 B.n280 B.n279 585
R101 B.n279 B.n278 585
R102 B.n85 B.n84 585
R103 B.n86 B.n85 585
R104 B.n271 B.n270 585
R105 B.n272 B.n271 585
R106 B.n269 B.n92 585
R107 B.n92 B.n91 585
R108 B.n268 B.n267 585
R109 B.n267 B.n266 585
R110 B.n94 B.n93 585
R111 B.n95 B.n94 585
R112 B.n259 B.n258 585
R113 B.n260 B.n259 585
R114 B.n257 B.n99 585
R115 B.n103 B.n99 585
R116 B.n256 B.n255 585
R117 B.n255 B.n254 585
R118 B.n101 B.n100 585
R119 B.n102 B.n101 585
R120 B.n247 B.n246 585
R121 B.n248 B.n247 585
R122 B.n245 B.n108 585
R123 B.n108 B.n107 585
R124 B.n244 B.n243 585
R125 B.n243 B.n242 585
R126 B.n110 B.n109 585
R127 B.n111 B.n110 585
R128 B.n235 B.n234 585
R129 B.n236 B.n235 585
R130 B.n233 B.n116 585
R131 B.n116 B.n115 585
R132 B.n232 B.n231 585
R133 B.n231 B.n230 585
R134 B.n118 B.n117 585
R135 B.n223 B.n118 585
R136 B.n222 B.n221 585
R137 B.n224 B.n222 585
R138 B.n220 B.n123 585
R139 B.n123 B.n122 585
R140 B.n219 B.n218 585
R141 B.n218 B.n217 585
R142 B.n125 B.n124 585
R143 B.n126 B.n125 585
R144 B.n210 B.n209 585
R145 B.n211 B.n210 585
R146 B.n208 B.n131 585
R147 B.n131 B.n130 585
R148 B.n207 B.n206 585
R149 B.n206 B.n205 585
R150 B.n202 B.n135 585
R151 B.n201 B.n200 585
R152 B.n198 B.n136 585
R153 B.n198 B.n134 585
R154 B.n197 B.n196 585
R155 B.n195 B.n194 585
R156 B.n193 B.n138 585
R157 B.n191 B.n190 585
R158 B.n189 B.n139 585
R159 B.n187 B.n186 585
R160 B.n184 B.n142 585
R161 B.n182 B.n181 585
R162 B.n180 B.n143 585
R163 B.n179 B.n178 585
R164 B.n176 B.n144 585
R165 B.n174 B.n173 585
R166 B.n172 B.n145 585
R167 B.n171 B.n170 585
R168 B.n168 B.n146 585
R169 B.n166 B.n165 585
R170 B.n164 B.n147 585
R171 B.n163 B.n162 585
R172 B.n160 B.n151 585
R173 B.n158 B.n157 585
R174 B.n156 B.n152 585
R175 B.n155 B.n154 585
R176 B.n133 B.n132 585
R177 B.n134 B.n133 585
R178 B.n204 B.n203 585
R179 B.n205 B.n204 585
R180 B.n129 B.n128 585
R181 B.n130 B.n129 585
R182 B.n213 B.n212 585
R183 B.n212 B.n211 585
R184 B.n214 B.n127 585
R185 B.n127 B.n126 585
R186 B.n216 B.n215 585
R187 B.n217 B.n216 585
R188 B.n121 B.n120 585
R189 B.n122 B.n121 585
R190 B.n226 B.n225 585
R191 B.n225 B.n224 585
R192 B.n227 B.n119 585
R193 B.n223 B.n119 585
R194 B.n229 B.n228 585
R195 B.n230 B.n229 585
R196 B.n114 B.n113 585
R197 B.n115 B.n114 585
R198 B.n238 B.n237 585
R199 B.n237 B.n236 585
R200 B.n239 B.n112 585
R201 B.n112 B.n111 585
R202 B.n241 B.n240 585
R203 B.n242 B.n241 585
R204 B.n106 B.n105 585
R205 B.n107 B.n106 585
R206 B.n250 B.n249 585
R207 B.n249 B.n248 585
R208 B.n251 B.n104 585
R209 B.n104 B.n102 585
R210 B.n253 B.n252 585
R211 B.n254 B.n253 585
R212 B.n98 B.n97 585
R213 B.n103 B.n98 585
R214 B.n262 B.n261 585
R215 B.n261 B.n260 585
R216 B.n263 B.n96 585
R217 B.n96 B.n95 585
R218 B.n265 B.n264 585
R219 B.n266 B.n265 585
R220 B.n90 B.n89 585
R221 B.n91 B.n90 585
R222 B.n274 B.n273 585
R223 B.n273 B.n272 585
R224 B.n275 B.n88 585
R225 B.n88 B.n86 585
R226 B.n277 B.n276 585
R227 B.n278 B.n277 585
R228 B.n82 B.n81 585
R229 B.n87 B.n82 585
R230 B.n287 B.n286 585
R231 B.n286 B.n285 585
R232 B.n288 B.n80 585
R233 B.n80 B.n79 585
R234 B.n290 B.n289 585
R235 B.n291 B.n290 585
R236 B.n3 B.n0 585
R237 B.n4 B.n3 585
R238 B.n446 B.n1 585
R239 B.n447 B.n446 585
R240 B.n445 B.n444 585
R241 B.n445 B.n8 585
R242 B.n443 B.n9 585
R243 B.n12 B.n9 585
R244 B.n442 B.n441 585
R245 B.n441 B.n440 585
R246 B.n11 B.n10 585
R247 B.n439 B.n11 585
R248 B.n437 B.n436 585
R249 B.n438 B.n437 585
R250 B.n435 B.n17 585
R251 B.n17 B.n16 585
R252 B.n434 B.n433 585
R253 B.n433 B.n432 585
R254 B.n19 B.n18 585
R255 B.n431 B.n19 585
R256 B.n429 B.n428 585
R257 B.n430 B.n429 585
R258 B.n427 B.n24 585
R259 B.n24 B.n23 585
R260 B.n426 B.n425 585
R261 B.n425 B.n424 585
R262 B.n26 B.n25 585
R263 B.n423 B.n26 585
R264 B.n421 B.n420 585
R265 B.n422 B.n421 585
R266 B.n419 B.n31 585
R267 B.n31 B.n30 585
R268 B.n418 B.n417 585
R269 B.n417 B.n416 585
R270 B.n33 B.n32 585
R271 B.n415 B.n33 585
R272 B.n413 B.n412 585
R273 B.n414 B.n413 585
R274 B.n411 B.n38 585
R275 B.n38 B.n37 585
R276 B.n410 B.n409 585
R277 B.n409 B.n408 585
R278 B.n40 B.n39 585
R279 B.n407 B.n40 585
R280 B.n405 B.n404 585
R281 B.n406 B.n405 585
R282 B.n403 B.n44 585
R283 B.n47 B.n44 585
R284 B.n402 B.n401 585
R285 B.n401 B.n400 585
R286 B.n46 B.n45 585
R287 B.n399 B.n46 585
R288 B.n397 B.n396 585
R289 B.n398 B.n397 585
R290 B.n395 B.n52 585
R291 B.n52 B.n51 585
R292 B.n394 B.n393 585
R293 B.n393 B.n392 585
R294 B.n54 B.n53 585
R295 B.n391 B.n54 585
R296 B.n389 B.n388 585
R297 B.n390 B.n389 585
R298 B.n450 B.n449 585
R299 B.n448 B.n2 585
R300 B.n389 B.n59 530.939
R301 B.n336 B.n57 530.939
R302 B.n206 B.n133 530.939
R303 B.n204 B.n135 530.939
R304 B.n64 B.t13 285.82
R305 B.n70 B.t6 285.82
R306 B.n148 B.t11 285.82
R307 B.n140 B.t17 285.82
R308 B.n337 B.n58 256.663
R309 B.n339 B.n58 256.663
R310 B.n345 B.n58 256.663
R311 B.n73 B.n58 256.663
R312 B.n351 B.n58 256.663
R313 B.n357 B.n58 256.663
R314 B.n359 B.n58 256.663
R315 B.n365 B.n58 256.663
R316 B.n367 B.n58 256.663
R317 B.n374 B.n58 256.663
R318 B.n376 B.n58 256.663
R319 B.n382 B.n58 256.663
R320 B.n384 B.n58 256.663
R321 B.n199 B.n134 256.663
R322 B.n137 B.n134 256.663
R323 B.n192 B.n134 256.663
R324 B.n185 B.n134 256.663
R325 B.n183 B.n134 256.663
R326 B.n177 B.n134 256.663
R327 B.n175 B.n134 256.663
R328 B.n169 B.n134 256.663
R329 B.n167 B.n134 256.663
R330 B.n161 B.n134 256.663
R331 B.n159 B.n134 256.663
R332 B.n153 B.n134 256.663
R333 B.n452 B.n451 256.663
R334 B.n65 B.t14 236.559
R335 B.n71 B.t7 236.559
R336 B.n149 B.t10 236.559
R337 B.n141 B.t16 236.559
R338 B.n205 B.n134 230.126
R339 B.n390 B.n58 230.126
R340 B.n64 B.t12 208.714
R341 B.n70 B.t4 208.714
R342 B.n148 B.t8 208.714
R343 B.n140 B.t15 208.714
R344 B.n385 B.n383 163.367
R345 B.n381 B.n61 163.367
R346 B.n377 B.n375 163.367
R347 B.n373 B.n63 163.367
R348 B.n368 B.n366 163.367
R349 B.n364 B.n67 163.367
R350 B.n360 B.n358 163.367
R351 B.n356 B.n69 163.367
R352 B.n352 B.n350 163.367
R353 B.n347 B.n346 163.367
R354 B.n344 B.n75 163.367
R355 B.n340 B.n338 163.367
R356 B.n206 B.n131 163.367
R357 B.n210 B.n131 163.367
R358 B.n210 B.n125 163.367
R359 B.n218 B.n125 163.367
R360 B.n218 B.n123 163.367
R361 B.n222 B.n123 163.367
R362 B.n222 B.n118 163.367
R363 B.n231 B.n118 163.367
R364 B.n231 B.n116 163.367
R365 B.n235 B.n116 163.367
R366 B.n235 B.n110 163.367
R367 B.n243 B.n110 163.367
R368 B.n243 B.n108 163.367
R369 B.n247 B.n108 163.367
R370 B.n247 B.n101 163.367
R371 B.n255 B.n101 163.367
R372 B.n255 B.n99 163.367
R373 B.n259 B.n99 163.367
R374 B.n259 B.n94 163.367
R375 B.n267 B.n94 163.367
R376 B.n267 B.n92 163.367
R377 B.n271 B.n92 163.367
R378 B.n271 B.n85 163.367
R379 B.n279 B.n85 163.367
R380 B.n279 B.n83 163.367
R381 B.n284 B.n83 163.367
R382 B.n284 B.n78 163.367
R383 B.n292 B.n78 163.367
R384 B.n293 B.n292 163.367
R385 B.n293 B.n5 163.367
R386 B.n6 B.n5 163.367
R387 B.n7 B.n6 163.367
R388 B.n299 B.n7 163.367
R389 B.n300 B.n299 163.367
R390 B.n300 B.n13 163.367
R391 B.n14 B.n13 163.367
R392 B.n15 B.n14 163.367
R393 B.n305 B.n15 163.367
R394 B.n305 B.n20 163.367
R395 B.n21 B.n20 163.367
R396 B.n22 B.n21 163.367
R397 B.n310 B.n22 163.367
R398 B.n310 B.n27 163.367
R399 B.n28 B.n27 163.367
R400 B.n29 B.n28 163.367
R401 B.n315 B.n29 163.367
R402 B.n315 B.n34 163.367
R403 B.n35 B.n34 163.367
R404 B.n36 B.n35 163.367
R405 B.n320 B.n36 163.367
R406 B.n320 B.n41 163.367
R407 B.n42 B.n41 163.367
R408 B.n43 B.n42 163.367
R409 B.n325 B.n43 163.367
R410 B.n325 B.n48 163.367
R411 B.n49 B.n48 163.367
R412 B.n50 B.n49 163.367
R413 B.n330 B.n50 163.367
R414 B.n330 B.n55 163.367
R415 B.n56 B.n55 163.367
R416 B.n57 B.n56 163.367
R417 B.n200 B.n198 163.367
R418 B.n198 B.n197 163.367
R419 B.n194 B.n193 163.367
R420 B.n191 B.n139 163.367
R421 B.n186 B.n184 163.367
R422 B.n182 B.n143 163.367
R423 B.n178 B.n176 163.367
R424 B.n174 B.n145 163.367
R425 B.n170 B.n168 163.367
R426 B.n166 B.n147 163.367
R427 B.n162 B.n160 163.367
R428 B.n158 B.n152 163.367
R429 B.n154 B.n133 163.367
R430 B.n204 B.n129 163.367
R431 B.n212 B.n129 163.367
R432 B.n212 B.n127 163.367
R433 B.n216 B.n127 163.367
R434 B.n216 B.n121 163.367
R435 B.n225 B.n121 163.367
R436 B.n225 B.n119 163.367
R437 B.n229 B.n119 163.367
R438 B.n229 B.n114 163.367
R439 B.n237 B.n114 163.367
R440 B.n237 B.n112 163.367
R441 B.n241 B.n112 163.367
R442 B.n241 B.n106 163.367
R443 B.n249 B.n106 163.367
R444 B.n249 B.n104 163.367
R445 B.n253 B.n104 163.367
R446 B.n253 B.n98 163.367
R447 B.n261 B.n98 163.367
R448 B.n261 B.n96 163.367
R449 B.n265 B.n96 163.367
R450 B.n265 B.n90 163.367
R451 B.n273 B.n90 163.367
R452 B.n273 B.n88 163.367
R453 B.n277 B.n88 163.367
R454 B.n277 B.n82 163.367
R455 B.n286 B.n82 163.367
R456 B.n286 B.n80 163.367
R457 B.n290 B.n80 163.367
R458 B.n290 B.n3 163.367
R459 B.n450 B.n3 163.367
R460 B.n446 B.n2 163.367
R461 B.n446 B.n445 163.367
R462 B.n445 B.n9 163.367
R463 B.n441 B.n9 163.367
R464 B.n441 B.n11 163.367
R465 B.n437 B.n11 163.367
R466 B.n437 B.n17 163.367
R467 B.n433 B.n17 163.367
R468 B.n433 B.n19 163.367
R469 B.n429 B.n19 163.367
R470 B.n429 B.n24 163.367
R471 B.n425 B.n24 163.367
R472 B.n425 B.n26 163.367
R473 B.n421 B.n26 163.367
R474 B.n421 B.n31 163.367
R475 B.n417 B.n31 163.367
R476 B.n417 B.n33 163.367
R477 B.n413 B.n33 163.367
R478 B.n413 B.n38 163.367
R479 B.n409 B.n38 163.367
R480 B.n409 B.n40 163.367
R481 B.n405 B.n40 163.367
R482 B.n405 B.n44 163.367
R483 B.n401 B.n44 163.367
R484 B.n401 B.n46 163.367
R485 B.n397 B.n46 163.367
R486 B.n397 B.n52 163.367
R487 B.n393 B.n52 163.367
R488 B.n393 B.n54 163.367
R489 B.n389 B.n54 163.367
R490 B.n205 B.n130 125.189
R491 B.n211 B.n130 125.189
R492 B.n211 B.n126 125.189
R493 B.n217 B.n126 125.189
R494 B.n217 B.n122 125.189
R495 B.n224 B.n122 125.189
R496 B.n224 B.n223 125.189
R497 B.n230 B.n115 125.189
R498 B.n236 B.n115 125.189
R499 B.n236 B.n111 125.189
R500 B.n242 B.n111 125.189
R501 B.n242 B.n107 125.189
R502 B.n248 B.n107 125.189
R503 B.n248 B.n102 125.189
R504 B.n254 B.n102 125.189
R505 B.n254 B.n103 125.189
R506 B.n260 B.n95 125.189
R507 B.n266 B.n95 125.189
R508 B.n266 B.n91 125.189
R509 B.n272 B.n91 125.189
R510 B.n272 B.n86 125.189
R511 B.n278 B.n86 125.189
R512 B.n278 B.n87 125.189
R513 B.n285 B.n79 125.189
R514 B.n291 B.n79 125.189
R515 B.n291 B.n4 125.189
R516 B.n449 B.n4 125.189
R517 B.n449 B.n448 125.189
R518 B.n448 B.n447 125.189
R519 B.n447 B.n8 125.189
R520 B.n12 B.n8 125.189
R521 B.n440 B.n12 125.189
R522 B.n439 B.n438 125.189
R523 B.n438 B.n16 125.189
R524 B.n432 B.n16 125.189
R525 B.n432 B.n431 125.189
R526 B.n431 B.n430 125.189
R527 B.n430 B.n23 125.189
R528 B.n424 B.n23 125.189
R529 B.n423 B.n422 125.189
R530 B.n422 B.n30 125.189
R531 B.n416 B.n30 125.189
R532 B.n416 B.n415 125.189
R533 B.n415 B.n414 125.189
R534 B.n414 B.n37 125.189
R535 B.n408 B.n37 125.189
R536 B.n408 B.n407 125.189
R537 B.n407 B.n406 125.189
R538 B.n400 B.n47 125.189
R539 B.n400 B.n399 125.189
R540 B.n399 B.n398 125.189
R541 B.n398 B.n51 125.189
R542 B.n392 B.n51 125.189
R543 B.n392 B.n391 125.189
R544 B.n391 B.n390 125.189
R545 B.n230 B.t9 123.347
R546 B.n406 B.t5 123.347
R547 B.n285 B.t2 104.938
R548 B.n440 B.t3 104.938
R549 B.n103 B.t0 86.5277
R550 B.t1 B.n423 86.5277
R551 B.n384 B.n59 71.676
R552 B.n383 B.n382 71.676
R553 B.n376 B.n61 71.676
R554 B.n375 B.n374 71.676
R555 B.n367 B.n63 71.676
R556 B.n366 B.n365 71.676
R557 B.n359 B.n67 71.676
R558 B.n358 B.n357 71.676
R559 B.n351 B.n69 71.676
R560 B.n350 B.n73 71.676
R561 B.n346 B.n345 71.676
R562 B.n339 B.n75 71.676
R563 B.n338 B.n337 71.676
R564 B.n337 B.n336 71.676
R565 B.n340 B.n339 71.676
R566 B.n345 B.n344 71.676
R567 B.n347 B.n73 71.676
R568 B.n352 B.n351 71.676
R569 B.n357 B.n356 71.676
R570 B.n360 B.n359 71.676
R571 B.n365 B.n364 71.676
R572 B.n368 B.n367 71.676
R573 B.n374 B.n373 71.676
R574 B.n377 B.n376 71.676
R575 B.n382 B.n381 71.676
R576 B.n385 B.n384 71.676
R577 B.n199 B.n135 71.676
R578 B.n197 B.n137 71.676
R579 B.n193 B.n192 71.676
R580 B.n185 B.n139 71.676
R581 B.n184 B.n183 71.676
R582 B.n177 B.n143 71.676
R583 B.n176 B.n175 71.676
R584 B.n169 B.n145 71.676
R585 B.n168 B.n167 71.676
R586 B.n161 B.n147 71.676
R587 B.n160 B.n159 71.676
R588 B.n153 B.n152 71.676
R589 B.n200 B.n199 71.676
R590 B.n194 B.n137 71.676
R591 B.n192 B.n191 71.676
R592 B.n186 B.n185 71.676
R593 B.n183 B.n182 71.676
R594 B.n178 B.n177 71.676
R595 B.n175 B.n174 71.676
R596 B.n170 B.n169 71.676
R597 B.n167 B.n166 71.676
R598 B.n162 B.n161 71.676
R599 B.n159 B.n158 71.676
R600 B.n154 B.n153 71.676
R601 B.n451 B.n450 71.676
R602 B.n451 B.n2 71.676
R603 B.n371 B.n65 59.5399
R604 B.n72 B.n71 59.5399
R605 B.n150 B.n149 59.5399
R606 B.n188 B.n141 59.5399
R607 B.n65 B.n64 49.2611
R608 B.n71 B.n70 49.2611
R609 B.n149 B.n148 49.2611
R610 B.n141 B.n140 49.2611
R611 B.n260 B.t0 38.6616
R612 B.n424 B.t1 38.6616
R613 B.n203 B.n202 34.4981
R614 B.n207 B.n132 34.4981
R615 B.n335 B.n334 34.4981
R616 B.n388 B.n387 34.4981
R617 B.n87 B.t2 20.2515
R618 B.t3 B.n439 20.2515
R619 B B.n452 18.0485
R620 B.n203 B.n128 10.6151
R621 B.n213 B.n128 10.6151
R622 B.n214 B.n213 10.6151
R623 B.n215 B.n214 10.6151
R624 B.n215 B.n120 10.6151
R625 B.n226 B.n120 10.6151
R626 B.n227 B.n226 10.6151
R627 B.n228 B.n227 10.6151
R628 B.n228 B.n113 10.6151
R629 B.n238 B.n113 10.6151
R630 B.n239 B.n238 10.6151
R631 B.n240 B.n239 10.6151
R632 B.n240 B.n105 10.6151
R633 B.n250 B.n105 10.6151
R634 B.n251 B.n250 10.6151
R635 B.n252 B.n251 10.6151
R636 B.n252 B.n97 10.6151
R637 B.n262 B.n97 10.6151
R638 B.n263 B.n262 10.6151
R639 B.n264 B.n263 10.6151
R640 B.n264 B.n89 10.6151
R641 B.n274 B.n89 10.6151
R642 B.n275 B.n274 10.6151
R643 B.n276 B.n275 10.6151
R644 B.n276 B.n81 10.6151
R645 B.n287 B.n81 10.6151
R646 B.n288 B.n287 10.6151
R647 B.n289 B.n288 10.6151
R648 B.n289 B.n0 10.6151
R649 B.n202 B.n201 10.6151
R650 B.n201 B.n136 10.6151
R651 B.n196 B.n136 10.6151
R652 B.n196 B.n195 10.6151
R653 B.n195 B.n138 10.6151
R654 B.n190 B.n138 10.6151
R655 B.n190 B.n189 10.6151
R656 B.n187 B.n142 10.6151
R657 B.n181 B.n142 10.6151
R658 B.n181 B.n180 10.6151
R659 B.n180 B.n179 10.6151
R660 B.n179 B.n144 10.6151
R661 B.n173 B.n144 10.6151
R662 B.n173 B.n172 10.6151
R663 B.n172 B.n171 10.6151
R664 B.n171 B.n146 10.6151
R665 B.n165 B.n164 10.6151
R666 B.n164 B.n163 10.6151
R667 B.n163 B.n151 10.6151
R668 B.n157 B.n151 10.6151
R669 B.n157 B.n156 10.6151
R670 B.n156 B.n155 10.6151
R671 B.n155 B.n132 10.6151
R672 B.n208 B.n207 10.6151
R673 B.n209 B.n208 10.6151
R674 B.n209 B.n124 10.6151
R675 B.n219 B.n124 10.6151
R676 B.n220 B.n219 10.6151
R677 B.n221 B.n220 10.6151
R678 B.n221 B.n117 10.6151
R679 B.n232 B.n117 10.6151
R680 B.n233 B.n232 10.6151
R681 B.n234 B.n233 10.6151
R682 B.n234 B.n109 10.6151
R683 B.n244 B.n109 10.6151
R684 B.n245 B.n244 10.6151
R685 B.n246 B.n245 10.6151
R686 B.n246 B.n100 10.6151
R687 B.n256 B.n100 10.6151
R688 B.n257 B.n256 10.6151
R689 B.n258 B.n257 10.6151
R690 B.n258 B.n93 10.6151
R691 B.n268 B.n93 10.6151
R692 B.n269 B.n268 10.6151
R693 B.n270 B.n269 10.6151
R694 B.n270 B.n84 10.6151
R695 B.n280 B.n84 10.6151
R696 B.n281 B.n280 10.6151
R697 B.n283 B.n281 10.6151
R698 B.n283 B.n282 10.6151
R699 B.n282 B.n77 10.6151
R700 B.n294 B.n77 10.6151
R701 B.n295 B.n294 10.6151
R702 B.n296 B.n295 10.6151
R703 B.n297 B.n296 10.6151
R704 B.n298 B.n297 10.6151
R705 B.n301 B.n298 10.6151
R706 B.n302 B.n301 10.6151
R707 B.n303 B.n302 10.6151
R708 B.n304 B.n303 10.6151
R709 B.n306 B.n304 10.6151
R710 B.n307 B.n306 10.6151
R711 B.n308 B.n307 10.6151
R712 B.n309 B.n308 10.6151
R713 B.n311 B.n309 10.6151
R714 B.n312 B.n311 10.6151
R715 B.n313 B.n312 10.6151
R716 B.n314 B.n313 10.6151
R717 B.n316 B.n314 10.6151
R718 B.n317 B.n316 10.6151
R719 B.n318 B.n317 10.6151
R720 B.n319 B.n318 10.6151
R721 B.n321 B.n319 10.6151
R722 B.n322 B.n321 10.6151
R723 B.n323 B.n322 10.6151
R724 B.n324 B.n323 10.6151
R725 B.n326 B.n324 10.6151
R726 B.n327 B.n326 10.6151
R727 B.n328 B.n327 10.6151
R728 B.n329 B.n328 10.6151
R729 B.n331 B.n329 10.6151
R730 B.n332 B.n331 10.6151
R731 B.n333 B.n332 10.6151
R732 B.n334 B.n333 10.6151
R733 B.n444 B.n1 10.6151
R734 B.n444 B.n443 10.6151
R735 B.n443 B.n442 10.6151
R736 B.n442 B.n10 10.6151
R737 B.n436 B.n10 10.6151
R738 B.n436 B.n435 10.6151
R739 B.n435 B.n434 10.6151
R740 B.n434 B.n18 10.6151
R741 B.n428 B.n18 10.6151
R742 B.n428 B.n427 10.6151
R743 B.n427 B.n426 10.6151
R744 B.n426 B.n25 10.6151
R745 B.n420 B.n25 10.6151
R746 B.n420 B.n419 10.6151
R747 B.n419 B.n418 10.6151
R748 B.n418 B.n32 10.6151
R749 B.n412 B.n32 10.6151
R750 B.n412 B.n411 10.6151
R751 B.n411 B.n410 10.6151
R752 B.n410 B.n39 10.6151
R753 B.n404 B.n39 10.6151
R754 B.n404 B.n403 10.6151
R755 B.n403 B.n402 10.6151
R756 B.n402 B.n45 10.6151
R757 B.n396 B.n45 10.6151
R758 B.n396 B.n395 10.6151
R759 B.n395 B.n394 10.6151
R760 B.n394 B.n53 10.6151
R761 B.n388 B.n53 10.6151
R762 B.n387 B.n386 10.6151
R763 B.n386 B.n60 10.6151
R764 B.n380 B.n60 10.6151
R765 B.n380 B.n379 10.6151
R766 B.n379 B.n378 10.6151
R767 B.n378 B.n62 10.6151
R768 B.n372 B.n62 10.6151
R769 B.n370 B.n369 10.6151
R770 B.n369 B.n66 10.6151
R771 B.n363 B.n66 10.6151
R772 B.n363 B.n362 10.6151
R773 B.n362 B.n361 10.6151
R774 B.n361 B.n68 10.6151
R775 B.n355 B.n68 10.6151
R776 B.n355 B.n354 10.6151
R777 B.n354 B.n353 10.6151
R778 B.n349 B.n348 10.6151
R779 B.n348 B.n74 10.6151
R780 B.n343 B.n74 10.6151
R781 B.n343 B.n342 10.6151
R782 B.n342 B.n341 10.6151
R783 B.n341 B.n76 10.6151
R784 B.n335 B.n76 10.6151
R785 B.n189 B.n188 9.36635
R786 B.n165 B.n150 9.36635
R787 B.n372 B.n371 9.36635
R788 B.n349 B.n72 9.36635
R789 B.n452 B.n0 8.11757
R790 B.n452 B.n1 8.11757
R791 B.n223 B.t9 1.8415
R792 B.n47 B.t5 1.8415
R793 B.n188 B.n187 1.24928
R794 B.n150 B.n146 1.24928
R795 B.n371 B.n370 1.24928
R796 B.n353 B.n72 1.24928
R797 VP.n12 VP.n0 161.3
R798 VP.n11 VP.n10 161.3
R799 VP.n9 VP.n1 161.3
R800 VP.n8 VP.n7 161.3
R801 VP.n6 VP.n2 161.3
R802 VP.n5 VP.n4 97.6287
R803 VP.n14 VP.n13 97.6287
R804 VP.n3 VP.t3 43.4633
R805 VP.n3 VP.t2 42.8245
R806 VP.n4 VP.n3 42.2806
R807 VP.n7 VP.n1 40.577
R808 VP.n11 VP.n1 40.577
R809 VP.n7 VP.n6 24.5923
R810 VP.n12 VP.n11 24.5923
R811 VP.n6 VP.n5 13.2801
R812 VP.n13 VP.n12 13.2801
R813 VP.n5 VP.t1 7.63398
R814 VP.n13 VP.t0 7.63398
R815 VP.n4 VP.n2 0.278335
R816 VP.n14 VP.n0 0.278335
R817 VP.n8 VP.n2 0.189894
R818 VP.n9 VP.n8 0.189894
R819 VP.n10 VP.n9 0.189894
R820 VP.n10 VP.n0 0.189894
R821 VP VP.n14 0.153485
R822 VTAIL.n7 VTAIL.t2 247.411
R823 VTAIL.n0 VTAIL.t1 247.411
R824 VTAIL.n1 VTAIL.t5 247.411
R825 VTAIL.n2 VTAIL.t7 247.411
R826 VTAIL.n6 VTAIL.t6 247.411
R827 VTAIL.n5 VTAIL.t4 247.411
R828 VTAIL.n4 VTAIL.t0 247.411
R829 VTAIL.n3 VTAIL.t3 247.411
R830 VTAIL.n7 VTAIL.n6 15.16
R831 VTAIL.n3 VTAIL.n2 15.16
R832 VTAIL.n4 VTAIL.n3 2.19016
R833 VTAIL.n6 VTAIL.n5 2.19016
R834 VTAIL.n2 VTAIL.n1 2.19016
R835 VTAIL VTAIL.n0 1.15352
R836 VTAIL VTAIL.n7 1.03714
R837 VTAIL.n5 VTAIL.n4 0.470328
R838 VTAIL.n1 VTAIL.n0 0.470328
R839 VDD1 VDD1.n1 267.216
R840 VDD1 VDD1.n0 235.862
R841 VDD1.n0 VDD1.t0 28.2862
R842 VDD1.n0 VDD1.t1 28.2862
R843 VDD1.n1 VDD1.t2 28.2862
R844 VDD1.n1 VDD1.t3 28.2862
R845 VN.n0 VN.t2 43.4633
R846 VN.n1 VN.t1 43.4633
R847 VN.n0 VN.t3 42.8245
R848 VN.n1 VN.t0 42.8245
R849 VN VN.n1 42.5594
R850 VN VN.n0 5.79803
R851 VDD2.n2 VDD2.n0 266.69
R852 VDD2.n2 VDD2.n1 235.804
R853 VDD2.n1 VDD2.t3 28.2862
R854 VDD2.n1 VDD2.t2 28.2862
R855 VDD2.n0 VDD2.t1 28.2862
R856 VDD2.n0 VDD2.t0 28.2862
R857 VDD2 VDD2.n2 0.0586897
C0 VDD1 VTAIL 2.50374f
C1 VDD2 VP 0.378753f
C2 VN VP 3.82591f
C3 VDD1 VDD2 0.93484f
C4 VTAIL VDD2 2.55534f
C5 VN VDD1 0.15633f
C6 VN VTAIL 1.21938f
C7 VN VDD2 0.578514f
C8 VDD1 VP 0.798518f
C9 VTAIL VP 1.23349f
C10 VDD2 B 2.641494f
C11 VDD1 B 4.99871f
C12 VTAIL B 2.681313f
C13 VN B 8.604599f
C14 VP B 7.082941f
C15 VDD2.t1 B 0.014546f
C16 VDD2.t0 B 0.014546f
C17 VDD2.n0 B 0.123103f
C18 VDD2.t3 B 0.014546f
C19 VDD2.t2 B 0.014546f
C20 VDD2.n1 B 0.035957f
C21 VDD2.n2 B 2.19156f
C22 VN.t2 B 0.256096f
C23 VN.t3 B 0.252701f
C24 VN.n0 B 0.170285f
C25 VN.t1 B 0.256096f
C26 VN.t0 B 0.252701f
C27 VN.n1 B 1.21264f
C28 VDD1.t0 B 0.013483f
C29 VDD1.t1 B 0.013483f
C30 VDD1.n0 B 0.03339f
C31 VDD1.t2 B 0.013483f
C32 VDD1.t3 B 0.013483f
C33 VDD1.n1 B 0.12116f
C34 VTAIL.t1 B 0.067436f
C35 VTAIL.n0 B 0.188348f
C36 VTAIL.t5 B 0.067436f
C37 VTAIL.n1 B 0.280241f
C38 VTAIL.t7 B 0.067436f
C39 VTAIL.n2 B 0.859888f
C40 VTAIL.t3 B 0.067436f
C41 VTAIL.n3 B 0.859888f
C42 VTAIL.t0 B 0.067436f
C43 VTAIL.n4 B 0.280241f
C44 VTAIL.t4 B 0.067436f
C45 VTAIL.n5 B 0.280241f
C46 VTAIL.t6 B 0.067436f
C47 VTAIL.n6 B 0.859888f
C48 VTAIL.t2 B 0.067436f
C49 VTAIL.n7 B 0.757678f
C50 VP.n0 B 0.038516f
C51 VP.t0 B 0.066348f
C52 VP.n1 B 0.023597f
C53 VP.n2 B 0.038516f
C54 VP.t1 B 0.066348f
C55 VP.t2 B 0.255432f
C56 VP.t3 B 0.258864f
C57 VP.n3 B 1.21028f
C58 VP.n4 B 1.16936f
C59 VP.n5 B 0.155923f
C60 VP.n6 B 0.041875f
C61 VP.n7 B 0.057761f
C62 VP.n8 B 0.029216f
C63 VP.n9 B 0.029216f
C64 VP.n10 B 0.029216f
C65 VP.n11 B 0.057761f
C66 VP.n12 B 0.041875f
C67 VP.n13 B 0.155923f
C68 VP.n14 B 0.041867f
.ends

