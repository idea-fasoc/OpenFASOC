* NGSPICE file created from diff_pair_sample_0881.ext - technology: sky130A

.subckt diff_pair_sample_0881 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0 ps=0 w=2.94 l=1.62
X1 VTAIL.t11 VP.t0 VDD1.t5 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=0.4851 ps=3.27 w=2.94 l=1.62
X2 B.t8 B.t6 B.t7 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0 ps=0 w=2.94 l=1.62
X3 B.t5 B.t3 B.t4 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0 ps=0 w=2.94 l=1.62
X4 B.t2 B.t0 B.t1 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0 ps=0 w=2.94 l=1.62
X5 VDD2.t5 VN.t0 VTAIL.t5 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=1.1466 ps=6.66 w=2.94 l=1.62
X6 VDD1.t0 VP.t1 VTAIL.t10 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0.4851 ps=3.27 w=2.94 l=1.62
X7 VDD2.t4 VN.t1 VTAIL.t1 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=1.1466 ps=6.66 w=2.94 l=1.62
X8 VTAIL.t3 VN.t2 VDD2.t3 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=0.4851 ps=3.27 w=2.94 l=1.62
X9 VDD2.t2 VN.t3 VTAIL.t4 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0.4851 ps=3.27 w=2.94 l=1.62
X10 VDD2.t1 VN.t4 VTAIL.t0 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0.4851 ps=3.27 w=2.94 l=1.62
X11 VDD1.t4 VP.t2 VTAIL.t9 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=1.1466 pd=6.66 as=0.4851 ps=3.27 w=2.94 l=1.62
X12 VDD1.t3 VP.t3 VTAIL.t8 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=1.1466 ps=6.66 w=2.94 l=1.62
X13 VTAIL.t7 VP.t4 VDD1.t2 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=0.4851 ps=3.27 w=2.94 l=1.62
X14 VDD1.t1 VP.t5 VTAIL.t6 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=1.1466 ps=6.66 w=2.94 l=1.62
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n2530_n1556# sky130_fd_pr__pfet_01v8 ad=0.4851 pd=3.27 as=0.4851 ps=3.27 w=2.94 l=1.62
R0 B.n312 B.n311 585
R1 B.n313 B.n40 585
R2 B.n315 B.n314 585
R3 B.n316 B.n39 585
R4 B.n318 B.n317 585
R5 B.n319 B.n38 585
R6 B.n321 B.n320 585
R7 B.n322 B.n37 585
R8 B.n324 B.n323 585
R9 B.n325 B.n36 585
R10 B.n327 B.n326 585
R11 B.n328 B.n35 585
R12 B.n330 B.n329 585
R13 B.n331 B.n34 585
R14 B.n333 B.n332 585
R15 B.n335 B.n31 585
R16 B.n337 B.n336 585
R17 B.n338 B.n30 585
R18 B.n340 B.n339 585
R19 B.n341 B.n29 585
R20 B.n343 B.n342 585
R21 B.n344 B.n28 585
R22 B.n346 B.n345 585
R23 B.n347 B.n25 585
R24 B.n350 B.n349 585
R25 B.n351 B.n24 585
R26 B.n353 B.n352 585
R27 B.n354 B.n23 585
R28 B.n356 B.n355 585
R29 B.n357 B.n22 585
R30 B.n359 B.n358 585
R31 B.n360 B.n21 585
R32 B.n362 B.n361 585
R33 B.n363 B.n20 585
R34 B.n365 B.n364 585
R35 B.n366 B.n19 585
R36 B.n368 B.n367 585
R37 B.n369 B.n18 585
R38 B.n371 B.n370 585
R39 B.n310 B.n41 585
R40 B.n309 B.n308 585
R41 B.n307 B.n42 585
R42 B.n306 B.n305 585
R43 B.n304 B.n43 585
R44 B.n303 B.n302 585
R45 B.n301 B.n44 585
R46 B.n300 B.n299 585
R47 B.n298 B.n45 585
R48 B.n297 B.n296 585
R49 B.n295 B.n46 585
R50 B.n294 B.n293 585
R51 B.n292 B.n47 585
R52 B.n291 B.n290 585
R53 B.n289 B.n48 585
R54 B.n288 B.n287 585
R55 B.n286 B.n49 585
R56 B.n285 B.n284 585
R57 B.n283 B.n50 585
R58 B.n282 B.n281 585
R59 B.n280 B.n51 585
R60 B.n279 B.n278 585
R61 B.n277 B.n52 585
R62 B.n276 B.n275 585
R63 B.n274 B.n53 585
R64 B.n273 B.n272 585
R65 B.n271 B.n54 585
R66 B.n270 B.n269 585
R67 B.n268 B.n55 585
R68 B.n267 B.n266 585
R69 B.n265 B.n56 585
R70 B.n264 B.n263 585
R71 B.n262 B.n57 585
R72 B.n261 B.n260 585
R73 B.n259 B.n58 585
R74 B.n258 B.n257 585
R75 B.n256 B.n59 585
R76 B.n255 B.n254 585
R77 B.n253 B.n60 585
R78 B.n252 B.n251 585
R79 B.n250 B.n61 585
R80 B.n249 B.n248 585
R81 B.n247 B.n62 585
R82 B.n246 B.n245 585
R83 B.n244 B.n63 585
R84 B.n243 B.n242 585
R85 B.n241 B.n64 585
R86 B.n240 B.n239 585
R87 B.n238 B.n65 585
R88 B.n237 B.n236 585
R89 B.n235 B.n66 585
R90 B.n234 B.n233 585
R91 B.n232 B.n67 585
R92 B.n231 B.n230 585
R93 B.n229 B.n68 585
R94 B.n228 B.n227 585
R95 B.n226 B.n69 585
R96 B.n225 B.n224 585
R97 B.n223 B.n70 585
R98 B.n222 B.n221 585
R99 B.n220 B.n71 585
R100 B.n219 B.n218 585
R101 B.n217 B.n72 585
R102 B.n157 B.n96 585
R103 B.n159 B.n158 585
R104 B.n160 B.n95 585
R105 B.n162 B.n161 585
R106 B.n163 B.n94 585
R107 B.n165 B.n164 585
R108 B.n166 B.n93 585
R109 B.n168 B.n167 585
R110 B.n169 B.n92 585
R111 B.n171 B.n170 585
R112 B.n172 B.n91 585
R113 B.n174 B.n173 585
R114 B.n175 B.n90 585
R115 B.n177 B.n176 585
R116 B.n178 B.n87 585
R117 B.n181 B.n180 585
R118 B.n182 B.n86 585
R119 B.n184 B.n183 585
R120 B.n185 B.n85 585
R121 B.n187 B.n186 585
R122 B.n188 B.n84 585
R123 B.n190 B.n189 585
R124 B.n191 B.n83 585
R125 B.n193 B.n192 585
R126 B.n195 B.n194 585
R127 B.n196 B.n79 585
R128 B.n198 B.n197 585
R129 B.n199 B.n78 585
R130 B.n201 B.n200 585
R131 B.n202 B.n77 585
R132 B.n204 B.n203 585
R133 B.n205 B.n76 585
R134 B.n207 B.n206 585
R135 B.n208 B.n75 585
R136 B.n210 B.n209 585
R137 B.n211 B.n74 585
R138 B.n213 B.n212 585
R139 B.n214 B.n73 585
R140 B.n216 B.n215 585
R141 B.n156 B.n155 585
R142 B.n154 B.n97 585
R143 B.n153 B.n152 585
R144 B.n151 B.n98 585
R145 B.n150 B.n149 585
R146 B.n148 B.n99 585
R147 B.n147 B.n146 585
R148 B.n145 B.n100 585
R149 B.n144 B.n143 585
R150 B.n142 B.n101 585
R151 B.n141 B.n140 585
R152 B.n139 B.n102 585
R153 B.n138 B.n137 585
R154 B.n136 B.n103 585
R155 B.n135 B.n134 585
R156 B.n133 B.n104 585
R157 B.n132 B.n131 585
R158 B.n130 B.n105 585
R159 B.n129 B.n128 585
R160 B.n127 B.n106 585
R161 B.n126 B.n125 585
R162 B.n124 B.n107 585
R163 B.n123 B.n122 585
R164 B.n121 B.n108 585
R165 B.n120 B.n119 585
R166 B.n118 B.n109 585
R167 B.n117 B.n116 585
R168 B.n115 B.n110 585
R169 B.n114 B.n113 585
R170 B.n112 B.n111 585
R171 B.n2 B.n0 585
R172 B.n417 B.n1 585
R173 B.n416 B.n415 585
R174 B.n414 B.n3 585
R175 B.n413 B.n412 585
R176 B.n411 B.n4 585
R177 B.n410 B.n409 585
R178 B.n408 B.n5 585
R179 B.n407 B.n406 585
R180 B.n405 B.n6 585
R181 B.n404 B.n403 585
R182 B.n402 B.n7 585
R183 B.n401 B.n400 585
R184 B.n399 B.n8 585
R185 B.n398 B.n397 585
R186 B.n396 B.n9 585
R187 B.n395 B.n394 585
R188 B.n393 B.n10 585
R189 B.n392 B.n391 585
R190 B.n390 B.n11 585
R191 B.n389 B.n388 585
R192 B.n387 B.n12 585
R193 B.n386 B.n385 585
R194 B.n384 B.n13 585
R195 B.n383 B.n382 585
R196 B.n381 B.n14 585
R197 B.n380 B.n379 585
R198 B.n378 B.n15 585
R199 B.n377 B.n376 585
R200 B.n375 B.n16 585
R201 B.n374 B.n373 585
R202 B.n372 B.n17 585
R203 B.n419 B.n418 585
R204 B.n157 B.n156 550.159
R205 B.n370 B.n17 550.159
R206 B.n217 B.n216 550.159
R207 B.n312 B.n41 550.159
R208 B.n80 B.t6 249.597
R209 B.n88 B.t3 249.597
R210 B.n26 B.t0 249.597
R211 B.n32 B.t9 249.597
R212 B.n80 B.t8 182.099
R213 B.n32 B.t10 182.099
R214 B.n88 B.t5 182.096
R215 B.n26 B.t1 182.096
R216 B.n156 B.n97 163.367
R217 B.n152 B.n97 163.367
R218 B.n152 B.n151 163.367
R219 B.n151 B.n150 163.367
R220 B.n150 B.n99 163.367
R221 B.n146 B.n99 163.367
R222 B.n146 B.n145 163.367
R223 B.n145 B.n144 163.367
R224 B.n144 B.n101 163.367
R225 B.n140 B.n101 163.367
R226 B.n140 B.n139 163.367
R227 B.n139 B.n138 163.367
R228 B.n138 B.n103 163.367
R229 B.n134 B.n103 163.367
R230 B.n134 B.n133 163.367
R231 B.n133 B.n132 163.367
R232 B.n132 B.n105 163.367
R233 B.n128 B.n105 163.367
R234 B.n128 B.n127 163.367
R235 B.n127 B.n126 163.367
R236 B.n126 B.n107 163.367
R237 B.n122 B.n107 163.367
R238 B.n122 B.n121 163.367
R239 B.n121 B.n120 163.367
R240 B.n120 B.n109 163.367
R241 B.n116 B.n109 163.367
R242 B.n116 B.n115 163.367
R243 B.n115 B.n114 163.367
R244 B.n114 B.n111 163.367
R245 B.n111 B.n2 163.367
R246 B.n418 B.n2 163.367
R247 B.n418 B.n417 163.367
R248 B.n417 B.n416 163.367
R249 B.n416 B.n3 163.367
R250 B.n412 B.n3 163.367
R251 B.n412 B.n411 163.367
R252 B.n411 B.n410 163.367
R253 B.n410 B.n5 163.367
R254 B.n406 B.n5 163.367
R255 B.n406 B.n405 163.367
R256 B.n405 B.n404 163.367
R257 B.n404 B.n7 163.367
R258 B.n400 B.n7 163.367
R259 B.n400 B.n399 163.367
R260 B.n399 B.n398 163.367
R261 B.n398 B.n9 163.367
R262 B.n394 B.n9 163.367
R263 B.n394 B.n393 163.367
R264 B.n393 B.n392 163.367
R265 B.n392 B.n11 163.367
R266 B.n388 B.n11 163.367
R267 B.n388 B.n387 163.367
R268 B.n387 B.n386 163.367
R269 B.n386 B.n13 163.367
R270 B.n382 B.n13 163.367
R271 B.n382 B.n381 163.367
R272 B.n381 B.n380 163.367
R273 B.n380 B.n15 163.367
R274 B.n376 B.n15 163.367
R275 B.n376 B.n375 163.367
R276 B.n375 B.n374 163.367
R277 B.n374 B.n17 163.367
R278 B.n158 B.n157 163.367
R279 B.n158 B.n95 163.367
R280 B.n162 B.n95 163.367
R281 B.n163 B.n162 163.367
R282 B.n164 B.n163 163.367
R283 B.n164 B.n93 163.367
R284 B.n168 B.n93 163.367
R285 B.n169 B.n168 163.367
R286 B.n170 B.n169 163.367
R287 B.n170 B.n91 163.367
R288 B.n174 B.n91 163.367
R289 B.n175 B.n174 163.367
R290 B.n176 B.n175 163.367
R291 B.n176 B.n87 163.367
R292 B.n181 B.n87 163.367
R293 B.n182 B.n181 163.367
R294 B.n183 B.n182 163.367
R295 B.n183 B.n85 163.367
R296 B.n187 B.n85 163.367
R297 B.n188 B.n187 163.367
R298 B.n189 B.n188 163.367
R299 B.n189 B.n83 163.367
R300 B.n193 B.n83 163.367
R301 B.n194 B.n193 163.367
R302 B.n194 B.n79 163.367
R303 B.n198 B.n79 163.367
R304 B.n199 B.n198 163.367
R305 B.n200 B.n199 163.367
R306 B.n200 B.n77 163.367
R307 B.n204 B.n77 163.367
R308 B.n205 B.n204 163.367
R309 B.n206 B.n205 163.367
R310 B.n206 B.n75 163.367
R311 B.n210 B.n75 163.367
R312 B.n211 B.n210 163.367
R313 B.n212 B.n211 163.367
R314 B.n212 B.n73 163.367
R315 B.n216 B.n73 163.367
R316 B.n218 B.n217 163.367
R317 B.n218 B.n71 163.367
R318 B.n222 B.n71 163.367
R319 B.n223 B.n222 163.367
R320 B.n224 B.n223 163.367
R321 B.n224 B.n69 163.367
R322 B.n228 B.n69 163.367
R323 B.n229 B.n228 163.367
R324 B.n230 B.n229 163.367
R325 B.n230 B.n67 163.367
R326 B.n234 B.n67 163.367
R327 B.n235 B.n234 163.367
R328 B.n236 B.n235 163.367
R329 B.n236 B.n65 163.367
R330 B.n240 B.n65 163.367
R331 B.n241 B.n240 163.367
R332 B.n242 B.n241 163.367
R333 B.n242 B.n63 163.367
R334 B.n246 B.n63 163.367
R335 B.n247 B.n246 163.367
R336 B.n248 B.n247 163.367
R337 B.n248 B.n61 163.367
R338 B.n252 B.n61 163.367
R339 B.n253 B.n252 163.367
R340 B.n254 B.n253 163.367
R341 B.n254 B.n59 163.367
R342 B.n258 B.n59 163.367
R343 B.n259 B.n258 163.367
R344 B.n260 B.n259 163.367
R345 B.n260 B.n57 163.367
R346 B.n264 B.n57 163.367
R347 B.n265 B.n264 163.367
R348 B.n266 B.n265 163.367
R349 B.n266 B.n55 163.367
R350 B.n270 B.n55 163.367
R351 B.n271 B.n270 163.367
R352 B.n272 B.n271 163.367
R353 B.n272 B.n53 163.367
R354 B.n276 B.n53 163.367
R355 B.n277 B.n276 163.367
R356 B.n278 B.n277 163.367
R357 B.n278 B.n51 163.367
R358 B.n282 B.n51 163.367
R359 B.n283 B.n282 163.367
R360 B.n284 B.n283 163.367
R361 B.n284 B.n49 163.367
R362 B.n288 B.n49 163.367
R363 B.n289 B.n288 163.367
R364 B.n290 B.n289 163.367
R365 B.n290 B.n47 163.367
R366 B.n294 B.n47 163.367
R367 B.n295 B.n294 163.367
R368 B.n296 B.n295 163.367
R369 B.n296 B.n45 163.367
R370 B.n300 B.n45 163.367
R371 B.n301 B.n300 163.367
R372 B.n302 B.n301 163.367
R373 B.n302 B.n43 163.367
R374 B.n306 B.n43 163.367
R375 B.n307 B.n306 163.367
R376 B.n308 B.n307 163.367
R377 B.n308 B.n41 163.367
R378 B.n370 B.n369 163.367
R379 B.n369 B.n368 163.367
R380 B.n368 B.n19 163.367
R381 B.n364 B.n19 163.367
R382 B.n364 B.n363 163.367
R383 B.n363 B.n362 163.367
R384 B.n362 B.n21 163.367
R385 B.n358 B.n21 163.367
R386 B.n358 B.n357 163.367
R387 B.n357 B.n356 163.367
R388 B.n356 B.n23 163.367
R389 B.n352 B.n23 163.367
R390 B.n352 B.n351 163.367
R391 B.n351 B.n350 163.367
R392 B.n350 B.n25 163.367
R393 B.n345 B.n25 163.367
R394 B.n345 B.n344 163.367
R395 B.n344 B.n343 163.367
R396 B.n343 B.n29 163.367
R397 B.n339 B.n29 163.367
R398 B.n339 B.n338 163.367
R399 B.n338 B.n337 163.367
R400 B.n337 B.n31 163.367
R401 B.n332 B.n31 163.367
R402 B.n332 B.n331 163.367
R403 B.n331 B.n330 163.367
R404 B.n330 B.n35 163.367
R405 B.n326 B.n35 163.367
R406 B.n326 B.n325 163.367
R407 B.n325 B.n324 163.367
R408 B.n324 B.n37 163.367
R409 B.n320 B.n37 163.367
R410 B.n320 B.n319 163.367
R411 B.n319 B.n318 163.367
R412 B.n318 B.n39 163.367
R413 B.n314 B.n39 163.367
R414 B.n314 B.n313 163.367
R415 B.n313 B.n312 163.367
R416 B.n81 B.t7 144.28
R417 B.n33 B.t11 144.28
R418 B.n89 B.t4 144.279
R419 B.n27 B.t2 144.279
R420 B.n82 B.n81 59.5399
R421 B.n179 B.n89 59.5399
R422 B.n348 B.n27 59.5399
R423 B.n334 B.n33 59.5399
R424 B.n81 B.n80 37.8187
R425 B.n89 B.n88 37.8187
R426 B.n27 B.n26 37.8187
R427 B.n33 B.n32 37.8187
R428 B.n372 B.n371 35.7468
R429 B.n311 B.n310 35.7468
R430 B.n215 B.n72 35.7468
R431 B.n155 B.n96 35.7468
R432 B B.n419 18.0485
R433 B.n371 B.n18 10.6151
R434 B.n367 B.n18 10.6151
R435 B.n367 B.n366 10.6151
R436 B.n366 B.n365 10.6151
R437 B.n365 B.n20 10.6151
R438 B.n361 B.n20 10.6151
R439 B.n361 B.n360 10.6151
R440 B.n360 B.n359 10.6151
R441 B.n359 B.n22 10.6151
R442 B.n355 B.n22 10.6151
R443 B.n355 B.n354 10.6151
R444 B.n354 B.n353 10.6151
R445 B.n353 B.n24 10.6151
R446 B.n349 B.n24 10.6151
R447 B.n347 B.n346 10.6151
R448 B.n346 B.n28 10.6151
R449 B.n342 B.n28 10.6151
R450 B.n342 B.n341 10.6151
R451 B.n341 B.n340 10.6151
R452 B.n340 B.n30 10.6151
R453 B.n336 B.n30 10.6151
R454 B.n336 B.n335 10.6151
R455 B.n333 B.n34 10.6151
R456 B.n329 B.n34 10.6151
R457 B.n329 B.n328 10.6151
R458 B.n328 B.n327 10.6151
R459 B.n327 B.n36 10.6151
R460 B.n323 B.n36 10.6151
R461 B.n323 B.n322 10.6151
R462 B.n322 B.n321 10.6151
R463 B.n321 B.n38 10.6151
R464 B.n317 B.n38 10.6151
R465 B.n317 B.n316 10.6151
R466 B.n316 B.n315 10.6151
R467 B.n315 B.n40 10.6151
R468 B.n311 B.n40 10.6151
R469 B.n219 B.n72 10.6151
R470 B.n220 B.n219 10.6151
R471 B.n221 B.n220 10.6151
R472 B.n221 B.n70 10.6151
R473 B.n225 B.n70 10.6151
R474 B.n226 B.n225 10.6151
R475 B.n227 B.n226 10.6151
R476 B.n227 B.n68 10.6151
R477 B.n231 B.n68 10.6151
R478 B.n232 B.n231 10.6151
R479 B.n233 B.n232 10.6151
R480 B.n233 B.n66 10.6151
R481 B.n237 B.n66 10.6151
R482 B.n238 B.n237 10.6151
R483 B.n239 B.n238 10.6151
R484 B.n239 B.n64 10.6151
R485 B.n243 B.n64 10.6151
R486 B.n244 B.n243 10.6151
R487 B.n245 B.n244 10.6151
R488 B.n245 B.n62 10.6151
R489 B.n249 B.n62 10.6151
R490 B.n250 B.n249 10.6151
R491 B.n251 B.n250 10.6151
R492 B.n251 B.n60 10.6151
R493 B.n255 B.n60 10.6151
R494 B.n256 B.n255 10.6151
R495 B.n257 B.n256 10.6151
R496 B.n257 B.n58 10.6151
R497 B.n261 B.n58 10.6151
R498 B.n262 B.n261 10.6151
R499 B.n263 B.n262 10.6151
R500 B.n263 B.n56 10.6151
R501 B.n267 B.n56 10.6151
R502 B.n268 B.n267 10.6151
R503 B.n269 B.n268 10.6151
R504 B.n269 B.n54 10.6151
R505 B.n273 B.n54 10.6151
R506 B.n274 B.n273 10.6151
R507 B.n275 B.n274 10.6151
R508 B.n275 B.n52 10.6151
R509 B.n279 B.n52 10.6151
R510 B.n280 B.n279 10.6151
R511 B.n281 B.n280 10.6151
R512 B.n281 B.n50 10.6151
R513 B.n285 B.n50 10.6151
R514 B.n286 B.n285 10.6151
R515 B.n287 B.n286 10.6151
R516 B.n287 B.n48 10.6151
R517 B.n291 B.n48 10.6151
R518 B.n292 B.n291 10.6151
R519 B.n293 B.n292 10.6151
R520 B.n293 B.n46 10.6151
R521 B.n297 B.n46 10.6151
R522 B.n298 B.n297 10.6151
R523 B.n299 B.n298 10.6151
R524 B.n299 B.n44 10.6151
R525 B.n303 B.n44 10.6151
R526 B.n304 B.n303 10.6151
R527 B.n305 B.n304 10.6151
R528 B.n305 B.n42 10.6151
R529 B.n309 B.n42 10.6151
R530 B.n310 B.n309 10.6151
R531 B.n159 B.n96 10.6151
R532 B.n160 B.n159 10.6151
R533 B.n161 B.n160 10.6151
R534 B.n161 B.n94 10.6151
R535 B.n165 B.n94 10.6151
R536 B.n166 B.n165 10.6151
R537 B.n167 B.n166 10.6151
R538 B.n167 B.n92 10.6151
R539 B.n171 B.n92 10.6151
R540 B.n172 B.n171 10.6151
R541 B.n173 B.n172 10.6151
R542 B.n173 B.n90 10.6151
R543 B.n177 B.n90 10.6151
R544 B.n178 B.n177 10.6151
R545 B.n180 B.n86 10.6151
R546 B.n184 B.n86 10.6151
R547 B.n185 B.n184 10.6151
R548 B.n186 B.n185 10.6151
R549 B.n186 B.n84 10.6151
R550 B.n190 B.n84 10.6151
R551 B.n191 B.n190 10.6151
R552 B.n192 B.n191 10.6151
R553 B.n196 B.n195 10.6151
R554 B.n197 B.n196 10.6151
R555 B.n197 B.n78 10.6151
R556 B.n201 B.n78 10.6151
R557 B.n202 B.n201 10.6151
R558 B.n203 B.n202 10.6151
R559 B.n203 B.n76 10.6151
R560 B.n207 B.n76 10.6151
R561 B.n208 B.n207 10.6151
R562 B.n209 B.n208 10.6151
R563 B.n209 B.n74 10.6151
R564 B.n213 B.n74 10.6151
R565 B.n214 B.n213 10.6151
R566 B.n215 B.n214 10.6151
R567 B.n155 B.n154 10.6151
R568 B.n154 B.n153 10.6151
R569 B.n153 B.n98 10.6151
R570 B.n149 B.n98 10.6151
R571 B.n149 B.n148 10.6151
R572 B.n148 B.n147 10.6151
R573 B.n147 B.n100 10.6151
R574 B.n143 B.n100 10.6151
R575 B.n143 B.n142 10.6151
R576 B.n142 B.n141 10.6151
R577 B.n141 B.n102 10.6151
R578 B.n137 B.n102 10.6151
R579 B.n137 B.n136 10.6151
R580 B.n136 B.n135 10.6151
R581 B.n135 B.n104 10.6151
R582 B.n131 B.n104 10.6151
R583 B.n131 B.n130 10.6151
R584 B.n130 B.n129 10.6151
R585 B.n129 B.n106 10.6151
R586 B.n125 B.n106 10.6151
R587 B.n125 B.n124 10.6151
R588 B.n124 B.n123 10.6151
R589 B.n123 B.n108 10.6151
R590 B.n119 B.n108 10.6151
R591 B.n119 B.n118 10.6151
R592 B.n118 B.n117 10.6151
R593 B.n117 B.n110 10.6151
R594 B.n113 B.n110 10.6151
R595 B.n113 B.n112 10.6151
R596 B.n112 B.n0 10.6151
R597 B.n415 B.n1 10.6151
R598 B.n415 B.n414 10.6151
R599 B.n414 B.n413 10.6151
R600 B.n413 B.n4 10.6151
R601 B.n409 B.n4 10.6151
R602 B.n409 B.n408 10.6151
R603 B.n408 B.n407 10.6151
R604 B.n407 B.n6 10.6151
R605 B.n403 B.n6 10.6151
R606 B.n403 B.n402 10.6151
R607 B.n402 B.n401 10.6151
R608 B.n401 B.n8 10.6151
R609 B.n397 B.n8 10.6151
R610 B.n397 B.n396 10.6151
R611 B.n396 B.n395 10.6151
R612 B.n395 B.n10 10.6151
R613 B.n391 B.n10 10.6151
R614 B.n391 B.n390 10.6151
R615 B.n390 B.n389 10.6151
R616 B.n389 B.n12 10.6151
R617 B.n385 B.n12 10.6151
R618 B.n385 B.n384 10.6151
R619 B.n384 B.n383 10.6151
R620 B.n383 B.n14 10.6151
R621 B.n379 B.n14 10.6151
R622 B.n379 B.n378 10.6151
R623 B.n378 B.n377 10.6151
R624 B.n377 B.n16 10.6151
R625 B.n373 B.n16 10.6151
R626 B.n373 B.n372 10.6151
R627 B.n348 B.n347 6.5566
R628 B.n335 B.n334 6.5566
R629 B.n180 B.n179 6.5566
R630 B.n192 B.n82 6.5566
R631 B.n349 B.n348 4.05904
R632 B.n334 B.n333 4.05904
R633 B.n179 B.n178 4.05904
R634 B.n195 B.n82 4.05904
R635 B.n419 B.n0 2.81026
R636 B.n419 B.n1 2.81026
R637 VP.n17 VP.n16 176.055
R638 VP.n32 VP.n31 176.055
R639 VP.n15 VP.n14 176.055
R640 VP.n9 VP.n8 161.3
R641 VP.n10 VP.n5 161.3
R642 VP.n12 VP.n11 161.3
R643 VP.n13 VP.n4 161.3
R644 VP.n30 VP.n0 161.3
R645 VP.n29 VP.n28 161.3
R646 VP.n27 VP.n1 161.3
R647 VP.n26 VP.n25 161.3
R648 VP.n23 VP.n2 161.3
R649 VP.n22 VP.n21 161.3
R650 VP.n20 VP.n3 161.3
R651 VP.n19 VP.n18 161.3
R652 VP.n6 VP.t2 77.4414
R653 VP.n22 VP.n3 56.5617
R654 VP.n29 VP.n1 56.5617
R655 VP.n12 VP.n5 56.5617
R656 VP.n7 VP.n6 54.2669
R657 VP.n17 VP.t1 43.7375
R658 VP.n24 VP.t0 43.7375
R659 VP.n31 VP.t5 43.7375
R660 VP.n14 VP.t3 43.7375
R661 VP.n7 VP.t4 43.7375
R662 VP.n16 VP.n15 37.921
R663 VP.n18 VP.n3 24.5923
R664 VP.n23 VP.n22 24.5923
R665 VP.n25 VP.n1 24.5923
R666 VP.n30 VP.n29 24.5923
R667 VP.n13 VP.n12 24.5923
R668 VP.n8 VP.n5 24.5923
R669 VP.n9 VP.n6 17.7808
R670 VP.n24 VP.n23 12.2964
R671 VP.n25 VP.n24 12.2964
R672 VP.n8 VP.n7 12.2964
R673 VP.n18 VP.n17 9.83723
R674 VP.n31 VP.n30 9.83723
R675 VP.n14 VP.n13 9.83723
R676 VP.n10 VP.n9 0.189894
R677 VP.n11 VP.n10 0.189894
R678 VP.n11 VP.n4 0.189894
R679 VP.n15 VP.n4 0.189894
R680 VP.n19 VP.n16 0.189894
R681 VP.n20 VP.n19 0.189894
R682 VP.n21 VP.n20 0.189894
R683 VP.n21 VP.n2 0.189894
R684 VP.n26 VP.n2 0.189894
R685 VP.n27 VP.n26 0.189894
R686 VP.n28 VP.n27 0.189894
R687 VP.n28 VP.n0 0.189894
R688 VP.n32 VP.n0 0.189894
R689 VP VP.n32 0.0516364
R690 VDD1 VDD1.t4 153.936
R691 VDD1.n1 VDD1.t0 153.822
R692 VDD1.n1 VDD1.n0 141.925
R693 VDD1.n3 VDD1.n2 141.561
R694 VDD1.n3 VDD1.n1 33.1367
R695 VDD1.n2 VDD1.t2 11.0566
R696 VDD1.n2 VDD1.t3 11.0566
R697 VDD1.n0 VDD1.t5 11.0566
R698 VDD1.n0 VDD1.t1 11.0566
R699 VDD1 VDD1.n3 0.362569
R700 VTAIL.n7 VTAIL.t1 135.939
R701 VTAIL.n11 VTAIL.t5 135.939
R702 VTAIL.n2 VTAIL.t6 135.939
R703 VTAIL.n10 VTAIL.t8 135.939
R704 VTAIL.n9 VTAIL.n8 124.882
R705 VTAIL.n6 VTAIL.n5 124.882
R706 VTAIL.n1 VTAIL.n0 124.882
R707 VTAIL.n4 VTAIL.n3 124.882
R708 VTAIL.n6 VTAIL.n4 18.2634
R709 VTAIL.n11 VTAIL.n10 16.5824
R710 VTAIL.n0 VTAIL.t0 11.0566
R711 VTAIL.n0 VTAIL.t2 11.0566
R712 VTAIL.n3 VTAIL.t10 11.0566
R713 VTAIL.n3 VTAIL.t11 11.0566
R714 VTAIL.n8 VTAIL.t9 11.0566
R715 VTAIL.n8 VTAIL.t7 11.0566
R716 VTAIL.n5 VTAIL.t4 11.0566
R717 VTAIL.n5 VTAIL.t3 11.0566
R718 VTAIL.n7 VTAIL.n6 1.68153
R719 VTAIL.n10 VTAIL.n9 1.68153
R720 VTAIL.n4 VTAIL.n2 1.68153
R721 VTAIL.n9 VTAIL.n7 1.31084
R722 VTAIL.n2 VTAIL.n1 1.31084
R723 VTAIL VTAIL.n11 1.20309
R724 VTAIL VTAIL.n1 0.478948
R725 VN.n11 VN.n10 176.055
R726 VN.n23 VN.n22 176.055
R727 VN.n21 VN.n12 161.3
R728 VN.n20 VN.n19 161.3
R729 VN.n18 VN.n13 161.3
R730 VN.n17 VN.n16 161.3
R731 VN.n9 VN.n0 161.3
R732 VN.n8 VN.n7 161.3
R733 VN.n6 VN.n1 161.3
R734 VN.n5 VN.n4 161.3
R735 VN.n2 VN.t4 77.4414
R736 VN.n14 VN.t1 77.4414
R737 VN.n8 VN.n1 56.5617
R738 VN.n20 VN.n13 56.5617
R739 VN.n3 VN.n2 54.2669
R740 VN.n15 VN.n14 54.2669
R741 VN.n3 VN.t5 43.7375
R742 VN.n10 VN.t0 43.7375
R743 VN.n15 VN.t2 43.7375
R744 VN.n22 VN.t3 43.7375
R745 VN VN.n23 38.3016
R746 VN.n4 VN.n1 24.5923
R747 VN.n9 VN.n8 24.5923
R748 VN.n16 VN.n13 24.5923
R749 VN.n21 VN.n20 24.5923
R750 VN.n17 VN.n14 17.7808
R751 VN.n5 VN.n2 17.7808
R752 VN.n4 VN.n3 12.2964
R753 VN.n16 VN.n15 12.2964
R754 VN.n10 VN.n9 9.83723
R755 VN.n22 VN.n21 9.83723
R756 VN.n23 VN.n12 0.189894
R757 VN.n19 VN.n12 0.189894
R758 VN.n19 VN.n18 0.189894
R759 VN.n18 VN.n17 0.189894
R760 VN.n6 VN.n5 0.189894
R761 VN.n7 VN.n6 0.189894
R762 VN.n7 VN.n0 0.189894
R763 VN.n11 VN.n0 0.189894
R764 VN VN.n11 0.0516364
R765 VDD2.n1 VDD2.t1 153.822
R766 VDD2.n2 VDD2.t2 152.618
R767 VDD2.n1 VDD2.n0 141.925
R768 VDD2 VDD2.n3 141.923
R769 VDD2.n2 VDD2.n1 31.7131
R770 VDD2.n3 VDD2.t3 11.0566
R771 VDD2.n3 VDD2.t4 11.0566
R772 VDD2.n0 VDD2.t0 11.0566
R773 VDD2.n0 VDD2.t5 11.0566
R774 VDD2 VDD2.n2 1.31947
C0 VP w_n2530_n1556# 4.68592f
C1 VTAIL w_n2530_n1556# 1.56335f
C2 VN B 0.855224f
C3 VTAIL VP 2.20835f
C4 VDD1 w_n2530_n1556# 1.4036f
C5 VDD1 VP 1.97139f
C6 VDD2 B 1.18413f
C7 VDD1 VTAIL 3.89146f
C8 VDD2 VN 1.74797f
C9 B w_n2530_n1556# 5.79368f
C10 VP B 1.3914f
C11 VN w_n2530_n1556# 4.36399f
C12 VTAIL B 1.345f
C13 VN VP 4.29722f
C14 VDD1 B 1.1333f
C15 VTAIL VN 2.19417f
C16 VDD2 w_n2530_n1556# 1.4567f
C17 VDD1 VN 0.15501f
C18 VDD2 VP 0.380578f
C19 VDD2 VTAIL 3.93744f
C20 VDD2 VDD1 1.05135f
C21 VDD2 VSUBS 0.870396f
C22 VDD1 VSUBS 1.221074f
C23 VTAIL VSUBS 0.449419f
C24 VN VSUBS 4.3703f
C25 VP VSUBS 1.675282f
C26 B VSUBS 2.747009f
C27 w_n2530_n1556# VSUBS 49.8815f
C28 VDD2.t1 VSUBS 0.267467f
C29 VDD2.t0 VSUBS 0.035744f
C30 VDD2.t5 VSUBS 0.035744f
C31 VDD2.n0 VSUBS 0.186512f
C32 VDD2.n1 VSUBS 1.31217f
C33 VDD2.t2 VSUBS 0.265291f
C34 VDD2.n2 VSUBS 1.1555f
C35 VDD2.t3 VSUBS 0.035744f
C36 VDD2.t4 VSUBS 0.035744f
C37 VDD2.n3 VSUBS 0.186503f
C38 VN.n0 VSUBS 0.048322f
C39 VN.t0 VSUBS 0.571858f
C40 VN.n1 VSUBS 0.066901f
C41 VN.t4 VSUBS 0.771323f
C42 VN.n2 VSUBS 0.349833f
C43 VN.t5 VSUBS 0.571858f
C44 VN.n3 VSUBS 0.353566f
C45 VN.n4 VSUBS 0.06749f
C46 VN.n5 VSUBS 0.309992f
C47 VN.n6 VSUBS 0.048322f
C48 VN.n7 VSUBS 0.048322f
C49 VN.n8 VSUBS 0.073586f
C50 VN.n9 VSUBS 0.063066f
C51 VN.n10 VSUBS 0.367271f
C52 VN.n11 VSUBS 0.047331f
C53 VN.n12 VSUBS 0.048322f
C54 VN.t3 VSUBS 0.571858f
C55 VN.n13 VSUBS 0.066901f
C56 VN.t1 VSUBS 0.771323f
C57 VN.n14 VSUBS 0.349833f
C58 VN.t2 VSUBS 0.571858f
C59 VN.n15 VSUBS 0.353566f
C60 VN.n16 VSUBS 0.06749f
C61 VN.n17 VSUBS 0.309992f
C62 VN.n18 VSUBS 0.048322f
C63 VN.n19 VSUBS 0.048322f
C64 VN.n20 VSUBS 0.073586f
C65 VN.n21 VSUBS 0.063066f
C66 VN.n22 VSUBS 0.367271f
C67 VN.n23 VSUBS 1.71329f
C68 VTAIL.t0 VSUBS 0.069134f
C69 VTAIL.t2 VSUBS 0.069134f
C70 VTAIL.n0 VSUBS 0.310001f
C71 VTAIL.n1 VSUBS 0.554604f
C72 VTAIL.t6 VSUBS 0.463622f
C73 VTAIL.n2 VSUBS 0.704837f
C74 VTAIL.t10 VSUBS 0.069134f
C75 VTAIL.t11 VSUBS 0.069134f
C76 VTAIL.n3 VSUBS 0.310001f
C77 VTAIL.n4 VSUBS 1.51387f
C78 VTAIL.t4 VSUBS 0.069134f
C79 VTAIL.t3 VSUBS 0.069134f
C80 VTAIL.n5 VSUBS 0.310002f
C81 VTAIL.n6 VSUBS 1.51386f
C82 VTAIL.t1 VSUBS 0.463623f
C83 VTAIL.n7 VSUBS 0.704836f
C84 VTAIL.t9 VSUBS 0.069134f
C85 VTAIL.t7 VSUBS 0.069134f
C86 VTAIL.n8 VSUBS 0.310002f
C87 VTAIL.n9 VSUBS 0.66991f
C88 VTAIL.t8 VSUBS 0.463622f
C89 VTAIL.n10 VSUBS 1.38761f
C90 VTAIL.t5 VSUBS 0.463622f
C91 VTAIL.n11 VSUBS 1.34173f
C92 VDD1.t4 VSUBS 0.263872f
C93 VDD1.t0 VSUBS 0.263626f
C94 VDD1.t5 VSUBS 0.035231f
C95 VDD1.t1 VSUBS 0.035231f
C96 VDD1.n0 VSUBS 0.183833f
C97 VDD1.n1 VSUBS 1.3491f
C98 VDD1.t2 VSUBS 0.035231f
C99 VDD1.t3 VSUBS 0.035231f
C100 VDD1.n2 VSUBS 0.183067f
C101 VDD1.n3 VSUBS 1.15686f
C102 VP.n0 VSUBS 0.049964f
C103 VP.t5 VSUBS 0.591282f
C104 VP.n1 VSUBS 0.069174f
C105 VP.n2 VSUBS 0.049964f
C106 VP.t0 VSUBS 0.591282f
C107 VP.n3 VSUBS 0.076086f
C108 VP.n4 VSUBS 0.049964f
C109 VP.t3 VSUBS 0.591282f
C110 VP.n5 VSUBS 0.069174f
C111 VP.t2 VSUBS 0.797523f
C112 VP.n6 VSUBS 0.361715f
C113 VP.t4 VSUBS 0.591282f
C114 VP.n7 VSUBS 0.365576f
C115 VP.n8 VSUBS 0.069783f
C116 VP.n9 VSUBS 0.320521f
C117 VP.n10 VSUBS 0.049964f
C118 VP.n11 VSUBS 0.049964f
C119 VP.n12 VSUBS 0.076086f
C120 VP.n13 VSUBS 0.065209f
C121 VP.n14 VSUBS 0.379746f
C122 VP.n15 VSUBS 1.73847f
C123 VP.n16 VSUBS 1.78596f
C124 VP.t1 VSUBS 0.591282f
C125 VP.n17 VSUBS 0.379746f
C126 VP.n18 VSUBS 0.065209f
C127 VP.n19 VSUBS 0.049964f
C128 VP.n20 VSUBS 0.049964f
C129 VP.n21 VSUBS 0.049964f
C130 VP.n22 VSUBS 0.069174f
C131 VP.n23 VSUBS 0.069783f
C132 VP.n24 VSUBS 0.268038f
C133 VP.n25 VSUBS 0.069783f
C134 VP.n26 VSUBS 0.049964f
C135 VP.n27 VSUBS 0.049964f
C136 VP.n28 VSUBS 0.049964f
C137 VP.n29 VSUBS 0.076086f
C138 VP.n30 VSUBS 0.065209f
C139 VP.n31 VSUBS 0.379746f
C140 VP.n32 VSUBS 0.048938f
C141 B.n0 VSUBS 0.004996f
C142 B.n1 VSUBS 0.004996f
C143 B.n2 VSUBS 0.007901f
C144 B.n3 VSUBS 0.007901f
C145 B.n4 VSUBS 0.007901f
C146 B.n5 VSUBS 0.007901f
C147 B.n6 VSUBS 0.007901f
C148 B.n7 VSUBS 0.007901f
C149 B.n8 VSUBS 0.007901f
C150 B.n9 VSUBS 0.007901f
C151 B.n10 VSUBS 0.007901f
C152 B.n11 VSUBS 0.007901f
C153 B.n12 VSUBS 0.007901f
C154 B.n13 VSUBS 0.007901f
C155 B.n14 VSUBS 0.007901f
C156 B.n15 VSUBS 0.007901f
C157 B.n16 VSUBS 0.007901f
C158 B.n17 VSUBS 0.019375f
C159 B.n18 VSUBS 0.007901f
C160 B.n19 VSUBS 0.007901f
C161 B.n20 VSUBS 0.007901f
C162 B.n21 VSUBS 0.007901f
C163 B.n22 VSUBS 0.007901f
C164 B.n23 VSUBS 0.007901f
C165 B.n24 VSUBS 0.007901f
C166 B.n25 VSUBS 0.007901f
C167 B.t2 VSUBS 0.079295f
C168 B.t1 VSUBS 0.091248f
C169 B.t0 VSUBS 0.257536f
C170 B.n26 VSUBS 0.082406f
C171 B.n27 VSUBS 0.068823f
C172 B.n28 VSUBS 0.007901f
C173 B.n29 VSUBS 0.007901f
C174 B.n30 VSUBS 0.007901f
C175 B.n31 VSUBS 0.007901f
C176 B.t11 VSUBS 0.079295f
C177 B.t10 VSUBS 0.091248f
C178 B.t9 VSUBS 0.257536f
C179 B.n32 VSUBS 0.082406f
C180 B.n33 VSUBS 0.068823f
C181 B.n34 VSUBS 0.007901f
C182 B.n35 VSUBS 0.007901f
C183 B.n36 VSUBS 0.007901f
C184 B.n37 VSUBS 0.007901f
C185 B.n38 VSUBS 0.007901f
C186 B.n39 VSUBS 0.007901f
C187 B.n40 VSUBS 0.007901f
C188 B.n41 VSUBS 0.019375f
C189 B.n42 VSUBS 0.007901f
C190 B.n43 VSUBS 0.007901f
C191 B.n44 VSUBS 0.007901f
C192 B.n45 VSUBS 0.007901f
C193 B.n46 VSUBS 0.007901f
C194 B.n47 VSUBS 0.007901f
C195 B.n48 VSUBS 0.007901f
C196 B.n49 VSUBS 0.007901f
C197 B.n50 VSUBS 0.007901f
C198 B.n51 VSUBS 0.007901f
C199 B.n52 VSUBS 0.007901f
C200 B.n53 VSUBS 0.007901f
C201 B.n54 VSUBS 0.007901f
C202 B.n55 VSUBS 0.007901f
C203 B.n56 VSUBS 0.007901f
C204 B.n57 VSUBS 0.007901f
C205 B.n58 VSUBS 0.007901f
C206 B.n59 VSUBS 0.007901f
C207 B.n60 VSUBS 0.007901f
C208 B.n61 VSUBS 0.007901f
C209 B.n62 VSUBS 0.007901f
C210 B.n63 VSUBS 0.007901f
C211 B.n64 VSUBS 0.007901f
C212 B.n65 VSUBS 0.007901f
C213 B.n66 VSUBS 0.007901f
C214 B.n67 VSUBS 0.007901f
C215 B.n68 VSUBS 0.007901f
C216 B.n69 VSUBS 0.007901f
C217 B.n70 VSUBS 0.007901f
C218 B.n71 VSUBS 0.007901f
C219 B.n72 VSUBS 0.019375f
C220 B.n73 VSUBS 0.007901f
C221 B.n74 VSUBS 0.007901f
C222 B.n75 VSUBS 0.007901f
C223 B.n76 VSUBS 0.007901f
C224 B.n77 VSUBS 0.007901f
C225 B.n78 VSUBS 0.007901f
C226 B.n79 VSUBS 0.007901f
C227 B.t7 VSUBS 0.079295f
C228 B.t8 VSUBS 0.091248f
C229 B.t6 VSUBS 0.257536f
C230 B.n80 VSUBS 0.082406f
C231 B.n81 VSUBS 0.068823f
C232 B.n82 VSUBS 0.018305f
C233 B.n83 VSUBS 0.007901f
C234 B.n84 VSUBS 0.007901f
C235 B.n85 VSUBS 0.007901f
C236 B.n86 VSUBS 0.007901f
C237 B.n87 VSUBS 0.007901f
C238 B.t4 VSUBS 0.079295f
C239 B.t5 VSUBS 0.091248f
C240 B.t3 VSUBS 0.257536f
C241 B.n88 VSUBS 0.082406f
C242 B.n89 VSUBS 0.068823f
C243 B.n90 VSUBS 0.007901f
C244 B.n91 VSUBS 0.007901f
C245 B.n92 VSUBS 0.007901f
C246 B.n93 VSUBS 0.007901f
C247 B.n94 VSUBS 0.007901f
C248 B.n95 VSUBS 0.007901f
C249 B.n96 VSUBS 0.019895f
C250 B.n97 VSUBS 0.007901f
C251 B.n98 VSUBS 0.007901f
C252 B.n99 VSUBS 0.007901f
C253 B.n100 VSUBS 0.007901f
C254 B.n101 VSUBS 0.007901f
C255 B.n102 VSUBS 0.007901f
C256 B.n103 VSUBS 0.007901f
C257 B.n104 VSUBS 0.007901f
C258 B.n105 VSUBS 0.007901f
C259 B.n106 VSUBS 0.007901f
C260 B.n107 VSUBS 0.007901f
C261 B.n108 VSUBS 0.007901f
C262 B.n109 VSUBS 0.007901f
C263 B.n110 VSUBS 0.007901f
C264 B.n111 VSUBS 0.007901f
C265 B.n112 VSUBS 0.007901f
C266 B.n113 VSUBS 0.007901f
C267 B.n114 VSUBS 0.007901f
C268 B.n115 VSUBS 0.007901f
C269 B.n116 VSUBS 0.007901f
C270 B.n117 VSUBS 0.007901f
C271 B.n118 VSUBS 0.007901f
C272 B.n119 VSUBS 0.007901f
C273 B.n120 VSUBS 0.007901f
C274 B.n121 VSUBS 0.007901f
C275 B.n122 VSUBS 0.007901f
C276 B.n123 VSUBS 0.007901f
C277 B.n124 VSUBS 0.007901f
C278 B.n125 VSUBS 0.007901f
C279 B.n126 VSUBS 0.007901f
C280 B.n127 VSUBS 0.007901f
C281 B.n128 VSUBS 0.007901f
C282 B.n129 VSUBS 0.007901f
C283 B.n130 VSUBS 0.007901f
C284 B.n131 VSUBS 0.007901f
C285 B.n132 VSUBS 0.007901f
C286 B.n133 VSUBS 0.007901f
C287 B.n134 VSUBS 0.007901f
C288 B.n135 VSUBS 0.007901f
C289 B.n136 VSUBS 0.007901f
C290 B.n137 VSUBS 0.007901f
C291 B.n138 VSUBS 0.007901f
C292 B.n139 VSUBS 0.007901f
C293 B.n140 VSUBS 0.007901f
C294 B.n141 VSUBS 0.007901f
C295 B.n142 VSUBS 0.007901f
C296 B.n143 VSUBS 0.007901f
C297 B.n144 VSUBS 0.007901f
C298 B.n145 VSUBS 0.007901f
C299 B.n146 VSUBS 0.007901f
C300 B.n147 VSUBS 0.007901f
C301 B.n148 VSUBS 0.007901f
C302 B.n149 VSUBS 0.007901f
C303 B.n150 VSUBS 0.007901f
C304 B.n151 VSUBS 0.007901f
C305 B.n152 VSUBS 0.007901f
C306 B.n153 VSUBS 0.007901f
C307 B.n154 VSUBS 0.007901f
C308 B.n155 VSUBS 0.019375f
C309 B.n156 VSUBS 0.019375f
C310 B.n157 VSUBS 0.019895f
C311 B.n158 VSUBS 0.007901f
C312 B.n159 VSUBS 0.007901f
C313 B.n160 VSUBS 0.007901f
C314 B.n161 VSUBS 0.007901f
C315 B.n162 VSUBS 0.007901f
C316 B.n163 VSUBS 0.007901f
C317 B.n164 VSUBS 0.007901f
C318 B.n165 VSUBS 0.007901f
C319 B.n166 VSUBS 0.007901f
C320 B.n167 VSUBS 0.007901f
C321 B.n168 VSUBS 0.007901f
C322 B.n169 VSUBS 0.007901f
C323 B.n170 VSUBS 0.007901f
C324 B.n171 VSUBS 0.007901f
C325 B.n172 VSUBS 0.007901f
C326 B.n173 VSUBS 0.007901f
C327 B.n174 VSUBS 0.007901f
C328 B.n175 VSUBS 0.007901f
C329 B.n176 VSUBS 0.007901f
C330 B.n177 VSUBS 0.007901f
C331 B.n178 VSUBS 0.005461f
C332 B.n179 VSUBS 0.018305f
C333 B.n180 VSUBS 0.00639f
C334 B.n181 VSUBS 0.007901f
C335 B.n182 VSUBS 0.007901f
C336 B.n183 VSUBS 0.007901f
C337 B.n184 VSUBS 0.007901f
C338 B.n185 VSUBS 0.007901f
C339 B.n186 VSUBS 0.007901f
C340 B.n187 VSUBS 0.007901f
C341 B.n188 VSUBS 0.007901f
C342 B.n189 VSUBS 0.007901f
C343 B.n190 VSUBS 0.007901f
C344 B.n191 VSUBS 0.007901f
C345 B.n192 VSUBS 0.00639f
C346 B.n193 VSUBS 0.007901f
C347 B.n194 VSUBS 0.007901f
C348 B.n195 VSUBS 0.005461f
C349 B.n196 VSUBS 0.007901f
C350 B.n197 VSUBS 0.007901f
C351 B.n198 VSUBS 0.007901f
C352 B.n199 VSUBS 0.007901f
C353 B.n200 VSUBS 0.007901f
C354 B.n201 VSUBS 0.007901f
C355 B.n202 VSUBS 0.007901f
C356 B.n203 VSUBS 0.007901f
C357 B.n204 VSUBS 0.007901f
C358 B.n205 VSUBS 0.007901f
C359 B.n206 VSUBS 0.007901f
C360 B.n207 VSUBS 0.007901f
C361 B.n208 VSUBS 0.007901f
C362 B.n209 VSUBS 0.007901f
C363 B.n210 VSUBS 0.007901f
C364 B.n211 VSUBS 0.007901f
C365 B.n212 VSUBS 0.007901f
C366 B.n213 VSUBS 0.007901f
C367 B.n214 VSUBS 0.007901f
C368 B.n215 VSUBS 0.019895f
C369 B.n216 VSUBS 0.019895f
C370 B.n217 VSUBS 0.019375f
C371 B.n218 VSUBS 0.007901f
C372 B.n219 VSUBS 0.007901f
C373 B.n220 VSUBS 0.007901f
C374 B.n221 VSUBS 0.007901f
C375 B.n222 VSUBS 0.007901f
C376 B.n223 VSUBS 0.007901f
C377 B.n224 VSUBS 0.007901f
C378 B.n225 VSUBS 0.007901f
C379 B.n226 VSUBS 0.007901f
C380 B.n227 VSUBS 0.007901f
C381 B.n228 VSUBS 0.007901f
C382 B.n229 VSUBS 0.007901f
C383 B.n230 VSUBS 0.007901f
C384 B.n231 VSUBS 0.007901f
C385 B.n232 VSUBS 0.007901f
C386 B.n233 VSUBS 0.007901f
C387 B.n234 VSUBS 0.007901f
C388 B.n235 VSUBS 0.007901f
C389 B.n236 VSUBS 0.007901f
C390 B.n237 VSUBS 0.007901f
C391 B.n238 VSUBS 0.007901f
C392 B.n239 VSUBS 0.007901f
C393 B.n240 VSUBS 0.007901f
C394 B.n241 VSUBS 0.007901f
C395 B.n242 VSUBS 0.007901f
C396 B.n243 VSUBS 0.007901f
C397 B.n244 VSUBS 0.007901f
C398 B.n245 VSUBS 0.007901f
C399 B.n246 VSUBS 0.007901f
C400 B.n247 VSUBS 0.007901f
C401 B.n248 VSUBS 0.007901f
C402 B.n249 VSUBS 0.007901f
C403 B.n250 VSUBS 0.007901f
C404 B.n251 VSUBS 0.007901f
C405 B.n252 VSUBS 0.007901f
C406 B.n253 VSUBS 0.007901f
C407 B.n254 VSUBS 0.007901f
C408 B.n255 VSUBS 0.007901f
C409 B.n256 VSUBS 0.007901f
C410 B.n257 VSUBS 0.007901f
C411 B.n258 VSUBS 0.007901f
C412 B.n259 VSUBS 0.007901f
C413 B.n260 VSUBS 0.007901f
C414 B.n261 VSUBS 0.007901f
C415 B.n262 VSUBS 0.007901f
C416 B.n263 VSUBS 0.007901f
C417 B.n264 VSUBS 0.007901f
C418 B.n265 VSUBS 0.007901f
C419 B.n266 VSUBS 0.007901f
C420 B.n267 VSUBS 0.007901f
C421 B.n268 VSUBS 0.007901f
C422 B.n269 VSUBS 0.007901f
C423 B.n270 VSUBS 0.007901f
C424 B.n271 VSUBS 0.007901f
C425 B.n272 VSUBS 0.007901f
C426 B.n273 VSUBS 0.007901f
C427 B.n274 VSUBS 0.007901f
C428 B.n275 VSUBS 0.007901f
C429 B.n276 VSUBS 0.007901f
C430 B.n277 VSUBS 0.007901f
C431 B.n278 VSUBS 0.007901f
C432 B.n279 VSUBS 0.007901f
C433 B.n280 VSUBS 0.007901f
C434 B.n281 VSUBS 0.007901f
C435 B.n282 VSUBS 0.007901f
C436 B.n283 VSUBS 0.007901f
C437 B.n284 VSUBS 0.007901f
C438 B.n285 VSUBS 0.007901f
C439 B.n286 VSUBS 0.007901f
C440 B.n287 VSUBS 0.007901f
C441 B.n288 VSUBS 0.007901f
C442 B.n289 VSUBS 0.007901f
C443 B.n290 VSUBS 0.007901f
C444 B.n291 VSUBS 0.007901f
C445 B.n292 VSUBS 0.007901f
C446 B.n293 VSUBS 0.007901f
C447 B.n294 VSUBS 0.007901f
C448 B.n295 VSUBS 0.007901f
C449 B.n296 VSUBS 0.007901f
C450 B.n297 VSUBS 0.007901f
C451 B.n298 VSUBS 0.007901f
C452 B.n299 VSUBS 0.007901f
C453 B.n300 VSUBS 0.007901f
C454 B.n301 VSUBS 0.007901f
C455 B.n302 VSUBS 0.007901f
C456 B.n303 VSUBS 0.007901f
C457 B.n304 VSUBS 0.007901f
C458 B.n305 VSUBS 0.007901f
C459 B.n306 VSUBS 0.007901f
C460 B.n307 VSUBS 0.007901f
C461 B.n308 VSUBS 0.007901f
C462 B.n309 VSUBS 0.007901f
C463 B.n310 VSUBS 0.020228f
C464 B.n311 VSUBS 0.019042f
C465 B.n312 VSUBS 0.019895f
C466 B.n313 VSUBS 0.007901f
C467 B.n314 VSUBS 0.007901f
C468 B.n315 VSUBS 0.007901f
C469 B.n316 VSUBS 0.007901f
C470 B.n317 VSUBS 0.007901f
C471 B.n318 VSUBS 0.007901f
C472 B.n319 VSUBS 0.007901f
C473 B.n320 VSUBS 0.007901f
C474 B.n321 VSUBS 0.007901f
C475 B.n322 VSUBS 0.007901f
C476 B.n323 VSUBS 0.007901f
C477 B.n324 VSUBS 0.007901f
C478 B.n325 VSUBS 0.007901f
C479 B.n326 VSUBS 0.007901f
C480 B.n327 VSUBS 0.007901f
C481 B.n328 VSUBS 0.007901f
C482 B.n329 VSUBS 0.007901f
C483 B.n330 VSUBS 0.007901f
C484 B.n331 VSUBS 0.007901f
C485 B.n332 VSUBS 0.007901f
C486 B.n333 VSUBS 0.005461f
C487 B.n334 VSUBS 0.018305f
C488 B.n335 VSUBS 0.00639f
C489 B.n336 VSUBS 0.007901f
C490 B.n337 VSUBS 0.007901f
C491 B.n338 VSUBS 0.007901f
C492 B.n339 VSUBS 0.007901f
C493 B.n340 VSUBS 0.007901f
C494 B.n341 VSUBS 0.007901f
C495 B.n342 VSUBS 0.007901f
C496 B.n343 VSUBS 0.007901f
C497 B.n344 VSUBS 0.007901f
C498 B.n345 VSUBS 0.007901f
C499 B.n346 VSUBS 0.007901f
C500 B.n347 VSUBS 0.00639f
C501 B.n348 VSUBS 0.018305f
C502 B.n349 VSUBS 0.005461f
C503 B.n350 VSUBS 0.007901f
C504 B.n351 VSUBS 0.007901f
C505 B.n352 VSUBS 0.007901f
C506 B.n353 VSUBS 0.007901f
C507 B.n354 VSUBS 0.007901f
C508 B.n355 VSUBS 0.007901f
C509 B.n356 VSUBS 0.007901f
C510 B.n357 VSUBS 0.007901f
C511 B.n358 VSUBS 0.007901f
C512 B.n359 VSUBS 0.007901f
C513 B.n360 VSUBS 0.007901f
C514 B.n361 VSUBS 0.007901f
C515 B.n362 VSUBS 0.007901f
C516 B.n363 VSUBS 0.007901f
C517 B.n364 VSUBS 0.007901f
C518 B.n365 VSUBS 0.007901f
C519 B.n366 VSUBS 0.007901f
C520 B.n367 VSUBS 0.007901f
C521 B.n368 VSUBS 0.007901f
C522 B.n369 VSUBS 0.007901f
C523 B.n370 VSUBS 0.019895f
C524 B.n371 VSUBS 0.019895f
C525 B.n372 VSUBS 0.019375f
C526 B.n373 VSUBS 0.007901f
C527 B.n374 VSUBS 0.007901f
C528 B.n375 VSUBS 0.007901f
C529 B.n376 VSUBS 0.007901f
C530 B.n377 VSUBS 0.007901f
C531 B.n378 VSUBS 0.007901f
C532 B.n379 VSUBS 0.007901f
C533 B.n380 VSUBS 0.007901f
C534 B.n381 VSUBS 0.007901f
C535 B.n382 VSUBS 0.007901f
C536 B.n383 VSUBS 0.007901f
C537 B.n384 VSUBS 0.007901f
C538 B.n385 VSUBS 0.007901f
C539 B.n386 VSUBS 0.007901f
C540 B.n387 VSUBS 0.007901f
C541 B.n388 VSUBS 0.007901f
C542 B.n389 VSUBS 0.007901f
C543 B.n390 VSUBS 0.007901f
C544 B.n391 VSUBS 0.007901f
C545 B.n392 VSUBS 0.007901f
C546 B.n393 VSUBS 0.007901f
C547 B.n394 VSUBS 0.007901f
C548 B.n395 VSUBS 0.007901f
C549 B.n396 VSUBS 0.007901f
C550 B.n397 VSUBS 0.007901f
C551 B.n398 VSUBS 0.007901f
C552 B.n399 VSUBS 0.007901f
C553 B.n400 VSUBS 0.007901f
C554 B.n401 VSUBS 0.007901f
C555 B.n402 VSUBS 0.007901f
C556 B.n403 VSUBS 0.007901f
C557 B.n404 VSUBS 0.007901f
C558 B.n405 VSUBS 0.007901f
C559 B.n406 VSUBS 0.007901f
C560 B.n407 VSUBS 0.007901f
C561 B.n408 VSUBS 0.007901f
C562 B.n409 VSUBS 0.007901f
C563 B.n410 VSUBS 0.007901f
C564 B.n411 VSUBS 0.007901f
C565 B.n412 VSUBS 0.007901f
C566 B.n413 VSUBS 0.007901f
C567 B.n414 VSUBS 0.007901f
C568 B.n415 VSUBS 0.007901f
C569 B.n416 VSUBS 0.007901f
C570 B.n417 VSUBS 0.007901f
C571 B.n418 VSUBS 0.007901f
C572 B.n419 VSUBS 0.01789f
.ends

