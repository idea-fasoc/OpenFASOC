* NGSPICE file created from diff_pair_sample_1118.ext - technology: sky130A

.subckt diff_pair_sample_1118 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t8 VP.t0 VDD1.t5 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=1.54275 ps=9.68 w=9.35 l=3.27
X1 B.t11 B.t9 B.t10 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=0 ps=0 w=9.35 l=3.27
X2 VDD1.t0 VP.t1 VTAIL.t7 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=3.6465 ps=19.48 w=9.35 l=3.27
X3 B.t8 B.t6 B.t7 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=0 ps=0 w=9.35 l=3.27
X4 VDD2.t5 VN.t0 VTAIL.t2 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=1.54275 ps=9.68 w=9.35 l=3.27
X5 B.t5 B.t3 B.t4 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=0 ps=0 w=9.35 l=3.27
X6 VDD2.t4 VN.t1 VTAIL.t0 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=3.6465 ps=19.48 w=9.35 l=3.27
X7 VDD2.t3 VN.t2 VTAIL.t1 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=3.6465 ps=19.48 w=9.35 l=3.27
X8 VDD2.t2 VN.t3 VTAIL.t11 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=1.54275 ps=9.68 w=9.35 l=3.27
X9 VTAIL.t6 VP.t2 VDD1.t4 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=1.54275 ps=9.68 w=9.35 l=3.27
X10 VDD1.t3 VP.t3 VTAIL.t5 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=3.6465 ps=19.48 w=9.35 l=3.27
X11 VTAIL.t10 VN.t4 VDD2.t1 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=1.54275 ps=9.68 w=9.35 l=3.27
X12 VDD1.t1 VP.t4 VTAIL.t4 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=1.54275 ps=9.68 w=9.35 l=3.27
X13 B.t2 B.t0 B.t1 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=0 ps=0 w=9.35 l=3.27
X14 VTAIL.t9 VN.t5 VDD2.t0 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=1.54275 pd=9.68 as=1.54275 ps=9.68 w=9.35 l=3.27
X15 VDD1.t2 VP.t5 VTAIL.t3 w_n3850_n2838# sky130_fd_pr__pfet_01v8 ad=3.6465 pd=19.48 as=1.54275 ps=9.68 w=9.35 l=3.27
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t5 102.09
R22 VP.n27 VP.n8 72.9405
R23 VP.n50 VP.n0 72.9405
R24 VP.n26 VP.n9 72.9405
R25 VP.n8 VP.t4 68.9103
R26 VP.n4 VP.t0 68.9103
R27 VP.n0 VP.t1 68.9103
R28 VP.n9 VP.t3 68.9103
R29 VP.n13 VP.t2 68.9103
R30 VP.n14 VP.n13 62.0537
R31 VP.n27 VP.n26 49.4387
R32 VP.n31 VP.n6 45.3497
R33 VP.n46 VP.n2 45.3497
R34 VP.n22 VP.n11 45.3497
R35 VP.n35 VP.n6 35.6371
R36 VP.n42 VP.n2 35.6371
R37 VP.n18 VP.n11 35.6371
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 17.1274
R51 VP.n48 VP.n0 17.1274
R52 VP.n24 VP.n9 17.1274
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 4.04078
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1.n44 VDD1.n0 756.745
R81 VDD1.n93 VDD1.n49 756.745
R82 VDD1.n45 VDD1.n44 585
R83 VDD1.n43 VDD1.n42 585
R84 VDD1.n4 VDD1.n3 585
R85 VDD1.n8 VDD1.n6 585
R86 VDD1.n37 VDD1.n36 585
R87 VDD1.n35 VDD1.n34 585
R88 VDD1.n10 VDD1.n9 585
R89 VDD1.n29 VDD1.n28 585
R90 VDD1.n27 VDD1.n26 585
R91 VDD1.n14 VDD1.n13 585
R92 VDD1.n21 VDD1.n20 585
R93 VDD1.n19 VDD1.n18 585
R94 VDD1.n66 VDD1.n65 585
R95 VDD1.n68 VDD1.n67 585
R96 VDD1.n61 VDD1.n60 585
R97 VDD1.n74 VDD1.n73 585
R98 VDD1.n76 VDD1.n75 585
R99 VDD1.n57 VDD1.n56 585
R100 VDD1.n83 VDD1.n82 585
R101 VDD1.n84 VDD1.n55 585
R102 VDD1.n86 VDD1.n85 585
R103 VDD1.n53 VDD1.n52 585
R104 VDD1.n92 VDD1.n91 585
R105 VDD1.n94 VDD1.n93 585
R106 VDD1.n17 VDD1.t2 329.038
R107 VDD1.n64 VDD1.t1 329.038
R108 VDD1.n44 VDD1.n43 171.744
R109 VDD1.n43 VDD1.n3 171.744
R110 VDD1.n8 VDD1.n3 171.744
R111 VDD1.n36 VDD1.n8 171.744
R112 VDD1.n36 VDD1.n35 171.744
R113 VDD1.n35 VDD1.n9 171.744
R114 VDD1.n28 VDD1.n9 171.744
R115 VDD1.n28 VDD1.n27 171.744
R116 VDD1.n27 VDD1.n13 171.744
R117 VDD1.n20 VDD1.n13 171.744
R118 VDD1.n20 VDD1.n19 171.744
R119 VDD1.n67 VDD1.n66 171.744
R120 VDD1.n67 VDD1.n60 171.744
R121 VDD1.n74 VDD1.n60 171.744
R122 VDD1.n75 VDD1.n74 171.744
R123 VDD1.n75 VDD1.n56 171.744
R124 VDD1.n83 VDD1.n56 171.744
R125 VDD1.n84 VDD1.n83 171.744
R126 VDD1.n85 VDD1.n84 171.744
R127 VDD1.n85 VDD1.n52 171.744
R128 VDD1.n92 VDD1.n52 171.744
R129 VDD1.n93 VDD1.n92 171.744
R130 VDD1.n19 VDD1.t2 85.8723
R131 VDD1.n66 VDD1.t1 85.8723
R132 VDD1.n99 VDD1.n98 81.4346
R133 VDD1.n101 VDD1.n100 80.714
R134 VDD1 VDD1.n48 53.3832
R135 VDD1.n99 VDD1.n97 53.2697
R136 VDD1.n101 VDD1.n99 43.9966
R137 VDD1.n6 VDD1.n4 13.1884
R138 VDD1.n86 VDD1.n53 13.1884
R139 VDD1.n42 VDD1.n41 12.8005
R140 VDD1.n38 VDD1.n37 12.8005
R141 VDD1.n87 VDD1.n55 12.8005
R142 VDD1.n91 VDD1.n90 12.8005
R143 VDD1.n45 VDD1.n2 12.0247
R144 VDD1.n34 VDD1.n7 12.0247
R145 VDD1.n82 VDD1.n81 12.0247
R146 VDD1.n94 VDD1.n51 12.0247
R147 VDD1.n46 VDD1.n0 11.249
R148 VDD1.n33 VDD1.n10 11.249
R149 VDD1.n80 VDD1.n57 11.249
R150 VDD1.n95 VDD1.n49 11.249
R151 VDD1.n18 VDD1.n17 10.7239
R152 VDD1.n65 VDD1.n64 10.7239
R153 VDD1.n30 VDD1.n29 10.4732
R154 VDD1.n77 VDD1.n76 10.4732
R155 VDD1.n26 VDD1.n12 9.69747
R156 VDD1.n73 VDD1.n59 9.69747
R157 VDD1.n48 VDD1.n47 9.45567
R158 VDD1.n97 VDD1.n96 9.45567
R159 VDD1.n16 VDD1.n15 9.3005
R160 VDD1.n23 VDD1.n22 9.3005
R161 VDD1.n25 VDD1.n24 9.3005
R162 VDD1.n12 VDD1.n11 9.3005
R163 VDD1.n31 VDD1.n30 9.3005
R164 VDD1.n33 VDD1.n32 9.3005
R165 VDD1.n7 VDD1.n5 9.3005
R166 VDD1.n39 VDD1.n38 9.3005
R167 VDD1.n47 VDD1.n46 9.3005
R168 VDD1.n2 VDD1.n1 9.3005
R169 VDD1.n41 VDD1.n40 9.3005
R170 VDD1.n96 VDD1.n95 9.3005
R171 VDD1.n51 VDD1.n50 9.3005
R172 VDD1.n90 VDD1.n89 9.3005
R173 VDD1.n63 VDD1.n62 9.3005
R174 VDD1.n70 VDD1.n69 9.3005
R175 VDD1.n72 VDD1.n71 9.3005
R176 VDD1.n59 VDD1.n58 9.3005
R177 VDD1.n78 VDD1.n77 9.3005
R178 VDD1.n80 VDD1.n79 9.3005
R179 VDD1.n81 VDD1.n54 9.3005
R180 VDD1.n88 VDD1.n87 9.3005
R181 VDD1.n25 VDD1.n14 8.92171
R182 VDD1.n72 VDD1.n61 8.92171
R183 VDD1.n22 VDD1.n21 8.14595
R184 VDD1.n69 VDD1.n68 8.14595
R185 VDD1.n18 VDD1.n16 7.3702
R186 VDD1.n65 VDD1.n63 7.3702
R187 VDD1.n21 VDD1.n16 5.81868
R188 VDD1.n68 VDD1.n63 5.81868
R189 VDD1.n22 VDD1.n14 5.04292
R190 VDD1.n69 VDD1.n61 5.04292
R191 VDD1.n26 VDD1.n25 4.26717
R192 VDD1.n73 VDD1.n72 4.26717
R193 VDD1.n29 VDD1.n12 3.49141
R194 VDD1.n76 VDD1.n59 3.49141
R195 VDD1.n100 VDD1.t4 3.47697
R196 VDD1.n100 VDD1.t3 3.47697
R197 VDD1.n98 VDD1.t5 3.47697
R198 VDD1.n98 VDD1.t0 3.47697
R199 VDD1.n48 VDD1.n0 2.71565
R200 VDD1.n30 VDD1.n10 2.71565
R201 VDD1.n77 VDD1.n57 2.71565
R202 VDD1.n97 VDD1.n49 2.71565
R203 VDD1.n17 VDD1.n15 2.41283
R204 VDD1.n64 VDD1.n62 2.41283
R205 VDD1.n46 VDD1.n45 1.93989
R206 VDD1.n34 VDD1.n33 1.93989
R207 VDD1.n82 VDD1.n80 1.93989
R208 VDD1.n95 VDD1.n94 1.93989
R209 VDD1.n42 VDD1.n2 1.16414
R210 VDD1.n37 VDD1.n7 1.16414
R211 VDD1.n81 VDD1.n55 1.16414
R212 VDD1.n91 VDD1.n51 1.16414
R213 VDD1 VDD1.n101 0.718172
R214 VDD1.n41 VDD1.n4 0.388379
R215 VDD1.n38 VDD1.n6 0.388379
R216 VDD1.n87 VDD1.n86 0.388379
R217 VDD1.n90 VDD1.n53 0.388379
R218 VDD1.n47 VDD1.n1 0.155672
R219 VDD1.n40 VDD1.n1 0.155672
R220 VDD1.n40 VDD1.n39 0.155672
R221 VDD1.n39 VDD1.n5 0.155672
R222 VDD1.n32 VDD1.n5 0.155672
R223 VDD1.n32 VDD1.n31 0.155672
R224 VDD1.n31 VDD1.n11 0.155672
R225 VDD1.n24 VDD1.n11 0.155672
R226 VDD1.n24 VDD1.n23 0.155672
R227 VDD1.n23 VDD1.n15 0.155672
R228 VDD1.n70 VDD1.n62 0.155672
R229 VDD1.n71 VDD1.n70 0.155672
R230 VDD1.n71 VDD1.n58 0.155672
R231 VDD1.n78 VDD1.n58 0.155672
R232 VDD1.n79 VDD1.n78 0.155672
R233 VDD1.n79 VDD1.n54 0.155672
R234 VDD1.n88 VDD1.n54 0.155672
R235 VDD1.n89 VDD1.n88 0.155672
R236 VDD1.n89 VDD1.n50 0.155672
R237 VDD1.n96 VDD1.n50 0.155672
R238 VTAIL.n202 VTAIL.n158 756.745
R239 VTAIL.n46 VTAIL.n2 756.745
R240 VTAIL.n152 VTAIL.n108 756.745
R241 VTAIL.n100 VTAIL.n56 756.745
R242 VTAIL.n175 VTAIL.n174 585
R243 VTAIL.n177 VTAIL.n176 585
R244 VTAIL.n170 VTAIL.n169 585
R245 VTAIL.n183 VTAIL.n182 585
R246 VTAIL.n185 VTAIL.n184 585
R247 VTAIL.n166 VTAIL.n165 585
R248 VTAIL.n192 VTAIL.n191 585
R249 VTAIL.n193 VTAIL.n164 585
R250 VTAIL.n195 VTAIL.n194 585
R251 VTAIL.n162 VTAIL.n161 585
R252 VTAIL.n201 VTAIL.n200 585
R253 VTAIL.n203 VTAIL.n202 585
R254 VTAIL.n19 VTAIL.n18 585
R255 VTAIL.n21 VTAIL.n20 585
R256 VTAIL.n14 VTAIL.n13 585
R257 VTAIL.n27 VTAIL.n26 585
R258 VTAIL.n29 VTAIL.n28 585
R259 VTAIL.n10 VTAIL.n9 585
R260 VTAIL.n36 VTAIL.n35 585
R261 VTAIL.n37 VTAIL.n8 585
R262 VTAIL.n39 VTAIL.n38 585
R263 VTAIL.n6 VTAIL.n5 585
R264 VTAIL.n45 VTAIL.n44 585
R265 VTAIL.n47 VTAIL.n46 585
R266 VTAIL.n153 VTAIL.n152 585
R267 VTAIL.n151 VTAIL.n150 585
R268 VTAIL.n112 VTAIL.n111 585
R269 VTAIL.n116 VTAIL.n114 585
R270 VTAIL.n145 VTAIL.n144 585
R271 VTAIL.n143 VTAIL.n142 585
R272 VTAIL.n118 VTAIL.n117 585
R273 VTAIL.n137 VTAIL.n136 585
R274 VTAIL.n135 VTAIL.n134 585
R275 VTAIL.n122 VTAIL.n121 585
R276 VTAIL.n129 VTAIL.n128 585
R277 VTAIL.n127 VTAIL.n126 585
R278 VTAIL.n101 VTAIL.n100 585
R279 VTAIL.n99 VTAIL.n98 585
R280 VTAIL.n60 VTAIL.n59 585
R281 VTAIL.n64 VTAIL.n62 585
R282 VTAIL.n93 VTAIL.n92 585
R283 VTAIL.n91 VTAIL.n90 585
R284 VTAIL.n66 VTAIL.n65 585
R285 VTAIL.n85 VTAIL.n84 585
R286 VTAIL.n83 VTAIL.n82 585
R287 VTAIL.n70 VTAIL.n69 585
R288 VTAIL.n77 VTAIL.n76 585
R289 VTAIL.n75 VTAIL.n74 585
R290 VTAIL.n173 VTAIL.t1 329.038
R291 VTAIL.n17 VTAIL.t7 329.038
R292 VTAIL.n125 VTAIL.t5 329.038
R293 VTAIL.n73 VTAIL.t0 329.038
R294 VTAIL.n176 VTAIL.n175 171.744
R295 VTAIL.n176 VTAIL.n169 171.744
R296 VTAIL.n183 VTAIL.n169 171.744
R297 VTAIL.n184 VTAIL.n183 171.744
R298 VTAIL.n184 VTAIL.n165 171.744
R299 VTAIL.n192 VTAIL.n165 171.744
R300 VTAIL.n193 VTAIL.n192 171.744
R301 VTAIL.n194 VTAIL.n193 171.744
R302 VTAIL.n194 VTAIL.n161 171.744
R303 VTAIL.n201 VTAIL.n161 171.744
R304 VTAIL.n202 VTAIL.n201 171.744
R305 VTAIL.n20 VTAIL.n19 171.744
R306 VTAIL.n20 VTAIL.n13 171.744
R307 VTAIL.n27 VTAIL.n13 171.744
R308 VTAIL.n28 VTAIL.n27 171.744
R309 VTAIL.n28 VTAIL.n9 171.744
R310 VTAIL.n36 VTAIL.n9 171.744
R311 VTAIL.n37 VTAIL.n36 171.744
R312 VTAIL.n38 VTAIL.n37 171.744
R313 VTAIL.n38 VTAIL.n5 171.744
R314 VTAIL.n45 VTAIL.n5 171.744
R315 VTAIL.n46 VTAIL.n45 171.744
R316 VTAIL.n152 VTAIL.n151 171.744
R317 VTAIL.n151 VTAIL.n111 171.744
R318 VTAIL.n116 VTAIL.n111 171.744
R319 VTAIL.n144 VTAIL.n116 171.744
R320 VTAIL.n144 VTAIL.n143 171.744
R321 VTAIL.n143 VTAIL.n117 171.744
R322 VTAIL.n136 VTAIL.n117 171.744
R323 VTAIL.n136 VTAIL.n135 171.744
R324 VTAIL.n135 VTAIL.n121 171.744
R325 VTAIL.n128 VTAIL.n121 171.744
R326 VTAIL.n128 VTAIL.n127 171.744
R327 VTAIL.n100 VTAIL.n99 171.744
R328 VTAIL.n99 VTAIL.n59 171.744
R329 VTAIL.n64 VTAIL.n59 171.744
R330 VTAIL.n92 VTAIL.n64 171.744
R331 VTAIL.n92 VTAIL.n91 171.744
R332 VTAIL.n91 VTAIL.n65 171.744
R333 VTAIL.n84 VTAIL.n65 171.744
R334 VTAIL.n84 VTAIL.n83 171.744
R335 VTAIL.n83 VTAIL.n69 171.744
R336 VTAIL.n76 VTAIL.n69 171.744
R337 VTAIL.n76 VTAIL.n75 171.744
R338 VTAIL.n175 VTAIL.t1 85.8723
R339 VTAIL.n19 VTAIL.t7 85.8723
R340 VTAIL.n127 VTAIL.t5 85.8723
R341 VTAIL.n75 VTAIL.t0 85.8723
R342 VTAIL.n107 VTAIL.n106 64.0354
R343 VTAIL.n55 VTAIL.n54 64.0354
R344 VTAIL.n1 VTAIL.n0 64.0353
R345 VTAIL.n53 VTAIL.n52 64.0353
R346 VTAIL.n207 VTAIL.n206 34.3187
R347 VTAIL.n51 VTAIL.n50 34.3187
R348 VTAIL.n157 VTAIL.n156 34.3187
R349 VTAIL.n105 VTAIL.n104 34.3187
R350 VTAIL.n55 VTAIL.n53 26.6341
R351 VTAIL.n207 VTAIL.n157 23.5307
R352 VTAIL.n195 VTAIL.n162 13.1884
R353 VTAIL.n39 VTAIL.n6 13.1884
R354 VTAIL.n114 VTAIL.n112 13.1884
R355 VTAIL.n62 VTAIL.n60 13.1884
R356 VTAIL.n196 VTAIL.n164 12.8005
R357 VTAIL.n200 VTAIL.n199 12.8005
R358 VTAIL.n40 VTAIL.n8 12.8005
R359 VTAIL.n44 VTAIL.n43 12.8005
R360 VTAIL.n150 VTAIL.n149 12.8005
R361 VTAIL.n146 VTAIL.n145 12.8005
R362 VTAIL.n98 VTAIL.n97 12.8005
R363 VTAIL.n94 VTAIL.n93 12.8005
R364 VTAIL.n191 VTAIL.n190 12.0247
R365 VTAIL.n203 VTAIL.n160 12.0247
R366 VTAIL.n35 VTAIL.n34 12.0247
R367 VTAIL.n47 VTAIL.n4 12.0247
R368 VTAIL.n153 VTAIL.n110 12.0247
R369 VTAIL.n142 VTAIL.n115 12.0247
R370 VTAIL.n101 VTAIL.n58 12.0247
R371 VTAIL.n90 VTAIL.n63 12.0247
R372 VTAIL.n189 VTAIL.n166 11.249
R373 VTAIL.n204 VTAIL.n158 11.249
R374 VTAIL.n33 VTAIL.n10 11.249
R375 VTAIL.n48 VTAIL.n2 11.249
R376 VTAIL.n154 VTAIL.n108 11.249
R377 VTAIL.n141 VTAIL.n118 11.249
R378 VTAIL.n102 VTAIL.n56 11.249
R379 VTAIL.n89 VTAIL.n66 11.249
R380 VTAIL.n174 VTAIL.n173 10.7239
R381 VTAIL.n18 VTAIL.n17 10.7239
R382 VTAIL.n126 VTAIL.n125 10.7239
R383 VTAIL.n74 VTAIL.n73 10.7239
R384 VTAIL.n186 VTAIL.n185 10.4732
R385 VTAIL.n30 VTAIL.n29 10.4732
R386 VTAIL.n138 VTAIL.n137 10.4732
R387 VTAIL.n86 VTAIL.n85 10.4732
R388 VTAIL.n182 VTAIL.n168 9.69747
R389 VTAIL.n26 VTAIL.n12 9.69747
R390 VTAIL.n134 VTAIL.n120 9.69747
R391 VTAIL.n82 VTAIL.n68 9.69747
R392 VTAIL.n206 VTAIL.n205 9.45567
R393 VTAIL.n50 VTAIL.n49 9.45567
R394 VTAIL.n156 VTAIL.n155 9.45567
R395 VTAIL.n104 VTAIL.n103 9.45567
R396 VTAIL.n205 VTAIL.n204 9.3005
R397 VTAIL.n160 VTAIL.n159 9.3005
R398 VTAIL.n199 VTAIL.n198 9.3005
R399 VTAIL.n172 VTAIL.n171 9.3005
R400 VTAIL.n179 VTAIL.n178 9.3005
R401 VTAIL.n181 VTAIL.n180 9.3005
R402 VTAIL.n168 VTAIL.n167 9.3005
R403 VTAIL.n187 VTAIL.n186 9.3005
R404 VTAIL.n189 VTAIL.n188 9.3005
R405 VTAIL.n190 VTAIL.n163 9.3005
R406 VTAIL.n197 VTAIL.n196 9.3005
R407 VTAIL.n49 VTAIL.n48 9.3005
R408 VTAIL.n4 VTAIL.n3 9.3005
R409 VTAIL.n43 VTAIL.n42 9.3005
R410 VTAIL.n16 VTAIL.n15 9.3005
R411 VTAIL.n23 VTAIL.n22 9.3005
R412 VTAIL.n25 VTAIL.n24 9.3005
R413 VTAIL.n12 VTAIL.n11 9.3005
R414 VTAIL.n31 VTAIL.n30 9.3005
R415 VTAIL.n33 VTAIL.n32 9.3005
R416 VTAIL.n34 VTAIL.n7 9.3005
R417 VTAIL.n41 VTAIL.n40 9.3005
R418 VTAIL.n124 VTAIL.n123 9.3005
R419 VTAIL.n131 VTAIL.n130 9.3005
R420 VTAIL.n133 VTAIL.n132 9.3005
R421 VTAIL.n120 VTAIL.n119 9.3005
R422 VTAIL.n139 VTAIL.n138 9.3005
R423 VTAIL.n141 VTAIL.n140 9.3005
R424 VTAIL.n115 VTAIL.n113 9.3005
R425 VTAIL.n147 VTAIL.n146 9.3005
R426 VTAIL.n155 VTAIL.n154 9.3005
R427 VTAIL.n110 VTAIL.n109 9.3005
R428 VTAIL.n149 VTAIL.n148 9.3005
R429 VTAIL.n72 VTAIL.n71 9.3005
R430 VTAIL.n79 VTAIL.n78 9.3005
R431 VTAIL.n81 VTAIL.n80 9.3005
R432 VTAIL.n68 VTAIL.n67 9.3005
R433 VTAIL.n87 VTAIL.n86 9.3005
R434 VTAIL.n89 VTAIL.n88 9.3005
R435 VTAIL.n63 VTAIL.n61 9.3005
R436 VTAIL.n95 VTAIL.n94 9.3005
R437 VTAIL.n103 VTAIL.n102 9.3005
R438 VTAIL.n58 VTAIL.n57 9.3005
R439 VTAIL.n97 VTAIL.n96 9.3005
R440 VTAIL.n181 VTAIL.n170 8.92171
R441 VTAIL.n25 VTAIL.n14 8.92171
R442 VTAIL.n133 VTAIL.n122 8.92171
R443 VTAIL.n81 VTAIL.n70 8.92171
R444 VTAIL.n178 VTAIL.n177 8.14595
R445 VTAIL.n22 VTAIL.n21 8.14595
R446 VTAIL.n130 VTAIL.n129 8.14595
R447 VTAIL.n78 VTAIL.n77 8.14595
R448 VTAIL.n174 VTAIL.n172 7.3702
R449 VTAIL.n18 VTAIL.n16 7.3702
R450 VTAIL.n126 VTAIL.n124 7.3702
R451 VTAIL.n74 VTAIL.n72 7.3702
R452 VTAIL.n177 VTAIL.n172 5.81868
R453 VTAIL.n21 VTAIL.n16 5.81868
R454 VTAIL.n129 VTAIL.n124 5.81868
R455 VTAIL.n77 VTAIL.n72 5.81868
R456 VTAIL.n178 VTAIL.n170 5.04292
R457 VTAIL.n22 VTAIL.n14 5.04292
R458 VTAIL.n130 VTAIL.n122 5.04292
R459 VTAIL.n78 VTAIL.n70 5.04292
R460 VTAIL.n182 VTAIL.n181 4.26717
R461 VTAIL.n26 VTAIL.n25 4.26717
R462 VTAIL.n134 VTAIL.n133 4.26717
R463 VTAIL.n82 VTAIL.n81 4.26717
R464 VTAIL.n185 VTAIL.n168 3.49141
R465 VTAIL.n29 VTAIL.n12 3.49141
R466 VTAIL.n137 VTAIL.n120 3.49141
R467 VTAIL.n85 VTAIL.n68 3.49141
R468 VTAIL.n0 VTAIL.t11 3.47697
R469 VTAIL.n0 VTAIL.t10 3.47697
R470 VTAIL.n52 VTAIL.t4 3.47697
R471 VTAIL.n52 VTAIL.t8 3.47697
R472 VTAIL.n106 VTAIL.t3 3.47697
R473 VTAIL.n106 VTAIL.t6 3.47697
R474 VTAIL.n54 VTAIL.t2 3.47697
R475 VTAIL.n54 VTAIL.t9 3.47697
R476 VTAIL.n105 VTAIL.n55 3.10395
R477 VTAIL.n157 VTAIL.n107 3.10395
R478 VTAIL.n53 VTAIL.n51 3.10395
R479 VTAIL.n186 VTAIL.n166 2.71565
R480 VTAIL.n206 VTAIL.n158 2.71565
R481 VTAIL.n30 VTAIL.n10 2.71565
R482 VTAIL.n50 VTAIL.n2 2.71565
R483 VTAIL.n156 VTAIL.n108 2.71565
R484 VTAIL.n138 VTAIL.n118 2.71565
R485 VTAIL.n104 VTAIL.n56 2.71565
R486 VTAIL.n86 VTAIL.n66 2.71565
R487 VTAIL.n173 VTAIL.n171 2.41283
R488 VTAIL.n17 VTAIL.n15 2.41283
R489 VTAIL.n125 VTAIL.n123 2.41283
R490 VTAIL.n73 VTAIL.n71 2.41283
R491 VTAIL VTAIL.n207 2.2699
R492 VTAIL.n107 VTAIL.n105 2.02205
R493 VTAIL.n51 VTAIL.n1 2.02205
R494 VTAIL.n191 VTAIL.n189 1.93989
R495 VTAIL.n204 VTAIL.n203 1.93989
R496 VTAIL.n35 VTAIL.n33 1.93989
R497 VTAIL.n48 VTAIL.n47 1.93989
R498 VTAIL.n154 VTAIL.n153 1.93989
R499 VTAIL.n142 VTAIL.n141 1.93989
R500 VTAIL.n102 VTAIL.n101 1.93989
R501 VTAIL.n90 VTAIL.n89 1.93989
R502 VTAIL.n190 VTAIL.n164 1.16414
R503 VTAIL.n200 VTAIL.n160 1.16414
R504 VTAIL.n34 VTAIL.n8 1.16414
R505 VTAIL.n44 VTAIL.n4 1.16414
R506 VTAIL.n150 VTAIL.n110 1.16414
R507 VTAIL.n145 VTAIL.n115 1.16414
R508 VTAIL.n98 VTAIL.n58 1.16414
R509 VTAIL.n93 VTAIL.n63 1.16414
R510 VTAIL VTAIL.n1 0.834552
R511 VTAIL.n196 VTAIL.n195 0.388379
R512 VTAIL.n199 VTAIL.n162 0.388379
R513 VTAIL.n40 VTAIL.n39 0.388379
R514 VTAIL.n43 VTAIL.n6 0.388379
R515 VTAIL.n149 VTAIL.n112 0.388379
R516 VTAIL.n146 VTAIL.n114 0.388379
R517 VTAIL.n97 VTAIL.n60 0.388379
R518 VTAIL.n94 VTAIL.n62 0.388379
R519 VTAIL.n179 VTAIL.n171 0.155672
R520 VTAIL.n180 VTAIL.n179 0.155672
R521 VTAIL.n180 VTAIL.n167 0.155672
R522 VTAIL.n187 VTAIL.n167 0.155672
R523 VTAIL.n188 VTAIL.n187 0.155672
R524 VTAIL.n188 VTAIL.n163 0.155672
R525 VTAIL.n197 VTAIL.n163 0.155672
R526 VTAIL.n198 VTAIL.n197 0.155672
R527 VTAIL.n198 VTAIL.n159 0.155672
R528 VTAIL.n205 VTAIL.n159 0.155672
R529 VTAIL.n23 VTAIL.n15 0.155672
R530 VTAIL.n24 VTAIL.n23 0.155672
R531 VTAIL.n24 VTAIL.n11 0.155672
R532 VTAIL.n31 VTAIL.n11 0.155672
R533 VTAIL.n32 VTAIL.n31 0.155672
R534 VTAIL.n32 VTAIL.n7 0.155672
R535 VTAIL.n41 VTAIL.n7 0.155672
R536 VTAIL.n42 VTAIL.n41 0.155672
R537 VTAIL.n42 VTAIL.n3 0.155672
R538 VTAIL.n49 VTAIL.n3 0.155672
R539 VTAIL.n155 VTAIL.n109 0.155672
R540 VTAIL.n148 VTAIL.n109 0.155672
R541 VTAIL.n148 VTAIL.n147 0.155672
R542 VTAIL.n147 VTAIL.n113 0.155672
R543 VTAIL.n140 VTAIL.n113 0.155672
R544 VTAIL.n140 VTAIL.n139 0.155672
R545 VTAIL.n139 VTAIL.n119 0.155672
R546 VTAIL.n132 VTAIL.n119 0.155672
R547 VTAIL.n132 VTAIL.n131 0.155672
R548 VTAIL.n131 VTAIL.n123 0.155672
R549 VTAIL.n103 VTAIL.n57 0.155672
R550 VTAIL.n96 VTAIL.n57 0.155672
R551 VTAIL.n96 VTAIL.n95 0.155672
R552 VTAIL.n95 VTAIL.n61 0.155672
R553 VTAIL.n88 VTAIL.n61 0.155672
R554 VTAIL.n88 VTAIL.n87 0.155672
R555 VTAIL.n87 VTAIL.n67 0.155672
R556 VTAIL.n80 VTAIL.n67 0.155672
R557 VTAIL.n80 VTAIL.n79 0.155672
R558 VTAIL.n79 VTAIL.n71 0.155672
R559 B.n378 B.n121 585
R560 B.n377 B.n376 585
R561 B.n375 B.n122 585
R562 B.n374 B.n373 585
R563 B.n372 B.n123 585
R564 B.n371 B.n370 585
R565 B.n369 B.n124 585
R566 B.n368 B.n367 585
R567 B.n366 B.n125 585
R568 B.n365 B.n364 585
R569 B.n363 B.n126 585
R570 B.n362 B.n361 585
R571 B.n360 B.n127 585
R572 B.n359 B.n358 585
R573 B.n357 B.n128 585
R574 B.n356 B.n355 585
R575 B.n354 B.n129 585
R576 B.n353 B.n352 585
R577 B.n351 B.n130 585
R578 B.n350 B.n349 585
R579 B.n348 B.n131 585
R580 B.n347 B.n346 585
R581 B.n345 B.n132 585
R582 B.n344 B.n343 585
R583 B.n342 B.n133 585
R584 B.n341 B.n340 585
R585 B.n339 B.n134 585
R586 B.n338 B.n337 585
R587 B.n336 B.n135 585
R588 B.n335 B.n334 585
R589 B.n333 B.n136 585
R590 B.n332 B.n331 585
R591 B.n330 B.n137 585
R592 B.n329 B.n328 585
R593 B.n327 B.n326 585
R594 B.n325 B.n141 585
R595 B.n324 B.n323 585
R596 B.n322 B.n142 585
R597 B.n321 B.n320 585
R598 B.n319 B.n143 585
R599 B.n318 B.n317 585
R600 B.n316 B.n144 585
R601 B.n315 B.n314 585
R602 B.n312 B.n145 585
R603 B.n311 B.n310 585
R604 B.n309 B.n148 585
R605 B.n308 B.n307 585
R606 B.n306 B.n149 585
R607 B.n305 B.n304 585
R608 B.n303 B.n150 585
R609 B.n302 B.n301 585
R610 B.n300 B.n151 585
R611 B.n299 B.n298 585
R612 B.n297 B.n152 585
R613 B.n296 B.n295 585
R614 B.n294 B.n153 585
R615 B.n293 B.n292 585
R616 B.n291 B.n154 585
R617 B.n290 B.n289 585
R618 B.n288 B.n155 585
R619 B.n287 B.n286 585
R620 B.n285 B.n156 585
R621 B.n284 B.n283 585
R622 B.n282 B.n157 585
R623 B.n281 B.n280 585
R624 B.n279 B.n158 585
R625 B.n278 B.n277 585
R626 B.n276 B.n159 585
R627 B.n275 B.n274 585
R628 B.n273 B.n160 585
R629 B.n272 B.n271 585
R630 B.n270 B.n161 585
R631 B.n269 B.n268 585
R632 B.n267 B.n162 585
R633 B.n266 B.n265 585
R634 B.n264 B.n163 585
R635 B.n263 B.n262 585
R636 B.n380 B.n379 585
R637 B.n381 B.n120 585
R638 B.n383 B.n382 585
R639 B.n384 B.n119 585
R640 B.n386 B.n385 585
R641 B.n387 B.n118 585
R642 B.n389 B.n388 585
R643 B.n390 B.n117 585
R644 B.n392 B.n391 585
R645 B.n393 B.n116 585
R646 B.n395 B.n394 585
R647 B.n396 B.n115 585
R648 B.n398 B.n397 585
R649 B.n399 B.n114 585
R650 B.n401 B.n400 585
R651 B.n402 B.n113 585
R652 B.n404 B.n403 585
R653 B.n405 B.n112 585
R654 B.n407 B.n406 585
R655 B.n408 B.n111 585
R656 B.n410 B.n409 585
R657 B.n411 B.n110 585
R658 B.n413 B.n412 585
R659 B.n414 B.n109 585
R660 B.n416 B.n415 585
R661 B.n417 B.n108 585
R662 B.n419 B.n418 585
R663 B.n420 B.n107 585
R664 B.n422 B.n421 585
R665 B.n423 B.n106 585
R666 B.n425 B.n424 585
R667 B.n426 B.n105 585
R668 B.n428 B.n427 585
R669 B.n429 B.n104 585
R670 B.n431 B.n430 585
R671 B.n432 B.n103 585
R672 B.n434 B.n433 585
R673 B.n435 B.n102 585
R674 B.n437 B.n436 585
R675 B.n438 B.n101 585
R676 B.n440 B.n439 585
R677 B.n441 B.n100 585
R678 B.n443 B.n442 585
R679 B.n444 B.n99 585
R680 B.n446 B.n445 585
R681 B.n447 B.n98 585
R682 B.n449 B.n448 585
R683 B.n450 B.n97 585
R684 B.n452 B.n451 585
R685 B.n453 B.n96 585
R686 B.n455 B.n454 585
R687 B.n456 B.n95 585
R688 B.n458 B.n457 585
R689 B.n459 B.n94 585
R690 B.n461 B.n460 585
R691 B.n462 B.n93 585
R692 B.n464 B.n463 585
R693 B.n465 B.n92 585
R694 B.n467 B.n466 585
R695 B.n468 B.n91 585
R696 B.n470 B.n469 585
R697 B.n471 B.n90 585
R698 B.n473 B.n472 585
R699 B.n474 B.n89 585
R700 B.n476 B.n475 585
R701 B.n477 B.n88 585
R702 B.n479 B.n478 585
R703 B.n480 B.n87 585
R704 B.n482 B.n481 585
R705 B.n483 B.n86 585
R706 B.n485 B.n484 585
R707 B.n486 B.n85 585
R708 B.n488 B.n487 585
R709 B.n489 B.n84 585
R710 B.n491 B.n490 585
R711 B.n492 B.n83 585
R712 B.n494 B.n493 585
R713 B.n495 B.n82 585
R714 B.n497 B.n496 585
R715 B.n498 B.n81 585
R716 B.n500 B.n499 585
R717 B.n501 B.n80 585
R718 B.n503 B.n502 585
R719 B.n504 B.n79 585
R720 B.n506 B.n505 585
R721 B.n507 B.n78 585
R722 B.n509 B.n508 585
R723 B.n510 B.n77 585
R724 B.n512 B.n511 585
R725 B.n513 B.n76 585
R726 B.n515 B.n514 585
R727 B.n516 B.n75 585
R728 B.n518 B.n517 585
R729 B.n519 B.n74 585
R730 B.n521 B.n520 585
R731 B.n522 B.n73 585
R732 B.n524 B.n523 585
R733 B.n525 B.n72 585
R734 B.n527 B.n526 585
R735 B.n528 B.n71 585
R736 B.n530 B.n529 585
R737 B.n531 B.n70 585
R738 B.n648 B.n27 585
R739 B.n647 B.n646 585
R740 B.n645 B.n28 585
R741 B.n644 B.n643 585
R742 B.n642 B.n29 585
R743 B.n641 B.n640 585
R744 B.n639 B.n30 585
R745 B.n638 B.n637 585
R746 B.n636 B.n31 585
R747 B.n635 B.n634 585
R748 B.n633 B.n32 585
R749 B.n632 B.n631 585
R750 B.n630 B.n33 585
R751 B.n629 B.n628 585
R752 B.n627 B.n34 585
R753 B.n626 B.n625 585
R754 B.n624 B.n35 585
R755 B.n623 B.n622 585
R756 B.n621 B.n36 585
R757 B.n620 B.n619 585
R758 B.n618 B.n37 585
R759 B.n617 B.n616 585
R760 B.n615 B.n38 585
R761 B.n614 B.n613 585
R762 B.n612 B.n39 585
R763 B.n611 B.n610 585
R764 B.n609 B.n40 585
R765 B.n608 B.n607 585
R766 B.n606 B.n41 585
R767 B.n605 B.n604 585
R768 B.n603 B.n42 585
R769 B.n602 B.n601 585
R770 B.n600 B.n43 585
R771 B.n599 B.n598 585
R772 B.n597 B.n596 585
R773 B.n595 B.n47 585
R774 B.n594 B.n593 585
R775 B.n592 B.n48 585
R776 B.n591 B.n590 585
R777 B.n589 B.n49 585
R778 B.n588 B.n587 585
R779 B.n586 B.n50 585
R780 B.n585 B.n584 585
R781 B.n582 B.n51 585
R782 B.n581 B.n580 585
R783 B.n579 B.n54 585
R784 B.n578 B.n577 585
R785 B.n576 B.n55 585
R786 B.n575 B.n574 585
R787 B.n573 B.n56 585
R788 B.n572 B.n571 585
R789 B.n570 B.n57 585
R790 B.n569 B.n568 585
R791 B.n567 B.n58 585
R792 B.n566 B.n565 585
R793 B.n564 B.n59 585
R794 B.n563 B.n562 585
R795 B.n561 B.n60 585
R796 B.n560 B.n559 585
R797 B.n558 B.n61 585
R798 B.n557 B.n556 585
R799 B.n555 B.n62 585
R800 B.n554 B.n553 585
R801 B.n552 B.n63 585
R802 B.n551 B.n550 585
R803 B.n549 B.n64 585
R804 B.n548 B.n547 585
R805 B.n546 B.n65 585
R806 B.n545 B.n544 585
R807 B.n543 B.n66 585
R808 B.n542 B.n541 585
R809 B.n540 B.n67 585
R810 B.n539 B.n538 585
R811 B.n537 B.n68 585
R812 B.n536 B.n535 585
R813 B.n534 B.n69 585
R814 B.n533 B.n532 585
R815 B.n650 B.n649 585
R816 B.n651 B.n26 585
R817 B.n653 B.n652 585
R818 B.n654 B.n25 585
R819 B.n656 B.n655 585
R820 B.n657 B.n24 585
R821 B.n659 B.n658 585
R822 B.n660 B.n23 585
R823 B.n662 B.n661 585
R824 B.n663 B.n22 585
R825 B.n665 B.n664 585
R826 B.n666 B.n21 585
R827 B.n668 B.n667 585
R828 B.n669 B.n20 585
R829 B.n671 B.n670 585
R830 B.n672 B.n19 585
R831 B.n674 B.n673 585
R832 B.n675 B.n18 585
R833 B.n677 B.n676 585
R834 B.n678 B.n17 585
R835 B.n680 B.n679 585
R836 B.n681 B.n16 585
R837 B.n683 B.n682 585
R838 B.n684 B.n15 585
R839 B.n686 B.n685 585
R840 B.n687 B.n14 585
R841 B.n689 B.n688 585
R842 B.n690 B.n13 585
R843 B.n692 B.n691 585
R844 B.n693 B.n12 585
R845 B.n695 B.n694 585
R846 B.n696 B.n11 585
R847 B.n698 B.n697 585
R848 B.n699 B.n10 585
R849 B.n701 B.n700 585
R850 B.n702 B.n9 585
R851 B.n704 B.n703 585
R852 B.n705 B.n8 585
R853 B.n707 B.n706 585
R854 B.n708 B.n7 585
R855 B.n710 B.n709 585
R856 B.n711 B.n6 585
R857 B.n713 B.n712 585
R858 B.n714 B.n5 585
R859 B.n716 B.n715 585
R860 B.n717 B.n4 585
R861 B.n719 B.n718 585
R862 B.n720 B.n3 585
R863 B.n722 B.n721 585
R864 B.n723 B.n0 585
R865 B.n2 B.n1 585
R866 B.n189 B.n188 585
R867 B.n191 B.n190 585
R868 B.n192 B.n187 585
R869 B.n194 B.n193 585
R870 B.n195 B.n186 585
R871 B.n197 B.n196 585
R872 B.n198 B.n185 585
R873 B.n200 B.n199 585
R874 B.n201 B.n184 585
R875 B.n203 B.n202 585
R876 B.n204 B.n183 585
R877 B.n206 B.n205 585
R878 B.n207 B.n182 585
R879 B.n209 B.n208 585
R880 B.n210 B.n181 585
R881 B.n212 B.n211 585
R882 B.n213 B.n180 585
R883 B.n215 B.n214 585
R884 B.n216 B.n179 585
R885 B.n218 B.n217 585
R886 B.n219 B.n178 585
R887 B.n221 B.n220 585
R888 B.n222 B.n177 585
R889 B.n224 B.n223 585
R890 B.n225 B.n176 585
R891 B.n227 B.n226 585
R892 B.n228 B.n175 585
R893 B.n230 B.n229 585
R894 B.n231 B.n174 585
R895 B.n233 B.n232 585
R896 B.n234 B.n173 585
R897 B.n236 B.n235 585
R898 B.n237 B.n172 585
R899 B.n239 B.n238 585
R900 B.n240 B.n171 585
R901 B.n242 B.n241 585
R902 B.n243 B.n170 585
R903 B.n245 B.n244 585
R904 B.n246 B.n169 585
R905 B.n248 B.n247 585
R906 B.n249 B.n168 585
R907 B.n251 B.n250 585
R908 B.n252 B.n167 585
R909 B.n254 B.n253 585
R910 B.n255 B.n166 585
R911 B.n257 B.n256 585
R912 B.n258 B.n165 585
R913 B.n260 B.n259 585
R914 B.n261 B.n164 585
R915 B.n262 B.n261 511.721
R916 B.n380 B.n121 511.721
R917 B.n532 B.n531 511.721
R918 B.n650 B.n27 511.721
R919 B.n138 B.t10 397.743
R920 B.n52 B.t2 397.743
R921 B.n146 B.t4 397.743
R922 B.n44 B.t8 397.743
R923 B.n139 B.t11 327.923
R924 B.n53 B.t1 327.923
R925 B.n147 B.t5 327.923
R926 B.n45 B.t7 327.923
R927 B.n146 B.t3 277.784
R928 B.n138 B.t9 277.784
R929 B.n52 B.t0 277.784
R930 B.n44 B.t6 277.784
R931 B.n725 B.n724 256.663
R932 B.n724 B.n723 235.042
R933 B.n724 B.n2 235.042
R934 B.n262 B.n163 163.367
R935 B.n266 B.n163 163.367
R936 B.n267 B.n266 163.367
R937 B.n268 B.n267 163.367
R938 B.n268 B.n161 163.367
R939 B.n272 B.n161 163.367
R940 B.n273 B.n272 163.367
R941 B.n274 B.n273 163.367
R942 B.n274 B.n159 163.367
R943 B.n278 B.n159 163.367
R944 B.n279 B.n278 163.367
R945 B.n280 B.n279 163.367
R946 B.n280 B.n157 163.367
R947 B.n284 B.n157 163.367
R948 B.n285 B.n284 163.367
R949 B.n286 B.n285 163.367
R950 B.n286 B.n155 163.367
R951 B.n290 B.n155 163.367
R952 B.n291 B.n290 163.367
R953 B.n292 B.n291 163.367
R954 B.n292 B.n153 163.367
R955 B.n296 B.n153 163.367
R956 B.n297 B.n296 163.367
R957 B.n298 B.n297 163.367
R958 B.n298 B.n151 163.367
R959 B.n302 B.n151 163.367
R960 B.n303 B.n302 163.367
R961 B.n304 B.n303 163.367
R962 B.n304 B.n149 163.367
R963 B.n308 B.n149 163.367
R964 B.n309 B.n308 163.367
R965 B.n310 B.n309 163.367
R966 B.n310 B.n145 163.367
R967 B.n315 B.n145 163.367
R968 B.n316 B.n315 163.367
R969 B.n317 B.n316 163.367
R970 B.n317 B.n143 163.367
R971 B.n321 B.n143 163.367
R972 B.n322 B.n321 163.367
R973 B.n323 B.n322 163.367
R974 B.n323 B.n141 163.367
R975 B.n327 B.n141 163.367
R976 B.n328 B.n327 163.367
R977 B.n328 B.n137 163.367
R978 B.n332 B.n137 163.367
R979 B.n333 B.n332 163.367
R980 B.n334 B.n333 163.367
R981 B.n334 B.n135 163.367
R982 B.n338 B.n135 163.367
R983 B.n339 B.n338 163.367
R984 B.n340 B.n339 163.367
R985 B.n340 B.n133 163.367
R986 B.n344 B.n133 163.367
R987 B.n345 B.n344 163.367
R988 B.n346 B.n345 163.367
R989 B.n346 B.n131 163.367
R990 B.n350 B.n131 163.367
R991 B.n351 B.n350 163.367
R992 B.n352 B.n351 163.367
R993 B.n352 B.n129 163.367
R994 B.n356 B.n129 163.367
R995 B.n357 B.n356 163.367
R996 B.n358 B.n357 163.367
R997 B.n358 B.n127 163.367
R998 B.n362 B.n127 163.367
R999 B.n363 B.n362 163.367
R1000 B.n364 B.n363 163.367
R1001 B.n364 B.n125 163.367
R1002 B.n368 B.n125 163.367
R1003 B.n369 B.n368 163.367
R1004 B.n370 B.n369 163.367
R1005 B.n370 B.n123 163.367
R1006 B.n374 B.n123 163.367
R1007 B.n375 B.n374 163.367
R1008 B.n376 B.n375 163.367
R1009 B.n376 B.n121 163.367
R1010 B.n531 B.n530 163.367
R1011 B.n530 B.n71 163.367
R1012 B.n526 B.n71 163.367
R1013 B.n526 B.n525 163.367
R1014 B.n525 B.n524 163.367
R1015 B.n524 B.n73 163.367
R1016 B.n520 B.n73 163.367
R1017 B.n520 B.n519 163.367
R1018 B.n519 B.n518 163.367
R1019 B.n518 B.n75 163.367
R1020 B.n514 B.n75 163.367
R1021 B.n514 B.n513 163.367
R1022 B.n513 B.n512 163.367
R1023 B.n512 B.n77 163.367
R1024 B.n508 B.n77 163.367
R1025 B.n508 B.n507 163.367
R1026 B.n507 B.n506 163.367
R1027 B.n506 B.n79 163.367
R1028 B.n502 B.n79 163.367
R1029 B.n502 B.n501 163.367
R1030 B.n501 B.n500 163.367
R1031 B.n500 B.n81 163.367
R1032 B.n496 B.n81 163.367
R1033 B.n496 B.n495 163.367
R1034 B.n495 B.n494 163.367
R1035 B.n494 B.n83 163.367
R1036 B.n490 B.n83 163.367
R1037 B.n490 B.n489 163.367
R1038 B.n489 B.n488 163.367
R1039 B.n488 B.n85 163.367
R1040 B.n484 B.n85 163.367
R1041 B.n484 B.n483 163.367
R1042 B.n483 B.n482 163.367
R1043 B.n482 B.n87 163.367
R1044 B.n478 B.n87 163.367
R1045 B.n478 B.n477 163.367
R1046 B.n477 B.n476 163.367
R1047 B.n476 B.n89 163.367
R1048 B.n472 B.n89 163.367
R1049 B.n472 B.n471 163.367
R1050 B.n471 B.n470 163.367
R1051 B.n470 B.n91 163.367
R1052 B.n466 B.n91 163.367
R1053 B.n466 B.n465 163.367
R1054 B.n465 B.n464 163.367
R1055 B.n464 B.n93 163.367
R1056 B.n460 B.n93 163.367
R1057 B.n460 B.n459 163.367
R1058 B.n459 B.n458 163.367
R1059 B.n458 B.n95 163.367
R1060 B.n454 B.n95 163.367
R1061 B.n454 B.n453 163.367
R1062 B.n453 B.n452 163.367
R1063 B.n452 B.n97 163.367
R1064 B.n448 B.n97 163.367
R1065 B.n448 B.n447 163.367
R1066 B.n447 B.n446 163.367
R1067 B.n446 B.n99 163.367
R1068 B.n442 B.n99 163.367
R1069 B.n442 B.n441 163.367
R1070 B.n441 B.n440 163.367
R1071 B.n440 B.n101 163.367
R1072 B.n436 B.n101 163.367
R1073 B.n436 B.n435 163.367
R1074 B.n435 B.n434 163.367
R1075 B.n434 B.n103 163.367
R1076 B.n430 B.n103 163.367
R1077 B.n430 B.n429 163.367
R1078 B.n429 B.n428 163.367
R1079 B.n428 B.n105 163.367
R1080 B.n424 B.n105 163.367
R1081 B.n424 B.n423 163.367
R1082 B.n423 B.n422 163.367
R1083 B.n422 B.n107 163.367
R1084 B.n418 B.n107 163.367
R1085 B.n418 B.n417 163.367
R1086 B.n417 B.n416 163.367
R1087 B.n416 B.n109 163.367
R1088 B.n412 B.n109 163.367
R1089 B.n412 B.n411 163.367
R1090 B.n411 B.n410 163.367
R1091 B.n410 B.n111 163.367
R1092 B.n406 B.n111 163.367
R1093 B.n406 B.n405 163.367
R1094 B.n405 B.n404 163.367
R1095 B.n404 B.n113 163.367
R1096 B.n400 B.n113 163.367
R1097 B.n400 B.n399 163.367
R1098 B.n399 B.n398 163.367
R1099 B.n398 B.n115 163.367
R1100 B.n394 B.n115 163.367
R1101 B.n394 B.n393 163.367
R1102 B.n393 B.n392 163.367
R1103 B.n392 B.n117 163.367
R1104 B.n388 B.n117 163.367
R1105 B.n388 B.n387 163.367
R1106 B.n387 B.n386 163.367
R1107 B.n386 B.n119 163.367
R1108 B.n382 B.n119 163.367
R1109 B.n382 B.n381 163.367
R1110 B.n381 B.n380 163.367
R1111 B.n646 B.n27 163.367
R1112 B.n646 B.n645 163.367
R1113 B.n645 B.n644 163.367
R1114 B.n644 B.n29 163.367
R1115 B.n640 B.n29 163.367
R1116 B.n640 B.n639 163.367
R1117 B.n639 B.n638 163.367
R1118 B.n638 B.n31 163.367
R1119 B.n634 B.n31 163.367
R1120 B.n634 B.n633 163.367
R1121 B.n633 B.n632 163.367
R1122 B.n632 B.n33 163.367
R1123 B.n628 B.n33 163.367
R1124 B.n628 B.n627 163.367
R1125 B.n627 B.n626 163.367
R1126 B.n626 B.n35 163.367
R1127 B.n622 B.n35 163.367
R1128 B.n622 B.n621 163.367
R1129 B.n621 B.n620 163.367
R1130 B.n620 B.n37 163.367
R1131 B.n616 B.n37 163.367
R1132 B.n616 B.n615 163.367
R1133 B.n615 B.n614 163.367
R1134 B.n614 B.n39 163.367
R1135 B.n610 B.n39 163.367
R1136 B.n610 B.n609 163.367
R1137 B.n609 B.n608 163.367
R1138 B.n608 B.n41 163.367
R1139 B.n604 B.n41 163.367
R1140 B.n604 B.n603 163.367
R1141 B.n603 B.n602 163.367
R1142 B.n602 B.n43 163.367
R1143 B.n598 B.n43 163.367
R1144 B.n598 B.n597 163.367
R1145 B.n597 B.n47 163.367
R1146 B.n593 B.n47 163.367
R1147 B.n593 B.n592 163.367
R1148 B.n592 B.n591 163.367
R1149 B.n591 B.n49 163.367
R1150 B.n587 B.n49 163.367
R1151 B.n587 B.n586 163.367
R1152 B.n586 B.n585 163.367
R1153 B.n585 B.n51 163.367
R1154 B.n580 B.n51 163.367
R1155 B.n580 B.n579 163.367
R1156 B.n579 B.n578 163.367
R1157 B.n578 B.n55 163.367
R1158 B.n574 B.n55 163.367
R1159 B.n574 B.n573 163.367
R1160 B.n573 B.n572 163.367
R1161 B.n572 B.n57 163.367
R1162 B.n568 B.n57 163.367
R1163 B.n568 B.n567 163.367
R1164 B.n567 B.n566 163.367
R1165 B.n566 B.n59 163.367
R1166 B.n562 B.n59 163.367
R1167 B.n562 B.n561 163.367
R1168 B.n561 B.n560 163.367
R1169 B.n560 B.n61 163.367
R1170 B.n556 B.n61 163.367
R1171 B.n556 B.n555 163.367
R1172 B.n555 B.n554 163.367
R1173 B.n554 B.n63 163.367
R1174 B.n550 B.n63 163.367
R1175 B.n550 B.n549 163.367
R1176 B.n549 B.n548 163.367
R1177 B.n548 B.n65 163.367
R1178 B.n544 B.n65 163.367
R1179 B.n544 B.n543 163.367
R1180 B.n543 B.n542 163.367
R1181 B.n542 B.n67 163.367
R1182 B.n538 B.n67 163.367
R1183 B.n538 B.n537 163.367
R1184 B.n537 B.n536 163.367
R1185 B.n536 B.n69 163.367
R1186 B.n532 B.n69 163.367
R1187 B.n651 B.n650 163.367
R1188 B.n652 B.n651 163.367
R1189 B.n652 B.n25 163.367
R1190 B.n656 B.n25 163.367
R1191 B.n657 B.n656 163.367
R1192 B.n658 B.n657 163.367
R1193 B.n658 B.n23 163.367
R1194 B.n662 B.n23 163.367
R1195 B.n663 B.n662 163.367
R1196 B.n664 B.n663 163.367
R1197 B.n664 B.n21 163.367
R1198 B.n668 B.n21 163.367
R1199 B.n669 B.n668 163.367
R1200 B.n670 B.n669 163.367
R1201 B.n670 B.n19 163.367
R1202 B.n674 B.n19 163.367
R1203 B.n675 B.n674 163.367
R1204 B.n676 B.n675 163.367
R1205 B.n676 B.n17 163.367
R1206 B.n680 B.n17 163.367
R1207 B.n681 B.n680 163.367
R1208 B.n682 B.n681 163.367
R1209 B.n682 B.n15 163.367
R1210 B.n686 B.n15 163.367
R1211 B.n687 B.n686 163.367
R1212 B.n688 B.n687 163.367
R1213 B.n688 B.n13 163.367
R1214 B.n692 B.n13 163.367
R1215 B.n693 B.n692 163.367
R1216 B.n694 B.n693 163.367
R1217 B.n694 B.n11 163.367
R1218 B.n698 B.n11 163.367
R1219 B.n699 B.n698 163.367
R1220 B.n700 B.n699 163.367
R1221 B.n700 B.n9 163.367
R1222 B.n704 B.n9 163.367
R1223 B.n705 B.n704 163.367
R1224 B.n706 B.n705 163.367
R1225 B.n706 B.n7 163.367
R1226 B.n710 B.n7 163.367
R1227 B.n711 B.n710 163.367
R1228 B.n712 B.n711 163.367
R1229 B.n712 B.n5 163.367
R1230 B.n716 B.n5 163.367
R1231 B.n717 B.n716 163.367
R1232 B.n718 B.n717 163.367
R1233 B.n718 B.n3 163.367
R1234 B.n722 B.n3 163.367
R1235 B.n723 B.n722 163.367
R1236 B.n189 B.n2 163.367
R1237 B.n190 B.n189 163.367
R1238 B.n190 B.n187 163.367
R1239 B.n194 B.n187 163.367
R1240 B.n195 B.n194 163.367
R1241 B.n196 B.n195 163.367
R1242 B.n196 B.n185 163.367
R1243 B.n200 B.n185 163.367
R1244 B.n201 B.n200 163.367
R1245 B.n202 B.n201 163.367
R1246 B.n202 B.n183 163.367
R1247 B.n206 B.n183 163.367
R1248 B.n207 B.n206 163.367
R1249 B.n208 B.n207 163.367
R1250 B.n208 B.n181 163.367
R1251 B.n212 B.n181 163.367
R1252 B.n213 B.n212 163.367
R1253 B.n214 B.n213 163.367
R1254 B.n214 B.n179 163.367
R1255 B.n218 B.n179 163.367
R1256 B.n219 B.n218 163.367
R1257 B.n220 B.n219 163.367
R1258 B.n220 B.n177 163.367
R1259 B.n224 B.n177 163.367
R1260 B.n225 B.n224 163.367
R1261 B.n226 B.n225 163.367
R1262 B.n226 B.n175 163.367
R1263 B.n230 B.n175 163.367
R1264 B.n231 B.n230 163.367
R1265 B.n232 B.n231 163.367
R1266 B.n232 B.n173 163.367
R1267 B.n236 B.n173 163.367
R1268 B.n237 B.n236 163.367
R1269 B.n238 B.n237 163.367
R1270 B.n238 B.n171 163.367
R1271 B.n242 B.n171 163.367
R1272 B.n243 B.n242 163.367
R1273 B.n244 B.n243 163.367
R1274 B.n244 B.n169 163.367
R1275 B.n248 B.n169 163.367
R1276 B.n249 B.n248 163.367
R1277 B.n250 B.n249 163.367
R1278 B.n250 B.n167 163.367
R1279 B.n254 B.n167 163.367
R1280 B.n255 B.n254 163.367
R1281 B.n256 B.n255 163.367
R1282 B.n256 B.n165 163.367
R1283 B.n260 B.n165 163.367
R1284 B.n261 B.n260 163.367
R1285 B.n147 B.n146 69.8187
R1286 B.n139 B.n138 69.8187
R1287 B.n53 B.n52 69.8187
R1288 B.n45 B.n44 69.8187
R1289 B.n313 B.n147 59.5399
R1290 B.n140 B.n139 59.5399
R1291 B.n583 B.n53 59.5399
R1292 B.n46 B.n45 59.5399
R1293 B.n649 B.n648 33.2493
R1294 B.n533 B.n70 33.2493
R1295 B.n379 B.n378 33.2493
R1296 B.n263 B.n164 33.2493
R1297 B B.n725 18.0485
R1298 B.n649 B.n26 10.6151
R1299 B.n653 B.n26 10.6151
R1300 B.n654 B.n653 10.6151
R1301 B.n655 B.n654 10.6151
R1302 B.n655 B.n24 10.6151
R1303 B.n659 B.n24 10.6151
R1304 B.n660 B.n659 10.6151
R1305 B.n661 B.n660 10.6151
R1306 B.n661 B.n22 10.6151
R1307 B.n665 B.n22 10.6151
R1308 B.n666 B.n665 10.6151
R1309 B.n667 B.n666 10.6151
R1310 B.n667 B.n20 10.6151
R1311 B.n671 B.n20 10.6151
R1312 B.n672 B.n671 10.6151
R1313 B.n673 B.n672 10.6151
R1314 B.n673 B.n18 10.6151
R1315 B.n677 B.n18 10.6151
R1316 B.n678 B.n677 10.6151
R1317 B.n679 B.n678 10.6151
R1318 B.n679 B.n16 10.6151
R1319 B.n683 B.n16 10.6151
R1320 B.n684 B.n683 10.6151
R1321 B.n685 B.n684 10.6151
R1322 B.n685 B.n14 10.6151
R1323 B.n689 B.n14 10.6151
R1324 B.n690 B.n689 10.6151
R1325 B.n691 B.n690 10.6151
R1326 B.n691 B.n12 10.6151
R1327 B.n695 B.n12 10.6151
R1328 B.n696 B.n695 10.6151
R1329 B.n697 B.n696 10.6151
R1330 B.n697 B.n10 10.6151
R1331 B.n701 B.n10 10.6151
R1332 B.n702 B.n701 10.6151
R1333 B.n703 B.n702 10.6151
R1334 B.n703 B.n8 10.6151
R1335 B.n707 B.n8 10.6151
R1336 B.n708 B.n707 10.6151
R1337 B.n709 B.n708 10.6151
R1338 B.n709 B.n6 10.6151
R1339 B.n713 B.n6 10.6151
R1340 B.n714 B.n713 10.6151
R1341 B.n715 B.n714 10.6151
R1342 B.n715 B.n4 10.6151
R1343 B.n719 B.n4 10.6151
R1344 B.n720 B.n719 10.6151
R1345 B.n721 B.n720 10.6151
R1346 B.n721 B.n0 10.6151
R1347 B.n648 B.n647 10.6151
R1348 B.n647 B.n28 10.6151
R1349 B.n643 B.n28 10.6151
R1350 B.n643 B.n642 10.6151
R1351 B.n642 B.n641 10.6151
R1352 B.n641 B.n30 10.6151
R1353 B.n637 B.n30 10.6151
R1354 B.n637 B.n636 10.6151
R1355 B.n636 B.n635 10.6151
R1356 B.n635 B.n32 10.6151
R1357 B.n631 B.n32 10.6151
R1358 B.n631 B.n630 10.6151
R1359 B.n630 B.n629 10.6151
R1360 B.n629 B.n34 10.6151
R1361 B.n625 B.n34 10.6151
R1362 B.n625 B.n624 10.6151
R1363 B.n624 B.n623 10.6151
R1364 B.n623 B.n36 10.6151
R1365 B.n619 B.n36 10.6151
R1366 B.n619 B.n618 10.6151
R1367 B.n618 B.n617 10.6151
R1368 B.n617 B.n38 10.6151
R1369 B.n613 B.n38 10.6151
R1370 B.n613 B.n612 10.6151
R1371 B.n612 B.n611 10.6151
R1372 B.n611 B.n40 10.6151
R1373 B.n607 B.n40 10.6151
R1374 B.n607 B.n606 10.6151
R1375 B.n606 B.n605 10.6151
R1376 B.n605 B.n42 10.6151
R1377 B.n601 B.n42 10.6151
R1378 B.n601 B.n600 10.6151
R1379 B.n600 B.n599 10.6151
R1380 B.n596 B.n595 10.6151
R1381 B.n595 B.n594 10.6151
R1382 B.n594 B.n48 10.6151
R1383 B.n590 B.n48 10.6151
R1384 B.n590 B.n589 10.6151
R1385 B.n589 B.n588 10.6151
R1386 B.n588 B.n50 10.6151
R1387 B.n584 B.n50 10.6151
R1388 B.n582 B.n581 10.6151
R1389 B.n581 B.n54 10.6151
R1390 B.n577 B.n54 10.6151
R1391 B.n577 B.n576 10.6151
R1392 B.n576 B.n575 10.6151
R1393 B.n575 B.n56 10.6151
R1394 B.n571 B.n56 10.6151
R1395 B.n571 B.n570 10.6151
R1396 B.n570 B.n569 10.6151
R1397 B.n569 B.n58 10.6151
R1398 B.n565 B.n58 10.6151
R1399 B.n565 B.n564 10.6151
R1400 B.n564 B.n563 10.6151
R1401 B.n563 B.n60 10.6151
R1402 B.n559 B.n60 10.6151
R1403 B.n559 B.n558 10.6151
R1404 B.n558 B.n557 10.6151
R1405 B.n557 B.n62 10.6151
R1406 B.n553 B.n62 10.6151
R1407 B.n553 B.n552 10.6151
R1408 B.n552 B.n551 10.6151
R1409 B.n551 B.n64 10.6151
R1410 B.n547 B.n64 10.6151
R1411 B.n547 B.n546 10.6151
R1412 B.n546 B.n545 10.6151
R1413 B.n545 B.n66 10.6151
R1414 B.n541 B.n66 10.6151
R1415 B.n541 B.n540 10.6151
R1416 B.n540 B.n539 10.6151
R1417 B.n539 B.n68 10.6151
R1418 B.n535 B.n68 10.6151
R1419 B.n535 B.n534 10.6151
R1420 B.n534 B.n533 10.6151
R1421 B.n529 B.n70 10.6151
R1422 B.n529 B.n528 10.6151
R1423 B.n528 B.n527 10.6151
R1424 B.n527 B.n72 10.6151
R1425 B.n523 B.n72 10.6151
R1426 B.n523 B.n522 10.6151
R1427 B.n522 B.n521 10.6151
R1428 B.n521 B.n74 10.6151
R1429 B.n517 B.n74 10.6151
R1430 B.n517 B.n516 10.6151
R1431 B.n516 B.n515 10.6151
R1432 B.n515 B.n76 10.6151
R1433 B.n511 B.n76 10.6151
R1434 B.n511 B.n510 10.6151
R1435 B.n510 B.n509 10.6151
R1436 B.n509 B.n78 10.6151
R1437 B.n505 B.n78 10.6151
R1438 B.n505 B.n504 10.6151
R1439 B.n504 B.n503 10.6151
R1440 B.n503 B.n80 10.6151
R1441 B.n499 B.n80 10.6151
R1442 B.n499 B.n498 10.6151
R1443 B.n498 B.n497 10.6151
R1444 B.n497 B.n82 10.6151
R1445 B.n493 B.n82 10.6151
R1446 B.n493 B.n492 10.6151
R1447 B.n492 B.n491 10.6151
R1448 B.n491 B.n84 10.6151
R1449 B.n487 B.n84 10.6151
R1450 B.n487 B.n486 10.6151
R1451 B.n486 B.n485 10.6151
R1452 B.n485 B.n86 10.6151
R1453 B.n481 B.n86 10.6151
R1454 B.n481 B.n480 10.6151
R1455 B.n480 B.n479 10.6151
R1456 B.n479 B.n88 10.6151
R1457 B.n475 B.n88 10.6151
R1458 B.n475 B.n474 10.6151
R1459 B.n474 B.n473 10.6151
R1460 B.n473 B.n90 10.6151
R1461 B.n469 B.n90 10.6151
R1462 B.n469 B.n468 10.6151
R1463 B.n468 B.n467 10.6151
R1464 B.n467 B.n92 10.6151
R1465 B.n463 B.n92 10.6151
R1466 B.n463 B.n462 10.6151
R1467 B.n462 B.n461 10.6151
R1468 B.n461 B.n94 10.6151
R1469 B.n457 B.n94 10.6151
R1470 B.n457 B.n456 10.6151
R1471 B.n456 B.n455 10.6151
R1472 B.n455 B.n96 10.6151
R1473 B.n451 B.n96 10.6151
R1474 B.n451 B.n450 10.6151
R1475 B.n450 B.n449 10.6151
R1476 B.n449 B.n98 10.6151
R1477 B.n445 B.n98 10.6151
R1478 B.n445 B.n444 10.6151
R1479 B.n444 B.n443 10.6151
R1480 B.n443 B.n100 10.6151
R1481 B.n439 B.n100 10.6151
R1482 B.n439 B.n438 10.6151
R1483 B.n438 B.n437 10.6151
R1484 B.n437 B.n102 10.6151
R1485 B.n433 B.n102 10.6151
R1486 B.n433 B.n432 10.6151
R1487 B.n432 B.n431 10.6151
R1488 B.n431 B.n104 10.6151
R1489 B.n427 B.n104 10.6151
R1490 B.n427 B.n426 10.6151
R1491 B.n426 B.n425 10.6151
R1492 B.n425 B.n106 10.6151
R1493 B.n421 B.n106 10.6151
R1494 B.n421 B.n420 10.6151
R1495 B.n420 B.n419 10.6151
R1496 B.n419 B.n108 10.6151
R1497 B.n415 B.n108 10.6151
R1498 B.n415 B.n414 10.6151
R1499 B.n414 B.n413 10.6151
R1500 B.n413 B.n110 10.6151
R1501 B.n409 B.n110 10.6151
R1502 B.n409 B.n408 10.6151
R1503 B.n408 B.n407 10.6151
R1504 B.n407 B.n112 10.6151
R1505 B.n403 B.n112 10.6151
R1506 B.n403 B.n402 10.6151
R1507 B.n402 B.n401 10.6151
R1508 B.n401 B.n114 10.6151
R1509 B.n397 B.n114 10.6151
R1510 B.n397 B.n396 10.6151
R1511 B.n396 B.n395 10.6151
R1512 B.n395 B.n116 10.6151
R1513 B.n391 B.n116 10.6151
R1514 B.n391 B.n390 10.6151
R1515 B.n390 B.n389 10.6151
R1516 B.n389 B.n118 10.6151
R1517 B.n385 B.n118 10.6151
R1518 B.n385 B.n384 10.6151
R1519 B.n384 B.n383 10.6151
R1520 B.n383 B.n120 10.6151
R1521 B.n379 B.n120 10.6151
R1522 B.n188 B.n1 10.6151
R1523 B.n191 B.n188 10.6151
R1524 B.n192 B.n191 10.6151
R1525 B.n193 B.n192 10.6151
R1526 B.n193 B.n186 10.6151
R1527 B.n197 B.n186 10.6151
R1528 B.n198 B.n197 10.6151
R1529 B.n199 B.n198 10.6151
R1530 B.n199 B.n184 10.6151
R1531 B.n203 B.n184 10.6151
R1532 B.n204 B.n203 10.6151
R1533 B.n205 B.n204 10.6151
R1534 B.n205 B.n182 10.6151
R1535 B.n209 B.n182 10.6151
R1536 B.n210 B.n209 10.6151
R1537 B.n211 B.n210 10.6151
R1538 B.n211 B.n180 10.6151
R1539 B.n215 B.n180 10.6151
R1540 B.n216 B.n215 10.6151
R1541 B.n217 B.n216 10.6151
R1542 B.n217 B.n178 10.6151
R1543 B.n221 B.n178 10.6151
R1544 B.n222 B.n221 10.6151
R1545 B.n223 B.n222 10.6151
R1546 B.n223 B.n176 10.6151
R1547 B.n227 B.n176 10.6151
R1548 B.n228 B.n227 10.6151
R1549 B.n229 B.n228 10.6151
R1550 B.n229 B.n174 10.6151
R1551 B.n233 B.n174 10.6151
R1552 B.n234 B.n233 10.6151
R1553 B.n235 B.n234 10.6151
R1554 B.n235 B.n172 10.6151
R1555 B.n239 B.n172 10.6151
R1556 B.n240 B.n239 10.6151
R1557 B.n241 B.n240 10.6151
R1558 B.n241 B.n170 10.6151
R1559 B.n245 B.n170 10.6151
R1560 B.n246 B.n245 10.6151
R1561 B.n247 B.n246 10.6151
R1562 B.n247 B.n168 10.6151
R1563 B.n251 B.n168 10.6151
R1564 B.n252 B.n251 10.6151
R1565 B.n253 B.n252 10.6151
R1566 B.n253 B.n166 10.6151
R1567 B.n257 B.n166 10.6151
R1568 B.n258 B.n257 10.6151
R1569 B.n259 B.n258 10.6151
R1570 B.n259 B.n164 10.6151
R1571 B.n264 B.n263 10.6151
R1572 B.n265 B.n264 10.6151
R1573 B.n265 B.n162 10.6151
R1574 B.n269 B.n162 10.6151
R1575 B.n270 B.n269 10.6151
R1576 B.n271 B.n270 10.6151
R1577 B.n271 B.n160 10.6151
R1578 B.n275 B.n160 10.6151
R1579 B.n276 B.n275 10.6151
R1580 B.n277 B.n276 10.6151
R1581 B.n277 B.n158 10.6151
R1582 B.n281 B.n158 10.6151
R1583 B.n282 B.n281 10.6151
R1584 B.n283 B.n282 10.6151
R1585 B.n283 B.n156 10.6151
R1586 B.n287 B.n156 10.6151
R1587 B.n288 B.n287 10.6151
R1588 B.n289 B.n288 10.6151
R1589 B.n289 B.n154 10.6151
R1590 B.n293 B.n154 10.6151
R1591 B.n294 B.n293 10.6151
R1592 B.n295 B.n294 10.6151
R1593 B.n295 B.n152 10.6151
R1594 B.n299 B.n152 10.6151
R1595 B.n300 B.n299 10.6151
R1596 B.n301 B.n300 10.6151
R1597 B.n301 B.n150 10.6151
R1598 B.n305 B.n150 10.6151
R1599 B.n306 B.n305 10.6151
R1600 B.n307 B.n306 10.6151
R1601 B.n307 B.n148 10.6151
R1602 B.n311 B.n148 10.6151
R1603 B.n312 B.n311 10.6151
R1604 B.n314 B.n144 10.6151
R1605 B.n318 B.n144 10.6151
R1606 B.n319 B.n318 10.6151
R1607 B.n320 B.n319 10.6151
R1608 B.n320 B.n142 10.6151
R1609 B.n324 B.n142 10.6151
R1610 B.n325 B.n324 10.6151
R1611 B.n326 B.n325 10.6151
R1612 B.n330 B.n329 10.6151
R1613 B.n331 B.n330 10.6151
R1614 B.n331 B.n136 10.6151
R1615 B.n335 B.n136 10.6151
R1616 B.n336 B.n335 10.6151
R1617 B.n337 B.n336 10.6151
R1618 B.n337 B.n134 10.6151
R1619 B.n341 B.n134 10.6151
R1620 B.n342 B.n341 10.6151
R1621 B.n343 B.n342 10.6151
R1622 B.n343 B.n132 10.6151
R1623 B.n347 B.n132 10.6151
R1624 B.n348 B.n347 10.6151
R1625 B.n349 B.n348 10.6151
R1626 B.n349 B.n130 10.6151
R1627 B.n353 B.n130 10.6151
R1628 B.n354 B.n353 10.6151
R1629 B.n355 B.n354 10.6151
R1630 B.n355 B.n128 10.6151
R1631 B.n359 B.n128 10.6151
R1632 B.n360 B.n359 10.6151
R1633 B.n361 B.n360 10.6151
R1634 B.n361 B.n126 10.6151
R1635 B.n365 B.n126 10.6151
R1636 B.n366 B.n365 10.6151
R1637 B.n367 B.n366 10.6151
R1638 B.n367 B.n124 10.6151
R1639 B.n371 B.n124 10.6151
R1640 B.n372 B.n371 10.6151
R1641 B.n373 B.n372 10.6151
R1642 B.n373 B.n122 10.6151
R1643 B.n377 B.n122 10.6151
R1644 B.n378 B.n377 10.6151
R1645 B.n725 B.n0 8.11757
R1646 B.n725 B.n1 8.11757
R1647 B.n596 B.n46 6.5566
R1648 B.n584 B.n583 6.5566
R1649 B.n314 B.n313 6.5566
R1650 B.n326 B.n140 6.5566
R1651 B.n599 B.n46 4.05904
R1652 B.n583 B.n582 4.05904
R1653 B.n313 B.n312 4.05904
R1654 B.n329 B.n140 4.05904
R1655 VN.n34 VN.n33 161.3
R1656 VN.n32 VN.n19 161.3
R1657 VN.n31 VN.n30 161.3
R1658 VN.n29 VN.n20 161.3
R1659 VN.n28 VN.n27 161.3
R1660 VN.n26 VN.n21 161.3
R1661 VN.n25 VN.n24 161.3
R1662 VN.n16 VN.n15 161.3
R1663 VN.n14 VN.n1 161.3
R1664 VN.n13 VN.n12 161.3
R1665 VN.n11 VN.n2 161.3
R1666 VN.n10 VN.n9 161.3
R1667 VN.n8 VN.n3 161.3
R1668 VN.n7 VN.n6 161.3
R1669 VN.n23 VN.t1 102.091
R1670 VN.n5 VN.t3 102.091
R1671 VN.n17 VN.n0 72.9405
R1672 VN.n35 VN.n18 72.9405
R1673 VN.n4 VN.t4 68.9103
R1674 VN.n0 VN.t2 68.9103
R1675 VN.n22 VN.t5 68.9103
R1676 VN.n18 VN.t0 68.9103
R1677 VN.n5 VN.n4 62.0536
R1678 VN.n23 VN.n22 62.0536
R1679 VN VN.n35 49.6041
R1680 VN.n13 VN.n2 45.3497
R1681 VN.n31 VN.n20 45.3497
R1682 VN.n9 VN.n2 35.6371
R1683 VN.n27 VN.n20 35.6371
R1684 VN.n8 VN.n7 24.4675
R1685 VN.n9 VN.n8 24.4675
R1686 VN.n14 VN.n13 24.4675
R1687 VN.n15 VN.n14 24.4675
R1688 VN.n27 VN.n26 24.4675
R1689 VN.n26 VN.n25 24.4675
R1690 VN.n33 VN.n32 24.4675
R1691 VN.n32 VN.n31 24.4675
R1692 VN.n15 VN.n0 17.1274
R1693 VN.n33 VN.n18 17.1274
R1694 VN.n7 VN.n4 12.234
R1695 VN.n25 VN.n22 12.234
R1696 VN.n24 VN.n23 4.04081
R1697 VN.n6 VN.n5 4.04081
R1698 VN.n35 VN.n34 0.354971
R1699 VN.n17 VN.n16 0.354971
R1700 VN VN.n17 0.26696
R1701 VN.n34 VN.n19 0.189894
R1702 VN.n30 VN.n19 0.189894
R1703 VN.n30 VN.n29 0.189894
R1704 VN.n29 VN.n28 0.189894
R1705 VN.n28 VN.n21 0.189894
R1706 VN.n24 VN.n21 0.189894
R1707 VN.n6 VN.n3 0.189894
R1708 VN.n10 VN.n3 0.189894
R1709 VN.n11 VN.n10 0.189894
R1710 VN.n12 VN.n11 0.189894
R1711 VN.n12 VN.n1 0.189894
R1712 VN.n16 VN.n1 0.189894
R1713 VDD2.n95 VDD2.n51 756.745
R1714 VDD2.n44 VDD2.n0 756.745
R1715 VDD2.n96 VDD2.n95 585
R1716 VDD2.n94 VDD2.n93 585
R1717 VDD2.n55 VDD2.n54 585
R1718 VDD2.n59 VDD2.n57 585
R1719 VDD2.n88 VDD2.n87 585
R1720 VDD2.n86 VDD2.n85 585
R1721 VDD2.n61 VDD2.n60 585
R1722 VDD2.n80 VDD2.n79 585
R1723 VDD2.n78 VDD2.n77 585
R1724 VDD2.n65 VDD2.n64 585
R1725 VDD2.n72 VDD2.n71 585
R1726 VDD2.n70 VDD2.n69 585
R1727 VDD2.n17 VDD2.n16 585
R1728 VDD2.n19 VDD2.n18 585
R1729 VDD2.n12 VDD2.n11 585
R1730 VDD2.n25 VDD2.n24 585
R1731 VDD2.n27 VDD2.n26 585
R1732 VDD2.n8 VDD2.n7 585
R1733 VDD2.n34 VDD2.n33 585
R1734 VDD2.n35 VDD2.n6 585
R1735 VDD2.n37 VDD2.n36 585
R1736 VDD2.n4 VDD2.n3 585
R1737 VDD2.n43 VDD2.n42 585
R1738 VDD2.n45 VDD2.n44 585
R1739 VDD2.n68 VDD2.t5 329.038
R1740 VDD2.n15 VDD2.t2 329.038
R1741 VDD2.n95 VDD2.n94 171.744
R1742 VDD2.n94 VDD2.n54 171.744
R1743 VDD2.n59 VDD2.n54 171.744
R1744 VDD2.n87 VDD2.n59 171.744
R1745 VDD2.n87 VDD2.n86 171.744
R1746 VDD2.n86 VDD2.n60 171.744
R1747 VDD2.n79 VDD2.n60 171.744
R1748 VDD2.n79 VDD2.n78 171.744
R1749 VDD2.n78 VDD2.n64 171.744
R1750 VDD2.n71 VDD2.n64 171.744
R1751 VDD2.n71 VDD2.n70 171.744
R1752 VDD2.n18 VDD2.n17 171.744
R1753 VDD2.n18 VDD2.n11 171.744
R1754 VDD2.n25 VDD2.n11 171.744
R1755 VDD2.n26 VDD2.n25 171.744
R1756 VDD2.n26 VDD2.n7 171.744
R1757 VDD2.n34 VDD2.n7 171.744
R1758 VDD2.n35 VDD2.n34 171.744
R1759 VDD2.n36 VDD2.n35 171.744
R1760 VDD2.n36 VDD2.n3 171.744
R1761 VDD2.n43 VDD2.n3 171.744
R1762 VDD2.n44 VDD2.n43 171.744
R1763 VDD2.n70 VDD2.t5 85.8723
R1764 VDD2.n17 VDD2.t2 85.8723
R1765 VDD2.n50 VDD2.n49 81.4346
R1766 VDD2 VDD2.n101 81.4317
R1767 VDD2.n50 VDD2.n48 53.2697
R1768 VDD2.n100 VDD2.n99 50.9975
R1769 VDD2.n100 VDD2.n50 41.8618
R1770 VDD2.n57 VDD2.n55 13.1884
R1771 VDD2.n37 VDD2.n4 13.1884
R1772 VDD2.n93 VDD2.n92 12.8005
R1773 VDD2.n89 VDD2.n88 12.8005
R1774 VDD2.n38 VDD2.n6 12.8005
R1775 VDD2.n42 VDD2.n41 12.8005
R1776 VDD2.n96 VDD2.n53 12.0247
R1777 VDD2.n85 VDD2.n58 12.0247
R1778 VDD2.n33 VDD2.n32 12.0247
R1779 VDD2.n45 VDD2.n2 12.0247
R1780 VDD2.n97 VDD2.n51 11.249
R1781 VDD2.n84 VDD2.n61 11.249
R1782 VDD2.n31 VDD2.n8 11.249
R1783 VDD2.n46 VDD2.n0 11.249
R1784 VDD2.n69 VDD2.n68 10.7239
R1785 VDD2.n16 VDD2.n15 10.7239
R1786 VDD2.n81 VDD2.n80 10.4732
R1787 VDD2.n28 VDD2.n27 10.4732
R1788 VDD2.n77 VDD2.n63 9.69747
R1789 VDD2.n24 VDD2.n10 9.69747
R1790 VDD2.n99 VDD2.n98 9.45567
R1791 VDD2.n48 VDD2.n47 9.45567
R1792 VDD2.n67 VDD2.n66 9.3005
R1793 VDD2.n74 VDD2.n73 9.3005
R1794 VDD2.n76 VDD2.n75 9.3005
R1795 VDD2.n63 VDD2.n62 9.3005
R1796 VDD2.n82 VDD2.n81 9.3005
R1797 VDD2.n84 VDD2.n83 9.3005
R1798 VDD2.n58 VDD2.n56 9.3005
R1799 VDD2.n90 VDD2.n89 9.3005
R1800 VDD2.n98 VDD2.n97 9.3005
R1801 VDD2.n53 VDD2.n52 9.3005
R1802 VDD2.n92 VDD2.n91 9.3005
R1803 VDD2.n47 VDD2.n46 9.3005
R1804 VDD2.n2 VDD2.n1 9.3005
R1805 VDD2.n41 VDD2.n40 9.3005
R1806 VDD2.n14 VDD2.n13 9.3005
R1807 VDD2.n21 VDD2.n20 9.3005
R1808 VDD2.n23 VDD2.n22 9.3005
R1809 VDD2.n10 VDD2.n9 9.3005
R1810 VDD2.n29 VDD2.n28 9.3005
R1811 VDD2.n31 VDD2.n30 9.3005
R1812 VDD2.n32 VDD2.n5 9.3005
R1813 VDD2.n39 VDD2.n38 9.3005
R1814 VDD2.n76 VDD2.n65 8.92171
R1815 VDD2.n23 VDD2.n12 8.92171
R1816 VDD2.n73 VDD2.n72 8.14595
R1817 VDD2.n20 VDD2.n19 8.14595
R1818 VDD2.n69 VDD2.n67 7.3702
R1819 VDD2.n16 VDD2.n14 7.3702
R1820 VDD2.n72 VDD2.n67 5.81868
R1821 VDD2.n19 VDD2.n14 5.81868
R1822 VDD2.n73 VDD2.n65 5.04292
R1823 VDD2.n20 VDD2.n12 5.04292
R1824 VDD2.n77 VDD2.n76 4.26717
R1825 VDD2.n24 VDD2.n23 4.26717
R1826 VDD2.n80 VDD2.n63 3.49141
R1827 VDD2.n27 VDD2.n10 3.49141
R1828 VDD2.n101 VDD2.t0 3.47697
R1829 VDD2.n101 VDD2.t4 3.47697
R1830 VDD2.n49 VDD2.t1 3.47697
R1831 VDD2.n49 VDD2.t3 3.47697
R1832 VDD2.n99 VDD2.n51 2.71565
R1833 VDD2.n81 VDD2.n61 2.71565
R1834 VDD2.n28 VDD2.n8 2.71565
R1835 VDD2.n48 VDD2.n0 2.71565
R1836 VDD2.n68 VDD2.n66 2.41283
R1837 VDD2.n15 VDD2.n13 2.41283
R1838 VDD2 VDD2.n100 2.38628
R1839 VDD2.n97 VDD2.n96 1.93989
R1840 VDD2.n85 VDD2.n84 1.93989
R1841 VDD2.n33 VDD2.n31 1.93989
R1842 VDD2.n46 VDD2.n45 1.93989
R1843 VDD2.n93 VDD2.n53 1.16414
R1844 VDD2.n88 VDD2.n58 1.16414
R1845 VDD2.n32 VDD2.n6 1.16414
R1846 VDD2.n42 VDD2.n2 1.16414
R1847 VDD2.n92 VDD2.n55 0.388379
R1848 VDD2.n89 VDD2.n57 0.388379
R1849 VDD2.n38 VDD2.n37 0.388379
R1850 VDD2.n41 VDD2.n4 0.388379
R1851 VDD2.n98 VDD2.n52 0.155672
R1852 VDD2.n91 VDD2.n52 0.155672
R1853 VDD2.n91 VDD2.n90 0.155672
R1854 VDD2.n90 VDD2.n56 0.155672
R1855 VDD2.n83 VDD2.n56 0.155672
R1856 VDD2.n83 VDD2.n82 0.155672
R1857 VDD2.n82 VDD2.n62 0.155672
R1858 VDD2.n75 VDD2.n62 0.155672
R1859 VDD2.n75 VDD2.n74 0.155672
R1860 VDD2.n74 VDD2.n66 0.155672
R1861 VDD2.n21 VDD2.n13 0.155672
R1862 VDD2.n22 VDD2.n21 0.155672
R1863 VDD2.n22 VDD2.n9 0.155672
R1864 VDD2.n29 VDD2.n9 0.155672
R1865 VDD2.n30 VDD2.n29 0.155672
R1866 VDD2.n30 VDD2.n5 0.155672
R1867 VDD2.n39 VDD2.n5 0.155672
R1868 VDD2.n40 VDD2.n39 0.155672
R1869 VDD2.n40 VDD2.n1 0.155672
R1870 VDD2.n47 VDD2.n1 0.155672
C0 VDD2 VDD1 1.66723f
C1 VDD2 VTAIL 7.0965f
C2 w_n3850_n2838# B 9.85847f
C3 VP VN 7.08694f
C4 VDD1 w_n3850_n2838# 2.26993f
C5 w_n3850_n2838# VTAIL 2.6665f
C6 VP B 2.115f
C7 VN B 1.27746f
C8 VDD1 VP 5.89938f
C9 VP VTAIL 5.9964f
C10 VDD1 VN 0.151534f
C11 VDD2 w_n3850_n2838# 2.37641f
C12 VN VTAIL 5.98219f
C13 VDD1 B 2.05576f
C14 VTAIL B 3.33379f
C15 VDD2 VP 0.514834f
C16 VDD2 VN 5.53877f
C17 VDD1 VTAIL 7.04008f
C18 VP w_n3850_n2838# 7.90707f
C19 VN w_n3850_n2838# 7.407451f
C20 VDD2 B 2.14592f
C21 VDD2 VSUBS 2.008884f
C22 VDD1 VSUBS 2.004393f
C23 VTAIL VSUBS 1.230729f
C24 VN VSUBS 6.43372f
C25 VP VSUBS 3.371769f
C26 B VSUBS 5.077041f
C27 w_n3850_n2838# VSUBS 0.135135p
C28 VDD2.n0 VSUBS 0.031266f
C29 VDD2.n1 VSUBS 0.029128f
C30 VDD2.n2 VSUBS 0.015652f
C31 VDD2.n3 VSUBS 0.036995f
C32 VDD2.n4 VSUBS 0.016112f
C33 VDD2.n5 VSUBS 0.029128f
C34 VDD2.n6 VSUBS 0.016573f
C35 VDD2.n7 VSUBS 0.036995f
C36 VDD2.n8 VSUBS 0.016573f
C37 VDD2.n9 VSUBS 0.029128f
C38 VDD2.n10 VSUBS 0.015652f
C39 VDD2.n11 VSUBS 0.036995f
C40 VDD2.n12 VSUBS 0.016573f
C41 VDD2.n13 VSUBS 1.09283f
C42 VDD2.n14 VSUBS 0.015652f
C43 VDD2.t2 VSUBS 0.079506f
C44 VDD2.n15 VSUBS 0.194534f
C45 VDD2.n16 VSUBS 0.02783f
C46 VDD2.n17 VSUBS 0.027746f
C47 VDD2.n18 VSUBS 0.036995f
C48 VDD2.n19 VSUBS 0.016573f
C49 VDD2.n20 VSUBS 0.015652f
C50 VDD2.n21 VSUBS 0.029128f
C51 VDD2.n22 VSUBS 0.029128f
C52 VDD2.n23 VSUBS 0.015652f
C53 VDD2.n24 VSUBS 0.016573f
C54 VDD2.n25 VSUBS 0.036995f
C55 VDD2.n26 VSUBS 0.036995f
C56 VDD2.n27 VSUBS 0.016573f
C57 VDD2.n28 VSUBS 0.015652f
C58 VDD2.n29 VSUBS 0.029128f
C59 VDD2.n30 VSUBS 0.029128f
C60 VDD2.n31 VSUBS 0.015652f
C61 VDD2.n32 VSUBS 0.015652f
C62 VDD2.n33 VSUBS 0.016573f
C63 VDD2.n34 VSUBS 0.036995f
C64 VDD2.n35 VSUBS 0.036995f
C65 VDD2.n36 VSUBS 0.036995f
C66 VDD2.n37 VSUBS 0.016112f
C67 VDD2.n38 VSUBS 0.015652f
C68 VDD2.n39 VSUBS 0.029128f
C69 VDD2.n40 VSUBS 0.029128f
C70 VDD2.n41 VSUBS 0.015652f
C71 VDD2.n42 VSUBS 0.016573f
C72 VDD2.n43 VSUBS 0.036995f
C73 VDD2.n44 VSUBS 0.087044f
C74 VDD2.n45 VSUBS 0.016573f
C75 VDD2.n46 VSUBS 0.015652f
C76 VDD2.n47 VSUBS 0.071704f
C77 VDD2.n48 VSUBS 0.075481f
C78 VDD2.t1 VSUBS 0.215213f
C79 VDD2.t3 VSUBS 0.215213f
C80 VDD2.n49 VSUBS 1.61803f
C81 VDD2.n50 VSUBS 3.54089f
C82 VDD2.n51 VSUBS 0.031266f
C83 VDD2.n52 VSUBS 0.029128f
C84 VDD2.n53 VSUBS 0.015652f
C85 VDD2.n54 VSUBS 0.036995f
C86 VDD2.n55 VSUBS 0.016112f
C87 VDD2.n56 VSUBS 0.029128f
C88 VDD2.n57 VSUBS 0.016112f
C89 VDD2.n58 VSUBS 0.015652f
C90 VDD2.n59 VSUBS 0.036995f
C91 VDD2.n60 VSUBS 0.036995f
C92 VDD2.n61 VSUBS 0.016573f
C93 VDD2.n62 VSUBS 0.029128f
C94 VDD2.n63 VSUBS 0.015652f
C95 VDD2.n64 VSUBS 0.036995f
C96 VDD2.n65 VSUBS 0.016573f
C97 VDD2.n66 VSUBS 1.09283f
C98 VDD2.n67 VSUBS 0.015652f
C99 VDD2.t5 VSUBS 0.079506f
C100 VDD2.n68 VSUBS 0.194534f
C101 VDD2.n69 VSUBS 0.02783f
C102 VDD2.n70 VSUBS 0.027746f
C103 VDD2.n71 VSUBS 0.036995f
C104 VDD2.n72 VSUBS 0.016573f
C105 VDD2.n73 VSUBS 0.015652f
C106 VDD2.n74 VSUBS 0.029128f
C107 VDD2.n75 VSUBS 0.029128f
C108 VDD2.n76 VSUBS 0.015652f
C109 VDD2.n77 VSUBS 0.016573f
C110 VDD2.n78 VSUBS 0.036995f
C111 VDD2.n79 VSUBS 0.036995f
C112 VDD2.n80 VSUBS 0.016573f
C113 VDD2.n81 VSUBS 0.015652f
C114 VDD2.n82 VSUBS 0.029128f
C115 VDD2.n83 VSUBS 0.029128f
C116 VDD2.n84 VSUBS 0.015652f
C117 VDD2.n85 VSUBS 0.016573f
C118 VDD2.n86 VSUBS 0.036995f
C119 VDD2.n87 VSUBS 0.036995f
C120 VDD2.n88 VSUBS 0.016573f
C121 VDD2.n89 VSUBS 0.015652f
C122 VDD2.n90 VSUBS 0.029128f
C123 VDD2.n91 VSUBS 0.029128f
C124 VDD2.n92 VSUBS 0.015652f
C125 VDD2.n93 VSUBS 0.016573f
C126 VDD2.n94 VSUBS 0.036995f
C127 VDD2.n95 VSUBS 0.087044f
C128 VDD2.n96 VSUBS 0.016573f
C129 VDD2.n97 VSUBS 0.015652f
C130 VDD2.n98 VSUBS 0.071704f
C131 VDD2.n99 VSUBS 0.063872f
C132 VDD2.n100 VSUBS 2.96113f
C133 VDD2.t0 VSUBS 0.215213f
C134 VDD2.t4 VSUBS 0.215213f
C135 VDD2.n101 VSUBS 1.61799f
C136 VN.t2 VSUBS 2.41897f
C137 VN.n0 VSUBS 0.982012f
C138 VN.n1 VSUBS 0.029275f
C139 VN.n2 VSUBS 0.02462f
C140 VN.n3 VSUBS 0.029275f
C141 VN.t4 VSUBS 2.41897f
C142 VN.n4 VSUBS 0.960321f
C143 VN.t3 VSUBS 2.76814f
C144 VN.n5 VSUBS 0.91248f
C145 VN.n6 VSUBS 0.341557f
C146 VN.n7 VSUBS 0.041093f
C147 VN.n8 VSUBS 0.054561f
C148 VN.n9 VSUBS 0.059118f
C149 VN.n10 VSUBS 0.029275f
C150 VN.n11 VSUBS 0.029275f
C151 VN.n12 VSUBS 0.029275f
C152 VN.n13 VSUBS 0.056295f
C153 VN.n14 VSUBS 0.054561f
C154 VN.n15 VSUBS 0.04648f
C155 VN.n16 VSUBS 0.047249f
C156 VN.n17 VSUBS 0.067472f
C157 VN.t0 VSUBS 2.41897f
C158 VN.n18 VSUBS 0.982012f
C159 VN.n19 VSUBS 0.029275f
C160 VN.n20 VSUBS 0.02462f
C161 VN.n21 VSUBS 0.029275f
C162 VN.t5 VSUBS 2.41897f
C163 VN.n22 VSUBS 0.960321f
C164 VN.t1 VSUBS 2.76814f
C165 VN.n23 VSUBS 0.91248f
C166 VN.n24 VSUBS 0.341557f
C167 VN.n25 VSUBS 0.041093f
C168 VN.n26 VSUBS 0.054561f
C169 VN.n27 VSUBS 0.059118f
C170 VN.n28 VSUBS 0.029275f
C171 VN.n29 VSUBS 0.029275f
C172 VN.n30 VSUBS 0.029275f
C173 VN.n31 VSUBS 0.056295f
C174 VN.n32 VSUBS 0.054561f
C175 VN.n33 VSUBS 0.04648f
C176 VN.n34 VSUBS 0.047249f
C177 VN.n35 VSUBS 1.648f
C178 B.n0 VSUBS 0.008347f
C179 B.n1 VSUBS 0.008347f
C180 B.n2 VSUBS 0.012344f
C181 B.n3 VSUBS 0.00946f
C182 B.n4 VSUBS 0.00946f
C183 B.n5 VSUBS 0.00946f
C184 B.n6 VSUBS 0.00946f
C185 B.n7 VSUBS 0.00946f
C186 B.n8 VSUBS 0.00946f
C187 B.n9 VSUBS 0.00946f
C188 B.n10 VSUBS 0.00946f
C189 B.n11 VSUBS 0.00946f
C190 B.n12 VSUBS 0.00946f
C191 B.n13 VSUBS 0.00946f
C192 B.n14 VSUBS 0.00946f
C193 B.n15 VSUBS 0.00946f
C194 B.n16 VSUBS 0.00946f
C195 B.n17 VSUBS 0.00946f
C196 B.n18 VSUBS 0.00946f
C197 B.n19 VSUBS 0.00946f
C198 B.n20 VSUBS 0.00946f
C199 B.n21 VSUBS 0.00946f
C200 B.n22 VSUBS 0.00946f
C201 B.n23 VSUBS 0.00946f
C202 B.n24 VSUBS 0.00946f
C203 B.n25 VSUBS 0.00946f
C204 B.n26 VSUBS 0.00946f
C205 B.n27 VSUBS 0.022785f
C206 B.n28 VSUBS 0.00946f
C207 B.n29 VSUBS 0.00946f
C208 B.n30 VSUBS 0.00946f
C209 B.n31 VSUBS 0.00946f
C210 B.n32 VSUBS 0.00946f
C211 B.n33 VSUBS 0.00946f
C212 B.n34 VSUBS 0.00946f
C213 B.n35 VSUBS 0.00946f
C214 B.n36 VSUBS 0.00946f
C215 B.n37 VSUBS 0.00946f
C216 B.n38 VSUBS 0.00946f
C217 B.n39 VSUBS 0.00946f
C218 B.n40 VSUBS 0.00946f
C219 B.n41 VSUBS 0.00946f
C220 B.n42 VSUBS 0.00946f
C221 B.n43 VSUBS 0.00946f
C222 B.t7 VSUBS 0.208001f
C223 B.t8 VSUBS 0.256849f
C224 B.t6 VSUBS 1.93559f
C225 B.n44 VSUBS 0.416325f
C226 B.n45 VSUBS 0.291773f
C227 B.n46 VSUBS 0.021917f
C228 B.n47 VSUBS 0.00946f
C229 B.n48 VSUBS 0.00946f
C230 B.n49 VSUBS 0.00946f
C231 B.n50 VSUBS 0.00946f
C232 B.n51 VSUBS 0.00946f
C233 B.t1 VSUBS 0.208004f
C234 B.t2 VSUBS 0.256852f
C235 B.t0 VSUBS 1.93559f
C236 B.n52 VSUBS 0.416322f
C237 B.n53 VSUBS 0.291769f
C238 B.n54 VSUBS 0.00946f
C239 B.n55 VSUBS 0.00946f
C240 B.n56 VSUBS 0.00946f
C241 B.n57 VSUBS 0.00946f
C242 B.n58 VSUBS 0.00946f
C243 B.n59 VSUBS 0.00946f
C244 B.n60 VSUBS 0.00946f
C245 B.n61 VSUBS 0.00946f
C246 B.n62 VSUBS 0.00946f
C247 B.n63 VSUBS 0.00946f
C248 B.n64 VSUBS 0.00946f
C249 B.n65 VSUBS 0.00946f
C250 B.n66 VSUBS 0.00946f
C251 B.n67 VSUBS 0.00946f
C252 B.n68 VSUBS 0.00946f
C253 B.n69 VSUBS 0.00946f
C254 B.n70 VSUBS 0.022009f
C255 B.n71 VSUBS 0.00946f
C256 B.n72 VSUBS 0.00946f
C257 B.n73 VSUBS 0.00946f
C258 B.n74 VSUBS 0.00946f
C259 B.n75 VSUBS 0.00946f
C260 B.n76 VSUBS 0.00946f
C261 B.n77 VSUBS 0.00946f
C262 B.n78 VSUBS 0.00946f
C263 B.n79 VSUBS 0.00946f
C264 B.n80 VSUBS 0.00946f
C265 B.n81 VSUBS 0.00946f
C266 B.n82 VSUBS 0.00946f
C267 B.n83 VSUBS 0.00946f
C268 B.n84 VSUBS 0.00946f
C269 B.n85 VSUBS 0.00946f
C270 B.n86 VSUBS 0.00946f
C271 B.n87 VSUBS 0.00946f
C272 B.n88 VSUBS 0.00946f
C273 B.n89 VSUBS 0.00946f
C274 B.n90 VSUBS 0.00946f
C275 B.n91 VSUBS 0.00946f
C276 B.n92 VSUBS 0.00946f
C277 B.n93 VSUBS 0.00946f
C278 B.n94 VSUBS 0.00946f
C279 B.n95 VSUBS 0.00946f
C280 B.n96 VSUBS 0.00946f
C281 B.n97 VSUBS 0.00946f
C282 B.n98 VSUBS 0.00946f
C283 B.n99 VSUBS 0.00946f
C284 B.n100 VSUBS 0.00946f
C285 B.n101 VSUBS 0.00946f
C286 B.n102 VSUBS 0.00946f
C287 B.n103 VSUBS 0.00946f
C288 B.n104 VSUBS 0.00946f
C289 B.n105 VSUBS 0.00946f
C290 B.n106 VSUBS 0.00946f
C291 B.n107 VSUBS 0.00946f
C292 B.n108 VSUBS 0.00946f
C293 B.n109 VSUBS 0.00946f
C294 B.n110 VSUBS 0.00946f
C295 B.n111 VSUBS 0.00946f
C296 B.n112 VSUBS 0.00946f
C297 B.n113 VSUBS 0.00946f
C298 B.n114 VSUBS 0.00946f
C299 B.n115 VSUBS 0.00946f
C300 B.n116 VSUBS 0.00946f
C301 B.n117 VSUBS 0.00946f
C302 B.n118 VSUBS 0.00946f
C303 B.n119 VSUBS 0.00946f
C304 B.n120 VSUBS 0.00946f
C305 B.n121 VSUBS 0.022785f
C306 B.n122 VSUBS 0.00946f
C307 B.n123 VSUBS 0.00946f
C308 B.n124 VSUBS 0.00946f
C309 B.n125 VSUBS 0.00946f
C310 B.n126 VSUBS 0.00946f
C311 B.n127 VSUBS 0.00946f
C312 B.n128 VSUBS 0.00946f
C313 B.n129 VSUBS 0.00946f
C314 B.n130 VSUBS 0.00946f
C315 B.n131 VSUBS 0.00946f
C316 B.n132 VSUBS 0.00946f
C317 B.n133 VSUBS 0.00946f
C318 B.n134 VSUBS 0.00946f
C319 B.n135 VSUBS 0.00946f
C320 B.n136 VSUBS 0.00946f
C321 B.n137 VSUBS 0.00946f
C322 B.t11 VSUBS 0.208004f
C323 B.t10 VSUBS 0.256852f
C324 B.t9 VSUBS 1.93559f
C325 B.n138 VSUBS 0.416322f
C326 B.n139 VSUBS 0.291769f
C327 B.n140 VSUBS 0.021917f
C328 B.n141 VSUBS 0.00946f
C329 B.n142 VSUBS 0.00946f
C330 B.n143 VSUBS 0.00946f
C331 B.n144 VSUBS 0.00946f
C332 B.n145 VSUBS 0.00946f
C333 B.t5 VSUBS 0.208001f
C334 B.t4 VSUBS 0.256849f
C335 B.t3 VSUBS 1.93559f
C336 B.n146 VSUBS 0.416325f
C337 B.n147 VSUBS 0.291773f
C338 B.n148 VSUBS 0.00946f
C339 B.n149 VSUBS 0.00946f
C340 B.n150 VSUBS 0.00946f
C341 B.n151 VSUBS 0.00946f
C342 B.n152 VSUBS 0.00946f
C343 B.n153 VSUBS 0.00946f
C344 B.n154 VSUBS 0.00946f
C345 B.n155 VSUBS 0.00946f
C346 B.n156 VSUBS 0.00946f
C347 B.n157 VSUBS 0.00946f
C348 B.n158 VSUBS 0.00946f
C349 B.n159 VSUBS 0.00946f
C350 B.n160 VSUBS 0.00946f
C351 B.n161 VSUBS 0.00946f
C352 B.n162 VSUBS 0.00946f
C353 B.n163 VSUBS 0.00946f
C354 B.n164 VSUBS 0.022009f
C355 B.n165 VSUBS 0.00946f
C356 B.n166 VSUBS 0.00946f
C357 B.n167 VSUBS 0.00946f
C358 B.n168 VSUBS 0.00946f
C359 B.n169 VSUBS 0.00946f
C360 B.n170 VSUBS 0.00946f
C361 B.n171 VSUBS 0.00946f
C362 B.n172 VSUBS 0.00946f
C363 B.n173 VSUBS 0.00946f
C364 B.n174 VSUBS 0.00946f
C365 B.n175 VSUBS 0.00946f
C366 B.n176 VSUBS 0.00946f
C367 B.n177 VSUBS 0.00946f
C368 B.n178 VSUBS 0.00946f
C369 B.n179 VSUBS 0.00946f
C370 B.n180 VSUBS 0.00946f
C371 B.n181 VSUBS 0.00946f
C372 B.n182 VSUBS 0.00946f
C373 B.n183 VSUBS 0.00946f
C374 B.n184 VSUBS 0.00946f
C375 B.n185 VSUBS 0.00946f
C376 B.n186 VSUBS 0.00946f
C377 B.n187 VSUBS 0.00946f
C378 B.n188 VSUBS 0.00946f
C379 B.n189 VSUBS 0.00946f
C380 B.n190 VSUBS 0.00946f
C381 B.n191 VSUBS 0.00946f
C382 B.n192 VSUBS 0.00946f
C383 B.n193 VSUBS 0.00946f
C384 B.n194 VSUBS 0.00946f
C385 B.n195 VSUBS 0.00946f
C386 B.n196 VSUBS 0.00946f
C387 B.n197 VSUBS 0.00946f
C388 B.n198 VSUBS 0.00946f
C389 B.n199 VSUBS 0.00946f
C390 B.n200 VSUBS 0.00946f
C391 B.n201 VSUBS 0.00946f
C392 B.n202 VSUBS 0.00946f
C393 B.n203 VSUBS 0.00946f
C394 B.n204 VSUBS 0.00946f
C395 B.n205 VSUBS 0.00946f
C396 B.n206 VSUBS 0.00946f
C397 B.n207 VSUBS 0.00946f
C398 B.n208 VSUBS 0.00946f
C399 B.n209 VSUBS 0.00946f
C400 B.n210 VSUBS 0.00946f
C401 B.n211 VSUBS 0.00946f
C402 B.n212 VSUBS 0.00946f
C403 B.n213 VSUBS 0.00946f
C404 B.n214 VSUBS 0.00946f
C405 B.n215 VSUBS 0.00946f
C406 B.n216 VSUBS 0.00946f
C407 B.n217 VSUBS 0.00946f
C408 B.n218 VSUBS 0.00946f
C409 B.n219 VSUBS 0.00946f
C410 B.n220 VSUBS 0.00946f
C411 B.n221 VSUBS 0.00946f
C412 B.n222 VSUBS 0.00946f
C413 B.n223 VSUBS 0.00946f
C414 B.n224 VSUBS 0.00946f
C415 B.n225 VSUBS 0.00946f
C416 B.n226 VSUBS 0.00946f
C417 B.n227 VSUBS 0.00946f
C418 B.n228 VSUBS 0.00946f
C419 B.n229 VSUBS 0.00946f
C420 B.n230 VSUBS 0.00946f
C421 B.n231 VSUBS 0.00946f
C422 B.n232 VSUBS 0.00946f
C423 B.n233 VSUBS 0.00946f
C424 B.n234 VSUBS 0.00946f
C425 B.n235 VSUBS 0.00946f
C426 B.n236 VSUBS 0.00946f
C427 B.n237 VSUBS 0.00946f
C428 B.n238 VSUBS 0.00946f
C429 B.n239 VSUBS 0.00946f
C430 B.n240 VSUBS 0.00946f
C431 B.n241 VSUBS 0.00946f
C432 B.n242 VSUBS 0.00946f
C433 B.n243 VSUBS 0.00946f
C434 B.n244 VSUBS 0.00946f
C435 B.n245 VSUBS 0.00946f
C436 B.n246 VSUBS 0.00946f
C437 B.n247 VSUBS 0.00946f
C438 B.n248 VSUBS 0.00946f
C439 B.n249 VSUBS 0.00946f
C440 B.n250 VSUBS 0.00946f
C441 B.n251 VSUBS 0.00946f
C442 B.n252 VSUBS 0.00946f
C443 B.n253 VSUBS 0.00946f
C444 B.n254 VSUBS 0.00946f
C445 B.n255 VSUBS 0.00946f
C446 B.n256 VSUBS 0.00946f
C447 B.n257 VSUBS 0.00946f
C448 B.n258 VSUBS 0.00946f
C449 B.n259 VSUBS 0.00946f
C450 B.n260 VSUBS 0.00946f
C451 B.n261 VSUBS 0.022009f
C452 B.n262 VSUBS 0.022785f
C453 B.n263 VSUBS 0.022785f
C454 B.n264 VSUBS 0.00946f
C455 B.n265 VSUBS 0.00946f
C456 B.n266 VSUBS 0.00946f
C457 B.n267 VSUBS 0.00946f
C458 B.n268 VSUBS 0.00946f
C459 B.n269 VSUBS 0.00946f
C460 B.n270 VSUBS 0.00946f
C461 B.n271 VSUBS 0.00946f
C462 B.n272 VSUBS 0.00946f
C463 B.n273 VSUBS 0.00946f
C464 B.n274 VSUBS 0.00946f
C465 B.n275 VSUBS 0.00946f
C466 B.n276 VSUBS 0.00946f
C467 B.n277 VSUBS 0.00946f
C468 B.n278 VSUBS 0.00946f
C469 B.n279 VSUBS 0.00946f
C470 B.n280 VSUBS 0.00946f
C471 B.n281 VSUBS 0.00946f
C472 B.n282 VSUBS 0.00946f
C473 B.n283 VSUBS 0.00946f
C474 B.n284 VSUBS 0.00946f
C475 B.n285 VSUBS 0.00946f
C476 B.n286 VSUBS 0.00946f
C477 B.n287 VSUBS 0.00946f
C478 B.n288 VSUBS 0.00946f
C479 B.n289 VSUBS 0.00946f
C480 B.n290 VSUBS 0.00946f
C481 B.n291 VSUBS 0.00946f
C482 B.n292 VSUBS 0.00946f
C483 B.n293 VSUBS 0.00946f
C484 B.n294 VSUBS 0.00946f
C485 B.n295 VSUBS 0.00946f
C486 B.n296 VSUBS 0.00946f
C487 B.n297 VSUBS 0.00946f
C488 B.n298 VSUBS 0.00946f
C489 B.n299 VSUBS 0.00946f
C490 B.n300 VSUBS 0.00946f
C491 B.n301 VSUBS 0.00946f
C492 B.n302 VSUBS 0.00946f
C493 B.n303 VSUBS 0.00946f
C494 B.n304 VSUBS 0.00946f
C495 B.n305 VSUBS 0.00946f
C496 B.n306 VSUBS 0.00946f
C497 B.n307 VSUBS 0.00946f
C498 B.n308 VSUBS 0.00946f
C499 B.n309 VSUBS 0.00946f
C500 B.n310 VSUBS 0.00946f
C501 B.n311 VSUBS 0.00946f
C502 B.n312 VSUBS 0.006538f
C503 B.n313 VSUBS 0.021917f
C504 B.n314 VSUBS 0.007651f
C505 B.n315 VSUBS 0.00946f
C506 B.n316 VSUBS 0.00946f
C507 B.n317 VSUBS 0.00946f
C508 B.n318 VSUBS 0.00946f
C509 B.n319 VSUBS 0.00946f
C510 B.n320 VSUBS 0.00946f
C511 B.n321 VSUBS 0.00946f
C512 B.n322 VSUBS 0.00946f
C513 B.n323 VSUBS 0.00946f
C514 B.n324 VSUBS 0.00946f
C515 B.n325 VSUBS 0.00946f
C516 B.n326 VSUBS 0.007651f
C517 B.n327 VSUBS 0.00946f
C518 B.n328 VSUBS 0.00946f
C519 B.n329 VSUBS 0.006538f
C520 B.n330 VSUBS 0.00946f
C521 B.n331 VSUBS 0.00946f
C522 B.n332 VSUBS 0.00946f
C523 B.n333 VSUBS 0.00946f
C524 B.n334 VSUBS 0.00946f
C525 B.n335 VSUBS 0.00946f
C526 B.n336 VSUBS 0.00946f
C527 B.n337 VSUBS 0.00946f
C528 B.n338 VSUBS 0.00946f
C529 B.n339 VSUBS 0.00946f
C530 B.n340 VSUBS 0.00946f
C531 B.n341 VSUBS 0.00946f
C532 B.n342 VSUBS 0.00946f
C533 B.n343 VSUBS 0.00946f
C534 B.n344 VSUBS 0.00946f
C535 B.n345 VSUBS 0.00946f
C536 B.n346 VSUBS 0.00946f
C537 B.n347 VSUBS 0.00946f
C538 B.n348 VSUBS 0.00946f
C539 B.n349 VSUBS 0.00946f
C540 B.n350 VSUBS 0.00946f
C541 B.n351 VSUBS 0.00946f
C542 B.n352 VSUBS 0.00946f
C543 B.n353 VSUBS 0.00946f
C544 B.n354 VSUBS 0.00946f
C545 B.n355 VSUBS 0.00946f
C546 B.n356 VSUBS 0.00946f
C547 B.n357 VSUBS 0.00946f
C548 B.n358 VSUBS 0.00946f
C549 B.n359 VSUBS 0.00946f
C550 B.n360 VSUBS 0.00946f
C551 B.n361 VSUBS 0.00946f
C552 B.n362 VSUBS 0.00946f
C553 B.n363 VSUBS 0.00946f
C554 B.n364 VSUBS 0.00946f
C555 B.n365 VSUBS 0.00946f
C556 B.n366 VSUBS 0.00946f
C557 B.n367 VSUBS 0.00946f
C558 B.n368 VSUBS 0.00946f
C559 B.n369 VSUBS 0.00946f
C560 B.n370 VSUBS 0.00946f
C561 B.n371 VSUBS 0.00946f
C562 B.n372 VSUBS 0.00946f
C563 B.n373 VSUBS 0.00946f
C564 B.n374 VSUBS 0.00946f
C565 B.n375 VSUBS 0.00946f
C566 B.n376 VSUBS 0.00946f
C567 B.n377 VSUBS 0.00946f
C568 B.n378 VSUBS 0.021688f
C569 B.n379 VSUBS 0.023107f
C570 B.n380 VSUBS 0.022009f
C571 B.n381 VSUBS 0.00946f
C572 B.n382 VSUBS 0.00946f
C573 B.n383 VSUBS 0.00946f
C574 B.n384 VSUBS 0.00946f
C575 B.n385 VSUBS 0.00946f
C576 B.n386 VSUBS 0.00946f
C577 B.n387 VSUBS 0.00946f
C578 B.n388 VSUBS 0.00946f
C579 B.n389 VSUBS 0.00946f
C580 B.n390 VSUBS 0.00946f
C581 B.n391 VSUBS 0.00946f
C582 B.n392 VSUBS 0.00946f
C583 B.n393 VSUBS 0.00946f
C584 B.n394 VSUBS 0.00946f
C585 B.n395 VSUBS 0.00946f
C586 B.n396 VSUBS 0.00946f
C587 B.n397 VSUBS 0.00946f
C588 B.n398 VSUBS 0.00946f
C589 B.n399 VSUBS 0.00946f
C590 B.n400 VSUBS 0.00946f
C591 B.n401 VSUBS 0.00946f
C592 B.n402 VSUBS 0.00946f
C593 B.n403 VSUBS 0.00946f
C594 B.n404 VSUBS 0.00946f
C595 B.n405 VSUBS 0.00946f
C596 B.n406 VSUBS 0.00946f
C597 B.n407 VSUBS 0.00946f
C598 B.n408 VSUBS 0.00946f
C599 B.n409 VSUBS 0.00946f
C600 B.n410 VSUBS 0.00946f
C601 B.n411 VSUBS 0.00946f
C602 B.n412 VSUBS 0.00946f
C603 B.n413 VSUBS 0.00946f
C604 B.n414 VSUBS 0.00946f
C605 B.n415 VSUBS 0.00946f
C606 B.n416 VSUBS 0.00946f
C607 B.n417 VSUBS 0.00946f
C608 B.n418 VSUBS 0.00946f
C609 B.n419 VSUBS 0.00946f
C610 B.n420 VSUBS 0.00946f
C611 B.n421 VSUBS 0.00946f
C612 B.n422 VSUBS 0.00946f
C613 B.n423 VSUBS 0.00946f
C614 B.n424 VSUBS 0.00946f
C615 B.n425 VSUBS 0.00946f
C616 B.n426 VSUBS 0.00946f
C617 B.n427 VSUBS 0.00946f
C618 B.n428 VSUBS 0.00946f
C619 B.n429 VSUBS 0.00946f
C620 B.n430 VSUBS 0.00946f
C621 B.n431 VSUBS 0.00946f
C622 B.n432 VSUBS 0.00946f
C623 B.n433 VSUBS 0.00946f
C624 B.n434 VSUBS 0.00946f
C625 B.n435 VSUBS 0.00946f
C626 B.n436 VSUBS 0.00946f
C627 B.n437 VSUBS 0.00946f
C628 B.n438 VSUBS 0.00946f
C629 B.n439 VSUBS 0.00946f
C630 B.n440 VSUBS 0.00946f
C631 B.n441 VSUBS 0.00946f
C632 B.n442 VSUBS 0.00946f
C633 B.n443 VSUBS 0.00946f
C634 B.n444 VSUBS 0.00946f
C635 B.n445 VSUBS 0.00946f
C636 B.n446 VSUBS 0.00946f
C637 B.n447 VSUBS 0.00946f
C638 B.n448 VSUBS 0.00946f
C639 B.n449 VSUBS 0.00946f
C640 B.n450 VSUBS 0.00946f
C641 B.n451 VSUBS 0.00946f
C642 B.n452 VSUBS 0.00946f
C643 B.n453 VSUBS 0.00946f
C644 B.n454 VSUBS 0.00946f
C645 B.n455 VSUBS 0.00946f
C646 B.n456 VSUBS 0.00946f
C647 B.n457 VSUBS 0.00946f
C648 B.n458 VSUBS 0.00946f
C649 B.n459 VSUBS 0.00946f
C650 B.n460 VSUBS 0.00946f
C651 B.n461 VSUBS 0.00946f
C652 B.n462 VSUBS 0.00946f
C653 B.n463 VSUBS 0.00946f
C654 B.n464 VSUBS 0.00946f
C655 B.n465 VSUBS 0.00946f
C656 B.n466 VSUBS 0.00946f
C657 B.n467 VSUBS 0.00946f
C658 B.n468 VSUBS 0.00946f
C659 B.n469 VSUBS 0.00946f
C660 B.n470 VSUBS 0.00946f
C661 B.n471 VSUBS 0.00946f
C662 B.n472 VSUBS 0.00946f
C663 B.n473 VSUBS 0.00946f
C664 B.n474 VSUBS 0.00946f
C665 B.n475 VSUBS 0.00946f
C666 B.n476 VSUBS 0.00946f
C667 B.n477 VSUBS 0.00946f
C668 B.n478 VSUBS 0.00946f
C669 B.n479 VSUBS 0.00946f
C670 B.n480 VSUBS 0.00946f
C671 B.n481 VSUBS 0.00946f
C672 B.n482 VSUBS 0.00946f
C673 B.n483 VSUBS 0.00946f
C674 B.n484 VSUBS 0.00946f
C675 B.n485 VSUBS 0.00946f
C676 B.n486 VSUBS 0.00946f
C677 B.n487 VSUBS 0.00946f
C678 B.n488 VSUBS 0.00946f
C679 B.n489 VSUBS 0.00946f
C680 B.n490 VSUBS 0.00946f
C681 B.n491 VSUBS 0.00946f
C682 B.n492 VSUBS 0.00946f
C683 B.n493 VSUBS 0.00946f
C684 B.n494 VSUBS 0.00946f
C685 B.n495 VSUBS 0.00946f
C686 B.n496 VSUBS 0.00946f
C687 B.n497 VSUBS 0.00946f
C688 B.n498 VSUBS 0.00946f
C689 B.n499 VSUBS 0.00946f
C690 B.n500 VSUBS 0.00946f
C691 B.n501 VSUBS 0.00946f
C692 B.n502 VSUBS 0.00946f
C693 B.n503 VSUBS 0.00946f
C694 B.n504 VSUBS 0.00946f
C695 B.n505 VSUBS 0.00946f
C696 B.n506 VSUBS 0.00946f
C697 B.n507 VSUBS 0.00946f
C698 B.n508 VSUBS 0.00946f
C699 B.n509 VSUBS 0.00946f
C700 B.n510 VSUBS 0.00946f
C701 B.n511 VSUBS 0.00946f
C702 B.n512 VSUBS 0.00946f
C703 B.n513 VSUBS 0.00946f
C704 B.n514 VSUBS 0.00946f
C705 B.n515 VSUBS 0.00946f
C706 B.n516 VSUBS 0.00946f
C707 B.n517 VSUBS 0.00946f
C708 B.n518 VSUBS 0.00946f
C709 B.n519 VSUBS 0.00946f
C710 B.n520 VSUBS 0.00946f
C711 B.n521 VSUBS 0.00946f
C712 B.n522 VSUBS 0.00946f
C713 B.n523 VSUBS 0.00946f
C714 B.n524 VSUBS 0.00946f
C715 B.n525 VSUBS 0.00946f
C716 B.n526 VSUBS 0.00946f
C717 B.n527 VSUBS 0.00946f
C718 B.n528 VSUBS 0.00946f
C719 B.n529 VSUBS 0.00946f
C720 B.n530 VSUBS 0.00946f
C721 B.n531 VSUBS 0.022009f
C722 B.n532 VSUBS 0.022785f
C723 B.n533 VSUBS 0.022785f
C724 B.n534 VSUBS 0.00946f
C725 B.n535 VSUBS 0.00946f
C726 B.n536 VSUBS 0.00946f
C727 B.n537 VSUBS 0.00946f
C728 B.n538 VSUBS 0.00946f
C729 B.n539 VSUBS 0.00946f
C730 B.n540 VSUBS 0.00946f
C731 B.n541 VSUBS 0.00946f
C732 B.n542 VSUBS 0.00946f
C733 B.n543 VSUBS 0.00946f
C734 B.n544 VSUBS 0.00946f
C735 B.n545 VSUBS 0.00946f
C736 B.n546 VSUBS 0.00946f
C737 B.n547 VSUBS 0.00946f
C738 B.n548 VSUBS 0.00946f
C739 B.n549 VSUBS 0.00946f
C740 B.n550 VSUBS 0.00946f
C741 B.n551 VSUBS 0.00946f
C742 B.n552 VSUBS 0.00946f
C743 B.n553 VSUBS 0.00946f
C744 B.n554 VSUBS 0.00946f
C745 B.n555 VSUBS 0.00946f
C746 B.n556 VSUBS 0.00946f
C747 B.n557 VSUBS 0.00946f
C748 B.n558 VSUBS 0.00946f
C749 B.n559 VSUBS 0.00946f
C750 B.n560 VSUBS 0.00946f
C751 B.n561 VSUBS 0.00946f
C752 B.n562 VSUBS 0.00946f
C753 B.n563 VSUBS 0.00946f
C754 B.n564 VSUBS 0.00946f
C755 B.n565 VSUBS 0.00946f
C756 B.n566 VSUBS 0.00946f
C757 B.n567 VSUBS 0.00946f
C758 B.n568 VSUBS 0.00946f
C759 B.n569 VSUBS 0.00946f
C760 B.n570 VSUBS 0.00946f
C761 B.n571 VSUBS 0.00946f
C762 B.n572 VSUBS 0.00946f
C763 B.n573 VSUBS 0.00946f
C764 B.n574 VSUBS 0.00946f
C765 B.n575 VSUBS 0.00946f
C766 B.n576 VSUBS 0.00946f
C767 B.n577 VSUBS 0.00946f
C768 B.n578 VSUBS 0.00946f
C769 B.n579 VSUBS 0.00946f
C770 B.n580 VSUBS 0.00946f
C771 B.n581 VSUBS 0.00946f
C772 B.n582 VSUBS 0.006538f
C773 B.n583 VSUBS 0.021917f
C774 B.n584 VSUBS 0.007651f
C775 B.n585 VSUBS 0.00946f
C776 B.n586 VSUBS 0.00946f
C777 B.n587 VSUBS 0.00946f
C778 B.n588 VSUBS 0.00946f
C779 B.n589 VSUBS 0.00946f
C780 B.n590 VSUBS 0.00946f
C781 B.n591 VSUBS 0.00946f
C782 B.n592 VSUBS 0.00946f
C783 B.n593 VSUBS 0.00946f
C784 B.n594 VSUBS 0.00946f
C785 B.n595 VSUBS 0.00946f
C786 B.n596 VSUBS 0.007651f
C787 B.n597 VSUBS 0.00946f
C788 B.n598 VSUBS 0.00946f
C789 B.n599 VSUBS 0.006538f
C790 B.n600 VSUBS 0.00946f
C791 B.n601 VSUBS 0.00946f
C792 B.n602 VSUBS 0.00946f
C793 B.n603 VSUBS 0.00946f
C794 B.n604 VSUBS 0.00946f
C795 B.n605 VSUBS 0.00946f
C796 B.n606 VSUBS 0.00946f
C797 B.n607 VSUBS 0.00946f
C798 B.n608 VSUBS 0.00946f
C799 B.n609 VSUBS 0.00946f
C800 B.n610 VSUBS 0.00946f
C801 B.n611 VSUBS 0.00946f
C802 B.n612 VSUBS 0.00946f
C803 B.n613 VSUBS 0.00946f
C804 B.n614 VSUBS 0.00946f
C805 B.n615 VSUBS 0.00946f
C806 B.n616 VSUBS 0.00946f
C807 B.n617 VSUBS 0.00946f
C808 B.n618 VSUBS 0.00946f
C809 B.n619 VSUBS 0.00946f
C810 B.n620 VSUBS 0.00946f
C811 B.n621 VSUBS 0.00946f
C812 B.n622 VSUBS 0.00946f
C813 B.n623 VSUBS 0.00946f
C814 B.n624 VSUBS 0.00946f
C815 B.n625 VSUBS 0.00946f
C816 B.n626 VSUBS 0.00946f
C817 B.n627 VSUBS 0.00946f
C818 B.n628 VSUBS 0.00946f
C819 B.n629 VSUBS 0.00946f
C820 B.n630 VSUBS 0.00946f
C821 B.n631 VSUBS 0.00946f
C822 B.n632 VSUBS 0.00946f
C823 B.n633 VSUBS 0.00946f
C824 B.n634 VSUBS 0.00946f
C825 B.n635 VSUBS 0.00946f
C826 B.n636 VSUBS 0.00946f
C827 B.n637 VSUBS 0.00946f
C828 B.n638 VSUBS 0.00946f
C829 B.n639 VSUBS 0.00946f
C830 B.n640 VSUBS 0.00946f
C831 B.n641 VSUBS 0.00946f
C832 B.n642 VSUBS 0.00946f
C833 B.n643 VSUBS 0.00946f
C834 B.n644 VSUBS 0.00946f
C835 B.n645 VSUBS 0.00946f
C836 B.n646 VSUBS 0.00946f
C837 B.n647 VSUBS 0.00946f
C838 B.n648 VSUBS 0.022785f
C839 B.n649 VSUBS 0.022009f
C840 B.n650 VSUBS 0.022009f
C841 B.n651 VSUBS 0.00946f
C842 B.n652 VSUBS 0.00946f
C843 B.n653 VSUBS 0.00946f
C844 B.n654 VSUBS 0.00946f
C845 B.n655 VSUBS 0.00946f
C846 B.n656 VSUBS 0.00946f
C847 B.n657 VSUBS 0.00946f
C848 B.n658 VSUBS 0.00946f
C849 B.n659 VSUBS 0.00946f
C850 B.n660 VSUBS 0.00946f
C851 B.n661 VSUBS 0.00946f
C852 B.n662 VSUBS 0.00946f
C853 B.n663 VSUBS 0.00946f
C854 B.n664 VSUBS 0.00946f
C855 B.n665 VSUBS 0.00946f
C856 B.n666 VSUBS 0.00946f
C857 B.n667 VSUBS 0.00946f
C858 B.n668 VSUBS 0.00946f
C859 B.n669 VSUBS 0.00946f
C860 B.n670 VSUBS 0.00946f
C861 B.n671 VSUBS 0.00946f
C862 B.n672 VSUBS 0.00946f
C863 B.n673 VSUBS 0.00946f
C864 B.n674 VSUBS 0.00946f
C865 B.n675 VSUBS 0.00946f
C866 B.n676 VSUBS 0.00946f
C867 B.n677 VSUBS 0.00946f
C868 B.n678 VSUBS 0.00946f
C869 B.n679 VSUBS 0.00946f
C870 B.n680 VSUBS 0.00946f
C871 B.n681 VSUBS 0.00946f
C872 B.n682 VSUBS 0.00946f
C873 B.n683 VSUBS 0.00946f
C874 B.n684 VSUBS 0.00946f
C875 B.n685 VSUBS 0.00946f
C876 B.n686 VSUBS 0.00946f
C877 B.n687 VSUBS 0.00946f
C878 B.n688 VSUBS 0.00946f
C879 B.n689 VSUBS 0.00946f
C880 B.n690 VSUBS 0.00946f
C881 B.n691 VSUBS 0.00946f
C882 B.n692 VSUBS 0.00946f
C883 B.n693 VSUBS 0.00946f
C884 B.n694 VSUBS 0.00946f
C885 B.n695 VSUBS 0.00946f
C886 B.n696 VSUBS 0.00946f
C887 B.n697 VSUBS 0.00946f
C888 B.n698 VSUBS 0.00946f
C889 B.n699 VSUBS 0.00946f
C890 B.n700 VSUBS 0.00946f
C891 B.n701 VSUBS 0.00946f
C892 B.n702 VSUBS 0.00946f
C893 B.n703 VSUBS 0.00946f
C894 B.n704 VSUBS 0.00946f
C895 B.n705 VSUBS 0.00946f
C896 B.n706 VSUBS 0.00946f
C897 B.n707 VSUBS 0.00946f
C898 B.n708 VSUBS 0.00946f
C899 B.n709 VSUBS 0.00946f
C900 B.n710 VSUBS 0.00946f
C901 B.n711 VSUBS 0.00946f
C902 B.n712 VSUBS 0.00946f
C903 B.n713 VSUBS 0.00946f
C904 B.n714 VSUBS 0.00946f
C905 B.n715 VSUBS 0.00946f
C906 B.n716 VSUBS 0.00946f
C907 B.n717 VSUBS 0.00946f
C908 B.n718 VSUBS 0.00946f
C909 B.n719 VSUBS 0.00946f
C910 B.n720 VSUBS 0.00946f
C911 B.n721 VSUBS 0.00946f
C912 B.n722 VSUBS 0.00946f
C913 B.n723 VSUBS 0.012344f
C914 B.n724 VSUBS 0.01315f
C915 B.n725 VSUBS 0.02615f
C916 VTAIL.t11 VSUBS 0.228954f
C917 VTAIL.t10 VSUBS 0.228954f
C918 VTAIL.n0 VSUBS 1.57278f
C919 VTAIL.n1 VSUBS 0.92761f
C920 VTAIL.n2 VSUBS 0.033262f
C921 VTAIL.n3 VSUBS 0.030987f
C922 VTAIL.n4 VSUBS 0.016651f
C923 VTAIL.n5 VSUBS 0.039357f
C924 VTAIL.n6 VSUBS 0.017141f
C925 VTAIL.n7 VSUBS 0.030987f
C926 VTAIL.n8 VSUBS 0.017631f
C927 VTAIL.n9 VSUBS 0.039357f
C928 VTAIL.n10 VSUBS 0.017631f
C929 VTAIL.n11 VSUBS 0.030987f
C930 VTAIL.n12 VSUBS 0.016651f
C931 VTAIL.n13 VSUBS 0.039357f
C932 VTAIL.n14 VSUBS 0.017631f
C933 VTAIL.n15 VSUBS 1.16261f
C934 VTAIL.n16 VSUBS 0.016651f
C935 VTAIL.t7 VSUBS 0.084583f
C936 VTAIL.n17 VSUBS 0.206955f
C937 VTAIL.n18 VSUBS 0.029607f
C938 VTAIL.n19 VSUBS 0.029518f
C939 VTAIL.n20 VSUBS 0.039357f
C940 VTAIL.n21 VSUBS 0.017631f
C941 VTAIL.n22 VSUBS 0.016651f
C942 VTAIL.n23 VSUBS 0.030987f
C943 VTAIL.n24 VSUBS 0.030987f
C944 VTAIL.n25 VSUBS 0.016651f
C945 VTAIL.n26 VSUBS 0.017631f
C946 VTAIL.n27 VSUBS 0.039357f
C947 VTAIL.n28 VSUBS 0.039357f
C948 VTAIL.n29 VSUBS 0.017631f
C949 VTAIL.n30 VSUBS 0.016651f
C950 VTAIL.n31 VSUBS 0.030987f
C951 VTAIL.n32 VSUBS 0.030987f
C952 VTAIL.n33 VSUBS 0.016651f
C953 VTAIL.n34 VSUBS 0.016651f
C954 VTAIL.n35 VSUBS 0.017631f
C955 VTAIL.n36 VSUBS 0.039357f
C956 VTAIL.n37 VSUBS 0.039357f
C957 VTAIL.n38 VSUBS 0.039357f
C958 VTAIL.n39 VSUBS 0.017141f
C959 VTAIL.n40 VSUBS 0.016651f
C960 VTAIL.n41 VSUBS 0.030987f
C961 VTAIL.n42 VSUBS 0.030987f
C962 VTAIL.n43 VSUBS 0.016651f
C963 VTAIL.n44 VSUBS 0.017631f
C964 VTAIL.n45 VSUBS 0.039357f
C965 VTAIL.n46 VSUBS 0.092602f
C966 VTAIL.n47 VSUBS 0.017631f
C967 VTAIL.n48 VSUBS 0.016651f
C968 VTAIL.n49 VSUBS 0.076282f
C969 VTAIL.n50 VSUBS 0.046589f
C970 VTAIL.n51 VSUBS 0.540818f
C971 VTAIL.t4 VSUBS 0.228954f
C972 VTAIL.t8 VSUBS 0.228954f
C973 VTAIL.n52 VSUBS 1.57278f
C974 VTAIL.n53 VSUBS 2.79784f
C975 VTAIL.t2 VSUBS 0.228954f
C976 VTAIL.t9 VSUBS 0.228954f
C977 VTAIL.n54 VSUBS 1.57279f
C978 VTAIL.n55 VSUBS 2.79783f
C979 VTAIL.n56 VSUBS 0.033262f
C980 VTAIL.n57 VSUBS 0.030987f
C981 VTAIL.n58 VSUBS 0.016651f
C982 VTAIL.n59 VSUBS 0.039357f
C983 VTAIL.n60 VSUBS 0.017141f
C984 VTAIL.n61 VSUBS 0.030987f
C985 VTAIL.n62 VSUBS 0.017141f
C986 VTAIL.n63 VSUBS 0.016651f
C987 VTAIL.n64 VSUBS 0.039357f
C988 VTAIL.n65 VSUBS 0.039357f
C989 VTAIL.n66 VSUBS 0.017631f
C990 VTAIL.n67 VSUBS 0.030987f
C991 VTAIL.n68 VSUBS 0.016651f
C992 VTAIL.n69 VSUBS 0.039357f
C993 VTAIL.n70 VSUBS 0.017631f
C994 VTAIL.n71 VSUBS 1.16261f
C995 VTAIL.n72 VSUBS 0.016651f
C996 VTAIL.t0 VSUBS 0.084583f
C997 VTAIL.n73 VSUBS 0.206955f
C998 VTAIL.n74 VSUBS 0.029607f
C999 VTAIL.n75 VSUBS 0.029518f
C1000 VTAIL.n76 VSUBS 0.039357f
C1001 VTAIL.n77 VSUBS 0.017631f
C1002 VTAIL.n78 VSUBS 0.016651f
C1003 VTAIL.n79 VSUBS 0.030987f
C1004 VTAIL.n80 VSUBS 0.030987f
C1005 VTAIL.n81 VSUBS 0.016651f
C1006 VTAIL.n82 VSUBS 0.017631f
C1007 VTAIL.n83 VSUBS 0.039357f
C1008 VTAIL.n84 VSUBS 0.039357f
C1009 VTAIL.n85 VSUBS 0.017631f
C1010 VTAIL.n86 VSUBS 0.016651f
C1011 VTAIL.n87 VSUBS 0.030987f
C1012 VTAIL.n88 VSUBS 0.030987f
C1013 VTAIL.n89 VSUBS 0.016651f
C1014 VTAIL.n90 VSUBS 0.017631f
C1015 VTAIL.n91 VSUBS 0.039357f
C1016 VTAIL.n92 VSUBS 0.039357f
C1017 VTAIL.n93 VSUBS 0.017631f
C1018 VTAIL.n94 VSUBS 0.016651f
C1019 VTAIL.n95 VSUBS 0.030987f
C1020 VTAIL.n96 VSUBS 0.030987f
C1021 VTAIL.n97 VSUBS 0.016651f
C1022 VTAIL.n98 VSUBS 0.017631f
C1023 VTAIL.n99 VSUBS 0.039357f
C1024 VTAIL.n100 VSUBS 0.092602f
C1025 VTAIL.n101 VSUBS 0.017631f
C1026 VTAIL.n102 VSUBS 0.016651f
C1027 VTAIL.n103 VSUBS 0.076282f
C1028 VTAIL.n104 VSUBS 0.046589f
C1029 VTAIL.n105 VSUBS 0.540818f
C1030 VTAIL.t3 VSUBS 0.228954f
C1031 VTAIL.t6 VSUBS 0.228954f
C1032 VTAIL.n106 VSUBS 1.57279f
C1033 VTAIL.n107 VSUBS 1.15419f
C1034 VTAIL.n108 VSUBS 0.033262f
C1035 VTAIL.n109 VSUBS 0.030987f
C1036 VTAIL.n110 VSUBS 0.016651f
C1037 VTAIL.n111 VSUBS 0.039357f
C1038 VTAIL.n112 VSUBS 0.017141f
C1039 VTAIL.n113 VSUBS 0.030987f
C1040 VTAIL.n114 VSUBS 0.017141f
C1041 VTAIL.n115 VSUBS 0.016651f
C1042 VTAIL.n116 VSUBS 0.039357f
C1043 VTAIL.n117 VSUBS 0.039357f
C1044 VTAIL.n118 VSUBS 0.017631f
C1045 VTAIL.n119 VSUBS 0.030987f
C1046 VTAIL.n120 VSUBS 0.016651f
C1047 VTAIL.n121 VSUBS 0.039357f
C1048 VTAIL.n122 VSUBS 0.017631f
C1049 VTAIL.n123 VSUBS 1.16261f
C1050 VTAIL.n124 VSUBS 0.016651f
C1051 VTAIL.t5 VSUBS 0.084583f
C1052 VTAIL.n125 VSUBS 0.206955f
C1053 VTAIL.n126 VSUBS 0.029607f
C1054 VTAIL.n127 VSUBS 0.029518f
C1055 VTAIL.n128 VSUBS 0.039357f
C1056 VTAIL.n129 VSUBS 0.017631f
C1057 VTAIL.n130 VSUBS 0.016651f
C1058 VTAIL.n131 VSUBS 0.030987f
C1059 VTAIL.n132 VSUBS 0.030987f
C1060 VTAIL.n133 VSUBS 0.016651f
C1061 VTAIL.n134 VSUBS 0.017631f
C1062 VTAIL.n135 VSUBS 0.039357f
C1063 VTAIL.n136 VSUBS 0.039357f
C1064 VTAIL.n137 VSUBS 0.017631f
C1065 VTAIL.n138 VSUBS 0.016651f
C1066 VTAIL.n139 VSUBS 0.030987f
C1067 VTAIL.n140 VSUBS 0.030987f
C1068 VTAIL.n141 VSUBS 0.016651f
C1069 VTAIL.n142 VSUBS 0.017631f
C1070 VTAIL.n143 VSUBS 0.039357f
C1071 VTAIL.n144 VSUBS 0.039357f
C1072 VTAIL.n145 VSUBS 0.017631f
C1073 VTAIL.n146 VSUBS 0.016651f
C1074 VTAIL.n147 VSUBS 0.030987f
C1075 VTAIL.n148 VSUBS 0.030987f
C1076 VTAIL.n149 VSUBS 0.016651f
C1077 VTAIL.n150 VSUBS 0.017631f
C1078 VTAIL.n151 VSUBS 0.039357f
C1079 VTAIL.n152 VSUBS 0.092602f
C1080 VTAIL.n153 VSUBS 0.017631f
C1081 VTAIL.n154 VSUBS 0.016651f
C1082 VTAIL.n155 VSUBS 0.076282f
C1083 VTAIL.n156 VSUBS 0.046589f
C1084 VTAIL.n157 VSUBS 1.87458f
C1085 VTAIL.n158 VSUBS 0.033262f
C1086 VTAIL.n159 VSUBS 0.030987f
C1087 VTAIL.n160 VSUBS 0.016651f
C1088 VTAIL.n161 VSUBS 0.039357f
C1089 VTAIL.n162 VSUBS 0.017141f
C1090 VTAIL.n163 VSUBS 0.030987f
C1091 VTAIL.n164 VSUBS 0.017631f
C1092 VTAIL.n165 VSUBS 0.039357f
C1093 VTAIL.n166 VSUBS 0.017631f
C1094 VTAIL.n167 VSUBS 0.030987f
C1095 VTAIL.n168 VSUBS 0.016651f
C1096 VTAIL.n169 VSUBS 0.039357f
C1097 VTAIL.n170 VSUBS 0.017631f
C1098 VTAIL.n171 VSUBS 1.16261f
C1099 VTAIL.n172 VSUBS 0.016651f
C1100 VTAIL.t1 VSUBS 0.084583f
C1101 VTAIL.n173 VSUBS 0.206955f
C1102 VTAIL.n174 VSUBS 0.029607f
C1103 VTAIL.n175 VSUBS 0.029518f
C1104 VTAIL.n176 VSUBS 0.039357f
C1105 VTAIL.n177 VSUBS 0.017631f
C1106 VTAIL.n178 VSUBS 0.016651f
C1107 VTAIL.n179 VSUBS 0.030987f
C1108 VTAIL.n180 VSUBS 0.030987f
C1109 VTAIL.n181 VSUBS 0.016651f
C1110 VTAIL.n182 VSUBS 0.017631f
C1111 VTAIL.n183 VSUBS 0.039357f
C1112 VTAIL.n184 VSUBS 0.039357f
C1113 VTAIL.n185 VSUBS 0.017631f
C1114 VTAIL.n186 VSUBS 0.016651f
C1115 VTAIL.n187 VSUBS 0.030987f
C1116 VTAIL.n188 VSUBS 0.030987f
C1117 VTAIL.n189 VSUBS 0.016651f
C1118 VTAIL.n190 VSUBS 0.016651f
C1119 VTAIL.n191 VSUBS 0.017631f
C1120 VTAIL.n192 VSUBS 0.039357f
C1121 VTAIL.n193 VSUBS 0.039357f
C1122 VTAIL.n194 VSUBS 0.039357f
C1123 VTAIL.n195 VSUBS 0.017141f
C1124 VTAIL.n196 VSUBS 0.016651f
C1125 VTAIL.n197 VSUBS 0.030987f
C1126 VTAIL.n198 VSUBS 0.030987f
C1127 VTAIL.n199 VSUBS 0.016651f
C1128 VTAIL.n200 VSUBS 0.017631f
C1129 VTAIL.n201 VSUBS 0.039357f
C1130 VTAIL.n202 VSUBS 0.092602f
C1131 VTAIL.n203 VSUBS 0.017631f
C1132 VTAIL.n204 VSUBS 0.016651f
C1133 VTAIL.n205 VSUBS 0.076282f
C1134 VTAIL.n206 VSUBS 0.046589f
C1135 VTAIL.n207 VSUBS 1.7913f
C1136 VDD1.n0 VSUBS 0.031434f
C1137 VDD1.n1 VSUBS 0.029284f
C1138 VDD1.n2 VSUBS 0.015736f
C1139 VDD1.n3 VSUBS 0.037194f
C1140 VDD1.n4 VSUBS 0.016199f
C1141 VDD1.n5 VSUBS 0.029284f
C1142 VDD1.n6 VSUBS 0.016199f
C1143 VDD1.n7 VSUBS 0.015736f
C1144 VDD1.n8 VSUBS 0.037194f
C1145 VDD1.n9 VSUBS 0.037194f
C1146 VDD1.n10 VSUBS 0.016662f
C1147 VDD1.n11 VSUBS 0.029284f
C1148 VDD1.n12 VSUBS 0.015736f
C1149 VDD1.n13 VSUBS 0.037194f
C1150 VDD1.n14 VSUBS 0.016662f
C1151 VDD1.n15 VSUBS 1.0987f
C1152 VDD1.n16 VSUBS 0.015736f
C1153 VDD1.t2 VSUBS 0.079933f
C1154 VDD1.n17 VSUBS 0.195579f
C1155 VDD1.n18 VSUBS 0.027979f
C1156 VDD1.n19 VSUBS 0.027895f
C1157 VDD1.n20 VSUBS 0.037194f
C1158 VDD1.n21 VSUBS 0.016662f
C1159 VDD1.n22 VSUBS 0.015736f
C1160 VDD1.n23 VSUBS 0.029284f
C1161 VDD1.n24 VSUBS 0.029284f
C1162 VDD1.n25 VSUBS 0.015736f
C1163 VDD1.n26 VSUBS 0.016662f
C1164 VDD1.n27 VSUBS 0.037194f
C1165 VDD1.n28 VSUBS 0.037194f
C1166 VDD1.n29 VSUBS 0.016662f
C1167 VDD1.n30 VSUBS 0.015736f
C1168 VDD1.n31 VSUBS 0.029284f
C1169 VDD1.n32 VSUBS 0.029284f
C1170 VDD1.n33 VSUBS 0.015736f
C1171 VDD1.n34 VSUBS 0.016662f
C1172 VDD1.n35 VSUBS 0.037194f
C1173 VDD1.n36 VSUBS 0.037194f
C1174 VDD1.n37 VSUBS 0.016662f
C1175 VDD1.n38 VSUBS 0.015736f
C1176 VDD1.n39 VSUBS 0.029284f
C1177 VDD1.n40 VSUBS 0.029284f
C1178 VDD1.n41 VSUBS 0.015736f
C1179 VDD1.n42 VSUBS 0.016662f
C1180 VDD1.n43 VSUBS 0.037194f
C1181 VDD1.n44 VSUBS 0.087511f
C1182 VDD1.n45 VSUBS 0.016662f
C1183 VDD1.n46 VSUBS 0.015736f
C1184 VDD1.n47 VSUBS 0.072089f
C1185 VDD1.n48 VSUBS 0.076909f
C1186 VDD1.n49 VSUBS 0.031434f
C1187 VDD1.n50 VSUBS 0.029284f
C1188 VDD1.n51 VSUBS 0.015736f
C1189 VDD1.n52 VSUBS 0.037194f
C1190 VDD1.n53 VSUBS 0.016199f
C1191 VDD1.n54 VSUBS 0.029284f
C1192 VDD1.n55 VSUBS 0.016662f
C1193 VDD1.n56 VSUBS 0.037194f
C1194 VDD1.n57 VSUBS 0.016662f
C1195 VDD1.n58 VSUBS 0.029284f
C1196 VDD1.n59 VSUBS 0.015736f
C1197 VDD1.n60 VSUBS 0.037194f
C1198 VDD1.n61 VSUBS 0.016662f
C1199 VDD1.n62 VSUBS 1.0987f
C1200 VDD1.n63 VSUBS 0.015736f
C1201 VDD1.t1 VSUBS 0.079933f
C1202 VDD1.n64 VSUBS 0.195579f
C1203 VDD1.n65 VSUBS 0.027979f
C1204 VDD1.n66 VSUBS 0.027895f
C1205 VDD1.n67 VSUBS 0.037194f
C1206 VDD1.n68 VSUBS 0.016662f
C1207 VDD1.n69 VSUBS 0.015736f
C1208 VDD1.n70 VSUBS 0.029284f
C1209 VDD1.n71 VSUBS 0.029284f
C1210 VDD1.n72 VSUBS 0.015736f
C1211 VDD1.n73 VSUBS 0.016662f
C1212 VDD1.n74 VSUBS 0.037194f
C1213 VDD1.n75 VSUBS 0.037194f
C1214 VDD1.n76 VSUBS 0.016662f
C1215 VDD1.n77 VSUBS 0.015736f
C1216 VDD1.n78 VSUBS 0.029284f
C1217 VDD1.n79 VSUBS 0.029284f
C1218 VDD1.n80 VSUBS 0.015736f
C1219 VDD1.n81 VSUBS 0.015736f
C1220 VDD1.n82 VSUBS 0.016662f
C1221 VDD1.n83 VSUBS 0.037194f
C1222 VDD1.n84 VSUBS 0.037194f
C1223 VDD1.n85 VSUBS 0.037194f
C1224 VDD1.n86 VSUBS 0.016199f
C1225 VDD1.n87 VSUBS 0.015736f
C1226 VDD1.n88 VSUBS 0.029284f
C1227 VDD1.n89 VSUBS 0.029284f
C1228 VDD1.n90 VSUBS 0.015736f
C1229 VDD1.n91 VSUBS 0.016662f
C1230 VDD1.n92 VSUBS 0.037194f
C1231 VDD1.n93 VSUBS 0.087511f
C1232 VDD1.n94 VSUBS 0.016662f
C1233 VDD1.n95 VSUBS 0.015736f
C1234 VDD1.n96 VSUBS 0.072089f
C1235 VDD1.n97 VSUBS 0.075886f
C1236 VDD1.t5 VSUBS 0.216369f
C1237 VDD1.t0 VSUBS 0.216369f
C1238 VDD1.n98 VSUBS 1.62672f
C1239 VDD1.n99 VSUBS 3.72311f
C1240 VDD1.t4 VSUBS 0.216369f
C1241 VDD1.t3 VSUBS 0.216369f
C1242 VDD1.n100 VSUBS 1.61886f
C1243 VDD1.n101 VSUBS 3.52474f
C1244 VP.t1 VSUBS 2.70236f
C1245 VP.n0 VSUBS 1.09706f
C1246 VP.n1 VSUBS 0.032705f
C1247 VP.n2 VSUBS 0.027504f
C1248 VP.n3 VSUBS 0.032705f
C1249 VP.t0 VSUBS 2.70236f
C1250 VP.n4 VSUBS 0.96418f
C1251 VP.n5 VSUBS 0.032705f
C1252 VP.n6 VSUBS 0.027504f
C1253 VP.n7 VSUBS 0.032705f
C1254 VP.t4 VSUBS 2.70236f
C1255 VP.n8 VSUBS 1.09706f
C1256 VP.t3 VSUBS 2.70236f
C1257 VP.n9 VSUBS 1.09706f
C1258 VP.n10 VSUBS 0.032705f
C1259 VP.n11 VSUBS 0.027504f
C1260 VP.n12 VSUBS 0.032705f
C1261 VP.t2 VSUBS 2.70236f
C1262 VP.n13 VSUBS 1.07283f
C1263 VP.t5 VSUBS 3.09243f
C1264 VP.n14 VSUBS 1.01938f
C1265 VP.n15 VSUBS 0.381572f
C1266 VP.n16 VSUBS 0.045907f
C1267 VP.n17 VSUBS 0.060953f
C1268 VP.n18 VSUBS 0.066044f
C1269 VP.n19 VSUBS 0.032705f
C1270 VP.n20 VSUBS 0.032705f
C1271 VP.n21 VSUBS 0.032705f
C1272 VP.n22 VSUBS 0.06289f
C1273 VP.n23 VSUBS 0.060953f
C1274 VP.n24 VSUBS 0.051925f
C1275 VP.n25 VSUBS 0.052784f
C1276 VP.n26 VSUBS 1.82764f
C1277 VP.n27 VSUBS 1.85142f
C1278 VP.n28 VSUBS 0.052784f
C1279 VP.n29 VSUBS 0.051925f
C1280 VP.n30 VSUBS 0.060953f
C1281 VP.n31 VSUBS 0.06289f
C1282 VP.n32 VSUBS 0.032705f
C1283 VP.n33 VSUBS 0.032705f
C1284 VP.n34 VSUBS 0.032705f
C1285 VP.n35 VSUBS 0.066044f
C1286 VP.n36 VSUBS 0.060953f
C1287 VP.n37 VSUBS 0.045907f
C1288 VP.n38 VSUBS 0.032705f
C1289 VP.n39 VSUBS 0.032705f
C1290 VP.n40 VSUBS 0.045907f
C1291 VP.n41 VSUBS 0.060953f
C1292 VP.n42 VSUBS 0.066044f
C1293 VP.n43 VSUBS 0.032705f
C1294 VP.n44 VSUBS 0.032705f
C1295 VP.n45 VSUBS 0.032705f
C1296 VP.n46 VSUBS 0.06289f
C1297 VP.n47 VSUBS 0.060953f
C1298 VP.n48 VSUBS 0.051925f
C1299 VP.n49 VSUBS 0.052784f
C1300 VP.n50 VSUBS 0.075376f
.ends

