* NGSPICE file created from diff_pair_sample_0273.ext - technology: sky130A

.subckt diff_pair_sample_0273 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X1 VDD1.t7 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X2 VDD1.t6 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X3 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=4.6215 ps=24.48 w=11.85 l=2.26
X4 VTAIL.t14 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X5 VDD2.t5 VN.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=4.6215 ps=24.48 w=11.85 l=2.26
X6 VTAIL.t3 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=1.95525 ps=12.18 w=11.85 l=2.26
X7 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=0 ps=0 w=11.85 l=2.26
X8 VTAIL.t7 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X9 VDD2.t4 VN.t3 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=4.6215 ps=24.48 w=11.85 l=2.26
X10 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=0 ps=0 w=11.85 l=2.26
X11 VTAIL.t15 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=1.95525 ps=12.18 w=11.85 l=2.26
X12 VTAIL.t10 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X13 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=4.6215 ps=24.48 w=11.85 l=2.26
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=0 ps=0 w=11.85 l=2.26
X15 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=1.95525 ps=12.18 w=11.85 l=2.26
X16 VDD2.t1 VN.t6 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X17 VTAIL.t6 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.95525 pd=12.18 as=1.95525 ps=12.18 w=11.85 l=2.26
X18 VTAIL.t8 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=1.95525 ps=12.18 w=11.85 l=2.26
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6215 pd=24.48 as=0 ps=0 w=11.85 l=2.26
R0 VN.n47 VN.n25 161.3
R1 VN.n46 VN.n45 161.3
R2 VN.n44 VN.n26 161.3
R3 VN.n43 VN.n42 161.3
R4 VN.n41 VN.n27 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n28 161.3
R7 VN.n36 VN.n35 161.3
R8 VN.n34 VN.n29 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n22 VN.n0 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n1 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n2 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n12 VN.n3 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n6 VN.t7 160.131
R21 VN.n31 VN.t3 160.131
R22 VN.n5 VN.t6 126.365
R23 VN.n15 VN.t5 126.365
R24 VN.n23 VN.t2 126.365
R25 VN.n30 VN.t1 126.365
R26 VN.n40 VN.t0 126.365
R27 VN.n48 VN.t4 126.365
R28 VN.n24 VN.n23 91.9169
R29 VN.n49 VN.n48 91.9169
R30 VN.n6 VN.n5 56.8068
R31 VN.n31 VN.n30 56.8068
R32 VN VN.n49 49.5436
R33 VN.n21 VN.n1 49.2348
R34 VN.n46 VN.n26 49.2348
R35 VN.n10 VN.n9 40.4934
R36 VN.n10 VN.n3 40.4934
R37 VN.n35 VN.n34 40.4934
R38 VN.n35 VN.n28 40.4934
R39 VN.n17 VN.n1 31.752
R40 VN.n42 VN.n26 31.752
R41 VN.n9 VN.n8 24.4675
R42 VN.n14 VN.n3 24.4675
R43 VN.n17 VN.n16 24.4675
R44 VN.n22 VN.n21 24.4675
R45 VN.n34 VN.n33 24.4675
R46 VN.n42 VN.n41 24.4675
R47 VN.n39 VN.n28 24.4675
R48 VN.n47 VN.n46 24.4675
R49 VN.n23 VN.n22 18.8401
R50 VN.n48 VN.n47 18.8401
R51 VN.n8 VN.n5 14.436
R52 VN.n15 VN.n14 14.436
R53 VN.n33 VN.n30 14.436
R54 VN.n40 VN.n39 14.436
R55 VN.n16 VN.n15 10.032
R56 VN.n41 VN.n40 10.032
R57 VN.n32 VN.n31 9.08053
R58 VN.n7 VN.n6 9.08053
R59 VN.n49 VN.n25 0.278367
R60 VN.n24 VN.n0 0.278367
R61 VN.n45 VN.n25 0.189894
R62 VN.n45 VN.n44 0.189894
R63 VN.n44 VN.n43 0.189894
R64 VN.n43 VN.n27 0.189894
R65 VN.n38 VN.n27 0.189894
R66 VN.n38 VN.n37 0.189894
R67 VN.n37 VN.n36 0.189894
R68 VN.n36 VN.n29 0.189894
R69 VN.n32 VN.n29 0.189894
R70 VN.n7 VN.n4 0.189894
R71 VN.n11 VN.n4 0.189894
R72 VN.n12 VN.n11 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n13 VN.n2 0.189894
R75 VN.n18 VN.n2 0.189894
R76 VN.n19 VN.n18 0.189894
R77 VN.n20 VN.n19 0.189894
R78 VN.n20 VN.n0 0.189894
R79 VN VN.n24 0.153454
R80 VTAIL.n11 VTAIL.t3 48.7176
R81 VTAIL.n10 VTAIL.t13 48.7176
R82 VTAIL.n7 VTAIL.t15 48.7176
R83 VTAIL.n15 VTAIL.t9 48.7174
R84 VTAIL.n2 VTAIL.t8 48.7174
R85 VTAIL.n3 VTAIL.t5 48.7174
R86 VTAIL.n6 VTAIL.t1 48.7174
R87 VTAIL.n14 VTAIL.t2 48.7174
R88 VTAIL.n13 VTAIL.n12 47.0467
R89 VTAIL.n9 VTAIL.n8 47.0467
R90 VTAIL.n1 VTAIL.n0 47.0465
R91 VTAIL.n5 VTAIL.n4 47.0465
R92 VTAIL.n15 VTAIL.n14 24.8152
R93 VTAIL.n7 VTAIL.n6 24.8152
R94 VTAIL.n9 VTAIL.n7 2.23326
R95 VTAIL.n10 VTAIL.n9 2.23326
R96 VTAIL.n13 VTAIL.n11 2.23326
R97 VTAIL.n14 VTAIL.n13 2.23326
R98 VTAIL.n6 VTAIL.n5 2.23326
R99 VTAIL.n5 VTAIL.n3 2.23326
R100 VTAIL.n2 VTAIL.n1 2.23326
R101 VTAIL VTAIL.n15 2.17507
R102 VTAIL.n0 VTAIL.t11 1.67139
R103 VTAIL.n0 VTAIL.t10 1.67139
R104 VTAIL.n4 VTAIL.t0 1.67139
R105 VTAIL.n4 VTAIL.t7 1.67139
R106 VTAIL.n12 VTAIL.t4 1.67139
R107 VTAIL.n12 VTAIL.t6 1.67139
R108 VTAIL.n8 VTAIL.t12 1.67139
R109 VTAIL.n8 VTAIL.t14 1.67139
R110 VTAIL.n11 VTAIL.n10 0.470328
R111 VTAIL.n3 VTAIL.n2 0.470328
R112 VTAIL VTAIL.n1 0.0586897
R113 VDD2.n2 VDD2.n1 64.7863
R114 VDD2.n2 VDD2.n0 64.7863
R115 VDD2 VDD2.n5 64.7835
R116 VDD2.n4 VDD2.n3 63.7255
R117 VDD2.n4 VDD2.n2 43.9782
R118 VDD2.n5 VDD2.t6 1.67139
R119 VDD2.n5 VDD2.t4 1.67139
R120 VDD2.n3 VDD2.t3 1.67139
R121 VDD2.n3 VDD2.t7 1.67139
R122 VDD2.n1 VDD2.t2 1.67139
R123 VDD2.n1 VDD2.t5 1.67139
R124 VDD2.n0 VDD2.t0 1.67139
R125 VDD2.n0 VDD2.t1 1.67139
R126 VDD2 VDD2.n4 1.17507
R127 B.n659 B.n658 585
R128 B.n661 B.n136 585
R129 B.n664 B.n663 585
R130 B.n665 B.n135 585
R131 B.n667 B.n666 585
R132 B.n669 B.n134 585
R133 B.n672 B.n671 585
R134 B.n673 B.n133 585
R135 B.n675 B.n674 585
R136 B.n677 B.n132 585
R137 B.n680 B.n679 585
R138 B.n681 B.n131 585
R139 B.n683 B.n682 585
R140 B.n685 B.n130 585
R141 B.n688 B.n687 585
R142 B.n689 B.n129 585
R143 B.n691 B.n690 585
R144 B.n693 B.n128 585
R145 B.n696 B.n695 585
R146 B.n697 B.n127 585
R147 B.n699 B.n698 585
R148 B.n701 B.n126 585
R149 B.n704 B.n703 585
R150 B.n705 B.n125 585
R151 B.n707 B.n706 585
R152 B.n709 B.n124 585
R153 B.n712 B.n711 585
R154 B.n713 B.n123 585
R155 B.n715 B.n714 585
R156 B.n717 B.n122 585
R157 B.n720 B.n719 585
R158 B.n721 B.n121 585
R159 B.n723 B.n722 585
R160 B.n725 B.n120 585
R161 B.n728 B.n727 585
R162 B.n729 B.n119 585
R163 B.n731 B.n730 585
R164 B.n733 B.n118 585
R165 B.n736 B.n735 585
R166 B.n737 B.n114 585
R167 B.n739 B.n738 585
R168 B.n741 B.n113 585
R169 B.n744 B.n743 585
R170 B.n745 B.n112 585
R171 B.n747 B.n746 585
R172 B.n749 B.n111 585
R173 B.n752 B.n751 585
R174 B.n753 B.n110 585
R175 B.n755 B.n754 585
R176 B.n757 B.n109 585
R177 B.n760 B.n759 585
R178 B.n762 B.n106 585
R179 B.n764 B.n763 585
R180 B.n766 B.n105 585
R181 B.n769 B.n768 585
R182 B.n770 B.n104 585
R183 B.n772 B.n771 585
R184 B.n774 B.n103 585
R185 B.n777 B.n776 585
R186 B.n778 B.n102 585
R187 B.n780 B.n779 585
R188 B.n782 B.n101 585
R189 B.n785 B.n784 585
R190 B.n786 B.n100 585
R191 B.n788 B.n787 585
R192 B.n790 B.n99 585
R193 B.n793 B.n792 585
R194 B.n794 B.n98 585
R195 B.n796 B.n795 585
R196 B.n798 B.n97 585
R197 B.n801 B.n800 585
R198 B.n802 B.n96 585
R199 B.n804 B.n803 585
R200 B.n806 B.n95 585
R201 B.n809 B.n808 585
R202 B.n810 B.n94 585
R203 B.n812 B.n811 585
R204 B.n814 B.n93 585
R205 B.n817 B.n816 585
R206 B.n818 B.n92 585
R207 B.n820 B.n819 585
R208 B.n822 B.n91 585
R209 B.n825 B.n824 585
R210 B.n826 B.n90 585
R211 B.n828 B.n827 585
R212 B.n830 B.n89 585
R213 B.n833 B.n832 585
R214 B.n834 B.n88 585
R215 B.n836 B.n835 585
R216 B.n838 B.n87 585
R217 B.n841 B.n840 585
R218 B.n842 B.n86 585
R219 B.n657 B.n84 585
R220 B.n845 B.n84 585
R221 B.n656 B.n83 585
R222 B.n846 B.n83 585
R223 B.n655 B.n82 585
R224 B.n847 B.n82 585
R225 B.n654 B.n653 585
R226 B.n653 B.n78 585
R227 B.n652 B.n77 585
R228 B.n853 B.n77 585
R229 B.n651 B.n76 585
R230 B.n854 B.n76 585
R231 B.n650 B.n75 585
R232 B.n855 B.n75 585
R233 B.n649 B.n648 585
R234 B.n648 B.n71 585
R235 B.n647 B.n70 585
R236 B.n861 B.n70 585
R237 B.n646 B.n69 585
R238 B.n862 B.n69 585
R239 B.n645 B.n68 585
R240 B.n863 B.n68 585
R241 B.n644 B.n643 585
R242 B.n643 B.n64 585
R243 B.n642 B.n63 585
R244 B.n869 B.n63 585
R245 B.n641 B.n62 585
R246 B.n870 B.n62 585
R247 B.n640 B.n61 585
R248 B.n871 B.n61 585
R249 B.n639 B.n638 585
R250 B.n638 B.n57 585
R251 B.n637 B.n56 585
R252 B.n877 B.n56 585
R253 B.n636 B.n55 585
R254 B.n878 B.n55 585
R255 B.n635 B.n54 585
R256 B.n879 B.n54 585
R257 B.n634 B.n633 585
R258 B.n633 B.n50 585
R259 B.n632 B.n49 585
R260 B.n885 B.n49 585
R261 B.n631 B.n48 585
R262 B.n886 B.n48 585
R263 B.n630 B.n47 585
R264 B.n887 B.n47 585
R265 B.n629 B.n628 585
R266 B.n628 B.n43 585
R267 B.n627 B.n42 585
R268 B.n893 B.n42 585
R269 B.n626 B.n41 585
R270 B.n894 B.n41 585
R271 B.n625 B.n40 585
R272 B.n895 B.n40 585
R273 B.n624 B.n623 585
R274 B.n623 B.n36 585
R275 B.n622 B.n35 585
R276 B.n901 B.n35 585
R277 B.n621 B.n34 585
R278 B.n902 B.n34 585
R279 B.n620 B.n33 585
R280 B.n903 B.n33 585
R281 B.n619 B.n618 585
R282 B.n618 B.n29 585
R283 B.n617 B.n28 585
R284 B.n909 B.n28 585
R285 B.n616 B.n27 585
R286 B.n910 B.n27 585
R287 B.n615 B.n26 585
R288 B.n911 B.n26 585
R289 B.n614 B.n613 585
R290 B.n613 B.n22 585
R291 B.n612 B.n21 585
R292 B.n917 B.n21 585
R293 B.n611 B.n20 585
R294 B.n918 B.n20 585
R295 B.n610 B.n19 585
R296 B.n919 B.n19 585
R297 B.n609 B.n608 585
R298 B.n608 B.n15 585
R299 B.n607 B.n14 585
R300 B.n925 B.n14 585
R301 B.n606 B.n13 585
R302 B.n926 B.n13 585
R303 B.n605 B.n12 585
R304 B.n927 B.n12 585
R305 B.n604 B.n603 585
R306 B.n603 B.n8 585
R307 B.n602 B.n7 585
R308 B.n933 B.n7 585
R309 B.n601 B.n6 585
R310 B.n934 B.n6 585
R311 B.n600 B.n5 585
R312 B.n935 B.n5 585
R313 B.n599 B.n598 585
R314 B.n598 B.n4 585
R315 B.n597 B.n137 585
R316 B.n597 B.n596 585
R317 B.n587 B.n138 585
R318 B.n139 B.n138 585
R319 B.n589 B.n588 585
R320 B.n590 B.n589 585
R321 B.n586 B.n144 585
R322 B.n144 B.n143 585
R323 B.n585 B.n584 585
R324 B.n584 B.n583 585
R325 B.n146 B.n145 585
R326 B.n147 B.n146 585
R327 B.n576 B.n575 585
R328 B.n577 B.n576 585
R329 B.n574 B.n152 585
R330 B.n152 B.n151 585
R331 B.n573 B.n572 585
R332 B.n572 B.n571 585
R333 B.n154 B.n153 585
R334 B.n155 B.n154 585
R335 B.n564 B.n563 585
R336 B.n565 B.n564 585
R337 B.n562 B.n160 585
R338 B.n160 B.n159 585
R339 B.n561 B.n560 585
R340 B.n560 B.n559 585
R341 B.n162 B.n161 585
R342 B.n163 B.n162 585
R343 B.n552 B.n551 585
R344 B.n553 B.n552 585
R345 B.n550 B.n168 585
R346 B.n168 B.n167 585
R347 B.n549 B.n548 585
R348 B.n548 B.n547 585
R349 B.n170 B.n169 585
R350 B.n171 B.n170 585
R351 B.n540 B.n539 585
R352 B.n541 B.n540 585
R353 B.n538 B.n175 585
R354 B.n179 B.n175 585
R355 B.n537 B.n536 585
R356 B.n536 B.n535 585
R357 B.n177 B.n176 585
R358 B.n178 B.n177 585
R359 B.n528 B.n527 585
R360 B.n529 B.n528 585
R361 B.n526 B.n184 585
R362 B.n184 B.n183 585
R363 B.n525 B.n524 585
R364 B.n524 B.n523 585
R365 B.n186 B.n185 585
R366 B.n187 B.n186 585
R367 B.n516 B.n515 585
R368 B.n517 B.n516 585
R369 B.n514 B.n191 585
R370 B.n195 B.n191 585
R371 B.n513 B.n512 585
R372 B.n512 B.n511 585
R373 B.n193 B.n192 585
R374 B.n194 B.n193 585
R375 B.n504 B.n503 585
R376 B.n505 B.n504 585
R377 B.n502 B.n200 585
R378 B.n200 B.n199 585
R379 B.n501 B.n500 585
R380 B.n500 B.n499 585
R381 B.n202 B.n201 585
R382 B.n203 B.n202 585
R383 B.n492 B.n491 585
R384 B.n493 B.n492 585
R385 B.n490 B.n208 585
R386 B.n208 B.n207 585
R387 B.n489 B.n488 585
R388 B.n488 B.n487 585
R389 B.n210 B.n209 585
R390 B.n211 B.n210 585
R391 B.n480 B.n479 585
R392 B.n481 B.n480 585
R393 B.n478 B.n216 585
R394 B.n216 B.n215 585
R395 B.n477 B.n476 585
R396 B.n476 B.n475 585
R397 B.n218 B.n217 585
R398 B.n219 B.n218 585
R399 B.n468 B.n467 585
R400 B.n469 B.n468 585
R401 B.n466 B.n224 585
R402 B.n224 B.n223 585
R403 B.n465 B.n464 585
R404 B.n464 B.n463 585
R405 B.n460 B.n228 585
R406 B.n459 B.n458 585
R407 B.n456 B.n229 585
R408 B.n456 B.n227 585
R409 B.n455 B.n454 585
R410 B.n453 B.n452 585
R411 B.n451 B.n231 585
R412 B.n449 B.n448 585
R413 B.n447 B.n232 585
R414 B.n446 B.n445 585
R415 B.n443 B.n233 585
R416 B.n441 B.n440 585
R417 B.n439 B.n234 585
R418 B.n438 B.n437 585
R419 B.n435 B.n235 585
R420 B.n433 B.n432 585
R421 B.n431 B.n236 585
R422 B.n430 B.n429 585
R423 B.n427 B.n237 585
R424 B.n425 B.n424 585
R425 B.n423 B.n238 585
R426 B.n422 B.n421 585
R427 B.n419 B.n239 585
R428 B.n417 B.n416 585
R429 B.n415 B.n240 585
R430 B.n414 B.n413 585
R431 B.n411 B.n241 585
R432 B.n409 B.n408 585
R433 B.n407 B.n242 585
R434 B.n406 B.n405 585
R435 B.n403 B.n243 585
R436 B.n401 B.n400 585
R437 B.n399 B.n244 585
R438 B.n398 B.n397 585
R439 B.n395 B.n245 585
R440 B.n393 B.n392 585
R441 B.n391 B.n246 585
R442 B.n390 B.n389 585
R443 B.n387 B.n247 585
R444 B.n385 B.n384 585
R445 B.n383 B.n248 585
R446 B.n382 B.n381 585
R447 B.n379 B.n378 585
R448 B.n377 B.n376 585
R449 B.n375 B.n253 585
R450 B.n373 B.n372 585
R451 B.n371 B.n254 585
R452 B.n370 B.n369 585
R453 B.n367 B.n255 585
R454 B.n365 B.n364 585
R455 B.n363 B.n256 585
R456 B.n362 B.n361 585
R457 B.n359 B.n358 585
R458 B.n357 B.n356 585
R459 B.n355 B.n261 585
R460 B.n353 B.n352 585
R461 B.n351 B.n262 585
R462 B.n350 B.n349 585
R463 B.n347 B.n263 585
R464 B.n345 B.n344 585
R465 B.n343 B.n264 585
R466 B.n342 B.n341 585
R467 B.n339 B.n265 585
R468 B.n337 B.n336 585
R469 B.n335 B.n266 585
R470 B.n334 B.n333 585
R471 B.n331 B.n267 585
R472 B.n329 B.n328 585
R473 B.n327 B.n268 585
R474 B.n326 B.n325 585
R475 B.n323 B.n269 585
R476 B.n321 B.n320 585
R477 B.n319 B.n270 585
R478 B.n318 B.n317 585
R479 B.n315 B.n271 585
R480 B.n313 B.n312 585
R481 B.n311 B.n272 585
R482 B.n310 B.n309 585
R483 B.n307 B.n273 585
R484 B.n305 B.n304 585
R485 B.n303 B.n274 585
R486 B.n302 B.n301 585
R487 B.n299 B.n275 585
R488 B.n297 B.n296 585
R489 B.n295 B.n276 585
R490 B.n294 B.n293 585
R491 B.n291 B.n277 585
R492 B.n289 B.n288 585
R493 B.n287 B.n278 585
R494 B.n286 B.n285 585
R495 B.n283 B.n279 585
R496 B.n281 B.n280 585
R497 B.n226 B.n225 585
R498 B.n227 B.n226 585
R499 B.n462 B.n461 585
R500 B.n463 B.n462 585
R501 B.n222 B.n221 585
R502 B.n223 B.n222 585
R503 B.n471 B.n470 585
R504 B.n470 B.n469 585
R505 B.n472 B.n220 585
R506 B.n220 B.n219 585
R507 B.n474 B.n473 585
R508 B.n475 B.n474 585
R509 B.n214 B.n213 585
R510 B.n215 B.n214 585
R511 B.n483 B.n482 585
R512 B.n482 B.n481 585
R513 B.n484 B.n212 585
R514 B.n212 B.n211 585
R515 B.n486 B.n485 585
R516 B.n487 B.n486 585
R517 B.n206 B.n205 585
R518 B.n207 B.n206 585
R519 B.n495 B.n494 585
R520 B.n494 B.n493 585
R521 B.n496 B.n204 585
R522 B.n204 B.n203 585
R523 B.n498 B.n497 585
R524 B.n499 B.n498 585
R525 B.n198 B.n197 585
R526 B.n199 B.n198 585
R527 B.n507 B.n506 585
R528 B.n506 B.n505 585
R529 B.n508 B.n196 585
R530 B.n196 B.n194 585
R531 B.n510 B.n509 585
R532 B.n511 B.n510 585
R533 B.n190 B.n189 585
R534 B.n195 B.n190 585
R535 B.n519 B.n518 585
R536 B.n518 B.n517 585
R537 B.n520 B.n188 585
R538 B.n188 B.n187 585
R539 B.n522 B.n521 585
R540 B.n523 B.n522 585
R541 B.n182 B.n181 585
R542 B.n183 B.n182 585
R543 B.n531 B.n530 585
R544 B.n530 B.n529 585
R545 B.n532 B.n180 585
R546 B.n180 B.n178 585
R547 B.n534 B.n533 585
R548 B.n535 B.n534 585
R549 B.n174 B.n173 585
R550 B.n179 B.n174 585
R551 B.n543 B.n542 585
R552 B.n542 B.n541 585
R553 B.n544 B.n172 585
R554 B.n172 B.n171 585
R555 B.n546 B.n545 585
R556 B.n547 B.n546 585
R557 B.n166 B.n165 585
R558 B.n167 B.n166 585
R559 B.n555 B.n554 585
R560 B.n554 B.n553 585
R561 B.n556 B.n164 585
R562 B.n164 B.n163 585
R563 B.n558 B.n557 585
R564 B.n559 B.n558 585
R565 B.n158 B.n157 585
R566 B.n159 B.n158 585
R567 B.n567 B.n566 585
R568 B.n566 B.n565 585
R569 B.n568 B.n156 585
R570 B.n156 B.n155 585
R571 B.n570 B.n569 585
R572 B.n571 B.n570 585
R573 B.n150 B.n149 585
R574 B.n151 B.n150 585
R575 B.n579 B.n578 585
R576 B.n578 B.n577 585
R577 B.n580 B.n148 585
R578 B.n148 B.n147 585
R579 B.n582 B.n581 585
R580 B.n583 B.n582 585
R581 B.n142 B.n141 585
R582 B.n143 B.n142 585
R583 B.n592 B.n591 585
R584 B.n591 B.n590 585
R585 B.n593 B.n140 585
R586 B.n140 B.n139 585
R587 B.n595 B.n594 585
R588 B.n596 B.n595 585
R589 B.n2 B.n0 585
R590 B.n4 B.n2 585
R591 B.n3 B.n1 585
R592 B.n934 B.n3 585
R593 B.n932 B.n931 585
R594 B.n933 B.n932 585
R595 B.n930 B.n9 585
R596 B.n9 B.n8 585
R597 B.n929 B.n928 585
R598 B.n928 B.n927 585
R599 B.n11 B.n10 585
R600 B.n926 B.n11 585
R601 B.n924 B.n923 585
R602 B.n925 B.n924 585
R603 B.n922 B.n16 585
R604 B.n16 B.n15 585
R605 B.n921 B.n920 585
R606 B.n920 B.n919 585
R607 B.n18 B.n17 585
R608 B.n918 B.n18 585
R609 B.n916 B.n915 585
R610 B.n917 B.n916 585
R611 B.n914 B.n23 585
R612 B.n23 B.n22 585
R613 B.n913 B.n912 585
R614 B.n912 B.n911 585
R615 B.n25 B.n24 585
R616 B.n910 B.n25 585
R617 B.n908 B.n907 585
R618 B.n909 B.n908 585
R619 B.n906 B.n30 585
R620 B.n30 B.n29 585
R621 B.n905 B.n904 585
R622 B.n904 B.n903 585
R623 B.n32 B.n31 585
R624 B.n902 B.n32 585
R625 B.n900 B.n899 585
R626 B.n901 B.n900 585
R627 B.n898 B.n37 585
R628 B.n37 B.n36 585
R629 B.n897 B.n896 585
R630 B.n896 B.n895 585
R631 B.n39 B.n38 585
R632 B.n894 B.n39 585
R633 B.n892 B.n891 585
R634 B.n893 B.n892 585
R635 B.n890 B.n44 585
R636 B.n44 B.n43 585
R637 B.n889 B.n888 585
R638 B.n888 B.n887 585
R639 B.n46 B.n45 585
R640 B.n886 B.n46 585
R641 B.n884 B.n883 585
R642 B.n885 B.n884 585
R643 B.n882 B.n51 585
R644 B.n51 B.n50 585
R645 B.n881 B.n880 585
R646 B.n880 B.n879 585
R647 B.n53 B.n52 585
R648 B.n878 B.n53 585
R649 B.n876 B.n875 585
R650 B.n877 B.n876 585
R651 B.n874 B.n58 585
R652 B.n58 B.n57 585
R653 B.n873 B.n872 585
R654 B.n872 B.n871 585
R655 B.n60 B.n59 585
R656 B.n870 B.n60 585
R657 B.n868 B.n867 585
R658 B.n869 B.n868 585
R659 B.n866 B.n65 585
R660 B.n65 B.n64 585
R661 B.n865 B.n864 585
R662 B.n864 B.n863 585
R663 B.n67 B.n66 585
R664 B.n862 B.n67 585
R665 B.n860 B.n859 585
R666 B.n861 B.n860 585
R667 B.n858 B.n72 585
R668 B.n72 B.n71 585
R669 B.n857 B.n856 585
R670 B.n856 B.n855 585
R671 B.n74 B.n73 585
R672 B.n854 B.n74 585
R673 B.n852 B.n851 585
R674 B.n853 B.n852 585
R675 B.n850 B.n79 585
R676 B.n79 B.n78 585
R677 B.n849 B.n848 585
R678 B.n848 B.n847 585
R679 B.n81 B.n80 585
R680 B.n846 B.n81 585
R681 B.n844 B.n843 585
R682 B.n845 B.n844 585
R683 B.n937 B.n936 585
R684 B.n936 B.n935 585
R685 B.n462 B.n228 526.135
R686 B.n844 B.n86 526.135
R687 B.n464 B.n226 526.135
R688 B.n659 B.n84 526.135
R689 B.n257 B.t16 333.834
R690 B.n249 B.t12 333.834
R691 B.n107 B.t19 333.834
R692 B.n115 B.t8 333.834
R693 B.n660 B.n85 256.663
R694 B.n662 B.n85 256.663
R695 B.n668 B.n85 256.663
R696 B.n670 B.n85 256.663
R697 B.n676 B.n85 256.663
R698 B.n678 B.n85 256.663
R699 B.n684 B.n85 256.663
R700 B.n686 B.n85 256.663
R701 B.n692 B.n85 256.663
R702 B.n694 B.n85 256.663
R703 B.n700 B.n85 256.663
R704 B.n702 B.n85 256.663
R705 B.n708 B.n85 256.663
R706 B.n710 B.n85 256.663
R707 B.n716 B.n85 256.663
R708 B.n718 B.n85 256.663
R709 B.n724 B.n85 256.663
R710 B.n726 B.n85 256.663
R711 B.n732 B.n85 256.663
R712 B.n734 B.n85 256.663
R713 B.n740 B.n85 256.663
R714 B.n742 B.n85 256.663
R715 B.n748 B.n85 256.663
R716 B.n750 B.n85 256.663
R717 B.n756 B.n85 256.663
R718 B.n758 B.n85 256.663
R719 B.n765 B.n85 256.663
R720 B.n767 B.n85 256.663
R721 B.n773 B.n85 256.663
R722 B.n775 B.n85 256.663
R723 B.n781 B.n85 256.663
R724 B.n783 B.n85 256.663
R725 B.n789 B.n85 256.663
R726 B.n791 B.n85 256.663
R727 B.n797 B.n85 256.663
R728 B.n799 B.n85 256.663
R729 B.n805 B.n85 256.663
R730 B.n807 B.n85 256.663
R731 B.n813 B.n85 256.663
R732 B.n815 B.n85 256.663
R733 B.n821 B.n85 256.663
R734 B.n823 B.n85 256.663
R735 B.n829 B.n85 256.663
R736 B.n831 B.n85 256.663
R737 B.n837 B.n85 256.663
R738 B.n839 B.n85 256.663
R739 B.n457 B.n227 256.663
R740 B.n230 B.n227 256.663
R741 B.n450 B.n227 256.663
R742 B.n444 B.n227 256.663
R743 B.n442 B.n227 256.663
R744 B.n436 B.n227 256.663
R745 B.n434 B.n227 256.663
R746 B.n428 B.n227 256.663
R747 B.n426 B.n227 256.663
R748 B.n420 B.n227 256.663
R749 B.n418 B.n227 256.663
R750 B.n412 B.n227 256.663
R751 B.n410 B.n227 256.663
R752 B.n404 B.n227 256.663
R753 B.n402 B.n227 256.663
R754 B.n396 B.n227 256.663
R755 B.n394 B.n227 256.663
R756 B.n388 B.n227 256.663
R757 B.n386 B.n227 256.663
R758 B.n380 B.n227 256.663
R759 B.n252 B.n227 256.663
R760 B.n374 B.n227 256.663
R761 B.n368 B.n227 256.663
R762 B.n366 B.n227 256.663
R763 B.n360 B.n227 256.663
R764 B.n260 B.n227 256.663
R765 B.n354 B.n227 256.663
R766 B.n348 B.n227 256.663
R767 B.n346 B.n227 256.663
R768 B.n340 B.n227 256.663
R769 B.n338 B.n227 256.663
R770 B.n332 B.n227 256.663
R771 B.n330 B.n227 256.663
R772 B.n324 B.n227 256.663
R773 B.n322 B.n227 256.663
R774 B.n316 B.n227 256.663
R775 B.n314 B.n227 256.663
R776 B.n308 B.n227 256.663
R777 B.n306 B.n227 256.663
R778 B.n300 B.n227 256.663
R779 B.n298 B.n227 256.663
R780 B.n292 B.n227 256.663
R781 B.n290 B.n227 256.663
R782 B.n284 B.n227 256.663
R783 B.n282 B.n227 256.663
R784 B.n462 B.n222 163.367
R785 B.n470 B.n222 163.367
R786 B.n470 B.n220 163.367
R787 B.n474 B.n220 163.367
R788 B.n474 B.n214 163.367
R789 B.n482 B.n214 163.367
R790 B.n482 B.n212 163.367
R791 B.n486 B.n212 163.367
R792 B.n486 B.n206 163.367
R793 B.n494 B.n206 163.367
R794 B.n494 B.n204 163.367
R795 B.n498 B.n204 163.367
R796 B.n498 B.n198 163.367
R797 B.n506 B.n198 163.367
R798 B.n506 B.n196 163.367
R799 B.n510 B.n196 163.367
R800 B.n510 B.n190 163.367
R801 B.n518 B.n190 163.367
R802 B.n518 B.n188 163.367
R803 B.n522 B.n188 163.367
R804 B.n522 B.n182 163.367
R805 B.n530 B.n182 163.367
R806 B.n530 B.n180 163.367
R807 B.n534 B.n180 163.367
R808 B.n534 B.n174 163.367
R809 B.n542 B.n174 163.367
R810 B.n542 B.n172 163.367
R811 B.n546 B.n172 163.367
R812 B.n546 B.n166 163.367
R813 B.n554 B.n166 163.367
R814 B.n554 B.n164 163.367
R815 B.n558 B.n164 163.367
R816 B.n558 B.n158 163.367
R817 B.n566 B.n158 163.367
R818 B.n566 B.n156 163.367
R819 B.n570 B.n156 163.367
R820 B.n570 B.n150 163.367
R821 B.n578 B.n150 163.367
R822 B.n578 B.n148 163.367
R823 B.n582 B.n148 163.367
R824 B.n582 B.n142 163.367
R825 B.n591 B.n142 163.367
R826 B.n591 B.n140 163.367
R827 B.n595 B.n140 163.367
R828 B.n595 B.n2 163.367
R829 B.n936 B.n2 163.367
R830 B.n936 B.n3 163.367
R831 B.n932 B.n3 163.367
R832 B.n932 B.n9 163.367
R833 B.n928 B.n9 163.367
R834 B.n928 B.n11 163.367
R835 B.n924 B.n11 163.367
R836 B.n924 B.n16 163.367
R837 B.n920 B.n16 163.367
R838 B.n920 B.n18 163.367
R839 B.n916 B.n18 163.367
R840 B.n916 B.n23 163.367
R841 B.n912 B.n23 163.367
R842 B.n912 B.n25 163.367
R843 B.n908 B.n25 163.367
R844 B.n908 B.n30 163.367
R845 B.n904 B.n30 163.367
R846 B.n904 B.n32 163.367
R847 B.n900 B.n32 163.367
R848 B.n900 B.n37 163.367
R849 B.n896 B.n37 163.367
R850 B.n896 B.n39 163.367
R851 B.n892 B.n39 163.367
R852 B.n892 B.n44 163.367
R853 B.n888 B.n44 163.367
R854 B.n888 B.n46 163.367
R855 B.n884 B.n46 163.367
R856 B.n884 B.n51 163.367
R857 B.n880 B.n51 163.367
R858 B.n880 B.n53 163.367
R859 B.n876 B.n53 163.367
R860 B.n876 B.n58 163.367
R861 B.n872 B.n58 163.367
R862 B.n872 B.n60 163.367
R863 B.n868 B.n60 163.367
R864 B.n868 B.n65 163.367
R865 B.n864 B.n65 163.367
R866 B.n864 B.n67 163.367
R867 B.n860 B.n67 163.367
R868 B.n860 B.n72 163.367
R869 B.n856 B.n72 163.367
R870 B.n856 B.n74 163.367
R871 B.n852 B.n74 163.367
R872 B.n852 B.n79 163.367
R873 B.n848 B.n79 163.367
R874 B.n848 B.n81 163.367
R875 B.n844 B.n81 163.367
R876 B.n458 B.n456 163.367
R877 B.n456 B.n455 163.367
R878 B.n452 B.n451 163.367
R879 B.n449 B.n232 163.367
R880 B.n445 B.n443 163.367
R881 B.n441 B.n234 163.367
R882 B.n437 B.n435 163.367
R883 B.n433 B.n236 163.367
R884 B.n429 B.n427 163.367
R885 B.n425 B.n238 163.367
R886 B.n421 B.n419 163.367
R887 B.n417 B.n240 163.367
R888 B.n413 B.n411 163.367
R889 B.n409 B.n242 163.367
R890 B.n405 B.n403 163.367
R891 B.n401 B.n244 163.367
R892 B.n397 B.n395 163.367
R893 B.n393 B.n246 163.367
R894 B.n389 B.n387 163.367
R895 B.n385 B.n248 163.367
R896 B.n381 B.n379 163.367
R897 B.n376 B.n375 163.367
R898 B.n373 B.n254 163.367
R899 B.n369 B.n367 163.367
R900 B.n365 B.n256 163.367
R901 B.n361 B.n359 163.367
R902 B.n356 B.n355 163.367
R903 B.n353 B.n262 163.367
R904 B.n349 B.n347 163.367
R905 B.n345 B.n264 163.367
R906 B.n341 B.n339 163.367
R907 B.n337 B.n266 163.367
R908 B.n333 B.n331 163.367
R909 B.n329 B.n268 163.367
R910 B.n325 B.n323 163.367
R911 B.n321 B.n270 163.367
R912 B.n317 B.n315 163.367
R913 B.n313 B.n272 163.367
R914 B.n309 B.n307 163.367
R915 B.n305 B.n274 163.367
R916 B.n301 B.n299 163.367
R917 B.n297 B.n276 163.367
R918 B.n293 B.n291 163.367
R919 B.n289 B.n278 163.367
R920 B.n285 B.n283 163.367
R921 B.n281 B.n226 163.367
R922 B.n464 B.n224 163.367
R923 B.n468 B.n224 163.367
R924 B.n468 B.n218 163.367
R925 B.n476 B.n218 163.367
R926 B.n476 B.n216 163.367
R927 B.n480 B.n216 163.367
R928 B.n480 B.n210 163.367
R929 B.n488 B.n210 163.367
R930 B.n488 B.n208 163.367
R931 B.n492 B.n208 163.367
R932 B.n492 B.n202 163.367
R933 B.n500 B.n202 163.367
R934 B.n500 B.n200 163.367
R935 B.n504 B.n200 163.367
R936 B.n504 B.n193 163.367
R937 B.n512 B.n193 163.367
R938 B.n512 B.n191 163.367
R939 B.n516 B.n191 163.367
R940 B.n516 B.n186 163.367
R941 B.n524 B.n186 163.367
R942 B.n524 B.n184 163.367
R943 B.n528 B.n184 163.367
R944 B.n528 B.n177 163.367
R945 B.n536 B.n177 163.367
R946 B.n536 B.n175 163.367
R947 B.n540 B.n175 163.367
R948 B.n540 B.n170 163.367
R949 B.n548 B.n170 163.367
R950 B.n548 B.n168 163.367
R951 B.n552 B.n168 163.367
R952 B.n552 B.n162 163.367
R953 B.n560 B.n162 163.367
R954 B.n560 B.n160 163.367
R955 B.n564 B.n160 163.367
R956 B.n564 B.n154 163.367
R957 B.n572 B.n154 163.367
R958 B.n572 B.n152 163.367
R959 B.n576 B.n152 163.367
R960 B.n576 B.n146 163.367
R961 B.n584 B.n146 163.367
R962 B.n584 B.n144 163.367
R963 B.n589 B.n144 163.367
R964 B.n589 B.n138 163.367
R965 B.n597 B.n138 163.367
R966 B.n598 B.n597 163.367
R967 B.n598 B.n5 163.367
R968 B.n6 B.n5 163.367
R969 B.n7 B.n6 163.367
R970 B.n603 B.n7 163.367
R971 B.n603 B.n12 163.367
R972 B.n13 B.n12 163.367
R973 B.n14 B.n13 163.367
R974 B.n608 B.n14 163.367
R975 B.n608 B.n19 163.367
R976 B.n20 B.n19 163.367
R977 B.n21 B.n20 163.367
R978 B.n613 B.n21 163.367
R979 B.n613 B.n26 163.367
R980 B.n27 B.n26 163.367
R981 B.n28 B.n27 163.367
R982 B.n618 B.n28 163.367
R983 B.n618 B.n33 163.367
R984 B.n34 B.n33 163.367
R985 B.n35 B.n34 163.367
R986 B.n623 B.n35 163.367
R987 B.n623 B.n40 163.367
R988 B.n41 B.n40 163.367
R989 B.n42 B.n41 163.367
R990 B.n628 B.n42 163.367
R991 B.n628 B.n47 163.367
R992 B.n48 B.n47 163.367
R993 B.n49 B.n48 163.367
R994 B.n633 B.n49 163.367
R995 B.n633 B.n54 163.367
R996 B.n55 B.n54 163.367
R997 B.n56 B.n55 163.367
R998 B.n638 B.n56 163.367
R999 B.n638 B.n61 163.367
R1000 B.n62 B.n61 163.367
R1001 B.n63 B.n62 163.367
R1002 B.n643 B.n63 163.367
R1003 B.n643 B.n68 163.367
R1004 B.n69 B.n68 163.367
R1005 B.n70 B.n69 163.367
R1006 B.n648 B.n70 163.367
R1007 B.n648 B.n75 163.367
R1008 B.n76 B.n75 163.367
R1009 B.n77 B.n76 163.367
R1010 B.n653 B.n77 163.367
R1011 B.n653 B.n82 163.367
R1012 B.n83 B.n82 163.367
R1013 B.n84 B.n83 163.367
R1014 B.n840 B.n838 163.367
R1015 B.n836 B.n88 163.367
R1016 B.n832 B.n830 163.367
R1017 B.n828 B.n90 163.367
R1018 B.n824 B.n822 163.367
R1019 B.n820 B.n92 163.367
R1020 B.n816 B.n814 163.367
R1021 B.n812 B.n94 163.367
R1022 B.n808 B.n806 163.367
R1023 B.n804 B.n96 163.367
R1024 B.n800 B.n798 163.367
R1025 B.n796 B.n98 163.367
R1026 B.n792 B.n790 163.367
R1027 B.n788 B.n100 163.367
R1028 B.n784 B.n782 163.367
R1029 B.n780 B.n102 163.367
R1030 B.n776 B.n774 163.367
R1031 B.n772 B.n104 163.367
R1032 B.n768 B.n766 163.367
R1033 B.n764 B.n106 163.367
R1034 B.n759 B.n757 163.367
R1035 B.n755 B.n110 163.367
R1036 B.n751 B.n749 163.367
R1037 B.n747 B.n112 163.367
R1038 B.n743 B.n741 163.367
R1039 B.n739 B.n114 163.367
R1040 B.n735 B.n733 163.367
R1041 B.n731 B.n119 163.367
R1042 B.n727 B.n725 163.367
R1043 B.n723 B.n121 163.367
R1044 B.n719 B.n717 163.367
R1045 B.n715 B.n123 163.367
R1046 B.n711 B.n709 163.367
R1047 B.n707 B.n125 163.367
R1048 B.n703 B.n701 163.367
R1049 B.n699 B.n127 163.367
R1050 B.n695 B.n693 163.367
R1051 B.n691 B.n129 163.367
R1052 B.n687 B.n685 163.367
R1053 B.n683 B.n131 163.367
R1054 B.n679 B.n677 163.367
R1055 B.n675 B.n133 163.367
R1056 B.n671 B.n669 163.367
R1057 B.n667 B.n135 163.367
R1058 B.n663 B.n661 163.367
R1059 B.n257 B.t18 123.665
R1060 B.n115 B.t10 123.665
R1061 B.n249 B.t15 123.65
R1062 B.n107 B.t20 123.65
R1063 B.n463 B.n227 88.0005
R1064 B.n845 B.n85 88.0005
R1065 B.n258 B.t17 73.4345
R1066 B.n116 B.t11 73.4345
R1067 B.n250 B.t14 73.4198
R1068 B.n108 B.t21 73.4198
R1069 B.n457 B.n228 71.676
R1070 B.n455 B.n230 71.676
R1071 B.n451 B.n450 71.676
R1072 B.n444 B.n232 71.676
R1073 B.n443 B.n442 71.676
R1074 B.n436 B.n234 71.676
R1075 B.n435 B.n434 71.676
R1076 B.n428 B.n236 71.676
R1077 B.n427 B.n426 71.676
R1078 B.n420 B.n238 71.676
R1079 B.n419 B.n418 71.676
R1080 B.n412 B.n240 71.676
R1081 B.n411 B.n410 71.676
R1082 B.n404 B.n242 71.676
R1083 B.n403 B.n402 71.676
R1084 B.n396 B.n244 71.676
R1085 B.n395 B.n394 71.676
R1086 B.n388 B.n246 71.676
R1087 B.n387 B.n386 71.676
R1088 B.n380 B.n248 71.676
R1089 B.n379 B.n252 71.676
R1090 B.n375 B.n374 71.676
R1091 B.n368 B.n254 71.676
R1092 B.n367 B.n366 71.676
R1093 B.n360 B.n256 71.676
R1094 B.n359 B.n260 71.676
R1095 B.n355 B.n354 71.676
R1096 B.n348 B.n262 71.676
R1097 B.n347 B.n346 71.676
R1098 B.n340 B.n264 71.676
R1099 B.n339 B.n338 71.676
R1100 B.n332 B.n266 71.676
R1101 B.n331 B.n330 71.676
R1102 B.n324 B.n268 71.676
R1103 B.n323 B.n322 71.676
R1104 B.n316 B.n270 71.676
R1105 B.n315 B.n314 71.676
R1106 B.n308 B.n272 71.676
R1107 B.n307 B.n306 71.676
R1108 B.n300 B.n274 71.676
R1109 B.n299 B.n298 71.676
R1110 B.n292 B.n276 71.676
R1111 B.n291 B.n290 71.676
R1112 B.n284 B.n278 71.676
R1113 B.n283 B.n282 71.676
R1114 B.n839 B.n86 71.676
R1115 B.n838 B.n837 71.676
R1116 B.n831 B.n88 71.676
R1117 B.n830 B.n829 71.676
R1118 B.n823 B.n90 71.676
R1119 B.n822 B.n821 71.676
R1120 B.n815 B.n92 71.676
R1121 B.n814 B.n813 71.676
R1122 B.n807 B.n94 71.676
R1123 B.n806 B.n805 71.676
R1124 B.n799 B.n96 71.676
R1125 B.n798 B.n797 71.676
R1126 B.n791 B.n98 71.676
R1127 B.n790 B.n789 71.676
R1128 B.n783 B.n100 71.676
R1129 B.n782 B.n781 71.676
R1130 B.n775 B.n102 71.676
R1131 B.n774 B.n773 71.676
R1132 B.n767 B.n104 71.676
R1133 B.n766 B.n765 71.676
R1134 B.n758 B.n106 71.676
R1135 B.n757 B.n756 71.676
R1136 B.n750 B.n110 71.676
R1137 B.n749 B.n748 71.676
R1138 B.n742 B.n112 71.676
R1139 B.n741 B.n740 71.676
R1140 B.n734 B.n114 71.676
R1141 B.n733 B.n732 71.676
R1142 B.n726 B.n119 71.676
R1143 B.n725 B.n724 71.676
R1144 B.n718 B.n121 71.676
R1145 B.n717 B.n716 71.676
R1146 B.n710 B.n123 71.676
R1147 B.n709 B.n708 71.676
R1148 B.n702 B.n125 71.676
R1149 B.n701 B.n700 71.676
R1150 B.n694 B.n127 71.676
R1151 B.n693 B.n692 71.676
R1152 B.n686 B.n129 71.676
R1153 B.n685 B.n684 71.676
R1154 B.n678 B.n131 71.676
R1155 B.n677 B.n676 71.676
R1156 B.n670 B.n133 71.676
R1157 B.n669 B.n668 71.676
R1158 B.n662 B.n135 71.676
R1159 B.n661 B.n660 71.676
R1160 B.n660 B.n659 71.676
R1161 B.n663 B.n662 71.676
R1162 B.n668 B.n667 71.676
R1163 B.n671 B.n670 71.676
R1164 B.n676 B.n675 71.676
R1165 B.n679 B.n678 71.676
R1166 B.n684 B.n683 71.676
R1167 B.n687 B.n686 71.676
R1168 B.n692 B.n691 71.676
R1169 B.n695 B.n694 71.676
R1170 B.n700 B.n699 71.676
R1171 B.n703 B.n702 71.676
R1172 B.n708 B.n707 71.676
R1173 B.n711 B.n710 71.676
R1174 B.n716 B.n715 71.676
R1175 B.n719 B.n718 71.676
R1176 B.n724 B.n723 71.676
R1177 B.n727 B.n726 71.676
R1178 B.n732 B.n731 71.676
R1179 B.n735 B.n734 71.676
R1180 B.n740 B.n739 71.676
R1181 B.n743 B.n742 71.676
R1182 B.n748 B.n747 71.676
R1183 B.n751 B.n750 71.676
R1184 B.n756 B.n755 71.676
R1185 B.n759 B.n758 71.676
R1186 B.n765 B.n764 71.676
R1187 B.n768 B.n767 71.676
R1188 B.n773 B.n772 71.676
R1189 B.n776 B.n775 71.676
R1190 B.n781 B.n780 71.676
R1191 B.n784 B.n783 71.676
R1192 B.n789 B.n788 71.676
R1193 B.n792 B.n791 71.676
R1194 B.n797 B.n796 71.676
R1195 B.n800 B.n799 71.676
R1196 B.n805 B.n804 71.676
R1197 B.n808 B.n807 71.676
R1198 B.n813 B.n812 71.676
R1199 B.n816 B.n815 71.676
R1200 B.n821 B.n820 71.676
R1201 B.n824 B.n823 71.676
R1202 B.n829 B.n828 71.676
R1203 B.n832 B.n831 71.676
R1204 B.n837 B.n836 71.676
R1205 B.n840 B.n839 71.676
R1206 B.n458 B.n457 71.676
R1207 B.n452 B.n230 71.676
R1208 B.n450 B.n449 71.676
R1209 B.n445 B.n444 71.676
R1210 B.n442 B.n441 71.676
R1211 B.n437 B.n436 71.676
R1212 B.n434 B.n433 71.676
R1213 B.n429 B.n428 71.676
R1214 B.n426 B.n425 71.676
R1215 B.n421 B.n420 71.676
R1216 B.n418 B.n417 71.676
R1217 B.n413 B.n412 71.676
R1218 B.n410 B.n409 71.676
R1219 B.n405 B.n404 71.676
R1220 B.n402 B.n401 71.676
R1221 B.n397 B.n396 71.676
R1222 B.n394 B.n393 71.676
R1223 B.n389 B.n388 71.676
R1224 B.n386 B.n385 71.676
R1225 B.n381 B.n380 71.676
R1226 B.n376 B.n252 71.676
R1227 B.n374 B.n373 71.676
R1228 B.n369 B.n368 71.676
R1229 B.n366 B.n365 71.676
R1230 B.n361 B.n360 71.676
R1231 B.n356 B.n260 71.676
R1232 B.n354 B.n353 71.676
R1233 B.n349 B.n348 71.676
R1234 B.n346 B.n345 71.676
R1235 B.n341 B.n340 71.676
R1236 B.n338 B.n337 71.676
R1237 B.n333 B.n332 71.676
R1238 B.n330 B.n329 71.676
R1239 B.n325 B.n324 71.676
R1240 B.n322 B.n321 71.676
R1241 B.n317 B.n316 71.676
R1242 B.n314 B.n313 71.676
R1243 B.n309 B.n308 71.676
R1244 B.n306 B.n305 71.676
R1245 B.n301 B.n300 71.676
R1246 B.n298 B.n297 71.676
R1247 B.n293 B.n292 71.676
R1248 B.n290 B.n289 71.676
R1249 B.n285 B.n284 71.676
R1250 B.n282 B.n281 71.676
R1251 B.n259 B.n258 59.5399
R1252 B.n251 B.n250 59.5399
R1253 B.n761 B.n108 59.5399
R1254 B.n117 B.n116 59.5399
R1255 B.n258 B.n257 50.2308
R1256 B.n250 B.n249 50.2308
R1257 B.n108 B.n107 50.2308
R1258 B.n116 B.n115 50.2308
R1259 B.n463 B.n223 43.6793
R1260 B.n469 B.n223 43.6793
R1261 B.n469 B.n219 43.6793
R1262 B.n475 B.n219 43.6793
R1263 B.n475 B.n215 43.6793
R1264 B.n481 B.n215 43.6793
R1265 B.n487 B.n211 43.6793
R1266 B.n487 B.n207 43.6793
R1267 B.n493 B.n207 43.6793
R1268 B.n493 B.n203 43.6793
R1269 B.n499 B.n203 43.6793
R1270 B.n499 B.n199 43.6793
R1271 B.n505 B.n199 43.6793
R1272 B.n505 B.n194 43.6793
R1273 B.n511 B.n194 43.6793
R1274 B.n511 B.n195 43.6793
R1275 B.n517 B.n187 43.6793
R1276 B.n523 B.n187 43.6793
R1277 B.n523 B.n183 43.6793
R1278 B.n529 B.n183 43.6793
R1279 B.n529 B.n178 43.6793
R1280 B.n535 B.n178 43.6793
R1281 B.n535 B.n179 43.6793
R1282 B.n541 B.n171 43.6793
R1283 B.n547 B.n171 43.6793
R1284 B.n547 B.n167 43.6793
R1285 B.n553 B.n167 43.6793
R1286 B.n553 B.n163 43.6793
R1287 B.n559 B.n163 43.6793
R1288 B.n565 B.n159 43.6793
R1289 B.n565 B.n155 43.6793
R1290 B.n571 B.n155 43.6793
R1291 B.n571 B.n151 43.6793
R1292 B.n577 B.n151 43.6793
R1293 B.n577 B.n147 43.6793
R1294 B.n583 B.n147 43.6793
R1295 B.n590 B.n143 43.6793
R1296 B.n590 B.n139 43.6793
R1297 B.n596 B.n139 43.6793
R1298 B.n596 B.n4 43.6793
R1299 B.n935 B.n4 43.6793
R1300 B.n935 B.n934 43.6793
R1301 B.n934 B.n933 43.6793
R1302 B.n933 B.n8 43.6793
R1303 B.n927 B.n8 43.6793
R1304 B.n927 B.n926 43.6793
R1305 B.n925 B.n15 43.6793
R1306 B.n919 B.n15 43.6793
R1307 B.n919 B.n918 43.6793
R1308 B.n918 B.n917 43.6793
R1309 B.n917 B.n22 43.6793
R1310 B.n911 B.n22 43.6793
R1311 B.n911 B.n910 43.6793
R1312 B.n909 B.n29 43.6793
R1313 B.n903 B.n29 43.6793
R1314 B.n903 B.n902 43.6793
R1315 B.n902 B.n901 43.6793
R1316 B.n901 B.n36 43.6793
R1317 B.n895 B.n36 43.6793
R1318 B.n894 B.n893 43.6793
R1319 B.n893 B.n43 43.6793
R1320 B.n887 B.n43 43.6793
R1321 B.n887 B.n886 43.6793
R1322 B.n886 B.n885 43.6793
R1323 B.n885 B.n50 43.6793
R1324 B.n879 B.n50 43.6793
R1325 B.n878 B.n877 43.6793
R1326 B.n877 B.n57 43.6793
R1327 B.n871 B.n57 43.6793
R1328 B.n871 B.n870 43.6793
R1329 B.n870 B.n869 43.6793
R1330 B.n869 B.n64 43.6793
R1331 B.n863 B.n64 43.6793
R1332 B.n863 B.n862 43.6793
R1333 B.n862 B.n861 43.6793
R1334 B.n861 B.n71 43.6793
R1335 B.n855 B.n854 43.6793
R1336 B.n854 B.n853 43.6793
R1337 B.n853 B.n78 43.6793
R1338 B.n847 B.n78 43.6793
R1339 B.n847 B.n846 43.6793
R1340 B.n846 B.n845 43.6793
R1341 B.n559 B.t7 42.3947
R1342 B.t4 B.n909 42.3947
R1343 B.n481 B.t13 39.8253
R1344 B.n855 B.t9 39.8253
R1345 B.n843 B.n842 34.1859
R1346 B.n658 B.n657 34.1859
R1347 B.n465 B.n225 34.1859
R1348 B.n461 B.n460 34.1859
R1349 B.n195 B.t1 32.1173
R1350 B.t2 B.n878 32.1173
R1351 B.n541 B.t0 28.2633
R1352 B.n895 B.t6 28.2633
R1353 B.n583 B.t5 25.6939
R1354 B.t3 B.n925 25.6939
R1355 B B.n937 18.0485
R1356 B.t5 B.n143 17.9859
R1357 B.n926 B.t3 17.9859
R1358 B.n179 B.t0 15.4166
R1359 B.t6 B.n894 15.4166
R1360 B.n517 B.t1 11.5625
R1361 B.n879 B.t2 11.5625
R1362 B.n842 B.n841 10.6151
R1363 B.n841 B.n87 10.6151
R1364 B.n835 B.n87 10.6151
R1365 B.n835 B.n834 10.6151
R1366 B.n834 B.n833 10.6151
R1367 B.n833 B.n89 10.6151
R1368 B.n827 B.n89 10.6151
R1369 B.n827 B.n826 10.6151
R1370 B.n826 B.n825 10.6151
R1371 B.n825 B.n91 10.6151
R1372 B.n819 B.n91 10.6151
R1373 B.n819 B.n818 10.6151
R1374 B.n818 B.n817 10.6151
R1375 B.n817 B.n93 10.6151
R1376 B.n811 B.n93 10.6151
R1377 B.n811 B.n810 10.6151
R1378 B.n810 B.n809 10.6151
R1379 B.n809 B.n95 10.6151
R1380 B.n803 B.n95 10.6151
R1381 B.n803 B.n802 10.6151
R1382 B.n802 B.n801 10.6151
R1383 B.n801 B.n97 10.6151
R1384 B.n795 B.n97 10.6151
R1385 B.n795 B.n794 10.6151
R1386 B.n794 B.n793 10.6151
R1387 B.n793 B.n99 10.6151
R1388 B.n787 B.n99 10.6151
R1389 B.n787 B.n786 10.6151
R1390 B.n786 B.n785 10.6151
R1391 B.n785 B.n101 10.6151
R1392 B.n779 B.n101 10.6151
R1393 B.n779 B.n778 10.6151
R1394 B.n778 B.n777 10.6151
R1395 B.n777 B.n103 10.6151
R1396 B.n771 B.n103 10.6151
R1397 B.n771 B.n770 10.6151
R1398 B.n770 B.n769 10.6151
R1399 B.n769 B.n105 10.6151
R1400 B.n763 B.n105 10.6151
R1401 B.n763 B.n762 10.6151
R1402 B.n760 B.n109 10.6151
R1403 B.n754 B.n109 10.6151
R1404 B.n754 B.n753 10.6151
R1405 B.n753 B.n752 10.6151
R1406 B.n752 B.n111 10.6151
R1407 B.n746 B.n111 10.6151
R1408 B.n746 B.n745 10.6151
R1409 B.n745 B.n744 10.6151
R1410 B.n744 B.n113 10.6151
R1411 B.n738 B.n737 10.6151
R1412 B.n737 B.n736 10.6151
R1413 B.n736 B.n118 10.6151
R1414 B.n730 B.n118 10.6151
R1415 B.n730 B.n729 10.6151
R1416 B.n729 B.n728 10.6151
R1417 B.n728 B.n120 10.6151
R1418 B.n722 B.n120 10.6151
R1419 B.n722 B.n721 10.6151
R1420 B.n721 B.n720 10.6151
R1421 B.n720 B.n122 10.6151
R1422 B.n714 B.n122 10.6151
R1423 B.n714 B.n713 10.6151
R1424 B.n713 B.n712 10.6151
R1425 B.n712 B.n124 10.6151
R1426 B.n706 B.n124 10.6151
R1427 B.n706 B.n705 10.6151
R1428 B.n705 B.n704 10.6151
R1429 B.n704 B.n126 10.6151
R1430 B.n698 B.n126 10.6151
R1431 B.n698 B.n697 10.6151
R1432 B.n697 B.n696 10.6151
R1433 B.n696 B.n128 10.6151
R1434 B.n690 B.n128 10.6151
R1435 B.n690 B.n689 10.6151
R1436 B.n689 B.n688 10.6151
R1437 B.n688 B.n130 10.6151
R1438 B.n682 B.n130 10.6151
R1439 B.n682 B.n681 10.6151
R1440 B.n681 B.n680 10.6151
R1441 B.n680 B.n132 10.6151
R1442 B.n674 B.n132 10.6151
R1443 B.n674 B.n673 10.6151
R1444 B.n673 B.n672 10.6151
R1445 B.n672 B.n134 10.6151
R1446 B.n666 B.n134 10.6151
R1447 B.n666 B.n665 10.6151
R1448 B.n665 B.n664 10.6151
R1449 B.n664 B.n136 10.6151
R1450 B.n658 B.n136 10.6151
R1451 B.n466 B.n465 10.6151
R1452 B.n467 B.n466 10.6151
R1453 B.n467 B.n217 10.6151
R1454 B.n477 B.n217 10.6151
R1455 B.n478 B.n477 10.6151
R1456 B.n479 B.n478 10.6151
R1457 B.n479 B.n209 10.6151
R1458 B.n489 B.n209 10.6151
R1459 B.n490 B.n489 10.6151
R1460 B.n491 B.n490 10.6151
R1461 B.n491 B.n201 10.6151
R1462 B.n501 B.n201 10.6151
R1463 B.n502 B.n501 10.6151
R1464 B.n503 B.n502 10.6151
R1465 B.n503 B.n192 10.6151
R1466 B.n513 B.n192 10.6151
R1467 B.n514 B.n513 10.6151
R1468 B.n515 B.n514 10.6151
R1469 B.n515 B.n185 10.6151
R1470 B.n525 B.n185 10.6151
R1471 B.n526 B.n525 10.6151
R1472 B.n527 B.n526 10.6151
R1473 B.n527 B.n176 10.6151
R1474 B.n537 B.n176 10.6151
R1475 B.n538 B.n537 10.6151
R1476 B.n539 B.n538 10.6151
R1477 B.n539 B.n169 10.6151
R1478 B.n549 B.n169 10.6151
R1479 B.n550 B.n549 10.6151
R1480 B.n551 B.n550 10.6151
R1481 B.n551 B.n161 10.6151
R1482 B.n561 B.n161 10.6151
R1483 B.n562 B.n561 10.6151
R1484 B.n563 B.n562 10.6151
R1485 B.n563 B.n153 10.6151
R1486 B.n573 B.n153 10.6151
R1487 B.n574 B.n573 10.6151
R1488 B.n575 B.n574 10.6151
R1489 B.n575 B.n145 10.6151
R1490 B.n585 B.n145 10.6151
R1491 B.n586 B.n585 10.6151
R1492 B.n588 B.n586 10.6151
R1493 B.n588 B.n587 10.6151
R1494 B.n587 B.n137 10.6151
R1495 B.n599 B.n137 10.6151
R1496 B.n600 B.n599 10.6151
R1497 B.n601 B.n600 10.6151
R1498 B.n602 B.n601 10.6151
R1499 B.n604 B.n602 10.6151
R1500 B.n605 B.n604 10.6151
R1501 B.n606 B.n605 10.6151
R1502 B.n607 B.n606 10.6151
R1503 B.n609 B.n607 10.6151
R1504 B.n610 B.n609 10.6151
R1505 B.n611 B.n610 10.6151
R1506 B.n612 B.n611 10.6151
R1507 B.n614 B.n612 10.6151
R1508 B.n615 B.n614 10.6151
R1509 B.n616 B.n615 10.6151
R1510 B.n617 B.n616 10.6151
R1511 B.n619 B.n617 10.6151
R1512 B.n620 B.n619 10.6151
R1513 B.n621 B.n620 10.6151
R1514 B.n622 B.n621 10.6151
R1515 B.n624 B.n622 10.6151
R1516 B.n625 B.n624 10.6151
R1517 B.n626 B.n625 10.6151
R1518 B.n627 B.n626 10.6151
R1519 B.n629 B.n627 10.6151
R1520 B.n630 B.n629 10.6151
R1521 B.n631 B.n630 10.6151
R1522 B.n632 B.n631 10.6151
R1523 B.n634 B.n632 10.6151
R1524 B.n635 B.n634 10.6151
R1525 B.n636 B.n635 10.6151
R1526 B.n637 B.n636 10.6151
R1527 B.n639 B.n637 10.6151
R1528 B.n640 B.n639 10.6151
R1529 B.n641 B.n640 10.6151
R1530 B.n642 B.n641 10.6151
R1531 B.n644 B.n642 10.6151
R1532 B.n645 B.n644 10.6151
R1533 B.n646 B.n645 10.6151
R1534 B.n647 B.n646 10.6151
R1535 B.n649 B.n647 10.6151
R1536 B.n650 B.n649 10.6151
R1537 B.n651 B.n650 10.6151
R1538 B.n652 B.n651 10.6151
R1539 B.n654 B.n652 10.6151
R1540 B.n655 B.n654 10.6151
R1541 B.n656 B.n655 10.6151
R1542 B.n657 B.n656 10.6151
R1543 B.n460 B.n459 10.6151
R1544 B.n459 B.n229 10.6151
R1545 B.n454 B.n229 10.6151
R1546 B.n454 B.n453 10.6151
R1547 B.n453 B.n231 10.6151
R1548 B.n448 B.n231 10.6151
R1549 B.n448 B.n447 10.6151
R1550 B.n447 B.n446 10.6151
R1551 B.n446 B.n233 10.6151
R1552 B.n440 B.n233 10.6151
R1553 B.n440 B.n439 10.6151
R1554 B.n439 B.n438 10.6151
R1555 B.n438 B.n235 10.6151
R1556 B.n432 B.n235 10.6151
R1557 B.n432 B.n431 10.6151
R1558 B.n431 B.n430 10.6151
R1559 B.n430 B.n237 10.6151
R1560 B.n424 B.n237 10.6151
R1561 B.n424 B.n423 10.6151
R1562 B.n423 B.n422 10.6151
R1563 B.n422 B.n239 10.6151
R1564 B.n416 B.n239 10.6151
R1565 B.n416 B.n415 10.6151
R1566 B.n415 B.n414 10.6151
R1567 B.n414 B.n241 10.6151
R1568 B.n408 B.n241 10.6151
R1569 B.n408 B.n407 10.6151
R1570 B.n407 B.n406 10.6151
R1571 B.n406 B.n243 10.6151
R1572 B.n400 B.n243 10.6151
R1573 B.n400 B.n399 10.6151
R1574 B.n399 B.n398 10.6151
R1575 B.n398 B.n245 10.6151
R1576 B.n392 B.n245 10.6151
R1577 B.n392 B.n391 10.6151
R1578 B.n391 B.n390 10.6151
R1579 B.n390 B.n247 10.6151
R1580 B.n384 B.n247 10.6151
R1581 B.n384 B.n383 10.6151
R1582 B.n383 B.n382 10.6151
R1583 B.n378 B.n377 10.6151
R1584 B.n377 B.n253 10.6151
R1585 B.n372 B.n253 10.6151
R1586 B.n372 B.n371 10.6151
R1587 B.n371 B.n370 10.6151
R1588 B.n370 B.n255 10.6151
R1589 B.n364 B.n255 10.6151
R1590 B.n364 B.n363 10.6151
R1591 B.n363 B.n362 10.6151
R1592 B.n358 B.n357 10.6151
R1593 B.n357 B.n261 10.6151
R1594 B.n352 B.n261 10.6151
R1595 B.n352 B.n351 10.6151
R1596 B.n351 B.n350 10.6151
R1597 B.n350 B.n263 10.6151
R1598 B.n344 B.n263 10.6151
R1599 B.n344 B.n343 10.6151
R1600 B.n343 B.n342 10.6151
R1601 B.n342 B.n265 10.6151
R1602 B.n336 B.n265 10.6151
R1603 B.n336 B.n335 10.6151
R1604 B.n335 B.n334 10.6151
R1605 B.n334 B.n267 10.6151
R1606 B.n328 B.n267 10.6151
R1607 B.n328 B.n327 10.6151
R1608 B.n327 B.n326 10.6151
R1609 B.n326 B.n269 10.6151
R1610 B.n320 B.n269 10.6151
R1611 B.n320 B.n319 10.6151
R1612 B.n319 B.n318 10.6151
R1613 B.n318 B.n271 10.6151
R1614 B.n312 B.n271 10.6151
R1615 B.n312 B.n311 10.6151
R1616 B.n311 B.n310 10.6151
R1617 B.n310 B.n273 10.6151
R1618 B.n304 B.n273 10.6151
R1619 B.n304 B.n303 10.6151
R1620 B.n303 B.n302 10.6151
R1621 B.n302 B.n275 10.6151
R1622 B.n296 B.n275 10.6151
R1623 B.n296 B.n295 10.6151
R1624 B.n295 B.n294 10.6151
R1625 B.n294 B.n277 10.6151
R1626 B.n288 B.n277 10.6151
R1627 B.n288 B.n287 10.6151
R1628 B.n287 B.n286 10.6151
R1629 B.n286 B.n279 10.6151
R1630 B.n280 B.n279 10.6151
R1631 B.n280 B.n225 10.6151
R1632 B.n461 B.n221 10.6151
R1633 B.n471 B.n221 10.6151
R1634 B.n472 B.n471 10.6151
R1635 B.n473 B.n472 10.6151
R1636 B.n473 B.n213 10.6151
R1637 B.n483 B.n213 10.6151
R1638 B.n484 B.n483 10.6151
R1639 B.n485 B.n484 10.6151
R1640 B.n485 B.n205 10.6151
R1641 B.n495 B.n205 10.6151
R1642 B.n496 B.n495 10.6151
R1643 B.n497 B.n496 10.6151
R1644 B.n497 B.n197 10.6151
R1645 B.n507 B.n197 10.6151
R1646 B.n508 B.n507 10.6151
R1647 B.n509 B.n508 10.6151
R1648 B.n509 B.n189 10.6151
R1649 B.n519 B.n189 10.6151
R1650 B.n520 B.n519 10.6151
R1651 B.n521 B.n520 10.6151
R1652 B.n521 B.n181 10.6151
R1653 B.n531 B.n181 10.6151
R1654 B.n532 B.n531 10.6151
R1655 B.n533 B.n532 10.6151
R1656 B.n533 B.n173 10.6151
R1657 B.n543 B.n173 10.6151
R1658 B.n544 B.n543 10.6151
R1659 B.n545 B.n544 10.6151
R1660 B.n545 B.n165 10.6151
R1661 B.n555 B.n165 10.6151
R1662 B.n556 B.n555 10.6151
R1663 B.n557 B.n556 10.6151
R1664 B.n557 B.n157 10.6151
R1665 B.n567 B.n157 10.6151
R1666 B.n568 B.n567 10.6151
R1667 B.n569 B.n568 10.6151
R1668 B.n569 B.n149 10.6151
R1669 B.n579 B.n149 10.6151
R1670 B.n580 B.n579 10.6151
R1671 B.n581 B.n580 10.6151
R1672 B.n581 B.n141 10.6151
R1673 B.n592 B.n141 10.6151
R1674 B.n593 B.n592 10.6151
R1675 B.n594 B.n593 10.6151
R1676 B.n594 B.n0 10.6151
R1677 B.n931 B.n1 10.6151
R1678 B.n931 B.n930 10.6151
R1679 B.n930 B.n929 10.6151
R1680 B.n929 B.n10 10.6151
R1681 B.n923 B.n10 10.6151
R1682 B.n923 B.n922 10.6151
R1683 B.n922 B.n921 10.6151
R1684 B.n921 B.n17 10.6151
R1685 B.n915 B.n17 10.6151
R1686 B.n915 B.n914 10.6151
R1687 B.n914 B.n913 10.6151
R1688 B.n913 B.n24 10.6151
R1689 B.n907 B.n24 10.6151
R1690 B.n907 B.n906 10.6151
R1691 B.n906 B.n905 10.6151
R1692 B.n905 B.n31 10.6151
R1693 B.n899 B.n31 10.6151
R1694 B.n899 B.n898 10.6151
R1695 B.n898 B.n897 10.6151
R1696 B.n897 B.n38 10.6151
R1697 B.n891 B.n38 10.6151
R1698 B.n891 B.n890 10.6151
R1699 B.n890 B.n889 10.6151
R1700 B.n889 B.n45 10.6151
R1701 B.n883 B.n45 10.6151
R1702 B.n883 B.n882 10.6151
R1703 B.n882 B.n881 10.6151
R1704 B.n881 B.n52 10.6151
R1705 B.n875 B.n52 10.6151
R1706 B.n875 B.n874 10.6151
R1707 B.n874 B.n873 10.6151
R1708 B.n873 B.n59 10.6151
R1709 B.n867 B.n59 10.6151
R1710 B.n867 B.n866 10.6151
R1711 B.n866 B.n865 10.6151
R1712 B.n865 B.n66 10.6151
R1713 B.n859 B.n66 10.6151
R1714 B.n859 B.n858 10.6151
R1715 B.n858 B.n857 10.6151
R1716 B.n857 B.n73 10.6151
R1717 B.n851 B.n73 10.6151
R1718 B.n851 B.n850 10.6151
R1719 B.n850 B.n849 10.6151
R1720 B.n849 B.n80 10.6151
R1721 B.n843 B.n80 10.6151
R1722 B.n762 B.n761 9.36635
R1723 B.n738 B.n117 9.36635
R1724 B.n382 B.n251 9.36635
R1725 B.n358 B.n259 9.36635
R1726 B.t13 B.n211 3.85451
R1727 B.t9 B.n71 3.85451
R1728 B.n937 B.n0 2.81026
R1729 B.n937 B.n1 2.81026
R1730 B.t7 B.n159 1.28517
R1731 B.n910 B.t4 1.28517
R1732 B.n761 B.n760 1.24928
R1733 B.n117 B.n113 1.24928
R1734 B.n378 B.n251 1.24928
R1735 B.n362 B.n259 1.24928
R1736 VP.n16 VP.n15 161.3
R1737 VP.n17 VP.n12 161.3
R1738 VP.n19 VP.n18 161.3
R1739 VP.n20 VP.n11 161.3
R1740 VP.n22 VP.n21 161.3
R1741 VP.n24 VP.n10 161.3
R1742 VP.n26 VP.n25 161.3
R1743 VP.n27 VP.n9 161.3
R1744 VP.n29 VP.n28 161.3
R1745 VP.n30 VP.n8 161.3
R1746 VP.n58 VP.n0 161.3
R1747 VP.n57 VP.n56 161.3
R1748 VP.n55 VP.n1 161.3
R1749 VP.n54 VP.n53 161.3
R1750 VP.n52 VP.n2 161.3
R1751 VP.n50 VP.n49 161.3
R1752 VP.n48 VP.n3 161.3
R1753 VP.n47 VP.n46 161.3
R1754 VP.n45 VP.n4 161.3
R1755 VP.n44 VP.n43 161.3
R1756 VP.n42 VP.n41 161.3
R1757 VP.n40 VP.n6 161.3
R1758 VP.n39 VP.n38 161.3
R1759 VP.n37 VP.n7 161.3
R1760 VP.n36 VP.n35 161.3
R1761 VP.n14 VP.t3 160.131
R1762 VP.n34 VP.t6 126.365
R1763 VP.n5 VP.t0 126.365
R1764 VP.n51 VP.t4 126.365
R1765 VP.n59 VP.t5 126.365
R1766 VP.n31 VP.t2 126.365
R1767 VP.n23 VP.t7 126.365
R1768 VP.n13 VP.t1 126.365
R1769 VP.n34 VP.n33 91.9169
R1770 VP.n60 VP.n59 91.9169
R1771 VP.n32 VP.n31 91.9169
R1772 VP.n14 VP.n13 56.8068
R1773 VP.n33 VP.n32 49.2647
R1774 VP.n39 VP.n7 49.2348
R1775 VP.n57 VP.n1 49.2348
R1776 VP.n29 VP.n9 49.2348
R1777 VP.n46 VP.n45 40.4934
R1778 VP.n46 VP.n3 40.4934
R1779 VP.n18 VP.n11 40.4934
R1780 VP.n18 VP.n17 40.4934
R1781 VP.n40 VP.n39 31.752
R1782 VP.n53 VP.n1 31.752
R1783 VP.n25 VP.n9 31.752
R1784 VP.n35 VP.n7 24.4675
R1785 VP.n41 VP.n40 24.4675
R1786 VP.n45 VP.n44 24.4675
R1787 VP.n50 VP.n3 24.4675
R1788 VP.n53 VP.n52 24.4675
R1789 VP.n58 VP.n57 24.4675
R1790 VP.n30 VP.n29 24.4675
R1791 VP.n22 VP.n11 24.4675
R1792 VP.n25 VP.n24 24.4675
R1793 VP.n17 VP.n16 24.4675
R1794 VP.n35 VP.n34 18.8401
R1795 VP.n59 VP.n58 18.8401
R1796 VP.n31 VP.n30 18.8401
R1797 VP.n44 VP.n5 14.436
R1798 VP.n51 VP.n50 14.436
R1799 VP.n23 VP.n22 14.436
R1800 VP.n16 VP.n13 14.436
R1801 VP.n41 VP.n5 10.032
R1802 VP.n52 VP.n51 10.032
R1803 VP.n24 VP.n23 10.032
R1804 VP.n15 VP.n14 9.08053
R1805 VP.n32 VP.n8 0.278367
R1806 VP.n36 VP.n33 0.278367
R1807 VP.n60 VP.n0 0.278367
R1808 VP.n15 VP.n12 0.189894
R1809 VP.n19 VP.n12 0.189894
R1810 VP.n20 VP.n19 0.189894
R1811 VP.n21 VP.n20 0.189894
R1812 VP.n21 VP.n10 0.189894
R1813 VP.n26 VP.n10 0.189894
R1814 VP.n27 VP.n26 0.189894
R1815 VP.n28 VP.n27 0.189894
R1816 VP.n28 VP.n8 0.189894
R1817 VP.n37 VP.n36 0.189894
R1818 VP.n38 VP.n37 0.189894
R1819 VP.n38 VP.n6 0.189894
R1820 VP.n42 VP.n6 0.189894
R1821 VP.n43 VP.n42 0.189894
R1822 VP.n43 VP.n4 0.189894
R1823 VP.n47 VP.n4 0.189894
R1824 VP.n48 VP.n47 0.189894
R1825 VP.n49 VP.n48 0.189894
R1826 VP.n49 VP.n2 0.189894
R1827 VP.n54 VP.n2 0.189894
R1828 VP.n55 VP.n54 0.189894
R1829 VP.n56 VP.n55 0.189894
R1830 VP.n56 VP.n0 0.189894
R1831 VP VP.n60 0.153454
R1832 VDD1 VDD1.n0 64.9
R1833 VDD1.n3 VDD1.n2 64.7863
R1834 VDD1.n3 VDD1.n1 64.7863
R1835 VDD1.n5 VDD1.n4 63.7253
R1836 VDD1.n5 VDD1.n3 44.5612
R1837 VDD1.n4 VDD1.t0 1.67139
R1838 VDD1.n4 VDD1.t5 1.67139
R1839 VDD1.n0 VDD1.t4 1.67139
R1840 VDD1.n0 VDD1.t6 1.67139
R1841 VDD1.n2 VDD1.t3 1.67139
R1842 VDD1.n2 VDD1.t2 1.67139
R1843 VDD1.n1 VDD1.t1 1.67139
R1844 VDD1.n1 VDD1.t7 1.67139
R1845 VDD1 VDD1.n5 1.05869
C0 VDD2 VN 8.343901f
C1 VDD2 VDD1 1.59913f
C2 VTAIL VN 8.63781f
C3 VTAIL VDD1 7.99977f
C4 VN VP 7.21721f
C5 VDD1 VP 8.67505f
C6 VTAIL VDD2 8.05191f
C7 VDD2 VP 0.483302f
C8 VTAIL VP 8.651919f
C9 VDD1 VN 0.150924f
C10 VDD2 B 5.00594f
C11 VDD1 B 5.407413f
C12 VTAIL B 10.152764f
C13 VN B 14.19514f
C14 VP B 12.747399f
C15 VDD1.t4 B 0.231672f
C16 VDD1.t6 B 0.231672f
C17 VDD1.n0 B 2.07312f
C18 VDD1.t1 B 0.231672f
C19 VDD1.t7 B 0.231672f
C20 VDD1.n1 B 2.07214f
C21 VDD1.t3 B 0.231672f
C22 VDD1.t2 B 0.231672f
C23 VDD1.n2 B 2.07214f
C24 VDD1.n3 B 3.09019f
C25 VDD1.t0 B 0.231672f
C26 VDD1.t5 B 0.231672f
C27 VDD1.n4 B 2.06434f
C28 VDD1.n5 B 2.82089f
C29 VP.n0 B 0.032543f
C30 VP.t5 B 1.80049f
C31 VP.n1 B 0.022648f
C32 VP.n2 B 0.024684f
C33 VP.t4 B 1.80049f
C34 VP.n3 B 0.049059f
C35 VP.n4 B 0.024684f
C36 VP.t0 B 1.80049f
C37 VP.n5 B 0.640244f
C38 VP.n6 B 0.024684f
C39 VP.n7 B 0.045774f
C40 VP.n8 B 0.032543f
C41 VP.t2 B 1.80049f
C42 VP.n9 B 0.022648f
C43 VP.n10 B 0.024684f
C44 VP.t7 B 1.80049f
C45 VP.n11 B 0.049059f
C46 VP.n12 B 0.024684f
C47 VP.t1 B 1.80049f
C48 VP.n13 B 0.706829f
C49 VP.t3 B 1.96492f
C50 VP.n14 B 0.693367f
C51 VP.n15 B 0.211449f
C52 VP.n16 B 0.036691f
C53 VP.n17 B 0.049059f
C54 VP.n18 B 0.019955f
C55 VP.n19 B 0.024684f
C56 VP.n20 B 0.024684f
C57 VP.n21 B 0.024684f
C58 VP.n22 B 0.036691f
C59 VP.n23 B 0.640244f
C60 VP.n24 B 0.032603f
C61 VP.n25 B 0.049651f
C62 VP.n26 B 0.024684f
C63 VP.n27 B 0.024684f
C64 VP.n28 B 0.024684f
C65 VP.n29 B 0.045774f
C66 VP.n30 B 0.04078f
C67 VP.n31 B 0.724138f
C68 VP.n32 B 1.33566f
C69 VP.n33 B 1.35367f
C70 VP.t6 B 1.80049f
C71 VP.n34 B 0.724138f
C72 VP.n35 B 0.04078f
C73 VP.n36 B 0.032543f
C74 VP.n37 B 0.024684f
C75 VP.n38 B 0.024684f
C76 VP.n39 B 0.022648f
C77 VP.n40 B 0.049651f
C78 VP.n41 B 0.032603f
C79 VP.n42 B 0.024684f
C80 VP.n43 B 0.024684f
C81 VP.n44 B 0.036691f
C82 VP.n45 B 0.049059f
C83 VP.n46 B 0.019955f
C84 VP.n47 B 0.024684f
C85 VP.n48 B 0.024684f
C86 VP.n49 B 0.024684f
C87 VP.n50 B 0.036691f
C88 VP.n51 B 0.640244f
C89 VP.n52 B 0.032603f
C90 VP.n53 B 0.049651f
C91 VP.n54 B 0.024684f
C92 VP.n55 B 0.024684f
C93 VP.n56 B 0.024684f
C94 VP.n57 B 0.045774f
C95 VP.n58 B 0.04078f
C96 VP.n59 B 0.724138f
C97 VP.n60 B 0.031777f
C98 VDD2.t0 B 0.228762f
C99 VDD2.t1 B 0.228762f
C100 VDD2.n0 B 2.04611f
C101 VDD2.t2 B 0.228762f
C102 VDD2.t5 B 0.228762f
C103 VDD2.n1 B 2.04611f
C104 VDD2.n2 B 3.00029f
C105 VDD2.t3 B 0.228762f
C106 VDD2.t7 B 0.228762f
C107 VDD2.n3 B 2.03841f
C108 VDD2.n4 B 2.75547f
C109 VDD2.t6 B 0.228762f
C110 VDD2.t4 B 0.228762f
C111 VDD2.n5 B 2.04607f
C112 VTAIL.t11 B 0.184129f
C113 VTAIL.t10 B 0.184129f
C114 VTAIL.n0 B 1.58483f
C115 VTAIL.n1 B 0.335644f
C116 VTAIL.t8 B 2.02174f
C117 VTAIL.n2 B 0.426989f
C118 VTAIL.t5 B 2.02174f
C119 VTAIL.n3 B 0.426989f
C120 VTAIL.t0 B 0.184129f
C121 VTAIL.t7 B 0.184129f
C122 VTAIL.n4 B 1.58483f
C123 VTAIL.n5 B 0.473422f
C124 VTAIL.t1 B 2.02174f
C125 VTAIL.n6 B 1.45303f
C126 VTAIL.t15 B 2.02174f
C127 VTAIL.n7 B 1.45302f
C128 VTAIL.t12 B 0.184129f
C129 VTAIL.t14 B 0.184129f
C130 VTAIL.n8 B 1.58484f
C131 VTAIL.n9 B 0.473417f
C132 VTAIL.t13 B 2.02174f
C133 VTAIL.n10 B 0.426984f
C134 VTAIL.t3 B 2.02174f
C135 VTAIL.n11 B 0.426984f
C136 VTAIL.t4 B 0.184129f
C137 VTAIL.t6 B 0.184129f
C138 VTAIL.n12 B 1.58484f
C139 VTAIL.n13 B 0.473417f
C140 VTAIL.t2 B 2.02174f
C141 VTAIL.n14 B 1.45303f
C142 VTAIL.t9 B 2.02174f
C143 VTAIL.n15 B 1.44934f
C144 VN.n0 B 0.031837f
C145 VN.t2 B 1.76141f
C146 VN.n1 B 0.022156f
C147 VN.n2 B 0.024148f
C148 VN.t5 B 1.76141f
C149 VN.n3 B 0.047994f
C150 VN.n4 B 0.024148f
C151 VN.t6 B 1.76141f
C152 VN.n5 B 0.691487f
C153 VN.t7 B 1.92227f
C154 VN.n6 B 0.678317f
C155 VN.n7 B 0.20686f
C156 VN.n8 B 0.035895f
C157 VN.n9 B 0.047994f
C158 VN.n10 B 0.019521f
C159 VN.n11 B 0.024148f
C160 VN.n12 B 0.024148f
C161 VN.n13 B 0.024148f
C162 VN.n14 B 0.035895f
C163 VN.n15 B 0.626347f
C164 VN.n16 B 0.031895f
C165 VN.n17 B 0.048573f
C166 VN.n18 B 0.024148f
C167 VN.n19 B 0.024148f
C168 VN.n20 B 0.024148f
C169 VN.n21 B 0.044781f
C170 VN.n22 B 0.039894f
C171 VN.n23 B 0.70842f
C172 VN.n24 B 0.031087f
C173 VN.n25 B 0.031837f
C174 VN.t4 B 1.76141f
C175 VN.n26 B 0.022156f
C176 VN.n27 B 0.024148f
C177 VN.t0 B 1.76141f
C178 VN.n28 B 0.047994f
C179 VN.n29 B 0.024148f
C180 VN.t1 B 1.76141f
C181 VN.n30 B 0.691487f
C182 VN.t3 B 1.92227f
C183 VN.n31 B 0.678317f
C184 VN.n32 B 0.20686f
C185 VN.n33 B 0.035895f
C186 VN.n34 B 0.047994f
C187 VN.n35 B 0.019521f
C188 VN.n36 B 0.024148f
C189 VN.n37 B 0.024148f
C190 VN.n38 B 0.024148f
C191 VN.n39 B 0.035895f
C192 VN.n40 B 0.626347f
C193 VN.n41 B 0.031895f
C194 VN.n42 B 0.048573f
C195 VN.n43 B 0.024148f
C196 VN.n44 B 0.024148f
C197 VN.n45 B 0.024148f
C198 VN.n46 B 0.044781f
C199 VN.n47 B 0.039894f
C200 VN.n48 B 0.70842f
C201 VN.n49 B 1.31967f
.ends

