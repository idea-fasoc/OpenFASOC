* NGSPICE file created from diff_pair_sample_0747.ext - technology: sky130A

.subckt diff_pair_sample_0747 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=0 ps=0 w=19.22 l=1.5
X1 B.t8 B.t6 B.t7 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=0 ps=0 w=19.22 l=1.5
X2 VTAIL.t11 VP.t0 VDD1.t3 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=3.1713 ps=19.55 w=19.22 l=1.5
X3 VTAIL.t3 VN.t0 VDD2.t5 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=3.1713 ps=19.55 w=19.22 l=1.5
X4 VDD1.t4 VP.t1 VTAIL.t10 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=3.1713 ps=19.55 w=19.22 l=1.5
X5 VDD2.t4 VN.t1 VTAIL.t2 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=7.4958 ps=39.22 w=19.22 l=1.5
X6 B.t5 B.t3 B.t4 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=0 ps=0 w=19.22 l=1.5
X7 B.t2 B.t0 B.t1 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=0 ps=0 w=19.22 l=1.5
X8 VTAIL.t9 VP.t2 VDD1.t5 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=3.1713 ps=19.55 w=19.22 l=1.5
X9 VTAIL.t4 VN.t2 VDD2.t3 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=3.1713 ps=19.55 w=19.22 l=1.5
X10 VDD1.t1 VP.t3 VTAIL.t8 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=7.4958 ps=39.22 w=19.22 l=1.5
X11 VDD2.t2 VN.t3 VTAIL.t5 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=7.4958 ps=39.22 w=19.22 l=1.5
X12 VDD2.t1 VN.t4 VTAIL.t1 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=3.1713 ps=19.55 w=19.22 l=1.5
X13 VDD1.t2 VP.t4 VTAIL.t7 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=3.1713 ps=19.55 w=19.22 l=1.5
X14 VDD1.t0 VP.t5 VTAIL.t6 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=3.1713 pd=19.55 as=7.4958 ps=39.22 w=19.22 l=1.5
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n2434_n4812# sky130_fd_pr__pfet_01v8 ad=7.4958 pd=39.22 as=3.1713 ps=19.55 w=19.22 l=1.5
R0 B.n450 B.n449 585
R1 B.n448 B.n119 585
R2 B.n447 B.n446 585
R3 B.n445 B.n120 585
R4 B.n444 B.n443 585
R5 B.n442 B.n121 585
R6 B.n441 B.n440 585
R7 B.n439 B.n122 585
R8 B.n438 B.n437 585
R9 B.n436 B.n123 585
R10 B.n435 B.n434 585
R11 B.n433 B.n124 585
R12 B.n432 B.n431 585
R13 B.n430 B.n125 585
R14 B.n429 B.n428 585
R15 B.n427 B.n126 585
R16 B.n426 B.n425 585
R17 B.n424 B.n127 585
R18 B.n423 B.n422 585
R19 B.n421 B.n128 585
R20 B.n420 B.n419 585
R21 B.n418 B.n129 585
R22 B.n417 B.n416 585
R23 B.n415 B.n130 585
R24 B.n414 B.n413 585
R25 B.n412 B.n131 585
R26 B.n411 B.n410 585
R27 B.n409 B.n132 585
R28 B.n408 B.n407 585
R29 B.n406 B.n133 585
R30 B.n405 B.n404 585
R31 B.n403 B.n134 585
R32 B.n402 B.n401 585
R33 B.n400 B.n135 585
R34 B.n399 B.n398 585
R35 B.n397 B.n136 585
R36 B.n396 B.n395 585
R37 B.n394 B.n137 585
R38 B.n393 B.n392 585
R39 B.n391 B.n138 585
R40 B.n390 B.n389 585
R41 B.n388 B.n139 585
R42 B.n387 B.n386 585
R43 B.n385 B.n140 585
R44 B.n384 B.n383 585
R45 B.n382 B.n141 585
R46 B.n381 B.n380 585
R47 B.n379 B.n142 585
R48 B.n378 B.n377 585
R49 B.n376 B.n143 585
R50 B.n375 B.n374 585
R51 B.n373 B.n144 585
R52 B.n372 B.n371 585
R53 B.n370 B.n145 585
R54 B.n369 B.n368 585
R55 B.n367 B.n146 585
R56 B.n366 B.n365 585
R57 B.n364 B.n147 585
R58 B.n363 B.n362 585
R59 B.n361 B.n148 585
R60 B.n360 B.n359 585
R61 B.n358 B.n149 585
R62 B.n357 B.n356 585
R63 B.n355 B.n354 585
R64 B.n353 B.n153 585
R65 B.n352 B.n351 585
R66 B.n350 B.n154 585
R67 B.n349 B.n348 585
R68 B.n347 B.n155 585
R69 B.n346 B.n345 585
R70 B.n344 B.n156 585
R71 B.n343 B.n342 585
R72 B.n340 B.n157 585
R73 B.n339 B.n338 585
R74 B.n337 B.n160 585
R75 B.n336 B.n335 585
R76 B.n334 B.n161 585
R77 B.n333 B.n332 585
R78 B.n331 B.n162 585
R79 B.n330 B.n329 585
R80 B.n328 B.n163 585
R81 B.n327 B.n326 585
R82 B.n325 B.n164 585
R83 B.n324 B.n323 585
R84 B.n322 B.n165 585
R85 B.n321 B.n320 585
R86 B.n319 B.n166 585
R87 B.n318 B.n317 585
R88 B.n316 B.n167 585
R89 B.n315 B.n314 585
R90 B.n313 B.n168 585
R91 B.n312 B.n311 585
R92 B.n310 B.n169 585
R93 B.n309 B.n308 585
R94 B.n307 B.n170 585
R95 B.n306 B.n305 585
R96 B.n304 B.n171 585
R97 B.n303 B.n302 585
R98 B.n301 B.n172 585
R99 B.n300 B.n299 585
R100 B.n298 B.n173 585
R101 B.n297 B.n296 585
R102 B.n295 B.n174 585
R103 B.n294 B.n293 585
R104 B.n292 B.n175 585
R105 B.n291 B.n290 585
R106 B.n289 B.n176 585
R107 B.n288 B.n287 585
R108 B.n286 B.n177 585
R109 B.n285 B.n284 585
R110 B.n283 B.n178 585
R111 B.n282 B.n281 585
R112 B.n280 B.n179 585
R113 B.n279 B.n278 585
R114 B.n277 B.n180 585
R115 B.n276 B.n275 585
R116 B.n274 B.n181 585
R117 B.n273 B.n272 585
R118 B.n271 B.n182 585
R119 B.n270 B.n269 585
R120 B.n268 B.n183 585
R121 B.n267 B.n266 585
R122 B.n265 B.n184 585
R123 B.n264 B.n263 585
R124 B.n262 B.n185 585
R125 B.n261 B.n260 585
R126 B.n259 B.n186 585
R127 B.n258 B.n257 585
R128 B.n256 B.n187 585
R129 B.n255 B.n254 585
R130 B.n253 B.n188 585
R131 B.n252 B.n251 585
R132 B.n250 B.n189 585
R133 B.n249 B.n248 585
R134 B.n247 B.n190 585
R135 B.n451 B.n118 585
R136 B.n453 B.n452 585
R137 B.n454 B.n117 585
R138 B.n456 B.n455 585
R139 B.n457 B.n116 585
R140 B.n459 B.n458 585
R141 B.n460 B.n115 585
R142 B.n462 B.n461 585
R143 B.n463 B.n114 585
R144 B.n465 B.n464 585
R145 B.n466 B.n113 585
R146 B.n468 B.n467 585
R147 B.n469 B.n112 585
R148 B.n471 B.n470 585
R149 B.n472 B.n111 585
R150 B.n474 B.n473 585
R151 B.n475 B.n110 585
R152 B.n477 B.n476 585
R153 B.n478 B.n109 585
R154 B.n480 B.n479 585
R155 B.n481 B.n108 585
R156 B.n483 B.n482 585
R157 B.n484 B.n107 585
R158 B.n486 B.n485 585
R159 B.n487 B.n106 585
R160 B.n489 B.n488 585
R161 B.n490 B.n105 585
R162 B.n492 B.n491 585
R163 B.n493 B.n104 585
R164 B.n495 B.n494 585
R165 B.n496 B.n103 585
R166 B.n498 B.n497 585
R167 B.n499 B.n102 585
R168 B.n501 B.n500 585
R169 B.n502 B.n101 585
R170 B.n504 B.n503 585
R171 B.n505 B.n100 585
R172 B.n507 B.n506 585
R173 B.n508 B.n99 585
R174 B.n510 B.n509 585
R175 B.n511 B.n98 585
R176 B.n513 B.n512 585
R177 B.n514 B.n97 585
R178 B.n516 B.n515 585
R179 B.n517 B.n96 585
R180 B.n519 B.n518 585
R181 B.n520 B.n95 585
R182 B.n522 B.n521 585
R183 B.n523 B.n94 585
R184 B.n525 B.n524 585
R185 B.n526 B.n93 585
R186 B.n528 B.n527 585
R187 B.n529 B.n92 585
R188 B.n531 B.n530 585
R189 B.n532 B.n91 585
R190 B.n534 B.n533 585
R191 B.n535 B.n90 585
R192 B.n537 B.n536 585
R193 B.n538 B.n89 585
R194 B.n540 B.n539 585
R195 B.n744 B.n743 585
R196 B.n742 B.n17 585
R197 B.n741 B.n740 585
R198 B.n739 B.n18 585
R199 B.n738 B.n737 585
R200 B.n736 B.n19 585
R201 B.n735 B.n734 585
R202 B.n733 B.n20 585
R203 B.n732 B.n731 585
R204 B.n730 B.n21 585
R205 B.n729 B.n728 585
R206 B.n727 B.n22 585
R207 B.n726 B.n725 585
R208 B.n724 B.n23 585
R209 B.n723 B.n722 585
R210 B.n721 B.n24 585
R211 B.n720 B.n719 585
R212 B.n718 B.n25 585
R213 B.n717 B.n716 585
R214 B.n715 B.n26 585
R215 B.n714 B.n713 585
R216 B.n712 B.n27 585
R217 B.n711 B.n710 585
R218 B.n709 B.n28 585
R219 B.n708 B.n707 585
R220 B.n706 B.n29 585
R221 B.n705 B.n704 585
R222 B.n703 B.n30 585
R223 B.n702 B.n701 585
R224 B.n700 B.n31 585
R225 B.n699 B.n698 585
R226 B.n697 B.n32 585
R227 B.n696 B.n695 585
R228 B.n694 B.n33 585
R229 B.n693 B.n692 585
R230 B.n691 B.n34 585
R231 B.n690 B.n689 585
R232 B.n688 B.n35 585
R233 B.n687 B.n686 585
R234 B.n685 B.n36 585
R235 B.n684 B.n683 585
R236 B.n682 B.n37 585
R237 B.n681 B.n680 585
R238 B.n679 B.n38 585
R239 B.n678 B.n677 585
R240 B.n676 B.n39 585
R241 B.n675 B.n674 585
R242 B.n673 B.n40 585
R243 B.n672 B.n671 585
R244 B.n670 B.n41 585
R245 B.n669 B.n668 585
R246 B.n667 B.n42 585
R247 B.n666 B.n665 585
R248 B.n664 B.n43 585
R249 B.n663 B.n662 585
R250 B.n661 B.n44 585
R251 B.n660 B.n659 585
R252 B.n658 B.n45 585
R253 B.n657 B.n656 585
R254 B.n655 B.n46 585
R255 B.n654 B.n653 585
R256 B.n652 B.n47 585
R257 B.n651 B.n650 585
R258 B.n649 B.n648 585
R259 B.n647 B.n51 585
R260 B.n646 B.n645 585
R261 B.n644 B.n52 585
R262 B.n643 B.n642 585
R263 B.n641 B.n53 585
R264 B.n640 B.n639 585
R265 B.n638 B.n54 585
R266 B.n637 B.n636 585
R267 B.n634 B.n55 585
R268 B.n633 B.n632 585
R269 B.n631 B.n58 585
R270 B.n630 B.n629 585
R271 B.n628 B.n59 585
R272 B.n627 B.n626 585
R273 B.n625 B.n60 585
R274 B.n624 B.n623 585
R275 B.n622 B.n61 585
R276 B.n621 B.n620 585
R277 B.n619 B.n62 585
R278 B.n618 B.n617 585
R279 B.n616 B.n63 585
R280 B.n615 B.n614 585
R281 B.n613 B.n64 585
R282 B.n612 B.n611 585
R283 B.n610 B.n65 585
R284 B.n609 B.n608 585
R285 B.n607 B.n66 585
R286 B.n606 B.n605 585
R287 B.n604 B.n67 585
R288 B.n603 B.n602 585
R289 B.n601 B.n68 585
R290 B.n600 B.n599 585
R291 B.n598 B.n69 585
R292 B.n597 B.n596 585
R293 B.n595 B.n70 585
R294 B.n594 B.n593 585
R295 B.n592 B.n71 585
R296 B.n591 B.n590 585
R297 B.n589 B.n72 585
R298 B.n588 B.n587 585
R299 B.n586 B.n73 585
R300 B.n585 B.n584 585
R301 B.n583 B.n74 585
R302 B.n582 B.n581 585
R303 B.n580 B.n75 585
R304 B.n579 B.n578 585
R305 B.n577 B.n76 585
R306 B.n576 B.n575 585
R307 B.n574 B.n77 585
R308 B.n573 B.n572 585
R309 B.n571 B.n78 585
R310 B.n570 B.n569 585
R311 B.n568 B.n79 585
R312 B.n567 B.n566 585
R313 B.n565 B.n80 585
R314 B.n564 B.n563 585
R315 B.n562 B.n81 585
R316 B.n561 B.n560 585
R317 B.n559 B.n82 585
R318 B.n558 B.n557 585
R319 B.n556 B.n83 585
R320 B.n555 B.n554 585
R321 B.n553 B.n84 585
R322 B.n552 B.n551 585
R323 B.n550 B.n85 585
R324 B.n549 B.n548 585
R325 B.n547 B.n86 585
R326 B.n546 B.n545 585
R327 B.n544 B.n87 585
R328 B.n543 B.n542 585
R329 B.n541 B.n88 585
R330 B.n745 B.n16 585
R331 B.n747 B.n746 585
R332 B.n748 B.n15 585
R333 B.n750 B.n749 585
R334 B.n751 B.n14 585
R335 B.n753 B.n752 585
R336 B.n754 B.n13 585
R337 B.n756 B.n755 585
R338 B.n757 B.n12 585
R339 B.n759 B.n758 585
R340 B.n760 B.n11 585
R341 B.n762 B.n761 585
R342 B.n763 B.n10 585
R343 B.n765 B.n764 585
R344 B.n766 B.n9 585
R345 B.n768 B.n767 585
R346 B.n769 B.n8 585
R347 B.n771 B.n770 585
R348 B.n772 B.n7 585
R349 B.n774 B.n773 585
R350 B.n775 B.n6 585
R351 B.n777 B.n776 585
R352 B.n778 B.n5 585
R353 B.n780 B.n779 585
R354 B.n781 B.n4 585
R355 B.n783 B.n782 585
R356 B.n784 B.n3 585
R357 B.n786 B.n785 585
R358 B.n787 B.n0 585
R359 B.n2 B.n1 585
R360 B.n205 B.n204 585
R361 B.n207 B.n206 585
R362 B.n208 B.n203 585
R363 B.n210 B.n209 585
R364 B.n211 B.n202 585
R365 B.n213 B.n212 585
R366 B.n214 B.n201 585
R367 B.n216 B.n215 585
R368 B.n217 B.n200 585
R369 B.n219 B.n218 585
R370 B.n220 B.n199 585
R371 B.n222 B.n221 585
R372 B.n223 B.n198 585
R373 B.n225 B.n224 585
R374 B.n226 B.n197 585
R375 B.n228 B.n227 585
R376 B.n229 B.n196 585
R377 B.n231 B.n230 585
R378 B.n232 B.n195 585
R379 B.n234 B.n233 585
R380 B.n235 B.n194 585
R381 B.n237 B.n236 585
R382 B.n238 B.n193 585
R383 B.n240 B.n239 585
R384 B.n241 B.n192 585
R385 B.n243 B.n242 585
R386 B.n244 B.n191 585
R387 B.n246 B.n245 585
R388 B.n247 B.n246 545.355
R389 B.n451 B.n450 545.355
R390 B.n541 B.n540 545.355
R391 B.n745 B.n744 545.355
R392 B.n158 B.t6 514.241
R393 B.n150 B.t3 514.241
R394 B.n56 B.t9 514.241
R395 B.n48 B.t0 514.241
R396 B.n789 B.n788 256.663
R397 B.n788 B.n787 235.042
R398 B.n788 B.n2 235.042
R399 B.n248 B.n247 163.367
R400 B.n248 B.n189 163.367
R401 B.n252 B.n189 163.367
R402 B.n253 B.n252 163.367
R403 B.n254 B.n253 163.367
R404 B.n254 B.n187 163.367
R405 B.n258 B.n187 163.367
R406 B.n259 B.n258 163.367
R407 B.n260 B.n259 163.367
R408 B.n260 B.n185 163.367
R409 B.n264 B.n185 163.367
R410 B.n265 B.n264 163.367
R411 B.n266 B.n265 163.367
R412 B.n266 B.n183 163.367
R413 B.n270 B.n183 163.367
R414 B.n271 B.n270 163.367
R415 B.n272 B.n271 163.367
R416 B.n272 B.n181 163.367
R417 B.n276 B.n181 163.367
R418 B.n277 B.n276 163.367
R419 B.n278 B.n277 163.367
R420 B.n278 B.n179 163.367
R421 B.n282 B.n179 163.367
R422 B.n283 B.n282 163.367
R423 B.n284 B.n283 163.367
R424 B.n284 B.n177 163.367
R425 B.n288 B.n177 163.367
R426 B.n289 B.n288 163.367
R427 B.n290 B.n289 163.367
R428 B.n290 B.n175 163.367
R429 B.n294 B.n175 163.367
R430 B.n295 B.n294 163.367
R431 B.n296 B.n295 163.367
R432 B.n296 B.n173 163.367
R433 B.n300 B.n173 163.367
R434 B.n301 B.n300 163.367
R435 B.n302 B.n301 163.367
R436 B.n302 B.n171 163.367
R437 B.n306 B.n171 163.367
R438 B.n307 B.n306 163.367
R439 B.n308 B.n307 163.367
R440 B.n308 B.n169 163.367
R441 B.n312 B.n169 163.367
R442 B.n313 B.n312 163.367
R443 B.n314 B.n313 163.367
R444 B.n314 B.n167 163.367
R445 B.n318 B.n167 163.367
R446 B.n319 B.n318 163.367
R447 B.n320 B.n319 163.367
R448 B.n320 B.n165 163.367
R449 B.n324 B.n165 163.367
R450 B.n325 B.n324 163.367
R451 B.n326 B.n325 163.367
R452 B.n326 B.n163 163.367
R453 B.n330 B.n163 163.367
R454 B.n331 B.n330 163.367
R455 B.n332 B.n331 163.367
R456 B.n332 B.n161 163.367
R457 B.n336 B.n161 163.367
R458 B.n337 B.n336 163.367
R459 B.n338 B.n337 163.367
R460 B.n338 B.n157 163.367
R461 B.n343 B.n157 163.367
R462 B.n344 B.n343 163.367
R463 B.n345 B.n344 163.367
R464 B.n345 B.n155 163.367
R465 B.n349 B.n155 163.367
R466 B.n350 B.n349 163.367
R467 B.n351 B.n350 163.367
R468 B.n351 B.n153 163.367
R469 B.n355 B.n153 163.367
R470 B.n356 B.n355 163.367
R471 B.n356 B.n149 163.367
R472 B.n360 B.n149 163.367
R473 B.n361 B.n360 163.367
R474 B.n362 B.n361 163.367
R475 B.n362 B.n147 163.367
R476 B.n366 B.n147 163.367
R477 B.n367 B.n366 163.367
R478 B.n368 B.n367 163.367
R479 B.n368 B.n145 163.367
R480 B.n372 B.n145 163.367
R481 B.n373 B.n372 163.367
R482 B.n374 B.n373 163.367
R483 B.n374 B.n143 163.367
R484 B.n378 B.n143 163.367
R485 B.n379 B.n378 163.367
R486 B.n380 B.n379 163.367
R487 B.n380 B.n141 163.367
R488 B.n384 B.n141 163.367
R489 B.n385 B.n384 163.367
R490 B.n386 B.n385 163.367
R491 B.n386 B.n139 163.367
R492 B.n390 B.n139 163.367
R493 B.n391 B.n390 163.367
R494 B.n392 B.n391 163.367
R495 B.n392 B.n137 163.367
R496 B.n396 B.n137 163.367
R497 B.n397 B.n396 163.367
R498 B.n398 B.n397 163.367
R499 B.n398 B.n135 163.367
R500 B.n402 B.n135 163.367
R501 B.n403 B.n402 163.367
R502 B.n404 B.n403 163.367
R503 B.n404 B.n133 163.367
R504 B.n408 B.n133 163.367
R505 B.n409 B.n408 163.367
R506 B.n410 B.n409 163.367
R507 B.n410 B.n131 163.367
R508 B.n414 B.n131 163.367
R509 B.n415 B.n414 163.367
R510 B.n416 B.n415 163.367
R511 B.n416 B.n129 163.367
R512 B.n420 B.n129 163.367
R513 B.n421 B.n420 163.367
R514 B.n422 B.n421 163.367
R515 B.n422 B.n127 163.367
R516 B.n426 B.n127 163.367
R517 B.n427 B.n426 163.367
R518 B.n428 B.n427 163.367
R519 B.n428 B.n125 163.367
R520 B.n432 B.n125 163.367
R521 B.n433 B.n432 163.367
R522 B.n434 B.n433 163.367
R523 B.n434 B.n123 163.367
R524 B.n438 B.n123 163.367
R525 B.n439 B.n438 163.367
R526 B.n440 B.n439 163.367
R527 B.n440 B.n121 163.367
R528 B.n444 B.n121 163.367
R529 B.n445 B.n444 163.367
R530 B.n446 B.n445 163.367
R531 B.n446 B.n119 163.367
R532 B.n450 B.n119 163.367
R533 B.n540 B.n89 163.367
R534 B.n536 B.n89 163.367
R535 B.n536 B.n535 163.367
R536 B.n535 B.n534 163.367
R537 B.n534 B.n91 163.367
R538 B.n530 B.n91 163.367
R539 B.n530 B.n529 163.367
R540 B.n529 B.n528 163.367
R541 B.n528 B.n93 163.367
R542 B.n524 B.n93 163.367
R543 B.n524 B.n523 163.367
R544 B.n523 B.n522 163.367
R545 B.n522 B.n95 163.367
R546 B.n518 B.n95 163.367
R547 B.n518 B.n517 163.367
R548 B.n517 B.n516 163.367
R549 B.n516 B.n97 163.367
R550 B.n512 B.n97 163.367
R551 B.n512 B.n511 163.367
R552 B.n511 B.n510 163.367
R553 B.n510 B.n99 163.367
R554 B.n506 B.n99 163.367
R555 B.n506 B.n505 163.367
R556 B.n505 B.n504 163.367
R557 B.n504 B.n101 163.367
R558 B.n500 B.n101 163.367
R559 B.n500 B.n499 163.367
R560 B.n499 B.n498 163.367
R561 B.n498 B.n103 163.367
R562 B.n494 B.n103 163.367
R563 B.n494 B.n493 163.367
R564 B.n493 B.n492 163.367
R565 B.n492 B.n105 163.367
R566 B.n488 B.n105 163.367
R567 B.n488 B.n487 163.367
R568 B.n487 B.n486 163.367
R569 B.n486 B.n107 163.367
R570 B.n482 B.n107 163.367
R571 B.n482 B.n481 163.367
R572 B.n481 B.n480 163.367
R573 B.n480 B.n109 163.367
R574 B.n476 B.n109 163.367
R575 B.n476 B.n475 163.367
R576 B.n475 B.n474 163.367
R577 B.n474 B.n111 163.367
R578 B.n470 B.n111 163.367
R579 B.n470 B.n469 163.367
R580 B.n469 B.n468 163.367
R581 B.n468 B.n113 163.367
R582 B.n464 B.n113 163.367
R583 B.n464 B.n463 163.367
R584 B.n463 B.n462 163.367
R585 B.n462 B.n115 163.367
R586 B.n458 B.n115 163.367
R587 B.n458 B.n457 163.367
R588 B.n457 B.n456 163.367
R589 B.n456 B.n117 163.367
R590 B.n452 B.n117 163.367
R591 B.n452 B.n451 163.367
R592 B.n744 B.n17 163.367
R593 B.n740 B.n17 163.367
R594 B.n740 B.n739 163.367
R595 B.n739 B.n738 163.367
R596 B.n738 B.n19 163.367
R597 B.n734 B.n19 163.367
R598 B.n734 B.n733 163.367
R599 B.n733 B.n732 163.367
R600 B.n732 B.n21 163.367
R601 B.n728 B.n21 163.367
R602 B.n728 B.n727 163.367
R603 B.n727 B.n726 163.367
R604 B.n726 B.n23 163.367
R605 B.n722 B.n23 163.367
R606 B.n722 B.n721 163.367
R607 B.n721 B.n720 163.367
R608 B.n720 B.n25 163.367
R609 B.n716 B.n25 163.367
R610 B.n716 B.n715 163.367
R611 B.n715 B.n714 163.367
R612 B.n714 B.n27 163.367
R613 B.n710 B.n27 163.367
R614 B.n710 B.n709 163.367
R615 B.n709 B.n708 163.367
R616 B.n708 B.n29 163.367
R617 B.n704 B.n29 163.367
R618 B.n704 B.n703 163.367
R619 B.n703 B.n702 163.367
R620 B.n702 B.n31 163.367
R621 B.n698 B.n31 163.367
R622 B.n698 B.n697 163.367
R623 B.n697 B.n696 163.367
R624 B.n696 B.n33 163.367
R625 B.n692 B.n33 163.367
R626 B.n692 B.n691 163.367
R627 B.n691 B.n690 163.367
R628 B.n690 B.n35 163.367
R629 B.n686 B.n35 163.367
R630 B.n686 B.n685 163.367
R631 B.n685 B.n684 163.367
R632 B.n684 B.n37 163.367
R633 B.n680 B.n37 163.367
R634 B.n680 B.n679 163.367
R635 B.n679 B.n678 163.367
R636 B.n678 B.n39 163.367
R637 B.n674 B.n39 163.367
R638 B.n674 B.n673 163.367
R639 B.n673 B.n672 163.367
R640 B.n672 B.n41 163.367
R641 B.n668 B.n41 163.367
R642 B.n668 B.n667 163.367
R643 B.n667 B.n666 163.367
R644 B.n666 B.n43 163.367
R645 B.n662 B.n43 163.367
R646 B.n662 B.n661 163.367
R647 B.n661 B.n660 163.367
R648 B.n660 B.n45 163.367
R649 B.n656 B.n45 163.367
R650 B.n656 B.n655 163.367
R651 B.n655 B.n654 163.367
R652 B.n654 B.n47 163.367
R653 B.n650 B.n47 163.367
R654 B.n650 B.n649 163.367
R655 B.n649 B.n51 163.367
R656 B.n645 B.n51 163.367
R657 B.n645 B.n644 163.367
R658 B.n644 B.n643 163.367
R659 B.n643 B.n53 163.367
R660 B.n639 B.n53 163.367
R661 B.n639 B.n638 163.367
R662 B.n638 B.n637 163.367
R663 B.n637 B.n55 163.367
R664 B.n632 B.n55 163.367
R665 B.n632 B.n631 163.367
R666 B.n631 B.n630 163.367
R667 B.n630 B.n59 163.367
R668 B.n626 B.n59 163.367
R669 B.n626 B.n625 163.367
R670 B.n625 B.n624 163.367
R671 B.n624 B.n61 163.367
R672 B.n620 B.n61 163.367
R673 B.n620 B.n619 163.367
R674 B.n619 B.n618 163.367
R675 B.n618 B.n63 163.367
R676 B.n614 B.n63 163.367
R677 B.n614 B.n613 163.367
R678 B.n613 B.n612 163.367
R679 B.n612 B.n65 163.367
R680 B.n608 B.n65 163.367
R681 B.n608 B.n607 163.367
R682 B.n607 B.n606 163.367
R683 B.n606 B.n67 163.367
R684 B.n602 B.n67 163.367
R685 B.n602 B.n601 163.367
R686 B.n601 B.n600 163.367
R687 B.n600 B.n69 163.367
R688 B.n596 B.n69 163.367
R689 B.n596 B.n595 163.367
R690 B.n595 B.n594 163.367
R691 B.n594 B.n71 163.367
R692 B.n590 B.n71 163.367
R693 B.n590 B.n589 163.367
R694 B.n589 B.n588 163.367
R695 B.n588 B.n73 163.367
R696 B.n584 B.n73 163.367
R697 B.n584 B.n583 163.367
R698 B.n583 B.n582 163.367
R699 B.n582 B.n75 163.367
R700 B.n578 B.n75 163.367
R701 B.n578 B.n577 163.367
R702 B.n577 B.n576 163.367
R703 B.n576 B.n77 163.367
R704 B.n572 B.n77 163.367
R705 B.n572 B.n571 163.367
R706 B.n571 B.n570 163.367
R707 B.n570 B.n79 163.367
R708 B.n566 B.n79 163.367
R709 B.n566 B.n565 163.367
R710 B.n565 B.n564 163.367
R711 B.n564 B.n81 163.367
R712 B.n560 B.n81 163.367
R713 B.n560 B.n559 163.367
R714 B.n559 B.n558 163.367
R715 B.n558 B.n83 163.367
R716 B.n554 B.n83 163.367
R717 B.n554 B.n553 163.367
R718 B.n553 B.n552 163.367
R719 B.n552 B.n85 163.367
R720 B.n548 B.n85 163.367
R721 B.n548 B.n547 163.367
R722 B.n547 B.n546 163.367
R723 B.n546 B.n87 163.367
R724 B.n542 B.n87 163.367
R725 B.n542 B.n541 163.367
R726 B.n746 B.n745 163.367
R727 B.n746 B.n15 163.367
R728 B.n750 B.n15 163.367
R729 B.n751 B.n750 163.367
R730 B.n752 B.n751 163.367
R731 B.n752 B.n13 163.367
R732 B.n756 B.n13 163.367
R733 B.n757 B.n756 163.367
R734 B.n758 B.n757 163.367
R735 B.n758 B.n11 163.367
R736 B.n762 B.n11 163.367
R737 B.n763 B.n762 163.367
R738 B.n764 B.n763 163.367
R739 B.n764 B.n9 163.367
R740 B.n768 B.n9 163.367
R741 B.n769 B.n768 163.367
R742 B.n770 B.n769 163.367
R743 B.n770 B.n7 163.367
R744 B.n774 B.n7 163.367
R745 B.n775 B.n774 163.367
R746 B.n776 B.n775 163.367
R747 B.n776 B.n5 163.367
R748 B.n780 B.n5 163.367
R749 B.n781 B.n780 163.367
R750 B.n782 B.n781 163.367
R751 B.n782 B.n3 163.367
R752 B.n786 B.n3 163.367
R753 B.n787 B.n786 163.367
R754 B.n205 B.n2 163.367
R755 B.n206 B.n205 163.367
R756 B.n206 B.n203 163.367
R757 B.n210 B.n203 163.367
R758 B.n211 B.n210 163.367
R759 B.n212 B.n211 163.367
R760 B.n212 B.n201 163.367
R761 B.n216 B.n201 163.367
R762 B.n217 B.n216 163.367
R763 B.n218 B.n217 163.367
R764 B.n218 B.n199 163.367
R765 B.n222 B.n199 163.367
R766 B.n223 B.n222 163.367
R767 B.n224 B.n223 163.367
R768 B.n224 B.n197 163.367
R769 B.n228 B.n197 163.367
R770 B.n229 B.n228 163.367
R771 B.n230 B.n229 163.367
R772 B.n230 B.n195 163.367
R773 B.n234 B.n195 163.367
R774 B.n235 B.n234 163.367
R775 B.n236 B.n235 163.367
R776 B.n236 B.n193 163.367
R777 B.n240 B.n193 163.367
R778 B.n241 B.n240 163.367
R779 B.n242 B.n241 163.367
R780 B.n242 B.n191 163.367
R781 B.n246 B.n191 163.367
R782 B.n150 B.t4 145.072
R783 B.n56 B.t11 145.072
R784 B.n158 B.t7 145.048
R785 B.n48 B.t2 145.048
R786 B.n151 B.t5 109.582
R787 B.n57 B.t10 109.582
R788 B.n159 B.t8 109.558
R789 B.n49 B.t1 109.558
R790 B.n341 B.n159 59.5399
R791 B.n152 B.n151 59.5399
R792 B.n635 B.n57 59.5399
R793 B.n50 B.n49 59.5399
R794 B.n159 B.n158 35.4914
R795 B.n151 B.n150 35.4914
R796 B.n57 B.n56 35.4914
R797 B.n49 B.n48 35.4914
R798 B.n743 B.n16 35.4346
R799 B.n539 B.n88 35.4346
R800 B.n245 B.n190 35.4346
R801 B.n449 B.n118 35.4346
R802 B B.n789 18.0485
R803 B.n747 B.n16 10.6151
R804 B.n748 B.n747 10.6151
R805 B.n749 B.n748 10.6151
R806 B.n749 B.n14 10.6151
R807 B.n753 B.n14 10.6151
R808 B.n754 B.n753 10.6151
R809 B.n755 B.n754 10.6151
R810 B.n755 B.n12 10.6151
R811 B.n759 B.n12 10.6151
R812 B.n760 B.n759 10.6151
R813 B.n761 B.n760 10.6151
R814 B.n761 B.n10 10.6151
R815 B.n765 B.n10 10.6151
R816 B.n766 B.n765 10.6151
R817 B.n767 B.n766 10.6151
R818 B.n767 B.n8 10.6151
R819 B.n771 B.n8 10.6151
R820 B.n772 B.n771 10.6151
R821 B.n773 B.n772 10.6151
R822 B.n773 B.n6 10.6151
R823 B.n777 B.n6 10.6151
R824 B.n778 B.n777 10.6151
R825 B.n779 B.n778 10.6151
R826 B.n779 B.n4 10.6151
R827 B.n783 B.n4 10.6151
R828 B.n784 B.n783 10.6151
R829 B.n785 B.n784 10.6151
R830 B.n785 B.n0 10.6151
R831 B.n743 B.n742 10.6151
R832 B.n742 B.n741 10.6151
R833 B.n741 B.n18 10.6151
R834 B.n737 B.n18 10.6151
R835 B.n737 B.n736 10.6151
R836 B.n736 B.n735 10.6151
R837 B.n735 B.n20 10.6151
R838 B.n731 B.n20 10.6151
R839 B.n731 B.n730 10.6151
R840 B.n730 B.n729 10.6151
R841 B.n729 B.n22 10.6151
R842 B.n725 B.n22 10.6151
R843 B.n725 B.n724 10.6151
R844 B.n724 B.n723 10.6151
R845 B.n723 B.n24 10.6151
R846 B.n719 B.n24 10.6151
R847 B.n719 B.n718 10.6151
R848 B.n718 B.n717 10.6151
R849 B.n717 B.n26 10.6151
R850 B.n713 B.n26 10.6151
R851 B.n713 B.n712 10.6151
R852 B.n712 B.n711 10.6151
R853 B.n711 B.n28 10.6151
R854 B.n707 B.n28 10.6151
R855 B.n707 B.n706 10.6151
R856 B.n706 B.n705 10.6151
R857 B.n705 B.n30 10.6151
R858 B.n701 B.n30 10.6151
R859 B.n701 B.n700 10.6151
R860 B.n700 B.n699 10.6151
R861 B.n699 B.n32 10.6151
R862 B.n695 B.n32 10.6151
R863 B.n695 B.n694 10.6151
R864 B.n694 B.n693 10.6151
R865 B.n693 B.n34 10.6151
R866 B.n689 B.n34 10.6151
R867 B.n689 B.n688 10.6151
R868 B.n688 B.n687 10.6151
R869 B.n687 B.n36 10.6151
R870 B.n683 B.n36 10.6151
R871 B.n683 B.n682 10.6151
R872 B.n682 B.n681 10.6151
R873 B.n681 B.n38 10.6151
R874 B.n677 B.n38 10.6151
R875 B.n677 B.n676 10.6151
R876 B.n676 B.n675 10.6151
R877 B.n675 B.n40 10.6151
R878 B.n671 B.n40 10.6151
R879 B.n671 B.n670 10.6151
R880 B.n670 B.n669 10.6151
R881 B.n669 B.n42 10.6151
R882 B.n665 B.n42 10.6151
R883 B.n665 B.n664 10.6151
R884 B.n664 B.n663 10.6151
R885 B.n663 B.n44 10.6151
R886 B.n659 B.n44 10.6151
R887 B.n659 B.n658 10.6151
R888 B.n658 B.n657 10.6151
R889 B.n657 B.n46 10.6151
R890 B.n653 B.n46 10.6151
R891 B.n653 B.n652 10.6151
R892 B.n652 B.n651 10.6151
R893 B.n648 B.n647 10.6151
R894 B.n647 B.n646 10.6151
R895 B.n646 B.n52 10.6151
R896 B.n642 B.n52 10.6151
R897 B.n642 B.n641 10.6151
R898 B.n641 B.n640 10.6151
R899 B.n640 B.n54 10.6151
R900 B.n636 B.n54 10.6151
R901 B.n634 B.n633 10.6151
R902 B.n633 B.n58 10.6151
R903 B.n629 B.n58 10.6151
R904 B.n629 B.n628 10.6151
R905 B.n628 B.n627 10.6151
R906 B.n627 B.n60 10.6151
R907 B.n623 B.n60 10.6151
R908 B.n623 B.n622 10.6151
R909 B.n622 B.n621 10.6151
R910 B.n621 B.n62 10.6151
R911 B.n617 B.n62 10.6151
R912 B.n617 B.n616 10.6151
R913 B.n616 B.n615 10.6151
R914 B.n615 B.n64 10.6151
R915 B.n611 B.n64 10.6151
R916 B.n611 B.n610 10.6151
R917 B.n610 B.n609 10.6151
R918 B.n609 B.n66 10.6151
R919 B.n605 B.n66 10.6151
R920 B.n605 B.n604 10.6151
R921 B.n604 B.n603 10.6151
R922 B.n603 B.n68 10.6151
R923 B.n599 B.n68 10.6151
R924 B.n599 B.n598 10.6151
R925 B.n598 B.n597 10.6151
R926 B.n597 B.n70 10.6151
R927 B.n593 B.n70 10.6151
R928 B.n593 B.n592 10.6151
R929 B.n592 B.n591 10.6151
R930 B.n591 B.n72 10.6151
R931 B.n587 B.n72 10.6151
R932 B.n587 B.n586 10.6151
R933 B.n586 B.n585 10.6151
R934 B.n585 B.n74 10.6151
R935 B.n581 B.n74 10.6151
R936 B.n581 B.n580 10.6151
R937 B.n580 B.n579 10.6151
R938 B.n579 B.n76 10.6151
R939 B.n575 B.n76 10.6151
R940 B.n575 B.n574 10.6151
R941 B.n574 B.n573 10.6151
R942 B.n573 B.n78 10.6151
R943 B.n569 B.n78 10.6151
R944 B.n569 B.n568 10.6151
R945 B.n568 B.n567 10.6151
R946 B.n567 B.n80 10.6151
R947 B.n563 B.n80 10.6151
R948 B.n563 B.n562 10.6151
R949 B.n562 B.n561 10.6151
R950 B.n561 B.n82 10.6151
R951 B.n557 B.n82 10.6151
R952 B.n557 B.n556 10.6151
R953 B.n556 B.n555 10.6151
R954 B.n555 B.n84 10.6151
R955 B.n551 B.n84 10.6151
R956 B.n551 B.n550 10.6151
R957 B.n550 B.n549 10.6151
R958 B.n549 B.n86 10.6151
R959 B.n545 B.n86 10.6151
R960 B.n545 B.n544 10.6151
R961 B.n544 B.n543 10.6151
R962 B.n543 B.n88 10.6151
R963 B.n539 B.n538 10.6151
R964 B.n538 B.n537 10.6151
R965 B.n537 B.n90 10.6151
R966 B.n533 B.n90 10.6151
R967 B.n533 B.n532 10.6151
R968 B.n532 B.n531 10.6151
R969 B.n531 B.n92 10.6151
R970 B.n527 B.n92 10.6151
R971 B.n527 B.n526 10.6151
R972 B.n526 B.n525 10.6151
R973 B.n525 B.n94 10.6151
R974 B.n521 B.n94 10.6151
R975 B.n521 B.n520 10.6151
R976 B.n520 B.n519 10.6151
R977 B.n519 B.n96 10.6151
R978 B.n515 B.n96 10.6151
R979 B.n515 B.n514 10.6151
R980 B.n514 B.n513 10.6151
R981 B.n513 B.n98 10.6151
R982 B.n509 B.n98 10.6151
R983 B.n509 B.n508 10.6151
R984 B.n508 B.n507 10.6151
R985 B.n507 B.n100 10.6151
R986 B.n503 B.n100 10.6151
R987 B.n503 B.n502 10.6151
R988 B.n502 B.n501 10.6151
R989 B.n501 B.n102 10.6151
R990 B.n497 B.n102 10.6151
R991 B.n497 B.n496 10.6151
R992 B.n496 B.n495 10.6151
R993 B.n495 B.n104 10.6151
R994 B.n491 B.n104 10.6151
R995 B.n491 B.n490 10.6151
R996 B.n490 B.n489 10.6151
R997 B.n489 B.n106 10.6151
R998 B.n485 B.n106 10.6151
R999 B.n485 B.n484 10.6151
R1000 B.n484 B.n483 10.6151
R1001 B.n483 B.n108 10.6151
R1002 B.n479 B.n108 10.6151
R1003 B.n479 B.n478 10.6151
R1004 B.n478 B.n477 10.6151
R1005 B.n477 B.n110 10.6151
R1006 B.n473 B.n110 10.6151
R1007 B.n473 B.n472 10.6151
R1008 B.n472 B.n471 10.6151
R1009 B.n471 B.n112 10.6151
R1010 B.n467 B.n112 10.6151
R1011 B.n467 B.n466 10.6151
R1012 B.n466 B.n465 10.6151
R1013 B.n465 B.n114 10.6151
R1014 B.n461 B.n114 10.6151
R1015 B.n461 B.n460 10.6151
R1016 B.n460 B.n459 10.6151
R1017 B.n459 B.n116 10.6151
R1018 B.n455 B.n116 10.6151
R1019 B.n455 B.n454 10.6151
R1020 B.n454 B.n453 10.6151
R1021 B.n453 B.n118 10.6151
R1022 B.n204 B.n1 10.6151
R1023 B.n207 B.n204 10.6151
R1024 B.n208 B.n207 10.6151
R1025 B.n209 B.n208 10.6151
R1026 B.n209 B.n202 10.6151
R1027 B.n213 B.n202 10.6151
R1028 B.n214 B.n213 10.6151
R1029 B.n215 B.n214 10.6151
R1030 B.n215 B.n200 10.6151
R1031 B.n219 B.n200 10.6151
R1032 B.n220 B.n219 10.6151
R1033 B.n221 B.n220 10.6151
R1034 B.n221 B.n198 10.6151
R1035 B.n225 B.n198 10.6151
R1036 B.n226 B.n225 10.6151
R1037 B.n227 B.n226 10.6151
R1038 B.n227 B.n196 10.6151
R1039 B.n231 B.n196 10.6151
R1040 B.n232 B.n231 10.6151
R1041 B.n233 B.n232 10.6151
R1042 B.n233 B.n194 10.6151
R1043 B.n237 B.n194 10.6151
R1044 B.n238 B.n237 10.6151
R1045 B.n239 B.n238 10.6151
R1046 B.n239 B.n192 10.6151
R1047 B.n243 B.n192 10.6151
R1048 B.n244 B.n243 10.6151
R1049 B.n245 B.n244 10.6151
R1050 B.n249 B.n190 10.6151
R1051 B.n250 B.n249 10.6151
R1052 B.n251 B.n250 10.6151
R1053 B.n251 B.n188 10.6151
R1054 B.n255 B.n188 10.6151
R1055 B.n256 B.n255 10.6151
R1056 B.n257 B.n256 10.6151
R1057 B.n257 B.n186 10.6151
R1058 B.n261 B.n186 10.6151
R1059 B.n262 B.n261 10.6151
R1060 B.n263 B.n262 10.6151
R1061 B.n263 B.n184 10.6151
R1062 B.n267 B.n184 10.6151
R1063 B.n268 B.n267 10.6151
R1064 B.n269 B.n268 10.6151
R1065 B.n269 B.n182 10.6151
R1066 B.n273 B.n182 10.6151
R1067 B.n274 B.n273 10.6151
R1068 B.n275 B.n274 10.6151
R1069 B.n275 B.n180 10.6151
R1070 B.n279 B.n180 10.6151
R1071 B.n280 B.n279 10.6151
R1072 B.n281 B.n280 10.6151
R1073 B.n281 B.n178 10.6151
R1074 B.n285 B.n178 10.6151
R1075 B.n286 B.n285 10.6151
R1076 B.n287 B.n286 10.6151
R1077 B.n287 B.n176 10.6151
R1078 B.n291 B.n176 10.6151
R1079 B.n292 B.n291 10.6151
R1080 B.n293 B.n292 10.6151
R1081 B.n293 B.n174 10.6151
R1082 B.n297 B.n174 10.6151
R1083 B.n298 B.n297 10.6151
R1084 B.n299 B.n298 10.6151
R1085 B.n299 B.n172 10.6151
R1086 B.n303 B.n172 10.6151
R1087 B.n304 B.n303 10.6151
R1088 B.n305 B.n304 10.6151
R1089 B.n305 B.n170 10.6151
R1090 B.n309 B.n170 10.6151
R1091 B.n310 B.n309 10.6151
R1092 B.n311 B.n310 10.6151
R1093 B.n311 B.n168 10.6151
R1094 B.n315 B.n168 10.6151
R1095 B.n316 B.n315 10.6151
R1096 B.n317 B.n316 10.6151
R1097 B.n317 B.n166 10.6151
R1098 B.n321 B.n166 10.6151
R1099 B.n322 B.n321 10.6151
R1100 B.n323 B.n322 10.6151
R1101 B.n323 B.n164 10.6151
R1102 B.n327 B.n164 10.6151
R1103 B.n328 B.n327 10.6151
R1104 B.n329 B.n328 10.6151
R1105 B.n329 B.n162 10.6151
R1106 B.n333 B.n162 10.6151
R1107 B.n334 B.n333 10.6151
R1108 B.n335 B.n334 10.6151
R1109 B.n335 B.n160 10.6151
R1110 B.n339 B.n160 10.6151
R1111 B.n340 B.n339 10.6151
R1112 B.n342 B.n156 10.6151
R1113 B.n346 B.n156 10.6151
R1114 B.n347 B.n346 10.6151
R1115 B.n348 B.n347 10.6151
R1116 B.n348 B.n154 10.6151
R1117 B.n352 B.n154 10.6151
R1118 B.n353 B.n352 10.6151
R1119 B.n354 B.n353 10.6151
R1120 B.n358 B.n357 10.6151
R1121 B.n359 B.n358 10.6151
R1122 B.n359 B.n148 10.6151
R1123 B.n363 B.n148 10.6151
R1124 B.n364 B.n363 10.6151
R1125 B.n365 B.n364 10.6151
R1126 B.n365 B.n146 10.6151
R1127 B.n369 B.n146 10.6151
R1128 B.n370 B.n369 10.6151
R1129 B.n371 B.n370 10.6151
R1130 B.n371 B.n144 10.6151
R1131 B.n375 B.n144 10.6151
R1132 B.n376 B.n375 10.6151
R1133 B.n377 B.n376 10.6151
R1134 B.n377 B.n142 10.6151
R1135 B.n381 B.n142 10.6151
R1136 B.n382 B.n381 10.6151
R1137 B.n383 B.n382 10.6151
R1138 B.n383 B.n140 10.6151
R1139 B.n387 B.n140 10.6151
R1140 B.n388 B.n387 10.6151
R1141 B.n389 B.n388 10.6151
R1142 B.n389 B.n138 10.6151
R1143 B.n393 B.n138 10.6151
R1144 B.n394 B.n393 10.6151
R1145 B.n395 B.n394 10.6151
R1146 B.n395 B.n136 10.6151
R1147 B.n399 B.n136 10.6151
R1148 B.n400 B.n399 10.6151
R1149 B.n401 B.n400 10.6151
R1150 B.n401 B.n134 10.6151
R1151 B.n405 B.n134 10.6151
R1152 B.n406 B.n405 10.6151
R1153 B.n407 B.n406 10.6151
R1154 B.n407 B.n132 10.6151
R1155 B.n411 B.n132 10.6151
R1156 B.n412 B.n411 10.6151
R1157 B.n413 B.n412 10.6151
R1158 B.n413 B.n130 10.6151
R1159 B.n417 B.n130 10.6151
R1160 B.n418 B.n417 10.6151
R1161 B.n419 B.n418 10.6151
R1162 B.n419 B.n128 10.6151
R1163 B.n423 B.n128 10.6151
R1164 B.n424 B.n423 10.6151
R1165 B.n425 B.n424 10.6151
R1166 B.n425 B.n126 10.6151
R1167 B.n429 B.n126 10.6151
R1168 B.n430 B.n429 10.6151
R1169 B.n431 B.n430 10.6151
R1170 B.n431 B.n124 10.6151
R1171 B.n435 B.n124 10.6151
R1172 B.n436 B.n435 10.6151
R1173 B.n437 B.n436 10.6151
R1174 B.n437 B.n122 10.6151
R1175 B.n441 B.n122 10.6151
R1176 B.n442 B.n441 10.6151
R1177 B.n443 B.n442 10.6151
R1178 B.n443 B.n120 10.6151
R1179 B.n447 B.n120 10.6151
R1180 B.n448 B.n447 10.6151
R1181 B.n449 B.n448 10.6151
R1182 B.n789 B.n0 8.11757
R1183 B.n789 B.n1 8.11757
R1184 B.n648 B.n50 6.5566
R1185 B.n636 B.n635 6.5566
R1186 B.n342 B.n341 6.5566
R1187 B.n354 B.n152 6.5566
R1188 B.n651 B.n50 4.05904
R1189 B.n635 B.n634 4.05904
R1190 B.n341 B.n340 4.05904
R1191 B.n357 B.n152 4.05904
R1192 VP.n6 VP.t1 339.288
R1193 VP.n17 VP.t4 308.801
R1194 VP.n24 VP.t2 308.801
R1195 VP.n31 VP.t3 308.801
R1196 VP.n14 VP.t5 308.801
R1197 VP.n7 VP.t0 308.801
R1198 VP.n17 VP.n16 181.958
R1199 VP.n32 VP.n31 181.958
R1200 VP.n15 VP.n14 181.958
R1201 VP.n9 VP.n8 161.3
R1202 VP.n10 VP.n5 161.3
R1203 VP.n12 VP.n11 161.3
R1204 VP.n13 VP.n4 161.3
R1205 VP.n30 VP.n0 161.3
R1206 VP.n29 VP.n28 161.3
R1207 VP.n27 VP.n1 161.3
R1208 VP.n26 VP.n25 161.3
R1209 VP.n23 VP.n2 161.3
R1210 VP.n22 VP.n21 161.3
R1211 VP.n20 VP.n3 161.3
R1212 VP.n19 VP.n18 161.3
R1213 VP.n22 VP.n3 56.5617
R1214 VP.n29 VP.n1 56.5617
R1215 VP.n12 VP.n5 56.5617
R1216 VP.n7 VP.n6 53.6855
R1217 VP.n16 VP.n15 49.6634
R1218 VP.n18 VP.n3 24.5923
R1219 VP.n23 VP.n22 24.5923
R1220 VP.n25 VP.n1 24.5923
R1221 VP.n30 VP.n29 24.5923
R1222 VP.n13 VP.n12 24.5923
R1223 VP.n8 VP.n5 24.5923
R1224 VP.n9 VP.n6 18.3622
R1225 VP.n24 VP.n23 12.2964
R1226 VP.n25 VP.n24 12.2964
R1227 VP.n8 VP.n7 12.2964
R1228 VP.n18 VP.n17 3.93519
R1229 VP.n31 VP.n30 3.93519
R1230 VP.n14 VP.n13 3.93519
R1231 VP.n10 VP.n9 0.189894
R1232 VP.n11 VP.n10 0.189894
R1233 VP.n11 VP.n4 0.189894
R1234 VP.n15 VP.n4 0.189894
R1235 VP.n19 VP.n16 0.189894
R1236 VP.n20 VP.n19 0.189894
R1237 VP.n21 VP.n20 0.189894
R1238 VP.n21 VP.n2 0.189894
R1239 VP.n26 VP.n2 0.189894
R1240 VP.n27 VP.n26 0.189894
R1241 VP.n28 VP.n27 0.189894
R1242 VP.n28 VP.n0 0.189894
R1243 VP.n32 VP.n0 0.189894
R1244 VP VP.n32 0.0516364
R1245 VDD1 VDD1.t4 69.2371
R1246 VDD1.n1 VDD1.t2 69.1233
R1247 VDD1.n1 VDD1.n0 66.6435
R1248 VDD1.n3 VDD1.n2 66.3043
R1249 VDD1.n3 VDD1.n1 46.7832
R1250 VDD1.n2 VDD1.t3 1.69171
R1251 VDD1.n2 VDD1.t0 1.69171
R1252 VDD1.n0 VDD1.t5 1.69171
R1253 VDD1.n0 VDD1.t1 1.69171
R1254 VDD1 VDD1.n3 0.336707
R1255 VTAIL.n7 VTAIL.t2 51.3169
R1256 VTAIL.n11 VTAIL.t5 51.3167
R1257 VTAIL.n2 VTAIL.t8 51.3167
R1258 VTAIL.n10 VTAIL.t6 51.3167
R1259 VTAIL.n9 VTAIL.n8 49.6257
R1260 VTAIL.n6 VTAIL.n5 49.6257
R1261 VTAIL.n1 VTAIL.n0 49.6257
R1262 VTAIL.n4 VTAIL.n3 49.6257
R1263 VTAIL.n6 VTAIL.n4 32.091
R1264 VTAIL.n11 VTAIL.n10 30.5134
R1265 VTAIL.n0 VTAIL.t1 1.69171
R1266 VTAIL.n0 VTAIL.t4 1.69171
R1267 VTAIL.n3 VTAIL.t7 1.69171
R1268 VTAIL.n3 VTAIL.t9 1.69171
R1269 VTAIL.n8 VTAIL.t10 1.69171
R1270 VTAIL.n8 VTAIL.t11 1.69171
R1271 VTAIL.n5 VTAIL.t0 1.69171
R1272 VTAIL.n5 VTAIL.t3 1.69171
R1273 VTAIL.n7 VTAIL.n6 1.57809
R1274 VTAIL.n10 VTAIL.n9 1.57809
R1275 VTAIL.n4 VTAIL.n2 1.57809
R1276 VTAIL.n9 VTAIL.n7 1.25912
R1277 VTAIL.n2 VTAIL.n1 1.25912
R1278 VTAIL VTAIL.n11 1.1255
R1279 VTAIL VTAIL.n1 0.453086
R1280 VN.n2 VN.t4 339.288
R1281 VN.n14 VN.t1 339.288
R1282 VN.n3 VN.t2 308.801
R1283 VN.n10 VN.t3 308.801
R1284 VN.n15 VN.t0 308.801
R1285 VN.n22 VN.t5 308.801
R1286 VN.n11 VN.n10 181.958
R1287 VN.n23 VN.n22 181.958
R1288 VN.n21 VN.n12 161.3
R1289 VN.n20 VN.n19 161.3
R1290 VN.n18 VN.n13 161.3
R1291 VN.n17 VN.n16 161.3
R1292 VN.n9 VN.n0 161.3
R1293 VN.n8 VN.n7 161.3
R1294 VN.n6 VN.n1 161.3
R1295 VN.n5 VN.n4 161.3
R1296 VN.n8 VN.n1 56.5617
R1297 VN.n20 VN.n13 56.5617
R1298 VN.n3 VN.n2 53.6855
R1299 VN.n15 VN.n14 53.6855
R1300 VN VN.n23 50.0441
R1301 VN.n4 VN.n1 24.5923
R1302 VN.n9 VN.n8 24.5923
R1303 VN.n16 VN.n13 24.5923
R1304 VN.n21 VN.n20 24.5923
R1305 VN.n17 VN.n14 18.3622
R1306 VN.n5 VN.n2 18.3622
R1307 VN.n4 VN.n3 12.2964
R1308 VN.n16 VN.n15 12.2964
R1309 VN.n10 VN.n9 3.93519
R1310 VN.n22 VN.n21 3.93519
R1311 VN.n23 VN.n12 0.189894
R1312 VN.n19 VN.n12 0.189894
R1313 VN.n19 VN.n18 0.189894
R1314 VN.n18 VN.n17 0.189894
R1315 VN.n6 VN.n5 0.189894
R1316 VN.n7 VN.n6 0.189894
R1317 VN.n7 VN.n0 0.189894
R1318 VN.n11 VN.n0 0.189894
R1319 VN VN.n11 0.0516364
R1320 VDD2.n1 VDD2.t1 69.1233
R1321 VDD2.n2 VDD2.t0 67.9957
R1322 VDD2.n1 VDD2.n0 66.6435
R1323 VDD2 VDD2.n3 66.6405
R1324 VDD2.n2 VDD2.n1 45.4114
R1325 VDD2.n3 VDD2.t5 1.69171
R1326 VDD2.n3 VDD2.t4 1.69171
R1327 VDD2.n0 VDD2.t3 1.69171
R1328 VDD2.n0 VDD2.t2 1.69171
R1329 VDD2 VDD2.n2 1.24188
C0 VDD1 w_n2434_n4812# 2.53686f
C1 w_n2434_n4812# B 10.1814f
C2 VDD2 VN 9.196879f
C3 w_n2434_n4812# VN 4.48242f
C4 VDD1 B 2.34526f
C5 VDD1 VN 0.149626f
C6 VN B 1.02208f
C7 VDD2 VP 0.36639f
C8 VDD2 VTAIL 11.339299f
C9 w_n2434_n4812# VP 4.79403f
C10 w_n2434_n4812# VTAIL 3.96737f
C11 VDD1 VP 9.40812f
C12 VP B 1.53682f
C13 VDD1 VTAIL 11.300099f
C14 VTAIL B 4.64547f
C15 VP VN 7.19489f
C16 VN VTAIL 8.80895f
C17 VDD2 w_n2434_n4812# 2.58652f
C18 VP VTAIL 8.823559f
C19 VDD2 VDD1 1.00888f
C20 VDD2 B 2.39309f
C21 VDD2 VSUBS 1.85124f
C22 VDD1 VSUBS 2.241148f
C23 VTAIL VSUBS 1.230127f
C24 VN VSUBS 5.30379f
C25 VP VSUBS 2.337616f
C26 B VSUBS 4.16202f
C27 w_n2434_n4812# VSUBS 0.14309p
C28 VDD2.t1 VSUBS 4.41906f
C29 VDD2.t3 VSUBS 0.407235f
C30 VDD2.t2 VSUBS 0.407235f
C31 VDD2.n0 VSUBS 3.40179f
C32 VDD2.n1 VSUBS 3.76311f
C33 VDD2.t0 VSUBS 4.40673f
C34 VDD2.n2 VSUBS 3.6248f
C35 VDD2.t5 VSUBS 0.407235f
C36 VDD2.t4 VSUBS 0.407235f
C37 VDD2.n3 VSUBS 3.40173f
C38 VN.n0 VSUBS 0.03708f
C39 VN.t3 VSUBS 2.94394f
C40 VN.n1 VSUBS 0.045181f
C41 VN.t4 VSUBS 3.04938f
C42 VN.n2 VSUBS 1.12799f
C43 VN.t2 VSUBS 2.94394f
C44 VN.n3 VSUBS 1.10111f
C45 VN.n4 VSUBS 0.051789f
C46 VN.n5 VSUBS 0.230787f
C47 VN.n6 VSUBS 0.03708f
C48 VN.n7 VSUBS 0.03708f
C49 VN.n8 VSUBS 0.062622f
C50 VN.n9 VSUBS 0.040247f
C51 VN.n10 VSUBS 1.09835f
C52 VN.n11 VSUBS 0.037159f
C53 VN.n12 VSUBS 0.03708f
C54 VN.t5 VSUBS 2.94394f
C55 VN.n13 VSUBS 0.045181f
C56 VN.t1 VSUBS 3.04938f
C57 VN.n14 VSUBS 1.12799f
C58 VN.t0 VSUBS 2.94394f
C59 VN.n15 VSUBS 1.10111f
C60 VN.n16 VSUBS 0.051789f
C61 VN.n17 VSUBS 0.230787f
C62 VN.n18 VSUBS 0.03708f
C63 VN.n19 VSUBS 0.03708f
C64 VN.n20 VSUBS 0.062622f
C65 VN.n21 VSUBS 0.040247f
C66 VN.n22 VSUBS 1.09835f
C67 VN.n23 VSUBS 2.02802f
C68 VTAIL.t1 VSUBS 0.409924f
C69 VTAIL.t4 VSUBS 0.409924f
C70 VTAIL.n0 VSUBS 3.23789f
C71 VTAIL.n1 VSUBS 0.843411f
C72 VTAIL.t8 VSUBS 4.22581f
C73 VTAIL.n2 VSUBS 1.0713f
C74 VTAIL.t7 VSUBS 0.409924f
C75 VTAIL.t9 VSUBS 0.409924f
C76 VTAIL.n3 VSUBS 3.23789f
C77 VTAIL.n4 VSUBS 2.91375f
C78 VTAIL.t0 VSUBS 0.409924f
C79 VTAIL.t3 VSUBS 0.409924f
C80 VTAIL.n5 VSUBS 3.23789f
C81 VTAIL.n6 VSUBS 2.91375f
C82 VTAIL.t2 VSUBS 4.22582f
C83 VTAIL.n7 VSUBS 1.07129f
C84 VTAIL.t10 VSUBS 0.409924f
C85 VTAIL.t11 VSUBS 0.409924f
C86 VTAIL.n8 VSUBS 3.23789f
C87 VTAIL.n9 VSUBS 0.941248f
C88 VTAIL.t6 VSUBS 4.22581f
C89 VTAIL.n10 VSUBS 2.90661f
C90 VTAIL.t5 VSUBS 4.22581f
C91 VTAIL.n11 VSUBS 2.86725f
C92 VDD1.t4 VSUBS 4.40335f
C93 VDD1.t2 VSUBS 4.40197f
C94 VDD1.t5 VSUBS 0.405659f
C95 VDD1.t1 VSUBS 0.405659f
C96 VDD1.n0 VSUBS 3.38863f
C97 VDD1.n1 VSUBS 3.8548f
C98 VDD1.t3 VSUBS 0.405659f
C99 VDD1.t0 VSUBS 0.405659f
C100 VDD1.n2 VSUBS 3.38495f
C101 VDD1.n3 VSUBS 3.55944f
C102 VP.n0 VSUBS 0.037771f
C103 VP.t3 VSUBS 2.99876f
C104 VP.n1 VSUBS 0.046023f
C105 VP.n2 VSUBS 0.037771f
C106 VP.t2 VSUBS 2.99876f
C107 VP.n3 VSUBS 0.063788f
C108 VP.n4 VSUBS 0.037771f
C109 VP.t5 VSUBS 2.99876f
C110 VP.n5 VSUBS 0.046023f
C111 VP.t1 VSUBS 3.10617f
C112 VP.n6 VSUBS 1.14899f
C113 VP.t0 VSUBS 2.99876f
C114 VP.n7 VSUBS 1.12162f
C115 VP.n8 VSUBS 0.052753f
C116 VP.n9 VSUBS 0.235084f
C117 VP.n10 VSUBS 0.037771f
C118 VP.n11 VSUBS 0.037771f
C119 VP.n12 VSUBS 0.063788f
C120 VP.n13 VSUBS 0.040997f
C121 VP.n14 VSUBS 1.1188f
C122 VP.n15 VSUBS 2.04122f
C123 VP.n16 VSUBS 2.06864f
C124 VP.t4 VSUBS 2.99876f
C125 VP.n17 VSUBS 1.1188f
C126 VP.n18 VSUBS 0.040997f
C127 VP.n19 VSUBS 0.037771f
C128 VP.n20 VSUBS 0.037771f
C129 VP.n21 VSUBS 0.037771f
C130 VP.n22 VSUBS 0.046023f
C131 VP.n23 VSUBS 0.052753f
C132 VP.n24 VSUBS 1.05181f
C133 VP.n25 VSUBS 0.052753f
C134 VP.n26 VSUBS 0.037771f
C135 VP.n27 VSUBS 0.037771f
C136 VP.n28 VSUBS 0.037771f
C137 VP.n29 VSUBS 0.063788f
C138 VP.n30 VSUBS 0.040997f
C139 VP.n31 VSUBS 1.1188f
C140 VP.n32 VSUBS 0.037851f
C141 B.n0 VSUBS 0.006971f
C142 B.n1 VSUBS 0.006971f
C143 B.n2 VSUBS 0.01031f
C144 B.n3 VSUBS 0.007901f
C145 B.n4 VSUBS 0.007901f
C146 B.n5 VSUBS 0.007901f
C147 B.n6 VSUBS 0.007901f
C148 B.n7 VSUBS 0.007901f
C149 B.n8 VSUBS 0.007901f
C150 B.n9 VSUBS 0.007901f
C151 B.n10 VSUBS 0.007901f
C152 B.n11 VSUBS 0.007901f
C153 B.n12 VSUBS 0.007901f
C154 B.n13 VSUBS 0.007901f
C155 B.n14 VSUBS 0.007901f
C156 B.n15 VSUBS 0.007901f
C157 B.n16 VSUBS 0.019111f
C158 B.n17 VSUBS 0.007901f
C159 B.n18 VSUBS 0.007901f
C160 B.n19 VSUBS 0.007901f
C161 B.n20 VSUBS 0.007901f
C162 B.n21 VSUBS 0.007901f
C163 B.n22 VSUBS 0.007901f
C164 B.n23 VSUBS 0.007901f
C165 B.n24 VSUBS 0.007901f
C166 B.n25 VSUBS 0.007901f
C167 B.n26 VSUBS 0.007901f
C168 B.n27 VSUBS 0.007901f
C169 B.n28 VSUBS 0.007901f
C170 B.n29 VSUBS 0.007901f
C171 B.n30 VSUBS 0.007901f
C172 B.n31 VSUBS 0.007901f
C173 B.n32 VSUBS 0.007901f
C174 B.n33 VSUBS 0.007901f
C175 B.n34 VSUBS 0.007901f
C176 B.n35 VSUBS 0.007901f
C177 B.n36 VSUBS 0.007901f
C178 B.n37 VSUBS 0.007901f
C179 B.n38 VSUBS 0.007901f
C180 B.n39 VSUBS 0.007901f
C181 B.n40 VSUBS 0.007901f
C182 B.n41 VSUBS 0.007901f
C183 B.n42 VSUBS 0.007901f
C184 B.n43 VSUBS 0.007901f
C185 B.n44 VSUBS 0.007901f
C186 B.n45 VSUBS 0.007901f
C187 B.n46 VSUBS 0.007901f
C188 B.n47 VSUBS 0.007901f
C189 B.t1 VSUBS 0.735641f
C190 B.t2 VSUBS 0.751551f
C191 B.t0 VSUBS 1.37766f
C192 B.n48 VSUBS 0.328782f
C193 B.n49 VSUBS 0.07629f
C194 B.n50 VSUBS 0.018306f
C195 B.n51 VSUBS 0.007901f
C196 B.n52 VSUBS 0.007901f
C197 B.n53 VSUBS 0.007901f
C198 B.n54 VSUBS 0.007901f
C199 B.n55 VSUBS 0.007901f
C200 B.t10 VSUBS 0.735611f
C201 B.t11 VSUBS 0.751525f
C202 B.t9 VSUBS 1.37766f
C203 B.n56 VSUBS 0.328808f
C204 B.n57 VSUBS 0.07632f
C205 B.n58 VSUBS 0.007901f
C206 B.n59 VSUBS 0.007901f
C207 B.n60 VSUBS 0.007901f
C208 B.n61 VSUBS 0.007901f
C209 B.n62 VSUBS 0.007901f
C210 B.n63 VSUBS 0.007901f
C211 B.n64 VSUBS 0.007901f
C212 B.n65 VSUBS 0.007901f
C213 B.n66 VSUBS 0.007901f
C214 B.n67 VSUBS 0.007901f
C215 B.n68 VSUBS 0.007901f
C216 B.n69 VSUBS 0.007901f
C217 B.n70 VSUBS 0.007901f
C218 B.n71 VSUBS 0.007901f
C219 B.n72 VSUBS 0.007901f
C220 B.n73 VSUBS 0.007901f
C221 B.n74 VSUBS 0.007901f
C222 B.n75 VSUBS 0.007901f
C223 B.n76 VSUBS 0.007901f
C224 B.n77 VSUBS 0.007901f
C225 B.n78 VSUBS 0.007901f
C226 B.n79 VSUBS 0.007901f
C227 B.n80 VSUBS 0.007901f
C228 B.n81 VSUBS 0.007901f
C229 B.n82 VSUBS 0.007901f
C230 B.n83 VSUBS 0.007901f
C231 B.n84 VSUBS 0.007901f
C232 B.n85 VSUBS 0.007901f
C233 B.n86 VSUBS 0.007901f
C234 B.n87 VSUBS 0.007901f
C235 B.n88 VSUBS 0.019929f
C236 B.n89 VSUBS 0.007901f
C237 B.n90 VSUBS 0.007901f
C238 B.n91 VSUBS 0.007901f
C239 B.n92 VSUBS 0.007901f
C240 B.n93 VSUBS 0.007901f
C241 B.n94 VSUBS 0.007901f
C242 B.n95 VSUBS 0.007901f
C243 B.n96 VSUBS 0.007901f
C244 B.n97 VSUBS 0.007901f
C245 B.n98 VSUBS 0.007901f
C246 B.n99 VSUBS 0.007901f
C247 B.n100 VSUBS 0.007901f
C248 B.n101 VSUBS 0.007901f
C249 B.n102 VSUBS 0.007901f
C250 B.n103 VSUBS 0.007901f
C251 B.n104 VSUBS 0.007901f
C252 B.n105 VSUBS 0.007901f
C253 B.n106 VSUBS 0.007901f
C254 B.n107 VSUBS 0.007901f
C255 B.n108 VSUBS 0.007901f
C256 B.n109 VSUBS 0.007901f
C257 B.n110 VSUBS 0.007901f
C258 B.n111 VSUBS 0.007901f
C259 B.n112 VSUBS 0.007901f
C260 B.n113 VSUBS 0.007901f
C261 B.n114 VSUBS 0.007901f
C262 B.n115 VSUBS 0.007901f
C263 B.n116 VSUBS 0.007901f
C264 B.n117 VSUBS 0.007901f
C265 B.n118 VSUBS 0.019971f
C266 B.n119 VSUBS 0.007901f
C267 B.n120 VSUBS 0.007901f
C268 B.n121 VSUBS 0.007901f
C269 B.n122 VSUBS 0.007901f
C270 B.n123 VSUBS 0.007901f
C271 B.n124 VSUBS 0.007901f
C272 B.n125 VSUBS 0.007901f
C273 B.n126 VSUBS 0.007901f
C274 B.n127 VSUBS 0.007901f
C275 B.n128 VSUBS 0.007901f
C276 B.n129 VSUBS 0.007901f
C277 B.n130 VSUBS 0.007901f
C278 B.n131 VSUBS 0.007901f
C279 B.n132 VSUBS 0.007901f
C280 B.n133 VSUBS 0.007901f
C281 B.n134 VSUBS 0.007901f
C282 B.n135 VSUBS 0.007901f
C283 B.n136 VSUBS 0.007901f
C284 B.n137 VSUBS 0.007901f
C285 B.n138 VSUBS 0.007901f
C286 B.n139 VSUBS 0.007901f
C287 B.n140 VSUBS 0.007901f
C288 B.n141 VSUBS 0.007901f
C289 B.n142 VSUBS 0.007901f
C290 B.n143 VSUBS 0.007901f
C291 B.n144 VSUBS 0.007901f
C292 B.n145 VSUBS 0.007901f
C293 B.n146 VSUBS 0.007901f
C294 B.n147 VSUBS 0.007901f
C295 B.n148 VSUBS 0.007901f
C296 B.n149 VSUBS 0.007901f
C297 B.t5 VSUBS 0.735611f
C298 B.t4 VSUBS 0.751525f
C299 B.t3 VSUBS 1.37766f
C300 B.n150 VSUBS 0.328808f
C301 B.n151 VSUBS 0.07632f
C302 B.n152 VSUBS 0.018306f
C303 B.n153 VSUBS 0.007901f
C304 B.n154 VSUBS 0.007901f
C305 B.n155 VSUBS 0.007901f
C306 B.n156 VSUBS 0.007901f
C307 B.n157 VSUBS 0.007901f
C308 B.t8 VSUBS 0.735641f
C309 B.t7 VSUBS 0.751551f
C310 B.t6 VSUBS 1.37766f
C311 B.n158 VSUBS 0.328782f
C312 B.n159 VSUBS 0.07629f
C313 B.n160 VSUBS 0.007901f
C314 B.n161 VSUBS 0.007901f
C315 B.n162 VSUBS 0.007901f
C316 B.n163 VSUBS 0.007901f
C317 B.n164 VSUBS 0.007901f
C318 B.n165 VSUBS 0.007901f
C319 B.n166 VSUBS 0.007901f
C320 B.n167 VSUBS 0.007901f
C321 B.n168 VSUBS 0.007901f
C322 B.n169 VSUBS 0.007901f
C323 B.n170 VSUBS 0.007901f
C324 B.n171 VSUBS 0.007901f
C325 B.n172 VSUBS 0.007901f
C326 B.n173 VSUBS 0.007901f
C327 B.n174 VSUBS 0.007901f
C328 B.n175 VSUBS 0.007901f
C329 B.n176 VSUBS 0.007901f
C330 B.n177 VSUBS 0.007901f
C331 B.n178 VSUBS 0.007901f
C332 B.n179 VSUBS 0.007901f
C333 B.n180 VSUBS 0.007901f
C334 B.n181 VSUBS 0.007901f
C335 B.n182 VSUBS 0.007901f
C336 B.n183 VSUBS 0.007901f
C337 B.n184 VSUBS 0.007901f
C338 B.n185 VSUBS 0.007901f
C339 B.n186 VSUBS 0.007901f
C340 B.n187 VSUBS 0.007901f
C341 B.n188 VSUBS 0.007901f
C342 B.n189 VSUBS 0.007901f
C343 B.n190 VSUBS 0.019929f
C344 B.n191 VSUBS 0.007901f
C345 B.n192 VSUBS 0.007901f
C346 B.n193 VSUBS 0.007901f
C347 B.n194 VSUBS 0.007901f
C348 B.n195 VSUBS 0.007901f
C349 B.n196 VSUBS 0.007901f
C350 B.n197 VSUBS 0.007901f
C351 B.n198 VSUBS 0.007901f
C352 B.n199 VSUBS 0.007901f
C353 B.n200 VSUBS 0.007901f
C354 B.n201 VSUBS 0.007901f
C355 B.n202 VSUBS 0.007901f
C356 B.n203 VSUBS 0.007901f
C357 B.n204 VSUBS 0.007901f
C358 B.n205 VSUBS 0.007901f
C359 B.n206 VSUBS 0.007901f
C360 B.n207 VSUBS 0.007901f
C361 B.n208 VSUBS 0.007901f
C362 B.n209 VSUBS 0.007901f
C363 B.n210 VSUBS 0.007901f
C364 B.n211 VSUBS 0.007901f
C365 B.n212 VSUBS 0.007901f
C366 B.n213 VSUBS 0.007901f
C367 B.n214 VSUBS 0.007901f
C368 B.n215 VSUBS 0.007901f
C369 B.n216 VSUBS 0.007901f
C370 B.n217 VSUBS 0.007901f
C371 B.n218 VSUBS 0.007901f
C372 B.n219 VSUBS 0.007901f
C373 B.n220 VSUBS 0.007901f
C374 B.n221 VSUBS 0.007901f
C375 B.n222 VSUBS 0.007901f
C376 B.n223 VSUBS 0.007901f
C377 B.n224 VSUBS 0.007901f
C378 B.n225 VSUBS 0.007901f
C379 B.n226 VSUBS 0.007901f
C380 B.n227 VSUBS 0.007901f
C381 B.n228 VSUBS 0.007901f
C382 B.n229 VSUBS 0.007901f
C383 B.n230 VSUBS 0.007901f
C384 B.n231 VSUBS 0.007901f
C385 B.n232 VSUBS 0.007901f
C386 B.n233 VSUBS 0.007901f
C387 B.n234 VSUBS 0.007901f
C388 B.n235 VSUBS 0.007901f
C389 B.n236 VSUBS 0.007901f
C390 B.n237 VSUBS 0.007901f
C391 B.n238 VSUBS 0.007901f
C392 B.n239 VSUBS 0.007901f
C393 B.n240 VSUBS 0.007901f
C394 B.n241 VSUBS 0.007901f
C395 B.n242 VSUBS 0.007901f
C396 B.n243 VSUBS 0.007901f
C397 B.n244 VSUBS 0.007901f
C398 B.n245 VSUBS 0.019111f
C399 B.n246 VSUBS 0.019111f
C400 B.n247 VSUBS 0.019929f
C401 B.n248 VSUBS 0.007901f
C402 B.n249 VSUBS 0.007901f
C403 B.n250 VSUBS 0.007901f
C404 B.n251 VSUBS 0.007901f
C405 B.n252 VSUBS 0.007901f
C406 B.n253 VSUBS 0.007901f
C407 B.n254 VSUBS 0.007901f
C408 B.n255 VSUBS 0.007901f
C409 B.n256 VSUBS 0.007901f
C410 B.n257 VSUBS 0.007901f
C411 B.n258 VSUBS 0.007901f
C412 B.n259 VSUBS 0.007901f
C413 B.n260 VSUBS 0.007901f
C414 B.n261 VSUBS 0.007901f
C415 B.n262 VSUBS 0.007901f
C416 B.n263 VSUBS 0.007901f
C417 B.n264 VSUBS 0.007901f
C418 B.n265 VSUBS 0.007901f
C419 B.n266 VSUBS 0.007901f
C420 B.n267 VSUBS 0.007901f
C421 B.n268 VSUBS 0.007901f
C422 B.n269 VSUBS 0.007901f
C423 B.n270 VSUBS 0.007901f
C424 B.n271 VSUBS 0.007901f
C425 B.n272 VSUBS 0.007901f
C426 B.n273 VSUBS 0.007901f
C427 B.n274 VSUBS 0.007901f
C428 B.n275 VSUBS 0.007901f
C429 B.n276 VSUBS 0.007901f
C430 B.n277 VSUBS 0.007901f
C431 B.n278 VSUBS 0.007901f
C432 B.n279 VSUBS 0.007901f
C433 B.n280 VSUBS 0.007901f
C434 B.n281 VSUBS 0.007901f
C435 B.n282 VSUBS 0.007901f
C436 B.n283 VSUBS 0.007901f
C437 B.n284 VSUBS 0.007901f
C438 B.n285 VSUBS 0.007901f
C439 B.n286 VSUBS 0.007901f
C440 B.n287 VSUBS 0.007901f
C441 B.n288 VSUBS 0.007901f
C442 B.n289 VSUBS 0.007901f
C443 B.n290 VSUBS 0.007901f
C444 B.n291 VSUBS 0.007901f
C445 B.n292 VSUBS 0.007901f
C446 B.n293 VSUBS 0.007901f
C447 B.n294 VSUBS 0.007901f
C448 B.n295 VSUBS 0.007901f
C449 B.n296 VSUBS 0.007901f
C450 B.n297 VSUBS 0.007901f
C451 B.n298 VSUBS 0.007901f
C452 B.n299 VSUBS 0.007901f
C453 B.n300 VSUBS 0.007901f
C454 B.n301 VSUBS 0.007901f
C455 B.n302 VSUBS 0.007901f
C456 B.n303 VSUBS 0.007901f
C457 B.n304 VSUBS 0.007901f
C458 B.n305 VSUBS 0.007901f
C459 B.n306 VSUBS 0.007901f
C460 B.n307 VSUBS 0.007901f
C461 B.n308 VSUBS 0.007901f
C462 B.n309 VSUBS 0.007901f
C463 B.n310 VSUBS 0.007901f
C464 B.n311 VSUBS 0.007901f
C465 B.n312 VSUBS 0.007901f
C466 B.n313 VSUBS 0.007901f
C467 B.n314 VSUBS 0.007901f
C468 B.n315 VSUBS 0.007901f
C469 B.n316 VSUBS 0.007901f
C470 B.n317 VSUBS 0.007901f
C471 B.n318 VSUBS 0.007901f
C472 B.n319 VSUBS 0.007901f
C473 B.n320 VSUBS 0.007901f
C474 B.n321 VSUBS 0.007901f
C475 B.n322 VSUBS 0.007901f
C476 B.n323 VSUBS 0.007901f
C477 B.n324 VSUBS 0.007901f
C478 B.n325 VSUBS 0.007901f
C479 B.n326 VSUBS 0.007901f
C480 B.n327 VSUBS 0.007901f
C481 B.n328 VSUBS 0.007901f
C482 B.n329 VSUBS 0.007901f
C483 B.n330 VSUBS 0.007901f
C484 B.n331 VSUBS 0.007901f
C485 B.n332 VSUBS 0.007901f
C486 B.n333 VSUBS 0.007901f
C487 B.n334 VSUBS 0.007901f
C488 B.n335 VSUBS 0.007901f
C489 B.n336 VSUBS 0.007901f
C490 B.n337 VSUBS 0.007901f
C491 B.n338 VSUBS 0.007901f
C492 B.n339 VSUBS 0.007901f
C493 B.n340 VSUBS 0.005461f
C494 B.n341 VSUBS 0.018306f
C495 B.n342 VSUBS 0.006391f
C496 B.n343 VSUBS 0.007901f
C497 B.n344 VSUBS 0.007901f
C498 B.n345 VSUBS 0.007901f
C499 B.n346 VSUBS 0.007901f
C500 B.n347 VSUBS 0.007901f
C501 B.n348 VSUBS 0.007901f
C502 B.n349 VSUBS 0.007901f
C503 B.n350 VSUBS 0.007901f
C504 B.n351 VSUBS 0.007901f
C505 B.n352 VSUBS 0.007901f
C506 B.n353 VSUBS 0.007901f
C507 B.n354 VSUBS 0.006391f
C508 B.n355 VSUBS 0.007901f
C509 B.n356 VSUBS 0.007901f
C510 B.n357 VSUBS 0.005461f
C511 B.n358 VSUBS 0.007901f
C512 B.n359 VSUBS 0.007901f
C513 B.n360 VSUBS 0.007901f
C514 B.n361 VSUBS 0.007901f
C515 B.n362 VSUBS 0.007901f
C516 B.n363 VSUBS 0.007901f
C517 B.n364 VSUBS 0.007901f
C518 B.n365 VSUBS 0.007901f
C519 B.n366 VSUBS 0.007901f
C520 B.n367 VSUBS 0.007901f
C521 B.n368 VSUBS 0.007901f
C522 B.n369 VSUBS 0.007901f
C523 B.n370 VSUBS 0.007901f
C524 B.n371 VSUBS 0.007901f
C525 B.n372 VSUBS 0.007901f
C526 B.n373 VSUBS 0.007901f
C527 B.n374 VSUBS 0.007901f
C528 B.n375 VSUBS 0.007901f
C529 B.n376 VSUBS 0.007901f
C530 B.n377 VSUBS 0.007901f
C531 B.n378 VSUBS 0.007901f
C532 B.n379 VSUBS 0.007901f
C533 B.n380 VSUBS 0.007901f
C534 B.n381 VSUBS 0.007901f
C535 B.n382 VSUBS 0.007901f
C536 B.n383 VSUBS 0.007901f
C537 B.n384 VSUBS 0.007901f
C538 B.n385 VSUBS 0.007901f
C539 B.n386 VSUBS 0.007901f
C540 B.n387 VSUBS 0.007901f
C541 B.n388 VSUBS 0.007901f
C542 B.n389 VSUBS 0.007901f
C543 B.n390 VSUBS 0.007901f
C544 B.n391 VSUBS 0.007901f
C545 B.n392 VSUBS 0.007901f
C546 B.n393 VSUBS 0.007901f
C547 B.n394 VSUBS 0.007901f
C548 B.n395 VSUBS 0.007901f
C549 B.n396 VSUBS 0.007901f
C550 B.n397 VSUBS 0.007901f
C551 B.n398 VSUBS 0.007901f
C552 B.n399 VSUBS 0.007901f
C553 B.n400 VSUBS 0.007901f
C554 B.n401 VSUBS 0.007901f
C555 B.n402 VSUBS 0.007901f
C556 B.n403 VSUBS 0.007901f
C557 B.n404 VSUBS 0.007901f
C558 B.n405 VSUBS 0.007901f
C559 B.n406 VSUBS 0.007901f
C560 B.n407 VSUBS 0.007901f
C561 B.n408 VSUBS 0.007901f
C562 B.n409 VSUBS 0.007901f
C563 B.n410 VSUBS 0.007901f
C564 B.n411 VSUBS 0.007901f
C565 B.n412 VSUBS 0.007901f
C566 B.n413 VSUBS 0.007901f
C567 B.n414 VSUBS 0.007901f
C568 B.n415 VSUBS 0.007901f
C569 B.n416 VSUBS 0.007901f
C570 B.n417 VSUBS 0.007901f
C571 B.n418 VSUBS 0.007901f
C572 B.n419 VSUBS 0.007901f
C573 B.n420 VSUBS 0.007901f
C574 B.n421 VSUBS 0.007901f
C575 B.n422 VSUBS 0.007901f
C576 B.n423 VSUBS 0.007901f
C577 B.n424 VSUBS 0.007901f
C578 B.n425 VSUBS 0.007901f
C579 B.n426 VSUBS 0.007901f
C580 B.n427 VSUBS 0.007901f
C581 B.n428 VSUBS 0.007901f
C582 B.n429 VSUBS 0.007901f
C583 B.n430 VSUBS 0.007901f
C584 B.n431 VSUBS 0.007901f
C585 B.n432 VSUBS 0.007901f
C586 B.n433 VSUBS 0.007901f
C587 B.n434 VSUBS 0.007901f
C588 B.n435 VSUBS 0.007901f
C589 B.n436 VSUBS 0.007901f
C590 B.n437 VSUBS 0.007901f
C591 B.n438 VSUBS 0.007901f
C592 B.n439 VSUBS 0.007901f
C593 B.n440 VSUBS 0.007901f
C594 B.n441 VSUBS 0.007901f
C595 B.n442 VSUBS 0.007901f
C596 B.n443 VSUBS 0.007901f
C597 B.n444 VSUBS 0.007901f
C598 B.n445 VSUBS 0.007901f
C599 B.n446 VSUBS 0.007901f
C600 B.n447 VSUBS 0.007901f
C601 B.n448 VSUBS 0.007901f
C602 B.n449 VSUBS 0.019069f
C603 B.n450 VSUBS 0.019929f
C604 B.n451 VSUBS 0.019111f
C605 B.n452 VSUBS 0.007901f
C606 B.n453 VSUBS 0.007901f
C607 B.n454 VSUBS 0.007901f
C608 B.n455 VSUBS 0.007901f
C609 B.n456 VSUBS 0.007901f
C610 B.n457 VSUBS 0.007901f
C611 B.n458 VSUBS 0.007901f
C612 B.n459 VSUBS 0.007901f
C613 B.n460 VSUBS 0.007901f
C614 B.n461 VSUBS 0.007901f
C615 B.n462 VSUBS 0.007901f
C616 B.n463 VSUBS 0.007901f
C617 B.n464 VSUBS 0.007901f
C618 B.n465 VSUBS 0.007901f
C619 B.n466 VSUBS 0.007901f
C620 B.n467 VSUBS 0.007901f
C621 B.n468 VSUBS 0.007901f
C622 B.n469 VSUBS 0.007901f
C623 B.n470 VSUBS 0.007901f
C624 B.n471 VSUBS 0.007901f
C625 B.n472 VSUBS 0.007901f
C626 B.n473 VSUBS 0.007901f
C627 B.n474 VSUBS 0.007901f
C628 B.n475 VSUBS 0.007901f
C629 B.n476 VSUBS 0.007901f
C630 B.n477 VSUBS 0.007901f
C631 B.n478 VSUBS 0.007901f
C632 B.n479 VSUBS 0.007901f
C633 B.n480 VSUBS 0.007901f
C634 B.n481 VSUBS 0.007901f
C635 B.n482 VSUBS 0.007901f
C636 B.n483 VSUBS 0.007901f
C637 B.n484 VSUBS 0.007901f
C638 B.n485 VSUBS 0.007901f
C639 B.n486 VSUBS 0.007901f
C640 B.n487 VSUBS 0.007901f
C641 B.n488 VSUBS 0.007901f
C642 B.n489 VSUBS 0.007901f
C643 B.n490 VSUBS 0.007901f
C644 B.n491 VSUBS 0.007901f
C645 B.n492 VSUBS 0.007901f
C646 B.n493 VSUBS 0.007901f
C647 B.n494 VSUBS 0.007901f
C648 B.n495 VSUBS 0.007901f
C649 B.n496 VSUBS 0.007901f
C650 B.n497 VSUBS 0.007901f
C651 B.n498 VSUBS 0.007901f
C652 B.n499 VSUBS 0.007901f
C653 B.n500 VSUBS 0.007901f
C654 B.n501 VSUBS 0.007901f
C655 B.n502 VSUBS 0.007901f
C656 B.n503 VSUBS 0.007901f
C657 B.n504 VSUBS 0.007901f
C658 B.n505 VSUBS 0.007901f
C659 B.n506 VSUBS 0.007901f
C660 B.n507 VSUBS 0.007901f
C661 B.n508 VSUBS 0.007901f
C662 B.n509 VSUBS 0.007901f
C663 B.n510 VSUBS 0.007901f
C664 B.n511 VSUBS 0.007901f
C665 B.n512 VSUBS 0.007901f
C666 B.n513 VSUBS 0.007901f
C667 B.n514 VSUBS 0.007901f
C668 B.n515 VSUBS 0.007901f
C669 B.n516 VSUBS 0.007901f
C670 B.n517 VSUBS 0.007901f
C671 B.n518 VSUBS 0.007901f
C672 B.n519 VSUBS 0.007901f
C673 B.n520 VSUBS 0.007901f
C674 B.n521 VSUBS 0.007901f
C675 B.n522 VSUBS 0.007901f
C676 B.n523 VSUBS 0.007901f
C677 B.n524 VSUBS 0.007901f
C678 B.n525 VSUBS 0.007901f
C679 B.n526 VSUBS 0.007901f
C680 B.n527 VSUBS 0.007901f
C681 B.n528 VSUBS 0.007901f
C682 B.n529 VSUBS 0.007901f
C683 B.n530 VSUBS 0.007901f
C684 B.n531 VSUBS 0.007901f
C685 B.n532 VSUBS 0.007901f
C686 B.n533 VSUBS 0.007901f
C687 B.n534 VSUBS 0.007901f
C688 B.n535 VSUBS 0.007901f
C689 B.n536 VSUBS 0.007901f
C690 B.n537 VSUBS 0.007901f
C691 B.n538 VSUBS 0.007901f
C692 B.n539 VSUBS 0.019111f
C693 B.n540 VSUBS 0.019111f
C694 B.n541 VSUBS 0.019929f
C695 B.n542 VSUBS 0.007901f
C696 B.n543 VSUBS 0.007901f
C697 B.n544 VSUBS 0.007901f
C698 B.n545 VSUBS 0.007901f
C699 B.n546 VSUBS 0.007901f
C700 B.n547 VSUBS 0.007901f
C701 B.n548 VSUBS 0.007901f
C702 B.n549 VSUBS 0.007901f
C703 B.n550 VSUBS 0.007901f
C704 B.n551 VSUBS 0.007901f
C705 B.n552 VSUBS 0.007901f
C706 B.n553 VSUBS 0.007901f
C707 B.n554 VSUBS 0.007901f
C708 B.n555 VSUBS 0.007901f
C709 B.n556 VSUBS 0.007901f
C710 B.n557 VSUBS 0.007901f
C711 B.n558 VSUBS 0.007901f
C712 B.n559 VSUBS 0.007901f
C713 B.n560 VSUBS 0.007901f
C714 B.n561 VSUBS 0.007901f
C715 B.n562 VSUBS 0.007901f
C716 B.n563 VSUBS 0.007901f
C717 B.n564 VSUBS 0.007901f
C718 B.n565 VSUBS 0.007901f
C719 B.n566 VSUBS 0.007901f
C720 B.n567 VSUBS 0.007901f
C721 B.n568 VSUBS 0.007901f
C722 B.n569 VSUBS 0.007901f
C723 B.n570 VSUBS 0.007901f
C724 B.n571 VSUBS 0.007901f
C725 B.n572 VSUBS 0.007901f
C726 B.n573 VSUBS 0.007901f
C727 B.n574 VSUBS 0.007901f
C728 B.n575 VSUBS 0.007901f
C729 B.n576 VSUBS 0.007901f
C730 B.n577 VSUBS 0.007901f
C731 B.n578 VSUBS 0.007901f
C732 B.n579 VSUBS 0.007901f
C733 B.n580 VSUBS 0.007901f
C734 B.n581 VSUBS 0.007901f
C735 B.n582 VSUBS 0.007901f
C736 B.n583 VSUBS 0.007901f
C737 B.n584 VSUBS 0.007901f
C738 B.n585 VSUBS 0.007901f
C739 B.n586 VSUBS 0.007901f
C740 B.n587 VSUBS 0.007901f
C741 B.n588 VSUBS 0.007901f
C742 B.n589 VSUBS 0.007901f
C743 B.n590 VSUBS 0.007901f
C744 B.n591 VSUBS 0.007901f
C745 B.n592 VSUBS 0.007901f
C746 B.n593 VSUBS 0.007901f
C747 B.n594 VSUBS 0.007901f
C748 B.n595 VSUBS 0.007901f
C749 B.n596 VSUBS 0.007901f
C750 B.n597 VSUBS 0.007901f
C751 B.n598 VSUBS 0.007901f
C752 B.n599 VSUBS 0.007901f
C753 B.n600 VSUBS 0.007901f
C754 B.n601 VSUBS 0.007901f
C755 B.n602 VSUBS 0.007901f
C756 B.n603 VSUBS 0.007901f
C757 B.n604 VSUBS 0.007901f
C758 B.n605 VSUBS 0.007901f
C759 B.n606 VSUBS 0.007901f
C760 B.n607 VSUBS 0.007901f
C761 B.n608 VSUBS 0.007901f
C762 B.n609 VSUBS 0.007901f
C763 B.n610 VSUBS 0.007901f
C764 B.n611 VSUBS 0.007901f
C765 B.n612 VSUBS 0.007901f
C766 B.n613 VSUBS 0.007901f
C767 B.n614 VSUBS 0.007901f
C768 B.n615 VSUBS 0.007901f
C769 B.n616 VSUBS 0.007901f
C770 B.n617 VSUBS 0.007901f
C771 B.n618 VSUBS 0.007901f
C772 B.n619 VSUBS 0.007901f
C773 B.n620 VSUBS 0.007901f
C774 B.n621 VSUBS 0.007901f
C775 B.n622 VSUBS 0.007901f
C776 B.n623 VSUBS 0.007901f
C777 B.n624 VSUBS 0.007901f
C778 B.n625 VSUBS 0.007901f
C779 B.n626 VSUBS 0.007901f
C780 B.n627 VSUBS 0.007901f
C781 B.n628 VSUBS 0.007901f
C782 B.n629 VSUBS 0.007901f
C783 B.n630 VSUBS 0.007901f
C784 B.n631 VSUBS 0.007901f
C785 B.n632 VSUBS 0.007901f
C786 B.n633 VSUBS 0.007901f
C787 B.n634 VSUBS 0.005461f
C788 B.n635 VSUBS 0.018306f
C789 B.n636 VSUBS 0.006391f
C790 B.n637 VSUBS 0.007901f
C791 B.n638 VSUBS 0.007901f
C792 B.n639 VSUBS 0.007901f
C793 B.n640 VSUBS 0.007901f
C794 B.n641 VSUBS 0.007901f
C795 B.n642 VSUBS 0.007901f
C796 B.n643 VSUBS 0.007901f
C797 B.n644 VSUBS 0.007901f
C798 B.n645 VSUBS 0.007901f
C799 B.n646 VSUBS 0.007901f
C800 B.n647 VSUBS 0.007901f
C801 B.n648 VSUBS 0.006391f
C802 B.n649 VSUBS 0.007901f
C803 B.n650 VSUBS 0.007901f
C804 B.n651 VSUBS 0.005461f
C805 B.n652 VSUBS 0.007901f
C806 B.n653 VSUBS 0.007901f
C807 B.n654 VSUBS 0.007901f
C808 B.n655 VSUBS 0.007901f
C809 B.n656 VSUBS 0.007901f
C810 B.n657 VSUBS 0.007901f
C811 B.n658 VSUBS 0.007901f
C812 B.n659 VSUBS 0.007901f
C813 B.n660 VSUBS 0.007901f
C814 B.n661 VSUBS 0.007901f
C815 B.n662 VSUBS 0.007901f
C816 B.n663 VSUBS 0.007901f
C817 B.n664 VSUBS 0.007901f
C818 B.n665 VSUBS 0.007901f
C819 B.n666 VSUBS 0.007901f
C820 B.n667 VSUBS 0.007901f
C821 B.n668 VSUBS 0.007901f
C822 B.n669 VSUBS 0.007901f
C823 B.n670 VSUBS 0.007901f
C824 B.n671 VSUBS 0.007901f
C825 B.n672 VSUBS 0.007901f
C826 B.n673 VSUBS 0.007901f
C827 B.n674 VSUBS 0.007901f
C828 B.n675 VSUBS 0.007901f
C829 B.n676 VSUBS 0.007901f
C830 B.n677 VSUBS 0.007901f
C831 B.n678 VSUBS 0.007901f
C832 B.n679 VSUBS 0.007901f
C833 B.n680 VSUBS 0.007901f
C834 B.n681 VSUBS 0.007901f
C835 B.n682 VSUBS 0.007901f
C836 B.n683 VSUBS 0.007901f
C837 B.n684 VSUBS 0.007901f
C838 B.n685 VSUBS 0.007901f
C839 B.n686 VSUBS 0.007901f
C840 B.n687 VSUBS 0.007901f
C841 B.n688 VSUBS 0.007901f
C842 B.n689 VSUBS 0.007901f
C843 B.n690 VSUBS 0.007901f
C844 B.n691 VSUBS 0.007901f
C845 B.n692 VSUBS 0.007901f
C846 B.n693 VSUBS 0.007901f
C847 B.n694 VSUBS 0.007901f
C848 B.n695 VSUBS 0.007901f
C849 B.n696 VSUBS 0.007901f
C850 B.n697 VSUBS 0.007901f
C851 B.n698 VSUBS 0.007901f
C852 B.n699 VSUBS 0.007901f
C853 B.n700 VSUBS 0.007901f
C854 B.n701 VSUBS 0.007901f
C855 B.n702 VSUBS 0.007901f
C856 B.n703 VSUBS 0.007901f
C857 B.n704 VSUBS 0.007901f
C858 B.n705 VSUBS 0.007901f
C859 B.n706 VSUBS 0.007901f
C860 B.n707 VSUBS 0.007901f
C861 B.n708 VSUBS 0.007901f
C862 B.n709 VSUBS 0.007901f
C863 B.n710 VSUBS 0.007901f
C864 B.n711 VSUBS 0.007901f
C865 B.n712 VSUBS 0.007901f
C866 B.n713 VSUBS 0.007901f
C867 B.n714 VSUBS 0.007901f
C868 B.n715 VSUBS 0.007901f
C869 B.n716 VSUBS 0.007901f
C870 B.n717 VSUBS 0.007901f
C871 B.n718 VSUBS 0.007901f
C872 B.n719 VSUBS 0.007901f
C873 B.n720 VSUBS 0.007901f
C874 B.n721 VSUBS 0.007901f
C875 B.n722 VSUBS 0.007901f
C876 B.n723 VSUBS 0.007901f
C877 B.n724 VSUBS 0.007901f
C878 B.n725 VSUBS 0.007901f
C879 B.n726 VSUBS 0.007901f
C880 B.n727 VSUBS 0.007901f
C881 B.n728 VSUBS 0.007901f
C882 B.n729 VSUBS 0.007901f
C883 B.n730 VSUBS 0.007901f
C884 B.n731 VSUBS 0.007901f
C885 B.n732 VSUBS 0.007901f
C886 B.n733 VSUBS 0.007901f
C887 B.n734 VSUBS 0.007901f
C888 B.n735 VSUBS 0.007901f
C889 B.n736 VSUBS 0.007901f
C890 B.n737 VSUBS 0.007901f
C891 B.n738 VSUBS 0.007901f
C892 B.n739 VSUBS 0.007901f
C893 B.n740 VSUBS 0.007901f
C894 B.n741 VSUBS 0.007901f
C895 B.n742 VSUBS 0.007901f
C896 B.n743 VSUBS 0.019929f
C897 B.n744 VSUBS 0.019929f
C898 B.n745 VSUBS 0.019111f
C899 B.n746 VSUBS 0.007901f
C900 B.n747 VSUBS 0.007901f
C901 B.n748 VSUBS 0.007901f
C902 B.n749 VSUBS 0.007901f
C903 B.n750 VSUBS 0.007901f
C904 B.n751 VSUBS 0.007901f
C905 B.n752 VSUBS 0.007901f
C906 B.n753 VSUBS 0.007901f
C907 B.n754 VSUBS 0.007901f
C908 B.n755 VSUBS 0.007901f
C909 B.n756 VSUBS 0.007901f
C910 B.n757 VSUBS 0.007901f
C911 B.n758 VSUBS 0.007901f
C912 B.n759 VSUBS 0.007901f
C913 B.n760 VSUBS 0.007901f
C914 B.n761 VSUBS 0.007901f
C915 B.n762 VSUBS 0.007901f
C916 B.n763 VSUBS 0.007901f
C917 B.n764 VSUBS 0.007901f
C918 B.n765 VSUBS 0.007901f
C919 B.n766 VSUBS 0.007901f
C920 B.n767 VSUBS 0.007901f
C921 B.n768 VSUBS 0.007901f
C922 B.n769 VSUBS 0.007901f
C923 B.n770 VSUBS 0.007901f
C924 B.n771 VSUBS 0.007901f
C925 B.n772 VSUBS 0.007901f
C926 B.n773 VSUBS 0.007901f
C927 B.n774 VSUBS 0.007901f
C928 B.n775 VSUBS 0.007901f
C929 B.n776 VSUBS 0.007901f
C930 B.n777 VSUBS 0.007901f
C931 B.n778 VSUBS 0.007901f
C932 B.n779 VSUBS 0.007901f
C933 B.n780 VSUBS 0.007901f
C934 B.n781 VSUBS 0.007901f
C935 B.n782 VSUBS 0.007901f
C936 B.n783 VSUBS 0.007901f
C937 B.n784 VSUBS 0.007901f
C938 B.n785 VSUBS 0.007901f
C939 B.n786 VSUBS 0.007901f
C940 B.n787 VSUBS 0.01031f
C941 B.n788 VSUBS 0.010983f
C942 B.n789 VSUBS 0.021841f
.ends

