* NGSPICE file created from diff_pair_sample_0487.ext - technology: sky130A

.subckt diff_pair_sample_0487 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=0 ps=0 w=8.13 l=2.38
X1 VDD1.t7 VP.t0 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=3.1707 ps=17.04 w=8.13 l=2.38
X2 VTAIL.t5 VN.t0 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X3 VDD2.t6 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=3.1707 ps=17.04 w=8.13 l=2.38
X4 VTAIL.t2 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=1.34145 ps=8.46 w=8.13 l=2.38
X5 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=0 ps=0 w=8.13 l=2.38
X7 VTAIL.t1 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=1.34145 ps=8.46 w=8.13 l=2.38
X8 VDD1.t6 VP.t1 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X9 VTAIL.t3 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=0 ps=0 w=8.13 l=2.38
X11 VDD2.t1 VN.t6 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=3.1707 ps=17.04 w=8.13 l=2.38
X12 VDD2.t0 VN.t7 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X13 VTAIL.t11 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X14 VTAIL.t8 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
X15 VDD1.t3 VP.t4 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=3.1707 ps=17.04 w=8.13 l=2.38
X16 VTAIL.t9 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=1.34145 ps=8.46 w=8.13 l=2.38
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=0 ps=0 w=8.13 l=2.38
X18 VTAIL.t10 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1707 pd=17.04 as=1.34145 ps=8.46 w=8.13 l=2.38
X19 VDD1.t0 VP.t7 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=1.34145 pd=8.46 as=1.34145 ps=8.46 w=8.13 l=2.38
R0 B.n746 B.n745 585
R1 B.n265 B.n124 585
R2 B.n264 B.n263 585
R3 B.n262 B.n261 585
R4 B.n260 B.n259 585
R5 B.n258 B.n257 585
R6 B.n256 B.n255 585
R7 B.n254 B.n253 585
R8 B.n252 B.n251 585
R9 B.n250 B.n249 585
R10 B.n248 B.n247 585
R11 B.n246 B.n245 585
R12 B.n244 B.n243 585
R13 B.n242 B.n241 585
R14 B.n240 B.n239 585
R15 B.n238 B.n237 585
R16 B.n236 B.n235 585
R17 B.n234 B.n233 585
R18 B.n232 B.n231 585
R19 B.n230 B.n229 585
R20 B.n228 B.n227 585
R21 B.n226 B.n225 585
R22 B.n224 B.n223 585
R23 B.n222 B.n221 585
R24 B.n220 B.n219 585
R25 B.n218 B.n217 585
R26 B.n216 B.n215 585
R27 B.n214 B.n213 585
R28 B.n212 B.n211 585
R29 B.n210 B.n209 585
R30 B.n208 B.n207 585
R31 B.n206 B.n205 585
R32 B.n204 B.n203 585
R33 B.n202 B.n201 585
R34 B.n200 B.n199 585
R35 B.n198 B.n197 585
R36 B.n196 B.n195 585
R37 B.n194 B.n193 585
R38 B.n192 B.n191 585
R39 B.n190 B.n189 585
R40 B.n188 B.n187 585
R41 B.n186 B.n185 585
R42 B.n184 B.n183 585
R43 B.n182 B.n181 585
R44 B.n180 B.n179 585
R45 B.n178 B.n177 585
R46 B.n176 B.n175 585
R47 B.n174 B.n173 585
R48 B.n172 B.n171 585
R49 B.n170 B.n169 585
R50 B.n168 B.n167 585
R51 B.n166 B.n165 585
R52 B.n164 B.n163 585
R53 B.n162 B.n161 585
R54 B.n160 B.n159 585
R55 B.n158 B.n157 585
R56 B.n156 B.n155 585
R57 B.n154 B.n153 585
R58 B.n152 B.n151 585
R59 B.n150 B.n149 585
R60 B.n148 B.n147 585
R61 B.n146 B.n145 585
R62 B.n144 B.n143 585
R63 B.n142 B.n141 585
R64 B.n140 B.n139 585
R65 B.n138 B.n137 585
R66 B.n136 B.n135 585
R67 B.n134 B.n133 585
R68 B.n132 B.n131 585
R69 B.n88 B.n87 585
R70 B.n744 B.n89 585
R71 B.n749 B.n89 585
R72 B.n743 B.n742 585
R73 B.n742 B.n85 585
R74 B.n741 B.n84 585
R75 B.n755 B.n84 585
R76 B.n740 B.n83 585
R77 B.n756 B.n83 585
R78 B.n739 B.n82 585
R79 B.n757 B.n82 585
R80 B.n738 B.n737 585
R81 B.n737 B.n78 585
R82 B.n736 B.n77 585
R83 B.n763 B.n77 585
R84 B.n735 B.n76 585
R85 B.n764 B.n76 585
R86 B.n734 B.n75 585
R87 B.n765 B.n75 585
R88 B.n733 B.n732 585
R89 B.n732 B.n71 585
R90 B.n731 B.n70 585
R91 B.n771 B.n70 585
R92 B.n730 B.n69 585
R93 B.n772 B.n69 585
R94 B.n729 B.n68 585
R95 B.n773 B.n68 585
R96 B.n728 B.n727 585
R97 B.n727 B.n64 585
R98 B.n726 B.n63 585
R99 B.n779 B.n63 585
R100 B.n725 B.n62 585
R101 B.n780 B.n62 585
R102 B.n724 B.n61 585
R103 B.n781 B.n61 585
R104 B.n723 B.n722 585
R105 B.n722 B.n57 585
R106 B.n721 B.n56 585
R107 B.n787 B.n56 585
R108 B.n720 B.n55 585
R109 B.n788 B.n55 585
R110 B.n719 B.n54 585
R111 B.n789 B.n54 585
R112 B.n718 B.n717 585
R113 B.n717 B.n50 585
R114 B.n716 B.n49 585
R115 B.n795 B.n49 585
R116 B.n715 B.n48 585
R117 B.n796 B.n48 585
R118 B.n714 B.n47 585
R119 B.n797 B.n47 585
R120 B.n713 B.n712 585
R121 B.n712 B.n43 585
R122 B.n711 B.n42 585
R123 B.n803 B.n42 585
R124 B.n710 B.n41 585
R125 B.n804 B.n41 585
R126 B.n709 B.n40 585
R127 B.n805 B.n40 585
R128 B.n708 B.n707 585
R129 B.n707 B.n36 585
R130 B.n706 B.n35 585
R131 B.n811 B.n35 585
R132 B.n705 B.n34 585
R133 B.n812 B.n34 585
R134 B.n704 B.n33 585
R135 B.n813 B.n33 585
R136 B.n703 B.n702 585
R137 B.n702 B.n29 585
R138 B.n701 B.n28 585
R139 B.n819 B.n28 585
R140 B.n700 B.n27 585
R141 B.n820 B.n27 585
R142 B.n699 B.n26 585
R143 B.n821 B.n26 585
R144 B.n698 B.n697 585
R145 B.n697 B.n22 585
R146 B.n696 B.n21 585
R147 B.n827 B.n21 585
R148 B.n695 B.n20 585
R149 B.n828 B.n20 585
R150 B.n694 B.n19 585
R151 B.n829 B.n19 585
R152 B.n693 B.n692 585
R153 B.n692 B.n15 585
R154 B.n691 B.n14 585
R155 B.n835 B.n14 585
R156 B.n690 B.n13 585
R157 B.n836 B.n13 585
R158 B.n689 B.n12 585
R159 B.n837 B.n12 585
R160 B.n688 B.n687 585
R161 B.n687 B.n8 585
R162 B.n686 B.n7 585
R163 B.n843 B.n7 585
R164 B.n685 B.n6 585
R165 B.n844 B.n6 585
R166 B.n684 B.n5 585
R167 B.n845 B.n5 585
R168 B.n683 B.n682 585
R169 B.n682 B.n4 585
R170 B.n681 B.n266 585
R171 B.n681 B.n680 585
R172 B.n671 B.n267 585
R173 B.n268 B.n267 585
R174 B.n673 B.n672 585
R175 B.n674 B.n673 585
R176 B.n670 B.n273 585
R177 B.n273 B.n272 585
R178 B.n669 B.n668 585
R179 B.n668 B.n667 585
R180 B.n275 B.n274 585
R181 B.n276 B.n275 585
R182 B.n660 B.n659 585
R183 B.n661 B.n660 585
R184 B.n658 B.n281 585
R185 B.n281 B.n280 585
R186 B.n657 B.n656 585
R187 B.n656 B.n655 585
R188 B.n283 B.n282 585
R189 B.n284 B.n283 585
R190 B.n648 B.n647 585
R191 B.n649 B.n648 585
R192 B.n646 B.n289 585
R193 B.n289 B.n288 585
R194 B.n645 B.n644 585
R195 B.n644 B.n643 585
R196 B.n291 B.n290 585
R197 B.n292 B.n291 585
R198 B.n636 B.n635 585
R199 B.n637 B.n636 585
R200 B.n634 B.n297 585
R201 B.n297 B.n296 585
R202 B.n633 B.n632 585
R203 B.n632 B.n631 585
R204 B.n299 B.n298 585
R205 B.n300 B.n299 585
R206 B.n624 B.n623 585
R207 B.n625 B.n624 585
R208 B.n622 B.n305 585
R209 B.n305 B.n304 585
R210 B.n621 B.n620 585
R211 B.n620 B.n619 585
R212 B.n307 B.n306 585
R213 B.n308 B.n307 585
R214 B.n612 B.n611 585
R215 B.n613 B.n612 585
R216 B.n610 B.n313 585
R217 B.n313 B.n312 585
R218 B.n609 B.n608 585
R219 B.n608 B.n607 585
R220 B.n315 B.n314 585
R221 B.n316 B.n315 585
R222 B.n600 B.n599 585
R223 B.n601 B.n600 585
R224 B.n598 B.n321 585
R225 B.n321 B.n320 585
R226 B.n597 B.n596 585
R227 B.n596 B.n595 585
R228 B.n323 B.n322 585
R229 B.n324 B.n323 585
R230 B.n588 B.n587 585
R231 B.n589 B.n588 585
R232 B.n586 B.n329 585
R233 B.n329 B.n328 585
R234 B.n585 B.n584 585
R235 B.n584 B.n583 585
R236 B.n331 B.n330 585
R237 B.n332 B.n331 585
R238 B.n576 B.n575 585
R239 B.n577 B.n576 585
R240 B.n574 B.n337 585
R241 B.n337 B.n336 585
R242 B.n573 B.n572 585
R243 B.n572 B.n571 585
R244 B.n339 B.n338 585
R245 B.n340 B.n339 585
R246 B.n564 B.n563 585
R247 B.n565 B.n564 585
R248 B.n562 B.n344 585
R249 B.n348 B.n344 585
R250 B.n561 B.n560 585
R251 B.n560 B.n559 585
R252 B.n346 B.n345 585
R253 B.n347 B.n346 585
R254 B.n552 B.n551 585
R255 B.n553 B.n552 585
R256 B.n550 B.n353 585
R257 B.n353 B.n352 585
R258 B.n549 B.n548 585
R259 B.n548 B.n547 585
R260 B.n355 B.n354 585
R261 B.n356 B.n355 585
R262 B.n540 B.n539 585
R263 B.n541 B.n540 585
R264 B.n359 B.n358 585
R265 B.n400 B.n398 585
R266 B.n401 B.n397 585
R267 B.n401 B.n360 585
R268 B.n404 B.n403 585
R269 B.n405 B.n396 585
R270 B.n407 B.n406 585
R271 B.n409 B.n395 585
R272 B.n412 B.n411 585
R273 B.n413 B.n394 585
R274 B.n415 B.n414 585
R275 B.n417 B.n393 585
R276 B.n420 B.n419 585
R277 B.n421 B.n392 585
R278 B.n423 B.n422 585
R279 B.n425 B.n391 585
R280 B.n428 B.n427 585
R281 B.n429 B.n390 585
R282 B.n431 B.n430 585
R283 B.n433 B.n389 585
R284 B.n436 B.n435 585
R285 B.n437 B.n388 585
R286 B.n439 B.n438 585
R287 B.n441 B.n387 585
R288 B.n444 B.n443 585
R289 B.n445 B.n386 585
R290 B.n447 B.n446 585
R291 B.n449 B.n385 585
R292 B.n452 B.n451 585
R293 B.n453 B.n384 585
R294 B.n458 B.n457 585
R295 B.n460 B.n383 585
R296 B.n463 B.n462 585
R297 B.n464 B.n382 585
R298 B.n466 B.n465 585
R299 B.n468 B.n381 585
R300 B.n471 B.n470 585
R301 B.n472 B.n380 585
R302 B.n474 B.n473 585
R303 B.n476 B.n379 585
R304 B.n479 B.n478 585
R305 B.n481 B.n376 585
R306 B.n483 B.n482 585
R307 B.n485 B.n375 585
R308 B.n488 B.n487 585
R309 B.n489 B.n374 585
R310 B.n491 B.n490 585
R311 B.n493 B.n373 585
R312 B.n496 B.n495 585
R313 B.n497 B.n372 585
R314 B.n499 B.n498 585
R315 B.n501 B.n371 585
R316 B.n504 B.n503 585
R317 B.n505 B.n370 585
R318 B.n507 B.n506 585
R319 B.n509 B.n369 585
R320 B.n512 B.n511 585
R321 B.n513 B.n368 585
R322 B.n515 B.n514 585
R323 B.n517 B.n367 585
R324 B.n520 B.n519 585
R325 B.n521 B.n366 585
R326 B.n523 B.n522 585
R327 B.n525 B.n365 585
R328 B.n528 B.n527 585
R329 B.n529 B.n364 585
R330 B.n531 B.n530 585
R331 B.n533 B.n363 585
R332 B.n534 B.n362 585
R333 B.n537 B.n536 585
R334 B.n538 B.n361 585
R335 B.n361 B.n360 585
R336 B.n543 B.n542 585
R337 B.n542 B.n541 585
R338 B.n544 B.n357 585
R339 B.n357 B.n356 585
R340 B.n546 B.n545 585
R341 B.n547 B.n546 585
R342 B.n351 B.n350 585
R343 B.n352 B.n351 585
R344 B.n555 B.n554 585
R345 B.n554 B.n553 585
R346 B.n556 B.n349 585
R347 B.n349 B.n347 585
R348 B.n558 B.n557 585
R349 B.n559 B.n558 585
R350 B.n343 B.n342 585
R351 B.n348 B.n343 585
R352 B.n567 B.n566 585
R353 B.n566 B.n565 585
R354 B.n568 B.n341 585
R355 B.n341 B.n340 585
R356 B.n570 B.n569 585
R357 B.n571 B.n570 585
R358 B.n335 B.n334 585
R359 B.n336 B.n335 585
R360 B.n579 B.n578 585
R361 B.n578 B.n577 585
R362 B.n580 B.n333 585
R363 B.n333 B.n332 585
R364 B.n582 B.n581 585
R365 B.n583 B.n582 585
R366 B.n327 B.n326 585
R367 B.n328 B.n327 585
R368 B.n591 B.n590 585
R369 B.n590 B.n589 585
R370 B.n592 B.n325 585
R371 B.n325 B.n324 585
R372 B.n594 B.n593 585
R373 B.n595 B.n594 585
R374 B.n319 B.n318 585
R375 B.n320 B.n319 585
R376 B.n603 B.n602 585
R377 B.n602 B.n601 585
R378 B.n604 B.n317 585
R379 B.n317 B.n316 585
R380 B.n606 B.n605 585
R381 B.n607 B.n606 585
R382 B.n311 B.n310 585
R383 B.n312 B.n311 585
R384 B.n615 B.n614 585
R385 B.n614 B.n613 585
R386 B.n616 B.n309 585
R387 B.n309 B.n308 585
R388 B.n618 B.n617 585
R389 B.n619 B.n618 585
R390 B.n303 B.n302 585
R391 B.n304 B.n303 585
R392 B.n627 B.n626 585
R393 B.n626 B.n625 585
R394 B.n628 B.n301 585
R395 B.n301 B.n300 585
R396 B.n630 B.n629 585
R397 B.n631 B.n630 585
R398 B.n295 B.n294 585
R399 B.n296 B.n295 585
R400 B.n639 B.n638 585
R401 B.n638 B.n637 585
R402 B.n640 B.n293 585
R403 B.n293 B.n292 585
R404 B.n642 B.n641 585
R405 B.n643 B.n642 585
R406 B.n287 B.n286 585
R407 B.n288 B.n287 585
R408 B.n651 B.n650 585
R409 B.n650 B.n649 585
R410 B.n652 B.n285 585
R411 B.n285 B.n284 585
R412 B.n654 B.n653 585
R413 B.n655 B.n654 585
R414 B.n279 B.n278 585
R415 B.n280 B.n279 585
R416 B.n663 B.n662 585
R417 B.n662 B.n661 585
R418 B.n664 B.n277 585
R419 B.n277 B.n276 585
R420 B.n666 B.n665 585
R421 B.n667 B.n666 585
R422 B.n271 B.n270 585
R423 B.n272 B.n271 585
R424 B.n676 B.n675 585
R425 B.n675 B.n674 585
R426 B.n677 B.n269 585
R427 B.n269 B.n268 585
R428 B.n679 B.n678 585
R429 B.n680 B.n679 585
R430 B.n2 B.n0 585
R431 B.n4 B.n2 585
R432 B.n3 B.n1 585
R433 B.n844 B.n3 585
R434 B.n842 B.n841 585
R435 B.n843 B.n842 585
R436 B.n840 B.n9 585
R437 B.n9 B.n8 585
R438 B.n839 B.n838 585
R439 B.n838 B.n837 585
R440 B.n11 B.n10 585
R441 B.n836 B.n11 585
R442 B.n834 B.n833 585
R443 B.n835 B.n834 585
R444 B.n832 B.n16 585
R445 B.n16 B.n15 585
R446 B.n831 B.n830 585
R447 B.n830 B.n829 585
R448 B.n18 B.n17 585
R449 B.n828 B.n18 585
R450 B.n826 B.n825 585
R451 B.n827 B.n826 585
R452 B.n824 B.n23 585
R453 B.n23 B.n22 585
R454 B.n823 B.n822 585
R455 B.n822 B.n821 585
R456 B.n25 B.n24 585
R457 B.n820 B.n25 585
R458 B.n818 B.n817 585
R459 B.n819 B.n818 585
R460 B.n816 B.n30 585
R461 B.n30 B.n29 585
R462 B.n815 B.n814 585
R463 B.n814 B.n813 585
R464 B.n32 B.n31 585
R465 B.n812 B.n32 585
R466 B.n810 B.n809 585
R467 B.n811 B.n810 585
R468 B.n808 B.n37 585
R469 B.n37 B.n36 585
R470 B.n807 B.n806 585
R471 B.n806 B.n805 585
R472 B.n39 B.n38 585
R473 B.n804 B.n39 585
R474 B.n802 B.n801 585
R475 B.n803 B.n802 585
R476 B.n800 B.n44 585
R477 B.n44 B.n43 585
R478 B.n799 B.n798 585
R479 B.n798 B.n797 585
R480 B.n46 B.n45 585
R481 B.n796 B.n46 585
R482 B.n794 B.n793 585
R483 B.n795 B.n794 585
R484 B.n792 B.n51 585
R485 B.n51 B.n50 585
R486 B.n791 B.n790 585
R487 B.n790 B.n789 585
R488 B.n53 B.n52 585
R489 B.n788 B.n53 585
R490 B.n786 B.n785 585
R491 B.n787 B.n786 585
R492 B.n784 B.n58 585
R493 B.n58 B.n57 585
R494 B.n783 B.n782 585
R495 B.n782 B.n781 585
R496 B.n60 B.n59 585
R497 B.n780 B.n60 585
R498 B.n778 B.n777 585
R499 B.n779 B.n778 585
R500 B.n776 B.n65 585
R501 B.n65 B.n64 585
R502 B.n775 B.n774 585
R503 B.n774 B.n773 585
R504 B.n67 B.n66 585
R505 B.n772 B.n67 585
R506 B.n770 B.n769 585
R507 B.n771 B.n770 585
R508 B.n768 B.n72 585
R509 B.n72 B.n71 585
R510 B.n767 B.n766 585
R511 B.n766 B.n765 585
R512 B.n74 B.n73 585
R513 B.n764 B.n74 585
R514 B.n762 B.n761 585
R515 B.n763 B.n762 585
R516 B.n760 B.n79 585
R517 B.n79 B.n78 585
R518 B.n759 B.n758 585
R519 B.n758 B.n757 585
R520 B.n81 B.n80 585
R521 B.n756 B.n81 585
R522 B.n754 B.n753 585
R523 B.n755 B.n754 585
R524 B.n752 B.n86 585
R525 B.n86 B.n85 585
R526 B.n751 B.n750 585
R527 B.n750 B.n749 585
R528 B.n847 B.n846 585
R529 B.n846 B.n845 585
R530 B.n542 B.n359 497.305
R531 B.n750 B.n88 497.305
R532 B.n540 B.n361 497.305
R533 B.n746 B.n89 497.305
R534 B.n377 B.t19 290.014
R535 B.n454 B.t8 290.014
R536 B.n128 B.t12 290.014
R537 B.n125 B.t16 290.014
R538 B.n377 B.t21 268.37
R539 B.n125 B.t17 268.37
R540 B.n454 B.t11 268.37
R541 B.n128 B.t14 268.37
R542 B.n748 B.n747 256.663
R543 B.n748 B.n123 256.663
R544 B.n748 B.n122 256.663
R545 B.n748 B.n121 256.663
R546 B.n748 B.n120 256.663
R547 B.n748 B.n119 256.663
R548 B.n748 B.n118 256.663
R549 B.n748 B.n117 256.663
R550 B.n748 B.n116 256.663
R551 B.n748 B.n115 256.663
R552 B.n748 B.n114 256.663
R553 B.n748 B.n113 256.663
R554 B.n748 B.n112 256.663
R555 B.n748 B.n111 256.663
R556 B.n748 B.n110 256.663
R557 B.n748 B.n109 256.663
R558 B.n748 B.n108 256.663
R559 B.n748 B.n107 256.663
R560 B.n748 B.n106 256.663
R561 B.n748 B.n105 256.663
R562 B.n748 B.n104 256.663
R563 B.n748 B.n103 256.663
R564 B.n748 B.n102 256.663
R565 B.n748 B.n101 256.663
R566 B.n748 B.n100 256.663
R567 B.n748 B.n99 256.663
R568 B.n748 B.n98 256.663
R569 B.n748 B.n97 256.663
R570 B.n748 B.n96 256.663
R571 B.n748 B.n95 256.663
R572 B.n748 B.n94 256.663
R573 B.n748 B.n93 256.663
R574 B.n748 B.n92 256.663
R575 B.n748 B.n91 256.663
R576 B.n748 B.n90 256.663
R577 B.n399 B.n360 256.663
R578 B.n402 B.n360 256.663
R579 B.n408 B.n360 256.663
R580 B.n410 B.n360 256.663
R581 B.n416 B.n360 256.663
R582 B.n418 B.n360 256.663
R583 B.n424 B.n360 256.663
R584 B.n426 B.n360 256.663
R585 B.n432 B.n360 256.663
R586 B.n434 B.n360 256.663
R587 B.n440 B.n360 256.663
R588 B.n442 B.n360 256.663
R589 B.n448 B.n360 256.663
R590 B.n450 B.n360 256.663
R591 B.n459 B.n360 256.663
R592 B.n461 B.n360 256.663
R593 B.n467 B.n360 256.663
R594 B.n469 B.n360 256.663
R595 B.n475 B.n360 256.663
R596 B.n477 B.n360 256.663
R597 B.n484 B.n360 256.663
R598 B.n486 B.n360 256.663
R599 B.n492 B.n360 256.663
R600 B.n494 B.n360 256.663
R601 B.n500 B.n360 256.663
R602 B.n502 B.n360 256.663
R603 B.n508 B.n360 256.663
R604 B.n510 B.n360 256.663
R605 B.n516 B.n360 256.663
R606 B.n518 B.n360 256.663
R607 B.n524 B.n360 256.663
R608 B.n526 B.n360 256.663
R609 B.n532 B.n360 256.663
R610 B.n535 B.n360 256.663
R611 B.n378 B.t20 215.812
R612 B.n126 B.t18 215.812
R613 B.n455 B.t10 215.812
R614 B.n129 B.t15 215.812
R615 B.n542 B.n357 163.367
R616 B.n546 B.n357 163.367
R617 B.n546 B.n351 163.367
R618 B.n554 B.n351 163.367
R619 B.n554 B.n349 163.367
R620 B.n558 B.n349 163.367
R621 B.n558 B.n343 163.367
R622 B.n566 B.n343 163.367
R623 B.n566 B.n341 163.367
R624 B.n570 B.n341 163.367
R625 B.n570 B.n335 163.367
R626 B.n578 B.n335 163.367
R627 B.n578 B.n333 163.367
R628 B.n582 B.n333 163.367
R629 B.n582 B.n327 163.367
R630 B.n590 B.n327 163.367
R631 B.n590 B.n325 163.367
R632 B.n594 B.n325 163.367
R633 B.n594 B.n319 163.367
R634 B.n602 B.n319 163.367
R635 B.n602 B.n317 163.367
R636 B.n606 B.n317 163.367
R637 B.n606 B.n311 163.367
R638 B.n614 B.n311 163.367
R639 B.n614 B.n309 163.367
R640 B.n618 B.n309 163.367
R641 B.n618 B.n303 163.367
R642 B.n626 B.n303 163.367
R643 B.n626 B.n301 163.367
R644 B.n630 B.n301 163.367
R645 B.n630 B.n295 163.367
R646 B.n638 B.n295 163.367
R647 B.n638 B.n293 163.367
R648 B.n642 B.n293 163.367
R649 B.n642 B.n287 163.367
R650 B.n650 B.n287 163.367
R651 B.n650 B.n285 163.367
R652 B.n654 B.n285 163.367
R653 B.n654 B.n279 163.367
R654 B.n662 B.n279 163.367
R655 B.n662 B.n277 163.367
R656 B.n666 B.n277 163.367
R657 B.n666 B.n271 163.367
R658 B.n675 B.n271 163.367
R659 B.n675 B.n269 163.367
R660 B.n679 B.n269 163.367
R661 B.n679 B.n2 163.367
R662 B.n846 B.n2 163.367
R663 B.n846 B.n3 163.367
R664 B.n842 B.n3 163.367
R665 B.n842 B.n9 163.367
R666 B.n838 B.n9 163.367
R667 B.n838 B.n11 163.367
R668 B.n834 B.n11 163.367
R669 B.n834 B.n16 163.367
R670 B.n830 B.n16 163.367
R671 B.n830 B.n18 163.367
R672 B.n826 B.n18 163.367
R673 B.n826 B.n23 163.367
R674 B.n822 B.n23 163.367
R675 B.n822 B.n25 163.367
R676 B.n818 B.n25 163.367
R677 B.n818 B.n30 163.367
R678 B.n814 B.n30 163.367
R679 B.n814 B.n32 163.367
R680 B.n810 B.n32 163.367
R681 B.n810 B.n37 163.367
R682 B.n806 B.n37 163.367
R683 B.n806 B.n39 163.367
R684 B.n802 B.n39 163.367
R685 B.n802 B.n44 163.367
R686 B.n798 B.n44 163.367
R687 B.n798 B.n46 163.367
R688 B.n794 B.n46 163.367
R689 B.n794 B.n51 163.367
R690 B.n790 B.n51 163.367
R691 B.n790 B.n53 163.367
R692 B.n786 B.n53 163.367
R693 B.n786 B.n58 163.367
R694 B.n782 B.n58 163.367
R695 B.n782 B.n60 163.367
R696 B.n778 B.n60 163.367
R697 B.n778 B.n65 163.367
R698 B.n774 B.n65 163.367
R699 B.n774 B.n67 163.367
R700 B.n770 B.n67 163.367
R701 B.n770 B.n72 163.367
R702 B.n766 B.n72 163.367
R703 B.n766 B.n74 163.367
R704 B.n762 B.n74 163.367
R705 B.n762 B.n79 163.367
R706 B.n758 B.n79 163.367
R707 B.n758 B.n81 163.367
R708 B.n754 B.n81 163.367
R709 B.n754 B.n86 163.367
R710 B.n750 B.n86 163.367
R711 B.n401 B.n400 163.367
R712 B.n403 B.n401 163.367
R713 B.n407 B.n396 163.367
R714 B.n411 B.n409 163.367
R715 B.n415 B.n394 163.367
R716 B.n419 B.n417 163.367
R717 B.n423 B.n392 163.367
R718 B.n427 B.n425 163.367
R719 B.n431 B.n390 163.367
R720 B.n435 B.n433 163.367
R721 B.n439 B.n388 163.367
R722 B.n443 B.n441 163.367
R723 B.n447 B.n386 163.367
R724 B.n451 B.n449 163.367
R725 B.n458 B.n384 163.367
R726 B.n462 B.n460 163.367
R727 B.n466 B.n382 163.367
R728 B.n470 B.n468 163.367
R729 B.n474 B.n380 163.367
R730 B.n478 B.n476 163.367
R731 B.n483 B.n376 163.367
R732 B.n487 B.n485 163.367
R733 B.n491 B.n374 163.367
R734 B.n495 B.n493 163.367
R735 B.n499 B.n372 163.367
R736 B.n503 B.n501 163.367
R737 B.n507 B.n370 163.367
R738 B.n511 B.n509 163.367
R739 B.n515 B.n368 163.367
R740 B.n519 B.n517 163.367
R741 B.n523 B.n366 163.367
R742 B.n527 B.n525 163.367
R743 B.n531 B.n364 163.367
R744 B.n534 B.n533 163.367
R745 B.n536 B.n361 163.367
R746 B.n540 B.n355 163.367
R747 B.n548 B.n355 163.367
R748 B.n548 B.n353 163.367
R749 B.n552 B.n353 163.367
R750 B.n552 B.n346 163.367
R751 B.n560 B.n346 163.367
R752 B.n560 B.n344 163.367
R753 B.n564 B.n344 163.367
R754 B.n564 B.n339 163.367
R755 B.n572 B.n339 163.367
R756 B.n572 B.n337 163.367
R757 B.n576 B.n337 163.367
R758 B.n576 B.n331 163.367
R759 B.n584 B.n331 163.367
R760 B.n584 B.n329 163.367
R761 B.n588 B.n329 163.367
R762 B.n588 B.n323 163.367
R763 B.n596 B.n323 163.367
R764 B.n596 B.n321 163.367
R765 B.n600 B.n321 163.367
R766 B.n600 B.n315 163.367
R767 B.n608 B.n315 163.367
R768 B.n608 B.n313 163.367
R769 B.n612 B.n313 163.367
R770 B.n612 B.n307 163.367
R771 B.n620 B.n307 163.367
R772 B.n620 B.n305 163.367
R773 B.n624 B.n305 163.367
R774 B.n624 B.n299 163.367
R775 B.n632 B.n299 163.367
R776 B.n632 B.n297 163.367
R777 B.n636 B.n297 163.367
R778 B.n636 B.n291 163.367
R779 B.n644 B.n291 163.367
R780 B.n644 B.n289 163.367
R781 B.n648 B.n289 163.367
R782 B.n648 B.n283 163.367
R783 B.n656 B.n283 163.367
R784 B.n656 B.n281 163.367
R785 B.n660 B.n281 163.367
R786 B.n660 B.n275 163.367
R787 B.n668 B.n275 163.367
R788 B.n668 B.n273 163.367
R789 B.n673 B.n273 163.367
R790 B.n673 B.n267 163.367
R791 B.n681 B.n267 163.367
R792 B.n682 B.n681 163.367
R793 B.n682 B.n5 163.367
R794 B.n6 B.n5 163.367
R795 B.n7 B.n6 163.367
R796 B.n687 B.n7 163.367
R797 B.n687 B.n12 163.367
R798 B.n13 B.n12 163.367
R799 B.n14 B.n13 163.367
R800 B.n692 B.n14 163.367
R801 B.n692 B.n19 163.367
R802 B.n20 B.n19 163.367
R803 B.n21 B.n20 163.367
R804 B.n697 B.n21 163.367
R805 B.n697 B.n26 163.367
R806 B.n27 B.n26 163.367
R807 B.n28 B.n27 163.367
R808 B.n702 B.n28 163.367
R809 B.n702 B.n33 163.367
R810 B.n34 B.n33 163.367
R811 B.n35 B.n34 163.367
R812 B.n707 B.n35 163.367
R813 B.n707 B.n40 163.367
R814 B.n41 B.n40 163.367
R815 B.n42 B.n41 163.367
R816 B.n712 B.n42 163.367
R817 B.n712 B.n47 163.367
R818 B.n48 B.n47 163.367
R819 B.n49 B.n48 163.367
R820 B.n717 B.n49 163.367
R821 B.n717 B.n54 163.367
R822 B.n55 B.n54 163.367
R823 B.n56 B.n55 163.367
R824 B.n722 B.n56 163.367
R825 B.n722 B.n61 163.367
R826 B.n62 B.n61 163.367
R827 B.n63 B.n62 163.367
R828 B.n727 B.n63 163.367
R829 B.n727 B.n68 163.367
R830 B.n69 B.n68 163.367
R831 B.n70 B.n69 163.367
R832 B.n732 B.n70 163.367
R833 B.n732 B.n75 163.367
R834 B.n76 B.n75 163.367
R835 B.n77 B.n76 163.367
R836 B.n737 B.n77 163.367
R837 B.n737 B.n82 163.367
R838 B.n83 B.n82 163.367
R839 B.n84 B.n83 163.367
R840 B.n742 B.n84 163.367
R841 B.n742 B.n89 163.367
R842 B.n133 B.n132 163.367
R843 B.n137 B.n136 163.367
R844 B.n141 B.n140 163.367
R845 B.n145 B.n144 163.367
R846 B.n149 B.n148 163.367
R847 B.n153 B.n152 163.367
R848 B.n157 B.n156 163.367
R849 B.n161 B.n160 163.367
R850 B.n165 B.n164 163.367
R851 B.n169 B.n168 163.367
R852 B.n173 B.n172 163.367
R853 B.n177 B.n176 163.367
R854 B.n181 B.n180 163.367
R855 B.n185 B.n184 163.367
R856 B.n189 B.n188 163.367
R857 B.n193 B.n192 163.367
R858 B.n197 B.n196 163.367
R859 B.n201 B.n200 163.367
R860 B.n205 B.n204 163.367
R861 B.n209 B.n208 163.367
R862 B.n213 B.n212 163.367
R863 B.n217 B.n216 163.367
R864 B.n221 B.n220 163.367
R865 B.n225 B.n224 163.367
R866 B.n229 B.n228 163.367
R867 B.n233 B.n232 163.367
R868 B.n237 B.n236 163.367
R869 B.n241 B.n240 163.367
R870 B.n245 B.n244 163.367
R871 B.n249 B.n248 163.367
R872 B.n253 B.n252 163.367
R873 B.n257 B.n256 163.367
R874 B.n261 B.n260 163.367
R875 B.n263 B.n124 163.367
R876 B.n541 B.n360 99.2918
R877 B.n749 B.n748 99.2918
R878 B.n399 B.n359 71.676
R879 B.n403 B.n402 71.676
R880 B.n408 B.n407 71.676
R881 B.n411 B.n410 71.676
R882 B.n416 B.n415 71.676
R883 B.n419 B.n418 71.676
R884 B.n424 B.n423 71.676
R885 B.n427 B.n426 71.676
R886 B.n432 B.n431 71.676
R887 B.n435 B.n434 71.676
R888 B.n440 B.n439 71.676
R889 B.n443 B.n442 71.676
R890 B.n448 B.n447 71.676
R891 B.n451 B.n450 71.676
R892 B.n459 B.n458 71.676
R893 B.n462 B.n461 71.676
R894 B.n467 B.n466 71.676
R895 B.n470 B.n469 71.676
R896 B.n475 B.n474 71.676
R897 B.n478 B.n477 71.676
R898 B.n484 B.n483 71.676
R899 B.n487 B.n486 71.676
R900 B.n492 B.n491 71.676
R901 B.n495 B.n494 71.676
R902 B.n500 B.n499 71.676
R903 B.n503 B.n502 71.676
R904 B.n508 B.n507 71.676
R905 B.n511 B.n510 71.676
R906 B.n516 B.n515 71.676
R907 B.n519 B.n518 71.676
R908 B.n524 B.n523 71.676
R909 B.n527 B.n526 71.676
R910 B.n532 B.n531 71.676
R911 B.n535 B.n534 71.676
R912 B.n90 B.n88 71.676
R913 B.n133 B.n91 71.676
R914 B.n137 B.n92 71.676
R915 B.n141 B.n93 71.676
R916 B.n145 B.n94 71.676
R917 B.n149 B.n95 71.676
R918 B.n153 B.n96 71.676
R919 B.n157 B.n97 71.676
R920 B.n161 B.n98 71.676
R921 B.n165 B.n99 71.676
R922 B.n169 B.n100 71.676
R923 B.n173 B.n101 71.676
R924 B.n177 B.n102 71.676
R925 B.n181 B.n103 71.676
R926 B.n185 B.n104 71.676
R927 B.n189 B.n105 71.676
R928 B.n193 B.n106 71.676
R929 B.n197 B.n107 71.676
R930 B.n201 B.n108 71.676
R931 B.n205 B.n109 71.676
R932 B.n209 B.n110 71.676
R933 B.n213 B.n111 71.676
R934 B.n217 B.n112 71.676
R935 B.n221 B.n113 71.676
R936 B.n225 B.n114 71.676
R937 B.n229 B.n115 71.676
R938 B.n233 B.n116 71.676
R939 B.n237 B.n117 71.676
R940 B.n241 B.n118 71.676
R941 B.n245 B.n119 71.676
R942 B.n249 B.n120 71.676
R943 B.n253 B.n121 71.676
R944 B.n257 B.n122 71.676
R945 B.n261 B.n123 71.676
R946 B.n747 B.n124 71.676
R947 B.n747 B.n746 71.676
R948 B.n263 B.n123 71.676
R949 B.n260 B.n122 71.676
R950 B.n256 B.n121 71.676
R951 B.n252 B.n120 71.676
R952 B.n248 B.n119 71.676
R953 B.n244 B.n118 71.676
R954 B.n240 B.n117 71.676
R955 B.n236 B.n116 71.676
R956 B.n232 B.n115 71.676
R957 B.n228 B.n114 71.676
R958 B.n224 B.n113 71.676
R959 B.n220 B.n112 71.676
R960 B.n216 B.n111 71.676
R961 B.n212 B.n110 71.676
R962 B.n208 B.n109 71.676
R963 B.n204 B.n108 71.676
R964 B.n200 B.n107 71.676
R965 B.n196 B.n106 71.676
R966 B.n192 B.n105 71.676
R967 B.n188 B.n104 71.676
R968 B.n184 B.n103 71.676
R969 B.n180 B.n102 71.676
R970 B.n176 B.n101 71.676
R971 B.n172 B.n100 71.676
R972 B.n168 B.n99 71.676
R973 B.n164 B.n98 71.676
R974 B.n160 B.n97 71.676
R975 B.n156 B.n96 71.676
R976 B.n152 B.n95 71.676
R977 B.n148 B.n94 71.676
R978 B.n144 B.n93 71.676
R979 B.n140 B.n92 71.676
R980 B.n136 B.n91 71.676
R981 B.n132 B.n90 71.676
R982 B.n400 B.n399 71.676
R983 B.n402 B.n396 71.676
R984 B.n409 B.n408 71.676
R985 B.n410 B.n394 71.676
R986 B.n417 B.n416 71.676
R987 B.n418 B.n392 71.676
R988 B.n425 B.n424 71.676
R989 B.n426 B.n390 71.676
R990 B.n433 B.n432 71.676
R991 B.n434 B.n388 71.676
R992 B.n441 B.n440 71.676
R993 B.n442 B.n386 71.676
R994 B.n449 B.n448 71.676
R995 B.n450 B.n384 71.676
R996 B.n460 B.n459 71.676
R997 B.n461 B.n382 71.676
R998 B.n468 B.n467 71.676
R999 B.n469 B.n380 71.676
R1000 B.n476 B.n475 71.676
R1001 B.n477 B.n376 71.676
R1002 B.n485 B.n484 71.676
R1003 B.n486 B.n374 71.676
R1004 B.n493 B.n492 71.676
R1005 B.n494 B.n372 71.676
R1006 B.n501 B.n500 71.676
R1007 B.n502 B.n370 71.676
R1008 B.n509 B.n508 71.676
R1009 B.n510 B.n368 71.676
R1010 B.n517 B.n516 71.676
R1011 B.n518 B.n366 71.676
R1012 B.n525 B.n524 71.676
R1013 B.n526 B.n364 71.676
R1014 B.n533 B.n532 71.676
R1015 B.n536 B.n535 71.676
R1016 B.n480 B.n378 59.5399
R1017 B.n456 B.n455 59.5399
R1018 B.n130 B.n129 59.5399
R1019 B.n127 B.n126 59.5399
R1020 B.n541 B.n356 55.8006
R1021 B.n547 B.n356 55.8006
R1022 B.n547 B.n352 55.8006
R1023 B.n553 B.n352 55.8006
R1024 B.n553 B.n347 55.8006
R1025 B.n559 B.n347 55.8006
R1026 B.n559 B.n348 55.8006
R1027 B.n565 B.n340 55.8006
R1028 B.n571 B.n340 55.8006
R1029 B.n571 B.n336 55.8006
R1030 B.n577 B.n336 55.8006
R1031 B.n577 B.n332 55.8006
R1032 B.n583 B.n332 55.8006
R1033 B.n583 B.n328 55.8006
R1034 B.n589 B.n328 55.8006
R1035 B.n589 B.n324 55.8006
R1036 B.n595 B.n324 55.8006
R1037 B.n601 B.n320 55.8006
R1038 B.n601 B.n316 55.8006
R1039 B.n607 B.n316 55.8006
R1040 B.n607 B.n312 55.8006
R1041 B.n613 B.n312 55.8006
R1042 B.n613 B.n308 55.8006
R1043 B.n619 B.n308 55.8006
R1044 B.n625 B.n304 55.8006
R1045 B.n625 B.n300 55.8006
R1046 B.n631 B.n300 55.8006
R1047 B.n631 B.n296 55.8006
R1048 B.n637 B.n296 55.8006
R1049 B.n637 B.n292 55.8006
R1050 B.n643 B.n292 55.8006
R1051 B.n649 B.n288 55.8006
R1052 B.n649 B.n284 55.8006
R1053 B.n655 B.n284 55.8006
R1054 B.n655 B.n280 55.8006
R1055 B.n661 B.n280 55.8006
R1056 B.n661 B.n276 55.8006
R1057 B.n667 B.n276 55.8006
R1058 B.n674 B.n272 55.8006
R1059 B.n674 B.n268 55.8006
R1060 B.n680 B.n268 55.8006
R1061 B.n680 B.n4 55.8006
R1062 B.n845 B.n4 55.8006
R1063 B.n845 B.n844 55.8006
R1064 B.n844 B.n843 55.8006
R1065 B.n843 B.n8 55.8006
R1066 B.n837 B.n8 55.8006
R1067 B.n837 B.n836 55.8006
R1068 B.n835 B.n15 55.8006
R1069 B.n829 B.n15 55.8006
R1070 B.n829 B.n828 55.8006
R1071 B.n828 B.n827 55.8006
R1072 B.n827 B.n22 55.8006
R1073 B.n821 B.n22 55.8006
R1074 B.n821 B.n820 55.8006
R1075 B.n819 B.n29 55.8006
R1076 B.n813 B.n29 55.8006
R1077 B.n813 B.n812 55.8006
R1078 B.n812 B.n811 55.8006
R1079 B.n811 B.n36 55.8006
R1080 B.n805 B.n36 55.8006
R1081 B.n805 B.n804 55.8006
R1082 B.n803 B.n43 55.8006
R1083 B.n797 B.n43 55.8006
R1084 B.n797 B.n796 55.8006
R1085 B.n796 B.n795 55.8006
R1086 B.n795 B.n50 55.8006
R1087 B.n789 B.n50 55.8006
R1088 B.n789 B.n788 55.8006
R1089 B.n787 B.n57 55.8006
R1090 B.n781 B.n57 55.8006
R1091 B.n781 B.n780 55.8006
R1092 B.n780 B.n779 55.8006
R1093 B.n779 B.n64 55.8006
R1094 B.n773 B.n64 55.8006
R1095 B.n773 B.n772 55.8006
R1096 B.n772 B.n771 55.8006
R1097 B.n771 B.n71 55.8006
R1098 B.n765 B.n71 55.8006
R1099 B.n764 B.n763 55.8006
R1100 B.n763 B.n78 55.8006
R1101 B.n757 B.n78 55.8006
R1102 B.n757 B.n756 55.8006
R1103 B.n756 B.n755 55.8006
R1104 B.n755 B.n85 55.8006
R1105 B.n749 B.n85 55.8006
R1106 B.n378 B.n377 52.5581
R1107 B.n455 B.n454 52.5581
R1108 B.n129 B.n128 52.5581
R1109 B.n126 B.n125 52.5581
R1110 B.n565 B.t9 37.7476
R1111 B.n765 B.t13 37.7476
R1112 B.t6 B.n272 32.8241
R1113 B.n836 B.t1 32.8241
R1114 B.n751 B.n87 32.3127
R1115 B.n745 B.n744 32.3127
R1116 B.n539 B.n538 32.3127
R1117 B.n543 B.n358 32.3127
R1118 B.t4 B.n288 31.1829
R1119 B.n820 B.t0 31.1829
R1120 B.t2 B.n304 29.5417
R1121 B.n804 B.t3 29.5417
R1122 B.n595 B.t5 27.9005
R1123 B.t5 B.n320 27.9005
R1124 B.n788 B.t7 27.9005
R1125 B.t7 B.n787 27.9005
R1126 B.n619 B.t2 26.2594
R1127 B.t3 B.n803 26.2594
R1128 B.n643 B.t4 24.6182
R1129 B.t0 B.n819 24.6182
R1130 B.n667 B.t6 22.977
R1131 B.t1 B.n835 22.977
R1132 B.n348 B.t9 18.0535
R1133 B.t13 B.n764 18.0535
R1134 B B.n847 18.0485
R1135 B.n131 B.n87 10.6151
R1136 B.n134 B.n131 10.6151
R1137 B.n135 B.n134 10.6151
R1138 B.n138 B.n135 10.6151
R1139 B.n139 B.n138 10.6151
R1140 B.n142 B.n139 10.6151
R1141 B.n143 B.n142 10.6151
R1142 B.n146 B.n143 10.6151
R1143 B.n147 B.n146 10.6151
R1144 B.n150 B.n147 10.6151
R1145 B.n151 B.n150 10.6151
R1146 B.n154 B.n151 10.6151
R1147 B.n155 B.n154 10.6151
R1148 B.n158 B.n155 10.6151
R1149 B.n159 B.n158 10.6151
R1150 B.n162 B.n159 10.6151
R1151 B.n163 B.n162 10.6151
R1152 B.n166 B.n163 10.6151
R1153 B.n167 B.n166 10.6151
R1154 B.n170 B.n167 10.6151
R1155 B.n171 B.n170 10.6151
R1156 B.n174 B.n171 10.6151
R1157 B.n175 B.n174 10.6151
R1158 B.n178 B.n175 10.6151
R1159 B.n179 B.n178 10.6151
R1160 B.n182 B.n179 10.6151
R1161 B.n183 B.n182 10.6151
R1162 B.n186 B.n183 10.6151
R1163 B.n187 B.n186 10.6151
R1164 B.n191 B.n190 10.6151
R1165 B.n194 B.n191 10.6151
R1166 B.n195 B.n194 10.6151
R1167 B.n198 B.n195 10.6151
R1168 B.n199 B.n198 10.6151
R1169 B.n202 B.n199 10.6151
R1170 B.n203 B.n202 10.6151
R1171 B.n206 B.n203 10.6151
R1172 B.n207 B.n206 10.6151
R1173 B.n211 B.n210 10.6151
R1174 B.n214 B.n211 10.6151
R1175 B.n215 B.n214 10.6151
R1176 B.n218 B.n215 10.6151
R1177 B.n219 B.n218 10.6151
R1178 B.n222 B.n219 10.6151
R1179 B.n223 B.n222 10.6151
R1180 B.n226 B.n223 10.6151
R1181 B.n227 B.n226 10.6151
R1182 B.n230 B.n227 10.6151
R1183 B.n231 B.n230 10.6151
R1184 B.n234 B.n231 10.6151
R1185 B.n235 B.n234 10.6151
R1186 B.n238 B.n235 10.6151
R1187 B.n239 B.n238 10.6151
R1188 B.n242 B.n239 10.6151
R1189 B.n243 B.n242 10.6151
R1190 B.n246 B.n243 10.6151
R1191 B.n247 B.n246 10.6151
R1192 B.n250 B.n247 10.6151
R1193 B.n251 B.n250 10.6151
R1194 B.n254 B.n251 10.6151
R1195 B.n255 B.n254 10.6151
R1196 B.n258 B.n255 10.6151
R1197 B.n259 B.n258 10.6151
R1198 B.n262 B.n259 10.6151
R1199 B.n264 B.n262 10.6151
R1200 B.n265 B.n264 10.6151
R1201 B.n745 B.n265 10.6151
R1202 B.n539 B.n354 10.6151
R1203 B.n549 B.n354 10.6151
R1204 B.n550 B.n549 10.6151
R1205 B.n551 B.n550 10.6151
R1206 B.n551 B.n345 10.6151
R1207 B.n561 B.n345 10.6151
R1208 B.n562 B.n561 10.6151
R1209 B.n563 B.n562 10.6151
R1210 B.n563 B.n338 10.6151
R1211 B.n573 B.n338 10.6151
R1212 B.n574 B.n573 10.6151
R1213 B.n575 B.n574 10.6151
R1214 B.n575 B.n330 10.6151
R1215 B.n585 B.n330 10.6151
R1216 B.n586 B.n585 10.6151
R1217 B.n587 B.n586 10.6151
R1218 B.n587 B.n322 10.6151
R1219 B.n597 B.n322 10.6151
R1220 B.n598 B.n597 10.6151
R1221 B.n599 B.n598 10.6151
R1222 B.n599 B.n314 10.6151
R1223 B.n609 B.n314 10.6151
R1224 B.n610 B.n609 10.6151
R1225 B.n611 B.n610 10.6151
R1226 B.n611 B.n306 10.6151
R1227 B.n621 B.n306 10.6151
R1228 B.n622 B.n621 10.6151
R1229 B.n623 B.n622 10.6151
R1230 B.n623 B.n298 10.6151
R1231 B.n633 B.n298 10.6151
R1232 B.n634 B.n633 10.6151
R1233 B.n635 B.n634 10.6151
R1234 B.n635 B.n290 10.6151
R1235 B.n645 B.n290 10.6151
R1236 B.n646 B.n645 10.6151
R1237 B.n647 B.n646 10.6151
R1238 B.n647 B.n282 10.6151
R1239 B.n657 B.n282 10.6151
R1240 B.n658 B.n657 10.6151
R1241 B.n659 B.n658 10.6151
R1242 B.n659 B.n274 10.6151
R1243 B.n669 B.n274 10.6151
R1244 B.n670 B.n669 10.6151
R1245 B.n672 B.n670 10.6151
R1246 B.n672 B.n671 10.6151
R1247 B.n671 B.n266 10.6151
R1248 B.n683 B.n266 10.6151
R1249 B.n684 B.n683 10.6151
R1250 B.n685 B.n684 10.6151
R1251 B.n686 B.n685 10.6151
R1252 B.n688 B.n686 10.6151
R1253 B.n689 B.n688 10.6151
R1254 B.n690 B.n689 10.6151
R1255 B.n691 B.n690 10.6151
R1256 B.n693 B.n691 10.6151
R1257 B.n694 B.n693 10.6151
R1258 B.n695 B.n694 10.6151
R1259 B.n696 B.n695 10.6151
R1260 B.n698 B.n696 10.6151
R1261 B.n699 B.n698 10.6151
R1262 B.n700 B.n699 10.6151
R1263 B.n701 B.n700 10.6151
R1264 B.n703 B.n701 10.6151
R1265 B.n704 B.n703 10.6151
R1266 B.n705 B.n704 10.6151
R1267 B.n706 B.n705 10.6151
R1268 B.n708 B.n706 10.6151
R1269 B.n709 B.n708 10.6151
R1270 B.n710 B.n709 10.6151
R1271 B.n711 B.n710 10.6151
R1272 B.n713 B.n711 10.6151
R1273 B.n714 B.n713 10.6151
R1274 B.n715 B.n714 10.6151
R1275 B.n716 B.n715 10.6151
R1276 B.n718 B.n716 10.6151
R1277 B.n719 B.n718 10.6151
R1278 B.n720 B.n719 10.6151
R1279 B.n721 B.n720 10.6151
R1280 B.n723 B.n721 10.6151
R1281 B.n724 B.n723 10.6151
R1282 B.n725 B.n724 10.6151
R1283 B.n726 B.n725 10.6151
R1284 B.n728 B.n726 10.6151
R1285 B.n729 B.n728 10.6151
R1286 B.n730 B.n729 10.6151
R1287 B.n731 B.n730 10.6151
R1288 B.n733 B.n731 10.6151
R1289 B.n734 B.n733 10.6151
R1290 B.n735 B.n734 10.6151
R1291 B.n736 B.n735 10.6151
R1292 B.n738 B.n736 10.6151
R1293 B.n739 B.n738 10.6151
R1294 B.n740 B.n739 10.6151
R1295 B.n741 B.n740 10.6151
R1296 B.n743 B.n741 10.6151
R1297 B.n744 B.n743 10.6151
R1298 B.n398 B.n358 10.6151
R1299 B.n398 B.n397 10.6151
R1300 B.n404 B.n397 10.6151
R1301 B.n405 B.n404 10.6151
R1302 B.n406 B.n405 10.6151
R1303 B.n406 B.n395 10.6151
R1304 B.n412 B.n395 10.6151
R1305 B.n413 B.n412 10.6151
R1306 B.n414 B.n413 10.6151
R1307 B.n414 B.n393 10.6151
R1308 B.n420 B.n393 10.6151
R1309 B.n421 B.n420 10.6151
R1310 B.n422 B.n421 10.6151
R1311 B.n422 B.n391 10.6151
R1312 B.n428 B.n391 10.6151
R1313 B.n429 B.n428 10.6151
R1314 B.n430 B.n429 10.6151
R1315 B.n430 B.n389 10.6151
R1316 B.n436 B.n389 10.6151
R1317 B.n437 B.n436 10.6151
R1318 B.n438 B.n437 10.6151
R1319 B.n438 B.n387 10.6151
R1320 B.n444 B.n387 10.6151
R1321 B.n445 B.n444 10.6151
R1322 B.n446 B.n445 10.6151
R1323 B.n446 B.n385 10.6151
R1324 B.n452 B.n385 10.6151
R1325 B.n453 B.n452 10.6151
R1326 B.n457 B.n453 10.6151
R1327 B.n463 B.n383 10.6151
R1328 B.n464 B.n463 10.6151
R1329 B.n465 B.n464 10.6151
R1330 B.n465 B.n381 10.6151
R1331 B.n471 B.n381 10.6151
R1332 B.n472 B.n471 10.6151
R1333 B.n473 B.n472 10.6151
R1334 B.n473 B.n379 10.6151
R1335 B.n479 B.n379 10.6151
R1336 B.n482 B.n481 10.6151
R1337 B.n482 B.n375 10.6151
R1338 B.n488 B.n375 10.6151
R1339 B.n489 B.n488 10.6151
R1340 B.n490 B.n489 10.6151
R1341 B.n490 B.n373 10.6151
R1342 B.n496 B.n373 10.6151
R1343 B.n497 B.n496 10.6151
R1344 B.n498 B.n497 10.6151
R1345 B.n498 B.n371 10.6151
R1346 B.n504 B.n371 10.6151
R1347 B.n505 B.n504 10.6151
R1348 B.n506 B.n505 10.6151
R1349 B.n506 B.n369 10.6151
R1350 B.n512 B.n369 10.6151
R1351 B.n513 B.n512 10.6151
R1352 B.n514 B.n513 10.6151
R1353 B.n514 B.n367 10.6151
R1354 B.n520 B.n367 10.6151
R1355 B.n521 B.n520 10.6151
R1356 B.n522 B.n521 10.6151
R1357 B.n522 B.n365 10.6151
R1358 B.n528 B.n365 10.6151
R1359 B.n529 B.n528 10.6151
R1360 B.n530 B.n529 10.6151
R1361 B.n530 B.n363 10.6151
R1362 B.n363 B.n362 10.6151
R1363 B.n537 B.n362 10.6151
R1364 B.n538 B.n537 10.6151
R1365 B.n544 B.n543 10.6151
R1366 B.n545 B.n544 10.6151
R1367 B.n545 B.n350 10.6151
R1368 B.n555 B.n350 10.6151
R1369 B.n556 B.n555 10.6151
R1370 B.n557 B.n556 10.6151
R1371 B.n557 B.n342 10.6151
R1372 B.n567 B.n342 10.6151
R1373 B.n568 B.n567 10.6151
R1374 B.n569 B.n568 10.6151
R1375 B.n569 B.n334 10.6151
R1376 B.n579 B.n334 10.6151
R1377 B.n580 B.n579 10.6151
R1378 B.n581 B.n580 10.6151
R1379 B.n581 B.n326 10.6151
R1380 B.n591 B.n326 10.6151
R1381 B.n592 B.n591 10.6151
R1382 B.n593 B.n592 10.6151
R1383 B.n593 B.n318 10.6151
R1384 B.n603 B.n318 10.6151
R1385 B.n604 B.n603 10.6151
R1386 B.n605 B.n604 10.6151
R1387 B.n605 B.n310 10.6151
R1388 B.n615 B.n310 10.6151
R1389 B.n616 B.n615 10.6151
R1390 B.n617 B.n616 10.6151
R1391 B.n617 B.n302 10.6151
R1392 B.n627 B.n302 10.6151
R1393 B.n628 B.n627 10.6151
R1394 B.n629 B.n628 10.6151
R1395 B.n629 B.n294 10.6151
R1396 B.n639 B.n294 10.6151
R1397 B.n640 B.n639 10.6151
R1398 B.n641 B.n640 10.6151
R1399 B.n641 B.n286 10.6151
R1400 B.n651 B.n286 10.6151
R1401 B.n652 B.n651 10.6151
R1402 B.n653 B.n652 10.6151
R1403 B.n653 B.n278 10.6151
R1404 B.n663 B.n278 10.6151
R1405 B.n664 B.n663 10.6151
R1406 B.n665 B.n664 10.6151
R1407 B.n665 B.n270 10.6151
R1408 B.n676 B.n270 10.6151
R1409 B.n677 B.n676 10.6151
R1410 B.n678 B.n677 10.6151
R1411 B.n678 B.n0 10.6151
R1412 B.n841 B.n1 10.6151
R1413 B.n841 B.n840 10.6151
R1414 B.n840 B.n839 10.6151
R1415 B.n839 B.n10 10.6151
R1416 B.n833 B.n10 10.6151
R1417 B.n833 B.n832 10.6151
R1418 B.n832 B.n831 10.6151
R1419 B.n831 B.n17 10.6151
R1420 B.n825 B.n17 10.6151
R1421 B.n825 B.n824 10.6151
R1422 B.n824 B.n823 10.6151
R1423 B.n823 B.n24 10.6151
R1424 B.n817 B.n24 10.6151
R1425 B.n817 B.n816 10.6151
R1426 B.n816 B.n815 10.6151
R1427 B.n815 B.n31 10.6151
R1428 B.n809 B.n31 10.6151
R1429 B.n809 B.n808 10.6151
R1430 B.n808 B.n807 10.6151
R1431 B.n807 B.n38 10.6151
R1432 B.n801 B.n38 10.6151
R1433 B.n801 B.n800 10.6151
R1434 B.n800 B.n799 10.6151
R1435 B.n799 B.n45 10.6151
R1436 B.n793 B.n45 10.6151
R1437 B.n793 B.n792 10.6151
R1438 B.n792 B.n791 10.6151
R1439 B.n791 B.n52 10.6151
R1440 B.n785 B.n52 10.6151
R1441 B.n785 B.n784 10.6151
R1442 B.n784 B.n783 10.6151
R1443 B.n783 B.n59 10.6151
R1444 B.n777 B.n59 10.6151
R1445 B.n777 B.n776 10.6151
R1446 B.n776 B.n775 10.6151
R1447 B.n775 B.n66 10.6151
R1448 B.n769 B.n66 10.6151
R1449 B.n769 B.n768 10.6151
R1450 B.n768 B.n767 10.6151
R1451 B.n767 B.n73 10.6151
R1452 B.n761 B.n73 10.6151
R1453 B.n761 B.n760 10.6151
R1454 B.n760 B.n759 10.6151
R1455 B.n759 B.n80 10.6151
R1456 B.n753 B.n80 10.6151
R1457 B.n753 B.n752 10.6151
R1458 B.n752 B.n751 10.6151
R1459 B.n187 B.n130 9.36635
R1460 B.n210 B.n127 9.36635
R1461 B.n457 B.n456 9.36635
R1462 B.n481 B.n480 9.36635
R1463 B.n847 B.n0 2.81026
R1464 B.n847 B.n1 2.81026
R1465 B.n190 B.n130 1.24928
R1466 B.n207 B.n127 1.24928
R1467 B.n456 B.n383 1.24928
R1468 B.n480 B.n479 1.24928
R1469 VP.n16 VP.n13 161.3
R1470 VP.n18 VP.n17 161.3
R1471 VP.n19 VP.n12 161.3
R1472 VP.n21 VP.n20 161.3
R1473 VP.n22 VP.n11 161.3
R1474 VP.n24 VP.n23 161.3
R1475 VP.n26 VP.n10 161.3
R1476 VP.n28 VP.n27 161.3
R1477 VP.n29 VP.n9 161.3
R1478 VP.n31 VP.n30 161.3
R1479 VP.n32 VP.n8 161.3
R1480 VP.n62 VP.n0 161.3
R1481 VP.n61 VP.n60 161.3
R1482 VP.n59 VP.n1 161.3
R1483 VP.n58 VP.n57 161.3
R1484 VP.n56 VP.n2 161.3
R1485 VP.n54 VP.n53 161.3
R1486 VP.n52 VP.n3 161.3
R1487 VP.n51 VP.n50 161.3
R1488 VP.n49 VP.n4 161.3
R1489 VP.n48 VP.n47 161.3
R1490 VP.n46 VP.n5 161.3
R1491 VP.n45 VP.n44 161.3
R1492 VP.n42 VP.n6 161.3
R1493 VP.n41 VP.n40 161.3
R1494 VP.n39 VP.n7 161.3
R1495 VP.n38 VP.n37 161.3
R1496 VP.n15 VP.t5 114.957
R1497 VP.n36 VP.n35 95.3422
R1498 VP.n64 VP.n63 95.3422
R1499 VP.n34 VP.n33 95.3422
R1500 VP.n36 VP.t6 82.3253
R1501 VP.n43 VP.t7 82.3253
R1502 VP.n55 VP.t3 82.3253
R1503 VP.n63 VP.t4 82.3253
R1504 VP.n33 VP.t0 82.3253
R1505 VP.n25 VP.t2 82.3253
R1506 VP.n14 VP.t1 82.3253
R1507 VP.n15 VP.n14 66.9989
R1508 VP.n50 VP.n49 56.5193
R1509 VP.n20 VP.n19 56.5193
R1510 VP.n35 VP.n34 46.9844
R1511 VP.n42 VP.n41 44.3785
R1512 VP.n57 VP.n1 44.3785
R1513 VP.n27 VP.n9 44.3785
R1514 VP.n41 VP.n7 36.6083
R1515 VP.n61 VP.n1 36.6083
R1516 VP.n31 VP.n9 36.6083
R1517 VP.n37 VP.n7 24.4675
R1518 VP.n44 VP.n42 24.4675
R1519 VP.n48 VP.n5 24.4675
R1520 VP.n49 VP.n48 24.4675
R1521 VP.n50 VP.n3 24.4675
R1522 VP.n54 VP.n3 24.4675
R1523 VP.n57 VP.n56 24.4675
R1524 VP.n62 VP.n61 24.4675
R1525 VP.n32 VP.n31 24.4675
R1526 VP.n20 VP.n11 24.4675
R1527 VP.n24 VP.n11 24.4675
R1528 VP.n27 VP.n26 24.4675
R1529 VP.n18 VP.n13 24.4675
R1530 VP.n19 VP.n18 24.4675
R1531 VP.n44 VP.n43 19.3294
R1532 VP.n56 VP.n55 19.3294
R1533 VP.n26 VP.n25 19.3294
R1534 VP.n37 VP.n36 15.4147
R1535 VP.n63 VP.n62 15.4147
R1536 VP.n33 VP.n32 15.4147
R1537 VP.n16 VP.n15 9.45072
R1538 VP.n43 VP.n5 5.13857
R1539 VP.n55 VP.n54 5.13857
R1540 VP.n25 VP.n24 5.13857
R1541 VP.n14 VP.n13 5.13857
R1542 VP.n34 VP.n8 0.278367
R1543 VP.n38 VP.n35 0.278367
R1544 VP.n64 VP.n0 0.278367
R1545 VP.n17 VP.n16 0.189894
R1546 VP.n17 VP.n12 0.189894
R1547 VP.n21 VP.n12 0.189894
R1548 VP.n22 VP.n21 0.189894
R1549 VP.n23 VP.n22 0.189894
R1550 VP.n23 VP.n10 0.189894
R1551 VP.n28 VP.n10 0.189894
R1552 VP.n29 VP.n28 0.189894
R1553 VP.n30 VP.n29 0.189894
R1554 VP.n30 VP.n8 0.189894
R1555 VP.n39 VP.n38 0.189894
R1556 VP.n40 VP.n39 0.189894
R1557 VP.n40 VP.n6 0.189894
R1558 VP.n45 VP.n6 0.189894
R1559 VP.n46 VP.n45 0.189894
R1560 VP.n47 VP.n46 0.189894
R1561 VP.n47 VP.n4 0.189894
R1562 VP.n51 VP.n4 0.189894
R1563 VP.n52 VP.n51 0.189894
R1564 VP.n53 VP.n52 0.189894
R1565 VP.n53 VP.n2 0.189894
R1566 VP.n58 VP.n2 0.189894
R1567 VP.n59 VP.n58 0.189894
R1568 VP.n60 VP.n59 0.189894
R1569 VP.n60 VP.n0 0.189894
R1570 VP VP.n64 0.153454
R1571 VTAIL.n354 VTAIL.n316 289.615
R1572 VTAIL.n40 VTAIL.n2 289.615
R1573 VTAIL.n84 VTAIL.n46 289.615
R1574 VTAIL.n130 VTAIL.n92 289.615
R1575 VTAIL.n310 VTAIL.n272 289.615
R1576 VTAIL.n264 VTAIL.n226 289.615
R1577 VTAIL.n220 VTAIL.n182 289.615
R1578 VTAIL.n174 VTAIL.n136 289.615
R1579 VTAIL.n331 VTAIL.n330 185
R1580 VTAIL.n328 VTAIL.n327 185
R1581 VTAIL.n337 VTAIL.n336 185
R1582 VTAIL.n339 VTAIL.n338 185
R1583 VTAIL.n324 VTAIL.n323 185
R1584 VTAIL.n345 VTAIL.n344 185
R1585 VTAIL.n347 VTAIL.n346 185
R1586 VTAIL.n320 VTAIL.n319 185
R1587 VTAIL.n353 VTAIL.n352 185
R1588 VTAIL.n355 VTAIL.n354 185
R1589 VTAIL.n17 VTAIL.n16 185
R1590 VTAIL.n14 VTAIL.n13 185
R1591 VTAIL.n23 VTAIL.n22 185
R1592 VTAIL.n25 VTAIL.n24 185
R1593 VTAIL.n10 VTAIL.n9 185
R1594 VTAIL.n31 VTAIL.n30 185
R1595 VTAIL.n33 VTAIL.n32 185
R1596 VTAIL.n6 VTAIL.n5 185
R1597 VTAIL.n39 VTAIL.n38 185
R1598 VTAIL.n41 VTAIL.n40 185
R1599 VTAIL.n61 VTAIL.n60 185
R1600 VTAIL.n58 VTAIL.n57 185
R1601 VTAIL.n67 VTAIL.n66 185
R1602 VTAIL.n69 VTAIL.n68 185
R1603 VTAIL.n54 VTAIL.n53 185
R1604 VTAIL.n75 VTAIL.n74 185
R1605 VTAIL.n77 VTAIL.n76 185
R1606 VTAIL.n50 VTAIL.n49 185
R1607 VTAIL.n83 VTAIL.n82 185
R1608 VTAIL.n85 VTAIL.n84 185
R1609 VTAIL.n107 VTAIL.n106 185
R1610 VTAIL.n104 VTAIL.n103 185
R1611 VTAIL.n113 VTAIL.n112 185
R1612 VTAIL.n115 VTAIL.n114 185
R1613 VTAIL.n100 VTAIL.n99 185
R1614 VTAIL.n121 VTAIL.n120 185
R1615 VTAIL.n123 VTAIL.n122 185
R1616 VTAIL.n96 VTAIL.n95 185
R1617 VTAIL.n129 VTAIL.n128 185
R1618 VTAIL.n131 VTAIL.n130 185
R1619 VTAIL.n311 VTAIL.n310 185
R1620 VTAIL.n309 VTAIL.n308 185
R1621 VTAIL.n276 VTAIL.n275 185
R1622 VTAIL.n303 VTAIL.n302 185
R1623 VTAIL.n301 VTAIL.n300 185
R1624 VTAIL.n280 VTAIL.n279 185
R1625 VTAIL.n295 VTAIL.n294 185
R1626 VTAIL.n293 VTAIL.n292 185
R1627 VTAIL.n284 VTAIL.n283 185
R1628 VTAIL.n287 VTAIL.n286 185
R1629 VTAIL.n265 VTAIL.n264 185
R1630 VTAIL.n263 VTAIL.n262 185
R1631 VTAIL.n230 VTAIL.n229 185
R1632 VTAIL.n257 VTAIL.n256 185
R1633 VTAIL.n255 VTAIL.n254 185
R1634 VTAIL.n234 VTAIL.n233 185
R1635 VTAIL.n249 VTAIL.n248 185
R1636 VTAIL.n247 VTAIL.n246 185
R1637 VTAIL.n238 VTAIL.n237 185
R1638 VTAIL.n241 VTAIL.n240 185
R1639 VTAIL.n221 VTAIL.n220 185
R1640 VTAIL.n219 VTAIL.n218 185
R1641 VTAIL.n186 VTAIL.n185 185
R1642 VTAIL.n213 VTAIL.n212 185
R1643 VTAIL.n211 VTAIL.n210 185
R1644 VTAIL.n190 VTAIL.n189 185
R1645 VTAIL.n205 VTAIL.n204 185
R1646 VTAIL.n203 VTAIL.n202 185
R1647 VTAIL.n194 VTAIL.n193 185
R1648 VTAIL.n197 VTAIL.n196 185
R1649 VTAIL.n175 VTAIL.n174 185
R1650 VTAIL.n173 VTAIL.n172 185
R1651 VTAIL.n140 VTAIL.n139 185
R1652 VTAIL.n167 VTAIL.n166 185
R1653 VTAIL.n165 VTAIL.n164 185
R1654 VTAIL.n144 VTAIL.n143 185
R1655 VTAIL.n159 VTAIL.n158 185
R1656 VTAIL.n157 VTAIL.n156 185
R1657 VTAIL.n148 VTAIL.n147 185
R1658 VTAIL.n151 VTAIL.n150 185
R1659 VTAIL.t7 VTAIL.n329 147.659
R1660 VTAIL.t1 VTAIL.n15 147.659
R1661 VTAIL.t12 VTAIL.n59 147.659
R1662 VTAIL.t10 VTAIL.n105 147.659
R1663 VTAIL.t14 VTAIL.n285 147.659
R1664 VTAIL.t9 VTAIL.n239 147.659
R1665 VTAIL.t4 VTAIL.n195 147.659
R1666 VTAIL.t2 VTAIL.n149 147.659
R1667 VTAIL.n330 VTAIL.n327 104.615
R1668 VTAIL.n337 VTAIL.n327 104.615
R1669 VTAIL.n338 VTAIL.n337 104.615
R1670 VTAIL.n338 VTAIL.n323 104.615
R1671 VTAIL.n345 VTAIL.n323 104.615
R1672 VTAIL.n346 VTAIL.n345 104.615
R1673 VTAIL.n346 VTAIL.n319 104.615
R1674 VTAIL.n353 VTAIL.n319 104.615
R1675 VTAIL.n354 VTAIL.n353 104.615
R1676 VTAIL.n16 VTAIL.n13 104.615
R1677 VTAIL.n23 VTAIL.n13 104.615
R1678 VTAIL.n24 VTAIL.n23 104.615
R1679 VTAIL.n24 VTAIL.n9 104.615
R1680 VTAIL.n31 VTAIL.n9 104.615
R1681 VTAIL.n32 VTAIL.n31 104.615
R1682 VTAIL.n32 VTAIL.n5 104.615
R1683 VTAIL.n39 VTAIL.n5 104.615
R1684 VTAIL.n40 VTAIL.n39 104.615
R1685 VTAIL.n60 VTAIL.n57 104.615
R1686 VTAIL.n67 VTAIL.n57 104.615
R1687 VTAIL.n68 VTAIL.n67 104.615
R1688 VTAIL.n68 VTAIL.n53 104.615
R1689 VTAIL.n75 VTAIL.n53 104.615
R1690 VTAIL.n76 VTAIL.n75 104.615
R1691 VTAIL.n76 VTAIL.n49 104.615
R1692 VTAIL.n83 VTAIL.n49 104.615
R1693 VTAIL.n84 VTAIL.n83 104.615
R1694 VTAIL.n106 VTAIL.n103 104.615
R1695 VTAIL.n113 VTAIL.n103 104.615
R1696 VTAIL.n114 VTAIL.n113 104.615
R1697 VTAIL.n114 VTAIL.n99 104.615
R1698 VTAIL.n121 VTAIL.n99 104.615
R1699 VTAIL.n122 VTAIL.n121 104.615
R1700 VTAIL.n122 VTAIL.n95 104.615
R1701 VTAIL.n129 VTAIL.n95 104.615
R1702 VTAIL.n130 VTAIL.n129 104.615
R1703 VTAIL.n310 VTAIL.n309 104.615
R1704 VTAIL.n309 VTAIL.n275 104.615
R1705 VTAIL.n302 VTAIL.n275 104.615
R1706 VTAIL.n302 VTAIL.n301 104.615
R1707 VTAIL.n301 VTAIL.n279 104.615
R1708 VTAIL.n294 VTAIL.n279 104.615
R1709 VTAIL.n294 VTAIL.n293 104.615
R1710 VTAIL.n293 VTAIL.n283 104.615
R1711 VTAIL.n286 VTAIL.n283 104.615
R1712 VTAIL.n264 VTAIL.n263 104.615
R1713 VTAIL.n263 VTAIL.n229 104.615
R1714 VTAIL.n256 VTAIL.n229 104.615
R1715 VTAIL.n256 VTAIL.n255 104.615
R1716 VTAIL.n255 VTAIL.n233 104.615
R1717 VTAIL.n248 VTAIL.n233 104.615
R1718 VTAIL.n248 VTAIL.n247 104.615
R1719 VTAIL.n247 VTAIL.n237 104.615
R1720 VTAIL.n240 VTAIL.n237 104.615
R1721 VTAIL.n220 VTAIL.n219 104.615
R1722 VTAIL.n219 VTAIL.n185 104.615
R1723 VTAIL.n212 VTAIL.n185 104.615
R1724 VTAIL.n212 VTAIL.n211 104.615
R1725 VTAIL.n211 VTAIL.n189 104.615
R1726 VTAIL.n204 VTAIL.n189 104.615
R1727 VTAIL.n204 VTAIL.n203 104.615
R1728 VTAIL.n203 VTAIL.n193 104.615
R1729 VTAIL.n196 VTAIL.n193 104.615
R1730 VTAIL.n174 VTAIL.n173 104.615
R1731 VTAIL.n173 VTAIL.n139 104.615
R1732 VTAIL.n166 VTAIL.n139 104.615
R1733 VTAIL.n166 VTAIL.n165 104.615
R1734 VTAIL.n165 VTAIL.n143 104.615
R1735 VTAIL.n158 VTAIL.n143 104.615
R1736 VTAIL.n158 VTAIL.n157 104.615
R1737 VTAIL.n157 VTAIL.n147 104.615
R1738 VTAIL.n150 VTAIL.n147 104.615
R1739 VTAIL.n330 VTAIL.t7 52.3082
R1740 VTAIL.n16 VTAIL.t1 52.3082
R1741 VTAIL.n60 VTAIL.t12 52.3082
R1742 VTAIL.n106 VTAIL.t10 52.3082
R1743 VTAIL.n286 VTAIL.t14 52.3082
R1744 VTAIL.n240 VTAIL.t9 52.3082
R1745 VTAIL.n196 VTAIL.t4 52.3082
R1746 VTAIL.n150 VTAIL.t2 52.3082
R1747 VTAIL.n271 VTAIL.n270 47.2427
R1748 VTAIL.n181 VTAIL.n180 47.2427
R1749 VTAIL.n1 VTAIL.n0 47.2426
R1750 VTAIL.n91 VTAIL.n90 47.2426
R1751 VTAIL.n359 VTAIL.n358 31.6035
R1752 VTAIL.n45 VTAIL.n44 31.6035
R1753 VTAIL.n89 VTAIL.n88 31.6035
R1754 VTAIL.n135 VTAIL.n134 31.6035
R1755 VTAIL.n315 VTAIL.n314 31.6035
R1756 VTAIL.n269 VTAIL.n268 31.6035
R1757 VTAIL.n225 VTAIL.n224 31.6035
R1758 VTAIL.n179 VTAIL.n178 31.6035
R1759 VTAIL.n359 VTAIL.n315 21.7117
R1760 VTAIL.n179 VTAIL.n135 21.7117
R1761 VTAIL.n331 VTAIL.n329 15.6677
R1762 VTAIL.n17 VTAIL.n15 15.6677
R1763 VTAIL.n61 VTAIL.n59 15.6677
R1764 VTAIL.n107 VTAIL.n105 15.6677
R1765 VTAIL.n287 VTAIL.n285 15.6677
R1766 VTAIL.n241 VTAIL.n239 15.6677
R1767 VTAIL.n197 VTAIL.n195 15.6677
R1768 VTAIL.n151 VTAIL.n149 15.6677
R1769 VTAIL.n332 VTAIL.n328 12.8005
R1770 VTAIL.n18 VTAIL.n14 12.8005
R1771 VTAIL.n62 VTAIL.n58 12.8005
R1772 VTAIL.n108 VTAIL.n104 12.8005
R1773 VTAIL.n288 VTAIL.n284 12.8005
R1774 VTAIL.n242 VTAIL.n238 12.8005
R1775 VTAIL.n198 VTAIL.n194 12.8005
R1776 VTAIL.n152 VTAIL.n148 12.8005
R1777 VTAIL.n336 VTAIL.n335 12.0247
R1778 VTAIL.n22 VTAIL.n21 12.0247
R1779 VTAIL.n66 VTAIL.n65 12.0247
R1780 VTAIL.n112 VTAIL.n111 12.0247
R1781 VTAIL.n292 VTAIL.n291 12.0247
R1782 VTAIL.n246 VTAIL.n245 12.0247
R1783 VTAIL.n202 VTAIL.n201 12.0247
R1784 VTAIL.n156 VTAIL.n155 12.0247
R1785 VTAIL.n339 VTAIL.n326 11.249
R1786 VTAIL.n25 VTAIL.n12 11.249
R1787 VTAIL.n69 VTAIL.n56 11.249
R1788 VTAIL.n115 VTAIL.n102 11.249
R1789 VTAIL.n295 VTAIL.n282 11.249
R1790 VTAIL.n249 VTAIL.n236 11.249
R1791 VTAIL.n205 VTAIL.n192 11.249
R1792 VTAIL.n159 VTAIL.n146 11.249
R1793 VTAIL.n340 VTAIL.n324 10.4732
R1794 VTAIL.n26 VTAIL.n10 10.4732
R1795 VTAIL.n70 VTAIL.n54 10.4732
R1796 VTAIL.n116 VTAIL.n100 10.4732
R1797 VTAIL.n296 VTAIL.n280 10.4732
R1798 VTAIL.n250 VTAIL.n234 10.4732
R1799 VTAIL.n206 VTAIL.n190 10.4732
R1800 VTAIL.n160 VTAIL.n144 10.4732
R1801 VTAIL.n344 VTAIL.n343 9.69747
R1802 VTAIL.n30 VTAIL.n29 9.69747
R1803 VTAIL.n74 VTAIL.n73 9.69747
R1804 VTAIL.n120 VTAIL.n119 9.69747
R1805 VTAIL.n300 VTAIL.n299 9.69747
R1806 VTAIL.n254 VTAIL.n253 9.69747
R1807 VTAIL.n210 VTAIL.n209 9.69747
R1808 VTAIL.n164 VTAIL.n163 9.69747
R1809 VTAIL.n358 VTAIL.n357 9.45567
R1810 VTAIL.n44 VTAIL.n43 9.45567
R1811 VTAIL.n88 VTAIL.n87 9.45567
R1812 VTAIL.n134 VTAIL.n133 9.45567
R1813 VTAIL.n314 VTAIL.n313 9.45567
R1814 VTAIL.n268 VTAIL.n267 9.45567
R1815 VTAIL.n224 VTAIL.n223 9.45567
R1816 VTAIL.n178 VTAIL.n177 9.45567
R1817 VTAIL.n318 VTAIL.n317 9.3005
R1818 VTAIL.n357 VTAIL.n356 9.3005
R1819 VTAIL.n349 VTAIL.n348 9.3005
R1820 VTAIL.n322 VTAIL.n321 9.3005
R1821 VTAIL.n343 VTAIL.n342 9.3005
R1822 VTAIL.n341 VTAIL.n340 9.3005
R1823 VTAIL.n326 VTAIL.n325 9.3005
R1824 VTAIL.n335 VTAIL.n334 9.3005
R1825 VTAIL.n333 VTAIL.n332 9.3005
R1826 VTAIL.n351 VTAIL.n350 9.3005
R1827 VTAIL.n4 VTAIL.n3 9.3005
R1828 VTAIL.n43 VTAIL.n42 9.3005
R1829 VTAIL.n35 VTAIL.n34 9.3005
R1830 VTAIL.n8 VTAIL.n7 9.3005
R1831 VTAIL.n29 VTAIL.n28 9.3005
R1832 VTAIL.n27 VTAIL.n26 9.3005
R1833 VTAIL.n12 VTAIL.n11 9.3005
R1834 VTAIL.n21 VTAIL.n20 9.3005
R1835 VTAIL.n19 VTAIL.n18 9.3005
R1836 VTAIL.n37 VTAIL.n36 9.3005
R1837 VTAIL.n48 VTAIL.n47 9.3005
R1838 VTAIL.n87 VTAIL.n86 9.3005
R1839 VTAIL.n79 VTAIL.n78 9.3005
R1840 VTAIL.n52 VTAIL.n51 9.3005
R1841 VTAIL.n73 VTAIL.n72 9.3005
R1842 VTAIL.n71 VTAIL.n70 9.3005
R1843 VTAIL.n56 VTAIL.n55 9.3005
R1844 VTAIL.n65 VTAIL.n64 9.3005
R1845 VTAIL.n63 VTAIL.n62 9.3005
R1846 VTAIL.n81 VTAIL.n80 9.3005
R1847 VTAIL.n94 VTAIL.n93 9.3005
R1848 VTAIL.n133 VTAIL.n132 9.3005
R1849 VTAIL.n125 VTAIL.n124 9.3005
R1850 VTAIL.n98 VTAIL.n97 9.3005
R1851 VTAIL.n119 VTAIL.n118 9.3005
R1852 VTAIL.n117 VTAIL.n116 9.3005
R1853 VTAIL.n102 VTAIL.n101 9.3005
R1854 VTAIL.n111 VTAIL.n110 9.3005
R1855 VTAIL.n109 VTAIL.n108 9.3005
R1856 VTAIL.n127 VTAIL.n126 9.3005
R1857 VTAIL.n274 VTAIL.n273 9.3005
R1858 VTAIL.n307 VTAIL.n306 9.3005
R1859 VTAIL.n305 VTAIL.n304 9.3005
R1860 VTAIL.n278 VTAIL.n277 9.3005
R1861 VTAIL.n299 VTAIL.n298 9.3005
R1862 VTAIL.n297 VTAIL.n296 9.3005
R1863 VTAIL.n282 VTAIL.n281 9.3005
R1864 VTAIL.n291 VTAIL.n290 9.3005
R1865 VTAIL.n289 VTAIL.n288 9.3005
R1866 VTAIL.n313 VTAIL.n312 9.3005
R1867 VTAIL.n267 VTAIL.n266 9.3005
R1868 VTAIL.n228 VTAIL.n227 9.3005
R1869 VTAIL.n261 VTAIL.n260 9.3005
R1870 VTAIL.n259 VTAIL.n258 9.3005
R1871 VTAIL.n232 VTAIL.n231 9.3005
R1872 VTAIL.n253 VTAIL.n252 9.3005
R1873 VTAIL.n251 VTAIL.n250 9.3005
R1874 VTAIL.n236 VTAIL.n235 9.3005
R1875 VTAIL.n245 VTAIL.n244 9.3005
R1876 VTAIL.n243 VTAIL.n242 9.3005
R1877 VTAIL.n223 VTAIL.n222 9.3005
R1878 VTAIL.n184 VTAIL.n183 9.3005
R1879 VTAIL.n217 VTAIL.n216 9.3005
R1880 VTAIL.n215 VTAIL.n214 9.3005
R1881 VTAIL.n188 VTAIL.n187 9.3005
R1882 VTAIL.n209 VTAIL.n208 9.3005
R1883 VTAIL.n207 VTAIL.n206 9.3005
R1884 VTAIL.n192 VTAIL.n191 9.3005
R1885 VTAIL.n201 VTAIL.n200 9.3005
R1886 VTAIL.n199 VTAIL.n198 9.3005
R1887 VTAIL.n177 VTAIL.n176 9.3005
R1888 VTAIL.n138 VTAIL.n137 9.3005
R1889 VTAIL.n171 VTAIL.n170 9.3005
R1890 VTAIL.n169 VTAIL.n168 9.3005
R1891 VTAIL.n142 VTAIL.n141 9.3005
R1892 VTAIL.n163 VTAIL.n162 9.3005
R1893 VTAIL.n161 VTAIL.n160 9.3005
R1894 VTAIL.n146 VTAIL.n145 9.3005
R1895 VTAIL.n155 VTAIL.n154 9.3005
R1896 VTAIL.n153 VTAIL.n152 9.3005
R1897 VTAIL.n347 VTAIL.n322 8.92171
R1898 VTAIL.n33 VTAIL.n8 8.92171
R1899 VTAIL.n77 VTAIL.n52 8.92171
R1900 VTAIL.n123 VTAIL.n98 8.92171
R1901 VTAIL.n303 VTAIL.n278 8.92171
R1902 VTAIL.n257 VTAIL.n232 8.92171
R1903 VTAIL.n213 VTAIL.n188 8.92171
R1904 VTAIL.n167 VTAIL.n142 8.92171
R1905 VTAIL.n348 VTAIL.n320 8.14595
R1906 VTAIL.n358 VTAIL.n316 8.14595
R1907 VTAIL.n34 VTAIL.n6 8.14595
R1908 VTAIL.n44 VTAIL.n2 8.14595
R1909 VTAIL.n78 VTAIL.n50 8.14595
R1910 VTAIL.n88 VTAIL.n46 8.14595
R1911 VTAIL.n124 VTAIL.n96 8.14595
R1912 VTAIL.n134 VTAIL.n92 8.14595
R1913 VTAIL.n314 VTAIL.n272 8.14595
R1914 VTAIL.n304 VTAIL.n276 8.14595
R1915 VTAIL.n268 VTAIL.n226 8.14595
R1916 VTAIL.n258 VTAIL.n230 8.14595
R1917 VTAIL.n224 VTAIL.n182 8.14595
R1918 VTAIL.n214 VTAIL.n186 8.14595
R1919 VTAIL.n178 VTAIL.n136 8.14595
R1920 VTAIL.n168 VTAIL.n140 8.14595
R1921 VTAIL.n352 VTAIL.n351 7.3702
R1922 VTAIL.n356 VTAIL.n355 7.3702
R1923 VTAIL.n38 VTAIL.n37 7.3702
R1924 VTAIL.n42 VTAIL.n41 7.3702
R1925 VTAIL.n82 VTAIL.n81 7.3702
R1926 VTAIL.n86 VTAIL.n85 7.3702
R1927 VTAIL.n128 VTAIL.n127 7.3702
R1928 VTAIL.n132 VTAIL.n131 7.3702
R1929 VTAIL.n312 VTAIL.n311 7.3702
R1930 VTAIL.n308 VTAIL.n307 7.3702
R1931 VTAIL.n266 VTAIL.n265 7.3702
R1932 VTAIL.n262 VTAIL.n261 7.3702
R1933 VTAIL.n222 VTAIL.n221 7.3702
R1934 VTAIL.n218 VTAIL.n217 7.3702
R1935 VTAIL.n176 VTAIL.n175 7.3702
R1936 VTAIL.n172 VTAIL.n171 7.3702
R1937 VTAIL.n352 VTAIL.n318 6.59444
R1938 VTAIL.n355 VTAIL.n318 6.59444
R1939 VTAIL.n38 VTAIL.n4 6.59444
R1940 VTAIL.n41 VTAIL.n4 6.59444
R1941 VTAIL.n82 VTAIL.n48 6.59444
R1942 VTAIL.n85 VTAIL.n48 6.59444
R1943 VTAIL.n128 VTAIL.n94 6.59444
R1944 VTAIL.n131 VTAIL.n94 6.59444
R1945 VTAIL.n311 VTAIL.n274 6.59444
R1946 VTAIL.n308 VTAIL.n274 6.59444
R1947 VTAIL.n265 VTAIL.n228 6.59444
R1948 VTAIL.n262 VTAIL.n228 6.59444
R1949 VTAIL.n221 VTAIL.n184 6.59444
R1950 VTAIL.n218 VTAIL.n184 6.59444
R1951 VTAIL.n175 VTAIL.n138 6.59444
R1952 VTAIL.n172 VTAIL.n138 6.59444
R1953 VTAIL.n351 VTAIL.n320 5.81868
R1954 VTAIL.n356 VTAIL.n316 5.81868
R1955 VTAIL.n37 VTAIL.n6 5.81868
R1956 VTAIL.n42 VTAIL.n2 5.81868
R1957 VTAIL.n81 VTAIL.n50 5.81868
R1958 VTAIL.n86 VTAIL.n46 5.81868
R1959 VTAIL.n127 VTAIL.n96 5.81868
R1960 VTAIL.n132 VTAIL.n92 5.81868
R1961 VTAIL.n312 VTAIL.n272 5.81868
R1962 VTAIL.n307 VTAIL.n276 5.81868
R1963 VTAIL.n266 VTAIL.n226 5.81868
R1964 VTAIL.n261 VTAIL.n230 5.81868
R1965 VTAIL.n222 VTAIL.n182 5.81868
R1966 VTAIL.n217 VTAIL.n186 5.81868
R1967 VTAIL.n176 VTAIL.n136 5.81868
R1968 VTAIL.n171 VTAIL.n140 5.81868
R1969 VTAIL.n348 VTAIL.n347 5.04292
R1970 VTAIL.n34 VTAIL.n33 5.04292
R1971 VTAIL.n78 VTAIL.n77 5.04292
R1972 VTAIL.n124 VTAIL.n123 5.04292
R1973 VTAIL.n304 VTAIL.n303 5.04292
R1974 VTAIL.n258 VTAIL.n257 5.04292
R1975 VTAIL.n214 VTAIL.n213 5.04292
R1976 VTAIL.n168 VTAIL.n167 5.04292
R1977 VTAIL.n333 VTAIL.n329 4.38564
R1978 VTAIL.n19 VTAIL.n15 4.38564
R1979 VTAIL.n63 VTAIL.n59 4.38564
R1980 VTAIL.n109 VTAIL.n105 4.38564
R1981 VTAIL.n243 VTAIL.n239 4.38564
R1982 VTAIL.n199 VTAIL.n195 4.38564
R1983 VTAIL.n153 VTAIL.n149 4.38564
R1984 VTAIL.n289 VTAIL.n285 4.38564
R1985 VTAIL.n344 VTAIL.n322 4.26717
R1986 VTAIL.n30 VTAIL.n8 4.26717
R1987 VTAIL.n74 VTAIL.n52 4.26717
R1988 VTAIL.n120 VTAIL.n98 4.26717
R1989 VTAIL.n300 VTAIL.n278 4.26717
R1990 VTAIL.n254 VTAIL.n232 4.26717
R1991 VTAIL.n210 VTAIL.n188 4.26717
R1992 VTAIL.n164 VTAIL.n142 4.26717
R1993 VTAIL.n343 VTAIL.n324 3.49141
R1994 VTAIL.n29 VTAIL.n10 3.49141
R1995 VTAIL.n73 VTAIL.n54 3.49141
R1996 VTAIL.n119 VTAIL.n100 3.49141
R1997 VTAIL.n299 VTAIL.n280 3.49141
R1998 VTAIL.n253 VTAIL.n234 3.49141
R1999 VTAIL.n209 VTAIL.n190 3.49141
R2000 VTAIL.n163 VTAIL.n144 3.49141
R2001 VTAIL.n340 VTAIL.n339 2.71565
R2002 VTAIL.n26 VTAIL.n25 2.71565
R2003 VTAIL.n70 VTAIL.n69 2.71565
R2004 VTAIL.n116 VTAIL.n115 2.71565
R2005 VTAIL.n296 VTAIL.n295 2.71565
R2006 VTAIL.n250 VTAIL.n249 2.71565
R2007 VTAIL.n206 VTAIL.n205 2.71565
R2008 VTAIL.n160 VTAIL.n159 2.71565
R2009 VTAIL.n0 VTAIL.t0 2.43592
R2010 VTAIL.n0 VTAIL.t3 2.43592
R2011 VTAIL.n90 VTAIL.t15 2.43592
R2012 VTAIL.n90 VTAIL.t8 2.43592
R2013 VTAIL.n270 VTAIL.t13 2.43592
R2014 VTAIL.n270 VTAIL.t11 2.43592
R2015 VTAIL.n180 VTAIL.t6 2.43592
R2016 VTAIL.n180 VTAIL.t5 2.43592
R2017 VTAIL.n181 VTAIL.n179 2.33671
R2018 VTAIL.n225 VTAIL.n181 2.33671
R2019 VTAIL.n271 VTAIL.n269 2.33671
R2020 VTAIL.n315 VTAIL.n271 2.33671
R2021 VTAIL.n135 VTAIL.n91 2.33671
R2022 VTAIL.n91 VTAIL.n89 2.33671
R2023 VTAIL.n45 VTAIL.n1 2.33671
R2024 VTAIL VTAIL.n359 2.27852
R2025 VTAIL.n336 VTAIL.n326 1.93989
R2026 VTAIL.n22 VTAIL.n12 1.93989
R2027 VTAIL.n66 VTAIL.n56 1.93989
R2028 VTAIL.n112 VTAIL.n102 1.93989
R2029 VTAIL.n292 VTAIL.n282 1.93989
R2030 VTAIL.n246 VTAIL.n236 1.93989
R2031 VTAIL.n202 VTAIL.n192 1.93989
R2032 VTAIL.n156 VTAIL.n146 1.93989
R2033 VTAIL.n335 VTAIL.n328 1.16414
R2034 VTAIL.n21 VTAIL.n14 1.16414
R2035 VTAIL.n65 VTAIL.n58 1.16414
R2036 VTAIL.n111 VTAIL.n104 1.16414
R2037 VTAIL.n291 VTAIL.n284 1.16414
R2038 VTAIL.n245 VTAIL.n238 1.16414
R2039 VTAIL.n201 VTAIL.n194 1.16414
R2040 VTAIL.n155 VTAIL.n148 1.16414
R2041 VTAIL.n269 VTAIL.n225 0.470328
R2042 VTAIL.n89 VTAIL.n45 0.470328
R2043 VTAIL.n332 VTAIL.n331 0.388379
R2044 VTAIL.n18 VTAIL.n17 0.388379
R2045 VTAIL.n62 VTAIL.n61 0.388379
R2046 VTAIL.n108 VTAIL.n107 0.388379
R2047 VTAIL.n288 VTAIL.n287 0.388379
R2048 VTAIL.n242 VTAIL.n241 0.388379
R2049 VTAIL.n198 VTAIL.n197 0.388379
R2050 VTAIL.n152 VTAIL.n151 0.388379
R2051 VTAIL.n334 VTAIL.n333 0.155672
R2052 VTAIL.n334 VTAIL.n325 0.155672
R2053 VTAIL.n341 VTAIL.n325 0.155672
R2054 VTAIL.n342 VTAIL.n341 0.155672
R2055 VTAIL.n342 VTAIL.n321 0.155672
R2056 VTAIL.n349 VTAIL.n321 0.155672
R2057 VTAIL.n350 VTAIL.n349 0.155672
R2058 VTAIL.n350 VTAIL.n317 0.155672
R2059 VTAIL.n357 VTAIL.n317 0.155672
R2060 VTAIL.n20 VTAIL.n19 0.155672
R2061 VTAIL.n20 VTAIL.n11 0.155672
R2062 VTAIL.n27 VTAIL.n11 0.155672
R2063 VTAIL.n28 VTAIL.n27 0.155672
R2064 VTAIL.n28 VTAIL.n7 0.155672
R2065 VTAIL.n35 VTAIL.n7 0.155672
R2066 VTAIL.n36 VTAIL.n35 0.155672
R2067 VTAIL.n36 VTAIL.n3 0.155672
R2068 VTAIL.n43 VTAIL.n3 0.155672
R2069 VTAIL.n64 VTAIL.n63 0.155672
R2070 VTAIL.n64 VTAIL.n55 0.155672
R2071 VTAIL.n71 VTAIL.n55 0.155672
R2072 VTAIL.n72 VTAIL.n71 0.155672
R2073 VTAIL.n72 VTAIL.n51 0.155672
R2074 VTAIL.n79 VTAIL.n51 0.155672
R2075 VTAIL.n80 VTAIL.n79 0.155672
R2076 VTAIL.n80 VTAIL.n47 0.155672
R2077 VTAIL.n87 VTAIL.n47 0.155672
R2078 VTAIL.n110 VTAIL.n109 0.155672
R2079 VTAIL.n110 VTAIL.n101 0.155672
R2080 VTAIL.n117 VTAIL.n101 0.155672
R2081 VTAIL.n118 VTAIL.n117 0.155672
R2082 VTAIL.n118 VTAIL.n97 0.155672
R2083 VTAIL.n125 VTAIL.n97 0.155672
R2084 VTAIL.n126 VTAIL.n125 0.155672
R2085 VTAIL.n126 VTAIL.n93 0.155672
R2086 VTAIL.n133 VTAIL.n93 0.155672
R2087 VTAIL.n313 VTAIL.n273 0.155672
R2088 VTAIL.n306 VTAIL.n273 0.155672
R2089 VTAIL.n306 VTAIL.n305 0.155672
R2090 VTAIL.n305 VTAIL.n277 0.155672
R2091 VTAIL.n298 VTAIL.n277 0.155672
R2092 VTAIL.n298 VTAIL.n297 0.155672
R2093 VTAIL.n297 VTAIL.n281 0.155672
R2094 VTAIL.n290 VTAIL.n281 0.155672
R2095 VTAIL.n290 VTAIL.n289 0.155672
R2096 VTAIL.n267 VTAIL.n227 0.155672
R2097 VTAIL.n260 VTAIL.n227 0.155672
R2098 VTAIL.n260 VTAIL.n259 0.155672
R2099 VTAIL.n259 VTAIL.n231 0.155672
R2100 VTAIL.n252 VTAIL.n231 0.155672
R2101 VTAIL.n252 VTAIL.n251 0.155672
R2102 VTAIL.n251 VTAIL.n235 0.155672
R2103 VTAIL.n244 VTAIL.n235 0.155672
R2104 VTAIL.n244 VTAIL.n243 0.155672
R2105 VTAIL.n223 VTAIL.n183 0.155672
R2106 VTAIL.n216 VTAIL.n183 0.155672
R2107 VTAIL.n216 VTAIL.n215 0.155672
R2108 VTAIL.n215 VTAIL.n187 0.155672
R2109 VTAIL.n208 VTAIL.n187 0.155672
R2110 VTAIL.n208 VTAIL.n207 0.155672
R2111 VTAIL.n207 VTAIL.n191 0.155672
R2112 VTAIL.n200 VTAIL.n191 0.155672
R2113 VTAIL.n200 VTAIL.n199 0.155672
R2114 VTAIL.n177 VTAIL.n137 0.155672
R2115 VTAIL.n170 VTAIL.n137 0.155672
R2116 VTAIL.n170 VTAIL.n169 0.155672
R2117 VTAIL.n169 VTAIL.n141 0.155672
R2118 VTAIL.n162 VTAIL.n141 0.155672
R2119 VTAIL.n162 VTAIL.n161 0.155672
R2120 VTAIL.n161 VTAIL.n145 0.155672
R2121 VTAIL.n154 VTAIL.n145 0.155672
R2122 VTAIL.n154 VTAIL.n153 0.155672
R2123 VTAIL VTAIL.n1 0.0586897
R2124 VDD1 VDD1.n0 65.1478
R2125 VDD1.n3 VDD1.n2 65.0341
R2126 VDD1.n3 VDD1.n1 65.0341
R2127 VDD1.n5 VDD1.n4 63.9215
R2128 VDD1.n5 VDD1.n3 41.8199
R2129 VDD1.n4 VDD1.t5 2.43592
R2130 VDD1.n4 VDD1.t7 2.43592
R2131 VDD1.n0 VDD1.t2 2.43592
R2132 VDD1.n0 VDD1.t6 2.43592
R2133 VDD1.n2 VDD1.t4 2.43592
R2134 VDD1.n2 VDD1.t3 2.43592
R2135 VDD1.n1 VDD1.t1 2.43592
R2136 VDD1.n1 VDD1.t0 2.43592
R2137 VDD1 VDD1.n5 1.11041
R2138 VN.n51 VN.n27 161.3
R2139 VN.n50 VN.n49 161.3
R2140 VN.n48 VN.n28 161.3
R2141 VN.n47 VN.n46 161.3
R2142 VN.n45 VN.n29 161.3
R2143 VN.n43 VN.n42 161.3
R2144 VN.n41 VN.n30 161.3
R2145 VN.n40 VN.n39 161.3
R2146 VN.n38 VN.n31 161.3
R2147 VN.n37 VN.n36 161.3
R2148 VN.n35 VN.n32 161.3
R2149 VN.n24 VN.n0 161.3
R2150 VN.n23 VN.n22 161.3
R2151 VN.n21 VN.n1 161.3
R2152 VN.n20 VN.n19 161.3
R2153 VN.n18 VN.n2 161.3
R2154 VN.n16 VN.n15 161.3
R2155 VN.n14 VN.n3 161.3
R2156 VN.n13 VN.n12 161.3
R2157 VN.n11 VN.n4 161.3
R2158 VN.n10 VN.n9 161.3
R2159 VN.n8 VN.n5 161.3
R2160 VN.n7 VN.t4 114.957
R2161 VN.n34 VN.t6 114.957
R2162 VN.n26 VN.n25 95.3422
R2163 VN.n53 VN.n52 95.3422
R2164 VN.n6 VN.t3 82.3253
R2165 VN.n17 VN.t5 82.3253
R2166 VN.n25 VN.t1 82.3253
R2167 VN.n33 VN.t0 82.3253
R2168 VN.n44 VN.t7 82.3253
R2169 VN.n52 VN.t2 82.3253
R2170 VN.n7 VN.n6 66.9989
R2171 VN.n34 VN.n33 66.9989
R2172 VN.n12 VN.n11 56.5193
R2173 VN.n39 VN.n38 56.5193
R2174 VN VN.n53 47.2633
R2175 VN.n19 VN.n1 44.3785
R2176 VN.n46 VN.n28 44.3785
R2177 VN.n23 VN.n1 36.6083
R2178 VN.n50 VN.n28 36.6083
R2179 VN.n10 VN.n5 24.4675
R2180 VN.n11 VN.n10 24.4675
R2181 VN.n12 VN.n3 24.4675
R2182 VN.n16 VN.n3 24.4675
R2183 VN.n19 VN.n18 24.4675
R2184 VN.n24 VN.n23 24.4675
R2185 VN.n38 VN.n37 24.4675
R2186 VN.n37 VN.n32 24.4675
R2187 VN.n46 VN.n45 24.4675
R2188 VN.n43 VN.n30 24.4675
R2189 VN.n39 VN.n30 24.4675
R2190 VN.n51 VN.n50 24.4675
R2191 VN.n18 VN.n17 19.3294
R2192 VN.n45 VN.n44 19.3294
R2193 VN.n25 VN.n24 15.4147
R2194 VN.n52 VN.n51 15.4147
R2195 VN.n35 VN.n34 9.45072
R2196 VN.n8 VN.n7 9.45072
R2197 VN.n6 VN.n5 5.13857
R2198 VN.n17 VN.n16 5.13857
R2199 VN.n33 VN.n32 5.13857
R2200 VN.n44 VN.n43 5.13857
R2201 VN.n53 VN.n27 0.278367
R2202 VN.n26 VN.n0 0.278367
R2203 VN.n49 VN.n27 0.189894
R2204 VN.n49 VN.n48 0.189894
R2205 VN.n48 VN.n47 0.189894
R2206 VN.n47 VN.n29 0.189894
R2207 VN.n42 VN.n29 0.189894
R2208 VN.n42 VN.n41 0.189894
R2209 VN.n41 VN.n40 0.189894
R2210 VN.n40 VN.n31 0.189894
R2211 VN.n36 VN.n31 0.189894
R2212 VN.n36 VN.n35 0.189894
R2213 VN.n9 VN.n8 0.189894
R2214 VN.n9 VN.n4 0.189894
R2215 VN.n13 VN.n4 0.189894
R2216 VN.n14 VN.n13 0.189894
R2217 VN.n15 VN.n14 0.189894
R2218 VN.n15 VN.n2 0.189894
R2219 VN.n20 VN.n2 0.189894
R2220 VN.n21 VN.n20 0.189894
R2221 VN.n22 VN.n21 0.189894
R2222 VN.n22 VN.n0 0.189894
R2223 VN VN.n26 0.153454
R2224 VDD2.n2 VDD2.n1 65.0341
R2225 VDD2.n2 VDD2.n0 65.0341
R2226 VDD2 VDD2.n5 65.0314
R2227 VDD2.n4 VDD2.n3 63.9215
R2228 VDD2.n4 VDD2.n2 41.2368
R2229 VDD2.n5 VDD2.t7 2.43592
R2230 VDD2.n5 VDD2.t1 2.43592
R2231 VDD2.n3 VDD2.t5 2.43592
R2232 VDD2.n3 VDD2.t0 2.43592
R2233 VDD2.n1 VDD2.t2 2.43592
R2234 VDD2.n1 VDD2.t6 2.43592
R2235 VDD2.n0 VDD2.t3 2.43592
R2236 VDD2.n0 VDD2.t4 2.43592
R2237 VDD2 VDD2.n4 1.22679
C0 VTAIL VDD2 6.73952f
C1 VDD1 VP 6.27611f
C2 VN VP 6.67549f
C3 VDD1 VDD2 1.66038f
C4 VN VDD2 5.93246f
C5 VDD1 VTAIL 6.68658f
C6 VTAIL VN 6.41542f
C7 VDD2 VP 0.495899f
C8 VDD1 VN 0.150969f
C9 VTAIL VP 6.42952f
C10 VDD2 B 4.829567f
C11 VDD1 B 5.251309f
C12 VTAIL B 8.033463f
C13 VN B 14.3497f
C14 VP B 12.965909f
C15 VDD2.t3 B 0.155496f
C16 VDD2.t4 B 0.155496f
C17 VDD2.n0 B 1.34727f
C18 VDD2.t2 B 0.155496f
C19 VDD2.t6 B 0.155496f
C20 VDD2.n1 B 1.34727f
C21 VDD2.n2 B 2.82438f
C22 VDD2.t5 B 0.155496f
C23 VDD2.t0 B 0.155496f
C24 VDD2.n3 B 1.33904f
C25 VDD2.n4 B 2.49619f
C26 VDD2.t7 B 0.155496f
C27 VDD2.t1 B 0.155496f
C28 VDD2.n5 B 1.34725f
C29 VN.n0 B 0.032402f
C30 VN.t1 B 1.27806f
C31 VN.n1 B 0.020378f
C32 VN.n2 B 0.024577f
C33 VN.t5 B 1.27806f
C34 VN.n3 B 0.045805f
C35 VN.n4 B 0.024577f
C36 VN.n5 B 0.027939f
C37 VN.t4 B 1.45048f
C38 VN.t3 B 1.27806f
C39 VN.n6 B 0.52782f
C40 VN.n7 B 0.52067f
C41 VN.n8 B 0.213603f
C42 VN.n9 B 0.024577f
C43 VN.n10 B 0.045805f
C44 VN.n11 B 0.035878f
C45 VN.n12 B 0.035878f
C46 VN.n13 B 0.024577f
C47 VN.n14 B 0.024577f
C48 VN.n15 B 0.024577f
C49 VN.n16 B 0.027939f
C50 VN.n17 B 0.466846f
C51 VN.n18 B 0.041055f
C52 VN.n19 B 0.047629f
C53 VN.n20 B 0.024577f
C54 VN.n21 B 0.024577f
C55 VN.n22 B 0.024577f
C56 VN.n23 B 0.049553f
C57 VN.n24 B 0.037437f
C58 VN.n25 B 0.549528f
C59 VN.n26 B 0.034826f
C60 VN.n27 B 0.032402f
C61 VN.t2 B 1.27806f
C62 VN.n28 B 0.020378f
C63 VN.n29 B 0.024577f
C64 VN.t7 B 1.27806f
C65 VN.n30 B 0.045805f
C66 VN.n31 B 0.024577f
C67 VN.n32 B 0.027939f
C68 VN.t6 B 1.45048f
C69 VN.t0 B 1.27806f
C70 VN.n33 B 0.52782f
C71 VN.n34 B 0.52067f
C72 VN.n35 B 0.213603f
C73 VN.n36 B 0.024577f
C74 VN.n37 B 0.045805f
C75 VN.n38 B 0.035878f
C76 VN.n39 B 0.035878f
C77 VN.n40 B 0.024577f
C78 VN.n41 B 0.024577f
C79 VN.n42 B 0.024577f
C80 VN.n43 B 0.027939f
C81 VN.n44 B 0.466846f
C82 VN.n45 B 0.041055f
C83 VN.n46 B 0.047629f
C84 VN.n47 B 0.024577f
C85 VN.n48 B 0.024577f
C86 VN.n49 B 0.024577f
C87 VN.n50 B 0.049553f
C88 VN.n51 B 0.037437f
C89 VN.n52 B 0.549528f
C90 VN.n53 B 1.25465f
C91 VDD1.t2 B 0.159303f
C92 VDD1.t6 B 0.159303f
C93 VDD1.n0 B 1.38126f
C94 VDD1.t1 B 0.159303f
C95 VDD1.t0 B 0.159303f
C96 VDD1.n1 B 1.38025f
C97 VDD1.t4 B 0.159303f
C98 VDD1.t3 B 0.159303f
C99 VDD1.n2 B 1.38025f
C100 VDD1.n3 B 2.94542f
C101 VDD1.t5 B 0.159303f
C102 VDD1.t7 B 0.159303f
C103 VDD1.n4 B 1.37182f
C104 VDD1.n5 B 2.58767f
C105 VTAIL.t0 B 0.135675f
C106 VTAIL.t3 B 0.135675f
C107 VTAIL.n0 B 1.1075f
C108 VTAIL.n1 B 0.371427f
C109 VTAIL.n2 B 0.030966f
C110 VTAIL.n3 B 0.021118f
C111 VTAIL.n4 B 0.011348f
C112 VTAIL.n5 B 0.026822f
C113 VTAIL.n6 B 0.012016f
C114 VTAIL.n7 B 0.021118f
C115 VTAIL.n8 B 0.011348f
C116 VTAIL.n9 B 0.026822f
C117 VTAIL.n10 B 0.012016f
C118 VTAIL.n11 B 0.021118f
C119 VTAIL.n12 B 0.011348f
C120 VTAIL.n13 B 0.026822f
C121 VTAIL.n14 B 0.012016f
C122 VTAIL.n15 B 0.101404f
C123 VTAIL.t1 B 0.043749f
C124 VTAIL.n16 B 0.020117f
C125 VTAIL.n17 B 0.015845f
C126 VTAIL.n18 B 0.011348f
C127 VTAIL.n19 B 0.709001f
C128 VTAIL.n20 B 0.021118f
C129 VTAIL.n21 B 0.011348f
C130 VTAIL.n22 B 0.012016f
C131 VTAIL.n23 B 0.026822f
C132 VTAIL.n24 B 0.026822f
C133 VTAIL.n25 B 0.012016f
C134 VTAIL.n26 B 0.011348f
C135 VTAIL.n27 B 0.021118f
C136 VTAIL.n28 B 0.021118f
C137 VTAIL.n29 B 0.011348f
C138 VTAIL.n30 B 0.012016f
C139 VTAIL.n31 B 0.026822f
C140 VTAIL.n32 B 0.026822f
C141 VTAIL.n33 B 0.012016f
C142 VTAIL.n34 B 0.011348f
C143 VTAIL.n35 B 0.021118f
C144 VTAIL.n36 B 0.021118f
C145 VTAIL.n37 B 0.011348f
C146 VTAIL.n38 B 0.012016f
C147 VTAIL.n39 B 0.026822f
C148 VTAIL.n40 B 0.060334f
C149 VTAIL.n41 B 0.012016f
C150 VTAIL.n42 B 0.011348f
C151 VTAIL.n43 B 0.047948f
C152 VTAIL.n44 B 0.033965f
C153 VTAIL.n45 B 0.208491f
C154 VTAIL.n46 B 0.030966f
C155 VTAIL.n47 B 0.021118f
C156 VTAIL.n48 B 0.011348f
C157 VTAIL.n49 B 0.026822f
C158 VTAIL.n50 B 0.012016f
C159 VTAIL.n51 B 0.021118f
C160 VTAIL.n52 B 0.011348f
C161 VTAIL.n53 B 0.026822f
C162 VTAIL.n54 B 0.012016f
C163 VTAIL.n55 B 0.021118f
C164 VTAIL.n56 B 0.011348f
C165 VTAIL.n57 B 0.026822f
C166 VTAIL.n58 B 0.012016f
C167 VTAIL.n59 B 0.101404f
C168 VTAIL.t12 B 0.043749f
C169 VTAIL.n60 B 0.020117f
C170 VTAIL.n61 B 0.015845f
C171 VTAIL.n62 B 0.011348f
C172 VTAIL.n63 B 0.709001f
C173 VTAIL.n64 B 0.021118f
C174 VTAIL.n65 B 0.011348f
C175 VTAIL.n66 B 0.012016f
C176 VTAIL.n67 B 0.026822f
C177 VTAIL.n68 B 0.026822f
C178 VTAIL.n69 B 0.012016f
C179 VTAIL.n70 B 0.011348f
C180 VTAIL.n71 B 0.021118f
C181 VTAIL.n72 B 0.021118f
C182 VTAIL.n73 B 0.011348f
C183 VTAIL.n74 B 0.012016f
C184 VTAIL.n75 B 0.026822f
C185 VTAIL.n76 B 0.026822f
C186 VTAIL.n77 B 0.012016f
C187 VTAIL.n78 B 0.011348f
C188 VTAIL.n79 B 0.021118f
C189 VTAIL.n80 B 0.021118f
C190 VTAIL.n81 B 0.011348f
C191 VTAIL.n82 B 0.012016f
C192 VTAIL.n83 B 0.026822f
C193 VTAIL.n84 B 0.060334f
C194 VTAIL.n85 B 0.012016f
C195 VTAIL.n86 B 0.011348f
C196 VTAIL.n87 B 0.047948f
C197 VTAIL.n88 B 0.033965f
C198 VTAIL.n89 B 0.208491f
C199 VTAIL.t15 B 0.135675f
C200 VTAIL.t8 B 0.135675f
C201 VTAIL.n90 B 1.1075f
C202 VTAIL.n91 B 0.52644f
C203 VTAIL.n92 B 0.030966f
C204 VTAIL.n93 B 0.021118f
C205 VTAIL.n94 B 0.011348f
C206 VTAIL.n95 B 0.026822f
C207 VTAIL.n96 B 0.012016f
C208 VTAIL.n97 B 0.021118f
C209 VTAIL.n98 B 0.011348f
C210 VTAIL.n99 B 0.026822f
C211 VTAIL.n100 B 0.012016f
C212 VTAIL.n101 B 0.021118f
C213 VTAIL.n102 B 0.011348f
C214 VTAIL.n103 B 0.026822f
C215 VTAIL.n104 B 0.012016f
C216 VTAIL.n105 B 0.101404f
C217 VTAIL.t10 B 0.043749f
C218 VTAIL.n106 B 0.020117f
C219 VTAIL.n107 B 0.015845f
C220 VTAIL.n108 B 0.011348f
C221 VTAIL.n109 B 0.709001f
C222 VTAIL.n110 B 0.021118f
C223 VTAIL.n111 B 0.011348f
C224 VTAIL.n112 B 0.012016f
C225 VTAIL.n113 B 0.026822f
C226 VTAIL.n114 B 0.026822f
C227 VTAIL.n115 B 0.012016f
C228 VTAIL.n116 B 0.011348f
C229 VTAIL.n117 B 0.021118f
C230 VTAIL.n118 B 0.021118f
C231 VTAIL.n119 B 0.011348f
C232 VTAIL.n120 B 0.012016f
C233 VTAIL.n121 B 0.026822f
C234 VTAIL.n122 B 0.026822f
C235 VTAIL.n123 B 0.012016f
C236 VTAIL.n124 B 0.011348f
C237 VTAIL.n125 B 0.021118f
C238 VTAIL.n126 B 0.021118f
C239 VTAIL.n127 B 0.011348f
C240 VTAIL.n128 B 0.012016f
C241 VTAIL.n129 B 0.026822f
C242 VTAIL.n130 B 0.060334f
C243 VTAIL.n131 B 0.012016f
C244 VTAIL.n132 B 0.011348f
C245 VTAIL.n133 B 0.047948f
C246 VTAIL.n134 B 0.033965f
C247 VTAIL.n135 B 1.09927f
C248 VTAIL.n136 B 0.030966f
C249 VTAIL.n137 B 0.021118f
C250 VTAIL.n138 B 0.011348f
C251 VTAIL.n139 B 0.026822f
C252 VTAIL.n140 B 0.012016f
C253 VTAIL.n141 B 0.021118f
C254 VTAIL.n142 B 0.011348f
C255 VTAIL.n143 B 0.026822f
C256 VTAIL.n144 B 0.012016f
C257 VTAIL.n145 B 0.021118f
C258 VTAIL.n146 B 0.011348f
C259 VTAIL.n147 B 0.026822f
C260 VTAIL.n148 B 0.012016f
C261 VTAIL.n149 B 0.101404f
C262 VTAIL.t2 B 0.043749f
C263 VTAIL.n150 B 0.020117f
C264 VTAIL.n151 B 0.015845f
C265 VTAIL.n152 B 0.011348f
C266 VTAIL.n153 B 0.709001f
C267 VTAIL.n154 B 0.021118f
C268 VTAIL.n155 B 0.011348f
C269 VTAIL.n156 B 0.012016f
C270 VTAIL.n157 B 0.026822f
C271 VTAIL.n158 B 0.026822f
C272 VTAIL.n159 B 0.012016f
C273 VTAIL.n160 B 0.011348f
C274 VTAIL.n161 B 0.021118f
C275 VTAIL.n162 B 0.021118f
C276 VTAIL.n163 B 0.011348f
C277 VTAIL.n164 B 0.012016f
C278 VTAIL.n165 B 0.026822f
C279 VTAIL.n166 B 0.026822f
C280 VTAIL.n167 B 0.012016f
C281 VTAIL.n168 B 0.011348f
C282 VTAIL.n169 B 0.021118f
C283 VTAIL.n170 B 0.021118f
C284 VTAIL.n171 B 0.011348f
C285 VTAIL.n172 B 0.012016f
C286 VTAIL.n173 B 0.026822f
C287 VTAIL.n174 B 0.060334f
C288 VTAIL.n175 B 0.012016f
C289 VTAIL.n176 B 0.011348f
C290 VTAIL.n177 B 0.047948f
C291 VTAIL.n178 B 0.033965f
C292 VTAIL.n179 B 1.09927f
C293 VTAIL.t6 B 0.135675f
C294 VTAIL.t5 B 0.135675f
C295 VTAIL.n180 B 1.10751f
C296 VTAIL.n181 B 0.526432f
C297 VTAIL.n182 B 0.030966f
C298 VTAIL.n183 B 0.021118f
C299 VTAIL.n184 B 0.011348f
C300 VTAIL.n185 B 0.026822f
C301 VTAIL.n186 B 0.012016f
C302 VTAIL.n187 B 0.021118f
C303 VTAIL.n188 B 0.011348f
C304 VTAIL.n189 B 0.026822f
C305 VTAIL.n190 B 0.012016f
C306 VTAIL.n191 B 0.021118f
C307 VTAIL.n192 B 0.011348f
C308 VTAIL.n193 B 0.026822f
C309 VTAIL.n194 B 0.012016f
C310 VTAIL.n195 B 0.101404f
C311 VTAIL.t4 B 0.043749f
C312 VTAIL.n196 B 0.020117f
C313 VTAIL.n197 B 0.015845f
C314 VTAIL.n198 B 0.011348f
C315 VTAIL.n199 B 0.709001f
C316 VTAIL.n200 B 0.021118f
C317 VTAIL.n201 B 0.011348f
C318 VTAIL.n202 B 0.012016f
C319 VTAIL.n203 B 0.026822f
C320 VTAIL.n204 B 0.026822f
C321 VTAIL.n205 B 0.012016f
C322 VTAIL.n206 B 0.011348f
C323 VTAIL.n207 B 0.021118f
C324 VTAIL.n208 B 0.021118f
C325 VTAIL.n209 B 0.011348f
C326 VTAIL.n210 B 0.012016f
C327 VTAIL.n211 B 0.026822f
C328 VTAIL.n212 B 0.026822f
C329 VTAIL.n213 B 0.012016f
C330 VTAIL.n214 B 0.011348f
C331 VTAIL.n215 B 0.021118f
C332 VTAIL.n216 B 0.021118f
C333 VTAIL.n217 B 0.011348f
C334 VTAIL.n218 B 0.012016f
C335 VTAIL.n219 B 0.026822f
C336 VTAIL.n220 B 0.060334f
C337 VTAIL.n221 B 0.012016f
C338 VTAIL.n222 B 0.011348f
C339 VTAIL.n223 B 0.047948f
C340 VTAIL.n224 B 0.033965f
C341 VTAIL.n225 B 0.208491f
C342 VTAIL.n226 B 0.030966f
C343 VTAIL.n227 B 0.021118f
C344 VTAIL.n228 B 0.011348f
C345 VTAIL.n229 B 0.026822f
C346 VTAIL.n230 B 0.012016f
C347 VTAIL.n231 B 0.021118f
C348 VTAIL.n232 B 0.011348f
C349 VTAIL.n233 B 0.026822f
C350 VTAIL.n234 B 0.012016f
C351 VTAIL.n235 B 0.021118f
C352 VTAIL.n236 B 0.011348f
C353 VTAIL.n237 B 0.026822f
C354 VTAIL.n238 B 0.012016f
C355 VTAIL.n239 B 0.101404f
C356 VTAIL.t9 B 0.043749f
C357 VTAIL.n240 B 0.020117f
C358 VTAIL.n241 B 0.015845f
C359 VTAIL.n242 B 0.011348f
C360 VTAIL.n243 B 0.709001f
C361 VTAIL.n244 B 0.021118f
C362 VTAIL.n245 B 0.011348f
C363 VTAIL.n246 B 0.012016f
C364 VTAIL.n247 B 0.026822f
C365 VTAIL.n248 B 0.026822f
C366 VTAIL.n249 B 0.012016f
C367 VTAIL.n250 B 0.011348f
C368 VTAIL.n251 B 0.021118f
C369 VTAIL.n252 B 0.021118f
C370 VTAIL.n253 B 0.011348f
C371 VTAIL.n254 B 0.012016f
C372 VTAIL.n255 B 0.026822f
C373 VTAIL.n256 B 0.026822f
C374 VTAIL.n257 B 0.012016f
C375 VTAIL.n258 B 0.011348f
C376 VTAIL.n259 B 0.021118f
C377 VTAIL.n260 B 0.021118f
C378 VTAIL.n261 B 0.011348f
C379 VTAIL.n262 B 0.012016f
C380 VTAIL.n263 B 0.026822f
C381 VTAIL.n264 B 0.060334f
C382 VTAIL.n265 B 0.012016f
C383 VTAIL.n266 B 0.011348f
C384 VTAIL.n267 B 0.047948f
C385 VTAIL.n268 B 0.033965f
C386 VTAIL.n269 B 0.208491f
C387 VTAIL.t13 B 0.135675f
C388 VTAIL.t11 B 0.135675f
C389 VTAIL.n270 B 1.10751f
C390 VTAIL.n271 B 0.526432f
C391 VTAIL.n272 B 0.030966f
C392 VTAIL.n273 B 0.021118f
C393 VTAIL.n274 B 0.011348f
C394 VTAIL.n275 B 0.026822f
C395 VTAIL.n276 B 0.012016f
C396 VTAIL.n277 B 0.021118f
C397 VTAIL.n278 B 0.011348f
C398 VTAIL.n279 B 0.026822f
C399 VTAIL.n280 B 0.012016f
C400 VTAIL.n281 B 0.021118f
C401 VTAIL.n282 B 0.011348f
C402 VTAIL.n283 B 0.026822f
C403 VTAIL.n284 B 0.012016f
C404 VTAIL.n285 B 0.101404f
C405 VTAIL.t14 B 0.043749f
C406 VTAIL.n286 B 0.020117f
C407 VTAIL.n287 B 0.015845f
C408 VTAIL.n288 B 0.011348f
C409 VTAIL.n289 B 0.709001f
C410 VTAIL.n290 B 0.021118f
C411 VTAIL.n291 B 0.011348f
C412 VTAIL.n292 B 0.012016f
C413 VTAIL.n293 B 0.026822f
C414 VTAIL.n294 B 0.026822f
C415 VTAIL.n295 B 0.012016f
C416 VTAIL.n296 B 0.011348f
C417 VTAIL.n297 B 0.021118f
C418 VTAIL.n298 B 0.021118f
C419 VTAIL.n299 B 0.011348f
C420 VTAIL.n300 B 0.012016f
C421 VTAIL.n301 B 0.026822f
C422 VTAIL.n302 B 0.026822f
C423 VTAIL.n303 B 0.012016f
C424 VTAIL.n304 B 0.011348f
C425 VTAIL.n305 B 0.021118f
C426 VTAIL.n306 B 0.021118f
C427 VTAIL.n307 B 0.011348f
C428 VTAIL.n308 B 0.012016f
C429 VTAIL.n309 B 0.026822f
C430 VTAIL.n310 B 0.060334f
C431 VTAIL.n311 B 0.012016f
C432 VTAIL.n312 B 0.011348f
C433 VTAIL.n313 B 0.047948f
C434 VTAIL.n314 B 0.033965f
C435 VTAIL.n315 B 1.09927f
C436 VTAIL.n316 B 0.030966f
C437 VTAIL.n317 B 0.021118f
C438 VTAIL.n318 B 0.011348f
C439 VTAIL.n319 B 0.026822f
C440 VTAIL.n320 B 0.012016f
C441 VTAIL.n321 B 0.021118f
C442 VTAIL.n322 B 0.011348f
C443 VTAIL.n323 B 0.026822f
C444 VTAIL.n324 B 0.012016f
C445 VTAIL.n325 B 0.021118f
C446 VTAIL.n326 B 0.011348f
C447 VTAIL.n327 B 0.026822f
C448 VTAIL.n328 B 0.012016f
C449 VTAIL.n329 B 0.101404f
C450 VTAIL.t7 B 0.043749f
C451 VTAIL.n330 B 0.020117f
C452 VTAIL.n331 B 0.015845f
C453 VTAIL.n332 B 0.011348f
C454 VTAIL.n333 B 0.709001f
C455 VTAIL.n334 B 0.021118f
C456 VTAIL.n335 B 0.011348f
C457 VTAIL.n336 B 0.012016f
C458 VTAIL.n337 B 0.026822f
C459 VTAIL.n338 B 0.026822f
C460 VTAIL.n339 B 0.012016f
C461 VTAIL.n340 B 0.011348f
C462 VTAIL.n341 B 0.021118f
C463 VTAIL.n342 B 0.021118f
C464 VTAIL.n343 B 0.011348f
C465 VTAIL.n344 B 0.012016f
C466 VTAIL.n345 B 0.026822f
C467 VTAIL.n346 B 0.026822f
C468 VTAIL.n347 B 0.012016f
C469 VTAIL.n348 B 0.011348f
C470 VTAIL.n349 B 0.021118f
C471 VTAIL.n350 B 0.021118f
C472 VTAIL.n351 B 0.011348f
C473 VTAIL.n352 B 0.012016f
C474 VTAIL.n353 B 0.026822f
C475 VTAIL.n354 B 0.060334f
C476 VTAIL.n355 B 0.012016f
C477 VTAIL.n356 B 0.011348f
C478 VTAIL.n357 B 0.047948f
C479 VTAIL.n358 B 0.033965f
C480 VTAIL.n359 B 1.09531f
C481 VP.n0 B 0.033144f
C482 VP.t4 B 1.30734f
C483 VP.n1 B 0.020845f
C484 VP.n2 B 0.02514f
C485 VP.t3 B 1.30734f
C486 VP.n3 B 0.046854f
C487 VP.n4 B 0.02514f
C488 VP.n5 B 0.028579f
C489 VP.n6 B 0.02514f
C490 VP.n7 B 0.050689f
C491 VP.n8 B 0.033144f
C492 VP.t0 B 1.30734f
C493 VP.n9 B 0.020845f
C494 VP.n10 B 0.02514f
C495 VP.t2 B 1.30734f
C496 VP.n11 B 0.046854f
C497 VP.n12 B 0.02514f
C498 VP.n13 B 0.028579f
C499 VP.t5 B 1.48371f
C500 VP.t1 B 1.30734f
C501 VP.n14 B 0.539914f
C502 VP.n15 B 0.5326f
C503 VP.n16 B 0.218498f
C504 VP.n17 B 0.02514f
C505 VP.n18 B 0.046854f
C506 VP.n19 B 0.0367f
C507 VP.n20 B 0.0367f
C508 VP.n21 B 0.02514f
C509 VP.n22 B 0.02514f
C510 VP.n23 B 0.02514f
C511 VP.n24 B 0.028579f
C512 VP.n25 B 0.477542f
C513 VP.n26 B 0.041995f
C514 VP.n27 B 0.048721f
C515 VP.n28 B 0.02514f
C516 VP.n29 B 0.02514f
C517 VP.n30 B 0.02514f
C518 VP.n31 B 0.050689f
C519 VP.n32 B 0.038294f
C520 VP.n33 B 0.56212f
C521 VP.n34 B 1.26975f
C522 VP.n35 B 1.28899f
C523 VP.t6 B 1.30734f
C524 VP.n36 B 0.56212f
C525 VP.n37 B 0.038294f
C526 VP.n38 B 0.033144f
C527 VP.n39 B 0.02514f
C528 VP.n40 B 0.02514f
C529 VP.n41 B 0.020845f
C530 VP.n42 B 0.048721f
C531 VP.t7 B 1.30734f
C532 VP.n43 B 0.477542f
C533 VP.n44 B 0.041995f
C534 VP.n45 B 0.02514f
C535 VP.n46 B 0.02514f
C536 VP.n47 B 0.02514f
C537 VP.n48 B 0.046854f
C538 VP.n49 B 0.0367f
C539 VP.n50 B 0.0367f
C540 VP.n51 B 0.02514f
C541 VP.n52 B 0.02514f
C542 VP.n53 B 0.02514f
C543 VP.n54 B 0.028579f
C544 VP.n55 B 0.477542f
C545 VP.n56 B 0.041995f
C546 VP.n57 B 0.048721f
C547 VP.n58 B 0.02514f
C548 VP.n59 B 0.02514f
C549 VP.n60 B 0.02514f
C550 VP.n61 B 0.050689f
C551 VP.n62 B 0.038294f
C552 VP.n63 B 0.56212f
C553 VP.n64 B 0.035624f
.ends

