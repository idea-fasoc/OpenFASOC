* NGSPICE file created from diff_pair_sample_1237.ext - technology: sky130A

.subckt diff_pair_sample_1237 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=0 ps=0 w=6.4 l=0.27
X2 VTAIL.t4 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X3 VDD2.t6 VN.t1 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=2.496 ps=13.58 w=6.4 l=0.27
X4 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X5 VTAIL.t6 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=1.056 ps=6.73 w=6.4 l=0.27
X6 VTAIL.t10 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=1.056 ps=6.73 w=6.4 l=0.27
X7 VDD2.t4 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=0 ps=0 w=6.4 l=0.27
X9 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X10 VDD2.t3 VN.t4 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=2.496 ps=13.58 w=6.4 l=0.27
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=0 ps=0 w=6.4 l=0.27
X12 VDD1.t3 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X13 VTAIL.t8 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=1.056 ps=6.73 w=6.4 l=0.27
X14 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=2.496 ps=13.58 w=6.4 l=0.27
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=0 ps=0 w=6.4 l=0.27
X16 VTAIL.t14 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X17 VDD1.t1 VP.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=2.496 ps=13.58 w=6.4 l=0.27
X18 VTAIL.t15 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.056 pd=6.73 as=1.056 ps=6.73 w=6.4 l=0.27
X19 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.496 pd=13.58 as=1.056 ps=6.73 w=6.4 l=0.27
R0 VN.n5 VN.t1 745.721
R1 VN.n1 VN.t5 745.721
R2 VN.n12 VN.t2 745.721
R3 VN.n8 VN.t4 745.721
R4 VN.n4 VN.t7 687.297
R5 VN.n2 VN.t3 687.297
R6 VN.n11 VN.t0 687.297
R7 VN.n9 VN.t6 687.297
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN.n3 VN.n2 43.8187
R15 VN.n4 VN.n3 43.8187
R16 VN.n11 VN.n10 43.8187
R17 VN.n10 VN.n9 43.8187
R18 VN VN.n13 36.2827
R19 VN.n2 VN.n1 29.2126
R20 VN.n5 VN.n4 29.2126
R21 VN.n12 VN.n11 29.2126
R22 VN.n9 VN.n8 29.2126
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VTAIL.n11 VTAIL.t3 53.7867
R27 VTAIL.n10 VTAIL.t13 53.7867
R28 VTAIL.n7 VTAIL.t10 53.7867
R29 VTAIL.n15 VTAIL.t9 53.7866
R30 VTAIL.n2 VTAIL.t8 53.7866
R31 VTAIL.n3 VTAIL.t2 53.7866
R32 VTAIL.n6 VTAIL.t6 53.7866
R33 VTAIL.n14 VTAIL.t0 53.7866
R34 VTAIL.n13 VTAIL.n12 50.693
R35 VTAIL.n9 VTAIL.n8 50.693
R36 VTAIL.n1 VTAIL.n0 50.6928
R37 VTAIL.n5 VTAIL.n4 50.6928
R38 VTAIL.n15 VTAIL.n14 18.4014
R39 VTAIL.n7 VTAIL.n6 18.4014
R40 VTAIL.n0 VTAIL.t12 3.09425
R41 VTAIL.n0 VTAIL.t15 3.09425
R42 VTAIL.n4 VTAIL.t1 3.09425
R43 VTAIL.n4 VTAIL.t4 3.09425
R44 VTAIL.n12 VTAIL.t5 3.09425
R45 VTAIL.n12 VTAIL.t7 3.09425
R46 VTAIL.n8 VTAIL.t11 3.09425
R47 VTAIL.n8 VTAIL.t14 3.09425
R48 VTAIL.n9 VTAIL.n7 0.517741
R49 VTAIL.n10 VTAIL.n9 0.517741
R50 VTAIL.n13 VTAIL.n11 0.517741
R51 VTAIL.n14 VTAIL.n13 0.517741
R52 VTAIL.n6 VTAIL.n5 0.517741
R53 VTAIL.n5 VTAIL.n3 0.517741
R54 VTAIL.n2 VTAIL.n1 0.517741
R55 VTAIL.n11 VTAIL.n10 0.470328
R56 VTAIL.n3 VTAIL.n2 0.470328
R57 VTAIL VTAIL.n15 0.459552
R58 VTAIL VTAIL.n1 0.0586897
R59 VDD2.n2 VDD2.n1 67.5749
R60 VDD2.n2 VDD2.n0 67.5749
R61 VDD2 VDD2.n5 67.5721
R62 VDD2.n4 VDD2.n3 67.3718
R63 VDD2.n4 VDD2.n2 31.5601
R64 VDD2.n5 VDD2.t1 3.09425
R65 VDD2.n5 VDD2.t3 3.09425
R66 VDD2.n3 VDD2.t5 3.09425
R67 VDD2.n3 VDD2.t7 3.09425
R68 VDD2.n1 VDD2.t0 3.09425
R69 VDD2.n1 VDD2.t6 3.09425
R70 VDD2.n0 VDD2.t2 3.09425
R71 VDD2.n0 VDD2.t4 3.09425
R72 VDD2 VDD2.n4 0.31731
R73 B.n252 B.t8 791.99
R74 B.n249 B.t19 791.99
R75 B.n66 B.t16 791.99
R76 B.n64 B.t12 791.99
R77 B.n449 B.n448 585
R78 B.n186 B.n63 585
R79 B.n185 B.n184 585
R80 B.n183 B.n182 585
R81 B.n181 B.n180 585
R82 B.n179 B.n178 585
R83 B.n177 B.n176 585
R84 B.n175 B.n174 585
R85 B.n173 B.n172 585
R86 B.n171 B.n170 585
R87 B.n169 B.n168 585
R88 B.n167 B.n166 585
R89 B.n165 B.n164 585
R90 B.n163 B.n162 585
R91 B.n161 B.n160 585
R92 B.n159 B.n158 585
R93 B.n157 B.n156 585
R94 B.n155 B.n154 585
R95 B.n153 B.n152 585
R96 B.n151 B.n150 585
R97 B.n149 B.n148 585
R98 B.n147 B.n146 585
R99 B.n145 B.n144 585
R100 B.n143 B.n142 585
R101 B.n141 B.n140 585
R102 B.n138 B.n137 585
R103 B.n136 B.n135 585
R104 B.n134 B.n133 585
R105 B.n132 B.n131 585
R106 B.n130 B.n129 585
R107 B.n128 B.n127 585
R108 B.n126 B.n125 585
R109 B.n124 B.n123 585
R110 B.n122 B.n121 585
R111 B.n120 B.n119 585
R112 B.n117 B.n116 585
R113 B.n115 B.n114 585
R114 B.n113 B.n112 585
R115 B.n111 B.n110 585
R116 B.n109 B.n108 585
R117 B.n107 B.n106 585
R118 B.n105 B.n104 585
R119 B.n103 B.n102 585
R120 B.n101 B.n100 585
R121 B.n99 B.n98 585
R122 B.n97 B.n96 585
R123 B.n95 B.n94 585
R124 B.n93 B.n92 585
R125 B.n91 B.n90 585
R126 B.n89 B.n88 585
R127 B.n87 B.n86 585
R128 B.n85 B.n84 585
R129 B.n83 B.n82 585
R130 B.n81 B.n80 585
R131 B.n79 B.n78 585
R132 B.n77 B.n76 585
R133 B.n75 B.n74 585
R134 B.n73 B.n72 585
R135 B.n71 B.n70 585
R136 B.n69 B.n68 585
R137 B.n447 B.n33 585
R138 B.n452 B.n33 585
R139 B.n446 B.n32 585
R140 B.n453 B.n32 585
R141 B.n445 B.n444 585
R142 B.n444 B.n28 585
R143 B.n443 B.n27 585
R144 B.n459 B.n27 585
R145 B.n442 B.n26 585
R146 B.n460 B.n26 585
R147 B.n441 B.n25 585
R148 B.n461 B.n25 585
R149 B.n440 B.n439 585
R150 B.n439 B.n21 585
R151 B.n438 B.n20 585
R152 B.n467 B.n20 585
R153 B.n437 B.n19 585
R154 B.n468 B.n19 585
R155 B.n436 B.n18 585
R156 B.n469 B.n18 585
R157 B.n435 B.n434 585
R158 B.n434 B.n433 585
R159 B.n432 B.n14 585
R160 B.n475 B.n14 585
R161 B.n431 B.n13 585
R162 B.n476 B.n13 585
R163 B.n430 B.n12 585
R164 B.n477 B.n12 585
R165 B.n429 B.n428 585
R166 B.n428 B.n11 585
R167 B.n427 B.n7 585
R168 B.n483 B.n7 585
R169 B.n426 B.n6 585
R170 B.n484 B.n6 585
R171 B.n425 B.n5 585
R172 B.n485 B.n5 585
R173 B.n424 B.n423 585
R174 B.n423 B.n4 585
R175 B.n422 B.n187 585
R176 B.n422 B.n421 585
R177 B.n411 B.n188 585
R178 B.n414 B.n188 585
R179 B.n413 B.n412 585
R180 B.n415 B.n413 585
R181 B.n410 B.n192 585
R182 B.n195 B.n192 585
R183 B.n409 B.n408 585
R184 B.n408 B.n407 585
R185 B.n194 B.n193 585
R186 B.n400 B.n194 585
R187 B.n399 B.n398 585
R188 B.n401 B.n399 585
R189 B.n397 B.n200 585
R190 B.n200 B.n199 585
R191 B.n396 B.n395 585
R192 B.n395 B.n394 585
R193 B.n202 B.n201 585
R194 B.n203 B.n202 585
R195 B.n387 B.n386 585
R196 B.n388 B.n387 585
R197 B.n385 B.n207 585
R198 B.n211 B.n207 585
R199 B.n384 B.n383 585
R200 B.n383 B.n382 585
R201 B.n209 B.n208 585
R202 B.n210 B.n209 585
R203 B.n375 B.n374 585
R204 B.n376 B.n375 585
R205 B.n373 B.n216 585
R206 B.n216 B.n215 585
R207 B.n368 B.n367 585
R208 B.n366 B.n248 585
R209 B.n365 B.n247 585
R210 B.n370 B.n247 585
R211 B.n364 B.n363 585
R212 B.n362 B.n361 585
R213 B.n360 B.n359 585
R214 B.n358 B.n357 585
R215 B.n356 B.n355 585
R216 B.n354 B.n353 585
R217 B.n352 B.n351 585
R218 B.n350 B.n349 585
R219 B.n348 B.n347 585
R220 B.n346 B.n345 585
R221 B.n344 B.n343 585
R222 B.n342 B.n341 585
R223 B.n340 B.n339 585
R224 B.n338 B.n337 585
R225 B.n336 B.n335 585
R226 B.n334 B.n333 585
R227 B.n332 B.n331 585
R228 B.n330 B.n329 585
R229 B.n328 B.n327 585
R230 B.n326 B.n325 585
R231 B.n324 B.n323 585
R232 B.n322 B.n321 585
R233 B.n320 B.n319 585
R234 B.n318 B.n317 585
R235 B.n316 B.n315 585
R236 B.n314 B.n313 585
R237 B.n312 B.n311 585
R238 B.n310 B.n309 585
R239 B.n308 B.n307 585
R240 B.n306 B.n305 585
R241 B.n304 B.n303 585
R242 B.n302 B.n301 585
R243 B.n300 B.n299 585
R244 B.n298 B.n297 585
R245 B.n296 B.n295 585
R246 B.n294 B.n293 585
R247 B.n292 B.n291 585
R248 B.n290 B.n289 585
R249 B.n288 B.n287 585
R250 B.n286 B.n285 585
R251 B.n284 B.n283 585
R252 B.n282 B.n281 585
R253 B.n280 B.n279 585
R254 B.n278 B.n277 585
R255 B.n276 B.n275 585
R256 B.n274 B.n273 585
R257 B.n272 B.n271 585
R258 B.n270 B.n269 585
R259 B.n268 B.n267 585
R260 B.n266 B.n265 585
R261 B.n264 B.n263 585
R262 B.n262 B.n261 585
R263 B.n260 B.n259 585
R264 B.n258 B.n257 585
R265 B.n256 B.n255 585
R266 B.n218 B.n217 585
R267 B.n372 B.n371 585
R268 B.n371 B.n370 585
R269 B.n214 B.n213 585
R270 B.n215 B.n214 585
R271 B.n378 B.n377 585
R272 B.n377 B.n376 585
R273 B.n379 B.n212 585
R274 B.n212 B.n210 585
R275 B.n381 B.n380 585
R276 B.n382 B.n381 585
R277 B.n206 B.n205 585
R278 B.n211 B.n206 585
R279 B.n390 B.n389 585
R280 B.n389 B.n388 585
R281 B.n391 B.n204 585
R282 B.n204 B.n203 585
R283 B.n393 B.n392 585
R284 B.n394 B.n393 585
R285 B.n198 B.n197 585
R286 B.n199 B.n198 585
R287 B.n403 B.n402 585
R288 B.n402 B.n401 585
R289 B.n404 B.n196 585
R290 B.n400 B.n196 585
R291 B.n406 B.n405 585
R292 B.n407 B.n406 585
R293 B.n191 B.n190 585
R294 B.n195 B.n191 585
R295 B.n417 B.n416 585
R296 B.n416 B.n415 585
R297 B.n418 B.n189 585
R298 B.n414 B.n189 585
R299 B.n420 B.n419 585
R300 B.n421 B.n420 585
R301 B.n2 B.n0 585
R302 B.n4 B.n2 585
R303 B.n3 B.n1 585
R304 B.n484 B.n3 585
R305 B.n482 B.n481 585
R306 B.n483 B.n482 585
R307 B.n480 B.n8 585
R308 B.n11 B.n8 585
R309 B.n479 B.n478 585
R310 B.n478 B.n477 585
R311 B.n10 B.n9 585
R312 B.n476 B.n10 585
R313 B.n474 B.n473 585
R314 B.n475 B.n474 585
R315 B.n472 B.n15 585
R316 B.n433 B.n15 585
R317 B.n471 B.n470 585
R318 B.n470 B.n469 585
R319 B.n17 B.n16 585
R320 B.n468 B.n17 585
R321 B.n466 B.n465 585
R322 B.n467 B.n466 585
R323 B.n464 B.n22 585
R324 B.n22 B.n21 585
R325 B.n463 B.n462 585
R326 B.n462 B.n461 585
R327 B.n24 B.n23 585
R328 B.n460 B.n24 585
R329 B.n458 B.n457 585
R330 B.n459 B.n458 585
R331 B.n456 B.n29 585
R332 B.n29 B.n28 585
R333 B.n455 B.n454 585
R334 B.n454 B.n453 585
R335 B.n31 B.n30 585
R336 B.n452 B.n31 585
R337 B.n487 B.n486 585
R338 B.n486 B.n485 585
R339 B.n368 B.n214 478.086
R340 B.n68 B.n31 478.086
R341 B.n371 B.n216 478.086
R342 B.n449 B.n33 478.086
R343 B.n451 B.n450 256.663
R344 B.n451 B.n62 256.663
R345 B.n451 B.n61 256.663
R346 B.n451 B.n60 256.663
R347 B.n451 B.n59 256.663
R348 B.n451 B.n58 256.663
R349 B.n451 B.n57 256.663
R350 B.n451 B.n56 256.663
R351 B.n451 B.n55 256.663
R352 B.n451 B.n54 256.663
R353 B.n451 B.n53 256.663
R354 B.n451 B.n52 256.663
R355 B.n451 B.n51 256.663
R356 B.n451 B.n50 256.663
R357 B.n451 B.n49 256.663
R358 B.n451 B.n48 256.663
R359 B.n451 B.n47 256.663
R360 B.n451 B.n46 256.663
R361 B.n451 B.n45 256.663
R362 B.n451 B.n44 256.663
R363 B.n451 B.n43 256.663
R364 B.n451 B.n42 256.663
R365 B.n451 B.n41 256.663
R366 B.n451 B.n40 256.663
R367 B.n451 B.n39 256.663
R368 B.n451 B.n38 256.663
R369 B.n451 B.n37 256.663
R370 B.n451 B.n36 256.663
R371 B.n451 B.n35 256.663
R372 B.n451 B.n34 256.663
R373 B.n370 B.n369 256.663
R374 B.n370 B.n219 256.663
R375 B.n370 B.n220 256.663
R376 B.n370 B.n221 256.663
R377 B.n370 B.n222 256.663
R378 B.n370 B.n223 256.663
R379 B.n370 B.n224 256.663
R380 B.n370 B.n225 256.663
R381 B.n370 B.n226 256.663
R382 B.n370 B.n227 256.663
R383 B.n370 B.n228 256.663
R384 B.n370 B.n229 256.663
R385 B.n370 B.n230 256.663
R386 B.n370 B.n231 256.663
R387 B.n370 B.n232 256.663
R388 B.n370 B.n233 256.663
R389 B.n370 B.n234 256.663
R390 B.n370 B.n235 256.663
R391 B.n370 B.n236 256.663
R392 B.n370 B.n237 256.663
R393 B.n370 B.n238 256.663
R394 B.n370 B.n239 256.663
R395 B.n370 B.n240 256.663
R396 B.n370 B.n241 256.663
R397 B.n370 B.n242 256.663
R398 B.n370 B.n243 256.663
R399 B.n370 B.n244 256.663
R400 B.n370 B.n245 256.663
R401 B.n370 B.n246 256.663
R402 B.n377 B.n214 163.367
R403 B.n377 B.n212 163.367
R404 B.n381 B.n212 163.367
R405 B.n381 B.n206 163.367
R406 B.n389 B.n206 163.367
R407 B.n389 B.n204 163.367
R408 B.n393 B.n204 163.367
R409 B.n393 B.n198 163.367
R410 B.n402 B.n198 163.367
R411 B.n402 B.n196 163.367
R412 B.n406 B.n196 163.367
R413 B.n406 B.n191 163.367
R414 B.n416 B.n191 163.367
R415 B.n416 B.n189 163.367
R416 B.n420 B.n189 163.367
R417 B.n420 B.n2 163.367
R418 B.n486 B.n2 163.367
R419 B.n486 B.n3 163.367
R420 B.n482 B.n3 163.367
R421 B.n482 B.n8 163.367
R422 B.n478 B.n8 163.367
R423 B.n478 B.n10 163.367
R424 B.n474 B.n10 163.367
R425 B.n474 B.n15 163.367
R426 B.n470 B.n15 163.367
R427 B.n470 B.n17 163.367
R428 B.n466 B.n17 163.367
R429 B.n466 B.n22 163.367
R430 B.n462 B.n22 163.367
R431 B.n462 B.n24 163.367
R432 B.n458 B.n24 163.367
R433 B.n458 B.n29 163.367
R434 B.n454 B.n29 163.367
R435 B.n454 B.n31 163.367
R436 B.n248 B.n247 163.367
R437 B.n363 B.n247 163.367
R438 B.n361 B.n360 163.367
R439 B.n357 B.n356 163.367
R440 B.n353 B.n352 163.367
R441 B.n349 B.n348 163.367
R442 B.n345 B.n344 163.367
R443 B.n341 B.n340 163.367
R444 B.n337 B.n336 163.367
R445 B.n333 B.n332 163.367
R446 B.n329 B.n328 163.367
R447 B.n325 B.n324 163.367
R448 B.n321 B.n320 163.367
R449 B.n317 B.n316 163.367
R450 B.n313 B.n312 163.367
R451 B.n309 B.n308 163.367
R452 B.n305 B.n304 163.367
R453 B.n301 B.n300 163.367
R454 B.n297 B.n296 163.367
R455 B.n293 B.n292 163.367
R456 B.n289 B.n288 163.367
R457 B.n285 B.n284 163.367
R458 B.n281 B.n280 163.367
R459 B.n277 B.n276 163.367
R460 B.n273 B.n272 163.367
R461 B.n269 B.n268 163.367
R462 B.n265 B.n264 163.367
R463 B.n261 B.n260 163.367
R464 B.n257 B.n256 163.367
R465 B.n371 B.n218 163.367
R466 B.n375 B.n216 163.367
R467 B.n375 B.n209 163.367
R468 B.n383 B.n209 163.367
R469 B.n383 B.n207 163.367
R470 B.n387 B.n207 163.367
R471 B.n387 B.n202 163.367
R472 B.n395 B.n202 163.367
R473 B.n395 B.n200 163.367
R474 B.n399 B.n200 163.367
R475 B.n399 B.n194 163.367
R476 B.n408 B.n194 163.367
R477 B.n408 B.n192 163.367
R478 B.n413 B.n192 163.367
R479 B.n413 B.n188 163.367
R480 B.n422 B.n188 163.367
R481 B.n423 B.n422 163.367
R482 B.n423 B.n5 163.367
R483 B.n6 B.n5 163.367
R484 B.n7 B.n6 163.367
R485 B.n428 B.n7 163.367
R486 B.n428 B.n12 163.367
R487 B.n13 B.n12 163.367
R488 B.n14 B.n13 163.367
R489 B.n434 B.n14 163.367
R490 B.n434 B.n18 163.367
R491 B.n19 B.n18 163.367
R492 B.n20 B.n19 163.367
R493 B.n439 B.n20 163.367
R494 B.n439 B.n25 163.367
R495 B.n26 B.n25 163.367
R496 B.n27 B.n26 163.367
R497 B.n444 B.n27 163.367
R498 B.n444 B.n32 163.367
R499 B.n33 B.n32 163.367
R500 B.n72 B.n71 163.367
R501 B.n76 B.n75 163.367
R502 B.n80 B.n79 163.367
R503 B.n84 B.n83 163.367
R504 B.n88 B.n87 163.367
R505 B.n92 B.n91 163.367
R506 B.n96 B.n95 163.367
R507 B.n100 B.n99 163.367
R508 B.n104 B.n103 163.367
R509 B.n108 B.n107 163.367
R510 B.n112 B.n111 163.367
R511 B.n116 B.n115 163.367
R512 B.n121 B.n120 163.367
R513 B.n125 B.n124 163.367
R514 B.n129 B.n128 163.367
R515 B.n133 B.n132 163.367
R516 B.n137 B.n136 163.367
R517 B.n142 B.n141 163.367
R518 B.n146 B.n145 163.367
R519 B.n150 B.n149 163.367
R520 B.n154 B.n153 163.367
R521 B.n158 B.n157 163.367
R522 B.n162 B.n161 163.367
R523 B.n166 B.n165 163.367
R524 B.n170 B.n169 163.367
R525 B.n174 B.n173 163.367
R526 B.n178 B.n177 163.367
R527 B.n182 B.n181 163.367
R528 B.n184 B.n63 163.367
R529 B.n370 B.n215 112.121
R530 B.n452 B.n451 112.121
R531 B.n252 B.t11 86.3035
R532 B.n64 B.t14 86.3035
R533 B.n249 B.t21 86.2968
R534 B.n66 B.t17 86.2968
R535 B.n253 B.t10 74.6672
R536 B.n65 B.t15 74.6672
R537 B.n250 B.t20 74.6604
R538 B.n67 B.t18 74.6604
R539 B.n369 B.n368 71.676
R540 B.n363 B.n219 71.676
R541 B.n360 B.n220 71.676
R542 B.n356 B.n221 71.676
R543 B.n352 B.n222 71.676
R544 B.n348 B.n223 71.676
R545 B.n344 B.n224 71.676
R546 B.n340 B.n225 71.676
R547 B.n336 B.n226 71.676
R548 B.n332 B.n227 71.676
R549 B.n328 B.n228 71.676
R550 B.n324 B.n229 71.676
R551 B.n320 B.n230 71.676
R552 B.n316 B.n231 71.676
R553 B.n312 B.n232 71.676
R554 B.n308 B.n233 71.676
R555 B.n304 B.n234 71.676
R556 B.n300 B.n235 71.676
R557 B.n296 B.n236 71.676
R558 B.n292 B.n237 71.676
R559 B.n288 B.n238 71.676
R560 B.n284 B.n239 71.676
R561 B.n280 B.n240 71.676
R562 B.n276 B.n241 71.676
R563 B.n272 B.n242 71.676
R564 B.n268 B.n243 71.676
R565 B.n264 B.n244 71.676
R566 B.n260 B.n245 71.676
R567 B.n256 B.n246 71.676
R568 B.n68 B.n34 71.676
R569 B.n72 B.n35 71.676
R570 B.n76 B.n36 71.676
R571 B.n80 B.n37 71.676
R572 B.n84 B.n38 71.676
R573 B.n88 B.n39 71.676
R574 B.n92 B.n40 71.676
R575 B.n96 B.n41 71.676
R576 B.n100 B.n42 71.676
R577 B.n104 B.n43 71.676
R578 B.n108 B.n44 71.676
R579 B.n112 B.n45 71.676
R580 B.n116 B.n46 71.676
R581 B.n121 B.n47 71.676
R582 B.n125 B.n48 71.676
R583 B.n129 B.n49 71.676
R584 B.n133 B.n50 71.676
R585 B.n137 B.n51 71.676
R586 B.n142 B.n52 71.676
R587 B.n146 B.n53 71.676
R588 B.n150 B.n54 71.676
R589 B.n154 B.n55 71.676
R590 B.n158 B.n56 71.676
R591 B.n162 B.n57 71.676
R592 B.n166 B.n58 71.676
R593 B.n170 B.n59 71.676
R594 B.n174 B.n60 71.676
R595 B.n178 B.n61 71.676
R596 B.n182 B.n62 71.676
R597 B.n450 B.n63 71.676
R598 B.n450 B.n449 71.676
R599 B.n184 B.n62 71.676
R600 B.n181 B.n61 71.676
R601 B.n177 B.n60 71.676
R602 B.n173 B.n59 71.676
R603 B.n169 B.n58 71.676
R604 B.n165 B.n57 71.676
R605 B.n161 B.n56 71.676
R606 B.n157 B.n55 71.676
R607 B.n153 B.n54 71.676
R608 B.n149 B.n53 71.676
R609 B.n145 B.n52 71.676
R610 B.n141 B.n51 71.676
R611 B.n136 B.n50 71.676
R612 B.n132 B.n49 71.676
R613 B.n128 B.n48 71.676
R614 B.n124 B.n47 71.676
R615 B.n120 B.n46 71.676
R616 B.n115 B.n45 71.676
R617 B.n111 B.n44 71.676
R618 B.n107 B.n43 71.676
R619 B.n103 B.n42 71.676
R620 B.n99 B.n41 71.676
R621 B.n95 B.n40 71.676
R622 B.n91 B.n39 71.676
R623 B.n87 B.n38 71.676
R624 B.n83 B.n37 71.676
R625 B.n79 B.n36 71.676
R626 B.n75 B.n35 71.676
R627 B.n71 B.n34 71.676
R628 B.n369 B.n248 71.676
R629 B.n361 B.n219 71.676
R630 B.n357 B.n220 71.676
R631 B.n353 B.n221 71.676
R632 B.n349 B.n222 71.676
R633 B.n345 B.n223 71.676
R634 B.n341 B.n224 71.676
R635 B.n337 B.n225 71.676
R636 B.n333 B.n226 71.676
R637 B.n329 B.n227 71.676
R638 B.n325 B.n228 71.676
R639 B.n321 B.n229 71.676
R640 B.n317 B.n230 71.676
R641 B.n313 B.n231 71.676
R642 B.n309 B.n232 71.676
R643 B.n305 B.n233 71.676
R644 B.n301 B.n234 71.676
R645 B.n297 B.n235 71.676
R646 B.n293 B.n236 71.676
R647 B.n289 B.n237 71.676
R648 B.n285 B.n238 71.676
R649 B.n281 B.n239 71.676
R650 B.n277 B.n240 71.676
R651 B.n273 B.n241 71.676
R652 B.n269 B.n242 71.676
R653 B.n265 B.n243 71.676
R654 B.n261 B.n244 71.676
R655 B.n257 B.n245 71.676
R656 B.n246 B.n218 71.676
R657 B.n376 B.n215 64.069
R658 B.n376 B.n210 64.069
R659 B.n382 B.n210 64.069
R660 B.n382 B.n211 64.069
R661 B.n388 B.n203 64.069
R662 B.n394 B.n203 64.069
R663 B.n394 B.n199 64.069
R664 B.n401 B.n199 64.069
R665 B.n407 B.n195 64.069
R666 B.n415 B.n414 64.069
R667 B.n421 B.n4 64.069
R668 B.n485 B.n4 64.069
R669 B.n485 B.n484 64.069
R670 B.n484 B.n483 64.069
R671 B.n477 B.n11 64.069
R672 B.n476 B.n475 64.069
R673 B.n469 B.n468 64.069
R674 B.n468 B.n467 64.069
R675 B.n467 B.n21 64.069
R676 B.n461 B.n21 64.069
R677 B.n460 B.n459 64.069
R678 B.n459 B.n28 64.069
R679 B.n453 B.n28 64.069
R680 B.n453 B.n452 64.069
R681 B.n400 B.t1 63.1268
R682 B.n433 B.t7 63.1268
R683 B.n254 B.n253 59.5399
R684 B.n251 B.n250 59.5399
R685 B.n118 B.n67 59.5399
R686 B.n139 B.n65 59.5399
R687 B.t6 B.n400 49.9363
R688 B.n433 B.t0 49.9363
R689 B.n388 B.t9 48.0519
R690 B.n195 B.t4 48.0519
R691 B.t5 B.n476 48.0519
R692 B.n461 B.t13 48.0519
R693 B.n414 B.t2 32.9769
R694 B.n11 B.t3 32.9769
R695 B.n421 B.t2 31.0926
R696 B.n483 B.t3 31.0926
R697 B.n69 B.n30 31.0639
R698 B.n448 B.n447 31.0639
R699 B.n373 B.n372 31.0639
R700 B.n367 B.n213 31.0639
R701 B B.n487 18.0485
R702 B.n211 B.t9 16.0176
R703 B.n415 B.t4 16.0176
R704 B.n477 B.t5 16.0176
R705 B.t13 B.n460 16.0176
R706 B.n401 B.t6 14.1333
R707 B.n469 B.t0 14.1333
R708 B.n253 B.n252 11.6369
R709 B.n250 B.n249 11.6369
R710 B.n67 B.n66 11.6369
R711 B.n65 B.n64 11.6369
R712 B.n70 B.n69 10.6151
R713 B.n73 B.n70 10.6151
R714 B.n74 B.n73 10.6151
R715 B.n77 B.n74 10.6151
R716 B.n78 B.n77 10.6151
R717 B.n81 B.n78 10.6151
R718 B.n82 B.n81 10.6151
R719 B.n85 B.n82 10.6151
R720 B.n86 B.n85 10.6151
R721 B.n89 B.n86 10.6151
R722 B.n90 B.n89 10.6151
R723 B.n93 B.n90 10.6151
R724 B.n94 B.n93 10.6151
R725 B.n97 B.n94 10.6151
R726 B.n98 B.n97 10.6151
R727 B.n101 B.n98 10.6151
R728 B.n102 B.n101 10.6151
R729 B.n105 B.n102 10.6151
R730 B.n106 B.n105 10.6151
R731 B.n109 B.n106 10.6151
R732 B.n110 B.n109 10.6151
R733 B.n113 B.n110 10.6151
R734 B.n114 B.n113 10.6151
R735 B.n117 B.n114 10.6151
R736 B.n122 B.n119 10.6151
R737 B.n123 B.n122 10.6151
R738 B.n126 B.n123 10.6151
R739 B.n127 B.n126 10.6151
R740 B.n130 B.n127 10.6151
R741 B.n131 B.n130 10.6151
R742 B.n134 B.n131 10.6151
R743 B.n135 B.n134 10.6151
R744 B.n138 B.n135 10.6151
R745 B.n143 B.n140 10.6151
R746 B.n144 B.n143 10.6151
R747 B.n147 B.n144 10.6151
R748 B.n148 B.n147 10.6151
R749 B.n151 B.n148 10.6151
R750 B.n152 B.n151 10.6151
R751 B.n155 B.n152 10.6151
R752 B.n156 B.n155 10.6151
R753 B.n159 B.n156 10.6151
R754 B.n160 B.n159 10.6151
R755 B.n163 B.n160 10.6151
R756 B.n164 B.n163 10.6151
R757 B.n167 B.n164 10.6151
R758 B.n168 B.n167 10.6151
R759 B.n171 B.n168 10.6151
R760 B.n172 B.n171 10.6151
R761 B.n175 B.n172 10.6151
R762 B.n176 B.n175 10.6151
R763 B.n179 B.n176 10.6151
R764 B.n180 B.n179 10.6151
R765 B.n183 B.n180 10.6151
R766 B.n185 B.n183 10.6151
R767 B.n186 B.n185 10.6151
R768 B.n448 B.n186 10.6151
R769 B.n374 B.n373 10.6151
R770 B.n374 B.n208 10.6151
R771 B.n384 B.n208 10.6151
R772 B.n385 B.n384 10.6151
R773 B.n386 B.n385 10.6151
R774 B.n386 B.n201 10.6151
R775 B.n396 B.n201 10.6151
R776 B.n397 B.n396 10.6151
R777 B.n398 B.n397 10.6151
R778 B.n398 B.n193 10.6151
R779 B.n409 B.n193 10.6151
R780 B.n410 B.n409 10.6151
R781 B.n412 B.n410 10.6151
R782 B.n412 B.n411 10.6151
R783 B.n411 B.n187 10.6151
R784 B.n424 B.n187 10.6151
R785 B.n425 B.n424 10.6151
R786 B.n426 B.n425 10.6151
R787 B.n427 B.n426 10.6151
R788 B.n429 B.n427 10.6151
R789 B.n430 B.n429 10.6151
R790 B.n431 B.n430 10.6151
R791 B.n432 B.n431 10.6151
R792 B.n435 B.n432 10.6151
R793 B.n436 B.n435 10.6151
R794 B.n437 B.n436 10.6151
R795 B.n438 B.n437 10.6151
R796 B.n440 B.n438 10.6151
R797 B.n441 B.n440 10.6151
R798 B.n442 B.n441 10.6151
R799 B.n443 B.n442 10.6151
R800 B.n445 B.n443 10.6151
R801 B.n446 B.n445 10.6151
R802 B.n447 B.n446 10.6151
R803 B.n367 B.n366 10.6151
R804 B.n366 B.n365 10.6151
R805 B.n365 B.n364 10.6151
R806 B.n364 B.n362 10.6151
R807 B.n362 B.n359 10.6151
R808 B.n359 B.n358 10.6151
R809 B.n358 B.n355 10.6151
R810 B.n355 B.n354 10.6151
R811 B.n354 B.n351 10.6151
R812 B.n351 B.n350 10.6151
R813 B.n350 B.n347 10.6151
R814 B.n347 B.n346 10.6151
R815 B.n346 B.n343 10.6151
R816 B.n343 B.n342 10.6151
R817 B.n342 B.n339 10.6151
R818 B.n339 B.n338 10.6151
R819 B.n338 B.n335 10.6151
R820 B.n335 B.n334 10.6151
R821 B.n334 B.n331 10.6151
R822 B.n331 B.n330 10.6151
R823 B.n330 B.n327 10.6151
R824 B.n327 B.n326 10.6151
R825 B.n326 B.n323 10.6151
R826 B.n323 B.n322 10.6151
R827 B.n319 B.n318 10.6151
R828 B.n318 B.n315 10.6151
R829 B.n315 B.n314 10.6151
R830 B.n314 B.n311 10.6151
R831 B.n311 B.n310 10.6151
R832 B.n310 B.n307 10.6151
R833 B.n307 B.n306 10.6151
R834 B.n306 B.n303 10.6151
R835 B.n303 B.n302 10.6151
R836 B.n299 B.n298 10.6151
R837 B.n298 B.n295 10.6151
R838 B.n295 B.n294 10.6151
R839 B.n294 B.n291 10.6151
R840 B.n291 B.n290 10.6151
R841 B.n290 B.n287 10.6151
R842 B.n287 B.n286 10.6151
R843 B.n286 B.n283 10.6151
R844 B.n283 B.n282 10.6151
R845 B.n282 B.n279 10.6151
R846 B.n279 B.n278 10.6151
R847 B.n278 B.n275 10.6151
R848 B.n275 B.n274 10.6151
R849 B.n274 B.n271 10.6151
R850 B.n271 B.n270 10.6151
R851 B.n270 B.n267 10.6151
R852 B.n267 B.n266 10.6151
R853 B.n266 B.n263 10.6151
R854 B.n263 B.n262 10.6151
R855 B.n262 B.n259 10.6151
R856 B.n259 B.n258 10.6151
R857 B.n258 B.n255 10.6151
R858 B.n255 B.n217 10.6151
R859 B.n372 B.n217 10.6151
R860 B.n378 B.n213 10.6151
R861 B.n379 B.n378 10.6151
R862 B.n380 B.n379 10.6151
R863 B.n380 B.n205 10.6151
R864 B.n390 B.n205 10.6151
R865 B.n391 B.n390 10.6151
R866 B.n392 B.n391 10.6151
R867 B.n392 B.n197 10.6151
R868 B.n403 B.n197 10.6151
R869 B.n404 B.n403 10.6151
R870 B.n405 B.n404 10.6151
R871 B.n405 B.n190 10.6151
R872 B.n417 B.n190 10.6151
R873 B.n418 B.n417 10.6151
R874 B.n419 B.n418 10.6151
R875 B.n419 B.n0 10.6151
R876 B.n481 B.n1 10.6151
R877 B.n481 B.n480 10.6151
R878 B.n480 B.n479 10.6151
R879 B.n479 B.n9 10.6151
R880 B.n473 B.n9 10.6151
R881 B.n473 B.n472 10.6151
R882 B.n472 B.n471 10.6151
R883 B.n471 B.n16 10.6151
R884 B.n465 B.n16 10.6151
R885 B.n465 B.n464 10.6151
R886 B.n464 B.n463 10.6151
R887 B.n463 B.n23 10.6151
R888 B.n457 B.n23 10.6151
R889 B.n457 B.n456 10.6151
R890 B.n456 B.n455 10.6151
R891 B.n455 B.n30 10.6151
R892 B.n118 B.n117 9.36635
R893 B.n140 B.n139 9.36635
R894 B.n322 B.n251 9.36635
R895 B.n299 B.n254 9.36635
R896 B.n487 B.n0 2.81026
R897 B.n487 B.n1 2.81026
R898 B.n119 B.n118 1.24928
R899 B.n139 B.n138 1.24928
R900 B.n319 B.n251 1.24928
R901 B.n302 B.n254 1.24928
R902 B.n407 B.t1 0.942684
R903 B.n475 B.t7 0.942684
R904 VP.n13 VP.t6 745.721
R905 VP.n9 VP.t2 745.721
R906 VP.n2 VP.t7 745.721
R907 VP.n6 VP.t5 745.721
R908 VP.n12 VP.t0 687.297
R909 VP.n10 VP.t4 687.297
R910 VP.n3 VP.t1 687.297
R911 VP.n5 VP.t3 687.297
R912 VP.n2 VP.n1 161.489
R913 VP.n14 VP.n13 161.3
R914 VP.n4 VP.n1 161.3
R915 VP.n7 VP.n6 161.3
R916 VP.n11 VP.n0 161.3
R917 VP.n9 VP.n8 161.3
R918 VP.n11 VP.n10 43.8187
R919 VP.n12 VP.n11 43.8187
R920 VP.n4 VP.n3 43.8187
R921 VP.n5 VP.n4 43.8187
R922 VP.n8 VP.n7 35.902
R923 VP.n10 VP.n9 29.2126
R924 VP.n13 VP.n12 29.2126
R925 VP.n3 VP.n2 29.2126
R926 VP.n6 VP.n5 29.2126
R927 VP.n7 VP.n1 0.189894
R928 VP.n8 VP.n0 0.189894
R929 VP.n14 VP.n0 0.189894
R930 VP VP.n14 0.0516364
R931 VDD1 VDD1.n0 67.6886
R932 VDD1.n3 VDD1.n2 67.5749
R933 VDD1.n3 VDD1.n1 67.5749
R934 VDD1.n5 VDD1.n4 67.3716
R935 VDD1.n5 VDD1.n3 32.1431
R936 VDD1.n4 VDD1.t4 3.09425
R937 VDD1.n4 VDD1.t2 3.09425
R938 VDD1.n0 VDD1.t0 3.09425
R939 VDD1.n0 VDD1.t6 3.09425
R940 VDD1.n2 VDD1.t7 3.09425
R941 VDD1.n2 VDD1.t1 3.09425
R942 VDD1.n1 VDD1.t5 3.09425
R943 VDD1.n1 VDD1.t3 3.09425
R944 VDD1 VDD1.n5 0.200931
C0 VTAIL VDD2 10.029901f
C1 VDD1 VN 0.14763f
C2 VP VN 3.76971f
C3 VDD1 VDD2 0.616831f
C4 VP VDD2 0.271849f
C5 VTAIL VDD1 9.99115f
C6 VTAIL VP 1.6825f
C7 VP VDD1 1.95732f
C8 VN VDD2 1.83332f
C9 VTAIL VN 1.6684f
C10 VDD2 B 2.605263f
C11 VDD1 B 2.775693f
C12 VTAIL B 5.297028f
C13 VN B 5.527513f
C14 VP B 4.497422f
C15 VDD1.t0 B 0.1413f
C16 VDD1.t6 B 0.1413f
C17 VDD1.n0 B 1.18929f
C18 VDD1.t5 B 0.1413f
C19 VDD1.t3 B 0.1413f
C20 VDD1.n1 B 1.18874f
C21 VDD1.t7 B 0.1413f
C22 VDD1.t1 B 0.1413f
C23 VDD1.n2 B 1.18874f
C24 VDD1.n3 B 1.82993f
C25 VDD1.t4 B 0.1413f
C26 VDD1.t2 B 0.1413f
C27 VDD1.n4 B 1.18781f
C28 VDD1.n5 B 1.92589f
C29 VP.n0 B 0.029597f
C30 VP.t0 B 0.145569f
C31 VP.t4 B 0.145569f
C32 VP.t2 B 0.15103f
C33 VP.n1 B 0.069549f
C34 VP.t3 B 0.145569f
C35 VP.t1 B 0.145569f
C36 VP.t7 B 0.15103f
C37 VP.n2 B 0.075936f
C38 VP.n3 B 0.066605f
C39 VP.n4 B 0.011643f
C40 VP.n5 B 0.066605f
C41 VP.t5 B 0.15103f
C42 VP.n6 B 0.075889f
C43 VP.n7 B 0.925717f
C44 VP.n8 B 0.955437f
C45 VP.n9 B 0.075889f
C46 VP.n10 B 0.066605f
C47 VP.n11 B 0.011643f
C48 VP.n12 B 0.066605f
C49 VP.t6 B 0.15103f
C50 VP.n13 B 0.075889f
C51 VP.n14 B 0.022937f
C52 VDD2.t2 B 0.142774f
C53 VDD2.t4 B 0.142774f
C54 VDD2.n0 B 1.20113f
C55 VDD2.t0 B 0.142774f
C56 VDD2.t6 B 0.142774f
C57 VDD2.n1 B 1.20113f
C58 VDD2.n2 B 1.7881f
C59 VDD2.t5 B 0.142774f
C60 VDD2.t7 B 0.142774f
C61 VDD2.n3 B 1.2002f
C62 VDD2.n4 B 1.9132f
C63 VDD2.t1 B 0.142774f
C64 VDD2.t3 B 0.142774f
C65 VDD2.n5 B 1.20111f
C66 VTAIL.t12 B 0.11148f
C67 VTAIL.t15 B 0.11148f
C68 VTAIL.n0 B 0.879386f
C69 VTAIL.n1 B 0.248359f
C70 VTAIL.t8 B 1.12176f
C71 VTAIL.n2 B 0.339254f
C72 VTAIL.t2 B 1.12176f
C73 VTAIL.n3 B 0.339254f
C74 VTAIL.t1 B 0.11148f
C75 VTAIL.t4 B 0.11148f
C76 VTAIL.n4 B 0.879386f
C77 VTAIL.n5 B 0.280963f
C78 VTAIL.t6 B 1.12176f
C79 VTAIL.n6 B 1.03391f
C80 VTAIL.t10 B 1.12177f
C81 VTAIL.n7 B 1.03391f
C82 VTAIL.t11 B 0.11148f
C83 VTAIL.t14 B 0.11148f
C84 VTAIL.n8 B 0.879391f
C85 VTAIL.n9 B 0.280959f
C86 VTAIL.t13 B 1.12177f
C87 VTAIL.n10 B 0.339248f
C88 VTAIL.t3 B 1.12177f
C89 VTAIL.n11 B 0.339248f
C90 VTAIL.t5 B 0.11148f
C91 VTAIL.t7 B 0.11148f
C92 VTAIL.n12 B 0.879391f
C93 VTAIL.n13 B 0.280959f
C94 VTAIL.t0 B 1.12176f
C95 VTAIL.n14 B 1.03391f
C96 VTAIL.t9 B 1.12176f
C97 VTAIL.n15 B 1.02978f
C98 VN.n0 B 0.068795f
C99 VN.t7 B 0.143992f
C100 VN.t3 B 0.143992f
C101 VN.t5 B 0.149394f
C102 VN.n1 B 0.075113f
C103 VN.n2 B 0.065884f
C104 VN.n3 B 0.011517f
C105 VN.n4 B 0.065884f
C106 VN.t1 B 0.149394f
C107 VN.n5 B 0.075067f
C108 VN.n6 B 0.022688f
C109 VN.n7 B 0.068795f
C110 VN.t2 B 0.149394f
C111 VN.t0 B 0.143992f
C112 VN.t6 B 0.143992f
C113 VN.t4 B 0.149394f
C114 VN.n8 B 0.075113f
C115 VN.n9 B 0.065884f
C116 VN.n10 B 0.011517f
C117 VN.n11 B 0.065884f
C118 VN.n12 B 0.075067f
C119 VN.n13 B 0.935115f
.ends

