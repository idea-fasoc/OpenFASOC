* NGSPICE file created from diff_pair_sample_1172.ext - technology: sky130A

.subckt diff_pair_sample_1172 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X1 VTAIL.t11 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X2 VDD1.t7 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=2.1138 ps=11.62 w=5.42 l=2.37
X3 VTAIL.t3 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X4 VDD2.t5 VN.t2 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=2.1138 ps=11.62 w=5.42 l=2.37
X5 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X6 VTAIL.t12 VN.t3 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0.8943 ps=5.75 w=5.42 l=2.37
X7 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0 ps=0 w=5.42 l=2.37
X8 VTAIL.t5 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0.8943 ps=5.75 w=5.42 l=2.37
X9 VTAIL.t13 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0.8943 ps=5.75 w=5.42 l=2.37
X10 VTAIL.t6 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X11 VDD2.t1 VN.t6 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=2.1138 ps=11.62 w=5.42 l=2.37
X12 VTAIL.t15 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X13 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0 ps=0 w=5.42 l=2.37
X14 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0 ps=0 w=5.42 l=2.37
X15 VDD1.t2 VP.t5 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=2.1138 ps=11.62 w=5.42 l=2.37
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0 ps=0 w=5.42 l=2.37
X17 VDD1.t1 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X18 VDD2.t0 VN.t7 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8943 pd=5.75 as=0.8943 ps=5.75 w=5.42 l=2.37
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1138 pd=11.62 as=0.8943 ps=5.75 w=5.42 l=2.37
R0 VN.n51 VN.n27 161.3
R1 VN.n50 VN.n49 161.3
R2 VN.n48 VN.n28 161.3
R3 VN.n47 VN.n46 161.3
R4 VN.n45 VN.n29 161.3
R5 VN.n43 VN.n42 161.3
R6 VN.n41 VN.n30 161.3
R7 VN.n40 VN.n39 161.3
R8 VN.n38 VN.n31 161.3
R9 VN.n37 VN.n36 161.3
R10 VN.n35 VN.n32 161.3
R11 VN.n24 VN.n0 161.3
R12 VN.n23 VN.n22 161.3
R13 VN.n21 VN.n1 161.3
R14 VN.n20 VN.n19 161.3
R15 VN.n18 VN.n2 161.3
R16 VN.n16 VN.n15 161.3
R17 VN.n14 VN.n3 161.3
R18 VN.n13 VN.n12 161.3
R19 VN.n11 VN.n4 161.3
R20 VN.n10 VN.n9 161.3
R21 VN.n8 VN.n5 161.3
R22 VN.n26 VN.n25 96.1531
R23 VN.n53 VN.n52 96.1531
R24 VN.n7 VN.t4 87.6179
R25 VN.n34 VN.t6 87.6179
R26 VN.n7 VN.n6 67.4531
R27 VN.n34 VN.n33 67.4531
R28 VN.n12 VN.n11 56.5617
R29 VN.n39 VN.n38 56.5617
R30 VN.n6 VN.t0 55.1153
R31 VN.n17 VN.t5 55.1153
R32 VN.n25 VN.t2 55.1153
R33 VN.n33 VN.t1 55.1153
R34 VN.n44 VN.t7 55.1153
R35 VN.n52 VN.t3 55.1153
R36 VN.n19 VN.n1 45.4209
R37 VN.n46 VN.n28 45.4209
R38 VN VN.n53 45.1497
R39 VN.n23 VN.n1 35.7332
R40 VN.n50 VN.n28 35.7332
R41 VN.n10 VN.n5 24.5923
R42 VN.n11 VN.n10 24.5923
R43 VN.n12 VN.n3 24.5923
R44 VN.n16 VN.n3 24.5923
R45 VN.n19 VN.n18 24.5923
R46 VN.n24 VN.n23 24.5923
R47 VN.n38 VN.n37 24.5923
R48 VN.n37 VN.n32 24.5923
R49 VN.n46 VN.n45 24.5923
R50 VN.n43 VN.n30 24.5923
R51 VN.n39 VN.n30 24.5923
R52 VN.n51 VN.n50 24.5923
R53 VN.n18 VN.n17 19.674
R54 VN.n45 VN.n44 19.674
R55 VN.n25 VN.n24 14.7556
R56 VN.n52 VN.n51 14.7556
R57 VN.n35 VN.n34 9.50446
R58 VN.n8 VN.n7 9.50446
R59 VN.n6 VN.n5 4.91887
R60 VN.n17 VN.n16 4.91887
R61 VN.n33 VN.n32 4.91887
R62 VN.n44 VN.n43 4.91887
R63 VN.n53 VN.n27 0.278335
R64 VN.n26 VN.n0 0.278335
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n42 VN.n29 0.189894
R70 VN.n42 VN.n41 0.189894
R71 VN.n41 VN.n40 0.189894
R72 VN.n40 VN.n31 0.189894
R73 VN.n36 VN.n31 0.189894
R74 VN.n36 VN.n35 0.189894
R75 VN.n9 VN.n8 0.189894
R76 VN.n9 VN.n4 0.189894
R77 VN.n13 VN.n4 0.189894
R78 VN.n14 VN.n13 0.189894
R79 VN.n15 VN.n14 0.189894
R80 VN.n15 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153485
R86 VTAIL.n226 VTAIL.n204 289.615
R87 VTAIL.n24 VTAIL.n2 289.615
R88 VTAIL.n52 VTAIL.n30 289.615
R89 VTAIL.n82 VTAIL.n60 289.615
R90 VTAIL.n198 VTAIL.n176 289.615
R91 VTAIL.n168 VTAIL.n146 289.615
R92 VTAIL.n140 VTAIL.n118 289.615
R93 VTAIL.n110 VTAIL.n88 289.615
R94 VTAIL.n212 VTAIL.n211 185
R95 VTAIL.n217 VTAIL.n216 185
R96 VTAIL.n219 VTAIL.n218 185
R97 VTAIL.n208 VTAIL.n207 185
R98 VTAIL.n225 VTAIL.n224 185
R99 VTAIL.n227 VTAIL.n226 185
R100 VTAIL.n10 VTAIL.n9 185
R101 VTAIL.n15 VTAIL.n14 185
R102 VTAIL.n17 VTAIL.n16 185
R103 VTAIL.n6 VTAIL.n5 185
R104 VTAIL.n23 VTAIL.n22 185
R105 VTAIL.n25 VTAIL.n24 185
R106 VTAIL.n38 VTAIL.n37 185
R107 VTAIL.n43 VTAIL.n42 185
R108 VTAIL.n45 VTAIL.n44 185
R109 VTAIL.n34 VTAIL.n33 185
R110 VTAIL.n51 VTAIL.n50 185
R111 VTAIL.n53 VTAIL.n52 185
R112 VTAIL.n68 VTAIL.n67 185
R113 VTAIL.n73 VTAIL.n72 185
R114 VTAIL.n75 VTAIL.n74 185
R115 VTAIL.n64 VTAIL.n63 185
R116 VTAIL.n81 VTAIL.n80 185
R117 VTAIL.n83 VTAIL.n82 185
R118 VTAIL.n199 VTAIL.n198 185
R119 VTAIL.n197 VTAIL.n196 185
R120 VTAIL.n180 VTAIL.n179 185
R121 VTAIL.n191 VTAIL.n190 185
R122 VTAIL.n189 VTAIL.n188 185
R123 VTAIL.n184 VTAIL.n183 185
R124 VTAIL.n169 VTAIL.n168 185
R125 VTAIL.n167 VTAIL.n166 185
R126 VTAIL.n150 VTAIL.n149 185
R127 VTAIL.n161 VTAIL.n160 185
R128 VTAIL.n159 VTAIL.n158 185
R129 VTAIL.n154 VTAIL.n153 185
R130 VTAIL.n141 VTAIL.n140 185
R131 VTAIL.n139 VTAIL.n138 185
R132 VTAIL.n122 VTAIL.n121 185
R133 VTAIL.n133 VTAIL.n132 185
R134 VTAIL.n131 VTAIL.n130 185
R135 VTAIL.n126 VTAIL.n125 185
R136 VTAIL.n111 VTAIL.n110 185
R137 VTAIL.n109 VTAIL.n108 185
R138 VTAIL.n92 VTAIL.n91 185
R139 VTAIL.n103 VTAIL.n102 185
R140 VTAIL.n101 VTAIL.n100 185
R141 VTAIL.n96 VTAIL.n95 185
R142 VTAIL.n213 VTAIL.t8 147.672
R143 VTAIL.n11 VTAIL.t5 147.672
R144 VTAIL.n39 VTAIL.t4 147.672
R145 VTAIL.n69 VTAIL.t0 147.672
R146 VTAIL.n185 VTAIL.t14 147.672
R147 VTAIL.n155 VTAIL.t13 147.672
R148 VTAIL.n127 VTAIL.t7 147.672
R149 VTAIL.n97 VTAIL.t12 147.672
R150 VTAIL.n217 VTAIL.n211 104.615
R151 VTAIL.n218 VTAIL.n217 104.615
R152 VTAIL.n218 VTAIL.n207 104.615
R153 VTAIL.n225 VTAIL.n207 104.615
R154 VTAIL.n226 VTAIL.n225 104.615
R155 VTAIL.n15 VTAIL.n9 104.615
R156 VTAIL.n16 VTAIL.n15 104.615
R157 VTAIL.n16 VTAIL.n5 104.615
R158 VTAIL.n23 VTAIL.n5 104.615
R159 VTAIL.n24 VTAIL.n23 104.615
R160 VTAIL.n43 VTAIL.n37 104.615
R161 VTAIL.n44 VTAIL.n43 104.615
R162 VTAIL.n44 VTAIL.n33 104.615
R163 VTAIL.n51 VTAIL.n33 104.615
R164 VTAIL.n52 VTAIL.n51 104.615
R165 VTAIL.n73 VTAIL.n67 104.615
R166 VTAIL.n74 VTAIL.n73 104.615
R167 VTAIL.n74 VTAIL.n63 104.615
R168 VTAIL.n81 VTAIL.n63 104.615
R169 VTAIL.n82 VTAIL.n81 104.615
R170 VTAIL.n198 VTAIL.n197 104.615
R171 VTAIL.n197 VTAIL.n179 104.615
R172 VTAIL.n190 VTAIL.n179 104.615
R173 VTAIL.n190 VTAIL.n189 104.615
R174 VTAIL.n189 VTAIL.n183 104.615
R175 VTAIL.n168 VTAIL.n167 104.615
R176 VTAIL.n167 VTAIL.n149 104.615
R177 VTAIL.n160 VTAIL.n149 104.615
R178 VTAIL.n160 VTAIL.n159 104.615
R179 VTAIL.n159 VTAIL.n153 104.615
R180 VTAIL.n140 VTAIL.n139 104.615
R181 VTAIL.n139 VTAIL.n121 104.615
R182 VTAIL.n132 VTAIL.n121 104.615
R183 VTAIL.n132 VTAIL.n131 104.615
R184 VTAIL.n131 VTAIL.n125 104.615
R185 VTAIL.n110 VTAIL.n109 104.615
R186 VTAIL.n109 VTAIL.n91 104.615
R187 VTAIL.n102 VTAIL.n91 104.615
R188 VTAIL.n102 VTAIL.n101 104.615
R189 VTAIL.n101 VTAIL.n95 104.615
R190 VTAIL.n175 VTAIL.n174 54.6916
R191 VTAIL.n117 VTAIL.n116 54.6916
R192 VTAIL.n1 VTAIL.n0 54.6915
R193 VTAIL.n59 VTAIL.n58 54.6915
R194 VTAIL.t8 VTAIL.n211 52.3082
R195 VTAIL.t5 VTAIL.n9 52.3082
R196 VTAIL.t4 VTAIL.n37 52.3082
R197 VTAIL.t0 VTAIL.n67 52.3082
R198 VTAIL.t14 VTAIL.n183 52.3082
R199 VTAIL.t13 VTAIL.n153 52.3082
R200 VTAIL.t7 VTAIL.n125 52.3082
R201 VTAIL.t12 VTAIL.n95 52.3082
R202 VTAIL.n231 VTAIL.n230 34.9005
R203 VTAIL.n29 VTAIL.n28 34.9005
R204 VTAIL.n57 VTAIL.n56 34.9005
R205 VTAIL.n87 VTAIL.n86 34.9005
R206 VTAIL.n203 VTAIL.n202 34.9005
R207 VTAIL.n173 VTAIL.n172 34.9005
R208 VTAIL.n145 VTAIL.n144 34.9005
R209 VTAIL.n115 VTAIL.n114 34.9005
R210 VTAIL.n231 VTAIL.n203 19.3669
R211 VTAIL.n115 VTAIL.n87 19.3669
R212 VTAIL.n213 VTAIL.n212 15.6666
R213 VTAIL.n11 VTAIL.n10 15.6666
R214 VTAIL.n39 VTAIL.n38 15.6666
R215 VTAIL.n69 VTAIL.n68 15.6666
R216 VTAIL.n185 VTAIL.n184 15.6666
R217 VTAIL.n155 VTAIL.n154 15.6666
R218 VTAIL.n127 VTAIL.n126 15.6666
R219 VTAIL.n97 VTAIL.n96 15.6666
R220 VTAIL.n216 VTAIL.n215 12.8005
R221 VTAIL.n14 VTAIL.n13 12.8005
R222 VTAIL.n42 VTAIL.n41 12.8005
R223 VTAIL.n72 VTAIL.n71 12.8005
R224 VTAIL.n188 VTAIL.n187 12.8005
R225 VTAIL.n158 VTAIL.n157 12.8005
R226 VTAIL.n130 VTAIL.n129 12.8005
R227 VTAIL.n100 VTAIL.n99 12.8005
R228 VTAIL.n219 VTAIL.n210 12.0247
R229 VTAIL.n17 VTAIL.n8 12.0247
R230 VTAIL.n45 VTAIL.n36 12.0247
R231 VTAIL.n75 VTAIL.n66 12.0247
R232 VTAIL.n191 VTAIL.n182 12.0247
R233 VTAIL.n161 VTAIL.n152 12.0247
R234 VTAIL.n133 VTAIL.n124 12.0247
R235 VTAIL.n103 VTAIL.n94 12.0247
R236 VTAIL.n220 VTAIL.n208 11.249
R237 VTAIL.n18 VTAIL.n6 11.249
R238 VTAIL.n46 VTAIL.n34 11.249
R239 VTAIL.n76 VTAIL.n64 11.249
R240 VTAIL.n192 VTAIL.n180 11.249
R241 VTAIL.n162 VTAIL.n150 11.249
R242 VTAIL.n134 VTAIL.n122 11.249
R243 VTAIL.n104 VTAIL.n92 11.249
R244 VTAIL.n224 VTAIL.n223 10.4732
R245 VTAIL.n22 VTAIL.n21 10.4732
R246 VTAIL.n50 VTAIL.n49 10.4732
R247 VTAIL.n80 VTAIL.n79 10.4732
R248 VTAIL.n196 VTAIL.n195 10.4732
R249 VTAIL.n166 VTAIL.n165 10.4732
R250 VTAIL.n138 VTAIL.n137 10.4732
R251 VTAIL.n108 VTAIL.n107 10.4732
R252 VTAIL.n227 VTAIL.n206 9.69747
R253 VTAIL.n25 VTAIL.n4 9.69747
R254 VTAIL.n53 VTAIL.n32 9.69747
R255 VTAIL.n83 VTAIL.n62 9.69747
R256 VTAIL.n199 VTAIL.n178 9.69747
R257 VTAIL.n169 VTAIL.n148 9.69747
R258 VTAIL.n141 VTAIL.n120 9.69747
R259 VTAIL.n111 VTAIL.n90 9.69747
R260 VTAIL.n230 VTAIL.n229 9.45567
R261 VTAIL.n28 VTAIL.n27 9.45567
R262 VTAIL.n56 VTAIL.n55 9.45567
R263 VTAIL.n86 VTAIL.n85 9.45567
R264 VTAIL.n202 VTAIL.n201 9.45567
R265 VTAIL.n172 VTAIL.n171 9.45567
R266 VTAIL.n144 VTAIL.n143 9.45567
R267 VTAIL.n114 VTAIL.n113 9.45567
R268 VTAIL.n229 VTAIL.n228 9.3005
R269 VTAIL.n206 VTAIL.n205 9.3005
R270 VTAIL.n223 VTAIL.n222 9.3005
R271 VTAIL.n221 VTAIL.n220 9.3005
R272 VTAIL.n210 VTAIL.n209 9.3005
R273 VTAIL.n215 VTAIL.n214 9.3005
R274 VTAIL.n27 VTAIL.n26 9.3005
R275 VTAIL.n4 VTAIL.n3 9.3005
R276 VTAIL.n21 VTAIL.n20 9.3005
R277 VTAIL.n19 VTAIL.n18 9.3005
R278 VTAIL.n8 VTAIL.n7 9.3005
R279 VTAIL.n13 VTAIL.n12 9.3005
R280 VTAIL.n55 VTAIL.n54 9.3005
R281 VTAIL.n32 VTAIL.n31 9.3005
R282 VTAIL.n49 VTAIL.n48 9.3005
R283 VTAIL.n47 VTAIL.n46 9.3005
R284 VTAIL.n36 VTAIL.n35 9.3005
R285 VTAIL.n41 VTAIL.n40 9.3005
R286 VTAIL.n85 VTAIL.n84 9.3005
R287 VTAIL.n62 VTAIL.n61 9.3005
R288 VTAIL.n79 VTAIL.n78 9.3005
R289 VTAIL.n77 VTAIL.n76 9.3005
R290 VTAIL.n66 VTAIL.n65 9.3005
R291 VTAIL.n71 VTAIL.n70 9.3005
R292 VTAIL.n201 VTAIL.n200 9.3005
R293 VTAIL.n178 VTAIL.n177 9.3005
R294 VTAIL.n195 VTAIL.n194 9.3005
R295 VTAIL.n193 VTAIL.n192 9.3005
R296 VTAIL.n182 VTAIL.n181 9.3005
R297 VTAIL.n187 VTAIL.n186 9.3005
R298 VTAIL.n171 VTAIL.n170 9.3005
R299 VTAIL.n148 VTAIL.n147 9.3005
R300 VTAIL.n165 VTAIL.n164 9.3005
R301 VTAIL.n163 VTAIL.n162 9.3005
R302 VTAIL.n152 VTAIL.n151 9.3005
R303 VTAIL.n157 VTAIL.n156 9.3005
R304 VTAIL.n143 VTAIL.n142 9.3005
R305 VTAIL.n120 VTAIL.n119 9.3005
R306 VTAIL.n137 VTAIL.n136 9.3005
R307 VTAIL.n135 VTAIL.n134 9.3005
R308 VTAIL.n124 VTAIL.n123 9.3005
R309 VTAIL.n129 VTAIL.n128 9.3005
R310 VTAIL.n113 VTAIL.n112 9.3005
R311 VTAIL.n90 VTAIL.n89 9.3005
R312 VTAIL.n107 VTAIL.n106 9.3005
R313 VTAIL.n105 VTAIL.n104 9.3005
R314 VTAIL.n94 VTAIL.n93 9.3005
R315 VTAIL.n99 VTAIL.n98 9.3005
R316 VTAIL.n228 VTAIL.n204 8.92171
R317 VTAIL.n26 VTAIL.n2 8.92171
R318 VTAIL.n54 VTAIL.n30 8.92171
R319 VTAIL.n84 VTAIL.n60 8.92171
R320 VTAIL.n200 VTAIL.n176 8.92171
R321 VTAIL.n170 VTAIL.n146 8.92171
R322 VTAIL.n142 VTAIL.n118 8.92171
R323 VTAIL.n112 VTAIL.n88 8.92171
R324 VTAIL.n230 VTAIL.n204 5.04292
R325 VTAIL.n28 VTAIL.n2 5.04292
R326 VTAIL.n56 VTAIL.n30 5.04292
R327 VTAIL.n86 VTAIL.n60 5.04292
R328 VTAIL.n202 VTAIL.n176 5.04292
R329 VTAIL.n172 VTAIL.n146 5.04292
R330 VTAIL.n144 VTAIL.n118 5.04292
R331 VTAIL.n114 VTAIL.n88 5.04292
R332 VTAIL.n214 VTAIL.n213 4.38687
R333 VTAIL.n12 VTAIL.n11 4.38687
R334 VTAIL.n40 VTAIL.n39 4.38687
R335 VTAIL.n70 VTAIL.n69 4.38687
R336 VTAIL.n186 VTAIL.n185 4.38687
R337 VTAIL.n156 VTAIL.n155 4.38687
R338 VTAIL.n128 VTAIL.n127 4.38687
R339 VTAIL.n98 VTAIL.n97 4.38687
R340 VTAIL.n228 VTAIL.n227 4.26717
R341 VTAIL.n26 VTAIL.n25 4.26717
R342 VTAIL.n54 VTAIL.n53 4.26717
R343 VTAIL.n84 VTAIL.n83 4.26717
R344 VTAIL.n200 VTAIL.n199 4.26717
R345 VTAIL.n170 VTAIL.n169 4.26717
R346 VTAIL.n142 VTAIL.n141 4.26717
R347 VTAIL.n112 VTAIL.n111 4.26717
R348 VTAIL.n0 VTAIL.t10 3.65364
R349 VTAIL.n0 VTAIL.t6 3.65364
R350 VTAIL.n58 VTAIL.t2 3.65364
R351 VTAIL.n58 VTAIL.t15 3.65364
R352 VTAIL.n174 VTAIL.t1 3.65364
R353 VTAIL.n174 VTAIL.t3 3.65364
R354 VTAIL.n116 VTAIL.t9 3.65364
R355 VTAIL.n116 VTAIL.t11 3.65364
R356 VTAIL.n224 VTAIL.n206 3.49141
R357 VTAIL.n22 VTAIL.n4 3.49141
R358 VTAIL.n50 VTAIL.n32 3.49141
R359 VTAIL.n80 VTAIL.n62 3.49141
R360 VTAIL.n196 VTAIL.n178 3.49141
R361 VTAIL.n166 VTAIL.n148 3.49141
R362 VTAIL.n138 VTAIL.n120 3.49141
R363 VTAIL.n108 VTAIL.n90 3.49141
R364 VTAIL.n223 VTAIL.n208 2.71565
R365 VTAIL.n21 VTAIL.n6 2.71565
R366 VTAIL.n49 VTAIL.n34 2.71565
R367 VTAIL.n79 VTAIL.n64 2.71565
R368 VTAIL.n195 VTAIL.n180 2.71565
R369 VTAIL.n165 VTAIL.n150 2.71565
R370 VTAIL.n137 VTAIL.n122 2.71565
R371 VTAIL.n107 VTAIL.n92 2.71565
R372 VTAIL.n117 VTAIL.n115 2.32809
R373 VTAIL.n145 VTAIL.n117 2.32809
R374 VTAIL.n175 VTAIL.n173 2.32809
R375 VTAIL.n203 VTAIL.n175 2.32809
R376 VTAIL.n87 VTAIL.n59 2.32809
R377 VTAIL.n59 VTAIL.n57 2.32809
R378 VTAIL.n29 VTAIL.n1 2.32809
R379 VTAIL VTAIL.n231 2.2699
R380 VTAIL.n220 VTAIL.n219 1.93989
R381 VTAIL.n18 VTAIL.n17 1.93989
R382 VTAIL.n46 VTAIL.n45 1.93989
R383 VTAIL.n76 VTAIL.n75 1.93989
R384 VTAIL.n192 VTAIL.n191 1.93989
R385 VTAIL.n162 VTAIL.n161 1.93989
R386 VTAIL.n134 VTAIL.n133 1.93989
R387 VTAIL.n104 VTAIL.n103 1.93989
R388 VTAIL.n216 VTAIL.n210 1.16414
R389 VTAIL.n14 VTAIL.n8 1.16414
R390 VTAIL.n42 VTAIL.n36 1.16414
R391 VTAIL.n72 VTAIL.n66 1.16414
R392 VTAIL.n188 VTAIL.n182 1.16414
R393 VTAIL.n158 VTAIL.n152 1.16414
R394 VTAIL.n130 VTAIL.n124 1.16414
R395 VTAIL.n100 VTAIL.n94 1.16414
R396 VTAIL.n173 VTAIL.n145 0.470328
R397 VTAIL.n57 VTAIL.n29 0.470328
R398 VTAIL.n215 VTAIL.n212 0.388379
R399 VTAIL.n13 VTAIL.n10 0.388379
R400 VTAIL.n41 VTAIL.n38 0.388379
R401 VTAIL.n71 VTAIL.n68 0.388379
R402 VTAIL.n187 VTAIL.n184 0.388379
R403 VTAIL.n157 VTAIL.n154 0.388379
R404 VTAIL.n129 VTAIL.n126 0.388379
R405 VTAIL.n99 VTAIL.n96 0.388379
R406 VTAIL.n214 VTAIL.n209 0.155672
R407 VTAIL.n221 VTAIL.n209 0.155672
R408 VTAIL.n222 VTAIL.n221 0.155672
R409 VTAIL.n222 VTAIL.n205 0.155672
R410 VTAIL.n229 VTAIL.n205 0.155672
R411 VTAIL.n12 VTAIL.n7 0.155672
R412 VTAIL.n19 VTAIL.n7 0.155672
R413 VTAIL.n20 VTAIL.n19 0.155672
R414 VTAIL.n20 VTAIL.n3 0.155672
R415 VTAIL.n27 VTAIL.n3 0.155672
R416 VTAIL.n40 VTAIL.n35 0.155672
R417 VTAIL.n47 VTAIL.n35 0.155672
R418 VTAIL.n48 VTAIL.n47 0.155672
R419 VTAIL.n48 VTAIL.n31 0.155672
R420 VTAIL.n55 VTAIL.n31 0.155672
R421 VTAIL.n70 VTAIL.n65 0.155672
R422 VTAIL.n77 VTAIL.n65 0.155672
R423 VTAIL.n78 VTAIL.n77 0.155672
R424 VTAIL.n78 VTAIL.n61 0.155672
R425 VTAIL.n85 VTAIL.n61 0.155672
R426 VTAIL.n201 VTAIL.n177 0.155672
R427 VTAIL.n194 VTAIL.n177 0.155672
R428 VTAIL.n194 VTAIL.n193 0.155672
R429 VTAIL.n193 VTAIL.n181 0.155672
R430 VTAIL.n186 VTAIL.n181 0.155672
R431 VTAIL.n171 VTAIL.n147 0.155672
R432 VTAIL.n164 VTAIL.n147 0.155672
R433 VTAIL.n164 VTAIL.n163 0.155672
R434 VTAIL.n163 VTAIL.n151 0.155672
R435 VTAIL.n156 VTAIL.n151 0.155672
R436 VTAIL.n143 VTAIL.n119 0.155672
R437 VTAIL.n136 VTAIL.n119 0.155672
R438 VTAIL.n136 VTAIL.n135 0.155672
R439 VTAIL.n135 VTAIL.n123 0.155672
R440 VTAIL.n128 VTAIL.n123 0.155672
R441 VTAIL.n113 VTAIL.n89 0.155672
R442 VTAIL.n106 VTAIL.n89 0.155672
R443 VTAIL.n106 VTAIL.n105 0.155672
R444 VTAIL.n105 VTAIL.n93 0.155672
R445 VTAIL.n98 VTAIL.n93 0.155672
R446 VTAIL VTAIL.n1 0.0586897
R447 VDD2.n2 VDD2.n1 72.4787
R448 VDD2.n2 VDD2.n0 72.4787
R449 VDD2 VDD2.n5 72.4759
R450 VDD2.n4 VDD2.n3 71.3704
R451 VDD2.n4 VDD2.n2 38.8618
R452 VDD2.n5 VDD2.t6 3.65364
R453 VDD2.n5 VDD2.t1 3.65364
R454 VDD2.n3 VDD2.t4 3.65364
R455 VDD2.n3 VDD2.t0 3.65364
R456 VDD2.n1 VDD2.t2 3.65364
R457 VDD2.n1 VDD2.t5 3.65364
R458 VDD2.n0 VDD2.t3 3.65364
R459 VDD2.n0 VDD2.t7 3.65364
R460 VDD2 VDD2.n4 1.22248
R461 B.n666 B.n665 585
R462 B.n225 B.n116 585
R463 B.n224 B.n223 585
R464 B.n222 B.n221 585
R465 B.n220 B.n219 585
R466 B.n218 B.n217 585
R467 B.n216 B.n215 585
R468 B.n214 B.n213 585
R469 B.n212 B.n211 585
R470 B.n210 B.n209 585
R471 B.n208 B.n207 585
R472 B.n206 B.n205 585
R473 B.n204 B.n203 585
R474 B.n202 B.n201 585
R475 B.n200 B.n199 585
R476 B.n198 B.n197 585
R477 B.n196 B.n195 585
R478 B.n194 B.n193 585
R479 B.n192 B.n191 585
R480 B.n190 B.n189 585
R481 B.n188 B.n187 585
R482 B.n186 B.n185 585
R483 B.n184 B.n183 585
R484 B.n182 B.n181 585
R485 B.n180 B.n179 585
R486 B.n178 B.n177 585
R487 B.n176 B.n175 585
R488 B.n174 B.n173 585
R489 B.n172 B.n171 585
R490 B.n170 B.n169 585
R491 B.n168 B.n167 585
R492 B.n166 B.n165 585
R493 B.n164 B.n163 585
R494 B.n162 B.n161 585
R495 B.n160 B.n159 585
R496 B.n158 B.n157 585
R497 B.n156 B.n155 585
R498 B.n154 B.n153 585
R499 B.n152 B.n151 585
R500 B.n150 B.n149 585
R501 B.n148 B.n147 585
R502 B.n146 B.n145 585
R503 B.n144 B.n143 585
R504 B.n142 B.n141 585
R505 B.n140 B.n139 585
R506 B.n138 B.n137 585
R507 B.n136 B.n135 585
R508 B.n134 B.n133 585
R509 B.n132 B.n131 585
R510 B.n130 B.n129 585
R511 B.n128 B.n127 585
R512 B.n126 B.n125 585
R513 B.n124 B.n123 585
R514 B.n88 B.n87 585
R515 B.n664 B.n89 585
R516 B.n669 B.n89 585
R517 B.n663 B.n662 585
R518 B.n662 B.n85 585
R519 B.n661 B.n84 585
R520 B.n675 B.n84 585
R521 B.n660 B.n83 585
R522 B.n676 B.n83 585
R523 B.n659 B.n82 585
R524 B.n677 B.n82 585
R525 B.n658 B.n657 585
R526 B.n657 B.n78 585
R527 B.n656 B.n77 585
R528 B.n683 B.n77 585
R529 B.n655 B.n76 585
R530 B.n684 B.n76 585
R531 B.n654 B.n75 585
R532 B.n685 B.n75 585
R533 B.n653 B.n652 585
R534 B.n652 B.n71 585
R535 B.n651 B.n70 585
R536 B.n691 B.n70 585
R537 B.n650 B.n69 585
R538 B.n692 B.n69 585
R539 B.n649 B.n68 585
R540 B.n693 B.n68 585
R541 B.n648 B.n647 585
R542 B.n647 B.n64 585
R543 B.n646 B.n63 585
R544 B.n699 B.n63 585
R545 B.n645 B.n62 585
R546 B.n700 B.n62 585
R547 B.n644 B.n61 585
R548 B.n701 B.n61 585
R549 B.n643 B.n642 585
R550 B.n642 B.n57 585
R551 B.n641 B.n56 585
R552 B.n707 B.n56 585
R553 B.n640 B.n55 585
R554 B.n708 B.n55 585
R555 B.n639 B.n54 585
R556 B.n709 B.n54 585
R557 B.n638 B.n637 585
R558 B.n637 B.n50 585
R559 B.n636 B.n49 585
R560 B.n715 B.n49 585
R561 B.n635 B.n48 585
R562 B.n716 B.n48 585
R563 B.n634 B.n47 585
R564 B.n717 B.n47 585
R565 B.n633 B.n632 585
R566 B.n632 B.n43 585
R567 B.n631 B.n42 585
R568 B.n723 B.n42 585
R569 B.n630 B.n41 585
R570 B.n724 B.n41 585
R571 B.n629 B.n40 585
R572 B.n725 B.n40 585
R573 B.n628 B.n627 585
R574 B.n627 B.n36 585
R575 B.n626 B.n35 585
R576 B.n731 B.n35 585
R577 B.n625 B.n34 585
R578 B.n732 B.n34 585
R579 B.n624 B.n33 585
R580 B.n733 B.n33 585
R581 B.n623 B.n622 585
R582 B.n622 B.n29 585
R583 B.n621 B.n28 585
R584 B.n739 B.n28 585
R585 B.n620 B.n27 585
R586 B.n740 B.n27 585
R587 B.n619 B.n26 585
R588 B.n741 B.n26 585
R589 B.n618 B.n617 585
R590 B.n617 B.n22 585
R591 B.n616 B.n21 585
R592 B.n747 B.n21 585
R593 B.n615 B.n20 585
R594 B.n748 B.n20 585
R595 B.n614 B.n19 585
R596 B.n749 B.n19 585
R597 B.n613 B.n612 585
R598 B.n612 B.n15 585
R599 B.n611 B.n14 585
R600 B.n755 B.n14 585
R601 B.n610 B.n13 585
R602 B.n756 B.n13 585
R603 B.n609 B.n12 585
R604 B.n757 B.n12 585
R605 B.n608 B.n607 585
R606 B.n607 B.n8 585
R607 B.n606 B.n7 585
R608 B.n763 B.n7 585
R609 B.n605 B.n6 585
R610 B.n764 B.n6 585
R611 B.n604 B.n5 585
R612 B.n765 B.n5 585
R613 B.n603 B.n602 585
R614 B.n602 B.n4 585
R615 B.n601 B.n226 585
R616 B.n601 B.n600 585
R617 B.n591 B.n227 585
R618 B.n228 B.n227 585
R619 B.n593 B.n592 585
R620 B.n594 B.n593 585
R621 B.n590 B.n233 585
R622 B.n233 B.n232 585
R623 B.n589 B.n588 585
R624 B.n588 B.n587 585
R625 B.n235 B.n234 585
R626 B.n236 B.n235 585
R627 B.n580 B.n579 585
R628 B.n581 B.n580 585
R629 B.n578 B.n241 585
R630 B.n241 B.n240 585
R631 B.n577 B.n576 585
R632 B.n576 B.n575 585
R633 B.n243 B.n242 585
R634 B.n244 B.n243 585
R635 B.n568 B.n567 585
R636 B.n569 B.n568 585
R637 B.n566 B.n249 585
R638 B.n249 B.n248 585
R639 B.n565 B.n564 585
R640 B.n564 B.n563 585
R641 B.n251 B.n250 585
R642 B.n252 B.n251 585
R643 B.n556 B.n555 585
R644 B.n557 B.n556 585
R645 B.n554 B.n257 585
R646 B.n257 B.n256 585
R647 B.n553 B.n552 585
R648 B.n552 B.n551 585
R649 B.n259 B.n258 585
R650 B.n260 B.n259 585
R651 B.n544 B.n543 585
R652 B.n545 B.n544 585
R653 B.n542 B.n265 585
R654 B.n265 B.n264 585
R655 B.n541 B.n540 585
R656 B.n540 B.n539 585
R657 B.n267 B.n266 585
R658 B.n268 B.n267 585
R659 B.n532 B.n531 585
R660 B.n533 B.n532 585
R661 B.n530 B.n273 585
R662 B.n273 B.n272 585
R663 B.n529 B.n528 585
R664 B.n528 B.n527 585
R665 B.n275 B.n274 585
R666 B.n276 B.n275 585
R667 B.n520 B.n519 585
R668 B.n521 B.n520 585
R669 B.n518 B.n281 585
R670 B.n281 B.n280 585
R671 B.n517 B.n516 585
R672 B.n516 B.n515 585
R673 B.n283 B.n282 585
R674 B.n284 B.n283 585
R675 B.n508 B.n507 585
R676 B.n509 B.n508 585
R677 B.n506 B.n289 585
R678 B.n289 B.n288 585
R679 B.n505 B.n504 585
R680 B.n504 B.n503 585
R681 B.n291 B.n290 585
R682 B.n292 B.n291 585
R683 B.n496 B.n495 585
R684 B.n497 B.n496 585
R685 B.n494 B.n297 585
R686 B.n297 B.n296 585
R687 B.n493 B.n492 585
R688 B.n492 B.n491 585
R689 B.n299 B.n298 585
R690 B.n300 B.n299 585
R691 B.n484 B.n483 585
R692 B.n485 B.n484 585
R693 B.n482 B.n304 585
R694 B.n308 B.n304 585
R695 B.n481 B.n480 585
R696 B.n480 B.n479 585
R697 B.n306 B.n305 585
R698 B.n307 B.n306 585
R699 B.n472 B.n471 585
R700 B.n473 B.n472 585
R701 B.n470 B.n313 585
R702 B.n313 B.n312 585
R703 B.n469 B.n468 585
R704 B.n468 B.n467 585
R705 B.n315 B.n314 585
R706 B.n316 B.n315 585
R707 B.n460 B.n459 585
R708 B.n461 B.n460 585
R709 B.n319 B.n318 585
R710 B.n352 B.n350 585
R711 B.n353 B.n349 585
R712 B.n353 B.n320 585
R713 B.n356 B.n355 585
R714 B.n357 B.n348 585
R715 B.n359 B.n358 585
R716 B.n361 B.n347 585
R717 B.n364 B.n363 585
R718 B.n365 B.n346 585
R719 B.n367 B.n366 585
R720 B.n369 B.n345 585
R721 B.n372 B.n371 585
R722 B.n373 B.n344 585
R723 B.n375 B.n374 585
R724 B.n377 B.n343 585
R725 B.n380 B.n379 585
R726 B.n381 B.n342 585
R727 B.n383 B.n382 585
R728 B.n385 B.n341 585
R729 B.n388 B.n387 585
R730 B.n389 B.n340 585
R731 B.n394 B.n393 585
R732 B.n396 B.n339 585
R733 B.n399 B.n398 585
R734 B.n400 B.n338 585
R735 B.n402 B.n401 585
R736 B.n404 B.n337 585
R737 B.n407 B.n406 585
R738 B.n408 B.n336 585
R739 B.n410 B.n409 585
R740 B.n412 B.n335 585
R741 B.n415 B.n414 585
R742 B.n417 B.n332 585
R743 B.n419 B.n418 585
R744 B.n421 B.n331 585
R745 B.n424 B.n423 585
R746 B.n425 B.n330 585
R747 B.n427 B.n426 585
R748 B.n429 B.n329 585
R749 B.n432 B.n431 585
R750 B.n433 B.n328 585
R751 B.n435 B.n434 585
R752 B.n437 B.n327 585
R753 B.n440 B.n439 585
R754 B.n441 B.n326 585
R755 B.n443 B.n442 585
R756 B.n445 B.n325 585
R757 B.n448 B.n447 585
R758 B.n449 B.n324 585
R759 B.n451 B.n450 585
R760 B.n453 B.n323 585
R761 B.n454 B.n322 585
R762 B.n457 B.n456 585
R763 B.n458 B.n321 585
R764 B.n321 B.n320 585
R765 B.n463 B.n462 585
R766 B.n462 B.n461 585
R767 B.n464 B.n317 585
R768 B.n317 B.n316 585
R769 B.n466 B.n465 585
R770 B.n467 B.n466 585
R771 B.n311 B.n310 585
R772 B.n312 B.n311 585
R773 B.n475 B.n474 585
R774 B.n474 B.n473 585
R775 B.n476 B.n309 585
R776 B.n309 B.n307 585
R777 B.n478 B.n477 585
R778 B.n479 B.n478 585
R779 B.n303 B.n302 585
R780 B.n308 B.n303 585
R781 B.n487 B.n486 585
R782 B.n486 B.n485 585
R783 B.n488 B.n301 585
R784 B.n301 B.n300 585
R785 B.n490 B.n489 585
R786 B.n491 B.n490 585
R787 B.n295 B.n294 585
R788 B.n296 B.n295 585
R789 B.n499 B.n498 585
R790 B.n498 B.n497 585
R791 B.n500 B.n293 585
R792 B.n293 B.n292 585
R793 B.n502 B.n501 585
R794 B.n503 B.n502 585
R795 B.n287 B.n286 585
R796 B.n288 B.n287 585
R797 B.n511 B.n510 585
R798 B.n510 B.n509 585
R799 B.n512 B.n285 585
R800 B.n285 B.n284 585
R801 B.n514 B.n513 585
R802 B.n515 B.n514 585
R803 B.n279 B.n278 585
R804 B.n280 B.n279 585
R805 B.n523 B.n522 585
R806 B.n522 B.n521 585
R807 B.n524 B.n277 585
R808 B.n277 B.n276 585
R809 B.n526 B.n525 585
R810 B.n527 B.n526 585
R811 B.n271 B.n270 585
R812 B.n272 B.n271 585
R813 B.n535 B.n534 585
R814 B.n534 B.n533 585
R815 B.n536 B.n269 585
R816 B.n269 B.n268 585
R817 B.n538 B.n537 585
R818 B.n539 B.n538 585
R819 B.n263 B.n262 585
R820 B.n264 B.n263 585
R821 B.n547 B.n546 585
R822 B.n546 B.n545 585
R823 B.n548 B.n261 585
R824 B.n261 B.n260 585
R825 B.n550 B.n549 585
R826 B.n551 B.n550 585
R827 B.n255 B.n254 585
R828 B.n256 B.n255 585
R829 B.n559 B.n558 585
R830 B.n558 B.n557 585
R831 B.n560 B.n253 585
R832 B.n253 B.n252 585
R833 B.n562 B.n561 585
R834 B.n563 B.n562 585
R835 B.n247 B.n246 585
R836 B.n248 B.n247 585
R837 B.n571 B.n570 585
R838 B.n570 B.n569 585
R839 B.n572 B.n245 585
R840 B.n245 B.n244 585
R841 B.n574 B.n573 585
R842 B.n575 B.n574 585
R843 B.n239 B.n238 585
R844 B.n240 B.n239 585
R845 B.n583 B.n582 585
R846 B.n582 B.n581 585
R847 B.n584 B.n237 585
R848 B.n237 B.n236 585
R849 B.n586 B.n585 585
R850 B.n587 B.n586 585
R851 B.n231 B.n230 585
R852 B.n232 B.n231 585
R853 B.n596 B.n595 585
R854 B.n595 B.n594 585
R855 B.n597 B.n229 585
R856 B.n229 B.n228 585
R857 B.n599 B.n598 585
R858 B.n600 B.n599 585
R859 B.n2 B.n0 585
R860 B.n4 B.n2 585
R861 B.n3 B.n1 585
R862 B.n764 B.n3 585
R863 B.n762 B.n761 585
R864 B.n763 B.n762 585
R865 B.n760 B.n9 585
R866 B.n9 B.n8 585
R867 B.n759 B.n758 585
R868 B.n758 B.n757 585
R869 B.n11 B.n10 585
R870 B.n756 B.n11 585
R871 B.n754 B.n753 585
R872 B.n755 B.n754 585
R873 B.n752 B.n16 585
R874 B.n16 B.n15 585
R875 B.n751 B.n750 585
R876 B.n750 B.n749 585
R877 B.n18 B.n17 585
R878 B.n748 B.n18 585
R879 B.n746 B.n745 585
R880 B.n747 B.n746 585
R881 B.n744 B.n23 585
R882 B.n23 B.n22 585
R883 B.n743 B.n742 585
R884 B.n742 B.n741 585
R885 B.n25 B.n24 585
R886 B.n740 B.n25 585
R887 B.n738 B.n737 585
R888 B.n739 B.n738 585
R889 B.n736 B.n30 585
R890 B.n30 B.n29 585
R891 B.n735 B.n734 585
R892 B.n734 B.n733 585
R893 B.n32 B.n31 585
R894 B.n732 B.n32 585
R895 B.n730 B.n729 585
R896 B.n731 B.n730 585
R897 B.n728 B.n37 585
R898 B.n37 B.n36 585
R899 B.n727 B.n726 585
R900 B.n726 B.n725 585
R901 B.n39 B.n38 585
R902 B.n724 B.n39 585
R903 B.n722 B.n721 585
R904 B.n723 B.n722 585
R905 B.n720 B.n44 585
R906 B.n44 B.n43 585
R907 B.n719 B.n718 585
R908 B.n718 B.n717 585
R909 B.n46 B.n45 585
R910 B.n716 B.n46 585
R911 B.n714 B.n713 585
R912 B.n715 B.n714 585
R913 B.n712 B.n51 585
R914 B.n51 B.n50 585
R915 B.n711 B.n710 585
R916 B.n710 B.n709 585
R917 B.n53 B.n52 585
R918 B.n708 B.n53 585
R919 B.n706 B.n705 585
R920 B.n707 B.n706 585
R921 B.n704 B.n58 585
R922 B.n58 B.n57 585
R923 B.n703 B.n702 585
R924 B.n702 B.n701 585
R925 B.n60 B.n59 585
R926 B.n700 B.n60 585
R927 B.n698 B.n697 585
R928 B.n699 B.n698 585
R929 B.n696 B.n65 585
R930 B.n65 B.n64 585
R931 B.n695 B.n694 585
R932 B.n694 B.n693 585
R933 B.n67 B.n66 585
R934 B.n692 B.n67 585
R935 B.n690 B.n689 585
R936 B.n691 B.n690 585
R937 B.n688 B.n72 585
R938 B.n72 B.n71 585
R939 B.n687 B.n686 585
R940 B.n686 B.n685 585
R941 B.n74 B.n73 585
R942 B.n684 B.n74 585
R943 B.n682 B.n681 585
R944 B.n683 B.n682 585
R945 B.n680 B.n79 585
R946 B.n79 B.n78 585
R947 B.n679 B.n678 585
R948 B.n678 B.n677 585
R949 B.n81 B.n80 585
R950 B.n676 B.n81 585
R951 B.n674 B.n673 585
R952 B.n675 B.n674 585
R953 B.n672 B.n86 585
R954 B.n86 B.n85 585
R955 B.n671 B.n670 585
R956 B.n670 B.n669 585
R957 B.n767 B.n766 585
R958 B.n766 B.n765 585
R959 B.n462 B.n319 478.086
R960 B.n670 B.n88 478.086
R961 B.n460 B.n321 478.086
R962 B.n666 B.n89 478.086
R963 B.n333 B.t15 262.786
R964 B.n390 B.t19 262.786
R965 B.n120 B.t12 262.786
R966 B.n117 B.t8 262.786
R967 B.n668 B.n667 256.663
R968 B.n668 B.n115 256.663
R969 B.n668 B.n114 256.663
R970 B.n668 B.n113 256.663
R971 B.n668 B.n112 256.663
R972 B.n668 B.n111 256.663
R973 B.n668 B.n110 256.663
R974 B.n668 B.n109 256.663
R975 B.n668 B.n108 256.663
R976 B.n668 B.n107 256.663
R977 B.n668 B.n106 256.663
R978 B.n668 B.n105 256.663
R979 B.n668 B.n104 256.663
R980 B.n668 B.n103 256.663
R981 B.n668 B.n102 256.663
R982 B.n668 B.n101 256.663
R983 B.n668 B.n100 256.663
R984 B.n668 B.n99 256.663
R985 B.n668 B.n98 256.663
R986 B.n668 B.n97 256.663
R987 B.n668 B.n96 256.663
R988 B.n668 B.n95 256.663
R989 B.n668 B.n94 256.663
R990 B.n668 B.n93 256.663
R991 B.n668 B.n92 256.663
R992 B.n668 B.n91 256.663
R993 B.n668 B.n90 256.663
R994 B.n351 B.n320 256.663
R995 B.n354 B.n320 256.663
R996 B.n360 B.n320 256.663
R997 B.n362 B.n320 256.663
R998 B.n368 B.n320 256.663
R999 B.n370 B.n320 256.663
R1000 B.n376 B.n320 256.663
R1001 B.n378 B.n320 256.663
R1002 B.n384 B.n320 256.663
R1003 B.n386 B.n320 256.663
R1004 B.n395 B.n320 256.663
R1005 B.n397 B.n320 256.663
R1006 B.n403 B.n320 256.663
R1007 B.n405 B.n320 256.663
R1008 B.n411 B.n320 256.663
R1009 B.n413 B.n320 256.663
R1010 B.n420 B.n320 256.663
R1011 B.n422 B.n320 256.663
R1012 B.n428 B.n320 256.663
R1013 B.n430 B.n320 256.663
R1014 B.n436 B.n320 256.663
R1015 B.n438 B.n320 256.663
R1016 B.n444 B.n320 256.663
R1017 B.n446 B.n320 256.663
R1018 B.n452 B.n320 256.663
R1019 B.n455 B.n320 256.663
R1020 B.n333 B.t18 221.653
R1021 B.n117 B.t10 221.653
R1022 B.n390 B.t21 221.653
R1023 B.n120 B.t13 221.653
R1024 B.n334 B.t17 169.29
R1025 B.n118 B.t11 169.29
R1026 B.n391 B.t20 169.288
R1027 B.n121 B.t14 169.288
R1028 B.n462 B.n317 163.367
R1029 B.n466 B.n317 163.367
R1030 B.n466 B.n311 163.367
R1031 B.n474 B.n311 163.367
R1032 B.n474 B.n309 163.367
R1033 B.n478 B.n309 163.367
R1034 B.n478 B.n303 163.367
R1035 B.n486 B.n303 163.367
R1036 B.n486 B.n301 163.367
R1037 B.n490 B.n301 163.367
R1038 B.n490 B.n295 163.367
R1039 B.n498 B.n295 163.367
R1040 B.n498 B.n293 163.367
R1041 B.n502 B.n293 163.367
R1042 B.n502 B.n287 163.367
R1043 B.n510 B.n287 163.367
R1044 B.n510 B.n285 163.367
R1045 B.n514 B.n285 163.367
R1046 B.n514 B.n279 163.367
R1047 B.n522 B.n279 163.367
R1048 B.n522 B.n277 163.367
R1049 B.n526 B.n277 163.367
R1050 B.n526 B.n271 163.367
R1051 B.n534 B.n271 163.367
R1052 B.n534 B.n269 163.367
R1053 B.n538 B.n269 163.367
R1054 B.n538 B.n263 163.367
R1055 B.n546 B.n263 163.367
R1056 B.n546 B.n261 163.367
R1057 B.n550 B.n261 163.367
R1058 B.n550 B.n255 163.367
R1059 B.n558 B.n255 163.367
R1060 B.n558 B.n253 163.367
R1061 B.n562 B.n253 163.367
R1062 B.n562 B.n247 163.367
R1063 B.n570 B.n247 163.367
R1064 B.n570 B.n245 163.367
R1065 B.n574 B.n245 163.367
R1066 B.n574 B.n239 163.367
R1067 B.n582 B.n239 163.367
R1068 B.n582 B.n237 163.367
R1069 B.n586 B.n237 163.367
R1070 B.n586 B.n231 163.367
R1071 B.n595 B.n231 163.367
R1072 B.n595 B.n229 163.367
R1073 B.n599 B.n229 163.367
R1074 B.n599 B.n2 163.367
R1075 B.n766 B.n2 163.367
R1076 B.n766 B.n3 163.367
R1077 B.n762 B.n3 163.367
R1078 B.n762 B.n9 163.367
R1079 B.n758 B.n9 163.367
R1080 B.n758 B.n11 163.367
R1081 B.n754 B.n11 163.367
R1082 B.n754 B.n16 163.367
R1083 B.n750 B.n16 163.367
R1084 B.n750 B.n18 163.367
R1085 B.n746 B.n18 163.367
R1086 B.n746 B.n23 163.367
R1087 B.n742 B.n23 163.367
R1088 B.n742 B.n25 163.367
R1089 B.n738 B.n25 163.367
R1090 B.n738 B.n30 163.367
R1091 B.n734 B.n30 163.367
R1092 B.n734 B.n32 163.367
R1093 B.n730 B.n32 163.367
R1094 B.n730 B.n37 163.367
R1095 B.n726 B.n37 163.367
R1096 B.n726 B.n39 163.367
R1097 B.n722 B.n39 163.367
R1098 B.n722 B.n44 163.367
R1099 B.n718 B.n44 163.367
R1100 B.n718 B.n46 163.367
R1101 B.n714 B.n46 163.367
R1102 B.n714 B.n51 163.367
R1103 B.n710 B.n51 163.367
R1104 B.n710 B.n53 163.367
R1105 B.n706 B.n53 163.367
R1106 B.n706 B.n58 163.367
R1107 B.n702 B.n58 163.367
R1108 B.n702 B.n60 163.367
R1109 B.n698 B.n60 163.367
R1110 B.n698 B.n65 163.367
R1111 B.n694 B.n65 163.367
R1112 B.n694 B.n67 163.367
R1113 B.n690 B.n67 163.367
R1114 B.n690 B.n72 163.367
R1115 B.n686 B.n72 163.367
R1116 B.n686 B.n74 163.367
R1117 B.n682 B.n74 163.367
R1118 B.n682 B.n79 163.367
R1119 B.n678 B.n79 163.367
R1120 B.n678 B.n81 163.367
R1121 B.n674 B.n81 163.367
R1122 B.n674 B.n86 163.367
R1123 B.n670 B.n86 163.367
R1124 B.n353 B.n352 163.367
R1125 B.n355 B.n353 163.367
R1126 B.n359 B.n348 163.367
R1127 B.n363 B.n361 163.367
R1128 B.n367 B.n346 163.367
R1129 B.n371 B.n369 163.367
R1130 B.n375 B.n344 163.367
R1131 B.n379 B.n377 163.367
R1132 B.n383 B.n342 163.367
R1133 B.n387 B.n385 163.367
R1134 B.n394 B.n340 163.367
R1135 B.n398 B.n396 163.367
R1136 B.n402 B.n338 163.367
R1137 B.n406 B.n404 163.367
R1138 B.n410 B.n336 163.367
R1139 B.n414 B.n412 163.367
R1140 B.n419 B.n332 163.367
R1141 B.n423 B.n421 163.367
R1142 B.n427 B.n330 163.367
R1143 B.n431 B.n429 163.367
R1144 B.n435 B.n328 163.367
R1145 B.n439 B.n437 163.367
R1146 B.n443 B.n326 163.367
R1147 B.n447 B.n445 163.367
R1148 B.n451 B.n324 163.367
R1149 B.n454 B.n453 163.367
R1150 B.n456 B.n321 163.367
R1151 B.n460 B.n315 163.367
R1152 B.n468 B.n315 163.367
R1153 B.n468 B.n313 163.367
R1154 B.n472 B.n313 163.367
R1155 B.n472 B.n306 163.367
R1156 B.n480 B.n306 163.367
R1157 B.n480 B.n304 163.367
R1158 B.n484 B.n304 163.367
R1159 B.n484 B.n299 163.367
R1160 B.n492 B.n299 163.367
R1161 B.n492 B.n297 163.367
R1162 B.n496 B.n297 163.367
R1163 B.n496 B.n291 163.367
R1164 B.n504 B.n291 163.367
R1165 B.n504 B.n289 163.367
R1166 B.n508 B.n289 163.367
R1167 B.n508 B.n283 163.367
R1168 B.n516 B.n283 163.367
R1169 B.n516 B.n281 163.367
R1170 B.n520 B.n281 163.367
R1171 B.n520 B.n275 163.367
R1172 B.n528 B.n275 163.367
R1173 B.n528 B.n273 163.367
R1174 B.n532 B.n273 163.367
R1175 B.n532 B.n267 163.367
R1176 B.n540 B.n267 163.367
R1177 B.n540 B.n265 163.367
R1178 B.n544 B.n265 163.367
R1179 B.n544 B.n259 163.367
R1180 B.n552 B.n259 163.367
R1181 B.n552 B.n257 163.367
R1182 B.n556 B.n257 163.367
R1183 B.n556 B.n251 163.367
R1184 B.n564 B.n251 163.367
R1185 B.n564 B.n249 163.367
R1186 B.n568 B.n249 163.367
R1187 B.n568 B.n243 163.367
R1188 B.n576 B.n243 163.367
R1189 B.n576 B.n241 163.367
R1190 B.n580 B.n241 163.367
R1191 B.n580 B.n235 163.367
R1192 B.n588 B.n235 163.367
R1193 B.n588 B.n233 163.367
R1194 B.n593 B.n233 163.367
R1195 B.n593 B.n227 163.367
R1196 B.n601 B.n227 163.367
R1197 B.n602 B.n601 163.367
R1198 B.n602 B.n5 163.367
R1199 B.n6 B.n5 163.367
R1200 B.n7 B.n6 163.367
R1201 B.n607 B.n7 163.367
R1202 B.n607 B.n12 163.367
R1203 B.n13 B.n12 163.367
R1204 B.n14 B.n13 163.367
R1205 B.n612 B.n14 163.367
R1206 B.n612 B.n19 163.367
R1207 B.n20 B.n19 163.367
R1208 B.n21 B.n20 163.367
R1209 B.n617 B.n21 163.367
R1210 B.n617 B.n26 163.367
R1211 B.n27 B.n26 163.367
R1212 B.n28 B.n27 163.367
R1213 B.n622 B.n28 163.367
R1214 B.n622 B.n33 163.367
R1215 B.n34 B.n33 163.367
R1216 B.n35 B.n34 163.367
R1217 B.n627 B.n35 163.367
R1218 B.n627 B.n40 163.367
R1219 B.n41 B.n40 163.367
R1220 B.n42 B.n41 163.367
R1221 B.n632 B.n42 163.367
R1222 B.n632 B.n47 163.367
R1223 B.n48 B.n47 163.367
R1224 B.n49 B.n48 163.367
R1225 B.n637 B.n49 163.367
R1226 B.n637 B.n54 163.367
R1227 B.n55 B.n54 163.367
R1228 B.n56 B.n55 163.367
R1229 B.n642 B.n56 163.367
R1230 B.n642 B.n61 163.367
R1231 B.n62 B.n61 163.367
R1232 B.n63 B.n62 163.367
R1233 B.n647 B.n63 163.367
R1234 B.n647 B.n68 163.367
R1235 B.n69 B.n68 163.367
R1236 B.n70 B.n69 163.367
R1237 B.n652 B.n70 163.367
R1238 B.n652 B.n75 163.367
R1239 B.n76 B.n75 163.367
R1240 B.n77 B.n76 163.367
R1241 B.n657 B.n77 163.367
R1242 B.n657 B.n82 163.367
R1243 B.n83 B.n82 163.367
R1244 B.n84 B.n83 163.367
R1245 B.n662 B.n84 163.367
R1246 B.n662 B.n89 163.367
R1247 B.n125 B.n124 163.367
R1248 B.n129 B.n128 163.367
R1249 B.n133 B.n132 163.367
R1250 B.n137 B.n136 163.367
R1251 B.n141 B.n140 163.367
R1252 B.n145 B.n144 163.367
R1253 B.n149 B.n148 163.367
R1254 B.n153 B.n152 163.367
R1255 B.n157 B.n156 163.367
R1256 B.n161 B.n160 163.367
R1257 B.n165 B.n164 163.367
R1258 B.n169 B.n168 163.367
R1259 B.n173 B.n172 163.367
R1260 B.n177 B.n176 163.367
R1261 B.n181 B.n180 163.367
R1262 B.n185 B.n184 163.367
R1263 B.n189 B.n188 163.367
R1264 B.n193 B.n192 163.367
R1265 B.n197 B.n196 163.367
R1266 B.n201 B.n200 163.367
R1267 B.n205 B.n204 163.367
R1268 B.n209 B.n208 163.367
R1269 B.n213 B.n212 163.367
R1270 B.n217 B.n216 163.367
R1271 B.n221 B.n220 163.367
R1272 B.n223 B.n116 163.367
R1273 B.n461 B.n320 114.165
R1274 B.n669 B.n668 114.165
R1275 B.n351 B.n319 71.676
R1276 B.n355 B.n354 71.676
R1277 B.n360 B.n359 71.676
R1278 B.n363 B.n362 71.676
R1279 B.n368 B.n367 71.676
R1280 B.n371 B.n370 71.676
R1281 B.n376 B.n375 71.676
R1282 B.n379 B.n378 71.676
R1283 B.n384 B.n383 71.676
R1284 B.n387 B.n386 71.676
R1285 B.n395 B.n394 71.676
R1286 B.n398 B.n397 71.676
R1287 B.n403 B.n402 71.676
R1288 B.n406 B.n405 71.676
R1289 B.n411 B.n410 71.676
R1290 B.n414 B.n413 71.676
R1291 B.n420 B.n419 71.676
R1292 B.n423 B.n422 71.676
R1293 B.n428 B.n427 71.676
R1294 B.n431 B.n430 71.676
R1295 B.n436 B.n435 71.676
R1296 B.n439 B.n438 71.676
R1297 B.n444 B.n443 71.676
R1298 B.n447 B.n446 71.676
R1299 B.n452 B.n451 71.676
R1300 B.n455 B.n454 71.676
R1301 B.n90 B.n88 71.676
R1302 B.n125 B.n91 71.676
R1303 B.n129 B.n92 71.676
R1304 B.n133 B.n93 71.676
R1305 B.n137 B.n94 71.676
R1306 B.n141 B.n95 71.676
R1307 B.n145 B.n96 71.676
R1308 B.n149 B.n97 71.676
R1309 B.n153 B.n98 71.676
R1310 B.n157 B.n99 71.676
R1311 B.n161 B.n100 71.676
R1312 B.n165 B.n101 71.676
R1313 B.n169 B.n102 71.676
R1314 B.n173 B.n103 71.676
R1315 B.n177 B.n104 71.676
R1316 B.n181 B.n105 71.676
R1317 B.n185 B.n106 71.676
R1318 B.n189 B.n107 71.676
R1319 B.n193 B.n108 71.676
R1320 B.n197 B.n109 71.676
R1321 B.n201 B.n110 71.676
R1322 B.n205 B.n111 71.676
R1323 B.n209 B.n112 71.676
R1324 B.n213 B.n113 71.676
R1325 B.n217 B.n114 71.676
R1326 B.n221 B.n115 71.676
R1327 B.n667 B.n116 71.676
R1328 B.n667 B.n666 71.676
R1329 B.n223 B.n115 71.676
R1330 B.n220 B.n114 71.676
R1331 B.n216 B.n113 71.676
R1332 B.n212 B.n112 71.676
R1333 B.n208 B.n111 71.676
R1334 B.n204 B.n110 71.676
R1335 B.n200 B.n109 71.676
R1336 B.n196 B.n108 71.676
R1337 B.n192 B.n107 71.676
R1338 B.n188 B.n106 71.676
R1339 B.n184 B.n105 71.676
R1340 B.n180 B.n104 71.676
R1341 B.n176 B.n103 71.676
R1342 B.n172 B.n102 71.676
R1343 B.n168 B.n101 71.676
R1344 B.n164 B.n100 71.676
R1345 B.n160 B.n99 71.676
R1346 B.n156 B.n98 71.676
R1347 B.n152 B.n97 71.676
R1348 B.n148 B.n96 71.676
R1349 B.n144 B.n95 71.676
R1350 B.n140 B.n94 71.676
R1351 B.n136 B.n93 71.676
R1352 B.n132 B.n92 71.676
R1353 B.n128 B.n91 71.676
R1354 B.n124 B.n90 71.676
R1355 B.n352 B.n351 71.676
R1356 B.n354 B.n348 71.676
R1357 B.n361 B.n360 71.676
R1358 B.n362 B.n346 71.676
R1359 B.n369 B.n368 71.676
R1360 B.n370 B.n344 71.676
R1361 B.n377 B.n376 71.676
R1362 B.n378 B.n342 71.676
R1363 B.n385 B.n384 71.676
R1364 B.n386 B.n340 71.676
R1365 B.n396 B.n395 71.676
R1366 B.n397 B.n338 71.676
R1367 B.n404 B.n403 71.676
R1368 B.n405 B.n336 71.676
R1369 B.n412 B.n411 71.676
R1370 B.n413 B.n332 71.676
R1371 B.n421 B.n420 71.676
R1372 B.n422 B.n330 71.676
R1373 B.n429 B.n428 71.676
R1374 B.n430 B.n328 71.676
R1375 B.n437 B.n436 71.676
R1376 B.n438 B.n326 71.676
R1377 B.n445 B.n444 71.676
R1378 B.n446 B.n324 71.676
R1379 B.n453 B.n452 71.676
R1380 B.n456 B.n455 71.676
R1381 B.n461 B.n316 69.9397
R1382 B.n467 B.n316 69.9397
R1383 B.n467 B.n312 69.9397
R1384 B.n473 B.n312 69.9397
R1385 B.n473 B.n307 69.9397
R1386 B.n479 B.n307 69.9397
R1387 B.n479 B.n308 69.9397
R1388 B.n485 B.n300 69.9397
R1389 B.n491 B.n300 69.9397
R1390 B.n491 B.n296 69.9397
R1391 B.n497 B.n296 69.9397
R1392 B.n497 B.n292 69.9397
R1393 B.n503 B.n292 69.9397
R1394 B.n503 B.n288 69.9397
R1395 B.n509 B.n288 69.9397
R1396 B.n509 B.n284 69.9397
R1397 B.n515 B.n284 69.9397
R1398 B.n521 B.n280 69.9397
R1399 B.n521 B.n276 69.9397
R1400 B.n527 B.n276 69.9397
R1401 B.n527 B.n272 69.9397
R1402 B.n533 B.n272 69.9397
R1403 B.n533 B.n268 69.9397
R1404 B.n539 B.n268 69.9397
R1405 B.n545 B.n264 69.9397
R1406 B.n545 B.n260 69.9397
R1407 B.n551 B.n260 69.9397
R1408 B.n551 B.n256 69.9397
R1409 B.n557 B.n256 69.9397
R1410 B.n557 B.n252 69.9397
R1411 B.n563 B.n252 69.9397
R1412 B.n569 B.n248 69.9397
R1413 B.n569 B.n244 69.9397
R1414 B.n575 B.n244 69.9397
R1415 B.n575 B.n240 69.9397
R1416 B.n581 B.n240 69.9397
R1417 B.n581 B.n236 69.9397
R1418 B.n587 B.n236 69.9397
R1419 B.n594 B.n232 69.9397
R1420 B.n594 B.n228 69.9397
R1421 B.n600 B.n228 69.9397
R1422 B.n600 B.n4 69.9397
R1423 B.n765 B.n4 69.9397
R1424 B.n765 B.n764 69.9397
R1425 B.n764 B.n763 69.9397
R1426 B.n763 B.n8 69.9397
R1427 B.n757 B.n8 69.9397
R1428 B.n757 B.n756 69.9397
R1429 B.n755 B.n15 69.9397
R1430 B.n749 B.n15 69.9397
R1431 B.n749 B.n748 69.9397
R1432 B.n748 B.n747 69.9397
R1433 B.n747 B.n22 69.9397
R1434 B.n741 B.n22 69.9397
R1435 B.n741 B.n740 69.9397
R1436 B.n739 B.n29 69.9397
R1437 B.n733 B.n29 69.9397
R1438 B.n733 B.n732 69.9397
R1439 B.n732 B.n731 69.9397
R1440 B.n731 B.n36 69.9397
R1441 B.n725 B.n36 69.9397
R1442 B.n725 B.n724 69.9397
R1443 B.n723 B.n43 69.9397
R1444 B.n717 B.n43 69.9397
R1445 B.n717 B.n716 69.9397
R1446 B.n716 B.n715 69.9397
R1447 B.n715 B.n50 69.9397
R1448 B.n709 B.n50 69.9397
R1449 B.n709 B.n708 69.9397
R1450 B.n707 B.n57 69.9397
R1451 B.n701 B.n57 69.9397
R1452 B.n701 B.n700 69.9397
R1453 B.n700 B.n699 69.9397
R1454 B.n699 B.n64 69.9397
R1455 B.n693 B.n64 69.9397
R1456 B.n693 B.n692 69.9397
R1457 B.n692 B.n691 69.9397
R1458 B.n691 B.n71 69.9397
R1459 B.n685 B.n71 69.9397
R1460 B.n684 B.n683 69.9397
R1461 B.n683 B.n78 69.9397
R1462 B.n677 B.n78 69.9397
R1463 B.n677 B.n676 69.9397
R1464 B.n676 B.n675 69.9397
R1465 B.n675 B.n85 69.9397
R1466 B.n669 B.n85 69.9397
R1467 B.n416 B.n334 59.5399
R1468 B.n392 B.n391 59.5399
R1469 B.n122 B.n121 59.5399
R1470 B.n119 B.n118 59.5399
R1471 B.n334 B.n333 52.3641
R1472 B.n391 B.n390 52.3641
R1473 B.n121 B.n120 52.3641
R1474 B.n118 B.n117 52.3641
R1475 B.n515 B.t0 42.1697
R1476 B.t6 B.n707 42.1697
R1477 B.t4 B.n232 40.1127
R1478 B.n756 B.t5 40.1127
R1479 B.n485 B.t16 38.0557
R1480 B.n539 B.t2 38.0557
R1481 B.t3 B.n723 38.0557
R1482 B.n685 B.t9 38.0557
R1483 B.t7 B.n248 35.9986
R1484 B.n740 B.t1 35.9986
R1485 B.n563 B.t7 33.9416
R1486 B.t1 B.n739 33.9416
R1487 B.n308 B.t16 31.8846
R1488 B.t2 B.n264 31.8846
R1489 B.n724 B.t3 31.8846
R1490 B.t9 B.n684 31.8846
R1491 B.n671 B.n87 31.0639
R1492 B.n665 B.n664 31.0639
R1493 B.n459 B.n458 31.0639
R1494 B.n463 B.n318 31.0639
R1495 B.n587 B.t4 29.8275
R1496 B.t5 B.n755 29.8275
R1497 B.t0 B.n280 27.7705
R1498 B.n708 B.t6 27.7705
R1499 B B.n767 18.0485
R1500 B.n123 B.n87 10.6151
R1501 B.n126 B.n123 10.6151
R1502 B.n127 B.n126 10.6151
R1503 B.n130 B.n127 10.6151
R1504 B.n131 B.n130 10.6151
R1505 B.n134 B.n131 10.6151
R1506 B.n135 B.n134 10.6151
R1507 B.n138 B.n135 10.6151
R1508 B.n139 B.n138 10.6151
R1509 B.n142 B.n139 10.6151
R1510 B.n143 B.n142 10.6151
R1511 B.n146 B.n143 10.6151
R1512 B.n147 B.n146 10.6151
R1513 B.n150 B.n147 10.6151
R1514 B.n151 B.n150 10.6151
R1515 B.n154 B.n151 10.6151
R1516 B.n155 B.n154 10.6151
R1517 B.n158 B.n155 10.6151
R1518 B.n159 B.n158 10.6151
R1519 B.n162 B.n159 10.6151
R1520 B.n163 B.n162 10.6151
R1521 B.n167 B.n166 10.6151
R1522 B.n170 B.n167 10.6151
R1523 B.n171 B.n170 10.6151
R1524 B.n174 B.n171 10.6151
R1525 B.n175 B.n174 10.6151
R1526 B.n178 B.n175 10.6151
R1527 B.n179 B.n178 10.6151
R1528 B.n182 B.n179 10.6151
R1529 B.n183 B.n182 10.6151
R1530 B.n187 B.n186 10.6151
R1531 B.n190 B.n187 10.6151
R1532 B.n191 B.n190 10.6151
R1533 B.n194 B.n191 10.6151
R1534 B.n195 B.n194 10.6151
R1535 B.n198 B.n195 10.6151
R1536 B.n199 B.n198 10.6151
R1537 B.n202 B.n199 10.6151
R1538 B.n203 B.n202 10.6151
R1539 B.n206 B.n203 10.6151
R1540 B.n207 B.n206 10.6151
R1541 B.n210 B.n207 10.6151
R1542 B.n211 B.n210 10.6151
R1543 B.n214 B.n211 10.6151
R1544 B.n215 B.n214 10.6151
R1545 B.n218 B.n215 10.6151
R1546 B.n219 B.n218 10.6151
R1547 B.n222 B.n219 10.6151
R1548 B.n224 B.n222 10.6151
R1549 B.n225 B.n224 10.6151
R1550 B.n665 B.n225 10.6151
R1551 B.n459 B.n314 10.6151
R1552 B.n469 B.n314 10.6151
R1553 B.n470 B.n469 10.6151
R1554 B.n471 B.n470 10.6151
R1555 B.n471 B.n305 10.6151
R1556 B.n481 B.n305 10.6151
R1557 B.n482 B.n481 10.6151
R1558 B.n483 B.n482 10.6151
R1559 B.n483 B.n298 10.6151
R1560 B.n493 B.n298 10.6151
R1561 B.n494 B.n493 10.6151
R1562 B.n495 B.n494 10.6151
R1563 B.n495 B.n290 10.6151
R1564 B.n505 B.n290 10.6151
R1565 B.n506 B.n505 10.6151
R1566 B.n507 B.n506 10.6151
R1567 B.n507 B.n282 10.6151
R1568 B.n517 B.n282 10.6151
R1569 B.n518 B.n517 10.6151
R1570 B.n519 B.n518 10.6151
R1571 B.n519 B.n274 10.6151
R1572 B.n529 B.n274 10.6151
R1573 B.n530 B.n529 10.6151
R1574 B.n531 B.n530 10.6151
R1575 B.n531 B.n266 10.6151
R1576 B.n541 B.n266 10.6151
R1577 B.n542 B.n541 10.6151
R1578 B.n543 B.n542 10.6151
R1579 B.n543 B.n258 10.6151
R1580 B.n553 B.n258 10.6151
R1581 B.n554 B.n553 10.6151
R1582 B.n555 B.n554 10.6151
R1583 B.n555 B.n250 10.6151
R1584 B.n565 B.n250 10.6151
R1585 B.n566 B.n565 10.6151
R1586 B.n567 B.n566 10.6151
R1587 B.n567 B.n242 10.6151
R1588 B.n577 B.n242 10.6151
R1589 B.n578 B.n577 10.6151
R1590 B.n579 B.n578 10.6151
R1591 B.n579 B.n234 10.6151
R1592 B.n589 B.n234 10.6151
R1593 B.n590 B.n589 10.6151
R1594 B.n592 B.n590 10.6151
R1595 B.n592 B.n591 10.6151
R1596 B.n591 B.n226 10.6151
R1597 B.n603 B.n226 10.6151
R1598 B.n604 B.n603 10.6151
R1599 B.n605 B.n604 10.6151
R1600 B.n606 B.n605 10.6151
R1601 B.n608 B.n606 10.6151
R1602 B.n609 B.n608 10.6151
R1603 B.n610 B.n609 10.6151
R1604 B.n611 B.n610 10.6151
R1605 B.n613 B.n611 10.6151
R1606 B.n614 B.n613 10.6151
R1607 B.n615 B.n614 10.6151
R1608 B.n616 B.n615 10.6151
R1609 B.n618 B.n616 10.6151
R1610 B.n619 B.n618 10.6151
R1611 B.n620 B.n619 10.6151
R1612 B.n621 B.n620 10.6151
R1613 B.n623 B.n621 10.6151
R1614 B.n624 B.n623 10.6151
R1615 B.n625 B.n624 10.6151
R1616 B.n626 B.n625 10.6151
R1617 B.n628 B.n626 10.6151
R1618 B.n629 B.n628 10.6151
R1619 B.n630 B.n629 10.6151
R1620 B.n631 B.n630 10.6151
R1621 B.n633 B.n631 10.6151
R1622 B.n634 B.n633 10.6151
R1623 B.n635 B.n634 10.6151
R1624 B.n636 B.n635 10.6151
R1625 B.n638 B.n636 10.6151
R1626 B.n639 B.n638 10.6151
R1627 B.n640 B.n639 10.6151
R1628 B.n641 B.n640 10.6151
R1629 B.n643 B.n641 10.6151
R1630 B.n644 B.n643 10.6151
R1631 B.n645 B.n644 10.6151
R1632 B.n646 B.n645 10.6151
R1633 B.n648 B.n646 10.6151
R1634 B.n649 B.n648 10.6151
R1635 B.n650 B.n649 10.6151
R1636 B.n651 B.n650 10.6151
R1637 B.n653 B.n651 10.6151
R1638 B.n654 B.n653 10.6151
R1639 B.n655 B.n654 10.6151
R1640 B.n656 B.n655 10.6151
R1641 B.n658 B.n656 10.6151
R1642 B.n659 B.n658 10.6151
R1643 B.n660 B.n659 10.6151
R1644 B.n661 B.n660 10.6151
R1645 B.n663 B.n661 10.6151
R1646 B.n664 B.n663 10.6151
R1647 B.n350 B.n318 10.6151
R1648 B.n350 B.n349 10.6151
R1649 B.n356 B.n349 10.6151
R1650 B.n357 B.n356 10.6151
R1651 B.n358 B.n357 10.6151
R1652 B.n358 B.n347 10.6151
R1653 B.n364 B.n347 10.6151
R1654 B.n365 B.n364 10.6151
R1655 B.n366 B.n365 10.6151
R1656 B.n366 B.n345 10.6151
R1657 B.n372 B.n345 10.6151
R1658 B.n373 B.n372 10.6151
R1659 B.n374 B.n373 10.6151
R1660 B.n374 B.n343 10.6151
R1661 B.n380 B.n343 10.6151
R1662 B.n381 B.n380 10.6151
R1663 B.n382 B.n381 10.6151
R1664 B.n382 B.n341 10.6151
R1665 B.n388 B.n341 10.6151
R1666 B.n389 B.n388 10.6151
R1667 B.n393 B.n389 10.6151
R1668 B.n399 B.n339 10.6151
R1669 B.n400 B.n399 10.6151
R1670 B.n401 B.n400 10.6151
R1671 B.n401 B.n337 10.6151
R1672 B.n407 B.n337 10.6151
R1673 B.n408 B.n407 10.6151
R1674 B.n409 B.n408 10.6151
R1675 B.n409 B.n335 10.6151
R1676 B.n415 B.n335 10.6151
R1677 B.n418 B.n417 10.6151
R1678 B.n418 B.n331 10.6151
R1679 B.n424 B.n331 10.6151
R1680 B.n425 B.n424 10.6151
R1681 B.n426 B.n425 10.6151
R1682 B.n426 B.n329 10.6151
R1683 B.n432 B.n329 10.6151
R1684 B.n433 B.n432 10.6151
R1685 B.n434 B.n433 10.6151
R1686 B.n434 B.n327 10.6151
R1687 B.n440 B.n327 10.6151
R1688 B.n441 B.n440 10.6151
R1689 B.n442 B.n441 10.6151
R1690 B.n442 B.n325 10.6151
R1691 B.n448 B.n325 10.6151
R1692 B.n449 B.n448 10.6151
R1693 B.n450 B.n449 10.6151
R1694 B.n450 B.n323 10.6151
R1695 B.n323 B.n322 10.6151
R1696 B.n457 B.n322 10.6151
R1697 B.n458 B.n457 10.6151
R1698 B.n464 B.n463 10.6151
R1699 B.n465 B.n464 10.6151
R1700 B.n465 B.n310 10.6151
R1701 B.n475 B.n310 10.6151
R1702 B.n476 B.n475 10.6151
R1703 B.n477 B.n476 10.6151
R1704 B.n477 B.n302 10.6151
R1705 B.n487 B.n302 10.6151
R1706 B.n488 B.n487 10.6151
R1707 B.n489 B.n488 10.6151
R1708 B.n489 B.n294 10.6151
R1709 B.n499 B.n294 10.6151
R1710 B.n500 B.n499 10.6151
R1711 B.n501 B.n500 10.6151
R1712 B.n501 B.n286 10.6151
R1713 B.n511 B.n286 10.6151
R1714 B.n512 B.n511 10.6151
R1715 B.n513 B.n512 10.6151
R1716 B.n513 B.n278 10.6151
R1717 B.n523 B.n278 10.6151
R1718 B.n524 B.n523 10.6151
R1719 B.n525 B.n524 10.6151
R1720 B.n525 B.n270 10.6151
R1721 B.n535 B.n270 10.6151
R1722 B.n536 B.n535 10.6151
R1723 B.n537 B.n536 10.6151
R1724 B.n537 B.n262 10.6151
R1725 B.n547 B.n262 10.6151
R1726 B.n548 B.n547 10.6151
R1727 B.n549 B.n548 10.6151
R1728 B.n549 B.n254 10.6151
R1729 B.n559 B.n254 10.6151
R1730 B.n560 B.n559 10.6151
R1731 B.n561 B.n560 10.6151
R1732 B.n561 B.n246 10.6151
R1733 B.n571 B.n246 10.6151
R1734 B.n572 B.n571 10.6151
R1735 B.n573 B.n572 10.6151
R1736 B.n573 B.n238 10.6151
R1737 B.n583 B.n238 10.6151
R1738 B.n584 B.n583 10.6151
R1739 B.n585 B.n584 10.6151
R1740 B.n585 B.n230 10.6151
R1741 B.n596 B.n230 10.6151
R1742 B.n597 B.n596 10.6151
R1743 B.n598 B.n597 10.6151
R1744 B.n598 B.n0 10.6151
R1745 B.n761 B.n1 10.6151
R1746 B.n761 B.n760 10.6151
R1747 B.n760 B.n759 10.6151
R1748 B.n759 B.n10 10.6151
R1749 B.n753 B.n10 10.6151
R1750 B.n753 B.n752 10.6151
R1751 B.n752 B.n751 10.6151
R1752 B.n751 B.n17 10.6151
R1753 B.n745 B.n17 10.6151
R1754 B.n745 B.n744 10.6151
R1755 B.n744 B.n743 10.6151
R1756 B.n743 B.n24 10.6151
R1757 B.n737 B.n24 10.6151
R1758 B.n737 B.n736 10.6151
R1759 B.n736 B.n735 10.6151
R1760 B.n735 B.n31 10.6151
R1761 B.n729 B.n31 10.6151
R1762 B.n729 B.n728 10.6151
R1763 B.n728 B.n727 10.6151
R1764 B.n727 B.n38 10.6151
R1765 B.n721 B.n38 10.6151
R1766 B.n721 B.n720 10.6151
R1767 B.n720 B.n719 10.6151
R1768 B.n719 B.n45 10.6151
R1769 B.n713 B.n45 10.6151
R1770 B.n713 B.n712 10.6151
R1771 B.n712 B.n711 10.6151
R1772 B.n711 B.n52 10.6151
R1773 B.n705 B.n52 10.6151
R1774 B.n705 B.n704 10.6151
R1775 B.n704 B.n703 10.6151
R1776 B.n703 B.n59 10.6151
R1777 B.n697 B.n59 10.6151
R1778 B.n697 B.n696 10.6151
R1779 B.n696 B.n695 10.6151
R1780 B.n695 B.n66 10.6151
R1781 B.n689 B.n66 10.6151
R1782 B.n689 B.n688 10.6151
R1783 B.n688 B.n687 10.6151
R1784 B.n687 B.n73 10.6151
R1785 B.n681 B.n73 10.6151
R1786 B.n681 B.n680 10.6151
R1787 B.n680 B.n679 10.6151
R1788 B.n679 B.n80 10.6151
R1789 B.n673 B.n80 10.6151
R1790 B.n673 B.n672 10.6151
R1791 B.n672 B.n671 10.6151
R1792 B.n163 B.n122 9.36635
R1793 B.n186 B.n119 9.36635
R1794 B.n393 B.n392 9.36635
R1795 B.n417 B.n416 9.36635
R1796 B.n767 B.n0 2.81026
R1797 B.n767 B.n1 2.81026
R1798 B.n166 B.n122 1.24928
R1799 B.n183 B.n119 1.24928
R1800 B.n392 B.n339 1.24928
R1801 B.n416 B.n415 1.24928
R1802 VP.n16 VP.n13 161.3
R1803 VP.n18 VP.n17 161.3
R1804 VP.n19 VP.n12 161.3
R1805 VP.n21 VP.n20 161.3
R1806 VP.n22 VP.n11 161.3
R1807 VP.n24 VP.n23 161.3
R1808 VP.n26 VP.n10 161.3
R1809 VP.n28 VP.n27 161.3
R1810 VP.n29 VP.n9 161.3
R1811 VP.n31 VP.n30 161.3
R1812 VP.n32 VP.n8 161.3
R1813 VP.n62 VP.n0 161.3
R1814 VP.n61 VP.n60 161.3
R1815 VP.n59 VP.n1 161.3
R1816 VP.n58 VP.n57 161.3
R1817 VP.n56 VP.n2 161.3
R1818 VP.n54 VP.n53 161.3
R1819 VP.n52 VP.n3 161.3
R1820 VP.n51 VP.n50 161.3
R1821 VP.n49 VP.n4 161.3
R1822 VP.n48 VP.n47 161.3
R1823 VP.n46 VP.n5 161.3
R1824 VP.n45 VP.n44 161.3
R1825 VP.n42 VP.n6 161.3
R1826 VP.n41 VP.n40 161.3
R1827 VP.n39 VP.n7 161.3
R1828 VP.n38 VP.n37 161.3
R1829 VP.n36 VP.n35 96.1531
R1830 VP.n64 VP.n63 96.1531
R1831 VP.n34 VP.n33 96.1531
R1832 VP.n15 VP.t3 87.6179
R1833 VP.n15 VP.n14 67.4531
R1834 VP.n50 VP.n49 56.5617
R1835 VP.n20 VP.n19 56.5617
R1836 VP.n36 VP.t7 55.1153
R1837 VP.n43 VP.t2 55.1153
R1838 VP.n55 VP.t4 55.1153
R1839 VP.n63 VP.t0 55.1153
R1840 VP.n33 VP.t5 55.1153
R1841 VP.n25 VP.t1 55.1153
R1842 VP.n14 VP.t6 55.1153
R1843 VP.n42 VP.n41 45.4209
R1844 VP.n57 VP.n1 45.4209
R1845 VP.n27 VP.n9 45.4209
R1846 VP.n35 VP.n34 44.8709
R1847 VP.n41 VP.n7 35.7332
R1848 VP.n61 VP.n1 35.7332
R1849 VP.n31 VP.n9 35.7332
R1850 VP.n37 VP.n7 24.5923
R1851 VP.n44 VP.n42 24.5923
R1852 VP.n48 VP.n5 24.5923
R1853 VP.n49 VP.n48 24.5923
R1854 VP.n50 VP.n3 24.5923
R1855 VP.n54 VP.n3 24.5923
R1856 VP.n57 VP.n56 24.5923
R1857 VP.n62 VP.n61 24.5923
R1858 VP.n32 VP.n31 24.5923
R1859 VP.n20 VP.n11 24.5923
R1860 VP.n24 VP.n11 24.5923
R1861 VP.n27 VP.n26 24.5923
R1862 VP.n18 VP.n13 24.5923
R1863 VP.n19 VP.n18 24.5923
R1864 VP.n44 VP.n43 19.674
R1865 VP.n56 VP.n55 19.674
R1866 VP.n26 VP.n25 19.674
R1867 VP.n37 VP.n36 14.7556
R1868 VP.n63 VP.n62 14.7556
R1869 VP.n33 VP.n32 14.7556
R1870 VP.n16 VP.n15 9.50446
R1871 VP.n43 VP.n5 4.91887
R1872 VP.n55 VP.n54 4.91887
R1873 VP.n25 VP.n24 4.91887
R1874 VP.n14 VP.n13 4.91887
R1875 VP.n34 VP.n8 0.278335
R1876 VP.n38 VP.n35 0.278335
R1877 VP.n64 VP.n0 0.278335
R1878 VP.n17 VP.n16 0.189894
R1879 VP.n17 VP.n12 0.189894
R1880 VP.n21 VP.n12 0.189894
R1881 VP.n22 VP.n21 0.189894
R1882 VP.n23 VP.n22 0.189894
R1883 VP.n23 VP.n10 0.189894
R1884 VP.n28 VP.n10 0.189894
R1885 VP.n29 VP.n28 0.189894
R1886 VP.n30 VP.n29 0.189894
R1887 VP.n30 VP.n8 0.189894
R1888 VP.n39 VP.n38 0.189894
R1889 VP.n40 VP.n39 0.189894
R1890 VP.n40 VP.n6 0.189894
R1891 VP.n45 VP.n6 0.189894
R1892 VP.n46 VP.n45 0.189894
R1893 VP.n47 VP.n46 0.189894
R1894 VP.n47 VP.n4 0.189894
R1895 VP.n51 VP.n4 0.189894
R1896 VP.n52 VP.n51 0.189894
R1897 VP.n53 VP.n52 0.189894
R1898 VP.n53 VP.n2 0.189894
R1899 VP.n58 VP.n2 0.189894
R1900 VP.n59 VP.n58 0.189894
R1901 VP.n60 VP.n59 0.189894
R1902 VP.n60 VP.n0 0.189894
R1903 VP VP.n64 0.153485
R1904 VDD1 VDD1.n0 72.5924
R1905 VDD1.n3 VDD1.n2 72.4787
R1906 VDD1.n3 VDD1.n1 72.4787
R1907 VDD1.n5 VDD1.n4 71.3703
R1908 VDD1.n5 VDD1.n3 39.4449
R1909 VDD1.n4 VDD1.t6 3.65364
R1910 VDD1.n4 VDD1.t2 3.65364
R1911 VDD1.n0 VDD1.t4 3.65364
R1912 VDD1.n0 VDD1.t1 3.65364
R1913 VDD1.n2 VDD1.t3 3.65364
R1914 VDD1.n2 VDD1.t7 3.65364
R1915 VDD1.n1 VDD1.t0 3.65364
R1916 VDD1.n1 VDD1.t5 3.65364
R1917 VDD1 VDD1.n5 1.1061
C0 VP VDD2 0.499104f
C1 VN VTAIL 4.87013f
C2 VN VDD1 0.151319f
C3 VDD1 VTAIL 5.72367f
C4 VN VDD2 4.10465f
C5 VDD2 VTAIL 5.77655f
C6 VDD2 VDD1 1.65542f
C7 VP VN 6.1565f
C8 VP VTAIL 4.88424f
C9 VP VDD1 4.44721f
C10 VDD2 B 4.599407f
C11 VDD1 B 5.015725f
C12 VTAIL B 6.053076f
C13 VN B 13.95651f
C14 VP B 12.558646f
C15 VDD1.t4 B 0.105473f
C16 VDD1.t1 B 0.105473f
C17 VDD1.n0 B 0.876982f
C18 VDD1.t0 B 0.105473f
C19 VDD1.t5 B 0.105473f
C20 VDD1.n1 B 0.876094f
C21 VDD1.t3 B 0.105473f
C22 VDD1.t7 B 0.105473f
C23 VDD1.n2 B 0.876094f
C24 VDD1.n3 B 2.74324f
C25 VDD1.t6 B 0.105473f
C26 VDD1.t2 B 0.105473f
C27 VDD1.n4 B 0.868745f
C28 VDD1.n5 B 2.34953f
C29 VP.n0 B 0.035864f
C30 VP.t0 B 0.919103f
C31 VP.n1 B 0.022852f
C32 VP.n2 B 0.027205f
C33 VP.t4 B 0.919103f
C34 VP.n3 B 0.050448f
C35 VP.n4 B 0.027205f
C36 VP.n5 B 0.030524f
C37 VP.n6 B 0.027205f
C38 VP.n7 B 0.054642f
C39 VP.n8 B 0.035864f
C40 VP.t5 B 0.919103f
C41 VP.n9 B 0.022852f
C42 VP.n10 B 0.027205f
C43 VP.t1 B 0.919103f
C44 VP.n11 B 0.050448f
C45 VP.n12 B 0.027205f
C46 VP.n13 B 0.030524f
C47 VP.t3 B 1.10636f
C48 VP.t6 B 0.919103f
C49 VP.n14 B 0.418052f
C50 VP.n15 B 0.411596f
C51 VP.n16 B 0.236171f
C52 VP.n17 B 0.027205f
C53 VP.n18 B 0.050448f
C54 VP.n19 B 0.039546f
C55 VP.n20 B 0.039546f
C56 VP.n21 B 0.027205f
C57 VP.n22 B 0.027205f
C58 VP.n23 B 0.027205f
C59 VP.n24 B 0.030524f
C60 VP.n25 B 0.351349f
C61 VP.n26 B 0.045467f
C62 VP.n27 B 0.052047f
C63 VP.n28 B 0.027205f
C64 VP.n29 B 0.027205f
C65 VP.n30 B 0.027205f
C66 VP.n31 B 0.054642f
C67 VP.n32 B 0.040486f
C68 VP.n33 B 0.440754f
C69 VP.n34 B 1.28024f
C70 VP.n35 B 1.3021f
C71 VP.t7 B 0.919103f
C72 VP.n36 B 0.440754f
C73 VP.n37 B 0.040486f
C74 VP.n38 B 0.035864f
C75 VP.n39 B 0.027205f
C76 VP.n40 B 0.027205f
C77 VP.n41 B 0.022852f
C78 VP.n42 B 0.052047f
C79 VP.t2 B 0.919103f
C80 VP.n43 B 0.351349f
C81 VP.n44 B 0.045467f
C82 VP.n45 B 0.027205f
C83 VP.n46 B 0.027205f
C84 VP.n47 B 0.027205f
C85 VP.n48 B 0.050448f
C86 VP.n49 B 0.039546f
C87 VP.n50 B 0.039546f
C88 VP.n51 B 0.027205f
C89 VP.n52 B 0.027205f
C90 VP.n53 B 0.027205f
C91 VP.n54 B 0.030524f
C92 VP.n55 B 0.351349f
C93 VP.n56 B 0.045467f
C94 VP.n57 B 0.052047f
C95 VP.n58 B 0.027205f
C96 VP.n59 B 0.027205f
C97 VP.n60 B 0.027205f
C98 VP.n61 B 0.054642f
C99 VP.n62 B 0.040486f
C100 VP.n63 B 0.440754f
C101 VP.n64 B 0.039046f
C102 VDD2.t3 B 0.104324f
C103 VDD2.t7 B 0.104324f
C104 VDD2.n0 B 0.86655f
C105 VDD2.t2 B 0.104324f
C106 VDD2.t5 B 0.104324f
C107 VDD2.n1 B 0.86655f
C108 VDD2.n2 B 2.6623f
C109 VDD2.t4 B 0.104324f
C110 VDD2.t0 B 0.104324f
C111 VDD2.n3 B 0.859284f
C112 VDD2.n4 B 2.29415f
C113 VDD2.t6 B 0.104324f
C114 VDD2.t1 B 0.104324f
C115 VDD2.n5 B 0.86652f
C116 VTAIL.t10 B 0.101186f
C117 VTAIL.t6 B 0.101186f
C118 VTAIL.n0 B 0.777024f
C119 VTAIL.n1 B 0.395395f
C120 VTAIL.n2 B 0.034801f
C121 VTAIL.n3 B 0.023625f
C122 VTAIL.n4 B 0.012695f
C123 VTAIL.n5 B 0.030006f
C124 VTAIL.n6 B 0.013442f
C125 VTAIL.n7 B 0.023625f
C126 VTAIL.n8 B 0.012695f
C127 VTAIL.n9 B 0.022505f
C128 VTAIL.n10 B 0.017721f
C129 VTAIL.t5 B 0.049082f
C130 VTAIL.n11 B 0.098099f
C131 VTAIL.n12 B 0.498674f
C132 VTAIL.n13 B 0.012695f
C133 VTAIL.n14 B 0.013442f
C134 VTAIL.n15 B 0.030006f
C135 VTAIL.n16 B 0.030006f
C136 VTAIL.n17 B 0.013442f
C137 VTAIL.n18 B 0.012695f
C138 VTAIL.n19 B 0.023625f
C139 VTAIL.n20 B 0.023625f
C140 VTAIL.n21 B 0.012695f
C141 VTAIL.n22 B 0.013442f
C142 VTAIL.n23 B 0.030006f
C143 VTAIL.n24 B 0.067777f
C144 VTAIL.n25 B 0.013442f
C145 VTAIL.n26 B 0.012695f
C146 VTAIL.n27 B 0.059126f
C147 VTAIL.n28 B 0.038348f
C148 VTAIL.n29 B 0.235683f
C149 VTAIL.n30 B 0.034801f
C150 VTAIL.n31 B 0.023625f
C151 VTAIL.n32 B 0.012695f
C152 VTAIL.n33 B 0.030006f
C153 VTAIL.n34 B 0.013442f
C154 VTAIL.n35 B 0.023625f
C155 VTAIL.n36 B 0.012695f
C156 VTAIL.n37 B 0.022505f
C157 VTAIL.n38 B 0.017721f
C158 VTAIL.t4 B 0.049082f
C159 VTAIL.n39 B 0.098099f
C160 VTAIL.n40 B 0.498674f
C161 VTAIL.n41 B 0.012695f
C162 VTAIL.n42 B 0.013442f
C163 VTAIL.n43 B 0.030006f
C164 VTAIL.n44 B 0.030006f
C165 VTAIL.n45 B 0.013442f
C166 VTAIL.n46 B 0.012695f
C167 VTAIL.n47 B 0.023625f
C168 VTAIL.n48 B 0.023625f
C169 VTAIL.n49 B 0.012695f
C170 VTAIL.n50 B 0.013442f
C171 VTAIL.n51 B 0.030006f
C172 VTAIL.n52 B 0.067777f
C173 VTAIL.n53 B 0.013442f
C174 VTAIL.n54 B 0.012695f
C175 VTAIL.n55 B 0.059126f
C176 VTAIL.n56 B 0.038348f
C177 VTAIL.n57 B 0.235683f
C178 VTAIL.t2 B 0.101186f
C179 VTAIL.t15 B 0.101186f
C180 VTAIL.n58 B 0.777024f
C181 VTAIL.n59 B 0.568151f
C182 VTAIL.n60 B 0.034801f
C183 VTAIL.n61 B 0.023625f
C184 VTAIL.n62 B 0.012695f
C185 VTAIL.n63 B 0.030006f
C186 VTAIL.n64 B 0.013442f
C187 VTAIL.n65 B 0.023625f
C188 VTAIL.n66 B 0.012695f
C189 VTAIL.n67 B 0.022505f
C190 VTAIL.n68 B 0.017721f
C191 VTAIL.t0 B 0.049082f
C192 VTAIL.n69 B 0.098099f
C193 VTAIL.n70 B 0.498674f
C194 VTAIL.n71 B 0.012695f
C195 VTAIL.n72 B 0.013442f
C196 VTAIL.n73 B 0.030006f
C197 VTAIL.n74 B 0.030006f
C198 VTAIL.n75 B 0.013442f
C199 VTAIL.n76 B 0.012695f
C200 VTAIL.n77 B 0.023625f
C201 VTAIL.n78 B 0.023625f
C202 VTAIL.n79 B 0.012695f
C203 VTAIL.n80 B 0.013442f
C204 VTAIL.n81 B 0.030006f
C205 VTAIL.n82 B 0.067777f
C206 VTAIL.n83 B 0.013442f
C207 VTAIL.n84 B 0.012695f
C208 VTAIL.n85 B 0.059126f
C209 VTAIL.n86 B 0.038348f
C210 VTAIL.n87 B 1.0537f
C211 VTAIL.n88 B 0.034801f
C212 VTAIL.n89 B 0.023625f
C213 VTAIL.n90 B 0.012695f
C214 VTAIL.n91 B 0.030006f
C215 VTAIL.n92 B 0.013442f
C216 VTAIL.n93 B 0.023625f
C217 VTAIL.n94 B 0.012695f
C218 VTAIL.n95 B 0.022505f
C219 VTAIL.n96 B 0.017721f
C220 VTAIL.t12 B 0.049082f
C221 VTAIL.n97 B 0.098099f
C222 VTAIL.n98 B 0.498674f
C223 VTAIL.n99 B 0.012695f
C224 VTAIL.n100 B 0.013442f
C225 VTAIL.n101 B 0.030006f
C226 VTAIL.n102 B 0.030006f
C227 VTAIL.n103 B 0.013442f
C228 VTAIL.n104 B 0.012695f
C229 VTAIL.n105 B 0.023625f
C230 VTAIL.n106 B 0.023625f
C231 VTAIL.n107 B 0.012695f
C232 VTAIL.n108 B 0.013442f
C233 VTAIL.n109 B 0.030006f
C234 VTAIL.n110 B 0.067777f
C235 VTAIL.n111 B 0.013442f
C236 VTAIL.n112 B 0.012695f
C237 VTAIL.n113 B 0.059126f
C238 VTAIL.n114 B 0.038348f
C239 VTAIL.n115 B 1.0537f
C240 VTAIL.t9 B 0.101186f
C241 VTAIL.t11 B 0.101186f
C242 VTAIL.n116 B 0.777029f
C243 VTAIL.n117 B 0.568146f
C244 VTAIL.n118 B 0.034801f
C245 VTAIL.n119 B 0.023625f
C246 VTAIL.n120 B 0.012695f
C247 VTAIL.n121 B 0.030006f
C248 VTAIL.n122 B 0.013442f
C249 VTAIL.n123 B 0.023625f
C250 VTAIL.n124 B 0.012695f
C251 VTAIL.n125 B 0.022505f
C252 VTAIL.n126 B 0.017721f
C253 VTAIL.t7 B 0.049082f
C254 VTAIL.n127 B 0.098099f
C255 VTAIL.n128 B 0.498674f
C256 VTAIL.n129 B 0.012695f
C257 VTAIL.n130 B 0.013442f
C258 VTAIL.n131 B 0.030006f
C259 VTAIL.n132 B 0.030006f
C260 VTAIL.n133 B 0.013442f
C261 VTAIL.n134 B 0.012695f
C262 VTAIL.n135 B 0.023625f
C263 VTAIL.n136 B 0.023625f
C264 VTAIL.n137 B 0.012695f
C265 VTAIL.n138 B 0.013442f
C266 VTAIL.n139 B 0.030006f
C267 VTAIL.n140 B 0.067777f
C268 VTAIL.n141 B 0.013442f
C269 VTAIL.n142 B 0.012695f
C270 VTAIL.n143 B 0.059126f
C271 VTAIL.n144 B 0.038348f
C272 VTAIL.n145 B 0.235683f
C273 VTAIL.n146 B 0.034801f
C274 VTAIL.n147 B 0.023625f
C275 VTAIL.n148 B 0.012695f
C276 VTAIL.n149 B 0.030006f
C277 VTAIL.n150 B 0.013442f
C278 VTAIL.n151 B 0.023625f
C279 VTAIL.n152 B 0.012695f
C280 VTAIL.n153 B 0.022505f
C281 VTAIL.n154 B 0.017721f
C282 VTAIL.t13 B 0.049082f
C283 VTAIL.n155 B 0.098099f
C284 VTAIL.n156 B 0.498674f
C285 VTAIL.n157 B 0.012695f
C286 VTAIL.n158 B 0.013442f
C287 VTAIL.n159 B 0.030006f
C288 VTAIL.n160 B 0.030006f
C289 VTAIL.n161 B 0.013442f
C290 VTAIL.n162 B 0.012695f
C291 VTAIL.n163 B 0.023625f
C292 VTAIL.n164 B 0.023625f
C293 VTAIL.n165 B 0.012695f
C294 VTAIL.n166 B 0.013442f
C295 VTAIL.n167 B 0.030006f
C296 VTAIL.n168 B 0.067777f
C297 VTAIL.n169 B 0.013442f
C298 VTAIL.n170 B 0.012695f
C299 VTAIL.n171 B 0.059126f
C300 VTAIL.n172 B 0.038348f
C301 VTAIL.n173 B 0.235683f
C302 VTAIL.t1 B 0.101186f
C303 VTAIL.t3 B 0.101186f
C304 VTAIL.n174 B 0.777029f
C305 VTAIL.n175 B 0.568146f
C306 VTAIL.n176 B 0.034801f
C307 VTAIL.n177 B 0.023625f
C308 VTAIL.n178 B 0.012695f
C309 VTAIL.n179 B 0.030006f
C310 VTAIL.n180 B 0.013442f
C311 VTAIL.n181 B 0.023625f
C312 VTAIL.n182 B 0.012695f
C313 VTAIL.n183 B 0.022505f
C314 VTAIL.n184 B 0.017721f
C315 VTAIL.t14 B 0.049082f
C316 VTAIL.n185 B 0.098099f
C317 VTAIL.n186 B 0.498674f
C318 VTAIL.n187 B 0.012695f
C319 VTAIL.n188 B 0.013442f
C320 VTAIL.n189 B 0.030006f
C321 VTAIL.n190 B 0.030006f
C322 VTAIL.n191 B 0.013442f
C323 VTAIL.n192 B 0.012695f
C324 VTAIL.n193 B 0.023625f
C325 VTAIL.n194 B 0.023625f
C326 VTAIL.n195 B 0.012695f
C327 VTAIL.n196 B 0.013442f
C328 VTAIL.n197 B 0.030006f
C329 VTAIL.n198 B 0.067777f
C330 VTAIL.n199 B 0.013442f
C331 VTAIL.n200 B 0.012695f
C332 VTAIL.n201 B 0.059126f
C333 VTAIL.n202 B 0.038348f
C334 VTAIL.n203 B 1.0537f
C335 VTAIL.n204 B 0.034801f
C336 VTAIL.n205 B 0.023625f
C337 VTAIL.n206 B 0.012695f
C338 VTAIL.n207 B 0.030006f
C339 VTAIL.n208 B 0.013442f
C340 VTAIL.n209 B 0.023625f
C341 VTAIL.n210 B 0.012695f
C342 VTAIL.n211 B 0.022505f
C343 VTAIL.n212 B 0.017721f
C344 VTAIL.t8 B 0.049082f
C345 VTAIL.n213 B 0.098099f
C346 VTAIL.n214 B 0.498674f
C347 VTAIL.n215 B 0.012695f
C348 VTAIL.n216 B 0.013442f
C349 VTAIL.n217 B 0.030006f
C350 VTAIL.n218 B 0.030006f
C351 VTAIL.n219 B 0.013442f
C352 VTAIL.n220 B 0.012695f
C353 VTAIL.n221 B 0.023625f
C354 VTAIL.n222 B 0.023625f
C355 VTAIL.n223 B 0.012695f
C356 VTAIL.n224 B 0.013442f
C357 VTAIL.n225 B 0.030006f
C358 VTAIL.n226 B 0.067777f
C359 VTAIL.n227 B 0.013442f
C360 VTAIL.n228 B 0.012695f
C361 VTAIL.n229 B 0.059126f
C362 VTAIL.n230 B 0.038348f
C363 VTAIL.n231 B 1.04927f
C364 VN.n0 B 0.035084f
C365 VN.t2 B 0.899096f
C366 VN.n1 B 0.022354f
C367 VN.n2 B 0.026612f
C368 VN.t5 B 0.899096f
C369 VN.n3 B 0.04935f
C370 VN.n4 B 0.026612f
C371 VN.n5 B 0.02986f
C372 VN.t4 B 1.08228f
C373 VN.t0 B 0.899096f
C374 VN.n6 B 0.408951f
C375 VN.n7 B 0.402636f
C376 VN.n8 B 0.23103f
C377 VN.n9 B 0.026612f
C378 VN.n10 B 0.04935f
C379 VN.n11 B 0.038685f
C380 VN.n12 B 0.038685f
C381 VN.n13 B 0.026612f
C382 VN.n14 B 0.026612f
C383 VN.n15 B 0.026612f
C384 VN.n16 B 0.02986f
C385 VN.n17 B 0.343701f
C386 VN.n18 B 0.044478f
C387 VN.n19 B 0.050914f
C388 VN.n20 B 0.026612f
C389 VN.n21 B 0.026612f
C390 VN.n22 B 0.026612f
C391 VN.n23 B 0.053452f
C392 VN.n24 B 0.039605f
C393 VN.n25 B 0.43116f
C394 VN.n26 B 0.038196f
C395 VN.n27 B 0.035084f
C396 VN.t3 B 0.899096f
C397 VN.n28 B 0.022354f
C398 VN.n29 B 0.026612f
C399 VN.t7 B 0.899096f
C400 VN.n30 B 0.04935f
C401 VN.n31 B 0.026612f
C402 VN.n32 B 0.02986f
C403 VN.t6 B 1.08228f
C404 VN.t1 B 0.899096f
C405 VN.n33 B 0.408951f
C406 VN.n34 B 0.402636f
C407 VN.n35 B 0.23103f
C408 VN.n36 B 0.026612f
C409 VN.n37 B 0.04935f
C410 VN.n38 B 0.038685f
C411 VN.n39 B 0.038685f
C412 VN.n40 B 0.026612f
C413 VN.n41 B 0.026612f
C414 VN.n42 B 0.026612f
C415 VN.n43 B 0.02986f
C416 VN.n44 B 0.343701f
C417 VN.n45 B 0.044478f
C418 VN.n46 B 0.050914f
C419 VN.n47 B 0.026612f
C420 VN.n48 B 0.026612f
C421 VN.n49 B 0.026612f
C422 VN.n50 B 0.053452f
C423 VN.n51 B 0.039605f
C424 VN.n52 B 0.43116f
C425 VN.n53 B 1.26693f
.ends

