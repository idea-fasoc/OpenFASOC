* NGSPICE file created from diff_pair_sample_0224.ext - technology: sky130A

.subckt diff_pair_sample_0224 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X1 VDD1.t9 VP.t0 VTAIL.t19 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X2 VTAIL.t18 VN.t1 VDD2.t8 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X3 VTAIL.t2 VP.t1 VDD1.t8 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X4 VDD1.t7 VP.t2 VTAIL.t5 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=4
X5 VTAIL.t7 VP.t3 VDD1.t6 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X6 VTAIL.t0 VP.t4 VDD1.t5 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X7 VDD2.t7 VN.t2 VTAIL.t11 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=4
X8 VDD1.t4 VP.t5 VTAIL.t1 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=4
X9 VDD2.t6 VN.t3 VTAIL.t16 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=4
X10 VDD2.t5 VN.t4 VTAIL.t14 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X11 VDD2.t4 VN.t5 VTAIL.t17 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=4
X12 B.t11 B.t9 B.t10 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=4
X13 B.t8 B.t6 B.t7 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=4
X14 B.t5 B.t3 B.t4 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=4
X15 VDD2.t3 VN.t6 VTAIL.t9 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=4
X16 VTAIL.t12 VN.t7 VDD2.t2 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X17 B.t2 B.t0 B.t1 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=0 ps=0 w=9.05 l=4
X18 VTAIL.t13 VN.t8 VDD2.t1 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X19 VDD1.t3 VP.t6 VTAIL.t3 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=3.5295 pd=18.88 as=1.49325 ps=9.38 w=9.05 l=4
X20 VTAIL.t15 VN.t9 VDD2.t0 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X21 VDD1.t2 VP.t7 VTAIL.t4 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X22 VTAIL.t6 VP.t8 VDD1.t1 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=1.49325 ps=9.38 w=9.05 l=4
X23 VDD1.t0 VP.t9 VTAIL.t8 w_n6166_n2778# sky130_fd_pr__pfet_01v8 ad=1.49325 pd=9.38 as=3.5295 ps=18.88 w=9.05 l=4
R0 VN.n113 VN.n58 161.3
R1 VN.n112 VN.n111 161.3
R2 VN.n110 VN.n59 161.3
R3 VN.n109 VN.n108 161.3
R4 VN.n107 VN.n60 161.3
R5 VN.n106 VN.n105 161.3
R6 VN.n104 VN.n61 161.3
R7 VN.n103 VN.n102 161.3
R8 VN.n100 VN.n62 161.3
R9 VN.n99 VN.n98 161.3
R10 VN.n97 VN.n63 161.3
R11 VN.n96 VN.n95 161.3
R12 VN.n94 VN.n64 161.3
R13 VN.n93 VN.n92 161.3
R14 VN.n91 VN.n65 161.3
R15 VN.n90 VN.n89 161.3
R16 VN.n88 VN.n66 161.3
R17 VN.n86 VN.n85 161.3
R18 VN.n84 VN.n67 161.3
R19 VN.n83 VN.n82 161.3
R20 VN.n81 VN.n68 161.3
R21 VN.n80 VN.n79 161.3
R22 VN.n78 VN.n69 161.3
R23 VN.n77 VN.n76 161.3
R24 VN.n75 VN.n70 161.3
R25 VN.n74 VN.n73 161.3
R26 VN.n55 VN.n0 161.3
R27 VN.n54 VN.n53 161.3
R28 VN.n52 VN.n1 161.3
R29 VN.n51 VN.n50 161.3
R30 VN.n49 VN.n2 161.3
R31 VN.n48 VN.n47 161.3
R32 VN.n46 VN.n3 161.3
R33 VN.n45 VN.n44 161.3
R34 VN.n42 VN.n4 161.3
R35 VN.n41 VN.n40 161.3
R36 VN.n39 VN.n5 161.3
R37 VN.n38 VN.n37 161.3
R38 VN.n36 VN.n6 161.3
R39 VN.n35 VN.n34 161.3
R40 VN.n33 VN.n7 161.3
R41 VN.n32 VN.n31 161.3
R42 VN.n30 VN.n8 161.3
R43 VN.n28 VN.n27 161.3
R44 VN.n26 VN.n9 161.3
R45 VN.n25 VN.n24 161.3
R46 VN.n23 VN.n10 161.3
R47 VN.n22 VN.n21 161.3
R48 VN.n20 VN.n11 161.3
R49 VN.n19 VN.n18 161.3
R50 VN.n17 VN.n12 161.3
R51 VN.n16 VN.n15 161.3
R52 VN.n14 VN.t5 86.7962
R53 VN.n72 VN.t3 86.7962
R54 VN.n14 VN.n13 71.1462
R55 VN.n72 VN.n71 71.1462
R56 VN.n57 VN.n56 62.1188
R57 VN.n115 VN.n114 62.1188
R58 VN VN.n115 58.7731
R59 VN.n50 VN.n49 56.5193
R60 VN.n108 VN.n107 56.5193
R61 VN.n13 VN.t8 54.5267
R62 VN.n29 VN.t4 54.5267
R63 VN.n43 VN.t7 54.5267
R64 VN.n56 VN.t6 54.5267
R65 VN.n71 VN.t9 54.5267
R66 VN.n87 VN.t0 54.5267
R67 VN.n101 VN.t1 54.5267
R68 VN.n114 VN.t2 54.5267
R69 VN.n23 VN.n22 48.7492
R70 VN.n36 VN.n35 48.7492
R71 VN.n81 VN.n80 48.7492
R72 VN.n94 VN.n93 48.7492
R73 VN.n22 VN.n11 32.2376
R74 VN.n37 VN.n36 32.2376
R75 VN.n80 VN.n69 32.2376
R76 VN.n95 VN.n94 32.2376
R77 VN.n17 VN.n16 24.4675
R78 VN.n18 VN.n17 24.4675
R79 VN.n18 VN.n11 24.4675
R80 VN.n24 VN.n23 24.4675
R81 VN.n24 VN.n9 24.4675
R82 VN.n28 VN.n9 24.4675
R83 VN.n31 VN.n30 24.4675
R84 VN.n31 VN.n7 24.4675
R85 VN.n35 VN.n7 24.4675
R86 VN.n37 VN.n5 24.4675
R87 VN.n41 VN.n5 24.4675
R88 VN.n42 VN.n41 24.4675
R89 VN.n44 VN.n3 24.4675
R90 VN.n48 VN.n3 24.4675
R91 VN.n49 VN.n48 24.4675
R92 VN.n50 VN.n1 24.4675
R93 VN.n54 VN.n1 24.4675
R94 VN.n55 VN.n54 24.4675
R95 VN.n76 VN.n69 24.4675
R96 VN.n76 VN.n75 24.4675
R97 VN.n75 VN.n74 24.4675
R98 VN.n93 VN.n65 24.4675
R99 VN.n89 VN.n65 24.4675
R100 VN.n89 VN.n88 24.4675
R101 VN.n86 VN.n67 24.4675
R102 VN.n82 VN.n67 24.4675
R103 VN.n82 VN.n81 24.4675
R104 VN.n107 VN.n106 24.4675
R105 VN.n106 VN.n61 24.4675
R106 VN.n102 VN.n61 24.4675
R107 VN.n100 VN.n99 24.4675
R108 VN.n99 VN.n63 24.4675
R109 VN.n95 VN.n63 24.4675
R110 VN.n113 VN.n112 24.4675
R111 VN.n112 VN.n59 24.4675
R112 VN.n108 VN.n59 24.4675
R113 VN.n44 VN.n43 20.5528
R114 VN.n102 VN.n101 20.5528
R115 VN.n56 VN.n55 20.0634
R116 VN.n114 VN.n113 20.0634
R117 VN.n29 VN.n28 12.234
R118 VN.n30 VN.n29 12.234
R119 VN.n88 VN.n87 12.234
R120 VN.n87 VN.n86 12.234
R121 VN.n16 VN.n13 3.91522
R122 VN.n43 VN.n42 3.91522
R123 VN.n74 VN.n71 3.91522
R124 VN.n101 VN.n100 3.91522
R125 VN.n73 VN.n72 2.69184
R126 VN.n15 VN.n14 2.69184
R127 VN.n115 VN.n58 0.417535
R128 VN.n57 VN.n0 0.417535
R129 VN VN.n57 0.394291
R130 VN.n111 VN.n58 0.189894
R131 VN.n111 VN.n110 0.189894
R132 VN.n110 VN.n109 0.189894
R133 VN.n109 VN.n60 0.189894
R134 VN.n105 VN.n60 0.189894
R135 VN.n105 VN.n104 0.189894
R136 VN.n104 VN.n103 0.189894
R137 VN.n103 VN.n62 0.189894
R138 VN.n98 VN.n62 0.189894
R139 VN.n98 VN.n97 0.189894
R140 VN.n97 VN.n96 0.189894
R141 VN.n96 VN.n64 0.189894
R142 VN.n92 VN.n64 0.189894
R143 VN.n92 VN.n91 0.189894
R144 VN.n91 VN.n90 0.189894
R145 VN.n90 VN.n66 0.189894
R146 VN.n85 VN.n66 0.189894
R147 VN.n85 VN.n84 0.189894
R148 VN.n84 VN.n83 0.189894
R149 VN.n83 VN.n68 0.189894
R150 VN.n79 VN.n68 0.189894
R151 VN.n79 VN.n78 0.189894
R152 VN.n78 VN.n77 0.189894
R153 VN.n77 VN.n70 0.189894
R154 VN.n73 VN.n70 0.189894
R155 VN.n15 VN.n12 0.189894
R156 VN.n19 VN.n12 0.189894
R157 VN.n20 VN.n19 0.189894
R158 VN.n21 VN.n20 0.189894
R159 VN.n21 VN.n10 0.189894
R160 VN.n25 VN.n10 0.189894
R161 VN.n26 VN.n25 0.189894
R162 VN.n27 VN.n26 0.189894
R163 VN.n27 VN.n8 0.189894
R164 VN.n32 VN.n8 0.189894
R165 VN.n33 VN.n32 0.189894
R166 VN.n34 VN.n33 0.189894
R167 VN.n34 VN.n6 0.189894
R168 VN.n38 VN.n6 0.189894
R169 VN.n39 VN.n38 0.189894
R170 VN.n40 VN.n39 0.189894
R171 VN.n40 VN.n4 0.189894
R172 VN.n45 VN.n4 0.189894
R173 VN.n46 VN.n45 0.189894
R174 VN.n47 VN.n46 0.189894
R175 VN.n47 VN.n2 0.189894
R176 VN.n51 VN.n2 0.189894
R177 VN.n52 VN.n51 0.189894
R178 VN.n53 VN.n52 0.189894
R179 VN.n53 VN.n0 0.189894
R180 VTAIL.n11 VTAIL.t16 69.6154
R181 VTAIL.n16 VTAIL.t1 69.6152
R182 VTAIL.n17 VTAIL.t9 69.6152
R183 VTAIL.n2 VTAIL.t8 69.6152
R184 VTAIL.n15 VTAIL.n14 66.0237
R185 VTAIL.n13 VTAIL.n12 66.0237
R186 VTAIL.n10 VTAIL.n9 66.0237
R187 VTAIL.n8 VTAIL.n7 66.0237
R188 VTAIL.n19 VTAIL.n18 66.0234
R189 VTAIL.n1 VTAIL.n0 66.0234
R190 VTAIL.n4 VTAIL.n3 66.0234
R191 VTAIL.n6 VTAIL.n5 66.0234
R192 VTAIL.n8 VTAIL.n6 27.6341
R193 VTAIL.n17 VTAIL.n16 23.9014
R194 VTAIL.n10 VTAIL.n8 3.73326
R195 VTAIL.n11 VTAIL.n10 3.73326
R196 VTAIL.n15 VTAIL.n13 3.73326
R197 VTAIL.n16 VTAIL.n15 3.73326
R198 VTAIL.n6 VTAIL.n4 3.73326
R199 VTAIL.n4 VTAIL.n2 3.73326
R200 VTAIL.n19 VTAIL.n17 3.73326
R201 VTAIL.n18 VTAIL.t14 3.59221
R202 VTAIL.n18 VTAIL.t12 3.59221
R203 VTAIL.n0 VTAIL.t17 3.59221
R204 VTAIL.n0 VTAIL.t13 3.59221
R205 VTAIL.n3 VTAIL.t4 3.59221
R206 VTAIL.n3 VTAIL.t2 3.59221
R207 VTAIL.n5 VTAIL.t5 3.59221
R208 VTAIL.n5 VTAIL.t6 3.59221
R209 VTAIL.n14 VTAIL.t19 3.59221
R210 VTAIL.n14 VTAIL.t7 3.59221
R211 VTAIL.n12 VTAIL.t3 3.59221
R212 VTAIL.n12 VTAIL.t0 3.59221
R213 VTAIL.n9 VTAIL.t10 3.59221
R214 VTAIL.n9 VTAIL.t15 3.59221
R215 VTAIL.n7 VTAIL.t11 3.59221
R216 VTAIL.n7 VTAIL.t18 3.59221
R217 VTAIL VTAIL.n1 2.85826
R218 VTAIL.n13 VTAIL.n11 2.33671
R219 VTAIL.n2 VTAIL.n1 2.33671
R220 VTAIL VTAIL.n19 0.8755
R221 VDD2.n1 VDD2.t4 90.0267
R222 VDD2.n4 VDD2.t7 86.2942
R223 VDD2.n3 VDD2.n2 85.4465
R224 VDD2 VDD2.n7 85.4437
R225 VDD2.n6 VDD2.n5 82.7025
R226 VDD2.n1 VDD2.n0 82.7022
R227 VDD2.n4 VDD2.n3 49.2476
R228 VDD2.n6 VDD2.n4 3.73326
R229 VDD2.n7 VDD2.t0 3.59221
R230 VDD2.n7 VDD2.t6 3.59221
R231 VDD2.n5 VDD2.t8 3.59221
R232 VDD2.n5 VDD2.t9 3.59221
R233 VDD2.n2 VDD2.t2 3.59221
R234 VDD2.n2 VDD2.t3 3.59221
R235 VDD2.n0 VDD2.t1 3.59221
R236 VDD2.n0 VDD2.t5 3.59221
R237 VDD2 VDD2.n6 0.991879
R238 VDD2.n3 VDD2.n1 0.878344
R239 VP.n34 VP.n33 161.3
R240 VP.n35 VP.n30 161.3
R241 VP.n37 VP.n36 161.3
R242 VP.n38 VP.n29 161.3
R243 VP.n40 VP.n39 161.3
R244 VP.n41 VP.n28 161.3
R245 VP.n43 VP.n42 161.3
R246 VP.n44 VP.n27 161.3
R247 VP.n46 VP.n45 161.3
R248 VP.n48 VP.n26 161.3
R249 VP.n50 VP.n49 161.3
R250 VP.n51 VP.n25 161.3
R251 VP.n53 VP.n52 161.3
R252 VP.n54 VP.n24 161.3
R253 VP.n56 VP.n55 161.3
R254 VP.n57 VP.n23 161.3
R255 VP.n59 VP.n58 161.3
R256 VP.n60 VP.n22 161.3
R257 VP.n63 VP.n62 161.3
R258 VP.n64 VP.n21 161.3
R259 VP.n66 VP.n65 161.3
R260 VP.n67 VP.n20 161.3
R261 VP.n69 VP.n68 161.3
R262 VP.n70 VP.n19 161.3
R263 VP.n72 VP.n71 161.3
R264 VP.n73 VP.n18 161.3
R265 VP.n130 VP.n0 161.3
R266 VP.n129 VP.n128 161.3
R267 VP.n127 VP.n1 161.3
R268 VP.n126 VP.n125 161.3
R269 VP.n124 VP.n2 161.3
R270 VP.n123 VP.n122 161.3
R271 VP.n121 VP.n3 161.3
R272 VP.n120 VP.n119 161.3
R273 VP.n117 VP.n4 161.3
R274 VP.n116 VP.n115 161.3
R275 VP.n114 VP.n5 161.3
R276 VP.n113 VP.n112 161.3
R277 VP.n111 VP.n6 161.3
R278 VP.n110 VP.n109 161.3
R279 VP.n108 VP.n7 161.3
R280 VP.n107 VP.n106 161.3
R281 VP.n105 VP.n8 161.3
R282 VP.n103 VP.n102 161.3
R283 VP.n101 VP.n9 161.3
R284 VP.n100 VP.n99 161.3
R285 VP.n98 VP.n10 161.3
R286 VP.n97 VP.n96 161.3
R287 VP.n95 VP.n11 161.3
R288 VP.n94 VP.n93 161.3
R289 VP.n92 VP.n12 161.3
R290 VP.n91 VP.n90 161.3
R291 VP.n89 VP.n88 161.3
R292 VP.n87 VP.n14 161.3
R293 VP.n86 VP.n85 161.3
R294 VP.n84 VP.n15 161.3
R295 VP.n83 VP.n82 161.3
R296 VP.n81 VP.n16 161.3
R297 VP.n80 VP.n79 161.3
R298 VP.n78 VP.n17 161.3
R299 VP.n32 VP.t6 86.7958
R300 VP.n32 VP.n31 71.1463
R301 VP.n77 VP.n76 62.1188
R302 VP.n132 VP.n131 62.1188
R303 VP.n75 VP.n74 62.1188
R304 VP.n77 VP.n75 58.7351
R305 VP.n82 VP.n15 56.5193
R306 VP.n125 VP.n124 56.5193
R307 VP.n68 VP.n67 56.5193
R308 VP.n76 VP.t2 54.5267
R309 VP.n13 VP.t8 54.5267
R310 VP.n104 VP.t7 54.5267
R311 VP.n118 VP.t1 54.5267
R312 VP.n131 VP.t9 54.5267
R313 VP.n74 VP.t5 54.5267
R314 VP.n61 VP.t3 54.5267
R315 VP.n47 VP.t0 54.5267
R316 VP.n31 VP.t4 54.5267
R317 VP.n98 VP.n97 48.7492
R318 VP.n111 VP.n110 48.7492
R319 VP.n54 VP.n53 48.7492
R320 VP.n41 VP.n40 48.7492
R321 VP.n97 VP.n11 32.2376
R322 VP.n112 VP.n111 32.2376
R323 VP.n55 VP.n54 32.2376
R324 VP.n40 VP.n29 32.2376
R325 VP.n80 VP.n17 24.4675
R326 VP.n81 VP.n80 24.4675
R327 VP.n82 VP.n81 24.4675
R328 VP.n86 VP.n15 24.4675
R329 VP.n87 VP.n86 24.4675
R330 VP.n88 VP.n87 24.4675
R331 VP.n92 VP.n91 24.4675
R332 VP.n93 VP.n92 24.4675
R333 VP.n93 VP.n11 24.4675
R334 VP.n99 VP.n98 24.4675
R335 VP.n99 VP.n9 24.4675
R336 VP.n103 VP.n9 24.4675
R337 VP.n106 VP.n105 24.4675
R338 VP.n106 VP.n7 24.4675
R339 VP.n110 VP.n7 24.4675
R340 VP.n112 VP.n5 24.4675
R341 VP.n116 VP.n5 24.4675
R342 VP.n117 VP.n116 24.4675
R343 VP.n119 VP.n3 24.4675
R344 VP.n123 VP.n3 24.4675
R345 VP.n124 VP.n123 24.4675
R346 VP.n125 VP.n1 24.4675
R347 VP.n129 VP.n1 24.4675
R348 VP.n130 VP.n129 24.4675
R349 VP.n68 VP.n19 24.4675
R350 VP.n72 VP.n19 24.4675
R351 VP.n73 VP.n72 24.4675
R352 VP.n55 VP.n23 24.4675
R353 VP.n59 VP.n23 24.4675
R354 VP.n60 VP.n59 24.4675
R355 VP.n62 VP.n21 24.4675
R356 VP.n66 VP.n21 24.4675
R357 VP.n67 VP.n66 24.4675
R358 VP.n42 VP.n41 24.4675
R359 VP.n42 VP.n27 24.4675
R360 VP.n46 VP.n27 24.4675
R361 VP.n49 VP.n48 24.4675
R362 VP.n49 VP.n25 24.4675
R363 VP.n53 VP.n25 24.4675
R364 VP.n35 VP.n34 24.4675
R365 VP.n36 VP.n35 24.4675
R366 VP.n36 VP.n29 24.4675
R367 VP.n88 VP.n13 20.5528
R368 VP.n119 VP.n118 20.5528
R369 VP.n62 VP.n61 20.5528
R370 VP.n76 VP.n17 20.0634
R371 VP.n131 VP.n130 20.0634
R372 VP.n74 VP.n73 20.0634
R373 VP.n104 VP.n103 12.234
R374 VP.n105 VP.n104 12.234
R375 VP.n47 VP.n46 12.234
R376 VP.n48 VP.n47 12.234
R377 VP.n91 VP.n13 3.91522
R378 VP.n118 VP.n117 3.91522
R379 VP.n61 VP.n60 3.91522
R380 VP.n34 VP.n31 3.91522
R381 VP.n33 VP.n32 2.69182
R382 VP.n75 VP.n18 0.417535
R383 VP.n78 VP.n77 0.417535
R384 VP.n132 VP.n0 0.417535
R385 VP VP.n132 0.394291
R386 VP.n33 VP.n30 0.189894
R387 VP.n37 VP.n30 0.189894
R388 VP.n38 VP.n37 0.189894
R389 VP.n39 VP.n38 0.189894
R390 VP.n39 VP.n28 0.189894
R391 VP.n43 VP.n28 0.189894
R392 VP.n44 VP.n43 0.189894
R393 VP.n45 VP.n44 0.189894
R394 VP.n45 VP.n26 0.189894
R395 VP.n50 VP.n26 0.189894
R396 VP.n51 VP.n50 0.189894
R397 VP.n52 VP.n51 0.189894
R398 VP.n52 VP.n24 0.189894
R399 VP.n56 VP.n24 0.189894
R400 VP.n57 VP.n56 0.189894
R401 VP.n58 VP.n57 0.189894
R402 VP.n58 VP.n22 0.189894
R403 VP.n63 VP.n22 0.189894
R404 VP.n64 VP.n63 0.189894
R405 VP.n65 VP.n64 0.189894
R406 VP.n65 VP.n20 0.189894
R407 VP.n69 VP.n20 0.189894
R408 VP.n70 VP.n69 0.189894
R409 VP.n71 VP.n70 0.189894
R410 VP.n71 VP.n18 0.189894
R411 VP.n79 VP.n78 0.189894
R412 VP.n79 VP.n16 0.189894
R413 VP.n83 VP.n16 0.189894
R414 VP.n84 VP.n83 0.189894
R415 VP.n85 VP.n84 0.189894
R416 VP.n85 VP.n14 0.189894
R417 VP.n89 VP.n14 0.189894
R418 VP.n90 VP.n89 0.189894
R419 VP.n90 VP.n12 0.189894
R420 VP.n94 VP.n12 0.189894
R421 VP.n95 VP.n94 0.189894
R422 VP.n96 VP.n95 0.189894
R423 VP.n96 VP.n10 0.189894
R424 VP.n100 VP.n10 0.189894
R425 VP.n101 VP.n100 0.189894
R426 VP.n102 VP.n101 0.189894
R427 VP.n102 VP.n8 0.189894
R428 VP.n107 VP.n8 0.189894
R429 VP.n108 VP.n107 0.189894
R430 VP.n109 VP.n108 0.189894
R431 VP.n109 VP.n6 0.189894
R432 VP.n113 VP.n6 0.189894
R433 VP.n114 VP.n113 0.189894
R434 VP.n115 VP.n114 0.189894
R435 VP.n115 VP.n4 0.189894
R436 VP.n120 VP.n4 0.189894
R437 VP.n121 VP.n120 0.189894
R438 VP.n122 VP.n121 0.189894
R439 VP.n122 VP.n2 0.189894
R440 VP.n126 VP.n2 0.189894
R441 VP.n127 VP.n126 0.189894
R442 VP.n128 VP.n127 0.189894
R443 VP.n128 VP.n0 0.189894
R444 VDD1.n1 VDD1.t3 90.027
R445 VDD1.n3 VDD1.t7 90.0267
R446 VDD1.n5 VDD1.n4 85.4465
R447 VDD1.n1 VDD1.n0 82.7025
R448 VDD1.n7 VDD1.n6 82.7023
R449 VDD1.n3 VDD1.n2 82.7022
R450 VDD1.n7 VDD1.n5 51.697
R451 VDD1.n6 VDD1.t6 3.59221
R452 VDD1.n6 VDD1.t4 3.59221
R453 VDD1.n0 VDD1.t5 3.59221
R454 VDD1.n0 VDD1.t9 3.59221
R455 VDD1.n4 VDD1.t8 3.59221
R456 VDD1.n4 VDD1.t0 3.59221
R457 VDD1.n2 VDD1.t1 3.59221
R458 VDD1.n2 VDD1.t2 3.59221
R459 VDD1 VDD1.n7 2.74188
R460 VDD1 VDD1.n1 0.991879
R461 VDD1.n5 VDD1.n3 0.878344
R462 B.n493 B.n492 585
R463 B.n491 B.n172 585
R464 B.n490 B.n489 585
R465 B.n488 B.n173 585
R466 B.n487 B.n486 585
R467 B.n485 B.n174 585
R468 B.n484 B.n483 585
R469 B.n482 B.n175 585
R470 B.n481 B.n480 585
R471 B.n479 B.n176 585
R472 B.n478 B.n477 585
R473 B.n476 B.n177 585
R474 B.n475 B.n474 585
R475 B.n473 B.n178 585
R476 B.n472 B.n471 585
R477 B.n470 B.n179 585
R478 B.n469 B.n468 585
R479 B.n467 B.n180 585
R480 B.n466 B.n465 585
R481 B.n464 B.n181 585
R482 B.n463 B.n462 585
R483 B.n461 B.n182 585
R484 B.n460 B.n459 585
R485 B.n458 B.n183 585
R486 B.n457 B.n456 585
R487 B.n455 B.n184 585
R488 B.n454 B.n453 585
R489 B.n452 B.n185 585
R490 B.n451 B.n450 585
R491 B.n449 B.n186 585
R492 B.n448 B.n447 585
R493 B.n446 B.n187 585
R494 B.n445 B.n444 585
R495 B.n442 B.n188 585
R496 B.n441 B.n440 585
R497 B.n439 B.n191 585
R498 B.n438 B.n437 585
R499 B.n436 B.n192 585
R500 B.n435 B.n434 585
R501 B.n433 B.n193 585
R502 B.n432 B.n431 585
R503 B.n430 B.n194 585
R504 B.n428 B.n427 585
R505 B.n426 B.n197 585
R506 B.n425 B.n424 585
R507 B.n423 B.n198 585
R508 B.n422 B.n421 585
R509 B.n420 B.n199 585
R510 B.n419 B.n418 585
R511 B.n417 B.n200 585
R512 B.n416 B.n415 585
R513 B.n414 B.n201 585
R514 B.n413 B.n412 585
R515 B.n411 B.n202 585
R516 B.n410 B.n409 585
R517 B.n408 B.n203 585
R518 B.n407 B.n406 585
R519 B.n405 B.n204 585
R520 B.n404 B.n403 585
R521 B.n402 B.n205 585
R522 B.n401 B.n400 585
R523 B.n399 B.n206 585
R524 B.n398 B.n397 585
R525 B.n396 B.n207 585
R526 B.n395 B.n394 585
R527 B.n393 B.n208 585
R528 B.n392 B.n391 585
R529 B.n390 B.n209 585
R530 B.n389 B.n388 585
R531 B.n387 B.n210 585
R532 B.n386 B.n385 585
R533 B.n384 B.n211 585
R534 B.n383 B.n382 585
R535 B.n381 B.n212 585
R536 B.n380 B.n379 585
R537 B.n494 B.n171 585
R538 B.n496 B.n495 585
R539 B.n497 B.n170 585
R540 B.n499 B.n498 585
R541 B.n500 B.n169 585
R542 B.n502 B.n501 585
R543 B.n503 B.n168 585
R544 B.n505 B.n504 585
R545 B.n506 B.n167 585
R546 B.n508 B.n507 585
R547 B.n509 B.n166 585
R548 B.n511 B.n510 585
R549 B.n512 B.n165 585
R550 B.n514 B.n513 585
R551 B.n515 B.n164 585
R552 B.n517 B.n516 585
R553 B.n518 B.n163 585
R554 B.n520 B.n519 585
R555 B.n521 B.n162 585
R556 B.n523 B.n522 585
R557 B.n524 B.n161 585
R558 B.n526 B.n525 585
R559 B.n527 B.n160 585
R560 B.n529 B.n528 585
R561 B.n530 B.n159 585
R562 B.n532 B.n531 585
R563 B.n533 B.n158 585
R564 B.n535 B.n534 585
R565 B.n536 B.n157 585
R566 B.n538 B.n537 585
R567 B.n539 B.n156 585
R568 B.n541 B.n540 585
R569 B.n542 B.n155 585
R570 B.n544 B.n543 585
R571 B.n545 B.n154 585
R572 B.n547 B.n546 585
R573 B.n548 B.n153 585
R574 B.n550 B.n549 585
R575 B.n551 B.n152 585
R576 B.n553 B.n552 585
R577 B.n554 B.n151 585
R578 B.n556 B.n555 585
R579 B.n557 B.n150 585
R580 B.n559 B.n558 585
R581 B.n560 B.n149 585
R582 B.n562 B.n561 585
R583 B.n563 B.n148 585
R584 B.n565 B.n564 585
R585 B.n566 B.n147 585
R586 B.n568 B.n567 585
R587 B.n569 B.n146 585
R588 B.n571 B.n570 585
R589 B.n572 B.n145 585
R590 B.n574 B.n573 585
R591 B.n575 B.n144 585
R592 B.n577 B.n576 585
R593 B.n578 B.n143 585
R594 B.n580 B.n579 585
R595 B.n581 B.n142 585
R596 B.n583 B.n582 585
R597 B.n584 B.n141 585
R598 B.n586 B.n585 585
R599 B.n587 B.n140 585
R600 B.n589 B.n588 585
R601 B.n590 B.n139 585
R602 B.n592 B.n591 585
R603 B.n593 B.n138 585
R604 B.n595 B.n594 585
R605 B.n596 B.n137 585
R606 B.n598 B.n597 585
R607 B.n599 B.n136 585
R608 B.n601 B.n600 585
R609 B.n602 B.n135 585
R610 B.n604 B.n603 585
R611 B.n605 B.n134 585
R612 B.n607 B.n606 585
R613 B.n608 B.n133 585
R614 B.n610 B.n609 585
R615 B.n611 B.n132 585
R616 B.n613 B.n612 585
R617 B.n614 B.n131 585
R618 B.n616 B.n615 585
R619 B.n617 B.n130 585
R620 B.n619 B.n618 585
R621 B.n620 B.n129 585
R622 B.n622 B.n621 585
R623 B.n623 B.n128 585
R624 B.n625 B.n624 585
R625 B.n626 B.n127 585
R626 B.n628 B.n627 585
R627 B.n629 B.n126 585
R628 B.n631 B.n630 585
R629 B.n632 B.n125 585
R630 B.n634 B.n633 585
R631 B.n635 B.n124 585
R632 B.n637 B.n636 585
R633 B.n638 B.n123 585
R634 B.n640 B.n639 585
R635 B.n641 B.n122 585
R636 B.n643 B.n642 585
R637 B.n644 B.n121 585
R638 B.n646 B.n645 585
R639 B.n647 B.n120 585
R640 B.n649 B.n648 585
R641 B.n650 B.n119 585
R642 B.n652 B.n651 585
R643 B.n653 B.n118 585
R644 B.n655 B.n654 585
R645 B.n656 B.n117 585
R646 B.n658 B.n657 585
R647 B.n659 B.n116 585
R648 B.n661 B.n660 585
R649 B.n662 B.n115 585
R650 B.n664 B.n663 585
R651 B.n665 B.n114 585
R652 B.n667 B.n666 585
R653 B.n668 B.n113 585
R654 B.n670 B.n669 585
R655 B.n671 B.n112 585
R656 B.n673 B.n672 585
R657 B.n674 B.n111 585
R658 B.n676 B.n675 585
R659 B.n677 B.n110 585
R660 B.n679 B.n678 585
R661 B.n680 B.n109 585
R662 B.n682 B.n681 585
R663 B.n683 B.n108 585
R664 B.n685 B.n684 585
R665 B.n686 B.n107 585
R666 B.n688 B.n687 585
R667 B.n689 B.n106 585
R668 B.n691 B.n690 585
R669 B.n692 B.n105 585
R670 B.n694 B.n693 585
R671 B.n695 B.n104 585
R672 B.n697 B.n696 585
R673 B.n698 B.n103 585
R674 B.n700 B.n699 585
R675 B.n701 B.n102 585
R676 B.n703 B.n702 585
R677 B.n704 B.n101 585
R678 B.n706 B.n705 585
R679 B.n707 B.n100 585
R680 B.n709 B.n708 585
R681 B.n710 B.n99 585
R682 B.n712 B.n711 585
R683 B.n713 B.n98 585
R684 B.n715 B.n714 585
R685 B.n716 B.n97 585
R686 B.n718 B.n717 585
R687 B.n719 B.n96 585
R688 B.n721 B.n720 585
R689 B.n722 B.n95 585
R690 B.n724 B.n723 585
R691 B.n725 B.n94 585
R692 B.n727 B.n726 585
R693 B.n728 B.n93 585
R694 B.n730 B.n729 585
R695 B.n731 B.n92 585
R696 B.n733 B.n732 585
R697 B.n734 B.n91 585
R698 B.n736 B.n735 585
R699 B.n737 B.n90 585
R700 B.n739 B.n738 585
R701 B.n740 B.n89 585
R702 B.n742 B.n741 585
R703 B.n743 B.n88 585
R704 B.n745 B.n744 585
R705 B.n746 B.n87 585
R706 B.n748 B.n747 585
R707 B.n861 B.n44 585
R708 B.n860 B.n859 585
R709 B.n858 B.n45 585
R710 B.n857 B.n856 585
R711 B.n855 B.n46 585
R712 B.n854 B.n853 585
R713 B.n852 B.n47 585
R714 B.n851 B.n850 585
R715 B.n849 B.n48 585
R716 B.n848 B.n847 585
R717 B.n846 B.n49 585
R718 B.n845 B.n844 585
R719 B.n843 B.n50 585
R720 B.n842 B.n841 585
R721 B.n840 B.n51 585
R722 B.n839 B.n838 585
R723 B.n837 B.n52 585
R724 B.n836 B.n835 585
R725 B.n834 B.n53 585
R726 B.n833 B.n832 585
R727 B.n831 B.n54 585
R728 B.n830 B.n829 585
R729 B.n828 B.n55 585
R730 B.n827 B.n826 585
R731 B.n825 B.n56 585
R732 B.n824 B.n823 585
R733 B.n822 B.n57 585
R734 B.n821 B.n820 585
R735 B.n819 B.n58 585
R736 B.n818 B.n817 585
R737 B.n816 B.n59 585
R738 B.n815 B.n814 585
R739 B.n813 B.n60 585
R740 B.n812 B.n811 585
R741 B.n810 B.n61 585
R742 B.n809 B.n808 585
R743 B.n807 B.n65 585
R744 B.n806 B.n805 585
R745 B.n804 B.n66 585
R746 B.n803 B.n802 585
R747 B.n801 B.n67 585
R748 B.n800 B.n799 585
R749 B.n797 B.n68 585
R750 B.n796 B.n795 585
R751 B.n794 B.n71 585
R752 B.n793 B.n792 585
R753 B.n791 B.n72 585
R754 B.n790 B.n789 585
R755 B.n788 B.n73 585
R756 B.n787 B.n786 585
R757 B.n785 B.n74 585
R758 B.n784 B.n783 585
R759 B.n782 B.n75 585
R760 B.n781 B.n780 585
R761 B.n779 B.n76 585
R762 B.n778 B.n777 585
R763 B.n776 B.n77 585
R764 B.n775 B.n774 585
R765 B.n773 B.n78 585
R766 B.n772 B.n771 585
R767 B.n770 B.n79 585
R768 B.n769 B.n768 585
R769 B.n767 B.n80 585
R770 B.n766 B.n765 585
R771 B.n764 B.n81 585
R772 B.n763 B.n762 585
R773 B.n761 B.n82 585
R774 B.n760 B.n759 585
R775 B.n758 B.n83 585
R776 B.n757 B.n756 585
R777 B.n755 B.n84 585
R778 B.n754 B.n753 585
R779 B.n752 B.n85 585
R780 B.n751 B.n750 585
R781 B.n749 B.n86 585
R782 B.n863 B.n862 585
R783 B.n864 B.n43 585
R784 B.n866 B.n865 585
R785 B.n867 B.n42 585
R786 B.n869 B.n868 585
R787 B.n870 B.n41 585
R788 B.n872 B.n871 585
R789 B.n873 B.n40 585
R790 B.n875 B.n874 585
R791 B.n876 B.n39 585
R792 B.n878 B.n877 585
R793 B.n879 B.n38 585
R794 B.n881 B.n880 585
R795 B.n882 B.n37 585
R796 B.n884 B.n883 585
R797 B.n885 B.n36 585
R798 B.n887 B.n886 585
R799 B.n888 B.n35 585
R800 B.n890 B.n889 585
R801 B.n891 B.n34 585
R802 B.n893 B.n892 585
R803 B.n894 B.n33 585
R804 B.n896 B.n895 585
R805 B.n897 B.n32 585
R806 B.n899 B.n898 585
R807 B.n900 B.n31 585
R808 B.n902 B.n901 585
R809 B.n903 B.n30 585
R810 B.n905 B.n904 585
R811 B.n906 B.n29 585
R812 B.n908 B.n907 585
R813 B.n909 B.n28 585
R814 B.n911 B.n910 585
R815 B.n912 B.n27 585
R816 B.n914 B.n913 585
R817 B.n915 B.n26 585
R818 B.n917 B.n916 585
R819 B.n918 B.n25 585
R820 B.n920 B.n919 585
R821 B.n921 B.n24 585
R822 B.n923 B.n922 585
R823 B.n924 B.n23 585
R824 B.n926 B.n925 585
R825 B.n927 B.n22 585
R826 B.n929 B.n928 585
R827 B.n930 B.n21 585
R828 B.n932 B.n931 585
R829 B.n933 B.n20 585
R830 B.n935 B.n934 585
R831 B.n936 B.n19 585
R832 B.n938 B.n937 585
R833 B.n939 B.n18 585
R834 B.n941 B.n940 585
R835 B.n942 B.n17 585
R836 B.n944 B.n943 585
R837 B.n945 B.n16 585
R838 B.n947 B.n946 585
R839 B.n948 B.n15 585
R840 B.n950 B.n949 585
R841 B.n951 B.n14 585
R842 B.n953 B.n952 585
R843 B.n954 B.n13 585
R844 B.n956 B.n955 585
R845 B.n957 B.n12 585
R846 B.n959 B.n958 585
R847 B.n960 B.n11 585
R848 B.n962 B.n961 585
R849 B.n963 B.n10 585
R850 B.n965 B.n964 585
R851 B.n966 B.n9 585
R852 B.n968 B.n967 585
R853 B.n969 B.n8 585
R854 B.n971 B.n970 585
R855 B.n972 B.n7 585
R856 B.n974 B.n973 585
R857 B.n975 B.n6 585
R858 B.n977 B.n976 585
R859 B.n978 B.n5 585
R860 B.n980 B.n979 585
R861 B.n981 B.n4 585
R862 B.n983 B.n982 585
R863 B.n984 B.n3 585
R864 B.n986 B.n985 585
R865 B.n987 B.n0 585
R866 B.n2 B.n1 585
R867 B.n255 B.n254 585
R868 B.n257 B.n256 585
R869 B.n258 B.n253 585
R870 B.n260 B.n259 585
R871 B.n261 B.n252 585
R872 B.n263 B.n262 585
R873 B.n264 B.n251 585
R874 B.n266 B.n265 585
R875 B.n267 B.n250 585
R876 B.n269 B.n268 585
R877 B.n270 B.n249 585
R878 B.n272 B.n271 585
R879 B.n273 B.n248 585
R880 B.n275 B.n274 585
R881 B.n276 B.n247 585
R882 B.n278 B.n277 585
R883 B.n279 B.n246 585
R884 B.n281 B.n280 585
R885 B.n282 B.n245 585
R886 B.n284 B.n283 585
R887 B.n285 B.n244 585
R888 B.n287 B.n286 585
R889 B.n288 B.n243 585
R890 B.n290 B.n289 585
R891 B.n291 B.n242 585
R892 B.n293 B.n292 585
R893 B.n294 B.n241 585
R894 B.n296 B.n295 585
R895 B.n297 B.n240 585
R896 B.n299 B.n298 585
R897 B.n300 B.n239 585
R898 B.n302 B.n301 585
R899 B.n303 B.n238 585
R900 B.n305 B.n304 585
R901 B.n306 B.n237 585
R902 B.n308 B.n307 585
R903 B.n309 B.n236 585
R904 B.n311 B.n310 585
R905 B.n312 B.n235 585
R906 B.n314 B.n313 585
R907 B.n315 B.n234 585
R908 B.n317 B.n316 585
R909 B.n318 B.n233 585
R910 B.n320 B.n319 585
R911 B.n321 B.n232 585
R912 B.n323 B.n322 585
R913 B.n324 B.n231 585
R914 B.n326 B.n325 585
R915 B.n327 B.n230 585
R916 B.n329 B.n328 585
R917 B.n330 B.n229 585
R918 B.n332 B.n331 585
R919 B.n333 B.n228 585
R920 B.n335 B.n334 585
R921 B.n336 B.n227 585
R922 B.n338 B.n337 585
R923 B.n339 B.n226 585
R924 B.n341 B.n340 585
R925 B.n342 B.n225 585
R926 B.n344 B.n343 585
R927 B.n345 B.n224 585
R928 B.n347 B.n346 585
R929 B.n348 B.n223 585
R930 B.n350 B.n349 585
R931 B.n351 B.n222 585
R932 B.n353 B.n352 585
R933 B.n354 B.n221 585
R934 B.n356 B.n355 585
R935 B.n357 B.n220 585
R936 B.n359 B.n358 585
R937 B.n360 B.n219 585
R938 B.n362 B.n361 585
R939 B.n363 B.n218 585
R940 B.n365 B.n364 585
R941 B.n366 B.n217 585
R942 B.n368 B.n367 585
R943 B.n369 B.n216 585
R944 B.n371 B.n370 585
R945 B.n372 B.n215 585
R946 B.n374 B.n373 585
R947 B.n375 B.n214 585
R948 B.n377 B.n376 585
R949 B.n378 B.n213 585
R950 B.n379 B.n378 540.549
R951 B.n494 B.n493 540.549
R952 B.n747 B.n86 540.549
R953 B.n862 B.n861 540.549
R954 B.n195 B.t0 264.017
R955 B.n189 B.t9 264.017
R956 B.n69 B.t3 264.017
R957 B.n62 B.t6 264.017
R958 B.n989 B.n988 256.663
R959 B.n988 B.n987 235.042
R960 B.n988 B.n2 235.042
R961 B.n189 B.t10 196.123
R962 B.n69 B.t5 196.123
R963 B.n195 B.t1 196.113
R964 B.n62 B.t8 196.113
R965 B.n379 B.n212 163.367
R966 B.n383 B.n212 163.367
R967 B.n384 B.n383 163.367
R968 B.n385 B.n384 163.367
R969 B.n385 B.n210 163.367
R970 B.n389 B.n210 163.367
R971 B.n390 B.n389 163.367
R972 B.n391 B.n390 163.367
R973 B.n391 B.n208 163.367
R974 B.n395 B.n208 163.367
R975 B.n396 B.n395 163.367
R976 B.n397 B.n396 163.367
R977 B.n397 B.n206 163.367
R978 B.n401 B.n206 163.367
R979 B.n402 B.n401 163.367
R980 B.n403 B.n402 163.367
R981 B.n403 B.n204 163.367
R982 B.n407 B.n204 163.367
R983 B.n408 B.n407 163.367
R984 B.n409 B.n408 163.367
R985 B.n409 B.n202 163.367
R986 B.n413 B.n202 163.367
R987 B.n414 B.n413 163.367
R988 B.n415 B.n414 163.367
R989 B.n415 B.n200 163.367
R990 B.n419 B.n200 163.367
R991 B.n420 B.n419 163.367
R992 B.n421 B.n420 163.367
R993 B.n421 B.n198 163.367
R994 B.n425 B.n198 163.367
R995 B.n426 B.n425 163.367
R996 B.n427 B.n426 163.367
R997 B.n427 B.n194 163.367
R998 B.n432 B.n194 163.367
R999 B.n433 B.n432 163.367
R1000 B.n434 B.n433 163.367
R1001 B.n434 B.n192 163.367
R1002 B.n438 B.n192 163.367
R1003 B.n439 B.n438 163.367
R1004 B.n440 B.n439 163.367
R1005 B.n440 B.n188 163.367
R1006 B.n445 B.n188 163.367
R1007 B.n446 B.n445 163.367
R1008 B.n447 B.n446 163.367
R1009 B.n447 B.n186 163.367
R1010 B.n451 B.n186 163.367
R1011 B.n452 B.n451 163.367
R1012 B.n453 B.n452 163.367
R1013 B.n453 B.n184 163.367
R1014 B.n457 B.n184 163.367
R1015 B.n458 B.n457 163.367
R1016 B.n459 B.n458 163.367
R1017 B.n459 B.n182 163.367
R1018 B.n463 B.n182 163.367
R1019 B.n464 B.n463 163.367
R1020 B.n465 B.n464 163.367
R1021 B.n465 B.n180 163.367
R1022 B.n469 B.n180 163.367
R1023 B.n470 B.n469 163.367
R1024 B.n471 B.n470 163.367
R1025 B.n471 B.n178 163.367
R1026 B.n475 B.n178 163.367
R1027 B.n476 B.n475 163.367
R1028 B.n477 B.n476 163.367
R1029 B.n477 B.n176 163.367
R1030 B.n481 B.n176 163.367
R1031 B.n482 B.n481 163.367
R1032 B.n483 B.n482 163.367
R1033 B.n483 B.n174 163.367
R1034 B.n487 B.n174 163.367
R1035 B.n488 B.n487 163.367
R1036 B.n489 B.n488 163.367
R1037 B.n489 B.n172 163.367
R1038 B.n493 B.n172 163.367
R1039 B.n747 B.n746 163.367
R1040 B.n746 B.n745 163.367
R1041 B.n745 B.n88 163.367
R1042 B.n741 B.n88 163.367
R1043 B.n741 B.n740 163.367
R1044 B.n740 B.n739 163.367
R1045 B.n739 B.n90 163.367
R1046 B.n735 B.n90 163.367
R1047 B.n735 B.n734 163.367
R1048 B.n734 B.n733 163.367
R1049 B.n733 B.n92 163.367
R1050 B.n729 B.n92 163.367
R1051 B.n729 B.n728 163.367
R1052 B.n728 B.n727 163.367
R1053 B.n727 B.n94 163.367
R1054 B.n723 B.n94 163.367
R1055 B.n723 B.n722 163.367
R1056 B.n722 B.n721 163.367
R1057 B.n721 B.n96 163.367
R1058 B.n717 B.n96 163.367
R1059 B.n717 B.n716 163.367
R1060 B.n716 B.n715 163.367
R1061 B.n715 B.n98 163.367
R1062 B.n711 B.n98 163.367
R1063 B.n711 B.n710 163.367
R1064 B.n710 B.n709 163.367
R1065 B.n709 B.n100 163.367
R1066 B.n705 B.n100 163.367
R1067 B.n705 B.n704 163.367
R1068 B.n704 B.n703 163.367
R1069 B.n703 B.n102 163.367
R1070 B.n699 B.n102 163.367
R1071 B.n699 B.n698 163.367
R1072 B.n698 B.n697 163.367
R1073 B.n697 B.n104 163.367
R1074 B.n693 B.n104 163.367
R1075 B.n693 B.n692 163.367
R1076 B.n692 B.n691 163.367
R1077 B.n691 B.n106 163.367
R1078 B.n687 B.n106 163.367
R1079 B.n687 B.n686 163.367
R1080 B.n686 B.n685 163.367
R1081 B.n685 B.n108 163.367
R1082 B.n681 B.n108 163.367
R1083 B.n681 B.n680 163.367
R1084 B.n680 B.n679 163.367
R1085 B.n679 B.n110 163.367
R1086 B.n675 B.n110 163.367
R1087 B.n675 B.n674 163.367
R1088 B.n674 B.n673 163.367
R1089 B.n673 B.n112 163.367
R1090 B.n669 B.n112 163.367
R1091 B.n669 B.n668 163.367
R1092 B.n668 B.n667 163.367
R1093 B.n667 B.n114 163.367
R1094 B.n663 B.n114 163.367
R1095 B.n663 B.n662 163.367
R1096 B.n662 B.n661 163.367
R1097 B.n661 B.n116 163.367
R1098 B.n657 B.n116 163.367
R1099 B.n657 B.n656 163.367
R1100 B.n656 B.n655 163.367
R1101 B.n655 B.n118 163.367
R1102 B.n651 B.n118 163.367
R1103 B.n651 B.n650 163.367
R1104 B.n650 B.n649 163.367
R1105 B.n649 B.n120 163.367
R1106 B.n645 B.n120 163.367
R1107 B.n645 B.n644 163.367
R1108 B.n644 B.n643 163.367
R1109 B.n643 B.n122 163.367
R1110 B.n639 B.n122 163.367
R1111 B.n639 B.n638 163.367
R1112 B.n638 B.n637 163.367
R1113 B.n637 B.n124 163.367
R1114 B.n633 B.n124 163.367
R1115 B.n633 B.n632 163.367
R1116 B.n632 B.n631 163.367
R1117 B.n631 B.n126 163.367
R1118 B.n627 B.n126 163.367
R1119 B.n627 B.n626 163.367
R1120 B.n626 B.n625 163.367
R1121 B.n625 B.n128 163.367
R1122 B.n621 B.n128 163.367
R1123 B.n621 B.n620 163.367
R1124 B.n620 B.n619 163.367
R1125 B.n619 B.n130 163.367
R1126 B.n615 B.n130 163.367
R1127 B.n615 B.n614 163.367
R1128 B.n614 B.n613 163.367
R1129 B.n613 B.n132 163.367
R1130 B.n609 B.n132 163.367
R1131 B.n609 B.n608 163.367
R1132 B.n608 B.n607 163.367
R1133 B.n607 B.n134 163.367
R1134 B.n603 B.n134 163.367
R1135 B.n603 B.n602 163.367
R1136 B.n602 B.n601 163.367
R1137 B.n601 B.n136 163.367
R1138 B.n597 B.n136 163.367
R1139 B.n597 B.n596 163.367
R1140 B.n596 B.n595 163.367
R1141 B.n595 B.n138 163.367
R1142 B.n591 B.n138 163.367
R1143 B.n591 B.n590 163.367
R1144 B.n590 B.n589 163.367
R1145 B.n589 B.n140 163.367
R1146 B.n585 B.n140 163.367
R1147 B.n585 B.n584 163.367
R1148 B.n584 B.n583 163.367
R1149 B.n583 B.n142 163.367
R1150 B.n579 B.n142 163.367
R1151 B.n579 B.n578 163.367
R1152 B.n578 B.n577 163.367
R1153 B.n577 B.n144 163.367
R1154 B.n573 B.n144 163.367
R1155 B.n573 B.n572 163.367
R1156 B.n572 B.n571 163.367
R1157 B.n571 B.n146 163.367
R1158 B.n567 B.n146 163.367
R1159 B.n567 B.n566 163.367
R1160 B.n566 B.n565 163.367
R1161 B.n565 B.n148 163.367
R1162 B.n561 B.n148 163.367
R1163 B.n561 B.n560 163.367
R1164 B.n560 B.n559 163.367
R1165 B.n559 B.n150 163.367
R1166 B.n555 B.n150 163.367
R1167 B.n555 B.n554 163.367
R1168 B.n554 B.n553 163.367
R1169 B.n553 B.n152 163.367
R1170 B.n549 B.n152 163.367
R1171 B.n549 B.n548 163.367
R1172 B.n548 B.n547 163.367
R1173 B.n547 B.n154 163.367
R1174 B.n543 B.n154 163.367
R1175 B.n543 B.n542 163.367
R1176 B.n542 B.n541 163.367
R1177 B.n541 B.n156 163.367
R1178 B.n537 B.n156 163.367
R1179 B.n537 B.n536 163.367
R1180 B.n536 B.n535 163.367
R1181 B.n535 B.n158 163.367
R1182 B.n531 B.n158 163.367
R1183 B.n531 B.n530 163.367
R1184 B.n530 B.n529 163.367
R1185 B.n529 B.n160 163.367
R1186 B.n525 B.n160 163.367
R1187 B.n525 B.n524 163.367
R1188 B.n524 B.n523 163.367
R1189 B.n523 B.n162 163.367
R1190 B.n519 B.n162 163.367
R1191 B.n519 B.n518 163.367
R1192 B.n518 B.n517 163.367
R1193 B.n517 B.n164 163.367
R1194 B.n513 B.n164 163.367
R1195 B.n513 B.n512 163.367
R1196 B.n512 B.n511 163.367
R1197 B.n511 B.n166 163.367
R1198 B.n507 B.n166 163.367
R1199 B.n507 B.n506 163.367
R1200 B.n506 B.n505 163.367
R1201 B.n505 B.n168 163.367
R1202 B.n501 B.n168 163.367
R1203 B.n501 B.n500 163.367
R1204 B.n500 B.n499 163.367
R1205 B.n499 B.n170 163.367
R1206 B.n495 B.n170 163.367
R1207 B.n495 B.n494 163.367
R1208 B.n861 B.n860 163.367
R1209 B.n860 B.n45 163.367
R1210 B.n856 B.n45 163.367
R1211 B.n856 B.n855 163.367
R1212 B.n855 B.n854 163.367
R1213 B.n854 B.n47 163.367
R1214 B.n850 B.n47 163.367
R1215 B.n850 B.n849 163.367
R1216 B.n849 B.n848 163.367
R1217 B.n848 B.n49 163.367
R1218 B.n844 B.n49 163.367
R1219 B.n844 B.n843 163.367
R1220 B.n843 B.n842 163.367
R1221 B.n842 B.n51 163.367
R1222 B.n838 B.n51 163.367
R1223 B.n838 B.n837 163.367
R1224 B.n837 B.n836 163.367
R1225 B.n836 B.n53 163.367
R1226 B.n832 B.n53 163.367
R1227 B.n832 B.n831 163.367
R1228 B.n831 B.n830 163.367
R1229 B.n830 B.n55 163.367
R1230 B.n826 B.n55 163.367
R1231 B.n826 B.n825 163.367
R1232 B.n825 B.n824 163.367
R1233 B.n824 B.n57 163.367
R1234 B.n820 B.n57 163.367
R1235 B.n820 B.n819 163.367
R1236 B.n819 B.n818 163.367
R1237 B.n818 B.n59 163.367
R1238 B.n814 B.n59 163.367
R1239 B.n814 B.n813 163.367
R1240 B.n813 B.n812 163.367
R1241 B.n812 B.n61 163.367
R1242 B.n808 B.n61 163.367
R1243 B.n808 B.n807 163.367
R1244 B.n807 B.n806 163.367
R1245 B.n806 B.n66 163.367
R1246 B.n802 B.n66 163.367
R1247 B.n802 B.n801 163.367
R1248 B.n801 B.n800 163.367
R1249 B.n800 B.n68 163.367
R1250 B.n795 B.n68 163.367
R1251 B.n795 B.n794 163.367
R1252 B.n794 B.n793 163.367
R1253 B.n793 B.n72 163.367
R1254 B.n789 B.n72 163.367
R1255 B.n789 B.n788 163.367
R1256 B.n788 B.n787 163.367
R1257 B.n787 B.n74 163.367
R1258 B.n783 B.n74 163.367
R1259 B.n783 B.n782 163.367
R1260 B.n782 B.n781 163.367
R1261 B.n781 B.n76 163.367
R1262 B.n777 B.n76 163.367
R1263 B.n777 B.n776 163.367
R1264 B.n776 B.n775 163.367
R1265 B.n775 B.n78 163.367
R1266 B.n771 B.n78 163.367
R1267 B.n771 B.n770 163.367
R1268 B.n770 B.n769 163.367
R1269 B.n769 B.n80 163.367
R1270 B.n765 B.n80 163.367
R1271 B.n765 B.n764 163.367
R1272 B.n764 B.n763 163.367
R1273 B.n763 B.n82 163.367
R1274 B.n759 B.n82 163.367
R1275 B.n759 B.n758 163.367
R1276 B.n758 B.n757 163.367
R1277 B.n757 B.n84 163.367
R1278 B.n753 B.n84 163.367
R1279 B.n753 B.n752 163.367
R1280 B.n752 B.n751 163.367
R1281 B.n751 B.n86 163.367
R1282 B.n862 B.n43 163.367
R1283 B.n866 B.n43 163.367
R1284 B.n867 B.n866 163.367
R1285 B.n868 B.n867 163.367
R1286 B.n868 B.n41 163.367
R1287 B.n872 B.n41 163.367
R1288 B.n873 B.n872 163.367
R1289 B.n874 B.n873 163.367
R1290 B.n874 B.n39 163.367
R1291 B.n878 B.n39 163.367
R1292 B.n879 B.n878 163.367
R1293 B.n880 B.n879 163.367
R1294 B.n880 B.n37 163.367
R1295 B.n884 B.n37 163.367
R1296 B.n885 B.n884 163.367
R1297 B.n886 B.n885 163.367
R1298 B.n886 B.n35 163.367
R1299 B.n890 B.n35 163.367
R1300 B.n891 B.n890 163.367
R1301 B.n892 B.n891 163.367
R1302 B.n892 B.n33 163.367
R1303 B.n896 B.n33 163.367
R1304 B.n897 B.n896 163.367
R1305 B.n898 B.n897 163.367
R1306 B.n898 B.n31 163.367
R1307 B.n902 B.n31 163.367
R1308 B.n903 B.n902 163.367
R1309 B.n904 B.n903 163.367
R1310 B.n904 B.n29 163.367
R1311 B.n908 B.n29 163.367
R1312 B.n909 B.n908 163.367
R1313 B.n910 B.n909 163.367
R1314 B.n910 B.n27 163.367
R1315 B.n914 B.n27 163.367
R1316 B.n915 B.n914 163.367
R1317 B.n916 B.n915 163.367
R1318 B.n916 B.n25 163.367
R1319 B.n920 B.n25 163.367
R1320 B.n921 B.n920 163.367
R1321 B.n922 B.n921 163.367
R1322 B.n922 B.n23 163.367
R1323 B.n926 B.n23 163.367
R1324 B.n927 B.n926 163.367
R1325 B.n928 B.n927 163.367
R1326 B.n928 B.n21 163.367
R1327 B.n932 B.n21 163.367
R1328 B.n933 B.n932 163.367
R1329 B.n934 B.n933 163.367
R1330 B.n934 B.n19 163.367
R1331 B.n938 B.n19 163.367
R1332 B.n939 B.n938 163.367
R1333 B.n940 B.n939 163.367
R1334 B.n940 B.n17 163.367
R1335 B.n944 B.n17 163.367
R1336 B.n945 B.n944 163.367
R1337 B.n946 B.n945 163.367
R1338 B.n946 B.n15 163.367
R1339 B.n950 B.n15 163.367
R1340 B.n951 B.n950 163.367
R1341 B.n952 B.n951 163.367
R1342 B.n952 B.n13 163.367
R1343 B.n956 B.n13 163.367
R1344 B.n957 B.n956 163.367
R1345 B.n958 B.n957 163.367
R1346 B.n958 B.n11 163.367
R1347 B.n962 B.n11 163.367
R1348 B.n963 B.n962 163.367
R1349 B.n964 B.n963 163.367
R1350 B.n964 B.n9 163.367
R1351 B.n968 B.n9 163.367
R1352 B.n969 B.n968 163.367
R1353 B.n970 B.n969 163.367
R1354 B.n970 B.n7 163.367
R1355 B.n974 B.n7 163.367
R1356 B.n975 B.n974 163.367
R1357 B.n976 B.n975 163.367
R1358 B.n976 B.n5 163.367
R1359 B.n980 B.n5 163.367
R1360 B.n981 B.n980 163.367
R1361 B.n982 B.n981 163.367
R1362 B.n982 B.n3 163.367
R1363 B.n986 B.n3 163.367
R1364 B.n987 B.n986 163.367
R1365 B.n254 B.n2 163.367
R1366 B.n257 B.n254 163.367
R1367 B.n258 B.n257 163.367
R1368 B.n259 B.n258 163.367
R1369 B.n259 B.n252 163.367
R1370 B.n263 B.n252 163.367
R1371 B.n264 B.n263 163.367
R1372 B.n265 B.n264 163.367
R1373 B.n265 B.n250 163.367
R1374 B.n269 B.n250 163.367
R1375 B.n270 B.n269 163.367
R1376 B.n271 B.n270 163.367
R1377 B.n271 B.n248 163.367
R1378 B.n275 B.n248 163.367
R1379 B.n276 B.n275 163.367
R1380 B.n277 B.n276 163.367
R1381 B.n277 B.n246 163.367
R1382 B.n281 B.n246 163.367
R1383 B.n282 B.n281 163.367
R1384 B.n283 B.n282 163.367
R1385 B.n283 B.n244 163.367
R1386 B.n287 B.n244 163.367
R1387 B.n288 B.n287 163.367
R1388 B.n289 B.n288 163.367
R1389 B.n289 B.n242 163.367
R1390 B.n293 B.n242 163.367
R1391 B.n294 B.n293 163.367
R1392 B.n295 B.n294 163.367
R1393 B.n295 B.n240 163.367
R1394 B.n299 B.n240 163.367
R1395 B.n300 B.n299 163.367
R1396 B.n301 B.n300 163.367
R1397 B.n301 B.n238 163.367
R1398 B.n305 B.n238 163.367
R1399 B.n306 B.n305 163.367
R1400 B.n307 B.n306 163.367
R1401 B.n307 B.n236 163.367
R1402 B.n311 B.n236 163.367
R1403 B.n312 B.n311 163.367
R1404 B.n313 B.n312 163.367
R1405 B.n313 B.n234 163.367
R1406 B.n317 B.n234 163.367
R1407 B.n318 B.n317 163.367
R1408 B.n319 B.n318 163.367
R1409 B.n319 B.n232 163.367
R1410 B.n323 B.n232 163.367
R1411 B.n324 B.n323 163.367
R1412 B.n325 B.n324 163.367
R1413 B.n325 B.n230 163.367
R1414 B.n329 B.n230 163.367
R1415 B.n330 B.n329 163.367
R1416 B.n331 B.n330 163.367
R1417 B.n331 B.n228 163.367
R1418 B.n335 B.n228 163.367
R1419 B.n336 B.n335 163.367
R1420 B.n337 B.n336 163.367
R1421 B.n337 B.n226 163.367
R1422 B.n341 B.n226 163.367
R1423 B.n342 B.n341 163.367
R1424 B.n343 B.n342 163.367
R1425 B.n343 B.n224 163.367
R1426 B.n347 B.n224 163.367
R1427 B.n348 B.n347 163.367
R1428 B.n349 B.n348 163.367
R1429 B.n349 B.n222 163.367
R1430 B.n353 B.n222 163.367
R1431 B.n354 B.n353 163.367
R1432 B.n355 B.n354 163.367
R1433 B.n355 B.n220 163.367
R1434 B.n359 B.n220 163.367
R1435 B.n360 B.n359 163.367
R1436 B.n361 B.n360 163.367
R1437 B.n361 B.n218 163.367
R1438 B.n365 B.n218 163.367
R1439 B.n366 B.n365 163.367
R1440 B.n367 B.n366 163.367
R1441 B.n367 B.n216 163.367
R1442 B.n371 B.n216 163.367
R1443 B.n372 B.n371 163.367
R1444 B.n373 B.n372 163.367
R1445 B.n373 B.n214 163.367
R1446 B.n377 B.n214 163.367
R1447 B.n378 B.n377 163.367
R1448 B.n190 B.t11 112.147
R1449 B.n70 B.t4 112.147
R1450 B.n196 B.t2 112.136
R1451 B.n63 B.t7 112.136
R1452 B.n196 B.n195 83.9763
R1453 B.n190 B.n189 83.9763
R1454 B.n70 B.n69 83.9763
R1455 B.n63 B.n62 83.9763
R1456 B.n429 B.n196 59.5399
R1457 B.n443 B.n190 59.5399
R1458 B.n798 B.n70 59.5399
R1459 B.n64 B.n63 59.5399
R1460 B.n863 B.n44 35.1225
R1461 B.n749 B.n748 35.1225
R1462 B.n492 B.n171 35.1225
R1463 B.n380 B.n213 35.1225
R1464 B B.n989 18.0485
R1465 B.n864 B.n863 10.6151
R1466 B.n865 B.n864 10.6151
R1467 B.n865 B.n42 10.6151
R1468 B.n869 B.n42 10.6151
R1469 B.n870 B.n869 10.6151
R1470 B.n871 B.n870 10.6151
R1471 B.n871 B.n40 10.6151
R1472 B.n875 B.n40 10.6151
R1473 B.n876 B.n875 10.6151
R1474 B.n877 B.n876 10.6151
R1475 B.n877 B.n38 10.6151
R1476 B.n881 B.n38 10.6151
R1477 B.n882 B.n881 10.6151
R1478 B.n883 B.n882 10.6151
R1479 B.n883 B.n36 10.6151
R1480 B.n887 B.n36 10.6151
R1481 B.n888 B.n887 10.6151
R1482 B.n889 B.n888 10.6151
R1483 B.n889 B.n34 10.6151
R1484 B.n893 B.n34 10.6151
R1485 B.n894 B.n893 10.6151
R1486 B.n895 B.n894 10.6151
R1487 B.n895 B.n32 10.6151
R1488 B.n899 B.n32 10.6151
R1489 B.n900 B.n899 10.6151
R1490 B.n901 B.n900 10.6151
R1491 B.n901 B.n30 10.6151
R1492 B.n905 B.n30 10.6151
R1493 B.n906 B.n905 10.6151
R1494 B.n907 B.n906 10.6151
R1495 B.n907 B.n28 10.6151
R1496 B.n911 B.n28 10.6151
R1497 B.n912 B.n911 10.6151
R1498 B.n913 B.n912 10.6151
R1499 B.n913 B.n26 10.6151
R1500 B.n917 B.n26 10.6151
R1501 B.n918 B.n917 10.6151
R1502 B.n919 B.n918 10.6151
R1503 B.n919 B.n24 10.6151
R1504 B.n923 B.n24 10.6151
R1505 B.n924 B.n923 10.6151
R1506 B.n925 B.n924 10.6151
R1507 B.n925 B.n22 10.6151
R1508 B.n929 B.n22 10.6151
R1509 B.n930 B.n929 10.6151
R1510 B.n931 B.n930 10.6151
R1511 B.n931 B.n20 10.6151
R1512 B.n935 B.n20 10.6151
R1513 B.n936 B.n935 10.6151
R1514 B.n937 B.n936 10.6151
R1515 B.n937 B.n18 10.6151
R1516 B.n941 B.n18 10.6151
R1517 B.n942 B.n941 10.6151
R1518 B.n943 B.n942 10.6151
R1519 B.n943 B.n16 10.6151
R1520 B.n947 B.n16 10.6151
R1521 B.n948 B.n947 10.6151
R1522 B.n949 B.n948 10.6151
R1523 B.n949 B.n14 10.6151
R1524 B.n953 B.n14 10.6151
R1525 B.n954 B.n953 10.6151
R1526 B.n955 B.n954 10.6151
R1527 B.n955 B.n12 10.6151
R1528 B.n959 B.n12 10.6151
R1529 B.n960 B.n959 10.6151
R1530 B.n961 B.n960 10.6151
R1531 B.n961 B.n10 10.6151
R1532 B.n965 B.n10 10.6151
R1533 B.n966 B.n965 10.6151
R1534 B.n967 B.n966 10.6151
R1535 B.n967 B.n8 10.6151
R1536 B.n971 B.n8 10.6151
R1537 B.n972 B.n971 10.6151
R1538 B.n973 B.n972 10.6151
R1539 B.n973 B.n6 10.6151
R1540 B.n977 B.n6 10.6151
R1541 B.n978 B.n977 10.6151
R1542 B.n979 B.n978 10.6151
R1543 B.n979 B.n4 10.6151
R1544 B.n983 B.n4 10.6151
R1545 B.n984 B.n983 10.6151
R1546 B.n985 B.n984 10.6151
R1547 B.n985 B.n0 10.6151
R1548 B.n859 B.n44 10.6151
R1549 B.n859 B.n858 10.6151
R1550 B.n858 B.n857 10.6151
R1551 B.n857 B.n46 10.6151
R1552 B.n853 B.n46 10.6151
R1553 B.n853 B.n852 10.6151
R1554 B.n852 B.n851 10.6151
R1555 B.n851 B.n48 10.6151
R1556 B.n847 B.n48 10.6151
R1557 B.n847 B.n846 10.6151
R1558 B.n846 B.n845 10.6151
R1559 B.n845 B.n50 10.6151
R1560 B.n841 B.n50 10.6151
R1561 B.n841 B.n840 10.6151
R1562 B.n840 B.n839 10.6151
R1563 B.n839 B.n52 10.6151
R1564 B.n835 B.n52 10.6151
R1565 B.n835 B.n834 10.6151
R1566 B.n834 B.n833 10.6151
R1567 B.n833 B.n54 10.6151
R1568 B.n829 B.n54 10.6151
R1569 B.n829 B.n828 10.6151
R1570 B.n828 B.n827 10.6151
R1571 B.n827 B.n56 10.6151
R1572 B.n823 B.n56 10.6151
R1573 B.n823 B.n822 10.6151
R1574 B.n822 B.n821 10.6151
R1575 B.n821 B.n58 10.6151
R1576 B.n817 B.n58 10.6151
R1577 B.n817 B.n816 10.6151
R1578 B.n816 B.n815 10.6151
R1579 B.n815 B.n60 10.6151
R1580 B.n811 B.n810 10.6151
R1581 B.n810 B.n809 10.6151
R1582 B.n809 B.n65 10.6151
R1583 B.n805 B.n65 10.6151
R1584 B.n805 B.n804 10.6151
R1585 B.n804 B.n803 10.6151
R1586 B.n803 B.n67 10.6151
R1587 B.n799 B.n67 10.6151
R1588 B.n797 B.n796 10.6151
R1589 B.n796 B.n71 10.6151
R1590 B.n792 B.n71 10.6151
R1591 B.n792 B.n791 10.6151
R1592 B.n791 B.n790 10.6151
R1593 B.n790 B.n73 10.6151
R1594 B.n786 B.n73 10.6151
R1595 B.n786 B.n785 10.6151
R1596 B.n785 B.n784 10.6151
R1597 B.n784 B.n75 10.6151
R1598 B.n780 B.n75 10.6151
R1599 B.n780 B.n779 10.6151
R1600 B.n779 B.n778 10.6151
R1601 B.n778 B.n77 10.6151
R1602 B.n774 B.n77 10.6151
R1603 B.n774 B.n773 10.6151
R1604 B.n773 B.n772 10.6151
R1605 B.n772 B.n79 10.6151
R1606 B.n768 B.n79 10.6151
R1607 B.n768 B.n767 10.6151
R1608 B.n767 B.n766 10.6151
R1609 B.n766 B.n81 10.6151
R1610 B.n762 B.n81 10.6151
R1611 B.n762 B.n761 10.6151
R1612 B.n761 B.n760 10.6151
R1613 B.n760 B.n83 10.6151
R1614 B.n756 B.n83 10.6151
R1615 B.n756 B.n755 10.6151
R1616 B.n755 B.n754 10.6151
R1617 B.n754 B.n85 10.6151
R1618 B.n750 B.n85 10.6151
R1619 B.n750 B.n749 10.6151
R1620 B.n748 B.n87 10.6151
R1621 B.n744 B.n87 10.6151
R1622 B.n744 B.n743 10.6151
R1623 B.n743 B.n742 10.6151
R1624 B.n742 B.n89 10.6151
R1625 B.n738 B.n89 10.6151
R1626 B.n738 B.n737 10.6151
R1627 B.n737 B.n736 10.6151
R1628 B.n736 B.n91 10.6151
R1629 B.n732 B.n91 10.6151
R1630 B.n732 B.n731 10.6151
R1631 B.n731 B.n730 10.6151
R1632 B.n730 B.n93 10.6151
R1633 B.n726 B.n93 10.6151
R1634 B.n726 B.n725 10.6151
R1635 B.n725 B.n724 10.6151
R1636 B.n724 B.n95 10.6151
R1637 B.n720 B.n95 10.6151
R1638 B.n720 B.n719 10.6151
R1639 B.n719 B.n718 10.6151
R1640 B.n718 B.n97 10.6151
R1641 B.n714 B.n97 10.6151
R1642 B.n714 B.n713 10.6151
R1643 B.n713 B.n712 10.6151
R1644 B.n712 B.n99 10.6151
R1645 B.n708 B.n99 10.6151
R1646 B.n708 B.n707 10.6151
R1647 B.n707 B.n706 10.6151
R1648 B.n706 B.n101 10.6151
R1649 B.n702 B.n101 10.6151
R1650 B.n702 B.n701 10.6151
R1651 B.n701 B.n700 10.6151
R1652 B.n700 B.n103 10.6151
R1653 B.n696 B.n103 10.6151
R1654 B.n696 B.n695 10.6151
R1655 B.n695 B.n694 10.6151
R1656 B.n694 B.n105 10.6151
R1657 B.n690 B.n105 10.6151
R1658 B.n690 B.n689 10.6151
R1659 B.n689 B.n688 10.6151
R1660 B.n688 B.n107 10.6151
R1661 B.n684 B.n107 10.6151
R1662 B.n684 B.n683 10.6151
R1663 B.n683 B.n682 10.6151
R1664 B.n682 B.n109 10.6151
R1665 B.n678 B.n109 10.6151
R1666 B.n678 B.n677 10.6151
R1667 B.n677 B.n676 10.6151
R1668 B.n676 B.n111 10.6151
R1669 B.n672 B.n111 10.6151
R1670 B.n672 B.n671 10.6151
R1671 B.n671 B.n670 10.6151
R1672 B.n670 B.n113 10.6151
R1673 B.n666 B.n113 10.6151
R1674 B.n666 B.n665 10.6151
R1675 B.n665 B.n664 10.6151
R1676 B.n664 B.n115 10.6151
R1677 B.n660 B.n115 10.6151
R1678 B.n660 B.n659 10.6151
R1679 B.n659 B.n658 10.6151
R1680 B.n658 B.n117 10.6151
R1681 B.n654 B.n117 10.6151
R1682 B.n654 B.n653 10.6151
R1683 B.n653 B.n652 10.6151
R1684 B.n652 B.n119 10.6151
R1685 B.n648 B.n119 10.6151
R1686 B.n648 B.n647 10.6151
R1687 B.n647 B.n646 10.6151
R1688 B.n646 B.n121 10.6151
R1689 B.n642 B.n121 10.6151
R1690 B.n642 B.n641 10.6151
R1691 B.n641 B.n640 10.6151
R1692 B.n640 B.n123 10.6151
R1693 B.n636 B.n123 10.6151
R1694 B.n636 B.n635 10.6151
R1695 B.n635 B.n634 10.6151
R1696 B.n634 B.n125 10.6151
R1697 B.n630 B.n125 10.6151
R1698 B.n630 B.n629 10.6151
R1699 B.n629 B.n628 10.6151
R1700 B.n628 B.n127 10.6151
R1701 B.n624 B.n127 10.6151
R1702 B.n624 B.n623 10.6151
R1703 B.n623 B.n622 10.6151
R1704 B.n622 B.n129 10.6151
R1705 B.n618 B.n129 10.6151
R1706 B.n618 B.n617 10.6151
R1707 B.n617 B.n616 10.6151
R1708 B.n616 B.n131 10.6151
R1709 B.n612 B.n131 10.6151
R1710 B.n612 B.n611 10.6151
R1711 B.n611 B.n610 10.6151
R1712 B.n610 B.n133 10.6151
R1713 B.n606 B.n133 10.6151
R1714 B.n606 B.n605 10.6151
R1715 B.n605 B.n604 10.6151
R1716 B.n604 B.n135 10.6151
R1717 B.n600 B.n135 10.6151
R1718 B.n600 B.n599 10.6151
R1719 B.n599 B.n598 10.6151
R1720 B.n598 B.n137 10.6151
R1721 B.n594 B.n137 10.6151
R1722 B.n594 B.n593 10.6151
R1723 B.n593 B.n592 10.6151
R1724 B.n592 B.n139 10.6151
R1725 B.n588 B.n139 10.6151
R1726 B.n588 B.n587 10.6151
R1727 B.n587 B.n586 10.6151
R1728 B.n586 B.n141 10.6151
R1729 B.n582 B.n141 10.6151
R1730 B.n582 B.n581 10.6151
R1731 B.n581 B.n580 10.6151
R1732 B.n580 B.n143 10.6151
R1733 B.n576 B.n143 10.6151
R1734 B.n576 B.n575 10.6151
R1735 B.n575 B.n574 10.6151
R1736 B.n574 B.n145 10.6151
R1737 B.n570 B.n145 10.6151
R1738 B.n570 B.n569 10.6151
R1739 B.n569 B.n568 10.6151
R1740 B.n568 B.n147 10.6151
R1741 B.n564 B.n147 10.6151
R1742 B.n564 B.n563 10.6151
R1743 B.n563 B.n562 10.6151
R1744 B.n562 B.n149 10.6151
R1745 B.n558 B.n149 10.6151
R1746 B.n558 B.n557 10.6151
R1747 B.n557 B.n556 10.6151
R1748 B.n556 B.n151 10.6151
R1749 B.n552 B.n151 10.6151
R1750 B.n552 B.n551 10.6151
R1751 B.n551 B.n550 10.6151
R1752 B.n550 B.n153 10.6151
R1753 B.n546 B.n153 10.6151
R1754 B.n546 B.n545 10.6151
R1755 B.n545 B.n544 10.6151
R1756 B.n544 B.n155 10.6151
R1757 B.n540 B.n155 10.6151
R1758 B.n540 B.n539 10.6151
R1759 B.n539 B.n538 10.6151
R1760 B.n538 B.n157 10.6151
R1761 B.n534 B.n157 10.6151
R1762 B.n534 B.n533 10.6151
R1763 B.n533 B.n532 10.6151
R1764 B.n532 B.n159 10.6151
R1765 B.n528 B.n159 10.6151
R1766 B.n528 B.n527 10.6151
R1767 B.n527 B.n526 10.6151
R1768 B.n526 B.n161 10.6151
R1769 B.n522 B.n161 10.6151
R1770 B.n522 B.n521 10.6151
R1771 B.n521 B.n520 10.6151
R1772 B.n520 B.n163 10.6151
R1773 B.n516 B.n163 10.6151
R1774 B.n516 B.n515 10.6151
R1775 B.n515 B.n514 10.6151
R1776 B.n514 B.n165 10.6151
R1777 B.n510 B.n165 10.6151
R1778 B.n510 B.n509 10.6151
R1779 B.n509 B.n508 10.6151
R1780 B.n508 B.n167 10.6151
R1781 B.n504 B.n167 10.6151
R1782 B.n504 B.n503 10.6151
R1783 B.n503 B.n502 10.6151
R1784 B.n502 B.n169 10.6151
R1785 B.n498 B.n169 10.6151
R1786 B.n498 B.n497 10.6151
R1787 B.n497 B.n496 10.6151
R1788 B.n496 B.n171 10.6151
R1789 B.n255 B.n1 10.6151
R1790 B.n256 B.n255 10.6151
R1791 B.n256 B.n253 10.6151
R1792 B.n260 B.n253 10.6151
R1793 B.n261 B.n260 10.6151
R1794 B.n262 B.n261 10.6151
R1795 B.n262 B.n251 10.6151
R1796 B.n266 B.n251 10.6151
R1797 B.n267 B.n266 10.6151
R1798 B.n268 B.n267 10.6151
R1799 B.n268 B.n249 10.6151
R1800 B.n272 B.n249 10.6151
R1801 B.n273 B.n272 10.6151
R1802 B.n274 B.n273 10.6151
R1803 B.n274 B.n247 10.6151
R1804 B.n278 B.n247 10.6151
R1805 B.n279 B.n278 10.6151
R1806 B.n280 B.n279 10.6151
R1807 B.n280 B.n245 10.6151
R1808 B.n284 B.n245 10.6151
R1809 B.n285 B.n284 10.6151
R1810 B.n286 B.n285 10.6151
R1811 B.n286 B.n243 10.6151
R1812 B.n290 B.n243 10.6151
R1813 B.n291 B.n290 10.6151
R1814 B.n292 B.n291 10.6151
R1815 B.n292 B.n241 10.6151
R1816 B.n296 B.n241 10.6151
R1817 B.n297 B.n296 10.6151
R1818 B.n298 B.n297 10.6151
R1819 B.n298 B.n239 10.6151
R1820 B.n302 B.n239 10.6151
R1821 B.n303 B.n302 10.6151
R1822 B.n304 B.n303 10.6151
R1823 B.n304 B.n237 10.6151
R1824 B.n308 B.n237 10.6151
R1825 B.n309 B.n308 10.6151
R1826 B.n310 B.n309 10.6151
R1827 B.n310 B.n235 10.6151
R1828 B.n314 B.n235 10.6151
R1829 B.n315 B.n314 10.6151
R1830 B.n316 B.n315 10.6151
R1831 B.n316 B.n233 10.6151
R1832 B.n320 B.n233 10.6151
R1833 B.n321 B.n320 10.6151
R1834 B.n322 B.n321 10.6151
R1835 B.n322 B.n231 10.6151
R1836 B.n326 B.n231 10.6151
R1837 B.n327 B.n326 10.6151
R1838 B.n328 B.n327 10.6151
R1839 B.n328 B.n229 10.6151
R1840 B.n332 B.n229 10.6151
R1841 B.n333 B.n332 10.6151
R1842 B.n334 B.n333 10.6151
R1843 B.n334 B.n227 10.6151
R1844 B.n338 B.n227 10.6151
R1845 B.n339 B.n338 10.6151
R1846 B.n340 B.n339 10.6151
R1847 B.n340 B.n225 10.6151
R1848 B.n344 B.n225 10.6151
R1849 B.n345 B.n344 10.6151
R1850 B.n346 B.n345 10.6151
R1851 B.n346 B.n223 10.6151
R1852 B.n350 B.n223 10.6151
R1853 B.n351 B.n350 10.6151
R1854 B.n352 B.n351 10.6151
R1855 B.n352 B.n221 10.6151
R1856 B.n356 B.n221 10.6151
R1857 B.n357 B.n356 10.6151
R1858 B.n358 B.n357 10.6151
R1859 B.n358 B.n219 10.6151
R1860 B.n362 B.n219 10.6151
R1861 B.n363 B.n362 10.6151
R1862 B.n364 B.n363 10.6151
R1863 B.n364 B.n217 10.6151
R1864 B.n368 B.n217 10.6151
R1865 B.n369 B.n368 10.6151
R1866 B.n370 B.n369 10.6151
R1867 B.n370 B.n215 10.6151
R1868 B.n374 B.n215 10.6151
R1869 B.n375 B.n374 10.6151
R1870 B.n376 B.n375 10.6151
R1871 B.n376 B.n213 10.6151
R1872 B.n381 B.n380 10.6151
R1873 B.n382 B.n381 10.6151
R1874 B.n382 B.n211 10.6151
R1875 B.n386 B.n211 10.6151
R1876 B.n387 B.n386 10.6151
R1877 B.n388 B.n387 10.6151
R1878 B.n388 B.n209 10.6151
R1879 B.n392 B.n209 10.6151
R1880 B.n393 B.n392 10.6151
R1881 B.n394 B.n393 10.6151
R1882 B.n394 B.n207 10.6151
R1883 B.n398 B.n207 10.6151
R1884 B.n399 B.n398 10.6151
R1885 B.n400 B.n399 10.6151
R1886 B.n400 B.n205 10.6151
R1887 B.n404 B.n205 10.6151
R1888 B.n405 B.n404 10.6151
R1889 B.n406 B.n405 10.6151
R1890 B.n406 B.n203 10.6151
R1891 B.n410 B.n203 10.6151
R1892 B.n411 B.n410 10.6151
R1893 B.n412 B.n411 10.6151
R1894 B.n412 B.n201 10.6151
R1895 B.n416 B.n201 10.6151
R1896 B.n417 B.n416 10.6151
R1897 B.n418 B.n417 10.6151
R1898 B.n418 B.n199 10.6151
R1899 B.n422 B.n199 10.6151
R1900 B.n423 B.n422 10.6151
R1901 B.n424 B.n423 10.6151
R1902 B.n424 B.n197 10.6151
R1903 B.n428 B.n197 10.6151
R1904 B.n431 B.n430 10.6151
R1905 B.n431 B.n193 10.6151
R1906 B.n435 B.n193 10.6151
R1907 B.n436 B.n435 10.6151
R1908 B.n437 B.n436 10.6151
R1909 B.n437 B.n191 10.6151
R1910 B.n441 B.n191 10.6151
R1911 B.n442 B.n441 10.6151
R1912 B.n444 B.n187 10.6151
R1913 B.n448 B.n187 10.6151
R1914 B.n449 B.n448 10.6151
R1915 B.n450 B.n449 10.6151
R1916 B.n450 B.n185 10.6151
R1917 B.n454 B.n185 10.6151
R1918 B.n455 B.n454 10.6151
R1919 B.n456 B.n455 10.6151
R1920 B.n456 B.n183 10.6151
R1921 B.n460 B.n183 10.6151
R1922 B.n461 B.n460 10.6151
R1923 B.n462 B.n461 10.6151
R1924 B.n462 B.n181 10.6151
R1925 B.n466 B.n181 10.6151
R1926 B.n467 B.n466 10.6151
R1927 B.n468 B.n467 10.6151
R1928 B.n468 B.n179 10.6151
R1929 B.n472 B.n179 10.6151
R1930 B.n473 B.n472 10.6151
R1931 B.n474 B.n473 10.6151
R1932 B.n474 B.n177 10.6151
R1933 B.n478 B.n177 10.6151
R1934 B.n479 B.n478 10.6151
R1935 B.n480 B.n479 10.6151
R1936 B.n480 B.n175 10.6151
R1937 B.n484 B.n175 10.6151
R1938 B.n485 B.n484 10.6151
R1939 B.n486 B.n485 10.6151
R1940 B.n486 B.n173 10.6151
R1941 B.n490 B.n173 10.6151
R1942 B.n491 B.n490 10.6151
R1943 B.n492 B.n491 10.6151
R1944 B.n989 B.n0 8.11757
R1945 B.n989 B.n1 8.11757
R1946 B.n811 B.n64 6.5566
R1947 B.n799 B.n798 6.5566
R1948 B.n430 B.n429 6.5566
R1949 B.n443 B.n442 6.5566
R1950 B.n64 B.n60 4.05904
R1951 B.n798 B.n797 4.05904
R1952 B.n429 B.n428 4.05904
R1953 B.n444 B.n443 4.05904
C0 VDD1 VP 9.374539f
C1 VDD2 B 2.95622f
C2 VDD1 VDD2 3.08666f
C3 w_n6166_n2778# B 12.0732f
C4 VN VP 9.918981f
C5 VDD1 w_n6166_n2778# 3.11603f
C6 VN VDD2 8.77274f
C7 VTAIL VP 10.1733f
C8 w_n6166_n2778# VN 13.562599f
C9 VDD1 B 2.78379f
C10 VTAIL VDD2 10.1078f
C11 VN B 1.60485f
C12 w_n6166_n2778# VTAIL 3.01853f
C13 VDD1 VN 0.156594f
C14 VTAIL B 3.53913f
C15 VP VDD2 0.761612f
C16 VDD1 VTAIL 10.046f
C17 w_n6166_n2778# VP 14.3697f
C18 VTAIL VN 10.1586f
C19 w_n6166_n2778# VDD2 3.33234f
C20 VP B 2.96976f
C21 VDD2 VSUBS 2.67429f
C22 VDD1 VSUBS 2.496707f
C23 VTAIL VSUBS 1.552105f
C24 VN VSUBS 10.06764f
C25 VP VSUBS 5.938691f
C26 B VSUBS 6.852836f
C27 w_n6166_n2778# VSUBS 0.211987p
C28 B.n0 VSUBS 0.008672f
C29 B.n1 VSUBS 0.008672f
C30 B.n2 VSUBS 0.012825f
C31 B.n3 VSUBS 0.009828f
C32 B.n4 VSUBS 0.009828f
C33 B.n5 VSUBS 0.009828f
C34 B.n6 VSUBS 0.009828f
C35 B.n7 VSUBS 0.009828f
C36 B.n8 VSUBS 0.009828f
C37 B.n9 VSUBS 0.009828f
C38 B.n10 VSUBS 0.009828f
C39 B.n11 VSUBS 0.009828f
C40 B.n12 VSUBS 0.009828f
C41 B.n13 VSUBS 0.009828f
C42 B.n14 VSUBS 0.009828f
C43 B.n15 VSUBS 0.009828f
C44 B.n16 VSUBS 0.009828f
C45 B.n17 VSUBS 0.009828f
C46 B.n18 VSUBS 0.009828f
C47 B.n19 VSUBS 0.009828f
C48 B.n20 VSUBS 0.009828f
C49 B.n21 VSUBS 0.009828f
C50 B.n22 VSUBS 0.009828f
C51 B.n23 VSUBS 0.009828f
C52 B.n24 VSUBS 0.009828f
C53 B.n25 VSUBS 0.009828f
C54 B.n26 VSUBS 0.009828f
C55 B.n27 VSUBS 0.009828f
C56 B.n28 VSUBS 0.009828f
C57 B.n29 VSUBS 0.009828f
C58 B.n30 VSUBS 0.009828f
C59 B.n31 VSUBS 0.009828f
C60 B.n32 VSUBS 0.009828f
C61 B.n33 VSUBS 0.009828f
C62 B.n34 VSUBS 0.009828f
C63 B.n35 VSUBS 0.009828f
C64 B.n36 VSUBS 0.009828f
C65 B.n37 VSUBS 0.009828f
C66 B.n38 VSUBS 0.009828f
C67 B.n39 VSUBS 0.009828f
C68 B.n40 VSUBS 0.009828f
C69 B.n41 VSUBS 0.009828f
C70 B.n42 VSUBS 0.009828f
C71 B.n43 VSUBS 0.009828f
C72 B.n44 VSUBS 0.024465f
C73 B.n45 VSUBS 0.009828f
C74 B.n46 VSUBS 0.009828f
C75 B.n47 VSUBS 0.009828f
C76 B.n48 VSUBS 0.009828f
C77 B.n49 VSUBS 0.009828f
C78 B.n50 VSUBS 0.009828f
C79 B.n51 VSUBS 0.009828f
C80 B.n52 VSUBS 0.009828f
C81 B.n53 VSUBS 0.009828f
C82 B.n54 VSUBS 0.009828f
C83 B.n55 VSUBS 0.009828f
C84 B.n56 VSUBS 0.009828f
C85 B.n57 VSUBS 0.009828f
C86 B.n58 VSUBS 0.009828f
C87 B.n59 VSUBS 0.009828f
C88 B.n60 VSUBS 0.006793f
C89 B.n61 VSUBS 0.009828f
C90 B.t7 VSUBS 0.399655f
C91 B.t8 VSUBS 0.440151f
C92 B.t6 VSUBS 2.40914f
C93 B.n62 VSUBS 0.255137f
C94 B.n63 VSUBS 0.108589f
C95 B.n64 VSUBS 0.02277f
C96 B.n65 VSUBS 0.009828f
C97 B.n66 VSUBS 0.009828f
C98 B.n67 VSUBS 0.009828f
C99 B.n68 VSUBS 0.009828f
C100 B.t4 VSUBS 0.399651f
C101 B.t5 VSUBS 0.440147f
C102 B.t3 VSUBS 2.40914f
C103 B.n69 VSUBS 0.255141f
C104 B.n70 VSUBS 0.108594f
C105 B.n71 VSUBS 0.009828f
C106 B.n72 VSUBS 0.009828f
C107 B.n73 VSUBS 0.009828f
C108 B.n74 VSUBS 0.009828f
C109 B.n75 VSUBS 0.009828f
C110 B.n76 VSUBS 0.009828f
C111 B.n77 VSUBS 0.009828f
C112 B.n78 VSUBS 0.009828f
C113 B.n79 VSUBS 0.009828f
C114 B.n80 VSUBS 0.009828f
C115 B.n81 VSUBS 0.009828f
C116 B.n82 VSUBS 0.009828f
C117 B.n83 VSUBS 0.009828f
C118 B.n84 VSUBS 0.009828f
C119 B.n85 VSUBS 0.009828f
C120 B.n86 VSUBS 0.024465f
C121 B.n87 VSUBS 0.009828f
C122 B.n88 VSUBS 0.009828f
C123 B.n89 VSUBS 0.009828f
C124 B.n90 VSUBS 0.009828f
C125 B.n91 VSUBS 0.009828f
C126 B.n92 VSUBS 0.009828f
C127 B.n93 VSUBS 0.009828f
C128 B.n94 VSUBS 0.009828f
C129 B.n95 VSUBS 0.009828f
C130 B.n96 VSUBS 0.009828f
C131 B.n97 VSUBS 0.009828f
C132 B.n98 VSUBS 0.009828f
C133 B.n99 VSUBS 0.009828f
C134 B.n100 VSUBS 0.009828f
C135 B.n101 VSUBS 0.009828f
C136 B.n102 VSUBS 0.009828f
C137 B.n103 VSUBS 0.009828f
C138 B.n104 VSUBS 0.009828f
C139 B.n105 VSUBS 0.009828f
C140 B.n106 VSUBS 0.009828f
C141 B.n107 VSUBS 0.009828f
C142 B.n108 VSUBS 0.009828f
C143 B.n109 VSUBS 0.009828f
C144 B.n110 VSUBS 0.009828f
C145 B.n111 VSUBS 0.009828f
C146 B.n112 VSUBS 0.009828f
C147 B.n113 VSUBS 0.009828f
C148 B.n114 VSUBS 0.009828f
C149 B.n115 VSUBS 0.009828f
C150 B.n116 VSUBS 0.009828f
C151 B.n117 VSUBS 0.009828f
C152 B.n118 VSUBS 0.009828f
C153 B.n119 VSUBS 0.009828f
C154 B.n120 VSUBS 0.009828f
C155 B.n121 VSUBS 0.009828f
C156 B.n122 VSUBS 0.009828f
C157 B.n123 VSUBS 0.009828f
C158 B.n124 VSUBS 0.009828f
C159 B.n125 VSUBS 0.009828f
C160 B.n126 VSUBS 0.009828f
C161 B.n127 VSUBS 0.009828f
C162 B.n128 VSUBS 0.009828f
C163 B.n129 VSUBS 0.009828f
C164 B.n130 VSUBS 0.009828f
C165 B.n131 VSUBS 0.009828f
C166 B.n132 VSUBS 0.009828f
C167 B.n133 VSUBS 0.009828f
C168 B.n134 VSUBS 0.009828f
C169 B.n135 VSUBS 0.009828f
C170 B.n136 VSUBS 0.009828f
C171 B.n137 VSUBS 0.009828f
C172 B.n138 VSUBS 0.009828f
C173 B.n139 VSUBS 0.009828f
C174 B.n140 VSUBS 0.009828f
C175 B.n141 VSUBS 0.009828f
C176 B.n142 VSUBS 0.009828f
C177 B.n143 VSUBS 0.009828f
C178 B.n144 VSUBS 0.009828f
C179 B.n145 VSUBS 0.009828f
C180 B.n146 VSUBS 0.009828f
C181 B.n147 VSUBS 0.009828f
C182 B.n148 VSUBS 0.009828f
C183 B.n149 VSUBS 0.009828f
C184 B.n150 VSUBS 0.009828f
C185 B.n151 VSUBS 0.009828f
C186 B.n152 VSUBS 0.009828f
C187 B.n153 VSUBS 0.009828f
C188 B.n154 VSUBS 0.009828f
C189 B.n155 VSUBS 0.009828f
C190 B.n156 VSUBS 0.009828f
C191 B.n157 VSUBS 0.009828f
C192 B.n158 VSUBS 0.009828f
C193 B.n159 VSUBS 0.009828f
C194 B.n160 VSUBS 0.009828f
C195 B.n161 VSUBS 0.009828f
C196 B.n162 VSUBS 0.009828f
C197 B.n163 VSUBS 0.009828f
C198 B.n164 VSUBS 0.009828f
C199 B.n165 VSUBS 0.009828f
C200 B.n166 VSUBS 0.009828f
C201 B.n167 VSUBS 0.009828f
C202 B.n168 VSUBS 0.009828f
C203 B.n169 VSUBS 0.009828f
C204 B.n170 VSUBS 0.009828f
C205 B.n171 VSUBS 0.024887f
C206 B.n172 VSUBS 0.009828f
C207 B.n173 VSUBS 0.009828f
C208 B.n174 VSUBS 0.009828f
C209 B.n175 VSUBS 0.009828f
C210 B.n176 VSUBS 0.009828f
C211 B.n177 VSUBS 0.009828f
C212 B.n178 VSUBS 0.009828f
C213 B.n179 VSUBS 0.009828f
C214 B.n180 VSUBS 0.009828f
C215 B.n181 VSUBS 0.009828f
C216 B.n182 VSUBS 0.009828f
C217 B.n183 VSUBS 0.009828f
C218 B.n184 VSUBS 0.009828f
C219 B.n185 VSUBS 0.009828f
C220 B.n186 VSUBS 0.009828f
C221 B.n187 VSUBS 0.009828f
C222 B.n188 VSUBS 0.009828f
C223 B.t11 VSUBS 0.399651f
C224 B.t10 VSUBS 0.440147f
C225 B.t9 VSUBS 2.40914f
C226 B.n189 VSUBS 0.255141f
C227 B.n190 VSUBS 0.108594f
C228 B.n191 VSUBS 0.009828f
C229 B.n192 VSUBS 0.009828f
C230 B.n193 VSUBS 0.009828f
C231 B.n194 VSUBS 0.009828f
C232 B.t2 VSUBS 0.399655f
C233 B.t1 VSUBS 0.440151f
C234 B.t0 VSUBS 2.40914f
C235 B.n195 VSUBS 0.255137f
C236 B.n196 VSUBS 0.108589f
C237 B.n197 VSUBS 0.009828f
C238 B.n198 VSUBS 0.009828f
C239 B.n199 VSUBS 0.009828f
C240 B.n200 VSUBS 0.009828f
C241 B.n201 VSUBS 0.009828f
C242 B.n202 VSUBS 0.009828f
C243 B.n203 VSUBS 0.009828f
C244 B.n204 VSUBS 0.009828f
C245 B.n205 VSUBS 0.009828f
C246 B.n206 VSUBS 0.009828f
C247 B.n207 VSUBS 0.009828f
C248 B.n208 VSUBS 0.009828f
C249 B.n209 VSUBS 0.009828f
C250 B.n210 VSUBS 0.009828f
C251 B.n211 VSUBS 0.009828f
C252 B.n212 VSUBS 0.009828f
C253 B.n213 VSUBS 0.023807f
C254 B.n214 VSUBS 0.009828f
C255 B.n215 VSUBS 0.009828f
C256 B.n216 VSUBS 0.009828f
C257 B.n217 VSUBS 0.009828f
C258 B.n218 VSUBS 0.009828f
C259 B.n219 VSUBS 0.009828f
C260 B.n220 VSUBS 0.009828f
C261 B.n221 VSUBS 0.009828f
C262 B.n222 VSUBS 0.009828f
C263 B.n223 VSUBS 0.009828f
C264 B.n224 VSUBS 0.009828f
C265 B.n225 VSUBS 0.009828f
C266 B.n226 VSUBS 0.009828f
C267 B.n227 VSUBS 0.009828f
C268 B.n228 VSUBS 0.009828f
C269 B.n229 VSUBS 0.009828f
C270 B.n230 VSUBS 0.009828f
C271 B.n231 VSUBS 0.009828f
C272 B.n232 VSUBS 0.009828f
C273 B.n233 VSUBS 0.009828f
C274 B.n234 VSUBS 0.009828f
C275 B.n235 VSUBS 0.009828f
C276 B.n236 VSUBS 0.009828f
C277 B.n237 VSUBS 0.009828f
C278 B.n238 VSUBS 0.009828f
C279 B.n239 VSUBS 0.009828f
C280 B.n240 VSUBS 0.009828f
C281 B.n241 VSUBS 0.009828f
C282 B.n242 VSUBS 0.009828f
C283 B.n243 VSUBS 0.009828f
C284 B.n244 VSUBS 0.009828f
C285 B.n245 VSUBS 0.009828f
C286 B.n246 VSUBS 0.009828f
C287 B.n247 VSUBS 0.009828f
C288 B.n248 VSUBS 0.009828f
C289 B.n249 VSUBS 0.009828f
C290 B.n250 VSUBS 0.009828f
C291 B.n251 VSUBS 0.009828f
C292 B.n252 VSUBS 0.009828f
C293 B.n253 VSUBS 0.009828f
C294 B.n254 VSUBS 0.009828f
C295 B.n255 VSUBS 0.009828f
C296 B.n256 VSUBS 0.009828f
C297 B.n257 VSUBS 0.009828f
C298 B.n258 VSUBS 0.009828f
C299 B.n259 VSUBS 0.009828f
C300 B.n260 VSUBS 0.009828f
C301 B.n261 VSUBS 0.009828f
C302 B.n262 VSUBS 0.009828f
C303 B.n263 VSUBS 0.009828f
C304 B.n264 VSUBS 0.009828f
C305 B.n265 VSUBS 0.009828f
C306 B.n266 VSUBS 0.009828f
C307 B.n267 VSUBS 0.009828f
C308 B.n268 VSUBS 0.009828f
C309 B.n269 VSUBS 0.009828f
C310 B.n270 VSUBS 0.009828f
C311 B.n271 VSUBS 0.009828f
C312 B.n272 VSUBS 0.009828f
C313 B.n273 VSUBS 0.009828f
C314 B.n274 VSUBS 0.009828f
C315 B.n275 VSUBS 0.009828f
C316 B.n276 VSUBS 0.009828f
C317 B.n277 VSUBS 0.009828f
C318 B.n278 VSUBS 0.009828f
C319 B.n279 VSUBS 0.009828f
C320 B.n280 VSUBS 0.009828f
C321 B.n281 VSUBS 0.009828f
C322 B.n282 VSUBS 0.009828f
C323 B.n283 VSUBS 0.009828f
C324 B.n284 VSUBS 0.009828f
C325 B.n285 VSUBS 0.009828f
C326 B.n286 VSUBS 0.009828f
C327 B.n287 VSUBS 0.009828f
C328 B.n288 VSUBS 0.009828f
C329 B.n289 VSUBS 0.009828f
C330 B.n290 VSUBS 0.009828f
C331 B.n291 VSUBS 0.009828f
C332 B.n292 VSUBS 0.009828f
C333 B.n293 VSUBS 0.009828f
C334 B.n294 VSUBS 0.009828f
C335 B.n295 VSUBS 0.009828f
C336 B.n296 VSUBS 0.009828f
C337 B.n297 VSUBS 0.009828f
C338 B.n298 VSUBS 0.009828f
C339 B.n299 VSUBS 0.009828f
C340 B.n300 VSUBS 0.009828f
C341 B.n301 VSUBS 0.009828f
C342 B.n302 VSUBS 0.009828f
C343 B.n303 VSUBS 0.009828f
C344 B.n304 VSUBS 0.009828f
C345 B.n305 VSUBS 0.009828f
C346 B.n306 VSUBS 0.009828f
C347 B.n307 VSUBS 0.009828f
C348 B.n308 VSUBS 0.009828f
C349 B.n309 VSUBS 0.009828f
C350 B.n310 VSUBS 0.009828f
C351 B.n311 VSUBS 0.009828f
C352 B.n312 VSUBS 0.009828f
C353 B.n313 VSUBS 0.009828f
C354 B.n314 VSUBS 0.009828f
C355 B.n315 VSUBS 0.009828f
C356 B.n316 VSUBS 0.009828f
C357 B.n317 VSUBS 0.009828f
C358 B.n318 VSUBS 0.009828f
C359 B.n319 VSUBS 0.009828f
C360 B.n320 VSUBS 0.009828f
C361 B.n321 VSUBS 0.009828f
C362 B.n322 VSUBS 0.009828f
C363 B.n323 VSUBS 0.009828f
C364 B.n324 VSUBS 0.009828f
C365 B.n325 VSUBS 0.009828f
C366 B.n326 VSUBS 0.009828f
C367 B.n327 VSUBS 0.009828f
C368 B.n328 VSUBS 0.009828f
C369 B.n329 VSUBS 0.009828f
C370 B.n330 VSUBS 0.009828f
C371 B.n331 VSUBS 0.009828f
C372 B.n332 VSUBS 0.009828f
C373 B.n333 VSUBS 0.009828f
C374 B.n334 VSUBS 0.009828f
C375 B.n335 VSUBS 0.009828f
C376 B.n336 VSUBS 0.009828f
C377 B.n337 VSUBS 0.009828f
C378 B.n338 VSUBS 0.009828f
C379 B.n339 VSUBS 0.009828f
C380 B.n340 VSUBS 0.009828f
C381 B.n341 VSUBS 0.009828f
C382 B.n342 VSUBS 0.009828f
C383 B.n343 VSUBS 0.009828f
C384 B.n344 VSUBS 0.009828f
C385 B.n345 VSUBS 0.009828f
C386 B.n346 VSUBS 0.009828f
C387 B.n347 VSUBS 0.009828f
C388 B.n348 VSUBS 0.009828f
C389 B.n349 VSUBS 0.009828f
C390 B.n350 VSUBS 0.009828f
C391 B.n351 VSUBS 0.009828f
C392 B.n352 VSUBS 0.009828f
C393 B.n353 VSUBS 0.009828f
C394 B.n354 VSUBS 0.009828f
C395 B.n355 VSUBS 0.009828f
C396 B.n356 VSUBS 0.009828f
C397 B.n357 VSUBS 0.009828f
C398 B.n358 VSUBS 0.009828f
C399 B.n359 VSUBS 0.009828f
C400 B.n360 VSUBS 0.009828f
C401 B.n361 VSUBS 0.009828f
C402 B.n362 VSUBS 0.009828f
C403 B.n363 VSUBS 0.009828f
C404 B.n364 VSUBS 0.009828f
C405 B.n365 VSUBS 0.009828f
C406 B.n366 VSUBS 0.009828f
C407 B.n367 VSUBS 0.009828f
C408 B.n368 VSUBS 0.009828f
C409 B.n369 VSUBS 0.009828f
C410 B.n370 VSUBS 0.009828f
C411 B.n371 VSUBS 0.009828f
C412 B.n372 VSUBS 0.009828f
C413 B.n373 VSUBS 0.009828f
C414 B.n374 VSUBS 0.009828f
C415 B.n375 VSUBS 0.009828f
C416 B.n376 VSUBS 0.009828f
C417 B.n377 VSUBS 0.009828f
C418 B.n378 VSUBS 0.023807f
C419 B.n379 VSUBS 0.024465f
C420 B.n380 VSUBS 0.024465f
C421 B.n381 VSUBS 0.009828f
C422 B.n382 VSUBS 0.009828f
C423 B.n383 VSUBS 0.009828f
C424 B.n384 VSUBS 0.009828f
C425 B.n385 VSUBS 0.009828f
C426 B.n386 VSUBS 0.009828f
C427 B.n387 VSUBS 0.009828f
C428 B.n388 VSUBS 0.009828f
C429 B.n389 VSUBS 0.009828f
C430 B.n390 VSUBS 0.009828f
C431 B.n391 VSUBS 0.009828f
C432 B.n392 VSUBS 0.009828f
C433 B.n393 VSUBS 0.009828f
C434 B.n394 VSUBS 0.009828f
C435 B.n395 VSUBS 0.009828f
C436 B.n396 VSUBS 0.009828f
C437 B.n397 VSUBS 0.009828f
C438 B.n398 VSUBS 0.009828f
C439 B.n399 VSUBS 0.009828f
C440 B.n400 VSUBS 0.009828f
C441 B.n401 VSUBS 0.009828f
C442 B.n402 VSUBS 0.009828f
C443 B.n403 VSUBS 0.009828f
C444 B.n404 VSUBS 0.009828f
C445 B.n405 VSUBS 0.009828f
C446 B.n406 VSUBS 0.009828f
C447 B.n407 VSUBS 0.009828f
C448 B.n408 VSUBS 0.009828f
C449 B.n409 VSUBS 0.009828f
C450 B.n410 VSUBS 0.009828f
C451 B.n411 VSUBS 0.009828f
C452 B.n412 VSUBS 0.009828f
C453 B.n413 VSUBS 0.009828f
C454 B.n414 VSUBS 0.009828f
C455 B.n415 VSUBS 0.009828f
C456 B.n416 VSUBS 0.009828f
C457 B.n417 VSUBS 0.009828f
C458 B.n418 VSUBS 0.009828f
C459 B.n419 VSUBS 0.009828f
C460 B.n420 VSUBS 0.009828f
C461 B.n421 VSUBS 0.009828f
C462 B.n422 VSUBS 0.009828f
C463 B.n423 VSUBS 0.009828f
C464 B.n424 VSUBS 0.009828f
C465 B.n425 VSUBS 0.009828f
C466 B.n426 VSUBS 0.009828f
C467 B.n427 VSUBS 0.009828f
C468 B.n428 VSUBS 0.006793f
C469 B.n429 VSUBS 0.02277f
C470 B.n430 VSUBS 0.007949f
C471 B.n431 VSUBS 0.009828f
C472 B.n432 VSUBS 0.009828f
C473 B.n433 VSUBS 0.009828f
C474 B.n434 VSUBS 0.009828f
C475 B.n435 VSUBS 0.009828f
C476 B.n436 VSUBS 0.009828f
C477 B.n437 VSUBS 0.009828f
C478 B.n438 VSUBS 0.009828f
C479 B.n439 VSUBS 0.009828f
C480 B.n440 VSUBS 0.009828f
C481 B.n441 VSUBS 0.009828f
C482 B.n442 VSUBS 0.007949f
C483 B.n443 VSUBS 0.02277f
C484 B.n444 VSUBS 0.006793f
C485 B.n445 VSUBS 0.009828f
C486 B.n446 VSUBS 0.009828f
C487 B.n447 VSUBS 0.009828f
C488 B.n448 VSUBS 0.009828f
C489 B.n449 VSUBS 0.009828f
C490 B.n450 VSUBS 0.009828f
C491 B.n451 VSUBS 0.009828f
C492 B.n452 VSUBS 0.009828f
C493 B.n453 VSUBS 0.009828f
C494 B.n454 VSUBS 0.009828f
C495 B.n455 VSUBS 0.009828f
C496 B.n456 VSUBS 0.009828f
C497 B.n457 VSUBS 0.009828f
C498 B.n458 VSUBS 0.009828f
C499 B.n459 VSUBS 0.009828f
C500 B.n460 VSUBS 0.009828f
C501 B.n461 VSUBS 0.009828f
C502 B.n462 VSUBS 0.009828f
C503 B.n463 VSUBS 0.009828f
C504 B.n464 VSUBS 0.009828f
C505 B.n465 VSUBS 0.009828f
C506 B.n466 VSUBS 0.009828f
C507 B.n467 VSUBS 0.009828f
C508 B.n468 VSUBS 0.009828f
C509 B.n469 VSUBS 0.009828f
C510 B.n470 VSUBS 0.009828f
C511 B.n471 VSUBS 0.009828f
C512 B.n472 VSUBS 0.009828f
C513 B.n473 VSUBS 0.009828f
C514 B.n474 VSUBS 0.009828f
C515 B.n475 VSUBS 0.009828f
C516 B.n476 VSUBS 0.009828f
C517 B.n477 VSUBS 0.009828f
C518 B.n478 VSUBS 0.009828f
C519 B.n479 VSUBS 0.009828f
C520 B.n480 VSUBS 0.009828f
C521 B.n481 VSUBS 0.009828f
C522 B.n482 VSUBS 0.009828f
C523 B.n483 VSUBS 0.009828f
C524 B.n484 VSUBS 0.009828f
C525 B.n485 VSUBS 0.009828f
C526 B.n486 VSUBS 0.009828f
C527 B.n487 VSUBS 0.009828f
C528 B.n488 VSUBS 0.009828f
C529 B.n489 VSUBS 0.009828f
C530 B.n490 VSUBS 0.009828f
C531 B.n491 VSUBS 0.009828f
C532 B.n492 VSUBS 0.023386f
C533 B.n493 VSUBS 0.024465f
C534 B.n494 VSUBS 0.023807f
C535 B.n495 VSUBS 0.009828f
C536 B.n496 VSUBS 0.009828f
C537 B.n497 VSUBS 0.009828f
C538 B.n498 VSUBS 0.009828f
C539 B.n499 VSUBS 0.009828f
C540 B.n500 VSUBS 0.009828f
C541 B.n501 VSUBS 0.009828f
C542 B.n502 VSUBS 0.009828f
C543 B.n503 VSUBS 0.009828f
C544 B.n504 VSUBS 0.009828f
C545 B.n505 VSUBS 0.009828f
C546 B.n506 VSUBS 0.009828f
C547 B.n507 VSUBS 0.009828f
C548 B.n508 VSUBS 0.009828f
C549 B.n509 VSUBS 0.009828f
C550 B.n510 VSUBS 0.009828f
C551 B.n511 VSUBS 0.009828f
C552 B.n512 VSUBS 0.009828f
C553 B.n513 VSUBS 0.009828f
C554 B.n514 VSUBS 0.009828f
C555 B.n515 VSUBS 0.009828f
C556 B.n516 VSUBS 0.009828f
C557 B.n517 VSUBS 0.009828f
C558 B.n518 VSUBS 0.009828f
C559 B.n519 VSUBS 0.009828f
C560 B.n520 VSUBS 0.009828f
C561 B.n521 VSUBS 0.009828f
C562 B.n522 VSUBS 0.009828f
C563 B.n523 VSUBS 0.009828f
C564 B.n524 VSUBS 0.009828f
C565 B.n525 VSUBS 0.009828f
C566 B.n526 VSUBS 0.009828f
C567 B.n527 VSUBS 0.009828f
C568 B.n528 VSUBS 0.009828f
C569 B.n529 VSUBS 0.009828f
C570 B.n530 VSUBS 0.009828f
C571 B.n531 VSUBS 0.009828f
C572 B.n532 VSUBS 0.009828f
C573 B.n533 VSUBS 0.009828f
C574 B.n534 VSUBS 0.009828f
C575 B.n535 VSUBS 0.009828f
C576 B.n536 VSUBS 0.009828f
C577 B.n537 VSUBS 0.009828f
C578 B.n538 VSUBS 0.009828f
C579 B.n539 VSUBS 0.009828f
C580 B.n540 VSUBS 0.009828f
C581 B.n541 VSUBS 0.009828f
C582 B.n542 VSUBS 0.009828f
C583 B.n543 VSUBS 0.009828f
C584 B.n544 VSUBS 0.009828f
C585 B.n545 VSUBS 0.009828f
C586 B.n546 VSUBS 0.009828f
C587 B.n547 VSUBS 0.009828f
C588 B.n548 VSUBS 0.009828f
C589 B.n549 VSUBS 0.009828f
C590 B.n550 VSUBS 0.009828f
C591 B.n551 VSUBS 0.009828f
C592 B.n552 VSUBS 0.009828f
C593 B.n553 VSUBS 0.009828f
C594 B.n554 VSUBS 0.009828f
C595 B.n555 VSUBS 0.009828f
C596 B.n556 VSUBS 0.009828f
C597 B.n557 VSUBS 0.009828f
C598 B.n558 VSUBS 0.009828f
C599 B.n559 VSUBS 0.009828f
C600 B.n560 VSUBS 0.009828f
C601 B.n561 VSUBS 0.009828f
C602 B.n562 VSUBS 0.009828f
C603 B.n563 VSUBS 0.009828f
C604 B.n564 VSUBS 0.009828f
C605 B.n565 VSUBS 0.009828f
C606 B.n566 VSUBS 0.009828f
C607 B.n567 VSUBS 0.009828f
C608 B.n568 VSUBS 0.009828f
C609 B.n569 VSUBS 0.009828f
C610 B.n570 VSUBS 0.009828f
C611 B.n571 VSUBS 0.009828f
C612 B.n572 VSUBS 0.009828f
C613 B.n573 VSUBS 0.009828f
C614 B.n574 VSUBS 0.009828f
C615 B.n575 VSUBS 0.009828f
C616 B.n576 VSUBS 0.009828f
C617 B.n577 VSUBS 0.009828f
C618 B.n578 VSUBS 0.009828f
C619 B.n579 VSUBS 0.009828f
C620 B.n580 VSUBS 0.009828f
C621 B.n581 VSUBS 0.009828f
C622 B.n582 VSUBS 0.009828f
C623 B.n583 VSUBS 0.009828f
C624 B.n584 VSUBS 0.009828f
C625 B.n585 VSUBS 0.009828f
C626 B.n586 VSUBS 0.009828f
C627 B.n587 VSUBS 0.009828f
C628 B.n588 VSUBS 0.009828f
C629 B.n589 VSUBS 0.009828f
C630 B.n590 VSUBS 0.009828f
C631 B.n591 VSUBS 0.009828f
C632 B.n592 VSUBS 0.009828f
C633 B.n593 VSUBS 0.009828f
C634 B.n594 VSUBS 0.009828f
C635 B.n595 VSUBS 0.009828f
C636 B.n596 VSUBS 0.009828f
C637 B.n597 VSUBS 0.009828f
C638 B.n598 VSUBS 0.009828f
C639 B.n599 VSUBS 0.009828f
C640 B.n600 VSUBS 0.009828f
C641 B.n601 VSUBS 0.009828f
C642 B.n602 VSUBS 0.009828f
C643 B.n603 VSUBS 0.009828f
C644 B.n604 VSUBS 0.009828f
C645 B.n605 VSUBS 0.009828f
C646 B.n606 VSUBS 0.009828f
C647 B.n607 VSUBS 0.009828f
C648 B.n608 VSUBS 0.009828f
C649 B.n609 VSUBS 0.009828f
C650 B.n610 VSUBS 0.009828f
C651 B.n611 VSUBS 0.009828f
C652 B.n612 VSUBS 0.009828f
C653 B.n613 VSUBS 0.009828f
C654 B.n614 VSUBS 0.009828f
C655 B.n615 VSUBS 0.009828f
C656 B.n616 VSUBS 0.009828f
C657 B.n617 VSUBS 0.009828f
C658 B.n618 VSUBS 0.009828f
C659 B.n619 VSUBS 0.009828f
C660 B.n620 VSUBS 0.009828f
C661 B.n621 VSUBS 0.009828f
C662 B.n622 VSUBS 0.009828f
C663 B.n623 VSUBS 0.009828f
C664 B.n624 VSUBS 0.009828f
C665 B.n625 VSUBS 0.009828f
C666 B.n626 VSUBS 0.009828f
C667 B.n627 VSUBS 0.009828f
C668 B.n628 VSUBS 0.009828f
C669 B.n629 VSUBS 0.009828f
C670 B.n630 VSUBS 0.009828f
C671 B.n631 VSUBS 0.009828f
C672 B.n632 VSUBS 0.009828f
C673 B.n633 VSUBS 0.009828f
C674 B.n634 VSUBS 0.009828f
C675 B.n635 VSUBS 0.009828f
C676 B.n636 VSUBS 0.009828f
C677 B.n637 VSUBS 0.009828f
C678 B.n638 VSUBS 0.009828f
C679 B.n639 VSUBS 0.009828f
C680 B.n640 VSUBS 0.009828f
C681 B.n641 VSUBS 0.009828f
C682 B.n642 VSUBS 0.009828f
C683 B.n643 VSUBS 0.009828f
C684 B.n644 VSUBS 0.009828f
C685 B.n645 VSUBS 0.009828f
C686 B.n646 VSUBS 0.009828f
C687 B.n647 VSUBS 0.009828f
C688 B.n648 VSUBS 0.009828f
C689 B.n649 VSUBS 0.009828f
C690 B.n650 VSUBS 0.009828f
C691 B.n651 VSUBS 0.009828f
C692 B.n652 VSUBS 0.009828f
C693 B.n653 VSUBS 0.009828f
C694 B.n654 VSUBS 0.009828f
C695 B.n655 VSUBS 0.009828f
C696 B.n656 VSUBS 0.009828f
C697 B.n657 VSUBS 0.009828f
C698 B.n658 VSUBS 0.009828f
C699 B.n659 VSUBS 0.009828f
C700 B.n660 VSUBS 0.009828f
C701 B.n661 VSUBS 0.009828f
C702 B.n662 VSUBS 0.009828f
C703 B.n663 VSUBS 0.009828f
C704 B.n664 VSUBS 0.009828f
C705 B.n665 VSUBS 0.009828f
C706 B.n666 VSUBS 0.009828f
C707 B.n667 VSUBS 0.009828f
C708 B.n668 VSUBS 0.009828f
C709 B.n669 VSUBS 0.009828f
C710 B.n670 VSUBS 0.009828f
C711 B.n671 VSUBS 0.009828f
C712 B.n672 VSUBS 0.009828f
C713 B.n673 VSUBS 0.009828f
C714 B.n674 VSUBS 0.009828f
C715 B.n675 VSUBS 0.009828f
C716 B.n676 VSUBS 0.009828f
C717 B.n677 VSUBS 0.009828f
C718 B.n678 VSUBS 0.009828f
C719 B.n679 VSUBS 0.009828f
C720 B.n680 VSUBS 0.009828f
C721 B.n681 VSUBS 0.009828f
C722 B.n682 VSUBS 0.009828f
C723 B.n683 VSUBS 0.009828f
C724 B.n684 VSUBS 0.009828f
C725 B.n685 VSUBS 0.009828f
C726 B.n686 VSUBS 0.009828f
C727 B.n687 VSUBS 0.009828f
C728 B.n688 VSUBS 0.009828f
C729 B.n689 VSUBS 0.009828f
C730 B.n690 VSUBS 0.009828f
C731 B.n691 VSUBS 0.009828f
C732 B.n692 VSUBS 0.009828f
C733 B.n693 VSUBS 0.009828f
C734 B.n694 VSUBS 0.009828f
C735 B.n695 VSUBS 0.009828f
C736 B.n696 VSUBS 0.009828f
C737 B.n697 VSUBS 0.009828f
C738 B.n698 VSUBS 0.009828f
C739 B.n699 VSUBS 0.009828f
C740 B.n700 VSUBS 0.009828f
C741 B.n701 VSUBS 0.009828f
C742 B.n702 VSUBS 0.009828f
C743 B.n703 VSUBS 0.009828f
C744 B.n704 VSUBS 0.009828f
C745 B.n705 VSUBS 0.009828f
C746 B.n706 VSUBS 0.009828f
C747 B.n707 VSUBS 0.009828f
C748 B.n708 VSUBS 0.009828f
C749 B.n709 VSUBS 0.009828f
C750 B.n710 VSUBS 0.009828f
C751 B.n711 VSUBS 0.009828f
C752 B.n712 VSUBS 0.009828f
C753 B.n713 VSUBS 0.009828f
C754 B.n714 VSUBS 0.009828f
C755 B.n715 VSUBS 0.009828f
C756 B.n716 VSUBS 0.009828f
C757 B.n717 VSUBS 0.009828f
C758 B.n718 VSUBS 0.009828f
C759 B.n719 VSUBS 0.009828f
C760 B.n720 VSUBS 0.009828f
C761 B.n721 VSUBS 0.009828f
C762 B.n722 VSUBS 0.009828f
C763 B.n723 VSUBS 0.009828f
C764 B.n724 VSUBS 0.009828f
C765 B.n725 VSUBS 0.009828f
C766 B.n726 VSUBS 0.009828f
C767 B.n727 VSUBS 0.009828f
C768 B.n728 VSUBS 0.009828f
C769 B.n729 VSUBS 0.009828f
C770 B.n730 VSUBS 0.009828f
C771 B.n731 VSUBS 0.009828f
C772 B.n732 VSUBS 0.009828f
C773 B.n733 VSUBS 0.009828f
C774 B.n734 VSUBS 0.009828f
C775 B.n735 VSUBS 0.009828f
C776 B.n736 VSUBS 0.009828f
C777 B.n737 VSUBS 0.009828f
C778 B.n738 VSUBS 0.009828f
C779 B.n739 VSUBS 0.009828f
C780 B.n740 VSUBS 0.009828f
C781 B.n741 VSUBS 0.009828f
C782 B.n742 VSUBS 0.009828f
C783 B.n743 VSUBS 0.009828f
C784 B.n744 VSUBS 0.009828f
C785 B.n745 VSUBS 0.009828f
C786 B.n746 VSUBS 0.009828f
C787 B.n747 VSUBS 0.023807f
C788 B.n748 VSUBS 0.023807f
C789 B.n749 VSUBS 0.024465f
C790 B.n750 VSUBS 0.009828f
C791 B.n751 VSUBS 0.009828f
C792 B.n752 VSUBS 0.009828f
C793 B.n753 VSUBS 0.009828f
C794 B.n754 VSUBS 0.009828f
C795 B.n755 VSUBS 0.009828f
C796 B.n756 VSUBS 0.009828f
C797 B.n757 VSUBS 0.009828f
C798 B.n758 VSUBS 0.009828f
C799 B.n759 VSUBS 0.009828f
C800 B.n760 VSUBS 0.009828f
C801 B.n761 VSUBS 0.009828f
C802 B.n762 VSUBS 0.009828f
C803 B.n763 VSUBS 0.009828f
C804 B.n764 VSUBS 0.009828f
C805 B.n765 VSUBS 0.009828f
C806 B.n766 VSUBS 0.009828f
C807 B.n767 VSUBS 0.009828f
C808 B.n768 VSUBS 0.009828f
C809 B.n769 VSUBS 0.009828f
C810 B.n770 VSUBS 0.009828f
C811 B.n771 VSUBS 0.009828f
C812 B.n772 VSUBS 0.009828f
C813 B.n773 VSUBS 0.009828f
C814 B.n774 VSUBS 0.009828f
C815 B.n775 VSUBS 0.009828f
C816 B.n776 VSUBS 0.009828f
C817 B.n777 VSUBS 0.009828f
C818 B.n778 VSUBS 0.009828f
C819 B.n779 VSUBS 0.009828f
C820 B.n780 VSUBS 0.009828f
C821 B.n781 VSUBS 0.009828f
C822 B.n782 VSUBS 0.009828f
C823 B.n783 VSUBS 0.009828f
C824 B.n784 VSUBS 0.009828f
C825 B.n785 VSUBS 0.009828f
C826 B.n786 VSUBS 0.009828f
C827 B.n787 VSUBS 0.009828f
C828 B.n788 VSUBS 0.009828f
C829 B.n789 VSUBS 0.009828f
C830 B.n790 VSUBS 0.009828f
C831 B.n791 VSUBS 0.009828f
C832 B.n792 VSUBS 0.009828f
C833 B.n793 VSUBS 0.009828f
C834 B.n794 VSUBS 0.009828f
C835 B.n795 VSUBS 0.009828f
C836 B.n796 VSUBS 0.009828f
C837 B.n797 VSUBS 0.006793f
C838 B.n798 VSUBS 0.02277f
C839 B.n799 VSUBS 0.007949f
C840 B.n800 VSUBS 0.009828f
C841 B.n801 VSUBS 0.009828f
C842 B.n802 VSUBS 0.009828f
C843 B.n803 VSUBS 0.009828f
C844 B.n804 VSUBS 0.009828f
C845 B.n805 VSUBS 0.009828f
C846 B.n806 VSUBS 0.009828f
C847 B.n807 VSUBS 0.009828f
C848 B.n808 VSUBS 0.009828f
C849 B.n809 VSUBS 0.009828f
C850 B.n810 VSUBS 0.009828f
C851 B.n811 VSUBS 0.007949f
C852 B.n812 VSUBS 0.009828f
C853 B.n813 VSUBS 0.009828f
C854 B.n814 VSUBS 0.009828f
C855 B.n815 VSUBS 0.009828f
C856 B.n816 VSUBS 0.009828f
C857 B.n817 VSUBS 0.009828f
C858 B.n818 VSUBS 0.009828f
C859 B.n819 VSUBS 0.009828f
C860 B.n820 VSUBS 0.009828f
C861 B.n821 VSUBS 0.009828f
C862 B.n822 VSUBS 0.009828f
C863 B.n823 VSUBS 0.009828f
C864 B.n824 VSUBS 0.009828f
C865 B.n825 VSUBS 0.009828f
C866 B.n826 VSUBS 0.009828f
C867 B.n827 VSUBS 0.009828f
C868 B.n828 VSUBS 0.009828f
C869 B.n829 VSUBS 0.009828f
C870 B.n830 VSUBS 0.009828f
C871 B.n831 VSUBS 0.009828f
C872 B.n832 VSUBS 0.009828f
C873 B.n833 VSUBS 0.009828f
C874 B.n834 VSUBS 0.009828f
C875 B.n835 VSUBS 0.009828f
C876 B.n836 VSUBS 0.009828f
C877 B.n837 VSUBS 0.009828f
C878 B.n838 VSUBS 0.009828f
C879 B.n839 VSUBS 0.009828f
C880 B.n840 VSUBS 0.009828f
C881 B.n841 VSUBS 0.009828f
C882 B.n842 VSUBS 0.009828f
C883 B.n843 VSUBS 0.009828f
C884 B.n844 VSUBS 0.009828f
C885 B.n845 VSUBS 0.009828f
C886 B.n846 VSUBS 0.009828f
C887 B.n847 VSUBS 0.009828f
C888 B.n848 VSUBS 0.009828f
C889 B.n849 VSUBS 0.009828f
C890 B.n850 VSUBS 0.009828f
C891 B.n851 VSUBS 0.009828f
C892 B.n852 VSUBS 0.009828f
C893 B.n853 VSUBS 0.009828f
C894 B.n854 VSUBS 0.009828f
C895 B.n855 VSUBS 0.009828f
C896 B.n856 VSUBS 0.009828f
C897 B.n857 VSUBS 0.009828f
C898 B.n858 VSUBS 0.009828f
C899 B.n859 VSUBS 0.009828f
C900 B.n860 VSUBS 0.009828f
C901 B.n861 VSUBS 0.024465f
C902 B.n862 VSUBS 0.023807f
C903 B.n863 VSUBS 0.023807f
C904 B.n864 VSUBS 0.009828f
C905 B.n865 VSUBS 0.009828f
C906 B.n866 VSUBS 0.009828f
C907 B.n867 VSUBS 0.009828f
C908 B.n868 VSUBS 0.009828f
C909 B.n869 VSUBS 0.009828f
C910 B.n870 VSUBS 0.009828f
C911 B.n871 VSUBS 0.009828f
C912 B.n872 VSUBS 0.009828f
C913 B.n873 VSUBS 0.009828f
C914 B.n874 VSUBS 0.009828f
C915 B.n875 VSUBS 0.009828f
C916 B.n876 VSUBS 0.009828f
C917 B.n877 VSUBS 0.009828f
C918 B.n878 VSUBS 0.009828f
C919 B.n879 VSUBS 0.009828f
C920 B.n880 VSUBS 0.009828f
C921 B.n881 VSUBS 0.009828f
C922 B.n882 VSUBS 0.009828f
C923 B.n883 VSUBS 0.009828f
C924 B.n884 VSUBS 0.009828f
C925 B.n885 VSUBS 0.009828f
C926 B.n886 VSUBS 0.009828f
C927 B.n887 VSUBS 0.009828f
C928 B.n888 VSUBS 0.009828f
C929 B.n889 VSUBS 0.009828f
C930 B.n890 VSUBS 0.009828f
C931 B.n891 VSUBS 0.009828f
C932 B.n892 VSUBS 0.009828f
C933 B.n893 VSUBS 0.009828f
C934 B.n894 VSUBS 0.009828f
C935 B.n895 VSUBS 0.009828f
C936 B.n896 VSUBS 0.009828f
C937 B.n897 VSUBS 0.009828f
C938 B.n898 VSUBS 0.009828f
C939 B.n899 VSUBS 0.009828f
C940 B.n900 VSUBS 0.009828f
C941 B.n901 VSUBS 0.009828f
C942 B.n902 VSUBS 0.009828f
C943 B.n903 VSUBS 0.009828f
C944 B.n904 VSUBS 0.009828f
C945 B.n905 VSUBS 0.009828f
C946 B.n906 VSUBS 0.009828f
C947 B.n907 VSUBS 0.009828f
C948 B.n908 VSUBS 0.009828f
C949 B.n909 VSUBS 0.009828f
C950 B.n910 VSUBS 0.009828f
C951 B.n911 VSUBS 0.009828f
C952 B.n912 VSUBS 0.009828f
C953 B.n913 VSUBS 0.009828f
C954 B.n914 VSUBS 0.009828f
C955 B.n915 VSUBS 0.009828f
C956 B.n916 VSUBS 0.009828f
C957 B.n917 VSUBS 0.009828f
C958 B.n918 VSUBS 0.009828f
C959 B.n919 VSUBS 0.009828f
C960 B.n920 VSUBS 0.009828f
C961 B.n921 VSUBS 0.009828f
C962 B.n922 VSUBS 0.009828f
C963 B.n923 VSUBS 0.009828f
C964 B.n924 VSUBS 0.009828f
C965 B.n925 VSUBS 0.009828f
C966 B.n926 VSUBS 0.009828f
C967 B.n927 VSUBS 0.009828f
C968 B.n928 VSUBS 0.009828f
C969 B.n929 VSUBS 0.009828f
C970 B.n930 VSUBS 0.009828f
C971 B.n931 VSUBS 0.009828f
C972 B.n932 VSUBS 0.009828f
C973 B.n933 VSUBS 0.009828f
C974 B.n934 VSUBS 0.009828f
C975 B.n935 VSUBS 0.009828f
C976 B.n936 VSUBS 0.009828f
C977 B.n937 VSUBS 0.009828f
C978 B.n938 VSUBS 0.009828f
C979 B.n939 VSUBS 0.009828f
C980 B.n940 VSUBS 0.009828f
C981 B.n941 VSUBS 0.009828f
C982 B.n942 VSUBS 0.009828f
C983 B.n943 VSUBS 0.009828f
C984 B.n944 VSUBS 0.009828f
C985 B.n945 VSUBS 0.009828f
C986 B.n946 VSUBS 0.009828f
C987 B.n947 VSUBS 0.009828f
C988 B.n948 VSUBS 0.009828f
C989 B.n949 VSUBS 0.009828f
C990 B.n950 VSUBS 0.009828f
C991 B.n951 VSUBS 0.009828f
C992 B.n952 VSUBS 0.009828f
C993 B.n953 VSUBS 0.009828f
C994 B.n954 VSUBS 0.009828f
C995 B.n955 VSUBS 0.009828f
C996 B.n956 VSUBS 0.009828f
C997 B.n957 VSUBS 0.009828f
C998 B.n958 VSUBS 0.009828f
C999 B.n959 VSUBS 0.009828f
C1000 B.n960 VSUBS 0.009828f
C1001 B.n961 VSUBS 0.009828f
C1002 B.n962 VSUBS 0.009828f
C1003 B.n963 VSUBS 0.009828f
C1004 B.n964 VSUBS 0.009828f
C1005 B.n965 VSUBS 0.009828f
C1006 B.n966 VSUBS 0.009828f
C1007 B.n967 VSUBS 0.009828f
C1008 B.n968 VSUBS 0.009828f
C1009 B.n969 VSUBS 0.009828f
C1010 B.n970 VSUBS 0.009828f
C1011 B.n971 VSUBS 0.009828f
C1012 B.n972 VSUBS 0.009828f
C1013 B.n973 VSUBS 0.009828f
C1014 B.n974 VSUBS 0.009828f
C1015 B.n975 VSUBS 0.009828f
C1016 B.n976 VSUBS 0.009828f
C1017 B.n977 VSUBS 0.009828f
C1018 B.n978 VSUBS 0.009828f
C1019 B.n979 VSUBS 0.009828f
C1020 B.n980 VSUBS 0.009828f
C1021 B.n981 VSUBS 0.009828f
C1022 B.n982 VSUBS 0.009828f
C1023 B.n983 VSUBS 0.009828f
C1024 B.n984 VSUBS 0.009828f
C1025 B.n985 VSUBS 0.009828f
C1026 B.n986 VSUBS 0.009828f
C1027 B.n987 VSUBS 0.012825f
C1028 B.n988 VSUBS 0.013662f
C1029 B.n989 VSUBS 0.027168f
C1030 VDD1.t3 VSUBS 2.36529f
C1031 VDD1.t5 VSUBS 0.236948f
C1032 VDD1.t9 VSUBS 0.236948f
C1033 VDD1.n0 VSUBS 1.76493f
C1034 VDD1.n1 VSUBS 2.11f
C1035 VDD1.t7 VSUBS 2.36528f
C1036 VDD1.t1 VSUBS 0.236948f
C1037 VDD1.t2 VSUBS 0.236948f
C1038 VDD1.n2 VSUBS 1.76493f
C1039 VDD1.n3 VSUBS 2.09877f
C1040 VDD1.t8 VSUBS 0.236948f
C1041 VDD1.t0 VSUBS 0.236948f
C1042 VDD1.n4 VSUBS 1.80601f
C1043 VDD1.n5 VSUBS 5.08642f
C1044 VDD1.t6 VSUBS 0.236948f
C1045 VDD1.t4 VSUBS 0.236948f
C1046 VDD1.n6 VSUBS 1.76493f
C1047 VDD1.n7 VSUBS 4.97935f
C1048 VP.n0 VSUBS 0.052331f
C1049 VP.t9 VSUBS 2.71844f
C1050 VP.n1 VSUBS 0.051851f
C1051 VP.n2 VSUBS 0.027821f
C1052 VP.n3 VSUBS 0.051851f
C1053 VP.n4 VSUBS 0.027821f
C1054 VP.t1 VSUBS 2.71844f
C1055 VP.n5 VSUBS 0.051851f
C1056 VP.n6 VSUBS 0.027821f
C1057 VP.n7 VSUBS 0.051851f
C1058 VP.n8 VSUBS 0.027821f
C1059 VP.t7 VSUBS 2.71844f
C1060 VP.n9 VSUBS 0.051851f
C1061 VP.n10 VSUBS 0.027821f
C1062 VP.n11 VSUBS 0.056047f
C1063 VP.n12 VSUBS 0.027821f
C1064 VP.t8 VSUBS 2.71844f
C1065 VP.n13 VSUBS 0.966398f
C1066 VP.n14 VSUBS 0.027821f
C1067 VP.n15 VSUBS 0.040228f
C1068 VP.n16 VSUBS 0.027821f
C1069 VP.n17 VSUBS 0.047243f
C1070 VP.n18 VSUBS 0.052331f
C1071 VP.t5 VSUBS 2.71844f
C1072 VP.n19 VSUBS 0.051851f
C1073 VP.n20 VSUBS 0.027821f
C1074 VP.n21 VSUBS 0.051851f
C1075 VP.n22 VSUBS 0.027821f
C1076 VP.t3 VSUBS 2.71844f
C1077 VP.n23 VSUBS 0.051851f
C1078 VP.n24 VSUBS 0.027821f
C1079 VP.n25 VSUBS 0.051851f
C1080 VP.n26 VSUBS 0.027821f
C1081 VP.t0 VSUBS 2.71844f
C1082 VP.n27 VSUBS 0.051851f
C1083 VP.n28 VSUBS 0.027821f
C1084 VP.n29 VSUBS 0.056047f
C1085 VP.n30 VSUBS 0.027821f
C1086 VP.t4 VSUBS 2.71844f
C1087 VP.n31 VSUBS 1.06006f
C1088 VP.t6 VSUBS 3.15964f
C1089 VP.n32 VSUBS 1.01282f
C1090 VP.n33 VSUBS 0.372309f
C1091 VP.n34 VSUBS 0.030348f
C1092 VP.n35 VSUBS 0.051851f
C1093 VP.n36 VSUBS 0.051851f
C1094 VP.n37 VSUBS 0.027821f
C1095 VP.n38 VSUBS 0.027821f
C1096 VP.n39 VSUBS 0.027821f
C1097 VP.n40 VSUBS 0.025185f
C1098 VP.n41 VSUBS 0.051851f
C1099 VP.n42 VSUBS 0.051851f
C1100 VP.n43 VSUBS 0.027821f
C1101 VP.n44 VSUBS 0.027821f
C1102 VP.n45 VSUBS 0.027821f
C1103 VP.n46 VSUBS 0.039051f
C1104 VP.n47 VSUBS 0.966398f
C1105 VP.n48 VSUBS 0.039051f
C1106 VP.n49 VSUBS 0.051851f
C1107 VP.n50 VSUBS 0.027821f
C1108 VP.n51 VSUBS 0.027821f
C1109 VP.n52 VSUBS 0.027821f
C1110 VP.n53 VSUBS 0.051851f
C1111 VP.n54 VSUBS 0.025185f
C1112 VP.n55 VSUBS 0.056047f
C1113 VP.n56 VSUBS 0.027821f
C1114 VP.n57 VSUBS 0.027821f
C1115 VP.n58 VSUBS 0.027821f
C1116 VP.n59 VSUBS 0.051851f
C1117 VP.n60 VSUBS 0.030348f
C1118 VP.n61 VSUBS 0.966398f
C1119 VP.n62 VSUBS 0.047755f
C1120 VP.n63 VSUBS 0.027821f
C1121 VP.n64 VSUBS 0.027821f
C1122 VP.n65 VSUBS 0.027821f
C1123 VP.n66 VSUBS 0.051851f
C1124 VP.n67 VSUBS 0.040228f
C1125 VP.n68 VSUBS 0.041004f
C1126 VP.n69 VSUBS 0.027821f
C1127 VP.n70 VSUBS 0.027821f
C1128 VP.n71 VSUBS 0.027821f
C1129 VP.n72 VSUBS 0.051851f
C1130 VP.n73 VSUBS 0.047243f
C1131 VP.n74 VSUBS 1.08873f
C1132 VP.n75 VSUBS 2.01794f
C1133 VP.t2 VSUBS 2.71844f
C1134 VP.n76 VSUBS 1.08873f
C1135 VP.n77 VSUBS 2.03497f
C1136 VP.n78 VSUBS 0.052331f
C1137 VP.n79 VSUBS 0.027821f
C1138 VP.n80 VSUBS 0.051851f
C1139 VP.n81 VSUBS 0.051851f
C1140 VP.n82 VSUBS 0.041004f
C1141 VP.n83 VSUBS 0.027821f
C1142 VP.n84 VSUBS 0.027821f
C1143 VP.n85 VSUBS 0.027821f
C1144 VP.n86 VSUBS 0.051851f
C1145 VP.n87 VSUBS 0.051851f
C1146 VP.n88 VSUBS 0.047755f
C1147 VP.n89 VSUBS 0.027821f
C1148 VP.n90 VSUBS 0.027821f
C1149 VP.n91 VSUBS 0.030348f
C1150 VP.n92 VSUBS 0.051851f
C1151 VP.n93 VSUBS 0.051851f
C1152 VP.n94 VSUBS 0.027821f
C1153 VP.n95 VSUBS 0.027821f
C1154 VP.n96 VSUBS 0.027821f
C1155 VP.n97 VSUBS 0.025185f
C1156 VP.n98 VSUBS 0.051851f
C1157 VP.n99 VSUBS 0.051851f
C1158 VP.n100 VSUBS 0.027821f
C1159 VP.n101 VSUBS 0.027821f
C1160 VP.n102 VSUBS 0.027821f
C1161 VP.n103 VSUBS 0.039051f
C1162 VP.n104 VSUBS 0.966398f
C1163 VP.n105 VSUBS 0.039051f
C1164 VP.n106 VSUBS 0.051851f
C1165 VP.n107 VSUBS 0.027821f
C1166 VP.n108 VSUBS 0.027821f
C1167 VP.n109 VSUBS 0.027821f
C1168 VP.n110 VSUBS 0.051851f
C1169 VP.n111 VSUBS 0.025185f
C1170 VP.n112 VSUBS 0.056047f
C1171 VP.n113 VSUBS 0.027821f
C1172 VP.n114 VSUBS 0.027821f
C1173 VP.n115 VSUBS 0.027821f
C1174 VP.n116 VSUBS 0.051851f
C1175 VP.n117 VSUBS 0.030348f
C1176 VP.n118 VSUBS 0.966398f
C1177 VP.n119 VSUBS 0.047755f
C1178 VP.n120 VSUBS 0.027821f
C1179 VP.n121 VSUBS 0.027821f
C1180 VP.n122 VSUBS 0.027821f
C1181 VP.n123 VSUBS 0.051851f
C1182 VP.n124 VSUBS 0.040228f
C1183 VP.n125 VSUBS 0.041004f
C1184 VP.n126 VSUBS 0.027821f
C1185 VP.n127 VSUBS 0.027821f
C1186 VP.n128 VSUBS 0.027821f
C1187 VP.n129 VSUBS 0.051851f
C1188 VP.n130 VSUBS 0.047243f
C1189 VP.n131 VSUBS 1.08873f
C1190 VP.n132 VSUBS 0.089294f
C1191 VDD2.t4 VSUBS 2.36716f
C1192 VDD2.t1 VSUBS 0.237135f
C1193 VDD2.t5 VSUBS 0.237135f
C1194 VDD2.n0 VSUBS 1.76633f
C1195 VDD2.n1 VSUBS 2.10043f
C1196 VDD2.t2 VSUBS 0.237135f
C1197 VDD2.t3 VSUBS 0.237135f
C1198 VDD2.n2 VSUBS 1.80744f
C1199 VDD2.n3 VSUBS 4.87652f
C1200 VDD2.t7 VSUBS 2.3225f
C1201 VDD2.n4 VSUBS 4.87241f
C1202 VDD2.t8 VSUBS 0.237135f
C1203 VDD2.t9 VSUBS 0.237135f
C1204 VDD2.n5 VSUBS 1.76633f
C1205 VDD2.n6 VSUBS 1.07917f
C1206 VDD2.t0 VSUBS 0.237135f
C1207 VDD2.t6 VSUBS 0.237135f
C1208 VDD2.n7 VSUBS 1.80737f
C1209 VTAIL.t17 VSUBS 0.228212f
C1210 VTAIL.t13 VSUBS 0.228212f
C1211 VTAIL.n0 VSUBS 1.56174f
C1212 VTAIL.n1 VSUBS 1.18162f
C1213 VTAIL.t8 VSUBS 2.08322f
C1214 VTAIL.n2 VSUBS 1.3725f
C1215 VTAIL.t4 VSUBS 0.228212f
C1216 VTAIL.t2 VSUBS 0.228212f
C1217 VTAIL.n3 VSUBS 1.56174f
C1218 VTAIL.n4 VSUBS 1.41518f
C1219 VTAIL.t5 VSUBS 0.228212f
C1220 VTAIL.t6 VSUBS 0.228212f
C1221 VTAIL.n5 VSUBS 1.56174f
C1222 VTAIL.n6 VSUBS 3.03467f
C1223 VTAIL.t11 VSUBS 0.228212f
C1224 VTAIL.t18 VSUBS 0.228212f
C1225 VTAIL.n7 VSUBS 1.56175f
C1226 VTAIL.n8 VSUBS 3.03466f
C1227 VTAIL.t10 VSUBS 0.228212f
C1228 VTAIL.t15 VSUBS 0.228212f
C1229 VTAIL.n9 VSUBS 1.56175f
C1230 VTAIL.n10 VSUBS 1.41518f
C1231 VTAIL.t16 VSUBS 2.08323f
C1232 VTAIL.n11 VSUBS 1.37249f
C1233 VTAIL.t3 VSUBS 0.228212f
C1234 VTAIL.t0 VSUBS 0.228212f
C1235 VTAIL.n12 VSUBS 1.56175f
C1236 VTAIL.n13 VSUBS 1.27158f
C1237 VTAIL.t19 VSUBS 0.228212f
C1238 VTAIL.t7 VSUBS 0.228212f
C1239 VTAIL.n14 VSUBS 1.56175f
C1240 VTAIL.n15 VSUBS 1.41518f
C1241 VTAIL.t1 VSUBS 2.08322f
C1242 VTAIL.n16 VSUBS 2.75177f
C1243 VTAIL.t9 VSUBS 2.08322f
C1244 VTAIL.n17 VSUBS 2.75177f
C1245 VTAIL.t14 VSUBS 0.228212f
C1246 VTAIL.t12 VSUBS 0.228212f
C1247 VTAIL.n18 VSUBS 1.56174f
C1248 VTAIL.n19 VSUBS 1.12134f
C1249 VN.n0 VSUBS 0.047382f
C1250 VN.t6 VSUBS 2.46135f
C1251 VN.n1 VSUBS 0.046947f
C1252 VN.n2 VSUBS 0.02519f
C1253 VN.n3 VSUBS 0.046947f
C1254 VN.n4 VSUBS 0.02519f
C1255 VN.t7 VSUBS 2.46135f
C1256 VN.n5 VSUBS 0.046947f
C1257 VN.n6 VSUBS 0.02519f
C1258 VN.n7 VSUBS 0.046947f
C1259 VN.n8 VSUBS 0.02519f
C1260 VN.t4 VSUBS 2.46135f
C1261 VN.n9 VSUBS 0.046947f
C1262 VN.n10 VSUBS 0.02519f
C1263 VN.n11 VSUBS 0.050746f
C1264 VN.n12 VSUBS 0.02519f
C1265 VN.t8 VSUBS 2.46135f
C1266 VN.n13 VSUBS 0.959808f
C1267 VN.t5 VSUBS 2.86083f
C1268 VN.n14 VSUBS 0.917029f
C1269 VN.n15 VSUBS 0.337098f
C1270 VN.n16 VSUBS 0.027478f
C1271 VN.n17 VSUBS 0.046947f
C1272 VN.n18 VSUBS 0.046947f
C1273 VN.n19 VSUBS 0.02519f
C1274 VN.n20 VSUBS 0.02519f
C1275 VN.n21 VSUBS 0.02519f
C1276 VN.n22 VSUBS 0.022803f
C1277 VN.n23 VSUBS 0.046947f
C1278 VN.n24 VSUBS 0.046947f
C1279 VN.n25 VSUBS 0.02519f
C1280 VN.n26 VSUBS 0.02519f
C1281 VN.n27 VSUBS 0.02519f
C1282 VN.n28 VSUBS 0.035358f
C1283 VN.n29 VSUBS 0.875004f
C1284 VN.n30 VSUBS 0.035358f
C1285 VN.n31 VSUBS 0.046947f
C1286 VN.n32 VSUBS 0.02519f
C1287 VN.n33 VSUBS 0.02519f
C1288 VN.n34 VSUBS 0.02519f
C1289 VN.n35 VSUBS 0.046947f
C1290 VN.n36 VSUBS 0.022803f
C1291 VN.n37 VSUBS 0.050746f
C1292 VN.n38 VSUBS 0.02519f
C1293 VN.n39 VSUBS 0.02519f
C1294 VN.n40 VSUBS 0.02519f
C1295 VN.n41 VSUBS 0.046947f
C1296 VN.n42 VSUBS 0.027478f
C1297 VN.n43 VSUBS 0.875004f
C1298 VN.n44 VSUBS 0.043239f
C1299 VN.n45 VSUBS 0.02519f
C1300 VN.n46 VSUBS 0.02519f
C1301 VN.n47 VSUBS 0.02519f
C1302 VN.n48 VSUBS 0.046947f
C1303 VN.n49 VSUBS 0.036424f
C1304 VN.n50 VSUBS 0.037126f
C1305 VN.n51 VSUBS 0.02519f
C1306 VN.n52 VSUBS 0.02519f
C1307 VN.n53 VSUBS 0.02519f
C1308 VN.n54 VSUBS 0.046947f
C1309 VN.n55 VSUBS 0.042775f
C1310 VN.n56 VSUBS 0.985767f
C1311 VN.n57 VSUBS 0.080849f
C1312 VN.n58 VSUBS 0.047382f
C1313 VN.t2 VSUBS 2.46135f
C1314 VN.n59 VSUBS 0.046947f
C1315 VN.n60 VSUBS 0.02519f
C1316 VN.n61 VSUBS 0.046947f
C1317 VN.n62 VSUBS 0.02519f
C1318 VN.t1 VSUBS 2.46135f
C1319 VN.n63 VSUBS 0.046947f
C1320 VN.n64 VSUBS 0.02519f
C1321 VN.n65 VSUBS 0.046947f
C1322 VN.n66 VSUBS 0.02519f
C1323 VN.t0 VSUBS 2.46135f
C1324 VN.n67 VSUBS 0.046947f
C1325 VN.n68 VSUBS 0.02519f
C1326 VN.n69 VSUBS 0.050746f
C1327 VN.n70 VSUBS 0.02519f
C1328 VN.t9 VSUBS 2.46135f
C1329 VN.n71 VSUBS 0.959808f
C1330 VN.t3 VSUBS 2.86083f
C1331 VN.n72 VSUBS 0.917029f
C1332 VN.n73 VSUBS 0.337098f
C1333 VN.n74 VSUBS 0.027478f
C1334 VN.n75 VSUBS 0.046947f
C1335 VN.n76 VSUBS 0.046947f
C1336 VN.n77 VSUBS 0.02519f
C1337 VN.n78 VSUBS 0.02519f
C1338 VN.n79 VSUBS 0.02519f
C1339 VN.n80 VSUBS 0.022803f
C1340 VN.n81 VSUBS 0.046947f
C1341 VN.n82 VSUBS 0.046947f
C1342 VN.n83 VSUBS 0.02519f
C1343 VN.n84 VSUBS 0.02519f
C1344 VN.n85 VSUBS 0.02519f
C1345 VN.n86 VSUBS 0.035358f
C1346 VN.n87 VSUBS 0.875004f
C1347 VN.n88 VSUBS 0.035358f
C1348 VN.n89 VSUBS 0.046947f
C1349 VN.n90 VSUBS 0.02519f
C1350 VN.n91 VSUBS 0.02519f
C1351 VN.n92 VSUBS 0.02519f
C1352 VN.n93 VSUBS 0.046947f
C1353 VN.n94 VSUBS 0.022803f
C1354 VN.n95 VSUBS 0.050746f
C1355 VN.n96 VSUBS 0.02519f
C1356 VN.n97 VSUBS 0.02519f
C1357 VN.n98 VSUBS 0.02519f
C1358 VN.n99 VSUBS 0.046947f
C1359 VN.n100 VSUBS 0.027478f
C1360 VN.n101 VSUBS 0.875004f
C1361 VN.n102 VSUBS 0.043239f
C1362 VN.n103 VSUBS 0.02519f
C1363 VN.n104 VSUBS 0.02519f
C1364 VN.n105 VSUBS 0.02519f
C1365 VN.n106 VSUBS 0.046947f
C1366 VN.n107 VSUBS 0.036424f
C1367 VN.n108 VSUBS 0.037126f
C1368 VN.n109 VSUBS 0.02519f
C1369 VN.n110 VSUBS 0.02519f
C1370 VN.n111 VSUBS 0.02519f
C1371 VN.n112 VSUBS 0.046947f
C1372 VN.n113 VSUBS 0.042775f
C1373 VN.n114 VSUBS 0.985767f
C1374 VN.n115 VSUBS 1.83294f
.ends

