* NGSPICE file created from diff_pair_sample_1744.ext - technology: sky130A

.subckt diff_pair_sample_1744 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=2.7225 ps=16.83 w=16.5 l=1.18
X1 B.t11 B.t9 B.t10 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=0 ps=0 w=16.5 l=1.18
X2 VTAIL.t6 VP.t1 VDD1.t4 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=2.7225 ps=16.83 w=16.5 l=1.18
X3 B.t8 B.t6 B.t7 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=0 ps=0 w=16.5 l=1.18
X4 VDD1.t3 VP.t2 VTAIL.t7 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=2.7225 ps=16.83 w=16.5 l=1.18
X5 VDD2.t5 VN.t0 VTAIL.t1 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=2.7225 ps=16.83 w=16.5 l=1.18
X6 VDD2.t4 VN.t1 VTAIL.t2 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=6.435 ps=33.78 w=16.5 l=1.18
X7 B.t5 B.t3 B.t4 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=0 ps=0 w=16.5 l=1.18
X8 VTAIL.t8 VP.t3 VDD1.t2 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=2.7225 ps=16.83 w=16.5 l=1.18
X9 VDD2.t3 VN.t2 VTAIL.t4 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=2.7225 ps=16.83 w=16.5 l=1.18
X10 VDD2.t2 VN.t3 VTAIL.t5 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=6.435 ps=33.78 w=16.5 l=1.18
X11 VTAIL.t3 VN.t4 VDD2.t1 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=2.7225 ps=16.83 w=16.5 l=1.18
X12 VDD1.t1 VP.t4 VTAIL.t11 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=6.435 ps=33.78 w=16.5 l=1.18
X13 VTAIL.t0 VN.t5 VDD2.t0 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=2.7225 ps=16.83 w=16.5 l=1.18
X14 B.t2 B.t0 B.t1 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=6.435 pd=33.78 as=0 ps=0 w=16.5 l=1.18
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n2178_n4268# sky130_fd_pr__pfet_01v8 ad=2.7225 pd=16.83 as=6.435 ps=33.78 w=16.5 l=1.18
R0 VP.n7 VP.t0 367.483
R1 VP.n3 VP.t2 336.993
R2 VP.n18 VP.t1 336.993
R3 VP.n25 VP.t5 336.993
R4 VP.n12 VP.t4 336.993
R5 VP.n6 VP.t3 336.993
R6 VP.n14 VP.n3 173.105
R7 VP.n26 VP.n25 173.105
R8 VP.n13 VP.n12 173.105
R9 VP.n8 VP.n5 161.3
R10 VP.n10 VP.n9 161.3
R11 VP.n11 VP.n4 161.3
R12 VP.n24 VP.n0 161.3
R13 VP.n23 VP.n22 161.3
R14 VP.n21 VP.n1 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n17 VP.n2 161.3
R17 VP.n16 VP.n15 161.3
R18 VP.n7 VP.n6 51.5093
R19 VP.n14 VP.n13 46.4058
R20 VP.n17 VP.n16 41.0614
R21 VP.n24 VP.n23 41.0614
R22 VP.n11 VP.n10 41.0614
R23 VP.n19 VP.n17 40.0926
R24 VP.n23 VP.n1 40.0926
R25 VP.n10 VP.n5 40.0926
R26 VP.n8 VP.n7 26.9198
R27 VP.n16 VP.n3 12.7883
R28 VP.n25 VP.n24 12.7883
R29 VP.n12 VP.n11 12.7883
R30 VP.n19 VP.n18 12.2964
R31 VP.n18 VP.n1 12.2964
R32 VP.n6 VP.n5 12.2964
R33 VP.n9 VP.n8 0.189894
R34 VP.n9 VP.n4 0.189894
R35 VP.n13 VP.n4 0.189894
R36 VP.n15 VP.n14 0.189894
R37 VP.n15 VP.n2 0.189894
R38 VP.n20 VP.n2 0.189894
R39 VP.n21 VP.n20 0.189894
R40 VP.n22 VP.n21 0.189894
R41 VP.n22 VP.n0 0.189894
R42 VP.n26 VP.n0 0.189894
R43 VP VP.n26 0.0516364
R44 VTAIL.n7 VTAIL.t2 56.0463
R45 VTAIL.n11 VTAIL.t5 56.0461
R46 VTAIL.n2 VTAIL.t9 56.0461
R47 VTAIL.n10 VTAIL.t11 56.0461
R48 VTAIL.n9 VTAIL.n8 54.0763
R49 VTAIL.n6 VTAIL.n5 54.0763
R50 VTAIL.n1 VTAIL.n0 54.0761
R51 VTAIL.n4 VTAIL.n3 54.0761
R52 VTAIL.n6 VTAIL.n4 29.1945
R53 VTAIL.n11 VTAIL.n10 27.8927
R54 VTAIL.n0 VTAIL.t4 1.9705
R55 VTAIL.n0 VTAIL.t3 1.9705
R56 VTAIL.n3 VTAIL.t7 1.9705
R57 VTAIL.n3 VTAIL.t6 1.9705
R58 VTAIL.n8 VTAIL.t10 1.9705
R59 VTAIL.n8 VTAIL.t8 1.9705
R60 VTAIL.n5 VTAIL.t1 1.9705
R61 VTAIL.n5 VTAIL.t0 1.9705
R62 VTAIL.n7 VTAIL.n6 1.30222
R63 VTAIL.n10 VTAIL.n9 1.30222
R64 VTAIL.n4 VTAIL.n2 1.30222
R65 VTAIL.n9 VTAIL.n7 1.12119
R66 VTAIL.n2 VTAIL.n1 1.12119
R67 VTAIL VTAIL.n11 0.918603
R68 VTAIL VTAIL.n1 0.384121
R69 VDD1 VDD1.t5 73.7596
R70 VDD1.n1 VDD1.t3 73.6458
R71 VDD1.n1 VDD1.n0 71.0249
R72 VDD1.n3 VDD1.n2 70.7549
R73 VDD1.n3 VDD1.n1 43.4039
R74 VDD1.n2 VDD1.t2 1.9705
R75 VDD1.n2 VDD1.t1 1.9705
R76 VDD1.n0 VDD1.t4 1.9705
R77 VDD1.n0 VDD1.t0 1.9705
R78 VDD1 VDD1.n3 0.267741
R79 B.n480 B.n79 585
R80 B.n482 B.n481 585
R81 B.n483 B.n78 585
R82 B.n485 B.n484 585
R83 B.n486 B.n77 585
R84 B.n488 B.n487 585
R85 B.n489 B.n76 585
R86 B.n491 B.n490 585
R87 B.n492 B.n75 585
R88 B.n494 B.n493 585
R89 B.n495 B.n74 585
R90 B.n497 B.n496 585
R91 B.n498 B.n73 585
R92 B.n500 B.n499 585
R93 B.n501 B.n72 585
R94 B.n503 B.n502 585
R95 B.n504 B.n71 585
R96 B.n506 B.n505 585
R97 B.n507 B.n70 585
R98 B.n509 B.n508 585
R99 B.n510 B.n69 585
R100 B.n512 B.n511 585
R101 B.n513 B.n68 585
R102 B.n515 B.n514 585
R103 B.n516 B.n67 585
R104 B.n518 B.n517 585
R105 B.n519 B.n66 585
R106 B.n521 B.n520 585
R107 B.n522 B.n65 585
R108 B.n524 B.n523 585
R109 B.n525 B.n64 585
R110 B.n527 B.n526 585
R111 B.n528 B.n63 585
R112 B.n530 B.n529 585
R113 B.n531 B.n62 585
R114 B.n533 B.n532 585
R115 B.n534 B.n61 585
R116 B.n536 B.n535 585
R117 B.n537 B.n60 585
R118 B.n539 B.n538 585
R119 B.n540 B.n59 585
R120 B.n542 B.n541 585
R121 B.n543 B.n58 585
R122 B.n545 B.n544 585
R123 B.n546 B.n57 585
R124 B.n548 B.n547 585
R125 B.n549 B.n56 585
R126 B.n551 B.n550 585
R127 B.n552 B.n55 585
R128 B.n554 B.n553 585
R129 B.n555 B.n54 585
R130 B.n557 B.n556 585
R131 B.n558 B.n53 585
R132 B.n560 B.n559 585
R133 B.n561 B.n50 585
R134 B.n564 B.n563 585
R135 B.n565 B.n49 585
R136 B.n567 B.n566 585
R137 B.n568 B.n48 585
R138 B.n570 B.n569 585
R139 B.n571 B.n47 585
R140 B.n573 B.n572 585
R141 B.n574 B.n43 585
R142 B.n576 B.n575 585
R143 B.n577 B.n42 585
R144 B.n579 B.n578 585
R145 B.n580 B.n41 585
R146 B.n582 B.n581 585
R147 B.n583 B.n40 585
R148 B.n585 B.n584 585
R149 B.n586 B.n39 585
R150 B.n588 B.n587 585
R151 B.n589 B.n38 585
R152 B.n591 B.n590 585
R153 B.n592 B.n37 585
R154 B.n594 B.n593 585
R155 B.n595 B.n36 585
R156 B.n597 B.n596 585
R157 B.n598 B.n35 585
R158 B.n600 B.n599 585
R159 B.n601 B.n34 585
R160 B.n603 B.n602 585
R161 B.n604 B.n33 585
R162 B.n606 B.n605 585
R163 B.n607 B.n32 585
R164 B.n609 B.n608 585
R165 B.n610 B.n31 585
R166 B.n612 B.n611 585
R167 B.n613 B.n30 585
R168 B.n615 B.n614 585
R169 B.n616 B.n29 585
R170 B.n618 B.n617 585
R171 B.n619 B.n28 585
R172 B.n621 B.n620 585
R173 B.n622 B.n27 585
R174 B.n624 B.n623 585
R175 B.n625 B.n26 585
R176 B.n627 B.n626 585
R177 B.n628 B.n25 585
R178 B.n630 B.n629 585
R179 B.n631 B.n24 585
R180 B.n633 B.n632 585
R181 B.n634 B.n23 585
R182 B.n636 B.n635 585
R183 B.n637 B.n22 585
R184 B.n639 B.n638 585
R185 B.n640 B.n21 585
R186 B.n642 B.n641 585
R187 B.n643 B.n20 585
R188 B.n645 B.n644 585
R189 B.n646 B.n19 585
R190 B.n648 B.n647 585
R191 B.n649 B.n18 585
R192 B.n651 B.n650 585
R193 B.n652 B.n17 585
R194 B.n654 B.n653 585
R195 B.n655 B.n16 585
R196 B.n657 B.n656 585
R197 B.n658 B.n15 585
R198 B.n479 B.n478 585
R199 B.n477 B.n80 585
R200 B.n476 B.n475 585
R201 B.n474 B.n81 585
R202 B.n473 B.n472 585
R203 B.n471 B.n82 585
R204 B.n470 B.n469 585
R205 B.n468 B.n83 585
R206 B.n467 B.n466 585
R207 B.n465 B.n84 585
R208 B.n464 B.n463 585
R209 B.n462 B.n85 585
R210 B.n461 B.n460 585
R211 B.n459 B.n86 585
R212 B.n458 B.n457 585
R213 B.n456 B.n87 585
R214 B.n455 B.n454 585
R215 B.n453 B.n88 585
R216 B.n452 B.n451 585
R217 B.n450 B.n89 585
R218 B.n449 B.n448 585
R219 B.n447 B.n90 585
R220 B.n446 B.n445 585
R221 B.n444 B.n91 585
R222 B.n443 B.n442 585
R223 B.n441 B.n92 585
R224 B.n440 B.n439 585
R225 B.n438 B.n93 585
R226 B.n437 B.n436 585
R227 B.n435 B.n94 585
R228 B.n434 B.n433 585
R229 B.n432 B.n95 585
R230 B.n431 B.n430 585
R231 B.n429 B.n96 585
R232 B.n428 B.n427 585
R233 B.n426 B.n97 585
R234 B.n425 B.n424 585
R235 B.n423 B.n98 585
R236 B.n422 B.n421 585
R237 B.n420 B.n99 585
R238 B.n419 B.n418 585
R239 B.n417 B.n100 585
R240 B.n416 B.n415 585
R241 B.n414 B.n101 585
R242 B.n413 B.n412 585
R243 B.n411 B.n102 585
R244 B.n410 B.n409 585
R245 B.n408 B.n103 585
R246 B.n407 B.n406 585
R247 B.n405 B.n104 585
R248 B.n404 B.n403 585
R249 B.n402 B.n105 585
R250 B.n401 B.n400 585
R251 B.n218 B.n167 585
R252 B.n220 B.n219 585
R253 B.n221 B.n166 585
R254 B.n223 B.n222 585
R255 B.n224 B.n165 585
R256 B.n226 B.n225 585
R257 B.n227 B.n164 585
R258 B.n229 B.n228 585
R259 B.n230 B.n163 585
R260 B.n232 B.n231 585
R261 B.n233 B.n162 585
R262 B.n235 B.n234 585
R263 B.n236 B.n161 585
R264 B.n238 B.n237 585
R265 B.n239 B.n160 585
R266 B.n241 B.n240 585
R267 B.n242 B.n159 585
R268 B.n244 B.n243 585
R269 B.n245 B.n158 585
R270 B.n247 B.n246 585
R271 B.n248 B.n157 585
R272 B.n250 B.n249 585
R273 B.n251 B.n156 585
R274 B.n253 B.n252 585
R275 B.n254 B.n155 585
R276 B.n256 B.n255 585
R277 B.n257 B.n154 585
R278 B.n259 B.n258 585
R279 B.n260 B.n153 585
R280 B.n262 B.n261 585
R281 B.n263 B.n152 585
R282 B.n265 B.n264 585
R283 B.n266 B.n151 585
R284 B.n268 B.n267 585
R285 B.n269 B.n150 585
R286 B.n271 B.n270 585
R287 B.n272 B.n149 585
R288 B.n274 B.n273 585
R289 B.n275 B.n148 585
R290 B.n277 B.n276 585
R291 B.n278 B.n147 585
R292 B.n280 B.n279 585
R293 B.n281 B.n146 585
R294 B.n283 B.n282 585
R295 B.n284 B.n145 585
R296 B.n286 B.n285 585
R297 B.n287 B.n144 585
R298 B.n289 B.n288 585
R299 B.n290 B.n143 585
R300 B.n292 B.n291 585
R301 B.n293 B.n142 585
R302 B.n295 B.n294 585
R303 B.n296 B.n141 585
R304 B.n298 B.n297 585
R305 B.n299 B.n138 585
R306 B.n302 B.n301 585
R307 B.n303 B.n137 585
R308 B.n305 B.n304 585
R309 B.n306 B.n136 585
R310 B.n308 B.n307 585
R311 B.n309 B.n135 585
R312 B.n311 B.n310 585
R313 B.n312 B.n134 585
R314 B.n317 B.n316 585
R315 B.n318 B.n133 585
R316 B.n320 B.n319 585
R317 B.n321 B.n132 585
R318 B.n323 B.n322 585
R319 B.n324 B.n131 585
R320 B.n326 B.n325 585
R321 B.n327 B.n130 585
R322 B.n329 B.n328 585
R323 B.n330 B.n129 585
R324 B.n332 B.n331 585
R325 B.n333 B.n128 585
R326 B.n335 B.n334 585
R327 B.n336 B.n127 585
R328 B.n338 B.n337 585
R329 B.n339 B.n126 585
R330 B.n341 B.n340 585
R331 B.n342 B.n125 585
R332 B.n344 B.n343 585
R333 B.n345 B.n124 585
R334 B.n347 B.n346 585
R335 B.n348 B.n123 585
R336 B.n350 B.n349 585
R337 B.n351 B.n122 585
R338 B.n353 B.n352 585
R339 B.n354 B.n121 585
R340 B.n356 B.n355 585
R341 B.n357 B.n120 585
R342 B.n359 B.n358 585
R343 B.n360 B.n119 585
R344 B.n362 B.n361 585
R345 B.n363 B.n118 585
R346 B.n365 B.n364 585
R347 B.n366 B.n117 585
R348 B.n368 B.n367 585
R349 B.n369 B.n116 585
R350 B.n371 B.n370 585
R351 B.n372 B.n115 585
R352 B.n374 B.n373 585
R353 B.n375 B.n114 585
R354 B.n377 B.n376 585
R355 B.n378 B.n113 585
R356 B.n380 B.n379 585
R357 B.n381 B.n112 585
R358 B.n383 B.n382 585
R359 B.n384 B.n111 585
R360 B.n386 B.n385 585
R361 B.n387 B.n110 585
R362 B.n389 B.n388 585
R363 B.n390 B.n109 585
R364 B.n392 B.n391 585
R365 B.n393 B.n108 585
R366 B.n395 B.n394 585
R367 B.n396 B.n107 585
R368 B.n398 B.n397 585
R369 B.n399 B.n106 585
R370 B.n217 B.n216 585
R371 B.n215 B.n168 585
R372 B.n214 B.n213 585
R373 B.n212 B.n169 585
R374 B.n211 B.n210 585
R375 B.n209 B.n170 585
R376 B.n208 B.n207 585
R377 B.n206 B.n171 585
R378 B.n205 B.n204 585
R379 B.n203 B.n172 585
R380 B.n202 B.n201 585
R381 B.n200 B.n173 585
R382 B.n199 B.n198 585
R383 B.n197 B.n174 585
R384 B.n196 B.n195 585
R385 B.n194 B.n175 585
R386 B.n193 B.n192 585
R387 B.n191 B.n176 585
R388 B.n190 B.n189 585
R389 B.n188 B.n177 585
R390 B.n187 B.n186 585
R391 B.n185 B.n178 585
R392 B.n184 B.n183 585
R393 B.n182 B.n179 585
R394 B.n181 B.n180 585
R395 B.n2 B.n0 585
R396 B.n697 B.n1 585
R397 B.n696 B.n695 585
R398 B.n694 B.n3 585
R399 B.n693 B.n692 585
R400 B.n691 B.n4 585
R401 B.n690 B.n689 585
R402 B.n688 B.n5 585
R403 B.n687 B.n686 585
R404 B.n685 B.n6 585
R405 B.n684 B.n683 585
R406 B.n682 B.n7 585
R407 B.n681 B.n680 585
R408 B.n679 B.n8 585
R409 B.n678 B.n677 585
R410 B.n676 B.n9 585
R411 B.n675 B.n674 585
R412 B.n673 B.n10 585
R413 B.n672 B.n671 585
R414 B.n670 B.n11 585
R415 B.n669 B.n668 585
R416 B.n667 B.n12 585
R417 B.n666 B.n665 585
R418 B.n664 B.n13 585
R419 B.n663 B.n662 585
R420 B.n661 B.n14 585
R421 B.n660 B.n659 585
R422 B.n699 B.n698 585
R423 B.n313 B.t6 541.003
R424 B.n139 B.t3 541.003
R425 B.n44 B.t9 541.003
R426 B.n51 B.t0 541.003
R427 B.n218 B.n217 502.111
R428 B.n660 B.n15 502.111
R429 B.n401 B.n106 502.111
R430 B.n480 B.n479 502.111
R431 B.n217 B.n168 163.367
R432 B.n213 B.n168 163.367
R433 B.n213 B.n212 163.367
R434 B.n212 B.n211 163.367
R435 B.n211 B.n170 163.367
R436 B.n207 B.n170 163.367
R437 B.n207 B.n206 163.367
R438 B.n206 B.n205 163.367
R439 B.n205 B.n172 163.367
R440 B.n201 B.n172 163.367
R441 B.n201 B.n200 163.367
R442 B.n200 B.n199 163.367
R443 B.n199 B.n174 163.367
R444 B.n195 B.n174 163.367
R445 B.n195 B.n194 163.367
R446 B.n194 B.n193 163.367
R447 B.n193 B.n176 163.367
R448 B.n189 B.n176 163.367
R449 B.n189 B.n188 163.367
R450 B.n188 B.n187 163.367
R451 B.n187 B.n178 163.367
R452 B.n183 B.n178 163.367
R453 B.n183 B.n182 163.367
R454 B.n182 B.n181 163.367
R455 B.n181 B.n2 163.367
R456 B.n698 B.n2 163.367
R457 B.n698 B.n697 163.367
R458 B.n697 B.n696 163.367
R459 B.n696 B.n3 163.367
R460 B.n692 B.n3 163.367
R461 B.n692 B.n691 163.367
R462 B.n691 B.n690 163.367
R463 B.n690 B.n5 163.367
R464 B.n686 B.n5 163.367
R465 B.n686 B.n685 163.367
R466 B.n685 B.n684 163.367
R467 B.n684 B.n7 163.367
R468 B.n680 B.n7 163.367
R469 B.n680 B.n679 163.367
R470 B.n679 B.n678 163.367
R471 B.n678 B.n9 163.367
R472 B.n674 B.n9 163.367
R473 B.n674 B.n673 163.367
R474 B.n673 B.n672 163.367
R475 B.n672 B.n11 163.367
R476 B.n668 B.n11 163.367
R477 B.n668 B.n667 163.367
R478 B.n667 B.n666 163.367
R479 B.n666 B.n13 163.367
R480 B.n662 B.n13 163.367
R481 B.n662 B.n661 163.367
R482 B.n661 B.n660 163.367
R483 B.n219 B.n218 163.367
R484 B.n219 B.n166 163.367
R485 B.n223 B.n166 163.367
R486 B.n224 B.n223 163.367
R487 B.n225 B.n224 163.367
R488 B.n225 B.n164 163.367
R489 B.n229 B.n164 163.367
R490 B.n230 B.n229 163.367
R491 B.n231 B.n230 163.367
R492 B.n231 B.n162 163.367
R493 B.n235 B.n162 163.367
R494 B.n236 B.n235 163.367
R495 B.n237 B.n236 163.367
R496 B.n237 B.n160 163.367
R497 B.n241 B.n160 163.367
R498 B.n242 B.n241 163.367
R499 B.n243 B.n242 163.367
R500 B.n243 B.n158 163.367
R501 B.n247 B.n158 163.367
R502 B.n248 B.n247 163.367
R503 B.n249 B.n248 163.367
R504 B.n249 B.n156 163.367
R505 B.n253 B.n156 163.367
R506 B.n254 B.n253 163.367
R507 B.n255 B.n254 163.367
R508 B.n255 B.n154 163.367
R509 B.n259 B.n154 163.367
R510 B.n260 B.n259 163.367
R511 B.n261 B.n260 163.367
R512 B.n261 B.n152 163.367
R513 B.n265 B.n152 163.367
R514 B.n266 B.n265 163.367
R515 B.n267 B.n266 163.367
R516 B.n267 B.n150 163.367
R517 B.n271 B.n150 163.367
R518 B.n272 B.n271 163.367
R519 B.n273 B.n272 163.367
R520 B.n273 B.n148 163.367
R521 B.n277 B.n148 163.367
R522 B.n278 B.n277 163.367
R523 B.n279 B.n278 163.367
R524 B.n279 B.n146 163.367
R525 B.n283 B.n146 163.367
R526 B.n284 B.n283 163.367
R527 B.n285 B.n284 163.367
R528 B.n285 B.n144 163.367
R529 B.n289 B.n144 163.367
R530 B.n290 B.n289 163.367
R531 B.n291 B.n290 163.367
R532 B.n291 B.n142 163.367
R533 B.n295 B.n142 163.367
R534 B.n296 B.n295 163.367
R535 B.n297 B.n296 163.367
R536 B.n297 B.n138 163.367
R537 B.n302 B.n138 163.367
R538 B.n303 B.n302 163.367
R539 B.n304 B.n303 163.367
R540 B.n304 B.n136 163.367
R541 B.n308 B.n136 163.367
R542 B.n309 B.n308 163.367
R543 B.n310 B.n309 163.367
R544 B.n310 B.n134 163.367
R545 B.n317 B.n134 163.367
R546 B.n318 B.n317 163.367
R547 B.n319 B.n318 163.367
R548 B.n319 B.n132 163.367
R549 B.n323 B.n132 163.367
R550 B.n324 B.n323 163.367
R551 B.n325 B.n324 163.367
R552 B.n325 B.n130 163.367
R553 B.n329 B.n130 163.367
R554 B.n330 B.n329 163.367
R555 B.n331 B.n330 163.367
R556 B.n331 B.n128 163.367
R557 B.n335 B.n128 163.367
R558 B.n336 B.n335 163.367
R559 B.n337 B.n336 163.367
R560 B.n337 B.n126 163.367
R561 B.n341 B.n126 163.367
R562 B.n342 B.n341 163.367
R563 B.n343 B.n342 163.367
R564 B.n343 B.n124 163.367
R565 B.n347 B.n124 163.367
R566 B.n348 B.n347 163.367
R567 B.n349 B.n348 163.367
R568 B.n349 B.n122 163.367
R569 B.n353 B.n122 163.367
R570 B.n354 B.n353 163.367
R571 B.n355 B.n354 163.367
R572 B.n355 B.n120 163.367
R573 B.n359 B.n120 163.367
R574 B.n360 B.n359 163.367
R575 B.n361 B.n360 163.367
R576 B.n361 B.n118 163.367
R577 B.n365 B.n118 163.367
R578 B.n366 B.n365 163.367
R579 B.n367 B.n366 163.367
R580 B.n367 B.n116 163.367
R581 B.n371 B.n116 163.367
R582 B.n372 B.n371 163.367
R583 B.n373 B.n372 163.367
R584 B.n373 B.n114 163.367
R585 B.n377 B.n114 163.367
R586 B.n378 B.n377 163.367
R587 B.n379 B.n378 163.367
R588 B.n379 B.n112 163.367
R589 B.n383 B.n112 163.367
R590 B.n384 B.n383 163.367
R591 B.n385 B.n384 163.367
R592 B.n385 B.n110 163.367
R593 B.n389 B.n110 163.367
R594 B.n390 B.n389 163.367
R595 B.n391 B.n390 163.367
R596 B.n391 B.n108 163.367
R597 B.n395 B.n108 163.367
R598 B.n396 B.n395 163.367
R599 B.n397 B.n396 163.367
R600 B.n397 B.n106 163.367
R601 B.n402 B.n401 163.367
R602 B.n403 B.n402 163.367
R603 B.n403 B.n104 163.367
R604 B.n407 B.n104 163.367
R605 B.n408 B.n407 163.367
R606 B.n409 B.n408 163.367
R607 B.n409 B.n102 163.367
R608 B.n413 B.n102 163.367
R609 B.n414 B.n413 163.367
R610 B.n415 B.n414 163.367
R611 B.n415 B.n100 163.367
R612 B.n419 B.n100 163.367
R613 B.n420 B.n419 163.367
R614 B.n421 B.n420 163.367
R615 B.n421 B.n98 163.367
R616 B.n425 B.n98 163.367
R617 B.n426 B.n425 163.367
R618 B.n427 B.n426 163.367
R619 B.n427 B.n96 163.367
R620 B.n431 B.n96 163.367
R621 B.n432 B.n431 163.367
R622 B.n433 B.n432 163.367
R623 B.n433 B.n94 163.367
R624 B.n437 B.n94 163.367
R625 B.n438 B.n437 163.367
R626 B.n439 B.n438 163.367
R627 B.n439 B.n92 163.367
R628 B.n443 B.n92 163.367
R629 B.n444 B.n443 163.367
R630 B.n445 B.n444 163.367
R631 B.n445 B.n90 163.367
R632 B.n449 B.n90 163.367
R633 B.n450 B.n449 163.367
R634 B.n451 B.n450 163.367
R635 B.n451 B.n88 163.367
R636 B.n455 B.n88 163.367
R637 B.n456 B.n455 163.367
R638 B.n457 B.n456 163.367
R639 B.n457 B.n86 163.367
R640 B.n461 B.n86 163.367
R641 B.n462 B.n461 163.367
R642 B.n463 B.n462 163.367
R643 B.n463 B.n84 163.367
R644 B.n467 B.n84 163.367
R645 B.n468 B.n467 163.367
R646 B.n469 B.n468 163.367
R647 B.n469 B.n82 163.367
R648 B.n473 B.n82 163.367
R649 B.n474 B.n473 163.367
R650 B.n475 B.n474 163.367
R651 B.n475 B.n80 163.367
R652 B.n479 B.n80 163.367
R653 B.n656 B.n15 163.367
R654 B.n656 B.n655 163.367
R655 B.n655 B.n654 163.367
R656 B.n654 B.n17 163.367
R657 B.n650 B.n17 163.367
R658 B.n650 B.n649 163.367
R659 B.n649 B.n648 163.367
R660 B.n648 B.n19 163.367
R661 B.n644 B.n19 163.367
R662 B.n644 B.n643 163.367
R663 B.n643 B.n642 163.367
R664 B.n642 B.n21 163.367
R665 B.n638 B.n21 163.367
R666 B.n638 B.n637 163.367
R667 B.n637 B.n636 163.367
R668 B.n636 B.n23 163.367
R669 B.n632 B.n23 163.367
R670 B.n632 B.n631 163.367
R671 B.n631 B.n630 163.367
R672 B.n630 B.n25 163.367
R673 B.n626 B.n25 163.367
R674 B.n626 B.n625 163.367
R675 B.n625 B.n624 163.367
R676 B.n624 B.n27 163.367
R677 B.n620 B.n27 163.367
R678 B.n620 B.n619 163.367
R679 B.n619 B.n618 163.367
R680 B.n618 B.n29 163.367
R681 B.n614 B.n29 163.367
R682 B.n614 B.n613 163.367
R683 B.n613 B.n612 163.367
R684 B.n612 B.n31 163.367
R685 B.n608 B.n31 163.367
R686 B.n608 B.n607 163.367
R687 B.n607 B.n606 163.367
R688 B.n606 B.n33 163.367
R689 B.n602 B.n33 163.367
R690 B.n602 B.n601 163.367
R691 B.n601 B.n600 163.367
R692 B.n600 B.n35 163.367
R693 B.n596 B.n35 163.367
R694 B.n596 B.n595 163.367
R695 B.n595 B.n594 163.367
R696 B.n594 B.n37 163.367
R697 B.n590 B.n37 163.367
R698 B.n590 B.n589 163.367
R699 B.n589 B.n588 163.367
R700 B.n588 B.n39 163.367
R701 B.n584 B.n39 163.367
R702 B.n584 B.n583 163.367
R703 B.n583 B.n582 163.367
R704 B.n582 B.n41 163.367
R705 B.n578 B.n41 163.367
R706 B.n578 B.n577 163.367
R707 B.n577 B.n576 163.367
R708 B.n576 B.n43 163.367
R709 B.n572 B.n43 163.367
R710 B.n572 B.n571 163.367
R711 B.n571 B.n570 163.367
R712 B.n570 B.n48 163.367
R713 B.n566 B.n48 163.367
R714 B.n566 B.n565 163.367
R715 B.n565 B.n564 163.367
R716 B.n564 B.n50 163.367
R717 B.n559 B.n50 163.367
R718 B.n559 B.n558 163.367
R719 B.n558 B.n557 163.367
R720 B.n557 B.n54 163.367
R721 B.n553 B.n54 163.367
R722 B.n553 B.n552 163.367
R723 B.n552 B.n551 163.367
R724 B.n551 B.n56 163.367
R725 B.n547 B.n56 163.367
R726 B.n547 B.n546 163.367
R727 B.n546 B.n545 163.367
R728 B.n545 B.n58 163.367
R729 B.n541 B.n58 163.367
R730 B.n541 B.n540 163.367
R731 B.n540 B.n539 163.367
R732 B.n539 B.n60 163.367
R733 B.n535 B.n60 163.367
R734 B.n535 B.n534 163.367
R735 B.n534 B.n533 163.367
R736 B.n533 B.n62 163.367
R737 B.n529 B.n62 163.367
R738 B.n529 B.n528 163.367
R739 B.n528 B.n527 163.367
R740 B.n527 B.n64 163.367
R741 B.n523 B.n64 163.367
R742 B.n523 B.n522 163.367
R743 B.n522 B.n521 163.367
R744 B.n521 B.n66 163.367
R745 B.n517 B.n66 163.367
R746 B.n517 B.n516 163.367
R747 B.n516 B.n515 163.367
R748 B.n515 B.n68 163.367
R749 B.n511 B.n68 163.367
R750 B.n511 B.n510 163.367
R751 B.n510 B.n509 163.367
R752 B.n509 B.n70 163.367
R753 B.n505 B.n70 163.367
R754 B.n505 B.n504 163.367
R755 B.n504 B.n503 163.367
R756 B.n503 B.n72 163.367
R757 B.n499 B.n72 163.367
R758 B.n499 B.n498 163.367
R759 B.n498 B.n497 163.367
R760 B.n497 B.n74 163.367
R761 B.n493 B.n74 163.367
R762 B.n493 B.n492 163.367
R763 B.n492 B.n491 163.367
R764 B.n491 B.n76 163.367
R765 B.n487 B.n76 163.367
R766 B.n487 B.n486 163.367
R767 B.n486 B.n485 163.367
R768 B.n485 B.n78 163.367
R769 B.n481 B.n78 163.367
R770 B.n481 B.n480 163.367
R771 B.n313 B.t8 139.142
R772 B.n51 B.t1 139.142
R773 B.n139 B.t5 139.12
R774 B.n44 B.t10 139.12
R775 B.n314 B.t7 109.856
R776 B.n52 B.t2 109.856
R777 B.n140 B.t4 109.835
R778 B.n45 B.t11 109.835
R779 B.n315 B.n314 59.5399
R780 B.n300 B.n140 59.5399
R781 B.n46 B.n45 59.5399
R782 B.n562 B.n52 59.5399
R783 B.n659 B.n658 32.6249
R784 B.n478 B.n79 32.6249
R785 B.n400 B.n399 32.6249
R786 B.n216 B.n167 32.6249
R787 B.n314 B.n313 29.2853
R788 B.n140 B.n139 29.2853
R789 B.n45 B.n44 29.2853
R790 B.n52 B.n51 29.2853
R791 B B.n699 18.0485
R792 B.n658 B.n657 10.6151
R793 B.n657 B.n16 10.6151
R794 B.n653 B.n16 10.6151
R795 B.n653 B.n652 10.6151
R796 B.n652 B.n651 10.6151
R797 B.n651 B.n18 10.6151
R798 B.n647 B.n18 10.6151
R799 B.n647 B.n646 10.6151
R800 B.n646 B.n645 10.6151
R801 B.n645 B.n20 10.6151
R802 B.n641 B.n20 10.6151
R803 B.n641 B.n640 10.6151
R804 B.n640 B.n639 10.6151
R805 B.n639 B.n22 10.6151
R806 B.n635 B.n22 10.6151
R807 B.n635 B.n634 10.6151
R808 B.n634 B.n633 10.6151
R809 B.n633 B.n24 10.6151
R810 B.n629 B.n24 10.6151
R811 B.n629 B.n628 10.6151
R812 B.n628 B.n627 10.6151
R813 B.n627 B.n26 10.6151
R814 B.n623 B.n26 10.6151
R815 B.n623 B.n622 10.6151
R816 B.n622 B.n621 10.6151
R817 B.n621 B.n28 10.6151
R818 B.n617 B.n28 10.6151
R819 B.n617 B.n616 10.6151
R820 B.n616 B.n615 10.6151
R821 B.n615 B.n30 10.6151
R822 B.n611 B.n30 10.6151
R823 B.n611 B.n610 10.6151
R824 B.n610 B.n609 10.6151
R825 B.n609 B.n32 10.6151
R826 B.n605 B.n32 10.6151
R827 B.n605 B.n604 10.6151
R828 B.n604 B.n603 10.6151
R829 B.n603 B.n34 10.6151
R830 B.n599 B.n34 10.6151
R831 B.n599 B.n598 10.6151
R832 B.n598 B.n597 10.6151
R833 B.n597 B.n36 10.6151
R834 B.n593 B.n36 10.6151
R835 B.n593 B.n592 10.6151
R836 B.n592 B.n591 10.6151
R837 B.n591 B.n38 10.6151
R838 B.n587 B.n38 10.6151
R839 B.n587 B.n586 10.6151
R840 B.n586 B.n585 10.6151
R841 B.n585 B.n40 10.6151
R842 B.n581 B.n40 10.6151
R843 B.n581 B.n580 10.6151
R844 B.n580 B.n579 10.6151
R845 B.n579 B.n42 10.6151
R846 B.n575 B.n574 10.6151
R847 B.n574 B.n573 10.6151
R848 B.n573 B.n47 10.6151
R849 B.n569 B.n47 10.6151
R850 B.n569 B.n568 10.6151
R851 B.n568 B.n567 10.6151
R852 B.n567 B.n49 10.6151
R853 B.n563 B.n49 10.6151
R854 B.n561 B.n560 10.6151
R855 B.n560 B.n53 10.6151
R856 B.n556 B.n53 10.6151
R857 B.n556 B.n555 10.6151
R858 B.n555 B.n554 10.6151
R859 B.n554 B.n55 10.6151
R860 B.n550 B.n55 10.6151
R861 B.n550 B.n549 10.6151
R862 B.n549 B.n548 10.6151
R863 B.n548 B.n57 10.6151
R864 B.n544 B.n57 10.6151
R865 B.n544 B.n543 10.6151
R866 B.n543 B.n542 10.6151
R867 B.n542 B.n59 10.6151
R868 B.n538 B.n59 10.6151
R869 B.n538 B.n537 10.6151
R870 B.n537 B.n536 10.6151
R871 B.n536 B.n61 10.6151
R872 B.n532 B.n61 10.6151
R873 B.n532 B.n531 10.6151
R874 B.n531 B.n530 10.6151
R875 B.n530 B.n63 10.6151
R876 B.n526 B.n63 10.6151
R877 B.n526 B.n525 10.6151
R878 B.n525 B.n524 10.6151
R879 B.n524 B.n65 10.6151
R880 B.n520 B.n65 10.6151
R881 B.n520 B.n519 10.6151
R882 B.n519 B.n518 10.6151
R883 B.n518 B.n67 10.6151
R884 B.n514 B.n67 10.6151
R885 B.n514 B.n513 10.6151
R886 B.n513 B.n512 10.6151
R887 B.n512 B.n69 10.6151
R888 B.n508 B.n69 10.6151
R889 B.n508 B.n507 10.6151
R890 B.n507 B.n506 10.6151
R891 B.n506 B.n71 10.6151
R892 B.n502 B.n71 10.6151
R893 B.n502 B.n501 10.6151
R894 B.n501 B.n500 10.6151
R895 B.n500 B.n73 10.6151
R896 B.n496 B.n73 10.6151
R897 B.n496 B.n495 10.6151
R898 B.n495 B.n494 10.6151
R899 B.n494 B.n75 10.6151
R900 B.n490 B.n75 10.6151
R901 B.n490 B.n489 10.6151
R902 B.n489 B.n488 10.6151
R903 B.n488 B.n77 10.6151
R904 B.n484 B.n77 10.6151
R905 B.n484 B.n483 10.6151
R906 B.n483 B.n482 10.6151
R907 B.n482 B.n79 10.6151
R908 B.n400 B.n105 10.6151
R909 B.n404 B.n105 10.6151
R910 B.n405 B.n404 10.6151
R911 B.n406 B.n405 10.6151
R912 B.n406 B.n103 10.6151
R913 B.n410 B.n103 10.6151
R914 B.n411 B.n410 10.6151
R915 B.n412 B.n411 10.6151
R916 B.n412 B.n101 10.6151
R917 B.n416 B.n101 10.6151
R918 B.n417 B.n416 10.6151
R919 B.n418 B.n417 10.6151
R920 B.n418 B.n99 10.6151
R921 B.n422 B.n99 10.6151
R922 B.n423 B.n422 10.6151
R923 B.n424 B.n423 10.6151
R924 B.n424 B.n97 10.6151
R925 B.n428 B.n97 10.6151
R926 B.n429 B.n428 10.6151
R927 B.n430 B.n429 10.6151
R928 B.n430 B.n95 10.6151
R929 B.n434 B.n95 10.6151
R930 B.n435 B.n434 10.6151
R931 B.n436 B.n435 10.6151
R932 B.n436 B.n93 10.6151
R933 B.n440 B.n93 10.6151
R934 B.n441 B.n440 10.6151
R935 B.n442 B.n441 10.6151
R936 B.n442 B.n91 10.6151
R937 B.n446 B.n91 10.6151
R938 B.n447 B.n446 10.6151
R939 B.n448 B.n447 10.6151
R940 B.n448 B.n89 10.6151
R941 B.n452 B.n89 10.6151
R942 B.n453 B.n452 10.6151
R943 B.n454 B.n453 10.6151
R944 B.n454 B.n87 10.6151
R945 B.n458 B.n87 10.6151
R946 B.n459 B.n458 10.6151
R947 B.n460 B.n459 10.6151
R948 B.n460 B.n85 10.6151
R949 B.n464 B.n85 10.6151
R950 B.n465 B.n464 10.6151
R951 B.n466 B.n465 10.6151
R952 B.n466 B.n83 10.6151
R953 B.n470 B.n83 10.6151
R954 B.n471 B.n470 10.6151
R955 B.n472 B.n471 10.6151
R956 B.n472 B.n81 10.6151
R957 B.n476 B.n81 10.6151
R958 B.n477 B.n476 10.6151
R959 B.n478 B.n477 10.6151
R960 B.n220 B.n167 10.6151
R961 B.n221 B.n220 10.6151
R962 B.n222 B.n221 10.6151
R963 B.n222 B.n165 10.6151
R964 B.n226 B.n165 10.6151
R965 B.n227 B.n226 10.6151
R966 B.n228 B.n227 10.6151
R967 B.n228 B.n163 10.6151
R968 B.n232 B.n163 10.6151
R969 B.n233 B.n232 10.6151
R970 B.n234 B.n233 10.6151
R971 B.n234 B.n161 10.6151
R972 B.n238 B.n161 10.6151
R973 B.n239 B.n238 10.6151
R974 B.n240 B.n239 10.6151
R975 B.n240 B.n159 10.6151
R976 B.n244 B.n159 10.6151
R977 B.n245 B.n244 10.6151
R978 B.n246 B.n245 10.6151
R979 B.n246 B.n157 10.6151
R980 B.n250 B.n157 10.6151
R981 B.n251 B.n250 10.6151
R982 B.n252 B.n251 10.6151
R983 B.n252 B.n155 10.6151
R984 B.n256 B.n155 10.6151
R985 B.n257 B.n256 10.6151
R986 B.n258 B.n257 10.6151
R987 B.n258 B.n153 10.6151
R988 B.n262 B.n153 10.6151
R989 B.n263 B.n262 10.6151
R990 B.n264 B.n263 10.6151
R991 B.n264 B.n151 10.6151
R992 B.n268 B.n151 10.6151
R993 B.n269 B.n268 10.6151
R994 B.n270 B.n269 10.6151
R995 B.n270 B.n149 10.6151
R996 B.n274 B.n149 10.6151
R997 B.n275 B.n274 10.6151
R998 B.n276 B.n275 10.6151
R999 B.n276 B.n147 10.6151
R1000 B.n280 B.n147 10.6151
R1001 B.n281 B.n280 10.6151
R1002 B.n282 B.n281 10.6151
R1003 B.n282 B.n145 10.6151
R1004 B.n286 B.n145 10.6151
R1005 B.n287 B.n286 10.6151
R1006 B.n288 B.n287 10.6151
R1007 B.n288 B.n143 10.6151
R1008 B.n292 B.n143 10.6151
R1009 B.n293 B.n292 10.6151
R1010 B.n294 B.n293 10.6151
R1011 B.n294 B.n141 10.6151
R1012 B.n298 B.n141 10.6151
R1013 B.n299 B.n298 10.6151
R1014 B.n301 B.n137 10.6151
R1015 B.n305 B.n137 10.6151
R1016 B.n306 B.n305 10.6151
R1017 B.n307 B.n306 10.6151
R1018 B.n307 B.n135 10.6151
R1019 B.n311 B.n135 10.6151
R1020 B.n312 B.n311 10.6151
R1021 B.n316 B.n312 10.6151
R1022 B.n320 B.n133 10.6151
R1023 B.n321 B.n320 10.6151
R1024 B.n322 B.n321 10.6151
R1025 B.n322 B.n131 10.6151
R1026 B.n326 B.n131 10.6151
R1027 B.n327 B.n326 10.6151
R1028 B.n328 B.n327 10.6151
R1029 B.n328 B.n129 10.6151
R1030 B.n332 B.n129 10.6151
R1031 B.n333 B.n332 10.6151
R1032 B.n334 B.n333 10.6151
R1033 B.n334 B.n127 10.6151
R1034 B.n338 B.n127 10.6151
R1035 B.n339 B.n338 10.6151
R1036 B.n340 B.n339 10.6151
R1037 B.n340 B.n125 10.6151
R1038 B.n344 B.n125 10.6151
R1039 B.n345 B.n344 10.6151
R1040 B.n346 B.n345 10.6151
R1041 B.n346 B.n123 10.6151
R1042 B.n350 B.n123 10.6151
R1043 B.n351 B.n350 10.6151
R1044 B.n352 B.n351 10.6151
R1045 B.n352 B.n121 10.6151
R1046 B.n356 B.n121 10.6151
R1047 B.n357 B.n356 10.6151
R1048 B.n358 B.n357 10.6151
R1049 B.n358 B.n119 10.6151
R1050 B.n362 B.n119 10.6151
R1051 B.n363 B.n362 10.6151
R1052 B.n364 B.n363 10.6151
R1053 B.n364 B.n117 10.6151
R1054 B.n368 B.n117 10.6151
R1055 B.n369 B.n368 10.6151
R1056 B.n370 B.n369 10.6151
R1057 B.n370 B.n115 10.6151
R1058 B.n374 B.n115 10.6151
R1059 B.n375 B.n374 10.6151
R1060 B.n376 B.n375 10.6151
R1061 B.n376 B.n113 10.6151
R1062 B.n380 B.n113 10.6151
R1063 B.n381 B.n380 10.6151
R1064 B.n382 B.n381 10.6151
R1065 B.n382 B.n111 10.6151
R1066 B.n386 B.n111 10.6151
R1067 B.n387 B.n386 10.6151
R1068 B.n388 B.n387 10.6151
R1069 B.n388 B.n109 10.6151
R1070 B.n392 B.n109 10.6151
R1071 B.n393 B.n392 10.6151
R1072 B.n394 B.n393 10.6151
R1073 B.n394 B.n107 10.6151
R1074 B.n398 B.n107 10.6151
R1075 B.n399 B.n398 10.6151
R1076 B.n216 B.n215 10.6151
R1077 B.n215 B.n214 10.6151
R1078 B.n214 B.n169 10.6151
R1079 B.n210 B.n169 10.6151
R1080 B.n210 B.n209 10.6151
R1081 B.n209 B.n208 10.6151
R1082 B.n208 B.n171 10.6151
R1083 B.n204 B.n171 10.6151
R1084 B.n204 B.n203 10.6151
R1085 B.n203 B.n202 10.6151
R1086 B.n202 B.n173 10.6151
R1087 B.n198 B.n173 10.6151
R1088 B.n198 B.n197 10.6151
R1089 B.n197 B.n196 10.6151
R1090 B.n196 B.n175 10.6151
R1091 B.n192 B.n175 10.6151
R1092 B.n192 B.n191 10.6151
R1093 B.n191 B.n190 10.6151
R1094 B.n190 B.n177 10.6151
R1095 B.n186 B.n177 10.6151
R1096 B.n186 B.n185 10.6151
R1097 B.n185 B.n184 10.6151
R1098 B.n184 B.n179 10.6151
R1099 B.n180 B.n179 10.6151
R1100 B.n180 B.n0 10.6151
R1101 B.n695 B.n1 10.6151
R1102 B.n695 B.n694 10.6151
R1103 B.n694 B.n693 10.6151
R1104 B.n693 B.n4 10.6151
R1105 B.n689 B.n4 10.6151
R1106 B.n689 B.n688 10.6151
R1107 B.n688 B.n687 10.6151
R1108 B.n687 B.n6 10.6151
R1109 B.n683 B.n6 10.6151
R1110 B.n683 B.n682 10.6151
R1111 B.n682 B.n681 10.6151
R1112 B.n681 B.n8 10.6151
R1113 B.n677 B.n8 10.6151
R1114 B.n677 B.n676 10.6151
R1115 B.n676 B.n675 10.6151
R1116 B.n675 B.n10 10.6151
R1117 B.n671 B.n10 10.6151
R1118 B.n671 B.n670 10.6151
R1119 B.n670 B.n669 10.6151
R1120 B.n669 B.n12 10.6151
R1121 B.n665 B.n12 10.6151
R1122 B.n665 B.n664 10.6151
R1123 B.n664 B.n663 10.6151
R1124 B.n663 B.n14 10.6151
R1125 B.n659 B.n14 10.6151
R1126 B.n575 B.n46 6.5566
R1127 B.n563 B.n562 6.5566
R1128 B.n301 B.n300 6.5566
R1129 B.n316 B.n315 6.5566
R1130 B.n46 B.n42 4.05904
R1131 B.n562 B.n561 4.05904
R1132 B.n300 B.n299 4.05904
R1133 B.n315 B.n133 4.05904
R1134 B.n699 B.n0 2.81026
R1135 B.n699 B.n1 2.81026
R1136 VN.n3 VN.t2 367.483
R1137 VN.n13 VN.t1 367.483
R1138 VN.n2 VN.t4 336.993
R1139 VN.n8 VN.t3 336.993
R1140 VN.n12 VN.t5 336.993
R1141 VN.n18 VN.t0 336.993
R1142 VN.n9 VN.n8 173.105
R1143 VN.n19 VN.n18 173.105
R1144 VN.n17 VN.n10 161.3
R1145 VN.n16 VN.n15 161.3
R1146 VN.n14 VN.n11 161.3
R1147 VN.n7 VN.n0 161.3
R1148 VN.n6 VN.n5 161.3
R1149 VN.n4 VN.n1 161.3
R1150 VN.n3 VN.n2 51.5093
R1151 VN.n13 VN.n12 51.5093
R1152 VN VN.n19 46.7865
R1153 VN.n7 VN.n6 41.0614
R1154 VN.n17 VN.n16 41.0614
R1155 VN.n6 VN.n1 40.0926
R1156 VN.n16 VN.n11 40.0926
R1157 VN.n14 VN.n13 26.9198
R1158 VN.n4 VN.n3 26.9198
R1159 VN.n8 VN.n7 12.7883
R1160 VN.n18 VN.n17 12.7883
R1161 VN.n2 VN.n1 12.2964
R1162 VN.n12 VN.n11 12.2964
R1163 VN.n19 VN.n10 0.189894
R1164 VN.n15 VN.n10 0.189894
R1165 VN.n15 VN.n14 0.189894
R1166 VN.n5 VN.n4 0.189894
R1167 VN.n5 VN.n0 0.189894
R1168 VN.n9 VN.n0 0.189894
R1169 VN VN.n9 0.0516364
R1170 VDD2.n1 VDD2.t3 73.6458
R1171 VDD2.n2 VDD2.t5 72.7251
R1172 VDD2.n1 VDD2.n0 71.0249
R1173 VDD2 VDD2.n3 71.0222
R1174 VDD2.n2 VDD2.n1 42.17
R1175 VDD2.n3 VDD2.t0 1.9705
R1176 VDD2.n3 VDD2.t4 1.9705
R1177 VDD2.n0 VDD2.t1 1.9705
R1178 VDD2.n0 VDD2.t2 1.9705
R1179 VDD2 VDD2.n2 1.03498
C0 VDD1 VDD2 0.886533f
C1 VP w_n2178_n4268# 4.15273f
C2 VN B 0.92205f
C3 VP VTAIL 6.99554f
C4 VDD2 w_n2178_n4268# 2.29909f
C5 VDD1 VN 0.148902f
C6 VTAIL VDD2 10.7634f
C7 VN w_n2178_n4268# 3.8751f
C8 VP VDD2 0.338811f
C9 VDD1 B 2.04092f
C10 VTAIL VN 6.98092f
C11 VP VN 6.37974f
C12 w_n2178_n4268# B 8.976919f
C13 VDD1 w_n2178_n4268# 2.25984f
C14 VTAIL B 3.87922f
C15 VN VDD2 7.33313f
C16 VP B 1.37843f
C17 VTAIL VDD1 10.7265f
C18 VP VDD1 7.51779f
C19 VDD2 B 2.08119f
C20 VTAIL w_n2178_n4268# 3.56499f
C21 VDD2 VSUBS 1.683068f
C22 VDD1 VSUBS 2.03744f
C23 VTAIL VSUBS 1.046914f
C24 VN VSUBS 4.95376f
C25 VP VSUBS 1.992214f
C26 B VSUBS 3.617272f
C27 w_n2178_n4268# VSUBS 0.113822p
C28 VDD2.t3 VSUBS 3.82043f
C29 VDD2.t1 VSUBS 0.3566f
C30 VDD2.t2 VSUBS 0.3566f
C31 VDD2.n0 VSUBS 2.9377f
C32 VDD2.n1 VSUBS 3.43684f
C33 VDD2.t5 VSUBS 3.81147f
C34 VDD2.n2 VSUBS 3.34049f
C35 VDD2.t0 VSUBS 0.3566f
C36 VDD2.t4 VSUBS 0.3566f
C37 VDD2.n3 VSUBS 2.93765f
C38 VN.n0 VSUBS 0.043065f
C39 VN.t3 VSUBS 2.30232f
C40 VN.n1 VSUBS 0.065634f
C41 VN.t2 VSUBS 2.38099f
C42 VN.t4 VSUBS 2.30232f
C43 VN.n2 VSUBS 0.885643f
C44 VN.n3 VSUBS 0.919643f
C45 VN.n4 VSUBS 0.223609f
C46 VN.n5 VSUBS 0.043065f
C47 VN.n6 VSUBS 0.034796f
C48 VN.n7 VSUBS 0.065996f
C49 VN.n8 VSUBS 0.892693f
C50 VN.n9 VSUBS 0.038497f
C51 VN.n10 VSUBS 0.043065f
C52 VN.t0 VSUBS 2.30232f
C53 VN.n11 VSUBS 0.065634f
C54 VN.t1 VSUBS 2.38099f
C55 VN.t5 VSUBS 2.30232f
C56 VN.n12 VSUBS 0.885643f
C57 VN.n13 VSUBS 0.919643f
C58 VN.n14 VSUBS 0.223609f
C59 VN.n15 VSUBS 0.043065f
C60 VN.n16 VSUBS 0.034796f
C61 VN.n17 VSUBS 0.065996f
C62 VN.n18 VSUBS 0.892693f
C63 VN.n19 VSUBS 2.12134f
C64 B.n0 VSUBS 0.005402f
C65 B.n1 VSUBS 0.005402f
C66 B.n2 VSUBS 0.008543f
C67 B.n3 VSUBS 0.008543f
C68 B.n4 VSUBS 0.008543f
C69 B.n5 VSUBS 0.008543f
C70 B.n6 VSUBS 0.008543f
C71 B.n7 VSUBS 0.008543f
C72 B.n8 VSUBS 0.008543f
C73 B.n9 VSUBS 0.008543f
C74 B.n10 VSUBS 0.008543f
C75 B.n11 VSUBS 0.008543f
C76 B.n12 VSUBS 0.008543f
C77 B.n13 VSUBS 0.008543f
C78 B.n14 VSUBS 0.008543f
C79 B.n15 VSUBS 0.020235f
C80 B.n16 VSUBS 0.008543f
C81 B.n17 VSUBS 0.008543f
C82 B.n18 VSUBS 0.008543f
C83 B.n19 VSUBS 0.008543f
C84 B.n20 VSUBS 0.008543f
C85 B.n21 VSUBS 0.008543f
C86 B.n22 VSUBS 0.008543f
C87 B.n23 VSUBS 0.008543f
C88 B.n24 VSUBS 0.008543f
C89 B.n25 VSUBS 0.008543f
C90 B.n26 VSUBS 0.008543f
C91 B.n27 VSUBS 0.008543f
C92 B.n28 VSUBS 0.008543f
C93 B.n29 VSUBS 0.008543f
C94 B.n30 VSUBS 0.008543f
C95 B.n31 VSUBS 0.008543f
C96 B.n32 VSUBS 0.008543f
C97 B.n33 VSUBS 0.008543f
C98 B.n34 VSUBS 0.008543f
C99 B.n35 VSUBS 0.008543f
C100 B.n36 VSUBS 0.008543f
C101 B.n37 VSUBS 0.008543f
C102 B.n38 VSUBS 0.008543f
C103 B.n39 VSUBS 0.008543f
C104 B.n40 VSUBS 0.008543f
C105 B.n41 VSUBS 0.008543f
C106 B.n42 VSUBS 0.005905f
C107 B.n43 VSUBS 0.008543f
C108 B.t11 VSUBS 0.675529f
C109 B.t10 VSUBS 0.68996f
C110 B.t9 VSUBS 0.997916f
C111 B.n44 VSUBS 0.271363f
C112 B.n45 VSUBS 0.080743f
C113 B.n46 VSUBS 0.019793f
C114 B.n47 VSUBS 0.008543f
C115 B.n48 VSUBS 0.008543f
C116 B.n49 VSUBS 0.008543f
C117 B.n50 VSUBS 0.008543f
C118 B.t2 VSUBS 0.675507f
C119 B.t1 VSUBS 0.689941f
C120 B.t0 VSUBS 0.997916f
C121 B.n51 VSUBS 0.271383f
C122 B.n52 VSUBS 0.080765f
C123 B.n53 VSUBS 0.008543f
C124 B.n54 VSUBS 0.008543f
C125 B.n55 VSUBS 0.008543f
C126 B.n56 VSUBS 0.008543f
C127 B.n57 VSUBS 0.008543f
C128 B.n58 VSUBS 0.008543f
C129 B.n59 VSUBS 0.008543f
C130 B.n60 VSUBS 0.008543f
C131 B.n61 VSUBS 0.008543f
C132 B.n62 VSUBS 0.008543f
C133 B.n63 VSUBS 0.008543f
C134 B.n64 VSUBS 0.008543f
C135 B.n65 VSUBS 0.008543f
C136 B.n66 VSUBS 0.008543f
C137 B.n67 VSUBS 0.008543f
C138 B.n68 VSUBS 0.008543f
C139 B.n69 VSUBS 0.008543f
C140 B.n70 VSUBS 0.008543f
C141 B.n71 VSUBS 0.008543f
C142 B.n72 VSUBS 0.008543f
C143 B.n73 VSUBS 0.008543f
C144 B.n74 VSUBS 0.008543f
C145 B.n75 VSUBS 0.008543f
C146 B.n76 VSUBS 0.008543f
C147 B.n77 VSUBS 0.008543f
C148 B.n78 VSUBS 0.008543f
C149 B.n79 VSUBS 0.019224f
C150 B.n80 VSUBS 0.008543f
C151 B.n81 VSUBS 0.008543f
C152 B.n82 VSUBS 0.008543f
C153 B.n83 VSUBS 0.008543f
C154 B.n84 VSUBS 0.008543f
C155 B.n85 VSUBS 0.008543f
C156 B.n86 VSUBS 0.008543f
C157 B.n87 VSUBS 0.008543f
C158 B.n88 VSUBS 0.008543f
C159 B.n89 VSUBS 0.008543f
C160 B.n90 VSUBS 0.008543f
C161 B.n91 VSUBS 0.008543f
C162 B.n92 VSUBS 0.008543f
C163 B.n93 VSUBS 0.008543f
C164 B.n94 VSUBS 0.008543f
C165 B.n95 VSUBS 0.008543f
C166 B.n96 VSUBS 0.008543f
C167 B.n97 VSUBS 0.008543f
C168 B.n98 VSUBS 0.008543f
C169 B.n99 VSUBS 0.008543f
C170 B.n100 VSUBS 0.008543f
C171 B.n101 VSUBS 0.008543f
C172 B.n102 VSUBS 0.008543f
C173 B.n103 VSUBS 0.008543f
C174 B.n104 VSUBS 0.008543f
C175 B.n105 VSUBS 0.008543f
C176 B.n106 VSUBS 0.020235f
C177 B.n107 VSUBS 0.008543f
C178 B.n108 VSUBS 0.008543f
C179 B.n109 VSUBS 0.008543f
C180 B.n110 VSUBS 0.008543f
C181 B.n111 VSUBS 0.008543f
C182 B.n112 VSUBS 0.008543f
C183 B.n113 VSUBS 0.008543f
C184 B.n114 VSUBS 0.008543f
C185 B.n115 VSUBS 0.008543f
C186 B.n116 VSUBS 0.008543f
C187 B.n117 VSUBS 0.008543f
C188 B.n118 VSUBS 0.008543f
C189 B.n119 VSUBS 0.008543f
C190 B.n120 VSUBS 0.008543f
C191 B.n121 VSUBS 0.008543f
C192 B.n122 VSUBS 0.008543f
C193 B.n123 VSUBS 0.008543f
C194 B.n124 VSUBS 0.008543f
C195 B.n125 VSUBS 0.008543f
C196 B.n126 VSUBS 0.008543f
C197 B.n127 VSUBS 0.008543f
C198 B.n128 VSUBS 0.008543f
C199 B.n129 VSUBS 0.008543f
C200 B.n130 VSUBS 0.008543f
C201 B.n131 VSUBS 0.008543f
C202 B.n132 VSUBS 0.008543f
C203 B.n133 VSUBS 0.005905f
C204 B.n134 VSUBS 0.008543f
C205 B.n135 VSUBS 0.008543f
C206 B.n136 VSUBS 0.008543f
C207 B.n137 VSUBS 0.008543f
C208 B.n138 VSUBS 0.008543f
C209 B.t4 VSUBS 0.675529f
C210 B.t5 VSUBS 0.68996f
C211 B.t3 VSUBS 0.997916f
C212 B.n139 VSUBS 0.271363f
C213 B.n140 VSUBS 0.080743f
C214 B.n141 VSUBS 0.008543f
C215 B.n142 VSUBS 0.008543f
C216 B.n143 VSUBS 0.008543f
C217 B.n144 VSUBS 0.008543f
C218 B.n145 VSUBS 0.008543f
C219 B.n146 VSUBS 0.008543f
C220 B.n147 VSUBS 0.008543f
C221 B.n148 VSUBS 0.008543f
C222 B.n149 VSUBS 0.008543f
C223 B.n150 VSUBS 0.008543f
C224 B.n151 VSUBS 0.008543f
C225 B.n152 VSUBS 0.008543f
C226 B.n153 VSUBS 0.008543f
C227 B.n154 VSUBS 0.008543f
C228 B.n155 VSUBS 0.008543f
C229 B.n156 VSUBS 0.008543f
C230 B.n157 VSUBS 0.008543f
C231 B.n158 VSUBS 0.008543f
C232 B.n159 VSUBS 0.008543f
C233 B.n160 VSUBS 0.008543f
C234 B.n161 VSUBS 0.008543f
C235 B.n162 VSUBS 0.008543f
C236 B.n163 VSUBS 0.008543f
C237 B.n164 VSUBS 0.008543f
C238 B.n165 VSUBS 0.008543f
C239 B.n166 VSUBS 0.008543f
C240 B.n167 VSUBS 0.020235f
C241 B.n168 VSUBS 0.008543f
C242 B.n169 VSUBS 0.008543f
C243 B.n170 VSUBS 0.008543f
C244 B.n171 VSUBS 0.008543f
C245 B.n172 VSUBS 0.008543f
C246 B.n173 VSUBS 0.008543f
C247 B.n174 VSUBS 0.008543f
C248 B.n175 VSUBS 0.008543f
C249 B.n176 VSUBS 0.008543f
C250 B.n177 VSUBS 0.008543f
C251 B.n178 VSUBS 0.008543f
C252 B.n179 VSUBS 0.008543f
C253 B.n180 VSUBS 0.008543f
C254 B.n181 VSUBS 0.008543f
C255 B.n182 VSUBS 0.008543f
C256 B.n183 VSUBS 0.008543f
C257 B.n184 VSUBS 0.008543f
C258 B.n185 VSUBS 0.008543f
C259 B.n186 VSUBS 0.008543f
C260 B.n187 VSUBS 0.008543f
C261 B.n188 VSUBS 0.008543f
C262 B.n189 VSUBS 0.008543f
C263 B.n190 VSUBS 0.008543f
C264 B.n191 VSUBS 0.008543f
C265 B.n192 VSUBS 0.008543f
C266 B.n193 VSUBS 0.008543f
C267 B.n194 VSUBS 0.008543f
C268 B.n195 VSUBS 0.008543f
C269 B.n196 VSUBS 0.008543f
C270 B.n197 VSUBS 0.008543f
C271 B.n198 VSUBS 0.008543f
C272 B.n199 VSUBS 0.008543f
C273 B.n200 VSUBS 0.008543f
C274 B.n201 VSUBS 0.008543f
C275 B.n202 VSUBS 0.008543f
C276 B.n203 VSUBS 0.008543f
C277 B.n204 VSUBS 0.008543f
C278 B.n205 VSUBS 0.008543f
C279 B.n206 VSUBS 0.008543f
C280 B.n207 VSUBS 0.008543f
C281 B.n208 VSUBS 0.008543f
C282 B.n209 VSUBS 0.008543f
C283 B.n210 VSUBS 0.008543f
C284 B.n211 VSUBS 0.008543f
C285 B.n212 VSUBS 0.008543f
C286 B.n213 VSUBS 0.008543f
C287 B.n214 VSUBS 0.008543f
C288 B.n215 VSUBS 0.008543f
C289 B.n216 VSUBS 0.019717f
C290 B.n217 VSUBS 0.019717f
C291 B.n218 VSUBS 0.020235f
C292 B.n219 VSUBS 0.008543f
C293 B.n220 VSUBS 0.008543f
C294 B.n221 VSUBS 0.008543f
C295 B.n222 VSUBS 0.008543f
C296 B.n223 VSUBS 0.008543f
C297 B.n224 VSUBS 0.008543f
C298 B.n225 VSUBS 0.008543f
C299 B.n226 VSUBS 0.008543f
C300 B.n227 VSUBS 0.008543f
C301 B.n228 VSUBS 0.008543f
C302 B.n229 VSUBS 0.008543f
C303 B.n230 VSUBS 0.008543f
C304 B.n231 VSUBS 0.008543f
C305 B.n232 VSUBS 0.008543f
C306 B.n233 VSUBS 0.008543f
C307 B.n234 VSUBS 0.008543f
C308 B.n235 VSUBS 0.008543f
C309 B.n236 VSUBS 0.008543f
C310 B.n237 VSUBS 0.008543f
C311 B.n238 VSUBS 0.008543f
C312 B.n239 VSUBS 0.008543f
C313 B.n240 VSUBS 0.008543f
C314 B.n241 VSUBS 0.008543f
C315 B.n242 VSUBS 0.008543f
C316 B.n243 VSUBS 0.008543f
C317 B.n244 VSUBS 0.008543f
C318 B.n245 VSUBS 0.008543f
C319 B.n246 VSUBS 0.008543f
C320 B.n247 VSUBS 0.008543f
C321 B.n248 VSUBS 0.008543f
C322 B.n249 VSUBS 0.008543f
C323 B.n250 VSUBS 0.008543f
C324 B.n251 VSUBS 0.008543f
C325 B.n252 VSUBS 0.008543f
C326 B.n253 VSUBS 0.008543f
C327 B.n254 VSUBS 0.008543f
C328 B.n255 VSUBS 0.008543f
C329 B.n256 VSUBS 0.008543f
C330 B.n257 VSUBS 0.008543f
C331 B.n258 VSUBS 0.008543f
C332 B.n259 VSUBS 0.008543f
C333 B.n260 VSUBS 0.008543f
C334 B.n261 VSUBS 0.008543f
C335 B.n262 VSUBS 0.008543f
C336 B.n263 VSUBS 0.008543f
C337 B.n264 VSUBS 0.008543f
C338 B.n265 VSUBS 0.008543f
C339 B.n266 VSUBS 0.008543f
C340 B.n267 VSUBS 0.008543f
C341 B.n268 VSUBS 0.008543f
C342 B.n269 VSUBS 0.008543f
C343 B.n270 VSUBS 0.008543f
C344 B.n271 VSUBS 0.008543f
C345 B.n272 VSUBS 0.008543f
C346 B.n273 VSUBS 0.008543f
C347 B.n274 VSUBS 0.008543f
C348 B.n275 VSUBS 0.008543f
C349 B.n276 VSUBS 0.008543f
C350 B.n277 VSUBS 0.008543f
C351 B.n278 VSUBS 0.008543f
C352 B.n279 VSUBS 0.008543f
C353 B.n280 VSUBS 0.008543f
C354 B.n281 VSUBS 0.008543f
C355 B.n282 VSUBS 0.008543f
C356 B.n283 VSUBS 0.008543f
C357 B.n284 VSUBS 0.008543f
C358 B.n285 VSUBS 0.008543f
C359 B.n286 VSUBS 0.008543f
C360 B.n287 VSUBS 0.008543f
C361 B.n288 VSUBS 0.008543f
C362 B.n289 VSUBS 0.008543f
C363 B.n290 VSUBS 0.008543f
C364 B.n291 VSUBS 0.008543f
C365 B.n292 VSUBS 0.008543f
C366 B.n293 VSUBS 0.008543f
C367 B.n294 VSUBS 0.008543f
C368 B.n295 VSUBS 0.008543f
C369 B.n296 VSUBS 0.008543f
C370 B.n297 VSUBS 0.008543f
C371 B.n298 VSUBS 0.008543f
C372 B.n299 VSUBS 0.005905f
C373 B.n300 VSUBS 0.019793f
C374 B.n301 VSUBS 0.00691f
C375 B.n302 VSUBS 0.008543f
C376 B.n303 VSUBS 0.008543f
C377 B.n304 VSUBS 0.008543f
C378 B.n305 VSUBS 0.008543f
C379 B.n306 VSUBS 0.008543f
C380 B.n307 VSUBS 0.008543f
C381 B.n308 VSUBS 0.008543f
C382 B.n309 VSUBS 0.008543f
C383 B.n310 VSUBS 0.008543f
C384 B.n311 VSUBS 0.008543f
C385 B.n312 VSUBS 0.008543f
C386 B.t7 VSUBS 0.675507f
C387 B.t8 VSUBS 0.689941f
C388 B.t6 VSUBS 0.997916f
C389 B.n313 VSUBS 0.271383f
C390 B.n314 VSUBS 0.080765f
C391 B.n315 VSUBS 0.019793f
C392 B.n316 VSUBS 0.00691f
C393 B.n317 VSUBS 0.008543f
C394 B.n318 VSUBS 0.008543f
C395 B.n319 VSUBS 0.008543f
C396 B.n320 VSUBS 0.008543f
C397 B.n321 VSUBS 0.008543f
C398 B.n322 VSUBS 0.008543f
C399 B.n323 VSUBS 0.008543f
C400 B.n324 VSUBS 0.008543f
C401 B.n325 VSUBS 0.008543f
C402 B.n326 VSUBS 0.008543f
C403 B.n327 VSUBS 0.008543f
C404 B.n328 VSUBS 0.008543f
C405 B.n329 VSUBS 0.008543f
C406 B.n330 VSUBS 0.008543f
C407 B.n331 VSUBS 0.008543f
C408 B.n332 VSUBS 0.008543f
C409 B.n333 VSUBS 0.008543f
C410 B.n334 VSUBS 0.008543f
C411 B.n335 VSUBS 0.008543f
C412 B.n336 VSUBS 0.008543f
C413 B.n337 VSUBS 0.008543f
C414 B.n338 VSUBS 0.008543f
C415 B.n339 VSUBS 0.008543f
C416 B.n340 VSUBS 0.008543f
C417 B.n341 VSUBS 0.008543f
C418 B.n342 VSUBS 0.008543f
C419 B.n343 VSUBS 0.008543f
C420 B.n344 VSUBS 0.008543f
C421 B.n345 VSUBS 0.008543f
C422 B.n346 VSUBS 0.008543f
C423 B.n347 VSUBS 0.008543f
C424 B.n348 VSUBS 0.008543f
C425 B.n349 VSUBS 0.008543f
C426 B.n350 VSUBS 0.008543f
C427 B.n351 VSUBS 0.008543f
C428 B.n352 VSUBS 0.008543f
C429 B.n353 VSUBS 0.008543f
C430 B.n354 VSUBS 0.008543f
C431 B.n355 VSUBS 0.008543f
C432 B.n356 VSUBS 0.008543f
C433 B.n357 VSUBS 0.008543f
C434 B.n358 VSUBS 0.008543f
C435 B.n359 VSUBS 0.008543f
C436 B.n360 VSUBS 0.008543f
C437 B.n361 VSUBS 0.008543f
C438 B.n362 VSUBS 0.008543f
C439 B.n363 VSUBS 0.008543f
C440 B.n364 VSUBS 0.008543f
C441 B.n365 VSUBS 0.008543f
C442 B.n366 VSUBS 0.008543f
C443 B.n367 VSUBS 0.008543f
C444 B.n368 VSUBS 0.008543f
C445 B.n369 VSUBS 0.008543f
C446 B.n370 VSUBS 0.008543f
C447 B.n371 VSUBS 0.008543f
C448 B.n372 VSUBS 0.008543f
C449 B.n373 VSUBS 0.008543f
C450 B.n374 VSUBS 0.008543f
C451 B.n375 VSUBS 0.008543f
C452 B.n376 VSUBS 0.008543f
C453 B.n377 VSUBS 0.008543f
C454 B.n378 VSUBS 0.008543f
C455 B.n379 VSUBS 0.008543f
C456 B.n380 VSUBS 0.008543f
C457 B.n381 VSUBS 0.008543f
C458 B.n382 VSUBS 0.008543f
C459 B.n383 VSUBS 0.008543f
C460 B.n384 VSUBS 0.008543f
C461 B.n385 VSUBS 0.008543f
C462 B.n386 VSUBS 0.008543f
C463 B.n387 VSUBS 0.008543f
C464 B.n388 VSUBS 0.008543f
C465 B.n389 VSUBS 0.008543f
C466 B.n390 VSUBS 0.008543f
C467 B.n391 VSUBS 0.008543f
C468 B.n392 VSUBS 0.008543f
C469 B.n393 VSUBS 0.008543f
C470 B.n394 VSUBS 0.008543f
C471 B.n395 VSUBS 0.008543f
C472 B.n396 VSUBS 0.008543f
C473 B.n397 VSUBS 0.008543f
C474 B.n398 VSUBS 0.008543f
C475 B.n399 VSUBS 0.020235f
C476 B.n400 VSUBS 0.019717f
C477 B.n401 VSUBS 0.019717f
C478 B.n402 VSUBS 0.008543f
C479 B.n403 VSUBS 0.008543f
C480 B.n404 VSUBS 0.008543f
C481 B.n405 VSUBS 0.008543f
C482 B.n406 VSUBS 0.008543f
C483 B.n407 VSUBS 0.008543f
C484 B.n408 VSUBS 0.008543f
C485 B.n409 VSUBS 0.008543f
C486 B.n410 VSUBS 0.008543f
C487 B.n411 VSUBS 0.008543f
C488 B.n412 VSUBS 0.008543f
C489 B.n413 VSUBS 0.008543f
C490 B.n414 VSUBS 0.008543f
C491 B.n415 VSUBS 0.008543f
C492 B.n416 VSUBS 0.008543f
C493 B.n417 VSUBS 0.008543f
C494 B.n418 VSUBS 0.008543f
C495 B.n419 VSUBS 0.008543f
C496 B.n420 VSUBS 0.008543f
C497 B.n421 VSUBS 0.008543f
C498 B.n422 VSUBS 0.008543f
C499 B.n423 VSUBS 0.008543f
C500 B.n424 VSUBS 0.008543f
C501 B.n425 VSUBS 0.008543f
C502 B.n426 VSUBS 0.008543f
C503 B.n427 VSUBS 0.008543f
C504 B.n428 VSUBS 0.008543f
C505 B.n429 VSUBS 0.008543f
C506 B.n430 VSUBS 0.008543f
C507 B.n431 VSUBS 0.008543f
C508 B.n432 VSUBS 0.008543f
C509 B.n433 VSUBS 0.008543f
C510 B.n434 VSUBS 0.008543f
C511 B.n435 VSUBS 0.008543f
C512 B.n436 VSUBS 0.008543f
C513 B.n437 VSUBS 0.008543f
C514 B.n438 VSUBS 0.008543f
C515 B.n439 VSUBS 0.008543f
C516 B.n440 VSUBS 0.008543f
C517 B.n441 VSUBS 0.008543f
C518 B.n442 VSUBS 0.008543f
C519 B.n443 VSUBS 0.008543f
C520 B.n444 VSUBS 0.008543f
C521 B.n445 VSUBS 0.008543f
C522 B.n446 VSUBS 0.008543f
C523 B.n447 VSUBS 0.008543f
C524 B.n448 VSUBS 0.008543f
C525 B.n449 VSUBS 0.008543f
C526 B.n450 VSUBS 0.008543f
C527 B.n451 VSUBS 0.008543f
C528 B.n452 VSUBS 0.008543f
C529 B.n453 VSUBS 0.008543f
C530 B.n454 VSUBS 0.008543f
C531 B.n455 VSUBS 0.008543f
C532 B.n456 VSUBS 0.008543f
C533 B.n457 VSUBS 0.008543f
C534 B.n458 VSUBS 0.008543f
C535 B.n459 VSUBS 0.008543f
C536 B.n460 VSUBS 0.008543f
C537 B.n461 VSUBS 0.008543f
C538 B.n462 VSUBS 0.008543f
C539 B.n463 VSUBS 0.008543f
C540 B.n464 VSUBS 0.008543f
C541 B.n465 VSUBS 0.008543f
C542 B.n466 VSUBS 0.008543f
C543 B.n467 VSUBS 0.008543f
C544 B.n468 VSUBS 0.008543f
C545 B.n469 VSUBS 0.008543f
C546 B.n470 VSUBS 0.008543f
C547 B.n471 VSUBS 0.008543f
C548 B.n472 VSUBS 0.008543f
C549 B.n473 VSUBS 0.008543f
C550 B.n474 VSUBS 0.008543f
C551 B.n475 VSUBS 0.008543f
C552 B.n476 VSUBS 0.008543f
C553 B.n477 VSUBS 0.008543f
C554 B.n478 VSUBS 0.020727f
C555 B.n479 VSUBS 0.019717f
C556 B.n480 VSUBS 0.020235f
C557 B.n481 VSUBS 0.008543f
C558 B.n482 VSUBS 0.008543f
C559 B.n483 VSUBS 0.008543f
C560 B.n484 VSUBS 0.008543f
C561 B.n485 VSUBS 0.008543f
C562 B.n486 VSUBS 0.008543f
C563 B.n487 VSUBS 0.008543f
C564 B.n488 VSUBS 0.008543f
C565 B.n489 VSUBS 0.008543f
C566 B.n490 VSUBS 0.008543f
C567 B.n491 VSUBS 0.008543f
C568 B.n492 VSUBS 0.008543f
C569 B.n493 VSUBS 0.008543f
C570 B.n494 VSUBS 0.008543f
C571 B.n495 VSUBS 0.008543f
C572 B.n496 VSUBS 0.008543f
C573 B.n497 VSUBS 0.008543f
C574 B.n498 VSUBS 0.008543f
C575 B.n499 VSUBS 0.008543f
C576 B.n500 VSUBS 0.008543f
C577 B.n501 VSUBS 0.008543f
C578 B.n502 VSUBS 0.008543f
C579 B.n503 VSUBS 0.008543f
C580 B.n504 VSUBS 0.008543f
C581 B.n505 VSUBS 0.008543f
C582 B.n506 VSUBS 0.008543f
C583 B.n507 VSUBS 0.008543f
C584 B.n508 VSUBS 0.008543f
C585 B.n509 VSUBS 0.008543f
C586 B.n510 VSUBS 0.008543f
C587 B.n511 VSUBS 0.008543f
C588 B.n512 VSUBS 0.008543f
C589 B.n513 VSUBS 0.008543f
C590 B.n514 VSUBS 0.008543f
C591 B.n515 VSUBS 0.008543f
C592 B.n516 VSUBS 0.008543f
C593 B.n517 VSUBS 0.008543f
C594 B.n518 VSUBS 0.008543f
C595 B.n519 VSUBS 0.008543f
C596 B.n520 VSUBS 0.008543f
C597 B.n521 VSUBS 0.008543f
C598 B.n522 VSUBS 0.008543f
C599 B.n523 VSUBS 0.008543f
C600 B.n524 VSUBS 0.008543f
C601 B.n525 VSUBS 0.008543f
C602 B.n526 VSUBS 0.008543f
C603 B.n527 VSUBS 0.008543f
C604 B.n528 VSUBS 0.008543f
C605 B.n529 VSUBS 0.008543f
C606 B.n530 VSUBS 0.008543f
C607 B.n531 VSUBS 0.008543f
C608 B.n532 VSUBS 0.008543f
C609 B.n533 VSUBS 0.008543f
C610 B.n534 VSUBS 0.008543f
C611 B.n535 VSUBS 0.008543f
C612 B.n536 VSUBS 0.008543f
C613 B.n537 VSUBS 0.008543f
C614 B.n538 VSUBS 0.008543f
C615 B.n539 VSUBS 0.008543f
C616 B.n540 VSUBS 0.008543f
C617 B.n541 VSUBS 0.008543f
C618 B.n542 VSUBS 0.008543f
C619 B.n543 VSUBS 0.008543f
C620 B.n544 VSUBS 0.008543f
C621 B.n545 VSUBS 0.008543f
C622 B.n546 VSUBS 0.008543f
C623 B.n547 VSUBS 0.008543f
C624 B.n548 VSUBS 0.008543f
C625 B.n549 VSUBS 0.008543f
C626 B.n550 VSUBS 0.008543f
C627 B.n551 VSUBS 0.008543f
C628 B.n552 VSUBS 0.008543f
C629 B.n553 VSUBS 0.008543f
C630 B.n554 VSUBS 0.008543f
C631 B.n555 VSUBS 0.008543f
C632 B.n556 VSUBS 0.008543f
C633 B.n557 VSUBS 0.008543f
C634 B.n558 VSUBS 0.008543f
C635 B.n559 VSUBS 0.008543f
C636 B.n560 VSUBS 0.008543f
C637 B.n561 VSUBS 0.005905f
C638 B.n562 VSUBS 0.019793f
C639 B.n563 VSUBS 0.00691f
C640 B.n564 VSUBS 0.008543f
C641 B.n565 VSUBS 0.008543f
C642 B.n566 VSUBS 0.008543f
C643 B.n567 VSUBS 0.008543f
C644 B.n568 VSUBS 0.008543f
C645 B.n569 VSUBS 0.008543f
C646 B.n570 VSUBS 0.008543f
C647 B.n571 VSUBS 0.008543f
C648 B.n572 VSUBS 0.008543f
C649 B.n573 VSUBS 0.008543f
C650 B.n574 VSUBS 0.008543f
C651 B.n575 VSUBS 0.00691f
C652 B.n576 VSUBS 0.008543f
C653 B.n577 VSUBS 0.008543f
C654 B.n578 VSUBS 0.008543f
C655 B.n579 VSUBS 0.008543f
C656 B.n580 VSUBS 0.008543f
C657 B.n581 VSUBS 0.008543f
C658 B.n582 VSUBS 0.008543f
C659 B.n583 VSUBS 0.008543f
C660 B.n584 VSUBS 0.008543f
C661 B.n585 VSUBS 0.008543f
C662 B.n586 VSUBS 0.008543f
C663 B.n587 VSUBS 0.008543f
C664 B.n588 VSUBS 0.008543f
C665 B.n589 VSUBS 0.008543f
C666 B.n590 VSUBS 0.008543f
C667 B.n591 VSUBS 0.008543f
C668 B.n592 VSUBS 0.008543f
C669 B.n593 VSUBS 0.008543f
C670 B.n594 VSUBS 0.008543f
C671 B.n595 VSUBS 0.008543f
C672 B.n596 VSUBS 0.008543f
C673 B.n597 VSUBS 0.008543f
C674 B.n598 VSUBS 0.008543f
C675 B.n599 VSUBS 0.008543f
C676 B.n600 VSUBS 0.008543f
C677 B.n601 VSUBS 0.008543f
C678 B.n602 VSUBS 0.008543f
C679 B.n603 VSUBS 0.008543f
C680 B.n604 VSUBS 0.008543f
C681 B.n605 VSUBS 0.008543f
C682 B.n606 VSUBS 0.008543f
C683 B.n607 VSUBS 0.008543f
C684 B.n608 VSUBS 0.008543f
C685 B.n609 VSUBS 0.008543f
C686 B.n610 VSUBS 0.008543f
C687 B.n611 VSUBS 0.008543f
C688 B.n612 VSUBS 0.008543f
C689 B.n613 VSUBS 0.008543f
C690 B.n614 VSUBS 0.008543f
C691 B.n615 VSUBS 0.008543f
C692 B.n616 VSUBS 0.008543f
C693 B.n617 VSUBS 0.008543f
C694 B.n618 VSUBS 0.008543f
C695 B.n619 VSUBS 0.008543f
C696 B.n620 VSUBS 0.008543f
C697 B.n621 VSUBS 0.008543f
C698 B.n622 VSUBS 0.008543f
C699 B.n623 VSUBS 0.008543f
C700 B.n624 VSUBS 0.008543f
C701 B.n625 VSUBS 0.008543f
C702 B.n626 VSUBS 0.008543f
C703 B.n627 VSUBS 0.008543f
C704 B.n628 VSUBS 0.008543f
C705 B.n629 VSUBS 0.008543f
C706 B.n630 VSUBS 0.008543f
C707 B.n631 VSUBS 0.008543f
C708 B.n632 VSUBS 0.008543f
C709 B.n633 VSUBS 0.008543f
C710 B.n634 VSUBS 0.008543f
C711 B.n635 VSUBS 0.008543f
C712 B.n636 VSUBS 0.008543f
C713 B.n637 VSUBS 0.008543f
C714 B.n638 VSUBS 0.008543f
C715 B.n639 VSUBS 0.008543f
C716 B.n640 VSUBS 0.008543f
C717 B.n641 VSUBS 0.008543f
C718 B.n642 VSUBS 0.008543f
C719 B.n643 VSUBS 0.008543f
C720 B.n644 VSUBS 0.008543f
C721 B.n645 VSUBS 0.008543f
C722 B.n646 VSUBS 0.008543f
C723 B.n647 VSUBS 0.008543f
C724 B.n648 VSUBS 0.008543f
C725 B.n649 VSUBS 0.008543f
C726 B.n650 VSUBS 0.008543f
C727 B.n651 VSUBS 0.008543f
C728 B.n652 VSUBS 0.008543f
C729 B.n653 VSUBS 0.008543f
C730 B.n654 VSUBS 0.008543f
C731 B.n655 VSUBS 0.008543f
C732 B.n656 VSUBS 0.008543f
C733 B.n657 VSUBS 0.008543f
C734 B.n658 VSUBS 0.020235f
C735 B.n659 VSUBS 0.019717f
C736 B.n660 VSUBS 0.019717f
C737 B.n661 VSUBS 0.008543f
C738 B.n662 VSUBS 0.008543f
C739 B.n663 VSUBS 0.008543f
C740 B.n664 VSUBS 0.008543f
C741 B.n665 VSUBS 0.008543f
C742 B.n666 VSUBS 0.008543f
C743 B.n667 VSUBS 0.008543f
C744 B.n668 VSUBS 0.008543f
C745 B.n669 VSUBS 0.008543f
C746 B.n670 VSUBS 0.008543f
C747 B.n671 VSUBS 0.008543f
C748 B.n672 VSUBS 0.008543f
C749 B.n673 VSUBS 0.008543f
C750 B.n674 VSUBS 0.008543f
C751 B.n675 VSUBS 0.008543f
C752 B.n676 VSUBS 0.008543f
C753 B.n677 VSUBS 0.008543f
C754 B.n678 VSUBS 0.008543f
C755 B.n679 VSUBS 0.008543f
C756 B.n680 VSUBS 0.008543f
C757 B.n681 VSUBS 0.008543f
C758 B.n682 VSUBS 0.008543f
C759 B.n683 VSUBS 0.008543f
C760 B.n684 VSUBS 0.008543f
C761 B.n685 VSUBS 0.008543f
C762 B.n686 VSUBS 0.008543f
C763 B.n687 VSUBS 0.008543f
C764 B.n688 VSUBS 0.008543f
C765 B.n689 VSUBS 0.008543f
C766 B.n690 VSUBS 0.008543f
C767 B.n691 VSUBS 0.008543f
C768 B.n692 VSUBS 0.008543f
C769 B.n693 VSUBS 0.008543f
C770 B.n694 VSUBS 0.008543f
C771 B.n695 VSUBS 0.008543f
C772 B.n696 VSUBS 0.008543f
C773 B.n697 VSUBS 0.008543f
C774 B.n698 VSUBS 0.008543f
C775 B.n699 VSUBS 0.019345f
C776 VDD1.t5 VSUBS 3.80457f
C777 VDD1.t3 VSUBS 3.80335f
C778 VDD1.t4 VSUBS 0.355006f
C779 VDD1.t0 VSUBS 0.355006f
C780 VDD1.n0 VSUBS 2.92457f
C781 VDD1.n1 VSUBS 3.5198f
C782 VDD1.t2 VSUBS 0.355006f
C783 VDD1.t1 VSUBS 0.355006f
C784 VDD1.n2 VSUBS 2.92198f
C785 VDD1.n3 VSUBS 3.27893f
C786 VTAIL.t4 VSUBS 0.359541f
C787 VTAIL.t3 VSUBS 0.359541f
C788 VTAIL.n0 VSUBS 2.79688f
C789 VTAIL.n1 VSUBS 0.790561f
C790 VTAIL.t9 VSUBS 3.6573f
C791 VTAIL.n2 VSUBS 0.992275f
C792 VTAIL.t7 VSUBS 0.359541f
C793 VTAIL.t6 VSUBS 0.359541f
C794 VTAIL.n3 VSUBS 2.79688f
C795 VTAIL.n4 VSUBS 2.64229f
C796 VTAIL.t1 VSUBS 0.359541f
C797 VTAIL.t0 VSUBS 0.359541f
C798 VTAIL.n5 VSUBS 2.79688f
C799 VTAIL.n6 VSUBS 2.64229f
C800 VTAIL.t2 VSUBS 3.65731f
C801 VTAIL.n7 VSUBS 0.992269f
C802 VTAIL.t10 VSUBS 0.359541f
C803 VTAIL.t8 VSUBS 0.359541f
C804 VTAIL.n8 VSUBS 2.79688f
C805 VTAIL.n9 VSUBS 0.87213f
C806 VTAIL.t11 VSUBS 3.6573f
C807 VTAIL.n10 VSUBS 2.64677f
C808 VTAIL.t5 VSUBS 3.6573f
C809 VTAIL.n11 VSUBS 2.61269f
C810 VP.n0 VSUBS 0.044048f
C811 VP.t5 VSUBS 2.35491f
C812 VP.n1 VSUBS 0.067134f
C813 VP.n2 VSUBS 0.044048f
C814 VP.t2 VSUBS 2.35491f
C815 VP.n3 VSUBS 0.913085f
C816 VP.n4 VSUBS 0.044048f
C817 VP.t4 VSUBS 2.35491f
C818 VP.n5 VSUBS 0.067134f
C819 VP.t0 VSUBS 2.43538f
C820 VP.t3 VSUBS 2.35491f
C821 VP.n6 VSUBS 0.905873f
C822 VP.n7 VSUBS 0.94065f
C823 VP.n8 VSUBS 0.228717f
C824 VP.n9 VSUBS 0.044048f
C825 VP.n10 VSUBS 0.03559f
C826 VP.n11 VSUBS 0.067503f
C827 VP.n12 VSUBS 0.913085f
C828 VP.n13 VSUBS 2.14105f
C829 VP.n14 VSUBS 2.17527f
C830 VP.n15 VSUBS 0.044048f
C831 VP.n16 VSUBS 0.067503f
C832 VP.n17 VSUBS 0.03559f
C833 VP.t1 VSUBS 2.35491f
C834 VP.n18 VSUBS 0.84148f
C835 VP.n19 VSUBS 0.067134f
C836 VP.n20 VSUBS 0.044048f
C837 VP.n21 VSUBS 0.044048f
C838 VP.n22 VSUBS 0.044048f
C839 VP.n23 VSUBS 0.03559f
C840 VP.n24 VSUBS 0.067503f
C841 VP.n25 VSUBS 0.913085f
C842 VP.n26 VSUBS 0.039376f
.ends

