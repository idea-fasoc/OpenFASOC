* NGSPICE file created from diff_pair_sample_0839.ext - technology: sky130A

.subckt diff_pair_sample_0839 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.51
X1 VDD2.t9 VN.t0 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=7.1565 ps=37.48 w=18.35 l=1.51
X2 VTAIL.t11 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X3 VDD1.t9 VP.t0 VTAIL.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X4 VDD2.t7 VN.t2 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X5 VTAIL.t10 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X6 VTAIL.t5 VP.t1 VDD1.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X7 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.51
X8 VTAIL.t18 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X9 VDD2.t4 VN.t5 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=3.02775 ps=18.68 w=18.35 l=1.51
X10 VTAIL.t1 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X11 VDD2.t3 VN.t6 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=3.02775 ps=18.68 w=18.35 l=1.51
X12 VDD1.t6 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=3.02775 ps=18.68 w=18.35 l=1.51
X13 VTAIL.t3 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X14 VDD1.t4 VP.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=7.1565 ps=37.48 w=18.35 l=1.51
X15 VDD2.t2 VN.t7 VTAIL.t19 B.t6 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=7.1565 ps=37.48 w=18.35 l=1.51
X16 VDD1.t3 VP.t6 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X17 VDD2.t1 VN.t8 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.51
X19 VTAIL.t6 VP.t7 VDD1.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X20 VTAIL.t16 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=3.02775 ps=18.68 w=18.35 l=1.51
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.51
X22 VDD1.t1 VP.t8 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=3.02775 pd=18.68 as=7.1565 ps=37.48 w=18.35 l=1.51
X23 VDD1.t0 VP.t9 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=3.02775 ps=18.68 w=18.35 l=1.51
R0 B.n985 B.n984 585
R1 B.n401 B.n140 585
R2 B.n400 B.n399 585
R3 B.n398 B.n397 585
R4 B.n396 B.n395 585
R5 B.n394 B.n393 585
R6 B.n392 B.n391 585
R7 B.n390 B.n389 585
R8 B.n388 B.n387 585
R9 B.n386 B.n385 585
R10 B.n384 B.n383 585
R11 B.n382 B.n381 585
R12 B.n380 B.n379 585
R13 B.n378 B.n377 585
R14 B.n376 B.n375 585
R15 B.n374 B.n373 585
R16 B.n372 B.n371 585
R17 B.n370 B.n369 585
R18 B.n368 B.n367 585
R19 B.n366 B.n365 585
R20 B.n364 B.n363 585
R21 B.n362 B.n361 585
R22 B.n360 B.n359 585
R23 B.n358 B.n357 585
R24 B.n356 B.n355 585
R25 B.n354 B.n353 585
R26 B.n352 B.n351 585
R27 B.n350 B.n349 585
R28 B.n348 B.n347 585
R29 B.n346 B.n345 585
R30 B.n344 B.n343 585
R31 B.n342 B.n341 585
R32 B.n340 B.n339 585
R33 B.n338 B.n337 585
R34 B.n336 B.n335 585
R35 B.n334 B.n333 585
R36 B.n332 B.n331 585
R37 B.n330 B.n329 585
R38 B.n328 B.n327 585
R39 B.n326 B.n325 585
R40 B.n324 B.n323 585
R41 B.n322 B.n321 585
R42 B.n320 B.n319 585
R43 B.n318 B.n317 585
R44 B.n316 B.n315 585
R45 B.n314 B.n313 585
R46 B.n312 B.n311 585
R47 B.n310 B.n309 585
R48 B.n308 B.n307 585
R49 B.n306 B.n305 585
R50 B.n304 B.n303 585
R51 B.n302 B.n301 585
R52 B.n300 B.n299 585
R53 B.n298 B.n297 585
R54 B.n296 B.n295 585
R55 B.n294 B.n293 585
R56 B.n292 B.n291 585
R57 B.n290 B.n289 585
R58 B.n288 B.n287 585
R59 B.n286 B.n285 585
R60 B.n284 B.n283 585
R61 B.n282 B.n281 585
R62 B.n280 B.n279 585
R63 B.n278 B.n277 585
R64 B.n276 B.n275 585
R65 B.n274 B.n273 585
R66 B.n272 B.n271 585
R67 B.n270 B.n269 585
R68 B.n268 B.n267 585
R69 B.n266 B.n265 585
R70 B.n264 B.n263 585
R71 B.n262 B.n261 585
R72 B.n260 B.n259 585
R73 B.n258 B.n257 585
R74 B.n256 B.n255 585
R75 B.n254 B.n253 585
R76 B.n252 B.n251 585
R77 B.n250 B.n249 585
R78 B.n248 B.n247 585
R79 B.n246 B.n245 585
R80 B.n244 B.n243 585
R81 B.n242 B.n241 585
R82 B.n240 B.n239 585
R83 B.n238 B.n237 585
R84 B.n236 B.n235 585
R85 B.n234 B.n233 585
R86 B.n232 B.n231 585
R87 B.n230 B.n229 585
R88 B.n228 B.n227 585
R89 B.n226 B.n225 585
R90 B.n224 B.n223 585
R91 B.n222 B.n221 585
R92 B.n220 B.n219 585
R93 B.n218 B.n217 585
R94 B.n216 B.n215 585
R95 B.n214 B.n213 585
R96 B.n212 B.n211 585
R97 B.n210 B.n209 585
R98 B.n208 B.n207 585
R99 B.n206 B.n205 585
R100 B.n204 B.n203 585
R101 B.n202 B.n201 585
R102 B.n200 B.n199 585
R103 B.n198 B.n197 585
R104 B.n196 B.n195 585
R105 B.n194 B.n193 585
R106 B.n192 B.n191 585
R107 B.n190 B.n189 585
R108 B.n188 B.n187 585
R109 B.n186 B.n185 585
R110 B.n184 B.n183 585
R111 B.n182 B.n181 585
R112 B.n180 B.n179 585
R113 B.n178 B.n177 585
R114 B.n176 B.n175 585
R115 B.n174 B.n173 585
R116 B.n172 B.n171 585
R117 B.n170 B.n169 585
R118 B.n168 B.n167 585
R119 B.n166 B.n165 585
R120 B.n164 B.n163 585
R121 B.n162 B.n161 585
R122 B.n160 B.n159 585
R123 B.n158 B.n157 585
R124 B.n156 B.n155 585
R125 B.n154 B.n153 585
R126 B.n152 B.n151 585
R127 B.n150 B.n149 585
R128 B.n148 B.n147 585
R129 B.n74 B.n73 585
R130 B.n983 B.n75 585
R131 B.n988 B.n75 585
R132 B.n982 B.n981 585
R133 B.n981 B.n71 585
R134 B.n980 B.n70 585
R135 B.n994 B.n70 585
R136 B.n979 B.n69 585
R137 B.n995 B.n69 585
R138 B.n978 B.n68 585
R139 B.n996 B.n68 585
R140 B.n977 B.n976 585
R141 B.n976 B.n67 585
R142 B.n975 B.n63 585
R143 B.n1002 B.n63 585
R144 B.n974 B.n62 585
R145 B.n1003 B.n62 585
R146 B.n973 B.n61 585
R147 B.n1004 B.n61 585
R148 B.n972 B.n971 585
R149 B.n971 B.n57 585
R150 B.n970 B.n56 585
R151 B.n1010 B.n56 585
R152 B.n969 B.n55 585
R153 B.n1011 B.n55 585
R154 B.n968 B.n54 585
R155 B.n1012 B.n54 585
R156 B.n967 B.n966 585
R157 B.n966 B.n50 585
R158 B.n965 B.n49 585
R159 B.n1018 B.n49 585
R160 B.n964 B.n48 585
R161 B.n1019 B.n48 585
R162 B.n963 B.n47 585
R163 B.n1020 B.n47 585
R164 B.n962 B.n961 585
R165 B.n961 B.n43 585
R166 B.n960 B.n42 585
R167 B.n1026 B.n42 585
R168 B.n959 B.n41 585
R169 B.n1027 B.n41 585
R170 B.n958 B.n40 585
R171 B.n1028 B.n40 585
R172 B.n957 B.n956 585
R173 B.n956 B.n36 585
R174 B.n955 B.n35 585
R175 B.n1034 B.n35 585
R176 B.n954 B.n34 585
R177 B.n1035 B.n34 585
R178 B.n953 B.n33 585
R179 B.n1036 B.n33 585
R180 B.n952 B.n951 585
R181 B.n951 B.n32 585
R182 B.n950 B.n28 585
R183 B.n1042 B.n28 585
R184 B.n949 B.n27 585
R185 B.n1043 B.n27 585
R186 B.n948 B.n26 585
R187 B.n1044 B.n26 585
R188 B.n947 B.n946 585
R189 B.n946 B.n22 585
R190 B.n945 B.n21 585
R191 B.n1050 B.n21 585
R192 B.n944 B.n20 585
R193 B.n1051 B.n20 585
R194 B.n943 B.n19 585
R195 B.n1052 B.n19 585
R196 B.n942 B.n941 585
R197 B.n941 B.n15 585
R198 B.n940 B.n14 585
R199 B.n1058 B.n14 585
R200 B.n939 B.n13 585
R201 B.n1059 B.n13 585
R202 B.n938 B.n12 585
R203 B.n1060 B.n12 585
R204 B.n937 B.n936 585
R205 B.n936 B.n935 585
R206 B.n934 B.n933 585
R207 B.n934 B.n8 585
R208 B.n932 B.n7 585
R209 B.n1067 B.n7 585
R210 B.n931 B.n6 585
R211 B.n1068 B.n6 585
R212 B.n930 B.n5 585
R213 B.n1069 B.n5 585
R214 B.n929 B.n928 585
R215 B.n928 B.n4 585
R216 B.n927 B.n402 585
R217 B.n927 B.n926 585
R218 B.n917 B.n403 585
R219 B.n404 B.n403 585
R220 B.n919 B.n918 585
R221 B.n920 B.n919 585
R222 B.n916 B.n409 585
R223 B.n409 B.n408 585
R224 B.n915 B.n914 585
R225 B.n914 B.n913 585
R226 B.n411 B.n410 585
R227 B.n412 B.n411 585
R228 B.n906 B.n905 585
R229 B.n907 B.n906 585
R230 B.n904 B.n417 585
R231 B.n417 B.n416 585
R232 B.n903 B.n902 585
R233 B.n902 B.n901 585
R234 B.n419 B.n418 585
R235 B.n420 B.n419 585
R236 B.n894 B.n893 585
R237 B.n895 B.n894 585
R238 B.n892 B.n425 585
R239 B.n425 B.n424 585
R240 B.n891 B.n890 585
R241 B.n890 B.n889 585
R242 B.n427 B.n426 585
R243 B.n882 B.n427 585
R244 B.n881 B.n880 585
R245 B.n883 B.n881 585
R246 B.n879 B.n432 585
R247 B.n432 B.n431 585
R248 B.n878 B.n877 585
R249 B.n877 B.n876 585
R250 B.n434 B.n433 585
R251 B.n435 B.n434 585
R252 B.n869 B.n868 585
R253 B.n870 B.n869 585
R254 B.n867 B.n439 585
R255 B.n443 B.n439 585
R256 B.n866 B.n865 585
R257 B.n865 B.n864 585
R258 B.n441 B.n440 585
R259 B.n442 B.n441 585
R260 B.n857 B.n856 585
R261 B.n858 B.n857 585
R262 B.n855 B.n448 585
R263 B.n448 B.n447 585
R264 B.n854 B.n853 585
R265 B.n853 B.n852 585
R266 B.n450 B.n449 585
R267 B.n451 B.n450 585
R268 B.n845 B.n844 585
R269 B.n846 B.n845 585
R270 B.n843 B.n456 585
R271 B.n456 B.n455 585
R272 B.n842 B.n841 585
R273 B.n841 B.n840 585
R274 B.n458 B.n457 585
R275 B.n459 B.n458 585
R276 B.n833 B.n832 585
R277 B.n834 B.n833 585
R278 B.n831 B.n464 585
R279 B.n464 B.n463 585
R280 B.n830 B.n829 585
R281 B.n829 B.n828 585
R282 B.n466 B.n465 585
R283 B.n821 B.n466 585
R284 B.n820 B.n819 585
R285 B.n822 B.n820 585
R286 B.n818 B.n471 585
R287 B.n471 B.n470 585
R288 B.n817 B.n816 585
R289 B.n816 B.n815 585
R290 B.n473 B.n472 585
R291 B.n474 B.n473 585
R292 B.n808 B.n807 585
R293 B.n809 B.n808 585
R294 B.n477 B.n476 585
R295 B.n548 B.n546 585
R296 B.n549 B.n545 585
R297 B.n549 B.n478 585
R298 B.n552 B.n551 585
R299 B.n553 B.n544 585
R300 B.n555 B.n554 585
R301 B.n557 B.n543 585
R302 B.n560 B.n559 585
R303 B.n561 B.n542 585
R304 B.n563 B.n562 585
R305 B.n565 B.n541 585
R306 B.n568 B.n567 585
R307 B.n569 B.n540 585
R308 B.n571 B.n570 585
R309 B.n573 B.n539 585
R310 B.n576 B.n575 585
R311 B.n577 B.n538 585
R312 B.n579 B.n578 585
R313 B.n581 B.n537 585
R314 B.n584 B.n583 585
R315 B.n585 B.n536 585
R316 B.n587 B.n586 585
R317 B.n589 B.n535 585
R318 B.n592 B.n591 585
R319 B.n593 B.n534 585
R320 B.n595 B.n594 585
R321 B.n597 B.n533 585
R322 B.n600 B.n599 585
R323 B.n601 B.n532 585
R324 B.n603 B.n602 585
R325 B.n605 B.n531 585
R326 B.n608 B.n607 585
R327 B.n609 B.n530 585
R328 B.n611 B.n610 585
R329 B.n613 B.n529 585
R330 B.n616 B.n615 585
R331 B.n617 B.n528 585
R332 B.n619 B.n618 585
R333 B.n621 B.n527 585
R334 B.n624 B.n623 585
R335 B.n625 B.n526 585
R336 B.n627 B.n626 585
R337 B.n629 B.n525 585
R338 B.n632 B.n631 585
R339 B.n633 B.n524 585
R340 B.n635 B.n634 585
R341 B.n637 B.n523 585
R342 B.n640 B.n639 585
R343 B.n641 B.n522 585
R344 B.n643 B.n642 585
R345 B.n645 B.n521 585
R346 B.n648 B.n647 585
R347 B.n649 B.n520 585
R348 B.n651 B.n650 585
R349 B.n653 B.n519 585
R350 B.n656 B.n655 585
R351 B.n657 B.n518 585
R352 B.n659 B.n658 585
R353 B.n661 B.n517 585
R354 B.n664 B.n663 585
R355 B.n666 B.n514 585
R356 B.n668 B.n667 585
R357 B.n670 B.n513 585
R358 B.n673 B.n672 585
R359 B.n674 B.n512 585
R360 B.n676 B.n675 585
R361 B.n678 B.n511 585
R362 B.n681 B.n680 585
R363 B.n682 B.n510 585
R364 B.n687 B.n686 585
R365 B.n689 B.n509 585
R366 B.n692 B.n691 585
R367 B.n693 B.n508 585
R368 B.n695 B.n694 585
R369 B.n697 B.n507 585
R370 B.n700 B.n699 585
R371 B.n701 B.n506 585
R372 B.n703 B.n702 585
R373 B.n705 B.n505 585
R374 B.n708 B.n707 585
R375 B.n709 B.n504 585
R376 B.n711 B.n710 585
R377 B.n713 B.n503 585
R378 B.n716 B.n715 585
R379 B.n717 B.n502 585
R380 B.n719 B.n718 585
R381 B.n721 B.n501 585
R382 B.n724 B.n723 585
R383 B.n725 B.n500 585
R384 B.n727 B.n726 585
R385 B.n729 B.n499 585
R386 B.n732 B.n731 585
R387 B.n733 B.n498 585
R388 B.n735 B.n734 585
R389 B.n737 B.n497 585
R390 B.n740 B.n739 585
R391 B.n741 B.n496 585
R392 B.n743 B.n742 585
R393 B.n745 B.n495 585
R394 B.n748 B.n747 585
R395 B.n749 B.n494 585
R396 B.n751 B.n750 585
R397 B.n753 B.n493 585
R398 B.n756 B.n755 585
R399 B.n757 B.n492 585
R400 B.n759 B.n758 585
R401 B.n761 B.n491 585
R402 B.n764 B.n763 585
R403 B.n765 B.n490 585
R404 B.n767 B.n766 585
R405 B.n769 B.n489 585
R406 B.n772 B.n771 585
R407 B.n773 B.n488 585
R408 B.n775 B.n774 585
R409 B.n777 B.n487 585
R410 B.n780 B.n779 585
R411 B.n781 B.n486 585
R412 B.n783 B.n782 585
R413 B.n785 B.n485 585
R414 B.n788 B.n787 585
R415 B.n789 B.n484 585
R416 B.n791 B.n790 585
R417 B.n793 B.n483 585
R418 B.n796 B.n795 585
R419 B.n797 B.n482 585
R420 B.n799 B.n798 585
R421 B.n801 B.n481 585
R422 B.n802 B.n480 585
R423 B.n805 B.n804 585
R424 B.n806 B.n479 585
R425 B.n479 B.n478 585
R426 B.n811 B.n810 585
R427 B.n810 B.n809 585
R428 B.n812 B.n475 585
R429 B.n475 B.n474 585
R430 B.n814 B.n813 585
R431 B.n815 B.n814 585
R432 B.n469 B.n468 585
R433 B.n470 B.n469 585
R434 B.n824 B.n823 585
R435 B.n823 B.n822 585
R436 B.n825 B.n467 585
R437 B.n821 B.n467 585
R438 B.n827 B.n826 585
R439 B.n828 B.n827 585
R440 B.n462 B.n461 585
R441 B.n463 B.n462 585
R442 B.n836 B.n835 585
R443 B.n835 B.n834 585
R444 B.n837 B.n460 585
R445 B.n460 B.n459 585
R446 B.n839 B.n838 585
R447 B.n840 B.n839 585
R448 B.n454 B.n453 585
R449 B.n455 B.n454 585
R450 B.n848 B.n847 585
R451 B.n847 B.n846 585
R452 B.n849 B.n452 585
R453 B.n452 B.n451 585
R454 B.n851 B.n850 585
R455 B.n852 B.n851 585
R456 B.n446 B.n445 585
R457 B.n447 B.n446 585
R458 B.n860 B.n859 585
R459 B.n859 B.n858 585
R460 B.n861 B.n444 585
R461 B.n444 B.n442 585
R462 B.n863 B.n862 585
R463 B.n864 B.n863 585
R464 B.n438 B.n437 585
R465 B.n443 B.n438 585
R466 B.n872 B.n871 585
R467 B.n871 B.n870 585
R468 B.n873 B.n436 585
R469 B.n436 B.n435 585
R470 B.n875 B.n874 585
R471 B.n876 B.n875 585
R472 B.n430 B.n429 585
R473 B.n431 B.n430 585
R474 B.n885 B.n884 585
R475 B.n884 B.n883 585
R476 B.n886 B.n428 585
R477 B.n882 B.n428 585
R478 B.n888 B.n887 585
R479 B.n889 B.n888 585
R480 B.n423 B.n422 585
R481 B.n424 B.n423 585
R482 B.n897 B.n896 585
R483 B.n896 B.n895 585
R484 B.n898 B.n421 585
R485 B.n421 B.n420 585
R486 B.n900 B.n899 585
R487 B.n901 B.n900 585
R488 B.n415 B.n414 585
R489 B.n416 B.n415 585
R490 B.n909 B.n908 585
R491 B.n908 B.n907 585
R492 B.n910 B.n413 585
R493 B.n413 B.n412 585
R494 B.n912 B.n911 585
R495 B.n913 B.n912 585
R496 B.n407 B.n406 585
R497 B.n408 B.n407 585
R498 B.n922 B.n921 585
R499 B.n921 B.n920 585
R500 B.n923 B.n405 585
R501 B.n405 B.n404 585
R502 B.n925 B.n924 585
R503 B.n926 B.n925 585
R504 B.n3 B.n0 585
R505 B.n4 B.n3 585
R506 B.n1066 B.n1 585
R507 B.n1067 B.n1066 585
R508 B.n1065 B.n1064 585
R509 B.n1065 B.n8 585
R510 B.n1063 B.n9 585
R511 B.n935 B.n9 585
R512 B.n1062 B.n1061 585
R513 B.n1061 B.n1060 585
R514 B.n11 B.n10 585
R515 B.n1059 B.n11 585
R516 B.n1057 B.n1056 585
R517 B.n1058 B.n1057 585
R518 B.n1055 B.n16 585
R519 B.n16 B.n15 585
R520 B.n1054 B.n1053 585
R521 B.n1053 B.n1052 585
R522 B.n18 B.n17 585
R523 B.n1051 B.n18 585
R524 B.n1049 B.n1048 585
R525 B.n1050 B.n1049 585
R526 B.n1047 B.n23 585
R527 B.n23 B.n22 585
R528 B.n1046 B.n1045 585
R529 B.n1045 B.n1044 585
R530 B.n25 B.n24 585
R531 B.n1043 B.n25 585
R532 B.n1041 B.n1040 585
R533 B.n1042 B.n1041 585
R534 B.n1039 B.n29 585
R535 B.n32 B.n29 585
R536 B.n1038 B.n1037 585
R537 B.n1037 B.n1036 585
R538 B.n31 B.n30 585
R539 B.n1035 B.n31 585
R540 B.n1033 B.n1032 585
R541 B.n1034 B.n1033 585
R542 B.n1031 B.n37 585
R543 B.n37 B.n36 585
R544 B.n1030 B.n1029 585
R545 B.n1029 B.n1028 585
R546 B.n39 B.n38 585
R547 B.n1027 B.n39 585
R548 B.n1025 B.n1024 585
R549 B.n1026 B.n1025 585
R550 B.n1023 B.n44 585
R551 B.n44 B.n43 585
R552 B.n1022 B.n1021 585
R553 B.n1021 B.n1020 585
R554 B.n46 B.n45 585
R555 B.n1019 B.n46 585
R556 B.n1017 B.n1016 585
R557 B.n1018 B.n1017 585
R558 B.n1015 B.n51 585
R559 B.n51 B.n50 585
R560 B.n1014 B.n1013 585
R561 B.n1013 B.n1012 585
R562 B.n53 B.n52 585
R563 B.n1011 B.n53 585
R564 B.n1009 B.n1008 585
R565 B.n1010 B.n1009 585
R566 B.n1007 B.n58 585
R567 B.n58 B.n57 585
R568 B.n1006 B.n1005 585
R569 B.n1005 B.n1004 585
R570 B.n60 B.n59 585
R571 B.n1003 B.n60 585
R572 B.n1001 B.n1000 585
R573 B.n1002 B.n1001 585
R574 B.n999 B.n64 585
R575 B.n67 B.n64 585
R576 B.n998 B.n997 585
R577 B.n997 B.n996 585
R578 B.n66 B.n65 585
R579 B.n995 B.n66 585
R580 B.n993 B.n992 585
R581 B.n994 B.n993 585
R582 B.n991 B.n72 585
R583 B.n72 B.n71 585
R584 B.n990 B.n989 585
R585 B.n989 B.n988 585
R586 B.n1070 B.n1069 585
R587 B.n1068 B.n2 585
R588 B.n989 B.n74 526.135
R589 B.n985 B.n75 526.135
R590 B.n808 B.n479 526.135
R591 B.n810 B.n477 526.135
R592 B.n144 B.t21 498.349
R593 B.n141 B.t14 498.349
R594 B.n683 B.t18 498.349
R595 B.n515 B.t10 498.349
R596 B.n141 B.t16 427.565
R597 B.n683 B.t20 427.565
R598 B.n144 B.t22 427.565
R599 B.n515 B.t13 427.565
R600 B.n142 B.t17 391.88
R601 B.n684 B.t19 391.88
R602 B.n145 B.t23 391.88
R603 B.n516 B.t12 391.88
R604 B.n987 B.n986 256.663
R605 B.n987 B.n139 256.663
R606 B.n987 B.n138 256.663
R607 B.n987 B.n137 256.663
R608 B.n987 B.n136 256.663
R609 B.n987 B.n135 256.663
R610 B.n987 B.n134 256.663
R611 B.n987 B.n133 256.663
R612 B.n987 B.n132 256.663
R613 B.n987 B.n131 256.663
R614 B.n987 B.n130 256.663
R615 B.n987 B.n129 256.663
R616 B.n987 B.n128 256.663
R617 B.n987 B.n127 256.663
R618 B.n987 B.n126 256.663
R619 B.n987 B.n125 256.663
R620 B.n987 B.n124 256.663
R621 B.n987 B.n123 256.663
R622 B.n987 B.n122 256.663
R623 B.n987 B.n121 256.663
R624 B.n987 B.n120 256.663
R625 B.n987 B.n119 256.663
R626 B.n987 B.n118 256.663
R627 B.n987 B.n117 256.663
R628 B.n987 B.n116 256.663
R629 B.n987 B.n115 256.663
R630 B.n987 B.n114 256.663
R631 B.n987 B.n113 256.663
R632 B.n987 B.n112 256.663
R633 B.n987 B.n111 256.663
R634 B.n987 B.n110 256.663
R635 B.n987 B.n109 256.663
R636 B.n987 B.n108 256.663
R637 B.n987 B.n107 256.663
R638 B.n987 B.n106 256.663
R639 B.n987 B.n105 256.663
R640 B.n987 B.n104 256.663
R641 B.n987 B.n103 256.663
R642 B.n987 B.n102 256.663
R643 B.n987 B.n101 256.663
R644 B.n987 B.n100 256.663
R645 B.n987 B.n99 256.663
R646 B.n987 B.n98 256.663
R647 B.n987 B.n97 256.663
R648 B.n987 B.n96 256.663
R649 B.n987 B.n95 256.663
R650 B.n987 B.n94 256.663
R651 B.n987 B.n93 256.663
R652 B.n987 B.n92 256.663
R653 B.n987 B.n91 256.663
R654 B.n987 B.n90 256.663
R655 B.n987 B.n89 256.663
R656 B.n987 B.n88 256.663
R657 B.n987 B.n87 256.663
R658 B.n987 B.n86 256.663
R659 B.n987 B.n85 256.663
R660 B.n987 B.n84 256.663
R661 B.n987 B.n83 256.663
R662 B.n987 B.n82 256.663
R663 B.n987 B.n81 256.663
R664 B.n987 B.n80 256.663
R665 B.n987 B.n79 256.663
R666 B.n987 B.n78 256.663
R667 B.n987 B.n77 256.663
R668 B.n987 B.n76 256.663
R669 B.n547 B.n478 256.663
R670 B.n550 B.n478 256.663
R671 B.n556 B.n478 256.663
R672 B.n558 B.n478 256.663
R673 B.n564 B.n478 256.663
R674 B.n566 B.n478 256.663
R675 B.n572 B.n478 256.663
R676 B.n574 B.n478 256.663
R677 B.n580 B.n478 256.663
R678 B.n582 B.n478 256.663
R679 B.n588 B.n478 256.663
R680 B.n590 B.n478 256.663
R681 B.n596 B.n478 256.663
R682 B.n598 B.n478 256.663
R683 B.n604 B.n478 256.663
R684 B.n606 B.n478 256.663
R685 B.n612 B.n478 256.663
R686 B.n614 B.n478 256.663
R687 B.n620 B.n478 256.663
R688 B.n622 B.n478 256.663
R689 B.n628 B.n478 256.663
R690 B.n630 B.n478 256.663
R691 B.n636 B.n478 256.663
R692 B.n638 B.n478 256.663
R693 B.n644 B.n478 256.663
R694 B.n646 B.n478 256.663
R695 B.n652 B.n478 256.663
R696 B.n654 B.n478 256.663
R697 B.n660 B.n478 256.663
R698 B.n662 B.n478 256.663
R699 B.n669 B.n478 256.663
R700 B.n671 B.n478 256.663
R701 B.n677 B.n478 256.663
R702 B.n679 B.n478 256.663
R703 B.n688 B.n478 256.663
R704 B.n690 B.n478 256.663
R705 B.n696 B.n478 256.663
R706 B.n698 B.n478 256.663
R707 B.n704 B.n478 256.663
R708 B.n706 B.n478 256.663
R709 B.n712 B.n478 256.663
R710 B.n714 B.n478 256.663
R711 B.n720 B.n478 256.663
R712 B.n722 B.n478 256.663
R713 B.n728 B.n478 256.663
R714 B.n730 B.n478 256.663
R715 B.n736 B.n478 256.663
R716 B.n738 B.n478 256.663
R717 B.n744 B.n478 256.663
R718 B.n746 B.n478 256.663
R719 B.n752 B.n478 256.663
R720 B.n754 B.n478 256.663
R721 B.n760 B.n478 256.663
R722 B.n762 B.n478 256.663
R723 B.n768 B.n478 256.663
R724 B.n770 B.n478 256.663
R725 B.n776 B.n478 256.663
R726 B.n778 B.n478 256.663
R727 B.n784 B.n478 256.663
R728 B.n786 B.n478 256.663
R729 B.n792 B.n478 256.663
R730 B.n794 B.n478 256.663
R731 B.n800 B.n478 256.663
R732 B.n803 B.n478 256.663
R733 B.n1072 B.n1071 256.663
R734 B.n149 B.n148 163.367
R735 B.n153 B.n152 163.367
R736 B.n157 B.n156 163.367
R737 B.n161 B.n160 163.367
R738 B.n165 B.n164 163.367
R739 B.n169 B.n168 163.367
R740 B.n173 B.n172 163.367
R741 B.n177 B.n176 163.367
R742 B.n181 B.n180 163.367
R743 B.n185 B.n184 163.367
R744 B.n189 B.n188 163.367
R745 B.n193 B.n192 163.367
R746 B.n197 B.n196 163.367
R747 B.n201 B.n200 163.367
R748 B.n205 B.n204 163.367
R749 B.n209 B.n208 163.367
R750 B.n213 B.n212 163.367
R751 B.n217 B.n216 163.367
R752 B.n221 B.n220 163.367
R753 B.n225 B.n224 163.367
R754 B.n229 B.n228 163.367
R755 B.n233 B.n232 163.367
R756 B.n237 B.n236 163.367
R757 B.n241 B.n240 163.367
R758 B.n245 B.n244 163.367
R759 B.n249 B.n248 163.367
R760 B.n253 B.n252 163.367
R761 B.n257 B.n256 163.367
R762 B.n261 B.n260 163.367
R763 B.n265 B.n264 163.367
R764 B.n269 B.n268 163.367
R765 B.n273 B.n272 163.367
R766 B.n277 B.n276 163.367
R767 B.n281 B.n280 163.367
R768 B.n285 B.n284 163.367
R769 B.n289 B.n288 163.367
R770 B.n293 B.n292 163.367
R771 B.n297 B.n296 163.367
R772 B.n301 B.n300 163.367
R773 B.n305 B.n304 163.367
R774 B.n309 B.n308 163.367
R775 B.n313 B.n312 163.367
R776 B.n317 B.n316 163.367
R777 B.n321 B.n320 163.367
R778 B.n325 B.n324 163.367
R779 B.n329 B.n328 163.367
R780 B.n333 B.n332 163.367
R781 B.n337 B.n336 163.367
R782 B.n341 B.n340 163.367
R783 B.n345 B.n344 163.367
R784 B.n349 B.n348 163.367
R785 B.n353 B.n352 163.367
R786 B.n357 B.n356 163.367
R787 B.n361 B.n360 163.367
R788 B.n365 B.n364 163.367
R789 B.n369 B.n368 163.367
R790 B.n373 B.n372 163.367
R791 B.n377 B.n376 163.367
R792 B.n381 B.n380 163.367
R793 B.n385 B.n384 163.367
R794 B.n389 B.n388 163.367
R795 B.n393 B.n392 163.367
R796 B.n397 B.n396 163.367
R797 B.n399 B.n140 163.367
R798 B.n808 B.n473 163.367
R799 B.n816 B.n473 163.367
R800 B.n816 B.n471 163.367
R801 B.n820 B.n471 163.367
R802 B.n820 B.n466 163.367
R803 B.n829 B.n466 163.367
R804 B.n829 B.n464 163.367
R805 B.n833 B.n464 163.367
R806 B.n833 B.n458 163.367
R807 B.n841 B.n458 163.367
R808 B.n841 B.n456 163.367
R809 B.n845 B.n456 163.367
R810 B.n845 B.n450 163.367
R811 B.n853 B.n450 163.367
R812 B.n853 B.n448 163.367
R813 B.n857 B.n448 163.367
R814 B.n857 B.n441 163.367
R815 B.n865 B.n441 163.367
R816 B.n865 B.n439 163.367
R817 B.n869 B.n439 163.367
R818 B.n869 B.n434 163.367
R819 B.n877 B.n434 163.367
R820 B.n877 B.n432 163.367
R821 B.n881 B.n432 163.367
R822 B.n881 B.n427 163.367
R823 B.n890 B.n427 163.367
R824 B.n890 B.n425 163.367
R825 B.n894 B.n425 163.367
R826 B.n894 B.n419 163.367
R827 B.n902 B.n419 163.367
R828 B.n902 B.n417 163.367
R829 B.n906 B.n417 163.367
R830 B.n906 B.n411 163.367
R831 B.n914 B.n411 163.367
R832 B.n914 B.n409 163.367
R833 B.n919 B.n409 163.367
R834 B.n919 B.n403 163.367
R835 B.n927 B.n403 163.367
R836 B.n928 B.n927 163.367
R837 B.n928 B.n5 163.367
R838 B.n6 B.n5 163.367
R839 B.n7 B.n6 163.367
R840 B.n934 B.n7 163.367
R841 B.n936 B.n934 163.367
R842 B.n936 B.n12 163.367
R843 B.n13 B.n12 163.367
R844 B.n14 B.n13 163.367
R845 B.n941 B.n14 163.367
R846 B.n941 B.n19 163.367
R847 B.n20 B.n19 163.367
R848 B.n21 B.n20 163.367
R849 B.n946 B.n21 163.367
R850 B.n946 B.n26 163.367
R851 B.n27 B.n26 163.367
R852 B.n28 B.n27 163.367
R853 B.n951 B.n28 163.367
R854 B.n951 B.n33 163.367
R855 B.n34 B.n33 163.367
R856 B.n35 B.n34 163.367
R857 B.n956 B.n35 163.367
R858 B.n956 B.n40 163.367
R859 B.n41 B.n40 163.367
R860 B.n42 B.n41 163.367
R861 B.n961 B.n42 163.367
R862 B.n961 B.n47 163.367
R863 B.n48 B.n47 163.367
R864 B.n49 B.n48 163.367
R865 B.n966 B.n49 163.367
R866 B.n966 B.n54 163.367
R867 B.n55 B.n54 163.367
R868 B.n56 B.n55 163.367
R869 B.n971 B.n56 163.367
R870 B.n971 B.n61 163.367
R871 B.n62 B.n61 163.367
R872 B.n63 B.n62 163.367
R873 B.n976 B.n63 163.367
R874 B.n976 B.n68 163.367
R875 B.n69 B.n68 163.367
R876 B.n70 B.n69 163.367
R877 B.n981 B.n70 163.367
R878 B.n981 B.n75 163.367
R879 B.n549 B.n548 163.367
R880 B.n551 B.n549 163.367
R881 B.n555 B.n544 163.367
R882 B.n559 B.n557 163.367
R883 B.n563 B.n542 163.367
R884 B.n567 B.n565 163.367
R885 B.n571 B.n540 163.367
R886 B.n575 B.n573 163.367
R887 B.n579 B.n538 163.367
R888 B.n583 B.n581 163.367
R889 B.n587 B.n536 163.367
R890 B.n591 B.n589 163.367
R891 B.n595 B.n534 163.367
R892 B.n599 B.n597 163.367
R893 B.n603 B.n532 163.367
R894 B.n607 B.n605 163.367
R895 B.n611 B.n530 163.367
R896 B.n615 B.n613 163.367
R897 B.n619 B.n528 163.367
R898 B.n623 B.n621 163.367
R899 B.n627 B.n526 163.367
R900 B.n631 B.n629 163.367
R901 B.n635 B.n524 163.367
R902 B.n639 B.n637 163.367
R903 B.n643 B.n522 163.367
R904 B.n647 B.n645 163.367
R905 B.n651 B.n520 163.367
R906 B.n655 B.n653 163.367
R907 B.n659 B.n518 163.367
R908 B.n663 B.n661 163.367
R909 B.n668 B.n514 163.367
R910 B.n672 B.n670 163.367
R911 B.n676 B.n512 163.367
R912 B.n680 B.n678 163.367
R913 B.n687 B.n510 163.367
R914 B.n691 B.n689 163.367
R915 B.n695 B.n508 163.367
R916 B.n699 B.n697 163.367
R917 B.n703 B.n506 163.367
R918 B.n707 B.n705 163.367
R919 B.n711 B.n504 163.367
R920 B.n715 B.n713 163.367
R921 B.n719 B.n502 163.367
R922 B.n723 B.n721 163.367
R923 B.n727 B.n500 163.367
R924 B.n731 B.n729 163.367
R925 B.n735 B.n498 163.367
R926 B.n739 B.n737 163.367
R927 B.n743 B.n496 163.367
R928 B.n747 B.n745 163.367
R929 B.n751 B.n494 163.367
R930 B.n755 B.n753 163.367
R931 B.n759 B.n492 163.367
R932 B.n763 B.n761 163.367
R933 B.n767 B.n490 163.367
R934 B.n771 B.n769 163.367
R935 B.n775 B.n488 163.367
R936 B.n779 B.n777 163.367
R937 B.n783 B.n486 163.367
R938 B.n787 B.n785 163.367
R939 B.n791 B.n484 163.367
R940 B.n795 B.n793 163.367
R941 B.n799 B.n482 163.367
R942 B.n802 B.n801 163.367
R943 B.n804 B.n479 163.367
R944 B.n810 B.n475 163.367
R945 B.n814 B.n475 163.367
R946 B.n814 B.n469 163.367
R947 B.n823 B.n469 163.367
R948 B.n823 B.n467 163.367
R949 B.n827 B.n467 163.367
R950 B.n827 B.n462 163.367
R951 B.n835 B.n462 163.367
R952 B.n835 B.n460 163.367
R953 B.n839 B.n460 163.367
R954 B.n839 B.n454 163.367
R955 B.n847 B.n454 163.367
R956 B.n847 B.n452 163.367
R957 B.n851 B.n452 163.367
R958 B.n851 B.n446 163.367
R959 B.n859 B.n446 163.367
R960 B.n859 B.n444 163.367
R961 B.n863 B.n444 163.367
R962 B.n863 B.n438 163.367
R963 B.n871 B.n438 163.367
R964 B.n871 B.n436 163.367
R965 B.n875 B.n436 163.367
R966 B.n875 B.n430 163.367
R967 B.n884 B.n430 163.367
R968 B.n884 B.n428 163.367
R969 B.n888 B.n428 163.367
R970 B.n888 B.n423 163.367
R971 B.n896 B.n423 163.367
R972 B.n896 B.n421 163.367
R973 B.n900 B.n421 163.367
R974 B.n900 B.n415 163.367
R975 B.n908 B.n415 163.367
R976 B.n908 B.n413 163.367
R977 B.n912 B.n413 163.367
R978 B.n912 B.n407 163.367
R979 B.n921 B.n407 163.367
R980 B.n921 B.n405 163.367
R981 B.n925 B.n405 163.367
R982 B.n925 B.n3 163.367
R983 B.n1070 B.n3 163.367
R984 B.n1066 B.n2 163.367
R985 B.n1066 B.n1065 163.367
R986 B.n1065 B.n9 163.367
R987 B.n1061 B.n9 163.367
R988 B.n1061 B.n11 163.367
R989 B.n1057 B.n11 163.367
R990 B.n1057 B.n16 163.367
R991 B.n1053 B.n16 163.367
R992 B.n1053 B.n18 163.367
R993 B.n1049 B.n18 163.367
R994 B.n1049 B.n23 163.367
R995 B.n1045 B.n23 163.367
R996 B.n1045 B.n25 163.367
R997 B.n1041 B.n25 163.367
R998 B.n1041 B.n29 163.367
R999 B.n1037 B.n29 163.367
R1000 B.n1037 B.n31 163.367
R1001 B.n1033 B.n31 163.367
R1002 B.n1033 B.n37 163.367
R1003 B.n1029 B.n37 163.367
R1004 B.n1029 B.n39 163.367
R1005 B.n1025 B.n39 163.367
R1006 B.n1025 B.n44 163.367
R1007 B.n1021 B.n44 163.367
R1008 B.n1021 B.n46 163.367
R1009 B.n1017 B.n46 163.367
R1010 B.n1017 B.n51 163.367
R1011 B.n1013 B.n51 163.367
R1012 B.n1013 B.n53 163.367
R1013 B.n1009 B.n53 163.367
R1014 B.n1009 B.n58 163.367
R1015 B.n1005 B.n58 163.367
R1016 B.n1005 B.n60 163.367
R1017 B.n1001 B.n60 163.367
R1018 B.n1001 B.n64 163.367
R1019 B.n997 B.n64 163.367
R1020 B.n997 B.n66 163.367
R1021 B.n993 B.n66 163.367
R1022 B.n993 B.n72 163.367
R1023 B.n989 B.n72 163.367
R1024 B.n76 B.n74 71.676
R1025 B.n149 B.n77 71.676
R1026 B.n153 B.n78 71.676
R1027 B.n157 B.n79 71.676
R1028 B.n161 B.n80 71.676
R1029 B.n165 B.n81 71.676
R1030 B.n169 B.n82 71.676
R1031 B.n173 B.n83 71.676
R1032 B.n177 B.n84 71.676
R1033 B.n181 B.n85 71.676
R1034 B.n185 B.n86 71.676
R1035 B.n189 B.n87 71.676
R1036 B.n193 B.n88 71.676
R1037 B.n197 B.n89 71.676
R1038 B.n201 B.n90 71.676
R1039 B.n205 B.n91 71.676
R1040 B.n209 B.n92 71.676
R1041 B.n213 B.n93 71.676
R1042 B.n217 B.n94 71.676
R1043 B.n221 B.n95 71.676
R1044 B.n225 B.n96 71.676
R1045 B.n229 B.n97 71.676
R1046 B.n233 B.n98 71.676
R1047 B.n237 B.n99 71.676
R1048 B.n241 B.n100 71.676
R1049 B.n245 B.n101 71.676
R1050 B.n249 B.n102 71.676
R1051 B.n253 B.n103 71.676
R1052 B.n257 B.n104 71.676
R1053 B.n261 B.n105 71.676
R1054 B.n265 B.n106 71.676
R1055 B.n269 B.n107 71.676
R1056 B.n273 B.n108 71.676
R1057 B.n277 B.n109 71.676
R1058 B.n281 B.n110 71.676
R1059 B.n285 B.n111 71.676
R1060 B.n289 B.n112 71.676
R1061 B.n293 B.n113 71.676
R1062 B.n297 B.n114 71.676
R1063 B.n301 B.n115 71.676
R1064 B.n305 B.n116 71.676
R1065 B.n309 B.n117 71.676
R1066 B.n313 B.n118 71.676
R1067 B.n317 B.n119 71.676
R1068 B.n321 B.n120 71.676
R1069 B.n325 B.n121 71.676
R1070 B.n329 B.n122 71.676
R1071 B.n333 B.n123 71.676
R1072 B.n337 B.n124 71.676
R1073 B.n341 B.n125 71.676
R1074 B.n345 B.n126 71.676
R1075 B.n349 B.n127 71.676
R1076 B.n353 B.n128 71.676
R1077 B.n357 B.n129 71.676
R1078 B.n361 B.n130 71.676
R1079 B.n365 B.n131 71.676
R1080 B.n369 B.n132 71.676
R1081 B.n373 B.n133 71.676
R1082 B.n377 B.n134 71.676
R1083 B.n381 B.n135 71.676
R1084 B.n385 B.n136 71.676
R1085 B.n389 B.n137 71.676
R1086 B.n393 B.n138 71.676
R1087 B.n397 B.n139 71.676
R1088 B.n986 B.n140 71.676
R1089 B.n986 B.n985 71.676
R1090 B.n399 B.n139 71.676
R1091 B.n396 B.n138 71.676
R1092 B.n392 B.n137 71.676
R1093 B.n388 B.n136 71.676
R1094 B.n384 B.n135 71.676
R1095 B.n380 B.n134 71.676
R1096 B.n376 B.n133 71.676
R1097 B.n372 B.n132 71.676
R1098 B.n368 B.n131 71.676
R1099 B.n364 B.n130 71.676
R1100 B.n360 B.n129 71.676
R1101 B.n356 B.n128 71.676
R1102 B.n352 B.n127 71.676
R1103 B.n348 B.n126 71.676
R1104 B.n344 B.n125 71.676
R1105 B.n340 B.n124 71.676
R1106 B.n336 B.n123 71.676
R1107 B.n332 B.n122 71.676
R1108 B.n328 B.n121 71.676
R1109 B.n324 B.n120 71.676
R1110 B.n320 B.n119 71.676
R1111 B.n316 B.n118 71.676
R1112 B.n312 B.n117 71.676
R1113 B.n308 B.n116 71.676
R1114 B.n304 B.n115 71.676
R1115 B.n300 B.n114 71.676
R1116 B.n296 B.n113 71.676
R1117 B.n292 B.n112 71.676
R1118 B.n288 B.n111 71.676
R1119 B.n284 B.n110 71.676
R1120 B.n280 B.n109 71.676
R1121 B.n276 B.n108 71.676
R1122 B.n272 B.n107 71.676
R1123 B.n268 B.n106 71.676
R1124 B.n264 B.n105 71.676
R1125 B.n260 B.n104 71.676
R1126 B.n256 B.n103 71.676
R1127 B.n252 B.n102 71.676
R1128 B.n248 B.n101 71.676
R1129 B.n244 B.n100 71.676
R1130 B.n240 B.n99 71.676
R1131 B.n236 B.n98 71.676
R1132 B.n232 B.n97 71.676
R1133 B.n228 B.n96 71.676
R1134 B.n224 B.n95 71.676
R1135 B.n220 B.n94 71.676
R1136 B.n216 B.n93 71.676
R1137 B.n212 B.n92 71.676
R1138 B.n208 B.n91 71.676
R1139 B.n204 B.n90 71.676
R1140 B.n200 B.n89 71.676
R1141 B.n196 B.n88 71.676
R1142 B.n192 B.n87 71.676
R1143 B.n188 B.n86 71.676
R1144 B.n184 B.n85 71.676
R1145 B.n180 B.n84 71.676
R1146 B.n176 B.n83 71.676
R1147 B.n172 B.n82 71.676
R1148 B.n168 B.n81 71.676
R1149 B.n164 B.n80 71.676
R1150 B.n160 B.n79 71.676
R1151 B.n156 B.n78 71.676
R1152 B.n152 B.n77 71.676
R1153 B.n148 B.n76 71.676
R1154 B.n547 B.n477 71.676
R1155 B.n551 B.n550 71.676
R1156 B.n556 B.n555 71.676
R1157 B.n559 B.n558 71.676
R1158 B.n564 B.n563 71.676
R1159 B.n567 B.n566 71.676
R1160 B.n572 B.n571 71.676
R1161 B.n575 B.n574 71.676
R1162 B.n580 B.n579 71.676
R1163 B.n583 B.n582 71.676
R1164 B.n588 B.n587 71.676
R1165 B.n591 B.n590 71.676
R1166 B.n596 B.n595 71.676
R1167 B.n599 B.n598 71.676
R1168 B.n604 B.n603 71.676
R1169 B.n607 B.n606 71.676
R1170 B.n612 B.n611 71.676
R1171 B.n615 B.n614 71.676
R1172 B.n620 B.n619 71.676
R1173 B.n623 B.n622 71.676
R1174 B.n628 B.n627 71.676
R1175 B.n631 B.n630 71.676
R1176 B.n636 B.n635 71.676
R1177 B.n639 B.n638 71.676
R1178 B.n644 B.n643 71.676
R1179 B.n647 B.n646 71.676
R1180 B.n652 B.n651 71.676
R1181 B.n655 B.n654 71.676
R1182 B.n660 B.n659 71.676
R1183 B.n663 B.n662 71.676
R1184 B.n669 B.n668 71.676
R1185 B.n672 B.n671 71.676
R1186 B.n677 B.n676 71.676
R1187 B.n680 B.n679 71.676
R1188 B.n688 B.n687 71.676
R1189 B.n691 B.n690 71.676
R1190 B.n696 B.n695 71.676
R1191 B.n699 B.n698 71.676
R1192 B.n704 B.n703 71.676
R1193 B.n707 B.n706 71.676
R1194 B.n712 B.n711 71.676
R1195 B.n715 B.n714 71.676
R1196 B.n720 B.n719 71.676
R1197 B.n723 B.n722 71.676
R1198 B.n728 B.n727 71.676
R1199 B.n731 B.n730 71.676
R1200 B.n736 B.n735 71.676
R1201 B.n739 B.n738 71.676
R1202 B.n744 B.n743 71.676
R1203 B.n747 B.n746 71.676
R1204 B.n752 B.n751 71.676
R1205 B.n755 B.n754 71.676
R1206 B.n760 B.n759 71.676
R1207 B.n763 B.n762 71.676
R1208 B.n768 B.n767 71.676
R1209 B.n771 B.n770 71.676
R1210 B.n776 B.n775 71.676
R1211 B.n779 B.n778 71.676
R1212 B.n784 B.n783 71.676
R1213 B.n787 B.n786 71.676
R1214 B.n792 B.n791 71.676
R1215 B.n795 B.n794 71.676
R1216 B.n800 B.n799 71.676
R1217 B.n803 B.n802 71.676
R1218 B.n548 B.n547 71.676
R1219 B.n550 B.n544 71.676
R1220 B.n557 B.n556 71.676
R1221 B.n558 B.n542 71.676
R1222 B.n565 B.n564 71.676
R1223 B.n566 B.n540 71.676
R1224 B.n573 B.n572 71.676
R1225 B.n574 B.n538 71.676
R1226 B.n581 B.n580 71.676
R1227 B.n582 B.n536 71.676
R1228 B.n589 B.n588 71.676
R1229 B.n590 B.n534 71.676
R1230 B.n597 B.n596 71.676
R1231 B.n598 B.n532 71.676
R1232 B.n605 B.n604 71.676
R1233 B.n606 B.n530 71.676
R1234 B.n613 B.n612 71.676
R1235 B.n614 B.n528 71.676
R1236 B.n621 B.n620 71.676
R1237 B.n622 B.n526 71.676
R1238 B.n629 B.n628 71.676
R1239 B.n630 B.n524 71.676
R1240 B.n637 B.n636 71.676
R1241 B.n638 B.n522 71.676
R1242 B.n645 B.n644 71.676
R1243 B.n646 B.n520 71.676
R1244 B.n653 B.n652 71.676
R1245 B.n654 B.n518 71.676
R1246 B.n661 B.n660 71.676
R1247 B.n662 B.n514 71.676
R1248 B.n670 B.n669 71.676
R1249 B.n671 B.n512 71.676
R1250 B.n678 B.n677 71.676
R1251 B.n679 B.n510 71.676
R1252 B.n689 B.n688 71.676
R1253 B.n690 B.n508 71.676
R1254 B.n697 B.n696 71.676
R1255 B.n698 B.n506 71.676
R1256 B.n705 B.n704 71.676
R1257 B.n706 B.n504 71.676
R1258 B.n713 B.n712 71.676
R1259 B.n714 B.n502 71.676
R1260 B.n721 B.n720 71.676
R1261 B.n722 B.n500 71.676
R1262 B.n729 B.n728 71.676
R1263 B.n730 B.n498 71.676
R1264 B.n737 B.n736 71.676
R1265 B.n738 B.n496 71.676
R1266 B.n745 B.n744 71.676
R1267 B.n746 B.n494 71.676
R1268 B.n753 B.n752 71.676
R1269 B.n754 B.n492 71.676
R1270 B.n761 B.n760 71.676
R1271 B.n762 B.n490 71.676
R1272 B.n769 B.n768 71.676
R1273 B.n770 B.n488 71.676
R1274 B.n777 B.n776 71.676
R1275 B.n778 B.n486 71.676
R1276 B.n785 B.n784 71.676
R1277 B.n786 B.n484 71.676
R1278 B.n793 B.n792 71.676
R1279 B.n794 B.n482 71.676
R1280 B.n801 B.n800 71.676
R1281 B.n804 B.n803 71.676
R1282 B.n1071 B.n1070 71.676
R1283 B.n1071 B.n2 71.676
R1284 B.n809 B.n478 60.064
R1285 B.n988 B.n987 60.064
R1286 B.n146 B.n145 59.5399
R1287 B.n143 B.n142 59.5399
R1288 B.n685 B.n684 59.5399
R1289 B.n665 B.n516 59.5399
R1290 B.n145 B.n144 35.6853
R1291 B.n142 B.n141 35.6853
R1292 B.n684 B.n683 35.6853
R1293 B.n516 B.n515 35.6853
R1294 B.n811 B.n476 34.1859
R1295 B.n807 B.n806 34.1859
R1296 B.n984 B.n983 34.1859
R1297 B.n990 B.n73 34.1859
R1298 B.n809 B.n474 31.6619
R1299 B.n815 B.n474 31.6619
R1300 B.n815 B.n470 31.6619
R1301 B.n822 B.n470 31.6619
R1302 B.n822 B.n821 31.6619
R1303 B.n828 B.n463 31.6619
R1304 B.n834 B.n463 31.6619
R1305 B.n834 B.n459 31.6619
R1306 B.n840 B.n459 31.6619
R1307 B.n840 B.n455 31.6619
R1308 B.n846 B.n455 31.6619
R1309 B.n846 B.n451 31.6619
R1310 B.n852 B.n451 31.6619
R1311 B.n858 B.n447 31.6619
R1312 B.n858 B.n442 31.6619
R1313 B.n864 B.n442 31.6619
R1314 B.n864 B.n443 31.6619
R1315 B.n870 B.n435 31.6619
R1316 B.n876 B.n435 31.6619
R1317 B.n876 B.n431 31.6619
R1318 B.n883 B.n431 31.6619
R1319 B.n883 B.n882 31.6619
R1320 B.n889 B.n424 31.6619
R1321 B.n895 B.n424 31.6619
R1322 B.n895 B.n420 31.6619
R1323 B.n901 B.n420 31.6619
R1324 B.n907 B.n416 31.6619
R1325 B.n907 B.n412 31.6619
R1326 B.n913 B.n412 31.6619
R1327 B.n913 B.n408 31.6619
R1328 B.n920 B.n408 31.6619
R1329 B.n926 B.n404 31.6619
R1330 B.n926 B.n4 31.6619
R1331 B.n1069 B.n4 31.6619
R1332 B.n1069 B.n1068 31.6619
R1333 B.n1068 B.n1067 31.6619
R1334 B.n1067 B.n8 31.6619
R1335 B.n935 B.n8 31.6619
R1336 B.n1060 B.n1059 31.6619
R1337 B.n1059 B.n1058 31.6619
R1338 B.n1058 B.n15 31.6619
R1339 B.n1052 B.n15 31.6619
R1340 B.n1052 B.n1051 31.6619
R1341 B.n1050 B.n22 31.6619
R1342 B.n1044 B.n22 31.6619
R1343 B.n1044 B.n1043 31.6619
R1344 B.n1043 B.n1042 31.6619
R1345 B.n1036 B.n32 31.6619
R1346 B.n1036 B.n1035 31.6619
R1347 B.n1035 B.n1034 31.6619
R1348 B.n1034 B.n36 31.6619
R1349 B.n1028 B.n36 31.6619
R1350 B.n1027 B.n1026 31.6619
R1351 B.n1026 B.n43 31.6619
R1352 B.n1020 B.n43 31.6619
R1353 B.n1020 B.n1019 31.6619
R1354 B.n1018 B.n50 31.6619
R1355 B.n1012 B.n50 31.6619
R1356 B.n1012 B.n1011 31.6619
R1357 B.n1011 B.n1010 31.6619
R1358 B.n1010 B.n57 31.6619
R1359 B.n1004 B.n57 31.6619
R1360 B.n1004 B.n1003 31.6619
R1361 B.n1003 B.n1002 31.6619
R1362 B.n996 B.n67 31.6619
R1363 B.n996 B.n995 31.6619
R1364 B.n995 B.n994 31.6619
R1365 B.n994 B.n71 31.6619
R1366 B.n988 B.n71 31.6619
R1367 B.n443 B.t5 30.2651
R1368 B.t4 B.n1027 30.2651
R1369 B.n821 B.t11 29.3338
R1370 B.n67 B.t15 29.3338
R1371 B.t6 B.n404 25.609
R1372 B.n935 B.t1 25.609
R1373 B.n901 B.t8 24.6777
R1374 B.t7 B.n1050 24.6777
R1375 B.n889 B.t3 20.0217
R1376 B.n1042 B.t9 20.0217
R1377 B B.n1072 18.0485
R1378 B.n852 B.t2 17.228
R1379 B.t0 B.n1018 17.228
R1380 B.t2 B.n447 14.4344
R1381 B.n1019 B.t0 14.4344
R1382 B.n882 B.t3 11.6407
R1383 B.n32 B.t9 11.6407
R1384 B.n812 B.n811 10.6151
R1385 B.n813 B.n812 10.6151
R1386 B.n813 B.n468 10.6151
R1387 B.n824 B.n468 10.6151
R1388 B.n825 B.n824 10.6151
R1389 B.n826 B.n825 10.6151
R1390 B.n826 B.n461 10.6151
R1391 B.n836 B.n461 10.6151
R1392 B.n837 B.n836 10.6151
R1393 B.n838 B.n837 10.6151
R1394 B.n838 B.n453 10.6151
R1395 B.n848 B.n453 10.6151
R1396 B.n849 B.n848 10.6151
R1397 B.n850 B.n849 10.6151
R1398 B.n850 B.n445 10.6151
R1399 B.n860 B.n445 10.6151
R1400 B.n861 B.n860 10.6151
R1401 B.n862 B.n861 10.6151
R1402 B.n862 B.n437 10.6151
R1403 B.n872 B.n437 10.6151
R1404 B.n873 B.n872 10.6151
R1405 B.n874 B.n873 10.6151
R1406 B.n874 B.n429 10.6151
R1407 B.n885 B.n429 10.6151
R1408 B.n886 B.n885 10.6151
R1409 B.n887 B.n886 10.6151
R1410 B.n887 B.n422 10.6151
R1411 B.n897 B.n422 10.6151
R1412 B.n898 B.n897 10.6151
R1413 B.n899 B.n898 10.6151
R1414 B.n899 B.n414 10.6151
R1415 B.n909 B.n414 10.6151
R1416 B.n910 B.n909 10.6151
R1417 B.n911 B.n910 10.6151
R1418 B.n911 B.n406 10.6151
R1419 B.n922 B.n406 10.6151
R1420 B.n923 B.n922 10.6151
R1421 B.n924 B.n923 10.6151
R1422 B.n924 B.n0 10.6151
R1423 B.n546 B.n476 10.6151
R1424 B.n546 B.n545 10.6151
R1425 B.n552 B.n545 10.6151
R1426 B.n553 B.n552 10.6151
R1427 B.n554 B.n553 10.6151
R1428 B.n554 B.n543 10.6151
R1429 B.n560 B.n543 10.6151
R1430 B.n561 B.n560 10.6151
R1431 B.n562 B.n561 10.6151
R1432 B.n562 B.n541 10.6151
R1433 B.n568 B.n541 10.6151
R1434 B.n569 B.n568 10.6151
R1435 B.n570 B.n569 10.6151
R1436 B.n570 B.n539 10.6151
R1437 B.n576 B.n539 10.6151
R1438 B.n577 B.n576 10.6151
R1439 B.n578 B.n577 10.6151
R1440 B.n578 B.n537 10.6151
R1441 B.n584 B.n537 10.6151
R1442 B.n585 B.n584 10.6151
R1443 B.n586 B.n585 10.6151
R1444 B.n586 B.n535 10.6151
R1445 B.n592 B.n535 10.6151
R1446 B.n593 B.n592 10.6151
R1447 B.n594 B.n593 10.6151
R1448 B.n594 B.n533 10.6151
R1449 B.n600 B.n533 10.6151
R1450 B.n601 B.n600 10.6151
R1451 B.n602 B.n601 10.6151
R1452 B.n602 B.n531 10.6151
R1453 B.n608 B.n531 10.6151
R1454 B.n609 B.n608 10.6151
R1455 B.n610 B.n609 10.6151
R1456 B.n610 B.n529 10.6151
R1457 B.n616 B.n529 10.6151
R1458 B.n617 B.n616 10.6151
R1459 B.n618 B.n617 10.6151
R1460 B.n618 B.n527 10.6151
R1461 B.n624 B.n527 10.6151
R1462 B.n625 B.n624 10.6151
R1463 B.n626 B.n625 10.6151
R1464 B.n626 B.n525 10.6151
R1465 B.n632 B.n525 10.6151
R1466 B.n633 B.n632 10.6151
R1467 B.n634 B.n633 10.6151
R1468 B.n634 B.n523 10.6151
R1469 B.n640 B.n523 10.6151
R1470 B.n641 B.n640 10.6151
R1471 B.n642 B.n641 10.6151
R1472 B.n642 B.n521 10.6151
R1473 B.n648 B.n521 10.6151
R1474 B.n649 B.n648 10.6151
R1475 B.n650 B.n649 10.6151
R1476 B.n650 B.n519 10.6151
R1477 B.n656 B.n519 10.6151
R1478 B.n657 B.n656 10.6151
R1479 B.n658 B.n657 10.6151
R1480 B.n658 B.n517 10.6151
R1481 B.n664 B.n517 10.6151
R1482 B.n667 B.n666 10.6151
R1483 B.n667 B.n513 10.6151
R1484 B.n673 B.n513 10.6151
R1485 B.n674 B.n673 10.6151
R1486 B.n675 B.n674 10.6151
R1487 B.n675 B.n511 10.6151
R1488 B.n681 B.n511 10.6151
R1489 B.n682 B.n681 10.6151
R1490 B.n686 B.n682 10.6151
R1491 B.n692 B.n509 10.6151
R1492 B.n693 B.n692 10.6151
R1493 B.n694 B.n693 10.6151
R1494 B.n694 B.n507 10.6151
R1495 B.n700 B.n507 10.6151
R1496 B.n701 B.n700 10.6151
R1497 B.n702 B.n701 10.6151
R1498 B.n702 B.n505 10.6151
R1499 B.n708 B.n505 10.6151
R1500 B.n709 B.n708 10.6151
R1501 B.n710 B.n709 10.6151
R1502 B.n710 B.n503 10.6151
R1503 B.n716 B.n503 10.6151
R1504 B.n717 B.n716 10.6151
R1505 B.n718 B.n717 10.6151
R1506 B.n718 B.n501 10.6151
R1507 B.n724 B.n501 10.6151
R1508 B.n725 B.n724 10.6151
R1509 B.n726 B.n725 10.6151
R1510 B.n726 B.n499 10.6151
R1511 B.n732 B.n499 10.6151
R1512 B.n733 B.n732 10.6151
R1513 B.n734 B.n733 10.6151
R1514 B.n734 B.n497 10.6151
R1515 B.n740 B.n497 10.6151
R1516 B.n741 B.n740 10.6151
R1517 B.n742 B.n741 10.6151
R1518 B.n742 B.n495 10.6151
R1519 B.n748 B.n495 10.6151
R1520 B.n749 B.n748 10.6151
R1521 B.n750 B.n749 10.6151
R1522 B.n750 B.n493 10.6151
R1523 B.n756 B.n493 10.6151
R1524 B.n757 B.n756 10.6151
R1525 B.n758 B.n757 10.6151
R1526 B.n758 B.n491 10.6151
R1527 B.n764 B.n491 10.6151
R1528 B.n765 B.n764 10.6151
R1529 B.n766 B.n765 10.6151
R1530 B.n766 B.n489 10.6151
R1531 B.n772 B.n489 10.6151
R1532 B.n773 B.n772 10.6151
R1533 B.n774 B.n773 10.6151
R1534 B.n774 B.n487 10.6151
R1535 B.n780 B.n487 10.6151
R1536 B.n781 B.n780 10.6151
R1537 B.n782 B.n781 10.6151
R1538 B.n782 B.n485 10.6151
R1539 B.n788 B.n485 10.6151
R1540 B.n789 B.n788 10.6151
R1541 B.n790 B.n789 10.6151
R1542 B.n790 B.n483 10.6151
R1543 B.n796 B.n483 10.6151
R1544 B.n797 B.n796 10.6151
R1545 B.n798 B.n797 10.6151
R1546 B.n798 B.n481 10.6151
R1547 B.n481 B.n480 10.6151
R1548 B.n805 B.n480 10.6151
R1549 B.n806 B.n805 10.6151
R1550 B.n807 B.n472 10.6151
R1551 B.n817 B.n472 10.6151
R1552 B.n818 B.n817 10.6151
R1553 B.n819 B.n818 10.6151
R1554 B.n819 B.n465 10.6151
R1555 B.n830 B.n465 10.6151
R1556 B.n831 B.n830 10.6151
R1557 B.n832 B.n831 10.6151
R1558 B.n832 B.n457 10.6151
R1559 B.n842 B.n457 10.6151
R1560 B.n843 B.n842 10.6151
R1561 B.n844 B.n843 10.6151
R1562 B.n844 B.n449 10.6151
R1563 B.n854 B.n449 10.6151
R1564 B.n855 B.n854 10.6151
R1565 B.n856 B.n855 10.6151
R1566 B.n856 B.n440 10.6151
R1567 B.n866 B.n440 10.6151
R1568 B.n867 B.n866 10.6151
R1569 B.n868 B.n867 10.6151
R1570 B.n868 B.n433 10.6151
R1571 B.n878 B.n433 10.6151
R1572 B.n879 B.n878 10.6151
R1573 B.n880 B.n879 10.6151
R1574 B.n880 B.n426 10.6151
R1575 B.n891 B.n426 10.6151
R1576 B.n892 B.n891 10.6151
R1577 B.n893 B.n892 10.6151
R1578 B.n893 B.n418 10.6151
R1579 B.n903 B.n418 10.6151
R1580 B.n904 B.n903 10.6151
R1581 B.n905 B.n904 10.6151
R1582 B.n905 B.n410 10.6151
R1583 B.n915 B.n410 10.6151
R1584 B.n916 B.n915 10.6151
R1585 B.n918 B.n916 10.6151
R1586 B.n918 B.n917 10.6151
R1587 B.n917 B.n402 10.6151
R1588 B.n929 B.n402 10.6151
R1589 B.n930 B.n929 10.6151
R1590 B.n931 B.n930 10.6151
R1591 B.n932 B.n931 10.6151
R1592 B.n933 B.n932 10.6151
R1593 B.n937 B.n933 10.6151
R1594 B.n938 B.n937 10.6151
R1595 B.n939 B.n938 10.6151
R1596 B.n940 B.n939 10.6151
R1597 B.n942 B.n940 10.6151
R1598 B.n943 B.n942 10.6151
R1599 B.n944 B.n943 10.6151
R1600 B.n945 B.n944 10.6151
R1601 B.n947 B.n945 10.6151
R1602 B.n948 B.n947 10.6151
R1603 B.n949 B.n948 10.6151
R1604 B.n950 B.n949 10.6151
R1605 B.n952 B.n950 10.6151
R1606 B.n953 B.n952 10.6151
R1607 B.n954 B.n953 10.6151
R1608 B.n955 B.n954 10.6151
R1609 B.n957 B.n955 10.6151
R1610 B.n958 B.n957 10.6151
R1611 B.n959 B.n958 10.6151
R1612 B.n960 B.n959 10.6151
R1613 B.n962 B.n960 10.6151
R1614 B.n963 B.n962 10.6151
R1615 B.n964 B.n963 10.6151
R1616 B.n965 B.n964 10.6151
R1617 B.n967 B.n965 10.6151
R1618 B.n968 B.n967 10.6151
R1619 B.n969 B.n968 10.6151
R1620 B.n970 B.n969 10.6151
R1621 B.n972 B.n970 10.6151
R1622 B.n973 B.n972 10.6151
R1623 B.n974 B.n973 10.6151
R1624 B.n975 B.n974 10.6151
R1625 B.n977 B.n975 10.6151
R1626 B.n978 B.n977 10.6151
R1627 B.n979 B.n978 10.6151
R1628 B.n980 B.n979 10.6151
R1629 B.n982 B.n980 10.6151
R1630 B.n983 B.n982 10.6151
R1631 B.n1064 B.n1 10.6151
R1632 B.n1064 B.n1063 10.6151
R1633 B.n1063 B.n1062 10.6151
R1634 B.n1062 B.n10 10.6151
R1635 B.n1056 B.n10 10.6151
R1636 B.n1056 B.n1055 10.6151
R1637 B.n1055 B.n1054 10.6151
R1638 B.n1054 B.n17 10.6151
R1639 B.n1048 B.n17 10.6151
R1640 B.n1048 B.n1047 10.6151
R1641 B.n1047 B.n1046 10.6151
R1642 B.n1046 B.n24 10.6151
R1643 B.n1040 B.n24 10.6151
R1644 B.n1040 B.n1039 10.6151
R1645 B.n1039 B.n1038 10.6151
R1646 B.n1038 B.n30 10.6151
R1647 B.n1032 B.n30 10.6151
R1648 B.n1032 B.n1031 10.6151
R1649 B.n1031 B.n1030 10.6151
R1650 B.n1030 B.n38 10.6151
R1651 B.n1024 B.n38 10.6151
R1652 B.n1024 B.n1023 10.6151
R1653 B.n1023 B.n1022 10.6151
R1654 B.n1022 B.n45 10.6151
R1655 B.n1016 B.n45 10.6151
R1656 B.n1016 B.n1015 10.6151
R1657 B.n1015 B.n1014 10.6151
R1658 B.n1014 B.n52 10.6151
R1659 B.n1008 B.n52 10.6151
R1660 B.n1008 B.n1007 10.6151
R1661 B.n1007 B.n1006 10.6151
R1662 B.n1006 B.n59 10.6151
R1663 B.n1000 B.n59 10.6151
R1664 B.n1000 B.n999 10.6151
R1665 B.n999 B.n998 10.6151
R1666 B.n998 B.n65 10.6151
R1667 B.n992 B.n65 10.6151
R1668 B.n992 B.n991 10.6151
R1669 B.n991 B.n990 10.6151
R1670 B.n147 B.n73 10.6151
R1671 B.n150 B.n147 10.6151
R1672 B.n151 B.n150 10.6151
R1673 B.n154 B.n151 10.6151
R1674 B.n155 B.n154 10.6151
R1675 B.n158 B.n155 10.6151
R1676 B.n159 B.n158 10.6151
R1677 B.n162 B.n159 10.6151
R1678 B.n163 B.n162 10.6151
R1679 B.n166 B.n163 10.6151
R1680 B.n167 B.n166 10.6151
R1681 B.n170 B.n167 10.6151
R1682 B.n171 B.n170 10.6151
R1683 B.n174 B.n171 10.6151
R1684 B.n175 B.n174 10.6151
R1685 B.n178 B.n175 10.6151
R1686 B.n179 B.n178 10.6151
R1687 B.n182 B.n179 10.6151
R1688 B.n183 B.n182 10.6151
R1689 B.n186 B.n183 10.6151
R1690 B.n187 B.n186 10.6151
R1691 B.n190 B.n187 10.6151
R1692 B.n191 B.n190 10.6151
R1693 B.n194 B.n191 10.6151
R1694 B.n195 B.n194 10.6151
R1695 B.n198 B.n195 10.6151
R1696 B.n199 B.n198 10.6151
R1697 B.n202 B.n199 10.6151
R1698 B.n203 B.n202 10.6151
R1699 B.n206 B.n203 10.6151
R1700 B.n207 B.n206 10.6151
R1701 B.n210 B.n207 10.6151
R1702 B.n211 B.n210 10.6151
R1703 B.n214 B.n211 10.6151
R1704 B.n215 B.n214 10.6151
R1705 B.n218 B.n215 10.6151
R1706 B.n219 B.n218 10.6151
R1707 B.n222 B.n219 10.6151
R1708 B.n223 B.n222 10.6151
R1709 B.n226 B.n223 10.6151
R1710 B.n227 B.n226 10.6151
R1711 B.n230 B.n227 10.6151
R1712 B.n231 B.n230 10.6151
R1713 B.n234 B.n231 10.6151
R1714 B.n235 B.n234 10.6151
R1715 B.n238 B.n235 10.6151
R1716 B.n239 B.n238 10.6151
R1717 B.n242 B.n239 10.6151
R1718 B.n243 B.n242 10.6151
R1719 B.n246 B.n243 10.6151
R1720 B.n247 B.n246 10.6151
R1721 B.n250 B.n247 10.6151
R1722 B.n251 B.n250 10.6151
R1723 B.n254 B.n251 10.6151
R1724 B.n255 B.n254 10.6151
R1725 B.n258 B.n255 10.6151
R1726 B.n259 B.n258 10.6151
R1727 B.n262 B.n259 10.6151
R1728 B.n263 B.n262 10.6151
R1729 B.n267 B.n266 10.6151
R1730 B.n270 B.n267 10.6151
R1731 B.n271 B.n270 10.6151
R1732 B.n274 B.n271 10.6151
R1733 B.n275 B.n274 10.6151
R1734 B.n278 B.n275 10.6151
R1735 B.n279 B.n278 10.6151
R1736 B.n282 B.n279 10.6151
R1737 B.n283 B.n282 10.6151
R1738 B.n287 B.n286 10.6151
R1739 B.n290 B.n287 10.6151
R1740 B.n291 B.n290 10.6151
R1741 B.n294 B.n291 10.6151
R1742 B.n295 B.n294 10.6151
R1743 B.n298 B.n295 10.6151
R1744 B.n299 B.n298 10.6151
R1745 B.n302 B.n299 10.6151
R1746 B.n303 B.n302 10.6151
R1747 B.n306 B.n303 10.6151
R1748 B.n307 B.n306 10.6151
R1749 B.n310 B.n307 10.6151
R1750 B.n311 B.n310 10.6151
R1751 B.n314 B.n311 10.6151
R1752 B.n315 B.n314 10.6151
R1753 B.n318 B.n315 10.6151
R1754 B.n319 B.n318 10.6151
R1755 B.n322 B.n319 10.6151
R1756 B.n323 B.n322 10.6151
R1757 B.n326 B.n323 10.6151
R1758 B.n327 B.n326 10.6151
R1759 B.n330 B.n327 10.6151
R1760 B.n331 B.n330 10.6151
R1761 B.n334 B.n331 10.6151
R1762 B.n335 B.n334 10.6151
R1763 B.n338 B.n335 10.6151
R1764 B.n339 B.n338 10.6151
R1765 B.n342 B.n339 10.6151
R1766 B.n343 B.n342 10.6151
R1767 B.n346 B.n343 10.6151
R1768 B.n347 B.n346 10.6151
R1769 B.n350 B.n347 10.6151
R1770 B.n351 B.n350 10.6151
R1771 B.n354 B.n351 10.6151
R1772 B.n355 B.n354 10.6151
R1773 B.n358 B.n355 10.6151
R1774 B.n359 B.n358 10.6151
R1775 B.n362 B.n359 10.6151
R1776 B.n363 B.n362 10.6151
R1777 B.n366 B.n363 10.6151
R1778 B.n367 B.n366 10.6151
R1779 B.n370 B.n367 10.6151
R1780 B.n371 B.n370 10.6151
R1781 B.n374 B.n371 10.6151
R1782 B.n375 B.n374 10.6151
R1783 B.n378 B.n375 10.6151
R1784 B.n379 B.n378 10.6151
R1785 B.n382 B.n379 10.6151
R1786 B.n383 B.n382 10.6151
R1787 B.n386 B.n383 10.6151
R1788 B.n387 B.n386 10.6151
R1789 B.n390 B.n387 10.6151
R1790 B.n391 B.n390 10.6151
R1791 B.n394 B.n391 10.6151
R1792 B.n395 B.n394 10.6151
R1793 B.n398 B.n395 10.6151
R1794 B.n400 B.n398 10.6151
R1795 B.n401 B.n400 10.6151
R1796 B.n984 B.n401 10.6151
R1797 B.n665 B.n664 9.36635
R1798 B.n685 B.n509 9.36635
R1799 B.n263 B.n146 9.36635
R1800 B.n286 B.n143 9.36635
R1801 B.n1072 B.n0 8.11757
R1802 B.n1072 B.n1 8.11757
R1803 B.t8 B.n416 6.98463
R1804 B.n1051 B.t7 6.98463
R1805 B.n920 B.t6 6.05341
R1806 B.n1060 B.t1 6.05341
R1807 B.n828 B.t11 2.32854
R1808 B.n1002 B.t15 2.32854
R1809 B.n870 B.t5 1.39733
R1810 B.n1028 B.t4 1.39733
R1811 B.n666 B.n665 1.24928
R1812 B.n686 B.n685 1.24928
R1813 B.n266 B.n146 1.24928
R1814 B.n283 B.n143 1.24928
R1815 VN.n7 VN.t5 325.976
R1816 VN.n34 VN.t7 325.976
R1817 VN.n12 VN.t2 292.872
R1818 VN.n6 VN.t4 292.872
R1819 VN.n18 VN.t1 292.872
R1820 VN.n25 VN.t0 292.872
R1821 VN.n39 VN.t8 292.872
R1822 VN.n33 VN.t9 292.872
R1823 VN.n45 VN.t3 292.872
R1824 VN.n52 VN.t6 292.872
R1825 VN.n26 VN.n25 176.959
R1826 VN.n53 VN.n52 176.959
R1827 VN.n51 VN.n27 161.3
R1828 VN.n50 VN.n49 161.3
R1829 VN.n48 VN.n28 161.3
R1830 VN.n47 VN.n46 161.3
R1831 VN.n44 VN.n29 161.3
R1832 VN.n43 VN.n42 161.3
R1833 VN.n41 VN.n30 161.3
R1834 VN.n40 VN.n39 161.3
R1835 VN.n38 VN.n31 161.3
R1836 VN.n37 VN.n36 161.3
R1837 VN.n35 VN.n32 161.3
R1838 VN.n24 VN.n0 161.3
R1839 VN.n23 VN.n22 161.3
R1840 VN.n21 VN.n1 161.3
R1841 VN.n20 VN.n19 161.3
R1842 VN.n17 VN.n2 161.3
R1843 VN.n16 VN.n15 161.3
R1844 VN.n14 VN.n3 161.3
R1845 VN.n13 VN.n12 161.3
R1846 VN.n11 VN.n4 161.3
R1847 VN.n10 VN.n9 161.3
R1848 VN.n8 VN.n5 161.3
R1849 VN.n23 VN.n1 56.5193
R1850 VN.n50 VN.n28 56.5193
R1851 VN VN.n53 52.2903
R1852 VN.n7 VN.n6 49.6167
R1853 VN.n34 VN.n33 49.6167
R1854 VN.n11 VN.n10 48.2635
R1855 VN.n16 VN.n3 48.2635
R1856 VN.n38 VN.n37 48.2635
R1857 VN.n43 VN.n30 48.2635
R1858 VN.n10 VN.n5 32.7233
R1859 VN.n17 VN.n16 32.7233
R1860 VN.n37 VN.n32 32.7233
R1861 VN.n44 VN.n43 32.7233
R1862 VN.n12 VN.n11 24.4675
R1863 VN.n12 VN.n3 24.4675
R1864 VN.n19 VN.n1 24.4675
R1865 VN.n24 VN.n23 24.4675
R1866 VN.n39 VN.n30 24.4675
R1867 VN.n39 VN.n38 24.4675
R1868 VN.n46 VN.n28 24.4675
R1869 VN.n51 VN.n50 24.4675
R1870 VN.n35 VN.n34 17.9026
R1871 VN.n8 VN.n7 17.9026
R1872 VN.n6 VN.n5 16.6381
R1873 VN.n18 VN.n17 16.6381
R1874 VN.n33 VN.n32 16.6381
R1875 VN.n45 VN.n44 16.6381
R1876 VN.n25 VN.n24 8.80862
R1877 VN.n52 VN.n51 8.80862
R1878 VN.n19 VN.n18 7.82994
R1879 VN.n46 VN.n45 7.82994
R1880 VN.n53 VN.n27 0.189894
R1881 VN.n49 VN.n27 0.189894
R1882 VN.n49 VN.n48 0.189894
R1883 VN.n48 VN.n47 0.189894
R1884 VN.n47 VN.n29 0.189894
R1885 VN.n42 VN.n29 0.189894
R1886 VN.n42 VN.n41 0.189894
R1887 VN.n41 VN.n40 0.189894
R1888 VN.n40 VN.n31 0.189894
R1889 VN.n36 VN.n31 0.189894
R1890 VN.n36 VN.n35 0.189894
R1891 VN.n9 VN.n8 0.189894
R1892 VN.n9 VN.n4 0.189894
R1893 VN.n13 VN.n4 0.189894
R1894 VN.n14 VN.n13 0.189894
R1895 VN.n15 VN.n14 0.189894
R1896 VN.n15 VN.n2 0.189894
R1897 VN.n20 VN.n2 0.189894
R1898 VN.n21 VN.n20 0.189894
R1899 VN.n22 VN.n21 0.189894
R1900 VN.n22 VN.n0 0.189894
R1901 VN.n26 VN.n0 0.189894
R1902 VN VN.n26 0.0516364
R1903 VTAIL.n416 VTAIL.n320 289.615
R1904 VTAIL.n98 VTAIL.n2 289.615
R1905 VTAIL.n314 VTAIL.n218 289.615
R1906 VTAIL.n208 VTAIL.n112 289.615
R1907 VTAIL.n352 VTAIL.n351 185
R1908 VTAIL.n357 VTAIL.n356 185
R1909 VTAIL.n359 VTAIL.n358 185
R1910 VTAIL.n348 VTAIL.n347 185
R1911 VTAIL.n365 VTAIL.n364 185
R1912 VTAIL.n367 VTAIL.n366 185
R1913 VTAIL.n344 VTAIL.n343 185
R1914 VTAIL.n373 VTAIL.n372 185
R1915 VTAIL.n375 VTAIL.n374 185
R1916 VTAIL.n340 VTAIL.n339 185
R1917 VTAIL.n381 VTAIL.n380 185
R1918 VTAIL.n383 VTAIL.n382 185
R1919 VTAIL.n336 VTAIL.n335 185
R1920 VTAIL.n389 VTAIL.n388 185
R1921 VTAIL.n391 VTAIL.n390 185
R1922 VTAIL.n332 VTAIL.n331 185
R1923 VTAIL.n398 VTAIL.n397 185
R1924 VTAIL.n399 VTAIL.n330 185
R1925 VTAIL.n401 VTAIL.n400 185
R1926 VTAIL.n328 VTAIL.n327 185
R1927 VTAIL.n407 VTAIL.n406 185
R1928 VTAIL.n409 VTAIL.n408 185
R1929 VTAIL.n324 VTAIL.n323 185
R1930 VTAIL.n415 VTAIL.n414 185
R1931 VTAIL.n417 VTAIL.n416 185
R1932 VTAIL.n34 VTAIL.n33 185
R1933 VTAIL.n39 VTAIL.n38 185
R1934 VTAIL.n41 VTAIL.n40 185
R1935 VTAIL.n30 VTAIL.n29 185
R1936 VTAIL.n47 VTAIL.n46 185
R1937 VTAIL.n49 VTAIL.n48 185
R1938 VTAIL.n26 VTAIL.n25 185
R1939 VTAIL.n55 VTAIL.n54 185
R1940 VTAIL.n57 VTAIL.n56 185
R1941 VTAIL.n22 VTAIL.n21 185
R1942 VTAIL.n63 VTAIL.n62 185
R1943 VTAIL.n65 VTAIL.n64 185
R1944 VTAIL.n18 VTAIL.n17 185
R1945 VTAIL.n71 VTAIL.n70 185
R1946 VTAIL.n73 VTAIL.n72 185
R1947 VTAIL.n14 VTAIL.n13 185
R1948 VTAIL.n80 VTAIL.n79 185
R1949 VTAIL.n81 VTAIL.n12 185
R1950 VTAIL.n83 VTAIL.n82 185
R1951 VTAIL.n10 VTAIL.n9 185
R1952 VTAIL.n89 VTAIL.n88 185
R1953 VTAIL.n91 VTAIL.n90 185
R1954 VTAIL.n6 VTAIL.n5 185
R1955 VTAIL.n97 VTAIL.n96 185
R1956 VTAIL.n99 VTAIL.n98 185
R1957 VTAIL.n315 VTAIL.n314 185
R1958 VTAIL.n313 VTAIL.n312 185
R1959 VTAIL.n222 VTAIL.n221 185
R1960 VTAIL.n307 VTAIL.n306 185
R1961 VTAIL.n305 VTAIL.n304 185
R1962 VTAIL.n226 VTAIL.n225 185
R1963 VTAIL.n299 VTAIL.n298 185
R1964 VTAIL.n297 VTAIL.n228 185
R1965 VTAIL.n296 VTAIL.n295 185
R1966 VTAIL.n231 VTAIL.n229 185
R1967 VTAIL.n290 VTAIL.n289 185
R1968 VTAIL.n288 VTAIL.n287 185
R1969 VTAIL.n235 VTAIL.n234 185
R1970 VTAIL.n282 VTAIL.n281 185
R1971 VTAIL.n280 VTAIL.n279 185
R1972 VTAIL.n239 VTAIL.n238 185
R1973 VTAIL.n274 VTAIL.n273 185
R1974 VTAIL.n272 VTAIL.n271 185
R1975 VTAIL.n243 VTAIL.n242 185
R1976 VTAIL.n266 VTAIL.n265 185
R1977 VTAIL.n264 VTAIL.n263 185
R1978 VTAIL.n247 VTAIL.n246 185
R1979 VTAIL.n258 VTAIL.n257 185
R1980 VTAIL.n256 VTAIL.n255 185
R1981 VTAIL.n251 VTAIL.n250 185
R1982 VTAIL.n209 VTAIL.n208 185
R1983 VTAIL.n207 VTAIL.n206 185
R1984 VTAIL.n116 VTAIL.n115 185
R1985 VTAIL.n201 VTAIL.n200 185
R1986 VTAIL.n199 VTAIL.n198 185
R1987 VTAIL.n120 VTAIL.n119 185
R1988 VTAIL.n193 VTAIL.n192 185
R1989 VTAIL.n191 VTAIL.n122 185
R1990 VTAIL.n190 VTAIL.n189 185
R1991 VTAIL.n125 VTAIL.n123 185
R1992 VTAIL.n184 VTAIL.n183 185
R1993 VTAIL.n182 VTAIL.n181 185
R1994 VTAIL.n129 VTAIL.n128 185
R1995 VTAIL.n176 VTAIL.n175 185
R1996 VTAIL.n174 VTAIL.n173 185
R1997 VTAIL.n133 VTAIL.n132 185
R1998 VTAIL.n168 VTAIL.n167 185
R1999 VTAIL.n166 VTAIL.n165 185
R2000 VTAIL.n137 VTAIL.n136 185
R2001 VTAIL.n160 VTAIL.n159 185
R2002 VTAIL.n158 VTAIL.n157 185
R2003 VTAIL.n141 VTAIL.n140 185
R2004 VTAIL.n152 VTAIL.n151 185
R2005 VTAIL.n150 VTAIL.n149 185
R2006 VTAIL.n145 VTAIL.n144 185
R2007 VTAIL.n353 VTAIL.t17 147.659
R2008 VTAIL.n35 VTAIL.t4 147.659
R2009 VTAIL.n252 VTAIL.t9 147.659
R2010 VTAIL.n146 VTAIL.t19 147.659
R2011 VTAIL.n357 VTAIL.n351 104.615
R2012 VTAIL.n358 VTAIL.n357 104.615
R2013 VTAIL.n358 VTAIL.n347 104.615
R2014 VTAIL.n365 VTAIL.n347 104.615
R2015 VTAIL.n366 VTAIL.n365 104.615
R2016 VTAIL.n366 VTAIL.n343 104.615
R2017 VTAIL.n373 VTAIL.n343 104.615
R2018 VTAIL.n374 VTAIL.n373 104.615
R2019 VTAIL.n374 VTAIL.n339 104.615
R2020 VTAIL.n381 VTAIL.n339 104.615
R2021 VTAIL.n382 VTAIL.n381 104.615
R2022 VTAIL.n382 VTAIL.n335 104.615
R2023 VTAIL.n389 VTAIL.n335 104.615
R2024 VTAIL.n390 VTAIL.n389 104.615
R2025 VTAIL.n390 VTAIL.n331 104.615
R2026 VTAIL.n398 VTAIL.n331 104.615
R2027 VTAIL.n399 VTAIL.n398 104.615
R2028 VTAIL.n400 VTAIL.n399 104.615
R2029 VTAIL.n400 VTAIL.n327 104.615
R2030 VTAIL.n407 VTAIL.n327 104.615
R2031 VTAIL.n408 VTAIL.n407 104.615
R2032 VTAIL.n408 VTAIL.n323 104.615
R2033 VTAIL.n415 VTAIL.n323 104.615
R2034 VTAIL.n416 VTAIL.n415 104.615
R2035 VTAIL.n39 VTAIL.n33 104.615
R2036 VTAIL.n40 VTAIL.n39 104.615
R2037 VTAIL.n40 VTAIL.n29 104.615
R2038 VTAIL.n47 VTAIL.n29 104.615
R2039 VTAIL.n48 VTAIL.n47 104.615
R2040 VTAIL.n48 VTAIL.n25 104.615
R2041 VTAIL.n55 VTAIL.n25 104.615
R2042 VTAIL.n56 VTAIL.n55 104.615
R2043 VTAIL.n56 VTAIL.n21 104.615
R2044 VTAIL.n63 VTAIL.n21 104.615
R2045 VTAIL.n64 VTAIL.n63 104.615
R2046 VTAIL.n64 VTAIL.n17 104.615
R2047 VTAIL.n71 VTAIL.n17 104.615
R2048 VTAIL.n72 VTAIL.n71 104.615
R2049 VTAIL.n72 VTAIL.n13 104.615
R2050 VTAIL.n80 VTAIL.n13 104.615
R2051 VTAIL.n81 VTAIL.n80 104.615
R2052 VTAIL.n82 VTAIL.n81 104.615
R2053 VTAIL.n82 VTAIL.n9 104.615
R2054 VTAIL.n89 VTAIL.n9 104.615
R2055 VTAIL.n90 VTAIL.n89 104.615
R2056 VTAIL.n90 VTAIL.n5 104.615
R2057 VTAIL.n97 VTAIL.n5 104.615
R2058 VTAIL.n98 VTAIL.n97 104.615
R2059 VTAIL.n314 VTAIL.n313 104.615
R2060 VTAIL.n313 VTAIL.n221 104.615
R2061 VTAIL.n306 VTAIL.n221 104.615
R2062 VTAIL.n306 VTAIL.n305 104.615
R2063 VTAIL.n305 VTAIL.n225 104.615
R2064 VTAIL.n298 VTAIL.n225 104.615
R2065 VTAIL.n298 VTAIL.n297 104.615
R2066 VTAIL.n297 VTAIL.n296 104.615
R2067 VTAIL.n296 VTAIL.n229 104.615
R2068 VTAIL.n289 VTAIL.n229 104.615
R2069 VTAIL.n289 VTAIL.n288 104.615
R2070 VTAIL.n288 VTAIL.n234 104.615
R2071 VTAIL.n281 VTAIL.n234 104.615
R2072 VTAIL.n281 VTAIL.n280 104.615
R2073 VTAIL.n280 VTAIL.n238 104.615
R2074 VTAIL.n273 VTAIL.n238 104.615
R2075 VTAIL.n273 VTAIL.n272 104.615
R2076 VTAIL.n272 VTAIL.n242 104.615
R2077 VTAIL.n265 VTAIL.n242 104.615
R2078 VTAIL.n265 VTAIL.n264 104.615
R2079 VTAIL.n264 VTAIL.n246 104.615
R2080 VTAIL.n257 VTAIL.n246 104.615
R2081 VTAIL.n257 VTAIL.n256 104.615
R2082 VTAIL.n256 VTAIL.n250 104.615
R2083 VTAIL.n208 VTAIL.n207 104.615
R2084 VTAIL.n207 VTAIL.n115 104.615
R2085 VTAIL.n200 VTAIL.n115 104.615
R2086 VTAIL.n200 VTAIL.n199 104.615
R2087 VTAIL.n199 VTAIL.n119 104.615
R2088 VTAIL.n192 VTAIL.n119 104.615
R2089 VTAIL.n192 VTAIL.n191 104.615
R2090 VTAIL.n191 VTAIL.n190 104.615
R2091 VTAIL.n190 VTAIL.n123 104.615
R2092 VTAIL.n183 VTAIL.n123 104.615
R2093 VTAIL.n183 VTAIL.n182 104.615
R2094 VTAIL.n182 VTAIL.n128 104.615
R2095 VTAIL.n175 VTAIL.n128 104.615
R2096 VTAIL.n175 VTAIL.n174 104.615
R2097 VTAIL.n174 VTAIL.n132 104.615
R2098 VTAIL.n167 VTAIL.n132 104.615
R2099 VTAIL.n167 VTAIL.n166 104.615
R2100 VTAIL.n166 VTAIL.n136 104.615
R2101 VTAIL.n159 VTAIL.n136 104.615
R2102 VTAIL.n159 VTAIL.n158 104.615
R2103 VTAIL.n158 VTAIL.n140 104.615
R2104 VTAIL.n151 VTAIL.n140 104.615
R2105 VTAIL.n151 VTAIL.n150 104.615
R2106 VTAIL.n150 VTAIL.n144 104.615
R2107 VTAIL.t17 VTAIL.n351 52.3082
R2108 VTAIL.t4 VTAIL.n33 52.3082
R2109 VTAIL.t9 VTAIL.n250 52.3082
R2110 VTAIL.t19 VTAIL.n144 52.3082
R2111 VTAIL.n217 VTAIL.n216 46.1028
R2112 VTAIL.n215 VTAIL.n214 46.1028
R2113 VTAIL.n111 VTAIL.n110 46.1028
R2114 VTAIL.n109 VTAIL.n108 46.1028
R2115 VTAIL.n423 VTAIL.n422 46.1027
R2116 VTAIL.n1 VTAIL.n0 46.1027
R2117 VTAIL.n105 VTAIL.n104 46.1027
R2118 VTAIL.n107 VTAIL.n106 46.1027
R2119 VTAIL.n421 VTAIL.n420 34.3187
R2120 VTAIL.n103 VTAIL.n102 34.3187
R2121 VTAIL.n319 VTAIL.n318 34.3187
R2122 VTAIL.n213 VTAIL.n212 34.3187
R2123 VTAIL.n109 VTAIL.n107 31.3583
R2124 VTAIL.n421 VTAIL.n319 29.7721
R2125 VTAIL.n353 VTAIL.n352 15.6677
R2126 VTAIL.n35 VTAIL.n34 15.6677
R2127 VTAIL.n252 VTAIL.n251 15.6677
R2128 VTAIL.n146 VTAIL.n145 15.6677
R2129 VTAIL.n401 VTAIL.n330 13.1884
R2130 VTAIL.n83 VTAIL.n12 13.1884
R2131 VTAIL.n299 VTAIL.n228 13.1884
R2132 VTAIL.n193 VTAIL.n122 13.1884
R2133 VTAIL.n356 VTAIL.n355 12.8005
R2134 VTAIL.n397 VTAIL.n396 12.8005
R2135 VTAIL.n402 VTAIL.n328 12.8005
R2136 VTAIL.n38 VTAIL.n37 12.8005
R2137 VTAIL.n79 VTAIL.n78 12.8005
R2138 VTAIL.n84 VTAIL.n10 12.8005
R2139 VTAIL.n300 VTAIL.n226 12.8005
R2140 VTAIL.n295 VTAIL.n230 12.8005
R2141 VTAIL.n255 VTAIL.n254 12.8005
R2142 VTAIL.n194 VTAIL.n120 12.8005
R2143 VTAIL.n189 VTAIL.n124 12.8005
R2144 VTAIL.n149 VTAIL.n148 12.8005
R2145 VTAIL.n359 VTAIL.n350 12.0247
R2146 VTAIL.n395 VTAIL.n332 12.0247
R2147 VTAIL.n406 VTAIL.n405 12.0247
R2148 VTAIL.n41 VTAIL.n32 12.0247
R2149 VTAIL.n77 VTAIL.n14 12.0247
R2150 VTAIL.n88 VTAIL.n87 12.0247
R2151 VTAIL.n304 VTAIL.n303 12.0247
R2152 VTAIL.n294 VTAIL.n231 12.0247
R2153 VTAIL.n258 VTAIL.n249 12.0247
R2154 VTAIL.n198 VTAIL.n197 12.0247
R2155 VTAIL.n188 VTAIL.n125 12.0247
R2156 VTAIL.n152 VTAIL.n143 12.0247
R2157 VTAIL.n360 VTAIL.n348 11.249
R2158 VTAIL.n392 VTAIL.n391 11.249
R2159 VTAIL.n409 VTAIL.n326 11.249
R2160 VTAIL.n42 VTAIL.n30 11.249
R2161 VTAIL.n74 VTAIL.n73 11.249
R2162 VTAIL.n91 VTAIL.n8 11.249
R2163 VTAIL.n307 VTAIL.n224 11.249
R2164 VTAIL.n291 VTAIL.n290 11.249
R2165 VTAIL.n259 VTAIL.n247 11.249
R2166 VTAIL.n201 VTAIL.n118 11.249
R2167 VTAIL.n185 VTAIL.n184 11.249
R2168 VTAIL.n153 VTAIL.n141 11.249
R2169 VTAIL.n364 VTAIL.n363 10.4732
R2170 VTAIL.n388 VTAIL.n334 10.4732
R2171 VTAIL.n410 VTAIL.n324 10.4732
R2172 VTAIL.n46 VTAIL.n45 10.4732
R2173 VTAIL.n70 VTAIL.n16 10.4732
R2174 VTAIL.n92 VTAIL.n6 10.4732
R2175 VTAIL.n308 VTAIL.n222 10.4732
R2176 VTAIL.n287 VTAIL.n233 10.4732
R2177 VTAIL.n263 VTAIL.n262 10.4732
R2178 VTAIL.n202 VTAIL.n116 10.4732
R2179 VTAIL.n181 VTAIL.n127 10.4732
R2180 VTAIL.n157 VTAIL.n156 10.4732
R2181 VTAIL.n367 VTAIL.n346 9.69747
R2182 VTAIL.n387 VTAIL.n336 9.69747
R2183 VTAIL.n414 VTAIL.n413 9.69747
R2184 VTAIL.n49 VTAIL.n28 9.69747
R2185 VTAIL.n69 VTAIL.n18 9.69747
R2186 VTAIL.n96 VTAIL.n95 9.69747
R2187 VTAIL.n312 VTAIL.n311 9.69747
R2188 VTAIL.n286 VTAIL.n235 9.69747
R2189 VTAIL.n266 VTAIL.n245 9.69747
R2190 VTAIL.n206 VTAIL.n205 9.69747
R2191 VTAIL.n180 VTAIL.n129 9.69747
R2192 VTAIL.n160 VTAIL.n139 9.69747
R2193 VTAIL.n420 VTAIL.n419 9.45567
R2194 VTAIL.n102 VTAIL.n101 9.45567
R2195 VTAIL.n318 VTAIL.n317 9.45567
R2196 VTAIL.n212 VTAIL.n211 9.45567
R2197 VTAIL.n419 VTAIL.n418 9.3005
R2198 VTAIL.n322 VTAIL.n321 9.3005
R2199 VTAIL.n413 VTAIL.n412 9.3005
R2200 VTAIL.n411 VTAIL.n410 9.3005
R2201 VTAIL.n326 VTAIL.n325 9.3005
R2202 VTAIL.n405 VTAIL.n404 9.3005
R2203 VTAIL.n403 VTAIL.n402 9.3005
R2204 VTAIL.n342 VTAIL.n341 9.3005
R2205 VTAIL.n371 VTAIL.n370 9.3005
R2206 VTAIL.n369 VTAIL.n368 9.3005
R2207 VTAIL.n346 VTAIL.n345 9.3005
R2208 VTAIL.n363 VTAIL.n362 9.3005
R2209 VTAIL.n361 VTAIL.n360 9.3005
R2210 VTAIL.n350 VTAIL.n349 9.3005
R2211 VTAIL.n355 VTAIL.n354 9.3005
R2212 VTAIL.n377 VTAIL.n376 9.3005
R2213 VTAIL.n379 VTAIL.n378 9.3005
R2214 VTAIL.n338 VTAIL.n337 9.3005
R2215 VTAIL.n385 VTAIL.n384 9.3005
R2216 VTAIL.n387 VTAIL.n386 9.3005
R2217 VTAIL.n334 VTAIL.n333 9.3005
R2218 VTAIL.n393 VTAIL.n392 9.3005
R2219 VTAIL.n395 VTAIL.n394 9.3005
R2220 VTAIL.n396 VTAIL.n329 9.3005
R2221 VTAIL.n101 VTAIL.n100 9.3005
R2222 VTAIL.n4 VTAIL.n3 9.3005
R2223 VTAIL.n95 VTAIL.n94 9.3005
R2224 VTAIL.n93 VTAIL.n92 9.3005
R2225 VTAIL.n8 VTAIL.n7 9.3005
R2226 VTAIL.n87 VTAIL.n86 9.3005
R2227 VTAIL.n85 VTAIL.n84 9.3005
R2228 VTAIL.n24 VTAIL.n23 9.3005
R2229 VTAIL.n53 VTAIL.n52 9.3005
R2230 VTAIL.n51 VTAIL.n50 9.3005
R2231 VTAIL.n28 VTAIL.n27 9.3005
R2232 VTAIL.n45 VTAIL.n44 9.3005
R2233 VTAIL.n43 VTAIL.n42 9.3005
R2234 VTAIL.n32 VTAIL.n31 9.3005
R2235 VTAIL.n37 VTAIL.n36 9.3005
R2236 VTAIL.n59 VTAIL.n58 9.3005
R2237 VTAIL.n61 VTAIL.n60 9.3005
R2238 VTAIL.n20 VTAIL.n19 9.3005
R2239 VTAIL.n67 VTAIL.n66 9.3005
R2240 VTAIL.n69 VTAIL.n68 9.3005
R2241 VTAIL.n16 VTAIL.n15 9.3005
R2242 VTAIL.n75 VTAIL.n74 9.3005
R2243 VTAIL.n77 VTAIL.n76 9.3005
R2244 VTAIL.n78 VTAIL.n11 9.3005
R2245 VTAIL.n278 VTAIL.n277 9.3005
R2246 VTAIL.n237 VTAIL.n236 9.3005
R2247 VTAIL.n284 VTAIL.n283 9.3005
R2248 VTAIL.n286 VTAIL.n285 9.3005
R2249 VTAIL.n233 VTAIL.n232 9.3005
R2250 VTAIL.n292 VTAIL.n291 9.3005
R2251 VTAIL.n294 VTAIL.n293 9.3005
R2252 VTAIL.n230 VTAIL.n227 9.3005
R2253 VTAIL.n317 VTAIL.n316 9.3005
R2254 VTAIL.n220 VTAIL.n219 9.3005
R2255 VTAIL.n311 VTAIL.n310 9.3005
R2256 VTAIL.n309 VTAIL.n308 9.3005
R2257 VTAIL.n224 VTAIL.n223 9.3005
R2258 VTAIL.n303 VTAIL.n302 9.3005
R2259 VTAIL.n301 VTAIL.n300 9.3005
R2260 VTAIL.n276 VTAIL.n275 9.3005
R2261 VTAIL.n241 VTAIL.n240 9.3005
R2262 VTAIL.n270 VTAIL.n269 9.3005
R2263 VTAIL.n268 VTAIL.n267 9.3005
R2264 VTAIL.n245 VTAIL.n244 9.3005
R2265 VTAIL.n262 VTAIL.n261 9.3005
R2266 VTAIL.n260 VTAIL.n259 9.3005
R2267 VTAIL.n249 VTAIL.n248 9.3005
R2268 VTAIL.n254 VTAIL.n253 9.3005
R2269 VTAIL.n172 VTAIL.n171 9.3005
R2270 VTAIL.n131 VTAIL.n130 9.3005
R2271 VTAIL.n178 VTAIL.n177 9.3005
R2272 VTAIL.n180 VTAIL.n179 9.3005
R2273 VTAIL.n127 VTAIL.n126 9.3005
R2274 VTAIL.n186 VTAIL.n185 9.3005
R2275 VTAIL.n188 VTAIL.n187 9.3005
R2276 VTAIL.n124 VTAIL.n121 9.3005
R2277 VTAIL.n211 VTAIL.n210 9.3005
R2278 VTAIL.n114 VTAIL.n113 9.3005
R2279 VTAIL.n205 VTAIL.n204 9.3005
R2280 VTAIL.n203 VTAIL.n202 9.3005
R2281 VTAIL.n118 VTAIL.n117 9.3005
R2282 VTAIL.n197 VTAIL.n196 9.3005
R2283 VTAIL.n195 VTAIL.n194 9.3005
R2284 VTAIL.n170 VTAIL.n169 9.3005
R2285 VTAIL.n135 VTAIL.n134 9.3005
R2286 VTAIL.n164 VTAIL.n163 9.3005
R2287 VTAIL.n162 VTAIL.n161 9.3005
R2288 VTAIL.n139 VTAIL.n138 9.3005
R2289 VTAIL.n156 VTAIL.n155 9.3005
R2290 VTAIL.n154 VTAIL.n153 9.3005
R2291 VTAIL.n143 VTAIL.n142 9.3005
R2292 VTAIL.n148 VTAIL.n147 9.3005
R2293 VTAIL.n368 VTAIL.n344 8.92171
R2294 VTAIL.n384 VTAIL.n383 8.92171
R2295 VTAIL.n417 VTAIL.n322 8.92171
R2296 VTAIL.n50 VTAIL.n26 8.92171
R2297 VTAIL.n66 VTAIL.n65 8.92171
R2298 VTAIL.n99 VTAIL.n4 8.92171
R2299 VTAIL.n315 VTAIL.n220 8.92171
R2300 VTAIL.n283 VTAIL.n282 8.92171
R2301 VTAIL.n267 VTAIL.n243 8.92171
R2302 VTAIL.n209 VTAIL.n114 8.92171
R2303 VTAIL.n177 VTAIL.n176 8.92171
R2304 VTAIL.n161 VTAIL.n137 8.92171
R2305 VTAIL.n372 VTAIL.n371 8.14595
R2306 VTAIL.n380 VTAIL.n338 8.14595
R2307 VTAIL.n418 VTAIL.n320 8.14595
R2308 VTAIL.n54 VTAIL.n53 8.14595
R2309 VTAIL.n62 VTAIL.n20 8.14595
R2310 VTAIL.n100 VTAIL.n2 8.14595
R2311 VTAIL.n316 VTAIL.n218 8.14595
R2312 VTAIL.n279 VTAIL.n237 8.14595
R2313 VTAIL.n271 VTAIL.n270 8.14595
R2314 VTAIL.n210 VTAIL.n112 8.14595
R2315 VTAIL.n173 VTAIL.n131 8.14595
R2316 VTAIL.n165 VTAIL.n164 8.14595
R2317 VTAIL.n375 VTAIL.n342 7.3702
R2318 VTAIL.n379 VTAIL.n340 7.3702
R2319 VTAIL.n57 VTAIL.n24 7.3702
R2320 VTAIL.n61 VTAIL.n22 7.3702
R2321 VTAIL.n278 VTAIL.n239 7.3702
R2322 VTAIL.n274 VTAIL.n241 7.3702
R2323 VTAIL.n172 VTAIL.n133 7.3702
R2324 VTAIL.n168 VTAIL.n135 7.3702
R2325 VTAIL.n376 VTAIL.n375 6.59444
R2326 VTAIL.n376 VTAIL.n340 6.59444
R2327 VTAIL.n58 VTAIL.n57 6.59444
R2328 VTAIL.n58 VTAIL.n22 6.59444
R2329 VTAIL.n275 VTAIL.n239 6.59444
R2330 VTAIL.n275 VTAIL.n274 6.59444
R2331 VTAIL.n169 VTAIL.n133 6.59444
R2332 VTAIL.n169 VTAIL.n168 6.59444
R2333 VTAIL.n372 VTAIL.n342 5.81868
R2334 VTAIL.n380 VTAIL.n379 5.81868
R2335 VTAIL.n420 VTAIL.n320 5.81868
R2336 VTAIL.n54 VTAIL.n24 5.81868
R2337 VTAIL.n62 VTAIL.n61 5.81868
R2338 VTAIL.n102 VTAIL.n2 5.81868
R2339 VTAIL.n318 VTAIL.n218 5.81868
R2340 VTAIL.n279 VTAIL.n278 5.81868
R2341 VTAIL.n271 VTAIL.n241 5.81868
R2342 VTAIL.n212 VTAIL.n112 5.81868
R2343 VTAIL.n173 VTAIL.n172 5.81868
R2344 VTAIL.n165 VTAIL.n135 5.81868
R2345 VTAIL.n371 VTAIL.n344 5.04292
R2346 VTAIL.n383 VTAIL.n338 5.04292
R2347 VTAIL.n418 VTAIL.n417 5.04292
R2348 VTAIL.n53 VTAIL.n26 5.04292
R2349 VTAIL.n65 VTAIL.n20 5.04292
R2350 VTAIL.n100 VTAIL.n99 5.04292
R2351 VTAIL.n316 VTAIL.n315 5.04292
R2352 VTAIL.n282 VTAIL.n237 5.04292
R2353 VTAIL.n270 VTAIL.n243 5.04292
R2354 VTAIL.n210 VTAIL.n209 5.04292
R2355 VTAIL.n176 VTAIL.n131 5.04292
R2356 VTAIL.n164 VTAIL.n137 5.04292
R2357 VTAIL.n354 VTAIL.n353 4.38563
R2358 VTAIL.n36 VTAIL.n35 4.38563
R2359 VTAIL.n253 VTAIL.n252 4.38563
R2360 VTAIL.n147 VTAIL.n146 4.38563
R2361 VTAIL.n368 VTAIL.n367 4.26717
R2362 VTAIL.n384 VTAIL.n336 4.26717
R2363 VTAIL.n414 VTAIL.n322 4.26717
R2364 VTAIL.n50 VTAIL.n49 4.26717
R2365 VTAIL.n66 VTAIL.n18 4.26717
R2366 VTAIL.n96 VTAIL.n4 4.26717
R2367 VTAIL.n312 VTAIL.n220 4.26717
R2368 VTAIL.n283 VTAIL.n235 4.26717
R2369 VTAIL.n267 VTAIL.n266 4.26717
R2370 VTAIL.n206 VTAIL.n114 4.26717
R2371 VTAIL.n177 VTAIL.n129 4.26717
R2372 VTAIL.n161 VTAIL.n160 4.26717
R2373 VTAIL.n364 VTAIL.n346 3.49141
R2374 VTAIL.n388 VTAIL.n387 3.49141
R2375 VTAIL.n413 VTAIL.n324 3.49141
R2376 VTAIL.n46 VTAIL.n28 3.49141
R2377 VTAIL.n70 VTAIL.n69 3.49141
R2378 VTAIL.n95 VTAIL.n6 3.49141
R2379 VTAIL.n311 VTAIL.n222 3.49141
R2380 VTAIL.n287 VTAIL.n286 3.49141
R2381 VTAIL.n263 VTAIL.n245 3.49141
R2382 VTAIL.n205 VTAIL.n116 3.49141
R2383 VTAIL.n181 VTAIL.n180 3.49141
R2384 VTAIL.n157 VTAIL.n139 3.49141
R2385 VTAIL.n363 VTAIL.n348 2.71565
R2386 VTAIL.n391 VTAIL.n334 2.71565
R2387 VTAIL.n410 VTAIL.n409 2.71565
R2388 VTAIL.n45 VTAIL.n30 2.71565
R2389 VTAIL.n73 VTAIL.n16 2.71565
R2390 VTAIL.n92 VTAIL.n91 2.71565
R2391 VTAIL.n308 VTAIL.n307 2.71565
R2392 VTAIL.n290 VTAIL.n233 2.71565
R2393 VTAIL.n262 VTAIL.n247 2.71565
R2394 VTAIL.n202 VTAIL.n201 2.71565
R2395 VTAIL.n184 VTAIL.n127 2.71565
R2396 VTAIL.n156 VTAIL.n141 2.71565
R2397 VTAIL.n360 VTAIL.n359 1.93989
R2398 VTAIL.n392 VTAIL.n332 1.93989
R2399 VTAIL.n406 VTAIL.n326 1.93989
R2400 VTAIL.n42 VTAIL.n41 1.93989
R2401 VTAIL.n74 VTAIL.n14 1.93989
R2402 VTAIL.n88 VTAIL.n8 1.93989
R2403 VTAIL.n304 VTAIL.n224 1.93989
R2404 VTAIL.n291 VTAIL.n231 1.93989
R2405 VTAIL.n259 VTAIL.n258 1.93989
R2406 VTAIL.n198 VTAIL.n118 1.93989
R2407 VTAIL.n185 VTAIL.n125 1.93989
R2408 VTAIL.n153 VTAIL.n152 1.93989
R2409 VTAIL.n111 VTAIL.n109 1.58671
R2410 VTAIL.n213 VTAIL.n111 1.58671
R2411 VTAIL.n217 VTAIL.n215 1.58671
R2412 VTAIL.n319 VTAIL.n217 1.58671
R2413 VTAIL.n107 VTAIL.n105 1.58671
R2414 VTAIL.n105 VTAIL.n103 1.58671
R2415 VTAIL.n423 VTAIL.n421 1.58671
R2416 VTAIL.n215 VTAIL.n213 1.26343
R2417 VTAIL.n103 VTAIL.n1 1.26343
R2418 VTAIL VTAIL.n1 1.24834
R2419 VTAIL.n356 VTAIL.n350 1.16414
R2420 VTAIL.n397 VTAIL.n395 1.16414
R2421 VTAIL.n405 VTAIL.n328 1.16414
R2422 VTAIL.n38 VTAIL.n32 1.16414
R2423 VTAIL.n79 VTAIL.n77 1.16414
R2424 VTAIL.n87 VTAIL.n10 1.16414
R2425 VTAIL.n303 VTAIL.n226 1.16414
R2426 VTAIL.n295 VTAIL.n294 1.16414
R2427 VTAIL.n255 VTAIL.n249 1.16414
R2428 VTAIL.n197 VTAIL.n120 1.16414
R2429 VTAIL.n189 VTAIL.n188 1.16414
R2430 VTAIL.n149 VTAIL.n143 1.16414
R2431 VTAIL.n422 VTAIL.t12 1.07952
R2432 VTAIL.n422 VTAIL.t11 1.07952
R2433 VTAIL.n0 VTAIL.t15 1.07952
R2434 VTAIL.n0 VTAIL.t18 1.07952
R2435 VTAIL.n104 VTAIL.t0 1.07952
R2436 VTAIL.n104 VTAIL.t6 1.07952
R2437 VTAIL.n106 VTAIL.t8 1.07952
R2438 VTAIL.n106 VTAIL.t3 1.07952
R2439 VTAIL.n216 VTAIL.t7 1.07952
R2440 VTAIL.n216 VTAIL.t1 1.07952
R2441 VTAIL.n214 VTAIL.t2 1.07952
R2442 VTAIL.n214 VTAIL.t5 1.07952
R2443 VTAIL.n110 VTAIL.t13 1.07952
R2444 VTAIL.n110 VTAIL.t16 1.07952
R2445 VTAIL.n108 VTAIL.t14 1.07952
R2446 VTAIL.n108 VTAIL.t10 1.07952
R2447 VTAIL.n355 VTAIL.n352 0.388379
R2448 VTAIL.n396 VTAIL.n330 0.388379
R2449 VTAIL.n402 VTAIL.n401 0.388379
R2450 VTAIL.n37 VTAIL.n34 0.388379
R2451 VTAIL.n78 VTAIL.n12 0.388379
R2452 VTAIL.n84 VTAIL.n83 0.388379
R2453 VTAIL.n300 VTAIL.n299 0.388379
R2454 VTAIL.n230 VTAIL.n228 0.388379
R2455 VTAIL.n254 VTAIL.n251 0.388379
R2456 VTAIL.n194 VTAIL.n193 0.388379
R2457 VTAIL.n124 VTAIL.n122 0.388379
R2458 VTAIL.n148 VTAIL.n145 0.388379
R2459 VTAIL VTAIL.n423 0.338862
R2460 VTAIL.n354 VTAIL.n349 0.155672
R2461 VTAIL.n361 VTAIL.n349 0.155672
R2462 VTAIL.n362 VTAIL.n361 0.155672
R2463 VTAIL.n362 VTAIL.n345 0.155672
R2464 VTAIL.n369 VTAIL.n345 0.155672
R2465 VTAIL.n370 VTAIL.n369 0.155672
R2466 VTAIL.n370 VTAIL.n341 0.155672
R2467 VTAIL.n377 VTAIL.n341 0.155672
R2468 VTAIL.n378 VTAIL.n377 0.155672
R2469 VTAIL.n378 VTAIL.n337 0.155672
R2470 VTAIL.n385 VTAIL.n337 0.155672
R2471 VTAIL.n386 VTAIL.n385 0.155672
R2472 VTAIL.n386 VTAIL.n333 0.155672
R2473 VTAIL.n393 VTAIL.n333 0.155672
R2474 VTAIL.n394 VTAIL.n393 0.155672
R2475 VTAIL.n394 VTAIL.n329 0.155672
R2476 VTAIL.n403 VTAIL.n329 0.155672
R2477 VTAIL.n404 VTAIL.n403 0.155672
R2478 VTAIL.n404 VTAIL.n325 0.155672
R2479 VTAIL.n411 VTAIL.n325 0.155672
R2480 VTAIL.n412 VTAIL.n411 0.155672
R2481 VTAIL.n412 VTAIL.n321 0.155672
R2482 VTAIL.n419 VTAIL.n321 0.155672
R2483 VTAIL.n36 VTAIL.n31 0.155672
R2484 VTAIL.n43 VTAIL.n31 0.155672
R2485 VTAIL.n44 VTAIL.n43 0.155672
R2486 VTAIL.n44 VTAIL.n27 0.155672
R2487 VTAIL.n51 VTAIL.n27 0.155672
R2488 VTAIL.n52 VTAIL.n51 0.155672
R2489 VTAIL.n52 VTAIL.n23 0.155672
R2490 VTAIL.n59 VTAIL.n23 0.155672
R2491 VTAIL.n60 VTAIL.n59 0.155672
R2492 VTAIL.n60 VTAIL.n19 0.155672
R2493 VTAIL.n67 VTAIL.n19 0.155672
R2494 VTAIL.n68 VTAIL.n67 0.155672
R2495 VTAIL.n68 VTAIL.n15 0.155672
R2496 VTAIL.n75 VTAIL.n15 0.155672
R2497 VTAIL.n76 VTAIL.n75 0.155672
R2498 VTAIL.n76 VTAIL.n11 0.155672
R2499 VTAIL.n85 VTAIL.n11 0.155672
R2500 VTAIL.n86 VTAIL.n85 0.155672
R2501 VTAIL.n86 VTAIL.n7 0.155672
R2502 VTAIL.n93 VTAIL.n7 0.155672
R2503 VTAIL.n94 VTAIL.n93 0.155672
R2504 VTAIL.n94 VTAIL.n3 0.155672
R2505 VTAIL.n101 VTAIL.n3 0.155672
R2506 VTAIL.n317 VTAIL.n219 0.155672
R2507 VTAIL.n310 VTAIL.n219 0.155672
R2508 VTAIL.n310 VTAIL.n309 0.155672
R2509 VTAIL.n309 VTAIL.n223 0.155672
R2510 VTAIL.n302 VTAIL.n223 0.155672
R2511 VTAIL.n302 VTAIL.n301 0.155672
R2512 VTAIL.n301 VTAIL.n227 0.155672
R2513 VTAIL.n293 VTAIL.n227 0.155672
R2514 VTAIL.n293 VTAIL.n292 0.155672
R2515 VTAIL.n292 VTAIL.n232 0.155672
R2516 VTAIL.n285 VTAIL.n232 0.155672
R2517 VTAIL.n285 VTAIL.n284 0.155672
R2518 VTAIL.n284 VTAIL.n236 0.155672
R2519 VTAIL.n277 VTAIL.n236 0.155672
R2520 VTAIL.n277 VTAIL.n276 0.155672
R2521 VTAIL.n276 VTAIL.n240 0.155672
R2522 VTAIL.n269 VTAIL.n240 0.155672
R2523 VTAIL.n269 VTAIL.n268 0.155672
R2524 VTAIL.n268 VTAIL.n244 0.155672
R2525 VTAIL.n261 VTAIL.n244 0.155672
R2526 VTAIL.n261 VTAIL.n260 0.155672
R2527 VTAIL.n260 VTAIL.n248 0.155672
R2528 VTAIL.n253 VTAIL.n248 0.155672
R2529 VTAIL.n211 VTAIL.n113 0.155672
R2530 VTAIL.n204 VTAIL.n113 0.155672
R2531 VTAIL.n204 VTAIL.n203 0.155672
R2532 VTAIL.n203 VTAIL.n117 0.155672
R2533 VTAIL.n196 VTAIL.n117 0.155672
R2534 VTAIL.n196 VTAIL.n195 0.155672
R2535 VTAIL.n195 VTAIL.n121 0.155672
R2536 VTAIL.n187 VTAIL.n121 0.155672
R2537 VTAIL.n187 VTAIL.n186 0.155672
R2538 VTAIL.n186 VTAIL.n126 0.155672
R2539 VTAIL.n179 VTAIL.n126 0.155672
R2540 VTAIL.n179 VTAIL.n178 0.155672
R2541 VTAIL.n178 VTAIL.n130 0.155672
R2542 VTAIL.n171 VTAIL.n130 0.155672
R2543 VTAIL.n171 VTAIL.n170 0.155672
R2544 VTAIL.n170 VTAIL.n134 0.155672
R2545 VTAIL.n163 VTAIL.n134 0.155672
R2546 VTAIL.n163 VTAIL.n162 0.155672
R2547 VTAIL.n162 VTAIL.n138 0.155672
R2548 VTAIL.n155 VTAIL.n138 0.155672
R2549 VTAIL.n155 VTAIL.n154 0.155672
R2550 VTAIL.n154 VTAIL.n142 0.155672
R2551 VTAIL.n147 VTAIL.n142 0.155672
R2552 VDD2.n201 VDD2.n105 289.615
R2553 VDD2.n96 VDD2.n0 289.615
R2554 VDD2.n202 VDD2.n201 185
R2555 VDD2.n200 VDD2.n199 185
R2556 VDD2.n109 VDD2.n108 185
R2557 VDD2.n194 VDD2.n193 185
R2558 VDD2.n192 VDD2.n191 185
R2559 VDD2.n113 VDD2.n112 185
R2560 VDD2.n186 VDD2.n185 185
R2561 VDD2.n184 VDD2.n115 185
R2562 VDD2.n183 VDD2.n182 185
R2563 VDD2.n118 VDD2.n116 185
R2564 VDD2.n177 VDD2.n176 185
R2565 VDD2.n175 VDD2.n174 185
R2566 VDD2.n122 VDD2.n121 185
R2567 VDD2.n169 VDD2.n168 185
R2568 VDD2.n167 VDD2.n166 185
R2569 VDD2.n126 VDD2.n125 185
R2570 VDD2.n161 VDD2.n160 185
R2571 VDD2.n159 VDD2.n158 185
R2572 VDD2.n130 VDD2.n129 185
R2573 VDD2.n153 VDD2.n152 185
R2574 VDD2.n151 VDD2.n150 185
R2575 VDD2.n134 VDD2.n133 185
R2576 VDD2.n145 VDD2.n144 185
R2577 VDD2.n143 VDD2.n142 185
R2578 VDD2.n138 VDD2.n137 185
R2579 VDD2.n32 VDD2.n31 185
R2580 VDD2.n37 VDD2.n36 185
R2581 VDD2.n39 VDD2.n38 185
R2582 VDD2.n28 VDD2.n27 185
R2583 VDD2.n45 VDD2.n44 185
R2584 VDD2.n47 VDD2.n46 185
R2585 VDD2.n24 VDD2.n23 185
R2586 VDD2.n53 VDD2.n52 185
R2587 VDD2.n55 VDD2.n54 185
R2588 VDD2.n20 VDD2.n19 185
R2589 VDD2.n61 VDD2.n60 185
R2590 VDD2.n63 VDD2.n62 185
R2591 VDD2.n16 VDD2.n15 185
R2592 VDD2.n69 VDD2.n68 185
R2593 VDD2.n71 VDD2.n70 185
R2594 VDD2.n12 VDD2.n11 185
R2595 VDD2.n78 VDD2.n77 185
R2596 VDD2.n79 VDD2.n10 185
R2597 VDD2.n81 VDD2.n80 185
R2598 VDD2.n8 VDD2.n7 185
R2599 VDD2.n87 VDD2.n86 185
R2600 VDD2.n89 VDD2.n88 185
R2601 VDD2.n4 VDD2.n3 185
R2602 VDD2.n95 VDD2.n94 185
R2603 VDD2.n97 VDD2.n96 185
R2604 VDD2.n139 VDD2.t3 147.659
R2605 VDD2.n33 VDD2.t4 147.659
R2606 VDD2.n201 VDD2.n200 104.615
R2607 VDD2.n200 VDD2.n108 104.615
R2608 VDD2.n193 VDD2.n108 104.615
R2609 VDD2.n193 VDD2.n192 104.615
R2610 VDD2.n192 VDD2.n112 104.615
R2611 VDD2.n185 VDD2.n112 104.615
R2612 VDD2.n185 VDD2.n184 104.615
R2613 VDD2.n184 VDD2.n183 104.615
R2614 VDD2.n183 VDD2.n116 104.615
R2615 VDD2.n176 VDD2.n116 104.615
R2616 VDD2.n176 VDD2.n175 104.615
R2617 VDD2.n175 VDD2.n121 104.615
R2618 VDD2.n168 VDD2.n121 104.615
R2619 VDD2.n168 VDD2.n167 104.615
R2620 VDD2.n167 VDD2.n125 104.615
R2621 VDD2.n160 VDD2.n125 104.615
R2622 VDD2.n160 VDD2.n159 104.615
R2623 VDD2.n159 VDD2.n129 104.615
R2624 VDD2.n152 VDD2.n129 104.615
R2625 VDD2.n152 VDD2.n151 104.615
R2626 VDD2.n151 VDD2.n133 104.615
R2627 VDD2.n144 VDD2.n133 104.615
R2628 VDD2.n144 VDD2.n143 104.615
R2629 VDD2.n143 VDD2.n137 104.615
R2630 VDD2.n37 VDD2.n31 104.615
R2631 VDD2.n38 VDD2.n37 104.615
R2632 VDD2.n38 VDD2.n27 104.615
R2633 VDD2.n45 VDD2.n27 104.615
R2634 VDD2.n46 VDD2.n45 104.615
R2635 VDD2.n46 VDD2.n23 104.615
R2636 VDD2.n53 VDD2.n23 104.615
R2637 VDD2.n54 VDD2.n53 104.615
R2638 VDD2.n54 VDD2.n19 104.615
R2639 VDD2.n61 VDD2.n19 104.615
R2640 VDD2.n62 VDD2.n61 104.615
R2641 VDD2.n62 VDD2.n15 104.615
R2642 VDD2.n69 VDD2.n15 104.615
R2643 VDD2.n70 VDD2.n69 104.615
R2644 VDD2.n70 VDD2.n11 104.615
R2645 VDD2.n78 VDD2.n11 104.615
R2646 VDD2.n79 VDD2.n78 104.615
R2647 VDD2.n80 VDD2.n79 104.615
R2648 VDD2.n80 VDD2.n7 104.615
R2649 VDD2.n87 VDD2.n7 104.615
R2650 VDD2.n88 VDD2.n87 104.615
R2651 VDD2.n88 VDD2.n3 104.615
R2652 VDD2.n95 VDD2.n3 104.615
R2653 VDD2.n96 VDD2.n95 104.615
R2654 VDD2.n104 VDD2.n103 63.9158
R2655 VDD2 VDD2.n209 63.9129
R2656 VDD2.n208 VDD2.n207 62.7816
R2657 VDD2.n102 VDD2.n101 62.7814
R2658 VDD2.n102 VDD2.n100 52.5837
R2659 VDD2.t3 VDD2.n137 52.3082
R2660 VDD2.t4 VDD2.n31 52.3082
R2661 VDD2.n206 VDD2.n205 50.9975
R2662 VDD2.n206 VDD2.n104 47.0687
R2663 VDD2.n139 VDD2.n138 15.6677
R2664 VDD2.n33 VDD2.n32 15.6677
R2665 VDD2.n186 VDD2.n115 13.1884
R2666 VDD2.n81 VDD2.n10 13.1884
R2667 VDD2.n187 VDD2.n113 12.8005
R2668 VDD2.n182 VDD2.n117 12.8005
R2669 VDD2.n142 VDD2.n141 12.8005
R2670 VDD2.n36 VDD2.n35 12.8005
R2671 VDD2.n77 VDD2.n76 12.8005
R2672 VDD2.n82 VDD2.n8 12.8005
R2673 VDD2.n191 VDD2.n190 12.0247
R2674 VDD2.n181 VDD2.n118 12.0247
R2675 VDD2.n145 VDD2.n136 12.0247
R2676 VDD2.n39 VDD2.n30 12.0247
R2677 VDD2.n75 VDD2.n12 12.0247
R2678 VDD2.n86 VDD2.n85 12.0247
R2679 VDD2.n194 VDD2.n111 11.249
R2680 VDD2.n178 VDD2.n177 11.249
R2681 VDD2.n146 VDD2.n134 11.249
R2682 VDD2.n40 VDD2.n28 11.249
R2683 VDD2.n72 VDD2.n71 11.249
R2684 VDD2.n89 VDD2.n6 11.249
R2685 VDD2.n195 VDD2.n109 10.4732
R2686 VDD2.n174 VDD2.n120 10.4732
R2687 VDD2.n150 VDD2.n149 10.4732
R2688 VDD2.n44 VDD2.n43 10.4732
R2689 VDD2.n68 VDD2.n14 10.4732
R2690 VDD2.n90 VDD2.n4 10.4732
R2691 VDD2.n199 VDD2.n198 9.69747
R2692 VDD2.n173 VDD2.n122 9.69747
R2693 VDD2.n153 VDD2.n132 9.69747
R2694 VDD2.n47 VDD2.n26 9.69747
R2695 VDD2.n67 VDD2.n16 9.69747
R2696 VDD2.n94 VDD2.n93 9.69747
R2697 VDD2.n205 VDD2.n204 9.45567
R2698 VDD2.n100 VDD2.n99 9.45567
R2699 VDD2.n165 VDD2.n164 9.3005
R2700 VDD2.n124 VDD2.n123 9.3005
R2701 VDD2.n171 VDD2.n170 9.3005
R2702 VDD2.n173 VDD2.n172 9.3005
R2703 VDD2.n120 VDD2.n119 9.3005
R2704 VDD2.n179 VDD2.n178 9.3005
R2705 VDD2.n181 VDD2.n180 9.3005
R2706 VDD2.n117 VDD2.n114 9.3005
R2707 VDD2.n204 VDD2.n203 9.3005
R2708 VDD2.n107 VDD2.n106 9.3005
R2709 VDD2.n198 VDD2.n197 9.3005
R2710 VDD2.n196 VDD2.n195 9.3005
R2711 VDD2.n111 VDD2.n110 9.3005
R2712 VDD2.n190 VDD2.n189 9.3005
R2713 VDD2.n188 VDD2.n187 9.3005
R2714 VDD2.n163 VDD2.n162 9.3005
R2715 VDD2.n128 VDD2.n127 9.3005
R2716 VDD2.n157 VDD2.n156 9.3005
R2717 VDD2.n155 VDD2.n154 9.3005
R2718 VDD2.n132 VDD2.n131 9.3005
R2719 VDD2.n149 VDD2.n148 9.3005
R2720 VDD2.n147 VDD2.n146 9.3005
R2721 VDD2.n136 VDD2.n135 9.3005
R2722 VDD2.n141 VDD2.n140 9.3005
R2723 VDD2.n99 VDD2.n98 9.3005
R2724 VDD2.n2 VDD2.n1 9.3005
R2725 VDD2.n93 VDD2.n92 9.3005
R2726 VDD2.n91 VDD2.n90 9.3005
R2727 VDD2.n6 VDD2.n5 9.3005
R2728 VDD2.n85 VDD2.n84 9.3005
R2729 VDD2.n83 VDD2.n82 9.3005
R2730 VDD2.n22 VDD2.n21 9.3005
R2731 VDD2.n51 VDD2.n50 9.3005
R2732 VDD2.n49 VDD2.n48 9.3005
R2733 VDD2.n26 VDD2.n25 9.3005
R2734 VDD2.n43 VDD2.n42 9.3005
R2735 VDD2.n41 VDD2.n40 9.3005
R2736 VDD2.n30 VDD2.n29 9.3005
R2737 VDD2.n35 VDD2.n34 9.3005
R2738 VDD2.n57 VDD2.n56 9.3005
R2739 VDD2.n59 VDD2.n58 9.3005
R2740 VDD2.n18 VDD2.n17 9.3005
R2741 VDD2.n65 VDD2.n64 9.3005
R2742 VDD2.n67 VDD2.n66 9.3005
R2743 VDD2.n14 VDD2.n13 9.3005
R2744 VDD2.n73 VDD2.n72 9.3005
R2745 VDD2.n75 VDD2.n74 9.3005
R2746 VDD2.n76 VDD2.n9 9.3005
R2747 VDD2.n202 VDD2.n107 8.92171
R2748 VDD2.n170 VDD2.n169 8.92171
R2749 VDD2.n154 VDD2.n130 8.92171
R2750 VDD2.n48 VDD2.n24 8.92171
R2751 VDD2.n64 VDD2.n63 8.92171
R2752 VDD2.n97 VDD2.n2 8.92171
R2753 VDD2.n203 VDD2.n105 8.14595
R2754 VDD2.n166 VDD2.n124 8.14595
R2755 VDD2.n158 VDD2.n157 8.14595
R2756 VDD2.n52 VDD2.n51 8.14595
R2757 VDD2.n60 VDD2.n18 8.14595
R2758 VDD2.n98 VDD2.n0 8.14595
R2759 VDD2.n165 VDD2.n126 7.3702
R2760 VDD2.n161 VDD2.n128 7.3702
R2761 VDD2.n55 VDD2.n22 7.3702
R2762 VDD2.n59 VDD2.n20 7.3702
R2763 VDD2.n162 VDD2.n126 6.59444
R2764 VDD2.n162 VDD2.n161 6.59444
R2765 VDD2.n56 VDD2.n55 6.59444
R2766 VDD2.n56 VDD2.n20 6.59444
R2767 VDD2.n205 VDD2.n105 5.81868
R2768 VDD2.n166 VDD2.n165 5.81868
R2769 VDD2.n158 VDD2.n128 5.81868
R2770 VDD2.n52 VDD2.n22 5.81868
R2771 VDD2.n60 VDD2.n59 5.81868
R2772 VDD2.n100 VDD2.n0 5.81868
R2773 VDD2.n203 VDD2.n202 5.04292
R2774 VDD2.n169 VDD2.n124 5.04292
R2775 VDD2.n157 VDD2.n130 5.04292
R2776 VDD2.n51 VDD2.n24 5.04292
R2777 VDD2.n63 VDD2.n18 5.04292
R2778 VDD2.n98 VDD2.n97 5.04292
R2779 VDD2.n140 VDD2.n139 4.38563
R2780 VDD2.n34 VDD2.n33 4.38563
R2781 VDD2.n199 VDD2.n107 4.26717
R2782 VDD2.n170 VDD2.n122 4.26717
R2783 VDD2.n154 VDD2.n153 4.26717
R2784 VDD2.n48 VDD2.n47 4.26717
R2785 VDD2.n64 VDD2.n16 4.26717
R2786 VDD2.n94 VDD2.n2 4.26717
R2787 VDD2.n198 VDD2.n109 3.49141
R2788 VDD2.n174 VDD2.n173 3.49141
R2789 VDD2.n150 VDD2.n132 3.49141
R2790 VDD2.n44 VDD2.n26 3.49141
R2791 VDD2.n68 VDD2.n67 3.49141
R2792 VDD2.n93 VDD2.n4 3.49141
R2793 VDD2.n195 VDD2.n194 2.71565
R2794 VDD2.n177 VDD2.n120 2.71565
R2795 VDD2.n149 VDD2.n134 2.71565
R2796 VDD2.n43 VDD2.n28 2.71565
R2797 VDD2.n71 VDD2.n14 2.71565
R2798 VDD2.n90 VDD2.n89 2.71565
R2799 VDD2.n191 VDD2.n111 1.93989
R2800 VDD2.n178 VDD2.n118 1.93989
R2801 VDD2.n146 VDD2.n145 1.93989
R2802 VDD2.n40 VDD2.n39 1.93989
R2803 VDD2.n72 VDD2.n12 1.93989
R2804 VDD2.n86 VDD2.n6 1.93989
R2805 VDD2.n208 VDD2.n206 1.58671
R2806 VDD2.n190 VDD2.n113 1.16414
R2807 VDD2.n182 VDD2.n181 1.16414
R2808 VDD2.n142 VDD2.n136 1.16414
R2809 VDD2.n36 VDD2.n30 1.16414
R2810 VDD2.n77 VDD2.n75 1.16414
R2811 VDD2.n85 VDD2.n8 1.16414
R2812 VDD2.n209 VDD2.t0 1.07952
R2813 VDD2.n209 VDD2.t2 1.07952
R2814 VDD2.n207 VDD2.t6 1.07952
R2815 VDD2.n207 VDD2.t1 1.07952
R2816 VDD2.n103 VDD2.t8 1.07952
R2817 VDD2.n103 VDD2.t9 1.07952
R2818 VDD2.n101 VDD2.t5 1.07952
R2819 VDD2.n101 VDD2.t7 1.07952
R2820 VDD2 VDD2.n208 0.455241
R2821 VDD2.n187 VDD2.n186 0.388379
R2822 VDD2.n117 VDD2.n115 0.388379
R2823 VDD2.n141 VDD2.n138 0.388379
R2824 VDD2.n35 VDD2.n32 0.388379
R2825 VDD2.n76 VDD2.n10 0.388379
R2826 VDD2.n82 VDD2.n81 0.388379
R2827 VDD2.n104 VDD2.n102 0.341706
R2828 VDD2.n204 VDD2.n106 0.155672
R2829 VDD2.n197 VDD2.n106 0.155672
R2830 VDD2.n197 VDD2.n196 0.155672
R2831 VDD2.n196 VDD2.n110 0.155672
R2832 VDD2.n189 VDD2.n110 0.155672
R2833 VDD2.n189 VDD2.n188 0.155672
R2834 VDD2.n188 VDD2.n114 0.155672
R2835 VDD2.n180 VDD2.n114 0.155672
R2836 VDD2.n180 VDD2.n179 0.155672
R2837 VDD2.n179 VDD2.n119 0.155672
R2838 VDD2.n172 VDD2.n119 0.155672
R2839 VDD2.n172 VDD2.n171 0.155672
R2840 VDD2.n171 VDD2.n123 0.155672
R2841 VDD2.n164 VDD2.n123 0.155672
R2842 VDD2.n164 VDD2.n163 0.155672
R2843 VDD2.n163 VDD2.n127 0.155672
R2844 VDD2.n156 VDD2.n127 0.155672
R2845 VDD2.n156 VDD2.n155 0.155672
R2846 VDD2.n155 VDD2.n131 0.155672
R2847 VDD2.n148 VDD2.n131 0.155672
R2848 VDD2.n148 VDD2.n147 0.155672
R2849 VDD2.n147 VDD2.n135 0.155672
R2850 VDD2.n140 VDD2.n135 0.155672
R2851 VDD2.n34 VDD2.n29 0.155672
R2852 VDD2.n41 VDD2.n29 0.155672
R2853 VDD2.n42 VDD2.n41 0.155672
R2854 VDD2.n42 VDD2.n25 0.155672
R2855 VDD2.n49 VDD2.n25 0.155672
R2856 VDD2.n50 VDD2.n49 0.155672
R2857 VDD2.n50 VDD2.n21 0.155672
R2858 VDD2.n57 VDD2.n21 0.155672
R2859 VDD2.n58 VDD2.n57 0.155672
R2860 VDD2.n58 VDD2.n17 0.155672
R2861 VDD2.n65 VDD2.n17 0.155672
R2862 VDD2.n66 VDD2.n65 0.155672
R2863 VDD2.n66 VDD2.n13 0.155672
R2864 VDD2.n73 VDD2.n13 0.155672
R2865 VDD2.n74 VDD2.n73 0.155672
R2866 VDD2.n74 VDD2.n9 0.155672
R2867 VDD2.n83 VDD2.n9 0.155672
R2868 VDD2.n84 VDD2.n83 0.155672
R2869 VDD2.n84 VDD2.n5 0.155672
R2870 VDD2.n91 VDD2.n5 0.155672
R2871 VDD2.n92 VDD2.n91 0.155672
R2872 VDD2.n92 VDD2.n1 0.155672
R2873 VDD2.n99 VDD2.n1 0.155672
R2874 VP.n15 VP.t9 325.976
R2875 VP.n48 VP.t6 292.872
R2876 VP.n35 VP.t3 292.872
R2877 VP.n41 VP.t4 292.872
R2878 VP.n54 VP.t7 292.872
R2879 VP.n61 VP.t8 292.872
R2880 VP.n20 VP.t0 292.872
R2881 VP.n33 VP.t5 292.872
R2882 VP.n26 VP.t2 292.872
R2883 VP.n14 VP.t1 292.872
R2884 VP.n36 VP.n35 176.959
R2885 VP.n62 VP.n61 176.959
R2886 VP.n34 VP.n33 176.959
R2887 VP.n16 VP.n13 161.3
R2888 VP.n18 VP.n17 161.3
R2889 VP.n19 VP.n12 161.3
R2890 VP.n21 VP.n20 161.3
R2891 VP.n22 VP.n11 161.3
R2892 VP.n24 VP.n23 161.3
R2893 VP.n25 VP.n10 161.3
R2894 VP.n28 VP.n27 161.3
R2895 VP.n29 VP.n9 161.3
R2896 VP.n31 VP.n30 161.3
R2897 VP.n32 VP.n8 161.3
R2898 VP.n60 VP.n0 161.3
R2899 VP.n59 VP.n58 161.3
R2900 VP.n57 VP.n1 161.3
R2901 VP.n56 VP.n55 161.3
R2902 VP.n53 VP.n2 161.3
R2903 VP.n52 VP.n51 161.3
R2904 VP.n50 VP.n3 161.3
R2905 VP.n49 VP.n48 161.3
R2906 VP.n47 VP.n4 161.3
R2907 VP.n46 VP.n45 161.3
R2908 VP.n44 VP.n5 161.3
R2909 VP.n43 VP.n42 161.3
R2910 VP.n40 VP.n6 161.3
R2911 VP.n39 VP.n38 161.3
R2912 VP.n37 VP.n7 161.3
R2913 VP.n40 VP.n39 56.5193
R2914 VP.n59 VP.n1 56.5193
R2915 VP.n31 VP.n9 56.5193
R2916 VP.n36 VP.n34 51.9096
R2917 VP.n15 VP.n14 49.6167
R2918 VP.n47 VP.n46 48.2635
R2919 VP.n52 VP.n3 48.2635
R2920 VP.n24 VP.n11 48.2635
R2921 VP.n19 VP.n18 48.2635
R2922 VP.n46 VP.n5 32.7233
R2923 VP.n53 VP.n52 32.7233
R2924 VP.n25 VP.n24 32.7233
R2925 VP.n18 VP.n13 32.7233
R2926 VP.n39 VP.n7 24.4675
R2927 VP.n42 VP.n40 24.4675
R2928 VP.n48 VP.n47 24.4675
R2929 VP.n48 VP.n3 24.4675
R2930 VP.n55 VP.n1 24.4675
R2931 VP.n60 VP.n59 24.4675
R2932 VP.n32 VP.n31 24.4675
R2933 VP.n27 VP.n9 24.4675
R2934 VP.n20 VP.n19 24.4675
R2935 VP.n20 VP.n11 24.4675
R2936 VP.n16 VP.n15 17.9026
R2937 VP.n41 VP.n5 16.6381
R2938 VP.n54 VP.n53 16.6381
R2939 VP.n26 VP.n25 16.6381
R2940 VP.n14 VP.n13 16.6381
R2941 VP.n35 VP.n7 8.80862
R2942 VP.n61 VP.n60 8.80862
R2943 VP.n33 VP.n32 8.80862
R2944 VP.n42 VP.n41 7.82994
R2945 VP.n55 VP.n54 7.82994
R2946 VP.n27 VP.n26 7.82994
R2947 VP.n17 VP.n16 0.189894
R2948 VP.n17 VP.n12 0.189894
R2949 VP.n21 VP.n12 0.189894
R2950 VP.n22 VP.n21 0.189894
R2951 VP.n23 VP.n22 0.189894
R2952 VP.n23 VP.n10 0.189894
R2953 VP.n28 VP.n10 0.189894
R2954 VP.n29 VP.n28 0.189894
R2955 VP.n30 VP.n29 0.189894
R2956 VP.n30 VP.n8 0.189894
R2957 VP.n34 VP.n8 0.189894
R2958 VP.n37 VP.n36 0.189894
R2959 VP.n38 VP.n37 0.189894
R2960 VP.n38 VP.n6 0.189894
R2961 VP.n43 VP.n6 0.189894
R2962 VP.n44 VP.n43 0.189894
R2963 VP.n45 VP.n44 0.189894
R2964 VP.n45 VP.n4 0.189894
R2965 VP.n49 VP.n4 0.189894
R2966 VP.n50 VP.n49 0.189894
R2967 VP.n51 VP.n50 0.189894
R2968 VP.n51 VP.n2 0.189894
R2969 VP.n56 VP.n2 0.189894
R2970 VP.n57 VP.n56 0.189894
R2971 VP.n58 VP.n57 0.189894
R2972 VP.n58 VP.n0 0.189894
R2973 VP.n62 VP.n0 0.189894
R2974 VP VP.n62 0.0516364
R2975 VDD1.n96 VDD1.n0 289.615
R2976 VDD1.n199 VDD1.n103 289.615
R2977 VDD1.n97 VDD1.n96 185
R2978 VDD1.n95 VDD1.n94 185
R2979 VDD1.n4 VDD1.n3 185
R2980 VDD1.n89 VDD1.n88 185
R2981 VDD1.n87 VDD1.n86 185
R2982 VDD1.n8 VDD1.n7 185
R2983 VDD1.n81 VDD1.n80 185
R2984 VDD1.n79 VDD1.n10 185
R2985 VDD1.n78 VDD1.n77 185
R2986 VDD1.n13 VDD1.n11 185
R2987 VDD1.n72 VDD1.n71 185
R2988 VDD1.n70 VDD1.n69 185
R2989 VDD1.n17 VDD1.n16 185
R2990 VDD1.n64 VDD1.n63 185
R2991 VDD1.n62 VDD1.n61 185
R2992 VDD1.n21 VDD1.n20 185
R2993 VDD1.n56 VDD1.n55 185
R2994 VDD1.n54 VDD1.n53 185
R2995 VDD1.n25 VDD1.n24 185
R2996 VDD1.n48 VDD1.n47 185
R2997 VDD1.n46 VDD1.n45 185
R2998 VDD1.n29 VDD1.n28 185
R2999 VDD1.n40 VDD1.n39 185
R3000 VDD1.n38 VDD1.n37 185
R3001 VDD1.n33 VDD1.n32 185
R3002 VDD1.n135 VDD1.n134 185
R3003 VDD1.n140 VDD1.n139 185
R3004 VDD1.n142 VDD1.n141 185
R3005 VDD1.n131 VDD1.n130 185
R3006 VDD1.n148 VDD1.n147 185
R3007 VDD1.n150 VDD1.n149 185
R3008 VDD1.n127 VDD1.n126 185
R3009 VDD1.n156 VDD1.n155 185
R3010 VDD1.n158 VDD1.n157 185
R3011 VDD1.n123 VDD1.n122 185
R3012 VDD1.n164 VDD1.n163 185
R3013 VDD1.n166 VDD1.n165 185
R3014 VDD1.n119 VDD1.n118 185
R3015 VDD1.n172 VDD1.n171 185
R3016 VDD1.n174 VDD1.n173 185
R3017 VDD1.n115 VDD1.n114 185
R3018 VDD1.n181 VDD1.n180 185
R3019 VDD1.n182 VDD1.n113 185
R3020 VDD1.n184 VDD1.n183 185
R3021 VDD1.n111 VDD1.n110 185
R3022 VDD1.n190 VDD1.n189 185
R3023 VDD1.n192 VDD1.n191 185
R3024 VDD1.n107 VDD1.n106 185
R3025 VDD1.n198 VDD1.n197 185
R3026 VDD1.n200 VDD1.n199 185
R3027 VDD1.n34 VDD1.t0 147.659
R3028 VDD1.n136 VDD1.t6 147.659
R3029 VDD1.n96 VDD1.n95 104.615
R3030 VDD1.n95 VDD1.n3 104.615
R3031 VDD1.n88 VDD1.n3 104.615
R3032 VDD1.n88 VDD1.n87 104.615
R3033 VDD1.n87 VDD1.n7 104.615
R3034 VDD1.n80 VDD1.n7 104.615
R3035 VDD1.n80 VDD1.n79 104.615
R3036 VDD1.n79 VDD1.n78 104.615
R3037 VDD1.n78 VDD1.n11 104.615
R3038 VDD1.n71 VDD1.n11 104.615
R3039 VDD1.n71 VDD1.n70 104.615
R3040 VDD1.n70 VDD1.n16 104.615
R3041 VDD1.n63 VDD1.n16 104.615
R3042 VDD1.n63 VDD1.n62 104.615
R3043 VDD1.n62 VDD1.n20 104.615
R3044 VDD1.n55 VDD1.n20 104.615
R3045 VDD1.n55 VDD1.n54 104.615
R3046 VDD1.n54 VDD1.n24 104.615
R3047 VDD1.n47 VDD1.n24 104.615
R3048 VDD1.n47 VDD1.n46 104.615
R3049 VDD1.n46 VDD1.n28 104.615
R3050 VDD1.n39 VDD1.n28 104.615
R3051 VDD1.n39 VDD1.n38 104.615
R3052 VDD1.n38 VDD1.n32 104.615
R3053 VDD1.n140 VDD1.n134 104.615
R3054 VDD1.n141 VDD1.n140 104.615
R3055 VDD1.n141 VDD1.n130 104.615
R3056 VDD1.n148 VDD1.n130 104.615
R3057 VDD1.n149 VDD1.n148 104.615
R3058 VDD1.n149 VDD1.n126 104.615
R3059 VDD1.n156 VDD1.n126 104.615
R3060 VDD1.n157 VDD1.n156 104.615
R3061 VDD1.n157 VDD1.n122 104.615
R3062 VDD1.n164 VDD1.n122 104.615
R3063 VDD1.n165 VDD1.n164 104.615
R3064 VDD1.n165 VDD1.n118 104.615
R3065 VDD1.n172 VDD1.n118 104.615
R3066 VDD1.n173 VDD1.n172 104.615
R3067 VDD1.n173 VDD1.n114 104.615
R3068 VDD1.n181 VDD1.n114 104.615
R3069 VDD1.n182 VDD1.n181 104.615
R3070 VDD1.n183 VDD1.n182 104.615
R3071 VDD1.n183 VDD1.n110 104.615
R3072 VDD1.n190 VDD1.n110 104.615
R3073 VDD1.n191 VDD1.n190 104.615
R3074 VDD1.n191 VDD1.n106 104.615
R3075 VDD1.n198 VDD1.n106 104.615
R3076 VDD1.n199 VDD1.n198 104.615
R3077 VDD1.n207 VDD1.n206 63.9158
R3078 VDD1.n102 VDD1.n101 62.7816
R3079 VDD1.n209 VDD1.n208 62.7814
R3080 VDD1.n205 VDD1.n204 62.7814
R3081 VDD1.n102 VDD1.n100 52.5837
R3082 VDD1.n205 VDD1.n203 52.5837
R3083 VDD1.t0 VDD1.n32 52.3082
R3084 VDD1.t6 VDD1.n134 52.3082
R3085 VDD1.n209 VDD1.n207 48.4449
R3086 VDD1.n34 VDD1.n33 15.6677
R3087 VDD1.n136 VDD1.n135 15.6677
R3088 VDD1.n81 VDD1.n10 13.1884
R3089 VDD1.n184 VDD1.n113 13.1884
R3090 VDD1.n82 VDD1.n8 12.8005
R3091 VDD1.n77 VDD1.n12 12.8005
R3092 VDD1.n37 VDD1.n36 12.8005
R3093 VDD1.n139 VDD1.n138 12.8005
R3094 VDD1.n180 VDD1.n179 12.8005
R3095 VDD1.n185 VDD1.n111 12.8005
R3096 VDD1.n86 VDD1.n85 12.0247
R3097 VDD1.n76 VDD1.n13 12.0247
R3098 VDD1.n40 VDD1.n31 12.0247
R3099 VDD1.n142 VDD1.n133 12.0247
R3100 VDD1.n178 VDD1.n115 12.0247
R3101 VDD1.n189 VDD1.n188 12.0247
R3102 VDD1.n89 VDD1.n6 11.249
R3103 VDD1.n73 VDD1.n72 11.249
R3104 VDD1.n41 VDD1.n29 11.249
R3105 VDD1.n143 VDD1.n131 11.249
R3106 VDD1.n175 VDD1.n174 11.249
R3107 VDD1.n192 VDD1.n109 11.249
R3108 VDD1.n90 VDD1.n4 10.4732
R3109 VDD1.n69 VDD1.n15 10.4732
R3110 VDD1.n45 VDD1.n44 10.4732
R3111 VDD1.n147 VDD1.n146 10.4732
R3112 VDD1.n171 VDD1.n117 10.4732
R3113 VDD1.n193 VDD1.n107 10.4732
R3114 VDD1.n94 VDD1.n93 9.69747
R3115 VDD1.n68 VDD1.n17 9.69747
R3116 VDD1.n48 VDD1.n27 9.69747
R3117 VDD1.n150 VDD1.n129 9.69747
R3118 VDD1.n170 VDD1.n119 9.69747
R3119 VDD1.n197 VDD1.n196 9.69747
R3120 VDD1.n100 VDD1.n99 9.45567
R3121 VDD1.n203 VDD1.n202 9.45567
R3122 VDD1.n60 VDD1.n59 9.3005
R3123 VDD1.n19 VDD1.n18 9.3005
R3124 VDD1.n66 VDD1.n65 9.3005
R3125 VDD1.n68 VDD1.n67 9.3005
R3126 VDD1.n15 VDD1.n14 9.3005
R3127 VDD1.n74 VDD1.n73 9.3005
R3128 VDD1.n76 VDD1.n75 9.3005
R3129 VDD1.n12 VDD1.n9 9.3005
R3130 VDD1.n99 VDD1.n98 9.3005
R3131 VDD1.n2 VDD1.n1 9.3005
R3132 VDD1.n93 VDD1.n92 9.3005
R3133 VDD1.n91 VDD1.n90 9.3005
R3134 VDD1.n6 VDD1.n5 9.3005
R3135 VDD1.n85 VDD1.n84 9.3005
R3136 VDD1.n83 VDD1.n82 9.3005
R3137 VDD1.n58 VDD1.n57 9.3005
R3138 VDD1.n23 VDD1.n22 9.3005
R3139 VDD1.n52 VDD1.n51 9.3005
R3140 VDD1.n50 VDD1.n49 9.3005
R3141 VDD1.n27 VDD1.n26 9.3005
R3142 VDD1.n44 VDD1.n43 9.3005
R3143 VDD1.n42 VDD1.n41 9.3005
R3144 VDD1.n31 VDD1.n30 9.3005
R3145 VDD1.n36 VDD1.n35 9.3005
R3146 VDD1.n202 VDD1.n201 9.3005
R3147 VDD1.n105 VDD1.n104 9.3005
R3148 VDD1.n196 VDD1.n195 9.3005
R3149 VDD1.n194 VDD1.n193 9.3005
R3150 VDD1.n109 VDD1.n108 9.3005
R3151 VDD1.n188 VDD1.n187 9.3005
R3152 VDD1.n186 VDD1.n185 9.3005
R3153 VDD1.n125 VDD1.n124 9.3005
R3154 VDD1.n154 VDD1.n153 9.3005
R3155 VDD1.n152 VDD1.n151 9.3005
R3156 VDD1.n129 VDD1.n128 9.3005
R3157 VDD1.n146 VDD1.n145 9.3005
R3158 VDD1.n144 VDD1.n143 9.3005
R3159 VDD1.n133 VDD1.n132 9.3005
R3160 VDD1.n138 VDD1.n137 9.3005
R3161 VDD1.n160 VDD1.n159 9.3005
R3162 VDD1.n162 VDD1.n161 9.3005
R3163 VDD1.n121 VDD1.n120 9.3005
R3164 VDD1.n168 VDD1.n167 9.3005
R3165 VDD1.n170 VDD1.n169 9.3005
R3166 VDD1.n117 VDD1.n116 9.3005
R3167 VDD1.n176 VDD1.n175 9.3005
R3168 VDD1.n178 VDD1.n177 9.3005
R3169 VDD1.n179 VDD1.n112 9.3005
R3170 VDD1.n97 VDD1.n2 8.92171
R3171 VDD1.n65 VDD1.n64 8.92171
R3172 VDD1.n49 VDD1.n25 8.92171
R3173 VDD1.n151 VDD1.n127 8.92171
R3174 VDD1.n167 VDD1.n166 8.92171
R3175 VDD1.n200 VDD1.n105 8.92171
R3176 VDD1.n98 VDD1.n0 8.14595
R3177 VDD1.n61 VDD1.n19 8.14595
R3178 VDD1.n53 VDD1.n52 8.14595
R3179 VDD1.n155 VDD1.n154 8.14595
R3180 VDD1.n163 VDD1.n121 8.14595
R3181 VDD1.n201 VDD1.n103 8.14595
R3182 VDD1.n60 VDD1.n21 7.3702
R3183 VDD1.n56 VDD1.n23 7.3702
R3184 VDD1.n158 VDD1.n125 7.3702
R3185 VDD1.n162 VDD1.n123 7.3702
R3186 VDD1.n57 VDD1.n21 6.59444
R3187 VDD1.n57 VDD1.n56 6.59444
R3188 VDD1.n159 VDD1.n158 6.59444
R3189 VDD1.n159 VDD1.n123 6.59444
R3190 VDD1.n100 VDD1.n0 5.81868
R3191 VDD1.n61 VDD1.n60 5.81868
R3192 VDD1.n53 VDD1.n23 5.81868
R3193 VDD1.n155 VDD1.n125 5.81868
R3194 VDD1.n163 VDD1.n162 5.81868
R3195 VDD1.n203 VDD1.n103 5.81868
R3196 VDD1.n98 VDD1.n97 5.04292
R3197 VDD1.n64 VDD1.n19 5.04292
R3198 VDD1.n52 VDD1.n25 5.04292
R3199 VDD1.n154 VDD1.n127 5.04292
R3200 VDD1.n166 VDD1.n121 5.04292
R3201 VDD1.n201 VDD1.n200 5.04292
R3202 VDD1.n35 VDD1.n34 4.38563
R3203 VDD1.n137 VDD1.n136 4.38563
R3204 VDD1.n94 VDD1.n2 4.26717
R3205 VDD1.n65 VDD1.n17 4.26717
R3206 VDD1.n49 VDD1.n48 4.26717
R3207 VDD1.n151 VDD1.n150 4.26717
R3208 VDD1.n167 VDD1.n119 4.26717
R3209 VDD1.n197 VDD1.n105 4.26717
R3210 VDD1.n93 VDD1.n4 3.49141
R3211 VDD1.n69 VDD1.n68 3.49141
R3212 VDD1.n45 VDD1.n27 3.49141
R3213 VDD1.n147 VDD1.n129 3.49141
R3214 VDD1.n171 VDD1.n170 3.49141
R3215 VDD1.n196 VDD1.n107 3.49141
R3216 VDD1.n90 VDD1.n89 2.71565
R3217 VDD1.n72 VDD1.n15 2.71565
R3218 VDD1.n44 VDD1.n29 2.71565
R3219 VDD1.n146 VDD1.n131 2.71565
R3220 VDD1.n174 VDD1.n117 2.71565
R3221 VDD1.n193 VDD1.n192 2.71565
R3222 VDD1.n86 VDD1.n6 1.93989
R3223 VDD1.n73 VDD1.n13 1.93989
R3224 VDD1.n41 VDD1.n40 1.93989
R3225 VDD1.n143 VDD1.n142 1.93989
R3226 VDD1.n175 VDD1.n115 1.93989
R3227 VDD1.n189 VDD1.n109 1.93989
R3228 VDD1.n85 VDD1.n8 1.16414
R3229 VDD1.n77 VDD1.n76 1.16414
R3230 VDD1.n37 VDD1.n31 1.16414
R3231 VDD1.n139 VDD1.n133 1.16414
R3232 VDD1.n180 VDD1.n178 1.16414
R3233 VDD1.n188 VDD1.n111 1.16414
R3234 VDD1 VDD1.n209 1.13197
R3235 VDD1.n208 VDD1.t7 1.07952
R3236 VDD1.n208 VDD1.t4 1.07952
R3237 VDD1.n101 VDD1.t8 1.07952
R3238 VDD1.n101 VDD1.t9 1.07952
R3239 VDD1.n206 VDD1.t2 1.07952
R3240 VDD1.n206 VDD1.t1 1.07952
R3241 VDD1.n204 VDD1.t5 1.07952
R3242 VDD1.n204 VDD1.t3 1.07952
R3243 VDD1 VDD1.n102 0.455241
R3244 VDD1.n82 VDD1.n81 0.388379
R3245 VDD1.n12 VDD1.n10 0.388379
R3246 VDD1.n36 VDD1.n33 0.388379
R3247 VDD1.n138 VDD1.n135 0.388379
R3248 VDD1.n179 VDD1.n113 0.388379
R3249 VDD1.n185 VDD1.n184 0.388379
R3250 VDD1.n207 VDD1.n205 0.341706
R3251 VDD1.n99 VDD1.n1 0.155672
R3252 VDD1.n92 VDD1.n1 0.155672
R3253 VDD1.n92 VDD1.n91 0.155672
R3254 VDD1.n91 VDD1.n5 0.155672
R3255 VDD1.n84 VDD1.n5 0.155672
R3256 VDD1.n84 VDD1.n83 0.155672
R3257 VDD1.n83 VDD1.n9 0.155672
R3258 VDD1.n75 VDD1.n9 0.155672
R3259 VDD1.n75 VDD1.n74 0.155672
R3260 VDD1.n74 VDD1.n14 0.155672
R3261 VDD1.n67 VDD1.n14 0.155672
R3262 VDD1.n67 VDD1.n66 0.155672
R3263 VDD1.n66 VDD1.n18 0.155672
R3264 VDD1.n59 VDD1.n18 0.155672
R3265 VDD1.n59 VDD1.n58 0.155672
R3266 VDD1.n58 VDD1.n22 0.155672
R3267 VDD1.n51 VDD1.n22 0.155672
R3268 VDD1.n51 VDD1.n50 0.155672
R3269 VDD1.n50 VDD1.n26 0.155672
R3270 VDD1.n43 VDD1.n26 0.155672
R3271 VDD1.n43 VDD1.n42 0.155672
R3272 VDD1.n42 VDD1.n30 0.155672
R3273 VDD1.n35 VDD1.n30 0.155672
R3274 VDD1.n137 VDD1.n132 0.155672
R3275 VDD1.n144 VDD1.n132 0.155672
R3276 VDD1.n145 VDD1.n144 0.155672
R3277 VDD1.n145 VDD1.n128 0.155672
R3278 VDD1.n152 VDD1.n128 0.155672
R3279 VDD1.n153 VDD1.n152 0.155672
R3280 VDD1.n153 VDD1.n124 0.155672
R3281 VDD1.n160 VDD1.n124 0.155672
R3282 VDD1.n161 VDD1.n160 0.155672
R3283 VDD1.n161 VDD1.n120 0.155672
R3284 VDD1.n168 VDD1.n120 0.155672
R3285 VDD1.n169 VDD1.n168 0.155672
R3286 VDD1.n169 VDD1.n116 0.155672
R3287 VDD1.n176 VDD1.n116 0.155672
R3288 VDD1.n177 VDD1.n176 0.155672
R3289 VDD1.n177 VDD1.n112 0.155672
R3290 VDD1.n186 VDD1.n112 0.155672
R3291 VDD1.n187 VDD1.n186 0.155672
R3292 VDD1.n187 VDD1.n108 0.155672
R3293 VDD1.n194 VDD1.n108 0.155672
R3294 VDD1.n195 VDD1.n194 0.155672
R3295 VDD1.n195 VDD1.n104 0.155672
R3296 VDD1.n202 VDD1.n104 0.155672
C0 VN VDD2 13.933599f
C1 VDD1 VN 0.15085f
C2 VP VN 7.96785f
C3 VTAIL VDD2 14.867101f
C4 VTAIL VDD1 14.8274f
C5 VDD1 VDD2 1.46678f
C6 VTAIL VP 13.878599f
C7 VP VDD2 0.445339f
C8 VDD1 VP 14.2225f
C9 VTAIL VN 13.863999f
C10 VDD2 B 7.05859f
C11 VDD1 B 7.031467f
C12 VTAIL B 9.741656f
C13 VN B 13.66369f
C14 VP B 11.830511f
C15 VDD1.n0 B 0.033205f
C16 VDD1.n1 B 0.022439f
C17 VDD1.n2 B 0.012058f
C18 VDD1.n3 B 0.0285f
C19 VDD1.n4 B 0.012767f
C20 VDD1.n5 B 0.022439f
C21 VDD1.n6 B 0.012058f
C22 VDD1.n7 B 0.0285f
C23 VDD1.n8 B 0.012767f
C24 VDD1.n9 B 0.022439f
C25 VDD1.n10 B 0.012412f
C26 VDD1.n11 B 0.0285f
C27 VDD1.n12 B 0.012058f
C28 VDD1.n13 B 0.012767f
C29 VDD1.n14 B 0.022439f
C30 VDD1.n15 B 0.012058f
C31 VDD1.n16 B 0.0285f
C32 VDD1.n17 B 0.012767f
C33 VDD1.n18 B 0.022439f
C34 VDD1.n19 B 0.012058f
C35 VDD1.n20 B 0.0285f
C36 VDD1.n21 B 0.012767f
C37 VDD1.n22 B 0.022439f
C38 VDD1.n23 B 0.012058f
C39 VDD1.n24 B 0.0285f
C40 VDD1.n25 B 0.012767f
C41 VDD1.n26 B 0.022439f
C42 VDD1.n27 B 0.012058f
C43 VDD1.n28 B 0.0285f
C44 VDD1.n29 B 0.012767f
C45 VDD1.n30 B 0.022439f
C46 VDD1.n31 B 0.012058f
C47 VDD1.n32 B 0.021375f
C48 VDD1.n33 B 0.016836f
C49 VDD1.t0 B 0.04725f
C50 VDD1.n34 B 0.165197f
C51 VDD1.n35 B 1.8044f
C52 VDD1.n36 B 0.012058f
C53 VDD1.n37 B 0.012767f
C54 VDD1.n38 B 0.0285f
C55 VDD1.n39 B 0.0285f
C56 VDD1.n40 B 0.012767f
C57 VDD1.n41 B 0.012058f
C58 VDD1.n42 B 0.022439f
C59 VDD1.n43 B 0.022439f
C60 VDD1.n44 B 0.012058f
C61 VDD1.n45 B 0.012767f
C62 VDD1.n46 B 0.0285f
C63 VDD1.n47 B 0.0285f
C64 VDD1.n48 B 0.012767f
C65 VDD1.n49 B 0.012058f
C66 VDD1.n50 B 0.022439f
C67 VDD1.n51 B 0.022439f
C68 VDD1.n52 B 0.012058f
C69 VDD1.n53 B 0.012767f
C70 VDD1.n54 B 0.0285f
C71 VDD1.n55 B 0.0285f
C72 VDD1.n56 B 0.012767f
C73 VDD1.n57 B 0.012058f
C74 VDD1.n58 B 0.022439f
C75 VDD1.n59 B 0.022439f
C76 VDD1.n60 B 0.012058f
C77 VDD1.n61 B 0.012767f
C78 VDD1.n62 B 0.0285f
C79 VDD1.n63 B 0.0285f
C80 VDD1.n64 B 0.012767f
C81 VDD1.n65 B 0.012058f
C82 VDD1.n66 B 0.022439f
C83 VDD1.n67 B 0.022439f
C84 VDD1.n68 B 0.012058f
C85 VDD1.n69 B 0.012767f
C86 VDD1.n70 B 0.0285f
C87 VDD1.n71 B 0.0285f
C88 VDD1.n72 B 0.012767f
C89 VDD1.n73 B 0.012058f
C90 VDD1.n74 B 0.022439f
C91 VDD1.n75 B 0.022439f
C92 VDD1.n76 B 0.012058f
C93 VDD1.n77 B 0.012767f
C94 VDD1.n78 B 0.0285f
C95 VDD1.n79 B 0.0285f
C96 VDD1.n80 B 0.0285f
C97 VDD1.n81 B 0.012412f
C98 VDD1.n82 B 0.012058f
C99 VDD1.n83 B 0.022439f
C100 VDD1.n84 B 0.022439f
C101 VDD1.n85 B 0.012058f
C102 VDD1.n86 B 0.012767f
C103 VDD1.n87 B 0.0285f
C104 VDD1.n88 B 0.0285f
C105 VDD1.n89 B 0.012767f
C106 VDD1.n90 B 0.012058f
C107 VDD1.n91 B 0.022439f
C108 VDD1.n92 B 0.022439f
C109 VDD1.n93 B 0.012058f
C110 VDD1.n94 B 0.012767f
C111 VDD1.n95 B 0.0285f
C112 VDD1.n96 B 0.064642f
C113 VDD1.n97 B 0.012767f
C114 VDD1.n98 B 0.012058f
C115 VDD1.n99 B 0.055238f
C116 VDD1.n100 B 0.056863f
C117 VDD1.t8 B 0.325377f
C118 VDD1.t9 B 0.325377f
C119 VDD1.n101 B 2.96847f
C120 VDD1.n102 B 0.487205f
C121 VDD1.n103 B 0.033205f
C122 VDD1.n104 B 0.022439f
C123 VDD1.n105 B 0.012058f
C124 VDD1.n106 B 0.0285f
C125 VDD1.n107 B 0.012767f
C126 VDD1.n108 B 0.022439f
C127 VDD1.n109 B 0.012058f
C128 VDD1.n110 B 0.0285f
C129 VDD1.n111 B 0.012767f
C130 VDD1.n112 B 0.022439f
C131 VDD1.n113 B 0.012412f
C132 VDD1.n114 B 0.0285f
C133 VDD1.n115 B 0.012767f
C134 VDD1.n116 B 0.022439f
C135 VDD1.n117 B 0.012058f
C136 VDD1.n118 B 0.0285f
C137 VDD1.n119 B 0.012767f
C138 VDD1.n120 B 0.022439f
C139 VDD1.n121 B 0.012058f
C140 VDD1.n122 B 0.0285f
C141 VDD1.n123 B 0.012767f
C142 VDD1.n124 B 0.022439f
C143 VDD1.n125 B 0.012058f
C144 VDD1.n126 B 0.0285f
C145 VDD1.n127 B 0.012767f
C146 VDD1.n128 B 0.022439f
C147 VDD1.n129 B 0.012058f
C148 VDD1.n130 B 0.0285f
C149 VDD1.n131 B 0.012767f
C150 VDD1.n132 B 0.022439f
C151 VDD1.n133 B 0.012058f
C152 VDD1.n134 B 0.021375f
C153 VDD1.n135 B 0.016836f
C154 VDD1.t6 B 0.04725f
C155 VDD1.n136 B 0.165197f
C156 VDD1.n137 B 1.80439f
C157 VDD1.n138 B 0.012058f
C158 VDD1.n139 B 0.012767f
C159 VDD1.n140 B 0.0285f
C160 VDD1.n141 B 0.0285f
C161 VDD1.n142 B 0.012767f
C162 VDD1.n143 B 0.012058f
C163 VDD1.n144 B 0.022439f
C164 VDD1.n145 B 0.022439f
C165 VDD1.n146 B 0.012058f
C166 VDD1.n147 B 0.012767f
C167 VDD1.n148 B 0.0285f
C168 VDD1.n149 B 0.0285f
C169 VDD1.n150 B 0.012767f
C170 VDD1.n151 B 0.012058f
C171 VDD1.n152 B 0.022439f
C172 VDD1.n153 B 0.022439f
C173 VDD1.n154 B 0.012058f
C174 VDD1.n155 B 0.012767f
C175 VDD1.n156 B 0.0285f
C176 VDD1.n157 B 0.0285f
C177 VDD1.n158 B 0.012767f
C178 VDD1.n159 B 0.012058f
C179 VDD1.n160 B 0.022439f
C180 VDD1.n161 B 0.022439f
C181 VDD1.n162 B 0.012058f
C182 VDD1.n163 B 0.012767f
C183 VDD1.n164 B 0.0285f
C184 VDD1.n165 B 0.0285f
C185 VDD1.n166 B 0.012767f
C186 VDD1.n167 B 0.012058f
C187 VDD1.n168 B 0.022439f
C188 VDD1.n169 B 0.022439f
C189 VDD1.n170 B 0.012058f
C190 VDD1.n171 B 0.012767f
C191 VDD1.n172 B 0.0285f
C192 VDD1.n173 B 0.0285f
C193 VDD1.n174 B 0.012767f
C194 VDD1.n175 B 0.012058f
C195 VDD1.n176 B 0.022439f
C196 VDD1.n177 B 0.022439f
C197 VDD1.n178 B 0.012058f
C198 VDD1.n179 B 0.012058f
C199 VDD1.n180 B 0.012767f
C200 VDD1.n181 B 0.0285f
C201 VDD1.n182 B 0.0285f
C202 VDD1.n183 B 0.0285f
C203 VDD1.n184 B 0.012412f
C204 VDD1.n185 B 0.012058f
C205 VDD1.n186 B 0.022439f
C206 VDD1.n187 B 0.022439f
C207 VDD1.n188 B 0.012058f
C208 VDD1.n189 B 0.012767f
C209 VDD1.n190 B 0.0285f
C210 VDD1.n191 B 0.0285f
C211 VDD1.n192 B 0.012767f
C212 VDD1.n193 B 0.012058f
C213 VDD1.n194 B 0.022439f
C214 VDD1.n195 B 0.022439f
C215 VDD1.n196 B 0.012058f
C216 VDD1.n197 B 0.012767f
C217 VDD1.n198 B 0.0285f
C218 VDD1.n199 B 0.064642f
C219 VDD1.n200 B 0.012767f
C220 VDD1.n201 B 0.012058f
C221 VDD1.n202 B 0.055238f
C222 VDD1.n203 B 0.056863f
C223 VDD1.t5 B 0.325377f
C224 VDD1.t3 B 0.325377f
C225 VDD1.n204 B 2.96846f
C226 VDD1.n205 B 0.48053f
C227 VDD1.t2 B 0.325377f
C228 VDD1.t1 B 0.325377f
C229 VDD1.n206 B 2.9754f
C230 VDD1.n207 B 2.53821f
C231 VDD1.t7 B 0.325377f
C232 VDD1.t4 B 0.325377f
C233 VDD1.n208 B 2.96846f
C234 VDD1.n209 B 2.87712f
C235 VP.n0 B 0.029373f
C236 VP.t8 B 2.23946f
C237 VP.n1 B 0.043698f
C238 VP.n2 B 0.029373f
C239 VP.t7 B 2.23946f
C240 VP.n3 B 0.055009f
C241 VP.n4 B 0.029373f
C242 VP.t6 B 2.23946f
C243 VP.n5 B 0.050594f
C244 VP.n6 B 0.029373f
C245 VP.n7 B 0.037447f
C246 VP.n8 B 0.029373f
C247 VP.t5 B 2.23946f
C248 VP.n9 B 0.043698f
C249 VP.n10 B 0.029373f
C250 VP.t2 B 2.23946f
C251 VP.n11 B 0.055009f
C252 VP.n12 B 0.029373f
C253 VP.t0 B 2.23946f
C254 VP.n13 B 0.050594f
C255 VP.t9 B 2.331f
C256 VP.t1 B 2.23946f
C257 VP.n14 B 0.846956f
C258 VP.n15 B 0.858129f
C259 VP.n16 B 0.185554f
C260 VP.n17 B 0.029373f
C261 VP.n18 B 0.026252f
C262 VP.n19 B 0.055009f
C263 VP.n20 B 0.815043f
C264 VP.n21 B 0.029373f
C265 VP.n22 B 0.029373f
C266 VP.n23 B 0.029373f
C267 VP.n24 B 0.026252f
C268 VP.n25 B 0.050594f
C269 VP.n26 B 0.787326f
C270 VP.n27 B 0.036366f
C271 VP.n28 B 0.029373f
C272 VP.n29 B 0.029373f
C273 VP.n30 B 0.029373f
C274 VP.n31 B 0.042061f
C275 VP.n32 B 0.037447f
C276 VP.n33 B 0.846588f
C277 VP.n34 B 1.69437f
C278 VP.t3 B 2.23946f
C279 VP.n35 B 0.846588f
C280 VP.n36 B 1.71471f
C281 VP.n37 B 0.029373f
C282 VP.n38 B 0.029373f
C283 VP.n39 B 0.042061f
C284 VP.n40 B 0.043698f
C285 VP.t4 B 2.23946f
C286 VP.n41 B 0.787326f
C287 VP.n42 B 0.036366f
C288 VP.n43 B 0.029373f
C289 VP.n44 B 0.029373f
C290 VP.n45 B 0.029373f
C291 VP.n46 B 0.026252f
C292 VP.n47 B 0.055009f
C293 VP.n48 B 0.815043f
C294 VP.n49 B 0.029373f
C295 VP.n50 B 0.029373f
C296 VP.n51 B 0.029373f
C297 VP.n52 B 0.026252f
C298 VP.n53 B 0.050594f
C299 VP.n54 B 0.787326f
C300 VP.n55 B 0.036366f
C301 VP.n56 B 0.029373f
C302 VP.n57 B 0.029373f
C303 VP.n58 B 0.029373f
C304 VP.n59 B 0.042061f
C305 VP.n60 B 0.037447f
C306 VP.n61 B 0.846588f
C307 VP.n62 B 0.028516f
C308 VDD2.n0 B 0.03307f
C309 VDD2.n1 B 0.022348f
C310 VDD2.n2 B 0.012009f
C311 VDD2.n3 B 0.028384f
C312 VDD2.n4 B 0.012715f
C313 VDD2.n5 B 0.022348f
C314 VDD2.n6 B 0.012009f
C315 VDD2.n7 B 0.028384f
C316 VDD2.n8 B 0.012715f
C317 VDD2.n9 B 0.022348f
C318 VDD2.n10 B 0.012362f
C319 VDD2.n11 B 0.028384f
C320 VDD2.n12 B 0.012715f
C321 VDD2.n13 B 0.022348f
C322 VDD2.n14 B 0.012009f
C323 VDD2.n15 B 0.028384f
C324 VDD2.n16 B 0.012715f
C325 VDD2.n17 B 0.022348f
C326 VDD2.n18 B 0.012009f
C327 VDD2.n19 B 0.028384f
C328 VDD2.n20 B 0.012715f
C329 VDD2.n21 B 0.022348f
C330 VDD2.n22 B 0.012009f
C331 VDD2.n23 B 0.028384f
C332 VDD2.n24 B 0.012715f
C333 VDD2.n25 B 0.022348f
C334 VDD2.n26 B 0.012009f
C335 VDD2.n27 B 0.028384f
C336 VDD2.n28 B 0.012715f
C337 VDD2.n29 B 0.022348f
C338 VDD2.n30 B 0.012009f
C339 VDD2.n31 B 0.021288f
C340 VDD2.n32 B 0.016767f
C341 VDD2.t4 B 0.047059f
C342 VDD2.n33 B 0.164528f
C343 VDD2.n34 B 1.79709f
C344 VDD2.n35 B 0.012009f
C345 VDD2.n36 B 0.012715f
C346 VDD2.n37 B 0.028384f
C347 VDD2.n38 B 0.028384f
C348 VDD2.n39 B 0.012715f
C349 VDD2.n40 B 0.012009f
C350 VDD2.n41 B 0.022348f
C351 VDD2.n42 B 0.022348f
C352 VDD2.n43 B 0.012009f
C353 VDD2.n44 B 0.012715f
C354 VDD2.n45 B 0.028384f
C355 VDD2.n46 B 0.028384f
C356 VDD2.n47 B 0.012715f
C357 VDD2.n48 B 0.012009f
C358 VDD2.n49 B 0.022348f
C359 VDD2.n50 B 0.022348f
C360 VDD2.n51 B 0.012009f
C361 VDD2.n52 B 0.012715f
C362 VDD2.n53 B 0.028384f
C363 VDD2.n54 B 0.028384f
C364 VDD2.n55 B 0.012715f
C365 VDD2.n56 B 0.012009f
C366 VDD2.n57 B 0.022348f
C367 VDD2.n58 B 0.022348f
C368 VDD2.n59 B 0.012009f
C369 VDD2.n60 B 0.012715f
C370 VDD2.n61 B 0.028384f
C371 VDD2.n62 B 0.028384f
C372 VDD2.n63 B 0.012715f
C373 VDD2.n64 B 0.012009f
C374 VDD2.n65 B 0.022348f
C375 VDD2.n66 B 0.022348f
C376 VDD2.n67 B 0.012009f
C377 VDD2.n68 B 0.012715f
C378 VDD2.n69 B 0.028384f
C379 VDD2.n70 B 0.028384f
C380 VDD2.n71 B 0.012715f
C381 VDD2.n72 B 0.012009f
C382 VDD2.n73 B 0.022348f
C383 VDD2.n74 B 0.022348f
C384 VDD2.n75 B 0.012009f
C385 VDD2.n76 B 0.012009f
C386 VDD2.n77 B 0.012715f
C387 VDD2.n78 B 0.028384f
C388 VDD2.n79 B 0.028384f
C389 VDD2.n80 B 0.028384f
C390 VDD2.n81 B 0.012362f
C391 VDD2.n82 B 0.012009f
C392 VDD2.n83 B 0.022348f
C393 VDD2.n84 B 0.022348f
C394 VDD2.n85 B 0.012009f
C395 VDD2.n86 B 0.012715f
C396 VDD2.n87 B 0.028384f
C397 VDD2.n88 B 0.028384f
C398 VDD2.n89 B 0.012715f
C399 VDD2.n90 B 0.012009f
C400 VDD2.n91 B 0.022348f
C401 VDD2.n92 B 0.022348f
C402 VDD2.n93 B 0.012009f
C403 VDD2.n94 B 0.012715f
C404 VDD2.n95 B 0.028384f
C405 VDD2.n96 B 0.06438f
C406 VDD2.n97 B 0.012715f
C407 VDD2.n98 B 0.012009f
C408 VDD2.n99 B 0.055014f
C409 VDD2.n100 B 0.056633f
C410 VDD2.t5 B 0.324059f
C411 VDD2.t7 B 0.324059f
C412 VDD2.n101 B 2.95644f
C413 VDD2.n102 B 0.478584f
C414 VDD2.t8 B 0.324059f
C415 VDD2.t9 B 0.324059f
C416 VDD2.n103 B 2.96335f
C417 VDD2.n104 B 2.43906f
C418 VDD2.n105 B 0.03307f
C419 VDD2.n106 B 0.022348f
C420 VDD2.n107 B 0.012009f
C421 VDD2.n108 B 0.028384f
C422 VDD2.n109 B 0.012715f
C423 VDD2.n110 B 0.022348f
C424 VDD2.n111 B 0.012009f
C425 VDD2.n112 B 0.028384f
C426 VDD2.n113 B 0.012715f
C427 VDD2.n114 B 0.022348f
C428 VDD2.n115 B 0.012362f
C429 VDD2.n116 B 0.028384f
C430 VDD2.n117 B 0.012009f
C431 VDD2.n118 B 0.012715f
C432 VDD2.n119 B 0.022348f
C433 VDD2.n120 B 0.012009f
C434 VDD2.n121 B 0.028384f
C435 VDD2.n122 B 0.012715f
C436 VDD2.n123 B 0.022348f
C437 VDD2.n124 B 0.012009f
C438 VDD2.n125 B 0.028384f
C439 VDD2.n126 B 0.012715f
C440 VDD2.n127 B 0.022348f
C441 VDD2.n128 B 0.012009f
C442 VDD2.n129 B 0.028384f
C443 VDD2.n130 B 0.012715f
C444 VDD2.n131 B 0.022348f
C445 VDD2.n132 B 0.012009f
C446 VDD2.n133 B 0.028384f
C447 VDD2.n134 B 0.012715f
C448 VDD2.n135 B 0.022348f
C449 VDD2.n136 B 0.012009f
C450 VDD2.n137 B 0.021288f
C451 VDD2.n138 B 0.016767f
C452 VDD2.t3 B 0.047059f
C453 VDD2.n139 B 0.164528f
C454 VDD2.n140 B 1.79709f
C455 VDD2.n141 B 0.012009f
C456 VDD2.n142 B 0.012715f
C457 VDD2.n143 B 0.028384f
C458 VDD2.n144 B 0.028384f
C459 VDD2.n145 B 0.012715f
C460 VDD2.n146 B 0.012009f
C461 VDD2.n147 B 0.022348f
C462 VDD2.n148 B 0.022348f
C463 VDD2.n149 B 0.012009f
C464 VDD2.n150 B 0.012715f
C465 VDD2.n151 B 0.028384f
C466 VDD2.n152 B 0.028384f
C467 VDD2.n153 B 0.012715f
C468 VDD2.n154 B 0.012009f
C469 VDD2.n155 B 0.022348f
C470 VDD2.n156 B 0.022348f
C471 VDD2.n157 B 0.012009f
C472 VDD2.n158 B 0.012715f
C473 VDD2.n159 B 0.028384f
C474 VDD2.n160 B 0.028384f
C475 VDD2.n161 B 0.012715f
C476 VDD2.n162 B 0.012009f
C477 VDD2.n163 B 0.022348f
C478 VDD2.n164 B 0.022348f
C479 VDD2.n165 B 0.012009f
C480 VDD2.n166 B 0.012715f
C481 VDD2.n167 B 0.028384f
C482 VDD2.n168 B 0.028384f
C483 VDD2.n169 B 0.012715f
C484 VDD2.n170 B 0.012009f
C485 VDD2.n171 B 0.022348f
C486 VDD2.n172 B 0.022348f
C487 VDD2.n173 B 0.012009f
C488 VDD2.n174 B 0.012715f
C489 VDD2.n175 B 0.028384f
C490 VDD2.n176 B 0.028384f
C491 VDD2.n177 B 0.012715f
C492 VDD2.n178 B 0.012009f
C493 VDD2.n179 B 0.022348f
C494 VDD2.n180 B 0.022348f
C495 VDD2.n181 B 0.012009f
C496 VDD2.n182 B 0.012715f
C497 VDD2.n183 B 0.028384f
C498 VDD2.n184 B 0.028384f
C499 VDD2.n185 B 0.028384f
C500 VDD2.n186 B 0.012362f
C501 VDD2.n187 B 0.012009f
C502 VDD2.n188 B 0.022348f
C503 VDD2.n189 B 0.022348f
C504 VDD2.n190 B 0.012009f
C505 VDD2.n191 B 0.012715f
C506 VDD2.n192 B 0.028384f
C507 VDD2.n193 B 0.028384f
C508 VDD2.n194 B 0.012715f
C509 VDD2.n195 B 0.012009f
C510 VDD2.n196 B 0.022348f
C511 VDD2.n197 B 0.022348f
C512 VDD2.n198 B 0.012009f
C513 VDD2.n199 B 0.012715f
C514 VDD2.n200 B 0.028384f
C515 VDD2.n201 B 0.06438f
C516 VDD2.n202 B 0.012715f
C517 VDD2.n203 B 0.012009f
C518 VDD2.n204 B 0.055014f
C519 VDD2.n205 B 0.051831f
C520 VDD2.n206 B 2.64236f
C521 VDD2.t6 B 0.324059f
C522 VDD2.t1 B 0.324059f
C523 VDD2.n207 B 2.95645f
C524 VDD2.n208 B 0.330856f
C525 VDD2.t0 B 0.324059f
C526 VDD2.t2 B 0.324059f
C527 VDD2.n209 B 2.96332f
C528 VTAIL.t15 B 0.340728f
C529 VTAIL.t18 B 0.340728f
C530 VTAIL.n0 B 3.04018f
C531 VTAIL.n1 B 0.419853f
C532 VTAIL.n2 B 0.034771f
C533 VTAIL.n3 B 0.023497f
C534 VTAIL.n4 B 0.012626f
C535 VTAIL.n5 B 0.029844f
C536 VTAIL.n6 B 0.013369f
C537 VTAIL.n7 B 0.023497f
C538 VTAIL.n8 B 0.012626f
C539 VTAIL.n9 B 0.029844f
C540 VTAIL.n10 B 0.013369f
C541 VTAIL.n11 B 0.023497f
C542 VTAIL.n12 B 0.012998f
C543 VTAIL.n13 B 0.029844f
C544 VTAIL.n14 B 0.013369f
C545 VTAIL.n15 B 0.023497f
C546 VTAIL.n16 B 0.012626f
C547 VTAIL.n17 B 0.029844f
C548 VTAIL.n18 B 0.013369f
C549 VTAIL.n19 B 0.023497f
C550 VTAIL.n20 B 0.012626f
C551 VTAIL.n21 B 0.029844f
C552 VTAIL.n22 B 0.013369f
C553 VTAIL.n23 B 0.023497f
C554 VTAIL.n24 B 0.012626f
C555 VTAIL.n25 B 0.029844f
C556 VTAIL.n26 B 0.013369f
C557 VTAIL.n27 B 0.023497f
C558 VTAIL.n28 B 0.012626f
C559 VTAIL.n29 B 0.029844f
C560 VTAIL.n30 B 0.013369f
C561 VTAIL.n31 B 0.023497f
C562 VTAIL.n32 B 0.012626f
C563 VTAIL.n33 B 0.022383f
C564 VTAIL.n34 B 0.01763f
C565 VTAIL.t4 B 0.04948f
C566 VTAIL.n35 B 0.17299f
C567 VTAIL.n36 B 1.88952f
C568 VTAIL.n37 B 0.012626f
C569 VTAIL.n38 B 0.013369f
C570 VTAIL.n39 B 0.029844f
C571 VTAIL.n40 B 0.029844f
C572 VTAIL.n41 B 0.013369f
C573 VTAIL.n42 B 0.012626f
C574 VTAIL.n43 B 0.023497f
C575 VTAIL.n44 B 0.023497f
C576 VTAIL.n45 B 0.012626f
C577 VTAIL.n46 B 0.013369f
C578 VTAIL.n47 B 0.029844f
C579 VTAIL.n48 B 0.029844f
C580 VTAIL.n49 B 0.013369f
C581 VTAIL.n50 B 0.012626f
C582 VTAIL.n51 B 0.023497f
C583 VTAIL.n52 B 0.023497f
C584 VTAIL.n53 B 0.012626f
C585 VTAIL.n54 B 0.013369f
C586 VTAIL.n55 B 0.029844f
C587 VTAIL.n56 B 0.029844f
C588 VTAIL.n57 B 0.013369f
C589 VTAIL.n58 B 0.012626f
C590 VTAIL.n59 B 0.023497f
C591 VTAIL.n60 B 0.023497f
C592 VTAIL.n61 B 0.012626f
C593 VTAIL.n62 B 0.013369f
C594 VTAIL.n63 B 0.029844f
C595 VTAIL.n64 B 0.029844f
C596 VTAIL.n65 B 0.013369f
C597 VTAIL.n66 B 0.012626f
C598 VTAIL.n67 B 0.023497f
C599 VTAIL.n68 B 0.023497f
C600 VTAIL.n69 B 0.012626f
C601 VTAIL.n70 B 0.013369f
C602 VTAIL.n71 B 0.029844f
C603 VTAIL.n72 B 0.029844f
C604 VTAIL.n73 B 0.013369f
C605 VTAIL.n74 B 0.012626f
C606 VTAIL.n75 B 0.023497f
C607 VTAIL.n76 B 0.023497f
C608 VTAIL.n77 B 0.012626f
C609 VTAIL.n78 B 0.012626f
C610 VTAIL.n79 B 0.013369f
C611 VTAIL.n80 B 0.029844f
C612 VTAIL.n81 B 0.029844f
C613 VTAIL.n82 B 0.029844f
C614 VTAIL.n83 B 0.012998f
C615 VTAIL.n84 B 0.012626f
C616 VTAIL.n85 B 0.023497f
C617 VTAIL.n86 B 0.023497f
C618 VTAIL.n87 B 0.012626f
C619 VTAIL.n88 B 0.013369f
C620 VTAIL.n89 B 0.029844f
C621 VTAIL.n90 B 0.029844f
C622 VTAIL.n91 B 0.013369f
C623 VTAIL.n92 B 0.012626f
C624 VTAIL.n93 B 0.023497f
C625 VTAIL.n94 B 0.023497f
C626 VTAIL.n95 B 0.012626f
C627 VTAIL.n96 B 0.013369f
C628 VTAIL.n97 B 0.029844f
C629 VTAIL.n98 B 0.067692f
C630 VTAIL.n99 B 0.013369f
C631 VTAIL.n100 B 0.012626f
C632 VTAIL.n101 B 0.057844f
C633 VTAIL.n102 B 0.038299f
C634 VTAIL.n103 B 0.237783f
C635 VTAIL.t0 B 0.340728f
C636 VTAIL.t6 B 0.340728f
C637 VTAIL.n104 B 3.04018f
C638 VTAIL.n105 B 0.469947f
C639 VTAIL.t8 B 0.340728f
C640 VTAIL.t3 B 0.340728f
C641 VTAIL.n106 B 3.04018f
C642 VTAIL.n107 B 2.10694f
C643 VTAIL.t14 B 0.340728f
C644 VTAIL.t10 B 0.340728f
C645 VTAIL.n108 B 3.04019f
C646 VTAIL.n109 B 2.10692f
C647 VTAIL.t13 B 0.340728f
C648 VTAIL.t16 B 0.340728f
C649 VTAIL.n110 B 3.04019f
C650 VTAIL.n111 B 0.469934f
C651 VTAIL.n112 B 0.034771f
C652 VTAIL.n113 B 0.023497f
C653 VTAIL.n114 B 0.012626f
C654 VTAIL.n115 B 0.029844f
C655 VTAIL.n116 B 0.013369f
C656 VTAIL.n117 B 0.023497f
C657 VTAIL.n118 B 0.012626f
C658 VTAIL.n119 B 0.029844f
C659 VTAIL.n120 B 0.013369f
C660 VTAIL.n121 B 0.023497f
C661 VTAIL.n122 B 0.012998f
C662 VTAIL.n123 B 0.029844f
C663 VTAIL.n124 B 0.012626f
C664 VTAIL.n125 B 0.013369f
C665 VTAIL.n126 B 0.023497f
C666 VTAIL.n127 B 0.012626f
C667 VTAIL.n128 B 0.029844f
C668 VTAIL.n129 B 0.013369f
C669 VTAIL.n130 B 0.023497f
C670 VTAIL.n131 B 0.012626f
C671 VTAIL.n132 B 0.029844f
C672 VTAIL.n133 B 0.013369f
C673 VTAIL.n134 B 0.023497f
C674 VTAIL.n135 B 0.012626f
C675 VTAIL.n136 B 0.029844f
C676 VTAIL.n137 B 0.013369f
C677 VTAIL.n138 B 0.023497f
C678 VTAIL.n139 B 0.012626f
C679 VTAIL.n140 B 0.029844f
C680 VTAIL.n141 B 0.013369f
C681 VTAIL.n142 B 0.023497f
C682 VTAIL.n143 B 0.012626f
C683 VTAIL.n144 B 0.022383f
C684 VTAIL.n145 B 0.01763f
C685 VTAIL.t19 B 0.04948f
C686 VTAIL.n146 B 0.17299f
C687 VTAIL.n147 B 1.88952f
C688 VTAIL.n148 B 0.012626f
C689 VTAIL.n149 B 0.013369f
C690 VTAIL.n150 B 0.029844f
C691 VTAIL.n151 B 0.029844f
C692 VTAIL.n152 B 0.013369f
C693 VTAIL.n153 B 0.012626f
C694 VTAIL.n154 B 0.023497f
C695 VTAIL.n155 B 0.023497f
C696 VTAIL.n156 B 0.012626f
C697 VTAIL.n157 B 0.013369f
C698 VTAIL.n158 B 0.029844f
C699 VTAIL.n159 B 0.029844f
C700 VTAIL.n160 B 0.013369f
C701 VTAIL.n161 B 0.012626f
C702 VTAIL.n162 B 0.023497f
C703 VTAIL.n163 B 0.023497f
C704 VTAIL.n164 B 0.012626f
C705 VTAIL.n165 B 0.013369f
C706 VTAIL.n166 B 0.029844f
C707 VTAIL.n167 B 0.029844f
C708 VTAIL.n168 B 0.013369f
C709 VTAIL.n169 B 0.012626f
C710 VTAIL.n170 B 0.023497f
C711 VTAIL.n171 B 0.023497f
C712 VTAIL.n172 B 0.012626f
C713 VTAIL.n173 B 0.013369f
C714 VTAIL.n174 B 0.029844f
C715 VTAIL.n175 B 0.029844f
C716 VTAIL.n176 B 0.013369f
C717 VTAIL.n177 B 0.012626f
C718 VTAIL.n178 B 0.023497f
C719 VTAIL.n179 B 0.023497f
C720 VTAIL.n180 B 0.012626f
C721 VTAIL.n181 B 0.013369f
C722 VTAIL.n182 B 0.029844f
C723 VTAIL.n183 B 0.029844f
C724 VTAIL.n184 B 0.013369f
C725 VTAIL.n185 B 0.012626f
C726 VTAIL.n186 B 0.023497f
C727 VTAIL.n187 B 0.023497f
C728 VTAIL.n188 B 0.012626f
C729 VTAIL.n189 B 0.013369f
C730 VTAIL.n190 B 0.029844f
C731 VTAIL.n191 B 0.029844f
C732 VTAIL.n192 B 0.029844f
C733 VTAIL.n193 B 0.012998f
C734 VTAIL.n194 B 0.012626f
C735 VTAIL.n195 B 0.023497f
C736 VTAIL.n196 B 0.023497f
C737 VTAIL.n197 B 0.012626f
C738 VTAIL.n198 B 0.013369f
C739 VTAIL.n199 B 0.029844f
C740 VTAIL.n200 B 0.029844f
C741 VTAIL.n201 B 0.013369f
C742 VTAIL.n202 B 0.012626f
C743 VTAIL.n203 B 0.023497f
C744 VTAIL.n204 B 0.023497f
C745 VTAIL.n205 B 0.012626f
C746 VTAIL.n206 B 0.013369f
C747 VTAIL.n207 B 0.029844f
C748 VTAIL.n208 B 0.067692f
C749 VTAIL.n209 B 0.013369f
C750 VTAIL.n210 B 0.012626f
C751 VTAIL.n211 B 0.057844f
C752 VTAIL.n212 B 0.038299f
C753 VTAIL.n213 B 0.237783f
C754 VTAIL.t2 B 0.340728f
C755 VTAIL.t5 B 0.340728f
C756 VTAIL.n214 B 3.04019f
C757 VTAIL.n215 B 0.445458f
C758 VTAIL.t7 B 0.340728f
C759 VTAIL.t1 B 0.340728f
C760 VTAIL.n216 B 3.04019f
C761 VTAIL.n217 B 0.469934f
C762 VTAIL.n218 B 0.034771f
C763 VTAIL.n219 B 0.023497f
C764 VTAIL.n220 B 0.012626f
C765 VTAIL.n221 B 0.029844f
C766 VTAIL.n222 B 0.013369f
C767 VTAIL.n223 B 0.023497f
C768 VTAIL.n224 B 0.012626f
C769 VTAIL.n225 B 0.029844f
C770 VTAIL.n226 B 0.013369f
C771 VTAIL.n227 B 0.023497f
C772 VTAIL.n228 B 0.012998f
C773 VTAIL.n229 B 0.029844f
C774 VTAIL.n230 B 0.012626f
C775 VTAIL.n231 B 0.013369f
C776 VTAIL.n232 B 0.023497f
C777 VTAIL.n233 B 0.012626f
C778 VTAIL.n234 B 0.029844f
C779 VTAIL.n235 B 0.013369f
C780 VTAIL.n236 B 0.023497f
C781 VTAIL.n237 B 0.012626f
C782 VTAIL.n238 B 0.029844f
C783 VTAIL.n239 B 0.013369f
C784 VTAIL.n240 B 0.023497f
C785 VTAIL.n241 B 0.012626f
C786 VTAIL.n242 B 0.029844f
C787 VTAIL.n243 B 0.013369f
C788 VTAIL.n244 B 0.023497f
C789 VTAIL.n245 B 0.012626f
C790 VTAIL.n246 B 0.029844f
C791 VTAIL.n247 B 0.013369f
C792 VTAIL.n248 B 0.023497f
C793 VTAIL.n249 B 0.012626f
C794 VTAIL.n250 B 0.022383f
C795 VTAIL.n251 B 0.01763f
C796 VTAIL.t9 B 0.04948f
C797 VTAIL.n252 B 0.17299f
C798 VTAIL.n253 B 1.88952f
C799 VTAIL.n254 B 0.012626f
C800 VTAIL.n255 B 0.013369f
C801 VTAIL.n256 B 0.029844f
C802 VTAIL.n257 B 0.029844f
C803 VTAIL.n258 B 0.013369f
C804 VTAIL.n259 B 0.012626f
C805 VTAIL.n260 B 0.023497f
C806 VTAIL.n261 B 0.023497f
C807 VTAIL.n262 B 0.012626f
C808 VTAIL.n263 B 0.013369f
C809 VTAIL.n264 B 0.029844f
C810 VTAIL.n265 B 0.029844f
C811 VTAIL.n266 B 0.013369f
C812 VTAIL.n267 B 0.012626f
C813 VTAIL.n268 B 0.023497f
C814 VTAIL.n269 B 0.023497f
C815 VTAIL.n270 B 0.012626f
C816 VTAIL.n271 B 0.013369f
C817 VTAIL.n272 B 0.029844f
C818 VTAIL.n273 B 0.029844f
C819 VTAIL.n274 B 0.013369f
C820 VTAIL.n275 B 0.012626f
C821 VTAIL.n276 B 0.023497f
C822 VTAIL.n277 B 0.023497f
C823 VTAIL.n278 B 0.012626f
C824 VTAIL.n279 B 0.013369f
C825 VTAIL.n280 B 0.029844f
C826 VTAIL.n281 B 0.029844f
C827 VTAIL.n282 B 0.013369f
C828 VTAIL.n283 B 0.012626f
C829 VTAIL.n284 B 0.023497f
C830 VTAIL.n285 B 0.023497f
C831 VTAIL.n286 B 0.012626f
C832 VTAIL.n287 B 0.013369f
C833 VTAIL.n288 B 0.029844f
C834 VTAIL.n289 B 0.029844f
C835 VTAIL.n290 B 0.013369f
C836 VTAIL.n291 B 0.012626f
C837 VTAIL.n292 B 0.023497f
C838 VTAIL.n293 B 0.023497f
C839 VTAIL.n294 B 0.012626f
C840 VTAIL.n295 B 0.013369f
C841 VTAIL.n296 B 0.029844f
C842 VTAIL.n297 B 0.029844f
C843 VTAIL.n298 B 0.029844f
C844 VTAIL.n299 B 0.012998f
C845 VTAIL.n300 B 0.012626f
C846 VTAIL.n301 B 0.023497f
C847 VTAIL.n302 B 0.023497f
C848 VTAIL.n303 B 0.012626f
C849 VTAIL.n304 B 0.013369f
C850 VTAIL.n305 B 0.029844f
C851 VTAIL.n306 B 0.029844f
C852 VTAIL.n307 B 0.013369f
C853 VTAIL.n308 B 0.012626f
C854 VTAIL.n309 B 0.023497f
C855 VTAIL.n310 B 0.023497f
C856 VTAIL.n311 B 0.012626f
C857 VTAIL.n312 B 0.013369f
C858 VTAIL.n313 B 0.029844f
C859 VTAIL.n314 B 0.067692f
C860 VTAIL.n315 B 0.013369f
C861 VTAIL.n316 B 0.012626f
C862 VTAIL.n317 B 0.057844f
C863 VTAIL.n318 B 0.038299f
C864 VTAIL.n319 B 1.77915f
C865 VTAIL.n320 B 0.034771f
C866 VTAIL.n321 B 0.023497f
C867 VTAIL.n322 B 0.012626f
C868 VTAIL.n323 B 0.029844f
C869 VTAIL.n324 B 0.013369f
C870 VTAIL.n325 B 0.023497f
C871 VTAIL.n326 B 0.012626f
C872 VTAIL.n327 B 0.029844f
C873 VTAIL.n328 B 0.013369f
C874 VTAIL.n329 B 0.023497f
C875 VTAIL.n330 B 0.012998f
C876 VTAIL.n331 B 0.029844f
C877 VTAIL.n332 B 0.013369f
C878 VTAIL.n333 B 0.023497f
C879 VTAIL.n334 B 0.012626f
C880 VTAIL.n335 B 0.029844f
C881 VTAIL.n336 B 0.013369f
C882 VTAIL.n337 B 0.023497f
C883 VTAIL.n338 B 0.012626f
C884 VTAIL.n339 B 0.029844f
C885 VTAIL.n340 B 0.013369f
C886 VTAIL.n341 B 0.023497f
C887 VTAIL.n342 B 0.012626f
C888 VTAIL.n343 B 0.029844f
C889 VTAIL.n344 B 0.013369f
C890 VTAIL.n345 B 0.023497f
C891 VTAIL.n346 B 0.012626f
C892 VTAIL.n347 B 0.029844f
C893 VTAIL.n348 B 0.013369f
C894 VTAIL.n349 B 0.023497f
C895 VTAIL.n350 B 0.012626f
C896 VTAIL.n351 B 0.022383f
C897 VTAIL.n352 B 0.01763f
C898 VTAIL.t17 B 0.04948f
C899 VTAIL.n353 B 0.17299f
C900 VTAIL.n354 B 1.88952f
C901 VTAIL.n355 B 0.012626f
C902 VTAIL.n356 B 0.013369f
C903 VTAIL.n357 B 0.029844f
C904 VTAIL.n358 B 0.029844f
C905 VTAIL.n359 B 0.013369f
C906 VTAIL.n360 B 0.012626f
C907 VTAIL.n361 B 0.023497f
C908 VTAIL.n362 B 0.023497f
C909 VTAIL.n363 B 0.012626f
C910 VTAIL.n364 B 0.013369f
C911 VTAIL.n365 B 0.029844f
C912 VTAIL.n366 B 0.029844f
C913 VTAIL.n367 B 0.013369f
C914 VTAIL.n368 B 0.012626f
C915 VTAIL.n369 B 0.023497f
C916 VTAIL.n370 B 0.023497f
C917 VTAIL.n371 B 0.012626f
C918 VTAIL.n372 B 0.013369f
C919 VTAIL.n373 B 0.029844f
C920 VTAIL.n374 B 0.029844f
C921 VTAIL.n375 B 0.013369f
C922 VTAIL.n376 B 0.012626f
C923 VTAIL.n377 B 0.023497f
C924 VTAIL.n378 B 0.023497f
C925 VTAIL.n379 B 0.012626f
C926 VTAIL.n380 B 0.013369f
C927 VTAIL.n381 B 0.029844f
C928 VTAIL.n382 B 0.029844f
C929 VTAIL.n383 B 0.013369f
C930 VTAIL.n384 B 0.012626f
C931 VTAIL.n385 B 0.023497f
C932 VTAIL.n386 B 0.023497f
C933 VTAIL.n387 B 0.012626f
C934 VTAIL.n388 B 0.013369f
C935 VTAIL.n389 B 0.029844f
C936 VTAIL.n390 B 0.029844f
C937 VTAIL.n391 B 0.013369f
C938 VTAIL.n392 B 0.012626f
C939 VTAIL.n393 B 0.023497f
C940 VTAIL.n394 B 0.023497f
C941 VTAIL.n395 B 0.012626f
C942 VTAIL.n396 B 0.012626f
C943 VTAIL.n397 B 0.013369f
C944 VTAIL.n398 B 0.029844f
C945 VTAIL.n399 B 0.029844f
C946 VTAIL.n400 B 0.029844f
C947 VTAIL.n401 B 0.012998f
C948 VTAIL.n402 B 0.012626f
C949 VTAIL.n403 B 0.023497f
C950 VTAIL.n404 B 0.023497f
C951 VTAIL.n405 B 0.012626f
C952 VTAIL.n406 B 0.013369f
C953 VTAIL.n407 B 0.029844f
C954 VTAIL.n408 B 0.029844f
C955 VTAIL.n409 B 0.013369f
C956 VTAIL.n410 B 0.012626f
C957 VTAIL.n411 B 0.023497f
C958 VTAIL.n412 B 0.023497f
C959 VTAIL.n413 B 0.012626f
C960 VTAIL.n414 B 0.013369f
C961 VTAIL.n415 B 0.029844f
C962 VTAIL.n416 B 0.067692f
C963 VTAIL.n417 B 0.013369f
C964 VTAIL.n418 B 0.012626f
C965 VTAIL.n419 B 0.057844f
C966 VTAIL.n420 B 0.038299f
C967 VTAIL.n421 B 1.77915f
C968 VTAIL.t12 B 0.340728f
C969 VTAIL.t11 B 0.340728f
C970 VTAIL.n422 B 3.04018f
C971 VTAIL.n423 B 0.375469f
C972 VN.n0 B 0.029096f
C973 VN.t0 B 2.21831f
C974 VN.n1 B 0.043286f
C975 VN.n2 B 0.029096f
C976 VN.t1 B 2.21831f
C977 VN.n3 B 0.054489f
C978 VN.n4 B 0.029096f
C979 VN.t2 B 2.21831f
C980 VN.n5 B 0.050116f
C981 VN.t5 B 2.30899f
C982 VN.t4 B 2.21831f
C983 VN.n6 B 0.838958f
C984 VN.n7 B 0.850025f
C985 VN.n8 B 0.183802f
C986 VN.n9 B 0.029096f
C987 VN.n10 B 0.026004f
C988 VN.n11 B 0.054489f
C989 VN.n12 B 0.807346f
C990 VN.n13 B 0.029096f
C991 VN.n14 B 0.029096f
C992 VN.n15 B 0.029096f
C993 VN.n16 B 0.026004f
C994 VN.n17 B 0.050116f
C995 VN.n18 B 0.779891f
C996 VN.n19 B 0.036022f
C997 VN.n20 B 0.029096f
C998 VN.n21 B 0.029096f
C999 VN.n22 B 0.029096f
C1000 VN.n23 B 0.041664f
C1001 VN.n24 B 0.037093f
C1002 VN.n25 B 0.838593f
C1003 VN.n26 B 0.028247f
C1004 VN.n27 B 0.029096f
C1005 VN.t6 B 2.21831f
C1006 VN.n28 B 0.043286f
C1007 VN.n29 B 0.029096f
C1008 VN.t3 B 2.21831f
C1009 VN.n30 B 0.054489f
C1010 VN.n31 B 0.029096f
C1011 VN.t8 B 2.21831f
C1012 VN.n32 B 0.050116f
C1013 VN.t7 B 2.30899f
C1014 VN.t9 B 2.21831f
C1015 VN.n33 B 0.838958f
C1016 VN.n34 B 0.850025f
C1017 VN.n35 B 0.183802f
C1018 VN.n36 B 0.029096f
C1019 VN.n37 B 0.026004f
C1020 VN.n38 B 0.054489f
C1021 VN.n39 B 0.807346f
C1022 VN.n40 B 0.029096f
C1023 VN.n41 B 0.029096f
C1024 VN.n42 B 0.029096f
C1025 VN.n43 B 0.026004f
C1026 VN.n44 B 0.050116f
C1027 VN.n45 B 0.779891f
C1028 VN.n46 B 0.036022f
C1029 VN.n47 B 0.029096f
C1030 VN.n48 B 0.029096f
C1031 VN.n49 B 0.029096f
C1032 VN.n50 B 0.041664f
C1033 VN.n51 B 0.037093f
C1034 VN.n52 B 0.838593f
C1035 VN.n53 B 1.69725f
.ends

