* NGSPICE file created from diff_pair_sample_1352.ext - technology: sky130A

.subckt diff_pair_sample_1352 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.77
X1 VTAIL.t14 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X2 VDD1.t5 VP.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.77
X3 VDD2.t7 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X4 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.77
X6 VDD1.t7 VP.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X7 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.77
X8 VDD1.t6 VP.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X9 VDD1.t2 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.77
X10 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.77
X11 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.77
X12 VTAIL.t9 VP.t6 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.77
X13 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.77
X14 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X15 VTAIL.t8 VP.t7 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.77
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.77
X18 VTAIL.t6 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.77
X19 VTAIL.t2 VN.t7 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.49335 pd=3.32 as=0.49335 ps=3.32 w=2.99 l=1.77
R0 VP.n31 VP.n30 178.428
R1 VP.n54 VP.n53 178.428
R2 VP.n29 VP.n28 178.428
R3 VP.n14 VP.n11 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n10 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n20 VP.n9 161.3
R8 VP.n23 VP.n22 161.3
R9 VP.n24 VP.n8 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n27 VP.n7 161.3
R12 VP.n52 VP.n0 161.3
R13 VP.n51 VP.n50 161.3
R14 VP.n49 VP.n1 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n45 VP.n2 161.3
R17 VP.n44 VP.n43 161.3
R18 VP.n42 VP.n3 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n4 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n5 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n6 161.3
R25 VP.n12 VP.t0 72.6378
R26 VP.n13 VP.n12 65.2126
R27 VP.n33 VP.n5 50.2061
R28 VP.n51 VP.n1 50.2061
R29 VP.n26 VP.n8 50.2061
R30 VP.n31 VP.t6 40.7118
R31 VP.n38 VP.t3 40.7118
R32 VP.n46 VP.t1 40.7118
R33 VP.n53 VP.t5 40.7118
R34 VP.n28 VP.t2 40.7118
R35 VP.n21 VP.t7 40.7118
R36 VP.n13 VP.t4 40.7118
R37 VP.n40 VP.n3 40.4934
R38 VP.n44 VP.n3 40.4934
R39 VP.n19 VP.n10 40.4934
R40 VP.n15 VP.n10 40.4934
R41 VP.n30 VP.n29 40.1369
R42 VP.n37 VP.n5 30.7807
R43 VP.n47 VP.n1 30.7807
R44 VP.n22 VP.n8 30.7807
R45 VP.n33 VP.n32 24.4675
R46 VP.n40 VP.n39 24.4675
R47 VP.n45 VP.n44 24.4675
R48 VP.n52 VP.n51 24.4675
R49 VP.n27 VP.n26 24.4675
R50 VP.n20 VP.n19 24.4675
R51 VP.n15 VP.n14 24.4675
R52 VP.n38 VP.n37 22.0208
R53 VP.n47 VP.n46 22.0208
R54 VP.n22 VP.n21 22.0208
R55 VP.n12 VP.n11 18.1539
R56 VP.n32 VP.n31 7.3406
R57 VP.n53 VP.n52 7.3406
R58 VP.n28 VP.n27 7.3406
R59 VP.n39 VP.n38 2.4472
R60 VP.n46 VP.n45 2.4472
R61 VP.n21 VP.n20 2.4472
R62 VP.n14 VP.n13 2.4472
R63 VP.n16 VP.n11 0.189894
R64 VP.n17 VP.n16 0.189894
R65 VP.n18 VP.n17 0.189894
R66 VP.n18 VP.n9 0.189894
R67 VP.n23 VP.n9 0.189894
R68 VP.n24 VP.n23 0.189894
R69 VP.n25 VP.n24 0.189894
R70 VP.n25 VP.n7 0.189894
R71 VP.n29 VP.n7 0.189894
R72 VP.n30 VP.n6 0.189894
R73 VP.n34 VP.n6 0.189894
R74 VP.n35 VP.n34 0.189894
R75 VP.n36 VP.n35 0.189894
R76 VP.n36 VP.n4 0.189894
R77 VP.n41 VP.n4 0.189894
R78 VP.n42 VP.n41 0.189894
R79 VP.n43 VP.n42 0.189894
R80 VP.n43 VP.n2 0.189894
R81 VP.n48 VP.n2 0.189894
R82 VP.n49 VP.n48 0.189894
R83 VP.n50 VP.n49 0.189894
R84 VP.n50 VP.n0 0.189894
R85 VP.n54 VP.n0 0.189894
R86 VP VP.n54 0.0516364
R87 VDD1 VDD1.n0 86.2526
R88 VDD1.n3 VDD1.n2 86.1388
R89 VDD1.n3 VDD1.n1 86.1388
R90 VDD1.n5 VDD1.n4 85.2891
R91 VDD1.n5 VDD1.n3 35.0224
R92 VDD1.n4 VDD1.t3 6.62257
R93 VDD1.n4 VDD1.t5 6.62257
R94 VDD1.n0 VDD1.t1 6.62257
R95 VDD1.n0 VDD1.t6 6.62257
R96 VDD1.n2 VDD1.t4 6.62257
R97 VDD1.n2 VDD1.t2 6.62257
R98 VDD1.n1 VDD1.t0 6.62257
R99 VDD1.n1 VDD1.t7 6.62257
R100 VDD1 VDD1.n5 0.847483
R101 VTAIL.n11 VTAIL.t15 75.2325
R102 VTAIL.n10 VTAIL.t1 75.2325
R103 VTAIL.n7 VTAIL.t6 75.2325
R104 VTAIL.n15 VTAIL.t3 75.2322
R105 VTAIL.n2 VTAIL.t0 75.2322
R106 VTAIL.n3 VTAIL.t10 75.2322
R107 VTAIL.n6 VTAIL.t9 75.2322
R108 VTAIL.n14 VTAIL.t13 75.2322
R109 VTAIL.n13 VTAIL.n12 68.6104
R110 VTAIL.n9 VTAIL.n8 68.6104
R111 VTAIL.n1 VTAIL.n0 68.6102
R112 VTAIL.n5 VTAIL.n4 68.6102
R113 VTAIL.n15 VTAIL.n14 16.7548
R114 VTAIL.n7 VTAIL.n6 16.7548
R115 VTAIL.n0 VTAIL.t4 6.62257
R116 VTAIL.n0 VTAIL.t7 6.62257
R117 VTAIL.n4 VTAIL.t12 6.62257
R118 VTAIL.n4 VTAIL.t14 6.62257
R119 VTAIL.n12 VTAIL.t11 6.62257
R120 VTAIL.n12 VTAIL.t8 6.62257
R121 VTAIL.n8 VTAIL.t5 6.62257
R122 VTAIL.n8 VTAIL.t2 6.62257
R123 VTAIL.n9 VTAIL.n7 1.81084
R124 VTAIL.n10 VTAIL.n9 1.81084
R125 VTAIL.n13 VTAIL.n11 1.81084
R126 VTAIL.n14 VTAIL.n13 1.81084
R127 VTAIL.n6 VTAIL.n5 1.81084
R128 VTAIL.n5 VTAIL.n3 1.81084
R129 VTAIL.n2 VTAIL.n1 1.81084
R130 VTAIL VTAIL.n15 1.75266
R131 VTAIL.n11 VTAIL.n10 0.470328
R132 VTAIL.n3 VTAIL.n2 0.470328
R133 VTAIL VTAIL.n1 0.0586897
R134 B.n522 B.n521 585
R135 B.n173 B.n93 585
R136 B.n172 B.n171 585
R137 B.n170 B.n169 585
R138 B.n168 B.n167 585
R139 B.n166 B.n165 585
R140 B.n164 B.n163 585
R141 B.n162 B.n161 585
R142 B.n160 B.n159 585
R143 B.n158 B.n157 585
R144 B.n156 B.n155 585
R145 B.n154 B.n153 585
R146 B.n152 B.n151 585
R147 B.n150 B.n149 585
R148 B.n148 B.n147 585
R149 B.n145 B.n144 585
R150 B.n143 B.n142 585
R151 B.n141 B.n140 585
R152 B.n139 B.n138 585
R153 B.n137 B.n136 585
R154 B.n135 B.n134 585
R155 B.n133 B.n132 585
R156 B.n131 B.n130 585
R157 B.n129 B.n128 585
R158 B.n127 B.n126 585
R159 B.n124 B.n123 585
R160 B.n122 B.n121 585
R161 B.n120 B.n119 585
R162 B.n118 B.n117 585
R163 B.n116 B.n115 585
R164 B.n114 B.n113 585
R165 B.n112 B.n111 585
R166 B.n110 B.n109 585
R167 B.n108 B.n107 585
R168 B.n106 B.n105 585
R169 B.n104 B.n103 585
R170 B.n102 B.n101 585
R171 B.n100 B.n99 585
R172 B.n74 B.n73 585
R173 B.n527 B.n526 585
R174 B.n520 B.n94 585
R175 B.n94 B.n71 585
R176 B.n519 B.n70 585
R177 B.n531 B.n70 585
R178 B.n518 B.n69 585
R179 B.n532 B.n69 585
R180 B.n517 B.n68 585
R181 B.n533 B.n68 585
R182 B.n516 B.n515 585
R183 B.n515 B.n64 585
R184 B.n514 B.n63 585
R185 B.n539 B.n63 585
R186 B.n513 B.n62 585
R187 B.n540 B.n62 585
R188 B.n512 B.n61 585
R189 B.n541 B.n61 585
R190 B.n511 B.n510 585
R191 B.n510 B.n57 585
R192 B.n509 B.n56 585
R193 B.n547 B.n56 585
R194 B.n508 B.n55 585
R195 B.n548 B.n55 585
R196 B.n507 B.n54 585
R197 B.n549 B.n54 585
R198 B.n506 B.n505 585
R199 B.n505 B.n50 585
R200 B.n504 B.n49 585
R201 B.n555 B.n49 585
R202 B.n503 B.n48 585
R203 B.n556 B.n48 585
R204 B.n502 B.n47 585
R205 B.n557 B.n47 585
R206 B.n501 B.n500 585
R207 B.n500 B.n43 585
R208 B.n499 B.n42 585
R209 B.n563 B.n42 585
R210 B.n498 B.n41 585
R211 B.n564 B.n41 585
R212 B.n497 B.n40 585
R213 B.n565 B.n40 585
R214 B.n496 B.n495 585
R215 B.n495 B.n36 585
R216 B.n494 B.n35 585
R217 B.n571 B.n35 585
R218 B.n493 B.n34 585
R219 B.n572 B.n34 585
R220 B.n492 B.n33 585
R221 B.n573 B.n33 585
R222 B.n491 B.n490 585
R223 B.n490 B.n29 585
R224 B.n489 B.n28 585
R225 B.n579 B.n28 585
R226 B.n488 B.n27 585
R227 B.n580 B.n27 585
R228 B.n487 B.n26 585
R229 B.n581 B.n26 585
R230 B.n486 B.n485 585
R231 B.n485 B.n25 585
R232 B.n484 B.n21 585
R233 B.n587 B.n21 585
R234 B.n483 B.n20 585
R235 B.n588 B.n20 585
R236 B.n482 B.n19 585
R237 B.n589 B.n19 585
R238 B.n481 B.n480 585
R239 B.n480 B.n15 585
R240 B.n479 B.n14 585
R241 B.n595 B.n14 585
R242 B.n478 B.n13 585
R243 B.n596 B.n13 585
R244 B.n477 B.n12 585
R245 B.n597 B.n12 585
R246 B.n476 B.n475 585
R247 B.n475 B.n8 585
R248 B.n474 B.n7 585
R249 B.n603 B.n7 585
R250 B.n473 B.n6 585
R251 B.n604 B.n6 585
R252 B.n472 B.n5 585
R253 B.n605 B.n5 585
R254 B.n471 B.n470 585
R255 B.n470 B.n4 585
R256 B.n469 B.n174 585
R257 B.n469 B.n468 585
R258 B.n459 B.n175 585
R259 B.n176 B.n175 585
R260 B.n461 B.n460 585
R261 B.n462 B.n461 585
R262 B.n458 B.n180 585
R263 B.n184 B.n180 585
R264 B.n457 B.n456 585
R265 B.n456 B.n455 585
R266 B.n182 B.n181 585
R267 B.n183 B.n182 585
R268 B.n448 B.n447 585
R269 B.n449 B.n448 585
R270 B.n446 B.n189 585
R271 B.n189 B.n188 585
R272 B.n445 B.n444 585
R273 B.n444 B.n443 585
R274 B.n191 B.n190 585
R275 B.n436 B.n191 585
R276 B.n435 B.n434 585
R277 B.n437 B.n435 585
R278 B.n433 B.n196 585
R279 B.n196 B.n195 585
R280 B.n432 B.n431 585
R281 B.n431 B.n430 585
R282 B.n198 B.n197 585
R283 B.n199 B.n198 585
R284 B.n423 B.n422 585
R285 B.n424 B.n423 585
R286 B.n421 B.n204 585
R287 B.n204 B.n203 585
R288 B.n420 B.n419 585
R289 B.n419 B.n418 585
R290 B.n206 B.n205 585
R291 B.n207 B.n206 585
R292 B.n411 B.n410 585
R293 B.n412 B.n411 585
R294 B.n409 B.n212 585
R295 B.n212 B.n211 585
R296 B.n408 B.n407 585
R297 B.n407 B.n406 585
R298 B.n214 B.n213 585
R299 B.n215 B.n214 585
R300 B.n399 B.n398 585
R301 B.n400 B.n399 585
R302 B.n397 B.n220 585
R303 B.n220 B.n219 585
R304 B.n396 B.n395 585
R305 B.n395 B.n394 585
R306 B.n222 B.n221 585
R307 B.n223 B.n222 585
R308 B.n387 B.n386 585
R309 B.n388 B.n387 585
R310 B.n385 B.n228 585
R311 B.n228 B.n227 585
R312 B.n384 B.n383 585
R313 B.n383 B.n382 585
R314 B.n230 B.n229 585
R315 B.n231 B.n230 585
R316 B.n375 B.n374 585
R317 B.n376 B.n375 585
R318 B.n373 B.n235 585
R319 B.n239 B.n235 585
R320 B.n372 B.n371 585
R321 B.n371 B.n370 585
R322 B.n237 B.n236 585
R323 B.n238 B.n237 585
R324 B.n363 B.n362 585
R325 B.n364 B.n363 585
R326 B.n361 B.n244 585
R327 B.n244 B.n243 585
R328 B.n360 B.n359 585
R329 B.n359 B.n358 585
R330 B.n246 B.n245 585
R331 B.n247 B.n246 585
R332 B.n354 B.n353 585
R333 B.n250 B.n249 585
R334 B.n350 B.n349 585
R335 B.n351 B.n350 585
R336 B.n348 B.n270 585
R337 B.n347 B.n346 585
R338 B.n345 B.n344 585
R339 B.n343 B.n342 585
R340 B.n341 B.n340 585
R341 B.n339 B.n338 585
R342 B.n337 B.n336 585
R343 B.n335 B.n334 585
R344 B.n333 B.n332 585
R345 B.n331 B.n330 585
R346 B.n329 B.n328 585
R347 B.n327 B.n326 585
R348 B.n325 B.n324 585
R349 B.n323 B.n322 585
R350 B.n321 B.n320 585
R351 B.n319 B.n318 585
R352 B.n317 B.n316 585
R353 B.n315 B.n314 585
R354 B.n313 B.n312 585
R355 B.n311 B.n310 585
R356 B.n309 B.n308 585
R357 B.n307 B.n306 585
R358 B.n305 B.n304 585
R359 B.n303 B.n302 585
R360 B.n301 B.n300 585
R361 B.n299 B.n298 585
R362 B.n297 B.n296 585
R363 B.n295 B.n294 585
R364 B.n293 B.n292 585
R365 B.n291 B.n290 585
R366 B.n289 B.n288 585
R367 B.n287 B.n286 585
R368 B.n285 B.n284 585
R369 B.n283 B.n282 585
R370 B.n281 B.n280 585
R371 B.n279 B.n278 585
R372 B.n277 B.n269 585
R373 B.n351 B.n269 585
R374 B.n355 B.n248 585
R375 B.n248 B.n247 585
R376 B.n357 B.n356 585
R377 B.n358 B.n357 585
R378 B.n242 B.n241 585
R379 B.n243 B.n242 585
R380 B.n366 B.n365 585
R381 B.n365 B.n364 585
R382 B.n367 B.n240 585
R383 B.n240 B.n238 585
R384 B.n369 B.n368 585
R385 B.n370 B.n369 585
R386 B.n234 B.n233 585
R387 B.n239 B.n234 585
R388 B.n378 B.n377 585
R389 B.n377 B.n376 585
R390 B.n379 B.n232 585
R391 B.n232 B.n231 585
R392 B.n381 B.n380 585
R393 B.n382 B.n381 585
R394 B.n226 B.n225 585
R395 B.n227 B.n226 585
R396 B.n390 B.n389 585
R397 B.n389 B.n388 585
R398 B.n391 B.n224 585
R399 B.n224 B.n223 585
R400 B.n393 B.n392 585
R401 B.n394 B.n393 585
R402 B.n218 B.n217 585
R403 B.n219 B.n218 585
R404 B.n402 B.n401 585
R405 B.n401 B.n400 585
R406 B.n403 B.n216 585
R407 B.n216 B.n215 585
R408 B.n405 B.n404 585
R409 B.n406 B.n405 585
R410 B.n210 B.n209 585
R411 B.n211 B.n210 585
R412 B.n414 B.n413 585
R413 B.n413 B.n412 585
R414 B.n415 B.n208 585
R415 B.n208 B.n207 585
R416 B.n417 B.n416 585
R417 B.n418 B.n417 585
R418 B.n202 B.n201 585
R419 B.n203 B.n202 585
R420 B.n426 B.n425 585
R421 B.n425 B.n424 585
R422 B.n427 B.n200 585
R423 B.n200 B.n199 585
R424 B.n429 B.n428 585
R425 B.n430 B.n429 585
R426 B.n194 B.n193 585
R427 B.n195 B.n194 585
R428 B.n439 B.n438 585
R429 B.n438 B.n437 585
R430 B.n440 B.n192 585
R431 B.n436 B.n192 585
R432 B.n442 B.n441 585
R433 B.n443 B.n442 585
R434 B.n187 B.n186 585
R435 B.n188 B.n187 585
R436 B.n451 B.n450 585
R437 B.n450 B.n449 585
R438 B.n452 B.n185 585
R439 B.n185 B.n183 585
R440 B.n454 B.n453 585
R441 B.n455 B.n454 585
R442 B.n179 B.n178 585
R443 B.n184 B.n179 585
R444 B.n464 B.n463 585
R445 B.n463 B.n462 585
R446 B.n465 B.n177 585
R447 B.n177 B.n176 585
R448 B.n467 B.n466 585
R449 B.n468 B.n467 585
R450 B.n2 B.n0 585
R451 B.n4 B.n2 585
R452 B.n3 B.n1 585
R453 B.n604 B.n3 585
R454 B.n602 B.n601 585
R455 B.n603 B.n602 585
R456 B.n600 B.n9 585
R457 B.n9 B.n8 585
R458 B.n599 B.n598 585
R459 B.n598 B.n597 585
R460 B.n11 B.n10 585
R461 B.n596 B.n11 585
R462 B.n594 B.n593 585
R463 B.n595 B.n594 585
R464 B.n592 B.n16 585
R465 B.n16 B.n15 585
R466 B.n591 B.n590 585
R467 B.n590 B.n589 585
R468 B.n18 B.n17 585
R469 B.n588 B.n18 585
R470 B.n586 B.n585 585
R471 B.n587 B.n586 585
R472 B.n584 B.n22 585
R473 B.n25 B.n22 585
R474 B.n583 B.n582 585
R475 B.n582 B.n581 585
R476 B.n24 B.n23 585
R477 B.n580 B.n24 585
R478 B.n578 B.n577 585
R479 B.n579 B.n578 585
R480 B.n576 B.n30 585
R481 B.n30 B.n29 585
R482 B.n575 B.n574 585
R483 B.n574 B.n573 585
R484 B.n32 B.n31 585
R485 B.n572 B.n32 585
R486 B.n570 B.n569 585
R487 B.n571 B.n570 585
R488 B.n568 B.n37 585
R489 B.n37 B.n36 585
R490 B.n567 B.n566 585
R491 B.n566 B.n565 585
R492 B.n39 B.n38 585
R493 B.n564 B.n39 585
R494 B.n562 B.n561 585
R495 B.n563 B.n562 585
R496 B.n560 B.n44 585
R497 B.n44 B.n43 585
R498 B.n559 B.n558 585
R499 B.n558 B.n557 585
R500 B.n46 B.n45 585
R501 B.n556 B.n46 585
R502 B.n554 B.n553 585
R503 B.n555 B.n554 585
R504 B.n552 B.n51 585
R505 B.n51 B.n50 585
R506 B.n551 B.n550 585
R507 B.n550 B.n549 585
R508 B.n53 B.n52 585
R509 B.n548 B.n53 585
R510 B.n546 B.n545 585
R511 B.n547 B.n546 585
R512 B.n544 B.n58 585
R513 B.n58 B.n57 585
R514 B.n543 B.n542 585
R515 B.n542 B.n541 585
R516 B.n60 B.n59 585
R517 B.n540 B.n60 585
R518 B.n538 B.n537 585
R519 B.n539 B.n538 585
R520 B.n536 B.n65 585
R521 B.n65 B.n64 585
R522 B.n535 B.n534 585
R523 B.n534 B.n533 585
R524 B.n67 B.n66 585
R525 B.n532 B.n67 585
R526 B.n530 B.n529 585
R527 B.n531 B.n530 585
R528 B.n528 B.n72 585
R529 B.n72 B.n71 585
R530 B.n607 B.n606 585
R531 B.n606 B.n605 585
R532 B.n353 B.n248 482.89
R533 B.n526 B.n72 482.89
R534 B.n269 B.n246 482.89
R535 B.n522 B.n94 482.89
R536 B.n524 B.n523 256.663
R537 B.n524 B.n92 256.663
R538 B.n524 B.n91 256.663
R539 B.n524 B.n90 256.663
R540 B.n524 B.n89 256.663
R541 B.n524 B.n88 256.663
R542 B.n524 B.n87 256.663
R543 B.n524 B.n86 256.663
R544 B.n524 B.n85 256.663
R545 B.n524 B.n84 256.663
R546 B.n524 B.n83 256.663
R547 B.n524 B.n82 256.663
R548 B.n524 B.n81 256.663
R549 B.n524 B.n80 256.663
R550 B.n524 B.n79 256.663
R551 B.n524 B.n78 256.663
R552 B.n524 B.n77 256.663
R553 B.n524 B.n76 256.663
R554 B.n524 B.n75 256.663
R555 B.n525 B.n524 256.663
R556 B.n352 B.n351 256.663
R557 B.n351 B.n251 256.663
R558 B.n351 B.n252 256.663
R559 B.n351 B.n253 256.663
R560 B.n351 B.n254 256.663
R561 B.n351 B.n255 256.663
R562 B.n351 B.n256 256.663
R563 B.n351 B.n257 256.663
R564 B.n351 B.n258 256.663
R565 B.n351 B.n259 256.663
R566 B.n351 B.n260 256.663
R567 B.n351 B.n261 256.663
R568 B.n351 B.n262 256.663
R569 B.n351 B.n263 256.663
R570 B.n351 B.n264 256.663
R571 B.n351 B.n265 256.663
R572 B.n351 B.n266 256.663
R573 B.n351 B.n267 256.663
R574 B.n351 B.n268 256.663
R575 B.n274 B.t8 247.032
R576 B.n271 B.t19 247.032
R577 B.n97 B.t16 247.032
R578 B.n95 B.t12 247.032
R579 B.n351 B.n247 163.702
R580 B.n524 B.n71 163.702
R581 B.n357 B.n248 163.367
R582 B.n357 B.n242 163.367
R583 B.n365 B.n242 163.367
R584 B.n365 B.n240 163.367
R585 B.n369 B.n240 163.367
R586 B.n369 B.n234 163.367
R587 B.n377 B.n234 163.367
R588 B.n377 B.n232 163.367
R589 B.n381 B.n232 163.367
R590 B.n381 B.n226 163.367
R591 B.n389 B.n226 163.367
R592 B.n389 B.n224 163.367
R593 B.n393 B.n224 163.367
R594 B.n393 B.n218 163.367
R595 B.n401 B.n218 163.367
R596 B.n401 B.n216 163.367
R597 B.n405 B.n216 163.367
R598 B.n405 B.n210 163.367
R599 B.n413 B.n210 163.367
R600 B.n413 B.n208 163.367
R601 B.n417 B.n208 163.367
R602 B.n417 B.n202 163.367
R603 B.n425 B.n202 163.367
R604 B.n425 B.n200 163.367
R605 B.n429 B.n200 163.367
R606 B.n429 B.n194 163.367
R607 B.n438 B.n194 163.367
R608 B.n438 B.n192 163.367
R609 B.n442 B.n192 163.367
R610 B.n442 B.n187 163.367
R611 B.n450 B.n187 163.367
R612 B.n450 B.n185 163.367
R613 B.n454 B.n185 163.367
R614 B.n454 B.n179 163.367
R615 B.n463 B.n179 163.367
R616 B.n463 B.n177 163.367
R617 B.n467 B.n177 163.367
R618 B.n467 B.n2 163.367
R619 B.n606 B.n2 163.367
R620 B.n606 B.n3 163.367
R621 B.n602 B.n3 163.367
R622 B.n602 B.n9 163.367
R623 B.n598 B.n9 163.367
R624 B.n598 B.n11 163.367
R625 B.n594 B.n11 163.367
R626 B.n594 B.n16 163.367
R627 B.n590 B.n16 163.367
R628 B.n590 B.n18 163.367
R629 B.n586 B.n18 163.367
R630 B.n586 B.n22 163.367
R631 B.n582 B.n22 163.367
R632 B.n582 B.n24 163.367
R633 B.n578 B.n24 163.367
R634 B.n578 B.n30 163.367
R635 B.n574 B.n30 163.367
R636 B.n574 B.n32 163.367
R637 B.n570 B.n32 163.367
R638 B.n570 B.n37 163.367
R639 B.n566 B.n37 163.367
R640 B.n566 B.n39 163.367
R641 B.n562 B.n39 163.367
R642 B.n562 B.n44 163.367
R643 B.n558 B.n44 163.367
R644 B.n558 B.n46 163.367
R645 B.n554 B.n46 163.367
R646 B.n554 B.n51 163.367
R647 B.n550 B.n51 163.367
R648 B.n550 B.n53 163.367
R649 B.n546 B.n53 163.367
R650 B.n546 B.n58 163.367
R651 B.n542 B.n58 163.367
R652 B.n542 B.n60 163.367
R653 B.n538 B.n60 163.367
R654 B.n538 B.n65 163.367
R655 B.n534 B.n65 163.367
R656 B.n534 B.n67 163.367
R657 B.n530 B.n67 163.367
R658 B.n530 B.n72 163.367
R659 B.n350 B.n250 163.367
R660 B.n350 B.n270 163.367
R661 B.n346 B.n345 163.367
R662 B.n342 B.n341 163.367
R663 B.n338 B.n337 163.367
R664 B.n334 B.n333 163.367
R665 B.n330 B.n329 163.367
R666 B.n326 B.n325 163.367
R667 B.n322 B.n321 163.367
R668 B.n318 B.n317 163.367
R669 B.n314 B.n313 163.367
R670 B.n310 B.n309 163.367
R671 B.n306 B.n305 163.367
R672 B.n302 B.n301 163.367
R673 B.n298 B.n297 163.367
R674 B.n294 B.n293 163.367
R675 B.n290 B.n289 163.367
R676 B.n286 B.n285 163.367
R677 B.n282 B.n281 163.367
R678 B.n278 B.n269 163.367
R679 B.n359 B.n246 163.367
R680 B.n359 B.n244 163.367
R681 B.n363 B.n244 163.367
R682 B.n363 B.n237 163.367
R683 B.n371 B.n237 163.367
R684 B.n371 B.n235 163.367
R685 B.n375 B.n235 163.367
R686 B.n375 B.n230 163.367
R687 B.n383 B.n230 163.367
R688 B.n383 B.n228 163.367
R689 B.n387 B.n228 163.367
R690 B.n387 B.n222 163.367
R691 B.n395 B.n222 163.367
R692 B.n395 B.n220 163.367
R693 B.n399 B.n220 163.367
R694 B.n399 B.n214 163.367
R695 B.n407 B.n214 163.367
R696 B.n407 B.n212 163.367
R697 B.n411 B.n212 163.367
R698 B.n411 B.n206 163.367
R699 B.n419 B.n206 163.367
R700 B.n419 B.n204 163.367
R701 B.n423 B.n204 163.367
R702 B.n423 B.n198 163.367
R703 B.n431 B.n198 163.367
R704 B.n431 B.n196 163.367
R705 B.n435 B.n196 163.367
R706 B.n435 B.n191 163.367
R707 B.n444 B.n191 163.367
R708 B.n444 B.n189 163.367
R709 B.n448 B.n189 163.367
R710 B.n448 B.n182 163.367
R711 B.n456 B.n182 163.367
R712 B.n456 B.n180 163.367
R713 B.n461 B.n180 163.367
R714 B.n461 B.n175 163.367
R715 B.n469 B.n175 163.367
R716 B.n470 B.n469 163.367
R717 B.n470 B.n5 163.367
R718 B.n6 B.n5 163.367
R719 B.n7 B.n6 163.367
R720 B.n475 B.n7 163.367
R721 B.n475 B.n12 163.367
R722 B.n13 B.n12 163.367
R723 B.n14 B.n13 163.367
R724 B.n480 B.n14 163.367
R725 B.n480 B.n19 163.367
R726 B.n20 B.n19 163.367
R727 B.n21 B.n20 163.367
R728 B.n485 B.n21 163.367
R729 B.n485 B.n26 163.367
R730 B.n27 B.n26 163.367
R731 B.n28 B.n27 163.367
R732 B.n490 B.n28 163.367
R733 B.n490 B.n33 163.367
R734 B.n34 B.n33 163.367
R735 B.n35 B.n34 163.367
R736 B.n495 B.n35 163.367
R737 B.n495 B.n40 163.367
R738 B.n41 B.n40 163.367
R739 B.n42 B.n41 163.367
R740 B.n500 B.n42 163.367
R741 B.n500 B.n47 163.367
R742 B.n48 B.n47 163.367
R743 B.n49 B.n48 163.367
R744 B.n505 B.n49 163.367
R745 B.n505 B.n54 163.367
R746 B.n55 B.n54 163.367
R747 B.n56 B.n55 163.367
R748 B.n510 B.n56 163.367
R749 B.n510 B.n61 163.367
R750 B.n62 B.n61 163.367
R751 B.n63 B.n62 163.367
R752 B.n515 B.n63 163.367
R753 B.n515 B.n68 163.367
R754 B.n69 B.n68 163.367
R755 B.n70 B.n69 163.367
R756 B.n94 B.n70 163.367
R757 B.n99 B.n74 163.367
R758 B.n103 B.n102 163.367
R759 B.n107 B.n106 163.367
R760 B.n111 B.n110 163.367
R761 B.n115 B.n114 163.367
R762 B.n119 B.n118 163.367
R763 B.n123 B.n122 163.367
R764 B.n128 B.n127 163.367
R765 B.n132 B.n131 163.367
R766 B.n136 B.n135 163.367
R767 B.n140 B.n139 163.367
R768 B.n144 B.n143 163.367
R769 B.n149 B.n148 163.367
R770 B.n153 B.n152 163.367
R771 B.n157 B.n156 163.367
R772 B.n161 B.n160 163.367
R773 B.n165 B.n164 163.367
R774 B.n169 B.n168 163.367
R775 B.n171 B.n93 163.367
R776 B.n274 B.t11 121.171
R777 B.n95 B.t14 121.171
R778 B.n271 B.t21 121.168
R779 B.n97 B.t17 121.168
R780 B.n358 B.n247 90.5026
R781 B.n358 B.n243 90.5026
R782 B.n364 B.n243 90.5026
R783 B.n364 B.n238 90.5026
R784 B.n370 B.n238 90.5026
R785 B.n370 B.n239 90.5026
R786 B.n376 B.n231 90.5026
R787 B.n382 B.n231 90.5026
R788 B.n382 B.n227 90.5026
R789 B.n388 B.n227 90.5026
R790 B.n388 B.n223 90.5026
R791 B.n394 B.n223 90.5026
R792 B.n394 B.n219 90.5026
R793 B.n400 B.n219 90.5026
R794 B.n406 B.n215 90.5026
R795 B.n406 B.n211 90.5026
R796 B.n412 B.n211 90.5026
R797 B.n412 B.n207 90.5026
R798 B.n418 B.n207 90.5026
R799 B.n424 B.n203 90.5026
R800 B.n424 B.n199 90.5026
R801 B.n430 B.n199 90.5026
R802 B.n430 B.n195 90.5026
R803 B.n437 B.n195 90.5026
R804 B.n437 B.n436 90.5026
R805 B.n443 B.n188 90.5026
R806 B.n449 B.n188 90.5026
R807 B.n449 B.n183 90.5026
R808 B.n455 B.n183 90.5026
R809 B.n455 B.n184 90.5026
R810 B.n462 B.n176 90.5026
R811 B.n468 B.n176 90.5026
R812 B.n468 B.n4 90.5026
R813 B.n605 B.n4 90.5026
R814 B.n605 B.n604 90.5026
R815 B.n604 B.n603 90.5026
R816 B.n603 B.n8 90.5026
R817 B.n597 B.n8 90.5026
R818 B.n596 B.n595 90.5026
R819 B.n595 B.n15 90.5026
R820 B.n589 B.n15 90.5026
R821 B.n589 B.n588 90.5026
R822 B.n588 B.n587 90.5026
R823 B.n581 B.n25 90.5026
R824 B.n581 B.n580 90.5026
R825 B.n580 B.n579 90.5026
R826 B.n579 B.n29 90.5026
R827 B.n573 B.n29 90.5026
R828 B.n573 B.n572 90.5026
R829 B.n571 B.n36 90.5026
R830 B.n565 B.n36 90.5026
R831 B.n565 B.n564 90.5026
R832 B.n564 B.n563 90.5026
R833 B.n563 B.n43 90.5026
R834 B.n557 B.n556 90.5026
R835 B.n556 B.n555 90.5026
R836 B.n555 B.n50 90.5026
R837 B.n549 B.n50 90.5026
R838 B.n549 B.n548 90.5026
R839 B.n548 B.n547 90.5026
R840 B.n547 B.n57 90.5026
R841 B.n541 B.n57 90.5026
R842 B.n540 B.n539 90.5026
R843 B.n539 B.n64 90.5026
R844 B.n533 B.n64 90.5026
R845 B.n533 B.n532 90.5026
R846 B.n532 B.n531 90.5026
R847 B.n531 B.n71 90.5026
R848 B.n418 B.t5 86.5099
R849 B.t7 B.n571 86.5099
R850 B.n275 B.t10 80.4429
R851 B.n96 B.t15 80.4429
R852 B.n272 B.t20 80.4411
R853 B.n98 B.t18 80.4411
R854 B.n443 B.t2 78.5244
R855 B.n587 B.t4 78.5244
R856 B.n353 B.n352 71.676
R857 B.n270 B.n251 71.676
R858 B.n345 B.n252 71.676
R859 B.n341 B.n253 71.676
R860 B.n337 B.n254 71.676
R861 B.n333 B.n255 71.676
R862 B.n329 B.n256 71.676
R863 B.n325 B.n257 71.676
R864 B.n321 B.n258 71.676
R865 B.n317 B.n259 71.676
R866 B.n313 B.n260 71.676
R867 B.n309 B.n261 71.676
R868 B.n305 B.n262 71.676
R869 B.n301 B.n263 71.676
R870 B.n297 B.n264 71.676
R871 B.n293 B.n265 71.676
R872 B.n289 B.n266 71.676
R873 B.n285 B.n267 71.676
R874 B.n281 B.n268 71.676
R875 B.n526 B.n525 71.676
R876 B.n99 B.n75 71.676
R877 B.n103 B.n76 71.676
R878 B.n107 B.n77 71.676
R879 B.n111 B.n78 71.676
R880 B.n115 B.n79 71.676
R881 B.n119 B.n80 71.676
R882 B.n123 B.n81 71.676
R883 B.n128 B.n82 71.676
R884 B.n132 B.n83 71.676
R885 B.n136 B.n84 71.676
R886 B.n140 B.n85 71.676
R887 B.n144 B.n86 71.676
R888 B.n149 B.n87 71.676
R889 B.n153 B.n88 71.676
R890 B.n157 B.n89 71.676
R891 B.n161 B.n90 71.676
R892 B.n165 B.n91 71.676
R893 B.n169 B.n92 71.676
R894 B.n523 B.n93 71.676
R895 B.n523 B.n522 71.676
R896 B.n171 B.n92 71.676
R897 B.n168 B.n91 71.676
R898 B.n164 B.n90 71.676
R899 B.n160 B.n89 71.676
R900 B.n156 B.n88 71.676
R901 B.n152 B.n87 71.676
R902 B.n148 B.n86 71.676
R903 B.n143 B.n85 71.676
R904 B.n139 B.n84 71.676
R905 B.n135 B.n83 71.676
R906 B.n131 B.n82 71.676
R907 B.n127 B.n81 71.676
R908 B.n122 B.n80 71.676
R909 B.n118 B.n79 71.676
R910 B.n114 B.n78 71.676
R911 B.n110 B.n77 71.676
R912 B.n106 B.n76 71.676
R913 B.n102 B.n75 71.676
R914 B.n525 B.n74 71.676
R915 B.n352 B.n250 71.676
R916 B.n346 B.n251 71.676
R917 B.n342 B.n252 71.676
R918 B.n338 B.n253 71.676
R919 B.n334 B.n254 71.676
R920 B.n330 B.n255 71.676
R921 B.n326 B.n256 71.676
R922 B.n322 B.n257 71.676
R923 B.n318 B.n258 71.676
R924 B.n314 B.n259 71.676
R925 B.n310 B.n260 71.676
R926 B.n306 B.n261 71.676
R927 B.n302 B.n262 71.676
R928 B.n298 B.n263 71.676
R929 B.n294 B.n264 71.676
R930 B.n290 B.n265 71.676
R931 B.n286 B.n266 71.676
R932 B.n282 B.n267 71.676
R933 B.n278 B.n268 71.676
R934 B.n400 B.t6 70.5389
R935 B.n557 B.t3 70.5389
R936 B.n462 B.t1 62.5534
R937 B.n597 B.t0 62.5534
R938 B.n276 B.n275 59.5399
R939 B.n273 B.n272 59.5399
R940 B.n125 B.n98 59.5399
R941 B.n146 B.n96 59.5399
R942 B.n376 B.t9 54.568
R943 B.n541 B.t13 54.568
R944 B.n275 B.n274 40.7278
R945 B.n272 B.n271 40.7278
R946 B.n98 B.n97 40.7278
R947 B.n96 B.n95 40.7278
R948 B.n239 B.t9 35.9352
R949 B.t13 B.n540 35.9352
R950 B.n528 B.n527 31.3761
R951 B.n521 B.n520 31.3761
R952 B.n277 B.n245 31.3761
R953 B.n355 B.n354 31.3761
R954 B.n184 B.t1 27.9497
R955 B.t0 B.n596 27.9497
R956 B.t6 B.n215 19.9642
R957 B.t3 B.n43 19.9642
R958 B B.n607 18.0485
R959 B.n436 B.t2 11.9787
R960 B.n25 B.t4 11.9787
R961 B.n527 B.n73 10.6151
R962 B.n100 B.n73 10.6151
R963 B.n101 B.n100 10.6151
R964 B.n104 B.n101 10.6151
R965 B.n105 B.n104 10.6151
R966 B.n108 B.n105 10.6151
R967 B.n109 B.n108 10.6151
R968 B.n112 B.n109 10.6151
R969 B.n113 B.n112 10.6151
R970 B.n116 B.n113 10.6151
R971 B.n117 B.n116 10.6151
R972 B.n120 B.n117 10.6151
R973 B.n121 B.n120 10.6151
R974 B.n124 B.n121 10.6151
R975 B.n129 B.n126 10.6151
R976 B.n130 B.n129 10.6151
R977 B.n133 B.n130 10.6151
R978 B.n134 B.n133 10.6151
R979 B.n137 B.n134 10.6151
R980 B.n138 B.n137 10.6151
R981 B.n141 B.n138 10.6151
R982 B.n142 B.n141 10.6151
R983 B.n145 B.n142 10.6151
R984 B.n150 B.n147 10.6151
R985 B.n151 B.n150 10.6151
R986 B.n154 B.n151 10.6151
R987 B.n155 B.n154 10.6151
R988 B.n158 B.n155 10.6151
R989 B.n159 B.n158 10.6151
R990 B.n162 B.n159 10.6151
R991 B.n163 B.n162 10.6151
R992 B.n166 B.n163 10.6151
R993 B.n167 B.n166 10.6151
R994 B.n170 B.n167 10.6151
R995 B.n172 B.n170 10.6151
R996 B.n173 B.n172 10.6151
R997 B.n521 B.n173 10.6151
R998 B.n360 B.n245 10.6151
R999 B.n361 B.n360 10.6151
R1000 B.n362 B.n361 10.6151
R1001 B.n362 B.n236 10.6151
R1002 B.n372 B.n236 10.6151
R1003 B.n373 B.n372 10.6151
R1004 B.n374 B.n373 10.6151
R1005 B.n374 B.n229 10.6151
R1006 B.n384 B.n229 10.6151
R1007 B.n385 B.n384 10.6151
R1008 B.n386 B.n385 10.6151
R1009 B.n386 B.n221 10.6151
R1010 B.n396 B.n221 10.6151
R1011 B.n397 B.n396 10.6151
R1012 B.n398 B.n397 10.6151
R1013 B.n398 B.n213 10.6151
R1014 B.n408 B.n213 10.6151
R1015 B.n409 B.n408 10.6151
R1016 B.n410 B.n409 10.6151
R1017 B.n410 B.n205 10.6151
R1018 B.n420 B.n205 10.6151
R1019 B.n421 B.n420 10.6151
R1020 B.n422 B.n421 10.6151
R1021 B.n422 B.n197 10.6151
R1022 B.n432 B.n197 10.6151
R1023 B.n433 B.n432 10.6151
R1024 B.n434 B.n433 10.6151
R1025 B.n434 B.n190 10.6151
R1026 B.n445 B.n190 10.6151
R1027 B.n446 B.n445 10.6151
R1028 B.n447 B.n446 10.6151
R1029 B.n447 B.n181 10.6151
R1030 B.n457 B.n181 10.6151
R1031 B.n458 B.n457 10.6151
R1032 B.n460 B.n458 10.6151
R1033 B.n460 B.n459 10.6151
R1034 B.n459 B.n174 10.6151
R1035 B.n471 B.n174 10.6151
R1036 B.n472 B.n471 10.6151
R1037 B.n473 B.n472 10.6151
R1038 B.n474 B.n473 10.6151
R1039 B.n476 B.n474 10.6151
R1040 B.n477 B.n476 10.6151
R1041 B.n478 B.n477 10.6151
R1042 B.n479 B.n478 10.6151
R1043 B.n481 B.n479 10.6151
R1044 B.n482 B.n481 10.6151
R1045 B.n483 B.n482 10.6151
R1046 B.n484 B.n483 10.6151
R1047 B.n486 B.n484 10.6151
R1048 B.n487 B.n486 10.6151
R1049 B.n488 B.n487 10.6151
R1050 B.n489 B.n488 10.6151
R1051 B.n491 B.n489 10.6151
R1052 B.n492 B.n491 10.6151
R1053 B.n493 B.n492 10.6151
R1054 B.n494 B.n493 10.6151
R1055 B.n496 B.n494 10.6151
R1056 B.n497 B.n496 10.6151
R1057 B.n498 B.n497 10.6151
R1058 B.n499 B.n498 10.6151
R1059 B.n501 B.n499 10.6151
R1060 B.n502 B.n501 10.6151
R1061 B.n503 B.n502 10.6151
R1062 B.n504 B.n503 10.6151
R1063 B.n506 B.n504 10.6151
R1064 B.n507 B.n506 10.6151
R1065 B.n508 B.n507 10.6151
R1066 B.n509 B.n508 10.6151
R1067 B.n511 B.n509 10.6151
R1068 B.n512 B.n511 10.6151
R1069 B.n513 B.n512 10.6151
R1070 B.n514 B.n513 10.6151
R1071 B.n516 B.n514 10.6151
R1072 B.n517 B.n516 10.6151
R1073 B.n518 B.n517 10.6151
R1074 B.n519 B.n518 10.6151
R1075 B.n520 B.n519 10.6151
R1076 B.n354 B.n249 10.6151
R1077 B.n349 B.n249 10.6151
R1078 B.n349 B.n348 10.6151
R1079 B.n348 B.n347 10.6151
R1080 B.n347 B.n344 10.6151
R1081 B.n344 B.n343 10.6151
R1082 B.n343 B.n340 10.6151
R1083 B.n340 B.n339 10.6151
R1084 B.n339 B.n336 10.6151
R1085 B.n336 B.n335 10.6151
R1086 B.n335 B.n332 10.6151
R1087 B.n332 B.n331 10.6151
R1088 B.n331 B.n328 10.6151
R1089 B.n328 B.n327 10.6151
R1090 B.n324 B.n323 10.6151
R1091 B.n323 B.n320 10.6151
R1092 B.n320 B.n319 10.6151
R1093 B.n319 B.n316 10.6151
R1094 B.n316 B.n315 10.6151
R1095 B.n315 B.n312 10.6151
R1096 B.n312 B.n311 10.6151
R1097 B.n311 B.n308 10.6151
R1098 B.n308 B.n307 10.6151
R1099 B.n304 B.n303 10.6151
R1100 B.n303 B.n300 10.6151
R1101 B.n300 B.n299 10.6151
R1102 B.n299 B.n296 10.6151
R1103 B.n296 B.n295 10.6151
R1104 B.n295 B.n292 10.6151
R1105 B.n292 B.n291 10.6151
R1106 B.n291 B.n288 10.6151
R1107 B.n288 B.n287 10.6151
R1108 B.n287 B.n284 10.6151
R1109 B.n284 B.n283 10.6151
R1110 B.n283 B.n280 10.6151
R1111 B.n280 B.n279 10.6151
R1112 B.n279 B.n277 10.6151
R1113 B.n356 B.n355 10.6151
R1114 B.n356 B.n241 10.6151
R1115 B.n366 B.n241 10.6151
R1116 B.n367 B.n366 10.6151
R1117 B.n368 B.n367 10.6151
R1118 B.n368 B.n233 10.6151
R1119 B.n378 B.n233 10.6151
R1120 B.n379 B.n378 10.6151
R1121 B.n380 B.n379 10.6151
R1122 B.n380 B.n225 10.6151
R1123 B.n390 B.n225 10.6151
R1124 B.n391 B.n390 10.6151
R1125 B.n392 B.n391 10.6151
R1126 B.n392 B.n217 10.6151
R1127 B.n402 B.n217 10.6151
R1128 B.n403 B.n402 10.6151
R1129 B.n404 B.n403 10.6151
R1130 B.n404 B.n209 10.6151
R1131 B.n414 B.n209 10.6151
R1132 B.n415 B.n414 10.6151
R1133 B.n416 B.n415 10.6151
R1134 B.n416 B.n201 10.6151
R1135 B.n426 B.n201 10.6151
R1136 B.n427 B.n426 10.6151
R1137 B.n428 B.n427 10.6151
R1138 B.n428 B.n193 10.6151
R1139 B.n439 B.n193 10.6151
R1140 B.n440 B.n439 10.6151
R1141 B.n441 B.n440 10.6151
R1142 B.n441 B.n186 10.6151
R1143 B.n451 B.n186 10.6151
R1144 B.n452 B.n451 10.6151
R1145 B.n453 B.n452 10.6151
R1146 B.n453 B.n178 10.6151
R1147 B.n464 B.n178 10.6151
R1148 B.n465 B.n464 10.6151
R1149 B.n466 B.n465 10.6151
R1150 B.n466 B.n0 10.6151
R1151 B.n601 B.n1 10.6151
R1152 B.n601 B.n600 10.6151
R1153 B.n600 B.n599 10.6151
R1154 B.n599 B.n10 10.6151
R1155 B.n593 B.n10 10.6151
R1156 B.n593 B.n592 10.6151
R1157 B.n592 B.n591 10.6151
R1158 B.n591 B.n17 10.6151
R1159 B.n585 B.n17 10.6151
R1160 B.n585 B.n584 10.6151
R1161 B.n584 B.n583 10.6151
R1162 B.n583 B.n23 10.6151
R1163 B.n577 B.n23 10.6151
R1164 B.n577 B.n576 10.6151
R1165 B.n576 B.n575 10.6151
R1166 B.n575 B.n31 10.6151
R1167 B.n569 B.n31 10.6151
R1168 B.n569 B.n568 10.6151
R1169 B.n568 B.n567 10.6151
R1170 B.n567 B.n38 10.6151
R1171 B.n561 B.n38 10.6151
R1172 B.n561 B.n560 10.6151
R1173 B.n560 B.n559 10.6151
R1174 B.n559 B.n45 10.6151
R1175 B.n553 B.n45 10.6151
R1176 B.n553 B.n552 10.6151
R1177 B.n552 B.n551 10.6151
R1178 B.n551 B.n52 10.6151
R1179 B.n545 B.n52 10.6151
R1180 B.n545 B.n544 10.6151
R1181 B.n544 B.n543 10.6151
R1182 B.n543 B.n59 10.6151
R1183 B.n537 B.n59 10.6151
R1184 B.n537 B.n536 10.6151
R1185 B.n536 B.n535 10.6151
R1186 B.n535 B.n66 10.6151
R1187 B.n529 B.n66 10.6151
R1188 B.n529 B.n528 10.6151
R1189 B.n125 B.n124 9.36635
R1190 B.n147 B.n146 9.36635
R1191 B.n327 B.n273 9.36635
R1192 B.n304 B.n276 9.36635
R1193 B.t5 B.n203 3.99324
R1194 B.n572 B.t7 3.99324
R1195 B.n607 B.n0 2.81026
R1196 B.n607 B.n1 2.81026
R1197 B.n126 B.n125 1.24928
R1198 B.n146 B.n145 1.24928
R1199 B.n324 B.n273 1.24928
R1200 B.n307 B.n276 1.24928
R1201 VN.n22 VN.n21 178.428
R1202 VN.n45 VN.n44 178.428
R1203 VN.n43 VN.n23 161.3
R1204 VN.n42 VN.n41 161.3
R1205 VN.n40 VN.n24 161.3
R1206 VN.n39 VN.n38 161.3
R1207 VN.n36 VN.n25 161.3
R1208 VN.n35 VN.n34 161.3
R1209 VN.n33 VN.n26 161.3
R1210 VN.n32 VN.n31 161.3
R1211 VN.n30 VN.n27 161.3
R1212 VN.n20 VN.n0 161.3
R1213 VN.n19 VN.n18 161.3
R1214 VN.n17 VN.n1 161.3
R1215 VN.n16 VN.n15 161.3
R1216 VN.n13 VN.n2 161.3
R1217 VN.n12 VN.n11 161.3
R1218 VN.n10 VN.n3 161.3
R1219 VN.n9 VN.n8 161.3
R1220 VN.n7 VN.n4 161.3
R1221 VN.n5 VN.t2 72.6378
R1222 VN.n28 VN.t3 72.6378
R1223 VN.n6 VN.n5 65.2126
R1224 VN.n29 VN.n28 65.2126
R1225 VN.n19 VN.n1 50.2061
R1226 VN.n42 VN.n24 50.2061
R1227 VN.n6 VN.t5 40.7118
R1228 VN.n14 VN.t1 40.7118
R1229 VN.n21 VN.t4 40.7118
R1230 VN.n29 VN.t7 40.7118
R1231 VN.n37 VN.t0 40.7118
R1232 VN.n44 VN.t6 40.7118
R1233 VN VN.n45 40.5175
R1234 VN.n8 VN.n3 40.4934
R1235 VN.n12 VN.n3 40.4934
R1236 VN.n31 VN.n26 40.4934
R1237 VN.n35 VN.n26 40.4934
R1238 VN.n15 VN.n1 30.7807
R1239 VN.n38 VN.n24 30.7807
R1240 VN.n8 VN.n7 24.4675
R1241 VN.n13 VN.n12 24.4675
R1242 VN.n20 VN.n19 24.4675
R1243 VN.n31 VN.n30 24.4675
R1244 VN.n36 VN.n35 24.4675
R1245 VN.n43 VN.n42 24.4675
R1246 VN.n15 VN.n14 22.0208
R1247 VN.n38 VN.n37 22.0208
R1248 VN.n28 VN.n27 18.1539
R1249 VN.n5 VN.n4 18.1539
R1250 VN.n21 VN.n20 7.3406
R1251 VN.n44 VN.n43 7.3406
R1252 VN.n7 VN.n6 2.4472
R1253 VN.n14 VN.n13 2.4472
R1254 VN.n30 VN.n29 2.4472
R1255 VN.n37 VN.n36 2.4472
R1256 VN.n45 VN.n23 0.189894
R1257 VN.n41 VN.n23 0.189894
R1258 VN.n41 VN.n40 0.189894
R1259 VN.n40 VN.n39 0.189894
R1260 VN.n39 VN.n25 0.189894
R1261 VN.n34 VN.n25 0.189894
R1262 VN.n34 VN.n33 0.189894
R1263 VN.n33 VN.n32 0.189894
R1264 VN.n32 VN.n27 0.189894
R1265 VN.n9 VN.n4 0.189894
R1266 VN.n10 VN.n9 0.189894
R1267 VN.n11 VN.n10 0.189894
R1268 VN.n11 VN.n2 0.189894
R1269 VN.n16 VN.n2 0.189894
R1270 VN.n17 VN.n16 0.189894
R1271 VN.n18 VN.n17 0.189894
R1272 VN.n18 VN.n0 0.189894
R1273 VN.n22 VN.n0 0.189894
R1274 VN VN.n22 0.0516364
R1275 VDD2.n2 VDD2.n1 86.1388
R1276 VDD2.n2 VDD2.n0 86.1388
R1277 VDD2 VDD2.n5 86.1361
R1278 VDD2.n4 VDD2.n3 85.2892
R1279 VDD2.n4 VDD2.n2 34.4394
R1280 VDD2.n5 VDD2.t0 6.62257
R1281 VDD2.n5 VDD2.t4 6.62257
R1282 VDD2.n3 VDD2.t1 6.62257
R1283 VDD2.n3 VDD2.t7 6.62257
R1284 VDD2.n1 VDD2.t6 6.62257
R1285 VDD2.n1 VDD2.t3 6.62257
R1286 VDD2.n0 VDD2.t5 6.62257
R1287 VDD2.n0 VDD2.t2 6.62257
R1288 VDD2 VDD2.n4 0.963862
C0 VDD2 VDD1 1.3444f
C1 VDD2 VP 0.43681f
C2 VDD2 VN 2.30484f
C3 VDD2 VTAIL 4.4917f
C4 VP VDD1 2.58488f
C5 VDD1 VN 0.155015f
C6 VP VN 4.98269f
C7 VTAIL VDD1 4.44285f
C8 VTAIL VP 2.99549f
C9 VTAIL VN 2.98138f
C10 VDD2 B 3.824444f
C11 VDD1 B 4.176732f
C12 VTAIL B 4.250404f
C13 VN B 11.465031f
C14 VP B 10.011031f
C15 VDD2.t5 B 0.057829f
C16 VDD2.t2 B 0.057829f
C17 VDD2.n0 B 0.430251f
C18 VDD2.t6 B 0.057829f
C19 VDD2.t3 B 0.057829f
C20 VDD2.n1 B 0.430251f
C21 VDD2.n2 B 2.17825f
C22 VDD2.t1 B 0.057829f
C23 VDD2.t7 B 0.057829f
C24 VDD2.n3 B 0.42624f
C25 VDD2.n4 B 1.89764f
C26 VDD2.t0 B 0.057829f
C27 VDD2.t4 B 0.057829f
C28 VDD2.n5 B 0.430228f
C29 VN.n0 B 0.033475f
C30 VN.t4 B 0.441139f
C31 VN.n1 B 0.031624f
C32 VN.n2 B 0.033475f
C33 VN.t1 B 0.441139f
C34 VN.n3 B 0.027062f
C35 VN.n4 B 0.217428f
C36 VN.t5 B 0.441139f
C37 VN.t2 B 0.592492f
C38 VN.n5 B 0.266144f
C39 VN.n6 B 0.256425f
C40 VN.n7 B 0.034668f
C41 VN.n8 B 0.066532f
C42 VN.n9 B 0.033475f
C43 VN.n10 B 0.033475f
C44 VN.n11 B 0.033475f
C45 VN.n12 B 0.066532f
C46 VN.n13 B 0.034668f
C47 VN.n14 B 0.196299f
C48 VN.n15 B 0.063983f
C49 VN.n16 B 0.033475f
C50 VN.n17 B 0.033475f
C51 VN.n18 B 0.033475f
C52 VN.n19 B 0.061439f
C53 VN.n20 B 0.040828f
C54 VN.n21 B 0.27609f
C55 VN.n22 B 0.034414f
C56 VN.n23 B 0.033475f
C57 VN.t6 B 0.441139f
C58 VN.n24 B 0.031624f
C59 VN.n25 B 0.033475f
C60 VN.t0 B 0.441139f
C61 VN.n26 B 0.027062f
C62 VN.n27 B 0.217428f
C63 VN.t7 B 0.441139f
C64 VN.t3 B 0.592492f
C65 VN.n28 B 0.266144f
C66 VN.n29 B 0.256425f
C67 VN.n30 B 0.034668f
C68 VN.n31 B 0.066532f
C69 VN.n32 B 0.033475f
C70 VN.n33 B 0.033475f
C71 VN.n34 B 0.033475f
C72 VN.n35 B 0.066532f
C73 VN.n36 B 0.034668f
C74 VN.n37 B 0.196299f
C75 VN.n38 B 0.063983f
C76 VN.n39 B 0.033475f
C77 VN.n40 B 0.033475f
C78 VN.n41 B 0.033475f
C79 VN.n42 B 0.061439f
C80 VN.n43 B 0.040828f
C81 VN.n44 B 0.27609f
C82 VN.n45 B 1.31009f
C83 VTAIL.t4 B 0.062339f
C84 VTAIL.t7 B 0.062339f
C85 VTAIL.n0 B 0.411878f
C86 VTAIL.n1 B 0.37141f
C87 VTAIL.t0 B 0.53616f
C88 VTAIL.n2 B 0.452138f
C89 VTAIL.t10 B 0.53616f
C90 VTAIL.n3 B 0.452138f
C91 VTAIL.t12 B 0.062339f
C92 VTAIL.t14 B 0.062339f
C93 VTAIL.n4 B 0.411878f
C94 VTAIL.n5 B 0.520368f
C95 VTAIL.t9 B 0.53616f
C96 VTAIL.n6 B 1.14362f
C97 VTAIL.t6 B 0.536162f
C98 VTAIL.n7 B 1.14362f
C99 VTAIL.t5 B 0.062339f
C100 VTAIL.t2 B 0.062339f
C101 VTAIL.n8 B 0.411879f
C102 VTAIL.n9 B 0.520366f
C103 VTAIL.t1 B 0.536162f
C104 VTAIL.n10 B 0.452136f
C105 VTAIL.t15 B 0.536162f
C106 VTAIL.n11 B 0.452136f
C107 VTAIL.t11 B 0.062339f
C108 VTAIL.t8 B 0.062339f
C109 VTAIL.n12 B 0.411879f
C110 VTAIL.n13 B 0.520366f
C111 VTAIL.t13 B 0.53616f
C112 VTAIL.n14 B 1.14362f
C113 VTAIL.t3 B 0.53616f
C114 VTAIL.n15 B 1.13867f
C115 VDD1.t1 B 0.058749f
C116 VDD1.t6 B 0.058749f
C117 VDD1.n0 B 0.437728f
C118 VDD1.t0 B 0.058749f
C119 VDD1.t7 B 0.058749f
C120 VDD1.n1 B 0.437094f
C121 VDD1.t4 B 0.058749f
C122 VDD1.t2 B 0.058749f
C123 VDD1.n2 B 0.437094f
C124 VDD1.n3 B 2.26542f
C125 VDD1.t3 B 0.058749f
C126 VDD1.t5 B 0.058749f
C127 VDD1.n4 B 0.433018f
C128 VDD1.n5 B 1.95782f
C129 VP.n0 B 0.034608f
C130 VP.t5 B 0.456072f
C131 VP.n1 B 0.032694f
C132 VP.n2 B 0.034608f
C133 VP.t1 B 0.456072f
C134 VP.n3 B 0.027978f
C135 VP.n4 B 0.034608f
C136 VP.t3 B 0.456072f
C137 VP.n5 B 0.032694f
C138 VP.n6 B 0.034608f
C139 VP.t6 B 0.456072f
C140 VP.n7 B 0.034608f
C141 VP.t2 B 0.456072f
C142 VP.n8 B 0.032694f
C143 VP.n9 B 0.034608f
C144 VP.t7 B 0.456072f
C145 VP.n10 B 0.027978f
C146 VP.n11 B 0.224788f
C147 VP.t4 B 0.456072f
C148 VP.t0 B 0.612548f
C149 VP.n12 B 0.275152f
C150 VP.n13 B 0.265105f
C151 VP.n14 B 0.035841f
C152 VP.n15 B 0.068784f
C153 VP.n16 B 0.034608f
C154 VP.n17 B 0.034608f
C155 VP.n18 B 0.034608f
C156 VP.n19 B 0.068784f
C157 VP.n20 B 0.035841f
C158 VP.n21 B 0.202943f
C159 VP.n22 B 0.066148f
C160 VP.n23 B 0.034608f
C161 VP.n24 B 0.034608f
C162 VP.n25 B 0.034608f
C163 VP.n26 B 0.063519f
C164 VP.n27 B 0.04221f
C165 VP.n28 B 0.285435f
C166 VP.n29 B 1.33165f
C167 VP.n30 B 1.36264f
C168 VP.n31 B 0.285435f
C169 VP.n32 B 0.04221f
C170 VP.n33 B 0.063519f
C171 VP.n34 B 0.034608f
C172 VP.n35 B 0.034608f
C173 VP.n36 B 0.034608f
C174 VP.n37 B 0.066148f
C175 VP.n38 B 0.202943f
C176 VP.n39 B 0.035841f
C177 VP.n40 B 0.068784f
C178 VP.n41 B 0.034608f
C179 VP.n42 B 0.034608f
C180 VP.n43 B 0.034608f
C181 VP.n44 B 0.068784f
C182 VP.n45 B 0.035841f
C183 VP.n46 B 0.202943f
C184 VP.n47 B 0.066148f
C185 VP.n48 B 0.034608f
C186 VP.n49 B 0.034608f
C187 VP.n50 B 0.034608f
C188 VP.n51 B 0.063519f
C189 VP.n52 B 0.04221f
C190 VP.n53 B 0.285435f
C191 VP.n54 B 0.035579f
.ends

