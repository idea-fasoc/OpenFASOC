* NGSPICE file created from diff_pair_sample_0458.ext - technology: sky130A

.subckt diff_pair_sample_0458 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4486 pd=15.17 as=5.7876 ps=30.46 w=14.84 l=3.68
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=0 ps=0 w=14.84 l=3.68
X2 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4486 pd=15.17 as=5.7876 ps=30.46 w=14.84 l=3.68
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=0 ps=0 w=14.84 l=3.68
X4 VTAIL.t5 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=2.4486 ps=15.17 w=14.84 l=3.68
X5 VTAIL.t7 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=2.4486 ps=15.17 w=14.84 l=3.68
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=0 ps=0 w=14.84 l=3.68
X7 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4486 pd=15.17 as=5.7876 ps=30.46 w=14.84 l=3.68
X8 VDD2.t0 VN.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4486 pd=15.17 as=5.7876 ps=30.46 w=14.84 l=3.68
X9 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=2.4486 ps=15.17 w=14.84 l=3.68
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=0 ps=0 w=14.84 l=3.68
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7876 pd=30.46 as=2.4486 ps=15.17 w=14.84 l=3.68
R0 VN.n1 VN.t3 130.389
R1 VN.n0 VN.t1 130.389
R2 VN.n0 VN.t0 129.067
R3 VN.n1 VN.t2 129.067
R4 VN VN.n1 53.8502
R5 VN VN.n0 1.94492
R6 VTAIL.n650 VTAIL.n574 289.615
R7 VTAIL.n76 VTAIL.n0 289.615
R8 VTAIL.n158 VTAIL.n82 289.615
R9 VTAIL.n240 VTAIL.n164 289.615
R10 VTAIL.n568 VTAIL.n492 289.615
R11 VTAIL.n486 VTAIL.n410 289.615
R12 VTAIL.n404 VTAIL.n328 289.615
R13 VTAIL.n322 VTAIL.n246 289.615
R14 VTAIL.n601 VTAIL.n600 185
R15 VTAIL.n598 VTAIL.n597 185
R16 VTAIL.n607 VTAIL.n606 185
R17 VTAIL.n609 VTAIL.n608 185
R18 VTAIL.n594 VTAIL.n593 185
R19 VTAIL.n615 VTAIL.n614 185
R20 VTAIL.n617 VTAIL.n616 185
R21 VTAIL.n590 VTAIL.n589 185
R22 VTAIL.n623 VTAIL.n622 185
R23 VTAIL.n625 VTAIL.n624 185
R24 VTAIL.n586 VTAIL.n585 185
R25 VTAIL.n631 VTAIL.n630 185
R26 VTAIL.n633 VTAIL.n632 185
R27 VTAIL.n582 VTAIL.n581 185
R28 VTAIL.n639 VTAIL.n638 185
R29 VTAIL.n642 VTAIL.n641 185
R30 VTAIL.n640 VTAIL.n578 185
R31 VTAIL.n647 VTAIL.n577 185
R32 VTAIL.n649 VTAIL.n648 185
R33 VTAIL.n651 VTAIL.n650 185
R34 VTAIL.n27 VTAIL.n26 185
R35 VTAIL.n24 VTAIL.n23 185
R36 VTAIL.n33 VTAIL.n32 185
R37 VTAIL.n35 VTAIL.n34 185
R38 VTAIL.n20 VTAIL.n19 185
R39 VTAIL.n41 VTAIL.n40 185
R40 VTAIL.n43 VTAIL.n42 185
R41 VTAIL.n16 VTAIL.n15 185
R42 VTAIL.n49 VTAIL.n48 185
R43 VTAIL.n51 VTAIL.n50 185
R44 VTAIL.n12 VTAIL.n11 185
R45 VTAIL.n57 VTAIL.n56 185
R46 VTAIL.n59 VTAIL.n58 185
R47 VTAIL.n8 VTAIL.n7 185
R48 VTAIL.n65 VTAIL.n64 185
R49 VTAIL.n68 VTAIL.n67 185
R50 VTAIL.n66 VTAIL.n4 185
R51 VTAIL.n73 VTAIL.n3 185
R52 VTAIL.n75 VTAIL.n74 185
R53 VTAIL.n77 VTAIL.n76 185
R54 VTAIL.n109 VTAIL.n108 185
R55 VTAIL.n106 VTAIL.n105 185
R56 VTAIL.n115 VTAIL.n114 185
R57 VTAIL.n117 VTAIL.n116 185
R58 VTAIL.n102 VTAIL.n101 185
R59 VTAIL.n123 VTAIL.n122 185
R60 VTAIL.n125 VTAIL.n124 185
R61 VTAIL.n98 VTAIL.n97 185
R62 VTAIL.n131 VTAIL.n130 185
R63 VTAIL.n133 VTAIL.n132 185
R64 VTAIL.n94 VTAIL.n93 185
R65 VTAIL.n139 VTAIL.n138 185
R66 VTAIL.n141 VTAIL.n140 185
R67 VTAIL.n90 VTAIL.n89 185
R68 VTAIL.n147 VTAIL.n146 185
R69 VTAIL.n150 VTAIL.n149 185
R70 VTAIL.n148 VTAIL.n86 185
R71 VTAIL.n155 VTAIL.n85 185
R72 VTAIL.n157 VTAIL.n156 185
R73 VTAIL.n159 VTAIL.n158 185
R74 VTAIL.n191 VTAIL.n190 185
R75 VTAIL.n188 VTAIL.n187 185
R76 VTAIL.n197 VTAIL.n196 185
R77 VTAIL.n199 VTAIL.n198 185
R78 VTAIL.n184 VTAIL.n183 185
R79 VTAIL.n205 VTAIL.n204 185
R80 VTAIL.n207 VTAIL.n206 185
R81 VTAIL.n180 VTAIL.n179 185
R82 VTAIL.n213 VTAIL.n212 185
R83 VTAIL.n215 VTAIL.n214 185
R84 VTAIL.n176 VTAIL.n175 185
R85 VTAIL.n221 VTAIL.n220 185
R86 VTAIL.n223 VTAIL.n222 185
R87 VTAIL.n172 VTAIL.n171 185
R88 VTAIL.n229 VTAIL.n228 185
R89 VTAIL.n232 VTAIL.n231 185
R90 VTAIL.n230 VTAIL.n168 185
R91 VTAIL.n237 VTAIL.n167 185
R92 VTAIL.n239 VTAIL.n238 185
R93 VTAIL.n241 VTAIL.n240 185
R94 VTAIL.n569 VTAIL.n568 185
R95 VTAIL.n567 VTAIL.n566 185
R96 VTAIL.n565 VTAIL.n495 185
R97 VTAIL.n499 VTAIL.n496 185
R98 VTAIL.n560 VTAIL.n559 185
R99 VTAIL.n558 VTAIL.n557 185
R100 VTAIL.n501 VTAIL.n500 185
R101 VTAIL.n552 VTAIL.n551 185
R102 VTAIL.n550 VTAIL.n549 185
R103 VTAIL.n505 VTAIL.n504 185
R104 VTAIL.n544 VTAIL.n543 185
R105 VTAIL.n542 VTAIL.n541 185
R106 VTAIL.n509 VTAIL.n508 185
R107 VTAIL.n536 VTAIL.n535 185
R108 VTAIL.n534 VTAIL.n533 185
R109 VTAIL.n513 VTAIL.n512 185
R110 VTAIL.n528 VTAIL.n527 185
R111 VTAIL.n526 VTAIL.n525 185
R112 VTAIL.n517 VTAIL.n516 185
R113 VTAIL.n520 VTAIL.n519 185
R114 VTAIL.n487 VTAIL.n486 185
R115 VTAIL.n485 VTAIL.n484 185
R116 VTAIL.n483 VTAIL.n413 185
R117 VTAIL.n417 VTAIL.n414 185
R118 VTAIL.n478 VTAIL.n477 185
R119 VTAIL.n476 VTAIL.n475 185
R120 VTAIL.n419 VTAIL.n418 185
R121 VTAIL.n470 VTAIL.n469 185
R122 VTAIL.n468 VTAIL.n467 185
R123 VTAIL.n423 VTAIL.n422 185
R124 VTAIL.n462 VTAIL.n461 185
R125 VTAIL.n460 VTAIL.n459 185
R126 VTAIL.n427 VTAIL.n426 185
R127 VTAIL.n454 VTAIL.n453 185
R128 VTAIL.n452 VTAIL.n451 185
R129 VTAIL.n431 VTAIL.n430 185
R130 VTAIL.n446 VTAIL.n445 185
R131 VTAIL.n444 VTAIL.n443 185
R132 VTAIL.n435 VTAIL.n434 185
R133 VTAIL.n438 VTAIL.n437 185
R134 VTAIL.n405 VTAIL.n404 185
R135 VTAIL.n403 VTAIL.n402 185
R136 VTAIL.n401 VTAIL.n331 185
R137 VTAIL.n335 VTAIL.n332 185
R138 VTAIL.n396 VTAIL.n395 185
R139 VTAIL.n394 VTAIL.n393 185
R140 VTAIL.n337 VTAIL.n336 185
R141 VTAIL.n388 VTAIL.n387 185
R142 VTAIL.n386 VTAIL.n385 185
R143 VTAIL.n341 VTAIL.n340 185
R144 VTAIL.n380 VTAIL.n379 185
R145 VTAIL.n378 VTAIL.n377 185
R146 VTAIL.n345 VTAIL.n344 185
R147 VTAIL.n372 VTAIL.n371 185
R148 VTAIL.n370 VTAIL.n369 185
R149 VTAIL.n349 VTAIL.n348 185
R150 VTAIL.n364 VTAIL.n363 185
R151 VTAIL.n362 VTAIL.n361 185
R152 VTAIL.n353 VTAIL.n352 185
R153 VTAIL.n356 VTAIL.n355 185
R154 VTAIL.n323 VTAIL.n322 185
R155 VTAIL.n321 VTAIL.n320 185
R156 VTAIL.n319 VTAIL.n249 185
R157 VTAIL.n253 VTAIL.n250 185
R158 VTAIL.n314 VTAIL.n313 185
R159 VTAIL.n312 VTAIL.n311 185
R160 VTAIL.n255 VTAIL.n254 185
R161 VTAIL.n306 VTAIL.n305 185
R162 VTAIL.n304 VTAIL.n303 185
R163 VTAIL.n259 VTAIL.n258 185
R164 VTAIL.n298 VTAIL.n297 185
R165 VTAIL.n296 VTAIL.n295 185
R166 VTAIL.n263 VTAIL.n262 185
R167 VTAIL.n290 VTAIL.n289 185
R168 VTAIL.n288 VTAIL.n287 185
R169 VTAIL.n267 VTAIL.n266 185
R170 VTAIL.n282 VTAIL.n281 185
R171 VTAIL.n280 VTAIL.n279 185
R172 VTAIL.n271 VTAIL.n270 185
R173 VTAIL.n274 VTAIL.n273 185
R174 VTAIL.t0 VTAIL.n518 147.659
R175 VTAIL.t2 VTAIL.n436 147.659
R176 VTAIL.t6 VTAIL.n354 147.659
R177 VTAIL.t7 VTAIL.n272 147.659
R178 VTAIL.t4 VTAIL.n599 147.659
R179 VTAIL.t5 VTAIL.n25 147.659
R180 VTAIL.t3 VTAIL.n107 147.659
R181 VTAIL.t1 VTAIL.n189 147.659
R182 VTAIL.n600 VTAIL.n597 104.615
R183 VTAIL.n607 VTAIL.n597 104.615
R184 VTAIL.n608 VTAIL.n607 104.615
R185 VTAIL.n608 VTAIL.n593 104.615
R186 VTAIL.n615 VTAIL.n593 104.615
R187 VTAIL.n616 VTAIL.n615 104.615
R188 VTAIL.n616 VTAIL.n589 104.615
R189 VTAIL.n623 VTAIL.n589 104.615
R190 VTAIL.n624 VTAIL.n623 104.615
R191 VTAIL.n624 VTAIL.n585 104.615
R192 VTAIL.n631 VTAIL.n585 104.615
R193 VTAIL.n632 VTAIL.n631 104.615
R194 VTAIL.n632 VTAIL.n581 104.615
R195 VTAIL.n639 VTAIL.n581 104.615
R196 VTAIL.n641 VTAIL.n639 104.615
R197 VTAIL.n641 VTAIL.n640 104.615
R198 VTAIL.n640 VTAIL.n577 104.615
R199 VTAIL.n649 VTAIL.n577 104.615
R200 VTAIL.n650 VTAIL.n649 104.615
R201 VTAIL.n26 VTAIL.n23 104.615
R202 VTAIL.n33 VTAIL.n23 104.615
R203 VTAIL.n34 VTAIL.n33 104.615
R204 VTAIL.n34 VTAIL.n19 104.615
R205 VTAIL.n41 VTAIL.n19 104.615
R206 VTAIL.n42 VTAIL.n41 104.615
R207 VTAIL.n42 VTAIL.n15 104.615
R208 VTAIL.n49 VTAIL.n15 104.615
R209 VTAIL.n50 VTAIL.n49 104.615
R210 VTAIL.n50 VTAIL.n11 104.615
R211 VTAIL.n57 VTAIL.n11 104.615
R212 VTAIL.n58 VTAIL.n57 104.615
R213 VTAIL.n58 VTAIL.n7 104.615
R214 VTAIL.n65 VTAIL.n7 104.615
R215 VTAIL.n67 VTAIL.n65 104.615
R216 VTAIL.n67 VTAIL.n66 104.615
R217 VTAIL.n66 VTAIL.n3 104.615
R218 VTAIL.n75 VTAIL.n3 104.615
R219 VTAIL.n76 VTAIL.n75 104.615
R220 VTAIL.n108 VTAIL.n105 104.615
R221 VTAIL.n115 VTAIL.n105 104.615
R222 VTAIL.n116 VTAIL.n115 104.615
R223 VTAIL.n116 VTAIL.n101 104.615
R224 VTAIL.n123 VTAIL.n101 104.615
R225 VTAIL.n124 VTAIL.n123 104.615
R226 VTAIL.n124 VTAIL.n97 104.615
R227 VTAIL.n131 VTAIL.n97 104.615
R228 VTAIL.n132 VTAIL.n131 104.615
R229 VTAIL.n132 VTAIL.n93 104.615
R230 VTAIL.n139 VTAIL.n93 104.615
R231 VTAIL.n140 VTAIL.n139 104.615
R232 VTAIL.n140 VTAIL.n89 104.615
R233 VTAIL.n147 VTAIL.n89 104.615
R234 VTAIL.n149 VTAIL.n147 104.615
R235 VTAIL.n149 VTAIL.n148 104.615
R236 VTAIL.n148 VTAIL.n85 104.615
R237 VTAIL.n157 VTAIL.n85 104.615
R238 VTAIL.n158 VTAIL.n157 104.615
R239 VTAIL.n190 VTAIL.n187 104.615
R240 VTAIL.n197 VTAIL.n187 104.615
R241 VTAIL.n198 VTAIL.n197 104.615
R242 VTAIL.n198 VTAIL.n183 104.615
R243 VTAIL.n205 VTAIL.n183 104.615
R244 VTAIL.n206 VTAIL.n205 104.615
R245 VTAIL.n206 VTAIL.n179 104.615
R246 VTAIL.n213 VTAIL.n179 104.615
R247 VTAIL.n214 VTAIL.n213 104.615
R248 VTAIL.n214 VTAIL.n175 104.615
R249 VTAIL.n221 VTAIL.n175 104.615
R250 VTAIL.n222 VTAIL.n221 104.615
R251 VTAIL.n222 VTAIL.n171 104.615
R252 VTAIL.n229 VTAIL.n171 104.615
R253 VTAIL.n231 VTAIL.n229 104.615
R254 VTAIL.n231 VTAIL.n230 104.615
R255 VTAIL.n230 VTAIL.n167 104.615
R256 VTAIL.n239 VTAIL.n167 104.615
R257 VTAIL.n240 VTAIL.n239 104.615
R258 VTAIL.n568 VTAIL.n567 104.615
R259 VTAIL.n567 VTAIL.n495 104.615
R260 VTAIL.n499 VTAIL.n495 104.615
R261 VTAIL.n559 VTAIL.n499 104.615
R262 VTAIL.n559 VTAIL.n558 104.615
R263 VTAIL.n558 VTAIL.n500 104.615
R264 VTAIL.n551 VTAIL.n500 104.615
R265 VTAIL.n551 VTAIL.n550 104.615
R266 VTAIL.n550 VTAIL.n504 104.615
R267 VTAIL.n543 VTAIL.n504 104.615
R268 VTAIL.n543 VTAIL.n542 104.615
R269 VTAIL.n542 VTAIL.n508 104.615
R270 VTAIL.n535 VTAIL.n508 104.615
R271 VTAIL.n535 VTAIL.n534 104.615
R272 VTAIL.n534 VTAIL.n512 104.615
R273 VTAIL.n527 VTAIL.n512 104.615
R274 VTAIL.n527 VTAIL.n526 104.615
R275 VTAIL.n526 VTAIL.n516 104.615
R276 VTAIL.n519 VTAIL.n516 104.615
R277 VTAIL.n486 VTAIL.n485 104.615
R278 VTAIL.n485 VTAIL.n413 104.615
R279 VTAIL.n417 VTAIL.n413 104.615
R280 VTAIL.n477 VTAIL.n417 104.615
R281 VTAIL.n477 VTAIL.n476 104.615
R282 VTAIL.n476 VTAIL.n418 104.615
R283 VTAIL.n469 VTAIL.n418 104.615
R284 VTAIL.n469 VTAIL.n468 104.615
R285 VTAIL.n468 VTAIL.n422 104.615
R286 VTAIL.n461 VTAIL.n422 104.615
R287 VTAIL.n461 VTAIL.n460 104.615
R288 VTAIL.n460 VTAIL.n426 104.615
R289 VTAIL.n453 VTAIL.n426 104.615
R290 VTAIL.n453 VTAIL.n452 104.615
R291 VTAIL.n452 VTAIL.n430 104.615
R292 VTAIL.n445 VTAIL.n430 104.615
R293 VTAIL.n445 VTAIL.n444 104.615
R294 VTAIL.n444 VTAIL.n434 104.615
R295 VTAIL.n437 VTAIL.n434 104.615
R296 VTAIL.n404 VTAIL.n403 104.615
R297 VTAIL.n403 VTAIL.n331 104.615
R298 VTAIL.n335 VTAIL.n331 104.615
R299 VTAIL.n395 VTAIL.n335 104.615
R300 VTAIL.n395 VTAIL.n394 104.615
R301 VTAIL.n394 VTAIL.n336 104.615
R302 VTAIL.n387 VTAIL.n336 104.615
R303 VTAIL.n387 VTAIL.n386 104.615
R304 VTAIL.n386 VTAIL.n340 104.615
R305 VTAIL.n379 VTAIL.n340 104.615
R306 VTAIL.n379 VTAIL.n378 104.615
R307 VTAIL.n378 VTAIL.n344 104.615
R308 VTAIL.n371 VTAIL.n344 104.615
R309 VTAIL.n371 VTAIL.n370 104.615
R310 VTAIL.n370 VTAIL.n348 104.615
R311 VTAIL.n363 VTAIL.n348 104.615
R312 VTAIL.n363 VTAIL.n362 104.615
R313 VTAIL.n362 VTAIL.n352 104.615
R314 VTAIL.n355 VTAIL.n352 104.615
R315 VTAIL.n322 VTAIL.n321 104.615
R316 VTAIL.n321 VTAIL.n249 104.615
R317 VTAIL.n253 VTAIL.n249 104.615
R318 VTAIL.n313 VTAIL.n253 104.615
R319 VTAIL.n313 VTAIL.n312 104.615
R320 VTAIL.n312 VTAIL.n254 104.615
R321 VTAIL.n305 VTAIL.n254 104.615
R322 VTAIL.n305 VTAIL.n304 104.615
R323 VTAIL.n304 VTAIL.n258 104.615
R324 VTAIL.n297 VTAIL.n258 104.615
R325 VTAIL.n297 VTAIL.n296 104.615
R326 VTAIL.n296 VTAIL.n262 104.615
R327 VTAIL.n289 VTAIL.n262 104.615
R328 VTAIL.n289 VTAIL.n288 104.615
R329 VTAIL.n288 VTAIL.n266 104.615
R330 VTAIL.n281 VTAIL.n266 104.615
R331 VTAIL.n281 VTAIL.n280 104.615
R332 VTAIL.n280 VTAIL.n270 104.615
R333 VTAIL.n273 VTAIL.n270 104.615
R334 VTAIL.n600 VTAIL.t4 52.3082
R335 VTAIL.n26 VTAIL.t5 52.3082
R336 VTAIL.n108 VTAIL.t3 52.3082
R337 VTAIL.n190 VTAIL.t1 52.3082
R338 VTAIL.n519 VTAIL.t0 52.3082
R339 VTAIL.n437 VTAIL.t2 52.3082
R340 VTAIL.n355 VTAIL.t6 52.3082
R341 VTAIL.n273 VTAIL.t7 52.3082
R342 VTAIL.n655 VTAIL.n654 36.0641
R343 VTAIL.n81 VTAIL.n80 36.0641
R344 VTAIL.n163 VTAIL.n162 36.0641
R345 VTAIL.n245 VTAIL.n244 36.0641
R346 VTAIL.n573 VTAIL.n572 36.0641
R347 VTAIL.n491 VTAIL.n490 36.0641
R348 VTAIL.n409 VTAIL.n408 36.0641
R349 VTAIL.n327 VTAIL.n326 36.0641
R350 VTAIL.n655 VTAIL.n573 28.6169
R351 VTAIL.n327 VTAIL.n245 28.6169
R352 VTAIL.n601 VTAIL.n599 15.6677
R353 VTAIL.n27 VTAIL.n25 15.6677
R354 VTAIL.n109 VTAIL.n107 15.6677
R355 VTAIL.n191 VTAIL.n189 15.6677
R356 VTAIL.n520 VTAIL.n518 15.6677
R357 VTAIL.n438 VTAIL.n436 15.6677
R358 VTAIL.n356 VTAIL.n354 15.6677
R359 VTAIL.n274 VTAIL.n272 15.6677
R360 VTAIL.n648 VTAIL.n647 13.1884
R361 VTAIL.n74 VTAIL.n73 13.1884
R362 VTAIL.n156 VTAIL.n155 13.1884
R363 VTAIL.n238 VTAIL.n237 13.1884
R364 VTAIL.n566 VTAIL.n565 13.1884
R365 VTAIL.n484 VTAIL.n483 13.1884
R366 VTAIL.n402 VTAIL.n401 13.1884
R367 VTAIL.n320 VTAIL.n319 13.1884
R368 VTAIL.n602 VTAIL.n598 12.8005
R369 VTAIL.n646 VTAIL.n578 12.8005
R370 VTAIL.n651 VTAIL.n576 12.8005
R371 VTAIL.n28 VTAIL.n24 12.8005
R372 VTAIL.n72 VTAIL.n4 12.8005
R373 VTAIL.n77 VTAIL.n2 12.8005
R374 VTAIL.n110 VTAIL.n106 12.8005
R375 VTAIL.n154 VTAIL.n86 12.8005
R376 VTAIL.n159 VTAIL.n84 12.8005
R377 VTAIL.n192 VTAIL.n188 12.8005
R378 VTAIL.n236 VTAIL.n168 12.8005
R379 VTAIL.n241 VTAIL.n166 12.8005
R380 VTAIL.n569 VTAIL.n494 12.8005
R381 VTAIL.n564 VTAIL.n496 12.8005
R382 VTAIL.n521 VTAIL.n517 12.8005
R383 VTAIL.n487 VTAIL.n412 12.8005
R384 VTAIL.n482 VTAIL.n414 12.8005
R385 VTAIL.n439 VTAIL.n435 12.8005
R386 VTAIL.n405 VTAIL.n330 12.8005
R387 VTAIL.n400 VTAIL.n332 12.8005
R388 VTAIL.n357 VTAIL.n353 12.8005
R389 VTAIL.n323 VTAIL.n248 12.8005
R390 VTAIL.n318 VTAIL.n250 12.8005
R391 VTAIL.n275 VTAIL.n271 12.8005
R392 VTAIL.n606 VTAIL.n605 12.0247
R393 VTAIL.n643 VTAIL.n642 12.0247
R394 VTAIL.n652 VTAIL.n574 12.0247
R395 VTAIL.n32 VTAIL.n31 12.0247
R396 VTAIL.n69 VTAIL.n68 12.0247
R397 VTAIL.n78 VTAIL.n0 12.0247
R398 VTAIL.n114 VTAIL.n113 12.0247
R399 VTAIL.n151 VTAIL.n150 12.0247
R400 VTAIL.n160 VTAIL.n82 12.0247
R401 VTAIL.n196 VTAIL.n195 12.0247
R402 VTAIL.n233 VTAIL.n232 12.0247
R403 VTAIL.n242 VTAIL.n164 12.0247
R404 VTAIL.n570 VTAIL.n492 12.0247
R405 VTAIL.n561 VTAIL.n560 12.0247
R406 VTAIL.n525 VTAIL.n524 12.0247
R407 VTAIL.n488 VTAIL.n410 12.0247
R408 VTAIL.n479 VTAIL.n478 12.0247
R409 VTAIL.n443 VTAIL.n442 12.0247
R410 VTAIL.n406 VTAIL.n328 12.0247
R411 VTAIL.n397 VTAIL.n396 12.0247
R412 VTAIL.n361 VTAIL.n360 12.0247
R413 VTAIL.n324 VTAIL.n246 12.0247
R414 VTAIL.n315 VTAIL.n314 12.0247
R415 VTAIL.n279 VTAIL.n278 12.0247
R416 VTAIL.n609 VTAIL.n596 11.249
R417 VTAIL.n638 VTAIL.n580 11.249
R418 VTAIL.n35 VTAIL.n22 11.249
R419 VTAIL.n64 VTAIL.n6 11.249
R420 VTAIL.n117 VTAIL.n104 11.249
R421 VTAIL.n146 VTAIL.n88 11.249
R422 VTAIL.n199 VTAIL.n186 11.249
R423 VTAIL.n228 VTAIL.n170 11.249
R424 VTAIL.n557 VTAIL.n498 11.249
R425 VTAIL.n528 VTAIL.n515 11.249
R426 VTAIL.n475 VTAIL.n416 11.249
R427 VTAIL.n446 VTAIL.n433 11.249
R428 VTAIL.n393 VTAIL.n334 11.249
R429 VTAIL.n364 VTAIL.n351 11.249
R430 VTAIL.n311 VTAIL.n252 11.249
R431 VTAIL.n282 VTAIL.n269 11.249
R432 VTAIL.n610 VTAIL.n594 10.4732
R433 VTAIL.n637 VTAIL.n582 10.4732
R434 VTAIL.n36 VTAIL.n20 10.4732
R435 VTAIL.n63 VTAIL.n8 10.4732
R436 VTAIL.n118 VTAIL.n102 10.4732
R437 VTAIL.n145 VTAIL.n90 10.4732
R438 VTAIL.n200 VTAIL.n184 10.4732
R439 VTAIL.n227 VTAIL.n172 10.4732
R440 VTAIL.n556 VTAIL.n501 10.4732
R441 VTAIL.n529 VTAIL.n513 10.4732
R442 VTAIL.n474 VTAIL.n419 10.4732
R443 VTAIL.n447 VTAIL.n431 10.4732
R444 VTAIL.n392 VTAIL.n337 10.4732
R445 VTAIL.n365 VTAIL.n349 10.4732
R446 VTAIL.n310 VTAIL.n255 10.4732
R447 VTAIL.n283 VTAIL.n267 10.4732
R448 VTAIL.n614 VTAIL.n613 9.69747
R449 VTAIL.n634 VTAIL.n633 9.69747
R450 VTAIL.n40 VTAIL.n39 9.69747
R451 VTAIL.n60 VTAIL.n59 9.69747
R452 VTAIL.n122 VTAIL.n121 9.69747
R453 VTAIL.n142 VTAIL.n141 9.69747
R454 VTAIL.n204 VTAIL.n203 9.69747
R455 VTAIL.n224 VTAIL.n223 9.69747
R456 VTAIL.n553 VTAIL.n552 9.69747
R457 VTAIL.n533 VTAIL.n532 9.69747
R458 VTAIL.n471 VTAIL.n470 9.69747
R459 VTAIL.n451 VTAIL.n450 9.69747
R460 VTAIL.n389 VTAIL.n388 9.69747
R461 VTAIL.n369 VTAIL.n368 9.69747
R462 VTAIL.n307 VTAIL.n306 9.69747
R463 VTAIL.n287 VTAIL.n286 9.69747
R464 VTAIL.n654 VTAIL.n653 9.45567
R465 VTAIL.n80 VTAIL.n79 9.45567
R466 VTAIL.n162 VTAIL.n161 9.45567
R467 VTAIL.n244 VTAIL.n243 9.45567
R468 VTAIL.n572 VTAIL.n571 9.45567
R469 VTAIL.n490 VTAIL.n489 9.45567
R470 VTAIL.n408 VTAIL.n407 9.45567
R471 VTAIL.n326 VTAIL.n325 9.45567
R472 VTAIL.n653 VTAIL.n652 9.3005
R473 VTAIL.n576 VTAIL.n575 9.3005
R474 VTAIL.n621 VTAIL.n620 9.3005
R475 VTAIL.n619 VTAIL.n618 9.3005
R476 VTAIL.n592 VTAIL.n591 9.3005
R477 VTAIL.n613 VTAIL.n612 9.3005
R478 VTAIL.n611 VTAIL.n610 9.3005
R479 VTAIL.n596 VTAIL.n595 9.3005
R480 VTAIL.n605 VTAIL.n604 9.3005
R481 VTAIL.n603 VTAIL.n602 9.3005
R482 VTAIL.n588 VTAIL.n587 9.3005
R483 VTAIL.n627 VTAIL.n626 9.3005
R484 VTAIL.n629 VTAIL.n628 9.3005
R485 VTAIL.n584 VTAIL.n583 9.3005
R486 VTAIL.n635 VTAIL.n634 9.3005
R487 VTAIL.n637 VTAIL.n636 9.3005
R488 VTAIL.n580 VTAIL.n579 9.3005
R489 VTAIL.n644 VTAIL.n643 9.3005
R490 VTAIL.n646 VTAIL.n645 9.3005
R491 VTAIL.n79 VTAIL.n78 9.3005
R492 VTAIL.n2 VTAIL.n1 9.3005
R493 VTAIL.n47 VTAIL.n46 9.3005
R494 VTAIL.n45 VTAIL.n44 9.3005
R495 VTAIL.n18 VTAIL.n17 9.3005
R496 VTAIL.n39 VTAIL.n38 9.3005
R497 VTAIL.n37 VTAIL.n36 9.3005
R498 VTAIL.n22 VTAIL.n21 9.3005
R499 VTAIL.n31 VTAIL.n30 9.3005
R500 VTAIL.n29 VTAIL.n28 9.3005
R501 VTAIL.n14 VTAIL.n13 9.3005
R502 VTAIL.n53 VTAIL.n52 9.3005
R503 VTAIL.n55 VTAIL.n54 9.3005
R504 VTAIL.n10 VTAIL.n9 9.3005
R505 VTAIL.n61 VTAIL.n60 9.3005
R506 VTAIL.n63 VTAIL.n62 9.3005
R507 VTAIL.n6 VTAIL.n5 9.3005
R508 VTAIL.n70 VTAIL.n69 9.3005
R509 VTAIL.n72 VTAIL.n71 9.3005
R510 VTAIL.n161 VTAIL.n160 9.3005
R511 VTAIL.n84 VTAIL.n83 9.3005
R512 VTAIL.n129 VTAIL.n128 9.3005
R513 VTAIL.n127 VTAIL.n126 9.3005
R514 VTAIL.n100 VTAIL.n99 9.3005
R515 VTAIL.n121 VTAIL.n120 9.3005
R516 VTAIL.n119 VTAIL.n118 9.3005
R517 VTAIL.n104 VTAIL.n103 9.3005
R518 VTAIL.n113 VTAIL.n112 9.3005
R519 VTAIL.n111 VTAIL.n110 9.3005
R520 VTAIL.n96 VTAIL.n95 9.3005
R521 VTAIL.n135 VTAIL.n134 9.3005
R522 VTAIL.n137 VTAIL.n136 9.3005
R523 VTAIL.n92 VTAIL.n91 9.3005
R524 VTAIL.n143 VTAIL.n142 9.3005
R525 VTAIL.n145 VTAIL.n144 9.3005
R526 VTAIL.n88 VTAIL.n87 9.3005
R527 VTAIL.n152 VTAIL.n151 9.3005
R528 VTAIL.n154 VTAIL.n153 9.3005
R529 VTAIL.n243 VTAIL.n242 9.3005
R530 VTAIL.n166 VTAIL.n165 9.3005
R531 VTAIL.n211 VTAIL.n210 9.3005
R532 VTAIL.n209 VTAIL.n208 9.3005
R533 VTAIL.n182 VTAIL.n181 9.3005
R534 VTAIL.n203 VTAIL.n202 9.3005
R535 VTAIL.n201 VTAIL.n200 9.3005
R536 VTAIL.n186 VTAIL.n185 9.3005
R537 VTAIL.n195 VTAIL.n194 9.3005
R538 VTAIL.n193 VTAIL.n192 9.3005
R539 VTAIL.n178 VTAIL.n177 9.3005
R540 VTAIL.n217 VTAIL.n216 9.3005
R541 VTAIL.n219 VTAIL.n218 9.3005
R542 VTAIL.n174 VTAIL.n173 9.3005
R543 VTAIL.n225 VTAIL.n224 9.3005
R544 VTAIL.n227 VTAIL.n226 9.3005
R545 VTAIL.n170 VTAIL.n169 9.3005
R546 VTAIL.n234 VTAIL.n233 9.3005
R547 VTAIL.n236 VTAIL.n235 9.3005
R548 VTAIL.n546 VTAIL.n545 9.3005
R549 VTAIL.n548 VTAIL.n547 9.3005
R550 VTAIL.n503 VTAIL.n502 9.3005
R551 VTAIL.n554 VTAIL.n553 9.3005
R552 VTAIL.n556 VTAIL.n555 9.3005
R553 VTAIL.n498 VTAIL.n497 9.3005
R554 VTAIL.n562 VTAIL.n561 9.3005
R555 VTAIL.n564 VTAIL.n563 9.3005
R556 VTAIL.n571 VTAIL.n570 9.3005
R557 VTAIL.n494 VTAIL.n493 9.3005
R558 VTAIL.n507 VTAIL.n506 9.3005
R559 VTAIL.n540 VTAIL.n539 9.3005
R560 VTAIL.n538 VTAIL.n537 9.3005
R561 VTAIL.n511 VTAIL.n510 9.3005
R562 VTAIL.n532 VTAIL.n531 9.3005
R563 VTAIL.n530 VTAIL.n529 9.3005
R564 VTAIL.n515 VTAIL.n514 9.3005
R565 VTAIL.n524 VTAIL.n523 9.3005
R566 VTAIL.n522 VTAIL.n521 9.3005
R567 VTAIL.n464 VTAIL.n463 9.3005
R568 VTAIL.n466 VTAIL.n465 9.3005
R569 VTAIL.n421 VTAIL.n420 9.3005
R570 VTAIL.n472 VTAIL.n471 9.3005
R571 VTAIL.n474 VTAIL.n473 9.3005
R572 VTAIL.n416 VTAIL.n415 9.3005
R573 VTAIL.n480 VTAIL.n479 9.3005
R574 VTAIL.n482 VTAIL.n481 9.3005
R575 VTAIL.n489 VTAIL.n488 9.3005
R576 VTAIL.n412 VTAIL.n411 9.3005
R577 VTAIL.n425 VTAIL.n424 9.3005
R578 VTAIL.n458 VTAIL.n457 9.3005
R579 VTAIL.n456 VTAIL.n455 9.3005
R580 VTAIL.n429 VTAIL.n428 9.3005
R581 VTAIL.n450 VTAIL.n449 9.3005
R582 VTAIL.n448 VTAIL.n447 9.3005
R583 VTAIL.n433 VTAIL.n432 9.3005
R584 VTAIL.n442 VTAIL.n441 9.3005
R585 VTAIL.n440 VTAIL.n439 9.3005
R586 VTAIL.n382 VTAIL.n381 9.3005
R587 VTAIL.n384 VTAIL.n383 9.3005
R588 VTAIL.n339 VTAIL.n338 9.3005
R589 VTAIL.n390 VTAIL.n389 9.3005
R590 VTAIL.n392 VTAIL.n391 9.3005
R591 VTAIL.n334 VTAIL.n333 9.3005
R592 VTAIL.n398 VTAIL.n397 9.3005
R593 VTAIL.n400 VTAIL.n399 9.3005
R594 VTAIL.n407 VTAIL.n406 9.3005
R595 VTAIL.n330 VTAIL.n329 9.3005
R596 VTAIL.n343 VTAIL.n342 9.3005
R597 VTAIL.n376 VTAIL.n375 9.3005
R598 VTAIL.n374 VTAIL.n373 9.3005
R599 VTAIL.n347 VTAIL.n346 9.3005
R600 VTAIL.n368 VTAIL.n367 9.3005
R601 VTAIL.n366 VTAIL.n365 9.3005
R602 VTAIL.n351 VTAIL.n350 9.3005
R603 VTAIL.n360 VTAIL.n359 9.3005
R604 VTAIL.n358 VTAIL.n357 9.3005
R605 VTAIL.n300 VTAIL.n299 9.3005
R606 VTAIL.n302 VTAIL.n301 9.3005
R607 VTAIL.n257 VTAIL.n256 9.3005
R608 VTAIL.n308 VTAIL.n307 9.3005
R609 VTAIL.n310 VTAIL.n309 9.3005
R610 VTAIL.n252 VTAIL.n251 9.3005
R611 VTAIL.n316 VTAIL.n315 9.3005
R612 VTAIL.n318 VTAIL.n317 9.3005
R613 VTAIL.n325 VTAIL.n324 9.3005
R614 VTAIL.n248 VTAIL.n247 9.3005
R615 VTAIL.n261 VTAIL.n260 9.3005
R616 VTAIL.n294 VTAIL.n293 9.3005
R617 VTAIL.n292 VTAIL.n291 9.3005
R618 VTAIL.n265 VTAIL.n264 9.3005
R619 VTAIL.n286 VTAIL.n285 9.3005
R620 VTAIL.n284 VTAIL.n283 9.3005
R621 VTAIL.n269 VTAIL.n268 9.3005
R622 VTAIL.n278 VTAIL.n277 9.3005
R623 VTAIL.n276 VTAIL.n275 9.3005
R624 VTAIL.n617 VTAIL.n592 8.92171
R625 VTAIL.n630 VTAIL.n584 8.92171
R626 VTAIL.n43 VTAIL.n18 8.92171
R627 VTAIL.n56 VTAIL.n10 8.92171
R628 VTAIL.n125 VTAIL.n100 8.92171
R629 VTAIL.n138 VTAIL.n92 8.92171
R630 VTAIL.n207 VTAIL.n182 8.92171
R631 VTAIL.n220 VTAIL.n174 8.92171
R632 VTAIL.n549 VTAIL.n503 8.92171
R633 VTAIL.n536 VTAIL.n511 8.92171
R634 VTAIL.n467 VTAIL.n421 8.92171
R635 VTAIL.n454 VTAIL.n429 8.92171
R636 VTAIL.n385 VTAIL.n339 8.92171
R637 VTAIL.n372 VTAIL.n347 8.92171
R638 VTAIL.n303 VTAIL.n257 8.92171
R639 VTAIL.n290 VTAIL.n265 8.92171
R640 VTAIL.n618 VTAIL.n590 8.14595
R641 VTAIL.n629 VTAIL.n586 8.14595
R642 VTAIL.n44 VTAIL.n16 8.14595
R643 VTAIL.n55 VTAIL.n12 8.14595
R644 VTAIL.n126 VTAIL.n98 8.14595
R645 VTAIL.n137 VTAIL.n94 8.14595
R646 VTAIL.n208 VTAIL.n180 8.14595
R647 VTAIL.n219 VTAIL.n176 8.14595
R648 VTAIL.n548 VTAIL.n505 8.14595
R649 VTAIL.n537 VTAIL.n509 8.14595
R650 VTAIL.n466 VTAIL.n423 8.14595
R651 VTAIL.n455 VTAIL.n427 8.14595
R652 VTAIL.n384 VTAIL.n341 8.14595
R653 VTAIL.n373 VTAIL.n345 8.14595
R654 VTAIL.n302 VTAIL.n259 8.14595
R655 VTAIL.n291 VTAIL.n263 8.14595
R656 VTAIL.n622 VTAIL.n621 7.3702
R657 VTAIL.n626 VTAIL.n625 7.3702
R658 VTAIL.n48 VTAIL.n47 7.3702
R659 VTAIL.n52 VTAIL.n51 7.3702
R660 VTAIL.n130 VTAIL.n129 7.3702
R661 VTAIL.n134 VTAIL.n133 7.3702
R662 VTAIL.n212 VTAIL.n211 7.3702
R663 VTAIL.n216 VTAIL.n215 7.3702
R664 VTAIL.n545 VTAIL.n544 7.3702
R665 VTAIL.n541 VTAIL.n540 7.3702
R666 VTAIL.n463 VTAIL.n462 7.3702
R667 VTAIL.n459 VTAIL.n458 7.3702
R668 VTAIL.n381 VTAIL.n380 7.3702
R669 VTAIL.n377 VTAIL.n376 7.3702
R670 VTAIL.n299 VTAIL.n298 7.3702
R671 VTAIL.n295 VTAIL.n294 7.3702
R672 VTAIL.n622 VTAIL.n588 6.59444
R673 VTAIL.n625 VTAIL.n588 6.59444
R674 VTAIL.n48 VTAIL.n14 6.59444
R675 VTAIL.n51 VTAIL.n14 6.59444
R676 VTAIL.n130 VTAIL.n96 6.59444
R677 VTAIL.n133 VTAIL.n96 6.59444
R678 VTAIL.n212 VTAIL.n178 6.59444
R679 VTAIL.n215 VTAIL.n178 6.59444
R680 VTAIL.n544 VTAIL.n507 6.59444
R681 VTAIL.n541 VTAIL.n507 6.59444
R682 VTAIL.n462 VTAIL.n425 6.59444
R683 VTAIL.n459 VTAIL.n425 6.59444
R684 VTAIL.n380 VTAIL.n343 6.59444
R685 VTAIL.n377 VTAIL.n343 6.59444
R686 VTAIL.n298 VTAIL.n261 6.59444
R687 VTAIL.n295 VTAIL.n261 6.59444
R688 VTAIL.n621 VTAIL.n590 5.81868
R689 VTAIL.n626 VTAIL.n586 5.81868
R690 VTAIL.n47 VTAIL.n16 5.81868
R691 VTAIL.n52 VTAIL.n12 5.81868
R692 VTAIL.n129 VTAIL.n98 5.81868
R693 VTAIL.n134 VTAIL.n94 5.81868
R694 VTAIL.n211 VTAIL.n180 5.81868
R695 VTAIL.n216 VTAIL.n176 5.81868
R696 VTAIL.n545 VTAIL.n505 5.81868
R697 VTAIL.n540 VTAIL.n509 5.81868
R698 VTAIL.n463 VTAIL.n423 5.81868
R699 VTAIL.n458 VTAIL.n427 5.81868
R700 VTAIL.n381 VTAIL.n341 5.81868
R701 VTAIL.n376 VTAIL.n345 5.81868
R702 VTAIL.n299 VTAIL.n259 5.81868
R703 VTAIL.n294 VTAIL.n263 5.81868
R704 VTAIL.n618 VTAIL.n617 5.04292
R705 VTAIL.n630 VTAIL.n629 5.04292
R706 VTAIL.n44 VTAIL.n43 5.04292
R707 VTAIL.n56 VTAIL.n55 5.04292
R708 VTAIL.n126 VTAIL.n125 5.04292
R709 VTAIL.n138 VTAIL.n137 5.04292
R710 VTAIL.n208 VTAIL.n207 5.04292
R711 VTAIL.n220 VTAIL.n219 5.04292
R712 VTAIL.n549 VTAIL.n548 5.04292
R713 VTAIL.n537 VTAIL.n536 5.04292
R714 VTAIL.n467 VTAIL.n466 5.04292
R715 VTAIL.n455 VTAIL.n454 5.04292
R716 VTAIL.n385 VTAIL.n384 5.04292
R717 VTAIL.n373 VTAIL.n372 5.04292
R718 VTAIL.n303 VTAIL.n302 5.04292
R719 VTAIL.n291 VTAIL.n290 5.04292
R720 VTAIL.n522 VTAIL.n518 4.38563
R721 VTAIL.n440 VTAIL.n436 4.38563
R722 VTAIL.n358 VTAIL.n354 4.38563
R723 VTAIL.n276 VTAIL.n272 4.38563
R724 VTAIL.n603 VTAIL.n599 4.38563
R725 VTAIL.n29 VTAIL.n25 4.38563
R726 VTAIL.n111 VTAIL.n107 4.38563
R727 VTAIL.n193 VTAIL.n189 4.38563
R728 VTAIL.n614 VTAIL.n592 4.26717
R729 VTAIL.n633 VTAIL.n584 4.26717
R730 VTAIL.n40 VTAIL.n18 4.26717
R731 VTAIL.n59 VTAIL.n10 4.26717
R732 VTAIL.n122 VTAIL.n100 4.26717
R733 VTAIL.n141 VTAIL.n92 4.26717
R734 VTAIL.n204 VTAIL.n182 4.26717
R735 VTAIL.n223 VTAIL.n174 4.26717
R736 VTAIL.n552 VTAIL.n503 4.26717
R737 VTAIL.n533 VTAIL.n511 4.26717
R738 VTAIL.n470 VTAIL.n421 4.26717
R739 VTAIL.n451 VTAIL.n429 4.26717
R740 VTAIL.n388 VTAIL.n339 4.26717
R741 VTAIL.n369 VTAIL.n347 4.26717
R742 VTAIL.n306 VTAIL.n257 4.26717
R743 VTAIL.n287 VTAIL.n265 4.26717
R744 VTAIL.n613 VTAIL.n594 3.49141
R745 VTAIL.n634 VTAIL.n582 3.49141
R746 VTAIL.n39 VTAIL.n20 3.49141
R747 VTAIL.n60 VTAIL.n8 3.49141
R748 VTAIL.n121 VTAIL.n102 3.49141
R749 VTAIL.n142 VTAIL.n90 3.49141
R750 VTAIL.n203 VTAIL.n184 3.49141
R751 VTAIL.n224 VTAIL.n172 3.49141
R752 VTAIL.n553 VTAIL.n501 3.49141
R753 VTAIL.n532 VTAIL.n513 3.49141
R754 VTAIL.n471 VTAIL.n419 3.49141
R755 VTAIL.n450 VTAIL.n431 3.49141
R756 VTAIL.n389 VTAIL.n337 3.49141
R757 VTAIL.n368 VTAIL.n349 3.49141
R758 VTAIL.n307 VTAIL.n255 3.49141
R759 VTAIL.n286 VTAIL.n267 3.49141
R760 VTAIL.n409 VTAIL.n327 3.4574
R761 VTAIL.n573 VTAIL.n491 3.4574
R762 VTAIL.n245 VTAIL.n163 3.4574
R763 VTAIL.n610 VTAIL.n609 2.71565
R764 VTAIL.n638 VTAIL.n637 2.71565
R765 VTAIL.n36 VTAIL.n35 2.71565
R766 VTAIL.n64 VTAIL.n63 2.71565
R767 VTAIL.n118 VTAIL.n117 2.71565
R768 VTAIL.n146 VTAIL.n145 2.71565
R769 VTAIL.n200 VTAIL.n199 2.71565
R770 VTAIL.n228 VTAIL.n227 2.71565
R771 VTAIL.n557 VTAIL.n556 2.71565
R772 VTAIL.n529 VTAIL.n528 2.71565
R773 VTAIL.n475 VTAIL.n474 2.71565
R774 VTAIL.n447 VTAIL.n446 2.71565
R775 VTAIL.n393 VTAIL.n392 2.71565
R776 VTAIL.n365 VTAIL.n364 2.71565
R777 VTAIL.n311 VTAIL.n310 2.71565
R778 VTAIL.n283 VTAIL.n282 2.71565
R779 VTAIL.n606 VTAIL.n596 1.93989
R780 VTAIL.n642 VTAIL.n580 1.93989
R781 VTAIL.n654 VTAIL.n574 1.93989
R782 VTAIL.n32 VTAIL.n22 1.93989
R783 VTAIL.n68 VTAIL.n6 1.93989
R784 VTAIL.n80 VTAIL.n0 1.93989
R785 VTAIL.n114 VTAIL.n104 1.93989
R786 VTAIL.n150 VTAIL.n88 1.93989
R787 VTAIL.n162 VTAIL.n82 1.93989
R788 VTAIL.n196 VTAIL.n186 1.93989
R789 VTAIL.n232 VTAIL.n170 1.93989
R790 VTAIL.n244 VTAIL.n164 1.93989
R791 VTAIL.n572 VTAIL.n492 1.93989
R792 VTAIL.n560 VTAIL.n498 1.93989
R793 VTAIL.n525 VTAIL.n515 1.93989
R794 VTAIL.n490 VTAIL.n410 1.93989
R795 VTAIL.n478 VTAIL.n416 1.93989
R796 VTAIL.n443 VTAIL.n433 1.93989
R797 VTAIL.n408 VTAIL.n328 1.93989
R798 VTAIL.n396 VTAIL.n334 1.93989
R799 VTAIL.n361 VTAIL.n351 1.93989
R800 VTAIL.n326 VTAIL.n246 1.93989
R801 VTAIL.n314 VTAIL.n252 1.93989
R802 VTAIL.n279 VTAIL.n269 1.93989
R803 VTAIL VTAIL.n81 1.78714
R804 VTAIL VTAIL.n655 1.67076
R805 VTAIL.n605 VTAIL.n598 1.16414
R806 VTAIL.n643 VTAIL.n578 1.16414
R807 VTAIL.n652 VTAIL.n651 1.16414
R808 VTAIL.n31 VTAIL.n24 1.16414
R809 VTAIL.n69 VTAIL.n4 1.16414
R810 VTAIL.n78 VTAIL.n77 1.16414
R811 VTAIL.n113 VTAIL.n106 1.16414
R812 VTAIL.n151 VTAIL.n86 1.16414
R813 VTAIL.n160 VTAIL.n159 1.16414
R814 VTAIL.n195 VTAIL.n188 1.16414
R815 VTAIL.n233 VTAIL.n168 1.16414
R816 VTAIL.n242 VTAIL.n241 1.16414
R817 VTAIL.n570 VTAIL.n569 1.16414
R818 VTAIL.n561 VTAIL.n496 1.16414
R819 VTAIL.n524 VTAIL.n517 1.16414
R820 VTAIL.n488 VTAIL.n487 1.16414
R821 VTAIL.n479 VTAIL.n414 1.16414
R822 VTAIL.n442 VTAIL.n435 1.16414
R823 VTAIL.n406 VTAIL.n405 1.16414
R824 VTAIL.n397 VTAIL.n332 1.16414
R825 VTAIL.n360 VTAIL.n353 1.16414
R826 VTAIL.n324 VTAIL.n323 1.16414
R827 VTAIL.n315 VTAIL.n250 1.16414
R828 VTAIL.n278 VTAIL.n271 1.16414
R829 VTAIL.n491 VTAIL.n409 0.470328
R830 VTAIL.n163 VTAIL.n81 0.470328
R831 VTAIL.n602 VTAIL.n601 0.388379
R832 VTAIL.n647 VTAIL.n646 0.388379
R833 VTAIL.n648 VTAIL.n576 0.388379
R834 VTAIL.n28 VTAIL.n27 0.388379
R835 VTAIL.n73 VTAIL.n72 0.388379
R836 VTAIL.n74 VTAIL.n2 0.388379
R837 VTAIL.n110 VTAIL.n109 0.388379
R838 VTAIL.n155 VTAIL.n154 0.388379
R839 VTAIL.n156 VTAIL.n84 0.388379
R840 VTAIL.n192 VTAIL.n191 0.388379
R841 VTAIL.n237 VTAIL.n236 0.388379
R842 VTAIL.n238 VTAIL.n166 0.388379
R843 VTAIL.n566 VTAIL.n494 0.388379
R844 VTAIL.n565 VTAIL.n564 0.388379
R845 VTAIL.n521 VTAIL.n520 0.388379
R846 VTAIL.n484 VTAIL.n412 0.388379
R847 VTAIL.n483 VTAIL.n482 0.388379
R848 VTAIL.n439 VTAIL.n438 0.388379
R849 VTAIL.n402 VTAIL.n330 0.388379
R850 VTAIL.n401 VTAIL.n400 0.388379
R851 VTAIL.n357 VTAIL.n356 0.388379
R852 VTAIL.n320 VTAIL.n248 0.388379
R853 VTAIL.n319 VTAIL.n318 0.388379
R854 VTAIL.n275 VTAIL.n274 0.388379
R855 VTAIL.n604 VTAIL.n603 0.155672
R856 VTAIL.n604 VTAIL.n595 0.155672
R857 VTAIL.n611 VTAIL.n595 0.155672
R858 VTAIL.n612 VTAIL.n611 0.155672
R859 VTAIL.n612 VTAIL.n591 0.155672
R860 VTAIL.n619 VTAIL.n591 0.155672
R861 VTAIL.n620 VTAIL.n619 0.155672
R862 VTAIL.n620 VTAIL.n587 0.155672
R863 VTAIL.n627 VTAIL.n587 0.155672
R864 VTAIL.n628 VTAIL.n627 0.155672
R865 VTAIL.n628 VTAIL.n583 0.155672
R866 VTAIL.n635 VTAIL.n583 0.155672
R867 VTAIL.n636 VTAIL.n635 0.155672
R868 VTAIL.n636 VTAIL.n579 0.155672
R869 VTAIL.n644 VTAIL.n579 0.155672
R870 VTAIL.n645 VTAIL.n644 0.155672
R871 VTAIL.n645 VTAIL.n575 0.155672
R872 VTAIL.n653 VTAIL.n575 0.155672
R873 VTAIL.n30 VTAIL.n29 0.155672
R874 VTAIL.n30 VTAIL.n21 0.155672
R875 VTAIL.n37 VTAIL.n21 0.155672
R876 VTAIL.n38 VTAIL.n37 0.155672
R877 VTAIL.n38 VTAIL.n17 0.155672
R878 VTAIL.n45 VTAIL.n17 0.155672
R879 VTAIL.n46 VTAIL.n45 0.155672
R880 VTAIL.n46 VTAIL.n13 0.155672
R881 VTAIL.n53 VTAIL.n13 0.155672
R882 VTAIL.n54 VTAIL.n53 0.155672
R883 VTAIL.n54 VTAIL.n9 0.155672
R884 VTAIL.n61 VTAIL.n9 0.155672
R885 VTAIL.n62 VTAIL.n61 0.155672
R886 VTAIL.n62 VTAIL.n5 0.155672
R887 VTAIL.n70 VTAIL.n5 0.155672
R888 VTAIL.n71 VTAIL.n70 0.155672
R889 VTAIL.n71 VTAIL.n1 0.155672
R890 VTAIL.n79 VTAIL.n1 0.155672
R891 VTAIL.n112 VTAIL.n111 0.155672
R892 VTAIL.n112 VTAIL.n103 0.155672
R893 VTAIL.n119 VTAIL.n103 0.155672
R894 VTAIL.n120 VTAIL.n119 0.155672
R895 VTAIL.n120 VTAIL.n99 0.155672
R896 VTAIL.n127 VTAIL.n99 0.155672
R897 VTAIL.n128 VTAIL.n127 0.155672
R898 VTAIL.n128 VTAIL.n95 0.155672
R899 VTAIL.n135 VTAIL.n95 0.155672
R900 VTAIL.n136 VTAIL.n135 0.155672
R901 VTAIL.n136 VTAIL.n91 0.155672
R902 VTAIL.n143 VTAIL.n91 0.155672
R903 VTAIL.n144 VTAIL.n143 0.155672
R904 VTAIL.n144 VTAIL.n87 0.155672
R905 VTAIL.n152 VTAIL.n87 0.155672
R906 VTAIL.n153 VTAIL.n152 0.155672
R907 VTAIL.n153 VTAIL.n83 0.155672
R908 VTAIL.n161 VTAIL.n83 0.155672
R909 VTAIL.n194 VTAIL.n193 0.155672
R910 VTAIL.n194 VTAIL.n185 0.155672
R911 VTAIL.n201 VTAIL.n185 0.155672
R912 VTAIL.n202 VTAIL.n201 0.155672
R913 VTAIL.n202 VTAIL.n181 0.155672
R914 VTAIL.n209 VTAIL.n181 0.155672
R915 VTAIL.n210 VTAIL.n209 0.155672
R916 VTAIL.n210 VTAIL.n177 0.155672
R917 VTAIL.n217 VTAIL.n177 0.155672
R918 VTAIL.n218 VTAIL.n217 0.155672
R919 VTAIL.n218 VTAIL.n173 0.155672
R920 VTAIL.n225 VTAIL.n173 0.155672
R921 VTAIL.n226 VTAIL.n225 0.155672
R922 VTAIL.n226 VTAIL.n169 0.155672
R923 VTAIL.n234 VTAIL.n169 0.155672
R924 VTAIL.n235 VTAIL.n234 0.155672
R925 VTAIL.n235 VTAIL.n165 0.155672
R926 VTAIL.n243 VTAIL.n165 0.155672
R927 VTAIL.n571 VTAIL.n493 0.155672
R928 VTAIL.n563 VTAIL.n493 0.155672
R929 VTAIL.n563 VTAIL.n562 0.155672
R930 VTAIL.n562 VTAIL.n497 0.155672
R931 VTAIL.n555 VTAIL.n497 0.155672
R932 VTAIL.n555 VTAIL.n554 0.155672
R933 VTAIL.n554 VTAIL.n502 0.155672
R934 VTAIL.n547 VTAIL.n502 0.155672
R935 VTAIL.n547 VTAIL.n546 0.155672
R936 VTAIL.n546 VTAIL.n506 0.155672
R937 VTAIL.n539 VTAIL.n506 0.155672
R938 VTAIL.n539 VTAIL.n538 0.155672
R939 VTAIL.n538 VTAIL.n510 0.155672
R940 VTAIL.n531 VTAIL.n510 0.155672
R941 VTAIL.n531 VTAIL.n530 0.155672
R942 VTAIL.n530 VTAIL.n514 0.155672
R943 VTAIL.n523 VTAIL.n514 0.155672
R944 VTAIL.n523 VTAIL.n522 0.155672
R945 VTAIL.n489 VTAIL.n411 0.155672
R946 VTAIL.n481 VTAIL.n411 0.155672
R947 VTAIL.n481 VTAIL.n480 0.155672
R948 VTAIL.n480 VTAIL.n415 0.155672
R949 VTAIL.n473 VTAIL.n415 0.155672
R950 VTAIL.n473 VTAIL.n472 0.155672
R951 VTAIL.n472 VTAIL.n420 0.155672
R952 VTAIL.n465 VTAIL.n420 0.155672
R953 VTAIL.n465 VTAIL.n464 0.155672
R954 VTAIL.n464 VTAIL.n424 0.155672
R955 VTAIL.n457 VTAIL.n424 0.155672
R956 VTAIL.n457 VTAIL.n456 0.155672
R957 VTAIL.n456 VTAIL.n428 0.155672
R958 VTAIL.n449 VTAIL.n428 0.155672
R959 VTAIL.n449 VTAIL.n448 0.155672
R960 VTAIL.n448 VTAIL.n432 0.155672
R961 VTAIL.n441 VTAIL.n432 0.155672
R962 VTAIL.n441 VTAIL.n440 0.155672
R963 VTAIL.n407 VTAIL.n329 0.155672
R964 VTAIL.n399 VTAIL.n329 0.155672
R965 VTAIL.n399 VTAIL.n398 0.155672
R966 VTAIL.n398 VTAIL.n333 0.155672
R967 VTAIL.n391 VTAIL.n333 0.155672
R968 VTAIL.n391 VTAIL.n390 0.155672
R969 VTAIL.n390 VTAIL.n338 0.155672
R970 VTAIL.n383 VTAIL.n338 0.155672
R971 VTAIL.n383 VTAIL.n382 0.155672
R972 VTAIL.n382 VTAIL.n342 0.155672
R973 VTAIL.n375 VTAIL.n342 0.155672
R974 VTAIL.n375 VTAIL.n374 0.155672
R975 VTAIL.n374 VTAIL.n346 0.155672
R976 VTAIL.n367 VTAIL.n346 0.155672
R977 VTAIL.n367 VTAIL.n366 0.155672
R978 VTAIL.n366 VTAIL.n350 0.155672
R979 VTAIL.n359 VTAIL.n350 0.155672
R980 VTAIL.n359 VTAIL.n358 0.155672
R981 VTAIL.n325 VTAIL.n247 0.155672
R982 VTAIL.n317 VTAIL.n247 0.155672
R983 VTAIL.n317 VTAIL.n316 0.155672
R984 VTAIL.n316 VTAIL.n251 0.155672
R985 VTAIL.n309 VTAIL.n251 0.155672
R986 VTAIL.n309 VTAIL.n308 0.155672
R987 VTAIL.n308 VTAIL.n256 0.155672
R988 VTAIL.n301 VTAIL.n256 0.155672
R989 VTAIL.n301 VTAIL.n300 0.155672
R990 VTAIL.n300 VTAIL.n260 0.155672
R991 VTAIL.n293 VTAIL.n260 0.155672
R992 VTAIL.n293 VTAIL.n292 0.155672
R993 VTAIL.n292 VTAIL.n264 0.155672
R994 VTAIL.n285 VTAIL.n264 0.155672
R995 VTAIL.n285 VTAIL.n284 0.155672
R996 VTAIL.n284 VTAIL.n268 0.155672
R997 VTAIL.n277 VTAIL.n268 0.155672
R998 VTAIL.n277 VTAIL.n276 0.155672
R999 VDD2.n2 VDD2.n0 111.678
R1000 VDD2.n2 VDD2.n1 64.7997
R1001 VDD2.n1 VDD2.t1 1.33473
R1002 VDD2.n1 VDD2.t0 1.33473
R1003 VDD2.n0 VDD2.t2 1.33473
R1004 VDD2.n0 VDD2.t3 1.33473
R1005 VDD2 VDD2.n2 0.0586897
R1006 B.n905 B.n904 585
R1007 B.n355 B.n135 585
R1008 B.n354 B.n353 585
R1009 B.n352 B.n351 585
R1010 B.n350 B.n349 585
R1011 B.n348 B.n347 585
R1012 B.n346 B.n345 585
R1013 B.n344 B.n343 585
R1014 B.n342 B.n341 585
R1015 B.n340 B.n339 585
R1016 B.n338 B.n337 585
R1017 B.n336 B.n335 585
R1018 B.n334 B.n333 585
R1019 B.n332 B.n331 585
R1020 B.n330 B.n329 585
R1021 B.n328 B.n327 585
R1022 B.n326 B.n325 585
R1023 B.n324 B.n323 585
R1024 B.n322 B.n321 585
R1025 B.n320 B.n319 585
R1026 B.n318 B.n317 585
R1027 B.n316 B.n315 585
R1028 B.n314 B.n313 585
R1029 B.n312 B.n311 585
R1030 B.n310 B.n309 585
R1031 B.n308 B.n307 585
R1032 B.n306 B.n305 585
R1033 B.n304 B.n303 585
R1034 B.n302 B.n301 585
R1035 B.n300 B.n299 585
R1036 B.n298 B.n297 585
R1037 B.n296 B.n295 585
R1038 B.n294 B.n293 585
R1039 B.n292 B.n291 585
R1040 B.n290 B.n289 585
R1041 B.n288 B.n287 585
R1042 B.n286 B.n285 585
R1043 B.n284 B.n283 585
R1044 B.n282 B.n281 585
R1045 B.n280 B.n279 585
R1046 B.n278 B.n277 585
R1047 B.n276 B.n275 585
R1048 B.n274 B.n273 585
R1049 B.n272 B.n271 585
R1050 B.n270 B.n269 585
R1051 B.n268 B.n267 585
R1052 B.n266 B.n265 585
R1053 B.n264 B.n263 585
R1054 B.n262 B.n261 585
R1055 B.n260 B.n259 585
R1056 B.n258 B.n257 585
R1057 B.n256 B.n255 585
R1058 B.n254 B.n253 585
R1059 B.n252 B.n251 585
R1060 B.n250 B.n249 585
R1061 B.n248 B.n247 585
R1062 B.n246 B.n245 585
R1063 B.n244 B.n243 585
R1064 B.n242 B.n241 585
R1065 B.n240 B.n239 585
R1066 B.n238 B.n237 585
R1067 B.n236 B.n235 585
R1068 B.n234 B.n233 585
R1069 B.n232 B.n231 585
R1070 B.n230 B.n229 585
R1071 B.n228 B.n227 585
R1072 B.n226 B.n225 585
R1073 B.n224 B.n223 585
R1074 B.n222 B.n221 585
R1075 B.n220 B.n219 585
R1076 B.n218 B.n217 585
R1077 B.n216 B.n215 585
R1078 B.n214 B.n213 585
R1079 B.n212 B.n211 585
R1080 B.n210 B.n209 585
R1081 B.n208 B.n207 585
R1082 B.n206 B.n205 585
R1083 B.n204 B.n203 585
R1084 B.n202 B.n201 585
R1085 B.n200 B.n199 585
R1086 B.n198 B.n197 585
R1087 B.n196 B.n195 585
R1088 B.n194 B.n193 585
R1089 B.n192 B.n191 585
R1090 B.n190 B.n189 585
R1091 B.n188 B.n187 585
R1092 B.n186 B.n185 585
R1093 B.n184 B.n183 585
R1094 B.n182 B.n181 585
R1095 B.n180 B.n179 585
R1096 B.n178 B.n177 585
R1097 B.n176 B.n175 585
R1098 B.n174 B.n173 585
R1099 B.n172 B.n171 585
R1100 B.n170 B.n169 585
R1101 B.n168 B.n167 585
R1102 B.n166 B.n165 585
R1103 B.n164 B.n163 585
R1104 B.n162 B.n161 585
R1105 B.n160 B.n159 585
R1106 B.n158 B.n157 585
R1107 B.n156 B.n155 585
R1108 B.n154 B.n153 585
R1109 B.n152 B.n151 585
R1110 B.n150 B.n149 585
R1111 B.n148 B.n147 585
R1112 B.n146 B.n145 585
R1113 B.n144 B.n143 585
R1114 B.n81 B.n80 585
R1115 B.n910 B.n909 585
R1116 B.n903 B.n136 585
R1117 B.n136 B.n78 585
R1118 B.n902 B.n77 585
R1119 B.n914 B.n77 585
R1120 B.n901 B.n76 585
R1121 B.n915 B.n76 585
R1122 B.n900 B.n75 585
R1123 B.n916 B.n75 585
R1124 B.n899 B.n898 585
R1125 B.n898 B.n71 585
R1126 B.n897 B.n70 585
R1127 B.n922 B.n70 585
R1128 B.n896 B.n69 585
R1129 B.n923 B.n69 585
R1130 B.n895 B.n68 585
R1131 B.n924 B.n68 585
R1132 B.n894 B.n893 585
R1133 B.n893 B.n64 585
R1134 B.n892 B.n63 585
R1135 B.n930 B.n63 585
R1136 B.n891 B.n62 585
R1137 B.n931 B.n62 585
R1138 B.n890 B.n61 585
R1139 B.n932 B.n61 585
R1140 B.n889 B.n888 585
R1141 B.n888 B.n57 585
R1142 B.n887 B.n56 585
R1143 B.n938 B.n56 585
R1144 B.n886 B.n55 585
R1145 B.n939 B.n55 585
R1146 B.n885 B.n54 585
R1147 B.n940 B.n54 585
R1148 B.n884 B.n883 585
R1149 B.n883 B.n50 585
R1150 B.n882 B.n49 585
R1151 B.n946 B.n49 585
R1152 B.n881 B.n48 585
R1153 B.n947 B.n48 585
R1154 B.n880 B.n47 585
R1155 B.n948 B.n47 585
R1156 B.n879 B.n878 585
R1157 B.n878 B.n43 585
R1158 B.n877 B.n42 585
R1159 B.n954 B.n42 585
R1160 B.n876 B.n41 585
R1161 B.n955 B.n41 585
R1162 B.n875 B.n40 585
R1163 B.n956 B.n40 585
R1164 B.n874 B.n873 585
R1165 B.n873 B.n39 585
R1166 B.n872 B.n35 585
R1167 B.n962 B.n35 585
R1168 B.n871 B.n34 585
R1169 B.n963 B.n34 585
R1170 B.n870 B.n33 585
R1171 B.n964 B.n33 585
R1172 B.n869 B.n868 585
R1173 B.n868 B.n29 585
R1174 B.n867 B.n28 585
R1175 B.n970 B.n28 585
R1176 B.n866 B.n27 585
R1177 B.n971 B.n27 585
R1178 B.n865 B.n26 585
R1179 B.n972 B.n26 585
R1180 B.n864 B.n863 585
R1181 B.n863 B.n22 585
R1182 B.n862 B.n21 585
R1183 B.n978 B.n21 585
R1184 B.n861 B.n20 585
R1185 B.n979 B.n20 585
R1186 B.n860 B.n19 585
R1187 B.n980 B.n19 585
R1188 B.n859 B.n858 585
R1189 B.n858 B.t2 585
R1190 B.n857 B.n15 585
R1191 B.n986 B.n15 585
R1192 B.n856 B.n14 585
R1193 B.n987 B.n14 585
R1194 B.n855 B.n13 585
R1195 B.n988 B.n13 585
R1196 B.n854 B.n853 585
R1197 B.n853 B.n12 585
R1198 B.n852 B.n851 585
R1199 B.n852 B.n8 585
R1200 B.n850 B.n7 585
R1201 B.n995 B.n7 585
R1202 B.n849 B.n6 585
R1203 B.n996 B.n6 585
R1204 B.n848 B.n5 585
R1205 B.n997 B.n5 585
R1206 B.n847 B.n846 585
R1207 B.n846 B.n4 585
R1208 B.n845 B.n356 585
R1209 B.n845 B.n844 585
R1210 B.n835 B.n357 585
R1211 B.n358 B.n357 585
R1212 B.n837 B.n836 585
R1213 B.n838 B.n837 585
R1214 B.n834 B.n363 585
R1215 B.n363 B.n362 585
R1216 B.n833 B.n832 585
R1217 B.n832 B.n831 585
R1218 B.n365 B.n364 585
R1219 B.t3 B.n365 585
R1220 B.n824 B.n823 585
R1221 B.n825 B.n824 585
R1222 B.n822 B.n370 585
R1223 B.n370 B.n369 585
R1224 B.n821 B.n820 585
R1225 B.n820 B.n819 585
R1226 B.n372 B.n371 585
R1227 B.n373 B.n372 585
R1228 B.n812 B.n811 585
R1229 B.n813 B.n812 585
R1230 B.n810 B.n378 585
R1231 B.n378 B.n377 585
R1232 B.n809 B.n808 585
R1233 B.n808 B.n807 585
R1234 B.n380 B.n379 585
R1235 B.n381 B.n380 585
R1236 B.n800 B.n799 585
R1237 B.n801 B.n800 585
R1238 B.n798 B.n386 585
R1239 B.n386 B.n385 585
R1240 B.n797 B.n796 585
R1241 B.n796 B.n795 585
R1242 B.n388 B.n387 585
R1243 B.n788 B.n388 585
R1244 B.n787 B.n786 585
R1245 B.n789 B.n787 585
R1246 B.n785 B.n393 585
R1247 B.n393 B.n392 585
R1248 B.n784 B.n783 585
R1249 B.n783 B.n782 585
R1250 B.n395 B.n394 585
R1251 B.n396 B.n395 585
R1252 B.n775 B.n774 585
R1253 B.n776 B.n775 585
R1254 B.n773 B.n401 585
R1255 B.n401 B.n400 585
R1256 B.n772 B.n771 585
R1257 B.n771 B.n770 585
R1258 B.n403 B.n402 585
R1259 B.n404 B.n403 585
R1260 B.n763 B.n762 585
R1261 B.n764 B.n763 585
R1262 B.n761 B.n409 585
R1263 B.n409 B.n408 585
R1264 B.n760 B.n759 585
R1265 B.n759 B.n758 585
R1266 B.n411 B.n410 585
R1267 B.n412 B.n411 585
R1268 B.n751 B.n750 585
R1269 B.n752 B.n751 585
R1270 B.n749 B.n417 585
R1271 B.n417 B.n416 585
R1272 B.n748 B.n747 585
R1273 B.n747 B.n746 585
R1274 B.n419 B.n418 585
R1275 B.n420 B.n419 585
R1276 B.n739 B.n738 585
R1277 B.n740 B.n739 585
R1278 B.n737 B.n425 585
R1279 B.n425 B.n424 585
R1280 B.n736 B.n735 585
R1281 B.n735 B.n734 585
R1282 B.n427 B.n426 585
R1283 B.n428 B.n427 585
R1284 B.n727 B.n726 585
R1285 B.n728 B.n727 585
R1286 B.n725 B.n433 585
R1287 B.n433 B.n432 585
R1288 B.n724 B.n723 585
R1289 B.n723 B.n722 585
R1290 B.n435 B.n434 585
R1291 B.n436 B.n435 585
R1292 B.n718 B.n717 585
R1293 B.n439 B.n438 585
R1294 B.n714 B.n713 585
R1295 B.n715 B.n714 585
R1296 B.n712 B.n494 585
R1297 B.n711 B.n710 585
R1298 B.n709 B.n708 585
R1299 B.n707 B.n706 585
R1300 B.n705 B.n704 585
R1301 B.n703 B.n702 585
R1302 B.n701 B.n700 585
R1303 B.n699 B.n698 585
R1304 B.n697 B.n696 585
R1305 B.n695 B.n694 585
R1306 B.n693 B.n692 585
R1307 B.n691 B.n690 585
R1308 B.n689 B.n688 585
R1309 B.n687 B.n686 585
R1310 B.n685 B.n684 585
R1311 B.n683 B.n682 585
R1312 B.n681 B.n680 585
R1313 B.n679 B.n678 585
R1314 B.n677 B.n676 585
R1315 B.n675 B.n674 585
R1316 B.n673 B.n672 585
R1317 B.n671 B.n670 585
R1318 B.n669 B.n668 585
R1319 B.n667 B.n666 585
R1320 B.n665 B.n664 585
R1321 B.n663 B.n662 585
R1322 B.n661 B.n660 585
R1323 B.n659 B.n658 585
R1324 B.n657 B.n656 585
R1325 B.n655 B.n654 585
R1326 B.n653 B.n652 585
R1327 B.n651 B.n650 585
R1328 B.n649 B.n648 585
R1329 B.n647 B.n646 585
R1330 B.n645 B.n644 585
R1331 B.n643 B.n642 585
R1332 B.n641 B.n640 585
R1333 B.n639 B.n638 585
R1334 B.n637 B.n636 585
R1335 B.n635 B.n634 585
R1336 B.n633 B.n632 585
R1337 B.n631 B.n630 585
R1338 B.n629 B.n628 585
R1339 B.n627 B.n626 585
R1340 B.n625 B.n624 585
R1341 B.n623 B.n622 585
R1342 B.n621 B.n620 585
R1343 B.n618 B.n617 585
R1344 B.n616 B.n615 585
R1345 B.n614 B.n613 585
R1346 B.n612 B.n611 585
R1347 B.n610 B.n609 585
R1348 B.n608 B.n607 585
R1349 B.n606 B.n605 585
R1350 B.n604 B.n603 585
R1351 B.n602 B.n601 585
R1352 B.n600 B.n599 585
R1353 B.n597 B.n596 585
R1354 B.n595 B.n594 585
R1355 B.n593 B.n592 585
R1356 B.n591 B.n590 585
R1357 B.n589 B.n588 585
R1358 B.n587 B.n586 585
R1359 B.n585 B.n584 585
R1360 B.n583 B.n582 585
R1361 B.n581 B.n580 585
R1362 B.n579 B.n578 585
R1363 B.n577 B.n576 585
R1364 B.n575 B.n574 585
R1365 B.n573 B.n572 585
R1366 B.n571 B.n570 585
R1367 B.n569 B.n568 585
R1368 B.n567 B.n566 585
R1369 B.n565 B.n564 585
R1370 B.n563 B.n562 585
R1371 B.n561 B.n560 585
R1372 B.n559 B.n558 585
R1373 B.n557 B.n556 585
R1374 B.n555 B.n554 585
R1375 B.n553 B.n552 585
R1376 B.n551 B.n550 585
R1377 B.n549 B.n548 585
R1378 B.n547 B.n546 585
R1379 B.n545 B.n544 585
R1380 B.n543 B.n542 585
R1381 B.n541 B.n540 585
R1382 B.n539 B.n538 585
R1383 B.n537 B.n536 585
R1384 B.n535 B.n534 585
R1385 B.n533 B.n532 585
R1386 B.n531 B.n530 585
R1387 B.n529 B.n528 585
R1388 B.n527 B.n526 585
R1389 B.n525 B.n524 585
R1390 B.n523 B.n522 585
R1391 B.n521 B.n520 585
R1392 B.n519 B.n518 585
R1393 B.n517 B.n516 585
R1394 B.n515 B.n514 585
R1395 B.n513 B.n512 585
R1396 B.n511 B.n510 585
R1397 B.n509 B.n508 585
R1398 B.n507 B.n506 585
R1399 B.n505 B.n504 585
R1400 B.n503 B.n502 585
R1401 B.n501 B.n500 585
R1402 B.n499 B.n493 585
R1403 B.n715 B.n493 585
R1404 B.n719 B.n437 585
R1405 B.n437 B.n436 585
R1406 B.n721 B.n720 585
R1407 B.n722 B.n721 585
R1408 B.n431 B.n430 585
R1409 B.n432 B.n431 585
R1410 B.n730 B.n729 585
R1411 B.n729 B.n728 585
R1412 B.n731 B.n429 585
R1413 B.n429 B.n428 585
R1414 B.n733 B.n732 585
R1415 B.n734 B.n733 585
R1416 B.n423 B.n422 585
R1417 B.n424 B.n423 585
R1418 B.n742 B.n741 585
R1419 B.n741 B.n740 585
R1420 B.n743 B.n421 585
R1421 B.n421 B.n420 585
R1422 B.n745 B.n744 585
R1423 B.n746 B.n745 585
R1424 B.n415 B.n414 585
R1425 B.n416 B.n415 585
R1426 B.n754 B.n753 585
R1427 B.n753 B.n752 585
R1428 B.n755 B.n413 585
R1429 B.n413 B.n412 585
R1430 B.n757 B.n756 585
R1431 B.n758 B.n757 585
R1432 B.n407 B.n406 585
R1433 B.n408 B.n407 585
R1434 B.n766 B.n765 585
R1435 B.n765 B.n764 585
R1436 B.n767 B.n405 585
R1437 B.n405 B.n404 585
R1438 B.n769 B.n768 585
R1439 B.n770 B.n769 585
R1440 B.n399 B.n398 585
R1441 B.n400 B.n399 585
R1442 B.n778 B.n777 585
R1443 B.n777 B.n776 585
R1444 B.n779 B.n397 585
R1445 B.n397 B.n396 585
R1446 B.n781 B.n780 585
R1447 B.n782 B.n781 585
R1448 B.n391 B.n390 585
R1449 B.n392 B.n391 585
R1450 B.n791 B.n790 585
R1451 B.n790 B.n789 585
R1452 B.n792 B.n389 585
R1453 B.n788 B.n389 585
R1454 B.n794 B.n793 585
R1455 B.n795 B.n794 585
R1456 B.n384 B.n383 585
R1457 B.n385 B.n384 585
R1458 B.n803 B.n802 585
R1459 B.n802 B.n801 585
R1460 B.n804 B.n382 585
R1461 B.n382 B.n381 585
R1462 B.n806 B.n805 585
R1463 B.n807 B.n806 585
R1464 B.n376 B.n375 585
R1465 B.n377 B.n376 585
R1466 B.n815 B.n814 585
R1467 B.n814 B.n813 585
R1468 B.n816 B.n374 585
R1469 B.n374 B.n373 585
R1470 B.n818 B.n817 585
R1471 B.n819 B.n818 585
R1472 B.n368 B.n367 585
R1473 B.n369 B.n368 585
R1474 B.n827 B.n826 585
R1475 B.n826 B.n825 585
R1476 B.n828 B.n366 585
R1477 B.n366 B.t3 585
R1478 B.n830 B.n829 585
R1479 B.n831 B.n830 585
R1480 B.n361 B.n360 585
R1481 B.n362 B.n361 585
R1482 B.n840 B.n839 585
R1483 B.n839 B.n838 585
R1484 B.n841 B.n359 585
R1485 B.n359 B.n358 585
R1486 B.n843 B.n842 585
R1487 B.n844 B.n843 585
R1488 B.n3 B.n0 585
R1489 B.n4 B.n3 585
R1490 B.n994 B.n1 585
R1491 B.n995 B.n994 585
R1492 B.n993 B.n992 585
R1493 B.n993 B.n8 585
R1494 B.n991 B.n9 585
R1495 B.n12 B.n9 585
R1496 B.n990 B.n989 585
R1497 B.n989 B.n988 585
R1498 B.n11 B.n10 585
R1499 B.n987 B.n11 585
R1500 B.n985 B.n984 585
R1501 B.n986 B.n985 585
R1502 B.n983 B.n16 585
R1503 B.n16 B.t2 585
R1504 B.n982 B.n981 585
R1505 B.n981 B.n980 585
R1506 B.n18 B.n17 585
R1507 B.n979 B.n18 585
R1508 B.n977 B.n976 585
R1509 B.n978 B.n977 585
R1510 B.n975 B.n23 585
R1511 B.n23 B.n22 585
R1512 B.n974 B.n973 585
R1513 B.n973 B.n972 585
R1514 B.n25 B.n24 585
R1515 B.n971 B.n25 585
R1516 B.n969 B.n968 585
R1517 B.n970 B.n969 585
R1518 B.n967 B.n30 585
R1519 B.n30 B.n29 585
R1520 B.n966 B.n965 585
R1521 B.n965 B.n964 585
R1522 B.n32 B.n31 585
R1523 B.n963 B.n32 585
R1524 B.n961 B.n960 585
R1525 B.n962 B.n961 585
R1526 B.n959 B.n36 585
R1527 B.n39 B.n36 585
R1528 B.n958 B.n957 585
R1529 B.n957 B.n956 585
R1530 B.n38 B.n37 585
R1531 B.n955 B.n38 585
R1532 B.n953 B.n952 585
R1533 B.n954 B.n953 585
R1534 B.n951 B.n44 585
R1535 B.n44 B.n43 585
R1536 B.n950 B.n949 585
R1537 B.n949 B.n948 585
R1538 B.n46 B.n45 585
R1539 B.n947 B.n46 585
R1540 B.n945 B.n944 585
R1541 B.n946 B.n945 585
R1542 B.n943 B.n51 585
R1543 B.n51 B.n50 585
R1544 B.n942 B.n941 585
R1545 B.n941 B.n940 585
R1546 B.n53 B.n52 585
R1547 B.n939 B.n53 585
R1548 B.n937 B.n936 585
R1549 B.n938 B.n937 585
R1550 B.n935 B.n58 585
R1551 B.n58 B.n57 585
R1552 B.n934 B.n933 585
R1553 B.n933 B.n932 585
R1554 B.n60 B.n59 585
R1555 B.n931 B.n60 585
R1556 B.n929 B.n928 585
R1557 B.n930 B.n929 585
R1558 B.n927 B.n65 585
R1559 B.n65 B.n64 585
R1560 B.n926 B.n925 585
R1561 B.n925 B.n924 585
R1562 B.n67 B.n66 585
R1563 B.n923 B.n67 585
R1564 B.n921 B.n920 585
R1565 B.n922 B.n921 585
R1566 B.n919 B.n72 585
R1567 B.n72 B.n71 585
R1568 B.n918 B.n917 585
R1569 B.n917 B.n916 585
R1570 B.n74 B.n73 585
R1571 B.n915 B.n74 585
R1572 B.n913 B.n912 585
R1573 B.n914 B.n913 585
R1574 B.n911 B.n79 585
R1575 B.n79 B.n78 585
R1576 B.n998 B.n997 585
R1577 B.n996 B.n2 585
R1578 B.n909 B.n79 458.866
R1579 B.n905 B.n136 458.866
R1580 B.n493 B.n435 458.866
R1581 B.n717 B.n437 458.866
R1582 B.n140 B.t6 408.954
R1583 B.n137 B.t9 408.954
R1584 B.n497 B.t14 408.954
R1585 B.n495 B.t17 408.954
R1586 B.n138 B.t10 331.185
R1587 B.n498 B.t13 331.185
R1588 B.n141 B.t7 331.185
R1589 B.n496 B.t16 331.185
R1590 B.n140 B.t4 306.435
R1591 B.n137 B.t8 306.435
R1592 B.n497 B.t11 306.435
R1593 B.n495 B.t15 306.435
R1594 B.n907 B.n906 256.663
R1595 B.n907 B.n134 256.663
R1596 B.n907 B.n133 256.663
R1597 B.n907 B.n132 256.663
R1598 B.n907 B.n131 256.663
R1599 B.n907 B.n130 256.663
R1600 B.n907 B.n129 256.663
R1601 B.n907 B.n128 256.663
R1602 B.n907 B.n127 256.663
R1603 B.n907 B.n126 256.663
R1604 B.n907 B.n125 256.663
R1605 B.n907 B.n124 256.663
R1606 B.n907 B.n123 256.663
R1607 B.n907 B.n122 256.663
R1608 B.n907 B.n121 256.663
R1609 B.n907 B.n120 256.663
R1610 B.n907 B.n119 256.663
R1611 B.n907 B.n118 256.663
R1612 B.n907 B.n117 256.663
R1613 B.n907 B.n116 256.663
R1614 B.n907 B.n115 256.663
R1615 B.n907 B.n114 256.663
R1616 B.n907 B.n113 256.663
R1617 B.n907 B.n112 256.663
R1618 B.n907 B.n111 256.663
R1619 B.n907 B.n110 256.663
R1620 B.n907 B.n109 256.663
R1621 B.n907 B.n108 256.663
R1622 B.n907 B.n107 256.663
R1623 B.n907 B.n106 256.663
R1624 B.n907 B.n105 256.663
R1625 B.n907 B.n104 256.663
R1626 B.n907 B.n103 256.663
R1627 B.n907 B.n102 256.663
R1628 B.n907 B.n101 256.663
R1629 B.n907 B.n100 256.663
R1630 B.n907 B.n99 256.663
R1631 B.n907 B.n98 256.663
R1632 B.n907 B.n97 256.663
R1633 B.n907 B.n96 256.663
R1634 B.n907 B.n95 256.663
R1635 B.n907 B.n94 256.663
R1636 B.n907 B.n93 256.663
R1637 B.n907 B.n92 256.663
R1638 B.n907 B.n91 256.663
R1639 B.n907 B.n90 256.663
R1640 B.n907 B.n89 256.663
R1641 B.n907 B.n88 256.663
R1642 B.n907 B.n87 256.663
R1643 B.n907 B.n86 256.663
R1644 B.n907 B.n85 256.663
R1645 B.n907 B.n84 256.663
R1646 B.n907 B.n83 256.663
R1647 B.n907 B.n82 256.663
R1648 B.n908 B.n907 256.663
R1649 B.n716 B.n715 256.663
R1650 B.n715 B.n440 256.663
R1651 B.n715 B.n441 256.663
R1652 B.n715 B.n442 256.663
R1653 B.n715 B.n443 256.663
R1654 B.n715 B.n444 256.663
R1655 B.n715 B.n445 256.663
R1656 B.n715 B.n446 256.663
R1657 B.n715 B.n447 256.663
R1658 B.n715 B.n448 256.663
R1659 B.n715 B.n449 256.663
R1660 B.n715 B.n450 256.663
R1661 B.n715 B.n451 256.663
R1662 B.n715 B.n452 256.663
R1663 B.n715 B.n453 256.663
R1664 B.n715 B.n454 256.663
R1665 B.n715 B.n455 256.663
R1666 B.n715 B.n456 256.663
R1667 B.n715 B.n457 256.663
R1668 B.n715 B.n458 256.663
R1669 B.n715 B.n459 256.663
R1670 B.n715 B.n460 256.663
R1671 B.n715 B.n461 256.663
R1672 B.n715 B.n462 256.663
R1673 B.n715 B.n463 256.663
R1674 B.n715 B.n464 256.663
R1675 B.n715 B.n465 256.663
R1676 B.n715 B.n466 256.663
R1677 B.n715 B.n467 256.663
R1678 B.n715 B.n468 256.663
R1679 B.n715 B.n469 256.663
R1680 B.n715 B.n470 256.663
R1681 B.n715 B.n471 256.663
R1682 B.n715 B.n472 256.663
R1683 B.n715 B.n473 256.663
R1684 B.n715 B.n474 256.663
R1685 B.n715 B.n475 256.663
R1686 B.n715 B.n476 256.663
R1687 B.n715 B.n477 256.663
R1688 B.n715 B.n478 256.663
R1689 B.n715 B.n479 256.663
R1690 B.n715 B.n480 256.663
R1691 B.n715 B.n481 256.663
R1692 B.n715 B.n482 256.663
R1693 B.n715 B.n483 256.663
R1694 B.n715 B.n484 256.663
R1695 B.n715 B.n485 256.663
R1696 B.n715 B.n486 256.663
R1697 B.n715 B.n487 256.663
R1698 B.n715 B.n488 256.663
R1699 B.n715 B.n489 256.663
R1700 B.n715 B.n490 256.663
R1701 B.n715 B.n491 256.663
R1702 B.n715 B.n492 256.663
R1703 B.n1000 B.n999 256.663
R1704 B.n143 B.n81 163.367
R1705 B.n147 B.n146 163.367
R1706 B.n151 B.n150 163.367
R1707 B.n155 B.n154 163.367
R1708 B.n159 B.n158 163.367
R1709 B.n163 B.n162 163.367
R1710 B.n167 B.n166 163.367
R1711 B.n171 B.n170 163.367
R1712 B.n175 B.n174 163.367
R1713 B.n179 B.n178 163.367
R1714 B.n183 B.n182 163.367
R1715 B.n187 B.n186 163.367
R1716 B.n191 B.n190 163.367
R1717 B.n195 B.n194 163.367
R1718 B.n199 B.n198 163.367
R1719 B.n203 B.n202 163.367
R1720 B.n207 B.n206 163.367
R1721 B.n211 B.n210 163.367
R1722 B.n215 B.n214 163.367
R1723 B.n219 B.n218 163.367
R1724 B.n223 B.n222 163.367
R1725 B.n227 B.n226 163.367
R1726 B.n231 B.n230 163.367
R1727 B.n235 B.n234 163.367
R1728 B.n239 B.n238 163.367
R1729 B.n243 B.n242 163.367
R1730 B.n247 B.n246 163.367
R1731 B.n251 B.n250 163.367
R1732 B.n255 B.n254 163.367
R1733 B.n259 B.n258 163.367
R1734 B.n263 B.n262 163.367
R1735 B.n267 B.n266 163.367
R1736 B.n271 B.n270 163.367
R1737 B.n275 B.n274 163.367
R1738 B.n279 B.n278 163.367
R1739 B.n283 B.n282 163.367
R1740 B.n287 B.n286 163.367
R1741 B.n291 B.n290 163.367
R1742 B.n295 B.n294 163.367
R1743 B.n299 B.n298 163.367
R1744 B.n303 B.n302 163.367
R1745 B.n307 B.n306 163.367
R1746 B.n311 B.n310 163.367
R1747 B.n315 B.n314 163.367
R1748 B.n319 B.n318 163.367
R1749 B.n323 B.n322 163.367
R1750 B.n327 B.n326 163.367
R1751 B.n331 B.n330 163.367
R1752 B.n335 B.n334 163.367
R1753 B.n339 B.n338 163.367
R1754 B.n343 B.n342 163.367
R1755 B.n347 B.n346 163.367
R1756 B.n351 B.n350 163.367
R1757 B.n353 B.n135 163.367
R1758 B.n723 B.n435 163.367
R1759 B.n723 B.n433 163.367
R1760 B.n727 B.n433 163.367
R1761 B.n727 B.n427 163.367
R1762 B.n735 B.n427 163.367
R1763 B.n735 B.n425 163.367
R1764 B.n739 B.n425 163.367
R1765 B.n739 B.n419 163.367
R1766 B.n747 B.n419 163.367
R1767 B.n747 B.n417 163.367
R1768 B.n751 B.n417 163.367
R1769 B.n751 B.n411 163.367
R1770 B.n759 B.n411 163.367
R1771 B.n759 B.n409 163.367
R1772 B.n763 B.n409 163.367
R1773 B.n763 B.n403 163.367
R1774 B.n771 B.n403 163.367
R1775 B.n771 B.n401 163.367
R1776 B.n775 B.n401 163.367
R1777 B.n775 B.n395 163.367
R1778 B.n783 B.n395 163.367
R1779 B.n783 B.n393 163.367
R1780 B.n787 B.n393 163.367
R1781 B.n787 B.n388 163.367
R1782 B.n796 B.n388 163.367
R1783 B.n796 B.n386 163.367
R1784 B.n800 B.n386 163.367
R1785 B.n800 B.n380 163.367
R1786 B.n808 B.n380 163.367
R1787 B.n808 B.n378 163.367
R1788 B.n812 B.n378 163.367
R1789 B.n812 B.n372 163.367
R1790 B.n820 B.n372 163.367
R1791 B.n820 B.n370 163.367
R1792 B.n824 B.n370 163.367
R1793 B.n824 B.n365 163.367
R1794 B.n832 B.n365 163.367
R1795 B.n832 B.n363 163.367
R1796 B.n837 B.n363 163.367
R1797 B.n837 B.n357 163.367
R1798 B.n845 B.n357 163.367
R1799 B.n846 B.n845 163.367
R1800 B.n846 B.n5 163.367
R1801 B.n6 B.n5 163.367
R1802 B.n7 B.n6 163.367
R1803 B.n852 B.n7 163.367
R1804 B.n853 B.n852 163.367
R1805 B.n853 B.n13 163.367
R1806 B.n14 B.n13 163.367
R1807 B.n15 B.n14 163.367
R1808 B.n858 B.n15 163.367
R1809 B.n858 B.n19 163.367
R1810 B.n20 B.n19 163.367
R1811 B.n21 B.n20 163.367
R1812 B.n863 B.n21 163.367
R1813 B.n863 B.n26 163.367
R1814 B.n27 B.n26 163.367
R1815 B.n28 B.n27 163.367
R1816 B.n868 B.n28 163.367
R1817 B.n868 B.n33 163.367
R1818 B.n34 B.n33 163.367
R1819 B.n35 B.n34 163.367
R1820 B.n873 B.n35 163.367
R1821 B.n873 B.n40 163.367
R1822 B.n41 B.n40 163.367
R1823 B.n42 B.n41 163.367
R1824 B.n878 B.n42 163.367
R1825 B.n878 B.n47 163.367
R1826 B.n48 B.n47 163.367
R1827 B.n49 B.n48 163.367
R1828 B.n883 B.n49 163.367
R1829 B.n883 B.n54 163.367
R1830 B.n55 B.n54 163.367
R1831 B.n56 B.n55 163.367
R1832 B.n888 B.n56 163.367
R1833 B.n888 B.n61 163.367
R1834 B.n62 B.n61 163.367
R1835 B.n63 B.n62 163.367
R1836 B.n893 B.n63 163.367
R1837 B.n893 B.n68 163.367
R1838 B.n69 B.n68 163.367
R1839 B.n70 B.n69 163.367
R1840 B.n898 B.n70 163.367
R1841 B.n898 B.n75 163.367
R1842 B.n76 B.n75 163.367
R1843 B.n77 B.n76 163.367
R1844 B.n136 B.n77 163.367
R1845 B.n714 B.n439 163.367
R1846 B.n714 B.n494 163.367
R1847 B.n710 B.n709 163.367
R1848 B.n706 B.n705 163.367
R1849 B.n702 B.n701 163.367
R1850 B.n698 B.n697 163.367
R1851 B.n694 B.n693 163.367
R1852 B.n690 B.n689 163.367
R1853 B.n686 B.n685 163.367
R1854 B.n682 B.n681 163.367
R1855 B.n678 B.n677 163.367
R1856 B.n674 B.n673 163.367
R1857 B.n670 B.n669 163.367
R1858 B.n666 B.n665 163.367
R1859 B.n662 B.n661 163.367
R1860 B.n658 B.n657 163.367
R1861 B.n654 B.n653 163.367
R1862 B.n650 B.n649 163.367
R1863 B.n646 B.n645 163.367
R1864 B.n642 B.n641 163.367
R1865 B.n638 B.n637 163.367
R1866 B.n634 B.n633 163.367
R1867 B.n630 B.n629 163.367
R1868 B.n626 B.n625 163.367
R1869 B.n622 B.n621 163.367
R1870 B.n617 B.n616 163.367
R1871 B.n613 B.n612 163.367
R1872 B.n609 B.n608 163.367
R1873 B.n605 B.n604 163.367
R1874 B.n601 B.n600 163.367
R1875 B.n596 B.n595 163.367
R1876 B.n592 B.n591 163.367
R1877 B.n588 B.n587 163.367
R1878 B.n584 B.n583 163.367
R1879 B.n580 B.n579 163.367
R1880 B.n576 B.n575 163.367
R1881 B.n572 B.n571 163.367
R1882 B.n568 B.n567 163.367
R1883 B.n564 B.n563 163.367
R1884 B.n560 B.n559 163.367
R1885 B.n556 B.n555 163.367
R1886 B.n552 B.n551 163.367
R1887 B.n548 B.n547 163.367
R1888 B.n544 B.n543 163.367
R1889 B.n540 B.n539 163.367
R1890 B.n536 B.n535 163.367
R1891 B.n532 B.n531 163.367
R1892 B.n528 B.n527 163.367
R1893 B.n524 B.n523 163.367
R1894 B.n520 B.n519 163.367
R1895 B.n516 B.n515 163.367
R1896 B.n512 B.n511 163.367
R1897 B.n508 B.n507 163.367
R1898 B.n504 B.n503 163.367
R1899 B.n500 B.n493 163.367
R1900 B.n721 B.n437 163.367
R1901 B.n721 B.n431 163.367
R1902 B.n729 B.n431 163.367
R1903 B.n729 B.n429 163.367
R1904 B.n733 B.n429 163.367
R1905 B.n733 B.n423 163.367
R1906 B.n741 B.n423 163.367
R1907 B.n741 B.n421 163.367
R1908 B.n745 B.n421 163.367
R1909 B.n745 B.n415 163.367
R1910 B.n753 B.n415 163.367
R1911 B.n753 B.n413 163.367
R1912 B.n757 B.n413 163.367
R1913 B.n757 B.n407 163.367
R1914 B.n765 B.n407 163.367
R1915 B.n765 B.n405 163.367
R1916 B.n769 B.n405 163.367
R1917 B.n769 B.n399 163.367
R1918 B.n777 B.n399 163.367
R1919 B.n777 B.n397 163.367
R1920 B.n781 B.n397 163.367
R1921 B.n781 B.n391 163.367
R1922 B.n790 B.n391 163.367
R1923 B.n790 B.n389 163.367
R1924 B.n794 B.n389 163.367
R1925 B.n794 B.n384 163.367
R1926 B.n802 B.n384 163.367
R1927 B.n802 B.n382 163.367
R1928 B.n806 B.n382 163.367
R1929 B.n806 B.n376 163.367
R1930 B.n814 B.n376 163.367
R1931 B.n814 B.n374 163.367
R1932 B.n818 B.n374 163.367
R1933 B.n818 B.n368 163.367
R1934 B.n826 B.n368 163.367
R1935 B.n826 B.n366 163.367
R1936 B.n830 B.n366 163.367
R1937 B.n830 B.n361 163.367
R1938 B.n839 B.n361 163.367
R1939 B.n839 B.n359 163.367
R1940 B.n843 B.n359 163.367
R1941 B.n843 B.n3 163.367
R1942 B.n998 B.n3 163.367
R1943 B.n994 B.n2 163.367
R1944 B.n994 B.n993 163.367
R1945 B.n993 B.n9 163.367
R1946 B.n989 B.n9 163.367
R1947 B.n989 B.n11 163.367
R1948 B.n985 B.n11 163.367
R1949 B.n985 B.n16 163.367
R1950 B.n981 B.n16 163.367
R1951 B.n981 B.n18 163.367
R1952 B.n977 B.n18 163.367
R1953 B.n977 B.n23 163.367
R1954 B.n973 B.n23 163.367
R1955 B.n973 B.n25 163.367
R1956 B.n969 B.n25 163.367
R1957 B.n969 B.n30 163.367
R1958 B.n965 B.n30 163.367
R1959 B.n965 B.n32 163.367
R1960 B.n961 B.n32 163.367
R1961 B.n961 B.n36 163.367
R1962 B.n957 B.n36 163.367
R1963 B.n957 B.n38 163.367
R1964 B.n953 B.n38 163.367
R1965 B.n953 B.n44 163.367
R1966 B.n949 B.n44 163.367
R1967 B.n949 B.n46 163.367
R1968 B.n945 B.n46 163.367
R1969 B.n945 B.n51 163.367
R1970 B.n941 B.n51 163.367
R1971 B.n941 B.n53 163.367
R1972 B.n937 B.n53 163.367
R1973 B.n937 B.n58 163.367
R1974 B.n933 B.n58 163.367
R1975 B.n933 B.n60 163.367
R1976 B.n929 B.n60 163.367
R1977 B.n929 B.n65 163.367
R1978 B.n925 B.n65 163.367
R1979 B.n925 B.n67 163.367
R1980 B.n921 B.n67 163.367
R1981 B.n921 B.n72 163.367
R1982 B.n917 B.n72 163.367
R1983 B.n917 B.n74 163.367
R1984 B.n913 B.n74 163.367
R1985 B.n913 B.n79 163.367
R1986 B.n141 B.n140 77.7702
R1987 B.n138 B.n137 77.7702
R1988 B.n498 B.n497 77.7702
R1989 B.n496 B.n495 77.7702
R1990 B.n909 B.n908 71.676
R1991 B.n143 B.n82 71.676
R1992 B.n147 B.n83 71.676
R1993 B.n151 B.n84 71.676
R1994 B.n155 B.n85 71.676
R1995 B.n159 B.n86 71.676
R1996 B.n163 B.n87 71.676
R1997 B.n167 B.n88 71.676
R1998 B.n171 B.n89 71.676
R1999 B.n175 B.n90 71.676
R2000 B.n179 B.n91 71.676
R2001 B.n183 B.n92 71.676
R2002 B.n187 B.n93 71.676
R2003 B.n191 B.n94 71.676
R2004 B.n195 B.n95 71.676
R2005 B.n199 B.n96 71.676
R2006 B.n203 B.n97 71.676
R2007 B.n207 B.n98 71.676
R2008 B.n211 B.n99 71.676
R2009 B.n215 B.n100 71.676
R2010 B.n219 B.n101 71.676
R2011 B.n223 B.n102 71.676
R2012 B.n227 B.n103 71.676
R2013 B.n231 B.n104 71.676
R2014 B.n235 B.n105 71.676
R2015 B.n239 B.n106 71.676
R2016 B.n243 B.n107 71.676
R2017 B.n247 B.n108 71.676
R2018 B.n251 B.n109 71.676
R2019 B.n255 B.n110 71.676
R2020 B.n259 B.n111 71.676
R2021 B.n263 B.n112 71.676
R2022 B.n267 B.n113 71.676
R2023 B.n271 B.n114 71.676
R2024 B.n275 B.n115 71.676
R2025 B.n279 B.n116 71.676
R2026 B.n283 B.n117 71.676
R2027 B.n287 B.n118 71.676
R2028 B.n291 B.n119 71.676
R2029 B.n295 B.n120 71.676
R2030 B.n299 B.n121 71.676
R2031 B.n303 B.n122 71.676
R2032 B.n307 B.n123 71.676
R2033 B.n311 B.n124 71.676
R2034 B.n315 B.n125 71.676
R2035 B.n319 B.n126 71.676
R2036 B.n323 B.n127 71.676
R2037 B.n327 B.n128 71.676
R2038 B.n331 B.n129 71.676
R2039 B.n335 B.n130 71.676
R2040 B.n339 B.n131 71.676
R2041 B.n343 B.n132 71.676
R2042 B.n347 B.n133 71.676
R2043 B.n351 B.n134 71.676
R2044 B.n906 B.n135 71.676
R2045 B.n906 B.n905 71.676
R2046 B.n353 B.n134 71.676
R2047 B.n350 B.n133 71.676
R2048 B.n346 B.n132 71.676
R2049 B.n342 B.n131 71.676
R2050 B.n338 B.n130 71.676
R2051 B.n334 B.n129 71.676
R2052 B.n330 B.n128 71.676
R2053 B.n326 B.n127 71.676
R2054 B.n322 B.n126 71.676
R2055 B.n318 B.n125 71.676
R2056 B.n314 B.n124 71.676
R2057 B.n310 B.n123 71.676
R2058 B.n306 B.n122 71.676
R2059 B.n302 B.n121 71.676
R2060 B.n298 B.n120 71.676
R2061 B.n294 B.n119 71.676
R2062 B.n290 B.n118 71.676
R2063 B.n286 B.n117 71.676
R2064 B.n282 B.n116 71.676
R2065 B.n278 B.n115 71.676
R2066 B.n274 B.n114 71.676
R2067 B.n270 B.n113 71.676
R2068 B.n266 B.n112 71.676
R2069 B.n262 B.n111 71.676
R2070 B.n258 B.n110 71.676
R2071 B.n254 B.n109 71.676
R2072 B.n250 B.n108 71.676
R2073 B.n246 B.n107 71.676
R2074 B.n242 B.n106 71.676
R2075 B.n238 B.n105 71.676
R2076 B.n234 B.n104 71.676
R2077 B.n230 B.n103 71.676
R2078 B.n226 B.n102 71.676
R2079 B.n222 B.n101 71.676
R2080 B.n218 B.n100 71.676
R2081 B.n214 B.n99 71.676
R2082 B.n210 B.n98 71.676
R2083 B.n206 B.n97 71.676
R2084 B.n202 B.n96 71.676
R2085 B.n198 B.n95 71.676
R2086 B.n194 B.n94 71.676
R2087 B.n190 B.n93 71.676
R2088 B.n186 B.n92 71.676
R2089 B.n182 B.n91 71.676
R2090 B.n178 B.n90 71.676
R2091 B.n174 B.n89 71.676
R2092 B.n170 B.n88 71.676
R2093 B.n166 B.n87 71.676
R2094 B.n162 B.n86 71.676
R2095 B.n158 B.n85 71.676
R2096 B.n154 B.n84 71.676
R2097 B.n150 B.n83 71.676
R2098 B.n146 B.n82 71.676
R2099 B.n908 B.n81 71.676
R2100 B.n717 B.n716 71.676
R2101 B.n494 B.n440 71.676
R2102 B.n709 B.n441 71.676
R2103 B.n705 B.n442 71.676
R2104 B.n701 B.n443 71.676
R2105 B.n697 B.n444 71.676
R2106 B.n693 B.n445 71.676
R2107 B.n689 B.n446 71.676
R2108 B.n685 B.n447 71.676
R2109 B.n681 B.n448 71.676
R2110 B.n677 B.n449 71.676
R2111 B.n673 B.n450 71.676
R2112 B.n669 B.n451 71.676
R2113 B.n665 B.n452 71.676
R2114 B.n661 B.n453 71.676
R2115 B.n657 B.n454 71.676
R2116 B.n653 B.n455 71.676
R2117 B.n649 B.n456 71.676
R2118 B.n645 B.n457 71.676
R2119 B.n641 B.n458 71.676
R2120 B.n637 B.n459 71.676
R2121 B.n633 B.n460 71.676
R2122 B.n629 B.n461 71.676
R2123 B.n625 B.n462 71.676
R2124 B.n621 B.n463 71.676
R2125 B.n616 B.n464 71.676
R2126 B.n612 B.n465 71.676
R2127 B.n608 B.n466 71.676
R2128 B.n604 B.n467 71.676
R2129 B.n600 B.n468 71.676
R2130 B.n595 B.n469 71.676
R2131 B.n591 B.n470 71.676
R2132 B.n587 B.n471 71.676
R2133 B.n583 B.n472 71.676
R2134 B.n579 B.n473 71.676
R2135 B.n575 B.n474 71.676
R2136 B.n571 B.n475 71.676
R2137 B.n567 B.n476 71.676
R2138 B.n563 B.n477 71.676
R2139 B.n559 B.n478 71.676
R2140 B.n555 B.n479 71.676
R2141 B.n551 B.n480 71.676
R2142 B.n547 B.n481 71.676
R2143 B.n543 B.n482 71.676
R2144 B.n539 B.n483 71.676
R2145 B.n535 B.n484 71.676
R2146 B.n531 B.n485 71.676
R2147 B.n527 B.n486 71.676
R2148 B.n523 B.n487 71.676
R2149 B.n519 B.n488 71.676
R2150 B.n515 B.n489 71.676
R2151 B.n511 B.n490 71.676
R2152 B.n507 B.n491 71.676
R2153 B.n503 B.n492 71.676
R2154 B.n716 B.n439 71.676
R2155 B.n710 B.n440 71.676
R2156 B.n706 B.n441 71.676
R2157 B.n702 B.n442 71.676
R2158 B.n698 B.n443 71.676
R2159 B.n694 B.n444 71.676
R2160 B.n690 B.n445 71.676
R2161 B.n686 B.n446 71.676
R2162 B.n682 B.n447 71.676
R2163 B.n678 B.n448 71.676
R2164 B.n674 B.n449 71.676
R2165 B.n670 B.n450 71.676
R2166 B.n666 B.n451 71.676
R2167 B.n662 B.n452 71.676
R2168 B.n658 B.n453 71.676
R2169 B.n654 B.n454 71.676
R2170 B.n650 B.n455 71.676
R2171 B.n646 B.n456 71.676
R2172 B.n642 B.n457 71.676
R2173 B.n638 B.n458 71.676
R2174 B.n634 B.n459 71.676
R2175 B.n630 B.n460 71.676
R2176 B.n626 B.n461 71.676
R2177 B.n622 B.n462 71.676
R2178 B.n617 B.n463 71.676
R2179 B.n613 B.n464 71.676
R2180 B.n609 B.n465 71.676
R2181 B.n605 B.n466 71.676
R2182 B.n601 B.n467 71.676
R2183 B.n596 B.n468 71.676
R2184 B.n592 B.n469 71.676
R2185 B.n588 B.n470 71.676
R2186 B.n584 B.n471 71.676
R2187 B.n580 B.n472 71.676
R2188 B.n576 B.n473 71.676
R2189 B.n572 B.n474 71.676
R2190 B.n568 B.n475 71.676
R2191 B.n564 B.n476 71.676
R2192 B.n560 B.n477 71.676
R2193 B.n556 B.n478 71.676
R2194 B.n552 B.n479 71.676
R2195 B.n548 B.n480 71.676
R2196 B.n544 B.n481 71.676
R2197 B.n540 B.n482 71.676
R2198 B.n536 B.n483 71.676
R2199 B.n532 B.n484 71.676
R2200 B.n528 B.n485 71.676
R2201 B.n524 B.n486 71.676
R2202 B.n520 B.n487 71.676
R2203 B.n516 B.n488 71.676
R2204 B.n512 B.n489 71.676
R2205 B.n508 B.n490 71.676
R2206 B.n504 B.n491 71.676
R2207 B.n500 B.n492 71.676
R2208 B.n999 B.n998 71.676
R2209 B.n999 B.n2 71.676
R2210 B.n715 B.n436 67.2637
R2211 B.n907 B.n78 67.2637
R2212 B.n142 B.n141 59.5399
R2213 B.n139 B.n138 59.5399
R2214 B.n598 B.n498 59.5399
R2215 B.n619 B.n496 59.5399
R2216 B.n722 B.n436 37.1867
R2217 B.n722 B.n432 37.1867
R2218 B.n728 B.n432 37.1867
R2219 B.n728 B.n428 37.1867
R2220 B.n734 B.n428 37.1867
R2221 B.n734 B.n424 37.1867
R2222 B.n740 B.n424 37.1867
R2223 B.n740 B.n420 37.1867
R2224 B.n746 B.n420 37.1867
R2225 B.n752 B.n416 37.1867
R2226 B.n752 B.n412 37.1867
R2227 B.n758 B.n412 37.1867
R2228 B.n758 B.n408 37.1867
R2229 B.n764 B.n408 37.1867
R2230 B.n764 B.n404 37.1867
R2231 B.n770 B.n404 37.1867
R2232 B.n770 B.n400 37.1867
R2233 B.n776 B.n400 37.1867
R2234 B.n776 B.n396 37.1867
R2235 B.n782 B.n396 37.1867
R2236 B.n782 B.n392 37.1867
R2237 B.n789 B.n392 37.1867
R2238 B.n789 B.n788 37.1867
R2239 B.n795 B.n385 37.1867
R2240 B.n801 B.n385 37.1867
R2241 B.n801 B.n381 37.1867
R2242 B.n807 B.n381 37.1867
R2243 B.n807 B.n377 37.1867
R2244 B.n813 B.n377 37.1867
R2245 B.n813 B.n373 37.1867
R2246 B.n819 B.n373 37.1867
R2247 B.n819 B.n369 37.1867
R2248 B.n825 B.n369 37.1867
R2249 B.n825 B.t3 37.1867
R2250 B.n831 B.t3 37.1867
R2251 B.n831 B.n362 37.1867
R2252 B.n838 B.n362 37.1867
R2253 B.n838 B.n358 37.1867
R2254 B.n844 B.n358 37.1867
R2255 B.n844 B.n4 37.1867
R2256 B.n997 B.n4 37.1867
R2257 B.n997 B.n996 37.1867
R2258 B.n996 B.n995 37.1867
R2259 B.n995 B.n8 37.1867
R2260 B.n12 B.n8 37.1867
R2261 B.n988 B.n12 37.1867
R2262 B.n988 B.n987 37.1867
R2263 B.n987 B.n986 37.1867
R2264 B.n986 B.t2 37.1867
R2265 B.n980 B.t2 37.1867
R2266 B.n980 B.n979 37.1867
R2267 B.n979 B.n978 37.1867
R2268 B.n978 B.n22 37.1867
R2269 B.n972 B.n22 37.1867
R2270 B.n972 B.n971 37.1867
R2271 B.n971 B.n970 37.1867
R2272 B.n970 B.n29 37.1867
R2273 B.n964 B.n29 37.1867
R2274 B.n964 B.n963 37.1867
R2275 B.n963 B.n962 37.1867
R2276 B.n956 B.n39 37.1867
R2277 B.n956 B.n955 37.1867
R2278 B.n955 B.n954 37.1867
R2279 B.n954 B.n43 37.1867
R2280 B.n948 B.n43 37.1867
R2281 B.n948 B.n947 37.1867
R2282 B.n947 B.n946 37.1867
R2283 B.n946 B.n50 37.1867
R2284 B.n940 B.n50 37.1867
R2285 B.n940 B.n939 37.1867
R2286 B.n939 B.n938 37.1867
R2287 B.n938 B.n57 37.1867
R2288 B.n932 B.n57 37.1867
R2289 B.n932 B.n931 37.1867
R2290 B.n930 B.n64 37.1867
R2291 B.n924 B.n64 37.1867
R2292 B.n924 B.n923 37.1867
R2293 B.n923 B.n922 37.1867
R2294 B.n922 B.n71 37.1867
R2295 B.n916 B.n71 37.1867
R2296 B.n916 B.n915 37.1867
R2297 B.n915 B.n914 37.1867
R2298 B.n914 B.n78 37.1867
R2299 B.n904 B.n903 29.8151
R2300 B.n719 B.n718 29.8151
R2301 B.n499 B.n434 29.8151
R2302 B.n911 B.n910 29.8151
R2303 B.t12 B.n416 29.5307
R2304 B.n795 B.t1 29.5307
R2305 B.n962 B.t0 29.5307
R2306 B.n931 B.t5 29.5307
R2307 B B.n1000 18.0485
R2308 B.n720 B.n719 10.6151
R2309 B.n720 B.n430 10.6151
R2310 B.n730 B.n430 10.6151
R2311 B.n731 B.n730 10.6151
R2312 B.n732 B.n731 10.6151
R2313 B.n732 B.n422 10.6151
R2314 B.n742 B.n422 10.6151
R2315 B.n743 B.n742 10.6151
R2316 B.n744 B.n743 10.6151
R2317 B.n744 B.n414 10.6151
R2318 B.n754 B.n414 10.6151
R2319 B.n755 B.n754 10.6151
R2320 B.n756 B.n755 10.6151
R2321 B.n756 B.n406 10.6151
R2322 B.n766 B.n406 10.6151
R2323 B.n767 B.n766 10.6151
R2324 B.n768 B.n767 10.6151
R2325 B.n768 B.n398 10.6151
R2326 B.n778 B.n398 10.6151
R2327 B.n779 B.n778 10.6151
R2328 B.n780 B.n779 10.6151
R2329 B.n780 B.n390 10.6151
R2330 B.n791 B.n390 10.6151
R2331 B.n792 B.n791 10.6151
R2332 B.n793 B.n792 10.6151
R2333 B.n793 B.n383 10.6151
R2334 B.n803 B.n383 10.6151
R2335 B.n804 B.n803 10.6151
R2336 B.n805 B.n804 10.6151
R2337 B.n805 B.n375 10.6151
R2338 B.n815 B.n375 10.6151
R2339 B.n816 B.n815 10.6151
R2340 B.n817 B.n816 10.6151
R2341 B.n817 B.n367 10.6151
R2342 B.n827 B.n367 10.6151
R2343 B.n828 B.n827 10.6151
R2344 B.n829 B.n828 10.6151
R2345 B.n829 B.n360 10.6151
R2346 B.n840 B.n360 10.6151
R2347 B.n841 B.n840 10.6151
R2348 B.n842 B.n841 10.6151
R2349 B.n842 B.n0 10.6151
R2350 B.n718 B.n438 10.6151
R2351 B.n713 B.n438 10.6151
R2352 B.n713 B.n712 10.6151
R2353 B.n712 B.n711 10.6151
R2354 B.n711 B.n708 10.6151
R2355 B.n708 B.n707 10.6151
R2356 B.n707 B.n704 10.6151
R2357 B.n704 B.n703 10.6151
R2358 B.n703 B.n700 10.6151
R2359 B.n700 B.n699 10.6151
R2360 B.n699 B.n696 10.6151
R2361 B.n696 B.n695 10.6151
R2362 B.n695 B.n692 10.6151
R2363 B.n692 B.n691 10.6151
R2364 B.n691 B.n688 10.6151
R2365 B.n688 B.n687 10.6151
R2366 B.n687 B.n684 10.6151
R2367 B.n684 B.n683 10.6151
R2368 B.n683 B.n680 10.6151
R2369 B.n680 B.n679 10.6151
R2370 B.n679 B.n676 10.6151
R2371 B.n676 B.n675 10.6151
R2372 B.n675 B.n672 10.6151
R2373 B.n672 B.n671 10.6151
R2374 B.n671 B.n668 10.6151
R2375 B.n668 B.n667 10.6151
R2376 B.n667 B.n664 10.6151
R2377 B.n664 B.n663 10.6151
R2378 B.n663 B.n660 10.6151
R2379 B.n660 B.n659 10.6151
R2380 B.n659 B.n656 10.6151
R2381 B.n656 B.n655 10.6151
R2382 B.n655 B.n652 10.6151
R2383 B.n652 B.n651 10.6151
R2384 B.n651 B.n648 10.6151
R2385 B.n648 B.n647 10.6151
R2386 B.n647 B.n644 10.6151
R2387 B.n644 B.n643 10.6151
R2388 B.n643 B.n640 10.6151
R2389 B.n640 B.n639 10.6151
R2390 B.n639 B.n636 10.6151
R2391 B.n636 B.n635 10.6151
R2392 B.n635 B.n632 10.6151
R2393 B.n632 B.n631 10.6151
R2394 B.n631 B.n628 10.6151
R2395 B.n628 B.n627 10.6151
R2396 B.n627 B.n624 10.6151
R2397 B.n624 B.n623 10.6151
R2398 B.n623 B.n620 10.6151
R2399 B.n618 B.n615 10.6151
R2400 B.n615 B.n614 10.6151
R2401 B.n614 B.n611 10.6151
R2402 B.n611 B.n610 10.6151
R2403 B.n610 B.n607 10.6151
R2404 B.n607 B.n606 10.6151
R2405 B.n606 B.n603 10.6151
R2406 B.n603 B.n602 10.6151
R2407 B.n602 B.n599 10.6151
R2408 B.n597 B.n594 10.6151
R2409 B.n594 B.n593 10.6151
R2410 B.n593 B.n590 10.6151
R2411 B.n590 B.n589 10.6151
R2412 B.n589 B.n586 10.6151
R2413 B.n586 B.n585 10.6151
R2414 B.n585 B.n582 10.6151
R2415 B.n582 B.n581 10.6151
R2416 B.n581 B.n578 10.6151
R2417 B.n578 B.n577 10.6151
R2418 B.n577 B.n574 10.6151
R2419 B.n574 B.n573 10.6151
R2420 B.n573 B.n570 10.6151
R2421 B.n570 B.n569 10.6151
R2422 B.n569 B.n566 10.6151
R2423 B.n566 B.n565 10.6151
R2424 B.n565 B.n562 10.6151
R2425 B.n562 B.n561 10.6151
R2426 B.n561 B.n558 10.6151
R2427 B.n558 B.n557 10.6151
R2428 B.n557 B.n554 10.6151
R2429 B.n554 B.n553 10.6151
R2430 B.n553 B.n550 10.6151
R2431 B.n550 B.n549 10.6151
R2432 B.n549 B.n546 10.6151
R2433 B.n546 B.n545 10.6151
R2434 B.n545 B.n542 10.6151
R2435 B.n542 B.n541 10.6151
R2436 B.n541 B.n538 10.6151
R2437 B.n538 B.n537 10.6151
R2438 B.n537 B.n534 10.6151
R2439 B.n534 B.n533 10.6151
R2440 B.n533 B.n530 10.6151
R2441 B.n530 B.n529 10.6151
R2442 B.n529 B.n526 10.6151
R2443 B.n526 B.n525 10.6151
R2444 B.n525 B.n522 10.6151
R2445 B.n522 B.n521 10.6151
R2446 B.n521 B.n518 10.6151
R2447 B.n518 B.n517 10.6151
R2448 B.n517 B.n514 10.6151
R2449 B.n514 B.n513 10.6151
R2450 B.n513 B.n510 10.6151
R2451 B.n510 B.n509 10.6151
R2452 B.n509 B.n506 10.6151
R2453 B.n506 B.n505 10.6151
R2454 B.n505 B.n502 10.6151
R2455 B.n502 B.n501 10.6151
R2456 B.n501 B.n499 10.6151
R2457 B.n724 B.n434 10.6151
R2458 B.n725 B.n724 10.6151
R2459 B.n726 B.n725 10.6151
R2460 B.n726 B.n426 10.6151
R2461 B.n736 B.n426 10.6151
R2462 B.n737 B.n736 10.6151
R2463 B.n738 B.n737 10.6151
R2464 B.n738 B.n418 10.6151
R2465 B.n748 B.n418 10.6151
R2466 B.n749 B.n748 10.6151
R2467 B.n750 B.n749 10.6151
R2468 B.n750 B.n410 10.6151
R2469 B.n760 B.n410 10.6151
R2470 B.n761 B.n760 10.6151
R2471 B.n762 B.n761 10.6151
R2472 B.n762 B.n402 10.6151
R2473 B.n772 B.n402 10.6151
R2474 B.n773 B.n772 10.6151
R2475 B.n774 B.n773 10.6151
R2476 B.n774 B.n394 10.6151
R2477 B.n784 B.n394 10.6151
R2478 B.n785 B.n784 10.6151
R2479 B.n786 B.n785 10.6151
R2480 B.n786 B.n387 10.6151
R2481 B.n797 B.n387 10.6151
R2482 B.n798 B.n797 10.6151
R2483 B.n799 B.n798 10.6151
R2484 B.n799 B.n379 10.6151
R2485 B.n809 B.n379 10.6151
R2486 B.n810 B.n809 10.6151
R2487 B.n811 B.n810 10.6151
R2488 B.n811 B.n371 10.6151
R2489 B.n821 B.n371 10.6151
R2490 B.n822 B.n821 10.6151
R2491 B.n823 B.n822 10.6151
R2492 B.n823 B.n364 10.6151
R2493 B.n833 B.n364 10.6151
R2494 B.n834 B.n833 10.6151
R2495 B.n836 B.n834 10.6151
R2496 B.n836 B.n835 10.6151
R2497 B.n835 B.n356 10.6151
R2498 B.n847 B.n356 10.6151
R2499 B.n848 B.n847 10.6151
R2500 B.n849 B.n848 10.6151
R2501 B.n850 B.n849 10.6151
R2502 B.n851 B.n850 10.6151
R2503 B.n854 B.n851 10.6151
R2504 B.n855 B.n854 10.6151
R2505 B.n856 B.n855 10.6151
R2506 B.n857 B.n856 10.6151
R2507 B.n859 B.n857 10.6151
R2508 B.n860 B.n859 10.6151
R2509 B.n861 B.n860 10.6151
R2510 B.n862 B.n861 10.6151
R2511 B.n864 B.n862 10.6151
R2512 B.n865 B.n864 10.6151
R2513 B.n866 B.n865 10.6151
R2514 B.n867 B.n866 10.6151
R2515 B.n869 B.n867 10.6151
R2516 B.n870 B.n869 10.6151
R2517 B.n871 B.n870 10.6151
R2518 B.n872 B.n871 10.6151
R2519 B.n874 B.n872 10.6151
R2520 B.n875 B.n874 10.6151
R2521 B.n876 B.n875 10.6151
R2522 B.n877 B.n876 10.6151
R2523 B.n879 B.n877 10.6151
R2524 B.n880 B.n879 10.6151
R2525 B.n881 B.n880 10.6151
R2526 B.n882 B.n881 10.6151
R2527 B.n884 B.n882 10.6151
R2528 B.n885 B.n884 10.6151
R2529 B.n886 B.n885 10.6151
R2530 B.n887 B.n886 10.6151
R2531 B.n889 B.n887 10.6151
R2532 B.n890 B.n889 10.6151
R2533 B.n891 B.n890 10.6151
R2534 B.n892 B.n891 10.6151
R2535 B.n894 B.n892 10.6151
R2536 B.n895 B.n894 10.6151
R2537 B.n896 B.n895 10.6151
R2538 B.n897 B.n896 10.6151
R2539 B.n899 B.n897 10.6151
R2540 B.n900 B.n899 10.6151
R2541 B.n901 B.n900 10.6151
R2542 B.n902 B.n901 10.6151
R2543 B.n903 B.n902 10.6151
R2544 B.n992 B.n1 10.6151
R2545 B.n992 B.n991 10.6151
R2546 B.n991 B.n990 10.6151
R2547 B.n990 B.n10 10.6151
R2548 B.n984 B.n10 10.6151
R2549 B.n984 B.n983 10.6151
R2550 B.n983 B.n982 10.6151
R2551 B.n982 B.n17 10.6151
R2552 B.n976 B.n17 10.6151
R2553 B.n976 B.n975 10.6151
R2554 B.n975 B.n974 10.6151
R2555 B.n974 B.n24 10.6151
R2556 B.n968 B.n24 10.6151
R2557 B.n968 B.n967 10.6151
R2558 B.n967 B.n966 10.6151
R2559 B.n966 B.n31 10.6151
R2560 B.n960 B.n31 10.6151
R2561 B.n960 B.n959 10.6151
R2562 B.n959 B.n958 10.6151
R2563 B.n958 B.n37 10.6151
R2564 B.n952 B.n37 10.6151
R2565 B.n952 B.n951 10.6151
R2566 B.n951 B.n950 10.6151
R2567 B.n950 B.n45 10.6151
R2568 B.n944 B.n45 10.6151
R2569 B.n944 B.n943 10.6151
R2570 B.n943 B.n942 10.6151
R2571 B.n942 B.n52 10.6151
R2572 B.n936 B.n52 10.6151
R2573 B.n936 B.n935 10.6151
R2574 B.n935 B.n934 10.6151
R2575 B.n934 B.n59 10.6151
R2576 B.n928 B.n59 10.6151
R2577 B.n928 B.n927 10.6151
R2578 B.n927 B.n926 10.6151
R2579 B.n926 B.n66 10.6151
R2580 B.n920 B.n66 10.6151
R2581 B.n920 B.n919 10.6151
R2582 B.n919 B.n918 10.6151
R2583 B.n918 B.n73 10.6151
R2584 B.n912 B.n73 10.6151
R2585 B.n912 B.n911 10.6151
R2586 B.n910 B.n80 10.6151
R2587 B.n144 B.n80 10.6151
R2588 B.n145 B.n144 10.6151
R2589 B.n148 B.n145 10.6151
R2590 B.n149 B.n148 10.6151
R2591 B.n152 B.n149 10.6151
R2592 B.n153 B.n152 10.6151
R2593 B.n156 B.n153 10.6151
R2594 B.n157 B.n156 10.6151
R2595 B.n160 B.n157 10.6151
R2596 B.n161 B.n160 10.6151
R2597 B.n164 B.n161 10.6151
R2598 B.n165 B.n164 10.6151
R2599 B.n168 B.n165 10.6151
R2600 B.n169 B.n168 10.6151
R2601 B.n172 B.n169 10.6151
R2602 B.n173 B.n172 10.6151
R2603 B.n176 B.n173 10.6151
R2604 B.n177 B.n176 10.6151
R2605 B.n180 B.n177 10.6151
R2606 B.n181 B.n180 10.6151
R2607 B.n184 B.n181 10.6151
R2608 B.n185 B.n184 10.6151
R2609 B.n188 B.n185 10.6151
R2610 B.n189 B.n188 10.6151
R2611 B.n192 B.n189 10.6151
R2612 B.n193 B.n192 10.6151
R2613 B.n196 B.n193 10.6151
R2614 B.n197 B.n196 10.6151
R2615 B.n200 B.n197 10.6151
R2616 B.n201 B.n200 10.6151
R2617 B.n204 B.n201 10.6151
R2618 B.n205 B.n204 10.6151
R2619 B.n208 B.n205 10.6151
R2620 B.n209 B.n208 10.6151
R2621 B.n212 B.n209 10.6151
R2622 B.n213 B.n212 10.6151
R2623 B.n216 B.n213 10.6151
R2624 B.n217 B.n216 10.6151
R2625 B.n220 B.n217 10.6151
R2626 B.n221 B.n220 10.6151
R2627 B.n224 B.n221 10.6151
R2628 B.n225 B.n224 10.6151
R2629 B.n228 B.n225 10.6151
R2630 B.n229 B.n228 10.6151
R2631 B.n232 B.n229 10.6151
R2632 B.n233 B.n232 10.6151
R2633 B.n236 B.n233 10.6151
R2634 B.n237 B.n236 10.6151
R2635 B.n241 B.n240 10.6151
R2636 B.n244 B.n241 10.6151
R2637 B.n245 B.n244 10.6151
R2638 B.n248 B.n245 10.6151
R2639 B.n249 B.n248 10.6151
R2640 B.n252 B.n249 10.6151
R2641 B.n253 B.n252 10.6151
R2642 B.n256 B.n253 10.6151
R2643 B.n257 B.n256 10.6151
R2644 B.n261 B.n260 10.6151
R2645 B.n264 B.n261 10.6151
R2646 B.n265 B.n264 10.6151
R2647 B.n268 B.n265 10.6151
R2648 B.n269 B.n268 10.6151
R2649 B.n272 B.n269 10.6151
R2650 B.n273 B.n272 10.6151
R2651 B.n276 B.n273 10.6151
R2652 B.n277 B.n276 10.6151
R2653 B.n280 B.n277 10.6151
R2654 B.n281 B.n280 10.6151
R2655 B.n284 B.n281 10.6151
R2656 B.n285 B.n284 10.6151
R2657 B.n288 B.n285 10.6151
R2658 B.n289 B.n288 10.6151
R2659 B.n292 B.n289 10.6151
R2660 B.n293 B.n292 10.6151
R2661 B.n296 B.n293 10.6151
R2662 B.n297 B.n296 10.6151
R2663 B.n300 B.n297 10.6151
R2664 B.n301 B.n300 10.6151
R2665 B.n304 B.n301 10.6151
R2666 B.n305 B.n304 10.6151
R2667 B.n308 B.n305 10.6151
R2668 B.n309 B.n308 10.6151
R2669 B.n312 B.n309 10.6151
R2670 B.n313 B.n312 10.6151
R2671 B.n316 B.n313 10.6151
R2672 B.n317 B.n316 10.6151
R2673 B.n320 B.n317 10.6151
R2674 B.n321 B.n320 10.6151
R2675 B.n324 B.n321 10.6151
R2676 B.n325 B.n324 10.6151
R2677 B.n328 B.n325 10.6151
R2678 B.n329 B.n328 10.6151
R2679 B.n332 B.n329 10.6151
R2680 B.n333 B.n332 10.6151
R2681 B.n336 B.n333 10.6151
R2682 B.n337 B.n336 10.6151
R2683 B.n340 B.n337 10.6151
R2684 B.n341 B.n340 10.6151
R2685 B.n344 B.n341 10.6151
R2686 B.n345 B.n344 10.6151
R2687 B.n348 B.n345 10.6151
R2688 B.n349 B.n348 10.6151
R2689 B.n352 B.n349 10.6151
R2690 B.n354 B.n352 10.6151
R2691 B.n355 B.n354 10.6151
R2692 B.n904 B.n355 10.6151
R2693 B.n620 B.n619 9.36635
R2694 B.n598 B.n597 9.36635
R2695 B.n237 B.n142 9.36635
R2696 B.n260 B.n139 9.36635
R2697 B.n1000 B.n0 8.11757
R2698 B.n1000 B.n1 8.11757
R2699 B.n746 B.t12 7.65648
R2700 B.n788 B.t1 7.65648
R2701 B.n39 B.t0 7.65648
R2702 B.t5 B.n930 7.65648
R2703 B.n619 B.n618 1.24928
R2704 B.n599 B.n598 1.24928
R2705 B.n240 B.n142 1.24928
R2706 B.n257 B.n139 1.24928
R2707 VP.n21 VP.n20 161.3
R2708 VP.n19 VP.n1 161.3
R2709 VP.n18 VP.n17 161.3
R2710 VP.n16 VP.n2 161.3
R2711 VP.n15 VP.n14 161.3
R2712 VP.n13 VP.n3 161.3
R2713 VP.n12 VP.n11 161.3
R2714 VP.n10 VP.n4 161.3
R2715 VP.n9 VP.n8 161.3
R2716 VP.n5 VP.t2 130.389
R2717 VP.n5 VP.t1 129.067
R2718 VP.n7 VP.t3 97.1864
R2719 VP.n0 VP.t0 97.1864
R2720 VP.n7 VP.n6 89.9996
R2721 VP.n22 VP.n0 89.9996
R2722 VP.n6 VP.n5 53.685
R2723 VP.n14 VP.n13 40.577
R2724 VP.n14 VP.n2 40.577
R2725 VP.n8 VP.n4 24.5923
R2726 VP.n12 VP.n4 24.5923
R2727 VP.n13 VP.n12 24.5923
R2728 VP.n18 VP.n2 24.5923
R2729 VP.n19 VP.n18 24.5923
R2730 VP.n20 VP.n19 24.5923
R2731 VP.n9 VP.n6 0.354861
R2732 VP.n22 VP.n21 0.354861
R2733 VP VP.n22 0.267071
R2734 VP.n8 VP.n7 0.246418
R2735 VP.n20 VP.n0 0.246418
R2736 VP.n10 VP.n9 0.189894
R2737 VP.n11 VP.n10 0.189894
R2738 VP.n11 VP.n3 0.189894
R2739 VP.n15 VP.n3 0.189894
R2740 VP.n16 VP.n15 0.189894
R2741 VP.n17 VP.n16 0.189894
R2742 VP.n17 VP.n1 0.189894
R2743 VP.n21 VP.n1 0.189894
R2744 VDD1 VDD1.n1 112.204
R2745 VDD1 VDD1.n0 64.8579
R2746 VDD1.n0 VDD1.t1 1.33473
R2747 VDD1.n0 VDD1.t2 1.33473
R2748 VDD1.n1 VDD1.t0 1.33473
R2749 VDD1.n1 VDD1.t3 1.33473
C0 VN VDD1 0.150163f
C1 VDD1 VP 6.43683f
C2 VDD1 VDD2 1.28638f
C3 VTAIL VDD1 6.30116f
C4 VN VP 7.49471f
C5 VN VDD2 6.12479f
C6 VN VTAIL 6.05615f
C7 VDD2 VP 0.463215f
C8 VTAIL VP 6.07026f
C9 VTAIL VDD2 6.36261f
C10 VDD2 B 4.597123f
C11 VDD1 B 9.41948f
C12 VTAIL B 12.394438f
C13 VN B 13.013169f
C14 VP B 11.430575f
C15 VDD1.t1 B 0.31915f
C16 VDD1.t2 B 0.31915f
C17 VDD1.n0 B 2.8882f
C18 VDD1.t0 B 0.31915f
C19 VDD1.t3 B 0.31915f
C20 VDD1.n1 B 3.73843f
C21 VP.t0 B 2.98997f
C22 VP.n0 B 1.10748f
C23 VP.n1 B 0.019985f
C24 VP.n2 B 0.039512f
C25 VP.n3 B 0.019985f
C26 VP.n4 B 0.037061f
C27 VP.t2 B 3.29521f
C28 VP.t1 B 3.28351f
C29 VP.n5 B 3.3692f
C30 VP.n6 B 1.27311f
C31 VP.t3 B 2.98997f
C32 VP.n7 B 1.10748f
C33 VP.n8 B 0.018948f
C34 VP.n9 B 0.032251f
C35 VP.n10 B 0.019985f
C36 VP.n11 B 0.019985f
C37 VP.n12 B 0.037061f
C38 VP.n13 B 0.039512f
C39 VP.n14 B 0.016142f
C40 VP.n15 B 0.019985f
C41 VP.n16 B 0.019985f
C42 VP.n17 B 0.019985f
C43 VP.n18 B 0.037061f
C44 VP.n19 B 0.037061f
C45 VP.n20 B 0.018948f
C46 VP.n21 B 0.032251f
C47 VP.n22 B 0.061383f
C48 VDD2.t2 B 0.31663f
C49 VDD2.t3 B 0.31663f
C50 VDD2.n0 B 3.68127f
C51 VDD2.t1 B 0.31663f
C52 VDD2.t0 B 0.31663f
C53 VDD2.n1 B 2.86492f
C54 VDD2.n2 B 4.38073f
C55 VTAIL.n0 B 0.023072f
C56 VTAIL.n1 B 0.016414f
C57 VTAIL.n2 B 0.00882f
C58 VTAIL.n3 B 0.020848f
C59 VTAIL.n4 B 0.009339f
C60 VTAIL.n5 B 0.016414f
C61 VTAIL.n6 B 0.00882f
C62 VTAIL.n7 B 0.020848f
C63 VTAIL.n8 B 0.009339f
C64 VTAIL.n9 B 0.016414f
C65 VTAIL.n10 B 0.00882f
C66 VTAIL.n11 B 0.020848f
C67 VTAIL.n12 B 0.009339f
C68 VTAIL.n13 B 0.016414f
C69 VTAIL.n14 B 0.00882f
C70 VTAIL.n15 B 0.020848f
C71 VTAIL.n16 B 0.009339f
C72 VTAIL.n17 B 0.016414f
C73 VTAIL.n18 B 0.00882f
C74 VTAIL.n19 B 0.020848f
C75 VTAIL.n20 B 0.009339f
C76 VTAIL.n21 B 0.016414f
C77 VTAIL.n22 B 0.00882f
C78 VTAIL.n23 B 0.020848f
C79 VTAIL.n24 B 0.009339f
C80 VTAIL.n25 B 0.106399f
C81 VTAIL.t5 B 0.034367f
C82 VTAIL.n26 B 0.015636f
C83 VTAIL.n27 B 0.012316f
C84 VTAIL.n28 B 0.00882f
C85 VTAIL.n29 B 1.0559f
C86 VTAIL.n30 B 0.016414f
C87 VTAIL.n31 B 0.00882f
C88 VTAIL.n32 B 0.009339f
C89 VTAIL.n33 B 0.020848f
C90 VTAIL.n34 B 0.020848f
C91 VTAIL.n35 B 0.009339f
C92 VTAIL.n36 B 0.00882f
C93 VTAIL.n37 B 0.016414f
C94 VTAIL.n38 B 0.016414f
C95 VTAIL.n39 B 0.00882f
C96 VTAIL.n40 B 0.009339f
C97 VTAIL.n41 B 0.020848f
C98 VTAIL.n42 B 0.020848f
C99 VTAIL.n43 B 0.009339f
C100 VTAIL.n44 B 0.00882f
C101 VTAIL.n45 B 0.016414f
C102 VTAIL.n46 B 0.016414f
C103 VTAIL.n47 B 0.00882f
C104 VTAIL.n48 B 0.009339f
C105 VTAIL.n49 B 0.020848f
C106 VTAIL.n50 B 0.020848f
C107 VTAIL.n51 B 0.009339f
C108 VTAIL.n52 B 0.00882f
C109 VTAIL.n53 B 0.016414f
C110 VTAIL.n54 B 0.016414f
C111 VTAIL.n55 B 0.00882f
C112 VTAIL.n56 B 0.009339f
C113 VTAIL.n57 B 0.020848f
C114 VTAIL.n58 B 0.020848f
C115 VTAIL.n59 B 0.009339f
C116 VTAIL.n60 B 0.00882f
C117 VTAIL.n61 B 0.016414f
C118 VTAIL.n62 B 0.016414f
C119 VTAIL.n63 B 0.00882f
C120 VTAIL.n64 B 0.009339f
C121 VTAIL.n65 B 0.020848f
C122 VTAIL.n66 B 0.020848f
C123 VTAIL.n67 B 0.020848f
C124 VTAIL.n68 B 0.009339f
C125 VTAIL.n69 B 0.00882f
C126 VTAIL.n70 B 0.016414f
C127 VTAIL.n71 B 0.016414f
C128 VTAIL.n72 B 0.00882f
C129 VTAIL.n73 B 0.00908f
C130 VTAIL.n74 B 0.00908f
C131 VTAIL.n75 B 0.020848f
C132 VTAIL.n76 B 0.045133f
C133 VTAIL.n77 B 0.009339f
C134 VTAIL.n78 B 0.00882f
C135 VTAIL.n79 B 0.042426f
C136 VTAIL.n80 B 0.025385f
C137 VTAIL.n81 B 0.135903f
C138 VTAIL.n82 B 0.023072f
C139 VTAIL.n83 B 0.016414f
C140 VTAIL.n84 B 0.00882f
C141 VTAIL.n85 B 0.020848f
C142 VTAIL.n86 B 0.009339f
C143 VTAIL.n87 B 0.016414f
C144 VTAIL.n88 B 0.00882f
C145 VTAIL.n89 B 0.020848f
C146 VTAIL.n90 B 0.009339f
C147 VTAIL.n91 B 0.016414f
C148 VTAIL.n92 B 0.00882f
C149 VTAIL.n93 B 0.020848f
C150 VTAIL.n94 B 0.009339f
C151 VTAIL.n95 B 0.016414f
C152 VTAIL.n96 B 0.00882f
C153 VTAIL.n97 B 0.020848f
C154 VTAIL.n98 B 0.009339f
C155 VTAIL.n99 B 0.016414f
C156 VTAIL.n100 B 0.00882f
C157 VTAIL.n101 B 0.020848f
C158 VTAIL.n102 B 0.009339f
C159 VTAIL.n103 B 0.016414f
C160 VTAIL.n104 B 0.00882f
C161 VTAIL.n105 B 0.020848f
C162 VTAIL.n106 B 0.009339f
C163 VTAIL.n107 B 0.106399f
C164 VTAIL.t3 B 0.034367f
C165 VTAIL.n108 B 0.015636f
C166 VTAIL.n109 B 0.012316f
C167 VTAIL.n110 B 0.00882f
C168 VTAIL.n111 B 1.0559f
C169 VTAIL.n112 B 0.016414f
C170 VTAIL.n113 B 0.00882f
C171 VTAIL.n114 B 0.009339f
C172 VTAIL.n115 B 0.020848f
C173 VTAIL.n116 B 0.020848f
C174 VTAIL.n117 B 0.009339f
C175 VTAIL.n118 B 0.00882f
C176 VTAIL.n119 B 0.016414f
C177 VTAIL.n120 B 0.016414f
C178 VTAIL.n121 B 0.00882f
C179 VTAIL.n122 B 0.009339f
C180 VTAIL.n123 B 0.020848f
C181 VTAIL.n124 B 0.020848f
C182 VTAIL.n125 B 0.009339f
C183 VTAIL.n126 B 0.00882f
C184 VTAIL.n127 B 0.016414f
C185 VTAIL.n128 B 0.016414f
C186 VTAIL.n129 B 0.00882f
C187 VTAIL.n130 B 0.009339f
C188 VTAIL.n131 B 0.020848f
C189 VTAIL.n132 B 0.020848f
C190 VTAIL.n133 B 0.009339f
C191 VTAIL.n134 B 0.00882f
C192 VTAIL.n135 B 0.016414f
C193 VTAIL.n136 B 0.016414f
C194 VTAIL.n137 B 0.00882f
C195 VTAIL.n138 B 0.009339f
C196 VTAIL.n139 B 0.020848f
C197 VTAIL.n140 B 0.020848f
C198 VTAIL.n141 B 0.009339f
C199 VTAIL.n142 B 0.00882f
C200 VTAIL.n143 B 0.016414f
C201 VTAIL.n144 B 0.016414f
C202 VTAIL.n145 B 0.00882f
C203 VTAIL.n146 B 0.009339f
C204 VTAIL.n147 B 0.020848f
C205 VTAIL.n148 B 0.020848f
C206 VTAIL.n149 B 0.020848f
C207 VTAIL.n150 B 0.009339f
C208 VTAIL.n151 B 0.00882f
C209 VTAIL.n152 B 0.016414f
C210 VTAIL.n153 B 0.016414f
C211 VTAIL.n154 B 0.00882f
C212 VTAIL.n155 B 0.00908f
C213 VTAIL.n156 B 0.00908f
C214 VTAIL.n157 B 0.020848f
C215 VTAIL.n158 B 0.045133f
C216 VTAIL.n159 B 0.009339f
C217 VTAIL.n160 B 0.00882f
C218 VTAIL.n161 B 0.042426f
C219 VTAIL.n162 B 0.025385f
C220 VTAIL.n163 B 0.224244f
C221 VTAIL.n164 B 0.023072f
C222 VTAIL.n165 B 0.016414f
C223 VTAIL.n166 B 0.00882f
C224 VTAIL.n167 B 0.020848f
C225 VTAIL.n168 B 0.009339f
C226 VTAIL.n169 B 0.016414f
C227 VTAIL.n170 B 0.00882f
C228 VTAIL.n171 B 0.020848f
C229 VTAIL.n172 B 0.009339f
C230 VTAIL.n173 B 0.016414f
C231 VTAIL.n174 B 0.00882f
C232 VTAIL.n175 B 0.020848f
C233 VTAIL.n176 B 0.009339f
C234 VTAIL.n177 B 0.016414f
C235 VTAIL.n178 B 0.00882f
C236 VTAIL.n179 B 0.020848f
C237 VTAIL.n180 B 0.009339f
C238 VTAIL.n181 B 0.016414f
C239 VTAIL.n182 B 0.00882f
C240 VTAIL.n183 B 0.020848f
C241 VTAIL.n184 B 0.009339f
C242 VTAIL.n185 B 0.016414f
C243 VTAIL.n186 B 0.00882f
C244 VTAIL.n187 B 0.020848f
C245 VTAIL.n188 B 0.009339f
C246 VTAIL.n189 B 0.106399f
C247 VTAIL.t1 B 0.034367f
C248 VTAIL.n190 B 0.015636f
C249 VTAIL.n191 B 0.012316f
C250 VTAIL.n192 B 0.00882f
C251 VTAIL.n193 B 1.0559f
C252 VTAIL.n194 B 0.016414f
C253 VTAIL.n195 B 0.00882f
C254 VTAIL.n196 B 0.009339f
C255 VTAIL.n197 B 0.020848f
C256 VTAIL.n198 B 0.020848f
C257 VTAIL.n199 B 0.009339f
C258 VTAIL.n200 B 0.00882f
C259 VTAIL.n201 B 0.016414f
C260 VTAIL.n202 B 0.016414f
C261 VTAIL.n203 B 0.00882f
C262 VTAIL.n204 B 0.009339f
C263 VTAIL.n205 B 0.020848f
C264 VTAIL.n206 B 0.020848f
C265 VTAIL.n207 B 0.009339f
C266 VTAIL.n208 B 0.00882f
C267 VTAIL.n209 B 0.016414f
C268 VTAIL.n210 B 0.016414f
C269 VTAIL.n211 B 0.00882f
C270 VTAIL.n212 B 0.009339f
C271 VTAIL.n213 B 0.020848f
C272 VTAIL.n214 B 0.020848f
C273 VTAIL.n215 B 0.009339f
C274 VTAIL.n216 B 0.00882f
C275 VTAIL.n217 B 0.016414f
C276 VTAIL.n218 B 0.016414f
C277 VTAIL.n219 B 0.00882f
C278 VTAIL.n220 B 0.009339f
C279 VTAIL.n221 B 0.020848f
C280 VTAIL.n222 B 0.020848f
C281 VTAIL.n223 B 0.009339f
C282 VTAIL.n224 B 0.00882f
C283 VTAIL.n225 B 0.016414f
C284 VTAIL.n226 B 0.016414f
C285 VTAIL.n227 B 0.00882f
C286 VTAIL.n228 B 0.009339f
C287 VTAIL.n229 B 0.020848f
C288 VTAIL.n230 B 0.020848f
C289 VTAIL.n231 B 0.020848f
C290 VTAIL.n232 B 0.009339f
C291 VTAIL.n233 B 0.00882f
C292 VTAIL.n234 B 0.016414f
C293 VTAIL.n235 B 0.016414f
C294 VTAIL.n236 B 0.00882f
C295 VTAIL.n237 B 0.00908f
C296 VTAIL.n238 B 0.00908f
C297 VTAIL.n239 B 0.020848f
C298 VTAIL.n240 B 0.045133f
C299 VTAIL.n241 B 0.009339f
C300 VTAIL.n242 B 0.00882f
C301 VTAIL.n243 B 0.042426f
C302 VTAIL.n244 B 0.025385f
C303 VTAIL.n245 B 1.28184f
C304 VTAIL.n246 B 0.023072f
C305 VTAIL.n247 B 0.016414f
C306 VTAIL.n248 B 0.00882f
C307 VTAIL.n249 B 0.020848f
C308 VTAIL.n250 B 0.009339f
C309 VTAIL.n251 B 0.016414f
C310 VTAIL.n252 B 0.00882f
C311 VTAIL.n253 B 0.020848f
C312 VTAIL.n254 B 0.020848f
C313 VTAIL.n255 B 0.009339f
C314 VTAIL.n256 B 0.016414f
C315 VTAIL.n257 B 0.00882f
C316 VTAIL.n258 B 0.020848f
C317 VTAIL.n259 B 0.009339f
C318 VTAIL.n260 B 0.016414f
C319 VTAIL.n261 B 0.00882f
C320 VTAIL.n262 B 0.020848f
C321 VTAIL.n263 B 0.009339f
C322 VTAIL.n264 B 0.016414f
C323 VTAIL.n265 B 0.00882f
C324 VTAIL.n266 B 0.020848f
C325 VTAIL.n267 B 0.009339f
C326 VTAIL.n268 B 0.016414f
C327 VTAIL.n269 B 0.00882f
C328 VTAIL.n270 B 0.020848f
C329 VTAIL.n271 B 0.009339f
C330 VTAIL.n272 B 0.106399f
C331 VTAIL.t7 B 0.034367f
C332 VTAIL.n273 B 0.015636f
C333 VTAIL.n274 B 0.012316f
C334 VTAIL.n275 B 0.00882f
C335 VTAIL.n276 B 1.0559f
C336 VTAIL.n277 B 0.016414f
C337 VTAIL.n278 B 0.00882f
C338 VTAIL.n279 B 0.009339f
C339 VTAIL.n280 B 0.020848f
C340 VTAIL.n281 B 0.020848f
C341 VTAIL.n282 B 0.009339f
C342 VTAIL.n283 B 0.00882f
C343 VTAIL.n284 B 0.016414f
C344 VTAIL.n285 B 0.016414f
C345 VTAIL.n286 B 0.00882f
C346 VTAIL.n287 B 0.009339f
C347 VTAIL.n288 B 0.020848f
C348 VTAIL.n289 B 0.020848f
C349 VTAIL.n290 B 0.009339f
C350 VTAIL.n291 B 0.00882f
C351 VTAIL.n292 B 0.016414f
C352 VTAIL.n293 B 0.016414f
C353 VTAIL.n294 B 0.00882f
C354 VTAIL.n295 B 0.009339f
C355 VTAIL.n296 B 0.020848f
C356 VTAIL.n297 B 0.020848f
C357 VTAIL.n298 B 0.009339f
C358 VTAIL.n299 B 0.00882f
C359 VTAIL.n300 B 0.016414f
C360 VTAIL.n301 B 0.016414f
C361 VTAIL.n302 B 0.00882f
C362 VTAIL.n303 B 0.009339f
C363 VTAIL.n304 B 0.020848f
C364 VTAIL.n305 B 0.020848f
C365 VTAIL.n306 B 0.009339f
C366 VTAIL.n307 B 0.00882f
C367 VTAIL.n308 B 0.016414f
C368 VTAIL.n309 B 0.016414f
C369 VTAIL.n310 B 0.00882f
C370 VTAIL.n311 B 0.009339f
C371 VTAIL.n312 B 0.020848f
C372 VTAIL.n313 B 0.020848f
C373 VTAIL.n314 B 0.009339f
C374 VTAIL.n315 B 0.00882f
C375 VTAIL.n316 B 0.016414f
C376 VTAIL.n317 B 0.016414f
C377 VTAIL.n318 B 0.00882f
C378 VTAIL.n319 B 0.00908f
C379 VTAIL.n320 B 0.00908f
C380 VTAIL.n321 B 0.020848f
C381 VTAIL.n322 B 0.045133f
C382 VTAIL.n323 B 0.009339f
C383 VTAIL.n324 B 0.00882f
C384 VTAIL.n325 B 0.042426f
C385 VTAIL.n326 B 0.025385f
C386 VTAIL.n327 B 1.28184f
C387 VTAIL.n328 B 0.023072f
C388 VTAIL.n329 B 0.016414f
C389 VTAIL.n330 B 0.00882f
C390 VTAIL.n331 B 0.020848f
C391 VTAIL.n332 B 0.009339f
C392 VTAIL.n333 B 0.016414f
C393 VTAIL.n334 B 0.00882f
C394 VTAIL.n335 B 0.020848f
C395 VTAIL.n336 B 0.020848f
C396 VTAIL.n337 B 0.009339f
C397 VTAIL.n338 B 0.016414f
C398 VTAIL.n339 B 0.00882f
C399 VTAIL.n340 B 0.020848f
C400 VTAIL.n341 B 0.009339f
C401 VTAIL.n342 B 0.016414f
C402 VTAIL.n343 B 0.00882f
C403 VTAIL.n344 B 0.020848f
C404 VTAIL.n345 B 0.009339f
C405 VTAIL.n346 B 0.016414f
C406 VTAIL.n347 B 0.00882f
C407 VTAIL.n348 B 0.020848f
C408 VTAIL.n349 B 0.009339f
C409 VTAIL.n350 B 0.016414f
C410 VTAIL.n351 B 0.00882f
C411 VTAIL.n352 B 0.020848f
C412 VTAIL.n353 B 0.009339f
C413 VTAIL.n354 B 0.106399f
C414 VTAIL.t6 B 0.034367f
C415 VTAIL.n355 B 0.015636f
C416 VTAIL.n356 B 0.012316f
C417 VTAIL.n357 B 0.00882f
C418 VTAIL.n358 B 1.0559f
C419 VTAIL.n359 B 0.016414f
C420 VTAIL.n360 B 0.00882f
C421 VTAIL.n361 B 0.009339f
C422 VTAIL.n362 B 0.020848f
C423 VTAIL.n363 B 0.020848f
C424 VTAIL.n364 B 0.009339f
C425 VTAIL.n365 B 0.00882f
C426 VTAIL.n366 B 0.016414f
C427 VTAIL.n367 B 0.016414f
C428 VTAIL.n368 B 0.00882f
C429 VTAIL.n369 B 0.009339f
C430 VTAIL.n370 B 0.020848f
C431 VTAIL.n371 B 0.020848f
C432 VTAIL.n372 B 0.009339f
C433 VTAIL.n373 B 0.00882f
C434 VTAIL.n374 B 0.016414f
C435 VTAIL.n375 B 0.016414f
C436 VTAIL.n376 B 0.00882f
C437 VTAIL.n377 B 0.009339f
C438 VTAIL.n378 B 0.020848f
C439 VTAIL.n379 B 0.020848f
C440 VTAIL.n380 B 0.009339f
C441 VTAIL.n381 B 0.00882f
C442 VTAIL.n382 B 0.016414f
C443 VTAIL.n383 B 0.016414f
C444 VTAIL.n384 B 0.00882f
C445 VTAIL.n385 B 0.009339f
C446 VTAIL.n386 B 0.020848f
C447 VTAIL.n387 B 0.020848f
C448 VTAIL.n388 B 0.009339f
C449 VTAIL.n389 B 0.00882f
C450 VTAIL.n390 B 0.016414f
C451 VTAIL.n391 B 0.016414f
C452 VTAIL.n392 B 0.00882f
C453 VTAIL.n393 B 0.009339f
C454 VTAIL.n394 B 0.020848f
C455 VTAIL.n395 B 0.020848f
C456 VTAIL.n396 B 0.009339f
C457 VTAIL.n397 B 0.00882f
C458 VTAIL.n398 B 0.016414f
C459 VTAIL.n399 B 0.016414f
C460 VTAIL.n400 B 0.00882f
C461 VTAIL.n401 B 0.00908f
C462 VTAIL.n402 B 0.00908f
C463 VTAIL.n403 B 0.020848f
C464 VTAIL.n404 B 0.045133f
C465 VTAIL.n405 B 0.009339f
C466 VTAIL.n406 B 0.00882f
C467 VTAIL.n407 B 0.042426f
C468 VTAIL.n408 B 0.025385f
C469 VTAIL.n409 B 0.224244f
C470 VTAIL.n410 B 0.023072f
C471 VTAIL.n411 B 0.016414f
C472 VTAIL.n412 B 0.00882f
C473 VTAIL.n413 B 0.020848f
C474 VTAIL.n414 B 0.009339f
C475 VTAIL.n415 B 0.016414f
C476 VTAIL.n416 B 0.00882f
C477 VTAIL.n417 B 0.020848f
C478 VTAIL.n418 B 0.020848f
C479 VTAIL.n419 B 0.009339f
C480 VTAIL.n420 B 0.016414f
C481 VTAIL.n421 B 0.00882f
C482 VTAIL.n422 B 0.020848f
C483 VTAIL.n423 B 0.009339f
C484 VTAIL.n424 B 0.016414f
C485 VTAIL.n425 B 0.00882f
C486 VTAIL.n426 B 0.020848f
C487 VTAIL.n427 B 0.009339f
C488 VTAIL.n428 B 0.016414f
C489 VTAIL.n429 B 0.00882f
C490 VTAIL.n430 B 0.020848f
C491 VTAIL.n431 B 0.009339f
C492 VTAIL.n432 B 0.016414f
C493 VTAIL.n433 B 0.00882f
C494 VTAIL.n434 B 0.020848f
C495 VTAIL.n435 B 0.009339f
C496 VTAIL.n436 B 0.106399f
C497 VTAIL.t2 B 0.034367f
C498 VTAIL.n437 B 0.015636f
C499 VTAIL.n438 B 0.012316f
C500 VTAIL.n439 B 0.00882f
C501 VTAIL.n440 B 1.0559f
C502 VTAIL.n441 B 0.016414f
C503 VTAIL.n442 B 0.00882f
C504 VTAIL.n443 B 0.009339f
C505 VTAIL.n444 B 0.020848f
C506 VTAIL.n445 B 0.020848f
C507 VTAIL.n446 B 0.009339f
C508 VTAIL.n447 B 0.00882f
C509 VTAIL.n448 B 0.016414f
C510 VTAIL.n449 B 0.016414f
C511 VTAIL.n450 B 0.00882f
C512 VTAIL.n451 B 0.009339f
C513 VTAIL.n452 B 0.020848f
C514 VTAIL.n453 B 0.020848f
C515 VTAIL.n454 B 0.009339f
C516 VTAIL.n455 B 0.00882f
C517 VTAIL.n456 B 0.016414f
C518 VTAIL.n457 B 0.016414f
C519 VTAIL.n458 B 0.00882f
C520 VTAIL.n459 B 0.009339f
C521 VTAIL.n460 B 0.020848f
C522 VTAIL.n461 B 0.020848f
C523 VTAIL.n462 B 0.009339f
C524 VTAIL.n463 B 0.00882f
C525 VTAIL.n464 B 0.016414f
C526 VTAIL.n465 B 0.016414f
C527 VTAIL.n466 B 0.00882f
C528 VTAIL.n467 B 0.009339f
C529 VTAIL.n468 B 0.020848f
C530 VTAIL.n469 B 0.020848f
C531 VTAIL.n470 B 0.009339f
C532 VTAIL.n471 B 0.00882f
C533 VTAIL.n472 B 0.016414f
C534 VTAIL.n473 B 0.016414f
C535 VTAIL.n474 B 0.00882f
C536 VTAIL.n475 B 0.009339f
C537 VTAIL.n476 B 0.020848f
C538 VTAIL.n477 B 0.020848f
C539 VTAIL.n478 B 0.009339f
C540 VTAIL.n479 B 0.00882f
C541 VTAIL.n480 B 0.016414f
C542 VTAIL.n481 B 0.016414f
C543 VTAIL.n482 B 0.00882f
C544 VTAIL.n483 B 0.00908f
C545 VTAIL.n484 B 0.00908f
C546 VTAIL.n485 B 0.020848f
C547 VTAIL.n486 B 0.045133f
C548 VTAIL.n487 B 0.009339f
C549 VTAIL.n488 B 0.00882f
C550 VTAIL.n489 B 0.042426f
C551 VTAIL.n490 B 0.025385f
C552 VTAIL.n491 B 0.224244f
C553 VTAIL.n492 B 0.023072f
C554 VTAIL.n493 B 0.016414f
C555 VTAIL.n494 B 0.00882f
C556 VTAIL.n495 B 0.020848f
C557 VTAIL.n496 B 0.009339f
C558 VTAIL.n497 B 0.016414f
C559 VTAIL.n498 B 0.00882f
C560 VTAIL.n499 B 0.020848f
C561 VTAIL.n500 B 0.020848f
C562 VTAIL.n501 B 0.009339f
C563 VTAIL.n502 B 0.016414f
C564 VTAIL.n503 B 0.00882f
C565 VTAIL.n504 B 0.020848f
C566 VTAIL.n505 B 0.009339f
C567 VTAIL.n506 B 0.016414f
C568 VTAIL.n507 B 0.00882f
C569 VTAIL.n508 B 0.020848f
C570 VTAIL.n509 B 0.009339f
C571 VTAIL.n510 B 0.016414f
C572 VTAIL.n511 B 0.00882f
C573 VTAIL.n512 B 0.020848f
C574 VTAIL.n513 B 0.009339f
C575 VTAIL.n514 B 0.016414f
C576 VTAIL.n515 B 0.00882f
C577 VTAIL.n516 B 0.020848f
C578 VTAIL.n517 B 0.009339f
C579 VTAIL.n518 B 0.106399f
C580 VTAIL.t0 B 0.034367f
C581 VTAIL.n519 B 0.015636f
C582 VTAIL.n520 B 0.012316f
C583 VTAIL.n521 B 0.00882f
C584 VTAIL.n522 B 1.0559f
C585 VTAIL.n523 B 0.016414f
C586 VTAIL.n524 B 0.00882f
C587 VTAIL.n525 B 0.009339f
C588 VTAIL.n526 B 0.020848f
C589 VTAIL.n527 B 0.020848f
C590 VTAIL.n528 B 0.009339f
C591 VTAIL.n529 B 0.00882f
C592 VTAIL.n530 B 0.016414f
C593 VTAIL.n531 B 0.016414f
C594 VTAIL.n532 B 0.00882f
C595 VTAIL.n533 B 0.009339f
C596 VTAIL.n534 B 0.020848f
C597 VTAIL.n535 B 0.020848f
C598 VTAIL.n536 B 0.009339f
C599 VTAIL.n537 B 0.00882f
C600 VTAIL.n538 B 0.016414f
C601 VTAIL.n539 B 0.016414f
C602 VTAIL.n540 B 0.00882f
C603 VTAIL.n541 B 0.009339f
C604 VTAIL.n542 B 0.020848f
C605 VTAIL.n543 B 0.020848f
C606 VTAIL.n544 B 0.009339f
C607 VTAIL.n545 B 0.00882f
C608 VTAIL.n546 B 0.016414f
C609 VTAIL.n547 B 0.016414f
C610 VTAIL.n548 B 0.00882f
C611 VTAIL.n549 B 0.009339f
C612 VTAIL.n550 B 0.020848f
C613 VTAIL.n551 B 0.020848f
C614 VTAIL.n552 B 0.009339f
C615 VTAIL.n553 B 0.00882f
C616 VTAIL.n554 B 0.016414f
C617 VTAIL.n555 B 0.016414f
C618 VTAIL.n556 B 0.00882f
C619 VTAIL.n557 B 0.009339f
C620 VTAIL.n558 B 0.020848f
C621 VTAIL.n559 B 0.020848f
C622 VTAIL.n560 B 0.009339f
C623 VTAIL.n561 B 0.00882f
C624 VTAIL.n562 B 0.016414f
C625 VTAIL.n563 B 0.016414f
C626 VTAIL.n564 B 0.00882f
C627 VTAIL.n565 B 0.00908f
C628 VTAIL.n566 B 0.00908f
C629 VTAIL.n567 B 0.020848f
C630 VTAIL.n568 B 0.045133f
C631 VTAIL.n569 B 0.009339f
C632 VTAIL.n570 B 0.00882f
C633 VTAIL.n571 B 0.042426f
C634 VTAIL.n572 B 0.025385f
C635 VTAIL.n573 B 1.28184f
C636 VTAIL.n574 B 0.023072f
C637 VTAIL.n575 B 0.016414f
C638 VTAIL.n576 B 0.00882f
C639 VTAIL.n577 B 0.020848f
C640 VTAIL.n578 B 0.009339f
C641 VTAIL.n579 B 0.016414f
C642 VTAIL.n580 B 0.00882f
C643 VTAIL.n581 B 0.020848f
C644 VTAIL.n582 B 0.009339f
C645 VTAIL.n583 B 0.016414f
C646 VTAIL.n584 B 0.00882f
C647 VTAIL.n585 B 0.020848f
C648 VTAIL.n586 B 0.009339f
C649 VTAIL.n587 B 0.016414f
C650 VTAIL.n588 B 0.00882f
C651 VTAIL.n589 B 0.020848f
C652 VTAIL.n590 B 0.009339f
C653 VTAIL.n591 B 0.016414f
C654 VTAIL.n592 B 0.00882f
C655 VTAIL.n593 B 0.020848f
C656 VTAIL.n594 B 0.009339f
C657 VTAIL.n595 B 0.016414f
C658 VTAIL.n596 B 0.00882f
C659 VTAIL.n597 B 0.020848f
C660 VTAIL.n598 B 0.009339f
C661 VTAIL.n599 B 0.106399f
C662 VTAIL.t4 B 0.034367f
C663 VTAIL.n600 B 0.015636f
C664 VTAIL.n601 B 0.012316f
C665 VTAIL.n602 B 0.00882f
C666 VTAIL.n603 B 1.0559f
C667 VTAIL.n604 B 0.016414f
C668 VTAIL.n605 B 0.00882f
C669 VTAIL.n606 B 0.009339f
C670 VTAIL.n607 B 0.020848f
C671 VTAIL.n608 B 0.020848f
C672 VTAIL.n609 B 0.009339f
C673 VTAIL.n610 B 0.00882f
C674 VTAIL.n611 B 0.016414f
C675 VTAIL.n612 B 0.016414f
C676 VTAIL.n613 B 0.00882f
C677 VTAIL.n614 B 0.009339f
C678 VTAIL.n615 B 0.020848f
C679 VTAIL.n616 B 0.020848f
C680 VTAIL.n617 B 0.009339f
C681 VTAIL.n618 B 0.00882f
C682 VTAIL.n619 B 0.016414f
C683 VTAIL.n620 B 0.016414f
C684 VTAIL.n621 B 0.00882f
C685 VTAIL.n622 B 0.009339f
C686 VTAIL.n623 B 0.020848f
C687 VTAIL.n624 B 0.020848f
C688 VTAIL.n625 B 0.009339f
C689 VTAIL.n626 B 0.00882f
C690 VTAIL.n627 B 0.016414f
C691 VTAIL.n628 B 0.016414f
C692 VTAIL.n629 B 0.00882f
C693 VTAIL.n630 B 0.009339f
C694 VTAIL.n631 B 0.020848f
C695 VTAIL.n632 B 0.020848f
C696 VTAIL.n633 B 0.009339f
C697 VTAIL.n634 B 0.00882f
C698 VTAIL.n635 B 0.016414f
C699 VTAIL.n636 B 0.016414f
C700 VTAIL.n637 B 0.00882f
C701 VTAIL.n638 B 0.009339f
C702 VTAIL.n639 B 0.020848f
C703 VTAIL.n640 B 0.020848f
C704 VTAIL.n641 B 0.020848f
C705 VTAIL.n642 B 0.009339f
C706 VTAIL.n643 B 0.00882f
C707 VTAIL.n644 B 0.016414f
C708 VTAIL.n645 B 0.016414f
C709 VTAIL.n646 B 0.00882f
C710 VTAIL.n647 B 0.00908f
C711 VTAIL.n648 B 0.00908f
C712 VTAIL.n649 B 0.020848f
C713 VTAIL.n650 B 0.045133f
C714 VTAIL.n651 B 0.009339f
C715 VTAIL.n652 B 0.00882f
C716 VTAIL.n653 B 0.042426f
C717 VTAIL.n654 B 0.025385f
C718 VTAIL.n655 B 1.18734f
C719 VN.t0 B 3.22972f
C720 VN.t1 B 3.24123f
C721 VN.n0 B 1.9766f
C722 VN.t2 B 3.22972f
C723 VN.t3 B 3.24123f
C724 VN.n1 B 3.32183f
.ends

