* NGSPICE file created from diff_pair_sample_1449.ext - technology: sky130A

.subckt diff_pair_sample_1449 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=0 ps=0 w=5.28 l=1.23
X1 B.t8 B.t6 B.t7 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=0 ps=0 w=5.28 l=1.23
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=2.0592 ps=11.34 w=5.28 l=1.23
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=2.0592 ps=11.34 w=5.28 l=1.23
X4 B.t5 B.t3 B.t4 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=0 ps=0 w=5.28 l=1.23
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=2.0592 ps=11.34 w=5.28 l=1.23
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=2.0592 ps=11.34 w=5.28 l=1.23
X7 B.t2 B.t0 B.t1 w_n1594_n2024# sky130_fd_pr__pfet_01v8 ad=2.0592 pd=11.34 as=0 ps=0 w=5.28 l=1.23
R0 B.n203 B.n202 585
R1 B.n201 B.n60 585
R2 B.n200 B.n199 585
R3 B.n198 B.n61 585
R4 B.n197 B.n196 585
R5 B.n195 B.n62 585
R6 B.n194 B.n193 585
R7 B.n192 B.n63 585
R8 B.n191 B.n190 585
R9 B.n189 B.n64 585
R10 B.n188 B.n187 585
R11 B.n186 B.n65 585
R12 B.n185 B.n184 585
R13 B.n183 B.n66 585
R14 B.n182 B.n181 585
R15 B.n180 B.n67 585
R16 B.n179 B.n178 585
R17 B.n177 B.n68 585
R18 B.n176 B.n175 585
R19 B.n174 B.n69 585
R20 B.n173 B.n172 585
R21 B.n171 B.n70 585
R22 B.n170 B.n169 585
R23 B.n165 B.n71 585
R24 B.n164 B.n163 585
R25 B.n162 B.n72 585
R26 B.n161 B.n160 585
R27 B.n159 B.n73 585
R28 B.n158 B.n157 585
R29 B.n156 B.n74 585
R30 B.n155 B.n154 585
R31 B.n152 B.n75 585
R32 B.n151 B.n150 585
R33 B.n149 B.n78 585
R34 B.n148 B.n147 585
R35 B.n146 B.n79 585
R36 B.n145 B.n144 585
R37 B.n143 B.n80 585
R38 B.n142 B.n141 585
R39 B.n140 B.n81 585
R40 B.n139 B.n138 585
R41 B.n137 B.n82 585
R42 B.n136 B.n135 585
R43 B.n134 B.n83 585
R44 B.n133 B.n132 585
R45 B.n131 B.n84 585
R46 B.n130 B.n129 585
R47 B.n128 B.n85 585
R48 B.n127 B.n126 585
R49 B.n125 B.n86 585
R50 B.n124 B.n123 585
R51 B.n122 B.n87 585
R52 B.n121 B.n120 585
R53 B.n204 B.n59 585
R54 B.n206 B.n205 585
R55 B.n207 B.n58 585
R56 B.n209 B.n208 585
R57 B.n210 B.n57 585
R58 B.n212 B.n211 585
R59 B.n213 B.n56 585
R60 B.n215 B.n214 585
R61 B.n216 B.n55 585
R62 B.n218 B.n217 585
R63 B.n219 B.n54 585
R64 B.n221 B.n220 585
R65 B.n222 B.n53 585
R66 B.n224 B.n223 585
R67 B.n225 B.n52 585
R68 B.n227 B.n226 585
R69 B.n228 B.n51 585
R70 B.n230 B.n229 585
R71 B.n231 B.n50 585
R72 B.n233 B.n232 585
R73 B.n234 B.n49 585
R74 B.n236 B.n235 585
R75 B.n237 B.n48 585
R76 B.n239 B.n238 585
R77 B.n240 B.n47 585
R78 B.n242 B.n241 585
R79 B.n243 B.n46 585
R80 B.n245 B.n244 585
R81 B.n246 B.n45 585
R82 B.n248 B.n247 585
R83 B.n249 B.n44 585
R84 B.n251 B.n250 585
R85 B.n252 B.n43 585
R86 B.n254 B.n253 585
R87 B.n255 B.n42 585
R88 B.n257 B.n256 585
R89 B.n338 B.n337 585
R90 B.n336 B.n11 585
R91 B.n335 B.n334 585
R92 B.n333 B.n12 585
R93 B.n332 B.n331 585
R94 B.n330 B.n13 585
R95 B.n329 B.n328 585
R96 B.n327 B.n14 585
R97 B.n326 B.n325 585
R98 B.n324 B.n15 585
R99 B.n323 B.n322 585
R100 B.n321 B.n16 585
R101 B.n320 B.n319 585
R102 B.n318 B.n17 585
R103 B.n317 B.n316 585
R104 B.n315 B.n18 585
R105 B.n314 B.n313 585
R106 B.n312 B.n19 585
R107 B.n311 B.n310 585
R108 B.n309 B.n20 585
R109 B.n308 B.n307 585
R110 B.n306 B.n21 585
R111 B.n304 B.n303 585
R112 B.n302 B.n24 585
R113 B.n301 B.n300 585
R114 B.n299 B.n25 585
R115 B.n298 B.n297 585
R116 B.n296 B.n26 585
R117 B.n295 B.n294 585
R118 B.n293 B.n27 585
R119 B.n292 B.n291 585
R120 B.n290 B.n289 585
R121 B.n288 B.n31 585
R122 B.n287 B.n286 585
R123 B.n285 B.n32 585
R124 B.n284 B.n283 585
R125 B.n282 B.n33 585
R126 B.n281 B.n280 585
R127 B.n279 B.n34 585
R128 B.n278 B.n277 585
R129 B.n276 B.n35 585
R130 B.n275 B.n274 585
R131 B.n273 B.n36 585
R132 B.n272 B.n271 585
R133 B.n270 B.n37 585
R134 B.n269 B.n268 585
R135 B.n267 B.n38 585
R136 B.n266 B.n265 585
R137 B.n264 B.n39 585
R138 B.n263 B.n262 585
R139 B.n261 B.n40 585
R140 B.n260 B.n259 585
R141 B.n258 B.n41 585
R142 B.n339 B.n10 585
R143 B.n341 B.n340 585
R144 B.n342 B.n9 585
R145 B.n344 B.n343 585
R146 B.n345 B.n8 585
R147 B.n347 B.n346 585
R148 B.n348 B.n7 585
R149 B.n350 B.n349 585
R150 B.n351 B.n6 585
R151 B.n353 B.n352 585
R152 B.n354 B.n5 585
R153 B.n356 B.n355 585
R154 B.n357 B.n4 585
R155 B.n359 B.n358 585
R156 B.n360 B.n3 585
R157 B.n362 B.n361 585
R158 B.n363 B.n0 585
R159 B.n2 B.n1 585
R160 B.n97 B.n96 585
R161 B.n98 B.n95 585
R162 B.n100 B.n99 585
R163 B.n101 B.n94 585
R164 B.n103 B.n102 585
R165 B.n104 B.n93 585
R166 B.n106 B.n105 585
R167 B.n107 B.n92 585
R168 B.n109 B.n108 585
R169 B.n110 B.n91 585
R170 B.n112 B.n111 585
R171 B.n113 B.n90 585
R172 B.n115 B.n114 585
R173 B.n116 B.n89 585
R174 B.n118 B.n117 585
R175 B.n119 B.n88 585
R176 B.n120 B.n119 487.695
R177 B.n202 B.n59 487.695
R178 B.n256 B.n41 487.695
R179 B.n339 B.n338 487.695
R180 B.n76 B.t3 307.724
R181 B.n166 B.t0 307.724
R182 B.n28 B.t6 307.724
R183 B.n22 B.t9 307.724
R184 B.n166 B.t1 285.902
R185 B.n28 B.t8 285.902
R186 B.n76 B.t4 285.902
R187 B.n22 B.t11 285.902
R188 B.n365 B.n364 256.663
R189 B.n167 B.t2 255.649
R190 B.n29 B.t7 255.649
R191 B.n77 B.t5 255.649
R192 B.n23 B.t10 255.649
R193 B.n364 B.n363 235.042
R194 B.n364 B.n2 235.042
R195 B.n120 B.n87 163.367
R196 B.n124 B.n87 163.367
R197 B.n125 B.n124 163.367
R198 B.n126 B.n125 163.367
R199 B.n126 B.n85 163.367
R200 B.n130 B.n85 163.367
R201 B.n131 B.n130 163.367
R202 B.n132 B.n131 163.367
R203 B.n132 B.n83 163.367
R204 B.n136 B.n83 163.367
R205 B.n137 B.n136 163.367
R206 B.n138 B.n137 163.367
R207 B.n138 B.n81 163.367
R208 B.n142 B.n81 163.367
R209 B.n143 B.n142 163.367
R210 B.n144 B.n143 163.367
R211 B.n144 B.n79 163.367
R212 B.n148 B.n79 163.367
R213 B.n149 B.n148 163.367
R214 B.n150 B.n149 163.367
R215 B.n150 B.n75 163.367
R216 B.n155 B.n75 163.367
R217 B.n156 B.n155 163.367
R218 B.n157 B.n156 163.367
R219 B.n157 B.n73 163.367
R220 B.n161 B.n73 163.367
R221 B.n162 B.n161 163.367
R222 B.n163 B.n162 163.367
R223 B.n163 B.n71 163.367
R224 B.n170 B.n71 163.367
R225 B.n171 B.n170 163.367
R226 B.n172 B.n171 163.367
R227 B.n172 B.n69 163.367
R228 B.n176 B.n69 163.367
R229 B.n177 B.n176 163.367
R230 B.n178 B.n177 163.367
R231 B.n178 B.n67 163.367
R232 B.n182 B.n67 163.367
R233 B.n183 B.n182 163.367
R234 B.n184 B.n183 163.367
R235 B.n184 B.n65 163.367
R236 B.n188 B.n65 163.367
R237 B.n189 B.n188 163.367
R238 B.n190 B.n189 163.367
R239 B.n190 B.n63 163.367
R240 B.n194 B.n63 163.367
R241 B.n195 B.n194 163.367
R242 B.n196 B.n195 163.367
R243 B.n196 B.n61 163.367
R244 B.n200 B.n61 163.367
R245 B.n201 B.n200 163.367
R246 B.n202 B.n201 163.367
R247 B.n256 B.n255 163.367
R248 B.n255 B.n254 163.367
R249 B.n254 B.n43 163.367
R250 B.n250 B.n43 163.367
R251 B.n250 B.n249 163.367
R252 B.n249 B.n248 163.367
R253 B.n248 B.n45 163.367
R254 B.n244 B.n45 163.367
R255 B.n244 B.n243 163.367
R256 B.n243 B.n242 163.367
R257 B.n242 B.n47 163.367
R258 B.n238 B.n47 163.367
R259 B.n238 B.n237 163.367
R260 B.n237 B.n236 163.367
R261 B.n236 B.n49 163.367
R262 B.n232 B.n49 163.367
R263 B.n232 B.n231 163.367
R264 B.n231 B.n230 163.367
R265 B.n230 B.n51 163.367
R266 B.n226 B.n51 163.367
R267 B.n226 B.n225 163.367
R268 B.n225 B.n224 163.367
R269 B.n224 B.n53 163.367
R270 B.n220 B.n53 163.367
R271 B.n220 B.n219 163.367
R272 B.n219 B.n218 163.367
R273 B.n218 B.n55 163.367
R274 B.n214 B.n55 163.367
R275 B.n214 B.n213 163.367
R276 B.n213 B.n212 163.367
R277 B.n212 B.n57 163.367
R278 B.n208 B.n57 163.367
R279 B.n208 B.n207 163.367
R280 B.n207 B.n206 163.367
R281 B.n206 B.n59 163.367
R282 B.n338 B.n11 163.367
R283 B.n334 B.n11 163.367
R284 B.n334 B.n333 163.367
R285 B.n333 B.n332 163.367
R286 B.n332 B.n13 163.367
R287 B.n328 B.n13 163.367
R288 B.n328 B.n327 163.367
R289 B.n327 B.n326 163.367
R290 B.n326 B.n15 163.367
R291 B.n322 B.n15 163.367
R292 B.n322 B.n321 163.367
R293 B.n321 B.n320 163.367
R294 B.n320 B.n17 163.367
R295 B.n316 B.n17 163.367
R296 B.n316 B.n315 163.367
R297 B.n315 B.n314 163.367
R298 B.n314 B.n19 163.367
R299 B.n310 B.n19 163.367
R300 B.n310 B.n309 163.367
R301 B.n309 B.n308 163.367
R302 B.n308 B.n21 163.367
R303 B.n303 B.n21 163.367
R304 B.n303 B.n302 163.367
R305 B.n302 B.n301 163.367
R306 B.n301 B.n25 163.367
R307 B.n297 B.n25 163.367
R308 B.n297 B.n296 163.367
R309 B.n296 B.n295 163.367
R310 B.n295 B.n27 163.367
R311 B.n291 B.n27 163.367
R312 B.n291 B.n290 163.367
R313 B.n290 B.n31 163.367
R314 B.n286 B.n31 163.367
R315 B.n286 B.n285 163.367
R316 B.n285 B.n284 163.367
R317 B.n284 B.n33 163.367
R318 B.n280 B.n33 163.367
R319 B.n280 B.n279 163.367
R320 B.n279 B.n278 163.367
R321 B.n278 B.n35 163.367
R322 B.n274 B.n35 163.367
R323 B.n274 B.n273 163.367
R324 B.n273 B.n272 163.367
R325 B.n272 B.n37 163.367
R326 B.n268 B.n37 163.367
R327 B.n268 B.n267 163.367
R328 B.n267 B.n266 163.367
R329 B.n266 B.n39 163.367
R330 B.n262 B.n39 163.367
R331 B.n262 B.n261 163.367
R332 B.n261 B.n260 163.367
R333 B.n260 B.n41 163.367
R334 B.n340 B.n339 163.367
R335 B.n340 B.n9 163.367
R336 B.n344 B.n9 163.367
R337 B.n345 B.n344 163.367
R338 B.n346 B.n345 163.367
R339 B.n346 B.n7 163.367
R340 B.n350 B.n7 163.367
R341 B.n351 B.n350 163.367
R342 B.n352 B.n351 163.367
R343 B.n352 B.n5 163.367
R344 B.n356 B.n5 163.367
R345 B.n357 B.n356 163.367
R346 B.n358 B.n357 163.367
R347 B.n358 B.n3 163.367
R348 B.n362 B.n3 163.367
R349 B.n363 B.n362 163.367
R350 B.n96 B.n2 163.367
R351 B.n96 B.n95 163.367
R352 B.n100 B.n95 163.367
R353 B.n101 B.n100 163.367
R354 B.n102 B.n101 163.367
R355 B.n102 B.n93 163.367
R356 B.n106 B.n93 163.367
R357 B.n107 B.n106 163.367
R358 B.n108 B.n107 163.367
R359 B.n108 B.n91 163.367
R360 B.n112 B.n91 163.367
R361 B.n113 B.n112 163.367
R362 B.n114 B.n113 163.367
R363 B.n114 B.n89 163.367
R364 B.n118 B.n89 163.367
R365 B.n119 B.n118 163.367
R366 B.n153 B.n77 59.5399
R367 B.n168 B.n167 59.5399
R368 B.n30 B.n29 59.5399
R369 B.n305 B.n23 59.5399
R370 B.n337 B.n10 31.6883
R371 B.n258 B.n257 31.6883
R372 B.n204 B.n203 31.6883
R373 B.n121 B.n88 31.6883
R374 B.n77 B.n76 30.255
R375 B.n167 B.n166 30.255
R376 B.n29 B.n28 30.255
R377 B.n23 B.n22 30.255
R378 B B.n365 18.0485
R379 B.n341 B.n10 10.6151
R380 B.n342 B.n341 10.6151
R381 B.n343 B.n342 10.6151
R382 B.n343 B.n8 10.6151
R383 B.n347 B.n8 10.6151
R384 B.n348 B.n347 10.6151
R385 B.n349 B.n348 10.6151
R386 B.n349 B.n6 10.6151
R387 B.n353 B.n6 10.6151
R388 B.n354 B.n353 10.6151
R389 B.n355 B.n354 10.6151
R390 B.n355 B.n4 10.6151
R391 B.n359 B.n4 10.6151
R392 B.n360 B.n359 10.6151
R393 B.n361 B.n360 10.6151
R394 B.n361 B.n0 10.6151
R395 B.n337 B.n336 10.6151
R396 B.n336 B.n335 10.6151
R397 B.n335 B.n12 10.6151
R398 B.n331 B.n12 10.6151
R399 B.n331 B.n330 10.6151
R400 B.n330 B.n329 10.6151
R401 B.n329 B.n14 10.6151
R402 B.n325 B.n14 10.6151
R403 B.n325 B.n324 10.6151
R404 B.n324 B.n323 10.6151
R405 B.n323 B.n16 10.6151
R406 B.n319 B.n16 10.6151
R407 B.n319 B.n318 10.6151
R408 B.n318 B.n317 10.6151
R409 B.n317 B.n18 10.6151
R410 B.n313 B.n18 10.6151
R411 B.n313 B.n312 10.6151
R412 B.n312 B.n311 10.6151
R413 B.n311 B.n20 10.6151
R414 B.n307 B.n20 10.6151
R415 B.n307 B.n306 10.6151
R416 B.n304 B.n24 10.6151
R417 B.n300 B.n24 10.6151
R418 B.n300 B.n299 10.6151
R419 B.n299 B.n298 10.6151
R420 B.n298 B.n26 10.6151
R421 B.n294 B.n26 10.6151
R422 B.n294 B.n293 10.6151
R423 B.n293 B.n292 10.6151
R424 B.n289 B.n288 10.6151
R425 B.n288 B.n287 10.6151
R426 B.n287 B.n32 10.6151
R427 B.n283 B.n32 10.6151
R428 B.n283 B.n282 10.6151
R429 B.n282 B.n281 10.6151
R430 B.n281 B.n34 10.6151
R431 B.n277 B.n34 10.6151
R432 B.n277 B.n276 10.6151
R433 B.n276 B.n275 10.6151
R434 B.n275 B.n36 10.6151
R435 B.n271 B.n36 10.6151
R436 B.n271 B.n270 10.6151
R437 B.n270 B.n269 10.6151
R438 B.n269 B.n38 10.6151
R439 B.n265 B.n38 10.6151
R440 B.n265 B.n264 10.6151
R441 B.n264 B.n263 10.6151
R442 B.n263 B.n40 10.6151
R443 B.n259 B.n40 10.6151
R444 B.n259 B.n258 10.6151
R445 B.n257 B.n42 10.6151
R446 B.n253 B.n42 10.6151
R447 B.n253 B.n252 10.6151
R448 B.n252 B.n251 10.6151
R449 B.n251 B.n44 10.6151
R450 B.n247 B.n44 10.6151
R451 B.n247 B.n246 10.6151
R452 B.n246 B.n245 10.6151
R453 B.n245 B.n46 10.6151
R454 B.n241 B.n46 10.6151
R455 B.n241 B.n240 10.6151
R456 B.n240 B.n239 10.6151
R457 B.n239 B.n48 10.6151
R458 B.n235 B.n48 10.6151
R459 B.n235 B.n234 10.6151
R460 B.n234 B.n233 10.6151
R461 B.n233 B.n50 10.6151
R462 B.n229 B.n50 10.6151
R463 B.n229 B.n228 10.6151
R464 B.n228 B.n227 10.6151
R465 B.n227 B.n52 10.6151
R466 B.n223 B.n52 10.6151
R467 B.n223 B.n222 10.6151
R468 B.n222 B.n221 10.6151
R469 B.n221 B.n54 10.6151
R470 B.n217 B.n54 10.6151
R471 B.n217 B.n216 10.6151
R472 B.n216 B.n215 10.6151
R473 B.n215 B.n56 10.6151
R474 B.n211 B.n56 10.6151
R475 B.n211 B.n210 10.6151
R476 B.n210 B.n209 10.6151
R477 B.n209 B.n58 10.6151
R478 B.n205 B.n58 10.6151
R479 B.n205 B.n204 10.6151
R480 B.n97 B.n1 10.6151
R481 B.n98 B.n97 10.6151
R482 B.n99 B.n98 10.6151
R483 B.n99 B.n94 10.6151
R484 B.n103 B.n94 10.6151
R485 B.n104 B.n103 10.6151
R486 B.n105 B.n104 10.6151
R487 B.n105 B.n92 10.6151
R488 B.n109 B.n92 10.6151
R489 B.n110 B.n109 10.6151
R490 B.n111 B.n110 10.6151
R491 B.n111 B.n90 10.6151
R492 B.n115 B.n90 10.6151
R493 B.n116 B.n115 10.6151
R494 B.n117 B.n116 10.6151
R495 B.n117 B.n88 10.6151
R496 B.n122 B.n121 10.6151
R497 B.n123 B.n122 10.6151
R498 B.n123 B.n86 10.6151
R499 B.n127 B.n86 10.6151
R500 B.n128 B.n127 10.6151
R501 B.n129 B.n128 10.6151
R502 B.n129 B.n84 10.6151
R503 B.n133 B.n84 10.6151
R504 B.n134 B.n133 10.6151
R505 B.n135 B.n134 10.6151
R506 B.n135 B.n82 10.6151
R507 B.n139 B.n82 10.6151
R508 B.n140 B.n139 10.6151
R509 B.n141 B.n140 10.6151
R510 B.n141 B.n80 10.6151
R511 B.n145 B.n80 10.6151
R512 B.n146 B.n145 10.6151
R513 B.n147 B.n146 10.6151
R514 B.n147 B.n78 10.6151
R515 B.n151 B.n78 10.6151
R516 B.n152 B.n151 10.6151
R517 B.n154 B.n74 10.6151
R518 B.n158 B.n74 10.6151
R519 B.n159 B.n158 10.6151
R520 B.n160 B.n159 10.6151
R521 B.n160 B.n72 10.6151
R522 B.n164 B.n72 10.6151
R523 B.n165 B.n164 10.6151
R524 B.n169 B.n165 10.6151
R525 B.n173 B.n70 10.6151
R526 B.n174 B.n173 10.6151
R527 B.n175 B.n174 10.6151
R528 B.n175 B.n68 10.6151
R529 B.n179 B.n68 10.6151
R530 B.n180 B.n179 10.6151
R531 B.n181 B.n180 10.6151
R532 B.n181 B.n66 10.6151
R533 B.n185 B.n66 10.6151
R534 B.n186 B.n185 10.6151
R535 B.n187 B.n186 10.6151
R536 B.n187 B.n64 10.6151
R537 B.n191 B.n64 10.6151
R538 B.n192 B.n191 10.6151
R539 B.n193 B.n192 10.6151
R540 B.n193 B.n62 10.6151
R541 B.n197 B.n62 10.6151
R542 B.n198 B.n197 10.6151
R543 B.n199 B.n198 10.6151
R544 B.n199 B.n60 10.6151
R545 B.n203 B.n60 10.6151
R546 B.n365 B.n0 8.11757
R547 B.n365 B.n1 8.11757
R548 B.n305 B.n304 6.5566
R549 B.n292 B.n30 6.5566
R550 B.n154 B.n153 6.5566
R551 B.n169 B.n168 6.5566
R552 B.n306 B.n305 4.05904
R553 B.n289 B.n30 4.05904
R554 B.n153 B.n152 4.05904
R555 B.n168 B.n70 4.05904
R556 VN VN.t0 252.213
R557 VN VN.t1 216.142
R558 VTAIL.n106 VTAIL.n84 756.745
R559 VTAIL.n22 VTAIL.n0 756.745
R560 VTAIL.n78 VTAIL.n56 756.745
R561 VTAIL.n50 VTAIL.n28 756.745
R562 VTAIL.n92 VTAIL.n91 585
R563 VTAIL.n97 VTAIL.n96 585
R564 VTAIL.n99 VTAIL.n98 585
R565 VTAIL.n88 VTAIL.n87 585
R566 VTAIL.n105 VTAIL.n104 585
R567 VTAIL.n107 VTAIL.n106 585
R568 VTAIL.n8 VTAIL.n7 585
R569 VTAIL.n13 VTAIL.n12 585
R570 VTAIL.n15 VTAIL.n14 585
R571 VTAIL.n4 VTAIL.n3 585
R572 VTAIL.n21 VTAIL.n20 585
R573 VTAIL.n23 VTAIL.n22 585
R574 VTAIL.n79 VTAIL.n78 585
R575 VTAIL.n77 VTAIL.n76 585
R576 VTAIL.n60 VTAIL.n59 585
R577 VTAIL.n71 VTAIL.n70 585
R578 VTAIL.n69 VTAIL.n68 585
R579 VTAIL.n64 VTAIL.n63 585
R580 VTAIL.n51 VTAIL.n50 585
R581 VTAIL.n49 VTAIL.n48 585
R582 VTAIL.n32 VTAIL.n31 585
R583 VTAIL.n43 VTAIL.n42 585
R584 VTAIL.n41 VTAIL.n40 585
R585 VTAIL.n36 VTAIL.n35 585
R586 VTAIL.n93 VTAIL.t2 327.856
R587 VTAIL.n9 VTAIL.t1 327.856
R588 VTAIL.n65 VTAIL.t0 327.856
R589 VTAIL.n37 VTAIL.t3 327.856
R590 VTAIL.n97 VTAIL.n91 171.744
R591 VTAIL.n98 VTAIL.n97 171.744
R592 VTAIL.n98 VTAIL.n87 171.744
R593 VTAIL.n105 VTAIL.n87 171.744
R594 VTAIL.n106 VTAIL.n105 171.744
R595 VTAIL.n13 VTAIL.n7 171.744
R596 VTAIL.n14 VTAIL.n13 171.744
R597 VTAIL.n14 VTAIL.n3 171.744
R598 VTAIL.n21 VTAIL.n3 171.744
R599 VTAIL.n22 VTAIL.n21 171.744
R600 VTAIL.n78 VTAIL.n77 171.744
R601 VTAIL.n77 VTAIL.n59 171.744
R602 VTAIL.n70 VTAIL.n59 171.744
R603 VTAIL.n70 VTAIL.n69 171.744
R604 VTAIL.n69 VTAIL.n63 171.744
R605 VTAIL.n50 VTAIL.n49 171.744
R606 VTAIL.n49 VTAIL.n31 171.744
R607 VTAIL.n42 VTAIL.n31 171.744
R608 VTAIL.n42 VTAIL.n41 171.744
R609 VTAIL.n41 VTAIL.n35 171.744
R610 VTAIL.t2 VTAIL.n91 85.8723
R611 VTAIL.t1 VTAIL.n7 85.8723
R612 VTAIL.t0 VTAIL.n63 85.8723
R613 VTAIL.t3 VTAIL.n35 85.8723
R614 VTAIL.n111 VTAIL.n110 32.1853
R615 VTAIL.n27 VTAIL.n26 32.1853
R616 VTAIL.n83 VTAIL.n82 32.1853
R617 VTAIL.n55 VTAIL.n54 32.1853
R618 VTAIL.n55 VTAIL.n27 19.6083
R619 VTAIL.n111 VTAIL.n83 18.2634
R620 VTAIL.n93 VTAIL.n92 16.381
R621 VTAIL.n9 VTAIL.n8 16.381
R622 VTAIL.n65 VTAIL.n64 16.381
R623 VTAIL.n37 VTAIL.n36 16.381
R624 VTAIL.n96 VTAIL.n95 12.8005
R625 VTAIL.n12 VTAIL.n11 12.8005
R626 VTAIL.n68 VTAIL.n67 12.8005
R627 VTAIL.n40 VTAIL.n39 12.8005
R628 VTAIL.n99 VTAIL.n90 12.0247
R629 VTAIL.n15 VTAIL.n6 12.0247
R630 VTAIL.n71 VTAIL.n62 12.0247
R631 VTAIL.n43 VTAIL.n34 12.0247
R632 VTAIL.n100 VTAIL.n88 11.249
R633 VTAIL.n16 VTAIL.n4 11.249
R634 VTAIL.n72 VTAIL.n60 11.249
R635 VTAIL.n44 VTAIL.n32 11.249
R636 VTAIL.n104 VTAIL.n103 10.4732
R637 VTAIL.n20 VTAIL.n19 10.4732
R638 VTAIL.n76 VTAIL.n75 10.4732
R639 VTAIL.n48 VTAIL.n47 10.4732
R640 VTAIL.n107 VTAIL.n86 9.69747
R641 VTAIL.n23 VTAIL.n2 9.69747
R642 VTAIL.n79 VTAIL.n58 9.69747
R643 VTAIL.n51 VTAIL.n30 9.69747
R644 VTAIL.n110 VTAIL.n109 9.45567
R645 VTAIL.n26 VTAIL.n25 9.45567
R646 VTAIL.n82 VTAIL.n81 9.45567
R647 VTAIL.n54 VTAIL.n53 9.45567
R648 VTAIL.n109 VTAIL.n108 9.3005
R649 VTAIL.n86 VTAIL.n85 9.3005
R650 VTAIL.n103 VTAIL.n102 9.3005
R651 VTAIL.n101 VTAIL.n100 9.3005
R652 VTAIL.n90 VTAIL.n89 9.3005
R653 VTAIL.n95 VTAIL.n94 9.3005
R654 VTAIL.n25 VTAIL.n24 9.3005
R655 VTAIL.n2 VTAIL.n1 9.3005
R656 VTAIL.n19 VTAIL.n18 9.3005
R657 VTAIL.n17 VTAIL.n16 9.3005
R658 VTAIL.n6 VTAIL.n5 9.3005
R659 VTAIL.n11 VTAIL.n10 9.3005
R660 VTAIL.n81 VTAIL.n80 9.3005
R661 VTAIL.n58 VTAIL.n57 9.3005
R662 VTAIL.n75 VTAIL.n74 9.3005
R663 VTAIL.n73 VTAIL.n72 9.3005
R664 VTAIL.n62 VTAIL.n61 9.3005
R665 VTAIL.n67 VTAIL.n66 9.3005
R666 VTAIL.n53 VTAIL.n52 9.3005
R667 VTAIL.n30 VTAIL.n29 9.3005
R668 VTAIL.n47 VTAIL.n46 9.3005
R669 VTAIL.n45 VTAIL.n44 9.3005
R670 VTAIL.n34 VTAIL.n33 9.3005
R671 VTAIL.n39 VTAIL.n38 9.3005
R672 VTAIL.n108 VTAIL.n84 8.92171
R673 VTAIL.n24 VTAIL.n0 8.92171
R674 VTAIL.n80 VTAIL.n56 8.92171
R675 VTAIL.n52 VTAIL.n28 8.92171
R676 VTAIL.n110 VTAIL.n84 5.04292
R677 VTAIL.n26 VTAIL.n0 5.04292
R678 VTAIL.n82 VTAIL.n56 5.04292
R679 VTAIL.n54 VTAIL.n28 5.04292
R680 VTAIL.n108 VTAIL.n107 4.26717
R681 VTAIL.n24 VTAIL.n23 4.26717
R682 VTAIL.n80 VTAIL.n79 4.26717
R683 VTAIL.n52 VTAIL.n51 4.26717
R684 VTAIL.n66 VTAIL.n65 3.71853
R685 VTAIL.n38 VTAIL.n37 3.71853
R686 VTAIL.n94 VTAIL.n93 3.71853
R687 VTAIL.n10 VTAIL.n9 3.71853
R688 VTAIL.n104 VTAIL.n86 3.49141
R689 VTAIL.n20 VTAIL.n2 3.49141
R690 VTAIL.n76 VTAIL.n58 3.49141
R691 VTAIL.n48 VTAIL.n30 3.49141
R692 VTAIL.n103 VTAIL.n88 2.71565
R693 VTAIL.n19 VTAIL.n4 2.71565
R694 VTAIL.n75 VTAIL.n60 2.71565
R695 VTAIL.n47 VTAIL.n32 2.71565
R696 VTAIL.n100 VTAIL.n99 1.93989
R697 VTAIL.n16 VTAIL.n15 1.93989
R698 VTAIL.n72 VTAIL.n71 1.93989
R699 VTAIL.n44 VTAIL.n43 1.93989
R700 VTAIL.n96 VTAIL.n90 1.16414
R701 VTAIL.n12 VTAIL.n6 1.16414
R702 VTAIL.n68 VTAIL.n62 1.16414
R703 VTAIL.n40 VTAIL.n34 1.16414
R704 VTAIL.n83 VTAIL.n55 1.14274
R705 VTAIL VTAIL.n27 0.864724
R706 VTAIL.n95 VTAIL.n92 0.388379
R707 VTAIL.n11 VTAIL.n8 0.388379
R708 VTAIL.n67 VTAIL.n64 0.388379
R709 VTAIL.n39 VTAIL.n36 0.388379
R710 VTAIL VTAIL.n111 0.278517
R711 VTAIL.n94 VTAIL.n89 0.155672
R712 VTAIL.n101 VTAIL.n89 0.155672
R713 VTAIL.n102 VTAIL.n101 0.155672
R714 VTAIL.n102 VTAIL.n85 0.155672
R715 VTAIL.n109 VTAIL.n85 0.155672
R716 VTAIL.n10 VTAIL.n5 0.155672
R717 VTAIL.n17 VTAIL.n5 0.155672
R718 VTAIL.n18 VTAIL.n17 0.155672
R719 VTAIL.n18 VTAIL.n1 0.155672
R720 VTAIL.n25 VTAIL.n1 0.155672
R721 VTAIL.n81 VTAIL.n57 0.155672
R722 VTAIL.n74 VTAIL.n57 0.155672
R723 VTAIL.n74 VTAIL.n73 0.155672
R724 VTAIL.n73 VTAIL.n61 0.155672
R725 VTAIL.n66 VTAIL.n61 0.155672
R726 VTAIL.n53 VTAIL.n29 0.155672
R727 VTAIL.n46 VTAIL.n29 0.155672
R728 VTAIL.n46 VTAIL.n45 0.155672
R729 VTAIL.n45 VTAIL.n33 0.155672
R730 VTAIL.n38 VTAIL.n33 0.155672
R731 VDD2.n49 VDD2.n27 756.745
R732 VDD2.n22 VDD2.n0 756.745
R733 VDD2.n50 VDD2.n49 585
R734 VDD2.n48 VDD2.n47 585
R735 VDD2.n31 VDD2.n30 585
R736 VDD2.n42 VDD2.n41 585
R737 VDD2.n40 VDD2.n39 585
R738 VDD2.n35 VDD2.n34 585
R739 VDD2.n8 VDD2.n7 585
R740 VDD2.n13 VDD2.n12 585
R741 VDD2.n15 VDD2.n14 585
R742 VDD2.n4 VDD2.n3 585
R743 VDD2.n21 VDD2.n20 585
R744 VDD2.n23 VDD2.n22 585
R745 VDD2.n36 VDD2.t1 327.856
R746 VDD2.n9 VDD2.t0 327.856
R747 VDD2.n49 VDD2.n48 171.744
R748 VDD2.n48 VDD2.n30 171.744
R749 VDD2.n41 VDD2.n30 171.744
R750 VDD2.n41 VDD2.n40 171.744
R751 VDD2.n40 VDD2.n34 171.744
R752 VDD2.n13 VDD2.n7 171.744
R753 VDD2.n14 VDD2.n13 171.744
R754 VDD2.n14 VDD2.n3 171.744
R755 VDD2.n21 VDD2.n3 171.744
R756 VDD2.n22 VDD2.n21 171.744
R757 VDD2.t1 VDD2.n34 85.8723
R758 VDD2.t0 VDD2.n7 85.8723
R759 VDD2.n54 VDD2.n26 79.765
R760 VDD2.n54 VDD2.n53 48.8641
R761 VDD2.n36 VDD2.n35 16.381
R762 VDD2.n9 VDD2.n8 16.381
R763 VDD2.n39 VDD2.n38 12.8005
R764 VDD2.n12 VDD2.n11 12.8005
R765 VDD2.n42 VDD2.n33 12.0247
R766 VDD2.n15 VDD2.n6 12.0247
R767 VDD2.n43 VDD2.n31 11.249
R768 VDD2.n16 VDD2.n4 11.249
R769 VDD2.n47 VDD2.n46 10.4732
R770 VDD2.n20 VDD2.n19 10.4732
R771 VDD2.n50 VDD2.n29 9.69747
R772 VDD2.n23 VDD2.n2 9.69747
R773 VDD2.n53 VDD2.n52 9.45567
R774 VDD2.n26 VDD2.n25 9.45567
R775 VDD2.n52 VDD2.n51 9.3005
R776 VDD2.n29 VDD2.n28 9.3005
R777 VDD2.n46 VDD2.n45 9.3005
R778 VDD2.n44 VDD2.n43 9.3005
R779 VDD2.n33 VDD2.n32 9.3005
R780 VDD2.n38 VDD2.n37 9.3005
R781 VDD2.n25 VDD2.n24 9.3005
R782 VDD2.n2 VDD2.n1 9.3005
R783 VDD2.n19 VDD2.n18 9.3005
R784 VDD2.n17 VDD2.n16 9.3005
R785 VDD2.n6 VDD2.n5 9.3005
R786 VDD2.n11 VDD2.n10 9.3005
R787 VDD2.n51 VDD2.n27 8.92171
R788 VDD2.n24 VDD2.n0 8.92171
R789 VDD2.n53 VDD2.n27 5.04292
R790 VDD2.n26 VDD2.n0 5.04292
R791 VDD2.n51 VDD2.n50 4.26717
R792 VDD2.n24 VDD2.n23 4.26717
R793 VDD2.n37 VDD2.n36 3.71853
R794 VDD2.n10 VDD2.n9 3.71853
R795 VDD2.n47 VDD2.n29 3.49141
R796 VDD2.n20 VDD2.n2 3.49141
R797 VDD2.n46 VDD2.n31 2.71565
R798 VDD2.n19 VDD2.n4 2.71565
R799 VDD2.n43 VDD2.n42 1.93989
R800 VDD2.n16 VDD2.n15 1.93989
R801 VDD2.n39 VDD2.n33 1.16414
R802 VDD2.n12 VDD2.n6 1.16414
R803 VDD2 VDD2.n54 0.394897
R804 VDD2.n38 VDD2.n35 0.388379
R805 VDD2.n11 VDD2.n8 0.388379
R806 VDD2.n52 VDD2.n28 0.155672
R807 VDD2.n45 VDD2.n28 0.155672
R808 VDD2.n45 VDD2.n44 0.155672
R809 VDD2.n44 VDD2.n32 0.155672
R810 VDD2.n37 VDD2.n32 0.155672
R811 VDD2.n10 VDD2.n5 0.155672
R812 VDD2.n17 VDD2.n5 0.155672
R813 VDD2.n18 VDD2.n17 0.155672
R814 VDD2.n18 VDD2.n1 0.155672
R815 VDD2.n25 VDD2.n1 0.155672
R816 VP.n0 VP.t1 251.928
R817 VP.n0 VP.t0 215.994
R818 VP VP.n0 0.146778
R819 VDD1.n22 VDD1.n0 756.745
R820 VDD1.n49 VDD1.n27 756.745
R821 VDD1.n23 VDD1.n22 585
R822 VDD1.n21 VDD1.n20 585
R823 VDD1.n4 VDD1.n3 585
R824 VDD1.n15 VDD1.n14 585
R825 VDD1.n13 VDD1.n12 585
R826 VDD1.n8 VDD1.n7 585
R827 VDD1.n35 VDD1.n34 585
R828 VDD1.n40 VDD1.n39 585
R829 VDD1.n42 VDD1.n41 585
R830 VDD1.n31 VDD1.n30 585
R831 VDD1.n48 VDD1.n47 585
R832 VDD1.n50 VDD1.n49 585
R833 VDD1.n9 VDD1.t0 327.856
R834 VDD1.n36 VDD1.t1 327.856
R835 VDD1.n22 VDD1.n21 171.744
R836 VDD1.n21 VDD1.n3 171.744
R837 VDD1.n14 VDD1.n3 171.744
R838 VDD1.n14 VDD1.n13 171.744
R839 VDD1.n13 VDD1.n7 171.744
R840 VDD1.n40 VDD1.n34 171.744
R841 VDD1.n41 VDD1.n40 171.744
R842 VDD1.n41 VDD1.n30 171.744
R843 VDD1.n48 VDD1.n30 171.744
R844 VDD1.n49 VDD1.n48 171.744
R845 VDD1.t0 VDD1.n7 85.8723
R846 VDD1.t1 VDD1.n34 85.8723
R847 VDD1 VDD1.n53 80.626
R848 VDD1 VDD1.n26 49.2585
R849 VDD1.n9 VDD1.n8 16.381
R850 VDD1.n36 VDD1.n35 16.381
R851 VDD1.n12 VDD1.n11 12.8005
R852 VDD1.n39 VDD1.n38 12.8005
R853 VDD1.n15 VDD1.n6 12.0247
R854 VDD1.n42 VDD1.n33 12.0247
R855 VDD1.n16 VDD1.n4 11.249
R856 VDD1.n43 VDD1.n31 11.249
R857 VDD1.n20 VDD1.n19 10.4732
R858 VDD1.n47 VDD1.n46 10.4732
R859 VDD1.n23 VDD1.n2 9.69747
R860 VDD1.n50 VDD1.n29 9.69747
R861 VDD1.n26 VDD1.n25 9.45567
R862 VDD1.n53 VDD1.n52 9.45567
R863 VDD1.n25 VDD1.n24 9.3005
R864 VDD1.n2 VDD1.n1 9.3005
R865 VDD1.n19 VDD1.n18 9.3005
R866 VDD1.n17 VDD1.n16 9.3005
R867 VDD1.n6 VDD1.n5 9.3005
R868 VDD1.n11 VDD1.n10 9.3005
R869 VDD1.n52 VDD1.n51 9.3005
R870 VDD1.n29 VDD1.n28 9.3005
R871 VDD1.n46 VDD1.n45 9.3005
R872 VDD1.n44 VDD1.n43 9.3005
R873 VDD1.n33 VDD1.n32 9.3005
R874 VDD1.n38 VDD1.n37 9.3005
R875 VDD1.n24 VDD1.n0 8.92171
R876 VDD1.n51 VDD1.n27 8.92171
R877 VDD1.n26 VDD1.n0 5.04292
R878 VDD1.n53 VDD1.n27 5.04292
R879 VDD1.n24 VDD1.n23 4.26717
R880 VDD1.n51 VDD1.n50 4.26717
R881 VDD1.n10 VDD1.n9 3.71853
R882 VDD1.n37 VDD1.n36 3.71853
R883 VDD1.n20 VDD1.n2 3.49141
R884 VDD1.n47 VDD1.n29 3.49141
R885 VDD1.n19 VDD1.n4 2.71565
R886 VDD1.n46 VDD1.n31 2.71565
R887 VDD1.n16 VDD1.n15 1.93989
R888 VDD1.n43 VDD1.n42 1.93989
R889 VDD1.n12 VDD1.n6 1.16414
R890 VDD1.n39 VDD1.n33 1.16414
R891 VDD1.n11 VDD1.n8 0.388379
R892 VDD1.n38 VDD1.n35 0.388379
R893 VDD1.n25 VDD1.n1 0.155672
R894 VDD1.n18 VDD1.n1 0.155672
R895 VDD1.n18 VDD1.n17 0.155672
R896 VDD1.n17 VDD1.n5 0.155672
R897 VDD1.n10 VDD1.n5 0.155672
R898 VDD1.n37 VDD1.n32 0.155672
R899 VDD1.n44 VDD1.n32 0.155672
R900 VDD1.n45 VDD1.n44 0.155672
R901 VDD1.n45 VDD1.n28 0.155672
R902 VDD1.n52 VDD1.n28 0.155672
C0 VP w_n1594_n2024# 2.15394f
C1 VN VDD1 0.147828f
C2 VTAIL B 1.68784f
C3 VN VDD2 1.18199f
C4 VTAIL VDD1 3.05911f
C5 VTAIL VDD2 3.10104f
C6 VN VP 3.5677f
C7 VDD1 B 1.00003f
C8 VDD2 B 1.01851f
C9 VN w_n1594_n2024# 1.95393f
C10 VP VTAIL 1.10931f
C11 VDD2 VDD1 0.515086f
C12 VP B 1.06475f
C13 VTAIL w_n1594_n2024# 1.77468f
C14 w_n1594_n2024# B 5.44825f
C15 VP VDD1 1.30763f
C16 VP VDD2 0.279122f
C17 w_n1594_n2024# VDD1 1.14348f
C18 w_n1594_n2024# VDD2 1.15313f
C19 VN VTAIL 1.09504f
C20 VN B 0.741301f
C21 VDD2 VSUBS 0.537048f
C22 VDD1 VSUBS 1.97485f
C23 VTAIL VSUBS 0.428194f
C24 VN VSUBS 3.66701f
C25 VP VSUBS 0.948092f
C26 B VSUBS 2.211889f
C27 w_n1594_n2024# VSUBS 40.3792f
C28 VDD1.n0 VSUBS 0.015981f
C29 VDD1.n1 VSUBS 0.014829f
C30 VDD1.n2 VSUBS 0.007969f
C31 VDD1.n3 VSUBS 0.018835f
C32 VDD1.n4 VSUBS 0.008437f
C33 VDD1.n5 VSUBS 0.014829f
C34 VDD1.n6 VSUBS 0.007969f
C35 VDD1.n7 VSUBS 0.014126f
C36 VDD1.n8 VSUBS 0.011964f
C37 VDD1.t0 VSUBS 0.040614f
C38 VDD1.n9 VSUBS 0.062602f
C39 VDD1.n10 VSUBS 0.291306f
C40 VDD1.n11 VSUBS 0.007969f
C41 VDD1.n12 VSUBS 0.008437f
C42 VDD1.n13 VSUBS 0.018835f
C43 VDD1.n14 VSUBS 0.018835f
C44 VDD1.n15 VSUBS 0.008437f
C45 VDD1.n16 VSUBS 0.007969f
C46 VDD1.n17 VSUBS 0.014829f
C47 VDD1.n18 VSUBS 0.014829f
C48 VDD1.n19 VSUBS 0.007969f
C49 VDD1.n20 VSUBS 0.008437f
C50 VDD1.n21 VSUBS 0.018835f
C51 VDD1.n22 VSUBS 0.04453f
C52 VDD1.n23 VSUBS 0.008437f
C53 VDD1.n24 VSUBS 0.007969f
C54 VDD1.n25 VSUBS 0.034277f
C55 VDD1.n26 VSUBS 0.032965f
C56 VDD1.n27 VSUBS 0.015981f
C57 VDD1.n28 VSUBS 0.014829f
C58 VDD1.n29 VSUBS 0.007969f
C59 VDD1.n30 VSUBS 0.018835f
C60 VDD1.n31 VSUBS 0.008437f
C61 VDD1.n32 VSUBS 0.014829f
C62 VDD1.n33 VSUBS 0.007969f
C63 VDD1.n34 VSUBS 0.014126f
C64 VDD1.n35 VSUBS 0.011964f
C65 VDD1.t1 VSUBS 0.040614f
C66 VDD1.n36 VSUBS 0.062602f
C67 VDD1.n37 VSUBS 0.291306f
C68 VDD1.n38 VSUBS 0.007969f
C69 VDD1.n39 VSUBS 0.008437f
C70 VDD1.n40 VSUBS 0.018835f
C71 VDD1.n41 VSUBS 0.018835f
C72 VDD1.n42 VSUBS 0.008437f
C73 VDD1.n43 VSUBS 0.007969f
C74 VDD1.n44 VSUBS 0.014829f
C75 VDD1.n45 VSUBS 0.014829f
C76 VDD1.n46 VSUBS 0.007969f
C77 VDD1.n47 VSUBS 0.008437f
C78 VDD1.n48 VSUBS 0.018835f
C79 VDD1.n49 VSUBS 0.04453f
C80 VDD1.n50 VSUBS 0.008437f
C81 VDD1.n51 VSUBS 0.007969f
C82 VDD1.n52 VSUBS 0.034277f
C83 VDD1.n53 VSUBS 0.277452f
C84 VP.t1 VSUBS 1.32458f
C85 VP.t0 VSUBS 1.06651f
C86 VP.n0 VSUBS 3.36704f
C87 VDD2.n0 VSUBS 0.016268f
C88 VDD2.n1 VSUBS 0.015096f
C89 VDD2.n2 VSUBS 0.008112f
C90 VDD2.n3 VSUBS 0.019174f
C91 VDD2.n4 VSUBS 0.008589f
C92 VDD2.n5 VSUBS 0.015096f
C93 VDD2.n6 VSUBS 0.008112f
C94 VDD2.n7 VSUBS 0.01438f
C95 VDD2.n8 VSUBS 0.012179f
C96 VDD2.t0 VSUBS 0.041344f
C97 VDD2.n9 VSUBS 0.063728f
C98 VDD2.n10 VSUBS 0.296545f
C99 VDD2.n11 VSUBS 0.008112f
C100 VDD2.n12 VSUBS 0.008589f
C101 VDD2.n13 VSUBS 0.019174f
C102 VDD2.n14 VSUBS 0.019174f
C103 VDD2.n15 VSUBS 0.008589f
C104 VDD2.n16 VSUBS 0.008112f
C105 VDD2.n17 VSUBS 0.015096f
C106 VDD2.n18 VSUBS 0.015096f
C107 VDD2.n19 VSUBS 0.008112f
C108 VDD2.n20 VSUBS 0.008589f
C109 VDD2.n21 VSUBS 0.019174f
C110 VDD2.n22 VSUBS 0.045331f
C111 VDD2.n23 VSUBS 0.008589f
C112 VDD2.n24 VSUBS 0.008112f
C113 VDD2.n25 VSUBS 0.034894f
C114 VDD2.n26 VSUBS 0.262756f
C115 VDD2.n27 VSUBS 0.016268f
C116 VDD2.n28 VSUBS 0.015096f
C117 VDD2.n29 VSUBS 0.008112f
C118 VDD2.n30 VSUBS 0.019174f
C119 VDD2.n31 VSUBS 0.008589f
C120 VDD2.n32 VSUBS 0.015096f
C121 VDD2.n33 VSUBS 0.008112f
C122 VDD2.n34 VSUBS 0.01438f
C123 VDD2.n35 VSUBS 0.012179f
C124 VDD2.t1 VSUBS 0.041344f
C125 VDD2.n36 VSUBS 0.063728f
C126 VDD2.n37 VSUBS 0.296545f
C127 VDD2.n38 VSUBS 0.008112f
C128 VDD2.n39 VSUBS 0.008589f
C129 VDD2.n40 VSUBS 0.019174f
C130 VDD2.n41 VSUBS 0.019174f
C131 VDD2.n42 VSUBS 0.008589f
C132 VDD2.n43 VSUBS 0.008112f
C133 VDD2.n44 VSUBS 0.015096f
C134 VDD2.n45 VSUBS 0.015096f
C135 VDD2.n46 VSUBS 0.008112f
C136 VDD2.n47 VSUBS 0.008589f
C137 VDD2.n48 VSUBS 0.019174f
C138 VDD2.n49 VSUBS 0.045331f
C139 VDD2.n50 VSUBS 0.008589f
C140 VDD2.n51 VSUBS 0.008112f
C141 VDD2.n52 VSUBS 0.034894f
C142 VDD2.n53 VSUBS 0.033172f
C143 VDD2.n54 VSUBS 1.24503f
C144 VTAIL.n0 VSUBS 0.018417f
C145 VTAIL.n1 VSUBS 0.01709f
C146 VTAIL.n2 VSUBS 0.009183f
C147 VTAIL.n3 VSUBS 0.021706f
C148 VTAIL.n4 VSUBS 0.009724f
C149 VTAIL.n5 VSUBS 0.01709f
C150 VTAIL.n6 VSUBS 0.009183f
C151 VTAIL.n7 VSUBS 0.01628f
C152 VTAIL.n8 VSUBS 0.013788f
C153 VTAIL.t1 VSUBS 0.046805f
C154 VTAIL.n9 VSUBS 0.072145f
C155 VTAIL.n10 VSUBS 0.335712f
C156 VTAIL.n11 VSUBS 0.009183f
C157 VTAIL.n12 VSUBS 0.009724f
C158 VTAIL.n13 VSUBS 0.021706f
C159 VTAIL.n14 VSUBS 0.021706f
C160 VTAIL.n15 VSUBS 0.009724f
C161 VTAIL.n16 VSUBS 0.009183f
C162 VTAIL.n17 VSUBS 0.01709f
C163 VTAIL.n18 VSUBS 0.01709f
C164 VTAIL.n19 VSUBS 0.009183f
C165 VTAIL.n20 VSUBS 0.009724f
C166 VTAIL.n21 VSUBS 0.021706f
C167 VTAIL.n22 VSUBS 0.051318f
C168 VTAIL.n23 VSUBS 0.009724f
C169 VTAIL.n24 VSUBS 0.009183f
C170 VTAIL.n25 VSUBS 0.039503f
C171 VTAIL.n26 VSUBS 0.025753f
C172 VTAIL.n27 VSUBS 0.693097f
C173 VTAIL.n28 VSUBS 0.018417f
C174 VTAIL.n29 VSUBS 0.01709f
C175 VTAIL.n30 VSUBS 0.009183f
C176 VTAIL.n31 VSUBS 0.021706f
C177 VTAIL.n32 VSUBS 0.009724f
C178 VTAIL.n33 VSUBS 0.01709f
C179 VTAIL.n34 VSUBS 0.009183f
C180 VTAIL.n35 VSUBS 0.01628f
C181 VTAIL.n36 VSUBS 0.013788f
C182 VTAIL.t3 VSUBS 0.046805f
C183 VTAIL.n37 VSUBS 0.072145f
C184 VTAIL.n38 VSUBS 0.335712f
C185 VTAIL.n39 VSUBS 0.009183f
C186 VTAIL.n40 VSUBS 0.009724f
C187 VTAIL.n41 VSUBS 0.021706f
C188 VTAIL.n42 VSUBS 0.021706f
C189 VTAIL.n43 VSUBS 0.009724f
C190 VTAIL.n44 VSUBS 0.009183f
C191 VTAIL.n45 VSUBS 0.01709f
C192 VTAIL.n46 VSUBS 0.01709f
C193 VTAIL.n47 VSUBS 0.009183f
C194 VTAIL.n48 VSUBS 0.009724f
C195 VTAIL.n49 VSUBS 0.021706f
C196 VTAIL.n50 VSUBS 0.051318f
C197 VTAIL.n51 VSUBS 0.009724f
C198 VTAIL.n52 VSUBS 0.009183f
C199 VTAIL.n53 VSUBS 0.039503f
C200 VTAIL.n54 VSUBS 0.025753f
C201 VTAIL.n55 VSUBS 0.708407f
C202 VTAIL.n56 VSUBS 0.018417f
C203 VTAIL.n57 VSUBS 0.01709f
C204 VTAIL.n58 VSUBS 0.009183f
C205 VTAIL.n59 VSUBS 0.021706f
C206 VTAIL.n60 VSUBS 0.009724f
C207 VTAIL.n61 VSUBS 0.01709f
C208 VTAIL.n62 VSUBS 0.009183f
C209 VTAIL.n63 VSUBS 0.01628f
C210 VTAIL.n64 VSUBS 0.013788f
C211 VTAIL.t0 VSUBS 0.046805f
C212 VTAIL.n65 VSUBS 0.072145f
C213 VTAIL.n66 VSUBS 0.335712f
C214 VTAIL.n67 VSUBS 0.009183f
C215 VTAIL.n68 VSUBS 0.009724f
C216 VTAIL.n69 VSUBS 0.021706f
C217 VTAIL.n70 VSUBS 0.021706f
C218 VTAIL.n71 VSUBS 0.009724f
C219 VTAIL.n72 VSUBS 0.009183f
C220 VTAIL.n73 VSUBS 0.01709f
C221 VTAIL.n74 VSUBS 0.01709f
C222 VTAIL.n75 VSUBS 0.009183f
C223 VTAIL.n76 VSUBS 0.009724f
C224 VTAIL.n77 VSUBS 0.021706f
C225 VTAIL.n78 VSUBS 0.051318f
C226 VTAIL.n79 VSUBS 0.009724f
C227 VTAIL.n80 VSUBS 0.009183f
C228 VTAIL.n81 VSUBS 0.039503f
C229 VTAIL.n82 VSUBS 0.025753f
C230 VTAIL.n83 VSUBS 0.63435f
C231 VTAIL.n84 VSUBS 0.018417f
C232 VTAIL.n85 VSUBS 0.01709f
C233 VTAIL.n86 VSUBS 0.009183f
C234 VTAIL.n87 VSUBS 0.021706f
C235 VTAIL.n88 VSUBS 0.009724f
C236 VTAIL.n89 VSUBS 0.01709f
C237 VTAIL.n90 VSUBS 0.009183f
C238 VTAIL.n91 VSUBS 0.01628f
C239 VTAIL.n92 VSUBS 0.013788f
C240 VTAIL.t2 VSUBS 0.046805f
C241 VTAIL.n93 VSUBS 0.072145f
C242 VTAIL.n94 VSUBS 0.335712f
C243 VTAIL.n95 VSUBS 0.009183f
C244 VTAIL.n96 VSUBS 0.009724f
C245 VTAIL.n97 VSUBS 0.021706f
C246 VTAIL.n98 VSUBS 0.021706f
C247 VTAIL.n99 VSUBS 0.009724f
C248 VTAIL.n100 VSUBS 0.009183f
C249 VTAIL.n101 VSUBS 0.01709f
C250 VTAIL.n102 VSUBS 0.01709f
C251 VTAIL.n103 VSUBS 0.009183f
C252 VTAIL.n104 VSUBS 0.009724f
C253 VTAIL.n105 VSUBS 0.021706f
C254 VTAIL.n106 VSUBS 0.051318f
C255 VTAIL.n107 VSUBS 0.009724f
C256 VTAIL.n108 VSUBS 0.009183f
C257 VTAIL.n109 VSUBS 0.039503f
C258 VTAIL.n110 VSUBS 0.025753f
C259 VTAIL.n111 VSUBS 0.58676f
C260 VN.t1 VSUBS 0.654487f
C261 VN.t0 VSUBS 0.816213f
C262 B.n0 VSUBS 0.005798f
C263 B.n1 VSUBS 0.005798f
C264 B.n2 VSUBS 0.008575f
C265 B.n3 VSUBS 0.006571f
C266 B.n4 VSUBS 0.006571f
C267 B.n5 VSUBS 0.006571f
C268 B.n6 VSUBS 0.006571f
C269 B.n7 VSUBS 0.006571f
C270 B.n8 VSUBS 0.006571f
C271 B.n9 VSUBS 0.006571f
C272 B.n10 VSUBS 0.014929f
C273 B.n11 VSUBS 0.006571f
C274 B.n12 VSUBS 0.006571f
C275 B.n13 VSUBS 0.006571f
C276 B.n14 VSUBS 0.006571f
C277 B.n15 VSUBS 0.006571f
C278 B.n16 VSUBS 0.006571f
C279 B.n17 VSUBS 0.006571f
C280 B.n18 VSUBS 0.006571f
C281 B.n19 VSUBS 0.006571f
C282 B.n20 VSUBS 0.006571f
C283 B.n21 VSUBS 0.006571f
C284 B.t10 VSUBS 0.072519f
C285 B.t11 VSUBS 0.085134f
C286 B.t9 VSUBS 0.277942f
C287 B.n22 VSUBS 0.152069f
C288 B.n23 VSUBS 0.128584f
C289 B.n24 VSUBS 0.006571f
C290 B.n25 VSUBS 0.006571f
C291 B.n26 VSUBS 0.006571f
C292 B.n27 VSUBS 0.006571f
C293 B.t7 VSUBS 0.072521f
C294 B.t8 VSUBS 0.085135f
C295 B.t6 VSUBS 0.277942f
C296 B.n28 VSUBS 0.152068f
C297 B.n29 VSUBS 0.128583f
C298 B.n30 VSUBS 0.015225f
C299 B.n31 VSUBS 0.006571f
C300 B.n32 VSUBS 0.006571f
C301 B.n33 VSUBS 0.006571f
C302 B.n34 VSUBS 0.006571f
C303 B.n35 VSUBS 0.006571f
C304 B.n36 VSUBS 0.006571f
C305 B.n37 VSUBS 0.006571f
C306 B.n38 VSUBS 0.006571f
C307 B.n39 VSUBS 0.006571f
C308 B.n40 VSUBS 0.006571f
C309 B.n41 VSUBS 0.015222f
C310 B.n42 VSUBS 0.006571f
C311 B.n43 VSUBS 0.006571f
C312 B.n44 VSUBS 0.006571f
C313 B.n45 VSUBS 0.006571f
C314 B.n46 VSUBS 0.006571f
C315 B.n47 VSUBS 0.006571f
C316 B.n48 VSUBS 0.006571f
C317 B.n49 VSUBS 0.006571f
C318 B.n50 VSUBS 0.006571f
C319 B.n51 VSUBS 0.006571f
C320 B.n52 VSUBS 0.006571f
C321 B.n53 VSUBS 0.006571f
C322 B.n54 VSUBS 0.006571f
C323 B.n55 VSUBS 0.006571f
C324 B.n56 VSUBS 0.006571f
C325 B.n57 VSUBS 0.006571f
C326 B.n58 VSUBS 0.006571f
C327 B.n59 VSUBS 0.014929f
C328 B.n60 VSUBS 0.006571f
C329 B.n61 VSUBS 0.006571f
C330 B.n62 VSUBS 0.006571f
C331 B.n63 VSUBS 0.006571f
C332 B.n64 VSUBS 0.006571f
C333 B.n65 VSUBS 0.006571f
C334 B.n66 VSUBS 0.006571f
C335 B.n67 VSUBS 0.006571f
C336 B.n68 VSUBS 0.006571f
C337 B.n69 VSUBS 0.006571f
C338 B.n70 VSUBS 0.004542f
C339 B.n71 VSUBS 0.006571f
C340 B.n72 VSUBS 0.006571f
C341 B.n73 VSUBS 0.006571f
C342 B.n74 VSUBS 0.006571f
C343 B.n75 VSUBS 0.006571f
C344 B.t5 VSUBS 0.072519f
C345 B.t4 VSUBS 0.085134f
C346 B.t3 VSUBS 0.277942f
C347 B.n76 VSUBS 0.152069f
C348 B.n77 VSUBS 0.128584f
C349 B.n78 VSUBS 0.006571f
C350 B.n79 VSUBS 0.006571f
C351 B.n80 VSUBS 0.006571f
C352 B.n81 VSUBS 0.006571f
C353 B.n82 VSUBS 0.006571f
C354 B.n83 VSUBS 0.006571f
C355 B.n84 VSUBS 0.006571f
C356 B.n85 VSUBS 0.006571f
C357 B.n86 VSUBS 0.006571f
C358 B.n87 VSUBS 0.006571f
C359 B.n88 VSUBS 0.014929f
C360 B.n89 VSUBS 0.006571f
C361 B.n90 VSUBS 0.006571f
C362 B.n91 VSUBS 0.006571f
C363 B.n92 VSUBS 0.006571f
C364 B.n93 VSUBS 0.006571f
C365 B.n94 VSUBS 0.006571f
C366 B.n95 VSUBS 0.006571f
C367 B.n96 VSUBS 0.006571f
C368 B.n97 VSUBS 0.006571f
C369 B.n98 VSUBS 0.006571f
C370 B.n99 VSUBS 0.006571f
C371 B.n100 VSUBS 0.006571f
C372 B.n101 VSUBS 0.006571f
C373 B.n102 VSUBS 0.006571f
C374 B.n103 VSUBS 0.006571f
C375 B.n104 VSUBS 0.006571f
C376 B.n105 VSUBS 0.006571f
C377 B.n106 VSUBS 0.006571f
C378 B.n107 VSUBS 0.006571f
C379 B.n108 VSUBS 0.006571f
C380 B.n109 VSUBS 0.006571f
C381 B.n110 VSUBS 0.006571f
C382 B.n111 VSUBS 0.006571f
C383 B.n112 VSUBS 0.006571f
C384 B.n113 VSUBS 0.006571f
C385 B.n114 VSUBS 0.006571f
C386 B.n115 VSUBS 0.006571f
C387 B.n116 VSUBS 0.006571f
C388 B.n117 VSUBS 0.006571f
C389 B.n118 VSUBS 0.006571f
C390 B.n119 VSUBS 0.014929f
C391 B.n120 VSUBS 0.015222f
C392 B.n121 VSUBS 0.015222f
C393 B.n122 VSUBS 0.006571f
C394 B.n123 VSUBS 0.006571f
C395 B.n124 VSUBS 0.006571f
C396 B.n125 VSUBS 0.006571f
C397 B.n126 VSUBS 0.006571f
C398 B.n127 VSUBS 0.006571f
C399 B.n128 VSUBS 0.006571f
C400 B.n129 VSUBS 0.006571f
C401 B.n130 VSUBS 0.006571f
C402 B.n131 VSUBS 0.006571f
C403 B.n132 VSUBS 0.006571f
C404 B.n133 VSUBS 0.006571f
C405 B.n134 VSUBS 0.006571f
C406 B.n135 VSUBS 0.006571f
C407 B.n136 VSUBS 0.006571f
C408 B.n137 VSUBS 0.006571f
C409 B.n138 VSUBS 0.006571f
C410 B.n139 VSUBS 0.006571f
C411 B.n140 VSUBS 0.006571f
C412 B.n141 VSUBS 0.006571f
C413 B.n142 VSUBS 0.006571f
C414 B.n143 VSUBS 0.006571f
C415 B.n144 VSUBS 0.006571f
C416 B.n145 VSUBS 0.006571f
C417 B.n146 VSUBS 0.006571f
C418 B.n147 VSUBS 0.006571f
C419 B.n148 VSUBS 0.006571f
C420 B.n149 VSUBS 0.006571f
C421 B.n150 VSUBS 0.006571f
C422 B.n151 VSUBS 0.006571f
C423 B.n152 VSUBS 0.004542f
C424 B.n153 VSUBS 0.015225f
C425 B.n154 VSUBS 0.005315f
C426 B.n155 VSUBS 0.006571f
C427 B.n156 VSUBS 0.006571f
C428 B.n157 VSUBS 0.006571f
C429 B.n158 VSUBS 0.006571f
C430 B.n159 VSUBS 0.006571f
C431 B.n160 VSUBS 0.006571f
C432 B.n161 VSUBS 0.006571f
C433 B.n162 VSUBS 0.006571f
C434 B.n163 VSUBS 0.006571f
C435 B.n164 VSUBS 0.006571f
C436 B.n165 VSUBS 0.006571f
C437 B.t2 VSUBS 0.072521f
C438 B.t1 VSUBS 0.085135f
C439 B.t0 VSUBS 0.277942f
C440 B.n166 VSUBS 0.152068f
C441 B.n167 VSUBS 0.128583f
C442 B.n168 VSUBS 0.015225f
C443 B.n169 VSUBS 0.005315f
C444 B.n170 VSUBS 0.006571f
C445 B.n171 VSUBS 0.006571f
C446 B.n172 VSUBS 0.006571f
C447 B.n173 VSUBS 0.006571f
C448 B.n174 VSUBS 0.006571f
C449 B.n175 VSUBS 0.006571f
C450 B.n176 VSUBS 0.006571f
C451 B.n177 VSUBS 0.006571f
C452 B.n178 VSUBS 0.006571f
C453 B.n179 VSUBS 0.006571f
C454 B.n180 VSUBS 0.006571f
C455 B.n181 VSUBS 0.006571f
C456 B.n182 VSUBS 0.006571f
C457 B.n183 VSUBS 0.006571f
C458 B.n184 VSUBS 0.006571f
C459 B.n185 VSUBS 0.006571f
C460 B.n186 VSUBS 0.006571f
C461 B.n187 VSUBS 0.006571f
C462 B.n188 VSUBS 0.006571f
C463 B.n189 VSUBS 0.006571f
C464 B.n190 VSUBS 0.006571f
C465 B.n191 VSUBS 0.006571f
C466 B.n192 VSUBS 0.006571f
C467 B.n193 VSUBS 0.006571f
C468 B.n194 VSUBS 0.006571f
C469 B.n195 VSUBS 0.006571f
C470 B.n196 VSUBS 0.006571f
C471 B.n197 VSUBS 0.006571f
C472 B.n198 VSUBS 0.006571f
C473 B.n199 VSUBS 0.006571f
C474 B.n200 VSUBS 0.006571f
C475 B.n201 VSUBS 0.006571f
C476 B.n202 VSUBS 0.015222f
C477 B.n203 VSUBS 0.014422f
C478 B.n204 VSUBS 0.015729f
C479 B.n205 VSUBS 0.006571f
C480 B.n206 VSUBS 0.006571f
C481 B.n207 VSUBS 0.006571f
C482 B.n208 VSUBS 0.006571f
C483 B.n209 VSUBS 0.006571f
C484 B.n210 VSUBS 0.006571f
C485 B.n211 VSUBS 0.006571f
C486 B.n212 VSUBS 0.006571f
C487 B.n213 VSUBS 0.006571f
C488 B.n214 VSUBS 0.006571f
C489 B.n215 VSUBS 0.006571f
C490 B.n216 VSUBS 0.006571f
C491 B.n217 VSUBS 0.006571f
C492 B.n218 VSUBS 0.006571f
C493 B.n219 VSUBS 0.006571f
C494 B.n220 VSUBS 0.006571f
C495 B.n221 VSUBS 0.006571f
C496 B.n222 VSUBS 0.006571f
C497 B.n223 VSUBS 0.006571f
C498 B.n224 VSUBS 0.006571f
C499 B.n225 VSUBS 0.006571f
C500 B.n226 VSUBS 0.006571f
C501 B.n227 VSUBS 0.006571f
C502 B.n228 VSUBS 0.006571f
C503 B.n229 VSUBS 0.006571f
C504 B.n230 VSUBS 0.006571f
C505 B.n231 VSUBS 0.006571f
C506 B.n232 VSUBS 0.006571f
C507 B.n233 VSUBS 0.006571f
C508 B.n234 VSUBS 0.006571f
C509 B.n235 VSUBS 0.006571f
C510 B.n236 VSUBS 0.006571f
C511 B.n237 VSUBS 0.006571f
C512 B.n238 VSUBS 0.006571f
C513 B.n239 VSUBS 0.006571f
C514 B.n240 VSUBS 0.006571f
C515 B.n241 VSUBS 0.006571f
C516 B.n242 VSUBS 0.006571f
C517 B.n243 VSUBS 0.006571f
C518 B.n244 VSUBS 0.006571f
C519 B.n245 VSUBS 0.006571f
C520 B.n246 VSUBS 0.006571f
C521 B.n247 VSUBS 0.006571f
C522 B.n248 VSUBS 0.006571f
C523 B.n249 VSUBS 0.006571f
C524 B.n250 VSUBS 0.006571f
C525 B.n251 VSUBS 0.006571f
C526 B.n252 VSUBS 0.006571f
C527 B.n253 VSUBS 0.006571f
C528 B.n254 VSUBS 0.006571f
C529 B.n255 VSUBS 0.006571f
C530 B.n256 VSUBS 0.014929f
C531 B.n257 VSUBS 0.014929f
C532 B.n258 VSUBS 0.015222f
C533 B.n259 VSUBS 0.006571f
C534 B.n260 VSUBS 0.006571f
C535 B.n261 VSUBS 0.006571f
C536 B.n262 VSUBS 0.006571f
C537 B.n263 VSUBS 0.006571f
C538 B.n264 VSUBS 0.006571f
C539 B.n265 VSUBS 0.006571f
C540 B.n266 VSUBS 0.006571f
C541 B.n267 VSUBS 0.006571f
C542 B.n268 VSUBS 0.006571f
C543 B.n269 VSUBS 0.006571f
C544 B.n270 VSUBS 0.006571f
C545 B.n271 VSUBS 0.006571f
C546 B.n272 VSUBS 0.006571f
C547 B.n273 VSUBS 0.006571f
C548 B.n274 VSUBS 0.006571f
C549 B.n275 VSUBS 0.006571f
C550 B.n276 VSUBS 0.006571f
C551 B.n277 VSUBS 0.006571f
C552 B.n278 VSUBS 0.006571f
C553 B.n279 VSUBS 0.006571f
C554 B.n280 VSUBS 0.006571f
C555 B.n281 VSUBS 0.006571f
C556 B.n282 VSUBS 0.006571f
C557 B.n283 VSUBS 0.006571f
C558 B.n284 VSUBS 0.006571f
C559 B.n285 VSUBS 0.006571f
C560 B.n286 VSUBS 0.006571f
C561 B.n287 VSUBS 0.006571f
C562 B.n288 VSUBS 0.006571f
C563 B.n289 VSUBS 0.004542f
C564 B.n290 VSUBS 0.006571f
C565 B.n291 VSUBS 0.006571f
C566 B.n292 VSUBS 0.005315f
C567 B.n293 VSUBS 0.006571f
C568 B.n294 VSUBS 0.006571f
C569 B.n295 VSUBS 0.006571f
C570 B.n296 VSUBS 0.006571f
C571 B.n297 VSUBS 0.006571f
C572 B.n298 VSUBS 0.006571f
C573 B.n299 VSUBS 0.006571f
C574 B.n300 VSUBS 0.006571f
C575 B.n301 VSUBS 0.006571f
C576 B.n302 VSUBS 0.006571f
C577 B.n303 VSUBS 0.006571f
C578 B.n304 VSUBS 0.005315f
C579 B.n305 VSUBS 0.015225f
C580 B.n306 VSUBS 0.004542f
C581 B.n307 VSUBS 0.006571f
C582 B.n308 VSUBS 0.006571f
C583 B.n309 VSUBS 0.006571f
C584 B.n310 VSUBS 0.006571f
C585 B.n311 VSUBS 0.006571f
C586 B.n312 VSUBS 0.006571f
C587 B.n313 VSUBS 0.006571f
C588 B.n314 VSUBS 0.006571f
C589 B.n315 VSUBS 0.006571f
C590 B.n316 VSUBS 0.006571f
C591 B.n317 VSUBS 0.006571f
C592 B.n318 VSUBS 0.006571f
C593 B.n319 VSUBS 0.006571f
C594 B.n320 VSUBS 0.006571f
C595 B.n321 VSUBS 0.006571f
C596 B.n322 VSUBS 0.006571f
C597 B.n323 VSUBS 0.006571f
C598 B.n324 VSUBS 0.006571f
C599 B.n325 VSUBS 0.006571f
C600 B.n326 VSUBS 0.006571f
C601 B.n327 VSUBS 0.006571f
C602 B.n328 VSUBS 0.006571f
C603 B.n329 VSUBS 0.006571f
C604 B.n330 VSUBS 0.006571f
C605 B.n331 VSUBS 0.006571f
C606 B.n332 VSUBS 0.006571f
C607 B.n333 VSUBS 0.006571f
C608 B.n334 VSUBS 0.006571f
C609 B.n335 VSUBS 0.006571f
C610 B.n336 VSUBS 0.006571f
C611 B.n337 VSUBS 0.015222f
C612 B.n338 VSUBS 0.015222f
C613 B.n339 VSUBS 0.014929f
C614 B.n340 VSUBS 0.006571f
C615 B.n341 VSUBS 0.006571f
C616 B.n342 VSUBS 0.006571f
C617 B.n343 VSUBS 0.006571f
C618 B.n344 VSUBS 0.006571f
C619 B.n345 VSUBS 0.006571f
C620 B.n346 VSUBS 0.006571f
C621 B.n347 VSUBS 0.006571f
C622 B.n348 VSUBS 0.006571f
C623 B.n349 VSUBS 0.006571f
C624 B.n350 VSUBS 0.006571f
C625 B.n351 VSUBS 0.006571f
C626 B.n352 VSUBS 0.006571f
C627 B.n353 VSUBS 0.006571f
C628 B.n354 VSUBS 0.006571f
C629 B.n355 VSUBS 0.006571f
C630 B.n356 VSUBS 0.006571f
C631 B.n357 VSUBS 0.006571f
C632 B.n358 VSUBS 0.006571f
C633 B.n359 VSUBS 0.006571f
C634 B.n360 VSUBS 0.006571f
C635 B.n361 VSUBS 0.006571f
C636 B.n362 VSUBS 0.006571f
C637 B.n363 VSUBS 0.008575f
C638 B.n364 VSUBS 0.009135f
C639 B.n365 VSUBS 0.018166f
.ends

