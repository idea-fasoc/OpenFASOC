# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_aoi21_1 0 0 ;
  SIZE 3.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 2.2 2.85 2.5 ;
      LAYER MET2 ;
        RECT 2.35 2.15 2.85 2.55 ;
      LAYER VIA12 ;
        RECT 2.47 2.22 2.73 2.48 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.9 6.15 ;
        RECT 1.4 4.25 1.65 6.15 ;
      LAYER MET2 ;
        RECT 2.85 5.6 3.35 5.9 ;
        RECT 2.9 5.55 3.3 5.95 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
        RECT 2.97 5.62 3.23 5.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.95 0 3.2 1.4 ;
        RECT 0.7 0 0.95 1.8 ;
      LAYER MET2 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 3.5 3.5 3.8 ;
        RECT 3.1 1.65 3.35 5.2 ;
        RECT 2.1 1.65 3.35 1.9 ;
        RECT 2.1 0.95 2.35 1.9 ;
      LAYER MET2 ;
        RECT 3 3.45 3.5 3.85 ;
      LAYER VIA12 ;
        RECT 3.12 3.52 3.38 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.25 3.75 2.5 5.2 ;
      RECT 0.55 3.75 0.8 5.2 ;
      RECT 0.55 3.75 2.5 4 ;
  END
END gf180mcu_osu_sc_9T_aoi21_1
