* NGSPICE file created from diff_pair_sample_0203.ext - technology: sky130A

.subckt diff_pair_sample_0203 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=0 ps=0 w=3.01 l=0.25
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=1.1739 ps=6.8 w=3.01 l=0.25
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=1.1739 ps=6.8 w=3.01 l=0.25
X3 VDD1.t0 VP.t1 VTAIL.t2 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=1.1739 ps=6.8 w=3.01 l=0.25
X4 B.t8 B.t6 B.t7 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=0 ps=0 w=3.01 l=0.25
X5 B.t5 B.t3 B.t4 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=0 ps=0 w=3.01 l=0.25
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=1.1739 ps=6.8 w=3.01 l=0.25
X7 B.t2 B.t0 B.t1 w_n1202_n1574# sky130_fd_pr__pfet_01v8 ad=1.1739 pd=6.8 as=0 ps=0 w=3.01 l=0.25
R0 B.n149 B.n44 585
R1 B.n148 B.n147 585
R2 B.n146 B.n45 585
R3 B.n145 B.n144 585
R4 B.n143 B.n46 585
R5 B.n142 B.n141 585
R6 B.n140 B.n47 585
R7 B.n139 B.n138 585
R8 B.n137 B.n48 585
R9 B.n136 B.n135 585
R10 B.n134 B.n49 585
R11 B.n133 B.n132 585
R12 B.n131 B.n50 585
R13 B.n130 B.n129 585
R14 B.n128 B.n51 585
R15 B.n126 B.n125 585
R16 B.n124 B.n54 585
R17 B.n123 B.n122 585
R18 B.n121 B.n55 585
R19 B.n120 B.n119 585
R20 B.n118 B.n56 585
R21 B.n117 B.n116 585
R22 B.n115 B.n57 585
R23 B.n114 B.n113 585
R24 B.n112 B.n58 585
R25 B.n111 B.n110 585
R26 B.n106 B.n59 585
R27 B.n105 B.n104 585
R28 B.n103 B.n60 585
R29 B.n102 B.n101 585
R30 B.n100 B.n61 585
R31 B.n99 B.n98 585
R32 B.n97 B.n62 585
R33 B.n96 B.n95 585
R34 B.n94 B.n63 585
R35 B.n93 B.n92 585
R36 B.n91 B.n64 585
R37 B.n90 B.n89 585
R38 B.n88 B.n65 585
R39 B.n87 B.n86 585
R40 B.n151 B.n150 585
R41 B.n152 B.n43 585
R42 B.n154 B.n153 585
R43 B.n155 B.n42 585
R44 B.n157 B.n156 585
R45 B.n158 B.n41 585
R46 B.n160 B.n159 585
R47 B.n161 B.n40 585
R48 B.n163 B.n162 585
R49 B.n164 B.n39 585
R50 B.n166 B.n165 585
R51 B.n167 B.n38 585
R52 B.n169 B.n168 585
R53 B.n170 B.n37 585
R54 B.n172 B.n171 585
R55 B.n173 B.n36 585
R56 B.n175 B.n174 585
R57 B.n176 B.n35 585
R58 B.n178 B.n177 585
R59 B.n179 B.n34 585
R60 B.n181 B.n180 585
R61 B.n182 B.n33 585
R62 B.n184 B.n183 585
R63 B.n185 B.n32 585
R64 B.n247 B.n246 585
R65 B.n245 B.n8 585
R66 B.n244 B.n243 585
R67 B.n242 B.n9 585
R68 B.n241 B.n240 585
R69 B.n239 B.n10 585
R70 B.n238 B.n237 585
R71 B.n236 B.n11 585
R72 B.n235 B.n234 585
R73 B.n233 B.n12 585
R74 B.n232 B.n231 585
R75 B.n230 B.n13 585
R76 B.n229 B.n228 585
R77 B.n227 B.n14 585
R78 B.n226 B.n225 585
R79 B.n223 B.n15 585
R80 B.n222 B.n221 585
R81 B.n220 B.n18 585
R82 B.n219 B.n218 585
R83 B.n217 B.n19 585
R84 B.n216 B.n215 585
R85 B.n214 B.n20 585
R86 B.n213 B.n212 585
R87 B.n211 B.n21 585
R88 B.n210 B.n209 585
R89 B.n208 B.n207 585
R90 B.n206 B.n25 585
R91 B.n205 B.n204 585
R92 B.n203 B.n26 585
R93 B.n202 B.n201 585
R94 B.n200 B.n27 585
R95 B.n199 B.n198 585
R96 B.n197 B.n28 585
R97 B.n196 B.n195 585
R98 B.n194 B.n29 585
R99 B.n193 B.n192 585
R100 B.n191 B.n30 585
R101 B.n190 B.n189 585
R102 B.n188 B.n31 585
R103 B.n187 B.n186 585
R104 B.n248 B.n7 585
R105 B.n250 B.n249 585
R106 B.n251 B.n6 585
R107 B.n253 B.n252 585
R108 B.n254 B.n5 585
R109 B.n256 B.n255 585
R110 B.n257 B.n4 585
R111 B.n259 B.n258 585
R112 B.n260 B.n3 585
R113 B.n262 B.n261 585
R114 B.n263 B.n0 585
R115 B.n2 B.n1 585
R116 B.n72 B.n71 585
R117 B.n73 B.n70 585
R118 B.n75 B.n74 585
R119 B.n76 B.n69 585
R120 B.n78 B.n77 585
R121 B.n79 B.n68 585
R122 B.n81 B.n80 585
R123 B.n82 B.n67 585
R124 B.n84 B.n83 585
R125 B.n85 B.n66 585
R126 B.n107 B.t3 514.465
R127 B.n52 B.t6 514.465
R128 B.n22 B.t9 514.465
R129 B.n16 B.t0 514.465
R130 B.n86 B.n85 506.916
R131 B.n150 B.n149 506.916
R132 B.n186 B.n185 506.916
R133 B.n246 B.n7 506.916
R134 B.n265 B.n264 256.663
R135 B.n264 B.n263 235.042
R136 B.n264 B.n2 235.042
R137 B.n86 B.n65 163.367
R138 B.n90 B.n65 163.367
R139 B.n91 B.n90 163.367
R140 B.n92 B.n91 163.367
R141 B.n92 B.n63 163.367
R142 B.n96 B.n63 163.367
R143 B.n97 B.n96 163.367
R144 B.n98 B.n97 163.367
R145 B.n98 B.n61 163.367
R146 B.n102 B.n61 163.367
R147 B.n103 B.n102 163.367
R148 B.n104 B.n103 163.367
R149 B.n104 B.n59 163.367
R150 B.n111 B.n59 163.367
R151 B.n112 B.n111 163.367
R152 B.n113 B.n112 163.367
R153 B.n113 B.n57 163.367
R154 B.n117 B.n57 163.367
R155 B.n118 B.n117 163.367
R156 B.n119 B.n118 163.367
R157 B.n119 B.n55 163.367
R158 B.n123 B.n55 163.367
R159 B.n124 B.n123 163.367
R160 B.n125 B.n124 163.367
R161 B.n125 B.n51 163.367
R162 B.n130 B.n51 163.367
R163 B.n131 B.n130 163.367
R164 B.n132 B.n131 163.367
R165 B.n132 B.n49 163.367
R166 B.n136 B.n49 163.367
R167 B.n137 B.n136 163.367
R168 B.n138 B.n137 163.367
R169 B.n138 B.n47 163.367
R170 B.n142 B.n47 163.367
R171 B.n143 B.n142 163.367
R172 B.n144 B.n143 163.367
R173 B.n144 B.n45 163.367
R174 B.n148 B.n45 163.367
R175 B.n149 B.n148 163.367
R176 B.n185 B.n184 163.367
R177 B.n184 B.n33 163.367
R178 B.n180 B.n33 163.367
R179 B.n180 B.n179 163.367
R180 B.n179 B.n178 163.367
R181 B.n178 B.n35 163.367
R182 B.n174 B.n35 163.367
R183 B.n174 B.n173 163.367
R184 B.n173 B.n172 163.367
R185 B.n172 B.n37 163.367
R186 B.n168 B.n37 163.367
R187 B.n168 B.n167 163.367
R188 B.n167 B.n166 163.367
R189 B.n166 B.n39 163.367
R190 B.n162 B.n39 163.367
R191 B.n162 B.n161 163.367
R192 B.n161 B.n160 163.367
R193 B.n160 B.n41 163.367
R194 B.n156 B.n41 163.367
R195 B.n156 B.n155 163.367
R196 B.n155 B.n154 163.367
R197 B.n154 B.n43 163.367
R198 B.n150 B.n43 163.367
R199 B.n246 B.n245 163.367
R200 B.n245 B.n244 163.367
R201 B.n244 B.n9 163.367
R202 B.n240 B.n9 163.367
R203 B.n240 B.n239 163.367
R204 B.n239 B.n238 163.367
R205 B.n238 B.n11 163.367
R206 B.n234 B.n11 163.367
R207 B.n234 B.n233 163.367
R208 B.n233 B.n232 163.367
R209 B.n232 B.n13 163.367
R210 B.n228 B.n13 163.367
R211 B.n228 B.n227 163.367
R212 B.n227 B.n226 163.367
R213 B.n226 B.n15 163.367
R214 B.n221 B.n15 163.367
R215 B.n221 B.n220 163.367
R216 B.n220 B.n219 163.367
R217 B.n219 B.n19 163.367
R218 B.n215 B.n19 163.367
R219 B.n215 B.n214 163.367
R220 B.n214 B.n213 163.367
R221 B.n213 B.n21 163.367
R222 B.n209 B.n21 163.367
R223 B.n209 B.n208 163.367
R224 B.n208 B.n25 163.367
R225 B.n204 B.n25 163.367
R226 B.n204 B.n203 163.367
R227 B.n203 B.n202 163.367
R228 B.n202 B.n27 163.367
R229 B.n198 B.n27 163.367
R230 B.n198 B.n197 163.367
R231 B.n197 B.n196 163.367
R232 B.n196 B.n29 163.367
R233 B.n192 B.n29 163.367
R234 B.n192 B.n191 163.367
R235 B.n191 B.n190 163.367
R236 B.n190 B.n31 163.367
R237 B.n186 B.n31 163.367
R238 B.n250 B.n7 163.367
R239 B.n251 B.n250 163.367
R240 B.n252 B.n251 163.367
R241 B.n252 B.n5 163.367
R242 B.n256 B.n5 163.367
R243 B.n257 B.n256 163.367
R244 B.n258 B.n257 163.367
R245 B.n258 B.n3 163.367
R246 B.n262 B.n3 163.367
R247 B.n263 B.n262 163.367
R248 B.n72 B.n2 163.367
R249 B.n73 B.n72 163.367
R250 B.n74 B.n73 163.367
R251 B.n74 B.n69 163.367
R252 B.n78 B.n69 163.367
R253 B.n79 B.n78 163.367
R254 B.n80 B.n79 163.367
R255 B.n80 B.n67 163.367
R256 B.n84 B.n67 163.367
R257 B.n85 B.n84 163.367
R258 B.n52 B.t7 156.63
R259 B.n22 B.t11 156.63
R260 B.n107 B.t4 156.627
R261 B.n16 B.t2 156.627
R262 B.n53 B.t8 145.381
R263 B.n23 B.t10 145.381
R264 B.n108 B.t5 145.38
R265 B.n17 B.t1 145.38
R266 B.n109 B.n108 59.5399
R267 B.n127 B.n53 59.5399
R268 B.n24 B.n23 59.5399
R269 B.n224 B.n17 59.5399
R270 B.n248 B.n247 32.9371
R271 B.n187 B.n32 32.9371
R272 B.n151 B.n44 32.9371
R273 B.n87 B.n66 32.9371
R274 B B.n265 18.0485
R275 B.n108 B.n107 11.249
R276 B.n53 B.n52 11.249
R277 B.n23 B.n22 11.249
R278 B.n17 B.n16 11.249
R279 B.n249 B.n248 10.6151
R280 B.n249 B.n6 10.6151
R281 B.n253 B.n6 10.6151
R282 B.n254 B.n253 10.6151
R283 B.n255 B.n254 10.6151
R284 B.n255 B.n4 10.6151
R285 B.n259 B.n4 10.6151
R286 B.n260 B.n259 10.6151
R287 B.n261 B.n260 10.6151
R288 B.n261 B.n0 10.6151
R289 B.n247 B.n8 10.6151
R290 B.n243 B.n8 10.6151
R291 B.n243 B.n242 10.6151
R292 B.n242 B.n241 10.6151
R293 B.n241 B.n10 10.6151
R294 B.n237 B.n10 10.6151
R295 B.n237 B.n236 10.6151
R296 B.n236 B.n235 10.6151
R297 B.n235 B.n12 10.6151
R298 B.n231 B.n12 10.6151
R299 B.n231 B.n230 10.6151
R300 B.n230 B.n229 10.6151
R301 B.n229 B.n14 10.6151
R302 B.n225 B.n14 10.6151
R303 B.n223 B.n222 10.6151
R304 B.n222 B.n18 10.6151
R305 B.n218 B.n18 10.6151
R306 B.n218 B.n217 10.6151
R307 B.n217 B.n216 10.6151
R308 B.n216 B.n20 10.6151
R309 B.n212 B.n20 10.6151
R310 B.n212 B.n211 10.6151
R311 B.n211 B.n210 10.6151
R312 B.n207 B.n206 10.6151
R313 B.n206 B.n205 10.6151
R314 B.n205 B.n26 10.6151
R315 B.n201 B.n26 10.6151
R316 B.n201 B.n200 10.6151
R317 B.n200 B.n199 10.6151
R318 B.n199 B.n28 10.6151
R319 B.n195 B.n28 10.6151
R320 B.n195 B.n194 10.6151
R321 B.n194 B.n193 10.6151
R322 B.n193 B.n30 10.6151
R323 B.n189 B.n30 10.6151
R324 B.n189 B.n188 10.6151
R325 B.n188 B.n187 10.6151
R326 B.n183 B.n32 10.6151
R327 B.n183 B.n182 10.6151
R328 B.n182 B.n181 10.6151
R329 B.n181 B.n34 10.6151
R330 B.n177 B.n34 10.6151
R331 B.n177 B.n176 10.6151
R332 B.n176 B.n175 10.6151
R333 B.n175 B.n36 10.6151
R334 B.n171 B.n36 10.6151
R335 B.n171 B.n170 10.6151
R336 B.n170 B.n169 10.6151
R337 B.n169 B.n38 10.6151
R338 B.n165 B.n38 10.6151
R339 B.n165 B.n164 10.6151
R340 B.n164 B.n163 10.6151
R341 B.n163 B.n40 10.6151
R342 B.n159 B.n40 10.6151
R343 B.n159 B.n158 10.6151
R344 B.n158 B.n157 10.6151
R345 B.n157 B.n42 10.6151
R346 B.n153 B.n42 10.6151
R347 B.n153 B.n152 10.6151
R348 B.n152 B.n151 10.6151
R349 B.n71 B.n1 10.6151
R350 B.n71 B.n70 10.6151
R351 B.n75 B.n70 10.6151
R352 B.n76 B.n75 10.6151
R353 B.n77 B.n76 10.6151
R354 B.n77 B.n68 10.6151
R355 B.n81 B.n68 10.6151
R356 B.n82 B.n81 10.6151
R357 B.n83 B.n82 10.6151
R358 B.n83 B.n66 10.6151
R359 B.n88 B.n87 10.6151
R360 B.n89 B.n88 10.6151
R361 B.n89 B.n64 10.6151
R362 B.n93 B.n64 10.6151
R363 B.n94 B.n93 10.6151
R364 B.n95 B.n94 10.6151
R365 B.n95 B.n62 10.6151
R366 B.n99 B.n62 10.6151
R367 B.n100 B.n99 10.6151
R368 B.n101 B.n100 10.6151
R369 B.n101 B.n60 10.6151
R370 B.n105 B.n60 10.6151
R371 B.n106 B.n105 10.6151
R372 B.n110 B.n106 10.6151
R373 B.n114 B.n58 10.6151
R374 B.n115 B.n114 10.6151
R375 B.n116 B.n115 10.6151
R376 B.n116 B.n56 10.6151
R377 B.n120 B.n56 10.6151
R378 B.n121 B.n120 10.6151
R379 B.n122 B.n121 10.6151
R380 B.n122 B.n54 10.6151
R381 B.n126 B.n54 10.6151
R382 B.n129 B.n128 10.6151
R383 B.n129 B.n50 10.6151
R384 B.n133 B.n50 10.6151
R385 B.n134 B.n133 10.6151
R386 B.n135 B.n134 10.6151
R387 B.n135 B.n48 10.6151
R388 B.n139 B.n48 10.6151
R389 B.n140 B.n139 10.6151
R390 B.n141 B.n140 10.6151
R391 B.n141 B.n46 10.6151
R392 B.n145 B.n46 10.6151
R393 B.n146 B.n145 10.6151
R394 B.n147 B.n146 10.6151
R395 B.n147 B.n44 10.6151
R396 B.n225 B.n224 8.74196
R397 B.n207 B.n24 8.74196
R398 B.n110 B.n109 8.74196
R399 B.n128 B.n127 8.74196
R400 B.n265 B.n0 8.11757
R401 B.n265 B.n1 8.11757
R402 B.n224 B.n223 1.87367
R403 B.n210 B.n24 1.87367
R404 B.n109 B.n58 1.87367
R405 B.n127 B.n126 1.87367
R406 VP.n0 VP.t1 633.477
R407 VP.n0 VP.t0 601.848
R408 VP VP.n0 0.0516364
R409 VTAIL.n2 VTAIL.t2 131.276
R410 VTAIL.n1 VTAIL.t0 131.276
R411 VTAIL.n3 VTAIL.t1 131.275
R412 VTAIL.n0 VTAIL.t3 131.275
R413 VTAIL.n1 VTAIL.n0 15.9789
R414 VTAIL.n3 VTAIL.n2 15.4789
R415 VTAIL.n2 VTAIL.n1 0.720328
R416 VTAIL VTAIL.n0 0.653517
R417 VTAIL VTAIL.n3 0.0673103
R418 VDD1 VDD1.t1 175.876
R419 VDD1 VDD1.t0 148.138
R420 VN VN.t1 633.857
R421 VN VN.t0 601.899
R422 VDD2.n0 VDD2.t1 175.226
R423 VDD2.n0 VDD2.t0 147.954
R424 VDD2 VDD2.n0 0.18369
C0 B VDD2 0.711288f
C1 B VN 0.538367f
C2 VTAIL B 0.923608f
C3 VDD1 VDD2 0.419075f
C4 B w_n1202_n1574# 3.76896f
C5 VDD1 VN 0.153399f
C6 VTAIL VDD1 2.64848f
C7 VP VDD2 0.240179f
C8 VP VN 2.70426f
C9 VDD1 w_n1202_n1574# 0.839435f
C10 VTAIL VP 0.419324f
C11 VP w_n1202_n1574# 1.45267f
C12 VDD2 VN 0.512367f
C13 VTAIL VDD2 2.68383f
C14 VDD1 B 0.699611f
C15 VTAIL VN 0.405048f
C16 VDD2 w_n1202_n1574# 0.839151f
C17 VN w_n1202_n1574# 1.30694f
C18 B VP 0.771911f
C19 VTAIL w_n1202_n1574# 1.39539f
C20 VDD1 VP 0.597383f
C21 VDD2 VSUBS 0.398605f
C22 VDD1 VSUBS 2.324562f
C23 VTAIL VSUBS 0.138294f
C24 VN VSUBS 3.46131f
C25 VP VSUBS 0.585223f
C26 B VSUBS 1.347603f
C27 w_n1202_n1574# VSUBS 23.958302f
C28 VDD2.t1 VSUBS 0.473713f
C29 VDD2.t0 VSUBS 0.341887f
C30 VDD2.n0 VSUBS 1.85628f
C31 VN.t0 VSUBS 0.121394f
C32 VN.t1 VSUBS 0.182005f
C33 VDD1.t0 VSUBS 0.320914f
C34 VDD1.t1 VSUBS 0.453337f
C35 VTAIL.t3 VSUBS 0.36021f
C36 VTAIL.n0 VSUBS 0.978502f
C37 VTAIL.t0 VSUBS 0.360211f
C38 VTAIL.n1 VSUBS 0.983501f
C39 VTAIL.t2 VSUBS 0.360211f
C40 VTAIL.n2 VSUBS 0.946077f
C41 VTAIL.t1 VSUBS 0.36021f
C42 VTAIL.n3 VSUBS 0.897202f
C43 VP.t1 VSUBS 0.184223f
C44 VP.t0 VSUBS 0.124397f
C45 VP.n0 VSUBS 2.38565f
C46 B.n0 VSUBS 0.007371f
C47 B.n1 VSUBS 0.007371f
C48 B.n2 VSUBS 0.010902f
C49 B.n3 VSUBS 0.008354f
C50 B.n4 VSUBS 0.008354f
C51 B.n5 VSUBS 0.008354f
C52 B.n6 VSUBS 0.008354f
C53 B.n7 VSUBS 0.019192f
C54 B.n8 VSUBS 0.008354f
C55 B.n9 VSUBS 0.008354f
C56 B.n10 VSUBS 0.008354f
C57 B.n11 VSUBS 0.008354f
C58 B.n12 VSUBS 0.008354f
C59 B.n13 VSUBS 0.008354f
C60 B.n14 VSUBS 0.008354f
C61 B.n15 VSUBS 0.008354f
C62 B.t1 VSUBS 0.08627f
C63 B.t2 VSUBS 0.090197f
C64 B.t0 VSUBS 0.038455f
C65 B.n16 VSUBS 0.069663f
C66 B.n17 VSUBS 0.066603f
C67 B.n18 VSUBS 0.008354f
C68 B.n19 VSUBS 0.008354f
C69 B.n20 VSUBS 0.008354f
C70 B.n21 VSUBS 0.008354f
C71 B.t10 VSUBS 0.08627f
C72 B.t11 VSUBS 0.090197f
C73 B.t9 VSUBS 0.038455f
C74 B.n22 VSUBS 0.069663f
C75 B.n23 VSUBS 0.066602f
C76 B.n24 VSUBS 0.019356f
C77 B.n25 VSUBS 0.008354f
C78 B.n26 VSUBS 0.008354f
C79 B.n27 VSUBS 0.008354f
C80 B.n28 VSUBS 0.008354f
C81 B.n29 VSUBS 0.008354f
C82 B.n30 VSUBS 0.008354f
C83 B.n31 VSUBS 0.008354f
C84 B.n32 VSUBS 0.019192f
C85 B.n33 VSUBS 0.008354f
C86 B.n34 VSUBS 0.008354f
C87 B.n35 VSUBS 0.008354f
C88 B.n36 VSUBS 0.008354f
C89 B.n37 VSUBS 0.008354f
C90 B.n38 VSUBS 0.008354f
C91 B.n39 VSUBS 0.008354f
C92 B.n40 VSUBS 0.008354f
C93 B.n41 VSUBS 0.008354f
C94 B.n42 VSUBS 0.008354f
C95 B.n43 VSUBS 0.008354f
C96 B.n44 VSUBS 0.019144f
C97 B.n45 VSUBS 0.008354f
C98 B.n46 VSUBS 0.008354f
C99 B.n47 VSUBS 0.008354f
C100 B.n48 VSUBS 0.008354f
C101 B.n49 VSUBS 0.008354f
C102 B.n50 VSUBS 0.008354f
C103 B.n51 VSUBS 0.008354f
C104 B.t8 VSUBS 0.08627f
C105 B.t7 VSUBS 0.090197f
C106 B.t6 VSUBS 0.038455f
C107 B.n52 VSUBS 0.069663f
C108 B.n53 VSUBS 0.066602f
C109 B.n54 VSUBS 0.008354f
C110 B.n55 VSUBS 0.008354f
C111 B.n56 VSUBS 0.008354f
C112 B.n57 VSUBS 0.008354f
C113 B.n58 VSUBS 0.004914f
C114 B.n59 VSUBS 0.008354f
C115 B.n60 VSUBS 0.008354f
C116 B.n61 VSUBS 0.008354f
C117 B.n62 VSUBS 0.008354f
C118 B.n63 VSUBS 0.008354f
C119 B.n64 VSUBS 0.008354f
C120 B.n65 VSUBS 0.008354f
C121 B.n66 VSUBS 0.019192f
C122 B.n67 VSUBS 0.008354f
C123 B.n68 VSUBS 0.008354f
C124 B.n69 VSUBS 0.008354f
C125 B.n70 VSUBS 0.008354f
C126 B.n71 VSUBS 0.008354f
C127 B.n72 VSUBS 0.008354f
C128 B.n73 VSUBS 0.008354f
C129 B.n74 VSUBS 0.008354f
C130 B.n75 VSUBS 0.008354f
C131 B.n76 VSUBS 0.008354f
C132 B.n77 VSUBS 0.008354f
C133 B.n78 VSUBS 0.008354f
C134 B.n79 VSUBS 0.008354f
C135 B.n80 VSUBS 0.008354f
C136 B.n81 VSUBS 0.008354f
C137 B.n82 VSUBS 0.008354f
C138 B.n83 VSUBS 0.008354f
C139 B.n84 VSUBS 0.008354f
C140 B.n85 VSUBS 0.019192f
C141 B.n86 VSUBS 0.020123f
C142 B.n87 VSUBS 0.020123f
C143 B.n88 VSUBS 0.008354f
C144 B.n89 VSUBS 0.008354f
C145 B.n90 VSUBS 0.008354f
C146 B.n91 VSUBS 0.008354f
C147 B.n92 VSUBS 0.008354f
C148 B.n93 VSUBS 0.008354f
C149 B.n94 VSUBS 0.008354f
C150 B.n95 VSUBS 0.008354f
C151 B.n96 VSUBS 0.008354f
C152 B.n97 VSUBS 0.008354f
C153 B.n98 VSUBS 0.008354f
C154 B.n99 VSUBS 0.008354f
C155 B.n100 VSUBS 0.008354f
C156 B.n101 VSUBS 0.008354f
C157 B.n102 VSUBS 0.008354f
C158 B.n103 VSUBS 0.008354f
C159 B.n104 VSUBS 0.008354f
C160 B.n105 VSUBS 0.008354f
C161 B.n106 VSUBS 0.008354f
C162 B.t5 VSUBS 0.08627f
C163 B.t4 VSUBS 0.090197f
C164 B.t3 VSUBS 0.038455f
C165 B.n107 VSUBS 0.069663f
C166 B.n108 VSUBS 0.066603f
C167 B.n109 VSUBS 0.019356f
C168 B.n110 VSUBS 0.007617f
C169 B.n111 VSUBS 0.008354f
C170 B.n112 VSUBS 0.008354f
C171 B.n113 VSUBS 0.008354f
C172 B.n114 VSUBS 0.008354f
C173 B.n115 VSUBS 0.008354f
C174 B.n116 VSUBS 0.008354f
C175 B.n117 VSUBS 0.008354f
C176 B.n118 VSUBS 0.008354f
C177 B.n119 VSUBS 0.008354f
C178 B.n120 VSUBS 0.008354f
C179 B.n121 VSUBS 0.008354f
C180 B.n122 VSUBS 0.008354f
C181 B.n123 VSUBS 0.008354f
C182 B.n124 VSUBS 0.008354f
C183 B.n125 VSUBS 0.008354f
C184 B.n126 VSUBS 0.004914f
C185 B.n127 VSUBS 0.019356f
C186 B.n128 VSUBS 0.007617f
C187 B.n129 VSUBS 0.008354f
C188 B.n130 VSUBS 0.008354f
C189 B.n131 VSUBS 0.008354f
C190 B.n132 VSUBS 0.008354f
C191 B.n133 VSUBS 0.008354f
C192 B.n134 VSUBS 0.008354f
C193 B.n135 VSUBS 0.008354f
C194 B.n136 VSUBS 0.008354f
C195 B.n137 VSUBS 0.008354f
C196 B.n138 VSUBS 0.008354f
C197 B.n139 VSUBS 0.008354f
C198 B.n140 VSUBS 0.008354f
C199 B.n141 VSUBS 0.008354f
C200 B.n142 VSUBS 0.008354f
C201 B.n143 VSUBS 0.008354f
C202 B.n144 VSUBS 0.008354f
C203 B.n145 VSUBS 0.008354f
C204 B.n146 VSUBS 0.008354f
C205 B.n147 VSUBS 0.008354f
C206 B.n148 VSUBS 0.008354f
C207 B.n149 VSUBS 0.020123f
C208 B.n150 VSUBS 0.019192f
C209 B.n151 VSUBS 0.020171f
C210 B.n152 VSUBS 0.008354f
C211 B.n153 VSUBS 0.008354f
C212 B.n154 VSUBS 0.008354f
C213 B.n155 VSUBS 0.008354f
C214 B.n156 VSUBS 0.008354f
C215 B.n157 VSUBS 0.008354f
C216 B.n158 VSUBS 0.008354f
C217 B.n159 VSUBS 0.008354f
C218 B.n160 VSUBS 0.008354f
C219 B.n161 VSUBS 0.008354f
C220 B.n162 VSUBS 0.008354f
C221 B.n163 VSUBS 0.008354f
C222 B.n164 VSUBS 0.008354f
C223 B.n165 VSUBS 0.008354f
C224 B.n166 VSUBS 0.008354f
C225 B.n167 VSUBS 0.008354f
C226 B.n168 VSUBS 0.008354f
C227 B.n169 VSUBS 0.008354f
C228 B.n170 VSUBS 0.008354f
C229 B.n171 VSUBS 0.008354f
C230 B.n172 VSUBS 0.008354f
C231 B.n173 VSUBS 0.008354f
C232 B.n174 VSUBS 0.008354f
C233 B.n175 VSUBS 0.008354f
C234 B.n176 VSUBS 0.008354f
C235 B.n177 VSUBS 0.008354f
C236 B.n178 VSUBS 0.008354f
C237 B.n179 VSUBS 0.008354f
C238 B.n180 VSUBS 0.008354f
C239 B.n181 VSUBS 0.008354f
C240 B.n182 VSUBS 0.008354f
C241 B.n183 VSUBS 0.008354f
C242 B.n184 VSUBS 0.008354f
C243 B.n185 VSUBS 0.019192f
C244 B.n186 VSUBS 0.020123f
C245 B.n187 VSUBS 0.020123f
C246 B.n188 VSUBS 0.008354f
C247 B.n189 VSUBS 0.008354f
C248 B.n190 VSUBS 0.008354f
C249 B.n191 VSUBS 0.008354f
C250 B.n192 VSUBS 0.008354f
C251 B.n193 VSUBS 0.008354f
C252 B.n194 VSUBS 0.008354f
C253 B.n195 VSUBS 0.008354f
C254 B.n196 VSUBS 0.008354f
C255 B.n197 VSUBS 0.008354f
C256 B.n198 VSUBS 0.008354f
C257 B.n199 VSUBS 0.008354f
C258 B.n200 VSUBS 0.008354f
C259 B.n201 VSUBS 0.008354f
C260 B.n202 VSUBS 0.008354f
C261 B.n203 VSUBS 0.008354f
C262 B.n204 VSUBS 0.008354f
C263 B.n205 VSUBS 0.008354f
C264 B.n206 VSUBS 0.008354f
C265 B.n207 VSUBS 0.007617f
C266 B.n208 VSUBS 0.008354f
C267 B.n209 VSUBS 0.008354f
C268 B.n210 VSUBS 0.004914f
C269 B.n211 VSUBS 0.008354f
C270 B.n212 VSUBS 0.008354f
C271 B.n213 VSUBS 0.008354f
C272 B.n214 VSUBS 0.008354f
C273 B.n215 VSUBS 0.008354f
C274 B.n216 VSUBS 0.008354f
C275 B.n217 VSUBS 0.008354f
C276 B.n218 VSUBS 0.008354f
C277 B.n219 VSUBS 0.008354f
C278 B.n220 VSUBS 0.008354f
C279 B.n221 VSUBS 0.008354f
C280 B.n222 VSUBS 0.008354f
C281 B.n223 VSUBS 0.004914f
C282 B.n224 VSUBS 0.019356f
C283 B.n225 VSUBS 0.007617f
C284 B.n226 VSUBS 0.008354f
C285 B.n227 VSUBS 0.008354f
C286 B.n228 VSUBS 0.008354f
C287 B.n229 VSUBS 0.008354f
C288 B.n230 VSUBS 0.008354f
C289 B.n231 VSUBS 0.008354f
C290 B.n232 VSUBS 0.008354f
C291 B.n233 VSUBS 0.008354f
C292 B.n234 VSUBS 0.008354f
C293 B.n235 VSUBS 0.008354f
C294 B.n236 VSUBS 0.008354f
C295 B.n237 VSUBS 0.008354f
C296 B.n238 VSUBS 0.008354f
C297 B.n239 VSUBS 0.008354f
C298 B.n240 VSUBS 0.008354f
C299 B.n241 VSUBS 0.008354f
C300 B.n242 VSUBS 0.008354f
C301 B.n243 VSUBS 0.008354f
C302 B.n244 VSUBS 0.008354f
C303 B.n245 VSUBS 0.008354f
C304 B.n246 VSUBS 0.020123f
C305 B.n247 VSUBS 0.020123f
C306 B.n248 VSUBS 0.019192f
C307 B.n249 VSUBS 0.008354f
C308 B.n250 VSUBS 0.008354f
C309 B.n251 VSUBS 0.008354f
C310 B.n252 VSUBS 0.008354f
C311 B.n253 VSUBS 0.008354f
C312 B.n254 VSUBS 0.008354f
C313 B.n255 VSUBS 0.008354f
C314 B.n256 VSUBS 0.008354f
C315 B.n257 VSUBS 0.008354f
C316 B.n258 VSUBS 0.008354f
C317 B.n259 VSUBS 0.008354f
C318 B.n260 VSUBS 0.008354f
C319 B.n261 VSUBS 0.008354f
C320 B.n262 VSUBS 0.008354f
C321 B.n263 VSUBS 0.010902f
C322 B.n264 VSUBS 0.011613f
C323 B.n265 VSUBS 0.023094f
.ends

