* NGSPICE file created from diff_pair_sample_0886.ext - technology: sky130A

.subckt diff_pair_sample_0886 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=0 ps=0 w=10.11 l=3.23
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=0 ps=0 w=10.11 l=3.23
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=0 ps=0 w=10.11 l=3.23
X3 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=3.9429 ps=21 w=10.11 l=3.23
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=0 ps=0 w=10.11 l=3.23
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=3.9429 ps=21 w=10.11 l=3.23
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=3.9429 ps=21 w=10.11 l=3.23
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.9429 pd=21 as=3.9429 ps=21 w=10.11 l=3.23
R0 B.n655 B.n654 585
R1 B.n263 B.n96 585
R2 B.n262 B.n261 585
R3 B.n260 B.n259 585
R4 B.n258 B.n257 585
R5 B.n256 B.n255 585
R6 B.n254 B.n253 585
R7 B.n252 B.n251 585
R8 B.n250 B.n249 585
R9 B.n248 B.n247 585
R10 B.n246 B.n245 585
R11 B.n244 B.n243 585
R12 B.n242 B.n241 585
R13 B.n240 B.n239 585
R14 B.n238 B.n237 585
R15 B.n236 B.n235 585
R16 B.n234 B.n233 585
R17 B.n232 B.n231 585
R18 B.n230 B.n229 585
R19 B.n228 B.n227 585
R20 B.n226 B.n225 585
R21 B.n224 B.n223 585
R22 B.n222 B.n221 585
R23 B.n220 B.n219 585
R24 B.n218 B.n217 585
R25 B.n216 B.n215 585
R26 B.n214 B.n213 585
R27 B.n212 B.n211 585
R28 B.n210 B.n209 585
R29 B.n208 B.n207 585
R30 B.n206 B.n205 585
R31 B.n204 B.n203 585
R32 B.n202 B.n201 585
R33 B.n200 B.n199 585
R34 B.n198 B.n197 585
R35 B.n196 B.n195 585
R36 B.n194 B.n193 585
R37 B.n192 B.n191 585
R38 B.n190 B.n189 585
R39 B.n188 B.n187 585
R40 B.n186 B.n185 585
R41 B.n184 B.n183 585
R42 B.n182 B.n181 585
R43 B.n180 B.n179 585
R44 B.n178 B.n177 585
R45 B.n176 B.n175 585
R46 B.n174 B.n173 585
R47 B.n172 B.n171 585
R48 B.n170 B.n169 585
R49 B.n168 B.n167 585
R50 B.n166 B.n165 585
R51 B.n164 B.n163 585
R52 B.n162 B.n161 585
R53 B.n160 B.n159 585
R54 B.n158 B.n157 585
R55 B.n156 B.n155 585
R56 B.n154 B.n153 585
R57 B.n152 B.n151 585
R58 B.n150 B.n149 585
R59 B.n148 B.n147 585
R60 B.n146 B.n145 585
R61 B.n144 B.n143 585
R62 B.n142 B.n141 585
R63 B.n140 B.n139 585
R64 B.n138 B.n137 585
R65 B.n136 B.n135 585
R66 B.n134 B.n133 585
R67 B.n132 B.n131 585
R68 B.n130 B.n129 585
R69 B.n128 B.n127 585
R70 B.n126 B.n125 585
R71 B.n124 B.n123 585
R72 B.n122 B.n121 585
R73 B.n120 B.n119 585
R74 B.n118 B.n117 585
R75 B.n116 B.n115 585
R76 B.n114 B.n113 585
R77 B.n112 B.n111 585
R78 B.n110 B.n109 585
R79 B.n108 B.n107 585
R80 B.n106 B.n105 585
R81 B.n104 B.n103 585
R82 B.n653 B.n55 585
R83 B.n658 B.n55 585
R84 B.n652 B.n54 585
R85 B.n659 B.n54 585
R86 B.n651 B.n650 585
R87 B.n650 B.n50 585
R88 B.n649 B.n49 585
R89 B.n665 B.n49 585
R90 B.n648 B.n48 585
R91 B.n666 B.n48 585
R92 B.n647 B.n47 585
R93 B.n667 B.n47 585
R94 B.n646 B.n645 585
R95 B.n645 B.n43 585
R96 B.n644 B.n42 585
R97 B.n673 B.n42 585
R98 B.n643 B.n41 585
R99 B.n674 B.n41 585
R100 B.n642 B.n40 585
R101 B.n675 B.n40 585
R102 B.n641 B.n640 585
R103 B.n640 B.n36 585
R104 B.n639 B.n35 585
R105 B.n681 B.n35 585
R106 B.n638 B.n34 585
R107 B.n682 B.n34 585
R108 B.n637 B.n33 585
R109 B.n683 B.n33 585
R110 B.n636 B.n635 585
R111 B.n635 B.n29 585
R112 B.n634 B.n28 585
R113 B.n689 B.n28 585
R114 B.n633 B.n27 585
R115 B.n690 B.n27 585
R116 B.n632 B.n26 585
R117 B.n691 B.n26 585
R118 B.n631 B.n630 585
R119 B.n630 B.n22 585
R120 B.n629 B.n21 585
R121 B.n697 B.n21 585
R122 B.n628 B.n20 585
R123 B.n698 B.n20 585
R124 B.n627 B.n19 585
R125 B.n699 B.n19 585
R126 B.n626 B.n625 585
R127 B.n625 B.n18 585
R128 B.n624 B.n14 585
R129 B.n705 B.n14 585
R130 B.n623 B.n13 585
R131 B.n706 B.n13 585
R132 B.n622 B.n12 585
R133 B.n707 B.n12 585
R134 B.n621 B.n620 585
R135 B.n620 B.n8 585
R136 B.n619 B.n7 585
R137 B.n713 B.n7 585
R138 B.n618 B.n6 585
R139 B.n714 B.n6 585
R140 B.n617 B.n5 585
R141 B.n715 B.n5 585
R142 B.n616 B.n615 585
R143 B.n615 B.n4 585
R144 B.n614 B.n264 585
R145 B.n614 B.n613 585
R146 B.n604 B.n265 585
R147 B.n266 B.n265 585
R148 B.n606 B.n605 585
R149 B.n607 B.n606 585
R150 B.n603 B.n271 585
R151 B.n271 B.n270 585
R152 B.n602 B.n601 585
R153 B.n601 B.n600 585
R154 B.n273 B.n272 585
R155 B.n593 B.n273 585
R156 B.n592 B.n591 585
R157 B.n594 B.n592 585
R158 B.n590 B.n278 585
R159 B.n278 B.n277 585
R160 B.n589 B.n588 585
R161 B.n588 B.n587 585
R162 B.n280 B.n279 585
R163 B.n281 B.n280 585
R164 B.n580 B.n579 585
R165 B.n581 B.n580 585
R166 B.n578 B.n286 585
R167 B.n286 B.n285 585
R168 B.n577 B.n576 585
R169 B.n576 B.n575 585
R170 B.n288 B.n287 585
R171 B.n289 B.n288 585
R172 B.n568 B.n567 585
R173 B.n569 B.n568 585
R174 B.n566 B.n294 585
R175 B.n294 B.n293 585
R176 B.n565 B.n564 585
R177 B.n564 B.n563 585
R178 B.n296 B.n295 585
R179 B.n297 B.n296 585
R180 B.n556 B.n555 585
R181 B.n557 B.n556 585
R182 B.n554 B.n301 585
R183 B.n305 B.n301 585
R184 B.n553 B.n552 585
R185 B.n552 B.n551 585
R186 B.n303 B.n302 585
R187 B.n304 B.n303 585
R188 B.n544 B.n543 585
R189 B.n545 B.n544 585
R190 B.n542 B.n310 585
R191 B.n310 B.n309 585
R192 B.n541 B.n540 585
R193 B.n540 B.n539 585
R194 B.n312 B.n311 585
R195 B.n313 B.n312 585
R196 B.n532 B.n531 585
R197 B.n533 B.n532 585
R198 B.n530 B.n318 585
R199 B.n318 B.n317 585
R200 B.n525 B.n524 585
R201 B.n523 B.n361 585
R202 B.n522 B.n360 585
R203 B.n527 B.n360 585
R204 B.n521 B.n520 585
R205 B.n519 B.n518 585
R206 B.n517 B.n516 585
R207 B.n515 B.n514 585
R208 B.n513 B.n512 585
R209 B.n511 B.n510 585
R210 B.n509 B.n508 585
R211 B.n507 B.n506 585
R212 B.n505 B.n504 585
R213 B.n503 B.n502 585
R214 B.n501 B.n500 585
R215 B.n499 B.n498 585
R216 B.n497 B.n496 585
R217 B.n495 B.n494 585
R218 B.n493 B.n492 585
R219 B.n491 B.n490 585
R220 B.n489 B.n488 585
R221 B.n487 B.n486 585
R222 B.n485 B.n484 585
R223 B.n483 B.n482 585
R224 B.n481 B.n480 585
R225 B.n479 B.n478 585
R226 B.n477 B.n476 585
R227 B.n475 B.n474 585
R228 B.n473 B.n472 585
R229 B.n471 B.n470 585
R230 B.n469 B.n468 585
R231 B.n467 B.n466 585
R232 B.n465 B.n464 585
R233 B.n463 B.n462 585
R234 B.n461 B.n460 585
R235 B.n459 B.n458 585
R236 B.n457 B.n456 585
R237 B.n454 B.n453 585
R238 B.n452 B.n451 585
R239 B.n450 B.n449 585
R240 B.n448 B.n447 585
R241 B.n446 B.n445 585
R242 B.n444 B.n443 585
R243 B.n442 B.n441 585
R244 B.n440 B.n439 585
R245 B.n438 B.n437 585
R246 B.n436 B.n435 585
R247 B.n433 B.n432 585
R248 B.n431 B.n430 585
R249 B.n429 B.n428 585
R250 B.n427 B.n426 585
R251 B.n425 B.n424 585
R252 B.n423 B.n422 585
R253 B.n421 B.n420 585
R254 B.n419 B.n418 585
R255 B.n417 B.n416 585
R256 B.n415 B.n414 585
R257 B.n413 B.n412 585
R258 B.n411 B.n410 585
R259 B.n409 B.n408 585
R260 B.n407 B.n406 585
R261 B.n405 B.n404 585
R262 B.n403 B.n402 585
R263 B.n401 B.n400 585
R264 B.n399 B.n398 585
R265 B.n397 B.n396 585
R266 B.n395 B.n394 585
R267 B.n393 B.n392 585
R268 B.n391 B.n390 585
R269 B.n389 B.n388 585
R270 B.n387 B.n386 585
R271 B.n385 B.n384 585
R272 B.n383 B.n382 585
R273 B.n381 B.n380 585
R274 B.n379 B.n378 585
R275 B.n377 B.n376 585
R276 B.n375 B.n374 585
R277 B.n373 B.n372 585
R278 B.n371 B.n370 585
R279 B.n369 B.n368 585
R280 B.n367 B.n366 585
R281 B.n320 B.n319 585
R282 B.n529 B.n528 585
R283 B.n528 B.n527 585
R284 B.n316 B.n315 585
R285 B.n317 B.n316 585
R286 B.n535 B.n534 585
R287 B.n534 B.n533 585
R288 B.n536 B.n314 585
R289 B.n314 B.n313 585
R290 B.n538 B.n537 585
R291 B.n539 B.n538 585
R292 B.n308 B.n307 585
R293 B.n309 B.n308 585
R294 B.n547 B.n546 585
R295 B.n546 B.n545 585
R296 B.n548 B.n306 585
R297 B.n306 B.n304 585
R298 B.n550 B.n549 585
R299 B.n551 B.n550 585
R300 B.n300 B.n299 585
R301 B.n305 B.n300 585
R302 B.n559 B.n558 585
R303 B.n558 B.n557 585
R304 B.n560 B.n298 585
R305 B.n298 B.n297 585
R306 B.n562 B.n561 585
R307 B.n563 B.n562 585
R308 B.n292 B.n291 585
R309 B.n293 B.n292 585
R310 B.n571 B.n570 585
R311 B.n570 B.n569 585
R312 B.n572 B.n290 585
R313 B.n290 B.n289 585
R314 B.n574 B.n573 585
R315 B.n575 B.n574 585
R316 B.n284 B.n283 585
R317 B.n285 B.n284 585
R318 B.n583 B.n582 585
R319 B.n582 B.n581 585
R320 B.n584 B.n282 585
R321 B.n282 B.n281 585
R322 B.n586 B.n585 585
R323 B.n587 B.n586 585
R324 B.n276 B.n275 585
R325 B.n277 B.n276 585
R326 B.n596 B.n595 585
R327 B.n595 B.n594 585
R328 B.n597 B.n274 585
R329 B.n593 B.n274 585
R330 B.n599 B.n598 585
R331 B.n600 B.n599 585
R332 B.n269 B.n268 585
R333 B.n270 B.n269 585
R334 B.n609 B.n608 585
R335 B.n608 B.n607 585
R336 B.n610 B.n267 585
R337 B.n267 B.n266 585
R338 B.n612 B.n611 585
R339 B.n613 B.n612 585
R340 B.n2 B.n0 585
R341 B.n4 B.n2 585
R342 B.n3 B.n1 585
R343 B.n714 B.n3 585
R344 B.n712 B.n711 585
R345 B.n713 B.n712 585
R346 B.n710 B.n9 585
R347 B.n9 B.n8 585
R348 B.n709 B.n708 585
R349 B.n708 B.n707 585
R350 B.n11 B.n10 585
R351 B.n706 B.n11 585
R352 B.n704 B.n703 585
R353 B.n705 B.n704 585
R354 B.n702 B.n15 585
R355 B.n18 B.n15 585
R356 B.n701 B.n700 585
R357 B.n700 B.n699 585
R358 B.n17 B.n16 585
R359 B.n698 B.n17 585
R360 B.n696 B.n695 585
R361 B.n697 B.n696 585
R362 B.n694 B.n23 585
R363 B.n23 B.n22 585
R364 B.n693 B.n692 585
R365 B.n692 B.n691 585
R366 B.n25 B.n24 585
R367 B.n690 B.n25 585
R368 B.n688 B.n687 585
R369 B.n689 B.n688 585
R370 B.n686 B.n30 585
R371 B.n30 B.n29 585
R372 B.n685 B.n684 585
R373 B.n684 B.n683 585
R374 B.n32 B.n31 585
R375 B.n682 B.n32 585
R376 B.n680 B.n679 585
R377 B.n681 B.n680 585
R378 B.n678 B.n37 585
R379 B.n37 B.n36 585
R380 B.n677 B.n676 585
R381 B.n676 B.n675 585
R382 B.n39 B.n38 585
R383 B.n674 B.n39 585
R384 B.n672 B.n671 585
R385 B.n673 B.n672 585
R386 B.n670 B.n44 585
R387 B.n44 B.n43 585
R388 B.n669 B.n668 585
R389 B.n668 B.n667 585
R390 B.n46 B.n45 585
R391 B.n666 B.n46 585
R392 B.n664 B.n663 585
R393 B.n665 B.n664 585
R394 B.n662 B.n51 585
R395 B.n51 B.n50 585
R396 B.n661 B.n660 585
R397 B.n660 B.n659 585
R398 B.n53 B.n52 585
R399 B.n658 B.n53 585
R400 B.n717 B.n716 585
R401 B.n716 B.n715 585
R402 B.n525 B.n316 482.89
R403 B.n103 B.n53 482.89
R404 B.n528 B.n318 482.89
R405 B.n655 B.n55 482.89
R406 B.n364 B.t15 318.822
R407 B.n97 B.t4 318.822
R408 B.n362 B.t12 318.822
R409 B.n100 B.t7 318.822
R410 B.n364 B.t13 284.267
R411 B.n362 B.t9 284.267
R412 B.n100 B.t6 284.267
R413 B.n97 B.t2 284.267
R414 B.n657 B.n656 256.663
R415 B.n657 B.n95 256.663
R416 B.n657 B.n94 256.663
R417 B.n657 B.n93 256.663
R418 B.n657 B.n92 256.663
R419 B.n657 B.n91 256.663
R420 B.n657 B.n90 256.663
R421 B.n657 B.n89 256.663
R422 B.n657 B.n88 256.663
R423 B.n657 B.n87 256.663
R424 B.n657 B.n86 256.663
R425 B.n657 B.n85 256.663
R426 B.n657 B.n84 256.663
R427 B.n657 B.n83 256.663
R428 B.n657 B.n82 256.663
R429 B.n657 B.n81 256.663
R430 B.n657 B.n80 256.663
R431 B.n657 B.n79 256.663
R432 B.n657 B.n78 256.663
R433 B.n657 B.n77 256.663
R434 B.n657 B.n76 256.663
R435 B.n657 B.n75 256.663
R436 B.n657 B.n74 256.663
R437 B.n657 B.n73 256.663
R438 B.n657 B.n72 256.663
R439 B.n657 B.n71 256.663
R440 B.n657 B.n70 256.663
R441 B.n657 B.n69 256.663
R442 B.n657 B.n68 256.663
R443 B.n657 B.n67 256.663
R444 B.n657 B.n66 256.663
R445 B.n657 B.n65 256.663
R446 B.n657 B.n64 256.663
R447 B.n657 B.n63 256.663
R448 B.n657 B.n62 256.663
R449 B.n657 B.n61 256.663
R450 B.n657 B.n60 256.663
R451 B.n657 B.n59 256.663
R452 B.n657 B.n58 256.663
R453 B.n657 B.n57 256.663
R454 B.n657 B.n56 256.663
R455 B.n527 B.n526 256.663
R456 B.n527 B.n321 256.663
R457 B.n527 B.n322 256.663
R458 B.n527 B.n323 256.663
R459 B.n527 B.n324 256.663
R460 B.n527 B.n325 256.663
R461 B.n527 B.n326 256.663
R462 B.n527 B.n327 256.663
R463 B.n527 B.n328 256.663
R464 B.n527 B.n329 256.663
R465 B.n527 B.n330 256.663
R466 B.n527 B.n331 256.663
R467 B.n527 B.n332 256.663
R468 B.n527 B.n333 256.663
R469 B.n527 B.n334 256.663
R470 B.n527 B.n335 256.663
R471 B.n527 B.n336 256.663
R472 B.n527 B.n337 256.663
R473 B.n527 B.n338 256.663
R474 B.n527 B.n339 256.663
R475 B.n527 B.n340 256.663
R476 B.n527 B.n341 256.663
R477 B.n527 B.n342 256.663
R478 B.n527 B.n343 256.663
R479 B.n527 B.n344 256.663
R480 B.n527 B.n345 256.663
R481 B.n527 B.n346 256.663
R482 B.n527 B.n347 256.663
R483 B.n527 B.n348 256.663
R484 B.n527 B.n349 256.663
R485 B.n527 B.n350 256.663
R486 B.n527 B.n351 256.663
R487 B.n527 B.n352 256.663
R488 B.n527 B.n353 256.663
R489 B.n527 B.n354 256.663
R490 B.n527 B.n355 256.663
R491 B.n527 B.n356 256.663
R492 B.n527 B.n357 256.663
R493 B.n527 B.n358 256.663
R494 B.n527 B.n359 256.663
R495 B.n365 B.t14 249.78
R496 B.n98 B.t5 249.78
R497 B.n363 B.t11 249.78
R498 B.n101 B.t8 249.78
R499 B.n534 B.n316 163.367
R500 B.n534 B.n314 163.367
R501 B.n538 B.n314 163.367
R502 B.n538 B.n308 163.367
R503 B.n546 B.n308 163.367
R504 B.n546 B.n306 163.367
R505 B.n550 B.n306 163.367
R506 B.n550 B.n300 163.367
R507 B.n558 B.n300 163.367
R508 B.n558 B.n298 163.367
R509 B.n562 B.n298 163.367
R510 B.n562 B.n292 163.367
R511 B.n570 B.n292 163.367
R512 B.n570 B.n290 163.367
R513 B.n574 B.n290 163.367
R514 B.n574 B.n284 163.367
R515 B.n582 B.n284 163.367
R516 B.n582 B.n282 163.367
R517 B.n586 B.n282 163.367
R518 B.n586 B.n276 163.367
R519 B.n595 B.n276 163.367
R520 B.n595 B.n274 163.367
R521 B.n599 B.n274 163.367
R522 B.n599 B.n269 163.367
R523 B.n608 B.n269 163.367
R524 B.n608 B.n267 163.367
R525 B.n612 B.n267 163.367
R526 B.n612 B.n2 163.367
R527 B.n716 B.n2 163.367
R528 B.n716 B.n3 163.367
R529 B.n712 B.n3 163.367
R530 B.n712 B.n9 163.367
R531 B.n708 B.n9 163.367
R532 B.n708 B.n11 163.367
R533 B.n704 B.n11 163.367
R534 B.n704 B.n15 163.367
R535 B.n700 B.n15 163.367
R536 B.n700 B.n17 163.367
R537 B.n696 B.n17 163.367
R538 B.n696 B.n23 163.367
R539 B.n692 B.n23 163.367
R540 B.n692 B.n25 163.367
R541 B.n688 B.n25 163.367
R542 B.n688 B.n30 163.367
R543 B.n684 B.n30 163.367
R544 B.n684 B.n32 163.367
R545 B.n680 B.n32 163.367
R546 B.n680 B.n37 163.367
R547 B.n676 B.n37 163.367
R548 B.n676 B.n39 163.367
R549 B.n672 B.n39 163.367
R550 B.n672 B.n44 163.367
R551 B.n668 B.n44 163.367
R552 B.n668 B.n46 163.367
R553 B.n664 B.n46 163.367
R554 B.n664 B.n51 163.367
R555 B.n660 B.n51 163.367
R556 B.n660 B.n53 163.367
R557 B.n361 B.n360 163.367
R558 B.n520 B.n360 163.367
R559 B.n518 B.n517 163.367
R560 B.n514 B.n513 163.367
R561 B.n510 B.n509 163.367
R562 B.n506 B.n505 163.367
R563 B.n502 B.n501 163.367
R564 B.n498 B.n497 163.367
R565 B.n494 B.n493 163.367
R566 B.n490 B.n489 163.367
R567 B.n486 B.n485 163.367
R568 B.n482 B.n481 163.367
R569 B.n478 B.n477 163.367
R570 B.n474 B.n473 163.367
R571 B.n470 B.n469 163.367
R572 B.n466 B.n465 163.367
R573 B.n462 B.n461 163.367
R574 B.n458 B.n457 163.367
R575 B.n453 B.n452 163.367
R576 B.n449 B.n448 163.367
R577 B.n445 B.n444 163.367
R578 B.n441 B.n440 163.367
R579 B.n437 B.n436 163.367
R580 B.n432 B.n431 163.367
R581 B.n428 B.n427 163.367
R582 B.n424 B.n423 163.367
R583 B.n420 B.n419 163.367
R584 B.n416 B.n415 163.367
R585 B.n412 B.n411 163.367
R586 B.n408 B.n407 163.367
R587 B.n404 B.n403 163.367
R588 B.n400 B.n399 163.367
R589 B.n396 B.n395 163.367
R590 B.n392 B.n391 163.367
R591 B.n388 B.n387 163.367
R592 B.n384 B.n383 163.367
R593 B.n380 B.n379 163.367
R594 B.n376 B.n375 163.367
R595 B.n372 B.n371 163.367
R596 B.n368 B.n367 163.367
R597 B.n528 B.n320 163.367
R598 B.n532 B.n318 163.367
R599 B.n532 B.n312 163.367
R600 B.n540 B.n312 163.367
R601 B.n540 B.n310 163.367
R602 B.n544 B.n310 163.367
R603 B.n544 B.n303 163.367
R604 B.n552 B.n303 163.367
R605 B.n552 B.n301 163.367
R606 B.n556 B.n301 163.367
R607 B.n556 B.n296 163.367
R608 B.n564 B.n296 163.367
R609 B.n564 B.n294 163.367
R610 B.n568 B.n294 163.367
R611 B.n568 B.n288 163.367
R612 B.n576 B.n288 163.367
R613 B.n576 B.n286 163.367
R614 B.n580 B.n286 163.367
R615 B.n580 B.n280 163.367
R616 B.n588 B.n280 163.367
R617 B.n588 B.n278 163.367
R618 B.n592 B.n278 163.367
R619 B.n592 B.n273 163.367
R620 B.n601 B.n273 163.367
R621 B.n601 B.n271 163.367
R622 B.n606 B.n271 163.367
R623 B.n606 B.n265 163.367
R624 B.n614 B.n265 163.367
R625 B.n615 B.n614 163.367
R626 B.n615 B.n5 163.367
R627 B.n6 B.n5 163.367
R628 B.n7 B.n6 163.367
R629 B.n620 B.n7 163.367
R630 B.n620 B.n12 163.367
R631 B.n13 B.n12 163.367
R632 B.n14 B.n13 163.367
R633 B.n625 B.n14 163.367
R634 B.n625 B.n19 163.367
R635 B.n20 B.n19 163.367
R636 B.n21 B.n20 163.367
R637 B.n630 B.n21 163.367
R638 B.n630 B.n26 163.367
R639 B.n27 B.n26 163.367
R640 B.n28 B.n27 163.367
R641 B.n635 B.n28 163.367
R642 B.n635 B.n33 163.367
R643 B.n34 B.n33 163.367
R644 B.n35 B.n34 163.367
R645 B.n640 B.n35 163.367
R646 B.n640 B.n40 163.367
R647 B.n41 B.n40 163.367
R648 B.n42 B.n41 163.367
R649 B.n645 B.n42 163.367
R650 B.n645 B.n47 163.367
R651 B.n48 B.n47 163.367
R652 B.n49 B.n48 163.367
R653 B.n650 B.n49 163.367
R654 B.n650 B.n54 163.367
R655 B.n55 B.n54 163.367
R656 B.n107 B.n106 163.367
R657 B.n111 B.n110 163.367
R658 B.n115 B.n114 163.367
R659 B.n119 B.n118 163.367
R660 B.n123 B.n122 163.367
R661 B.n127 B.n126 163.367
R662 B.n131 B.n130 163.367
R663 B.n135 B.n134 163.367
R664 B.n139 B.n138 163.367
R665 B.n143 B.n142 163.367
R666 B.n147 B.n146 163.367
R667 B.n151 B.n150 163.367
R668 B.n155 B.n154 163.367
R669 B.n159 B.n158 163.367
R670 B.n163 B.n162 163.367
R671 B.n167 B.n166 163.367
R672 B.n171 B.n170 163.367
R673 B.n175 B.n174 163.367
R674 B.n179 B.n178 163.367
R675 B.n183 B.n182 163.367
R676 B.n187 B.n186 163.367
R677 B.n191 B.n190 163.367
R678 B.n195 B.n194 163.367
R679 B.n199 B.n198 163.367
R680 B.n203 B.n202 163.367
R681 B.n207 B.n206 163.367
R682 B.n211 B.n210 163.367
R683 B.n215 B.n214 163.367
R684 B.n219 B.n218 163.367
R685 B.n223 B.n222 163.367
R686 B.n227 B.n226 163.367
R687 B.n231 B.n230 163.367
R688 B.n235 B.n234 163.367
R689 B.n239 B.n238 163.367
R690 B.n243 B.n242 163.367
R691 B.n247 B.n246 163.367
R692 B.n251 B.n250 163.367
R693 B.n255 B.n254 163.367
R694 B.n259 B.n258 163.367
R695 B.n261 B.n96 163.367
R696 B.n527 B.n317 90.8032
R697 B.n658 B.n657 90.8032
R698 B.n526 B.n525 71.676
R699 B.n520 B.n321 71.676
R700 B.n517 B.n322 71.676
R701 B.n513 B.n323 71.676
R702 B.n509 B.n324 71.676
R703 B.n505 B.n325 71.676
R704 B.n501 B.n326 71.676
R705 B.n497 B.n327 71.676
R706 B.n493 B.n328 71.676
R707 B.n489 B.n329 71.676
R708 B.n485 B.n330 71.676
R709 B.n481 B.n331 71.676
R710 B.n477 B.n332 71.676
R711 B.n473 B.n333 71.676
R712 B.n469 B.n334 71.676
R713 B.n465 B.n335 71.676
R714 B.n461 B.n336 71.676
R715 B.n457 B.n337 71.676
R716 B.n452 B.n338 71.676
R717 B.n448 B.n339 71.676
R718 B.n444 B.n340 71.676
R719 B.n440 B.n341 71.676
R720 B.n436 B.n342 71.676
R721 B.n431 B.n343 71.676
R722 B.n427 B.n344 71.676
R723 B.n423 B.n345 71.676
R724 B.n419 B.n346 71.676
R725 B.n415 B.n347 71.676
R726 B.n411 B.n348 71.676
R727 B.n407 B.n349 71.676
R728 B.n403 B.n350 71.676
R729 B.n399 B.n351 71.676
R730 B.n395 B.n352 71.676
R731 B.n391 B.n353 71.676
R732 B.n387 B.n354 71.676
R733 B.n383 B.n355 71.676
R734 B.n379 B.n356 71.676
R735 B.n375 B.n357 71.676
R736 B.n371 B.n358 71.676
R737 B.n367 B.n359 71.676
R738 B.n103 B.n56 71.676
R739 B.n107 B.n57 71.676
R740 B.n111 B.n58 71.676
R741 B.n115 B.n59 71.676
R742 B.n119 B.n60 71.676
R743 B.n123 B.n61 71.676
R744 B.n127 B.n62 71.676
R745 B.n131 B.n63 71.676
R746 B.n135 B.n64 71.676
R747 B.n139 B.n65 71.676
R748 B.n143 B.n66 71.676
R749 B.n147 B.n67 71.676
R750 B.n151 B.n68 71.676
R751 B.n155 B.n69 71.676
R752 B.n159 B.n70 71.676
R753 B.n163 B.n71 71.676
R754 B.n167 B.n72 71.676
R755 B.n171 B.n73 71.676
R756 B.n175 B.n74 71.676
R757 B.n179 B.n75 71.676
R758 B.n183 B.n76 71.676
R759 B.n187 B.n77 71.676
R760 B.n191 B.n78 71.676
R761 B.n195 B.n79 71.676
R762 B.n199 B.n80 71.676
R763 B.n203 B.n81 71.676
R764 B.n207 B.n82 71.676
R765 B.n211 B.n83 71.676
R766 B.n215 B.n84 71.676
R767 B.n219 B.n85 71.676
R768 B.n223 B.n86 71.676
R769 B.n227 B.n87 71.676
R770 B.n231 B.n88 71.676
R771 B.n235 B.n89 71.676
R772 B.n239 B.n90 71.676
R773 B.n243 B.n91 71.676
R774 B.n247 B.n92 71.676
R775 B.n251 B.n93 71.676
R776 B.n255 B.n94 71.676
R777 B.n259 B.n95 71.676
R778 B.n656 B.n96 71.676
R779 B.n656 B.n655 71.676
R780 B.n261 B.n95 71.676
R781 B.n258 B.n94 71.676
R782 B.n254 B.n93 71.676
R783 B.n250 B.n92 71.676
R784 B.n246 B.n91 71.676
R785 B.n242 B.n90 71.676
R786 B.n238 B.n89 71.676
R787 B.n234 B.n88 71.676
R788 B.n230 B.n87 71.676
R789 B.n226 B.n86 71.676
R790 B.n222 B.n85 71.676
R791 B.n218 B.n84 71.676
R792 B.n214 B.n83 71.676
R793 B.n210 B.n82 71.676
R794 B.n206 B.n81 71.676
R795 B.n202 B.n80 71.676
R796 B.n198 B.n79 71.676
R797 B.n194 B.n78 71.676
R798 B.n190 B.n77 71.676
R799 B.n186 B.n76 71.676
R800 B.n182 B.n75 71.676
R801 B.n178 B.n74 71.676
R802 B.n174 B.n73 71.676
R803 B.n170 B.n72 71.676
R804 B.n166 B.n71 71.676
R805 B.n162 B.n70 71.676
R806 B.n158 B.n69 71.676
R807 B.n154 B.n68 71.676
R808 B.n150 B.n67 71.676
R809 B.n146 B.n66 71.676
R810 B.n142 B.n65 71.676
R811 B.n138 B.n64 71.676
R812 B.n134 B.n63 71.676
R813 B.n130 B.n62 71.676
R814 B.n126 B.n61 71.676
R815 B.n122 B.n60 71.676
R816 B.n118 B.n59 71.676
R817 B.n114 B.n58 71.676
R818 B.n110 B.n57 71.676
R819 B.n106 B.n56 71.676
R820 B.n526 B.n361 71.676
R821 B.n518 B.n321 71.676
R822 B.n514 B.n322 71.676
R823 B.n510 B.n323 71.676
R824 B.n506 B.n324 71.676
R825 B.n502 B.n325 71.676
R826 B.n498 B.n326 71.676
R827 B.n494 B.n327 71.676
R828 B.n490 B.n328 71.676
R829 B.n486 B.n329 71.676
R830 B.n482 B.n330 71.676
R831 B.n478 B.n331 71.676
R832 B.n474 B.n332 71.676
R833 B.n470 B.n333 71.676
R834 B.n466 B.n334 71.676
R835 B.n462 B.n335 71.676
R836 B.n458 B.n336 71.676
R837 B.n453 B.n337 71.676
R838 B.n449 B.n338 71.676
R839 B.n445 B.n339 71.676
R840 B.n441 B.n340 71.676
R841 B.n437 B.n341 71.676
R842 B.n432 B.n342 71.676
R843 B.n428 B.n343 71.676
R844 B.n424 B.n344 71.676
R845 B.n420 B.n345 71.676
R846 B.n416 B.n346 71.676
R847 B.n412 B.n347 71.676
R848 B.n408 B.n348 71.676
R849 B.n404 B.n349 71.676
R850 B.n400 B.n350 71.676
R851 B.n396 B.n351 71.676
R852 B.n392 B.n352 71.676
R853 B.n388 B.n353 71.676
R854 B.n384 B.n354 71.676
R855 B.n380 B.n355 71.676
R856 B.n376 B.n356 71.676
R857 B.n372 B.n357 71.676
R858 B.n368 B.n358 71.676
R859 B.n359 B.n320 71.676
R860 B.n365 B.n364 69.0429
R861 B.n363 B.n362 69.0429
R862 B.n101 B.n100 69.0429
R863 B.n98 B.n97 69.0429
R864 B.n434 B.n365 59.5399
R865 B.n455 B.n363 59.5399
R866 B.n102 B.n101 59.5399
R867 B.n99 B.n98 59.5399
R868 B.n533 B.n317 48.6193
R869 B.n533 B.n313 48.6193
R870 B.n539 B.n313 48.6193
R871 B.n539 B.n309 48.6193
R872 B.n545 B.n309 48.6193
R873 B.n545 B.n304 48.6193
R874 B.n551 B.n304 48.6193
R875 B.n551 B.n305 48.6193
R876 B.n557 B.n297 48.6193
R877 B.n563 B.n297 48.6193
R878 B.n563 B.n293 48.6193
R879 B.n569 B.n293 48.6193
R880 B.n569 B.n289 48.6193
R881 B.n575 B.n289 48.6193
R882 B.n575 B.n285 48.6193
R883 B.n581 B.n285 48.6193
R884 B.n581 B.n281 48.6193
R885 B.n587 B.n281 48.6193
R886 B.n587 B.n277 48.6193
R887 B.n594 B.n277 48.6193
R888 B.n594 B.n593 48.6193
R889 B.n600 B.n270 48.6193
R890 B.n607 B.n270 48.6193
R891 B.n607 B.n266 48.6193
R892 B.n613 B.n266 48.6193
R893 B.n613 B.n4 48.6193
R894 B.n715 B.n4 48.6193
R895 B.n715 B.n714 48.6193
R896 B.n714 B.n713 48.6193
R897 B.n713 B.n8 48.6193
R898 B.n707 B.n8 48.6193
R899 B.n707 B.n706 48.6193
R900 B.n706 B.n705 48.6193
R901 B.n699 B.n18 48.6193
R902 B.n699 B.n698 48.6193
R903 B.n698 B.n697 48.6193
R904 B.n697 B.n22 48.6193
R905 B.n691 B.n22 48.6193
R906 B.n691 B.n690 48.6193
R907 B.n690 B.n689 48.6193
R908 B.n689 B.n29 48.6193
R909 B.n683 B.n29 48.6193
R910 B.n683 B.n682 48.6193
R911 B.n682 B.n681 48.6193
R912 B.n681 B.n36 48.6193
R913 B.n675 B.n36 48.6193
R914 B.n674 B.n673 48.6193
R915 B.n673 B.n43 48.6193
R916 B.n667 B.n43 48.6193
R917 B.n667 B.n666 48.6193
R918 B.n666 B.n665 48.6193
R919 B.n665 B.n50 48.6193
R920 B.n659 B.n50 48.6193
R921 B.n659 B.n658 48.6193
R922 B.n600 B.t0 40.7545
R923 B.n705 B.t1 40.7545
R924 B.n104 B.n52 31.3761
R925 B.n654 B.n653 31.3761
R926 B.n530 B.n529 31.3761
R927 B.n524 B.n315 31.3761
R928 B.n557 B.t10 25.0249
R929 B.n675 B.t3 25.0249
R930 B.n305 B.t10 23.5949
R931 B.t3 B.n674 23.5949
R932 B B.n717 18.0485
R933 B.n105 B.n104 10.6151
R934 B.n108 B.n105 10.6151
R935 B.n109 B.n108 10.6151
R936 B.n112 B.n109 10.6151
R937 B.n113 B.n112 10.6151
R938 B.n116 B.n113 10.6151
R939 B.n117 B.n116 10.6151
R940 B.n120 B.n117 10.6151
R941 B.n121 B.n120 10.6151
R942 B.n124 B.n121 10.6151
R943 B.n125 B.n124 10.6151
R944 B.n128 B.n125 10.6151
R945 B.n129 B.n128 10.6151
R946 B.n132 B.n129 10.6151
R947 B.n133 B.n132 10.6151
R948 B.n136 B.n133 10.6151
R949 B.n137 B.n136 10.6151
R950 B.n140 B.n137 10.6151
R951 B.n141 B.n140 10.6151
R952 B.n144 B.n141 10.6151
R953 B.n145 B.n144 10.6151
R954 B.n148 B.n145 10.6151
R955 B.n149 B.n148 10.6151
R956 B.n152 B.n149 10.6151
R957 B.n153 B.n152 10.6151
R958 B.n156 B.n153 10.6151
R959 B.n157 B.n156 10.6151
R960 B.n160 B.n157 10.6151
R961 B.n161 B.n160 10.6151
R962 B.n164 B.n161 10.6151
R963 B.n165 B.n164 10.6151
R964 B.n168 B.n165 10.6151
R965 B.n169 B.n168 10.6151
R966 B.n172 B.n169 10.6151
R967 B.n173 B.n172 10.6151
R968 B.n177 B.n176 10.6151
R969 B.n180 B.n177 10.6151
R970 B.n181 B.n180 10.6151
R971 B.n184 B.n181 10.6151
R972 B.n185 B.n184 10.6151
R973 B.n188 B.n185 10.6151
R974 B.n189 B.n188 10.6151
R975 B.n192 B.n189 10.6151
R976 B.n193 B.n192 10.6151
R977 B.n197 B.n196 10.6151
R978 B.n200 B.n197 10.6151
R979 B.n201 B.n200 10.6151
R980 B.n204 B.n201 10.6151
R981 B.n205 B.n204 10.6151
R982 B.n208 B.n205 10.6151
R983 B.n209 B.n208 10.6151
R984 B.n212 B.n209 10.6151
R985 B.n213 B.n212 10.6151
R986 B.n216 B.n213 10.6151
R987 B.n217 B.n216 10.6151
R988 B.n220 B.n217 10.6151
R989 B.n221 B.n220 10.6151
R990 B.n224 B.n221 10.6151
R991 B.n225 B.n224 10.6151
R992 B.n228 B.n225 10.6151
R993 B.n229 B.n228 10.6151
R994 B.n232 B.n229 10.6151
R995 B.n233 B.n232 10.6151
R996 B.n236 B.n233 10.6151
R997 B.n237 B.n236 10.6151
R998 B.n240 B.n237 10.6151
R999 B.n241 B.n240 10.6151
R1000 B.n244 B.n241 10.6151
R1001 B.n245 B.n244 10.6151
R1002 B.n248 B.n245 10.6151
R1003 B.n249 B.n248 10.6151
R1004 B.n252 B.n249 10.6151
R1005 B.n253 B.n252 10.6151
R1006 B.n256 B.n253 10.6151
R1007 B.n257 B.n256 10.6151
R1008 B.n260 B.n257 10.6151
R1009 B.n262 B.n260 10.6151
R1010 B.n263 B.n262 10.6151
R1011 B.n654 B.n263 10.6151
R1012 B.n531 B.n530 10.6151
R1013 B.n531 B.n311 10.6151
R1014 B.n541 B.n311 10.6151
R1015 B.n542 B.n541 10.6151
R1016 B.n543 B.n542 10.6151
R1017 B.n543 B.n302 10.6151
R1018 B.n553 B.n302 10.6151
R1019 B.n554 B.n553 10.6151
R1020 B.n555 B.n554 10.6151
R1021 B.n555 B.n295 10.6151
R1022 B.n565 B.n295 10.6151
R1023 B.n566 B.n565 10.6151
R1024 B.n567 B.n566 10.6151
R1025 B.n567 B.n287 10.6151
R1026 B.n577 B.n287 10.6151
R1027 B.n578 B.n577 10.6151
R1028 B.n579 B.n578 10.6151
R1029 B.n579 B.n279 10.6151
R1030 B.n589 B.n279 10.6151
R1031 B.n590 B.n589 10.6151
R1032 B.n591 B.n590 10.6151
R1033 B.n591 B.n272 10.6151
R1034 B.n602 B.n272 10.6151
R1035 B.n603 B.n602 10.6151
R1036 B.n605 B.n603 10.6151
R1037 B.n605 B.n604 10.6151
R1038 B.n604 B.n264 10.6151
R1039 B.n616 B.n264 10.6151
R1040 B.n617 B.n616 10.6151
R1041 B.n618 B.n617 10.6151
R1042 B.n619 B.n618 10.6151
R1043 B.n621 B.n619 10.6151
R1044 B.n622 B.n621 10.6151
R1045 B.n623 B.n622 10.6151
R1046 B.n624 B.n623 10.6151
R1047 B.n626 B.n624 10.6151
R1048 B.n627 B.n626 10.6151
R1049 B.n628 B.n627 10.6151
R1050 B.n629 B.n628 10.6151
R1051 B.n631 B.n629 10.6151
R1052 B.n632 B.n631 10.6151
R1053 B.n633 B.n632 10.6151
R1054 B.n634 B.n633 10.6151
R1055 B.n636 B.n634 10.6151
R1056 B.n637 B.n636 10.6151
R1057 B.n638 B.n637 10.6151
R1058 B.n639 B.n638 10.6151
R1059 B.n641 B.n639 10.6151
R1060 B.n642 B.n641 10.6151
R1061 B.n643 B.n642 10.6151
R1062 B.n644 B.n643 10.6151
R1063 B.n646 B.n644 10.6151
R1064 B.n647 B.n646 10.6151
R1065 B.n648 B.n647 10.6151
R1066 B.n649 B.n648 10.6151
R1067 B.n651 B.n649 10.6151
R1068 B.n652 B.n651 10.6151
R1069 B.n653 B.n652 10.6151
R1070 B.n524 B.n523 10.6151
R1071 B.n523 B.n522 10.6151
R1072 B.n522 B.n521 10.6151
R1073 B.n521 B.n519 10.6151
R1074 B.n519 B.n516 10.6151
R1075 B.n516 B.n515 10.6151
R1076 B.n515 B.n512 10.6151
R1077 B.n512 B.n511 10.6151
R1078 B.n511 B.n508 10.6151
R1079 B.n508 B.n507 10.6151
R1080 B.n507 B.n504 10.6151
R1081 B.n504 B.n503 10.6151
R1082 B.n503 B.n500 10.6151
R1083 B.n500 B.n499 10.6151
R1084 B.n499 B.n496 10.6151
R1085 B.n496 B.n495 10.6151
R1086 B.n495 B.n492 10.6151
R1087 B.n492 B.n491 10.6151
R1088 B.n491 B.n488 10.6151
R1089 B.n488 B.n487 10.6151
R1090 B.n487 B.n484 10.6151
R1091 B.n484 B.n483 10.6151
R1092 B.n483 B.n480 10.6151
R1093 B.n480 B.n479 10.6151
R1094 B.n479 B.n476 10.6151
R1095 B.n476 B.n475 10.6151
R1096 B.n475 B.n472 10.6151
R1097 B.n472 B.n471 10.6151
R1098 B.n471 B.n468 10.6151
R1099 B.n468 B.n467 10.6151
R1100 B.n467 B.n464 10.6151
R1101 B.n464 B.n463 10.6151
R1102 B.n463 B.n460 10.6151
R1103 B.n460 B.n459 10.6151
R1104 B.n459 B.n456 10.6151
R1105 B.n454 B.n451 10.6151
R1106 B.n451 B.n450 10.6151
R1107 B.n450 B.n447 10.6151
R1108 B.n447 B.n446 10.6151
R1109 B.n446 B.n443 10.6151
R1110 B.n443 B.n442 10.6151
R1111 B.n442 B.n439 10.6151
R1112 B.n439 B.n438 10.6151
R1113 B.n438 B.n435 10.6151
R1114 B.n433 B.n430 10.6151
R1115 B.n430 B.n429 10.6151
R1116 B.n429 B.n426 10.6151
R1117 B.n426 B.n425 10.6151
R1118 B.n425 B.n422 10.6151
R1119 B.n422 B.n421 10.6151
R1120 B.n421 B.n418 10.6151
R1121 B.n418 B.n417 10.6151
R1122 B.n417 B.n414 10.6151
R1123 B.n414 B.n413 10.6151
R1124 B.n413 B.n410 10.6151
R1125 B.n410 B.n409 10.6151
R1126 B.n409 B.n406 10.6151
R1127 B.n406 B.n405 10.6151
R1128 B.n405 B.n402 10.6151
R1129 B.n402 B.n401 10.6151
R1130 B.n401 B.n398 10.6151
R1131 B.n398 B.n397 10.6151
R1132 B.n397 B.n394 10.6151
R1133 B.n394 B.n393 10.6151
R1134 B.n393 B.n390 10.6151
R1135 B.n390 B.n389 10.6151
R1136 B.n389 B.n386 10.6151
R1137 B.n386 B.n385 10.6151
R1138 B.n385 B.n382 10.6151
R1139 B.n382 B.n381 10.6151
R1140 B.n381 B.n378 10.6151
R1141 B.n378 B.n377 10.6151
R1142 B.n377 B.n374 10.6151
R1143 B.n374 B.n373 10.6151
R1144 B.n373 B.n370 10.6151
R1145 B.n370 B.n369 10.6151
R1146 B.n369 B.n366 10.6151
R1147 B.n366 B.n319 10.6151
R1148 B.n529 B.n319 10.6151
R1149 B.n535 B.n315 10.6151
R1150 B.n536 B.n535 10.6151
R1151 B.n537 B.n536 10.6151
R1152 B.n537 B.n307 10.6151
R1153 B.n547 B.n307 10.6151
R1154 B.n548 B.n547 10.6151
R1155 B.n549 B.n548 10.6151
R1156 B.n549 B.n299 10.6151
R1157 B.n559 B.n299 10.6151
R1158 B.n560 B.n559 10.6151
R1159 B.n561 B.n560 10.6151
R1160 B.n561 B.n291 10.6151
R1161 B.n571 B.n291 10.6151
R1162 B.n572 B.n571 10.6151
R1163 B.n573 B.n572 10.6151
R1164 B.n573 B.n283 10.6151
R1165 B.n583 B.n283 10.6151
R1166 B.n584 B.n583 10.6151
R1167 B.n585 B.n584 10.6151
R1168 B.n585 B.n275 10.6151
R1169 B.n596 B.n275 10.6151
R1170 B.n597 B.n596 10.6151
R1171 B.n598 B.n597 10.6151
R1172 B.n598 B.n268 10.6151
R1173 B.n609 B.n268 10.6151
R1174 B.n610 B.n609 10.6151
R1175 B.n611 B.n610 10.6151
R1176 B.n611 B.n0 10.6151
R1177 B.n711 B.n1 10.6151
R1178 B.n711 B.n710 10.6151
R1179 B.n710 B.n709 10.6151
R1180 B.n709 B.n10 10.6151
R1181 B.n703 B.n10 10.6151
R1182 B.n703 B.n702 10.6151
R1183 B.n702 B.n701 10.6151
R1184 B.n701 B.n16 10.6151
R1185 B.n695 B.n16 10.6151
R1186 B.n695 B.n694 10.6151
R1187 B.n694 B.n693 10.6151
R1188 B.n693 B.n24 10.6151
R1189 B.n687 B.n24 10.6151
R1190 B.n687 B.n686 10.6151
R1191 B.n686 B.n685 10.6151
R1192 B.n685 B.n31 10.6151
R1193 B.n679 B.n31 10.6151
R1194 B.n679 B.n678 10.6151
R1195 B.n678 B.n677 10.6151
R1196 B.n677 B.n38 10.6151
R1197 B.n671 B.n38 10.6151
R1198 B.n671 B.n670 10.6151
R1199 B.n670 B.n669 10.6151
R1200 B.n669 B.n45 10.6151
R1201 B.n663 B.n45 10.6151
R1202 B.n663 B.n662 10.6151
R1203 B.n662 B.n661 10.6151
R1204 B.n661 B.n52 10.6151
R1205 B.n173 B.n102 9.36635
R1206 B.n196 B.n99 9.36635
R1207 B.n456 B.n455 9.36635
R1208 B.n434 B.n433 9.36635
R1209 B.n593 B.t0 7.8653
R1210 B.n18 B.t1 7.8653
R1211 B.n717 B.n0 2.81026
R1212 B.n717 B.n1 2.81026
R1213 B.n176 B.n102 1.24928
R1214 B.n193 B.n99 1.24928
R1215 B.n455 B.n454 1.24928
R1216 B.n435 B.n434 1.24928
R1217 VN VN.t0 159.024
R1218 VN VN.t1 114.748
R1219 VTAIL.n210 VTAIL.n162 289.615
R1220 VTAIL.n48 VTAIL.n0 289.615
R1221 VTAIL.n156 VTAIL.n108 289.615
R1222 VTAIL.n102 VTAIL.n54 289.615
R1223 VTAIL.n178 VTAIL.n177 185
R1224 VTAIL.n183 VTAIL.n182 185
R1225 VTAIL.n185 VTAIL.n184 185
R1226 VTAIL.n174 VTAIL.n173 185
R1227 VTAIL.n191 VTAIL.n190 185
R1228 VTAIL.n193 VTAIL.n192 185
R1229 VTAIL.n170 VTAIL.n169 185
R1230 VTAIL.n200 VTAIL.n199 185
R1231 VTAIL.n201 VTAIL.n168 185
R1232 VTAIL.n203 VTAIL.n202 185
R1233 VTAIL.n166 VTAIL.n165 185
R1234 VTAIL.n209 VTAIL.n208 185
R1235 VTAIL.n211 VTAIL.n210 185
R1236 VTAIL.n16 VTAIL.n15 185
R1237 VTAIL.n21 VTAIL.n20 185
R1238 VTAIL.n23 VTAIL.n22 185
R1239 VTAIL.n12 VTAIL.n11 185
R1240 VTAIL.n29 VTAIL.n28 185
R1241 VTAIL.n31 VTAIL.n30 185
R1242 VTAIL.n8 VTAIL.n7 185
R1243 VTAIL.n38 VTAIL.n37 185
R1244 VTAIL.n39 VTAIL.n6 185
R1245 VTAIL.n41 VTAIL.n40 185
R1246 VTAIL.n4 VTAIL.n3 185
R1247 VTAIL.n47 VTAIL.n46 185
R1248 VTAIL.n49 VTAIL.n48 185
R1249 VTAIL.n157 VTAIL.n156 185
R1250 VTAIL.n155 VTAIL.n154 185
R1251 VTAIL.n112 VTAIL.n111 185
R1252 VTAIL.n149 VTAIL.n148 185
R1253 VTAIL.n147 VTAIL.n114 185
R1254 VTAIL.n146 VTAIL.n145 185
R1255 VTAIL.n117 VTAIL.n115 185
R1256 VTAIL.n140 VTAIL.n139 185
R1257 VTAIL.n138 VTAIL.n137 185
R1258 VTAIL.n121 VTAIL.n120 185
R1259 VTAIL.n132 VTAIL.n131 185
R1260 VTAIL.n130 VTAIL.n129 185
R1261 VTAIL.n125 VTAIL.n124 185
R1262 VTAIL.n103 VTAIL.n102 185
R1263 VTAIL.n101 VTAIL.n100 185
R1264 VTAIL.n58 VTAIL.n57 185
R1265 VTAIL.n95 VTAIL.n94 185
R1266 VTAIL.n93 VTAIL.n60 185
R1267 VTAIL.n92 VTAIL.n91 185
R1268 VTAIL.n63 VTAIL.n61 185
R1269 VTAIL.n86 VTAIL.n85 185
R1270 VTAIL.n84 VTAIL.n83 185
R1271 VTAIL.n67 VTAIL.n66 185
R1272 VTAIL.n78 VTAIL.n77 185
R1273 VTAIL.n76 VTAIL.n75 185
R1274 VTAIL.n71 VTAIL.n70 185
R1275 VTAIL.n179 VTAIL.t3 149.524
R1276 VTAIL.n17 VTAIL.t0 149.524
R1277 VTAIL.n126 VTAIL.t1 149.524
R1278 VTAIL.n72 VTAIL.t2 149.524
R1279 VTAIL.n183 VTAIL.n177 104.615
R1280 VTAIL.n184 VTAIL.n183 104.615
R1281 VTAIL.n184 VTAIL.n173 104.615
R1282 VTAIL.n191 VTAIL.n173 104.615
R1283 VTAIL.n192 VTAIL.n191 104.615
R1284 VTAIL.n192 VTAIL.n169 104.615
R1285 VTAIL.n200 VTAIL.n169 104.615
R1286 VTAIL.n201 VTAIL.n200 104.615
R1287 VTAIL.n202 VTAIL.n201 104.615
R1288 VTAIL.n202 VTAIL.n165 104.615
R1289 VTAIL.n209 VTAIL.n165 104.615
R1290 VTAIL.n210 VTAIL.n209 104.615
R1291 VTAIL.n21 VTAIL.n15 104.615
R1292 VTAIL.n22 VTAIL.n21 104.615
R1293 VTAIL.n22 VTAIL.n11 104.615
R1294 VTAIL.n29 VTAIL.n11 104.615
R1295 VTAIL.n30 VTAIL.n29 104.615
R1296 VTAIL.n30 VTAIL.n7 104.615
R1297 VTAIL.n38 VTAIL.n7 104.615
R1298 VTAIL.n39 VTAIL.n38 104.615
R1299 VTAIL.n40 VTAIL.n39 104.615
R1300 VTAIL.n40 VTAIL.n3 104.615
R1301 VTAIL.n47 VTAIL.n3 104.615
R1302 VTAIL.n48 VTAIL.n47 104.615
R1303 VTAIL.n156 VTAIL.n155 104.615
R1304 VTAIL.n155 VTAIL.n111 104.615
R1305 VTAIL.n148 VTAIL.n111 104.615
R1306 VTAIL.n148 VTAIL.n147 104.615
R1307 VTAIL.n147 VTAIL.n146 104.615
R1308 VTAIL.n146 VTAIL.n115 104.615
R1309 VTAIL.n139 VTAIL.n115 104.615
R1310 VTAIL.n139 VTAIL.n138 104.615
R1311 VTAIL.n138 VTAIL.n120 104.615
R1312 VTAIL.n131 VTAIL.n120 104.615
R1313 VTAIL.n131 VTAIL.n130 104.615
R1314 VTAIL.n130 VTAIL.n124 104.615
R1315 VTAIL.n102 VTAIL.n101 104.615
R1316 VTAIL.n101 VTAIL.n57 104.615
R1317 VTAIL.n94 VTAIL.n57 104.615
R1318 VTAIL.n94 VTAIL.n93 104.615
R1319 VTAIL.n93 VTAIL.n92 104.615
R1320 VTAIL.n92 VTAIL.n61 104.615
R1321 VTAIL.n85 VTAIL.n61 104.615
R1322 VTAIL.n85 VTAIL.n84 104.615
R1323 VTAIL.n84 VTAIL.n66 104.615
R1324 VTAIL.n77 VTAIL.n66 104.615
R1325 VTAIL.n77 VTAIL.n76 104.615
R1326 VTAIL.n76 VTAIL.n70 104.615
R1327 VTAIL.t3 VTAIL.n177 52.3082
R1328 VTAIL.t0 VTAIL.n15 52.3082
R1329 VTAIL.t1 VTAIL.n124 52.3082
R1330 VTAIL.t2 VTAIL.n70 52.3082
R1331 VTAIL.n215 VTAIL.n214 35.0944
R1332 VTAIL.n53 VTAIL.n52 35.0944
R1333 VTAIL.n161 VTAIL.n160 35.0944
R1334 VTAIL.n107 VTAIL.n106 35.0944
R1335 VTAIL.n107 VTAIL.n53 27.2203
R1336 VTAIL.n215 VTAIL.n161 24.1514
R1337 VTAIL.n203 VTAIL.n168 13.1884
R1338 VTAIL.n41 VTAIL.n6 13.1884
R1339 VTAIL.n149 VTAIL.n114 13.1884
R1340 VTAIL.n95 VTAIL.n60 13.1884
R1341 VTAIL.n199 VTAIL.n198 12.8005
R1342 VTAIL.n204 VTAIL.n166 12.8005
R1343 VTAIL.n37 VTAIL.n36 12.8005
R1344 VTAIL.n42 VTAIL.n4 12.8005
R1345 VTAIL.n150 VTAIL.n112 12.8005
R1346 VTAIL.n145 VTAIL.n116 12.8005
R1347 VTAIL.n96 VTAIL.n58 12.8005
R1348 VTAIL.n91 VTAIL.n62 12.8005
R1349 VTAIL.n197 VTAIL.n170 12.0247
R1350 VTAIL.n208 VTAIL.n207 12.0247
R1351 VTAIL.n35 VTAIL.n8 12.0247
R1352 VTAIL.n46 VTAIL.n45 12.0247
R1353 VTAIL.n154 VTAIL.n153 12.0247
R1354 VTAIL.n144 VTAIL.n117 12.0247
R1355 VTAIL.n100 VTAIL.n99 12.0247
R1356 VTAIL.n90 VTAIL.n63 12.0247
R1357 VTAIL.n194 VTAIL.n193 11.249
R1358 VTAIL.n211 VTAIL.n164 11.249
R1359 VTAIL.n32 VTAIL.n31 11.249
R1360 VTAIL.n49 VTAIL.n2 11.249
R1361 VTAIL.n157 VTAIL.n110 11.249
R1362 VTAIL.n141 VTAIL.n140 11.249
R1363 VTAIL.n103 VTAIL.n56 11.249
R1364 VTAIL.n87 VTAIL.n86 11.249
R1365 VTAIL.n190 VTAIL.n172 10.4732
R1366 VTAIL.n212 VTAIL.n162 10.4732
R1367 VTAIL.n28 VTAIL.n10 10.4732
R1368 VTAIL.n50 VTAIL.n0 10.4732
R1369 VTAIL.n158 VTAIL.n108 10.4732
R1370 VTAIL.n137 VTAIL.n119 10.4732
R1371 VTAIL.n104 VTAIL.n54 10.4732
R1372 VTAIL.n83 VTAIL.n65 10.4732
R1373 VTAIL.n179 VTAIL.n178 10.2747
R1374 VTAIL.n17 VTAIL.n16 10.2747
R1375 VTAIL.n126 VTAIL.n125 10.2747
R1376 VTAIL.n72 VTAIL.n71 10.2747
R1377 VTAIL.n189 VTAIL.n174 9.69747
R1378 VTAIL.n27 VTAIL.n12 9.69747
R1379 VTAIL.n136 VTAIL.n121 9.69747
R1380 VTAIL.n82 VTAIL.n67 9.69747
R1381 VTAIL.n214 VTAIL.n213 9.45567
R1382 VTAIL.n52 VTAIL.n51 9.45567
R1383 VTAIL.n160 VTAIL.n159 9.45567
R1384 VTAIL.n106 VTAIL.n105 9.45567
R1385 VTAIL.n213 VTAIL.n212 9.3005
R1386 VTAIL.n164 VTAIL.n163 9.3005
R1387 VTAIL.n207 VTAIL.n206 9.3005
R1388 VTAIL.n205 VTAIL.n204 9.3005
R1389 VTAIL.n181 VTAIL.n180 9.3005
R1390 VTAIL.n176 VTAIL.n175 9.3005
R1391 VTAIL.n187 VTAIL.n186 9.3005
R1392 VTAIL.n189 VTAIL.n188 9.3005
R1393 VTAIL.n172 VTAIL.n171 9.3005
R1394 VTAIL.n195 VTAIL.n194 9.3005
R1395 VTAIL.n197 VTAIL.n196 9.3005
R1396 VTAIL.n198 VTAIL.n167 9.3005
R1397 VTAIL.n51 VTAIL.n50 9.3005
R1398 VTAIL.n2 VTAIL.n1 9.3005
R1399 VTAIL.n45 VTAIL.n44 9.3005
R1400 VTAIL.n43 VTAIL.n42 9.3005
R1401 VTAIL.n19 VTAIL.n18 9.3005
R1402 VTAIL.n14 VTAIL.n13 9.3005
R1403 VTAIL.n25 VTAIL.n24 9.3005
R1404 VTAIL.n27 VTAIL.n26 9.3005
R1405 VTAIL.n10 VTAIL.n9 9.3005
R1406 VTAIL.n33 VTAIL.n32 9.3005
R1407 VTAIL.n35 VTAIL.n34 9.3005
R1408 VTAIL.n36 VTAIL.n5 9.3005
R1409 VTAIL.n128 VTAIL.n127 9.3005
R1410 VTAIL.n123 VTAIL.n122 9.3005
R1411 VTAIL.n134 VTAIL.n133 9.3005
R1412 VTAIL.n136 VTAIL.n135 9.3005
R1413 VTAIL.n119 VTAIL.n118 9.3005
R1414 VTAIL.n142 VTAIL.n141 9.3005
R1415 VTAIL.n144 VTAIL.n143 9.3005
R1416 VTAIL.n116 VTAIL.n113 9.3005
R1417 VTAIL.n159 VTAIL.n158 9.3005
R1418 VTAIL.n110 VTAIL.n109 9.3005
R1419 VTAIL.n153 VTAIL.n152 9.3005
R1420 VTAIL.n151 VTAIL.n150 9.3005
R1421 VTAIL.n74 VTAIL.n73 9.3005
R1422 VTAIL.n69 VTAIL.n68 9.3005
R1423 VTAIL.n80 VTAIL.n79 9.3005
R1424 VTAIL.n82 VTAIL.n81 9.3005
R1425 VTAIL.n65 VTAIL.n64 9.3005
R1426 VTAIL.n88 VTAIL.n87 9.3005
R1427 VTAIL.n90 VTAIL.n89 9.3005
R1428 VTAIL.n62 VTAIL.n59 9.3005
R1429 VTAIL.n105 VTAIL.n104 9.3005
R1430 VTAIL.n56 VTAIL.n55 9.3005
R1431 VTAIL.n99 VTAIL.n98 9.3005
R1432 VTAIL.n97 VTAIL.n96 9.3005
R1433 VTAIL.n186 VTAIL.n185 8.92171
R1434 VTAIL.n24 VTAIL.n23 8.92171
R1435 VTAIL.n133 VTAIL.n132 8.92171
R1436 VTAIL.n79 VTAIL.n78 8.92171
R1437 VTAIL.n182 VTAIL.n176 8.14595
R1438 VTAIL.n20 VTAIL.n14 8.14595
R1439 VTAIL.n129 VTAIL.n123 8.14595
R1440 VTAIL.n75 VTAIL.n69 8.14595
R1441 VTAIL.n181 VTAIL.n178 7.3702
R1442 VTAIL.n19 VTAIL.n16 7.3702
R1443 VTAIL.n128 VTAIL.n125 7.3702
R1444 VTAIL.n74 VTAIL.n71 7.3702
R1445 VTAIL.n182 VTAIL.n181 5.81868
R1446 VTAIL.n20 VTAIL.n19 5.81868
R1447 VTAIL.n129 VTAIL.n128 5.81868
R1448 VTAIL.n75 VTAIL.n74 5.81868
R1449 VTAIL.n185 VTAIL.n176 5.04292
R1450 VTAIL.n23 VTAIL.n14 5.04292
R1451 VTAIL.n132 VTAIL.n123 5.04292
R1452 VTAIL.n78 VTAIL.n69 5.04292
R1453 VTAIL.n186 VTAIL.n174 4.26717
R1454 VTAIL.n24 VTAIL.n12 4.26717
R1455 VTAIL.n133 VTAIL.n121 4.26717
R1456 VTAIL.n79 VTAIL.n67 4.26717
R1457 VTAIL.n190 VTAIL.n189 3.49141
R1458 VTAIL.n214 VTAIL.n162 3.49141
R1459 VTAIL.n28 VTAIL.n27 3.49141
R1460 VTAIL.n52 VTAIL.n0 3.49141
R1461 VTAIL.n160 VTAIL.n108 3.49141
R1462 VTAIL.n137 VTAIL.n136 3.49141
R1463 VTAIL.n106 VTAIL.n54 3.49141
R1464 VTAIL.n83 VTAIL.n82 3.49141
R1465 VTAIL.n180 VTAIL.n179 2.84303
R1466 VTAIL.n18 VTAIL.n17 2.84303
R1467 VTAIL.n127 VTAIL.n126 2.84303
R1468 VTAIL.n73 VTAIL.n72 2.84303
R1469 VTAIL.n193 VTAIL.n172 2.71565
R1470 VTAIL.n212 VTAIL.n211 2.71565
R1471 VTAIL.n31 VTAIL.n10 2.71565
R1472 VTAIL.n50 VTAIL.n49 2.71565
R1473 VTAIL.n158 VTAIL.n157 2.71565
R1474 VTAIL.n140 VTAIL.n119 2.71565
R1475 VTAIL.n104 VTAIL.n103 2.71565
R1476 VTAIL.n86 VTAIL.n65 2.71565
R1477 VTAIL.n161 VTAIL.n107 2.00481
R1478 VTAIL.n194 VTAIL.n170 1.93989
R1479 VTAIL.n208 VTAIL.n164 1.93989
R1480 VTAIL.n32 VTAIL.n8 1.93989
R1481 VTAIL.n46 VTAIL.n2 1.93989
R1482 VTAIL.n154 VTAIL.n110 1.93989
R1483 VTAIL.n141 VTAIL.n117 1.93989
R1484 VTAIL.n100 VTAIL.n56 1.93989
R1485 VTAIL.n87 VTAIL.n63 1.93989
R1486 VTAIL VTAIL.n53 1.29576
R1487 VTAIL.n199 VTAIL.n197 1.16414
R1488 VTAIL.n207 VTAIL.n166 1.16414
R1489 VTAIL.n37 VTAIL.n35 1.16414
R1490 VTAIL.n45 VTAIL.n4 1.16414
R1491 VTAIL.n153 VTAIL.n112 1.16414
R1492 VTAIL.n145 VTAIL.n144 1.16414
R1493 VTAIL.n99 VTAIL.n58 1.16414
R1494 VTAIL.n91 VTAIL.n90 1.16414
R1495 VTAIL VTAIL.n215 0.709552
R1496 VTAIL.n198 VTAIL.n168 0.388379
R1497 VTAIL.n204 VTAIL.n203 0.388379
R1498 VTAIL.n36 VTAIL.n6 0.388379
R1499 VTAIL.n42 VTAIL.n41 0.388379
R1500 VTAIL.n150 VTAIL.n149 0.388379
R1501 VTAIL.n116 VTAIL.n114 0.388379
R1502 VTAIL.n96 VTAIL.n95 0.388379
R1503 VTAIL.n62 VTAIL.n60 0.388379
R1504 VTAIL.n180 VTAIL.n175 0.155672
R1505 VTAIL.n187 VTAIL.n175 0.155672
R1506 VTAIL.n188 VTAIL.n187 0.155672
R1507 VTAIL.n188 VTAIL.n171 0.155672
R1508 VTAIL.n195 VTAIL.n171 0.155672
R1509 VTAIL.n196 VTAIL.n195 0.155672
R1510 VTAIL.n196 VTAIL.n167 0.155672
R1511 VTAIL.n205 VTAIL.n167 0.155672
R1512 VTAIL.n206 VTAIL.n205 0.155672
R1513 VTAIL.n206 VTAIL.n163 0.155672
R1514 VTAIL.n213 VTAIL.n163 0.155672
R1515 VTAIL.n18 VTAIL.n13 0.155672
R1516 VTAIL.n25 VTAIL.n13 0.155672
R1517 VTAIL.n26 VTAIL.n25 0.155672
R1518 VTAIL.n26 VTAIL.n9 0.155672
R1519 VTAIL.n33 VTAIL.n9 0.155672
R1520 VTAIL.n34 VTAIL.n33 0.155672
R1521 VTAIL.n34 VTAIL.n5 0.155672
R1522 VTAIL.n43 VTAIL.n5 0.155672
R1523 VTAIL.n44 VTAIL.n43 0.155672
R1524 VTAIL.n44 VTAIL.n1 0.155672
R1525 VTAIL.n51 VTAIL.n1 0.155672
R1526 VTAIL.n159 VTAIL.n109 0.155672
R1527 VTAIL.n152 VTAIL.n109 0.155672
R1528 VTAIL.n152 VTAIL.n151 0.155672
R1529 VTAIL.n151 VTAIL.n113 0.155672
R1530 VTAIL.n143 VTAIL.n113 0.155672
R1531 VTAIL.n143 VTAIL.n142 0.155672
R1532 VTAIL.n142 VTAIL.n118 0.155672
R1533 VTAIL.n135 VTAIL.n118 0.155672
R1534 VTAIL.n135 VTAIL.n134 0.155672
R1535 VTAIL.n134 VTAIL.n122 0.155672
R1536 VTAIL.n127 VTAIL.n122 0.155672
R1537 VTAIL.n105 VTAIL.n55 0.155672
R1538 VTAIL.n98 VTAIL.n55 0.155672
R1539 VTAIL.n98 VTAIL.n97 0.155672
R1540 VTAIL.n97 VTAIL.n59 0.155672
R1541 VTAIL.n89 VTAIL.n59 0.155672
R1542 VTAIL.n89 VTAIL.n88 0.155672
R1543 VTAIL.n88 VTAIL.n64 0.155672
R1544 VTAIL.n81 VTAIL.n64 0.155672
R1545 VTAIL.n81 VTAIL.n80 0.155672
R1546 VTAIL.n80 VTAIL.n68 0.155672
R1547 VTAIL.n73 VTAIL.n68 0.155672
R1548 VDD2.n101 VDD2.n53 289.615
R1549 VDD2.n48 VDD2.n0 289.615
R1550 VDD2.n102 VDD2.n101 185
R1551 VDD2.n100 VDD2.n99 185
R1552 VDD2.n57 VDD2.n56 185
R1553 VDD2.n94 VDD2.n93 185
R1554 VDD2.n92 VDD2.n59 185
R1555 VDD2.n91 VDD2.n90 185
R1556 VDD2.n62 VDD2.n60 185
R1557 VDD2.n85 VDD2.n84 185
R1558 VDD2.n83 VDD2.n82 185
R1559 VDD2.n66 VDD2.n65 185
R1560 VDD2.n77 VDD2.n76 185
R1561 VDD2.n75 VDD2.n74 185
R1562 VDD2.n70 VDD2.n69 185
R1563 VDD2.n16 VDD2.n15 185
R1564 VDD2.n21 VDD2.n20 185
R1565 VDD2.n23 VDD2.n22 185
R1566 VDD2.n12 VDD2.n11 185
R1567 VDD2.n29 VDD2.n28 185
R1568 VDD2.n31 VDD2.n30 185
R1569 VDD2.n8 VDD2.n7 185
R1570 VDD2.n38 VDD2.n37 185
R1571 VDD2.n39 VDD2.n6 185
R1572 VDD2.n41 VDD2.n40 185
R1573 VDD2.n4 VDD2.n3 185
R1574 VDD2.n47 VDD2.n46 185
R1575 VDD2.n49 VDD2.n48 185
R1576 VDD2.n71 VDD2.t1 149.524
R1577 VDD2.n17 VDD2.t0 149.524
R1578 VDD2.n101 VDD2.n100 104.615
R1579 VDD2.n100 VDD2.n56 104.615
R1580 VDD2.n93 VDD2.n56 104.615
R1581 VDD2.n93 VDD2.n92 104.615
R1582 VDD2.n92 VDD2.n91 104.615
R1583 VDD2.n91 VDD2.n60 104.615
R1584 VDD2.n84 VDD2.n60 104.615
R1585 VDD2.n84 VDD2.n83 104.615
R1586 VDD2.n83 VDD2.n65 104.615
R1587 VDD2.n76 VDD2.n65 104.615
R1588 VDD2.n76 VDD2.n75 104.615
R1589 VDD2.n75 VDD2.n69 104.615
R1590 VDD2.n21 VDD2.n15 104.615
R1591 VDD2.n22 VDD2.n21 104.615
R1592 VDD2.n22 VDD2.n11 104.615
R1593 VDD2.n29 VDD2.n11 104.615
R1594 VDD2.n30 VDD2.n29 104.615
R1595 VDD2.n30 VDD2.n7 104.615
R1596 VDD2.n38 VDD2.n7 104.615
R1597 VDD2.n39 VDD2.n38 104.615
R1598 VDD2.n40 VDD2.n39 104.615
R1599 VDD2.n40 VDD2.n3 104.615
R1600 VDD2.n47 VDD2.n3 104.615
R1601 VDD2.n48 VDD2.n47 104.615
R1602 VDD2.n106 VDD2.n52 90.2861
R1603 VDD2.t1 VDD2.n69 52.3082
R1604 VDD2.t0 VDD2.n15 52.3082
R1605 VDD2.n106 VDD2.n105 51.7732
R1606 VDD2.n94 VDD2.n59 13.1884
R1607 VDD2.n41 VDD2.n6 13.1884
R1608 VDD2.n95 VDD2.n57 12.8005
R1609 VDD2.n90 VDD2.n61 12.8005
R1610 VDD2.n37 VDD2.n36 12.8005
R1611 VDD2.n42 VDD2.n4 12.8005
R1612 VDD2.n99 VDD2.n98 12.0247
R1613 VDD2.n89 VDD2.n62 12.0247
R1614 VDD2.n35 VDD2.n8 12.0247
R1615 VDD2.n46 VDD2.n45 12.0247
R1616 VDD2.n102 VDD2.n55 11.249
R1617 VDD2.n86 VDD2.n85 11.249
R1618 VDD2.n32 VDD2.n31 11.249
R1619 VDD2.n49 VDD2.n2 11.249
R1620 VDD2.n103 VDD2.n53 10.4732
R1621 VDD2.n82 VDD2.n64 10.4732
R1622 VDD2.n28 VDD2.n10 10.4732
R1623 VDD2.n50 VDD2.n0 10.4732
R1624 VDD2.n71 VDD2.n70 10.2747
R1625 VDD2.n17 VDD2.n16 10.2747
R1626 VDD2.n81 VDD2.n66 9.69747
R1627 VDD2.n27 VDD2.n12 9.69747
R1628 VDD2.n105 VDD2.n104 9.45567
R1629 VDD2.n52 VDD2.n51 9.45567
R1630 VDD2.n73 VDD2.n72 9.3005
R1631 VDD2.n68 VDD2.n67 9.3005
R1632 VDD2.n79 VDD2.n78 9.3005
R1633 VDD2.n81 VDD2.n80 9.3005
R1634 VDD2.n64 VDD2.n63 9.3005
R1635 VDD2.n87 VDD2.n86 9.3005
R1636 VDD2.n89 VDD2.n88 9.3005
R1637 VDD2.n61 VDD2.n58 9.3005
R1638 VDD2.n104 VDD2.n103 9.3005
R1639 VDD2.n55 VDD2.n54 9.3005
R1640 VDD2.n98 VDD2.n97 9.3005
R1641 VDD2.n96 VDD2.n95 9.3005
R1642 VDD2.n51 VDD2.n50 9.3005
R1643 VDD2.n2 VDD2.n1 9.3005
R1644 VDD2.n45 VDD2.n44 9.3005
R1645 VDD2.n43 VDD2.n42 9.3005
R1646 VDD2.n19 VDD2.n18 9.3005
R1647 VDD2.n14 VDD2.n13 9.3005
R1648 VDD2.n25 VDD2.n24 9.3005
R1649 VDD2.n27 VDD2.n26 9.3005
R1650 VDD2.n10 VDD2.n9 9.3005
R1651 VDD2.n33 VDD2.n32 9.3005
R1652 VDD2.n35 VDD2.n34 9.3005
R1653 VDD2.n36 VDD2.n5 9.3005
R1654 VDD2.n78 VDD2.n77 8.92171
R1655 VDD2.n24 VDD2.n23 8.92171
R1656 VDD2.n74 VDD2.n68 8.14595
R1657 VDD2.n20 VDD2.n14 8.14595
R1658 VDD2.n73 VDD2.n70 7.3702
R1659 VDD2.n19 VDD2.n16 7.3702
R1660 VDD2.n74 VDD2.n73 5.81868
R1661 VDD2.n20 VDD2.n19 5.81868
R1662 VDD2.n77 VDD2.n68 5.04292
R1663 VDD2.n23 VDD2.n14 5.04292
R1664 VDD2.n78 VDD2.n66 4.26717
R1665 VDD2.n24 VDD2.n12 4.26717
R1666 VDD2.n105 VDD2.n53 3.49141
R1667 VDD2.n82 VDD2.n81 3.49141
R1668 VDD2.n28 VDD2.n27 3.49141
R1669 VDD2.n52 VDD2.n0 3.49141
R1670 VDD2.n72 VDD2.n71 2.84303
R1671 VDD2.n18 VDD2.n17 2.84303
R1672 VDD2.n103 VDD2.n102 2.71565
R1673 VDD2.n85 VDD2.n64 2.71565
R1674 VDD2.n31 VDD2.n10 2.71565
R1675 VDD2.n50 VDD2.n49 2.71565
R1676 VDD2.n99 VDD2.n55 1.93989
R1677 VDD2.n86 VDD2.n62 1.93989
R1678 VDD2.n32 VDD2.n8 1.93989
R1679 VDD2.n46 VDD2.n2 1.93989
R1680 VDD2.n98 VDD2.n57 1.16414
R1681 VDD2.n90 VDD2.n89 1.16414
R1682 VDD2.n37 VDD2.n35 1.16414
R1683 VDD2.n45 VDD2.n4 1.16414
R1684 VDD2 VDD2.n106 0.825931
R1685 VDD2.n95 VDD2.n94 0.388379
R1686 VDD2.n61 VDD2.n59 0.388379
R1687 VDD2.n36 VDD2.n6 0.388379
R1688 VDD2.n42 VDD2.n41 0.388379
R1689 VDD2.n104 VDD2.n54 0.155672
R1690 VDD2.n97 VDD2.n54 0.155672
R1691 VDD2.n97 VDD2.n96 0.155672
R1692 VDD2.n96 VDD2.n58 0.155672
R1693 VDD2.n88 VDD2.n58 0.155672
R1694 VDD2.n88 VDD2.n87 0.155672
R1695 VDD2.n87 VDD2.n63 0.155672
R1696 VDD2.n80 VDD2.n63 0.155672
R1697 VDD2.n80 VDD2.n79 0.155672
R1698 VDD2.n79 VDD2.n67 0.155672
R1699 VDD2.n72 VDD2.n67 0.155672
R1700 VDD2.n18 VDD2.n13 0.155672
R1701 VDD2.n25 VDD2.n13 0.155672
R1702 VDD2.n26 VDD2.n25 0.155672
R1703 VDD2.n26 VDD2.n9 0.155672
R1704 VDD2.n33 VDD2.n9 0.155672
R1705 VDD2.n34 VDD2.n33 0.155672
R1706 VDD2.n34 VDD2.n5 0.155672
R1707 VDD2.n43 VDD2.n5 0.155672
R1708 VDD2.n44 VDD2.n43 0.155672
R1709 VDD2.n44 VDD2.n1 0.155672
R1710 VDD2.n51 VDD2.n1 0.155672
R1711 VP.n0 VP.t0 159.118
R1712 VP.n0 VP.t1 114.222
R1713 VP VP.n0 0.52637
R1714 VDD1.n48 VDD1.n0 289.615
R1715 VDD1.n101 VDD1.n53 289.615
R1716 VDD1.n49 VDD1.n48 185
R1717 VDD1.n47 VDD1.n46 185
R1718 VDD1.n4 VDD1.n3 185
R1719 VDD1.n41 VDD1.n40 185
R1720 VDD1.n39 VDD1.n6 185
R1721 VDD1.n38 VDD1.n37 185
R1722 VDD1.n9 VDD1.n7 185
R1723 VDD1.n32 VDD1.n31 185
R1724 VDD1.n30 VDD1.n29 185
R1725 VDD1.n13 VDD1.n12 185
R1726 VDD1.n24 VDD1.n23 185
R1727 VDD1.n22 VDD1.n21 185
R1728 VDD1.n17 VDD1.n16 185
R1729 VDD1.n69 VDD1.n68 185
R1730 VDD1.n74 VDD1.n73 185
R1731 VDD1.n76 VDD1.n75 185
R1732 VDD1.n65 VDD1.n64 185
R1733 VDD1.n82 VDD1.n81 185
R1734 VDD1.n84 VDD1.n83 185
R1735 VDD1.n61 VDD1.n60 185
R1736 VDD1.n91 VDD1.n90 185
R1737 VDD1.n92 VDD1.n59 185
R1738 VDD1.n94 VDD1.n93 185
R1739 VDD1.n57 VDD1.n56 185
R1740 VDD1.n100 VDD1.n99 185
R1741 VDD1.n102 VDD1.n101 185
R1742 VDD1.n18 VDD1.t1 149.524
R1743 VDD1.n70 VDD1.t0 149.524
R1744 VDD1.n48 VDD1.n47 104.615
R1745 VDD1.n47 VDD1.n3 104.615
R1746 VDD1.n40 VDD1.n3 104.615
R1747 VDD1.n40 VDD1.n39 104.615
R1748 VDD1.n39 VDD1.n38 104.615
R1749 VDD1.n38 VDD1.n7 104.615
R1750 VDD1.n31 VDD1.n7 104.615
R1751 VDD1.n31 VDD1.n30 104.615
R1752 VDD1.n30 VDD1.n12 104.615
R1753 VDD1.n23 VDD1.n12 104.615
R1754 VDD1.n23 VDD1.n22 104.615
R1755 VDD1.n22 VDD1.n16 104.615
R1756 VDD1.n74 VDD1.n68 104.615
R1757 VDD1.n75 VDD1.n74 104.615
R1758 VDD1.n75 VDD1.n64 104.615
R1759 VDD1.n82 VDD1.n64 104.615
R1760 VDD1.n83 VDD1.n82 104.615
R1761 VDD1.n83 VDD1.n60 104.615
R1762 VDD1.n91 VDD1.n60 104.615
R1763 VDD1.n92 VDD1.n91 104.615
R1764 VDD1.n93 VDD1.n92 104.615
R1765 VDD1.n93 VDD1.n56 104.615
R1766 VDD1.n100 VDD1.n56 104.615
R1767 VDD1.n101 VDD1.n100 104.615
R1768 VDD1 VDD1.n105 91.5782
R1769 VDD1 VDD1.n52 52.5987
R1770 VDD1.t1 VDD1.n16 52.3082
R1771 VDD1.t0 VDD1.n68 52.3082
R1772 VDD1.n41 VDD1.n6 13.1884
R1773 VDD1.n94 VDD1.n59 13.1884
R1774 VDD1.n42 VDD1.n4 12.8005
R1775 VDD1.n37 VDD1.n8 12.8005
R1776 VDD1.n90 VDD1.n89 12.8005
R1777 VDD1.n95 VDD1.n57 12.8005
R1778 VDD1.n46 VDD1.n45 12.0247
R1779 VDD1.n36 VDD1.n9 12.0247
R1780 VDD1.n88 VDD1.n61 12.0247
R1781 VDD1.n99 VDD1.n98 12.0247
R1782 VDD1.n49 VDD1.n2 11.249
R1783 VDD1.n33 VDD1.n32 11.249
R1784 VDD1.n85 VDD1.n84 11.249
R1785 VDD1.n102 VDD1.n55 11.249
R1786 VDD1.n50 VDD1.n0 10.4732
R1787 VDD1.n29 VDD1.n11 10.4732
R1788 VDD1.n81 VDD1.n63 10.4732
R1789 VDD1.n103 VDD1.n53 10.4732
R1790 VDD1.n18 VDD1.n17 10.2747
R1791 VDD1.n70 VDD1.n69 10.2747
R1792 VDD1.n28 VDD1.n13 9.69747
R1793 VDD1.n80 VDD1.n65 9.69747
R1794 VDD1.n52 VDD1.n51 9.45567
R1795 VDD1.n105 VDD1.n104 9.45567
R1796 VDD1.n20 VDD1.n19 9.3005
R1797 VDD1.n15 VDD1.n14 9.3005
R1798 VDD1.n26 VDD1.n25 9.3005
R1799 VDD1.n28 VDD1.n27 9.3005
R1800 VDD1.n11 VDD1.n10 9.3005
R1801 VDD1.n34 VDD1.n33 9.3005
R1802 VDD1.n36 VDD1.n35 9.3005
R1803 VDD1.n8 VDD1.n5 9.3005
R1804 VDD1.n51 VDD1.n50 9.3005
R1805 VDD1.n2 VDD1.n1 9.3005
R1806 VDD1.n45 VDD1.n44 9.3005
R1807 VDD1.n43 VDD1.n42 9.3005
R1808 VDD1.n104 VDD1.n103 9.3005
R1809 VDD1.n55 VDD1.n54 9.3005
R1810 VDD1.n98 VDD1.n97 9.3005
R1811 VDD1.n96 VDD1.n95 9.3005
R1812 VDD1.n72 VDD1.n71 9.3005
R1813 VDD1.n67 VDD1.n66 9.3005
R1814 VDD1.n78 VDD1.n77 9.3005
R1815 VDD1.n80 VDD1.n79 9.3005
R1816 VDD1.n63 VDD1.n62 9.3005
R1817 VDD1.n86 VDD1.n85 9.3005
R1818 VDD1.n88 VDD1.n87 9.3005
R1819 VDD1.n89 VDD1.n58 9.3005
R1820 VDD1.n25 VDD1.n24 8.92171
R1821 VDD1.n77 VDD1.n76 8.92171
R1822 VDD1.n21 VDD1.n15 8.14595
R1823 VDD1.n73 VDD1.n67 8.14595
R1824 VDD1.n20 VDD1.n17 7.3702
R1825 VDD1.n72 VDD1.n69 7.3702
R1826 VDD1.n21 VDD1.n20 5.81868
R1827 VDD1.n73 VDD1.n72 5.81868
R1828 VDD1.n24 VDD1.n15 5.04292
R1829 VDD1.n76 VDD1.n67 5.04292
R1830 VDD1.n25 VDD1.n13 4.26717
R1831 VDD1.n77 VDD1.n65 4.26717
R1832 VDD1.n52 VDD1.n0 3.49141
R1833 VDD1.n29 VDD1.n28 3.49141
R1834 VDD1.n81 VDD1.n80 3.49141
R1835 VDD1.n105 VDD1.n53 3.49141
R1836 VDD1.n19 VDD1.n18 2.84303
R1837 VDD1.n71 VDD1.n70 2.84303
R1838 VDD1.n50 VDD1.n49 2.71565
R1839 VDD1.n32 VDD1.n11 2.71565
R1840 VDD1.n84 VDD1.n63 2.71565
R1841 VDD1.n103 VDD1.n102 2.71565
R1842 VDD1.n46 VDD1.n2 1.93989
R1843 VDD1.n33 VDD1.n9 1.93989
R1844 VDD1.n85 VDD1.n61 1.93989
R1845 VDD1.n99 VDD1.n55 1.93989
R1846 VDD1.n45 VDD1.n4 1.16414
R1847 VDD1.n37 VDD1.n36 1.16414
R1848 VDD1.n90 VDD1.n88 1.16414
R1849 VDD1.n98 VDD1.n57 1.16414
R1850 VDD1.n42 VDD1.n41 0.388379
R1851 VDD1.n8 VDD1.n6 0.388379
R1852 VDD1.n89 VDD1.n59 0.388379
R1853 VDD1.n95 VDD1.n94 0.388379
R1854 VDD1.n51 VDD1.n1 0.155672
R1855 VDD1.n44 VDD1.n1 0.155672
R1856 VDD1.n44 VDD1.n43 0.155672
R1857 VDD1.n43 VDD1.n5 0.155672
R1858 VDD1.n35 VDD1.n5 0.155672
R1859 VDD1.n35 VDD1.n34 0.155672
R1860 VDD1.n34 VDD1.n10 0.155672
R1861 VDD1.n27 VDD1.n10 0.155672
R1862 VDD1.n27 VDD1.n26 0.155672
R1863 VDD1.n26 VDD1.n14 0.155672
R1864 VDD1.n19 VDD1.n14 0.155672
R1865 VDD1.n71 VDD1.n66 0.155672
R1866 VDD1.n78 VDD1.n66 0.155672
R1867 VDD1.n79 VDD1.n78 0.155672
R1868 VDD1.n79 VDD1.n62 0.155672
R1869 VDD1.n86 VDD1.n62 0.155672
R1870 VDD1.n87 VDD1.n86 0.155672
R1871 VDD1.n87 VDD1.n58 0.155672
R1872 VDD1.n96 VDD1.n58 0.155672
R1873 VDD1.n97 VDD1.n96 0.155672
R1874 VDD1.n97 VDD1.n54 0.155672
R1875 VDD1.n104 VDD1.n54 0.155672
C0 VTAIL VP 2.26446f
C1 VTAIL VN 2.25023f
C2 VDD1 VP 2.66267f
C3 VDD1 VN 0.148411f
C4 VDD2 VP 0.359403f
C5 VDD1 VTAIL 4.69795f
C6 VDD2 VN 2.45367f
C7 VDD2 VTAIL 4.75372f
C8 VDD2 VDD1 0.751153f
C9 VN VP 5.40439f
C10 VDD2 B 4.314431f
C11 VDD1 B 7.07909f
C12 VTAIL B 6.895871f
C13 VN B 10.96184f
C14 VP B 7.067708f
C15 VDD1.n0 B 0.029777f
C16 VDD1.n1 B 0.020884f
C17 VDD1.n2 B 0.011222f
C18 VDD1.n3 B 0.026525f
C19 VDD1.n4 B 0.011882f
C20 VDD1.n5 B 0.020884f
C21 VDD1.n6 B 0.011552f
C22 VDD1.n7 B 0.026525f
C23 VDD1.n8 B 0.011222f
C24 VDD1.n9 B 0.011882f
C25 VDD1.n10 B 0.020884f
C26 VDD1.n11 B 0.011222f
C27 VDD1.n12 B 0.026525f
C28 VDD1.n13 B 0.011882f
C29 VDD1.n14 B 0.020884f
C30 VDD1.n15 B 0.011222f
C31 VDD1.n16 B 0.019894f
C32 VDD1.n17 B 0.018752f
C33 VDD1.t1 B 0.044589f
C34 VDD1.n18 B 0.135423f
C35 VDD1.n19 B 0.87801f
C36 VDD1.n20 B 0.011222f
C37 VDD1.n21 B 0.011882f
C38 VDD1.n22 B 0.026525f
C39 VDD1.n23 B 0.026525f
C40 VDD1.n24 B 0.011882f
C41 VDD1.n25 B 0.011222f
C42 VDD1.n26 B 0.020884f
C43 VDD1.n27 B 0.020884f
C44 VDD1.n28 B 0.011222f
C45 VDD1.n29 B 0.011882f
C46 VDD1.n30 B 0.026525f
C47 VDD1.n31 B 0.026525f
C48 VDD1.n32 B 0.011882f
C49 VDD1.n33 B 0.011222f
C50 VDD1.n34 B 0.020884f
C51 VDD1.n35 B 0.020884f
C52 VDD1.n36 B 0.011222f
C53 VDD1.n37 B 0.011882f
C54 VDD1.n38 B 0.026525f
C55 VDD1.n39 B 0.026525f
C56 VDD1.n40 B 0.026525f
C57 VDD1.n41 B 0.011552f
C58 VDD1.n42 B 0.011222f
C59 VDD1.n43 B 0.020884f
C60 VDD1.n44 B 0.020884f
C61 VDD1.n45 B 0.011222f
C62 VDD1.n46 B 0.011882f
C63 VDD1.n47 B 0.026525f
C64 VDD1.n48 B 0.058171f
C65 VDD1.n49 B 0.011882f
C66 VDD1.n50 B 0.011222f
C67 VDD1.n51 B 0.052553f
C68 VDD1.n52 B 0.048683f
C69 VDD1.n53 B 0.029777f
C70 VDD1.n54 B 0.020884f
C71 VDD1.n55 B 0.011222f
C72 VDD1.n56 B 0.026525f
C73 VDD1.n57 B 0.011882f
C74 VDD1.n58 B 0.020884f
C75 VDD1.n59 B 0.011552f
C76 VDD1.n60 B 0.026525f
C77 VDD1.n61 B 0.011882f
C78 VDD1.n62 B 0.020884f
C79 VDD1.n63 B 0.011222f
C80 VDD1.n64 B 0.026525f
C81 VDD1.n65 B 0.011882f
C82 VDD1.n66 B 0.020884f
C83 VDD1.n67 B 0.011222f
C84 VDD1.n68 B 0.019894f
C85 VDD1.n69 B 0.018752f
C86 VDD1.t0 B 0.044589f
C87 VDD1.n70 B 0.135423f
C88 VDD1.n71 B 0.87801f
C89 VDD1.n72 B 0.011222f
C90 VDD1.n73 B 0.011882f
C91 VDD1.n74 B 0.026525f
C92 VDD1.n75 B 0.026525f
C93 VDD1.n76 B 0.011882f
C94 VDD1.n77 B 0.011222f
C95 VDD1.n78 B 0.020884f
C96 VDD1.n79 B 0.020884f
C97 VDD1.n80 B 0.011222f
C98 VDD1.n81 B 0.011882f
C99 VDD1.n82 B 0.026525f
C100 VDD1.n83 B 0.026525f
C101 VDD1.n84 B 0.011882f
C102 VDD1.n85 B 0.011222f
C103 VDD1.n86 B 0.020884f
C104 VDD1.n87 B 0.020884f
C105 VDD1.n88 B 0.011222f
C106 VDD1.n89 B 0.011222f
C107 VDD1.n90 B 0.011882f
C108 VDD1.n91 B 0.026525f
C109 VDD1.n92 B 0.026525f
C110 VDD1.n93 B 0.026525f
C111 VDD1.n94 B 0.011552f
C112 VDD1.n95 B 0.011222f
C113 VDD1.n96 B 0.020884f
C114 VDD1.n97 B 0.020884f
C115 VDD1.n98 B 0.011222f
C116 VDD1.n99 B 0.011882f
C117 VDD1.n100 B 0.026525f
C118 VDD1.n101 B 0.058171f
C119 VDD1.n102 B 0.011882f
C120 VDD1.n103 B 0.011222f
C121 VDD1.n104 B 0.052553f
C122 VDD1.n105 B 0.619893f
C123 VP.t0 B 3.56057f
C124 VP.t1 B 2.92069f
C125 VP.n0 B 3.82061f
C126 VDD2.n0 B 0.029685f
C127 VDD2.n1 B 0.020819f
C128 VDD2.n2 B 0.011187f
C129 VDD2.n3 B 0.026443f
C130 VDD2.n4 B 0.011845f
C131 VDD2.n5 B 0.020819f
C132 VDD2.n6 B 0.011516f
C133 VDD2.n7 B 0.026443f
C134 VDD2.n8 B 0.011845f
C135 VDD2.n9 B 0.020819f
C136 VDD2.n10 B 0.011187f
C137 VDD2.n11 B 0.026443f
C138 VDD2.n12 B 0.011845f
C139 VDD2.n13 B 0.020819f
C140 VDD2.n14 B 0.011187f
C141 VDD2.n15 B 0.019832f
C142 VDD2.n16 B 0.018693f
C143 VDD2.t0 B 0.04445f
C144 VDD2.n17 B 0.135001f
C145 VDD2.n18 B 0.875268f
C146 VDD2.n19 B 0.011187f
C147 VDD2.n20 B 0.011845f
C148 VDD2.n21 B 0.026443f
C149 VDD2.n22 B 0.026443f
C150 VDD2.n23 B 0.011845f
C151 VDD2.n24 B 0.011187f
C152 VDD2.n25 B 0.020819f
C153 VDD2.n26 B 0.020819f
C154 VDD2.n27 B 0.011187f
C155 VDD2.n28 B 0.011845f
C156 VDD2.n29 B 0.026443f
C157 VDD2.n30 B 0.026443f
C158 VDD2.n31 B 0.011845f
C159 VDD2.n32 B 0.011187f
C160 VDD2.n33 B 0.020819f
C161 VDD2.n34 B 0.020819f
C162 VDD2.n35 B 0.011187f
C163 VDD2.n36 B 0.011187f
C164 VDD2.n37 B 0.011845f
C165 VDD2.n38 B 0.026443f
C166 VDD2.n39 B 0.026443f
C167 VDD2.n40 B 0.026443f
C168 VDD2.n41 B 0.011516f
C169 VDD2.n42 B 0.011187f
C170 VDD2.n43 B 0.020819f
C171 VDD2.n44 B 0.020819f
C172 VDD2.n45 B 0.011187f
C173 VDD2.n46 B 0.011845f
C174 VDD2.n47 B 0.026443f
C175 VDD2.n48 B 0.057989f
C176 VDD2.n49 B 0.011845f
C177 VDD2.n50 B 0.011187f
C178 VDD2.n51 B 0.052389f
C179 VDD2.n52 B 0.575032f
C180 VDD2.n53 B 0.029685f
C181 VDD2.n54 B 0.020819f
C182 VDD2.n55 B 0.011187f
C183 VDD2.n56 B 0.026443f
C184 VDD2.n57 B 0.011845f
C185 VDD2.n58 B 0.020819f
C186 VDD2.n59 B 0.011516f
C187 VDD2.n60 B 0.026443f
C188 VDD2.n61 B 0.011187f
C189 VDD2.n62 B 0.011845f
C190 VDD2.n63 B 0.020819f
C191 VDD2.n64 B 0.011187f
C192 VDD2.n65 B 0.026443f
C193 VDD2.n66 B 0.011845f
C194 VDD2.n67 B 0.020819f
C195 VDD2.n68 B 0.011187f
C196 VDD2.n69 B 0.019832f
C197 VDD2.n70 B 0.018693f
C198 VDD2.t1 B 0.04445f
C199 VDD2.n71 B 0.135001f
C200 VDD2.n72 B 0.875268f
C201 VDD2.n73 B 0.011187f
C202 VDD2.n74 B 0.011845f
C203 VDD2.n75 B 0.026443f
C204 VDD2.n76 B 0.026443f
C205 VDD2.n77 B 0.011845f
C206 VDD2.n78 B 0.011187f
C207 VDD2.n79 B 0.020819f
C208 VDD2.n80 B 0.020819f
C209 VDD2.n81 B 0.011187f
C210 VDD2.n82 B 0.011845f
C211 VDD2.n83 B 0.026443f
C212 VDD2.n84 B 0.026443f
C213 VDD2.n85 B 0.011845f
C214 VDD2.n86 B 0.011187f
C215 VDD2.n87 B 0.020819f
C216 VDD2.n88 B 0.020819f
C217 VDD2.n89 B 0.011187f
C218 VDD2.n90 B 0.011845f
C219 VDD2.n91 B 0.026443f
C220 VDD2.n92 B 0.026443f
C221 VDD2.n93 B 0.026443f
C222 VDD2.n94 B 0.011516f
C223 VDD2.n95 B 0.011187f
C224 VDD2.n96 B 0.020819f
C225 VDD2.n97 B 0.020819f
C226 VDD2.n98 B 0.011187f
C227 VDD2.n99 B 0.011845f
C228 VDD2.n100 B 0.026443f
C229 VDD2.n101 B 0.057989f
C230 VDD2.n102 B 0.011845f
C231 VDD2.n103 B 0.011187f
C232 VDD2.n104 B 0.052389f
C233 VDD2.n105 B 0.046995f
C234 VDD2.n106 B 2.50288f
C235 VTAIL.n0 B 0.031034f
C236 VTAIL.n1 B 0.021766f
C237 VTAIL.n2 B 0.011696f
C238 VTAIL.n3 B 0.027645f
C239 VTAIL.n4 B 0.012384f
C240 VTAIL.n5 B 0.021766f
C241 VTAIL.n6 B 0.01204f
C242 VTAIL.n7 B 0.027645f
C243 VTAIL.n8 B 0.012384f
C244 VTAIL.n9 B 0.021766f
C245 VTAIL.n10 B 0.011696f
C246 VTAIL.n11 B 0.027645f
C247 VTAIL.n12 B 0.012384f
C248 VTAIL.n13 B 0.021766f
C249 VTAIL.n14 B 0.011696f
C250 VTAIL.n15 B 0.020734f
C251 VTAIL.n16 B 0.019543f
C252 VTAIL.t0 B 0.046471f
C253 VTAIL.n17 B 0.141139f
C254 VTAIL.n18 B 0.915066f
C255 VTAIL.n19 B 0.011696f
C256 VTAIL.n20 B 0.012384f
C257 VTAIL.n21 B 0.027645f
C258 VTAIL.n22 B 0.027645f
C259 VTAIL.n23 B 0.012384f
C260 VTAIL.n24 B 0.011696f
C261 VTAIL.n25 B 0.021766f
C262 VTAIL.n26 B 0.021766f
C263 VTAIL.n27 B 0.011696f
C264 VTAIL.n28 B 0.012384f
C265 VTAIL.n29 B 0.027645f
C266 VTAIL.n30 B 0.027645f
C267 VTAIL.n31 B 0.012384f
C268 VTAIL.n32 B 0.011696f
C269 VTAIL.n33 B 0.021766f
C270 VTAIL.n34 B 0.021766f
C271 VTAIL.n35 B 0.011696f
C272 VTAIL.n36 B 0.011696f
C273 VTAIL.n37 B 0.012384f
C274 VTAIL.n38 B 0.027645f
C275 VTAIL.n39 B 0.027645f
C276 VTAIL.n40 B 0.027645f
C277 VTAIL.n41 B 0.01204f
C278 VTAIL.n42 B 0.011696f
C279 VTAIL.n43 B 0.021766f
C280 VTAIL.n44 B 0.021766f
C281 VTAIL.n45 B 0.011696f
C282 VTAIL.n46 B 0.012384f
C283 VTAIL.n47 B 0.027645f
C284 VTAIL.n48 B 0.060626f
C285 VTAIL.n49 B 0.012384f
C286 VTAIL.n50 B 0.011696f
C287 VTAIL.n51 B 0.054771f
C288 VTAIL.n52 B 0.034134f
C289 VTAIL.n53 B 1.44935f
C290 VTAIL.n54 B 0.031034f
C291 VTAIL.n55 B 0.021766f
C292 VTAIL.n56 B 0.011696f
C293 VTAIL.n57 B 0.027645f
C294 VTAIL.n58 B 0.012384f
C295 VTAIL.n59 B 0.021766f
C296 VTAIL.n60 B 0.01204f
C297 VTAIL.n61 B 0.027645f
C298 VTAIL.n62 B 0.011696f
C299 VTAIL.n63 B 0.012384f
C300 VTAIL.n64 B 0.021766f
C301 VTAIL.n65 B 0.011696f
C302 VTAIL.n66 B 0.027645f
C303 VTAIL.n67 B 0.012384f
C304 VTAIL.n68 B 0.021766f
C305 VTAIL.n69 B 0.011696f
C306 VTAIL.n70 B 0.020734f
C307 VTAIL.n71 B 0.019543f
C308 VTAIL.t2 B 0.046471f
C309 VTAIL.n72 B 0.141139f
C310 VTAIL.n73 B 0.915066f
C311 VTAIL.n74 B 0.011696f
C312 VTAIL.n75 B 0.012384f
C313 VTAIL.n76 B 0.027645f
C314 VTAIL.n77 B 0.027645f
C315 VTAIL.n78 B 0.012384f
C316 VTAIL.n79 B 0.011696f
C317 VTAIL.n80 B 0.021766f
C318 VTAIL.n81 B 0.021766f
C319 VTAIL.n82 B 0.011696f
C320 VTAIL.n83 B 0.012384f
C321 VTAIL.n84 B 0.027645f
C322 VTAIL.n85 B 0.027645f
C323 VTAIL.n86 B 0.012384f
C324 VTAIL.n87 B 0.011696f
C325 VTAIL.n88 B 0.021766f
C326 VTAIL.n89 B 0.021766f
C327 VTAIL.n90 B 0.011696f
C328 VTAIL.n91 B 0.012384f
C329 VTAIL.n92 B 0.027645f
C330 VTAIL.n93 B 0.027645f
C331 VTAIL.n94 B 0.027645f
C332 VTAIL.n95 B 0.01204f
C333 VTAIL.n96 B 0.011696f
C334 VTAIL.n97 B 0.021766f
C335 VTAIL.n98 B 0.021766f
C336 VTAIL.n99 B 0.011696f
C337 VTAIL.n100 B 0.012384f
C338 VTAIL.n101 B 0.027645f
C339 VTAIL.n102 B 0.060626f
C340 VTAIL.n103 B 0.012384f
C341 VTAIL.n104 B 0.011696f
C342 VTAIL.n105 B 0.054771f
C343 VTAIL.n106 B 0.034134f
C344 VTAIL.n107 B 1.49908f
C345 VTAIL.n108 B 0.031034f
C346 VTAIL.n109 B 0.021766f
C347 VTAIL.n110 B 0.011696f
C348 VTAIL.n111 B 0.027645f
C349 VTAIL.n112 B 0.012384f
C350 VTAIL.n113 B 0.021766f
C351 VTAIL.n114 B 0.01204f
C352 VTAIL.n115 B 0.027645f
C353 VTAIL.n116 B 0.011696f
C354 VTAIL.n117 B 0.012384f
C355 VTAIL.n118 B 0.021766f
C356 VTAIL.n119 B 0.011696f
C357 VTAIL.n120 B 0.027645f
C358 VTAIL.n121 B 0.012384f
C359 VTAIL.n122 B 0.021766f
C360 VTAIL.n123 B 0.011696f
C361 VTAIL.n124 B 0.020734f
C362 VTAIL.n125 B 0.019543f
C363 VTAIL.t1 B 0.046471f
C364 VTAIL.n126 B 0.141139f
C365 VTAIL.n127 B 0.915066f
C366 VTAIL.n128 B 0.011696f
C367 VTAIL.n129 B 0.012384f
C368 VTAIL.n130 B 0.027645f
C369 VTAIL.n131 B 0.027645f
C370 VTAIL.n132 B 0.012384f
C371 VTAIL.n133 B 0.011696f
C372 VTAIL.n134 B 0.021766f
C373 VTAIL.n135 B 0.021766f
C374 VTAIL.n136 B 0.011696f
C375 VTAIL.n137 B 0.012384f
C376 VTAIL.n138 B 0.027645f
C377 VTAIL.n139 B 0.027645f
C378 VTAIL.n140 B 0.012384f
C379 VTAIL.n141 B 0.011696f
C380 VTAIL.n142 B 0.021766f
C381 VTAIL.n143 B 0.021766f
C382 VTAIL.n144 B 0.011696f
C383 VTAIL.n145 B 0.012384f
C384 VTAIL.n146 B 0.027645f
C385 VTAIL.n147 B 0.027645f
C386 VTAIL.n148 B 0.027645f
C387 VTAIL.n149 B 0.01204f
C388 VTAIL.n150 B 0.011696f
C389 VTAIL.n151 B 0.021766f
C390 VTAIL.n152 B 0.021766f
C391 VTAIL.n153 B 0.011696f
C392 VTAIL.n154 B 0.012384f
C393 VTAIL.n155 B 0.027645f
C394 VTAIL.n156 B 0.060626f
C395 VTAIL.n157 B 0.012384f
C396 VTAIL.n158 B 0.011696f
C397 VTAIL.n159 B 0.054771f
C398 VTAIL.n160 B 0.034134f
C399 VTAIL.n161 B 1.28384f
C400 VTAIL.n162 B 0.031034f
C401 VTAIL.n163 B 0.021766f
C402 VTAIL.n164 B 0.011696f
C403 VTAIL.n165 B 0.027645f
C404 VTAIL.n166 B 0.012384f
C405 VTAIL.n167 B 0.021766f
C406 VTAIL.n168 B 0.01204f
C407 VTAIL.n169 B 0.027645f
C408 VTAIL.n170 B 0.012384f
C409 VTAIL.n171 B 0.021766f
C410 VTAIL.n172 B 0.011696f
C411 VTAIL.n173 B 0.027645f
C412 VTAIL.n174 B 0.012384f
C413 VTAIL.n175 B 0.021766f
C414 VTAIL.n176 B 0.011696f
C415 VTAIL.n177 B 0.020734f
C416 VTAIL.n178 B 0.019543f
C417 VTAIL.t3 B 0.046471f
C418 VTAIL.n179 B 0.141139f
C419 VTAIL.n180 B 0.915066f
C420 VTAIL.n181 B 0.011696f
C421 VTAIL.n182 B 0.012384f
C422 VTAIL.n183 B 0.027645f
C423 VTAIL.n184 B 0.027645f
C424 VTAIL.n185 B 0.012384f
C425 VTAIL.n186 B 0.011696f
C426 VTAIL.n187 B 0.021766f
C427 VTAIL.n188 B 0.021766f
C428 VTAIL.n189 B 0.011696f
C429 VTAIL.n190 B 0.012384f
C430 VTAIL.n191 B 0.027645f
C431 VTAIL.n192 B 0.027645f
C432 VTAIL.n193 B 0.012384f
C433 VTAIL.n194 B 0.011696f
C434 VTAIL.n195 B 0.021766f
C435 VTAIL.n196 B 0.021766f
C436 VTAIL.n197 B 0.011696f
C437 VTAIL.n198 B 0.011696f
C438 VTAIL.n199 B 0.012384f
C439 VTAIL.n200 B 0.027645f
C440 VTAIL.n201 B 0.027645f
C441 VTAIL.n202 B 0.027645f
C442 VTAIL.n203 B 0.01204f
C443 VTAIL.n204 B 0.011696f
C444 VTAIL.n205 B 0.021766f
C445 VTAIL.n206 B 0.021766f
C446 VTAIL.n207 B 0.011696f
C447 VTAIL.n208 B 0.012384f
C448 VTAIL.n209 B 0.027645f
C449 VTAIL.n210 B 0.060626f
C450 VTAIL.n211 B 0.012384f
C451 VTAIL.n212 B 0.011696f
C452 VTAIL.n213 B 0.054771f
C453 VTAIL.n214 B 0.034134f
C454 VTAIL.n215 B 1.193f
C455 VN.t1 B 2.85759f
C456 VN.t0 B 3.47876f
.ends

