* NGSPICE file created from diff_pair_sample_0258.ext - technology: sky130A

.subckt diff_pair_sample_0258 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=0 ps=0 w=6.21 l=3.6
X1 B.t8 B.t6 B.t7 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=0 ps=0 w=6.21 l=3.6
X2 B.t5 B.t3 B.t4 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=0 ps=0 w=6.21 l=3.6
X3 VDD2.t1 VN.t0 VTAIL.t2 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=2.4219 ps=13.2 w=6.21 l=3.6
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=2.4219 ps=13.2 w=6.21 l=3.6
X5 B.t2 B.t0 B.t1 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=0 ps=0 w=6.21 l=3.6
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=2.4219 ps=13.2 w=6.21 l=3.6
X7 VDD2.t0 VN.t1 VTAIL.t3 w_n2542_n2210# sky130_fd_pr__pfet_01v8 ad=2.4219 pd=13.2 as=2.4219 ps=13.2 w=6.21 l=3.6
R0 B.n362 B.n51 585
R1 B.n364 B.n363 585
R2 B.n365 B.n50 585
R3 B.n367 B.n366 585
R4 B.n368 B.n49 585
R5 B.n370 B.n369 585
R6 B.n371 B.n48 585
R7 B.n373 B.n372 585
R8 B.n374 B.n47 585
R9 B.n376 B.n375 585
R10 B.n377 B.n46 585
R11 B.n379 B.n378 585
R12 B.n380 B.n45 585
R13 B.n382 B.n381 585
R14 B.n383 B.n44 585
R15 B.n385 B.n384 585
R16 B.n386 B.n43 585
R17 B.n388 B.n387 585
R18 B.n389 B.n42 585
R19 B.n391 B.n390 585
R20 B.n392 B.n41 585
R21 B.n394 B.n393 585
R22 B.n395 B.n40 585
R23 B.n397 B.n396 585
R24 B.n398 B.n37 585
R25 B.n401 B.n400 585
R26 B.n402 B.n36 585
R27 B.n404 B.n403 585
R28 B.n405 B.n35 585
R29 B.n407 B.n406 585
R30 B.n408 B.n34 585
R31 B.n410 B.n409 585
R32 B.n411 B.n33 585
R33 B.n413 B.n412 585
R34 B.n415 B.n414 585
R35 B.n416 B.n29 585
R36 B.n418 B.n417 585
R37 B.n419 B.n28 585
R38 B.n421 B.n420 585
R39 B.n422 B.n27 585
R40 B.n424 B.n423 585
R41 B.n425 B.n26 585
R42 B.n427 B.n426 585
R43 B.n428 B.n25 585
R44 B.n430 B.n429 585
R45 B.n431 B.n24 585
R46 B.n433 B.n432 585
R47 B.n434 B.n23 585
R48 B.n436 B.n435 585
R49 B.n437 B.n22 585
R50 B.n439 B.n438 585
R51 B.n440 B.n21 585
R52 B.n442 B.n441 585
R53 B.n443 B.n20 585
R54 B.n445 B.n444 585
R55 B.n446 B.n19 585
R56 B.n448 B.n447 585
R57 B.n449 B.n18 585
R58 B.n451 B.n450 585
R59 B.n361 B.n360 585
R60 B.n359 B.n52 585
R61 B.n358 B.n357 585
R62 B.n356 B.n53 585
R63 B.n355 B.n354 585
R64 B.n353 B.n54 585
R65 B.n352 B.n351 585
R66 B.n350 B.n55 585
R67 B.n349 B.n348 585
R68 B.n347 B.n56 585
R69 B.n346 B.n345 585
R70 B.n344 B.n57 585
R71 B.n343 B.n342 585
R72 B.n341 B.n58 585
R73 B.n340 B.n339 585
R74 B.n338 B.n59 585
R75 B.n337 B.n336 585
R76 B.n335 B.n60 585
R77 B.n334 B.n333 585
R78 B.n332 B.n61 585
R79 B.n331 B.n330 585
R80 B.n329 B.n62 585
R81 B.n328 B.n327 585
R82 B.n326 B.n63 585
R83 B.n325 B.n324 585
R84 B.n323 B.n64 585
R85 B.n322 B.n321 585
R86 B.n320 B.n65 585
R87 B.n319 B.n318 585
R88 B.n317 B.n66 585
R89 B.n316 B.n315 585
R90 B.n314 B.n67 585
R91 B.n313 B.n312 585
R92 B.n311 B.n68 585
R93 B.n310 B.n309 585
R94 B.n308 B.n69 585
R95 B.n307 B.n306 585
R96 B.n305 B.n70 585
R97 B.n304 B.n303 585
R98 B.n302 B.n71 585
R99 B.n301 B.n300 585
R100 B.n299 B.n72 585
R101 B.n298 B.n297 585
R102 B.n296 B.n73 585
R103 B.n295 B.n294 585
R104 B.n293 B.n74 585
R105 B.n292 B.n291 585
R106 B.n290 B.n75 585
R107 B.n289 B.n288 585
R108 B.n287 B.n76 585
R109 B.n286 B.n285 585
R110 B.n284 B.n77 585
R111 B.n283 B.n282 585
R112 B.n281 B.n78 585
R113 B.n280 B.n279 585
R114 B.n278 B.n79 585
R115 B.n277 B.n276 585
R116 B.n275 B.n80 585
R117 B.n274 B.n273 585
R118 B.n272 B.n81 585
R119 B.n271 B.n270 585
R120 B.n269 B.n82 585
R121 B.n268 B.n267 585
R122 B.n178 B.n177 585
R123 B.n179 B.n116 585
R124 B.n181 B.n180 585
R125 B.n182 B.n115 585
R126 B.n184 B.n183 585
R127 B.n185 B.n114 585
R128 B.n187 B.n186 585
R129 B.n188 B.n113 585
R130 B.n190 B.n189 585
R131 B.n191 B.n112 585
R132 B.n193 B.n192 585
R133 B.n194 B.n111 585
R134 B.n196 B.n195 585
R135 B.n197 B.n110 585
R136 B.n199 B.n198 585
R137 B.n200 B.n109 585
R138 B.n202 B.n201 585
R139 B.n203 B.n108 585
R140 B.n205 B.n204 585
R141 B.n206 B.n107 585
R142 B.n208 B.n207 585
R143 B.n209 B.n106 585
R144 B.n211 B.n210 585
R145 B.n212 B.n105 585
R146 B.n214 B.n213 585
R147 B.n216 B.n215 585
R148 B.n217 B.n101 585
R149 B.n219 B.n218 585
R150 B.n220 B.n100 585
R151 B.n222 B.n221 585
R152 B.n223 B.n99 585
R153 B.n225 B.n224 585
R154 B.n226 B.n98 585
R155 B.n228 B.n227 585
R156 B.n230 B.n95 585
R157 B.n232 B.n231 585
R158 B.n233 B.n94 585
R159 B.n235 B.n234 585
R160 B.n236 B.n93 585
R161 B.n238 B.n237 585
R162 B.n239 B.n92 585
R163 B.n241 B.n240 585
R164 B.n242 B.n91 585
R165 B.n244 B.n243 585
R166 B.n245 B.n90 585
R167 B.n247 B.n246 585
R168 B.n248 B.n89 585
R169 B.n250 B.n249 585
R170 B.n251 B.n88 585
R171 B.n253 B.n252 585
R172 B.n254 B.n87 585
R173 B.n256 B.n255 585
R174 B.n257 B.n86 585
R175 B.n259 B.n258 585
R176 B.n260 B.n85 585
R177 B.n262 B.n261 585
R178 B.n263 B.n84 585
R179 B.n265 B.n264 585
R180 B.n266 B.n83 585
R181 B.n176 B.n117 585
R182 B.n175 B.n174 585
R183 B.n173 B.n118 585
R184 B.n172 B.n171 585
R185 B.n170 B.n119 585
R186 B.n169 B.n168 585
R187 B.n167 B.n120 585
R188 B.n166 B.n165 585
R189 B.n164 B.n121 585
R190 B.n163 B.n162 585
R191 B.n161 B.n122 585
R192 B.n160 B.n159 585
R193 B.n158 B.n123 585
R194 B.n157 B.n156 585
R195 B.n155 B.n124 585
R196 B.n154 B.n153 585
R197 B.n152 B.n125 585
R198 B.n151 B.n150 585
R199 B.n149 B.n126 585
R200 B.n148 B.n147 585
R201 B.n146 B.n127 585
R202 B.n145 B.n144 585
R203 B.n143 B.n128 585
R204 B.n142 B.n141 585
R205 B.n140 B.n129 585
R206 B.n139 B.n138 585
R207 B.n137 B.n130 585
R208 B.n136 B.n135 585
R209 B.n134 B.n131 585
R210 B.n133 B.n132 585
R211 B.n2 B.n0 585
R212 B.n497 B.n1 585
R213 B.n496 B.n495 585
R214 B.n494 B.n3 585
R215 B.n493 B.n492 585
R216 B.n491 B.n4 585
R217 B.n490 B.n489 585
R218 B.n488 B.n5 585
R219 B.n487 B.n486 585
R220 B.n485 B.n6 585
R221 B.n484 B.n483 585
R222 B.n482 B.n7 585
R223 B.n481 B.n480 585
R224 B.n479 B.n8 585
R225 B.n478 B.n477 585
R226 B.n476 B.n9 585
R227 B.n475 B.n474 585
R228 B.n473 B.n10 585
R229 B.n472 B.n471 585
R230 B.n470 B.n11 585
R231 B.n469 B.n468 585
R232 B.n467 B.n12 585
R233 B.n466 B.n465 585
R234 B.n464 B.n13 585
R235 B.n463 B.n462 585
R236 B.n461 B.n14 585
R237 B.n460 B.n459 585
R238 B.n458 B.n15 585
R239 B.n457 B.n456 585
R240 B.n455 B.n16 585
R241 B.n454 B.n453 585
R242 B.n452 B.n17 585
R243 B.n499 B.n498 585
R244 B.n178 B.n117 516.524
R245 B.n450 B.n17 516.524
R246 B.n268 B.n83 516.524
R247 B.n360 B.n51 516.524
R248 B.n96 B.t6 250.754
R249 B.n102 B.t9 250.754
R250 B.n30 B.t3 250.754
R251 B.n38 B.t0 250.754
R252 B.n96 B.t8 188.66
R253 B.n38 B.t1 188.66
R254 B.n102 B.t11 188.654
R255 B.n30 B.t4 188.654
R256 B.n174 B.n117 163.367
R257 B.n174 B.n173 163.367
R258 B.n173 B.n172 163.367
R259 B.n172 B.n119 163.367
R260 B.n168 B.n119 163.367
R261 B.n168 B.n167 163.367
R262 B.n167 B.n166 163.367
R263 B.n166 B.n121 163.367
R264 B.n162 B.n121 163.367
R265 B.n162 B.n161 163.367
R266 B.n161 B.n160 163.367
R267 B.n160 B.n123 163.367
R268 B.n156 B.n123 163.367
R269 B.n156 B.n155 163.367
R270 B.n155 B.n154 163.367
R271 B.n154 B.n125 163.367
R272 B.n150 B.n125 163.367
R273 B.n150 B.n149 163.367
R274 B.n149 B.n148 163.367
R275 B.n148 B.n127 163.367
R276 B.n144 B.n127 163.367
R277 B.n144 B.n143 163.367
R278 B.n143 B.n142 163.367
R279 B.n142 B.n129 163.367
R280 B.n138 B.n129 163.367
R281 B.n138 B.n137 163.367
R282 B.n137 B.n136 163.367
R283 B.n136 B.n131 163.367
R284 B.n132 B.n131 163.367
R285 B.n132 B.n2 163.367
R286 B.n498 B.n2 163.367
R287 B.n498 B.n497 163.367
R288 B.n497 B.n496 163.367
R289 B.n496 B.n3 163.367
R290 B.n492 B.n3 163.367
R291 B.n492 B.n491 163.367
R292 B.n491 B.n490 163.367
R293 B.n490 B.n5 163.367
R294 B.n486 B.n5 163.367
R295 B.n486 B.n485 163.367
R296 B.n485 B.n484 163.367
R297 B.n484 B.n7 163.367
R298 B.n480 B.n7 163.367
R299 B.n480 B.n479 163.367
R300 B.n479 B.n478 163.367
R301 B.n478 B.n9 163.367
R302 B.n474 B.n9 163.367
R303 B.n474 B.n473 163.367
R304 B.n473 B.n472 163.367
R305 B.n472 B.n11 163.367
R306 B.n468 B.n11 163.367
R307 B.n468 B.n467 163.367
R308 B.n467 B.n466 163.367
R309 B.n466 B.n13 163.367
R310 B.n462 B.n13 163.367
R311 B.n462 B.n461 163.367
R312 B.n461 B.n460 163.367
R313 B.n460 B.n15 163.367
R314 B.n456 B.n15 163.367
R315 B.n456 B.n455 163.367
R316 B.n455 B.n454 163.367
R317 B.n454 B.n17 163.367
R318 B.n179 B.n178 163.367
R319 B.n180 B.n179 163.367
R320 B.n180 B.n115 163.367
R321 B.n184 B.n115 163.367
R322 B.n185 B.n184 163.367
R323 B.n186 B.n185 163.367
R324 B.n186 B.n113 163.367
R325 B.n190 B.n113 163.367
R326 B.n191 B.n190 163.367
R327 B.n192 B.n191 163.367
R328 B.n192 B.n111 163.367
R329 B.n196 B.n111 163.367
R330 B.n197 B.n196 163.367
R331 B.n198 B.n197 163.367
R332 B.n198 B.n109 163.367
R333 B.n202 B.n109 163.367
R334 B.n203 B.n202 163.367
R335 B.n204 B.n203 163.367
R336 B.n204 B.n107 163.367
R337 B.n208 B.n107 163.367
R338 B.n209 B.n208 163.367
R339 B.n210 B.n209 163.367
R340 B.n210 B.n105 163.367
R341 B.n214 B.n105 163.367
R342 B.n215 B.n214 163.367
R343 B.n215 B.n101 163.367
R344 B.n219 B.n101 163.367
R345 B.n220 B.n219 163.367
R346 B.n221 B.n220 163.367
R347 B.n221 B.n99 163.367
R348 B.n225 B.n99 163.367
R349 B.n226 B.n225 163.367
R350 B.n227 B.n226 163.367
R351 B.n227 B.n95 163.367
R352 B.n232 B.n95 163.367
R353 B.n233 B.n232 163.367
R354 B.n234 B.n233 163.367
R355 B.n234 B.n93 163.367
R356 B.n238 B.n93 163.367
R357 B.n239 B.n238 163.367
R358 B.n240 B.n239 163.367
R359 B.n240 B.n91 163.367
R360 B.n244 B.n91 163.367
R361 B.n245 B.n244 163.367
R362 B.n246 B.n245 163.367
R363 B.n246 B.n89 163.367
R364 B.n250 B.n89 163.367
R365 B.n251 B.n250 163.367
R366 B.n252 B.n251 163.367
R367 B.n252 B.n87 163.367
R368 B.n256 B.n87 163.367
R369 B.n257 B.n256 163.367
R370 B.n258 B.n257 163.367
R371 B.n258 B.n85 163.367
R372 B.n262 B.n85 163.367
R373 B.n263 B.n262 163.367
R374 B.n264 B.n263 163.367
R375 B.n264 B.n83 163.367
R376 B.n269 B.n268 163.367
R377 B.n270 B.n269 163.367
R378 B.n270 B.n81 163.367
R379 B.n274 B.n81 163.367
R380 B.n275 B.n274 163.367
R381 B.n276 B.n275 163.367
R382 B.n276 B.n79 163.367
R383 B.n280 B.n79 163.367
R384 B.n281 B.n280 163.367
R385 B.n282 B.n281 163.367
R386 B.n282 B.n77 163.367
R387 B.n286 B.n77 163.367
R388 B.n287 B.n286 163.367
R389 B.n288 B.n287 163.367
R390 B.n288 B.n75 163.367
R391 B.n292 B.n75 163.367
R392 B.n293 B.n292 163.367
R393 B.n294 B.n293 163.367
R394 B.n294 B.n73 163.367
R395 B.n298 B.n73 163.367
R396 B.n299 B.n298 163.367
R397 B.n300 B.n299 163.367
R398 B.n300 B.n71 163.367
R399 B.n304 B.n71 163.367
R400 B.n305 B.n304 163.367
R401 B.n306 B.n305 163.367
R402 B.n306 B.n69 163.367
R403 B.n310 B.n69 163.367
R404 B.n311 B.n310 163.367
R405 B.n312 B.n311 163.367
R406 B.n312 B.n67 163.367
R407 B.n316 B.n67 163.367
R408 B.n317 B.n316 163.367
R409 B.n318 B.n317 163.367
R410 B.n318 B.n65 163.367
R411 B.n322 B.n65 163.367
R412 B.n323 B.n322 163.367
R413 B.n324 B.n323 163.367
R414 B.n324 B.n63 163.367
R415 B.n328 B.n63 163.367
R416 B.n329 B.n328 163.367
R417 B.n330 B.n329 163.367
R418 B.n330 B.n61 163.367
R419 B.n334 B.n61 163.367
R420 B.n335 B.n334 163.367
R421 B.n336 B.n335 163.367
R422 B.n336 B.n59 163.367
R423 B.n340 B.n59 163.367
R424 B.n341 B.n340 163.367
R425 B.n342 B.n341 163.367
R426 B.n342 B.n57 163.367
R427 B.n346 B.n57 163.367
R428 B.n347 B.n346 163.367
R429 B.n348 B.n347 163.367
R430 B.n348 B.n55 163.367
R431 B.n352 B.n55 163.367
R432 B.n353 B.n352 163.367
R433 B.n354 B.n353 163.367
R434 B.n354 B.n53 163.367
R435 B.n358 B.n53 163.367
R436 B.n359 B.n358 163.367
R437 B.n360 B.n359 163.367
R438 B.n450 B.n449 163.367
R439 B.n449 B.n448 163.367
R440 B.n448 B.n19 163.367
R441 B.n444 B.n19 163.367
R442 B.n444 B.n443 163.367
R443 B.n443 B.n442 163.367
R444 B.n442 B.n21 163.367
R445 B.n438 B.n21 163.367
R446 B.n438 B.n437 163.367
R447 B.n437 B.n436 163.367
R448 B.n436 B.n23 163.367
R449 B.n432 B.n23 163.367
R450 B.n432 B.n431 163.367
R451 B.n431 B.n430 163.367
R452 B.n430 B.n25 163.367
R453 B.n426 B.n25 163.367
R454 B.n426 B.n425 163.367
R455 B.n425 B.n424 163.367
R456 B.n424 B.n27 163.367
R457 B.n420 B.n27 163.367
R458 B.n420 B.n419 163.367
R459 B.n419 B.n418 163.367
R460 B.n418 B.n29 163.367
R461 B.n414 B.n29 163.367
R462 B.n414 B.n413 163.367
R463 B.n413 B.n33 163.367
R464 B.n409 B.n33 163.367
R465 B.n409 B.n408 163.367
R466 B.n408 B.n407 163.367
R467 B.n407 B.n35 163.367
R468 B.n403 B.n35 163.367
R469 B.n403 B.n402 163.367
R470 B.n402 B.n401 163.367
R471 B.n401 B.n37 163.367
R472 B.n396 B.n37 163.367
R473 B.n396 B.n395 163.367
R474 B.n395 B.n394 163.367
R475 B.n394 B.n41 163.367
R476 B.n390 B.n41 163.367
R477 B.n390 B.n389 163.367
R478 B.n389 B.n388 163.367
R479 B.n388 B.n43 163.367
R480 B.n384 B.n43 163.367
R481 B.n384 B.n383 163.367
R482 B.n383 B.n382 163.367
R483 B.n382 B.n45 163.367
R484 B.n378 B.n45 163.367
R485 B.n378 B.n377 163.367
R486 B.n377 B.n376 163.367
R487 B.n376 B.n47 163.367
R488 B.n372 B.n47 163.367
R489 B.n372 B.n371 163.367
R490 B.n371 B.n370 163.367
R491 B.n370 B.n49 163.367
R492 B.n366 B.n49 163.367
R493 B.n366 B.n365 163.367
R494 B.n365 B.n364 163.367
R495 B.n364 B.n51 163.367
R496 B.n97 B.t7 112.442
R497 B.n39 B.t2 112.442
R498 B.n103 B.t10 112.436
R499 B.n31 B.t5 112.436
R500 B.n97 B.n96 76.2187
R501 B.n103 B.n102 76.2187
R502 B.n31 B.n30 76.2187
R503 B.n39 B.n38 76.2187
R504 B.n229 B.n97 59.5399
R505 B.n104 B.n103 59.5399
R506 B.n32 B.n31 59.5399
R507 B.n399 B.n39 59.5399
R508 B.n452 B.n451 33.5615
R509 B.n362 B.n361 33.5615
R510 B.n267 B.n266 33.5615
R511 B.n177 B.n176 33.5615
R512 B B.n499 18.0485
R513 B.n451 B.n18 10.6151
R514 B.n447 B.n18 10.6151
R515 B.n447 B.n446 10.6151
R516 B.n446 B.n445 10.6151
R517 B.n445 B.n20 10.6151
R518 B.n441 B.n20 10.6151
R519 B.n441 B.n440 10.6151
R520 B.n440 B.n439 10.6151
R521 B.n439 B.n22 10.6151
R522 B.n435 B.n22 10.6151
R523 B.n435 B.n434 10.6151
R524 B.n434 B.n433 10.6151
R525 B.n433 B.n24 10.6151
R526 B.n429 B.n24 10.6151
R527 B.n429 B.n428 10.6151
R528 B.n428 B.n427 10.6151
R529 B.n427 B.n26 10.6151
R530 B.n423 B.n26 10.6151
R531 B.n423 B.n422 10.6151
R532 B.n422 B.n421 10.6151
R533 B.n421 B.n28 10.6151
R534 B.n417 B.n28 10.6151
R535 B.n417 B.n416 10.6151
R536 B.n416 B.n415 10.6151
R537 B.n412 B.n411 10.6151
R538 B.n411 B.n410 10.6151
R539 B.n410 B.n34 10.6151
R540 B.n406 B.n34 10.6151
R541 B.n406 B.n405 10.6151
R542 B.n405 B.n404 10.6151
R543 B.n404 B.n36 10.6151
R544 B.n400 B.n36 10.6151
R545 B.n398 B.n397 10.6151
R546 B.n397 B.n40 10.6151
R547 B.n393 B.n40 10.6151
R548 B.n393 B.n392 10.6151
R549 B.n392 B.n391 10.6151
R550 B.n391 B.n42 10.6151
R551 B.n387 B.n42 10.6151
R552 B.n387 B.n386 10.6151
R553 B.n386 B.n385 10.6151
R554 B.n385 B.n44 10.6151
R555 B.n381 B.n44 10.6151
R556 B.n381 B.n380 10.6151
R557 B.n380 B.n379 10.6151
R558 B.n379 B.n46 10.6151
R559 B.n375 B.n46 10.6151
R560 B.n375 B.n374 10.6151
R561 B.n374 B.n373 10.6151
R562 B.n373 B.n48 10.6151
R563 B.n369 B.n48 10.6151
R564 B.n369 B.n368 10.6151
R565 B.n368 B.n367 10.6151
R566 B.n367 B.n50 10.6151
R567 B.n363 B.n50 10.6151
R568 B.n363 B.n362 10.6151
R569 B.n267 B.n82 10.6151
R570 B.n271 B.n82 10.6151
R571 B.n272 B.n271 10.6151
R572 B.n273 B.n272 10.6151
R573 B.n273 B.n80 10.6151
R574 B.n277 B.n80 10.6151
R575 B.n278 B.n277 10.6151
R576 B.n279 B.n278 10.6151
R577 B.n279 B.n78 10.6151
R578 B.n283 B.n78 10.6151
R579 B.n284 B.n283 10.6151
R580 B.n285 B.n284 10.6151
R581 B.n285 B.n76 10.6151
R582 B.n289 B.n76 10.6151
R583 B.n290 B.n289 10.6151
R584 B.n291 B.n290 10.6151
R585 B.n291 B.n74 10.6151
R586 B.n295 B.n74 10.6151
R587 B.n296 B.n295 10.6151
R588 B.n297 B.n296 10.6151
R589 B.n297 B.n72 10.6151
R590 B.n301 B.n72 10.6151
R591 B.n302 B.n301 10.6151
R592 B.n303 B.n302 10.6151
R593 B.n303 B.n70 10.6151
R594 B.n307 B.n70 10.6151
R595 B.n308 B.n307 10.6151
R596 B.n309 B.n308 10.6151
R597 B.n309 B.n68 10.6151
R598 B.n313 B.n68 10.6151
R599 B.n314 B.n313 10.6151
R600 B.n315 B.n314 10.6151
R601 B.n315 B.n66 10.6151
R602 B.n319 B.n66 10.6151
R603 B.n320 B.n319 10.6151
R604 B.n321 B.n320 10.6151
R605 B.n321 B.n64 10.6151
R606 B.n325 B.n64 10.6151
R607 B.n326 B.n325 10.6151
R608 B.n327 B.n326 10.6151
R609 B.n327 B.n62 10.6151
R610 B.n331 B.n62 10.6151
R611 B.n332 B.n331 10.6151
R612 B.n333 B.n332 10.6151
R613 B.n333 B.n60 10.6151
R614 B.n337 B.n60 10.6151
R615 B.n338 B.n337 10.6151
R616 B.n339 B.n338 10.6151
R617 B.n339 B.n58 10.6151
R618 B.n343 B.n58 10.6151
R619 B.n344 B.n343 10.6151
R620 B.n345 B.n344 10.6151
R621 B.n345 B.n56 10.6151
R622 B.n349 B.n56 10.6151
R623 B.n350 B.n349 10.6151
R624 B.n351 B.n350 10.6151
R625 B.n351 B.n54 10.6151
R626 B.n355 B.n54 10.6151
R627 B.n356 B.n355 10.6151
R628 B.n357 B.n356 10.6151
R629 B.n357 B.n52 10.6151
R630 B.n361 B.n52 10.6151
R631 B.n177 B.n116 10.6151
R632 B.n181 B.n116 10.6151
R633 B.n182 B.n181 10.6151
R634 B.n183 B.n182 10.6151
R635 B.n183 B.n114 10.6151
R636 B.n187 B.n114 10.6151
R637 B.n188 B.n187 10.6151
R638 B.n189 B.n188 10.6151
R639 B.n189 B.n112 10.6151
R640 B.n193 B.n112 10.6151
R641 B.n194 B.n193 10.6151
R642 B.n195 B.n194 10.6151
R643 B.n195 B.n110 10.6151
R644 B.n199 B.n110 10.6151
R645 B.n200 B.n199 10.6151
R646 B.n201 B.n200 10.6151
R647 B.n201 B.n108 10.6151
R648 B.n205 B.n108 10.6151
R649 B.n206 B.n205 10.6151
R650 B.n207 B.n206 10.6151
R651 B.n207 B.n106 10.6151
R652 B.n211 B.n106 10.6151
R653 B.n212 B.n211 10.6151
R654 B.n213 B.n212 10.6151
R655 B.n217 B.n216 10.6151
R656 B.n218 B.n217 10.6151
R657 B.n218 B.n100 10.6151
R658 B.n222 B.n100 10.6151
R659 B.n223 B.n222 10.6151
R660 B.n224 B.n223 10.6151
R661 B.n224 B.n98 10.6151
R662 B.n228 B.n98 10.6151
R663 B.n231 B.n230 10.6151
R664 B.n231 B.n94 10.6151
R665 B.n235 B.n94 10.6151
R666 B.n236 B.n235 10.6151
R667 B.n237 B.n236 10.6151
R668 B.n237 B.n92 10.6151
R669 B.n241 B.n92 10.6151
R670 B.n242 B.n241 10.6151
R671 B.n243 B.n242 10.6151
R672 B.n243 B.n90 10.6151
R673 B.n247 B.n90 10.6151
R674 B.n248 B.n247 10.6151
R675 B.n249 B.n248 10.6151
R676 B.n249 B.n88 10.6151
R677 B.n253 B.n88 10.6151
R678 B.n254 B.n253 10.6151
R679 B.n255 B.n254 10.6151
R680 B.n255 B.n86 10.6151
R681 B.n259 B.n86 10.6151
R682 B.n260 B.n259 10.6151
R683 B.n261 B.n260 10.6151
R684 B.n261 B.n84 10.6151
R685 B.n265 B.n84 10.6151
R686 B.n266 B.n265 10.6151
R687 B.n176 B.n175 10.6151
R688 B.n175 B.n118 10.6151
R689 B.n171 B.n118 10.6151
R690 B.n171 B.n170 10.6151
R691 B.n170 B.n169 10.6151
R692 B.n169 B.n120 10.6151
R693 B.n165 B.n120 10.6151
R694 B.n165 B.n164 10.6151
R695 B.n164 B.n163 10.6151
R696 B.n163 B.n122 10.6151
R697 B.n159 B.n122 10.6151
R698 B.n159 B.n158 10.6151
R699 B.n158 B.n157 10.6151
R700 B.n157 B.n124 10.6151
R701 B.n153 B.n124 10.6151
R702 B.n153 B.n152 10.6151
R703 B.n152 B.n151 10.6151
R704 B.n151 B.n126 10.6151
R705 B.n147 B.n126 10.6151
R706 B.n147 B.n146 10.6151
R707 B.n146 B.n145 10.6151
R708 B.n145 B.n128 10.6151
R709 B.n141 B.n128 10.6151
R710 B.n141 B.n140 10.6151
R711 B.n140 B.n139 10.6151
R712 B.n139 B.n130 10.6151
R713 B.n135 B.n130 10.6151
R714 B.n135 B.n134 10.6151
R715 B.n134 B.n133 10.6151
R716 B.n133 B.n0 10.6151
R717 B.n495 B.n1 10.6151
R718 B.n495 B.n494 10.6151
R719 B.n494 B.n493 10.6151
R720 B.n493 B.n4 10.6151
R721 B.n489 B.n4 10.6151
R722 B.n489 B.n488 10.6151
R723 B.n488 B.n487 10.6151
R724 B.n487 B.n6 10.6151
R725 B.n483 B.n6 10.6151
R726 B.n483 B.n482 10.6151
R727 B.n482 B.n481 10.6151
R728 B.n481 B.n8 10.6151
R729 B.n477 B.n8 10.6151
R730 B.n477 B.n476 10.6151
R731 B.n476 B.n475 10.6151
R732 B.n475 B.n10 10.6151
R733 B.n471 B.n10 10.6151
R734 B.n471 B.n470 10.6151
R735 B.n470 B.n469 10.6151
R736 B.n469 B.n12 10.6151
R737 B.n465 B.n12 10.6151
R738 B.n465 B.n464 10.6151
R739 B.n464 B.n463 10.6151
R740 B.n463 B.n14 10.6151
R741 B.n459 B.n14 10.6151
R742 B.n459 B.n458 10.6151
R743 B.n458 B.n457 10.6151
R744 B.n457 B.n16 10.6151
R745 B.n453 B.n16 10.6151
R746 B.n453 B.n452 10.6151
R747 B.n412 B.n32 6.5566
R748 B.n400 B.n399 6.5566
R749 B.n216 B.n104 6.5566
R750 B.n229 B.n228 6.5566
R751 B.n415 B.n32 4.05904
R752 B.n399 B.n398 4.05904
R753 B.n213 B.n104 4.05904
R754 B.n230 B.n229 4.05904
R755 B.n499 B.n0 2.81026
R756 B.n499 B.n1 2.81026
R757 VN VN.t0 123.189
R758 VN VN.t1 80.8866
R759 VTAIL.n1 VTAIL.t2 82.2531
R760 VTAIL.n3 VTAIL.t3 82.2521
R761 VTAIL.n0 VTAIL.t0 82.2521
R762 VTAIL.n2 VTAIL.t1 82.2521
R763 VTAIL.n1 VTAIL.n0 24.4962
R764 VTAIL.n3 VTAIL.n2 21.1083
R765 VTAIL.n2 VTAIL.n1 2.16429
R766 VTAIL VTAIL.n0 1.3755
R767 VTAIL VTAIL.n3 0.789293
R768 VDD2.n0 VDD2.t0 134.72
R769 VDD2.n0 VDD2.t1 98.9308
R770 VDD2 VDD2.n0 0.905672
R771 VP.n0 VP.t1 123.282
R772 VP.n0 VP.t0 80.3607
R773 VP VP.n0 0.52637
R774 VDD1 VDD1.t1 136.091
R775 VDD1 VDD1.t0 99.836
C0 VP B 1.68508f
C1 VDD1 VDD2 0.782139f
C2 VTAIL VDD2 3.87031f
C3 VN VDD2 1.62893f
C4 VTAIL VDD1 3.8112f
C5 VDD2 w_n2542_n2210# 1.53563f
C6 VN VDD1 0.148581f
C7 VDD1 w_n2542_n2210# 1.49741f
C8 VTAIL VN 1.73913f
C9 VTAIL w_n2542_n2210# 1.98357f
C10 VN w_n2542_n2210# 3.48971f
C11 VDD2 B 1.41047f
C12 VDD1 B 1.37145f
C13 VTAIL B 2.64228f
C14 VP VDD2 0.374692f
C15 VN B 1.14518f
C16 VP VDD1 1.85371f
C17 w_n2542_n2210# B 8.277889f
C18 VTAIL VP 1.75334f
C19 VN VP 4.84985f
C20 VP w_n2542_n2210# 3.81567f
C21 VDD2 VSUBS 0.764264f
C22 VDD1 VSUBS 3.160507f
C23 VTAIL VSUBS 0.580045f
C24 VN VSUBS 5.79374f
C25 VP VSUBS 1.629788f
C26 B VSUBS 4.153847f
C27 w_n2542_n2210# VSUBS 70.0677f
C28 VDD1.t0 VSUBS 0.651979f
C29 VDD1.t1 VSUBS 0.933407f
C30 VP.t1 VSUBS 2.96332f
C31 VP.t0 VSUBS 2.25619f
C32 VP.n0 VSUBS 3.26262f
C33 VDD2.t0 VSUBS 0.94876f
C34 VDD2.t1 VSUBS 0.675806f
C35 VDD2.n0 VSUBS 2.14848f
C36 VTAIL.t0 VSUBS 0.917675f
C37 VTAIL.n0 VSUBS 1.72238f
C38 VTAIL.t2 VSUBS 0.917679f
C39 VTAIL.n1 VSUBS 1.77907f
C40 VTAIL.t1 VSUBS 0.917672f
C41 VTAIL.n2 VSUBS 1.53558f
C42 VTAIL.t3 VSUBS 0.917675f
C43 VTAIL.n3 VSUBS 1.43675f
C44 VN.t1 VSUBS 2.17099f
C45 VN.t0 VSUBS 2.84629f
C46 B.n0 VSUBS 0.004685f
C47 B.n1 VSUBS 0.004685f
C48 B.n2 VSUBS 0.007409f
C49 B.n3 VSUBS 0.007409f
C50 B.n4 VSUBS 0.007409f
C51 B.n5 VSUBS 0.007409f
C52 B.n6 VSUBS 0.007409f
C53 B.n7 VSUBS 0.007409f
C54 B.n8 VSUBS 0.007409f
C55 B.n9 VSUBS 0.007409f
C56 B.n10 VSUBS 0.007409f
C57 B.n11 VSUBS 0.007409f
C58 B.n12 VSUBS 0.007409f
C59 B.n13 VSUBS 0.007409f
C60 B.n14 VSUBS 0.007409f
C61 B.n15 VSUBS 0.007409f
C62 B.n16 VSUBS 0.007409f
C63 B.n17 VSUBS 0.016997f
C64 B.n18 VSUBS 0.007409f
C65 B.n19 VSUBS 0.007409f
C66 B.n20 VSUBS 0.007409f
C67 B.n21 VSUBS 0.007409f
C68 B.n22 VSUBS 0.007409f
C69 B.n23 VSUBS 0.007409f
C70 B.n24 VSUBS 0.007409f
C71 B.n25 VSUBS 0.007409f
C72 B.n26 VSUBS 0.007409f
C73 B.n27 VSUBS 0.007409f
C74 B.n28 VSUBS 0.007409f
C75 B.n29 VSUBS 0.007409f
C76 B.t5 VSUBS 0.193327f
C77 B.t4 VSUBS 0.221134f
C78 B.t3 VSUBS 1.13377f
C79 B.n30 VSUBS 0.135721f
C80 B.n31 VSUBS 0.079395f
C81 B.n32 VSUBS 0.017166f
C82 B.n33 VSUBS 0.007409f
C83 B.n34 VSUBS 0.007409f
C84 B.n35 VSUBS 0.007409f
C85 B.n36 VSUBS 0.007409f
C86 B.n37 VSUBS 0.007409f
C87 B.t2 VSUBS 0.193326f
C88 B.t1 VSUBS 0.221133f
C89 B.t0 VSUBS 1.13377f
C90 B.n38 VSUBS 0.135722f
C91 B.n39 VSUBS 0.079396f
C92 B.n40 VSUBS 0.007409f
C93 B.n41 VSUBS 0.007409f
C94 B.n42 VSUBS 0.007409f
C95 B.n43 VSUBS 0.007409f
C96 B.n44 VSUBS 0.007409f
C97 B.n45 VSUBS 0.007409f
C98 B.n46 VSUBS 0.007409f
C99 B.n47 VSUBS 0.007409f
C100 B.n48 VSUBS 0.007409f
C101 B.n49 VSUBS 0.007409f
C102 B.n50 VSUBS 0.007409f
C103 B.n51 VSUBS 0.018306f
C104 B.n52 VSUBS 0.007409f
C105 B.n53 VSUBS 0.007409f
C106 B.n54 VSUBS 0.007409f
C107 B.n55 VSUBS 0.007409f
C108 B.n56 VSUBS 0.007409f
C109 B.n57 VSUBS 0.007409f
C110 B.n58 VSUBS 0.007409f
C111 B.n59 VSUBS 0.007409f
C112 B.n60 VSUBS 0.007409f
C113 B.n61 VSUBS 0.007409f
C114 B.n62 VSUBS 0.007409f
C115 B.n63 VSUBS 0.007409f
C116 B.n64 VSUBS 0.007409f
C117 B.n65 VSUBS 0.007409f
C118 B.n66 VSUBS 0.007409f
C119 B.n67 VSUBS 0.007409f
C120 B.n68 VSUBS 0.007409f
C121 B.n69 VSUBS 0.007409f
C122 B.n70 VSUBS 0.007409f
C123 B.n71 VSUBS 0.007409f
C124 B.n72 VSUBS 0.007409f
C125 B.n73 VSUBS 0.007409f
C126 B.n74 VSUBS 0.007409f
C127 B.n75 VSUBS 0.007409f
C128 B.n76 VSUBS 0.007409f
C129 B.n77 VSUBS 0.007409f
C130 B.n78 VSUBS 0.007409f
C131 B.n79 VSUBS 0.007409f
C132 B.n80 VSUBS 0.007409f
C133 B.n81 VSUBS 0.007409f
C134 B.n82 VSUBS 0.007409f
C135 B.n83 VSUBS 0.018306f
C136 B.n84 VSUBS 0.007409f
C137 B.n85 VSUBS 0.007409f
C138 B.n86 VSUBS 0.007409f
C139 B.n87 VSUBS 0.007409f
C140 B.n88 VSUBS 0.007409f
C141 B.n89 VSUBS 0.007409f
C142 B.n90 VSUBS 0.007409f
C143 B.n91 VSUBS 0.007409f
C144 B.n92 VSUBS 0.007409f
C145 B.n93 VSUBS 0.007409f
C146 B.n94 VSUBS 0.007409f
C147 B.n95 VSUBS 0.007409f
C148 B.t7 VSUBS 0.193326f
C149 B.t8 VSUBS 0.221133f
C150 B.t6 VSUBS 1.13377f
C151 B.n96 VSUBS 0.135722f
C152 B.n97 VSUBS 0.079396f
C153 B.n98 VSUBS 0.007409f
C154 B.n99 VSUBS 0.007409f
C155 B.n100 VSUBS 0.007409f
C156 B.n101 VSUBS 0.007409f
C157 B.t10 VSUBS 0.193327f
C158 B.t11 VSUBS 0.221134f
C159 B.t9 VSUBS 1.13377f
C160 B.n102 VSUBS 0.135721f
C161 B.n103 VSUBS 0.079395f
C162 B.n104 VSUBS 0.017166f
C163 B.n105 VSUBS 0.007409f
C164 B.n106 VSUBS 0.007409f
C165 B.n107 VSUBS 0.007409f
C166 B.n108 VSUBS 0.007409f
C167 B.n109 VSUBS 0.007409f
C168 B.n110 VSUBS 0.007409f
C169 B.n111 VSUBS 0.007409f
C170 B.n112 VSUBS 0.007409f
C171 B.n113 VSUBS 0.007409f
C172 B.n114 VSUBS 0.007409f
C173 B.n115 VSUBS 0.007409f
C174 B.n116 VSUBS 0.007409f
C175 B.n117 VSUBS 0.016997f
C176 B.n118 VSUBS 0.007409f
C177 B.n119 VSUBS 0.007409f
C178 B.n120 VSUBS 0.007409f
C179 B.n121 VSUBS 0.007409f
C180 B.n122 VSUBS 0.007409f
C181 B.n123 VSUBS 0.007409f
C182 B.n124 VSUBS 0.007409f
C183 B.n125 VSUBS 0.007409f
C184 B.n126 VSUBS 0.007409f
C185 B.n127 VSUBS 0.007409f
C186 B.n128 VSUBS 0.007409f
C187 B.n129 VSUBS 0.007409f
C188 B.n130 VSUBS 0.007409f
C189 B.n131 VSUBS 0.007409f
C190 B.n132 VSUBS 0.007409f
C191 B.n133 VSUBS 0.007409f
C192 B.n134 VSUBS 0.007409f
C193 B.n135 VSUBS 0.007409f
C194 B.n136 VSUBS 0.007409f
C195 B.n137 VSUBS 0.007409f
C196 B.n138 VSUBS 0.007409f
C197 B.n139 VSUBS 0.007409f
C198 B.n140 VSUBS 0.007409f
C199 B.n141 VSUBS 0.007409f
C200 B.n142 VSUBS 0.007409f
C201 B.n143 VSUBS 0.007409f
C202 B.n144 VSUBS 0.007409f
C203 B.n145 VSUBS 0.007409f
C204 B.n146 VSUBS 0.007409f
C205 B.n147 VSUBS 0.007409f
C206 B.n148 VSUBS 0.007409f
C207 B.n149 VSUBS 0.007409f
C208 B.n150 VSUBS 0.007409f
C209 B.n151 VSUBS 0.007409f
C210 B.n152 VSUBS 0.007409f
C211 B.n153 VSUBS 0.007409f
C212 B.n154 VSUBS 0.007409f
C213 B.n155 VSUBS 0.007409f
C214 B.n156 VSUBS 0.007409f
C215 B.n157 VSUBS 0.007409f
C216 B.n158 VSUBS 0.007409f
C217 B.n159 VSUBS 0.007409f
C218 B.n160 VSUBS 0.007409f
C219 B.n161 VSUBS 0.007409f
C220 B.n162 VSUBS 0.007409f
C221 B.n163 VSUBS 0.007409f
C222 B.n164 VSUBS 0.007409f
C223 B.n165 VSUBS 0.007409f
C224 B.n166 VSUBS 0.007409f
C225 B.n167 VSUBS 0.007409f
C226 B.n168 VSUBS 0.007409f
C227 B.n169 VSUBS 0.007409f
C228 B.n170 VSUBS 0.007409f
C229 B.n171 VSUBS 0.007409f
C230 B.n172 VSUBS 0.007409f
C231 B.n173 VSUBS 0.007409f
C232 B.n174 VSUBS 0.007409f
C233 B.n175 VSUBS 0.007409f
C234 B.n176 VSUBS 0.016997f
C235 B.n177 VSUBS 0.018306f
C236 B.n178 VSUBS 0.018306f
C237 B.n179 VSUBS 0.007409f
C238 B.n180 VSUBS 0.007409f
C239 B.n181 VSUBS 0.007409f
C240 B.n182 VSUBS 0.007409f
C241 B.n183 VSUBS 0.007409f
C242 B.n184 VSUBS 0.007409f
C243 B.n185 VSUBS 0.007409f
C244 B.n186 VSUBS 0.007409f
C245 B.n187 VSUBS 0.007409f
C246 B.n188 VSUBS 0.007409f
C247 B.n189 VSUBS 0.007409f
C248 B.n190 VSUBS 0.007409f
C249 B.n191 VSUBS 0.007409f
C250 B.n192 VSUBS 0.007409f
C251 B.n193 VSUBS 0.007409f
C252 B.n194 VSUBS 0.007409f
C253 B.n195 VSUBS 0.007409f
C254 B.n196 VSUBS 0.007409f
C255 B.n197 VSUBS 0.007409f
C256 B.n198 VSUBS 0.007409f
C257 B.n199 VSUBS 0.007409f
C258 B.n200 VSUBS 0.007409f
C259 B.n201 VSUBS 0.007409f
C260 B.n202 VSUBS 0.007409f
C261 B.n203 VSUBS 0.007409f
C262 B.n204 VSUBS 0.007409f
C263 B.n205 VSUBS 0.007409f
C264 B.n206 VSUBS 0.007409f
C265 B.n207 VSUBS 0.007409f
C266 B.n208 VSUBS 0.007409f
C267 B.n209 VSUBS 0.007409f
C268 B.n210 VSUBS 0.007409f
C269 B.n211 VSUBS 0.007409f
C270 B.n212 VSUBS 0.007409f
C271 B.n213 VSUBS 0.005121f
C272 B.n214 VSUBS 0.007409f
C273 B.n215 VSUBS 0.007409f
C274 B.n216 VSUBS 0.005993f
C275 B.n217 VSUBS 0.007409f
C276 B.n218 VSUBS 0.007409f
C277 B.n219 VSUBS 0.007409f
C278 B.n220 VSUBS 0.007409f
C279 B.n221 VSUBS 0.007409f
C280 B.n222 VSUBS 0.007409f
C281 B.n223 VSUBS 0.007409f
C282 B.n224 VSUBS 0.007409f
C283 B.n225 VSUBS 0.007409f
C284 B.n226 VSUBS 0.007409f
C285 B.n227 VSUBS 0.007409f
C286 B.n228 VSUBS 0.005993f
C287 B.n229 VSUBS 0.017166f
C288 B.n230 VSUBS 0.005121f
C289 B.n231 VSUBS 0.007409f
C290 B.n232 VSUBS 0.007409f
C291 B.n233 VSUBS 0.007409f
C292 B.n234 VSUBS 0.007409f
C293 B.n235 VSUBS 0.007409f
C294 B.n236 VSUBS 0.007409f
C295 B.n237 VSUBS 0.007409f
C296 B.n238 VSUBS 0.007409f
C297 B.n239 VSUBS 0.007409f
C298 B.n240 VSUBS 0.007409f
C299 B.n241 VSUBS 0.007409f
C300 B.n242 VSUBS 0.007409f
C301 B.n243 VSUBS 0.007409f
C302 B.n244 VSUBS 0.007409f
C303 B.n245 VSUBS 0.007409f
C304 B.n246 VSUBS 0.007409f
C305 B.n247 VSUBS 0.007409f
C306 B.n248 VSUBS 0.007409f
C307 B.n249 VSUBS 0.007409f
C308 B.n250 VSUBS 0.007409f
C309 B.n251 VSUBS 0.007409f
C310 B.n252 VSUBS 0.007409f
C311 B.n253 VSUBS 0.007409f
C312 B.n254 VSUBS 0.007409f
C313 B.n255 VSUBS 0.007409f
C314 B.n256 VSUBS 0.007409f
C315 B.n257 VSUBS 0.007409f
C316 B.n258 VSUBS 0.007409f
C317 B.n259 VSUBS 0.007409f
C318 B.n260 VSUBS 0.007409f
C319 B.n261 VSUBS 0.007409f
C320 B.n262 VSUBS 0.007409f
C321 B.n263 VSUBS 0.007409f
C322 B.n264 VSUBS 0.007409f
C323 B.n265 VSUBS 0.007409f
C324 B.n266 VSUBS 0.018306f
C325 B.n267 VSUBS 0.016997f
C326 B.n268 VSUBS 0.016997f
C327 B.n269 VSUBS 0.007409f
C328 B.n270 VSUBS 0.007409f
C329 B.n271 VSUBS 0.007409f
C330 B.n272 VSUBS 0.007409f
C331 B.n273 VSUBS 0.007409f
C332 B.n274 VSUBS 0.007409f
C333 B.n275 VSUBS 0.007409f
C334 B.n276 VSUBS 0.007409f
C335 B.n277 VSUBS 0.007409f
C336 B.n278 VSUBS 0.007409f
C337 B.n279 VSUBS 0.007409f
C338 B.n280 VSUBS 0.007409f
C339 B.n281 VSUBS 0.007409f
C340 B.n282 VSUBS 0.007409f
C341 B.n283 VSUBS 0.007409f
C342 B.n284 VSUBS 0.007409f
C343 B.n285 VSUBS 0.007409f
C344 B.n286 VSUBS 0.007409f
C345 B.n287 VSUBS 0.007409f
C346 B.n288 VSUBS 0.007409f
C347 B.n289 VSUBS 0.007409f
C348 B.n290 VSUBS 0.007409f
C349 B.n291 VSUBS 0.007409f
C350 B.n292 VSUBS 0.007409f
C351 B.n293 VSUBS 0.007409f
C352 B.n294 VSUBS 0.007409f
C353 B.n295 VSUBS 0.007409f
C354 B.n296 VSUBS 0.007409f
C355 B.n297 VSUBS 0.007409f
C356 B.n298 VSUBS 0.007409f
C357 B.n299 VSUBS 0.007409f
C358 B.n300 VSUBS 0.007409f
C359 B.n301 VSUBS 0.007409f
C360 B.n302 VSUBS 0.007409f
C361 B.n303 VSUBS 0.007409f
C362 B.n304 VSUBS 0.007409f
C363 B.n305 VSUBS 0.007409f
C364 B.n306 VSUBS 0.007409f
C365 B.n307 VSUBS 0.007409f
C366 B.n308 VSUBS 0.007409f
C367 B.n309 VSUBS 0.007409f
C368 B.n310 VSUBS 0.007409f
C369 B.n311 VSUBS 0.007409f
C370 B.n312 VSUBS 0.007409f
C371 B.n313 VSUBS 0.007409f
C372 B.n314 VSUBS 0.007409f
C373 B.n315 VSUBS 0.007409f
C374 B.n316 VSUBS 0.007409f
C375 B.n317 VSUBS 0.007409f
C376 B.n318 VSUBS 0.007409f
C377 B.n319 VSUBS 0.007409f
C378 B.n320 VSUBS 0.007409f
C379 B.n321 VSUBS 0.007409f
C380 B.n322 VSUBS 0.007409f
C381 B.n323 VSUBS 0.007409f
C382 B.n324 VSUBS 0.007409f
C383 B.n325 VSUBS 0.007409f
C384 B.n326 VSUBS 0.007409f
C385 B.n327 VSUBS 0.007409f
C386 B.n328 VSUBS 0.007409f
C387 B.n329 VSUBS 0.007409f
C388 B.n330 VSUBS 0.007409f
C389 B.n331 VSUBS 0.007409f
C390 B.n332 VSUBS 0.007409f
C391 B.n333 VSUBS 0.007409f
C392 B.n334 VSUBS 0.007409f
C393 B.n335 VSUBS 0.007409f
C394 B.n336 VSUBS 0.007409f
C395 B.n337 VSUBS 0.007409f
C396 B.n338 VSUBS 0.007409f
C397 B.n339 VSUBS 0.007409f
C398 B.n340 VSUBS 0.007409f
C399 B.n341 VSUBS 0.007409f
C400 B.n342 VSUBS 0.007409f
C401 B.n343 VSUBS 0.007409f
C402 B.n344 VSUBS 0.007409f
C403 B.n345 VSUBS 0.007409f
C404 B.n346 VSUBS 0.007409f
C405 B.n347 VSUBS 0.007409f
C406 B.n348 VSUBS 0.007409f
C407 B.n349 VSUBS 0.007409f
C408 B.n350 VSUBS 0.007409f
C409 B.n351 VSUBS 0.007409f
C410 B.n352 VSUBS 0.007409f
C411 B.n353 VSUBS 0.007409f
C412 B.n354 VSUBS 0.007409f
C413 B.n355 VSUBS 0.007409f
C414 B.n356 VSUBS 0.007409f
C415 B.n357 VSUBS 0.007409f
C416 B.n358 VSUBS 0.007409f
C417 B.n359 VSUBS 0.007409f
C418 B.n360 VSUBS 0.016997f
C419 B.n361 VSUBS 0.017848f
C420 B.n362 VSUBS 0.017454f
C421 B.n363 VSUBS 0.007409f
C422 B.n364 VSUBS 0.007409f
C423 B.n365 VSUBS 0.007409f
C424 B.n366 VSUBS 0.007409f
C425 B.n367 VSUBS 0.007409f
C426 B.n368 VSUBS 0.007409f
C427 B.n369 VSUBS 0.007409f
C428 B.n370 VSUBS 0.007409f
C429 B.n371 VSUBS 0.007409f
C430 B.n372 VSUBS 0.007409f
C431 B.n373 VSUBS 0.007409f
C432 B.n374 VSUBS 0.007409f
C433 B.n375 VSUBS 0.007409f
C434 B.n376 VSUBS 0.007409f
C435 B.n377 VSUBS 0.007409f
C436 B.n378 VSUBS 0.007409f
C437 B.n379 VSUBS 0.007409f
C438 B.n380 VSUBS 0.007409f
C439 B.n381 VSUBS 0.007409f
C440 B.n382 VSUBS 0.007409f
C441 B.n383 VSUBS 0.007409f
C442 B.n384 VSUBS 0.007409f
C443 B.n385 VSUBS 0.007409f
C444 B.n386 VSUBS 0.007409f
C445 B.n387 VSUBS 0.007409f
C446 B.n388 VSUBS 0.007409f
C447 B.n389 VSUBS 0.007409f
C448 B.n390 VSUBS 0.007409f
C449 B.n391 VSUBS 0.007409f
C450 B.n392 VSUBS 0.007409f
C451 B.n393 VSUBS 0.007409f
C452 B.n394 VSUBS 0.007409f
C453 B.n395 VSUBS 0.007409f
C454 B.n396 VSUBS 0.007409f
C455 B.n397 VSUBS 0.007409f
C456 B.n398 VSUBS 0.005121f
C457 B.n399 VSUBS 0.017166f
C458 B.n400 VSUBS 0.005993f
C459 B.n401 VSUBS 0.007409f
C460 B.n402 VSUBS 0.007409f
C461 B.n403 VSUBS 0.007409f
C462 B.n404 VSUBS 0.007409f
C463 B.n405 VSUBS 0.007409f
C464 B.n406 VSUBS 0.007409f
C465 B.n407 VSUBS 0.007409f
C466 B.n408 VSUBS 0.007409f
C467 B.n409 VSUBS 0.007409f
C468 B.n410 VSUBS 0.007409f
C469 B.n411 VSUBS 0.007409f
C470 B.n412 VSUBS 0.005993f
C471 B.n413 VSUBS 0.007409f
C472 B.n414 VSUBS 0.007409f
C473 B.n415 VSUBS 0.005121f
C474 B.n416 VSUBS 0.007409f
C475 B.n417 VSUBS 0.007409f
C476 B.n418 VSUBS 0.007409f
C477 B.n419 VSUBS 0.007409f
C478 B.n420 VSUBS 0.007409f
C479 B.n421 VSUBS 0.007409f
C480 B.n422 VSUBS 0.007409f
C481 B.n423 VSUBS 0.007409f
C482 B.n424 VSUBS 0.007409f
C483 B.n425 VSUBS 0.007409f
C484 B.n426 VSUBS 0.007409f
C485 B.n427 VSUBS 0.007409f
C486 B.n428 VSUBS 0.007409f
C487 B.n429 VSUBS 0.007409f
C488 B.n430 VSUBS 0.007409f
C489 B.n431 VSUBS 0.007409f
C490 B.n432 VSUBS 0.007409f
C491 B.n433 VSUBS 0.007409f
C492 B.n434 VSUBS 0.007409f
C493 B.n435 VSUBS 0.007409f
C494 B.n436 VSUBS 0.007409f
C495 B.n437 VSUBS 0.007409f
C496 B.n438 VSUBS 0.007409f
C497 B.n439 VSUBS 0.007409f
C498 B.n440 VSUBS 0.007409f
C499 B.n441 VSUBS 0.007409f
C500 B.n442 VSUBS 0.007409f
C501 B.n443 VSUBS 0.007409f
C502 B.n444 VSUBS 0.007409f
C503 B.n445 VSUBS 0.007409f
C504 B.n446 VSUBS 0.007409f
C505 B.n447 VSUBS 0.007409f
C506 B.n448 VSUBS 0.007409f
C507 B.n449 VSUBS 0.007409f
C508 B.n450 VSUBS 0.018306f
C509 B.n451 VSUBS 0.018306f
C510 B.n452 VSUBS 0.016997f
C511 B.n453 VSUBS 0.007409f
C512 B.n454 VSUBS 0.007409f
C513 B.n455 VSUBS 0.007409f
C514 B.n456 VSUBS 0.007409f
C515 B.n457 VSUBS 0.007409f
C516 B.n458 VSUBS 0.007409f
C517 B.n459 VSUBS 0.007409f
C518 B.n460 VSUBS 0.007409f
C519 B.n461 VSUBS 0.007409f
C520 B.n462 VSUBS 0.007409f
C521 B.n463 VSUBS 0.007409f
C522 B.n464 VSUBS 0.007409f
C523 B.n465 VSUBS 0.007409f
C524 B.n466 VSUBS 0.007409f
C525 B.n467 VSUBS 0.007409f
C526 B.n468 VSUBS 0.007409f
C527 B.n469 VSUBS 0.007409f
C528 B.n470 VSUBS 0.007409f
C529 B.n471 VSUBS 0.007409f
C530 B.n472 VSUBS 0.007409f
C531 B.n473 VSUBS 0.007409f
C532 B.n474 VSUBS 0.007409f
C533 B.n475 VSUBS 0.007409f
C534 B.n476 VSUBS 0.007409f
C535 B.n477 VSUBS 0.007409f
C536 B.n478 VSUBS 0.007409f
C537 B.n479 VSUBS 0.007409f
C538 B.n480 VSUBS 0.007409f
C539 B.n481 VSUBS 0.007409f
C540 B.n482 VSUBS 0.007409f
C541 B.n483 VSUBS 0.007409f
C542 B.n484 VSUBS 0.007409f
C543 B.n485 VSUBS 0.007409f
C544 B.n486 VSUBS 0.007409f
C545 B.n487 VSUBS 0.007409f
C546 B.n488 VSUBS 0.007409f
C547 B.n489 VSUBS 0.007409f
C548 B.n490 VSUBS 0.007409f
C549 B.n491 VSUBS 0.007409f
C550 B.n492 VSUBS 0.007409f
C551 B.n493 VSUBS 0.007409f
C552 B.n494 VSUBS 0.007409f
C553 B.n495 VSUBS 0.007409f
C554 B.n496 VSUBS 0.007409f
C555 B.n497 VSUBS 0.007409f
C556 B.n498 VSUBS 0.007409f
C557 B.n499 VSUBS 0.016777f
.ends

