* NGSPICE file created from diff_pair_sample_1543.ext - technology: sky130A

.subckt diff_pair_sample_1543 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.23595 pd=1.76 as=0.5577 ps=3.64 w=1.43 l=0.99
X1 B.t11 B.t9 B.t10 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0 ps=0 w=1.43 l=0.99
X2 VTAIL.t0 VN.t0 VDD2.t3 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0.23595 ps=1.76 w=1.43 l=0.99
X3 B.t8 B.t6 B.t7 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0 ps=0 w=1.43 l=0.99
X4 VTAIL.t6 VP.t1 VDD1.t2 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0.23595 ps=1.76 w=1.43 l=0.99
X5 VDD2.t2 VN.t1 VTAIL.t3 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.23595 pd=1.76 as=0.5577 ps=3.64 w=1.43 l=0.99
X6 VTAIL.t4 VP.t2 VDD1.t1 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0.23595 ps=1.76 w=1.43 l=0.99
X7 B.t5 B.t3 B.t4 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0 ps=0 w=1.43 l=0.99
X8 VDD2.t1 VN.t2 VTAIL.t1 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.23595 pd=1.76 as=0.5577 ps=3.64 w=1.43 l=0.99
X9 B.t2 B.t0 B.t1 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0 ps=0 w=1.43 l=0.99
X10 VTAIL.t2 VN.t3 VDD2.t0 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.5577 pd=3.64 as=0.23595 ps=1.76 w=1.43 l=0.99
X11 VDD1.t0 VP.t3 VTAIL.t7 w_n1762_n1254# sky130_fd_pr__pfet_01v8 ad=0.23595 pd=1.76 as=0.5577 ps=3.64 w=1.43 l=0.99
R0 VP.n0 VP.t1 93.3418
R1 VP.n0 VP.t0 93.2546
R2 VP.n4 VP.n3 80.6037
R3 VP.n2 VP.n1 80.6037
R4 VP.n2 VP.t2 74.7348
R5 VP.n3 VP.t3 74.7348
R6 VP.n1 VP.n0 64.6168
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VTAIL.n5 VTAIL.t6 255.647
R11 VTAIL.n4 VTAIL.t3 255.647
R12 VTAIL.n3 VTAIL.t0 255.647
R13 VTAIL.n7 VTAIL.t1 255.647
R14 VTAIL.n0 VTAIL.t2 255.647
R15 VTAIL.n1 VTAIL.t7 255.647
R16 VTAIL.n2 VTAIL.t4 255.647
R17 VTAIL.n6 VTAIL.t5 255.647
R18 VTAIL.n7 VTAIL.n6 14.7376
R19 VTAIL.n3 VTAIL.n2 14.7376
R20 VTAIL.n4 VTAIL.n3 1.13843
R21 VTAIL.n6 VTAIL.n5 1.13843
R22 VTAIL.n2 VTAIL.n1 1.13843
R23 VTAIL VTAIL.n0 0.627655
R24 VTAIL VTAIL.n7 0.511276
R25 VTAIL.n5 VTAIL.n4 0.470328
R26 VTAIL.n1 VTAIL.n0 0.470328
R27 VDD1 VDD1.n1 278.481
R28 VDD1 VDD1.n0 249.653
R29 VDD1.n0 VDD1.t2 22.7313
R30 VDD1.n0 VDD1.t3 22.7313
R31 VDD1.n1 VDD1.t1 22.7313
R32 VDD1.n1 VDD1.t0 22.7313
R33 B.n154 B.n51 585
R34 B.n153 B.n152 585
R35 B.n151 B.n52 585
R36 B.n150 B.n149 585
R37 B.n148 B.n53 585
R38 B.n147 B.n146 585
R39 B.n145 B.n54 585
R40 B.n144 B.n143 585
R41 B.n142 B.n55 585
R42 B.n141 B.n140 585
R43 B.n139 B.n56 585
R44 B.n138 B.n137 585
R45 B.n133 B.n57 585
R46 B.n132 B.n131 585
R47 B.n130 B.n58 585
R48 B.n129 B.n128 585
R49 B.n127 B.n59 585
R50 B.n126 B.n125 585
R51 B.n124 B.n60 585
R52 B.n123 B.n122 585
R53 B.n120 B.n61 585
R54 B.n119 B.n118 585
R55 B.n117 B.n64 585
R56 B.n116 B.n115 585
R57 B.n114 B.n65 585
R58 B.n113 B.n112 585
R59 B.n111 B.n66 585
R60 B.n110 B.n109 585
R61 B.n108 B.n67 585
R62 B.n107 B.n106 585
R63 B.n105 B.n68 585
R64 B.n156 B.n155 585
R65 B.n157 B.n50 585
R66 B.n159 B.n158 585
R67 B.n160 B.n49 585
R68 B.n162 B.n161 585
R69 B.n163 B.n48 585
R70 B.n165 B.n164 585
R71 B.n166 B.n47 585
R72 B.n168 B.n167 585
R73 B.n169 B.n46 585
R74 B.n171 B.n170 585
R75 B.n172 B.n45 585
R76 B.n174 B.n173 585
R77 B.n175 B.n44 585
R78 B.n177 B.n176 585
R79 B.n178 B.n43 585
R80 B.n180 B.n179 585
R81 B.n181 B.n42 585
R82 B.n183 B.n182 585
R83 B.n184 B.n41 585
R84 B.n186 B.n185 585
R85 B.n187 B.n40 585
R86 B.n189 B.n188 585
R87 B.n190 B.n39 585
R88 B.n192 B.n191 585
R89 B.n193 B.n38 585
R90 B.n195 B.n194 585
R91 B.n196 B.n37 585
R92 B.n198 B.n197 585
R93 B.n199 B.n36 585
R94 B.n201 B.n200 585
R95 B.n202 B.n35 585
R96 B.n204 B.n203 585
R97 B.n205 B.n34 585
R98 B.n207 B.n206 585
R99 B.n208 B.n33 585
R100 B.n210 B.n209 585
R101 B.n211 B.n32 585
R102 B.n213 B.n212 585
R103 B.n214 B.n31 585
R104 B.n263 B.n262 585
R105 B.n261 B.n12 585
R106 B.n260 B.n259 585
R107 B.n258 B.n13 585
R108 B.n257 B.n256 585
R109 B.n255 B.n14 585
R110 B.n254 B.n253 585
R111 B.n252 B.n15 585
R112 B.n251 B.n250 585
R113 B.n249 B.n16 585
R114 B.n248 B.n247 585
R115 B.n245 B.n17 585
R116 B.n244 B.n243 585
R117 B.n242 B.n20 585
R118 B.n241 B.n240 585
R119 B.n239 B.n21 585
R120 B.n238 B.n237 585
R121 B.n236 B.n22 585
R122 B.n235 B.n234 585
R123 B.n233 B.n23 585
R124 B.n231 B.n230 585
R125 B.n229 B.n26 585
R126 B.n228 B.n227 585
R127 B.n226 B.n27 585
R128 B.n225 B.n224 585
R129 B.n223 B.n28 585
R130 B.n222 B.n221 585
R131 B.n220 B.n29 585
R132 B.n219 B.n218 585
R133 B.n217 B.n30 585
R134 B.n216 B.n215 585
R135 B.n264 B.n11 585
R136 B.n266 B.n265 585
R137 B.n267 B.n10 585
R138 B.n269 B.n268 585
R139 B.n270 B.n9 585
R140 B.n272 B.n271 585
R141 B.n273 B.n8 585
R142 B.n275 B.n274 585
R143 B.n276 B.n7 585
R144 B.n278 B.n277 585
R145 B.n279 B.n6 585
R146 B.n281 B.n280 585
R147 B.n282 B.n5 585
R148 B.n284 B.n283 585
R149 B.n285 B.n4 585
R150 B.n287 B.n286 585
R151 B.n288 B.n3 585
R152 B.n290 B.n289 585
R153 B.n291 B.n0 585
R154 B.n2 B.n1 585
R155 B.n78 B.n77 585
R156 B.n80 B.n79 585
R157 B.n81 B.n76 585
R158 B.n83 B.n82 585
R159 B.n84 B.n75 585
R160 B.n86 B.n85 585
R161 B.n87 B.n74 585
R162 B.n89 B.n88 585
R163 B.n90 B.n73 585
R164 B.n92 B.n91 585
R165 B.n93 B.n72 585
R166 B.n95 B.n94 585
R167 B.n96 B.n71 585
R168 B.n98 B.n97 585
R169 B.n99 B.n70 585
R170 B.n101 B.n100 585
R171 B.n102 B.n69 585
R172 B.n104 B.n103 585
R173 B.n105 B.n104 511.721
R174 B.n156 B.n51 511.721
R175 B.n216 B.n31 511.721
R176 B.n262 B.n11 511.721
R177 B.n134 B.t1 274.75
R178 B.n24 B.t5 274.75
R179 B.n62 B.t10 274.75
R180 B.n18 B.t8 274.75
R181 B.n293 B.n292 256.663
R182 B.n135 B.t2 249.15
R183 B.n25 B.t4 249.15
R184 B.n63 B.t11 249.15
R185 B.n19 B.t7 249.15
R186 B.n62 B.t9 237.669
R187 B.n134 B.t0 237.669
R188 B.n24 B.t3 237.669
R189 B.n18 B.t6 237.669
R190 B.n292 B.n291 235.042
R191 B.n292 B.n2 235.042
R192 B.n106 B.n105 163.367
R193 B.n106 B.n67 163.367
R194 B.n110 B.n67 163.367
R195 B.n111 B.n110 163.367
R196 B.n112 B.n111 163.367
R197 B.n112 B.n65 163.367
R198 B.n116 B.n65 163.367
R199 B.n117 B.n116 163.367
R200 B.n118 B.n117 163.367
R201 B.n118 B.n61 163.367
R202 B.n123 B.n61 163.367
R203 B.n124 B.n123 163.367
R204 B.n125 B.n124 163.367
R205 B.n125 B.n59 163.367
R206 B.n129 B.n59 163.367
R207 B.n130 B.n129 163.367
R208 B.n131 B.n130 163.367
R209 B.n131 B.n57 163.367
R210 B.n138 B.n57 163.367
R211 B.n139 B.n138 163.367
R212 B.n140 B.n139 163.367
R213 B.n140 B.n55 163.367
R214 B.n144 B.n55 163.367
R215 B.n145 B.n144 163.367
R216 B.n146 B.n145 163.367
R217 B.n146 B.n53 163.367
R218 B.n150 B.n53 163.367
R219 B.n151 B.n150 163.367
R220 B.n152 B.n151 163.367
R221 B.n152 B.n51 163.367
R222 B.n212 B.n31 163.367
R223 B.n212 B.n211 163.367
R224 B.n211 B.n210 163.367
R225 B.n210 B.n33 163.367
R226 B.n206 B.n33 163.367
R227 B.n206 B.n205 163.367
R228 B.n205 B.n204 163.367
R229 B.n204 B.n35 163.367
R230 B.n200 B.n35 163.367
R231 B.n200 B.n199 163.367
R232 B.n199 B.n198 163.367
R233 B.n198 B.n37 163.367
R234 B.n194 B.n37 163.367
R235 B.n194 B.n193 163.367
R236 B.n193 B.n192 163.367
R237 B.n192 B.n39 163.367
R238 B.n188 B.n39 163.367
R239 B.n188 B.n187 163.367
R240 B.n187 B.n186 163.367
R241 B.n186 B.n41 163.367
R242 B.n182 B.n41 163.367
R243 B.n182 B.n181 163.367
R244 B.n181 B.n180 163.367
R245 B.n180 B.n43 163.367
R246 B.n176 B.n43 163.367
R247 B.n176 B.n175 163.367
R248 B.n175 B.n174 163.367
R249 B.n174 B.n45 163.367
R250 B.n170 B.n45 163.367
R251 B.n170 B.n169 163.367
R252 B.n169 B.n168 163.367
R253 B.n168 B.n47 163.367
R254 B.n164 B.n47 163.367
R255 B.n164 B.n163 163.367
R256 B.n163 B.n162 163.367
R257 B.n162 B.n49 163.367
R258 B.n158 B.n49 163.367
R259 B.n158 B.n157 163.367
R260 B.n157 B.n156 163.367
R261 B.n262 B.n261 163.367
R262 B.n261 B.n260 163.367
R263 B.n260 B.n13 163.367
R264 B.n256 B.n13 163.367
R265 B.n256 B.n255 163.367
R266 B.n255 B.n254 163.367
R267 B.n254 B.n15 163.367
R268 B.n250 B.n15 163.367
R269 B.n250 B.n249 163.367
R270 B.n249 B.n248 163.367
R271 B.n248 B.n17 163.367
R272 B.n243 B.n17 163.367
R273 B.n243 B.n242 163.367
R274 B.n242 B.n241 163.367
R275 B.n241 B.n21 163.367
R276 B.n237 B.n21 163.367
R277 B.n237 B.n236 163.367
R278 B.n236 B.n235 163.367
R279 B.n235 B.n23 163.367
R280 B.n230 B.n23 163.367
R281 B.n230 B.n229 163.367
R282 B.n229 B.n228 163.367
R283 B.n228 B.n27 163.367
R284 B.n224 B.n27 163.367
R285 B.n224 B.n223 163.367
R286 B.n223 B.n222 163.367
R287 B.n222 B.n29 163.367
R288 B.n218 B.n29 163.367
R289 B.n218 B.n217 163.367
R290 B.n217 B.n216 163.367
R291 B.n266 B.n11 163.367
R292 B.n267 B.n266 163.367
R293 B.n268 B.n267 163.367
R294 B.n268 B.n9 163.367
R295 B.n272 B.n9 163.367
R296 B.n273 B.n272 163.367
R297 B.n274 B.n273 163.367
R298 B.n274 B.n7 163.367
R299 B.n278 B.n7 163.367
R300 B.n279 B.n278 163.367
R301 B.n280 B.n279 163.367
R302 B.n280 B.n5 163.367
R303 B.n284 B.n5 163.367
R304 B.n285 B.n284 163.367
R305 B.n286 B.n285 163.367
R306 B.n286 B.n3 163.367
R307 B.n290 B.n3 163.367
R308 B.n291 B.n290 163.367
R309 B.n77 B.n2 163.367
R310 B.n80 B.n77 163.367
R311 B.n81 B.n80 163.367
R312 B.n82 B.n81 163.367
R313 B.n82 B.n75 163.367
R314 B.n86 B.n75 163.367
R315 B.n87 B.n86 163.367
R316 B.n88 B.n87 163.367
R317 B.n88 B.n73 163.367
R318 B.n92 B.n73 163.367
R319 B.n93 B.n92 163.367
R320 B.n94 B.n93 163.367
R321 B.n94 B.n71 163.367
R322 B.n98 B.n71 163.367
R323 B.n99 B.n98 163.367
R324 B.n100 B.n99 163.367
R325 B.n100 B.n69 163.367
R326 B.n104 B.n69 163.367
R327 B.n121 B.n63 59.5399
R328 B.n136 B.n135 59.5399
R329 B.n232 B.n25 59.5399
R330 B.n246 B.n19 59.5399
R331 B.n264 B.n263 33.2493
R332 B.n215 B.n214 33.2493
R333 B.n155 B.n154 33.2493
R334 B.n103 B.n68 33.2493
R335 B.n63 B.n62 25.6005
R336 B.n135 B.n134 25.6005
R337 B.n25 B.n24 25.6005
R338 B.n19 B.n18 25.6005
R339 B B.n293 18.0485
R340 B.n265 B.n264 10.6151
R341 B.n265 B.n10 10.6151
R342 B.n269 B.n10 10.6151
R343 B.n270 B.n269 10.6151
R344 B.n271 B.n270 10.6151
R345 B.n271 B.n8 10.6151
R346 B.n275 B.n8 10.6151
R347 B.n276 B.n275 10.6151
R348 B.n277 B.n276 10.6151
R349 B.n277 B.n6 10.6151
R350 B.n281 B.n6 10.6151
R351 B.n282 B.n281 10.6151
R352 B.n283 B.n282 10.6151
R353 B.n283 B.n4 10.6151
R354 B.n287 B.n4 10.6151
R355 B.n288 B.n287 10.6151
R356 B.n289 B.n288 10.6151
R357 B.n289 B.n0 10.6151
R358 B.n263 B.n12 10.6151
R359 B.n259 B.n12 10.6151
R360 B.n259 B.n258 10.6151
R361 B.n258 B.n257 10.6151
R362 B.n257 B.n14 10.6151
R363 B.n253 B.n14 10.6151
R364 B.n253 B.n252 10.6151
R365 B.n252 B.n251 10.6151
R366 B.n251 B.n16 10.6151
R367 B.n247 B.n16 10.6151
R368 B.n245 B.n244 10.6151
R369 B.n244 B.n20 10.6151
R370 B.n240 B.n20 10.6151
R371 B.n240 B.n239 10.6151
R372 B.n239 B.n238 10.6151
R373 B.n238 B.n22 10.6151
R374 B.n234 B.n22 10.6151
R375 B.n234 B.n233 10.6151
R376 B.n231 B.n26 10.6151
R377 B.n227 B.n26 10.6151
R378 B.n227 B.n226 10.6151
R379 B.n226 B.n225 10.6151
R380 B.n225 B.n28 10.6151
R381 B.n221 B.n28 10.6151
R382 B.n221 B.n220 10.6151
R383 B.n220 B.n219 10.6151
R384 B.n219 B.n30 10.6151
R385 B.n215 B.n30 10.6151
R386 B.n214 B.n213 10.6151
R387 B.n213 B.n32 10.6151
R388 B.n209 B.n32 10.6151
R389 B.n209 B.n208 10.6151
R390 B.n208 B.n207 10.6151
R391 B.n207 B.n34 10.6151
R392 B.n203 B.n34 10.6151
R393 B.n203 B.n202 10.6151
R394 B.n202 B.n201 10.6151
R395 B.n201 B.n36 10.6151
R396 B.n197 B.n36 10.6151
R397 B.n197 B.n196 10.6151
R398 B.n196 B.n195 10.6151
R399 B.n195 B.n38 10.6151
R400 B.n191 B.n38 10.6151
R401 B.n191 B.n190 10.6151
R402 B.n190 B.n189 10.6151
R403 B.n189 B.n40 10.6151
R404 B.n185 B.n40 10.6151
R405 B.n185 B.n184 10.6151
R406 B.n184 B.n183 10.6151
R407 B.n183 B.n42 10.6151
R408 B.n179 B.n42 10.6151
R409 B.n179 B.n178 10.6151
R410 B.n178 B.n177 10.6151
R411 B.n177 B.n44 10.6151
R412 B.n173 B.n44 10.6151
R413 B.n173 B.n172 10.6151
R414 B.n172 B.n171 10.6151
R415 B.n171 B.n46 10.6151
R416 B.n167 B.n46 10.6151
R417 B.n167 B.n166 10.6151
R418 B.n166 B.n165 10.6151
R419 B.n165 B.n48 10.6151
R420 B.n161 B.n48 10.6151
R421 B.n161 B.n160 10.6151
R422 B.n160 B.n159 10.6151
R423 B.n159 B.n50 10.6151
R424 B.n155 B.n50 10.6151
R425 B.n78 B.n1 10.6151
R426 B.n79 B.n78 10.6151
R427 B.n79 B.n76 10.6151
R428 B.n83 B.n76 10.6151
R429 B.n84 B.n83 10.6151
R430 B.n85 B.n84 10.6151
R431 B.n85 B.n74 10.6151
R432 B.n89 B.n74 10.6151
R433 B.n90 B.n89 10.6151
R434 B.n91 B.n90 10.6151
R435 B.n91 B.n72 10.6151
R436 B.n95 B.n72 10.6151
R437 B.n96 B.n95 10.6151
R438 B.n97 B.n96 10.6151
R439 B.n97 B.n70 10.6151
R440 B.n101 B.n70 10.6151
R441 B.n102 B.n101 10.6151
R442 B.n103 B.n102 10.6151
R443 B.n107 B.n68 10.6151
R444 B.n108 B.n107 10.6151
R445 B.n109 B.n108 10.6151
R446 B.n109 B.n66 10.6151
R447 B.n113 B.n66 10.6151
R448 B.n114 B.n113 10.6151
R449 B.n115 B.n114 10.6151
R450 B.n115 B.n64 10.6151
R451 B.n119 B.n64 10.6151
R452 B.n120 B.n119 10.6151
R453 B.n122 B.n60 10.6151
R454 B.n126 B.n60 10.6151
R455 B.n127 B.n126 10.6151
R456 B.n128 B.n127 10.6151
R457 B.n128 B.n58 10.6151
R458 B.n132 B.n58 10.6151
R459 B.n133 B.n132 10.6151
R460 B.n137 B.n133 10.6151
R461 B.n141 B.n56 10.6151
R462 B.n142 B.n141 10.6151
R463 B.n143 B.n142 10.6151
R464 B.n143 B.n54 10.6151
R465 B.n147 B.n54 10.6151
R466 B.n148 B.n147 10.6151
R467 B.n149 B.n148 10.6151
R468 B.n149 B.n52 10.6151
R469 B.n153 B.n52 10.6151
R470 B.n154 B.n153 10.6151
R471 B.n293 B.n0 8.11757
R472 B.n293 B.n1 8.11757
R473 B.n246 B.n245 6.5566
R474 B.n233 B.n232 6.5566
R475 B.n122 B.n121 6.5566
R476 B.n137 B.n136 6.5566
R477 B.n247 B.n246 4.05904
R478 B.n232 B.n231 4.05904
R479 B.n121 B.n120 4.05904
R480 B.n136 B.n56 4.05904
R481 VN.n0 VN.t3 93.3418
R482 VN.n1 VN.t1 93.3418
R483 VN.n1 VN.t0 93.2546
R484 VN.n0 VN.t2 93.2546
R485 VN VN.n1 64.9023
R486 VN VN.n0 31.2622
R487 VDD2.n2 VDD2.n0 277.957
R488 VDD2.n2 VDD2.n1 249.595
R489 VDD2.n1 VDD2.t3 22.7313
R490 VDD2.n1 VDD2.t2 22.7313
R491 VDD2.n0 VDD2.t0 22.7313
R492 VDD2.n0 VDD2.t1 22.7313
R493 VDD2 VDD2.n2 0.0586897
C0 VDD1 w_n1762_n1254# 0.839876f
C1 VDD1 VDD2 0.63663f
C2 VP B 1.01592f
C3 VP VTAIL 0.937352f
C4 VP VN 3.08265f
C5 VP w_n1762_n1254# 2.66573f
C6 VTAIL B 0.984551f
C7 VP VDD2 0.299299f
C8 VN B 0.655289f
C9 VP VDD1 0.838693f
C10 B w_n1762_n1254# 4.29222f
C11 VTAIL VN 0.923245f
C12 VDD2 B 0.717359f
C13 VTAIL w_n1762_n1254# 1.3956f
C14 VDD1 B 0.69115f
C15 VN w_n1762_n1254# 2.44966f
C16 VTAIL VDD2 2.20019f
C17 VN VDD2 0.694776f
C18 VDD1 VTAIL 2.15678f
C19 VDD1 VN 0.154061f
C20 VDD2 w_n1762_n1254# 0.859504f
C21 VDD2 VSUBS 0.428637f
C22 VDD1 VSUBS 2.448827f
C23 VTAIL VSUBS 0.297691f
C24 VN VSUBS 4.30843f
C25 VP VSUBS 0.97465f
C26 B VSUBS 1.884569f
C27 w_n1762_n1254# VSUBS 28.3541f
C28 VDD2.t0 VSUBS 0.023224f
C29 VDD2.t1 VSUBS 0.023224f
C30 VDD2.n0 VSUBS 0.16034f
C31 VDD2.t3 VSUBS 0.023224f
C32 VDD2.t2 VSUBS 0.023224f
C33 VDD2.n1 VSUBS 0.088362f
C34 VDD2.n2 VSUBS 1.77862f
C35 VN.t3 VSUBS 0.303745f
C36 VN.t2 VSUBS 0.303469f
C37 VN.n0 VSUBS 0.341175f
C38 VN.t1 VSUBS 0.303745f
C39 VN.t0 VSUBS 0.303469f
C40 VN.n1 VSUBS 1.25912f
C41 B.n0 VSUBS 0.008548f
C42 B.n1 VSUBS 0.008548f
C43 B.n2 VSUBS 0.012642f
C44 B.n3 VSUBS 0.009688f
C45 B.n4 VSUBS 0.009688f
C46 B.n5 VSUBS 0.009688f
C47 B.n6 VSUBS 0.009688f
C48 B.n7 VSUBS 0.009688f
C49 B.n8 VSUBS 0.009688f
C50 B.n9 VSUBS 0.009688f
C51 B.n10 VSUBS 0.009688f
C52 B.n11 VSUBS 0.021992f
C53 B.n12 VSUBS 0.009688f
C54 B.n13 VSUBS 0.009688f
C55 B.n14 VSUBS 0.009688f
C56 B.n15 VSUBS 0.009688f
C57 B.n16 VSUBS 0.009688f
C58 B.n17 VSUBS 0.009688f
C59 B.t7 VSUBS 0.03994f
C60 B.t8 VSUBS 0.044478f
C61 B.t6 VSUBS 0.096933f
C62 B.n18 VSUBS 0.068326f
C63 B.n19 VSUBS 0.06252f
C64 B.n20 VSUBS 0.009688f
C65 B.n21 VSUBS 0.009688f
C66 B.n22 VSUBS 0.009688f
C67 B.n23 VSUBS 0.009688f
C68 B.t4 VSUBS 0.03994f
C69 B.t5 VSUBS 0.044478f
C70 B.t3 VSUBS 0.096933f
C71 B.n24 VSUBS 0.068326f
C72 B.n25 VSUBS 0.06252f
C73 B.n26 VSUBS 0.009688f
C74 B.n27 VSUBS 0.009688f
C75 B.n28 VSUBS 0.009688f
C76 B.n29 VSUBS 0.009688f
C77 B.n30 VSUBS 0.009688f
C78 B.n31 VSUBS 0.021992f
C79 B.n32 VSUBS 0.009688f
C80 B.n33 VSUBS 0.009688f
C81 B.n34 VSUBS 0.009688f
C82 B.n35 VSUBS 0.009688f
C83 B.n36 VSUBS 0.009688f
C84 B.n37 VSUBS 0.009688f
C85 B.n38 VSUBS 0.009688f
C86 B.n39 VSUBS 0.009688f
C87 B.n40 VSUBS 0.009688f
C88 B.n41 VSUBS 0.009688f
C89 B.n42 VSUBS 0.009688f
C90 B.n43 VSUBS 0.009688f
C91 B.n44 VSUBS 0.009688f
C92 B.n45 VSUBS 0.009688f
C93 B.n46 VSUBS 0.009688f
C94 B.n47 VSUBS 0.009688f
C95 B.n48 VSUBS 0.009688f
C96 B.n49 VSUBS 0.009688f
C97 B.n50 VSUBS 0.009688f
C98 B.n51 VSUBS 0.023884f
C99 B.n52 VSUBS 0.009688f
C100 B.n53 VSUBS 0.009688f
C101 B.n54 VSUBS 0.009688f
C102 B.n55 VSUBS 0.009688f
C103 B.n56 VSUBS 0.006696f
C104 B.n57 VSUBS 0.009688f
C105 B.n58 VSUBS 0.009688f
C106 B.n59 VSUBS 0.009688f
C107 B.n60 VSUBS 0.009688f
C108 B.n61 VSUBS 0.009688f
C109 B.t11 VSUBS 0.03994f
C110 B.t10 VSUBS 0.044478f
C111 B.t9 VSUBS 0.096933f
C112 B.n62 VSUBS 0.068326f
C113 B.n63 VSUBS 0.06252f
C114 B.n64 VSUBS 0.009688f
C115 B.n65 VSUBS 0.009688f
C116 B.n66 VSUBS 0.009688f
C117 B.n67 VSUBS 0.009688f
C118 B.n68 VSUBS 0.023884f
C119 B.n69 VSUBS 0.009688f
C120 B.n70 VSUBS 0.009688f
C121 B.n71 VSUBS 0.009688f
C122 B.n72 VSUBS 0.009688f
C123 B.n73 VSUBS 0.009688f
C124 B.n74 VSUBS 0.009688f
C125 B.n75 VSUBS 0.009688f
C126 B.n76 VSUBS 0.009688f
C127 B.n77 VSUBS 0.009688f
C128 B.n78 VSUBS 0.009688f
C129 B.n79 VSUBS 0.009688f
C130 B.n80 VSUBS 0.009688f
C131 B.n81 VSUBS 0.009688f
C132 B.n82 VSUBS 0.009688f
C133 B.n83 VSUBS 0.009688f
C134 B.n84 VSUBS 0.009688f
C135 B.n85 VSUBS 0.009688f
C136 B.n86 VSUBS 0.009688f
C137 B.n87 VSUBS 0.009688f
C138 B.n88 VSUBS 0.009688f
C139 B.n89 VSUBS 0.009688f
C140 B.n90 VSUBS 0.009688f
C141 B.n91 VSUBS 0.009688f
C142 B.n92 VSUBS 0.009688f
C143 B.n93 VSUBS 0.009688f
C144 B.n94 VSUBS 0.009688f
C145 B.n95 VSUBS 0.009688f
C146 B.n96 VSUBS 0.009688f
C147 B.n97 VSUBS 0.009688f
C148 B.n98 VSUBS 0.009688f
C149 B.n99 VSUBS 0.009688f
C150 B.n100 VSUBS 0.009688f
C151 B.n101 VSUBS 0.009688f
C152 B.n102 VSUBS 0.009688f
C153 B.n103 VSUBS 0.021992f
C154 B.n104 VSUBS 0.021992f
C155 B.n105 VSUBS 0.023884f
C156 B.n106 VSUBS 0.009688f
C157 B.n107 VSUBS 0.009688f
C158 B.n108 VSUBS 0.009688f
C159 B.n109 VSUBS 0.009688f
C160 B.n110 VSUBS 0.009688f
C161 B.n111 VSUBS 0.009688f
C162 B.n112 VSUBS 0.009688f
C163 B.n113 VSUBS 0.009688f
C164 B.n114 VSUBS 0.009688f
C165 B.n115 VSUBS 0.009688f
C166 B.n116 VSUBS 0.009688f
C167 B.n117 VSUBS 0.009688f
C168 B.n118 VSUBS 0.009688f
C169 B.n119 VSUBS 0.009688f
C170 B.n120 VSUBS 0.006696f
C171 B.n121 VSUBS 0.022446f
C172 B.n122 VSUBS 0.007836f
C173 B.n123 VSUBS 0.009688f
C174 B.n124 VSUBS 0.009688f
C175 B.n125 VSUBS 0.009688f
C176 B.n126 VSUBS 0.009688f
C177 B.n127 VSUBS 0.009688f
C178 B.n128 VSUBS 0.009688f
C179 B.n129 VSUBS 0.009688f
C180 B.n130 VSUBS 0.009688f
C181 B.n131 VSUBS 0.009688f
C182 B.n132 VSUBS 0.009688f
C183 B.n133 VSUBS 0.009688f
C184 B.t2 VSUBS 0.03994f
C185 B.t1 VSUBS 0.044478f
C186 B.t0 VSUBS 0.096933f
C187 B.n134 VSUBS 0.068326f
C188 B.n135 VSUBS 0.06252f
C189 B.n136 VSUBS 0.022446f
C190 B.n137 VSUBS 0.007836f
C191 B.n138 VSUBS 0.009688f
C192 B.n139 VSUBS 0.009688f
C193 B.n140 VSUBS 0.009688f
C194 B.n141 VSUBS 0.009688f
C195 B.n142 VSUBS 0.009688f
C196 B.n143 VSUBS 0.009688f
C197 B.n144 VSUBS 0.009688f
C198 B.n145 VSUBS 0.009688f
C199 B.n146 VSUBS 0.009688f
C200 B.n147 VSUBS 0.009688f
C201 B.n148 VSUBS 0.009688f
C202 B.n149 VSUBS 0.009688f
C203 B.n150 VSUBS 0.009688f
C204 B.n151 VSUBS 0.009688f
C205 B.n152 VSUBS 0.009688f
C206 B.n153 VSUBS 0.009688f
C207 B.n154 VSUBS 0.02276f
C208 B.n155 VSUBS 0.023116f
C209 B.n156 VSUBS 0.021992f
C210 B.n157 VSUBS 0.009688f
C211 B.n158 VSUBS 0.009688f
C212 B.n159 VSUBS 0.009688f
C213 B.n160 VSUBS 0.009688f
C214 B.n161 VSUBS 0.009688f
C215 B.n162 VSUBS 0.009688f
C216 B.n163 VSUBS 0.009688f
C217 B.n164 VSUBS 0.009688f
C218 B.n165 VSUBS 0.009688f
C219 B.n166 VSUBS 0.009688f
C220 B.n167 VSUBS 0.009688f
C221 B.n168 VSUBS 0.009688f
C222 B.n169 VSUBS 0.009688f
C223 B.n170 VSUBS 0.009688f
C224 B.n171 VSUBS 0.009688f
C225 B.n172 VSUBS 0.009688f
C226 B.n173 VSUBS 0.009688f
C227 B.n174 VSUBS 0.009688f
C228 B.n175 VSUBS 0.009688f
C229 B.n176 VSUBS 0.009688f
C230 B.n177 VSUBS 0.009688f
C231 B.n178 VSUBS 0.009688f
C232 B.n179 VSUBS 0.009688f
C233 B.n180 VSUBS 0.009688f
C234 B.n181 VSUBS 0.009688f
C235 B.n182 VSUBS 0.009688f
C236 B.n183 VSUBS 0.009688f
C237 B.n184 VSUBS 0.009688f
C238 B.n185 VSUBS 0.009688f
C239 B.n186 VSUBS 0.009688f
C240 B.n187 VSUBS 0.009688f
C241 B.n188 VSUBS 0.009688f
C242 B.n189 VSUBS 0.009688f
C243 B.n190 VSUBS 0.009688f
C244 B.n191 VSUBS 0.009688f
C245 B.n192 VSUBS 0.009688f
C246 B.n193 VSUBS 0.009688f
C247 B.n194 VSUBS 0.009688f
C248 B.n195 VSUBS 0.009688f
C249 B.n196 VSUBS 0.009688f
C250 B.n197 VSUBS 0.009688f
C251 B.n198 VSUBS 0.009688f
C252 B.n199 VSUBS 0.009688f
C253 B.n200 VSUBS 0.009688f
C254 B.n201 VSUBS 0.009688f
C255 B.n202 VSUBS 0.009688f
C256 B.n203 VSUBS 0.009688f
C257 B.n204 VSUBS 0.009688f
C258 B.n205 VSUBS 0.009688f
C259 B.n206 VSUBS 0.009688f
C260 B.n207 VSUBS 0.009688f
C261 B.n208 VSUBS 0.009688f
C262 B.n209 VSUBS 0.009688f
C263 B.n210 VSUBS 0.009688f
C264 B.n211 VSUBS 0.009688f
C265 B.n212 VSUBS 0.009688f
C266 B.n213 VSUBS 0.009688f
C267 B.n214 VSUBS 0.021992f
C268 B.n215 VSUBS 0.023884f
C269 B.n216 VSUBS 0.023884f
C270 B.n217 VSUBS 0.009688f
C271 B.n218 VSUBS 0.009688f
C272 B.n219 VSUBS 0.009688f
C273 B.n220 VSUBS 0.009688f
C274 B.n221 VSUBS 0.009688f
C275 B.n222 VSUBS 0.009688f
C276 B.n223 VSUBS 0.009688f
C277 B.n224 VSUBS 0.009688f
C278 B.n225 VSUBS 0.009688f
C279 B.n226 VSUBS 0.009688f
C280 B.n227 VSUBS 0.009688f
C281 B.n228 VSUBS 0.009688f
C282 B.n229 VSUBS 0.009688f
C283 B.n230 VSUBS 0.009688f
C284 B.n231 VSUBS 0.006696f
C285 B.n232 VSUBS 0.022446f
C286 B.n233 VSUBS 0.007836f
C287 B.n234 VSUBS 0.009688f
C288 B.n235 VSUBS 0.009688f
C289 B.n236 VSUBS 0.009688f
C290 B.n237 VSUBS 0.009688f
C291 B.n238 VSUBS 0.009688f
C292 B.n239 VSUBS 0.009688f
C293 B.n240 VSUBS 0.009688f
C294 B.n241 VSUBS 0.009688f
C295 B.n242 VSUBS 0.009688f
C296 B.n243 VSUBS 0.009688f
C297 B.n244 VSUBS 0.009688f
C298 B.n245 VSUBS 0.007836f
C299 B.n246 VSUBS 0.022446f
C300 B.n247 VSUBS 0.006696f
C301 B.n248 VSUBS 0.009688f
C302 B.n249 VSUBS 0.009688f
C303 B.n250 VSUBS 0.009688f
C304 B.n251 VSUBS 0.009688f
C305 B.n252 VSUBS 0.009688f
C306 B.n253 VSUBS 0.009688f
C307 B.n254 VSUBS 0.009688f
C308 B.n255 VSUBS 0.009688f
C309 B.n256 VSUBS 0.009688f
C310 B.n257 VSUBS 0.009688f
C311 B.n258 VSUBS 0.009688f
C312 B.n259 VSUBS 0.009688f
C313 B.n260 VSUBS 0.009688f
C314 B.n261 VSUBS 0.009688f
C315 B.n262 VSUBS 0.023884f
C316 B.n263 VSUBS 0.023884f
C317 B.n264 VSUBS 0.021992f
C318 B.n265 VSUBS 0.009688f
C319 B.n266 VSUBS 0.009688f
C320 B.n267 VSUBS 0.009688f
C321 B.n268 VSUBS 0.009688f
C322 B.n269 VSUBS 0.009688f
C323 B.n270 VSUBS 0.009688f
C324 B.n271 VSUBS 0.009688f
C325 B.n272 VSUBS 0.009688f
C326 B.n273 VSUBS 0.009688f
C327 B.n274 VSUBS 0.009688f
C328 B.n275 VSUBS 0.009688f
C329 B.n276 VSUBS 0.009688f
C330 B.n277 VSUBS 0.009688f
C331 B.n278 VSUBS 0.009688f
C332 B.n279 VSUBS 0.009688f
C333 B.n280 VSUBS 0.009688f
C334 B.n281 VSUBS 0.009688f
C335 B.n282 VSUBS 0.009688f
C336 B.n283 VSUBS 0.009688f
C337 B.n284 VSUBS 0.009688f
C338 B.n285 VSUBS 0.009688f
C339 B.n286 VSUBS 0.009688f
C340 B.n287 VSUBS 0.009688f
C341 B.n288 VSUBS 0.009688f
C342 B.n289 VSUBS 0.009688f
C343 B.n290 VSUBS 0.009688f
C344 B.n291 VSUBS 0.012642f
C345 B.n292 VSUBS 0.013467f
C346 B.n293 VSUBS 0.026781f
C347 VDD1.t2 VSUBS 0.022449f
C348 VDD1.t3 VSUBS 0.022449f
C349 VDD1.n0 VSUBS 0.085476f
C350 VDD1.t1 VSUBS 0.022449f
C351 VDD1.t0 VSUBS 0.022449f
C352 VDD1.n1 VSUBS 0.160399f
C353 VTAIL.t2 VSUBS 0.114394f
C354 VTAIL.n0 VSUBS 0.225151f
C355 VTAIL.t7 VSUBS 0.114394f
C356 VTAIL.n1 VSUBS 0.25527f
C357 VTAIL.t4 VSUBS 0.114394f
C358 VTAIL.n2 VSUBS 0.615942f
C359 VTAIL.t0 VSUBS 0.114394f
C360 VTAIL.n3 VSUBS 0.615942f
C361 VTAIL.t3 VSUBS 0.114394f
C362 VTAIL.n4 VSUBS 0.25527f
C363 VTAIL.t6 VSUBS 0.114394f
C364 VTAIL.n5 VSUBS 0.25527f
C365 VTAIL.t5 VSUBS 0.114394f
C366 VTAIL.n6 VSUBS 0.615942f
C367 VTAIL.t1 VSUBS 0.114394f
C368 VTAIL.n7 VSUBS 0.57896f
C369 VP.t0 VSUBS 0.32478f
C370 VP.t1 VSUBS 0.325076f
C371 VP.n0 VSUBS 1.32489f
C372 VP.n1 VSUBS 2.67746f
C373 VP.t2 VSUBS 0.279703f
C374 VP.n2 VSUBS 0.226981f
C375 VP.t3 VSUBS 0.279703f
C376 VP.n3 VSUBS 0.226981f
C377 VP.n4 VSUBS 0.077967f
.ends

