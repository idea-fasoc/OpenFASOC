* NGSPICE file created from diff_pair_sample_0120.ext - technology: sky130A

.subckt diff_pair_sample_0120 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0.7029 ps=4.59 w=4.26 l=2.21
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0 ps=0 w=4.26 l=2.21
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0 ps=0 w=4.26 l=2.21
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0 ps=0 w=4.26 l=2.21
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0 ps=0 w=4.26 l=2.21
X5 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7029 pd=4.59 as=1.6614 ps=9.3 w=4.26 l=2.21
X6 VTAIL.t6 VN.t1 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0.7029 ps=4.59 w=4.26 l=2.21
X7 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0.7029 ps=4.59 w=4.26 l=2.21
X8 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6614 pd=9.3 as=0.7029 ps=4.59 w=4.26 l=2.21
X9 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7029 pd=4.59 as=1.6614 ps=9.3 w=4.26 l=2.21
X10 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7029 pd=4.59 as=1.6614 ps=9.3 w=4.26 l=2.21
X11 VDD2.t2 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7029 pd=4.59 as=1.6614 ps=9.3 w=4.26 l=2.21
R0 VN.n0 VN.t0 82.285
R1 VN.n1 VN.t2 82.285
R2 VN.n0 VN.t3 81.6462
R3 VN.n1 VN.t1 81.6462
R4 VN VN.n1 45.2564
R5 VN VN.n0 5.79803
R6 VDD2.n2 VDD2.n0 107.038
R7 VDD2.n2 VDD2.n1 73.0819
R8 VDD2.n1 VDD2.t1 4.64839
R9 VDD2.n1 VDD2.t3 4.64839
R10 VDD2.n0 VDD2.t0 4.64839
R11 VDD2.n0 VDD2.t2 4.64839
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t2 61.0512
R14 VTAIL.n4 VTAIL.t5 61.0512
R15 VTAIL.n3 VTAIL.t6 61.0512
R16 VTAIL.n7 VTAIL.t4 61.051
R17 VTAIL.n0 VTAIL.t7 61.051
R18 VTAIL.n1 VTAIL.t3 61.051
R19 VTAIL.n2 VTAIL.t1 61.051
R20 VTAIL.n6 VTAIL.t0 61.051
R21 VTAIL.n3 VTAIL.n2 18.2289
R22 VTAIL.n7 VTAIL.n6 18.2289
R23 VTAIL.n4 VTAIL.n3 2.19016
R24 VTAIL.n6 VTAIL.n5 2.19016
R25 VTAIL.n2 VTAIL.n1 2.19016
R26 VTAIL VTAIL.n0 1.15352
R27 VTAIL VTAIL.n7 1.03714
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n399 B.n398 585
R31 B.n399 B.n58 585
R32 B.n402 B.n401 585
R33 B.n403 B.n86 585
R34 B.n405 B.n404 585
R35 B.n407 B.n85 585
R36 B.n410 B.n409 585
R37 B.n411 B.n84 585
R38 B.n413 B.n412 585
R39 B.n415 B.n83 585
R40 B.n418 B.n417 585
R41 B.n419 B.n82 585
R42 B.n421 B.n420 585
R43 B.n423 B.n81 585
R44 B.n426 B.n425 585
R45 B.n427 B.n80 585
R46 B.n429 B.n428 585
R47 B.n431 B.n79 585
R48 B.n434 B.n433 585
R49 B.n435 B.n76 585
R50 B.n438 B.n437 585
R51 B.n440 B.n75 585
R52 B.n443 B.n442 585
R53 B.n444 B.n74 585
R54 B.n446 B.n445 585
R55 B.n448 B.n73 585
R56 B.n451 B.n450 585
R57 B.n452 B.n69 585
R58 B.n454 B.n453 585
R59 B.n456 B.n68 585
R60 B.n459 B.n458 585
R61 B.n460 B.n67 585
R62 B.n462 B.n461 585
R63 B.n464 B.n66 585
R64 B.n467 B.n466 585
R65 B.n468 B.n65 585
R66 B.n470 B.n469 585
R67 B.n472 B.n64 585
R68 B.n475 B.n474 585
R69 B.n476 B.n63 585
R70 B.n478 B.n477 585
R71 B.n480 B.n62 585
R72 B.n483 B.n482 585
R73 B.n484 B.n61 585
R74 B.n486 B.n485 585
R75 B.n488 B.n60 585
R76 B.n491 B.n490 585
R77 B.n492 B.n59 585
R78 B.n397 B.n57 585
R79 B.n495 B.n57 585
R80 B.n396 B.n56 585
R81 B.n496 B.n56 585
R82 B.n395 B.n55 585
R83 B.n497 B.n55 585
R84 B.n394 B.n393 585
R85 B.n393 B.n51 585
R86 B.n392 B.n50 585
R87 B.n503 B.n50 585
R88 B.n391 B.n49 585
R89 B.n504 B.n49 585
R90 B.n390 B.n48 585
R91 B.n505 B.n48 585
R92 B.n389 B.n388 585
R93 B.n388 B.n47 585
R94 B.n387 B.n43 585
R95 B.n511 B.n43 585
R96 B.n386 B.n42 585
R97 B.n512 B.n42 585
R98 B.n385 B.n41 585
R99 B.n513 B.n41 585
R100 B.n384 B.n383 585
R101 B.n383 B.n37 585
R102 B.n382 B.n36 585
R103 B.n519 B.n36 585
R104 B.n381 B.n35 585
R105 B.n520 B.n35 585
R106 B.n380 B.n34 585
R107 B.n521 B.n34 585
R108 B.n379 B.n378 585
R109 B.n378 B.n30 585
R110 B.n377 B.n29 585
R111 B.n527 B.n29 585
R112 B.n376 B.n28 585
R113 B.n528 B.n28 585
R114 B.n375 B.n27 585
R115 B.n529 B.n27 585
R116 B.n374 B.n373 585
R117 B.n373 B.n23 585
R118 B.n372 B.n22 585
R119 B.n535 B.n22 585
R120 B.n371 B.n21 585
R121 B.n536 B.n21 585
R122 B.n370 B.n20 585
R123 B.n537 B.n20 585
R124 B.n369 B.n368 585
R125 B.n368 B.n16 585
R126 B.n367 B.n15 585
R127 B.n543 B.n15 585
R128 B.n366 B.n14 585
R129 B.n544 B.n14 585
R130 B.n365 B.n13 585
R131 B.n545 B.n13 585
R132 B.n364 B.n363 585
R133 B.n363 B.n12 585
R134 B.n362 B.n361 585
R135 B.n362 B.n8 585
R136 B.n360 B.n7 585
R137 B.n552 B.n7 585
R138 B.n359 B.n6 585
R139 B.n553 B.n6 585
R140 B.n358 B.n5 585
R141 B.n554 B.n5 585
R142 B.n357 B.n356 585
R143 B.n356 B.n4 585
R144 B.n355 B.n87 585
R145 B.n355 B.n354 585
R146 B.n345 B.n88 585
R147 B.n89 B.n88 585
R148 B.n347 B.n346 585
R149 B.n348 B.n347 585
R150 B.n344 B.n93 585
R151 B.n97 B.n93 585
R152 B.n343 B.n342 585
R153 B.n342 B.n341 585
R154 B.n95 B.n94 585
R155 B.n96 B.n95 585
R156 B.n334 B.n333 585
R157 B.n335 B.n334 585
R158 B.n332 B.n102 585
R159 B.n102 B.n101 585
R160 B.n331 B.n330 585
R161 B.n330 B.n329 585
R162 B.n104 B.n103 585
R163 B.n105 B.n104 585
R164 B.n322 B.n321 585
R165 B.n323 B.n322 585
R166 B.n320 B.n109 585
R167 B.n113 B.n109 585
R168 B.n319 B.n318 585
R169 B.n318 B.n317 585
R170 B.n111 B.n110 585
R171 B.n112 B.n111 585
R172 B.n310 B.n309 585
R173 B.n311 B.n310 585
R174 B.n308 B.n118 585
R175 B.n118 B.n117 585
R176 B.n307 B.n306 585
R177 B.n306 B.n305 585
R178 B.n120 B.n119 585
R179 B.n121 B.n120 585
R180 B.n298 B.n297 585
R181 B.n299 B.n298 585
R182 B.n296 B.n126 585
R183 B.n126 B.n125 585
R184 B.n295 B.n294 585
R185 B.n294 B.n293 585
R186 B.n128 B.n127 585
R187 B.n286 B.n128 585
R188 B.n285 B.n284 585
R189 B.n287 B.n285 585
R190 B.n283 B.n133 585
R191 B.n133 B.n132 585
R192 B.n282 B.n281 585
R193 B.n281 B.n280 585
R194 B.n135 B.n134 585
R195 B.n136 B.n135 585
R196 B.n273 B.n272 585
R197 B.n274 B.n273 585
R198 B.n271 B.n141 585
R199 B.n141 B.n140 585
R200 B.n270 B.n269 585
R201 B.n269 B.n268 585
R202 B.n265 B.n145 585
R203 B.n264 B.n263 585
R204 B.n261 B.n146 585
R205 B.n261 B.n144 585
R206 B.n260 B.n259 585
R207 B.n258 B.n257 585
R208 B.n256 B.n148 585
R209 B.n254 B.n253 585
R210 B.n252 B.n149 585
R211 B.n251 B.n250 585
R212 B.n248 B.n150 585
R213 B.n246 B.n245 585
R214 B.n244 B.n151 585
R215 B.n243 B.n242 585
R216 B.n240 B.n152 585
R217 B.n238 B.n237 585
R218 B.n236 B.n153 585
R219 B.n235 B.n234 585
R220 B.n232 B.n154 585
R221 B.n230 B.n229 585
R222 B.n227 B.n155 585
R223 B.n226 B.n225 585
R224 B.n223 B.n158 585
R225 B.n221 B.n220 585
R226 B.n219 B.n159 585
R227 B.n218 B.n217 585
R228 B.n215 B.n160 585
R229 B.n213 B.n212 585
R230 B.n211 B.n161 585
R231 B.n209 B.n208 585
R232 B.n206 B.n164 585
R233 B.n204 B.n203 585
R234 B.n202 B.n165 585
R235 B.n201 B.n200 585
R236 B.n198 B.n166 585
R237 B.n196 B.n195 585
R238 B.n194 B.n167 585
R239 B.n193 B.n192 585
R240 B.n190 B.n168 585
R241 B.n188 B.n187 585
R242 B.n186 B.n169 585
R243 B.n185 B.n184 585
R244 B.n182 B.n170 585
R245 B.n180 B.n179 585
R246 B.n178 B.n171 585
R247 B.n177 B.n176 585
R248 B.n174 B.n172 585
R249 B.n143 B.n142 585
R250 B.n267 B.n266 585
R251 B.n268 B.n267 585
R252 B.n139 B.n138 585
R253 B.n140 B.n139 585
R254 B.n276 B.n275 585
R255 B.n275 B.n274 585
R256 B.n277 B.n137 585
R257 B.n137 B.n136 585
R258 B.n279 B.n278 585
R259 B.n280 B.n279 585
R260 B.n131 B.n130 585
R261 B.n132 B.n131 585
R262 B.n289 B.n288 585
R263 B.n288 B.n287 585
R264 B.n290 B.n129 585
R265 B.n286 B.n129 585
R266 B.n292 B.n291 585
R267 B.n293 B.n292 585
R268 B.n124 B.n123 585
R269 B.n125 B.n124 585
R270 B.n301 B.n300 585
R271 B.n300 B.n299 585
R272 B.n302 B.n122 585
R273 B.n122 B.n121 585
R274 B.n304 B.n303 585
R275 B.n305 B.n304 585
R276 B.n116 B.n115 585
R277 B.n117 B.n116 585
R278 B.n313 B.n312 585
R279 B.n312 B.n311 585
R280 B.n314 B.n114 585
R281 B.n114 B.n112 585
R282 B.n316 B.n315 585
R283 B.n317 B.n316 585
R284 B.n108 B.n107 585
R285 B.n113 B.n108 585
R286 B.n325 B.n324 585
R287 B.n324 B.n323 585
R288 B.n326 B.n106 585
R289 B.n106 B.n105 585
R290 B.n328 B.n327 585
R291 B.n329 B.n328 585
R292 B.n100 B.n99 585
R293 B.n101 B.n100 585
R294 B.n337 B.n336 585
R295 B.n336 B.n335 585
R296 B.n338 B.n98 585
R297 B.n98 B.n96 585
R298 B.n340 B.n339 585
R299 B.n341 B.n340 585
R300 B.n92 B.n91 585
R301 B.n97 B.n92 585
R302 B.n350 B.n349 585
R303 B.n349 B.n348 585
R304 B.n351 B.n90 585
R305 B.n90 B.n89 585
R306 B.n353 B.n352 585
R307 B.n354 B.n353 585
R308 B.n3 B.n0 585
R309 B.n4 B.n3 585
R310 B.n551 B.n1 585
R311 B.n552 B.n551 585
R312 B.n550 B.n549 585
R313 B.n550 B.n8 585
R314 B.n548 B.n9 585
R315 B.n12 B.n9 585
R316 B.n547 B.n546 585
R317 B.n546 B.n545 585
R318 B.n11 B.n10 585
R319 B.n544 B.n11 585
R320 B.n542 B.n541 585
R321 B.n543 B.n542 585
R322 B.n540 B.n17 585
R323 B.n17 B.n16 585
R324 B.n539 B.n538 585
R325 B.n538 B.n537 585
R326 B.n19 B.n18 585
R327 B.n536 B.n19 585
R328 B.n534 B.n533 585
R329 B.n535 B.n534 585
R330 B.n532 B.n24 585
R331 B.n24 B.n23 585
R332 B.n531 B.n530 585
R333 B.n530 B.n529 585
R334 B.n26 B.n25 585
R335 B.n528 B.n26 585
R336 B.n526 B.n525 585
R337 B.n527 B.n526 585
R338 B.n524 B.n31 585
R339 B.n31 B.n30 585
R340 B.n523 B.n522 585
R341 B.n522 B.n521 585
R342 B.n33 B.n32 585
R343 B.n520 B.n33 585
R344 B.n518 B.n517 585
R345 B.n519 B.n518 585
R346 B.n516 B.n38 585
R347 B.n38 B.n37 585
R348 B.n515 B.n514 585
R349 B.n514 B.n513 585
R350 B.n40 B.n39 585
R351 B.n512 B.n40 585
R352 B.n510 B.n509 585
R353 B.n511 B.n510 585
R354 B.n508 B.n44 585
R355 B.n47 B.n44 585
R356 B.n507 B.n506 585
R357 B.n506 B.n505 585
R358 B.n46 B.n45 585
R359 B.n504 B.n46 585
R360 B.n502 B.n501 585
R361 B.n503 B.n502 585
R362 B.n500 B.n52 585
R363 B.n52 B.n51 585
R364 B.n499 B.n498 585
R365 B.n498 B.n497 585
R366 B.n54 B.n53 585
R367 B.n496 B.n54 585
R368 B.n494 B.n493 585
R369 B.n495 B.n494 585
R370 B.n555 B.n554 585
R371 B.n553 B.n2 585
R372 B.n494 B.n59 526.135
R373 B.n399 B.n57 526.135
R374 B.n269 B.n143 526.135
R375 B.n267 B.n145 526.135
R376 B.n400 B.n58 256.663
R377 B.n406 B.n58 256.663
R378 B.n408 B.n58 256.663
R379 B.n414 B.n58 256.663
R380 B.n416 B.n58 256.663
R381 B.n422 B.n58 256.663
R382 B.n424 B.n58 256.663
R383 B.n430 B.n58 256.663
R384 B.n432 B.n58 256.663
R385 B.n439 B.n58 256.663
R386 B.n441 B.n58 256.663
R387 B.n447 B.n58 256.663
R388 B.n449 B.n58 256.663
R389 B.n455 B.n58 256.663
R390 B.n457 B.n58 256.663
R391 B.n463 B.n58 256.663
R392 B.n465 B.n58 256.663
R393 B.n471 B.n58 256.663
R394 B.n473 B.n58 256.663
R395 B.n479 B.n58 256.663
R396 B.n481 B.n58 256.663
R397 B.n487 B.n58 256.663
R398 B.n489 B.n58 256.663
R399 B.n262 B.n144 256.663
R400 B.n147 B.n144 256.663
R401 B.n255 B.n144 256.663
R402 B.n249 B.n144 256.663
R403 B.n247 B.n144 256.663
R404 B.n241 B.n144 256.663
R405 B.n239 B.n144 256.663
R406 B.n233 B.n144 256.663
R407 B.n231 B.n144 256.663
R408 B.n224 B.n144 256.663
R409 B.n222 B.n144 256.663
R410 B.n216 B.n144 256.663
R411 B.n214 B.n144 256.663
R412 B.n207 B.n144 256.663
R413 B.n205 B.n144 256.663
R414 B.n199 B.n144 256.663
R415 B.n197 B.n144 256.663
R416 B.n191 B.n144 256.663
R417 B.n189 B.n144 256.663
R418 B.n183 B.n144 256.663
R419 B.n181 B.n144 256.663
R420 B.n175 B.n144 256.663
R421 B.n173 B.n144 256.663
R422 B.n557 B.n556 256.663
R423 B.n70 B.t12 253.827
R424 B.n77 B.t8 253.827
R425 B.n162 B.t4 253.827
R426 B.n156 B.t15 253.827
R427 B.n490 B.n488 163.367
R428 B.n486 B.n61 163.367
R429 B.n482 B.n480 163.367
R430 B.n478 B.n63 163.367
R431 B.n474 B.n472 163.367
R432 B.n470 B.n65 163.367
R433 B.n466 B.n464 163.367
R434 B.n462 B.n67 163.367
R435 B.n458 B.n456 163.367
R436 B.n454 B.n69 163.367
R437 B.n450 B.n448 163.367
R438 B.n446 B.n74 163.367
R439 B.n442 B.n440 163.367
R440 B.n438 B.n76 163.367
R441 B.n433 B.n431 163.367
R442 B.n429 B.n80 163.367
R443 B.n425 B.n423 163.367
R444 B.n421 B.n82 163.367
R445 B.n417 B.n415 163.367
R446 B.n413 B.n84 163.367
R447 B.n409 B.n407 163.367
R448 B.n405 B.n86 163.367
R449 B.n401 B.n399 163.367
R450 B.n269 B.n141 163.367
R451 B.n273 B.n141 163.367
R452 B.n273 B.n135 163.367
R453 B.n281 B.n135 163.367
R454 B.n281 B.n133 163.367
R455 B.n285 B.n133 163.367
R456 B.n285 B.n128 163.367
R457 B.n294 B.n128 163.367
R458 B.n294 B.n126 163.367
R459 B.n298 B.n126 163.367
R460 B.n298 B.n120 163.367
R461 B.n306 B.n120 163.367
R462 B.n306 B.n118 163.367
R463 B.n310 B.n118 163.367
R464 B.n310 B.n111 163.367
R465 B.n318 B.n111 163.367
R466 B.n318 B.n109 163.367
R467 B.n322 B.n109 163.367
R468 B.n322 B.n104 163.367
R469 B.n330 B.n104 163.367
R470 B.n330 B.n102 163.367
R471 B.n334 B.n102 163.367
R472 B.n334 B.n95 163.367
R473 B.n342 B.n95 163.367
R474 B.n342 B.n93 163.367
R475 B.n347 B.n93 163.367
R476 B.n347 B.n88 163.367
R477 B.n355 B.n88 163.367
R478 B.n356 B.n355 163.367
R479 B.n356 B.n5 163.367
R480 B.n6 B.n5 163.367
R481 B.n7 B.n6 163.367
R482 B.n362 B.n7 163.367
R483 B.n363 B.n362 163.367
R484 B.n363 B.n13 163.367
R485 B.n14 B.n13 163.367
R486 B.n15 B.n14 163.367
R487 B.n368 B.n15 163.367
R488 B.n368 B.n20 163.367
R489 B.n21 B.n20 163.367
R490 B.n22 B.n21 163.367
R491 B.n373 B.n22 163.367
R492 B.n373 B.n27 163.367
R493 B.n28 B.n27 163.367
R494 B.n29 B.n28 163.367
R495 B.n378 B.n29 163.367
R496 B.n378 B.n34 163.367
R497 B.n35 B.n34 163.367
R498 B.n36 B.n35 163.367
R499 B.n383 B.n36 163.367
R500 B.n383 B.n41 163.367
R501 B.n42 B.n41 163.367
R502 B.n43 B.n42 163.367
R503 B.n388 B.n43 163.367
R504 B.n388 B.n48 163.367
R505 B.n49 B.n48 163.367
R506 B.n50 B.n49 163.367
R507 B.n393 B.n50 163.367
R508 B.n393 B.n55 163.367
R509 B.n56 B.n55 163.367
R510 B.n57 B.n56 163.367
R511 B.n263 B.n261 163.367
R512 B.n261 B.n260 163.367
R513 B.n257 B.n256 163.367
R514 B.n254 B.n149 163.367
R515 B.n250 B.n248 163.367
R516 B.n246 B.n151 163.367
R517 B.n242 B.n240 163.367
R518 B.n238 B.n153 163.367
R519 B.n234 B.n232 163.367
R520 B.n230 B.n155 163.367
R521 B.n225 B.n223 163.367
R522 B.n221 B.n159 163.367
R523 B.n217 B.n215 163.367
R524 B.n213 B.n161 163.367
R525 B.n208 B.n206 163.367
R526 B.n204 B.n165 163.367
R527 B.n200 B.n198 163.367
R528 B.n196 B.n167 163.367
R529 B.n192 B.n190 163.367
R530 B.n188 B.n169 163.367
R531 B.n184 B.n182 163.367
R532 B.n180 B.n171 163.367
R533 B.n176 B.n174 163.367
R534 B.n267 B.n139 163.367
R535 B.n275 B.n139 163.367
R536 B.n275 B.n137 163.367
R537 B.n279 B.n137 163.367
R538 B.n279 B.n131 163.367
R539 B.n288 B.n131 163.367
R540 B.n288 B.n129 163.367
R541 B.n292 B.n129 163.367
R542 B.n292 B.n124 163.367
R543 B.n300 B.n124 163.367
R544 B.n300 B.n122 163.367
R545 B.n304 B.n122 163.367
R546 B.n304 B.n116 163.367
R547 B.n312 B.n116 163.367
R548 B.n312 B.n114 163.367
R549 B.n316 B.n114 163.367
R550 B.n316 B.n108 163.367
R551 B.n324 B.n108 163.367
R552 B.n324 B.n106 163.367
R553 B.n328 B.n106 163.367
R554 B.n328 B.n100 163.367
R555 B.n336 B.n100 163.367
R556 B.n336 B.n98 163.367
R557 B.n340 B.n98 163.367
R558 B.n340 B.n92 163.367
R559 B.n349 B.n92 163.367
R560 B.n349 B.n90 163.367
R561 B.n353 B.n90 163.367
R562 B.n353 B.n3 163.367
R563 B.n555 B.n3 163.367
R564 B.n551 B.n2 163.367
R565 B.n551 B.n550 163.367
R566 B.n550 B.n9 163.367
R567 B.n546 B.n9 163.367
R568 B.n546 B.n11 163.367
R569 B.n542 B.n11 163.367
R570 B.n542 B.n17 163.367
R571 B.n538 B.n17 163.367
R572 B.n538 B.n19 163.367
R573 B.n534 B.n19 163.367
R574 B.n534 B.n24 163.367
R575 B.n530 B.n24 163.367
R576 B.n530 B.n26 163.367
R577 B.n526 B.n26 163.367
R578 B.n526 B.n31 163.367
R579 B.n522 B.n31 163.367
R580 B.n522 B.n33 163.367
R581 B.n518 B.n33 163.367
R582 B.n518 B.n38 163.367
R583 B.n514 B.n38 163.367
R584 B.n514 B.n40 163.367
R585 B.n510 B.n40 163.367
R586 B.n510 B.n44 163.367
R587 B.n506 B.n44 163.367
R588 B.n506 B.n46 163.367
R589 B.n502 B.n46 163.367
R590 B.n502 B.n52 163.367
R591 B.n498 B.n52 163.367
R592 B.n498 B.n54 163.367
R593 B.n494 B.n54 163.367
R594 B.n268 B.n144 144.207
R595 B.n495 B.n58 144.207
R596 B.n77 B.t10 123.814
R597 B.n162 B.t7 123.814
R598 B.n70 B.t13 123.811
R599 B.n156 B.t17 123.811
R600 B.n268 B.n140 78.4483
R601 B.n274 B.n140 78.4483
R602 B.n274 B.n136 78.4483
R603 B.n280 B.n136 78.4483
R604 B.n280 B.n132 78.4483
R605 B.n287 B.n132 78.4483
R606 B.n287 B.n286 78.4483
R607 B.n293 B.n125 78.4483
R608 B.n299 B.n125 78.4483
R609 B.n299 B.n121 78.4483
R610 B.n305 B.n121 78.4483
R611 B.n305 B.n117 78.4483
R612 B.n311 B.n117 78.4483
R613 B.n311 B.n112 78.4483
R614 B.n317 B.n112 78.4483
R615 B.n317 B.n113 78.4483
R616 B.n323 B.n105 78.4483
R617 B.n329 B.n105 78.4483
R618 B.n329 B.n101 78.4483
R619 B.n335 B.n101 78.4483
R620 B.n335 B.n96 78.4483
R621 B.n341 B.n96 78.4483
R622 B.n341 B.n97 78.4483
R623 B.n348 B.n89 78.4483
R624 B.n354 B.n89 78.4483
R625 B.n354 B.n4 78.4483
R626 B.n554 B.n4 78.4483
R627 B.n554 B.n553 78.4483
R628 B.n553 B.n552 78.4483
R629 B.n552 B.n8 78.4483
R630 B.n12 B.n8 78.4483
R631 B.n545 B.n12 78.4483
R632 B.n544 B.n543 78.4483
R633 B.n543 B.n16 78.4483
R634 B.n537 B.n16 78.4483
R635 B.n537 B.n536 78.4483
R636 B.n536 B.n535 78.4483
R637 B.n535 B.n23 78.4483
R638 B.n529 B.n23 78.4483
R639 B.n528 B.n527 78.4483
R640 B.n527 B.n30 78.4483
R641 B.n521 B.n30 78.4483
R642 B.n521 B.n520 78.4483
R643 B.n520 B.n519 78.4483
R644 B.n519 B.n37 78.4483
R645 B.n513 B.n37 78.4483
R646 B.n513 B.n512 78.4483
R647 B.n512 B.n511 78.4483
R648 B.n505 B.n47 78.4483
R649 B.n505 B.n504 78.4483
R650 B.n504 B.n503 78.4483
R651 B.n503 B.n51 78.4483
R652 B.n497 B.n51 78.4483
R653 B.n497 B.n496 78.4483
R654 B.n496 B.n495 78.4483
R655 B.n293 B.t5 77.2947
R656 B.n511 B.t9 77.2947
R657 B.n78 B.t11 74.5533
R658 B.n163 B.t6 74.5533
R659 B.n71 B.t14 74.5494
R660 B.n157 B.t16 74.5494
R661 B.n489 B.n59 71.676
R662 B.n488 B.n487 71.676
R663 B.n481 B.n61 71.676
R664 B.n480 B.n479 71.676
R665 B.n473 B.n63 71.676
R666 B.n472 B.n471 71.676
R667 B.n465 B.n65 71.676
R668 B.n464 B.n463 71.676
R669 B.n457 B.n67 71.676
R670 B.n456 B.n455 71.676
R671 B.n449 B.n69 71.676
R672 B.n448 B.n447 71.676
R673 B.n441 B.n74 71.676
R674 B.n440 B.n439 71.676
R675 B.n432 B.n76 71.676
R676 B.n431 B.n430 71.676
R677 B.n424 B.n80 71.676
R678 B.n423 B.n422 71.676
R679 B.n416 B.n82 71.676
R680 B.n415 B.n414 71.676
R681 B.n408 B.n84 71.676
R682 B.n407 B.n406 71.676
R683 B.n400 B.n86 71.676
R684 B.n401 B.n400 71.676
R685 B.n406 B.n405 71.676
R686 B.n409 B.n408 71.676
R687 B.n414 B.n413 71.676
R688 B.n417 B.n416 71.676
R689 B.n422 B.n421 71.676
R690 B.n425 B.n424 71.676
R691 B.n430 B.n429 71.676
R692 B.n433 B.n432 71.676
R693 B.n439 B.n438 71.676
R694 B.n442 B.n441 71.676
R695 B.n447 B.n446 71.676
R696 B.n450 B.n449 71.676
R697 B.n455 B.n454 71.676
R698 B.n458 B.n457 71.676
R699 B.n463 B.n462 71.676
R700 B.n466 B.n465 71.676
R701 B.n471 B.n470 71.676
R702 B.n474 B.n473 71.676
R703 B.n479 B.n478 71.676
R704 B.n482 B.n481 71.676
R705 B.n487 B.n486 71.676
R706 B.n490 B.n489 71.676
R707 B.n262 B.n145 71.676
R708 B.n260 B.n147 71.676
R709 B.n256 B.n255 71.676
R710 B.n249 B.n149 71.676
R711 B.n248 B.n247 71.676
R712 B.n241 B.n151 71.676
R713 B.n240 B.n239 71.676
R714 B.n233 B.n153 71.676
R715 B.n232 B.n231 71.676
R716 B.n224 B.n155 71.676
R717 B.n223 B.n222 71.676
R718 B.n216 B.n159 71.676
R719 B.n215 B.n214 71.676
R720 B.n207 B.n161 71.676
R721 B.n206 B.n205 71.676
R722 B.n199 B.n165 71.676
R723 B.n198 B.n197 71.676
R724 B.n191 B.n167 71.676
R725 B.n190 B.n189 71.676
R726 B.n183 B.n169 71.676
R727 B.n182 B.n181 71.676
R728 B.n175 B.n171 71.676
R729 B.n174 B.n173 71.676
R730 B.n263 B.n262 71.676
R731 B.n257 B.n147 71.676
R732 B.n255 B.n254 71.676
R733 B.n250 B.n249 71.676
R734 B.n247 B.n246 71.676
R735 B.n242 B.n241 71.676
R736 B.n239 B.n238 71.676
R737 B.n234 B.n233 71.676
R738 B.n231 B.n230 71.676
R739 B.n225 B.n224 71.676
R740 B.n222 B.n221 71.676
R741 B.n217 B.n216 71.676
R742 B.n214 B.n213 71.676
R743 B.n208 B.n207 71.676
R744 B.n205 B.n204 71.676
R745 B.n200 B.n199 71.676
R746 B.n197 B.n196 71.676
R747 B.n192 B.n191 71.676
R748 B.n189 B.n188 71.676
R749 B.n184 B.n183 71.676
R750 B.n181 B.n180 71.676
R751 B.n176 B.n175 71.676
R752 B.n173 B.n143 71.676
R753 B.n556 B.n555 71.676
R754 B.n556 B.n2 71.676
R755 B.n348 B.t3 65.7582
R756 B.n545 B.t2 65.7582
R757 B.n72 B.n71 59.5399
R758 B.n436 B.n78 59.5399
R759 B.n210 B.n163 59.5399
R760 B.n228 B.n157 59.5399
R761 B.n113 B.t1 54.2218
R762 B.t0 B.n528 54.2218
R763 B.n71 B.n70 49.2611
R764 B.n78 B.n77 49.2611
R765 B.n163 B.n162 49.2611
R766 B.n157 B.n156 49.2611
R767 B.n266 B.n265 34.1859
R768 B.n270 B.n142 34.1859
R769 B.n398 B.n397 34.1859
R770 B.n493 B.n492 34.1859
R771 B.n323 B.t1 24.227
R772 B.n529 B.t0 24.227
R773 B B.n557 18.0485
R774 B.n97 B.t3 12.6906
R775 B.t2 B.n544 12.6906
R776 B.n266 B.n138 10.6151
R777 B.n276 B.n138 10.6151
R778 B.n277 B.n276 10.6151
R779 B.n278 B.n277 10.6151
R780 B.n278 B.n130 10.6151
R781 B.n289 B.n130 10.6151
R782 B.n290 B.n289 10.6151
R783 B.n291 B.n290 10.6151
R784 B.n291 B.n123 10.6151
R785 B.n301 B.n123 10.6151
R786 B.n302 B.n301 10.6151
R787 B.n303 B.n302 10.6151
R788 B.n303 B.n115 10.6151
R789 B.n313 B.n115 10.6151
R790 B.n314 B.n313 10.6151
R791 B.n315 B.n314 10.6151
R792 B.n315 B.n107 10.6151
R793 B.n325 B.n107 10.6151
R794 B.n326 B.n325 10.6151
R795 B.n327 B.n326 10.6151
R796 B.n327 B.n99 10.6151
R797 B.n337 B.n99 10.6151
R798 B.n338 B.n337 10.6151
R799 B.n339 B.n338 10.6151
R800 B.n339 B.n91 10.6151
R801 B.n350 B.n91 10.6151
R802 B.n351 B.n350 10.6151
R803 B.n352 B.n351 10.6151
R804 B.n352 B.n0 10.6151
R805 B.n265 B.n264 10.6151
R806 B.n264 B.n146 10.6151
R807 B.n259 B.n146 10.6151
R808 B.n259 B.n258 10.6151
R809 B.n258 B.n148 10.6151
R810 B.n253 B.n148 10.6151
R811 B.n253 B.n252 10.6151
R812 B.n252 B.n251 10.6151
R813 B.n251 B.n150 10.6151
R814 B.n245 B.n150 10.6151
R815 B.n245 B.n244 10.6151
R816 B.n244 B.n243 10.6151
R817 B.n243 B.n152 10.6151
R818 B.n237 B.n152 10.6151
R819 B.n237 B.n236 10.6151
R820 B.n236 B.n235 10.6151
R821 B.n235 B.n154 10.6151
R822 B.n229 B.n154 10.6151
R823 B.n227 B.n226 10.6151
R824 B.n226 B.n158 10.6151
R825 B.n220 B.n158 10.6151
R826 B.n220 B.n219 10.6151
R827 B.n219 B.n218 10.6151
R828 B.n218 B.n160 10.6151
R829 B.n212 B.n160 10.6151
R830 B.n212 B.n211 10.6151
R831 B.n209 B.n164 10.6151
R832 B.n203 B.n164 10.6151
R833 B.n203 B.n202 10.6151
R834 B.n202 B.n201 10.6151
R835 B.n201 B.n166 10.6151
R836 B.n195 B.n166 10.6151
R837 B.n195 B.n194 10.6151
R838 B.n194 B.n193 10.6151
R839 B.n193 B.n168 10.6151
R840 B.n187 B.n168 10.6151
R841 B.n187 B.n186 10.6151
R842 B.n186 B.n185 10.6151
R843 B.n185 B.n170 10.6151
R844 B.n179 B.n170 10.6151
R845 B.n179 B.n178 10.6151
R846 B.n178 B.n177 10.6151
R847 B.n177 B.n172 10.6151
R848 B.n172 B.n142 10.6151
R849 B.n271 B.n270 10.6151
R850 B.n272 B.n271 10.6151
R851 B.n272 B.n134 10.6151
R852 B.n282 B.n134 10.6151
R853 B.n283 B.n282 10.6151
R854 B.n284 B.n283 10.6151
R855 B.n284 B.n127 10.6151
R856 B.n295 B.n127 10.6151
R857 B.n296 B.n295 10.6151
R858 B.n297 B.n296 10.6151
R859 B.n297 B.n119 10.6151
R860 B.n307 B.n119 10.6151
R861 B.n308 B.n307 10.6151
R862 B.n309 B.n308 10.6151
R863 B.n309 B.n110 10.6151
R864 B.n319 B.n110 10.6151
R865 B.n320 B.n319 10.6151
R866 B.n321 B.n320 10.6151
R867 B.n321 B.n103 10.6151
R868 B.n331 B.n103 10.6151
R869 B.n332 B.n331 10.6151
R870 B.n333 B.n332 10.6151
R871 B.n333 B.n94 10.6151
R872 B.n343 B.n94 10.6151
R873 B.n344 B.n343 10.6151
R874 B.n346 B.n344 10.6151
R875 B.n346 B.n345 10.6151
R876 B.n345 B.n87 10.6151
R877 B.n357 B.n87 10.6151
R878 B.n358 B.n357 10.6151
R879 B.n359 B.n358 10.6151
R880 B.n360 B.n359 10.6151
R881 B.n361 B.n360 10.6151
R882 B.n364 B.n361 10.6151
R883 B.n365 B.n364 10.6151
R884 B.n366 B.n365 10.6151
R885 B.n367 B.n366 10.6151
R886 B.n369 B.n367 10.6151
R887 B.n370 B.n369 10.6151
R888 B.n371 B.n370 10.6151
R889 B.n372 B.n371 10.6151
R890 B.n374 B.n372 10.6151
R891 B.n375 B.n374 10.6151
R892 B.n376 B.n375 10.6151
R893 B.n377 B.n376 10.6151
R894 B.n379 B.n377 10.6151
R895 B.n380 B.n379 10.6151
R896 B.n381 B.n380 10.6151
R897 B.n382 B.n381 10.6151
R898 B.n384 B.n382 10.6151
R899 B.n385 B.n384 10.6151
R900 B.n386 B.n385 10.6151
R901 B.n387 B.n386 10.6151
R902 B.n389 B.n387 10.6151
R903 B.n390 B.n389 10.6151
R904 B.n391 B.n390 10.6151
R905 B.n392 B.n391 10.6151
R906 B.n394 B.n392 10.6151
R907 B.n395 B.n394 10.6151
R908 B.n396 B.n395 10.6151
R909 B.n397 B.n396 10.6151
R910 B.n549 B.n1 10.6151
R911 B.n549 B.n548 10.6151
R912 B.n548 B.n547 10.6151
R913 B.n547 B.n10 10.6151
R914 B.n541 B.n10 10.6151
R915 B.n541 B.n540 10.6151
R916 B.n540 B.n539 10.6151
R917 B.n539 B.n18 10.6151
R918 B.n533 B.n18 10.6151
R919 B.n533 B.n532 10.6151
R920 B.n532 B.n531 10.6151
R921 B.n531 B.n25 10.6151
R922 B.n525 B.n25 10.6151
R923 B.n525 B.n524 10.6151
R924 B.n524 B.n523 10.6151
R925 B.n523 B.n32 10.6151
R926 B.n517 B.n32 10.6151
R927 B.n517 B.n516 10.6151
R928 B.n516 B.n515 10.6151
R929 B.n515 B.n39 10.6151
R930 B.n509 B.n39 10.6151
R931 B.n509 B.n508 10.6151
R932 B.n508 B.n507 10.6151
R933 B.n507 B.n45 10.6151
R934 B.n501 B.n45 10.6151
R935 B.n501 B.n500 10.6151
R936 B.n500 B.n499 10.6151
R937 B.n499 B.n53 10.6151
R938 B.n493 B.n53 10.6151
R939 B.n492 B.n491 10.6151
R940 B.n491 B.n60 10.6151
R941 B.n485 B.n60 10.6151
R942 B.n485 B.n484 10.6151
R943 B.n484 B.n483 10.6151
R944 B.n483 B.n62 10.6151
R945 B.n477 B.n62 10.6151
R946 B.n477 B.n476 10.6151
R947 B.n476 B.n475 10.6151
R948 B.n475 B.n64 10.6151
R949 B.n469 B.n64 10.6151
R950 B.n469 B.n468 10.6151
R951 B.n468 B.n467 10.6151
R952 B.n467 B.n66 10.6151
R953 B.n461 B.n66 10.6151
R954 B.n461 B.n460 10.6151
R955 B.n460 B.n459 10.6151
R956 B.n459 B.n68 10.6151
R957 B.n453 B.n452 10.6151
R958 B.n452 B.n451 10.6151
R959 B.n451 B.n73 10.6151
R960 B.n445 B.n73 10.6151
R961 B.n445 B.n444 10.6151
R962 B.n444 B.n443 10.6151
R963 B.n443 B.n75 10.6151
R964 B.n437 B.n75 10.6151
R965 B.n435 B.n434 10.6151
R966 B.n434 B.n79 10.6151
R967 B.n428 B.n79 10.6151
R968 B.n428 B.n427 10.6151
R969 B.n427 B.n426 10.6151
R970 B.n426 B.n81 10.6151
R971 B.n420 B.n81 10.6151
R972 B.n420 B.n419 10.6151
R973 B.n419 B.n418 10.6151
R974 B.n418 B.n83 10.6151
R975 B.n412 B.n83 10.6151
R976 B.n412 B.n411 10.6151
R977 B.n411 B.n410 10.6151
R978 B.n410 B.n85 10.6151
R979 B.n404 B.n85 10.6151
R980 B.n404 B.n403 10.6151
R981 B.n403 B.n402 10.6151
R982 B.n402 B.n398 10.6151
R983 B.n557 B.n0 8.11757
R984 B.n557 B.n1 8.11757
R985 B.n228 B.n227 6.5566
R986 B.n211 B.n210 6.5566
R987 B.n453 B.n72 6.5566
R988 B.n437 B.n436 6.5566
R989 B.n229 B.n228 4.05904
R990 B.n210 B.n209 4.05904
R991 B.n72 B.n68 4.05904
R992 B.n436 B.n435 4.05904
R993 B.n286 B.t5 1.15414
R994 B.n47 B.t9 1.15414
R995 VP.n12 VP.n0 161.3
R996 VP.n11 VP.n10 161.3
R997 VP.n9 VP.n1 161.3
R998 VP.n8 VP.n7 161.3
R999 VP.n6 VP.n2 161.3
R1000 VP.n5 VP.n4 97.6287
R1001 VP.n14 VP.n13 97.6287
R1002 VP.n3 VP.t2 82.285
R1003 VP.n3 VP.t0 81.6462
R1004 VP.n5 VP.t1 46.4557
R1005 VP.n13 VP.t3 46.4557
R1006 VP.n4 VP.n3 44.9775
R1007 VP.n7 VP.n1 40.577
R1008 VP.n11 VP.n1 40.577
R1009 VP.n7 VP.n6 24.5923
R1010 VP.n12 VP.n11 24.5923
R1011 VP.n6 VP.n5 13.2801
R1012 VP.n13 VP.n12 13.2801
R1013 VP.n4 VP.n2 0.278335
R1014 VP.n14 VP.n0 0.278335
R1015 VP.n8 VP.n2 0.189894
R1016 VP.n9 VP.n8 0.189894
R1017 VP.n10 VP.n9 0.189894
R1018 VP.n10 VP.n0 0.189894
R1019 VP VP.n14 0.153485
R1020 VDD1 VDD1.n1 107.562
R1021 VDD1 VDD1.n0 73.1401
R1022 VDD1.n0 VDD1.t1 4.64839
R1023 VDD1.n0 VDD1.t3 4.64839
R1024 VDD1.n1 VDD1.t2 4.64839
R1025 VDD1.n1 VDD1.t0 4.64839
C0 VN VDD2 1.84307f
C1 VN VDD1 0.152928f
C2 VN VTAIL 2.14884f
C3 VP VDD2 0.374169f
C4 VP VDD1 2.06324f
C5 VTAIL VP 2.16294f
C6 VDD1 VDD2 0.93437f
C7 VTAIL VDD2 3.45976f
C8 VTAIL VDD1 3.40817f
C9 VN VP 4.48102f
C10 VDD2 B 2.864832f
C11 VDD1 B 6.1965f
C12 VTAIL B 4.988487f
C13 VN B 8.901589f
C14 VP B 7.436295f
C15 VDD1.t1 B 0.094992f
C16 VDD1.t3 B 0.094992f
C17 VDD1.n0 B 0.755075f
C18 VDD1.t2 B 0.094992f
C19 VDD1.t0 B 0.094992f
C20 VDD1.n1 B 1.15442f
C21 VP.n0 B 0.04524f
C22 VP.t3 B 0.834561f
C23 VP.n1 B 0.027716f
C24 VP.n2 B 0.04524f
C25 VP.t1 B 0.834561f
C26 VP.t0 B 1.05976f
C27 VP.t2 B 1.06382f
C28 VP.n3 B 2.06383f
C29 VP.n4 B 1.53068f
C30 VP.n5 B 0.435353f
C31 VP.n6 B 0.049185f
C32 VP.n7 B 0.067844f
C33 VP.n8 B 0.034316f
C34 VP.n9 B 0.034316f
C35 VP.n10 B 0.034316f
C36 VP.n11 B 0.067844f
C37 VP.n12 B 0.049185f
C38 VP.n13 B 0.435353f
C39 VP.n14 B 0.049176f
C40 VTAIL.t7 B 0.660775f
C41 VTAIL.n0 B 0.342704f
C42 VTAIL.t3 B 0.660775f
C43 VTAIL.n1 B 0.413082f
C44 VTAIL.t1 B 0.660775f
C45 VTAIL.n2 B 1.06537f
C46 VTAIL.t6 B 0.660777f
C47 VTAIL.n3 B 1.06537f
C48 VTAIL.t5 B 0.660777f
C49 VTAIL.n4 B 0.41308f
C50 VTAIL.t2 B 0.660777f
C51 VTAIL.n5 B 0.41308f
C52 VTAIL.t0 B 0.660775f
C53 VTAIL.n6 B 1.06537f
C54 VTAIL.t4 B 0.660775f
C55 VTAIL.n7 B 0.987089f
C56 VDD2.t0 B 0.061617f
C57 VDD2.t2 B 0.061617f
C58 VDD2.n0 B 0.734352f
C59 VDD2.t1 B 0.061617f
C60 VDD2.t3 B 0.061617f
C61 VDD2.n1 B 0.489558f
C62 VDD2.n2 B 1.89654f
C63 VN.t0 B 0.793515f
C64 VN.t3 B 0.790485f
C65 VN.n0 B 0.522402f
C66 VN.t2 B 0.793515f
C67 VN.t1 B 0.790485f
C68 VN.n1 B 1.5529f
.ends

