* NGSPICE file created from diff_pair_sample_1017.ext - technology: sky130A

.subckt diff_pair_sample_1017 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X1 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=0 ps=0 w=9.44 l=1.12
X2 VDD1.t4 VP.t1 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=3.6816 ps=19.66 w=9.44 l=1.12
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=0 ps=0 w=9.44 l=1.12
X4 VTAIL.t17 VP.t2 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X5 VDD1.t3 VP.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=1.5576 ps=9.77 w=9.44 l=1.12
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=0 ps=0 w=9.44 l=1.12
X7 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=1.5576 ps=9.77 w=9.44 l=1.12
X8 VDD2.t8 VN.t1 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=3.6816 ps=19.66 w=9.44 l=1.12
X9 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X10 VTAIL.t5 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X11 VDD2.t5 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X12 VTAIL.t7 VN.t5 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X13 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=1.5576 ps=9.77 w=9.44 l=1.12
X14 VDD1.t5 VP.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=3.6816 ps=19.66 w=9.44 l=1.12
X15 VTAIL.t14 VP.t5 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X16 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=3.6816 ps=19.66 w=9.44 l=1.12
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=0 ps=0 w=9.44 l=1.12
X18 VDD1.t1 VP.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6816 pd=19.66 as=1.5576 ps=9.77 w=9.44 l=1.12
X19 VTAIL.t12 VP.t7 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X20 VTAIL.t4 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X21 VDD1.t0 VP.t8 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X22 VTAIL.t8 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
X23 VDD1.t9 VP.t9 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5576 pd=9.77 as=1.5576 ps=9.77 w=9.44 l=1.12
R0 VP.n10 VP.t3 260.755
R1 VP.n5 VP.t6 238.203
R2 VP.n41 VP.t1 238.203
R3 VP.n23 VP.t4 238.203
R4 VP.n34 VP.t9 203.13
R5 VP.n29 VP.t7 203.13
R6 VP.n1 VP.t0 203.13
R7 VP.n16 VP.t8 203.13
R8 VP.n7 VP.t2 203.13
R9 VP.n11 VP.t5 203.13
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n9 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n8 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n22 VP.n6 161.3
R17 VP.n40 VP.n0 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n2 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n3 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n28 VP.n4 161.3
R25 VP.n27 VP.n26 161.3
R26 VP.n24 VP.n23 80.6037
R27 VP.n42 VP.n41 80.6037
R28 VP.n25 VP.n5 80.6037
R29 VP.n30 VP.n3 56.5617
R30 VP.n36 VP.n35 56.5617
R31 VP.n18 VP.n17 56.5617
R32 VP.n12 VP.n9 56.5617
R33 VP.n27 VP.n5 48.6923
R34 VP.n41 VP.n40 48.6923
R35 VP.n23 VP.n22 48.6923
R36 VP.n25 VP.n24 43.3006
R37 VP.n11 VP.n10 34.7238
R38 VP.n13 VP.n10 28.3586
R39 VP.n28 VP.n27 24.5923
R40 VP.n34 VP.n3 24.5923
R41 VP.n35 VP.n34 24.5923
R42 VP.n40 VP.n39 24.5923
R43 VP.n22 VP.n21 24.5923
R44 VP.n16 VP.n9 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n30 VP.n29 22.1332
R47 VP.n36 VP.n1 22.1332
R48 VP.n18 VP.n7 22.1332
R49 VP.n12 VP.n11 22.1332
R50 VP.n29 VP.n28 2.45968
R51 VP.n39 VP.n1 2.45968
R52 VP.n21 VP.n7 2.45968
R53 VP.n24 VP.n6 0.285035
R54 VP.n26 VP.n25 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n14 VP.n13 0.189894
R57 VP.n15 VP.n14 0.189894
R58 VP.n15 VP.n8 0.189894
R59 VP.n19 VP.n8 0.189894
R60 VP.n20 VP.n19 0.189894
R61 VP.n20 VP.n6 0.189894
R62 VP.n26 VP.n4 0.189894
R63 VP.n31 VP.n4 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n33 VP.n2 0.189894
R67 VP.n37 VP.n2 0.189894
R68 VP.n38 VP.n37 0.189894
R69 VP.n38 VP.n0 0.189894
R70 VP VP.n42 0.146778
R71 VDD1.n44 VDD1.n0 289.615
R72 VDD1.n95 VDD1.n51 289.615
R73 VDD1.n45 VDD1.n44 185
R74 VDD1.n43 VDD1.n42 185
R75 VDD1.n4 VDD1.n3 185
R76 VDD1.n8 VDD1.n6 185
R77 VDD1.n37 VDD1.n36 185
R78 VDD1.n35 VDD1.n34 185
R79 VDD1.n10 VDD1.n9 185
R80 VDD1.n29 VDD1.n28 185
R81 VDD1.n27 VDD1.n26 185
R82 VDD1.n14 VDD1.n13 185
R83 VDD1.n21 VDD1.n20 185
R84 VDD1.n19 VDD1.n18 185
R85 VDD1.n68 VDD1.n67 185
R86 VDD1.n70 VDD1.n69 185
R87 VDD1.n63 VDD1.n62 185
R88 VDD1.n76 VDD1.n75 185
R89 VDD1.n78 VDD1.n77 185
R90 VDD1.n59 VDD1.n58 185
R91 VDD1.n85 VDD1.n84 185
R92 VDD1.n86 VDD1.n57 185
R93 VDD1.n88 VDD1.n87 185
R94 VDD1.n55 VDD1.n54 185
R95 VDD1.n94 VDD1.n93 185
R96 VDD1.n96 VDD1.n95 185
R97 VDD1.n17 VDD1.t3 149.524
R98 VDD1.n66 VDD1.t1 149.524
R99 VDD1.n44 VDD1.n43 104.615
R100 VDD1.n43 VDD1.n3 104.615
R101 VDD1.n8 VDD1.n3 104.615
R102 VDD1.n36 VDD1.n8 104.615
R103 VDD1.n36 VDD1.n35 104.615
R104 VDD1.n35 VDD1.n9 104.615
R105 VDD1.n28 VDD1.n9 104.615
R106 VDD1.n28 VDD1.n27 104.615
R107 VDD1.n27 VDD1.n13 104.615
R108 VDD1.n20 VDD1.n13 104.615
R109 VDD1.n20 VDD1.n19 104.615
R110 VDD1.n69 VDD1.n68 104.615
R111 VDD1.n69 VDD1.n62 104.615
R112 VDD1.n76 VDD1.n62 104.615
R113 VDD1.n77 VDD1.n76 104.615
R114 VDD1.n77 VDD1.n58 104.615
R115 VDD1.n85 VDD1.n58 104.615
R116 VDD1.n86 VDD1.n85 104.615
R117 VDD1.n87 VDD1.n86 104.615
R118 VDD1.n87 VDD1.n54 104.615
R119 VDD1.n94 VDD1.n54 104.615
R120 VDD1.n95 VDD1.n94 104.615
R121 VDD1.n103 VDD1.n102 67.7628
R122 VDD1.n50 VDD1.n49 66.8808
R123 VDD1.n105 VDD1.n104 66.8807
R124 VDD1.n101 VDD1.n100 66.8807
R125 VDD1.n50 VDD1.n48 53.9929
R126 VDD1.n101 VDD1.n99 53.9929
R127 VDD1.n19 VDD1.t3 52.3082
R128 VDD1.n68 VDD1.t1 52.3082
R129 VDD1.n105 VDD1.n103 38.9987
R130 VDD1.n6 VDD1.n4 13.1884
R131 VDD1.n88 VDD1.n55 13.1884
R132 VDD1.n42 VDD1.n41 12.8005
R133 VDD1.n38 VDD1.n37 12.8005
R134 VDD1.n89 VDD1.n57 12.8005
R135 VDD1.n93 VDD1.n92 12.8005
R136 VDD1.n45 VDD1.n2 12.0247
R137 VDD1.n34 VDD1.n7 12.0247
R138 VDD1.n84 VDD1.n83 12.0247
R139 VDD1.n96 VDD1.n53 12.0247
R140 VDD1.n46 VDD1.n0 11.249
R141 VDD1.n33 VDD1.n10 11.249
R142 VDD1.n82 VDD1.n59 11.249
R143 VDD1.n97 VDD1.n51 11.249
R144 VDD1.n30 VDD1.n29 10.4732
R145 VDD1.n79 VDD1.n78 10.4732
R146 VDD1.n18 VDD1.n17 10.2747
R147 VDD1.n67 VDD1.n66 10.2747
R148 VDD1.n26 VDD1.n12 9.69747
R149 VDD1.n75 VDD1.n61 9.69747
R150 VDD1.n48 VDD1.n47 9.45567
R151 VDD1.n99 VDD1.n98 9.45567
R152 VDD1.n16 VDD1.n15 9.3005
R153 VDD1.n23 VDD1.n22 9.3005
R154 VDD1.n25 VDD1.n24 9.3005
R155 VDD1.n12 VDD1.n11 9.3005
R156 VDD1.n31 VDD1.n30 9.3005
R157 VDD1.n33 VDD1.n32 9.3005
R158 VDD1.n7 VDD1.n5 9.3005
R159 VDD1.n39 VDD1.n38 9.3005
R160 VDD1.n47 VDD1.n46 9.3005
R161 VDD1.n2 VDD1.n1 9.3005
R162 VDD1.n41 VDD1.n40 9.3005
R163 VDD1.n98 VDD1.n97 9.3005
R164 VDD1.n53 VDD1.n52 9.3005
R165 VDD1.n92 VDD1.n91 9.3005
R166 VDD1.n65 VDD1.n64 9.3005
R167 VDD1.n72 VDD1.n71 9.3005
R168 VDD1.n74 VDD1.n73 9.3005
R169 VDD1.n61 VDD1.n60 9.3005
R170 VDD1.n80 VDD1.n79 9.3005
R171 VDD1.n82 VDD1.n81 9.3005
R172 VDD1.n83 VDD1.n56 9.3005
R173 VDD1.n90 VDD1.n89 9.3005
R174 VDD1.n25 VDD1.n14 8.92171
R175 VDD1.n74 VDD1.n63 8.92171
R176 VDD1.n22 VDD1.n21 8.14595
R177 VDD1.n71 VDD1.n70 8.14595
R178 VDD1.n18 VDD1.n16 7.3702
R179 VDD1.n67 VDD1.n65 7.3702
R180 VDD1.n21 VDD1.n16 5.81868
R181 VDD1.n70 VDD1.n65 5.81868
R182 VDD1.n22 VDD1.n14 5.04292
R183 VDD1.n71 VDD1.n63 5.04292
R184 VDD1.n26 VDD1.n25 4.26717
R185 VDD1.n75 VDD1.n74 4.26717
R186 VDD1.n29 VDD1.n12 3.49141
R187 VDD1.n78 VDD1.n61 3.49141
R188 VDD1.n17 VDD1.n15 2.84303
R189 VDD1.n66 VDD1.n64 2.84303
R190 VDD1.n48 VDD1.n0 2.71565
R191 VDD1.n30 VDD1.n10 2.71565
R192 VDD1.n79 VDD1.n59 2.71565
R193 VDD1.n99 VDD1.n51 2.71565
R194 VDD1.n104 VDD1.t8 2.09796
R195 VDD1.n104 VDD1.t5 2.09796
R196 VDD1.n49 VDD1.t2 2.09796
R197 VDD1.n49 VDD1.t0 2.09796
R198 VDD1.n102 VDD1.t7 2.09796
R199 VDD1.n102 VDD1.t4 2.09796
R200 VDD1.n100 VDD1.t6 2.09796
R201 VDD1.n100 VDD1.t9 2.09796
R202 VDD1.n46 VDD1.n45 1.93989
R203 VDD1.n34 VDD1.n33 1.93989
R204 VDD1.n84 VDD1.n82 1.93989
R205 VDD1.n97 VDD1.n96 1.93989
R206 VDD1.n42 VDD1.n2 1.16414
R207 VDD1.n37 VDD1.n7 1.16414
R208 VDD1.n83 VDD1.n57 1.16414
R209 VDD1.n93 VDD1.n53 1.16414
R210 VDD1 VDD1.n105 0.87981
R211 VDD1.n41 VDD1.n4 0.388379
R212 VDD1.n38 VDD1.n6 0.388379
R213 VDD1.n89 VDD1.n88 0.388379
R214 VDD1.n92 VDD1.n55 0.388379
R215 VDD1 VDD1.n50 0.37119
R216 VDD1.n103 VDD1.n101 0.257654
R217 VDD1.n47 VDD1.n1 0.155672
R218 VDD1.n40 VDD1.n1 0.155672
R219 VDD1.n40 VDD1.n39 0.155672
R220 VDD1.n39 VDD1.n5 0.155672
R221 VDD1.n32 VDD1.n5 0.155672
R222 VDD1.n32 VDD1.n31 0.155672
R223 VDD1.n31 VDD1.n11 0.155672
R224 VDD1.n24 VDD1.n11 0.155672
R225 VDD1.n24 VDD1.n23 0.155672
R226 VDD1.n23 VDD1.n15 0.155672
R227 VDD1.n72 VDD1.n64 0.155672
R228 VDD1.n73 VDD1.n72 0.155672
R229 VDD1.n73 VDD1.n60 0.155672
R230 VDD1.n80 VDD1.n60 0.155672
R231 VDD1.n81 VDD1.n80 0.155672
R232 VDD1.n81 VDD1.n56 0.155672
R233 VDD1.n90 VDD1.n56 0.155672
R234 VDD1.n91 VDD1.n90 0.155672
R235 VDD1.n91 VDD1.n52 0.155672
R236 VDD1.n98 VDD1.n52 0.155672
R237 VTAIL.n208 VTAIL.n164 289.615
R238 VTAIL.n46 VTAIL.n2 289.615
R239 VTAIL.n158 VTAIL.n114 289.615
R240 VTAIL.n104 VTAIL.n60 289.615
R241 VTAIL.n181 VTAIL.n180 185
R242 VTAIL.n183 VTAIL.n182 185
R243 VTAIL.n176 VTAIL.n175 185
R244 VTAIL.n189 VTAIL.n188 185
R245 VTAIL.n191 VTAIL.n190 185
R246 VTAIL.n172 VTAIL.n171 185
R247 VTAIL.n198 VTAIL.n197 185
R248 VTAIL.n199 VTAIL.n170 185
R249 VTAIL.n201 VTAIL.n200 185
R250 VTAIL.n168 VTAIL.n167 185
R251 VTAIL.n207 VTAIL.n206 185
R252 VTAIL.n209 VTAIL.n208 185
R253 VTAIL.n19 VTAIL.n18 185
R254 VTAIL.n21 VTAIL.n20 185
R255 VTAIL.n14 VTAIL.n13 185
R256 VTAIL.n27 VTAIL.n26 185
R257 VTAIL.n29 VTAIL.n28 185
R258 VTAIL.n10 VTAIL.n9 185
R259 VTAIL.n36 VTAIL.n35 185
R260 VTAIL.n37 VTAIL.n8 185
R261 VTAIL.n39 VTAIL.n38 185
R262 VTAIL.n6 VTAIL.n5 185
R263 VTAIL.n45 VTAIL.n44 185
R264 VTAIL.n47 VTAIL.n46 185
R265 VTAIL.n159 VTAIL.n158 185
R266 VTAIL.n157 VTAIL.n156 185
R267 VTAIL.n118 VTAIL.n117 185
R268 VTAIL.n122 VTAIL.n120 185
R269 VTAIL.n151 VTAIL.n150 185
R270 VTAIL.n149 VTAIL.n148 185
R271 VTAIL.n124 VTAIL.n123 185
R272 VTAIL.n143 VTAIL.n142 185
R273 VTAIL.n141 VTAIL.n140 185
R274 VTAIL.n128 VTAIL.n127 185
R275 VTAIL.n135 VTAIL.n134 185
R276 VTAIL.n133 VTAIL.n132 185
R277 VTAIL.n105 VTAIL.n104 185
R278 VTAIL.n103 VTAIL.n102 185
R279 VTAIL.n64 VTAIL.n63 185
R280 VTAIL.n68 VTAIL.n66 185
R281 VTAIL.n97 VTAIL.n96 185
R282 VTAIL.n95 VTAIL.n94 185
R283 VTAIL.n70 VTAIL.n69 185
R284 VTAIL.n89 VTAIL.n88 185
R285 VTAIL.n87 VTAIL.n86 185
R286 VTAIL.n74 VTAIL.n73 185
R287 VTAIL.n81 VTAIL.n80 185
R288 VTAIL.n79 VTAIL.n78 185
R289 VTAIL.n179 VTAIL.t9 149.524
R290 VTAIL.n17 VTAIL.t18 149.524
R291 VTAIL.n131 VTAIL.t15 149.524
R292 VTAIL.n77 VTAIL.t1 149.524
R293 VTAIL.n182 VTAIL.n181 104.615
R294 VTAIL.n182 VTAIL.n175 104.615
R295 VTAIL.n189 VTAIL.n175 104.615
R296 VTAIL.n190 VTAIL.n189 104.615
R297 VTAIL.n190 VTAIL.n171 104.615
R298 VTAIL.n198 VTAIL.n171 104.615
R299 VTAIL.n199 VTAIL.n198 104.615
R300 VTAIL.n200 VTAIL.n199 104.615
R301 VTAIL.n200 VTAIL.n167 104.615
R302 VTAIL.n207 VTAIL.n167 104.615
R303 VTAIL.n208 VTAIL.n207 104.615
R304 VTAIL.n20 VTAIL.n19 104.615
R305 VTAIL.n20 VTAIL.n13 104.615
R306 VTAIL.n27 VTAIL.n13 104.615
R307 VTAIL.n28 VTAIL.n27 104.615
R308 VTAIL.n28 VTAIL.n9 104.615
R309 VTAIL.n36 VTAIL.n9 104.615
R310 VTAIL.n37 VTAIL.n36 104.615
R311 VTAIL.n38 VTAIL.n37 104.615
R312 VTAIL.n38 VTAIL.n5 104.615
R313 VTAIL.n45 VTAIL.n5 104.615
R314 VTAIL.n46 VTAIL.n45 104.615
R315 VTAIL.n158 VTAIL.n157 104.615
R316 VTAIL.n157 VTAIL.n117 104.615
R317 VTAIL.n122 VTAIL.n117 104.615
R318 VTAIL.n150 VTAIL.n122 104.615
R319 VTAIL.n150 VTAIL.n149 104.615
R320 VTAIL.n149 VTAIL.n123 104.615
R321 VTAIL.n142 VTAIL.n123 104.615
R322 VTAIL.n142 VTAIL.n141 104.615
R323 VTAIL.n141 VTAIL.n127 104.615
R324 VTAIL.n134 VTAIL.n127 104.615
R325 VTAIL.n134 VTAIL.n133 104.615
R326 VTAIL.n104 VTAIL.n103 104.615
R327 VTAIL.n103 VTAIL.n63 104.615
R328 VTAIL.n68 VTAIL.n63 104.615
R329 VTAIL.n96 VTAIL.n68 104.615
R330 VTAIL.n96 VTAIL.n95 104.615
R331 VTAIL.n95 VTAIL.n69 104.615
R332 VTAIL.n88 VTAIL.n69 104.615
R333 VTAIL.n88 VTAIL.n87 104.615
R334 VTAIL.n87 VTAIL.n73 104.615
R335 VTAIL.n80 VTAIL.n73 104.615
R336 VTAIL.n80 VTAIL.n79 104.615
R337 VTAIL.n181 VTAIL.t9 52.3082
R338 VTAIL.n19 VTAIL.t18 52.3082
R339 VTAIL.n133 VTAIL.t15 52.3082
R340 VTAIL.n79 VTAIL.t1 52.3082
R341 VTAIL.n113 VTAIL.n112 50.202
R342 VTAIL.n111 VTAIL.n110 50.202
R343 VTAIL.n59 VTAIL.n58 50.202
R344 VTAIL.n57 VTAIL.n56 50.202
R345 VTAIL.n215 VTAIL.n214 50.2019
R346 VTAIL.n1 VTAIL.n0 50.2019
R347 VTAIL.n53 VTAIL.n52 50.2019
R348 VTAIL.n55 VTAIL.n54 50.2019
R349 VTAIL.n213 VTAIL.n212 36.0641
R350 VTAIL.n51 VTAIL.n50 36.0641
R351 VTAIL.n163 VTAIL.n162 36.0641
R352 VTAIL.n109 VTAIL.n108 36.0641
R353 VTAIL.n57 VTAIL.n55 23.0048
R354 VTAIL.n213 VTAIL.n163 21.7548
R355 VTAIL.n201 VTAIL.n168 13.1884
R356 VTAIL.n39 VTAIL.n6 13.1884
R357 VTAIL.n120 VTAIL.n118 13.1884
R358 VTAIL.n66 VTAIL.n64 13.1884
R359 VTAIL.n202 VTAIL.n170 12.8005
R360 VTAIL.n206 VTAIL.n205 12.8005
R361 VTAIL.n40 VTAIL.n8 12.8005
R362 VTAIL.n44 VTAIL.n43 12.8005
R363 VTAIL.n156 VTAIL.n155 12.8005
R364 VTAIL.n152 VTAIL.n151 12.8005
R365 VTAIL.n102 VTAIL.n101 12.8005
R366 VTAIL.n98 VTAIL.n97 12.8005
R367 VTAIL.n197 VTAIL.n196 12.0247
R368 VTAIL.n209 VTAIL.n166 12.0247
R369 VTAIL.n35 VTAIL.n34 12.0247
R370 VTAIL.n47 VTAIL.n4 12.0247
R371 VTAIL.n159 VTAIL.n116 12.0247
R372 VTAIL.n148 VTAIL.n121 12.0247
R373 VTAIL.n105 VTAIL.n62 12.0247
R374 VTAIL.n94 VTAIL.n67 12.0247
R375 VTAIL.n195 VTAIL.n172 11.249
R376 VTAIL.n210 VTAIL.n164 11.249
R377 VTAIL.n33 VTAIL.n10 11.249
R378 VTAIL.n48 VTAIL.n2 11.249
R379 VTAIL.n160 VTAIL.n114 11.249
R380 VTAIL.n147 VTAIL.n124 11.249
R381 VTAIL.n106 VTAIL.n60 11.249
R382 VTAIL.n93 VTAIL.n70 11.249
R383 VTAIL.n192 VTAIL.n191 10.4732
R384 VTAIL.n30 VTAIL.n29 10.4732
R385 VTAIL.n144 VTAIL.n143 10.4732
R386 VTAIL.n90 VTAIL.n89 10.4732
R387 VTAIL.n180 VTAIL.n179 10.2747
R388 VTAIL.n18 VTAIL.n17 10.2747
R389 VTAIL.n132 VTAIL.n131 10.2747
R390 VTAIL.n78 VTAIL.n77 10.2747
R391 VTAIL.n188 VTAIL.n174 9.69747
R392 VTAIL.n26 VTAIL.n12 9.69747
R393 VTAIL.n140 VTAIL.n126 9.69747
R394 VTAIL.n86 VTAIL.n72 9.69747
R395 VTAIL.n212 VTAIL.n211 9.45567
R396 VTAIL.n50 VTAIL.n49 9.45567
R397 VTAIL.n162 VTAIL.n161 9.45567
R398 VTAIL.n108 VTAIL.n107 9.45567
R399 VTAIL.n211 VTAIL.n210 9.3005
R400 VTAIL.n166 VTAIL.n165 9.3005
R401 VTAIL.n205 VTAIL.n204 9.3005
R402 VTAIL.n178 VTAIL.n177 9.3005
R403 VTAIL.n185 VTAIL.n184 9.3005
R404 VTAIL.n187 VTAIL.n186 9.3005
R405 VTAIL.n174 VTAIL.n173 9.3005
R406 VTAIL.n193 VTAIL.n192 9.3005
R407 VTAIL.n195 VTAIL.n194 9.3005
R408 VTAIL.n196 VTAIL.n169 9.3005
R409 VTAIL.n203 VTAIL.n202 9.3005
R410 VTAIL.n49 VTAIL.n48 9.3005
R411 VTAIL.n4 VTAIL.n3 9.3005
R412 VTAIL.n43 VTAIL.n42 9.3005
R413 VTAIL.n16 VTAIL.n15 9.3005
R414 VTAIL.n23 VTAIL.n22 9.3005
R415 VTAIL.n25 VTAIL.n24 9.3005
R416 VTAIL.n12 VTAIL.n11 9.3005
R417 VTAIL.n31 VTAIL.n30 9.3005
R418 VTAIL.n33 VTAIL.n32 9.3005
R419 VTAIL.n34 VTAIL.n7 9.3005
R420 VTAIL.n41 VTAIL.n40 9.3005
R421 VTAIL.n130 VTAIL.n129 9.3005
R422 VTAIL.n137 VTAIL.n136 9.3005
R423 VTAIL.n139 VTAIL.n138 9.3005
R424 VTAIL.n126 VTAIL.n125 9.3005
R425 VTAIL.n145 VTAIL.n144 9.3005
R426 VTAIL.n147 VTAIL.n146 9.3005
R427 VTAIL.n121 VTAIL.n119 9.3005
R428 VTAIL.n153 VTAIL.n152 9.3005
R429 VTAIL.n161 VTAIL.n160 9.3005
R430 VTAIL.n116 VTAIL.n115 9.3005
R431 VTAIL.n155 VTAIL.n154 9.3005
R432 VTAIL.n76 VTAIL.n75 9.3005
R433 VTAIL.n83 VTAIL.n82 9.3005
R434 VTAIL.n85 VTAIL.n84 9.3005
R435 VTAIL.n72 VTAIL.n71 9.3005
R436 VTAIL.n91 VTAIL.n90 9.3005
R437 VTAIL.n93 VTAIL.n92 9.3005
R438 VTAIL.n67 VTAIL.n65 9.3005
R439 VTAIL.n99 VTAIL.n98 9.3005
R440 VTAIL.n107 VTAIL.n106 9.3005
R441 VTAIL.n62 VTAIL.n61 9.3005
R442 VTAIL.n101 VTAIL.n100 9.3005
R443 VTAIL.n187 VTAIL.n176 8.92171
R444 VTAIL.n25 VTAIL.n14 8.92171
R445 VTAIL.n139 VTAIL.n128 8.92171
R446 VTAIL.n85 VTAIL.n74 8.92171
R447 VTAIL.n184 VTAIL.n183 8.14595
R448 VTAIL.n22 VTAIL.n21 8.14595
R449 VTAIL.n136 VTAIL.n135 8.14595
R450 VTAIL.n82 VTAIL.n81 8.14595
R451 VTAIL.n180 VTAIL.n178 7.3702
R452 VTAIL.n18 VTAIL.n16 7.3702
R453 VTAIL.n132 VTAIL.n130 7.3702
R454 VTAIL.n78 VTAIL.n76 7.3702
R455 VTAIL.n183 VTAIL.n178 5.81868
R456 VTAIL.n21 VTAIL.n16 5.81868
R457 VTAIL.n135 VTAIL.n130 5.81868
R458 VTAIL.n81 VTAIL.n76 5.81868
R459 VTAIL.n184 VTAIL.n176 5.04292
R460 VTAIL.n22 VTAIL.n14 5.04292
R461 VTAIL.n136 VTAIL.n128 5.04292
R462 VTAIL.n82 VTAIL.n74 5.04292
R463 VTAIL.n188 VTAIL.n187 4.26717
R464 VTAIL.n26 VTAIL.n25 4.26717
R465 VTAIL.n140 VTAIL.n139 4.26717
R466 VTAIL.n86 VTAIL.n85 4.26717
R467 VTAIL.n191 VTAIL.n174 3.49141
R468 VTAIL.n29 VTAIL.n12 3.49141
R469 VTAIL.n143 VTAIL.n126 3.49141
R470 VTAIL.n89 VTAIL.n72 3.49141
R471 VTAIL.n179 VTAIL.n177 2.84303
R472 VTAIL.n17 VTAIL.n15 2.84303
R473 VTAIL.n131 VTAIL.n129 2.84303
R474 VTAIL.n77 VTAIL.n75 2.84303
R475 VTAIL.n192 VTAIL.n172 2.71565
R476 VTAIL.n212 VTAIL.n164 2.71565
R477 VTAIL.n30 VTAIL.n10 2.71565
R478 VTAIL.n50 VTAIL.n2 2.71565
R479 VTAIL.n162 VTAIL.n114 2.71565
R480 VTAIL.n144 VTAIL.n124 2.71565
R481 VTAIL.n108 VTAIL.n60 2.71565
R482 VTAIL.n90 VTAIL.n70 2.71565
R483 VTAIL.n214 VTAIL.t2 2.09796
R484 VTAIL.n214 VTAIL.t5 2.09796
R485 VTAIL.n0 VTAIL.t6 2.09796
R486 VTAIL.n0 VTAIL.t7 2.09796
R487 VTAIL.n52 VTAIL.t10 2.09796
R488 VTAIL.n52 VTAIL.t19 2.09796
R489 VTAIL.n54 VTAIL.t13 2.09796
R490 VTAIL.n54 VTAIL.t12 2.09796
R491 VTAIL.n112 VTAIL.t11 2.09796
R492 VTAIL.n112 VTAIL.t17 2.09796
R493 VTAIL.n110 VTAIL.t16 2.09796
R494 VTAIL.n110 VTAIL.t14 2.09796
R495 VTAIL.n58 VTAIL.t3 2.09796
R496 VTAIL.n58 VTAIL.t8 2.09796
R497 VTAIL.n56 VTAIL.t0 2.09796
R498 VTAIL.n56 VTAIL.t4 2.09796
R499 VTAIL.n197 VTAIL.n195 1.93989
R500 VTAIL.n210 VTAIL.n209 1.93989
R501 VTAIL.n35 VTAIL.n33 1.93989
R502 VTAIL.n48 VTAIL.n47 1.93989
R503 VTAIL.n160 VTAIL.n159 1.93989
R504 VTAIL.n148 VTAIL.n147 1.93989
R505 VTAIL.n106 VTAIL.n105 1.93989
R506 VTAIL.n94 VTAIL.n93 1.93989
R507 VTAIL.n59 VTAIL.n57 1.2505
R508 VTAIL.n109 VTAIL.n59 1.2505
R509 VTAIL.n113 VTAIL.n111 1.2505
R510 VTAIL.n163 VTAIL.n113 1.2505
R511 VTAIL.n55 VTAIL.n53 1.2505
R512 VTAIL.n53 VTAIL.n51 1.2505
R513 VTAIL.n215 VTAIL.n213 1.2505
R514 VTAIL.n196 VTAIL.n170 1.16414
R515 VTAIL.n206 VTAIL.n166 1.16414
R516 VTAIL.n34 VTAIL.n8 1.16414
R517 VTAIL.n44 VTAIL.n4 1.16414
R518 VTAIL.n156 VTAIL.n116 1.16414
R519 VTAIL.n151 VTAIL.n121 1.16414
R520 VTAIL.n102 VTAIL.n62 1.16414
R521 VTAIL.n97 VTAIL.n67 1.16414
R522 VTAIL.n111 VTAIL.n109 1.09533
R523 VTAIL.n51 VTAIL.n1 1.09533
R524 VTAIL VTAIL.n1 0.99619
R525 VTAIL.n202 VTAIL.n201 0.388379
R526 VTAIL.n205 VTAIL.n168 0.388379
R527 VTAIL.n40 VTAIL.n39 0.388379
R528 VTAIL.n43 VTAIL.n6 0.388379
R529 VTAIL.n155 VTAIL.n118 0.388379
R530 VTAIL.n152 VTAIL.n120 0.388379
R531 VTAIL.n101 VTAIL.n64 0.388379
R532 VTAIL.n98 VTAIL.n66 0.388379
R533 VTAIL VTAIL.n215 0.25481
R534 VTAIL.n185 VTAIL.n177 0.155672
R535 VTAIL.n186 VTAIL.n185 0.155672
R536 VTAIL.n186 VTAIL.n173 0.155672
R537 VTAIL.n193 VTAIL.n173 0.155672
R538 VTAIL.n194 VTAIL.n193 0.155672
R539 VTAIL.n194 VTAIL.n169 0.155672
R540 VTAIL.n203 VTAIL.n169 0.155672
R541 VTAIL.n204 VTAIL.n203 0.155672
R542 VTAIL.n204 VTAIL.n165 0.155672
R543 VTAIL.n211 VTAIL.n165 0.155672
R544 VTAIL.n23 VTAIL.n15 0.155672
R545 VTAIL.n24 VTAIL.n23 0.155672
R546 VTAIL.n24 VTAIL.n11 0.155672
R547 VTAIL.n31 VTAIL.n11 0.155672
R548 VTAIL.n32 VTAIL.n31 0.155672
R549 VTAIL.n32 VTAIL.n7 0.155672
R550 VTAIL.n41 VTAIL.n7 0.155672
R551 VTAIL.n42 VTAIL.n41 0.155672
R552 VTAIL.n42 VTAIL.n3 0.155672
R553 VTAIL.n49 VTAIL.n3 0.155672
R554 VTAIL.n161 VTAIL.n115 0.155672
R555 VTAIL.n154 VTAIL.n115 0.155672
R556 VTAIL.n154 VTAIL.n153 0.155672
R557 VTAIL.n153 VTAIL.n119 0.155672
R558 VTAIL.n146 VTAIL.n119 0.155672
R559 VTAIL.n146 VTAIL.n145 0.155672
R560 VTAIL.n145 VTAIL.n125 0.155672
R561 VTAIL.n138 VTAIL.n125 0.155672
R562 VTAIL.n138 VTAIL.n137 0.155672
R563 VTAIL.n137 VTAIL.n129 0.155672
R564 VTAIL.n107 VTAIL.n61 0.155672
R565 VTAIL.n100 VTAIL.n61 0.155672
R566 VTAIL.n100 VTAIL.n99 0.155672
R567 VTAIL.n99 VTAIL.n65 0.155672
R568 VTAIL.n92 VTAIL.n65 0.155672
R569 VTAIL.n92 VTAIL.n91 0.155672
R570 VTAIL.n91 VTAIL.n71 0.155672
R571 VTAIL.n84 VTAIL.n71 0.155672
R572 VTAIL.n84 VTAIL.n83 0.155672
R573 VTAIL.n83 VTAIL.n75 0.155672
R574 B.n670 B.n669 585
R575 B.n260 B.n101 585
R576 B.n259 B.n258 585
R577 B.n257 B.n256 585
R578 B.n255 B.n254 585
R579 B.n253 B.n252 585
R580 B.n251 B.n250 585
R581 B.n249 B.n248 585
R582 B.n247 B.n246 585
R583 B.n245 B.n244 585
R584 B.n243 B.n242 585
R585 B.n241 B.n240 585
R586 B.n239 B.n238 585
R587 B.n237 B.n236 585
R588 B.n235 B.n234 585
R589 B.n233 B.n232 585
R590 B.n231 B.n230 585
R591 B.n229 B.n228 585
R592 B.n227 B.n226 585
R593 B.n225 B.n224 585
R594 B.n223 B.n222 585
R595 B.n221 B.n220 585
R596 B.n219 B.n218 585
R597 B.n217 B.n216 585
R598 B.n215 B.n214 585
R599 B.n213 B.n212 585
R600 B.n211 B.n210 585
R601 B.n209 B.n208 585
R602 B.n207 B.n206 585
R603 B.n205 B.n204 585
R604 B.n203 B.n202 585
R605 B.n201 B.n200 585
R606 B.n199 B.n198 585
R607 B.n197 B.n196 585
R608 B.n195 B.n194 585
R609 B.n193 B.n192 585
R610 B.n191 B.n190 585
R611 B.n189 B.n188 585
R612 B.n187 B.n186 585
R613 B.n185 B.n184 585
R614 B.n183 B.n182 585
R615 B.n181 B.n180 585
R616 B.n179 B.n178 585
R617 B.n177 B.n176 585
R618 B.n175 B.n174 585
R619 B.n173 B.n172 585
R620 B.n171 B.n170 585
R621 B.n169 B.n168 585
R622 B.n167 B.n166 585
R623 B.n165 B.n164 585
R624 B.n163 B.n162 585
R625 B.n161 B.n160 585
R626 B.n159 B.n158 585
R627 B.n157 B.n156 585
R628 B.n155 B.n154 585
R629 B.n153 B.n152 585
R630 B.n151 B.n150 585
R631 B.n149 B.n148 585
R632 B.n147 B.n146 585
R633 B.n145 B.n144 585
R634 B.n143 B.n142 585
R635 B.n141 B.n140 585
R636 B.n139 B.n138 585
R637 B.n137 B.n136 585
R638 B.n135 B.n134 585
R639 B.n133 B.n132 585
R640 B.n131 B.n130 585
R641 B.n129 B.n128 585
R642 B.n127 B.n126 585
R643 B.n125 B.n124 585
R644 B.n123 B.n122 585
R645 B.n121 B.n120 585
R646 B.n119 B.n118 585
R647 B.n117 B.n116 585
R648 B.n115 B.n114 585
R649 B.n113 B.n112 585
R650 B.n111 B.n110 585
R651 B.n109 B.n108 585
R652 B.n668 B.n62 585
R653 B.n673 B.n62 585
R654 B.n667 B.n61 585
R655 B.n674 B.n61 585
R656 B.n666 B.n665 585
R657 B.n665 B.n57 585
R658 B.n664 B.n56 585
R659 B.n680 B.n56 585
R660 B.n663 B.n55 585
R661 B.n681 B.n55 585
R662 B.n662 B.n54 585
R663 B.n682 B.n54 585
R664 B.n661 B.n660 585
R665 B.n660 B.n50 585
R666 B.n659 B.n49 585
R667 B.n688 B.n49 585
R668 B.n658 B.n48 585
R669 B.n689 B.n48 585
R670 B.n657 B.n47 585
R671 B.n690 B.n47 585
R672 B.n656 B.n655 585
R673 B.n655 B.n43 585
R674 B.n654 B.n42 585
R675 B.n696 B.n42 585
R676 B.n653 B.n41 585
R677 B.n697 B.n41 585
R678 B.n652 B.n40 585
R679 B.n698 B.n40 585
R680 B.n651 B.n650 585
R681 B.n650 B.n36 585
R682 B.n649 B.n35 585
R683 B.n704 B.n35 585
R684 B.n648 B.n34 585
R685 B.n705 B.n34 585
R686 B.n647 B.n33 585
R687 B.n706 B.n33 585
R688 B.n646 B.n645 585
R689 B.n645 B.n29 585
R690 B.n644 B.n28 585
R691 B.n712 B.n28 585
R692 B.n643 B.n27 585
R693 B.n713 B.n27 585
R694 B.n642 B.n26 585
R695 B.n714 B.n26 585
R696 B.n641 B.n640 585
R697 B.n640 B.n22 585
R698 B.n639 B.n21 585
R699 B.n720 B.n21 585
R700 B.n638 B.n20 585
R701 B.n721 B.n20 585
R702 B.n637 B.n19 585
R703 B.n722 B.n19 585
R704 B.n636 B.n635 585
R705 B.n635 B.n15 585
R706 B.n634 B.n14 585
R707 B.n728 B.n14 585
R708 B.n633 B.n13 585
R709 B.n729 B.n13 585
R710 B.n632 B.n12 585
R711 B.n730 B.n12 585
R712 B.n631 B.n630 585
R713 B.n630 B.n629 585
R714 B.n628 B.n627 585
R715 B.n628 B.n8 585
R716 B.n626 B.n7 585
R717 B.n737 B.n7 585
R718 B.n625 B.n6 585
R719 B.n738 B.n6 585
R720 B.n624 B.n5 585
R721 B.n739 B.n5 585
R722 B.n623 B.n622 585
R723 B.n622 B.n4 585
R724 B.n621 B.n261 585
R725 B.n621 B.n620 585
R726 B.n611 B.n262 585
R727 B.n263 B.n262 585
R728 B.n613 B.n612 585
R729 B.n614 B.n613 585
R730 B.n610 B.n268 585
R731 B.n268 B.n267 585
R732 B.n609 B.n608 585
R733 B.n608 B.n607 585
R734 B.n270 B.n269 585
R735 B.n271 B.n270 585
R736 B.n600 B.n599 585
R737 B.n601 B.n600 585
R738 B.n598 B.n276 585
R739 B.n276 B.n275 585
R740 B.n597 B.n596 585
R741 B.n596 B.n595 585
R742 B.n278 B.n277 585
R743 B.n279 B.n278 585
R744 B.n588 B.n587 585
R745 B.n589 B.n588 585
R746 B.n586 B.n284 585
R747 B.n284 B.n283 585
R748 B.n585 B.n584 585
R749 B.n584 B.n583 585
R750 B.n286 B.n285 585
R751 B.n287 B.n286 585
R752 B.n576 B.n575 585
R753 B.n577 B.n576 585
R754 B.n574 B.n291 585
R755 B.n295 B.n291 585
R756 B.n573 B.n572 585
R757 B.n572 B.n571 585
R758 B.n293 B.n292 585
R759 B.n294 B.n293 585
R760 B.n564 B.n563 585
R761 B.n565 B.n564 585
R762 B.n562 B.n299 585
R763 B.n303 B.n299 585
R764 B.n561 B.n560 585
R765 B.n560 B.n559 585
R766 B.n301 B.n300 585
R767 B.n302 B.n301 585
R768 B.n552 B.n551 585
R769 B.n553 B.n552 585
R770 B.n550 B.n308 585
R771 B.n308 B.n307 585
R772 B.n549 B.n548 585
R773 B.n548 B.n547 585
R774 B.n310 B.n309 585
R775 B.n311 B.n310 585
R776 B.n540 B.n539 585
R777 B.n541 B.n540 585
R778 B.n538 B.n316 585
R779 B.n316 B.n315 585
R780 B.n537 B.n536 585
R781 B.n536 B.n535 585
R782 B.n318 B.n317 585
R783 B.n319 B.n318 585
R784 B.n528 B.n527 585
R785 B.n529 B.n528 585
R786 B.n526 B.n324 585
R787 B.n324 B.n323 585
R788 B.n521 B.n520 585
R789 B.n519 B.n365 585
R790 B.n518 B.n364 585
R791 B.n523 B.n364 585
R792 B.n517 B.n516 585
R793 B.n515 B.n514 585
R794 B.n513 B.n512 585
R795 B.n511 B.n510 585
R796 B.n509 B.n508 585
R797 B.n507 B.n506 585
R798 B.n505 B.n504 585
R799 B.n503 B.n502 585
R800 B.n501 B.n500 585
R801 B.n499 B.n498 585
R802 B.n497 B.n496 585
R803 B.n495 B.n494 585
R804 B.n493 B.n492 585
R805 B.n491 B.n490 585
R806 B.n489 B.n488 585
R807 B.n487 B.n486 585
R808 B.n485 B.n484 585
R809 B.n483 B.n482 585
R810 B.n481 B.n480 585
R811 B.n479 B.n478 585
R812 B.n477 B.n476 585
R813 B.n475 B.n474 585
R814 B.n473 B.n472 585
R815 B.n471 B.n470 585
R816 B.n469 B.n468 585
R817 B.n467 B.n466 585
R818 B.n465 B.n464 585
R819 B.n463 B.n462 585
R820 B.n461 B.n460 585
R821 B.n459 B.n458 585
R822 B.n457 B.n456 585
R823 B.n454 B.n453 585
R824 B.n452 B.n451 585
R825 B.n450 B.n449 585
R826 B.n448 B.n447 585
R827 B.n446 B.n445 585
R828 B.n444 B.n443 585
R829 B.n442 B.n441 585
R830 B.n440 B.n439 585
R831 B.n438 B.n437 585
R832 B.n436 B.n435 585
R833 B.n433 B.n432 585
R834 B.n431 B.n430 585
R835 B.n429 B.n428 585
R836 B.n427 B.n426 585
R837 B.n425 B.n424 585
R838 B.n423 B.n422 585
R839 B.n421 B.n420 585
R840 B.n419 B.n418 585
R841 B.n417 B.n416 585
R842 B.n415 B.n414 585
R843 B.n413 B.n412 585
R844 B.n411 B.n410 585
R845 B.n409 B.n408 585
R846 B.n407 B.n406 585
R847 B.n405 B.n404 585
R848 B.n403 B.n402 585
R849 B.n401 B.n400 585
R850 B.n399 B.n398 585
R851 B.n397 B.n396 585
R852 B.n395 B.n394 585
R853 B.n393 B.n392 585
R854 B.n391 B.n390 585
R855 B.n389 B.n388 585
R856 B.n387 B.n386 585
R857 B.n385 B.n384 585
R858 B.n383 B.n382 585
R859 B.n381 B.n380 585
R860 B.n379 B.n378 585
R861 B.n377 B.n376 585
R862 B.n375 B.n374 585
R863 B.n373 B.n372 585
R864 B.n371 B.n370 585
R865 B.n326 B.n325 585
R866 B.n525 B.n524 585
R867 B.n524 B.n523 585
R868 B.n322 B.n321 585
R869 B.n323 B.n322 585
R870 B.n531 B.n530 585
R871 B.n530 B.n529 585
R872 B.n532 B.n320 585
R873 B.n320 B.n319 585
R874 B.n534 B.n533 585
R875 B.n535 B.n534 585
R876 B.n314 B.n313 585
R877 B.n315 B.n314 585
R878 B.n543 B.n542 585
R879 B.n542 B.n541 585
R880 B.n544 B.n312 585
R881 B.n312 B.n311 585
R882 B.n546 B.n545 585
R883 B.n547 B.n546 585
R884 B.n306 B.n305 585
R885 B.n307 B.n306 585
R886 B.n555 B.n554 585
R887 B.n554 B.n553 585
R888 B.n556 B.n304 585
R889 B.n304 B.n302 585
R890 B.n558 B.n557 585
R891 B.n559 B.n558 585
R892 B.n298 B.n297 585
R893 B.n303 B.n298 585
R894 B.n567 B.n566 585
R895 B.n566 B.n565 585
R896 B.n568 B.n296 585
R897 B.n296 B.n294 585
R898 B.n570 B.n569 585
R899 B.n571 B.n570 585
R900 B.n290 B.n289 585
R901 B.n295 B.n290 585
R902 B.n579 B.n578 585
R903 B.n578 B.n577 585
R904 B.n580 B.n288 585
R905 B.n288 B.n287 585
R906 B.n582 B.n581 585
R907 B.n583 B.n582 585
R908 B.n282 B.n281 585
R909 B.n283 B.n282 585
R910 B.n591 B.n590 585
R911 B.n590 B.n589 585
R912 B.n592 B.n280 585
R913 B.n280 B.n279 585
R914 B.n594 B.n593 585
R915 B.n595 B.n594 585
R916 B.n274 B.n273 585
R917 B.n275 B.n274 585
R918 B.n603 B.n602 585
R919 B.n602 B.n601 585
R920 B.n604 B.n272 585
R921 B.n272 B.n271 585
R922 B.n606 B.n605 585
R923 B.n607 B.n606 585
R924 B.n266 B.n265 585
R925 B.n267 B.n266 585
R926 B.n616 B.n615 585
R927 B.n615 B.n614 585
R928 B.n617 B.n264 585
R929 B.n264 B.n263 585
R930 B.n619 B.n618 585
R931 B.n620 B.n619 585
R932 B.n3 B.n0 585
R933 B.n4 B.n3 585
R934 B.n736 B.n1 585
R935 B.n737 B.n736 585
R936 B.n735 B.n734 585
R937 B.n735 B.n8 585
R938 B.n733 B.n9 585
R939 B.n629 B.n9 585
R940 B.n732 B.n731 585
R941 B.n731 B.n730 585
R942 B.n11 B.n10 585
R943 B.n729 B.n11 585
R944 B.n727 B.n726 585
R945 B.n728 B.n727 585
R946 B.n725 B.n16 585
R947 B.n16 B.n15 585
R948 B.n724 B.n723 585
R949 B.n723 B.n722 585
R950 B.n18 B.n17 585
R951 B.n721 B.n18 585
R952 B.n719 B.n718 585
R953 B.n720 B.n719 585
R954 B.n717 B.n23 585
R955 B.n23 B.n22 585
R956 B.n716 B.n715 585
R957 B.n715 B.n714 585
R958 B.n25 B.n24 585
R959 B.n713 B.n25 585
R960 B.n711 B.n710 585
R961 B.n712 B.n711 585
R962 B.n709 B.n30 585
R963 B.n30 B.n29 585
R964 B.n708 B.n707 585
R965 B.n707 B.n706 585
R966 B.n32 B.n31 585
R967 B.n705 B.n32 585
R968 B.n703 B.n702 585
R969 B.n704 B.n703 585
R970 B.n701 B.n37 585
R971 B.n37 B.n36 585
R972 B.n700 B.n699 585
R973 B.n699 B.n698 585
R974 B.n39 B.n38 585
R975 B.n697 B.n39 585
R976 B.n695 B.n694 585
R977 B.n696 B.n695 585
R978 B.n693 B.n44 585
R979 B.n44 B.n43 585
R980 B.n692 B.n691 585
R981 B.n691 B.n690 585
R982 B.n46 B.n45 585
R983 B.n689 B.n46 585
R984 B.n687 B.n686 585
R985 B.n688 B.n687 585
R986 B.n685 B.n51 585
R987 B.n51 B.n50 585
R988 B.n684 B.n683 585
R989 B.n683 B.n682 585
R990 B.n53 B.n52 585
R991 B.n681 B.n53 585
R992 B.n679 B.n678 585
R993 B.n680 B.n679 585
R994 B.n677 B.n58 585
R995 B.n58 B.n57 585
R996 B.n676 B.n675 585
R997 B.n675 B.n674 585
R998 B.n60 B.n59 585
R999 B.n673 B.n60 585
R1000 B.n740 B.n739 585
R1001 B.n738 B.n2 585
R1002 B.n108 B.n60 511.721
R1003 B.n670 B.n62 511.721
R1004 B.n524 B.n324 511.721
R1005 B.n521 B.n322 511.721
R1006 B.n105 B.t18 406.807
R1007 B.n102 B.t14 406.807
R1008 B.n368 B.t10 406.807
R1009 B.n366 B.t21 406.807
R1010 B.n102 B.t16 266.384
R1011 B.n368 B.t13 266.384
R1012 B.n105 B.t19 266.384
R1013 B.n366 B.t23 266.384
R1014 B.n672 B.n671 256.663
R1015 B.n672 B.n100 256.663
R1016 B.n672 B.n99 256.663
R1017 B.n672 B.n98 256.663
R1018 B.n672 B.n97 256.663
R1019 B.n672 B.n96 256.663
R1020 B.n672 B.n95 256.663
R1021 B.n672 B.n94 256.663
R1022 B.n672 B.n93 256.663
R1023 B.n672 B.n92 256.663
R1024 B.n672 B.n91 256.663
R1025 B.n672 B.n90 256.663
R1026 B.n672 B.n89 256.663
R1027 B.n672 B.n88 256.663
R1028 B.n672 B.n87 256.663
R1029 B.n672 B.n86 256.663
R1030 B.n672 B.n85 256.663
R1031 B.n672 B.n84 256.663
R1032 B.n672 B.n83 256.663
R1033 B.n672 B.n82 256.663
R1034 B.n672 B.n81 256.663
R1035 B.n672 B.n80 256.663
R1036 B.n672 B.n79 256.663
R1037 B.n672 B.n78 256.663
R1038 B.n672 B.n77 256.663
R1039 B.n672 B.n76 256.663
R1040 B.n672 B.n75 256.663
R1041 B.n672 B.n74 256.663
R1042 B.n672 B.n73 256.663
R1043 B.n672 B.n72 256.663
R1044 B.n672 B.n71 256.663
R1045 B.n672 B.n70 256.663
R1046 B.n672 B.n69 256.663
R1047 B.n672 B.n68 256.663
R1048 B.n672 B.n67 256.663
R1049 B.n672 B.n66 256.663
R1050 B.n672 B.n65 256.663
R1051 B.n672 B.n64 256.663
R1052 B.n672 B.n63 256.663
R1053 B.n523 B.n522 256.663
R1054 B.n523 B.n327 256.663
R1055 B.n523 B.n328 256.663
R1056 B.n523 B.n329 256.663
R1057 B.n523 B.n330 256.663
R1058 B.n523 B.n331 256.663
R1059 B.n523 B.n332 256.663
R1060 B.n523 B.n333 256.663
R1061 B.n523 B.n334 256.663
R1062 B.n523 B.n335 256.663
R1063 B.n523 B.n336 256.663
R1064 B.n523 B.n337 256.663
R1065 B.n523 B.n338 256.663
R1066 B.n523 B.n339 256.663
R1067 B.n523 B.n340 256.663
R1068 B.n523 B.n341 256.663
R1069 B.n523 B.n342 256.663
R1070 B.n523 B.n343 256.663
R1071 B.n523 B.n344 256.663
R1072 B.n523 B.n345 256.663
R1073 B.n523 B.n346 256.663
R1074 B.n523 B.n347 256.663
R1075 B.n523 B.n348 256.663
R1076 B.n523 B.n349 256.663
R1077 B.n523 B.n350 256.663
R1078 B.n523 B.n351 256.663
R1079 B.n523 B.n352 256.663
R1080 B.n523 B.n353 256.663
R1081 B.n523 B.n354 256.663
R1082 B.n523 B.n355 256.663
R1083 B.n523 B.n356 256.663
R1084 B.n523 B.n357 256.663
R1085 B.n523 B.n358 256.663
R1086 B.n523 B.n359 256.663
R1087 B.n523 B.n360 256.663
R1088 B.n523 B.n361 256.663
R1089 B.n523 B.n362 256.663
R1090 B.n523 B.n363 256.663
R1091 B.n742 B.n741 256.663
R1092 B.n103 B.t17 238.262
R1093 B.n369 B.t12 238.262
R1094 B.n106 B.t20 238.262
R1095 B.n367 B.t22 238.262
R1096 B.n112 B.n111 163.367
R1097 B.n116 B.n115 163.367
R1098 B.n120 B.n119 163.367
R1099 B.n124 B.n123 163.367
R1100 B.n128 B.n127 163.367
R1101 B.n132 B.n131 163.367
R1102 B.n136 B.n135 163.367
R1103 B.n140 B.n139 163.367
R1104 B.n144 B.n143 163.367
R1105 B.n148 B.n147 163.367
R1106 B.n152 B.n151 163.367
R1107 B.n156 B.n155 163.367
R1108 B.n160 B.n159 163.367
R1109 B.n164 B.n163 163.367
R1110 B.n168 B.n167 163.367
R1111 B.n172 B.n171 163.367
R1112 B.n176 B.n175 163.367
R1113 B.n180 B.n179 163.367
R1114 B.n184 B.n183 163.367
R1115 B.n188 B.n187 163.367
R1116 B.n192 B.n191 163.367
R1117 B.n196 B.n195 163.367
R1118 B.n200 B.n199 163.367
R1119 B.n204 B.n203 163.367
R1120 B.n208 B.n207 163.367
R1121 B.n212 B.n211 163.367
R1122 B.n216 B.n215 163.367
R1123 B.n220 B.n219 163.367
R1124 B.n224 B.n223 163.367
R1125 B.n228 B.n227 163.367
R1126 B.n232 B.n231 163.367
R1127 B.n236 B.n235 163.367
R1128 B.n240 B.n239 163.367
R1129 B.n244 B.n243 163.367
R1130 B.n248 B.n247 163.367
R1131 B.n252 B.n251 163.367
R1132 B.n256 B.n255 163.367
R1133 B.n258 B.n101 163.367
R1134 B.n528 B.n324 163.367
R1135 B.n528 B.n318 163.367
R1136 B.n536 B.n318 163.367
R1137 B.n536 B.n316 163.367
R1138 B.n540 B.n316 163.367
R1139 B.n540 B.n310 163.367
R1140 B.n548 B.n310 163.367
R1141 B.n548 B.n308 163.367
R1142 B.n552 B.n308 163.367
R1143 B.n552 B.n301 163.367
R1144 B.n560 B.n301 163.367
R1145 B.n560 B.n299 163.367
R1146 B.n564 B.n299 163.367
R1147 B.n564 B.n293 163.367
R1148 B.n572 B.n293 163.367
R1149 B.n572 B.n291 163.367
R1150 B.n576 B.n291 163.367
R1151 B.n576 B.n286 163.367
R1152 B.n584 B.n286 163.367
R1153 B.n584 B.n284 163.367
R1154 B.n588 B.n284 163.367
R1155 B.n588 B.n278 163.367
R1156 B.n596 B.n278 163.367
R1157 B.n596 B.n276 163.367
R1158 B.n600 B.n276 163.367
R1159 B.n600 B.n270 163.367
R1160 B.n608 B.n270 163.367
R1161 B.n608 B.n268 163.367
R1162 B.n613 B.n268 163.367
R1163 B.n613 B.n262 163.367
R1164 B.n621 B.n262 163.367
R1165 B.n622 B.n621 163.367
R1166 B.n622 B.n5 163.367
R1167 B.n6 B.n5 163.367
R1168 B.n7 B.n6 163.367
R1169 B.n628 B.n7 163.367
R1170 B.n630 B.n628 163.367
R1171 B.n630 B.n12 163.367
R1172 B.n13 B.n12 163.367
R1173 B.n14 B.n13 163.367
R1174 B.n635 B.n14 163.367
R1175 B.n635 B.n19 163.367
R1176 B.n20 B.n19 163.367
R1177 B.n21 B.n20 163.367
R1178 B.n640 B.n21 163.367
R1179 B.n640 B.n26 163.367
R1180 B.n27 B.n26 163.367
R1181 B.n28 B.n27 163.367
R1182 B.n645 B.n28 163.367
R1183 B.n645 B.n33 163.367
R1184 B.n34 B.n33 163.367
R1185 B.n35 B.n34 163.367
R1186 B.n650 B.n35 163.367
R1187 B.n650 B.n40 163.367
R1188 B.n41 B.n40 163.367
R1189 B.n42 B.n41 163.367
R1190 B.n655 B.n42 163.367
R1191 B.n655 B.n47 163.367
R1192 B.n48 B.n47 163.367
R1193 B.n49 B.n48 163.367
R1194 B.n660 B.n49 163.367
R1195 B.n660 B.n54 163.367
R1196 B.n55 B.n54 163.367
R1197 B.n56 B.n55 163.367
R1198 B.n665 B.n56 163.367
R1199 B.n665 B.n61 163.367
R1200 B.n62 B.n61 163.367
R1201 B.n365 B.n364 163.367
R1202 B.n516 B.n364 163.367
R1203 B.n514 B.n513 163.367
R1204 B.n510 B.n509 163.367
R1205 B.n506 B.n505 163.367
R1206 B.n502 B.n501 163.367
R1207 B.n498 B.n497 163.367
R1208 B.n494 B.n493 163.367
R1209 B.n490 B.n489 163.367
R1210 B.n486 B.n485 163.367
R1211 B.n482 B.n481 163.367
R1212 B.n478 B.n477 163.367
R1213 B.n474 B.n473 163.367
R1214 B.n470 B.n469 163.367
R1215 B.n466 B.n465 163.367
R1216 B.n462 B.n461 163.367
R1217 B.n458 B.n457 163.367
R1218 B.n453 B.n452 163.367
R1219 B.n449 B.n448 163.367
R1220 B.n445 B.n444 163.367
R1221 B.n441 B.n440 163.367
R1222 B.n437 B.n436 163.367
R1223 B.n432 B.n431 163.367
R1224 B.n428 B.n427 163.367
R1225 B.n424 B.n423 163.367
R1226 B.n420 B.n419 163.367
R1227 B.n416 B.n415 163.367
R1228 B.n412 B.n411 163.367
R1229 B.n408 B.n407 163.367
R1230 B.n404 B.n403 163.367
R1231 B.n400 B.n399 163.367
R1232 B.n396 B.n395 163.367
R1233 B.n392 B.n391 163.367
R1234 B.n388 B.n387 163.367
R1235 B.n384 B.n383 163.367
R1236 B.n380 B.n379 163.367
R1237 B.n376 B.n375 163.367
R1238 B.n372 B.n371 163.367
R1239 B.n524 B.n326 163.367
R1240 B.n530 B.n322 163.367
R1241 B.n530 B.n320 163.367
R1242 B.n534 B.n320 163.367
R1243 B.n534 B.n314 163.367
R1244 B.n542 B.n314 163.367
R1245 B.n542 B.n312 163.367
R1246 B.n546 B.n312 163.367
R1247 B.n546 B.n306 163.367
R1248 B.n554 B.n306 163.367
R1249 B.n554 B.n304 163.367
R1250 B.n558 B.n304 163.367
R1251 B.n558 B.n298 163.367
R1252 B.n566 B.n298 163.367
R1253 B.n566 B.n296 163.367
R1254 B.n570 B.n296 163.367
R1255 B.n570 B.n290 163.367
R1256 B.n578 B.n290 163.367
R1257 B.n578 B.n288 163.367
R1258 B.n582 B.n288 163.367
R1259 B.n582 B.n282 163.367
R1260 B.n590 B.n282 163.367
R1261 B.n590 B.n280 163.367
R1262 B.n594 B.n280 163.367
R1263 B.n594 B.n274 163.367
R1264 B.n602 B.n274 163.367
R1265 B.n602 B.n272 163.367
R1266 B.n606 B.n272 163.367
R1267 B.n606 B.n266 163.367
R1268 B.n615 B.n266 163.367
R1269 B.n615 B.n264 163.367
R1270 B.n619 B.n264 163.367
R1271 B.n619 B.n3 163.367
R1272 B.n740 B.n3 163.367
R1273 B.n736 B.n2 163.367
R1274 B.n736 B.n735 163.367
R1275 B.n735 B.n9 163.367
R1276 B.n731 B.n9 163.367
R1277 B.n731 B.n11 163.367
R1278 B.n727 B.n11 163.367
R1279 B.n727 B.n16 163.367
R1280 B.n723 B.n16 163.367
R1281 B.n723 B.n18 163.367
R1282 B.n719 B.n18 163.367
R1283 B.n719 B.n23 163.367
R1284 B.n715 B.n23 163.367
R1285 B.n715 B.n25 163.367
R1286 B.n711 B.n25 163.367
R1287 B.n711 B.n30 163.367
R1288 B.n707 B.n30 163.367
R1289 B.n707 B.n32 163.367
R1290 B.n703 B.n32 163.367
R1291 B.n703 B.n37 163.367
R1292 B.n699 B.n37 163.367
R1293 B.n699 B.n39 163.367
R1294 B.n695 B.n39 163.367
R1295 B.n695 B.n44 163.367
R1296 B.n691 B.n44 163.367
R1297 B.n691 B.n46 163.367
R1298 B.n687 B.n46 163.367
R1299 B.n687 B.n51 163.367
R1300 B.n683 B.n51 163.367
R1301 B.n683 B.n53 163.367
R1302 B.n679 B.n53 163.367
R1303 B.n679 B.n58 163.367
R1304 B.n675 B.n58 163.367
R1305 B.n675 B.n60 163.367
R1306 B.n523 B.n323 102.413
R1307 B.n673 B.n672 102.413
R1308 B.n108 B.n63 71.676
R1309 B.n112 B.n64 71.676
R1310 B.n116 B.n65 71.676
R1311 B.n120 B.n66 71.676
R1312 B.n124 B.n67 71.676
R1313 B.n128 B.n68 71.676
R1314 B.n132 B.n69 71.676
R1315 B.n136 B.n70 71.676
R1316 B.n140 B.n71 71.676
R1317 B.n144 B.n72 71.676
R1318 B.n148 B.n73 71.676
R1319 B.n152 B.n74 71.676
R1320 B.n156 B.n75 71.676
R1321 B.n160 B.n76 71.676
R1322 B.n164 B.n77 71.676
R1323 B.n168 B.n78 71.676
R1324 B.n172 B.n79 71.676
R1325 B.n176 B.n80 71.676
R1326 B.n180 B.n81 71.676
R1327 B.n184 B.n82 71.676
R1328 B.n188 B.n83 71.676
R1329 B.n192 B.n84 71.676
R1330 B.n196 B.n85 71.676
R1331 B.n200 B.n86 71.676
R1332 B.n204 B.n87 71.676
R1333 B.n208 B.n88 71.676
R1334 B.n212 B.n89 71.676
R1335 B.n216 B.n90 71.676
R1336 B.n220 B.n91 71.676
R1337 B.n224 B.n92 71.676
R1338 B.n228 B.n93 71.676
R1339 B.n232 B.n94 71.676
R1340 B.n236 B.n95 71.676
R1341 B.n240 B.n96 71.676
R1342 B.n244 B.n97 71.676
R1343 B.n248 B.n98 71.676
R1344 B.n252 B.n99 71.676
R1345 B.n256 B.n100 71.676
R1346 B.n671 B.n101 71.676
R1347 B.n671 B.n670 71.676
R1348 B.n258 B.n100 71.676
R1349 B.n255 B.n99 71.676
R1350 B.n251 B.n98 71.676
R1351 B.n247 B.n97 71.676
R1352 B.n243 B.n96 71.676
R1353 B.n239 B.n95 71.676
R1354 B.n235 B.n94 71.676
R1355 B.n231 B.n93 71.676
R1356 B.n227 B.n92 71.676
R1357 B.n223 B.n91 71.676
R1358 B.n219 B.n90 71.676
R1359 B.n215 B.n89 71.676
R1360 B.n211 B.n88 71.676
R1361 B.n207 B.n87 71.676
R1362 B.n203 B.n86 71.676
R1363 B.n199 B.n85 71.676
R1364 B.n195 B.n84 71.676
R1365 B.n191 B.n83 71.676
R1366 B.n187 B.n82 71.676
R1367 B.n183 B.n81 71.676
R1368 B.n179 B.n80 71.676
R1369 B.n175 B.n79 71.676
R1370 B.n171 B.n78 71.676
R1371 B.n167 B.n77 71.676
R1372 B.n163 B.n76 71.676
R1373 B.n159 B.n75 71.676
R1374 B.n155 B.n74 71.676
R1375 B.n151 B.n73 71.676
R1376 B.n147 B.n72 71.676
R1377 B.n143 B.n71 71.676
R1378 B.n139 B.n70 71.676
R1379 B.n135 B.n69 71.676
R1380 B.n131 B.n68 71.676
R1381 B.n127 B.n67 71.676
R1382 B.n123 B.n66 71.676
R1383 B.n119 B.n65 71.676
R1384 B.n115 B.n64 71.676
R1385 B.n111 B.n63 71.676
R1386 B.n522 B.n521 71.676
R1387 B.n516 B.n327 71.676
R1388 B.n513 B.n328 71.676
R1389 B.n509 B.n329 71.676
R1390 B.n505 B.n330 71.676
R1391 B.n501 B.n331 71.676
R1392 B.n497 B.n332 71.676
R1393 B.n493 B.n333 71.676
R1394 B.n489 B.n334 71.676
R1395 B.n485 B.n335 71.676
R1396 B.n481 B.n336 71.676
R1397 B.n477 B.n337 71.676
R1398 B.n473 B.n338 71.676
R1399 B.n469 B.n339 71.676
R1400 B.n465 B.n340 71.676
R1401 B.n461 B.n341 71.676
R1402 B.n457 B.n342 71.676
R1403 B.n452 B.n343 71.676
R1404 B.n448 B.n344 71.676
R1405 B.n444 B.n345 71.676
R1406 B.n440 B.n346 71.676
R1407 B.n436 B.n347 71.676
R1408 B.n431 B.n348 71.676
R1409 B.n427 B.n349 71.676
R1410 B.n423 B.n350 71.676
R1411 B.n419 B.n351 71.676
R1412 B.n415 B.n352 71.676
R1413 B.n411 B.n353 71.676
R1414 B.n407 B.n354 71.676
R1415 B.n403 B.n355 71.676
R1416 B.n399 B.n356 71.676
R1417 B.n395 B.n357 71.676
R1418 B.n391 B.n358 71.676
R1419 B.n387 B.n359 71.676
R1420 B.n383 B.n360 71.676
R1421 B.n379 B.n361 71.676
R1422 B.n375 B.n362 71.676
R1423 B.n371 B.n363 71.676
R1424 B.n522 B.n365 71.676
R1425 B.n514 B.n327 71.676
R1426 B.n510 B.n328 71.676
R1427 B.n506 B.n329 71.676
R1428 B.n502 B.n330 71.676
R1429 B.n498 B.n331 71.676
R1430 B.n494 B.n332 71.676
R1431 B.n490 B.n333 71.676
R1432 B.n486 B.n334 71.676
R1433 B.n482 B.n335 71.676
R1434 B.n478 B.n336 71.676
R1435 B.n474 B.n337 71.676
R1436 B.n470 B.n338 71.676
R1437 B.n466 B.n339 71.676
R1438 B.n462 B.n340 71.676
R1439 B.n458 B.n341 71.676
R1440 B.n453 B.n342 71.676
R1441 B.n449 B.n343 71.676
R1442 B.n445 B.n344 71.676
R1443 B.n441 B.n345 71.676
R1444 B.n437 B.n346 71.676
R1445 B.n432 B.n347 71.676
R1446 B.n428 B.n348 71.676
R1447 B.n424 B.n349 71.676
R1448 B.n420 B.n350 71.676
R1449 B.n416 B.n351 71.676
R1450 B.n412 B.n352 71.676
R1451 B.n408 B.n353 71.676
R1452 B.n404 B.n354 71.676
R1453 B.n400 B.n355 71.676
R1454 B.n396 B.n356 71.676
R1455 B.n392 B.n357 71.676
R1456 B.n388 B.n358 71.676
R1457 B.n384 B.n359 71.676
R1458 B.n380 B.n360 71.676
R1459 B.n376 B.n361 71.676
R1460 B.n372 B.n362 71.676
R1461 B.n363 B.n326 71.676
R1462 B.n741 B.n740 71.676
R1463 B.n741 B.n2 71.676
R1464 B.n107 B.n106 59.5399
R1465 B.n104 B.n103 59.5399
R1466 B.n434 B.n369 59.5399
R1467 B.n455 B.n367 59.5399
R1468 B.n529 B.n323 50.833
R1469 B.n529 B.n319 50.833
R1470 B.n535 B.n319 50.833
R1471 B.n535 B.n315 50.833
R1472 B.n541 B.n315 50.833
R1473 B.n547 B.n311 50.833
R1474 B.n547 B.n307 50.833
R1475 B.n553 B.n307 50.833
R1476 B.n553 B.n302 50.833
R1477 B.n559 B.n302 50.833
R1478 B.n559 B.n303 50.833
R1479 B.n565 B.n294 50.833
R1480 B.n571 B.n294 50.833
R1481 B.n571 B.n295 50.833
R1482 B.n577 B.n287 50.833
R1483 B.n583 B.n287 50.833
R1484 B.n583 B.n283 50.833
R1485 B.n589 B.n283 50.833
R1486 B.n595 B.n279 50.833
R1487 B.n595 B.n275 50.833
R1488 B.n601 B.n275 50.833
R1489 B.n607 B.n271 50.833
R1490 B.n607 B.n267 50.833
R1491 B.n614 B.n267 50.833
R1492 B.n620 B.n263 50.833
R1493 B.n620 B.n4 50.833
R1494 B.n739 B.n4 50.833
R1495 B.n739 B.n738 50.833
R1496 B.n738 B.n737 50.833
R1497 B.n737 B.n8 50.833
R1498 B.n629 B.n8 50.833
R1499 B.n730 B.n729 50.833
R1500 B.n729 B.n728 50.833
R1501 B.n728 B.n15 50.833
R1502 B.n722 B.n721 50.833
R1503 B.n721 B.n720 50.833
R1504 B.n720 B.n22 50.833
R1505 B.n714 B.n713 50.833
R1506 B.n713 B.n712 50.833
R1507 B.n712 B.n29 50.833
R1508 B.n706 B.n29 50.833
R1509 B.n705 B.n704 50.833
R1510 B.n704 B.n36 50.833
R1511 B.n698 B.n36 50.833
R1512 B.n697 B.n696 50.833
R1513 B.n696 B.n43 50.833
R1514 B.n690 B.n43 50.833
R1515 B.n690 B.n689 50.833
R1516 B.n689 B.n688 50.833
R1517 B.n688 B.n50 50.833
R1518 B.n682 B.n681 50.833
R1519 B.n681 B.n680 50.833
R1520 B.n680 B.n57 50.833
R1521 B.n674 B.n57 50.833
R1522 B.n674 B.n673 50.833
R1523 B.n295 B.t4 49.3379
R1524 B.t5 B.n705 49.3379
R1525 B.t11 B.n311 38.8724
R1526 B.t3 B.n279 38.8724
R1527 B.n614 B.t1 38.8724
R1528 B.n730 B.t6 38.8724
R1529 B.t2 B.n22 38.8724
R1530 B.t15 B.n50 38.8724
R1531 B.n303 B.t0 35.8823
R1532 B.t9 B.n697 35.8823
R1533 B.n520 B.n321 33.2493
R1534 B.n526 B.n525 33.2493
R1535 B.n669 B.n668 33.2493
R1536 B.n109 B.n59 33.2493
R1537 B.n106 B.n105 28.1217
R1538 B.n103 B.n102 28.1217
R1539 B.n369 B.n368 28.1217
R1540 B.n367 B.n366 28.1217
R1541 B.n601 B.t8 25.4167
R1542 B.t8 B.n271 25.4167
R1543 B.t7 B.n15 25.4167
R1544 B.n722 B.t7 25.4167
R1545 B B.n742 18.0485
R1546 B.n565 B.t0 14.9512
R1547 B.n698 B.t9 14.9512
R1548 B.n541 B.t11 11.9611
R1549 B.n589 B.t3 11.9611
R1550 B.t1 B.n263 11.9611
R1551 B.n629 B.t6 11.9611
R1552 B.n714 B.t2 11.9611
R1553 B.n682 B.t15 11.9611
R1554 B.n531 B.n321 10.6151
R1555 B.n532 B.n531 10.6151
R1556 B.n533 B.n532 10.6151
R1557 B.n533 B.n313 10.6151
R1558 B.n543 B.n313 10.6151
R1559 B.n544 B.n543 10.6151
R1560 B.n545 B.n544 10.6151
R1561 B.n545 B.n305 10.6151
R1562 B.n555 B.n305 10.6151
R1563 B.n556 B.n555 10.6151
R1564 B.n557 B.n556 10.6151
R1565 B.n557 B.n297 10.6151
R1566 B.n567 B.n297 10.6151
R1567 B.n568 B.n567 10.6151
R1568 B.n569 B.n568 10.6151
R1569 B.n569 B.n289 10.6151
R1570 B.n579 B.n289 10.6151
R1571 B.n580 B.n579 10.6151
R1572 B.n581 B.n580 10.6151
R1573 B.n581 B.n281 10.6151
R1574 B.n591 B.n281 10.6151
R1575 B.n592 B.n591 10.6151
R1576 B.n593 B.n592 10.6151
R1577 B.n593 B.n273 10.6151
R1578 B.n603 B.n273 10.6151
R1579 B.n604 B.n603 10.6151
R1580 B.n605 B.n604 10.6151
R1581 B.n605 B.n265 10.6151
R1582 B.n616 B.n265 10.6151
R1583 B.n617 B.n616 10.6151
R1584 B.n618 B.n617 10.6151
R1585 B.n618 B.n0 10.6151
R1586 B.n520 B.n519 10.6151
R1587 B.n519 B.n518 10.6151
R1588 B.n518 B.n517 10.6151
R1589 B.n517 B.n515 10.6151
R1590 B.n515 B.n512 10.6151
R1591 B.n512 B.n511 10.6151
R1592 B.n511 B.n508 10.6151
R1593 B.n508 B.n507 10.6151
R1594 B.n507 B.n504 10.6151
R1595 B.n504 B.n503 10.6151
R1596 B.n503 B.n500 10.6151
R1597 B.n500 B.n499 10.6151
R1598 B.n499 B.n496 10.6151
R1599 B.n496 B.n495 10.6151
R1600 B.n495 B.n492 10.6151
R1601 B.n492 B.n491 10.6151
R1602 B.n491 B.n488 10.6151
R1603 B.n488 B.n487 10.6151
R1604 B.n487 B.n484 10.6151
R1605 B.n484 B.n483 10.6151
R1606 B.n483 B.n480 10.6151
R1607 B.n480 B.n479 10.6151
R1608 B.n479 B.n476 10.6151
R1609 B.n476 B.n475 10.6151
R1610 B.n475 B.n472 10.6151
R1611 B.n472 B.n471 10.6151
R1612 B.n471 B.n468 10.6151
R1613 B.n468 B.n467 10.6151
R1614 B.n467 B.n464 10.6151
R1615 B.n464 B.n463 10.6151
R1616 B.n463 B.n460 10.6151
R1617 B.n460 B.n459 10.6151
R1618 B.n459 B.n456 10.6151
R1619 B.n454 B.n451 10.6151
R1620 B.n451 B.n450 10.6151
R1621 B.n450 B.n447 10.6151
R1622 B.n447 B.n446 10.6151
R1623 B.n446 B.n443 10.6151
R1624 B.n443 B.n442 10.6151
R1625 B.n442 B.n439 10.6151
R1626 B.n439 B.n438 10.6151
R1627 B.n438 B.n435 10.6151
R1628 B.n433 B.n430 10.6151
R1629 B.n430 B.n429 10.6151
R1630 B.n429 B.n426 10.6151
R1631 B.n426 B.n425 10.6151
R1632 B.n425 B.n422 10.6151
R1633 B.n422 B.n421 10.6151
R1634 B.n421 B.n418 10.6151
R1635 B.n418 B.n417 10.6151
R1636 B.n417 B.n414 10.6151
R1637 B.n414 B.n413 10.6151
R1638 B.n413 B.n410 10.6151
R1639 B.n410 B.n409 10.6151
R1640 B.n409 B.n406 10.6151
R1641 B.n406 B.n405 10.6151
R1642 B.n405 B.n402 10.6151
R1643 B.n402 B.n401 10.6151
R1644 B.n401 B.n398 10.6151
R1645 B.n398 B.n397 10.6151
R1646 B.n397 B.n394 10.6151
R1647 B.n394 B.n393 10.6151
R1648 B.n393 B.n390 10.6151
R1649 B.n390 B.n389 10.6151
R1650 B.n389 B.n386 10.6151
R1651 B.n386 B.n385 10.6151
R1652 B.n385 B.n382 10.6151
R1653 B.n382 B.n381 10.6151
R1654 B.n381 B.n378 10.6151
R1655 B.n378 B.n377 10.6151
R1656 B.n377 B.n374 10.6151
R1657 B.n374 B.n373 10.6151
R1658 B.n373 B.n370 10.6151
R1659 B.n370 B.n325 10.6151
R1660 B.n525 B.n325 10.6151
R1661 B.n527 B.n526 10.6151
R1662 B.n527 B.n317 10.6151
R1663 B.n537 B.n317 10.6151
R1664 B.n538 B.n537 10.6151
R1665 B.n539 B.n538 10.6151
R1666 B.n539 B.n309 10.6151
R1667 B.n549 B.n309 10.6151
R1668 B.n550 B.n549 10.6151
R1669 B.n551 B.n550 10.6151
R1670 B.n551 B.n300 10.6151
R1671 B.n561 B.n300 10.6151
R1672 B.n562 B.n561 10.6151
R1673 B.n563 B.n562 10.6151
R1674 B.n563 B.n292 10.6151
R1675 B.n573 B.n292 10.6151
R1676 B.n574 B.n573 10.6151
R1677 B.n575 B.n574 10.6151
R1678 B.n575 B.n285 10.6151
R1679 B.n585 B.n285 10.6151
R1680 B.n586 B.n585 10.6151
R1681 B.n587 B.n586 10.6151
R1682 B.n587 B.n277 10.6151
R1683 B.n597 B.n277 10.6151
R1684 B.n598 B.n597 10.6151
R1685 B.n599 B.n598 10.6151
R1686 B.n599 B.n269 10.6151
R1687 B.n609 B.n269 10.6151
R1688 B.n610 B.n609 10.6151
R1689 B.n612 B.n610 10.6151
R1690 B.n612 B.n611 10.6151
R1691 B.n611 B.n261 10.6151
R1692 B.n623 B.n261 10.6151
R1693 B.n624 B.n623 10.6151
R1694 B.n625 B.n624 10.6151
R1695 B.n626 B.n625 10.6151
R1696 B.n627 B.n626 10.6151
R1697 B.n631 B.n627 10.6151
R1698 B.n632 B.n631 10.6151
R1699 B.n633 B.n632 10.6151
R1700 B.n634 B.n633 10.6151
R1701 B.n636 B.n634 10.6151
R1702 B.n637 B.n636 10.6151
R1703 B.n638 B.n637 10.6151
R1704 B.n639 B.n638 10.6151
R1705 B.n641 B.n639 10.6151
R1706 B.n642 B.n641 10.6151
R1707 B.n643 B.n642 10.6151
R1708 B.n644 B.n643 10.6151
R1709 B.n646 B.n644 10.6151
R1710 B.n647 B.n646 10.6151
R1711 B.n648 B.n647 10.6151
R1712 B.n649 B.n648 10.6151
R1713 B.n651 B.n649 10.6151
R1714 B.n652 B.n651 10.6151
R1715 B.n653 B.n652 10.6151
R1716 B.n654 B.n653 10.6151
R1717 B.n656 B.n654 10.6151
R1718 B.n657 B.n656 10.6151
R1719 B.n658 B.n657 10.6151
R1720 B.n659 B.n658 10.6151
R1721 B.n661 B.n659 10.6151
R1722 B.n662 B.n661 10.6151
R1723 B.n663 B.n662 10.6151
R1724 B.n664 B.n663 10.6151
R1725 B.n666 B.n664 10.6151
R1726 B.n667 B.n666 10.6151
R1727 B.n668 B.n667 10.6151
R1728 B.n734 B.n1 10.6151
R1729 B.n734 B.n733 10.6151
R1730 B.n733 B.n732 10.6151
R1731 B.n732 B.n10 10.6151
R1732 B.n726 B.n10 10.6151
R1733 B.n726 B.n725 10.6151
R1734 B.n725 B.n724 10.6151
R1735 B.n724 B.n17 10.6151
R1736 B.n718 B.n17 10.6151
R1737 B.n718 B.n717 10.6151
R1738 B.n717 B.n716 10.6151
R1739 B.n716 B.n24 10.6151
R1740 B.n710 B.n24 10.6151
R1741 B.n710 B.n709 10.6151
R1742 B.n709 B.n708 10.6151
R1743 B.n708 B.n31 10.6151
R1744 B.n702 B.n31 10.6151
R1745 B.n702 B.n701 10.6151
R1746 B.n701 B.n700 10.6151
R1747 B.n700 B.n38 10.6151
R1748 B.n694 B.n38 10.6151
R1749 B.n694 B.n693 10.6151
R1750 B.n693 B.n692 10.6151
R1751 B.n692 B.n45 10.6151
R1752 B.n686 B.n45 10.6151
R1753 B.n686 B.n685 10.6151
R1754 B.n685 B.n684 10.6151
R1755 B.n684 B.n52 10.6151
R1756 B.n678 B.n52 10.6151
R1757 B.n678 B.n677 10.6151
R1758 B.n677 B.n676 10.6151
R1759 B.n676 B.n59 10.6151
R1760 B.n110 B.n109 10.6151
R1761 B.n113 B.n110 10.6151
R1762 B.n114 B.n113 10.6151
R1763 B.n117 B.n114 10.6151
R1764 B.n118 B.n117 10.6151
R1765 B.n121 B.n118 10.6151
R1766 B.n122 B.n121 10.6151
R1767 B.n125 B.n122 10.6151
R1768 B.n126 B.n125 10.6151
R1769 B.n129 B.n126 10.6151
R1770 B.n130 B.n129 10.6151
R1771 B.n133 B.n130 10.6151
R1772 B.n134 B.n133 10.6151
R1773 B.n137 B.n134 10.6151
R1774 B.n138 B.n137 10.6151
R1775 B.n141 B.n138 10.6151
R1776 B.n142 B.n141 10.6151
R1777 B.n145 B.n142 10.6151
R1778 B.n146 B.n145 10.6151
R1779 B.n149 B.n146 10.6151
R1780 B.n150 B.n149 10.6151
R1781 B.n153 B.n150 10.6151
R1782 B.n154 B.n153 10.6151
R1783 B.n157 B.n154 10.6151
R1784 B.n158 B.n157 10.6151
R1785 B.n161 B.n158 10.6151
R1786 B.n162 B.n161 10.6151
R1787 B.n165 B.n162 10.6151
R1788 B.n166 B.n165 10.6151
R1789 B.n169 B.n166 10.6151
R1790 B.n170 B.n169 10.6151
R1791 B.n173 B.n170 10.6151
R1792 B.n174 B.n173 10.6151
R1793 B.n178 B.n177 10.6151
R1794 B.n181 B.n178 10.6151
R1795 B.n182 B.n181 10.6151
R1796 B.n185 B.n182 10.6151
R1797 B.n186 B.n185 10.6151
R1798 B.n189 B.n186 10.6151
R1799 B.n190 B.n189 10.6151
R1800 B.n193 B.n190 10.6151
R1801 B.n194 B.n193 10.6151
R1802 B.n198 B.n197 10.6151
R1803 B.n201 B.n198 10.6151
R1804 B.n202 B.n201 10.6151
R1805 B.n205 B.n202 10.6151
R1806 B.n206 B.n205 10.6151
R1807 B.n209 B.n206 10.6151
R1808 B.n210 B.n209 10.6151
R1809 B.n213 B.n210 10.6151
R1810 B.n214 B.n213 10.6151
R1811 B.n217 B.n214 10.6151
R1812 B.n218 B.n217 10.6151
R1813 B.n221 B.n218 10.6151
R1814 B.n222 B.n221 10.6151
R1815 B.n225 B.n222 10.6151
R1816 B.n226 B.n225 10.6151
R1817 B.n229 B.n226 10.6151
R1818 B.n230 B.n229 10.6151
R1819 B.n233 B.n230 10.6151
R1820 B.n234 B.n233 10.6151
R1821 B.n237 B.n234 10.6151
R1822 B.n238 B.n237 10.6151
R1823 B.n241 B.n238 10.6151
R1824 B.n242 B.n241 10.6151
R1825 B.n245 B.n242 10.6151
R1826 B.n246 B.n245 10.6151
R1827 B.n249 B.n246 10.6151
R1828 B.n250 B.n249 10.6151
R1829 B.n253 B.n250 10.6151
R1830 B.n254 B.n253 10.6151
R1831 B.n257 B.n254 10.6151
R1832 B.n259 B.n257 10.6151
R1833 B.n260 B.n259 10.6151
R1834 B.n669 B.n260 10.6151
R1835 B.n456 B.n455 9.36635
R1836 B.n434 B.n433 9.36635
R1837 B.n174 B.n107 9.36635
R1838 B.n197 B.n104 9.36635
R1839 B.n742 B.n0 8.11757
R1840 B.n742 B.n1 8.11757
R1841 B.n577 B.t4 1.49557
R1842 B.n706 B.t5 1.49557
R1843 B.n455 B.n454 1.24928
R1844 B.n435 B.n434 1.24928
R1845 B.n177 B.n107 1.24928
R1846 B.n194 B.n104 1.24928
R1847 VN.n4 VN.t6 260.755
R1848 VN.n23 VN.t7 260.755
R1849 VN.n17 VN.t1 238.203
R1850 VN.n36 VN.t0 238.203
R1851 VN.n10 VN.t4 203.13
R1852 VN.n5 VN.t5 203.13
R1853 VN.n1 VN.t3 203.13
R1854 VN.n29 VN.t2 203.13
R1855 VN.n24 VN.t9 203.13
R1856 VN.n20 VN.t8 203.13
R1857 VN.n35 VN.n19 161.3
R1858 VN.n34 VN.n33 161.3
R1859 VN.n32 VN.n31 161.3
R1860 VN.n30 VN.n21 161.3
R1861 VN.n29 VN.n28 161.3
R1862 VN.n27 VN.n22 161.3
R1863 VN.n26 VN.n25 161.3
R1864 VN.n16 VN.n0 161.3
R1865 VN.n15 VN.n14 161.3
R1866 VN.n13 VN.n12 161.3
R1867 VN.n11 VN.n2 161.3
R1868 VN.n10 VN.n9 161.3
R1869 VN.n8 VN.n3 161.3
R1870 VN.n7 VN.n6 161.3
R1871 VN.n37 VN.n36 80.6037
R1872 VN.n18 VN.n17 80.6037
R1873 VN.n6 VN.n3 56.5617
R1874 VN.n12 VN.n11 56.5617
R1875 VN.n25 VN.n22 56.5617
R1876 VN.n31 VN.n30 56.5617
R1877 VN.n17 VN.n16 48.6923
R1878 VN.n36 VN.n35 48.6923
R1879 VN VN.n37 43.5862
R1880 VN.n5 VN.n4 34.7238
R1881 VN.n24 VN.n23 34.7238
R1882 VN.n26 VN.n23 28.3586
R1883 VN.n7 VN.n4 28.3586
R1884 VN.n10 VN.n3 24.5923
R1885 VN.n11 VN.n10 24.5923
R1886 VN.n16 VN.n15 24.5923
R1887 VN.n30 VN.n29 24.5923
R1888 VN.n29 VN.n22 24.5923
R1889 VN.n35 VN.n34 24.5923
R1890 VN.n6 VN.n5 22.1332
R1891 VN.n12 VN.n1 22.1332
R1892 VN.n25 VN.n24 22.1332
R1893 VN.n31 VN.n20 22.1332
R1894 VN.n15 VN.n1 2.45968
R1895 VN.n34 VN.n20 2.45968
R1896 VN.n37 VN.n19 0.285035
R1897 VN.n18 VN.n0 0.285035
R1898 VN.n33 VN.n19 0.189894
R1899 VN.n33 VN.n32 0.189894
R1900 VN.n32 VN.n21 0.189894
R1901 VN.n28 VN.n21 0.189894
R1902 VN.n28 VN.n27 0.189894
R1903 VN.n27 VN.n26 0.189894
R1904 VN.n8 VN.n7 0.189894
R1905 VN.n9 VN.n8 0.189894
R1906 VN.n9 VN.n2 0.189894
R1907 VN.n13 VN.n2 0.189894
R1908 VN.n14 VN.n13 0.189894
R1909 VN.n14 VN.n0 0.189894
R1910 VN VN.n18 0.146778
R1911 VDD2.n97 VDD2.n53 289.615
R1912 VDD2.n44 VDD2.n0 289.615
R1913 VDD2.n98 VDD2.n97 185
R1914 VDD2.n96 VDD2.n95 185
R1915 VDD2.n57 VDD2.n56 185
R1916 VDD2.n61 VDD2.n59 185
R1917 VDD2.n90 VDD2.n89 185
R1918 VDD2.n88 VDD2.n87 185
R1919 VDD2.n63 VDD2.n62 185
R1920 VDD2.n82 VDD2.n81 185
R1921 VDD2.n80 VDD2.n79 185
R1922 VDD2.n67 VDD2.n66 185
R1923 VDD2.n74 VDD2.n73 185
R1924 VDD2.n72 VDD2.n71 185
R1925 VDD2.n17 VDD2.n16 185
R1926 VDD2.n19 VDD2.n18 185
R1927 VDD2.n12 VDD2.n11 185
R1928 VDD2.n25 VDD2.n24 185
R1929 VDD2.n27 VDD2.n26 185
R1930 VDD2.n8 VDD2.n7 185
R1931 VDD2.n34 VDD2.n33 185
R1932 VDD2.n35 VDD2.n6 185
R1933 VDD2.n37 VDD2.n36 185
R1934 VDD2.n4 VDD2.n3 185
R1935 VDD2.n43 VDD2.n42 185
R1936 VDD2.n45 VDD2.n44 185
R1937 VDD2.n70 VDD2.t9 149.524
R1938 VDD2.n15 VDD2.t3 149.524
R1939 VDD2.n97 VDD2.n96 104.615
R1940 VDD2.n96 VDD2.n56 104.615
R1941 VDD2.n61 VDD2.n56 104.615
R1942 VDD2.n89 VDD2.n61 104.615
R1943 VDD2.n89 VDD2.n88 104.615
R1944 VDD2.n88 VDD2.n62 104.615
R1945 VDD2.n81 VDD2.n62 104.615
R1946 VDD2.n81 VDD2.n80 104.615
R1947 VDD2.n80 VDD2.n66 104.615
R1948 VDD2.n73 VDD2.n66 104.615
R1949 VDD2.n73 VDD2.n72 104.615
R1950 VDD2.n18 VDD2.n17 104.615
R1951 VDD2.n18 VDD2.n11 104.615
R1952 VDD2.n25 VDD2.n11 104.615
R1953 VDD2.n26 VDD2.n25 104.615
R1954 VDD2.n26 VDD2.n7 104.615
R1955 VDD2.n34 VDD2.n7 104.615
R1956 VDD2.n35 VDD2.n34 104.615
R1957 VDD2.n36 VDD2.n35 104.615
R1958 VDD2.n36 VDD2.n3 104.615
R1959 VDD2.n43 VDD2.n3 104.615
R1960 VDD2.n44 VDD2.n43 104.615
R1961 VDD2.n52 VDD2.n51 67.7628
R1962 VDD2 VDD2.n105 67.76
R1963 VDD2.n104 VDD2.n103 66.8808
R1964 VDD2.n50 VDD2.n49 66.8807
R1965 VDD2.n50 VDD2.n48 53.9929
R1966 VDD2.n102 VDD2.n101 52.7429
R1967 VDD2.n72 VDD2.t9 52.3082
R1968 VDD2.n17 VDD2.t3 52.3082
R1969 VDD2.n102 VDD2.n52 37.7907
R1970 VDD2.n59 VDD2.n57 13.1884
R1971 VDD2.n37 VDD2.n4 13.1884
R1972 VDD2.n95 VDD2.n94 12.8005
R1973 VDD2.n91 VDD2.n90 12.8005
R1974 VDD2.n38 VDD2.n6 12.8005
R1975 VDD2.n42 VDD2.n41 12.8005
R1976 VDD2.n98 VDD2.n55 12.0247
R1977 VDD2.n87 VDD2.n60 12.0247
R1978 VDD2.n33 VDD2.n32 12.0247
R1979 VDD2.n45 VDD2.n2 12.0247
R1980 VDD2.n99 VDD2.n53 11.249
R1981 VDD2.n86 VDD2.n63 11.249
R1982 VDD2.n31 VDD2.n8 11.249
R1983 VDD2.n46 VDD2.n0 11.249
R1984 VDD2.n83 VDD2.n82 10.4732
R1985 VDD2.n28 VDD2.n27 10.4732
R1986 VDD2.n71 VDD2.n70 10.2747
R1987 VDD2.n16 VDD2.n15 10.2747
R1988 VDD2.n79 VDD2.n65 9.69747
R1989 VDD2.n24 VDD2.n10 9.69747
R1990 VDD2.n101 VDD2.n100 9.45567
R1991 VDD2.n48 VDD2.n47 9.45567
R1992 VDD2.n69 VDD2.n68 9.3005
R1993 VDD2.n76 VDD2.n75 9.3005
R1994 VDD2.n78 VDD2.n77 9.3005
R1995 VDD2.n65 VDD2.n64 9.3005
R1996 VDD2.n84 VDD2.n83 9.3005
R1997 VDD2.n86 VDD2.n85 9.3005
R1998 VDD2.n60 VDD2.n58 9.3005
R1999 VDD2.n92 VDD2.n91 9.3005
R2000 VDD2.n100 VDD2.n99 9.3005
R2001 VDD2.n55 VDD2.n54 9.3005
R2002 VDD2.n94 VDD2.n93 9.3005
R2003 VDD2.n47 VDD2.n46 9.3005
R2004 VDD2.n2 VDD2.n1 9.3005
R2005 VDD2.n41 VDD2.n40 9.3005
R2006 VDD2.n14 VDD2.n13 9.3005
R2007 VDD2.n21 VDD2.n20 9.3005
R2008 VDD2.n23 VDD2.n22 9.3005
R2009 VDD2.n10 VDD2.n9 9.3005
R2010 VDD2.n29 VDD2.n28 9.3005
R2011 VDD2.n31 VDD2.n30 9.3005
R2012 VDD2.n32 VDD2.n5 9.3005
R2013 VDD2.n39 VDD2.n38 9.3005
R2014 VDD2.n78 VDD2.n67 8.92171
R2015 VDD2.n23 VDD2.n12 8.92171
R2016 VDD2.n75 VDD2.n74 8.14595
R2017 VDD2.n20 VDD2.n19 8.14595
R2018 VDD2.n71 VDD2.n69 7.3702
R2019 VDD2.n16 VDD2.n14 7.3702
R2020 VDD2.n74 VDD2.n69 5.81868
R2021 VDD2.n19 VDD2.n14 5.81868
R2022 VDD2.n75 VDD2.n67 5.04292
R2023 VDD2.n20 VDD2.n12 5.04292
R2024 VDD2.n79 VDD2.n78 4.26717
R2025 VDD2.n24 VDD2.n23 4.26717
R2026 VDD2.n82 VDD2.n65 3.49141
R2027 VDD2.n27 VDD2.n10 3.49141
R2028 VDD2.n70 VDD2.n68 2.84303
R2029 VDD2.n15 VDD2.n13 2.84303
R2030 VDD2.n101 VDD2.n53 2.71565
R2031 VDD2.n83 VDD2.n63 2.71565
R2032 VDD2.n28 VDD2.n8 2.71565
R2033 VDD2.n48 VDD2.n0 2.71565
R2034 VDD2.n105 VDD2.t0 2.09796
R2035 VDD2.n105 VDD2.t2 2.09796
R2036 VDD2.n103 VDD2.t1 2.09796
R2037 VDD2.n103 VDD2.t7 2.09796
R2038 VDD2.n51 VDD2.t6 2.09796
R2039 VDD2.n51 VDD2.t8 2.09796
R2040 VDD2.n49 VDD2.t4 2.09796
R2041 VDD2.n49 VDD2.t5 2.09796
R2042 VDD2.n99 VDD2.n98 1.93989
R2043 VDD2.n87 VDD2.n86 1.93989
R2044 VDD2.n33 VDD2.n31 1.93989
R2045 VDD2.n46 VDD2.n45 1.93989
R2046 VDD2.n104 VDD2.n102 1.2505
R2047 VDD2.n95 VDD2.n55 1.16414
R2048 VDD2.n90 VDD2.n60 1.16414
R2049 VDD2.n32 VDD2.n6 1.16414
R2050 VDD2.n42 VDD2.n2 1.16414
R2051 VDD2.n94 VDD2.n57 0.388379
R2052 VDD2.n91 VDD2.n59 0.388379
R2053 VDD2.n38 VDD2.n37 0.388379
R2054 VDD2.n41 VDD2.n4 0.388379
R2055 VDD2 VDD2.n104 0.37119
R2056 VDD2.n52 VDD2.n50 0.257654
R2057 VDD2.n100 VDD2.n54 0.155672
R2058 VDD2.n93 VDD2.n54 0.155672
R2059 VDD2.n93 VDD2.n92 0.155672
R2060 VDD2.n92 VDD2.n58 0.155672
R2061 VDD2.n85 VDD2.n58 0.155672
R2062 VDD2.n85 VDD2.n84 0.155672
R2063 VDD2.n84 VDD2.n64 0.155672
R2064 VDD2.n77 VDD2.n64 0.155672
R2065 VDD2.n77 VDD2.n76 0.155672
R2066 VDD2.n76 VDD2.n68 0.155672
R2067 VDD2.n21 VDD2.n13 0.155672
R2068 VDD2.n22 VDD2.n21 0.155672
R2069 VDD2.n22 VDD2.n9 0.155672
R2070 VDD2.n29 VDD2.n9 0.155672
R2071 VDD2.n30 VDD2.n29 0.155672
R2072 VDD2.n30 VDD2.n5 0.155672
R2073 VDD2.n39 VDD2.n5 0.155672
R2074 VDD2.n40 VDD2.n39 0.155672
R2075 VDD2.n40 VDD2.n1 0.155672
R2076 VDD2.n47 VDD2.n1 0.155672
C0 VP VDD1 6.88566f
C1 VN VDD1 0.150443f
C2 VP VTAIL 6.78287f
C3 VTAIL VN 6.76846f
C4 VDD2 VDD1 1.23152f
C5 VDD2 VTAIL 10.000799f
C6 VP VN 5.73759f
C7 VTAIL VDD1 9.96129f
C8 VDD2 VP 0.395127f
C9 VDD2 VN 6.64454f
C10 VDD2 B 5.008248f
C11 VDD1 B 4.967028f
C12 VTAIL B 5.992056f
C13 VN B 11.02986f
C14 VP B 9.358879f
C15 VDD2.n0 B 0.032965f
C16 VDD2.n1 B 0.023011f
C17 VDD2.n2 B 0.012365f
C18 VDD2.n3 B 0.029227f
C19 VDD2.n4 B 0.012729f
C20 VDD2.n5 B 0.023011f
C21 VDD2.n6 B 0.013093f
C22 VDD2.n7 B 0.029227f
C23 VDD2.n8 B 0.013093f
C24 VDD2.n9 B 0.023011f
C25 VDD2.n10 B 0.012365f
C26 VDD2.n11 B 0.029227f
C27 VDD2.n12 B 0.013093f
C28 VDD2.n13 B 0.898847f
C29 VDD2.n14 B 0.012365f
C30 VDD2.t3 B 0.04905f
C31 VDD2.n15 B 0.143301f
C32 VDD2.n16 B 0.020661f
C33 VDD2.n17 B 0.02192f
C34 VDD2.n18 B 0.029227f
C35 VDD2.n19 B 0.013093f
C36 VDD2.n20 B 0.012365f
C37 VDD2.n21 B 0.023011f
C38 VDD2.n22 B 0.023011f
C39 VDD2.n23 B 0.012365f
C40 VDD2.n24 B 0.013093f
C41 VDD2.n25 B 0.029227f
C42 VDD2.n26 B 0.029227f
C43 VDD2.n27 B 0.013093f
C44 VDD2.n28 B 0.012365f
C45 VDD2.n29 B 0.023011f
C46 VDD2.n30 B 0.023011f
C47 VDD2.n31 B 0.012365f
C48 VDD2.n32 B 0.012365f
C49 VDD2.n33 B 0.013093f
C50 VDD2.n34 B 0.029227f
C51 VDD2.n35 B 0.029227f
C52 VDD2.n36 B 0.029227f
C53 VDD2.n37 B 0.012729f
C54 VDD2.n38 B 0.012365f
C55 VDD2.n39 B 0.023011f
C56 VDD2.n40 B 0.023011f
C57 VDD2.n41 B 0.012365f
C58 VDD2.n42 B 0.013093f
C59 VDD2.n43 B 0.029227f
C60 VDD2.n44 B 0.06437f
C61 VDD2.n45 B 0.013093f
C62 VDD2.n46 B 0.012365f
C63 VDD2.n47 B 0.059477f
C64 VDD2.n48 B 0.055414f
C65 VDD2.t4 B 0.171659f
C66 VDD2.t5 B 0.171659f
C67 VDD2.n49 B 1.50781f
C68 VDD2.n50 B 0.435268f
C69 VDD2.t6 B 0.171659f
C70 VDD2.t8 B 0.171659f
C71 VDD2.n51 B 1.5124f
C72 VDD2.n52 B 1.81001f
C73 VDD2.n53 B 0.032965f
C74 VDD2.n54 B 0.023011f
C75 VDD2.n55 B 0.012365f
C76 VDD2.n56 B 0.029227f
C77 VDD2.n57 B 0.012729f
C78 VDD2.n58 B 0.023011f
C79 VDD2.n59 B 0.012729f
C80 VDD2.n60 B 0.012365f
C81 VDD2.n61 B 0.029227f
C82 VDD2.n62 B 0.029227f
C83 VDD2.n63 B 0.013093f
C84 VDD2.n64 B 0.023011f
C85 VDD2.n65 B 0.012365f
C86 VDD2.n66 B 0.029227f
C87 VDD2.n67 B 0.013093f
C88 VDD2.n68 B 0.898847f
C89 VDD2.n69 B 0.012365f
C90 VDD2.t9 B 0.04905f
C91 VDD2.n70 B 0.143301f
C92 VDD2.n71 B 0.020661f
C93 VDD2.n72 B 0.02192f
C94 VDD2.n73 B 0.029227f
C95 VDD2.n74 B 0.013093f
C96 VDD2.n75 B 0.012365f
C97 VDD2.n76 B 0.023011f
C98 VDD2.n77 B 0.023011f
C99 VDD2.n78 B 0.012365f
C100 VDD2.n79 B 0.013093f
C101 VDD2.n80 B 0.029227f
C102 VDD2.n81 B 0.029227f
C103 VDD2.n82 B 0.013093f
C104 VDD2.n83 B 0.012365f
C105 VDD2.n84 B 0.023011f
C106 VDD2.n85 B 0.023011f
C107 VDD2.n86 B 0.012365f
C108 VDD2.n87 B 0.013093f
C109 VDD2.n88 B 0.029227f
C110 VDD2.n89 B 0.029227f
C111 VDD2.n90 B 0.013093f
C112 VDD2.n91 B 0.012365f
C113 VDD2.n92 B 0.023011f
C114 VDD2.n93 B 0.023011f
C115 VDD2.n94 B 0.012365f
C116 VDD2.n95 B 0.013093f
C117 VDD2.n96 B 0.029227f
C118 VDD2.n97 B 0.06437f
C119 VDD2.n98 B 0.013093f
C120 VDD2.n99 B 0.012365f
C121 VDD2.n100 B 0.059477f
C122 VDD2.n101 B 0.052159f
C123 VDD2.n102 B 1.9513f
C124 VDD2.t1 B 0.171659f
C125 VDD2.t7 B 0.171659f
C126 VDD2.n103 B 1.50782f
C127 VDD2.n104 B 0.304265f
C128 VDD2.t0 B 0.171659f
C129 VDD2.t2 B 0.171659f
C130 VDD2.n105 B 1.51237f
C131 VN.n0 B 0.046986f
C132 VN.t3 B 1.00649f
C133 VN.n1 B 0.380011f
C134 VN.n2 B 0.035212f
C135 VN.t4 B 1.00649f
C136 VN.n3 B 0.04875f
C137 VN.t6 B 1.1054f
C138 VN.n4 B 0.427747f
C139 VN.t5 B 1.00649f
C140 VN.n5 B 0.433877f
C141 VN.n6 B 0.050398f
C142 VN.n7 B 0.183461f
C143 VN.n8 B 0.035212f
C144 VN.n9 B 0.035212f
C145 VN.n10 B 0.413073f
C146 VN.n11 B 0.04875f
C147 VN.n12 B 0.050398f
C148 VN.n13 B 0.035212f
C149 VN.n14 B 0.035212f
C150 VN.n15 B 0.036285f
C151 VN.n16 B 0.041436f
C152 VN.t1 B 1.06654f
C153 VN.n17 B 0.441036f
C154 VN.n18 B 0.032977f
C155 VN.n19 B 0.046986f
C156 VN.t8 B 1.00649f
C157 VN.n20 B 0.380011f
C158 VN.n21 B 0.035212f
C159 VN.t2 B 1.00649f
C160 VN.n22 B 0.04875f
C161 VN.t7 B 1.1054f
C162 VN.n23 B 0.427747f
C163 VN.t9 B 1.00649f
C164 VN.n24 B 0.433877f
C165 VN.n25 B 0.050398f
C166 VN.n26 B 0.183461f
C167 VN.n27 B 0.035212f
C168 VN.n28 B 0.035212f
C169 VN.n29 B 0.413073f
C170 VN.n30 B 0.04875f
C171 VN.n31 B 0.050398f
C172 VN.n32 B 0.035212f
C173 VN.n33 B 0.035212f
C174 VN.n34 B 0.036285f
C175 VN.n35 B 0.041436f
C176 VN.t0 B 1.06654f
C177 VN.n36 B 0.441036f
C178 VN.n37 B 1.56058f
C179 VTAIL.t6 B 0.188645f
C180 VTAIL.t7 B 0.188645f
C181 VTAIL.n0 B 1.5914f
C182 VTAIL.n1 B 0.40391f
C183 VTAIL.n2 B 0.036227f
C184 VTAIL.n3 B 0.025288f
C185 VTAIL.n4 B 0.013589f
C186 VTAIL.n5 B 0.032119f
C187 VTAIL.n6 B 0.013988f
C188 VTAIL.n7 B 0.025288f
C189 VTAIL.n8 B 0.014388f
C190 VTAIL.n9 B 0.032119f
C191 VTAIL.n10 B 0.014388f
C192 VTAIL.n11 B 0.025288f
C193 VTAIL.n12 B 0.013589f
C194 VTAIL.n13 B 0.032119f
C195 VTAIL.n14 B 0.014388f
C196 VTAIL.n15 B 0.987791f
C197 VTAIL.n16 B 0.013589f
C198 VTAIL.t18 B 0.053904f
C199 VTAIL.n17 B 0.157481f
C200 VTAIL.n18 B 0.022706f
C201 VTAIL.n19 B 0.024089f
C202 VTAIL.n20 B 0.032119f
C203 VTAIL.n21 B 0.014388f
C204 VTAIL.n22 B 0.013589f
C205 VTAIL.n23 B 0.025288f
C206 VTAIL.n24 B 0.025288f
C207 VTAIL.n25 B 0.013589f
C208 VTAIL.n26 B 0.014388f
C209 VTAIL.n27 B 0.032119f
C210 VTAIL.n28 B 0.032119f
C211 VTAIL.n29 B 0.014388f
C212 VTAIL.n30 B 0.013589f
C213 VTAIL.n31 B 0.025288f
C214 VTAIL.n32 B 0.025288f
C215 VTAIL.n33 B 0.013589f
C216 VTAIL.n34 B 0.013589f
C217 VTAIL.n35 B 0.014388f
C218 VTAIL.n36 B 0.032119f
C219 VTAIL.n37 B 0.032119f
C220 VTAIL.n38 B 0.032119f
C221 VTAIL.n39 B 0.013988f
C222 VTAIL.n40 B 0.013589f
C223 VTAIL.n41 B 0.025288f
C224 VTAIL.n42 B 0.025288f
C225 VTAIL.n43 B 0.013589f
C226 VTAIL.n44 B 0.014388f
C227 VTAIL.n45 B 0.032119f
C228 VTAIL.n46 B 0.070739f
C229 VTAIL.n47 B 0.014388f
C230 VTAIL.n48 B 0.013589f
C231 VTAIL.n49 B 0.065362f
C232 VTAIL.n50 B 0.039907f
C233 VTAIL.n51 B 0.216575f
C234 VTAIL.t10 B 0.188645f
C235 VTAIL.t19 B 0.188645f
C236 VTAIL.n52 B 1.5914f
C237 VTAIL.n53 B 0.437276f
C238 VTAIL.t13 B 0.188645f
C239 VTAIL.t12 B 0.188645f
C240 VTAIL.n54 B 1.5914f
C241 VTAIL.n55 B 1.54576f
C242 VTAIL.t0 B 0.188645f
C243 VTAIL.t4 B 0.188645f
C244 VTAIL.n56 B 1.59141f
C245 VTAIL.n57 B 1.54575f
C246 VTAIL.t3 B 0.188645f
C247 VTAIL.t8 B 0.188645f
C248 VTAIL.n58 B 1.59141f
C249 VTAIL.n59 B 0.437267f
C250 VTAIL.n60 B 0.036227f
C251 VTAIL.n61 B 0.025288f
C252 VTAIL.n62 B 0.013589f
C253 VTAIL.n63 B 0.032119f
C254 VTAIL.n64 B 0.013988f
C255 VTAIL.n65 B 0.025288f
C256 VTAIL.n66 B 0.013988f
C257 VTAIL.n67 B 0.013589f
C258 VTAIL.n68 B 0.032119f
C259 VTAIL.n69 B 0.032119f
C260 VTAIL.n70 B 0.014388f
C261 VTAIL.n71 B 0.025288f
C262 VTAIL.n72 B 0.013589f
C263 VTAIL.n73 B 0.032119f
C264 VTAIL.n74 B 0.014388f
C265 VTAIL.n75 B 0.987791f
C266 VTAIL.n76 B 0.013589f
C267 VTAIL.t1 B 0.053904f
C268 VTAIL.n77 B 0.157481f
C269 VTAIL.n78 B 0.022706f
C270 VTAIL.n79 B 0.024089f
C271 VTAIL.n80 B 0.032119f
C272 VTAIL.n81 B 0.014388f
C273 VTAIL.n82 B 0.013589f
C274 VTAIL.n83 B 0.025288f
C275 VTAIL.n84 B 0.025288f
C276 VTAIL.n85 B 0.013589f
C277 VTAIL.n86 B 0.014388f
C278 VTAIL.n87 B 0.032119f
C279 VTAIL.n88 B 0.032119f
C280 VTAIL.n89 B 0.014388f
C281 VTAIL.n90 B 0.013589f
C282 VTAIL.n91 B 0.025288f
C283 VTAIL.n92 B 0.025288f
C284 VTAIL.n93 B 0.013589f
C285 VTAIL.n94 B 0.014388f
C286 VTAIL.n95 B 0.032119f
C287 VTAIL.n96 B 0.032119f
C288 VTAIL.n97 B 0.014388f
C289 VTAIL.n98 B 0.013589f
C290 VTAIL.n99 B 0.025288f
C291 VTAIL.n100 B 0.025288f
C292 VTAIL.n101 B 0.013589f
C293 VTAIL.n102 B 0.014388f
C294 VTAIL.n103 B 0.032119f
C295 VTAIL.n104 B 0.070739f
C296 VTAIL.n105 B 0.014388f
C297 VTAIL.n106 B 0.013589f
C298 VTAIL.n107 B 0.065362f
C299 VTAIL.n108 B 0.039907f
C300 VTAIL.n109 B 0.216575f
C301 VTAIL.t16 B 0.188645f
C302 VTAIL.t14 B 0.188645f
C303 VTAIL.n110 B 1.59141f
C304 VTAIL.n111 B 0.424623f
C305 VTAIL.t11 B 0.188645f
C306 VTAIL.t17 B 0.188645f
C307 VTAIL.n112 B 1.59141f
C308 VTAIL.n113 B 0.437267f
C309 VTAIL.n114 B 0.036227f
C310 VTAIL.n115 B 0.025288f
C311 VTAIL.n116 B 0.013589f
C312 VTAIL.n117 B 0.032119f
C313 VTAIL.n118 B 0.013988f
C314 VTAIL.n119 B 0.025288f
C315 VTAIL.n120 B 0.013988f
C316 VTAIL.n121 B 0.013589f
C317 VTAIL.n122 B 0.032119f
C318 VTAIL.n123 B 0.032119f
C319 VTAIL.n124 B 0.014388f
C320 VTAIL.n125 B 0.025288f
C321 VTAIL.n126 B 0.013589f
C322 VTAIL.n127 B 0.032119f
C323 VTAIL.n128 B 0.014388f
C324 VTAIL.n129 B 0.987791f
C325 VTAIL.n130 B 0.013589f
C326 VTAIL.t15 B 0.053904f
C327 VTAIL.n131 B 0.157481f
C328 VTAIL.n132 B 0.022706f
C329 VTAIL.n133 B 0.024089f
C330 VTAIL.n134 B 0.032119f
C331 VTAIL.n135 B 0.014388f
C332 VTAIL.n136 B 0.013589f
C333 VTAIL.n137 B 0.025288f
C334 VTAIL.n138 B 0.025288f
C335 VTAIL.n139 B 0.013589f
C336 VTAIL.n140 B 0.014388f
C337 VTAIL.n141 B 0.032119f
C338 VTAIL.n142 B 0.032119f
C339 VTAIL.n143 B 0.014388f
C340 VTAIL.n144 B 0.013589f
C341 VTAIL.n145 B 0.025288f
C342 VTAIL.n146 B 0.025288f
C343 VTAIL.n147 B 0.013589f
C344 VTAIL.n148 B 0.014388f
C345 VTAIL.n149 B 0.032119f
C346 VTAIL.n150 B 0.032119f
C347 VTAIL.n151 B 0.014388f
C348 VTAIL.n152 B 0.013589f
C349 VTAIL.n153 B 0.025288f
C350 VTAIL.n154 B 0.025288f
C351 VTAIL.n155 B 0.013589f
C352 VTAIL.n156 B 0.014388f
C353 VTAIL.n157 B 0.032119f
C354 VTAIL.n158 B 0.070739f
C355 VTAIL.n159 B 0.014388f
C356 VTAIL.n160 B 0.013589f
C357 VTAIL.n161 B 0.065362f
C358 VTAIL.n162 B 0.039907f
C359 VTAIL.n163 B 1.23585f
C360 VTAIL.n164 B 0.036227f
C361 VTAIL.n165 B 0.025288f
C362 VTAIL.n166 B 0.013589f
C363 VTAIL.n167 B 0.032119f
C364 VTAIL.n168 B 0.013988f
C365 VTAIL.n169 B 0.025288f
C366 VTAIL.n170 B 0.014388f
C367 VTAIL.n171 B 0.032119f
C368 VTAIL.n172 B 0.014388f
C369 VTAIL.n173 B 0.025288f
C370 VTAIL.n174 B 0.013589f
C371 VTAIL.n175 B 0.032119f
C372 VTAIL.n176 B 0.014388f
C373 VTAIL.n177 B 0.987791f
C374 VTAIL.n178 B 0.013589f
C375 VTAIL.t9 B 0.053904f
C376 VTAIL.n179 B 0.157481f
C377 VTAIL.n180 B 0.022706f
C378 VTAIL.n181 B 0.024089f
C379 VTAIL.n182 B 0.032119f
C380 VTAIL.n183 B 0.014388f
C381 VTAIL.n184 B 0.013589f
C382 VTAIL.n185 B 0.025288f
C383 VTAIL.n186 B 0.025288f
C384 VTAIL.n187 B 0.013589f
C385 VTAIL.n188 B 0.014388f
C386 VTAIL.n189 B 0.032119f
C387 VTAIL.n190 B 0.032119f
C388 VTAIL.n191 B 0.014388f
C389 VTAIL.n192 B 0.013589f
C390 VTAIL.n193 B 0.025288f
C391 VTAIL.n194 B 0.025288f
C392 VTAIL.n195 B 0.013589f
C393 VTAIL.n196 B 0.013589f
C394 VTAIL.n197 B 0.014388f
C395 VTAIL.n198 B 0.032119f
C396 VTAIL.n199 B 0.032119f
C397 VTAIL.n200 B 0.032119f
C398 VTAIL.n201 B 0.013988f
C399 VTAIL.n202 B 0.013589f
C400 VTAIL.n203 B 0.025288f
C401 VTAIL.n204 B 0.025288f
C402 VTAIL.n205 B 0.013589f
C403 VTAIL.n206 B 0.014388f
C404 VTAIL.n207 B 0.032119f
C405 VTAIL.n208 B 0.070739f
C406 VTAIL.n209 B 0.014388f
C407 VTAIL.n210 B 0.013589f
C408 VTAIL.n211 B 0.065362f
C409 VTAIL.n212 B 0.039907f
C410 VTAIL.n213 B 1.23585f
C411 VTAIL.t2 B 0.188645f
C412 VTAIL.t5 B 0.188645f
C413 VTAIL.n214 B 1.5914f
C414 VTAIL.n215 B 0.356143f
C415 VDD1.n0 B 0.03339f
C416 VDD1.n1 B 0.023308f
C417 VDD1.n2 B 0.012525f
C418 VDD1.n3 B 0.029604f
C419 VDD1.n4 B 0.012893f
C420 VDD1.n5 B 0.023308f
C421 VDD1.n6 B 0.012893f
C422 VDD1.n7 B 0.012525f
C423 VDD1.n8 B 0.029604f
C424 VDD1.n9 B 0.029604f
C425 VDD1.n10 B 0.013261f
C426 VDD1.n11 B 0.023308f
C427 VDD1.n12 B 0.012525f
C428 VDD1.n13 B 0.029604f
C429 VDD1.n14 B 0.013261f
C430 VDD1.n15 B 0.910429f
C431 VDD1.n16 B 0.012525f
C432 VDD1.t3 B 0.049682f
C433 VDD1.n17 B 0.145148f
C434 VDD1.n18 B 0.020927f
C435 VDD1.n19 B 0.022203f
C436 VDD1.n20 B 0.029604f
C437 VDD1.n21 B 0.013261f
C438 VDD1.n22 B 0.012525f
C439 VDD1.n23 B 0.023308f
C440 VDD1.n24 B 0.023308f
C441 VDD1.n25 B 0.012525f
C442 VDD1.n26 B 0.013261f
C443 VDD1.n27 B 0.029604f
C444 VDD1.n28 B 0.029604f
C445 VDD1.n29 B 0.013261f
C446 VDD1.n30 B 0.012525f
C447 VDD1.n31 B 0.023308f
C448 VDD1.n32 B 0.023308f
C449 VDD1.n33 B 0.012525f
C450 VDD1.n34 B 0.013261f
C451 VDD1.n35 B 0.029604f
C452 VDD1.n36 B 0.029604f
C453 VDD1.n37 B 0.013261f
C454 VDD1.n38 B 0.012525f
C455 VDD1.n39 B 0.023308f
C456 VDD1.n40 B 0.023308f
C457 VDD1.n41 B 0.012525f
C458 VDD1.n42 B 0.013261f
C459 VDD1.n43 B 0.029604f
C460 VDD1.n44 B 0.065199f
C461 VDD1.n45 B 0.013261f
C462 VDD1.n46 B 0.012525f
C463 VDD1.n47 B 0.060243f
C464 VDD1.n48 B 0.056128f
C465 VDD1.t2 B 0.173871f
C466 VDD1.t0 B 0.173871f
C467 VDD1.n49 B 1.52725f
C468 VDD1.n50 B 0.447296f
C469 VDD1.n51 B 0.03339f
C470 VDD1.n52 B 0.023308f
C471 VDD1.n53 B 0.012525f
C472 VDD1.n54 B 0.029604f
C473 VDD1.n55 B 0.012893f
C474 VDD1.n56 B 0.023308f
C475 VDD1.n57 B 0.013261f
C476 VDD1.n58 B 0.029604f
C477 VDD1.n59 B 0.013261f
C478 VDD1.n60 B 0.023308f
C479 VDD1.n61 B 0.012525f
C480 VDD1.n62 B 0.029604f
C481 VDD1.n63 B 0.013261f
C482 VDD1.n64 B 0.910429f
C483 VDD1.n65 B 0.012525f
C484 VDD1.t1 B 0.049682f
C485 VDD1.n66 B 0.145148f
C486 VDD1.n67 B 0.020927f
C487 VDD1.n68 B 0.022203f
C488 VDD1.n69 B 0.029604f
C489 VDD1.n70 B 0.013261f
C490 VDD1.n71 B 0.012525f
C491 VDD1.n72 B 0.023308f
C492 VDD1.n73 B 0.023308f
C493 VDD1.n74 B 0.012525f
C494 VDD1.n75 B 0.013261f
C495 VDD1.n76 B 0.029604f
C496 VDD1.n77 B 0.029604f
C497 VDD1.n78 B 0.013261f
C498 VDD1.n79 B 0.012525f
C499 VDD1.n80 B 0.023308f
C500 VDD1.n81 B 0.023308f
C501 VDD1.n82 B 0.012525f
C502 VDD1.n83 B 0.012525f
C503 VDD1.n84 B 0.013261f
C504 VDD1.n85 B 0.029604f
C505 VDD1.n86 B 0.029604f
C506 VDD1.n87 B 0.029604f
C507 VDD1.n88 B 0.012893f
C508 VDD1.n89 B 0.012525f
C509 VDD1.n90 B 0.023308f
C510 VDD1.n91 B 0.023308f
C511 VDD1.n92 B 0.012525f
C512 VDD1.n93 B 0.013261f
C513 VDD1.n94 B 0.029604f
C514 VDD1.n95 B 0.065199f
C515 VDD1.n96 B 0.013261f
C516 VDD1.n97 B 0.012525f
C517 VDD1.n98 B 0.060243f
C518 VDD1.n99 B 0.056128f
C519 VDD1.t6 B 0.173871f
C520 VDD1.t9 B 0.173871f
C521 VDD1.n100 B 1.52724f
C522 VDD1.n101 B 0.440877f
C523 VDD1.t7 B 0.173871f
C524 VDD1.t4 B 0.173871f
C525 VDD1.n102 B 1.53188f
C526 VDD1.n103 B 1.91337f
C527 VDD1.t8 B 0.173871f
C528 VDD1.t5 B 0.173871f
C529 VDD1.n104 B 1.52724f
C530 VDD1.n105 B 2.19587f
C531 VP.n0 B 0.047848f
C532 VP.t0 B 1.02495f
C533 VP.n1 B 0.386983f
C534 VP.n2 B 0.035858f
C535 VP.t9 B 1.02495f
C536 VP.n3 B 0.049645f
C537 VP.n4 B 0.035858f
C538 VP.t7 B 1.02495f
C539 VP.t6 B 1.0861f
C540 VP.n5 B 0.449128f
C541 VP.n6 B 0.047848f
C542 VP.t4 B 1.0861f
C543 VP.t2 B 1.02495f
C544 VP.n7 B 0.386983f
C545 VP.n8 B 0.035858f
C546 VP.t8 B 1.02495f
C547 VP.n9 B 0.049645f
C548 VP.t3 B 1.12568f
C549 VP.n10 B 0.435594f
C550 VP.t5 B 1.02495f
C551 VP.n11 B 0.441837f
C552 VP.n12 B 0.051323f
C553 VP.n13 B 0.186827f
C554 VP.n14 B 0.035858f
C555 VP.n15 B 0.035858f
C556 VP.n16 B 0.420651f
C557 VP.n17 B 0.049645f
C558 VP.n18 B 0.051323f
C559 VP.n19 B 0.035858f
C560 VP.n20 B 0.035858f
C561 VP.n21 B 0.036951f
C562 VP.n22 B 0.042197f
C563 VP.n23 B 0.449128f
C564 VP.n24 B 1.5692f
C565 VP.n25 B 1.59905f
C566 VP.n26 B 0.047848f
C567 VP.n27 B 0.042197f
C568 VP.n28 B 0.036951f
C569 VP.n29 B 0.386983f
C570 VP.n30 B 0.051323f
C571 VP.n31 B 0.035858f
C572 VP.n32 B 0.035858f
C573 VP.n33 B 0.035858f
C574 VP.n34 B 0.420651f
C575 VP.n35 B 0.049645f
C576 VP.n36 B 0.051323f
C577 VP.n37 B 0.035858f
C578 VP.n38 B 0.035858f
C579 VP.n39 B 0.036951f
C580 VP.n40 B 0.042197f
C581 VP.t1 B 1.0861f
C582 VP.n41 B 0.449128f
C583 VP.n42 B 0.033582f
.ends

