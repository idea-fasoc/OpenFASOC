* NGSPICE file created from diff_pair_sample_0963.ext - technology: sky130A

.subckt diff_pair_sample_0963 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=6.3804 ps=33.5 w=16.36 l=1.85
X1 VDD2.t4 VN.t1 VTAIL.t9 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=2.6994 ps=16.69 w=16.36 l=1.85
X2 VTAIL.t8 VN.t2 VDD2.t3 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=2.6994 ps=16.69 w=16.36 l=1.85
X3 VDD2.t2 VN.t3 VTAIL.t7 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=6.3804 ps=33.5 w=16.36 l=1.85
X4 B.t11 B.t9 B.t10 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=0 ps=0 w=16.36 l=1.85
X5 VTAIL.t10 VN.t4 VDD2.t1 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=2.6994 ps=16.69 w=16.36 l=1.85
X6 VDD1.t5 VP.t0 VTAIL.t1 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=6.3804 ps=33.5 w=16.36 l=1.85
X7 B.t8 B.t6 B.t7 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=0 ps=0 w=16.36 l=1.85
X8 B.t5 B.t3 B.t4 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=0 ps=0 w=16.36 l=1.85
X9 VTAIL.t3 VP.t1 VDD1.t4 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=2.6994 ps=16.69 w=16.36 l=1.85
X10 VDD1.t3 VP.t2 VTAIL.t0 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=2.6994 ps=16.69 w=16.36 l=1.85
X11 B.t2 B.t0 B.t1 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=0 ps=0 w=16.36 l=1.85
X12 VDD1.t2 VP.t3 VTAIL.t2 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=2.6994 ps=16.69 w=16.36 l=1.85
X13 VDD2.t0 VN.t5 VTAIL.t11 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=6.3804 pd=33.5 as=2.6994 ps=16.69 w=16.36 l=1.85
X14 VDD1.t1 VP.t4 VTAIL.t4 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=6.3804 ps=33.5 w=16.36 l=1.85
X15 VTAIL.t5 VP.t5 VDD1.t0 w_n2714_n4240# sky130_fd_pr__pfet_01v8 ad=2.6994 pd=16.69 as=2.6994 ps=16.69 w=16.36 l=1.85
R0 VN.n2 VN.t1 243.796
R1 VN.n14 VN.t3 243.796
R2 VN.n3 VN.t2 213.123
R3 VN.n10 VN.t0 213.123
R4 VN.n15 VN.t4 213.123
R5 VN.n22 VN.t5 213.123
R6 VN.n21 VN.n12 161.3
R7 VN.n20 VN.n19 161.3
R8 VN.n18 VN.n13 161.3
R9 VN.n17 VN.n16 161.3
R10 VN.n9 VN.n0 161.3
R11 VN.n8 VN.n7 161.3
R12 VN.n6 VN.n1 161.3
R13 VN.n5 VN.n4 161.3
R14 VN.n11 VN.n10 89.7593
R15 VN.n23 VN.n22 89.7593
R16 VN.n3 VN.n2 57.8394
R17 VN.n15 VN.n14 57.8394
R18 VN.n8 VN.n1 56.0773
R19 VN.n20 VN.n13 56.0773
R20 VN VN.n23 49.3239
R21 VN.n9 VN.n8 25.0767
R22 VN.n21 VN.n20 25.0767
R23 VN.n4 VN.n1 24.5923
R24 VN.n16 VN.n13 24.5923
R25 VN.n10 VN.n9 21.1495
R26 VN.n22 VN.n21 21.1495
R27 VN.n17 VN.n14 13.1274
R28 VN.n5 VN.n2 13.1274
R29 VN.n4 VN.n3 12.2964
R30 VN.n16 VN.n15 12.2964
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n7 VTAIL.t7 53.348
R41 VTAIL.n11 VTAIL.t6 53.3478
R42 VTAIL.n2 VTAIL.t1 53.3478
R43 VTAIL.n10 VTAIL.t4 53.3478
R44 VTAIL.n9 VTAIL.n8 51.3612
R45 VTAIL.n6 VTAIL.n5 51.3612
R46 VTAIL.n1 VTAIL.n0 51.3609
R47 VTAIL.n4 VTAIL.n3 51.3609
R48 VTAIL.n6 VTAIL.n4 30.2289
R49 VTAIL.n11 VTAIL.n10 28.3496
R50 VTAIL.n0 VTAIL.t9 1.98736
R51 VTAIL.n0 VTAIL.t8 1.98736
R52 VTAIL.n3 VTAIL.t0 1.98736
R53 VTAIL.n3 VTAIL.t3 1.98736
R54 VTAIL.n8 VTAIL.t2 1.98736
R55 VTAIL.n8 VTAIL.t5 1.98736
R56 VTAIL.n5 VTAIL.t11 1.98736
R57 VTAIL.n5 VTAIL.t10 1.98736
R58 VTAIL.n7 VTAIL.n6 1.87981
R59 VTAIL.n10 VTAIL.n9 1.87981
R60 VTAIL.n4 VTAIL.n2 1.87981
R61 VTAIL.n9 VTAIL.n7 1.40998
R62 VTAIL.n2 VTAIL.n1 1.40998
R63 VTAIL VTAIL.n11 1.35179
R64 VTAIL VTAIL.n1 0.528517
R65 VDD2.n1 VDD2.t4 71.3807
R66 VDD2.n2 VDD2.t0 70.0268
R67 VDD2.n1 VDD2.n0 68.4542
R68 VDD2 VDD2.n3 68.4514
R69 VDD2.n2 VDD2.n1 43.9265
R70 VDD2.n3 VDD2.t1 1.98736
R71 VDD2.n3 VDD2.t2 1.98736
R72 VDD2.n0 VDD2.t3 1.98736
R73 VDD2.n0 VDD2.t5 1.98736
R74 VDD2 VDD2.n2 1.46817
R75 B.n422 B.n421 585
R76 B.n420 B.n117 585
R77 B.n419 B.n418 585
R78 B.n417 B.n118 585
R79 B.n416 B.n415 585
R80 B.n414 B.n119 585
R81 B.n413 B.n412 585
R82 B.n411 B.n120 585
R83 B.n410 B.n409 585
R84 B.n408 B.n121 585
R85 B.n407 B.n406 585
R86 B.n405 B.n122 585
R87 B.n404 B.n403 585
R88 B.n402 B.n123 585
R89 B.n401 B.n400 585
R90 B.n399 B.n124 585
R91 B.n398 B.n397 585
R92 B.n396 B.n125 585
R93 B.n395 B.n394 585
R94 B.n393 B.n126 585
R95 B.n392 B.n391 585
R96 B.n390 B.n127 585
R97 B.n389 B.n388 585
R98 B.n387 B.n128 585
R99 B.n386 B.n385 585
R100 B.n384 B.n129 585
R101 B.n383 B.n382 585
R102 B.n381 B.n130 585
R103 B.n380 B.n379 585
R104 B.n378 B.n131 585
R105 B.n377 B.n376 585
R106 B.n375 B.n132 585
R107 B.n374 B.n373 585
R108 B.n372 B.n133 585
R109 B.n371 B.n370 585
R110 B.n369 B.n134 585
R111 B.n368 B.n367 585
R112 B.n366 B.n135 585
R113 B.n365 B.n364 585
R114 B.n363 B.n136 585
R115 B.n362 B.n361 585
R116 B.n360 B.n137 585
R117 B.n359 B.n358 585
R118 B.n357 B.n138 585
R119 B.n356 B.n355 585
R120 B.n354 B.n139 585
R121 B.n353 B.n352 585
R122 B.n351 B.n140 585
R123 B.n350 B.n349 585
R124 B.n348 B.n141 585
R125 B.n347 B.n346 585
R126 B.n345 B.n142 585
R127 B.n344 B.n343 585
R128 B.n342 B.n143 585
R129 B.n341 B.n340 585
R130 B.n336 B.n144 585
R131 B.n335 B.n334 585
R132 B.n333 B.n145 585
R133 B.n332 B.n331 585
R134 B.n330 B.n146 585
R135 B.n329 B.n328 585
R136 B.n327 B.n147 585
R137 B.n326 B.n325 585
R138 B.n324 B.n148 585
R139 B.n322 B.n321 585
R140 B.n320 B.n151 585
R141 B.n319 B.n318 585
R142 B.n317 B.n152 585
R143 B.n316 B.n315 585
R144 B.n314 B.n153 585
R145 B.n313 B.n312 585
R146 B.n311 B.n154 585
R147 B.n310 B.n309 585
R148 B.n308 B.n155 585
R149 B.n307 B.n306 585
R150 B.n305 B.n156 585
R151 B.n304 B.n303 585
R152 B.n302 B.n157 585
R153 B.n301 B.n300 585
R154 B.n299 B.n158 585
R155 B.n298 B.n297 585
R156 B.n296 B.n159 585
R157 B.n295 B.n294 585
R158 B.n293 B.n160 585
R159 B.n292 B.n291 585
R160 B.n290 B.n161 585
R161 B.n289 B.n288 585
R162 B.n287 B.n162 585
R163 B.n286 B.n285 585
R164 B.n284 B.n163 585
R165 B.n283 B.n282 585
R166 B.n281 B.n164 585
R167 B.n280 B.n279 585
R168 B.n278 B.n165 585
R169 B.n277 B.n276 585
R170 B.n275 B.n166 585
R171 B.n274 B.n273 585
R172 B.n272 B.n167 585
R173 B.n271 B.n270 585
R174 B.n269 B.n168 585
R175 B.n268 B.n267 585
R176 B.n266 B.n169 585
R177 B.n265 B.n264 585
R178 B.n263 B.n170 585
R179 B.n262 B.n261 585
R180 B.n260 B.n171 585
R181 B.n259 B.n258 585
R182 B.n257 B.n172 585
R183 B.n256 B.n255 585
R184 B.n254 B.n173 585
R185 B.n253 B.n252 585
R186 B.n251 B.n174 585
R187 B.n250 B.n249 585
R188 B.n248 B.n175 585
R189 B.n247 B.n246 585
R190 B.n245 B.n176 585
R191 B.n244 B.n243 585
R192 B.n242 B.n177 585
R193 B.n423 B.n116 585
R194 B.n425 B.n424 585
R195 B.n426 B.n115 585
R196 B.n428 B.n427 585
R197 B.n429 B.n114 585
R198 B.n431 B.n430 585
R199 B.n432 B.n113 585
R200 B.n434 B.n433 585
R201 B.n435 B.n112 585
R202 B.n437 B.n436 585
R203 B.n438 B.n111 585
R204 B.n440 B.n439 585
R205 B.n441 B.n110 585
R206 B.n443 B.n442 585
R207 B.n444 B.n109 585
R208 B.n446 B.n445 585
R209 B.n447 B.n108 585
R210 B.n449 B.n448 585
R211 B.n450 B.n107 585
R212 B.n452 B.n451 585
R213 B.n453 B.n106 585
R214 B.n455 B.n454 585
R215 B.n456 B.n105 585
R216 B.n458 B.n457 585
R217 B.n459 B.n104 585
R218 B.n461 B.n460 585
R219 B.n462 B.n103 585
R220 B.n464 B.n463 585
R221 B.n465 B.n102 585
R222 B.n467 B.n466 585
R223 B.n468 B.n101 585
R224 B.n470 B.n469 585
R225 B.n471 B.n100 585
R226 B.n473 B.n472 585
R227 B.n474 B.n99 585
R228 B.n476 B.n475 585
R229 B.n477 B.n98 585
R230 B.n479 B.n478 585
R231 B.n480 B.n97 585
R232 B.n482 B.n481 585
R233 B.n483 B.n96 585
R234 B.n485 B.n484 585
R235 B.n486 B.n95 585
R236 B.n488 B.n487 585
R237 B.n489 B.n94 585
R238 B.n491 B.n490 585
R239 B.n492 B.n93 585
R240 B.n494 B.n493 585
R241 B.n495 B.n92 585
R242 B.n497 B.n496 585
R243 B.n498 B.n91 585
R244 B.n500 B.n499 585
R245 B.n501 B.n90 585
R246 B.n503 B.n502 585
R247 B.n504 B.n89 585
R248 B.n506 B.n505 585
R249 B.n507 B.n88 585
R250 B.n509 B.n508 585
R251 B.n510 B.n87 585
R252 B.n512 B.n511 585
R253 B.n513 B.n86 585
R254 B.n515 B.n514 585
R255 B.n516 B.n85 585
R256 B.n518 B.n517 585
R257 B.n519 B.n84 585
R258 B.n521 B.n520 585
R259 B.n522 B.n83 585
R260 B.n524 B.n523 585
R261 B.n702 B.n701 585
R262 B.n700 B.n19 585
R263 B.n699 B.n698 585
R264 B.n697 B.n20 585
R265 B.n696 B.n695 585
R266 B.n694 B.n21 585
R267 B.n693 B.n692 585
R268 B.n691 B.n22 585
R269 B.n690 B.n689 585
R270 B.n688 B.n23 585
R271 B.n687 B.n686 585
R272 B.n685 B.n24 585
R273 B.n684 B.n683 585
R274 B.n682 B.n25 585
R275 B.n681 B.n680 585
R276 B.n679 B.n26 585
R277 B.n678 B.n677 585
R278 B.n676 B.n27 585
R279 B.n675 B.n674 585
R280 B.n673 B.n28 585
R281 B.n672 B.n671 585
R282 B.n670 B.n29 585
R283 B.n669 B.n668 585
R284 B.n667 B.n30 585
R285 B.n666 B.n665 585
R286 B.n664 B.n31 585
R287 B.n663 B.n662 585
R288 B.n661 B.n32 585
R289 B.n660 B.n659 585
R290 B.n658 B.n33 585
R291 B.n657 B.n656 585
R292 B.n655 B.n34 585
R293 B.n654 B.n653 585
R294 B.n652 B.n35 585
R295 B.n651 B.n650 585
R296 B.n649 B.n36 585
R297 B.n648 B.n647 585
R298 B.n646 B.n37 585
R299 B.n645 B.n644 585
R300 B.n643 B.n38 585
R301 B.n642 B.n641 585
R302 B.n640 B.n39 585
R303 B.n639 B.n638 585
R304 B.n637 B.n40 585
R305 B.n636 B.n635 585
R306 B.n634 B.n41 585
R307 B.n633 B.n632 585
R308 B.n631 B.n42 585
R309 B.n630 B.n629 585
R310 B.n628 B.n43 585
R311 B.n627 B.n626 585
R312 B.n625 B.n44 585
R313 B.n624 B.n623 585
R314 B.n622 B.n45 585
R315 B.n620 B.n619 585
R316 B.n618 B.n48 585
R317 B.n617 B.n616 585
R318 B.n615 B.n49 585
R319 B.n614 B.n613 585
R320 B.n612 B.n50 585
R321 B.n611 B.n610 585
R322 B.n609 B.n51 585
R323 B.n608 B.n607 585
R324 B.n606 B.n52 585
R325 B.n605 B.n604 585
R326 B.n603 B.n53 585
R327 B.n602 B.n601 585
R328 B.n600 B.n57 585
R329 B.n599 B.n598 585
R330 B.n597 B.n58 585
R331 B.n596 B.n595 585
R332 B.n594 B.n59 585
R333 B.n593 B.n592 585
R334 B.n591 B.n60 585
R335 B.n590 B.n589 585
R336 B.n588 B.n61 585
R337 B.n587 B.n586 585
R338 B.n585 B.n62 585
R339 B.n584 B.n583 585
R340 B.n582 B.n63 585
R341 B.n581 B.n580 585
R342 B.n579 B.n64 585
R343 B.n578 B.n577 585
R344 B.n576 B.n65 585
R345 B.n575 B.n574 585
R346 B.n573 B.n66 585
R347 B.n572 B.n571 585
R348 B.n570 B.n67 585
R349 B.n569 B.n568 585
R350 B.n567 B.n68 585
R351 B.n566 B.n565 585
R352 B.n564 B.n69 585
R353 B.n563 B.n562 585
R354 B.n561 B.n70 585
R355 B.n560 B.n559 585
R356 B.n558 B.n71 585
R357 B.n557 B.n556 585
R358 B.n555 B.n72 585
R359 B.n554 B.n553 585
R360 B.n552 B.n73 585
R361 B.n551 B.n550 585
R362 B.n549 B.n74 585
R363 B.n548 B.n547 585
R364 B.n546 B.n75 585
R365 B.n545 B.n544 585
R366 B.n543 B.n76 585
R367 B.n542 B.n541 585
R368 B.n540 B.n77 585
R369 B.n539 B.n538 585
R370 B.n537 B.n78 585
R371 B.n536 B.n535 585
R372 B.n534 B.n79 585
R373 B.n533 B.n532 585
R374 B.n531 B.n80 585
R375 B.n530 B.n529 585
R376 B.n528 B.n81 585
R377 B.n527 B.n526 585
R378 B.n525 B.n82 585
R379 B.n703 B.n18 585
R380 B.n705 B.n704 585
R381 B.n706 B.n17 585
R382 B.n708 B.n707 585
R383 B.n709 B.n16 585
R384 B.n711 B.n710 585
R385 B.n712 B.n15 585
R386 B.n714 B.n713 585
R387 B.n715 B.n14 585
R388 B.n717 B.n716 585
R389 B.n718 B.n13 585
R390 B.n720 B.n719 585
R391 B.n721 B.n12 585
R392 B.n723 B.n722 585
R393 B.n724 B.n11 585
R394 B.n726 B.n725 585
R395 B.n727 B.n10 585
R396 B.n729 B.n728 585
R397 B.n730 B.n9 585
R398 B.n732 B.n731 585
R399 B.n733 B.n8 585
R400 B.n735 B.n734 585
R401 B.n736 B.n7 585
R402 B.n738 B.n737 585
R403 B.n739 B.n6 585
R404 B.n741 B.n740 585
R405 B.n742 B.n5 585
R406 B.n744 B.n743 585
R407 B.n745 B.n4 585
R408 B.n747 B.n746 585
R409 B.n748 B.n3 585
R410 B.n750 B.n749 585
R411 B.n751 B.n0 585
R412 B.n2 B.n1 585
R413 B.n194 B.n193 585
R414 B.n196 B.n195 585
R415 B.n197 B.n192 585
R416 B.n199 B.n198 585
R417 B.n200 B.n191 585
R418 B.n202 B.n201 585
R419 B.n203 B.n190 585
R420 B.n205 B.n204 585
R421 B.n206 B.n189 585
R422 B.n208 B.n207 585
R423 B.n209 B.n188 585
R424 B.n211 B.n210 585
R425 B.n212 B.n187 585
R426 B.n214 B.n213 585
R427 B.n215 B.n186 585
R428 B.n217 B.n216 585
R429 B.n218 B.n185 585
R430 B.n220 B.n219 585
R431 B.n221 B.n184 585
R432 B.n223 B.n222 585
R433 B.n224 B.n183 585
R434 B.n226 B.n225 585
R435 B.n227 B.n182 585
R436 B.n229 B.n228 585
R437 B.n230 B.n181 585
R438 B.n232 B.n231 585
R439 B.n233 B.n180 585
R440 B.n235 B.n234 585
R441 B.n236 B.n179 585
R442 B.n238 B.n237 585
R443 B.n239 B.n178 585
R444 B.n241 B.n240 585
R445 B.n242 B.n241 578.989
R446 B.n421 B.n116 578.989
R447 B.n523 B.n82 578.989
R448 B.n703 B.n702 578.989
R449 B.n149 B.t3 419.664
R450 B.n337 B.t9 419.664
R451 B.n54 B.t0 419.664
R452 B.n46 B.t6 419.664
R453 B.n753 B.n752 256.663
R454 B.n752 B.n751 235.042
R455 B.n752 B.n2 235.042
R456 B.n243 B.n242 163.367
R457 B.n243 B.n176 163.367
R458 B.n247 B.n176 163.367
R459 B.n248 B.n247 163.367
R460 B.n249 B.n248 163.367
R461 B.n249 B.n174 163.367
R462 B.n253 B.n174 163.367
R463 B.n254 B.n253 163.367
R464 B.n255 B.n254 163.367
R465 B.n255 B.n172 163.367
R466 B.n259 B.n172 163.367
R467 B.n260 B.n259 163.367
R468 B.n261 B.n260 163.367
R469 B.n261 B.n170 163.367
R470 B.n265 B.n170 163.367
R471 B.n266 B.n265 163.367
R472 B.n267 B.n266 163.367
R473 B.n267 B.n168 163.367
R474 B.n271 B.n168 163.367
R475 B.n272 B.n271 163.367
R476 B.n273 B.n272 163.367
R477 B.n273 B.n166 163.367
R478 B.n277 B.n166 163.367
R479 B.n278 B.n277 163.367
R480 B.n279 B.n278 163.367
R481 B.n279 B.n164 163.367
R482 B.n283 B.n164 163.367
R483 B.n284 B.n283 163.367
R484 B.n285 B.n284 163.367
R485 B.n285 B.n162 163.367
R486 B.n289 B.n162 163.367
R487 B.n290 B.n289 163.367
R488 B.n291 B.n290 163.367
R489 B.n291 B.n160 163.367
R490 B.n295 B.n160 163.367
R491 B.n296 B.n295 163.367
R492 B.n297 B.n296 163.367
R493 B.n297 B.n158 163.367
R494 B.n301 B.n158 163.367
R495 B.n302 B.n301 163.367
R496 B.n303 B.n302 163.367
R497 B.n303 B.n156 163.367
R498 B.n307 B.n156 163.367
R499 B.n308 B.n307 163.367
R500 B.n309 B.n308 163.367
R501 B.n309 B.n154 163.367
R502 B.n313 B.n154 163.367
R503 B.n314 B.n313 163.367
R504 B.n315 B.n314 163.367
R505 B.n315 B.n152 163.367
R506 B.n319 B.n152 163.367
R507 B.n320 B.n319 163.367
R508 B.n321 B.n320 163.367
R509 B.n321 B.n148 163.367
R510 B.n326 B.n148 163.367
R511 B.n327 B.n326 163.367
R512 B.n328 B.n327 163.367
R513 B.n328 B.n146 163.367
R514 B.n332 B.n146 163.367
R515 B.n333 B.n332 163.367
R516 B.n334 B.n333 163.367
R517 B.n334 B.n144 163.367
R518 B.n341 B.n144 163.367
R519 B.n342 B.n341 163.367
R520 B.n343 B.n342 163.367
R521 B.n343 B.n142 163.367
R522 B.n347 B.n142 163.367
R523 B.n348 B.n347 163.367
R524 B.n349 B.n348 163.367
R525 B.n349 B.n140 163.367
R526 B.n353 B.n140 163.367
R527 B.n354 B.n353 163.367
R528 B.n355 B.n354 163.367
R529 B.n355 B.n138 163.367
R530 B.n359 B.n138 163.367
R531 B.n360 B.n359 163.367
R532 B.n361 B.n360 163.367
R533 B.n361 B.n136 163.367
R534 B.n365 B.n136 163.367
R535 B.n366 B.n365 163.367
R536 B.n367 B.n366 163.367
R537 B.n367 B.n134 163.367
R538 B.n371 B.n134 163.367
R539 B.n372 B.n371 163.367
R540 B.n373 B.n372 163.367
R541 B.n373 B.n132 163.367
R542 B.n377 B.n132 163.367
R543 B.n378 B.n377 163.367
R544 B.n379 B.n378 163.367
R545 B.n379 B.n130 163.367
R546 B.n383 B.n130 163.367
R547 B.n384 B.n383 163.367
R548 B.n385 B.n384 163.367
R549 B.n385 B.n128 163.367
R550 B.n389 B.n128 163.367
R551 B.n390 B.n389 163.367
R552 B.n391 B.n390 163.367
R553 B.n391 B.n126 163.367
R554 B.n395 B.n126 163.367
R555 B.n396 B.n395 163.367
R556 B.n397 B.n396 163.367
R557 B.n397 B.n124 163.367
R558 B.n401 B.n124 163.367
R559 B.n402 B.n401 163.367
R560 B.n403 B.n402 163.367
R561 B.n403 B.n122 163.367
R562 B.n407 B.n122 163.367
R563 B.n408 B.n407 163.367
R564 B.n409 B.n408 163.367
R565 B.n409 B.n120 163.367
R566 B.n413 B.n120 163.367
R567 B.n414 B.n413 163.367
R568 B.n415 B.n414 163.367
R569 B.n415 B.n118 163.367
R570 B.n419 B.n118 163.367
R571 B.n420 B.n419 163.367
R572 B.n421 B.n420 163.367
R573 B.n523 B.n522 163.367
R574 B.n522 B.n521 163.367
R575 B.n521 B.n84 163.367
R576 B.n517 B.n84 163.367
R577 B.n517 B.n516 163.367
R578 B.n516 B.n515 163.367
R579 B.n515 B.n86 163.367
R580 B.n511 B.n86 163.367
R581 B.n511 B.n510 163.367
R582 B.n510 B.n509 163.367
R583 B.n509 B.n88 163.367
R584 B.n505 B.n88 163.367
R585 B.n505 B.n504 163.367
R586 B.n504 B.n503 163.367
R587 B.n503 B.n90 163.367
R588 B.n499 B.n90 163.367
R589 B.n499 B.n498 163.367
R590 B.n498 B.n497 163.367
R591 B.n497 B.n92 163.367
R592 B.n493 B.n92 163.367
R593 B.n493 B.n492 163.367
R594 B.n492 B.n491 163.367
R595 B.n491 B.n94 163.367
R596 B.n487 B.n94 163.367
R597 B.n487 B.n486 163.367
R598 B.n486 B.n485 163.367
R599 B.n485 B.n96 163.367
R600 B.n481 B.n96 163.367
R601 B.n481 B.n480 163.367
R602 B.n480 B.n479 163.367
R603 B.n479 B.n98 163.367
R604 B.n475 B.n98 163.367
R605 B.n475 B.n474 163.367
R606 B.n474 B.n473 163.367
R607 B.n473 B.n100 163.367
R608 B.n469 B.n100 163.367
R609 B.n469 B.n468 163.367
R610 B.n468 B.n467 163.367
R611 B.n467 B.n102 163.367
R612 B.n463 B.n102 163.367
R613 B.n463 B.n462 163.367
R614 B.n462 B.n461 163.367
R615 B.n461 B.n104 163.367
R616 B.n457 B.n104 163.367
R617 B.n457 B.n456 163.367
R618 B.n456 B.n455 163.367
R619 B.n455 B.n106 163.367
R620 B.n451 B.n106 163.367
R621 B.n451 B.n450 163.367
R622 B.n450 B.n449 163.367
R623 B.n449 B.n108 163.367
R624 B.n445 B.n108 163.367
R625 B.n445 B.n444 163.367
R626 B.n444 B.n443 163.367
R627 B.n443 B.n110 163.367
R628 B.n439 B.n110 163.367
R629 B.n439 B.n438 163.367
R630 B.n438 B.n437 163.367
R631 B.n437 B.n112 163.367
R632 B.n433 B.n112 163.367
R633 B.n433 B.n432 163.367
R634 B.n432 B.n431 163.367
R635 B.n431 B.n114 163.367
R636 B.n427 B.n114 163.367
R637 B.n427 B.n426 163.367
R638 B.n426 B.n425 163.367
R639 B.n425 B.n116 163.367
R640 B.n702 B.n19 163.367
R641 B.n698 B.n19 163.367
R642 B.n698 B.n697 163.367
R643 B.n697 B.n696 163.367
R644 B.n696 B.n21 163.367
R645 B.n692 B.n21 163.367
R646 B.n692 B.n691 163.367
R647 B.n691 B.n690 163.367
R648 B.n690 B.n23 163.367
R649 B.n686 B.n23 163.367
R650 B.n686 B.n685 163.367
R651 B.n685 B.n684 163.367
R652 B.n684 B.n25 163.367
R653 B.n680 B.n25 163.367
R654 B.n680 B.n679 163.367
R655 B.n679 B.n678 163.367
R656 B.n678 B.n27 163.367
R657 B.n674 B.n27 163.367
R658 B.n674 B.n673 163.367
R659 B.n673 B.n672 163.367
R660 B.n672 B.n29 163.367
R661 B.n668 B.n29 163.367
R662 B.n668 B.n667 163.367
R663 B.n667 B.n666 163.367
R664 B.n666 B.n31 163.367
R665 B.n662 B.n31 163.367
R666 B.n662 B.n661 163.367
R667 B.n661 B.n660 163.367
R668 B.n660 B.n33 163.367
R669 B.n656 B.n33 163.367
R670 B.n656 B.n655 163.367
R671 B.n655 B.n654 163.367
R672 B.n654 B.n35 163.367
R673 B.n650 B.n35 163.367
R674 B.n650 B.n649 163.367
R675 B.n649 B.n648 163.367
R676 B.n648 B.n37 163.367
R677 B.n644 B.n37 163.367
R678 B.n644 B.n643 163.367
R679 B.n643 B.n642 163.367
R680 B.n642 B.n39 163.367
R681 B.n638 B.n39 163.367
R682 B.n638 B.n637 163.367
R683 B.n637 B.n636 163.367
R684 B.n636 B.n41 163.367
R685 B.n632 B.n41 163.367
R686 B.n632 B.n631 163.367
R687 B.n631 B.n630 163.367
R688 B.n630 B.n43 163.367
R689 B.n626 B.n43 163.367
R690 B.n626 B.n625 163.367
R691 B.n625 B.n624 163.367
R692 B.n624 B.n45 163.367
R693 B.n619 B.n45 163.367
R694 B.n619 B.n618 163.367
R695 B.n618 B.n617 163.367
R696 B.n617 B.n49 163.367
R697 B.n613 B.n49 163.367
R698 B.n613 B.n612 163.367
R699 B.n612 B.n611 163.367
R700 B.n611 B.n51 163.367
R701 B.n607 B.n51 163.367
R702 B.n607 B.n606 163.367
R703 B.n606 B.n605 163.367
R704 B.n605 B.n53 163.367
R705 B.n601 B.n53 163.367
R706 B.n601 B.n600 163.367
R707 B.n600 B.n599 163.367
R708 B.n599 B.n58 163.367
R709 B.n595 B.n58 163.367
R710 B.n595 B.n594 163.367
R711 B.n594 B.n593 163.367
R712 B.n593 B.n60 163.367
R713 B.n589 B.n60 163.367
R714 B.n589 B.n588 163.367
R715 B.n588 B.n587 163.367
R716 B.n587 B.n62 163.367
R717 B.n583 B.n62 163.367
R718 B.n583 B.n582 163.367
R719 B.n582 B.n581 163.367
R720 B.n581 B.n64 163.367
R721 B.n577 B.n64 163.367
R722 B.n577 B.n576 163.367
R723 B.n576 B.n575 163.367
R724 B.n575 B.n66 163.367
R725 B.n571 B.n66 163.367
R726 B.n571 B.n570 163.367
R727 B.n570 B.n569 163.367
R728 B.n569 B.n68 163.367
R729 B.n565 B.n68 163.367
R730 B.n565 B.n564 163.367
R731 B.n564 B.n563 163.367
R732 B.n563 B.n70 163.367
R733 B.n559 B.n70 163.367
R734 B.n559 B.n558 163.367
R735 B.n558 B.n557 163.367
R736 B.n557 B.n72 163.367
R737 B.n553 B.n72 163.367
R738 B.n553 B.n552 163.367
R739 B.n552 B.n551 163.367
R740 B.n551 B.n74 163.367
R741 B.n547 B.n74 163.367
R742 B.n547 B.n546 163.367
R743 B.n546 B.n545 163.367
R744 B.n545 B.n76 163.367
R745 B.n541 B.n76 163.367
R746 B.n541 B.n540 163.367
R747 B.n540 B.n539 163.367
R748 B.n539 B.n78 163.367
R749 B.n535 B.n78 163.367
R750 B.n535 B.n534 163.367
R751 B.n534 B.n533 163.367
R752 B.n533 B.n80 163.367
R753 B.n529 B.n80 163.367
R754 B.n529 B.n528 163.367
R755 B.n528 B.n527 163.367
R756 B.n527 B.n82 163.367
R757 B.n704 B.n703 163.367
R758 B.n704 B.n17 163.367
R759 B.n708 B.n17 163.367
R760 B.n709 B.n708 163.367
R761 B.n710 B.n709 163.367
R762 B.n710 B.n15 163.367
R763 B.n714 B.n15 163.367
R764 B.n715 B.n714 163.367
R765 B.n716 B.n715 163.367
R766 B.n716 B.n13 163.367
R767 B.n720 B.n13 163.367
R768 B.n721 B.n720 163.367
R769 B.n722 B.n721 163.367
R770 B.n722 B.n11 163.367
R771 B.n726 B.n11 163.367
R772 B.n727 B.n726 163.367
R773 B.n728 B.n727 163.367
R774 B.n728 B.n9 163.367
R775 B.n732 B.n9 163.367
R776 B.n733 B.n732 163.367
R777 B.n734 B.n733 163.367
R778 B.n734 B.n7 163.367
R779 B.n738 B.n7 163.367
R780 B.n739 B.n738 163.367
R781 B.n740 B.n739 163.367
R782 B.n740 B.n5 163.367
R783 B.n744 B.n5 163.367
R784 B.n745 B.n744 163.367
R785 B.n746 B.n745 163.367
R786 B.n746 B.n3 163.367
R787 B.n750 B.n3 163.367
R788 B.n751 B.n750 163.367
R789 B.n194 B.n2 163.367
R790 B.n195 B.n194 163.367
R791 B.n195 B.n192 163.367
R792 B.n199 B.n192 163.367
R793 B.n200 B.n199 163.367
R794 B.n201 B.n200 163.367
R795 B.n201 B.n190 163.367
R796 B.n205 B.n190 163.367
R797 B.n206 B.n205 163.367
R798 B.n207 B.n206 163.367
R799 B.n207 B.n188 163.367
R800 B.n211 B.n188 163.367
R801 B.n212 B.n211 163.367
R802 B.n213 B.n212 163.367
R803 B.n213 B.n186 163.367
R804 B.n217 B.n186 163.367
R805 B.n218 B.n217 163.367
R806 B.n219 B.n218 163.367
R807 B.n219 B.n184 163.367
R808 B.n223 B.n184 163.367
R809 B.n224 B.n223 163.367
R810 B.n225 B.n224 163.367
R811 B.n225 B.n182 163.367
R812 B.n229 B.n182 163.367
R813 B.n230 B.n229 163.367
R814 B.n231 B.n230 163.367
R815 B.n231 B.n180 163.367
R816 B.n235 B.n180 163.367
R817 B.n236 B.n235 163.367
R818 B.n237 B.n236 163.367
R819 B.n237 B.n178 163.367
R820 B.n241 B.n178 163.367
R821 B.n337 B.t10 149.438
R822 B.n54 B.t2 149.438
R823 B.n149 B.t4 149.417
R824 B.n46 B.t8 149.417
R825 B.n338 B.t11 107.159
R826 B.n55 B.t1 107.159
R827 B.n150 B.t5 107.138
R828 B.n47 B.t7 107.138
R829 B.n323 B.n150 59.5399
R830 B.n339 B.n338 59.5399
R831 B.n56 B.n55 59.5399
R832 B.n621 B.n47 59.5399
R833 B.n150 B.n149 42.2793
R834 B.n338 B.n337 42.2793
R835 B.n55 B.n54 42.2793
R836 B.n47 B.n46 42.2793
R837 B.n701 B.n18 37.62
R838 B.n525 B.n524 37.62
R839 B.n423 B.n422 37.62
R840 B.n240 B.n177 37.62
R841 B B.n753 18.0485
R842 B.n705 B.n18 10.6151
R843 B.n706 B.n705 10.6151
R844 B.n707 B.n706 10.6151
R845 B.n707 B.n16 10.6151
R846 B.n711 B.n16 10.6151
R847 B.n712 B.n711 10.6151
R848 B.n713 B.n712 10.6151
R849 B.n713 B.n14 10.6151
R850 B.n717 B.n14 10.6151
R851 B.n718 B.n717 10.6151
R852 B.n719 B.n718 10.6151
R853 B.n719 B.n12 10.6151
R854 B.n723 B.n12 10.6151
R855 B.n724 B.n723 10.6151
R856 B.n725 B.n724 10.6151
R857 B.n725 B.n10 10.6151
R858 B.n729 B.n10 10.6151
R859 B.n730 B.n729 10.6151
R860 B.n731 B.n730 10.6151
R861 B.n731 B.n8 10.6151
R862 B.n735 B.n8 10.6151
R863 B.n736 B.n735 10.6151
R864 B.n737 B.n736 10.6151
R865 B.n737 B.n6 10.6151
R866 B.n741 B.n6 10.6151
R867 B.n742 B.n741 10.6151
R868 B.n743 B.n742 10.6151
R869 B.n743 B.n4 10.6151
R870 B.n747 B.n4 10.6151
R871 B.n748 B.n747 10.6151
R872 B.n749 B.n748 10.6151
R873 B.n749 B.n0 10.6151
R874 B.n701 B.n700 10.6151
R875 B.n700 B.n699 10.6151
R876 B.n699 B.n20 10.6151
R877 B.n695 B.n20 10.6151
R878 B.n695 B.n694 10.6151
R879 B.n694 B.n693 10.6151
R880 B.n693 B.n22 10.6151
R881 B.n689 B.n22 10.6151
R882 B.n689 B.n688 10.6151
R883 B.n688 B.n687 10.6151
R884 B.n687 B.n24 10.6151
R885 B.n683 B.n24 10.6151
R886 B.n683 B.n682 10.6151
R887 B.n682 B.n681 10.6151
R888 B.n681 B.n26 10.6151
R889 B.n677 B.n26 10.6151
R890 B.n677 B.n676 10.6151
R891 B.n676 B.n675 10.6151
R892 B.n675 B.n28 10.6151
R893 B.n671 B.n28 10.6151
R894 B.n671 B.n670 10.6151
R895 B.n670 B.n669 10.6151
R896 B.n669 B.n30 10.6151
R897 B.n665 B.n30 10.6151
R898 B.n665 B.n664 10.6151
R899 B.n664 B.n663 10.6151
R900 B.n663 B.n32 10.6151
R901 B.n659 B.n32 10.6151
R902 B.n659 B.n658 10.6151
R903 B.n658 B.n657 10.6151
R904 B.n657 B.n34 10.6151
R905 B.n653 B.n34 10.6151
R906 B.n653 B.n652 10.6151
R907 B.n652 B.n651 10.6151
R908 B.n651 B.n36 10.6151
R909 B.n647 B.n36 10.6151
R910 B.n647 B.n646 10.6151
R911 B.n646 B.n645 10.6151
R912 B.n645 B.n38 10.6151
R913 B.n641 B.n38 10.6151
R914 B.n641 B.n640 10.6151
R915 B.n640 B.n639 10.6151
R916 B.n639 B.n40 10.6151
R917 B.n635 B.n40 10.6151
R918 B.n635 B.n634 10.6151
R919 B.n634 B.n633 10.6151
R920 B.n633 B.n42 10.6151
R921 B.n629 B.n42 10.6151
R922 B.n629 B.n628 10.6151
R923 B.n628 B.n627 10.6151
R924 B.n627 B.n44 10.6151
R925 B.n623 B.n44 10.6151
R926 B.n623 B.n622 10.6151
R927 B.n620 B.n48 10.6151
R928 B.n616 B.n48 10.6151
R929 B.n616 B.n615 10.6151
R930 B.n615 B.n614 10.6151
R931 B.n614 B.n50 10.6151
R932 B.n610 B.n50 10.6151
R933 B.n610 B.n609 10.6151
R934 B.n609 B.n608 10.6151
R935 B.n608 B.n52 10.6151
R936 B.n604 B.n603 10.6151
R937 B.n603 B.n602 10.6151
R938 B.n602 B.n57 10.6151
R939 B.n598 B.n57 10.6151
R940 B.n598 B.n597 10.6151
R941 B.n597 B.n596 10.6151
R942 B.n596 B.n59 10.6151
R943 B.n592 B.n59 10.6151
R944 B.n592 B.n591 10.6151
R945 B.n591 B.n590 10.6151
R946 B.n590 B.n61 10.6151
R947 B.n586 B.n61 10.6151
R948 B.n586 B.n585 10.6151
R949 B.n585 B.n584 10.6151
R950 B.n584 B.n63 10.6151
R951 B.n580 B.n63 10.6151
R952 B.n580 B.n579 10.6151
R953 B.n579 B.n578 10.6151
R954 B.n578 B.n65 10.6151
R955 B.n574 B.n65 10.6151
R956 B.n574 B.n573 10.6151
R957 B.n573 B.n572 10.6151
R958 B.n572 B.n67 10.6151
R959 B.n568 B.n67 10.6151
R960 B.n568 B.n567 10.6151
R961 B.n567 B.n566 10.6151
R962 B.n566 B.n69 10.6151
R963 B.n562 B.n69 10.6151
R964 B.n562 B.n561 10.6151
R965 B.n561 B.n560 10.6151
R966 B.n560 B.n71 10.6151
R967 B.n556 B.n71 10.6151
R968 B.n556 B.n555 10.6151
R969 B.n555 B.n554 10.6151
R970 B.n554 B.n73 10.6151
R971 B.n550 B.n73 10.6151
R972 B.n550 B.n549 10.6151
R973 B.n549 B.n548 10.6151
R974 B.n548 B.n75 10.6151
R975 B.n544 B.n75 10.6151
R976 B.n544 B.n543 10.6151
R977 B.n543 B.n542 10.6151
R978 B.n542 B.n77 10.6151
R979 B.n538 B.n77 10.6151
R980 B.n538 B.n537 10.6151
R981 B.n537 B.n536 10.6151
R982 B.n536 B.n79 10.6151
R983 B.n532 B.n79 10.6151
R984 B.n532 B.n531 10.6151
R985 B.n531 B.n530 10.6151
R986 B.n530 B.n81 10.6151
R987 B.n526 B.n81 10.6151
R988 B.n526 B.n525 10.6151
R989 B.n524 B.n83 10.6151
R990 B.n520 B.n83 10.6151
R991 B.n520 B.n519 10.6151
R992 B.n519 B.n518 10.6151
R993 B.n518 B.n85 10.6151
R994 B.n514 B.n85 10.6151
R995 B.n514 B.n513 10.6151
R996 B.n513 B.n512 10.6151
R997 B.n512 B.n87 10.6151
R998 B.n508 B.n87 10.6151
R999 B.n508 B.n507 10.6151
R1000 B.n507 B.n506 10.6151
R1001 B.n506 B.n89 10.6151
R1002 B.n502 B.n89 10.6151
R1003 B.n502 B.n501 10.6151
R1004 B.n501 B.n500 10.6151
R1005 B.n500 B.n91 10.6151
R1006 B.n496 B.n91 10.6151
R1007 B.n496 B.n495 10.6151
R1008 B.n495 B.n494 10.6151
R1009 B.n494 B.n93 10.6151
R1010 B.n490 B.n93 10.6151
R1011 B.n490 B.n489 10.6151
R1012 B.n489 B.n488 10.6151
R1013 B.n488 B.n95 10.6151
R1014 B.n484 B.n95 10.6151
R1015 B.n484 B.n483 10.6151
R1016 B.n483 B.n482 10.6151
R1017 B.n482 B.n97 10.6151
R1018 B.n478 B.n97 10.6151
R1019 B.n478 B.n477 10.6151
R1020 B.n477 B.n476 10.6151
R1021 B.n476 B.n99 10.6151
R1022 B.n472 B.n99 10.6151
R1023 B.n472 B.n471 10.6151
R1024 B.n471 B.n470 10.6151
R1025 B.n470 B.n101 10.6151
R1026 B.n466 B.n101 10.6151
R1027 B.n466 B.n465 10.6151
R1028 B.n465 B.n464 10.6151
R1029 B.n464 B.n103 10.6151
R1030 B.n460 B.n103 10.6151
R1031 B.n460 B.n459 10.6151
R1032 B.n459 B.n458 10.6151
R1033 B.n458 B.n105 10.6151
R1034 B.n454 B.n105 10.6151
R1035 B.n454 B.n453 10.6151
R1036 B.n453 B.n452 10.6151
R1037 B.n452 B.n107 10.6151
R1038 B.n448 B.n107 10.6151
R1039 B.n448 B.n447 10.6151
R1040 B.n447 B.n446 10.6151
R1041 B.n446 B.n109 10.6151
R1042 B.n442 B.n109 10.6151
R1043 B.n442 B.n441 10.6151
R1044 B.n441 B.n440 10.6151
R1045 B.n440 B.n111 10.6151
R1046 B.n436 B.n111 10.6151
R1047 B.n436 B.n435 10.6151
R1048 B.n435 B.n434 10.6151
R1049 B.n434 B.n113 10.6151
R1050 B.n430 B.n113 10.6151
R1051 B.n430 B.n429 10.6151
R1052 B.n429 B.n428 10.6151
R1053 B.n428 B.n115 10.6151
R1054 B.n424 B.n115 10.6151
R1055 B.n424 B.n423 10.6151
R1056 B.n193 B.n1 10.6151
R1057 B.n196 B.n193 10.6151
R1058 B.n197 B.n196 10.6151
R1059 B.n198 B.n197 10.6151
R1060 B.n198 B.n191 10.6151
R1061 B.n202 B.n191 10.6151
R1062 B.n203 B.n202 10.6151
R1063 B.n204 B.n203 10.6151
R1064 B.n204 B.n189 10.6151
R1065 B.n208 B.n189 10.6151
R1066 B.n209 B.n208 10.6151
R1067 B.n210 B.n209 10.6151
R1068 B.n210 B.n187 10.6151
R1069 B.n214 B.n187 10.6151
R1070 B.n215 B.n214 10.6151
R1071 B.n216 B.n215 10.6151
R1072 B.n216 B.n185 10.6151
R1073 B.n220 B.n185 10.6151
R1074 B.n221 B.n220 10.6151
R1075 B.n222 B.n221 10.6151
R1076 B.n222 B.n183 10.6151
R1077 B.n226 B.n183 10.6151
R1078 B.n227 B.n226 10.6151
R1079 B.n228 B.n227 10.6151
R1080 B.n228 B.n181 10.6151
R1081 B.n232 B.n181 10.6151
R1082 B.n233 B.n232 10.6151
R1083 B.n234 B.n233 10.6151
R1084 B.n234 B.n179 10.6151
R1085 B.n238 B.n179 10.6151
R1086 B.n239 B.n238 10.6151
R1087 B.n240 B.n239 10.6151
R1088 B.n244 B.n177 10.6151
R1089 B.n245 B.n244 10.6151
R1090 B.n246 B.n245 10.6151
R1091 B.n246 B.n175 10.6151
R1092 B.n250 B.n175 10.6151
R1093 B.n251 B.n250 10.6151
R1094 B.n252 B.n251 10.6151
R1095 B.n252 B.n173 10.6151
R1096 B.n256 B.n173 10.6151
R1097 B.n257 B.n256 10.6151
R1098 B.n258 B.n257 10.6151
R1099 B.n258 B.n171 10.6151
R1100 B.n262 B.n171 10.6151
R1101 B.n263 B.n262 10.6151
R1102 B.n264 B.n263 10.6151
R1103 B.n264 B.n169 10.6151
R1104 B.n268 B.n169 10.6151
R1105 B.n269 B.n268 10.6151
R1106 B.n270 B.n269 10.6151
R1107 B.n270 B.n167 10.6151
R1108 B.n274 B.n167 10.6151
R1109 B.n275 B.n274 10.6151
R1110 B.n276 B.n275 10.6151
R1111 B.n276 B.n165 10.6151
R1112 B.n280 B.n165 10.6151
R1113 B.n281 B.n280 10.6151
R1114 B.n282 B.n281 10.6151
R1115 B.n282 B.n163 10.6151
R1116 B.n286 B.n163 10.6151
R1117 B.n287 B.n286 10.6151
R1118 B.n288 B.n287 10.6151
R1119 B.n288 B.n161 10.6151
R1120 B.n292 B.n161 10.6151
R1121 B.n293 B.n292 10.6151
R1122 B.n294 B.n293 10.6151
R1123 B.n294 B.n159 10.6151
R1124 B.n298 B.n159 10.6151
R1125 B.n299 B.n298 10.6151
R1126 B.n300 B.n299 10.6151
R1127 B.n300 B.n157 10.6151
R1128 B.n304 B.n157 10.6151
R1129 B.n305 B.n304 10.6151
R1130 B.n306 B.n305 10.6151
R1131 B.n306 B.n155 10.6151
R1132 B.n310 B.n155 10.6151
R1133 B.n311 B.n310 10.6151
R1134 B.n312 B.n311 10.6151
R1135 B.n312 B.n153 10.6151
R1136 B.n316 B.n153 10.6151
R1137 B.n317 B.n316 10.6151
R1138 B.n318 B.n317 10.6151
R1139 B.n318 B.n151 10.6151
R1140 B.n322 B.n151 10.6151
R1141 B.n325 B.n324 10.6151
R1142 B.n325 B.n147 10.6151
R1143 B.n329 B.n147 10.6151
R1144 B.n330 B.n329 10.6151
R1145 B.n331 B.n330 10.6151
R1146 B.n331 B.n145 10.6151
R1147 B.n335 B.n145 10.6151
R1148 B.n336 B.n335 10.6151
R1149 B.n340 B.n336 10.6151
R1150 B.n344 B.n143 10.6151
R1151 B.n345 B.n344 10.6151
R1152 B.n346 B.n345 10.6151
R1153 B.n346 B.n141 10.6151
R1154 B.n350 B.n141 10.6151
R1155 B.n351 B.n350 10.6151
R1156 B.n352 B.n351 10.6151
R1157 B.n352 B.n139 10.6151
R1158 B.n356 B.n139 10.6151
R1159 B.n357 B.n356 10.6151
R1160 B.n358 B.n357 10.6151
R1161 B.n358 B.n137 10.6151
R1162 B.n362 B.n137 10.6151
R1163 B.n363 B.n362 10.6151
R1164 B.n364 B.n363 10.6151
R1165 B.n364 B.n135 10.6151
R1166 B.n368 B.n135 10.6151
R1167 B.n369 B.n368 10.6151
R1168 B.n370 B.n369 10.6151
R1169 B.n370 B.n133 10.6151
R1170 B.n374 B.n133 10.6151
R1171 B.n375 B.n374 10.6151
R1172 B.n376 B.n375 10.6151
R1173 B.n376 B.n131 10.6151
R1174 B.n380 B.n131 10.6151
R1175 B.n381 B.n380 10.6151
R1176 B.n382 B.n381 10.6151
R1177 B.n382 B.n129 10.6151
R1178 B.n386 B.n129 10.6151
R1179 B.n387 B.n386 10.6151
R1180 B.n388 B.n387 10.6151
R1181 B.n388 B.n127 10.6151
R1182 B.n392 B.n127 10.6151
R1183 B.n393 B.n392 10.6151
R1184 B.n394 B.n393 10.6151
R1185 B.n394 B.n125 10.6151
R1186 B.n398 B.n125 10.6151
R1187 B.n399 B.n398 10.6151
R1188 B.n400 B.n399 10.6151
R1189 B.n400 B.n123 10.6151
R1190 B.n404 B.n123 10.6151
R1191 B.n405 B.n404 10.6151
R1192 B.n406 B.n405 10.6151
R1193 B.n406 B.n121 10.6151
R1194 B.n410 B.n121 10.6151
R1195 B.n411 B.n410 10.6151
R1196 B.n412 B.n411 10.6151
R1197 B.n412 B.n119 10.6151
R1198 B.n416 B.n119 10.6151
R1199 B.n417 B.n416 10.6151
R1200 B.n418 B.n417 10.6151
R1201 B.n418 B.n117 10.6151
R1202 B.n422 B.n117 10.6151
R1203 B.n622 B.n621 9.36635
R1204 B.n604 B.n56 9.36635
R1205 B.n323 B.n322 9.36635
R1206 B.n339 B.n143 9.36635
R1207 B.n753 B.n0 8.11757
R1208 B.n753 B.n1 8.11757
R1209 B.n621 B.n620 1.24928
R1210 B.n56 B.n52 1.24928
R1211 B.n324 B.n323 1.24928
R1212 B.n340 B.n339 1.24928
R1213 VP.n6 VP.t3 243.796
R1214 VP.n17 VP.t2 213.123
R1215 VP.n24 VP.t1 213.123
R1216 VP.n31 VP.t0 213.123
R1217 VP.n14 VP.t4 213.123
R1218 VP.n7 VP.t5 213.123
R1219 VP.n9 VP.n8 161.3
R1220 VP.n10 VP.n5 161.3
R1221 VP.n12 VP.n11 161.3
R1222 VP.n13 VP.n4 161.3
R1223 VP.n30 VP.n0 161.3
R1224 VP.n29 VP.n28 161.3
R1225 VP.n27 VP.n1 161.3
R1226 VP.n26 VP.n25 161.3
R1227 VP.n23 VP.n2 161.3
R1228 VP.n22 VP.n21 161.3
R1229 VP.n20 VP.n3 161.3
R1230 VP.n19 VP.n18 161.3
R1231 VP.n17 VP.n16 89.7593
R1232 VP.n32 VP.n31 89.7593
R1233 VP.n15 VP.n14 89.7593
R1234 VP.n7 VP.n6 57.8394
R1235 VP.n22 VP.n3 56.0773
R1236 VP.n29 VP.n1 56.0773
R1237 VP.n12 VP.n5 56.0773
R1238 VP.n16 VP.n15 49.0451
R1239 VP.n18 VP.n3 25.0767
R1240 VP.n30 VP.n29 25.0767
R1241 VP.n13 VP.n12 25.0767
R1242 VP.n23 VP.n22 24.5923
R1243 VP.n25 VP.n1 24.5923
R1244 VP.n8 VP.n5 24.5923
R1245 VP.n18 VP.n17 21.1495
R1246 VP.n31 VP.n30 21.1495
R1247 VP.n14 VP.n13 21.1495
R1248 VP.n9 VP.n6 13.1274
R1249 VP.n24 VP.n23 12.2964
R1250 VP.n25 VP.n24 12.2964
R1251 VP.n8 VP.n7 12.2964
R1252 VP.n15 VP.n4 0.278335
R1253 VP.n19 VP.n16 0.278335
R1254 VP.n32 VP.n0 0.278335
R1255 VP.n10 VP.n9 0.189894
R1256 VP.n11 VP.n10 0.189894
R1257 VP.n11 VP.n4 0.189894
R1258 VP.n20 VP.n19 0.189894
R1259 VP.n21 VP.n20 0.189894
R1260 VP.n21 VP.n2 0.189894
R1261 VP.n26 VP.n2 0.189894
R1262 VP.n27 VP.n26 0.189894
R1263 VP.n28 VP.n27 0.189894
R1264 VP.n28 VP.n0 0.189894
R1265 VP VP.n32 0.153485
R1266 VDD1 VDD1.t2 71.4945
R1267 VDD1.n1 VDD1.t3 71.3807
R1268 VDD1.n1 VDD1.n0 68.4542
R1269 VDD1.n3 VDD1.n2 68.0398
R1270 VDD1.n3 VDD1.n1 45.4492
R1271 VDD1.n2 VDD1.t0 1.98736
R1272 VDD1.n2 VDD1.t1 1.98736
R1273 VDD1.n0 VDD1.t4 1.98736
R1274 VDD1.n0 VDD1.t5 1.98736
R1275 VDD1 VDD1.n3 0.412138
C0 B VN 1.063f
C1 VP VN 7.0044f
C2 VTAIL B 4.27919f
C3 VDD2 B 2.28536f
C4 VTAIL VP 8.184791f
C5 B w_n2714_n4240# 9.86246f
C6 VDD2 VP 0.395619f
C7 VP w_n2714_n4240# 5.39065f
C8 VDD1 B 2.22923f
C9 VDD1 VP 8.60523f
C10 VTAIL VN 8.17033f
C11 VDD2 VN 8.36416f
C12 w_n2714_n4240# VN 5.04186f
C13 VTAIL VDD2 9.63519f
C14 VTAIL w_n2714_n4240# 3.5529f
C15 VDD1 VN 0.1501f
C16 VDD2 w_n2714_n4240# 2.47859f
C17 VP B 1.64157f
C18 VTAIL VDD1 9.59177f
C19 VDD2 VDD1 1.14076f
C20 VDD1 w_n2714_n4240# 2.41746f
C21 VDD2 VSUBS 1.835455f
C22 VDD1 VSUBS 2.253084f
C23 VTAIL VSUBS 1.212625f
C24 VN VSUBS 5.38985f
C25 VP VSUBS 2.522218f
C26 B VSUBS 4.264958f
C27 w_n2714_n4240# VSUBS 0.140922p
C28 VDD1.t2 VSUBS 3.73029f
C29 VDD1.t3 VSUBS 3.7289f
C30 VDD1.t4 VSUBS 0.349402f
C31 VDD1.t5 VSUBS 0.349402f
C32 VDD1.n0 VSUBS 2.86433f
C33 VDD1.n1 VSUBS 3.84259f
C34 VDD1.t0 VSUBS 0.349402f
C35 VDD1.t1 VSUBS 0.349402f
C36 VDD1.n2 VSUBS 2.85981f
C37 VDD1.n3 VSUBS 3.45811f
C38 VP.n0 VSUBS 0.045884f
C39 VP.t0 VSUBS 2.89198f
C40 VP.n1 VSUBS 0.059175f
C41 VP.n2 VSUBS 0.034805f
C42 VP.t1 VSUBS 2.89198f
C43 VP.n3 VSUBS 0.04141f
C44 VP.n4 VSUBS 0.045884f
C45 VP.t4 VSUBS 2.89198f
C46 VP.n5 VSUBS 0.059175f
C47 VP.t3 VSUBS 3.03998f
C48 VP.n6 VSUBS 1.10671f
C49 VP.t5 VSUBS 2.89198f
C50 VP.n7 VSUBS 1.09428f
C51 VP.n8 VSUBS 0.048611f
C52 VP.n9 VSUBS 0.255903f
C53 VP.n10 VSUBS 0.034805f
C54 VP.n11 VSUBS 0.034805f
C55 VP.n12 VSUBS 0.04141f
C56 VP.n13 VSUBS 0.060685f
C57 VP.n14 VSUBS 1.11664f
C58 VP.n15 VSUBS 1.86436f
C59 VP.n16 VSUBS 1.88995f
C60 VP.t2 VSUBS 2.89198f
C61 VP.n17 VSUBS 1.11664f
C62 VP.n18 VSUBS 0.060685f
C63 VP.n19 VSUBS 0.045884f
C64 VP.n20 VSUBS 0.034805f
C65 VP.n21 VSUBS 0.034805f
C66 VP.n22 VSUBS 0.059175f
C67 VP.n23 VSUBS 0.048611f
C68 VP.n24 VSUBS 1.0159f
C69 VP.n25 VSUBS 0.048611f
C70 VP.n26 VSUBS 0.034805f
C71 VP.n27 VSUBS 0.034805f
C72 VP.n28 VSUBS 0.034805f
C73 VP.n29 VSUBS 0.04141f
C74 VP.n30 VSUBS 0.060685f
C75 VP.n31 VSUBS 1.11664f
C76 VP.n32 VSUBS 0.040205f
C77 B.n0 VSUBS 0.006991f
C78 B.n1 VSUBS 0.006991f
C79 B.n2 VSUBS 0.01034f
C80 B.n3 VSUBS 0.007924f
C81 B.n4 VSUBS 0.007924f
C82 B.n5 VSUBS 0.007924f
C83 B.n6 VSUBS 0.007924f
C84 B.n7 VSUBS 0.007924f
C85 B.n8 VSUBS 0.007924f
C86 B.n9 VSUBS 0.007924f
C87 B.n10 VSUBS 0.007924f
C88 B.n11 VSUBS 0.007924f
C89 B.n12 VSUBS 0.007924f
C90 B.n13 VSUBS 0.007924f
C91 B.n14 VSUBS 0.007924f
C92 B.n15 VSUBS 0.007924f
C93 B.n16 VSUBS 0.007924f
C94 B.n17 VSUBS 0.007924f
C95 B.n18 VSUBS 0.019985f
C96 B.n19 VSUBS 0.007924f
C97 B.n20 VSUBS 0.007924f
C98 B.n21 VSUBS 0.007924f
C99 B.n22 VSUBS 0.007924f
C100 B.n23 VSUBS 0.007924f
C101 B.n24 VSUBS 0.007924f
C102 B.n25 VSUBS 0.007924f
C103 B.n26 VSUBS 0.007924f
C104 B.n27 VSUBS 0.007924f
C105 B.n28 VSUBS 0.007924f
C106 B.n29 VSUBS 0.007924f
C107 B.n30 VSUBS 0.007924f
C108 B.n31 VSUBS 0.007924f
C109 B.n32 VSUBS 0.007924f
C110 B.n33 VSUBS 0.007924f
C111 B.n34 VSUBS 0.007924f
C112 B.n35 VSUBS 0.007924f
C113 B.n36 VSUBS 0.007924f
C114 B.n37 VSUBS 0.007924f
C115 B.n38 VSUBS 0.007924f
C116 B.n39 VSUBS 0.007924f
C117 B.n40 VSUBS 0.007924f
C118 B.n41 VSUBS 0.007924f
C119 B.n42 VSUBS 0.007924f
C120 B.n43 VSUBS 0.007924f
C121 B.n44 VSUBS 0.007924f
C122 B.n45 VSUBS 0.007924f
C123 B.t7 VSUBS 0.62078f
C124 B.t8 VSUBS 0.639673f
C125 B.t6 VSUBS 1.4906f
C126 B.n46 VSUBS 0.304256f
C127 B.n47 VSUBS 0.07807f
C128 B.n48 VSUBS 0.007924f
C129 B.n49 VSUBS 0.007924f
C130 B.n50 VSUBS 0.007924f
C131 B.n51 VSUBS 0.007924f
C132 B.n52 VSUBS 0.004428f
C133 B.n53 VSUBS 0.007924f
C134 B.t1 VSUBS 0.62076f
C135 B.t2 VSUBS 0.639656f
C136 B.t0 VSUBS 1.4906f
C137 B.n54 VSUBS 0.304273f
C138 B.n55 VSUBS 0.07809f
C139 B.n56 VSUBS 0.018358f
C140 B.n57 VSUBS 0.007924f
C141 B.n58 VSUBS 0.007924f
C142 B.n59 VSUBS 0.007924f
C143 B.n60 VSUBS 0.007924f
C144 B.n61 VSUBS 0.007924f
C145 B.n62 VSUBS 0.007924f
C146 B.n63 VSUBS 0.007924f
C147 B.n64 VSUBS 0.007924f
C148 B.n65 VSUBS 0.007924f
C149 B.n66 VSUBS 0.007924f
C150 B.n67 VSUBS 0.007924f
C151 B.n68 VSUBS 0.007924f
C152 B.n69 VSUBS 0.007924f
C153 B.n70 VSUBS 0.007924f
C154 B.n71 VSUBS 0.007924f
C155 B.n72 VSUBS 0.007924f
C156 B.n73 VSUBS 0.007924f
C157 B.n74 VSUBS 0.007924f
C158 B.n75 VSUBS 0.007924f
C159 B.n76 VSUBS 0.007924f
C160 B.n77 VSUBS 0.007924f
C161 B.n78 VSUBS 0.007924f
C162 B.n79 VSUBS 0.007924f
C163 B.n80 VSUBS 0.007924f
C164 B.n81 VSUBS 0.007924f
C165 B.n82 VSUBS 0.020798f
C166 B.n83 VSUBS 0.007924f
C167 B.n84 VSUBS 0.007924f
C168 B.n85 VSUBS 0.007924f
C169 B.n86 VSUBS 0.007924f
C170 B.n87 VSUBS 0.007924f
C171 B.n88 VSUBS 0.007924f
C172 B.n89 VSUBS 0.007924f
C173 B.n90 VSUBS 0.007924f
C174 B.n91 VSUBS 0.007924f
C175 B.n92 VSUBS 0.007924f
C176 B.n93 VSUBS 0.007924f
C177 B.n94 VSUBS 0.007924f
C178 B.n95 VSUBS 0.007924f
C179 B.n96 VSUBS 0.007924f
C180 B.n97 VSUBS 0.007924f
C181 B.n98 VSUBS 0.007924f
C182 B.n99 VSUBS 0.007924f
C183 B.n100 VSUBS 0.007924f
C184 B.n101 VSUBS 0.007924f
C185 B.n102 VSUBS 0.007924f
C186 B.n103 VSUBS 0.007924f
C187 B.n104 VSUBS 0.007924f
C188 B.n105 VSUBS 0.007924f
C189 B.n106 VSUBS 0.007924f
C190 B.n107 VSUBS 0.007924f
C191 B.n108 VSUBS 0.007924f
C192 B.n109 VSUBS 0.007924f
C193 B.n110 VSUBS 0.007924f
C194 B.n111 VSUBS 0.007924f
C195 B.n112 VSUBS 0.007924f
C196 B.n113 VSUBS 0.007924f
C197 B.n114 VSUBS 0.007924f
C198 B.n115 VSUBS 0.007924f
C199 B.n116 VSUBS 0.019985f
C200 B.n117 VSUBS 0.007924f
C201 B.n118 VSUBS 0.007924f
C202 B.n119 VSUBS 0.007924f
C203 B.n120 VSUBS 0.007924f
C204 B.n121 VSUBS 0.007924f
C205 B.n122 VSUBS 0.007924f
C206 B.n123 VSUBS 0.007924f
C207 B.n124 VSUBS 0.007924f
C208 B.n125 VSUBS 0.007924f
C209 B.n126 VSUBS 0.007924f
C210 B.n127 VSUBS 0.007924f
C211 B.n128 VSUBS 0.007924f
C212 B.n129 VSUBS 0.007924f
C213 B.n130 VSUBS 0.007924f
C214 B.n131 VSUBS 0.007924f
C215 B.n132 VSUBS 0.007924f
C216 B.n133 VSUBS 0.007924f
C217 B.n134 VSUBS 0.007924f
C218 B.n135 VSUBS 0.007924f
C219 B.n136 VSUBS 0.007924f
C220 B.n137 VSUBS 0.007924f
C221 B.n138 VSUBS 0.007924f
C222 B.n139 VSUBS 0.007924f
C223 B.n140 VSUBS 0.007924f
C224 B.n141 VSUBS 0.007924f
C225 B.n142 VSUBS 0.007924f
C226 B.n143 VSUBS 0.007458f
C227 B.n144 VSUBS 0.007924f
C228 B.n145 VSUBS 0.007924f
C229 B.n146 VSUBS 0.007924f
C230 B.n147 VSUBS 0.007924f
C231 B.n148 VSUBS 0.007924f
C232 B.t5 VSUBS 0.62078f
C233 B.t4 VSUBS 0.639673f
C234 B.t3 VSUBS 1.4906f
C235 B.n149 VSUBS 0.304256f
C236 B.n150 VSUBS 0.07807f
C237 B.n151 VSUBS 0.007924f
C238 B.n152 VSUBS 0.007924f
C239 B.n153 VSUBS 0.007924f
C240 B.n154 VSUBS 0.007924f
C241 B.n155 VSUBS 0.007924f
C242 B.n156 VSUBS 0.007924f
C243 B.n157 VSUBS 0.007924f
C244 B.n158 VSUBS 0.007924f
C245 B.n159 VSUBS 0.007924f
C246 B.n160 VSUBS 0.007924f
C247 B.n161 VSUBS 0.007924f
C248 B.n162 VSUBS 0.007924f
C249 B.n163 VSUBS 0.007924f
C250 B.n164 VSUBS 0.007924f
C251 B.n165 VSUBS 0.007924f
C252 B.n166 VSUBS 0.007924f
C253 B.n167 VSUBS 0.007924f
C254 B.n168 VSUBS 0.007924f
C255 B.n169 VSUBS 0.007924f
C256 B.n170 VSUBS 0.007924f
C257 B.n171 VSUBS 0.007924f
C258 B.n172 VSUBS 0.007924f
C259 B.n173 VSUBS 0.007924f
C260 B.n174 VSUBS 0.007924f
C261 B.n175 VSUBS 0.007924f
C262 B.n176 VSUBS 0.007924f
C263 B.n177 VSUBS 0.020798f
C264 B.n178 VSUBS 0.007924f
C265 B.n179 VSUBS 0.007924f
C266 B.n180 VSUBS 0.007924f
C267 B.n181 VSUBS 0.007924f
C268 B.n182 VSUBS 0.007924f
C269 B.n183 VSUBS 0.007924f
C270 B.n184 VSUBS 0.007924f
C271 B.n185 VSUBS 0.007924f
C272 B.n186 VSUBS 0.007924f
C273 B.n187 VSUBS 0.007924f
C274 B.n188 VSUBS 0.007924f
C275 B.n189 VSUBS 0.007924f
C276 B.n190 VSUBS 0.007924f
C277 B.n191 VSUBS 0.007924f
C278 B.n192 VSUBS 0.007924f
C279 B.n193 VSUBS 0.007924f
C280 B.n194 VSUBS 0.007924f
C281 B.n195 VSUBS 0.007924f
C282 B.n196 VSUBS 0.007924f
C283 B.n197 VSUBS 0.007924f
C284 B.n198 VSUBS 0.007924f
C285 B.n199 VSUBS 0.007924f
C286 B.n200 VSUBS 0.007924f
C287 B.n201 VSUBS 0.007924f
C288 B.n202 VSUBS 0.007924f
C289 B.n203 VSUBS 0.007924f
C290 B.n204 VSUBS 0.007924f
C291 B.n205 VSUBS 0.007924f
C292 B.n206 VSUBS 0.007924f
C293 B.n207 VSUBS 0.007924f
C294 B.n208 VSUBS 0.007924f
C295 B.n209 VSUBS 0.007924f
C296 B.n210 VSUBS 0.007924f
C297 B.n211 VSUBS 0.007924f
C298 B.n212 VSUBS 0.007924f
C299 B.n213 VSUBS 0.007924f
C300 B.n214 VSUBS 0.007924f
C301 B.n215 VSUBS 0.007924f
C302 B.n216 VSUBS 0.007924f
C303 B.n217 VSUBS 0.007924f
C304 B.n218 VSUBS 0.007924f
C305 B.n219 VSUBS 0.007924f
C306 B.n220 VSUBS 0.007924f
C307 B.n221 VSUBS 0.007924f
C308 B.n222 VSUBS 0.007924f
C309 B.n223 VSUBS 0.007924f
C310 B.n224 VSUBS 0.007924f
C311 B.n225 VSUBS 0.007924f
C312 B.n226 VSUBS 0.007924f
C313 B.n227 VSUBS 0.007924f
C314 B.n228 VSUBS 0.007924f
C315 B.n229 VSUBS 0.007924f
C316 B.n230 VSUBS 0.007924f
C317 B.n231 VSUBS 0.007924f
C318 B.n232 VSUBS 0.007924f
C319 B.n233 VSUBS 0.007924f
C320 B.n234 VSUBS 0.007924f
C321 B.n235 VSUBS 0.007924f
C322 B.n236 VSUBS 0.007924f
C323 B.n237 VSUBS 0.007924f
C324 B.n238 VSUBS 0.007924f
C325 B.n239 VSUBS 0.007924f
C326 B.n240 VSUBS 0.019985f
C327 B.n241 VSUBS 0.019985f
C328 B.n242 VSUBS 0.020798f
C329 B.n243 VSUBS 0.007924f
C330 B.n244 VSUBS 0.007924f
C331 B.n245 VSUBS 0.007924f
C332 B.n246 VSUBS 0.007924f
C333 B.n247 VSUBS 0.007924f
C334 B.n248 VSUBS 0.007924f
C335 B.n249 VSUBS 0.007924f
C336 B.n250 VSUBS 0.007924f
C337 B.n251 VSUBS 0.007924f
C338 B.n252 VSUBS 0.007924f
C339 B.n253 VSUBS 0.007924f
C340 B.n254 VSUBS 0.007924f
C341 B.n255 VSUBS 0.007924f
C342 B.n256 VSUBS 0.007924f
C343 B.n257 VSUBS 0.007924f
C344 B.n258 VSUBS 0.007924f
C345 B.n259 VSUBS 0.007924f
C346 B.n260 VSUBS 0.007924f
C347 B.n261 VSUBS 0.007924f
C348 B.n262 VSUBS 0.007924f
C349 B.n263 VSUBS 0.007924f
C350 B.n264 VSUBS 0.007924f
C351 B.n265 VSUBS 0.007924f
C352 B.n266 VSUBS 0.007924f
C353 B.n267 VSUBS 0.007924f
C354 B.n268 VSUBS 0.007924f
C355 B.n269 VSUBS 0.007924f
C356 B.n270 VSUBS 0.007924f
C357 B.n271 VSUBS 0.007924f
C358 B.n272 VSUBS 0.007924f
C359 B.n273 VSUBS 0.007924f
C360 B.n274 VSUBS 0.007924f
C361 B.n275 VSUBS 0.007924f
C362 B.n276 VSUBS 0.007924f
C363 B.n277 VSUBS 0.007924f
C364 B.n278 VSUBS 0.007924f
C365 B.n279 VSUBS 0.007924f
C366 B.n280 VSUBS 0.007924f
C367 B.n281 VSUBS 0.007924f
C368 B.n282 VSUBS 0.007924f
C369 B.n283 VSUBS 0.007924f
C370 B.n284 VSUBS 0.007924f
C371 B.n285 VSUBS 0.007924f
C372 B.n286 VSUBS 0.007924f
C373 B.n287 VSUBS 0.007924f
C374 B.n288 VSUBS 0.007924f
C375 B.n289 VSUBS 0.007924f
C376 B.n290 VSUBS 0.007924f
C377 B.n291 VSUBS 0.007924f
C378 B.n292 VSUBS 0.007924f
C379 B.n293 VSUBS 0.007924f
C380 B.n294 VSUBS 0.007924f
C381 B.n295 VSUBS 0.007924f
C382 B.n296 VSUBS 0.007924f
C383 B.n297 VSUBS 0.007924f
C384 B.n298 VSUBS 0.007924f
C385 B.n299 VSUBS 0.007924f
C386 B.n300 VSUBS 0.007924f
C387 B.n301 VSUBS 0.007924f
C388 B.n302 VSUBS 0.007924f
C389 B.n303 VSUBS 0.007924f
C390 B.n304 VSUBS 0.007924f
C391 B.n305 VSUBS 0.007924f
C392 B.n306 VSUBS 0.007924f
C393 B.n307 VSUBS 0.007924f
C394 B.n308 VSUBS 0.007924f
C395 B.n309 VSUBS 0.007924f
C396 B.n310 VSUBS 0.007924f
C397 B.n311 VSUBS 0.007924f
C398 B.n312 VSUBS 0.007924f
C399 B.n313 VSUBS 0.007924f
C400 B.n314 VSUBS 0.007924f
C401 B.n315 VSUBS 0.007924f
C402 B.n316 VSUBS 0.007924f
C403 B.n317 VSUBS 0.007924f
C404 B.n318 VSUBS 0.007924f
C405 B.n319 VSUBS 0.007924f
C406 B.n320 VSUBS 0.007924f
C407 B.n321 VSUBS 0.007924f
C408 B.n322 VSUBS 0.007458f
C409 B.n323 VSUBS 0.018358f
C410 B.n324 VSUBS 0.004428f
C411 B.n325 VSUBS 0.007924f
C412 B.n326 VSUBS 0.007924f
C413 B.n327 VSUBS 0.007924f
C414 B.n328 VSUBS 0.007924f
C415 B.n329 VSUBS 0.007924f
C416 B.n330 VSUBS 0.007924f
C417 B.n331 VSUBS 0.007924f
C418 B.n332 VSUBS 0.007924f
C419 B.n333 VSUBS 0.007924f
C420 B.n334 VSUBS 0.007924f
C421 B.n335 VSUBS 0.007924f
C422 B.n336 VSUBS 0.007924f
C423 B.t11 VSUBS 0.62076f
C424 B.t10 VSUBS 0.639656f
C425 B.t9 VSUBS 1.4906f
C426 B.n337 VSUBS 0.304273f
C427 B.n338 VSUBS 0.07809f
C428 B.n339 VSUBS 0.018358f
C429 B.n340 VSUBS 0.004428f
C430 B.n341 VSUBS 0.007924f
C431 B.n342 VSUBS 0.007924f
C432 B.n343 VSUBS 0.007924f
C433 B.n344 VSUBS 0.007924f
C434 B.n345 VSUBS 0.007924f
C435 B.n346 VSUBS 0.007924f
C436 B.n347 VSUBS 0.007924f
C437 B.n348 VSUBS 0.007924f
C438 B.n349 VSUBS 0.007924f
C439 B.n350 VSUBS 0.007924f
C440 B.n351 VSUBS 0.007924f
C441 B.n352 VSUBS 0.007924f
C442 B.n353 VSUBS 0.007924f
C443 B.n354 VSUBS 0.007924f
C444 B.n355 VSUBS 0.007924f
C445 B.n356 VSUBS 0.007924f
C446 B.n357 VSUBS 0.007924f
C447 B.n358 VSUBS 0.007924f
C448 B.n359 VSUBS 0.007924f
C449 B.n360 VSUBS 0.007924f
C450 B.n361 VSUBS 0.007924f
C451 B.n362 VSUBS 0.007924f
C452 B.n363 VSUBS 0.007924f
C453 B.n364 VSUBS 0.007924f
C454 B.n365 VSUBS 0.007924f
C455 B.n366 VSUBS 0.007924f
C456 B.n367 VSUBS 0.007924f
C457 B.n368 VSUBS 0.007924f
C458 B.n369 VSUBS 0.007924f
C459 B.n370 VSUBS 0.007924f
C460 B.n371 VSUBS 0.007924f
C461 B.n372 VSUBS 0.007924f
C462 B.n373 VSUBS 0.007924f
C463 B.n374 VSUBS 0.007924f
C464 B.n375 VSUBS 0.007924f
C465 B.n376 VSUBS 0.007924f
C466 B.n377 VSUBS 0.007924f
C467 B.n378 VSUBS 0.007924f
C468 B.n379 VSUBS 0.007924f
C469 B.n380 VSUBS 0.007924f
C470 B.n381 VSUBS 0.007924f
C471 B.n382 VSUBS 0.007924f
C472 B.n383 VSUBS 0.007924f
C473 B.n384 VSUBS 0.007924f
C474 B.n385 VSUBS 0.007924f
C475 B.n386 VSUBS 0.007924f
C476 B.n387 VSUBS 0.007924f
C477 B.n388 VSUBS 0.007924f
C478 B.n389 VSUBS 0.007924f
C479 B.n390 VSUBS 0.007924f
C480 B.n391 VSUBS 0.007924f
C481 B.n392 VSUBS 0.007924f
C482 B.n393 VSUBS 0.007924f
C483 B.n394 VSUBS 0.007924f
C484 B.n395 VSUBS 0.007924f
C485 B.n396 VSUBS 0.007924f
C486 B.n397 VSUBS 0.007924f
C487 B.n398 VSUBS 0.007924f
C488 B.n399 VSUBS 0.007924f
C489 B.n400 VSUBS 0.007924f
C490 B.n401 VSUBS 0.007924f
C491 B.n402 VSUBS 0.007924f
C492 B.n403 VSUBS 0.007924f
C493 B.n404 VSUBS 0.007924f
C494 B.n405 VSUBS 0.007924f
C495 B.n406 VSUBS 0.007924f
C496 B.n407 VSUBS 0.007924f
C497 B.n408 VSUBS 0.007924f
C498 B.n409 VSUBS 0.007924f
C499 B.n410 VSUBS 0.007924f
C500 B.n411 VSUBS 0.007924f
C501 B.n412 VSUBS 0.007924f
C502 B.n413 VSUBS 0.007924f
C503 B.n414 VSUBS 0.007924f
C504 B.n415 VSUBS 0.007924f
C505 B.n416 VSUBS 0.007924f
C506 B.n417 VSUBS 0.007924f
C507 B.n418 VSUBS 0.007924f
C508 B.n419 VSUBS 0.007924f
C509 B.n420 VSUBS 0.007924f
C510 B.n421 VSUBS 0.020798f
C511 B.n422 VSUBS 0.019985f
C512 B.n423 VSUBS 0.020798f
C513 B.n424 VSUBS 0.007924f
C514 B.n425 VSUBS 0.007924f
C515 B.n426 VSUBS 0.007924f
C516 B.n427 VSUBS 0.007924f
C517 B.n428 VSUBS 0.007924f
C518 B.n429 VSUBS 0.007924f
C519 B.n430 VSUBS 0.007924f
C520 B.n431 VSUBS 0.007924f
C521 B.n432 VSUBS 0.007924f
C522 B.n433 VSUBS 0.007924f
C523 B.n434 VSUBS 0.007924f
C524 B.n435 VSUBS 0.007924f
C525 B.n436 VSUBS 0.007924f
C526 B.n437 VSUBS 0.007924f
C527 B.n438 VSUBS 0.007924f
C528 B.n439 VSUBS 0.007924f
C529 B.n440 VSUBS 0.007924f
C530 B.n441 VSUBS 0.007924f
C531 B.n442 VSUBS 0.007924f
C532 B.n443 VSUBS 0.007924f
C533 B.n444 VSUBS 0.007924f
C534 B.n445 VSUBS 0.007924f
C535 B.n446 VSUBS 0.007924f
C536 B.n447 VSUBS 0.007924f
C537 B.n448 VSUBS 0.007924f
C538 B.n449 VSUBS 0.007924f
C539 B.n450 VSUBS 0.007924f
C540 B.n451 VSUBS 0.007924f
C541 B.n452 VSUBS 0.007924f
C542 B.n453 VSUBS 0.007924f
C543 B.n454 VSUBS 0.007924f
C544 B.n455 VSUBS 0.007924f
C545 B.n456 VSUBS 0.007924f
C546 B.n457 VSUBS 0.007924f
C547 B.n458 VSUBS 0.007924f
C548 B.n459 VSUBS 0.007924f
C549 B.n460 VSUBS 0.007924f
C550 B.n461 VSUBS 0.007924f
C551 B.n462 VSUBS 0.007924f
C552 B.n463 VSUBS 0.007924f
C553 B.n464 VSUBS 0.007924f
C554 B.n465 VSUBS 0.007924f
C555 B.n466 VSUBS 0.007924f
C556 B.n467 VSUBS 0.007924f
C557 B.n468 VSUBS 0.007924f
C558 B.n469 VSUBS 0.007924f
C559 B.n470 VSUBS 0.007924f
C560 B.n471 VSUBS 0.007924f
C561 B.n472 VSUBS 0.007924f
C562 B.n473 VSUBS 0.007924f
C563 B.n474 VSUBS 0.007924f
C564 B.n475 VSUBS 0.007924f
C565 B.n476 VSUBS 0.007924f
C566 B.n477 VSUBS 0.007924f
C567 B.n478 VSUBS 0.007924f
C568 B.n479 VSUBS 0.007924f
C569 B.n480 VSUBS 0.007924f
C570 B.n481 VSUBS 0.007924f
C571 B.n482 VSUBS 0.007924f
C572 B.n483 VSUBS 0.007924f
C573 B.n484 VSUBS 0.007924f
C574 B.n485 VSUBS 0.007924f
C575 B.n486 VSUBS 0.007924f
C576 B.n487 VSUBS 0.007924f
C577 B.n488 VSUBS 0.007924f
C578 B.n489 VSUBS 0.007924f
C579 B.n490 VSUBS 0.007924f
C580 B.n491 VSUBS 0.007924f
C581 B.n492 VSUBS 0.007924f
C582 B.n493 VSUBS 0.007924f
C583 B.n494 VSUBS 0.007924f
C584 B.n495 VSUBS 0.007924f
C585 B.n496 VSUBS 0.007924f
C586 B.n497 VSUBS 0.007924f
C587 B.n498 VSUBS 0.007924f
C588 B.n499 VSUBS 0.007924f
C589 B.n500 VSUBS 0.007924f
C590 B.n501 VSUBS 0.007924f
C591 B.n502 VSUBS 0.007924f
C592 B.n503 VSUBS 0.007924f
C593 B.n504 VSUBS 0.007924f
C594 B.n505 VSUBS 0.007924f
C595 B.n506 VSUBS 0.007924f
C596 B.n507 VSUBS 0.007924f
C597 B.n508 VSUBS 0.007924f
C598 B.n509 VSUBS 0.007924f
C599 B.n510 VSUBS 0.007924f
C600 B.n511 VSUBS 0.007924f
C601 B.n512 VSUBS 0.007924f
C602 B.n513 VSUBS 0.007924f
C603 B.n514 VSUBS 0.007924f
C604 B.n515 VSUBS 0.007924f
C605 B.n516 VSUBS 0.007924f
C606 B.n517 VSUBS 0.007924f
C607 B.n518 VSUBS 0.007924f
C608 B.n519 VSUBS 0.007924f
C609 B.n520 VSUBS 0.007924f
C610 B.n521 VSUBS 0.007924f
C611 B.n522 VSUBS 0.007924f
C612 B.n523 VSUBS 0.019985f
C613 B.n524 VSUBS 0.019985f
C614 B.n525 VSUBS 0.020798f
C615 B.n526 VSUBS 0.007924f
C616 B.n527 VSUBS 0.007924f
C617 B.n528 VSUBS 0.007924f
C618 B.n529 VSUBS 0.007924f
C619 B.n530 VSUBS 0.007924f
C620 B.n531 VSUBS 0.007924f
C621 B.n532 VSUBS 0.007924f
C622 B.n533 VSUBS 0.007924f
C623 B.n534 VSUBS 0.007924f
C624 B.n535 VSUBS 0.007924f
C625 B.n536 VSUBS 0.007924f
C626 B.n537 VSUBS 0.007924f
C627 B.n538 VSUBS 0.007924f
C628 B.n539 VSUBS 0.007924f
C629 B.n540 VSUBS 0.007924f
C630 B.n541 VSUBS 0.007924f
C631 B.n542 VSUBS 0.007924f
C632 B.n543 VSUBS 0.007924f
C633 B.n544 VSUBS 0.007924f
C634 B.n545 VSUBS 0.007924f
C635 B.n546 VSUBS 0.007924f
C636 B.n547 VSUBS 0.007924f
C637 B.n548 VSUBS 0.007924f
C638 B.n549 VSUBS 0.007924f
C639 B.n550 VSUBS 0.007924f
C640 B.n551 VSUBS 0.007924f
C641 B.n552 VSUBS 0.007924f
C642 B.n553 VSUBS 0.007924f
C643 B.n554 VSUBS 0.007924f
C644 B.n555 VSUBS 0.007924f
C645 B.n556 VSUBS 0.007924f
C646 B.n557 VSUBS 0.007924f
C647 B.n558 VSUBS 0.007924f
C648 B.n559 VSUBS 0.007924f
C649 B.n560 VSUBS 0.007924f
C650 B.n561 VSUBS 0.007924f
C651 B.n562 VSUBS 0.007924f
C652 B.n563 VSUBS 0.007924f
C653 B.n564 VSUBS 0.007924f
C654 B.n565 VSUBS 0.007924f
C655 B.n566 VSUBS 0.007924f
C656 B.n567 VSUBS 0.007924f
C657 B.n568 VSUBS 0.007924f
C658 B.n569 VSUBS 0.007924f
C659 B.n570 VSUBS 0.007924f
C660 B.n571 VSUBS 0.007924f
C661 B.n572 VSUBS 0.007924f
C662 B.n573 VSUBS 0.007924f
C663 B.n574 VSUBS 0.007924f
C664 B.n575 VSUBS 0.007924f
C665 B.n576 VSUBS 0.007924f
C666 B.n577 VSUBS 0.007924f
C667 B.n578 VSUBS 0.007924f
C668 B.n579 VSUBS 0.007924f
C669 B.n580 VSUBS 0.007924f
C670 B.n581 VSUBS 0.007924f
C671 B.n582 VSUBS 0.007924f
C672 B.n583 VSUBS 0.007924f
C673 B.n584 VSUBS 0.007924f
C674 B.n585 VSUBS 0.007924f
C675 B.n586 VSUBS 0.007924f
C676 B.n587 VSUBS 0.007924f
C677 B.n588 VSUBS 0.007924f
C678 B.n589 VSUBS 0.007924f
C679 B.n590 VSUBS 0.007924f
C680 B.n591 VSUBS 0.007924f
C681 B.n592 VSUBS 0.007924f
C682 B.n593 VSUBS 0.007924f
C683 B.n594 VSUBS 0.007924f
C684 B.n595 VSUBS 0.007924f
C685 B.n596 VSUBS 0.007924f
C686 B.n597 VSUBS 0.007924f
C687 B.n598 VSUBS 0.007924f
C688 B.n599 VSUBS 0.007924f
C689 B.n600 VSUBS 0.007924f
C690 B.n601 VSUBS 0.007924f
C691 B.n602 VSUBS 0.007924f
C692 B.n603 VSUBS 0.007924f
C693 B.n604 VSUBS 0.007458f
C694 B.n605 VSUBS 0.007924f
C695 B.n606 VSUBS 0.007924f
C696 B.n607 VSUBS 0.007924f
C697 B.n608 VSUBS 0.007924f
C698 B.n609 VSUBS 0.007924f
C699 B.n610 VSUBS 0.007924f
C700 B.n611 VSUBS 0.007924f
C701 B.n612 VSUBS 0.007924f
C702 B.n613 VSUBS 0.007924f
C703 B.n614 VSUBS 0.007924f
C704 B.n615 VSUBS 0.007924f
C705 B.n616 VSUBS 0.007924f
C706 B.n617 VSUBS 0.007924f
C707 B.n618 VSUBS 0.007924f
C708 B.n619 VSUBS 0.007924f
C709 B.n620 VSUBS 0.004428f
C710 B.n621 VSUBS 0.018358f
C711 B.n622 VSUBS 0.007458f
C712 B.n623 VSUBS 0.007924f
C713 B.n624 VSUBS 0.007924f
C714 B.n625 VSUBS 0.007924f
C715 B.n626 VSUBS 0.007924f
C716 B.n627 VSUBS 0.007924f
C717 B.n628 VSUBS 0.007924f
C718 B.n629 VSUBS 0.007924f
C719 B.n630 VSUBS 0.007924f
C720 B.n631 VSUBS 0.007924f
C721 B.n632 VSUBS 0.007924f
C722 B.n633 VSUBS 0.007924f
C723 B.n634 VSUBS 0.007924f
C724 B.n635 VSUBS 0.007924f
C725 B.n636 VSUBS 0.007924f
C726 B.n637 VSUBS 0.007924f
C727 B.n638 VSUBS 0.007924f
C728 B.n639 VSUBS 0.007924f
C729 B.n640 VSUBS 0.007924f
C730 B.n641 VSUBS 0.007924f
C731 B.n642 VSUBS 0.007924f
C732 B.n643 VSUBS 0.007924f
C733 B.n644 VSUBS 0.007924f
C734 B.n645 VSUBS 0.007924f
C735 B.n646 VSUBS 0.007924f
C736 B.n647 VSUBS 0.007924f
C737 B.n648 VSUBS 0.007924f
C738 B.n649 VSUBS 0.007924f
C739 B.n650 VSUBS 0.007924f
C740 B.n651 VSUBS 0.007924f
C741 B.n652 VSUBS 0.007924f
C742 B.n653 VSUBS 0.007924f
C743 B.n654 VSUBS 0.007924f
C744 B.n655 VSUBS 0.007924f
C745 B.n656 VSUBS 0.007924f
C746 B.n657 VSUBS 0.007924f
C747 B.n658 VSUBS 0.007924f
C748 B.n659 VSUBS 0.007924f
C749 B.n660 VSUBS 0.007924f
C750 B.n661 VSUBS 0.007924f
C751 B.n662 VSUBS 0.007924f
C752 B.n663 VSUBS 0.007924f
C753 B.n664 VSUBS 0.007924f
C754 B.n665 VSUBS 0.007924f
C755 B.n666 VSUBS 0.007924f
C756 B.n667 VSUBS 0.007924f
C757 B.n668 VSUBS 0.007924f
C758 B.n669 VSUBS 0.007924f
C759 B.n670 VSUBS 0.007924f
C760 B.n671 VSUBS 0.007924f
C761 B.n672 VSUBS 0.007924f
C762 B.n673 VSUBS 0.007924f
C763 B.n674 VSUBS 0.007924f
C764 B.n675 VSUBS 0.007924f
C765 B.n676 VSUBS 0.007924f
C766 B.n677 VSUBS 0.007924f
C767 B.n678 VSUBS 0.007924f
C768 B.n679 VSUBS 0.007924f
C769 B.n680 VSUBS 0.007924f
C770 B.n681 VSUBS 0.007924f
C771 B.n682 VSUBS 0.007924f
C772 B.n683 VSUBS 0.007924f
C773 B.n684 VSUBS 0.007924f
C774 B.n685 VSUBS 0.007924f
C775 B.n686 VSUBS 0.007924f
C776 B.n687 VSUBS 0.007924f
C777 B.n688 VSUBS 0.007924f
C778 B.n689 VSUBS 0.007924f
C779 B.n690 VSUBS 0.007924f
C780 B.n691 VSUBS 0.007924f
C781 B.n692 VSUBS 0.007924f
C782 B.n693 VSUBS 0.007924f
C783 B.n694 VSUBS 0.007924f
C784 B.n695 VSUBS 0.007924f
C785 B.n696 VSUBS 0.007924f
C786 B.n697 VSUBS 0.007924f
C787 B.n698 VSUBS 0.007924f
C788 B.n699 VSUBS 0.007924f
C789 B.n700 VSUBS 0.007924f
C790 B.n701 VSUBS 0.020798f
C791 B.n702 VSUBS 0.020798f
C792 B.n703 VSUBS 0.019985f
C793 B.n704 VSUBS 0.007924f
C794 B.n705 VSUBS 0.007924f
C795 B.n706 VSUBS 0.007924f
C796 B.n707 VSUBS 0.007924f
C797 B.n708 VSUBS 0.007924f
C798 B.n709 VSUBS 0.007924f
C799 B.n710 VSUBS 0.007924f
C800 B.n711 VSUBS 0.007924f
C801 B.n712 VSUBS 0.007924f
C802 B.n713 VSUBS 0.007924f
C803 B.n714 VSUBS 0.007924f
C804 B.n715 VSUBS 0.007924f
C805 B.n716 VSUBS 0.007924f
C806 B.n717 VSUBS 0.007924f
C807 B.n718 VSUBS 0.007924f
C808 B.n719 VSUBS 0.007924f
C809 B.n720 VSUBS 0.007924f
C810 B.n721 VSUBS 0.007924f
C811 B.n722 VSUBS 0.007924f
C812 B.n723 VSUBS 0.007924f
C813 B.n724 VSUBS 0.007924f
C814 B.n725 VSUBS 0.007924f
C815 B.n726 VSUBS 0.007924f
C816 B.n727 VSUBS 0.007924f
C817 B.n728 VSUBS 0.007924f
C818 B.n729 VSUBS 0.007924f
C819 B.n730 VSUBS 0.007924f
C820 B.n731 VSUBS 0.007924f
C821 B.n732 VSUBS 0.007924f
C822 B.n733 VSUBS 0.007924f
C823 B.n734 VSUBS 0.007924f
C824 B.n735 VSUBS 0.007924f
C825 B.n736 VSUBS 0.007924f
C826 B.n737 VSUBS 0.007924f
C827 B.n738 VSUBS 0.007924f
C828 B.n739 VSUBS 0.007924f
C829 B.n740 VSUBS 0.007924f
C830 B.n741 VSUBS 0.007924f
C831 B.n742 VSUBS 0.007924f
C832 B.n743 VSUBS 0.007924f
C833 B.n744 VSUBS 0.007924f
C834 B.n745 VSUBS 0.007924f
C835 B.n746 VSUBS 0.007924f
C836 B.n747 VSUBS 0.007924f
C837 B.n748 VSUBS 0.007924f
C838 B.n749 VSUBS 0.007924f
C839 B.n750 VSUBS 0.007924f
C840 B.n751 VSUBS 0.01034f
C841 B.n752 VSUBS 0.011015f
C842 B.n753 VSUBS 0.021904f
C843 VDD2.t4 VSUBS 3.7453f
C844 VDD2.t3 VSUBS 0.350939f
C845 VDD2.t5 VSUBS 0.350939f
C846 VDD2.n0 VSUBS 2.87692f
C847 VDD2.n1 VSUBS 3.74292f
C848 VDD2.t0 VSUBS 3.7308f
C849 VDD2.n2 VSUBS 3.51629f
C850 VDD2.t1 VSUBS 0.350939f
C851 VDD2.t2 VSUBS 0.350939f
C852 VDD2.n3 VSUBS 2.87687f
C853 VTAIL.t9 VSUBS 0.356586f
C854 VTAIL.t8 VSUBS 0.356586f
C855 VTAIL.n0 VSUBS 2.74348f
C856 VTAIL.n1 VSUBS 0.85438f
C857 VTAIL.t1 VSUBS 3.59088f
C858 VTAIL.n2 VSUBS 1.09959f
C859 VTAIL.t0 VSUBS 0.356586f
C860 VTAIL.t3 VSUBS 0.356586f
C861 VTAIL.n3 VSUBS 2.74348f
C862 VTAIL.n4 VSUBS 2.81138f
C863 VTAIL.t11 VSUBS 0.356586f
C864 VTAIL.t10 VSUBS 0.356586f
C865 VTAIL.n5 VSUBS 2.74349f
C866 VTAIL.n6 VSUBS 2.81138f
C867 VTAIL.t7 VSUBS 3.59088f
C868 VTAIL.n7 VSUBS 1.09959f
C869 VTAIL.t2 VSUBS 0.356586f
C870 VTAIL.t5 VSUBS 0.356586f
C871 VTAIL.n8 VSUBS 2.74349f
C872 VTAIL.n9 VSUBS 0.974471f
C873 VTAIL.t4 VSUBS 3.59088f
C874 VTAIL.n10 VSUBS 2.76948f
C875 VTAIL.t6 VSUBS 3.59088f
C876 VTAIL.n11 VSUBS 2.72255f
C877 VN.n0 VSUBS 0.044866f
C878 VN.t0 VSUBS 2.82782f
C879 VN.n1 VSUBS 0.057863f
C880 VN.t1 VSUBS 2.97253f
C881 VN.n2 VSUBS 1.08216f
C882 VN.t2 VSUBS 2.82782f
C883 VN.n3 VSUBS 1.07001f
C884 VN.n4 VSUBS 0.047532f
C885 VN.n5 VSUBS 0.250226f
C886 VN.n6 VSUBS 0.034033f
C887 VN.n7 VSUBS 0.034033f
C888 VN.n8 VSUBS 0.040491f
C889 VN.n9 VSUBS 0.059338f
C890 VN.n10 VSUBS 1.09187f
C891 VN.n11 VSUBS 0.039313f
C892 VN.n12 VSUBS 0.044866f
C893 VN.t5 VSUBS 2.82782f
C894 VN.n13 VSUBS 0.057863f
C895 VN.t3 VSUBS 2.97253f
C896 VN.n14 VSUBS 1.08216f
C897 VN.t4 VSUBS 2.82782f
C898 VN.n15 VSUBS 1.07001f
C899 VN.n16 VSUBS 0.047532f
C900 VN.n17 VSUBS 0.250226f
C901 VN.n18 VSUBS 0.034033f
C902 VN.n19 VSUBS 0.034033f
C903 VN.n20 VSUBS 0.040491f
C904 VN.n21 VSUBS 0.059338f
C905 VN.n22 VSUBS 1.09187f
C906 VN.n23 VSUBS 1.84134f
.ends

