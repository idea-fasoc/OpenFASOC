* NGSPICE file created from diff_pair_sample_1324.ext - technology: sky130A

.subckt diff_pair_sample_1324 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0 ps=0 w=3.51 l=3.77
X1 B.t8 B.t6 B.t7 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0 ps=0 w=3.51 l=3.77
X2 VDD2.t7 VN.t0 VTAIL.t13 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=1.3689 ps=7.8 w=3.51 l=3.77
X3 VTAIL.t4 VP.t0 VDD1.t7 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X4 VDD2.t6 VN.t1 VTAIL.t14 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=1.3689 ps=7.8 w=3.51 l=3.77
X5 VTAIL.t11 VN.t2 VDD2.t5 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X6 VDD1.t6 VP.t1 VTAIL.t7 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=1.3689 ps=7.8 w=3.51 l=3.77
X7 B.t5 B.t3 B.t4 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0 ps=0 w=3.51 l=3.77
X8 VTAIL.t9 VN.t3 VDD2.t4 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X9 VDD1.t5 VP.t2 VTAIL.t2 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=1.3689 ps=7.8 w=3.51 l=3.77
X10 VTAIL.t3 VP.t3 VDD1.t4 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0.57915 ps=3.84 w=3.51 l=3.77
X11 VDD2.t3 VN.t4 VTAIL.t12 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X12 VTAIL.t5 VP.t4 VDD1.t3 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X13 VTAIL.t10 VN.t5 VDD2.t2 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0.57915 ps=3.84 w=3.51 l=3.77
X14 VTAIL.t8 VN.t6 VDD2.t1 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0.57915 ps=3.84 w=3.51 l=3.77
X15 B.t2 B.t0 B.t1 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0 ps=0 w=3.51 l=3.77
X16 VDD2.t0 VN.t7 VTAIL.t15 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X17 VDD1.t2 VP.t5 VTAIL.t6 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X18 VDD1.t1 VP.t6 VTAIL.t0 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=0.57915 pd=3.84 as=0.57915 ps=3.84 w=3.51 l=3.77
X19 VTAIL.t1 VP.t7 VDD1.t0 w_n5070_n1670# sky130_fd_pr__pfet_01v8 ad=1.3689 pd=7.8 as=0.57915 ps=3.84 w=3.51 l=3.77
R0 B.n357 B.n356 585
R1 B.n355 B.n132 585
R2 B.n354 B.n353 585
R3 B.n352 B.n133 585
R4 B.n351 B.n350 585
R5 B.n349 B.n134 585
R6 B.n348 B.n347 585
R7 B.n346 B.n135 585
R8 B.n345 B.n344 585
R9 B.n343 B.n136 585
R10 B.n342 B.n341 585
R11 B.n340 B.n137 585
R12 B.n339 B.n338 585
R13 B.n337 B.n138 585
R14 B.n336 B.n335 585
R15 B.n334 B.n139 585
R16 B.n333 B.n332 585
R17 B.n330 B.n140 585
R18 B.n329 B.n328 585
R19 B.n327 B.n143 585
R20 B.n326 B.n325 585
R21 B.n324 B.n144 585
R22 B.n323 B.n322 585
R23 B.n321 B.n145 585
R24 B.n320 B.n319 585
R25 B.n318 B.n146 585
R26 B.n316 B.n315 585
R27 B.n314 B.n149 585
R28 B.n313 B.n312 585
R29 B.n311 B.n150 585
R30 B.n310 B.n309 585
R31 B.n308 B.n151 585
R32 B.n307 B.n306 585
R33 B.n305 B.n152 585
R34 B.n304 B.n303 585
R35 B.n302 B.n153 585
R36 B.n301 B.n300 585
R37 B.n299 B.n154 585
R38 B.n298 B.n297 585
R39 B.n296 B.n155 585
R40 B.n295 B.n294 585
R41 B.n293 B.n156 585
R42 B.n292 B.n291 585
R43 B.n358 B.n131 585
R44 B.n360 B.n359 585
R45 B.n361 B.n130 585
R46 B.n363 B.n362 585
R47 B.n364 B.n129 585
R48 B.n366 B.n365 585
R49 B.n367 B.n128 585
R50 B.n369 B.n368 585
R51 B.n370 B.n127 585
R52 B.n372 B.n371 585
R53 B.n373 B.n126 585
R54 B.n375 B.n374 585
R55 B.n376 B.n125 585
R56 B.n378 B.n377 585
R57 B.n379 B.n124 585
R58 B.n381 B.n380 585
R59 B.n382 B.n123 585
R60 B.n384 B.n383 585
R61 B.n385 B.n122 585
R62 B.n387 B.n386 585
R63 B.n388 B.n121 585
R64 B.n390 B.n389 585
R65 B.n391 B.n120 585
R66 B.n393 B.n392 585
R67 B.n394 B.n119 585
R68 B.n396 B.n395 585
R69 B.n397 B.n118 585
R70 B.n399 B.n398 585
R71 B.n400 B.n117 585
R72 B.n402 B.n401 585
R73 B.n403 B.n116 585
R74 B.n405 B.n404 585
R75 B.n406 B.n115 585
R76 B.n408 B.n407 585
R77 B.n409 B.n114 585
R78 B.n411 B.n410 585
R79 B.n412 B.n113 585
R80 B.n414 B.n413 585
R81 B.n415 B.n112 585
R82 B.n417 B.n416 585
R83 B.n418 B.n111 585
R84 B.n420 B.n419 585
R85 B.n421 B.n110 585
R86 B.n423 B.n422 585
R87 B.n424 B.n109 585
R88 B.n426 B.n425 585
R89 B.n427 B.n108 585
R90 B.n429 B.n428 585
R91 B.n430 B.n107 585
R92 B.n432 B.n431 585
R93 B.n433 B.n106 585
R94 B.n435 B.n434 585
R95 B.n436 B.n105 585
R96 B.n438 B.n437 585
R97 B.n439 B.n104 585
R98 B.n441 B.n440 585
R99 B.n442 B.n103 585
R100 B.n444 B.n443 585
R101 B.n445 B.n102 585
R102 B.n447 B.n446 585
R103 B.n448 B.n101 585
R104 B.n450 B.n449 585
R105 B.n451 B.n100 585
R106 B.n453 B.n452 585
R107 B.n454 B.n99 585
R108 B.n456 B.n455 585
R109 B.n457 B.n98 585
R110 B.n459 B.n458 585
R111 B.n460 B.n97 585
R112 B.n462 B.n461 585
R113 B.n463 B.n96 585
R114 B.n465 B.n464 585
R115 B.n466 B.n95 585
R116 B.n468 B.n467 585
R117 B.n469 B.n94 585
R118 B.n471 B.n470 585
R119 B.n472 B.n93 585
R120 B.n474 B.n473 585
R121 B.n475 B.n92 585
R122 B.n477 B.n476 585
R123 B.n478 B.n91 585
R124 B.n480 B.n479 585
R125 B.n481 B.n90 585
R126 B.n483 B.n482 585
R127 B.n484 B.n89 585
R128 B.n486 B.n485 585
R129 B.n487 B.n88 585
R130 B.n489 B.n488 585
R131 B.n490 B.n87 585
R132 B.n492 B.n491 585
R133 B.n493 B.n86 585
R134 B.n495 B.n494 585
R135 B.n496 B.n85 585
R136 B.n498 B.n497 585
R137 B.n499 B.n84 585
R138 B.n501 B.n500 585
R139 B.n502 B.n83 585
R140 B.n504 B.n503 585
R141 B.n505 B.n82 585
R142 B.n507 B.n506 585
R143 B.n508 B.n81 585
R144 B.n510 B.n509 585
R145 B.n511 B.n80 585
R146 B.n513 B.n512 585
R147 B.n514 B.n79 585
R148 B.n516 B.n515 585
R149 B.n517 B.n78 585
R150 B.n519 B.n518 585
R151 B.n520 B.n77 585
R152 B.n522 B.n521 585
R153 B.n523 B.n76 585
R154 B.n525 B.n524 585
R155 B.n526 B.n75 585
R156 B.n528 B.n527 585
R157 B.n529 B.n74 585
R158 B.n531 B.n530 585
R159 B.n532 B.n73 585
R160 B.n534 B.n533 585
R161 B.n535 B.n72 585
R162 B.n537 B.n536 585
R163 B.n538 B.n71 585
R164 B.n540 B.n539 585
R165 B.n541 B.n70 585
R166 B.n543 B.n542 585
R167 B.n544 B.n69 585
R168 B.n546 B.n545 585
R169 B.n547 B.n68 585
R170 B.n549 B.n548 585
R171 B.n550 B.n67 585
R172 B.n552 B.n551 585
R173 B.n553 B.n66 585
R174 B.n555 B.n554 585
R175 B.n556 B.n65 585
R176 B.n558 B.n557 585
R177 B.n559 B.n64 585
R178 B.n561 B.n560 585
R179 B.n562 B.n63 585
R180 B.n564 B.n563 585
R181 B.n629 B.n36 585
R182 B.n628 B.n627 585
R183 B.n626 B.n37 585
R184 B.n625 B.n624 585
R185 B.n623 B.n38 585
R186 B.n622 B.n621 585
R187 B.n620 B.n39 585
R188 B.n619 B.n618 585
R189 B.n617 B.n40 585
R190 B.n616 B.n615 585
R191 B.n614 B.n41 585
R192 B.n613 B.n612 585
R193 B.n611 B.n42 585
R194 B.n610 B.n609 585
R195 B.n608 B.n43 585
R196 B.n607 B.n606 585
R197 B.n605 B.n44 585
R198 B.n604 B.n603 585
R199 B.n602 B.n45 585
R200 B.n601 B.n600 585
R201 B.n599 B.n49 585
R202 B.n598 B.n597 585
R203 B.n596 B.n50 585
R204 B.n595 B.n594 585
R205 B.n593 B.n51 585
R206 B.n592 B.n591 585
R207 B.n589 B.n52 585
R208 B.n588 B.n587 585
R209 B.n586 B.n55 585
R210 B.n585 B.n584 585
R211 B.n583 B.n56 585
R212 B.n582 B.n581 585
R213 B.n580 B.n57 585
R214 B.n579 B.n578 585
R215 B.n577 B.n58 585
R216 B.n576 B.n575 585
R217 B.n574 B.n59 585
R218 B.n573 B.n572 585
R219 B.n571 B.n60 585
R220 B.n570 B.n569 585
R221 B.n568 B.n61 585
R222 B.n567 B.n566 585
R223 B.n565 B.n62 585
R224 B.n631 B.n630 585
R225 B.n632 B.n35 585
R226 B.n634 B.n633 585
R227 B.n635 B.n34 585
R228 B.n637 B.n636 585
R229 B.n638 B.n33 585
R230 B.n640 B.n639 585
R231 B.n641 B.n32 585
R232 B.n643 B.n642 585
R233 B.n644 B.n31 585
R234 B.n646 B.n645 585
R235 B.n647 B.n30 585
R236 B.n649 B.n648 585
R237 B.n650 B.n29 585
R238 B.n652 B.n651 585
R239 B.n653 B.n28 585
R240 B.n655 B.n654 585
R241 B.n656 B.n27 585
R242 B.n658 B.n657 585
R243 B.n659 B.n26 585
R244 B.n661 B.n660 585
R245 B.n662 B.n25 585
R246 B.n664 B.n663 585
R247 B.n665 B.n24 585
R248 B.n667 B.n666 585
R249 B.n668 B.n23 585
R250 B.n670 B.n669 585
R251 B.n671 B.n22 585
R252 B.n673 B.n672 585
R253 B.n674 B.n21 585
R254 B.n676 B.n675 585
R255 B.n677 B.n20 585
R256 B.n679 B.n678 585
R257 B.n680 B.n19 585
R258 B.n682 B.n681 585
R259 B.n683 B.n18 585
R260 B.n685 B.n684 585
R261 B.n686 B.n17 585
R262 B.n688 B.n687 585
R263 B.n689 B.n16 585
R264 B.n691 B.n690 585
R265 B.n692 B.n15 585
R266 B.n694 B.n693 585
R267 B.n695 B.n14 585
R268 B.n697 B.n696 585
R269 B.n698 B.n13 585
R270 B.n700 B.n699 585
R271 B.n701 B.n12 585
R272 B.n703 B.n702 585
R273 B.n704 B.n11 585
R274 B.n706 B.n705 585
R275 B.n707 B.n10 585
R276 B.n709 B.n708 585
R277 B.n710 B.n9 585
R278 B.n712 B.n711 585
R279 B.n713 B.n8 585
R280 B.n715 B.n714 585
R281 B.n716 B.n7 585
R282 B.n718 B.n717 585
R283 B.n719 B.n6 585
R284 B.n721 B.n720 585
R285 B.n722 B.n5 585
R286 B.n724 B.n723 585
R287 B.n725 B.n4 585
R288 B.n727 B.n726 585
R289 B.n728 B.n3 585
R290 B.n730 B.n729 585
R291 B.n731 B.n0 585
R292 B.n2 B.n1 585
R293 B.n191 B.n190 585
R294 B.n193 B.n192 585
R295 B.n194 B.n189 585
R296 B.n196 B.n195 585
R297 B.n197 B.n188 585
R298 B.n199 B.n198 585
R299 B.n200 B.n187 585
R300 B.n202 B.n201 585
R301 B.n203 B.n186 585
R302 B.n205 B.n204 585
R303 B.n206 B.n185 585
R304 B.n208 B.n207 585
R305 B.n209 B.n184 585
R306 B.n211 B.n210 585
R307 B.n212 B.n183 585
R308 B.n214 B.n213 585
R309 B.n215 B.n182 585
R310 B.n217 B.n216 585
R311 B.n218 B.n181 585
R312 B.n220 B.n219 585
R313 B.n221 B.n180 585
R314 B.n223 B.n222 585
R315 B.n224 B.n179 585
R316 B.n226 B.n225 585
R317 B.n227 B.n178 585
R318 B.n229 B.n228 585
R319 B.n230 B.n177 585
R320 B.n232 B.n231 585
R321 B.n233 B.n176 585
R322 B.n235 B.n234 585
R323 B.n236 B.n175 585
R324 B.n238 B.n237 585
R325 B.n239 B.n174 585
R326 B.n241 B.n240 585
R327 B.n242 B.n173 585
R328 B.n244 B.n243 585
R329 B.n245 B.n172 585
R330 B.n247 B.n246 585
R331 B.n248 B.n171 585
R332 B.n250 B.n249 585
R333 B.n251 B.n170 585
R334 B.n253 B.n252 585
R335 B.n254 B.n169 585
R336 B.n256 B.n255 585
R337 B.n257 B.n168 585
R338 B.n259 B.n258 585
R339 B.n260 B.n167 585
R340 B.n262 B.n261 585
R341 B.n263 B.n166 585
R342 B.n265 B.n264 585
R343 B.n266 B.n165 585
R344 B.n268 B.n267 585
R345 B.n269 B.n164 585
R346 B.n271 B.n270 585
R347 B.n272 B.n163 585
R348 B.n274 B.n273 585
R349 B.n275 B.n162 585
R350 B.n277 B.n276 585
R351 B.n278 B.n161 585
R352 B.n280 B.n279 585
R353 B.n281 B.n160 585
R354 B.n283 B.n282 585
R355 B.n284 B.n159 585
R356 B.n286 B.n285 585
R357 B.n287 B.n158 585
R358 B.n289 B.n288 585
R359 B.n290 B.n157 585
R360 B.n291 B.n290 473.281
R361 B.n358 B.n357 473.281
R362 B.n563 B.n62 473.281
R363 B.n630 B.n629 473.281
R364 B.n733 B.n732 256.663
R365 B.n732 B.n731 235.042
R366 B.n732 B.n2 235.042
R367 B.n147 B.t9 231.758
R368 B.n141 B.t0 231.758
R369 B.n53 B.t3 231.758
R370 B.n46 B.t6 231.758
R371 B.n141 B.t1 207.977
R372 B.n53 B.t5 207.977
R373 B.n147 B.t10 207.976
R374 B.n46 B.t8 207.976
R375 B.n291 B.n156 163.367
R376 B.n295 B.n156 163.367
R377 B.n296 B.n295 163.367
R378 B.n297 B.n296 163.367
R379 B.n297 B.n154 163.367
R380 B.n301 B.n154 163.367
R381 B.n302 B.n301 163.367
R382 B.n303 B.n302 163.367
R383 B.n303 B.n152 163.367
R384 B.n307 B.n152 163.367
R385 B.n308 B.n307 163.367
R386 B.n309 B.n308 163.367
R387 B.n309 B.n150 163.367
R388 B.n313 B.n150 163.367
R389 B.n314 B.n313 163.367
R390 B.n315 B.n314 163.367
R391 B.n315 B.n146 163.367
R392 B.n320 B.n146 163.367
R393 B.n321 B.n320 163.367
R394 B.n322 B.n321 163.367
R395 B.n322 B.n144 163.367
R396 B.n326 B.n144 163.367
R397 B.n327 B.n326 163.367
R398 B.n328 B.n327 163.367
R399 B.n328 B.n140 163.367
R400 B.n333 B.n140 163.367
R401 B.n334 B.n333 163.367
R402 B.n335 B.n334 163.367
R403 B.n335 B.n138 163.367
R404 B.n339 B.n138 163.367
R405 B.n340 B.n339 163.367
R406 B.n341 B.n340 163.367
R407 B.n341 B.n136 163.367
R408 B.n345 B.n136 163.367
R409 B.n346 B.n345 163.367
R410 B.n347 B.n346 163.367
R411 B.n347 B.n134 163.367
R412 B.n351 B.n134 163.367
R413 B.n352 B.n351 163.367
R414 B.n353 B.n352 163.367
R415 B.n353 B.n132 163.367
R416 B.n357 B.n132 163.367
R417 B.n563 B.n562 163.367
R418 B.n562 B.n561 163.367
R419 B.n561 B.n64 163.367
R420 B.n557 B.n64 163.367
R421 B.n557 B.n556 163.367
R422 B.n556 B.n555 163.367
R423 B.n555 B.n66 163.367
R424 B.n551 B.n66 163.367
R425 B.n551 B.n550 163.367
R426 B.n550 B.n549 163.367
R427 B.n549 B.n68 163.367
R428 B.n545 B.n68 163.367
R429 B.n545 B.n544 163.367
R430 B.n544 B.n543 163.367
R431 B.n543 B.n70 163.367
R432 B.n539 B.n70 163.367
R433 B.n539 B.n538 163.367
R434 B.n538 B.n537 163.367
R435 B.n537 B.n72 163.367
R436 B.n533 B.n72 163.367
R437 B.n533 B.n532 163.367
R438 B.n532 B.n531 163.367
R439 B.n531 B.n74 163.367
R440 B.n527 B.n74 163.367
R441 B.n527 B.n526 163.367
R442 B.n526 B.n525 163.367
R443 B.n525 B.n76 163.367
R444 B.n521 B.n76 163.367
R445 B.n521 B.n520 163.367
R446 B.n520 B.n519 163.367
R447 B.n519 B.n78 163.367
R448 B.n515 B.n78 163.367
R449 B.n515 B.n514 163.367
R450 B.n514 B.n513 163.367
R451 B.n513 B.n80 163.367
R452 B.n509 B.n80 163.367
R453 B.n509 B.n508 163.367
R454 B.n508 B.n507 163.367
R455 B.n507 B.n82 163.367
R456 B.n503 B.n82 163.367
R457 B.n503 B.n502 163.367
R458 B.n502 B.n501 163.367
R459 B.n501 B.n84 163.367
R460 B.n497 B.n84 163.367
R461 B.n497 B.n496 163.367
R462 B.n496 B.n495 163.367
R463 B.n495 B.n86 163.367
R464 B.n491 B.n86 163.367
R465 B.n491 B.n490 163.367
R466 B.n490 B.n489 163.367
R467 B.n489 B.n88 163.367
R468 B.n485 B.n88 163.367
R469 B.n485 B.n484 163.367
R470 B.n484 B.n483 163.367
R471 B.n483 B.n90 163.367
R472 B.n479 B.n90 163.367
R473 B.n479 B.n478 163.367
R474 B.n478 B.n477 163.367
R475 B.n477 B.n92 163.367
R476 B.n473 B.n92 163.367
R477 B.n473 B.n472 163.367
R478 B.n472 B.n471 163.367
R479 B.n471 B.n94 163.367
R480 B.n467 B.n94 163.367
R481 B.n467 B.n466 163.367
R482 B.n466 B.n465 163.367
R483 B.n465 B.n96 163.367
R484 B.n461 B.n96 163.367
R485 B.n461 B.n460 163.367
R486 B.n460 B.n459 163.367
R487 B.n459 B.n98 163.367
R488 B.n455 B.n98 163.367
R489 B.n455 B.n454 163.367
R490 B.n454 B.n453 163.367
R491 B.n453 B.n100 163.367
R492 B.n449 B.n100 163.367
R493 B.n449 B.n448 163.367
R494 B.n448 B.n447 163.367
R495 B.n447 B.n102 163.367
R496 B.n443 B.n102 163.367
R497 B.n443 B.n442 163.367
R498 B.n442 B.n441 163.367
R499 B.n441 B.n104 163.367
R500 B.n437 B.n104 163.367
R501 B.n437 B.n436 163.367
R502 B.n436 B.n435 163.367
R503 B.n435 B.n106 163.367
R504 B.n431 B.n106 163.367
R505 B.n431 B.n430 163.367
R506 B.n430 B.n429 163.367
R507 B.n429 B.n108 163.367
R508 B.n425 B.n108 163.367
R509 B.n425 B.n424 163.367
R510 B.n424 B.n423 163.367
R511 B.n423 B.n110 163.367
R512 B.n419 B.n110 163.367
R513 B.n419 B.n418 163.367
R514 B.n418 B.n417 163.367
R515 B.n417 B.n112 163.367
R516 B.n413 B.n112 163.367
R517 B.n413 B.n412 163.367
R518 B.n412 B.n411 163.367
R519 B.n411 B.n114 163.367
R520 B.n407 B.n114 163.367
R521 B.n407 B.n406 163.367
R522 B.n406 B.n405 163.367
R523 B.n405 B.n116 163.367
R524 B.n401 B.n116 163.367
R525 B.n401 B.n400 163.367
R526 B.n400 B.n399 163.367
R527 B.n399 B.n118 163.367
R528 B.n395 B.n118 163.367
R529 B.n395 B.n394 163.367
R530 B.n394 B.n393 163.367
R531 B.n393 B.n120 163.367
R532 B.n389 B.n120 163.367
R533 B.n389 B.n388 163.367
R534 B.n388 B.n387 163.367
R535 B.n387 B.n122 163.367
R536 B.n383 B.n122 163.367
R537 B.n383 B.n382 163.367
R538 B.n382 B.n381 163.367
R539 B.n381 B.n124 163.367
R540 B.n377 B.n124 163.367
R541 B.n377 B.n376 163.367
R542 B.n376 B.n375 163.367
R543 B.n375 B.n126 163.367
R544 B.n371 B.n126 163.367
R545 B.n371 B.n370 163.367
R546 B.n370 B.n369 163.367
R547 B.n369 B.n128 163.367
R548 B.n365 B.n128 163.367
R549 B.n365 B.n364 163.367
R550 B.n364 B.n363 163.367
R551 B.n363 B.n130 163.367
R552 B.n359 B.n130 163.367
R553 B.n359 B.n358 163.367
R554 B.n629 B.n628 163.367
R555 B.n628 B.n37 163.367
R556 B.n624 B.n37 163.367
R557 B.n624 B.n623 163.367
R558 B.n623 B.n622 163.367
R559 B.n622 B.n39 163.367
R560 B.n618 B.n39 163.367
R561 B.n618 B.n617 163.367
R562 B.n617 B.n616 163.367
R563 B.n616 B.n41 163.367
R564 B.n612 B.n41 163.367
R565 B.n612 B.n611 163.367
R566 B.n611 B.n610 163.367
R567 B.n610 B.n43 163.367
R568 B.n606 B.n43 163.367
R569 B.n606 B.n605 163.367
R570 B.n605 B.n604 163.367
R571 B.n604 B.n45 163.367
R572 B.n600 B.n45 163.367
R573 B.n600 B.n599 163.367
R574 B.n599 B.n598 163.367
R575 B.n598 B.n50 163.367
R576 B.n594 B.n50 163.367
R577 B.n594 B.n593 163.367
R578 B.n593 B.n592 163.367
R579 B.n592 B.n52 163.367
R580 B.n587 B.n52 163.367
R581 B.n587 B.n586 163.367
R582 B.n586 B.n585 163.367
R583 B.n585 B.n56 163.367
R584 B.n581 B.n56 163.367
R585 B.n581 B.n580 163.367
R586 B.n580 B.n579 163.367
R587 B.n579 B.n58 163.367
R588 B.n575 B.n58 163.367
R589 B.n575 B.n574 163.367
R590 B.n574 B.n573 163.367
R591 B.n573 B.n60 163.367
R592 B.n569 B.n60 163.367
R593 B.n569 B.n568 163.367
R594 B.n568 B.n567 163.367
R595 B.n567 B.n62 163.367
R596 B.n630 B.n35 163.367
R597 B.n634 B.n35 163.367
R598 B.n635 B.n634 163.367
R599 B.n636 B.n635 163.367
R600 B.n636 B.n33 163.367
R601 B.n640 B.n33 163.367
R602 B.n641 B.n640 163.367
R603 B.n642 B.n641 163.367
R604 B.n642 B.n31 163.367
R605 B.n646 B.n31 163.367
R606 B.n647 B.n646 163.367
R607 B.n648 B.n647 163.367
R608 B.n648 B.n29 163.367
R609 B.n652 B.n29 163.367
R610 B.n653 B.n652 163.367
R611 B.n654 B.n653 163.367
R612 B.n654 B.n27 163.367
R613 B.n658 B.n27 163.367
R614 B.n659 B.n658 163.367
R615 B.n660 B.n659 163.367
R616 B.n660 B.n25 163.367
R617 B.n664 B.n25 163.367
R618 B.n665 B.n664 163.367
R619 B.n666 B.n665 163.367
R620 B.n666 B.n23 163.367
R621 B.n670 B.n23 163.367
R622 B.n671 B.n670 163.367
R623 B.n672 B.n671 163.367
R624 B.n672 B.n21 163.367
R625 B.n676 B.n21 163.367
R626 B.n677 B.n676 163.367
R627 B.n678 B.n677 163.367
R628 B.n678 B.n19 163.367
R629 B.n682 B.n19 163.367
R630 B.n683 B.n682 163.367
R631 B.n684 B.n683 163.367
R632 B.n684 B.n17 163.367
R633 B.n688 B.n17 163.367
R634 B.n689 B.n688 163.367
R635 B.n690 B.n689 163.367
R636 B.n690 B.n15 163.367
R637 B.n694 B.n15 163.367
R638 B.n695 B.n694 163.367
R639 B.n696 B.n695 163.367
R640 B.n696 B.n13 163.367
R641 B.n700 B.n13 163.367
R642 B.n701 B.n700 163.367
R643 B.n702 B.n701 163.367
R644 B.n702 B.n11 163.367
R645 B.n706 B.n11 163.367
R646 B.n707 B.n706 163.367
R647 B.n708 B.n707 163.367
R648 B.n708 B.n9 163.367
R649 B.n712 B.n9 163.367
R650 B.n713 B.n712 163.367
R651 B.n714 B.n713 163.367
R652 B.n714 B.n7 163.367
R653 B.n718 B.n7 163.367
R654 B.n719 B.n718 163.367
R655 B.n720 B.n719 163.367
R656 B.n720 B.n5 163.367
R657 B.n724 B.n5 163.367
R658 B.n725 B.n724 163.367
R659 B.n726 B.n725 163.367
R660 B.n726 B.n3 163.367
R661 B.n730 B.n3 163.367
R662 B.n731 B.n730 163.367
R663 B.n190 B.n2 163.367
R664 B.n193 B.n190 163.367
R665 B.n194 B.n193 163.367
R666 B.n195 B.n194 163.367
R667 B.n195 B.n188 163.367
R668 B.n199 B.n188 163.367
R669 B.n200 B.n199 163.367
R670 B.n201 B.n200 163.367
R671 B.n201 B.n186 163.367
R672 B.n205 B.n186 163.367
R673 B.n206 B.n205 163.367
R674 B.n207 B.n206 163.367
R675 B.n207 B.n184 163.367
R676 B.n211 B.n184 163.367
R677 B.n212 B.n211 163.367
R678 B.n213 B.n212 163.367
R679 B.n213 B.n182 163.367
R680 B.n217 B.n182 163.367
R681 B.n218 B.n217 163.367
R682 B.n219 B.n218 163.367
R683 B.n219 B.n180 163.367
R684 B.n223 B.n180 163.367
R685 B.n224 B.n223 163.367
R686 B.n225 B.n224 163.367
R687 B.n225 B.n178 163.367
R688 B.n229 B.n178 163.367
R689 B.n230 B.n229 163.367
R690 B.n231 B.n230 163.367
R691 B.n231 B.n176 163.367
R692 B.n235 B.n176 163.367
R693 B.n236 B.n235 163.367
R694 B.n237 B.n236 163.367
R695 B.n237 B.n174 163.367
R696 B.n241 B.n174 163.367
R697 B.n242 B.n241 163.367
R698 B.n243 B.n242 163.367
R699 B.n243 B.n172 163.367
R700 B.n247 B.n172 163.367
R701 B.n248 B.n247 163.367
R702 B.n249 B.n248 163.367
R703 B.n249 B.n170 163.367
R704 B.n253 B.n170 163.367
R705 B.n254 B.n253 163.367
R706 B.n255 B.n254 163.367
R707 B.n255 B.n168 163.367
R708 B.n259 B.n168 163.367
R709 B.n260 B.n259 163.367
R710 B.n261 B.n260 163.367
R711 B.n261 B.n166 163.367
R712 B.n265 B.n166 163.367
R713 B.n266 B.n265 163.367
R714 B.n267 B.n266 163.367
R715 B.n267 B.n164 163.367
R716 B.n271 B.n164 163.367
R717 B.n272 B.n271 163.367
R718 B.n273 B.n272 163.367
R719 B.n273 B.n162 163.367
R720 B.n277 B.n162 163.367
R721 B.n278 B.n277 163.367
R722 B.n279 B.n278 163.367
R723 B.n279 B.n160 163.367
R724 B.n283 B.n160 163.367
R725 B.n284 B.n283 163.367
R726 B.n285 B.n284 163.367
R727 B.n285 B.n158 163.367
R728 B.n289 B.n158 163.367
R729 B.n290 B.n289 163.367
R730 B.n142 B.t2 128.463
R731 B.n54 B.t4 128.463
R732 B.n148 B.t11 128.459
R733 B.n47 B.t7 128.459
R734 B.n148 B.n147 79.5157
R735 B.n142 B.n141 79.5157
R736 B.n54 B.n53 79.5157
R737 B.n47 B.n46 79.5157
R738 B.n317 B.n148 59.5399
R739 B.n331 B.n142 59.5399
R740 B.n590 B.n54 59.5399
R741 B.n48 B.n47 59.5399
R742 B.n631 B.n36 30.7517
R743 B.n565 B.n564 30.7517
R744 B.n356 B.n131 30.7517
R745 B.n292 B.n157 30.7517
R746 B B.n733 18.0485
R747 B.n632 B.n631 10.6151
R748 B.n633 B.n632 10.6151
R749 B.n633 B.n34 10.6151
R750 B.n637 B.n34 10.6151
R751 B.n638 B.n637 10.6151
R752 B.n639 B.n638 10.6151
R753 B.n639 B.n32 10.6151
R754 B.n643 B.n32 10.6151
R755 B.n644 B.n643 10.6151
R756 B.n645 B.n644 10.6151
R757 B.n645 B.n30 10.6151
R758 B.n649 B.n30 10.6151
R759 B.n650 B.n649 10.6151
R760 B.n651 B.n650 10.6151
R761 B.n651 B.n28 10.6151
R762 B.n655 B.n28 10.6151
R763 B.n656 B.n655 10.6151
R764 B.n657 B.n656 10.6151
R765 B.n657 B.n26 10.6151
R766 B.n661 B.n26 10.6151
R767 B.n662 B.n661 10.6151
R768 B.n663 B.n662 10.6151
R769 B.n663 B.n24 10.6151
R770 B.n667 B.n24 10.6151
R771 B.n668 B.n667 10.6151
R772 B.n669 B.n668 10.6151
R773 B.n669 B.n22 10.6151
R774 B.n673 B.n22 10.6151
R775 B.n674 B.n673 10.6151
R776 B.n675 B.n674 10.6151
R777 B.n675 B.n20 10.6151
R778 B.n679 B.n20 10.6151
R779 B.n680 B.n679 10.6151
R780 B.n681 B.n680 10.6151
R781 B.n681 B.n18 10.6151
R782 B.n685 B.n18 10.6151
R783 B.n686 B.n685 10.6151
R784 B.n687 B.n686 10.6151
R785 B.n687 B.n16 10.6151
R786 B.n691 B.n16 10.6151
R787 B.n692 B.n691 10.6151
R788 B.n693 B.n692 10.6151
R789 B.n693 B.n14 10.6151
R790 B.n697 B.n14 10.6151
R791 B.n698 B.n697 10.6151
R792 B.n699 B.n698 10.6151
R793 B.n699 B.n12 10.6151
R794 B.n703 B.n12 10.6151
R795 B.n704 B.n703 10.6151
R796 B.n705 B.n704 10.6151
R797 B.n705 B.n10 10.6151
R798 B.n709 B.n10 10.6151
R799 B.n710 B.n709 10.6151
R800 B.n711 B.n710 10.6151
R801 B.n711 B.n8 10.6151
R802 B.n715 B.n8 10.6151
R803 B.n716 B.n715 10.6151
R804 B.n717 B.n716 10.6151
R805 B.n717 B.n6 10.6151
R806 B.n721 B.n6 10.6151
R807 B.n722 B.n721 10.6151
R808 B.n723 B.n722 10.6151
R809 B.n723 B.n4 10.6151
R810 B.n727 B.n4 10.6151
R811 B.n728 B.n727 10.6151
R812 B.n729 B.n728 10.6151
R813 B.n729 B.n0 10.6151
R814 B.n627 B.n36 10.6151
R815 B.n627 B.n626 10.6151
R816 B.n626 B.n625 10.6151
R817 B.n625 B.n38 10.6151
R818 B.n621 B.n38 10.6151
R819 B.n621 B.n620 10.6151
R820 B.n620 B.n619 10.6151
R821 B.n619 B.n40 10.6151
R822 B.n615 B.n40 10.6151
R823 B.n615 B.n614 10.6151
R824 B.n614 B.n613 10.6151
R825 B.n613 B.n42 10.6151
R826 B.n609 B.n42 10.6151
R827 B.n609 B.n608 10.6151
R828 B.n608 B.n607 10.6151
R829 B.n607 B.n44 10.6151
R830 B.n603 B.n602 10.6151
R831 B.n602 B.n601 10.6151
R832 B.n601 B.n49 10.6151
R833 B.n597 B.n49 10.6151
R834 B.n597 B.n596 10.6151
R835 B.n596 B.n595 10.6151
R836 B.n595 B.n51 10.6151
R837 B.n591 B.n51 10.6151
R838 B.n589 B.n588 10.6151
R839 B.n588 B.n55 10.6151
R840 B.n584 B.n55 10.6151
R841 B.n584 B.n583 10.6151
R842 B.n583 B.n582 10.6151
R843 B.n582 B.n57 10.6151
R844 B.n578 B.n57 10.6151
R845 B.n578 B.n577 10.6151
R846 B.n577 B.n576 10.6151
R847 B.n576 B.n59 10.6151
R848 B.n572 B.n59 10.6151
R849 B.n572 B.n571 10.6151
R850 B.n571 B.n570 10.6151
R851 B.n570 B.n61 10.6151
R852 B.n566 B.n61 10.6151
R853 B.n566 B.n565 10.6151
R854 B.n564 B.n63 10.6151
R855 B.n560 B.n63 10.6151
R856 B.n560 B.n559 10.6151
R857 B.n559 B.n558 10.6151
R858 B.n558 B.n65 10.6151
R859 B.n554 B.n65 10.6151
R860 B.n554 B.n553 10.6151
R861 B.n553 B.n552 10.6151
R862 B.n552 B.n67 10.6151
R863 B.n548 B.n67 10.6151
R864 B.n548 B.n547 10.6151
R865 B.n547 B.n546 10.6151
R866 B.n546 B.n69 10.6151
R867 B.n542 B.n69 10.6151
R868 B.n542 B.n541 10.6151
R869 B.n541 B.n540 10.6151
R870 B.n540 B.n71 10.6151
R871 B.n536 B.n71 10.6151
R872 B.n536 B.n535 10.6151
R873 B.n535 B.n534 10.6151
R874 B.n534 B.n73 10.6151
R875 B.n530 B.n73 10.6151
R876 B.n530 B.n529 10.6151
R877 B.n529 B.n528 10.6151
R878 B.n528 B.n75 10.6151
R879 B.n524 B.n75 10.6151
R880 B.n524 B.n523 10.6151
R881 B.n523 B.n522 10.6151
R882 B.n522 B.n77 10.6151
R883 B.n518 B.n77 10.6151
R884 B.n518 B.n517 10.6151
R885 B.n517 B.n516 10.6151
R886 B.n516 B.n79 10.6151
R887 B.n512 B.n79 10.6151
R888 B.n512 B.n511 10.6151
R889 B.n511 B.n510 10.6151
R890 B.n510 B.n81 10.6151
R891 B.n506 B.n81 10.6151
R892 B.n506 B.n505 10.6151
R893 B.n505 B.n504 10.6151
R894 B.n504 B.n83 10.6151
R895 B.n500 B.n83 10.6151
R896 B.n500 B.n499 10.6151
R897 B.n499 B.n498 10.6151
R898 B.n498 B.n85 10.6151
R899 B.n494 B.n85 10.6151
R900 B.n494 B.n493 10.6151
R901 B.n493 B.n492 10.6151
R902 B.n492 B.n87 10.6151
R903 B.n488 B.n87 10.6151
R904 B.n488 B.n487 10.6151
R905 B.n487 B.n486 10.6151
R906 B.n486 B.n89 10.6151
R907 B.n482 B.n89 10.6151
R908 B.n482 B.n481 10.6151
R909 B.n481 B.n480 10.6151
R910 B.n480 B.n91 10.6151
R911 B.n476 B.n91 10.6151
R912 B.n476 B.n475 10.6151
R913 B.n475 B.n474 10.6151
R914 B.n474 B.n93 10.6151
R915 B.n470 B.n93 10.6151
R916 B.n470 B.n469 10.6151
R917 B.n469 B.n468 10.6151
R918 B.n468 B.n95 10.6151
R919 B.n464 B.n95 10.6151
R920 B.n464 B.n463 10.6151
R921 B.n463 B.n462 10.6151
R922 B.n462 B.n97 10.6151
R923 B.n458 B.n97 10.6151
R924 B.n458 B.n457 10.6151
R925 B.n457 B.n456 10.6151
R926 B.n456 B.n99 10.6151
R927 B.n452 B.n99 10.6151
R928 B.n452 B.n451 10.6151
R929 B.n451 B.n450 10.6151
R930 B.n450 B.n101 10.6151
R931 B.n446 B.n101 10.6151
R932 B.n446 B.n445 10.6151
R933 B.n445 B.n444 10.6151
R934 B.n444 B.n103 10.6151
R935 B.n440 B.n103 10.6151
R936 B.n440 B.n439 10.6151
R937 B.n439 B.n438 10.6151
R938 B.n438 B.n105 10.6151
R939 B.n434 B.n105 10.6151
R940 B.n434 B.n433 10.6151
R941 B.n433 B.n432 10.6151
R942 B.n432 B.n107 10.6151
R943 B.n428 B.n107 10.6151
R944 B.n428 B.n427 10.6151
R945 B.n427 B.n426 10.6151
R946 B.n426 B.n109 10.6151
R947 B.n422 B.n109 10.6151
R948 B.n422 B.n421 10.6151
R949 B.n421 B.n420 10.6151
R950 B.n420 B.n111 10.6151
R951 B.n416 B.n111 10.6151
R952 B.n416 B.n415 10.6151
R953 B.n415 B.n414 10.6151
R954 B.n414 B.n113 10.6151
R955 B.n410 B.n113 10.6151
R956 B.n410 B.n409 10.6151
R957 B.n409 B.n408 10.6151
R958 B.n408 B.n115 10.6151
R959 B.n404 B.n115 10.6151
R960 B.n404 B.n403 10.6151
R961 B.n403 B.n402 10.6151
R962 B.n402 B.n117 10.6151
R963 B.n398 B.n117 10.6151
R964 B.n398 B.n397 10.6151
R965 B.n397 B.n396 10.6151
R966 B.n396 B.n119 10.6151
R967 B.n392 B.n119 10.6151
R968 B.n392 B.n391 10.6151
R969 B.n391 B.n390 10.6151
R970 B.n390 B.n121 10.6151
R971 B.n386 B.n121 10.6151
R972 B.n386 B.n385 10.6151
R973 B.n385 B.n384 10.6151
R974 B.n384 B.n123 10.6151
R975 B.n380 B.n123 10.6151
R976 B.n380 B.n379 10.6151
R977 B.n379 B.n378 10.6151
R978 B.n378 B.n125 10.6151
R979 B.n374 B.n125 10.6151
R980 B.n374 B.n373 10.6151
R981 B.n373 B.n372 10.6151
R982 B.n372 B.n127 10.6151
R983 B.n368 B.n127 10.6151
R984 B.n368 B.n367 10.6151
R985 B.n367 B.n366 10.6151
R986 B.n366 B.n129 10.6151
R987 B.n362 B.n129 10.6151
R988 B.n362 B.n361 10.6151
R989 B.n361 B.n360 10.6151
R990 B.n360 B.n131 10.6151
R991 B.n191 B.n1 10.6151
R992 B.n192 B.n191 10.6151
R993 B.n192 B.n189 10.6151
R994 B.n196 B.n189 10.6151
R995 B.n197 B.n196 10.6151
R996 B.n198 B.n197 10.6151
R997 B.n198 B.n187 10.6151
R998 B.n202 B.n187 10.6151
R999 B.n203 B.n202 10.6151
R1000 B.n204 B.n203 10.6151
R1001 B.n204 B.n185 10.6151
R1002 B.n208 B.n185 10.6151
R1003 B.n209 B.n208 10.6151
R1004 B.n210 B.n209 10.6151
R1005 B.n210 B.n183 10.6151
R1006 B.n214 B.n183 10.6151
R1007 B.n215 B.n214 10.6151
R1008 B.n216 B.n215 10.6151
R1009 B.n216 B.n181 10.6151
R1010 B.n220 B.n181 10.6151
R1011 B.n221 B.n220 10.6151
R1012 B.n222 B.n221 10.6151
R1013 B.n222 B.n179 10.6151
R1014 B.n226 B.n179 10.6151
R1015 B.n227 B.n226 10.6151
R1016 B.n228 B.n227 10.6151
R1017 B.n228 B.n177 10.6151
R1018 B.n232 B.n177 10.6151
R1019 B.n233 B.n232 10.6151
R1020 B.n234 B.n233 10.6151
R1021 B.n234 B.n175 10.6151
R1022 B.n238 B.n175 10.6151
R1023 B.n239 B.n238 10.6151
R1024 B.n240 B.n239 10.6151
R1025 B.n240 B.n173 10.6151
R1026 B.n244 B.n173 10.6151
R1027 B.n245 B.n244 10.6151
R1028 B.n246 B.n245 10.6151
R1029 B.n246 B.n171 10.6151
R1030 B.n250 B.n171 10.6151
R1031 B.n251 B.n250 10.6151
R1032 B.n252 B.n251 10.6151
R1033 B.n252 B.n169 10.6151
R1034 B.n256 B.n169 10.6151
R1035 B.n257 B.n256 10.6151
R1036 B.n258 B.n257 10.6151
R1037 B.n258 B.n167 10.6151
R1038 B.n262 B.n167 10.6151
R1039 B.n263 B.n262 10.6151
R1040 B.n264 B.n263 10.6151
R1041 B.n264 B.n165 10.6151
R1042 B.n268 B.n165 10.6151
R1043 B.n269 B.n268 10.6151
R1044 B.n270 B.n269 10.6151
R1045 B.n270 B.n163 10.6151
R1046 B.n274 B.n163 10.6151
R1047 B.n275 B.n274 10.6151
R1048 B.n276 B.n275 10.6151
R1049 B.n276 B.n161 10.6151
R1050 B.n280 B.n161 10.6151
R1051 B.n281 B.n280 10.6151
R1052 B.n282 B.n281 10.6151
R1053 B.n282 B.n159 10.6151
R1054 B.n286 B.n159 10.6151
R1055 B.n287 B.n286 10.6151
R1056 B.n288 B.n287 10.6151
R1057 B.n288 B.n157 10.6151
R1058 B.n293 B.n292 10.6151
R1059 B.n294 B.n293 10.6151
R1060 B.n294 B.n155 10.6151
R1061 B.n298 B.n155 10.6151
R1062 B.n299 B.n298 10.6151
R1063 B.n300 B.n299 10.6151
R1064 B.n300 B.n153 10.6151
R1065 B.n304 B.n153 10.6151
R1066 B.n305 B.n304 10.6151
R1067 B.n306 B.n305 10.6151
R1068 B.n306 B.n151 10.6151
R1069 B.n310 B.n151 10.6151
R1070 B.n311 B.n310 10.6151
R1071 B.n312 B.n311 10.6151
R1072 B.n312 B.n149 10.6151
R1073 B.n316 B.n149 10.6151
R1074 B.n319 B.n318 10.6151
R1075 B.n319 B.n145 10.6151
R1076 B.n323 B.n145 10.6151
R1077 B.n324 B.n323 10.6151
R1078 B.n325 B.n324 10.6151
R1079 B.n325 B.n143 10.6151
R1080 B.n329 B.n143 10.6151
R1081 B.n330 B.n329 10.6151
R1082 B.n332 B.n139 10.6151
R1083 B.n336 B.n139 10.6151
R1084 B.n337 B.n336 10.6151
R1085 B.n338 B.n337 10.6151
R1086 B.n338 B.n137 10.6151
R1087 B.n342 B.n137 10.6151
R1088 B.n343 B.n342 10.6151
R1089 B.n344 B.n343 10.6151
R1090 B.n344 B.n135 10.6151
R1091 B.n348 B.n135 10.6151
R1092 B.n349 B.n348 10.6151
R1093 B.n350 B.n349 10.6151
R1094 B.n350 B.n133 10.6151
R1095 B.n354 B.n133 10.6151
R1096 B.n355 B.n354 10.6151
R1097 B.n356 B.n355 10.6151
R1098 B.n733 B.n0 8.11757
R1099 B.n733 B.n1 8.11757
R1100 B.n603 B.n48 6.5566
R1101 B.n591 B.n590 6.5566
R1102 B.n318 B.n317 6.5566
R1103 B.n331 B.n330 6.5566
R1104 B.n48 B.n44 4.05904
R1105 B.n590 B.n589 4.05904
R1106 B.n317 B.n316 4.05904
R1107 B.n332 B.n331 4.05904
R1108 VN.n76 VN.n75 161.3
R1109 VN.n74 VN.n40 161.3
R1110 VN.n73 VN.n72 161.3
R1111 VN.n71 VN.n41 161.3
R1112 VN.n70 VN.n69 161.3
R1113 VN.n68 VN.n42 161.3
R1114 VN.n67 VN.n66 161.3
R1115 VN.n65 VN.n43 161.3
R1116 VN.n64 VN.n63 161.3
R1117 VN.n62 VN.n44 161.3
R1118 VN.n61 VN.n60 161.3
R1119 VN.n59 VN.n46 161.3
R1120 VN.n58 VN.n57 161.3
R1121 VN.n56 VN.n47 161.3
R1122 VN.n55 VN.n54 161.3
R1123 VN.n53 VN.n48 161.3
R1124 VN.n52 VN.n51 161.3
R1125 VN.n37 VN.n36 161.3
R1126 VN.n35 VN.n1 161.3
R1127 VN.n34 VN.n33 161.3
R1128 VN.n32 VN.n2 161.3
R1129 VN.n31 VN.n30 161.3
R1130 VN.n29 VN.n3 161.3
R1131 VN.n28 VN.n27 161.3
R1132 VN.n26 VN.n4 161.3
R1133 VN.n25 VN.n24 161.3
R1134 VN.n22 VN.n5 161.3
R1135 VN.n21 VN.n20 161.3
R1136 VN.n19 VN.n6 161.3
R1137 VN.n18 VN.n17 161.3
R1138 VN.n16 VN.n7 161.3
R1139 VN.n15 VN.n14 161.3
R1140 VN.n13 VN.n8 161.3
R1141 VN.n12 VN.n11 161.3
R1142 VN.n38 VN.n0 82.7273
R1143 VN.n77 VN.n39 82.7273
R1144 VN.n50 VN.n49 72.3975
R1145 VN.n10 VN.n9 72.3975
R1146 VN.n49 VN.t1 55.3381
R1147 VN.n9 VN.t5 55.3381
R1148 VN VN.n77 50.2177
R1149 VN.n30 VN.n2 50.2061
R1150 VN.n69 VN.n41 50.2061
R1151 VN.n17 VN.n16 40.4934
R1152 VN.n17 VN.n6 40.4934
R1153 VN.n57 VN.n56 40.4934
R1154 VN.n57 VN.n46 40.4934
R1155 VN.n30 VN.n29 30.7807
R1156 VN.n69 VN.n68 30.7807
R1157 VN.n11 VN.n8 24.4675
R1158 VN.n15 VN.n8 24.4675
R1159 VN.n16 VN.n15 24.4675
R1160 VN.n21 VN.n6 24.4675
R1161 VN.n22 VN.n21 24.4675
R1162 VN.n24 VN.n22 24.4675
R1163 VN.n28 VN.n4 24.4675
R1164 VN.n29 VN.n28 24.4675
R1165 VN.n34 VN.n2 24.4675
R1166 VN.n35 VN.n34 24.4675
R1167 VN.n36 VN.n35 24.4675
R1168 VN.n56 VN.n55 24.4675
R1169 VN.n55 VN.n48 24.4675
R1170 VN.n51 VN.n48 24.4675
R1171 VN.n68 VN.n67 24.4675
R1172 VN.n67 VN.n43 24.4675
R1173 VN.n63 VN.n62 24.4675
R1174 VN.n62 VN.n61 24.4675
R1175 VN.n61 VN.n46 24.4675
R1176 VN.n75 VN.n74 24.4675
R1177 VN.n74 VN.n73 24.4675
R1178 VN.n73 VN.n41 24.4675
R1179 VN.n10 VN.t7 22.4384
R1180 VN.n23 VN.t3 22.4384
R1181 VN.n0 VN.t0 22.4384
R1182 VN.n50 VN.t2 22.4384
R1183 VN.n45 VN.t4 22.4384
R1184 VN.n39 VN.t6 22.4384
R1185 VN.n23 VN.n4 22.0208
R1186 VN.n45 VN.n43 22.0208
R1187 VN.n36 VN.n0 7.3406
R1188 VN.n75 VN.n39 7.3406
R1189 VN.n52 VN.n49 3.236
R1190 VN.n12 VN.n9 3.236
R1191 VN.n11 VN.n10 2.4472
R1192 VN.n24 VN.n23 2.4472
R1193 VN.n51 VN.n50 2.4472
R1194 VN.n63 VN.n45 2.4472
R1195 VN.n77 VN.n76 0.354971
R1196 VN.n38 VN.n37 0.354971
R1197 VN VN.n38 0.26696
R1198 VN.n76 VN.n40 0.189894
R1199 VN.n72 VN.n40 0.189894
R1200 VN.n72 VN.n71 0.189894
R1201 VN.n71 VN.n70 0.189894
R1202 VN.n70 VN.n42 0.189894
R1203 VN.n66 VN.n42 0.189894
R1204 VN.n66 VN.n65 0.189894
R1205 VN.n65 VN.n64 0.189894
R1206 VN.n64 VN.n44 0.189894
R1207 VN.n60 VN.n44 0.189894
R1208 VN.n60 VN.n59 0.189894
R1209 VN.n59 VN.n58 0.189894
R1210 VN.n58 VN.n47 0.189894
R1211 VN.n54 VN.n47 0.189894
R1212 VN.n54 VN.n53 0.189894
R1213 VN.n53 VN.n52 0.189894
R1214 VN.n13 VN.n12 0.189894
R1215 VN.n14 VN.n13 0.189894
R1216 VN.n14 VN.n7 0.189894
R1217 VN.n18 VN.n7 0.189894
R1218 VN.n19 VN.n18 0.189894
R1219 VN.n20 VN.n19 0.189894
R1220 VN.n20 VN.n5 0.189894
R1221 VN.n25 VN.n5 0.189894
R1222 VN.n26 VN.n25 0.189894
R1223 VN.n27 VN.n26 0.189894
R1224 VN.n27 VN.n3 0.189894
R1225 VN.n31 VN.n3 0.189894
R1226 VN.n32 VN.n31 0.189894
R1227 VN.n33 VN.n32 0.189894
R1228 VN.n33 VN.n1 0.189894
R1229 VN.n37 VN.n1 0.189894
R1230 VTAIL.n11 VTAIL.t3 113.072
R1231 VTAIL.n10 VTAIL.t14 113.072
R1232 VTAIL.n7 VTAIL.t8 113.072
R1233 VTAIL.n15 VTAIL.t13 113.072
R1234 VTAIL.n2 VTAIL.t10 113.072
R1235 VTAIL.n3 VTAIL.t7 113.072
R1236 VTAIL.n6 VTAIL.t1 113.072
R1237 VTAIL.n14 VTAIL.t2 113.072
R1238 VTAIL.n13 VTAIL.n12 103.811
R1239 VTAIL.n9 VTAIL.n8 103.811
R1240 VTAIL.n1 VTAIL.n0 103.811
R1241 VTAIL.n5 VTAIL.n4 103.811
R1242 VTAIL.n15 VTAIL.n14 18.9272
R1243 VTAIL.n7 VTAIL.n6 18.9272
R1244 VTAIL.n0 VTAIL.t15 9.26118
R1245 VTAIL.n0 VTAIL.t9 9.26118
R1246 VTAIL.n4 VTAIL.t6 9.26118
R1247 VTAIL.n4 VTAIL.t4 9.26118
R1248 VTAIL.n12 VTAIL.t0 9.26118
R1249 VTAIL.n12 VTAIL.t5 9.26118
R1250 VTAIL.n8 VTAIL.t12 9.26118
R1251 VTAIL.n8 VTAIL.t11 9.26118
R1252 VTAIL.n9 VTAIL.n7 3.53498
R1253 VTAIL.n10 VTAIL.n9 3.53498
R1254 VTAIL.n13 VTAIL.n11 3.53498
R1255 VTAIL.n14 VTAIL.n13 3.53498
R1256 VTAIL.n6 VTAIL.n5 3.53498
R1257 VTAIL.n5 VTAIL.n3 3.53498
R1258 VTAIL.n2 VTAIL.n1 3.53498
R1259 VTAIL VTAIL.n15 3.47679
R1260 VTAIL.n11 VTAIL.n10 0.470328
R1261 VTAIL.n3 VTAIL.n2 0.470328
R1262 VTAIL VTAIL.n1 0.0586897
R1263 VDD2.n2 VDD2.n1 122.201
R1264 VDD2.n2 VDD2.n0 122.201
R1265 VDD2 VDD2.n5 122.2
R1266 VDD2.n4 VDD2.n3 120.49
R1267 VDD2.n4 VDD2.n2 42.6463
R1268 VDD2.n5 VDD2.t5 9.26118
R1269 VDD2.n5 VDD2.t6 9.26118
R1270 VDD2.n3 VDD2.t1 9.26118
R1271 VDD2.n3 VDD2.t3 9.26118
R1272 VDD2.n1 VDD2.t4 9.26118
R1273 VDD2.n1 VDD2.t7 9.26118
R1274 VDD2.n0 VDD2.t2 9.26118
R1275 VDD2.n0 VDD2.t0 9.26118
R1276 VDD2 VDD2.n4 1.82593
R1277 VP.n25 VP.n24 161.3
R1278 VP.n26 VP.n21 161.3
R1279 VP.n28 VP.n27 161.3
R1280 VP.n29 VP.n20 161.3
R1281 VP.n31 VP.n30 161.3
R1282 VP.n32 VP.n19 161.3
R1283 VP.n34 VP.n33 161.3
R1284 VP.n35 VP.n18 161.3
R1285 VP.n38 VP.n37 161.3
R1286 VP.n39 VP.n17 161.3
R1287 VP.n41 VP.n40 161.3
R1288 VP.n42 VP.n16 161.3
R1289 VP.n44 VP.n43 161.3
R1290 VP.n45 VP.n15 161.3
R1291 VP.n47 VP.n46 161.3
R1292 VP.n48 VP.n14 161.3
R1293 VP.n50 VP.n49 161.3
R1294 VP.n93 VP.n92 161.3
R1295 VP.n91 VP.n1 161.3
R1296 VP.n90 VP.n89 161.3
R1297 VP.n88 VP.n2 161.3
R1298 VP.n87 VP.n86 161.3
R1299 VP.n85 VP.n3 161.3
R1300 VP.n84 VP.n83 161.3
R1301 VP.n82 VP.n4 161.3
R1302 VP.n81 VP.n80 161.3
R1303 VP.n78 VP.n5 161.3
R1304 VP.n77 VP.n76 161.3
R1305 VP.n75 VP.n6 161.3
R1306 VP.n74 VP.n73 161.3
R1307 VP.n72 VP.n7 161.3
R1308 VP.n71 VP.n70 161.3
R1309 VP.n69 VP.n8 161.3
R1310 VP.n68 VP.n67 161.3
R1311 VP.n65 VP.n9 161.3
R1312 VP.n64 VP.n63 161.3
R1313 VP.n62 VP.n10 161.3
R1314 VP.n61 VP.n60 161.3
R1315 VP.n59 VP.n11 161.3
R1316 VP.n58 VP.n57 161.3
R1317 VP.n56 VP.n12 161.3
R1318 VP.n55 VP.n54 161.3
R1319 VP.n53 VP.n52 82.7273
R1320 VP.n94 VP.n0 82.7273
R1321 VP.n51 VP.n13 82.7273
R1322 VP.n23 VP.n22 72.3975
R1323 VP.n22 VP.t3 55.3379
R1324 VP.n60 VP.n59 50.2061
R1325 VP.n86 VP.n2 50.2061
R1326 VP.n43 VP.n15 50.2061
R1327 VP.n52 VP.n51 50.0524
R1328 VP.n73 VP.n72 40.4934
R1329 VP.n73 VP.n6 40.4934
R1330 VP.n30 VP.n19 40.4934
R1331 VP.n30 VP.n29 40.4934
R1332 VP.n60 VP.n10 30.7807
R1333 VP.n86 VP.n85 30.7807
R1334 VP.n43 VP.n42 30.7807
R1335 VP.n54 VP.n12 24.4675
R1336 VP.n58 VP.n12 24.4675
R1337 VP.n59 VP.n58 24.4675
R1338 VP.n64 VP.n10 24.4675
R1339 VP.n65 VP.n64 24.4675
R1340 VP.n67 VP.n8 24.4675
R1341 VP.n71 VP.n8 24.4675
R1342 VP.n72 VP.n71 24.4675
R1343 VP.n77 VP.n6 24.4675
R1344 VP.n78 VP.n77 24.4675
R1345 VP.n80 VP.n78 24.4675
R1346 VP.n84 VP.n4 24.4675
R1347 VP.n85 VP.n84 24.4675
R1348 VP.n90 VP.n2 24.4675
R1349 VP.n91 VP.n90 24.4675
R1350 VP.n92 VP.n91 24.4675
R1351 VP.n47 VP.n15 24.4675
R1352 VP.n48 VP.n47 24.4675
R1353 VP.n49 VP.n48 24.4675
R1354 VP.n34 VP.n19 24.4675
R1355 VP.n35 VP.n34 24.4675
R1356 VP.n37 VP.n35 24.4675
R1357 VP.n41 VP.n17 24.4675
R1358 VP.n42 VP.n41 24.4675
R1359 VP.n24 VP.n21 24.4675
R1360 VP.n28 VP.n21 24.4675
R1361 VP.n29 VP.n28 24.4675
R1362 VP.n53 VP.t7 22.4384
R1363 VP.n66 VP.t5 22.4384
R1364 VP.n79 VP.t0 22.4384
R1365 VP.n0 VP.t1 22.4384
R1366 VP.n13 VP.t2 22.4384
R1367 VP.n36 VP.t4 22.4384
R1368 VP.n23 VP.t6 22.4384
R1369 VP.n66 VP.n65 22.0208
R1370 VP.n79 VP.n4 22.0208
R1371 VP.n36 VP.n17 22.0208
R1372 VP.n54 VP.n53 7.3406
R1373 VP.n92 VP.n0 7.3406
R1374 VP.n49 VP.n13 7.3406
R1375 VP.n25 VP.n22 3.23599
R1376 VP.n67 VP.n66 2.4472
R1377 VP.n80 VP.n79 2.4472
R1378 VP.n37 VP.n36 2.4472
R1379 VP.n24 VP.n23 2.4472
R1380 VP.n51 VP.n50 0.354971
R1381 VP.n55 VP.n52 0.354971
R1382 VP.n94 VP.n93 0.354971
R1383 VP VP.n94 0.26696
R1384 VP.n26 VP.n25 0.189894
R1385 VP.n27 VP.n26 0.189894
R1386 VP.n27 VP.n20 0.189894
R1387 VP.n31 VP.n20 0.189894
R1388 VP.n32 VP.n31 0.189894
R1389 VP.n33 VP.n32 0.189894
R1390 VP.n33 VP.n18 0.189894
R1391 VP.n38 VP.n18 0.189894
R1392 VP.n39 VP.n38 0.189894
R1393 VP.n40 VP.n39 0.189894
R1394 VP.n40 VP.n16 0.189894
R1395 VP.n44 VP.n16 0.189894
R1396 VP.n45 VP.n44 0.189894
R1397 VP.n46 VP.n45 0.189894
R1398 VP.n46 VP.n14 0.189894
R1399 VP.n50 VP.n14 0.189894
R1400 VP.n56 VP.n55 0.189894
R1401 VP.n57 VP.n56 0.189894
R1402 VP.n57 VP.n11 0.189894
R1403 VP.n61 VP.n11 0.189894
R1404 VP.n62 VP.n61 0.189894
R1405 VP.n63 VP.n62 0.189894
R1406 VP.n63 VP.n9 0.189894
R1407 VP.n68 VP.n9 0.189894
R1408 VP.n69 VP.n68 0.189894
R1409 VP.n70 VP.n69 0.189894
R1410 VP.n70 VP.n7 0.189894
R1411 VP.n74 VP.n7 0.189894
R1412 VP.n75 VP.n74 0.189894
R1413 VP.n76 VP.n75 0.189894
R1414 VP.n76 VP.n5 0.189894
R1415 VP.n81 VP.n5 0.189894
R1416 VP.n82 VP.n81 0.189894
R1417 VP.n83 VP.n82 0.189894
R1418 VP.n83 VP.n3 0.189894
R1419 VP.n87 VP.n3 0.189894
R1420 VP.n88 VP.n87 0.189894
R1421 VP.n89 VP.n88 0.189894
R1422 VP.n89 VP.n1 0.189894
R1423 VP.n93 VP.n1 0.189894
R1424 VDD1 VDD1.n0 122.316
R1425 VDD1.n3 VDD1.n2 122.201
R1426 VDD1.n3 VDD1.n1 122.201
R1427 VDD1.n5 VDD1.n4 120.49
R1428 VDD1.n5 VDD1.n3 43.2293
R1429 VDD1.n4 VDD1.t3 9.26118
R1430 VDD1.n4 VDD1.t5 9.26118
R1431 VDD1.n0 VDD1.t4 9.26118
R1432 VDD1.n0 VDD1.t1 9.26118
R1433 VDD1.n2 VDD1.t7 9.26118
R1434 VDD1.n2 VDD1.t6 9.26118
R1435 VDD1.n1 VDD1.t0 9.26118
R1436 VDD1.n1 VDD1.t2 9.26118
R1437 VDD1 VDD1.n5 1.70955
C0 B w_n5070_n1670# 9.5703f
C1 w_n5070_n1670# VP 11.164901f
C2 w_n5070_n1670# VDD1 2.0989f
C3 VTAIL VDD2 6.28492f
C4 B VN 1.4278f
C5 VP VN 7.52585f
C6 B VP 2.54287f
C7 VDD1 VN 0.158346f
C8 B VDD1 1.77782f
C9 w_n5070_n1670# VDD2 2.26227f
C10 VDD1 VP 3.53608f
C11 VDD2 VN 3.04795f
C12 w_n5070_n1670# VTAIL 2.44069f
C13 B VDD2 1.91091f
C14 VP VDD2 0.649499f
C15 VDD1 VDD2 2.38392f
C16 VTAIL VN 4.54447f
C17 B VTAIL 2.45692f
C18 VTAIL VP 4.55857f
C19 VDD1 VTAIL 6.22266f
C20 w_n5070_n1670# VN 10.5048f
C21 VDD2 VSUBS 2.251681f
C22 VDD1 VSUBS 3.10842f
C23 VTAIL VSUBS 0.756688f
C24 VN VSUBS 8.24504f
C25 VP VSUBS 4.140713f
C26 B VSUBS 5.250635f
C27 w_n5070_n1670# VSUBS 0.106896p
C28 VDD1.t4 VSUBS 0.100417f
C29 VDD1.t1 VSUBS 0.100417f
C30 VDD1.n0 VSUBS 0.577681f
C31 VDD1.t0 VSUBS 0.100417f
C32 VDD1.t2 VSUBS 0.100417f
C33 VDD1.n1 VSUBS 0.576469f
C34 VDD1.t7 VSUBS 0.100417f
C35 VDD1.t6 VSUBS 0.100417f
C36 VDD1.n2 VSUBS 0.576469f
C37 VDD1.n3 VSUBS 5.43319f
C38 VDD1.t3 VSUBS 0.100417f
C39 VDD1.t5 VSUBS 0.100417f
C40 VDD1.n4 VSUBS 0.560865f
C41 VDD1.n5 VSUBS 4.14992f
C42 VP.t1 VSUBS 1.51007f
C43 VP.n0 VSUBS 0.776324f
C44 VP.n1 VSUBS 0.044993f
C45 VP.n2 VSUBS 0.082578f
C46 VP.n3 VSUBS 0.044993f
C47 VP.n4 VSUBS 0.079715f
C48 VP.n5 VSUBS 0.044993f
C49 VP.n6 VSUBS 0.089423f
C50 VP.n7 VSUBS 0.044993f
C51 VP.n8 VSUBS 0.083855f
C52 VP.n9 VSUBS 0.044993f
C53 VP.t5 VSUBS 1.51007f
C54 VP.n10 VSUBS 0.090136f
C55 VP.n11 VSUBS 0.044993f
C56 VP.n12 VSUBS 0.083855f
C57 VP.t2 VSUBS 1.51007f
C58 VP.n13 VSUBS 0.776324f
C59 VP.n14 VSUBS 0.044993f
C60 VP.n15 VSUBS 0.082578f
C61 VP.n16 VSUBS 0.044993f
C62 VP.n17 VSUBS 0.079715f
C63 VP.n18 VSUBS 0.044993f
C64 VP.n19 VSUBS 0.089423f
C65 VP.n20 VSUBS 0.044993f
C66 VP.n21 VSUBS 0.083855f
C67 VP.t3 VSUBS 2.0731f
C68 VP.n22 VSUBS 0.759822f
C69 VP.t6 VSUBS 1.51007f
C70 VP.n23 VSUBS 0.742832f
C71 VP.n24 VSUBS 0.046595f
C72 VP.n25 VSUBS 0.572904f
C73 VP.n26 VSUBS 0.044993f
C74 VP.n27 VSUBS 0.044993f
C75 VP.n28 VSUBS 0.083855f
C76 VP.n29 VSUBS 0.089423f
C77 VP.n30 VSUBS 0.036373f
C78 VP.n31 VSUBS 0.044993f
C79 VP.n32 VSUBS 0.044993f
C80 VP.n33 VSUBS 0.044993f
C81 VP.n34 VSUBS 0.083855f
C82 VP.n35 VSUBS 0.083855f
C83 VP.t4 VSUBS 1.51007f
C84 VP.n36 VSUBS 0.597574f
C85 VP.n37 VSUBS 0.046595f
C86 VP.n38 VSUBS 0.044993f
C87 VP.n39 VSUBS 0.044993f
C88 VP.n40 VSUBS 0.044993f
C89 VP.n41 VSUBS 0.083855f
C90 VP.n42 VSUBS 0.090136f
C91 VP.n43 VSUBS 0.042504f
C92 VP.n44 VSUBS 0.044993f
C93 VP.n45 VSUBS 0.044993f
C94 VP.n46 VSUBS 0.044993f
C95 VP.n47 VSUBS 0.083855f
C96 VP.n48 VSUBS 0.083855f
C97 VP.n49 VSUBS 0.054875f
C98 VP.n50 VSUBS 0.072617f
C99 VP.n51 VSUBS 2.58838f
C100 VP.n52 VSUBS 2.62069f
C101 VP.t7 VSUBS 1.51007f
C102 VP.n53 VSUBS 0.776324f
C103 VP.n54 VSUBS 0.054875f
C104 VP.n55 VSUBS 0.072617f
C105 VP.n56 VSUBS 0.044993f
C106 VP.n57 VSUBS 0.044993f
C107 VP.n58 VSUBS 0.083855f
C108 VP.n59 VSUBS 0.082578f
C109 VP.n60 VSUBS 0.042504f
C110 VP.n61 VSUBS 0.044993f
C111 VP.n62 VSUBS 0.044993f
C112 VP.n63 VSUBS 0.044993f
C113 VP.n64 VSUBS 0.083855f
C114 VP.n65 VSUBS 0.079715f
C115 VP.n66 VSUBS 0.597574f
C116 VP.n67 VSUBS 0.046595f
C117 VP.n68 VSUBS 0.044993f
C118 VP.n69 VSUBS 0.044993f
C119 VP.n70 VSUBS 0.044993f
C120 VP.n71 VSUBS 0.083855f
C121 VP.n72 VSUBS 0.089423f
C122 VP.n73 VSUBS 0.036373f
C123 VP.n74 VSUBS 0.044993f
C124 VP.n75 VSUBS 0.044993f
C125 VP.n76 VSUBS 0.044993f
C126 VP.n77 VSUBS 0.083855f
C127 VP.n78 VSUBS 0.083855f
C128 VP.t0 VSUBS 1.51007f
C129 VP.n79 VSUBS 0.597574f
C130 VP.n80 VSUBS 0.046595f
C131 VP.n81 VSUBS 0.044993f
C132 VP.n82 VSUBS 0.044993f
C133 VP.n83 VSUBS 0.044993f
C134 VP.n84 VSUBS 0.083855f
C135 VP.n85 VSUBS 0.090136f
C136 VP.n86 VSUBS 0.042504f
C137 VP.n87 VSUBS 0.044993f
C138 VP.n88 VSUBS 0.044993f
C139 VP.n89 VSUBS 0.044993f
C140 VP.n90 VSUBS 0.083855f
C141 VP.n91 VSUBS 0.083855f
C142 VP.n92 VSUBS 0.054875f
C143 VP.n93 VSUBS 0.072617f
C144 VP.n94 VSUBS 0.131033f
C145 VDD2.t2 VSUBS 0.099944f
C146 VDD2.t0 VSUBS 0.099944f
C147 VDD2.n0 VSUBS 0.573753f
C148 VDD2.t4 VSUBS 0.099944f
C149 VDD2.t7 VSUBS 0.099944f
C150 VDD2.n1 VSUBS 0.573753f
C151 VDD2.n2 VSUBS 5.33314f
C152 VDD2.t1 VSUBS 0.099944f
C153 VDD2.t3 VSUBS 0.099944f
C154 VDD2.n3 VSUBS 0.558225f
C155 VDD2.n4 VSUBS 4.08524f
C156 VDD2.t5 VSUBS 0.099944f
C157 VDD2.t6 VSUBS 0.099944f
C158 VDD2.n5 VSUBS 0.573715f
C159 VTAIL.t15 VSUBS 0.099221f
C160 VTAIL.t9 VSUBS 0.099221f
C161 VTAIL.n0 VSUBS 0.478009f
C162 VTAIL.n1 VSUBS 0.9226f
C163 VTAIL.t10 VSUBS 0.695424f
C164 VTAIL.n2 VSUBS 1.02323f
C165 VTAIL.t7 VSUBS 0.695424f
C166 VTAIL.n3 VSUBS 1.02323f
C167 VTAIL.t6 VSUBS 0.099221f
C168 VTAIL.t4 VSUBS 0.099221f
C169 VTAIL.n4 VSUBS 0.478009f
C170 VTAIL.n5 VSUBS 1.32329f
C171 VTAIL.t1 VSUBS 0.695424f
C172 VTAIL.n6 VSUBS 2.21117f
C173 VTAIL.t8 VSUBS 0.695428f
C174 VTAIL.n7 VSUBS 2.21117f
C175 VTAIL.t12 VSUBS 0.099221f
C176 VTAIL.t11 VSUBS 0.099221f
C177 VTAIL.n8 VSUBS 0.478012f
C178 VTAIL.n9 VSUBS 1.32329f
C179 VTAIL.t14 VSUBS 0.695428f
C180 VTAIL.n10 VSUBS 1.02323f
C181 VTAIL.t3 VSUBS 0.695428f
C182 VTAIL.n11 VSUBS 1.02323f
C183 VTAIL.t0 VSUBS 0.099221f
C184 VTAIL.t5 VSUBS 0.099221f
C185 VTAIL.n12 VSUBS 0.478012f
C186 VTAIL.n13 VSUBS 1.32329f
C187 VTAIL.t2 VSUBS 0.695424f
C188 VTAIL.n14 VSUBS 2.21117f
C189 VTAIL.t13 VSUBS 0.695424f
C190 VTAIL.n15 VSUBS 2.20447f
C191 VN.t0 VSUBS 1.31139f
C192 VN.n0 VSUBS 0.674186f
C193 VN.n1 VSUBS 0.039073f
C194 VN.n2 VSUBS 0.071713f
C195 VN.n3 VSUBS 0.039073f
C196 VN.n4 VSUBS 0.069227f
C197 VN.n5 VSUBS 0.039073f
C198 VN.n6 VSUBS 0.077658f
C199 VN.n7 VSUBS 0.039073f
C200 VN.n8 VSUBS 0.072823f
C201 VN.t5 VSUBS 1.80035f
C202 VN.n9 VSUBS 0.659853f
C203 VN.t7 VSUBS 1.31139f
C204 VN.n10 VSUBS 0.6451f
C205 VN.n11 VSUBS 0.040465f
C206 VN.n12 VSUBS 0.497528f
C207 VN.n13 VSUBS 0.039073f
C208 VN.n14 VSUBS 0.039073f
C209 VN.n15 VSUBS 0.072823f
C210 VN.n16 VSUBS 0.077658f
C211 VN.n17 VSUBS 0.031587f
C212 VN.n18 VSUBS 0.039073f
C213 VN.n19 VSUBS 0.039073f
C214 VN.n20 VSUBS 0.039073f
C215 VN.n21 VSUBS 0.072823f
C216 VN.n22 VSUBS 0.072823f
C217 VN.t3 VSUBS 1.31139f
C218 VN.n23 VSUBS 0.518953f
C219 VN.n24 VSUBS 0.040465f
C220 VN.n25 VSUBS 0.039073f
C221 VN.n26 VSUBS 0.039073f
C222 VN.n27 VSUBS 0.039073f
C223 VN.n28 VSUBS 0.072823f
C224 VN.n29 VSUBS 0.078277f
C225 VN.n30 VSUBS 0.036912f
C226 VN.n31 VSUBS 0.039073f
C227 VN.n32 VSUBS 0.039073f
C228 VN.n33 VSUBS 0.039073f
C229 VN.n34 VSUBS 0.072823f
C230 VN.n35 VSUBS 0.072823f
C231 VN.n36 VSUBS 0.047656f
C232 VN.n37 VSUBS 0.063063f
C233 VN.n38 VSUBS 0.113793f
C234 VN.t6 VSUBS 1.31139f
C235 VN.n39 VSUBS 0.674186f
C236 VN.n40 VSUBS 0.039073f
C237 VN.n41 VSUBS 0.071713f
C238 VN.n42 VSUBS 0.039073f
C239 VN.n43 VSUBS 0.069227f
C240 VN.n44 VSUBS 0.039073f
C241 VN.t4 VSUBS 1.31139f
C242 VN.n45 VSUBS 0.518953f
C243 VN.n46 VSUBS 0.077658f
C244 VN.n47 VSUBS 0.039073f
C245 VN.n48 VSUBS 0.072823f
C246 VN.t1 VSUBS 1.80035f
C247 VN.n49 VSUBS 0.659853f
C248 VN.t2 VSUBS 1.31139f
C249 VN.n50 VSUBS 0.6451f
C250 VN.n51 VSUBS 0.040465f
C251 VN.n52 VSUBS 0.497528f
C252 VN.n53 VSUBS 0.039073f
C253 VN.n54 VSUBS 0.039073f
C254 VN.n55 VSUBS 0.072823f
C255 VN.n56 VSUBS 0.077658f
C256 VN.n57 VSUBS 0.031587f
C257 VN.n58 VSUBS 0.039073f
C258 VN.n59 VSUBS 0.039073f
C259 VN.n60 VSUBS 0.039073f
C260 VN.n61 VSUBS 0.072823f
C261 VN.n62 VSUBS 0.072823f
C262 VN.n63 VSUBS 0.040465f
C263 VN.n64 VSUBS 0.039073f
C264 VN.n65 VSUBS 0.039073f
C265 VN.n66 VSUBS 0.039073f
C266 VN.n67 VSUBS 0.072823f
C267 VN.n68 VSUBS 0.078277f
C268 VN.n69 VSUBS 0.036912f
C269 VN.n70 VSUBS 0.039073f
C270 VN.n71 VSUBS 0.039073f
C271 VN.n72 VSUBS 0.039073f
C272 VN.n73 VSUBS 0.072823f
C273 VN.n74 VSUBS 0.072823f
C274 VN.n75 VSUBS 0.047656f
C275 VN.n76 VSUBS 0.063063f
C276 VN.n77 VSUBS 2.2638f
C277 B.n0 VSUBS 0.009662f
C278 B.n1 VSUBS 0.009662f
C279 B.n2 VSUBS 0.014289f
C280 B.n3 VSUBS 0.01095f
C281 B.n4 VSUBS 0.01095f
C282 B.n5 VSUBS 0.01095f
C283 B.n6 VSUBS 0.01095f
C284 B.n7 VSUBS 0.01095f
C285 B.n8 VSUBS 0.01095f
C286 B.n9 VSUBS 0.01095f
C287 B.n10 VSUBS 0.01095f
C288 B.n11 VSUBS 0.01095f
C289 B.n12 VSUBS 0.01095f
C290 B.n13 VSUBS 0.01095f
C291 B.n14 VSUBS 0.01095f
C292 B.n15 VSUBS 0.01095f
C293 B.n16 VSUBS 0.01095f
C294 B.n17 VSUBS 0.01095f
C295 B.n18 VSUBS 0.01095f
C296 B.n19 VSUBS 0.01095f
C297 B.n20 VSUBS 0.01095f
C298 B.n21 VSUBS 0.01095f
C299 B.n22 VSUBS 0.01095f
C300 B.n23 VSUBS 0.01095f
C301 B.n24 VSUBS 0.01095f
C302 B.n25 VSUBS 0.01095f
C303 B.n26 VSUBS 0.01095f
C304 B.n27 VSUBS 0.01095f
C305 B.n28 VSUBS 0.01095f
C306 B.n29 VSUBS 0.01095f
C307 B.n30 VSUBS 0.01095f
C308 B.n31 VSUBS 0.01095f
C309 B.n32 VSUBS 0.01095f
C310 B.n33 VSUBS 0.01095f
C311 B.n34 VSUBS 0.01095f
C312 B.n35 VSUBS 0.01095f
C313 B.n36 VSUBS 0.025258f
C314 B.n37 VSUBS 0.01095f
C315 B.n38 VSUBS 0.01095f
C316 B.n39 VSUBS 0.01095f
C317 B.n40 VSUBS 0.01095f
C318 B.n41 VSUBS 0.01095f
C319 B.n42 VSUBS 0.01095f
C320 B.n43 VSUBS 0.01095f
C321 B.n44 VSUBS 0.007569f
C322 B.n45 VSUBS 0.01095f
C323 B.t7 VSUBS 0.138844f
C324 B.t8 VSUBS 0.175931f
C325 B.t6 VSUBS 1.01143f
C326 B.n46 VSUBS 0.149635f
C327 B.n47 VSUBS 0.112619f
C328 B.n48 VSUBS 0.02537f
C329 B.n49 VSUBS 0.01095f
C330 B.n50 VSUBS 0.01095f
C331 B.n51 VSUBS 0.01095f
C332 B.n52 VSUBS 0.01095f
C333 B.t4 VSUBS 0.138844f
C334 B.t5 VSUBS 0.17593f
C335 B.t3 VSUBS 1.01143f
C336 B.n53 VSUBS 0.149636f
C337 B.n54 VSUBS 0.112619f
C338 B.n55 VSUBS 0.01095f
C339 B.n56 VSUBS 0.01095f
C340 B.n57 VSUBS 0.01095f
C341 B.n58 VSUBS 0.01095f
C342 B.n59 VSUBS 0.01095f
C343 B.n60 VSUBS 0.01095f
C344 B.n61 VSUBS 0.01095f
C345 B.n62 VSUBS 0.025258f
C346 B.n63 VSUBS 0.01095f
C347 B.n64 VSUBS 0.01095f
C348 B.n65 VSUBS 0.01095f
C349 B.n66 VSUBS 0.01095f
C350 B.n67 VSUBS 0.01095f
C351 B.n68 VSUBS 0.01095f
C352 B.n69 VSUBS 0.01095f
C353 B.n70 VSUBS 0.01095f
C354 B.n71 VSUBS 0.01095f
C355 B.n72 VSUBS 0.01095f
C356 B.n73 VSUBS 0.01095f
C357 B.n74 VSUBS 0.01095f
C358 B.n75 VSUBS 0.01095f
C359 B.n76 VSUBS 0.01095f
C360 B.n77 VSUBS 0.01095f
C361 B.n78 VSUBS 0.01095f
C362 B.n79 VSUBS 0.01095f
C363 B.n80 VSUBS 0.01095f
C364 B.n81 VSUBS 0.01095f
C365 B.n82 VSUBS 0.01095f
C366 B.n83 VSUBS 0.01095f
C367 B.n84 VSUBS 0.01095f
C368 B.n85 VSUBS 0.01095f
C369 B.n86 VSUBS 0.01095f
C370 B.n87 VSUBS 0.01095f
C371 B.n88 VSUBS 0.01095f
C372 B.n89 VSUBS 0.01095f
C373 B.n90 VSUBS 0.01095f
C374 B.n91 VSUBS 0.01095f
C375 B.n92 VSUBS 0.01095f
C376 B.n93 VSUBS 0.01095f
C377 B.n94 VSUBS 0.01095f
C378 B.n95 VSUBS 0.01095f
C379 B.n96 VSUBS 0.01095f
C380 B.n97 VSUBS 0.01095f
C381 B.n98 VSUBS 0.01095f
C382 B.n99 VSUBS 0.01095f
C383 B.n100 VSUBS 0.01095f
C384 B.n101 VSUBS 0.01095f
C385 B.n102 VSUBS 0.01095f
C386 B.n103 VSUBS 0.01095f
C387 B.n104 VSUBS 0.01095f
C388 B.n105 VSUBS 0.01095f
C389 B.n106 VSUBS 0.01095f
C390 B.n107 VSUBS 0.01095f
C391 B.n108 VSUBS 0.01095f
C392 B.n109 VSUBS 0.01095f
C393 B.n110 VSUBS 0.01095f
C394 B.n111 VSUBS 0.01095f
C395 B.n112 VSUBS 0.01095f
C396 B.n113 VSUBS 0.01095f
C397 B.n114 VSUBS 0.01095f
C398 B.n115 VSUBS 0.01095f
C399 B.n116 VSUBS 0.01095f
C400 B.n117 VSUBS 0.01095f
C401 B.n118 VSUBS 0.01095f
C402 B.n119 VSUBS 0.01095f
C403 B.n120 VSUBS 0.01095f
C404 B.n121 VSUBS 0.01095f
C405 B.n122 VSUBS 0.01095f
C406 B.n123 VSUBS 0.01095f
C407 B.n124 VSUBS 0.01095f
C408 B.n125 VSUBS 0.01095f
C409 B.n126 VSUBS 0.01095f
C410 B.n127 VSUBS 0.01095f
C411 B.n128 VSUBS 0.01095f
C412 B.n129 VSUBS 0.01095f
C413 B.n130 VSUBS 0.01095f
C414 B.n131 VSUBS 0.025392f
C415 B.n132 VSUBS 0.01095f
C416 B.n133 VSUBS 0.01095f
C417 B.n134 VSUBS 0.01095f
C418 B.n135 VSUBS 0.01095f
C419 B.n136 VSUBS 0.01095f
C420 B.n137 VSUBS 0.01095f
C421 B.n138 VSUBS 0.01095f
C422 B.n139 VSUBS 0.01095f
C423 B.n140 VSUBS 0.01095f
C424 B.t2 VSUBS 0.138844f
C425 B.t1 VSUBS 0.17593f
C426 B.t0 VSUBS 1.01143f
C427 B.n141 VSUBS 0.149636f
C428 B.n142 VSUBS 0.112619f
C429 B.n143 VSUBS 0.01095f
C430 B.n144 VSUBS 0.01095f
C431 B.n145 VSUBS 0.01095f
C432 B.n146 VSUBS 0.01095f
C433 B.t11 VSUBS 0.138844f
C434 B.t10 VSUBS 0.175931f
C435 B.t9 VSUBS 1.01143f
C436 B.n147 VSUBS 0.149635f
C437 B.n148 VSUBS 0.112619f
C438 B.n149 VSUBS 0.01095f
C439 B.n150 VSUBS 0.01095f
C440 B.n151 VSUBS 0.01095f
C441 B.n152 VSUBS 0.01095f
C442 B.n153 VSUBS 0.01095f
C443 B.n154 VSUBS 0.01095f
C444 B.n155 VSUBS 0.01095f
C445 B.n156 VSUBS 0.01095f
C446 B.n157 VSUBS 0.024018f
C447 B.n158 VSUBS 0.01095f
C448 B.n159 VSUBS 0.01095f
C449 B.n160 VSUBS 0.01095f
C450 B.n161 VSUBS 0.01095f
C451 B.n162 VSUBS 0.01095f
C452 B.n163 VSUBS 0.01095f
C453 B.n164 VSUBS 0.01095f
C454 B.n165 VSUBS 0.01095f
C455 B.n166 VSUBS 0.01095f
C456 B.n167 VSUBS 0.01095f
C457 B.n168 VSUBS 0.01095f
C458 B.n169 VSUBS 0.01095f
C459 B.n170 VSUBS 0.01095f
C460 B.n171 VSUBS 0.01095f
C461 B.n172 VSUBS 0.01095f
C462 B.n173 VSUBS 0.01095f
C463 B.n174 VSUBS 0.01095f
C464 B.n175 VSUBS 0.01095f
C465 B.n176 VSUBS 0.01095f
C466 B.n177 VSUBS 0.01095f
C467 B.n178 VSUBS 0.01095f
C468 B.n179 VSUBS 0.01095f
C469 B.n180 VSUBS 0.01095f
C470 B.n181 VSUBS 0.01095f
C471 B.n182 VSUBS 0.01095f
C472 B.n183 VSUBS 0.01095f
C473 B.n184 VSUBS 0.01095f
C474 B.n185 VSUBS 0.01095f
C475 B.n186 VSUBS 0.01095f
C476 B.n187 VSUBS 0.01095f
C477 B.n188 VSUBS 0.01095f
C478 B.n189 VSUBS 0.01095f
C479 B.n190 VSUBS 0.01095f
C480 B.n191 VSUBS 0.01095f
C481 B.n192 VSUBS 0.01095f
C482 B.n193 VSUBS 0.01095f
C483 B.n194 VSUBS 0.01095f
C484 B.n195 VSUBS 0.01095f
C485 B.n196 VSUBS 0.01095f
C486 B.n197 VSUBS 0.01095f
C487 B.n198 VSUBS 0.01095f
C488 B.n199 VSUBS 0.01095f
C489 B.n200 VSUBS 0.01095f
C490 B.n201 VSUBS 0.01095f
C491 B.n202 VSUBS 0.01095f
C492 B.n203 VSUBS 0.01095f
C493 B.n204 VSUBS 0.01095f
C494 B.n205 VSUBS 0.01095f
C495 B.n206 VSUBS 0.01095f
C496 B.n207 VSUBS 0.01095f
C497 B.n208 VSUBS 0.01095f
C498 B.n209 VSUBS 0.01095f
C499 B.n210 VSUBS 0.01095f
C500 B.n211 VSUBS 0.01095f
C501 B.n212 VSUBS 0.01095f
C502 B.n213 VSUBS 0.01095f
C503 B.n214 VSUBS 0.01095f
C504 B.n215 VSUBS 0.01095f
C505 B.n216 VSUBS 0.01095f
C506 B.n217 VSUBS 0.01095f
C507 B.n218 VSUBS 0.01095f
C508 B.n219 VSUBS 0.01095f
C509 B.n220 VSUBS 0.01095f
C510 B.n221 VSUBS 0.01095f
C511 B.n222 VSUBS 0.01095f
C512 B.n223 VSUBS 0.01095f
C513 B.n224 VSUBS 0.01095f
C514 B.n225 VSUBS 0.01095f
C515 B.n226 VSUBS 0.01095f
C516 B.n227 VSUBS 0.01095f
C517 B.n228 VSUBS 0.01095f
C518 B.n229 VSUBS 0.01095f
C519 B.n230 VSUBS 0.01095f
C520 B.n231 VSUBS 0.01095f
C521 B.n232 VSUBS 0.01095f
C522 B.n233 VSUBS 0.01095f
C523 B.n234 VSUBS 0.01095f
C524 B.n235 VSUBS 0.01095f
C525 B.n236 VSUBS 0.01095f
C526 B.n237 VSUBS 0.01095f
C527 B.n238 VSUBS 0.01095f
C528 B.n239 VSUBS 0.01095f
C529 B.n240 VSUBS 0.01095f
C530 B.n241 VSUBS 0.01095f
C531 B.n242 VSUBS 0.01095f
C532 B.n243 VSUBS 0.01095f
C533 B.n244 VSUBS 0.01095f
C534 B.n245 VSUBS 0.01095f
C535 B.n246 VSUBS 0.01095f
C536 B.n247 VSUBS 0.01095f
C537 B.n248 VSUBS 0.01095f
C538 B.n249 VSUBS 0.01095f
C539 B.n250 VSUBS 0.01095f
C540 B.n251 VSUBS 0.01095f
C541 B.n252 VSUBS 0.01095f
C542 B.n253 VSUBS 0.01095f
C543 B.n254 VSUBS 0.01095f
C544 B.n255 VSUBS 0.01095f
C545 B.n256 VSUBS 0.01095f
C546 B.n257 VSUBS 0.01095f
C547 B.n258 VSUBS 0.01095f
C548 B.n259 VSUBS 0.01095f
C549 B.n260 VSUBS 0.01095f
C550 B.n261 VSUBS 0.01095f
C551 B.n262 VSUBS 0.01095f
C552 B.n263 VSUBS 0.01095f
C553 B.n264 VSUBS 0.01095f
C554 B.n265 VSUBS 0.01095f
C555 B.n266 VSUBS 0.01095f
C556 B.n267 VSUBS 0.01095f
C557 B.n268 VSUBS 0.01095f
C558 B.n269 VSUBS 0.01095f
C559 B.n270 VSUBS 0.01095f
C560 B.n271 VSUBS 0.01095f
C561 B.n272 VSUBS 0.01095f
C562 B.n273 VSUBS 0.01095f
C563 B.n274 VSUBS 0.01095f
C564 B.n275 VSUBS 0.01095f
C565 B.n276 VSUBS 0.01095f
C566 B.n277 VSUBS 0.01095f
C567 B.n278 VSUBS 0.01095f
C568 B.n279 VSUBS 0.01095f
C569 B.n280 VSUBS 0.01095f
C570 B.n281 VSUBS 0.01095f
C571 B.n282 VSUBS 0.01095f
C572 B.n283 VSUBS 0.01095f
C573 B.n284 VSUBS 0.01095f
C574 B.n285 VSUBS 0.01095f
C575 B.n286 VSUBS 0.01095f
C576 B.n287 VSUBS 0.01095f
C577 B.n288 VSUBS 0.01095f
C578 B.n289 VSUBS 0.01095f
C579 B.n290 VSUBS 0.024018f
C580 B.n291 VSUBS 0.025258f
C581 B.n292 VSUBS 0.025258f
C582 B.n293 VSUBS 0.01095f
C583 B.n294 VSUBS 0.01095f
C584 B.n295 VSUBS 0.01095f
C585 B.n296 VSUBS 0.01095f
C586 B.n297 VSUBS 0.01095f
C587 B.n298 VSUBS 0.01095f
C588 B.n299 VSUBS 0.01095f
C589 B.n300 VSUBS 0.01095f
C590 B.n301 VSUBS 0.01095f
C591 B.n302 VSUBS 0.01095f
C592 B.n303 VSUBS 0.01095f
C593 B.n304 VSUBS 0.01095f
C594 B.n305 VSUBS 0.01095f
C595 B.n306 VSUBS 0.01095f
C596 B.n307 VSUBS 0.01095f
C597 B.n308 VSUBS 0.01095f
C598 B.n309 VSUBS 0.01095f
C599 B.n310 VSUBS 0.01095f
C600 B.n311 VSUBS 0.01095f
C601 B.n312 VSUBS 0.01095f
C602 B.n313 VSUBS 0.01095f
C603 B.n314 VSUBS 0.01095f
C604 B.n315 VSUBS 0.01095f
C605 B.n316 VSUBS 0.007569f
C606 B.n317 VSUBS 0.02537f
C607 B.n318 VSUBS 0.008857f
C608 B.n319 VSUBS 0.01095f
C609 B.n320 VSUBS 0.01095f
C610 B.n321 VSUBS 0.01095f
C611 B.n322 VSUBS 0.01095f
C612 B.n323 VSUBS 0.01095f
C613 B.n324 VSUBS 0.01095f
C614 B.n325 VSUBS 0.01095f
C615 B.n326 VSUBS 0.01095f
C616 B.n327 VSUBS 0.01095f
C617 B.n328 VSUBS 0.01095f
C618 B.n329 VSUBS 0.01095f
C619 B.n330 VSUBS 0.008857f
C620 B.n331 VSUBS 0.02537f
C621 B.n332 VSUBS 0.007569f
C622 B.n333 VSUBS 0.01095f
C623 B.n334 VSUBS 0.01095f
C624 B.n335 VSUBS 0.01095f
C625 B.n336 VSUBS 0.01095f
C626 B.n337 VSUBS 0.01095f
C627 B.n338 VSUBS 0.01095f
C628 B.n339 VSUBS 0.01095f
C629 B.n340 VSUBS 0.01095f
C630 B.n341 VSUBS 0.01095f
C631 B.n342 VSUBS 0.01095f
C632 B.n343 VSUBS 0.01095f
C633 B.n344 VSUBS 0.01095f
C634 B.n345 VSUBS 0.01095f
C635 B.n346 VSUBS 0.01095f
C636 B.n347 VSUBS 0.01095f
C637 B.n348 VSUBS 0.01095f
C638 B.n349 VSUBS 0.01095f
C639 B.n350 VSUBS 0.01095f
C640 B.n351 VSUBS 0.01095f
C641 B.n352 VSUBS 0.01095f
C642 B.n353 VSUBS 0.01095f
C643 B.n354 VSUBS 0.01095f
C644 B.n355 VSUBS 0.01095f
C645 B.n356 VSUBS 0.023884f
C646 B.n357 VSUBS 0.025258f
C647 B.n358 VSUBS 0.024018f
C648 B.n359 VSUBS 0.01095f
C649 B.n360 VSUBS 0.01095f
C650 B.n361 VSUBS 0.01095f
C651 B.n362 VSUBS 0.01095f
C652 B.n363 VSUBS 0.01095f
C653 B.n364 VSUBS 0.01095f
C654 B.n365 VSUBS 0.01095f
C655 B.n366 VSUBS 0.01095f
C656 B.n367 VSUBS 0.01095f
C657 B.n368 VSUBS 0.01095f
C658 B.n369 VSUBS 0.01095f
C659 B.n370 VSUBS 0.01095f
C660 B.n371 VSUBS 0.01095f
C661 B.n372 VSUBS 0.01095f
C662 B.n373 VSUBS 0.01095f
C663 B.n374 VSUBS 0.01095f
C664 B.n375 VSUBS 0.01095f
C665 B.n376 VSUBS 0.01095f
C666 B.n377 VSUBS 0.01095f
C667 B.n378 VSUBS 0.01095f
C668 B.n379 VSUBS 0.01095f
C669 B.n380 VSUBS 0.01095f
C670 B.n381 VSUBS 0.01095f
C671 B.n382 VSUBS 0.01095f
C672 B.n383 VSUBS 0.01095f
C673 B.n384 VSUBS 0.01095f
C674 B.n385 VSUBS 0.01095f
C675 B.n386 VSUBS 0.01095f
C676 B.n387 VSUBS 0.01095f
C677 B.n388 VSUBS 0.01095f
C678 B.n389 VSUBS 0.01095f
C679 B.n390 VSUBS 0.01095f
C680 B.n391 VSUBS 0.01095f
C681 B.n392 VSUBS 0.01095f
C682 B.n393 VSUBS 0.01095f
C683 B.n394 VSUBS 0.01095f
C684 B.n395 VSUBS 0.01095f
C685 B.n396 VSUBS 0.01095f
C686 B.n397 VSUBS 0.01095f
C687 B.n398 VSUBS 0.01095f
C688 B.n399 VSUBS 0.01095f
C689 B.n400 VSUBS 0.01095f
C690 B.n401 VSUBS 0.01095f
C691 B.n402 VSUBS 0.01095f
C692 B.n403 VSUBS 0.01095f
C693 B.n404 VSUBS 0.01095f
C694 B.n405 VSUBS 0.01095f
C695 B.n406 VSUBS 0.01095f
C696 B.n407 VSUBS 0.01095f
C697 B.n408 VSUBS 0.01095f
C698 B.n409 VSUBS 0.01095f
C699 B.n410 VSUBS 0.01095f
C700 B.n411 VSUBS 0.01095f
C701 B.n412 VSUBS 0.01095f
C702 B.n413 VSUBS 0.01095f
C703 B.n414 VSUBS 0.01095f
C704 B.n415 VSUBS 0.01095f
C705 B.n416 VSUBS 0.01095f
C706 B.n417 VSUBS 0.01095f
C707 B.n418 VSUBS 0.01095f
C708 B.n419 VSUBS 0.01095f
C709 B.n420 VSUBS 0.01095f
C710 B.n421 VSUBS 0.01095f
C711 B.n422 VSUBS 0.01095f
C712 B.n423 VSUBS 0.01095f
C713 B.n424 VSUBS 0.01095f
C714 B.n425 VSUBS 0.01095f
C715 B.n426 VSUBS 0.01095f
C716 B.n427 VSUBS 0.01095f
C717 B.n428 VSUBS 0.01095f
C718 B.n429 VSUBS 0.01095f
C719 B.n430 VSUBS 0.01095f
C720 B.n431 VSUBS 0.01095f
C721 B.n432 VSUBS 0.01095f
C722 B.n433 VSUBS 0.01095f
C723 B.n434 VSUBS 0.01095f
C724 B.n435 VSUBS 0.01095f
C725 B.n436 VSUBS 0.01095f
C726 B.n437 VSUBS 0.01095f
C727 B.n438 VSUBS 0.01095f
C728 B.n439 VSUBS 0.01095f
C729 B.n440 VSUBS 0.01095f
C730 B.n441 VSUBS 0.01095f
C731 B.n442 VSUBS 0.01095f
C732 B.n443 VSUBS 0.01095f
C733 B.n444 VSUBS 0.01095f
C734 B.n445 VSUBS 0.01095f
C735 B.n446 VSUBS 0.01095f
C736 B.n447 VSUBS 0.01095f
C737 B.n448 VSUBS 0.01095f
C738 B.n449 VSUBS 0.01095f
C739 B.n450 VSUBS 0.01095f
C740 B.n451 VSUBS 0.01095f
C741 B.n452 VSUBS 0.01095f
C742 B.n453 VSUBS 0.01095f
C743 B.n454 VSUBS 0.01095f
C744 B.n455 VSUBS 0.01095f
C745 B.n456 VSUBS 0.01095f
C746 B.n457 VSUBS 0.01095f
C747 B.n458 VSUBS 0.01095f
C748 B.n459 VSUBS 0.01095f
C749 B.n460 VSUBS 0.01095f
C750 B.n461 VSUBS 0.01095f
C751 B.n462 VSUBS 0.01095f
C752 B.n463 VSUBS 0.01095f
C753 B.n464 VSUBS 0.01095f
C754 B.n465 VSUBS 0.01095f
C755 B.n466 VSUBS 0.01095f
C756 B.n467 VSUBS 0.01095f
C757 B.n468 VSUBS 0.01095f
C758 B.n469 VSUBS 0.01095f
C759 B.n470 VSUBS 0.01095f
C760 B.n471 VSUBS 0.01095f
C761 B.n472 VSUBS 0.01095f
C762 B.n473 VSUBS 0.01095f
C763 B.n474 VSUBS 0.01095f
C764 B.n475 VSUBS 0.01095f
C765 B.n476 VSUBS 0.01095f
C766 B.n477 VSUBS 0.01095f
C767 B.n478 VSUBS 0.01095f
C768 B.n479 VSUBS 0.01095f
C769 B.n480 VSUBS 0.01095f
C770 B.n481 VSUBS 0.01095f
C771 B.n482 VSUBS 0.01095f
C772 B.n483 VSUBS 0.01095f
C773 B.n484 VSUBS 0.01095f
C774 B.n485 VSUBS 0.01095f
C775 B.n486 VSUBS 0.01095f
C776 B.n487 VSUBS 0.01095f
C777 B.n488 VSUBS 0.01095f
C778 B.n489 VSUBS 0.01095f
C779 B.n490 VSUBS 0.01095f
C780 B.n491 VSUBS 0.01095f
C781 B.n492 VSUBS 0.01095f
C782 B.n493 VSUBS 0.01095f
C783 B.n494 VSUBS 0.01095f
C784 B.n495 VSUBS 0.01095f
C785 B.n496 VSUBS 0.01095f
C786 B.n497 VSUBS 0.01095f
C787 B.n498 VSUBS 0.01095f
C788 B.n499 VSUBS 0.01095f
C789 B.n500 VSUBS 0.01095f
C790 B.n501 VSUBS 0.01095f
C791 B.n502 VSUBS 0.01095f
C792 B.n503 VSUBS 0.01095f
C793 B.n504 VSUBS 0.01095f
C794 B.n505 VSUBS 0.01095f
C795 B.n506 VSUBS 0.01095f
C796 B.n507 VSUBS 0.01095f
C797 B.n508 VSUBS 0.01095f
C798 B.n509 VSUBS 0.01095f
C799 B.n510 VSUBS 0.01095f
C800 B.n511 VSUBS 0.01095f
C801 B.n512 VSUBS 0.01095f
C802 B.n513 VSUBS 0.01095f
C803 B.n514 VSUBS 0.01095f
C804 B.n515 VSUBS 0.01095f
C805 B.n516 VSUBS 0.01095f
C806 B.n517 VSUBS 0.01095f
C807 B.n518 VSUBS 0.01095f
C808 B.n519 VSUBS 0.01095f
C809 B.n520 VSUBS 0.01095f
C810 B.n521 VSUBS 0.01095f
C811 B.n522 VSUBS 0.01095f
C812 B.n523 VSUBS 0.01095f
C813 B.n524 VSUBS 0.01095f
C814 B.n525 VSUBS 0.01095f
C815 B.n526 VSUBS 0.01095f
C816 B.n527 VSUBS 0.01095f
C817 B.n528 VSUBS 0.01095f
C818 B.n529 VSUBS 0.01095f
C819 B.n530 VSUBS 0.01095f
C820 B.n531 VSUBS 0.01095f
C821 B.n532 VSUBS 0.01095f
C822 B.n533 VSUBS 0.01095f
C823 B.n534 VSUBS 0.01095f
C824 B.n535 VSUBS 0.01095f
C825 B.n536 VSUBS 0.01095f
C826 B.n537 VSUBS 0.01095f
C827 B.n538 VSUBS 0.01095f
C828 B.n539 VSUBS 0.01095f
C829 B.n540 VSUBS 0.01095f
C830 B.n541 VSUBS 0.01095f
C831 B.n542 VSUBS 0.01095f
C832 B.n543 VSUBS 0.01095f
C833 B.n544 VSUBS 0.01095f
C834 B.n545 VSUBS 0.01095f
C835 B.n546 VSUBS 0.01095f
C836 B.n547 VSUBS 0.01095f
C837 B.n548 VSUBS 0.01095f
C838 B.n549 VSUBS 0.01095f
C839 B.n550 VSUBS 0.01095f
C840 B.n551 VSUBS 0.01095f
C841 B.n552 VSUBS 0.01095f
C842 B.n553 VSUBS 0.01095f
C843 B.n554 VSUBS 0.01095f
C844 B.n555 VSUBS 0.01095f
C845 B.n556 VSUBS 0.01095f
C846 B.n557 VSUBS 0.01095f
C847 B.n558 VSUBS 0.01095f
C848 B.n559 VSUBS 0.01095f
C849 B.n560 VSUBS 0.01095f
C850 B.n561 VSUBS 0.01095f
C851 B.n562 VSUBS 0.01095f
C852 B.n563 VSUBS 0.024018f
C853 B.n564 VSUBS 0.024018f
C854 B.n565 VSUBS 0.025258f
C855 B.n566 VSUBS 0.01095f
C856 B.n567 VSUBS 0.01095f
C857 B.n568 VSUBS 0.01095f
C858 B.n569 VSUBS 0.01095f
C859 B.n570 VSUBS 0.01095f
C860 B.n571 VSUBS 0.01095f
C861 B.n572 VSUBS 0.01095f
C862 B.n573 VSUBS 0.01095f
C863 B.n574 VSUBS 0.01095f
C864 B.n575 VSUBS 0.01095f
C865 B.n576 VSUBS 0.01095f
C866 B.n577 VSUBS 0.01095f
C867 B.n578 VSUBS 0.01095f
C868 B.n579 VSUBS 0.01095f
C869 B.n580 VSUBS 0.01095f
C870 B.n581 VSUBS 0.01095f
C871 B.n582 VSUBS 0.01095f
C872 B.n583 VSUBS 0.01095f
C873 B.n584 VSUBS 0.01095f
C874 B.n585 VSUBS 0.01095f
C875 B.n586 VSUBS 0.01095f
C876 B.n587 VSUBS 0.01095f
C877 B.n588 VSUBS 0.01095f
C878 B.n589 VSUBS 0.007569f
C879 B.n590 VSUBS 0.02537f
C880 B.n591 VSUBS 0.008857f
C881 B.n592 VSUBS 0.01095f
C882 B.n593 VSUBS 0.01095f
C883 B.n594 VSUBS 0.01095f
C884 B.n595 VSUBS 0.01095f
C885 B.n596 VSUBS 0.01095f
C886 B.n597 VSUBS 0.01095f
C887 B.n598 VSUBS 0.01095f
C888 B.n599 VSUBS 0.01095f
C889 B.n600 VSUBS 0.01095f
C890 B.n601 VSUBS 0.01095f
C891 B.n602 VSUBS 0.01095f
C892 B.n603 VSUBS 0.008857f
C893 B.n604 VSUBS 0.01095f
C894 B.n605 VSUBS 0.01095f
C895 B.n606 VSUBS 0.01095f
C896 B.n607 VSUBS 0.01095f
C897 B.n608 VSUBS 0.01095f
C898 B.n609 VSUBS 0.01095f
C899 B.n610 VSUBS 0.01095f
C900 B.n611 VSUBS 0.01095f
C901 B.n612 VSUBS 0.01095f
C902 B.n613 VSUBS 0.01095f
C903 B.n614 VSUBS 0.01095f
C904 B.n615 VSUBS 0.01095f
C905 B.n616 VSUBS 0.01095f
C906 B.n617 VSUBS 0.01095f
C907 B.n618 VSUBS 0.01095f
C908 B.n619 VSUBS 0.01095f
C909 B.n620 VSUBS 0.01095f
C910 B.n621 VSUBS 0.01095f
C911 B.n622 VSUBS 0.01095f
C912 B.n623 VSUBS 0.01095f
C913 B.n624 VSUBS 0.01095f
C914 B.n625 VSUBS 0.01095f
C915 B.n626 VSUBS 0.01095f
C916 B.n627 VSUBS 0.01095f
C917 B.n628 VSUBS 0.01095f
C918 B.n629 VSUBS 0.025258f
C919 B.n630 VSUBS 0.024018f
C920 B.n631 VSUBS 0.024018f
C921 B.n632 VSUBS 0.01095f
C922 B.n633 VSUBS 0.01095f
C923 B.n634 VSUBS 0.01095f
C924 B.n635 VSUBS 0.01095f
C925 B.n636 VSUBS 0.01095f
C926 B.n637 VSUBS 0.01095f
C927 B.n638 VSUBS 0.01095f
C928 B.n639 VSUBS 0.01095f
C929 B.n640 VSUBS 0.01095f
C930 B.n641 VSUBS 0.01095f
C931 B.n642 VSUBS 0.01095f
C932 B.n643 VSUBS 0.01095f
C933 B.n644 VSUBS 0.01095f
C934 B.n645 VSUBS 0.01095f
C935 B.n646 VSUBS 0.01095f
C936 B.n647 VSUBS 0.01095f
C937 B.n648 VSUBS 0.01095f
C938 B.n649 VSUBS 0.01095f
C939 B.n650 VSUBS 0.01095f
C940 B.n651 VSUBS 0.01095f
C941 B.n652 VSUBS 0.01095f
C942 B.n653 VSUBS 0.01095f
C943 B.n654 VSUBS 0.01095f
C944 B.n655 VSUBS 0.01095f
C945 B.n656 VSUBS 0.01095f
C946 B.n657 VSUBS 0.01095f
C947 B.n658 VSUBS 0.01095f
C948 B.n659 VSUBS 0.01095f
C949 B.n660 VSUBS 0.01095f
C950 B.n661 VSUBS 0.01095f
C951 B.n662 VSUBS 0.01095f
C952 B.n663 VSUBS 0.01095f
C953 B.n664 VSUBS 0.01095f
C954 B.n665 VSUBS 0.01095f
C955 B.n666 VSUBS 0.01095f
C956 B.n667 VSUBS 0.01095f
C957 B.n668 VSUBS 0.01095f
C958 B.n669 VSUBS 0.01095f
C959 B.n670 VSUBS 0.01095f
C960 B.n671 VSUBS 0.01095f
C961 B.n672 VSUBS 0.01095f
C962 B.n673 VSUBS 0.01095f
C963 B.n674 VSUBS 0.01095f
C964 B.n675 VSUBS 0.01095f
C965 B.n676 VSUBS 0.01095f
C966 B.n677 VSUBS 0.01095f
C967 B.n678 VSUBS 0.01095f
C968 B.n679 VSUBS 0.01095f
C969 B.n680 VSUBS 0.01095f
C970 B.n681 VSUBS 0.01095f
C971 B.n682 VSUBS 0.01095f
C972 B.n683 VSUBS 0.01095f
C973 B.n684 VSUBS 0.01095f
C974 B.n685 VSUBS 0.01095f
C975 B.n686 VSUBS 0.01095f
C976 B.n687 VSUBS 0.01095f
C977 B.n688 VSUBS 0.01095f
C978 B.n689 VSUBS 0.01095f
C979 B.n690 VSUBS 0.01095f
C980 B.n691 VSUBS 0.01095f
C981 B.n692 VSUBS 0.01095f
C982 B.n693 VSUBS 0.01095f
C983 B.n694 VSUBS 0.01095f
C984 B.n695 VSUBS 0.01095f
C985 B.n696 VSUBS 0.01095f
C986 B.n697 VSUBS 0.01095f
C987 B.n698 VSUBS 0.01095f
C988 B.n699 VSUBS 0.01095f
C989 B.n700 VSUBS 0.01095f
C990 B.n701 VSUBS 0.01095f
C991 B.n702 VSUBS 0.01095f
C992 B.n703 VSUBS 0.01095f
C993 B.n704 VSUBS 0.01095f
C994 B.n705 VSUBS 0.01095f
C995 B.n706 VSUBS 0.01095f
C996 B.n707 VSUBS 0.01095f
C997 B.n708 VSUBS 0.01095f
C998 B.n709 VSUBS 0.01095f
C999 B.n710 VSUBS 0.01095f
C1000 B.n711 VSUBS 0.01095f
C1001 B.n712 VSUBS 0.01095f
C1002 B.n713 VSUBS 0.01095f
C1003 B.n714 VSUBS 0.01095f
C1004 B.n715 VSUBS 0.01095f
C1005 B.n716 VSUBS 0.01095f
C1006 B.n717 VSUBS 0.01095f
C1007 B.n718 VSUBS 0.01095f
C1008 B.n719 VSUBS 0.01095f
C1009 B.n720 VSUBS 0.01095f
C1010 B.n721 VSUBS 0.01095f
C1011 B.n722 VSUBS 0.01095f
C1012 B.n723 VSUBS 0.01095f
C1013 B.n724 VSUBS 0.01095f
C1014 B.n725 VSUBS 0.01095f
C1015 B.n726 VSUBS 0.01095f
C1016 B.n727 VSUBS 0.01095f
C1017 B.n728 VSUBS 0.01095f
C1018 B.n729 VSUBS 0.01095f
C1019 B.n730 VSUBS 0.01095f
C1020 B.n731 VSUBS 0.014289f
C1021 B.n732 VSUBS 0.015222f
C1022 B.n733 VSUBS 0.03027f
.ends

