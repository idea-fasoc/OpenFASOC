* NGSPICE file created from diff_pair_sample_0408.ext - technology: sky130A

.subckt diff_pair_sample_0408 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0 ps=0 w=0.83 l=1.56
X1 B.t8 B.t6 B.t7 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0 ps=0 w=0.83 l=1.56
X2 VTAIL.t7 VP.t0 VDD1.t0 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0.13695 ps=1.16 w=0.83 l=1.56
X3 B.t5 B.t3 B.t4 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0 ps=0 w=0.83 l=1.56
X4 VTAIL.t1 VN.t0 VDD2.t3 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0.13695 ps=1.16 w=0.83 l=1.56
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.13695 pd=1.16 as=0.3237 ps=2.44 w=0.83 l=1.56
X6 VDD1.t2 VP.t1 VTAIL.t6 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.13695 pd=1.16 as=0.3237 ps=2.44 w=0.83 l=1.56
X7 VTAIL.t5 VP.t2 VDD1.t3 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0.13695 ps=1.16 w=0.83 l=1.56
X8 VTAIL.t2 VN.t2 VDD2.t1 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0.13695 ps=1.16 w=0.83 l=1.56
X9 VDD2.t0 VN.t3 VTAIL.t3 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.13695 pd=1.16 as=0.3237 ps=2.44 w=0.83 l=1.56
X10 VDD1.t1 VP.t3 VTAIL.t4 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.13695 pd=1.16 as=0.3237 ps=2.44 w=0.83 l=1.56
X11 B.t2 B.t0 B.t1 w_n2104_n1134# sky130_fd_pr__pfet_01v8 ad=0.3237 pd=2.44 as=0 ps=0 w=0.83 l=1.56
R0 B.n69 B.t1 686.611
R1 B.n63 B.t7 686.611
R2 B.n27 B.t5 686.611
R3 B.n20 B.t11 686.611
R4 B.n70 B.t2 649.957
R5 B.n64 B.t8 649.957
R6 B.n28 B.t4 649.957
R7 B.n21 B.t10 649.957
R8 B.n163 B.n162 585
R9 B.n161 B.n58 585
R10 B.n160 B.n159 585
R11 B.n158 B.n59 585
R12 B.n157 B.n156 585
R13 B.n155 B.n60 585
R14 B.n154 B.n153 585
R15 B.n152 B.n61 585
R16 B.n151 B.n150 585
R17 B.n148 B.n62 585
R18 B.n147 B.n146 585
R19 B.n145 B.n65 585
R20 B.n144 B.n143 585
R21 B.n142 B.n66 585
R22 B.n141 B.n140 585
R23 B.n139 B.n67 585
R24 B.n138 B.n137 585
R25 B.n136 B.n68 585
R26 B.n134 B.n133 585
R27 B.n132 B.n71 585
R28 B.n131 B.n130 585
R29 B.n129 B.n72 585
R30 B.n128 B.n127 585
R31 B.n126 B.n73 585
R32 B.n125 B.n124 585
R33 B.n123 B.n74 585
R34 B.n122 B.n121 585
R35 B.n164 B.n57 585
R36 B.n166 B.n165 585
R37 B.n167 B.n56 585
R38 B.n169 B.n168 585
R39 B.n170 B.n55 585
R40 B.n172 B.n171 585
R41 B.n173 B.n54 585
R42 B.n175 B.n174 585
R43 B.n176 B.n53 585
R44 B.n178 B.n177 585
R45 B.n179 B.n52 585
R46 B.n181 B.n180 585
R47 B.n182 B.n51 585
R48 B.n184 B.n183 585
R49 B.n185 B.n50 585
R50 B.n187 B.n186 585
R51 B.n188 B.n49 585
R52 B.n190 B.n189 585
R53 B.n191 B.n48 585
R54 B.n193 B.n192 585
R55 B.n194 B.n47 585
R56 B.n196 B.n195 585
R57 B.n197 B.n46 585
R58 B.n199 B.n198 585
R59 B.n200 B.n45 585
R60 B.n202 B.n201 585
R61 B.n203 B.n44 585
R62 B.n205 B.n204 585
R63 B.n206 B.n43 585
R64 B.n208 B.n207 585
R65 B.n209 B.n42 585
R66 B.n211 B.n210 585
R67 B.n212 B.n41 585
R68 B.n214 B.n213 585
R69 B.n215 B.n40 585
R70 B.n217 B.n216 585
R71 B.n218 B.n39 585
R72 B.n220 B.n219 585
R73 B.n221 B.n38 585
R74 B.n223 B.n222 585
R75 B.n224 B.n37 585
R76 B.n226 B.n225 585
R77 B.n227 B.n36 585
R78 B.n229 B.n228 585
R79 B.n230 B.n35 585
R80 B.n232 B.n231 585
R81 B.n233 B.n34 585
R82 B.n235 B.n234 585
R83 B.n236 B.n33 585
R84 B.n238 B.n237 585
R85 B.n279 B.n14 585
R86 B.n278 B.n277 585
R87 B.n276 B.n15 585
R88 B.n275 B.n274 585
R89 B.n273 B.n16 585
R90 B.n272 B.n271 585
R91 B.n270 B.n17 585
R92 B.n269 B.n268 585
R93 B.n267 B.n18 585
R94 B.n266 B.n265 585
R95 B.n264 B.n19 585
R96 B.n263 B.n262 585
R97 B.n261 B.n23 585
R98 B.n260 B.n259 585
R99 B.n258 B.n24 585
R100 B.n257 B.n256 585
R101 B.n255 B.n25 585
R102 B.n254 B.n253 585
R103 B.n251 B.n26 585
R104 B.n250 B.n249 585
R105 B.n248 B.n29 585
R106 B.n247 B.n246 585
R107 B.n245 B.n30 585
R108 B.n244 B.n243 585
R109 B.n242 B.n31 585
R110 B.n241 B.n240 585
R111 B.n239 B.n32 585
R112 B.n281 B.n280 585
R113 B.n282 B.n13 585
R114 B.n284 B.n283 585
R115 B.n285 B.n12 585
R116 B.n287 B.n286 585
R117 B.n288 B.n11 585
R118 B.n290 B.n289 585
R119 B.n291 B.n10 585
R120 B.n293 B.n292 585
R121 B.n294 B.n9 585
R122 B.n296 B.n295 585
R123 B.n297 B.n8 585
R124 B.n299 B.n298 585
R125 B.n300 B.n7 585
R126 B.n302 B.n301 585
R127 B.n303 B.n6 585
R128 B.n305 B.n304 585
R129 B.n306 B.n5 585
R130 B.n308 B.n307 585
R131 B.n309 B.n4 585
R132 B.n311 B.n310 585
R133 B.n312 B.n3 585
R134 B.n314 B.n313 585
R135 B.n315 B.n0 585
R136 B.n2 B.n1 585
R137 B.n87 B.n86 585
R138 B.n89 B.n88 585
R139 B.n90 B.n85 585
R140 B.n92 B.n91 585
R141 B.n93 B.n84 585
R142 B.n95 B.n94 585
R143 B.n96 B.n83 585
R144 B.n98 B.n97 585
R145 B.n99 B.n82 585
R146 B.n101 B.n100 585
R147 B.n102 B.n81 585
R148 B.n104 B.n103 585
R149 B.n105 B.n80 585
R150 B.n107 B.n106 585
R151 B.n108 B.n79 585
R152 B.n110 B.n109 585
R153 B.n111 B.n78 585
R154 B.n113 B.n112 585
R155 B.n114 B.n77 585
R156 B.n116 B.n115 585
R157 B.n117 B.n76 585
R158 B.n119 B.n118 585
R159 B.n120 B.n75 585
R160 B.n121 B.n120 554.963
R161 B.n164 B.n163 554.963
R162 B.n237 B.n32 554.963
R163 B.n280 B.n279 554.963
R164 B.n317 B.n316 256.663
R165 B.n316 B.n315 235.042
R166 B.n316 B.n2 235.042
R167 B.n69 B.t0 207.206
R168 B.n63 B.t6 207.206
R169 B.n27 B.t3 207.206
R170 B.n20 B.t9 207.206
R171 B.n121 B.n74 163.367
R172 B.n125 B.n74 163.367
R173 B.n126 B.n125 163.367
R174 B.n127 B.n126 163.367
R175 B.n127 B.n72 163.367
R176 B.n131 B.n72 163.367
R177 B.n132 B.n131 163.367
R178 B.n133 B.n132 163.367
R179 B.n133 B.n68 163.367
R180 B.n138 B.n68 163.367
R181 B.n139 B.n138 163.367
R182 B.n140 B.n139 163.367
R183 B.n140 B.n66 163.367
R184 B.n144 B.n66 163.367
R185 B.n145 B.n144 163.367
R186 B.n146 B.n145 163.367
R187 B.n146 B.n62 163.367
R188 B.n151 B.n62 163.367
R189 B.n152 B.n151 163.367
R190 B.n153 B.n152 163.367
R191 B.n153 B.n60 163.367
R192 B.n157 B.n60 163.367
R193 B.n158 B.n157 163.367
R194 B.n159 B.n158 163.367
R195 B.n159 B.n58 163.367
R196 B.n163 B.n58 163.367
R197 B.n237 B.n236 163.367
R198 B.n236 B.n235 163.367
R199 B.n235 B.n34 163.367
R200 B.n231 B.n34 163.367
R201 B.n231 B.n230 163.367
R202 B.n230 B.n229 163.367
R203 B.n229 B.n36 163.367
R204 B.n225 B.n36 163.367
R205 B.n225 B.n224 163.367
R206 B.n224 B.n223 163.367
R207 B.n223 B.n38 163.367
R208 B.n219 B.n38 163.367
R209 B.n219 B.n218 163.367
R210 B.n218 B.n217 163.367
R211 B.n217 B.n40 163.367
R212 B.n213 B.n40 163.367
R213 B.n213 B.n212 163.367
R214 B.n212 B.n211 163.367
R215 B.n211 B.n42 163.367
R216 B.n207 B.n42 163.367
R217 B.n207 B.n206 163.367
R218 B.n206 B.n205 163.367
R219 B.n205 B.n44 163.367
R220 B.n201 B.n44 163.367
R221 B.n201 B.n200 163.367
R222 B.n200 B.n199 163.367
R223 B.n199 B.n46 163.367
R224 B.n195 B.n46 163.367
R225 B.n195 B.n194 163.367
R226 B.n194 B.n193 163.367
R227 B.n193 B.n48 163.367
R228 B.n189 B.n48 163.367
R229 B.n189 B.n188 163.367
R230 B.n188 B.n187 163.367
R231 B.n187 B.n50 163.367
R232 B.n183 B.n50 163.367
R233 B.n183 B.n182 163.367
R234 B.n182 B.n181 163.367
R235 B.n181 B.n52 163.367
R236 B.n177 B.n52 163.367
R237 B.n177 B.n176 163.367
R238 B.n176 B.n175 163.367
R239 B.n175 B.n54 163.367
R240 B.n171 B.n54 163.367
R241 B.n171 B.n170 163.367
R242 B.n170 B.n169 163.367
R243 B.n169 B.n56 163.367
R244 B.n165 B.n56 163.367
R245 B.n165 B.n164 163.367
R246 B.n279 B.n278 163.367
R247 B.n278 B.n15 163.367
R248 B.n274 B.n15 163.367
R249 B.n274 B.n273 163.367
R250 B.n273 B.n272 163.367
R251 B.n272 B.n17 163.367
R252 B.n268 B.n17 163.367
R253 B.n268 B.n267 163.367
R254 B.n267 B.n266 163.367
R255 B.n266 B.n19 163.367
R256 B.n262 B.n19 163.367
R257 B.n262 B.n261 163.367
R258 B.n261 B.n260 163.367
R259 B.n260 B.n24 163.367
R260 B.n256 B.n24 163.367
R261 B.n256 B.n255 163.367
R262 B.n255 B.n254 163.367
R263 B.n254 B.n26 163.367
R264 B.n249 B.n26 163.367
R265 B.n249 B.n248 163.367
R266 B.n248 B.n247 163.367
R267 B.n247 B.n30 163.367
R268 B.n243 B.n30 163.367
R269 B.n243 B.n242 163.367
R270 B.n242 B.n241 163.367
R271 B.n241 B.n32 163.367
R272 B.n280 B.n13 163.367
R273 B.n284 B.n13 163.367
R274 B.n285 B.n284 163.367
R275 B.n286 B.n285 163.367
R276 B.n286 B.n11 163.367
R277 B.n290 B.n11 163.367
R278 B.n291 B.n290 163.367
R279 B.n292 B.n291 163.367
R280 B.n292 B.n9 163.367
R281 B.n296 B.n9 163.367
R282 B.n297 B.n296 163.367
R283 B.n298 B.n297 163.367
R284 B.n298 B.n7 163.367
R285 B.n302 B.n7 163.367
R286 B.n303 B.n302 163.367
R287 B.n304 B.n303 163.367
R288 B.n304 B.n5 163.367
R289 B.n308 B.n5 163.367
R290 B.n309 B.n308 163.367
R291 B.n310 B.n309 163.367
R292 B.n310 B.n3 163.367
R293 B.n314 B.n3 163.367
R294 B.n315 B.n314 163.367
R295 B.n86 B.n2 163.367
R296 B.n89 B.n86 163.367
R297 B.n90 B.n89 163.367
R298 B.n91 B.n90 163.367
R299 B.n91 B.n84 163.367
R300 B.n95 B.n84 163.367
R301 B.n96 B.n95 163.367
R302 B.n97 B.n96 163.367
R303 B.n97 B.n82 163.367
R304 B.n101 B.n82 163.367
R305 B.n102 B.n101 163.367
R306 B.n103 B.n102 163.367
R307 B.n103 B.n80 163.367
R308 B.n107 B.n80 163.367
R309 B.n108 B.n107 163.367
R310 B.n109 B.n108 163.367
R311 B.n109 B.n78 163.367
R312 B.n113 B.n78 163.367
R313 B.n114 B.n113 163.367
R314 B.n115 B.n114 163.367
R315 B.n115 B.n76 163.367
R316 B.n119 B.n76 163.367
R317 B.n120 B.n119 163.367
R318 B.n135 B.n70 59.5399
R319 B.n149 B.n64 59.5399
R320 B.n252 B.n28 59.5399
R321 B.n22 B.n21 59.5399
R322 B.n70 B.n69 36.655
R323 B.n64 B.n63 36.655
R324 B.n28 B.n27 36.655
R325 B.n21 B.n20 36.655
R326 B.n162 B.n57 36.059
R327 B.n281 B.n14 36.059
R328 B.n239 B.n238 36.059
R329 B.n122 B.n75 36.059
R330 B B.n317 18.0485
R331 B.n282 B.n281 10.6151
R332 B.n283 B.n282 10.6151
R333 B.n283 B.n12 10.6151
R334 B.n287 B.n12 10.6151
R335 B.n288 B.n287 10.6151
R336 B.n289 B.n288 10.6151
R337 B.n289 B.n10 10.6151
R338 B.n293 B.n10 10.6151
R339 B.n294 B.n293 10.6151
R340 B.n295 B.n294 10.6151
R341 B.n295 B.n8 10.6151
R342 B.n299 B.n8 10.6151
R343 B.n300 B.n299 10.6151
R344 B.n301 B.n300 10.6151
R345 B.n301 B.n6 10.6151
R346 B.n305 B.n6 10.6151
R347 B.n306 B.n305 10.6151
R348 B.n307 B.n306 10.6151
R349 B.n307 B.n4 10.6151
R350 B.n311 B.n4 10.6151
R351 B.n312 B.n311 10.6151
R352 B.n313 B.n312 10.6151
R353 B.n313 B.n0 10.6151
R354 B.n277 B.n14 10.6151
R355 B.n277 B.n276 10.6151
R356 B.n276 B.n275 10.6151
R357 B.n275 B.n16 10.6151
R358 B.n271 B.n16 10.6151
R359 B.n271 B.n270 10.6151
R360 B.n270 B.n269 10.6151
R361 B.n269 B.n18 10.6151
R362 B.n265 B.n264 10.6151
R363 B.n264 B.n263 10.6151
R364 B.n263 B.n23 10.6151
R365 B.n259 B.n23 10.6151
R366 B.n259 B.n258 10.6151
R367 B.n258 B.n257 10.6151
R368 B.n257 B.n25 10.6151
R369 B.n253 B.n25 10.6151
R370 B.n251 B.n250 10.6151
R371 B.n250 B.n29 10.6151
R372 B.n246 B.n29 10.6151
R373 B.n246 B.n245 10.6151
R374 B.n245 B.n244 10.6151
R375 B.n244 B.n31 10.6151
R376 B.n240 B.n31 10.6151
R377 B.n240 B.n239 10.6151
R378 B.n238 B.n33 10.6151
R379 B.n234 B.n33 10.6151
R380 B.n234 B.n233 10.6151
R381 B.n233 B.n232 10.6151
R382 B.n232 B.n35 10.6151
R383 B.n228 B.n35 10.6151
R384 B.n228 B.n227 10.6151
R385 B.n227 B.n226 10.6151
R386 B.n226 B.n37 10.6151
R387 B.n222 B.n37 10.6151
R388 B.n222 B.n221 10.6151
R389 B.n221 B.n220 10.6151
R390 B.n220 B.n39 10.6151
R391 B.n216 B.n39 10.6151
R392 B.n216 B.n215 10.6151
R393 B.n215 B.n214 10.6151
R394 B.n214 B.n41 10.6151
R395 B.n210 B.n41 10.6151
R396 B.n210 B.n209 10.6151
R397 B.n209 B.n208 10.6151
R398 B.n208 B.n43 10.6151
R399 B.n204 B.n43 10.6151
R400 B.n204 B.n203 10.6151
R401 B.n203 B.n202 10.6151
R402 B.n202 B.n45 10.6151
R403 B.n198 B.n45 10.6151
R404 B.n198 B.n197 10.6151
R405 B.n197 B.n196 10.6151
R406 B.n196 B.n47 10.6151
R407 B.n192 B.n47 10.6151
R408 B.n192 B.n191 10.6151
R409 B.n191 B.n190 10.6151
R410 B.n190 B.n49 10.6151
R411 B.n186 B.n49 10.6151
R412 B.n186 B.n185 10.6151
R413 B.n185 B.n184 10.6151
R414 B.n184 B.n51 10.6151
R415 B.n180 B.n51 10.6151
R416 B.n180 B.n179 10.6151
R417 B.n179 B.n178 10.6151
R418 B.n178 B.n53 10.6151
R419 B.n174 B.n53 10.6151
R420 B.n174 B.n173 10.6151
R421 B.n173 B.n172 10.6151
R422 B.n172 B.n55 10.6151
R423 B.n168 B.n55 10.6151
R424 B.n168 B.n167 10.6151
R425 B.n167 B.n166 10.6151
R426 B.n166 B.n57 10.6151
R427 B.n87 B.n1 10.6151
R428 B.n88 B.n87 10.6151
R429 B.n88 B.n85 10.6151
R430 B.n92 B.n85 10.6151
R431 B.n93 B.n92 10.6151
R432 B.n94 B.n93 10.6151
R433 B.n94 B.n83 10.6151
R434 B.n98 B.n83 10.6151
R435 B.n99 B.n98 10.6151
R436 B.n100 B.n99 10.6151
R437 B.n100 B.n81 10.6151
R438 B.n104 B.n81 10.6151
R439 B.n105 B.n104 10.6151
R440 B.n106 B.n105 10.6151
R441 B.n106 B.n79 10.6151
R442 B.n110 B.n79 10.6151
R443 B.n111 B.n110 10.6151
R444 B.n112 B.n111 10.6151
R445 B.n112 B.n77 10.6151
R446 B.n116 B.n77 10.6151
R447 B.n117 B.n116 10.6151
R448 B.n118 B.n117 10.6151
R449 B.n118 B.n75 10.6151
R450 B.n123 B.n122 10.6151
R451 B.n124 B.n123 10.6151
R452 B.n124 B.n73 10.6151
R453 B.n128 B.n73 10.6151
R454 B.n129 B.n128 10.6151
R455 B.n130 B.n129 10.6151
R456 B.n130 B.n71 10.6151
R457 B.n134 B.n71 10.6151
R458 B.n137 B.n136 10.6151
R459 B.n137 B.n67 10.6151
R460 B.n141 B.n67 10.6151
R461 B.n142 B.n141 10.6151
R462 B.n143 B.n142 10.6151
R463 B.n143 B.n65 10.6151
R464 B.n147 B.n65 10.6151
R465 B.n148 B.n147 10.6151
R466 B.n150 B.n61 10.6151
R467 B.n154 B.n61 10.6151
R468 B.n155 B.n154 10.6151
R469 B.n156 B.n155 10.6151
R470 B.n156 B.n59 10.6151
R471 B.n160 B.n59 10.6151
R472 B.n161 B.n160 10.6151
R473 B.n162 B.n161 10.6151
R474 B.n317 B.n0 8.11757
R475 B.n317 B.n1 8.11757
R476 B.n265 B.n22 6.5566
R477 B.n253 B.n252 6.5566
R478 B.n136 B.n135 6.5566
R479 B.n149 B.n148 6.5566
R480 B.n22 B.n18 4.05904
R481 B.n252 B.n251 4.05904
R482 B.n135 B.n134 4.05904
R483 B.n150 B.n149 4.05904
R484 VP.n4 VP.n3 176.226
R485 VP.n12 VP.n11 176.226
R486 VP.n10 VP.n0 161.3
R487 VP.n9 VP.n8 161.3
R488 VP.n7 VP.n1 161.3
R489 VP.n6 VP.n5 161.3
R490 VP.n9 VP.n1 56.5193
R491 VP.n2 VP.t2 50.0485
R492 VP.n2 VP.t1 49.727
R493 VP.n3 VP.n2 47.4381
R494 VP.n5 VP.n1 24.4675
R495 VP.n10 VP.n9 24.4675
R496 VP.n4 VP.t0 12.8229
R497 VP.n11 VP.t3 12.8229
R498 VP.n5 VP.n4 9.54263
R499 VP.n11 VP.n10 9.54263
R500 VP.n6 VP.n3 0.189894
R501 VP.n7 VP.n6 0.189894
R502 VP.n8 VP.n7 0.189894
R503 VP.n8 VP.n0 0.189894
R504 VP.n12 VP.n0 0.189894
R505 VP VP.n12 0.0516364
R506 VDD1 VDD1.n1 668.168
R507 VDD1 VDD1.n0 638.383
R508 VDD1.n0 VDD1.t3 39.1632
R509 VDD1.n0 VDD1.t2 39.1632
R510 VDD1.n1 VDD1.t0 39.1632
R511 VDD1.n1 VDD1.t1 39.1632
R512 VTAIL.n7 VTAIL.t3 660.808
R513 VTAIL.n0 VTAIL.t2 660.808
R514 VTAIL.n1 VTAIL.t4 660.808
R515 VTAIL.n2 VTAIL.t7 660.808
R516 VTAIL.n6 VTAIL.t6 660.808
R517 VTAIL.n5 VTAIL.t5 660.808
R518 VTAIL.n4 VTAIL.t0 660.808
R519 VTAIL.n3 VTAIL.t1 660.808
R520 VTAIL.n7 VTAIL.n6 14.7117
R521 VTAIL.n3 VTAIL.n2 14.7117
R522 VTAIL.n4 VTAIL.n3 1.62981
R523 VTAIL.n6 VTAIL.n5 1.62981
R524 VTAIL.n2 VTAIL.n1 1.62981
R525 VTAIL VTAIL.n0 0.873345
R526 VTAIL VTAIL.n7 0.756965
R527 VTAIL.n5 VTAIL.n4 0.470328
R528 VTAIL.n1 VTAIL.n0 0.470328
R529 VN.n0 VN.t2 50.0485
R530 VN.n1 VN.t1 50.0485
R531 VN.n0 VN.t3 49.727
R532 VN.n1 VN.t0 49.727
R533 VN VN.n1 47.8188
R534 VN VN.n0 12.8529
R535 VDD2.n2 VDD2.n0 667.643
R536 VDD2.n2 VDD2.n1 638.324
R537 VDD2.n1 VDD2.t3 39.1632
R538 VDD2.n1 VDD2.t2 39.1632
R539 VDD2.n0 VDD2.t1 39.1632
R540 VDD2.n0 VDD2.t0 39.1632
R541 VDD2 VDD2.n2 0.0586897
C0 B VDD2 0.812281f
C1 VTAIL VDD2 2.24421f
C2 VTAIL B 0.909698f
C3 VDD1 VDD2 0.774965f
C4 B VDD1 0.77661f
C5 VTAIL VDD1 2.19698f
C6 VP VDD2 0.336876f
C7 B VP 1.17073f
C8 w_n2104_n1134# VDD2 0.972752f
C9 VTAIL VP 1.04245f
C10 B w_n2104_n1134# 4.85427f
C11 VDD1 VP 0.760476f
C12 VTAIL w_n2104_n1134# 1.27406f
C13 VDD1 w_n2104_n1134# 0.941046f
C14 VN VDD2 0.581034f
C15 VP w_n2104_n1134# 3.37495f
C16 B VN 0.732446f
C17 VTAIL VN 1.02834f
C18 VDD1 VN 0.155465f
C19 VP VN 3.38134f
C20 w_n2104_n1134# VN 3.11545f
C21 VDD2 VSUBS 0.502464f
C22 VDD1 VSUBS 2.701866f
C23 VTAIL VSUBS 0.344975f
C24 VN VSUBS 4.74609f
C25 VP VSUBS 1.195011f
C26 B VSUBS 2.302667f
C27 w_n2104_n1134# VSUBS 30.8278f
C28 VDD2.t1 VSUBS 0.015772f
C29 VDD2.t0 VSUBS 0.015772f
C30 VDD2.n0 VSUBS 0.063274f
C31 VDD2.t3 VSUBS 0.015772f
C32 VDD2.t2 VSUBS 0.015772f
C33 VDD2.n1 VSUBS 0.033873f
C34 VDD2.n2 VSUBS 1.90835f
C35 VN.t2 VSUBS 0.409435f
C36 VN.t3 VSUBS 0.407208f
C37 VN.n0 VSUBS 0.288559f
C38 VN.t1 VSUBS 0.409435f
C39 VN.t0 VSUBS 0.407208f
C40 VN.n1 VSUBS 1.83447f
C41 VTAIL.t2 VSUBS 0.07743f
C42 VTAIL.n0 VSUBS 0.154466f
C43 VTAIL.t4 VSUBS 0.07743f
C44 VTAIL.n1 VSUBS 0.217761f
C45 VTAIL.t7 VSUBS 0.07743f
C46 VTAIL.n2 VSUBS 0.72738f
C47 VTAIL.t1 VSUBS 0.07743f
C48 VTAIL.n3 VSUBS 0.72738f
C49 VTAIL.t0 VSUBS 0.07743f
C50 VTAIL.n4 VSUBS 0.217761f
C51 VTAIL.t5 VSUBS 0.07743f
C52 VTAIL.n5 VSUBS 0.217761f
C53 VTAIL.t6 VSUBS 0.07743f
C54 VTAIL.n6 VSUBS 0.72738f
C55 VTAIL.t3 VSUBS 0.07743f
C56 VTAIL.n7 VSUBS 0.654347f
C57 VDD1.t3 VSUBS 0.01516f
C58 VDD1.t2 VSUBS 0.01516f
C59 VDD1.n0 VSUBS 0.032577f
C60 VDD1.t0 VSUBS 0.01516f
C61 VDD1.t1 VSUBS 0.01516f
C62 VDD1.n1 VSUBS 0.063421f
C63 VP.n0 VSUBS 0.063209f
C64 VP.t3 VSUBS 0.137249f
C65 VP.n1 VSUBS 0.092274f
C66 VP.t2 VSUBS 0.433929f
C67 VP.t1 VSUBS 0.431569f
C68 VP.n2 VSUBS 1.9087f
C69 VP.n3 VSUBS 2.51686f
C70 VP.t0 VSUBS 0.137249f
C71 VP.n4 VSUBS 0.269585f
C72 VP.n5 VSUBS 0.082324f
C73 VP.n6 VSUBS 0.063209f
C74 VP.n7 VSUBS 0.063209f
C75 VP.n8 VSUBS 0.063209f
C76 VP.n9 VSUBS 0.092274f
C77 VP.n10 VSUBS 0.082324f
C78 VP.n11 VSUBS 0.269585f
C79 VP.n12 VSUBS 0.061474f
C80 B.n0 VSUBS 0.00967f
C81 B.n1 VSUBS 0.00967f
C82 B.n2 VSUBS 0.014302f
C83 B.n3 VSUBS 0.01096f
C84 B.n4 VSUBS 0.01096f
C85 B.n5 VSUBS 0.01096f
C86 B.n6 VSUBS 0.01096f
C87 B.n7 VSUBS 0.01096f
C88 B.n8 VSUBS 0.01096f
C89 B.n9 VSUBS 0.01096f
C90 B.n10 VSUBS 0.01096f
C91 B.n11 VSUBS 0.01096f
C92 B.n12 VSUBS 0.01096f
C93 B.n13 VSUBS 0.01096f
C94 B.n14 VSUBS 0.028186f
C95 B.n15 VSUBS 0.01096f
C96 B.n16 VSUBS 0.01096f
C97 B.n17 VSUBS 0.01096f
C98 B.n18 VSUBS 0.007575f
C99 B.n19 VSUBS 0.01096f
C100 B.t10 VSUBS 0.02501f
C101 B.t11 VSUBS 0.027412f
C102 B.t9 VSUBS 0.105759f
C103 B.n20 VSUBS 0.071714f
C104 B.n21 VSUBS 0.060631f
C105 B.n22 VSUBS 0.025392f
C106 B.n23 VSUBS 0.01096f
C107 B.n24 VSUBS 0.01096f
C108 B.n25 VSUBS 0.01096f
C109 B.n26 VSUBS 0.01096f
C110 B.t4 VSUBS 0.02501f
C111 B.t5 VSUBS 0.027412f
C112 B.t3 VSUBS 0.105759f
C113 B.n27 VSUBS 0.071714f
C114 B.n28 VSUBS 0.060631f
C115 B.n29 VSUBS 0.01096f
C116 B.n30 VSUBS 0.01096f
C117 B.n31 VSUBS 0.01096f
C118 B.n32 VSUBS 0.028186f
C119 B.n33 VSUBS 0.01096f
C120 B.n34 VSUBS 0.01096f
C121 B.n35 VSUBS 0.01096f
C122 B.n36 VSUBS 0.01096f
C123 B.n37 VSUBS 0.01096f
C124 B.n38 VSUBS 0.01096f
C125 B.n39 VSUBS 0.01096f
C126 B.n40 VSUBS 0.01096f
C127 B.n41 VSUBS 0.01096f
C128 B.n42 VSUBS 0.01096f
C129 B.n43 VSUBS 0.01096f
C130 B.n44 VSUBS 0.01096f
C131 B.n45 VSUBS 0.01096f
C132 B.n46 VSUBS 0.01096f
C133 B.n47 VSUBS 0.01096f
C134 B.n48 VSUBS 0.01096f
C135 B.n49 VSUBS 0.01096f
C136 B.n50 VSUBS 0.01096f
C137 B.n51 VSUBS 0.01096f
C138 B.n52 VSUBS 0.01096f
C139 B.n53 VSUBS 0.01096f
C140 B.n54 VSUBS 0.01096f
C141 B.n55 VSUBS 0.01096f
C142 B.n56 VSUBS 0.01096f
C143 B.n57 VSUBS 0.027785f
C144 B.n58 VSUBS 0.01096f
C145 B.n59 VSUBS 0.01096f
C146 B.n60 VSUBS 0.01096f
C147 B.n61 VSUBS 0.01096f
C148 B.n62 VSUBS 0.01096f
C149 B.t8 VSUBS 0.02501f
C150 B.t7 VSUBS 0.027412f
C151 B.t6 VSUBS 0.105759f
C152 B.n63 VSUBS 0.071714f
C153 B.n64 VSUBS 0.060631f
C154 B.n65 VSUBS 0.01096f
C155 B.n66 VSUBS 0.01096f
C156 B.n67 VSUBS 0.01096f
C157 B.n68 VSUBS 0.01096f
C158 B.t2 VSUBS 0.02501f
C159 B.t1 VSUBS 0.027412f
C160 B.t0 VSUBS 0.105759f
C161 B.n69 VSUBS 0.071714f
C162 B.n70 VSUBS 0.060631f
C163 B.n71 VSUBS 0.01096f
C164 B.n72 VSUBS 0.01096f
C165 B.n73 VSUBS 0.01096f
C166 B.n74 VSUBS 0.01096f
C167 B.n75 VSUBS 0.026612f
C168 B.n76 VSUBS 0.01096f
C169 B.n77 VSUBS 0.01096f
C170 B.n78 VSUBS 0.01096f
C171 B.n79 VSUBS 0.01096f
C172 B.n80 VSUBS 0.01096f
C173 B.n81 VSUBS 0.01096f
C174 B.n82 VSUBS 0.01096f
C175 B.n83 VSUBS 0.01096f
C176 B.n84 VSUBS 0.01096f
C177 B.n85 VSUBS 0.01096f
C178 B.n86 VSUBS 0.01096f
C179 B.n87 VSUBS 0.01096f
C180 B.n88 VSUBS 0.01096f
C181 B.n89 VSUBS 0.01096f
C182 B.n90 VSUBS 0.01096f
C183 B.n91 VSUBS 0.01096f
C184 B.n92 VSUBS 0.01096f
C185 B.n93 VSUBS 0.01096f
C186 B.n94 VSUBS 0.01096f
C187 B.n95 VSUBS 0.01096f
C188 B.n96 VSUBS 0.01096f
C189 B.n97 VSUBS 0.01096f
C190 B.n98 VSUBS 0.01096f
C191 B.n99 VSUBS 0.01096f
C192 B.n100 VSUBS 0.01096f
C193 B.n101 VSUBS 0.01096f
C194 B.n102 VSUBS 0.01096f
C195 B.n103 VSUBS 0.01096f
C196 B.n104 VSUBS 0.01096f
C197 B.n105 VSUBS 0.01096f
C198 B.n106 VSUBS 0.01096f
C199 B.n107 VSUBS 0.01096f
C200 B.n108 VSUBS 0.01096f
C201 B.n109 VSUBS 0.01096f
C202 B.n110 VSUBS 0.01096f
C203 B.n111 VSUBS 0.01096f
C204 B.n112 VSUBS 0.01096f
C205 B.n113 VSUBS 0.01096f
C206 B.n114 VSUBS 0.01096f
C207 B.n115 VSUBS 0.01096f
C208 B.n116 VSUBS 0.01096f
C209 B.n117 VSUBS 0.01096f
C210 B.n118 VSUBS 0.01096f
C211 B.n119 VSUBS 0.01096f
C212 B.n120 VSUBS 0.026612f
C213 B.n121 VSUBS 0.028186f
C214 B.n122 VSUBS 0.028186f
C215 B.n123 VSUBS 0.01096f
C216 B.n124 VSUBS 0.01096f
C217 B.n125 VSUBS 0.01096f
C218 B.n126 VSUBS 0.01096f
C219 B.n127 VSUBS 0.01096f
C220 B.n128 VSUBS 0.01096f
C221 B.n129 VSUBS 0.01096f
C222 B.n130 VSUBS 0.01096f
C223 B.n131 VSUBS 0.01096f
C224 B.n132 VSUBS 0.01096f
C225 B.n133 VSUBS 0.01096f
C226 B.n134 VSUBS 0.007575f
C227 B.n135 VSUBS 0.025392f
C228 B.n136 VSUBS 0.008864f
C229 B.n137 VSUBS 0.01096f
C230 B.n138 VSUBS 0.01096f
C231 B.n139 VSUBS 0.01096f
C232 B.n140 VSUBS 0.01096f
C233 B.n141 VSUBS 0.01096f
C234 B.n142 VSUBS 0.01096f
C235 B.n143 VSUBS 0.01096f
C236 B.n144 VSUBS 0.01096f
C237 B.n145 VSUBS 0.01096f
C238 B.n146 VSUBS 0.01096f
C239 B.n147 VSUBS 0.01096f
C240 B.n148 VSUBS 0.008864f
C241 B.n149 VSUBS 0.025392f
C242 B.n150 VSUBS 0.007575f
C243 B.n151 VSUBS 0.01096f
C244 B.n152 VSUBS 0.01096f
C245 B.n153 VSUBS 0.01096f
C246 B.n154 VSUBS 0.01096f
C247 B.n155 VSUBS 0.01096f
C248 B.n156 VSUBS 0.01096f
C249 B.n157 VSUBS 0.01096f
C250 B.n158 VSUBS 0.01096f
C251 B.n159 VSUBS 0.01096f
C252 B.n160 VSUBS 0.01096f
C253 B.n161 VSUBS 0.01096f
C254 B.n162 VSUBS 0.027013f
C255 B.n163 VSUBS 0.028186f
C256 B.n164 VSUBS 0.026612f
C257 B.n165 VSUBS 0.01096f
C258 B.n166 VSUBS 0.01096f
C259 B.n167 VSUBS 0.01096f
C260 B.n168 VSUBS 0.01096f
C261 B.n169 VSUBS 0.01096f
C262 B.n170 VSUBS 0.01096f
C263 B.n171 VSUBS 0.01096f
C264 B.n172 VSUBS 0.01096f
C265 B.n173 VSUBS 0.01096f
C266 B.n174 VSUBS 0.01096f
C267 B.n175 VSUBS 0.01096f
C268 B.n176 VSUBS 0.01096f
C269 B.n177 VSUBS 0.01096f
C270 B.n178 VSUBS 0.01096f
C271 B.n179 VSUBS 0.01096f
C272 B.n180 VSUBS 0.01096f
C273 B.n181 VSUBS 0.01096f
C274 B.n182 VSUBS 0.01096f
C275 B.n183 VSUBS 0.01096f
C276 B.n184 VSUBS 0.01096f
C277 B.n185 VSUBS 0.01096f
C278 B.n186 VSUBS 0.01096f
C279 B.n187 VSUBS 0.01096f
C280 B.n188 VSUBS 0.01096f
C281 B.n189 VSUBS 0.01096f
C282 B.n190 VSUBS 0.01096f
C283 B.n191 VSUBS 0.01096f
C284 B.n192 VSUBS 0.01096f
C285 B.n193 VSUBS 0.01096f
C286 B.n194 VSUBS 0.01096f
C287 B.n195 VSUBS 0.01096f
C288 B.n196 VSUBS 0.01096f
C289 B.n197 VSUBS 0.01096f
C290 B.n198 VSUBS 0.01096f
C291 B.n199 VSUBS 0.01096f
C292 B.n200 VSUBS 0.01096f
C293 B.n201 VSUBS 0.01096f
C294 B.n202 VSUBS 0.01096f
C295 B.n203 VSUBS 0.01096f
C296 B.n204 VSUBS 0.01096f
C297 B.n205 VSUBS 0.01096f
C298 B.n206 VSUBS 0.01096f
C299 B.n207 VSUBS 0.01096f
C300 B.n208 VSUBS 0.01096f
C301 B.n209 VSUBS 0.01096f
C302 B.n210 VSUBS 0.01096f
C303 B.n211 VSUBS 0.01096f
C304 B.n212 VSUBS 0.01096f
C305 B.n213 VSUBS 0.01096f
C306 B.n214 VSUBS 0.01096f
C307 B.n215 VSUBS 0.01096f
C308 B.n216 VSUBS 0.01096f
C309 B.n217 VSUBS 0.01096f
C310 B.n218 VSUBS 0.01096f
C311 B.n219 VSUBS 0.01096f
C312 B.n220 VSUBS 0.01096f
C313 B.n221 VSUBS 0.01096f
C314 B.n222 VSUBS 0.01096f
C315 B.n223 VSUBS 0.01096f
C316 B.n224 VSUBS 0.01096f
C317 B.n225 VSUBS 0.01096f
C318 B.n226 VSUBS 0.01096f
C319 B.n227 VSUBS 0.01096f
C320 B.n228 VSUBS 0.01096f
C321 B.n229 VSUBS 0.01096f
C322 B.n230 VSUBS 0.01096f
C323 B.n231 VSUBS 0.01096f
C324 B.n232 VSUBS 0.01096f
C325 B.n233 VSUBS 0.01096f
C326 B.n234 VSUBS 0.01096f
C327 B.n235 VSUBS 0.01096f
C328 B.n236 VSUBS 0.01096f
C329 B.n237 VSUBS 0.026612f
C330 B.n238 VSUBS 0.026612f
C331 B.n239 VSUBS 0.028186f
C332 B.n240 VSUBS 0.01096f
C333 B.n241 VSUBS 0.01096f
C334 B.n242 VSUBS 0.01096f
C335 B.n243 VSUBS 0.01096f
C336 B.n244 VSUBS 0.01096f
C337 B.n245 VSUBS 0.01096f
C338 B.n246 VSUBS 0.01096f
C339 B.n247 VSUBS 0.01096f
C340 B.n248 VSUBS 0.01096f
C341 B.n249 VSUBS 0.01096f
C342 B.n250 VSUBS 0.01096f
C343 B.n251 VSUBS 0.007575f
C344 B.n252 VSUBS 0.025392f
C345 B.n253 VSUBS 0.008864f
C346 B.n254 VSUBS 0.01096f
C347 B.n255 VSUBS 0.01096f
C348 B.n256 VSUBS 0.01096f
C349 B.n257 VSUBS 0.01096f
C350 B.n258 VSUBS 0.01096f
C351 B.n259 VSUBS 0.01096f
C352 B.n260 VSUBS 0.01096f
C353 B.n261 VSUBS 0.01096f
C354 B.n262 VSUBS 0.01096f
C355 B.n263 VSUBS 0.01096f
C356 B.n264 VSUBS 0.01096f
C357 B.n265 VSUBS 0.008864f
C358 B.n266 VSUBS 0.01096f
C359 B.n267 VSUBS 0.01096f
C360 B.n268 VSUBS 0.01096f
C361 B.n269 VSUBS 0.01096f
C362 B.n270 VSUBS 0.01096f
C363 B.n271 VSUBS 0.01096f
C364 B.n272 VSUBS 0.01096f
C365 B.n273 VSUBS 0.01096f
C366 B.n274 VSUBS 0.01096f
C367 B.n275 VSUBS 0.01096f
C368 B.n276 VSUBS 0.01096f
C369 B.n277 VSUBS 0.01096f
C370 B.n278 VSUBS 0.01096f
C371 B.n279 VSUBS 0.028186f
C372 B.n280 VSUBS 0.026612f
C373 B.n281 VSUBS 0.026612f
C374 B.n282 VSUBS 0.01096f
C375 B.n283 VSUBS 0.01096f
C376 B.n284 VSUBS 0.01096f
C377 B.n285 VSUBS 0.01096f
C378 B.n286 VSUBS 0.01096f
C379 B.n287 VSUBS 0.01096f
C380 B.n288 VSUBS 0.01096f
C381 B.n289 VSUBS 0.01096f
C382 B.n290 VSUBS 0.01096f
C383 B.n291 VSUBS 0.01096f
C384 B.n292 VSUBS 0.01096f
C385 B.n293 VSUBS 0.01096f
C386 B.n294 VSUBS 0.01096f
C387 B.n295 VSUBS 0.01096f
C388 B.n296 VSUBS 0.01096f
C389 B.n297 VSUBS 0.01096f
C390 B.n298 VSUBS 0.01096f
C391 B.n299 VSUBS 0.01096f
C392 B.n300 VSUBS 0.01096f
C393 B.n301 VSUBS 0.01096f
C394 B.n302 VSUBS 0.01096f
C395 B.n303 VSUBS 0.01096f
C396 B.n304 VSUBS 0.01096f
C397 B.n305 VSUBS 0.01096f
C398 B.n306 VSUBS 0.01096f
C399 B.n307 VSUBS 0.01096f
C400 B.n308 VSUBS 0.01096f
C401 B.n309 VSUBS 0.01096f
C402 B.n310 VSUBS 0.01096f
C403 B.n311 VSUBS 0.01096f
C404 B.n312 VSUBS 0.01096f
C405 B.n313 VSUBS 0.01096f
C406 B.n314 VSUBS 0.01096f
C407 B.n315 VSUBS 0.014302f
C408 B.n316 VSUBS 0.015235f
C409 B.n317 VSUBS 0.030296f
.ends

