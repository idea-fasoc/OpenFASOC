* NGSPICE file created from diff_pair_sample_0222.ext - technology: sky130A

.subckt diff_pair_sample_0222 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=1.34475 ps=8.48 w=8.15 l=2.2
X1 VDD1.t5 VP.t0 VTAIL.t2 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=1.34475 ps=8.48 w=8.15 l=2.2
X2 B.t11 B.t9 B.t10 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=0 ps=0 w=8.15 l=2.2
X3 VDD1.t4 VP.t1 VTAIL.t4 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=1.34475 ps=8.48 w=8.15 l=2.2
X4 VDD1.t3 VP.t2 VTAIL.t0 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=3.1785 ps=17.08 w=8.15 l=2.2
X5 VDD2.t0 VN.t1 VTAIL.t10 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=3.1785 ps=17.08 w=8.15 l=2.2
X6 B.t8 B.t6 B.t7 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=0 ps=0 w=8.15 l=2.2
X7 VDD2.t1 VN.t2 VTAIL.t9 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=3.1785 ps=17.08 w=8.15 l=2.2
X8 VTAIL.t3 VP.t3 VDD1.t2 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=1.34475 ps=8.48 w=8.15 l=2.2
X9 VDD2.t4 VN.t3 VTAIL.t8 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=1.34475 ps=8.48 w=8.15 l=2.2
X10 VTAIL.t7 VN.t4 VDD2.t3 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=1.34475 ps=8.48 w=8.15 l=2.2
X11 B.t5 B.t3 B.t4 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=0 ps=0 w=8.15 l=2.2
X12 VTAIL.t1 VP.t4 VDD1.t1 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=1.34475 ps=8.48 w=8.15 l=2.2
X13 B.t2 B.t0 B.t1 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=0 ps=0 w=8.15 l=2.2
X14 VDD2.t5 VN.t5 VTAIL.t6 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=3.1785 pd=17.08 as=1.34475 ps=8.48 w=8.15 l=2.2
X15 VDD1.t0 VP.t5 VTAIL.t5 w_n2994_n2598# sky130_fd_pr__pfet_01v8 ad=1.34475 pd=8.48 as=3.1785 ps=17.08 w=8.15 l=2.2
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n3 VN.t5 121.707
R11 VN.n17 VN.t2 121.707
R12 VN.n13 VN.n12 97.0549
R13 VN.n27 VN.n26 97.0549
R14 VN.n4 VN.t4 89.28
R15 VN.n12 VN.t1 89.28
R16 VN.n18 VN.t0 89.28
R17 VN.n26 VN.t3 89.28
R18 VN.n4 VN.n3 59.2585
R19 VN.n18 VN.n17 59.2585
R20 VN VN.n27 44.4489
R21 VN.n10 VN.n1 41.9503
R22 VN.n24 VN.n15 41.9503
R23 VN.n6 VN.n1 39.0365
R24 VN.n20 VN.n15 39.0365
R25 VN.n6 VN.n5 24.4675
R26 VN.n11 VN.n10 24.4675
R27 VN.n20 VN.n19 24.4675
R28 VN.n25 VN.n24 24.4675
R29 VN.n12 VN.n11 13.702
R30 VN.n26 VN.n25 13.702
R31 VN.n5 VN.n4 12.234
R32 VN.n19 VN.n18 12.234
R33 VN.n17 VN.n16 9.58252
R34 VN.n3 VN.n2 9.58252
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VDD2.n83 VDD2.n45 756.745
R47 VDD2.n38 VDD2.n0 756.745
R48 VDD2.n84 VDD2.n83 585
R49 VDD2.n82 VDD2.n81 585
R50 VDD2.n49 VDD2.n48 585
R51 VDD2.n76 VDD2.n75 585
R52 VDD2.n74 VDD2.n73 585
R53 VDD2.n53 VDD2.n52 585
R54 VDD2.n68 VDD2.n67 585
R55 VDD2.n66 VDD2.n65 585
R56 VDD2.n57 VDD2.n56 585
R57 VDD2.n60 VDD2.n59 585
R58 VDD2.n15 VDD2.n14 585
R59 VDD2.n12 VDD2.n11 585
R60 VDD2.n21 VDD2.n20 585
R61 VDD2.n23 VDD2.n22 585
R62 VDD2.n8 VDD2.n7 585
R63 VDD2.n29 VDD2.n28 585
R64 VDD2.n31 VDD2.n30 585
R65 VDD2.n4 VDD2.n3 585
R66 VDD2.n37 VDD2.n36 585
R67 VDD2.n39 VDD2.n38 585
R68 VDD2.t4 VDD2.n58 327.473
R69 VDD2.t5 VDD2.n13 327.473
R70 VDD2.n83 VDD2.n82 171.744
R71 VDD2.n82 VDD2.n48 171.744
R72 VDD2.n75 VDD2.n48 171.744
R73 VDD2.n75 VDD2.n74 171.744
R74 VDD2.n74 VDD2.n52 171.744
R75 VDD2.n67 VDD2.n52 171.744
R76 VDD2.n67 VDD2.n66 171.744
R77 VDD2.n66 VDD2.n56 171.744
R78 VDD2.n59 VDD2.n56 171.744
R79 VDD2.n14 VDD2.n11 171.744
R80 VDD2.n21 VDD2.n11 171.744
R81 VDD2.n22 VDD2.n21 171.744
R82 VDD2.n22 VDD2.n7 171.744
R83 VDD2.n29 VDD2.n7 171.744
R84 VDD2.n30 VDD2.n29 171.744
R85 VDD2.n30 VDD2.n3 171.744
R86 VDD2.n37 VDD2.n3 171.744
R87 VDD2.n38 VDD2.n37 171.744
R88 VDD2.n59 VDD2.t4 85.8723
R89 VDD2.n14 VDD2.t5 85.8723
R90 VDD2.n44 VDD2.n43 83.0828
R91 VDD2 VDD2.n89 83.0801
R92 VDD2.n44 VDD2.n42 50.2506
R93 VDD2.n88 VDD2.n87 48.6702
R94 VDD2.n88 VDD2.n44 37.8295
R95 VDD2.n60 VDD2.n58 16.3894
R96 VDD2.n15 VDD2.n13 16.3894
R97 VDD2.n61 VDD2.n57 12.8005
R98 VDD2.n16 VDD2.n12 12.8005
R99 VDD2.n65 VDD2.n64 12.0247
R100 VDD2.n20 VDD2.n19 12.0247
R101 VDD2.n68 VDD2.n55 11.249
R102 VDD2.n23 VDD2.n10 11.249
R103 VDD2.n69 VDD2.n53 10.4732
R104 VDD2.n24 VDD2.n8 10.4732
R105 VDD2.n73 VDD2.n72 9.69747
R106 VDD2.n28 VDD2.n27 9.69747
R107 VDD2.n87 VDD2.n86 9.45567
R108 VDD2.n42 VDD2.n41 9.45567
R109 VDD2.n86 VDD2.n85 9.3005
R110 VDD2.n47 VDD2.n46 9.3005
R111 VDD2.n80 VDD2.n79 9.3005
R112 VDD2.n78 VDD2.n77 9.3005
R113 VDD2.n51 VDD2.n50 9.3005
R114 VDD2.n72 VDD2.n71 9.3005
R115 VDD2.n70 VDD2.n69 9.3005
R116 VDD2.n55 VDD2.n54 9.3005
R117 VDD2.n64 VDD2.n63 9.3005
R118 VDD2.n62 VDD2.n61 9.3005
R119 VDD2.n2 VDD2.n1 9.3005
R120 VDD2.n41 VDD2.n40 9.3005
R121 VDD2.n33 VDD2.n32 9.3005
R122 VDD2.n6 VDD2.n5 9.3005
R123 VDD2.n27 VDD2.n26 9.3005
R124 VDD2.n25 VDD2.n24 9.3005
R125 VDD2.n10 VDD2.n9 9.3005
R126 VDD2.n19 VDD2.n18 9.3005
R127 VDD2.n17 VDD2.n16 9.3005
R128 VDD2.n35 VDD2.n34 9.3005
R129 VDD2.n76 VDD2.n51 8.92171
R130 VDD2.n31 VDD2.n6 8.92171
R131 VDD2.n87 VDD2.n45 8.14595
R132 VDD2.n77 VDD2.n49 8.14595
R133 VDD2.n32 VDD2.n4 8.14595
R134 VDD2.n42 VDD2.n0 8.14595
R135 VDD2.n85 VDD2.n84 7.3702
R136 VDD2.n81 VDD2.n80 7.3702
R137 VDD2.n36 VDD2.n35 7.3702
R138 VDD2.n40 VDD2.n39 7.3702
R139 VDD2.n84 VDD2.n47 6.59444
R140 VDD2.n81 VDD2.n47 6.59444
R141 VDD2.n36 VDD2.n2 6.59444
R142 VDD2.n39 VDD2.n2 6.59444
R143 VDD2.n85 VDD2.n45 5.81868
R144 VDD2.n80 VDD2.n49 5.81868
R145 VDD2.n35 VDD2.n4 5.81868
R146 VDD2.n40 VDD2.n0 5.81868
R147 VDD2.n77 VDD2.n76 5.04292
R148 VDD2.n32 VDD2.n31 5.04292
R149 VDD2.n73 VDD2.n51 4.26717
R150 VDD2.n28 VDD2.n6 4.26717
R151 VDD2.n89 VDD2.t2 3.98884
R152 VDD2.n89 VDD2.t1 3.98884
R153 VDD2.n43 VDD2.t3 3.98884
R154 VDD2.n43 VDD2.t0 3.98884
R155 VDD2.n62 VDD2.n58 3.70995
R156 VDD2.n17 VDD2.n13 3.70995
R157 VDD2.n72 VDD2.n53 3.49141
R158 VDD2.n27 VDD2.n8 3.49141
R159 VDD2.n69 VDD2.n68 2.71565
R160 VDD2.n24 VDD2.n23 2.71565
R161 VDD2.n65 VDD2.n55 1.93989
R162 VDD2.n20 VDD2.n10 1.93989
R163 VDD2 VDD2.n88 1.69447
R164 VDD2.n64 VDD2.n57 1.16414
R165 VDD2.n19 VDD2.n12 1.16414
R166 VDD2.n61 VDD2.n60 0.388379
R167 VDD2.n16 VDD2.n15 0.388379
R168 VDD2.n86 VDD2.n46 0.155672
R169 VDD2.n79 VDD2.n46 0.155672
R170 VDD2.n79 VDD2.n78 0.155672
R171 VDD2.n78 VDD2.n50 0.155672
R172 VDD2.n71 VDD2.n50 0.155672
R173 VDD2.n71 VDD2.n70 0.155672
R174 VDD2.n70 VDD2.n54 0.155672
R175 VDD2.n63 VDD2.n54 0.155672
R176 VDD2.n63 VDD2.n62 0.155672
R177 VDD2.n18 VDD2.n17 0.155672
R178 VDD2.n18 VDD2.n9 0.155672
R179 VDD2.n25 VDD2.n9 0.155672
R180 VDD2.n26 VDD2.n25 0.155672
R181 VDD2.n26 VDD2.n5 0.155672
R182 VDD2.n33 VDD2.n5 0.155672
R183 VDD2.n34 VDD2.n33 0.155672
R184 VDD2.n34 VDD2.n1 0.155672
R185 VDD2.n41 VDD2.n1 0.155672
R186 VTAIL.n178 VTAIL.n140 756.745
R187 VTAIL.n40 VTAIL.n2 756.745
R188 VTAIL.n134 VTAIL.n96 756.745
R189 VTAIL.n88 VTAIL.n50 756.745
R190 VTAIL.n155 VTAIL.n154 585
R191 VTAIL.n152 VTAIL.n151 585
R192 VTAIL.n161 VTAIL.n160 585
R193 VTAIL.n163 VTAIL.n162 585
R194 VTAIL.n148 VTAIL.n147 585
R195 VTAIL.n169 VTAIL.n168 585
R196 VTAIL.n171 VTAIL.n170 585
R197 VTAIL.n144 VTAIL.n143 585
R198 VTAIL.n177 VTAIL.n176 585
R199 VTAIL.n179 VTAIL.n178 585
R200 VTAIL.n17 VTAIL.n16 585
R201 VTAIL.n14 VTAIL.n13 585
R202 VTAIL.n23 VTAIL.n22 585
R203 VTAIL.n25 VTAIL.n24 585
R204 VTAIL.n10 VTAIL.n9 585
R205 VTAIL.n31 VTAIL.n30 585
R206 VTAIL.n33 VTAIL.n32 585
R207 VTAIL.n6 VTAIL.n5 585
R208 VTAIL.n39 VTAIL.n38 585
R209 VTAIL.n41 VTAIL.n40 585
R210 VTAIL.n135 VTAIL.n134 585
R211 VTAIL.n133 VTAIL.n132 585
R212 VTAIL.n100 VTAIL.n99 585
R213 VTAIL.n127 VTAIL.n126 585
R214 VTAIL.n125 VTAIL.n124 585
R215 VTAIL.n104 VTAIL.n103 585
R216 VTAIL.n119 VTAIL.n118 585
R217 VTAIL.n117 VTAIL.n116 585
R218 VTAIL.n108 VTAIL.n107 585
R219 VTAIL.n111 VTAIL.n110 585
R220 VTAIL.n89 VTAIL.n88 585
R221 VTAIL.n87 VTAIL.n86 585
R222 VTAIL.n54 VTAIL.n53 585
R223 VTAIL.n81 VTAIL.n80 585
R224 VTAIL.n79 VTAIL.n78 585
R225 VTAIL.n58 VTAIL.n57 585
R226 VTAIL.n73 VTAIL.n72 585
R227 VTAIL.n71 VTAIL.n70 585
R228 VTAIL.n62 VTAIL.n61 585
R229 VTAIL.n65 VTAIL.n64 585
R230 VTAIL.t10 VTAIL.n153 327.473
R231 VTAIL.t5 VTAIL.n15 327.473
R232 VTAIL.t0 VTAIL.n109 327.473
R233 VTAIL.t9 VTAIL.n63 327.473
R234 VTAIL.n154 VTAIL.n151 171.744
R235 VTAIL.n161 VTAIL.n151 171.744
R236 VTAIL.n162 VTAIL.n161 171.744
R237 VTAIL.n162 VTAIL.n147 171.744
R238 VTAIL.n169 VTAIL.n147 171.744
R239 VTAIL.n170 VTAIL.n169 171.744
R240 VTAIL.n170 VTAIL.n143 171.744
R241 VTAIL.n177 VTAIL.n143 171.744
R242 VTAIL.n178 VTAIL.n177 171.744
R243 VTAIL.n16 VTAIL.n13 171.744
R244 VTAIL.n23 VTAIL.n13 171.744
R245 VTAIL.n24 VTAIL.n23 171.744
R246 VTAIL.n24 VTAIL.n9 171.744
R247 VTAIL.n31 VTAIL.n9 171.744
R248 VTAIL.n32 VTAIL.n31 171.744
R249 VTAIL.n32 VTAIL.n5 171.744
R250 VTAIL.n39 VTAIL.n5 171.744
R251 VTAIL.n40 VTAIL.n39 171.744
R252 VTAIL.n134 VTAIL.n133 171.744
R253 VTAIL.n133 VTAIL.n99 171.744
R254 VTAIL.n126 VTAIL.n99 171.744
R255 VTAIL.n126 VTAIL.n125 171.744
R256 VTAIL.n125 VTAIL.n103 171.744
R257 VTAIL.n118 VTAIL.n103 171.744
R258 VTAIL.n118 VTAIL.n117 171.744
R259 VTAIL.n117 VTAIL.n107 171.744
R260 VTAIL.n110 VTAIL.n107 171.744
R261 VTAIL.n88 VTAIL.n87 171.744
R262 VTAIL.n87 VTAIL.n53 171.744
R263 VTAIL.n80 VTAIL.n53 171.744
R264 VTAIL.n80 VTAIL.n79 171.744
R265 VTAIL.n79 VTAIL.n57 171.744
R266 VTAIL.n72 VTAIL.n57 171.744
R267 VTAIL.n72 VTAIL.n71 171.744
R268 VTAIL.n71 VTAIL.n61 171.744
R269 VTAIL.n64 VTAIL.n61 171.744
R270 VTAIL.n154 VTAIL.t10 85.8723
R271 VTAIL.n16 VTAIL.t5 85.8723
R272 VTAIL.n110 VTAIL.t0 85.8723
R273 VTAIL.n64 VTAIL.t9 85.8723
R274 VTAIL.n95 VTAIL.n94 65.9142
R275 VTAIL.n49 VTAIL.n48 65.9142
R276 VTAIL.n1 VTAIL.n0 65.9141
R277 VTAIL.n47 VTAIL.n46 65.9141
R278 VTAIL.n183 VTAIL.n182 31.9914
R279 VTAIL.n45 VTAIL.n44 31.9914
R280 VTAIL.n139 VTAIL.n138 31.9914
R281 VTAIL.n93 VTAIL.n92 31.9914
R282 VTAIL.n49 VTAIL.n47 23.7548
R283 VTAIL.n183 VTAIL.n139 21.5738
R284 VTAIL.n155 VTAIL.n153 16.3894
R285 VTAIL.n17 VTAIL.n15 16.3894
R286 VTAIL.n111 VTAIL.n109 16.3894
R287 VTAIL.n65 VTAIL.n63 16.3894
R288 VTAIL.n156 VTAIL.n152 12.8005
R289 VTAIL.n18 VTAIL.n14 12.8005
R290 VTAIL.n112 VTAIL.n108 12.8005
R291 VTAIL.n66 VTAIL.n62 12.8005
R292 VTAIL.n160 VTAIL.n159 12.0247
R293 VTAIL.n22 VTAIL.n21 12.0247
R294 VTAIL.n116 VTAIL.n115 12.0247
R295 VTAIL.n70 VTAIL.n69 12.0247
R296 VTAIL.n163 VTAIL.n150 11.249
R297 VTAIL.n25 VTAIL.n12 11.249
R298 VTAIL.n119 VTAIL.n106 11.249
R299 VTAIL.n73 VTAIL.n60 11.249
R300 VTAIL.n164 VTAIL.n148 10.4732
R301 VTAIL.n26 VTAIL.n10 10.4732
R302 VTAIL.n120 VTAIL.n104 10.4732
R303 VTAIL.n74 VTAIL.n58 10.4732
R304 VTAIL.n168 VTAIL.n167 9.69747
R305 VTAIL.n30 VTAIL.n29 9.69747
R306 VTAIL.n124 VTAIL.n123 9.69747
R307 VTAIL.n78 VTAIL.n77 9.69747
R308 VTAIL.n182 VTAIL.n181 9.45567
R309 VTAIL.n44 VTAIL.n43 9.45567
R310 VTAIL.n138 VTAIL.n137 9.45567
R311 VTAIL.n92 VTAIL.n91 9.45567
R312 VTAIL.n142 VTAIL.n141 9.3005
R313 VTAIL.n181 VTAIL.n180 9.3005
R314 VTAIL.n173 VTAIL.n172 9.3005
R315 VTAIL.n146 VTAIL.n145 9.3005
R316 VTAIL.n167 VTAIL.n166 9.3005
R317 VTAIL.n165 VTAIL.n164 9.3005
R318 VTAIL.n150 VTAIL.n149 9.3005
R319 VTAIL.n159 VTAIL.n158 9.3005
R320 VTAIL.n157 VTAIL.n156 9.3005
R321 VTAIL.n175 VTAIL.n174 9.3005
R322 VTAIL.n4 VTAIL.n3 9.3005
R323 VTAIL.n43 VTAIL.n42 9.3005
R324 VTAIL.n35 VTAIL.n34 9.3005
R325 VTAIL.n8 VTAIL.n7 9.3005
R326 VTAIL.n29 VTAIL.n28 9.3005
R327 VTAIL.n27 VTAIL.n26 9.3005
R328 VTAIL.n12 VTAIL.n11 9.3005
R329 VTAIL.n21 VTAIL.n20 9.3005
R330 VTAIL.n19 VTAIL.n18 9.3005
R331 VTAIL.n37 VTAIL.n36 9.3005
R332 VTAIL.n98 VTAIL.n97 9.3005
R333 VTAIL.n131 VTAIL.n130 9.3005
R334 VTAIL.n129 VTAIL.n128 9.3005
R335 VTAIL.n102 VTAIL.n101 9.3005
R336 VTAIL.n123 VTAIL.n122 9.3005
R337 VTAIL.n121 VTAIL.n120 9.3005
R338 VTAIL.n106 VTAIL.n105 9.3005
R339 VTAIL.n115 VTAIL.n114 9.3005
R340 VTAIL.n113 VTAIL.n112 9.3005
R341 VTAIL.n137 VTAIL.n136 9.3005
R342 VTAIL.n91 VTAIL.n90 9.3005
R343 VTAIL.n52 VTAIL.n51 9.3005
R344 VTAIL.n85 VTAIL.n84 9.3005
R345 VTAIL.n83 VTAIL.n82 9.3005
R346 VTAIL.n56 VTAIL.n55 9.3005
R347 VTAIL.n77 VTAIL.n76 9.3005
R348 VTAIL.n75 VTAIL.n74 9.3005
R349 VTAIL.n60 VTAIL.n59 9.3005
R350 VTAIL.n69 VTAIL.n68 9.3005
R351 VTAIL.n67 VTAIL.n66 9.3005
R352 VTAIL.n171 VTAIL.n146 8.92171
R353 VTAIL.n33 VTAIL.n8 8.92171
R354 VTAIL.n127 VTAIL.n102 8.92171
R355 VTAIL.n81 VTAIL.n56 8.92171
R356 VTAIL.n172 VTAIL.n144 8.14595
R357 VTAIL.n182 VTAIL.n140 8.14595
R358 VTAIL.n34 VTAIL.n6 8.14595
R359 VTAIL.n44 VTAIL.n2 8.14595
R360 VTAIL.n138 VTAIL.n96 8.14595
R361 VTAIL.n128 VTAIL.n100 8.14595
R362 VTAIL.n92 VTAIL.n50 8.14595
R363 VTAIL.n82 VTAIL.n54 8.14595
R364 VTAIL.n176 VTAIL.n175 7.3702
R365 VTAIL.n180 VTAIL.n179 7.3702
R366 VTAIL.n38 VTAIL.n37 7.3702
R367 VTAIL.n42 VTAIL.n41 7.3702
R368 VTAIL.n136 VTAIL.n135 7.3702
R369 VTAIL.n132 VTAIL.n131 7.3702
R370 VTAIL.n90 VTAIL.n89 7.3702
R371 VTAIL.n86 VTAIL.n85 7.3702
R372 VTAIL.n176 VTAIL.n142 6.59444
R373 VTAIL.n179 VTAIL.n142 6.59444
R374 VTAIL.n38 VTAIL.n4 6.59444
R375 VTAIL.n41 VTAIL.n4 6.59444
R376 VTAIL.n135 VTAIL.n98 6.59444
R377 VTAIL.n132 VTAIL.n98 6.59444
R378 VTAIL.n89 VTAIL.n52 6.59444
R379 VTAIL.n86 VTAIL.n52 6.59444
R380 VTAIL.n175 VTAIL.n144 5.81868
R381 VTAIL.n180 VTAIL.n140 5.81868
R382 VTAIL.n37 VTAIL.n6 5.81868
R383 VTAIL.n42 VTAIL.n2 5.81868
R384 VTAIL.n136 VTAIL.n96 5.81868
R385 VTAIL.n131 VTAIL.n100 5.81868
R386 VTAIL.n90 VTAIL.n50 5.81868
R387 VTAIL.n85 VTAIL.n54 5.81868
R388 VTAIL.n172 VTAIL.n171 5.04292
R389 VTAIL.n34 VTAIL.n33 5.04292
R390 VTAIL.n128 VTAIL.n127 5.04292
R391 VTAIL.n82 VTAIL.n81 5.04292
R392 VTAIL.n168 VTAIL.n146 4.26717
R393 VTAIL.n30 VTAIL.n8 4.26717
R394 VTAIL.n124 VTAIL.n102 4.26717
R395 VTAIL.n78 VTAIL.n56 4.26717
R396 VTAIL.n0 VTAIL.t6 3.98884
R397 VTAIL.n0 VTAIL.t7 3.98884
R398 VTAIL.n46 VTAIL.t2 3.98884
R399 VTAIL.n46 VTAIL.t1 3.98884
R400 VTAIL.n94 VTAIL.t4 3.98884
R401 VTAIL.n94 VTAIL.t3 3.98884
R402 VTAIL.n48 VTAIL.t8 3.98884
R403 VTAIL.n48 VTAIL.t11 3.98884
R404 VTAIL.n157 VTAIL.n153 3.70995
R405 VTAIL.n19 VTAIL.n15 3.70995
R406 VTAIL.n67 VTAIL.n63 3.70995
R407 VTAIL.n113 VTAIL.n109 3.70995
R408 VTAIL.n167 VTAIL.n148 3.49141
R409 VTAIL.n29 VTAIL.n10 3.49141
R410 VTAIL.n123 VTAIL.n104 3.49141
R411 VTAIL.n77 VTAIL.n58 3.49141
R412 VTAIL.n164 VTAIL.n163 2.71565
R413 VTAIL.n26 VTAIL.n25 2.71565
R414 VTAIL.n120 VTAIL.n119 2.71565
R415 VTAIL.n74 VTAIL.n73 2.71565
R416 VTAIL.n93 VTAIL.n49 2.18153
R417 VTAIL.n139 VTAIL.n95 2.18153
R418 VTAIL.n47 VTAIL.n45 2.18153
R419 VTAIL.n160 VTAIL.n150 1.93989
R420 VTAIL.n22 VTAIL.n12 1.93989
R421 VTAIL.n116 VTAIL.n106 1.93989
R422 VTAIL.n70 VTAIL.n60 1.93989
R423 VTAIL VTAIL.n183 1.57809
R424 VTAIL.n95 VTAIL.n93 1.56084
R425 VTAIL.n45 VTAIL.n1 1.56084
R426 VTAIL.n159 VTAIL.n152 1.16414
R427 VTAIL.n21 VTAIL.n14 1.16414
R428 VTAIL.n115 VTAIL.n108 1.16414
R429 VTAIL.n69 VTAIL.n62 1.16414
R430 VTAIL VTAIL.n1 0.603948
R431 VTAIL.n156 VTAIL.n155 0.388379
R432 VTAIL.n18 VTAIL.n17 0.388379
R433 VTAIL.n112 VTAIL.n111 0.388379
R434 VTAIL.n66 VTAIL.n65 0.388379
R435 VTAIL.n158 VTAIL.n157 0.155672
R436 VTAIL.n158 VTAIL.n149 0.155672
R437 VTAIL.n165 VTAIL.n149 0.155672
R438 VTAIL.n166 VTAIL.n165 0.155672
R439 VTAIL.n166 VTAIL.n145 0.155672
R440 VTAIL.n173 VTAIL.n145 0.155672
R441 VTAIL.n174 VTAIL.n173 0.155672
R442 VTAIL.n174 VTAIL.n141 0.155672
R443 VTAIL.n181 VTAIL.n141 0.155672
R444 VTAIL.n20 VTAIL.n19 0.155672
R445 VTAIL.n20 VTAIL.n11 0.155672
R446 VTAIL.n27 VTAIL.n11 0.155672
R447 VTAIL.n28 VTAIL.n27 0.155672
R448 VTAIL.n28 VTAIL.n7 0.155672
R449 VTAIL.n35 VTAIL.n7 0.155672
R450 VTAIL.n36 VTAIL.n35 0.155672
R451 VTAIL.n36 VTAIL.n3 0.155672
R452 VTAIL.n43 VTAIL.n3 0.155672
R453 VTAIL.n137 VTAIL.n97 0.155672
R454 VTAIL.n130 VTAIL.n97 0.155672
R455 VTAIL.n130 VTAIL.n129 0.155672
R456 VTAIL.n129 VTAIL.n101 0.155672
R457 VTAIL.n122 VTAIL.n101 0.155672
R458 VTAIL.n122 VTAIL.n121 0.155672
R459 VTAIL.n121 VTAIL.n105 0.155672
R460 VTAIL.n114 VTAIL.n105 0.155672
R461 VTAIL.n114 VTAIL.n113 0.155672
R462 VTAIL.n91 VTAIL.n51 0.155672
R463 VTAIL.n84 VTAIL.n51 0.155672
R464 VTAIL.n84 VTAIL.n83 0.155672
R465 VTAIL.n83 VTAIL.n55 0.155672
R466 VTAIL.n76 VTAIL.n55 0.155672
R467 VTAIL.n76 VTAIL.n75 0.155672
R468 VTAIL.n75 VTAIL.n59 0.155672
R469 VTAIL.n68 VTAIL.n59 0.155672
R470 VTAIL.n68 VTAIL.n67 0.155672
R471 VP.n11 VP.n8 161.3
R472 VP.n13 VP.n12 161.3
R473 VP.n14 VP.n7 161.3
R474 VP.n16 VP.n15 161.3
R475 VP.n17 VP.n6 161.3
R476 VP.n36 VP.n0 161.3
R477 VP.n35 VP.n34 161.3
R478 VP.n33 VP.n1 161.3
R479 VP.n32 VP.n31 161.3
R480 VP.n30 VP.n2 161.3
R481 VP.n28 VP.n27 161.3
R482 VP.n26 VP.n3 161.3
R483 VP.n25 VP.n24 161.3
R484 VP.n23 VP.n4 161.3
R485 VP.n22 VP.n21 161.3
R486 VP.n9 VP.t1 121.707
R487 VP.n20 VP.n5 97.0549
R488 VP.n38 VP.n37 97.0549
R489 VP.n19 VP.n18 97.0549
R490 VP.n5 VP.t0 89.28
R491 VP.n29 VP.t4 89.28
R492 VP.n37 VP.t5 89.28
R493 VP.n18 VP.t2 89.28
R494 VP.n10 VP.t3 89.28
R495 VP.n10 VP.n9 59.2585
R496 VP.n20 VP.n19 44.17
R497 VP.n24 VP.n23 41.9503
R498 VP.n35 VP.n1 41.9503
R499 VP.n16 VP.n7 41.9503
R500 VP.n24 VP.n3 39.0365
R501 VP.n31 VP.n1 39.0365
R502 VP.n12 VP.n7 39.0365
R503 VP.n23 VP.n22 24.4675
R504 VP.n28 VP.n3 24.4675
R505 VP.n31 VP.n30 24.4675
R506 VP.n36 VP.n35 24.4675
R507 VP.n17 VP.n16 24.4675
R508 VP.n12 VP.n11 24.4675
R509 VP.n22 VP.n5 13.702
R510 VP.n37 VP.n36 13.702
R511 VP.n18 VP.n17 13.702
R512 VP.n29 VP.n28 12.234
R513 VP.n30 VP.n29 12.234
R514 VP.n11 VP.n10 12.234
R515 VP.n9 VP.n8 9.58252
R516 VP.n19 VP.n6 0.278367
R517 VP.n21 VP.n20 0.278367
R518 VP.n38 VP.n0 0.278367
R519 VP.n13 VP.n8 0.189894
R520 VP.n14 VP.n13 0.189894
R521 VP.n15 VP.n14 0.189894
R522 VP.n15 VP.n6 0.189894
R523 VP.n21 VP.n4 0.189894
R524 VP.n25 VP.n4 0.189894
R525 VP.n26 VP.n25 0.189894
R526 VP.n27 VP.n26 0.189894
R527 VP.n27 VP.n2 0.189894
R528 VP.n32 VP.n2 0.189894
R529 VP.n33 VP.n32 0.189894
R530 VP.n34 VP.n33 0.189894
R531 VP.n34 VP.n0 0.189894
R532 VP VP.n38 0.153454
R533 VDD1.n38 VDD1.n0 756.745
R534 VDD1.n81 VDD1.n43 756.745
R535 VDD1.n39 VDD1.n38 585
R536 VDD1.n37 VDD1.n36 585
R537 VDD1.n4 VDD1.n3 585
R538 VDD1.n31 VDD1.n30 585
R539 VDD1.n29 VDD1.n28 585
R540 VDD1.n8 VDD1.n7 585
R541 VDD1.n23 VDD1.n22 585
R542 VDD1.n21 VDD1.n20 585
R543 VDD1.n12 VDD1.n11 585
R544 VDD1.n15 VDD1.n14 585
R545 VDD1.n58 VDD1.n57 585
R546 VDD1.n55 VDD1.n54 585
R547 VDD1.n64 VDD1.n63 585
R548 VDD1.n66 VDD1.n65 585
R549 VDD1.n51 VDD1.n50 585
R550 VDD1.n72 VDD1.n71 585
R551 VDD1.n74 VDD1.n73 585
R552 VDD1.n47 VDD1.n46 585
R553 VDD1.n80 VDD1.n79 585
R554 VDD1.n82 VDD1.n81 585
R555 VDD1.t4 VDD1.n13 327.473
R556 VDD1.t5 VDD1.n56 327.473
R557 VDD1.n38 VDD1.n37 171.744
R558 VDD1.n37 VDD1.n3 171.744
R559 VDD1.n30 VDD1.n3 171.744
R560 VDD1.n30 VDD1.n29 171.744
R561 VDD1.n29 VDD1.n7 171.744
R562 VDD1.n22 VDD1.n7 171.744
R563 VDD1.n22 VDD1.n21 171.744
R564 VDD1.n21 VDD1.n11 171.744
R565 VDD1.n14 VDD1.n11 171.744
R566 VDD1.n57 VDD1.n54 171.744
R567 VDD1.n64 VDD1.n54 171.744
R568 VDD1.n65 VDD1.n64 171.744
R569 VDD1.n65 VDD1.n50 171.744
R570 VDD1.n72 VDD1.n50 171.744
R571 VDD1.n73 VDD1.n72 171.744
R572 VDD1.n73 VDD1.n46 171.744
R573 VDD1.n80 VDD1.n46 171.744
R574 VDD1.n81 VDD1.n80 171.744
R575 VDD1.n14 VDD1.t4 85.8723
R576 VDD1.n57 VDD1.t5 85.8723
R577 VDD1.n87 VDD1.n86 83.0828
R578 VDD1.n89 VDD1.n88 82.593
R579 VDD1 VDD1.n42 50.3642
R580 VDD1.n87 VDD1.n85 50.2506
R581 VDD1.n89 VDD1.n87 39.503
R582 VDD1.n15 VDD1.n13 16.3894
R583 VDD1.n58 VDD1.n56 16.3894
R584 VDD1.n16 VDD1.n12 12.8005
R585 VDD1.n59 VDD1.n55 12.8005
R586 VDD1.n20 VDD1.n19 12.0247
R587 VDD1.n63 VDD1.n62 12.0247
R588 VDD1.n23 VDD1.n10 11.249
R589 VDD1.n66 VDD1.n53 11.249
R590 VDD1.n24 VDD1.n8 10.4732
R591 VDD1.n67 VDD1.n51 10.4732
R592 VDD1.n28 VDD1.n27 9.69747
R593 VDD1.n71 VDD1.n70 9.69747
R594 VDD1.n42 VDD1.n41 9.45567
R595 VDD1.n85 VDD1.n84 9.45567
R596 VDD1.n41 VDD1.n40 9.3005
R597 VDD1.n2 VDD1.n1 9.3005
R598 VDD1.n35 VDD1.n34 9.3005
R599 VDD1.n33 VDD1.n32 9.3005
R600 VDD1.n6 VDD1.n5 9.3005
R601 VDD1.n27 VDD1.n26 9.3005
R602 VDD1.n25 VDD1.n24 9.3005
R603 VDD1.n10 VDD1.n9 9.3005
R604 VDD1.n19 VDD1.n18 9.3005
R605 VDD1.n17 VDD1.n16 9.3005
R606 VDD1.n45 VDD1.n44 9.3005
R607 VDD1.n84 VDD1.n83 9.3005
R608 VDD1.n76 VDD1.n75 9.3005
R609 VDD1.n49 VDD1.n48 9.3005
R610 VDD1.n70 VDD1.n69 9.3005
R611 VDD1.n68 VDD1.n67 9.3005
R612 VDD1.n53 VDD1.n52 9.3005
R613 VDD1.n62 VDD1.n61 9.3005
R614 VDD1.n60 VDD1.n59 9.3005
R615 VDD1.n78 VDD1.n77 9.3005
R616 VDD1.n31 VDD1.n6 8.92171
R617 VDD1.n74 VDD1.n49 8.92171
R618 VDD1.n42 VDD1.n0 8.14595
R619 VDD1.n32 VDD1.n4 8.14595
R620 VDD1.n75 VDD1.n47 8.14595
R621 VDD1.n85 VDD1.n43 8.14595
R622 VDD1.n40 VDD1.n39 7.3702
R623 VDD1.n36 VDD1.n35 7.3702
R624 VDD1.n79 VDD1.n78 7.3702
R625 VDD1.n83 VDD1.n82 7.3702
R626 VDD1.n39 VDD1.n2 6.59444
R627 VDD1.n36 VDD1.n2 6.59444
R628 VDD1.n79 VDD1.n45 6.59444
R629 VDD1.n82 VDD1.n45 6.59444
R630 VDD1.n40 VDD1.n0 5.81868
R631 VDD1.n35 VDD1.n4 5.81868
R632 VDD1.n78 VDD1.n47 5.81868
R633 VDD1.n83 VDD1.n43 5.81868
R634 VDD1.n32 VDD1.n31 5.04292
R635 VDD1.n75 VDD1.n74 5.04292
R636 VDD1.n28 VDD1.n6 4.26717
R637 VDD1.n71 VDD1.n49 4.26717
R638 VDD1.n88 VDD1.t2 3.98884
R639 VDD1.n88 VDD1.t3 3.98884
R640 VDD1.n86 VDD1.t1 3.98884
R641 VDD1.n86 VDD1.t0 3.98884
R642 VDD1.n17 VDD1.n13 3.70995
R643 VDD1.n60 VDD1.n56 3.70995
R644 VDD1.n27 VDD1.n8 3.49141
R645 VDD1.n70 VDD1.n51 3.49141
R646 VDD1.n24 VDD1.n23 2.71565
R647 VDD1.n67 VDD1.n66 2.71565
R648 VDD1.n20 VDD1.n10 1.93989
R649 VDD1.n63 VDD1.n53 1.93989
R650 VDD1.n19 VDD1.n12 1.16414
R651 VDD1.n62 VDD1.n55 1.16414
R652 VDD1 VDD1.n89 0.487569
R653 VDD1.n16 VDD1.n15 0.388379
R654 VDD1.n59 VDD1.n58 0.388379
R655 VDD1.n41 VDD1.n1 0.155672
R656 VDD1.n34 VDD1.n1 0.155672
R657 VDD1.n34 VDD1.n33 0.155672
R658 VDD1.n33 VDD1.n5 0.155672
R659 VDD1.n26 VDD1.n5 0.155672
R660 VDD1.n26 VDD1.n25 0.155672
R661 VDD1.n25 VDD1.n9 0.155672
R662 VDD1.n18 VDD1.n9 0.155672
R663 VDD1.n18 VDD1.n17 0.155672
R664 VDD1.n61 VDD1.n60 0.155672
R665 VDD1.n61 VDD1.n52 0.155672
R666 VDD1.n68 VDD1.n52 0.155672
R667 VDD1.n69 VDD1.n68 0.155672
R668 VDD1.n69 VDD1.n48 0.155672
R669 VDD1.n76 VDD1.n48 0.155672
R670 VDD1.n77 VDD1.n76 0.155672
R671 VDD1.n77 VDD1.n44 0.155672
R672 VDD1.n84 VDD1.n44 0.155672
R673 B.n435 B.n60 585
R674 B.n437 B.n436 585
R675 B.n438 B.n59 585
R676 B.n440 B.n439 585
R677 B.n441 B.n58 585
R678 B.n443 B.n442 585
R679 B.n444 B.n57 585
R680 B.n446 B.n445 585
R681 B.n447 B.n56 585
R682 B.n449 B.n448 585
R683 B.n450 B.n55 585
R684 B.n452 B.n451 585
R685 B.n453 B.n54 585
R686 B.n455 B.n454 585
R687 B.n456 B.n53 585
R688 B.n458 B.n457 585
R689 B.n459 B.n52 585
R690 B.n461 B.n460 585
R691 B.n462 B.n51 585
R692 B.n464 B.n463 585
R693 B.n465 B.n50 585
R694 B.n467 B.n466 585
R695 B.n468 B.n49 585
R696 B.n470 B.n469 585
R697 B.n471 B.n48 585
R698 B.n473 B.n472 585
R699 B.n474 B.n47 585
R700 B.n476 B.n475 585
R701 B.n477 B.n46 585
R702 B.n479 B.n478 585
R703 B.n481 B.n43 585
R704 B.n483 B.n482 585
R705 B.n484 B.n42 585
R706 B.n486 B.n485 585
R707 B.n487 B.n41 585
R708 B.n489 B.n488 585
R709 B.n490 B.n40 585
R710 B.n492 B.n491 585
R711 B.n493 B.n39 585
R712 B.n495 B.n494 585
R713 B.n497 B.n496 585
R714 B.n498 B.n35 585
R715 B.n500 B.n499 585
R716 B.n501 B.n34 585
R717 B.n503 B.n502 585
R718 B.n504 B.n33 585
R719 B.n506 B.n505 585
R720 B.n507 B.n32 585
R721 B.n509 B.n508 585
R722 B.n510 B.n31 585
R723 B.n512 B.n511 585
R724 B.n513 B.n30 585
R725 B.n515 B.n514 585
R726 B.n516 B.n29 585
R727 B.n518 B.n517 585
R728 B.n519 B.n28 585
R729 B.n521 B.n520 585
R730 B.n522 B.n27 585
R731 B.n524 B.n523 585
R732 B.n525 B.n26 585
R733 B.n527 B.n526 585
R734 B.n528 B.n25 585
R735 B.n530 B.n529 585
R736 B.n531 B.n24 585
R737 B.n533 B.n532 585
R738 B.n534 B.n23 585
R739 B.n536 B.n535 585
R740 B.n537 B.n22 585
R741 B.n539 B.n538 585
R742 B.n540 B.n21 585
R743 B.n434 B.n433 585
R744 B.n432 B.n61 585
R745 B.n431 B.n430 585
R746 B.n429 B.n62 585
R747 B.n428 B.n427 585
R748 B.n426 B.n63 585
R749 B.n425 B.n424 585
R750 B.n423 B.n64 585
R751 B.n422 B.n421 585
R752 B.n420 B.n65 585
R753 B.n419 B.n418 585
R754 B.n417 B.n66 585
R755 B.n416 B.n415 585
R756 B.n414 B.n67 585
R757 B.n413 B.n412 585
R758 B.n411 B.n68 585
R759 B.n410 B.n409 585
R760 B.n408 B.n69 585
R761 B.n407 B.n406 585
R762 B.n405 B.n70 585
R763 B.n404 B.n403 585
R764 B.n402 B.n71 585
R765 B.n401 B.n400 585
R766 B.n399 B.n72 585
R767 B.n398 B.n397 585
R768 B.n396 B.n73 585
R769 B.n395 B.n394 585
R770 B.n393 B.n74 585
R771 B.n392 B.n391 585
R772 B.n390 B.n75 585
R773 B.n389 B.n388 585
R774 B.n387 B.n76 585
R775 B.n386 B.n385 585
R776 B.n384 B.n77 585
R777 B.n383 B.n382 585
R778 B.n381 B.n78 585
R779 B.n380 B.n379 585
R780 B.n378 B.n79 585
R781 B.n377 B.n376 585
R782 B.n375 B.n80 585
R783 B.n374 B.n373 585
R784 B.n372 B.n81 585
R785 B.n371 B.n370 585
R786 B.n369 B.n82 585
R787 B.n368 B.n367 585
R788 B.n366 B.n83 585
R789 B.n365 B.n364 585
R790 B.n363 B.n84 585
R791 B.n362 B.n361 585
R792 B.n360 B.n85 585
R793 B.n359 B.n358 585
R794 B.n357 B.n86 585
R795 B.n356 B.n355 585
R796 B.n354 B.n87 585
R797 B.n353 B.n352 585
R798 B.n351 B.n88 585
R799 B.n350 B.n349 585
R800 B.n348 B.n89 585
R801 B.n347 B.n346 585
R802 B.n345 B.n90 585
R803 B.n344 B.n343 585
R804 B.n342 B.n91 585
R805 B.n341 B.n340 585
R806 B.n339 B.n92 585
R807 B.n338 B.n337 585
R808 B.n336 B.n93 585
R809 B.n335 B.n334 585
R810 B.n333 B.n94 585
R811 B.n332 B.n331 585
R812 B.n330 B.n95 585
R813 B.n329 B.n328 585
R814 B.n327 B.n96 585
R815 B.n326 B.n325 585
R816 B.n324 B.n97 585
R817 B.n323 B.n322 585
R818 B.n321 B.n98 585
R819 B.n320 B.n319 585
R820 B.n213 B.n138 585
R821 B.n215 B.n214 585
R822 B.n216 B.n137 585
R823 B.n218 B.n217 585
R824 B.n219 B.n136 585
R825 B.n221 B.n220 585
R826 B.n222 B.n135 585
R827 B.n224 B.n223 585
R828 B.n225 B.n134 585
R829 B.n227 B.n226 585
R830 B.n228 B.n133 585
R831 B.n230 B.n229 585
R832 B.n231 B.n132 585
R833 B.n233 B.n232 585
R834 B.n234 B.n131 585
R835 B.n236 B.n235 585
R836 B.n237 B.n130 585
R837 B.n239 B.n238 585
R838 B.n240 B.n129 585
R839 B.n242 B.n241 585
R840 B.n243 B.n128 585
R841 B.n245 B.n244 585
R842 B.n246 B.n127 585
R843 B.n248 B.n247 585
R844 B.n249 B.n126 585
R845 B.n251 B.n250 585
R846 B.n252 B.n125 585
R847 B.n254 B.n253 585
R848 B.n255 B.n124 585
R849 B.n257 B.n256 585
R850 B.n259 B.n121 585
R851 B.n261 B.n260 585
R852 B.n262 B.n120 585
R853 B.n264 B.n263 585
R854 B.n265 B.n119 585
R855 B.n267 B.n266 585
R856 B.n268 B.n118 585
R857 B.n270 B.n269 585
R858 B.n271 B.n117 585
R859 B.n273 B.n272 585
R860 B.n275 B.n274 585
R861 B.n276 B.n113 585
R862 B.n278 B.n277 585
R863 B.n279 B.n112 585
R864 B.n281 B.n280 585
R865 B.n282 B.n111 585
R866 B.n284 B.n283 585
R867 B.n285 B.n110 585
R868 B.n287 B.n286 585
R869 B.n288 B.n109 585
R870 B.n290 B.n289 585
R871 B.n291 B.n108 585
R872 B.n293 B.n292 585
R873 B.n294 B.n107 585
R874 B.n296 B.n295 585
R875 B.n297 B.n106 585
R876 B.n299 B.n298 585
R877 B.n300 B.n105 585
R878 B.n302 B.n301 585
R879 B.n303 B.n104 585
R880 B.n305 B.n304 585
R881 B.n306 B.n103 585
R882 B.n308 B.n307 585
R883 B.n309 B.n102 585
R884 B.n311 B.n310 585
R885 B.n312 B.n101 585
R886 B.n314 B.n313 585
R887 B.n315 B.n100 585
R888 B.n317 B.n316 585
R889 B.n318 B.n99 585
R890 B.n212 B.n211 585
R891 B.n210 B.n139 585
R892 B.n209 B.n208 585
R893 B.n207 B.n140 585
R894 B.n206 B.n205 585
R895 B.n204 B.n141 585
R896 B.n203 B.n202 585
R897 B.n201 B.n142 585
R898 B.n200 B.n199 585
R899 B.n198 B.n143 585
R900 B.n197 B.n196 585
R901 B.n195 B.n144 585
R902 B.n194 B.n193 585
R903 B.n192 B.n145 585
R904 B.n191 B.n190 585
R905 B.n189 B.n146 585
R906 B.n188 B.n187 585
R907 B.n186 B.n147 585
R908 B.n185 B.n184 585
R909 B.n183 B.n148 585
R910 B.n182 B.n181 585
R911 B.n180 B.n149 585
R912 B.n179 B.n178 585
R913 B.n177 B.n150 585
R914 B.n176 B.n175 585
R915 B.n174 B.n151 585
R916 B.n173 B.n172 585
R917 B.n171 B.n152 585
R918 B.n170 B.n169 585
R919 B.n168 B.n153 585
R920 B.n167 B.n166 585
R921 B.n165 B.n154 585
R922 B.n164 B.n163 585
R923 B.n162 B.n155 585
R924 B.n161 B.n160 585
R925 B.n159 B.n156 585
R926 B.n158 B.n157 585
R927 B.n2 B.n0 585
R928 B.n597 B.n1 585
R929 B.n596 B.n595 585
R930 B.n594 B.n3 585
R931 B.n593 B.n592 585
R932 B.n591 B.n4 585
R933 B.n590 B.n589 585
R934 B.n588 B.n5 585
R935 B.n587 B.n586 585
R936 B.n585 B.n6 585
R937 B.n584 B.n583 585
R938 B.n582 B.n7 585
R939 B.n581 B.n580 585
R940 B.n579 B.n8 585
R941 B.n578 B.n577 585
R942 B.n576 B.n9 585
R943 B.n575 B.n574 585
R944 B.n573 B.n10 585
R945 B.n572 B.n571 585
R946 B.n570 B.n11 585
R947 B.n569 B.n568 585
R948 B.n567 B.n12 585
R949 B.n566 B.n565 585
R950 B.n564 B.n13 585
R951 B.n563 B.n562 585
R952 B.n561 B.n14 585
R953 B.n560 B.n559 585
R954 B.n558 B.n15 585
R955 B.n557 B.n556 585
R956 B.n555 B.n16 585
R957 B.n554 B.n553 585
R958 B.n552 B.n17 585
R959 B.n551 B.n550 585
R960 B.n549 B.n18 585
R961 B.n548 B.n547 585
R962 B.n546 B.n19 585
R963 B.n545 B.n544 585
R964 B.n543 B.n20 585
R965 B.n542 B.n541 585
R966 B.n599 B.n598 585
R967 B.n213 B.n212 492.5
R968 B.n542 B.n21 492.5
R969 B.n320 B.n99 492.5
R970 B.n435 B.n434 492.5
R971 B.n114 B.t2 355.666
R972 B.n44 B.t10 355.666
R973 B.n122 B.t5 355.666
R974 B.n36 B.t7 355.666
R975 B.n115 B.t1 306.599
R976 B.n45 B.t11 306.599
R977 B.n123 B.t4 306.599
R978 B.n37 B.t8 306.599
R979 B.n114 B.t0 296.632
R980 B.n122 B.t3 296.632
R981 B.n36 B.t6 296.632
R982 B.n44 B.t9 296.632
R983 B.n212 B.n139 163.367
R984 B.n208 B.n139 163.367
R985 B.n208 B.n207 163.367
R986 B.n207 B.n206 163.367
R987 B.n206 B.n141 163.367
R988 B.n202 B.n141 163.367
R989 B.n202 B.n201 163.367
R990 B.n201 B.n200 163.367
R991 B.n200 B.n143 163.367
R992 B.n196 B.n143 163.367
R993 B.n196 B.n195 163.367
R994 B.n195 B.n194 163.367
R995 B.n194 B.n145 163.367
R996 B.n190 B.n145 163.367
R997 B.n190 B.n189 163.367
R998 B.n189 B.n188 163.367
R999 B.n188 B.n147 163.367
R1000 B.n184 B.n147 163.367
R1001 B.n184 B.n183 163.367
R1002 B.n183 B.n182 163.367
R1003 B.n182 B.n149 163.367
R1004 B.n178 B.n149 163.367
R1005 B.n178 B.n177 163.367
R1006 B.n177 B.n176 163.367
R1007 B.n176 B.n151 163.367
R1008 B.n172 B.n151 163.367
R1009 B.n172 B.n171 163.367
R1010 B.n171 B.n170 163.367
R1011 B.n170 B.n153 163.367
R1012 B.n166 B.n153 163.367
R1013 B.n166 B.n165 163.367
R1014 B.n165 B.n164 163.367
R1015 B.n164 B.n155 163.367
R1016 B.n160 B.n155 163.367
R1017 B.n160 B.n159 163.367
R1018 B.n159 B.n158 163.367
R1019 B.n158 B.n2 163.367
R1020 B.n598 B.n2 163.367
R1021 B.n598 B.n597 163.367
R1022 B.n597 B.n596 163.367
R1023 B.n596 B.n3 163.367
R1024 B.n592 B.n3 163.367
R1025 B.n592 B.n591 163.367
R1026 B.n591 B.n590 163.367
R1027 B.n590 B.n5 163.367
R1028 B.n586 B.n5 163.367
R1029 B.n586 B.n585 163.367
R1030 B.n585 B.n584 163.367
R1031 B.n584 B.n7 163.367
R1032 B.n580 B.n7 163.367
R1033 B.n580 B.n579 163.367
R1034 B.n579 B.n578 163.367
R1035 B.n578 B.n9 163.367
R1036 B.n574 B.n9 163.367
R1037 B.n574 B.n573 163.367
R1038 B.n573 B.n572 163.367
R1039 B.n572 B.n11 163.367
R1040 B.n568 B.n11 163.367
R1041 B.n568 B.n567 163.367
R1042 B.n567 B.n566 163.367
R1043 B.n566 B.n13 163.367
R1044 B.n562 B.n13 163.367
R1045 B.n562 B.n561 163.367
R1046 B.n561 B.n560 163.367
R1047 B.n560 B.n15 163.367
R1048 B.n556 B.n15 163.367
R1049 B.n556 B.n555 163.367
R1050 B.n555 B.n554 163.367
R1051 B.n554 B.n17 163.367
R1052 B.n550 B.n17 163.367
R1053 B.n550 B.n549 163.367
R1054 B.n549 B.n548 163.367
R1055 B.n548 B.n19 163.367
R1056 B.n544 B.n19 163.367
R1057 B.n544 B.n543 163.367
R1058 B.n543 B.n542 163.367
R1059 B.n214 B.n213 163.367
R1060 B.n214 B.n137 163.367
R1061 B.n218 B.n137 163.367
R1062 B.n219 B.n218 163.367
R1063 B.n220 B.n219 163.367
R1064 B.n220 B.n135 163.367
R1065 B.n224 B.n135 163.367
R1066 B.n225 B.n224 163.367
R1067 B.n226 B.n225 163.367
R1068 B.n226 B.n133 163.367
R1069 B.n230 B.n133 163.367
R1070 B.n231 B.n230 163.367
R1071 B.n232 B.n231 163.367
R1072 B.n232 B.n131 163.367
R1073 B.n236 B.n131 163.367
R1074 B.n237 B.n236 163.367
R1075 B.n238 B.n237 163.367
R1076 B.n238 B.n129 163.367
R1077 B.n242 B.n129 163.367
R1078 B.n243 B.n242 163.367
R1079 B.n244 B.n243 163.367
R1080 B.n244 B.n127 163.367
R1081 B.n248 B.n127 163.367
R1082 B.n249 B.n248 163.367
R1083 B.n250 B.n249 163.367
R1084 B.n250 B.n125 163.367
R1085 B.n254 B.n125 163.367
R1086 B.n255 B.n254 163.367
R1087 B.n256 B.n255 163.367
R1088 B.n256 B.n121 163.367
R1089 B.n261 B.n121 163.367
R1090 B.n262 B.n261 163.367
R1091 B.n263 B.n262 163.367
R1092 B.n263 B.n119 163.367
R1093 B.n267 B.n119 163.367
R1094 B.n268 B.n267 163.367
R1095 B.n269 B.n268 163.367
R1096 B.n269 B.n117 163.367
R1097 B.n273 B.n117 163.367
R1098 B.n274 B.n273 163.367
R1099 B.n274 B.n113 163.367
R1100 B.n278 B.n113 163.367
R1101 B.n279 B.n278 163.367
R1102 B.n280 B.n279 163.367
R1103 B.n280 B.n111 163.367
R1104 B.n284 B.n111 163.367
R1105 B.n285 B.n284 163.367
R1106 B.n286 B.n285 163.367
R1107 B.n286 B.n109 163.367
R1108 B.n290 B.n109 163.367
R1109 B.n291 B.n290 163.367
R1110 B.n292 B.n291 163.367
R1111 B.n292 B.n107 163.367
R1112 B.n296 B.n107 163.367
R1113 B.n297 B.n296 163.367
R1114 B.n298 B.n297 163.367
R1115 B.n298 B.n105 163.367
R1116 B.n302 B.n105 163.367
R1117 B.n303 B.n302 163.367
R1118 B.n304 B.n303 163.367
R1119 B.n304 B.n103 163.367
R1120 B.n308 B.n103 163.367
R1121 B.n309 B.n308 163.367
R1122 B.n310 B.n309 163.367
R1123 B.n310 B.n101 163.367
R1124 B.n314 B.n101 163.367
R1125 B.n315 B.n314 163.367
R1126 B.n316 B.n315 163.367
R1127 B.n316 B.n99 163.367
R1128 B.n321 B.n320 163.367
R1129 B.n322 B.n321 163.367
R1130 B.n322 B.n97 163.367
R1131 B.n326 B.n97 163.367
R1132 B.n327 B.n326 163.367
R1133 B.n328 B.n327 163.367
R1134 B.n328 B.n95 163.367
R1135 B.n332 B.n95 163.367
R1136 B.n333 B.n332 163.367
R1137 B.n334 B.n333 163.367
R1138 B.n334 B.n93 163.367
R1139 B.n338 B.n93 163.367
R1140 B.n339 B.n338 163.367
R1141 B.n340 B.n339 163.367
R1142 B.n340 B.n91 163.367
R1143 B.n344 B.n91 163.367
R1144 B.n345 B.n344 163.367
R1145 B.n346 B.n345 163.367
R1146 B.n346 B.n89 163.367
R1147 B.n350 B.n89 163.367
R1148 B.n351 B.n350 163.367
R1149 B.n352 B.n351 163.367
R1150 B.n352 B.n87 163.367
R1151 B.n356 B.n87 163.367
R1152 B.n357 B.n356 163.367
R1153 B.n358 B.n357 163.367
R1154 B.n358 B.n85 163.367
R1155 B.n362 B.n85 163.367
R1156 B.n363 B.n362 163.367
R1157 B.n364 B.n363 163.367
R1158 B.n364 B.n83 163.367
R1159 B.n368 B.n83 163.367
R1160 B.n369 B.n368 163.367
R1161 B.n370 B.n369 163.367
R1162 B.n370 B.n81 163.367
R1163 B.n374 B.n81 163.367
R1164 B.n375 B.n374 163.367
R1165 B.n376 B.n375 163.367
R1166 B.n376 B.n79 163.367
R1167 B.n380 B.n79 163.367
R1168 B.n381 B.n380 163.367
R1169 B.n382 B.n381 163.367
R1170 B.n382 B.n77 163.367
R1171 B.n386 B.n77 163.367
R1172 B.n387 B.n386 163.367
R1173 B.n388 B.n387 163.367
R1174 B.n388 B.n75 163.367
R1175 B.n392 B.n75 163.367
R1176 B.n393 B.n392 163.367
R1177 B.n394 B.n393 163.367
R1178 B.n394 B.n73 163.367
R1179 B.n398 B.n73 163.367
R1180 B.n399 B.n398 163.367
R1181 B.n400 B.n399 163.367
R1182 B.n400 B.n71 163.367
R1183 B.n404 B.n71 163.367
R1184 B.n405 B.n404 163.367
R1185 B.n406 B.n405 163.367
R1186 B.n406 B.n69 163.367
R1187 B.n410 B.n69 163.367
R1188 B.n411 B.n410 163.367
R1189 B.n412 B.n411 163.367
R1190 B.n412 B.n67 163.367
R1191 B.n416 B.n67 163.367
R1192 B.n417 B.n416 163.367
R1193 B.n418 B.n417 163.367
R1194 B.n418 B.n65 163.367
R1195 B.n422 B.n65 163.367
R1196 B.n423 B.n422 163.367
R1197 B.n424 B.n423 163.367
R1198 B.n424 B.n63 163.367
R1199 B.n428 B.n63 163.367
R1200 B.n429 B.n428 163.367
R1201 B.n430 B.n429 163.367
R1202 B.n430 B.n61 163.367
R1203 B.n434 B.n61 163.367
R1204 B.n538 B.n21 163.367
R1205 B.n538 B.n537 163.367
R1206 B.n537 B.n536 163.367
R1207 B.n536 B.n23 163.367
R1208 B.n532 B.n23 163.367
R1209 B.n532 B.n531 163.367
R1210 B.n531 B.n530 163.367
R1211 B.n530 B.n25 163.367
R1212 B.n526 B.n25 163.367
R1213 B.n526 B.n525 163.367
R1214 B.n525 B.n524 163.367
R1215 B.n524 B.n27 163.367
R1216 B.n520 B.n27 163.367
R1217 B.n520 B.n519 163.367
R1218 B.n519 B.n518 163.367
R1219 B.n518 B.n29 163.367
R1220 B.n514 B.n29 163.367
R1221 B.n514 B.n513 163.367
R1222 B.n513 B.n512 163.367
R1223 B.n512 B.n31 163.367
R1224 B.n508 B.n31 163.367
R1225 B.n508 B.n507 163.367
R1226 B.n507 B.n506 163.367
R1227 B.n506 B.n33 163.367
R1228 B.n502 B.n33 163.367
R1229 B.n502 B.n501 163.367
R1230 B.n501 B.n500 163.367
R1231 B.n500 B.n35 163.367
R1232 B.n496 B.n35 163.367
R1233 B.n496 B.n495 163.367
R1234 B.n495 B.n39 163.367
R1235 B.n491 B.n39 163.367
R1236 B.n491 B.n490 163.367
R1237 B.n490 B.n489 163.367
R1238 B.n489 B.n41 163.367
R1239 B.n485 B.n41 163.367
R1240 B.n485 B.n484 163.367
R1241 B.n484 B.n483 163.367
R1242 B.n483 B.n43 163.367
R1243 B.n478 B.n43 163.367
R1244 B.n478 B.n477 163.367
R1245 B.n477 B.n476 163.367
R1246 B.n476 B.n47 163.367
R1247 B.n472 B.n47 163.367
R1248 B.n472 B.n471 163.367
R1249 B.n471 B.n470 163.367
R1250 B.n470 B.n49 163.367
R1251 B.n466 B.n49 163.367
R1252 B.n466 B.n465 163.367
R1253 B.n465 B.n464 163.367
R1254 B.n464 B.n51 163.367
R1255 B.n460 B.n51 163.367
R1256 B.n460 B.n459 163.367
R1257 B.n459 B.n458 163.367
R1258 B.n458 B.n53 163.367
R1259 B.n454 B.n53 163.367
R1260 B.n454 B.n453 163.367
R1261 B.n453 B.n452 163.367
R1262 B.n452 B.n55 163.367
R1263 B.n448 B.n55 163.367
R1264 B.n448 B.n447 163.367
R1265 B.n447 B.n446 163.367
R1266 B.n446 B.n57 163.367
R1267 B.n442 B.n57 163.367
R1268 B.n442 B.n441 163.367
R1269 B.n441 B.n440 163.367
R1270 B.n440 B.n59 163.367
R1271 B.n436 B.n59 163.367
R1272 B.n436 B.n435 163.367
R1273 B.n116 B.n115 59.5399
R1274 B.n258 B.n123 59.5399
R1275 B.n38 B.n37 59.5399
R1276 B.n480 B.n45 59.5399
R1277 B.n115 B.n114 49.0672
R1278 B.n123 B.n122 49.0672
R1279 B.n37 B.n36 49.0672
R1280 B.n45 B.n44 49.0672
R1281 B.n541 B.n540 32.0005
R1282 B.n433 B.n60 32.0005
R1283 B.n319 B.n318 32.0005
R1284 B.n211 B.n138 32.0005
R1285 B B.n599 18.0485
R1286 B.n540 B.n539 10.6151
R1287 B.n539 B.n22 10.6151
R1288 B.n535 B.n22 10.6151
R1289 B.n535 B.n534 10.6151
R1290 B.n534 B.n533 10.6151
R1291 B.n533 B.n24 10.6151
R1292 B.n529 B.n24 10.6151
R1293 B.n529 B.n528 10.6151
R1294 B.n528 B.n527 10.6151
R1295 B.n527 B.n26 10.6151
R1296 B.n523 B.n26 10.6151
R1297 B.n523 B.n522 10.6151
R1298 B.n522 B.n521 10.6151
R1299 B.n521 B.n28 10.6151
R1300 B.n517 B.n28 10.6151
R1301 B.n517 B.n516 10.6151
R1302 B.n516 B.n515 10.6151
R1303 B.n515 B.n30 10.6151
R1304 B.n511 B.n30 10.6151
R1305 B.n511 B.n510 10.6151
R1306 B.n510 B.n509 10.6151
R1307 B.n509 B.n32 10.6151
R1308 B.n505 B.n32 10.6151
R1309 B.n505 B.n504 10.6151
R1310 B.n504 B.n503 10.6151
R1311 B.n503 B.n34 10.6151
R1312 B.n499 B.n34 10.6151
R1313 B.n499 B.n498 10.6151
R1314 B.n498 B.n497 10.6151
R1315 B.n494 B.n493 10.6151
R1316 B.n493 B.n492 10.6151
R1317 B.n492 B.n40 10.6151
R1318 B.n488 B.n40 10.6151
R1319 B.n488 B.n487 10.6151
R1320 B.n487 B.n486 10.6151
R1321 B.n486 B.n42 10.6151
R1322 B.n482 B.n42 10.6151
R1323 B.n482 B.n481 10.6151
R1324 B.n479 B.n46 10.6151
R1325 B.n475 B.n46 10.6151
R1326 B.n475 B.n474 10.6151
R1327 B.n474 B.n473 10.6151
R1328 B.n473 B.n48 10.6151
R1329 B.n469 B.n48 10.6151
R1330 B.n469 B.n468 10.6151
R1331 B.n468 B.n467 10.6151
R1332 B.n467 B.n50 10.6151
R1333 B.n463 B.n50 10.6151
R1334 B.n463 B.n462 10.6151
R1335 B.n462 B.n461 10.6151
R1336 B.n461 B.n52 10.6151
R1337 B.n457 B.n52 10.6151
R1338 B.n457 B.n456 10.6151
R1339 B.n456 B.n455 10.6151
R1340 B.n455 B.n54 10.6151
R1341 B.n451 B.n54 10.6151
R1342 B.n451 B.n450 10.6151
R1343 B.n450 B.n449 10.6151
R1344 B.n449 B.n56 10.6151
R1345 B.n445 B.n56 10.6151
R1346 B.n445 B.n444 10.6151
R1347 B.n444 B.n443 10.6151
R1348 B.n443 B.n58 10.6151
R1349 B.n439 B.n58 10.6151
R1350 B.n439 B.n438 10.6151
R1351 B.n438 B.n437 10.6151
R1352 B.n437 B.n60 10.6151
R1353 B.n319 B.n98 10.6151
R1354 B.n323 B.n98 10.6151
R1355 B.n324 B.n323 10.6151
R1356 B.n325 B.n324 10.6151
R1357 B.n325 B.n96 10.6151
R1358 B.n329 B.n96 10.6151
R1359 B.n330 B.n329 10.6151
R1360 B.n331 B.n330 10.6151
R1361 B.n331 B.n94 10.6151
R1362 B.n335 B.n94 10.6151
R1363 B.n336 B.n335 10.6151
R1364 B.n337 B.n336 10.6151
R1365 B.n337 B.n92 10.6151
R1366 B.n341 B.n92 10.6151
R1367 B.n342 B.n341 10.6151
R1368 B.n343 B.n342 10.6151
R1369 B.n343 B.n90 10.6151
R1370 B.n347 B.n90 10.6151
R1371 B.n348 B.n347 10.6151
R1372 B.n349 B.n348 10.6151
R1373 B.n349 B.n88 10.6151
R1374 B.n353 B.n88 10.6151
R1375 B.n354 B.n353 10.6151
R1376 B.n355 B.n354 10.6151
R1377 B.n355 B.n86 10.6151
R1378 B.n359 B.n86 10.6151
R1379 B.n360 B.n359 10.6151
R1380 B.n361 B.n360 10.6151
R1381 B.n361 B.n84 10.6151
R1382 B.n365 B.n84 10.6151
R1383 B.n366 B.n365 10.6151
R1384 B.n367 B.n366 10.6151
R1385 B.n367 B.n82 10.6151
R1386 B.n371 B.n82 10.6151
R1387 B.n372 B.n371 10.6151
R1388 B.n373 B.n372 10.6151
R1389 B.n373 B.n80 10.6151
R1390 B.n377 B.n80 10.6151
R1391 B.n378 B.n377 10.6151
R1392 B.n379 B.n378 10.6151
R1393 B.n379 B.n78 10.6151
R1394 B.n383 B.n78 10.6151
R1395 B.n384 B.n383 10.6151
R1396 B.n385 B.n384 10.6151
R1397 B.n385 B.n76 10.6151
R1398 B.n389 B.n76 10.6151
R1399 B.n390 B.n389 10.6151
R1400 B.n391 B.n390 10.6151
R1401 B.n391 B.n74 10.6151
R1402 B.n395 B.n74 10.6151
R1403 B.n396 B.n395 10.6151
R1404 B.n397 B.n396 10.6151
R1405 B.n397 B.n72 10.6151
R1406 B.n401 B.n72 10.6151
R1407 B.n402 B.n401 10.6151
R1408 B.n403 B.n402 10.6151
R1409 B.n403 B.n70 10.6151
R1410 B.n407 B.n70 10.6151
R1411 B.n408 B.n407 10.6151
R1412 B.n409 B.n408 10.6151
R1413 B.n409 B.n68 10.6151
R1414 B.n413 B.n68 10.6151
R1415 B.n414 B.n413 10.6151
R1416 B.n415 B.n414 10.6151
R1417 B.n415 B.n66 10.6151
R1418 B.n419 B.n66 10.6151
R1419 B.n420 B.n419 10.6151
R1420 B.n421 B.n420 10.6151
R1421 B.n421 B.n64 10.6151
R1422 B.n425 B.n64 10.6151
R1423 B.n426 B.n425 10.6151
R1424 B.n427 B.n426 10.6151
R1425 B.n427 B.n62 10.6151
R1426 B.n431 B.n62 10.6151
R1427 B.n432 B.n431 10.6151
R1428 B.n433 B.n432 10.6151
R1429 B.n215 B.n138 10.6151
R1430 B.n216 B.n215 10.6151
R1431 B.n217 B.n216 10.6151
R1432 B.n217 B.n136 10.6151
R1433 B.n221 B.n136 10.6151
R1434 B.n222 B.n221 10.6151
R1435 B.n223 B.n222 10.6151
R1436 B.n223 B.n134 10.6151
R1437 B.n227 B.n134 10.6151
R1438 B.n228 B.n227 10.6151
R1439 B.n229 B.n228 10.6151
R1440 B.n229 B.n132 10.6151
R1441 B.n233 B.n132 10.6151
R1442 B.n234 B.n233 10.6151
R1443 B.n235 B.n234 10.6151
R1444 B.n235 B.n130 10.6151
R1445 B.n239 B.n130 10.6151
R1446 B.n240 B.n239 10.6151
R1447 B.n241 B.n240 10.6151
R1448 B.n241 B.n128 10.6151
R1449 B.n245 B.n128 10.6151
R1450 B.n246 B.n245 10.6151
R1451 B.n247 B.n246 10.6151
R1452 B.n247 B.n126 10.6151
R1453 B.n251 B.n126 10.6151
R1454 B.n252 B.n251 10.6151
R1455 B.n253 B.n252 10.6151
R1456 B.n253 B.n124 10.6151
R1457 B.n257 B.n124 10.6151
R1458 B.n260 B.n259 10.6151
R1459 B.n260 B.n120 10.6151
R1460 B.n264 B.n120 10.6151
R1461 B.n265 B.n264 10.6151
R1462 B.n266 B.n265 10.6151
R1463 B.n266 B.n118 10.6151
R1464 B.n270 B.n118 10.6151
R1465 B.n271 B.n270 10.6151
R1466 B.n272 B.n271 10.6151
R1467 B.n276 B.n275 10.6151
R1468 B.n277 B.n276 10.6151
R1469 B.n277 B.n112 10.6151
R1470 B.n281 B.n112 10.6151
R1471 B.n282 B.n281 10.6151
R1472 B.n283 B.n282 10.6151
R1473 B.n283 B.n110 10.6151
R1474 B.n287 B.n110 10.6151
R1475 B.n288 B.n287 10.6151
R1476 B.n289 B.n288 10.6151
R1477 B.n289 B.n108 10.6151
R1478 B.n293 B.n108 10.6151
R1479 B.n294 B.n293 10.6151
R1480 B.n295 B.n294 10.6151
R1481 B.n295 B.n106 10.6151
R1482 B.n299 B.n106 10.6151
R1483 B.n300 B.n299 10.6151
R1484 B.n301 B.n300 10.6151
R1485 B.n301 B.n104 10.6151
R1486 B.n305 B.n104 10.6151
R1487 B.n306 B.n305 10.6151
R1488 B.n307 B.n306 10.6151
R1489 B.n307 B.n102 10.6151
R1490 B.n311 B.n102 10.6151
R1491 B.n312 B.n311 10.6151
R1492 B.n313 B.n312 10.6151
R1493 B.n313 B.n100 10.6151
R1494 B.n317 B.n100 10.6151
R1495 B.n318 B.n317 10.6151
R1496 B.n211 B.n210 10.6151
R1497 B.n210 B.n209 10.6151
R1498 B.n209 B.n140 10.6151
R1499 B.n205 B.n140 10.6151
R1500 B.n205 B.n204 10.6151
R1501 B.n204 B.n203 10.6151
R1502 B.n203 B.n142 10.6151
R1503 B.n199 B.n142 10.6151
R1504 B.n199 B.n198 10.6151
R1505 B.n198 B.n197 10.6151
R1506 B.n197 B.n144 10.6151
R1507 B.n193 B.n144 10.6151
R1508 B.n193 B.n192 10.6151
R1509 B.n192 B.n191 10.6151
R1510 B.n191 B.n146 10.6151
R1511 B.n187 B.n146 10.6151
R1512 B.n187 B.n186 10.6151
R1513 B.n186 B.n185 10.6151
R1514 B.n185 B.n148 10.6151
R1515 B.n181 B.n148 10.6151
R1516 B.n181 B.n180 10.6151
R1517 B.n180 B.n179 10.6151
R1518 B.n179 B.n150 10.6151
R1519 B.n175 B.n150 10.6151
R1520 B.n175 B.n174 10.6151
R1521 B.n174 B.n173 10.6151
R1522 B.n173 B.n152 10.6151
R1523 B.n169 B.n152 10.6151
R1524 B.n169 B.n168 10.6151
R1525 B.n168 B.n167 10.6151
R1526 B.n167 B.n154 10.6151
R1527 B.n163 B.n154 10.6151
R1528 B.n163 B.n162 10.6151
R1529 B.n162 B.n161 10.6151
R1530 B.n161 B.n156 10.6151
R1531 B.n157 B.n156 10.6151
R1532 B.n157 B.n0 10.6151
R1533 B.n595 B.n1 10.6151
R1534 B.n595 B.n594 10.6151
R1535 B.n594 B.n593 10.6151
R1536 B.n593 B.n4 10.6151
R1537 B.n589 B.n4 10.6151
R1538 B.n589 B.n588 10.6151
R1539 B.n588 B.n587 10.6151
R1540 B.n587 B.n6 10.6151
R1541 B.n583 B.n6 10.6151
R1542 B.n583 B.n582 10.6151
R1543 B.n582 B.n581 10.6151
R1544 B.n581 B.n8 10.6151
R1545 B.n577 B.n8 10.6151
R1546 B.n577 B.n576 10.6151
R1547 B.n576 B.n575 10.6151
R1548 B.n575 B.n10 10.6151
R1549 B.n571 B.n10 10.6151
R1550 B.n571 B.n570 10.6151
R1551 B.n570 B.n569 10.6151
R1552 B.n569 B.n12 10.6151
R1553 B.n565 B.n12 10.6151
R1554 B.n565 B.n564 10.6151
R1555 B.n564 B.n563 10.6151
R1556 B.n563 B.n14 10.6151
R1557 B.n559 B.n14 10.6151
R1558 B.n559 B.n558 10.6151
R1559 B.n558 B.n557 10.6151
R1560 B.n557 B.n16 10.6151
R1561 B.n553 B.n16 10.6151
R1562 B.n553 B.n552 10.6151
R1563 B.n552 B.n551 10.6151
R1564 B.n551 B.n18 10.6151
R1565 B.n547 B.n18 10.6151
R1566 B.n547 B.n546 10.6151
R1567 B.n546 B.n545 10.6151
R1568 B.n545 B.n20 10.6151
R1569 B.n541 B.n20 10.6151
R1570 B.n497 B.n38 9.36635
R1571 B.n480 B.n479 9.36635
R1572 B.n258 B.n257 9.36635
R1573 B.n275 B.n116 9.36635
R1574 B.n599 B.n0 2.81026
R1575 B.n599 B.n1 2.81026
R1576 B.n494 B.n38 1.24928
R1577 B.n481 B.n480 1.24928
R1578 B.n259 B.n258 1.24928
R1579 B.n272 B.n116 1.24928
C0 VDD1 VDD2 1.24933f
C1 VN VDD1 0.149994f
C2 w_n2994_n2598# VDD2 1.99417f
C3 VN w_n2994_n2598# 5.51445f
C4 VP VDD2 0.423885f
C5 VN VP 5.82769f
C6 B VDD2 1.75083f
C7 VTAIL VDD2 6.261549f
C8 VN B 1.03753f
C9 VN VTAIL 4.76692f
C10 VDD1 w_n2994_n2598# 1.92185f
C11 VDD1 VP 4.80784f
C12 VP w_n2994_n2598# 5.90042f
C13 VDD1 B 1.68633f
C14 VTAIL VDD1 6.21283f
C15 VN VDD2 4.53651f
C16 B w_n2994_n2598# 8.04383f
C17 VTAIL w_n2994_n2598# 2.39389f
C18 B VP 1.67993f
C19 VTAIL VP 4.78118f
C20 VTAIL B 2.68747f
C21 VDD2 VSUBS 1.457778f
C22 VDD1 VSUBS 1.493303f
C23 VTAIL VSUBS 0.979806f
C24 VN VSUBS 5.32115f
C25 VP VSUBS 2.484722f
C26 B VSUBS 3.91404f
C27 w_n2994_n2598# VSUBS 96.466705f
C28 B.n0 VSUBS 0.004481f
C29 B.n1 VSUBS 0.004481f
C30 B.n2 VSUBS 0.007087f
C31 B.n3 VSUBS 0.007087f
C32 B.n4 VSUBS 0.007087f
C33 B.n5 VSUBS 0.007087f
C34 B.n6 VSUBS 0.007087f
C35 B.n7 VSUBS 0.007087f
C36 B.n8 VSUBS 0.007087f
C37 B.n9 VSUBS 0.007087f
C38 B.n10 VSUBS 0.007087f
C39 B.n11 VSUBS 0.007087f
C40 B.n12 VSUBS 0.007087f
C41 B.n13 VSUBS 0.007087f
C42 B.n14 VSUBS 0.007087f
C43 B.n15 VSUBS 0.007087f
C44 B.n16 VSUBS 0.007087f
C45 B.n17 VSUBS 0.007087f
C46 B.n18 VSUBS 0.007087f
C47 B.n19 VSUBS 0.007087f
C48 B.n20 VSUBS 0.007087f
C49 B.n21 VSUBS 0.016622f
C50 B.n22 VSUBS 0.007087f
C51 B.n23 VSUBS 0.007087f
C52 B.n24 VSUBS 0.007087f
C53 B.n25 VSUBS 0.007087f
C54 B.n26 VSUBS 0.007087f
C55 B.n27 VSUBS 0.007087f
C56 B.n28 VSUBS 0.007087f
C57 B.n29 VSUBS 0.007087f
C58 B.n30 VSUBS 0.007087f
C59 B.n31 VSUBS 0.007087f
C60 B.n32 VSUBS 0.007087f
C61 B.n33 VSUBS 0.007087f
C62 B.n34 VSUBS 0.007087f
C63 B.n35 VSUBS 0.007087f
C64 B.t8 VSUBS 0.131478f
C65 B.t7 VSUBS 0.156918f
C66 B.t6 VSUBS 0.836981f
C67 B.n36 VSUBS 0.260234f
C68 B.n37 VSUBS 0.194509f
C69 B.n38 VSUBS 0.016419f
C70 B.n39 VSUBS 0.007087f
C71 B.n40 VSUBS 0.007087f
C72 B.n41 VSUBS 0.007087f
C73 B.n42 VSUBS 0.007087f
C74 B.n43 VSUBS 0.007087f
C75 B.t11 VSUBS 0.131481f
C76 B.t10 VSUBS 0.15692f
C77 B.t9 VSUBS 0.836981f
C78 B.n44 VSUBS 0.260232f
C79 B.n45 VSUBS 0.194507f
C80 B.n46 VSUBS 0.007087f
C81 B.n47 VSUBS 0.007087f
C82 B.n48 VSUBS 0.007087f
C83 B.n49 VSUBS 0.007087f
C84 B.n50 VSUBS 0.007087f
C85 B.n51 VSUBS 0.007087f
C86 B.n52 VSUBS 0.007087f
C87 B.n53 VSUBS 0.007087f
C88 B.n54 VSUBS 0.007087f
C89 B.n55 VSUBS 0.007087f
C90 B.n56 VSUBS 0.007087f
C91 B.n57 VSUBS 0.007087f
C92 B.n58 VSUBS 0.007087f
C93 B.n59 VSUBS 0.007087f
C94 B.n60 VSUBS 0.015768f
C95 B.n61 VSUBS 0.007087f
C96 B.n62 VSUBS 0.007087f
C97 B.n63 VSUBS 0.007087f
C98 B.n64 VSUBS 0.007087f
C99 B.n65 VSUBS 0.007087f
C100 B.n66 VSUBS 0.007087f
C101 B.n67 VSUBS 0.007087f
C102 B.n68 VSUBS 0.007087f
C103 B.n69 VSUBS 0.007087f
C104 B.n70 VSUBS 0.007087f
C105 B.n71 VSUBS 0.007087f
C106 B.n72 VSUBS 0.007087f
C107 B.n73 VSUBS 0.007087f
C108 B.n74 VSUBS 0.007087f
C109 B.n75 VSUBS 0.007087f
C110 B.n76 VSUBS 0.007087f
C111 B.n77 VSUBS 0.007087f
C112 B.n78 VSUBS 0.007087f
C113 B.n79 VSUBS 0.007087f
C114 B.n80 VSUBS 0.007087f
C115 B.n81 VSUBS 0.007087f
C116 B.n82 VSUBS 0.007087f
C117 B.n83 VSUBS 0.007087f
C118 B.n84 VSUBS 0.007087f
C119 B.n85 VSUBS 0.007087f
C120 B.n86 VSUBS 0.007087f
C121 B.n87 VSUBS 0.007087f
C122 B.n88 VSUBS 0.007087f
C123 B.n89 VSUBS 0.007087f
C124 B.n90 VSUBS 0.007087f
C125 B.n91 VSUBS 0.007087f
C126 B.n92 VSUBS 0.007087f
C127 B.n93 VSUBS 0.007087f
C128 B.n94 VSUBS 0.007087f
C129 B.n95 VSUBS 0.007087f
C130 B.n96 VSUBS 0.007087f
C131 B.n97 VSUBS 0.007087f
C132 B.n98 VSUBS 0.007087f
C133 B.n99 VSUBS 0.016622f
C134 B.n100 VSUBS 0.007087f
C135 B.n101 VSUBS 0.007087f
C136 B.n102 VSUBS 0.007087f
C137 B.n103 VSUBS 0.007087f
C138 B.n104 VSUBS 0.007087f
C139 B.n105 VSUBS 0.007087f
C140 B.n106 VSUBS 0.007087f
C141 B.n107 VSUBS 0.007087f
C142 B.n108 VSUBS 0.007087f
C143 B.n109 VSUBS 0.007087f
C144 B.n110 VSUBS 0.007087f
C145 B.n111 VSUBS 0.007087f
C146 B.n112 VSUBS 0.007087f
C147 B.n113 VSUBS 0.007087f
C148 B.t1 VSUBS 0.131481f
C149 B.t2 VSUBS 0.15692f
C150 B.t0 VSUBS 0.836981f
C151 B.n114 VSUBS 0.260232f
C152 B.n115 VSUBS 0.194507f
C153 B.n116 VSUBS 0.016419f
C154 B.n117 VSUBS 0.007087f
C155 B.n118 VSUBS 0.007087f
C156 B.n119 VSUBS 0.007087f
C157 B.n120 VSUBS 0.007087f
C158 B.n121 VSUBS 0.007087f
C159 B.t4 VSUBS 0.131478f
C160 B.t5 VSUBS 0.156918f
C161 B.t3 VSUBS 0.836981f
C162 B.n122 VSUBS 0.260234f
C163 B.n123 VSUBS 0.194509f
C164 B.n124 VSUBS 0.007087f
C165 B.n125 VSUBS 0.007087f
C166 B.n126 VSUBS 0.007087f
C167 B.n127 VSUBS 0.007087f
C168 B.n128 VSUBS 0.007087f
C169 B.n129 VSUBS 0.007087f
C170 B.n130 VSUBS 0.007087f
C171 B.n131 VSUBS 0.007087f
C172 B.n132 VSUBS 0.007087f
C173 B.n133 VSUBS 0.007087f
C174 B.n134 VSUBS 0.007087f
C175 B.n135 VSUBS 0.007087f
C176 B.n136 VSUBS 0.007087f
C177 B.n137 VSUBS 0.007087f
C178 B.n138 VSUBS 0.016622f
C179 B.n139 VSUBS 0.007087f
C180 B.n140 VSUBS 0.007087f
C181 B.n141 VSUBS 0.007087f
C182 B.n142 VSUBS 0.007087f
C183 B.n143 VSUBS 0.007087f
C184 B.n144 VSUBS 0.007087f
C185 B.n145 VSUBS 0.007087f
C186 B.n146 VSUBS 0.007087f
C187 B.n147 VSUBS 0.007087f
C188 B.n148 VSUBS 0.007087f
C189 B.n149 VSUBS 0.007087f
C190 B.n150 VSUBS 0.007087f
C191 B.n151 VSUBS 0.007087f
C192 B.n152 VSUBS 0.007087f
C193 B.n153 VSUBS 0.007087f
C194 B.n154 VSUBS 0.007087f
C195 B.n155 VSUBS 0.007087f
C196 B.n156 VSUBS 0.007087f
C197 B.n157 VSUBS 0.007087f
C198 B.n158 VSUBS 0.007087f
C199 B.n159 VSUBS 0.007087f
C200 B.n160 VSUBS 0.007087f
C201 B.n161 VSUBS 0.007087f
C202 B.n162 VSUBS 0.007087f
C203 B.n163 VSUBS 0.007087f
C204 B.n164 VSUBS 0.007087f
C205 B.n165 VSUBS 0.007087f
C206 B.n166 VSUBS 0.007087f
C207 B.n167 VSUBS 0.007087f
C208 B.n168 VSUBS 0.007087f
C209 B.n169 VSUBS 0.007087f
C210 B.n170 VSUBS 0.007087f
C211 B.n171 VSUBS 0.007087f
C212 B.n172 VSUBS 0.007087f
C213 B.n173 VSUBS 0.007087f
C214 B.n174 VSUBS 0.007087f
C215 B.n175 VSUBS 0.007087f
C216 B.n176 VSUBS 0.007087f
C217 B.n177 VSUBS 0.007087f
C218 B.n178 VSUBS 0.007087f
C219 B.n179 VSUBS 0.007087f
C220 B.n180 VSUBS 0.007087f
C221 B.n181 VSUBS 0.007087f
C222 B.n182 VSUBS 0.007087f
C223 B.n183 VSUBS 0.007087f
C224 B.n184 VSUBS 0.007087f
C225 B.n185 VSUBS 0.007087f
C226 B.n186 VSUBS 0.007087f
C227 B.n187 VSUBS 0.007087f
C228 B.n188 VSUBS 0.007087f
C229 B.n189 VSUBS 0.007087f
C230 B.n190 VSUBS 0.007087f
C231 B.n191 VSUBS 0.007087f
C232 B.n192 VSUBS 0.007087f
C233 B.n193 VSUBS 0.007087f
C234 B.n194 VSUBS 0.007087f
C235 B.n195 VSUBS 0.007087f
C236 B.n196 VSUBS 0.007087f
C237 B.n197 VSUBS 0.007087f
C238 B.n198 VSUBS 0.007087f
C239 B.n199 VSUBS 0.007087f
C240 B.n200 VSUBS 0.007087f
C241 B.n201 VSUBS 0.007087f
C242 B.n202 VSUBS 0.007087f
C243 B.n203 VSUBS 0.007087f
C244 B.n204 VSUBS 0.007087f
C245 B.n205 VSUBS 0.007087f
C246 B.n206 VSUBS 0.007087f
C247 B.n207 VSUBS 0.007087f
C248 B.n208 VSUBS 0.007087f
C249 B.n209 VSUBS 0.007087f
C250 B.n210 VSUBS 0.007087f
C251 B.n211 VSUBS 0.016101f
C252 B.n212 VSUBS 0.016101f
C253 B.n213 VSUBS 0.016622f
C254 B.n214 VSUBS 0.007087f
C255 B.n215 VSUBS 0.007087f
C256 B.n216 VSUBS 0.007087f
C257 B.n217 VSUBS 0.007087f
C258 B.n218 VSUBS 0.007087f
C259 B.n219 VSUBS 0.007087f
C260 B.n220 VSUBS 0.007087f
C261 B.n221 VSUBS 0.007087f
C262 B.n222 VSUBS 0.007087f
C263 B.n223 VSUBS 0.007087f
C264 B.n224 VSUBS 0.007087f
C265 B.n225 VSUBS 0.007087f
C266 B.n226 VSUBS 0.007087f
C267 B.n227 VSUBS 0.007087f
C268 B.n228 VSUBS 0.007087f
C269 B.n229 VSUBS 0.007087f
C270 B.n230 VSUBS 0.007087f
C271 B.n231 VSUBS 0.007087f
C272 B.n232 VSUBS 0.007087f
C273 B.n233 VSUBS 0.007087f
C274 B.n234 VSUBS 0.007087f
C275 B.n235 VSUBS 0.007087f
C276 B.n236 VSUBS 0.007087f
C277 B.n237 VSUBS 0.007087f
C278 B.n238 VSUBS 0.007087f
C279 B.n239 VSUBS 0.007087f
C280 B.n240 VSUBS 0.007087f
C281 B.n241 VSUBS 0.007087f
C282 B.n242 VSUBS 0.007087f
C283 B.n243 VSUBS 0.007087f
C284 B.n244 VSUBS 0.007087f
C285 B.n245 VSUBS 0.007087f
C286 B.n246 VSUBS 0.007087f
C287 B.n247 VSUBS 0.007087f
C288 B.n248 VSUBS 0.007087f
C289 B.n249 VSUBS 0.007087f
C290 B.n250 VSUBS 0.007087f
C291 B.n251 VSUBS 0.007087f
C292 B.n252 VSUBS 0.007087f
C293 B.n253 VSUBS 0.007087f
C294 B.n254 VSUBS 0.007087f
C295 B.n255 VSUBS 0.007087f
C296 B.n256 VSUBS 0.007087f
C297 B.n257 VSUBS 0.00667f
C298 B.n258 VSUBS 0.016419f
C299 B.n259 VSUBS 0.00396f
C300 B.n260 VSUBS 0.007087f
C301 B.n261 VSUBS 0.007087f
C302 B.n262 VSUBS 0.007087f
C303 B.n263 VSUBS 0.007087f
C304 B.n264 VSUBS 0.007087f
C305 B.n265 VSUBS 0.007087f
C306 B.n266 VSUBS 0.007087f
C307 B.n267 VSUBS 0.007087f
C308 B.n268 VSUBS 0.007087f
C309 B.n269 VSUBS 0.007087f
C310 B.n270 VSUBS 0.007087f
C311 B.n271 VSUBS 0.007087f
C312 B.n272 VSUBS 0.00396f
C313 B.n273 VSUBS 0.007087f
C314 B.n274 VSUBS 0.007087f
C315 B.n275 VSUBS 0.00667f
C316 B.n276 VSUBS 0.007087f
C317 B.n277 VSUBS 0.007087f
C318 B.n278 VSUBS 0.007087f
C319 B.n279 VSUBS 0.007087f
C320 B.n280 VSUBS 0.007087f
C321 B.n281 VSUBS 0.007087f
C322 B.n282 VSUBS 0.007087f
C323 B.n283 VSUBS 0.007087f
C324 B.n284 VSUBS 0.007087f
C325 B.n285 VSUBS 0.007087f
C326 B.n286 VSUBS 0.007087f
C327 B.n287 VSUBS 0.007087f
C328 B.n288 VSUBS 0.007087f
C329 B.n289 VSUBS 0.007087f
C330 B.n290 VSUBS 0.007087f
C331 B.n291 VSUBS 0.007087f
C332 B.n292 VSUBS 0.007087f
C333 B.n293 VSUBS 0.007087f
C334 B.n294 VSUBS 0.007087f
C335 B.n295 VSUBS 0.007087f
C336 B.n296 VSUBS 0.007087f
C337 B.n297 VSUBS 0.007087f
C338 B.n298 VSUBS 0.007087f
C339 B.n299 VSUBS 0.007087f
C340 B.n300 VSUBS 0.007087f
C341 B.n301 VSUBS 0.007087f
C342 B.n302 VSUBS 0.007087f
C343 B.n303 VSUBS 0.007087f
C344 B.n304 VSUBS 0.007087f
C345 B.n305 VSUBS 0.007087f
C346 B.n306 VSUBS 0.007087f
C347 B.n307 VSUBS 0.007087f
C348 B.n308 VSUBS 0.007087f
C349 B.n309 VSUBS 0.007087f
C350 B.n310 VSUBS 0.007087f
C351 B.n311 VSUBS 0.007087f
C352 B.n312 VSUBS 0.007087f
C353 B.n313 VSUBS 0.007087f
C354 B.n314 VSUBS 0.007087f
C355 B.n315 VSUBS 0.007087f
C356 B.n316 VSUBS 0.007087f
C357 B.n317 VSUBS 0.007087f
C358 B.n318 VSUBS 0.016622f
C359 B.n319 VSUBS 0.016101f
C360 B.n320 VSUBS 0.016101f
C361 B.n321 VSUBS 0.007087f
C362 B.n322 VSUBS 0.007087f
C363 B.n323 VSUBS 0.007087f
C364 B.n324 VSUBS 0.007087f
C365 B.n325 VSUBS 0.007087f
C366 B.n326 VSUBS 0.007087f
C367 B.n327 VSUBS 0.007087f
C368 B.n328 VSUBS 0.007087f
C369 B.n329 VSUBS 0.007087f
C370 B.n330 VSUBS 0.007087f
C371 B.n331 VSUBS 0.007087f
C372 B.n332 VSUBS 0.007087f
C373 B.n333 VSUBS 0.007087f
C374 B.n334 VSUBS 0.007087f
C375 B.n335 VSUBS 0.007087f
C376 B.n336 VSUBS 0.007087f
C377 B.n337 VSUBS 0.007087f
C378 B.n338 VSUBS 0.007087f
C379 B.n339 VSUBS 0.007087f
C380 B.n340 VSUBS 0.007087f
C381 B.n341 VSUBS 0.007087f
C382 B.n342 VSUBS 0.007087f
C383 B.n343 VSUBS 0.007087f
C384 B.n344 VSUBS 0.007087f
C385 B.n345 VSUBS 0.007087f
C386 B.n346 VSUBS 0.007087f
C387 B.n347 VSUBS 0.007087f
C388 B.n348 VSUBS 0.007087f
C389 B.n349 VSUBS 0.007087f
C390 B.n350 VSUBS 0.007087f
C391 B.n351 VSUBS 0.007087f
C392 B.n352 VSUBS 0.007087f
C393 B.n353 VSUBS 0.007087f
C394 B.n354 VSUBS 0.007087f
C395 B.n355 VSUBS 0.007087f
C396 B.n356 VSUBS 0.007087f
C397 B.n357 VSUBS 0.007087f
C398 B.n358 VSUBS 0.007087f
C399 B.n359 VSUBS 0.007087f
C400 B.n360 VSUBS 0.007087f
C401 B.n361 VSUBS 0.007087f
C402 B.n362 VSUBS 0.007087f
C403 B.n363 VSUBS 0.007087f
C404 B.n364 VSUBS 0.007087f
C405 B.n365 VSUBS 0.007087f
C406 B.n366 VSUBS 0.007087f
C407 B.n367 VSUBS 0.007087f
C408 B.n368 VSUBS 0.007087f
C409 B.n369 VSUBS 0.007087f
C410 B.n370 VSUBS 0.007087f
C411 B.n371 VSUBS 0.007087f
C412 B.n372 VSUBS 0.007087f
C413 B.n373 VSUBS 0.007087f
C414 B.n374 VSUBS 0.007087f
C415 B.n375 VSUBS 0.007087f
C416 B.n376 VSUBS 0.007087f
C417 B.n377 VSUBS 0.007087f
C418 B.n378 VSUBS 0.007087f
C419 B.n379 VSUBS 0.007087f
C420 B.n380 VSUBS 0.007087f
C421 B.n381 VSUBS 0.007087f
C422 B.n382 VSUBS 0.007087f
C423 B.n383 VSUBS 0.007087f
C424 B.n384 VSUBS 0.007087f
C425 B.n385 VSUBS 0.007087f
C426 B.n386 VSUBS 0.007087f
C427 B.n387 VSUBS 0.007087f
C428 B.n388 VSUBS 0.007087f
C429 B.n389 VSUBS 0.007087f
C430 B.n390 VSUBS 0.007087f
C431 B.n391 VSUBS 0.007087f
C432 B.n392 VSUBS 0.007087f
C433 B.n393 VSUBS 0.007087f
C434 B.n394 VSUBS 0.007087f
C435 B.n395 VSUBS 0.007087f
C436 B.n396 VSUBS 0.007087f
C437 B.n397 VSUBS 0.007087f
C438 B.n398 VSUBS 0.007087f
C439 B.n399 VSUBS 0.007087f
C440 B.n400 VSUBS 0.007087f
C441 B.n401 VSUBS 0.007087f
C442 B.n402 VSUBS 0.007087f
C443 B.n403 VSUBS 0.007087f
C444 B.n404 VSUBS 0.007087f
C445 B.n405 VSUBS 0.007087f
C446 B.n406 VSUBS 0.007087f
C447 B.n407 VSUBS 0.007087f
C448 B.n408 VSUBS 0.007087f
C449 B.n409 VSUBS 0.007087f
C450 B.n410 VSUBS 0.007087f
C451 B.n411 VSUBS 0.007087f
C452 B.n412 VSUBS 0.007087f
C453 B.n413 VSUBS 0.007087f
C454 B.n414 VSUBS 0.007087f
C455 B.n415 VSUBS 0.007087f
C456 B.n416 VSUBS 0.007087f
C457 B.n417 VSUBS 0.007087f
C458 B.n418 VSUBS 0.007087f
C459 B.n419 VSUBS 0.007087f
C460 B.n420 VSUBS 0.007087f
C461 B.n421 VSUBS 0.007087f
C462 B.n422 VSUBS 0.007087f
C463 B.n423 VSUBS 0.007087f
C464 B.n424 VSUBS 0.007087f
C465 B.n425 VSUBS 0.007087f
C466 B.n426 VSUBS 0.007087f
C467 B.n427 VSUBS 0.007087f
C468 B.n428 VSUBS 0.007087f
C469 B.n429 VSUBS 0.007087f
C470 B.n430 VSUBS 0.007087f
C471 B.n431 VSUBS 0.007087f
C472 B.n432 VSUBS 0.007087f
C473 B.n433 VSUBS 0.016956f
C474 B.n434 VSUBS 0.016101f
C475 B.n435 VSUBS 0.016622f
C476 B.n436 VSUBS 0.007087f
C477 B.n437 VSUBS 0.007087f
C478 B.n438 VSUBS 0.007087f
C479 B.n439 VSUBS 0.007087f
C480 B.n440 VSUBS 0.007087f
C481 B.n441 VSUBS 0.007087f
C482 B.n442 VSUBS 0.007087f
C483 B.n443 VSUBS 0.007087f
C484 B.n444 VSUBS 0.007087f
C485 B.n445 VSUBS 0.007087f
C486 B.n446 VSUBS 0.007087f
C487 B.n447 VSUBS 0.007087f
C488 B.n448 VSUBS 0.007087f
C489 B.n449 VSUBS 0.007087f
C490 B.n450 VSUBS 0.007087f
C491 B.n451 VSUBS 0.007087f
C492 B.n452 VSUBS 0.007087f
C493 B.n453 VSUBS 0.007087f
C494 B.n454 VSUBS 0.007087f
C495 B.n455 VSUBS 0.007087f
C496 B.n456 VSUBS 0.007087f
C497 B.n457 VSUBS 0.007087f
C498 B.n458 VSUBS 0.007087f
C499 B.n459 VSUBS 0.007087f
C500 B.n460 VSUBS 0.007087f
C501 B.n461 VSUBS 0.007087f
C502 B.n462 VSUBS 0.007087f
C503 B.n463 VSUBS 0.007087f
C504 B.n464 VSUBS 0.007087f
C505 B.n465 VSUBS 0.007087f
C506 B.n466 VSUBS 0.007087f
C507 B.n467 VSUBS 0.007087f
C508 B.n468 VSUBS 0.007087f
C509 B.n469 VSUBS 0.007087f
C510 B.n470 VSUBS 0.007087f
C511 B.n471 VSUBS 0.007087f
C512 B.n472 VSUBS 0.007087f
C513 B.n473 VSUBS 0.007087f
C514 B.n474 VSUBS 0.007087f
C515 B.n475 VSUBS 0.007087f
C516 B.n476 VSUBS 0.007087f
C517 B.n477 VSUBS 0.007087f
C518 B.n478 VSUBS 0.007087f
C519 B.n479 VSUBS 0.00667f
C520 B.n480 VSUBS 0.016419f
C521 B.n481 VSUBS 0.00396f
C522 B.n482 VSUBS 0.007087f
C523 B.n483 VSUBS 0.007087f
C524 B.n484 VSUBS 0.007087f
C525 B.n485 VSUBS 0.007087f
C526 B.n486 VSUBS 0.007087f
C527 B.n487 VSUBS 0.007087f
C528 B.n488 VSUBS 0.007087f
C529 B.n489 VSUBS 0.007087f
C530 B.n490 VSUBS 0.007087f
C531 B.n491 VSUBS 0.007087f
C532 B.n492 VSUBS 0.007087f
C533 B.n493 VSUBS 0.007087f
C534 B.n494 VSUBS 0.00396f
C535 B.n495 VSUBS 0.007087f
C536 B.n496 VSUBS 0.007087f
C537 B.n497 VSUBS 0.00667f
C538 B.n498 VSUBS 0.007087f
C539 B.n499 VSUBS 0.007087f
C540 B.n500 VSUBS 0.007087f
C541 B.n501 VSUBS 0.007087f
C542 B.n502 VSUBS 0.007087f
C543 B.n503 VSUBS 0.007087f
C544 B.n504 VSUBS 0.007087f
C545 B.n505 VSUBS 0.007087f
C546 B.n506 VSUBS 0.007087f
C547 B.n507 VSUBS 0.007087f
C548 B.n508 VSUBS 0.007087f
C549 B.n509 VSUBS 0.007087f
C550 B.n510 VSUBS 0.007087f
C551 B.n511 VSUBS 0.007087f
C552 B.n512 VSUBS 0.007087f
C553 B.n513 VSUBS 0.007087f
C554 B.n514 VSUBS 0.007087f
C555 B.n515 VSUBS 0.007087f
C556 B.n516 VSUBS 0.007087f
C557 B.n517 VSUBS 0.007087f
C558 B.n518 VSUBS 0.007087f
C559 B.n519 VSUBS 0.007087f
C560 B.n520 VSUBS 0.007087f
C561 B.n521 VSUBS 0.007087f
C562 B.n522 VSUBS 0.007087f
C563 B.n523 VSUBS 0.007087f
C564 B.n524 VSUBS 0.007087f
C565 B.n525 VSUBS 0.007087f
C566 B.n526 VSUBS 0.007087f
C567 B.n527 VSUBS 0.007087f
C568 B.n528 VSUBS 0.007087f
C569 B.n529 VSUBS 0.007087f
C570 B.n530 VSUBS 0.007087f
C571 B.n531 VSUBS 0.007087f
C572 B.n532 VSUBS 0.007087f
C573 B.n533 VSUBS 0.007087f
C574 B.n534 VSUBS 0.007087f
C575 B.n535 VSUBS 0.007087f
C576 B.n536 VSUBS 0.007087f
C577 B.n537 VSUBS 0.007087f
C578 B.n538 VSUBS 0.007087f
C579 B.n539 VSUBS 0.007087f
C580 B.n540 VSUBS 0.016622f
C581 B.n541 VSUBS 0.016101f
C582 B.n542 VSUBS 0.016101f
C583 B.n543 VSUBS 0.007087f
C584 B.n544 VSUBS 0.007087f
C585 B.n545 VSUBS 0.007087f
C586 B.n546 VSUBS 0.007087f
C587 B.n547 VSUBS 0.007087f
C588 B.n548 VSUBS 0.007087f
C589 B.n549 VSUBS 0.007087f
C590 B.n550 VSUBS 0.007087f
C591 B.n551 VSUBS 0.007087f
C592 B.n552 VSUBS 0.007087f
C593 B.n553 VSUBS 0.007087f
C594 B.n554 VSUBS 0.007087f
C595 B.n555 VSUBS 0.007087f
C596 B.n556 VSUBS 0.007087f
C597 B.n557 VSUBS 0.007087f
C598 B.n558 VSUBS 0.007087f
C599 B.n559 VSUBS 0.007087f
C600 B.n560 VSUBS 0.007087f
C601 B.n561 VSUBS 0.007087f
C602 B.n562 VSUBS 0.007087f
C603 B.n563 VSUBS 0.007087f
C604 B.n564 VSUBS 0.007087f
C605 B.n565 VSUBS 0.007087f
C606 B.n566 VSUBS 0.007087f
C607 B.n567 VSUBS 0.007087f
C608 B.n568 VSUBS 0.007087f
C609 B.n569 VSUBS 0.007087f
C610 B.n570 VSUBS 0.007087f
C611 B.n571 VSUBS 0.007087f
C612 B.n572 VSUBS 0.007087f
C613 B.n573 VSUBS 0.007087f
C614 B.n574 VSUBS 0.007087f
C615 B.n575 VSUBS 0.007087f
C616 B.n576 VSUBS 0.007087f
C617 B.n577 VSUBS 0.007087f
C618 B.n578 VSUBS 0.007087f
C619 B.n579 VSUBS 0.007087f
C620 B.n580 VSUBS 0.007087f
C621 B.n581 VSUBS 0.007087f
C622 B.n582 VSUBS 0.007087f
C623 B.n583 VSUBS 0.007087f
C624 B.n584 VSUBS 0.007087f
C625 B.n585 VSUBS 0.007087f
C626 B.n586 VSUBS 0.007087f
C627 B.n587 VSUBS 0.007087f
C628 B.n588 VSUBS 0.007087f
C629 B.n589 VSUBS 0.007087f
C630 B.n590 VSUBS 0.007087f
C631 B.n591 VSUBS 0.007087f
C632 B.n592 VSUBS 0.007087f
C633 B.n593 VSUBS 0.007087f
C634 B.n594 VSUBS 0.007087f
C635 B.n595 VSUBS 0.007087f
C636 B.n596 VSUBS 0.007087f
C637 B.n597 VSUBS 0.007087f
C638 B.n598 VSUBS 0.007087f
C639 B.n599 VSUBS 0.016046f
C640 VDD1.n0 VSUBS 0.025013f
C641 VDD1.n1 VSUBS 0.021917f
C642 VDD1.n2 VSUBS 0.011777f
C643 VDD1.n3 VSUBS 0.027837f
C644 VDD1.n4 VSUBS 0.01247f
C645 VDD1.n5 VSUBS 0.021917f
C646 VDD1.n6 VSUBS 0.011777f
C647 VDD1.n7 VSUBS 0.027837f
C648 VDD1.n8 VSUBS 0.01247f
C649 VDD1.n9 VSUBS 0.021917f
C650 VDD1.n10 VSUBS 0.011777f
C651 VDD1.n11 VSUBS 0.027837f
C652 VDD1.n12 VSUBS 0.01247f
C653 VDD1.n13 VSUBS 0.11037f
C654 VDD1.t4 VSUBS 0.059378f
C655 VDD1.n14 VSUBS 0.020878f
C656 VDD1.n15 VSUBS 0.017708f
C657 VDD1.n16 VSUBS 0.011777f
C658 VDD1.n17 VSUBS 0.717579f
C659 VDD1.n18 VSUBS 0.021917f
C660 VDD1.n19 VSUBS 0.011777f
C661 VDD1.n20 VSUBS 0.01247f
C662 VDD1.n21 VSUBS 0.027837f
C663 VDD1.n22 VSUBS 0.027837f
C664 VDD1.n23 VSUBS 0.01247f
C665 VDD1.n24 VSUBS 0.011777f
C666 VDD1.n25 VSUBS 0.021917f
C667 VDD1.n26 VSUBS 0.021917f
C668 VDD1.n27 VSUBS 0.011777f
C669 VDD1.n28 VSUBS 0.01247f
C670 VDD1.n29 VSUBS 0.027837f
C671 VDD1.n30 VSUBS 0.027837f
C672 VDD1.n31 VSUBS 0.01247f
C673 VDD1.n32 VSUBS 0.011777f
C674 VDD1.n33 VSUBS 0.021917f
C675 VDD1.n34 VSUBS 0.021917f
C676 VDD1.n35 VSUBS 0.011777f
C677 VDD1.n36 VSUBS 0.01247f
C678 VDD1.n37 VSUBS 0.027837f
C679 VDD1.n38 VSUBS 0.07056f
C680 VDD1.n39 VSUBS 0.01247f
C681 VDD1.n40 VSUBS 0.011777f
C682 VDD1.n41 VSUBS 0.050361f
C683 VDD1.n42 VSUBS 0.056188f
C684 VDD1.n43 VSUBS 0.025013f
C685 VDD1.n44 VSUBS 0.021917f
C686 VDD1.n45 VSUBS 0.011777f
C687 VDD1.n46 VSUBS 0.027837f
C688 VDD1.n47 VSUBS 0.01247f
C689 VDD1.n48 VSUBS 0.021917f
C690 VDD1.n49 VSUBS 0.011777f
C691 VDD1.n50 VSUBS 0.027837f
C692 VDD1.n51 VSUBS 0.01247f
C693 VDD1.n52 VSUBS 0.021917f
C694 VDD1.n53 VSUBS 0.011777f
C695 VDD1.n54 VSUBS 0.027837f
C696 VDD1.n55 VSUBS 0.01247f
C697 VDD1.n56 VSUBS 0.11037f
C698 VDD1.t5 VSUBS 0.059378f
C699 VDD1.n57 VSUBS 0.020878f
C700 VDD1.n58 VSUBS 0.017708f
C701 VDD1.n59 VSUBS 0.011777f
C702 VDD1.n60 VSUBS 0.717579f
C703 VDD1.n61 VSUBS 0.021917f
C704 VDD1.n62 VSUBS 0.011777f
C705 VDD1.n63 VSUBS 0.01247f
C706 VDD1.n64 VSUBS 0.027837f
C707 VDD1.n65 VSUBS 0.027837f
C708 VDD1.n66 VSUBS 0.01247f
C709 VDD1.n67 VSUBS 0.011777f
C710 VDD1.n68 VSUBS 0.021917f
C711 VDD1.n69 VSUBS 0.021917f
C712 VDD1.n70 VSUBS 0.011777f
C713 VDD1.n71 VSUBS 0.01247f
C714 VDD1.n72 VSUBS 0.027837f
C715 VDD1.n73 VSUBS 0.027837f
C716 VDD1.n74 VSUBS 0.01247f
C717 VDD1.n75 VSUBS 0.011777f
C718 VDD1.n76 VSUBS 0.021917f
C719 VDD1.n77 VSUBS 0.021917f
C720 VDD1.n78 VSUBS 0.011777f
C721 VDD1.n79 VSUBS 0.01247f
C722 VDD1.n80 VSUBS 0.027837f
C723 VDD1.n81 VSUBS 0.07056f
C724 VDD1.n82 VSUBS 0.01247f
C725 VDD1.n83 VSUBS 0.011777f
C726 VDD1.n84 VSUBS 0.050361f
C727 VDD1.n85 VSUBS 0.055593f
C728 VDD1.t1 VSUBS 0.141154f
C729 VDD1.t0 VSUBS 0.141154f
C730 VDD1.n86 VSUBS 1.01409f
C731 VDD1.n87 VSUBS 2.29514f
C732 VDD1.t2 VSUBS 0.141154f
C733 VDD1.t3 VSUBS 0.141154f
C734 VDD1.n88 VSUBS 1.01064f
C735 VDD1.n89 VSUBS 2.29371f
C736 VP.n0 VSUBS 0.050448f
C737 VP.t5 VSUBS 1.84407f
C738 VP.n1 VSUBS 0.031045f
C739 VP.n2 VSUBS 0.038264f
C740 VP.t4 VSUBS 1.84407f
C741 VP.n3 VSUBS 0.076571f
C742 VP.n4 VSUBS 0.038264f
C743 VP.t0 VSUBS 1.84407f
C744 VP.n5 VSUBS 0.791175f
C745 VP.n6 VSUBS 0.050448f
C746 VP.t2 VSUBS 1.84407f
C747 VP.n7 VSUBS 0.031045f
C748 VP.n8 VSUBS 0.325715f
C749 VP.t3 VSUBS 1.84407f
C750 VP.t1 VSUBS 2.07882f
C751 VP.n9 VSUBS 0.762975f
C752 VP.n10 VSUBS 0.774831f
C753 VP.n11 VSUBS 0.053711f
C754 VP.n12 VSUBS 0.076571f
C755 VP.n13 VSUBS 0.038264f
C756 VP.n14 VSUBS 0.038264f
C757 VP.n15 VSUBS 0.038264f
C758 VP.n16 VSUBS 0.075424f
C759 VP.n17 VSUBS 0.055823f
C760 VP.n18 VSUBS 0.791175f
C761 VP.n19 VSUBS 1.75495f
C762 VP.n20 VSUBS 1.78609f
C763 VP.n21 VSUBS 0.050448f
C764 VP.n22 VSUBS 0.055823f
C765 VP.n23 VSUBS 0.075424f
C766 VP.n24 VSUBS 0.031045f
C767 VP.n25 VSUBS 0.038264f
C768 VP.n26 VSUBS 0.038264f
C769 VP.n27 VSUBS 0.038264f
C770 VP.n28 VSUBS 0.053711f
C771 VP.n29 VSUBS 0.676113f
C772 VP.n30 VSUBS 0.053711f
C773 VP.n31 VSUBS 0.076571f
C774 VP.n32 VSUBS 0.038264f
C775 VP.n33 VSUBS 0.038264f
C776 VP.n34 VSUBS 0.038264f
C777 VP.n35 VSUBS 0.075424f
C778 VP.n36 VSUBS 0.055823f
C779 VP.n37 VSUBS 0.791175f
C780 VP.n38 VSUBS 0.054296f
C781 VTAIL.t6 VSUBS 0.197963f
C782 VTAIL.t7 VSUBS 0.197963f
C783 VTAIL.n0 VSUBS 1.28107f
C784 VTAIL.n1 VSUBS 0.853317f
C785 VTAIL.n2 VSUBS 0.035079f
C786 VTAIL.n3 VSUBS 0.030738f
C787 VTAIL.n4 VSUBS 0.016517f
C788 VTAIL.n5 VSUBS 0.03904f
C789 VTAIL.n6 VSUBS 0.017489f
C790 VTAIL.n7 VSUBS 0.030738f
C791 VTAIL.n8 VSUBS 0.016517f
C792 VTAIL.n9 VSUBS 0.03904f
C793 VTAIL.n10 VSUBS 0.017489f
C794 VTAIL.n11 VSUBS 0.030738f
C795 VTAIL.n12 VSUBS 0.016517f
C796 VTAIL.n13 VSUBS 0.03904f
C797 VTAIL.n14 VSUBS 0.017489f
C798 VTAIL.n15 VSUBS 0.154789f
C799 VTAIL.t5 VSUBS 0.083276f
C800 VTAIL.n16 VSUBS 0.02928f
C801 VTAIL.n17 VSUBS 0.024835f
C802 VTAIL.n18 VSUBS 0.016517f
C803 VTAIL.n19 VSUBS 1.00637f
C804 VTAIL.n20 VSUBS 0.030738f
C805 VTAIL.n21 VSUBS 0.016517f
C806 VTAIL.n22 VSUBS 0.017489f
C807 VTAIL.n23 VSUBS 0.03904f
C808 VTAIL.n24 VSUBS 0.03904f
C809 VTAIL.n25 VSUBS 0.017489f
C810 VTAIL.n26 VSUBS 0.016517f
C811 VTAIL.n27 VSUBS 0.030738f
C812 VTAIL.n28 VSUBS 0.030738f
C813 VTAIL.n29 VSUBS 0.016517f
C814 VTAIL.n30 VSUBS 0.017489f
C815 VTAIL.n31 VSUBS 0.03904f
C816 VTAIL.n32 VSUBS 0.03904f
C817 VTAIL.n33 VSUBS 0.017489f
C818 VTAIL.n34 VSUBS 0.016517f
C819 VTAIL.n35 VSUBS 0.030738f
C820 VTAIL.n36 VSUBS 0.030738f
C821 VTAIL.n37 VSUBS 0.016517f
C822 VTAIL.n38 VSUBS 0.017489f
C823 VTAIL.n39 VSUBS 0.03904f
C824 VTAIL.n40 VSUBS 0.098957f
C825 VTAIL.n41 VSUBS 0.017489f
C826 VTAIL.n42 VSUBS 0.016517f
C827 VTAIL.n43 VSUBS 0.070629f
C828 VTAIL.n44 VSUBS 0.049949f
C829 VTAIL.n45 VSUBS 0.396576f
C830 VTAIL.t2 VSUBS 0.197963f
C831 VTAIL.t1 VSUBS 0.197963f
C832 VTAIL.n46 VSUBS 1.28107f
C833 VTAIL.n47 VSUBS 2.40047f
C834 VTAIL.t8 VSUBS 0.197963f
C835 VTAIL.t11 VSUBS 0.197963f
C836 VTAIL.n48 VSUBS 1.28108f
C837 VTAIL.n49 VSUBS 2.40046f
C838 VTAIL.n50 VSUBS 0.035079f
C839 VTAIL.n51 VSUBS 0.030738f
C840 VTAIL.n52 VSUBS 0.016517f
C841 VTAIL.n53 VSUBS 0.03904f
C842 VTAIL.n54 VSUBS 0.017489f
C843 VTAIL.n55 VSUBS 0.030738f
C844 VTAIL.n56 VSUBS 0.016517f
C845 VTAIL.n57 VSUBS 0.03904f
C846 VTAIL.n58 VSUBS 0.017489f
C847 VTAIL.n59 VSUBS 0.030738f
C848 VTAIL.n60 VSUBS 0.016517f
C849 VTAIL.n61 VSUBS 0.03904f
C850 VTAIL.n62 VSUBS 0.017489f
C851 VTAIL.n63 VSUBS 0.154789f
C852 VTAIL.t9 VSUBS 0.083276f
C853 VTAIL.n64 VSUBS 0.02928f
C854 VTAIL.n65 VSUBS 0.024835f
C855 VTAIL.n66 VSUBS 0.016517f
C856 VTAIL.n67 VSUBS 1.00637f
C857 VTAIL.n68 VSUBS 0.030738f
C858 VTAIL.n69 VSUBS 0.016517f
C859 VTAIL.n70 VSUBS 0.017489f
C860 VTAIL.n71 VSUBS 0.03904f
C861 VTAIL.n72 VSUBS 0.03904f
C862 VTAIL.n73 VSUBS 0.017489f
C863 VTAIL.n74 VSUBS 0.016517f
C864 VTAIL.n75 VSUBS 0.030738f
C865 VTAIL.n76 VSUBS 0.030738f
C866 VTAIL.n77 VSUBS 0.016517f
C867 VTAIL.n78 VSUBS 0.017489f
C868 VTAIL.n79 VSUBS 0.03904f
C869 VTAIL.n80 VSUBS 0.03904f
C870 VTAIL.n81 VSUBS 0.017489f
C871 VTAIL.n82 VSUBS 0.016517f
C872 VTAIL.n83 VSUBS 0.030738f
C873 VTAIL.n84 VSUBS 0.030738f
C874 VTAIL.n85 VSUBS 0.016517f
C875 VTAIL.n86 VSUBS 0.017489f
C876 VTAIL.n87 VSUBS 0.03904f
C877 VTAIL.n88 VSUBS 0.098957f
C878 VTAIL.n89 VSUBS 0.017489f
C879 VTAIL.n90 VSUBS 0.016517f
C880 VTAIL.n91 VSUBS 0.070629f
C881 VTAIL.n92 VSUBS 0.049949f
C882 VTAIL.n93 VSUBS 0.396576f
C883 VTAIL.t4 VSUBS 0.197963f
C884 VTAIL.t3 VSUBS 0.197963f
C885 VTAIL.n94 VSUBS 1.28108f
C886 VTAIL.n95 VSUBS 1.00956f
C887 VTAIL.n96 VSUBS 0.035079f
C888 VTAIL.n97 VSUBS 0.030738f
C889 VTAIL.n98 VSUBS 0.016517f
C890 VTAIL.n99 VSUBS 0.03904f
C891 VTAIL.n100 VSUBS 0.017489f
C892 VTAIL.n101 VSUBS 0.030738f
C893 VTAIL.n102 VSUBS 0.016517f
C894 VTAIL.n103 VSUBS 0.03904f
C895 VTAIL.n104 VSUBS 0.017489f
C896 VTAIL.n105 VSUBS 0.030738f
C897 VTAIL.n106 VSUBS 0.016517f
C898 VTAIL.n107 VSUBS 0.03904f
C899 VTAIL.n108 VSUBS 0.017489f
C900 VTAIL.n109 VSUBS 0.154789f
C901 VTAIL.t0 VSUBS 0.083276f
C902 VTAIL.n110 VSUBS 0.02928f
C903 VTAIL.n111 VSUBS 0.024835f
C904 VTAIL.n112 VSUBS 0.016517f
C905 VTAIL.n113 VSUBS 1.00637f
C906 VTAIL.n114 VSUBS 0.030738f
C907 VTAIL.n115 VSUBS 0.016517f
C908 VTAIL.n116 VSUBS 0.017489f
C909 VTAIL.n117 VSUBS 0.03904f
C910 VTAIL.n118 VSUBS 0.03904f
C911 VTAIL.n119 VSUBS 0.017489f
C912 VTAIL.n120 VSUBS 0.016517f
C913 VTAIL.n121 VSUBS 0.030738f
C914 VTAIL.n122 VSUBS 0.030738f
C915 VTAIL.n123 VSUBS 0.016517f
C916 VTAIL.n124 VSUBS 0.017489f
C917 VTAIL.n125 VSUBS 0.03904f
C918 VTAIL.n126 VSUBS 0.03904f
C919 VTAIL.n127 VSUBS 0.017489f
C920 VTAIL.n128 VSUBS 0.016517f
C921 VTAIL.n129 VSUBS 0.030738f
C922 VTAIL.n130 VSUBS 0.030738f
C923 VTAIL.n131 VSUBS 0.016517f
C924 VTAIL.n132 VSUBS 0.017489f
C925 VTAIL.n133 VSUBS 0.03904f
C926 VTAIL.n134 VSUBS 0.098957f
C927 VTAIL.n135 VSUBS 0.017489f
C928 VTAIL.n136 VSUBS 0.016517f
C929 VTAIL.n137 VSUBS 0.070629f
C930 VTAIL.n138 VSUBS 0.049949f
C931 VTAIL.n139 VSUBS 1.57146f
C932 VTAIL.n140 VSUBS 0.035079f
C933 VTAIL.n141 VSUBS 0.030738f
C934 VTAIL.n142 VSUBS 0.016517f
C935 VTAIL.n143 VSUBS 0.03904f
C936 VTAIL.n144 VSUBS 0.017489f
C937 VTAIL.n145 VSUBS 0.030738f
C938 VTAIL.n146 VSUBS 0.016517f
C939 VTAIL.n147 VSUBS 0.03904f
C940 VTAIL.n148 VSUBS 0.017489f
C941 VTAIL.n149 VSUBS 0.030738f
C942 VTAIL.n150 VSUBS 0.016517f
C943 VTAIL.n151 VSUBS 0.03904f
C944 VTAIL.n152 VSUBS 0.017489f
C945 VTAIL.n153 VSUBS 0.154789f
C946 VTAIL.t10 VSUBS 0.083276f
C947 VTAIL.n154 VSUBS 0.02928f
C948 VTAIL.n155 VSUBS 0.024835f
C949 VTAIL.n156 VSUBS 0.016517f
C950 VTAIL.n157 VSUBS 1.00637f
C951 VTAIL.n158 VSUBS 0.030738f
C952 VTAIL.n159 VSUBS 0.016517f
C953 VTAIL.n160 VSUBS 0.017489f
C954 VTAIL.n161 VSUBS 0.03904f
C955 VTAIL.n162 VSUBS 0.03904f
C956 VTAIL.n163 VSUBS 0.017489f
C957 VTAIL.n164 VSUBS 0.016517f
C958 VTAIL.n165 VSUBS 0.030738f
C959 VTAIL.n166 VSUBS 0.030738f
C960 VTAIL.n167 VSUBS 0.016517f
C961 VTAIL.n168 VSUBS 0.017489f
C962 VTAIL.n169 VSUBS 0.03904f
C963 VTAIL.n170 VSUBS 0.03904f
C964 VTAIL.n171 VSUBS 0.017489f
C965 VTAIL.n172 VSUBS 0.016517f
C966 VTAIL.n173 VSUBS 0.030738f
C967 VTAIL.n174 VSUBS 0.030738f
C968 VTAIL.n175 VSUBS 0.016517f
C969 VTAIL.n176 VSUBS 0.017489f
C970 VTAIL.n177 VSUBS 0.03904f
C971 VTAIL.n178 VSUBS 0.098957f
C972 VTAIL.n179 VSUBS 0.017489f
C973 VTAIL.n180 VSUBS 0.016517f
C974 VTAIL.n181 VSUBS 0.070629f
C975 VTAIL.n182 VSUBS 0.049949f
C976 VTAIL.n183 VSUBS 1.51169f
C977 VDD2.n0 VSUBS 0.02474f
C978 VDD2.n1 VSUBS 0.021678f
C979 VDD2.n2 VSUBS 0.011649f
C980 VDD2.n3 VSUBS 0.027534f
C981 VDD2.n4 VSUBS 0.012334f
C982 VDD2.n5 VSUBS 0.021678f
C983 VDD2.n6 VSUBS 0.011649f
C984 VDD2.n7 VSUBS 0.027534f
C985 VDD2.n8 VSUBS 0.012334f
C986 VDD2.n9 VSUBS 0.021678f
C987 VDD2.n10 VSUBS 0.011649f
C988 VDD2.n11 VSUBS 0.027534f
C989 VDD2.n12 VSUBS 0.012334f
C990 VDD2.n13 VSUBS 0.109167f
C991 VDD2.t5 VSUBS 0.058731f
C992 VDD2.n14 VSUBS 0.02065f
C993 VDD2.n15 VSUBS 0.017515f
C994 VDD2.n16 VSUBS 0.011649f
C995 VDD2.n17 VSUBS 0.709755f
C996 VDD2.n18 VSUBS 0.021678f
C997 VDD2.n19 VSUBS 0.011649f
C998 VDD2.n20 VSUBS 0.012334f
C999 VDD2.n21 VSUBS 0.027534f
C1000 VDD2.n22 VSUBS 0.027534f
C1001 VDD2.n23 VSUBS 0.012334f
C1002 VDD2.n24 VSUBS 0.011649f
C1003 VDD2.n25 VSUBS 0.021678f
C1004 VDD2.n26 VSUBS 0.021678f
C1005 VDD2.n27 VSUBS 0.011649f
C1006 VDD2.n28 VSUBS 0.012334f
C1007 VDD2.n29 VSUBS 0.027534f
C1008 VDD2.n30 VSUBS 0.027534f
C1009 VDD2.n31 VSUBS 0.012334f
C1010 VDD2.n32 VSUBS 0.011649f
C1011 VDD2.n33 VSUBS 0.021678f
C1012 VDD2.n34 VSUBS 0.021678f
C1013 VDD2.n35 VSUBS 0.011649f
C1014 VDD2.n36 VSUBS 0.012334f
C1015 VDD2.n37 VSUBS 0.027534f
C1016 VDD2.n38 VSUBS 0.06979f
C1017 VDD2.n39 VSUBS 0.012334f
C1018 VDD2.n40 VSUBS 0.011649f
C1019 VDD2.n41 VSUBS 0.049812f
C1020 VDD2.n42 VSUBS 0.054987f
C1021 VDD2.t3 VSUBS 0.139615f
C1022 VDD2.t0 VSUBS 0.139615f
C1023 VDD2.n43 VSUBS 1.00304f
C1024 VDD2.n44 VSUBS 2.17407f
C1025 VDD2.n45 VSUBS 0.02474f
C1026 VDD2.n46 VSUBS 0.021678f
C1027 VDD2.n47 VSUBS 0.011649f
C1028 VDD2.n48 VSUBS 0.027534f
C1029 VDD2.n49 VSUBS 0.012334f
C1030 VDD2.n50 VSUBS 0.021678f
C1031 VDD2.n51 VSUBS 0.011649f
C1032 VDD2.n52 VSUBS 0.027534f
C1033 VDD2.n53 VSUBS 0.012334f
C1034 VDD2.n54 VSUBS 0.021678f
C1035 VDD2.n55 VSUBS 0.011649f
C1036 VDD2.n56 VSUBS 0.027534f
C1037 VDD2.n57 VSUBS 0.012334f
C1038 VDD2.n58 VSUBS 0.109167f
C1039 VDD2.t4 VSUBS 0.058731f
C1040 VDD2.n59 VSUBS 0.02065f
C1041 VDD2.n60 VSUBS 0.017515f
C1042 VDD2.n61 VSUBS 0.011649f
C1043 VDD2.n62 VSUBS 0.709755f
C1044 VDD2.n63 VSUBS 0.021678f
C1045 VDD2.n64 VSUBS 0.011649f
C1046 VDD2.n65 VSUBS 0.012334f
C1047 VDD2.n66 VSUBS 0.027534f
C1048 VDD2.n67 VSUBS 0.027534f
C1049 VDD2.n68 VSUBS 0.012334f
C1050 VDD2.n69 VSUBS 0.011649f
C1051 VDD2.n70 VSUBS 0.021678f
C1052 VDD2.n71 VSUBS 0.021678f
C1053 VDD2.n72 VSUBS 0.011649f
C1054 VDD2.n73 VSUBS 0.012334f
C1055 VDD2.n74 VSUBS 0.027534f
C1056 VDD2.n75 VSUBS 0.027534f
C1057 VDD2.n76 VSUBS 0.012334f
C1058 VDD2.n77 VSUBS 0.011649f
C1059 VDD2.n78 VSUBS 0.021678f
C1060 VDD2.n79 VSUBS 0.021678f
C1061 VDD2.n80 VSUBS 0.011649f
C1062 VDD2.n81 VSUBS 0.012334f
C1063 VDD2.n82 VSUBS 0.027534f
C1064 VDD2.n83 VSUBS 0.06979f
C1065 VDD2.n84 VSUBS 0.012334f
C1066 VDD2.n85 VSUBS 0.011649f
C1067 VDD2.n86 VSUBS 0.049812f
C1068 VDD2.n87 VSUBS 0.050198f
C1069 VDD2.n88 VSUBS 1.86546f
C1070 VDD2.t2 VSUBS 0.139615f
C1071 VDD2.t1 VSUBS 0.139615f
C1072 VDD2.n89 VSUBS 1.00302f
C1073 VN.n0 VSUBS 0.048667f
C1074 VN.t1 VSUBS 1.77898f
C1075 VN.n1 VSUBS 0.029949f
C1076 VN.n2 VSUBS 0.314217f
C1077 VN.t4 VSUBS 1.77898f
C1078 VN.t5 VSUBS 2.00544f
C1079 VN.n3 VSUBS 0.736041f
C1080 VN.n4 VSUBS 0.747479f
C1081 VN.n5 VSUBS 0.051815f
C1082 VN.n6 VSUBS 0.073868f
C1083 VN.n7 VSUBS 0.036913f
C1084 VN.n8 VSUBS 0.036913f
C1085 VN.n9 VSUBS 0.036913f
C1086 VN.n10 VSUBS 0.072761f
C1087 VN.n11 VSUBS 0.053853f
C1088 VN.n12 VSUBS 0.763247f
C1089 VN.n13 VSUBS 0.05238f
C1090 VN.n14 VSUBS 0.048667f
C1091 VN.t3 VSUBS 1.77898f
C1092 VN.n15 VSUBS 0.029949f
C1093 VN.n16 VSUBS 0.314217f
C1094 VN.t0 VSUBS 1.77898f
C1095 VN.t2 VSUBS 2.00544f
C1096 VN.n17 VSUBS 0.736041f
C1097 VN.n18 VSUBS 0.747479f
C1098 VN.n19 VSUBS 0.051815f
C1099 VN.n20 VSUBS 0.073868f
C1100 VN.n21 VSUBS 0.036913f
C1101 VN.n22 VSUBS 0.036913f
C1102 VN.n23 VSUBS 0.036913f
C1103 VN.n24 VSUBS 0.072761f
C1104 VN.n25 VSUBS 0.053853f
C1105 VN.n26 VSUBS 0.763247f
C1106 VN.n27 VSUBS 1.71325f
.ends

