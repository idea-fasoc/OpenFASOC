* NGSPICE file created from diff_pair_sample_1775.ext - technology: sky130A

.subckt diff_pair_sample_1775 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=0 ps=0 w=3.74 l=0.59
X1 B.t8 B.t6 B.t7 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=0 ps=0 w=3.74 l=0.59
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=1.4586 ps=8.26 w=3.74 l=0.59
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=1.4586 ps=8.26 w=3.74 l=0.59
X4 B.t5 B.t3 B.t4 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=0 ps=0 w=3.74 l=0.59
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=1.4586 ps=8.26 w=3.74 l=0.59
X6 B.t2 B.t0 B.t1 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=0 ps=0 w=3.74 l=0.59
X7 VDD2.t0 VN.t1 VTAIL.t2 w_n1338_n1720# sky130_fd_pr__pfet_01v8 ad=1.4586 pd=8.26 as=1.4586 ps=8.26 w=3.74 l=0.59
R0 B.n166 B.n49 585
R1 B.n165 B.n164 585
R2 B.n163 B.n50 585
R3 B.n162 B.n161 585
R4 B.n160 B.n51 585
R5 B.n159 B.n158 585
R6 B.n157 B.n52 585
R7 B.n156 B.n155 585
R8 B.n154 B.n53 585
R9 B.n153 B.n152 585
R10 B.n151 B.n54 585
R11 B.n150 B.n149 585
R12 B.n148 B.n55 585
R13 B.n147 B.n146 585
R14 B.n145 B.n56 585
R15 B.n144 B.n143 585
R16 B.n142 B.n57 585
R17 B.n140 B.n139 585
R18 B.n138 B.n60 585
R19 B.n137 B.n136 585
R20 B.n135 B.n61 585
R21 B.n134 B.n133 585
R22 B.n132 B.n62 585
R23 B.n131 B.n130 585
R24 B.n129 B.n63 585
R25 B.n128 B.n127 585
R26 B.n126 B.n64 585
R27 B.n125 B.n124 585
R28 B.n120 B.n65 585
R29 B.n119 B.n118 585
R30 B.n117 B.n66 585
R31 B.n116 B.n115 585
R32 B.n114 B.n67 585
R33 B.n113 B.n112 585
R34 B.n111 B.n68 585
R35 B.n110 B.n109 585
R36 B.n108 B.n69 585
R37 B.n107 B.n106 585
R38 B.n105 B.n70 585
R39 B.n104 B.n103 585
R40 B.n102 B.n71 585
R41 B.n101 B.n100 585
R42 B.n99 B.n72 585
R43 B.n98 B.n97 585
R44 B.n168 B.n167 585
R45 B.n169 B.n48 585
R46 B.n171 B.n170 585
R47 B.n172 B.n47 585
R48 B.n174 B.n173 585
R49 B.n175 B.n46 585
R50 B.n177 B.n176 585
R51 B.n178 B.n45 585
R52 B.n180 B.n179 585
R53 B.n181 B.n44 585
R54 B.n183 B.n182 585
R55 B.n184 B.n43 585
R56 B.n186 B.n185 585
R57 B.n187 B.n42 585
R58 B.n189 B.n188 585
R59 B.n190 B.n41 585
R60 B.n192 B.n191 585
R61 B.n193 B.n40 585
R62 B.n195 B.n194 585
R63 B.n196 B.n39 585
R64 B.n198 B.n197 585
R65 B.n199 B.n38 585
R66 B.n201 B.n200 585
R67 B.n202 B.n37 585
R68 B.n204 B.n203 585
R69 B.n205 B.n36 585
R70 B.n207 B.n206 585
R71 B.n208 B.n35 585
R72 B.n276 B.n275 585
R73 B.n274 B.n9 585
R74 B.n273 B.n272 585
R75 B.n271 B.n10 585
R76 B.n270 B.n269 585
R77 B.n268 B.n11 585
R78 B.n267 B.n266 585
R79 B.n265 B.n12 585
R80 B.n264 B.n263 585
R81 B.n262 B.n13 585
R82 B.n261 B.n260 585
R83 B.n259 B.n14 585
R84 B.n258 B.n257 585
R85 B.n256 B.n15 585
R86 B.n255 B.n254 585
R87 B.n253 B.n16 585
R88 B.n252 B.n251 585
R89 B.n249 B.n17 585
R90 B.n248 B.n247 585
R91 B.n246 B.n20 585
R92 B.n245 B.n244 585
R93 B.n243 B.n21 585
R94 B.n242 B.n241 585
R95 B.n240 B.n22 585
R96 B.n239 B.n238 585
R97 B.n237 B.n23 585
R98 B.n236 B.n235 585
R99 B.n234 B.n233 585
R100 B.n232 B.n27 585
R101 B.n231 B.n230 585
R102 B.n229 B.n28 585
R103 B.n228 B.n227 585
R104 B.n226 B.n29 585
R105 B.n225 B.n224 585
R106 B.n223 B.n30 585
R107 B.n222 B.n221 585
R108 B.n220 B.n31 585
R109 B.n219 B.n218 585
R110 B.n217 B.n32 585
R111 B.n216 B.n215 585
R112 B.n214 B.n33 585
R113 B.n213 B.n212 585
R114 B.n211 B.n34 585
R115 B.n210 B.n209 585
R116 B.n277 B.n8 585
R117 B.n279 B.n278 585
R118 B.n280 B.n7 585
R119 B.n282 B.n281 585
R120 B.n283 B.n6 585
R121 B.n285 B.n284 585
R122 B.n286 B.n5 585
R123 B.n288 B.n287 585
R124 B.n289 B.n4 585
R125 B.n291 B.n290 585
R126 B.n292 B.n3 585
R127 B.n294 B.n293 585
R128 B.n295 B.n0 585
R129 B.n2 B.n1 585
R130 B.n80 B.n79 585
R131 B.n81 B.n78 585
R132 B.n83 B.n82 585
R133 B.n84 B.n77 585
R134 B.n86 B.n85 585
R135 B.n87 B.n76 585
R136 B.n89 B.n88 585
R137 B.n90 B.n75 585
R138 B.n92 B.n91 585
R139 B.n93 B.n74 585
R140 B.n95 B.n94 585
R141 B.n96 B.n73 585
R142 B.n98 B.n73 530.939
R143 B.n168 B.n49 530.939
R144 B.n210 B.n35 530.939
R145 B.n277 B.n276 530.939
R146 B.n121 B.t3 357.339
R147 B.n58 B.t6 357.339
R148 B.n24 B.t0 357.339
R149 B.n18 B.t9 357.339
R150 B.n297 B.n296 256.663
R151 B.n58 B.t7 248.429
R152 B.n24 B.t2 248.429
R153 B.n121 B.t4 248.429
R154 B.n18 B.t11 248.429
R155 B.n296 B.n295 235.042
R156 B.n296 B.n2 235.042
R157 B.n59 B.t8 230.588
R158 B.n25 B.t1 230.588
R159 B.n122 B.t5 230.588
R160 B.n19 B.t10 230.588
R161 B.n99 B.n98 163.367
R162 B.n100 B.n99 163.367
R163 B.n100 B.n71 163.367
R164 B.n104 B.n71 163.367
R165 B.n105 B.n104 163.367
R166 B.n106 B.n105 163.367
R167 B.n106 B.n69 163.367
R168 B.n110 B.n69 163.367
R169 B.n111 B.n110 163.367
R170 B.n112 B.n111 163.367
R171 B.n112 B.n67 163.367
R172 B.n116 B.n67 163.367
R173 B.n117 B.n116 163.367
R174 B.n118 B.n117 163.367
R175 B.n118 B.n65 163.367
R176 B.n125 B.n65 163.367
R177 B.n126 B.n125 163.367
R178 B.n127 B.n126 163.367
R179 B.n127 B.n63 163.367
R180 B.n131 B.n63 163.367
R181 B.n132 B.n131 163.367
R182 B.n133 B.n132 163.367
R183 B.n133 B.n61 163.367
R184 B.n137 B.n61 163.367
R185 B.n138 B.n137 163.367
R186 B.n139 B.n138 163.367
R187 B.n139 B.n57 163.367
R188 B.n144 B.n57 163.367
R189 B.n145 B.n144 163.367
R190 B.n146 B.n145 163.367
R191 B.n146 B.n55 163.367
R192 B.n150 B.n55 163.367
R193 B.n151 B.n150 163.367
R194 B.n152 B.n151 163.367
R195 B.n152 B.n53 163.367
R196 B.n156 B.n53 163.367
R197 B.n157 B.n156 163.367
R198 B.n158 B.n157 163.367
R199 B.n158 B.n51 163.367
R200 B.n162 B.n51 163.367
R201 B.n163 B.n162 163.367
R202 B.n164 B.n163 163.367
R203 B.n164 B.n49 163.367
R204 B.n206 B.n35 163.367
R205 B.n206 B.n205 163.367
R206 B.n205 B.n204 163.367
R207 B.n204 B.n37 163.367
R208 B.n200 B.n37 163.367
R209 B.n200 B.n199 163.367
R210 B.n199 B.n198 163.367
R211 B.n198 B.n39 163.367
R212 B.n194 B.n39 163.367
R213 B.n194 B.n193 163.367
R214 B.n193 B.n192 163.367
R215 B.n192 B.n41 163.367
R216 B.n188 B.n41 163.367
R217 B.n188 B.n187 163.367
R218 B.n187 B.n186 163.367
R219 B.n186 B.n43 163.367
R220 B.n182 B.n43 163.367
R221 B.n182 B.n181 163.367
R222 B.n181 B.n180 163.367
R223 B.n180 B.n45 163.367
R224 B.n176 B.n45 163.367
R225 B.n176 B.n175 163.367
R226 B.n175 B.n174 163.367
R227 B.n174 B.n47 163.367
R228 B.n170 B.n47 163.367
R229 B.n170 B.n169 163.367
R230 B.n169 B.n168 163.367
R231 B.n276 B.n9 163.367
R232 B.n272 B.n9 163.367
R233 B.n272 B.n271 163.367
R234 B.n271 B.n270 163.367
R235 B.n270 B.n11 163.367
R236 B.n266 B.n11 163.367
R237 B.n266 B.n265 163.367
R238 B.n265 B.n264 163.367
R239 B.n264 B.n13 163.367
R240 B.n260 B.n13 163.367
R241 B.n260 B.n259 163.367
R242 B.n259 B.n258 163.367
R243 B.n258 B.n15 163.367
R244 B.n254 B.n15 163.367
R245 B.n254 B.n253 163.367
R246 B.n253 B.n252 163.367
R247 B.n252 B.n17 163.367
R248 B.n247 B.n17 163.367
R249 B.n247 B.n246 163.367
R250 B.n246 B.n245 163.367
R251 B.n245 B.n21 163.367
R252 B.n241 B.n21 163.367
R253 B.n241 B.n240 163.367
R254 B.n240 B.n239 163.367
R255 B.n239 B.n23 163.367
R256 B.n235 B.n23 163.367
R257 B.n235 B.n234 163.367
R258 B.n234 B.n27 163.367
R259 B.n230 B.n27 163.367
R260 B.n230 B.n229 163.367
R261 B.n229 B.n228 163.367
R262 B.n228 B.n29 163.367
R263 B.n224 B.n29 163.367
R264 B.n224 B.n223 163.367
R265 B.n223 B.n222 163.367
R266 B.n222 B.n31 163.367
R267 B.n218 B.n31 163.367
R268 B.n218 B.n217 163.367
R269 B.n217 B.n216 163.367
R270 B.n216 B.n33 163.367
R271 B.n212 B.n33 163.367
R272 B.n212 B.n211 163.367
R273 B.n211 B.n210 163.367
R274 B.n278 B.n277 163.367
R275 B.n278 B.n7 163.367
R276 B.n282 B.n7 163.367
R277 B.n283 B.n282 163.367
R278 B.n284 B.n283 163.367
R279 B.n284 B.n5 163.367
R280 B.n288 B.n5 163.367
R281 B.n289 B.n288 163.367
R282 B.n290 B.n289 163.367
R283 B.n290 B.n3 163.367
R284 B.n294 B.n3 163.367
R285 B.n295 B.n294 163.367
R286 B.n80 B.n2 163.367
R287 B.n81 B.n80 163.367
R288 B.n82 B.n81 163.367
R289 B.n82 B.n77 163.367
R290 B.n86 B.n77 163.367
R291 B.n87 B.n86 163.367
R292 B.n88 B.n87 163.367
R293 B.n88 B.n75 163.367
R294 B.n92 B.n75 163.367
R295 B.n93 B.n92 163.367
R296 B.n94 B.n93 163.367
R297 B.n94 B.n73 163.367
R298 B.n123 B.n122 59.5399
R299 B.n141 B.n59 59.5399
R300 B.n26 B.n25 59.5399
R301 B.n250 B.n19 59.5399
R302 B.n275 B.n8 34.4981
R303 B.n209 B.n208 34.4981
R304 B.n167 B.n166 34.4981
R305 B.n97 B.n96 34.4981
R306 B B.n297 18.0485
R307 B.n122 B.n121 17.8429
R308 B.n59 B.n58 17.8429
R309 B.n25 B.n24 17.8429
R310 B.n19 B.n18 17.8429
R311 B.n279 B.n8 10.6151
R312 B.n280 B.n279 10.6151
R313 B.n281 B.n280 10.6151
R314 B.n281 B.n6 10.6151
R315 B.n285 B.n6 10.6151
R316 B.n286 B.n285 10.6151
R317 B.n287 B.n286 10.6151
R318 B.n287 B.n4 10.6151
R319 B.n291 B.n4 10.6151
R320 B.n292 B.n291 10.6151
R321 B.n293 B.n292 10.6151
R322 B.n293 B.n0 10.6151
R323 B.n275 B.n274 10.6151
R324 B.n274 B.n273 10.6151
R325 B.n273 B.n10 10.6151
R326 B.n269 B.n10 10.6151
R327 B.n269 B.n268 10.6151
R328 B.n268 B.n267 10.6151
R329 B.n267 B.n12 10.6151
R330 B.n263 B.n12 10.6151
R331 B.n263 B.n262 10.6151
R332 B.n262 B.n261 10.6151
R333 B.n261 B.n14 10.6151
R334 B.n257 B.n14 10.6151
R335 B.n257 B.n256 10.6151
R336 B.n256 B.n255 10.6151
R337 B.n255 B.n16 10.6151
R338 B.n251 B.n16 10.6151
R339 B.n249 B.n248 10.6151
R340 B.n248 B.n20 10.6151
R341 B.n244 B.n20 10.6151
R342 B.n244 B.n243 10.6151
R343 B.n243 B.n242 10.6151
R344 B.n242 B.n22 10.6151
R345 B.n238 B.n22 10.6151
R346 B.n238 B.n237 10.6151
R347 B.n237 B.n236 10.6151
R348 B.n233 B.n232 10.6151
R349 B.n232 B.n231 10.6151
R350 B.n231 B.n28 10.6151
R351 B.n227 B.n28 10.6151
R352 B.n227 B.n226 10.6151
R353 B.n226 B.n225 10.6151
R354 B.n225 B.n30 10.6151
R355 B.n221 B.n30 10.6151
R356 B.n221 B.n220 10.6151
R357 B.n220 B.n219 10.6151
R358 B.n219 B.n32 10.6151
R359 B.n215 B.n32 10.6151
R360 B.n215 B.n214 10.6151
R361 B.n214 B.n213 10.6151
R362 B.n213 B.n34 10.6151
R363 B.n209 B.n34 10.6151
R364 B.n208 B.n207 10.6151
R365 B.n207 B.n36 10.6151
R366 B.n203 B.n36 10.6151
R367 B.n203 B.n202 10.6151
R368 B.n202 B.n201 10.6151
R369 B.n201 B.n38 10.6151
R370 B.n197 B.n38 10.6151
R371 B.n197 B.n196 10.6151
R372 B.n196 B.n195 10.6151
R373 B.n195 B.n40 10.6151
R374 B.n191 B.n40 10.6151
R375 B.n191 B.n190 10.6151
R376 B.n190 B.n189 10.6151
R377 B.n189 B.n42 10.6151
R378 B.n185 B.n42 10.6151
R379 B.n185 B.n184 10.6151
R380 B.n184 B.n183 10.6151
R381 B.n183 B.n44 10.6151
R382 B.n179 B.n44 10.6151
R383 B.n179 B.n178 10.6151
R384 B.n178 B.n177 10.6151
R385 B.n177 B.n46 10.6151
R386 B.n173 B.n46 10.6151
R387 B.n173 B.n172 10.6151
R388 B.n172 B.n171 10.6151
R389 B.n171 B.n48 10.6151
R390 B.n167 B.n48 10.6151
R391 B.n79 B.n1 10.6151
R392 B.n79 B.n78 10.6151
R393 B.n83 B.n78 10.6151
R394 B.n84 B.n83 10.6151
R395 B.n85 B.n84 10.6151
R396 B.n85 B.n76 10.6151
R397 B.n89 B.n76 10.6151
R398 B.n90 B.n89 10.6151
R399 B.n91 B.n90 10.6151
R400 B.n91 B.n74 10.6151
R401 B.n95 B.n74 10.6151
R402 B.n96 B.n95 10.6151
R403 B.n97 B.n72 10.6151
R404 B.n101 B.n72 10.6151
R405 B.n102 B.n101 10.6151
R406 B.n103 B.n102 10.6151
R407 B.n103 B.n70 10.6151
R408 B.n107 B.n70 10.6151
R409 B.n108 B.n107 10.6151
R410 B.n109 B.n108 10.6151
R411 B.n109 B.n68 10.6151
R412 B.n113 B.n68 10.6151
R413 B.n114 B.n113 10.6151
R414 B.n115 B.n114 10.6151
R415 B.n115 B.n66 10.6151
R416 B.n119 B.n66 10.6151
R417 B.n120 B.n119 10.6151
R418 B.n124 B.n120 10.6151
R419 B.n128 B.n64 10.6151
R420 B.n129 B.n128 10.6151
R421 B.n130 B.n129 10.6151
R422 B.n130 B.n62 10.6151
R423 B.n134 B.n62 10.6151
R424 B.n135 B.n134 10.6151
R425 B.n136 B.n135 10.6151
R426 B.n136 B.n60 10.6151
R427 B.n140 B.n60 10.6151
R428 B.n143 B.n142 10.6151
R429 B.n143 B.n56 10.6151
R430 B.n147 B.n56 10.6151
R431 B.n148 B.n147 10.6151
R432 B.n149 B.n148 10.6151
R433 B.n149 B.n54 10.6151
R434 B.n153 B.n54 10.6151
R435 B.n154 B.n153 10.6151
R436 B.n155 B.n154 10.6151
R437 B.n155 B.n52 10.6151
R438 B.n159 B.n52 10.6151
R439 B.n160 B.n159 10.6151
R440 B.n161 B.n160 10.6151
R441 B.n161 B.n50 10.6151
R442 B.n165 B.n50 10.6151
R443 B.n166 B.n165 10.6151
R444 B.n251 B.n250 8.74196
R445 B.n233 B.n26 8.74196
R446 B.n124 B.n123 8.74196
R447 B.n142 B.n141 8.74196
R448 B.n297 B.n0 8.11757
R449 B.n297 B.n1 8.11757
R450 B.n250 B.n249 1.87367
R451 B.n236 B.n26 1.87367
R452 B.n123 B.n64 1.87367
R453 B.n141 B.n140 1.87367
R454 VN VN.t1 414.115
R455 VN VN.t0 380.702
R456 VTAIL.n74 VTAIL.n60 756.745
R457 VTAIL.n14 VTAIL.n0 756.745
R458 VTAIL.n54 VTAIL.n40 756.745
R459 VTAIL.n34 VTAIL.n20 756.745
R460 VTAIL.n67 VTAIL.n66 585
R461 VTAIL.n64 VTAIL.n63 585
R462 VTAIL.n73 VTAIL.n72 585
R463 VTAIL.n75 VTAIL.n74 585
R464 VTAIL.n7 VTAIL.n6 585
R465 VTAIL.n4 VTAIL.n3 585
R466 VTAIL.n13 VTAIL.n12 585
R467 VTAIL.n15 VTAIL.n14 585
R468 VTAIL.n55 VTAIL.n54 585
R469 VTAIL.n53 VTAIL.n52 585
R470 VTAIL.n44 VTAIL.n43 585
R471 VTAIL.n47 VTAIL.n46 585
R472 VTAIL.n35 VTAIL.n34 585
R473 VTAIL.n33 VTAIL.n32 585
R474 VTAIL.n24 VTAIL.n23 585
R475 VTAIL.n27 VTAIL.n26 585
R476 VTAIL.t3 VTAIL.n65 330.707
R477 VTAIL.t0 VTAIL.n5 330.707
R478 VTAIL.t1 VTAIL.n45 330.707
R479 VTAIL.t2 VTAIL.n25 330.707
R480 VTAIL.n66 VTAIL.n63 171.744
R481 VTAIL.n73 VTAIL.n63 171.744
R482 VTAIL.n74 VTAIL.n73 171.744
R483 VTAIL.n6 VTAIL.n3 171.744
R484 VTAIL.n13 VTAIL.n3 171.744
R485 VTAIL.n14 VTAIL.n13 171.744
R486 VTAIL.n54 VTAIL.n53 171.744
R487 VTAIL.n53 VTAIL.n43 171.744
R488 VTAIL.n46 VTAIL.n43 171.744
R489 VTAIL.n34 VTAIL.n33 171.744
R490 VTAIL.n33 VTAIL.n23 171.744
R491 VTAIL.n26 VTAIL.n23 171.744
R492 VTAIL.n66 VTAIL.t3 85.8723
R493 VTAIL.n6 VTAIL.t0 85.8723
R494 VTAIL.n46 VTAIL.t1 85.8723
R495 VTAIL.n26 VTAIL.t2 85.8723
R496 VTAIL.n79 VTAIL.n78 30.246
R497 VTAIL.n19 VTAIL.n18 30.246
R498 VTAIL.n59 VTAIL.n58 30.246
R499 VTAIL.n39 VTAIL.n38 30.246
R500 VTAIL.n39 VTAIL.n19 17.1945
R501 VTAIL.n79 VTAIL.n59 16.4014
R502 VTAIL.n67 VTAIL.n65 16.3201
R503 VTAIL.n7 VTAIL.n5 16.3201
R504 VTAIL.n47 VTAIL.n45 16.3201
R505 VTAIL.n27 VTAIL.n25 16.3201
R506 VTAIL.n68 VTAIL.n64 12.8005
R507 VTAIL.n8 VTAIL.n4 12.8005
R508 VTAIL.n48 VTAIL.n44 12.8005
R509 VTAIL.n28 VTAIL.n24 12.8005
R510 VTAIL.n72 VTAIL.n71 12.0247
R511 VTAIL.n12 VTAIL.n11 12.0247
R512 VTAIL.n52 VTAIL.n51 12.0247
R513 VTAIL.n32 VTAIL.n31 12.0247
R514 VTAIL.n75 VTAIL.n62 11.249
R515 VTAIL.n15 VTAIL.n2 11.249
R516 VTAIL.n55 VTAIL.n42 11.249
R517 VTAIL.n35 VTAIL.n22 11.249
R518 VTAIL.n76 VTAIL.n60 10.4732
R519 VTAIL.n16 VTAIL.n0 10.4732
R520 VTAIL.n56 VTAIL.n40 10.4732
R521 VTAIL.n36 VTAIL.n20 10.4732
R522 VTAIL.n78 VTAIL.n77 9.45567
R523 VTAIL.n18 VTAIL.n17 9.45567
R524 VTAIL.n58 VTAIL.n57 9.45567
R525 VTAIL.n38 VTAIL.n37 9.45567
R526 VTAIL.n77 VTAIL.n76 9.3005
R527 VTAIL.n62 VTAIL.n61 9.3005
R528 VTAIL.n71 VTAIL.n70 9.3005
R529 VTAIL.n69 VTAIL.n68 9.3005
R530 VTAIL.n17 VTAIL.n16 9.3005
R531 VTAIL.n2 VTAIL.n1 9.3005
R532 VTAIL.n11 VTAIL.n10 9.3005
R533 VTAIL.n9 VTAIL.n8 9.3005
R534 VTAIL.n57 VTAIL.n56 9.3005
R535 VTAIL.n42 VTAIL.n41 9.3005
R536 VTAIL.n51 VTAIL.n50 9.3005
R537 VTAIL.n49 VTAIL.n48 9.3005
R538 VTAIL.n37 VTAIL.n36 9.3005
R539 VTAIL.n22 VTAIL.n21 9.3005
R540 VTAIL.n31 VTAIL.n30 9.3005
R541 VTAIL.n29 VTAIL.n28 9.3005
R542 VTAIL.n69 VTAIL.n65 3.78097
R543 VTAIL.n9 VTAIL.n5 3.78097
R544 VTAIL.n49 VTAIL.n45 3.78097
R545 VTAIL.n29 VTAIL.n25 3.78097
R546 VTAIL.n78 VTAIL.n60 3.49141
R547 VTAIL.n18 VTAIL.n0 3.49141
R548 VTAIL.n58 VTAIL.n40 3.49141
R549 VTAIL.n38 VTAIL.n20 3.49141
R550 VTAIL.n76 VTAIL.n75 2.71565
R551 VTAIL.n16 VTAIL.n15 2.71565
R552 VTAIL.n56 VTAIL.n55 2.71565
R553 VTAIL.n36 VTAIL.n35 2.71565
R554 VTAIL.n72 VTAIL.n62 1.93989
R555 VTAIL.n12 VTAIL.n2 1.93989
R556 VTAIL.n52 VTAIL.n42 1.93989
R557 VTAIL.n32 VTAIL.n22 1.93989
R558 VTAIL.n71 VTAIL.n64 1.16414
R559 VTAIL.n11 VTAIL.n4 1.16414
R560 VTAIL.n51 VTAIL.n44 1.16414
R561 VTAIL.n31 VTAIL.n24 1.16414
R562 VTAIL.n59 VTAIL.n39 0.866879
R563 VTAIL VTAIL.n19 0.726793
R564 VTAIL.n68 VTAIL.n67 0.388379
R565 VTAIL.n8 VTAIL.n7 0.388379
R566 VTAIL.n48 VTAIL.n47 0.388379
R567 VTAIL.n28 VTAIL.n27 0.388379
R568 VTAIL.n70 VTAIL.n69 0.155672
R569 VTAIL.n70 VTAIL.n61 0.155672
R570 VTAIL.n77 VTAIL.n61 0.155672
R571 VTAIL.n10 VTAIL.n9 0.155672
R572 VTAIL.n10 VTAIL.n1 0.155672
R573 VTAIL.n17 VTAIL.n1 0.155672
R574 VTAIL.n57 VTAIL.n41 0.155672
R575 VTAIL.n50 VTAIL.n41 0.155672
R576 VTAIL.n50 VTAIL.n49 0.155672
R577 VTAIL.n37 VTAIL.n21 0.155672
R578 VTAIL.n30 VTAIL.n21 0.155672
R579 VTAIL.n30 VTAIL.n29 0.155672
R580 VTAIL VTAIL.n79 0.140586
R581 VDD2.n33 VDD2.n19 756.745
R582 VDD2.n14 VDD2.n0 756.745
R583 VDD2.n34 VDD2.n33 585
R584 VDD2.n32 VDD2.n31 585
R585 VDD2.n23 VDD2.n22 585
R586 VDD2.n26 VDD2.n25 585
R587 VDD2.n7 VDD2.n6 585
R588 VDD2.n4 VDD2.n3 585
R589 VDD2.n13 VDD2.n12 585
R590 VDD2.n15 VDD2.n14 585
R591 VDD2.t0 VDD2.n24 330.707
R592 VDD2.t1 VDD2.n5 330.707
R593 VDD2.n33 VDD2.n32 171.744
R594 VDD2.n32 VDD2.n22 171.744
R595 VDD2.n25 VDD2.n22 171.744
R596 VDD2.n6 VDD2.n3 171.744
R597 VDD2.n13 VDD2.n3 171.744
R598 VDD2.n14 VDD2.n13 171.744
R599 VDD2.n25 VDD2.t0 85.8723
R600 VDD2.n6 VDD2.t1 85.8723
R601 VDD2.n38 VDD2.n18 75.4118
R602 VDD2.n38 VDD2.n37 46.9247
R603 VDD2.n26 VDD2.n24 16.3201
R604 VDD2.n7 VDD2.n5 16.3201
R605 VDD2.n27 VDD2.n23 12.8005
R606 VDD2.n8 VDD2.n4 12.8005
R607 VDD2.n31 VDD2.n30 12.0247
R608 VDD2.n12 VDD2.n11 12.0247
R609 VDD2.n34 VDD2.n21 11.249
R610 VDD2.n15 VDD2.n2 11.249
R611 VDD2.n35 VDD2.n19 10.4732
R612 VDD2.n16 VDD2.n0 10.4732
R613 VDD2.n37 VDD2.n36 9.45567
R614 VDD2.n18 VDD2.n17 9.45567
R615 VDD2.n36 VDD2.n35 9.3005
R616 VDD2.n21 VDD2.n20 9.3005
R617 VDD2.n30 VDD2.n29 9.3005
R618 VDD2.n28 VDD2.n27 9.3005
R619 VDD2.n17 VDD2.n16 9.3005
R620 VDD2.n2 VDD2.n1 9.3005
R621 VDD2.n11 VDD2.n10 9.3005
R622 VDD2.n9 VDD2.n8 9.3005
R623 VDD2.n28 VDD2.n24 3.78097
R624 VDD2.n9 VDD2.n5 3.78097
R625 VDD2.n37 VDD2.n19 3.49141
R626 VDD2.n18 VDD2.n0 3.49141
R627 VDD2.n35 VDD2.n34 2.71565
R628 VDD2.n16 VDD2.n15 2.71565
R629 VDD2.n31 VDD2.n21 1.93989
R630 VDD2.n12 VDD2.n2 1.93989
R631 VDD2.n30 VDD2.n23 1.16414
R632 VDD2.n11 VDD2.n4 1.16414
R633 VDD2.n27 VDD2.n26 0.388379
R634 VDD2.n8 VDD2.n7 0.388379
R635 VDD2 VDD2.n38 0.256966
R636 VDD2.n36 VDD2.n20 0.155672
R637 VDD2.n29 VDD2.n20 0.155672
R638 VDD2.n29 VDD2.n28 0.155672
R639 VDD2.n10 VDD2.n9 0.155672
R640 VDD2.n10 VDD2.n1 0.155672
R641 VDD2.n17 VDD2.n1 0.155672
R642 VP.n0 VP.t0 413.735
R643 VP.n0 VP.t1 380.651
R644 VP VP.n0 0.0516364
R645 VDD1.n14 VDD1.n0 756.745
R646 VDD1.n33 VDD1.n19 756.745
R647 VDD1.n15 VDD1.n14 585
R648 VDD1.n13 VDD1.n12 585
R649 VDD1.n4 VDD1.n3 585
R650 VDD1.n7 VDD1.n6 585
R651 VDD1.n26 VDD1.n25 585
R652 VDD1.n23 VDD1.n22 585
R653 VDD1.n32 VDD1.n31 585
R654 VDD1.n34 VDD1.n33 585
R655 VDD1.t1 VDD1.n5 330.707
R656 VDD1.t0 VDD1.n24 330.707
R657 VDD1.n14 VDD1.n13 171.744
R658 VDD1.n13 VDD1.n3 171.744
R659 VDD1.n6 VDD1.n3 171.744
R660 VDD1.n25 VDD1.n22 171.744
R661 VDD1.n32 VDD1.n22 171.744
R662 VDD1.n33 VDD1.n32 171.744
R663 VDD1.n6 VDD1.t1 85.8723
R664 VDD1.n25 VDD1.t0 85.8723
R665 VDD1 VDD1.n37 76.1349
R666 VDD1 VDD1.n18 47.1812
R667 VDD1.n7 VDD1.n5 16.3201
R668 VDD1.n26 VDD1.n24 16.3201
R669 VDD1.n8 VDD1.n4 12.8005
R670 VDD1.n27 VDD1.n23 12.8005
R671 VDD1.n12 VDD1.n11 12.0247
R672 VDD1.n31 VDD1.n30 12.0247
R673 VDD1.n15 VDD1.n2 11.249
R674 VDD1.n34 VDD1.n21 11.249
R675 VDD1.n16 VDD1.n0 10.4732
R676 VDD1.n35 VDD1.n19 10.4732
R677 VDD1.n18 VDD1.n17 9.45567
R678 VDD1.n37 VDD1.n36 9.45567
R679 VDD1.n17 VDD1.n16 9.3005
R680 VDD1.n2 VDD1.n1 9.3005
R681 VDD1.n11 VDD1.n10 9.3005
R682 VDD1.n9 VDD1.n8 9.3005
R683 VDD1.n36 VDD1.n35 9.3005
R684 VDD1.n21 VDD1.n20 9.3005
R685 VDD1.n30 VDD1.n29 9.3005
R686 VDD1.n28 VDD1.n27 9.3005
R687 VDD1.n9 VDD1.n5 3.78097
R688 VDD1.n28 VDD1.n24 3.78097
R689 VDD1.n18 VDD1.n0 3.49141
R690 VDD1.n37 VDD1.n19 3.49141
R691 VDD1.n16 VDD1.n15 2.71565
R692 VDD1.n35 VDD1.n34 2.71565
R693 VDD1.n12 VDD1.n2 1.93989
R694 VDD1.n31 VDD1.n21 1.93989
R695 VDD1.n11 VDD1.n4 1.16414
R696 VDD1.n30 VDD1.n23 1.16414
R697 VDD1.n8 VDD1.n7 0.388379
R698 VDD1.n27 VDD1.n26 0.388379
R699 VDD1.n17 VDD1.n1 0.155672
R700 VDD1.n10 VDD1.n1 0.155672
R701 VDD1.n10 VDD1.n9 0.155672
R702 VDD1.n29 VDD1.n28 0.155672
R703 VDD1.n29 VDD1.n20 0.155672
R704 VDD1.n36 VDD1.n20 0.155672
C0 VDD1 w_n1338_n1720# 0.945259f
C1 B w_n1338_n1720# 4.31867f
C2 VDD1 VN 0.153277f
C3 VN B 0.608519f
C4 VDD2 VP 0.25422f
C5 VP VTAIL 0.661738f
C6 VDD2 VTAIL 2.68839f
C7 VDD1 B 0.798809f
C8 VP w_n1338_n1720# 1.6755f
C9 VDD2 w_n1338_n1720# 0.948404f
C10 w_n1338_n1720# VTAIL 1.53192f
C11 VN VP 2.9861f
C12 VDD2 VN 0.743579f
C13 VN VTAIL 0.647464f
C14 VDD1 VP 0.842627f
C15 VDD1 VDD2 0.449343f
C16 VDD1 VTAIL 2.65083f
C17 VN w_n1338_n1720# 1.51063f
C18 VP B 0.873283f
C19 VDD2 B 0.812632f
C20 B VTAIL 1.17712f
C21 VDD2 VSUBS 0.445339f
C22 VDD1 VSUBS 1.792004f
C23 VTAIL VSUBS 0.355274f
C24 VN VSUBS 3.49804f
C25 VP VSUBS 0.695098f
C26 B VSUBS 1.643694f
C27 w_n1338_n1720# VSUBS 29.013199f
C28 VDD1.n0 VSUBS 0.016607f
C29 VDD1.n1 VSUBS 0.016584f
C30 VDD1.n2 VSUBS 0.008912f
C31 VDD1.n3 VSUBS 0.021064f
C32 VDD1.n4 VSUBS 0.009436f
C33 VDD1.n5 VSUBS 0.062375f
C34 VDD1.t1 VSUBS 0.045686f
C35 VDD1.n6 VSUBS 0.015798f
C36 VDD1.n7 VSUBS 0.013249f
C37 VDD1.n8 VSUBS 0.008912f
C38 VDD1.n9 VSUBS 0.209742f
C39 VDD1.n10 VSUBS 0.016584f
C40 VDD1.n11 VSUBS 0.008912f
C41 VDD1.n12 VSUBS 0.009436f
C42 VDD1.n13 VSUBS 0.021064f
C43 VDD1.n14 VSUBS 0.045489f
C44 VDD1.n15 VSUBS 0.009436f
C45 VDD1.n16 VSUBS 0.008912f
C46 VDD1.n17 VSUBS 0.036068f
C47 VDD1.n18 VSUBS 0.034272f
C48 VDD1.n19 VSUBS 0.016607f
C49 VDD1.n20 VSUBS 0.016584f
C50 VDD1.n21 VSUBS 0.008912f
C51 VDD1.n22 VSUBS 0.021064f
C52 VDD1.n23 VSUBS 0.009436f
C53 VDD1.n24 VSUBS 0.062375f
C54 VDD1.t0 VSUBS 0.045686f
C55 VDD1.n25 VSUBS 0.015798f
C56 VDD1.n26 VSUBS 0.013249f
C57 VDD1.n27 VSUBS 0.008912f
C58 VDD1.n28 VSUBS 0.209742f
C59 VDD1.n29 VSUBS 0.016584f
C60 VDD1.n30 VSUBS 0.008912f
C61 VDD1.n31 VSUBS 0.009436f
C62 VDD1.n32 VSUBS 0.021064f
C63 VDD1.n33 VSUBS 0.045489f
C64 VDD1.n34 VSUBS 0.009436f
C65 VDD1.n35 VSUBS 0.008912f
C66 VDD1.n36 VSUBS 0.036068f
C67 VDD1.n37 VSUBS 0.259361f
C68 VP.t0 VSUBS 0.413662f
C69 VP.t1 VSUBS 0.321181f
C70 VP.n0 VSUBS 2.25382f
C71 VDD2.n0 VSUBS 0.016992f
C72 VDD2.n1 VSUBS 0.016969f
C73 VDD2.n2 VSUBS 0.009119f
C74 VDD2.n3 VSUBS 0.021553f
C75 VDD2.n4 VSUBS 0.009655f
C76 VDD2.n5 VSUBS 0.063823f
C77 VDD2.t1 VSUBS 0.046746f
C78 VDD2.n6 VSUBS 0.016165f
C79 VDD2.n7 VSUBS 0.013557f
C80 VDD2.n8 VSUBS 0.009119f
C81 VDD2.n9 VSUBS 0.214611f
C82 VDD2.n10 VSUBS 0.016969f
C83 VDD2.n11 VSUBS 0.009119f
C84 VDD2.n12 VSUBS 0.009655f
C85 VDD2.n13 VSUBS 0.021553f
C86 VDD2.n14 VSUBS 0.046545f
C87 VDD2.n15 VSUBS 0.009655f
C88 VDD2.n16 VSUBS 0.009119f
C89 VDD2.n17 VSUBS 0.036906f
C90 VDD2.n18 VSUBS 0.246455f
C91 VDD2.n19 VSUBS 0.016992f
C92 VDD2.n20 VSUBS 0.016969f
C93 VDD2.n21 VSUBS 0.009119f
C94 VDD2.n22 VSUBS 0.021553f
C95 VDD2.n23 VSUBS 0.009655f
C96 VDD2.n24 VSUBS 0.063823f
C97 VDD2.t0 VSUBS 0.046746f
C98 VDD2.n25 VSUBS 0.016165f
C99 VDD2.n26 VSUBS 0.013557f
C100 VDD2.n27 VSUBS 0.009119f
C101 VDD2.n28 VSUBS 0.214611f
C102 VDD2.n29 VSUBS 0.016969f
C103 VDD2.n30 VSUBS 0.009119f
C104 VDD2.n31 VSUBS 0.009655f
C105 VDD2.n32 VSUBS 0.021553f
C106 VDD2.n33 VSUBS 0.046545f
C107 VDD2.n34 VSUBS 0.009655f
C108 VDD2.n35 VSUBS 0.009119f
C109 VDD2.n36 VSUBS 0.036906f
C110 VDD2.n37 VSUBS 0.034821f
C111 VDD2.n38 VSUBS 1.18689f
C112 VTAIL.n0 VSUBS 0.019874f
C113 VTAIL.n1 VSUBS 0.019847f
C114 VTAIL.n2 VSUBS 0.010665f
C115 VTAIL.n3 VSUBS 0.025208f
C116 VTAIL.n4 VSUBS 0.011292f
C117 VTAIL.n5 VSUBS 0.074646f
C118 VTAIL.t0 VSUBS 0.054673f
C119 VTAIL.n6 VSUBS 0.018906f
C120 VTAIL.n7 VSUBS 0.015855f
C121 VTAIL.n8 VSUBS 0.010665f
C122 VTAIL.n9 VSUBS 0.251003f
C123 VTAIL.n10 VSUBS 0.019847f
C124 VTAIL.n11 VSUBS 0.010665f
C125 VTAIL.n12 VSUBS 0.011292f
C126 VTAIL.n13 VSUBS 0.025208f
C127 VTAIL.n14 VSUBS 0.054438f
C128 VTAIL.n15 VSUBS 0.011292f
C129 VTAIL.n16 VSUBS 0.010665f
C130 VTAIL.n17 VSUBS 0.043164f
C131 VTAIL.n18 VSUBS 0.026998f
C132 VTAIL.n19 VSUBS 0.640197f
C133 VTAIL.n20 VSUBS 0.019874f
C134 VTAIL.n21 VSUBS 0.019847f
C135 VTAIL.n22 VSUBS 0.010665f
C136 VTAIL.n23 VSUBS 0.025208f
C137 VTAIL.n24 VSUBS 0.011292f
C138 VTAIL.n25 VSUBS 0.074646f
C139 VTAIL.t2 VSUBS 0.054673f
C140 VTAIL.n26 VSUBS 0.018906f
C141 VTAIL.n27 VSUBS 0.015855f
C142 VTAIL.n28 VSUBS 0.010665f
C143 VTAIL.n29 VSUBS 0.251003f
C144 VTAIL.n30 VSUBS 0.019847f
C145 VTAIL.n31 VSUBS 0.010665f
C146 VTAIL.n32 VSUBS 0.011292f
C147 VTAIL.n33 VSUBS 0.025208f
C148 VTAIL.n34 VSUBS 0.054438f
C149 VTAIL.n35 VSUBS 0.011292f
C150 VTAIL.n36 VSUBS 0.010665f
C151 VTAIL.n37 VSUBS 0.043164f
C152 VTAIL.n38 VSUBS 0.026998f
C153 VTAIL.n39 VSUBS 0.649156f
C154 VTAIL.n40 VSUBS 0.019874f
C155 VTAIL.n41 VSUBS 0.019847f
C156 VTAIL.n42 VSUBS 0.010665f
C157 VTAIL.n43 VSUBS 0.025208f
C158 VTAIL.n44 VSUBS 0.011292f
C159 VTAIL.n45 VSUBS 0.074646f
C160 VTAIL.t1 VSUBS 0.054673f
C161 VTAIL.n46 VSUBS 0.018906f
C162 VTAIL.n47 VSUBS 0.015855f
C163 VTAIL.n48 VSUBS 0.010665f
C164 VTAIL.n49 VSUBS 0.251003f
C165 VTAIL.n50 VSUBS 0.019847f
C166 VTAIL.n51 VSUBS 0.010665f
C167 VTAIL.n52 VSUBS 0.011292f
C168 VTAIL.n53 VSUBS 0.025208f
C169 VTAIL.n54 VSUBS 0.054438f
C170 VTAIL.n55 VSUBS 0.011292f
C171 VTAIL.n56 VSUBS 0.010665f
C172 VTAIL.n57 VSUBS 0.043164f
C173 VTAIL.n58 VSUBS 0.026998f
C174 VTAIL.n59 VSUBS 0.598436f
C175 VTAIL.n60 VSUBS 0.019874f
C176 VTAIL.n61 VSUBS 0.019847f
C177 VTAIL.n62 VSUBS 0.010665f
C178 VTAIL.n63 VSUBS 0.025208f
C179 VTAIL.n64 VSUBS 0.011292f
C180 VTAIL.n65 VSUBS 0.074646f
C181 VTAIL.t3 VSUBS 0.054673f
C182 VTAIL.n66 VSUBS 0.018906f
C183 VTAIL.n67 VSUBS 0.015855f
C184 VTAIL.n68 VSUBS 0.010665f
C185 VTAIL.n69 VSUBS 0.251003f
C186 VTAIL.n70 VSUBS 0.019847f
C187 VTAIL.n71 VSUBS 0.010665f
C188 VTAIL.n72 VSUBS 0.011292f
C189 VTAIL.n73 VSUBS 0.025208f
C190 VTAIL.n74 VSUBS 0.054438f
C191 VTAIL.n75 VSUBS 0.011292f
C192 VTAIL.n76 VSUBS 0.010665f
C193 VTAIL.n77 VSUBS 0.043164f
C194 VTAIL.n78 VSUBS 0.026998f
C195 VTAIL.n79 VSUBS 0.551989f
C196 VN.t0 VSUBS 0.315228f
C197 VN.t1 VSUBS 0.409076f
C198 B.n0 VSUBS 0.006737f
C199 B.n1 VSUBS 0.006737f
C200 B.n2 VSUBS 0.009964f
C201 B.n3 VSUBS 0.007636f
C202 B.n4 VSUBS 0.007636f
C203 B.n5 VSUBS 0.007636f
C204 B.n6 VSUBS 0.007636f
C205 B.n7 VSUBS 0.007636f
C206 B.n8 VSUBS 0.018226f
C207 B.n9 VSUBS 0.007636f
C208 B.n10 VSUBS 0.007636f
C209 B.n11 VSUBS 0.007636f
C210 B.n12 VSUBS 0.007636f
C211 B.n13 VSUBS 0.007636f
C212 B.n14 VSUBS 0.007636f
C213 B.n15 VSUBS 0.007636f
C214 B.n16 VSUBS 0.007636f
C215 B.n17 VSUBS 0.007636f
C216 B.t10 VSUBS 0.058491f
C217 B.t11 VSUBS 0.065721f
C218 B.t9 VSUBS 0.106903f
C219 B.n18 VSUBS 0.121684f
C220 B.n19 VSUBS 0.11156f
C221 B.n20 VSUBS 0.007636f
C222 B.n21 VSUBS 0.007636f
C223 B.n22 VSUBS 0.007636f
C224 B.n23 VSUBS 0.007636f
C225 B.t1 VSUBS 0.058492f
C226 B.t2 VSUBS 0.065722f
C227 B.t0 VSUBS 0.106903f
C228 B.n24 VSUBS 0.121683f
C229 B.n25 VSUBS 0.111559f
C230 B.n26 VSUBS 0.017691f
C231 B.n27 VSUBS 0.007636f
C232 B.n28 VSUBS 0.007636f
C233 B.n29 VSUBS 0.007636f
C234 B.n30 VSUBS 0.007636f
C235 B.n31 VSUBS 0.007636f
C236 B.n32 VSUBS 0.007636f
C237 B.n33 VSUBS 0.007636f
C238 B.n34 VSUBS 0.007636f
C239 B.n35 VSUBS 0.018226f
C240 B.n36 VSUBS 0.007636f
C241 B.n37 VSUBS 0.007636f
C242 B.n38 VSUBS 0.007636f
C243 B.n39 VSUBS 0.007636f
C244 B.n40 VSUBS 0.007636f
C245 B.n41 VSUBS 0.007636f
C246 B.n42 VSUBS 0.007636f
C247 B.n43 VSUBS 0.007636f
C248 B.n44 VSUBS 0.007636f
C249 B.n45 VSUBS 0.007636f
C250 B.n46 VSUBS 0.007636f
C251 B.n47 VSUBS 0.007636f
C252 B.n48 VSUBS 0.007636f
C253 B.n49 VSUBS 0.01883f
C254 B.n50 VSUBS 0.007636f
C255 B.n51 VSUBS 0.007636f
C256 B.n52 VSUBS 0.007636f
C257 B.n53 VSUBS 0.007636f
C258 B.n54 VSUBS 0.007636f
C259 B.n55 VSUBS 0.007636f
C260 B.n56 VSUBS 0.007636f
C261 B.n57 VSUBS 0.007636f
C262 B.t8 VSUBS 0.058492f
C263 B.t7 VSUBS 0.065722f
C264 B.t6 VSUBS 0.106903f
C265 B.n58 VSUBS 0.121683f
C266 B.n59 VSUBS 0.111559f
C267 B.n60 VSUBS 0.007636f
C268 B.n61 VSUBS 0.007636f
C269 B.n62 VSUBS 0.007636f
C270 B.n63 VSUBS 0.007636f
C271 B.n64 VSUBS 0.004492f
C272 B.n65 VSUBS 0.007636f
C273 B.n66 VSUBS 0.007636f
C274 B.n67 VSUBS 0.007636f
C275 B.n68 VSUBS 0.007636f
C276 B.n69 VSUBS 0.007636f
C277 B.n70 VSUBS 0.007636f
C278 B.n71 VSUBS 0.007636f
C279 B.n72 VSUBS 0.007636f
C280 B.n73 VSUBS 0.018226f
C281 B.n74 VSUBS 0.007636f
C282 B.n75 VSUBS 0.007636f
C283 B.n76 VSUBS 0.007636f
C284 B.n77 VSUBS 0.007636f
C285 B.n78 VSUBS 0.007636f
C286 B.n79 VSUBS 0.007636f
C287 B.n80 VSUBS 0.007636f
C288 B.n81 VSUBS 0.007636f
C289 B.n82 VSUBS 0.007636f
C290 B.n83 VSUBS 0.007636f
C291 B.n84 VSUBS 0.007636f
C292 B.n85 VSUBS 0.007636f
C293 B.n86 VSUBS 0.007636f
C294 B.n87 VSUBS 0.007636f
C295 B.n88 VSUBS 0.007636f
C296 B.n89 VSUBS 0.007636f
C297 B.n90 VSUBS 0.007636f
C298 B.n91 VSUBS 0.007636f
C299 B.n92 VSUBS 0.007636f
C300 B.n93 VSUBS 0.007636f
C301 B.n94 VSUBS 0.007636f
C302 B.n95 VSUBS 0.007636f
C303 B.n96 VSUBS 0.018226f
C304 B.n97 VSUBS 0.01883f
C305 B.n98 VSUBS 0.01883f
C306 B.n99 VSUBS 0.007636f
C307 B.n100 VSUBS 0.007636f
C308 B.n101 VSUBS 0.007636f
C309 B.n102 VSUBS 0.007636f
C310 B.n103 VSUBS 0.007636f
C311 B.n104 VSUBS 0.007636f
C312 B.n105 VSUBS 0.007636f
C313 B.n106 VSUBS 0.007636f
C314 B.n107 VSUBS 0.007636f
C315 B.n108 VSUBS 0.007636f
C316 B.n109 VSUBS 0.007636f
C317 B.n110 VSUBS 0.007636f
C318 B.n111 VSUBS 0.007636f
C319 B.n112 VSUBS 0.007636f
C320 B.n113 VSUBS 0.007636f
C321 B.n114 VSUBS 0.007636f
C322 B.n115 VSUBS 0.007636f
C323 B.n116 VSUBS 0.007636f
C324 B.n117 VSUBS 0.007636f
C325 B.n118 VSUBS 0.007636f
C326 B.n119 VSUBS 0.007636f
C327 B.n120 VSUBS 0.007636f
C328 B.t5 VSUBS 0.058491f
C329 B.t4 VSUBS 0.065721f
C330 B.t3 VSUBS 0.106903f
C331 B.n121 VSUBS 0.121684f
C332 B.n122 VSUBS 0.11156f
C333 B.n123 VSUBS 0.017691f
C334 B.n124 VSUBS 0.006962f
C335 B.n125 VSUBS 0.007636f
C336 B.n126 VSUBS 0.007636f
C337 B.n127 VSUBS 0.007636f
C338 B.n128 VSUBS 0.007636f
C339 B.n129 VSUBS 0.007636f
C340 B.n130 VSUBS 0.007636f
C341 B.n131 VSUBS 0.007636f
C342 B.n132 VSUBS 0.007636f
C343 B.n133 VSUBS 0.007636f
C344 B.n134 VSUBS 0.007636f
C345 B.n135 VSUBS 0.007636f
C346 B.n136 VSUBS 0.007636f
C347 B.n137 VSUBS 0.007636f
C348 B.n138 VSUBS 0.007636f
C349 B.n139 VSUBS 0.007636f
C350 B.n140 VSUBS 0.004492f
C351 B.n141 VSUBS 0.017691f
C352 B.n142 VSUBS 0.006962f
C353 B.n143 VSUBS 0.007636f
C354 B.n144 VSUBS 0.007636f
C355 B.n145 VSUBS 0.007636f
C356 B.n146 VSUBS 0.007636f
C357 B.n147 VSUBS 0.007636f
C358 B.n148 VSUBS 0.007636f
C359 B.n149 VSUBS 0.007636f
C360 B.n150 VSUBS 0.007636f
C361 B.n151 VSUBS 0.007636f
C362 B.n152 VSUBS 0.007636f
C363 B.n153 VSUBS 0.007636f
C364 B.n154 VSUBS 0.007636f
C365 B.n155 VSUBS 0.007636f
C366 B.n156 VSUBS 0.007636f
C367 B.n157 VSUBS 0.007636f
C368 B.n158 VSUBS 0.007636f
C369 B.n159 VSUBS 0.007636f
C370 B.n160 VSUBS 0.007636f
C371 B.n161 VSUBS 0.007636f
C372 B.n162 VSUBS 0.007636f
C373 B.n163 VSUBS 0.007636f
C374 B.n164 VSUBS 0.007636f
C375 B.n165 VSUBS 0.007636f
C376 B.n166 VSUBS 0.017976f
C377 B.n167 VSUBS 0.01908f
C378 B.n168 VSUBS 0.018226f
C379 B.n169 VSUBS 0.007636f
C380 B.n170 VSUBS 0.007636f
C381 B.n171 VSUBS 0.007636f
C382 B.n172 VSUBS 0.007636f
C383 B.n173 VSUBS 0.007636f
C384 B.n174 VSUBS 0.007636f
C385 B.n175 VSUBS 0.007636f
C386 B.n176 VSUBS 0.007636f
C387 B.n177 VSUBS 0.007636f
C388 B.n178 VSUBS 0.007636f
C389 B.n179 VSUBS 0.007636f
C390 B.n180 VSUBS 0.007636f
C391 B.n181 VSUBS 0.007636f
C392 B.n182 VSUBS 0.007636f
C393 B.n183 VSUBS 0.007636f
C394 B.n184 VSUBS 0.007636f
C395 B.n185 VSUBS 0.007636f
C396 B.n186 VSUBS 0.007636f
C397 B.n187 VSUBS 0.007636f
C398 B.n188 VSUBS 0.007636f
C399 B.n189 VSUBS 0.007636f
C400 B.n190 VSUBS 0.007636f
C401 B.n191 VSUBS 0.007636f
C402 B.n192 VSUBS 0.007636f
C403 B.n193 VSUBS 0.007636f
C404 B.n194 VSUBS 0.007636f
C405 B.n195 VSUBS 0.007636f
C406 B.n196 VSUBS 0.007636f
C407 B.n197 VSUBS 0.007636f
C408 B.n198 VSUBS 0.007636f
C409 B.n199 VSUBS 0.007636f
C410 B.n200 VSUBS 0.007636f
C411 B.n201 VSUBS 0.007636f
C412 B.n202 VSUBS 0.007636f
C413 B.n203 VSUBS 0.007636f
C414 B.n204 VSUBS 0.007636f
C415 B.n205 VSUBS 0.007636f
C416 B.n206 VSUBS 0.007636f
C417 B.n207 VSUBS 0.007636f
C418 B.n208 VSUBS 0.018226f
C419 B.n209 VSUBS 0.01883f
C420 B.n210 VSUBS 0.01883f
C421 B.n211 VSUBS 0.007636f
C422 B.n212 VSUBS 0.007636f
C423 B.n213 VSUBS 0.007636f
C424 B.n214 VSUBS 0.007636f
C425 B.n215 VSUBS 0.007636f
C426 B.n216 VSUBS 0.007636f
C427 B.n217 VSUBS 0.007636f
C428 B.n218 VSUBS 0.007636f
C429 B.n219 VSUBS 0.007636f
C430 B.n220 VSUBS 0.007636f
C431 B.n221 VSUBS 0.007636f
C432 B.n222 VSUBS 0.007636f
C433 B.n223 VSUBS 0.007636f
C434 B.n224 VSUBS 0.007636f
C435 B.n225 VSUBS 0.007636f
C436 B.n226 VSUBS 0.007636f
C437 B.n227 VSUBS 0.007636f
C438 B.n228 VSUBS 0.007636f
C439 B.n229 VSUBS 0.007636f
C440 B.n230 VSUBS 0.007636f
C441 B.n231 VSUBS 0.007636f
C442 B.n232 VSUBS 0.007636f
C443 B.n233 VSUBS 0.006962f
C444 B.n234 VSUBS 0.007636f
C445 B.n235 VSUBS 0.007636f
C446 B.n236 VSUBS 0.004492f
C447 B.n237 VSUBS 0.007636f
C448 B.n238 VSUBS 0.007636f
C449 B.n239 VSUBS 0.007636f
C450 B.n240 VSUBS 0.007636f
C451 B.n241 VSUBS 0.007636f
C452 B.n242 VSUBS 0.007636f
C453 B.n243 VSUBS 0.007636f
C454 B.n244 VSUBS 0.007636f
C455 B.n245 VSUBS 0.007636f
C456 B.n246 VSUBS 0.007636f
C457 B.n247 VSUBS 0.007636f
C458 B.n248 VSUBS 0.007636f
C459 B.n249 VSUBS 0.004492f
C460 B.n250 VSUBS 0.017691f
C461 B.n251 VSUBS 0.006962f
C462 B.n252 VSUBS 0.007636f
C463 B.n253 VSUBS 0.007636f
C464 B.n254 VSUBS 0.007636f
C465 B.n255 VSUBS 0.007636f
C466 B.n256 VSUBS 0.007636f
C467 B.n257 VSUBS 0.007636f
C468 B.n258 VSUBS 0.007636f
C469 B.n259 VSUBS 0.007636f
C470 B.n260 VSUBS 0.007636f
C471 B.n261 VSUBS 0.007636f
C472 B.n262 VSUBS 0.007636f
C473 B.n263 VSUBS 0.007636f
C474 B.n264 VSUBS 0.007636f
C475 B.n265 VSUBS 0.007636f
C476 B.n266 VSUBS 0.007636f
C477 B.n267 VSUBS 0.007636f
C478 B.n268 VSUBS 0.007636f
C479 B.n269 VSUBS 0.007636f
C480 B.n270 VSUBS 0.007636f
C481 B.n271 VSUBS 0.007636f
C482 B.n272 VSUBS 0.007636f
C483 B.n273 VSUBS 0.007636f
C484 B.n274 VSUBS 0.007636f
C485 B.n275 VSUBS 0.01883f
C486 B.n276 VSUBS 0.01883f
C487 B.n277 VSUBS 0.018226f
C488 B.n278 VSUBS 0.007636f
C489 B.n279 VSUBS 0.007636f
C490 B.n280 VSUBS 0.007636f
C491 B.n281 VSUBS 0.007636f
C492 B.n282 VSUBS 0.007636f
C493 B.n283 VSUBS 0.007636f
C494 B.n284 VSUBS 0.007636f
C495 B.n285 VSUBS 0.007636f
C496 B.n286 VSUBS 0.007636f
C497 B.n287 VSUBS 0.007636f
C498 B.n288 VSUBS 0.007636f
C499 B.n289 VSUBS 0.007636f
C500 B.n290 VSUBS 0.007636f
C501 B.n291 VSUBS 0.007636f
C502 B.n292 VSUBS 0.007636f
C503 B.n293 VSUBS 0.007636f
C504 B.n294 VSUBS 0.007636f
C505 B.n295 VSUBS 0.009964f
C506 B.n296 VSUBS 0.010614f
C507 B.n297 VSUBS 0.021108f
.ends

