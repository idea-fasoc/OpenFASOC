* NGSPICE file created from diff_pair_sample_0074.ext - technology: sky130A

.subckt diff_pair_sample_0074 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=0.83655 pd=5.4 as=1.9773 ps=10.92 w=5.07 l=1.48
X1 VTAIL.t5 VP.t1 VDD1.t2 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0.83655 ps=5.4 w=5.07 l=1.48
X2 B.t11 B.t9 B.t10 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0 ps=0 w=5.07 l=1.48
X3 B.t8 B.t6 B.t7 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0 ps=0 w=5.07 l=1.48
X4 VDD2.t3 VN.t0 VTAIL.t3 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=0.83655 pd=5.4 as=1.9773 ps=10.92 w=5.07 l=1.48
X5 B.t5 B.t3 B.t4 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0 ps=0 w=5.07 l=1.48
X6 VDD2.t2 VN.t1 VTAIL.t0 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=0.83655 pd=5.4 as=1.9773 ps=10.92 w=5.07 l=1.48
X7 B.t2 B.t0 B.t1 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0 ps=0 w=5.07 l=1.48
X8 VTAIL.t1 VN.t2 VDD2.t1 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0.83655 ps=5.4 w=5.07 l=1.48
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0.83655 ps=5.4 w=5.07 l=1.48
X10 VDD1.t1 VP.t2 VTAIL.t4 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=0.83655 pd=5.4 as=1.9773 ps=10.92 w=5.07 l=1.48
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n2056_n1982# sky130_fd_pr__pfet_01v8 ad=1.9773 pd=10.92 as=0.83655 ps=5.4 w=5.07 l=1.48
R0 VP.n4 VP.n3 178.183
R1 VP.n12 VP.n11 178.183
R2 VP.n10 VP.n0 161.3
R3 VP.n9 VP.n8 161.3
R4 VP.n7 VP.n1 161.3
R5 VP.n6 VP.n5 161.3
R6 VP.n2 VP.t3 118.626
R7 VP.n2 VP.t2 118.312
R8 VP.n4 VP.t1 82.5593
R9 VP.n11 VP.t0 82.5593
R10 VP.n9 VP.n1 56.5193
R11 VP.n3 VP.n2 50.6296
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 7.58527
R15 VP.n11 VP.n10 7.58527
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VTAIL.n5 VTAIL.t6 93.0823
R23 VTAIL.n4 VTAIL.t0 93.0823
R24 VTAIL.n3 VTAIL.t2 93.0823
R25 VTAIL.n6 VTAIL.t4 93.0822
R26 VTAIL.n7 VTAIL.t3 93.0822
R27 VTAIL.n0 VTAIL.t1 93.0822
R28 VTAIL.n1 VTAIL.t7 93.0822
R29 VTAIL.n2 VTAIL.t5 93.0822
R30 VTAIL.n7 VTAIL.n6 18.2979
R31 VTAIL.n3 VTAIL.n2 18.2979
R32 VTAIL.n4 VTAIL.n3 1.56084
R33 VTAIL.n6 VTAIL.n5 1.56084
R34 VTAIL.n2 VTAIL.n1 1.56084
R35 VTAIL VTAIL.n0 0.838862
R36 VTAIL VTAIL.n7 0.722483
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 136.641
R40 VDD1 VDD1.n0 103.407
R41 VDD1.n0 VDD1.t0 6.41174
R42 VDD1.n0 VDD1.t1 6.41174
R43 VDD1.n1 VDD1.t2 6.41174
R44 VDD1.n1 VDD1.t3 6.41174
R45 B.n300 B.n299 585
R46 B.n301 B.n44 585
R47 B.n303 B.n302 585
R48 B.n304 B.n43 585
R49 B.n306 B.n305 585
R50 B.n307 B.n42 585
R51 B.n309 B.n308 585
R52 B.n310 B.n41 585
R53 B.n312 B.n311 585
R54 B.n313 B.n40 585
R55 B.n315 B.n314 585
R56 B.n316 B.n39 585
R57 B.n318 B.n317 585
R58 B.n319 B.n38 585
R59 B.n321 B.n320 585
R60 B.n322 B.n37 585
R61 B.n324 B.n323 585
R62 B.n325 B.n36 585
R63 B.n327 B.n326 585
R64 B.n328 B.n35 585
R65 B.n330 B.n329 585
R66 B.n332 B.n32 585
R67 B.n334 B.n333 585
R68 B.n335 B.n31 585
R69 B.n337 B.n336 585
R70 B.n338 B.n30 585
R71 B.n340 B.n339 585
R72 B.n341 B.n29 585
R73 B.n343 B.n342 585
R74 B.n344 B.n25 585
R75 B.n346 B.n345 585
R76 B.n347 B.n24 585
R77 B.n349 B.n348 585
R78 B.n350 B.n23 585
R79 B.n352 B.n351 585
R80 B.n353 B.n22 585
R81 B.n355 B.n354 585
R82 B.n356 B.n21 585
R83 B.n358 B.n357 585
R84 B.n359 B.n20 585
R85 B.n361 B.n360 585
R86 B.n362 B.n19 585
R87 B.n364 B.n363 585
R88 B.n365 B.n18 585
R89 B.n367 B.n366 585
R90 B.n368 B.n17 585
R91 B.n370 B.n369 585
R92 B.n371 B.n16 585
R93 B.n373 B.n372 585
R94 B.n374 B.n15 585
R95 B.n376 B.n375 585
R96 B.n377 B.n14 585
R97 B.n298 B.n45 585
R98 B.n297 B.n296 585
R99 B.n295 B.n46 585
R100 B.n294 B.n293 585
R101 B.n292 B.n47 585
R102 B.n291 B.n290 585
R103 B.n289 B.n48 585
R104 B.n288 B.n287 585
R105 B.n286 B.n49 585
R106 B.n285 B.n284 585
R107 B.n283 B.n50 585
R108 B.n282 B.n281 585
R109 B.n280 B.n51 585
R110 B.n279 B.n278 585
R111 B.n277 B.n52 585
R112 B.n276 B.n275 585
R113 B.n274 B.n53 585
R114 B.n273 B.n272 585
R115 B.n271 B.n54 585
R116 B.n270 B.n269 585
R117 B.n268 B.n55 585
R118 B.n267 B.n266 585
R119 B.n265 B.n56 585
R120 B.n264 B.n263 585
R121 B.n262 B.n57 585
R122 B.n261 B.n260 585
R123 B.n259 B.n58 585
R124 B.n258 B.n257 585
R125 B.n256 B.n59 585
R126 B.n255 B.n254 585
R127 B.n253 B.n60 585
R128 B.n252 B.n251 585
R129 B.n250 B.n61 585
R130 B.n249 B.n248 585
R131 B.n247 B.n62 585
R132 B.n246 B.n245 585
R133 B.n244 B.n63 585
R134 B.n243 B.n242 585
R135 B.n241 B.n64 585
R136 B.n240 B.n239 585
R137 B.n238 B.n65 585
R138 B.n237 B.n236 585
R139 B.n235 B.n66 585
R140 B.n234 B.n233 585
R141 B.n232 B.n67 585
R142 B.n231 B.n230 585
R143 B.n229 B.n68 585
R144 B.n228 B.n227 585
R145 B.n226 B.n69 585
R146 B.n147 B.n146 585
R147 B.n148 B.n99 585
R148 B.n150 B.n149 585
R149 B.n151 B.n98 585
R150 B.n153 B.n152 585
R151 B.n154 B.n97 585
R152 B.n156 B.n155 585
R153 B.n157 B.n96 585
R154 B.n159 B.n158 585
R155 B.n160 B.n95 585
R156 B.n162 B.n161 585
R157 B.n163 B.n94 585
R158 B.n165 B.n164 585
R159 B.n166 B.n93 585
R160 B.n168 B.n167 585
R161 B.n169 B.n92 585
R162 B.n171 B.n170 585
R163 B.n172 B.n91 585
R164 B.n174 B.n173 585
R165 B.n175 B.n90 585
R166 B.n177 B.n176 585
R167 B.n179 B.n178 585
R168 B.n180 B.n86 585
R169 B.n182 B.n181 585
R170 B.n183 B.n85 585
R171 B.n185 B.n184 585
R172 B.n186 B.n84 585
R173 B.n188 B.n187 585
R174 B.n189 B.n83 585
R175 B.n191 B.n190 585
R176 B.n192 B.n80 585
R177 B.n195 B.n194 585
R178 B.n196 B.n79 585
R179 B.n198 B.n197 585
R180 B.n199 B.n78 585
R181 B.n201 B.n200 585
R182 B.n202 B.n77 585
R183 B.n204 B.n203 585
R184 B.n205 B.n76 585
R185 B.n207 B.n206 585
R186 B.n208 B.n75 585
R187 B.n210 B.n209 585
R188 B.n211 B.n74 585
R189 B.n213 B.n212 585
R190 B.n214 B.n73 585
R191 B.n216 B.n215 585
R192 B.n217 B.n72 585
R193 B.n219 B.n218 585
R194 B.n220 B.n71 585
R195 B.n222 B.n221 585
R196 B.n223 B.n70 585
R197 B.n225 B.n224 585
R198 B.n145 B.n100 585
R199 B.n144 B.n143 585
R200 B.n142 B.n101 585
R201 B.n141 B.n140 585
R202 B.n139 B.n102 585
R203 B.n138 B.n137 585
R204 B.n136 B.n103 585
R205 B.n135 B.n134 585
R206 B.n133 B.n104 585
R207 B.n132 B.n131 585
R208 B.n130 B.n105 585
R209 B.n129 B.n128 585
R210 B.n127 B.n106 585
R211 B.n126 B.n125 585
R212 B.n124 B.n107 585
R213 B.n123 B.n122 585
R214 B.n121 B.n108 585
R215 B.n120 B.n119 585
R216 B.n118 B.n109 585
R217 B.n117 B.n116 585
R218 B.n115 B.n110 585
R219 B.n114 B.n113 585
R220 B.n112 B.n111 585
R221 B.n2 B.n0 585
R222 B.n413 B.n1 585
R223 B.n412 B.n411 585
R224 B.n410 B.n3 585
R225 B.n409 B.n408 585
R226 B.n407 B.n4 585
R227 B.n406 B.n405 585
R228 B.n404 B.n5 585
R229 B.n403 B.n402 585
R230 B.n401 B.n6 585
R231 B.n400 B.n399 585
R232 B.n398 B.n7 585
R233 B.n397 B.n396 585
R234 B.n395 B.n8 585
R235 B.n394 B.n393 585
R236 B.n392 B.n9 585
R237 B.n391 B.n390 585
R238 B.n389 B.n10 585
R239 B.n388 B.n387 585
R240 B.n386 B.n11 585
R241 B.n385 B.n384 585
R242 B.n383 B.n12 585
R243 B.n382 B.n381 585
R244 B.n380 B.n13 585
R245 B.n379 B.n378 585
R246 B.n415 B.n414 585
R247 B.n147 B.n100 516.524
R248 B.n378 B.n377 516.524
R249 B.n226 B.n225 516.524
R250 B.n299 B.n298 516.524
R251 B.n81 B.t0 287.923
R252 B.n87 B.t6 287.923
R253 B.n26 B.t3 287.923
R254 B.n33 B.t9 287.923
R255 B.n143 B.n100 163.367
R256 B.n143 B.n142 163.367
R257 B.n142 B.n141 163.367
R258 B.n141 B.n102 163.367
R259 B.n137 B.n102 163.367
R260 B.n137 B.n136 163.367
R261 B.n136 B.n135 163.367
R262 B.n135 B.n104 163.367
R263 B.n131 B.n104 163.367
R264 B.n131 B.n130 163.367
R265 B.n130 B.n129 163.367
R266 B.n129 B.n106 163.367
R267 B.n125 B.n106 163.367
R268 B.n125 B.n124 163.367
R269 B.n124 B.n123 163.367
R270 B.n123 B.n108 163.367
R271 B.n119 B.n108 163.367
R272 B.n119 B.n118 163.367
R273 B.n118 B.n117 163.367
R274 B.n117 B.n110 163.367
R275 B.n113 B.n110 163.367
R276 B.n113 B.n112 163.367
R277 B.n112 B.n2 163.367
R278 B.n414 B.n2 163.367
R279 B.n414 B.n413 163.367
R280 B.n413 B.n412 163.367
R281 B.n412 B.n3 163.367
R282 B.n408 B.n3 163.367
R283 B.n408 B.n407 163.367
R284 B.n407 B.n406 163.367
R285 B.n406 B.n5 163.367
R286 B.n402 B.n5 163.367
R287 B.n402 B.n401 163.367
R288 B.n401 B.n400 163.367
R289 B.n400 B.n7 163.367
R290 B.n396 B.n7 163.367
R291 B.n396 B.n395 163.367
R292 B.n395 B.n394 163.367
R293 B.n394 B.n9 163.367
R294 B.n390 B.n9 163.367
R295 B.n390 B.n389 163.367
R296 B.n389 B.n388 163.367
R297 B.n388 B.n11 163.367
R298 B.n384 B.n11 163.367
R299 B.n384 B.n383 163.367
R300 B.n383 B.n382 163.367
R301 B.n382 B.n13 163.367
R302 B.n378 B.n13 163.367
R303 B.n148 B.n147 163.367
R304 B.n149 B.n148 163.367
R305 B.n149 B.n98 163.367
R306 B.n153 B.n98 163.367
R307 B.n154 B.n153 163.367
R308 B.n155 B.n154 163.367
R309 B.n155 B.n96 163.367
R310 B.n159 B.n96 163.367
R311 B.n160 B.n159 163.367
R312 B.n161 B.n160 163.367
R313 B.n161 B.n94 163.367
R314 B.n165 B.n94 163.367
R315 B.n166 B.n165 163.367
R316 B.n167 B.n166 163.367
R317 B.n167 B.n92 163.367
R318 B.n171 B.n92 163.367
R319 B.n172 B.n171 163.367
R320 B.n173 B.n172 163.367
R321 B.n173 B.n90 163.367
R322 B.n177 B.n90 163.367
R323 B.n178 B.n177 163.367
R324 B.n178 B.n86 163.367
R325 B.n182 B.n86 163.367
R326 B.n183 B.n182 163.367
R327 B.n184 B.n183 163.367
R328 B.n184 B.n84 163.367
R329 B.n188 B.n84 163.367
R330 B.n189 B.n188 163.367
R331 B.n190 B.n189 163.367
R332 B.n190 B.n80 163.367
R333 B.n195 B.n80 163.367
R334 B.n196 B.n195 163.367
R335 B.n197 B.n196 163.367
R336 B.n197 B.n78 163.367
R337 B.n201 B.n78 163.367
R338 B.n202 B.n201 163.367
R339 B.n203 B.n202 163.367
R340 B.n203 B.n76 163.367
R341 B.n207 B.n76 163.367
R342 B.n208 B.n207 163.367
R343 B.n209 B.n208 163.367
R344 B.n209 B.n74 163.367
R345 B.n213 B.n74 163.367
R346 B.n214 B.n213 163.367
R347 B.n215 B.n214 163.367
R348 B.n215 B.n72 163.367
R349 B.n219 B.n72 163.367
R350 B.n220 B.n219 163.367
R351 B.n221 B.n220 163.367
R352 B.n221 B.n70 163.367
R353 B.n225 B.n70 163.367
R354 B.n227 B.n226 163.367
R355 B.n227 B.n68 163.367
R356 B.n231 B.n68 163.367
R357 B.n232 B.n231 163.367
R358 B.n233 B.n232 163.367
R359 B.n233 B.n66 163.367
R360 B.n237 B.n66 163.367
R361 B.n238 B.n237 163.367
R362 B.n239 B.n238 163.367
R363 B.n239 B.n64 163.367
R364 B.n243 B.n64 163.367
R365 B.n244 B.n243 163.367
R366 B.n245 B.n244 163.367
R367 B.n245 B.n62 163.367
R368 B.n249 B.n62 163.367
R369 B.n250 B.n249 163.367
R370 B.n251 B.n250 163.367
R371 B.n251 B.n60 163.367
R372 B.n255 B.n60 163.367
R373 B.n256 B.n255 163.367
R374 B.n257 B.n256 163.367
R375 B.n257 B.n58 163.367
R376 B.n261 B.n58 163.367
R377 B.n262 B.n261 163.367
R378 B.n263 B.n262 163.367
R379 B.n263 B.n56 163.367
R380 B.n267 B.n56 163.367
R381 B.n268 B.n267 163.367
R382 B.n269 B.n268 163.367
R383 B.n269 B.n54 163.367
R384 B.n273 B.n54 163.367
R385 B.n274 B.n273 163.367
R386 B.n275 B.n274 163.367
R387 B.n275 B.n52 163.367
R388 B.n279 B.n52 163.367
R389 B.n280 B.n279 163.367
R390 B.n281 B.n280 163.367
R391 B.n281 B.n50 163.367
R392 B.n285 B.n50 163.367
R393 B.n286 B.n285 163.367
R394 B.n287 B.n286 163.367
R395 B.n287 B.n48 163.367
R396 B.n291 B.n48 163.367
R397 B.n292 B.n291 163.367
R398 B.n293 B.n292 163.367
R399 B.n293 B.n46 163.367
R400 B.n297 B.n46 163.367
R401 B.n298 B.n297 163.367
R402 B.n377 B.n376 163.367
R403 B.n376 B.n15 163.367
R404 B.n372 B.n15 163.367
R405 B.n372 B.n371 163.367
R406 B.n371 B.n370 163.367
R407 B.n370 B.n17 163.367
R408 B.n366 B.n17 163.367
R409 B.n366 B.n365 163.367
R410 B.n365 B.n364 163.367
R411 B.n364 B.n19 163.367
R412 B.n360 B.n19 163.367
R413 B.n360 B.n359 163.367
R414 B.n359 B.n358 163.367
R415 B.n358 B.n21 163.367
R416 B.n354 B.n21 163.367
R417 B.n354 B.n353 163.367
R418 B.n353 B.n352 163.367
R419 B.n352 B.n23 163.367
R420 B.n348 B.n23 163.367
R421 B.n348 B.n347 163.367
R422 B.n347 B.n346 163.367
R423 B.n346 B.n25 163.367
R424 B.n342 B.n25 163.367
R425 B.n342 B.n341 163.367
R426 B.n341 B.n340 163.367
R427 B.n340 B.n30 163.367
R428 B.n336 B.n30 163.367
R429 B.n336 B.n335 163.367
R430 B.n335 B.n334 163.367
R431 B.n334 B.n32 163.367
R432 B.n329 B.n32 163.367
R433 B.n329 B.n328 163.367
R434 B.n328 B.n327 163.367
R435 B.n327 B.n36 163.367
R436 B.n323 B.n36 163.367
R437 B.n323 B.n322 163.367
R438 B.n322 B.n321 163.367
R439 B.n321 B.n38 163.367
R440 B.n317 B.n38 163.367
R441 B.n317 B.n316 163.367
R442 B.n316 B.n315 163.367
R443 B.n315 B.n40 163.367
R444 B.n311 B.n40 163.367
R445 B.n311 B.n310 163.367
R446 B.n310 B.n309 163.367
R447 B.n309 B.n42 163.367
R448 B.n305 B.n42 163.367
R449 B.n305 B.n304 163.367
R450 B.n304 B.n303 163.367
R451 B.n303 B.n44 163.367
R452 B.n299 B.n44 163.367
R453 B.n81 B.t2 155.544
R454 B.n33 B.t10 155.544
R455 B.n87 B.t8 155.541
R456 B.n26 B.t4 155.541
R457 B.n82 B.t1 120.442
R458 B.n34 B.t11 120.442
R459 B.n88 B.t7 120.438
R460 B.n27 B.t5 120.438
R461 B.n193 B.n82 59.5399
R462 B.n89 B.n88 59.5399
R463 B.n28 B.n27 59.5399
R464 B.n331 B.n34 59.5399
R465 B.n82 B.n81 35.1035
R466 B.n88 B.n87 35.1035
R467 B.n27 B.n26 35.1035
R468 B.n34 B.n33 35.1035
R469 B.n379 B.n14 33.5615
R470 B.n300 B.n45 33.5615
R471 B.n224 B.n69 33.5615
R472 B.n146 B.n145 33.5615
R473 B B.n415 18.0485
R474 B.n375 B.n14 10.6151
R475 B.n375 B.n374 10.6151
R476 B.n374 B.n373 10.6151
R477 B.n373 B.n16 10.6151
R478 B.n369 B.n16 10.6151
R479 B.n369 B.n368 10.6151
R480 B.n368 B.n367 10.6151
R481 B.n367 B.n18 10.6151
R482 B.n363 B.n18 10.6151
R483 B.n363 B.n362 10.6151
R484 B.n362 B.n361 10.6151
R485 B.n361 B.n20 10.6151
R486 B.n357 B.n20 10.6151
R487 B.n357 B.n356 10.6151
R488 B.n356 B.n355 10.6151
R489 B.n355 B.n22 10.6151
R490 B.n351 B.n22 10.6151
R491 B.n351 B.n350 10.6151
R492 B.n350 B.n349 10.6151
R493 B.n349 B.n24 10.6151
R494 B.n345 B.n344 10.6151
R495 B.n344 B.n343 10.6151
R496 B.n343 B.n29 10.6151
R497 B.n339 B.n29 10.6151
R498 B.n339 B.n338 10.6151
R499 B.n338 B.n337 10.6151
R500 B.n337 B.n31 10.6151
R501 B.n333 B.n31 10.6151
R502 B.n333 B.n332 10.6151
R503 B.n330 B.n35 10.6151
R504 B.n326 B.n35 10.6151
R505 B.n326 B.n325 10.6151
R506 B.n325 B.n324 10.6151
R507 B.n324 B.n37 10.6151
R508 B.n320 B.n37 10.6151
R509 B.n320 B.n319 10.6151
R510 B.n319 B.n318 10.6151
R511 B.n318 B.n39 10.6151
R512 B.n314 B.n39 10.6151
R513 B.n314 B.n313 10.6151
R514 B.n313 B.n312 10.6151
R515 B.n312 B.n41 10.6151
R516 B.n308 B.n41 10.6151
R517 B.n308 B.n307 10.6151
R518 B.n307 B.n306 10.6151
R519 B.n306 B.n43 10.6151
R520 B.n302 B.n43 10.6151
R521 B.n302 B.n301 10.6151
R522 B.n301 B.n300 10.6151
R523 B.n228 B.n69 10.6151
R524 B.n229 B.n228 10.6151
R525 B.n230 B.n229 10.6151
R526 B.n230 B.n67 10.6151
R527 B.n234 B.n67 10.6151
R528 B.n235 B.n234 10.6151
R529 B.n236 B.n235 10.6151
R530 B.n236 B.n65 10.6151
R531 B.n240 B.n65 10.6151
R532 B.n241 B.n240 10.6151
R533 B.n242 B.n241 10.6151
R534 B.n242 B.n63 10.6151
R535 B.n246 B.n63 10.6151
R536 B.n247 B.n246 10.6151
R537 B.n248 B.n247 10.6151
R538 B.n248 B.n61 10.6151
R539 B.n252 B.n61 10.6151
R540 B.n253 B.n252 10.6151
R541 B.n254 B.n253 10.6151
R542 B.n254 B.n59 10.6151
R543 B.n258 B.n59 10.6151
R544 B.n259 B.n258 10.6151
R545 B.n260 B.n259 10.6151
R546 B.n260 B.n57 10.6151
R547 B.n264 B.n57 10.6151
R548 B.n265 B.n264 10.6151
R549 B.n266 B.n265 10.6151
R550 B.n266 B.n55 10.6151
R551 B.n270 B.n55 10.6151
R552 B.n271 B.n270 10.6151
R553 B.n272 B.n271 10.6151
R554 B.n272 B.n53 10.6151
R555 B.n276 B.n53 10.6151
R556 B.n277 B.n276 10.6151
R557 B.n278 B.n277 10.6151
R558 B.n278 B.n51 10.6151
R559 B.n282 B.n51 10.6151
R560 B.n283 B.n282 10.6151
R561 B.n284 B.n283 10.6151
R562 B.n284 B.n49 10.6151
R563 B.n288 B.n49 10.6151
R564 B.n289 B.n288 10.6151
R565 B.n290 B.n289 10.6151
R566 B.n290 B.n47 10.6151
R567 B.n294 B.n47 10.6151
R568 B.n295 B.n294 10.6151
R569 B.n296 B.n295 10.6151
R570 B.n296 B.n45 10.6151
R571 B.n146 B.n99 10.6151
R572 B.n150 B.n99 10.6151
R573 B.n151 B.n150 10.6151
R574 B.n152 B.n151 10.6151
R575 B.n152 B.n97 10.6151
R576 B.n156 B.n97 10.6151
R577 B.n157 B.n156 10.6151
R578 B.n158 B.n157 10.6151
R579 B.n158 B.n95 10.6151
R580 B.n162 B.n95 10.6151
R581 B.n163 B.n162 10.6151
R582 B.n164 B.n163 10.6151
R583 B.n164 B.n93 10.6151
R584 B.n168 B.n93 10.6151
R585 B.n169 B.n168 10.6151
R586 B.n170 B.n169 10.6151
R587 B.n170 B.n91 10.6151
R588 B.n174 B.n91 10.6151
R589 B.n175 B.n174 10.6151
R590 B.n176 B.n175 10.6151
R591 B.n180 B.n179 10.6151
R592 B.n181 B.n180 10.6151
R593 B.n181 B.n85 10.6151
R594 B.n185 B.n85 10.6151
R595 B.n186 B.n185 10.6151
R596 B.n187 B.n186 10.6151
R597 B.n187 B.n83 10.6151
R598 B.n191 B.n83 10.6151
R599 B.n192 B.n191 10.6151
R600 B.n194 B.n79 10.6151
R601 B.n198 B.n79 10.6151
R602 B.n199 B.n198 10.6151
R603 B.n200 B.n199 10.6151
R604 B.n200 B.n77 10.6151
R605 B.n204 B.n77 10.6151
R606 B.n205 B.n204 10.6151
R607 B.n206 B.n205 10.6151
R608 B.n206 B.n75 10.6151
R609 B.n210 B.n75 10.6151
R610 B.n211 B.n210 10.6151
R611 B.n212 B.n211 10.6151
R612 B.n212 B.n73 10.6151
R613 B.n216 B.n73 10.6151
R614 B.n217 B.n216 10.6151
R615 B.n218 B.n217 10.6151
R616 B.n218 B.n71 10.6151
R617 B.n222 B.n71 10.6151
R618 B.n223 B.n222 10.6151
R619 B.n224 B.n223 10.6151
R620 B.n145 B.n144 10.6151
R621 B.n144 B.n101 10.6151
R622 B.n140 B.n101 10.6151
R623 B.n140 B.n139 10.6151
R624 B.n139 B.n138 10.6151
R625 B.n138 B.n103 10.6151
R626 B.n134 B.n103 10.6151
R627 B.n134 B.n133 10.6151
R628 B.n133 B.n132 10.6151
R629 B.n132 B.n105 10.6151
R630 B.n128 B.n105 10.6151
R631 B.n128 B.n127 10.6151
R632 B.n127 B.n126 10.6151
R633 B.n126 B.n107 10.6151
R634 B.n122 B.n107 10.6151
R635 B.n122 B.n121 10.6151
R636 B.n121 B.n120 10.6151
R637 B.n120 B.n109 10.6151
R638 B.n116 B.n109 10.6151
R639 B.n116 B.n115 10.6151
R640 B.n115 B.n114 10.6151
R641 B.n114 B.n111 10.6151
R642 B.n111 B.n0 10.6151
R643 B.n411 B.n1 10.6151
R644 B.n411 B.n410 10.6151
R645 B.n410 B.n409 10.6151
R646 B.n409 B.n4 10.6151
R647 B.n405 B.n4 10.6151
R648 B.n405 B.n404 10.6151
R649 B.n404 B.n403 10.6151
R650 B.n403 B.n6 10.6151
R651 B.n399 B.n6 10.6151
R652 B.n399 B.n398 10.6151
R653 B.n398 B.n397 10.6151
R654 B.n397 B.n8 10.6151
R655 B.n393 B.n8 10.6151
R656 B.n393 B.n392 10.6151
R657 B.n392 B.n391 10.6151
R658 B.n391 B.n10 10.6151
R659 B.n387 B.n10 10.6151
R660 B.n387 B.n386 10.6151
R661 B.n386 B.n385 10.6151
R662 B.n385 B.n12 10.6151
R663 B.n381 B.n12 10.6151
R664 B.n381 B.n380 10.6151
R665 B.n380 B.n379 10.6151
R666 B.n28 B.n24 9.36635
R667 B.n331 B.n330 9.36635
R668 B.n176 B.n89 9.36635
R669 B.n194 B.n193 9.36635
R670 B.n415 B.n0 2.81026
R671 B.n415 B.n1 2.81026
R672 B.n345 B.n28 1.24928
R673 B.n332 B.n331 1.24928
R674 B.n179 B.n89 1.24928
R675 B.n193 B.n192 1.24928
R676 VN.n0 VN.t2 118.626
R677 VN.n1 VN.t1 118.626
R678 VN.n0 VN.t0 118.312
R679 VN.n1 VN.t3 118.312
R680 VN VN.n1 51.0103
R681 VN VN.n0 13.1353
R682 VDD2.n2 VDD2.n0 136.117
R683 VDD2.n2 VDD2.n1 103.35
R684 VDD2.n1 VDD2.t0 6.41174
R685 VDD2.n1 VDD2.t2 6.41174
R686 VDD2.n0 VDD2.t1 6.41174
R687 VDD2.n0 VDD2.t3 6.41174
R688 VDD2 VDD2.n2 0.0586897
C0 VN w_n2056_n1982# 3.14659f
C1 VP B 1.24905f
C2 VDD2 B 0.911759f
C3 B VTAIL 2.26809f
C4 VDD1 w_n2056_n1982# 1.04706f
C5 B w_n2056_n1982# 5.93033f
C6 VDD1 VN 0.148105f
C7 VN B 0.820413f
C8 VDD2 VP 0.327204f
C9 VP VTAIL 2.06286f
C10 VDD2 VTAIL 3.49035f
C11 VDD1 B 0.877807f
C12 VP w_n2056_n1982# 3.40798f
C13 VDD2 w_n2056_n1982# 1.07792f
C14 w_n2056_n1982# VTAIL 2.35936f
C15 VN VP 4.10219f
C16 VDD2 VN 1.93514f
C17 VN VTAIL 2.04876f
C18 VDD1 VP 2.10969f
C19 VDD1 VDD2 0.75481f
C20 VDD1 VTAIL 3.44365f
C21 VDD2 VSUBS 0.552442f
C22 VDD1 VSUBS 4.104718f
C23 VTAIL VSUBS 0.561838f
C24 VN VSUBS 4.36444f
C25 VP VSUBS 1.323712f
C26 B VSUBS 2.593269f
C27 w_n2056_n1982# VSUBS 51.0464f
C28 VDD2.t1 VSUBS 0.070001f
C29 VDD2.t3 VSUBS 0.070001f
C30 VDD2.n0 VSUBS 0.653015f
C31 VDD2.t0 VSUBS 0.070001f
C32 VDD2.t2 VSUBS 0.070001f
C33 VDD2.n1 VSUBS 0.442899f
C34 VDD2.n2 VSUBS 2.03248f
C35 VN.t2 VSUBS 1.01817f
C36 VN.t0 VSUBS 1.01674f
C37 VN.n0 VSUBS 0.787602f
C38 VN.t1 VSUBS 1.01817f
C39 VN.t3 VSUBS 1.01674f
C40 VN.n1 VSUBS 2.09197f
C41 B.n0 VSUBS 0.005801f
C42 B.n1 VSUBS 0.005801f
C43 B.n2 VSUBS 0.009174f
C44 B.n3 VSUBS 0.009174f
C45 B.n4 VSUBS 0.009174f
C46 B.n5 VSUBS 0.009174f
C47 B.n6 VSUBS 0.009174f
C48 B.n7 VSUBS 0.009174f
C49 B.n8 VSUBS 0.009174f
C50 B.n9 VSUBS 0.009174f
C51 B.n10 VSUBS 0.009174f
C52 B.n11 VSUBS 0.009174f
C53 B.n12 VSUBS 0.009174f
C54 B.n13 VSUBS 0.009174f
C55 B.n14 VSUBS 0.022409f
C56 B.n15 VSUBS 0.009174f
C57 B.n16 VSUBS 0.009174f
C58 B.n17 VSUBS 0.009174f
C59 B.n18 VSUBS 0.009174f
C60 B.n19 VSUBS 0.009174f
C61 B.n20 VSUBS 0.009174f
C62 B.n21 VSUBS 0.009174f
C63 B.n22 VSUBS 0.009174f
C64 B.n23 VSUBS 0.009174f
C65 B.n24 VSUBS 0.008635f
C66 B.n25 VSUBS 0.009174f
C67 B.t5 VSUBS 0.185923f
C68 B.t4 VSUBS 0.202434f
C69 B.t3 VSUBS 0.454956f
C70 B.n26 VSUBS 0.12234f
C71 B.n27 VSUBS 0.086242f
C72 B.n28 VSUBS 0.021256f
C73 B.n29 VSUBS 0.009174f
C74 B.n30 VSUBS 0.009174f
C75 B.n31 VSUBS 0.009174f
C76 B.n32 VSUBS 0.009174f
C77 B.t11 VSUBS 0.185923f
C78 B.t10 VSUBS 0.202433f
C79 B.t9 VSUBS 0.454956f
C80 B.n33 VSUBS 0.12234f
C81 B.n34 VSUBS 0.086243f
C82 B.n35 VSUBS 0.009174f
C83 B.n36 VSUBS 0.009174f
C84 B.n37 VSUBS 0.009174f
C85 B.n38 VSUBS 0.009174f
C86 B.n39 VSUBS 0.009174f
C87 B.n40 VSUBS 0.009174f
C88 B.n41 VSUBS 0.009174f
C89 B.n42 VSUBS 0.009174f
C90 B.n43 VSUBS 0.009174f
C91 B.n44 VSUBS 0.009174f
C92 B.n45 VSUBS 0.022358f
C93 B.n46 VSUBS 0.009174f
C94 B.n47 VSUBS 0.009174f
C95 B.n48 VSUBS 0.009174f
C96 B.n49 VSUBS 0.009174f
C97 B.n50 VSUBS 0.009174f
C98 B.n51 VSUBS 0.009174f
C99 B.n52 VSUBS 0.009174f
C100 B.n53 VSUBS 0.009174f
C101 B.n54 VSUBS 0.009174f
C102 B.n55 VSUBS 0.009174f
C103 B.n56 VSUBS 0.009174f
C104 B.n57 VSUBS 0.009174f
C105 B.n58 VSUBS 0.009174f
C106 B.n59 VSUBS 0.009174f
C107 B.n60 VSUBS 0.009174f
C108 B.n61 VSUBS 0.009174f
C109 B.n62 VSUBS 0.009174f
C110 B.n63 VSUBS 0.009174f
C111 B.n64 VSUBS 0.009174f
C112 B.n65 VSUBS 0.009174f
C113 B.n66 VSUBS 0.009174f
C114 B.n67 VSUBS 0.009174f
C115 B.n68 VSUBS 0.009174f
C116 B.n69 VSUBS 0.021303f
C117 B.n70 VSUBS 0.009174f
C118 B.n71 VSUBS 0.009174f
C119 B.n72 VSUBS 0.009174f
C120 B.n73 VSUBS 0.009174f
C121 B.n74 VSUBS 0.009174f
C122 B.n75 VSUBS 0.009174f
C123 B.n76 VSUBS 0.009174f
C124 B.n77 VSUBS 0.009174f
C125 B.n78 VSUBS 0.009174f
C126 B.n79 VSUBS 0.009174f
C127 B.n80 VSUBS 0.009174f
C128 B.t1 VSUBS 0.185923f
C129 B.t2 VSUBS 0.202433f
C130 B.t0 VSUBS 0.454956f
C131 B.n81 VSUBS 0.12234f
C132 B.n82 VSUBS 0.086243f
C133 B.n83 VSUBS 0.009174f
C134 B.n84 VSUBS 0.009174f
C135 B.n85 VSUBS 0.009174f
C136 B.n86 VSUBS 0.009174f
C137 B.t7 VSUBS 0.185923f
C138 B.t8 VSUBS 0.202434f
C139 B.t6 VSUBS 0.454956f
C140 B.n87 VSUBS 0.12234f
C141 B.n88 VSUBS 0.086242f
C142 B.n89 VSUBS 0.021256f
C143 B.n90 VSUBS 0.009174f
C144 B.n91 VSUBS 0.009174f
C145 B.n92 VSUBS 0.009174f
C146 B.n93 VSUBS 0.009174f
C147 B.n94 VSUBS 0.009174f
C148 B.n95 VSUBS 0.009174f
C149 B.n96 VSUBS 0.009174f
C150 B.n97 VSUBS 0.009174f
C151 B.n98 VSUBS 0.009174f
C152 B.n99 VSUBS 0.009174f
C153 B.n100 VSUBS 0.021303f
C154 B.n101 VSUBS 0.009174f
C155 B.n102 VSUBS 0.009174f
C156 B.n103 VSUBS 0.009174f
C157 B.n104 VSUBS 0.009174f
C158 B.n105 VSUBS 0.009174f
C159 B.n106 VSUBS 0.009174f
C160 B.n107 VSUBS 0.009174f
C161 B.n108 VSUBS 0.009174f
C162 B.n109 VSUBS 0.009174f
C163 B.n110 VSUBS 0.009174f
C164 B.n111 VSUBS 0.009174f
C165 B.n112 VSUBS 0.009174f
C166 B.n113 VSUBS 0.009174f
C167 B.n114 VSUBS 0.009174f
C168 B.n115 VSUBS 0.009174f
C169 B.n116 VSUBS 0.009174f
C170 B.n117 VSUBS 0.009174f
C171 B.n118 VSUBS 0.009174f
C172 B.n119 VSUBS 0.009174f
C173 B.n120 VSUBS 0.009174f
C174 B.n121 VSUBS 0.009174f
C175 B.n122 VSUBS 0.009174f
C176 B.n123 VSUBS 0.009174f
C177 B.n124 VSUBS 0.009174f
C178 B.n125 VSUBS 0.009174f
C179 B.n126 VSUBS 0.009174f
C180 B.n127 VSUBS 0.009174f
C181 B.n128 VSUBS 0.009174f
C182 B.n129 VSUBS 0.009174f
C183 B.n130 VSUBS 0.009174f
C184 B.n131 VSUBS 0.009174f
C185 B.n132 VSUBS 0.009174f
C186 B.n133 VSUBS 0.009174f
C187 B.n134 VSUBS 0.009174f
C188 B.n135 VSUBS 0.009174f
C189 B.n136 VSUBS 0.009174f
C190 B.n137 VSUBS 0.009174f
C191 B.n138 VSUBS 0.009174f
C192 B.n139 VSUBS 0.009174f
C193 B.n140 VSUBS 0.009174f
C194 B.n141 VSUBS 0.009174f
C195 B.n142 VSUBS 0.009174f
C196 B.n143 VSUBS 0.009174f
C197 B.n144 VSUBS 0.009174f
C198 B.n145 VSUBS 0.021303f
C199 B.n146 VSUBS 0.022409f
C200 B.n147 VSUBS 0.022409f
C201 B.n148 VSUBS 0.009174f
C202 B.n149 VSUBS 0.009174f
C203 B.n150 VSUBS 0.009174f
C204 B.n151 VSUBS 0.009174f
C205 B.n152 VSUBS 0.009174f
C206 B.n153 VSUBS 0.009174f
C207 B.n154 VSUBS 0.009174f
C208 B.n155 VSUBS 0.009174f
C209 B.n156 VSUBS 0.009174f
C210 B.n157 VSUBS 0.009174f
C211 B.n158 VSUBS 0.009174f
C212 B.n159 VSUBS 0.009174f
C213 B.n160 VSUBS 0.009174f
C214 B.n161 VSUBS 0.009174f
C215 B.n162 VSUBS 0.009174f
C216 B.n163 VSUBS 0.009174f
C217 B.n164 VSUBS 0.009174f
C218 B.n165 VSUBS 0.009174f
C219 B.n166 VSUBS 0.009174f
C220 B.n167 VSUBS 0.009174f
C221 B.n168 VSUBS 0.009174f
C222 B.n169 VSUBS 0.009174f
C223 B.n170 VSUBS 0.009174f
C224 B.n171 VSUBS 0.009174f
C225 B.n172 VSUBS 0.009174f
C226 B.n173 VSUBS 0.009174f
C227 B.n174 VSUBS 0.009174f
C228 B.n175 VSUBS 0.009174f
C229 B.n176 VSUBS 0.008635f
C230 B.n177 VSUBS 0.009174f
C231 B.n178 VSUBS 0.009174f
C232 B.n179 VSUBS 0.005127f
C233 B.n180 VSUBS 0.009174f
C234 B.n181 VSUBS 0.009174f
C235 B.n182 VSUBS 0.009174f
C236 B.n183 VSUBS 0.009174f
C237 B.n184 VSUBS 0.009174f
C238 B.n185 VSUBS 0.009174f
C239 B.n186 VSUBS 0.009174f
C240 B.n187 VSUBS 0.009174f
C241 B.n188 VSUBS 0.009174f
C242 B.n189 VSUBS 0.009174f
C243 B.n190 VSUBS 0.009174f
C244 B.n191 VSUBS 0.009174f
C245 B.n192 VSUBS 0.005127f
C246 B.n193 VSUBS 0.021256f
C247 B.n194 VSUBS 0.008635f
C248 B.n195 VSUBS 0.009174f
C249 B.n196 VSUBS 0.009174f
C250 B.n197 VSUBS 0.009174f
C251 B.n198 VSUBS 0.009174f
C252 B.n199 VSUBS 0.009174f
C253 B.n200 VSUBS 0.009174f
C254 B.n201 VSUBS 0.009174f
C255 B.n202 VSUBS 0.009174f
C256 B.n203 VSUBS 0.009174f
C257 B.n204 VSUBS 0.009174f
C258 B.n205 VSUBS 0.009174f
C259 B.n206 VSUBS 0.009174f
C260 B.n207 VSUBS 0.009174f
C261 B.n208 VSUBS 0.009174f
C262 B.n209 VSUBS 0.009174f
C263 B.n210 VSUBS 0.009174f
C264 B.n211 VSUBS 0.009174f
C265 B.n212 VSUBS 0.009174f
C266 B.n213 VSUBS 0.009174f
C267 B.n214 VSUBS 0.009174f
C268 B.n215 VSUBS 0.009174f
C269 B.n216 VSUBS 0.009174f
C270 B.n217 VSUBS 0.009174f
C271 B.n218 VSUBS 0.009174f
C272 B.n219 VSUBS 0.009174f
C273 B.n220 VSUBS 0.009174f
C274 B.n221 VSUBS 0.009174f
C275 B.n222 VSUBS 0.009174f
C276 B.n223 VSUBS 0.009174f
C277 B.n224 VSUBS 0.022409f
C278 B.n225 VSUBS 0.022409f
C279 B.n226 VSUBS 0.021303f
C280 B.n227 VSUBS 0.009174f
C281 B.n228 VSUBS 0.009174f
C282 B.n229 VSUBS 0.009174f
C283 B.n230 VSUBS 0.009174f
C284 B.n231 VSUBS 0.009174f
C285 B.n232 VSUBS 0.009174f
C286 B.n233 VSUBS 0.009174f
C287 B.n234 VSUBS 0.009174f
C288 B.n235 VSUBS 0.009174f
C289 B.n236 VSUBS 0.009174f
C290 B.n237 VSUBS 0.009174f
C291 B.n238 VSUBS 0.009174f
C292 B.n239 VSUBS 0.009174f
C293 B.n240 VSUBS 0.009174f
C294 B.n241 VSUBS 0.009174f
C295 B.n242 VSUBS 0.009174f
C296 B.n243 VSUBS 0.009174f
C297 B.n244 VSUBS 0.009174f
C298 B.n245 VSUBS 0.009174f
C299 B.n246 VSUBS 0.009174f
C300 B.n247 VSUBS 0.009174f
C301 B.n248 VSUBS 0.009174f
C302 B.n249 VSUBS 0.009174f
C303 B.n250 VSUBS 0.009174f
C304 B.n251 VSUBS 0.009174f
C305 B.n252 VSUBS 0.009174f
C306 B.n253 VSUBS 0.009174f
C307 B.n254 VSUBS 0.009174f
C308 B.n255 VSUBS 0.009174f
C309 B.n256 VSUBS 0.009174f
C310 B.n257 VSUBS 0.009174f
C311 B.n258 VSUBS 0.009174f
C312 B.n259 VSUBS 0.009174f
C313 B.n260 VSUBS 0.009174f
C314 B.n261 VSUBS 0.009174f
C315 B.n262 VSUBS 0.009174f
C316 B.n263 VSUBS 0.009174f
C317 B.n264 VSUBS 0.009174f
C318 B.n265 VSUBS 0.009174f
C319 B.n266 VSUBS 0.009174f
C320 B.n267 VSUBS 0.009174f
C321 B.n268 VSUBS 0.009174f
C322 B.n269 VSUBS 0.009174f
C323 B.n270 VSUBS 0.009174f
C324 B.n271 VSUBS 0.009174f
C325 B.n272 VSUBS 0.009174f
C326 B.n273 VSUBS 0.009174f
C327 B.n274 VSUBS 0.009174f
C328 B.n275 VSUBS 0.009174f
C329 B.n276 VSUBS 0.009174f
C330 B.n277 VSUBS 0.009174f
C331 B.n278 VSUBS 0.009174f
C332 B.n279 VSUBS 0.009174f
C333 B.n280 VSUBS 0.009174f
C334 B.n281 VSUBS 0.009174f
C335 B.n282 VSUBS 0.009174f
C336 B.n283 VSUBS 0.009174f
C337 B.n284 VSUBS 0.009174f
C338 B.n285 VSUBS 0.009174f
C339 B.n286 VSUBS 0.009174f
C340 B.n287 VSUBS 0.009174f
C341 B.n288 VSUBS 0.009174f
C342 B.n289 VSUBS 0.009174f
C343 B.n290 VSUBS 0.009174f
C344 B.n291 VSUBS 0.009174f
C345 B.n292 VSUBS 0.009174f
C346 B.n293 VSUBS 0.009174f
C347 B.n294 VSUBS 0.009174f
C348 B.n295 VSUBS 0.009174f
C349 B.n296 VSUBS 0.009174f
C350 B.n297 VSUBS 0.009174f
C351 B.n298 VSUBS 0.021303f
C352 B.n299 VSUBS 0.022409f
C353 B.n300 VSUBS 0.021355f
C354 B.n301 VSUBS 0.009174f
C355 B.n302 VSUBS 0.009174f
C356 B.n303 VSUBS 0.009174f
C357 B.n304 VSUBS 0.009174f
C358 B.n305 VSUBS 0.009174f
C359 B.n306 VSUBS 0.009174f
C360 B.n307 VSUBS 0.009174f
C361 B.n308 VSUBS 0.009174f
C362 B.n309 VSUBS 0.009174f
C363 B.n310 VSUBS 0.009174f
C364 B.n311 VSUBS 0.009174f
C365 B.n312 VSUBS 0.009174f
C366 B.n313 VSUBS 0.009174f
C367 B.n314 VSUBS 0.009174f
C368 B.n315 VSUBS 0.009174f
C369 B.n316 VSUBS 0.009174f
C370 B.n317 VSUBS 0.009174f
C371 B.n318 VSUBS 0.009174f
C372 B.n319 VSUBS 0.009174f
C373 B.n320 VSUBS 0.009174f
C374 B.n321 VSUBS 0.009174f
C375 B.n322 VSUBS 0.009174f
C376 B.n323 VSUBS 0.009174f
C377 B.n324 VSUBS 0.009174f
C378 B.n325 VSUBS 0.009174f
C379 B.n326 VSUBS 0.009174f
C380 B.n327 VSUBS 0.009174f
C381 B.n328 VSUBS 0.009174f
C382 B.n329 VSUBS 0.009174f
C383 B.n330 VSUBS 0.008635f
C384 B.n331 VSUBS 0.021256f
C385 B.n332 VSUBS 0.005127f
C386 B.n333 VSUBS 0.009174f
C387 B.n334 VSUBS 0.009174f
C388 B.n335 VSUBS 0.009174f
C389 B.n336 VSUBS 0.009174f
C390 B.n337 VSUBS 0.009174f
C391 B.n338 VSUBS 0.009174f
C392 B.n339 VSUBS 0.009174f
C393 B.n340 VSUBS 0.009174f
C394 B.n341 VSUBS 0.009174f
C395 B.n342 VSUBS 0.009174f
C396 B.n343 VSUBS 0.009174f
C397 B.n344 VSUBS 0.009174f
C398 B.n345 VSUBS 0.005127f
C399 B.n346 VSUBS 0.009174f
C400 B.n347 VSUBS 0.009174f
C401 B.n348 VSUBS 0.009174f
C402 B.n349 VSUBS 0.009174f
C403 B.n350 VSUBS 0.009174f
C404 B.n351 VSUBS 0.009174f
C405 B.n352 VSUBS 0.009174f
C406 B.n353 VSUBS 0.009174f
C407 B.n354 VSUBS 0.009174f
C408 B.n355 VSUBS 0.009174f
C409 B.n356 VSUBS 0.009174f
C410 B.n357 VSUBS 0.009174f
C411 B.n358 VSUBS 0.009174f
C412 B.n359 VSUBS 0.009174f
C413 B.n360 VSUBS 0.009174f
C414 B.n361 VSUBS 0.009174f
C415 B.n362 VSUBS 0.009174f
C416 B.n363 VSUBS 0.009174f
C417 B.n364 VSUBS 0.009174f
C418 B.n365 VSUBS 0.009174f
C419 B.n366 VSUBS 0.009174f
C420 B.n367 VSUBS 0.009174f
C421 B.n368 VSUBS 0.009174f
C422 B.n369 VSUBS 0.009174f
C423 B.n370 VSUBS 0.009174f
C424 B.n371 VSUBS 0.009174f
C425 B.n372 VSUBS 0.009174f
C426 B.n373 VSUBS 0.009174f
C427 B.n374 VSUBS 0.009174f
C428 B.n375 VSUBS 0.009174f
C429 B.n376 VSUBS 0.009174f
C430 B.n377 VSUBS 0.022409f
C431 B.n378 VSUBS 0.021303f
C432 B.n379 VSUBS 0.021303f
C433 B.n380 VSUBS 0.009174f
C434 B.n381 VSUBS 0.009174f
C435 B.n382 VSUBS 0.009174f
C436 B.n383 VSUBS 0.009174f
C437 B.n384 VSUBS 0.009174f
C438 B.n385 VSUBS 0.009174f
C439 B.n386 VSUBS 0.009174f
C440 B.n387 VSUBS 0.009174f
C441 B.n388 VSUBS 0.009174f
C442 B.n389 VSUBS 0.009174f
C443 B.n390 VSUBS 0.009174f
C444 B.n391 VSUBS 0.009174f
C445 B.n392 VSUBS 0.009174f
C446 B.n393 VSUBS 0.009174f
C447 B.n394 VSUBS 0.009174f
C448 B.n395 VSUBS 0.009174f
C449 B.n396 VSUBS 0.009174f
C450 B.n397 VSUBS 0.009174f
C451 B.n398 VSUBS 0.009174f
C452 B.n399 VSUBS 0.009174f
C453 B.n400 VSUBS 0.009174f
C454 B.n401 VSUBS 0.009174f
C455 B.n402 VSUBS 0.009174f
C456 B.n403 VSUBS 0.009174f
C457 B.n404 VSUBS 0.009174f
C458 B.n405 VSUBS 0.009174f
C459 B.n406 VSUBS 0.009174f
C460 B.n407 VSUBS 0.009174f
C461 B.n408 VSUBS 0.009174f
C462 B.n409 VSUBS 0.009174f
C463 B.n410 VSUBS 0.009174f
C464 B.n411 VSUBS 0.009174f
C465 B.n412 VSUBS 0.009174f
C466 B.n413 VSUBS 0.009174f
C467 B.n414 VSUBS 0.009174f
C468 B.n415 VSUBS 0.020774f
C469 VDD1.t0 VSUBS 0.108009f
C470 VDD1.t1 VSUBS 0.108009f
C471 VDD1.n0 VSUBS 0.683702f
C472 VDD1.t2 VSUBS 0.108009f
C473 VDD1.t3 VSUBS 0.108009f
C474 VDD1.n1 VSUBS 1.02492f
C475 VTAIL.t1 VSUBS 0.849984f
C476 VTAIL.n0 VSUBS 0.626628f
C477 VTAIL.t7 VSUBS 0.849984f
C478 VTAIL.n1 VSUBS 0.689718f
C479 VTAIL.t5 VSUBS 0.849984f
C480 VTAIL.n2 VSUBS 1.53531f
C481 VTAIL.t2 VSUBS 0.849989f
C482 VTAIL.n3 VSUBS 1.53531f
C483 VTAIL.t0 VSUBS 0.849989f
C484 VTAIL.n4 VSUBS 0.689713f
C485 VTAIL.t6 VSUBS 0.849989f
C486 VTAIL.n5 VSUBS 0.689713f
C487 VTAIL.t4 VSUBS 0.849984f
C488 VTAIL.n6 VSUBS 1.53531f
C489 VTAIL.t3 VSUBS 0.849984f
C490 VTAIL.n7 VSUBS 1.46206f
C491 VP.n0 VSUBS 0.056042f
C492 VP.t0 VSUBS 1.101f
C493 VP.n1 VSUBS 0.081811f
C494 VP.t3 VSUBS 1.30356f
C495 VP.t2 VSUBS 1.30174f
C496 VP.n2 VSUBS 2.64653f
C497 VP.n3 VSUBS 2.5403f
C498 VP.t1 VSUBS 1.101f
C499 VP.n4 VSUBS 0.551539f
C500 VP.n5 VSUBS 0.068864f
C501 VP.n6 VSUBS 0.056042f
C502 VP.n7 VSUBS 0.056042f
C503 VP.n8 VSUBS 0.056042f
C504 VP.n9 VSUBS 0.081811f
C505 VP.n10 VSUBS 0.068864f
C506 VP.n11 VSUBS 0.551539f
C507 VP.n12 VSUBS 0.054645f
.ends

