* NGSPICE file created from diff_pair_sample_0601.ext - technology: sky130A

.subckt diff_pair_sample_0601 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.1
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.1
X2 VDD2.t2 VN.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.1
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.1
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.1
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=0 ps=0 w=9.79 l=2.1
X6 VDD2.t0 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.1
X7 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.1
X8 VTAIL.t4 VN.t3 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.1
X9 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.1
X10 VDD1.t1 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.61535 pd=10.12 as=3.8181 ps=20.36 w=9.79 l=2.1
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8181 pd=20.36 as=1.61535 ps=10.12 w=9.79 l=2.1
R0 VN.n0 VN.t0 148.458
R1 VN.n1 VN.t2 148.458
R2 VN.n0 VN.t1 147.911
R3 VN.n1 VN.t3 147.911
R4 VN VN.n1 50.3258
R5 VN VN.n0 6.90537
R6 VDD2.n2 VDD2.n0 104.936
R7 VDD2.n2 VDD2.n1 66.4968
R8 VDD2.n1 VDD2.t1 2.02297
R9 VDD2.n1 VDD2.t0 2.02297
R10 VDD2.n0 VDD2.t3 2.02297
R11 VDD2.n0 VDD2.t2 2.02297
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t3 51.8406
R14 VTAIL.n4 VTAIL.t5 51.8406
R15 VTAIL.n3 VTAIL.t4 51.8406
R16 VTAIL.n7 VTAIL.t6 51.8405
R17 VTAIL.n0 VTAIL.t7 51.8405
R18 VTAIL.n1 VTAIL.t0 51.8405
R19 VTAIL.n2 VTAIL.t1 51.8405
R20 VTAIL.n6 VTAIL.t2 51.8405
R21 VTAIL.n7 VTAIL.n6 22.9014
R22 VTAIL.n3 VTAIL.n2 22.9014
R23 VTAIL.n4 VTAIL.n3 2.09533
R24 VTAIL.n6 VTAIL.n5 2.09533
R25 VTAIL.n2 VTAIL.n1 2.09533
R26 VTAIL VTAIL.n0 1.1061
R27 VTAIL VTAIL.n7 0.989724
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n648 B.n647 585
R31 B.n259 B.n96 585
R32 B.n258 B.n257 585
R33 B.n256 B.n255 585
R34 B.n254 B.n253 585
R35 B.n252 B.n251 585
R36 B.n250 B.n249 585
R37 B.n248 B.n247 585
R38 B.n246 B.n245 585
R39 B.n244 B.n243 585
R40 B.n242 B.n241 585
R41 B.n240 B.n239 585
R42 B.n238 B.n237 585
R43 B.n236 B.n235 585
R44 B.n234 B.n233 585
R45 B.n232 B.n231 585
R46 B.n230 B.n229 585
R47 B.n228 B.n227 585
R48 B.n226 B.n225 585
R49 B.n224 B.n223 585
R50 B.n222 B.n221 585
R51 B.n220 B.n219 585
R52 B.n218 B.n217 585
R53 B.n216 B.n215 585
R54 B.n214 B.n213 585
R55 B.n212 B.n211 585
R56 B.n210 B.n209 585
R57 B.n208 B.n207 585
R58 B.n206 B.n205 585
R59 B.n204 B.n203 585
R60 B.n202 B.n201 585
R61 B.n200 B.n199 585
R62 B.n198 B.n197 585
R63 B.n196 B.n195 585
R64 B.n194 B.n193 585
R65 B.n191 B.n190 585
R66 B.n189 B.n188 585
R67 B.n187 B.n186 585
R68 B.n185 B.n184 585
R69 B.n183 B.n182 585
R70 B.n181 B.n180 585
R71 B.n179 B.n178 585
R72 B.n177 B.n176 585
R73 B.n175 B.n174 585
R74 B.n173 B.n172 585
R75 B.n170 B.n169 585
R76 B.n168 B.n167 585
R77 B.n166 B.n165 585
R78 B.n164 B.n163 585
R79 B.n162 B.n161 585
R80 B.n160 B.n159 585
R81 B.n158 B.n157 585
R82 B.n156 B.n155 585
R83 B.n154 B.n153 585
R84 B.n152 B.n151 585
R85 B.n150 B.n149 585
R86 B.n148 B.n147 585
R87 B.n146 B.n145 585
R88 B.n144 B.n143 585
R89 B.n142 B.n141 585
R90 B.n140 B.n139 585
R91 B.n138 B.n137 585
R92 B.n136 B.n135 585
R93 B.n134 B.n133 585
R94 B.n132 B.n131 585
R95 B.n130 B.n129 585
R96 B.n128 B.n127 585
R97 B.n126 B.n125 585
R98 B.n124 B.n123 585
R99 B.n122 B.n121 585
R100 B.n120 B.n119 585
R101 B.n118 B.n117 585
R102 B.n116 B.n115 585
R103 B.n114 B.n113 585
R104 B.n112 B.n111 585
R105 B.n110 B.n109 585
R106 B.n108 B.n107 585
R107 B.n106 B.n105 585
R108 B.n104 B.n103 585
R109 B.n102 B.n101 585
R110 B.n646 B.n56 585
R111 B.n651 B.n56 585
R112 B.n645 B.n55 585
R113 B.n652 B.n55 585
R114 B.n644 B.n643 585
R115 B.n643 B.n51 585
R116 B.n642 B.n50 585
R117 B.n658 B.n50 585
R118 B.n641 B.n49 585
R119 B.n659 B.n49 585
R120 B.n640 B.n48 585
R121 B.n660 B.n48 585
R122 B.n639 B.n638 585
R123 B.n638 B.n47 585
R124 B.n637 B.n43 585
R125 B.n666 B.n43 585
R126 B.n636 B.n42 585
R127 B.n667 B.n42 585
R128 B.n635 B.n41 585
R129 B.n668 B.n41 585
R130 B.n634 B.n633 585
R131 B.n633 B.n37 585
R132 B.n632 B.n36 585
R133 B.n674 B.n36 585
R134 B.n631 B.n35 585
R135 B.n675 B.n35 585
R136 B.n630 B.n34 585
R137 B.n676 B.n34 585
R138 B.n629 B.n628 585
R139 B.n628 B.n30 585
R140 B.n627 B.n29 585
R141 B.n682 B.n29 585
R142 B.n626 B.n28 585
R143 B.n683 B.n28 585
R144 B.n625 B.n27 585
R145 B.n684 B.n27 585
R146 B.n624 B.n623 585
R147 B.n623 B.n23 585
R148 B.n622 B.n22 585
R149 B.n690 B.n22 585
R150 B.n621 B.n21 585
R151 B.n691 B.n21 585
R152 B.n620 B.n20 585
R153 B.n692 B.n20 585
R154 B.n619 B.n618 585
R155 B.n618 B.n16 585
R156 B.n617 B.n15 585
R157 B.n698 B.n15 585
R158 B.n616 B.n14 585
R159 B.n699 B.n14 585
R160 B.n615 B.n13 585
R161 B.n700 B.n13 585
R162 B.n614 B.n613 585
R163 B.n613 B.n12 585
R164 B.n612 B.n611 585
R165 B.n612 B.n8 585
R166 B.n610 B.n7 585
R167 B.n707 B.n7 585
R168 B.n609 B.n6 585
R169 B.n708 B.n6 585
R170 B.n608 B.n5 585
R171 B.n709 B.n5 585
R172 B.n607 B.n606 585
R173 B.n606 B.n4 585
R174 B.n605 B.n260 585
R175 B.n605 B.n604 585
R176 B.n595 B.n261 585
R177 B.n262 B.n261 585
R178 B.n597 B.n596 585
R179 B.n598 B.n597 585
R180 B.n594 B.n266 585
R181 B.n270 B.n266 585
R182 B.n593 B.n592 585
R183 B.n592 B.n591 585
R184 B.n268 B.n267 585
R185 B.n269 B.n268 585
R186 B.n584 B.n583 585
R187 B.n585 B.n584 585
R188 B.n582 B.n275 585
R189 B.n275 B.n274 585
R190 B.n581 B.n580 585
R191 B.n580 B.n579 585
R192 B.n277 B.n276 585
R193 B.n278 B.n277 585
R194 B.n572 B.n571 585
R195 B.n573 B.n572 585
R196 B.n570 B.n283 585
R197 B.n283 B.n282 585
R198 B.n569 B.n568 585
R199 B.n568 B.n567 585
R200 B.n285 B.n284 585
R201 B.n286 B.n285 585
R202 B.n560 B.n559 585
R203 B.n561 B.n560 585
R204 B.n558 B.n291 585
R205 B.n291 B.n290 585
R206 B.n557 B.n556 585
R207 B.n556 B.n555 585
R208 B.n293 B.n292 585
R209 B.n294 B.n293 585
R210 B.n548 B.n547 585
R211 B.n549 B.n548 585
R212 B.n546 B.n299 585
R213 B.n299 B.n298 585
R214 B.n545 B.n544 585
R215 B.n544 B.n543 585
R216 B.n301 B.n300 585
R217 B.n536 B.n301 585
R218 B.n535 B.n534 585
R219 B.n537 B.n535 585
R220 B.n533 B.n306 585
R221 B.n306 B.n305 585
R222 B.n532 B.n531 585
R223 B.n531 B.n530 585
R224 B.n308 B.n307 585
R225 B.n309 B.n308 585
R226 B.n523 B.n522 585
R227 B.n524 B.n523 585
R228 B.n521 B.n314 585
R229 B.n314 B.n313 585
R230 B.n516 B.n515 585
R231 B.n514 B.n356 585
R232 B.n513 B.n355 585
R233 B.n518 B.n355 585
R234 B.n512 B.n511 585
R235 B.n510 B.n509 585
R236 B.n508 B.n507 585
R237 B.n506 B.n505 585
R238 B.n504 B.n503 585
R239 B.n502 B.n501 585
R240 B.n500 B.n499 585
R241 B.n498 B.n497 585
R242 B.n496 B.n495 585
R243 B.n494 B.n493 585
R244 B.n492 B.n491 585
R245 B.n490 B.n489 585
R246 B.n488 B.n487 585
R247 B.n486 B.n485 585
R248 B.n484 B.n483 585
R249 B.n482 B.n481 585
R250 B.n480 B.n479 585
R251 B.n478 B.n477 585
R252 B.n476 B.n475 585
R253 B.n474 B.n473 585
R254 B.n472 B.n471 585
R255 B.n470 B.n469 585
R256 B.n468 B.n467 585
R257 B.n466 B.n465 585
R258 B.n464 B.n463 585
R259 B.n462 B.n461 585
R260 B.n460 B.n459 585
R261 B.n458 B.n457 585
R262 B.n456 B.n455 585
R263 B.n454 B.n453 585
R264 B.n452 B.n451 585
R265 B.n450 B.n449 585
R266 B.n448 B.n447 585
R267 B.n446 B.n445 585
R268 B.n444 B.n443 585
R269 B.n442 B.n441 585
R270 B.n440 B.n439 585
R271 B.n438 B.n437 585
R272 B.n436 B.n435 585
R273 B.n434 B.n433 585
R274 B.n432 B.n431 585
R275 B.n430 B.n429 585
R276 B.n428 B.n427 585
R277 B.n426 B.n425 585
R278 B.n424 B.n423 585
R279 B.n422 B.n421 585
R280 B.n420 B.n419 585
R281 B.n418 B.n417 585
R282 B.n416 B.n415 585
R283 B.n414 B.n413 585
R284 B.n412 B.n411 585
R285 B.n410 B.n409 585
R286 B.n408 B.n407 585
R287 B.n406 B.n405 585
R288 B.n404 B.n403 585
R289 B.n402 B.n401 585
R290 B.n400 B.n399 585
R291 B.n398 B.n397 585
R292 B.n396 B.n395 585
R293 B.n394 B.n393 585
R294 B.n392 B.n391 585
R295 B.n390 B.n389 585
R296 B.n388 B.n387 585
R297 B.n386 B.n385 585
R298 B.n384 B.n383 585
R299 B.n382 B.n381 585
R300 B.n380 B.n379 585
R301 B.n378 B.n377 585
R302 B.n376 B.n375 585
R303 B.n374 B.n373 585
R304 B.n372 B.n371 585
R305 B.n370 B.n369 585
R306 B.n368 B.n367 585
R307 B.n366 B.n365 585
R308 B.n364 B.n363 585
R309 B.n316 B.n315 585
R310 B.n520 B.n519 585
R311 B.n519 B.n518 585
R312 B.n312 B.n311 585
R313 B.n313 B.n312 585
R314 B.n526 B.n525 585
R315 B.n525 B.n524 585
R316 B.n527 B.n310 585
R317 B.n310 B.n309 585
R318 B.n529 B.n528 585
R319 B.n530 B.n529 585
R320 B.n304 B.n303 585
R321 B.n305 B.n304 585
R322 B.n539 B.n538 585
R323 B.n538 B.n537 585
R324 B.n540 B.n302 585
R325 B.n536 B.n302 585
R326 B.n542 B.n541 585
R327 B.n543 B.n542 585
R328 B.n297 B.n296 585
R329 B.n298 B.n297 585
R330 B.n551 B.n550 585
R331 B.n550 B.n549 585
R332 B.n552 B.n295 585
R333 B.n295 B.n294 585
R334 B.n554 B.n553 585
R335 B.n555 B.n554 585
R336 B.n289 B.n288 585
R337 B.n290 B.n289 585
R338 B.n563 B.n562 585
R339 B.n562 B.n561 585
R340 B.n564 B.n287 585
R341 B.n287 B.n286 585
R342 B.n566 B.n565 585
R343 B.n567 B.n566 585
R344 B.n281 B.n280 585
R345 B.n282 B.n281 585
R346 B.n575 B.n574 585
R347 B.n574 B.n573 585
R348 B.n576 B.n279 585
R349 B.n279 B.n278 585
R350 B.n578 B.n577 585
R351 B.n579 B.n578 585
R352 B.n273 B.n272 585
R353 B.n274 B.n273 585
R354 B.n587 B.n586 585
R355 B.n586 B.n585 585
R356 B.n588 B.n271 585
R357 B.n271 B.n269 585
R358 B.n590 B.n589 585
R359 B.n591 B.n590 585
R360 B.n265 B.n264 585
R361 B.n270 B.n265 585
R362 B.n600 B.n599 585
R363 B.n599 B.n598 585
R364 B.n601 B.n263 585
R365 B.n263 B.n262 585
R366 B.n603 B.n602 585
R367 B.n604 B.n603 585
R368 B.n3 B.n0 585
R369 B.n4 B.n3 585
R370 B.n706 B.n1 585
R371 B.n707 B.n706 585
R372 B.n705 B.n704 585
R373 B.n705 B.n8 585
R374 B.n703 B.n9 585
R375 B.n12 B.n9 585
R376 B.n702 B.n701 585
R377 B.n701 B.n700 585
R378 B.n11 B.n10 585
R379 B.n699 B.n11 585
R380 B.n697 B.n696 585
R381 B.n698 B.n697 585
R382 B.n695 B.n17 585
R383 B.n17 B.n16 585
R384 B.n694 B.n693 585
R385 B.n693 B.n692 585
R386 B.n19 B.n18 585
R387 B.n691 B.n19 585
R388 B.n689 B.n688 585
R389 B.n690 B.n689 585
R390 B.n687 B.n24 585
R391 B.n24 B.n23 585
R392 B.n686 B.n685 585
R393 B.n685 B.n684 585
R394 B.n26 B.n25 585
R395 B.n683 B.n26 585
R396 B.n681 B.n680 585
R397 B.n682 B.n681 585
R398 B.n679 B.n31 585
R399 B.n31 B.n30 585
R400 B.n678 B.n677 585
R401 B.n677 B.n676 585
R402 B.n33 B.n32 585
R403 B.n675 B.n33 585
R404 B.n673 B.n672 585
R405 B.n674 B.n673 585
R406 B.n671 B.n38 585
R407 B.n38 B.n37 585
R408 B.n670 B.n669 585
R409 B.n669 B.n668 585
R410 B.n40 B.n39 585
R411 B.n667 B.n40 585
R412 B.n665 B.n664 585
R413 B.n666 B.n665 585
R414 B.n663 B.n44 585
R415 B.n47 B.n44 585
R416 B.n662 B.n661 585
R417 B.n661 B.n660 585
R418 B.n46 B.n45 585
R419 B.n659 B.n46 585
R420 B.n657 B.n656 585
R421 B.n658 B.n657 585
R422 B.n655 B.n52 585
R423 B.n52 B.n51 585
R424 B.n654 B.n653 585
R425 B.n653 B.n652 585
R426 B.n54 B.n53 585
R427 B.n651 B.n54 585
R428 B.n710 B.n709 585
R429 B.n708 B.n2 585
R430 B.n101 B.n54 492.5
R431 B.n648 B.n56 492.5
R432 B.n519 B.n314 492.5
R433 B.n516 B.n312 492.5
R434 B.n99 B.t11 319.495
R435 B.n97 B.t15 319.495
R436 B.n360 B.t4 319.495
R437 B.n357 B.t8 319.495
R438 B.n650 B.n649 256.663
R439 B.n650 B.n95 256.663
R440 B.n650 B.n94 256.663
R441 B.n650 B.n93 256.663
R442 B.n650 B.n92 256.663
R443 B.n650 B.n91 256.663
R444 B.n650 B.n90 256.663
R445 B.n650 B.n89 256.663
R446 B.n650 B.n88 256.663
R447 B.n650 B.n87 256.663
R448 B.n650 B.n86 256.663
R449 B.n650 B.n85 256.663
R450 B.n650 B.n84 256.663
R451 B.n650 B.n83 256.663
R452 B.n650 B.n82 256.663
R453 B.n650 B.n81 256.663
R454 B.n650 B.n80 256.663
R455 B.n650 B.n79 256.663
R456 B.n650 B.n78 256.663
R457 B.n650 B.n77 256.663
R458 B.n650 B.n76 256.663
R459 B.n650 B.n75 256.663
R460 B.n650 B.n74 256.663
R461 B.n650 B.n73 256.663
R462 B.n650 B.n72 256.663
R463 B.n650 B.n71 256.663
R464 B.n650 B.n70 256.663
R465 B.n650 B.n69 256.663
R466 B.n650 B.n68 256.663
R467 B.n650 B.n67 256.663
R468 B.n650 B.n66 256.663
R469 B.n650 B.n65 256.663
R470 B.n650 B.n64 256.663
R471 B.n650 B.n63 256.663
R472 B.n650 B.n62 256.663
R473 B.n650 B.n61 256.663
R474 B.n650 B.n60 256.663
R475 B.n650 B.n59 256.663
R476 B.n650 B.n58 256.663
R477 B.n650 B.n57 256.663
R478 B.n518 B.n517 256.663
R479 B.n518 B.n317 256.663
R480 B.n518 B.n318 256.663
R481 B.n518 B.n319 256.663
R482 B.n518 B.n320 256.663
R483 B.n518 B.n321 256.663
R484 B.n518 B.n322 256.663
R485 B.n518 B.n323 256.663
R486 B.n518 B.n324 256.663
R487 B.n518 B.n325 256.663
R488 B.n518 B.n326 256.663
R489 B.n518 B.n327 256.663
R490 B.n518 B.n328 256.663
R491 B.n518 B.n329 256.663
R492 B.n518 B.n330 256.663
R493 B.n518 B.n331 256.663
R494 B.n518 B.n332 256.663
R495 B.n518 B.n333 256.663
R496 B.n518 B.n334 256.663
R497 B.n518 B.n335 256.663
R498 B.n518 B.n336 256.663
R499 B.n518 B.n337 256.663
R500 B.n518 B.n338 256.663
R501 B.n518 B.n339 256.663
R502 B.n518 B.n340 256.663
R503 B.n518 B.n341 256.663
R504 B.n518 B.n342 256.663
R505 B.n518 B.n343 256.663
R506 B.n518 B.n344 256.663
R507 B.n518 B.n345 256.663
R508 B.n518 B.n346 256.663
R509 B.n518 B.n347 256.663
R510 B.n518 B.n348 256.663
R511 B.n518 B.n349 256.663
R512 B.n518 B.n350 256.663
R513 B.n518 B.n351 256.663
R514 B.n518 B.n352 256.663
R515 B.n518 B.n353 256.663
R516 B.n518 B.n354 256.663
R517 B.n712 B.n711 256.663
R518 B.n105 B.n104 163.367
R519 B.n109 B.n108 163.367
R520 B.n113 B.n112 163.367
R521 B.n117 B.n116 163.367
R522 B.n121 B.n120 163.367
R523 B.n125 B.n124 163.367
R524 B.n129 B.n128 163.367
R525 B.n133 B.n132 163.367
R526 B.n137 B.n136 163.367
R527 B.n141 B.n140 163.367
R528 B.n145 B.n144 163.367
R529 B.n149 B.n148 163.367
R530 B.n153 B.n152 163.367
R531 B.n157 B.n156 163.367
R532 B.n161 B.n160 163.367
R533 B.n165 B.n164 163.367
R534 B.n169 B.n168 163.367
R535 B.n174 B.n173 163.367
R536 B.n178 B.n177 163.367
R537 B.n182 B.n181 163.367
R538 B.n186 B.n185 163.367
R539 B.n190 B.n189 163.367
R540 B.n195 B.n194 163.367
R541 B.n199 B.n198 163.367
R542 B.n203 B.n202 163.367
R543 B.n207 B.n206 163.367
R544 B.n211 B.n210 163.367
R545 B.n215 B.n214 163.367
R546 B.n219 B.n218 163.367
R547 B.n223 B.n222 163.367
R548 B.n227 B.n226 163.367
R549 B.n231 B.n230 163.367
R550 B.n235 B.n234 163.367
R551 B.n239 B.n238 163.367
R552 B.n243 B.n242 163.367
R553 B.n247 B.n246 163.367
R554 B.n251 B.n250 163.367
R555 B.n255 B.n254 163.367
R556 B.n257 B.n96 163.367
R557 B.n523 B.n314 163.367
R558 B.n523 B.n308 163.367
R559 B.n531 B.n308 163.367
R560 B.n531 B.n306 163.367
R561 B.n535 B.n306 163.367
R562 B.n535 B.n301 163.367
R563 B.n544 B.n301 163.367
R564 B.n544 B.n299 163.367
R565 B.n548 B.n299 163.367
R566 B.n548 B.n293 163.367
R567 B.n556 B.n293 163.367
R568 B.n556 B.n291 163.367
R569 B.n560 B.n291 163.367
R570 B.n560 B.n285 163.367
R571 B.n568 B.n285 163.367
R572 B.n568 B.n283 163.367
R573 B.n572 B.n283 163.367
R574 B.n572 B.n277 163.367
R575 B.n580 B.n277 163.367
R576 B.n580 B.n275 163.367
R577 B.n584 B.n275 163.367
R578 B.n584 B.n268 163.367
R579 B.n592 B.n268 163.367
R580 B.n592 B.n266 163.367
R581 B.n597 B.n266 163.367
R582 B.n597 B.n261 163.367
R583 B.n605 B.n261 163.367
R584 B.n606 B.n605 163.367
R585 B.n606 B.n5 163.367
R586 B.n6 B.n5 163.367
R587 B.n7 B.n6 163.367
R588 B.n612 B.n7 163.367
R589 B.n613 B.n612 163.367
R590 B.n613 B.n13 163.367
R591 B.n14 B.n13 163.367
R592 B.n15 B.n14 163.367
R593 B.n618 B.n15 163.367
R594 B.n618 B.n20 163.367
R595 B.n21 B.n20 163.367
R596 B.n22 B.n21 163.367
R597 B.n623 B.n22 163.367
R598 B.n623 B.n27 163.367
R599 B.n28 B.n27 163.367
R600 B.n29 B.n28 163.367
R601 B.n628 B.n29 163.367
R602 B.n628 B.n34 163.367
R603 B.n35 B.n34 163.367
R604 B.n36 B.n35 163.367
R605 B.n633 B.n36 163.367
R606 B.n633 B.n41 163.367
R607 B.n42 B.n41 163.367
R608 B.n43 B.n42 163.367
R609 B.n638 B.n43 163.367
R610 B.n638 B.n48 163.367
R611 B.n49 B.n48 163.367
R612 B.n50 B.n49 163.367
R613 B.n643 B.n50 163.367
R614 B.n643 B.n55 163.367
R615 B.n56 B.n55 163.367
R616 B.n356 B.n355 163.367
R617 B.n511 B.n355 163.367
R618 B.n509 B.n508 163.367
R619 B.n505 B.n504 163.367
R620 B.n501 B.n500 163.367
R621 B.n497 B.n496 163.367
R622 B.n493 B.n492 163.367
R623 B.n489 B.n488 163.367
R624 B.n485 B.n484 163.367
R625 B.n481 B.n480 163.367
R626 B.n477 B.n476 163.367
R627 B.n473 B.n472 163.367
R628 B.n469 B.n468 163.367
R629 B.n465 B.n464 163.367
R630 B.n461 B.n460 163.367
R631 B.n457 B.n456 163.367
R632 B.n453 B.n452 163.367
R633 B.n449 B.n448 163.367
R634 B.n445 B.n444 163.367
R635 B.n441 B.n440 163.367
R636 B.n437 B.n436 163.367
R637 B.n433 B.n432 163.367
R638 B.n429 B.n428 163.367
R639 B.n425 B.n424 163.367
R640 B.n421 B.n420 163.367
R641 B.n417 B.n416 163.367
R642 B.n413 B.n412 163.367
R643 B.n409 B.n408 163.367
R644 B.n405 B.n404 163.367
R645 B.n401 B.n400 163.367
R646 B.n397 B.n396 163.367
R647 B.n393 B.n392 163.367
R648 B.n389 B.n388 163.367
R649 B.n385 B.n384 163.367
R650 B.n381 B.n380 163.367
R651 B.n377 B.n376 163.367
R652 B.n373 B.n372 163.367
R653 B.n369 B.n368 163.367
R654 B.n365 B.n364 163.367
R655 B.n519 B.n316 163.367
R656 B.n525 B.n312 163.367
R657 B.n525 B.n310 163.367
R658 B.n529 B.n310 163.367
R659 B.n529 B.n304 163.367
R660 B.n538 B.n304 163.367
R661 B.n538 B.n302 163.367
R662 B.n542 B.n302 163.367
R663 B.n542 B.n297 163.367
R664 B.n550 B.n297 163.367
R665 B.n550 B.n295 163.367
R666 B.n554 B.n295 163.367
R667 B.n554 B.n289 163.367
R668 B.n562 B.n289 163.367
R669 B.n562 B.n287 163.367
R670 B.n566 B.n287 163.367
R671 B.n566 B.n281 163.367
R672 B.n574 B.n281 163.367
R673 B.n574 B.n279 163.367
R674 B.n578 B.n279 163.367
R675 B.n578 B.n273 163.367
R676 B.n586 B.n273 163.367
R677 B.n586 B.n271 163.367
R678 B.n590 B.n271 163.367
R679 B.n590 B.n265 163.367
R680 B.n599 B.n265 163.367
R681 B.n599 B.n263 163.367
R682 B.n603 B.n263 163.367
R683 B.n603 B.n3 163.367
R684 B.n710 B.n3 163.367
R685 B.n706 B.n2 163.367
R686 B.n706 B.n705 163.367
R687 B.n705 B.n9 163.367
R688 B.n701 B.n9 163.367
R689 B.n701 B.n11 163.367
R690 B.n697 B.n11 163.367
R691 B.n697 B.n17 163.367
R692 B.n693 B.n17 163.367
R693 B.n693 B.n19 163.367
R694 B.n689 B.n19 163.367
R695 B.n689 B.n24 163.367
R696 B.n685 B.n24 163.367
R697 B.n685 B.n26 163.367
R698 B.n681 B.n26 163.367
R699 B.n681 B.n31 163.367
R700 B.n677 B.n31 163.367
R701 B.n677 B.n33 163.367
R702 B.n673 B.n33 163.367
R703 B.n673 B.n38 163.367
R704 B.n669 B.n38 163.367
R705 B.n669 B.n40 163.367
R706 B.n665 B.n40 163.367
R707 B.n665 B.n44 163.367
R708 B.n661 B.n44 163.367
R709 B.n661 B.n46 163.367
R710 B.n657 B.n46 163.367
R711 B.n657 B.n52 163.367
R712 B.n653 B.n52 163.367
R713 B.n653 B.n54 163.367
R714 B.n97 B.t16 120.522
R715 B.n360 B.t7 120.522
R716 B.n99 B.t13 120.51
R717 B.n357 B.t10 120.51
R718 B.n518 B.n313 92.732
R719 B.n651 B.n650 92.732
R720 B.n98 B.t17 73.3953
R721 B.n361 B.t6 73.3953
R722 B.n100 B.t14 73.3836
R723 B.n358 B.t9 73.3836
R724 B.n101 B.n57 71.676
R725 B.n105 B.n58 71.676
R726 B.n109 B.n59 71.676
R727 B.n113 B.n60 71.676
R728 B.n117 B.n61 71.676
R729 B.n121 B.n62 71.676
R730 B.n125 B.n63 71.676
R731 B.n129 B.n64 71.676
R732 B.n133 B.n65 71.676
R733 B.n137 B.n66 71.676
R734 B.n141 B.n67 71.676
R735 B.n145 B.n68 71.676
R736 B.n149 B.n69 71.676
R737 B.n153 B.n70 71.676
R738 B.n157 B.n71 71.676
R739 B.n161 B.n72 71.676
R740 B.n165 B.n73 71.676
R741 B.n169 B.n74 71.676
R742 B.n174 B.n75 71.676
R743 B.n178 B.n76 71.676
R744 B.n182 B.n77 71.676
R745 B.n186 B.n78 71.676
R746 B.n190 B.n79 71.676
R747 B.n195 B.n80 71.676
R748 B.n199 B.n81 71.676
R749 B.n203 B.n82 71.676
R750 B.n207 B.n83 71.676
R751 B.n211 B.n84 71.676
R752 B.n215 B.n85 71.676
R753 B.n219 B.n86 71.676
R754 B.n223 B.n87 71.676
R755 B.n227 B.n88 71.676
R756 B.n231 B.n89 71.676
R757 B.n235 B.n90 71.676
R758 B.n239 B.n91 71.676
R759 B.n243 B.n92 71.676
R760 B.n247 B.n93 71.676
R761 B.n251 B.n94 71.676
R762 B.n255 B.n95 71.676
R763 B.n649 B.n96 71.676
R764 B.n649 B.n648 71.676
R765 B.n257 B.n95 71.676
R766 B.n254 B.n94 71.676
R767 B.n250 B.n93 71.676
R768 B.n246 B.n92 71.676
R769 B.n242 B.n91 71.676
R770 B.n238 B.n90 71.676
R771 B.n234 B.n89 71.676
R772 B.n230 B.n88 71.676
R773 B.n226 B.n87 71.676
R774 B.n222 B.n86 71.676
R775 B.n218 B.n85 71.676
R776 B.n214 B.n84 71.676
R777 B.n210 B.n83 71.676
R778 B.n206 B.n82 71.676
R779 B.n202 B.n81 71.676
R780 B.n198 B.n80 71.676
R781 B.n194 B.n79 71.676
R782 B.n189 B.n78 71.676
R783 B.n185 B.n77 71.676
R784 B.n181 B.n76 71.676
R785 B.n177 B.n75 71.676
R786 B.n173 B.n74 71.676
R787 B.n168 B.n73 71.676
R788 B.n164 B.n72 71.676
R789 B.n160 B.n71 71.676
R790 B.n156 B.n70 71.676
R791 B.n152 B.n69 71.676
R792 B.n148 B.n68 71.676
R793 B.n144 B.n67 71.676
R794 B.n140 B.n66 71.676
R795 B.n136 B.n65 71.676
R796 B.n132 B.n64 71.676
R797 B.n128 B.n63 71.676
R798 B.n124 B.n62 71.676
R799 B.n120 B.n61 71.676
R800 B.n116 B.n60 71.676
R801 B.n112 B.n59 71.676
R802 B.n108 B.n58 71.676
R803 B.n104 B.n57 71.676
R804 B.n517 B.n516 71.676
R805 B.n511 B.n317 71.676
R806 B.n508 B.n318 71.676
R807 B.n504 B.n319 71.676
R808 B.n500 B.n320 71.676
R809 B.n496 B.n321 71.676
R810 B.n492 B.n322 71.676
R811 B.n488 B.n323 71.676
R812 B.n484 B.n324 71.676
R813 B.n480 B.n325 71.676
R814 B.n476 B.n326 71.676
R815 B.n472 B.n327 71.676
R816 B.n468 B.n328 71.676
R817 B.n464 B.n329 71.676
R818 B.n460 B.n330 71.676
R819 B.n456 B.n331 71.676
R820 B.n452 B.n332 71.676
R821 B.n448 B.n333 71.676
R822 B.n444 B.n334 71.676
R823 B.n440 B.n335 71.676
R824 B.n436 B.n336 71.676
R825 B.n432 B.n337 71.676
R826 B.n428 B.n338 71.676
R827 B.n424 B.n339 71.676
R828 B.n420 B.n340 71.676
R829 B.n416 B.n341 71.676
R830 B.n412 B.n342 71.676
R831 B.n408 B.n343 71.676
R832 B.n404 B.n344 71.676
R833 B.n400 B.n345 71.676
R834 B.n396 B.n346 71.676
R835 B.n392 B.n347 71.676
R836 B.n388 B.n348 71.676
R837 B.n384 B.n349 71.676
R838 B.n380 B.n350 71.676
R839 B.n376 B.n351 71.676
R840 B.n372 B.n352 71.676
R841 B.n368 B.n353 71.676
R842 B.n364 B.n354 71.676
R843 B.n517 B.n356 71.676
R844 B.n509 B.n317 71.676
R845 B.n505 B.n318 71.676
R846 B.n501 B.n319 71.676
R847 B.n497 B.n320 71.676
R848 B.n493 B.n321 71.676
R849 B.n489 B.n322 71.676
R850 B.n485 B.n323 71.676
R851 B.n481 B.n324 71.676
R852 B.n477 B.n325 71.676
R853 B.n473 B.n326 71.676
R854 B.n469 B.n327 71.676
R855 B.n465 B.n328 71.676
R856 B.n461 B.n329 71.676
R857 B.n457 B.n330 71.676
R858 B.n453 B.n331 71.676
R859 B.n449 B.n332 71.676
R860 B.n445 B.n333 71.676
R861 B.n441 B.n334 71.676
R862 B.n437 B.n335 71.676
R863 B.n433 B.n336 71.676
R864 B.n429 B.n337 71.676
R865 B.n425 B.n338 71.676
R866 B.n421 B.n339 71.676
R867 B.n417 B.n340 71.676
R868 B.n413 B.n341 71.676
R869 B.n409 B.n342 71.676
R870 B.n405 B.n343 71.676
R871 B.n401 B.n344 71.676
R872 B.n397 B.n345 71.676
R873 B.n393 B.n346 71.676
R874 B.n389 B.n347 71.676
R875 B.n385 B.n348 71.676
R876 B.n381 B.n349 71.676
R877 B.n377 B.n350 71.676
R878 B.n373 B.n351 71.676
R879 B.n369 B.n352 71.676
R880 B.n365 B.n353 71.676
R881 B.n354 B.n316 71.676
R882 B.n711 B.n710 71.676
R883 B.n711 B.n2 71.676
R884 B.n171 B.n100 59.5399
R885 B.n192 B.n98 59.5399
R886 B.n362 B.n361 59.5399
R887 B.n359 B.n358 59.5399
R888 B.n524 B.n313 49.652
R889 B.n524 B.n309 49.652
R890 B.n530 B.n309 49.652
R891 B.n530 B.n305 49.652
R892 B.n537 B.n305 49.652
R893 B.n537 B.n536 49.652
R894 B.n543 B.n298 49.652
R895 B.n549 B.n298 49.652
R896 B.n549 B.n294 49.652
R897 B.n555 B.n294 49.652
R898 B.n555 B.n290 49.652
R899 B.n561 B.n290 49.652
R900 B.n561 B.n286 49.652
R901 B.n567 B.n286 49.652
R902 B.n567 B.n282 49.652
R903 B.n573 B.n282 49.652
R904 B.n579 B.n278 49.652
R905 B.n579 B.n274 49.652
R906 B.n585 B.n274 49.652
R907 B.n585 B.n269 49.652
R908 B.n591 B.n269 49.652
R909 B.n591 B.n270 49.652
R910 B.n598 B.n262 49.652
R911 B.n604 B.n262 49.652
R912 B.n604 B.n4 49.652
R913 B.n709 B.n4 49.652
R914 B.n709 B.n708 49.652
R915 B.n708 B.n707 49.652
R916 B.n707 B.n8 49.652
R917 B.n12 B.n8 49.652
R918 B.n700 B.n12 49.652
R919 B.n699 B.n698 49.652
R920 B.n698 B.n16 49.652
R921 B.n692 B.n16 49.652
R922 B.n692 B.n691 49.652
R923 B.n691 B.n690 49.652
R924 B.n690 B.n23 49.652
R925 B.n684 B.n683 49.652
R926 B.n683 B.n682 49.652
R927 B.n682 B.n30 49.652
R928 B.n676 B.n30 49.652
R929 B.n676 B.n675 49.652
R930 B.n675 B.n674 49.652
R931 B.n674 B.n37 49.652
R932 B.n668 B.n37 49.652
R933 B.n668 B.n667 49.652
R934 B.n667 B.n666 49.652
R935 B.n660 B.n47 49.652
R936 B.n660 B.n659 49.652
R937 B.n659 B.n658 49.652
R938 B.n658 B.n51 49.652
R939 B.n652 B.n51 49.652
R940 B.n652 B.n651 49.652
R941 B.n100 B.n99 47.1278
R942 B.n98 B.n97 47.1278
R943 B.n361 B.n360 47.1278
R944 B.n358 B.n357 47.1278
R945 B.n536 B.t5 40.89
R946 B.t1 B.n278 40.89
R947 B.t2 B.n23 40.89
R948 B.n47 B.t12 40.89
R949 B.n598 B.t0 33.5883
R950 B.n700 B.t3 33.5883
R951 B.n515 B.n311 32.0005
R952 B.n521 B.n520 32.0005
R953 B.n647 B.n646 32.0005
R954 B.n102 B.n53 32.0005
R955 B B.n712 18.0485
R956 B.n270 B.t0 16.0642
R957 B.t3 B.n699 16.0642
R958 B.n526 B.n311 10.6151
R959 B.n527 B.n526 10.6151
R960 B.n528 B.n527 10.6151
R961 B.n528 B.n303 10.6151
R962 B.n539 B.n303 10.6151
R963 B.n540 B.n539 10.6151
R964 B.n541 B.n540 10.6151
R965 B.n541 B.n296 10.6151
R966 B.n551 B.n296 10.6151
R967 B.n552 B.n551 10.6151
R968 B.n553 B.n552 10.6151
R969 B.n553 B.n288 10.6151
R970 B.n563 B.n288 10.6151
R971 B.n564 B.n563 10.6151
R972 B.n565 B.n564 10.6151
R973 B.n565 B.n280 10.6151
R974 B.n575 B.n280 10.6151
R975 B.n576 B.n575 10.6151
R976 B.n577 B.n576 10.6151
R977 B.n577 B.n272 10.6151
R978 B.n587 B.n272 10.6151
R979 B.n588 B.n587 10.6151
R980 B.n589 B.n588 10.6151
R981 B.n589 B.n264 10.6151
R982 B.n600 B.n264 10.6151
R983 B.n601 B.n600 10.6151
R984 B.n602 B.n601 10.6151
R985 B.n602 B.n0 10.6151
R986 B.n515 B.n514 10.6151
R987 B.n514 B.n513 10.6151
R988 B.n513 B.n512 10.6151
R989 B.n512 B.n510 10.6151
R990 B.n510 B.n507 10.6151
R991 B.n507 B.n506 10.6151
R992 B.n506 B.n503 10.6151
R993 B.n503 B.n502 10.6151
R994 B.n502 B.n499 10.6151
R995 B.n499 B.n498 10.6151
R996 B.n498 B.n495 10.6151
R997 B.n495 B.n494 10.6151
R998 B.n494 B.n491 10.6151
R999 B.n491 B.n490 10.6151
R1000 B.n490 B.n487 10.6151
R1001 B.n487 B.n486 10.6151
R1002 B.n486 B.n483 10.6151
R1003 B.n483 B.n482 10.6151
R1004 B.n482 B.n479 10.6151
R1005 B.n479 B.n478 10.6151
R1006 B.n478 B.n475 10.6151
R1007 B.n475 B.n474 10.6151
R1008 B.n474 B.n471 10.6151
R1009 B.n471 B.n470 10.6151
R1010 B.n470 B.n467 10.6151
R1011 B.n467 B.n466 10.6151
R1012 B.n466 B.n463 10.6151
R1013 B.n463 B.n462 10.6151
R1014 B.n462 B.n459 10.6151
R1015 B.n459 B.n458 10.6151
R1016 B.n458 B.n455 10.6151
R1017 B.n455 B.n454 10.6151
R1018 B.n454 B.n451 10.6151
R1019 B.n451 B.n450 10.6151
R1020 B.n447 B.n446 10.6151
R1021 B.n446 B.n443 10.6151
R1022 B.n443 B.n442 10.6151
R1023 B.n442 B.n439 10.6151
R1024 B.n439 B.n438 10.6151
R1025 B.n438 B.n435 10.6151
R1026 B.n435 B.n434 10.6151
R1027 B.n434 B.n431 10.6151
R1028 B.n431 B.n430 10.6151
R1029 B.n427 B.n426 10.6151
R1030 B.n426 B.n423 10.6151
R1031 B.n423 B.n422 10.6151
R1032 B.n422 B.n419 10.6151
R1033 B.n419 B.n418 10.6151
R1034 B.n418 B.n415 10.6151
R1035 B.n415 B.n414 10.6151
R1036 B.n414 B.n411 10.6151
R1037 B.n411 B.n410 10.6151
R1038 B.n410 B.n407 10.6151
R1039 B.n407 B.n406 10.6151
R1040 B.n406 B.n403 10.6151
R1041 B.n403 B.n402 10.6151
R1042 B.n402 B.n399 10.6151
R1043 B.n399 B.n398 10.6151
R1044 B.n398 B.n395 10.6151
R1045 B.n395 B.n394 10.6151
R1046 B.n394 B.n391 10.6151
R1047 B.n391 B.n390 10.6151
R1048 B.n390 B.n387 10.6151
R1049 B.n387 B.n386 10.6151
R1050 B.n386 B.n383 10.6151
R1051 B.n383 B.n382 10.6151
R1052 B.n382 B.n379 10.6151
R1053 B.n379 B.n378 10.6151
R1054 B.n378 B.n375 10.6151
R1055 B.n375 B.n374 10.6151
R1056 B.n374 B.n371 10.6151
R1057 B.n371 B.n370 10.6151
R1058 B.n370 B.n367 10.6151
R1059 B.n367 B.n366 10.6151
R1060 B.n366 B.n363 10.6151
R1061 B.n363 B.n315 10.6151
R1062 B.n520 B.n315 10.6151
R1063 B.n522 B.n521 10.6151
R1064 B.n522 B.n307 10.6151
R1065 B.n532 B.n307 10.6151
R1066 B.n533 B.n532 10.6151
R1067 B.n534 B.n533 10.6151
R1068 B.n534 B.n300 10.6151
R1069 B.n545 B.n300 10.6151
R1070 B.n546 B.n545 10.6151
R1071 B.n547 B.n546 10.6151
R1072 B.n547 B.n292 10.6151
R1073 B.n557 B.n292 10.6151
R1074 B.n558 B.n557 10.6151
R1075 B.n559 B.n558 10.6151
R1076 B.n559 B.n284 10.6151
R1077 B.n569 B.n284 10.6151
R1078 B.n570 B.n569 10.6151
R1079 B.n571 B.n570 10.6151
R1080 B.n571 B.n276 10.6151
R1081 B.n581 B.n276 10.6151
R1082 B.n582 B.n581 10.6151
R1083 B.n583 B.n582 10.6151
R1084 B.n583 B.n267 10.6151
R1085 B.n593 B.n267 10.6151
R1086 B.n594 B.n593 10.6151
R1087 B.n596 B.n594 10.6151
R1088 B.n596 B.n595 10.6151
R1089 B.n595 B.n260 10.6151
R1090 B.n607 B.n260 10.6151
R1091 B.n608 B.n607 10.6151
R1092 B.n609 B.n608 10.6151
R1093 B.n610 B.n609 10.6151
R1094 B.n611 B.n610 10.6151
R1095 B.n614 B.n611 10.6151
R1096 B.n615 B.n614 10.6151
R1097 B.n616 B.n615 10.6151
R1098 B.n617 B.n616 10.6151
R1099 B.n619 B.n617 10.6151
R1100 B.n620 B.n619 10.6151
R1101 B.n621 B.n620 10.6151
R1102 B.n622 B.n621 10.6151
R1103 B.n624 B.n622 10.6151
R1104 B.n625 B.n624 10.6151
R1105 B.n626 B.n625 10.6151
R1106 B.n627 B.n626 10.6151
R1107 B.n629 B.n627 10.6151
R1108 B.n630 B.n629 10.6151
R1109 B.n631 B.n630 10.6151
R1110 B.n632 B.n631 10.6151
R1111 B.n634 B.n632 10.6151
R1112 B.n635 B.n634 10.6151
R1113 B.n636 B.n635 10.6151
R1114 B.n637 B.n636 10.6151
R1115 B.n639 B.n637 10.6151
R1116 B.n640 B.n639 10.6151
R1117 B.n641 B.n640 10.6151
R1118 B.n642 B.n641 10.6151
R1119 B.n644 B.n642 10.6151
R1120 B.n645 B.n644 10.6151
R1121 B.n646 B.n645 10.6151
R1122 B.n704 B.n1 10.6151
R1123 B.n704 B.n703 10.6151
R1124 B.n703 B.n702 10.6151
R1125 B.n702 B.n10 10.6151
R1126 B.n696 B.n10 10.6151
R1127 B.n696 B.n695 10.6151
R1128 B.n695 B.n694 10.6151
R1129 B.n694 B.n18 10.6151
R1130 B.n688 B.n18 10.6151
R1131 B.n688 B.n687 10.6151
R1132 B.n687 B.n686 10.6151
R1133 B.n686 B.n25 10.6151
R1134 B.n680 B.n25 10.6151
R1135 B.n680 B.n679 10.6151
R1136 B.n679 B.n678 10.6151
R1137 B.n678 B.n32 10.6151
R1138 B.n672 B.n32 10.6151
R1139 B.n672 B.n671 10.6151
R1140 B.n671 B.n670 10.6151
R1141 B.n670 B.n39 10.6151
R1142 B.n664 B.n39 10.6151
R1143 B.n664 B.n663 10.6151
R1144 B.n663 B.n662 10.6151
R1145 B.n662 B.n45 10.6151
R1146 B.n656 B.n45 10.6151
R1147 B.n656 B.n655 10.6151
R1148 B.n655 B.n654 10.6151
R1149 B.n654 B.n53 10.6151
R1150 B.n103 B.n102 10.6151
R1151 B.n106 B.n103 10.6151
R1152 B.n107 B.n106 10.6151
R1153 B.n110 B.n107 10.6151
R1154 B.n111 B.n110 10.6151
R1155 B.n114 B.n111 10.6151
R1156 B.n115 B.n114 10.6151
R1157 B.n118 B.n115 10.6151
R1158 B.n119 B.n118 10.6151
R1159 B.n122 B.n119 10.6151
R1160 B.n123 B.n122 10.6151
R1161 B.n126 B.n123 10.6151
R1162 B.n127 B.n126 10.6151
R1163 B.n130 B.n127 10.6151
R1164 B.n131 B.n130 10.6151
R1165 B.n134 B.n131 10.6151
R1166 B.n135 B.n134 10.6151
R1167 B.n138 B.n135 10.6151
R1168 B.n139 B.n138 10.6151
R1169 B.n142 B.n139 10.6151
R1170 B.n143 B.n142 10.6151
R1171 B.n146 B.n143 10.6151
R1172 B.n147 B.n146 10.6151
R1173 B.n150 B.n147 10.6151
R1174 B.n151 B.n150 10.6151
R1175 B.n154 B.n151 10.6151
R1176 B.n155 B.n154 10.6151
R1177 B.n158 B.n155 10.6151
R1178 B.n159 B.n158 10.6151
R1179 B.n162 B.n159 10.6151
R1180 B.n163 B.n162 10.6151
R1181 B.n166 B.n163 10.6151
R1182 B.n167 B.n166 10.6151
R1183 B.n170 B.n167 10.6151
R1184 B.n175 B.n172 10.6151
R1185 B.n176 B.n175 10.6151
R1186 B.n179 B.n176 10.6151
R1187 B.n180 B.n179 10.6151
R1188 B.n183 B.n180 10.6151
R1189 B.n184 B.n183 10.6151
R1190 B.n187 B.n184 10.6151
R1191 B.n188 B.n187 10.6151
R1192 B.n191 B.n188 10.6151
R1193 B.n196 B.n193 10.6151
R1194 B.n197 B.n196 10.6151
R1195 B.n200 B.n197 10.6151
R1196 B.n201 B.n200 10.6151
R1197 B.n204 B.n201 10.6151
R1198 B.n205 B.n204 10.6151
R1199 B.n208 B.n205 10.6151
R1200 B.n209 B.n208 10.6151
R1201 B.n212 B.n209 10.6151
R1202 B.n213 B.n212 10.6151
R1203 B.n216 B.n213 10.6151
R1204 B.n217 B.n216 10.6151
R1205 B.n220 B.n217 10.6151
R1206 B.n221 B.n220 10.6151
R1207 B.n224 B.n221 10.6151
R1208 B.n225 B.n224 10.6151
R1209 B.n228 B.n225 10.6151
R1210 B.n229 B.n228 10.6151
R1211 B.n232 B.n229 10.6151
R1212 B.n233 B.n232 10.6151
R1213 B.n236 B.n233 10.6151
R1214 B.n237 B.n236 10.6151
R1215 B.n240 B.n237 10.6151
R1216 B.n241 B.n240 10.6151
R1217 B.n244 B.n241 10.6151
R1218 B.n245 B.n244 10.6151
R1219 B.n248 B.n245 10.6151
R1220 B.n249 B.n248 10.6151
R1221 B.n252 B.n249 10.6151
R1222 B.n253 B.n252 10.6151
R1223 B.n256 B.n253 10.6151
R1224 B.n258 B.n256 10.6151
R1225 B.n259 B.n258 10.6151
R1226 B.n647 B.n259 10.6151
R1227 B.n450 B.n359 9.36635
R1228 B.n427 B.n362 9.36635
R1229 B.n171 B.n170 9.36635
R1230 B.n193 B.n192 9.36635
R1231 B.n543 B.t5 8.76253
R1232 B.n573 B.t1 8.76253
R1233 B.n684 B.t2 8.76253
R1234 B.n666 B.t12 8.76253
R1235 B.n712 B.n0 8.11757
R1236 B.n712 B.n1 8.11757
R1237 B.n447 B.n359 1.24928
R1238 B.n430 B.n362 1.24928
R1239 B.n172 B.n171 1.24928
R1240 B.n192 B.n191 1.24928
R1241 VP.n10 VP.n0 161.3
R1242 VP.n9 VP.n8 161.3
R1243 VP.n7 VP.n1 161.3
R1244 VP.n6 VP.n5 161.3
R1245 VP.n2 VP.t1 148.458
R1246 VP.n2 VP.t2 147.911
R1247 VP.n4 VP.t3 112.353
R1248 VP.n11 VP.t0 112.353
R1249 VP.n4 VP.n3 88.0021
R1250 VP.n12 VP.n11 88.0021
R1251 VP.n9 VP.n1 56.5193
R1252 VP.n3 VP.n2 50.047
R1253 VP.n5 VP.n1 24.4675
R1254 VP.n10 VP.n9 24.4675
R1255 VP.n5 VP.n4 22.7548
R1256 VP.n11 VP.n10 22.7548
R1257 VP.n6 VP.n3 0.278367
R1258 VP.n12 VP.n0 0.278367
R1259 VP.n7 VP.n6 0.189894
R1260 VP.n8 VP.n7 0.189894
R1261 VP.n8 VP.n0 0.189894
R1262 VP VP.n12 0.153454
R1263 VDD1 VDD1.n1 105.46
R1264 VDD1 VDD1.n0 66.555
R1265 VDD1.n0 VDD1.t2 2.02297
R1266 VDD1.n0 VDD1.t1 2.02297
R1267 VDD1.n1 VDD1.t0 2.02297
R1268 VDD1.n1 VDD1.t3 2.02297
C0 VTAIL VDD2 4.85212f
C1 VN VDD1 0.148675f
C2 VP VDD1 3.98158f
C3 VDD2 VDD1 0.908845f
C4 VP VN 5.41941f
C5 VTAIL VDD1 4.80126f
C6 VN VDD2 3.76825f
C7 VTAIL VN 3.70706f
C8 VP VDD2 0.362617f
C9 VTAIL VP 3.72117f
C10 VDD2 B 3.313436f
C11 VDD1 B 7.06638f
C12 VTAIL B 8.468587f
C13 VN B 9.5797f
C14 VP B 7.724688f
C15 VDD1.t2 B 0.209638f
C16 VDD1.t1 B 0.209638f
C17 VDD1.n0 B 1.84655f
C18 VDD1.t0 B 0.209638f
C19 VDD1.t3 B 0.209638f
C20 VDD1.n1 B 2.42135f
C21 VP.n0 B 0.039872f
C22 VP.t0 B 1.68315f
C23 VP.n1 B 0.044149f
C24 VP.t2 B 1.86965f
C25 VP.t1 B 1.87248f
C26 VP.n2 B 2.58712f
C27 VP.n3 B 1.56971f
C28 VP.t3 B 1.68315f
C29 VP.n4 B 0.711643f
C30 VP.n5 B 0.054416f
C31 VP.n6 B 0.039872f
C32 VP.n7 B 0.030243f
C33 VP.n8 B 0.030243f
C34 VP.n9 B 0.044149f
C35 VP.n10 B 0.054416f
C36 VP.n11 B 0.711643f
C37 VP.n12 B 0.034274f
C38 VTAIL.t7 B 1.40399f
C39 VTAIL.n0 B 0.293216f
C40 VTAIL.t0 B 1.40399f
C41 VTAIL.n1 B 0.346793f
C42 VTAIL.t1 B 1.40399f
C43 VTAIL.n2 B 1.12022f
C44 VTAIL.t4 B 1.404f
C45 VTAIL.n3 B 1.12021f
C46 VTAIL.t5 B 1.404f
C47 VTAIL.n4 B 0.346784f
C48 VTAIL.t3 B 1.404f
C49 VTAIL.n5 B 0.346784f
C50 VTAIL.t2 B 1.40399f
C51 VTAIL.n6 B 1.12022f
C52 VTAIL.t6 B 1.40399f
C53 VTAIL.n7 B 1.06034f
C54 VDD2.t3 B 0.209641f
C55 VDD2.t2 B 0.209641f
C56 VDD2.n0 B 2.39653f
C57 VDD2.t1 B 0.209641f
C58 VDD2.t0 B 0.209641f
C59 VDD2.n1 B 1.8462f
C60 VDD2.n2 B 3.42996f
C61 VN.t0 B 1.83793f
C62 VN.t1 B 1.83515f
C63 VN.n0 B 1.23431f
C64 VN.t2 B 1.83793f
C65 VN.t3 B 1.83515f
C66 VN.n1 B 2.55466f
.ends

