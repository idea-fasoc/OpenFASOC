* NGSPICE file created from diff_pair_sample_1225.ext - technology: sky130A

.subckt diff_pair_sample_1225 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X1 VTAIL.t14 VP.t1 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X2 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X3 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.14
X4 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.14
X5 VDD1.t0 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.14
X7 VTAIL.t12 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.14
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.14
X9 VDD1.t3 VP.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.14
X10 VTAIL.t6 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X11 VDD1.t7 VP.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.14
X12 VTAIL.t5 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.14
X13 VDD1.t5 VP.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X14 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X15 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.14
X16 VDD2.t1 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.14
X17 VTAIL.t8 VP.t7 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.14
X18 VDD2.t0 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.14
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.14
R0 VP.n15 VP.n12 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n18 VP.n11 161.3
R3 VP.n20 VP.n19 161.3
R4 VP.n22 VP.n10 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n9 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n28 VP.n8 161.3
R9 VP.n54 VP.n0 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n1 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n2 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n3 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n41 VP.n4 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n5 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n6 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n13 VP.t3 157.587
R24 VP.n7 VP.t7 123.091
R25 VP.n40 VP.t2 123.091
R26 VP.n47 VP.t0 123.091
R27 VP.n55 VP.t5 123.091
R28 VP.n29 VP.t4 123.091
R29 VP.n21 VP.t1 123.091
R30 VP.n14 VP.t6 123.091
R31 VP.n31 VP.n7 88.4915
R32 VP.n56 VP.n55 88.4915
R33 VP.n30 VP.n29 88.4915
R34 VP.n35 VP.n34 56.5193
R35 VP.n42 VP.n3 56.5193
R36 VP.n53 VP.n1 56.5193
R37 VP.n27 VP.n9 56.5193
R38 VP.n16 VP.n11 56.5193
R39 VP.n31 VP.n30 48.0299
R40 VP.n14 VP.n13 47.0153
R41 VP.n34 VP.n33 24.4675
R42 VP.n35 VP.n5 24.4675
R43 VP.n39 VP.n5 24.4675
R44 VP.n42 VP.n41 24.4675
R45 VP.n46 VP.n3 24.4675
R46 VP.n49 VP.n48 24.4675
R47 VP.n49 VP.n1 24.4675
R48 VP.n54 VP.n53 24.4675
R49 VP.n28 VP.n27 24.4675
R50 VP.n20 VP.n11 24.4675
R51 VP.n23 VP.n22 24.4675
R52 VP.n23 VP.n9 24.4675
R53 VP.n16 VP.n15 24.4675
R54 VP.n41 VP.n40 23.7335
R55 VP.n47 VP.n46 23.7335
R56 VP.n21 VP.n20 23.7335
R57 VP.n15 VP.n14 23.7335
R58 VP.n33 VP.n7 22.2655
R59 VP.n55 VP.n54 22.2655
R60 VP.n29 VP.n28 22.2655
R61 VP.n13 VP.n12 8.75906
R62 VP.n40 VP.n39 0.73451
R63 VP.n48 VP.n47 0.73451
R64 VP.n22 VP.n21 0.73451
R65 VP.n30 VP.n8 0.278367
R66 VP.n32 VP.n31 0.278367
R67 VP.n56 VP.n0 0.278367
R68 VP.n17 VP.n12 0.189894
R69 VP.n18 VP.n17 0.189894
R70 VP.n19 VP.n18 0.189894
R71 VP.n19 VP.n10 0.189894
R72 VP.n24 VP.n10 0.189894
R73 VP.n25 VP.n24 0.189894
R74 VP.n26 VP.n25 0.189894
R75 VP.n26 VP.n8 0.189894
R76 VP.n32 VP.n6 0.189894
R77 VP.n36 VP.n6 0.189894
R78 VP.n37 VP.n36 0.189894
R79 VP.n38 VP.n37 0.189894
R80 VP.n38 VP.n4 0.189894
R81 VP.n43 VP.n4 0.189894
R82 VP.n44 VP.n43 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n45 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VP VP.n56 0.153454
R90 VDD1 VDD1.n0 61.1987
R91 VDD1.n3 VDD1.n2 61.0849
R92 VDD1.n3 VDD1.n1 61.0849
R93 VDD1.n5 VDD1.n4 60.0756
R94 VDD1.n5 VDD1.n3 43.3026
R95 VDD1.n4 VDD1.t1 1.81203
R96 VDD1.n4 VDD1.t3 1.81203
R97 VDD1.n0 VDD1.t6 1.81203
R98 VDD1.n0 VDD1.t5 1.81203
R99 VDD1.n2 VDD1.t2 1.81203
R100 VDD1.n2 VDD1.t7 1.81203
R101 VDD1.n1 VDD1.t4 1.81203
R102 VDD1.n1 VDD1.t0 1.81203
R103 VDD1 VDD1.n5 1.00697
R104 VTAIL.n11 VTAIL.t12 45.2085
R105 VTAIL.n10 VTAIL.t3 45.2085
R106 VTAIL.n7 VTAIL.t7 45.2085
R107 VTAIL.n15 VTAIL.t4 45.2084
R108 VTAIL.n2 VTAIL.t5 45.2084
R109 VTAIL.n3 VTAIL.t10 45.2084
R110 VTAIL.n6 VTAIL.t8 45.2084
R111 VTAIL.n14 VTAIL.t11 45.2084
R112 VTAIL.n13 VTAIL.n12 43.397
R113 VTAIL.n9 VTAIL.n8 43.397
R114 VTAIL.n1 VTAIL.n0 43.3968
R115 VTAIL.n5 VTAIL.n4 43.3968
R116 VTAIL.n15 VTAIL.n14 23.9186
R117 VTAIL.n7 VTAIL.n6 23.9186
R118 VTAIL.n9 VTAIL.n7 2.12981
R119 VTAIL.n10 VTAIL.n9 2.12981
R120 VTAIL.n13 VTAIL.n11 2.12981
R121 VTAIL.n14 VTAIL.n13 2.12981
R122 VTAIL.n6 VTAIL.n5 2.12981
R123 VTAIL.n5 VTAIL.n3 2.12981
R124 VTAIL.n2 VTAIL.n1 2.12981
R125 VTAIL VTAIL.n15 2.07162
R126 VTAIL.n0 VTAIL.t1 1.81203
R127 VTAIL.n0 VTAIL.t6 1.81203
R128 VTAIL.n4 VTAIL.t13 1.81203
R129 VTAIL.n4 VTAIL.t15 1.81203
R130 VTAIL.n12 VTAIL.t9 1.81203
R131 VTAIL.n12 VTAIL.t14 1.81203
R132 VTAIL.n8 VTAIL.t0 1.81203
R133 VTAIL.n8 VTAIL.t2 1.81203
R134 VTAIL.n11 VTAIL.n10 0.470328
R135 VTAIL.n3 VTAIL.n2 0.470328
R136 VTAIL VTAIL.n1 0.0586897
R137 B.n801 B.n800 585
R138 B.n802 B.n801 585
R139 B.n302 B.n127 585
R140 B.n301 B.n300 585
R141 B.n299 B.n298 585
R142 B.n297 B.n296 585
R143 B.n295 B.n294 585
R144 B.n293 B.n292 585
R145 B.n291 B.n290 585
R146 B.n289 B.n288 585
R147 B.n287 B.n286 585
R148 B.n285 B.n284 585
R149 B.n283 B.n282 585
R150 B.n281 B.n280 585
R151 B.n279 B.n278 585
R152 B.n277 B.n276 585
R153 B.n275 B.n274 585
R154 B.n273 B.n272 585
R155 B.n271 B.n270 585
R156 B.n269 B.n268 585
R157 B.n267 B.n266 585
R158 B.n265 B.n264 585
R159 B.n263 B.n262 585
R160 B.n261 B.n260 585
R161 B.n259 B.n258 585
R162 B.n257 B.n256 585
R163 B.n255 B.n254 585
R164 B.n253 B.n252 585
R165 B.n251 B.n250 585
R166 B.n249 B.n248 585
R167 B.n247 B.n246 585
R168 B.n245 B.n244 585
R169 B.n243 B.n242 585
R170 B.n241 B.n240 585
R171 B.n239 B.n238 585
R172 B.n237 B.n236 585
R173 B.n235 B.n234 585
R174 B.n233 B.n232 585
R175 B.n231 B.n230 585
R176 B.n229 B.n228 585
R177 B.n227 B.n226 585
R178 B.n225 B.n224 585
R179 B.n223 B.n222 585
R180 B.n221 B.n220 585
R181 B.n219 B.n218 585
R182 B.n217 B.n216 585
R183 B.n215 B.n214 585
R184 B.n213 B.n212 585
R185 B.n211 B.n210 585
R186 B.n208 B.n207 585
R187 B.n206 B.n205 585
R188 B.n204 B.n203 585
R189 B.n202 B.n201 585
R190 B.n200 B.n199 585
R191 B.n198 B.n197 585
R192 B.n196 B.n195 585
R193 B.n194 B.n193 585
R194 B.n192 B.n191 585
R195 B.n190 B.n189 585
R196 B.n188 B.n187 585
R197 B.n186 B.n185 585
R198 B.n184 B.n183 585
R199 B.n182 B.n181 585
R200 B.n180 B.n179 585
R201 B.n178 B.n177 585
R202 B.n176 B.n175 585
R203 B.n174 B.n173 585
R204 B.n172 B.n171 585
R205 B.n170 B.n169 585
R206 B.n168 B.n167 585
R207 B.n166 B.n165 585
R208 B.n164 B.n163 585
R209 B.n162 B.n161 585
R210 B.n160 B.n159 585
R211 B.n158 B.n157 585
R212 B.n156 B.n155 585
R213 B.n154 B.n153 585
R214 B.n152 B.n151 585
R215 B.n150 B.n149 585
R216 B.n148 B.n147 585
R217 B.n146 B.n145 585
R218 B.n144 B.n143 585
R219 B.n142 B.n141 585
R220 B.n140 B.n139 585
R221 B.n138 B.n137 585
R222 B.n136 B.n135 585
R223 B.n134 B.n133 585
R224 B.n82 B.n81 585
R225 B.n799 B.n83 585
R226 B.n803 B.n83 585
R227 B.n798 B.n797 585
R228 B.n797 B.n79 585
R229 B.n796 B.n78 585
R230 B.n809 B.n78 585
R231 B.n795 B.n77 585
R232 B.n810 B.n77 585
R233 B.n794 B.n76 585
R234 B.n811 B.n76 585
R235 B.n793 B.n792 585
R236 B.n792 B.n72 585
R237 B.n791 B.n71 585
R238 B.n817 B.n71 585
R239 B.n790 B.n70 585
R240 B.t13 B.n70 585
R241 B.n789 B.n69 585
R242 B.n818 B.n69 585
R243 B.n788 B.n787 585
R244 B.n787 B.n65 585
R245 B.n786 B.n64 585
R246 B.n824 B.n64 585
R247 B.n785 B.n63 585
R248 B.n825 B.n63 585
R249 B.n784 B.n62 585
R250 B.n826 B.n62 585
R251 B.n783 B.n782 585
R252 B.n782 B.n58 585
R253 B.n781 B.n57 585
R254 B.n832 B.n57 585
R255 B.n780 B.n56 585
R256 B.n833 B.n56 585
R257 B.n779 B.n55 585
R258 B.n834 B.n55 585
R259 B.n778 B.n777 585
R260 B.n777 B.n54 585
R261 B.n776 B.n50 585
R262 B.n840 B.n50 585
R263 B.n775 B.n49 585
R264 B.n841 B.n49 585
R265 B.n774 B.n48 585
R266 B.n842 B.n48 585
R267 B.n773 B.n772 585
R268 B.n772 B.n44 585
R269 B.n771 B.n43 585
R270 B.n848 B.n43 585
R271 B.n770 B.n42 585
R272 B.n849 B.n42 585
R273 B.n769 B.n41 585
R274 B.n850 B.n41 585
R275 B.n768 B.n767 585
R276 B.n767 B.n37 585
R277 B.n766 B.n36 585
R278 B.n856 B.n36 585
R279 B.n765 B.n35 585
R280 B.n857 B.n35 585
R281 B.n764 B.n34 585
R282 B.n858 B.n34 585
R283 B.n763 B.n762 585
R284 B.n762 B.n30 585
R285 B.n761 B.n29 585
R286 B.n864 B.n29 585
R287 B.n760 B.n28 585
R288 B.n865 B.n28 585
R289 B.n759 B.n27 585
R290 B.t1 B.n27 585
R291 B.n758 B.n757 585
R292 B.n757 B.n23 585
R293 B.n756 B.n22 585
R294 B.n871 B.n22 585
R295 B.n755 B.n21 585
R296 B.n872 B.n21 585
R297 B.n754 B.n20 585
R298 B.n873 B.n20 585
R299 B.n753 B.n752 585
R300 B.n752 B.n16 585
R301 B.n751 B.n15 585
R302 B.n879 B.n15 585
R303 B.n750 B.n14 585
R304 B.n880 B.n14 585
R305 B.n749 B.n13 585
R306 B.n881 B.n13 585
R307 B.n748 B.n747 585
R308 B.n747 B.n12 585
R309 B.n746 B.n745 585
R310 B.n746 B.n8 585
R311 B.n744 B.n7 585
R312 B.n888 B.n7 585
R313 B.n743 B.n6 585
R314 B.n889 B.n6 585
R315 B.n742 B.n5 585
R316 B.n890 B.n5 585
R317 B.n741 B.n740 585
R318 B.n740 B.n4 585
R319 B.n739 B.n303 585
R320 B.n739 B.n738 585
R321 B.n729 B.n304 585
R322 B.n305 B.n304 585
R323 B.n731 B.n730 585
R324 B.n732 B.n731 585
R325 B.n728 B.n309 585
R326 B.n313 B.n309 585
R327 B.n727 B.n726 585
R328 B.n726 B.n725 585
R329 B.n311 B.n310 585
R330 B.n312 B.n311 585
R331 B.n718 B.n717 585
R332 B.n719 B.n718 585
R333 B.n716 B.n318 585
R334 B.n318 B.n317 585
R335 B.n715 B.n714 585
R336 B.n714 B.n713 585
R337 B.n320 B.n319 585
R338 B.n321 B.n320 585
R339 B.n707 B.n706 585
R340 B.t2 B.n707 585
R341 B.n705 B.n326 585
R342 B.n326 B.n325 585
R343 B.n704 B.n703 585
R344 B.n703 B.n702 585
R345 B.n328 B.n327 585
R346 B.n329 B.n328 585
R347 B.n695 B.n694 585
R348 B.n696 B.n695 585
R349 B.n693 B.n334 585
R350 B.n334 B.n333 585
R351 B.n692 B.n691 585
R352 B.n691 B.n690 585
R353 B.n336 B.n335 585
R354 B.n337 B.n336 585
R355 B.n683 B.n682 585
R356 B.n684 B.n683 585
R357 B.n681 B.n342 585
R358 B.n342 B.n341 585
R359 B.n680 B.n679 585
R360 B.n679 B.n678 585
R361 B.n344 B.n343 585
R362 B.n345 B.n344 585
R363 B.n671 B.n670 585
R364 B.n672 B.n671 585
R365 B.n669 B.n350 585
R366 B.n350 B.n349 585
R367 B.n668 B.n667 585
R368 B.n667 B.n666 585
R369 B.n352 B.n351 585
R370 B.n659 B.n352 585
R371 B.n658 B.n657 585
R372 B.n660 B.n658 585
R373 B.n656 B.n357 585
R374 B.n357 B.n356 585
R375 B.n655 B.n654 585
R376 B.n654 B.n653 585
R377 B.n359 B.n358 585
R378 B.n360 B.n359 585
R379 B.n646 B.n645 585
R380 B.n647 B.n646 585
R381 B.n644 B.n365 585
R382 B.n365 B.n364 585
R383 B.n643 B.n642 585
R384 B.n642 B.n641 585
R385 B.n367 B.n366 585
R386 B.n368 B.n367 585
R387 B.n634 B.n633 585
R388 B.n635 B.n634 585
R389 B.n632 B.n372 585
R390 B.n372 B.t9 585
R391 B.n631 B.n630 585
R392 B.n630 B.n629 585
R393 B.n374 B.n373 585
R394 B.n375 B.n374 585
R395 B.n622 B.n621 585
R396 B.n623 B.n622 585
R397 B.n620 B.n380 585
R398 B.n380 B.n379 585
R399 B.n619 B.n618 585
R400 B.n618 B.n617 585
R401 B.n382 B.n381 585
R402 B.n383 B.n382 585
R403 B.n610 B.n609 585
R404 B.n611 B.n610 585
R405 B.n386 B.n385 585
R406 B.n435 B.n434 585
R407 B.n436 B.n432 585
R408 B.n432 B.n387 585
R409 B.n438 B.n437 585
R410 B.n440 B.n431 585
R411 B.n443 B.n442 585
R412 B.n444 B.n430 585
R413 B.n446 B.n445 585
R414 B.n448 B.n429 585
R415 B.n451 B.n450 585
R416 B.n452 B.n428 585
R417 B.n454 B.n453 585
R418 B.n456 B.n427 585
R419 B.n459 B.n458 585
R420 B.n460 B.n426 585
R421 B.n462 B.n461 585
R422 B.n464 B.n425 585
R423 B.n467 B.n466 585
R424 B.n468 B.n424 585
R425 B.n470 B.n469 585
R426 B.n472 B.n423 585
R427 B.n475 B.n474 585
R428 B.n476 B.n422 585
R429 B.n478 B.n477 585
R430 B.n480 B.n421 585
R431 B.n483 B.n482 585
R432 B.n484 B.n420 585
R433 B.n486 B.n485 585
R434 B.n488 B.n419 585
R435 B.n491 B.n490 585
R436 B.n492 B.n418 585
R437 B.n494 B.n493 585
R438 B.n496 B.n417 585
R439 B.n499 B.n498 585
R440 B.n500 B.n416 585
R441 B.n502 B.n501 585
R442 B.n504 B.n415 585
R443 B.n507 B.n506 585
R444 B.n508 B.n412 585
R445 B.n511 B.n510 585
R446 B.n513 B.n411 585
R447 B.n516 B.n515 585
R448 B.n517 B.n410 585
R449 B.n519 B.n518 585
R450 B.n521 B.n409 585
R451 B.n524 B.n523 585
R452 B.n525 B.n408 585
R453 B.n530 B.n529 585
R454 B.n532 B.n407 585
R455 B.n535 B.n534 585
R456 B.n536 B.n406 585
R457 B.n538 B.n537 585
R458 B.n540 B.n405 585
R459 B.n543 B.n542 585
R460 B.n544 B.n404 585
R461 B.n546 B.n545 585
R462 B.n548 B.n403 585
R463 B.n551 B.n550 585
R464 B.n552 B.n402 585
R465 B.n554 B.n553 585
R466 B.n556 B.n401 585
R467 B.n559 B.n558 585
R468 B.n560 B.n400 585
R469 B.n562 B.n561 585
R470 B.n564 B.n399 585
R471 B.n567 B.n566 585
R472 B.n568 B.n398 585
R473 B.n570 B.n569 585
R474 B.n572 B.n397 585
R475 B.n575 B.n574 585
R476 B.n576 B.n396 585
R477 B.n578 B.n577 585
R478 B.n580 B.n395 585
R479 B.n583 B.n582 585
R480 B.n584 B.n394 585
R481 B.n586 B.n585 585
R482 B.n588 B.n393 585
R483 B.n591 B.n590 585
R484 B.n592 B.n392 585
R485 B.n594 B.n593 585
R486 B.n596 B.n391 585
R487 B.n599 B.n598 585
R488 B.n600 B.n390 585
R489 B.n602 B.n601 585
R490 B.n604 B.n389 585
R491 B.n607 B.n606 585
R492 B.n608 B.n388 585
R493 B.n613 B.n612 585
R494 B.n612 B.n611 585
R495 B.n614 B.n384 585
R496 B.n384 B.n383 585
R497 B.n616 B.n615 585
R498 B.n617 B.n616 585
R499 B.n378 B.n377 585
R500 B.n379 B.n378 585
R501 B.n625 B.n624 585
R502 B.n624 B.n623 585
R503 B.n626 B.n376 585
R504 B.n376 B.n375 585
R505 B.n628 B.n627 585
R506 B.n629 B.n628 585
R507 B.n371 B.n370 585
R508 B.t9 B.n371 585
R509 B.n637 B.n636 585
R510 B.n636 B.n635 585
R511 B.n638 B.n369 585
R512 B.n369 B.n368 585
R513 B.n640 B.n639 585
R514 B.n641 B.n640 585
R515 B.n363 B.n362 585
R516 B.n364 B.n363 585
R517 B.n649 B.n648 585
R518 B.n648 B.n647 585
R519 B.n650 B.n361 585
R520 B.n361 B.n360 585
R521 B.n652 B.n651 585
R522 B.n653 B.n652 585
R523 B.n355 B.n354 585
R524 B.n356 B.n355 585
R525 B.n662 B.n661 585
R526 B.n661 B.n660 585
R527 B.n663 B.n353 585
R528 B.n659 B.n353 585
R529 B.n665 B.n664 585
R530 B.n666 B.n665 585
R531 B.n348 B.n347 585
R532 B.n349 B.n348 585
R533 B.n674 B.n673 585
R534 B.n673 B.n672 585
R535 B.n675 B.n346 585
R536 B.n346 B.n345 585
R537 B.n677 B.n676 585
R538 B.n678 B.n677 585
R539 B.n340 B.n339 585
R540 B.n341 B.n340 585
R541 B.n686 B.n685 585
R542 B.n685 B.n684 585
R543 B.n687 B.n338 585
R544 B.n338 B.n337 585
R545 B.n689 B.n688 585
R546 B.n690 B.n689 585
R547 B.n332 B.n331 585
R548 B.n333 B.n332 585
R549 B.n698 B.n697 585
R550 B.n697 B.n696 585
R551 B.n699 B.n330 585
R552 B.n330 B.n329 585
R553 B.n701 B.n700 585
R554 B.n702 B.n701 585
R555 B.n324 B.n323 585
R556 B.n325 B.n324 585
R557 B.n709 B.n708 585
R558 B.n708 B.t2 585
R559 B.n710 B.n322 585
R560 B.n322 B.n321 585
R561 B.n712 B.n711 585
R562 B.n713 B.n712 585
R563 B.n316 B.n315 585
R564 B.n317 B.n316 585
R565 B.n721 B.n720 585
R566 B.n720 B.n719 585
R567 B.n722 B.n314 585
R568 B.n314 B.n312 585
R569 B.n724 B.n723 585
R570 B.n725 B.n724 585
R571 B.n308 B.n307 585
R572 B.n313 B.n308 585
R573 B.n734 B.n733 585
R574 B.n733 B.n732 585
R575 B.n735 B.n306 585
R576 B.n306 B.n305 585
R577 B.n737 B.n736 585
R578 B.n738 B.n737 585
R579 B.n3 B.n0 585
R580 B.n4 B.n3 585
R581 B.n887 B.n1 585
R582 B.n888 B.n887 585
R583 B.n886 B.n885 585
R584 B.n886 B.n8 585
R585 B.n884 B.n9 585
R586 B.n12 B.n9 585
R587 B.n883 B.n882 585
R588 B.n882 B.n881 585
R589 B.n11 B.n10 585
R590 B.n880 B.n11 585
R591 B.n878 B.n877 585
R592 B.n879 B.n878 585
R593 B.n876 B.n17 585
R594 B.n17 B.n16 585
R595 B.n875 B.n874 585
R596 B.n874 B.n873 585
R597 B.n19 B.n18 585
R598 B.n872 B.n19 585
R599 B.n870 B.n869 585
R600 B.n871 B.n870 585
R601 B.n868 B.n24 585
R602 B.n24 B.n23 585
R603 B.n867 B.n866 585
R604 B.n866 B.t1 585
R605 B.n26 B.n25 585
R606 B.n865 B.n26 585
R607 B.n863 B.n862 585
R608 B.n864 B.n863 585
R609 B.n861 B.n31 585
R610 B.n31 B.n30 585
R611 B.n860 B.n859 585
R612 B.n859 B.n858 585
R613 B.n33 B.n32 585
R614 B.n857 B.n33 585
R615 B.n855 B.n854 585
R616 B.n856 B.n855 585
R617 B.n853 B.n38 585
R618 B.n38 B.n37 585
R619 B.n852 B.n851 585
R620 B.n851 B.n850 585
R621 B.n40 B.n39 585
R622 B.n849 B.n40 585
R623 B.n847 B.n846 585
R624 B.n848 B.n847 585
R625 B.n845 B.n45 585
R626 B.n45 B.n44 585
R627 B.n844 B.n843 585
R628 B.n843 B.n842 585
R629 B.n47 B.n46 585
R630 B.n841 B.n47 585
R631 B.n839 B.n838 585
R632 B.n840 B.n839 585
R633 B.n837 B.n51 585
R634 B.n54 B.n51 585
R635 B.n836 B.n835 585
R636 B.n835 B.n834 585
R637 B.n53 B.n52 585
R638 B.n833 B.n53 585
R639 B.n831 B.n830 585
R640 B.n832 B.n831 585
R641 B.n829 B.n59 585
R642 B.n59 B.n58 585
R643 B.n828 B.n827 585
R644 B.n827 B.n826 585
R645 B.n61 B.n60 585
R646 B.n825 B.n61 585
R647 B.n823 B.n822 585
R648 B.n824 B.n823 585
R649 B.n821 B.n66 585
R650 B.n66 B.n65 585
R651 B.n820 B.n819 585
R652 B.n819 B.n818 585
R653 B.n68 B.n67 585
R654 B.t13 B.n68 585
R655 B.n816 B.n815 585
R656 B.n817 B.n816 585
R657 B.n814 B.n73 585
R658 B.n73 B.n72 585
R659 B.n813 B.n812 585
R660 B.n812 B.n811 585
R661 B.n75 B.n74 585
R662 B.n810 B.n75 585
R663 B.n808 B.n807 585
R664 B.n809 B.n808 585
R665 B.n806 B.n80 585
R666 B.n80 B.n79 585
R667 B.n805 B.n804 585
R668 B.n804 B.n803 585
R669 B.n891 B.n890 585
R670 B.n889 B.n2 585
R671 B.n804 B.n82 449.257
R672 B.n801 B.n83 449.257
R673 B.n610 B.n388 449.257
R674 B.n612 B.n386 449.257
R675 B.n131 B.t12 330.318
R676 B.n128 B.t19 330.318
R677 B.n526 B.t16 330.318
R678 B.n413 B.t8 330.318
R679 B.n802 B.n126 256.663
R680 B.n802 B.n125 256.663
R681 B.n802 B.n124 256.663
R682 B.n802 B.n123 256.663
R683 B.n802 B.n122 256.663
R684 B.n802 B.n121 256.663
R685 B.n802 B.n120 256.663
R686 B.n802 B.n119 256.663
R687 B.n802 B.n118 256.663
R688 B.n802 B.n117 256.663
R689 B.n802 B.n116 256.663
R690 B.n802 B.n115 256.663
R691 B.n802 B.n114 256.663
R692 B.n802 B.n113 256.663
R693 B.n802 B.n112 256.663
R694 B.n802 B.n111 256.663
R695 B.n802 B.n110 256.663
R696 B.n802 B.n109 256.663
R697 B.n802 B.n108 256.663
R698 B.n802 B.n107 256.663
R699 B.n802 B.n106 256.663
R700 B.n802 B.n105 256.663
R701 B.n802 B.n104 256.663
R702 B.n802 B.n103 256.663
R703 B.n802 B.n102 256.663
R704 B.n802 B.n101 256.663
R705 B.n802 B.n100 256.663
R706 B.n802 B.n99 256.663
R707 B.n802 B.n98 256.663
R708 B.n802 B.n97 256.663
R709 B.n802 B.n96 256.663
R710 B.n802 B.n95 256.663
R711 B.n802 B.n94 256.663
R712 B.n802 B.n93 256.663
R713 B.n802 B.n92 256.663
R714 B.n802 B.n91 256.663
R715 B.n802 B.n90 256.663
R716 B.n802 B.n89 256.663
R717 B.n802 B.n88 256.663
R718 B.n802 B.n87 256.663
R719 B.n802 B.n86 256.663
R720 B.n802 B.n85 256.663
R721 B.n802 B.n84 256.663
R722 B.n433 B.n387 256.663
R723 B.n439 B.n387 256.663
R724 B.n441 B.n387 256.663
R725 B.n447 B.n387 256.663
R726 B.n449 B.n387 256.663
R727 B.n455 B.n387 256.663
R728 B.n457 B.n387 256.663
R729 B.n463 B.n387 256.663
R730 B.n465 B.n387 256.663
R731 B.n471 B.n387 256.663
R732 B.n473 B.n387 256.663
R733 B.n479 B.n387 256.663
R734 B.n481 B.n387 256.663
R735 B.n487 B.n387 256.663
R736 B.n489 B.n387 256.663
R737 B.n495 B.n387 256.663
R738 B.n497 B.n387 256.663
R739 B.n503 B.n387 256.663
R740 B.n505 B.n387 256.663
R741 B.n512 B.n387 256.663
R742 B.n514 B.n387 256.663
R743 B.n520 B.n387 256.663
R744 B.n522 B.n387 256.663
R745 B.n531 B.n387 256.663
R746 B.n533 B.n387 256.663
R747 B.n539 B.n387 256.663
R748 B.n541 B.n387 256.663
R749 B.n547 B.n387 256.663
R750 B.n549 B.n387 256.663
R751 B.n555 B.n387 256.663
R752 B.n557 B.n387 256.663
R753 B.n563 B.n387 256.663
R754 B.n565 B.n387 256.663
R755 B.n571 B.n387 256.663
R756 B.n573 B.n387 256.663
R757 B.n579 B.n387 256.663
R758 B.n581 B.n387 256.663
R759 B.n587 B.n387 256.663
R760 B.n589 B.n387 256.663
R761 B.n595 B.n387 256.663
R762 B.n597 B.n387 256.663
R763 B.n603 B.n387 256.663
R764 B.n605 B.n387 256.663
R765 B.n893 B.n892 256.663
R766 B.n135 B.n134 163.367
R767 B.n139 B.n138 163.367
R768 B.n143 B.n142 163.367
R769 B.n147 B.n146 163.367
R770 B.n151 B.n150 163.367
R771 B.n155 B.n154 163.367
R772 B.n159 B.n158 163.367
R773 B.n163 B.n162 163.367
R774 B.n167 B.n166 163.367
R775 B.n171 B.n170 163.367
R776 B.n175 B.n174 163.367
R777 B.n179 B.n178 163.367
R778 B.n183 B.n182 163.367
R779 B.n187 B.n186 163.367
R780 B.n191 B.n190 163.367
R781 B.n195 B.n194 163.367
R782 B.n199 B.n198 163.367
R783 B.n203 B.n202 163.367
R784 B.n207 B.n206 163.367
R785 B.n212 B.n211 163.367
R786 B.n216 B.n215 163.367
R787 B.n220 B.n219 163.367
R788 B.n224 B.n223 163.367
R789 B.n228 B.n227 163.367
R790 B.n232 B.n231 163.367
R791 B.n236 B.n235 163.367
R792 B.n240 B.n239 163.367
R793 B.n244 B.n243 163.367
R794 B.n248 B.n247 163.367
R795 B.n252 B.n251 163.367
R796 B.n256 B.n255 163.367
R797 B.n260 B.n259 163.367
R798 B.n264 B.n263 163.367
R799 B.n268 B.n267 163.367
R800 B.n272 B.n271 163.367
R801 B.n276 B.n275 163.367
R802 B.n280 B.n279 163.367
R803 B.n284 B.n283 163.367
R804 B.n288 B.n287 163.367
R805 B.n292 B.n291 163.367
R806 B.n296 B.n295 163.367
R807 B.n300 B.n299 163.367
R808 B.n801 B.n127 163.367
R809 B.n610 B.n382 163.367
R810 B.n618 B.n382 163.367
R811 B.n618 B.n380 163.367
R812 B.n622 B.n380 163.367
R813 B.n622 B.n374 163.367
R814 B.n630 B.n374 163.367
R815 B.n630 B.n372 163.367
R816 B.n634 B.n372 163.367
R817 B.n634 B.n367 163.367
R818 B.n642 B.n367 163.367
R819 B.n642 B.n365 163.367
R820 B.n646 B.n365 163.367
R821 B.n646 B.n359 163.367
R822 B.n654 B.n359 163.367
R823 B.n654 B.n357 163.367
R824 B.n658 B.n357 163.367
R825 B.n658 B.n352 163.367
R826 B.n667 B.n352 163.367
R827 B.n667 B.n350 163.367
R828 B.n671 B.n350 163.367
R829 B.n671 B.n344 163.367
R830 B.n679 B.n344 163.367
R831 B.n679 B.n342 163.367
R832 B.n683 B.n342 163.367
R833 B.n683 B.n336 163.367
R834 B.n691 B.n336 163.367
R835 B.n691 B.n334 163.367
R836 B.n695 B.n334 163.367
R837 B.n695 B.n328 163.367
R838 B.n703 B.n328 163.367
R839 B.n703 B.n326 163.367
R840 B.n707 B.n326 163.367
R841 B.n707 B.n320 163.367
R842 B.n714 B.n320 163.367
R843 B.n714 B.n318 163.367
R844 B.n718 B.n318 163.367
R845 B.n718 B.n311 163.367
R846 B.n726 B.n311 163.367
R847 B.n726 B.n309 163.367
R848 B.n731 B.n309 163.367
R849 B.n731 B.n304 163.367
R850 B.n739 B.n304 163.367
R851 B.n740 B.n739 163.367
R852 B.n740 B.n5 163.367
R853 B.n6 B.n5 163.367
R854 B.n7 B.n6 163.367
R855 B.n746 B.n7 163.367
R856 B.n747 B.n746 163.367
R857 B.n747 B.n13 163.367
R858 B.n14 B.n13 163.367
R859 B.n15 B.n14 163.367
R860 B.n752 B.n15 163.367
R861 B.n752 B.n20 163.367
R862 B.n21 B.n20 163.367
R863 B.n22 B.n21 163.367
R864 B.n757 B.n22 163.367
R865 B.n757 B.n27 163.367
R866 B.n28 B.n27 163.367
R867 B.n29 B.n28 163.367
R868 B.n762 B.n29 163.367
R869 B.n762 B.n34 163.367
R870 B.n35 B.n34 163.367
R871 B.n36 B.n35 163.367
R872 B.n767 B.n36 163.367
R873 B.n767 B.n41 163.367
R874 B.n42 B.n41 163.367
R875 B.n43 B.n42 163.367
R876 B.n772 B.n43 163.367
R877 B.n772 B.n48 163.367
R878 B.n49 B.n48 163.367
R879 B.n50 B.n49 163.367
R880 B.n777 B.n50 163.367
R881 B.n777 B.n55 163.367
R882 B.n56 B.n55 163.367
R883 B.n57 B.n56 163.367
R884 B.n782 B.n57 163.367
R885 B.n782 B.n62 163.367
R886 B.n63 B.n62 163.367
R887 B.n64 B.n63 163.367
R888 B.n787 B.n64 163.367
R889 B.n787 B.n69 163.367
R890 B.n70 B.n69 163.367
R891 B.n71 B.n70 163.367
R892 B.n792 B.n71 163.367
R893 B.n792 B.n76 163.367
R894 B.n77 B.n76 163.367
R895 B.n78 B.n77 163.367
R896 B.n797 B.n78 163.367
R897 B.n797 B.n83 163.367
R898 B.n434 B.n432 163.367
R899 B.n438 B.n432 163.367
R900 B.n442 B.n440 163.367
R901 B.n446 B.n430 163.367
R902 B.n450 B.n448 163.367
R903 B.n454 B.n428 163.367
R904 B.n458 B.n456 163.367
R905 B.n462 B.n426 163.367
R906 B.n466 B.n464 163.367
R907 B.n470 B.n424 163.367
R908 B.n474 B.n472 163.367
R909 B.n478 B.n422 163.367
R910 B.n482 B.n480 163.367
R911 B.n486 B.n420 163.367
R912 B.n490 B.n488 163.367
R913 B.n494 B.n418 163.367
R914 B.n498 B.n496 163.367
R915 B.n502 B.n416 163.367
R916 B.n506 B.n504 163.367
R917 B.n511 B.n412 163.367
R918 B.n515 B.n513 163.367
R919 B.n519 B.n410 163.367
R920 B.n523 B.n521 163.367
R921 B.n530 B.n408 163.367
R922 B.n534 B.n532 163.367
R923 B.n538 B.n406 163.367
R924 B.n542 B.n540 163.367
R925 B.n546 B.n404 163.367
R926 B.n550 B.n548 163.367
R927 B.n554 B.n402 163.367
R928 B.n558 B.n556 163.367
R929 B.n562 B.n400 163.367
R930 B.n566 B.n564 163.367
R931 B.n570 B.n398 163.367
R932 B.n574 B.n572 163.367
R933 B.n578 B.n396 163.367
R934 B.n582 B.n580 163.367
R935 B.n586 B.n394 163.367
R936 B.n590 B.n588 163.367
R937 B.n594 B.n392 163.367
R938 B.n598 B.n596 163.367
R939 B.n602 B.n390 163.367
R940 B.n606 B.n604 163.367
R941 B.n612 B.n384 163.367
R942 B.n616 B.n384 163.367
R943 B.n616 B.n378 163.367
R944 B.n624 B.n378 163.367
R945 B.n624 B.n376 163.367
R946 B.n628 B.n376 163.367
R947 B.n628 B.n371 163.367
R948 B.n636 B.n371 163.367
R949 B.n636 B.n369 163.367
R950 B.n640 B.n369 163.367
R951 B.n640 B.n363 163.367
R952 B.n648 B.n363 163.367
R953 B.n648 B.n361 163.367
R954 B.n652 B.n361 163.367
R955 B.n652 B.n355 163.367
R956 B.n661 B.n355 163.367
R957 B.n661 B.n353 163.367
R958 B.n665 B.n353 163.367
R959 B.n665 B.n348 163.367
R960 B.n673 B.n348 163.367
R961 B.n673 B.n346 163.367
R962 B.n677 B.n346 163.367
R963 B.n677 B.n340 163.367
R964 B.n685 B.n340 163.367
R965 B.n685 B.n338 163.367
R966 B.n689 B.n338 163.367
R967 B.n689 B.n332 163.367
R968 B.n697 B.n332 163.367
R969 B.n697 B.n330 163.367
R970 B.n701 B.n330 163.367
R971 B.n701 B.n324 163.367
R972 B.n708 B.n324 163.367
R973 B.n708 B.n322 163.367
R974 B.n712 B.n322 163.367
R975 B.n712 B.n316 163.367
R976 B.n720 B.n316 163.367
R977 B.n720 B.n314 163.367
R978 B.n724 B.n314 163.367
R979 B.n724 B.n308 163.367
R980 B.n733 B.n308 163.367
R981 B.n733 B.n306 163.367
R982 B.n737 B.n306 163.367
R983 B.n737 B.n3 163.367
R984 B.n891 B.n3 163.367
R985 B.n887 B.n2 163.367
R986 B.n887 B.n886 163.367
R987 B.n886 B.n9 163.367
R988 B.n882 B.n9 163.367
R989 B.n882 B.n11 163.367
R990 B.n878 B.n11 163.367
R991 B.n878 B.n17 163.367
R992 B.n874 B.n17 163.367
R993 B.n874 B.n19 163.367
R994 B.n870 B.n19 163.367
R995 B.n870 B.n24 163.367
R996 B.n866 B.n24 163.367
R997 B.n866 B.n26 163.367
R998 B.n863 B.n26 163.367
R999 B.n863 B.n31 163.367
R1000 B.n859 B.n31 163.367
R1001 B.n859 B.n33 163.367
R1002 B.n855 B.n33 163.367
R1003 B.n855 B.n38 163.367
R1004 B.n851 B.n38 163.367
R1005 B.n851 B.n40 163.367
R1006 B.n847 B.n40 163.367
R1007 B.n847 B.n45 163.367
R1008 B.n843 B.n45 163.367
R1009 B.n843 B.n47 163.367
R1010 B.n839 B.n47 163.367
R1011 B.n839 B.n51 163.367
R1012 B.n835 B.n51 163.367
R1013 B.n835 B.n53 163.367
R1014 B.n831 B.n53 163.367
R1015 B.n831 B.n59 163.367
R1016 B.n827 B.n59 163.367
R1017 B.n827 B.n61 163.367
R1018 B.n823 B.n61 163.367
R1019 B.n823 B.n66 163.367
R1020 B.n819 B.n66 163.367
R1021 B.n819 B.n68 163.367
R1022 B.n816 B.n68 163.367
R1023 B.n816 B.n73 163.367
R1024 B.n812 B.n73 163.367
R1025 B.n812 B.n75 163.367
R1026 B.n808 B.n75 163.367
R1027 B.n808 B.n80 163.367
R1028 B.n804 B.n80 163.367
R1029 B.n128 B.t20 116.823
R1030 B.n526 B.t18 116.823
R1031 B.n131 B.t14 116.808
R1032 B.n413 B.t11 116.808
R1033 B.n611 B.n387 80.778
R1034 B.n803 B.n802 80.778
R1035 B.n84 B.n82 71.676
R1036 B.n135 B.n85 71.676
R1037 B.n139 B.n86 71.676
R1038 B.n143 B.n87 71.676
R1039 B.n147 B.n88 71.676
R1040 B.n151 B.n89 71.676
R1041 B.n155 B.n90 71.676
R1042 B.n159 B.n91 71.676
R1043 B.n163 B.n92 71.676
R1044 B.n167 B.n93 71.676
R1045 B.n171 B.n94 71.676
R1046 B.n175 B.n95 71.676
R1047 B.n179 B.n96 71.676
R1048 B.n183 B.n97 71.676
R1049 B.n187 B.n98 71.676
R1050 B.n191 B.n99 71.676
R1051 B.n195 B.n100 71.676
R1052 B.n199 B.n101 71.676
R1053 B.n203 B.n102 71.676
R1054 B.n207 B.n103 71.676
R1055 B.n212 B.n104 71.676
R1056 B.n216 B.n105 71.676
R1057 B.n220 B.n106 71.676
R1058 B.n224 B.n107 71.676
R1059 B.n228 B.n108 71.676
R1060 B.n232 B.n109 71.676
R1061 B.n236 B.n110 71.676
R1062 B.n240 B.n111 71.676
R1063 B.n244 B.n112 71.676
R1064 B.n248 B.n113 71.676
R1065 B.n252 B.n114 71.676
R1066 B.n256 B.n115 71.676
R1067 B.n260 B.n116 71.676
R1068 B.n264 B.n117 71.676
R1069 B.n268 B.n118 71.676
R1070 B.n272 B.n119 71.676
R1071 B.n276 B.n120 71.676
R1072 B.n280 B.n121 71.676
R1073 B.n284 B.n122 71.676
R1074 B.n288 B.n123 71.676
R1075 B.n292 B.n124 71.676
R1076 B.n296 B.n125 71.676
R1077 B.n300 B.n126 71.676
R1078 B.n127 B.n126 71.676
R1079 B.n299 B.n125 71.676
R1080 B.n295 B.n124 71.676
R1081 B.n291 B.n123 71.676
R1082 B.n287 B.n122 71.676
R1083 B.n283 B.n121 71.676
R1084 B.n279 B.n120 71.676
R1085 B.n275 B.n119 71.676
R1086 B.n271 B.n118 71.676
R1087 B.n267 B.n117 71.676
R1088 B.n263 B.n116 71.676
R1089 B.n259 B.n115 71.676
R1090 B.n255 B.n114 71.676
R1091 B.n251 B.n113 71.676
R1092 B.n247 B.n112 71.676
R1093 B.n243 B.n111 71.676
R1094 B.n239 B.n110 71.676
R1095 B.n235 B.n109 71.676
R1096 B.n231 B.n108 71.676
R1097 B.n227 B.n107 71.676
R1098 B.n223 B.n106 71.676
R1099 B.n219 B.n105 71.676
R1100 B.n215 B.n104 71.676
R1101 B.n211 B.n103 71.676
R1102 B.n206 B.n102 71.676
R1103 B.n202 B.n101 71.676
R1104 B.n198 B.n100 71.676
R1105 B.n194 B.n99 71.676
R1106 B.n190 B.n98 71.676
R1107 B.n186 B.n97 71.676
R1108 B.n182 B.n96 71.676
R1109 B.n178 B.n95 71.676
R1110 B.n174 B.n94 71.676
R1111 B.n170 B.n93 71.676
R1112 B.n166 B.n92 71.676
R1113 B.n162 B.n91 71.676
R1114 B.n158 B.n90 71.676
R1115 B.n154 B.n89 71.676
R1116 B.n150 B.n88 71.676
R1117 B.n146 B.n87 71.676
R1118 B.n142 B.n86 71.676
R1119 B.n138 B.n85 71.676
R1120 B.n134 B.n84 71.676
R1121 B.n433 B.n386 71.676
R1122 B.n439 B.n438 71.676
R1123 B.n442 B.n441 71.676
R1124 B.n447 B.n446 71.676
R1125 B.n450 B.n449 71.676
R1126 B.n455 B.n454 71.676
R1127 B.n458 B.n457 71.676
R1128 B.n463 B.n462 71.676
R1129 B.n466 B.n465 71.676
R1130 B.n471 B.n470 71.676
R1131 B.n474 B.n473 71.676
R1132 B.n479 B.n478 71.676
R1133 B.n482 B.n481 71.676
R1134 B.n487 B.n486 71.676
R1135 B.n490 B.n489 71.676
R1136 B.n495 B.n494 71.676
R1137 B.n498 B.n497 71.676
R1138 B.n503 B.n502 71.676
R1139 B.n506 B.n505 71.676
R1140 B.n512 B.n511 71.676
R1141 B.n515 B.n514 71.676
R1142 B.n520 B.n519 71.676
R1143 B.n523 B.n522 71.676
R1144 B.n531 B.n530 71.676
R1145 B.n534 B.n533 71.676
R1146 B.n539 B.n538 71.676
R1147 B.n542 B.n541 71.676
R1148 B.n547 B.n546 71.676
R1149 B.n550 B.n549 71.676
R1150 B.n555 B.n554 71.676
R1151 B.n558 B.n557 71.676
R1152 B.n563 B.n562 71.676
R1153 B.n566 B.n565 71.676
R1154 B.n571 B.n570 71.676
R1155 B.n574 B.n573 71.676
R1156 B.n579 B.n578 71.676
R1157 B.n582 B.n581 71.676
R1158 B.n587 B.n586 71.676
R1159 B.n590 B.n589 71.676
R1160 B.n595 B.n594 71.676
R1161 B.n598 B.n597 71.676
R1162 B.n603 B.n602 71.676
R1163 B.n606 B.n605 71.676
R1164 B.n434 B.n433 71.676
R1165 B.n440 B.n439 71.676
R1166 B.n441 B.n430 71.676
R1167 B.n448 B.n447 71.676
R1168 B.n449 B.n428 71.676
R1169 B.n456 B.n455 71.676
R1170 B.n457 B.n426 71.676
R1171 B.n464 B.n463 71.676
R1172 B.n465 B.n424 71.676
R1173 B.n472 B.n471 71.676
R1174 B.n473 B.n422 71.676
R1175 B.n480 B.n479 71.676
R1176 B.n481 B.n420 71.676
R1177 B.n488 B.n487 71.676
R1178 B.n489 B.n418 71.676
R1179 B.n496 B.n495 71.676
R1180 B.n497 B.n416 71.676
R1181 B.n504 B.n503 71.676
R1182 B.n505 B.n412 71.676
R1183 B.n513 B.n512 71.676
R1184 B.n514 B.n410 71.676
R1185 B.n521 B.n520 71.676
R1186 B.n522 B.n408 71.676
R1187 B.n532 B.n531 71.676
R1188 B.n533 B.n406 71.676
R1189 B.n540 B.n539 71.676
R1190 B.n541 B.n404 71.676
R1191 B.n548 B.n547 71.676
R1192 B.n549 B.n402 71.676
R1193 B.n556 B.n555 71.676
R1194 B.n557 B.n400 71.676
R1195 B.n564 B.n563 71.676
R1196 B.n565 B.n398 71.676
R1197 B.n572 B.n571 71.676
R1198 B.n573 B.n396 71.676
R1199 B.n580 B.n579 71.676
R1200 B.n581 B.n394 71.676
R1201 B.n588 B.n587 71.676
R1202 B.n589 B.n392 71.676
R1203 B.n596 B.n595 71.676
R1204 B.n597 B.n390 71.676
R1205 B.n604 B.n603 71.676
R1206 B.n605 B.n388 71.676
R1207 B.n892 B.n891 71.676
R1208 B.n892 B.n2 71.676
R1209 B.n129 B.t21 68.9196
R1210 B.n527 B.t17 68.9196
R1211 B.n132 B.t15 68.9059
R1212 B.n414 B.t10 68.9059
R1213 B.n209 B.n132 59.5399
R1214 B.n130 B.n129 59.5399
R1215 B.n528 B.n527 59.5399
R1216 B.n509 B.n414 59.5399
R1217 B.n132 B.n131 47.9035
R1218 B.n129 B.n128 47.9035
R1219 B.n527 B.n526 47.9035
R1220 B.n414 B.n413 47.9035
R1221 B.n611 B.n383 46.1591
R1222 B.n617 B.n383 46.1591
R1223 B.n617 B.n379 46.1591
R1224 B.n623 B.n379 46.1591
R1225 B.n623 B.n375 46.1591
R1226 B.n629 B.n375 46.1591
R1227 B.n629 B.t9 46.1591
R1228 B.n635 B.t9 46.1591
R1229 B.n635 B.n368 46.1591
R1230 B.n641 B.n368 46.1591
R1231 B.n641 B.n364 46.1591
R1232 B.n647 B.n364 46.1591
R1233 B.n647 B.n360 46.1591
R1234 B.n653 B.n360 46.1591
R1235 B.n653 B.n356 46.1591
R1236 B.n660 B.n356 46.1591
R1237 B.n660 B.n659 46.1591
R1238 B.n666 B.n349 46.1591
R1239 B.n672 B.n349 46.1591
R1240 B.n672 B.n345 46.1591
R1241 B.n678 B.n345 46.1591
R1242 B.n678 B.n341 46.1591
R1243 B.n684 B.n341 46.1591
R1244 B.n690 B.n337 46.1591
R1245 B.n690 B.n333 46.1591
R1246 B.n696 B.n333 46.1591
R1247 B.n696 B.n329 46.1591
R1248 B.n702 B.n329 46.1591
R1249 B.n702 B.n325 46.1591
R1250 B.t2 B.n325 46.1591
R1251 B.t2 B.n321 46.1591
R1252 B.n713 B.n321 46.1591
R1253 B.n713 B.n317 46.1591
R1254 B.n719 B.n317 46.1591
R1255 B.n719 B.n312 46.1591
R1256 B.n725 B.n312 46.1591
R1257 B.n725 B.n313 46.1591
R1258 B.n732 B.n305 46.1591
R1259 B.n738 B.n305 46.1591
R1260 B.n738 B.n4 46.1591
R1261 B.n890 B.n4 46.1591
R1262 B.n890 B.n889 46.1591
R1263 B.n889 B.n888 46.1591
R1264 B.n888 B.n8 46.1591
R1265 B.n12 B.n8 46.1591
R1266 B.n881 B.n12 46.1591
R1267 B.n880 B.n879 46.1591
R1268 B.n879 B.n16 46.1591
R1269 B.n873 B.n16 46.1591
R1270 B.n873 B.n872 46.1591
R1271 B.n872 B.n871 46.1591
R1272 B.n871 B.n23 46.1591
R1273 B.t1 B.n23 46.1591
R1274 B.t1 B.n865 46.1591
R1275 B.n865 B.n864 46.1591
R1276 B.n864 B.n30 46.1591
R1277 B.n858 B.n30 46.1591
R1278 B.n858 B.n857 46.1591
R1279 B.n857 B.n856 46.1591
R1280 B.n856 B.n37 46.1591
R1281 B.n850 B.n849 46.1591
R1282 B.n849 B.n848 46.1591
R1283 B.n848 B.n44 46.1591
R1284 B.n842 B.n44 46.1591
R1285 B.n842 B.n841 46.1591
R1286 B.n841 B.n840 46.1591
R1287 B.n834 B.n54 46.1591
R1288 B.n834 B.n833 46.1591
R1289 B.n833 B.n832 46.1591
R1290 B.n832 B.n58 46.1591
R1291 B.n826 B.n58 46.1591
R1292 B.n826 B.n825 46.1591
R1293 B.n825 B.n824 46.1591
R1294 B.n824 B.n65 46.1591
R1295 B.n818 B.n65 46.1591
R1296 B.n818 B.t13 46.1591
R1297 B.t13 B.n817 46.1591
R1298 B.n817 B.n72 46.1591
R1299 B.n811 B.n72 46.1591
R1300 B.n811 B.n810 46.1591
R1301 B.n810 B.n809 46.1591
R1302 B.n809 B.n79 46.1591
R1303 B.n803 B.n79 46.1591
R1304 B.n684 B.t0 33.9406
R1305 B.n732 B.t3 33.9406
R1306 B.n881 B.t5 33.9406
R1307 B.n850 B.t6 33.9406
R1308 B.n800 B.n799 29.1907
R1309 B.n613 B.n385 29.1907
R1310 B.n609 B.n608 29.1907
R1311 B.n805 B.n81 29.1907
R1312 B.n666 B.t7 24.4374
R1313 B.n840 B.t4 24.4374
R1314 B.n659 B.t7 21.7222
R1315 B.n54 B.t4 21.7222
R1316 B B.n893 18.0485
R1317 B.t0 B.n337 12.219
R1318 B.n313 B.t3 12.219
R1319 B.t5 B.n880 12.219
R1320 B.t6 B.n37 12.219
R1321 B.n614 B.n613 10.6151
R1322 B.n615 B.n614 10.6151
R1323 B.n615 B.n377 10.6151
R1324 B.n625 B.n377 10.6151
R1325 B.n626 B.n625 10.6151
R1326 B.n627 B.n626 10.6151
R1327 B.n627 B.n370 10.6151
R1328 B.n637 B.n370 10.6151
R1329 B.n638 B.n637 10.6151
R1330 B.n639 B.n638 10.6151
R1331 B.n639 B.n362 10.6151
R1332 B.n649 B.n362 10.6151
R1333 B.n650 B.n649 10.6151
R1334 B.n651 B.n650 10.6151
R1335 B.n651 B.n354 10.6151
R1336 B.n662 B.n354 10.6151
R1337 B.n663 B.n662 10.6151
R1338 B.n664 B.n663 10.6151
R1339 B.n664 B.n347 10.6151
R1340 B.n674 B.n347 10.6151
R1341 B.n675 B.n674 10.6151
R1342 B.n676 B.n675 10.6151
R1343 B.n676 B.n339 10.6151
R1344 B.n686 B.n339 10.6151
R1345 B.n687 B.n686 10.6151
R1346 B.n688 B.n687 10.6151
R1347 B.n688 B.n331 10.6151
R1348 B.n698 B.n331 10.6151
R1349 B.n699 B.n698 10.6151
R1350 B.n700 B.n699 10.6151
R1351 B.n700 B.n323 10.6151
R1352 B.n709 B.n323 10.6151
R1353 B.n710 B.n709 10.6151
R1354 B.n711 B.n710 10.6151
R1355 B.n711 B.n315 10.6151
R1356 B.n721 B.n315 10.6151
R1357 B.n722 B.n721 10.6151
R1358 B.n723 B.n722 10.6151
R1359 B.n723 B.n307 10.6151
R1360 B.n734 B.n307 10.6151
R1361 B.n735 B.n734 10.6151
R1362 B.n736 B.n735 10.6151
R1363 B.n736 B.n0 10.6151
R1364 B.n435 B.n385 10.6151
R1365 B.n436 B.n435 10.6151
R1366 B.n437 B.n436 10.6151
R1367 B.n437 B.n431 10.6151
R1368 B.n443 B.n431 10.6151
R1369 B.n444 B.n443 10.6151
R1370 B.n445 B.n444 10.6151
R1371 B.n445 B.n429 10.6151
R1372 B.n451 B.n429 10.6151
R1373 B.n452 B.n451 10.6151
R1374 B.n453 B.n452 10.6151
R1375 B.n453 B.n427 10.6151
R1376 B.n459 B.n427 10.6151
R1377 B.n460 B.n459 10.6151
R1378 B.n461 B.n460 10.6151
R1379 B.n461 B.n425 10.6151
R1380 B.n467 B.n425 10.6151
R1381 B.n468 B.n467 10.6151
R1382 B.n469 B.n468 10.6151
R1383 B.n469 B.n423 10.6151
R1384 B.n475 B.n423 10.6151
R1385 B.n476 B.n475 10.6151
R1386 B.n477 B.n476 10.6151
R1387 B.n477 B.n421 10.6151
R1388 B.n483 B.n421 10.6151
R1389 B.n484 B.n483 10.6151
R1390 B.n485 B.n484 10.6151
R1391 B.n485 B.n419 10.6151
R1392 B.n491 B.n419 10.6151
R1393 B.n492 B.n491 10.6151
R1394 B.n493 B.n492 10.6151
R1395 B.n493 B.n417 10.6151
R1396 B.n499 B.n417 10.6151
R1397 B.n500 B.n499 10.6151
R1398 B.n501 B.n500 10.6151
R1399 B.n501 B.n415 10.6151
R1400 B.n507 B.n415 10.6151
R1401 B.n508 B.n507 10.6151
R1402 B.n510 B.n411 10.6151
R1403 B.n516 B.n411 10.6151
R1404 B.n517 B.n516 10.6151
R1405 B.n518 B.n517 10.6151
R1406 B.n518 B.n409 10.6151
R1407 B.n524 B.n409 10.6151
R1408 B.n525 B.n524 10.6151
R1409 B.n529 B.n525 10.6151
R1410 B.n535 B.n407 10.6151
R1411 B.n536 B.n535 10.6151
R1412 B.n537 B.n536 10.6151
R1413 B.n537 B.n405 10.6151
R1414 B.n543 B.n405 10.6151
R1415 B.n544 B.n543 10.6151
R1416 B.n545 B.n544 10.6151
R1417 B.n545 B.n403 10.6151
R1418 B.n551 B.n403 10.6151
R1419 B.n552 B.n551 10.6151
R1420 B.n553 B.n552 10.6151
R1421 B.n553 B.n401 10.6151
R1422 B.n559 B.n401 10.6151
R1423 B.n560 B.n559 10.6151
R1424 B.n561 B.n560 10.6151
R1425 B.n561 B.n399 10.6151
R1426 B.n567 B.n399 10.6151
R1427 B.n568 B.n567 10.6151
R1428 B.n569 B.n568 10.6151
R1429 B.n569 B.n397 10.6151
R1430 B.n575 B.n397 10.6151
R1431 B.n576 B.n575 10.6151
R1432 B.n577 B.n576 10.6151
R1433 B.n577 B.n395 10.6151
R1434 B.n583 B.n395 10.6151
R1435 B.n584 B.n583 10.6151
R1436 B.n585 B.n584 10.6151
R1437 B.n585 B.n393 10.6151
R1438 B.n591 B.n393 10.6151
R1439 B.n592 B.n591 10.6151
R1440 B.n593 B.n592 10.6151
R1441 B.n593 B.n391 10.6151
R1442 B.n599 B.n391 10.6151
R1443 B.n600 B.n599 10.6151
R1444 B.n601 B.n600 10.6151
R1445 B.n601 B.n389 10.6151
R1446 B.n607 B.n389 10.6151
R1447 B.n608 B.n607 10.6151
R1448 B.n609 B.n381 10.6151
R1449 B.n619 B.n381 10.6151
R1450 B.n620 B.n619 10.6151
R1451 B.n621 B.n620 10.6151
R1452 B.n621 B.n373 10.6151
R1453 B.n631 B.n373 10.6151
R1454 B.n632 B.n631 10.6151
R1455 B.n633 B.n632 10.6151
R1456 B.n633 B.n366 10.6151
R1457 B.n643 B.n366 10.6151
R1458 B.n644 B.n643 10.6151
R1459 B.n645 B.n644 10.6151
R1460 B.n645 B.n358 10.6151
R1461 B.n655 B.n358 10.6151
R1462 B.n656 B.n655 10.6151
R1463 B.n657 B.n656 10.6151
R1464 B.n657 B.n351 10.6151
R1465 B.n668 B.n351 10.6151
R1466 B.n669 B.n668 10.6151
R1467 B.n670 B.n669 10.6151
R1468 B.n670 B.n343 10.6151
R1469 B.n680 B.n343 10.6151
R1470 B.n681 B.n680 10.6151
R1471 B.n682 B.n681 10.6151
R1472 B.n682 B.n335 10.6151
R1473 B.n692 B.n335 10.6151
R1474 B.n693 B.n692 10.6151
R1475 B.n694 B.n693 10.6151
R1476 B.n694 B.n327 10.6151
R1477 B.n704 B.n327 10.6151
R1478 B.n705 B.n704 10.6151
R1479 B.n706 B.n705 10.6151
R1480 B.n706 B.n319 10.6151
R1481 B.n715 B.n319 10.6151
R1482 B.n716 B.n715 10.6151
R1483 B.n717 B.n716 10.6151
R1484 B.n717 B.n310 10.6151
R1485 B.n727 B.n310 10.6151
R1486 B.n728 B.n727 10.6151
R1487 B.n730 B.n728 10.6151
R1488 B.n730 B.n729 10.6151
R1489 B.n729 B.n303 10.6151
R1490 B.n741 B.n303 10.6151
R1491 B.n742 B.n741 10.6151
R1492 B.n743 B.n742 10.6151
R1493 B.n744 B.n743 10.6151
R1494 B.n745 B.n744 10.6151
R1495 B.n748 B.n745 10.6151
R1496 B.n749 B.n748 10.6151
R1497 B.n750 B.n749 10.6151
R1498 B.n751 B.n750 10.6151
R1499 B.n753 B.n751 10.6151
R1500 B.n754 B.n753 10.6151
R1501 B.n755 B.n754 10.6151
R1502 B.n756 B.n755 10.6151
R1503 B.n758 B.n756 10.6151
R1504 B.n759 B.n758 10.6151
R1505 B.n760 B.n759 10.6151
R1506 B.n761 B.n760 10.6151
R1507 B.n763 B.n761 10.6151
R1508 B.n764 B.n763 10.6151
R1509 B.n765 B.n764 10.6151
R1510 B.n766 B.n765 10.6151
R1511 B.n768 B.n766 10.6151
R1512 B.n769 B.n768 10.6151
R1513 B.n770 B.n769 10.6151
R1514 B.n771 B.n770 10.6151
R1515 B.n773 B.n771 10.6151
R1516 B.n774 B.n773 10.6151
R1517 B.n775 B.n774 10.6151
R1518 B.n776 B.n775 10.6151
R1519 B.n778 B.n776 10.6151
R1520 B.n779 B.n778 10.6151
R1521 B.n780 B.n779 10.6151
R1522 B.n781 B.n780 10.6151
R1523 B.n783 B.n781 10.6151
R1524 B.n784 B.n783 10.6151
R1525 B.n785 B.n784 10.6151
R1526 B.n786 B.n785 10.6151
R1527 B.n788 B.n786 10.6151
R1528 B.n789 B.n788 10.6151
R1529 B.n790 B.n789 10.6151
R1530 B.n791 B.n790 10.6151
R1531 B.n793 B.n791 10.6151
R1532 B.n794 B.n793 10.6151
R1533 B.n795 B.n794 10.6151
R1534 B.n796 B.n795 10.6151
R1535 B.n798 B.n796 10.6151
R1536 B.n799 B.n798 10.6151
R1537 B.n885 B.n1 10.6151
R1538 B.n885 B.n884 10.6151
R1539 B.n884 B.n883 10.6151
R1540 B.n883 B.n10 10.6151
R1541 B.n877 B.n10 10.6151
R1542 B.n877 B.n876 10.6151
R1543 B.n876 B.n875 10.6151
R1544 B.n875 B.n18 10.6151
R1545 B.n869 B.n18 10.6151
R1546 B.n869 B.n868 10.6151
R1547 B.n868 B.n867 10.6151
R1548 B.n867 B.n25 10.6151
R1549 B.n862 B.n25 10.6151
R1550 B.n862 B.n861 10.6151
R1551 B.n861 B.n860 10.6151
R1552 B.n860 B.n32 10.6151
R1553 B.n854 B.n32 10.6151
R1554 B.n854 B.n853 10.6151
R1555 B.n853 B.n852 10.6151
R1556 B.n852 B.n39 10.6151
R1557 B.n846 B.n39 10.6151
R1558 B.n846 B.n845 10.6151
R1559 B.n845 B.n844 10.6151
R1560 B.n844 B.n46 10.6151
R1561 B.n838 B.n46 10.6151
R1562 B.n838 B.n837 10.6151
R1563 B.n837 B.n836 10.6151
R1564 B.n836 B.n52 10.6151
R1565 B.n830 B.n52 10.6151
R1566 B.n830 B.n829 10.6151
R1567 B.n829 B.n828 10.6151
R1568 B.n828 B.n60 10.6151
R1569 B.n822 B.n60 10.6151
R1570 B.n822 B.n821 10.6151
R1571 B.n821 B.n820 10.6151
R1572 B.n820 B.n67 10.6151
R1573 B.n815 B.n67 10.6151
R1574 B.n815 B.n814 10.6151
R1575 B.n814 B.n813 10.6151
R1576 B.n813 B.n74 10.6151
R1577 B.n807 B.n74 10.6151
R1578 B.n807 B.n806 10.6151
R1579 B.n806 B.n805 10.6151
R1580 B.n133 B.n81 10.6151
R1581 B.n136 B.n133 10.6151
R1582 B.n137 B.n136 10.6151
R1583 B.n140 B.n137 10.6151
R1584 B.n141 B.n140 10.6151
R1585 B.n144 B.n141 10.6151
R1586 B.n145 B.n144 10.6151
R1587 B.n148 B.n145 10.6151
R1588 B.n149 B.n148 10.6151
R1589 B.n152 B.n149 10.6151
R1590 B.n153 B.n152 10.6151
R1591 B.n156 B.n153 10.6151
R1592 B.n157 B.n156 10.6151
R1593 B.n160 B.n157 10.6151
R1594 B.n161 B.n160 10.6151
R1595 B.n164 B.n161 10.6151
R1596 B.n165 B.n164 10.6151
R1597 B.n168 B.n165 10.6151
R1598 B.n169 B.n168 10.6151
R1599 B.n172 B.n169 10.6151
R1600 B.n173 B.n172 10.6151
R1601 B.n176 B.n173 10.6151
R1602 B.n177 B.n176 10.6151
R1603 B.n180 B.n177 10.6151
R1604 B.n181 B.n180 10.6151
R1605 B.n184 B.n181 10.6151
R1606 B.n185 B.n184 10.6151
R1607 B.n188 B.n185 10.6151
R1608 B.n189 B.n188 10.6151
R1609 B.n192 B.n189 10.6151
R1610 B.n193 B.n192 10.6151
R1611 B.n196 B.n193 10.6151
R1612 B.n197 B.n196 10.6151
R1613 B.n200 B.n197 10.6151
R1614 B.n201 B.n200 10.6151
R1615 B.n204 B.n201 10.6151
R1616 B.n205 B.n204 10.6151
R1617 B.n208 B.n205 10.6151
R1618 B.n213 B.n210 10.6151
R1619 B.n214 B.n213 10.6151
R1620 B.n217 B.n214 10.6151
R1621 B.n218 B.n217 10.6151
R1622 B.n221 B.n218 10.6151
R1623 B.n222 B.n221 10.6151
R1624 B.n225 B.n222 10.6151
R1625 B.n226 B.n225 10.6151
R1626 B.n230 B.n229 10.6151
R1627 B.n233 B.n230 10.6151
R1628 B.n234 B.n233 10.6151
R1629 B.n237 B.n234 10.6151
R1630 B.n238 B.n237 10.6151
R1631 B.n241 B.n238 10.6151
R1632 B.n242 B.n241 10.6151
R1633 B.n245 B.n242 10.6151
R1634 B.n246 B.n245 10.6151
R1635 B.n249 B.n246 10.6151
R1636 B.n250 B.n249 10.6151
R1637 B.n253 B.n250 10.6151
R1638 B.n254 B.n253 10.6151
R1639 B.n257 B.n254 10.6151
R1640 B.n258 B.n257 10.6151
R1641 B.n261 B.n258 10.6151
R1642 B.n262 B.n261 10.6151
R1643 B.n265 B.n262 10.6151
R1644 B.n266 B.n265 10.6151
R1645 B.n269 B.n266 10.6151
R1646 B.n270 B.n269 10.6151
R1647 B.n273 B.n270 10.6151
R1648 B.n274 B.n273 10.6151
R1649 B.n277 B.n274 10.6151
R1650 B.n278 B.n277 10.6151
R1651 B.n281 B.n278 10.6151
R1652 B.n282 B.n281 10.6151
R1653 B.n285 B.n282 10.6151
R1654 B.n286 B.n285 10.6151
R1655 B.n289 B.n286 10.6151
R1656 B.n290 B.n289 10.6151
R1657 B.n293 B.n290 10.6151
R1658 B.n294 B.n293 10.6151
R1659 B.n297 B.n294 10.6151
R1660 B.n298 B.n297 10.6151
R1661 B.n301 B.n298 10.6151
R1662 B.n302 B.n301 10.6151
R1663 B.n800 B.n302 10.6151
R1664 B.n893 B.n0 8.11757
R1665 B.n893 B.n1 8.11757
R1666 B.n510 B.n509 6.5566
R1667 B.n529 B.n528 6.5566
R1668 B.n210 B.n209 6.5566
R1669 B.n226 B.n130 6.5566
R1670 B.n509 B.n508 4.05904
R1671 B.n528 B.n407 4.05904
R1672 B.n209 B.n208 4.05904
R1673 B.n229 B.n130 4.05904
R1674 VN.n43 VN.n23 161.3
R1675 VN.n42 VN.n41 161.3
R1676 VN.n40 VN.n24 161.3
R1677 VN.n39 VN.n38 161.3
R1678 VN.n37 VN.n25 161.3
R1679 VN.n35 VN.n34 161.3
R1680 VN.n33 VN.n26 161.3
R1681 VN.n32 VN.n31 161.3
R1682 VN.n30 VN.n27 161.3
R1683 VN.n20 VN.n0 161.3
R1684 VN.n19 VN.n18 161.3
R1685 VN.n17 VN.n1 161.3
R1686 VN.n16 VN.n15 161.3
R1687 VN.n14 VN.n2 161.3
R1688 VN.n12 VN.n11 161.3
R1689 VN.n10 VN.n3 161.3
R1690 VN.n9 VN.n8 161.3
R1691 VN.n7 VN.n4 161.3
R1692 VN.n5 VN.t3 157.587
R1693 VN.n28 VN.t6 157.587
R1694 VN.n6 VN.t7 123.091
R1695 VN.n13 VN.t2 123.091
R1696 VN.n21 VN.t5 123.091
R1697 VN.n29 VN.t0 123.091
R1698 VN.n36 VN.t4 123.091
R1699 VN.n44 VN.t1 123.091
R1700 VN.n22 VN.n21 88.4915
R1701 VN.n45 VN.n44 88.4915
R1702 VN.n8 VN.n3 56.5193
R1703 VN.n19 VN.n1 56.5193
R1704 VN.n31 VN.n26 56.5193
R1705 VN.n42 VN.n24 56.5193
R1706 VN VN.n45 48.3088
R1707 VN.n6 VN.n5 47.0153
R1708 VN.n29 VN.n28 47.0153
R1709 VN.n8 VN.n7 24.4675
R1710 VN.n12 VN.n3 24.4675
R1711 VN.n15 VN.n14 24.4675
R1712 VN.n15 VN.n1 24.4675
R1713 VN.n20 VN.n19 24.4675
R1714 VN.n31 VN.n30 24.4675
R1715 VN.n38 VN.n24 24.4675
R1716 VN.n38 VN.n37 24.4675
R1717 VN.n35 VN.n26 24.4675
R1718 VN.n43 VN.n42 24.4675
R1719 VN.n7 VN.n6 23.7335
R1720 VN.n13 VN.n12 23.7335
R1721 VN.n30 VN.n29 23.7335
R1722 VN.n36 VN.n35 23.7335
R1723 VN.n21 VN.n20 22.2655
R1724 VN.n44 VN.n43 22.2655
R1725 VN.n28 VN.n27 8.75906
R1726 VN.n5 VN.n4 8.75906
R1727 VN.n14 VN.n13 0.73451
R1728 VN.n37 VN.n36 0.73451
R1729 VN.n45 VN.n23 0.278367
R1730 VN.n22 VN.n0 0.278367
R1731 VN.n41 VN.n23 0.189894
R1732 VN.n41 VN.n40 0.189894
R1733 VN.n40 VN.n39 0.189894
R1734 VN.n39 VN.n25 0.189894
R1735 VN.n34 VN.n25 0.189894
R1736 VN.n34 VN.n33 0.189894
R1737 VN.n33 VN.n32 0.189894
R1738 VN.n32 VN.n27 0.189894
R1739 VN.n9 VN.n4 0.189894
R1740 VN.n10 VN.n9 0.189894
R1741 VN.n11 VN.n10 0.189894
R1742 VN.n11 VN.n2 0.189894
R1743 VN.n16 VN.n2 0.189894
R1744 VN.n17 VN.n16 0.189894
R1745 VN.n18 VN.n17 0.189894
R1746 VN.n18 VN.n0 0.189894
R1747 VN VN.n22 0.153454
R1748 VDD2.n2 VDD2.n1 61.0849
R1749 VDD2.n2 VDD2.n0 61.0849
R1750 VDD2 VDD2.n5 61.0821
R1751 VDD2.n4 VDD2.n3 60.0758
R1752 VDD2.n4 VDD2.n2 42.7196
R1753 VDD2.n5 VDD2.t7 1.81203
R1754 VDD2.n5 VDD2.t1 1.81203
R1755 VDD2.n3 VDD2.t6 1.81203
R1756 VDD2.n3 VDD2.t3 1.81203
R1757 VDD2.n1 VDD2.t5 1.81203
R1758 VDD2.n1 VDD2.t2 1.81203
R1759 VDD2.n0 VDD2.t4 1.81203
R1760 VDD2.n0 VDD2.t0 1.81203
R1761 VDD2 VDD2.n4 1.12334
C0 VTAIL VDD2 7.71869f
C1 VTAIL VP 7.93637f
C2 VDD2 VN 7.627501f
C3 VP VN 6.89966f
C4 VTAIL VDD1 7.66736f
C5 VDD2 VP 0.470812f
C6 VDD1 VN 0.150987f
C7 VDD1 VDD2 1.53864f
C8 VDD1 VP 7.94616f
C9 VTAIL VN 7.922259f
C10 VDD2 B 4.824872f
C11 VDD1 B 5.214273f
C12 VTAIL B 9.5304f
C13 VN B 13.660871f
C14 VP B 12.210309f
C15 VDD2.t4 B 0.210633f
C16 VDD2.t0 B 0.210633f
C17 VDD2.n0 B 1.87117f
C18 VDD2.t5 B 0.210633f
C19 VDD2.t2 B 0.210633f
C20 VDD2.n1 B 1.87117f
C21 VDD2.n2 B 2.87561f
C22 VDD2.t6 B 0.210633f
C23 VDD2.t3 B 0.210633f
C24 VDD2.n3 B 1.86358f
C25 VDD2.n4 B 2.64362f
C26 VDD2.t7 B 0.210633f
C27 VDD2.t1 B 0.210633f
C28 VDD2.n5 B 1.87113f
C29 VN.n0 B 0.033258f
C30 VN.t5 B 1.60316f
C31 VN.n1 B 0.034717f
C32 VN.n2 B 0.025226f
C33 VN.t2 B 1.60316f
C34 VN.n3 B 0.036826f
C35 VN.n4 B 0.212932f
C36 VN.t7 B 1.60316f
C37 VN.t3 B 1.75965f
C38 VN.n5 B 0.628076f
C39 VN.n6 B 0.650204f
C40 VN.n7 B 0.046318f
C41 VN.n8 B 0.036826f
C42 VN.n9 B 0.025226f
C43 VN.n10 B 0.025226f
C44 VN.n11 B 0.025226f
C45 VN.n12 B 0.046318f
C46 VN.n13 B 0.574404f
C47 VN.n14 B 0.024499f
C48 VN.n15 B 0.047015f
C49 VN.n16 B 0.025226f
C50 VN.n17 B 0.025226f
C51 VN.n18 B 0.025226f
C52 VN.n19 B 0.038935f
C53 VN.n20 B 0.044925f
C54 VN.n21 B 0.661077f
C55 VN.n22 B 0.029136f
C56 VN.n23 B 0.033258f
C57 VN.t1 B 1.60316f
C58 VN.n24 B 0.034717f
C59 VN.n25 B 0.025226f
C60 VN.t4 B 1.60316f
C61 VN.n26 B 0.036826f
C62 VN.n27 B 0.212932f
C63 VN.t0 B 1.60316f
C64 VN.t6 B 1.75965f
C65 VN.n28 B 0.628076f
C66 VN.n29 B 0.650204f
C67 VN.n30 B 0.046318f
C68 VN.n31 B 0.036826f
C69 VN.n32 B 0.025226f
C70 VN.n33 B 0.025226f
C71 VN.n34 B 0.025226f
C72 VN.n35 B 0.046318f
C73 VN.n36 B 0.574404f
C74 VN.n37 B 0.024499f
C75 VN.n38 B 0.047015f
C76 VN.n39 B 0.025226f
C77 VN.n40 B 0.025226f
C78 VN.n41 B 0.025226f
C79 VN.n42 B 0.038935f
C80 VN.n43 B 0.044925f
C81 VN.n44 B 0.661077f
C82 VN.n45 B 1.32444f
C83 VTAIL.t1 B 0.170878f
C84 VTAIL.t6 B 0.170878f
C85 VTAIL.n0 B 1.45009f
C86 VTAIL.n1 B 0.338734f
C87 VTAIL.t5 B 1.84618f
C88 VTAIL.n2 B 0.434913f
C89 VTAIL.t10 B 1.84618f
C90 VTAIL.n3 B 0.434913f
C91 VTAIL.t13 B 0.170878f
C92 VTAIL.t15 B 0.170878f
C93 VTAIL.n4 B 1.45009f
C94 VTAIL.n5 B 0.470764f
C95 VTAIL.t8 B 1.84618f
C96 VTAIL.n6 B 1.4101f
C97 VTAIL.t7 B 1.8462f
C98 VTAIL.n7 B 1.41009f
C99 VTAIL.t0 B 0.170878f
C100 VTAIL.t2 B 0.170878f
C101 VTAIL.n8 B 1.4501f
C102 VTAIL.n9 B 0.470759f
C103 VTAIL.t3 B 1.8462f
C104 VTAIL.n10 B 0.4349f
C105 VTAIL.t12 B 1.8462f
C106 VTAIL.n11 B 0.4349f
C107 VTAIL.t9 B 0.170878f
C108 VTAIL.t14 B 0.170878f
C109 VTAIL.n12 B 1.4501f
C110 VTAIL.n13 B 0.470759f
C111 VTAIL.t11 B 1.84618f
C112 VTAIL.n14 B 1.4101f
C113 VTAIL.t4 B 1.84618f
C114 VTAIL.n15 B 1.40639f
C115 VDD1.t6 B 0.213506f
C116 VDD1.t5 B 0.213506f
C117 VDD1.n0 B 1.8977f
C118 VDD1.t4 B 0.213506f
C119 VDD1.t0 B 0.213506f
C120 VDD1.n1 B 1.89669f
C121 VDD1.t2 B 0.213506f
C122 VDD1.t7 B 0.213506f
C123 VDD1.n2 B 1.89669f
C124 VDD1.n3 B 2.96663f
C125 VDD1.t1 B 0.213506f
C126 VDD1.t3 B 0.213506f
C127 VDD1.n4 B 1.88899f
C128 VDD1.n5 B 2.70992f
C129 VP.n0 B 0.033757f
C130 VP.t5 B 1.6272f
C131 VP.n1 B 0.035238f
C132 VP.n2 B 0.025605f
C133 VP.t0 B 1.6272f
C134 VP.n3 B 0.037378f
C135 VP.n4 B 0.025605f
C136 VP.t2 B 1.6272f
C137 VP.n5 B 0.04772f
C138 VP.n6 B 0.025605f
C139 VP.t7 B 1.6272f
C140 VP.n7 B 0.670993f
C141 VP.n8 B 0.033757f
C142 VP.t4 B 1.6272f
C143 VP.n9 B 0.035238f
C144 VP.n10 B 0.025605f
C145 VP.t1 B 1.6272f
C146 VP.n11 B 0.037378f
C147 VP.n12 B 0.216126f
C148 VP.t6 B 1.6272f
C149 VP.t3 B 1.78604f
C150 VP.n13 B 0.637497f
C151 VP.n14 B 0.659957f
C152 VP.n15 B 0.047013f
C153 VP.n16 B 0.037378f
C154 VP.n17 B 0.025605f
C155 VP.n18 B 0.025605f
C156 VP.n19 B 0.025605f
C157 VP.n20 B 0.047013f
C158 VP.n21 B 0.58302f
C159 VP.n22 B 0.024866f
C160 VP.n23 B 0.04772f
C161 VP.n24 B 0.025605f
C162 VP.n25 B 0.025605f
C163 VP.n26 B 0.025605f
C164 VP.n27 B 0.039519f
C165 VP.n28 B 0.045599f
C166 VP.n29 B 0.670993f
C167 VP.n30 B 1.33046f
C168 VP.n31 B 1.34963f
C169 VP.n32 B 0.033757f
C170 VP.n33 B 0.045599f
C171 VP.n34 B 0.039519f
C172 VP.n35 B 0.035238f
C173 VP.n36 B 0.025605f
C174 VP.n37 B 0.025605f
C175 VP.n38 B 0.025605f
C176 VP.n39 B 0.024866f
C177 VP.n40 B 0.58302f
C178 VP.n41 B 0.047013f
C179 VP.n42 B 0.037378f
C180 VP.n43 B 0.025605f
C181 VP.n44 B 0.025605f
C182 VP.n45 B 0.025605f
C183 VP.n46 B 0.047013f
C184 VP.n47 B 0.58302f
C185 VP.n48 B 0.024866f
C186 VP.n49 B 0.04772f
C187 VP.n50 B 0.025605f
C188 VP.n51 B 0.025605f
C189 VP.n52 B 0.025605f
C190 VP.n53 B 0.039519f
C191 VP.n54 B 0.045599f
C192 VP.n55 B 0.670993f
C193 VP.n56 B 0.029573f
.ends

