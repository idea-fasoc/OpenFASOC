** sch_path: /home/chandru/Tools/OpenFASOC/generators/lc-dco/xschem_rundir/swcap_3M2C_scaled.sch
.subckt swcap_3M2C_scaled outn outp sw<7> sw<6> sw<5> sw<4> sw<3> sw<2> sw<1> sw<0> GND
*.PININFO outn:O outp:O sw[7:0]:I GND:B
XC2<7> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<6> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<5> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<4> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<3> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<2> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<1> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2<0> net2 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM6 net1 sw<0> net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 GND sw<0> net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 GND sw<0> net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1<7> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<6> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<5> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<4> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<3> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<2> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<1> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC1<0> outp net1 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<15> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<14> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<13> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<12> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<11> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<10> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<9> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<8> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<7> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<6> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<5> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<4> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<3> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<2> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<1> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC4<0> net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM3 net3 sw<1> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 GND sw<1> net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 GND sw<1> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC3<15> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<14> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<13> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<12> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<11> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<10> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<9> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<8> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<7> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<6> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<5> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<4> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<3> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<2> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<1> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3<0> outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<31> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<30> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<29> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<28> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<27> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<26> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<25> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<24> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<23> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<22> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<21> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<20> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<19> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<18> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<17> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<16> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<15> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<14> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<13> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<12> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<11> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<10> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<9> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<8> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<7> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<6> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<5> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<4> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<3> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<2> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<1> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC6<0> net6 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM7 net5 sw<2> net6 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 GND sw<2> net5 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 GND sw<2> net6 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC5<31> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<30> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<29> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<28> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<27> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<26> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<25> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<24> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<23> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<22> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<21> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<20> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<19> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<18> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<17> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<16> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<15> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<14> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<13> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<12> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<11> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<10> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<9> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<8> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<7> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<6> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<5> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<4> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<3> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<2> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<1> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC5<0> outp net5 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<63> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<62> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<61> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<60> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<59> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<58> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<57> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<56> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<55> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<54> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<53> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<52> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<51> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<50> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<49> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<48> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<47> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<46> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<45> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<44> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<43> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<42> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<41> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<40> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<39> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<38> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<37> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<36> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<35> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<34> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<33> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<32> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<31> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<30> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<29> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<28> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<27> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<26> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<25> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<24> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<23> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<22> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<21> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<20> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<19> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<18> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<17> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<16> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<15> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<14> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<13> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<12> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<11> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<10> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<9> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<8> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<7> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<6> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<5> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<4> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<3> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<2> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<1> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC8<0> net8 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM10 net7 sw<3> net8 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 GND sw<3> net7 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 GND sw<3> net8 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC7<63> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<62> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<61> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<60> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<59> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<58> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<57> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<56> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<55> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<54> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<53> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<52> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<51> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<50> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<49> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<48> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<47> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<46> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<45> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<44> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<43> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<42> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<41> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<40> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<39> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<38> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<37> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<36> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<35> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<34> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<33> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<32> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<31> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<30> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<29> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<28> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<27> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<26> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<25> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<24> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<23> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<22> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<21> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<20> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<19> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<18> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<17> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<16> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<15> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<14> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<13> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<12> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<11> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<10> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<9> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<8> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<7> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<6> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<5> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<4> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<3> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<2> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<1> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC7<0> outp net7 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<127> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<126> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<125> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<124> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<123> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<122> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<121> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<120> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<119> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<118> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<117> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<116> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<115> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<114> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<113> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<112> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<111> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<110> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<109> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<108> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<107> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<106> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<105> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<104> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<103> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<102> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<101> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<100> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<99> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<98> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<97> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<96> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<95> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<94> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<93> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<92> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<91> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<90> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<89> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<88> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<87> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<86> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<85> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<84> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<83> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<82> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<81> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<80> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<79> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<78> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<77> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<76> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<75> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<74> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<73> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<72> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<71> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<70> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<69> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<68> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<67> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<66> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<65> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<64> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<63> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<62> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<61> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<60> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<59> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<58> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<57> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<56> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<55> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<54> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<53> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<52> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<51> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<50> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<49> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<48> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<47> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<46> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<45> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<44> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<43> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<42> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<41> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<40> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<39> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<38> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<37> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<36> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<35> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<34> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<33> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<32> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<31> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<30> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<29> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<28> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<27> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<26> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<25> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<24> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<23> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<22> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<21> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<20> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<19> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<18> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<17> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<16> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<15> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<14> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<13> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<12> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<11> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<10> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<9> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<8> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<7> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<6> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<5> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<4> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<3> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<2> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<1> net10<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC10<0> net10<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM13<1> net9<1> sw<4> net10<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13<0> net9<0> sw<4> net10<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14<2> GND sw<4> net9<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14<1> GND sw<4> net9<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14<0> GND sw<4> net9<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15<2> GND sw<4> net10<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15<1> GND sw<4> net10<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15<0> GND sw<4> net10<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC9<127> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<126> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<125> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<124> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<123> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<122> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<121> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<120> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<119> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<118> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<117> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<116> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<115> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<114> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<113> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<112> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<111> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<110> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<109> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<108> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<107> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<106> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<105> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<104> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<103> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<102> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<101> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<100> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<99> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<98> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<97> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<96> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<95> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<94> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<93> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<92> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<91> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<90> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<89> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<88> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<87> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<86> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<85> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<84> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<83> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<82> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<81> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<80> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<79> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<78> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<77> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<76> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<75> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<74> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<73> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<72> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<71> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<70> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<69> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<68> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<67> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<66> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<65> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<64> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<63> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<62> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<61> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<60> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<59> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<58> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<57> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<56> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<55> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<54> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<53> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<52> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<51> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<50> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<49> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<48> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<47> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<46> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<45> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<44> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<43> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<42> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<41> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<40> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<39> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<38> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<37> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<36> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<35> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<34> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<33> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<32> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<31> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<30> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<29> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<28> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<27> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<26> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<25> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<24> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<23> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<22> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<21> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<20> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<19> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<18> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<17> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<16> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<15> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<14> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<13> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<12> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<11> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<10> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<9> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<8> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<7> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<6> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<5> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<4> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<3> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<2> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<1> outp net9<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC9<0> outp net9<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<255> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<254> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<253> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<252> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<251> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<250> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<249> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<248> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<247> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<246> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<245> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<244> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<243> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<242> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<241> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<240> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<239> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<238> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<237> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<236> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<235> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<234> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<233> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<232> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<231> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<230> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<229> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<228> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<227> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<226> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<225> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<224> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<223> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<222> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<221> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<220> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<219> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<218> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<217> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<216> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<215> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<214> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<213> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<212> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<211> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<210> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<209> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<208> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<207> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<206> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<205> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<204> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<203> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<202> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<201> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<200> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<199> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<198> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<197> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<196> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<195> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<194> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<193> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<192> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<191> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<190> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<189> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<188> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<187> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<186> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<185> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<184> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<183> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<182> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<181> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<180> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<179> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<178> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<177> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<176> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<175> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<174> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<173> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<172> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<171> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<170> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<169> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<168> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<167> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<166> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<165> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<164> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<163> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<162> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<161> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<160> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<159> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<158> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<157> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<156> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<155> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<154> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<153> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<152> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<151> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<150> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<149> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<148> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<147> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<146> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<145> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<144> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<143> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<142> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<141> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<140> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<139> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<138> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<137> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<136> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<135> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<134> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<133> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<132> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<131> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<130> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<129> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<128> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<127> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<126> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<125> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<124> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<123> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<122> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<121> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<120> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<119> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<118> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<117> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<116> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<115> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<114> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<113> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<112> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<111> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<110> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<109> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<108> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<107> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<106> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<105> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<104> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<103> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<102> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<101> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<100> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<99> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<98> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<97> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<96> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<95> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<94> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<93> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<92> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<91> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<90> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<89> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<88> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<87> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<86> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<85> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<84> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<83> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<82> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<81> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<80> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<79> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<78> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<77> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<76> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<75> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<74> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<73> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<72> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<71> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<70> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<69> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<68> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<67> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<66> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<65> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<64> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<63> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<62> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<61> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<60> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<59> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<58> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<57> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<56> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<55> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<54> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<53> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<52> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<51> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<50> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<49> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<48> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<47> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<46> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<45> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<44> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<43> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<42> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<41> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<40> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<39> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<38> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<37> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<36> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<35> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<34> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<33> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<32> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<31> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<30> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<29> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<28> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<27> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<26> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<25> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<24> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<23> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<22> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<21> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<20> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<19> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<18> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<17> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<16> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<15> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<14> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<13> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<12> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<11> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<10> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<9> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<8> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<7> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<6> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<5> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<4> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<3> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<2> net12<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<1> net12<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC12<0> net12<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM16<2> net11<2> sw<5> net12<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16<1> net11<1> sw<5> net12<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16<0> net11<0> sw<5> net12<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17<2> GND sw<5> net11<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17<1> GND sw<5> net11<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17<0> GND sw<5> net11<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18<2> GND sw<5> net12<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18<1> GND sw<5> net12<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18<0> GND sw<5> net12<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC11<255> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<254> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<253> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<252> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<251> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<250> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<249> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<248> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<247> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<246> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<245> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<244> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<243> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<242> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<241> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<240> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<239> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<238> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<237> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<236> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<235> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<234> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<233> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<232> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<231> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<230> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<229> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<228> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<227> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<226> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<225> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<224> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<223> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<222> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<221> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<220> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<219> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<218> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<217> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<216> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<215> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<214> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<213> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<212> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<211> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<210> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<209> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<208> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<207> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<206> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<205> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<204> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<203> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<202> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<201> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<200> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<199> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<198> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<197> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<196> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<195> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<194> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<193> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<192> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<191> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<190> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<189> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<188> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<187> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<186> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<185> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<184> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<183> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<182> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<181> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<180> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<179> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<178> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<177> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<176> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<175> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<174> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<173> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<172> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<171> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<170> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<169> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<168> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<167> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<166> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<165> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<164> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<163> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<162> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<161> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<160> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<159> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<158> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<157> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<156> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<155> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<154> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<153> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<152> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<151> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<150> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<149> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<148> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<147> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<146> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<145> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<144> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<143> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<142> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<141> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<140> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<139> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<138> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<137> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<136> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<135> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<134> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<133> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<132> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<131> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<130> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<129> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<128> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<127> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<126> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<125> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<124> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<123> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<122> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<121> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<120> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<119> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<118> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<117> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<116> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<115> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<114> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<113> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<112> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<111> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<110> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<109> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<108> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<107> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<106> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<105> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<104> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<103> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<102> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<101> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<100> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<99> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<98> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<97> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<96> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<95> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<94> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<93> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<92> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<91> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<90> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<89> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<88> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<87> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<86> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<85> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<84> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<83> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<82> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<81> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<80> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<79> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<78> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<77> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<76> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<75> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<74> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<73> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<72> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<71> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<70> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<69> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<68> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<67> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<66> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<65> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<64> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<63> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<62> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<61> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<60> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<59> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<58> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<57> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<56> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<55> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<54> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<53> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<52> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<51> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<50> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<49> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<48> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<47> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<46> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<45> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<44> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<43> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<42> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<41> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<40> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<39> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<38> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<37> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<36> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<35> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<34> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<33> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<32> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<31> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<30> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<29> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<28> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<27> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<26> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<25> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<24> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<23> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<22> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<21> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<20> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<19> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<18> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<17> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<16> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<15> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<14> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<13> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<12> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<11> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<10> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<9> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<8> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<7> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<6> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<5> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<4> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<3> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<2> outp net11<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<1> outp net11<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC11<0> outp net11<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<511> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<510> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<509> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<508> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<507> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<506> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<505> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<504> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<503> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<502> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<501> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<500> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<499> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<498> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<497> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<496> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<495> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<494> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<493> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<492> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<491> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<490> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<489> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<488> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<487> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<486> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<485> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<484> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<483> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<482> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<481> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<480> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<479> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<478> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<477> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<476> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<475> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<474> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<473> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<472> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<471> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<470> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<469> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<468> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<467> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<466> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<465> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<464> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<463> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<462> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<461> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<460> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<459> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<458> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<457> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<456> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<455> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<454> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<453> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<452> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<451> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<450> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<449> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<448> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<447> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<446> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<445> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<444> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<443> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<442> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<441> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<440> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<439> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<438> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<437> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<436> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<435> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<434> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<433> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<432> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<431> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<430> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<429> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<428> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<427> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<426> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<425> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<424> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<423> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<422> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<421> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<420> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<419> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<418> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<417> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<416> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<415> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<414> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<413> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<412> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<411> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<410> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<409> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<408> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<407> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<406> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<405> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<404> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<403> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<402> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<401> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<400> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<399> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<398> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<397> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<396> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<395> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<394> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<393> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<392> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<391> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<390> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<389> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<388> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<387> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<386> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<385> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<384> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<383> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<382> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<381> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<380> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<379> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<378> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<377> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<376> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<375> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<374> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<373> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<372> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<371> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<370> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<369> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<368> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<367> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<366> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<365> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<364> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<363> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<362> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<361> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<360> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<359> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<358> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<357> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<356> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<355> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<354> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<353> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<352> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<351> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<350> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<349> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<348> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<347> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<346> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<345> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<344> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<343> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<342> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<341> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<340> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<339> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<338> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<337> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<336> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<335> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<334> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<333> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<332> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<331> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<330> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<329> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<328> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<327> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<326> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<325> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<324> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<323> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<322> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<321> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<320> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<319> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<318> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<317> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<316> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<315> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<314> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<313> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<312> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<311> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<310> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<309> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<308> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<307> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<306> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<305> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<304> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<303> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<302> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<301> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<300> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<299> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<298> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<297> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<296> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<295> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<294> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<293> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<292> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<291> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<290> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<289> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<288> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<287> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<286> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<285> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<284> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<283> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<282> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<281> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<280> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<279> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<278> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<277> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<276> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<275> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<274> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<273> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<272> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<271> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<270> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<269> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<268> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<267> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<266> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<265> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<264> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<263> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<262> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<261> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<260> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<259> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<258> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<257> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<256> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<255> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<254> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<253> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<252> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<251> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<250> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<249> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<248> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<247> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<246> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<245> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<244> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<243> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<242> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<241> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<240> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<239> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<238> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<237> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<236> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<235> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<234> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<233> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<232> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<231> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<230> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<229> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<228> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<227> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<226> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<225> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<224> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<223> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<222> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<221> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<220> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<219> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<218> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<217> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<216> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<215> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<214> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<213> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<212> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<211> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<210> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<209> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<208> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<207> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<206> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<205> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<204> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<203> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<202> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<201> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<200> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<199> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<198> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<197> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<196> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<195> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<194> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<193> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<192> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<191> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<190> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<189> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<188> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<187> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<186> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<185> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<184> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<183> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<182> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<181> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<180> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<179> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<178> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<177> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<176> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<175> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<174> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<173> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<172> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<171> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<170> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<169> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<168> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<167> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<166> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<165> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<164> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<163> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<162> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<161> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<160> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<159> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<158> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<157> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<156> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<155> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<154> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<153> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<152> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<151> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<150> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<149> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<148> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<147> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<146> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<145> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<144> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<143> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<142> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<141> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<140> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<139> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<138> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<137> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<136> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<135> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<134> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<133> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<132> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<131> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<130> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<129> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<128> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<127> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<126> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<125> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<124> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<123> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<122> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<121> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<120> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<119> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<118> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<117> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<116> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<115> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<114> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<113> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<112> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<111> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<110> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<109> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<108> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<107> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<106> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<105> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<104> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<103> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<102> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<101> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<100> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<99> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<98> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<97> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<96> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<95> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<94> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<93> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<92> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<91> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<90> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<89> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<88> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<87> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<86> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<85> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<84> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<83> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<82> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<81> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<80> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<79> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<78> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<77> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<76> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<75> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<74> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<73> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<72> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<71> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<70> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<69> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<68> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<67> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<66> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<65> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<64> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<63> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<62> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<61> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<60> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<59> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<58> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<57> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<56> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<55> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<54> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<53> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<52> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<51> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<50> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<49> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<48> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<47> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<46> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<45> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<44> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<43> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<42> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<41> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<40> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<39> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<38> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<37> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<36> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<35> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<34> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<33> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<32> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<31> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<30> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<29> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<28> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<27> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<26> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<25> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<24> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<23> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<22> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<21> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<20> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<19> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<18> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<17> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<16> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<15> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<14> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<13> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<12> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<11> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<10> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<9> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<8> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<7> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<6> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<5> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<4> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<3> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<2> net14<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<1> net14<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC14<0> net14<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM19<2> net13<2> sw<6> net14<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM19<1> net13<1> sw<6> net14<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM19<0> net13<0> sw<6> net14<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM20<2> GND sw<6> net13<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20<1> GND sw<6> net13<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20<0> GND sw<6> net13<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21<2> GND sw<6> net14<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21<1> GND sw<6> net14<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21<0> GND sw<6> net14<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC13<511> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<510> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<509> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<508> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<507> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<506> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<505> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<504> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<503> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<502> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<501> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<500> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<499> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<498> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<497> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<496> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<495> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<494> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<493> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<492> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<491> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<490> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<489> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<488> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<487> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<486> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<485> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<484> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<483> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<482> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<481> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<480> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<479> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<478> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<477> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<476> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<475> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<474> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<473> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<472> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<471> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<470> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<469> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<468> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<467> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<466> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<465> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<464> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<463> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<462> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<461> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<460> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<459> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<458> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<457> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<456> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<455> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<454> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<453> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<452> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<451> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<450> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<449> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<448> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<447> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<446> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<445> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<444> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<443> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<442> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<441> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<440> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<439> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<438> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<437> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<436> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<435> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<434> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<433> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<432> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<431> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<430> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<429> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<428> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<427> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<426> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<425> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<424> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<423> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<422> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<421> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<420> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<419> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<418> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<417> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<416> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<415> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<414> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<413> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<412> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<411> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<410> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<409> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<408> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<407> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<406> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<405> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<404> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<403> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<402> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<401> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<400> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<399> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<398> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<397> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<396> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<395> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<394> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<393> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<392> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<391> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<390> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<389> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<388> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<387> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<386> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<385> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<384> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<383> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<382> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<381> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<380> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<379> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<378> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<377> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<376> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<375> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<374> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<373> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<372> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<371> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<370> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<369> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<368> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<367> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<366> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<365> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<364> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<363> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<362> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<361> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<360> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<359> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<358> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<357> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<356> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<355> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<354> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<353> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<352> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<351> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<350> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<349> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<348> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<347> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<346> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<345> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<344> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<343> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<342> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<341> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<340> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<339> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<338> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<337> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<336> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<335> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<334> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<333> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<332> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<331> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<330> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<329> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<328> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<327> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<326> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<325> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<324> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<323> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<322> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<321> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<320> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<319> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<318> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<317> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<316> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<315> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<314> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<313> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<312> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<311> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<310> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<309> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<308> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<307> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<306> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<305> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<304> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<303> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<302> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<301> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<300> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<299> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<298> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<297> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<296> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<295> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<294> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<293> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<292> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<291> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<290> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<289> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<288> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<287> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<286> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<285> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<284> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<283> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<282> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<281> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<280> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<279> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<278> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<277> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<276> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<275> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<274> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<273> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<272> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<271> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<270> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<269> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<268> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<267> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<266> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<265> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<264> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<263> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<262> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<261> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<260> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<259> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<258> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<257> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<256> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<255> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<254> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<253> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<252> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<251> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<250> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<249> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<248> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<247> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<246> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<245> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<244> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<243> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<242> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<241> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<240> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<239> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<238> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<237> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<236> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<235> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<234> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<233> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<232> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<231> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<230> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<229> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<228> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<227> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<226> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<225> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<224> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<223> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<222> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<221> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<220> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<219> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<218> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<217> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<216> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<215> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<214> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<213> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<212> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<211> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<210> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<209> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<208> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<207> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<206> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<205> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<204> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<203> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<202> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<201> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<200> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<199> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<198> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<197> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<196> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<195> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<194> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<193> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<192> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<191> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<190> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<189> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<188> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<187> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<186> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<185> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<184> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<183> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<182> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<181> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<180> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<179> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<178> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<177> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<176> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<175> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<174> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<173> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<172> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<171> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<170> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<169> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<168> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<167> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<166> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<165> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<164> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<163> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<162> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<161> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<160> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<159> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<158> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<157> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<156> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<155> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<154> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<153> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<152> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<151> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<150> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<149> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<148> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<147> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<146> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<145> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<144> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<143> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<142> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<141> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<140> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<139> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<138> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<137> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<136> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<135> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<134> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<133> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<132> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<131> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<130> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<129> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<128> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<127> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<126> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<125> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<124> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<123> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<122> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<121> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<120> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<119> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<118> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<117> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<116> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<115> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<114> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<113> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<112> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<111> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<110> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<109> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<108> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<107> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<106> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<105> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<104> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<103> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<102> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<101> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<100> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<99> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<98> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<97> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<96> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<95> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<94> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<93> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<92> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<91> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<90> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<89> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<88> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<87> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<86> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<85> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<84> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<83> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<82> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<81> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<80> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<79> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<78> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<77> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<76> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<75> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<74> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<73> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<72> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<71> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<70> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<69> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<68> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<67> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<66> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<65> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<64> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<63> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<62> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<61> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<60> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<59> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<58> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<57> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<56> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<55> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<54> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<53> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<52> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<51> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<50> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<49> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<48> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<47> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<46> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<45> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<44> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<43> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<42> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<41> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<40> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<39> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<38> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<37> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<36> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<35> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<34> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<33> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<32> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<31> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<30> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<29> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<28> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<27> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<26> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<25> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<24> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<23> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<22> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<21> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<20> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<19> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<18> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<17> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<16> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<15> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<14> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<13> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<12> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<11> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<10> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<9> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<8> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<7> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<6> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<5> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<4> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<3> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<2> outp net13<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<1> outp net13<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC13<0> outp net13<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1023> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1022> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1021> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1020> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1019> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1018> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1017> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1016> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1015> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1014> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1013> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1012> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1011> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1010> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1009> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1008> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1007> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1006> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1005> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1004> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1003> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1002> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1001> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1000> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<999> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<998> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<997> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<996> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<995> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<994> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<993> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<992> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<991> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<990> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<989> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<988> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<987> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<986> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<985> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<984> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<983> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<982> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<981> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<980> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<979> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<978> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<977> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<976> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<975> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<974> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<973> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<972> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<971> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<970> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<969> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<968> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<967> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<966> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<965> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<964> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<963> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<962> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<961> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<960> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<959> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<958> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<957> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<956> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<955> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<954> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<953> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<952> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<951> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<950> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<949> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<948> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<947> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<946> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<945> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<944> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<943> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<942> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<941> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<940> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<939> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<938> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<937> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<936> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<935> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<934> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<933> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<932> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<931> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<930> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<929> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<928> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<927> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<926> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<925> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<924> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<923> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<922> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<921> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<920> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<919> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<918> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<917> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<916> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<915> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<914> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<913> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<912> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<911> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<910> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<909> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<908> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<907> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<906> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<905> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<904> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<903> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<902> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<901> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<900> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<899> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<898> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<897> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<896> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<895> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<894> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<893> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<892> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<891> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<890> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<889> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<888> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<887> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<886> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<885> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<884> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<883> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<882> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<881> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<880> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<879> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<878> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<877> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<876> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<875> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<874> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<873> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<872> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<871> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<870> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<869> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<868> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<867> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<866> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<865> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<864> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<863> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<862> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<861> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<860> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<859> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<858> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<857> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<856> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<855> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<854> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<853> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<852> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<851> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<850> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<849> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<848> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<847> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<846> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<845> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<844> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<843> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<842> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<841> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<840> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<839> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<838> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<837> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<836> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<835> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<834> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<833> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<832> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<831> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<830> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<829> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<828> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<827> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<826> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<825> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<824> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<823> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<822> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<821> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<820> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<819> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<818> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<817> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<816> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<815> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<814> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<813> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<812> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<811> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<810> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<809> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<808> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<807> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<806> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<805> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<804> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<803> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<802> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<801> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<800> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<799> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<798> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<797> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<796> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<795> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<794> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<793> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<792> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<791> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<790> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<789> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<788> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<787> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<786> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<785> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<784> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<783> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<782> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<781> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<780> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<779> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<778> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<777> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<776> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<775> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<774> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<773> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<772> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<771> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<770> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<769> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<768> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<767> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<766> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<765> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<764> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<763> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<762> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<761> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<760> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<759> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<758> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<757> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<756> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<755> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<754> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<753> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<752> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<751> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<750> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<749> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<748> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<747> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<746> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<745> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<744> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<743> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<742> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<741> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<740> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<739> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<738> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<737> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<736> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<735> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<734> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<733> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<732> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<731> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<730> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<729> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<728> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<727> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<726> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<725> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<724> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<723> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<722> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<721> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<720> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<719> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<718> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<717> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<716> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<715> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<714> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<713> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<712> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<711> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<710> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<709> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<708> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<707> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<706> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<705> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<704> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<703> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<702> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<701> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<700> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<699> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<698> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<697> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<696> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<695> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<694> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<693> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<692> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<691> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<690> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<689> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<688> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<687> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<686> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<685> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<684> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<683> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<682> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<681> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<680> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<679> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<678> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<677> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<676> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<675> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<674> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<673> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<672> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<671> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<670> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<669> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<668> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<667> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<666> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<665> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<664> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<663> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<662> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<661> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<660> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<659> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<658> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<657> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<656> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<655> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<654> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<653> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<652> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<651> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<650> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<649> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<648> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<647> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<646> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<645> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<644> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<643> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<642> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<641> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<640> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<639> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<638> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<637> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<636> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<635> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<634> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<633> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<632> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<631> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<630> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<629> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<628> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<627> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<626> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<625> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<624> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<623> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<622> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<621> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<620> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<619> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<618> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<617> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<616> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<615> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<614> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<613> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<612> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<611> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<610> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<609> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<608> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<607> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<606> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<605> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<604> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<603> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<602> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<601> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<600> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<599> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<598> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<597> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<596> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<595> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<594> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<593> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<592> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<591> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<590> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<589> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<588> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<587> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<586> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<585> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<584> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<583> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<582> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<581> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<580> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<579> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<578> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<577> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<576> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<575> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<574> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<573> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<572> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<571> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<570> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<569> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<568> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<567> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<566> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<565> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<564> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<563> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<562> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<561> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<560> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<559> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<558> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<557> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<556> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<555> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<554> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<553> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<552> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<551> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<550> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<549> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<548> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<547> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<546> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<545> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<544> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<543> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<542> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<541> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<540> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<539> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<538> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<537> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<536> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<535> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<534> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<533> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<532> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<531> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<530> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<529> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<528> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<527> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<526> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<525> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<524> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<523> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<522> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<521> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<520> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<519> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<518> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<517> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<516> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<515> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<514> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<513> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<512> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<511> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<510> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<509> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<508> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<507> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<506> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<505> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<504> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<503> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<502> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<501> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<500> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<499> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<498> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<497> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<496> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<495> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<494> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<493> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<492> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<491> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<490> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<489> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<488> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<487> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<486> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<485> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<484> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<483> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<482> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<481> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<480> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<479> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<478> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<477> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<476> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<475> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<474> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<473> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<472> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<471> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<470> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<469> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<468> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<467> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<466> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<465> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<464> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<463> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<462> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<461> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<460> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<459> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<458> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<457> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<456> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<455> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<454> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<453> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<452> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<451> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<450> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<449> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<448> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<447> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<446> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<445> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<444> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<443> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<442> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<441> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<440> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<439> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<438> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<437> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<436> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<435> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<434> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<433> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<432> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<431> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<430> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<429> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<428> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<427> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<426> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<425> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<424> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<423> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<422> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<421> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<420> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<419> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<418> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<417> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<416> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<415> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<414> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<413> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<412> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<411> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<410> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<409> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<408> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<407> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<406> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<405> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<404> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<403> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<402> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<401> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<400> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<399> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<398> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<397> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<396> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<395> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<394> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<393> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<392> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<391> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<390> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<389> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<388> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<387> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<386> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<385> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<384> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<383> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<382> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<381> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<380> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<379> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<378> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<377> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<376> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<375> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<374> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<373> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<372> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<371> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<370> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<369> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<368> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<367> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<366> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<365> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<364> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<363> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<362> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<361> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<360> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<359> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<358> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<357> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<356> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<355> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<354> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<353> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<352> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<351> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<350> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<349> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<348> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<347> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<346> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<345> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<344> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<343> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<342> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<341> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<340> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<339> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<338> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<337> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<336> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<335> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<334> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<333> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<332> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<331> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<330> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<329> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<328> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<327> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<326> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<325> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<324> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<323> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<322> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<321> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<320> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<319> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<318> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<317> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<316> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<315> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<314> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<313> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<312> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<311> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<310> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<309> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<308> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<307> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<306> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<305> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<304> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<303> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<302> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<301> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<300> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<299> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<298> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<297> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<296> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<295> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<294> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<293> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<292> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<291> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<290> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<289> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<288> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<287> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<286> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<285> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<284> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<283> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<282> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<281> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<280> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<279> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<278> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<277> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<276> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<275> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<274> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<273> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<272> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<271> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<270> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<269> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<268> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<267> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<266> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<265> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<264> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<263> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<262> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<261> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<260> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<259> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<258> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<257> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<256> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<255> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<254> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<253> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<252> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<251> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<250> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<249> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<248> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<247> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<246> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<245> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<244> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<243> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<242> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<241> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<240> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<239> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<238> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<237> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<236> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<235> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<234> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<233> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<232> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<231> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<230> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<229> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<228> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<227> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<226> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<225> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<224> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<223> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<222> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<221> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<220> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<219> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<218> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<217> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<216> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<215> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<214> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<213> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<212> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<211> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<210> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<209> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<208> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<207> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<206> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<205> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<204> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<203> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<202> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<201> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<200> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<199> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<198> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<197> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<196> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<195> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<194> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<193> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<192> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<191> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<190> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<189> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<188> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<187> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<186> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<185> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<184> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<183> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<182> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<181> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<180> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<179> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<178> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<177> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<176> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<175> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<174> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<173> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<172> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<171> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<170> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<169> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<168> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<167> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<166> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<165> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<164> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<163> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<162> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<161> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<160> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<159> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<158> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<157> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<156> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<155> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<154> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<153> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<152> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<151> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<150> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<149> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<148> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<147> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<146> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<145> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<144> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<143> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<142> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<141> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<140> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<139> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<138> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<137> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<136> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<135> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<134> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<133> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<132> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<131> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<130> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<129> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<128> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<127> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<126> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<125> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<124> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<123> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<122> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<121> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<120> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<119> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<118> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<117> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<116> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<115> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<114> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<113> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<112> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<111> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<110> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<109> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<108> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<107> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<106> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<105> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<104> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<103> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<102> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<101> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<100> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<99> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<98> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<97> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<96> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<95> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<94> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<93> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<92> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<91> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<90> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<89> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<88> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<87> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<86> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<85> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<84> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<83> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<82> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<81> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<80> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<79> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<78> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<77> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<76> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<75> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<74> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<73> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<72> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<71> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<70> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<69> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<68> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<67> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<66> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<65> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<64> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<63> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<62> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<61> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<60> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<59> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<58> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<57> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<56> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<55> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<54> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<53> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<52> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<51> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<50> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<49> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<48> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<47> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<46> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<45> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<44> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<43> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<42> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<41> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<40> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<39> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<38> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<37> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<36> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<35> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<34> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<33> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<32> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<31> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<30> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<29> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<28> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<27> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<26> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<25> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<24> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<23> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<22> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<21> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<20> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<19> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<18> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<17> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<16> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<15> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<14> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<13> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<12> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<11> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<10> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<9> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<8> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<7> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<6> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<5> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<4> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<3> net16<3> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<2> net16<2> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<1> net16<1> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC16<0> net16<0> outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM22<3> net15<3> sw<7> net16<3> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22<2> net15<2> sw<7> net16<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22<1> net15<1> sw<7> net16<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22<0> net15<0> sw<7> net16<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=11 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23<3> GND sw<7> net15<3> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23<2> GND sw<7> net15<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23<1> GND sw<7> net15<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23<0> GND sw<7> net15<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24<3> GND sw<7> net16<3> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24<2> GND sw<7> net16<2> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24<1> GND sw<7> net16<1> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24<0> GND sw<7> net16<0> GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC15<1023> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1022> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1021> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1020> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1019> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1018> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1017> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1016> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1015> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1014> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1013> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1012> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1011> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1010> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1009> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1008> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1007> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1006> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1005> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1004> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1003> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1002> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1001> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1000> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<999> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<998> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<997> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<996> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<995> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<994> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<993> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<992> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<991> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<990> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<989> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<988> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<987> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<986> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<985> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<984> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<983> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<982> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<981> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<980> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<979> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<978> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<977> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<976> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<975> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<974> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<973> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<972> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<971> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<970> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<969> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<968> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<967> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<966> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<965> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<964> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<963> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<962> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<961> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<960> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<959> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<958> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<957> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<956> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<955> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<954> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<953> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<952> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<951> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<950> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<949> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<948> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<947> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<946> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<945> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<944> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<943> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<942> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<941> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<940> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<939> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<938> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<937> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<936> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<935> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<934> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<933> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<932> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<931> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<930> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<929> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<928> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<927> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<926> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<925> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<924> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<923> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<922> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<921> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<920> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<919> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<918> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<917> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<916> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<915> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<914> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<913> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<912> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<911> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<910> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<909> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<908> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<907> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<906> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<905> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<904> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<903> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<902> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<901> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<900> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<899> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<898> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<897> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<896> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<895> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<894> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<893> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<892> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<891> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<890> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<889> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<888> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<887> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<886> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<885> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<884> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<883> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<882> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<881> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<880> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<879> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<878> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<877> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<876> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<875> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<874> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<873> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<872> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<871> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<870> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<869> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<868> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<867> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<866> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<865> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<864> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<863> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<862> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<861> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<860> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<859> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<858> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<857> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<856> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<855> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<854> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<853> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<852> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<851> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<850> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<849> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<848> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<847> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<846> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<845> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<844> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<843> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<842> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<841> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<840> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<839> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<838> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<837> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<836> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<835> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<834> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<833> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<832> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<831> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<830> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<829> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<828> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<827> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<826> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<825> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<824> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<823> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<822> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<821> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<820> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<819> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<818> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<817> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<816> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<815> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<814> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<813> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<812> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<811> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<810> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<809> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<808> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<807> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<806> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<805> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<804> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<803> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<802> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<801> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<800> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<799> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<798> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<797> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<796> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<795> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<794> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<793> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<792> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<791> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<790> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<789> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<788> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<787> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<786> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<785> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<784> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<783> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<782> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<781> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<780> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<779> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<778> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<777> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<776> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<775> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<774> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<773> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<772> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<771> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<770> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<769> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<768> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<767> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<766> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<765> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<764> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<763> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<762> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<761> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<760> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<759> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<758> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<757> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<756> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<755> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<754> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<753> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<752> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<751> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<750> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<749> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<748> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<747> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<746> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<745> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<744> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<743> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<742> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<741> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<740> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<739> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<738> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<737> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<736> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<735> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<734> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<733> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<732> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<731> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<730> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<729> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<728> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<727> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<726> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<725> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<724> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<723> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<722> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<721> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<720> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<719> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<718> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<717> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<716> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<715> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<714> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<713> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<712> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<711> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<710> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<709> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<708> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<707> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<706> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<705> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<704> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<703> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<702> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<701> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<700> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<699> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<698> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<697> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<696> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<695> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<694> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<693> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<692> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<691> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<690> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<689> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<688> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<687> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<686> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<685> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<684> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<683> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<682> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<681> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<680> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<679> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<678> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<677> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<676> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<675> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<674> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<673> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<672> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<671> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<670> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<669> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<668> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<667> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<666> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<665> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<664> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<663> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<662> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<661> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<660> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<659> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<658> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<657> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<656> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<655> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<654> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<653> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<652> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<651> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<650> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<649> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<648> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<647> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<646> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<645> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<644> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<643> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<642> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<641> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<640> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<639> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<638> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<637> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<636> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<635> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<634> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<633> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<632> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<631> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<630> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<629> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<628> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<627> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<626> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<625> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<624> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<623> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<622> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<621> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<620> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<619> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<618> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<617> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<616> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<615> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<614> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<613> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<612> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<611> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<610> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<609> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<608> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<607> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<606> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<605> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<604> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<603> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<602> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<601> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<600> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<599> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<598> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<597> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<596> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<595> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<594> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<593> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<592> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<591> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<590> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<589> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<588> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<587> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<586> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<585> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<584> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<583> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<582> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<581> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<580> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<579> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<578> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<577> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<576> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<575> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<574> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<573> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<572> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<571> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<570> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<569> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<568> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<567> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<566> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<565> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<564> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<563> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<562> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<561> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<560> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<559> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<558> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<557> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<556> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<555> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<554> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<553> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<552> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<551> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<550> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<549> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<548> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<547> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<546> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<545> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<544> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<543> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<542> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<541> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<540> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<539> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<538> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<537> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<536> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<535> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<534> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<533> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<532> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<531> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<530> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<529> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<528> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<527> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<526> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<525> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<524> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<523> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<522> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<521> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<520> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<519> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<518> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<517> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<516> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<515> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<514> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<513> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<512> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<511> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<510> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<509> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<508> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<507> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<506> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<505> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<504> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<503> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<502> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<501> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<500> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<499> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<498> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<497> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<496> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<495> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<494> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<493> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<492> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<491> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<490> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<489> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<488> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<487> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<486> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<485> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<484> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<483> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<482> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<481> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<480> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<479> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<478> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<477> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<476> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<475> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<474> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<473> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<472> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<471> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<470> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<469> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<468> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<467> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<466> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<465> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<464> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<463> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<462> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<461> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<460> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<459> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<458> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<457> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<456> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<455> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<454> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<453> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<452> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<451> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<450> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<449> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<448> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<447> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<446> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<445> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<444> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<443> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<442> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<441> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<440> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<439> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<438> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<437> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<436> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<435> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<434> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<433> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<432> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<431> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<430> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<429> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<428> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<427> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<426> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<425> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<424> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<423> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<422> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<421> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<420> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<419> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<418> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<417> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<416> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<415> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<414> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<413> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<412> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<411> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<410> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<409> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<408> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<407> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<406> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<405> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<404> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<403> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<402> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<401> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<400> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<399> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<398> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<397> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<396> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<395> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<394> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<393> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<392> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<391> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<390> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<389> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<388> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<387> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<386> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<385> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<384> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<383> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<382> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<381> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<380> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<379> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<378> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<377> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<376> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<375> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<374> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<373> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<372> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<371> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<370> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<369> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<368> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<367> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<366> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<365> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<364> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<363> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<362> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<361> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<360> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<359> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<358> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<357> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<356> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<355> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<354> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<353> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<352> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<351> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<350> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<349> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<348> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<347> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<346> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<345> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<344> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<343> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<342> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<341> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<340> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<339> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<338> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<337> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<336> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<335> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<334> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<333> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<332> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<331> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<330> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<329> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<328> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<327> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<326> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<325> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<324> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<323> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<322> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<321> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<320> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<319> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<318> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<317> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<316> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<315> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<314> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<313> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<312> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<311> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<310> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<309> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<308> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<307> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<306> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<305> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<304> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<303> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<302> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<301> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<300> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<299> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<298> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<297> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<296> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<295> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<294> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<293> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<292> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<291> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<290> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<289> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<288> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<287> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<286> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<285> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<284> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<283> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<282> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<281> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<280> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<279> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<278> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<277> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<276> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<275> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<274> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<273> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<272> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<271> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<270> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<269> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<268> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<267> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<266> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<265> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<264> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<263> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<262> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<261> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<260> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<259> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<258> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<257> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<256> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<255> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<254> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<253> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<252> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<251> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<250> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<249> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<248> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<247> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<246> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<245> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<244> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<243> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<242> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<241> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<240> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<239> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<238> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<237> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<236> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<235> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<234> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<233> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<232> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<231> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<230> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<229> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<228> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<227> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<226> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<225> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<224> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<223> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<222> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<221> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<220> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<219> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<218> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<217> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<216> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<215> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<214> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<213> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<212> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<211> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<210> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<209> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<208> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<207> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<206> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<205> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<204> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<203> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<202> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<201> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<200> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<199> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<198> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<197> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<196> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<195> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<194> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<193> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<192> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<191> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<190> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<189> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<188> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<187> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<186> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<185> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<184> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<183> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<182> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<181> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<180> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<179> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<178> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<177> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<176> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<175> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<174> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<173> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<172> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<171> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<170> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<169> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<168> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<167> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<166> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<165> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<164> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<163> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<162> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<161> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<160> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<159> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<158> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<157> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<156> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<155> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<154> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<153> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<152> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<151> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<150> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<149> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<148> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<147> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<146> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<145> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<144> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<143> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<142> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<141> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<140> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<139> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<138> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<137> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<136> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<135> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<134> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<133> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<132> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<131> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<130> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<129> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<128> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<127> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<126> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<125> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<124> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<123> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<122> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<121> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<120> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<119> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<118> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<117> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<116> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<115> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<114> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<113> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<112> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<111> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<110> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<109> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<108> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<107> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<106> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<105> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<104> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<103> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<102> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<101> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<100> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<99> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<98> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<97> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<96> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<95> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<94> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<93> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<92> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<91> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<90> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<89> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<88> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<87> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<86> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<85> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<84> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<83> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<82> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<81> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<80> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<79> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<78> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<77> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<76> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<75> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<74> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<73> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<72> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<71> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<70> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<69> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<68> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<67> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<66> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<65> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<64> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<63> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<62> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<61> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<60> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<59> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<58> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<57> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<56> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<55> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<54> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<53> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<52> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<51> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<50> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<49> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<48> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<47> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<46> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<45> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<44> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<43> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<42> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<41> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<40> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<39> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<38> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<37> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<36> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<35> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<34> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<33> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<32> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<31> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<30> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<29> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<28> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<27> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<26> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<25> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<24> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<23> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<22> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<21> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<20> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<19> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<18> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<17> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<16> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<15> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<14> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<13> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<12> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<11> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<10> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<9> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<8> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<7> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<6> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<5> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<4> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<3> outp net15<3> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<2> outp net15<2> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<1> outp net15<1> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC15<0> outp net15<0> sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
.ends
