* NGSPICE file created from diff_pair_sample_1316.ext - technology: sky130A

.subckt diff_pair_sample_1316 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=0 ps=0 w=9.65 l=0.16
X1 VTAIL.t11 VP.t0 VDD1.t3 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=2.4125 ps=10.15 w=9.65 l=0.16
X2 VDD2.t5 VN.t0 VTAIL.t3 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=2.4125 ps=10.15 w=9.65 l=0.16
X3 VTAIL.t4 VN.t1 VDD2.t4 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=2.4125 ps=10.15 w=9.65 l=0.16
X4 VTAIL.t10 VP.t1 VDD1.t1 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=2.4125 ps=10.15 w=9.65 l=0.16
X5 VDD2.t3 VN.t2 VTAIL.t5 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=4.58375 ps=20.25 w=9.65 l=0.16
X6 VDD2.t2 VN.t3 VTAIL.t2 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=2.4125 ps=10.15 w=9.65 l=0.16
X7 B.t8 B.t6 B.t7 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=0 ps=0 w=9.65 l=0.16
X8 VTAIL.t1 VN.t4 VDD2.t1 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=2.4125 ps=10.15 w=9.65 l=0.16
X9 VDD1.t4 VP.t2 VTAIL.t9 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=4.58375 ps=20.25 w=9.65 l=0.16
X10 VDD1.t5 VP.t3 VTAIL.t8 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=4.58375 ps=20.25 w=9.65 l=0.16
X11 B.t5 B.t3 B.t4 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=0 ps=0 w=9.65 l=0.16
X12 B.t2 B.t0 B.t1 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=0 ps=0 w=9.65 l=0.16
X13 VDD1.t2 VP.t4 VTAIL.t7 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=2.4125 ps=10.15 w=9.65 l=0.16
X14 VDD2.t0 VN.t5 VTAIL.t0 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=2.4125 pd=10.15 as=4.58375 ps=20.25 w=9.65 l=0.16
X15 VDD1.t0 VP.t5 VTAIL.t6 w_n1498_n2898# sky130_fd_pr__pfet_01v8 ad=4.58375 pd=20.25 as=2.4125 ps=10.15 w=9.65 l=0.16
R0 B.n88 B.t6 1704.94
R1 B.n96 B.t9 1704.94
R2 B.n28 B.t3 1704.94
R3 B.n34 B.t0 1704.94
R4 B.n315 B.n314 585
R5 B.n316 B.n53 585
R6 B.n318 B.n317 585
R7 B.n319 B.n52 585
R8 B.n321 B.n320 585
R9 B.n322 B.n51 585
R10 B.n324 B.n323 585
R11 B.n325 B.n50 585
R12 B.n327 B.n326 585
R13 B.n328 B.n49 585
R14 B.n330 B.n329 585
R15 B.n331 B.n48 585
R16 B.n333 B.n332 585
R17 B.n334 B.n47 585
R18 B.n336 B.n335 585
R19 B.n337 B.n46 585
R20 B.n339 B.n338 585
R21 B.n340 B.n45 585
R22 B.n342 B.n341 585
R23 B.n343 B.n44 585
R24 B.n345 B.n344 585
R25 B.n346 B.n43 585
R26 B.n348 B.n347 585
R27 B.n349 B.n42 585
R28 B.n351 B.n350 585
R29 B.n352 B.n41 585
R30 B.n354 B.n353 585
R31 B.n355 B.n40 585
R32 B.n357 B.n356 585
R33 B.n358 B.n39 585
R34 B.n360 B.n359 585
R35 B.n361 B.n38 585
R36 B.n363 B.n362 585
R37 B.n364 B.n37 585
R38 B.n366 B.n365 585
R39 B.n368 B.n367 585
R40 B.n369 B.n33 585
R41 B.n371 B.n370 585
R42 B.n372 B.n32 585
R43 B.n374 B.n373 585
R44 B.n375 B.n31 585
R45 B.n377 B.n376 585
R46 B.n378 B.n30 585
R47 B.n380 B.n379 585
R48 B.n382 B.n27 585
R49 B.n384 B.n383 585
R50 B.n385 B.n26 585
R51 B.n387 B.n386 585
R52 B.n388 B.n25 585
R53 B.n390 B.n389 585
R54 B.n391 B.n24 585
R55 B.n393 B.n392 585
R56 B.n394 B.n23 585
R57 B.n396 B.n395 585
R58 B.n397 B.n22 585
R59 B.n399 B.n398 585
R60 B.n400 B.n21 585
R61 B.n402 B.n401 585
R62 B.n403 B.n20 585
R63 B.n405 B.n404 585
R64 B.n406 B.n19 585
R65 B.n408 B.n407 585
R66 B.n409 B.n18 585
R67 B.n411 B.n410 585
R68 B.n412 B.n17 585
R69 B.n414 B.n413 585
R70 B.n415 B.n16 585
R71 B.n417 B.n416 585
R72 B.n418 B.n15 585
R73 B.n420 B.n419 585
R74 B.n421 B.n14 585
R75 B.n423 B.n422 585
R76 B.n424 B.n13 585
R77 B.n426 B.n425 585
R78 B.n427 B.n12 585
R79 B.n429 B.n428 585
R80 B.n430 B.n11 585
R81 B.n432 B.n431 585
R82 B.n433 B.n10 585
R83 B.n313 B.n54 585
R84 B.n312 B.n311 585
R85 B.n310 B.n55 585
R86 B.n309 B.n308 585
R87 B.n307 B.n56 585
R88 B.n306 B.n305 585
R89 B.n304 B.n57 585
R90 B.n303 B.n302 585
R91 B.n301 B.n58 585
R92 B.n300 B.n299 585
R93 B.n298 B.n59 585
R94 B.n297 B.n296 585
R95 B.n295 B.n60 585
R96 B.n294 B.n293 585
R97 B.n292 B.n61 585
R98 B.n291 B.n290 585
R99 B.n289 B.n62 585
R100 B.n288 B.n287 585
R101 B.n286 B.n63 585
R102 B.n285 B.n284 585
R103 B.n283 B.n64 585
R104 B.n282 B.n281 585
R105 B.n280 B.n65 585
R106 B.n279 B.n278 585
R107 B.n277 B.n66 585
R108 B.n276 B.n275 585
R109 B.n274 B.n67 585
R110 B.n273 B.n272 585
R111 B.n271 B.n68 585
R112 B.n270 B.n269 585
R113 B.n268 B.n69 585
R114 B.n267 B.n266 585
R115 B.n265 B.n70 585
R116 B.n145 B.n114 585
R117 B.n147 B.n146 585
R118 B.n148 B.n113 585
R119 B.n150 B.n149 585
R120 B.n151 B.n112 585
R121 B.n153 B.n152 585
R122 B.n154 B.n111 585
R123 B.n156 B.n155 585
R124 B.n157 B.n110 585
R125 B.n159 B.n158 585
R126 B.n160 B.n109 585
R127 B.n162 B.n161 585
R128 B.n163 B.n108 585
R129 B.n165 B.n164 585
R130 B.n166 B.n107 585
R131 B.n168 B.n167 585
R132 B.n169 B.n106 585
R133 B.n171 B.n170 585
R134 B.n172 B.n105 585
R135 B.n174 B.n173 585
R136 B.n175 B.n104 585
R137 B.n177 B.n176 585
R138 B.n178 B.n103 585
R139 B.n180 B.n179 585
R140 B.n181 B.n102 585
R141 B.n183 B.n182 585
R142 B.n184 B.n101 585
R143 B.n186 B.n185 585
R144 B.n187 B.n100 585
R145 B.n189 B.n188 585
R146 B.n190 B.n99 585
R147 B.n192 B.n191 585
R148 B.n193 B.n98 585
R149 B.n195 B.n194 585
R150 B.n196 B.n95 585
R151 B.n199 B.n198 585
R152 B.n200 B.n94 585
R153 B.n202 B.n201 585
R154 B.n203 B.n93 585
R155 B.n205 B.n204 585
R156 B.n206 B.n92 585
R157 B.n208 B.n207 585
R158 B.n209 B.n91 585
R159 B.n211 B.n210 585
R160 B.n213 B.n212 585
R161 B.n214 B.n87 585
R162 B.n216 B.n215 585
R163 B.n217 B.n86 585
R164 B.n219 B.n218 585
R165 B.n220 B.n85 585
R166 B.n222 B.n221 585
R167 B.n223 B.n84 585
R168 B.n225 B.n224 585
R169 B.n226 B.n83 585
R170 B.n228 B.n227 585
R171 B.n229 B.n82 585
R172 B.n231 B.n230 585
R173 B.n232 B.n81 585
R174 B.n234 B.n233 585
R175 B.n235 B.n80 585
R176 B.n237 B.n236 585
R177 B.n238 B.n79 585
R178 B.n240 B.n239 585
R179 B.n241 B.n78 585
R180 B.n243 B.n242 585
R181 B.n244 B.n77 585
R182 B.n246 B.n245 585
R183 B.n247 B.n76 585
R184 B.n249 B.n248 585
R185 B.n250 B.n75 585
R186 B.n252 B.n251 585
R187 B.n253 B.n74 585
R188 B.n255 B.n254 585
R189 B.n256 B.n73 585
R190 B.n258 B.n257 585
R191 B.n259 B.n72 585
R192 B.n261 B.n260 585
R193 B.n262 B.n71 585
R194 B.n264 B.n263 585
R195 B.n144 B.n143 585
R196 B.n142 B.n115 585
R197 B.n141 B.n140 585
R198 B.n139 B.n116 585
R199 B.n138 B.n137 585
R200 B.n136 B.n117 585
R201 B.n135 B.n134 585
R202 B.n133 B.n118 585
R203 B.n132 B.n131 585
R204 B.n130 B.n119 585
R205 B.n129 B.n128 585
R206 B.n127 B.n120 585
R207 B.n126 B.n125 585
R208 B.n124 B.n121 585
R209 B.n123 B.n122 585
R210 B.n2 B.n0 585
R211 B.n457 B.n1 585
R212 B.n456 B.n455 585
R213 B.n454 B.n3 585
R214 B.n453 B.n452 585
R215 B.n451 B.n4 585
R216 B.n450 B.n449 585
R217 B.n448 B.n5 585
R218 B.n447 B.n446 585
R219 B.n445 B.n6 585
R220 B.n444 B.n443 585
R221 B.n442 B.n7 585
R222 B.n441 B.n440 585
R223 B.n439 B.n8 585
R224 B.n438 B.n437 585
R225 B.n436 B.n9 585
R226 B.n435 B.n434 585
R227 B.n459 B.n458 585
R228 B.n145 B.n144 478.086
R229 B.n434 B.n433 478.086
R230 B.n265 B.n264 478.086
R231 B.n314 B.n313 478.086
R232 B.n144 B.n115 163.367
R233 B.n140 B.n115 163.367
R234 B.n140 B.n139 163.367
R235 B.n139 B.n138 163.367
R236 B.n138 B.n117 163.367
R237 B.n134 B.n117 163.367
R238 B.n134 B.n133 163.367
R239 B.n133 B.n132 163.367
R240 B.n132 B.n119 163.367
R241 B.n128 B.n119 163.367
R242 B.n128 B.n127 163.367
R243 B.n127 B.n126 163.367
R244 B.n126 B.n121 163.367
R245 B.n122 B.n121 163.367
R246 B.n122 B.n2 163.367
R247 B.n458 B.n2 163.367
R248 B.n458 B.n457 163.367
R249 B.n457 B.n456 163.367
R250 B.n456 B.n3 163.367
R251 B.n452 B.n3 163.367
R252 B.n452 B.n451 163.367
R253 B.n451 B.n450 163.367
R254 B.n450 B.n5 163.367
R255 B.n446 B.n5 163.367
R256 B.n446 B.n445 163.367
R257 B.n445 B.n444 163.367
R258 B.n444 B.n7 163.367
R259 B.n440 B.n7 163.367
R260 B.n440 B.n439 163.367
R261 B.n439 B.n438 163.367
R262 B.n438 B.n9 163.367
R263 B.n434 B.n9 163.367
R264 B.n146 B.n145 163.367
R265 B.n146 B.n113 163.367
R266 B.n150 B.n113 163.367
R267 B.n151 B.n150 163.367
R268 B.n152 B.n151 163.367
R269 B.n152 B.n111 163.367
R270 B.n156 B.n111 163.367
R271 B.n157 B.n156 163.367
R272 B.n158 B.n157 163.367
R273 B.n158 B.n109 163.367
R274 B.n162 B.n109 163.367
R275 B.n163 B.n162 163.367
R276 B.n164 B.n163 163.367
R277 B.n164 B.n107 163.367
R278 B.n168 B.n107 163.367
R279 B.n169 B.n168 163.367
R280 B.n170 B.n169 163.367
R281 B.n170 B.n105 163.367
R282 B.n174 B.n105 163.367
R283 B.n175 B.n174 163.367
R284 B.n176 B.n175 163.367
R285 B.n176 B.n103 163.367
R286 B.n180 B.n103 163.367
R287 B.n181 B.n180 163.367
R288 B.n182 B.n181 163.367
R289 B.n182 B.n101 163.367
R290 B.n186 B.n101 163.367
R291 B.n187 B.n186 163.367
R292 B.n188 B.n187 163.367
R293 B.n188 B.n99 163.367
R294 B.n192 B.n99 163.367
R295 B.n193 B.n192 163.367
R296 B.n194 B.n193 163.367
R297 B.n194 B.n95 163.367
R298 B.n199 B.n95 163.367
R299 B.n200 B.n199 163.367
R300 B.n201 B.n200 163.367
R301 B.n201 B.n93 163.367
R302 B.n205 B.n93 163.367
R303 B.n206 B.n205 163.367
R304 B.n207 B.n206 163.367
R305 B.n207 B.n91 163.367
R306 B.n211 B.n91 163.367
R307 B.n212 B.n211 163.367
R308 B.n212 B.n87 163.367
R309 B.n216 B.n87 163.367
R310 B.n217 B.n216 163.367
R311 B.n218 B.n217 163.367
R312 B.n218 B.n85 163.367
R313 B.n222 B.n85 163.367
R314 B.n223 B.n222 163.367
R315 B.n224 B.n223 163.367
R316 B.n224 B.n83 163.367
R317 B.n228 B.n83 163.367
R318 B.n229 B.n228 163.367
R319 B.n230 B.n229 163.367
R320 B.n230 B.n81 163.367
R321 B.n234 B.n81 163.367
R322 B.n235 B.n234 163.367
R323 B.n236 B.n235 163.367
R324 B.n236 B.n79 163.367
R325 B.n240 B.n79 163.367
R326 B.n241 B.n240 163.367
R327 B.n242 B.n241 163.367
R328 B.n242 B.n77 163.367
R329 B.n246 B.n77 163.367
R330 B.n247 B.n246 163.367
R331 B.n248 B.n247 163.367
R332 B.n248 B.n75 163.367
R333 B.n252 B.n75 163.367
R334 B.n253 B.n252 163.367
R335 B.n254 B.n253 163.367
R336 B.n254 B.n73 163.367
R337 B.n258 B.n73 163.367
R338 B.n259 B.n258 163.367
R339 B.n260 B.n259 163.367
R340 B.n260 B.n71 163.367
R341 B.n264 B.n71 163.367
R342 B.n266 B.n265 163.367
R343 B.n266 B.n69 163.367
R344 B.n270 B.n69 163.367
R345 B.n271 B.n270 163.367
R346 B.n272 B.n271 163.367
R347 B.n272 B.n67 163.367
R348 B.n276 B.n67 163.367
R349 B.n277 B.n276 163.367
R350 B.n278 B.n277 163.367
R351 B.n278 B.n65 163.367
R352 B.n282 B.n65 163.367
R353 B.n283 B.n282 163.367
R354 B.n284 B.n283 163.367
R355 B.n284 B.n63 163.367
R356 B.n288 B.n63 163.367
R357 B.n289 B.n288 163.367
R358 B.n290 B.n289 163.367
R359 B.n290 B.n61 163.367
R360 B.n294 B.n61 163.367
R361 B.n295 B.n294 163.367
R362 B.n296 B.n295 163.367
R363 B.n296 B.n59 163.367
R364 B.n300 B.n59 163.367
R365 B.n301 B.n300 163.367
R366 B.n302 B.n301 163.367
R367 B.n302 B.n57 163.367
R368 B.n306 B.n57 163.367
R369 B.n307 B.n306 163.367
R370 B.n308 B.n307 163.367
R371 B.n308 B.n55 163.367
R372 B.n312 B.n55 163.367
R373 B.n313 B.n312 163.367
R374 B.n433 B.n432 163.367
R375 B.n432 B.n11 163.367
R376 B.n428 B.n11 163.367
R377 B.n428 B.n427 163.367
R378 B.n427 B.n426 163.367
R379 B.n426 B.n13 163.367
R380 B.n422 B.n13 163.367
R381 B.n422 B.n421 163.367
R382 B.n421 B.n420 163.367
R383 B.n420 B.n15 163.367
R384 B.n416 B.n15 163.367
R385 B.n416 B.n415 163.367
R386 B.n415 B.n414 163.367
R387 B.n414 B.n17 163.367
R388 B.n410 B.n17 163.367
R389 B.n410 B.n409 163.367
R390 B.n409 B.n408 163.367
R391 B.n408 B.n19 163.367
R392 B.n404 B.n19 163.367
R393 B.n404 B.n403 163.367
R394 B.n403 B.n402 163.367
R395 B.n402 B.n21 163.367
R396 B.n398 B.n21 163.367
R397 B.n398 B.n397 163.367
R398 B.n397 B.n396 163.367
R399 B.n396 B.n23 163.367
R400 B.n392 B.n23 163.367
R401 B.n392 B.n391 163.367
R402 B.n391 B.n390 163.367
R403 B.n390 B.n25 163.367
R404 B.n386 B.n25 163.367
R405 B.n386 B.n385 163.367
R406 B.n385 B.n384 163.367
R407 B.n384 B.n27 163.367
R408 B.n379 B.n27 163.367
R409 B.n379 B.n378 163.367
R410 B.n378 B.n377 163.367
R411 B.n377 B.n31 163.367
R412 B.n373 B.n31 163.367
R413 B.n373 B.n372 163.367
R414 B.n372 B.n371 163.367
R415 B.n371 B.n33 163.367
R416 B.n367 B.n33 163.367
R417 B.n367 B.n366 163.367
R418 B.n366 B.n37 163.367
R419 B.n362 B.n37 163.367
R420 B.n362 B.n361 163.367
R421 B.n361 B.n360 163.367
R422 B.n360 B.n39 163.367
R423 B.n356 B.n39 163.367
R424 B.n356 B.n355 163.367
R425 B.n355 B.n354 163.367
R426 B.n354 B.n41 163.367
R427 B.n350 B.n41 163.367
R428 B.n350 B.n349 163.367
R429 B.n349 B.n348 163.367
R430 B.n348 B.n43 163.367
R431 B.n344 B.n43 163.367
R432 B.n344 B.n343 163.367
R433 B.n343 B.n342 163.367
R434 B.n342 B.n45 163.367
R435 B.n338 B.n45 163.367
R436 B.n338 B.n337 163.367
R437 B.n337 B.n336 163.367
R438 B.n336 B.n47 163.367
R439 B.n332 B.n47 163.367
R440 B.n332 B.n331 163.367
R441 B.n331 B.n330 163.367
R442 B.n330 B.n49 163.367
R443 B.n326 B.n49 163.367
R444 B.n326 B.n325 163.367
R445 B.n325 B.n324 163.367
R446 B.n324 B.n51 163.367
R447 B.n320 B.n51 163.367
R448 B.n320 B.n319 163.367
R449 B.n319 B.n318 163.367
R450 B.n318 B.n53 163.367
R451 B.n314 B.n53 163.367
R452 B.n88 B.t8 124.865
R453 B.n34 B.t1 124.865
R454 B.n96 B.t11 124.853
R455 B.n28 B.t4 124.853
R456 B.n89 B.t7 112.064
R457 B.n35 B.t2 112.064
R458 B.n97 B.t10 112.053
R459 B.n29 B.t5 112.053
R460 B.n90 B.n89 59.5399
R461 B.n197 B.n97 59.5399
R462 B.n381 B.n29 59.5399
R463 B.n36 B.n35 59.5399
R464 B.n435 B.n10 31.0639
R465 B.n315 B.n54 31.0639
R466 B.n263 B.n70 31.0639
R467 B.n143 B.n114 31.0639
R468 B B.n459 18.0485
R469 B.n89 B.n88 12.8005
R470 B.n97 B.n96 12.8005
R471 B.n29 B.n28 12.8005
R472 B.n35 B.n34 12.8005
R473 B.n431 B.n10 10.6151
R474 B.n431 B.n430 10.6151
R475 B.n430 B.n429 10.6151
R476 B.n429 B.n12 10.6151
R477 B.n425 B.n12 10.6151
R478 B.n425 B.n424 10.6151
R479 B.n424 B.n423 10.6151
R480 B.n423 B.n14 10.6151
R481 B.n419 B.n14 10.6151
R482 B.n419 B.n418 10.6151
R483 B.n418 B.n417 10.6151
R484 B.n417 B.n16 10.6151
R485 B.n413 B.n16 10.6151
R486 B.n413 B.n412 10.6151
R487 B.n412 B.n411 10.6151
R488 B.n411 B.n18 10.6151
R489 B.n407 B.n18 10.6151
R490 B.n407 B.n406 10.6151
R491 B.n406 B.n405 10.6151
R492 B.n405 B.n20 10.6151
R493 B.n401 B.n20 10.6151
R494 B.n401 B.n400 10.6151
R495 B.n400 B.n399 10.6151
R496 B.n399 B.n22 10.6151
R497 B.n395 B.n22 10.6151
R498 B.n395 B.n394 10.6151
R499 B.n394 B.n393 10.6151
R500 B.n393 B.n24 10.6151
R501 B.n389 B.n24 10.6151
R502 B.n389 B.n388 10.6151
R503 B.n388 B.n387 10.6151
R504 B.n387 B.n26 10.6151
R505 B.n383 B.n26 10.6151
R506 B.n383 B.n382 10.6151
R507 B.n380 B.n30 10.6151
R508 B.n376 B.n30 10.6151
R509 B.n376 B.n375 10.6151
R510 B.n375 B.n374 10.6151
R511 B.n374 B.n32 10.6151
R512 B.n370 B.n32 10.6151
R513 B.n370 B.n369 10.6151
R514 B.n369 B.n368 10.6151
R515 B.n365 B.n364 10.6151
R516 B.n364 B.n363 10.6151
R517 B.n363 B.n38 10.6151
R518 B.n359 B.n38 10.6151
R519 B.n359 B.n358 10.6151
R520 B.n358 B.n357 10.6151
R521 B.n357 B.n40 10.6151
R522 B.n353 B.n40 10.6151
R523 B.n353 B.n352 10.6151
R524 B.n352 B.n351 10.6151
R525 B.n351 B.n42 10.6151
R526 B.n347 B.n42 10.6151
R527 B.n347 B.n346 10.6151
R528 B.n346 B.n345 10.6151
R529 B.n345 B.n44 10.6151
R530 B.n341 B.n44 10.6151
R531 B.n341 B.n340 10.6151
R532 B.n340 B.n339 10.6151
R533 B.n339 B.n46 10.6151
R534 B.n335 B.n46 10.6151
R535 B.n335 B.n334 10.6151
R536 B.n334 B.n333 10.6151
R537 B.n333 B.n48 10.6151
R538 B.n329 B.n48 10.6151
R539 B.n329 B.n328 10.6151
R540 B.n328 B.n327 10.6151
R541 B.n327 B.n50 10.6151
R542 B.n323 B.n50 10.6151
R543 B.n323 B.n322 10.6151
R544 B.n322 B.n321 10.6151
R545 B.n321 B.n52 10.6151
R546 B.n317 B.n52 10.6151
R547 B.n317 B.n316 10.6151
R548 B.n316 B.n315 10.6151
R549 B.n267 B.n70 10.6151
R550 B.n268 B.n267 10.6151
R551 B.n269 B.n268 10.6151
R552 B.n269 B.n68 10.6151
R553 B.n273 B.n68 10.6151
R554 B.n274 B.n273 10.6151
R555 B.n275 B.n274 10.6151
R556 B.n275 B.n66 10.6151
R557 B.n279 B.n66 10.6151
R558 B.n280 B.n279 10.6151
R559 B.n281 B.n280 10.6151
R560 B.n281 B.n64 10.6151
R561 B.n285 B.n64 10.6151
R562 B.n286 B.n285 10.6151
R563 B.n287 B.n286 10.6151
R564 B.n287 B.n62 10.6151
R565 B.n291 B.n62 10.6151
R566 B.n292 B.n291 10.6151
R567 B.n293 B.n292 10.6151
R568 B.n293 B.n60 10.6151
R569 B.n297 B.n60 10.6151
R570 B.n298 B.n297 10.6151
R571 B.n299 B.n298 10.6151
R572 B.n299 B.n58 10.6151
R573 B.n303 B.n58 10.6151
R574 B.n304 B.n303 10.6151
R575 B.n305 B.n304 10.6151
R576 B.n305 B.n56 10.6151
R577 B.n309 B.n56 10.6151
R578 B.n310 B.n309 10.6151
R579 B.n311 B.n310 10.6151
R580 B.n311 B.n54 10.6151
R581 B.n147 B.n114 10.6151
R582 B.n148 B.n147 10.6151
R583 B.n149 B.n148 10.6151
R584 B.n149 B.n112 10.6151
R585 B.n153 B.n112 10.6151
R586 B.n154 B.n153 10.6151
R587 B.n155 B.n154 10.6151
R588 B.n155 B.n110 10.6151
R589 B.n159 B.n110 10.6151
R590 B.n160 B.n159 10.6151
R591 B.n161 B.n160 10.6151
R592 B.n161 B.n108 10.6151
R593 B.n165 B.n108 10.6151
R594 B.n166 B.n165 10.6151
R595 B.n167 B.n166 10.6151
R596 B.n167 B.n106 10.6151
R597 B.n171 B.n106 10.6151
R598 B.n172 B.n171 10.6151
R599 B.n173 B.n172 10.6151
R600 B.n173 B.n104 10.6151
R601 B.n177 B.n104 10.6151
R602 B.n178 B.n177 10.6151
R603 B.n179 B.n178 10.6151
R604 B.n179 B.n102 10.6151
R605 B.n183 B.n102 10.6151
R606 B.n184 B.n183 10.6151
R607 B.n185 B.n184 10.6151
R608 B.n185 B.n100 10.6151
R609 B.n189 B.n100 10.6151
R610 B.n190 B.n189 10.6151
R611 B.n191 B.n190 10.6151
R612 B.n191 B.n98 10.6151
R613 B.n195 B.n98 10.6151
R614 B.n196 B.n195 10.6151
R615 B.n198 B.n94 10.6151
R616 B.n202 B.n94 10.6151
R617 B.n203 B.n202 10.6151
R618 B.n204 B.n203 10.6151
R619 B.n204 B.n92 10.6151
R620 B.n208 B.n92 10.6151
R621 B.n209 B.n208 10.6151
R622 B.n210 B.n209 10.6151
R623 B.n214 B.n213 10.6151
R624 B.n215 B.n214 10.6151
R625 B.n215 B.n86 10.6151
R626 B.n219 B.n86 10.6151
R627 B.n220 B.n219 10.6151
R628 B.n221 B.n220 10.6151
R629 B.n221 B.n84 10.6151
R630 B.n225 B.n84 10.6151
R631 B.n226 B.n225 10.6151
R632 B.n227 B.n226 10.6151
R633 B.n227 B.n82 10.6151
R634 B.n231 B.n82 10.6151
R635 B.n232 B.n231 10.6151
R636 B.n233 B.n232 10.6151
R637 B.n233 B.n80 10.6151
R638 B.n237 B.n80 10.6151
R639 B.n238 B.n237 10.6151
R640 B.n239 B.n238 10.6151
R641 B.n239 B.n78 10.6151
R642 B.n243 B.n78 10.6151
R643 B.n244 B.n243 10.6151
R644 B.n245 B.n244 10.6151
R645 B.n245 B.n76 10.6151
R646 B.n249 B.n76 10.6151
R647 B.n250 B.n249 10.6151
R648 B.n251 B.n250 10.6151
R649 B.n251 B.n74 10.6151
R650 B.n255 B.n74 10.6151
R651 B.n256 B.n255 10.6151
R652 B.n257 B.n256 10.6151
R653 B.n257 B.n72 10.6151
R654 B.n261 B.n72 10.6151
R655 B.n262 B.n261 10.6151
R656 B.n263 B.n262 10.6151
R657 B.n143 B.n142 10.6151
R658 B.n142 B.n141 10.6151
R659 B.n141 B.n116 10.6151
R660 B.n137 B.n116 10.6151
R661 B.n137 B.n136 10.6151
R662 B.n136 B.n135 10.6151
R663 B.n135 B.n118 10.6151
R664 B.n131 B.n118 10.6151
R665 B.n131 B.n130 10.6151
R666 B.n130 B.n129 10.6151
R667 B.n129 B.n120 10.6151
R668 B.n125 B.n120 10.6151
R669 B.n125 B.n124 10.6151
R670 B.n124 B.n123 10.6151
R671 B.n123 B.n0 10.6151
R672 B.n455 B.n1 10.6151
R673 B.n455 B.n454 10.6151
R674 B.n454 B.n453 10.6151
R675 B.n453 B.n4 10.6151
R676 B.n449 B.n4 10.6151
R677 B.n449 B.n448 10.6151
R678 B.n448 B.n447 10.6151
R679 B.n447 B.n6 10.6151
R680 B.n443 B.n6 10.6151
R681 B.n443 B.n442 10.6151
R682 B.n442 B.n441 10.6151
R683 B.n441 B.n8 10.6151
R684 B.n437 B.n8 10.6151
R685 B.n437 B.n436 10.6151
R686 B.n436 B.n435 10.6151
R687 B.n381 B.n380 6.5566
R688 B.n368 B.n36 6.5566
R689 B.n198 B.n197 6.5566
R690 B.n210 B.n90 6.5566
R691 B.n382 B.n381 4.05904
R692 B.n365 B.n36 4.05904
R693 B.n197 B.n196 4.05904
R694 B.n213 B.n90 4.05904
R695 B.n459 B.n0 2.81026
R696 B.n459 B.n1 2.81026
R697 VP.n7 VP.t3 1710.73
R698 VP.n5 VP.t5 1710.73
R699 VP.n0 VP.t4 1710.73
R700 VP.n2 VP.t2 1710.73
R701 VP.n6 VP.t0 1650.85
R702 VP.n1 VP.t1 1650.85
R703 VP.n3 VP.n0 161.489
R704 VP.n8 VP.n7 161.3
R705 VP.n3 VP.n2 161.3
R706 VP.n5 VP.n4 161.3
R707 VP.n4 VP.n3 38.1672
R708 VP.n6 VP.n5 36.5157
R709 VP.n7 VP.n6 36.5157
R710 VP.n1 VP.n0 36.5157
R711 VP.n2 VP.n1 36.5157
R712 VP.n8 VP.n4 0.189894
R713 VP VP.n8 0.0516364
R714 VDD1 VDD1.t2 84.3786
R715 VDD1.n1 VDD1.t0 84.2649
R716 VDD1.n1 VDD1.n0 78.8767
R717 VDD1.n3 VDD1.n2 78.7899
R718 VDD1.n3 VDD1.n1 34.7509
R719 VDD1.n2 VDD1.t1 5.10413
R720 VDD1.n2 VDD1.t4 5.10413
R721 VDD1.n0 VDD1.t3 5.10413
R722 VDD1.n0 VDD1.t5 5.10413
R723 VDD1 VDD1.n3 0.0845517
R724 VTAIL.n7 VTAIL.t5 67.2149
R725 VTAIL.n11 VTAIL.t0 67.2147
R726 VTAIL.n2 VTAIL.t8 67.2147
R727 VTAIL.n10 VTAIL.t9 67.2147
R728 VTAIL.n9 VTAIL.n8 62.1113
R729 VTAIL.n6 VTAIL.n5 62.1113
R730 VTAIL.n1 VTAIL.n0 62.111
R731 VTAIL.n4 VTAIL.n3 62.111
R732 VTAIL.n6 VTAIL.n4 21.8238
R733 VTAIL.n11 VTAIL.n10 21.2548
R734 VTAIL.n0 VTAIL.t2 5.10413
R735 VTAIL.n0 VTAIL.t4 5.10413
R736 VTAIL.n3 VTAIL.t6 5.10413
R737 VTAIL.n3 VTAIL.t11 5.10413
R738 VTAIL.n8 VTAIL.t7 5.10413
R739 VTAIL.n8 VTAIL.t10 5.10413
R740 VTAIL.n5 VTAIL.t3 5.10413
R741 VTAIL.n5 VTAIL.t1 5.10413
R742 VTAIL.n9 VTAIL.n7 0.75481
R743 VTAIL.n2 VTAIL.n1 0.75481
R744 VTAIL.n7 VTAIL.n6 0.569465
R745 VTAIL.n10 VTAIL.n9 0.569465
R746 VTAIL.n4 VTAIL.n2 0.569465
R747 VTAIL VTAIL.n11 0.369034
R748 VTAIL VTAIL.n1 0.200931
R749 VN.n2 VN.t5 1710.73
R750 VN.n0 VN.t3 1710.73
R751 VN.n6 VN.t0 1710.73
R752 VN.n4 VN.t2 1710.73
R753 VN.n1 VN.t1 1650.85
R754 VN.n5 VN.t4 1650.85
R755 VN.n7 VN.n4 161.489
R756 VN.n3 VN.n0 161.489
R757 VN.n3 VN.n2 161.3
R758 VN.n7 VN.n6 161.3
R759 VN VN.n7 38.5478
R760 VN.n1 VN.n0 36.5157
R761 VN.n2 VN.n1 36.5157
R762 VN.n6 VN.n5 36.5157
R763 VN.n5 VN.n4 36.5157
R764 VN VN.n3 0.0516364
R765 VDD2.n1 VDD2.t2 84.2649
R766 VDD2.n2 VDD2.t5 83.8936
R767 VDD2.n1 VDD2.n0 78.8767
R768 VDD2 VDD2.n3 78.874
R769 VDD2.n2 VDD2.n1 33.8834
R770 VDD2.n3 VDD2.t1 5.10413
R771 VDD2.n3 VDD2.t3 5.10413
R772 VDD2.n0 VDD2.t4 5.10413
R773 VDD2.n0 VDD2.t0 5.10413
R774 VDD2 VDD2.n2 0.485414
C0 VP w_n1498_n2898# 2.34906f
C1 VTAIL w_n1498_n2898# 2.63526f
C2 VN B 0.639703f
C3 VTAIL VP 1.13737f
C4 VDD1 w_n1498_n2898# 1.5316f
C5 VDD1 VP 1.68161f
C6 VDD2 B 1.29897f
C7 VDD1 VTAIL 11.5976f
C8 VDD2 VN 1.56724f
C9 B w_n1498_n2898# 5.88162f
C10 VN w_n1498_n2898# 2.16171f
C11 VP B 0.941018f
C12 VTAIL B 2.04167f
C13 VN VP 4.2687f
C14 VDD1 B 1.2782f
C15 VTAIL VN 1.12275f
C16 VDD2 w_n1498_n2898# 1.54454f
C17 VDD1 VN 0.147253f
C18 VDD2 VP 0.265626f
C19 VDD2 VTAIL 11.6291f
C20 VDD2 VDD1 0.57916f
C21 VDD2 VSUBS 1.09585f
C22 VDD1 VSUBS 1.362375f
C23 VTAIL VSUBS 0.537181f
C24 VN VSUBS 3.57723f
C25 VP VSUBS 0.984024f
C26 B VSUBS 2.102756f
C27 w_n1498_n2898# VSUBS 53.658398f
C28 VDD2.t2 VSUBS 1.73491f
C29 VDD2.t4 VSUBS 0.245894f
C30 VDD2.t0 VSUBS 0.245894f
C31 VDD2.n0 VSUBS 1.38685f
C32 VDD2.n1 VSUBS 1.96411f
C33 VDD2.t5 VSUBS 1.73267f
C34 VDD2.n2 VSUBS 1.93994f
C35 VDD2.t1 VSUBS 0.245894f
C36 VDD2.t3 VSUBS 0.245894f
C37 VDD2.n3 VSUBS 1.38682f
C38 VN.t3 VSUBS 0.251689f
C39 VN.n0 VSUBS 0.133227f
C40 VN.t1 VSUBS 0.247743f
C41 VN.n1 VSUBS 0.110261f
C42 VN.t5 VSUBS 0.251689f
C43 VN.n2 VSUBS 0.133141f
C44 VN.n3 VSUBS 0.117227f
C45 VN.t2 VSUBS 0.251689f
C46 VN.n4 VSUBS 0.133227f
C47 VN.t0 VSUBS 0.251689f
C48 VN.t4 VSUBS 0.247743f
C49 VN.n5 VSUBS 0.110261f
C50 VN.n6 VSUBS 0.133141f
C51 VN.n7 VSUBS 2.09318f
C52 VTAIL.t2 VSUBS 0.313253f
C53 VTAIL.t4 VSUBS 0.313253f
C54 VTAIL.n0 VSUBS 1.63779f
C55 VTAIL.n1 VSUBS 0.657988f
C56 VTAIL.t8 VSUBS 2.05826f
C57 VTAIL.n2 VSUBS 0.833574f
C58 VTAIL.t6 VSUBS 0.313253f
C59 VTAIL.t11 VSUBS 0.313253f
C60 VTAIL.n3 VSUBS 1.63779f
C61 VTAIL.n4 VSUBS 1.81872f
C62 VTAIL.t3 VSUBS 0.313253f
C63 VTAIL.t1 VSUBS 0.313253f
C64 VTAIL.n5 VSUBS 1.6378f
C65 VTAIL.n6 VSUBS 1.81872f
C66 VTAIL.t5 VSUBS 2.05827f
C67 VTAIL.n7 VSUBS 0.833561f
C68 VTAIL.t7 VSUBS 0.313253f
C69 VTAIL.t10 VSUBS 0.313253f
C70 VTAIL.n8 VSUBS 1.6378f
C71 VTAIL.n9 VSUBS 0.690177f
C72 VTAIL.t9 VSUBS 2.05826f
C73 VTAIL.n10 VSUBS 1.91241f
C74 VTAIL.t0 VSUBS 2.05826f
C75 VTAIL.n11 VSUBS 1.8949f
C76 VDD1.t2 VSUBS 1.72396f
C77 VDD1.t0 VSUBS 1.72324f
C78 VDD1.t3 VSUBS 0.244239f
C79 VDD1.t5 VSUBS 0.244239f
C80 VDD1.n0 VSUBS 1.37751f
C81 VDD1.n1 VSUBS 2.0085f
C82 VDD1.t1 VSUBS 0.244239f
C83 VDD1.t4 VSUBS 0.244239f
C84 VDD1.n2 VSUBS 1.37703f
C85 VDD1.n3 VSUBS 1.86315f
C86 VP.t4 VSUBS 0.25873f
C87 VP.n0 VSUBS 0.136954f
C88 VP.t1 VSUBS 0.254675f
C89 VP.n1 VSUBS 0.113346f
C90 VP.t2 VSUBS 0.25873f
C91 VP.n2 VSUBS 0.136866f
C92 VP.n3 VSUBS 2.11328f
C93 VP.n4 VSUBS 2.09274f
C94 VP.t0 VSUBS 0.254675f
C95 VP.t5 VSUBS 0.25873f
C96 VP.n5 VSUBS 0.136866f
C97 VP.n6 VSUBS 0.113346f
C98 VP.t3 VSUBS 0.25873f
C99 VP.n7 VSUBS 0.136866f
C100 VP.n8 VSUBS 0.045129f
C101 B.n0 VSUBS 0.005044f
C102 B.n1 VSUBS 0.005044f
C103 B.n2 VSUBS 0.007977f
C104 B.n3 VSUBS 0.007977f
C105 B.n4 VSUBS 0.007977f
C106 B.n5 VSUBS 0.007977f
C107 B.n6 VSUBS 0.007977f
C108 B.n7 VSUBS 0.007977f
C109 B.n8 VSUBS 0.007977f
C110 B.n9 VSUBS 0.007977f
C111 B.n10 VSUBS 0.01844f
C112 B.n11 VSUBS 0.007977f
C113 B.n12 VSUBS 0.007977f
C114 B.n13 VSUBS 0.007977f
C115 B.n14 VSUBS 0.007977f
C116 B.n15 VSUBS 0.007977f
C117 B.n16 VSUBS 0.007977f
C118 B.n17 VSUBS 0.007977f
C119 B.n18 VSUBS 0.007977f
C120 B.n19 VSUBS 0.007977f
C121 B.n20 VSUBS 0.007977f
C122 B.n21 VSUBS 0.007977f
C123 B.n22 VSUBS 0.007977f
C124 B.n23 VSUBS 0.007977f
C125 B.n24 VSUBS 0.007977f
C126 B.n25 VSUBS 0.007977f
C127 B.n26 VSUBS 0.007977f
C128 B.n27 VSUBS 0.007977f
C129 B.t5 VSUBS 0.390222f
C130 B.t4 VSUBS 0.396912f
C131 B.t3 VSUBS 0.068098f
C132 B.n28 VSUBS 0.091287f
C133 B.n29 VSUBS 0.076636f
C134 B.n30 VSUBS 0.007977f
C135 B.n31 VSUBS 0.007977f
C136 B.n32 VSUBS 0.007977f
C137 B.n33 VSUBS 0.007977f
C138 B.t2 VSUBS 0.390218f
C139 B.t1 VSUBS 0.396908f
C140 B.t0 VSUBS 0.068098f
C141 B.n34 VSUBS 0.091291f
C142 B.n35 VSUBS 0.07664f
C143 B.n36 VSUBS 0.018482f
C144 B.n37 VSUBS 0.007977f
C145 B.n38 VSUBS 0.007977f
C146 B.n39 VSUBS 0.007977f
C147 B.n40 VSUBS 0.007977f
C148 B.n41 VSUBS 0.007977f
C149 B.n42 VSUBS 0.007977f
C150 B.n43 VSUBS 0.007977f
C151 B.n44 VSUBS 0.007977f
C152 B.n45 VSUBS 0.007977f
C153 B.n46 VSUBS 0.007977f
C154 B.n47 VSUBS 0.007977f
C155 B.n48 VSUBS 0.007977f
C156 B.n49 VSUBS 0.007977f
C157 B.n50 VSUBS 0.007977f
C158 B.n51 VSUBS 0.007977f
C159 B.n52 VSUBS 0.007977f
C160 B.n53 VSUBS 0.007977f
C161 B.n54 VSUBS 0.018682f
C162 B.n55 VSUBS 0.007977f
C163 B.n56 VSUBS 0.007977f
C164 B.n57 VSUBS 0.007977f
C165 B.n58 VSUBS 0.007977f
C166 B.n59 VSUBS 0.007977f
C167 B.n60 VSUBS 0.007977f
C168 B.n61 VSUBS 0.007977f
C169 B.n62 VSUBS 0.007977f
C170 B.n63 VSUBS 0.007977f
C171 B.n64 VSUBS 0.007977f
C172 B.n65 VSUBS 0.007977f
C173 B.n66 VSUBS 0.007977f
C174 B.n67 VSUBS 0.007977f
C175 B.n68 VSUBS 0.007977f
C176 B.n69 VSUBS 0.007977f
C177 B.n70 VSUBS 0.017691f
C178 B.n71 VSUBS 0.007977f
C179 B.n72 VSUBS 0.007977f
C180 B.n73 VSUBS 0.007977f
C181 B.n74 VSUBS 0.007977f
C182 B.n75 VSUBS 0.007977f
C183 B.n76 VSUBS 0.007977f
C184 B.n77 VSUBS 0.007977f
C185 B.n78 VSUBS 0.007977f
C186 B.n79 VSUBS 0.007977f
C187 B.n80 VSUBS 0.007977f
C188 B.n81 VSUBS 0.007977f
C189 B.n82 VSUBS 0.007977f
C190 B.n83 VSUBS 0.007977f
C191 B.n84 VSUBS 0.007977f
C192 B.n85 VSUBS 0.007977f
C193 B.n86 VSUBS 0.007977f
C194 B.n87 VSUBS 0.007977f
C195 B.t7 VSUBS 0.390218f
C196 B.t8 VSUBS 0.396908f
C197 B.t6 VSUBS 0.068098f
C198 B.n88 VSUBS 0.091291f
C199 B.n89 VSUBS 0.07664f
C200 B.n90 VSUBS 0.018482f
C201 B.n91 VSUBS 0.007977f
C202 B.n92 VSUBS 0.007977f
C203 B.n93 VSUBS 0.007977f
C204 B.n94 VSUBS 0.007977f
C205 B.n95 VSUBS 0.007977f
C206 B.t10 VSUBS 0.390222f
C207 B.t11 VSUBS 0.396912f
C208 B.t9 VSUBS 0.068098f
C209 B.n96 VSUBS 0.091287f
C210 B.n97 VSUBS 0.076636f
C211 B.n98 VSUBS 0.007977f
C212 B.n99 VSUBS 0.007977f
C213 B.n100 VSUBS 0.007977f
C214 B.n101 VSUBS 0.007977f
C215 B.n102 VSUBS 0.007977f
C216 B.n103 VSUBS 0.007977f
C217 B.n104 VSUBS 0.007977f
C218 B.n105 VSUBS 0.007977f
C219 B.n106 VSUBS 0.007977f
C220 B.n107 VSUBS 0.007977f
C221 B.n108 VSUBS 0.007977f
C222 B.n109 VSUBS 0.007977f
C223 B.n110 VSUBS 0.007977f
C224 B.n111 VSUBS 0.007977f
C225 B.n112 VSUBS 0.007977f
C226 B.n113 VSUBS 0.007977f
C227 B.n114 VSUBS 0.01844f
C228 B.n115 VSUBS 0.007977f
C229 B.n116 VSUBS 0.007977f
C230 B.n117 VSUBS 0.007977f
C231 B.n118 VSUBS 0.007977f
C232 B.n119 VSUBS 0.007977f
C233 B.n120 VSUBS 0.007977f
C234 B.n121 VSUBS 0.007977f
C235 B.n122 VSUBS 0.007977f
C236 B.n123 VSUBS 0.007977f
C237 B.n124 VSUBS 0.007977f
C238 B.n125 VSUBS 0.007977f
C239 B.n126 VSUBS 0.007977f
C240 B.n127 VSUBS 0.007977f
C241 B.n128 VSUBS 0.007977f
C242 B.n129 VSUBS 0.007977f
C243 B.n130 VSUBS 0.007977f
C244 B.n131 VSUBS 0.007977f
C245 B.n132 VSUBS 0.007977f
C246 B.n133 VSUBS 0.007977f
C247 B.n134 VSUBS 0.007977f
C248 B.n135 VSUBS 0.007977f
C249 B.n136 VSUBS 0.007977f
C250 B.n137 VSUBS 0.007977f
C251 B.n138 VSUBS 0.007977f
C252 B.n139 VSUBS 0.007977f
C253 B.n140 VSUBS 0.007977f
C254 B.n141 VSUBS 0.007977f
C255 B.n142 VSUBS 0.007977f
C256 B.n143 VSUBS 0.017691f
C257 B.n144 VSUBS 0.017691f
C258 B.n145 VSUBS 0.01844f
C259 B.n146 VSUBS 0.007977f
C260 B.n147 VSUBS 0.007977f
C261 B.n148 VSUBS 0.007977f
C262 B.n149 VSUBS 0.007977f
C263 B.n150 VSUBS 0.007977f
C264 B.n151 VSUBS 0.007977f
C265 B.n152 VSUBS 0.007977f
C266 B.n153 VSUBS 0.007977f
C267 B.n154 VSUBS 0.007977f
C268 B.n155 VSUBS 0.007977f
C269 B.n156 VSUBS 0.007977f
C270 B.n157 VSUBS 0.007977f
C271 B.n158 VSUBS 0.007977f
C272 B.n159 VSUBS 0.007977f
C273 B.n160 VSUBS 0.007977f
C274 B.n161 VSUBS 0.007977f
C275 B.n162 VSUBS 0.007977f
C276 B.n163 VSUBS 0.007977f
C277 B.n164 VSUBS 0.007977f
C278 B.n165 VSUBS 0.007977f
C279 B.n166 VSUBS 0.007977f
C280 B.n167 VSUBS 0.007977f
C281 B.n168 VSUBS 0.007977f
C282 B.n169 VSUBS 0.007977f
C283 B.n170 VSUBS 0.007977f
C284 B.n171 VSUBS 0.007977f
C285 B.n172 VSUBS 0.007977f
C286 B.n173 VSUBS 0.007977f
C287 B.n174 VSUBS 0.007977f
C288 B.n175 VSUBS 0.007977f
C289 B.n176 VSUBS 0.007977f
C290 B.n177 VSUBS 0.007977f
C291 B.n178 VSUBS 0.007977f
C292 B.n179 VSUBS 0.007977f
C293 B.n180 VSUBS 0.007977f
C294 B.n181 VSUBS 0.007977f
C295 B.n182 VSUBS 0.007977f
C296 B.n183 VSUBS 0.007977f
C297 B.n184 VSUBS 0.007977f
C298 B.n185 VSUBS 0.007977f
C299 B.n186 VSUBS 0.007977f
C300 B.n187 VSUBS 0.007977f
C301 B.n188 VSUBS 0.007977f
C302 B.n189 VSUBS 0.007977f
C303 B.n190 VSUBS 0.007977f
C304 B.n191 VSUBS 0.007977f
C305 B.n192 VSUBS 0.007977f
C306 B.n193 VSUBS 0.007977f
C307 B.n194 VSUBS 0.007977f
C308 B.n195 VSUBS 0.007977f
C309 B.n196 VSUBS 0.005514f
C310 B.n197 VSUBS 0.018482f
C311 B.n198 VSUBS 0.006452f
C312 B.n199 VSUBS 0.007977f
C313 B.n200 VSUBS 0.007977f
C314 B.n201 VSUBS 0.007977f
C315 B.n202 VSUBS 0.007977f
C316 B.n203 VSUBS 0.007977f
C317 B.n204 VSUBS 0.007977f
C318 B.n205 VSUBS 0.007977f
C319 B.n206 VSUBS 0.007977f
C320 B.n207 VSUBS 0.007977f
C321 B.n208 VSUBS 0.007977f
C322 B.n209 VSUBS 0.007977f
C323 B.n210 VSUBS 0.006452f
C324 B.n211 VSUBS 0.007977f
C325 B.n212 VSUBS 0.007977f
C326 B.n213 VSUBS 0.005514f
C327 B.n214 VSUBS 0.007977f
C328 B.n215 VSUBS 0.007977f
C329 B.n216 VSUBS 0.007977f
C330 B.n217 VSUBS 0.007977f
C331 B.n218 VSUBS 0.007977f
C332 B.n219 VSUBS 0.007977f
C333 B.n220 VSUBS 0.007977f
C334 B.n221 VSUBS 0.007977f
C335 B.n222 VSUBS 0.007977f
C336 B.n223 VSUBS 0.007977f
C337 B.n224 VSUBS 0.007977f
C338 B.n225 VSUBS 0.007977f
C339 B.n226 VSUBS 0.007977f
C340 B.n227 VSUBS 0.007977f
C341 B.n228 VSUBS 0.007977f
C342 B.n229 VSUBS 0.007977f
C343 B.n230 VSUBS 0.007977f
C344 B.n231 VSUBS 0.007977f
C345 B.n232 VSUBS 0.007977f
C346 B.n233 VSUBS 0.007977f
C347 B.n234 VSUBS 0.007977f
C348 B.n235 VSUBS 0.007977f
C349 B.n236 VSUBS 0.007977f
C350 B.n237 VSUBS 0.007977f
C351 B.n238 VSUBS 0.007977f
C352 B.n239 VSUBS 0.007977f
C353 B.n240 VSUBS 0.007977f
C354 B.n241 VSUBS 0.007977f
C355 B.n242 VSUBS 0.007977f
C356 B.n243 VSUBS 0.007977f
C357 B.n244 VSUBS 0.007977f
C358 B.n245 VSUBS 0.007977f
C359 B.n246 VSUBS 0.007977f
C360 B.n247 VSUBS 0.007977f
C361 B.n248 VSUBS 0.007977f
C362 B.n249 VSUBS 0.007977f
C363 B.n250 VSUBS 0.007977f
C364 B.n251 VSUBS 0.007977f
C365 B.n252 VSUBS 0.007977f
C366 B.n253 VSUBS 0.007977f
C367 B.n254 VSUBS 0.007977f
C368 B.n255 VSUBS 0.007977f
C369 B.n256 VSUBS 0.007977f
C370 B.n257 VSUBS 0.007977f
C371 B.n258 VSUBS 0.007977f
C372 B.n259 VSUBS 0.007977f
C373 B.n260 VSUBS 0.007977f
C374 B.n261 VSUBS 0.007977f
C375 B.n262 VSUBS 0.007977f
C376 B.n263 VSUBS 0.01844f
C377 B.n264 VSUBS 0.01844f
C378 B.n265 VSUBS 0.017691f
C379 B.n266 VSUBS 0.007977f
C380 B.n267 VSUBS 0.007977f
C381 B.n268 VSUBS 0.007977f
C382 B.n269 VSUBS 0.007977f
C383 B.n270 VSUBS 0.007977f
C384 B.n271 VSUBS 0.007977f
C385 B.n272 VSUBS 0.007977f
C386 B.n273 VSUBS 0.007977f
C387 B.n274 VSUBS 0.007977f
C388 B.n275 VSUBS 0.007977f
C389 B.n276 VSUBS 0.007977f
C390 B.n277 VSUBS 0.007977f
C391 B.n278 VSUBS 0.007977f
C392 B.n279 VSUBS 0.007977f
C393 B.n280 VSUBS 0.007977f
C394 B.n281 VSUBS 0.007977f
C395 B.n282 VSUBS 0.007977f
C396 B.n283 VSUBS 0.007977f
C397 B.n284 VSUBS 0.007977f
C398 B.n285 VSUBS 0.007977f
C399 B.n286 VSUBS 0.007977f
C400 B.n287 VSUBS 0.007977f
C401 B.n288 VSUBS 0.007977f
C402 B.n289 VSUBS 0.007977f
C403 B.n290 VSUBS 0.007977f
C404 B.n291 VSUBS 0.007977f
C405 B.n292 VSUBS 0.007977f
C406 B.n293 VSUBS 0.007977f
C407 B.n294 VSUBS 0.007977f
C408 B.n295 VSUBS 0.007977f
C409 B.n296 VSUBS 0.007977f
C410 B.n297 VSUBS 0.007977f
C411 B.n298 VSUBS 0.007977f
C412 B.n299 VSUBS 0.007977f
C413 B.n300 VSUBS 0.007977f
C414 B.n301 VSUBS 0.007977f
C415 B.n302 VSUBS 0.007977f
C416 B.n303 VSUBS 0.007977f
C417 B.n304 VSUBS 0.007977f
C418 B.n305 VSUBS 0.007977f
C419 B.n306 VSUBS 0.007977f
C420 B.n307 VSUBS 0.007977f
C421 B.n308 VSUBS 0.007977f
C422 B.n309 VSUBS 0.007977f
C423 B.n310 VSUBS 0.007977f
C424 B.n311 VSUBS 0.007977f
C425 B.n312 VSUBS 0.007977f
C426 B.n313 VSUBS 0.017691f
C427 B.n314 VSUBS 0.01844f
C428 B.n315 VSUBS 0.017449f
C429 B.n316 VSUBS 0.007977f
C430 B.n317 VSUBS 0.007977f
C431 B.n318 VSUBS 0.007977f
C432 B.n319 VSUBS 0.007977f
C433 B.n320 VSUBS 0.007977f
C434 B.n321 VSUBS 0.007977f
C435 B.n322 VSUBS 0.007977f
C436 B.n323 VSUBS 0.007977f
C437 B.n324 VSUBS 0.007977f
C438 B.n325 VSUBS 0.007977f
C439 B.n326 VSUBS 0.007977f
C440 B.n327 VSUBS 0.007977f
C441 B.n328 VSUBS 0.007977f
C442 B.n329 VSUBS 0.007977f
C443 B.n330 VSUBS 0.007977f
C444 B.n331 VSUBS 0.007977f
C445 B.n332 VSUBS 0.007977f
C446 B.n333 VSUBS 0.007977f
C447 B.n334 VSUBS 0.007977f
C448 B.n335 VSUBS 0.007977f
C449 B.n336 VSUBS 0.007977f
C450 B.n337 VSUBS 0.007977f
C451 B.n338 VSUBS 0.007977f
C452 B.n339 VSUBS 0.007977f
C453 B.n340 VSUBS 0.007977f
C454 B.n341 VSUBS 0.007977f
C455 B.n342 VSUBS 0.007977f
C456 B.n343 VSUBS 0.007977f
C457 B.n344 VSUBS 0.007977f
C458 B.n345 VSUBS 0.007977f
C459 B.n346 VSUBS 0.007977f
C460 B.n347 VSUBS 0.007977f
C461 B.n348 VSUBS 0.007977f
C462 B.n349 VSUBS 0.007977f
C463 B.n350 VSUBS 0.007977f
C464 B.n351 VSUBS 0.007977f
C465 B.n352 VSUBS 0.007977f
C466 B.n353 VSUBS 0.007977f
C467 B.n354 VSUBS 0.007977f
C468 B.n355 VSUBS 0.007977f
C469 B.n356 VSUBS 0.007977f
C470 B.n357 VSUBS 0.007977f
C471 B.n358 VSUBS 0.007977f
C472 B.n359 VSUBS 0.007977f
C473 B.n360 VSUBS 0.007977f
C474 B.n361 VSUBS 0.007977f
C475 B.n362 VSUBS 0.007977f
C476 B.n363 VSUBS 0.007977f
C477 B.n364 VSUBS 0.007977f
C478 B.n365 VSUBS 0.005514f
C479 B.n366 VSUBS 0.007977f
C480 B.n367 VSUBS 0.007977f
C481 B.n368 VSUBS 0.006452f
C482 B.n369 VSUBS 0.007977f
C483 B.n370 VSUBS 0.007977f
C484 B.n371 VSUBS 0.007977f
C485 B.n372 VSUBS 0.007977f
C486 B.n373 VSUBS 0.007977f
C487 B.n374 VSUBS 0.007977f
C488 B.n375 VSUBS 0.007977f
C489 B.n376 VSUBS 0.007977f
C490 B.n377 VSUBS 0.007977f
C491 B.n378 VSUBS 0.007977f
C492 B.n379 VSUBS 0.007977f
C493 B.n380 VSUBS 0.006452f
C494 B.n381 VSUBS 0.018482f
C495 B.n382 VSUBS 0.005514f
C496 B.n383 VSUBS 0.007977f
C497 B.n384 VSUBS 0.007977f
C498 B.n385 VSUBS 0.007977f
C499 B.n386 VSUBS 0.007977f
C500 B.n387 VSUBS 0.007977f
C501 B.n388 VSUBS 0.007977f
C502 B.n389 VSUBS 0.007977f
C503 B.n390 VSUBS 0.007977f
C504 B.n391 VSUBS 0.007977f
C505 B.n392 VSUBS 0.007977f
C506 B.n393 VSUBS 0.007977f
C507 B.n394 VSUBS 0.007977f
C508 B.n395 VSUBS 0.007977f
C509 B.n396 VSUBS 0.007977f
C510 B.n397 VSUBS 0.007977f
C511 B.n398 VSUBS 0.007977f
C512 B.n399 VSUBS 0.007977f
C513 B.n400 VSUBS 0.007977f
C514 B.n401 VSUBS 0.007977f
C515 B.n402 VSUBS 0.007977f
C516 B.n403 VSUBS 0.007977f
C517 B.n404 VSUBS 0.007977f
C518 B.n405 VSUBS 0.007977f
C519 B.n406 VSUBS 0.007977f
C520 B.n407 VSUBS 0.007977f
C521 B.n408 VSUBS 0.007977f
C522 B.n409 VSUBS 0.007977f
C523 B.n410 VSUBS 0.007977f
C524 B.n411 VSUBS 0.007977f
C525 B.n412 VSUBS 0.007977f
C526 B.n413 VSUBS 0.007977f
C527 B.n414 VSUBS 0.007977f
C528 B.n415 VSUBS 0.007977f
C529 B.n416 VSUBS 0.007977f
C530 B.n417 VSUBS 0.007977f
C531 B.n418 VSUBS 0.007977f
C532 B.n419 VSUBS 0.007977f
C533 B.n420 VSUBS 0.007977f
C534 B.n421 VSUBS 0.007977f
C535 B.n422 VSUBS 0.007977f
C536 B.n423 VSUBS 0.007977f
C537 B.n424 VSUBS 0.007977f
C538 B.n425 VSUBS 0.007977f
C539 B.n426 VSUBS 0.007977f
C540 B.n427 VSUBS 0.007977f
C541 B.n428 VSUBS 0.007977f
C542 B.n429 VSUBS 0.007977f
C543 B.n430 VSUBS 0.007977f
C544 B.n431 VSUBS 0.007977f
C545 B.n432 VSUBS 0.007977f
C546 B.n433 VSUBS 0.01844f
C547 B.n434 VSUBS 0.017691f
C548 B.n435 VSUBS 0.017691f
C549 B.n436 VSUBS 0.007977f
C550 B.n437 VSUBS 0.007977f
C551 B.n438 VSUBS 0.007977f
C552 B.n439 VSUBS 0.007977f
C553 B.n440 VSUBS 0.007977f
C554 B.n441 VSUBS 0.007977f
C555 B.n442 VSUBS 0.007977f
C556 B.n443 VSUBS 0.007977f
C557 B.n444 VSUBS 0.007977f
C558 B.n445 VSUBS 0.007977f
C559 B.n446 VSUBS 0.007977f
C560 B.n447 VSUBS 0.007977f
C561 B.n448 VSUBS 0.007977f
C562 B.n449 VSUBS 0.007977f
C563 B.n450 VSUBS 0.007977f
C564 B.n451 VSUBS 0.007977f
C565 B.n452 VSUBS 0.007977f
C566 B.n453 VSUBS 0.007977f
C567 B.n454 VSUBS 0.007977f
C568 B.n455 VSUBS 0.007977f
C569 B.n456 VSUBS 0.007977f
C570 B.n457 VSUBS 0.007977f
C571 B.n458 VSUBS 0.007977f
C572 B.n459 VSUBS 0.018063f
.ends

