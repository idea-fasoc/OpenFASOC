* NGSPICE file created from diff_pair_sample_0347.ext - technology: sky130A

.subckt diff_pair_sample_0347 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=7.0512 ps=36.94 w=18.08 l=2.45
X1 VDD1.t4 VP.t1 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=2.9832 ps=18.41 w=18.08 l=2.45
X2 VDD1.t3 VP.t2 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=7.0512 ps=36.94 w=18.08 l=2.45
X3 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=2.9832 ps=18.41 w=18.08 l=2.45
X4 VDD1.t2 VP.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=2.9832 ps=18.41 w=18.08 l=2.45
X5 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=7.0512 ps=36.94 w=18.08 l=2.45
X6 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=0 ps=0 w=18.08 l=2.45
X7 VTAIL.t6 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=2.9832 ps=18.41 w=18.08 l=2.45
X8 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=2.9832 ps=18.41 w=18.08 l=2.45
X9 VTAIL.t9 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=2.9832 ps=18.41 w=18.08 l=2.45
X10 VDD2.t2 VN.t3 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=7.0512 ps=36.94 w=18.08 l=2.45
X11 VTAIL.t10 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=2.9832 ps=18.41 w=18.08 l=2.45
X12 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=0 ps=0 w=18.08 l=2.45
X13 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=0 ps=0 w=18.08 l=2.45
X14 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9832 pd=18.41 as=2.9832 ps=18.41 w=18.08 l=2.45
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0512 pd=36.94 as=0 ps=0 w=18.08 l=2.45
R0 VP.n9 VP.t3 212.732
R1 VP.n30 VP.t5 177.849
R2 VP.n20 VP.t1 177.849
R3 VP.n38 VP.t2 177.849
R4 VP.n10 VP.t4 177.849
R5 VP.n18 VP.t0 177.849
R6 VP.n11 VP.n8 161.3
R7 VP.n13 VP.n12 161.3
R8 VP.n14 VP.n7 161.3
R9 VP.n16 VP.n15 161.3
R10 VP.n17 VP.n6 161.3
R11 VP.n37 VP.n0 161.3
R12 VP.n36 VP.n35 161.3
R13 VP.n34 VP.n1 161.3
R14 VP.n33 VP.n32 161.3
R15 VP.n31 VP.n2 161.3
R16 VP.n30 VP.n29 161.3
R17 VP.n28 VP.n3 161.3
R18 VP.n27 VP.n26 161.3
R19 VP.n25 VP.n4 161.3
R20 VP.n24 VP.n23 161.3
R21 VP.n22 VP.n5 161.3
R22 VP.n21 VP.n20 97.1368
R23 VP.n39 VP.n38 97.1368
R24 VP.n19 VP.n18 97.1368
R25 VP.n21 VP.n19 52.7345
R26 VP.n26 VP.n25 51.2335
R27 VP.n32 VP.n1 51.2335
R28 VP.n12 VP.n7 51.2335
R29 VP.n10 VP.n9 48.154
R30 VP.n25 VP.n24 29.9206
R31 VP.n36 VP.n1 29.9206
R32 VP.n16 VP.n7 29.9206
R33 VP.n24 VP.n5 24.5923
R34 VP.n26 VP.n3 24.5923
R35 VP.n30 VP.n3 24.5923
R36 VP.n31 VP.n30 24.5923
R37 VP.n32 VP.n31 24.5923
R38 VP.n37 VP.n36 24.5923
R39 VP.n17 VP.n16 24.5923
R40 VP.n11 VP.n10 24.5923
R41 VP.n12 VP.n11 24.5923
R42 VP.n20 VP.n5 13.7719
R43 VP.n38 VP.n37 13.7719
R44 VP.n18 VP.n17 13.7719
R45 VP.n9 VP.n8 6.57284
R46 VP.n19 VP.n6 0.278335
R47 VP.n22 VP.n21 0.278335
R48 VP.n39 VP.n0 0.278335
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153485
R64 VTAIL.n406 VTAIL.n405 289.615
R65 VTAIL.n100 VTAIL.n99 289.615
R66 VTAIL.n306 VTAIL.n305 289.615
R67 VTAIL.n204 VTAIL.n203 289.615
R68 VTAIL.n341 VTAIL.n340 185
R69 VTAIL.n338 VTAIL.n337 185
R70 VTAIL.n347 VTAIL.n346 185
R71 VTAIL.n349 VTAIL.n348 185
R72 VTAIL.n334 VTAIL.n333 185
R73 VTAIL.n355 VTAIL.n354 185
R74 VTAIL.n358 VTAIL.n357 185
R75 VTAIL.n356 VTAIL.n330 185
R76 VTAIL.n363 VTAIL.n329 185
R77 VTAIL.n365 VTAIL.n364 185
R78 VTAIL.n367 VTAIL.n366 185
R79 VTAIL.n326 VTAIL.n325 185
R80 VTAIL.n373 VTAIL.n372 185
R81 VTAIL.n375 VTAIL.n374 185
R82 VTAIL.n322 VTAIL.n321 185
R83 VTAIL.n381 VTAIL.n380 185
R84 VTAIL.n383 VTAIL.n382 185
R85 VTAIL.n318 VTAIL.n317 185
R86 VTAIL.n389 VTAIL.n388 185
R87 VTAIL.n391 VTAIL.n390 185
R88 VTAIL.n314 VTAIL.n313 185
R89 VTAIL.n397 VTAIL.n396 185
R90 VTAIL.n399 VTAIL.n398 185
R91 VTAIL.n310 VTAIL.n309 185
R92 VTAIL.n405 VTAIL.n404 185
R93 VTAIL.n35 VTAIL.n34 185
R94 VTAIL.n32 VTAIL.n31 185
R95 VTAIL.n41 VTAIL.n40 185
R96 VTAIL.n43 VTAIL.n42 185
R97 VTAIL.n28 VTAIL.n27 185
R98 VTAIL.n49 VTAIL.n48 185
R99 VTAIL.n52 VTAIL.n51 185
R100 VTAIL.n50 VTAIL.n24 185
R101 VTAIL.n57 VTAIL.n23 185
R102 VTAIL.n59 VTAIL.n58 185
R103 VTAIL.n61 VTAIL.n60 185
R104 VTAIL.n20 VTAIL.n19 185
R105 VTAIL.n67 VTAIL.n66 185
R106 VTAIL.n69 VTAIL.n68 185
R107 VTAIL.n16 VTAIL.n15 185
R108 VTAIL.n75 VTAIL.n74 185
R109 VTAIL.n77 VTAIL.n76 185
R110 VTAIL.n12 VTAIL.n11 185
R111 VTAIL.n83 VTAIL.n82 185
R112 VTAIL.n85 VTAIL.n84 185
R113 VTAIL.n8 VTAIL.n7 185
R114 VTAIL.n91 VTAIL.n90 185
R115 VTAIL.n93 VTAIL.n92 185
R116 VTAIL.n4 VTAIL.n3 185
R117 VTAIL.n99 VTAIL.n98 185
R118 VTAIL.n305 VTAIL.n304 185
R119 VTAIL.n210 VTAIL.n209 185
R120 VTAIL.n299 VTAIL.n298 185
R121 VTAIL.n297 VTAIL.n296 185
R122 VTAIL.n214 VTAIL.n213 185
R123 VTAIL.n291 VTAIL.n290 185
R124 VTAIL.n289 VTAIL.n288 185
R125 VTAIL.n218 VTAIL.n217 185
R126 VTAIL.n283 VTAIL.n282 185
R127 VTAIL.n281 VTAIL.n280 185
R128 VTAIL.n222 VTAIL.n221 185
R129 VTAIL.n275 VTAIL.n274 185
R130 VTAIL.n273 VTAIL.n272 185
R131 VTAIL.n226 VTAIL.n225 185
R132 VTAIL.n267 VTAIL.n266 185
R133 VTAIL.n265 VTAIL.n264 185
R134 VTAIL.n263 VTAIL.n229 185
R135 VTAIL.n233 VTAIL.n230 185
R136 VTAIL.n258 VTAIL.n257 185
R137 VTAIL.n256 VTAIL.n255 185
R138 VTAIL.n235 VTAIL.n234 185
R139 VTAIL.n250 VTAIL.n249 185
R140 VTAIL.n248 VTAIL.n247 185
R141 VTAIL.n239 VTAIL.n238 185
R142 VTAIL.n242 VTAIL.n241 185
R143 VTAIL.n203 VTAIL.n202 185
R144 VTAIL.n108 VTAIL.n107 185
R145 VTAIL.n197 VTAIL.n196 185
R146 VTAIL.n195 VTAIL.n194 185
R147 VTAIL.n112 VTAIL.n111 185
R148 VTAIL.n189 VTAIL.n188 185
R149 VTAIL.n187 VTAIL.n186 185
R150 VTAIL.n116 VTAIL.n115 185
R151 VTAIL.n181 VTAIL.n180 185
R152 VTAIL.n179 VTAIL.n178 185
R153 VTAIL.n120 VTAIL.n119 185
R154 VTAIL.n173 VTAIL.n172 185
R155 VTAIL.n171 VTAIL.n170 185
R156 VTAIL.n124 VTAIL.n123 185
R157 VTAIL.n165 VTAIL.n164 185
R158 VTAIL.n163 VTAIL.n162 185
R159 VTAIL.n161 VTAIL.n127 185
R160 VTAIL.n131 VTAIL.n128 185
R161 VTAIL.n156 VTAIL.n155 185
R162 VTAIL.n154 VTAIL.n153 185
R163 VTAIL.n133 VTAIL.n132 185
R164 VTAIL.n148 VTAIL.n147 185
R165 VTAIL.n146 VTAIL.n145 185
R166 VTAIL.n137 VTAIL.n136 185
R167 VTAIL.n140 VTAIL.n139 185
R168 VTAIL.t0 VTAIL.n339 149.524
R169 VTAIL.t8 VTAIL.n33 149.524
R170 VTAIL.t4 VTAIL.n240 149.524
R171 VTAIL.t11 VTAIL.n138 149.524
R172 VTAIL.n340 VTAIL.n337 104.615
R173 VTAIL.n347 VTAIL.n337 104.615
R174 VTAIL.n348 VTAIL.n347 104.615
R175 VTAIL.n348 VTAIL.n333 104.615
R176 VTAIL.n355 VTAIL.n333 104.615
R177 VTAIL.n357 VTAIL.n355 104.615
R178 VTAIL.n357 VTAIL.n356 104.615
R179 VTAIL.n356 VTAIL.n329 104.615
R180 VTAIL.n365 VTAIL.n329 104.615
R181 VTAIL.n366 VTAIL.n365 104.615
R182 VTAIL.n366 VTAIL.n325 104.615
R183 VTAIL.n373 VTAIL.n325 104.615
R184 VTAIL.n374 VTAIL.n373 104.615
R185 VTAIL.n374 VTAIL.n321 104.615
R186 VTAIL.n381 VTAIL.n321 104.615
R187 VTAIL.n382 VTAIL.n381 104.615
R188 VTAIL.n382 VTAIL.n317 104.615
R189 VTAIL.n389 VTAIL.n317 104.615
R190 VTAIL.n390 VTAIL.n389 104.615
R191 VTAIL.n390 VTAIL.n313 104.615
R192 VTAIL.n397 VTAIL.n313 104.615
R193 VTAIL.n398 VTAIL.n397 104.615
R194 VTAIL.n398 VTAIL.n309 104.615
R195 VTAIL.n405 VTAIL.n309 104.615
R196 VTAIL.n34 VTAIL.n31 104.615
R197 VTAIL.n41 VTAIL.n31 104.615
R198 VTAIL.n42 VTAIL.n41 104.615
R199 VTAIL.n42 VTAIL.n27 104.615
R200 VTAIL.n49 VTAIL.n27 104.615
R201 VTAIL.n51 VTAIL.n49 104.615
R202 VTAIL.n51 VTAIL.n50 104.615
R203 VTAIL.n50 VTAIL.n23 104.615
R204 VTAIL.n59 VTAIL.n23 104.615
R205 VTAIL.n60 VTAIL.n59 104.615
R206 VTAIL.n60 VTAIL.n19 104.615
R207 VTAIL.n67 VTAIL.n19 104.615
R208 VTAIL.n68 VTAIL.n67 104.615
R209 VTAIL.n68 VTAIL.n15 104.615
R210 VTAIL.n75 VTAIL.n15 104.615
R211 VTAIL.n76 VTAIL.n75 104.615
R212 VTAIL.n76 VTAIL.n11 104.615
R213 VTAIL.n83 VTAIL.n11 104.615
R214 VTAIL.n84 VTAIL.n83 104.615
R215 VTAIL.n84 VTAIL.n7 104.615
R216 VTAIL.n91 VTAIL.n7 104.615
R217 VTAIL.n92 VTAIL.n91 104.615
R218 VTAIL.n92 VTAIL.n3 104.615
R219 VTAIL.n99 VTAIL.n3 104.615
R220 VTAIL.n305 VTAIL.n209 104.615
R221 VTAIL.n298 VTAIL.n209 104.615
R222 VTAIL.n298 VTAIL.n297 104.615
R223 VTAIL.n297 VTAIL.n213 104.615
R224 VTAIL.n290 VTAIL.n213 104.615
R225 VTAIL.n290 VTAIL.n289 104.615
R226 VTAIL.n289 VTAIL.n217 104.615
R227 VTAIL.n282 VTAIL.n217 104.615
R228 VTAIL.n282 VTAIL.n281 104.615
R229 VTAIL.n281 VTAIL.n221 104.615
R230 VTAIL.n274 VTAIL.n221 104.615
R231 VTAIL.n274 VTAIL.n273 104.615
R232 VTAIL.n273 VTAIL.n225 104.615
R233 VTAIL.n266 VTAIL.n225 104.615
R234 VTAIL.n266 VTAIL.n265 104.615
R235 VTAIL.n265 VTAIL.n229 104.615
R236 VTAIL.n233 VTAIL.n229 104.615
R237 VTAIL.n257 VTAIL.n233 104.615
R238 VTAIL.n257 VTAIL.n256 104.615
R239 VTAIL.n256 VTAIL.n234 104.615
R240 VTAIL.n249 VTAIL.n234 104.615
R241 VTAIL.n249 VTAIL.n248 104.615
R242 VTAIL.n248 VTAIL.n238 104.615
R243 VTAIL.n241 VTAIL.n238 104.615
R244 VTAIL.n203 VTAIL.n107 104.615
R245 VTAIL.n196 VTAIL.n107 104.615
R246 VTAIL.n196 VTAIL.n195 104.615
R247 VTAIL.n195 VTAIL.n111 104.615
R248 VTAIL.n188 VTAIL.n111 104.615
R249 VTAIL.n188 VTAIL.n187 104.615
R250 VTAIL.n187 VTAIL.n115 104.615
R251 VTAIL.n180 VTAIL.n115 104.615
R252 VTAIL.n180 VTAIL.n179 104.615
R253 VTAIL.n179 VTAIL.n119 104.615
R254 VTAIL.n172 VTAIL.n119 104.615
R255 VTAIL.n172 VTAIL.n171 104.615
R256 VTAIL.n171 VTAIL.n123 104.615
R257 VTAIL.n164 VTAIL.n123 104.615
R258 VTAIL.n164 VTAIL.n163 104.615
R259 VTAIL.n163 VTAIL.n127 104.615
R260 VTAIL.n131 VTAIL.n127 104.615
R261 VTAIL.n155 VTAIL.n131 104.615
R262 VTAIL.n155 VTAIL.n154 104.615
R263 VTAIL.n154 VTAIL.n132 104.615
R264 VTAIL.n147 VTAIL.n132 104.615
R265 VTAIL.n147 VTAIL.n146 104.615
R266 VTAIL.n146 VTAIL.n136 104.615
R267 VTAIL.n139 VTAIL.n136 104.615
R268 VTAIL.n340 VTAIL.t0 52.3082
R269 VTAIL.n34 VTAIL.t8 52.3082
R270 VTAIL.n241 VTAIL.t4 52.3082
R271 VTAIL.n139 VTAIL.t11 52.3082
R272 VTAIL.n207 VTAIL.n206 47.3069
R273 VTAIL.n105 VTAIL.n104 47.3069
R274 VTAIL.n1 VTAIL.n0 47.3068
R275 VTAIL.n103 VTAIL.n102 47.3068
R276 VTAIL.n407 VTAIL.n406 34.9005
R277 VTAIL.n101 VTAIL.n100 34.9005
R278 VTAIL.n307 VTAIL.n306 34.9005
R279 VTAIL.n205 VTAIL.n204 34.9005
R280 VTAIL.n105 VTAIL.n103 32.7462
R281 VTAIL.n407 VTAIL.n307 30.3496
R282 VTAIL.n364 VTAIL.n363 13.1884
R283 VTAIL.n58 VTAIL.n57 13.1884
R284 VTAIL.n264 VTAIL.n263 13.1884
R285 VTAIL.n162 VTAIL.n161 13.1884
R286 VTAIL.n362 VTAIL.n330 12.8005
R287 VTAIL.n367 VTAIL.n328 12.8005
R288 VTAIL.n56 VTAIL.n24 12.8005
R289 VTAIL.n61 VTAIL.n22 12.8005
R290 VTAIL.n267 VTAIL.n228 12.8005
R291 VTAIL.n262 VTAIL.n230 12.8005
R292 VTAIL.n165 VTAIL.n126 12.8005
R293 VTAIL.n160 VTAIL.n128 12.8005
R294 VTAIL.n359 VTAIL.n358 12.0247
R295 VTAIL.n368 VTAIL.n326 12.0247
R296 VTAIL.n404 VTAIL.n308 12.0247
R297 VTAIL.n53 VTAIL.n52 12.0247
R298 VTAIL.n62 VTAIL.n20 12.0247
R299 VTAIL.n98 VTAIL.n2 12.0247
R300 VTAIL.n304 VTAIL.n208 12.0247
R301 VTAIL.n268 VTAIL.n226 12.0247
R302 VTAIL.n259 VTAIL.n258 12.0247
R303 VTAIL.n202 VTAIL.n106 12.0247
R304 VTAIL.n166 VTAIL.n124 12.0247
R305 VTAIL.n157 VTAIL.n156 12.0247
R306 VTAIL.n354 VTAIL.n332 11.249
R307 VTAIL.n372 VTAIL.n371 11.249
R308 VTAIL.n403 VTAIL.n310 11.249
R309 VTAIL.n48 VTAIL.n26 11.249
R310 VTAIL.n66 VTAIL.n65 11.249
R311 VTAIL.n97 VTAIL.n4 11.249
R312 VTAIL.n303 VTAIL.n210 11.249
R313 VTAIL.n272 VTAIL.n271 11.249
R314 VTAIL.n255 VTAIL.n232 11.249
R315 VTAIL.n201 VTAIL.n108 11.249
R316 VTAIL.n170 VTAIL.n169 11.249
R317 VTAIL.n153 VTAIL.n130 11.249
R318 VTAIL.n353 VTAIL.n334 10.4732
R319 VTAIL.n375 VTAIL.n324 10.4732
R320 VTAIL.n400 VTAIL.n399 10.4732
R321 VTAIL.n47 VTAIL.n28 10.4732
R322 VTAIL.n69 VTAIL.n18 10.4732
R323 VTAIL.n94 VTAIL.n93 10.4732
R324 VTAIL.n300 VTAIL.n299 10.4732
R325 VTAIL.n275 VTAIL.n224 10.4732
R326 VTAIL.n254 VTAIL.n235 10.4732
R327 VTAIL.n198 VTAIL.n197 10.4732
R328 VTAIL.n173 VTAIL.n122 10.4732
R329 VTAIL.n152 VTAIL.n133 10.4732
R330 VTAIL.n341 VTAIL.n339 10.2747
R331 VTAIL.n35 VTAIL.n33 10.2747
R332 VTAIL.n242 VTAIL.n240 10.2747
R333 VTAIL.n140 VTAIL.n138 10.2747
R334 VTAIL.n350 VTAIL.n349 9.69747
R335 VTAIL.n376 VTAIL.n322 9.69747
R336 VTAIL.n396 VTAIL.n312 9.69747
R337 VTAIL.n44 VTAIL.n43 9.69747
R338 VTAIL.n70 VTAIL.n16 9.69747
R339 VTAIL.n90 VTAIL.n6 9.69747
R340 VTAIL.n296 VTAIL.n212 9.69747
R341 VTAIL.n276 VTAIL.n222 9.69747
R342 VTAIL.n251 VTAIL.n250 9.69747
R343 VTAIL.n194 VTAIL.n110 9.69747
R344 VTAIL.n174 VTAIL.n120 9.69747
R345 VTAIL.n149 VTAIL.n148 9.69747
R346 VTAIL.n402 VTAIL.n308 9.45567
R347 VTAIL.n96 VTAIL.n2 9.45567
R348 VTAIL.n302 VTAIL.n208 9.45567
R349 VTAIL.n200 VTAIL.n106 9.45567
R350 VTAIL.n387 VTAIL.n386 9.3005
R351 VTAIL.n316 VTAIL.n315 9.3005
R352 VTAIL.n393 VTAIL.n392 9.3005
R353 VTAIL.n395 VTAIL.n394 9.3005
R354 VTAIL.n312 VTAIL.n311 9.3005
R355 VTAIL.n401 VTAIL.n400 9.3005
R356 VTAIL.n403 VTAIL.n402 9.3005
R357 VTAIL.n320 VTAIL.n319 9.3005
R358 VTAIL.n379 VTAIL.n378 9.3005
R359 VTAIL.n377 VTAIL.n376 9.3005
R360 VTAIL.n324 VTAIL.n323 9.3005
R361 VTAIL.n371 VTAIL.n370 9.3005
R362 VTAIL.n369 VTAIL.n368 9.3005
R363 VTAIL.n328 VTAIL.n327 9.3005
R364 VTAIL.n343 VTAIL.n342 9.3005
R365 VTAIL.n345 VTAIL.n344 9.3005
R366 VTAIL.n336 VTAIL.n335 9.3005
R367 VTAIL.n351 VTAIL.n350 9.3005
R368 VTAIL.n353 VTAIL.n352 9.3005
R369 VTAIL.n332 VTAIL.n331 9.3005
R370 VTAIL.n360 VTAIL.n359 9.3005
R371 VTAIL.n362 VTAIL.n361 9.3005
R372 VTAIL.n385 VTAIL.n384 9.3005
R373 VTAIL.n81 VTAIL.n80 9.3005
R374 VTAIL.n10 VTAIL.n9 9.3005
R375 VTAIL.n87 VTAIL.n86 9.3005
R376 VTAIL.n89 VTAIL.n88 9.3005
R377 VTAIL.n6 VTAIL.n5 9.3005
R378 VTAIL.n95 VTAIL.n94 9.3005
R379 VTAIL.n97 VTAIL.n96 9.3005
R380 VTAIL.n14 VTAIL.n13 9.3005
R381 VTAIL.n73 VTAIL.n72 9.3005
R382 VTAIL.n71 VTAIL.n70 9.3005
R383 VTAIL.n18 VTAIL.n17 9.3005
R384 VTAIL.n65 VTAIL.n64 9.3005
R385 VTAIL.n63 VTAIL.n62 9.3005
R386 VTAIL.n22 VTAIL.n21 9.3005
R387 VTAIL.n37 VTAIL.n36 9.3005
R388 VTAIL.n39 VTAIL.n38 9.3005
R389 VTAIL.n30 VTAIL.n29 9.3005
R390 VTAIL.n45 VTAIL.n44 9.3005
R391 VTAIL.n47 VTAIL.n46 9.3005
R392 VTAIL.n26 VTAIL.n25 9.3005
R393 VTAIL.n54 VTAIL.n53 9.3005
R394 VTAIL.n56 VTAIL.n55 9.3005
R395 VTAIL.n79 VTAIL.n78 9.3005
R396 VTAIL.n303 VTAIL.n302 9.3005
R397 VTAIL.n301 VTAIL.n300 9.3005
R398 VTAIL.n212 VTAIL.n211 9.3005
R399 VTAIL.n295 VTAIL.n294 9.3005
R400 VTAIL.n293 VTAIL.n292 9.3005
R401 VTAIL.n216 VTAIL.n215 9.3005
R402 VTAIL.n287 VTAIL.n286 9.3005
R403 VTAIL.n285 VTAIL.n284 9.3005
R404 VTAIL.n220 VTAIL.n219 9.3005
R405 VTAIL.n279 VTAIL.n278 9.3005
R406 VTAIL.n277 VTAIL.n276 9.3005
R407 VTAIL.n224 VTAIL.n223 9.3005
R408 VTAIL.n271 VTAIL.n270 9.3005
R409 VTAIL.n269 VTAIL.n268 9.3005
R410 VTAIL.n228 VTAIL.n227 9.3005
R411 VTAIL.n262 VTAIL.n261 9.3005
R412 VTAIL.n260 VTAIL.n259 9.3005
R413 VTAIL.n232 VTAIL.n231 9.3005
R414 VTAIL.n254 VTAIL.n253 9.3005
R415 VTAIL.n252 VTAIL.n251 9.3005
R416 VTAIL.n237 VTAIL.n236 9.3005
R417 VTAIL.n246 VTAIL.n245 9.3005
R418 VTAIL.n244 VTAIL.n243 9.3005
R419 VTAIL.n142 VTAIL.n141 9.3005
R420 VTAIL.n144 VTAIL.n143 9.3005
R421 VTAIL.n135 VTAIL.n134 9.3005
R422 VTAIL.n150 VTAIL.n149 9.3005
R423 VTAIL.n152 VTAIL.n151 9.3005
R424 VTAIL.n130 VTAIL.n129 9.3005
R425 VTAIL.n158 VTAIL.n157 9.3005
R426 VTAIL.n160 VTAIL.n159 9.3005
R427 VTAIL.n114 VTAIL.n113 9.3005
R428 VTAIL.n191 VTAIL.n190 9.3005
R429 VTAIL.n193 VTAIL.n192 9.3005
R430 VTAIL.n110 VTAIL.n109 9.3005
R431 VTAIL.n199 VTAIL.n198 9.3005
R432 VTAIL.n201 VTAIL.n200 9.3005
R433 VTAIL.n185 VTAIL.n184 9.3005
R434 VTAIL.n183 VTAIL.n182 9.3005
R435 VTAIL.n118 VTAIL.n117 9.3005
R436 VTAIL.n177 VTAIL.n176 9.3005
R437 VTAIL.n175 VTAIL.n174 9.3005
R438 VTAIL.n122 VTAIL.n121 9.3005
R439 VTAIL.n169 VTAIL.n168 9.3005
R440 VTAIL.n167 VTAIL.n166 9.3005
R441 VTAIL.n126 VTAIL.n125 9.3005
R442 VTAIL.n346 VTAIL.n336 8.92171
R443 VTAIL.n380 VTAIL.n379 8.92171
R444 VTAIL.n395 VTAIL.n314 8.92171
R445 VTAIL.n40 VTAIL.n30 8.92171
R446 VTAIL.n74 VTAIL.n73 8.92171
R447 VTAIL.n89 VTAIL.n8 8.92171
R448 VTAIL.n295 VTAIL.n214 8.92171
R449 VTAIL.n280 VTAIL.n279 8.92171
R450 VTAIL.n247 VTAIL.n237 8.92171
R451 VTAIL.n193 VTAIL.n112 8.92171
R452 VTAIL.n178 VTAIL.n177 8.92171
R453 VTAIL.n145 VTAIL.n135 8.92171
R454 VTAIL.n345 VTAIL.n338 8.14595
R455 VTAIL.n383 VTAIL.n320 8.14595
R456 VTAIL.n392 VTAIL.n391 8.14595
R457 VTAIL.n39 VTAIL.n32 8.14595
R458 VTAIL.n77 VTAIL.n14 8.14595
R459 VTAIL.n86 VTAIL.n85 8.14595
R460 VTAIL.n292 VTAIL.n291 8.14595
R461 VTAIL.n283 VTAIL.n220 8.14595
R462 VTAIL.n246 VTAIL.n239 8.14595
R463 VTAIL.n190 VTAIL.n189 8.14595
R464 VTAIL.n181 VTAIL.n118 8.14595
R465 VTAIL.n144 VTAIL.n137 8.14595
R466 VTAIL.n342 VTAIL.n341 7.3702
R467 VTAIL.n384 VTAIL.n318 7.3702
R468 VTAIL.n388 VTAIL.n316 7.3702
R469 VTAIL.n36 VTAIL.n35 7.3702
R470 VTAIL.n78 VTAIL.n12 7.3702
R471 VTAIL.n82 VTAIL.n10 7.3702
R472 VTAIL.n288 VTAIL.n216 7.3702
R473 VTAIL.n284 VTAIL.n218 7.3702
R474 VTAIL.n243 VTAIL.n242 7.3702
R475 VTAIL.n186 VTAIL.n114 7.3702
R476 VTAIL.n182 VTAIL.n116 7.3702
R477 VTAIL.n141 VTAIL.n140 7.3702
R478 VTAIL.n387 VTAIL.n318 6.59444
R479 VTAIL.n388 VTAIL.n387 6.59444
R480 VTAIL.n81 VTAIL.n12 6.59444
R481 VTAIL.n82 VTAIL.n81 6.59444
R482 VTAIL.n288 VTAIL.n287 6.59444
R483 VTAIL.n287 VTAIL.n218 6.59444
R484 VTAIL.n186 VTAIL.n185 6.59444
R485 VTAIL.n185 VTAIL.n116 6.59444
R486 VTAIL.n342 VTAIL.n338 5.81868
R487 VTAIL.n384 VTAIL.n383 5.81868
R488 VTAIL.n391 VTAIL.n316 5.81868
R489 VTAIL.n36 VTAIL.n32 5.81868
R490 VTAIL.n78 VTAIL.n77 5.81868
R491 VTAIL.n85 VTAIL.n10 5.81868
R492 VTAIL.n291 VTAIL.n216 5.81868
R493 VTAIL.n284 VTAIL.n283 5.81868
R494 VTAIL.n243 VTAIL.n239 5.81868
R495 VTAIL.n189 VTAIL.n114 5.81868
R496 VTAIL.n182 VTAIL.n181 5.81868
R497 VTAIL.n141 VTAIL.n137 5.81868
R498 VTAIL.n346 VTAIL.n345 5.04292
R499 VTAIL.n380 VTAIL.n320 5.04292
R500 VTAIL.n392 VTAIL.n314 5.04292
R501 VTAIL.n40 VTAIL.n39 5.04292
R502 VTAIL.n74 VTAIL.n14 5.04292
R503 VTAIL.n86 VTAIL.n8 5.04292
R504 VTAIL.n292 VTAIL.n214 5.04292
R505 VTAIL.n280 VTAIL.n220 5.04292
R506 VTAIL.n247 VTAIL.n246 5.04292
R507 VTAIL.n190 VTAIL.n112 5.04292
R508 VTAIL.n178 VTAIL.n118 5.04292
R509 VTAIL.n145 VTAIL.n144 5.04292
R510 VTAIL.n349 VTAIL.n336 4.26717
R511 VTAIL.n379 VTAIL.n322 4.26717
R512 VTAIL.n396 VTAIL.n395 4.26717
R513 VTAIL.n43 VTAIL.n30 4.26717
R514 VTAIL.n73 VTAIL.n16 4.26717
R515 VTAIL.n90 VTAIL.n89 4.26717
R516 VTAIL.n296 VTAIL.n295 4.26717
R517 VTAIL.n279 VTAIL.n222 4.26717
R518 VTAIL.n250 VTAIL.n237 4.26717
R519 VTAIL.n194 VTAIL.n193 4.26717
R520 VTAIL.n177 VTAIL.n120 4.26717
R521 VTAIL.n148 VTAIL.n135 4.26717
R522 VTAIL.n350 VTAIL.n334 3.49141
R523 VTAIL.n376 VTAIL.n375 3.49141
R524 VTAIL.n399 VTAIL.n312 3.49141
R525 VTAIL.n44 VTAIL.n28 3.49141
R526 VTAIL.n70 VTAIL.n69 3.49141
R527 VTAIL.n93 VTAIL.n6 3.49141
R528 VTAIL.n299 VTAIL.n212 3.49141
R529 VTAIL.n276 VTAIL.n275 3.49141
R530 VTAIL.n251 VTAIL.n235 3.49141
R531 VTAIL.n197 VTAIL.n110 3.49141
R532 VTAIL.n174 VTAIL.n173 3.49141
R533 VTAIL.n149 VTAIL.n133 3.49141
R534 VTAIL.n142 VTAIL.n138 2.84303
R535 VTAIL.n343 VTAIL.n339 2.84303
R536 VTAIL.n37 VTAIL.n33 2.84303
R537 VTAIL.n244 VTAIL.n240 2.84303
R538 VTAIL.n354 VTAIL.n353 2.71565
R539 VTAIL.n372 VTAIL.n324 2.71565
R540 VTAIL.n400 VTAIL.n310 2.71565
R541 VTAIL.n48 VTAIL.n47 2.71565
R542 VTAIL.n66 VTAIL.n18 2.71565
R543 VTAIL.n94 VTAIL.n4 2.71565
R544 VTAIL.n300 VTAIL.n210 2.71565
R545 VTAIL.n272 VTAIL.n224 2.71565
R546 VTAIL.n255 VTAIL.n254 2.71565
R547 VTAIL.n198 VTAIL.n108 2.71565
R548 VTAIL.n170 VTAIL.n122 2.71565
R549 VTAIL.n153 VTAIL.n152 2.71565
R550 VTAIL.n205 VTAIL.n105 2.39705
R551 VTAIL.n307 VTAIL.n207 2.39705
R552 VTAIL.n103 VTAIL.n101 2.39705
R553 VTAIL.n358 VTAIL.n332 1.93989
R554 VTAIL.n371 VTAIL.n326 1.93989
R555 VTAIL.n404 VTAIL.n403 1.93989
R556 VTAIL.n52 VTAIL.n26 1.93989
R557 VTAIL.n65 VTAIL.n20 1.93989
R558 VTAIL.n98 VTAIL.n97 1.93989
R559 VTAIL.n304 VTAIL.n303 1.93989
R560 VTAIL.n271 VTAIL.n226 1.93989
R561 VTAIL.n258 VTAIL.n232 1.93989
R562 VTAIL.n202 VTAIL.n201 1.93989
R563 VTAIL.n169 VTAIL.n124 1.93989
R564 VTAIL.n156 VTAIL.n130 1.93989
R565 VTAIL VTAIL.n407 1.73972
R566 VTAIL.n207 VTAIL.n205 1.6686
R567 VTAIL.n101 VTAIL.n1 1.6686
R568 VTAIL.n359 VTAIL.n330 1.16414
R569 VTAIL.n368 VTAIL.n367 1.16414
R570 VTAIL.n406 VTAIL.n308 1.16414
R571 VTAIL.n53 VTAIL.n24 1.16414
R572 VTAIL.n62 VTAIL.n61 1.16414
R573 VTAIL.n100 VTAIL.n2 1.16414
R574 VTAIL.n306 VTAIL.n208 1.16414
R575 VTAIL.n268 VTAIL.n267 1.16414
R576 VTAIL.n259 VTAIL.n230 1.16414
R577 VTAIL.n204 VTAIL.n106 1.16414
R578 VTAIL.n166 VTAIL.n165 1.16414
R579 VTAIL.n157 VTAIL.n128 1.16414
R580 VTAIL.n0 VTAIL.t3 1.09563
R581 VTAIL.n0 VTAIL.t10 1.09563
R582 VTAIL.n102 VTAIL.t7 1.09563
R583 VTAIL.n102 VTAIL.t9 1.09563
R584 VTAIL.n206 VTAIL.t5 1.09563
R585 VTAIL.n206 VTAIL.t6 1.09563
R586 VTAIL.n104 VTAIL.t1 1.09563
R587 VTAIL.n104 VTAIL.t2 1.09563
R588 VTAIL VTAIL.n1 0.657828
R589 VTAIL.n363 VTAIL.n362 0.388379
R590 VTAIL.n364 VTAIL.n328 0.388379
R591 VTAIL.n57 VTAIL.n56 0.388379
R592 VTAIL.n58 VTAIL.n22 0.388379
R593 VTAIL.n264 VTAIL.n228 0.388379
R594 VTAIL.n263 VTAIL.n262 0.388379
R595 VTAIL.n162 VTAIL.n126 0.388379
R596 VTAIL.n161 VTAIL.n160 0.388379
R597 VTAIL.n344 VTAIL.n343 0.155672
R598 VTAIL.n344 VTAIL.n335 0.155672
R599 VTAIL.n351 VTAIL.n335 0.155672
R600 VTAIL.n352 VTAIL.n351 0.155672
R601 VTAIL.n352 VTAIL.n331 0.155672
R602 VTAIL.n360 VTAIL.n331 0.155672
R603 VTAIL.n361 VTAIL.n360 0.155672
R604 VTAIL.n361 VTAIL.n327 0.155672
R605 VTAIL.n369 VTAIL.n327 0.155672
R606 VTAIL.n370 VTAIL.n369 0.155672
R607 VTAIL.n370 VTAIL.n323 0.155672
R608 VTAIL.n377 VTAIL.n323 0.155672
R609 VTAIL.n378 VTAIL.n377 0.155672
R610 VTAIL.n378 VTAIL.n319 0.155672
R611 VTAIL.n385 VTAIL.n319 0.155672
R612 VTAIL.n386 VTAIL.n385 0.155672
R613 VTAIL.n386 VTAIL.n315 0.155672
R614 VTAIL.n393 VTAIL.n315 0.155672
R615 VTAIL.n394 VTAIL.n393 0.155672
R616 VTAIL.n394 VTAIL.n311 0.155672
R617 VTAIL.n401 VTAIL.n311 0.155672
R618 VTAIL.n402 VTAIL.n401 0.155672
R619 VTAIL.n38 VTAIL.n37 0.155672
R620 VTAIL.n38 VTAIL.n29 0.155672
R621 VTAIL.n45 VTAIL.n29 0.155672
R622 VTAIL.n46 VTAIL.n45 0.155672
R623 VTAIL.n46 VTAIL.n25 0.155672
R624 VTAIL.n54 VTAIL.n25 0.155672
R625 VTAIL.n55 VTAIL.n54 0.155672
R626 VTAIL.n55 VTAIL.n21 0.155672
R627 VTAIL.n63 VTAIL.n21 0.155672
R628 VTAIL.n64 VTAIL.n63 0.155672
R629 VTAIL.n64 VTAIL.n17 0.155672
R630 VTAIL.n71 VTAIL.n17 0.155672
R631 VTAIL.n72 VTAIL.n71 0.155672
R632 VTAIL.n72 VTAIL.n13 0.155672
R633 VTAIL.n79 VTAIL.n13 0.155672
R634 VTAIL.n80 VTAIL.n79 0.155672
R635 VTAIL.n80 VTAIL.n9 0.155672
R636 VTAIL.n87 VTAIL.n9 0.155672
R637 VTAIL.n88 VTAIL.n87 0.155672
R638 VTAIL.n88 VTAIL.n5 0.155672
R639 VTAIL.n95 VTAIL.n5 0.155672
R640 VTAIL.n96 VTAIL.n95 0.155672
R641 VTAIL.n302 VTAIL.n301 0.155672
R642 VTAIL.n301 VTAIL.n211 0.155672
R643 VTAIL.n294 VTAIL.n211 0.155672
R644 VTAIL.n294 VTAIL.n293 0.155672
R645 VTAIL.n293 VTAIL.n215 0.155672
R646 VTAIL.n286 VTAIL.n215 0.155672
R647 VTAIL.n286 VTAIL.n285 0.155672
R648 VTAIL.n285 VTAIL.n219 0.155672
R649 VTAIL.n278 VTAIL.n219 0.155672
R650 VTAIL.n278 VTAIL.n277 0.155672
R651 VTAIL.n277 VTAIL.n223 0.155672
R652 VTAIL.n270 VTAIL.n223 0.155672
R653 VTAIL.n270 VTAIL.n269 0.155672
R654 VTAIL.n269 VTAIL.n227 0.155672
R655 VTAIL.n261 VTAIL.n227 0.155672
R656 VTAIL.n261 VTAIL.n260 0.155672
R657 VTAIL.n260 VTAIL.n231 0.155672
R658 VTAIL.n253 VTAIL.n231 0.155672
R659 VTAIL.n253 VTAIL.n252 0.155672
R660 VTAIL.n252 VTAIL.n236 0.155672
R661 VTAIL.n245 VTAIL.n236 0.155672
R662 VTAIL.n245 VTAIL.n244 0.155672
R663 VTAIL.n200 VTAIL.n199 0.155672
R664 VTAIL.n199 VTAIL.n109 0.155672
R665 VTAIL.n192 VTAIL.n109 0.155672
R666 VTAIL.n192 VTAIL.n191 0.155672
R667 VTAIL.n191 VTAIL.n113 0.155672
R668 VTAIL.n184 VTAIL.n113 0.155672
R669 VTAIL.n184 VTAIL.n183 0.155672
R670 VTAIL.n183 VTAIL.n117 0.155672
R671 VTAIL.n176 VTAIL.n117 0.155672
R672 VTAIL.n176 VTAIL.n175 0.155672
R673 VTAIL.n175 VTAIL.n121 0.155672
R674 VTAIL.n168 VTAIL.n121 0.155672
R675 VTAIL.n168 VTAIL.n167 0.155672
R676 VTAIL.n167 VTAIL.n125 0.155672
R677 VTAIL.n159 VTAIL.n125 0.155672
R678 VTAIL.n159 VTAIL.n158 0.155672
R679 VTAIL.n158 VTAIL.n129 0.155672
R680 VTAIL.n151 VTAIL.n129 0.155672
R681 VTAIL.n151 VTAIL.n150 0.155672
R682 VTAIL.n150 VTAIL.n134 0.155672
R683 VTAIL.n143 VTAIL.n134 0.155672
R684 VTAIL.n143 VTAIL.n142 0.155672
R685 VDD1.n98 VDD1.n97 289.615
R686 VDD1.n197 VDD1.n196 289.615
R687 VDD1.n97 VDD1.n96 185
R688 VDD1.n2 VDD1.n1 185
R689 VDD1.n91 VDD1.n90 185
R690 VDD1.n89 VDD1.n88 185
R691 VDD1.n6 VDD1.n5 185
R692 VDD1.n83 VDD1.n82 185
R693 VDD1.n81 VDD1.n80 185
R694 VDD1.n10 VDD1.n9 185
R695 VDD1.n75 VDD1.n74 185
R696 VDD1.n73 VDD1.n72 185
R697 VDD1.n14 VDD1.n13 185
R698 VDD1.n67 VDD1.n66 185
R699 VDD1.n65 VDD1.n64 185
R700 VDD1.n18 VDD1.n17 185
R701 VDD1.n59 VDD1.n58 185
R702 VDD1.n57 VDD1.n56 185
R703 VDD1.n55 VDD1.n21 185
R704 VDD1.n25 VDD1.n22 185
R705 VDD1.n50 VDD1.n49 185
R706 VDD1.n48 VDD1.n47 185
R707 VDD1.n27 VDD1.n26 185
R708 VDD1.n42 VDD1.n41 185
R709 VDD1.n40 VDD1.n39 185
R710 VDD1.n31 VDD1.n30 185
R711 VDD1.n34 VDD1.n33 185
R712 VDD1.n132 VDD1.n131 185
R713 VDD1.n129 VDD1.n128 185
R714 VDD1.n138 VDD1.n137 185
R715 VDD1.n140 VDD1.n139 185
R716 VDD1.n125 VDD1.n124 185
R717 VDD1.n146 VDD1.n145 185
R718 VDD1.n149 VDD1.n148 185
R719 VDD1.n147 VDD1.n121 185
R720 VDD1.n154 VDD1.n120 185
R721 VDD1.n156 VDD1.n155 185
R722 VDD1.n158 VDD1.n157 185
R723 VDD1.n117 VDD1.n116 185
R724 VDD1.n164 VDD1.n163 185
R725 VDD1.n166 VDD1.n165 185
R726 VDD1.n113 VDD1.n112 185
R727 VDD1.n172 VDD1.n171 185
R728 VDD1.n174 VDD1.n173 185
R729 VDD1.n109 VDD1.n108 185
R730 VDD1.n180 VDD1.n179 185
R731 VDD1.n182 VDD1.n181 185
R732 VDD1.n105 VDD1.n104 185
R733 VDD1.n188 VDD1.n187 185
R734 VDD1.n190 VDD1.n189 185
R735 VDD1.n101 VDD1.n100 185
R736 VDD1.n196 VDD1.n195 185
R737 VDD1.t2 VDD1.n32 149.524
R738 VDD1.t4 VDD1.n130 149.524
R739 VDD1.n97 VDD1.n1 104.615
R740 VDD1.n90 VDD1.n1 104.615
R741 VDD1.n90 VDD1.n89 104.615
R742 VDD1.n89 VDD1.n5 104.615
R743 VDD1.n82 VDD1.n5 104.615
R744 VDD1.n82 VDD1.n81 104.615
R745 VDD1.n81 VDD1.n9 104.615
R746 VDD1.n74 VDD1.n9 104.615
R747 VDD1.n74 VDD1.n73 104.615
R748 VDD1.n73 VDD1.n13 104.615
R749 VDD1.n66 VDD1.n13 104.615
R750 VDD1.n66 VDD1.n65 104.615
R751 VDD1.n65 VDD1.n17 104.615
R752 VDD1.n58 VDD1.n17 104.615
R753 VDD1.n58 VDD1.n57 104.615
R754 VDD1.n57 VDD1.n21 104.615
R755 VDD1.n25 VDD1.n21 104.615
R756 VDD1.n49 VDD1.n25 104.615
R757 VDD1.n49 VDD1.n48 104.615
R758 VDD1.n48 VDD1.n26 104.615
R759 VDD1.n41 VDD1.n26 104.615
R760 VDD1.n41 VDD1.n40 104.615
R761 VDD1.n40 VDD1.n30 104.615
R762 VDD1.n33 VDD1.n30 104.615
R763 VDD1.n131 VDD1.n128 104.615
R764 VDD1.n138 VDD1.n128 104.615
R765 VDD1.n139 VDD1.n138 104.615
R766 VDD1.n139 VDD1.n124 104.615
R767 VDD1.n146 VDD1.n124 104.615
R768 VDD1.n148 VDD1.n146 104.615
R769 VDD1.n148 VDD1.n147 104.615
R770 VDD1.n147 VDD1.n120 104.615
R771 VDD1.n156 VDD1.n120 104.615
R772 VDD1.n157 VDD1.n156 104.615
R773 VDD1.n157 VDD1.n116 104.615
R774 VDD1.n164 VDD1.n116 104.615
R775 VDD1.n165 VDD1.n164 104.615
R776 VDD1.n165 VDD1.n112 104.615
R777 VDD1.n172 VDD1.n112 104.615
R778 VDD1.n173 VDD1.n172 104.615
R779 VDD1.n173 VDD1.n108 104.615
R780 VDD1.n180 VDD1.n108 104.615
R781 VDD1.n181 VDD1.n180 104.615
R782 VDD1.n181 VDD1.n104 104.615
R783 VDD1.n188 VDD1.n104 104.615
R784 VDD1.n189 VDD1.n188 104.615
R785 VDD1.n189 VDD1.n100 104.615
R786 VDD1.n196 VDD1.n100 104.615
R787 VDD1.n199 VDD1.n198 64.5293
R788 VDD1.n201 VDD1.n200 63.9845
R789 VDD1 VDD1.n98 53.4349
R790 VDD1.n199 VDD1.n197 53.3214
R791 VDD1.n33 VDD1.t2 52.3082
R792 VDD1.n131 VDD1.t4 52.3082
R793 VDD1.n201 VDD1.n199 48.8716
R794 VDD1.n56 VDD1.n55 13.1884
R795 VDD1.n155 VDD1.n154 13.1884
R796 VDD1.n59 VDD1.n20 12.8005
R797 VDD1.n54 VDD1.n22 12.8005
R798 VDD1.n153 VDD1.n121 12.8005
R799 VDD1.n158 VDD1.n119 12.8005
R800 VDD1.n96 VDD1.n0 12.0247
R801 VDD1.n60 VDD1.n18 12.0247
R802 VDD1.n51 VDD1.n50 12.0247
R803 VDD1.n150 VDD1.n149 12.0247
R804 VDD1.n159 VDD1.n117 12.0247
R805 VDD1.n195 VDD1.n99 12.0247
R806 VDD1.n95 VDD1.n2 11.249
R807 VDD1.n64 VDD1.n63 11.249
R808 VDD1.n47 VDD1.n24 11.249
R809 VDD1.n145 VDD1.n123 11.249
R810 VDD1.n163 VDD1.n162 11.249
R811 VDD1.n194 VDD1.n101 11.249
R812 VDD1.n92 VDD1.n91 10.4732
R813 VDD1.n67 VDD1.n16 10.4732
R814 VDD1.n46 VDD1.n27 10.4732
R815 VDD1.n144 VDD1.n125 10.4732
R816 VDD1.n166 VDD1.n115 10.4732
R817 VDD1.n191 VDD1.n190 10.4732
R818 VDD1.n34 VDD1.n32 10.2747
R819 VDD1.n132 VDD1.n130 10.2747
R820 VDD1.n88 VDD1.n4 9.69747
R821 VDD1.n68 VDD1.n14 9.69747
R822 VDD1.n43 VDD1.n42 9.69747
R823 VDD1.n141 VDD1.n140 9.69747
R824 VDD1.n167 VDD1.n113 9.69747
R825 VDD1.n187 VDD1.n103 9.69747
R826 VDD1.n94 VDD1.n0 9.45567
R827 VDD1.n193 VDD1.n99 9.45567
R828 VDD1.n36 VDD1.n35 9.3005
R829 VDD1.n38 VDD1.n37 9.3005
R830 VDD1.n29 VDD1.n28 9.3005
R831 VDD1.n44 VDD1.n43 9.3005
R832 VDD1.n46 VDD1.n45 9.3005
R833 VDD1.n24 VDD1.n23 9.3005
R834 VDD1.n52 VDD1.n51 9.3005
R835 VDD1.n54 VDD1.n53 9.3005
R836 VDD1.n8 VDD1.n7 9.3005
R837 VDD1.n85 VDD1.n84 9.3005
R838 VDD1.n87 VDD1.n86 9.3005
R839 VDD1.n4 VDD1.n3 9.3005
R840 VDD1.n93 VDD1.n92 9.3005
R841 VDD1.n95 VDD1.n94 9.3005
R842 VDD1.n79 VDD1.n78 9.3005
R843 VDD1.n77 VDD1.n76 9.3005
R844 VDD1.n12 VDD1.n11 9.3005
R845 VDD1.n71 VDD1.n70 9.3005
R846 VDD1.n69 VDD1.n68 9.3005
R847 VDD1.n16 VDD1.n15 9.3005
R848 VDD1.n63 VDD1.n62 9.3005
R849 VDD1.n61 VDD1.n60 9.3005
R850 VDD1.n20 VDD1.n19 9.3005
R851 VDD1.n178 VDD1.n177 9.3005
R852 VDD1.n107 VDD1.n106 9.3005
R853 VDD1.n184 VDD1.n183 9.3005
R854 VDD1.n186 VDD1.n185 9.3005
R855 VDD1.n103 VDD1.n102 9.3005
R856 VDD1.n192 VDD1.n191 9.3005
R857 VDD1.n194 VDD1.n193 9.3005
R858 VDD1.n111 VDD1.n110 9.3005
R859 VDD1.n170 VDD1.n169 9.3005
R860 VDD1.n168 VDD1.n167 9.3005
R861 VDD1.n115 VDD1.n114 9.3005
R862 VDD1.n162 VDD1.n161 9.3005
R863 VDD1.n160 VDD1.n159 9.3005
R864 VDD1.n119 VDD1.n118 9.3005
R865 VDD1.n134 VDD1.n133 9.3005
R866 VDD1.n136 VDD1.n135 9.3005
R867 VDD1.n127 VDD1.n126 9.3005
R868 VDD1.n142 VDD1.n141 9.3005
R869 VDD1.n144 VDD1.n143 9.3005
R870 VDD1.n123 VDD1.n122 9.3005
R871 VDD1.n151 VDD1.n150 9.3005
R872 VDD1.n153 VDD1.n152 9.3005
R873 VDD1.n176 VDD1.n175 9.3005
R874 VDD1.n87 VDD1.n6 8.92171
R875 VDD1.n72 VDD1.n71 8.92171
R876 VDD1.n39 VDD1.n29 8.92171
R877 VDD1.n137 VDD1.n127 8.92171
R878 VDD1.n171 VDD1.n170 8.92171
R879 VDD1.n186 VDD1.n105 8.92171
R880 VDD1.n84 VDD1.n83 8.14595
R881 VDD1.n75 VDD1.n12 8.14595
R882 VDD1.n38 VDD1.n31 8.14595
R883 VDD1.n136 VDD1.n129 8.14595
R884 VDD1.n174 VDD1.n111 8.14595
R885 VDD1.n183 VDD1.n182 8.14595
R886 VDD1.n80 VDD1.n8 7.3702
R887 VDD1.n76 VDD1.n10 7.3702
R888 VDD1.n35 VDD1.n34 7.3702
R889 VDD1.n133 VDD1.n132 7.3702
R890 VDD1.n175 VDD1.n109 7.3702
R891 VDD1.n179 VDD1.n107 7.3702
R892 VDD1.n80 VDD1.n79 6.59444
R893 VDD1.n79 VDD1.n10 6.59444
R894 VDD1.n178 VDD1.n109 6.59444
R895 VDD1.n179 VDD1.n178 6.59444
R896 VDD1.n83 VDD1.n8 5.81868
R897 VDD1.n76 VDD1.n75 5.81868
R898 VDD1.n35 VDD1.n31 5.81868
R899 VDD1.n133 VDD1.n129 5.81868
R900 VDD1.n175 VDD1.n174 5.81868
R901 VDD1.n182 VDD1.n107 5.81868
R902 VDD1.n84 VDD1.n6 5.04292
R903 VDD1.n72 VDD1.n12 5.04292
R904 VDD1.n39 VDD1.n38 5.04292
R905 VDD1.n137 VDD1.n136 5.04292
R906 VDD1.n171 VDD1.n111 5.04292
R907 VDD1.n183 VDD1.n105 5.04292
R908 VDD1.n88 VDD1.n87 4.26717
R909 VDD1.n71 VDD1.n14 4.26717
R910 VDD1.n42 VDD1.n29 4.26717
R911 VDD1.n140 VDD1.n127 4.26717
R912 VDD1.n170 VDD1.n113 4.26717
R913 VDD1.n187 VDD1.n186 4.26717
R914 VDD1.n91 VDD1.n4 3.49141
R915 VDD1.n68 VDD1.n67 3.49141
R916 VDD1.n43 VDD1.n27 3.49141
R917 VDD1.n141 VDD1.n125 3.49141
R918 VDD1.n167 VDD1.n166 3.49141
R919 VDD1.n190 VDD1.n103 3.49141
R920 VDD1.n36 VDD1.n32 2.84303
R921 VDD1.n134 VDD1.n130 2.84303
R922 VDD1.n92 VDD1.n2 2.71565
R923 VDD1.n64 VDD1.n16 2.71565
R924 VDD1.n47 VDD1.n46 2.71565
R925 VDD1.n145 VDD1.n144 2.71565
R926 VDD1.n163 VDD1.n115 2.71565
R927 VDD1.n191 VDD1.n101 2.71565
R928 VDD1.n96 VDD1.n95 1.93989
R929 VDD1.n63 VDD1.n18 1.93989
R930 VDD1.n50 VDD1.n24 1.93989
R931 VDD1.n149 VDD1.n123 1.93989
R932 VDD1.n162 VDD1.n117 1.93989
R933 VDD1.n195 VDD1.n194 1.93989
R934 VDD1.n98 VDD1.n0 1.16414
R935 VDD1.n60 VDD1.n59 1.16414
R936 VDD1.n51 VDD1.n22 1.16414
R937 VDD1.n150 VDD1.n121 1.16414
R938 VDD1.n159 VDD1.n158 1.16414
R939 VDD1.n197 VDD1.n99 1.16414
R940 VDD1.n200 VDD1.t1 1.09563
R941 VDD1.n200 VDD1.t5 1.09563
R942 VDD1.n198 VDD1.t0 1.09563
R943 VDD1.n198 VDD1.t3 1.09563
R944 VDD1 VDD1.n201 0.541448
R945 VDD1.n56 VDD1.n20 0.388379
R946 VDD1.n55 VDD1.n54 0.388379
R947 VDD1.n154 VDD1.n153 0.388379
R948 VDD1.n155 VDD1.n119 0.388379
R949 VDD1.n94 VDD1.n93 0.155672
R950 VDD1.n93 VDD1.n3 0.155672
R951 VDD1.n86 VDD1.n3 0.155672
R952 VDD1.n86 VDD1.n85 0.155672
R953 VDD1.n85 VDD1.n7 0.155672
R954 VDD1.n78 VDD1.n7 0.155672
R955 VDD1.n78 VDD1.n77 0.155672
R956 VDD1.n77 VDD1.n11 0.155672
R957 VDD1.n70 VDD1.n11 0.155672
R958 VDD1.n70 VDD1.n69 0.155672
R959 VDD1.n69 VDD1.n15 0.155672
R960 VDD1.n62 VDD1.n15 0.155672
R961 VDD1.n62 VDD1.n61 0.155672
R962 VDD1.n61 VDD1.n19 0.155672
R963 VDD1.n53 VDD1.n19 0.155672
R964 VDD1.n53 VDD1.n52 0.155672
R965 VDD1.n52 VDD1.n23 0.155672
R966 VDD1.n45 VDD1.n23 0.155672
R967 VDD1.n45 VDD1.n44 0.155672
R968 VDD1.n44 VDD1.n28 0.155672
R969 VDD1.n37 VDD1.n28 0.155672
R970 VDD1.n37 VDD1.n36 0.155672
R971 VDD1.n135 VDD1.n134 0.155672
R972 VDD1.n135 VDD1.n126 0.155672
R973 VDD1.n142 VDD1.n126 0.155672
R974 VDD1.n143 VDD1.n142 0.155672
R975 VDD1.n143 VDD1.n122 0.155672
R976 VDD1.n151 VDD1.n122 0.155672
R977 VDD1.n152 VDD1.n151 0.155672
R978 VDD1.n152 VDD1.n118 0.155672
R979 VDD1.n160 VDD1.n118 0.155672
R980 VDD1.n161 VDD1.n160 0.155672
R981 VDD1.n161 VDD1.n114 0.155672
R982 VDD1.n168 VDD1.n114 0.155672
R983 VDD1.n169 VDD1.n168 0.155672
R984 VDD1.n169 VDD1.n110 0.155672
R985 VDD1.n176 VDD1.n110 0.155672
R986 VDD1.n177 VDD1.n176 0.155672
R987 VDD1.n177 VDD1.n106 0.155672
R988 VDD1.n184 VDD1.n106 0.155672
R989 VDD1.n185 VDD1.n184 0.155672
R990 VDD1.n185 VDD1.n102 0.155672
R991 VDD1.n192 VDD1.n102 0.155672
R992 VDD1.n193 VDD1.n192 0.155672
R993 B.n987 B.n986 585
R994 B.n988 B.n987 585
R995 B.n402 B.n141 585
R996 B.n401 B.n400 585
R997 B.n399 B.n398 585
R998 B.n397 B.n396 585
R999 B.n395 B.n394 585
R1000 B.n393 B.n392 585
R1001 B.n391 B.n390 585
R1002 B.n389 B.n388 585
R1003 B.n387 B.n386 585
R1004 B.n385 B.n384 585
R1005 B.n383 B.n382 585
R1006 B.n381 B.n380 585
R1007 B.n379 B.n378 585
R1008 B.n377 B.n376 585
R1009 B.n375 B.n374 585
R1010 B.n373 B.n372 585
R1011 B.n371 B.n370 585
R1012 B.n369 B.n368 585
R1013 B.n367 B.n366 585
R1014 B.n365 B.n364 585
R1015 B.n363 B.n362 585
R1016 B.n361 B.n360 585
R1017 B.n359 B.n358 585
R1018 B.n357 B.n356 585
R1019 B.n355 B.n354 585
R1020 B.n353 B.n352 585
R1021 B.n351 B.n350 585
R1022 B.n349 B.n348 585
R1023 B.n347 B.n346 585
R1024 B.n345 B.n344 585
R1025 B.n343 B.n342 585
R1026 B.n341 B.n340 585
R1027 B.n339 B.n338 585
R1028 B.n337 B.n336 585
R1029 B.n335 B.n334 585
R1030 B.n333 B.n332 585
R1031 B.n331 B.n330 585
R1032 B.n329 B.n328 585
R1033 B.n327 B.n326 585
R1034 B.n325 B.n324 585
R1035 B.n323 B.n322 585
R1036 B.n321 B.n320 585
R1037 B.n319 B.n318 585
R1038 B.n317 B.n316 585
R1039 B.n315 B.n314 585
R1040 B.n313 B.n312 585
R1041 B.n311 B.n310 585
R1042 B.n309 B.n308 585
R1043 B.n307 B.n306 585
R1044 B.n305 B.n304 585
R1045 B.n303 B.n302 585
R1046 B.n301 B.n300 585
R1047 B.n299 B.n298 585
R1048 B.n297 B.n296 585
R1049 B.n295 B.n294 585
R1050 B.n293 B.n292 585
R1051 B.n291 B.n290 585
R1052 B.n289 B.n288 585
R1053 B.n287 B.n286 585
R1054 B.n284 B.n283 585
R1055 B.n282 B.n281 585
R1056 B.n280 B.n279 585
R1057 B.n278 B.n277 585
R1058 B.n276 B.n275 585
R1059 B.n274 B.n273 585
R1060 B.n272 B.n271 585
R1061 B.n270 B.n269 585
R1062 B.n268 B.n267 585
R1063 B.n266 B.n265 585
R1064 B.n264 B.n263 585
R1065 B.n262 B.n261 585
R1066 B.n260 B.n259 585
R1067 B.n258 B.n257 585
R1068 B.n256 B.n255 585
R1069 B.n254 B.n253 585
R1070 B.n252 B.n251 585
R1071 B.n250 B.n249 585
R1072 B.n248 B.n247 585
R1073 B.n246 B.n245 585
R1074 B.n244 B.n243 585
R1075 B.n242 B.n241 585
R1076 B.n240 B.n239 585
R1077 B.n238 B.n237 585
R1078 B.n236 B.n235 585
R1079 B.n234 B.n233 585
R1080 B.n232 B.n231 585
R1081 B.n230 B.n229 585
R1082 B.n228 B.n227 585
R1083 B.n226 B.n225 585
R1084 B.n224 B.n223 585
R1085 B.n222 B.n221 585
R1086 B.n220 B.n219 585
R1087 B.n218 B.n217 585
R1088 B.n216 B.n215 585
R1089 B.n214 B.n213 585
R1090 B.n212 B.n211 585
R1091 B.n210 B.n209 585
R1092 B.n208 B.n207 585
R1093 B.n206 B.n205 585
R1094 B.n204 B.n203 585
R1095 B.n202 B.n201 585
R1096 B.n200 B.n199 585
R1097 B.n198 B.n197 585
R1098 B.n196 B.n195 585
R1099 B.n194 B.n193 585
R1100 B.n192 B.n191 585
R1101 B.n190 B.n189 585
R1102 B.n188 B.n187 585
R1103 B.n186 B.n185 585
R1104 B.n184 B.n183 585
R1105 B.n182 B.n181 585
R1106 B.n180 B.n179 585
R1107 B.n178 B.n177 585
R1108 B.n176 B.n175 585
R1109 B.n174 B.n173 585
R1110 B.n172 B.n171 585
R1111 B.n170 B.n169 585
R1112 B.n168 B.n167 585
R1113 B.n166 B.n165 585
R1114 B.n164 B.n163 585
R1115 B.n162 B.n161 585
R1116 B.n160 B.n159 585
R1117 B.n158 B.n157 585
R1118 B.n156 B.n155 585
R1119 B.n154 B.n153 585
R1120 B.n152 B.n151 585
R1121 B.n150 B.n149 585
R1122 B.n148 B.n147 585
R1123 B.n985 B.n76 585
R1124 B.n989 B.n76 585
R1125 B.n984 B.n75 585
R1126 B.n990 B.n75 585
R1127 B.n983 B.n982 585
R1128 B.n982 B.n71 585
R1129 B.n981 B.n70 585
R1130 B.n996 B.n70 585
R1131 B.n980 B.n69 585
R1132 B.n997 B.n69 585
R1133 B.n979 B.n68 585
R1134 B.n998 B.n68 585
R1135 B.n978 B.n977 585
R1136 B.n977 B.n64 585
R1137 B.n976 B.n63 585
R1138 B.n1004 B.n63 585
R1139 B.n975 B.n62 585
R1140 B.n1005 B.n62 585
R1141 B.n974 B.n61 585
R1142 B.n1006 B.n61 585
R1143 B.n973 B.n972 585
R1144 B.n972 B.n57 585
R1145 B.n971 B.n56 585
R1146 B.n1012 B.n56 585
R1147 B.n970 B.n55 585
R1148 B.n1013 B.n55 585
R1149 B.n969 B.n54 585
R1150 B.n1014 B.n54 585
R1151 B.n968 B.n967 585
R1152 B.n967 B.n50 585
R1153 B.n966 B.n49 585
R1154 B.n1020 B.n49 585
R1155 B.n965 B.n48 585
R1156 B.n1021 B.n48 585
R1157 B.n964 B.n47 585
R1158 B.n1022 B.n47 585
R1159 B.n963 B.n962 585
R1160 B.n962 B.n46 585
R1161 B.n961 B.n42 585
R1162 B.n1028 B.n42 585
R1163 B.n960 B.n41 585
R1164 B.n1029 B.n41 585
R1165 B.n959 B.n40 585
R1166 B.n1030 B.n40 585
R1167 B.n958 B.n957 585
R1168 B.n957 B.n36 585
R1169 B.n956 B.n35 585
R1170 B.n1036 B.n35 585
R1171 B.n955 B.n34 585
R1172 B.n1037 B.n34 585
R1173 B.n954 B.n33 585
R1174 B.n1038 B.n33 585
R1175 B.n953 B.n952 585
R1176 B.n952 B.n29 585
R1177 B.n951 B.n28 585
R1178 B.n1044 B.n28 585
R1179 B.n950 B.n27 585
R1180 B.n1045 B.n27 585
R1181 B.n949 B.n26 585
R1182 B.n1046 B.n26 585
R1183 B.n948 B.n947 585
R1184 B.n947 B.n22 585
R1185 B.n946 B.n21 585
R1186 B.n1052 B.n21 585
R1187 B.n945 B.n20 585
R1188 B.n1053 B.n20 585
R1189 B.n944 B.n19 585
R1190 B.n1054 B.n19 585
R1191 B.n943 B.n942 585
R1192 B.n942 B.n15 585
R1193 B.n941 B.n14 585
R1194 B.n1060 B.n14 585
R1195 B.n940 B.n13 585
R1196 B.n1061 B.n13 585
R1197 B.n939 B.n12 585
R1198 B.n1062 B.n12 585
R1199 B.n938 B.n937 585
R1200 B.n937 B.n8 585
R1201 B.n936 B.n7 585
R1202 B.n1068 B.n7 585
R1203 B.n935 B.n6 585
R1204 B.n1069 B.n6 585
R1205 B.n934 B.n5 585
R1206 B.n1070 B.n5 585
R1207 B.n933 B.n932 585
R1208 B.n932 B.n4 585
R1209 B.n931 B.n403 585
R1210 B.n931 B.n930 585
R1211 B.n921 B.n404 585
R1212 B.n405 B.n404 585
R1213 B.n923 B.n922 585
R1214 B.n924 B.n923 585
R1215 B.n920 B.n410 585
R1216 B.n410 B.n409 585
R1217 B.n919 B.n918 585
R1218 B.n918 B.n917 585
R1219 B.n412 B.n411 585
R1220 B.n413 B.n412 585
R1221 B.n910 B.n909 585
R1222 B.n911 B.n910 585
R1223 B.n908 B.n418 585
R1224 B.n418 B.n417 585
R1225 B.n907 B.n906 585
R1226 B.n906 B.n905 585
R1227 B.n420 B.n419 585
R1228 B.n421 B.n420 585
R1229 B.n898 B.n897 585
R1230 B.n899 B.n898 585
R1231 B.n896 B.n426 585
R1232 B.n426 B.n425 585
R1233 B.n895 B.n894 585
R1234 B.n894 B.n893 585
R1235 B.n428 B.n427 585
R1236 B.n429 B.n428 585
R1237 B.n886 B.n885 585
R1238 B.n887 B.n886 585
R1239 B.n884 B.n434 585
R1240 B.n434 B.n433 585
R1241 B.n883 B.n882 585
R1242 B.n882 B.n881 585
R1243 B.n436 B.n435 585
R1244 B.n437 B.n436 585
R1245 B.n874 B.n873 585
R1246 B.n875 B.n874 585
R1247 B.n872 B.n442 585
R1248 B.n442 B.n441 585
R1249 B.n871 B.n870 585
R1250 B.n870 B.n869 585
R1251 B.n444 B.n443 585
R1252 B.n862 B.n444 585
R1253 B.n861 B.n860 585
R1254 B.n863 B.n861 585
R1255 B.n859 B.n449 585
R1256 B.n449 B.n448 585
R1257 B.n858 B.n857 585
R1258 B.n857 B.n856 585
R1259 B.n451 B.n450 585
R1260 B.n452 B.n451 585
R1261 B.n849 B.n848 585
R1262 B.n850 B.n849 585
R1263 B.n847 B.n457 585
R1264 B.n457 B.n456 585
R1265 B.n846 B.n845 585
R1266 B.n845 B.n844 585
R1267 B.n459 B.n458 585
R1268 B.n460 B.n459 585
R1269 B.n837 B.n836 585
R1270 B.n838 B.n837 585
R1271 B.n835 B.n465 585
R1272 B.n465 B.n464 585
R1273 B.n834 B.n833 585
R1274 B.n833 B.n832 585
R1275 B.n467 B.n466 585
R1276 B.n468 B.n467 585
R1277 B.n825 B.n824 585
R1278 B.n826 B.n825 585
R1279 B.n823 B.n473 585
R1280 B.n473 B.n472 585
R1281 B.n822 B.n821 585
R1282 B.n821 B.n820 585
R1283 B.n475 B.n474 585
R1284 B.n476 B.n475 585
R1285 B.n813 B.n812 585
R1286 B.n814 B.n813 585
R1287 B.n811 B.n481 585
R1288 B.n481 B.n480 585
R1289 B.n805 B.n804 585
R1290 B.n803 B.n547 585
R1291 B.n802 B.n546 585
R1292 B.n807 B.n546 585
R1293 B.n801 B.n800 585
R1294 B.n799 B.n798 585
R1295 B.n797 B.n796 585
R1296 B.n795 B.n794 585
R1297 B.n793 B.n792 585
R1298 B.n791 B.n790 585
R1299 B.n789 B.n788 585
R1300 B.n787 B.n786 585
R1301 B.n785 B.n784 585
R1302 B.n783 B.n782 585
R1303 B.n781 B.n780 585
R1304 B.n779 B.n778 585
R1305 B.n777 B.n776 585
R1306 B.n775 B.n774 585
R1307 B.n773 B.n772 585
R1308 B.n771 B.n770 585
R1309 B.n769 B.n768 585
R1310 B.n767 B.n766 585
R1311 B.n765 B.n764 585
R1312 B.n763 B.n762 585
R1313 B.n761 B.n760 585
R1314 B.n759 B.n758 585
R1315 B.n757 B.n756 585
R1316 B.n755 B.n754 585
R1317 B.n753 B.n752 585
R1318 B.n751 B.n750 585
R1319 B.n749 B.n748 585
R1320 B.n747 B.n746 585
R1321 B.n745 B.n744 585
R1322 B.n743 B.n742 585
R1323 B.n741 B.n740 585
R1324 B.n739 B.n738 585
R1325 B.n737 B.n736 585
R1326 B.n735 B.n734 585
R1327 B.n733 B.n732 585
R1328 B.n731 B.n730 585
R1329 B.n729 B.n728 585
R1330 B.n727 B.n726 585
R1331 B.n725 B.n724 585
R1332 B.n723 B.n722 585
R1333 B.n721 B.n720 585
R1334 B.n719 B.n718 585
R1335 B.n717 B.n716 585
R1336 B.n715 B.n714 585
R1337 B.n713 B.n712 585
R1338 B.n711 B.n710 585
R1339 B.n709 B.n708 585
R1340 B.n707 B.n706 585
R1341 B.n705 B.n704 585
R1342 B.n703 B.n702 585
R1343 B.n701 B.n700 585
R1344 B.n699 B.n698 585
R1345 B.n697 B.n696 585
R1346 B.n695 B.n694 585
R1347 B.n693 B.n692 585
R1348 B.n691 B.n690 585
R1349 B.n689 B.n688 585
R1350 B.n686 B.n685 585
R1351 B.n684 B.n683 585
R1352 B.n682 B.n681 585
R1353 B.n680 B.n679 585
R1354 B.n678 B.n677 585
R1355 B.n676 B.n675 585
R1356 B.n674 B.n673 585
R1357 B.n672 B.n671 585
R1358 B.n670 B.n669 585
R1359 B.n668 B.n667 585
R1360 B.n666 B.n665 585
R1361 B.n664 B.n663 585
R1362 B.n662 B.n661 585
R1363 B.n660 B.n659 585
R1364 B.n658 B.n657 585
R1365 B.n656 B.n655 585
R1366 B.n654 B.n653 585
R1367 B.n652 B.n651 585
R1368 B.n650 B.n649 585
R1369 B.n648 B.n647 585
R1370 B.n646 B.n645 585
R1371 B.n644 B.n643 585
R1372 B.n642 B.n641 585
R1373 B.n640 B.n639 585
R1374 B.n638 B.n637 585
R1375 B.n636 B.n635 585
R1376 B.n634 B.n633 585
R1377 B.n632 B.n631 585
R1378 B.n630 B.n629 585
R1379 B.n628 B.n627 585
R1380 B.n626 B.n625 585
R1381 B.n624 B.n623 585
R1382 B.n622 B.n621 585
R1383 B.n620 B.n619 585
R1384 B.n618 B.n617 585
R1385 B.n616 B.n615 585
R1386 B.n614 B.n613 585
R1387 B.n612 B.n611 585
R1388 B.n610 B.n609 585
R1389 B.n608 B.n607 585
R1390 B.n606 B.n605 585
R1391 B.n604 B.n603 585
R1392 B.n602 B.n601 585
R1393 B.n600 B.n599 585
R1394 B.n598 B.n597 585
R1395 B.n596 B.n595 585
R1396 B.n594 B.n593 585
R1397 B.n592 B.n591 585
R1398 B.n590 B.n589 585
R1399 B.n588 B.n587 585
R1400 B.n586 B.n585 585
R1401 B.n584 B.n583 585
R1402 B.n582 B.n581 585
R1403 B.n580 B.n579 585
R1404 B.n578 B.n577 585
R1405 B.n576 B.n575 585
R1406 B.n574 B.n573 585
R1407 B.n572 B.n571 585
R1408 B.n570 B.n569 585
R1409 B.n568 B.n567 585
R1410 B.n566 B.n565 585
R1411 B.n564 B.n563 585
R1412 B.n562 B.n561 585
R1413 B.n560 B.n559 585
R1414 B.n558 B.n557 585
R1415 B.n556 B.n555 585
R1416 B.n554 B.n553 585
R1417 B.n483 B.n482 585
R1418 B.n810 B.n809 585
R1419 B.n479 B.n478 585
R1420 B.n480 B.n479 585
R1421 B.n816 B.n815 585
R1422 B.n815 B.n814 585
R1423 B.n817 B.n477 585
R1424 B.n477 B.n476 585
R1425 B.n819 B.n818 585
R1426 B.n820 B.n819 585
R1427 B.n471 B.n470 585
R1428 B.n472 B.n471 585
R1429 B.n828 B.n827 585
R1430 B.n827 B.n826 585
R1431 B.n829 B.n469 585
R1432 B.n469 B.n468 585
R1433 B.n831 B.n830 585
R1434 B.n832 B.n831 585
R1435 B.n463 B.n462 585
R1436 B.n464 B.n463 585
R1437 B.n840 B.n839 585
R1438 B.n839 B.n838 585
R1439 B.n841 B.n461 585
R1440 B.n461 B.n460 585
R1441 B.n843 B.n842 585
R1442 B.n844 B.n843 585
R1443 B.n455 B.n454 585
R1444 B.n456 B.n455 585
R1445 B.n852 B.n851 585
R1446 B.n851 B.n850 585
R1447 B.n853 B.n453 585
R1448 B.n453 B.n452 585
R1449 B.n855 B.n854 585
R1450 B.n856 B.n855 585
R1451 B.n447 B.n446 585
R1452 B.n448 B.n447 585
R1453 B.n865 B.n864 585
R1454 B.n864 B.n863 585
R1455 B.n866 B.n445 585
R1456 B.n862 B.n445 585
R1457 B.n868 B.n867 585
R1458 B.n869 B.n868 585
R1459 B.n440 B.n439 585
R1460 B.n441 B.n440 585
R1461 B.n877 B.n876 585
R1462 B.n876 B.n875 585
R1463 B.n878 B.n438 585
R1464 B.n438 B.n437 585
R1465 B.n880 B.n879 585
R1466 B.n881 B.n880 585
R1467 B.n432 B.n431 585
R1468 B.n433 B.n432 585
R1469 B.n889 B.n888 585
R1470 B.n888 B.n887 585
R1471 B.n890 B.n430 585
R1472 B.n430 B.n429 585
R1473 B.n892 B.n891 585
R1474 B.n893 B.n892 585
R1475 B.n424 B.n423 585
R1476 B.n425 B.n424 585
R1477 B.n901 B.n900 585
R1478 B.n900 B.n899 585
R1479 B.n902 B.n422 585
R1480 B.n422 B.n421 585
R1481 B.n904 B.n903 585
R1482 B.n905 B.n904 585
R1483 B.n416 B.n415 585
R1484 B.n417 B.n416 585
R1485 B.n913 B.n912 585
R1486 B.n912 B.n911 585
R1487 B.n914 B.n414 585
R1488 B.n414 B.n413 585
R1489 B.n916 B.n915 585
R1490 B.n917 B.n916 585
R1491 B.n408 B.n407 585
R1492 B.n409 B.n408 585
R1493 B.n926 B.n925 585
R1494 B.n925 B.n924 585
R1495 B.n927 B.n406 585
R1496 B.n406 B.n405 585
R1497 B.n929 B.n928 585
R1498 B.n930 B.n929 585
R1499 B.n2 B.n0 585
R1500 B.n4 B.n2 585
R1501 B.n3 B.n1 585
R1502 B.n1069 B.n3 585
R1503 B.n1067 B.n1066 585
R1504 B.n1068 B.n1067 585
R1505 B.n1065 B.n9 585
R1506 B.n9 B.n8 585
R1507 B.n1064 B.n1063 585
R1508 B.n1063 B.n1062 585
R1509 B.n11 B.n10 585
R1510 B.n1061 B.n11 585
R1511 B.n1059 B.n1058 585
R1512 B.n1060 B.n1059 585
R1513 B.n1057 B.n16 585
R1514 B.n16 B.n15 585
R1515 B.n1056 B.n1055 585
R1516 B.n1055 B.n1054 585
R1517 B.n18 B.n17 585
R1518 B.n1053 B.n18 585
R1519 B.n1051 B.n1050 585
R1520 B.n1052 B.n1051 585
R1521 B.n1049 B.n23 585
R1522 B.n23 B.n22 585
R1523 B.n1048 B.n1047 585
R1524 B.n1047 B.n1046 585
R1525 B.n25 B.n24 585
R1526 B.n1045 B.n25 585
R1527 B.n1043 B.n1042 585
R1528 B.n1044 B.n1043 585
R1529 B.n1041 B.n30 585
R1530 B.n30 B.n29 585
R1531 B.n1040 B.n1039 585
R1532 B.n1039 B.n1038 585
R1533 B.n32 B.n31 585
R1534 B.n1037 B.n32 585
R1535 B.n1035 B.n1034 585
R1536 B.n1036 B.n1035 585
R1537 B.n1033 B.n37 585
R1538 B.n37 B.n36 585
R1539 B.n1032 B.n1031 585
R1540 B.n1031 B.n1030 585
R1541 B.n39 B.n38 585
R1542 B.n1029 B.n39 585
R1543 B.n1027 B.n1026 585
R1544 B.n1028 B.n1027 585
R1545 B.n1025 B.n43 585
R1546 B.n46 B.n43 585
R1547 B.n1024 B.n1023 585
R1548 B.n1023 B.n1022 585
R1549 B.n45 B.n44 585
R1550 B.n1021 B.n45 585
R1551 B.n1019 B.n1018 585
R1552 B.n1020 B.n1019 585
R1553 B.n1017 B.n51 585
R1554 B.n51 B.n50 585
R1555 B.n1016 B.n1015 585
R1556 B.n1015 B.n1014 585
R1557 B.n53 B.n52 585
R1558 B.n1013 B.n53 585
R1559 B.n1011 B.n1010 585
R1560 B.n1012 B.n1011 585
R1561 B.n1009 B.n58 585
R1562 B.n58 B.n57 585
R1563 B.n1008 B.n1007 585
R1564 B.n1007 B.n1006 585
R1565 B.n60 B.n59 585
R1566 B.n1005 B.n60 585
R1567 B.n1003 B.n1002 585
R1568 B.n1004 B.n1003 585
R1569 B.n1001 B.n65 585
R1570 B.n65 B.n64 585
R1571 B.n1000 B.n999 585
R1572 B.n999 B.n998 585
R1573 B.n67 B.n66 585
R1574 B.n997 B.n67 585
R1575 B.n995 B.n994 585
R1576 B.n996 B.n995 585
R1577 B.n993 B.n72 585
R1578 B.n72 B.n71 585
R1579 B.n992 B.n991 585
R1580 B.n991 B.n990 585
R1581 B.n74 B.n73 585
R1582 B.n989 B.n74 585
R1583 B.n1072 B.n1071 585
R1584 B.n1071 B.n1070 585
R1585 B.n550 B.t16 440.56
R1586 B.n548 B.t19 440.56
R1587 B.n144 B.t11 440.56
R1588 B.n142 B.t8 440.56
R1589 B.n805 B.n479 434.841
R1590 B.n147 B.n74 434.841
R1591 B.n809 B.n481 434.841
R1592 B.n987 B.n76 434.841
R1593 B.n551 B.t15 386.644
R1594 B.n143 B.t9 386.644
R1595 B.n549 B.t18 386.644
R1596 B.n145 B.t12 386.644
R1597 B.n550 B.t13 385.658
R1598 B.n548 B.t17 385.658
R1599 B.n144 B.t10 385.658
R1600 B.n142 B.t6 385.658
R1601 B.n988 B.n140 256.663
R1602 B.n988 B.n139 256.663
R1603 B.n988 B.n138 256.663
R1604 B.n988 B.n137 256.663
R1605 B.n988 B.n136 256.663
R1606 B.n988 B.n135 256.663
R1607 B.n988 B.n134 256.663
R1608 B.n988 B.n133 256.663
R1609 B.n988 B.n132 256.663
R1610 B.n988 B.n131 256.663
R1611 B.n988 B.n130 256.663
R1612 B.n988 B.n129 256.663
R1613 B.n988 B.n128 256.663
R1614 B.n988 B.n127 256.663
R1615 B.n988 B.n126 256.663
R1616 B.n988 B.n125 256.663
R1617 B.n988 B.n124 256.663
R1618 B.n988 B.n123 256.663
R1619 B.n988 B.n122 256.663
R1620 B.n988 B.n121 256.663
R1621 B.n988 B.n120 256.663
R1622 B.n988 B.n119 256.663
R1623 B.n988 B.n118 256.663
R1624 B.n988 B.n117 256.663
R1625 B.n988 B.n116 256.663
R1626 B.n988 B.n115 256.663
R1627 B.n988 B.n114 256.663
R1628 B.n988 B.n113 256.663
R1629 B.n988 B.n112 256.663
R1630 B.n988 B.n111 256.663
R1631 B.n988 B.n110 256.663
R1632 B.n988 B.n109 256.663
R1633 B.n988 B.n108 256.663
R1634 B.n988 B.n107 256.663
R1635 B.n988 B.n106 256.663
R1636 B.n988 B.n105 256.663
R1637 B.n988 B.n104 256.663
R1638 B.n988 B.n103 256.663
R1639 B.n988 B.n102 256.663
R1640 B.n988 B.n101 256.663
R1641 B.n988 B.n100 256.663
R1642 B.n988 B.n99 256.663
R1643 B.n988 B.n98 256.663
R1644 B.n988 B.n97 256.663
R1645 B.n988 B.n96 256.663
R1646 B.n988 B.n95 256.663
R1647 B.n988 B.n94 256.663
R1648 B.n988 B.n93 256.663
R1649 B.n988 B.n92 256.663
R1650 B.n988 B.n91 256.663
R1651 B.n988 B.n90 256.663
R1652 B.n988 B.n89 256.663
R1653 B.n988 B.n88 256.663
R1654 B.n988 B.n87 256.663
R1655 B.n988 B.n86 256.663
R1656 B.n988 B.n85 256.663
R1657 B.n988 B.n84 256.663
R1658 B.n988 B.n83 256.663
R1659 B.n988 B.n82 256.663
R1660 B.n988 B.n81 256.663
R1661 B.n988 B.n80 256.663
R1662 B.n988 B.n79 256.663
R1663 B.n988 B.n78 256.663
R1664 B.n988 B.n77 256.663
R1665 B.n807 B.n806 256.663
R1666 B.n807 B.n484 256.663
R1667 B.n807 B.n485 256.663
R1668 B.n807 B.n486 256.663
R1669 B.n807 B.n487 256.663
R1670 B.n807 B.n488 256.663
R1671 B.n807 B.n489 256.663
R1672 B.n807 B.n490 256.663
R1673 B.n807 B.n491 256.663
R1674 B.n807 B.n492 256.663
R1675 B.n807 B.n493 256.663
R1676 B.n807 B.n494 256.663
R1677 B.n807 B.n495 256.663
R1678 B.n807 B.n496 256.663
R1679 B.n807 B.n497 256.663
R1680 B.n807 B.n498 256.663
R1681 B.n807 B.n499 256.663
R1682 B.n807 B.n500 256.663
R1683 B.n807 B.n501 256.663
R1684 B.n807 B.n502 256.663
R1685 B.n807 B.n503 256.663
R1686 B.n807 B.n504 256.663
R1687 B.n807 B.n505 256.663
R1688 B.n807 B.n506 256.663
R1689 B.n807 B.n507 256.663
R1690 B.n807 B.n508 256.663
R1691 B.n807 B.n509 256.663
R1692 B.n807 B.n510 256.663
R1693 B.n807 B.n511 256.663
R1694 B.n807 B.n512 256.663
R1695 B.n807 B.n513 256.663
R1696 B.n807 B.n514 256.663
R1697 B.n807 B.n515 256.663
R1698 B.n807 B.n516 256.663
R1699 B.n807 B.n517 256.663
R1700 B.n807 B.n518 256.663
R1701 B.n807 B.n519 256.663
R1702 B.n807 B.n520 256.663
R1703 B.n807 B.n521 256.663
R1704 B.n807 B.n522 256.663
R1705 B.n807 B.n523 256.663
R1706 B.n807 B.n524 256.663
R1707 B.n807 B.n525 256.663
R1708 B.n807 B.n526 256.663
R1709 B.n807 B.n527 256.663
R1710 B.n807 B.n528 256.663
R1711 B.n807 B.n529 256.663
R1712 B.n807 B.n530 256.663
R1713 B.n807 B.n531 256.663
R1714 B.n807 B.n532 256.663
R1715 B.n807 B.n533 256.663
R1716 B.n807 B.n534 256.663
R1717 B.n807 B.n535 256.663
R1718 B.n807 B.n536 256.663
R1719 B.n807 B.n537 256.663
R1720 B.n807 B.n538 256.663
R1721 B.n807 B.n539 256.663
R1722 B.n807 B.n540 256.663
R1723 B.n807 B.n541 256.663
R1724 B.n807 B.n542 256.663
R1725 B.n807 B.n543 256.663
R1726 B.n807 B.n544 256.663
R1727 B.n807 B.n545 256.663
R1728 B.n808 B.n807 256.663
R1729 B.n815 B.n479 163.367
R1730 B.n815 B.n477 163.367
R1731 B.n819 B.n477 163.367
R1732 B.n819 B.n471 163.367
R1733 B.n827 B.n471 163.367
R1734 B.n827 B.n469 163.367
R1735 B.n831 B.n469 163.367
R1736 B.n831 B.n463 163.367
R1737 B.n839 B.n463 163.367
R1738 B.n839 B.n461 163.367
R1739 B.n843 B.n461 163.367
R1740 B.n843 B.n455 163.367
R1741 B.n851 B.n455 163.367
R1742 B.n851 B.n453 163.367
R1743 B.n855 B.n453 163.367
R1744 B.n855 B.n447 163.367
R1745 B.n864 B.n447 163.367
R1746 B.n864 B.n445 163.367
R1747 B.n868 B.n445 163.367
R1748 B.n868 B.n440 163.367
R1749 B.n876 B.n440 163.367
R1750 B.n876 B.n438 163.367
R1751 B.n880 B.n438 163.367
R1752 B.n880 B.n432 163.367
R1753 B.n888 B.n432 163.367
R1754 B.n888 B.n430 163.367
R1755 B.n892 B.n430 163.367
R1756 B.n892 B.n424 163.367
R1757 B.n900 B.n424 163.367
R1758 B.n900 B.n422 163.367
R1759 B.n904 B.n422 163.367
R1760 B.n904 B.n416 163.367
R1761 B.n912 B.n416 163.367
R1762 B.n912 B.n414 163.367
R1763 B.n916 B.n414 163.367
R1764 B.n916 B.n408 163.367
R1765 B.n925 B.n408 163.367
R1766 B.n925 B.n406 163.367
R1767 B.n929 B.n406 163.367
R1768 B.n929 B.n2 163.367
R1769 B.n1071 B.n2 163.367
R1770 B.n1071 B.n3 163.367
R1771 B.n1067 B.n3 163.367
R1772 B.n1067 B.n9 163.367
R1773 B.n1063 B.n9 163.367
R1774 B.n1063 B.n11 163.367
R1775 B.n1059 B.n11 163.367
R1776 B.n1059 B.n16 163.367
R1777 B.n1055 B.n16 163.367
R1778 B.n1055 B.n18 163.367
R1779 B.n1051 B.n18 163.367
R1780 B.n1051 B.n23 163.367
R1781 B.n1047 B.n23 163.367
R1782 B.n1047 B.n25 163.367
R1783 B.n1043 B.n25 163.367
R1784 B.n1043 B.n30 163.367
R1785 B.n1039 B.n30 163.367
R1786 B.n1039 B.n32 163.367
R1787 B.n1035 B.n32 163.367
R1788 B.n1035 B.n37 163.367
R1789 B.n1031 B.n37 163.367
R1790 B.n1031 B.n39 163.367
R1791 B.n1027 B.n39 163.367
R1792 B.n1027 B.n43 163.367
R1793 B.n1023 B.n43 163.367
R1794 B.n1023 B.n45 163.367
R1795 B.n1019 B.n45 163.367
R1796 B.n1019 B.n51 163.367
R1797 B.n1015 B.n51 163.367
R1798 B.n1015 B.n53 163.367
R1799 B.n1011 B.n53 163.367
R1800 B.n1011 B.n58 163.367
R1801 B.n1007 B.n58 163.367
R1802 B.n1007 B.n60 163.367
R1803 B.n1003 B.n60 163.367
R1804 B.n1003 B.n65 163.367
R1805 B.n999 B.n65 163.367
R1806 B.n999 B.n67 163.367
R1807 B.n995 B.n67 163.367
R1808 B.n995 B.n72 163.367
R1809 B.n991 B.n72 163.367
R1810 B.n991 B.n74 163.367
R1811 B.n547 B.n546 163.367
R1812 B.n800 B.n546 163.367
R1813 B.n798 B.n797 163.367
R1814 B.n794 B.n793 163.367
R1815 B.n790 B.n789 163.367
R1816 B.n786 B.n785 163.367
R1817 B.n782 B.n781 163.367
R1818 B.n778 B.n777 163.367
R1819 B.n774 B.n773 163.367
R1820 B.n770 B.n769 163.367
R1821 B.n766 B.n765 163.367
R1822 B.n762 B.n761 163.367
R1823 B.n758 B.n757 163.367
R1824 B.n754 B.n753 163.367
R1825 B.n750 B.n749 163.367
R1826 B.n746 B.n745 163.367
R1827 B.n742 B.n741 163.367
R1828 B.n738 B.n737 163.367
R1829 B.n734 B.n733 163.367
R1830 B.n730 B.n729 163.367
R1831 B.n726 B.n725 163.367
R1832 B.n722 B.n721 163.367
R1833 B.n718 B.n717 163.367
R1834 B.n714 B.n713 163.367
R1835 B.n710 B.n709 163.367
R1836 B.n706 B.n705 163.367
R1837 B.n702 B.n701 163.367
R1838 B.n698 B.n697 163.367
R1839 B.n694 B.n693 163.367
R1840 B.n690 B.n689 163.367
R1841 B.n685 B.n684 163.367
R1842 B.n681 B.n680 163.367
R1843 B.n677 B.n676 163.367
R1844 B.n673 B.n672 163.367
R1845 B.n669 B.n668 163.367
R1846 B.n665 B.n664 163.367
R1847 B.n661 B.n660 163.367
R1848 B.n657 B.n656 163.367
R1849 B.n653 B.n652 163.367
R1850 B.n649 B.n648 163.367
R1851 B.n645 B.n644 163.367
R1852 B.n641 B.n640 163.367
R1853 B.n637 B.n636 163.367
R1854 B.n633 B.n632 163.367
R1855 B.n629 B.n628 163.367
R1856 B.n625 B.n624 163.367
R1857 B.n621 B.n620 163.367
R1858 B.n617 B.n616 163.367
R1859 B.n613 B.n612 163.367
R1860 B.n609 B.n608 163.367
R1861 B.n605 B.n604 163.367
R1862 B.n601 B.n600 163.367
R1863 B.n597 B.n596 163.367
R1864 B.n593 B.n592 163.367
R1865 B.n589 B.n588 163.367
R1866 B.n585 B.n584 163.367
R1867 B.n581 B.n580 163.367
R1868 B.n577 B.n576 163.367
R1869 B.n573 B.n572 163.367
R1870 B.n569 B.n568 163.367
R1871 B.n565 B.n564 163.367
R1872 B.n561 B.n560 163.367
R1873 B.n557 B.n556 163.367
R1874 B.n553 B.n483 163.367
R1875 B.n813 B.n481 163.367
R1876 B.n813 B.n475 163.367
R1877 B.n821 B.n475 163.367
R1878 B.n821 B.n473 163.367
R1879 B.n825 B.n473 163.367
R1880 B.n825 B.n467 163.367
R1881 B.n833 B.n467 163.367
R1882 B.n833 B.n465 163.367
R1883 B.n837 B.n465 163.367
R1884 B.n837 B.n459 163.367
R1885 B.n845 B.n459 163.367
R1886 B.n845 B.n457 163.367
R1887 B.n849 B.n457 163.367
R1888 B.n849 B.n451 163.367
R1889 B.n857 B.n451 163.367
R1890 B.n857 B.n449 163.367
R1891 B.n861 B.n449 163.367
R1892 B.n861 B.n444 163.367
R1893 B.n870 B.n444 163.367
R1894 B.n870 B.n442 163.367
R1895 B.n874 B.n442 163.367
R1896 B.n874 B.n436 163.367
R1897 B.n882 B.n436 163.367
R1898 B.n882 B.n434 163.367
R1899 B.n886 B.n434 163.367
R1900 B.n886 B.n428 163.367
R1901 B.n894 B.n428 163.367
R1902 B.n894 B.n426 163.367
R1903 B.n898 B.n426 163.367
R1904 B.n898 B.n420 163.367
R1905 B.n906 B.n420 163.367
R1906 B.n906 B.n418 163.367
R1907 B.n910 B.n418 163.367
R1908 B.n910 B.n412 163.367
R1909 B.n918 B.n412 163.367
R1910 B.n918 B.n410 163.367
R1911 B.n923 B.n410 163.367
R1912 B.n923 B.n404 163.367
R1913 B.n931 B.n404 163.367
R1914 B.n932 B.n931 163.367
R1915 B.n932 B.n5 163.367
R1916 B.n6 B.n5 163.367
R1917 B.n7 B.n6 163.367
R1918 B.n937 B.n7 163.367
R1919 B.n937 B.n12 163.367
R1920 B.n13 B.n12 163.367
R1921 B.n14 B.n13 163.367
R1922 B.n942 B.n14 163.367
R1923 B.n942 B.n19 163.367
R1924 B.n20 B.n19 163.367
R1925 B.n21 B.n20 163.367
R1926 B.n947 B.n21 163.367
R1927 B.n947 B.n26 163.367
R1928 B.n27 B.n26 163.367
R1929 B.n28 B.n27 163.367
R1930 B.n952 B.n28 163.367
R1931 B.n952 B.n33 163.367
R1932 B.n34 B.n33 163.367
R1933 B.n35 B.n34 163.367
R1934 B.n957 B.n35 163.367
R1935 B.n957 B.n40 163.367
R1936 B.n41 B.n40 163.367
R1937 B.n42 B.n41 163.367
R1938 B.n962 B.n42 163.367
R1939 B.n962 B.n47 163.367
R1940 B.n48 B.n47 163.367
R1941 B.n49 B.n48 163.367
R1942 B.n967 B.n49 163.367
R1943 B.n967 B.n54 163.367
R1944 B.n55 B.n54 163.367
R1945 B.n56 B.n55 163.367
R1946 B.n972 B.n56 163.367
R1947 B.n972 B.n61 163.367
R1948 B.n62 B.n61 163.367
R1949 B.n63 B.n62 163.367
R1950 B.n977 B.n63 163.367
R1951 B.n977 B.n68 163.367
R1952 B.n69 B.n68 163.367
R1953 B.n70 B.n69 163.367
R1954 B.n982 B.n70 163.367
R1955 B.n982 B.n75 163.367
R1956 B.n76 B.n75 163.367
R1957 B.n151 B.n150 163.367
R1958 B.n155 B.n154 163.367
R1959 B.n159 B.n158 163.367
R1960 B.n163 B.n162 163.367
R1961 B.n167 B.n166 163.367
R1962 B.n171 B.n170 163.367
R1963 B.n175 B.n174 163.367
R1964 B.n179 B.n178 163.367
R1965 B.n183 B.n182 163.367
R1966 B.n187 B.n186 163.367
R1967 B.n191 B.n190 163.367
R1968 B.n195 B.n194 163.367
R1969 B.n199 B.n198 163.367
R1970 B.n203 B.n202 163.367
R1971 B.n207 B.n206 163.367
R1972 B.n211 B.n210 163.367
R1973 B.n215 B.n214 163.367
R1974 B.n219 B.n218 163.367
R1975 B.n223 B.n222 163.367
R1976 B.n227 B.n226 163.367
R1977 B.n231 B.n230 163.367
R1978 B.n235 B.n234 163.367
R1979 B.n239 B.n238 163.367
R1980 B.n243 B.n242 163.367
R1981 B.n247 B.n246 163.367
R1982 B.n251 B.n250 163.367
R1983 B.n255 B.n254 163.367
R1984 B.n259 B.n258 163.367
R1985 B.n263 B.n262 163.367
R1986 B.n267 B.n266 163.367
R1987 B.n271 B.n270 163.367
R1988 B.n275 B.n274 163.367
R1989 B.n279 B.n278 163.367
R1990 B.n283 B.n282 163.367
R1991 B.n288 B.n287 163.367
R1992 B.n292 B.n291 163.367
R1993 B.n296 B.n295 163.367
R1994 B.n300 B.n299 163.367
R1995 B.n304 B.n303 163.367
R1996 B.n308 B.n307 163.367
R1997 B.n312 B.n311 163.367
R1998 B.n316 B.n315 163.367
R1999 B.n320 B.n319 163.367
R2000 B.n324 B.n323 163.367
R2001 B.n328 B.n327 163.367
R2002 B.n332 B.n331 163.367
R2003 B.n336 B.n335 163.367
R2004 B.n340 B.n339 163.367
R2005 B.n344 B.n343 163.367
R2006 B.n348 B.n347 163.367
R2007 B.n352 B.n351 163.367
R2008 B.n356 B.n355 163.367
R2009 B.n360 B.n359 163.367
R2010 B.n364 B.n363 163.367
R2011 B.n368 B.n367 163.367
R2012 B.n372 B.n371 163.367
R2013 B.n376 B.n375 163.367
R2014 B.n380 B.n379 163.367
R2015 B.n384 B.n383 163.367
R2016 B.n388 B.n387 163.367
R2017 B.n392 B.n391 163.367
R2018 B.n396 B.n395 163.367
R2019 B.n400 B.n399 163.367
R2020 B.n987 B.n141 163.367
R2021 B.n806 B.n805 71.676
R2022 B.n800 B.n484 71.676
R2023 B.n797 B.n485 71.676
R2024 B.n793 B.n486 71.676
R2025 B.n789 B.n487 71.676
R2026 B.n785 B.n488 71.676
R2027 B.n781 B.n489 71.676
R2028 B.n777 B.n490 71.676
R2029 B.n773 B.n491 71.676
R2030 B.n769 B.n492 71.676
R2031 B.n765 B.n493 71.676
R2032 B.n761 B.n494 71.676
R2033 B.n757 B.n495 71.676
R2034 B.n753 B.n496 71.676
R2035 B.n749 B.n497 71.676
R2036 B.n745 B.n498 71.676
R2037 B.n741 B.n499 71.676
R2038 B.n737 B.n500 71.676
R2039 B.n733 B.n501 71.676
R2040 B.n729 B.n502 71.676
R2041 B.n725 B.n503 71.676
R2042 B.n721 B.n504 71.676
R2043 B.n717 B.n505 71.676
R2044 B.n713 B.n506 71.676
R2045 B.n709 B.n507 71.676
R2046 B.n705 B.n508 71.676
R2047 B.n701 B.n509 71.676
R2048 B.n697 B.n510 71.676
R2049 B.n693 B.n511 71.676
R2050 B.n689 B.n512 71.676
R2051 B.n684 B.n513 71.676
R2052 B.n680 B.n514 71.676
R2053 B.n676 B.n515 71.676
R2054 B.n672 B.n516 71.676
R2055 B.n668 B.n517 71.676
R2056 B.n664 B.n518 71.676
R2057 B.n660 B.n519 71.676
R2058 B.n656 B.n520 71.676
R2059 B.n652 B.n521 71.676
R2060 B.n648 B.n522 71.676
R2061 B.n644 B.n523 71.676
R2062 B.n640 B.n524 71.676
R2063 B.n636 B.n525 71.676
R2064 B.n632 B.n526 71.676
R2065 B.n628 B.n527 71.676
R2066 B.n624 B.n528 71.676
R2067 B.n620 B.n529 71.676
R2068 B.n616 B.n530 71.676
R2069 B.n612 B.n531 71.676
R2070 B.n608 B.n532 71.676
R2071 B.n604 B.n533 71.676
R2072 B.n600 B.n534 71.676
R2073 B.n596 B.n535 71.676
R2074 B.n592 B.n536 71.676
R2075 B.n588 B.n537 71.676
R2076 B.n584 B.n538 71.676
R2077 B.n580 B.n539 71.676
R2078 B.n576 B.n540 71.676
R2079 B.n572 B.n541 71.676
R2080 B.n568 B.n542 71.676
R2081 B.n564 B.n543 71.676
R2082 B.n560 B.n544 71.676
R2083 B.n556 B.n545 71.676
R2084 B.n808 B.n483 71.676
R2085 B.n147 B.n77 71.676
R2086 B.n151 B.n78 71.676
R2087 B.n155 B.n79 71.676
R2088 B.n159 B.n80 71.676
R2089 B.n163 B.n81 71.676
R2090 B.n167 B.n82 71.676
R2091 B.n171 B.n83 71.676
R2092 B.n175 B.n84 71.676
R2093 B.n179 B.n85 71.676
R2094 B.n183 B.n86 71.676
R2095 B.n187 B.n87 71.676
R2096 B.n191 B.n88 71.676
R2097 B.n195 B.n89 71.676
R2098 B.n199 B.n90 71.676
R2099 B.n203 B.n91 71.676
R2100 B.n207 B.n92 71.676
R2101 B.n211 B.n93 71.676
R2102 B.n215 B.n94 71.676
R2103 B.n219 B.n95 71.676
R2104 B.n223 B.n96 71.676
R2105 B.n227 B.n97 71.676
R2106 B.n231 B.n98 71.676
R2107 B.n235 B.n99 71.676
R2108 B.n239 B.n100 71.676
R2109 B.n243 B.n101 71.676
R2110 B.n247 B.n102 71.676
R2111 B.n251 B.n103 71.676
R2112 B.n255 B.n104 71.676
R2113 B.n259 B.n105 71.676
R2114 B.n263 B.n106 71.676
R2115 B.n267 B.n107 71.676
R2116 B.n271 B.n108 71.676
R2117 B.n275 B.n109 71.676
R2118 B.n279 B.n110 71.676
R2119 B.n283 B.n111 71.676
R2120 B.n288 B.n112 71.676
R2121 B.n292 B.n113 71.676
R2122 B.n296 B.n114 71.676
R2123 B.n300 B.n115 71.676
R2124 B.n304 B.n116 71.676
R2125 B.n308 B.n117 71.676
R2126 B.n312 B.n118 71.676
R2127 B.n316 B.n119 71.676
R2128 B.n320 B.n120 71.676
R2129 B.n324 B.n121 71.676
R2130 B.n328 B.n122 71.676
R2131 B.n332 B.n123 71.676
R2132 B.n336 B.n124 71.676
R2133 B.n340 B.n125 71.676
R2134 B.n344 B.n126 71.676
R2135 B.n348 B.n127 71.676
R2136 B.n352 B.n128 71.676
R2137 B.n356 B.n129 71.676
R2138 B.n360 B.n130 71.676
R2139 B.n364 B.n131 71.676
R2140 B.n368 B.n132 71.676
R2141 B.n372 B.n133 71.676
R2142 B.n376 B.n134 71.676
R2143 B.n380 B.n135 71.676
R2144 B.n384 B.n136 71.676
R2145 B.n388 B.n137 71.676
R2146 B.n392 B.n138 71.676
R2147 B.n396 B.n139 71.676
R2148 B.n400 B.n140 71.676
R2149 B.n141 B.n140 71.676
R2150 B.n399 B.n139 71.676
R2151 B.n395 B.n138 71.676
R2152 B.n391 B.n137 71.676
R2153 B.n387 B.n136 71.676
R2154 B.n383 B.n135 71.676
R2155 B.n379 B.n134 71.676
R2156 B.n375 B.n133 71.676
R2157 B.n371 B.n132 71.676
R2158 B.n367 B.n131 71.676
R2159 B.n363 B.n130 71.676
R2160 B.n359 B.n129 71.676
R2161 B.n355 B.n128 71.676
R2162 B.n351 B.n127 71.676
R2163 B.n347 B.n126 71.676
R2164 B.n343 B.n125 71.676
R2165 B.n339 B.n124 71.676
R2166 B.n335 B.n123 71.676
R2167 B.n331 B.n122 71.676
R2168 B.n327 B.n121 71.676
R2169 B.n323 B.n120 71.676
R2170 B.n319 B.n119 71.676
R2171 B.n315 B.n118 71.676
R2172 B.n311 B.n117 71.676
R2173 B.n307 B.n116 71.676
R2174 B.n303 B.n115 71.676
R2175 B.n299 B.n114 71.676
R2176 B.n295 B.n113 71.676
R2177 B.n291 B.n112 71.676
R2178 B.n287 B.n111 71.676
R2179 B.n282 B.n110 71.676
R2180 B.n278 B.n109 71.676
R2181 B.n274 B.n108 71.676
R2182 B.n270 B.n107 71.676
R2183 B.n266 B.n106 71.676
R2184 B.n262 B.n105 71.676
R2185 B.n258 B.n104 71.676
R2186 B.n254 B.n103 71.676
R2187 B.n250 B.n102 71.676
R2188 B.n246 B.n101 71.676
R2189 B.n242 B.n100 71.676
R2190 B.n238 B.n99 71.676
R2191 B.n234 B.n98 71.676
R2192 B.n230 B.n97 71.676
R2193 B.n226 B.n96 71.676
R2194 B.n222 B.n95 71.676
R2195 B.n218 B.n94 71.676
R2196 B.n214 B.n93 71.676
R2197 B.n210 B.n92 71.676
R2198 B.n206 B.n91 71.676
R2199 B.n202 B.n90 71.676
R2200 B.n198 B.n89 71.676
R2201 B.n194 B.n88 71.676
R2202 B.n190 B.n87 71.676
R2203 B.n186 B.n86 71.676
R2204 B.n182 B.n85 71.676
R2205 B.n178 B.n84 71.676
R2206 B.n174 B.n83 71.676
R2207 B.n170 B.n82 71.676
R2208 B.n166 B.n81 71.676
R2209 B.n162 B.n80 71.676
R2210 B.n158 B.n79 71.676
R2211 B.n154 B.n78 71.676
R2212 B.n150 B.n77 71.676
R2213 B.n806 B.n547 71.676
R2214 B.n798 B.n484 71.676
R2215 B.n794 B.n485 71.676
R2216 B.n790 B.n486 71.676
R2217 B.n786 B.n487 71.676
R2218 B.n782 B.n488 71.676
R2219 B.n778 B.n489 71.676
R2220 B.n774 B.n490 71.676
R2221 B.n770 B.n491 71.676
R2222 B.n766 B.n492 71.676
R2223 B.n762 B.n493 71.676
R2224 B.n758 B.n494 71.676
R2225 B.n754 B.n495 71.676
R2226 B.n750 B.n496 71.676
R2227 B.n746 B.n497 71.676
R2228 B.n742 B.n498 71.676
R2229 B.n738 B.n499 71.676
R2230 B.n734 B.n500 71.676
R2231 B.n730 B.n501 71.676
R2232 B.n726 B.n502 71.676
R2233 B.n722 B.n503 71.676
R2234 B.n718 B.n504 71.676
R2235 B.n714 B.n505 71.676
R2236 B.n710 B.n506 71.676
R2237 B.n706 B.n507 71.676
R2238 B.n702 B.n508 71.676
R2239 B.n698 B.n509 71.676
R2240 B.n694 B.n510 71.676
R2241 B.n690 B.n511 71.676
R2242 B.n685 B.n512 71.676
R2243 B.n681 B.n513 71.676
R2244 B.n677 B.n514 71.676
R2245 B.n673 B.n515 71.676
R2246 B.n669 B.n516 71.676
R2247 B.n665 B.n517 71.676
R2248 B.n661 B.n518 71.676
R2249 B.n657 B.n519 71.676
R2250 B.n653 B.n520 71.676
R2251 B.n649 B.n521 71.676
R2252 B.n645 B.n522 71.676
R2253 B.n641 B.n523 71.676
R2254 B.n637 B.n524 71.676
R2255 B.n633 B.n525 71.676
R2256 B.n629 B.n526 71.676
R2257 B.n625 B.n527 71.676
R2258 B.n621 B.n528 71.676
R2259 B.n617 B.n529 71.676
R2260 B.n613 B.n530 71.676
R2261 B.n609 B.n531 71.676
R2262 B.n605 B.n532 71.676
R2263 B.n601 B.n533 71.676
R2264 B.n597 B.n534 71.676
R2265 B.n593 B.n535 71.676
R2266 B.n589 B.n536 71.676
R2267 B.n585 B.n537 71.676
R2268 B.n581 B.n538 71.676
R2269 B.n577 B.n539 71.676
R2270 B.n573 B.n540 71.676
R2271 B.n569 B.n541 71.676
R2272 B.n565 B.n542 71.676
R2273 B.n561 B.n543 71.676
R2274 B.n557 B.n544 71.676
R2275 B.n553 B.n545 71.676
R2276 B.n809 B.n808 71.676
R2277 B.n552 B.n551 59.5399
R2278 B.n687 B.n549 59.5399
R2279 B.n146 B.n145 59.5399
R2280 B.n285 B.n143 59.5399
R2281 B.n551 B.n550 53.9157
R2282 B.n549 B.n548 53.9157
R2283 B.n145 B.n144 53.9157
R2284 B.n143 B.n142 53.9157
R2285 B.n807 B.n480 52.2805
R2286 B.n989 B.n988 52.2805
R2287 B.n814 B.n480 32.0279
R2288 B.n814 B.n476 32.0279
R2289 B.n820 B.n476 32.0279
R2290 B.n820 B.n472 32.0279
R2291 B.n826 B.n472 32.0279
R2292 B.n826 B.n468 32.0279
R2293 B.n832 B.n468 32.0279
R2294 B.n838 B.n464 32.0279
R2295 B.n838 B.n460 32.0279
R2296 B.n844 B.n460 32.0279
R2297 B.n844 B.n456 32.0279
R2298 B.n850 B.n456 32.0279
R2299 B.n850 B.n452 32.0279
R2300 B.n856 B.n452 32.0279
R2301 B.n856 B.n448 32.0279
R2302 B.n863 B.n448 32.0279
R2303 B.n863 B.n862 32.0279
R2304 B.n869 B.n441 32.0279
R2305 B.n875 B.n441 32.0279
R2306 B.n875 B.n437 32.0279
R2307 B.n881 B.n437 32.0279
R2308 B.n881 B.n433 32.0279
R2309 B.n887 B.n433 32.0279
R2310 B.n887 B.n429 32.0279
R2311 B.n893 B.n429 32.0279
R2312 B.n899 B.n425 32.0279
R2313 B.n899 B.n421 32.0279
R2314 B.n905 B.n421 32.0279
R2315 B.n905 B.n417 32.0279
R2316 B.n911 B.n417 32.0279
R2317 B.n911 B.n413 32.0279
R2318 B.n917 B.n413 32.0279
R2319 B.n924 B.n409 32.0279
R2320 B.n924 B.n405 32.0279
R2321 B.n930 B.n405 32.0279
R2322 B.n930 B.n4 32.0279
R2323 B.n1070 B.n4 32.0279
R2324 B.n1070 B.n1069 32.0279
R2325 B.n1069 B.n1068 32.0279
R2326 B.n1068 B.n8 32.0279
R2327 B.n1062 B.n8 32.0279
R2328 B.n1062 B.n1061 32.0279
R2329 B.n1060 B.n15 32.0279
R2330 B.n1054 B.n15 32.0279
R2331 B.n1054 B.n1053 32.0279
R2332 B.n1053 B.n1052 32.0279
R2333 B.n1052 B.n22 32.0279
R2334 B.n1046 B.n22 32.0279
R2335 B.n1046 B.n1045 32.0279
R2336 B.n1044 B.n29 32.0279
R2337 B.n1038 B.n29 32.0279
R2338 B.n1038 B.n1037 32.0279
R2339 B.n1037 B.n1036 32.0279
R2340 B.n1036 B.n36 32.0279
R2341 B.n1030 B.n36 32.0279
R2342 B.n1030 B.n1029 32.0279
R2343 B.n1029 B.n1028 32.0279
R2344 B.n1022 B.n46 32.0279
R2345 B.n1022 B.n1021 32.0279
R2346 B.n1021 B.n1020 32.0279
R2347 B.n1020 B.n50 32.0279
R2348 B.n1014 B.n50 32.0279
R2349 B.n1014 B.n1013 32.0279
R2350 B.n1013 B.n1012 32.0279
R2351 B.n1012 B.n57 32.0279
R2352 B.n1006 B.n57 32.0279
R2353 B.n1006 B.n1005 32.0279
R2354 B.n1004 B.n64 32.0279
R2355 B.n998 B.n64 32.0279
R2356 B.n998 B.n997 32.0279
R2357 B.n997 B.n996 32.0279
R2358 B.n996 B.n71 32.0279
R2359 B.n990 B.n71 32.0279
R2360 B.n990 B.n989 32.0279
R2361 B.n862 B.t1 30.6149
R2362 B.n46 B.t0 30.6149
R2363 B.n148 B.n73 28.2542
R2364 B.n986 B.n985 28.2542
R2365 B.n811 B.n810 28.2542
R2366 B.n804 B.n478 28.2542
R2367 B.t2 B.n425 27.789
R2368 B.n1045 B.t4 27.789
R2369 B.t5 B.n409 22.1371
R2370 B.n1061 B.t3 22.1371
R2371 B.n832 B.t14 18.3692
R2372 B.t7 B.n1004 18.3692
R2373 B B.n1072 18.0485
R2374 B.t14 B.n464 13.6592
R2375 B.n1005 B.t7 13.6592
R2376 B.n149 B.n148 10.6151
R2377 B.n152 B.n149 10.6151
R2378 B.n153 B.n152 10.6151
R2379 B.n156 B.n153 10.6151
R2380 B.n157 B.n156 10.6151
R2381 B.n160 B.n157 10.6151
R2382 B.n161 B.n160 10.6151
R2383 B.n164 B.n161 10.6151
R2384 B.n165 B.n164 10.6151
R2385 B.n168 B.n165 10.6151
R2386 B.n169 B.n168 10.6151
R2387 B.n172 B.n169 10.6151
R2388 B.n173 B.n172 10.6151
R2389 B.n176 B.n173 10.6151
R2390 B.n177 B.n176 10.6151
R2391 B.n180 B.n177 10.6151
R2392 B.n181 B.n180 10.6151
R2393 B.n184 B.n181 10.6151
R2394 B.n185 B.n184 10.6151
R2395 B.n188 B.n185 10.6151
R2396 B.n189 B.n188 10.6151
R2397 B.n192 B.n189 10.6151
R2398 B.n193 B.n192 10.6151
R2399 B.n196 B.n193 10.6151
R2400 B.n197 B.n196 10.6151
R2401 B.n200 B.n197 10.6151
R2402 B.n201 B.n200 10.6151
R2403 B.n204 B.n201 10.6151
R2404 B.n205 B.n204 10.6151
R2405 B.n208 B.n205 10.6151
R2406 B.n209 B.n208 10.6151
R2407 B.n212 B.n209 10.6151
R2408 B.n213 B.n212 10.6151
R2409 B.n216 B.n213 10.6151
R2410 B.n217 B.n216 10.6151
R2411 B.n220 B.n217 10.6151
R2412 B.n221 B.n220 10.6151
R2413 B.n224 B.n221 10.6151
R2414 B.n225 B.n224 10.6151
R2415 B.n228 B.n225 10.6151
R2416 B.n229 B.n228 10.6151
R2417 B.n232 B.n229 10.6151
R2418 B.n233 B.n232 10.6151
R2419 B.n236 B.n233 10.6151
R2420 B.n237 B.n236 10.6151
R2421 B.n240 B.n237 10.6151
R2422 B.n241 B.n240 10.6151
R2423 B.n244 B.n241 10.6151
R2424 B.n245 B.n244 10.6151
R2425 B.n248 B.n245 10.6151
R2426 B.n249 B.n248 10.6151
R2427 B.n252 B.n249 10.6151
R2428 B.n253 B.n252 10.6151
R2429 B.n256 B.n253 10.6151
R2430 B.n257 B.n256 10.6151
R2431 B.n260 B.n257 10.6151
R2432 B.n261 B.n260 10.6151
R2433 B.n264 B.n261 10.6151
R2434 B.n265 B.n264 10.6151
R2435 B.n269 B.n268 10.6151
R2436 B.n272 B.n269 10.6151
R2437 B.n273 B.n272 10.6151
R2438 B.n276 B.n273 10.6151
R2439 B.n277 B.n276 10.6151
R2440 B.n280 B.n277 10.6151
R2441 B.n281 B.n280 10.6151
R2442 B.n284 B.n281 10.6151
R2443 B.n289 B.n286 10.6151
R2444 B.n290 B.n289 10.6151
R2445 B.n293 B.n290 10.6151
R2446 B.n294 B.n293 10.6151
R2447 B.n297 B.n294 10.6151
R2448 B.n298 B.n297 10.6151
R2449 B.n301 B.n298 10.6151
R2450 B.n302 B.n301 10.6151
R2451 B.n305 B.n302 10.6151
R2452 B.n306 B.n305 10.6151
R2453 B.n309 B.n306 10.6151
R2454 B.n310 B.n309 10.6151
R2455 B.n313 B.n310 10.6151
R2456 B.n314 B.n313 10.6151
R2457 B.n317 B.n314 10.6151
R2458 B.n318 B.n317 10.6151
R2459 B.n321 B.n318 10.6151
R2460 B.n322 B.n321 10.6151
R2461 B.n325 B.n322 10.6151
R2462 B.n326 B.n325 10.6151
R2463 B.n329 B.n326 10.6151
R2464 B.n330 B.n329 10.6151
R2465 B.n333 B.n330 10.6151
R2466 B.n334 B.n333 10.6151
R2467 B.n337 B.n334 10.6151
R2468 B.n338 B.n337 10.6151
R2469 B.n341 B.n338 10.6151
R2470 B.n342 B.n341 10.6151
R2471 B.n345 B.n342 10.6151
R2472 B.n346 B.n345 10.6151
R2473 B.n349 B.n346 10.6151
R2474 B.n350 B.n349 10.6151
R2475 B.n353 B.n350 10.6151
R2476 B.n354 B.n353 10.6151
R2477 B.n357 B.n354 10.6151
R2478 B.n358 B.n357 10.6151
R2479 B.n361 B.n358 10.6151
R2480 B.n362 B.n361 10.6151
R2481 B.n365 B.n362 10.6151
R2482 B.n366 B.n365 10.6151
R2483 B.n369 B.n366 10.6151
R2484 B.n370 B.n369 10.6151
R2485 B.n373 B.n370 10.6151
R2486 B.n374 B.n373 10.6151
R2487 B.n377 B.n374 10.6151
R2488 B.n378 B.n377 10.6151
R2489 B.n381 B.n378 10.6151
R2490 B.n382 B.n381 10.6151
R2491 B.n385 B.n382 10.6151
R2492 B.n386 B.n385 10.6151
R2493 B.n389 B.n386 10.6151
R2494 B.n390 B.n389 10.6151
R2495 B.n393 B.n390 10.6151
R2496 B.n394 B.n393 10.6151
R2497 B.n397 B.n394 10.6151
R2498 B.n398 B.n397 10.6151
R2499 B.n401 B.n398 10.6151
R2500 B.n402 B.n401 10.6151
R2501 B.n986 B.n402 10.6151
R2502 B.n812 B.n811 10.6151
R2503 B.n812 B.n474 10.6151
R2504 B.n822 B.n474 10.6151
R2505 B.n823 B.n822 10.6151
R2506 B.n824 B.n823 10.6151
R2507 B.n824 B.n466 10.6151
R2508 B.n834 B.n466 10.6151
R2509 B.n835 B.n834 10.6151
R2510 B.n836 B.n835 10.6151
R2511 B.n836 B.n458 10.6151
R2512 B.n846 B.n458 10.6151
R2513 B.n847 B.n846 10.6151
R2514 B.n848 B.n847 10.6151
R2515 B.n848 B.n450 10.6151
R2516 B.n858 B.n450 10.6151
R2517 B.n859 B.n858 10.6151
R2518 B.n860 B.n859 10.6151
R2519 B.n860 B.n443 10.6151
R2520 B.n871 B.n443 10.6151
R2521 B.n872 B.n871 10.6151
R2522 B.n873 B.n872 10.6151
R2523 B.n873 B.n435 10.6151
R2524 B.n883 B.n435 10.6151
R2525 B.n884 B.n883 10.6151
R2526 B.n885 B.n884 10.6151
R2527 B.n885 B.n427 10.6151
R2528 B.n895 B.n427 10.6151
R2529 B.n896 B.n895 10.6151
R2530 B.n897 B.n896 10.6151
R2531 B.n897 B.n419 10.6151
R2532 B.n907 B.n419 10.6151
R2533 B.n908 B.n907 10.6151
R2534 B.n909 B.n908 10.6151
R2535 B.n909 B.n411 10.6151
R2536 B.n919 B.n411 10.6151
R2537 B.n920 B.n919 10.6151
R2538 B.n922 B.n920 10.6151
R2539 B.n922 B.n921 10.6151
R2540 B.n921 B.n403 10.6151
R2541 B.n933 B.n403 10.6151
R2542 B.n934 B.n933 10.6151
R2543 B.n935 B.n934 10.6151
R2544 B.n936 B.n935 10.6151
R2545 B.n938 B.n936 10.6151
R2546 B.n939 B.n938 10.6151
R2547 B.n940 B.n939 10.6151
R2548 B.n941 B.n940 10.6151
R2549 B.n943 B.n941 10.6151
R2550 B.n944 B.n943 10.6151
R2551 B.n945 B.n944 10.6151
R2552 B.n946 B.n945 10.6151
R2553 B.n948 B.n946 10.6151
R2554 B.n949 B.n948 10.6151
R2555 B.n950 B.n949 10.6151
R2556 B.n951 B.n950 10.6151
R2557 B.n953 B.n951 10.6151
R2558 B.n954 B.n953 10.6151
R2559 B.n955 B.n954 10.6151
R2560 B.n956 B.n955 10.6151
R2561 B.n958 B.n956 10.6151
R2562 B.n959 B.n958 10.6151
R2563 B.n960 B.n959 10.6151
R2564 B.n961 B.n960 10.6151
R2565 B.n963 B.n961 10.6151
R2566 B.n964 B.n963 10.6151
R2567 B.n965 B.n964 10.6151
R2568 B.n966 B.n965 10.6151
R2569 B.n968 B.n966 10.6151
R2570 B.n969 B.n968 10.6151
R2571 B.n970 B.n969 10.6151
R2572 B.n971 B.n970 10.6151
R2573 B.n973 B.n971 10.6151
R2574 B.n974 B.n973 10.6151
R2575 B.n975 B.n974 10.6151
R2576 B.n976 B.n975 10.6151
R2577 B.n978 B.n976 10.6151
R2578 B.n979 B.n978 10.6151
R2579 B.n980 B.n979 10.6151
R2580 B.n981 B.n980 10.6151
R2581 B.n983 B.n981 10.6151
R2582 B.n984 B.n983 10.6151
R2583 B.n985 B.n984 10.6151
R2584 B.n804 B.n803 10.6151
R2585 B.n803 B.n802 10.6151
R2586 B.n802 B.n801 10.6151
R2587 B.n801 B.n799 10.6151
R2588 B.n799 B.n796 10.6151
R2589 B.n796 B.n795 10.6151
R2590 B.n795 B.n792 10.6151
R2591 B.n792 B.n791 10.6151
R2592 B.n791 B.n788 10.6151
R2593 B.n788 B.n787 10.6151
R2594 B.n787 B.n784 10.6151
R2595 B.n784 B.n783 10.6151
R2596 B.n783 B.n780 10.6151
R2597 B.n780 B.n779 10.6151
R2598 B.n779 B.n776 10.6151
R2599 B.n776 B.n775 10.6151
R2600 B.n775 B.n772 10.6151
R2601 B.n772 B.n771 10.6151
R2602 B.n771 B.n768 10.6151
R2603 B.n768 B.n767 10.6151
R2604 B.n767 B.n764 10.6151
R2605 B.n764 B.n763 10.6151
R2606 B.n763 B.n760 10.6151
R2607 B.n760 B.n759 10.6151
R2608 B.n759 B.n756 10.6151
R2609 B.n756 B.n755 10.6151
R2610 B.n755 B.n752 10.6151
R2611 B.n752 B.n751 10.6151
R2612 B.n751 B.n748 10.6151
R2613 B.n748 B.n747 10.6151
R2614 B.n747 B.n744 10.6151
R2615 B.n744 B.n743 10.6151
R2616 B.n743 B.n740 10.6151
R2617 B.n740 B.n739 10.6151
R2618 B.n739 B.n736 10.6151
R2619 B.n736 B.n735 10.6151
R2620 B.n735 B.n732 10.6151
R2621 B.n732 B.n731 10.6151
R2622 B.n731 B.n728 10.6151
R2623 B.n728 B.n727 10.6151
R2624 B.n727 B.n724 10.6151
R2625 B.n724 B.n723 10.6151
R2626 B.n723 B.n720 10.6151
R2627 B.n720 B.n719 10.6151
R2628 B.n719 B.n716 10.6151
R2629 B.n716 B.n715 10.6151
R2630 B.n715 B.n712 10.6151
R2631 B.n712 B.n711 10.6151
R2632 B.n711 B.n708 10.6151
R2633 B.n708 B.n707 10.6151
R2634 B.n707 B.n704 10.6151
R2635 B.n704 B.n703 10.6151
R2636 B.n703 B.n700 10.6151
R2637 B.n700 B.n699 10.6151
R2638 B.n699 B.n696 10.6151
R2639 B.n696 B.n695 10.6151
R2640 B.n695 B.n692 10.6151
R2641 B.n692 B.n691 10.6151
R2642 B.n691 B.n688 10.6151
R2643 B.n686 B.n683 10.6151
R2644 B.n683 B.n682 10.6151
R2645 B.n682 B.n679 10.6151
R2646 B.n679 B.n678 10.6151
R2647 B.n678 B.n675 10.6151
R2648 B.n675 B.n674 10.6151
R2649 B.n674 B.n671 10.6151
R2650 B.n671 B.n670 10.6151
R2651 B.n667 B.n666 10.6151
R2652 B.n666 B.n663 10.6151
R2653 B.n663 B.n662 10.6151
R2654 B.n662 B.n659 10.6151
R2655 B.n659 B.n658 10.6151
R2656 B.n658 B.n655 10.6151
R2657 B.n655 B.n654 10.6151
R2658 B.n654 B.n651 10.6151
R2659 B.n651 B.n650 10.6151
R2660 B.n650 B.n647 10.6151
R2661 B.n647 B.n646 10.6151
R2662 B.n646 B.n643 10.6151
R2663 B.n643 B.n642 10.6151
R2664 B.n642 B.n639 10.6151
R2665 B.n639 B.n638 10.6151
R2666 B.n638 B.n635 10.6151
R2667 B.n635 B.n634 10.6151
R2668 B.n634 B.n631 10.6151
R2669 B.n631 B.n630 10.6151
R2670 B.n630 B.n627 10.6151
R2671 B.n627 B.n626 10.6151
R2672 B.n626 B.n623 10.6151
R2673 B.n623 B.n622 10.6151
R2674 B.n622 B.n619 10.6151
R2675 B.n619 B.n618 10.6151
R2676 B.n618 B.n615 10.6151
R2677 B.n615 B.n614 10.6151
R2678 B.n614 B.n611 10.6151
R2679 B.n611 B.n610 10.6151
R2680 B.n610 B.n607 10.6151
R2681 B.n607 B.n606 10.6151
R2682 B.n606 B.n603 10.6151
R2683 B.n603 B.n602 10.6151
R2684 B.n602 B.n599 10.6151
R2685 B.n599 B.n598 10.6151
R2686 B.n598 B.n595 10.6151
R2687 B.n595 B.n594 10.6151
R2688 B.n594 B.n591 10.6151
R2689 B.n591 B.n590 10.6151
R2690 B.n590 B.n587 10.6151
R2691 B.n587 B.n586 10.6151
R2692 B.n586 B.n583 10.6151
R2693 B.n583 B.n582 10.6151
R2694 B.n582 B.n579 10.6151
R2695 B.n579 B.n578 10.6151
R2696 B.n578 B.n575 10.6151
R2697 B.n575 B.n574 10.6151
R2698 B.n574 B.n571 10.6151
R2699 B.n571 B.n570 10.6151
R2700 B.n570 B.n567 10.6151
R2701 B.n567 B.n566 10.6151
R2702 B.n566 B.n563 10.6151
R2703 B.n563 B.n562 10.6151
R2704 B.n562 B.n559 10.6151
R2705 B.n559 B.n558 10.6151
R2706 B.n558 B.n555 10.6151
R2707 B.n555 B.n554 10.6151
R2708 B.n554 B.n482 10.6151
R2709 B.n810 B.n482 10.6151
R2710 B.n816 B.n478 10.6151
R2711 B.n817 B.n816 10.6151
R2712 B.n818 B.n817 10.6151
R2713 B.n818 B.n470 10.6151
R2714 B.n828 B.n470 10.6151
R2715 B.n829 B.n828 10.6151
R2716 B.n830 B.n829 10.6151
R2717 B.n830 B.n462 10.6151
R2718 B.n840 B.n462 10.6151
R2719 B.n841 B.n840 10.6151
R2720 B.n842 B.n841 10.6151
R2721 B.n842 B.n454 10.6151
R2722 B.n852 B.n454 10.6151
R2723 B.n853 B.n852 10.6151
R2724 B.n854 B.n853 10.6151
R2725 B.n854 B.n446 10.6151
R2726 B.n865 B.n446 10.6151
R2727 B.n866 B.n865 10.6151
R2728 B.n867 B.n866 10.6151
R2729 B.n867 B.n439 10.6151
R2730 B.n877 B.n439 10.6151
R2731 B.n878 B.n877 10.6151
R2732 B.n879 B.n878 10.6151
R2733 B.n879 B.n431 10.6151
R2734 B.n889 B.n431 10.6151
R2735 B.n890 B.n889 10.6151
R2736 B.n891 B.n890 10.6151
R2737 B.n891 B.n423 10.6151
R2738 B.n901 B.n423 10.6151
R2739 B.n902 B.n901 10.6151
R2740 B.n903 B.n902 10.6151
R2741 B.n903 B.n415 10.6151
R2742 B.n913 B.n415 10.6151
R2743 B.n914 B.n913 10.6151
R2744 B.n915 B.n914 10.6151
R2745 B.n915 B.n407 10.6151
R2746 B.n926 B.n407 10.6151
R2747 B.n927 B.n926 10.6151
R2748 B.n928 B.n927 10.6151
R2749 B.n928 B.n0 10.6151
R2750 B.n1066 B.n1 10.6151
R2751 B.n1066 B.n1065 10.6151
R2752 B.n1065 B.n1064 10.6151
R2753 B.n1064 B.n10 10.6151
R2754 B.n1058 B.n10 10.6151
R2755 B.n1058 B.n1057 10.6151
R2756 B.n1057 B.n1056 10.6151
R2757 B.n1056 B.n17 10.6151
R2758 B.n1050 B.n17 10.6151
R2759 B.n1050 B.n1049 10.6151
R2760 B.n1049 B.n1048 10.6151
R2761 B.n1048 B.n24 10.6151
R2762 B.n1042 B.n24 10.6151
R2763 B.n1042 B.n1041 10.6151
R2764 B.n1041 B.n1040 10.6151
R2765 B.n1040 B.n31 10.6151
R2766 B.n1034 B.n31 10.6151
R2767 B.n1034 B.n1033 10.6151
R2768 B.n1033 B.n1032 10.6151
R2769 B.n1032 B.n38 10.6151
R2770 B.n1026 B.n38 10.6151
R2771 B.n1026 B.n1025 10.6151
R2772 B.n1025 B.n1024 10.6151
R2773 B.n1024 B.n44 10.6151
R2774 B.n1018 B.n44 10.6151
R2775 B.n1018 B.n1017 10.6151
R2776 B.n1017 B.n1016 10.6151
R2777 B.n1016 B.n52 10.6151
R2778 B.n1010 B.n52 10.6151
R2779 B.n1010 B.n1009 10.6151
R2780 B.n1009 B.n1008 10.6151
R2781 B.n1008 B.n59 10.6151
R2782 B.n1002 B.n59 10.6151
R2783 B.n1002 B.n1001 10.6151
R2784 B.n1001 B.n1000 10.6151
R2785 B.n1000 B.n66 10.6151
R2786 B.n994 B.n66 10.6151
R2787 B.n994 B.n993 10.6151
R2788 B.n993 B.n992 10.6151
R2789 B.n992 B.n73 10.6151
R2790 B.n917 B.t5 9.89132
R2791 B.t3 B.n1060 9.89132
R2792 B.n268 B.n146 6.5566
R2793 B.n285 B.n284 6.5566
R2794 B.n687 B.n686 6.5566
R2795 B.n670 B.n552 6.5566
R2796 B.n893 B.t2 4.23942
R2797 B.t4 B.n1044 4.23942
R2798 B.n265 B.n146 4.05904
R2799 B.n286 B.n285 4.05904
R2800 B.n688 B.n687 4.05904
R2801 B.n667 B.n552 4.05904
R2802 B.n1072 B.n0 2.81026
R2803 B.n1072 B.n1 2.81026
R2804 B.n869 B.t1 1.41347
R2805 B.n1028 B.t0 1.41347
R2806 VN.n3 VN.t0 212.732
R2807 VN.n17 VN.t3 212.732
R2808 VN.n4 VN.t4 177.849
R2809 VN.n12 VN.t1 177.849
R2810 VN.n18 VN.t5 177.849
R2811 VN.n26 VN.t2 177.849
R2812 VN.n25 VN.n14 161.3
R2813 VN.n24 VN.n23 161.3
R2814 VN.n22 VN.n15 161.3
R2815 VN.n21 VN.n20 161.3
R2816 VN.n19 VN.n16 161.3
R2817 VN.n11 VN.n0 161.3
R2818 VN.n10 VN.n9 161.3
R2819 VN.n8 VN.n1 161.3
R2820 VN.n7 VN.n6 161.3
R2821 VN.n5 VN.n2 161.3
R2822 VN.n13 VN.n12 97.1368
R2823 VN.n27 VN.n26 97.1368
R2824 VN VN.n27 53.0133
R2825 VN.n6 VN.n1 51.2335
R2826 VN.n20 VN.n15 51.2335
R2827 VN.n4 VN.n3 48.154
R2828 VN.n18 VN.n17 48.154
R2829 VN.n10 VN.n1 29.9206
R2830 VN.n24 VN.n15 29.9206
R2831 VN.n5 VN.n4 24.5923
R2832 VN.n6 VN.n5 24.5923
R2833 VN.n11 VN.n10 24.5923
R2834 VN.n20 VN.n19 24.5923
R2835 VN.n19 VN.n18 24.5923
R2836 VN.n25 VN.n24 24.5923
R2837 VN.n12 VN.n11 13.7719
R2838 VN.n26 VN.n25 13.7719
R2839 VN.n17 VN.n16 6.57284
R2840 VN.n3 VN.n2 6.57284
R2841 VN.n27 VN.n14 0.278335
R2842 VN.n13 VN.n0 0.278335
R2843 VN.n23 VN.n14 0.189894
R2844 VN.n23 VN.n22 0.189894
R2845 VN.n22 VN.n21 0.189894
R2846 VN.n21 VN.n16 0.189894
R2847 VN.n7 VN.n2 0.189894
R2848 VN.n8 VN.n7 0.189894
R2849 VN.n9 VN.n8 0.189894
R2850 VN.n9 VN.n0 0.189894
R2851 VN VN.n13 0.153485
R2852 VDD2.n199 VDD2.n198 289.615
R2853 VDD2.n98 VDD2.n97 289.615
R2854 VDD2.n198 VDD2.n197 185
R2855 VDD2.n103 VDD2.n102 185
R2856 VDD2.n192 VDD2.n191 185
R2857 VDD2.n190 VDD2.n189 185
R2858 VDD2.n107 VDD2.n106 185
R2859 VDD2.n184 VDD2.n183 185
R2860 VDD2.n182 VDD2.n181 185
R2861 VDD2.n111 VDD2.n110 185
R2862 VDD2.n176 VDD2.n175 185
R2863 VDD2.n174 VDD2.n173 185
R2864 VDD2.n115 VDD2.n114 185
R2865 VDD2.n168 VDD2.n167 185
R2866 VDD2.n166 VDD2.n165 185
R2867 VDD2.n119 VDD2.n118 185
R2868 VDD2.n160 VDD2.n159 185
R2869 VDD2.n158 VDD2.n157 185
R2870 VDD2.n156 VDD2.n122 185
R2871 VDD2.n126 VDD2.n123 185
R2872 VDD2.n151 VDD2.n150 185
R2873 VDD2.n149 VDD2.n148 185
R2874 VDD2.n128 VDD2.n127 185
R2875 VDD2.n143 VDD2.n142 185
R2876 VDD2.n141 VDD2.n140 185
R2877 VDD2.n132 VDD2.n131 185
R2878 VDD2.n135 VDD2.n134 185
R2879 VDD2.n33 VDD2.n32 185
R2880 VDD2.n30 VDD2.n29 185
R2881 VDD2.n39 VDD2.n38 185
R2882 VDD2.n41 VDD2.n40 185
R2883 VDD2.n26 VDD2.n25 185
R2884 VDD2.n47 VDD2.n46 185
R2885 VDD2.n50 VDD2.n49 185
R2886 VDD2.n48 VDD2.n22 185
R2887 VDD2.n55 VDD2.n21 185
R2888 VDD2.n57 VDD2.n56 185
R2889 VDD2.n59 VDD2.n58 185
R2890 VDD2.n18 VDD2.n17 185
R2891 VDD2.n65 VDD2.n64 185
R2892 VDD2.n67 VDD2.n66 185
R2893 VDD2.n14 VDD2.n13 185
R2894 VDD2.n73 VDD2.n72 185
R2895 VDD2.n75 VDD2.n74 185
R2896 VDD2.n10 VDD2.n9 185
R2897 VDD2.n81 VDD2.n80 185
R2898 VDD2.n83 VDD2.n82 185
R2899 VDD2.n6 VDD2.n5 185
R2900 VDD2.n89 VDD2.n88 185
R2901 VDD2.n91 VDD2.n90 185
R2902 VDD2.n2 VDD2.n1 185
R2903 VDD2.n97 VDD2.n96 185
R2904 VDD2.t3 VDD2.n133 149.524
R2905 VDD2.t5 VDD2.n31 149.524
R2906 VDD2.n198 VDD2.n102 104.615
R2907 VDD2.n191 VDD2.n102 104.615
R2908 VDD2.n191 VDD2.n190 104.615
R2909 VDD2.n190 VDD2.n106 104.615
R2910 VDD2.n183 VDD2.n106 104.615
R2911 VDD2.n183 VDD2.n182 104.615
R2912 VDD2.n182 VDD2.n110 104.615
R2913 VDD2.n175 VDD2.n110 104.615
R2914 VDD2.n175 VDD2.n174 104.615
R2915 VDD2.n174 VDD2.n114 104.615
R2916 VDD2.n167 VDD2.n114 104.615
R2917 VDD2.n167 VDD2.n166 104.615
R2918 VDD2.n166 VDD2.n118 104.615
R2919 VDD2.n159 VDD2.n118 104.615
R2920 VDD2.n159 VDD2.n158 104.615
R2921 VDD2.n158 VDD2.n122 104.615
R2922 VDD2.n126 VDD2.n122 104.615
R2923 VDD2.n150 VDD2.n126 104.615
R2924 VDD2.n150 VDD2.n149 104.615
R2925 VDD2.n149 VDD2.n127 104.615
R2926 VDD2.n142 VDD2.n127 104.615
R2927 VDD2.n142 VDD2.n141 104.615
R2928 VDD2.n141 VDD2.n131 104.615
R2929 VDD2.n134 VDD2.n131 104.615
R2930 VDD2.n32 VDD2.n29 104.615
R2931 VDD2.n39 VDD2.n29 104.615
R2932 VDD2.n40 VDD2.n39 104.615
R2933 VDD2.n40 VDD2.n25 104.615
R2934 VDD2.n47 VDD2.n25 104.615
R2935 VDD2.n49 VDD2.n47 104.615
R2936 VDD2.n49 VDD2.n48 104.615
R2937 VDD2.n48 VDD2.n21 104.615
R2938 VDD2.n57 VDD2.n21 104.615
R2939 VDD2.n58 VDD2.n57 104.615
R2940 VDD2.n58 VDD2.n17 104.615
R2941 VDD2.n65 VDD2.n17 104.615
R2942 VDD2.n66 VDD2.n65 104.615
R2943 VDD2.n66 VDD2.n13 104.615
R2944 VDD2.n73 VDD2.n13 104.615
R2945 VDD2.n74 VDD2.n73 104.615
R2946 VDD2.n74 VDD2.n9 104.615
R2947 VDD2.n81 VDD2.n9 104.615
R2948 VDD2.n82 VDD2.n81 104.615
R2949 VDD2.n82 VDD2.n5 104.615
R2950 VDD2.n89 VDD2.n5 104.615
R2951 VDD2.n90 VDD2.n89 104.615
R2952 VDD2.n90 VDD2.n1 104.615
R2953 VDD2.n97 VDD2.n1 104.615
R2954 VDD2.n100 VDD2.n99 64.5293
R2955 VDD2 VDD2.n201 64.5255
R2956 VDD2.n100 VDD2.n98 53.3214
R2957 VDD2.n134 VDD2.t3 52.3082
R2958 VDD2.n32 VDD2.t5 52.3082
R2959 VDD2.n200 VDD2.n199 51.5793
R2960 VDD2.n200 VDD2.n100 47.0903
R2961 VDD2.n157 VDD2.n156 13.1884
R2962 VDD2.n56 VDD2.n55 13.1884
R2963 VDD2.n160 VDD2.n121 12.8005
R2964 VDD2.n155 VDD2.n123 12.8005
R2965 VDD2.n54 VDD2.n22 12.8005
R2966 VDD2.n59 VDD2.n20 12.8005
R2967 VDD2.n197 VDD2.n101 12.0247
R2968 VDD2.n161 VDD2.n119 12.0247
R2969 VDD2.n152 VDD2.n151 12.0247
R2970 VDD2.n51 VDD2.n50 12.0247
R2971 VDD2.n60 VDD2.n18 12.0247
R2972 VDD2.n96 VDD2.n0 12.0247
R2973 VDD2.n196 VDD2.n103 11.249
R2974 VDD2.n165 VDD2.n164 11.249
R2975 VDD2.n148 VDD2.n125 11.249
R2976 VDD2.n46 VDD2.n24 11.249
R2977 VDD2.n64 VDD2.n63 11.249
R2978 VDD2.n95 VDD2.n2 11.249
R2979 VDD2.n193 VDD2.n192 10.4732
R2980 VDD2.n168 VDD2.n117 10.4732
R2981 VDD2.n147 VDD2.n128 10.4732
R2982 VDD2.n45 VDD2.n26 10.4732
R2983 VDD2.n67 VDD2.n16 10.4732
R2984 VDD2.n92 VDD2.n91 10.4732
R2985 VDD2.n135 VDD2.n133 10.2747
R2986 VDD2.n33 VDD2.n31 10.2747
R2987 VDD2.n189 VDD2.n105 9.69747
R2988 VDD2.n169 VDD2.n115 9.69747
R2989 VDD2.n144 VDD2.n143 9.69747
R2990 VDD2.n42 VDD2.n41 9.69747
R2991 VDD2.n68 VDD2.n14 9.69747
R2992 VDD2.n88 VDD2.n4 9.69747
R2993 VDD2.n195 VDD2.n101 9.45567
R2994 VDD2.n94 VDD2.n0 9.45567
R2995 VDD2.n137 VDD2.n136 9.3005
R2996 VDD2.n139 VDD2.n138 9.3005
R2997 VDD2.n130 VDD2.n129 9.3005
R2998 VDD2.n145 VDD2.n144 9.3005
R2999 VDD2.n147 VDD2.n146 9.3005
R3000 VDD2.n125 VDD2.n124 9.3005
R3001 VDD2.n153 VDD2.n152 9.3005
R3002 VDD2.n155 VDD2.n154 9.3005
R3003 VDD2.n109 VDD2.n108 9.3005
R3004 VDD2.n186 VDD2.n185 9.3005
R3005 VDD2.n188 VDD2.n187 9.3005
R3006 VDD2.n105 VDD2.n104 9.3005
R3007 VDD2.n194 VDD2.n193 9.3005
R3008 VDD2.n196 VDD2.n195 9.3005
R3009 VDD2.n180 VDD2.n179 9.3005
R3010 VDD2.n178 VDD2.n177 9.3005
R3011 VDD2.n113 VDD2.n112 9.3005
R3012 VDD2.n172 VDD2.n171 9.3005
R3013 VDD2.n170 VDD2.n169 9.3005
R3014 VDD2.n117 VDD2.n116 9.3005
R3015 VDD2.n164 VDD2.n163 9.3005
R3016 VDD2.n162 VDD2.n161 9.3005
R3017 VDD2.n121 VDD2.n120 9.3005
R3018 VDD2.n79 VDD2.n78 9.3005
R3019 VDD2.n8 VDD2.n7 9.3005
R3020 VDD2.n85 VDD2.n84 9.3005
R3021 VDD2.n87 VDD2.n86 9.3005
R3022 VDD2.n4 VDD2.n3 9.3005
R3023 VDD2.n93 VDD2.n92 9.3005
R3024 VDD2.n95 VDD2.n94 9.3005
R3025 VDD2.n12 VDD2.n11 9.3005
R3026 VDD2.n71 VDD2.n70 9.3005
R3027 VDD2.n69 VDD2.n68 9.3005
R3028 VDD2.n16 VDD2.n15 9.3005
R3029 VDD2.n63 VDD2.n62 9.3005
R3030 VDD2.n61 VDD2.n60 9.3005
R3031 VDD2.n20 VDD2.n19 9.3005
R3032 VDD2.n35 VDD2.n34 9.3005
R3033 VDD2.n37 VDD2.n36 9.3005
R3034 VDD2.n28 VDD2.n27 9.3005
R3035 VDD2.n43 VDD2.n42 9.3005
R3036 VDD2.n45 VDD2.n44 9.3005
R3037 VDD2.n24 VDD2.n23 9.3005
R3038 VDD2.n52 VDD2.n51 9.3005
R3039 VDD2.n54 VDD2.n53 9.3005
R3040 VDD2.n77 VDD2.n76 9.3005
R3041 VDD2.n188 VDD2.n107 8.92171
R3042 VDD2.n173 VDD2.n172 8.92171
R3043 VDD2.n140 VDD2.n130 8.92171
R3044 VDD2.n38 VDD2.n28 8.92171
R3045 VDD2.n72 VDD2.n71 8.92171
R3046 VDD2.n87 VDD2.n6 8.92171
R3047 VDD2.n185 VDD2.n184 8.14595
R3048 VDD2.n176 VDD2.n113 8.14595
R3049 VDD2.n139 VDD2.n132 8.14595
R3050 VDD2.n37 VDD2.n30 8.14595
R3051 VDD2.n75 VDD2.n12 8.14595
R3052 VDD2.n84 VDD2.n83 8.14595
R3053 VDD2.n181 VDD2.n109 7.3702
R3054 VDD2.n177 VDD2.n111 7.3702
R3055 VDD2.n136 VDD2.n135 7.3702
R3056 VDD2.n34 VDD2.n33 7.3702
R3057 VDD2.n76 VDD2.n10 7.3702
R3058 VDD2.n80 VDD2.n8 7.3702
R3059 VDD2.n181 VDD2.n180 6.59444
R3060 VDD2.n180 VDD2.n111 6.59444
R3061 VDD2.n79 VDD2.n10 6.59444
R3062 VDD2.n80 VDD2.n79 6.59444
R3063 VDD2.n184 VDD2.n109 5.81868
R3064 VDD2.n177 VDD2.n176 5.81868
R3065 VDD2.n136 VDD2.n132 5.81868
R3066 VDD2.n34 VDD2.n30 5.81868
R3067 VDD2.n76 VDD2.n75 5.81868
R3068 VDD2.n83 VDD2.n8 5.81868
R3069 VDD2.n185 VDD2.n107 5.04292
R3070 VDD2.n173 VDD2.n113 5.04292
R3071 VDD2.n140 VDD2.n139 5.04292
R3072 VDD2.n38 VDD2.n37 5.04292
R3073 VDD2.n72 VDD2.n12 5.04292
R3074 VDD2.n84 VDD2.n6 5.04292
R3075 VDD2.n189 VDD2.n188 4.26717
R3076 VDD2.n172 VDD2.n115 4.26717
R3077 VDD2.n143 VDD2.n130 4.26717
R3078 VDD2.n41 VDD2.n28 4.26717
R3079 VDD2.n71 VDD2.n14 4.26717
R3080 VDD2.n88 VDD2.n87 4.26717
R3081 VDD2.n192 VDD2.n105 3.49141
R3082 VDD2.n169 VDD2.n168 3.49141
R3083 VDD2.n144 VDD2.n128 3.49141
R3084 VDD2.n42 VDD2.n26 3.49141
R3085 VDD2.n68 VDD2.n67 3.49141
R3086 VDD2.n91 VDD2.n4 3.49141
R3087 VDD2.n137 VDD2.n133 2.84303
R3088 VDD2.n35 VDD2.n31 2.84303
R3089 VDD2.n193 VDD2.n103 2.71565
R3090 VDD2.n165 VDD2.n117 2.71565
R3091 VDD2.n148 VDD2.n147 2.71565
R3092 VDD2.n46 VDD2.n45 2.71565
R3093 VDD2.n64 VDD2.n16 2.71565
R3094 VDD2.n92 VDD2.n2 2.71565
R3095 VDD2.n197 VDD2.n196 1.93989
R3096 VDD2.n164 VDD2.n119 1.93989
R3097 VDD2.n151 VDD2.n125 1.93989
R3098 VDD2.n50 VDD2.n24 1.93989
R3099 VDD2.n63 VDD2.n18 1.93989
R3100 VDD2.n96 VDD2.n95 1.93989
R3101 VDD2 VDD2.n200 1.8561
R3102 VDD2.n199 VDD2.n101 1.16414
R3103 VDD2.n161 VDD2.n160 1.16414
R3104 VDD2.n152 VDD2.n123 1.16414
R3105 VDD2.n51 VDD2.n22 1.16414
R3106 VDD2.n60 VDD2.n59 1.16414
R3107 VDD2.n98 VDD2.n0 1.16414
R3108 VDD2.n201 VDD2.t0 1.09563
R3109 VDD2.n201 VDD2.t2 1.09563
R3110 VDD2.n99 VDD2.t1 1.09563
R3111 VDD2.n99 VDD2.t4 1.09563
R3112 VDD2.n157 VDD2.n121 0.388379
R3113 VDD2.n156 VDD2.n155 0.388379
R3114 VDD2.n55 VDD2.n54 0.388379
R3115 VDD2.n56 VDD2.n20 0.388379
R3116 VDD2.n195 VDD2.n194 0.155672
R3117 VDD2.n194 VDD2.n104 0.155672
R3118 VDD2.n187 VDD2.n104 0.155672
R3119 VDD2.n187 VDD2.n186 0.155672
R3120 VDD2.n186 VDD2.n108 0.155672
R3121 VDD2.n179 VDD2.n108 0.155672
R3122 VDD2.n179 VDD2.n178 0.155672
R3123 VDD2.n178 VDD2.n112 0.155672
R3124 VDD2.n171 VDD2.n112 0.155672
R3125 VDD2.n171 VDD2.n170 0.155672
R3126 VDD2.n170 VDD2.n116 0.155672
R3127 VDD2.n163 VDD2.n116 0.155672
R3128 VDD2.n163 VDD2.n162 0.155672
R3129 VDD2.n162 VDD2.n120 0.155672
R3130 VDD2.n154 VDD2.n120 0.155672
R3131 VDD2.n154 VDD2.n153 0.155672
R3132 VDD2.n153 VDD2.n124 0.155672
R3133 VDD2.n146 VDD2.n124 0.155672
R3134 VDD2.n146 VDD2.n145 0.155672
R3135 VDD2.n145 VDD2.n129 0.155672
R3136 VDD2.n138 VDD2.n129 0.155672
R3137 VDD2.n138 VDD2.n137 0.155672
R3138 VDD2.n36 VDD2.n35 0.155672
R3139 VDD2.n36 VDD2.n27 0.155672
R3140 VDD2.n43 VDD2.n27 0.155672
R3141 VDD2.n44 VDD2.n43 0.155672
R3142 VDD2.n44 VDD2.n23 0.155672
R3143 VDD2.n52 VDD2.n23 0.155672
R3144 VDD2.n53 VDD2.n52 0.155672
R3145 VDD2.n53 VDD2.n19 0.155672
R3146 VDD2.n61 VDD2.n19 0.155672
R3147 VDD2.n62 VDD2.n61 0.155672
R3148 VDD2.n62 VDD2.n15 0.155672
R3149 VDD2.n69 VDD2.n15 0.155672
R3150 VDD2.n70 VDD2.n69 0.155672
R3151 VDD2.n70 VDD2.n11 0.155672
R3152 VDD2.n77 VDD2.n11 0.155672
R3153 VDD2.n78 VDD2.n77 0.155672
R3154 VDD2.n78 VDD2.n7 0.155672
R3155 VDD2.n85 VDD2.n7 0.155672
R3156 VDD2.n86 VDD2.n85 0.155672
R3157 VDD2.n86 VDD2.n3 0.155672
R3158 VDD2.n93 VDD2.n3 0.155672
R3159 VDD2.n94 VDD2.n93 0.155672
C0 VDD1 VDD2 1.34914f
C1 VN VTAIL 9.67654f
C2 VN VP 7.90076f
C3 VTAIL VP 9.69094f
C4 VDD1 VN 0.150841f
C5 VDD1 VTAIL 9.96515f
C6 VDD2 VN 9.82271f
C7 VDD2 VTAIL 10.0133f
C8 VDD1 VP 10.1139f
C9 VDD2 VP 0.446423f
C10 VDD2 B 6.947706f
C11 VDD1 B 7.077899f
C12 VTAIL B 10.137278f
C13 VN B 12.97726f
C14 VP B 11.462892f
C15 VDD2.n0 B 0.011941f
C16 VDD2.n1 B 0.0269f
C17 VDD2.n2 B 0.01205f
C18 VDD2.n3 B 0.021179f
C19 VDD2.n4 B 0.011381f
C20 VDD2.n5 B 0.0269f
C21 VDD2.n6 B 0.01205f
C22 VDD2.n7 B 0.021179f
C23 VDD2.n8 B 0.011381f
C24 VDD2.n9 B 0.0269f
C25 VDD2.n10 B 0.01205f
C26 VDD2.n11 B 0.021179f
C27 VDD2.n12 B 0.011381f
C28 VDD2.n13 B 0.0269f
C29 VDD2.n14 B 0.01205f
C30 VDD2.n15 B 0.021179f
C31 VDD2.n16 B 0.011381f
C32 VDD2.n17 B 0.0269f
C33 VDD2.n18 B 0.01205f
C34 VDD2.n19 B 0.021179f
C35 VDD2.n20 B 0.011381f
C36 VDD2.n21 B 0.0269f
C37 VDD2.n22 B 0.01205f
C38 VDD2.n23 B 0.021179f
C39 VDD2.n24 B 0.011381f
C40 VDD2.n25 B 0.0269f
C41 VDD2.n26 B 0.01205f
C42 VDD2.n27 B 0.021179f
C43 VDD2.n28 B 0.011381f
C44 VDD2.n29 B 0.0269f
C45 VDD2.n30 B 0.01205f
C46 VDD2.n31 B 0.202133f
C47 VDD2.t5 B 0.046125f
C48 VDD2.n32 B 0.020175f
C49 VDD2.n33 B 0.019016f
C50 VDD2.n34 B 0.011381f
C51 VDD2.n35 B 1.64117f
C52 VDD2.n36 B 0.021179f
C53 VDD2.n37 B 0.011381f
C54 VDD2.n38 B 0.01205f
C55 VDD2.n39 B 0.0269f
C56 VDD2.n40 B 0.0269f
C57 VDD2.n41 B 0.01205f
C58 VDD2.n42 B 0.011381f
C59 VDD2.n43 B 0.021179f
C60 VDD2.n44 B 0.021179f
C61 VDD2.n45 B 0.011381f
C62 VDD2.n46 B 0.01205f
C63 VDD2.n47 B 0.0269f
C64 VDD2.n48 B 0.0269f
C65 VDD2.n49 B 0.0269f
C66 VDD2.n50 B 0.01205f
C67 VDD2.n51 B 0.011381f
C68 VDD2.n52 B 0.021179f
C69 VDD2.n53 B 0.021179f
C70 VDD2.n54 B 0.011381f
C71 VDD2.n55 B 0.011715f
C72 VDD2.n56 B 0.011715f
C73 VDD2.n57 B 0.0269f
C74 VDD2.n58 B 0.0269f
C75 VDD2.n59 B 0.01205f
C76 VDD2.n60 B 0.011381f
C77 VDD2.n61 B 0.021179f
C78 VDD2.n62 B 0.021179f
C79 VDD2.n63 B 0.011381f
C80 VDD2.n64 B 0.01205f
C81 VDD2.n65 B 0.0269f
C82 VDD2.n66 B 0.0269f
C83 VDD2.n67 B 0.01205f
C84 VDD2.n68 B 0.011381f
C85 VDD2.n69 B 0.021179f
C86 VDD2.n70 B 0.021179f
C87 VDD2.n71 B 0.011381f
C88 VDD2.n72 B 0.01205f
C89 VDD2.n73 B 0.0269f
C90 VDD2.n74 B 0.0269f
C91 VDD2.n75 B 0.01205f
C92 VDD2.n76 B 0.011381f
C93 VDD2.n77 B 0.021179f
C94 VDD2.n78 B 0.021179f
C95 VDD2.n79 B 0.011381f
C96 VDD2.n80 B 0.01205f
C97 VDD2.n81 B 0.0269f
C98 VDD2.n82 B 0.0269f
C99 VDD2.n83 B 0.01205f
C100 VDD2.n84 B 0.011381f
C101 VDD2.n85 B 0.021179f
C102 VDD2.n86 B 0.021179f
C103 VDD2.n87 B 0.011381f
C104 VDD2.n88 B 0.01205f
C105 VDD2.n89 B 0.0269f
C106 VDD2.n90 B 0.0269f
C107 VDD2.n91 B 0.01205f
C108 VDD2.n92 B 0.011381f
C109 VDD2.n93 B 0.021179f
C110 VDD2.n94 B 0.05474f
C111 VDD2.n95 B 0.011381f
C112 VDD2.n96 B 0.01205f
C113 VDD2.n97 B 0.05419f
C114 VDD2.n98 B 0.065827f
C115 VDD2.t1 B 0.30259f
C116 VDD2.t4 B 0.30259f
C117 VDD2.n99 B 2.76871f
C118 VDD2.n100 B 2.53131f
C119 VDD2.n101 B 0.011941f
C120 VDD2.n102 B 0.0269f
C121 VDD2.n103 B 0.01205f
C122 VDD2.n104 B 0.021179f
C123 VDD2.n105 B 0.011381f
C124 VDD2.n106 B 0.0269f
C125 VDD2.n107 B 0.01205f
C126 VDD2.n108 B 0.021179f
C127 VDD2.n109 B 0.011381f
C128 VDD2.n110 B 0.0269f
C129 VDD2.n111 B 0.01205f
C130 VDD2.n112 B 0.021179f
C131 VDD2.n113 B 0.011381f
C132 VDD2.n114 B 0.0269f
C133 VDD2.n115 B 0.01205f
C134 VDD2.n116 B 0.021179f
C135 VDD2.n117 B 0.011381f
C136 VDD2.n118 B 0.0269f
C137 VDD2.n119 B 0.01205f
C138 VDD2.n120 B 0.021179f
C139 VDD2.n121 B 0.011381f
C140 VDD2.n122 B 0.0269f
C141 VDD2.n123 B 0.01205f
C142 VDD2.n124 B 0.021179f
C143 VDD2.n125 B 0.011381f
C144 VDD2.n126 B 0.0269f
C145 VDD2.n127 B 0.0269f
C146 VDD2.n128 B 0.01205f
C147 VDD2.n129 B 0.021179f
C148 VDD2.n130 B 0.011381f
C149 VDD2.n131 B 0.0269f
C150 VDD2.n132 B 0.01205f
C151 VDD2.n133 B 0.202133f
C152 VDD2.t3 B 0.046125f
C153 VDD2.n134 B 0.020175f
C154 VDD2.n135 B 0.019016f
C155 VDD2.n136 B 0.011381f
C156 VDD2.n137 B 1.64117f
C157 VDD2.n138 B 0.021179f
C158 VDD2.n139 B 0.011381f
C159 VDD2.n140 B 0.01205f
C160 VDD2.n141 B 0.0269f
C161 VDD2.n142 B 0.0269f
C162 VDD2.n143 B 0.01205f
C163 VDD2.n144 B 0.011381f
C164 VDD2.n145 B 0.021179f
C165 VDD2.n146 B 0.021179f
C166 VDD2.n147 B 0.011381f
C167 VDD2.n148 B 0.01205f
C168 VDD2.n149 B 0.0269f
C169 VDD2.n150 B 0.0269f
C170 VDD2.n151 B 0.01205f
C171 VDD2.n152 B 0.011381f
C172 VDD2.n153 B 0.021179f
C173 VDD2.n154 B 0.021179f
C174 VDD2.n155 B 0.011381f
C175 VDD2.n156 B 0.011715f
C176 VDD2.n157 B 0.011715f
C177 VDD2.n158 B 0.0269f
C178 VDD2.n159 B 0.0269f
C179 VDD2.n160 B 0.01205f
C180 VDD2.n161 B 0.011381f
C181 VDD2.n162 B 0.021179f
C182 VDD2.n163 B 0.021179f
C183 VDD2.n164 B 0.011381f
C184 VDD2.n165 B 0.01205f
C185 VDD2.n166 B 0.0269f
C186 VDD2.n167 B 0.0269f
C187 VDD2.n168 B 0.01205f
C188 VDD2.n169 B 0.011381f
C189 VDD2.n170 B 0.021179f
C190 VDD2.n171 B 0.021179f
C191 VDD2.n172 B 0.011381f
C192 VDD2.n173 B 0.01205f
C193 VDD2.n174 B 0.0269f
C194 VDD2.n175 B 0.0269f
C195 VDD2.n176 B 0.01205f
C196 VDD2.n177 B 0.011381f
C197 VDD2.n178 B 0.021179f
C198 VDD2.n179 B 0.021179f
C199 VDD2.n180 B 0.011381f
C200 VDD2.n181 B 0.01205f
C201 VDD2.n182 B 0.0269f
C202 VDD2.n183 B 0.0269f
C203 VDD2.n184 B 0.01205f
C204 VDD2.n185 B 0.011381f
C205 VDD2.n186 B 0.021179f
C206 VDD2.n187 B 0.021179f
C207 VDD2.n188 B 0.011381f
C208 VDD2.n189 B 0.01205f
C209 VDD2.n190 B 0.0269f
C210 VDD2.n191 B 0.0269f
C211 VDD2.n192 B 0.01205f
C212 VDD2.n193 B 0.011381f
C213 VDD2.n194 B 0.021179f
C214 VDD2.n195 B 0.05474f
C215 VDD2.n196 B 0.011381f
C216 VDD2.n197 B 0.01205f
C217 VDD2.n198 B 0.05419f
C218 VDD2.n199 B 0.060526f
C219 VDD2.n200 B 2.5312f
C220 VDD2.t0 B 0.30259f
C221 VDD2.t2 B 0.30259f
C222 VDD2.n201 B 2.76868f
C223 VN.n0 B 0.030528f
C224 VN.t1 B 2.82159f
C225 VN.n1 B 0.022539f
C226 VN.n2 B 0.220207f
C227 VN.t4 B 2.82159f
C228 VN.t0 B 3.00509f
C229 VN.n3 B 1.01899f
C230 VN.n4 B 1.05597f
C231 VN.n5 B 0.042941f
C232 VN.n6 B 0.041839f
C233 VN.n7 B 0.023156f
C234 VN.n8 B 0.023156f
C235 VN.n9 B 0.023156f
C236 VN.n10 B 0.045886f
C237 VN.n11 B 0.033614f
C238 VN.n12 B 1.05679f
C239 VN.n13 B 0.03434f
C240 VN.n14 B 0.030528f
C241 VN.t2 B 2.82159f
C242 VN.n15 B 0.022539f
C243 VN.n16 B 0.220207f
C244 VN.t5 B 2.82159f
C245 VN.t3 B 3.00509f
C246 VN.n17 B 1.01899f
C247 VN.n18 B 1.05597f
C248 VN.n19 B 0.042941f
C249 VN.n20 B 0.041839f
C250 VN.n21 B 0.023156f
C251 VN.n22 B 0.023156f
C252 VN.n23 B 0.023156f
C253 VN.n24 B 0.045886f
C254 VN.n25 B 0.033614f
C255 VN.n26 B 1.05679f
C256 VN.n27 B 1.4011f
C257 VDD1.n0 B 0.012074f
C258 VDD1.n1 B 0.0272f
C259 VDD1.n2 B 0.012184f
C260 VDD1.n3 B 0.021415f
C261 VDD1.n4 B 0.011508f
C262 VDD1.n5 B 0.0272f
C263 VDD1.n6 B 0.012184f
C264 VDD1.n7 B 0.021415f
C265 VDD1.n8 B 0.011508f
C266 VDD1.n9 B 0.0272f
C267 VDD1.n10 B 0.012184f
C268 VDD1.n11 B 0.021415f
C269 VDD1.n12 B 0.011508f
C270 VDD1.n13 B 0.0272f
C271 VDD1.n14 B 0.012184f
C272 VDD1.n15 B 0.021415f
C273 VDD1.n16 B 0.011508f
C274 VDD1.n17 B 0.0272f
C275 VDD1.n18 B 0.012184f
C276 VDD1.n19 B 0.021415f
C277 VDD1.n20 B 0.011508f
C278 VDD1.n21 B 0.0272f
C279 VDD1.n22 B 0.012184f
C280 VDD1.n23 B 0.021415f
C281 VDD1.n24 B 0.011508f
C282 VDD1.n25 B 0.0272f
C283 VDD1.n26 B 0.0272f
C284 VDD1.n27 B 0.012184f
C285 VDD1.n28 B 0.021415f
C286 VDD1.n29 B 0.011508f
C287 VDD1.n30 B 0.0272f
C288 VDD1.n31 B 0.012184f
C289 VDD1.n32 B 0.204388f
C290 VDD1.t2 B 0.04664f
C291 VDD1.n33 B 0.0204f
C292 VDD1.n34 B 0.019228f
C293 VDD1.n35 B 0.011508f
C294 VDD1.n36 B 1.65948f
C295 VDD1.n37 B 0.021415f
C296 VDD1.n38 B 0.011508f
C297 VDD1.n39 B 0.012184f
C298 VDD1.n40 B 0.0272f
C299 VDD1.n41 B 0.0272f
C300 VDD1.n42 B 0.012184f
C301 VDD1.n43 B 0.011508f
C302 VDD1.n44 B 0.021415f
C303 VDD1.n45 B 0.021415f
C304 VDD1.n46 B 0.011508f
C305 VDD1.n47 B 0.012184f
C306 VDD1.n48 B 0.0272f
C307 VDD1.n49 B 0.0272f
C308 VDD1.n50 B 0.012184f
C309 VDD1.n51 B 0.011508f
C310 VDD1.n52 B 0.021415f
C311 VDD1.n53 B 0.021415f
C312 VDD1.n54 B 0.011508f
C313 VDD1.n55 B 0.011846f
C314 VDD1.n56 B 0.011846f
C315 VDD1.n57 B 0.0272f
C316 VDD1.n58 B 0.0272f
C317 VDD1.n59 B 0.012184f
C318 VDD1.n60 B 0.011508f
C319 VDD1.n61 B 0.021415f
C320 VDD1.n62 B 0.021415f
C321 VDD1.n63 B 0.011508f
C322 VDD1.n64 B 0.012184f
C323 VDD1.n65 B 0.0272f
C324 VDD1.n66 B 0.0272f
C325 VDD1.n67 B 0.012184f
C326 VDD1.n68 B 0.011508f
C327 VDD1.n69 B 0.021415f
C328 VDD1.n70 B 0.021415f
C329 VDD1.n71 B 0.011508f
C330 VDD1.n72 B 0.012184f
C331 VDD1.n73 B 0.0272f
C332 VDD1.n74 B 0.0272f
C333 VDD1.n75 B 0.012184f
C334 VDD1.n76 B 0.011508f
C335 VDD1.n77 B 0.021415f
C336 VDD1.n78 B 0.021415f
C337 VDD1.n79 B 0.011508f
C338 VDD1.n80 B 0.012184f
C339 VDD1.n81 B 0.0272f
C340 VDD1.n82 B 0.0272f
C341 VDD1.n83 B 0.012184f
C342 VDD1.n84 B 0.011508f
C343 VDD1.n85 B 0.021415f
C344 VDD1.n86 B 0.021415f
C345 VDD1.n87 B 0.011508f
C346 VDD1.n88 B 0.012184f
C347 VDD1.n89 B 0.0272f
C348 VDD1.n90 B 0.0272f
C349 VDD1.n91 B 0.012184f
C350 VDD1.n92 B 0.011508f
C351 VDD1.n93 B 0.021415f
C352 VDD1.n94 B 0.055351f
C353 VDD1.n95 B 0.011508f
C354 VDD1.n96 B 0.012184f
C355 VDD1.n97 B 0.054794f
C356 VDD1.n98 B 0.067161f
C357 VDD1.n99 B 0.012074f
C358 VDD1.n100 B 0.0272f
C359 VDD1.n101 B 0.012184f
C360 VDD1.n102 B 0.021415f
C361 VDD1.n103 B 0.011508f
C362 VDD1.n104 B 0.0272f
C363 VDD1.n105 B 0.012184f
C364 VDD1.n106 B 0.021415f
C365 VDD1.n107 B 0.011508f
C366 VDD1.n108 B 0.0272f
C367 VDD1.n109 B 0.012184f
C368 VDD1.n110 B 0.021415f
C369 VDD1.n111 B 0.011508f
C370 VDD1.n112 B 0.0272f
C371 VDD1.n113 B 0.012184f
C372 VDD1.n114 B 0.021415f
C373 VDD1.n115 B 0.011508f
C374 VDD1.n116 B 0.0272f
C375 VDD1.n117 B 0.012184f
C376 VDD1.n118 B 0.021415f
C377 VDD1.n119 B 0.011508f
C378 VDD1.n120 B 0.0272f
C379 VDD1.n121 B 0.012184f
C380 VDD1.n122 B 0.021415f
C381 VDD1.n123 B 0.011508f
C382 VDD1.n124 B 0.0272f
C383 VDD1.n125 B 0.012184f
C384 VDD1.n126 B 0.021415f
C385 VDD1.n127 B 0.011508f
C386 VDD1.n128 B 0.0272f
C387 VDD1.n129 B 0.012184f
C388 VDD1.n130 B 0.204388f
C389 VDD1.t4 B 0.04664f
C390 VDD1.n131 B 0.0204f
C391 VDD1.n132 B 0.019228f
C392 VDD1.n133 B 0.011508f
C393 VDD1.n134 B 1.65948f
C394 VDD1.n135 B 0.021415f
C395 VDD1.n136 B 0.011508f
C396 VDD1.n137 B 0.012184f
C397 VDD1.n138 B 0.0272f
C398 VDD1.n139 B 0.0272f
C399 VDD1.n140 B 0.012184f
C400 VDD1.n141 B 0.011508f
C401 VDD1.n142 B 0.021415f
C402 VDD1.n143 B 0.021415f
C403 VDD1.n144 B 0.011508f
C404 VDD1.n145 B 0.012184f
C405 VDD1.n146 B 0.0272f
C406 VDD1.n147 B 0.0272f
C407 VDD1.n148 B 0.0272f
C408 VDD1.n149 B 0.012184f
C409 VDD1.n150 B 0.011508f
C410 VDD1.n151 B 0.021415f
C411 VDD1.n152 B 0.021415f
C412 VDD1.n153 B 0.011508f
C413 VDD1.n154 B 0.011846f
C414 VDD1.n155 B 0.011846f
C415 VDD1.n156 B 0.0272f
C416 VDD1.n157 B 0.0272f
C417 VDD1.n158 B 0.012184f
C418 VDD1.n159 B 0.011508f
C419 VDD1.n160 B 0.021415f
C420 VDD1.n161 B 0.021415f
C421 VDD1.n162 B 0.011508f
C422 VDD1.n163 B 0.012184f
C423 VDD1.n164 B 0.0272f
C424 VDD1.n165 B 0.0272f
C425 VDD1.n166 B 0.012184f
C426 VDD1.n167 B 0.011508f
C427 VDD1.n168 B 0.021415f
C428 VDD1.n169 B 0.021415f
C429 VDD1.n170 B 0.011508f
C430 VDD1.n171 B 0.012184f
C431 VDD1.n172 B 0.0272f
C432 VDD1.n173 B 0.0272f
C433 VDD1.n174 B 0.012184f
C434 VDD1.n175 B 0.011508f
C435 VDD1.n176 B 0.021415f
C436 VDD1.n177 B 0.021415f
C437 VDD1.n178 B 0.011508f
C438 VDD1.n179 B 0.012184f
C439 VDD1.n180 B 0.0272f
C440 VDD1.n181 B 0.0272f
C441 VDD1.n182 B 0.012184f
C442 VDD1.n183 B 0.011508f
C443 VDD1.n184 B 0.021415f
C444 VDD1.n185 B 0.021415f
C445 VDD1.n186 B 0.011508f
C446 VDD1.n187 B 0.012184f
C447 VDD1.n188 B 0.0272f
C448 VDD1.n189 B 0.0272f
C449 VDD1.n190 B 0.012184f
C450 VDD1.n191 B 0.011508f
C451 VDD1.n192 B 0.021415f
C452 VDD1.n193 B 0.055351f
C453 VDD1.n194 B 0.011508f
C454 VDD1.n195 B 0.012184f
C455 VDD1.n196 B 0.054794f
C456 VDD1.n197 B 0.066562f
C457 VDD1.t0 B 0.305965f
C458 VDD1.t3 B 0.305965f
C459 VDD1.n198 B 2.79959f
C460 VDD1.n199 B 2.66586f
C461 VDD1.t1 B 0.305965f
C462 VDD1.t5 B 0.305965f
C463 VDD1.n200 B 2.79638f
C464 VDD1.n201 B 2.74135f
C465 VTAIL.t3 B 0.321293f
C466 VTAIL.t10 B 0.321293f
C467 VTAIL.n0 B 2.87525f
C468 VTAIL.n1 B 0.377063f
C469 VTAIL.n2 B 0.012679f
C470 VTAIL.n3 B 0.028562f
C471 VTAIL.n4 B 0.012795f
C472 VTAIL.n5 B 0.022488f
C473 VTAIL.n6 B 0.012084f
C474 VTAIL.n7 B 0.028562f
C475 VTAIL.n8 B 0.012795f
C476 VTAIL.n9 B 0.022488f
C477 VTAIL.n10 B 0.012084f
C478 VTAIL.n11 B 0.028562f
C479 VTAIL.n12 B 0.012795f
C480 VTAIL.n13 B 0.022488f
C481 VTAIL.n14 B 0.012084f
C482 VTAIL.n15 B 0.028562f
C483 VTAIL.n16 B 0.012795f
C484 VTAIL.n17 B 0.022488f
C485 VTAIL.n18 B 0.012084f
C486 VTAIL.n19 B 0.028562f
C487 VTAIL.n20 B 0.012795f
C488 VTAIL.n21 B 0.022488f
C489 VTAIL.n22 B 0.012084f
C490 VTAIL.n23 B 0.028562f
C491 VTAIL.n24 B 0.012795f
C492 VTAIL.n25 B 0.022488f
C493 VTAIL.n26 B 0.012084f
C494 VTAIL.n27 B 0.028562f
C495 VTAIL.n28 B 0.012795f
C496 VTAIL.n29 B 0.022488f
C497 VTAIL.n30 B 0.012084f
C498 VTAIL.n31 B 0.028562f
C499 VTAIL.n32 B 0.012795f
C500 VTAIL.n33 B 0.214627f
C501 VTAIL.t8 B 0.048976f
C502 VTAIL.n34 B 0.021422f
C503 VTAIL.n35 B 0.020191f
C504 VTAIL.n36 B 0.012084f
C505 VTAIL.n37 B 1.74262f
C506 VTAIL.n38 B 0.022488f
C507 VTAIL.n39 B 0.012084f
C508 VTAIL.n40 B 0.012795f
C509 VTAIL.n41 B 0.028562f
C510 VTAIL.n42 B 0.028562f
C511 VTAIL.n43 B 0.012795f
C512 VTAIL.n44 B 0.012084f
C513 VTAIL.n45 B 0.022488f
C514 VTAIL.n46 B 0.022488f
C515 VTAIL.n47 B 0.012084f
C516 VTAIL.n48 B 0.012795f
C517 VTAIL.n49 B 0.028562f
C518 VTAIL.n50 B 0.028562f
C519 VTAIL.n51 B 0.028562f
C520 VTAIL.n52 B 0.012795f
C521 VTAIL.n53 B 0.012084f
C522 VTAIL.n54 B 0.022488f
C523 VTAIL.n55 B 0.022488f
C524 VTAIL.n56 B 0.012084f
C525 VTAIL.n57 B 0.01244f
C526 VTAIL.n58 B 0.01244f
C527 VTAIL.n59 B 0.028562f
C528 VTAIL.n60 B 0.028562f
C529 VTAIL.n61 B 0.012795f
C530 VTAIL.n62 B 0.012084f
C531 VTAIL.n63 B 0.022488f
C532 VTAIL.n64 B 0.022488f
C533 VTAIL.n65 B 0.012084f
C534 VTAIL.n66 B 0.012795f
C535 VTAIL.n67 B 0.028562f
C536 VTAIL.n68 B 0.028562f
C537 VTAIL.n69 B 0.012795f
C538 VTAIL.n70 B 0.012084f
C539 VTAIL.n71 B 0.022488f
C540 VTAIL.n72 B 0.022488f
C541 VTAIL.n73 B 0.012084f
C542 VTAIL.n74 B 0.012795f
C543 VTAIL.n75 B 0.028562f
C544 VTAIL.n76 B 0.028562f
C545 VTAIL.n77 B 0.012795f
C546 VTAIL.n78 B 0.012084f
C547 VTAIL.n79 B 0.022488f
C548 VTAIL.n80 B 0.022488f
C549 VTAIL.n81 B 0.012084f
C550 VTAIL.n82 B 0.012795f
C551 VTAIL.n83 B 0.028562f
C552 VTAIL.n84 B 0.028562f
C553 VTAIL.n85 B 0.012795f
C554 VTAIL.n86 B 0.012084f
C555 VTAIL.n87 B 0.022488f
C556 VTAIL.n88 B 0.022488f
C557 VTAIL.n89 B 0.012084f
C558 VTAIL.n90 B 0.012795f
C559 VTAIL.n91 B 0.028562f
C560 VTAIL.n92 B 0.028562f
C561 VTAIL.n93 B 0.012795f
C562 VTAIL.n94 B 0.012084f
C563 VTAIL.n95 B 0.022488f
C564 VTAIL.n96 B 0.058124f
C565 VTAIL.n97 B 0.012084f
C566 VTAIL.n98 B 0.012795f
C567 VTAIL.n99 B 0.05754f
C568 VTAIL.n100 B 0.048771f
C569 VTAIL.n101 B 0.316168f
C570 VTAIL.t7 B 0.321293f
C571 VTAIL.t9 B 0.321293f
C572 VTAIL.n102 B 2.87525f
C573 VTAIL.n103 B 2.1644f
C574 VTAIL.t1 B 0.321293f
C575 VTAIL.t2 B 0.321293f
C576 VTAIL.n104 B 2.87526f
C577 VTAIL.n105 B 2.16439f
C578 VTAIL.n106 B 0.012679f
C579 VTAIL.n107 B 0.028562f
C580 VTAIL.n108 B 0.012795f
C581 VTAIL.n109 B 0.022488f
C582 VTAIL.n110 B 0.012084f
C583 VTAIL.n111 B 0.028562f
C584 VTAIL.n112 B 0.012795f
C585 VTAIL.n113 B 0.022488f
C586 VTAIL.n114 B 0.012084f
C587 VTAIL.n115 B 0.028562f
C588 VTAIL.n116 B 0.012795f
C589 VTAIL.n117 B 0.022488f
C590 VTAIL.n118 B 0.012084f
C591 VTAIL.n119 B 0.028562f
C592 VTAIL.n120 B 0.012795f
C593 VTAIL.n121 B 0.022488f
C594 VTAIL.n122 B 0.012084f
C595 VTAIL.n123 B 0.028562f
C596 VTAIL.n124 B 0.012795f
C597 VTAIL.n125 B 0.022488f
C598 VTAIL.n126 B 0.012084f
C599 VTAIL.n127 B 0.028562f
C600 VTAIL.n128 B 0.012795f
C601 VTAIL.n129 B 0.022488f
C602 VTAIL.n130 B 0.012084f
C603 VTAIL.n131 B 0.028562f
C604 VTAIL.n132 B 0.028562f
C605 VTAIL.n133 B 0.012795f
C606 VTAIL.n134 B 0.022488f
C607 VTAIL.n135 B 0.012084f
C608 VTAIL.n136 B 0.028562f
C609 VTAIL.n137 B 0.012795f
C610 VTAIL.n138 B 0.214627f
C611 VTAIL.t11 B 0.048976f
C612 VTAIL.n139 B 0.021422f
C613 VTAIL.n140 B 0.020191f
C614 VTAIL.n141 B 0.012084f
C615 VTAIL.n142 B 1.74262f
C616 VTAIL.n143 B 0.022488f
C617 VTAIL.n144 B 0.012084f
C618 VTAIL.n145 B 0.012795f
C619 VTAIL.n146 B 0.028562f
C620 VTAIL.n147 B 0.028562f
C621 VTAIL.n148 B 0.012795f
C622 VTAIL.n149 B 0.012084f
C623 VTAIL.n150 B 0.022488f
C624 VTAIL.n151 B 0.022488f
C625 VTAIL.n152 B 0.012084f
C626 VTAIL.n153 B 0.012795f
C627 VTAIL.n154 B 0.028562f
C628 VTAIL.n155 B 0.028562f
C629 VTAIL.n156 B 0.012795f
C630 VTAIL.n157 B 0.012084f
C631 VTAIL.n158 B 0.022488f
C632 VTAIL.n159 B 0.022488f
C633 VTAIL.n160 B 0.012084f
C634 VTAIL.n161 B 0.01244f
C635 VTAIL.n162 B 0.01244f
C636 VTAIL.n163 B 0.028562f
C637 VTAIL.n164 B 0.028562f
C638 VTAIL.n165 B 0.012795f
C639 VTAIL.n166 B 0.012084f
C640 VTAIL.n167 B 0.022488f
C641 VTAIL.n168 B 0.022488f
C642 VTAIL.n169 B 0.012084f
C643 VTAIL.n170 B 0.012795f
C644 VTAIL.n171 B 0.028562f
C645 VTAIL.n172 B 0.028562f
C646 VTAIL.n173 B 0.012795f
C647 VTAIL.n174 B 0.012084f
C648 VTAIL.n175 B 0.022488f
C649 VTAIL.n176 B 0.022488f
C650 VTAIL.n177 B 0.012084f
C651 VTAIL.n178 B 0.012795f
C652 VTAIL.n179 B 0.028562f
C653 VTAIL.n180 B 0.028562f
C654 VTAIL.n181 B 0.012795f
C655 VTAIL.n182 B 0.012084f
C656 VTAIL.n183 B 0.022488f
C657 VTAIL.n184 B 0.022488f
C658 VTAIL.n185 B 0.012084f
C659 VTAIL.n186 B 0.012795f
C660 VTAIL.n187 B 0.028562f
C661 VTAIL.n188 B 0.028562f
C662 VTAIL.n189 B 0.012795f
C663 VTAIL.n190 B 0.012084f
C664 VTAIL.n191 B 0.022488f
C665 VTAIL.n192 B 0.022488f
C666 VTAIL.n193 B 0.012084f
C667 VTAIL.n194 B 0.012795f
C668 VTAIL.n195 B 0.028562f
C669 VTAIL.n196 B 0.028562f
C670 VTAIL.n197 B 0.012795f
C671 VTAIL.n198 B 0.012084f
C672 VTAIL.n199 B 0.022488f
C673 VTAIL.n200 B 0.058124f
C674 VTAIL.n201 B 0.012084f
C675 VTAIL.n202 B 0.012795f
C676 VTAIL.n203 B 0.05754f
C677 VTAIL.n204 B 0.048771f
C678 VTAIL.n205 B 0.316168f
C679 VTAIL.t5 B 0.321293f
C680 VTAIL.t6 B 0.321293f
C681 VTAIL.n206 B 2.87526f
C682 VTAIL.n207 B 0.503083f
C683 VTAIL.n208 B 0.012679f
C684 VTAIL.n209 B 0.028562f
C685 VTAIL.n210 B 0.012795f
C686 VTAIL.n211 B 0.022488f
C687 VTAIL.n212 B 0.012084f
C688 VTAIL.n213 B 0.028562f
C689 VTAIL.n214 B 0.012795f
C690 VTAIL.n215 B 0.022488f
C691 VTAIL.n216 B 0.012084f
C692 VTAIL.n217 B 0.028562f
C693 VTAIL.n218 B 0.012795f
C694 VTAIL.n219 B 0.022488f
C695 VTAIL.n220 B 0.012084f
C696 VTAIL.n221 B 0.028562f
C697 VTAIL.n222 B 0.012795f
C698 VTAIL.n223 B 0.022488f
C699 VTAIL.n224 B 0.012084f
C700 VTAIL.n225 B 0.028562f
C701 VTAIL.n226 B 0.012795f
C702 VTAIL.n227 B 0.022488f
C703 VTAIL.n228 B 0.012084f
C704 VTAIL.n229 B 0.028562f
C705 VTAIL.n230 B 0.012795f
C706 VTAIL.n231 B 0.022488f
C707 VTAIL.n232 B 0.012084f
C708 VTAIL.n233 B 0.028562f
C709 VTAIL.n234 B 0.028562f
C710 VTAIL.n235 B 0.012795f
C711 VTAIL.n236 B 0.022488f
C712 VTAIL.n237 B 0.012084f
C713 VTAIL.n238 B 0.028562f
C714 VTAIL.n239 B 0.012795f
C715 VTAIL.n240 B 0.214627f
C716 VTAIL.t4 B 0.048976f
C717 VTAIL.n241 B 0.021422f
C718 VTAIL.n242 B 0.020191f
C719 VTAIL.n243 B 0.012084f
C720 VTAIL.n244 B 1.74262f
C721 VTAIL.n245 B 0.022488f
C722 VTAIL.n246 B 0.012084f
C723 VTAIL.n247 B 0.012795f
C724 VTAIL.n248 B 0.028562f
C725 VTAIL.n249 B 0.028562f
C726 VTAIL.n250 B 0.012795f
C727 VTAIL.n251 B 0.012084f
C728 VTAIL.n252 B 0.022488f
C729 VTAIL.n253 B 0.022488f
C730 VTAIL.n254 B 0.012084f
C731 VTAIL.n255 B 0.012795f
C732 VTAIL.n256 B 0.028562f
C733 VTAIL.n257 B 0.028562f
C734 VTAIL.n258 B 0.012795f
C735 VTAIL.n259 B 0.012084f
C736 VTAIL.n260 B 0.022488f
C737 VTAIL.n261 B 0.022488f
C738 VTAIL.n262 B 0.012084f
C739 VTAIL.n263 B 0.01244f
C740 VTAIL.n264 B 0.01244f
C741 VTAIL.n265 B 0.028562f
C742 VTAIL.n266 B 0.028562f
C743 VTAIL.n267 B 0.012795f
C744 VTAIL.n268 B 0.012084f
C745 VTAIL.n269 B 0.022488f
C746 VTAIL.n270 B 0.022488f
C747 VTAIL.n271 B 0.012084f
C748 VTAIL.n272 B 0.012795f
C749 VTAIL.n273 B 0.028562f
C750 VTAIL.n274 B 0.028562f
C751 VTAIL.n275 B 0.012795f
C752 VTAIL.n276 B 0.012084f
C753 VTAIL.n277 B 0.022488f
C754 VTAIL.n278 B 0.022488f
C755 VTAIL.n279 B 0.012084f
C756 VTAIL.n280 B 0.012795f
C757 VTAIL.n281 B 0.028562f
C758 VTAIL.n282 B 0.028562f
C759 VTAIL.n283 B 0.012795f
C760 VTAIL.n284 B 0.012084f
C761 VTAIL.n285 B 0.022488f
C762 VTAIL.n286 B 0.022488f
C763 VTAIL.n287 B 0.012084f
C764 VTAIL.n288 B 0.012795f
C765 VTAIL.n289 B 0.028562f
C766 VTAIL.n290 B 0.028562f
C767 VTAIL.n291 B 0.012795f
C768 VTAIL.n292 B 0.012084f
C769 VTAIL.n293 B 0.022488f
C770 VTAIL.n294 B 0.022488f
C771 VTAIL.n295 B 0.012084f
C772 VTAIL.n296 B 0.012795f
C773 VTAIL.n297 B 0.028562f
C774 VTAIL.n298 B 0.028562f
C775 VTAIL.n299 B 0.012795f
C776 VTAIL.n300 B 0.012084f
C777 VTAIL.n301 B 0.022488f
C778 VTAIL.n302 B 0.058124f
C779 VTAIL.n303 B 0.012084f
C780 VTAIL.n304 B 0.012795f
C781 VTAIL.n305 B 0.05754f
C782 VTAIL.n306 B 0.048771f
C783 VTAIL.n307 B 1.80382f
C784 VTAIL.n308 B 0.012679f
C785 VTAIL.n309 B 0.028562f
C786 VTAIL.n310 B 0.012795f
C787 VTAIL.n311 B 0.022488f
C788 VTAIL.n312 B 0.012084f
C789 VTAIL.n313 B 0.028562f
C790 VTAIL.n314 B 0.012795f
C791 VTAIL.n315 B 0.022488f
C792 VTAIL.n316 B 0.012084f
C793 VTAIL.n317 B 0.028562f
C794 VTAIL.n318 B 0.012795f
C795 VTAIL.n319 B 0.022488f
C796 VTAIL.n320 B 0.012084f
C797 VTAIL.n321 B 0.028562f
C798 VTAIL.n322 B 0.012795f
C799 VTAIL.n323 B 0.022488f
C800 VTAIL.n324 B 0.012084f
C801 VTAIL.n325 B 0.028562f
C802 VTAIL.n326 B 0.012795f
C803 VTAIL.n327 B 0.022488f
C804 VTAIL.n328 B 0.012084f
C805 VTAIL.n329 B 0.028562f
C806 VTAIL.n330 B 0.012795f
C807 VTAIL.n331 B 0.022488f
C808 VTAIL.n332 B 0.012084f
C809 VTAIL.n333 B 0.028562f
C810 VTAIL.n334 B 0.012795f
C811 VTAIL.n335 B 0.022488f
C812 VTAIL.n336 B 0.012084f
C813 VTAIL.n337 B 0.028562f
C814 VTAIL.n338 B 0.012795f
C815 VTAIL.n339 B 0.214627f
C816 VTAIL.t0 B 0.048976f
C817 VTAIL.n340 B 0.021422f
C818 VTAIL.n341 B 0.020191f
C819 VTAIL.n342 B 0.012084f
C820 VTAIL.n343 B 1.74262f
C821 VTAIL.n344 B 0.022488f
C822 VTAIL.n345 B 0.012084f
C823 VTAIL.n346 B 0.012795f
C824 VTAIL.n347 B 0.028562f
C825 VTAIL.n348 B 0.028562f
C826 VTAIL.n349 B 0.012795f
C827 VTAIL.n350 B 0.012084f
C828 VTAIL.n351 B 0.022488f
C829 VTAIL.n352 B 0.022488f
C830 VTAIL.n353 B 0.012084f
C831 VTAIL.n354 B 0.012795f
C832 VTAIL.n355 B 0.028562f
C833 VTAIL.n356 B 0.028562f
C834 VTAIL.n357 B 0.028562f
C835 VTAIL.n358 B 0.012795f
C836 VTAIL.n359 B 0.012084f
C837 VTAIL.n360 B 0.022488f
C838 VTAIL.n361 B 0.022488f
C839 VTAIL.n362 B 0.012084f
C840 VTAIL.n363 B 0.01244f
C841 VTAIL.n364 B 0.01244f
C842 VTAIL.n365 B 0.028562f
C843 VTAIL.n366 B 0.028562f
C844 VTAIL.n367 B 0.012795f
C845 VTAIL.n368 B 0.012084f
C846 VTAIL.n369 B 0.022488f
C847 VTAIL.n370 B 0.022488f
C848 VTAIL.n371 B 0.012084f
C849 VTAIL.n372 B 0.012795f
C850 VTAIL.n373 B 0.028562f
C851 VTAIL.n374 B 0.028562f
C852 VTAIL.n375 B 0.012795f
C853 VTAIL.n376 B 0.012084f
C854 VTAIL.n377 B 0.022488f
C855 VTAIL.n378 B 0.022488f
C856 VTAIL.n379 B 0.012084f
C857 VTAIL.n380 B 0.012795f
C858 VTAIL.n381 B 0.028562f
C859 VTAIL.n382 B 0.028562f
C860 VTAIL.n383 B 0.012795f
C861 VTAIL.n384 B 0.012084f
C862 VTAIL.n385 B 0.022488f
C863 VTAIL.n386 B 0.022488f
C864 VTAIL.n387 B 0.012084f
C865 VTAIL.n388 B 0.012795f
C866 VTAIL.n389 B 0.028562f
C867 VTAIL.n390 B 0.028562f
C868 VTAIL.n391 B 0.012795f
C869 VTAIL.n392 B 0.012084f
C870 VTAIL.n393 B 0.022488f
C871 VTAIL.n394 B 0.022488f
C872 VTAIL.n395 B 0.012084f
C873 VTAIL.n396 B 0.012795f
C874 VTAIL.n397 B 0.028562f
C875 VTAIL.n398 B 0.028562f
C876 VTAIL.n399 B 0.012795f
C877 VTAIL.n400 B 0.012084f
C878 VTAIL.n401 B 0.022488f
C879 VTAIL.n402 B 0.058124f
C880 VTAIL.n403 B 0.012084f
C881 VTAIL.n404 B 0.012795f
C882 VTAIL.n405 B 0.05754f
C883 VTAIL.n406 B 0.048771f
C884 VTAIL.n407 B 1.75619f
C885 VP.n0 B 0.030899f
C886 VP.t2 B 2.85588f
C887 VP.n1 B 0.022813f
C888 VP.n2 B 0.023438f
C889 VP.t5 B 2.85588f
C890 VP.n3 B 0.043463f
C891 VP.n4 B 0.023438f
C892 VP.n5 B 0.034022f
C893 VP.n6 B 0.030899f
C894 VP.t0 B 2.85588f
C895 VP.n7 B 0.022813f
C896 VP.n8 B 0.222882f
C897 VP.t4 B 2.85588f
C898 VP.t3 B 3.04161f
C899 VP.n9 B 1.03137f
C900 VP.n10 B 1.06881f
C901 VP.n11 B 0.043463f
C902 VP.n12 B 0.042347f
C903 VP.n13 B 0.023438f
C904 VP.n14 B 0.023438f
C905 VP.n15 B 0.023438f
C906 VP.n16 B 0.046443f
C907 VP.n17 B 0.034022f
C908 VP.n18 B 1.06963f
C909 VP.n19 B 1.40564f
C910 VP.t1 B 2.85588f
C911 VP.n20 B 1.06963f
C912 VP.n21 B 1.42166f
C913 VP.n22 B 0.030899f
C914 VP.n23 B 0.023438f
C915 VP.n24 B 0.046443f
C916 VP.n25 B 0.022813f
C917 VP.n26 B 0.042347f
C918 VP.n27 B 0.023438f
C919 VP.n28 B 0.023438f
C920 VP.n29 B 0.023438f
C921 VP.n30 B 1.0133f
C922 VP.n31 B 0.043463f
C923 VP.n32 B 0.042347f
C924 VP.n33 B 0.023438f
C925 VP.n34 B 0.023438f
C926 VP.n35 B 0.023438f
C927 VP.n36 B 0.046443f
C928 VP.n37 B 0.034022f
C929 VP.n38 B 1.06963f
C930 VP.n39 B 0.034757f
.ends

