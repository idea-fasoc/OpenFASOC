* NGSPICE file created from diff_pair_sample_0145.ext - technology: sky130A

.subckt diff_pair_sample_0145 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=0 ps=0 w=6.85 l=0.73
X1 VTAIL.t7 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=1.13025 ps=7.18 w=6.85 l=0.73
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=0 ps=0 w=6.85 l=0.73
X3 VDD2.t2 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.13025 pd=7.18 as=2.6715 ps=14.48 w=6.85 l=0.73
X4 VTAIL.t0 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=1.13025 ps=7.18 w=6.85 l=0.73
X5 VTAIL.t5 VN.t2 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=1.13025 ps=7.18 w=6.85 l=0.73
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=0 ps=0 w=6.85 l=0.73
X7 VDD2.t1 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.13025 pd=7.18 as=2.6715 ps=14.48 w=6.85 l=0.73
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=0 ps=0 w=6.85 l=0.73
X9 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.13025 pd=7.18 as=2.6715 ps=14.48 w=6.85 l=0.73
X10 VTAIL.t2 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6715 pd=14.48 as=1.13025 ps=7.18 w=6.85 l=0.73
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.13025 pd=7.18 as=2.6715 ps=14.48 w=6.85 l=0.73
R0 B.n468 B.n467 585
R1 B.n469 B.n468 585
R2 B.n196 B.n67 585
R3 B.n195 B.n194 585
R4 B.n193 B.n192 585
R5 B.n191 B.n190 585
R6 B.n189 B.n188 585
R7 B.n187 B.n186 585
R8 B.n185 B.n184 585
R9 B.n183 B.n182 585
R10 B.n181 B.n180 585
R11 B.n179 B.n178 585
R12 B.n177 B.n176 585
R13 B.n175 B.n174 585
R14 B.n173 B.n172 585
R15 B.n171 B.n170 585
R16 B.n169 B.n168 585
R17 B.n167 B.n166 585
R18 B.n165 B.n164 585
R19 B.n163 B.n162 585
R20 B.n161 B.n160 585
R21 B.n159 B.n158 585
R22 B.n157 B.n156 585
R23 B.n155 B.n154 585
R24 B.n153 B.n152 585
R25 B.n151 B.n150 585
R26 B.n149 B.n148 585
R27 B.n147 B.n146 585
R28 B.n145 B.n144 585
R29 B.n143 B.n142 585
R30 B.n141 B.n140 585
R31 B.n139 B.n138 585
R32 B.n137 B.n136 585
R33 B.n135 B.n134 585
R34 B.n133 B.n132 585
R35 B.n131 B.n130 585
R36 B.n129 B.n128 585
R37 B.n126 B.n125 585
R38 B.n124 B.n123 585
R39 B.n122 B.n121 585
R40 B.n120 B.n119 585
R41 B.n118 B.n117 585
R42 B.n116 B.n115 585
R43 B.n114 B.n113 585
R44 B.n112 B.n111 585
R45 B.n110 B.n109 585
R46 B.n108 B.n107 585
R47 B.n106 B.n105 585
R48 B.n104 B.n103 585
R49 B.n102 B.n101 585
R50 B.n100 B.n99 585
R51 B.n98 B.n97 585
R52 B.n96 B.n95 585
R53 B.n94 B.n93 585
R54 B.n92 B.n91 585
R55 B.n90 B.n89 585
R56 B.n88 B.n87 585
R57 B.n86 B.n85 585
R58 B.n84 B.n83 585
R59 B.n82 B.n81 585
R60 B.n80 B.n79 585
R61 B.n78 B.n77 585
R62 B.n76 B.n75 585
R63 B.n74 B.n73 585
R64 B.n466 B.n35 585
R65 B.n470 B.n35 585
R66 B.n465 B.n34 585
R67 B.n471 B.n34 585
R68 B.n464 B.n463 585
R69 B.n463 B.n30 585
R70 B.n462 B.n29 585
R71 B.n477 B.n29 585
R72 B.n461 B.n28 585
R73 B.n478 B.n28 585
R74 B.n460 B.n27 585
R75 B.n479 B.n27 585
R76 B.n459 B.n458 585
R77 B.n458 B.n23 585
R78 B.n457 B.n22 585
R79 B.n485 B.n22 585
R80 B.n456 B.n21 585
R81 B.n486 B.n21 585
R82 B.n455 B.n20 585
R83 B.n487 B.n20 585
R84 B.n454 B.n453 585
R85 B.n453 B.n16 585
R86 B.n452 B.n15 585
R87 B.n493 B.n15 585
R88 B.n451 B.n14 585
R89 B.n494 B.n14 585
R90 B.n450 B.n13 585
R91 B.n495 B.n13 585
R92 B.n449 B.n448 585
R93 B.n448 B.n12 585
R94 B.n447 B.n446 585
R95 B.n447 B.n8 585
R96 B.n445 B.n7 585
R97 B.n502 B.n7 585
R98 B.n444 B.n6 585
R99 B.n503 B.n6 585
R100 B.n443 B.n5 585
R101 B.n504 B.n5 585
R102 B.n442 B.n441 585
R103 B.n441 B.n4 585
R104 B.n440 B.n197 585
R105 B.n440 B.n439 585
R106 B.n429 B.n198 585
R107 B.n432 B.n198 585
R108 B.n431 B.n430 585
R109 B.n433 B.n431 585
R110 B.n428 B.n203 585
R111 B.n203 B.n202 585
R112 B.n427 B.n426 585
R113 B.n426 B.n425 585
R114 B.n205 B.n204 585
R115 B.n206 B.n205 585
R116 B.n418 B.n417 585
R117 B.n419 B.n418 585
R118 B.n416 B.n211 585
R119 B.n211 B.n210 585
R120 B.n415 B.n414 585
R121 B.n414 B.n413 585
R122 B.n213 B.n212 585
R123 B.n214 B.n213 585
R124 B.n406 B.n405 585
R125 B.n407 B.n406 585
R126 B.n404 B.n218 585
R127 B.n222 B.n218 585
R128 B.n403 B.n402 585
R129 B.n402 B.n401 585
R130 B.n220 B.n219 585
R131 B.n221 B.n220 585
R132 B.n394 B.n393 585
R133 B.n395 B.n394 585
R134 B.n392 B.n227 585
R135 B.n227 B.n226 585
R136 B.n386 B.n385 585
R137 B.n384 B.n260 585
R138 B.n383 B.n259 585
R139 B.n388 B.n259 585
R140 B.n382 B.n381 585
R141 B.n380 B.n379 585
R142 B.n378 B.n377 585
R143 B.n376 B.n375 585
R144 B.n374 B.n373 585
R145 B.n372 B.n371 585
R146 B.n370 B.n369 585
R147 B.n368 B.n367 585
R148 B.n366 B.n365 585
R149 B.n364 B.n363 585
R150 B.n362 B.n361 585
R151 B.n360 B.n359 585
R152 B.n358 B.n357 585
R153 B.n356 B.n355 585
R154 B.n354 B.n353 585
R155 B.n352 B.n351 585
R156 B.n350 B.n349 585
R157 B.n348 B.n347 585
R158 B.n346 B.n345 585
R159 B.n344 B.n343 585
R160 B.n342 B.n341 585
R161 B.n340 B.n339 585
R162 B.n338 B.n337 585
R163 B.n336 B.n335 585
R164 B.n334 B.n333 585
R165 B.n332 B.n331 585
R166 B.n330 B.n329 585
R167 B.n328 B.n327 585
R168 B.n326 B.n325 585
R169 B.n324 B.n323 585
R170 B.n322 B.n321 585
R171 B.n320 B.n319 585
R172 B.n318 B.n317 585
R173 B.n315 B.n314 585
R174 B.n313 B.n312 585
R175 B.n311 B.n310 585
R176 B.n309 B.n308 585
R177 B.n307 B.n306 585
R178 B.n305 B.n304 585
R179 B.n303 B.n302 585
R180 B.n301 B.n300 585
R181 B.n299 B.n298 585
R182 B.n297 B.n296 585
R183 B.n295 B.n294 585
R184 B.n293 B.n292 585
R185 B.n291 B.n290 585
R186 B.n289 B.n288 585
R187 B.n287 B.n286 585
R188 B.n285 B.n284 585
R189 B.n283 B.n282 585
R190 B.n281 B.n280 585
R191 B.n279 B.n278 585
R192 B.n277 B.n276 585
R193 B.n275 B.n274 585
R194 B.n273 B.n272 585
R195 B.n271 B.n270 585
R196 B.n269 B.n268 585
R197 B.n267 B.n266 585
R198 B.n229 B.n228 585
R199 B.n391 B.n390 585
R200 B.n225 B.n224 585
R201 B.n226 B.n225 585
R202 B.n397 B.n396 585
R203 B.n396 B.n395 585
R204 B.n398 B.n223 585
R205 B.n223 B.n221 585
R206 B.n400 B.n399 585
R207 B.n401 B.n400 585
R208 B.n217 B.n216 585
R209 B.n222 B.n217 585
R210 B.n409 B.n408 585
R211 B.n408 B.n407 585
R212 B.n410 B.n215 585
R213 B.n215 B.n214 585
R214 B.n412 B.n411 585
R215 B.n413 B.n412 585
R216 B.n209 B.n208 585
R217 B.n210 B.n209 585
R218 B.n421 B.n420 585
R219 B.n420 B.n419 585
R220 B.n422 B.n207 585
R221 B.n207 B.n206 585
R222 B.n424 B.n423 585
R223 B.n425 B.n424 585
R224 B.n201 B.n200 585
R225 B.n202 B.n201 585
R226 B.n435 B.n434 585
R227 B.n434 B.n433 585
R228 B.n436 B.n199 585
R229 B.n432 B.n199 585
R230 B.n438 B.n437 585
R231 B.n439 B.n438 585
R232 B.n3 B.n0 585
R233 B.n4 B.n3 585
R234 B.n501 B.n1 585
R235 B.n502 B.n501 585
R236 B.n500 B.n499 585
R237 B.n500 B.n8 585
R238 B.n498 B.n9 585
R239 B.n12 B.n9 585
R240 B.n497 B.n496 585
R241 B.n496 B.n495 585
R242 B.n11 B.n10 585
R243 B.n494 B.n11 585
R244 B.n492 B.n491 585
R245 B.n493 B.n492 585
R246 B.n490 B.n17 585
R247 B.n17 B.n16 585
R248 B.n489 B.n488 585
R249 B.n488 B.n487 585
R250 B.n19 B.n18 585
R251 B.n486 B.n19 585
R252 B.n484 B.n483 585
R253 B.n485 B.n484 585
R254 B.n482 B.n24 585
R255 B.n24 B.n23 585
R256 B.n481 B.n480 585
R257 B.n480 B.n479 585
R258 B.n26 B.n25 585
R259 B.n478 B.n26 585
R260 B.n476 B.n475 585
R261 B.n477 B.n476 585
R262 B.n474 B.n31 585
R263 B.n31 B.n30 585
R264 B.n473 B.n472 585
R265 B.n472 B.n471 585
R266 B.n33 B.n32 585
R267 B.n470 B.n33 585
R268 B.n505 B.n504 585
R269 B.n503 B.n2 585
R270 B.n73 B.n33 454.062
R271 B.n468 B.n35 454.062
R272 B.n390 B.n227 454.062
R273 B.n386 B.n225 454.062
R274 B.n71 B.t15 428.755
R275 B.n68 B.t8 428.755
R276 B.n264 B.t4 428.755
R277 B.n261 B.t12 428.755
R278 B.n469 B.n66 256.663
R279 B.n469 B.n65 256.663
R280 B.n469 B.n64 256.663
R281 B.n469 B.n63 256.663
R282 B.n469 B.n62 256.663
R283 B.n469 B.n61 256.663
R284 B.n469 B.n60 256.663
R285 B.n469 B.n59 256.663
R286 B.n469 B.n58 256.663
R287 B.n469 B.n57 256.663
R288 B.n469 B.n56 256.663
R289 B.n469 B.n55 256.663
R290 B.n469 B.n54 256.663
R291 B.n469 B.n53 256.663
R292 B.n469 B.n52 256.663
R293 B.n469 B.n51 256.663
R294 B.n469 B.n50 256.663
R295 B.n469 B.n49 256.663
R296 B.n469 B.n48 256.663
R297 B.n469 B.n47 256.663
R298 B.n469 B.n46 256.663
R299 B.n469 B.n45 256.663
R300 B.n469 B.n44 256.663
R301 B.n469 B.n43 256.663
R302 B.n469 B.n42 256.663
R303 B.n469 B.n41 256.663
R304 B.n469 B.n40 256.663
R305 B.n469 B.n39 256.663
R306 B.n469 B.n38 256.663
R307 B.n469 B.n37 256.663
R308 B.n469 B.n36 256.663
R309 B.n388 B.n387 256.663
R310 B.n388 B.n230 256.663
R311 B.n388 B.n231 256.663
R312 B.n388 B.n232 256.663
R313 B.n388 B.n233 256.663
R314 B.n388 B.n234 256.663
R315 B.n388 B.n235 256.663
R316 B.n388 B.n236 256.663
R317 B.n388 B.n237 256.663
R318 B.n388 B.n238 256.663
R319 B.n388 B.n239 256.663
R320 B.n388 B.n240 256.663
R321 B.n388 B.n241 256.663
R322 B.n388 B.n242 256.663
R323 B.n388 B.n243 256.663
R324 B.n388 B.n244 256.663
R325 B.n388 B.n245 256.663
R326 B.n388 B.n246 256.663
R327 B.n388 B.n247 256.663
R328 B.n388 B.n248 256.663
R329 B.n388 B.n249 256.663
R330 B.n388 B.n250 256.663
R331 B.n388 B.n251 256.663
R332 B.n388 B.n252 256.663
R333 B.n388 B.n253 256.663
R334 B.n388 B.n254 256.663
R335 B.n388 B.n255 256.663
R336 B.n388 B.n256 256.663
R337 B.n388 B.n257 256.663
R338 B.n388 B.n258 256.663
R339 B.n389 B.n388 256.663
R340 B.n507 B.n506 256.663
R341 B.n77 B.n76 163.367
R342 B.n81 B.n80 163.367
R343 B.n85 B.n84 163.367
R344 B.n89 B.n88 163.367
R345 B.n93 B.n92 163.367
R346 B.n97 B.n96 163.367
R347 B.n101 B.n100 163.367
R348 B.n105 B.n104 163.367
R349 B.n109 B.n108 163.367
R350 B.n113 B.n112 163.367
R351 B.n117 B.n116 163.367
R352 B.n121 B.n120 163.367
R353 B.n125 B.n124 163.367
R354 B.n130 B.n129 163.367
R355 B.n134 B.n133 163.367
R356 B.n138 B.n137 163.367
R357 B.n142 B.n141 163.367
R358 B.n146 B.n145 163.367
R359 B.n150 B.n149 163.367
R360 B.n154 B.n153 163.367
R361 B.n158 B.n157 163.367
R362 B.n162 B.n161 163.367
R363 B.n166 B.n165 163.367
R364 B.n170 B.n169 163.367
R365 B.n174 B.n173 163.367
R366 B.n178 B.n177 163.367
R367 B.n182 B.n181 163.367
R368 B.n186 B.n185 163.367
R369 B.n190 B.n189 163.367
R370 B.n194 B.n193 163.367
R371 B.n468 B.n67 163.367
R372 B.n394 B.n227 163.367
R373 B.n394 B.n220 163.367
R374 B.n402 B.n220 163.367
R375 B.n402 B.n218 163.367
R376 B.n406 B.n218 163.367
R377 B.n406 B.n213 163.367
R378 B.n414 B.n213 163.367
R379 B.n414 B.n211 163.367
R380 B.n418 B.n211 163.367
R381 B.n418 B.n205 163.367
R382 B.n426 B.n205 163.367
R383 B.n426 B.n203 163.367
R384 B.n431 B.n203 163.367
R385 B.n431 B.n198 163.367
R386 B.n440 B.n198 163.367
R387 B.n441 B.n440 163.367
R388 B.n441 B.n5 163.367
R389 B.n6 B.n5 163.367
R390 B.n7 B.n6 163.367
R391 B.n447 B.n7 163.367
R392 B.n448 B.n447 163.367
R393 B.n448 B.n13 163.367
R394 B.n14 B.n13 163.367
R395 B.n15 B.n14 163.367
R396 B.n453 B.n15 163.367
R397 B.n453 B.n20 163.367
R398 B.n21 B.n20 163.367
R399 B.n22 B.n21 163.367
R400 B.n458 B.n22 163.367
R401 B.n458 B.n27 163.367
R402 B.n28 B.n27 163.367
R403 B.n29 B.n28 163.367
R404 B.n463 B.n29 163.367
R405 B.n463 B.n34 163.367
R406 B.n35 B.n34 163.367
R407 B.n260 B.n259 163.367
R408 B.n381 B.n259 163.367
R409 B.n379 B.n378 163.367
R410 B.n375 B.n374 163.367
R411 B.n371 B.n370 163.367
R412 B.n367 B.n366 163.367
R413 B.n363 B.n362 163.367
R414 B.n359 B.n358 163.367
R415 B.n355 B.n354 163.367
R416 B.n351 B.n350 163.367
R417 B.n347 B.n346 163.367
R418 B.n343 B.n342 163.367
R419 B.n339 B.n338 163.367
R420 B.n335 B.n334 163.367
R421 B.n331 B.n330 163.367
R422 B.n327 B.n326 163.367
R423 B.n323 B.n322 163.367
R424 B.n319 B.n318 163.367
R425 B.n314 B.n313 163.367
R426 B.n310 B.n309 163.367
R427 B.n306 B.n305 163.367
R428 B.n302 B.n301 163.367
R429 B.n298 B.n297 163.367
R430 B.n294 B.n293 163.367
R431 B.n290 B.n289 163.367
R432 B.n286 B.n285 163.367
R433 B.n282 B.n281 163.367
R434 B.n278 B.n277 163.367
R435 B.n274 B.n273 163.367
R436 B.n270 B.n269 163.367
R437 B.n266 B.n229 163.367
R438 B.n396 B.n225 163.367
R439 B.n396 B.n223 163.367
R440 B.n400 B.n223 163.367
R441 B.n400 B.n217 163.367
R442 B.n408 B.n217 163.367
R443 B.n408 B.n215 163.367
R444 B.n412 B.n215 163.367
R445 B.n412 B.n209 163.367
R446 B.n420 B.n209 163.367
R447 B.n420 B.n207 163.367
R448 B.n424 B.n207 163.367
R449 B.n424 B.n201 163.367
R450 B.n434 B.n201 163.367
R451 B.n434 B.n199 163.367
R452 B.n438 B.n199 163.367
R453 B.n438 B.n3 163.367
R454 B.n505 B.n3 163.367
R455 B.n501 B.n2 163.367
R456 B.n501 B.n500 163.367
R457 B.n500 B.n9 163.367
R458 B.n496 B.n9 163.367
R459 B.n496 B.n11 163.367
R460 B.n492 B.n11 163.367
R461 B.n492 B.n17 163.367
R462 B.n488 B.n17 163.367
R463 B.n488 B.n19 163.367
R464 B.n484 B.n19 163.367
R465 B.n484 B.n24 163.367
R466 B.n480 B.n24 163.367
R467 B.n480 B.n26 163.367
R468 B.n476 B.n26 163.367
R469 B.n476 B.n31 163.367
R470 B.n472 B.n31 163.367
R471 B.n472 B.n33 163.367
R472 B.n388 B.n226 109.773
R473 B.n470 B.n469 109.773
R474 B.n68 B.t10 90.5542
R475 B.n264 B.t7 90.5542
R476 B.n71 B.t16 90.5465
R477 B.n261 B.t14 90.5465
R478 B.n73 B.n36 71.676
R479 B.n77 B.n37 71.676
R480 B.n81 B.n38 71.676
R481 B.n85 B.n39 71.676
R482 B.n89 B.n40 71.676
R483 B.n93 B.n41 71.676
R484 B.n97 B.n42 71.676
R485 B.n101 B.n43 71.676
R486 B.n105 B.n44 71.676
R487 B.n109 B.n45 71.676
R488 B.n113 B.n46 71.676
R489 B.n117 B.n47 71.676
R490 B.n121 B.n48 71.676
R491 B.n125 B.n49 71.676
R492 B.n130 B.n50 71.676
R493 B.n134 B.n51 71.676
R494 B.n138 B.n52 71.676
R495 B.n142 B.n53 71.676
R496 B.n146 B.n54 71.676
R497 B.n150 B.n55 71.676
R498 B.n154 B.n56 71.676
R499 B.n158 B.n57 71.676
R500 B.n162 B.n58 71.676
R501 B.n166 B.n59 71.676
R502 B.n170 B.n60 71.676
R503 B.n174 B.n61 71.676
R504 B.n178 B.n62 71.676
R505 B.n182 B.n63 71.676
R506 B.n186 B.n64 71.676
R507 B.n190 B.n65 71.676
R508 B.n194 B.n66 71.676
R509 B.n67 B.n66 71.676
R510 B.n193 B.n65 71.676
R511 B.n189 B.n64 71.676
R512 B.n185 B.n63 71.676
R513 B.n181 B.n62 71.676
R514 B.n177 B.n61 71.676
R515 B.n173 B.n60 71.676
R516 B.n169 B.n59 71.676
R517 B.n165 B.n58 71.676
R518 B.n161 B.n57 71.676
R519 B.n157 B.n56 71.676
R520 B.n153 B.n55 71.676
R521 B.n149 B.n54 71.676
R522 B.n145 B.n53 71.676
R523 B.n141 B.n52 71.676
R524 B.n137 B.n51 71.676
R525 B.n133 B.n50 71.676
R526 B.n129 B.n49 71.676
R527 B.n124 B.n48 71.676
R528 B.n120 B.n47 71.676
R529 B.n116 B.n46 71.676
R530 B.n112 B.n45 71.676
R531 B.n108 B.n44 71.676
R532 B.n104 B.n43 71.676
R533 B.n100 B.n42 71.676
R534 B.n96 B.n41 71.676
R535 B.n92 B.n40 71.676
R536 B.n88 B.n39 71.676
R537 B.n84 B.n38 71.676
R538 B.n80 B.n37 71.676
R539 B.n76 B.n36 71.676
R540 B.n387 B.n386 71.676
R541 B.n381 B.n230 71.676
R542 B.n378 B.n231 71.676
R543 B.n374 B.n232 71.676
R544 B.n370 B.n233 71.676
R545 B.n366 B.n234 71.676
R546 B.n362 B.n235 71.676
R547 B.n358 B.n236 71.676
R548 B.n354 B.n237 71.676
R549 B.n350 B.n238 71.676
R550 B.n346 B.n239 71.676
R551 B.n342 B.n240 71.676
R552 B.n338 B.n241 71.676
R553 B.n334 B.n242 71.676
R554 B.n330 B.n243 71.676
R555 B.n326 B.n244 71.676
R556 B.n322 B.n245 71.676
R557 B.n318 B.n246 71.676
R558 B.n313 B.n247 71.676
R559 B.n309 B.n248 71.676
R560 B.n305 B.n249 71.676
R561 B.n301 B.n250 71.676
R562 B.n297 B.n251 71.676
R563 B.n293 B.n252 71.676
R564 B.n289 B.n253 71.676
R565 B.n285 B.n254 71.676
R566 B.n281 B.n255 71.676
R567 B.n277 B.n256 71.676
R568 B.n273 B.n257 71.676
R569 B.n269 B.n258 71.676
R570 B.n389 B.n229 71.676
R571 B.n387 B.n260 71.676
R572 B.n379 B.n230 71.676
R573 B.n375 B.n231 71.676
R574 B.n371 B.n232 71.676
R575 B.n367 B.n233 71.676
R576 B.n363 B.n234 71.676
R577 B.n359 B.n235 71.676
R578 B.n355 B.n236 71.676
R579 B.n351 B.n237 71.676
R580 B.n347 B.n238 71.676
R581 B.n343 B.n239 71.676
R582 B.n339 B.n240 71.676
R583 B.n335 B.n241 71.676
R584 B.n331 B.n242 71.676
R585 B.n327 B.n243 71.676
R586 B.n323 B.n244 71.676
R587 B.n319 B.n245 71.676
R588 B.n314 B.n246 71.676
R589 B.n310 B.n247 71.676
R590 B.n306 B.n248 71.676
R591 B.n302 B.n249 71.676
R592 B.n298 B.n250 71.676
R593 B.n294 B.n251 71.676
R594 B.n290 B.n252 71.676
R595 B.n286 B.n253 71.676
R596 B.n282 B.n254 71.676
R597 B.n278 B.n255 71.676
R598 B.n274 B.n256 71.676
R599 B.n270 B.n257 71.676
R600 B.n266 B.n258 71.676
R601 B.n390 B.n389 71.676
R602 B.n506 B.n505 71.676
R603 B.n506 B.n2 71.676
R604 B.n69 B.t11 69.9967
R605 B.n265 B.t6 69.9967
R606 B.n72 B.t17 69.9889
R607 B.n262 B.t13 69.9889
R608 B.n395 B.n226 61.6912
R609 B.n395 B.n221 61.6912
R610 B.n401 B.n221 61.6912
R611 B.n401 B.n222 61.6912
R612 B.n407 B.n214 61.6912
R613 B.n413 B.n214 61.6912
R614 B.n413 B.n210 61.6912
R615 B.n419 B.n210 61.6912
R616 B.n419 B.n206 61.6912
R617 B.n425 B.n206 61.6912
R618 B.n433 B.n202 61.6912
R619 B.n433 B.n432 61.6912
R620 B.n439 B.n4 61.6912
R621 B.n504 B.n4 61.6912
R622 B.n504 B.n503 61.6912
R623 B.n503 B.n502 61.6912
R624 B.n502 B.n8 61.6912
R625 B.n495 B.n12 61.6912
R626 B.n495 B.n494 61.6912
R627 B.n493 B.n16 61.6912
R628 B.n487 B.n16 61.6912
R629 B.n487 B.n486 61.6912
R630 B.n486 B.n485 61.6912
R631 B.n485 B.n23 61.6912
R632 B.n479 B.n23 61.6912
R633 B.n478 B.n477 61.6912
R634 B.n477 B.n30 61.6912
R635 B.n471 B.n30 61.6912
R636 B.n471 B.n470 61.6912
R637 B.n127 B.n72 59.5399
R638 B.n70 B.n69 59.5399
R639 B.n316 B.n265 59.5399
R640 B.n263 B.n262 59.5399
R641 B.n222 B.t5 55.3407
R642 B.t9 B.n478 55.3407
R643 B.t1 B.n202 48.083
R644 B.n494 B.t3 48.083
R645 B.n439 B.t0 40.8252
R646 B.t2 B.n8 40.8252
R647 B.n467 B.n466 29.5029
R648 B.n385 B.n224 29.5029
R649 B.n392 B.n391 29.5029
R650 B.n74 B.n32 29.5029
R651 B.n432 B.t0 20.8665
R652 B.n12 B.t2 20.8665
R653 B.n72 B.n71 20.5581
R654 B.n69 B.n68 20.5581
R655 B.n265 B.n264 20.5581
R656 B.n262 B.n261 20.5581
R657 B B.n507 18.0485
R658 B.n425 B.t1 13.6087
R659 B.t3 B.n493 13.6087
R660 B.n397 B.n224 10.6151
R661 B.n398 B.n397 10.6151
R662 B.n399 B.n398 10.6151
R663 B.n399 B.n216 10.6151
R664 B.n409 B.n216 10.6151
R665 B.n410 B.n409 10.6151
R666 B.n411 B.n410 10.6151
R667 B.n411 B.n208 10.6151
R668 B.n421 B.n208 10.6151
R669 B.n422 B.n421 10.6151
R670 B.n423 B.n422 10.6151
R671 B.n423 B.n200 10.6151
R672 B.n435 B.n200 10.6151
R673 B.n436 B.n435 10.6151
R674 B.n437 B.n436 10.6151
R675 B.n437 B.n0 10.6151
R676 B.n385 B.n384 10.6151
R677 B.n384 B.n383 10.6151
R678 B.n383 B.n382 10.6151
R679 B.n382 B.n380 10.6151
R680 B.n380 B.n377 10.6151
R681 B.n377 B.n376 10.6151
R682 B.n376 B.n373 10.6151
R683 B.n373 B.n372 10.6151
R684 B.n372 B.n369 10.6151
R685 B.n369 B.n368 10.6151
R686 B.n368 B.n365 10.6151
R687 B.n365 B.n364 10.6151
R688 B.n364 B.n361 10.6151
R689 B.n361 B.n360 10.6151
R690 B.n360 B.n357 10.6151
R691 B.n357 B.n356 10.6151
R692 B.n356 B.n353 10.6151
R693 B.n353 B.n352 10.6151
R694 B.n352 B.n349 10.6151
R695 B.n349 B.n348 10.6151
R696 B.n348 B.n345 10.6151
R697 B.n345 B.n344 10.6151
R698 B.n344 B.n341 10.6151
R699 B.n341 B.n340 10.6151
R700 B.n340 B.n337 10.6151
R701 B.n337 B.n336 10.6151
R702 B.n333 B.n332 10.6151
R703 B.n332 B.n329 10.6151
R704 B.n329 B.n328 10.6151
R705 B.n328 B.n325 10.6151
R706 B.n325 B.n324 10.6151
R707 B.n324 B.n321 10.6151
R708 B.n321 B.n320 10.6151
R709 B.n320 B.n317 10.6151
R710 B.n315 B.n312 10.6151
R711 B.n312 B.n311 10.6151
R712 B.n311 B.n308 10.6151
R713 B.n308 B.n307 10.6151
R714 B.n307 B.n304 10.6151
R715 B.n304 B.n303 10.6151
R716 B.n303 B.n300 10.6151
R717 B.n300 B.n299 10.6151
R718 B.n299 B.n296 10.6151
R719 B.n296 B.n295 10.6151
R720 B.n295 B.n292 10.6151
R721 B.n292 B.n291 10.6151
R722 B.n291 B.n288 10.6151
R723 B.n288 B.n287 10.6151
R724 B.n287 B.n284 10.6151
R725 B.n284 B.n283 10.6151
R726 B.n283 B.n280 10.6151
R727 B.n280 B.n279 10.6151
R728 B.n279 B.n276 10.6151
R729 B.n276 B.n275 10.6151
R730 B.n275 B.n272 10.6151
R731 B.n272 B.n271 10.6151
R732 B.n271 B.n268 10.6151
R733 B.n268 B.n267 10.6151
R734 B.n267 B.n228 10.6151
R735 B.n391 B.n228 10.6151
R736 B.n393 B.n392 10.6151
R737 B.n393 B.n219 10.6151
R738 B.n403 B.n219 10.6151
R739 B.n404 B.n403 10.6151
R740 B.n405 B.n404 10.6151
R741 B.n405 B.n212 10.6151
R742 B.n415 B.n212 10.6151
R743 B.n416 B.n415 10.6151
R744 B.n417 B.n416 10.6151
R745 B.n417 B.n204 10.6151
R746 B.n427 B.n204 10.6151
R747 B.n428 B.n427 10.6151
R748 B.n430 B.n428 10.6151
R749 B.n430 B.n429 10.6151
R750 B.n429 B.n197 10.6151
R751 B.n442 B.n197 10.6151
R752 B.n443 B.n442 10.6151
R753 B.n444 B.n443 10.6151
R754 B.n445 B.n444 10.6151
R755 B.n446 B.n445 10.6151
R756 B.n449 B.n446 10.6151
R757 B.n450 B.n449 10.6151
R758 B.n451 B.n450 10.6151
R759 B.n452 B.n451 10.6151
R760 B.n454 B.n452 10.6151
R761 B.n455 B.n454 10.6151
R762 B.n456 B.n455 10.6151
R763 B.n457 B.n456 10.6151
R764 B.n459 B.n457 10.6151
R765 B.n460 B.n459 10.6151
R766 B.n461 B.n460 10.6151
R767 B.n462 B.n461 10.6151
R768 B.n464 B.n462 10.6151
R769 B.n465 B.n464 10.6151
R770 B.n466 B.n465 10.6151
R771 B.n499 B.n1 10.6151
R772 B.n499 B.n498 10.6151
R773 B.n498 B.n497 10.6151
R774 B.n497 B.n10 10.6151
R775 B.n491 B.n10 10.6151
R776 B.n491 B.n490 10.6151
R777 B.n490 B.n489 10.6151
R778 B.n489 B.n18 10.6151
R779 B.n483 B.n18 10.6151
R780 B.n483 B.n482 10.6151
R781 B.n482 B.n481 10.6151
R782 B.n481 B.n25 10.6151
R783 B.n475 B.n25 10.6151
R784 B.n475 B.n474 10.6151
R785 B.n474 B.n473 10.6151
R786 B.n473 B.n32 10.6151
R787 B.n75 B.n74 10.6151
R788 B.n78 B.n75 10.6151
R789 B.n79 B.n78 10.6151
R790 B.n82 B.n79 10.6151
R791 B.n83 B.n82 10.6151
R792 B.n86 B.n83 10.6151
R793 B.n87 B.n86 10.6151
R794 B.n90 B.n87 10.6151
R795 B.n91 B.n90 10.6151
R796 B.n94 B.n91 10.6151
R797 B.n95 B.n94 10.6151
R798 B.n98 B.n95 10.6151
R799 B.n99 B.n98 10.6151
R800 B.n102 B.n99 10.6151
R801 B.n103 B.n102 10.6151
R802 B.n106 B.n103 10.6151
R803 B.n107 B.n106 10.6151
R804 B.n110 B.n107 10.6151
R805 B.n111 B.n110 10.6151
R806 B.n114 B.n111 10.6151
R807 B.n115 B.n114 10.6151
R808 B.n118 B.n115 10.6151
R809 B.n119 B.n118 10.6151
R810 B.n122 B.n119 10.6151
R811 B.n123 B.n122 10.6151
R812 B.n126 B.n123 10.6151
R813 B.n131 B.n128 10.6151
R814 B.n132 B.n131 10.6151
R815 B.n135 B.n132 10.6151
R816 B.n136 B.n135 10.6151
R817 B.n139 B.n136 10.6151
R818 B.n140 B.n139 10.6151
R819 B.n143 B.n140 10.6151
R820 B.n144 B.n143 10.6151
R821 B.n148 B.n147 10.6151
R822 B.n151 B.n148 10.6151
R823 B.n152 B.n151 10.6151
R824 B.n155 B.n152 10.6151
R825 B.n156 B.n155 10.6151
R826 B.n159 B.n156 10.6151
R827 B.n160 B.n159 10.6151
R828 B.n163 B.n160 10.6151
R829 B.n164 B.n163 10.6151
R830 B.n167 B.n164 10.6151
R831 B.n168 B.n167 10.6151
R832 B.n171 B.n168 10.6151
R833 B.n172 B.n171 10.6151
R834 B.n175 B.n172 10.6151
R835 B.n176 B.n175 10.6151
R836 B.n179 B.n176 10.6151
R837 B.n180 B.n179 10.6151
R838 B.n183 B.n180 10.6151
R839 B.n184 B.n183 10.6151
R840 B.n187 B.n184 10.6151
R841 B.n188 B.n187 10.6151
R842 B.n191 B.n188 10.6151
R843 B.n192 B.n191 10.6151
R844 B.n195 B.n192 10.6151
R845 B.n196 B.n195 10.6151
R846 B.n467 B.n196 10.6151
R847 B.n507 B.n0 8.11757
R848 B.n507 B.n1 8.11757
R849 B.n333 B.n263 6.5566
R850 B.n317 B.n316 6.5566
R851 B.n128 B.n127 6.5566
R852 B.n144 B.n70 6.5566
R853 B.n407 B.t5 6.35102
R854 B.n479 B.t9 6.35102
R855 B.n336 B.n263 4.05904
R856 B.n316 B.n315 4.05904
R857 B.n127 B.n126 4.05904
R858 B.n147 B.n70 4.05904
R859 VN.n0 VN.t2 301.284
R860 VN.n1 VN.t3 301.284
R861 VN.n0 VN.t1 301.233
R862 VN.n1 VN.t0 301.233
R863 VN VN.n1 81.664
R864 VN VN.n0 44.7132
R865 VDD2.n2 VDD2.n0 99.9014
R866 VDD2.n2 VDD2.n1 67.541
R867 VDD2.n1 VDD2.t3 2.89101
R868 VDD2.n1 VDD2.t1 2.89101
R869 VDD2.n0 VDD2.t0 2.89101
R870 VDD2.n0 VDD2.t2 2.89101
R871 VDD2 VDD2.n2 0.0586897
R872 VTAIL.n5 VTAIL.t0 53.7529
R873 VTAIL.n4 VTAIL.t4 53.7529
R874 VTAIL.n3 VTAIL.t7 53.7529
R875 VTAIL.n7 VTAIL.t6 53.7527
R876 VTAIL.n0 VTAIL.t5 53.7527
R877 VTAIL.n1 VTAIL.t1 53.7527
R878 VTAIL.n2 VTAIL.t2 53.7527
R879 VTAIL.n6 VTAIL.t3 53.7527
R880 VTAIL.n7 VTAIL.n6 19.1858
R881 VTAIL.n3 VTAIL.n2 19.1858
R882 VTAIL.n4 VTAIL.n3 0.914293
R883 VTAIL.n6 VTAIL.n5 0.914293
R884 VTAIL.n2 VTAIL.n1 0.914293
R885 VTAIL VTAIL.n0 0.515586
R886 VTAIL.n5 VTAIL.n4 0.470328
R887 VTAIL.n1 VTAIL.n0 0.470328
R888 VTAIL VTAIL.n7 0.399207
R889 VP.n1 VP.t0 301.284
R890 VP.n1 VP.t1 301.233
R891 VP.n3 VP.t2 280.286
R892 VP.n5 VP.t3 280.286
R893 VP.n6 VP.n5 161.3
R894 VP.n4 VP.n0 161.3
R895 VP.n3 VP.n2 161.3
R896 VP.n2 VP.n1 81.2833
R897 VP.n4 VP.n3 24.1005
R898 VP.n5 VP.n4 24.1005
R899 VP.n2 VP.n0 0.189894
R900 VP.n6 VP.n0 0.189894
R901 VP VP.n6 0.0516364
R902 VDD1 VDD1.n1 100.427
R903 VDD1 VDD1.n0 67.5992
R904 VDD1.n0 VDD1.t3 2.89101
R905 VDD1.n0 VDD1.t2 2.89101
R906 VDD1.n1 VDD1.t1 2.89101
R907 VDD1.n1 VDD1.t0 2.89101
C0 VDD2 VDD1 0.573313f
C1 VP VDD2 0.27512f
C2 VP VDD1 2.08917f
C3 VTAIL VN 1.82931f
C4 VN VDD2 1.96143f
C5 VN VDD1 0.147116f
C6 VP VN 3.89094f
C7 VTAIL VDD2 4.49706f
C8 VTAIL VDD1 4.45539f
C9 VP VTAIL 1.84341f
C10 VDD2 B 2.286608f
C11 VDD1 B 5.35993f
C12 VTAIL B 5.768237f
C13 VN B 6.03692f
C14 VP B 4.551667f
C15 VDD1.t3 B 0.151458f
C16 VDD1.t2 B 0.151458f
C17 VDD1.n0 B 1.29403f
C18 VDD1.t1 B 0.151458f
C19 VDD1.t0 B 0.151458f
C20 VDD1.n1 B 1.72481f
C21 VP.n0 B 0.038968f
C22 VP.t1 B 0.580534f
C23 VP.t0 B 0.580583f
C24 VP.n1 B 1.07825f
C25 VP.n2 B 2.04466f
C26 VP.t2 B 0.563092f
C27 VP.n3 B 0.248026f
C28 VP.n4 B 0.008843f
C29 VP.t3 B 0.563092f
C30 VP.n5 B 0.248026f
C31 VP.n6 B 0.030199f
C32 VTAIL.t5 B 0.703929f
C33 VTAIL.n0 B 0.189505f
C34 VTAIL.t1 B 0.703929f
C35 VTAIL.n1 B 0.205757f
C36 VTAIL.t2 B 0.703929f
C37 VTAIL.n2 B 0.636385f
C38 VTAIL.t7 B 0.703935f
C39 VTAIL.n3 B 0.636379f
C40 VTAIL.t4 B 0.703935f
C41 VTAIL.n4 B 0.205751f
C42 VTAIL.t0 B 0.703935f
C43 VTAIL.n5 B 0.205751f
C44 VTAIL.t3 B 0.703929f
C45 VTAIL.n6 B 0.636385f
C46 VTAIL.t6 B 0.703929f
C47 VTAIL.n7 B 0.61539f
C48 VDD2.t0 B 0.10491f
C49 VDD2.t2 B 0.10491f
C50 VDD2.n0 B 1.17862f
C51 VDD2.t3 B 0.10491f
C52 VDD2.t1 B 0.10491f
C53 VDD2.n1 B 0.89614f
C54 VDD2.n2 B 1.94437f
C55 VN.t2 B 0.373965f
C56 VN.t1 B 0.373933f
C57 VN.n0 B 0.302968f
C58 VN.t3 B 0.373965f
C59 VN.t0 B 0.373933f
C60 VN.n1 B 0.70428f
.ends

