* NGSPICE file created from diff_pair_sample_0054.ext - technology: sky130A

.subckt diff_pair_sample_0054 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=1.38
X1 VTAIL.t14 VN.t1 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=1.38
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=1.38
X4 VTAIL.t18 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X5 VTAIL.t15 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X6 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=1.38
X7 VTAIL.t3 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X8 VDD1.t8 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=1.38
X9 VDD1.t7 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=1.38
X10 VDD1.t6 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X11 VTAIL.t11 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X12 VTAIL.t6 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X13 VDD2.t4 VN.t5 VTAIL.t9 B.t22 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=1.38
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0 ps=0 w=2.49 l=1.38
X15 VDD2.t3 VN.t6 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=1.38
X16 VDD2.t2 VN.t7 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X17 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X18 VTAIL.t1 VP.t6 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X19 VTAIL.t0 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X20 VDD2.t1 VN.t8 VTAIL.t10 B.t23 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=1.38
X21 VDD2.t0 VN.t9 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.41085 ps=2.82 w=2.49 l=1.38
X22 VDD1.t1 VP.t8 VTAIL.t8 B.t22 sky130_fd_pr__nfet_01v8 ad=0.41085 pd=2.82 as=0.9711 ps=5.76 w=2.49 l=1.38
X23 VDD1.t0 VP.t9 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=0.9711 pd=5.76 as=0.41085 ps=2.82 w=2.49 l=1.38
R0 VN.n25 VN.n24 177.448
R1 VN.n51 VN.n50 177.448
R2 VN.n49 VN.n26 161.3
R3 VN.n48 VN.n47 161.3
R4 VN.n46 VN.n27 161.3
R5 VN.n45 VN.n44 161.3
R6 VN.n42 VN.n28 161.3
R7 VN.n41 VN.n40 161.3
R8 VN.n39 VN.n29 161.3
R9 VN.n38 VN.n37 161.3
R10 VN.n36 VN.n30 161.3
R11 VN.n35 VN.n34 161.3
R12 VN.n23 VN.n0 161.3
R13 VN.n22 VN.n21 161.3
R14 VN.n20 VN.n1 161.3
R15 VN.n19 VN.n18 161.3
R16 VN.n16 VN.n2 161.3
R17 VN.n15 VN.n14 161.3
R18 VN.n13 VN.n3 161.3
R19 VN.n12 VN.n11 161.3
R20 VN.n9 VN.n4 161.3
R21 VN.n8 VN.n7 161.3
R22 VN.n6 VN.t6 76.3298
R23 VN.n33 VN.t5 76.3298
R24 VN.n22 VN.n1 56.5193
R25 VN.n48 VN.n27 56.5193
R26 VN.n9 VN.n8 50.6917
R27 VN.n16 VN.n15 50.6917
R28 VN.n36 VN.n35 50.6917
R29 VN.n42 VN.n41 50.6917
R30 VN.n6 VN.n5 43.6963
R31 VN.n33 VN.n32 43.6963
R32 VN.n5 VN.t3 43.4853
R33 VN.n10 VN.t9 43.4853
R34 VN.n17 VN.t4 43.4853
R35 VN.n24 VN.t0 43.4853
R36 VN.n32 VN.t1 43.4853
R37 VN.n31 VN.t7 43.4853
R38 VN.n43 VN.t2 43.4853
R39 VN.n50 VN.t8 43.4853
R40 VN VN.n51 39.5289
R41 VN.n11 VN.n9 30.2951
R42 VN.n15 VN.n3 30.2951
R43 VN.n37 VN.n36 30.2951
R44 VN.n41 VN.n29 30.2951
R45 VN.n18 VN.n1 24.4675
R46 VN.n23 VN.n22 24.4675
R47 VN.n44 VN.n27 24.4675
R48 VN.n49 VN.n48 24.4675
R49 VN.n8 VN.n5 22.5101
R50 VN.n17 VN.n16 22.5101
R51 VN.n35 VN.n32 22.5101
R52 VN.n43 VN.n42 22.5101
R53 VN.n34 VN.n33 17.9509
R54 VN.n7 VN.n6 17.9509
R55 VN.n11 VN.n10 12.234
R56 VN.n10 VN.n3 12.234
R57 VN.n31 VN.n29 12.234
R58 VN.n37 VN.n31 12.234
R59 VN.n24 VN.n23 8.31928
R60 VN.n50 VN.n49 8.31928
R61 VN.n18 VN.n17 1.95786
R62 VN.n44 VN.n43 1.95786
R63 VN.n51 VN.n26 0.189894
R64 VN.n47 VN.n26 0.189894
R65 VN.n47 VN.n46 0.189894
R66 VN.n46 VN.n45 0.189894
R67 VN.n45 VN.n28 0.189894
R68 VN.n40 VN.n28 0.189894
R69 VN.n40 VN.n39 0.189894
R70 VN.n39 VN.n38 0.189894
R71 VN.n38 VN.n30 0.189894
R72 VN.n34 VN.n30 0.189894
R73 VN.n7 VN.n4 0.189894
R74 VN.n12 VN.n4 0.189894
R75 VN.n13 VN.n12 0.189894
R76 VN.n14 VN.n13 0.189894
R77 VN.n14 VN.n2 0.189894
R78 VN.n19 VN.n2 0.189894
R79 VN.n20 VN.n19 0.189894
R80 VN.n21 VN.n20 0.189894
R81 VN.n21 VN.n0 0.189894
R82 VN.n25 VN.n0 0.189894
R83 VN VN.n25 0.0516364
R84 VTAIL.n56 VTAIL.n50 289.615
R85 VTAIL.n8 VTAIL.n2 289.615
R86 VTAIL.n44 VTAIL.n38 289.615
R87 VTAIL.n28 VTAIL.n22 289.615
R88 VTAIL.n55 VTAIL.n54 185
R89 VTAIL.n57 VTAIL.n56 185
R90 VTAIL.n7 VTAIL.n6 185
R91 VTAIL.n9 VTAIL.n8 185
R92 VTAIL.n45 VTAIL.n44 185
R93 VTAIL.n43 VTAIL.n42 185
R94 VTAIL.n29 VTAIL.n28 185
R95 VTAIL.n27 VTAIL.n26 185
R96 VTAIL.n53 VTAIL.t13 151.613
R97 VTAIL.n5 VTAIL.t8 151.613
R98 VTAIL.n41 VTAIL.t7 151.613
R99 VTAIL.n25 VTAIL.t9 151.613
R100 VTAIL.n56 VTAIL.n55 104.615
R101 VTAIL.n8 VTAIL.n7 104.615
R102 VTAIL.n44 VTAIL.n43 104.615
R103 VTAIL.n28 VTAIL.n27 104.615
R104 VTAIL.n37 VTAIL.n36 70.0259
R105 VTAIL.n35 VTAIL.n34 70.0259
R106 VTAIL.n21 VTAIL.n20 70.0259
R107 VTAIL.n19 VTAIL.n18 70.0259
R108 VTAIL.n63 VTAIL.n62 70.0259
R109 VTAIL.n1 VTAIL.n0 70.0259
R110 VTAIL.n15 VTAIL.n14 70.0259
R111 VTAIL.n17 VTAIL.n16 70.0259
R112 VTAIL.n55 VTAIL.t13 52.3082
R113 VTAIL.n7 VTAIL.t8 52.3082
R114 VTAIL.n43 VTAIL.t7 52.3082
R115 VTAIL.n27 VTAIL.t9 52.3082
R116 VTAIL.n61 VTAIL.n60 33.9308
R117 VTAIL.n13 VTAIL.n12 33.9308
R118 VTAIL.n49 VTAIL.n48 33.9308
R119 VTAIL.n33 VTAIL.n32 33.9308
R120 VTAIL.n19 VTAIL.n17 17.4617
R121 VTAIL.n61 VTAIL.n49 15.9876
R122 VTAIL.n54 VTAIL.n53 15.3979
R123 VTAIL.n6 VTAIL.n5 15.3979
R124 VTAIL.n42 VTAIL.n41 15.3979
R125 VTAIL.n26 VTAIL.n25 15.3979
R126 VTAIL.n57 VTAIL.n52 12.8005
R127 VTAIL.n9 VTAIL.n4 12.8005
R128 VTAIL.n45 VTAIL.n40 12.8005
R129 VTAIL.n29 VTAIL.n24 12.8005
R130 VTAIL.n58 VTAIL.n50 12.0247
R131 VTAIL.n10 VTAIL.n2 12.0247
R132 VTAIL.n46 VTAIL.n38 12.0247
R133 VTAIL.n30 VTAIL.n22 12.0247
R134 VTAIL.n60 VTAIL.n59 9.45567
R135 VTAIL.n12 VTAIL.n11 9.45567
R136 VTAIL.n48 VTAIL.n47 9.45567
R137 VTAIL.n32 VTAIL.n31 9.45567
R138 VTAIL.n59 VTAIL.n58 9.3005
R139 VTAIL.n52 VTAIL.n51 9.3005
R140 VTAIL.n11 VTAIL.n10 9.3005
R141 VTAIL.n4 VTAIL.n3 9.3005
R142 VTAIL.n47 VTAIL.n46 9.3005
R143 VTAIL.n40 VTAIL.n39 9.3005
R144 VTAIL.n31 VTAIL.n30 9.3005
R145 VTAIL.n24 VTAIL.n23 9.3005
R146 VTAIL.n62 VTAIL.t17 7.95231
R147 VTAIL.n62 VTAIL.t11 7.95231
R148 VTAIL.n0 VTAIL.t12 7.95231
R149 VTAIL.n0 VTAIL.t15 7.95231
R150 VTAIL.n14 VTAIL.t2 7.95231
R151 VTAIL.n14 VTAIL.t6 7.95231
R152 VTAIL.n16 VTAIL.t19 7.95231
R153 VTAIL.n16 VTAIL.t3 7.95231
R154 VTAIL.n36 VTAIL.t4 7.95231
R155 VTAIL.n36 VTAIL.t0 7.95231
R156 VTAIL.n34 VTAIL.t5 7.95231
R157 VTAIL.n34 VTAIL.t1 7.95231
R158 VTAIL.n20 VTAIL.t16 7.95231
R159 VTAIL.n20 VTAIL.t14 7.95231
R160 VTAIL.n18 VTAIL.t10 7.95231
R161 VTAIL.n18 VTAIL.t18 7.95231
R162 VTAIL.n53 VTAIL.n51 4.69785
R163 VTAIL.n5 VTAIL.n3 4.69785
R164 VTAIL.n41 VTAIL.n39 4.69785
R165 VTAIL.n25 VTAIL.n23 4.69785
R166 VTAIL.n60 VTAIL.n50 1.93989
R167 VTAIL.n12 VTAIL.n2 1.93989
R168 VTAIL.n48 VTAIL.n38 1.93989
R169 VTAIL.n32 VTAIL.n22 1.93989
R170 VTAIL.n21 VTAIL.n19 1.47464
R171 VTAIL.n33 VTAIL.n21 1.47464
R172 VTAIL.n37 VTAIL.n35 1.47464
R173 VTAIL.n49 VTAIL.n37 1.47464
R174 VTAIL.n17 VTAIL.n15 1.47464
R175 VTAIL.n15 VTAIL.n13 1.47464
R176 VTAIL.n63 VTAIL.n61 1.47464
R177 VTAIL.n35 VTAIL.n33 1.2074
R178 VTAIL.n13 VTAIL.n1 1.2074
R179 VTAIL VTAIL.n1 1.16429
R180 VTAIL.n58 VTAIL.n57 1.16414
R181 VTAIL.n10 VTAIL.n9 1.16414
R182 VTAIL.n46 VTAIL.n45 1.16414
R183 VTAIL.n30 VTAIL.n29 1.16414
R184 VTAIL.n54 VTAIL.n52 0.388379
R185 VTAIL.n6 VTAIL.n4 0.388379
R186 VTAIL.n42 VTAIL.n40 0.388379
R187 VTAIL.n26 VTAIL.n24 0.388379
R188 VTAIL VTAIL.n63 0.310845
R189 VTAIL.n59 VTAIL.n51 0.155672
R190 VTAIL.n11 VTAIL.n3 0.155672
R191 VTAIL.n47 VTAIL.n39 0.155672
R192 VTAIL.n31 VTAIL.n23 0.155672
R193 VDD2.n21 VDD2.n15 289.615
R194 VDD2.n6 VDD2.n0 289.615
R195 VDD2.n22 VDD2.n21 185
R196 VDD2.n20 VDD2.n19 185
R197 VDD2.n5 VDD2.n4 185
R198 VDD2.n7 VDD2.n6 185
R199 VDD2.n18 VDD2.t1 151.613
R200 VDD2.n3 VDD2.t3 151.613
R201 VDD2.n21 VDD2.n20 104.615
R202 VDD2.n6 VDD2.n5 104.615
R203 VDD2.n14 VDD2.n13 87.7549
R204 VDD2 VDD2.n29 87.752
R205 VDD2.n28 VDD2.n27 86.7047
R206 VDD2.n12 VDD2.n11 86.7046
R207 VDD2.n20 VDD2.t1 52.3082
R208 VDD2.n5 VDD2.t3 52.3082
R209 VDD2.n12 VDD2.n10 52.0837
R210 VDD2.n26 VDD2.n25 50.6096
R211 VDD2.n26 VDD2.n14 32.864
R212 VDD2.n19 VDD2.n18 15.3979
R213 VDD2.n4 VDD2.n3 15.3979
R214 VDD2.n22 VDD2.n17 12.8005
R215 VDD2.n7 VDD2.n2 12.8005
R216 VDD2.n23 VDD2.n15 12.0247
R217 VDD2.n8 VDD2.n0 12.0247
R218 VDD2.n25 VDD2.n24 9.45567
R219 VDD2.n10 VDD2.n9 9.45567
R220 VDD2.n24 VDD2.n23 9.3005
R221 VDD2.n17 VDD2.n16 9.3005
R222 VDD2.n9 VDD2.n8 9.3005
R223 VDD2.n2 VDD2.n1 9.3005
R224 VDD2.n29 VDD2.t8 7.95231
R225 VDD2.n29 VDD2.t4 7.95231
R226 VDD2.n27 VDD2.t7 7.95231
R227 VDD2.n27 VDD2.t2 7.95231
R228 VDD2.n13 VDD2.t5 7.95231
R229 VDD2.n13 VDD2.t9 7.95231
R230 VDD2.n11 VDD2.t6 7.95231
R231 VDD2.n11 VDD2.t0 7.95231
R232 VDD2.n18 VDD2.n16 4.69785
R233 VDD2.n3 VDD2.n1 4.69785
R234 VDD2.n25 VDD2.n15 1.93989
R235 VDD2.n10 VDD2.n0 1.93989
R236 VDD2.n28 VDD2.n26 1.47464
R237 VDD2.n23 VDD2.n22 1.16414
R238 VDD2.n8 VDD2.n7 1.16414
R239 VDD2 VDD2.n28 0.427224
R240 VDD2.n19 VDD2.n17 0.388379
R241 VDD2.n4 VDD2.n2 0.388379
R242 VDD2.n14 VDD2.n12 0.313688
R243 VDD2.n24 VDD2.n16 0.155672
R244 VDD2.n9 VDD2.n1 0.155672
R245 B.n430 B.n429 585
R246 B.n430 B.n71 585
R247 B.n433 B.n432 585
R248 B.n434 B.n94 585
R249 B.n436 B.n435 585
R250 B.n438 B.n93 585
R251 B.n441 B.n440 585
R252 B.n442 B.n92 585
R253 B.n444 B.n443 585
R254 B.n446 B.n91 585
R255 B.n449 B.n448 585
R256 B.n450 B.n90 585
R257 B.n452 B.n451 585
R258 B.n454 B.n89 585
R259 B.n457 B.n456 585
R260 B.n459 B.n86 585
R261 B.n461 B.n460 585
R262 B.n463 B.n85 585
R263 B.n466 B.n465 585
R264 B.n467 B.n84 585
R265 B.n469 B.n468 585
R266 B.n471 B.n83 585
R267 B.n473 B.n472 585
R268 B.n475 B.n474 585
R269 B.n478 B.n477 585
R270 B.n479 B.n78 585
R271 B.n481 B.n480 585
R272 B.n483 B.n77 585
R273 B.n486 B.n485 585
R274 B.n487 B.n76 585
R275 B.n489 B.n488 585
R276 B.n491 B.n75 585
R277 B.n494 B.n493 585
R278 B.n495 B.n74 585
R279 B.n497 B.n496 585
R280 B.n499 B.n73 585
R281 B.n502 B.n501 585
R282 B.n503 B.n72 585
R283 B.n428 B.n70 585
R284 B.n506 B.n70 585
R285 B.n427 B.n69 585
R286 B.n507 B.n69 585
R287 B.n426 B.n68 585
R288 B.n508 B.n68 585
R289 B.n425 B.n424 585
R290 B.n424 B.n64 585
R291 B.n423 B.n63 585
R292 B.n514 B.n63 585
R293 B.n422 B.n62 585
R294 B.n515 B.n62 585
R295 B.n421 B.n61 585
R296 B.n516 B.n61 585
R297 B.n420 B.n419 585
R298 B.n419 B.n57 585
R299 B.n418 B.n56 585
R300 B.n522 B.n56 585
R301 B.n417 B.n55 585
R302 B.n523 B.n55 585
R303 B.n416 B.n54 585
R304 B.n524 B.n54 585
R305 B.n415 B.n414 585
R306 B.n414 B.n50 585
R307 B.n413 B.n49 585
R308 B.n530 B.n49 585
R309 B.n412 B.n48 585
R310 B.n531 B.n48 585
R311 B.n411 B.n47 585
R312 B.n532 B.n47 585
R313 B.n410 B.n409 585
R314 B.n409 B.n43 585
R315 B.n408 B.n42 585
R316 B.n538 B.n42 585
R317 B.n407 B.n41 585
R318 B.n539 B.n41 585
R319 B.n406 B.n40 585
R320 B.n540 B.n40 585
R321 B.n405 B.n404 585
R322 B.n404 B.n36 585
R323 B.n403 B.n35 585
R324 B.n546 B.n35 585
R325 B.n402 B.n34 585
R326 B.n547 B.n34 585
R327 B.n401 B.n33 585
R328 B.n548 B.n33 585
R329 B.n400 B.n399 585
R330 B.n399 B.n32 585
R331 B.n398 B.n28 585
R332 B.n554 B.n28 585
R333 B.n397 B.n27 585
R334 B.n555 B.n27 585
R335 B.n396 B.n26 585
R336 B.n556 B.n26 585
R337 B.n395 B.n394 585
R338 B.n394 B.n22 585
R339 B.n393 B.n21 585
R340 B.n562 B.n21 585
R341 B.n392 B.n20 585
R342 B.n563 B.n20 585
R343 B.n391 B.n19 585
R344 B.n564 B.n19 585
R345 B.n390 B.n389 585
R346 B.n389 B.n15 585
R347 B.n388 B.n14 585
R348 B.n570 B.n14 585
R349 B.n387 B.n13 585
R350 B.n571 B.n13 585
R351 B.n386 B.n12 585
R352 B.n572 B.n12 585
R353 B.n385 B.n384 585
R354 B.n384 B.n8 585
R355 B.n383 B.n7 585
R356 B.n578 B.n7 585
R357 B.n382 B.n6 585
R358 B.n579 B.n6 585
R359 B.n381 B.n5 585
R360 B.n580 B.n5 585
R361 B.n380 B.n379 585
R362 B.n379 B.n4 585
R363 B.n378 B.n95 585
R364 B.n378 B.n377 585
R365 B.n368 B.n96 585
R366 B.n97 B.n96 585
R367 B.n370 B.n369 585
R368 B.n371 B.n370 585
R369 B.n367 B.n101 585
R370 B.n105 B.n101 585
R371 B.n366 B.n365 585
R372 B.n365 B.n364 585
R373 B.n103 B.n102 585
R374 B.n104 B.n103 585
R375 B.n357 B.n356 585
R376 B.n358 B.n357 585
R377 B.n355 B.n110 585
R378 B.n110 B.n109 585
R379 B.n354 B.n353 585
R380 B.n353 B.n352 585
R381 B.n112 B.n111 585
R382 B.n113 B.n112 585
R383 B.n345 B.n344 585
R384 B.n346 B.n345 585
R385 B.n343 B.n118 585
R386 B.n118 B.n117 585
R387 B.n342 B.n341 585
R388 B.n341 B.n340 585
R389 B.n120 B.n119 585
R390 B.n333 B.n120 585
R391 B.n332 B.n331 585
R392 B.n334 B.n332 585
R393 B.n330 B.n125 585
R394 B.n125 B.n124 585
R395 B.n329 B.n328 585
R396 B.n328 B.n327 585
R397 B.n127 B.n126 585
R398 B.n128 B.n127 585
R399 B.n320 B.n319 585
R400 B.n321 B.n320 585
R401 B.n318 B.n133 585
R402 B.n133 B.n132 585
R403 B.n317 B.n316 585
R404 B.n316 B.n315 585
R405 B.n135 B.n134 585
R406 B.n136 B.n135 585
R407 B.n308 B.n307 585
R408 B.n309 B.n308 585
R409 B.n306 B.n140 585
R410 B.n144 B.n140 585
R411 B.n305 B.n304 585
R412 B.n304 B.n303 585
R413 B.n142 B.n141 585
R414 B.n143 B.n142 585
R415 B.n296 B.n295 585
R416 B.n297 B.n296 585
R417 B.n294 B.n149 585
R418 B.n149 B.n148 585
R419 B.n293 B.n292 585
R420 B.n292 B.n291 585
R421 B.n151 B.n150 585
R422 B.n152 B.n151 585
R423 B.n284 B.n283 585
R424 B.n285 B.n284 585
R425 B.n282 B.n156 585
R426 B.n160 B.n156 585
R427 B.n281 B.n280 585
R428 B.n280 B.n279 585
R429 B.n158 B.n157 585
R430 B.n159 B.n158 585
R431 B.n272 B.n271 585
R432 B.n273 B.n272 585
R433 B.n270 B.n165 585
R434 B.n165 B.n164 585
R435 B.n269 B.n268 585
R436 B.n268 B.n267 585
R437 B.n264 B.n169 585
R438 B.n263 B.n262 585
R439 B.n260 B.n170 585
R440 B.n260 B.n168 585
R441 B.n259 B.n258 585
R442 B.n257 B.n256 585
R443 B.n255 B.n172 585
R444 B.n253 B.n252 585
R445 B.n251 B.n173 585
R446 B.n250 B.n249 585
R447 B.n247 B.n174 585
R448 B.n245 B.n244 585
R449 B.n243 B.n175 585
R450 B.n242 B.n241 585
R451 B.n239 B.n176 585
R452 B.n237 B.n236 585
R453 B.n235 B.n177 585
R454 B.n234 B.n233 585
R455 B.n231 B.n181 585
R456 B.n229 B.n228 585
R457 B.n227 B.n182 585
R458 B.n226 B.n225 585
R459 B.n223 B.n183 585
R460 B.n221 B.n220 585
R461 B.n218 B.n184 585
R462 B.n217 B.n216 585
R463 B.n214 B.n187 585
R464 B.n212 B.n211 585
R465 B.n210 B.n188 585
R466 B.n209 B.n208 585
R467 B.n206 B.n189 585
R468 B.n204 B.n203 585
R469 B.n202 B.n190 585
R470 B.n201 B.n200 585
R471 B.n198 B.n191 585
R472 B.n196 B.n195 585
R473 B.n194 B.n193 585
R474 B.n167 B.n166 585
R475 B.n266 B.n265 585
R476 B.n267 B.n266 585
R477 B.n163 B.n162 585
R478 B.n164 B.n163 585
R479 B.n275 B.n274 585
R480 B.n274 B.n273 585
R481 B.n276 B.n161 585
R482 B.n161 B.n159 585
R483 B.n278 B.n277 585
R484 B.n279 B.n278 585
R485 B.n155 B.n154 585
R486 B.n160 B.n155 585
R487 B.n287 B.n286 585
R488 B.n286 B.n285 585
R489 B.n288 B.n153 585
R490 B.n153 B.n152 585
R491 B.n290 B.n289 585
R492 B.n291 B.n290 585
R493 B.n147 B.n146 585
R494 B.n148 B.n147 585
R495 B.n299 B.n298 585
R496 B.n298 B.n297 585
R497 B.n300 B.n145 585
R498 B.n145 B.n143 585
R499 B.n302 B.n301 585
R500 B.n303 B.n302 585
R501 B.n139 B.n138 585
R502 B.n144 B.n139 585
R503 B.n311 B.n310 585
R504 B.n310 B.n309 585
R505 B.n312 B.n137 585
R506 B.n137 B.n136 585
R507 B.n314 B.n313 585
R508 B.n315 B.n314 585
R509 B.n131 B.n130 585
R510 B.n132 B.n131 585
R511 B.n323 B.n322 585
R512 B.n322 B.n321 585
R513 B.n324 B.n129 585
R514 B.n129 B.n128 585
R515 B.n326 B.n325 585
R516 B.n327 B.n326 585
R517 B.n123 B.n122 585
R518 B.n124 B.n123 585
R519 B.n336 B.n335 585
R520 B.n335 B.n334 585
R521 B.n337 B.n121 585
R522 B.n333 B.n121 585
R523 B.n339 B.n338 585
R524 B.n340 B.n339 585
R525 B.n116 B.n115 585
R526 B.n117 B.n116 585
R527 B.n348 B.n347 585
R528 B.n347 B.n346 585
R529 B.n349 B.n114 585
R530 B.n114 B.n113 585
R531 B.n351 B.n350 585
R532 B.n352 B.n351 585
R533 B.n108 B.n107 585
R534 B.n109 B.n108 585
R535 B.n360 B.n359 585
R536 B.n359 B.n358 585
R537 B.n361 B.n106 585
R538 B.n106 B.n104 585
R539 B.n363 B.n362 585
R540 B.n364 B.n363 585
R541 B.n100 B.n99 585
R542 B.n105 B.n100 585
R543 B.n373 B.n372 585
R544 B.n372 B.n371 585
R545 B.n374 B.n98 585
R546 B.n98 B.n97 585
R547 B.n376 B.n375 585
R548 B.n377 B.n376 585
R549 B.n2 B.n0 585
R550 B.n4 B.n2 585
R551 B.n3 B.n1 585
R552 B.n579 B.n3 585
R553 B.n577 B.n576 585
R554 B.n578 B.n577 585
R555 B.n575 B.n9 585
R556 B.n9 B.n8 585
R557 B.n574 B.n573 585
R558 B.n573 B.n572 585
R559 B.n11 B.n10 585
R560 B.n571 B.n11 585
R561 B.n569 B.n568 585
R562 B.n570 B.n569 585
R563 B.n567 B.n16 585
R564 B.n16 B.n15 585
R565 B.n566 B.n565 585
R566 B.n565 B.n564 585
R567 B.n18 B.n17 585
R568 B.n563 B.n18 585
R569 B.n561 B.n560 585
R570 B.n562 B.n561 585
R571 B.n559 B.n23 585
R572 B.n23 B.n22 585
R573 B.n558 B.n557 585
R574 B.n557 B.n556 585
R575 B.n25 B.n24 585
R576 B.n555 B.n25 585
R577 B.n553 B.n552 585
R578 B.n554 B.n553 585
R579 B.n551 B.n29 585
R580 B.n32 B.n29 585
R581 B.n550 B.n549 585
R582 B.n549 B.n548 585
R583 B.n31 B.n30 585
R584 B.n547 B.n31 585
R585 B.n545 B.n544 585
R586 B.n546 B.n545 585
R587 B.n543 B.n37 585
R588 B.n37 B.n36 585
R589 B.n542 B.n541 585
R590 B.n541 B.n540 585
R591 B.n39 B.n38 585
R592 B.n539 B.n39 585
R593 B.n537 B.n536 585
R594 B.n538 B.n537 585
R595 B.n535 B.n44 585
R596 B.n44 B.n43 585
R597 B.n534 B.n533 585
R598 B.n533 B.n532 585
R599 B.n46 B.n45 585
R600 B.n531 B.n46 585
R601 B.n529 B.n528 585
R602 B.n530 B.n529 585
R603 B.n527 B.n51 585
R604 B.n51 B.n50 585
R605 B.n526 B.n525 585
R606 B.n525 B.n524 585
R607 B.n53 B.n52 585
R608 B.n523 B.n53 585
R609 B.n521 B.n520 585
R610 B.n522 B.n521 585
R611 B.n519 B.n58 585
R612 B.n58 B.n57 585
R613 B.n518 B.n517 585
R614 B.n517 B.n516 585
R615 B.n60 B.n59 585
R616 B.n515 B.n60 585
R617 B.n513 B.n512 585
R618 B.n514 B.n513 585
R619 B.n511 B.n65 585
R620 B.n65 B.n64 585
R621 B.n510 B.n509 585
R622 B.n509 B.n508 585
R623 B.n67 B.n66 585
R624 B.n507 B.n67 585
R625 B.n505 B.n504 585
R626 B.n506 B.n505 585
R627 B.n582 B.n581 585
R628 B.n581 B.n580 585
R629 B.n266 B.n169 535.745
R630 B.n505 B.n72 535.745
R631 B.n268 B.n167 535.745
R632 B.n430 B.n70 535.745
R633 B.n431 B.n71 256.663
R634 B.n437 B.n71 256.663
R635 B.n439 B.n71 256.663
R636 B.n445 B.n71 256.663
R637 B.n447 B.n71 256.663
R638 B.n453 B.n71 256.663
R639 B.n455 B.n71 256.663
R640 B.n462 B.n71 256.663
R641 B.n464 B.n71 256.663
R642 B.n470 B.n71 256.663
R643 B.n82 B.n71 256.663
R644 B.n476 B.n71 256.663
R645 B.n482 B.n71 256.663
R646 B.n484 B.n71 256.663
R647 B.n490 B.n71 256.663
R648 B.n492 B.n71 256.663
R649 B.n498 B.n71 256.663
R650 B.n500 B.n71 256.663
R651 B.n261 B.n168 256.663
R652 B.n171 B.n168 256.663
R653 B.n254 B.n168 256.663
R654 B.n248 B.n168 256.663
R655 B.n246 B.n168 256.663
R656 B.n240 B.n168 256.663
R657 B.n238 B.n168 256.663
R658 B.n232 B.n168 256.663
R659 B.n230 B.n168 256.663
R660 B.n224 B.n168 256.663
R661 B.n222 B.n168 256.663
R662 B.n215 B.n168 256.663
R663 B.n213 B.n168 256.663
R664 B.n207 B.n168 256.663
R665 B.n205 B.n168 256.663
R666 B.n199 B.n168 256.663
R667 B.n197 B.n168 256.663
R668 B.n192 B.n168 256.663
R669 B.n185 B.t16 248.448
R670 B.n178 B.t8 248.448
R671 B.n79 B.t12 248.448
R672 B.n87 B.t19 248.448
R673 B.n267 B.n168 202.577
R674 B.n506 B.n71 202.577
R675 B.n266 B.n163 163.367
R676 B.n274 B.n163 163.367
R677 B.n274 B.n161 163.367
R678 B.n278 B.n161 163.367
R679 B.n278 B.n155 163.367
R680 B.n286 B.n155 163.367
R681 B.n286 B.n153 163.367
R682 B.n290 B.n153 163.367
R683 B.n290 B.n147 163.367
R684 B.n298 B.n147 163.367
R685 B.n298 B.n145 163.367
R686 B.n302 B.n145 163.367
R687 B.n302 B.n139 163.367
R688 B.n310 B.n139 163.367
R689 B.n310 B.n137 163.367
R690 B.n314 B.n137 163.367
R691 B.n314 B.n131 163.367
R692 B.n322 B.n131 163.367
R693 B.n322 B.n129 163.367
R694 B.n326 B.n129 163.367
R695 B.n326 B.n123 163.367
R696 B.n335 B.n123 163.367
R697 B.n335 B.n121 163.367
R698 B.n339 B.n121 163.367
R699 B.n339 B.n116 163.367
R700 B.n347 B.n116 163.367
R701 B.n347 B.n114 163.367
R702 B.n351 B.n114 163.367
R703 B.n351 B.n108 163.367
R704 B.n359 B.n108 163.367
R705 B.n359 B.n106 163.367
R706 B.n363 B.n106 163.367
R707 B.n363 B.n100 163.367
R708 B.n372 B.n100 163.367
R709 B.n372 B.n98 163.367
R710 B.n376 B.n98 163.367
R711 B.n376 B.n2 163.367
R712 B.n581 B.n2 163.367
R713 B.n581 B.n3 163.367
R714 B.n577 B.n3 163.367
R715 B.n577 B.n9 163.367
R716 B.n573 B.n9 163.367
R717 B.n573 B.n11 163.367
R718 B.n569 B.n11 163.367
R719 B.n569 B.n16 163.367
R720 B.n565 B.n16 163.367
R721 B.n565 B.n18 163.367
R722 B.n561 B.n18 163.367
R723 B.n561 B.n23 163.367
R724 B.n557 B.n23 163.367
R725 B.n557 B.n25 163.367
R726 B.n553 B.n25 163.367
R727 B.n553 B.n29 163.367
R728 B.n549 B.n29 163.367
R729 B.n549 B.n31 163.367
R730 B.n545 B.n31 163.367
R731 B.n545 B.n37 163.367
R732 B.n541 B.n37 163.367
R733 B.n541 B.n39 163.367
R734 B.n537 B.n39 163.367
R735 B.n537 B.n44 163.367
R736 B.n533 B.n44 163.367
R737 B.n533 B.n46 163.367
R738 B.n529 B.n46 163.367
R739 B.n529 B.n51 163.367
R740 B.n525 B.n51 163.367
R741 B.n525 B.n53 163.367
R742 B.n521 B.n53 163.367
R743 B.n521 B.n58 163.367
R744 B.n517 B.n58 163.367
R745 B.n517 B.n60 163.367
R746 B.n513 B.n60 163.367
R747 B.n513 B.n65 163.367
R748 B.n509 B.n65 163.367
R749 B.n509 B.n67 163.367
R750 B.n505 B.n67 163.367
R751 B.n262 B.n260 163.367
R752 B.n260 B.n259 163.367
R753 B.n256 B.n255 163.367
R754 B.n253 B.n173 163.367
R755 B.n249 B.n247 163.367
R756 B.n245 B.n175 163.367
R757 B.n241 B.n239 163.367
R758 B.n237 B.n177 163.367
R759 B.n233 B.n231 163.367
R760 B.n229 B.n182 163.367
R761 B.n225 B.n223 163.367
R762 B.n221 B.n184 163.367
R763 B.n216 B.n214 163.367
R764 B.n212 B.n188 163.367
R765 B.n208 B.n206 163.367
R766 B.n204 B.n190 163.367
R767 B.n200 B.n198 163.367
R768 B.n196 B.n193 163.367
R769 B.n268 B.n165 163.367
R770 B.n272 B.n165 163.367
R771 B.n272 B.n158 163.367
R772 B.n280 B.n158 163.367
R773 B.n280 B.n156 163.367
R774 B.n284 B.n156 163.367
R775 B.n284 B.n151 163.367
R776 B.n292 B.n151 163.367
R777 B.n292 B.n149 163.367
R778 B.n296 B.n149 163.367
R779 B.n296 B.n142 163.367
R780 B.n304 B.n142 163.367
R781 B.n304 B.n140 163.367
R782 B.n308 B.n140 163.367
R783 B.n308 B.n135 163.367
R784 B.n316 B.n135 163.367
R785 B.n316 B.n133 163.367
R786 B.n320 B.n133 163.367
R787 B.n320 B.n127 163.367
R788 B.n328 B.n127 163.367
R789 B.n328 B.n125 163.367
R790 B.n332 B.n125 163.367
R791 B.n332 B.n120 163.367
R792 B.n341 B.n120 163.367
R793 B.n341 B.n118 163.367
R794 B.n345 B.n118 163.367
R795 B.n345 B.n112 163.367
R796 B.n353 B.n112 163.367
R797 B.n353 B.n110 163.367
R798 B.n357 B.n110 163.367
R799 B.n357 B.n103 163.367
R800 B.n365 B.n103 163.367
R801 B.n365 B.n101 163.367
R802 B.n370 B.n101 163.367
R803 B.n370 B.n96 163.367
R804 B.n378 B.n96 163.367
R805 B.n379 B.n378 163.367
R806 B.n379 B.n5 163.367
R807 B.n6 B.n5 163.367
R808 B.n7 B.n6 163.367
R809 B.n384 B.n7 163.367
R810 B.n384 B.n12 163.367
R811 B.n13 B.n12 163.367
R812 B.n14 B.n13 163.367
R813 B.n389 B.n14 163.367
R814 B.n389 B.n19 163.367
R815 B.n20 B.n19 163.367
R816 B.n21 B.n20 163.367
R817 B.n394 B.n21 163.367
R818 B.n394 B.n26 163.367
R819 B.n27 B.n26 163.367
R820 B.n28 B.n27 163.367
R821 B.n399 B.n28 163.367
R822 B.n399 B.n33 163.367
R823 B.n34 B.n33 163.367
R824 B.n35 B.n34 163.367
R825 B.n404 B.n35 163.367
R826 B.n404 B.n40 163.367
R827 B.n41 B.n40 163.367
R828 B.n42 B.n41 163.367
R829 B.n409 B.n42 163.367
R830 B.n409 B.n47 163.367
R831 B.n48 B.n47 163.367
R832 B.n49 B.n48 163.367
R833 B.n414 B.n49 163.367
R834 B.n414 B.n54 163.367
R835 B.n55 B.n54 163.367
R836 B.n56 B.n55 163.367
R837 B.n419 B.n56 163.367
R838 B.n419 B.n61 163.367
R839 B.n62 B.n61 163.367
R840 B.n63 B.n62 163.367
R841 B.n424 B.n63 163.367
R842 B.n424 B.n68 163.367
R843 B.n69 B.n68 163.367
R844 B.n70 B.n69 163.367
R845 B.n501 B.n499 163.367
R846 B.n497 B.n74 163.367
R847 B.n493 B.n491 163.367
R848 B.n489 B.n76 163.367
R849 B.n485 B.n483 163.367
R850 B.n481 B.n78 163.367
R851 B.n477 B.n475 163.367
R852 B.n472 B.n471 163.367
R853 B.n469 B.n84 163.367
R854 B.n465 B.n463 163.367
R855 B.n461 B.n86 163.367
R856 B.n456 B.n454 163.367
R857 B.n452 B.n90 163.367
R858 B.n448 B.n446 163.367
R859 B.n444 B.n92 163.367
R860 B.n440 B.n438 163.367
R861 B.n436 B.n94 163.367
R862 B.n432 B.n430 163.367
R863 B.n185 B.t18 155.668
R864 B.n87 B.t20 155.668
R865 B.n178 B.t11 155.668
R866 B.n79 B.t14 155.668
R867 B.n186 B.t17 122.505
R868 B.n88 B.t21 122.505
R869 B.n179 B.t10 122.505
R870 B.n80 B.t15 122.505
R871 B.n267 B.n164 96.3302
R872 B.n273 B.n164 96.3302
R873 B.n273 B.n159 96.3302
R874 B.n279 B.n159 96.3302
R875 B.n279 B.n160 96.3302
R876 B.n285 B.n152 96.3302
R877 B.n291 B.n152 96.3302
R878 B.n291 B.n148 96.3302
R879 B.n297 B.n148 96.3302
R880 B.n297 B.n143 96.3302
R881 B.n303 B.n143 96.3302
R882 B.n303 B.n144 96.3302
R883 B.n309 B.n136 96.3302
R884 B.n315 B.n136 96.3302
R885 B.n315 B.n132 96.3302
R886 B.n321 B.n132 96.3302
R887 B.n327 B.n128 96.3302
R888 B.n327 B.n124 96.3302
R889 B.n334 B.n124 96.3302
R890 B.n334 B.n333 96.3302
R891 B.n340 B.n117 96.3302
R892 B.n346 B.n117 96.3302
R893 B.n346 B.n113 96.3302
R894 B.n352 B.n113 96.3302
R895 B.n358 B.n109 96.3302
R896 B.n358 B.n104 96.3302
R897 B.n364 B.n104 96.3302
R898 B.n364 B.n105 96.3302
R899 B.n371 B.n97 96.3302
R900 B.n377 B.n97 96.3302
R901 B.n377 B.n4 96.3302
R902 B.n580 B.n4 96.3302
R903 B.n580 B.n579 96.3302
R904 B.n579 B.n578 96.3302
R905 B.n578 B.n8 96.3302
R906 B.n572 B.n8 96.3302
R907 B.n571 B.n570 96.3302
R908 B.n570 B.n15 96.3302
R909 B.n564 B.n15 96.3302
R910 B.n564 B.n563 96.3302
R911 B.n562 B.n22 96.3302
R912 B.n556 B.n22 96.3302
R913 B.n556 B.n555 96.3302
R914 B.n555 B.n554 96.3302
R915 B.n548 B.n32 96.3302
R916 B.n548 B.n547 96.3302
R917 B.n547 B.n546 96.3302
R918 B.n546 B.n36 96.3302
R919 B.n540 B.n539 96.3302
R920 B.n539 B.n538 96.3302
R921 B.n538 B.n43 96.3302
R922 B.n532 B.n43 96.3302
R923 B.n531 B.n530 96.3302
R924 B.n530 B.n50 96.3302
R925 B.n524 B.n50 96.3302
R926 B.n524 B.n523 96.3302
R927 B.n523 B.n522 96.3302
R928 B.n522 B.n57 96.3302
R929 B.n516 B.n57 96.3302
R930 B.n515 B.n514 96.3302
R931 B.n514 B.n64 96.3302
R932 B.n508 B.n64 96.3302
R933 B.n508 B.n507 96.3302
R934 B.n507 B.n506 96.3302
R935 B.n105 B.t22 84.9973
R936 B.t5 B.n571 84.9973
R937 B.n352 B.t6 82.1641
R938 B.t1 B.n562 82.1641
R939 B.n333 B.t2 79.3308
R940 B.n32 B.t4 79.3308
R941 B.n321 B.t3 76.4976
R942 B.n540 B.t0 76.4976
R943 B.n144 B.t23 73.6644
R944 B.t7 B.n531 73.6644
R945 B.n261 B.n169 71.676
R946 B.n259 B.n171 71.676
R947 B.n255 B.n254 71.676
R948 B.n248 B.n173 71.676
R949 B.n247 B.n246 71.676
R950 B.n240 B.n175 71.676
R951 B.n239 B.n238 71.676
R952 B.n232 B.n177 71.676
R953 B.n231 B.n230 71.676
R954 B.n224 B.n182 71.676
R955 B.n223 B.n222 71.676
R956 B.n215 B.n184 71.676
R957 B.n214 B.n213 71.676
R958 B.n207 B.n188 71.676
R959 B.n206 B.n205 71.676
R960 B.n199 B.n190 71.676
R961 B.n198 B.n197 71.676
R962 B.n193 B.n192 71.676
R963 B.n500 B.n72 71.676
R964 B.n499 B.n498 71.676
R965 B.n492 B.n74 71.676
R966 B.n491 B.n490 71.676
R967 B.n484 B.n76 71.676
R968 B.n483 B.n482 71.676
R969 B.n476 B.n78 71.676
R970 B.n475 B.n82 71.676
R971 B.n471 B.n470 71.676
R972 B.n464 B.n84 71.676
R973 B.n463 B.n462 71.676
R974 B.n455 B.n86 71.676
R975 B.n454 B.n453 71.676
R976 B.n447 B.n90 71.676
R977 B.n446 B.n445 71.676
R978 B.n439 B.n92 71.676
R979 B.n438 B.n437 71.676
R980 B.n431 B.n94 71.676
R981 B.n432 B.n431 71.676
R982 B.n437 B.n436 71.676
R983 B.n440 B.n439 71.676
R984 B.n445 B.n444 71.676
R985 B.n448 B.n447 71.676
R986 B.n453 B.n452 71.676
R987 B.n456 B.n455 71.676
R988 B.n462 B.n461 71.676
R989 B.n465 B.n464 71.676
R990 B.n470 B.n469 71.676
R991 B.n472 B.n82 71.676
R992 B.n477 B.n476 71.676
R993 B.n482 B.n481 71.676
R994 B.n485 B.n484 71.676
R995 B.n490 B.n489 71.676
R996 B.n493 B.n492 71.676
R997 B.n498 B.n497 71.676
R998 B.n501 B.n500 71.676
R999 B.n262 B.n261 71.676
R1000 B.n256 B.n171 71.676
R1001 B.n254 B.n253 71.676
R1002 B.n249 B.n248 71.676
R1003 B.n246 B.n245 71.676
R1004 B.n241 B.n240 71.676
R1005 B.n238 B.n237 71.676
R1006 B.n233 B.n232 71.676
R1007 B.n230 B.n229 71.676
R1008 B.n225 B.n224 71.676
R1009 B.n222 B.n221 71.676
R1010 B.n216 B.n215 71.676
R1011 B.n213 B.n212 71.676
R1012 B.n208 B.n207 71.676
R1013 B.n205 B.n204 71.676
R1014 B.n200 B.n199 71.676
R1015 B.n197 B.n196 71.676
R1016 B.n192 B.n167 71.676
R1017 B.n219 B.n186 59.5399
R1018 B.n180 B.n179 59.5399
R1019 B.n81 B.n80 59.5399
R1020 B.n458 B.n88 59.5399
R1021 B.n160 B.t9 50.9986
R1022 B.t13 B.n515 50.9986
R1023 B.n285 B.t9 45.3321
R1024 B.n516 B.t13 45.3321
R1025 B.n504 B.n503 34.8103
R1026 B.n429 B.n428 34.8103
R1027 B.n269 B.n166 34.8103
R1028 B.n265 B.n264 34.8103
R1029 B.n186 B.n185 33.1641
R1030 B.n179 B.n178 33.1641
R1031 B.n80 B.n79 33.1641
R1032 B.n88 B.n87 33.1641
R1033 B.n309 B.t23 22.6663
R1034 B.n532 B.t7 22.6663
R1035 B.t3 B.n128 19.8331
R1036 B.t0 B.n36 19.8331
R1037 B B.n582 18.0485
R1038 B.n340 B.t2 16.9999
R1039 B.n554 B.t4 16.9999
R1040 B.t6 B.n109 14.1666
R1041 B.n563 B.t1 14.1666
R1042 B.n371 B.t22 11.3334
R1043 B.n572 B.t5 11.3334
R1044 B.n503 B.n502 10.6151
R1045 B.n502 B.n73 10.6151
R1046 B.n496 B.n73 10.6151
R1047 B.n496 B.n495 10.6151
R1048 B.n495 B.n494 10.6151
R1049 B.n494 B.n75 10.6151
R1050 B.n488 B.n75 10.6151
R1051 B.n488 B.n487 10.6151
R1052 B.n487 B.n486 10.6151
R1053 B.n486 B.n77 10.6151
R1054 B.n480 B.n77 10.6151
R1055 B.n480 B.n479 10.6151
R1056 B.n479 B.n478 10.6151
R1057 B.n474 B.n473 10.6151
R1058 B.n473 B.n83 10.6151
R1059 B.n468 B.n83 10.6151
R1060 B.n468 B.n467 10.6151
R1061 B.n467 B.n466 10.6151
R1062 B.n466 B.n85 10.6151
R1063 B.n460 B.n85 10.6151
R1064 B.n460 B.n459 10.6151
R1065 B.n457 B.n89 10.6151
R1066 B.n451 B.n89 10.6151
R1067 B.n451 B.n450 10.6151
R1068 B.n450 B.n449 10.6151
R1069 B.n449 B.n91 10.6151
R1070 B.n443 B.n91 10.6151
R1071 B.n443 B.n442 10.6151
R1072 B.n442 B.n441 10.6151
R1073 B.n441 B.n93 10.6151
R1074 B.n435 B.n93 10.6151
R1075 B.n435 B.n434 10.6151
R1076 B.n434 B.n433 10.6151
R1077 B.n433 B.n429 10.6151
R1078 B.n270 B.n269 10.6151
R1079 B.n271 B.n270 10.6151
R1080 B.n271 B.n157 10.6151
R1081 B.n281 B.n157 10.6151
R1082 B.n282 B.n281 10.6151
R1083 B.n283 B.n282 10.6151
R1084 B.n283 B.n150 10.6151
R1085 B.n293 B.n150 10.6151
R1086 B.n294 B.n293 10.6151
R1087 B.n295 B.n294 10.6151
R1088 B.n295 B.n141 10.6151
R1089 B.n305 B.n141 10.6151
R1090 B.n306 B.n305 10.6151
R1091 B.n307 B.n306 10.6151
R1092 B.n307 B.n134 10.6151
R1093 B.n317 B.n134 10.6151
R1094 B.n318 B.n317 10.6151
R1095 B.n319 B.n318 10.6151
R1096 B.n319 B.n126 10.6151
R1097 B.n329 B.n126 10.6151
R1098 B.n330 B.n329 10.6151
R1099 B.n331 B.n330 10.6151
R1100 B.n331 B.n119 10.6151
R1101 B.n342 B.n119 10.6151
R1102 B.n343 B.n342 10.6151
R1103 B.n344 B.n343 10.6151
R1104 B.n344 B.n111 10.6151
R1105 B.n354 B.n111 10.6151
R1106 B.n355 B.n354 10.6151
R1107 B.n356 B.n355 10.6151
R1108 B.n356 B.n102 10.6151
R1109 B.n366 B.n102 10.6151
R1110 B.n367 B.n366 10.6151
R1111 B.n369 B.n367 10.6151
R1112 B.n369 B.n368 10.6151
R1113 B.n368 B.n95 10.6151
R1114 B.n380 B.n95 10.6151
R1115 B.n381 B.n380 10.6151
R1116 B.n382 B.n381 10.6151
R1117 B.n383 B.n382 10.6151
R1118 B.n385 B.n383 10.6151
R1119 B.n386 B.n385 10.6151
R1120 B.n387 B.n386 10.6151
R1121 B.n388 B.n387 10.6151
R1122 B.n390 B.n388 10.6151
R1123 B.n391 B.n390 10.6151
R1124 B.n392 B.n391 10.6151
R1125 B.n393 B.n392 10.6151
R1126 B.n395 B.n393 10.6151
R1127 B.n396 B.n395 10.6151
R1128 B.n397 B.n396 10.6151
R1129 B.n398 B.n397 10.6151
R1130 B.n400 B.n398 10.6151
R1131 B.n401 B.n400 10.6151
R1132 B.n402 B.n401 10.6151
R1133 B.n403 B.n402 10.6151
R1134 B.n405 B.n403 10.6151
R1135 B.n406 B.n405 10.6151
R1136 B.n407 B.n406 10.6151
R1137 B.n408 B.n407 10.6151
R1138 B.n410 B.n408 10.6151
R1139 B.n411 B.n410 10.6151
R1140 B.n412 B.n411 10.6151
R1141 B.n413 B.n412 10.6151
R1142 B.n415 B.n413 10.6151
R1143 B.n416 B.n415 10.6151
R1144 B.n417 B.n416 10.6151
R1145 B.n418 B.n417 10.6151
R1146 B.n420 B.n418 10.6151
R1147 B.n421 B.n420 10.6151
R1148 B.n422 B.n421 10.6151
R1149 B.n423 B.n422 10.6151
R1150 B.n425 B.n423 10.6151
R1151 B.n426 B.n425 10.6151
R1152 B.n427 B.n426 10.6151
R1153 B.n428 B.n427 10.6151
R1154 B.n264 B.n263 10.6151
R1155 B.n263 B.n170 10.6151
R1156 B.n258 B.n170 10.6151
R1157 B.n258 B.n257 10.6151
R1158 B.n257 B.n172 10.6151
R1159 B.n252 B.n172 10.6151
R1160 B.n252 B.n251 10.6151
R1161 B.n251 B.n250 10.6151
R1162 B.n250 B.n174 10.6151
R1163 B.n244 B.n174 10.6151
R1164 B.n244 B.n243 10.6151
R1165 B.n243 B.n242 10.6151
R1166 B.n242 B.n176 10.6151
R1167 B.n236 B.n235 10.6151
R1168 B.n235 B.n234 10.6151
R1169 B.n234 B.n181 10.6151
R1170 B.n228 B.n181 10.6151
R1171 B.n228 B.n227 10.6151
R1172 B.n227 B.n226 10.6151
R1173 B.n226 B.n183 10.6151
R1174 B.n220 B.n183 10.6151
R1175 B.n218 B.n217 10.6151
R1176 B.n217 B.n187 10.6151
R1177 B.n211 B.n187 10.6151
R1178 B.n211 B.n210 10.6151
R1179 B.n210 B.n209 10.6151
R1180 B.n209 B.n189 10.6151
R1181 B.n203 B.n189 10.6151
R1182 B.n203 B.n202 10.6151
R1183 B.n202 B.n201 10.6151
R1184 B.n201 B.n191 10.6151
R1185 B.n195 B.n191 10.6151
R1186 B.n195 B.n194 10.6151
R1187 B.n194 B.n166 10.6151
R1188 B.n265 B.n162 10.6151
R1189 B.n275 B.n162 10.6151
R1190 B.n276 B.n275 10.6151
R1191 B.n277 B.n276 10.6151
R1192 B.n277 B.n154 10.6151
R1193 B.n287 B.n154 10.6151
R1194 B.n288 B.n287 10.6151
R1195 B.n289 B.n288 10.6151
R1196 B.n289 B.n146 10.6151
R1197 B.n299 B.n146 10.6151
R1198 B.n300 B.n299 10.6151
R1199 B.n301 B.n300 10.6151
R1200 B.n301 B.n138 10.6151
R1201 B.n311 B.n138 10.6151
R1202 B.n312 B.n311 10.6151
R1203 B.n313 B.n312 10.6151
R1204 B.n313 B.n130 10.6151
R1205 B.n323 B.n130 10.6151
R1206 B.n324 B.n323 10.6151
R1207 B.n325 B.n324 10.6151
R1208 B.n325 B.n122 10.6151
R1209 B.n336 B.n122 10.6151
R1210 B.n337 B.n336 10.6151
R1211 B.n338 B.n337 10.6151
R1212 B.n338 B.n115 10.6151
R1213 B.n348 B.n115 10.6151
R1214 B.n349 B.n348 10.6151
R1215 B.n350 B.n349 10.6151
R1216 B.n350 B.n107 10.6151
R1217 B.n360 B.n107 10.6151
R1218 B.n361 B.n360 10.6151
R1219 B.n362 B.n361 10.6151
R1220 B.n362 B.n99 10.6151
R1221 B.n373 B.n99 10.6151
R1222 B.n374 B.n373 10.6151
R1223 B.n375 B.n374 10.6151
R1224 B.n375 B.n0 10.6151
R1225 B.n576 B.n1 10.6151
R1226 B.n576 B.n575 10.6151
R1227 B.n575 B.n574 10.6151
R1228 B.n574 B.n10 10.6151
R1229 B.n568 B.n10 10.6151
R1230 B.n568 B.n567 10.6151
R1231 B.n567 B.n566 10.6151
R1232 B.n566 B.n17 10.6151
R1233 B.n560 B.n17 10.6151
R1234 B.n560 B.n559 10.6151
R1235 B.n559 B.n558 10.6151
R1236 B.n558 B.n24 10.6151
R1237 B.n552 B.n24 10.6151
R1238 B.n552 B.n551 10.6151
R1239 B.n551 B.n550 10.6151
R1240 B.n550 B.n30 10.6151
R1241 B.n544 B.n30 10.6151
R1242 B.n544 B.n543 10.6151
R1243 B.n543 B.n542 10.6151
R1244 B.n542 B.n38 10.6151
R1245 B.n536 B.n38 10.6151
R1246 B.n536 B.n535 10.6151
R1247 B.n535 B.n534 10.6151
R1248 B.n534 B.n45 10.6151
R1249 B.n528 B.n45 10.6151
R1250 B.n528 B.n527 10.6151
R1251 B.n527 B.n526 10.6151
R1252 B.n526 B.n52 10.6151
R1253 B.n520 B.n52 10.6151
R1254 B.n520 B.n519 10.6151
R1255 B.n519 B.n518 10.6151
R1256 B.n518 B.n59 10.6151
R1257 B.n512 B.n59 10.6151
R1258 B.n512 B.n511 10.6151
R1259 B.n511 B.n510 10.6151
R1260 B.n510 B.n66 10.6151
R1261 B.n504 B.n66 10.6151
R1262 B.n474 B.n81 6.5566
R1263 B.n459 B.n458 6.5566
R1264 B.n236 B.n180 6.5566
R1265 B.n220 B.n219 6.5566
R1266 B.n478 B.n81 4.05904
R1267 B.n458 B.n457 4.05904
R1268 B.n180 B.n176 4.05904
R1269 B.n219 B.n218 4.05904
R1270 B.n582 B.n0 2.81026
R1271 B.n582 B.n1 2.81026
R1272 VP.n35 VP.n34 177.448
R1273 VP.n60 VP.n59 177.448
R1274 VP.n33 VP.n32 177.448
R1275 VP.n16 VP.n15 161.3
R1276 VP.n17 VP.n12 161.3
R1277 VP.n20 VP.n19 161.3
R1278 VP.n21 VP.n11 161.3
R1279 VP.n23 VP.n22 161.3
R1280 VP.n24 VP.n10 161.3
R1281 VP.n27 VP.n26 161.3
R1282 VP.n28 VP.n9 161.3
R1283 VP.n30 VP.n29 161.3
R1284 VP.n31 VP.n8 161.3
R1285 VP.n58 VP.n0 161.3
R1286 VP.n57 VP.n56 161.3
R1287 VP.n55 VP.n1 161.3
R1288 VP.n54 VP.n53 161.3
R1289 VP.n51 VP.n2 161.3
R1290 VP.n50 VP.n49 161.3
R1291 VP.n48 VP.n3 161.3
R1292 VP.n47 VP.n46 161.3
R1293 VP.n44 VP.n4 161.3
R1294 VP.n43 VP.n42 161.3
R1295 VP.n41 VP.n40 161.3
R1296 VP.n39 VP.n6 161.3
R1297 VP.n38 VP.n37 161.3
R1298 VP.n36 VP.n7 161.3
R1299 VP.n14 VP.t2 76.3298
R1300 VP.n39 VP.n38 56.5193
R1301 VP.n57 VP.n1 56.5193
R1302 VP.n30 VP.n9 56.5193
R1303 VP.n44 VP.n43 50.6917
R1304 VP.n51 VP.n50 50.6917
R1305 VP.n24 VP.n23 50.6917
R1306 VP.n17 VP.n16 50.6917
R1307 VP.n14 VP.n13 43.6963
R1308 VP.n34 VP.t9 43.4853
R1309 VP.n5 VP.t0 43.4853
R1310 VP.n45 VP.t5 43.4853
R1311 VP.n52 VP.t4 43.4853
R1312 VP.n59 VP.t8 43.4853
R1313 VP.n32 VP.t1 43.4853
R1314 VP.n25 VP.t7 43.4853
R1315 VP.n18 VP.t3 43.4853
R1316 VP.n13 VP.t6 43.4853
R1317 VP.n35 VP.n33 39.1482
R1318 VP.n46 VP.n44 30.2951
R1319 VP.n50 VP.n3 30.2951
R1320 VP.n23 VP.n11 30.2951
R1321 VP.n19 VP.n17 30.2951
R1322 VP.n38 VP.n7 24.4675
R1323 VP.n40 VP.n39 24.4675
R1324 VP.n53 VP.n1 24.4675
R1325 VP.n58 VP.n57 24.4675
R1326 VP.n31 VP.n30 24.4675
R1327 VP.n26 VP.n9 24.4675
R1328 VP.n43 VP.n5 22.5101
R1329 VP.n52 VP.n51 22.5101
R1330 VP.n25 VP.n24 22.5101
R1331 VP.n16 VP.n13 22.5101
R1332 VP.n15 VP.n14 17.9509
R1333 VP.n46 VP.n45 12.234
R1334 VP.n45 VP.n3 12.234
R1335 VP.n19 VP.n18 12.234
R1336 VP.n18 VP.n11 12.234
R1337 VP.n34 VP.n7 8.31928
R1338 VP.n59 VP.n58 8.31928
R1339 VP.n32 VP.n31 8.31928
R1340 VP.n40 VP.n5 1.95786
R1341 VP.n53 VP.n52 1.95786
R1342 VP.n26 VP.n25 1.95786
R1343 VP.n15 VP.n12 0.189894
R1344 VP.n20 VP.n12 0.189894
R1345 VP.n21 VP.n20 0.189894
R1346 VP.n22 VP.n21 0.189894
R1347 VP.n22 VP.n10 0.189894
R1348 VP.n27 VP.n10 0.189894
R1349 VP.n28 VP.n27 0.189894
R1350 VP.n29 VP.n28 0.189894
R1351 VP.n29 VP.n8 0.189894
R1352 VP.n33 VP.n8 0.189894
R1353 VP.n36 VP.n35 0.189894
R1354 VP.n37 VP.n36 0.189894
R1355 VP.n37 VP.n6 0.189894
R1356 VP.n41 VP.n6 0.189894
R1357 VP.n42 VP.n41 0.189894
R1358 VP.n42 VP.n4 0.189894
R1359 VP.n47 VP.n4 0.189894
R1360 VP.n48 VP.n47 0.189894
R1361 VP.n49 VP.n48 0.189894
R1362 VP.n49 VP.n2 0.189894
R1363 VP.n54 VP.n2 0.189894
R1364 VP.n55 VP.n54 0.189894
R1365 VP.n56 VP.n55 0.189894
R1366 VP.n56 VP.n0 0.189894
R1367 VP.n60 VP.n0 0.189894
R1368 VP VP.n60 0.0516364
R1369 VDD1.n6 VDD1.n0 289.615
R1370 VDD1.n19 VDD1.n13 289.615
R1371 VDD1.n7 VDD1.n6 185
R1372 VDD1.n5 VDD1.n4 185
R1373 VDD1.n18 VDD1.n17 185
R1374 VDD1.n20 VDD1.n19 185
R1375 VDD1.n3 VDD1.t7 151.613
R1376 VDD1.n16 VDD1.t0 151.613
R1377 VDD1.n6 VDD1.n5 104.615
R1378 VDD1.n19 VDD1.n18 104.615
R1379 VDD1.n27 VDD1.n26 87.7549
R1380 VDD1.n12 VDD1.n11 86.7047
R1381 VDD1.n29 VDD1.n28 86.7046
R1382 VDD1.n25 VDD1.n24 86.7046
R1383 VDD1.n5 VDD1.t7 52.3082
R1384 VDD1.n18 VDD1.t0 52.3082
R1385 VDD1.n12 VDD1.n10 52.0837
R1386 VDD1.n25 VDD1.n23 52.0837
R1387 VDD1.n29 VDD1.n27 34.1841
R1388 VDD1.n4 VDD1.n3 15.3979
R1389 VDD1.n17 VDD1.n16 15.3979
R1390 VDD1.n7 VDD1.n2 12.8005
R1391 VDD1.n20 VDD1.n15 12.8005
R1392 VDD1.n8 VDD1.n0 12.0247
R1393 VDD1.n21 VDD1.n13 12.0247
R1394 VDD1.n10 VDD1.n9 9.45567
R1395 VDD1.n23 VDD1.n22 9.45567
R1396 VDD1.n9 VDD1.n8 9.3005
R1397 VDD1.n2 VDD1.n1 9.3005
R1398 VDD1.n22 VDD1.n21 9.3005
R1399 VDD1.n15 VDD1.n14 9.3005
R1400 VDD1.n28 VDD1.t2 7.95231
R1401 VDD1.n28 VDD1.t8 7.95231
R1402 VDD1.n11 VDD1.t3 7.95231
R1403 VDD1.n11 VDD1.t6 7.95231
R1404 VDD1.n26 VDD1.t5 7.95231
R1405 VDD1.n26 VDD1.t1 7.95231
R1406 VDD1.n24 VDD1.t9 7.95231
R1407 VDD1.n24 VDD1.t4 7.95231
R1408 VDD1.n3 VDD1.n1 4.69785
R1409 VDD1.n16 VDD1.n14 4.69785
R1410 VDD1.n10 VDD1.n0 1.93989
R1411 VDD1.n23 VDD1.n13 1.93989
R1412 VDD1.n8 VDD1.n7 1.16414
R1413 VDD1.n21 VDD1.n20 1.16414
R1414 VDD1 VDD1.n29 1.04791
R1415 VDD1 VDD1.n12 0.427224
R1416 VDD1.n4 VDD1.n2 0.388379
R1417 VDD1.n17 VDD1.n15 0.388379
R1418 VDD1.n27 VDD1.n25 0.313688
R1419 VDD1.n9 VDD1.n1 0.155672
R1420 VDD1.n22 VDD1.n14 0.155672
C0 VP VN 4.8486f
C1 VP VDD1 2.5176f
C2 VTAIL VN 2.93857f
C3 VTAIL VDD1 4.95807f
C4 VDD2 VP 0.433597f
C5 VDD2 VTAIL 5.0026f
C6 VN VDD1 0.156373f
C7 VTAIL VP 2.95275f
C8 VDD2 VN 2.24301f
C9 VDD2 VDD1 1.37971f
C10 VDD2 B 4.072138f
C11 VDD1 B 4.049158f
C12 VTAIL B 3.258985f
C13 VN B 11.43835f
C14 VP B 9.942533f
C15 VDD1.n0 B 0.031891f
C16 VDD1.n1 B 0.179336f
C17 VDD1.n2 B 0.012872f
C18 VDD1.t7 B 0.05246f
C19 VDD1.n3 B 0.084298f
C20 VDD1.n4 B 0.017222f
C21 VDD1.n5 B 0.022818f
C22 VDD1.n6 B 0.062718f
C23 VDD1.n7 B 0.013629f
C24 VDD1.n8 B 0.012872f
C25 VDD1.n9 B 0.058312f
C26 VDD1.n10 B 0.055949f
C27 VDD1.t3 B 0.047132f
C28 VDD1.t6 B 0.047132f
C29 VDD1.n11 B 0.334225f
C30 VDD1.n12 B 0.478926f
C31 VDD1.n13 B 0.031891f
C32 VDD1.n14 B 0.179336f
C33 VDD1.n15 B 0.012872f
C34 VDD1.t0 B 0.05246f
C35 VDD1.n16 B 0.084298f
C36 VDD1.n17 B 0.017222f
C37 VDD1.n18 B 0.022818f
C38 VDD1.n19 B 0.062718f
C39 VDD1.n20 B 0.013629f
C40 VDD1.n21 B 0.012872f
C41 VDD1.n22 B 0.058312f
C42 VDD1.n23 B 0.055949f
C43 VDD1.t9 B 0.047132f
C44 VDD1.t4 B 0.047132f
C45 VDD1.n24 B 0.334224f
C46 VDD1.n25 B 0.471937f
C47 VDD1.t5 B 0.047132f
C48 VDD1.t1 B 0.047132f
C49 VDD1.n26 B 0.338774f
C50 VDD1.n27 B 1.69395f
C51 VDD1.t2 B 0.047132f
C52 VDD1.t8 B 0.047132f
C53 VDD1.n28 B 0.334223f
C54 VDD1.n29 B 1.81416f
C55 VP.n0 B 0.037495f
C56 VP.t8 B 0.312736f
C57 VP.n1 B 0.061531f
C58 VP.n2 B 0.037495f
C59 VP.t4 B 0.312736f
C60 VP.n3 B 0.057675f
C61 VP.n4 B 0.037495f
C62 VP.t0 B 0.312736f
C63 VP.n5 B 0.154858f
C64 VP.n6 B 0.037495f
C65 VP.n7 B 0.047111f
C66 VP.n8 B 0.037495f
C67 VP.t1 B 0.312736f
C68 VP.n9 B 0.061531f
C69 VP.n10 B 0.037495f
C70 VP.t7 B 0.312736f
C71 VP.n11 B 0.057675f
C72 VP.n12 B 0.037495f
C73 VP.t6 B 0.312736f
C74 VP.n13 B 0.235812f
C75 VP.t2 B 0.437207f
C76 VP.n14 B 0.214719f
C77 VP.n15 B 0.232835f
C78 VP.n16 B 0.065694f
C79 VP.n17 B 0.035982f
C80 VP.t3 B 0.312736f
C81 VP.n18 B 0.154858f
C82 VP.n19 B 0.057675f
C83 VP.n20 B 0.037495f
C84 VP.n21 B 0.037495f
C85 VP.n22 B 0.037495f
C86 VP.n23 B 0.035982f
C87 VP.n24 B 0.065694f
C88 VP.n25 B 0.154858f
C89 VP.n26 B 0.038141f
C90 VP.n27 B 0.037495f
C91 VP.n28 B 0.037495f
C92 VP.n29 B 0.037495f
C93 VP.n30 B 0.047948f
C94 VP.n31 B 0.047111f
C95 VP.n32 B 0.221517f
C96 VP.n33 B 1.37915f
C97 VP.t9 B 0.312736f
C98 VP.n34 B 0.221517f
C99 VP.n35 B 1.41357f
C100 VP.n36 B 0.037495f
C101 VP.n37 B 0.037495f
C102 VP.n38 B 0.047948f
C103 VP.n39 B 0.061531f
C104 VP.n40 B 0.038141f
C105 VP.n41 B 0.037495f
C106 VP.n42 B 0.037495f
C107 VP.n43 B 0.065694f
C108 VP.n44 B 0.035982f
C109 VP.t5 B 0.312736f
C110 VP.n45 B 0.154858f
C111 VP.n46 B 0.057675f
C112 VP.n47 B 0.037495f
C113 VP.n48 B 0.037495f
C114 VP.n49 B 0.037495f
C115 VP.n50 B 0.035982f
C116 VP.n51 B 0.065694f
C117 VP.n52 B 0.154858f
C118 VP.n53 B 0.038141f
C119 VP.n54 B 0.037495f
C120 VP.n55 B 0.037495f
C121 VP.n56 B 0.037495f
C122 VP.n57 B 0.047948f
C123 VP.n58 B 0.047111f
C124 VP.n59 B 0.221517f
C125 VP.n60 B 0.035731f
C126 VDD2.n0 B 0.030981f
C127 VDD2.n1 B 0.174218f
C128 VDD2.n2 B 0.012504f
C129 VDD2.t3 B 0.050963f
C130 VDD2.n3 B 0.081892f
C131 VDD2.n4 B 0.01673f
C132 VDD2.n5 B 0.022166f
C133 VDD2.n6 B 0.060928f
C134 VDD2.n7 B 0.01324f
C135 VDD2.n8 B 0.012504f
C136 VDD2.n9 B 0.056648f
C137 VDD2.n10 B 0.054352f
C138 VDD2.t6 B 0.045787f
C139 VDD2.t0 B 0.045787f
C140 VDD2.n11 B 0.324685f
C141 VDD2.n12 B 0.458468f
C142 VDD2.t5 B 0.045787f
C143 VDD2.t9 B 0.045787f
C144 VDD2.n13 B 0.329105f
C145 VDD2.n14 B 1.56466f
C146 VDD2.n15 B 0.030981f
C147 VDD2.n16 B 0.174218f
C148 VDD2.n17 B 0.012504f
C149 VDD2.t1 B 0.050963f
C150 VDD2.n18 B 0.081892f
C151 VDD2.n19 B 0.01673f
C152 VDD2.n20 B 0.022166f
C153 VDD2.n21 B 0.060928f
C154 VDD2.n22 B 0.01324f
C155 VDD2.n23 B 0.012504f
C156 VDD2.n24 B 0.056648f
C157 VDD2.n25 B 0.049909f
C158 VDD2.n26 B 1.54571f
C159 VDD2.t7 B 0.045787f
C160 VDD2.t2 B 0.045787f
C161 VDD2.n27 B 0.324686f
C162 VDD2.n28 B 0.312723f
C163 VDD2.t8 B 0.045787f
C164 VDD2.t4 B 0.045787f
C165 VDD2.n29 B 0.329085f
C166 VTAIL.t12 B 0.063345f
C167 VTAIL.t15 B 0.063345f
C168 VTAIL.n0 B 0.394564f
C169 VTAIL.n1 B 0.492243f
C170 VTAIL.n2 B 0.04286f
C171 VTAIL.n3 B 0.241022f
C172 VTAIL.n4 B 0.017299f
C173 VTAIL.t8 B 0.070505f
C174 VTAIL.n5 B 0.113294f
C175 VTAIL.n6 B 0.023146f
C176 VTAIL.n7 B 0.030666f
C177 VTAIL.n8 B 0.084291f
C178 VTAIL.n9 B 0.018316f
C179 VTAIL.n10 B 0.017299f
C180 VTAIL.n11 B 0.07837f
C181 VTAIL.n12 B 0.046849f
C182 VTAIL.n13 B 0.30784f
C183 VTAIL.t2 B 0.063345f
C184 VTAIL.t6 B 0.063345f
C185 VTAIL.n14 B 0.394564f
C186 VTAIL.n15 B 0.552157f
C187 VTAIL.t19 B 0.063345f
C188 VTAIL.t3 B 0.063345f
C189 VTAIL.n16 B 0.394564f
C190 VTAIL.n17 B 1.36504f
C191 VTAIL.t10 B 0.063345f
C192 VTAIL.t18 B 0.063345f
C193 VTAIL.n18 B 0.394567f
C194 VTAIL.n19 B 1.36503f
C195 VTAIL.t16 B 0.063345f
C196 VTAIL.t14 B 0.063345f
C197 VTAIL.n20 B 0.394567f
C198 VTAIL.n21 B 0.552155f
C199 VTAIL.n22 B 0.04286f
C200 VTAIL.n23 B 0.241022f
C201 VTAIL.n24 B 0.017299f
C202 VTAIL.t9 B 0.070505f
C203 VTAIL.n25 B 0.113294f
C204 VTAIL.n26 B 0.023146f
C205 VTAIL.n27 B 0.030666f
C206 VTAIL.n28 B 0.084291f
C207 VTAIL.n29 B 0.018316f
C208 VTAIL.n30 B 0.017299f
C209 VTAIL.n31 B 0.07837f
C210 VTAIL.n32 B 0.046849f
C211 VTAIL.n33 B 0.30784f
C212 VTAIL.t5 B 0.063345f
C213 VTAIL.t1 B 0.063345f
C214 VTAIL.n34 B 0.394567f
C215 VTAIL.n35 B 0.524433f
C216 VTAIL.t4 B 0.063345f
C217 VTAIL.t0 B 0.063345f
C218 VTAIL.n36 B 0.394567f
C219 VTAIL.n37 B 0.552155f
C220 VTAIL.n38 B 0.04286f
C221 VTAIL.n39 B 0.241022f
C222 VTAIL.n40 B 0.017299f
C223 VTAIL.t7 B 0.070505f
C224 VTAIL.n41 B 0.113294f
C225 VTAIL.n42 B 0.023146f
C226 VTAIL.n43 B 0.030666f
C227 VTAIL.n44 B 0.084291f
C228 VTAIL.n45 B 0.018316f
C229 VTAIL.n46 B 0.017299f
C230 VTAIL.n47 B 0.07837f
C231 VTAIL.n48 B 0.046849f
C232 VTAIL.n49 B 0.995525f
C233 VTAIL.n50 B 0.04286f
C234 VTAIL.n51 B 0.241022f
C235 VTAIL.n52 B 0.017299f
C236 VTAIL.t13 B 0.070505f
C237 VTAIL.n53 B 0.113294f
C238 VTAIL.n54 B 0.023146f
C239 VTAIL.n55 B 0.030666f
C240 VTAIL.n56 B 0.084291f
C241 VTAIL.n57 B 0.018316f
C242 VTAIL.n58 B 0.017299f
C243 VTAIL.n59 B 0.07837f
C244 VTAIL.n60 B 0.046849f
C245 VTAIL.n61 B 0.995525f
C246 VTAIL.t17 B 0.063345f
C247 VTAIL.t11 B 0.063345f
C248 VTAIL.n62 B 0.394564f
C249 VTAIL.n63 B 0.431435f
C250 VN.n0 B 0.035856f
C251 VN.t0 B 0.299061f
C252 VN.n1 B 0.05884f
C253 VN.n2 B 0.035856f
C254 VN.t4 B 0.299061f
C255 VN.n3 B 0.055153f
C256 VN.n4 B 0.035856f
C257 VN.t3 B 0.299061f
C258 VN.n5 B 0.2255f
C259 VN.t6 B 0.418088f
C260 VN.n6 B 0.20533f
C261 VN.n7 B 0.222653f
C262 VN.n8 B 0.062821f
C263 VN.n9 B 0.034408f
C264 VN.t9 B 0.299061f
C265 VN.n10 B 0.148087f
C266 VN.n11 B 0.055153f
C267 VN.n12 B 0.035856f
C268 VN.n13 B 0.035856f
C269 VN.n14 B 0.035856f
C270 VN.n15 B 0.034408f
C271 VN.n16 B 0.062821f
C272 VN.n17 B 0.148087f
C273 VN.n18 B 0.036473f
C274 VN.n19 B 0.035856f
C275 VN.n20 B 0.035856f
C276 VN.n21 B 0.035856f
C277 VN.n22 B 0.045852f
C278 VN.n23 B 0.045051f
C279 VN.n24 B 0.21183f
C280 VN.n25 B 0.034168f
C281 VN.n26 B 0.035856f
C282 VN.t8 B 0.299061f
C283 VN.n27 B 0.05884f
C284 VN.n28 B 0.035856f
C285 VN.t2 B 0.299061f
C286 VN.n29 B 0.055153f
C287 VN.n30 B 0.035856f
C288 VN.t7 B 0.299061f
C289 VN.n31 B 0.148087f
C290 VN.t1 B 0.299061f
C291 VN.n32 B 0.2255f
C292 VN.t5 B 0.418088f
C293 VN.n33 B 0.20533f
C294 VN.n34 B 0.222653f
C295 VN.n35 B 0.062821f
C296 VN.n36 B 0.034408f
C297 VN.n37 B 0.055153f
C298 VN.n38 B 0.035856f
C299 VN.n39 B 0.035856f
C300 VN.n40 B 0.035856f
C301 VN.n41 B 0.034408f
C302 VN.n42 B 0.062821f
C303 VN.n43 B 0.148087f
C304 VN.n44 B 0.036473f
C305 VN.n45 B 0.035856f
C306 VN.n46 B 0.035856f
C307 VN.n47 B 0.035856f
C308 VN.n48 B 0.045852f
C309 VN.n49 B 0.045051f
C310 VN.n50 B 0.21183f
C311 VN.n51 B 1.34248f
.ends

