* NGSPICE file created from diff_pair_sample_1391.ext - technology: sky130A

.subckt diff_pair_sample_1391 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t8 VN.t0 VDD2.t0 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.64
X1 VDD1.t5 VP.t0 VTAIL.t2 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.64
X2 VDD2.t4 VN.t1 VTAIL.t7 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.64
X3 VTAIL.t6 VN.t2 VDD2.t3 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.64
X4 VDD2.t2 VN.t3 VTAIL.t5 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.64
X5 VDD1.t4 VP.t1 VTAIL.t1 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.64
X6 VDD2.t1 VN.t4 VTAIL.t4 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.64
X7 B.t11 B.t9 B.t10 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.64
X8 VTAIL.t11 VP.t2 VDD1.t3 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.64
X9 B.t8 B.t6 B.t7 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.64
X10 VDD2.t5 VN.t5 VTAIL.t3 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.64
X11 VDD1.t2 VP.t3 VTAIL.t10 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=3.20265 ps=19.74 w=19.41 l=3.64
X12 VTAIL.t9 VP.t4 VDD1.t1 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=3.20265 ps=19.74 w=19.41 l=3.64
X13 B.t5 B.t3 B.t4 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.64
X14 B.t2 B.t0 B.t1 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=7.5699 pd=39.6 as=0 ps=0 w=19.41 l=3.64
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n4146_n4850# sky130_fd_pr__pfet_01v8 ad=3.20265 pd=19.74 as=7.5699 ps=39.6 w=19.41 l=3.64
R0 VN.n26 VN.t3 162.023
R1 VN.n6 VN.t1 162.023
R2 VN.n38 VN.n37 161.3
R3 VN.n36 VN.n21 161.3
R4 VN.n35 VN.n34 161.3
R5 VN.n33 VN.n22 161.3
R6 VN.n32 VN.n31 161.3
R7 VN.n30 VN.n23 161.3
R8 VN.n29 VN.n28 161.3
R9 VN.n27 VN.n24 161.3
R10 VN.n18 VN.n17 161.3
R11 VN.n16 VN.n1 161.3
R12 VN.n15 VN.n14 161.3
R13 VN.n13 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n5 VN.t2 128.512
R19 VN.n0 VN.t4 128.512
R20 VN.n25 VN.t0 128.512
R21 VN.n20 VN.t5 128.512
R22 VN.n19 VN.n0 79.3019
R23 VN.n39 VN.n20 79.3019
R24 VN.n6 VN.n5 62.396
R25 VN.n26 VN.n25 62.396
R26 VN VN.n39 58.6685
R27 VN.n11 VN.n2 56.5193
R28 VN.n31 VN.n22 56.5193
R29 VN.n9 VN.n4 24.4675
R30 VN.n10 VN.n9 24.4675
R31 VN.n11 VN.n10 24.4675
R32 VN.n15 VN.n2 24.4675
R33 VN.n16 VN.n15 24.4675
R34 VN.n17 VN.n16 24.4675
R35 VN.n31 VN.n30 24.4675
R36 VN.n30 VN.n29 24.4675
R37 VN.n29 VN.n24 24.4675
R38 VN.n37 VN.n36 24.4675
R39 VN.n36 VN.n35 24.4675
R40 VN.n35 VN.n22 24.4675
R41 VN.n5 VN.n4 12.234
R42 VN.n25 VN.n24 12.234
R43 VN.n17 VN.n0 10.766
R44 VN.n37 VN.n20 10.766
R45 VN.n27 VN.n26 3.13206
R46 VN.n7 VN.n6 3.13206
R47 VN.n39 VN.n38 0.354971
R48 VN.n19 VN.n18 0.354971
R49 VN VN.n19 0.26696
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VDD2.n208 VDD2.n207 585
R65 VDD2.n206 VDD2.n205 585
R66 VDD2.n111 VDD2.n110 585
R67 VDD2.n200 VDD2.n199 585
R68 VDD2.n198 VDD2.n197 585
R69 VDD2.n115 VDD2.n114 585
R70 VDD2.n192 VDD2.n191 585
R71 VDD2.n190 VDD2.n189 585
R72 VDD2.n119 VDD2.n118 585
R73 VDD2.n184 VDD2.n183 585
R74 VDD2.n182 VDD2.n181 585
R75 VDD2.n123 VDD2.n122 585
R76 VDD2.n176 VDD2.n175 585
R77 VDD2.n174 VDD2.n173 585
R78 VDD2.n127 VDD2.n126 585
R79 VDD2.n168 VDD2.n167 585
R80 VDD2.n166 VDD2.n165 585
R81 VDD2.n164 VDD2.n130 585
R82 VDD2.n134 VDD2.n131 585
R83 VDD2.n159 VDD2.n158 585
R84 VDD2.n157 VDD2.n156 585
R85 VDD2.n136 VDD2.n135 585
R86 VDD2.n151 VDD2.n150 585
R87 VDD2.n149 VDD2.n148 585
R88 VDD2.n140 VDD2.n139 585
R89 VDD2.n143 VDD2.n142 585
R90 VDD2.n35 VDD2.n34 585
R91 VDD2.n32 VDD2.n31 585
R92 VDD2.n41 VDD2.n40 585
R93 VDD2.n43 VDD2.n42 585
R94 VDD2.n28 VDD2.n27 585
R95 VDD2.n49 VDD2.n48 585
R96 VDD2.n52 VDD2.n51 585
R97 VDD2.n50 VDD2.n24 585
R98 VDD2.n57 VDD2.n23 585
R99 VDD2.n59 VDD2.n58 585
R100 VDD2.n61 VDD2.n60 585
R101 VDD2.n20 VDD2.n19 585
R102 VDD2.n67 VDD2.n66 585
R103 VDD2.n69 VDD2.n68 585
R104 VDD2.n16 VDD2.n15 585
R105 VDD2.n75 VDD2.n74 585
R106 VDD2.n77 VDD2.n76 585
R107 VDD2.n12 VDD2.n11 585
R108 VDD2.n83 VDD2.n82 585
R109 VDD2.n85 VDD2.n84 585
R110 VDD2.n8 VDD2.n7 585
R111 VDD2.n91 VDD2.n90 585
R112 VDD2.n93 VDD2.n92 585
R113 VDD2.n4 VDD2.n3 585
R114 VDD2.n99 VDD2.n98 585
R115 VDD2.n101 VDD2.n100 585
R116 VDD2.n207 VDD2.n107 498.474
R117 VDD2.n100 VDD2.n0 498.474
R118 VDD2.t5 VDD2.n141 329.036
R119 VDD2.t4 VDD2.n33 329.036
R120 VDD2.n207 VDD2.n206 171.744
R121 VDD2.n206 VDD2.n110 171.744
R122 VDD2.n199 VDD2.n110 171.744
R123 VDD2.n199 VDD2.n198 171.744
R124 VDD2.n198 VDD2.n114 171.744
R125 VDD2.n191 VDD2.n114 171.744
R126 VDD2.n191 VDD2.n190 171.744
R127 VDD2.n190 VDD2.n118 171.744
R128 VDD2.n183 VDD2.n118 171.744
R129 VDD2.n183 VDD2.n182 171.744
R130 VDD2.n182 VDD2.n122 171.744
R131 VDD2.n175 VDD2.n122 171.744
R132 VDD2.n175 VDD2.n174 171.744
R133 VDD2.n174 VDD2.n126 171.744
R134 VDD2.n167 VDD2.n126 171.744
R135 VDD2.n167 VDD2.n166 171.744
R136 VDD2.n166 VDD2.n130 171.744
R137 VDD2.n134 VDD2.n130 171.744
R138 VDD2.n158 VDD2.n134 171.744
R139 VDD2.n158 VDD2.n157 171.744
R140 VDD2.n157 VDD2.n135 171.744
R141 VDD2.n150 VDD2.n135 171.744
R142 VDD2.n150 VDD2.n149 171.744
R143 VDD2.n149 VDD2.n139 171.744
R144 VDD2.n142 VDD2.n139 171.744
R145 VDD2.n34 VDD2.n31 171.744
R146 VDD2.n41 VDD2.n31 171.744
R147 VDD2.n42 VDD2.n41 171.744
R148 VDD2.n42 VDD2.n27 171.744
R149 VDD2.n49 VDD2.n27 171.744
R150 VDD2.n51 VDD2.n49 171.744
R151 VDD2.n51 VDD2.n50 171.744
R152 VDD2.n50 VDD2.n23 171.744
R153 VDD2.n59 VDD2.n23 171.744
R154 VDD2.n60 VDD2.n59 171.744
R155 VDD2.n60 VDD2.n19 171.744
R156 VDD2.n67 VDD2.n19 171.744
R157 VDD2.n68 VDD2.n67 171.744
R158 VDD2.n68 VDD2.n15 171.744
R159 VDD2.n75 VDD2.n15 171.744
R160 VDD2.n76 VDD2.n75 171.744
R161 VDD2.n76 VDD2.n11 171.744
R162 VDD2.n83 VDD2.n11 171.744
R163 VDD2.n84 VDD2.n83 171.744
R164 VDD2.n84 VDD2.n7 171.744
R165 VDD2.n91 VDD2.n7 171.744
R166 VDD2.n92 VDD2.n91 171.744
R167 VDD2.n92 VDD2.n3 171.744
R168 VDD2.n99 VDD2.n3 171.744
R169 VDD2.n100 VDD2.n99 171.744
R170 VDD2.n142 VDD2.t5 85.8723
R171 VDD2.n34 VDD2.t4 85.8723
R172 VDD2.n106 VDD2.n105 70.3888
R173 VDD2 VDD2.n213 70.3859
R174 VDD2.n106 VDD2.n104 53.1211
R175 VDD2.n212 VDD2.n106 51.5709
R176 VDD2.n212 VDD2.n211 50.6096
R177 VDD2.n165 VDD2.n164 13.1884
R178 VDD2.n58 VDD2.n57 13.1884
R179 VDD2.n209 VDD2.n208 12.8005
R180 VDD2.n168 VDD2.n129 12.8005
R181 VDD2.n163 VDD2.n131 12.8005
R182 VDD2.n56 VDD2.n24 12.8005
R183 VDD2.n61 VDD2.n22 12.8005
R184 VDD2.n102 VDD2.n101 12.8005
R185 VDD2.n205 VDD2.n109 12.0247
R186 VDD2.n169 VDD2.n127 12.0247
R187 VDD2.n160 VDD2.n159 12.0247
R188 VDD2.n53 VDD2.n52 12.0247
R189 VDD2.n62 VDD2.n20 12.0247
R190 VDD2.n98 VDD2.n2 12.0247
R191 VDD2.n204 VDD2.n111 11.249
R192 VDD2.n173 VDD2.n172 11.249
R193 VDD2.n156 VDD2.n133 11.249
R194 VDD2.n48 VDD2.n26 11.249
R195 VDD2.n66 VDD2.n65 11.249
R196 VDD2.n97 VDD2.n4 11.249
R197 VDD2.n143 VDD2.n141 10.7239
R198 VDD2.n35 VDD2.n33 10.7239
R199 VDD2.n201 VDD2.n200 10.4732
R200 VDD2.n176 VDD2.n125 10.4732
R201 VDD2.n155 VDD2.n136 10.4732
R202 VDD2.n47 VDD2.n28 10.4732
R203 VDD2.n69 VDD2.n18 10.4732
R204 VDD2.n94 VDD2.n93 10.4732
R205 VDD2.n197 VDD2.n113 9.69747
R206 VDD2.n177 VDD2.n123 9.69747
R207 VDD2.n152 VDD2.n151 9.69747
R208 VDD2.n44 VDD2.n43 9.69747
R209 VDD2.n70 VDD2.n16 9.69747
R210 VDD2.n90 VDD2.n6 9.69747
R211 VDD2.n211 VDD2.n210 9.45567
R212 VDD2.n104 VDD2.n103 9.45567
R213 VDD2.n145 VDD2.n144 9.3005
R214 VDD2.n147 VDD2.n146 9.3005
R215 VDD2.n138 VDD2.n137 9.3005
R216 VDD2.n153 VDD2.n152 9.3005
R217 VDD2.n155 VDD2.n154 9.3005
R218 VDD2.n133 VDD2.n132 9.3005
R219 VDD2.n161 VDD2.n160 9.3005
R220 VDD2.n163 VDD2.n162 9.3005
R221 VDD2.n117 VDD2.n116 9.3005
R222 VDD2.n194 VDD2.n193 9.3005
R223 VDD2.n196 VDD2.n195 9.3005
R224 VDD2.n113 VDD2.n112 9.3005
R225 VDD2.n202 VDD2.n201 9.3005
R226 VDD2.n204 VDD2.n203 9.3005
R227 VDD2.n109 VDD2.n108 9.3005
R228 VDD2.n210 VDD2.n209 9.3005
R229 VDD2.n188 VDD2.n187 9.3005
R230 VDD2.n186 VDD2.n185 9.3005
R231 VDD2.n121 VDD2.n120 9.3005
R232 VDD2.n180 VDD2.n179 9.3005
R233 VDD2.n178 VDD2.n177 9.3005
R234 VDD2.n125 VDD2.n124 9.3005
R235 VDD2.n172 VDD2.n171 9.3005
R236 VDD2.n170 VDD2.n169 9.3005
R237 VDD2.n129 VDD2.n128 9.3005
R238 VDD2.n79 VDD2.n78 9.3005
R239 VDD2.n14 VDD2.n13 9.3005
R240 VDD2.n73 VDD2.n72 9.3005
R241 VDD2.n71 VDD2.n70 9.3005
R242 VDD2.n18 VDD2.n17 9.3005
R243 VDD2.n65 VDD2.n64 9.3005
R244 VDD2.n63 VDD2.n62 9.3005
R245 VDD2.n22 VDD2.n21 9.3005
R246 VDD2.n37 VDD2.n36 9.3005
R247 VDD2.n39 VDD2.n38 9.3005
R248 VDD2.n30 VDD2.n29 9.3005
R249 VDD2.n45 VDD2.n44 9.3005
R250 VDD2.n47 VDD2.n46 9.3005
R251 VDD2.n26 VDD2.n25 9.3005
R252 VDD2.n54 VDD2.n53 9.3005
R253 VDD2.n56 VDD2.n55 9.3005
R254 VDD2.n81 VDD2.n80 9.3005
R255 VDD2.n10 VDD2.n9 9.3005
R256 VDD2.n87 VDD2.n86 9.3005
R257 VDD2.n89 VDD2.n88 9.3005
R258 VDD2.n6 VDD2.n5 9.3005
R259 VDD2.n95 VDD2.n94 9.3005
R260 VDD2.n97 VDD2.n96 9.3005
R261 VDD2.n2 VDD2.n1 9.3005
R262 VDD2.n103 VDD2.n102 9.3005
R263 VDD2.n196 VDD2.n115 8.92171
R264 VDD2.n181 VDD2.n180 8.92171
R265 VDD2.n148 VDD2.n138 8.92171
R266 VDD2.n40 VDD2.n30 8.92171
R267 VDD2.n74 VDD2.n73 8.92171
R268 VDD2.n89 VDD2.n8 8.92171
R269 VDD2.n193 VDD2.n192 8.14595
R270 VDD2.n184 VDD2.n121 8.14595
R271 VDD2.n147 VDD2.n140 8.14595
R272 VDD2.n39 VDD2.n32 8.14595
R273 VDD2.n77 VDD2.n14 8.14595
R274 VDD2.n86 VDD2.n85 8.14595
R275 VDD2.n211 VDD2.n107 7.75445
R276 VDD2.n104 VDD2.n0 7.75445
R277 VDD2.n189 VDD2.n117 7.3702
R278 VDD2.n185 VDD2.n119 7.3702
R279 VDD2.n144 VDD2.n143 7.3702
R280 VDD2.n36 VDD2.n35 7.3702
R281 VDD2.n78 VDD2.n12 7.3702
R282 VDD2.n82 VDD2.n10 7.3702
R283 VDD2.n189 VDD2.n188 6.59444
R284 VDD2.n188 VDD2.n119 6.59444
R285 VDD2.n81 VDD2.n12 6.59444
R286 VDD2.n82 VDD2.n81 6.59444
R287 VDD2.n209 VDD2.n107 6.08283
R288 VDD2.n102 VDD2.n0 6.08283
R289 VDD2.n192 VDD2.n117 5.81868
R290 VDD2.n185 VDD2.n184 5.81868
R291 VDD2.n144 VDD2.n140 5.81868
R292 VDD2.n36 VDD2.n32 5.81868
R293 VDD2.n78 VDD2.n77 5.81868
R294 VDD2.n85 VDD2.n10 5.81868
R295 VDD2.n193 VDD2.n115 5.04292
R296 VDD2.n181 VDD2.n121 5.04292
R297 VDD2.n148 VDD2.n147 5.04292
R298 VDD2.n40 VDD2.n39 5.04292
R299 VDD2.n74 VDD2.n14 5.04292
R300 VDD2.n86 VDD2.n8 5.04292
R301 VDD2.n197 VDD2.n196 4.26717
R302 VDD2.n180 VDD2.n123 4.26717
R303 VDD2.n151 VDD2.n138 4.26717
R304 VDD2.n43 VDD2.n30 4.26717
R305 VDD2.n73 VDD2.n16 4.26717
R306 VDD2.n90 VDD2.n89 4.26717
R307 VDD2.n200 VDD2.n113 3.49141
R308 VDD2.n177 VDD2.n176 3.49141
R309 VDD2.n152 VDD2.n136 3.49141
R310 VDD2.n44 VDD2.n28 3.49141
R311 VDD2.n70 VDD2.n69 3.49141
R312 VDD2.n93 VDD2.n6 3.49141
R313 VDD2.n201 VDD2.n111 2.71565
R314 VDD2.n173 VDD2.n125 2.71565
R315 VDD2.n156 VDD2.n155 2.71565
R316 VDD2.n48 VDD2.n47 2.71565
R317 VDD2.n66 VDD2.n18 2.71565
R318 VDD2.n94 VDD2.n4 2.71565
R319 VDD2 VDD2.n212 2.6255
R320 VDD2.n145 VDD2.n141 2.41282
R321 VDD2.n37 VDD2.n33 2.41282
R322 VDD2.n205 VDD2.n204 1.93989
R323 VDD2.n172 VDD2.n127 1.93989
R324 VDD2.n159 VDD2.n133 1.93989
R325 VDD2.n52 VDD2.n26 1.93989
R326 VDD2.n65 VDD2.n20 1.93989
R327 VDD2.n98 VDD2.n97 1.93989
R328 VDD2.n213 VDD2.t0 1.67515
R329 VDD2.n213 VDD2.t2 1.67515
R330 VDD2.n105 VDD2.t3 1.67515
R331 VDD2.n105 VDD2.t1 1.67515
R332 VDD2.n208 VDD2.n109 1.16414
R333 VDD2.n169 VDD2.n168 1.16414
R334 VDD2.n160 VDD2.n131 1.16414
R335 VDD2.n53 VDD2.n24 1.16414
R336 VDD2.n62 VDD2.n61 1.16414
R337 VDD2.n101 VDD2.n2 1.16414
R338 VDD2.n165 VDD2.n129 0.388379
R339 VDD2.n164 VDD2.n163 0.388379
R340 VDD2.n57 VDD2.n56 0.388379
R341 VDD2.n58 VDD2.n22 0.388379
R342 VDD2.n210 VDD2.n108 0.155672
R343 VDD2.n203 VDD2.n108 0.155672
R344 VDD2.n203 VDD2.n202 0.155672
R345 VDD2.n202 VDD2.n112 0.155672
R346 VDD2.n195 VDD2.n112 0.155672
R347 VDD2.n195 VDD2.n194 0.155672
R348 VDD2.n194 VDD2.n116 0.155672
R349 VDD2.n187 VDD2.n116 0.155672
R350 VDD2.n187 VDD2.n186 0.155672
R351 VDD2.n186 VDD2.n120 0.155672
R352 VDD2.n179 VDD2.n120 0.155672
R353 VDD2.n179 VDD2.n178 0.155672
R354 VDD2.n178 VDD2.n124 0.155672
R355 VDD2.n171 VDD2.n124 0.155672
R356 VDD2.n171 VDD2.n170 0.155672
R357 VDD2.n170 VDD2.n128 0.155672
R358 VDD2.n162 VDD2.n128 0.155672
R359 VDD2.n162 VDD2.n161 0.155672
R360 VDD2.n161 VDD2.n132 0.155672
R361 VDD2.n154 VDD2.n132 0.155672
R362 VDD2.n154 VDD2.n153 0.155672
R363 VDD2.n153 VDD2.n137 0.155672
R364 VDD2.n146 VDD2.n137 0.155672
R365 VDD2.n146 VDD2.n145 0.155672
R366 VDD2.n38 VDD2.n37 0.155672
R367 VDD2.n38 VDD2.n29 0.155672
R368 VDD2.n45 VDD2.n29 0.155672
R369 VDD2.n46 VDD2.n45 0.155672
R370 VDD2.n46 VDD2.n25 0.155672
R371 VDD2.n54 VDD2.n25 0.155672
R372 VDD2.n55 VDD2.n54 0.155672
R373 VDD2.n55 VDD2.n21 0.155672
R374 VDD2.n63 VDD2.n21 0.155672
R375 VDD2.n64 VDD2.n63 0.155672
R376 VDD2.n64 VDD2.n17 0.155672
R377 VDD2.n71 VDD2.n17 0.155672
R378 VDD2.n72 VDD2.n71 0.155672
R379 VDD2.n72 VDD2.n13 0.155672
R380 VDD2.n79 VDD2.n13 0.155672
R381 VDD2.n80 VDD2.n79 0.155672
R382 VDD2.n80 VDD2.n9 0.155672
R383 VDD2.n87 VDD2.n9 0.155672
R384 VDD2.n88 VDD2.n87 0.155672
R385 VDD2.n88 VDD2.n5 0.155672
R386 VDD2.n95 VDD2.n5 0.155672
R387 VDD2.n96 VDD2.n95 0.155672
R388 VDD2.n96 VDD2.n1 0.155672
R389 VDD2.n103 VDD2.n1 0.155672
R390 VTAIL.n361 VTAIL.n360 585
R391 VTAIL.n358 VTAIL.n357 585
R392 VTAIL.n367 VTAIL.n366 585
R393 VTAIL.n369 VTAIL.n368 585
R394 VTAIL.n354 VTAIL.n353 585
R395 VTAIL.n375 VTAIL.n374 585
R396 VTAIL.n378 VTAIL.n377 585
R397 VTAIL.n376 VTAIL.n350 585
R398 VTAIL.n383 VTAIL.n349 585
R399 VTAIL.n385 VTAIL.n384 585
R400 VTAIL.n387 VTAIL.n386 585
R401 VTAIL.n346 VTAIL.n345 585
R402 VTAIL.n393 VTAIL.n392 585
R403 VTAIL.n395 VTAIL.n394 585
R404 VTAIL.n342 VTAIL.n341 585
R405 VTAIL.n401 VTAIL.n400 585
R406 VTAIL.n403 VTAIL.n402 585
R407 VTAIL.n338 VTAIL.n337 585
R408 VTAIL.n409 VTAIL.n408 585
R409 VTAIL.n411 VTAIL.n410 585
R410 VTAIL.n334 VTAIL.n333 585
R411 VTAIL.n417 VTAIL.n416 585
R412 VTAIL.n419 VTAIL.n418 585
R413 VTAIL.n330 VTAIL.n329 585
R414 VTAIL.n425 VTAIL.n424 585
R415 VTAIL.n427 VTAIL.n426 585
R416 VTAIL.n37 VTAIL.n36 585
R417 VTAIL.n34 VTAIL.n33 585
R418 VTAIL.n43 VTAIL.n42 585
R419 VTAIL.n45 VTAIL.n44 585
R420 VTAIL.n30 VTAIL.n29 585
R421 VTAIL.n51 VTAIL.n50 585
R422 VTAIL.n54 VTAIL.n53 585
R423 VTAIL.n52 VTAIL.n26 585
R424 VTAIL.n59 VTAIL.n25 585
R425 VTAIL.n61 VTAIL.n60 585
R426 VTAIL.n63 VTAIL.n62 585
R427 VTAIL.n22 VTAIL.n21 585
R428 VTAIL.n69 VTAIL.n68 585
R429 VTAIL.n71 VTAIL.n70 585
R430 VTAIL.n18 VTAIL.n17 585
R431 VTAIL.n77 VTAIL.n76 585
R432 VTAIL.n79 VTAIL.n78 585
R433 VTAIL.n14 VTAIL.n13 585
R434 VTAIL.n85 VTAIL.n84 585
R435 VTAIL.n87 VTAIL.n86 585
R436 VTAIL.n10 VTAIL.n9 585
R437 VTAIL.n93 VTAIL.n92 585
R438 VTAIL.n95 VTAIL.n94 585
R439 VTAIL.n6 VTAIL.n5 585
R440 VTAIL.n101 VTAIL.n100 585
R441 VTAIL.n103 VTAIL.n102 585
R442 VTAIL.n321 VTAIL.n320 585
R443 VTAIL.n319 VTAIL.n318 585
R444 VTAIL.n224 VTAIL.n223 585
R445 VTAIL.n313 VTAIL.n312 585
R446 VTAIL.n311 VTAIL.n310 585
R447 VTAIL.n228 VTAIL.n227 585
R448 VTAIL.n305 VTAIL.n304 585
R449 VTAIL.n303 VTAIL.n302 585
R450 VTAIL.n232 VTAIL.n231 585
R451 VTAIL.n297 VTAIL.n296 585
R452 VTAIL.n295 VTAIL.n294 585
R453 VTAIL.n236 VTAIL.n235 585
R454 VTAIL.n289 VTAIL.n288 585
R455 VTAIL.n287 VTAIL.n286 585
R456 VTAIL.n240 VTAIL.n239 585
R457 VTAIL.n281 VTAIL.n280 585
R458 VTAIL.n279 VTAIL.n278 585
R459 VTAIL.n277 VTAIL.n243 585
R460 VTAIL.n247 VTAIL.n244 585
R461 VTAIL.n272 VTAIL.n271 585
R462 VTAIL.n270 VTAIL.n269 585
R463 VTAIL.n249 VTAIL.n248 585
R464 VTAIL.n264 VTAIL.n263 585
R465 VTAIL.n262 VTAIL.n261 585
R466 VTAIL.n253 VTAIL.n252 585
R467 VTAIL.n256 VTAIL.n255 585
R468 VTAIL.n213 VTAIL.n212 585
R469 VTAIL.n211 VTAIL.n210 585
R470 VTAIL.n116 VTAIL.n115 585
R471 VTAIL.n205 VTAIL.n204 585
R472 VTAIL.n203 VTAIL.n202 585
R473 VTAIL.n120 VTAIL.n119 585
R474 VTAIL.n197 VTAIL.n196 585
R475 VTAIL.n195 VTAIL.n194 585
R476 VTAIL.n124 VTAIL.n123 585
R477 VTAIL.n189 VTAIL.n188 585
R478 VTAIL.n187 VTAIL.n186 585
R479 VTAIL.n128 VTAIL.n127 585
R480 VTAIL.n181 VTAIL.n180 585
R481 VTAIL.n179 VTAIL.n178 585
R482 VTAIL.n132 VTAIL.n131 585
R483 VTAIL.n173 VTAIL.n172 585
R484 VTAIL.n171 VTAIL.n170 585
R485 VTAIL.n169 VTAIL.n135 585
R486 VTAIL.n139 VTAIL.n136 585
R487 VTAIL.n164 VTAIL.n163 585
R488 VTAIL.n162 VTAIL.n161 585
R489 VTAIL.n141 VTAIL.n140 585
R490 VTAIL.n156 VTAIL.n155 585
R491 VTAIL.n154 VTAIL.n153 585
R492 VTAIL.n145 VTAIL.n144 585
R493 VTAIL.n148 VTAIL.n147 585
R494 VTAIL.n426 VTAIL.n326 498.474
R495 VTAIL.n102 VTAIL.n2 498.474
R496 VTAIL.n320 VTAIL.n220 498.474
R497 VTAIL.n212 VTAIL.n112 498.474
R498 VTAIL.t4 VTAIL.n359 329.036
R499 VTAIL.t1 VTAIL.n35 329.036
R500 VTAIL.t0 VTAIL.n254 329.036
R501 VTAIL.t5 VTAIL.n146 329.036
R502 VTAIL.n360 VTAIL.n357 171.744
R503 VTAIL.n367 VTAIL.n357 171.744
R504 VTAIL.n368 VTAIL.n367 171.744
R505 VTAIL.n368 VTAIL.n353 171.744
R506 VTAIL.n375 VTAIL.n353 171.744
R507 VTAIL.n377 VTAIL.n375 171.744
R508 VTAIL.n377 VTAIL.n376 171.744
R509 VTAIL.n376 VTAIL.n349 171.744
R510 VTAIL.n385 VTAIL.n349 171.744
R511 VTAIL.n386 VTAIL.n385 171.744
R512 VTAIL.n386 VTAIL.n345 171.744
R513 VTAIL.n393 VTAIL.n345 171.744
R514 VTAIL.n394 VTAIL.n393 171.744
R515 VTAIL.n394 VTAIL.n341 171.744
R516 VTAIL.n401 VTAIL.n341 171.744
R517 VTAIL.n402 VTAIL.n401 171.744
R518 VTAIL.n402 VTAIL.n337 171.744
R519 VTAIL.n409 VTAIL.n337 171.744
R520 VTAIL.n410 VTAIL.n409 171.744
R521 VTAIL.n410 VTAIL.n333 171.744
R522 VTAIL.n417 VTAIL.n333 171.744
R523 VTAIL.n418 VTAIL.n417 171.744
R524 VTAIL.n418 VTAIL.n329 171.744
R525 VTAIL.n425 VTAIL.n329 171.744
R526 VTAIL.n426 VTAIL.n425 171.744
R527 VTAIL.n36 VTAIL.n33 171.744
R528 VTAIL.n43 VTAIL.n33 171.744
R529 VTAIL.n44 VTAIL.n43 171.744
R530 VTAIL.n44 VTAIL.n29 171.744
R531 VTAIL.n51 VTAIL.n29 171.744
R532 VTAIL.n53 VTAIL.n51 171.744
R533 VTAIL.n53 VTAIL.n52 171.744
R534 VTAIL.n52 VTAIL.n25 171.744
R535 VTAIL.n61 VTAIL.n25 171.744
R536 VTAIL.n62 VTAIL.n61 171.744
R537 VTAIL.n62 VTAIL.n21 171.744
R538 VTAIL.n69 VTAIL.n21 171.744
R539 VTAIL.n70 VTAIL.n69 171.744
R540 VTAIL.n70 VTAIL.n17 171.744
R541 VTAIL.n77 VTAIL.n17 171.744
R542 VTAIL.n78 VTAIL.n77 171.744
R543 VTAIL.n78 VTAIL.n13 171.744
R544 VTAIL.n85 VTAIL.n13 171.744
R545 VTAIL.n86 VTAIL.n85 171.744
R546 VTAIL.n86 VTAIL.n9 171.744
R547 VTAIL.n93 VTAIL.n9 171.744
R548 VTAIL.n94 VTAIL.n93 171.744
R549 VTAIL.n94 VTAIL.n5 171.744
R550 VTAIL.n101 VTAIL.n5 171.744
R551 VTAIL.n102 VTAIL.n101 171.744
R552 VTAIL.n320 VTAIL.n319 171.744
R553 VTAIL.n319 VTAIL.n223 171.744
R554 VTAIL.n312 VTAIL.n223 171.744
R555 VTAIL.n312 VTAIL.n311 171.744
R556 VTAIL.n311 VTAIL.n227 171.744
R557 VTAIL.n304 VTAIL.n227 171.744
R558 VTAIL.n304 VTAIL.n303 171.744
R559 VTAIL.n303 VTAIL.n231 171.744
R560 VTAIL.n296 VTAIL.n231 171.744
R561 VTAIL.n296 VTAIL.n295 171.744
R562 VTAIL.n295 VTAIL.n235 171.744
R563 VTAIL.n288 VTAIL.n235 171.744
R564 VTAIL.n288 VTAIL.n287 171.744
R565 VTAIL.n287 VTAIL.n239 171.744
R566 VTAIL.n280 VTAIL.n239 171.744
R567 VTAIL.n280 VTAIL.n279 171.744
R568 VTAIL.n279 VTAIL.n243 171.744
R569 VTAIL.n247 VTAIL.n243 171.744
R570 VTAIL.n271 VTAIL.n247 171.744
R571 VTAIL.n271 VTAIL.n270 171.744
R572 VTAIL.n270 VTAIL.n248 171.744
R573 VTAIL.n263 VTAIL.n248 171.744
R574 VTAIL.n263 VTAIL.n262 171.744
R575 VTAIL.n262 VTAIL.n252 171.744
R576 VTAIL.n255 VTAIL.n252 171.744
R577 VTAIL.n212 VTAIL.n211 171.744
R578 VTAIL.n211 VTAIL.n115 171.744
R579 VTAIL.n204 VTAIL.n115 171.744
R580 VTAIL.n204 VTAIL.n203 171.744
R581 VTAIL.n203 VTAIL.n119 171.744
R582 VTAIL.n196 VTAIL.n119 171.744
R583 VTAIL.n196 VTAIL.n195 171.744
R584 VTAIL.n195 VTAIL.n123 171.744
R585 VTAIL.n188 VTAIL.n123 171.744
R586 VTAIL.n188 VTAIL.n187 171.744
R587 VTAIL.n187 VTAIL.n127 171.744
R588 VTAIL.n180 VTAIL.n127 171.744
R589 VTAIL.n180 VTAIL.n179 171.744
R590 VTAIL.n179 VTAIL.n131 171.744
R591 VTAIL.n172 VTAIL.n131 171.744
R592 VTAIL.n172 VTAIL.n171 171.744
R593 VTAIL.n171 VTAIL.n135 171.744
R594 VTAIL.n139 VTAIL.n135 171.744
R595 VTAIL.n163 VTAIL.n139 171.744
R596 VTAIL.n163 VTAIL.n162 171.744
R597 VTAIL.n162 VTAIL.n140 171.744
R598 VTAIL.n155 VTAIL.n140 171.744
R599 VTAIL.n155 VTAIL.n154 171.744
R600 VTAIL.n154 VTAIL.n144 171.744
R601 VTAIL.n147 VTAIL.n144 171.744
R602 VTAIL.n360 VTAIL.t4 85.8723
R603 VTAIL.n36 VTAIL.t1 85.8723
R604 VTAIL.n255 VTAIL.t0 85.8723
R605 VTAIL.n147 VTAIL.t5 85.8723
R606 VTAIL.n219 VTAIL.n218 52.9099
R607 VTAIL.n111 VTAIL.n110 52.9099
R608 VTAIL.n1 VTAIL.n0 52.9097
R609 VTAIL.n109 VTAIL.n108 52.9097
R610 VTAIL.n111 VTAIL.n109 35.9445
R611 VTAIL.n431 VTAIL.n430 33.9308
R612 VTAIL.n107 VTAIL.n106 33.9308
R613 VTAIL.n325 VTAIL.n324 33.9308
R614 VTAIL.n217 VTAIL.n216 33.9308
R615 VTAIL.n431 VTAIL.n325 32.5221
R616 VTAIL.n384 VTAIL.n383 13.1884
R617 VTAIL.n60 VTAIL.n59 13.1884
R618 VTAIL.n278 VTAIL.n277 13.1884
R619 VTAIL.n170 VTAIL.n169 13.1884
R620 VTAIL.n382 VTAIL.n350 12.8005
R621 VTAIL.n387 VTAIL.n348 12.8005
R622 VTAIL.n428 VTAIL.n427 12.8005
R623 VTAIL.n58 VTAIL.n26 12.8005
R624 VTAIL.n63 VTAIL.n24 12.8005
R625 VTAIL.n104 VTAIL.n103 12.8005
R626 VTAIL.n322 VTAIL.n321 12.8005
R627 VTAIL.n281 VTAIL.n242 12.8005
R628 VTAIL.n276 VTAIL.n244 12.8005
R629 VTAIL.n214 VTAIL.n213 12.8005
R630 VTAIL.n173 VTAIL.n134 12.8005
R631 VTAIL.n168 VTAIL.n136 12.8005
R632 VTAIL.n379 VTAIL.n378 12.0247
R633 VTAIL.n388 VTAIL.n346 12.0247
R634 VTAIL.n424 VTAIL.n328 12.0247
R635 VTAIL.n55 VTAIL.n54 12.0247
R636 VTAIL.n64 VTAIL.n22 12.0247
R637 VTAIL.n100 VTAIL.n4 12.0247
R638 VTAIL.n318 VTAIL.n222 12.0247
R639 VTAIL.n282 VTAIL.n240 12.0247
R640 VTAIL.n273 VTAIL.n272 12.0247
R641 VTAIL.n210 VTAIL.n114 12.0247
R642 VTAIL.n174 VTAIL.n132 12.0247
R643 VTAIL.n165 VTAIL.n164 12.0247
R644 VTAIL.n374 VTAIL.n352 11.249
R645 VTAIL.n392 VTAIL.n391 11.249
R646 VTAIL.n423 VTAIL.n330 11.249
R647 VTAIL.n50 VTAIL.n28 11.249
R648 VTAIL.n68 VTAIL.n67 11.249
R649 VTAIL.n99 VTAIL.n6 11.249
R650 VTAIL.n317 VTAIL.n224 11.249
R651 VTAIL.n286 VTAIL.n285 11.249
R652 VTAIL.n269 VTAIL.n246 11.249
R653 VTAIL.n209 VTAIL.n116 11.249
R654 VTAIL.n178 VTAIL.n177 11.249
R655 VTAIL.n161 VTAIL.n138 11.249
R656 VTAIL.n361 VTAIL.n359 10.7239
R657 VTAIL.n37 VTAIL.n35 10.7239
R658 VTAIL.n256 VTAIL.n254 10.7239
R659 VTAIL.n148 VTAIL.n146 10.7239
R660 VTAIL.n373 VTAIL.n354 10.4732
R661 VTAIL.n395 VTAIL.n344 10.4732
R662 VTAIL.n420 VTAIL.n419 10.4732
R663 VTAIL.n49 VTAIL.n30 10.4732
R664 VTAIL.n71 VTAIL.n20 10.4732
R665 VTAIL.n96 VTAIL.n95 10.4732
R666 VTAIL.n314 VTAIL.n313 10.4732
R667 VTAIL.n289 VTAIL.n238 10.4732
R668 VTAIL.n268 VTAIL.n249 10.4732
R669 VTAIL.n206 VTAIL.n205 10.4732
R670 VTAIL.n181 VTAIL.n130 10.4732
R671 VTAIL.n160 VTAIL.n141 10.4732
R672 VTAIL.n370 VTAIL.n369 9.69747
R673 VTAIL.n396 VTAIL.n342 9.69747
R674 VTAIL.n416 VTAIL.n332 9.69747
R675 VTAIL.n46 VTAIL.n45 9.69747
R676 VTAIL.n72 VTAIL.n18 9.69747
R677 VTAIL.n92 VTAIL.n8 9.69747
R678 VTAIL.n310 VTAIL.n226 9.69747
R679 VTAIL.n290 VTAIL.n236 9.69747
R680 VTAIL.n265 VTAIL.n264 9.69747
R681 VTAIL.n202 VTAIL.n118 9.69747
R682 VTAIL.n182 VTAIL.n128 9.69747
R683 VTAIL.n157 VTAIL.n156 9.69747
R684 VTAIL.n430 VTAIL.n429 9.45567
R685 VTAIL.n106 VTAIL.n105 9.45567
R686 VTAIL.n324 VTAIL.n323 9.45567
R687 VTAIL.n216 VTAIL.n215 9.45567
R688 VTAIL.n405 VTAIL.n404 9.3005
R689 VTAIL.n340 VTAIL.n339 9.3005
R690 VTAIL.n399 VTAIL.n398 9.3005
R691 VTAIL.n397 VTAIL.n396 9.3005
R692 VTAIL.n344 VTAIL.n343 9.3005
R693 VTAIL.n391 VTAIL.n390 9.3005
R694 VTAIL.n389 VTAIL.n388 9.3005
R695 VTAIL.n348 VTAIL.n347 9.3005
R696 VTAIL.n363 VTAIL.n362 9.3005
R697 VTAIL.n365 VTAIL.n364 9.3005
R698 VTAIL.n356 VTAIL.n355 9.3005
R699 VTAIL.n371 VTAIL.n370 9.3005
R700 VTAIL.n373 VTAIL.n372 9.3005
R701 VTAIL.n352 VTAIL.n351 9.3005
R702 VTAIL.n380 VTAIL.n379 9.3005
R703 VTAIL.n382 VTAIL.n381 9.3005
R704 VTAIL.n407 VTAIL.n406 9.3005
R705 VTAIL.n336 VTAIL.n335 9.3005
R706 VTAIL.n413 VTAIL.n412 9.3005
R707 VTAIL.n415 VTAIL.n414 9.3005
R708 VTAIL.n332 VTAIL.n331 9.3005
R709 VTAIL.n421 VTAIL.n420 9.3005
R710 VTAIL.n423 VTAIL.n422 9.3005
R711 VTAIL.n328 VTAIL.n327 9.3005
R712 VTAIL.n429 VTAIL.n428 9.3005
R713 VTAIL.n81 VTAIL.n80 9.3005
R714 VTAIL.n16 VTAIL.n15 9.3005
R715 VTAIL.n75 VTAIL.n74 9.3005
R716 VTAIL.n73 VTAIL.n72 9.3005
R717 VTAIL.n20 VTAIL.n19 9.3005
R718 VTAIL.n67 VTAIL.n66 9.3005
R719 VTAIL.n65 VTAIL.n64 9.3005
R720 VTAIL.n24 VTAIL.n23 9.3005
R721 VTAIL.n39 VTAIL.n38 9.3005
R722 VTAIL.n41 VTAIL.n40 9.3005
R723 VTAIL.n32 VTAIL.n31 9.3005
R724 VTAIL.n47 VTAIL.n46 9.3005
R725 VTAIL.n49 VTAIL.n48 9.3005
R726 VTAIL.n28 VTAIL.n27 9.3005
R727 VTAIL.n56 VTAIL.n55 9.3005
R728 VTAIL.n58 VTAIL.n57 9.3005
R729 VTAIL.n83 VTAIL.n82 9.3005
R730 VTAIL.n12 VTAIL.n11 9.3005
R731 VTAIL.n89 VTAIL.n88 9.3005
R732 VTAIL.n91 VTAIL.n90 9.3005
R733 VTAIL.n8 VTAIL.n7 9.3005
R734 VTAIL.n97 VTAIL.n96 9.3005
R735 VTAIL.n99 VTAIL.n98 9.3005
R736 VTAIL.n4 VTAIL.n3 9.3005
R737 VTAIL.n105 VTAIL.n104 9.3005
R738 VTAIL.n258 VTAIL.n257 9.3005
R739 VTAIL.n260 VTAIL.n259 9.3005
R740 VTAIL.n251 VTAIL.n250 9.3005
R741 VTAIL.n266 VTAIL.n265 9.3005
R742 VTAIL.n268 VTAIL.n267 9.3005
R743 VTAIL.n246 VTAIL.n245 9.3005
R744 VTAIL.n274 VTAIL.n273 9.3005
R745 VTAIL.n276 VTAIL.n275 9.3005
R746 VTAIL.n230 VTAIL.n229 9.3005
R747 VTAIL.n307 VTAIL.n306 9.3005
R748 VTAIL.n309 VTAIL.n308 9.3005
R749 VTAIL.n226 VTAIL.n225 9.3005
R750 VTAIL.n315 VTAIL.n314 9.3005
R751 VTAIL.n317 VTAIL.n316 9.3005
R752 VTAIL.n222 VTAIL.n221 9.3005
R753 VTAIL.n323 VTAIL.n322 9.3005
R754 VTAIL.n301 VTAIL.n300 9.3005
R755 VTAIL.n299 VTAIL.n298 9.3005
R756 VTAIL.n234 VTAIL.n233 9.3005
R757 VTAIL.n293 VTAIL.n292 9.3005
R758 VTAIL.n291 VTAIL.n290 9.3005
R759 VTAIL.n238 VTAIL.n237 9.3005
R760 VTAIL.n285 VTAIL.n284 9.3005
R761 VTAIL.n283 VTAIL.n282 9.3005
R762 VTAIL.n242 VTAIL.n241 9.3005
R763 VTAIL.n150 VTAIL.n149 9.3005
R764 VTAIL.n152 VTAIL.n151 9.3005
R765 VTAIL.n143 VTAIL.n142 9.3005
R766 VTAIL.n158 VTAIL.n157 9.3005
R767 VTAIL.n160 VTAIL.n159 9.3005
R768 VTAIL.n138 VTAIL.n137 9.3005
R769 VTAIL.n166 VTAIL.n165 9.3005
R770 VTAIL.n168 VTAIL.n167 9.3005
R771 VTAIL.n122 VTAIL.n121 9.3005
R772 VTAIL.n199 VTAIL.n198 9.3005
R773 VTAIL.n201 VTAIL.n200 9.3005
R774 VTAIL.n118 VTAIL.n117 9.3005
R775 VTAIL.n207 VTAIL.n206 9.3005
R776 VTAIL.n209 VTAIL.n208 9.3005
R777 VTAIL.n114 VTAIL.n113 9.3005
R778 VTAIL.n215 VTAIL.n214 9.3005
R779 VTAIL.n193 VTAIL.n192 9.3005
R780 VTAIL.n191 VTAIL.n190 9.3005
R781 VTAIL.n126 VTAIL.n125 9.3005
R782 VTAIL.n185 VTAIL.n184 9.3005
R783 VTAIL.n183 VTAIL.n182 9.3005
R784 VTAIL.n130 VTAIL.n129 9.3005
R785 VTAIL.n177 VTAIL.n176 9.3005
R786 VTAIL.n175 VTAIL.n174 9.3005
R787 VTAIL.n134 VTAIL.n133 9.3005
R788 VTAIL.n366 VTAIL.n356 8.92171
R789 VTAIL.n400 VTAIL.n399 8.92171
R790 VTAIL.n415 VTAIL.n334 8.92171
R791 VTAIL.n42 VTAIL.n32 8.92171
R792 VTAIL.n76 VTAIL.n75 8.92171
R793 VTAIL.n91 VTAIL.n10 8.92171
R794 VTAIL.n309 VTAIL.n228 8.92171
R795 VTAIL.n294 VTAIL.n293 8.92171
R796 VTAIL.n261 VTAIL.n251 8.92171
R797 VTAIL.n201 VTAIL.n120 8.92171
R798 VTAIL.n186 VTAIL.n185 8.92171
R799 VTAIL.n153 VTAIL.n143 8.92171
R800 VTAIL.n365 VTAIL.n358 8.14595
R801 VTAIL.n403 VTAIL.n340 8.14595
R802 VTAIL.n412 VTAIL.n411 8.14595
R803 VTAIL.n41 VTAIL.n34 8.14595
R804 VTAIL.n79 VTAIL.n16 8.14595
R805 VTAIL.n88 VTAIL.n87 8.14595
R806 VTAIL.n306 VTAIL.n305 8.14595
R807 VTAIL.n297 VTAIL.n234 8.14595
R808 VTAIL.n260 VTAIL.n253 8.14595
R809 VTAIL.n198 VTAIL.n197 8.14595
R810 VTAIL.n189 VTAIL.n126 8.14595
R811 VTAIL.n152 VTAIL.n145 8.14595
R812 VTAIL.n430 VTAIL.n326 7.75445
R813 VTAIL.n106 VTAIL.n2 7.75445
R814 VTAIL.n324 VTAIL.n220 7.75445
R815 VTAIL.n216 VTAIL.n112 7.75445
R816 VTAIL.n362 VTAIL.n361 7.3702
R817 VTAIL.n404 VTAIL.n338 7.3702
R818 VTAIL.n408 VTAIL.n336 7.3702
R819 VTAIL.n38 VTAIL.n37 7.3702
R820 VTAIL.n80 VTAIL.n14 7.3702
R821 VTAIL.n84 VTAIL.n12 7.3702
R822 VTAIL.n302 VTAIL.n230 7.3702
R823 VTAIL.n298 VTAIL.n232 7.3702
R824 VTAIL.n257 VTAIL.n256 7.3702
R825 VTAIL.n194 VTAIL.n122 7.3702
R826 VTAIL.n190 VTAIL.n124 7.3702
R827 VTAIL.n149 VTAIL.n148 7.3702
R828 VTAIL.n407 VTAIL.n338 6.59444
R829 VTAIL.n408 VTAIL.n407 6.59444
R830 VTAIL.n83 VTAIL.n14 6.59444
R831 VTAIL.n84 VTAIL.n83 6.59444
R832 VTAIL.n302 VTAIL.n301 6.59444
R833 VTAIL.n301 VTAIL.n232 6.59444
R834 VTAIL.n194 VTAIL.n193 6.59444
R835 VTAIL.n193 VTAIL.n124 6.59444
R836 VTAIL.n428 VTAIL.n326 6.08283
R837 VTAIL.n104 VTAIL.n2 6.08283
R838 VTAIL.n322 VTAIL.n220 6.08283
R839 VTAIL.n214 VTAIL.n112 6.08283
R840 VTAIL.n362 VTAIL.n358 5.81868
R841 VTAIL.n404 VTAIL.n403 5.81868
R842 VTAIL.n411 VTAIL.n336 5.81868
R843 VTAIL.n38 VTAIL.n34 5.81868
R844 VTAIL.n80 VTAIL.n79 5.81868
R845 VTAIL.n87 VTAIL.n12 5.81868
R846 VTAIL.n305 VTAIL.n230 5.81868
R847 VTAIL.n298 VTAIL.n297 5.81868
R848 VTAIL.n257 VTAIL.n253 5.81868
R849 VTAIL.n197 VTAIL.n122 5.81868
R850 VTAIL.n190 VTAIL.n189 5.81868
R851 VTAIL.n149 VTAIL.n145 5.81868
R852 VTAIL.n366 VTAIL.n365 5.04292
R853 VTAIL.n400 VTAIL.n340 5.04292
R854 VTAIL.n412 VTAIL.n334 5.04292
R855 VTAIL.n42 VTAIL.n41 5.04292
R856 VTAIL.n76 VTAIL.n16 5.04292
R857 VTAIL.n88 VTAIL.n10 5.04292
R858 VTAIL.n306 VTAIL.n228 5.04292
R859 VTAIL.n294 VTAIL.n234 5.04292
R860 VTAIL.n261 VTAIL.n260 5.04292
R861 VTAIL.n198 VTAIL.n120 5.04292
R862 VTAIL.n186 VTAIL.n126 5.04292
R863 VTAIL.n153 VTAIL.n152 5.04292
R864 VTAIL.n369 VTAIL.n356 4.26717
R865 VTAIL.n399 VTAIL.n342 4.26717
R866 VTAIL.n416 VTAIL.n415 4.26717
R867 VTAIL.n45 VTAIL.n32 4.26717
R868 VTAIL.n75 VTAIL.n18 4.26717
R869 VTAIL.n92 VTAIL.n91 4.26717
R870 VTAIL.n310 VTAIL.n309 4.26717
R871 VTAIL.n293 VTAIL.n236 4.26717
R872 VTAIL.n264 VTAIL.n251 4.26717
R873 VTAIL.n202 VTAIL.n201 4.26717
R874 VTAIL.n185 VTAIL.n128 4.26717
R875 VTAIL.n156 VTAIL.n143 4.26717
R876 VTAIL.n370 VTAIL.n354 3.49141
R877 VTAIL.n396 VTAIL.n395 3.49141
R878 VTAIL.n419 VTAIL.n332 3.49141
R879 VTAIL.n46 VTAIL.n30 3.49141
R880 VTAIL.n72 VTAIL.n71 3.49141
R881 VTAIL.n95 VTAIL.n8 3.49141
R882 VTAIL.n313 VTAIL.n226 3.49141
R883 VTAIL.n290 VTAIL.n289 3.49141
R884 VTAIL.n265 VTAIL.n249 3.49141
R885 VTAIL.n205 VTAIL.n118 3.49141
R886 VTAIL.n182 VTAIL.n181 3.49141
R887 VTAIL.n157 VTAIL.n141 3.49141
R888 VTAIL.n217 VTAIL.n111 3.42291
R889 VTAIL.n325 VTAIL.n219 3.42291
R890 VTAIL.n109 VTAIL.n107 3.42291
R891 VTAIL.n374 VTAIL.n373 2.71565
R892 VTAIL.n392 VTAIL.n344 2.71565
R893 VTAIL.n420 VTAIL.n330 2.71565
R894 VTAIL.n50 VTAIL.n49 2.71565
R895 VTAIL.n68 VTAIL.n20 2.71565
R896 VTAIL.n96 VTAIL.n6 2.71565
R897 VTAIL.n314 VTAIL.n224 2.71565
R898 VTAIL.n286 VTAIL.n238 2.71565
R899 VTAIL.n269 VTAIL.n268 2.71565
R900 VTAIL.n206 VTAIL.n116 2.71565
R901 VTAIL.n178 VTAIL.n130 2.71565
R902 VTAIL.n161 VTAIL.n160 2.71565
R903 VTAIL VTAIL.n431 2.50912
R904 VTAIL.n258 VTAIL.n254 2.41282
R905 VTAIL.n150 VTAIL.n146 2.41282
R906 VTAIL.n363 VTAIL.n359 2.41282
R907 VTAIL.n39 VTAIL.n35 2.41282
R908 VTAIL.n219 VTAIL.n217 2.18153
R909 VTAIL.n107 VTAIL.n1 2.18153
R910 VTAIL.n378 VTAIL.n352 1.93989
R911 VTAIL.n391 VTAIL.n346 1.93989
R912 VTAIL.n424 VTAIL.n423 1.93989
R913 VTAIL.n54 VTAIL.n28 1.93989
R914 VTAIL.n67 VTAIL.n22 1.93989
R915 VTAIL.n100 VTAIL.n99 1.93989
R916 VTAIL.n318 VTAIL.n317 1.93989
R917 VTAIL.n285 VTAIL.n240 1.93989
R918 VTAIL.n272 VTAIL.n246 1.93989
R919 VTAIL.n210 VTAIL.n209 1.93989
R920 VTAIL.n177 VTAIL.n132 1.93989
R921 VTAIL.n164 VTAIL.n138 1.93989
R922 VTAIL.n0 VTAIL.t7 1.67515
R923 VTAIL.n0 VTAIL.t6 1.67515
R924 VTAIL.n108 VTAIL.t10 1.67515
R925 VTAIL.n108 VTAIL.t9 1.67515
R926 VTAIL.n218 VTAIL.t2 1.67515
R927 VTAIL.n218 VTAIL.t11 1.67515
R928 VTAIL.n110 VTAIL.t3 1.67515
R929 VTAIL.n110 VTAIL.t8 1.67515
R930 VTAIL.n379 VTAIL.n350 1.16414
R931 VTAIL.n388 VTAIL.n387 1.16414
R932 VTAIL.n427 VTAIL.n328 1.16414
R933 VTAIL.n55 VTAIL.n26 1.16414
R934 VTAIL.n64 VTAIL.n63 1.16414
R935 VTAIL.n103 VTAIL.n4 1.16414
R936 VTAIL.n321 VTAIL.n222 1.16414
R937 VTAIL.n282 VTAIL.n281 1.16414
R938 VTAIL.n273 VTAIL.n244 1.16414
R939 VTAIL.n213 VTAIL.n114 1.16414
R940 VTAIL.n174 VTAIL.n173 1.16414
R941 VTAIL.n165 VTAIL.n136 1.16414
R942 VTAIL VTAIL.n1 0.914293
R943 VTAIL.n383 VTAIL.n382 0.388379
R944 VTAIL.n384 VTAIL.n348 0.388379
R945 VTAIL.n59 VTAIL.n58 0.388379
R946 VTAIL.n60 VTAIL.n24 0.388379
R947 VTAIL.n278 VTAIL.n242 0.388379
R948 VTAIL.n277 VTAIL.n276 0.388379
R949 VTAIL.n170 VTAIL.n134 0.388379
R950 VTAIL.n169 VTAIL.n168 0.388379
R951 VTAIL.n364 VTAIL.n363 0.155672
R952 VTAIL.n364 VTAIL.n355 0.155672
R953 VTAIL.n371 VTAIL.n355 0.155672
R954 VTAIL.n372 VTAIL.n371 0.155672
R955 VTAIL.n372 VTAIL.n351 0.155672
R956 VTAIL.n380 VTAIL.n351 0.155672
R957 VTAIL.n381 VTAIL.n380 0.155672
R958 VTAIL.n381 VTAIL.n347 0.155672
R959 VTAIL.n389 VTAIL.n347 0.155672
R960 VTAIL.n390 VTAIL.n389 0.155672
R961 VTAIL.n390 VTAIL.n343 0.155672
R962 VTAIL.n397 VTAIL.n343 0.155672
R963 VTAIL.n398 VTAIL.n397 0.155672
R964 VTAIL.n398 VTAIL.n339 0.155672
R965 VTAIL.n405 VTAIL.n339 0.155672
R966 VTAIL.n406 VTAIL.n405 0.155672
R967 VTAIL.n406 VTAIL.n335 0.155672
R968 VTAIL.n413 VTAIL.n335 0.155672
R969 VTAIL.n414 VTAIL.n413 0.155672
R970 VTAIL.n414 VTAIL.n331 0.155672
R971 VTAIL.n421 VTAIL.n331 0.155672
R972 VTAIL.n422 VTAIL.n421 0.155672
R973 VTAIL.n422 VTAIL.n327 0.155672
R974 VTAIL.n429 VTAIL.n327 0.155672
R975 VTAIL.n40 VTAIL.n39 0.155672
R976 VTAIL.n40 VTAIL.n31 0.155672
R977 VTAIL.n47 VTAIL.n31 0.155672
R978 VTAIL.n48 VTAIL.n47 0.155672
R979 VTAIL.n48 VTAIL.n27 0.155672
R980 VTAIL.n56 VTAIL.n27 0.155672
R981 VTAIL.n57 VTAIL.n56 0.155672
R982 VTAIL.n57 VTAIL.n23 0.155672
R983 VTAIL.n65 VTAIL.n23 0.155672
R984 VTAIL.n66 VTAIL.n65 0.155672
R985 VTAIL.n66 VTAIL.n19 0.155672
R986 VTAIL.n73 VTAIL.n19 0.155672
R987 VTAIL.n74 VTAIL.n73 0.155672
R988 VTAIL.n74 VTAIL.n15 0.155672
R989 VTAIL.n81 VTAIL.n15 0.155672
R990 VTAIL.n82 VTAIL.n81 0.155672
R991 VTAIL.n82 VTAIL.n11 0.155672
R992 VTAIL.n89 VTAIL.n11 0.155672
R993 VTAIL.n90 VTAIL.n89 0.155672
R994 VTAIL.n90 VTAIL.n7 0.155672
R995 VTAIL.n97 VTAIL.n7 0.155672
R996 VTAIL.n98 VTAIL.n97 0.155672
R997 VTAIL.n98 VTAIL.n3 0.155672
R998 VTAIL.n105 VTAIL.n3 0.155672
R999 VTAIL.n323 VTAIL.n221 0.155672
R1000 VTAIL.n316 VTAIL.n221 0.155672
R1001 VTAIL.n316 VTAIL.n315 0.155672
R1002 VTAIL.n315 VTAIL.n225 0.155672
R1003 VTAIL.n308 VTAIL.n225 0.155672
R1004 VTAIL.n308 VTAIL.n307 0.155672
R1005 VTAIL.n307 VTAIL.n229 0.155672
R1006 VTAIL.n300 VTAIL.n229 0.155672
R1007 VTAIL.n300 VTAIL.n299 0.155672
R1008 VTAIL.n299 VTAIL.n233 0.155672
R1009 VTAIL.n292 VTAIL.n233 0.155672
R1010 VTAIL.n292 VTAIL.n291 0.155672
R1011 VTAIL.n291 VTAIL.n237 0.155672
R1012 VTAIL.n284 VTAIL.n237 0.155672
R1013 VTAIL.n284 VTAIL.n283 0.155672
R1014 VTAIL.n283 VTAIL.n241 0.155672
R1015 VTAIL.n275 VTAIL.n241 0.155672
R1016 VTAIL.n275 VTAIL.n274 0.155672
R1017 VTAIL.n274 VTAIL.n245 0.155672
R1018 VTAIL.n267 VTAIL.n245 0.155672
R1019 VTAIL.n267 VTAIL.n266 0.155672
R1020 VTAIL.n266 VTAIL.n250 0.155672
R1021 VTAIL.n259 VTAIL.n250 0.155672
R1022 VTAIL.n259 VTAIL.n258 0.155672
R1023 VTAIL.n215 VTAIL.n113 0.155672
R1024 VTAIL.n208 VTAIL.n113 0.155672
R1025 VTAIL.n208 VTAIL.n207 0.155672
R1026 VTAIL.n207 VTAIL.n117 0.155672
R1027 VTAIL.n200 VTAIL.n117 0.155672
R1028 VTAIL.n200 VTAIL.n199 0.155672
R1029 VTAIL.n199 VTAIL.n121 0.155672
R1030 VTAIL.n192 VTAIL.n121 0.155672
R1031 VTAIL.n192 VTAIL.n191 0.155672
R1032 VTAIL.n191 VTAIL.n125 0.155672
R1033 VTAIL.n184 VTAIL.n125 0.155672
R1034 VTAIL.n184 VTAIL.n183 0.155672
R1035 VTAIL.n183 VTAIL.n129 0.155672
R1036 VTAIL.n176 VTAIL.n129 0.155672
R1037 VTAIL.n176 VTAIL.n175 0.155672
R1038 VTAIL.n175 VTAIL.n133 0.155672
R1039 VTAIL.n167 VTAIL.n133 0.155672
R1040 VTAIL.n167 VTAIL.n166 0.155672
R1041 VTAIL.n166 VTAIL.n137 0.155672
R1042 VTAIL.n159 VTAIL.n137 0.155672
R1043 VTAIL.n159 VTAIL.n158 0.155672
R1044 VTAIL.n158 VTAIL.n142 0.155672
R1045 VTAIL.n151 VTAIL.n142 0.155672
R1046 VTAIL.n151 VTAIL.n150 0.155672
R1047 VP.n15 VP.t0 162.023
R1048 VP.n16 VP.n13 161.3
R1049 VP.n18 VP.n17 161.3
R1050 VP.n19 VP.n12 161.3
R1051 VP.n21 VP.n20 161.3
R1052 VP.n22 VP.n11 161.3
R1053 VP.n24 VP.n23 161.3
R1054 VP.n25 VP.n10 161.3
R1055 VP.n27 VP.n26 161.3
R1056 VP.n55 VP.n54 161.3
R1057 VP.n53 VP.n1 161.3
R1058 VP.n52 VP.n51 161.3
R1059 VP.n50 VP.n2 161.3
R1060 VP.n49 VP.n48 161.3
R1061 VP.n47 VP.n3 161.3
R1062 VP.n46 VP.n45 161.3
R1063 VP.n44 VP.n4 161.3
R1064 VP.n43 VP.n42 161.3
R1065 VP.n40 VP.n5 161.3
R1066 VP.n39 VP.n38 161.3
R1067 VP.n37 VP.n6 161.3
R1068 VP.n36 VP.n35 161.3
R1069 VP.n34 VP.n7 161.3
R1070 VP.n33 VP.n32 161.3
R1071 VP.n31 VP.n8 161.3
R1072 VP.n29 VP.t3 128.512
R1073 VP.n41 VP.t4 128.512
R1074 VP.n0 VP.t1 128.512
R1075 VP.n9 VP.t5 128.512
R1076 VP.n14 VP.t2 128.512
R1077 VP.n30 VP.n29 79.3019
R1078 VP.n56 VP.n0 79.3019
R1079 VP.n28 VP.n9 79.3019
R1080 VP.n15 VP.n14 62.396
R1081 VP.n30 VP.n28 58.5031
R1082 VP.n35 VP.n6 56.5193
R1083 VP.n48 VP.n2 56.5193
R1084 VP.n20 VP.n11 56.5193
R1085 VP.n33 VP.n8 24.4675
R1086 VP.n34 VP.n33 24.4675
R1087 VP.n35 VP.n34 24.4675
R1088 VP.n39 VP.n6 24.4675
R1089 VP.n40 VP.n39 24.4675
R1090 VP.n42 VP.n40 24.4675
R1091 VP.n46 VP.n4 24.4675
R1092 VP.n47 VP.n46 24.4675
R1093 VP.n48 VP.n47 24.4675
R1094 VP.n52 VP.n2 24.4675
R1095 VP.n53 VP.n52 24.4675
R1096 VP.n54 VP.n53 24.4675
R1097 VP.n24 VP.n11 24.4675
R1098 VP.n25 VP.n24 24.4675
R1099 VP.n26 VP.n25 24.4675
R1100 VP.n18 VP.n13 24.4675
R1101 VP.n19 VP.n18 24.4675
R1102 VP.n20 VP.n19 24.4675
R1103 VP.n42 VP.n41 12.234
R1104 VP.n41 VP.n4 12.234
R1105 VP.n14 VP.n13 12.234
R1106 VP.n29 VP.n8 10.766
R1107 VP.n54 VP.n0 10.766
R1108 VP.n26 VP.n9 10.766
R1109 VP.n16 VP.n15 3.13204
R1110 VP.n28 VP.n27 0.354971
R1111 VP.n31 VP.n30 0.354971
R1112 VP.n56 VP.n55 0.354971
R1113 VP VP.n56 0.26696
R1114 VP.n17 VP.n16 0.189894
R1115 VP.n17 VP.n12 0.189894
R1116 VP.n21 VP.n12 0.189894
R1117 VP.n22 VP.n21 0.189894
R1118 VP.n23 VP.n22 0.189894
R1119 VP.n23 VP.n10 0.189894
R1120 VP.n27 VP.n10 0.189894
R1121 VP.n32 VP.n31 0.189894
R1122 VP.n32 VP.n7 0.189894
R1123 VP.n36 VP.n7 0.189894
R1124 VP.n37 VP.n36 0.189894
R1125 VP.n38 VP.n37 0.189894
R1126 VP.n38 VP.n5 0.189894
R1127 VP.n43 VP.n5 0.189894
R1128 VP.n44 VP.n43 0.189894
R1129 VP.n45 VP.n44 0.189894
R1130 VP.n45 VP.n3 0.189894
R1131 VP.n49 VP.n3 0.189894
R1132 VP.n50 VP.n49 0.189894
R1133 VP.n51 VP.n50 0.189894
R1134 VP.n51 VP.n1 0.189894
R1135 VP.n55 VP.n1 0.189894
R1136 VDD1.n101 VDD1.n100 585
R1137 VDD1.n99 VDD1.n98 585
R1138 VDD1.n4 VDD1.n3 585
R1139 VDD1.n93 VDD1.n92 585
R1140 VDD1.n91 VDD1.n90 585
R1141 VDD1.n8 VDD1.n7 585
R1142 VDD1.n85 VDD1.n84 585
R1143 VDD1.n83 VDD1.n82 585
R1144 VDD1.n12 VDD1.n11 585
R1145 VDD1.n77 VDD1.n76 585
R1146 VDD1.n75 VDD1.n74 585
R1147 VDD1.n16 VDD1.n15 585
R1148 VDD1.n69 VDD1.n68 585
R1149 VDD1.n67 VDD1.n66 585
R1150 VDD1.n20 VDD1.n19 585
R1151 VDD1.n61 VDD1.n60 585
R1152 VDD1.n59 VDD1.n58 585
R1153 VDD1.n57 VDD1.n23 585
R1154 VDD1.n27 VDD1.n24 585
R1155 VDD1.n52 VDD1.n51 585
R1156 VDD1.n50 VDD1.n49 585
R1157 VDD1.n29 VDD1.n28 585
R1158 VDD1.n44 VDD1.n43 585
R1159 VDD1.n42 VDD1.n41 585
R1160 VDD1.n33 VDD1.n32 585
R1161 VDD1.n36 VDD1.n35 585
R1162 VDD1.n140 VDD1.n139 585
R1163 VDD1.n137 VDD1.n136 585
R1164 VDD1.n146 VDD1.n145 585
R1165 VDD1.n148 VDD1.n147 585
R1166 VDD1.n133 VDD1.n132 585
R1167 VDD1.n154 VDD1.n153 585
R1168 VDD1.n157 VDD1.n156 585
R1169 VDD1.n155 VDD1.n129 585
R1170 VDD1.n162 VDD1.n128 585
R1171 VDD1.n164 VDD1.n163 585
R1172 VDD1.n166 VDD1.n165 585
R1173 VDD1.n125 VDD1.n124 585
R1174 VDD1.n172 VDD1.n171 585
R1175 VDD1.n174 VDD1.n173 585
R1176 VDD1.n121 VDD1.n120 585
R1177 VDD1.n180 VDD1.n179 585
R1178 VDD1.n182 VDD1.n181 585
R1179 VDD1.n117 VDD1.n116 585
R1180 VDD1.n188 VDD1.n187 585
R1181 VDD1.n190 VDD1.n189 585
R1182 VDD1.n113 VDD1.n112 585
R1183 VDD1.n196 VDD1.n195 585
R1184 VDD1.n198 VDD1.n197 585
R1185 VDD1.n109 VDD1.n108 585
R1186 VDD1.n204 VDD1.n203 585
R1187 VDD1.n206 VDD1.n205 585
R1188 VDD1.n100 VDD1.n0 498.474
R1189 VDD1.n205 VDD1.n105 498.474
R1190 VDD1.t5 VDD1.n34 329.036
R1191 VDD1.t2 VDD1.n138 329.036
R1192 VDD1.n100 VDD1.n99 171.744
R1193 VDD1.n99 VDD1.n3 171.744
R1194 VDD1.n92 VDD1.n3 171.744
R1195 VDD1.n92 VDD1.n91 171.744
R1196 VDD1.n91 VDD1.n7 171.744
R1197 VDD1.n84 VDD1.n7 171.744
R1198 VDD1.n84 VDD1.n83 171.744
R1199 VDD1.n83 VDD1.n11 171.744
R1200 VDD1.n76 VDD1.n11 171.744
R1201 VDD1.n76 VDD1.n75 171.744
R1202 VDD1.n75 VDD1.n15 171.744
R1203 VDD1.n68 VDD1.n15 171.744
R1204 VDD1.n68 VDD1.n67 171.744
R1205 VDD1.n67 VDD1.n19 171.744
R1206 VDD1.n60 VDD1.n19 171.744
R1207 VDD1.n60 VDD1.n59 171.744
R1208 VDD1.n59 VDD1.n23 171.744
R1209 VDD1.n27 VDD1.n23 171.744
R1210 VDD1.n51 VDD1.n27 171.744
R1211 VDD1.n51 VDD1.n50 171.744
R1212 VDD1.n50 VDD1.n28 171.744
R1213 VDD1.n43 VDD1.n28 171.744
R1214 VDD1.n43 VDD1.n42 171.744
R1215 VDD1.n42 VDD1.n32 171.744
R1216 VDD1.n35 VDD1.n32 171.744
R1217 VDD1.n139 VDD1.n136 171.744
R1218 VDD1.n146 VDD1.n136 171.744
R1219 VDD1.n147 VDD1.n146 171.744
R1220 VDD1.n147 VDD1.n132 171.744
R1221 VDD1.n154 VDD1.n132 171.744
R1222 VDD1.n156 VDD1.n154 171.744
R1223 VDD1.n156 VDD1.n155 171.744
R1224 VDD1.n155 VDD1.n128 171.744
R1225 VDD1.n164 VDD1.n128 171.744
R1226 VDD1.n165 VDD1.n164 171.744
R1227 VDD1.n165 VDD1.n124 171.744
R1228 VDD1.n172 VDD1.n124 171.744
R1229 VDD1.n173 VDD1.n172 171.744
R1230 VDD1.n173 VDD1.n120 171.744
R1231 VDD1.n180 VDD1.n120 171.744
R1232 VDD1.n181 VDD1.n180 171.744
R1233 VDD1.n181 VDD1.n116 171.744
R1234 VDD1.n188 VDD1.n116 171.744
R1235 VDD1.n189 VDD1.n188 171.744
R1236 VDD1.n189 VDD1.n112 171.744
R1237 VDD1.n196 VDD1.n112 171.744
R1238 VDD1.n197 VDD1.n196 171.744
R1239 VDD1.n197 VDD1.n108 171.744
R1240 VDD1.n204 VDD1.n108 171.744
R1241 VDD1.n205 VDD1.n204 171.744
R1242 VDD1.n35 VDD1.t5 85.8723
R1243 VDD1.n139 VDD1.t2 85.8723
R1244 VDD1.n211 VDD1.n210 70.3888
R1245 VDD1.n213 VDD1.n212 69.5885
R1246 VDD1.n213 VDD1.n211 53.8651
R1247 VDD1 VDD1.n104 53.2346
R1248 VDD1.n211 VDD1.n209 53.1211
R1249 VDD1.n58 VDD1.n57 13.1884
R1250 VDD1.n163 VDD1.n162 13.1884
R1251 VDD1.n102 VDD1.n101 12.8005
R1252 VDD1.n61 VDD1.n22 12.8005
R1253 VDD1.n56 VDD1.n24 12.8005
R1254 VDD1.n161 VDD1.n129 12.8005
R1255 VDD1.n166 VDD1.n127 12.8005
R1256 VDD1.n207 VDD1.n206 12.8005
R1257 VDD1.n98 VDD1.n2 12.0247
R1258 VDD1.n62 VDD1.n20 12.0247
R1259 VDD1.n53 VDD1.n52 12.0247
R1260 VDD1.n158 VDD1.n157 12.0247
R1261 VDD1.n167 VDD1.n125 12.0247
R1262 VDD1.n203 VDD1.n107 12.0247
R1263 VDD1.n97 VDD1.n4 11.249
R1264 VDD1.n66 VDD1.n65 11.249
R1265 VDD1.n49 VDD1.n26 11.249
R1266 VDD1.n153 VDD1.n131 11.249
R1267 VDD1.n171 VDD1.n170 11.249
R1268 VDD1.n202 VDD1.n109 11.249
R1269 VDD1.n36 VDD1.n34 10.7239
R1270 VDD1.n140 VDD1.n138 10.7239
R1271 VDD1.n94 VDD1.n93 10.4732
R1272 VDD1.n69 VDD1.n18 10.4732
R1273 VDD1.n48 VDD1.n29 10.4732
R1274 VDD1.n152 VDD1.n133 10.4732
R1275 VDD1.n174 VDD1.n123 10.4732
R1276 VDD1.n199 VDD1.n198 10.4732
R1277 VDD1.n90 VDD1.n6 9.69747
R1278 VDD1.n70 VDD1.n16 9.69747
R1279 VDD1.n45 VDD1.n44 9.69747
R1280 VDD1.n149 VDD1.n148 9.69747
R1281 VDD1.n175 VDD1.n121 9.69747
R1282 VDD1.n195 VDD1.n111 9.69747
R1283 VDD1.n104 VDD1.n103 9.45567
R1284 VDD1.n209 VDD1.n208 9.45567
R1285 VDD1.n38 VDD1.n37 9.3005
R1286 VDD1.n40 VDD1.n39 9.3005
R1287 VDD1.n31 VDD1.n30 9.3005
R1288 VDD1.n46 VDD1.n45 9.3005
R1289 VDD1.n48 VDD1.n47 9.3005
R1290 VDD1.n26 VDD1.n25 9.3005
R1291 VDD1.n54 VDD1.n53 9.3005
R1292 VDD1.n56 VDD1.n55 9.3005
R1293 VDD1.n10 VDD1.n9 9.3005
R1294 VDD1.n87 VDD1.n86 9.3005
R1295 VDD1.n89 VDD1.n88 9.3005
R1296 VDD1.n6 VDD1.n5 9.3005
R1297 VDD1.n95 VDD1.n94 9.3005
R1298 VDD1.n97 VDD1.n96 9.3005
R1299 VDD1.n2 VDD1.n1 9.3005
R1300 VDD1.n103 VDD1.n102 9.3005
R1301 VDD1.n81 VDD1.n80 9.3005
R1302 VDD1.n79 VDD1.n78 9.3005
R1303 VDD1.n14 VDD1.n13 9.3005
R1304 VDD1.n73 VDD1.n72 9.3005
R1305 VDD1.n71 VDD1.n70 9.3005
R1306 VDD1.n18 VDD1.n17 9.3005
R1307 VDD1.n65 VDD1.n64 9.3005
R1308 VDD1.n63 VDD1.n62 9.3005
R1309 VDD1.n22 VDD1.n21 9.3005
R1310 VDD1.n184 VDD1.n183 9.3005
R1311 VDD1.n119 VDD1.n118 9.3005
R1312 VDD1.n178 VDD1.n177 9.3005
R1313 VDD1.n176 VDD1.n175 9.3005
R1314 VDD1.n123 VDD1.n122 9.3005
R1315 VDD1.n170 VDD1.n169 9.3005
R1316 VDD1.n168 VDD1.n167 9.3005
R1317 VDD1.n127 VDD1.n126 9.3005
R1318 VDD1.n142 VDD1.n141 9.3005
R1319 VDD1.n144 VDD1.n143 9.3005
R1320 VDD1.n135 VDD1.n134 9.3005
R1321 VDD1.n150 VDD1.n149 9.3005
R1322 VDD1.n152 VDD1.n151 9.3005
R1323 VDD1.n131 VDD1.n130 9.3005
R1324 VDD1.n159 VDD1.n158 9.3005
R1325 VDD1.n161 VDD1.n160 9.3005
R1326 VDD1.n186 VDD1.n185 9.3005
R1327 VDD1.n115 VDD1.n114 9.3005
R1328 VDD1.n192 VDD1.n191 9.3005
R1329 VDD1.n194 VDD1.n193 9.3005
R1330 VDD1.n111 VDD1.n110 9.3005
R1331 VDD1.n200 VDD1.n199 9.3005
R1332 VDD1.n202 VDD1.n201 9.3005
R1333 VDD1.n107 VDD1.n106 9.3005
R1334 VDD1.n208 VDD1.n207 9.3005
R1335 VDD1.n89 VDD1.n8 8.92171
R1336 VDD1.n74 VDD1.n73 8.92171
R1337 VDD1.n41 VDD1.n31 8.92171
R1338 VDD1.n145 VDD1.n135 8.92171
R1339 VDD1.n179 VDD1.n178 8.92171
R1340 VDD1.n194 VDD1.n113 8.92171
R1341 VDD1.n86 VDD1.n85 8.14595
R1342 VDD1.n77 VDD1.n14 8.14595
R1343 VDD1.n40 VDD1.n33 8.14595
R1344 VDD1.n144 VDD1.n137 8.14595
R1345 VDD1.n182 VDD1.n119 8.14595
R1346 VDD1.n191 VDD1.n190 8.14595
R1347 VDD1.n104 VDD1.n0 7.75445
R1348 VDD1.n209 VDD1.n105 7.75445
R1349 VDD1.n82 VDD1.n10 7.3702
R1350 VDD1.n78 VDD1.n12 7.3702
R1351 VDD1.n37 VDD1.n36 7.3702
R1352 VDD1.n141 VDD1.n140 7.3702
R1353 VDD1.n183 VDD1.n117 7.3702
R1354 VDD1.n187 VDD1.n115 7.3702
R1355 VDD1.n82 VDD1.n81 6.59444
R1356 VDD1.n81 VDD1.n12 6.59444
R1357 VDD1.n186 VDD1.n117 6.59444
R1358 VDD1.n187 VDD1.n186 6.59444
R1359 VDD1.n102 VDD1.n0 6.08283
R1360 VDD1.n207 VDD1.n105 6.08283
R1361 VDD1.n85 VDD1.n10 5.81868
R1362 VDD1.n78 VDD1.n77 5.81868
R1363 VDD1.n37 VDD1.n33 5.81868
R1364 VDD1.n141 VDD1.n137 5.81868
R1365 VDD1.n183 VDD1.n182 5.81868
R1366 VDD1.n190 VDD1.n115 5.81868
R1367 VDD1.n86 VDD1.n8 5.04292
R1368 VDD1.n74 VDD1.n14 5.04292
R1369 VDD1.n41 VDD1.n40 5.04292
R1370 VDD1.n145 VDD1.n144 5.04292
R1371 VDD1.n179 VDD1.n119 5.04292
R1372 VDD1.n191 VDD1.n113 5.04292
R1373 VDD1.n90 VDD1.n89 4.26717
R1374 VDD1.n73 VDD1.n16 4.26717
R1375 VDD1.n44 VDD1.n31 4.26717
R1376 VDD1.n148 VDD1.n135 4.26717
R1377 VDD1.n178 VDD1.n121 4.26717
R1378 VDD1.n195 VDD1.n194 4.26717
R1379 VDD1.n93 VDD1.n6 3.49141
R1380 VDD1.n70 VDD1.n69 3.49141
R1381 VDD1.n45 VDD1.n29 3.49141
R1382 VDD1.n149 VDD1.n133 3.49141
R1383 VDD1.n175 VDD1.n174 3.49141
R1384 VDD1.n198 VDD1.n111 3.49141
R1385 VDD1.n94 VDD1.n4 2.71565
R1386 VDD1.n66 VDD1.n18 2.71565
R1387 VDD1.n49 VDD1.n48 2.71565
R1388 VDD1.n153 VDD1.n152 2.71565
R1389 VDD1.n171 VDD1.n123 2.71565
R1390 VDD1.n199 VDD1.n109 2.71565
R1391 VDD1.n38 VDD1.n34 2.41282
R1392 VDD1.n142 VDD1.n138 2.41282
R1393 VDD1.n98 VDD1.n97 1.93989
R1394 VDD1.n65 VDD1.n20 1.93989
R1395 VDD1.n52 VDD1.n26 1.93989
R1396 VDD1.n157 VDD1.n131 1.93989
R1397 VDD1.n170 VDD1.n125 1.93989
R1398 VDD1.n203 VDD1.n202 1.93989
R1399 VDD1.n212 VDD1.t3 1.67515
R1400 VDD1.n212 VDD1.t0 1.67515
R1401 VDD1.n210 VDD1.t1 1.67515
R1402 VDD1.n210 VDD1.t4 1.67515
R1403 VDD1.n101 VDD1.n2 1.16414
R1404 VDD1.n62 VDD1.n61 1.16414
R1405 VDD1.n53 VDD1.n24 1.16414
R1406 VDD1.n158 VDD1.n129 1.16414
R1407 VDD1.n167 VDD1.n166 1.16414
R1408 VDD1.n206 VDD1.n107 1.16414
R1409 VDD1 VDD1.n213 0.797914
R1410 VDD1.n58 VDD1.n22 0.388379
R1411 VDD1.n57 VDD1.n56 0.388379
R1412 VDD1.n162 VDD1.n161 0.388379
R1413 VDD1.n163 VDD1.n127 0.388379
R1414 VDD1.n103 VDD1.n1 0.155672
R1415 VDD1.n96 VDD1.n1 0.155672
R1416 VDD1.n96 VDD1.n95 0.155672
R1417 VDD1.n95 VDD1.n5 0.155672
R1418 VDD1.n88 VDD1.n5 0.155672
R1419 VDD1.n88 VDD1.n87 0.155672
R1420 VDD1.n87 VDD1.n9 0.155672
R1421 VDD1.n80 VDD1.n9 0.155672
R1422 VDD1.n80 VDD1.n79 0.155672
R1423 VDD1.n79 VDD1.n13 0.155672
R1424 VDD1.n72 VDD1.n13 0.155672
R1425 VDD1.n72 VDD1.n71 0.155672
R1426 VDD1.n71 VDD1.n17 0.155672
R1427 VDD1.n64 VDD1.n17 0.155672
R1428 VDD1.n64 VDD1.n63 0.155672
R1429 VDD1.n63 VDD1.n21 0.155672
R1430 VDD1.n55 VDD1.n21 0.155672
R1431 VDD1.n55 VDD1.n54 0.155672
R1432 VDD1.n54 VDD1.n25 0.155672
R1433 VDD1.n47 VDD1.n25 0.155672
R1434 VDD1.n47 VDD1.n46 0.155672
R1435 VDD1.n46 VDD1.n30 0.155672
R1436 VDD1.n39 VDD1.n30 0.155672
R1437 VDD1.n39 VDD1.n38 0.155672
R1438 VDD1.n143 VDD1.n142 0.155672
R1439 VDD1.n143 VDD1.n134 0.155672
R1440 VDD1.n150 VDD1.n134 0.155672
R1441 VDD1.n151 VDD1.n150 0.155672
R1442 VDD1.n151 VDD1.n130 0.155672
R1443 VDD1.n159 VDD1.n130 0.155672
R1444 VDD1.n160 VDD1.n159 0.155672
R1445 VDD1.n160 VDD1.n126 0.155672
R1446 VDD1.n168 VDD1.n126 0.155672
R1447 VDD1.n169 VDD1.n168 0.155672
R1448 VDD1.n169 VDD1.n122 0.155672
R1449 VDD1.n176 VDD1.n122 0.155672
R1450 VDD1.n177 VDD1.n176 0.155672
R1451 VDD1.n177 VDD1.n118 0.155672
R1452 VDD1.n184 VDD1.n118 0.155672
R1453 VDD1.n185 VDD1.n184 0.155672
R1454 VDD1.n185 VDD1.n114 0.155672
R1455 VDD1.n192 VDD1.n114 0.155672
R1456 VDD1.n193 VDD1.n192 0.155672
R1457 VDD1.n193 VDD1.n110 0.155672
R1458 VDD1.n200 VDD1.n110 0.155672
R1459 VDD1.n201 VDD1.n200 0.155672
R1460 VDD1.n201 VDD1.n106 0.155672
R1461 VDD1.n208 VDD1.n106 0.155672
R1462 B.n190 B.t5 585.894
R1463 B.n68 B.t7 585.894
R1464 B.n196 B.t11 585.894
R1465 B.n62 B.t1 585.894
R1466 B.n711 B.n710 585
R1467 B.n712 B.n101 585
R1468 B.n714 B.n713 585
R1469 B.n715 B.n100 585
R1470 B.n717 B.n716 585
R1471 B.n718 B.n99 585
R1472 B.n720 B.n719 585
R1473 B.n721 B.n98 585
R1474 B.n723 B.n722 585
R1475 B.n724 B.n97 585
R1476 B.n726 B.n725 585
R1477 B.n727 B.n96 585
R1478 B.n729 B.n728 585
R1479 B.n730 B.n95 585
R1480 B.n732 B.n731 585
R1481 B.n733 B.n94 585
R1482 B.n735 B.n734 585
R1483 B.n736 B.n93 585
R1484 B.n738 B.n737 585
R1485 B.n739 B.n92 585
R1486 B.n741 B.n740 585
R1487 B.n742 B.n91 585
R1488 B.n744 B.n743 585
R1489 B.n745 B.n90 585
R1490 B.n747 B.n746 585
R1491 B.n748 B.n89 585
R1492 B.n750 B.n749 585
R1493 B.n751 B.n88 585
R1494 B.n753 B.n752 585
R1495 B.n754 B.n87 585
R1496 B.n756 B.n755 585
R1497 B.n757 B.n86 585
R1498 B.n759 B.n758 585
R1499 B.n760 B.n85 585
R1500 B.n762 B.n761 585
R1501 B.n763 B.n84 585
R1502 B.n765 B.n764 585
R1503 B.n766 B.n83 585
R1504 B.n768 B.n767 585
R1505 B.n769 B.n82 585
R1506 B.n771 B.n770 585
R1507 B.n772 B.n81 585
R1508 B.n774 B.n773 585
R1509 B.n775 B.n80 585
R1510 B.n777 B.n776 585
R1511 B.n778 B.n79 585
R1512 B.n780 B.n779 585
R1513 B.n781 B.n78 585
R1514 B.n783 B.n782 585
R1515 B.n784 B.n77 585
R1516 B.n786 B.n785 585
R1517 B.n787 B.n76 585
R1518 B.n789 B.n788 585
R1519 B.n790 B.n75 585
R1520 B.n792 B.n791 585
R1521 B.n793 B.n74 585
R1522 B.n795 B.n794 585
R1523 B.n796 B.n73 585
R1524 B.n798 B.n797 585
R1525 B.n799 B.n72 585
R1526 B.n801 B.n800 585
R1527 B.n802 B.n71 585
R1528 B.n804 B.n803 585
R1529 B.n806 B.n805 585
R1530 B.n807 B.n67 585
R1531 B.n809 B.n808 585
R1532 B.n810 B.n66 585
R1533 B.n812 B.n811 585
R1534 B.n813 B.n65 585
R1535 B.n815 B.n814 585
R1536 B.n816 B.n64 585
R1537 B.n818 B.n817 585
R1538 B.n819 B.n61 585
R1539 B.n822 B.n821 585
R1540 B.n823 B.n60 585
R1541 B.n825 B.n824 585
R1542 B.n826 B.n59 585
R1543 B.n828 B.n827 585
R1544 B.n829 B.n58 585
R1545 B.n831 B.n830 585
R1546 B.n832 B.n57 585
R1547 B.n834 B.n833 585
R1548 B.n835 B.n56 585
R1549 B.n837 B.n836 585
R1550 B.n838 B.n55 585
R1551 B.n840 B.n839 585
R1552 B.n841 B.n54 585
R1553 B.n843 B.n842 585
R1554 B.n844 B.n53 585
R1555 B.n846 B.n845 585
R1556 B.n847 B.n52 585
R1557 B.n849 B.n848 585
R1558 B.n850 B.n51 585
R1559 B.n852 B.n851 585
R1560 B.n853 B.n50 585
R1561 B.n855 B.n854 585
R1562 B.n856 B.n49 585
R1563 B.n858 B.n857 585
R1564 B.n859 B.n48 585
R1565 B.n861 B.n860 585
R1566 B.n862 B.n47 585
R1567 B.n864 B.n863 585
R1568 B.n865 B.n46 585
R1569 B.n867 B.n866 585
R1570 B.n868 B.n45 585
R1571 B.n870 B.n869 585
R1572 B.n871 B.n44 585
R1573 B.n873 B.n872 585
R1574 B.n874 B.n43 585
R1575 B.n876 B.n875 585
R1576 B.n877 B.n42 585
R1577 B.n879 B.n878 585
R1578 B.n880 B.n41 585
R1579 B.n882 B.n881 585
R1580 B.n883 B.n40 585
R1581 B.n885 B.n884 585
R1582 B.n886 B.n39 585
R1583 B.n888 B.n887 585
R1584 B.n889 B.n38 585
R1585 B.n891 B.n890 585
R1586 B.n892 B.n37 585
R1587 B.n894 B.n893 585
R1588 B.n895 B.n36 585
R1589 B.n897 B.n896 585
R1590 B.n898 B.n35 585
R1591 B.n900 B.n899 585
R1592 B.n901 B.n34 585
R1593 B.n903 B.n902 585
R1594 B.n904 B.n33 585
R1595 B.n906 B.n905 585
R1596 B.n907 B.n32 585
R1597 B.n909 B.n908 585
R1598 B.n910 B.n31 585
R1599 B.n912 B.n911 585
R1600 B.n913 B.n30 585
R1601 B.n915 B.n914 585
R1602 B.n709 B.n102 585
R1603 B.n708 B.n707 585
R1604 B.n706 B.n103 585
R1605 B.n705 B.n704 585
R1606 B.n703 B.n104 585
R1607 B.n702 B.n701 585
R1608 B.n700 B.n105 585
R1609 B.n699 B.n698 585
R1610 B.n697 B.n106 585
R1611 B.n696 B.n695 585
R1612 B.n694 B.n107 585
R1613 B.n693 B.n692 585
R1614 B.n691 B.n108 585
R1615 B.n690 B.n689 585
R1616 B.n688 B.n109 585
R1617 B.n687 B.n686 585
R1618 B.n685 B.n110 585
R1619 B.n684 B.n683 585
R1620 B.n682 B.n111 585
R1621 B.n681 B.n680 585
R1622 B.n679 B.n112 585
R1623 B.n678 B.n677 585
R1624 B.n676 B.n113 585
R1625 B.n675 B.n674 585
R1626 B.n673 B.n114 585
R1627 B.n672 B.n671 585
R1628 B.n670 B.n115 585
R1629 B.n669 B.n668 585
R1630 B.n667 B.n116 585
R1631 B.n666 B.n665 585
R1632 B.n664 B.n117 585
R1633 B.n663 B.n662 585
R1634 B.n661 B.n118 585
R1635 B.n660 B.n659 585
R1636 B.n658 B.n119 585
R1637 B.n657 B.n656 585
R1638 B.n655 B.n120 585
R1639 B.n654 B.n653 585
R1640 B.n652 B.n121 585
R1641 B.n651 B.n650 585
R1642 B.n649 B.n122 585
R1643 B.n648 B.n647 585
R1644 B.n646 B.n123 585
R1645 B.n645 B.n644 585
R1646 B.n643 B.n124 585
R1647 B.n642 B.n641 585
R1648 B.n640 B.n125 585
R1649 B.n639 B.n638 585
R1650 B.n637 B.n126 585
R1651 B.n636 B.n635 585
R1652 B.n634 B.n127 585
R1653 B.n633 B.n632 585
R1654 B.n631 B.n128 585
R1655 B.n630 B.n629 585
R1656 B.n628 B.n129 585
R1657 B.n627 B.n626 585
R1658 B.n625 B.n130 585
R1659 B.n624 B.n623 585
R1660 B.n622 B.n131 585
R1661 B.n621 B.n620 585
R1662 B.n619 B.n132 585
R1663 B.n618 B.n617 585
R1664 B.n616 B.n133 585
R1665 B.n615 B.n614 585
R1666 B.n613 B.n134 585
R1667 B.n612 B.n611 585
R1668 B.n610 B.n135 585
R1669 B.n609 B.n608 585
R1670 B.n607 B.n136 585
R1671 B.n606 B.n605 585
R1672 B.n604 B.n137 585
R1673 B.n603 B.n602 585
R1674 B.n601 B.n138 585
R1675 B.n600 B.n599 585
R1676 B.n598 B.n139 585
R1677 B.n597 B.n596 585
R1678 B.n595 B.n140 585
R1679 B.n594 B.n593 585
R1680 B.n592 B.n141 585
R1681 B.n591 B.n590 585
R1682 B.n589 B.n142 585
R1683 B.n588 B.n587 585
R1684 B.n586 B.n143 585
R1685 B.n585 B.n584 585
R1686 B.n583 B.n144 585
R1687 B.n582 B.n581 585
R1688 B.n580 B.n145 585
R1689 B.n579 B.n578 585
R1690 B.n577 B.n146 585
R1691 B.n576 B.n575 585
R1692 B.n574 B.n147 585
R1693 B.n573 B.n572 585
R1694 B.n571 B.n148 585
R1695 B.n570 B.n569 585
R1696 B.n568 B.n149 585
R1697 B.n567 B.n566 585
R1698 B.n565 B.n150 585
R1699 B.n564 B.n563 585
R1700 B.n562 B.n151 585
R1701 B.n561 B.n560 585
R1702 B.n559 B.n152 585
R1703 B.n558 B.n557 585
R1704 B.n556 B.n153 585
R1705 B.n555 B.n554 585
R1706 B.n553 B.n154 585
R1707 B.n552 B.n551 585
R1708 B.n550 B.n155 585
R1709 B.n549 B.n548 585
R1710 B.n547 B.n156 585
R1711 B.n546 B.n545 585
R1712 B.n544 B.n157 585
R1713 B.n339 B.n338 585
R1714 B.n340 B.n229 585
R1715 B.n342 B.n341 585
R1716 B.n343 B.n228 585
R1717 B.n345 B.n344 585
R1718 B.n346 B.n227 585
R1719 B.n348 B.n347 585
R1720 B.n349 B.n226 585
R1721 B.n351 B.n350 585
R1722 B.n352 B.n225 585
R1723 B.n354 B.n353 585
R1724 B.n355 B.n224 585
R1725 B.n357 B.n356 585
R1726 B.n358 B.n223 585
R1727 B.n360 B.n359 585
R1728 B.n361 B.n222 585
R1729 B.n363 B.n362 585
R1730 B.n364 B.n221 585
R1731 B.n366 B.n365 585
R1732 B.n367 B.n220 585
R1733 B.n369 B.n368 585
R1734 B.n370 B.n219 585
R1735 B.n372 B.n371 585
R1736 B.n373 B.n218 585
R1737 B.n375 B.n374 585
R1738 B.n376 B.n217 585
R1739 B.n378 B.n377 585
R1740 B.n379 B.n216 585
R1741 B.n381 B.n380 585
R1742 B.n382 B.n215 585
R1743 B.n384 B.n383 585
R1744 B.n385 B.n214 585
R1745 B.n387 B.n386 585
R1746 B.n388 B.n213 585
R1747 B.n390 B.n389 585
R1748 B.n391 B.n212 585
R1749 B.n393 B.n392 585
R1750 B.n394 B.n211 585
R1751 B.n396 B.n395 585
R1752 B.n397 B.n210 585
R1753 B.n399 B.n398 585
R1754 B.n400 B.n209 585
R1755 B.n402 B.n401 585
R1756 B.n403 B.n208 585
R1757 B.n405 B.n404 585
R1758 B.n406 B.n207 585
R1759 B.n408 B.n407 585
R1760 B.n409 B.n206 585
R1761 B.n411 B.n410 585
R1762 B.n412 B.n205 585
R1763 B.n414 B.n413 585
R1764 B.n415 B.n204 585
R1765 B.n417 B.n416 585
R1766 B.n418 B.n203 585
R1767 B.n420 B.n419 585
R1768 B.n421 B.n202 585
R1769 B.n423 B.n422 585
R1770 B.n424 B.n201 585
R1771 B.n426 B.n425 585
R1772 B.n427 B.n200 585
R1773 B.n429 B.n428 585
R1774 B.n430 B.n199 585
R1775 B.n432 B.n431 585
R1776 B.n434 B.n433 585
R1777 B.n435 B.n195 585
R1778 B.n437 B.n436 585
R1779 B.n438 B.n194 585
R1780 B.n440 B.n439 585
R1781 B.n441 B.n193 585
R1782 B.n443 B.n442 585
R1783 B.n444 B.n192 585
R1784 B.n446 B.n445 585
R1785 B.n447 B.n189 585
R1786 B.n450 B.n449 585
R1787 B.n451 B.n188 585
R1788 B.n453 B.n452 585
R1789 B.n454 B.n187 585
R1790 B.n456 B.n455 585
R1791 B.n457 B.n186 585
R1792 B.n459 B.n458 585
R1793 B.n460 B.n185 585
R1794 B.n462 B.n461 585
R1795 B.n463 B.n184 585
R1796 B.n465 B.n464 585
R1797 B.n466 B.n183 585
R1798 B.n468 B.n467 585
R1799 B.n469 B.n182 585
R1800 B.n471 B.n470 585
R1801 B.n472 B.n181 585
R1802 B.n474 B.n473 585
R1803 B.n475 B.n180 585
R1804 B.n477 B.n476 585
R1805 B.n478 B.n179 585
R1806 B.n480 B.n479 585
R1807 B.n481 B.n178 585
R1808 B.n483 B.n482 585
R1809 B.n484 B.n177 585
R1810 B.n486 B.n485 585
R1811 B.n487 B.n176 585
R1812 B.n489 B.n488 585
R1813 B.n490 B.n175 585
R1814 B.n492 B.n491 585
R1815 B.n493 B.n174 585
R1816 B.n495 B.n494 585
R1817 B.n496 B.n173 585
R1818 B.n498 B.n497 585
R1819 B.n499 B.n172 585
R1820 B.n501 B.n500 585
R1821 B.n502 B.n171 585
R1822 B.n504 B.n503 585
R1823 B.n505 B.n170 585
R1824 B.n507 B.n506 585
R1825 B.n508 B.n169 585
R1826 B.n510 B.n509 585
R1827 B.n511 B.n168 585
R1828 B.n513 B.n512 585
R1829 B.n514 B.n167 585
R1830 B.n516 B.n515 585
R1831 B.n517 B.n166 585
R1832 B.n519 B.n518 585
R1833 B.n520 B.n165 585
R1834 B.n522 B.n521 585
R1835 B.n523 B.n164 585
R1836 B.n525 B.n524 585
R1837 B.n526 B.n163 585
R1838 B.n528 B.n527 585
R1839 B.n529 B.n162 585
R1840 B.n531 B.n530 585
R1841 B.n532 B.n161 585
R1842 B.n534 B.n533 585
R1843 B.n535 B.n160 585
R1844 B.n537 B.n536 585
R1845 B.n538 B.n159 585
R1846 B.n540 B.n539 585
R1847 B.n541 B.n158 585
R1848 B.n543 B.n542 585
R1849 B.n337 B.n230 585
R1850 B.n336 B.n335 585
R1851 B.n334 B.n231 585
R1852 B.n333 B.n332 585
R1853 B.n331 B.n232 585
R1854 B.n330 B.n329 585
R1855 B.n328 B.n233 585
R1856 B.n327 B.n326 585
R1857 B.n325 B.n234 585
R1858 B.n324 B.n323 585
R1859 B.n322 B.n235 585
R1860 B.n321 B.n320 585
R1861 B.n319 B.n236 585
R1862 B.n318 B.n317 585
R1863 B.n316 B.n237 585
R1864 B.n315 B.n314 585
R1865 B.n313 B.n238 585
R1866 B.n312 B.n311 585
R1867 B.n310 B.n239 585
R1868 B.n309 B.n308 585
R1869 B.n307 B.n240 585
R1870 B.n306 B.n305 585
R1871 B.n304 B.n241 585
R1872 B.n303 B.n302 585
R1873 B.n301 B.n242 585
R1874 B.n300 B.n299 585
R1875 B.n298 B.n243 585
R1876 B.n297 B.n296 585
R1877 B.n295 B.n244 585
R1878 B.n294 B.n293 585
R1879 B.n292 B.n245 585
R1880 B.n291 B.n290 585
R1881 B.n289 B.n246 585
R1882 B.n288 B.n287 585
R1883 B.n286 B.n247 585
R1884 B.n285 B.n284 585
R1885 B.n283 B.n248 585
R1886 B.n282 B.n281 585
R1887 B.n280 B.n249 585
R1888 B.n279 B.n278 585
R1889 B.n277 B.n250 585
R1890 B.n276 B.n275 585
R1891 B.n274 B.n251 585
R1892 B.n273 B.n272 585
R1893 B.n271 B.n252 585
R1894 B.n270 B.n269 585
R1895 B.n268 B.n253 585
R1896 B.n267 B.n266 585
R1897 B.n265 B.n254 585
R1898 B.n264 B.n263 585
R1899 B.n262 B.n255 585
R1900 B.n261 B.n260 585
R1901 B.n259 B.n256 585
R1902 B.n258 B.n257 585
R1903 B.n2 B.n0 585
R1904 B.n997 B.n1 585
R1905 B.n996 B.n995 585
R1906 B.n994 B.n3 585
R1907 B.n993 B.n992 585
R1908 B.n991 B.n4 585
R1909 B.n990 B.n989 585
R1910 B.n988 B.n5 585
R1911 B.n987 B.n986 585
R1912 B.n985 B.n6 585
R1913 B.n984 B.n983 585
R1914 B.n982 B.n7 585
R1915 B.n981 B.n980 585
R1916 B.n979 B.n8 585
R1917 B.n978 B.n977 585
R1918 B.n976 B.n9 585
R1919 B.n975 B.n974 585
R1920 B.n973 B.n10 585
R1921 B.n972 B.n971 585
R1922 B.n970 B.n11 585
R1923 B.n969 B.n968 585
R1924 B.n967 B.n12 585
R1925 B.n966 B.n965 585
R1926 B.n964 B.n13 585
R1927 B.n963 B.n962 585
R1928 B.n961 B.n14 585
R1929 B.n960 B.n959 585
R1930 B.n958 B.n15 585
R1931 B.n957 B.n956 585
R1932 B.n955 B.n16 585
R1933 B.n954 B.n953 585
R1934 B.n952 B.n17 585
R1935 B.n951 B.n950 585
R1936 B.n949 B.n18 585
R1937 B.n948 B.n947 585
R1938 B.n946 B.n19 585
R1939 B.n945 B.n944 585
R1940 B.n943 B.n20 585
R1941 B.n942 B.n941 585
R1942 B.n940 B.n21 585
R1943 B.n939 B.n938 585
R1944 B.n937 B.n22 585
R1945 B.n936 B.n935 585
R1946 B.n934 B.n23 585
R1947 B.n933 B.n932 585
R1948 B.n931 B.n24 585
R1949 B.n930 B.n929 585
R1950 B.n928 B.n25 585
R1951 B.n927 B.n926 585
R1952 B.n925 B.n26 585
R1953 B.n924 B.n923 585
R1954 B.n922 B.n27 585
R1955 B.n921 B.n920 585
R1956 B.n919 B.n28 585
R1957 B.n918 B.n917 585
R1958 B.n916 B.n29 585
R1959 B.n999 B.n998 585
R1960 B.n191 B.t4 508.901
R1961 B.n69 B.t8 508.901
R1962 B.n197 B.t10 508.901
R1963 B.n63 B.t2 508.901
R1964 B.n338 B.n337 502.111
R1965 B.n914 B.n29 502.111
R1966 B.n542 B.n157 502.111
R1967 B.n710 B.n709 502.111
R1968 B.n190 B.t3 337.726
R1969 B.n196 B.t9 337.726
R1970 B.n62 B.t0 337.726
R1971 B.n68 B.t6 337.726
R1972 B.n337 B.n336 163.367
R1973 B.n336 B.n231 163.367
R1974 B.n332 B.n231 163.367
R1975 B.n332 B.n331 163.367
R1976 B.n331 B.n330 163.367
R1977 B.n330 B.n233 163.367
R1978 B.n326 B.n233 163.367
R1979 B.n326 B.n325 163.367
R1980 B.n325 B.n324 163.367
R1981 B.n324 B.n235 163.367
R1982 B.n320 B.n235 163.367
R1983 B.n320 B.n319 163.367
R1984 B.n319 B.n318 163.367
R1985 B.n318 B.n237 163.367
R1986 B.n314 B.n237 163.367
R1987 B.n314 B.n313 163.367
R1988 B.n313 B.n312 163.367
R1989 B.n312 B.n239 163.367
R1990 B.n308 B.n239 163.367
R1991 B.n308 B.n307 163.367
R1992 B.n307 B.n306 163.367
R1993 B.n306 B.n241 163.367
R1994 B.n302 B.n241 163.367
R1995 B.n302 B.n301 163.367
R1996 B.n301 B.n300 163.367
R1997 B.n300 B.n243 163.367
R1998 B.n296 B.n243 163.367
R1999 B.n296 B.n295 163.367
R2000 B.n295 B.n294 163.367
R2001 B.n294 B.n245 163.367
R2002 B.n290 B.n245 163.367
R2003 B.n290 B.n289 163.367
R2004 B.n289 B.n288 163.367
R2005 B.n288 B.n247 163.367
R2006 B.n284 B.n247 163.367
R2007 B.n284 B.n283 163.367
R2008 B.n283 B.n282 163.367
R2009 B.n282 B.n249 163.367
R2010 B.n278 B.n249 163.367
R2011 B.n278 B.n277 163.367
R2012 B.n277 B.n276 163.367
R2013 B.n276 B.n251 163.367
R2014 B.n272 B.n251 163.367
R2015 B.n272 B.n271 163.367
R2016 B.n271 B.n270 163.367
R2017 B.n270 B.n253 163.367
R2018 B.n266 B.n253 163.367
R2019 B.n266 B.n265 163.367
R2020 B.n265 B.n264 163.367
R2021 B.n264 B.n255 163.367
R2022 B.n260 B.n255 163.367
R2023 B.n260 B.n259 163.367
R2024 B.n259 B.n258 163.367
R2025 B.n258 B.n2 163.367
R2026 B.n998 B.n2 163.367
R2027 B.n998 B.n997 163.367
R2028 B.n997 B.n996 163.367
R2029 B.n996 B.n3 163.367
R2030 B.n992 B.n3 163.367
R2031 B.n992 B.n991 163.367
R2032 B.n991 B.n990 163.367
R2033 B.n990 B.n5 163.367
R2034 B.n986 B.n5 163.367
R2035 B.n986 B.n985 163.367
R2036 B.n985 B.n984 163.367
R2037 B.n984 B.n7 163.367
R2038 B.n980 B.n7 163.367
R2039 B.n980 B.n979 163.367
R2040 B.n979 B.n978 163.367
R2041 B.n978 B.n9 163.367
R2042 B.n974 B.n9 163.367
R2043 B.n974 B.n973 163.367
R2044 B.n973 B.n972 163.367
R2045 B.n972 B.n11 163.367
R2046 B.n968 B.n11 163.367
R2047 B.n968 B.n967 163.367
R2048 B.n967 B.n966 163.367
R2049 B.n966 B.n13 163.367
R2050 B.n962 B.n13 163.367
R2051 B.n962 B.n961 163.367
R2052 B.n961 B.n960 163.367
R2053 B.n960 B.n15 163.367
R2054 B.n956 B.n15 163.367
R2055 B.n956 B.n955 163.367
R2056 B.n955 B.n954 163.367
R2057 B.n954 B.n17 163.367
R2058 B.n950 B.n17 163.367
R2059 B.n950 B.n949 163.367
R2060 B.n949 B.n948 163.367
R2061 B.n948 B.n19 163.367
R2062 B.n944 B.n19 163.367
R2063 B.n944 B.n943 163.367
R2064 B.n943 B.n942 163.367
R2065 B.n942 B.n21 163.367
R2066 B.n938 B.n21 163.367
R2067 B.n938 B.n937 163.367
R2068 B.n937 B.n936 163.367
R2069 B.n936 B.n23 163.367
R2070 B.n932 B.n23 163.367
R2071 B.n932 B.n931 163.367
R2072 B.n931 B.n930 163.367
R2073 B.n930 B.n25 163.367
R2074 B.n926 B.n25 163.367
R2075 B.n926 B.n925 163.367
R2076 B.n925 B.n924 163.367
R2077 B.n924 B.n27 163.367
R2078 B.n920 B.n27 163.367
R2079 B.n920 B.n919 163.367
R2080 B.n919 B.n918 163.367
R2081 B.n918 B.n29 163.367
R2082 B.n338 B.n229 163.367
R2083 B.n342 B.n229 163.367
R2084 B.n343 B.n342 163.367
R2085 B.n344 B.n343 163.367
R2086 B.n344 B.n227 163.367
R2087 B.n348 B.n227 163.367
R2088 B.n349 B.n348 163.367
R2089 B.n350 B.n349 163.367
R2090 B.n350 B.n225 163.367
R2091 B.n354 B.n225 163.367
R2092 B.n355 B.n354 163.367
R2093 B.n356 B.n355 163.367
R2094 B.n356 B.n223 163.367
R2095 B.n360 B.n223 163.367
R2096 B.n361 B.n360 163.367
R2097 B.n362 B.n361 163.367
R2098 B.n362 B.n221 163.367
R2099 B.n366 B.n221 163.367
R2100 B.n367 B.n366 163.367
R2101 B.n368 B.n367 163.367
R2102 B.n368 B.n219 163.367
R2103 B.n372 B.n219 163.367
R2104 B.n373 B.n372 163.367
R2105 B.n374 B.n373 163.367
R2106 B.n374 B.n217 163.367
R2107 B.n378 B.n217 163.367
R2108 B.n379 B.n378 163.367
R2109 B.n380 B.n379 163.367
R2110 B.n380 B.n215 163.367
R2111 B.n384 B.n215 163.367
R2112 B.n385 B.n384 163.367
R2113 B.n386 B.n385 163.367
R2114 B.n386 B.n213 163.367
R2115 B.n390 B.n213 163.367
R2116 B.n391 B.n390 163.367
R2117 B.n392 B.n391 163.367
R2118 B.n392 B.n211 163.367
R2119 B.n396 B.n211 163.367
R2120 B.n397 B.n396 163.367
R2121 B.n398 B.n397 163.367
R2122 B.n398 B.n209 163.367
R2123 B.n402 B.n209 163.367
R2124 B.n403 B.n402 163.367
R2125 B.n404 B.n403 163.367
R2126 B.n404 B.n207 163.367
R2127 B.n408 B.n207 163.367
R2128 B.n409 B.n408 163.367
R2129 B.n410 B.n409 163.367
R2130 B.n410 B.n205 163.367
R2131 B.n414 B.n205 163.367
R2132 B.n415 B.n414 163.367
R2133 B.n416 B.n415 163.367
R2134 B.n416 B.n203 163.367
R2135 B.n420 B.n203 163.367
R2136 B.n421 B.n420 163.367
R2137 B.n422 B.n421 163.367
R2138 B.n422 B.n201 163.367
R2139 B.n426 B.n201 163.367
R2140 B.n427 B.n426 163.367
R2141 B.n428 B.n427 163.367
R2142 B.n428 B.n199 163.367
R2143 B.n432 B.n199 163.367
R2144 B.n433 B.n432 163.367
R2145 B.n433 B.n195 163.367
R2146 B.n437 B.n195 163.367
R2147 B.n438 B.n437 163.367
R2148 B.n439 B.n438 163.367
R2149 B.n439 B.n193 163.367
R2150 B.n443 B.n193 163.367
R2151 B.n444 B.n443 163.367
R2152 B.n445 B.n444 163.367
R2153 B.n445 B.n189 163.367
R2154 B.n450 B.n189 163.367
R2155 B.n451 B.n450 163.367
R2156 B.n452 B.n451 163.367
R2157 B.n452 B.n187 163.367
R2158 B.n456 B.n187 163.367
R2159 B.n457 B.n456 163.367
R2160 B.n458 B.n457 163.367
R2161 B.n458 B.n185 163.367
R2162 B.n462 B.n185 163.367
R2163 B.n463 B.n462 163.367
R2164 B.n464 B.n463 163.367
R2165 B.n464 B.n183 163.367
R2166 B.n468 B.n183 163.367
R2167 B.n469 B.n468 163.367
R2168 B.n470 B.n469 163.367
R2169 B.n470 B.n181 163.367
R2170 B.n474 B.n181 163.367
R2171 B.n475 B.n474 163.367
R2172 B.n476 B.n475 163.367
R2173 B.n476 B.n179 163.367
R2174 B.n480 B.n179 163.367
R2175 B.n481 B.n480 163.367
R2176 B.n482 B.n481 163.367
R2177 B.n482 B.n177 163.367
R2178 B.n486 B.n177 163.367
R2179 B.n487 B.n486 163.367
R2180 B.n488 B.n487 163.367
R2181 B.n488 B.n175 163.367
R2182 B.n492 B.n175 163.367
R2183 B.n493 B.n492 163.367
R2184 B.n494 B.n493 163.367
R2185 B.n494 B.n173 163.367
R2186 B.n498 B.n173 163.367
R2187 B.n499 B.n498 163.367
R2188 B.n500 B.n499 163.367
R2189 B.n500 B.n171 163.367
R2190 B.n504 B.n171 163.367
R2191 B.n505 B.n504 163.367
R2192 B.n506 B.n505 163.367
R2193 B.n506 B.n169 163.367
R2194 B.n510 B.n169 163.367
R2195 B.n511 B.n510 163.367
R2196 B.n512 B.n511 163.367
R2197 B.n512 B.n167 163.367
R2198 B.n516 B.n167 163.367
R2199 B.n517 B.n516 163.367
R2200 B.n518 B.n517 163.367
R2201 B.n518 B.n165 163.367
R2202 B.n522 B.n165 163.367
R2203 B.n523 B.n522 163.367
R2204 B.n524 B.n523 163.367
R2205 B.n524 B.n163 163.367
R2206 B.n528 B.n163 163.367
R2207 B.n529 B.n528 163.367
R2208 B.n530 B.n529 163.367
R2209 B.n530 B.n161 163.367
R2210 B.n534 B.n161 163.367
R2211 B.n535 B.n534 163.367
R2212 B.n536 B.n535 163.367
R2213 B.n536 B.n159 163.367
R2214 B.n540 B.n159 163.367
R2215 B.n541 B.n540 163.367
R2216 B.n542 B.n541 163.367
R2217 B.n546 B.n157 163.367
R2218 B.n547 B.n546 163.367
R2219 B.n548 B.n547 163.367
R2220 B.n548 B.n155 163.367
R2221 B.n552 B.n155 163.367
R2222 B.n553 B.n552 163.367
R2223 B.n554 B.n553 163.367
R2224 B.n554 B.n153 163.367
R2225 B.n558 B.n153 163.367
R2226 B.n559 B.n558 163.367
R2227 B.n560 B.n559 163.367
R2228 B.n560 B.n151 163.367
R2229 B.n564 B.n151 163.367
R2230 B.n565 B.n564 163.367
R2231 B.n566 B.n565 163.367
R2232 B.n566 B.n149 163.367
R2233 B.n570 B.n149 163.367
R2234 B.n571 B.n570 163.367
R2235 B.n572 B.n571 163.367
R2236 B.n572 B.n147 163.367
R2237 B.n576 B.n147 163.367
R2238 B.n577 B.n576 163.367
R2239 B.n578 B.n577 163.367
R2240 B.n578 B.n145 163.367
R2241 B.n582 B.n145 163.367
R2242 B.n583 B.n582 163.367
R2243 B.n584 B.n583 163.367
R2244 B.n584 B.n143 163.367
R2245 B.n588 B.n143 163.367
R2246 B.n589 B.n588 163.367
R2247 B.n590 B.n589 163.367
R2248 B.n590 B.n141 163.367
R2249 B.n594 B.n141 163.367
R2250 B.n595 B.n594 163.367
R2251 B.n596 B.n595 163.367
R2252 B.n596 B.n139 163.367
R2253 B.n600 B.n139 163.367
R2254 B.n601 B.n600 163.367
R2255 B.n602 B.n601 163.367
R2256 B.n602 B.n137 163.367
R2257 B.n606 B.n137 163.367
R2258 B.n607 B.n606 163.367
R2259 B.n608 B.n607 163.367
R2260 B.n608 B.n135 163.367
R2261 B.n612 B.n135 163.367
R2262 B.n613 B.n612 163.367
R2263 B.n614 B.n613 163.367
R2264 B.n614 B.n133 163.367
R2265 B.n618 B.n133 163.367
R2266 B.n619 B.n618 163.367
R2267 B.n620 B.n619 163.367
R2268 B.n620 B.n131 163.367
R2269 B.n624 B.n131 163.367
R2270 B.n625 B.n624 163.367
R2271 B.n626 B.n625 163.367
R2272 B.n626 B.n129 163.367
R2273 B.n630 B.n129 163.367
R2274 B.n631 B.n630 163.367
R2275 B.n632 B.n631 163.367
R2276 B.n632 B.n127 163.367
R2277 B.n636 B.n127 163.367
R2278 B.n637 B.n636 163.367
R2279 B.n638 B.n637 163.367
R2280 B.n638 B.n125 163.367
R2281 B.n642 B.n125 163.367
R2282 B.n643 B.n642 163.367
R2283 B.n644 B.n643 163.367
R2284 B.n644 B.n123 163.367
R2285 B.n648 B.n123 163.367
R2286 B.n649 B.n648 163.367
R2287 B.n650 B.n649 163.367
R2288 B.n650 B.n121 163.367
R2289 B.n654 B.n121 163.367
R2290 B.n655 B.n654 163.367
R2291 B.n656 B.n655 163.367
R2292 B.n656 B.n119 163.367
R2293 B.n660 B.n119 163.367
R2294 B.n661 B.n660 163.367
R2295 B.n662 B.n661 163.367
R2296 B.n662 B.n117 163.367
R2297 B.n666 B.n117 163.367
R2298 B.n667 B.n666 163.367
R2299 B.n668 B.n667 163.367
R2300 B.n668 B.n115 163.367
R2301 B.n672 B.n115 163.367
R2302 B.n673 B.n672 163.367
R2303 B.n674 B.n673 163.367
R2304 B.n674 B.n113 163.367
R2305 B.n678 B.n113 163.367
R2306 B.n679 B.n678 163.367
R2307 B.n680 B.n679 163.367
R2308 B.n680 B.n111 163.367
R2309 B.n684 B.n111 163.367
R2310 B.n685 B.n684 163.367
R2311 B.n686 B.n685 163.367
R2312 B.n686 B.n109 163.367
R2313 B.n690 B.n109 163.367
R2314 B.n691 B.n690 163.367
R2315 B.n692 B.n691 163.367
R2316 B.n692 B.n107 163.367
R2317 B.n696 B.n107 163.367
R2318 B.n697 B.n696 163.367
R2319 B.n698 B.n697 163.367
R2320 B.n698 B.n105 163.367
R2321 B.n702 B.n105 163.367
R2322 B.n703 B.n702 163.367
R2323 B.n704 B.n703 163.367
R2324 B.n704 B.n103 163.367
R2325 B.n708 B.n103 163.367
R2326 B.n709 B.n708 163.367
R2327 B.n914 B.n913 163.367
R2328 B.n913 B.n912 163.367
R2329 B.n912 B.n31 163.367
R2330 B.n908 B.n31 163.367
R2331 B.n908 B.n907 163.367
R2332 B.n907 B.n906 163.367
R2333 B.n906 B.n33 163.367
R2334 B.n902 B.n33 163.367
R2335 B.n902 B.n901 163.367
R2336 B.n901 B.n900 163.367
R2337 B.n900 B.n35 163.367
R2338 B.n896 B.n35 163.367
R2339 B.n896 B.n895 163.367
R2340 B.n895 B.n894 163.367
R2341 B.n894 B.n37 163.367
R2342 B.n890 B.n37 163.367
R2343 B.n890 B.n889 163.367
R2344 B.n889 B.n888 163.367
R2345 B.n888 B.n39 163.367
R2346 B.n884 B.n39 163.367
R2347 B.n884 B.n883 163.367
R2348 B.n883 B.n882 163.367
R2349 B.n882 B.n41 163.367
R2350 B.n878 B.n41 163.367
R2351 B.n878 B.n877 163.367
R2352 B.n877 B.n876 163.367
R2353 B.n876 B.n43 163.367
R2354 B.n872 B.n43 163.367
R2355 B.n872 B.n871 163.367
R2356 B.n871 B.n870 163.367
R2357 B.n870 B.n45 163.367
R2358 B.n866 B.n45 163.367
R2359 B.n866 B.n865 163.367
R2360 B.n865 B.n864 163.367
R2361 B.n864 B.n47 163.367
R2362 B.n860 B.n47 163.367
R2363 B.n860 B.n859 163.367
R2364 B.n859 B.n858 163.367
R2365 B.n858 B.n49 163.367
R2366 B.n854 B.n49 163.367
R2367 B.n854 B.n853 163.367
R2368 B.n853 B.n852 163.367
R2369 B.n852 B.n51 163.367
R2370 B.n848 B.n51 163.367
R2371 B.n848 B.n847 163.367
R2372 B.n847 B.n846 163.367
R2373 B.n846 B.n53 163.367
R2374 B.n842 B.n53 163.367
R2375 B.n842 B.n841 163.367
R2376 B.n841 B.n840 163.367
R2377 B.n840 B.n55 163.367
R2378 B.n836 B.n55 163.367
R2379 B.n836 B.n835 163.367
R2380 B.n835 B.n834 163.367
R2381 B.n834 B.n57 163.367
R2382 B.n830 B.n57 163.367
R2383 B.n830 B.n829 163.367
R2384 B.n829 B.n828 163.367
R2385 B.n828 B.n59 163.367
R2386 B.n824 B.n59 163.367
R2387 B.n824 B.n823 163.367
R2388 B.n823 B.n822 163.367
R2389 B.n822 B.n61 163.367
R2390 B.n817 B.n61 163.367
R2391 B.n817 B.n816 163.367
R2392 B.n816 B.n815 163.367
R2393 B.n815 B.n65 163.367
R2394 B.n811 B.n65 163.367
R2395 B.n811 B.n810 163.367
R2396 B.n810 B.n809 163.367
R2397 B.n809 B.n67 163.367
R2398 B.n805 B.n67 163.367
R2399 B.n805 B.n804 163.367
R2400 B.n804 B.n71 163.367
R2401 B.n800 B.n71 163.367
R2402 B.n800 B.n799 163.367
R2403 B.n799 B.n798 163.367
R2404 B.n798 B.n73 163.367
R2405 B.n794 B.n73 163.367
R2406 B.n794 B.n793 163.367
R2407 B.n793 B.n792 163.367
R2408 B.n792 B.n75 163.367
R2409 B.n788 B.n75 163.367
R2410 B.n788 B.n787 163.367
R2411 B.n787 B.n786 163.367
R2412 B.n786 B.n77 163.367
R2413 B.n782 B.n77 163.367
R2414 B.n782 B.n781 163.367
R2415 B.n781 B.n780 163.367
R2416 B.n780 B.n79 163.367
R2417 B.n776 B.n79 163.367
R2418 B.n776 B.n775 163.367
R2419 B.n775 B.n774 163.367
R2420 B.n774 B.n81 163.367
R2421 B.n770 B.n81 163.367
R2422 B.n770 B.n769 163.367
R2423 B.n769 B.n768 163.367
R2424 B.n768 B.n83 163.367
R2425 B.n764 B.n83 163.367
R2426 B.n764 B.n763 163.367
R2427 B.n763 B.n762 163.367
R2428 B.n762 B.n85 163.367
R2429 B.n758 B.n85 163.367
R2430 B.n758 B.n757 163.367
R2431 B.n757 B.n756 163.367
R2432 B.n756 B.n87 163.367
R2433 B.n752 B.n87 163.367
R2434 B.n752 B.n751 163.367
R2435 B.n751 B.n750 163.367
R2436 B.n750 B.n89 163.367
R2437 B.n746 B.n89 163.367
R2438 B.n746 B.n745 163.367
R2439 B.n745 B.n744 163.367
R2440 B.n744 B.n91 163.367
R2441 B.n740 B.n91 163.367
R2442 B.n740 B.n739 163.367
R2443 B.n739 B.n738 163.367
R2444 B.n738 B.n93 163.367
R2445 B.n734 B.n93 163.367
R2446 B.n734 B.n733 163.367
R2447 B.n733 B.n732 163.367
R2448 B.n732 B.n95 163.367
R2449 B.n728 B.n95 163.367
R2450 B.n728 B.n727 163.367
R2451 B.n727 B.n726 163.367
R2452 B.n726 B.n97 163.367
R2453 B.n722 B.n97 163.367
R2454 B.n722 B.n721 163.367
R2455 B.n721 B.n720 163.367
R2456 B.n720 B.n99 163.367
R2457 B.n716 B.n99 163.367
R2458 B.n716 B.n715 163.367
R2459 B.n715 B.n714 163.367
R2460 B.n714 B.n101 163.367
R2461 B.n710 B.n101 163.367
R2462 B.n191 B.n190 76.9944
R2463 B.n197 B.n196 76.9944
R2464 B.n63 B.n62 76.9944
R2465 B.n69 B.n68 76.9944
R2466 B.n448 B.n191 59.5399
R2467 B.n198 B.n197 59.5399
R2468 B.n820 B.n63 59.5399
R2469 B.n70 B.n69 59.5399
R2470 B.n916 B.n915 32.6249
R2471 B.n711 B.n102 32.6249
R2472 B.n544 B.n543 32.6249
R2473 B.n339 B.n230 32.6249
R2474 B B.n999 18.0485
R2475 B.n915 B.n30 10.6151
R2476 B.n911 B.n30 10.6151
R2477 B.n911 B.n910 10.6151
R2478 B.n910 B.n909 10.6151
R2479 B.n909 B.n32 10.6151
R2480 B.n905 B.n32 10.6151
R2481 B.n905 B.n904 10.6151
R2482 B.n904 B.n903 10.6151
R2483 B.n903 B.n34 10.6151
R2484 B.n899 B.n34 10.6151
R2485 B.n899 B.n898 10.6151
R2486 B.n898 B.n897 10.6151
R2487 B.n897 B.n36 10.6151
R2488 B.n893 B.n36 10.6151
R2489 B.n893 B.n892 10.6151
R2490 B.n892 B.n891 10.6151
R2491 B.n891 B.n38 10.6151
R2492 B.n887 B.n38 10.6151
R2493 B.n887 B.n886 10.6151
R2494 B.n886 B.n885 10.6151
R2495 B.n885 B.n40 10.6151
R2496 B.n881 B.n40 10.6151
R2497 B.n881 B.n880 10.6151
R2498 B.n880 B.n879 10.6151
R2499 B.n879 B.n42 10.6151
R2500 B.n875 B.n42 10.6151
R2501 B.n875 B.n874 10.6151
R2502 B.n874 B.n873 10.6151
R2503 B.n873 B.n44 10.6151
R2504 B.n869 B.n44 10.6151
R2505 B.n869 B.n868 10.6151
R2506 B.n868 B.n867 10.6151
R2507 B.n867 B.n46 10.6151
R2508 B.n863 B.n46 10.6151
R2509 B.n863 B.n862 10.6151
R2510 B.n862 B.n861 10.6151
R2511 B.n861 B.n48 10.6151
R2512 B.n857 B.n48 10.6151
R2513 B.n857 B.n856 10.6151
R2514 B.n856 B.n855 10.6151
R2515 B.n855 B.n50 10.6151
R2516 B.n851 B.n50 10.6151
R2517 B.n851 B.n850 10.6151
R2518 B.n850 B.n849 10.6151
R2519 B.n849 B.n52 10.6151
R2520 B.n845 B.n52 10.6151
R2521 B.n845 B.n844 10.6151
R2522 B.n844 B.n843 10.6151
R2523 B.n843 B.n54 10.6151
R2524 B.n839 B.n54 10.6151
R2525 B.n839 B.n838 10.6151
R2526 B.n838 B.n837 10.6151
R2527 B.n837 B.n56 10.6151
R2528 B.n833 B.n56 10.6151
R2529 B.n833 B.n832 10.6151
R2530 B.n832 B.n831 10.6151
R2531 B.n831 B.n58 10.6151
R2532 B.n827 B.n58 10.6151
R2533 B.n827 B.n826 10.6151
R2534 B.n826 B.n825 10.6151
R2535 B.n825 B.n60 10.6151
R2536 B.n821 B.n60 10.6151
R2537 B.n819 B.n818 10.6151
R2538 B.n818 B.n64 10.6151
R2539 B.n814 B.n64 10.6151
R2540 B.n814 B.n813 10.6151
R2541 B.n813 B.n812 10.6151
R2542 B.n812 B.n66 10.6151
R2543 B.n808 B.n66 10.6151
R2544 B.n808 B.n807 10.6151
R2545 B.n807 B.n806 10.6151
R2546 B.n803 B.n802 10.6151
R2547 B.n802 B.n801 10.6151
R2548 B.n801 B.n72 10.6151
R2549 B.n797 B.n72 10.6151
R2550 B.n797 B.n796 10.6151
R2551 B.n796 B.n795 10.6151
R2552 B.n795 B.n74 10.6151
R2553 B.n791 B.n74 10.6151
R2554 B.n791 B.n790 10.6151
R2555 B.n790 B.n789 10.6151
R2556 B.n789 B.n76 10.6151
R2557 B.n785 B.n76 10.6151
R2558 B.n785 B.n784 10.6151
R2559 B.n784 B.n783 10.6151
R2560 B.n783 B.n78 10.6151
R2561 B.n779 B.n78 10.6151
R2562 B.n779 B.n778 10.6151
R2563 B.n778 B.n777 10.6151
R2564 B.n777 B.n80 10.6151
R2565 B.n773 B.n80 10.6151
R2566 B.n773 B.n772 10.6151
R2567 B.n772 B.n771 10.6151
R2568 B.n771 B.n82 10.6151
R2569 B.n767 B.n82 10.6151
R2570 B.n767 B.n766 10.6151
R2571 B.n766 B.n765 10.6151
R2572 B.n765 B.n84 10.6151
R2573 B.n761 B.n84 10.6151
R2574 B.n761 B.n760 10.6151
R2575 B.n760 B.n759 10.6151
R2576 B.n759 B.n86 10.6151
R2577 B.n755 B.n86 10.6151
R2578 B.n755 B.n754 10.6151
R2579 B.n754 B.n753 10.6151
R2580 B.n753 B.n88 10.6151
R2581 B.n749 B.n88 10.6151
R2582 B.n749 B.n748 10.6151
R2583 B.n748 B.n747 10.6151
R2584 B.n747 B.n90 10.6151
R2585 B.n743 B.n90 10.6151
R2586 B.n743 B.n742 10.6151
R2587 B.n742 B.n741 10.6151
R2588 B.n741 B.n92 10.6151
R2589 B.n737 B.n92 10.6151
R2590 B.n737 B.n736 10.6151
R2591 B.n736 B.n735 10.6151
R2592 B.n735 B.n94 10.6151
R2593 B.n731 B.n94 10.6151
R2594 B.n731 B.n730 10.6151
R2595 B.n730 B.n729 10.6151
R2596 B.n729 B.n96 10.6151
R2597 B.n725 B.n96 10.6151
R2598 B.n725 B.n724 10.6151
R2599 B.n724 B.n723 10.6151
R2600 B.n723 B.n98 10.6151
R2601 B.n719 B.n98 10.6151
R2602 B.n719 B.n718 10.6151
R2603 B.n718 B.n717 10.6151
R2604 B.n717 B.n100 10.6151
R2605 B.n713 B.n100 10.6151
R2606 B.n713 B.n712 10.6151
R2607 B.n712 B.n711 10.6151
R2608 B.n545 B.n544 10.6151
R2609 B.n545 B.n156 10.6151
R2610 B.n549 B.n156 10.6151
R2611 B.n550 B.n549 10.6151
R2612 B.n551 B.n550 10.6151
R2613 B.n551 B.n154 10.6151
R2614 B.n555 B.n154 10.6151
R2615 B.n556 B.n555 10.6151
R2616 B.n557 B.n556 10.6151
R2617 B.n557 B.n152 10.6151
R2618 B.n561 B.n152 10.6151
R2619 B.n562 B.n561 10.6151
R2620 B.n563 B.n562 10.6151
R2621 B.n563 B.n150 10.6151
R2622 B.n567 B.n150 10.6151
R2623 B.n568 B.n567 10.6151
R2624 B.n569 B.n568 10.6151
R2625 B.n569 B.n148 10.6151
R2626 B.n573 B.n148 10.6151
R2627 B.n574 B.n573 10.6151
R2628 B.n575 B.n574 10.6151
R2629 B.n575 B.n146 10.6151
R2630 B.n579 B.n146 10.6151
R2631 B.n580 B.n579 10.6151
R2632 B.n581 B.n580 10.6151
R2633 B.n581 B.n144 10.6151
R2634 B.n585 B.n144 10.6151
R2635 B.n586 B.n585 10.6151
R2636 B.n587 B.n586 10.6151
R2637 B.n587 B.n142 10.6151
R2638 B.n591 B.n142 10.6151
R2639 B.n592 B.n591 10.6151
R2640 B.n593 B.n592 10.6151
R2641 B.n593 B.n140 10.6151
R2642 B.n597 B.n140 10.6151
R2643 B.n598 B.n597 10.6151
R2644 B.n599 B.n598 10.6151
R2645 B.n599 B.n138 10.6151
R2646 B.n603 B.n138 10.6151
R2647 B.n604 B.n603 10.6151
R2648 B.n605 B.n604 10.6151
R2649 B.n605 B.n136 10.6151
R2650 B.n609 B.n136 10.6151
R2651 B.n610 B.n609 10.6151
R2652 B.n611 B.n610 10.6151
R2653 B.n611 B.n134 10.6151
R2654 B.n615 B.n134 10.6151
R2655 B.n616 B.n615 10.6151
R2656 B.n617 B.n616 10.6151
R2657 B.n617 B.n132 10.6151
R2658 B.n621 B.n132 10.6151
R2659 B.n622 B.n621 10.6151
R2660 B.n623 B.n622 10.6151
R2661 B.n623 B.n130 10.6151
R2662 B.n627 B.n130 10.6151
R2663 B.n628 B.n627 10.6151
R2664 B.n629 B.n628 10.6151
R2665 B.n629 B.n128 10.6151
R2666 B.n633 B.n128 10.6151
R2667 B.n634 B.n633 10.6151
R2668 B.n635 B.n634 10.6151
R2669 B.n635 B.n126 10.6151
R2670 B.n639 B.n126 10.6151
R2671 B.n640 B.n639 10.6151
R2672 B.n641 B.n640 10.6151
R2673 B.n641 B.n124 10.6151
R2674 B.n645 B.n124 10.6151
R2675 B.n646 B.n645 10.6151
R2676 B.n647 B.n646 10.6151
R2677 B.n647 B.n122 10.6151
R2678 B.n651 B.n122 10.6151
R2679 B.n652 B.n651 10.6151
R2680 B.n653 B.n652 10.6151
R2681 B.n653 B.n120 10.6151
R2682 B.n657 B.n120 10.6151
R2683 B.n658 B.n657 10.6151
R2684 B.n659 B.n658 10.6151
R2685 B.n659 B.n118 10.6151
R2686 B.n663 B.n118 10.6151
R2687 B.n664 B.n663 10.6151
R2688 B.n665 B.n664 10.6151
R2689 B.n665 B.n116 10.6151
R2690 B.n669 B.n116 10.6151
R2691 B.n670 B.n669 10.6151
R2692 B.n671 B.n670 10.6151
R2693 B.n671 B.n114 10.6151
R2694 B.n675 B.n114 10.6151
R2695 B.n676 B.n675 10.6151
R2696 B.n677 B.n676 10.6151
R2697 B.n677 B.n112 10.6151
R2698 B.n681 B.n112 10.6151
R2699 B.n682 B.n681 10.6151
R2700 B.n683 B.n682 10.6151
R2701 B.n683 B.n110 10.6151
R2702 B.n687 B.n110 10.6151
R2703 B.n688 B.n687 10.6151
R2704 B.n689 B.n688 10.6151
R2705 B.n689 B.n108 10.6151
R2706 B.n693 B.n108 10.6151
R2707 B.n694 B.n693 10.6151
R2708 B.n695 B.n694 10.6151
R2709 B.n695 B.n106 10.6151
R2710 B.n699 B.n106 10.6151
R2711 B.n700 B.n699 10.6151
R2712 B.n701 B.n700 10.6151
R2713 B.n701 B.n104 10.6151
R2714 B.n705 B.n104 10.6151
R2715 B.n706 B.n705 10.6151
R2716 B.n707 B.n706 10.6151
R2717 B.n707 B.n102 10.6151
R2718 B.n340 B.n339 10.6151
R2719 B.n341 B.n340 10.6151
R2720 B.n341 B.n228 10.6151
R2721 B.n345 B.n228 10.6151
R2722 B.n346 B.n345 10.6151
R2723 B.n347 B.n346 10.6151
R2724 B.n347 B.n226 10.6151
R2725 B.n351 B.n226 10.6151
R2726 B.n352 B.n351 10.6151
R2727 B.n353 B.n352 10.6151
R2728 B.n353 B.n224 10.6151
R2729 B.n357 B.n224 10.6151
R2730 B.n358 B.n357 10.6151
R2731 B.n359 B.n358 10.6151
R2732 B.n359 B.n222 10.6151
R2733 B.n363 B.n222 10.6151
R2734 B.n364 B.n363 10.6151
R2735 B.n365 B.n364 10.6151
R2736 B.n365 B.n220 10.6151
R2737 B.n369 B.n220 10.6151
R2738 B.n370 B.n369 10.6151
R2739 B.n371 B.n370 10.6151
R2740 B.n371 B.n218 10.6151
R2741 B.n375 B.n218 10.6151
R2742 B.n376 B.n375 10.6151
R2743 B.n377 B.n376 10.6151
R2744 B.n377 B.n216 10.6151
R2745 B.n381 B.n216 10.6151
R2746 B.n382 B.n381 10.6151
R2747 B.n383 B.n382 10.6151
R2748 B.n383 B.n214 10.6151
R2749 B.n387 B.n214 10.6151
R2750 B.n388 B.n387 10.6151
R2751 B.n389 B.n388 10.6151
R2752 B.n389 B.n212 10.6151
R2753 B.n393 B.n212 10.6151
R2754 B.n394 B.n393 10.6151
R2755 B.n395 B.n394 10.6151
R2756 B.n395 B.n210 10.6151
R2757 B.n399 B.n210 10.6151
R2758 B.n400 B.n399 10.6151
R2759 B.n401 B.n400 10.6151
R2760 B.n401 B.n208 10.6151
R2761 B.n405 B.n208 10.6151
R2762 B.n406 B.n405 10.6151
R2763 B.n407 B.n406 10.6151
R2764 B.n407 B.n206 10.6151
R2765 B.n411 B.n206 10.6151
R2766 B.n412 B.n411 10.6151
R2767 B.n413 B.n412 10.6151
R2768 B.n413 B.n204 10.6151
R2769 B.n417 B.n204 10.6151
R2770 B.n418 B.n417 10.6151
R2771 B.n419 B.n418 10.6151
R2772 B.n419 B.n202 10.6151
R2773 B.n423 B.n202 10.6151
R2774 B.n424 B.n423 10.6151
R2775 B.n425 B.n424 10.6151
R2776 B.n425 B.n200 10.6151
R2777 B.n429 B.n200 10.6151
R2778 B.n430 B.n429 10.6151
R2779 B.n431 B.n430 10.6151
R2780 B.n435 B.n434 10.6151
R2781 B.n436 B.n435 10.6151
R2782 B.n436 B.n194 10.6151
R2783 B.n440 B.n194 10.6151
R2784 B.n441 B.n440 10.6151
R2785 B.n442 B.n441 10.6151
R2786 B.n442 B.n192 10.6151
R2787 B.n446 B.n192 10.6151
R2788 B.n447 B.n446 10.6151
R2789 B.n449 B.n188 10.6151
R2790 B.n453 B.n188 10.6151
R2791 B.n454 B.n453 10.6151
R2792 B.n455 B.n454 10.6151
R2793 B.n455 B.n186 10.6151
R2794 B.n459 B.n186 10.6151
R2795 B.n460 B.n459 10.6151
R2796 B.n461 B.n460 10.6151
R2797 B.n461 B.n184 10.6151
R2798 B.n465 B.n184 10.6151
R2799 B.n466 B.n465 10.6151
R2800 B.n467 B.n466 10.6151
R2801 B.n467 B.n182 10.6151
R2802 B.n471 B.n182 10.6151
R2803 B.n472 B.n471 10.6151
R2804 B.n473 B.n472 10.6151
R2805 B.n473 B.n180 10.6151
R2806 B.n477 B.n180 10.6151
R2807 B.n478 B.n477 10.6151
R2808 B.n479 B.n478 10.6151
R2809 B.n479 B.n178 10.6151
R2810 B.n483 B.n178 10.6151
R2811 B.n484 B.n483 10.6151
R2812 B.n485 B.n484 10.6151
R2813 B.n485 B.n176 10.6151
R2814 B.n489 B.n176 10.6151
R2815 B.n490 B.n489 10.6151
R2816 B.n491 B.n490 10.6151
R2817 B.n491 B.n174 10.6151
R2818 B.n495 B.n174 10.6151
R2819 B.n496 B.n495 10.6151
R2820 B.n497 B.n496 10.6151
R2821 B.n497 B.n172 10.6151
R2822 B.n501 B.n172 10.6151
R2823 B.n502 B.n501 10.6151
R2824 B.n503 B.n502 10.6151
R2825 B.n503 B.n170 10.6151
R2826 B.n507 B.n170 10.6151
R2827 B.n508 B.n507 10.6151
R2828 B.n509 B.n508 10.6151
R2829 B.n509 B.n168 10.6151
R2830 B.n513 B.n168 10.6151
R2831 B.n514 B.n513 10.6151
R2832 B.n515 B.n514 10.6151
R2833 B.n515 B.n166 10.6151
R2834 B.n519 B.n166 10.6151
R2835 B.n520 B.n519 10.6151
R2836 B.n521 B.n520 10.6151
R2837 B.n521 B.n164 10.6151
R2838 B.n525 B.n164 10.6151
R2839 B.n526 B.n525 10.6151
R2840 B.n527 B.n526 10.6151
R2841 B.n527 B.n162 10.6151
R2842 B.n531 B.n162 10.6151
R2843 B.n532 B.n531 10.6151
R2844 B.n533 B.n532 10.6151
R2845 B.n533 B.n160 10.6151
R2846 B.n537 B.n160 10.6151
R2847 B.n538 B.n537 10.6151
R2848 B.n539 B.n538 10.6151
R2849 B.n539 B.n158 10.6151
R2850 B.n543 B.n158 10.6151
R2851 B.n335 B.n230 10.6151
R2852 B.n335 B.n334 10.6151
R2853 B.n334 B.n333 10.6151
R2854 B.n333 B.n232 10.6151
R2855 B.n329 B.n232 10.6151
R2856 B.n329 B.n328 10.6151
R2857 B.n328 B.n327 10.6151
R2858 B.n327 B.n234 10.6151
R2859 B.n323 B.n234 10.6151
R2860 B.n323 B.n322 10.6151
R2861 B.n322 B.n321 10.6151
R2862 B.n321 B.n236 10.6151
R2863 B.n317 B.n236 10.6151
R2864 B.n317 B.n316 10.6151
R2865 B.n316 B.n315 10.6151
R2866 B.n315 B.n238 10.6151
R2867 B.n311 B.n238 10.6151
R2868 B.n311 B.n310 10.6151
R2869 B.n310 B.n309 10.6151
R2870 B.n309 B.n240 10.6151
R2871 B.n305 B.n240 10.6151
R2872 B.n305 B.n304 10.6151
R2873 B.n304 B.n303 10.6151
R2874 B.n303 B.n242 10.6151
R2875 B.n299 B.n242 10.6151
R2876 B.n299 B.n298 10.6151
R2877 B.n298 B.n297 10.6151
R2878 B.n297 B.n244 10.6151
R2879 B.n293 B.n244 10.6151
R2880 B.n293 B.n292 10.6151
R2881 B.n292 B.n291 10.6151
R2882 B.n291 B.n246 10.6151
R2883 B.n287 B.n246 10.6151
R2884 B.n287 B.n286 10.6151
R2885 B.n286 B.n285 10.6151
R2886 B.n285 B.n248 10.6151
R2887 B.n281 B.n248 10.6151
R2888 B.n281 B.n280 10.6151
R2889 B.n280 B.n279 10.6151
R2890 B.n279 B.n250 10.6151
R2891 B.n275 B.n250 10.6151
R2892 B.n275 B.n274 10.6151
R2893 B.n274 B.n273 10.6151
R2894 B.n273 B.n252 10.6151
R2895 B.n269 B.n252 10.6151
R2896 B.n269 B.n268 10.6151
R2897 B.n268 B.n267 10.6151
R2898 B.n267 B.n254 10.6151
R2899 B.n263 B.n254 10.6151
R2900 B.n263 B.n262 10.6151
R2901 B.n262 B.n261 10.6151
R2902 B.n261 B.n256 10.6151
R2903 B.n257 B.n256 10.6151
R2904 B.n257 B.n0 10.6151
R2905 B.n995 B.n1 10.6151
R2906 B.n995 B.n994 10.6151
R2907 B.n994 B.n993 10.6151
R2908 B.n993 B.n4 10.6151
R2909 B.n989 B.n4 10.6151
R2910 B.n989 B.n988 10.6151
R2911 B.n988 B.n987 10.6151
R2912 B.n987 B.n6 10.6151
R2913 B.n983 B.n6 10.6151
R2914 B.n983 B.n982 10.6151
R2915 B.n982 B.n981 10.6151
R2916 B.n981 B.n8 10.6151
R2917 B.n977 B.n8 10.6151
R2918 B.n977 B.n976 10.6151
R2919 B.n976 B.n975 10.6151
R2920 B.n975 B.n10 10.6151
R2921 B.n971 B.n10 10.6151
R2922 B.n971 B.n970 10.6151
R2923 B.n970 B.n969 10.6151
R2924 B.n969 B.n12 10.6151
R2925 B.n965 B.n12 10.6151
R2926 B.n965 B.n964 10.6151
R2927 B.n964 B.n963 10.6151
R2928 B.n963 B.n14 10.6151
R2929 B.n959 B.n14 10.6151
R2930 B.n959 B.n958 10.6151
R2931 B.n958 B.n957 10.6151
R2932 B.n957 B.n16 10.6151
R2933 B.n953 B.n16 10.6151
R2934 B.n953 B.n952 10.6151
R2935 B.n952 B.n951 10.6151
R2936 B.n951 B.n18 10.6151
R2937 B.n947 B.n18 10.6151
R2938 B.n947 B.n946 10.6151
R2939 B.n946 B.n945 10.6151
R2940 B.n945 B.n20 10.6151
R2941 B.n941 B.n20 10.6151
R2942 B.n941 B.n940 10.6151
R2943 B.n940 B.n939 10.6151
R2944 B.n939 B.n22 10.6151
R2945 B.n935 B.n22 10.6151
R2946 B.n935 B.n934 10.6151
R2947 B.n934 B.n933 10.6151
R2948 B.n933 B.n24 10.6151
R2949 B.n929 B.n24 10.6151
R2950 B.n929 B.n928 10.6151
R2951 B.n928 B.n927 10.6151
R2952 B.n927 B.n26 10.6151
R2953 B.n923 B.n26 10.6151
R2954 B.n923 B.n922 10.6151
R2955 B.n922 B.n921 10.6151
R2956 B.n921 B.n28 10.6151
R2957 B.n917 B.n28 10.6151
R2958 B.n917 B.n916 10.6151
R2959 B.n821 B.n820 9.36635
R2960 B.n803 B.n70 9.36635
R2961 B.n431 B.n198 9.36635
R2962 B.n449 B.n448 9.36635
R2963 B.n999 B.n0 2.81026
R2964 B.n999 B.n1 2.81026
R2965 B.n820 B.n819 1.24928
R2966 B.n806 B.n70 1.24928
R2967 B.n434 B.n198 1.24928
R2968 B.n448 B.n447 1.24928
C0 VDD1 w_n4146_n4850# 3.05028f
C1 VN w_n4146_n4850# 8.235379f
C2 VDD1 VN 0.152258f
C3 VDD2 w_n4146_n4850# 3.1686f
C4 VDD1 VDD2 1.81407f
C5 B w_n4146_n4850# 13.19f
C6 VDD1 B 2.96076f
C7 VTAIL w_n4146_n4850# 4.06986f
C8 VDD2 VN 11.2435f
C9 VDD1 VTAIL 10.4748f
C10 VN B 1.47367f
C11 VP w_n4146_n4850# 8.7743f
C12 VDD2 B 3.0598f
C13 VN VTAIL 11.3008f
C14 VDD1 VP 11.6343f
C15 VDD2 VTAIL 10.5322f
C16 VTAIL B 5.84063f
C17 VN VP 9.30781f
C18 VDD2 VP 0.546788f
C19 B VP 2.37869f
C20 VTAIL VP 11.3154f
C21 VDD2 VSUBS 2.35795f
C22 VDD1 VSUBS 2.383412f
C23 VTAIL VSUBS 1.654719f
C24 VN VSUBS 7.12449f
C25 VP VSUBS 4.014655f
C26 B VSUBS 6.290131f
C27 w_n4146_n4850# VSUBS 0.245626p
C28 B.n0 VSUBS 0.004457f
C29 B.n1 VSUBS 0.004457f
C30 B.n2 VSUBS 0.007047f
C31 B.n3 VSUBS 0.007047f
C32 B.n4 VSUBS 0.007047f
C33 B.n5 VSUBS 0.007047f
C34 B.n6 VSUBS 0.007047f
C35 B.n7 VSUBS 0.007047f
C36 B.n8 VSUBS 0.007047f
C37 B.n9 VSUBS 0.007047f
C38 B.n10 VSUBS 0.007047f
C39 B.n11 VSUBS 0.007047f
C40 B.n12 VSUBS 0.007047f
C41 B.n13 VSUBS 0.007047f
C42 B.n14 VSUBS 0.007047f
C43 B.n15 VSUBS 0.007047f
C44 B.n16 VSUBS 0.007047f
C45 B.n17 VSUBS 0.007047f
C46 B.n18 VSUBS 0.007047f
C47 B.n19 VSUBS 0.007047f
C48 B.n20 VSUBS 0.007047f
C49 B.n21 VSUBS 0.007047f
C50 B.n22 VSUBS 0.007047f
C51 B.n23 VSUBS 0.007047f
C52 B.n24 VSUBS 0.007047f
C53 B.n25 VSUBS 0.007047f
C54 B.n26 VSUBS 0.007047f
C55 B.n27 VSUBS 0.007047f
C56 B.n28 VSUBS 0.007047f
C57 B.n29 VSUBS 0.016346f
C58 B.n30 VSUBS 0.007047f
C59 B.n31 VSUBS 0.007047f
C60 B.n32 VSUBS 0.007047f
C61 B.n33 VSUBS 0.007047f
C62 B.n34 VSUBS 0.007047f
C63 B.n35 VSUBS 0.007047f
C64 B.n36 VSUBS 0.007047f
C65 B.n37 VSUBS 0.007047f
C66 B.n38 VSUBS 0.007047f
C67 B.n39 VSUBS 0.007047f
C68 B.n40 VSUBS 0.007047f
C69 B.n41 VSUBS 0.007047f
C70 B.n42 VSUBS 0.007047f
C71 B.n43 VSUBS 0.007047f
C72 B.n44 VSUBS 0.007047f
C73 B.n45 VSUBS 0.007047f
C74 B.n46 VSUBS 0.007047f
C75 B.n47 VSUBS 0.007047f
C76 B.n48 VSUBS 0.007047f
C77 B.n49 VSUBS 0.007047f
C78 B.n50 VSUBS 0.007047f
C79 B.n51 VSUBS 0.007047f
C80 B.n52 VSUBS 0.007047f
C81 B.n53 VSUBS 0.007047f
C82 B.n54 VSUBS 0.007047f
C83 B.n55 VSUBS 0.007047f
C84 B.n56 VSUBS 0.007047f
C85 B.n57 VSUBS 0.007047f
C86 B.n58 VSUBS 0.007047f
C87 B.n59 VSUBS 0.007047f
C88 B.n60 VSUBS 0.007047f
C89 B.n61 VSUBS 0.007047f
C90 B.t2 VSUBS 0.387793f
C91 B.t1 VSUBS 0.432765f
C92 B.t0 VSUBS 3.21651f
C93 B.n62 VSUBS 0.691244f
C94 B.n63 VSUBS 0.352268f
C95 B.n64 VSUBS 0.007047f
C96 B.n65 VSUBS 0.007047f
C97 B.n66 VSUBS 0.007047f
C98 B.n67 VSUBS 0.007047f
C99 B.t8 VSUBS 0.387797f
C100 B.t7 VSUBS 0.432768f
C101 B.t6 VSUBS 3.21651f
C102 B.n68 VSUBS 0.691241f
C103 B.n69 VSUBS 0.352264f
C104 B.n70 VSUBS 0.016328f
C105 B.n71 VSUBS 0.007047f
C106 B.n72 VSUBS 0.007047f
C107 B.n73 VSUBS 0.007047f
C108 B.n74 VSUBS 0.007047f
C109 B.n75 VSUBS 0.007047f
C110 B.n76 VSUBS 0.007047f
C111 B.n77 VSUBS 0.007047f
C112 B.n78 VSUBS 0.007047f
C113 B.n79 VSUBS 0.007047f
C114 B.n80 VSUBS 0.007047f
C115 B.n81 VSUBS 0.007047f
C116 B.n82 VSUBS 0.007047f
C117 B.n83 VSUBS 0.007047f
C118 B.n84 VSUBS 0.007047f
C119 B.n85 VSUBS 0.007047f
C120 B.n86 VSUBS 0.007047f
C121 B.n87 VSUBS 0.007047f
C122 B.n88 VSUBS 0.007047f
C123 B.n89 VSUBS 0.007047f
C124 B.n90 VSUBS 0.007047f
C125 B.n91 VSUBS 0.007047f
C126 B.n92 VSUBS 0.007047f
C127 B.n93 VSUBS 0.007047f
C128 B.n94 VSUBS 0.007047f
C129 B.n95 VSUBS 0.007047f
C130 B.n96 VSUBS 0.007047f
C131 B.n97 VSUBS 0.007047f
C132 B.n98 VSUBS 0.007047f
C133 B.n99 VSUBS 0.007047f
C134 B.n100 VSUBS 0.007047f
C135 B.n101 VSUBS 0.007047f
C136 B.n102 VSUBS 0.01718f
C137 B.n103 VSUBS 0.007047f
C138 B.n104 VSUBS 0.007047f
C139 B.n105 VSUBS 0.007047f
C140 B.n106 VSUBS 0.007047f
C141 B.n107 VSUBS 0.007047f
C142 B.n108 VSUBS 0.007047f
C143 B.n109 VSUBS 0.007047f
C144 B.n110 VSUBS 0.007047f
C145 B.n111 VSUBS 0.007047f
C146 B.n112 VSUBS 0.007047f
C147 B.n113 VSUBS 0.007047f
C148 B.n114 VSUBS 0.007047f
C149 B.n115 VSUBS 0.007047f
C150 B.n116 VSUBS 0.007047f
C151 B.n117 VSUBS 0.007047f
C152 B.n118 VSUBS 0.007047f
C153 B.n119 VSUBS 0.007047f
C154 B.n120 VSUBS 0.007047f
C155 B.n121 VSUBS 0.007047f
C156 B.n122 VSUBS 0.007047f
C157 B.n123 VSUBS 0.007047f
C158 B.n124 VSUBS 0.007047f
C159 B.n125 VSUBS 0.007047f
C160 B.n126 VSUBS 0.007047f
C161 B.n127 VSUBS 0.007047f
C162 B.n128 VSUBS 0.007047f
C163 B.n129 VSUBS 0.007047f
C164 B.n130 VSUBS 0.007047f
C165 B.n131 VSUBS 0.007047f
C166 B.n132 VSUBS 0.007047f
C167 B.n133 VSUBS 0.007047f
C168 B.n134 VSUBS 0.007047f
C169 B.n135 VSUBS 0.007047f
C170 B.n136 VSUBS 0.007047f
C171 B.n137 VSUBS 0.007047f
C172 B.n138 VSUBS 0.007047f
C173 B.n139 VSUBS 0.007047f
C174 B.n140 VSUBS 0.007047f
C175 B.n141 VSUBS 0.007047f
C176 B.n142 VSUBS 0.007047f
C177 B.n143 VSUBS 0.007047f
C178 B.n144 VSUBS 0.007047f
C179 B.n145 VSUBS 0.007047f
C180 B.n146 VSUBS 0.007047f
C181 B.n147 VSUBS 0.007047f
C182 B.n148 VSUBS 0.007047f
C183 B.n149 VSUBS 0.007047f
C184 B.n150 VSUBS 0.007047f
C185 B.n151 VSUBS 0.007047f
C186 B.n152 VSUBS 0.007047f
C187 B.n153 VSUBS 0.007047f
C188 B.n154 VSUBS 0.007047f
C189 B.n155 VSUBS 0.007047f
C190 B.n156 VSUBS 0.007047f
C191 B.n157 VSUBS 0.016346f
C192 B.n158 VSUBS 0.007047f
C193 B.n159 VSUBS 0.007047f
C194 B.n160 VSUBS 0.007047f
C195 B.n161 VSUBS 0.007047f
C196 B.n162 VSUBS 0.007047f
C197 B.n163 VSUBS 0.007047f
C198 B.n164 VSUBS 0.007047f
C199 B.n165 VSUBS 0.007047f
C200 B.n166 VSUBS 0.007047f
C201 B.n167 VSUBS 0.007047f
C202 B.n168 VSUBS 0.007047f
C203 B.n169 VSUBS 0.007047f
C204 B.n170 VSUBS 0.007047f
C205 B.n171 VSUBS 0.007047f
C206 B.n172 VSUBS 0.007047f
C207 B.n173 VSUBS 0.007047f
C208 B.n174 VSUBS 0.007047f
C209 B.n175 VSUBS 0.007047f
C210 B.n176 VSUBS 0.007047f
C211 B.n177 VSUBS 0.007047f
C212 B.n178 VSUBS 0.007047f
C213 B.n179 VSUBS 0.007047f
C214 B.n180 VSUBS 0.007047f
C215 B.n181 VSUBS 0.007047f
C216 B.n182 VSUBS 0.007047f
C217 B.n183 VSUBS 0.007047f
C218 B.n184 VSUBS 0.007047f
C219 B.n185 VSUBS 0.007047f
C220 B.n186 VSUBS 0.007047f
C221 B.n187 VSUBS 0.007047f
C222 B.n188 VSUBS 0.007047f
C223 B.n189 VSUBS 0.007047f
C224 B.t4 VSUBS 0.387797f
C225 B.t5 VSUBS 0.432768f
C226 B.t3 VSUBS 3.21651f
C227 B.n190 VSUBS 0.691241f
C228 B.n191 VSUBS 0.352264f
C229 B.n192 VSUBS 0.007047f
C230 B.n193 VSUBS 0.007047f
C231 B.n194 VSUBS 0.007047f
C232 B.n195 VSUBS 0.007047f
C233 B.t10 VSUBS 0.387793f
C234 B.t11 VSUBS 0.432765f
C235 B.t9 VSUBS 3.21651f
C236 B.n196 VSUBS 0.691244f
C237 B.n197 VSUBS 0.352268f
C238 B.n198 VSUBS 0.016328f
C239 B.n199 VSUBS 0.007047f
C240 B.n200 VSUBS 0.007047f
C241 B.n201 VSUBS 0.007047f
C242 B.n202 VSUBS 0.007047f
C243 B.n203 VSUBS 0.007047f
C244 B.n204 VSUBS 0.007047f
C245 B.n205 VSUBS 0.007047f
C246 B.n206 VSUBS 0.007047f
C247 B.n207 VSUBS 0.007047f
C248 B.n208 VSUBS 0.007047f
C249 B.n209 VSUBS 0.007047f
C250 B.n210 VSUBS 0.007047f
C251 B.n211 VSUBS 0.007047f
C252 B.n212 VSUBS 0.007047f
C253 B.n213 VSUBS 0.007047f
C254 B.n214 VSUBS 0.007047f
C255 B.n215 VSUBS 0.007047f
C256 B.n216 VSUBS 0.007047f
C257 B.n217 VSUBS 0.007047f
C258 B.n218 VSUBS 0.007047f
C259 B.n219 VSUBS 0.007047f
C260 B.n220 VSUBS 0.007047f
C261 B.n221 VSUBS 0.007047f
C262 B.n222 VSUBS 0.007047f
C263 B.n223 VSUBS 0.007047f
C264 B.n224 VSUBS 0.007047f
C265 B.n225 VSUBS 0.007047f
C266 B.n226 VSUBS 0.007047f
C267 B.n227 VSUBS 0.007047f
C268 B.n228 VSUBS 0.007047f
C269 B.n229 VSUBS 0.007047f
C270 B.n230 VSUBS 0.016346f
C271 B.n231 VSUBS 0.007047f
C272 B.n232 VSUBS 0.007047f
C273 B.n233 VSUBS 0.007047f
C274 B.n234 VSUBS 0.007047f
C275 B.n235 VSUBS 0.007047f
C276 B.n236 VSUBS 0.007047f
C277 B.n237 VSUBS 0.007047f
C278 B.n238 VSUBS 0.007047f
C279 B.n239 VSUBS 0.007047f
C280 B.n240 VSUBS 0.007047f
C281 B.n241 VSUBS 0.007047f
C282 B.n242 VSUBS 0.007047f
C283 B.n243 VSUBS 0.007047f
C284 B.n244 VSUBS 0.007047f
C285 B.n245 VSUBS 0.007047f
C286 B.n246 VSUBS 0.007047f
C287 B.n247 VSUBS 0.007047f
C288 B.n248 VSUBS 0.007047f
C289 B.n249 VSUBS 0.007047f
C290 B.n250 VSUBS 0.007047f
C291 B.n251 VSUBS 0.007047f
C292 B.n252 VSUBS 0.007047f
C293 B.n253 VSUBS 0.007047f
C294 B.n254 VSUBS 0.007047f
C295 B.n255 VSUBS 0.007047f
C296 B.n256 VSUBS 0.007047f
C297 B.n257 VSUBS 0.007047f
C298 B.n258 VSUBS 0.007047f
C299 B.n259 VSUBS 0.007047f
C300 B.n260 VSUBS 0.007047f
C301 B.n261 VSUBS 0.007047f
C302 B.n262 VSUBS 0.007047f
C303 B.n263 VSUBS 0.007047f
C304 B.n264 VSUBS 0.007047f
C305 B.n265 VSUBS 0.007047f
C306 B.n266 VSUBS 0.007047f
C307 B.n267 VSUBS 0.007047f
C308 B.n268 VSUBS 0.007047f
C309 B.n269 VSUBS 0.007047f
C310 B.n270 VSUBS 0.007047f
C311 B.n271 VSUBS 0.007047f
C312 B.n272 VSUBS 0.007047f
C313 B.n273 VSUBS 0.007047f
C314 B.n274 VSUBS 0.007047f
C315 B.n275 VSUBS 0.007047f
C316 B.n276 VSUBS 0.007047f
C317 B.n277 VSUBS 0.007047f
C318 B.n278 VSUBS 0.007047f
C319 B.n279 VSUBS 0.007047f
C320 B.n280 VSUBS 0.007047f
C321 B.n281 VSUBS 0.007047f
C322 B.n282 VSUBS 0.007047f
C323 B.n283 VSUBS 0.007047f
C324 B.n284 VSUBS 0.007047f
C325 B.n285 VSUBS 0.007047f
C326 B.n286 VSUBS 0.007047f
C327 B.n287 VSUBS 0.007047f
C328 B.n288 VSUBS 0.007047f
C329 B.n289 VSUBS 0.007047f
C330 B.n290 VSUBS 0.007047f
C331 B.n291 VSUBS 0.007047f
C332 B.n292 VSUBS 0.007047f
C333 B.n293 VSUBS 0.007047f
C334 B.n294 VSUBS 0.007047f
C335 B.n295 VSUBS 0.007047f
C336 B.n296 VSUBS 0.007047f
C337 B.n297 VSUBS 0.007047f
C338 B.n298 VSUBS 0.007047f
C339 B.n299 VSUBS 0.007047f
C340 B.n300 VSUBS 0.007047f
C341 B.n301 VSUBS 0.007047f
C342 B.n302 VSUBS 0.007047f
C343 B.n303 VSUBS 0.007047f
C344 B.n304 VSUBS 0.007047f
C345 B.n305 VSUBS 0.007047f
C346 B.n306 VSUBS 0.007047f
C347 B.n307 VSUBS 0.007047f
C348 B.n308 VSUBS 0.007047f
C349 B.n309 VSUBS 0.007047f
C350 B.n310 VSUBS 0.007047f
C351 B.n311 VSUBS 0.007047f
C352 B.n312 VSUBS 0.007047f
C353 B.n313 VSUBS 0.007047f
C354 B.n314 VSUBS 0.007047f
C355 B.n315 VSUBS 0.007047f
C356 B.n316 VSUBS 0.007047f
C357 B.n317 VSUBS 0.007047f
C358 B.n318 VSUBS 0.007047f
C359 B.n319 VSUBS 0.007047f
C360 B.n320 VSUBS 0.007047f
C361 B.n321 VSUBS 0.007047f
C362 B.n322 VSUBS 0.007047f
C363 B.n323 VSUBS 0.007047f
C364 B.n324 VSUBS 0.007047f
C365 B.n325 VSUBS 0.007047f
C366 B.n326 VSUBS 0.007047f
C367 B.n327 VSUBS 0.007047f
C368 B.n328 VSUBS 0.007047f
C369 B.n329 VSUBS 0.007047f
C370 B.n330 VSUBS 0.007047f
C371 B.n331 VSUBS 0.007047f
C372 B.n332 VSUBS 0.007047f
C373 B.n333 VSUBS 0.007047f
C374 B.n334 VSUBS 0.007047f
C375 B.n335 VSUBS 0.007047f
C376 B.n336 VSUBS 0.007047f
C377 B.n337 VSUBS 0.016346f
C378 B.n338 VSUBS 0.016611f
C379 B.n339 VSUBS 0.016611f
C380 B.n340 VSUBS 0.007047f
C381 B.n341 VSUBS 0.007047f
C382 B.n342 VSUBS 0.007047f
C383 B.n343 VSUBS 0.007047f
C384 B.n344 VSUBS 0.007047f
C385 B.n345 VSUBS 0.007047f
C386 B.n346 VSUBS 0.007047f
C387 B.n347 VSUBS 0.007047f
C388 B.n348 VSUBS 0.007047f
C389 B.n349 VSUBS 0.007047f
C390 B.n350 VSUBS 0.007047f
C391 B.n351 VSUBS 0.007047f
C392 B.n352 VSUBS 0.007047f
C393 B.n353 VSUBS 0.007047f
C394 B.n354 VSUBS 0.007047f
C395 B.n355 VSUBS 0.007047f
C396 B.n356 VSUBS 0.007047f
C397 B.n357 VSUBS 0.007047f
C398 B.n358 VSUBS 0.007047f
C399 B.n359 VSUBS 0.007047f
C400 B.n360 VSUBS 0.007047f
C401 B.n361 VSUBS 0.007047f
C402 B.n362 VSUBS 0.007047f
C403 B.n363 VSUBS 0.007047f
C404 B.n364 VSUBS 0.007047f
C405 B.n365 VSUBS 0.007047f
C406 B.n366 VSUBS 0.007047f
C407 B.n367 VSUBS 0.007047f
C408 B.n368 VSUBS 0.007047f
C409 B.n369 VSUBS 0.007047f
C410 B.n370 VSUBS 0.007047f
C411 B.n371 VSUBS 0.007047f
C412 B.n372 VSUBS 0.007047f
C413 B.n373 VSUBS 0.007047f
C414 B.n374 VSUBS 0.007047f
C415 B.n375 VSUBS 0.007047f
C416 B.n376 VSUBS 0.007047f
C417 B.n377 VSUBS 0.007047f
C418 B.n378 VSUBS 0.007047f
C419 B.n379 VSUBS 0.007047f
C420 B.n380 VSUBS 0.007047f
C421 B.n381 VSUBS 0.007047f
C422 B.n382 VSUBS 0.007047f
C423 B.n383 VSUBS 0.007047f
C424 B.n384 VSUBS 0.007047f
C425 B.n385 VSUBS 0.007047f
C426 B.n386 VSUBS 0.007047f
C427 B.n387 VSUBS 0.007047f
C428 B.n388 VSUBS 0.007047f
C429 B.n389 VSUBS 0.007047f
C430 B.n390 VSUBS 0.007047f
C431 B.n391 VSUBS 0.007047f
C432 B.n392 VSUBS 0.007047f
C433 B.n393 VSUBS 0.007047f
C434 B.n394 VSUBS 0.007047f
C435 B.n395 VSUBS 0.007047f
C436 B.n396 VSUBS 0.007047f
C437 B.n397 VSUBS 0.007047f
C438 B.n398 VSUBS 0.007047f
C439 B.n399 VSUBS 0.007047f
C440 B.n400 VSUBS 0.007047f
C441 B.n401 VSUBS 0.007047f
C442 B.n402 VSUBS 0.007047f
C443 B.n403 VSUBS 0.007047f
C444 B.n404 VSUBS 0.007047f
C445 B.n405 VSUBS 0.007047f
C446 B.n406 VSUBS 0.007047f
C447 B.n407 VSUBS 0.007047f
C448 B.n408 VSUBS 0.007047f
C449 B.n409 VSUBS 0.007047f
C450 B.n410 VSUBS 0.007047f
C451 B.n411 VSUBS 0.007047f
C452 B.n412 VSUBS 0.007047f
C453 B.n413 VSUBS 0.007047f
C454 B.n414 VSUBS 0.007047f
C455 B.n415 VSUBS 0.007047f
C456 B.n416 VSUBS 0.007047f
C457 B.n417 VSUBS 0.007047f
C458 B.n418 VSUBS 0.007047f
C459 B.n419 VSUBS 0.007047f
C460 B.n420 VSUBS 0.007047f
C461 B.n421 VSUBS 0.007047f
C462 B.n422 VSUBS 0.007047f
C463 B.n423 VSUBS 0.007047f
C464 B.n424 VSUBS 0.007047f
C465 B.n425 VSUBS 0.007047f
C466 B.n426 VSUBS 0.007047f
C467 B.n427 VSUBS 0.007047f
C468 B.n428 VSUBS 0.007047f
C469 B.n429 VSUBS 0.007047f
C470 B.n430 VSUBS 0.007047f
C471 B.n431 VSUBS 0.006633f
C472 B.n432 VSUBS 0.007047f
C473 B.n433 VSUBS 0.007047f
C474 B.n434 VSUBS 0.003938f
C475 B.n435 VSUBS 0.007047f
C476 B.n436 VSUBS 0.007047f
C477 B.n437 VSUBS 0.007047f
C478 B.n438 VSUBS 0.007047f
C479 B.n439 VSUBS 0.007047f
C480 B.n440 VSUBS 0.007047f
C481 B.n441 VSUBS 0.007047f
C482 B.n442 VSUBS 0.007047f
C483 B.n443 VSUBS 0.007047f
C484 B.n444 VSUBS 0.007047f
C485 B.n445 VSUBS 0.007047f
C486 B.n446 VSUBS 0.007047f
C487 B.n447 VSUBS 0.003938f
C488 B.n448 VSUBS 0.016328f
C489 B.n449 VSUBS 0.006633f
C490 B.n450 VSUBS 0.007047f
C491 B.n451 VSUBS 0.007047f
C492 B.n452 VSUBS 0.007047f
C493 B.n453 VSUBS 0.007047f
C494 B.n454 VSUBS 0.007047f
C495 B.n455 VSUBS 0.007047f
C496 B.n456 VSUBS 0.007047f
C497 B.n457 VSUBS 0.007047f
C498 B.n458 VSUBS 0.007047f
C499 B.n459 VSUBS 0.007047f
C500 B.n460 VSUBS 0.007047f
C501 B.n461 VSUBS 0.007047f
C502 B.n462 VSUBS 0.007047f
C503 B.n463 VSUBS 0.007047f
C504 B.n464 VSUBS 0.007047f
C505 B.n465 VSUBS 0.007047f
C506 B.n466 VSUBS 0.007047f
C507 B.n467 VSUBS 0.007047f
C508 B.n468 VSUBS 0.007047f
C509 B.n469 VSUBS 0.007047f
C510 B.n470 VSUBS 0.007047f
C511 B.n471 VSUBS 0.007047f
C512 B.n472 VSUBS 0.007047f
C513 B.n473 VSUBS 0.007047f
C514 B.n474 VSUBS 0.007047f
C515 B.n475 VSUBS 0.007047f
C516 B.n476 VSUBS 0.007047f
C517 B.n477 VSUBS 0.007047f
C518 B.n478 VSUBS 0.007047f
C519 B.n479 VSUBS 0.007047f
C520 B.n480 VSUBS 0.007047f
C521 B.n481 VSUBS 0.007047f
C522 B.n482 VSUBS 0.007047f
C523 B.n483 VSUBS 0.007047f
C524 B.n484 VSUBS 0.007047f
C525 B.n485 VSUBS 0.007047f
C526 B.n486 VSUBS 0.007047f
C527 B.n487 VSUBS 0.007047f
C528 B.n488 VSUBS 0.007047f
C529 B.n489 VSUBS 0.007047f
C530 B.n490 VSUBS 0.007047f
C531 B.n491 VSUBS 0.007047f
C532 B.n492 VSUBS 0.007047f
C533 B.n493 VSUBS 0.007047f
C534 B.n494 VSUBS 0.007047f
C535 B.n495 VSUBS 0.007047f
C536 B.n496 VSUBS 0.007047f
C537 B.n497 VSUBS 0.007047f
C538 B.n498 VSUBS 0.007047f
C539 B.n499 VSUBS 0.007047f
C540 B.n500 VSUBS 0.007047f
C541 B.n501 VSUBS 0.007047f
C542 B.n502 VSUBS 0.007047f
C543 B.n503 VSUBS 0.007047f
C544 B.n504 VSUBS 0.007047f
C545 B.n505 VSUBS 0.007047f
C546 B.n506 VSUBS 0.007047f
C547 B.n507 VSUBS 0.007047f
C548 B.n508 VSUBS 0.007047f
C549 B.n509 VSUBS 0.007047f
C550 B.n510 VSUBS 0.007047f
C551 B.n511 VSUBS 0.007047f
C552 B.n512 VSUBS 0.007047f
C553 B.n513 VSUBS 0.007047f
C554 B.n514 VSUBS 0.007047f
C555 B.n515 VSUBS 0.007047f
C556 B.n516 VSUBS 0.007047f
C557 B.n517 VSUBS 0.007047f
C558 B.n518 VSUBS 0.007047f
C559 B.n519 VSUBS 0.007047f
C560 B.n520 VSUBS 0.007047f
C561 B.n521 VSUBS 0.007047f
C562 B.n522 VSUBS 0.007047f
C563 B.n523 VSUBS 0.007047f
C564 B.n524 VSUBS 0.007047f
C565 B.n525 VSUBS 0.007047f
C566 B.n526 VSUBS 0.007047f
C567 B.n527 VSUBS 0.007047f
C568 B.n528 VSUBS 0.007047f
C569 B.n529 VSUBS 0.007047f
C570 B.n530 VSUBS 0.007047f
C571 B.n531 VSUBS 0.007047f
C572 B.n532 VSUBS 0.007047f
C573 B.n533 VSUBS 0.007047f
C574 B.n534 VSUBS 0.007047f
C575 B.n535 VSUBS 0.007047f
C576 B.n536 VSUBS 0.007047f
C577 B.n537 VSUBS 0.007047f
C578 B.n538 VSUBS 0.007047f
C579 B.n539 VSUBS 0.007047f
C580 B.n540 VSUBS 0.007047f
C581 B.n541 VSUBS 0.007047f
C582 B.n542 VSUBS 0.016611f
C583 B.n543 VSUBS 0.016611f
C584 B.n544 VSUBS 0.016346f
C585 B.n545 VSUBS 0.007047f
C586 B.n546 VSUBS 0.007047f
C587 B.n547 VSUBS 0.007047f
C588 B.n548 VSUBS 0.007047f
C589 B.n549 VSUBS 0.007047f
C590 B.n550 VSUBS 0.007047f
C591 B.n551 VSUBS 0.007047f
C592 B.n552 VSUBS 0.007047f
C593 B.n553 VSUBS 0.007047f
C594 B.n554 VSUBS 0.007047f
C595 B.n555 VSUBS 0.007047f
C596 B.n556 VSUBS 0.007047f
C597 B.n557 VSUBS 0.007047f
C598 B.n558 VSUBS 0.007047f
C599 B.n559 VSUBS 0.007047f
C600 B.n560 VSUBS 0.007047f
C601 B.n561 VSUBS 0.007047f
C602 B.n562 VSUBS 0.007047f
C603 B.n563 VSUBS 0.007047f
C604 B.n564 VSUBS 0.007047f
C605 B.n565 VSUBS 0.007047f
C606 B.n566 VSUBS 0.007047f
C607 B.n567 VSUBS 0.007047f
C608 B.n568 VSUBS 0.007047f
C609 B.n569 VSUBS 0.007047f
C610 B.n570 VSUBS 0.007047f
C611 B.n571 VSUBS 0.007047f
C612 B.n572 VSUBS 0.007047f
C613 B.n573 VSUBS 0.007047f
C614 B.n574 VSUBS 0.007047f
C615 B.n575 VSUBS 0.007047f
C616 B.n576 VSUBS 0.007047f
C617 B.n577 VSUBS 0.007047f
C618 B.n578 VSUBS 0.007047f
C619 B.n579 VSUBS 0.007047f
C620 B.n580 VSUBS 0.007047f
C621 B.n581 VSUBS 0.007047f
C622 B.n582 VSUBS 0.007047f
C623 B.n583 VSUBS 0.007047f
C624 B.n584 VSUBS 0.007047f
C625 B.n585 VSUBS 0.007047f
C626 B.n586 VSUBS 0.007047f
C627 B.n587 VSUBS 0.007047f
C628 B.n588 VSUBS 0.007047f
C629 B.n589 VSUBS 0.007047f
C630 B.n590 VSUBS 0.007047f
C631 B.n591 VSUBS 0.007047f
C632 B.n592 VSUBS 0.007047f
C633 B.n593 VSUBS 0.007047f
C634 B.n594 VSUBS 0.007047f
C635 B.n595 VSUBS 0.007047f
C636 B.n596 VSUBS 0.007047f
C637 B.n597 VSUBS 0.007047f
C638 B.n598 VSUBS 0.007047f
C639 B.n599 VSUBS 0.007047f
C640 B.n600 VSUBS 0.007047f
C641 B.n601 VSUBS 0.007047f
C642 B.n602 VSUBS 0.007047f
C643 B.n603 VSUBS 0.007047f
C644 B.n604 VSUBS 0.007047f
C645 B.n605 VSUBS 0.007047f
C646 B.n606 VSUBS 0.007047f
C647 B.n607 VSUBS 0.007047f
C648 B.n608 VSUBS 0.007047f
C649 B.n609 VSUBS 0.007047f
C650 B.n610 VSUBS 0.007047f
C651 B.n611 VSUBS 0.007047f
C652 B.n612 VSUBS 0.007047f
C653 B.n613 VSUBS 0.007047f
C654 B.n614 VSUBS 0.007047f
C655 B.n615 VSUBS 0.007047f
C656 B.n616 VSUBS 0.007047f
C657 B.n617 VSUBS 0.007047f
C658 B.n618 VSUBS 0.007047f
C659 B.n619 VSUBS 0.007047f
C660 B.n620 VSUBS 0.007047f
C661 B.n621 VSUBS 0.007047f
C662 B.n622 VSUBS 0.007047f
C663 B.n623 VSUBS 0.007047f
C664 B.n624 VSUBS 0.007047f
C665 B.n625 VSUBS 0.007047f
C666 B.n626 VSUBS 0.007047f
C667 B.n627 VSUBS 0.007047f
C668 B.n628 VSUBS 0.007047f
C669 B.n629 VSUBS 0.007047f
C670 B.n630 VSUBS 0.007047f
C671 B.n631 VSUBS 0.007047f
C672 B.n632 VSUBS 0.007047f
C673 B.n633 VSUBS 0.007047f
C674 B.n634 VSUBS 0.007047f
C675 B.n635 VSUBS 0.007047f
C676 B.n636 VSUBS 0.007047f
C677 B.n637 VSUBS 0.007047f
C678 B.n638 VSUBS 0.007047f
C679 B.n639 VSUBS 0.007047f
C680 B.n640 VSUBS 0.007047f
C681 B.n641 VSUBS 0.007047f
C682 B.n642 VSUBS 0.007047f
C683 B.n643 VSUBS 0.007047f
C684 B.n644 VSUBS 0.007047f
C685 B.n645 VSUBS 0.007047f
C686 B.n646 VSUBS 0.007047f
C687 B.n647 VSUBS 0.007047f
C688 B.n648 VSUBS 0.007047f
C689 B.n649 VSUBS 0.007047f
C690 B.n650 VSUBS 0.007047f
C691 B.n651 VSUBS 0.007047f
C692 B.n652 VSUBS 0.007047f
C693 B.n653 VSUBS 0.007047f
C694 B.n654 VSUBS 0.007047f
C695 B.n655 VSUBS 0.007047f
C696 B.n656 VSUBS 0.007047f
C697 B.n657 VSUBS 0.007047f
C698 B.n658 VSUBS 0.007047f
C699 B.n659 VSUBS 0.007047f
C700 B.n660 VSUBS 0.007047f
C701 B.n661 VSUBS 0.007047f
C702 B.n662 VSUBS 0.007047f
C703 B.n663 VSUBS 0.007047f
C704 B.n664 VSUBS 0.007047f
C705 B.n665 VSUBS 0.007047f
C706 B.n666 VSUBS 0.007047f
C707 B.n667 VSUBS 0.007047f
C708 B.n668 VSUBS 0.007047f
C709 B.n669 VSUBS 0.007047f
C710 B.n670 VSUBS 0.007047f
C711 B.n671 VSUBS 0.007047f
C712 B.n672 VSUBS 0.007047f
C713 B.n673 VSUBS 0.007047f
C714 B.n674 VSUBS 0.007047f
C715 B.n675 VSUBS 0.007047f
C716 B.n676 VSUBS 0.007047f
C717 B.n677 VSUBS 0.007047f
C718 B.n678 VSUBS 0.007047f
C719 B.n679 VSUBS 0.007047f
C720 B.n680 VSUBS 0.007047f
C721 B.n681 VSUBS 0.007047f
C722 B.n682 VSUBS 0.007047f
C723 B.n683 VSUBS 0.007047f
C724 B.n684 VSUBS 0.007047f
C725 B.n685 VSUBS 0.007047f
C726 B.n686 VSUBS 0.007047f
C727 B.n687 VSUBS 0.007047f
C728 B.n688 VSUBS 0.007047f
C729 B.n689 VSUBS 0.007047f
C730 B.n690 VSUBS 0.007047f
C731 B.n691 VSUBS 0.007047f
C732 B.n692 VSUBS 0.007047f
C733 B.n693 VSUBS 0.007047f
C734 B.n694 VSUBS 0.007047f
C735 B.n695 VSUBS 0.007047f
C736 B.n696 VSUBS 0.007047f
C737 B.n697 VSUBS 0.007047f
C738 B.n698 VSUBS 0.007047f
C739 B.n699 VSUBS 0.007047f
C740 B.n700 VSUBS 0.007047f
C741 B.n701 VSUBS 0.007047f
C742 B.n702 VSUBS 0.007047f
C743 B.n703 VSUBS 0.007047f
C744 B.n704 VSUBS 0.007047f
C745 B.n705 VSUBS 0.007047f
C746 B.n706 VSUBS 0.007047f
C747 B.n707 VSUBS 0.007047f
C748 B.n708 VSUBS 0.007047f
C749 B.n709 VSUBS 0.016346f
C750 B.n710 VSUBS 0.016611f
C751 B.n711 VSUBS 0.015777f
C752 B.n712 VSUBS 0.007047f
C753 B.n713 VSUBS 0.007047f
C754 B.n714 VSUBS 0.007047f
C755 B.n715 VSUBS 0.007047f
C756 B.n716 VSUBS 0.007047f
C757 B.n717 VSUBS 0.007047f
C758 B.n718 VSUBS 0.007047f
C759 B.n719 VSUBS 0.007047f
C760 B.n720 VSUBS 0.007047f
C761 B.n721 VSUBS 0.007047f
C762 B.n722 VSUBS 0.007047f
C763 B.n723 VSUBS 0.007047f
C764 B.n724 VSUBS 0.007047f
C765 B.n725 VSUBS 0.007047f
C766 B.n726 VSUBS 0.007047f
C767 B.n727 VSUBS 0.007047f
C768 B.n728 VSUBS 0.007047f
C769 B.n729 VSUBS 0.007047f
C770 B.n730 VSUBS 0.007047f
C771 B.n731 VSUBS 0.007047f
C772 B.n732 VSUBS 0.007047f
C773 B.n733 VSUBS 0.007047f
C774 B.n734 VSUBS 0.007047f
C775 B.n735 VSUBS 0.007047f
C776 B.n736 VSUBS 0.007047f
C777 B.n737 VSUBS 0.007047f
C778 B.n738 VSUBS 0.007047f
C779 B.n739 VSUBS 0.007047f
C780 B.n740 VSUBS 0.007047f
C781 B.n741 VSUBS 0.007047f
C782 B.n742 VSUBS 0.007047f
C783 B.n743 VSUBS 0.007047f
C784 B.n744 VSUBS 0.007047f
C785 B.n745 VSUBS 0.007047f
C786 B.n746 VSUBS 0.007047f
C787 B.n747 VSUBS 0.007047f
C788 B.n748 VSUBS 0.007047f
C789 B.n749 VSUBS 0.007047f
C790 B.n750 VSUBS 0.007047f
C791 B.n751 VSUBS 0.007047f
C792 B.n752 VSUBS 0.007047f
C793 B.n753 VSUBS 0.007047f
C794 B.n754 VSUBS 0.007047f
C795 B.n755 VSUBS 0.007047f
C796 B.n756 VSUBS 0.007047f
C797 B.n757 VSUBS 0.007047f
C798 B.n758 VSUBS 0.007047f
C799 B.n759 VSUBS 0.007047f
C800 B.n760 VSUBS 0.007047f
C801 B.n761 VSUBS 0.007047f
C802 B.n762 VSUBS 0.007047f
C803 B.n763 VSUBS 0.007047f
C804 B.n764 VSUBS 0.007047f
C805 B.n765 VSUBS 0.007047f
C806 B.n766 VSUBS 0.007047f
C807 B.n767 VSUBS 0.007047f
C808 B.n768 VSUBS 0.007047f
C809 B.n769 VSUBS 0.007047f
C810 B.n770 VSUBS 0.007047f
C811 B.n771 VSUBS 0.007047f
C812 B.n772 VSUBS 0.007047f
C813 B.n773 VSUBS 0.007047f
C814 B.n774 VSUBS 0.007047f
C815 B.n775 VSUBS 0.007047f
C816 B.n776 VSUBS 0.007047f
C817 B.n777 VSUBS 0.007047f
C818 B.n778 VSUBS 0.007047f
C819 B.n779 VSUBS 0.007047f
C820 B.n780 VSUBS 0.007047f
C821 B.n781 VSUBS 0.007047f
C822 B.n782 VSUBS 0.007047f
C823 B.n783 VSUBS 0.007047f
C824 B.n784 VSUBS 0.007047f
C825 B.n785 VSUBS 0.007047f
C826 B.n786 VSUBS 0.007047f
C827 B.n787 VSUBS 0.007047f
C828 B.n788 VSUBS 0.007047f
C829 B.n789 VSUBS 0.007047f
C830 B.n790 VSUBS 0.007047f
C831 B.n791 VSUBS 0.007047f
C832 B.n792 VSUBS 0.007047f
C833 B.n793 VSUBS 0.007047f
C834 B.n794 VSUBS 0.007047f
C835 B.n795 VSUBS 0.007047f
C836 B.n796 VSUBS 0.007047f
C837 B.n797 VSUBS 0.007047f
C838 B.n798 VSUBS 0.007047f
C839 B.n799 VSUBS 0.007047f
C840 B.n800 VSUBS 0.007047f
C841 B.n801 VSUBS 0.007047f
C842 B.n802 VSUBS 0.007047f
C843 B.n803 VSUBS 0.006633f
C844 B.n804 VSUBS 0.007047f
C845 B.n805 VSUBS 0.007047f
C846 B.n806 VSUBS 0.003938f
C847 B.n807 VSUBS 0.007047f
C848 B.n808 VSUBS 0.007047f
C849 B.n809 VSUBS 0.007047f
C850 B.n810 VSUBS 0.007047f
C851 B.n811 VSUBS 0.007047f
C852 B.n812 VSUBS 0.007047f
C853 B.n813 VSUBS 0.007047f
C854 B.n814 VSUBS 0.007047f
C855 B.n815 VSUBS 0.007047f
C856 B.n816 VSUBS 0.007047f
C857 B.n817 VSUBS 0.007047f
C858 B.n818 VSUBS 0.007047f
C859 B.n819 VSUBS 0.003938f
C860 B.n820 VSUBS 0.016328f
C861 B.n821 VSUBS 0.006633f
C862 B.n822 VSUBS 0.007047f
C863 B.n823 VSUBS 0.007047f
C864 B.n824 VSUBS 0.007047f
C865 B.n825 VSUBS 0.007047f
C866 B.n826 VSUBS 0.007047f
C867 B.n827 VSUBS 0.007047f
C868 B.n828 VSUBS 0.007047f
C869 B.n829 VSUBS 0.007047f
C870 B.n830 VSUBS 0.007047f
C871 B.n831 VSUBS 0.007047f
C872 B.n832 VSUBS 0.007047f
C873 B.n833 VSUBS 0.007047f
C874 B.n834 VSUBS 0.007047f
C875 B.n835 VSUBS 0.007047f
C876 B.n836 VSUBS 0.007047f
C877 B.n837 VSUBS 0.007047f
C878 B.n838 VSUBS 0.007047f
C879 B.n839 VSUBS 0.007047f
C880 B.n840 VSUBS 0.007047f
C881 B.n841 VSUBS 0.007047f
C882 B.n842 VSUBS 0.007047f
C883 B.n843 VSUBS 0.007047f
C884 B.n844 VSUBS 0.007047f
C885 B.n845 VSUBS 0.007047f
C886 B.n846 VSUBS 0.007047f
C887 B.n847 VSUBS 0.007047f
C888 B.n848 VSUBS 0.007047f
C889 B.n849 VSUBS 0.007047f
C890 B.n850 VSUBS 0.007047f
C891 B.n851 VSUBS 0.007047f
C892 B.n852 VSUBS 0.007047f
C893 B.n853 VSUBS 0.007047f
C894 B.n854 VSUBS 0.007047f
C895 B.n855 VSUBS 0.007047f
C896 B.n856 VSUBS 0.007047f
C897 B.n857 VSUBS 0.007047f
C898 B.n858 VSUBS 0.007047f
C899 B.n859 VSUBS 0.007047f
C900 B.n860 VSUBS 0.007047f
C901 B.n861 VSUBS 0.007047f
C902 B.n862 VSUBS 0.007047f
C903 B.n863 VSUBS 0.007047f
C904 B.n864 VSUBS 0.007047f
C905 B.n865 VSUBS 0.007047f
C906 B.n866 VSUBS 0.007047f
C907 B.n867 VSUBS 0.007047f
C908 B.n868 VSUBS 0.007047f
C909 B.n869 VSUBS 0.007047f
C910 B.n870 VSUBS 0.007047f
C911 B.n871 VSUBS 0.007047f
C912 B.n872 VSUBS 0.007047f
C913 B.n873 VSUBS 0.007047f
C914 B.n874 VSUBS 0.007047f
C915 B.n875 VSUBS 0.007047f
C916 B.n876 VSUBS 0.007047f
C917 B.n877 VSUBS 0.007047f
C918 B.n878 VSUBS 0.007047f
C919 B.n879 VSUBS 0.007047f
C920 B.n880 VSUBS 0.007047f
C921 B.n881 VSUBS 0.007047f
C922 B.n882 VSUBS 0.007047f
C923 B.n883 VSUBS 0.007047f
C924 B.n884 VSUBS 0.007047f
C925 B.n885 VSUBS 0.007047f
C926 B.n886 VSUBS 0.007047f
C927 B.n887 VSUBS 0.007047f
C928 B.n888 VSUBS 0.007047f
C929 B.n889 VSUBS 0.007047f
C930 B.n890 VSUBS 0.007047f
C931 B.n891 VSUBS 0.007047f
C932 B.n892 VSUBS 0.007047f
C933 B.n893 VSUBS 0.007047f
C934 B.n894 VSUBS 0.007047f
C935 B.n895 VSUBS 0.007047f
C936 B.n896 VSUBS 0.007047f
C937 B.n897 VSUBS 0.007047f
C938 B.n898 VSUBS 0.007047f
C939 B.n899 VSUBS 0.007047f
C940 B.n900 VSUBS 0.007047f
C941 B.n901 VSUBS 0.007047f
C942 B.n902 VSUBS 0.007047f
C943 B.n903 VSUBS 0.007047f
C944 B.n904 VSUBS 0.007047f
C945 B.n905 VSUBS 0.007047f
C946 B.n906 VSUBS 0.007047f
C947 B.n907 VSUBS 0.007047f
C948 B.n908 VSUBS 0.007047f
C949 B.n909 VSUBS 0.007047f
C950 B.n910 VSUBS 0.007047f
C951 B.n911 VSUBS 0.007047f
C952 B.n912 VSUBS 0.007047f
C953 B.n913 VSUBS 0.007047f
C954 B.n914 VSUBS 0.016611f
C955 B.n915 VSUBS 0.016611f
C956 B.n916 VSUBS 0.016346f
C957 B.n917 VSUBS 0.007047f
C958 B.n918 VSUBS 0.007047f
C959 B.n919 VSUBS 0.007047f
C960 B.n920 VSUBS 0.007047f
C961 B.n921 VSUBS 0.007047f
C962 B.n922 VSUBS 0.007047f
C963 B.n923 VSUBS 0.007047f
C964 B.n924 VSUBS 0.007047f
C965 B.n925 VSUBS 0.007047f
C966 B.n926 VSUBS 0.007047f
C967 B.n927 VSUBS 0.007047f
C968 B.n928 VSUBS 0.007047f
C969 B.n929 VSUBS 0.007047f
C970 B.n930 VSUBS 0.007047f
C971 B.n931 VSUBS 0.007047f
C972 B.n932 VSUBS 0.007047f
C973 B.n933 VSUBS 0.007047f
C974 B.n934 VSUBS 0.007047f
C975 B.n935 VSUBS 0.007047f
C976 B.n936 VSUBS 0.007047f
C977 B.n937 VSUBS 0.007047f
C978 B.n938 VSUBS 0.007047f
C979 B.n939 VSUBS 0.007047f
C980 B.n940 VSUBS 0.007047f
C981 B.n941 VSUBS 0.007047f
C982 B.n942 VSUBS 0.007047f
C983 B.n943 VSUBS 0.007047f
C984 B.n944 VSUBS 0.007047f
C985 B.n945 VSUBS 0.007047f
C986 B.n946 VSUBS 0.007047f
C987 B.n947 VSUBS 0.007047f
C988 B.n948 VSUBS 0.007047f
C989 B.n949 VSUBS 0.007047f
C990 B.n950 VSUBS 0.007047f
C991 B.n951 VSUBS 0.007047f
C992 B.n952 VSUBS 0.007047f
C993 B.n953 VSUBS 0.007047f
C994 B.n954 VSUBS 0.007047f
C995 B.n955 VSUBS 0.007047f
C996 B.n956 VSUBS 0.007047f
C997 B.n957 VSUBS 0.007047f
C998 B.n958 VSUBS 0.007047f
C999 B.n959 VSUBS 0.007047f
C1000 B.n960 VSUBS 0.007047f
C1001 B.n961 VSUBS 0.007047f
C1002 B.n962 VSUBS 0.007047f
C1003 B.n963 VSUBS 0.007047f
C1004 B.n964 VSUBS 0.007047f
C1005 B.n965 VSUBS 0.007047f
C1006 B.n966 VSUBS 0.007047f
C1007 B.n967 VSUBS 0.007047f
C1008 B.n968 VSUBS 0.007047f
C1009 B.n969 VSUBS 0.007047f
C1010 B.n970 VSUBS 0.007047f
C1011 B.n971 VSUBS 0.007047f
C1012 B.n972 VSUBS 0.007047f
C1013 B.n973 VSUBS 0.007047f
C1014 B.n974 VSUBS 0.007047f
C1015 B.n975 VSUBS 0.007047f
C1016 B.n976 VSUBS 0.007047f
C1017 B.n977 VSUBS 0.007047f
C1018 B.n978 VSUBS 0.007047f
C1019 B.n979 VSUBS 0.007047f
C1020 B.n980 VSUBS 0.007047f
C1021 B.n981 VSUBS 0.007047f
C1022 B.n982 VSUBS 0.007047f
C1023 B.n983 VSUBS 0.007047f
C1024 B.n984 VSUBS 0.007047f
C1025 B.n985 VSUBS 0.007047f
C1026 B.n986 VSUBS 0.007047f
C1027 B.n987 VSUBS 0.007047f
C1028 B.n988 VSUBS 0.007047f
C1029 B.n989 VSUBS 0.007047f
C1030 B.n990 VSUBS 0.007047f
C1031 B.n991 VSUBS 0.007047f
C1032 B.n992 VSUBS 0.007047f
C1033 B.n993 VSUBS 0.007047f
C1034 B.n994 VSUBS 0.007047f
C1035 B.n995 VSUBS 0.007047f
C1036 B.n996 VSUBS 0.007047f
C1037 B.n997 VSUBS 0.007047f
C1038 B.n998 VSUBS 0.007047f
C1039 B.n999 VSUBS 0.015958f
C1040 VDD1.n0 VSUBS 0.028416f
C1041 VDD1.n1 VSUBS 0.027188f
C1042 VDD1.n2 VSUBS 0.014609f
C1043 VDD1.n3 VSUBS 0.034531f
C1044 VDD1.n4 VSUBS 0.015469f
C1045 VDD1.n5 VSUBS 0.027188f
C1046 VDD1.n6 VSUBS 0.014609f
C1047 VDD1.n7 VSUBS 0.034531f
C1048 VDD1.n8 VSUBS 0.015469f
C1049 VDD1.n9 VSUBS 0.027188f
C1050 VDD1.n10 VSUBS 0.014609f
C1051 VDD1.n11 VSUBS 0.034531f
C1052 VDD1.n12 VSUBS 0.015469f
C1053 VDD1.n13 VSUBS 0.027188f
C1054 VDD1.n14 VSUBS 0.014609f
C1055 VDD1.n15 VSUBS 0.034531f
C1056 VDD1.n16 VSUBS 0.015469f
C1057 VDD1.n17 VSUBS 0.027188f
C1058 VDD1.n18 VSUBS 0.014609f
C1059 VDD1.n19 VSUBS 0.034531f
C1060 VDD1.n20 VSUBS 0.015469f
C1061 VDD1.n21 VSUBS 0.027188f
C1062 VDD1.n22 VSUBS 0.014609f
C1063 VDD1.n23 VSUBS 0.034531f
C1064 VDD1.n24 VSUBS 0.015469f
C1065 VDD1.n25 VSUBS 0.027188f
C1066 VDD1.n26 VSUBS 0.014609f
C1067 VDD1.n27 VSUBS 0.034531f
C1068 VDD1.n28 VSUBS 0.034531f
C1069 VDD1.n29 VSUBS 0.015469f
C1070 VDD1.n30 VSUBS 0.027188f
C1071 VDD1.n31 VSUBS 0.014609f
C1072 VDD1.n32 VSUBS 0.034531f
C1073 VDD1.n33 VSUBS 0.015469f
C1074 VDD1.n34 VSUBS 0.30521f
C1075 VDD1.t5 VSUBS 0.075092f
C1076 VDD1.n35 VSUBS 0.025899f
C1077 VDD1.n36 VSUBS 0.025976f
C1078 VDD1.n37 VSUBS 0.014609f
C1079 VDD1.n38 VSUBS 2.21854f
C1080 VDD1.n39 VSUBS 0.027188f
C1081 VDD1.n40 VSUBS 0.014609f
C1082 VDD1.n41 VSUBS 0.015469f
C1083 VDD1.n42 VSUBS 0.034531f
C1084 VDD1.n43 VSUBS 0.034531f
C1085 VDD1.n44 VSUBS 0.015469f
C1086 VDD1.n45 VSUBS 0.014609f
C1087 VDD1.n46 VSUBS 0.027188f
C1088 VDD1.n47 VSUBS 0.027188f
C1089 VDD1.n48 VSUBS 0.014609f
C1090 VDD1.n49 VSUBS 0.015469f
C1091 VDD1.n50 VSUBS 0.034531f
C1092 VDD1.n51 VSUBS 0.034531f
C1093 VDD1.n52 VSUBS 0.015469f
C1094 VDD1.n53 VSUBS 0.014609f
C1095 VDD1.n54 VSUBS 0.027188f
C1096 VDD1.n55 VSUBS 0.027188f
C1097 VDD1.n56 VSUBS 0.014609f
C1098 VDD1.n57 VSUBS 0.015039f
C1099 VDD1.n58 VSUBS 0.015039f
C1100 VDD1.n59 VSUBS 0.034531f
C1101 VDD1.n60 VSUBS 0.034531f
C1102 VDD1.n61 VSUBS 0.015469f
C1103 VDD1.n62 VSUBS 0.014609f
C1104 VDD1.n63 VSUBS 0.027188f
C1105 VDD1.n64 VSUBS 0.027188f
C1106 VDD1.n65 VSUBS 0.014609f
C1107 VDD1.n66 VSUBS 0.015469f
C1108 VDD1.n67 VSUBS 0.034531f
C1109 VDD1.n68 VSUBS 0.034531f
C1110 VDD1.n69 VSUBS 0.015469f
C1111 VDD1.n70 VSUBS 0.014609f
C1112 VDD1.n71 VSUBS 0.027188f
C1113 VDD1.n72 VSUBS 0.027188f
C1114 VDD1.n73 VSUBS 0.014609f
C1115 VDD1.n74 VSUBS 0.015469f
C1116 VDD1.n75 VSUBS 0.034531f
C1117 VDD1.n76 VSUBS 0.034531f
C1118 VDD1.n77 VSUBS 0.015469f
C1119 VDD1.n78 VSUBS 0.014609f
C1120 VDD1.n79 VSUBS 0.027188f
C1121 VDD1.n80 VSUBS 0.027188f
C1122 VDD1.n81 VSUBS 0.014609f
C1123 VDD1.n82 VSUBS 0.015469f
C1124 VDD1.n83 VSUBS 0.034531f
C1125 VDD1.n84 VSUBS 0.034531f
C1126 VDD1.n85 VSUBS 0.015469f
C1127 VDD1.n86 VSUBS 0.014609f
C1128 VDD1.n87 VSUBS 0.027188f
C1129 VDD1.n88 VSUBS 0.027188f
C1130 VDD1.n89 VSUBS 0.014609f
C1131 VDD1.n90 VSUBS 0.015469f
C1132 VDD1.n91 VSUBS 0.034531f
C1133 VDD1.n92 VSUBS 0.034531f
C1134 VDD1.n93 VSUBS 0.015469f
C1135 VDD1.n94 VSUBS 0.014609f
C1136 VDD1.n95 VSUBS 0.027188f
C1137 VDD1.n96 VSUBS 0.027188f
C1138 VDD1.n97 VSUBS 0.014609f
C1139 VDD1.n98 VSUBS 0.015469f
C1140 VDD1.n99 VSUBS 0.034531f
C1141 VDD1.n100 VSUBS 0.084183f
C1142 VDD1.n101 VSUBS 0.015469f
C1143 VDD1.n102 VSUBS 0.02869f
C1144 VDD1.n103 VSUBS 0.066186f
C1145 VDD1.n104 VSUBS 0.096392f
C1146 VDD1.n105 VSUBS 0.028416f
C1147 VDD1.n106 VSUBS 0.027188f
C1148 VDD1.n107 VSUBS 0.014609f
C1149 VDD1.n108 VSUBS 0.034531f
C1150 VDD1.n109 VSUBS 0.015469f
C1151 VDD1.n110 VSUBS 0.027188f
C1152 VDD1.n111 VSUBS 0.014609f
C1153 VDD1.n112 VSUBS 0.034531f
C1154 VDD1.n113 VSUBS 0.015469f
C1155 VDD1.n114 VSUBS 0.027188f
C1156 VDD1.n115 VSUBS 0.014609f
C1157 VDD1.n116 VSUBS 0.034531f
C1158 VDD1.n117 VSUBS 0.015469f
C1159 VDD1.n118 VSUBS 0.027188f
C1160 VDD1.n119 VSUBS 0.014609f
C1161 VDD1.n120 VSUBS 0.034531f
C1162 VDD1.n121 VSUBS 0.015469f
C1163 VDD1.n122 VSUBS 0.027188f
C1164 VDD1.n123 VSUBS 0.014609f
C1165 VDD1.n124 VSUBS 0.034531f
C1166 VDD1.n125 VSUBS 0.015469f
C1167 VDD1.n126 VSUBS 0.027188f
C1168 VDD1.n127 VSUBS 0.014609f
C1169 VDD1.n128 VSUBS 0.034531f
C1170 VDD1.n129 VSUBS 0.015469f
C1171 VDD1.n130 VSUBS 0.027188f
C1172 VDD1.n131 VSUBS 0.014609f
C1173 VDD1.n132 VSUBS 0.034531f
C1174 VDD1.n133 VSUBS 0.015469f
C1175 VDD1.n134 VSUBS 0.027188f
C1176 VDD1.n135 VSUBS 0.014609f
C1177 VDD1.n136 VSUBS 0.034531f
C1178 VDD1.n137 VSUBS 0.015469f
C1179 VDD1.n138 VSUBS 0.30521f
C1180 VDD1.t2 VSUBS 0.075092f
C1181 VDD1.n139 VSUBS 0.025899f
C1182 VDD1.n140 VSUBS 0.025976f
C1183 VDD1.n141 VSUBS 0.014609f
C1184 VDD1.n142 VSUBS 2.21854f
C1185 VDD1.n143 VSUBS 0.027188f
C1186 VDD1.n144 VSUBS 0.014609f
C1187 VDD1.n145 VSUBS 0.015469f
C1188 VDD1.n146 VSUBS 0.034531f
C1189 VDD1.n147 VSUBS 0.034531f
C1190 VDD1.n148 VSUBS 0.015469f
C1191 VDD1.n149 VSUBS 0.014609f
C1192 VDD1.n150 VSUBS 0.027188f
C1193 VDD1.n151 VSUBS 0.027188f
C1194 VDD1.n152 VSUBS 0.014609f
C1195 VDD1.n153 VSUBS 0.015469f
C1196 VDD1.n154 VSUBS 0.034531f
C1197 VDD1.n155 VSUBS 0.034531f
C1198 VDD1.n156 VSUBS 0.034531f
C1199 VDD1.n157 VSUBS 0.015469f
C1200 VDD1.n158 VSUBS 0.014609f
C1201 VDD1.n159 VSUBS 0.027188f
C1202 VDD1.n160 VSUBS 0.027188f
C1203 VDD1.n161 VSUBS 0.014609f
C1204 VDD1.n162 VSUBS 0.015039f
C1205 VDD1.n163 VSUBS 0.015039f
C1206 VDD1.n164 VSUBS 0.034531f
C1207 VDD1.n165 VSUBS 0.034531f
C1208 VDD1.n166 VSUBS 0.015469f
C1209 VDD1.n167 VSUBS 0.014609f
C1210 VDD1.n168 VSUBS 0.027188f
C1211 VDD1.n169 VSUBS 0.027188f
C1212 VDD1.n170 VSUBS 0.014609f
C1213 VDD1.n171 VSUBS 0.015469f
C1214 VDD1.n172 VSUBS 0.034531f
C1215 VDD1.n173 VSUBS 0.034531f
C1216 VDD1.n174 VSUBS 0.015469f
C1217 VDD1.n175 VSUBS 0.014609f
C1218 VDD1.n176 VSUBS 0.027188f
C1219 VDD1.n177 VSUBS 0.027188f
C1220 VDD1.n178 VSUBS 0.014609f
C1221 VDD1.n179 VSUBS 0.015469f
C1222 VDD1.n180 VSUBS 0.034531f
C1223 VDD1.n181 VSUBS 0.034531f
C1224 VDD1.n182 VSUBS 0.015469f
C1225 VDD1.n183 VSUBS 0.014609f
C1226 VDD1.n184 VSUBS 0.027188f
C1227 VDD1.n185 VSUBS 0.027188f
C1228 VDD1.n186 VSUBS 0.014609f
C1229 VDD1.n187 VSUBS 0.015469f
C1230 VDD1.n188 VSUBS 0.034531f
C1231 VDD1.n189 VSUBS 0.034531f
C1232 VDD1.n190 VSUBS 0.015469f
C1233 VDD1.n191 VSUBS 0.014609f
C1234 VDD1.n192 VSUBS 0.027188f
C1235 VDD1.n193 VSUBS 0.027188f
C1236 VDD1.n194 VSUBS 0.014609f
C1237 VDD1.n195 VSUBS 0.015469f
C1238 VDD1.n196 VSUBS 0.034531f
C1239 VDD1.n197 VSUBS 0.034531f
C1240 VDD1.n198 VSUBS 0.015469f
C1241 VDD1.n199 VSUBS 0.014609f
C1242 VDD1.n200 VSUBS 0.027188f
C1243 VDD1.n201 VSUBS 0.027188f
C1244 VDD1.n202 VSUBS 0.014609f
C1245 VDD1.n203 VSUBS 0.015469f
C1246 VDD1.n204 VSUBS 0.034531f
C1247 VDD1.n205 VSUBS 0.084183f
C1248 VDD1.n206 VSUBS 0.015469f
C1249 VDD1.n207 VSUBS 0.02869f
C1250 VDD1.n208 VSUBS 0.066186f
C1251 VDD1.n209 VSUBS 0.095356f
C1252 VDD1.t1 VSUBS 0.417014f
C1253 VDD1.t4 VSUBS 0.417014f
C1254 VDD1.n210 VSUBS 3.52232f
C1255 VDD1.n211 VSUBS 4.37949f
C1256 VDD1.t3 VSUBS 0.417014f
C1257 VDD1.t0 VSUBS 0.417014f
C1258 VDD1.n212 VSUBS 3.51201f
C1259 VDD1.n213 VSUBS 4.25886f
C1260 VP.t1 VSUBS 4.62752f
C1261 VP.n0 VSUBS 1.68761f
C1262 VP.n1 VSUBS 0.02378f
C1263 VP.n2 VSUBS 0.03571f
C1264 VP.n3 VSUBS 0.02378f
C1265 VP.n4 VSUBS 0.033379f
C1266 VP.n5 VSUBS 0.02378f
C1267 VP.n6 VSUBS 0.033722f
C1268 VP.n7 VSUBS 0.02378f
C1269 VP.n8 VSUBS 0.032066f
C1270 VP.t5 VSUBS 4.62752f
C1271 VP.n9 VSUBS 1.68761f
C1272 VP.n10 VSUBS 0.02378f
C1273 VP.n11 VSUBS 0.03571f
C1274 VP.n12 VSUBS 0.02378f
C1275 VP.n13 VSUBS 0.033379f
C1276 VP.t0 VSUBS 4.9945f
C1277 VP.t2 VSUBS 4.62752f
C1278 VP.n14 VSUBS 1.67438f
C1279 VP.n15 VSUBS 1.5986f
C1280 VP.n16 VSUBS 0.297447f
C1281 VP.n17 VSUBS 0.02378f
C1282 VP.n18 VSUBS 0.044319f
C1283 VP.n19 VSUBS 0.044319f
C1284 VP.n20 VSUBS 0.033722f
C1285 VP.n21 VSUBS 0.02378f
C1286 VP.n22 VSUBS 0.02378f
C1287 VP.n23 VSUBS 0.02378f
C1288 VP.n24 VSUBS 0.044319f
C1289 VP.n25 VSUBS 0.044319f
C1290 VP.n26 VSUBS 0.032066f
C1291 VP.n27 VSUBS 0.03838f
C1292 VP.n28 VSUBS 1.69191f
C1293 VP.t3 VSUBS 4.62752f
C1294 VP.n29 VSUBS 1.68761f
C1295 VP.n30 VSUBS 1.70652f
C1296 VP.n31 VSUBS 0.03838f
C1297 VP.n32 VSUBS 0.02378f
C1298 VP.n33 VSUBS 0.044319f
C1299 VP.n34 VSUBS 0.044319f
C1300 VP.n35 VSUBS 0.03571f
C1301 VP.n36 VSUBS 0.02378f
C1302 VP.n37 VSUBS 0.02378f
C1303 VP.n38 VSUBS 0.02378f
C1304 VP.n39 VSUBS 0.044319f
C1305 VP.n40 VSUBS 0.044319f
C1306 VP.t4 VSUBS 4.62752f
C1307 VP.n41 VSUBS 1.59134f
C1308 VP.n42 VSUBS 0.033379f
C1309 VP.n43 VSUBS 0.02378f
C1310 VP.n44 VSUBS 0.02378f
C1311 VP.n45 VSUBS 0.02378f
C1312 VP.n46 VSUBS 0.044319f
C1313 VP.n47 VSUBS 0.044319f
C1314 VP.n48 VSUBS 0.033722f
C1315 VP.n49 VSUBS 0.02378f
C1316 VP.n50 VSUBS 0.02378f
C1317 VP.n51 VSUBS 0.02378f
C1318 VP.n52 VSUBS 0.044319f
C1319 VP.n53 VSUBS 0.044319f
C1320 VP.n54 VSUBS 0.032066f
C1321 VP.n55 VSUBS 0.03838f
C1322 VP.n56 VSUBS 0.064754f
C1323 VTAIL.t7 VSUBS 0.427487f
C1324 VTAIL.t6 VSUBS 0.427487f
C1325 VTAIL.n0 VSUBS 3.43219f
C1326 VTAIL.n1 VSUBS 0.946383f
C1327 VTAIL.n2 VSUBS 0.02913f
C1328 VTAIL.n3 VSUBS 0.027871f
C1329 VTAIL.n4 VSUBS 0.014976f
C1330 VTAIL.n5 VSUBS 0.035399f
C1331 VTAIL.n6 VSUBS 0.015857f
C1332 VTAIL.n7 VSUBS 0.027871f
C1333 VTAIL.n8 VSUBS 0.014976f
C1334 VTAIL.n9 VSUBS 0.035399f
C1335 VTAIL.n10 VSUBS 0.015857f
C1336 VTAIL.n11 VSUBS 0.027871f
C1337 VTAIL.n12 VSUBS 0.014976f
C1338 VTAIL.n13 VSUBS 0.035399f
C1339 VTAIL.n14 VSUBS 0.015857f
C1340 VTAIL.n15 VSUBS 0.027871f
C1341 VTAIL.n16 VSUBS 0.014976f
C1342 VTAIL.n17 VSUBS 0.035399f
C1343 VTAIL.n18 VSUBS 0.015857f
C1344 VTAIL.n19 VSUBS 0.027871f
C1345 VTAIL.n20 VSUBS 0.014976f
C1346 VTAIL.n21 VSUBS 0.035399f
C1347 VTAIL.n22 VSUBS 0.015857f
C1348 VTAIL.n23 VSUBS 0.027871f
C1349 VTAIL.n24 VSUBS 0.014976f
C1350 VTAIL.n25 VSUBS 0.035399f
C1351 VTAIL.n26 VSUBS 0.015857f
C1352 VTAIL.n27 VSUBS 0.027871f
C1353 VTAIL.n28 VSUBS 0.014976f
C1354 VTAIL.n29 VSUBS 0.035399f
C1355 VTAIL.n30 VSUBS 0.015857f
C1356 VTAIL.n31 VSUBS 0.027871f
C1357 VTAIL.n32 VSUBS 0.014976f
C1358 VTAIL.n33 VSUBS 0.035399f
C1359 VTAIL.n34 VSUBS 0.015857f
C1360 VTAIL.n35 VSUBS 0.312876f
C1361 VTAIL.t1 VSUBS 0.076978f
C1362 VTAIL.n36 VSUBS 0.026549f
C1363 VTAIL.n37 VSUBS 0.026629f
C1364 VTAIL.n38 VSUBS 0.014976f
C1365 VTAIL.n39 VSUBS 2.27426f
C1366 VTAIL.n40 VSUBS 0.027871f
C1367 VTAIL.n41 VSUBS 0.014976f
C1368 VTAIL.n42 VSUBS 0.015857f
C1369 VTAIL.n43 VSUBS 0.035399f
C1370 VTAIL.n44 VSUBS 0.035399f
C1371 VTAIL.n45 VSUBS 0.015857f
C1372 VTAIL.n46 VSUBS 0.014976f
C1373 VTAIL.n47 VSUBS 0.027871f
C1374 VTAIL.n48 VSUBS 0.027871f
C1375 VTAIL.n49 VSUBS 0.014976f
C1376 VTAIL.n50 VSUBS 0.015857f
C1377 VTAIL.n51 VSUBS 0.035399f
C1378 VTAIL.n52 VSUBS 0.035399f
C1379 VTAIL.n53 VSUBS 0.035399f
C1380 VTAIL.n54 VSUBS 0.015857f
C1381 VTAIL.n55 VSUBS 0.014976f
C1382 VTAIL.n56 VSUBS 0.027871f
C1383 VTAIL.n57 VSUBS 0.027871f
C1384 VTAIL.n58 VSUBS 0.014976f
C1385 VTAIL.n59 VSUBS 0.015417f
C1386 VTAIL.n60 VSUBS 0.015417f
C1387 VTAIL.n61 VSUBS 0.035399f
C1388 VTAIL.n62 VSUBS 0.035399f
C1389 VTAIL.n63 VSUBS 0.015857f
C1390 VTAIL.n64 VSUBS 0.014976f
C1391 VTAIL.n65 VSUBS 0.027871f
C1392 VTAIL.n66 VSUBS 0.027871f
C1393 VTAIL.n67 VSUBS 0.014976f
C1394 VTAIL.n68 VSUBS 0.015857f
C1395 VTAIL.n69 VSUBS 0.035399f
C1396 VTAIL.n70 VSUBS 0.035399f
C1397 VTAIL.n71 VSUBS 0.015857f
C1398 VTAIL.n72 VSUBS 0.014976f
C1399 VTAIL.n73 VSUBS 0.027871f
C1400 VTAIL.n74 VSUBS 0.027871f
C1401 VTAIL.n75 VSUBS 0.014976f
C1402 VTAIL.n76 VSUBS 0.015857f
C1403 VTAIL.n77 VSUBS 0.035399f
C1404 VTAIL.n78 VSUBS 0.035399f
C1405 VTAIL.n79 VSUBS 0.015857f
C1406 VTAIL.n80 VSUBS 0.014976f
C1407 VTAIL.n81 VSUBS 0.027871f
C1408 VTAIL.n82 VSUBS 0.027871f
C1409 VTAIL.n83 VSUBS 0.014976f
C1410 VTAIL.n84 VSUBS 0.015857f
C1411 VTAIL.n85 VSUBS 0.035399f
C1412 VTAIL.n86 VSUBS 0.035399f
C1413 VTAIL.n87 VSUBS 0.015857f
C1414 VTAIL.n88 VSUBS 0.014976f
C1415 VTAIL.n89 VSUBS 0.027871f
C1416 VTAIL.n90 VSUBS 0.027871f
C1417 VTAIL.n91 VSUBS 0.014976f
C1418 VTAIL.n92 VSUBS 0.015857f
C1419 VTAIL.n93 VSUBS 0.035399f
C1420 VTAIL.n94 VSUBS 0.035399f
C1421 VTAIL.n95 VSUBS 0.015857f
C1422 VTAIL.n96 VSUBS 0.014976f
C1423 VTAIL.n97 VSUBS 0.027871f
C1424 VTAIL.n98 VSUBS 0.027871f
C1425 VTAIL.n99 VSUBS 0.014976f
C1426 VTAIL.n100 VSUBS 0.015857f
C1427 VTAIL.n101 VSUBS 0.035399f
C1428 VTAIL.n102 VSUBS 0.086297f
C1429 VTAIL.n103 VSUBS 0.015857f
C1430 VTAIL.n104 VSUBS 0.02941f
C1431 VTAIL.n105 VSUBS 0.067848f
C1432 VTAIL.n106 VSUBS 0.065227f
C1433 VTAIL.n107 VSUBS 0.528957f
C1434 VTAIL.t10 VSUBS 0.427487f
C1435 VTAIL.t9 VSUBS 0.427487f
C1436 VTAIL.n108 VSUBS 3.43219f
C1437 VTAIL.n109 VSUBS 3.47177f
C1438 VTAIL.t3 VSUBS 0.427487f
C1439 VTAIL.t8 VSUBS 0.427487f
C1440 VTAIL.n110 VSUBS 3.43221f
C1441 VTAIL.n111 VSUBS 3.47175f
C1442 VTAIL.n112 VSUBS 0.02913f
C1443 VTAIL.n113 VSUBS 0.027871f
C1444 VTAIL.n114 VSUBS 0.014976f
C1445 VTAIL.n115 VSUBS 0.035399f
C1446 VTAIL.n116 VSUBS 0.015857f
C1447 VTAIL.n117 VSUBS 0.027871f
C1448 VTAIL.n118 VSUBS 0.014976f
C1449 VTAIL.n119 VSUBS 0.035399f
C1450 VTAIL.n120 VSUBS 0.015857f
C1451 VTAIL.n121 VSUBS 0.027871f
C1452 VTAIL.n122 VSUBS 0.014976f
C1453 VTAIL.n123 VSUBS 0.035399f
C1454 VTAIL.n124 VSUBS 0.015857f
C1455 VTAIL.n125 VSUBS 0.027871f
C1456 VTAIL.n126 VSUBS 0.014976f
C1457 VTAIL.n127 VSUBS 0.035399f
C1458 VTAIL.n128 VSUBS 0.015857f
C1459 VTAIL.n129 VSUBS 0.027871f
C1460 VTAIL.n130 VSUBS 0.014976f
C1461 VTAIL.n131 VSUBS 0.035399f
C1462 VTAIL.n132 VSUBS 0.015857f
C1463 VTAIL.n133 VSUBS 0.027871f
C1464 VTAIL.n134 VSUBS 0.014976f
C1465 VTAIL.n135 VSUBS 0.035399f
C1466 VTAIL.n136 VSUBS 0.015857f
C1467 VTAIL.n137 VSUBS 0.027871f
C1468 VTAIL.n138 VSUBS 0.014976f
C1469 VTAIL.n139 VSUBS 0.035399f
C1470 VTAIL.n140 VSUBS 0.035399f
C1471 VTAIL.n141 VSUBS 0.015857f
C1472 VTAIL.n142 VSUBS 0.027871f
C1473 VTAIL.n143 VSUBS 0.014976f
C1474 VTAIL.n144 VSUBS 0.035399f
C1475 VTAIL.n145 VSUBS 0.015857f
C1476 VTAIL.n146 VSUBS 0.312876f
C1477 VTAIL.t5 VSUBS 0.076978f
C1478 VTAIL.n147 VSUBS 0.026549f
C1479 VTAIL.n148 VSUBS 0.026629f
C1480 VTAIL.n149 VSUBS 0.014976f
C1481 VTAIL.n150 VSUBS 2.27426f
C1482 VTAIL.n151 VSUBS 0.027871f
C1483 VTAIL.n152 VSUBS 0.014976f
C1484 VTAIL.n153 VSUBS 0.015857f
C1485 VTAIL.n154 VSUBS 0.035399f
C1486 VTAIL.n155 VSUBS 0.035399f
C1487 VTAIL.n156 VSUBS 0.015857f
C1488 VTAIL.n157 VSUBS 0.014976f
C1489 VTAIL.n158 VSUBS 0.027871f
C1490 VTAIL.n159 VSUBS 0.027871f
C1491 VTAIL.n160 VSUBS 0.014976f
C1492 VTAIL.n161 VSUBS 0.015857f
C1493 VTAIL.n162 VSUBS 0.035399f
C1494 VTAIL.n163 VSUBS 0.035399f
C1495 VTAIL.n164 VSUBS 0.015857f
C1496 VTAIL.n165 VSUBS 0.014976f
C1497 VTAIL.n166 VSUBS 0.027871f
C1498 VTAIL.n167 VSUBS 0.027871f
C1499 VTAIL.n168 VSUBS 0.014976f
C1500 VTAIL.n169 VSUBS 0.015417f
C1501 VTAIL.n170 VSUBS 0.015417f
C1502 VTAIL.n171 VSUBS 0.035399f
C1503 VTAIL.n172 VSUBS 0.035399f
C1504 VTAIL.n173 VSUBS 0.015857f
C1505 VTAIL.n174 VSUBS 0.014976f
C1506 VTAIL.n175 VSUBS 0.027871f
C1507 VTAIL.n176 VSUBS 0.027871f
C1508 VTAIL.n177 VSUBS 0.014976f
C1509 VTAIL.n178 VSUBS 0.015857f
C1510 VTAIL.n179 VSUBS 0.035399f
C1511 VTAIL.n180 VSUBS 0.035399f
C1512 VTAIL.n181 VSUBS 0.015857f
C1513 VTAIL.n182 VSUBS 0.014976f
C1514 VTAIL.n183 VSUBS 0.027871f
C1515 VTAIL.n184 VSUBS 0.027871f
C1516 VTAIL.n185 VSUBS 0.014976f
C1517 VTAIL.n186 VSUBS 0.015857f
C1518 VTAIL.n187 VSUBS 0.035399f
C1519 VTAIL.n188 VSUBS 0.035399f
C1520 VTAIL.n189 VSUBS 0.015857f
C1521 VTAIL.n190 VSUBS 0.014976f
C1522 VTAIL.n191 VSUBS 0.027871f
C1523 VTAIL.n192 VSUBS 0.027871f
C1524 VTAIL.n193 VSUBS 0.014976f
C1525 VTAIL.n194 VSUBS 0.015857f
C1526 VTAIL.n195 VSUBS 0.035399f
C1527 VTAIL.n196 VSUBS 0.035399f
C1528 VTAIL.n197 VSUBS 0.015857f
C1529 VTAIL.n198 VSUBS 0.014976f
C1530 VTAIL.n199 VSUBS 0.027871f
C1531 VTAIL.n200 VSUBS 0.027871f
C1532 VTAIL.n201 VSUBS 0.014976f
C1533 VTAIL.n202 VSUBS 0.015857f
C1534 VTAIL.n203 VSUBS 0.035399f
C1535 VTAIL.n204 VSUBS 0.035399f
C1536 VTAIL.n205 VSUBS 0.015857f
C1537 VTAIL.n206 VSUBS 0.014976f
C1538 VTAIL.n207 VSUBS 0.027871f
C1539 VTAIL.n208 VSUBS 0.027871f
C1540 VTAIL.n209 VSUBS 0.014976f
C1541 VTAIL.n210 VSUBS 0.015857f
C1542 VTAIL.n211 VSUBS 0.035399f
C1543 VTAIL.n212 VSUBS 0.086297f
C1544 VTAIL.n213 VSUBS 0.015857f
C1545 VTAIL.n214 VSUBS 0.02941f
C1546 VTAIL.n215 VSUBS 0.067848f
C1547 VTAIL.n216 VSUBS 0.065227f
C1548 VTAIL.n217 VSUBS 0.528957f
C1549 VTAIL.t2 VSUBS 0.427487f
C1550 VTAIL.t11 VSUBS 0.427487f
C1551 VTAIL.n218 VSUBS 3.43221f
C1552 VTAIL.n219 VSUBS 1.17165f
C1553 VTAIL.n220 VSUBS 0.02913f
C1554 VTAIL.n221 VSUBS 0.027871f
C1555 VTAIL.n222 VSUBS 0.014976f
C1556 VTAIL.n223 VSUBS 0.035399f
C1557 VTAIL.n224 VSUBS 0.015857f
C1558 VTAIL.n225 VSUBS 0.027871f
C1559 VTAIL.n226 VSUBS 0.014976f
C1560 VTAIL.n227 VSUBS 0.035399f
C1561 VTAIL.n228 VSUBS 0.015857f
C1562 VTAIL.n229 VSUBS 0.027871f
C1563 VTAIL.n230 VSUBS 0.014976f
C1564 VTAIL.n231 VSUBS 0.035399f
C1565 VTAIL.n232 VSUBS 0.015857f
C1566 VTAIL.n233 VSUBS 0.027871f
C1567 VTAIL.n234 VSUBS 0.014976f
C1568 VTAIL.n235 VSUBS 0.035399f
C1569 VTAIL.n236 VSUBS 0.015857f
C1570 VTAIL.n237 VSUBS 0.027871f
C1571 VTAIL.n238 VSUBS 0.014976f
C1572 VTAIL.n239 VSUBS 0.035399f
C1573 VTAIL.n240 VSUBS 0.015857f
C1574 VTAIL.n241 VSUBS 0.027871f
C1575 VTAIL.n242 VSUBS 0.014976f
C1576 VTAIL.n243 VSUBS 0.035399f
C1577 VTAIL.n244 VSUBS 0.015857f
C1578 VTAIL.n245 VSUBS 0.027871f
C1579 VTAIL.n246 VSUBS 0.014976f
C1580 VTAIL.n247 VSUBS 0.035399f
C1581 VTAIL.n248 VSUBS 0.035399f
C1582 VTAIL.n249 VSUBS 0.015857f
C1583 VTAIL.n250 VSUBS 0.027871f
C1584 VTAIL.n251 VSUBS 0.014976f
C1585 VTAIL.n252 VSUBS 0.035399f
C1586 VTAIL.n253 VSUBS 0.015857f
C1587 VTAIL.n254 VSUBS 0.312876f
C1588 VTAIL.t0 VSUBS 0.076978f
C1589 VTAIL.n255 VSUBS 0.026549f
C1590 VTAIL.n256 VSUBS 0.026629f
C1591 VTAIL.n257 VSUBS 0.014976f
C1592 VTAIL.n258 VSUBS 2.27426f
C1593 VTAIL.n259 VSUBS 0.027871f
C1594 VTAIL.n260 VSUBS 0.014976f
C1595 VTAIL.n261 VSUBS 0.015857f
C1596 VTAIL.n262 VSUBS 0.035399f
C1597 VTAIL.n263 VSUBS 0.035399f
C1598 VTAIL.n264 VSUBS 0.015857f
C1599 VTAIL.n265 VSUBS 0.014976f
C1600 VTAIL.n266 VSUBS 0.027871f
C1601 VTAIL.n267 VSUBS 0.027871f
C1602 VTAIL.n268 VSUBS 0.014976f
C1603 VTAIL.n269 VSUBS 0.015857f
C1604 VTAIL.n270 VSUBS 0.035399f
C1605 VTAIL.n271 VSUBS 0.035399f
C1606 VTAIL.n272 VSUBS 0.015857f
C1607 VTAIL.n273 VSUBS 0.014976f
C1608 VTAIL.n274 VSUBS 0.027871f
C1609 VTAIL.n275 VSUBS 0.027871f
C1610 VTAIL.n276 VSUBS 0.014976f
C1611 VTAIL.n277 VSUBS 0.015417f
C1612 VTAIL.n278 VSUBS 0.015417f
C1613 VTAIL.n279 VSUBS 0.035399f
C1614 VTAIL.n280 VSUBS 0.035399f
C1615 VTAIL.n281 VSUBS 0.015857f
C1616 VTAIL.n282 VSUBS 0.014976f
C1617 VTAIL.n283 VSUBS 0.027871f
C1618 VTAIL.n284 VSUBS 0.027871f
C1619 VTAIL.n285 VSUBS 0.014976f
C1620 VTAIL.n286 VSUBS 0.015857f
C1621 VTAIL.n287 VSUBS 0.035399f
C1622 VTAIL.n288 VSUBS 0.035399f
C1623 VTAIL.n289 VSUBS 0.015857f
C1624 VTAIL.n290 VSUBS 0.014976f
C1625 VTAIL.n291 VSUBS 0.027871f
C1626 VTAIL.n292 VSUBS 0.027871f
C1627 VTAIL.n293 VSUBS 0.014976f
C1628 VTAIL.n294 VSUBS 0.015857f
C1629 VTAIL.n295 VSUBS 0.035399f
C1630 VTAIL.n296 VSUBS 0.035399f
C1631 VTAIL.n297 VSUBS 0.015857f
C1632 VTAIL.n298 VSUBS 0.014976f
C1633 VTAIL.n299 VSUBS 0.027871f
C1634 VTAIL.n300 VSUBS 0.027871f
C1635 VTAIL.n301 VSUBS 0.014976f
C1636 VTAIL.n302 VSUBS 0.015857f
C1637 VTAIL.n303 VSUBS 0.035399f
C1638 VTAIL.n304 VSUBS 0.035399f
C1639 VTAIL.n305 VSUBS 0.015857f
C1640 VTAIL.n306 VSUBS 0.014976f
C1641 VTAIL.n307 VSUBS 0.027871f
C1642 VTAIL.n308 VSUBS 0.027871f
C1643 VTAIL.n309 VSUBS 0.014976f
C1644 VTAIL.n310 VSUBS 0.015857f
C1645 VTAIL.n311 VSUBS 0.035399f
C1646 VTAIL.n312 VSUBS 0.035399f
C1647 VTAIL.n313 VSUBS 0.015857f
C1648 VTAIL.n314 VSUBS 0.014976f
C1649 VTAIL.n315 VSUBS 0.027871f
C1650 VTAIL.n316 VSUBS 0.027871f
C1651 VTAIL.n317 VSUBS 0.014976f
C1652 VTAIL.n318 VSUBS 0.015857f
C1653 VTAIL.n319 VSUBS 0.035399f
C1654 VTAIL.n320 VSUBS 0.086297f
C1655 VTAIL.n321 VSUBS 0.015857f
C1656 VTAIL.n322 VSUBS 0.02941f
C1657 VTAIL.n323 VSUBS 0.067848f
C1658 VTAIL.n324 VSUBS 0.065227f
C1659 VTAIL.n325 VSUBS 2.52171f
C1660 VTAIL.n326 VSUBS 0.02913f
C1661 VTAIL.n327 VSUBS 0.027871f
C1662 VTAIL.n328 VSUBS 0.014976f
C1663 VTAIL.n329 VSUBS 0.035399f
C1664 VTAIL.n330 VSUBS 0.015857f
C1665 VTAIL.n331 VSUBS 0.027871f
C1666 VTAIL.n332 VSUBS 0.014976f
C1667 VTAIL.n333 VSUBS 0.035399f
C1668 VTAIL.n334 VSUBS 0.015857f
C1669 VTAIL.n335 VSUBS 0.027871f
C1670 VTAIL.n336 VSUBS 0.014976f
C1671 VTAIL.n337 VSUBS 0.035399f
C1672 VTAIL.n338 VSUBS 0.015857f
C1673 VTAIL.n339 VSUBS 0.027871f
C1674 VTAIL.n340 VSUBS 0.014976f
C1675 VTAIL.n341 VSUBS 0.035399f
C1676 VTAIL.n342 VSUBS 0.015857f
C1677 VTAIL.n343 VSUBS 0.027871f
C1678 VTAIL.n344 VSUBS 0.014976f
C1679 VTAIL.n345 VSUBS 0.035399f
C1680 VTAIL.n346 VSUBS 0.015857f
C1681 VTAIL.n347 VSUBS 0.027871f
C1682 VTAIL.n348 VSUBS 0.014976f
C1683 VTAIL.n349 VSUBS 0.035399f
C1684 VTAIL.n350 VSUBS 0.015857f
C1685 VTAIL.n351 VSUBS 0.027871f
C1686 VTAIL.n352 VSUBS 0.014976f
C1687 VTAIL.n353 VSUBS 0.035399f
C1688 VTAIL.n354 VSUBS 0.015857f
C1689 VTAIL.n355 VSUBS 0.027871f
C1690 VTAIL.n356 VSUBS 0.014976f
C1691 VTAIL.n357 VSUBS 0.035399f
C1692 VTAIL.n358 VSUBS 0.015857f
C1693 VTAIL.n359 VSUBS 0.312876f
C1694 VTAIL.t4 VSUBS 0.076978f
C1695 VTAIL.n360 VSUBS 0.026549f
C1696 VTAIL.n361 VSUBS 0.026629f
C1697 VTAIL.n362 VSUBS 0.014976f
C1698 VTAIL.n363 VSUBS 2.27426f
C1699 VTAIL.n364 VSUBS 0.027871f
C1700 VTAIL.n365 VSUBS 0.014976f
C1701 VTAIL.n366 VSUBS 0.015857f
C1702 VTAIL.n367 VSUBS 0.035399f
C1703 VTAIL.n368 VSUBS 0.035399f
C1704 VTAIL.n369 VSUBS 0.015857f
C1705 VTAIL.n370 VSUBS 0.014976f
C1706 VTAIL.n371 VSUBS 0.027871f
C1707 VTAIL.n372 VSUBS 0.027871f
C1708 VTAIL.n373 VSUBS 0.014976f
C1709 VTAIL.n374 VSUBS 0.015857f
C1710 VTAIL.n375 VSUBS 0.035399f
C1711 VTAIL.n376 VSUBS 0.035399f
C1712 VTAIL.n377 VSUBS 0.035399f
C1713 VTAIL.n378 VSUBS 0.015857f
C1714 VTAIL.n379 VSUBS 0.014976f
C1715 VTAIL.n380 VSUBS 0.027871f
C1716 VTAIL.n381 VSUBS 0.027871f
C1717 VTAIL.n382 VSUBS 0.014976f
C1718 VTAIL.n383 VSUBS 0.015417f
C1719 VTAIL.n384 VSUBS 0.015417f
C1720 VTAIL.n385 VSUBS 0.035399f
C1721 VTAIL.n386 VSUBS 0.035399f
C1722 VTAIL.n387 VSUBS 0.015857f
C1723 VTAIL.n388 VSUBS 0.014976f
C1724 VTAIL.n389 VSUBS 0.027871f
C1725 VTAIL.n390 VSUBS 0.027871f
C1726 VTAIL.n391 VSUBS 0.014976f
C1727 VTAIL.n392 VSUBS 0.015857f
C1728 VTAIL.n393 VSUBS 0.035399f
C1729 VTAIL.n394 VSUBS 0.035399f
C1730 VTAIL.n395 VSUBS 0.015857f
C1731 VTAIL.n396 VSUBS 0.014976f
C1732 VTAIL.n397 VSUBS 0.027871f
C1733 VTAIL.n398 VSUBS 0.027871f
C1734 VTAIL.n399 VSUBS 0.014976f
C1735 VTAIL.n400 VSUBS 0.015857f
C1736 VTAIL.n401 VSUBS 0.035399f
C1737 VTAIL.n402 VSUBS 0.035399f
C1738 VTAIL.n403 VSUBS 0.015857f
C1739 VTAIL.n404 VSUBS 0.014976f
C1740 VTAIL.n405 VSUBS 0.027871f
C1741 VTAIL.n406 VSUBS 0.027871f
C1742 VTAIL.n407 VSUBS 0.014976f
C1743 VTAIL.n408 VSUBS 0.015857f
C1744 VTAIL.n409 VSUBS 0.035399f
C1745 VTAIL.n410 VSUBS 0.035399f
C1746 VTAIL.n411 VSUBS 0.015857f
C1747 VTAIL.n412 VSUBS 0.014976f
C1748 VTAIL.n413 VSUBS 0.027871f
C1749 VTAIL.n414 VSUBS 0.027871f
C1750 VTAIL.n415 VSUBS 0.014976f
C1751 VTAIL.n416 VSUBS 0.015857f
C1752 VTAIL.n417 VSUBS 0.035399f
C1753 VTAIL.n418 VSUBS 0.035399f
C1754 VTAIL.n419 VSUBS 0.015857f
C1755 VTAIL.n420 VSUBS 0.014976f
C1756 VTAIL.n421 VSUBS 0.027871f
C1757 VTAIL.n422 VSUBS 0.027871f
C1758 VTAIL.n423 VSUBS 0.014976f
C1759 VTAIL.n424 VSUBS 0.015857f
C1760 VTAIL.n425 VSUBS 0.035399f
C1761 VTAIL.n426 VSUBS 0.086297f
C1762 VTAIL.n427 VSUBS 0.015857f
C1763 VTAIL.n428 VSUBS 0.02941f
C1764 VTAIL.n429 VSUBS 0.067848f
C1765 VTAIL.n430 VSUBS 0.065227f
C1766 VTAIL.n431 VSUBS 2.43965f
C1767 VDD2.n0 VSUBS 0.028315f
C1768 VDD2.n1 VSUBS 0.027091f
C1769 VDD2.n2 VSUBS 0.014558f
C1770 VDD2.n3 VSUBS 0.034409f
C1771 VDD2.n4 VSUBS 0.015414f
C1772 VDD2.n5 VSUBS 0.027091f
C1773 VDD2.n6 VSUBS 0.014558f
C1774 VDD2.n7 VSUBS 0.034409f
C1775 VDD2.n8 VSUBS 0.015414f
C1776 VDD2.n9 VSUBS 0.027091f
C1777 VDD2.n10 VSUBS 0.014558f
C1778 VDD2.n11 VSUBS 0.034409f
C1779 VDD2.n12 VSUBS 0.015414f
C1780 VDD2.n13 VSUBS 0.027091f
C1781 VDD2.n14 VSUBS 0.014558f
C1782 VDD2.n15 VSUBS 0.034409f
C1783 VDD2.n16 VSUBS 0.015414f
C1784 VDD2.n17 VSUBS 0.027091f
C1785 VDD2.n18 VSUBS 0.014558f
C1786 VDD2.n19 VSUBS 0.034409f
C1787 VDD2.n20 VSUBS 0.015414f
C1788 VDD2.n21 VSUBS 0.027091f
C1789 VDD2.n22 VSUBS 0.014558f
C1790 VDD2.n23 VSUBS 0.034409f
C1791 VDD2.n24 VSUBS 0.015414f
C1792 VDD2.n25 VSUBS 0.027091f
C1793 VDD2.n26 VSUBS 0.014558f
C1794 VDD2.n27 VSUBS 0.034409f
C1795 VDD2.n28 VSUBS 0.015414f
C1796 VDD2.n29 VSUBS 0.027091f
C1797 VDD2.n30 VSUBS 0.014558f
C1798 VDD2.n31 VSUBS 0.034409f
C1799 VDD2.n32 VSUBS 0.015414f
C1800 VDD2.n33 VSUBS 0.304129f
C1801 VDD2.t4 VSUBS 0.074826f
C1802 VDD2.n34 VSUBS 0.025807f
C1803 VDD2.n35 VSUBS 0.025884f
C1804 VDD2.n36 VSUBS 0.014558f
C1805 VDD2.n37 VSUBS 2.21068f
C1806 VDD2.n38 VSUBS 0.027091f
C1807 VDD2.n39 VSUBS 0.014558f
C1808 VDD2.n40 VSUBS 0.015414f
C1809 VDD2.n41 VSUBS 0.034409f
C1810 VDD2.n42 VSUBS 0.034409f
C1811 VDD2.n43 VSUBS 0.015414f
C1812 VDD2.n44 VSUBS 0.014558f
C1813 VDD2.n45 VSUBS 0.027091f
C1814 VDD2.n46 VSUBS 0.027091f
C1815 VDD2.n47 VSUBS 0.014558f
C1816 VDD2.n48 VSUBS 0.015414f
C1817 VDD2.n49 VSUBS 0.034409f
C1818 VDD2.n50 VSUBS 0.034409f
C1819 VDD2.n51 VSUBS 0.034409f
C1820 VDD2.n52 VSUBS 0.015414f
C1821 VDD2.n53 VSUBS 0.014558f
C1822 VDD2.n54 VSUBS 0.027091f
C1823 VDD2.n55 VSUBS 0.027091f
C1824 VDD2.n56 VSUBS 0.014558f
C1825 VDD2.n57 VSUBS 0.014986f
C1826 VDD2.n58 VSUBS 0.014986f
C1827 VDD2.n59 VSUBS 0.034409f
C1828 VDD2.n60 VSUBS 0.034409f
C1829 VDD2.n61 VSUBS 0.015414f
C1830 VDD2.n62 VSUBS 0.014558f
C1831 VDD2.n63 VSUBS 0.027091f
C1832 VDD2.n64 VSUBS 0.027091f
C1833 VDD2.n65 VSUBS 0.014558f
C1834 VDD2.n66 VSUBS 0.015414f
C1835 VDD2.n67 VSUBS 0.034409f
C1836 VDD2.n68 VSUBS 0.034409f
C1837 VDD2.n69 VSUBS 0.015414f
C1838 VDD2.n70 VSUBS 0.014558f
C1839 VDD2.n71 VSUBS 0.027091f
C1840 VDD2.n72 VSUBS 0.027091f
C1841 VDD2.n73 VSUBS 0.014558f
C1842 VDD2.n74 VSUBS 0.015414f
C1843 VDD2.n75 VSUBS 0.034409f
C1844 VDD2.n76 VSUBS 0.034409f
C1845 VDD2.n77 VSUBS 0.015414f
C1846 VDD2.n78 VSUBS 0.014558f
C1847 VDD2.n79 VSUBS 0.027091f
C1848 VDD2.n80 VSUBS 0.027091f
C1849 VDD2.n81 VSUBS 0.014558f
C1850 VDD2.n82 VSUBS 0.015414f
C1851 VDD2.n83 VSUBS 0.034409f
C1852 VDD2.n84 VSUBS 0.034409f
C1853 VDD2.n85 VSUBS 0.015414f
C1854 VDD2.n86 VSUBS 0.014558f
C1855 VDD2.n87 VSUBS 0.027091f
C1856 VDD2.n88 VSUBS 0.027091f
C1857 VDD2.n89 VSUBS 0.014558f
C1858 VDD2.n90 VSUBS 0.015414f
C1859 VDD2.n91 VSUBS 0.034409f
C1860 VDD2.n92 VSUBS 0.034409f
C1861 VDD2.n93 VSUBS 0.015414f
C1862 VDD2.n94 VSUBS 0.014558f
C1863 VDD2.n95 VSUBS 0.027091f
C1864 VDD2.n96 VSUBS 0.027091f
C1865 VDD2.n97 VSUBS 0.014558f
C1866 VDD2.n98 VSUBS 0.015414f
C1867 VDD2.n99 VSUBS 0.034409f
C1868 VDD2.n100 VSUBS 0.083885f
C1869 VDD2.n101 VSUBS 0.015414f
C1870 VDD2.n102 VSUBS 0.028588f
C1871 VDD2.n103 VSUBS 0.065951f
C1872 VDD2.n104 VSUBS 0.095018f
C1873 VDD2.t3 VSUBS 0.415536f
C1874 VDD2.t1 VSUBS 0.415536f
C1875 VDD2.n105 VSUBS 3.50983f
C1876 VDD2.n106 VSUBS 4.1932f
C1877 VDD2.n107 VSUBS 0.028315f
C1878 VDD2.n108 VSUBS 0.027091f
C1879 VDD2.n109 VSUBS 0.014558f
C1880 VDD2.n110 VSUBS 0.034409f
C1881 VDD2.n111 VSUBS 0.015414f
C1882 VDD2.n112 VSUBS 0.027091f
C1883 VDD2.n113 VSUBS 0.014558f
C1884 VDD2.n114 VSUBS 0.034409f
C1885 VDD2.n115 VSUBS 0.015414f
C1886 VDD2.n116 VSUBS 0.027091f
C1887 VDD2.n117 VSUBS 0.014558f
C1888 VDD2.n118 VSUBS 0.034409f
C1889 VDD2.n119 VSUBS 0.015414f
C1890 VDD2.n120 VSUBS 0.027091f
C1891 VDD2.n121 VSUBS 0.014558f
C1892 VDD2.n122 VSUBS 0.034409f
C1893 VDD2.n123 VSUBS 0.015414f
C1894 VDD2.n124 VSUBS 0.027091f
C1895 VDD2.n125 VSUBS 0.014558f
C1896 VDD2.n126 VSUBS 0.034409f
C1897 VDD2.n127 VSUBS 0.015414f
C1898 VDD2.n128 VSUBS 0.027091f
C1899 VDD2.n129 VSUBS 0.014558f
C1900 VDD2.n130 VSUBS 0.034409f
C1901 VDD2.n131 VSUBS 0.015414f
C1902 VDD2.n132 VSUBS 0.027091f
C1903 VDD2.n133 VSUBS 0.014558f
C1904 VDD2.n134 VSUBS 0.034409f
C1905 VDD2.n135 VSUBS 0.034409f
C1906 VDD2.n136 VSUBS 0.015414f
C1907 VDD2.n137 VSUBS 0.027091f
C1908 VDD2.n138 VSUBS 0.014558f
C1909 VDD2.n139 VSUBS 0.034409f
C1910 VDD2.n140 VSUBS 0.015414f
C1911 VDD2.n141 VSUBS 0.304128f
C1912 VDD2.t5 VSUBS 0.074826f
C1913 VDD2.n142 VSUBS 0.025807f
C1914 VDD2.n143 VSUBS 0.025884f
C1915 VDD2.n144 VSUBS 0.014558f
C1916 VDD2.n145 VSUBS 2.21068f
C1917 VDD2.n146 VSUBS 0.027091f
C1918 VDD2.n147 VSUBS 0.014558f
C1919 VDD2.n148 VSUBS 0.015414f
C1920 VDD2.n149 VSUBS 0.034409f
C1921 VDD2.n150 VSUBS 0.034409f
C1922 VDD2.n151 VSUBS 0.015414f
C1923 VDD2.n152 VSUBS 0.014558f
C1924 VDD2.n153 VSUBS 0.027091f
C1925 VDD2.n154 VSUBS 0.027091f
C1926 VDD2.n155 VSUBS 0.014558f
C1927 VDD2.n156 VSUBS 0.015414f
C1928 VDD2.n157 VSUBS 0.034409f
C1929 VDD2.n158 VSUBS 0.034409f
C1930 VDD2.n159 VSUBS 0.015414f
C1931 VDD2.n160 VSUBS 0.014558f
C1932 VDD2.n161 VSUBS 0.027091f
C1933 VDD2.n162 VSUBS 0.027091f
C1934 VDD2.n163 VSUBS 0.014558f
C1935 VDD2.n164 VSUBS 0.014986f
C1936 VDD2.n165 VSUBS 0.014986f
C1937 VDD2.n166 VSUBS 0.034409f
C1938 VDD2.n167 VSUBS 0.034409f
C1939 VDD2.n168 VSUBS 0.015414f
C1940 VDD2.n169 VSUBS 0.014558f
C1941 VDD2.n170 VSUBS 0.027091f
C1942 VDD2.n171 VSUBS 0.027091f
C1943 VDD2.n172 VSUBS 0.014558f
C1944 VDD2.n173 VSUBS 0.015414f
C1945 VDD2.n174 VSUBS 0.034409f
C1946 VDD2.n175 VSUBS 0.034409f
C1947 VDD2.n176 VSUBS 0.015414f
C1948 VDD2.n177 VSUBS 0.014558f
C1949 VDD2.n178 VSUBS 0.027091f
C1950 VDD2.n179 VSUBS 0.027091f
C1951 VDD2.n180 VSUBS 0.014558f
C1952 VDD2.n181 VSUBS 0.015414f
C1953 VDD2.n182 VSUBS 0.034409f
C1954 VDD2.n183 VSUBS 0.034409f
C1955 VDD2.n184 VSUBS 0.015414f
C1956 VDD2.n185 VSUBS 0.014558f
C1957 VDD2.n186 VSUBS 0.027091f
C1958 VDD2.n187 VSUBS 0.027091f
C1959 VDD2.n188 VSUBS 0.014558f
C1960 VDD2.n189 VSUBS 0.015414f
C1961 VDD2.n190 VSUBS 0.034409f
C1962 VDD2.n191 VSUBS 0.034409f
C1963 VDD2.n192 VSUBS 0.015414f
C1964 VDD2.n193 VSUBS 0.014558f
C1965 VDD2.n194 VSUBS 0.027091f
C1966 VDD2.n195 VSUBS 0.027091f
C1967 VDD2.n196 VSUBS 0.014558f
C1968 VDD2.n197 VSUBS 0.015414f
C1969 VDD2.n198 VSUBS 0.034409f
C1970 VDD2.n199 VSUBS 0.034409f
C1971 VDD2.n200 VSUBS 0.015414f
C1972 VDD2.n201 VSUBS 0.014558f
C1973 VDD2.n202 VSUBS 0.027091f
C1974 VDD2.n203 VSUBS 0.027091f
C1975 VDD2.n204 VSUBS 0.014558f
C1976 VDD2.n205 VSUBS 0.015414f
C1977 VDD2.n206 VSUBS 0.034409f
C1978 VDD2.n207 VSUBS 0.083885f
C1979 VDD2.n208 VSUBS 0.015414f
C1980 VDD2.n209 VSUBS 0.028588f
C1981 VDD2.n210 VSUBS 0.065951f
C1982 VDD2.n211 VSUBS 0.082085f
C1983 VDD2.n212 VSUBS 3.69515f
C1984 VDD2.t0 VSUBS 0.415536f
C1985 VDD2.t2 VSUBS 0.415536f
C1986 VDD2.n213 VSUBS 3.50978f
C1987 VN.t4 VSUBS 4.26171f
C1988 VN.n0 VSUBS 1.5542f
C1989 VN.n1 VSUBS 0.0219f
C1990 VN.n2 VSUBS 0.032887f
C1991 VN.n3 VSUBS 0.0219f
C1992 VN.n4 VSUBS 0.03074f
C1993 VN.t2 VSUBS 4.26171f
C1994 VN.n5 VSUBS 1.54202f
C1995 VN.t1 VSUBS 4.59968f
C1996 VN.n6 VSUBS 1.47223f
C1997 VN.n7 VSUBS 0.273933f
C1998 VN.n8 VSUBS 0.0219f
C1999 VN.n9 VSUBS 0.040816f
C2000 VN.n10 VSUBS 0.040816f
C2001 VN.n11 VSUBS 0.031056f
C2002 VN.n12 VSUBS 0.0219f
C2003 VN.n13 VSUBS 0.0219f
C2004 VN.n14 VSUBS 0.0219f
C2005 VN.n15 VSUBS 0.040816f
C2006 VN.n16 VSUBS 0.040816f
C2007 VN.n17 VSUBS 0.029531f
C2008 VN.n18 VSUBS 0.035346f
C2009 VN.n19 VSUBS 0.059635f
C2010 VN.t5 VSUBS 4.26171f
C2011 VN.n20 VSUBS 1.5542f
C2012 VN.n21 VSUBS 0.0219f
C2013 VN.n22 VSUBS 0.032887f
C2014 VN.n23 VSUBS 0.0219f
C2015 VN.n24 VSUBS 0.03074f
C2016 VN.t3 VSUBS 4.59968f
C2017 VN.t0 VSUBS 4.26171f
C2018 VN.n25 VSUBS 1.54202f
C2019 VN.n26 VSUBS 1.47223f
C2020 VN.n27 VSUBS 0.273933f
C2021 VN.n28 VSUBS 0.0219f
C2022 VN.n29 VSUBS 0.040816f
C2023 VN.n30 VSUBS 0.040816f
C2024 VN.n31 VSUBS 0.031056f
C2025 VN.n32 VSUBS 0.0219f
C2026 VN.n33 VSUBS 0.0219f
C2027 VN.n34 VSUBS 0.0219f
C2028 VN.n35 VSUBS 0.040816f
C2029 VN.n36 VSUBS 0.040816f
C2030 VN.n37 VSUBS 0.029531f
C2031 VN.n38 VSUBS 0.035346f
C2032 VN.n39 VSUBS 1.56667f
.ends

