* NGSPICE file created from diff_pair_sample_0205.ext - technology: sky130A

.subckt diff_pair_sample_0205 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X1 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=0 ps=0 w=16.82 l=0.64
X2 VDD2.t6 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=2.7753 ps=17.15 w=16.82 l=0.64
X3 VTAIL.t2 VP.t0 VDD1.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X4 VDD2.t9 VN.t2 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=2.7753 ps=17.15 w=16.82 l=0.64
X5 VTAIL.t12 VN.t3 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X6 VDD1.t8 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=2.7753 ps=17.15 w=16.82 l=0.64
X7 VTAIL.t3 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X8 VDD1.t6 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X9 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=0 ps=0 w=16.82 l=0.64
X10 VDD2.t3 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X11 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=0 ps=0 w=16.82 l=0.64
X12 VDD1.t5 VP.t4 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=6.5598 ps=34.42 w=16.82 l=0.64
X13 VTAIL.t4 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X14 VDD2.t2 VN.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X15 VTAIL.t18 VP.t6 VDD1.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X16 VDD2.t1 VN.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=6.5598 ps=34.42 w=16.82 l=0.64
X17 VTAIL.t8 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X18 VTAIL.t7 VN.t8 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X19 VDD1.t2 VP.t7 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=6.5598 ps=34.42 w=16.82 l=0.64
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=0 ps=0 w=16.82 l=0.64
X21 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=2.7753 ps=17.15 w=16.82 l=0.64
X22 VDD1.t0 VP.t9 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5598 pd=34.42 as=2.7753 ps=17.15 w=16.82 l=0.64
X23 VDD2.t4 VN.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7753 pd=17.15 as=6.5598 ps=34.42 w=16.82 l=0.64
R0 VN.n2 VN.t1 721.58
R1 VN.n10 VN.t6 721.58
R2 VN.n1 VN.t7 694.759
R3 VN.n4 VN.t5 694.759
R4 VN.n5 VN.t3 694.759
R5 VN.n6 VN.t9 694.759
R6 VN.n9 VN.t0 694.759
R7 VN.n12 VN.t4 694.759
R8 VN.n13 VN.t8 694.759
R9 VN.n14 VN.t2 694.759
R10 VN.n7 VN.n6 161.3
R11 VN.n15 VN.n14 161.3
R12 VN.n13 VN.n8 80.6037
R13 VN.n12 VN.n11 80.6037
R14 VN.n5 VN.n0 80.6037
R15 VN.n4 VN.n3 80.6037
R16 VN.n4 VN.n1 48.2005
R17 VN.n5 VN.n4 48.2005
R18 VN.n6 VN.n5 48.2005
R19 VN.n12 VN.n9 48.2005
R20 VN.n13 VN.n12 48.2005
R21 VN.n14 VN.n13 48.2005
R22 VN VN.n15 46.5744
R23 VN.n11 VN.n10 45.2318
R24 VN.n3 VN.n2 45.2318
R25 VN.n10 VN.n9 13.3799
R26 VN.n2 VN.n1 13.3799
R27 VN.n11 VN.n8 0.380177
R28 VN.n3 VN.n0 0.380177
R29 VN.n15 VN.n8 0.285035
R30 VN.n7 VN.n0 0.285035
R31 VN VN.n7 0.0516364
R32 VDD2.n185 VDD2.n97 289.615
R33 VDD2.n88 VDD2.n0 289.615
R34 VDD2.n186 VDD2.n185 185
R35 VDD2.n184 VDD2.n183 185
R36 VDD2.n101 VDD2.n100 185
R37 VDD2.n178 VDD2.n177 185
R38 VDD2.n176 VDD2.n175 185
R39 VDD2.n174 VDD2.n104 185
R40 VDD2.n108 VDD2.n105 185
R41 VDD2.n169 VDD2.n168 185
R42 VDD2.n167 VDD2.n166 185
R43 VDD2.n110 VDD2.n109 185
R44 VDD2.n161 VDD2.n160 185
R45 VDD2.n159 VDD2.n158 185
R46 VDD2.n114 VDD2.n113 185
R47 VDD2.n153 VDD2.n152 185
R48 VDD2.n151 VDD2.n150 185
R49 VDD2.n118 VDD2.n117 185
R50 VDD2.n145 VDD2.n144 185
R51 VDD2.n143 VDD2.n142 185
R52 VDD2.n122 VDD2.n121 185
R53 VDD2.n137 VDD2.n136 185
R54 VDD2.n135 VDD2.n134 185
R55 VDD2.n126 VDD2.n125 185
R56 VDD2.n129 VDD2.n128 185
R57 VDD2.n31 VDD2.n30 185
R58 VDD2.n28 VDD2.n27 185
R59 VDD2.n37 VDD2.n36 185
R60 VDD2.n39 VDD2.n38 185
R61 VDD2.n24 VDD2.n23 185
R62 VDD2.n45 VDD2.n44 185
R63 VDD2.n47 VDD2.n46 185
R64 VDD2.n20 VDD2.n19 185
R65 VDD2.n53 VDD2.n52 185
R66 VDD2.n55 VDD2.n54 185
R67 VDD2.n16 VDD2.n15 185
R68 VDD2.n61 VDD2.n60 185
R69 VDD2.n63 VDD2.n62 185
R70 VDD2.n12 VDD2.n11 185
R71 VDD2.n69 VDD2.n68 185
R72 VDD2.n72 VDD2.n71 185
R73 VDD2.n70 VDD2.n8 185
R74 VDD2.n77 VDD2.n7 185
R75 VDD2.n79 VDD2.n78 185
R76 VDD2.n81 VDD2.n80 185
R77 VDD2.n4 VDD2.n3 185
R78 VDD2.n87 VDD2.n86 185
R79 VDD2.n89 VDD2.n88 185
R80 VDD2.t9 VDD2.n127 147.659
R81 VDD2.t6 VDD2.n29 147.659
R82 VDD2.n185 VDD2.n184 104.615
R83 VDD2.n184 VDD2.n100 104.615
R84 VDD2.n177 VDD2.n100 104.615
R85 VDD2.n177 VDD2.n176 104.615
R86 VDD2.n176 VDD2.n104 104.615
R87 VDD2.n108 VDD2.n104 104.615
R88 VDD2.n168 VDD2.n108 104.615
R89 VDD2.n168 VDD2.n167 104.615
R90 VDD2.n167 VDD2.n109 104.615
R91 VDD2.n160 VDD2.n109 104.615
R92 VDD2.n160 VDD2.n159 104.615
R93 VDD2.n159 VDD2.n113 104.615
R94 VDD2.n152 VDD2.n113 104.615
R95 VDD2.n152 VDD2.n151 104.615
R96 VDD2.n151 VDD2.n117 104.615
R97 VDD2.n144 VDD2.n117 104.615
R98 VDD2.n144 VDD2.n143 104.615
R99 VDD2.n143 VDD2.n121 104.615
R100 VDD2.n136 VDD2.n121 104.615
R101 VDD2.n136 VDD2.n135 104.615
R102 VDD2.n135 VDD2.n125 104.615
R103 VDD2.n128 VDD2.n125 104.615
R104 VDD2.n30 VDD2.n27 104.615
R105 VDD2.n37 VDD2.n27 104.615
R106 VDD2.n38 VDD2.n37 104.615
R107 VDD2.n38 VDD2.n23 104.615
R108 VDD2.n45 VDD2.n23 104.615
R109 VDD2.n46 VDD2.n45 104.615
R110 VDD2.n46 VDD2.n19 104.615
R111 VDD2.n53 VDD2.n19 104.615
R112 VDD2.n54 VDD2.n53 104.615
R113 VDD2.n54 VDD2.n15 104.615
R114 VDD2.n61 VDD2.n15 104.615
R115 VDD2.n62 VDD2.n61 104.615
R116 VDD2.n62 VDD2.n11 104.615
R117 VDD2.n69 VDD2.n11 104.615
R118 VDD2.n71 VDD2.n69 104.615
R119 VDD2.n71 VDD2.n70 104.615
R120 VDD2.n70 VDD2.n7 104.615
R121 VDD2.n79 VDD2.n7 104.615
R122 VDD2.n80 VDD2.n79 104.615
R123 VDD2.n80 VDD2.n3 104.615
R124 VDD2.n87 VDD2.n3 104.615
R125 VDD2.n88 VDD2.n87 104.615
R126 VDD2.n96 VDD2.n95 61.6843
R127 VDD2 VDD2.n193 61.6815
R128 VDD2.n192 VDD2.n191 61.1127
R129 VDD2.n94 VDD2.n93 61.1125
R130 VDD2.n128 VDD2.t9 52.3082
R131 VDD2.n30 VDD2.t6 52.3082
R132 VDD2.n94 VDD2.n92 50.0882
R133 VDD2.n190 VDD2.n189 49.252
R134 VDD2.n190 VDD2.n96 42.1873
R135 VDD2.n129 VDD2.n127 15.6677
R136 VDD2.n31 VDD2.n29 15.6677
R137 VDD2.n175 VDD2.n174 13.1884
R138 VDD2.n78 VDD2.n77 13.1884
R139 VDD2.n178 VDD2.n103 12.8005
R140 VDD2.n173 VDD2.n105 12.8005
R141 VDD2.n130 VDD2.n126 12.8005
R142 VDD2.n32 VDD2.n28 12.8005
R143 VDD2.n76 VDD2.n8 12.8005
R144 VDD2.n81 VDD2.n6 12.8005
R145 VDD2.n179 VDD2.n101 12.0247
R146 VDD2.n170 VDD2.n169 12.0247
R147 VDD2.n134 VDD2.n133 12.0247
R148 VDD2.n36 VDD2.n35 12.0247
R149 VDD2.n73 VDD2.n72 12.0247
R150 VDD2.n82 VDD2.n4 12.0247
R151 VDD2.n183 VDD2.n182 11.249
R152 VDD2.n166 VDD2.n107 11.249
R153 VDD2.n137 VDD2.n124 11.249
R154 VDD2.n39 VDD2.n26 11.249
R155 VDD2.n68 VDD2.n10 11.249
R156 VDD2.n86 VDD2.n85 11.249
R157 VDD2.n186 VDD2.n99 10.4732
R158 VDD2.n165 VDD2.n110 10.4732
R159 VDD2.n138 VDD2.n122 10.4732
R160 VDD2.n40 VDD2.n24 10.4732
R161 VDD2.n67 VDD2.n12 10.4732
R162 VDD2.n89 VDD2.n2 10.4732
R163 VDD2.n187 VDD2.n97 9.69747
R164 VDD2.n162 VDD2.n161 9.69747
R165 VDD2.n142 VDD2.n141 9.69747
R166 VDD2.n44 VDD2.n43 9.69747
R167 VDD2.n64 VDD2.n63 9.69747
R168 VDD2.n90 VDD2.n0 9.69747
R169 VDD2.n189 VDD2.n188 9.45567
R170 VDD2.n92 VDD2.n91 9.45567
R171 VDD2.n155 VDD2.n154 9.3005
R172 VDD2.n157 VDD2.n156 9.3005
R173 VDD2.n112 VDD2.n111 9.3005
R174 VDD2.n163 VDD2.n162 9.3005
R175 VDD2.n165 VDD2.n164 9.3005
R176 VDD2.n107 VDD2.n106 9.3005
R177 VDD2.n171 VDD2.n170 9.3005
R178 VDD2.n173 VDD2.n172 9.3005
R179 VDD2.n188 VDD2.n187 9.3005
R180 VDD2.n99 VDD2.n98 9.3005
R181 VDD2.n182 VDD2.n181 9.3005
R182 VDD2.n180 VDD2.n179 9.3005
R183 VDD2.n103 VDD2.n102 9.3005
R184 VDD2.n116 VDD2.n115 9.3005
R185 VDD2.n149 VDD2.n148 9.3005
R186 VDD2.n147 VDD2.n146 9.3005
R187 VDD2.n120 VDD2.n119 9.3005
R188 VDD2.n141 VDD2.n140 9.3005
R189 VDD2.n139 VDD2.n138 9.3005
R190 VDD2.n124 VDD2.n123 9.3005
R191 VDD2.n133 VDD2.n132 9.3005
R192 VDD2.n131 VDD2.n130 9.3005
R193 VDD2.n91 VDD2.n90 9.3005
R194 VDD2.n2 VDD2.n1 9.3005
R195 VDD2.n85 VDD2.n84 9.3005
R196 VDD2.n83 VDD2.n82 9.3005
R197 VDD2.n6 VDD2.n5 9.3005
R198 VDD2.n51 VDD2.n50 9.3005
R199 VDD2.n49 VDD2.n48 9.3005
R200 VDD2.n22 VDD2.n21 9.3005
R201 VDD2.n43 VDD2.n42 9.3005
R202 VDD2.n41 VDD2.n40 9.3005
R203 VDD2.n26 VDD2.n25 9.3005
R204 VDD2.n35 VDD2.n34 9.3005
R205 VDD2.n33 VDD2.n32 9.3005
R206 VDD2.n18 VDD2.n17 9.3005
R207 VDD2.n57 VDD2.n56 9.3005
R208 VDD2.n59 VDD2.n58 9.3005
R209 VDD2.n14 VDD2.n13 9.3005
R210 VDD2.n65 VDD2.n64 9.3005
R211 VDD2.n67 VDD2.n66 9.3005
R212 VDD2.n10 VDD2.n9 9.3005
R213 VDD2.n74 VDD2.n73 9.3005
R214 VDD2.n76 VDD2.n75 9.3005
R215 VDD2.n158 VDD2.n112 8.92171
R216 VDD2.n145 VDD2.n120 8.92171
R217 VDD2.n47 VDD2.n22 8.92171
R218 VDD2.n60 VDD2.n14 8.92171
R219 VDD2.n157 VDD2.n114 8.14595
R220 VDD2.n146 VDD2.n118 8.14595
R221 VDD2.n48 VDD2.n20 8.14595
R222 VDD2.n59 VDD2.n16 8.14595
R223 VDD2.n154 VDD2.n153 7.3702
R224 VDD2.n150 VDD2.n149 7.3702
R225 VDD2.n52 VDD2.n51 7.3702
R226 VDD2.n56 VDD2.n55 7.3702
R227 VDD2.n153 VDD2.n116 6.59444
R228 VDD2.n150 VDD2.n116 6.59444
R229 VDD2.n52 VDD2.n18 6.59444
R230 VDD2.n55 VDD2.n18 6.59444
R231 VDD2.n154 VDD2.n114 5.81868
R232 VDD2.n149 VDD2.n118 5.81868
R233 VDD2.n51 VDD2.n20 5.81868
R234 VDD2.n56 VDD2.n16 5.81868
R235 VDD2.n158 VDD2.n157 5.04292
R236 VDD2.n146 VDD2.n145 5.04292
R237 VDD2.n48 VDD2.n47 5.04292
R238 VDD2.n60 VDD2.n59 5.04292
R239 VDD2.n131 VDD2.n127 4.38563
R240 VDD2.n33 VDD2.n29 4.38563
R241 VDD2.n189 VDD2.n97 4.26717
R242 VDD2.n161 VDD2.n112 4.26717
R243 VDD2.n142 VDD2.n120 4.26717
R244 VDD2.n44 VDD2.n22 4.26717
R245 VDD2.n63 VDD2.n14 4.26717
R246 VDD2.n92 VDD2.n0 4.26717
R247 VDD2.n187 VDD2.n186 3.49141
R248 VDD2.n162 VDD2.n110 3.49141
R249 VDD2.n141 VDD2.n122 3.49141
R250 VDD2.n43 VDD2.n24 3.49141
R251 VDD2.n64 VDD2.n12 3.49141
R252 VDD2.n90 VDD2.n89 3.49141
R253 VDD2.n183 VDD2.n99 2.71565
R254 VDD2.n166 VDD2.n165 2.71565
R255 VDD2.n138 VDD2.n137 2.71565
R256 VDD2.n40 VDD2.n39 2.71565
R257 VDD2.n68 VDD2.n67 2.71565
R258 VDD2.n86 VDD2.n2 2.71565
R259 VDD2.n182 VDD2.n101 1.93989
R260 VDD2.n169 VDD2.n107 1.93989
R261 VDD2.n134 VDD2.n124 1.93989
R262 VDD2.n36 VDD2.n26 1.93989
R263 VDD2.n72 VDD2.n10 1.93989
R264 VDD2.n85 VDD2.n4 1.93989
R265 VDD2.n193 VDD2.t7 1.17767
R266 VDD2.n193 VDD2.t1 1.17767
R267 VDD2.n191 VDD2.t5 1.17767
R268 VDD2.n191 VDD2.t3 1.17767
R269 VDD2.n95 VDD2.t8 1.17767
R270 VDD2.n95 VDD2.t4 1.17767
R271 VDD2.n93 VDD2.t0 1.17767
R272 VDD2.n93 VDD2.t2 1.17767
R273 VDD2.n179 VDD2.n178 1.16414
R274 VDD2.n170 VDD2.n105 1.16414
R275 VDD2.n133 VDD2.n126 1.16414
R276 VDD2.n35 VDD2.n28 1.16414
R277 VDD2.n73 VDD2.n8 1.16414
R278 VDD2.n82 VDD2.n81 1.16414
R279 VDD2.n192 VDD2.n190 0.836707
R280 VDD2.n175 VDD2.n103 0.388379
R281 VDD2.n174 VDD2.n173 0.388379
R282 VDD2.n130 VDD2.n129 0.388379
R283 VDD2.n32 VDD2.n31 0.388379
R284 VDD2.n77 VDD2.n76 0.388379
R285 VDD2.n78 VDD2.n6 0.388379
R286 VDD2 VDD2.n192 0.267741
R287 VDD2.n188 VDD2.n98 0.155672
R288 VDD2.n181 VDD2.n98 0.155672
R289 VDD2.n181 VDD2.n180 0.155672
R290 VDD2.n180 VDD2.n102 0.155672
R291 VDD2.n172 VDD2.n102 0.155672
R292 VDD2.n172 VDD2.n171 0.155672
R293 VDD2.n171 VDD2.n106 0.155672
R294 VDD2.n164 VDD2.n106 0.155672
R295 VDD2.n164 VDD2.n163 0.155672
R296 VDD2.n163 VDD2.n111 0.155672
R297 VDD2.n156 VDD2.n111 0.155672
R298 VDD2.n156 VDD2.n155 0.155672
R299 VDD2.n155 VDD2.n115 0.155672
R300 VDD2.n148 VDD2.n115 0.155672
R301 VDD2.n148 VDD2.n147 0.155672
R302 VDD2.n147 VDD2.n119 0.155672
R303 VDD2.n140 VDD2.n119 0.155672
R304 VDD2.n140 VDD2.n139 0.155672
R305 VDD2.n139 VDD2.n123 0.155672
R306 VDD2.n132 VDD2.n123 0.155672
R307 VDD2.n132 VDD2.n131 0.155672
R308 VDD2.n34 VDD2.n33 0.155672
R309 VDD2.n34 VDD2.n25 0.155672
R310 VDD2.n41 VDD2.n25 0.155672
R311 VDD2.n42 VDD2.n41 0.155672
R312 VDD2.n42 VDD2.n21 0.155672
R313 VDD2.n49 VDD2.n21 0.155672
R314 VDD2.n50 VDD2.n49 0.155672
R315 VDD2.n50 VDD2.n17 0.155672
R316 VDD2.n57 VDD2.n17 0.155672
R317 VDD2.n58 VDD2.n57 0.155672
R318 VDD2.n58 VDD2.n13 0.155672
R319 VDD2.n65 VDD2.n13 0.155672
R320 VDD2.n66 VDD2.n65 0.155672
R321 VDD2.n66 VDD2.n9 0.155672
R322 VDD2.n74 VDD2.n9 0.155672
R323 VDD2.n75 VDD2.n74 0.155672
R324 VDD2.n75 VDD2.n5 0.155672
R325 VDD2.n83 VDD2.n5 0.155672
R326 VDD2.n84 VDD2.n83 0.155672
R327 VDD2.n84 VDD2.n1 0.155672
R328 VDD2.n91 VDD2.n1 0.155672
R329 VDD2.n96 VDD2.n94 0.154206
R330 VTAIL.n384 VTAIL.n296 289.615
R331 VTAIL.n90 VTAIL.n2 289.615
R332 VTAIL.n290 VTAIL.n202 289.615
R333 VTAIL.n192 VTAIL.n104 289.615
R334 VTAIL.n327 VTAIL.n326 185
R335 VTAIL.n324 VTAIL.n323 185
R336 VTAIL.n333 VTAIL.n332 185
R337 VTAIL.n335 VTAIL.n334 185
R338 VTAIL.n320 VTAIL.n319 185
R339 VTAIL.n341 VTAIL.n340 185
R340 VTAIL.n343 VTAIL.n342 185
R341 VTAIL.n316 VTAIL.n315 185
R342 VTAIL.n349 VTAIL.n348 185
R343 VTAIL.n351 VTAIL.n350 185
R344 VTAIL.n312 VTAIL.n311 185
R345 VTAIL.n357 VTAIL.n356 185
R346 VTAIL.n359 VTAIL.n358 185
R347 VTAIL.n308 VTAIL.n307 185
R348 VTAIL.n365 VTAIL.n364 185
R349 VTAIL.n368 VTAIL.n367 185
R350 VTAIL.n366 VTAIL.n304 185
R351 VTAIL.n373 VTAIL.n303 185
R352 VTAIL.n375 VTAIL.n374 185
R353 VTAIL.n377 VTAIL.n376 185
R354 VTAIL.n300 VTAIL.n299 185
R355 VTAIL.n383 VTAIL.n382 185
R356 VTAIL.n385 VTAIL.n384 185
R357 VTAIL.n33 VTAIL.n32 185
R358 VTAIL.n30 VTAIL.n29 185
R359 VTAIL.n39 VTAIL.n38 185
R360 VTAIL.n41 VTAIL.n40 185
R361 VTAIL.n26 VTAIL.n25 185
R362 VTAIL.n47 VTAIL.n46 185
R363 VTAIL.n49 VTAIL.n48 185
R364 VTAIL.n22 VTAIL.n21 185
R365 VTAIL.n55 VTAIL.n54 185
R366 VTAIL.n57 VTAIL.n56 185
R367 VTAIL.n18 VTAIL.n17 185
R368 VTAIL.n63 VTAIL.n62 185
R369 VTAIL.n65 VTAIL.n64 185
R370 VTAIL.n14 VTAIL.n13 185
R371 VTAIL.n71 VTAIL.n70 185
R372 VTAIL.n74 VTAIL.n73 185
R373 VTAIL.n72 VTAIL.n10 185
R374 VTAIL.n79 VTAIL.n9 185
R375 VTAIL.n81 VTAIL.n80 185
R376 VTAIL.n83 VTAIL.n82 185
R377 VTAIL.n6 VTAIL.n5 185
R378 VTAIL.n89 VTAIL.n88 185
R379 VTAIL.n91 VTAIL.n90 185
R380 VTAIL.n291 VTAIL.n290 185
R381 VTAIL.n289 VTAIL.n288 185
R382 VTAIL.n206 VTAIL.n205 185
R383 VTAIL.n283 VTAIL.n282 185
R384 VTAIL.n281 VTAIL.n280 185
R385 VTAIL.n279 VTAIL.n209 185
R386 VTAIL.n213 VTAIL.n210 185
R387 VTAIL.n274 VTAIL.n273 185
R388 VTAIL.n272 VTAIL.n271 185
R389 VTAIL.n215 VTAIL.n214 185
R390 VTAIL.n266 VTAIL.n265 185
R391 VTAIL.n264 VTAIL.n263 185
R392 VTAIL.n219 VTAIL.n218 185
R393 VTAIL.n258 VTAIL.n257 185
R394 VTAIL.n256 VTAIL.n255 185
R395 VTAIL.n223 VTAIL.n222 185
R396 VTAIL.n250 VTAIL.n249 185
R397 VTAIL.n248 VTAIL.n247 185
R398 VTAIL.n227 VTAIL.n226 185
R399 VTAIL.n242 VTAIL.n241 185
R400 VTAIL.n240 VTAIL.n239 185
R401 VTAIL.n231 VTAIL.n230 185
R402 VTAIL.n234 VTAIL.n233 185
R403 VTAIL.n193 VTAIL.n192 185
R404 VTAIL.n191 VTAIL.n190 185
R405 VTAIL.n108 VTAIL.n107 185
R406 VTAIL.n185 VTAIL.n184 185
R407 VTAIL.n183 VTAIL.n182 185
R408 VTAIL.n181 VTAIL.n111 185
R409 VTAIL.n115 VTAIL.n112 185
R410 VTAIL.n176 VTAIL.n175 185
R411 VTAIL.n174 VTAIL.n173 185
R412 VTAIL.n117 VTAIL.n116 185
R413 VTAIL.n168 VTAIL.n167 185
R414 VTAIL.n166 VTAIL.n165 185
R415 VTAIL.n121 VTAIL.n120 185
R416 VTAIL.n160 VTAIL.n159 185
R417 VTAIL.n158 VTAIL.n157 185
R418 VTAIL.n125 VTAIL.n124 185
R419 VTAIL.n152 VTAIL.n151 185
R420 VTAIL.n150 VTAIL.n149 185
R421 VTAIL.n129 VTAIL.n128 185
R422 VTAIL.n144 VTAIL.n143 185
R423 VTAIL.n142 VTAIL.n141 185
R424 VTAIL.n133 VTAIL.n132 185
R425 VTAIL.n136 VTAIL.n135 185
R426 VTAIL.t17 VTAIL.n232 147.659
R427 VTAIL.t9 VTAIL.n134 147.659
R428 VTAIL.t6 VTAIL.n325 147.659
R429 VTAIL.t16 VTAIL.n31 147.659
R430 VTAIL.n326 VTAIL.n323 104.615
R431 VTAIL.n333 VTAIL.n323 104.615
R432 VTAIL.n334 VTAIL.n333 104.615
R433 VTAIL.n334 VTAIL.n319 104.615
R434 VTAIL.n341 VTAIL.n319 104.615
R435 VTAIL.n342 VTAIL.n341 104.615
R436 VTAIL.n342 VTAIL.n315 104.615
R437 VTAIL.n349 VTAIL.n315 104.615
R438 VTAIL.n350 VTAIL.n349 104.615
R439 VTAIL.n350 VTAIL.n311 104.615
R440 VTAIL.n357 VTAIL.n311 104.615
R441 VTAIL.n358 VTAIL.n357 104.615
R442 VTAIL.n358 VTAIL.n307 104.615
R443 VTAIL.n365 VTAIL.n307 104.615
R444 VTAIL.n367 VTAIL.n365 104.615
R445 VTAIL.n367 VTAIL.n366 104.615
R446 VTAIL.n366 VTAIL.n303 104.615
R447 VTAIL.n375 VTAIL.n303 104.615
R448 VTAIL.n376 VTAIL.n375 104.615
R449 VTAIL.n376 VTAIL.n299 104.615
R450 VTAIL.n383 VTAIL.n299 104.615
R451 VTAIL.n384 VTAIL.n383 104.615
R452 VTAIL.n32 VTAIL.n29 104.615
R453 VTAIL.n39 VTAIL.n29 104.615
R454 VTAIL.n40 VTAIL.n39 104.615
R455 VTAIL.n40 VTAIL.n25 104.615
R456 VTAIL.n47 VTAIL.n25 104.615
R457 VTAIL.n48 VTAIL.n47 104.615
R458 VTAIL.n48 VTAIL.n21 104.615
R459 VTAIL.n55 VTAIL.n21 104.615
R460 VTAIL.n56 VTAIL.n55 104.615
R461 VTAIL.n56 VTAIL.n17 104.615
R462 VTAIL.n63 VTAIL.n17 104.615
R463 VTAIL.n64 VTAIL.n63 104.615
R464 VTAIL.n64 VTAIL.n13 104.615
R465 VTAIL.n71 VTAIL.n13 104.615
R466 VTAIL.n73 VTAIL.n71 104.615
R467 VTAIL.n73 VTAIL.n72 104.615
R468 VTAIL.n72 VTAIL.n9 104.615
R469 VTAIL.n81 VTAIL.n9 104.615
R470 VTAIL.n82 VTAIL.n81 104.615
R471 VTAIL.n82 VTAIL.n5 104.615
R472 VTAIL.n89 VTAIL.n5 104.615
R473 VTAIL.n90 VTAIL.n89 104.615
R474 VTAIL.n290 VTAIL.n289 104.615
R475 VTAIL.n289 VTAIL.n205 104.615
R476 VTAIL.n282 VTAIL.n205 104.615
R477 VTAIL.n282 VTAIL.n281 104.615
R478 VTAIL.n281 VTAIL.n209 104.615
R479 VTAIL.n213 VTAIL.n209 104.615
R480 VTAIL.n273 VTAIL.n213 104.615
R481 VTAIL.n273 VTAIL.n272 104.615
R482 VTAIL.n272 VTAIL.n214 104.615
R483 VTAIL.n265 VTAIL.n214 104.615
R484 VTAIL.n265 VTAIL.n264 104.615
R485 VTAIL.n264 VTAIL.n218 104.615
R486 VTAIL.n257 VTAIL.n218 104.615
R487 VTAIL.n257 VTAIL.n256 104.615
R488 VTAIL.n256 VTAIL.n222 104.615
R489 VTAIL.n249 VTAIL.n222 104.615
R490 VTAIL.n249 VTAIL.n248 104.615
R491 VTAIL.n248 VTAIL.n226 104.615
R492 VTAIL.n241 VTAIL.n226 104.615
R493 VTAIL.n241 VTAIL.n240 104.615
R494 VTAIL.n240 VTAIL.n230 104.615
R495 VTAIL.n233 VTAIL.n230 104.615
R496 VTAIL.n192 VTAIL.n191 104.615
R497 VTAIL.n191 VTAIL.n107 104.615
R498 VTAIL.n184 VTAIL.n107 104.615
R499 VTAIL.n184 VTAIL.n183 104.615
R500 VTAIL.n183 VTAIL.n111 104.615
R501 VTAIL.n115 VTAIL.n111 104.615
R502 VTAIL.n175 VTAIL.n115 104.615
R503 VTAIL.n175 VTAIL.n174 104.615
R504 VTAIL.n174 VTAIL.n116 104.615
R505 VTAIL.n167 VTAIL.n116 104.615
R506 VTAIL.n167 VTAIL.n166 104.615
R507 VTAIL.n166 VTAIL.n120 104.615
R508 VTAIL.n159 VTAIL.n120 104.615
R509 VTAIL.n159 VTAIL.n158 104.615
R510 VTAIL.n158 VTAIL.n124 104.615
R511 VTAIL.n151 VTAIL.n124 104.615
R512 VTAIL.n151 VTAIL.n150 104.615
R513 VTAIL.n150 VTAIL.n128 104.615
R514 VTAIL.n143 VTAIL.n128 104.615
R515 VTAIL.n143 VTAIL.n142 104.615
R516 VTAIL.n142 VTAIL.n132 104.615
R517 VTAIL.n135 VTAIL.n132 104.615
R518 VTAIL.n326 VTAIL.t6 52.3082
R519 VTAIL.n32 VTAIL.t16 52.3082
R520 VTAIL.n233 VTAIL.t17 52.3082
R521 VTAIL.n135 VTAIL.t9 52.3082
R522 VTAIL.n201 VTAIL.n200 44.4339
R523 VTAIL.n199 VTAIL.n198 44.4339
R524 VTAIL.n103 VTAIL.n102 44.4339
R525 VTAIL.n101 VTAIL.n100 44.4339
R526 VTAIL.n391 VTAIL.n390 44.4337
R527 VTAIL.n1 VTAIL.n0 44.4337
R528 VTAIL.n97 VTAIL.n96 44.4337
R529 VTAIL.n99 VTAIL.n98 44.4337
R530 VTAIL.n389 VTAIL.n388 32.5732
R531 VTAIL.n95 VTAIL.n94 32.5732
R532 VTAIL.n295 VTAIL.n294 32.5732
R533 VTAIL.n197 VTAIL.n196 32.5732
R534 VTAIL.n101 VTAIL.n99 28.5393
R535 VTAIL.n389 VTAIL.n295 27.7031
R536 VTAIL.n327 VTAIL.n325 15.6677
R537 VTAIL.n33 VTAIL.n31 15.6677
R538 VTAIL.n234 VTAIL.n232 15.6677
R539 VTAIL.n136 VTAIL.n134 15.6677
R540 VTAIL.n374 VTAIL.n373 13.1884
R541 VTAIL.n80 VTAIL.n79 13.1884
R542 VTAIL.n280 VTAIL.n279 13.1884
R543 VTAIL.n182 VTAIL.n181 13.1884
R544 VTAIL.n328 VTAIL.n324 12.8005
R545 VTAIL.n372 VTAIL.n304 12.8005
R546 VTAIL.n377 VTAIL.n302 12.8005
R547 VTAIL.n34 VTAIL.n30 12.8005
R548 VTAIL.n78 VTAIL.n10 12.8005
R549 VTAIL.n83 VTAIL.n8 12.8005
R550 VTAIL.n283 VTAIL.n208 12.8005
R551 VTAIL.n278 VTAIL.n210 12.8005
R552 VTAIL.n235 VTAIL.n231 12.8005
R553 VTAIL.n185 VTAIL.n110 12.8005
R554 VTAIL.n180 VTAIL.n112 12.8005
R555 VTAIL.n137 VTAIL.n133 12.8005
R556 VTAIL.n332 VTAIL.n331 12.0247
R557 VTAIL.n369 VTAIL.n368 12.0247
R558 VTAIL.n378 VTAIL.n300 12.0247
R559 VTAIL.n38 VTAIL.n37 12.0247
R560 VTAIL.n75 VTAIL.n74 12.0247
R561 VTAIL.n84 VTAIL.n6 12.0247
R562 VTAIL.n284 VTAIL.n206 12.0247
R563 VTAIL.n275 VTAIL.n274 12.0247
R564 VTAIL.n239 VTAIL.n238 12.0247
R565 VTAIL.n186 VTAIL.n108 12.0247
R566 VTAIL.n177 VTAIL.n176 12.0247
R567 VTAIL.n141 VTAIL.n140 12.0247
R568 VTAIL.n335 VTAIL.n322 11.249
R569 VTAIL.n364 VTAIL.n306 11.249
R570 VTAIL.n382 VTAIL.n381 11.249
R571 VTAIL.n41 VTAIL.n28 11.249
R572 VTAIL.n70 VTAIL.n12 11.249
R573 VTAIL.n88 VTAIL.n87 11.249
R574 VTAIL.n288 VTAIL.n287 11.249
R575 VTAIL.n271 VTAIL.n212 11.249
R576 VTAIL.n242 VTAIL.n229 11.249
R577 VTAIL.n190 VTAIL.n189 11.249
R578 VTAIL.n173 VTAIL.n114 11.249
R579 VTAIL.n144 VTAIL.n131 11.249
R580 VTAIL.n336 VTAIL.n320 10.4732
R581 VTAIL.n363 VTAIL.n308 10.4732
R582 VTAIL.n385 VTAIL.n298 10.4732
R583 VTAIL.n42 VTAIL.n26 10.4732
R584 VTAIL.n69 VTAIL.n14 10.4732
R585 VTAIL.n91 VTAIL.n4 10.4732
R586 VTAIL.n291 VTAIL.n204 10.4732
R587 VTAIL.n270 VTAIL.n215 10.4732
R588 VTAIL.n243 VTAIL.n227 10.4732
R589 VTAIL.n193 VTAIL.n106 10.4732
R590 VTAIL.n172 VTAIL.n117 10.4732
R591 VTAIL.n145 VTAIL.n129 10.4732
R592 VTAIL.n340 VTAIL.n339 9.69747
R593 VTAIL.n360 VTAIL.n359 9.69747
R594 VTAIL.n386 VTAIL.n296 9.69747
R595 VTAIL.n46 VTAIL.n45 9.69747
R596 VTAIL.n66 VTAIL.n65 9.69747
R597 VTAIL.n92 VTAIL.n2 9.69747
R598 VTAIL.n292 VTAIL.n202 9.69747
R599 VTAIL.n267 VTAIL.n266 9.69747
R600 VTAIL.n247 VTAIL.n246 9.69747
R601 VTAIL.n194 VTAIL.n104 9.69747
R602 VTAIL.n169 VTAIL.n168 9.69747
R603 VTAIL.n149 VTAIL.n148 9.69747
R604 VTAIL.n388 VTAIL.n387 9.45567
R605 VTAIL.n94 VTAIL.n93 9.45567
R606 VTAIL.n294 VTAIL.n293 9.45567
R607 VTAIL.n196 VTAIL.n195 9.45567
R608 VTAIL.n387 VTAIL.n386 9.3005
R609 VTAIL.n298 VTAIL.n297 9.3005
R610 VTAIL.n381 VTAIL.n380 9.3005
R611 VTAIL.n379 VTAIL.n378 9.3005
R612 VTAIL.n302 VTAIL.n301 9.3005
R613 VTAIL.n347 VTAIL.n346 9.3005
R614 VTAIL.n345 VTAIL.n344 9.3005
R615 VTAIL.n318 VTAIL.n317 9.3005
R616 VTAIL.n339 VTAIL.n338 9.3005
R617 VTAIL.n337 VTAIL.n336 9.3005
R618 VTAIL.n322 VTAIL.n321 9.3005
R619 VTAIL.n331 VTAIL.n330 9.3005
R620 VTAIL.n329 VTAIL.n328 9.3005
R621 VTAIL.n314 VTAIL.n313 9.3005
R622 VTAIL.n353 VTAIL.n352 9.3005
R623 VTAIL.n355 VTAIL.n354 9.3005
R624 VTAIL.n310 VTAIL.n309 9.3005
R625 VTAIL.n361 VTAIL.n360 9.3005
R626 VTAIL.n363 VTAIL.n362 9.3005
R627 VTAIL.n306 VTAIL.n305 9.3005
R628 VTAIL.n370 VTAIL.n369 9.3005
R629 VTAIL.n372 VTAIL.n371 9.3005
R630 VTAIL.n93 VTAIL.n92 9.3005
R631 VTAIL.n4 VTAIL.n3 9.3005
R632 VTAIL.n87 VTAIL.n86 9.3005
R633 VTAIL.n85 VTAIL.n84 9.3005
R634 VTAIL.n8 VTAIL.n7 9.3005
R635 VTAIL.n53 VTAIL.n52 9.3005
R636 VTAIL.n51 VTAIL.n50 9.3005
R637 VTAIL.n24 VTAIL.n23 9.3005
R638 VTAIL.n45 VTAIL.n44 9.3005
R639 VTAIL.n43 VTAIL.n42 9.3005
R640 VTAIL.n28 VTAIL.n27 9.3005
R641 VTAIL.n37 VTAIL.n36 9.3005
R642 VTAIL.n35 VTAIL.n34 9.3005
R643 VTAIL.n20 VTAIL.n19 9.3005
R644 VTAIL.n59 VTAIL.n58 9.3005
R645 VTAIL.n61 VTAIL.n60 9.3005
R646 VTAIL.n16 VTAIL.n15 9.3005
R647 VTAIL.n67 VTAIL.n66 9.3005
R648 VTAIL.n69 VTAIL.n68 9.3005
R649 VTAIL.n12 VTAIL.n11 9.3005
R650 VTAIL.n76 VTAIL.n75 9.3005
R651 VTAIL.n78 VTAIL.n77 9.3005
R652 VTAIL.n260 VTAIL.n259 9.3005
R653 VTAIL.n262 VTAIL.n261 9.3005
R654 VTAIL.n217 VTAIL.n216 9.3005
R655 VTAIL.n268 VTAIL.n267 9.3005
R656 VTAIL.n270 VTAIL.n269 9.3005
R657 VTAIL.n212 VTAIL.n211 9.3005
R658 VTAIL.n276 VTAIL.n275 9.3005
R659 VTAIL.n278 VTAIL.n277 9.3005
R660 VTAIL.n293 VTAIL.n292 9.3005
R661 VTAIL.n204 VTAIL.n203 9.3005
R662 VTAIL.n287 VTAIL.n286 9.3005
R663 VTAIL.n285 VTAIL.n284 9.3005
R664 VTAIL.n208 VTAIL.n207 9.3005
R665 VTAIL.n221 VTAIL.n220 9.3005
R666 VTAIL.n254 VTAIL.n253 9.3005
R667 VTAIL.n252 VTAIL.n251 9.3005
R668 VTAIL.n225 VTAIL.n224 9.3005
R669 VTAIL.n246 VTAIL.n245 9.3005
R670 VTAIL.n244 VTAIL.n243 9.3005
R671 VTAIL.n229 VTAIL.n228 9.3005
R672 VTAIL.n238 VTAIL.n237 9.3005
R673 VTAIL.n236 VTAIL.n235 9.3005
R674 VTAIL.n162 VTAIL.n161 9.3005
R675 VTAIL.n164 VTAIL.n163 9.3005
R676 VTAIL.n119 VTAIL.n118 9.3005
R677 VTAIL.n170 VTAIL.n169 9.3005
R678 VTAIL.n172 VTAIL.n171 9.3005
R679 VTAIL.n114 VTAIL.n113 9.3005
R680 VTAIL.n178 VTAIL.n177 9.3005
R681 VTAIL.n180 VTAIL.n179 9.3005
R682 VTAIL.n195 VTAIL.n194 9.3005
R683 VTAIL.n106 VTAIL.n105 9.3005
R684 VTAIL.n189 VTAIL.n188 9.3005
R685 VTAIL.n187 VTAIL.n186 9.3005
R686 VTAIL.n110 VTAIL.n109 9.3005
R687 VTAIL.n123 VTAIL.n122 9.3005
R688 VTAIL.n156 VTAIL.n155 9.3005
R689 VTAIL.n154 VTAIL.n153 9.3005
R690 VTAIL.n127 VTAIL.n126 9.3005
R691 VTAIL.n148 VTAIL.n147 9.3005
R692 VTAIL.n146 VTAIL.n145 9.3005
R693 VTAIL.n131 VTAIL.n130 9.3005
R694 VTAIL.n140 VTAIL.n139 9.3005
R695 VTAIL.n138 VTAIL.n137 9.3005
R696 VTAIL.n343 VTAIL.n318 8.92171
R697 VTAIL.n356 VTAIL.n310 8.92171
R698 VTAIL.n49 VTAIL.n24 8.92171
R699 VTAIL.n62 VTAIL.n16 8.92171
R700 VTAIL.n263 VTAIL.n217 8.92171
R701 VTAIL.n250 VTAIL.n225 8.92171
R702 VTAIL.n165 VTAIL.n119 8.92171
R703 VTAIL.n152 VTAIL.n127 8.92171
R704 VTAIL.n344 VTAIL.n316 8.14595
R705 VTAIL.n355 VTAIL.n312 8.14595
R706 VTAIL.n50 VTAIL.n22 8.14595
R707 VTAIL.n61 VTAIL.n18 8.14595
R708 VTAIL.n262 VTAIL.n219 8.14595
R709 VTAIL.n251 VTAIL.n223 8.14595
R710 VTAIL.n164 VTAIL.n121 8.14595
R711 VTAIL.n153 VTAIL.n125 8.14595
R712 VTAIL.n348 VTAIL.n347 7.3702
R713 VTAIL.n352 VTAIL.n351 7.3702
R714 VTAIL.n54 VTAIL.n53 7.3702
R715 VTAIL.n58 VTAIL.n57 7.3702
R716 VTAIL.n259 VTAIL.n258 7.3702
R717 VTAIL.n255 VTAIL.n254 7.3702
R718 VTAIL.n161 VTAIL.n160 7.3702
R719 VTAIL.n157 VTAIL.n156 7.3702
R720 VTAIL.n348 VTAIL.n314 6.59444
R721 VTAIL.n351 VTAIL.n314 6.59444
R722 VTAIL.n54 VTAIL.n20 6.59444
R723 VTAIL.n57 VTAIL.n20 6.59444
R724 VTAIL.n258 VTAIL.n221 6.59444
R725 VTAIL.n255 VTAIL.n221 6.59444
R726 VTAIL.n160 VTAIL.n123 6.59444
R727 VTAIL.n157 VTAIL.n123 6.59444
R728 VTAIL.n347 VTAIL.n316 5.81868
R729 VTAIL.n352 VTAIL.n312 5.81868
R730 VTAIL.n53 VTAIL.n22 5.81868
R731 VTAIL.n58 VTAIL.n18 5.81868
R732 VTAIL.n259 VTAIL.n219 5.81868
R733 VTAIL.n254 VTAIL.n223 5.81868
R734 VTAIL.n161 VTAIL.n121 5.81868
R735 VTAIL.n156 VTAIL.n125 5.81868
R736 VTAIL.n344 VTAIL.n343 5.04292
R737 VTAIL.n356 VTAIL.n355 5.04292
R738 VTAIL.n50 VTAIL.n49 5.04292
R739 VTAIL.n62 VTAIL.n61 5.04292
R740 VTAIL.n263 VTAIL.n262 5.04292
R741 VTAIL.n251 VTAIL.n250 5.04292
R742 VTAIL.n165 VTAIL.n164 5.04292
R743 VTAIL.n153 VTAIL.n152 5.04292
R744 VTAIL.n236 VTAIL.n232 4.38563
R745 VTAIL.n138 VTAIL.n134 4.38563
R746 VTAIL.n329 VTAIL.n325 4.38563
R747 VTAIL.n35 VTAIL.n31 4.38563
R748 VTAIL.n340 VTAIL.n318 4.26717
R749 VTAIL.n359 VTAIL.n310 4.26717
R750 VTAIL.n388 VTAIL.n296 4.26717
R751 VTAIL.n46 VTAIL.n24 4.26717
R752 VTAIL.n65 VTAIL.n16 4.26717
R753 VTAIL.n94 VTAIL.n2 4.26717
R754 VTAIL.n294 VTAIL.n202 4.26717
R755 VTAIL.n266 VTAIL.n217 4.26717
R756 VTAIL.n247 VTAIL.n225 4.26717
R757 VTAIL.n196 VTAIL.n104 4.26717
R758 VTAIL.n168 VTAIL.n119 4.26717
R759 VTAIL.n149 VTAIL.n127 4.26717
R760 VTAIL.n339 VTAIL.n320 3.49141
R761 VTAIL.n360 VTAIL.n308 3.49141
R762 VTAIL.n386 VTAIL.n385 3.49141
R763 VTAIL.n45 VTAIL.n26 3.49141
R764 VTAIL.n66 VTAIL.n14 3.49141
R765 VTAIL.n92 VTAIL.n91 3.49141
R766 VTAIL.n292 VTAIL.n291 3.49141
R767 VTAIL.n267 VTAIL.n215 3.49141
R768 VTAIL.n246 VTAIL.n227 3.49141
R769 VTAIL.n194 VTAIL.n193 3.49141
R770 VTAIL.n169 VTAIL.n117 3.49141
R771 VTAIL.n148 VTAIL.n129 3.49141
R772 VTAIL.n336 VTAIL.n335 2.71565
R773 VTAIL.n364 VTAIL.n363 2.71565
R774 VTAIL.n382 VTAIL.n298 2.71565
R775 VTAIL.n42 VTAIL.n41 2.71565
R776 VTAIL.n70 VTAIL.n69 2.71565
R777 VTAIL.n88 VTAIL.n4 2.71565
R778 VTAIL.n288 VTAIL.n204 2.71565
R779 VTAIL.n271 VTAIL.n270 2.71565
R780 VTAIL.n243 VTAIL.n242 2.71565
R781 VTAIL.n190 VTAIL.n106 2.71565
R782 VTAIL.n173 VTAIL.n172 2.71565
R783 VTAIL.n145 VTAIL.n144 2.71565
R784 VTAIL.n332 VTAIL.n322 1.93989
R785 VTAIL.n368 VTAIL.n306 1.93989
R786 VTAIL.n381 VTAIL.n300 1.93989
R787 VTAIL.n38 VTAIL.n28 1.93989
R788 VTAIL.n74 VTAIL.n12 1.93989
R789 VTAIL.n87 VTAIL.n6 1.93989
R790 VTAIL.n287 VTAIL.n206 1.93989
R791 VTAIL.n274 VTAIL.n212 1.93989
R792 VTAIL.n239 VTAIL.n229 1.93989
R793 VTAIL.n189 VTAIL.n108 1.93989
R794 VTAIL.n176 VTAIL.n114 1.93989
R795 VTAIL.n141 VTAIL.n131 1.93989
R796 VTAIL.n390 VTAIL.t10 1.17767
R797 VTAIL.n390 VTAIL.t12 1.17767
R798 VTAIL.n0 VTAIL.t14 1.17767
R799 VTAIL.n0 VTAIL.t8 1.17767
R800 VTAIL.n96 VTAIL.t5 1.17767
R801 VTAIL.n96 VTAIL.t18 1.17767
R802 VTAIL.n98 VTAIL.t19 1.17767
R803 VTAIL.n98 VTAIL.t2 1.17767
R804 VTAIL.n200 VTAIL.t0 1.17767
R805 VTAIL.n200 VTAIL.t3 1.17767
R806 VTAIL.n198 VTAIL.t1 1.17767
R807 VTAIL.n198 VTAIL.t4 1.17767
R808 VTAIL.n102 VTAIL.t11 1.17767
R809 VTAIL.n102 VTAIL.t15 1.17767
R810 VTAIL.n100 VTAIL.t13 1.17767
R811 VTAIL.n100 VTAIL.t7 1.17767
R812 VTAIL.n331 VTAIL.n324 1.16414
R813 VTAIL.n369 VTAIL.n304 1.16414
R814 VTAIL.n378 VTAIL.n377 1.16414
R815 VTAIL.n37 VTAIL.n30 1.16414
R816 VTAIL.n75 VTAIL.n10 1.16414
R817 VTAIL.n84 VTAIL.n83 1.16414
R818 VTAIL.n284 VTAIL.n283 1.16414
R819 VTAIL.n275 VTAIL.n210 1.16414
R820 VTAIL.n238 VTAIL.n231 1.16414
R821 VTAIL.n186 VTAIL.n185 1.16414
R822 VTAIL.n177 VTAIL.n112 1.16414
R823 VTAIL.n140 VTAIL.n133 1.16414
R824 VTAIL.n199 VTAIL.n197 0.888431
R825 VTAIL.n95 VTAIL.n1 0.888431
R826 VTAIL.n103 VTAIL.n101 0.836707
R827 VTAIL.n197 VTAIL.n103 0.836707
R828 VTAIL.n201 VTAIL.n199 0.836707
R829 VTAIL.n295 VTAIL.n201 0.836707
R830 VTAIL.n99 VTAIL.n97 0.836707
R831 VTAIL.n97 VTAIL.n95 0.836707
R832 VTAIL.n391 VTAIL.n389 0.836707
R833 VTAIL VTAIL.n1 0.685845
R834 VTAIL.n328 VTAIL.n327 0.388379
R835 VTAIL.n373 VTAIL.n372 0.388379
R836 VTAIL.n374 VTAIL.n302 0.388379
R837 VTAIL.n34 VTAIL.n33 0.388379
R838 VTAIL.n79 VTAIL.n78 0.388379
R839 VTAIL.n80 VTAIL.n8 0.388379
R840 VTAIL.n280 VTAIL.n208 0.388379
R841 VTAIL.n279 VTAIL.n278 0.388379
R842 VTAIL.n235 VTAIL.n234 0.388379
R843 VTAIL.n182 VTAIL.n110 0.388379
R844 VTAIL.n181 VTAIL.n180 0.388379
R845 VTAIL.n137 VTAIL.n136 0.388379
R846 VTAIL.n330 VTAIL.n329 0.155672
R847 VTAIL.n330 VTAIL.n321 0.155672
R848 VTAIL.n337 VTAIL.n321 0.155672
R849 VTAIL.n338 VTAIL.n337 0.155672
R850 VTAIL.n338 VTAIL.n317 0.155672
R851 VTAIL.n345 VTAIL.n317 0.155672
R852 VTAIL.n346 VTAIL.n345 0.155672
R853 VTAIL.n346 VTAIL.n313 0.155672
R854 VTAIL.n353 VTAIL.n313 0.155672
R855 VTAIL.n354 VTAIL.n353 0.155672
R856 VTAIL.n354 VTAIL.n309 0.155672
R857 VTAIL.n361 VTAIL.n309 0.155672
R858 VTAIL.n362 VTAIL.n361 0.155672
R859 VTAIL.n362 VTAIL.n305 0.155672
R860 VTAIL.n370 VTAIL.n305 0.155672
R861 VTAIL.n371 VTAIL.n370 0.155672
R862 VTAIL.n371 VTAIL.n301 0.155672
R863 VTAIL.n379 VTAIL.n301 0.155672
R864 VTAIL.n380 VTAIL.n379 0.155672
R865 VTAIL.n380 VTAIL.n297 0.155672
R866 VTAIL.n387 VTAIL.n297 0.155672
R867 VTAIL.n36 VTAIL.n35 0.155672
R868 VTAIL.n36 VTAIL.n27 0.155672
R869 VTAIL.n43 VTAIL.n27 0.155672
R870 VTAIL.n44 VTAIL.n43 0.155672
R871 VTAIL.n44 VTAIL.n23 0.155672
R872 VTAIL.n51 VTAIL.n23 0.155672
R873 VTAIL.n52 VTAIL.n51 0.155672
R874 VTAIL.n52 VTAIL.n19 0.155672
R875 VTAIL.n59 VTAIL.n19 0.155672
R876 VTAIL.n60 VTAIL.n59 0.155672
R877 VTAIL.n60 VTAIL.n15 0.155672
R878 VTAIL.n67 VTAIL.n15 0.155672
R879 VTAIL.n68 VTAIL.n67 0.155672
R880 VTAIL.n68 VTAIL.n11 0.155672
R881 VTAIL.n76 VTAIL.n11 0.155672
R882 VTAIL.n77 VTAIL.n76 0.155672
R883 VTAIL.n77 VTAIL.n7 0.155672
R884 VTAIL.n85 VTAIL.n7 0.155672
R885 VTAIL.n86 VTAIL.n85 0.155672
R886 VTAIL.n86 VTAIL.n3 0.155672
R887 VTAIL.n93 VTAIL.n3 0.155672
R888 VTAIL.n293 VTAIL.n203 0.155672
R889 VTAIL.n286 VTAIL.n203 0.155672
R890 VTAIL.n286 VTAIL.n285 0.155672
R891 VTAIL.n285 VTAIL.n207 0.155672
R892 VTAIL.n277 VTAIL.n207 0.155672
R893 VTAIL.n277 VTAIL.n276 0.155672
R894 VTAIL.n276 VTAIL.n211 0.155672
R895 VTAIL.n269 VTAIL.n211 0.155672
R896 VTAIL.n269 VTAIL.n268 0.155672
R897 VTAIL.n268 VTAIL.n216 0.155672
R898 VTAIL.n261 VTAIL.n216 0.155672
R899 VTAIL.n261 VTAIL.n260 0.155672
R900 VTAIL.n260 VTAIL.n220 0.155672
R901 VTAIL.n253 VTAIL.n220 0.155672
R902 VTAIL.n253 VTAIL.n252 0.155672
R903 VTAIL.n252 VTAIL.n224 0.155672
R904 VTAIL.n245 VTAIL.n224 0.155672
R905 VTAIL.n245 VTAIL.n244 0.155672
R906 VTAIL.n244 VTAIL.n228 0.155672
R907 VTAIL.n237 VTAIL.n228 0.155672
R908 VTAIL.n237 VTAIL.n236 0.155672
R909 VTAIL.n195 VTAIL.n105 0.155672
R910 VTAIL.n188 VTAIL.n105 0.155672
R911 VTAIL.n188 VTAIL.n187 0.155672
R912 VTAIL.n187 VTAIL.n109 0.155672
R913 VTAIL.n179 VTAIL.n109 0.155672
R914 VTAIL.n179 VTAIL.n178 0.155672
R915 VTAIL.n178 VTAIL.n113 0.155672
R916 VTAIL.n171 VTAIL.n113 0.155672
R917 VTAIL.n171 VTAIL.n170 0.155672
R918 VTAIL.n170 VTAIL.n118 0.155672
R919 VTAIL.n163 VTAIL.n118 0.155672
R920 VTAIL.n163 VTAIL.n162 0.155672
R921 VTAIL.n162 VTAIL.n122 0.155672
R922 VTAIL.n155 VTAIL.n122 0.155672
R923 VTAIL.n155 VTAIL.n154 0.155672
R924 VTAIL.n154 VTAIL.n126 0.155672
R925 VTAIL.n147 VTAIL.n126 0.155672
R926 VTAIL.n147 VTAIL.n146 0.155672
R927 VTAIL.n146 VTAIL.n130 0.155672
R928 VTAIL.n139 VTAIL.n130 0.155672
R929 VTAIL.n139 VTAIL.n138 0.155672
R930 VTAIL VTAIL.n391 0.151362
R931 B.n466 B.t17 837.15
R932 B.n464 B.t21 837.15
R933 B.n112 B.t14 837.15
R934 B.n110 B.t10 837.15
R935 B.n819 B.n818 585
R936 B.n820 B.n819 585
R937 B.n354 B.n109 585
R938 B.n353 B.n352 585
R939 B.n351 B.n350 585
R940 B.n349 B.n348 585
R941 B.n347 B.n346 585
R942 B.n345 B.n344 585
R943 B.n343 B.n342 585
R944 B.n341 B.n340 585
R945 B.n339 B.n338 585
R946 B.n337 B.n336 585
R947 B.n335 B.n334 585
R948 B.n333 B.n332 585
R949 B.n331 B.n330 585
R950 B.n329 B.n328 585
R951 B.n327 B.n326 585
R952 B.n325 B.n324 585
R953 B.n323 B.n322 585
R954 B.n321 B.n320 585
R955 B.n319 B.n318 585
R956 B.n317 B.n316 585
R957 B.n315 B.n314 585
R958 B.n313 B.n312 585
R959 B.n311 B.n310 585
R960 B.n309 B.n308 585
R961 B.n307 B.n306 585
R962 B.n305 B.n304 585
R963 B.n303 B.n302 585
R964 B.n301 B.n300 585
R965 B.n299 B.n298 585
R966 B.n297 B.n296 585
R967 B.n295 B.n294 585
R968 B.n293 B.n292 585
R969 B.n291 B.n290 585
R970 B.n289 B.n288 585
R971 B.n287 B.n286 585
R972 B.n285 B.n284 585
R973 B.n283 B.n282 585
R974 B.n281 B.n280 585
R975 B.n279 B.n278 585
R976 B.n277 B.n276 585
R977 B.n275 B.n274 585
R978 B.n273 B.n272 585
R979 B.n271 B.n270 585
R980 B.n269 B.n268 585
R981 B.n267 B.n266 585
R982 B.n265 B.n264 585
R983 B.n263 B.n262 585
R984 B.n261 B.n260 585
R985 B.n259 B.n258 585
R986 B.n257 B.n256 585
R987 B.n255 B.n254 585
R988 B.n253 B.n252 585
R989 B.n251 B.n250 585
R990 B.n249 B.n248 585
R991 B.n247 B.n246 585
R992 B.n244 B.n243 585
R993 B.n242 B.n241 585
R994 B.n240 B.n239 585
R995 B.n238 B.n237 585
R996 B.n236 B.n235 585
R997 B.n234 B.n233 585
R998 B.n232 B.n231 585
R999 B.n230 B.n229 585
R1000 B.n228 B.n227 585
R1001 B.n226 B.n225 585
R1002 B.n224 B.n223 585
R1003 B.n222 B.n221 585
R1004 B.n220 B.n219 585
R1005 B.n218 B.n217 585
R1006 B.n216 B.n215 585
R1007 B.n214 B.n213 585
R1008 B.n212 B.n211 585
R1009 B.n210 B.n209 585
R1010 B.n208 B.n207 585
R1011 B.n206 B.n205 585
R1012 B.n204 B.n203 585
R1013 B.n202 B.n201 585
R1014 B.n200 B.n199 585
R1015 B.n198 B.n197 585
R1016 B.n196 B.n195 585
R1017 B.n194 B.n193 585
R1018 B.n192 B.n191 585
R1019 B.n190 B.n189 585
R1020 B.n188 B.n187 585
R1021 B.n186 B.n185 585
R1022 B.n184 B.n183 585
R1023 B.n182 B.n181 585
R1024 B.n180 B.n179 585
R1025 B.n178 B.n177 585
R1026 B.n176 B.n175 585
R1027 B.n174 B.n173 585
R1028 B.n172 B.n171 585
R1029 B.n170 B.n169 585
R1030 B.n168 B.n167 585
R1031 B.n166 B.n165 585
R1032 B.n164 B.n163 585
R1033 B.n162 B.n161 585
R1034 B.n160 B.n159 585
R1035 B.n158 B.n157 585
R1036 B.n156 B.n155 585
R1037 B.n154 B.n153 585
R1038 B.n152 B.n151 585
R1039 B.n150 B.n149 585
R1040 B.n148 B.n147 585
R1041 B.n146 B.n145 585
R1042 B.n144 B.n143 585
R1043 B.n142 B.n141 585
R1044 B.n140 B.n139 585
R1045 B.n138 B.n137 585
R1046 B.n136 B.n135 585
R1047 B.n134 B.n133 585
R1048 B.n132 B.n131 585
R1049 B.n130 B.n129 585
R1050 B.n128 B.n127 585
R1051 B.n126 B.n125 585
R1052 B.n124 B.n123 585
R1053 B.n122 B.n121 585
R1054 B.n120 B.n119 585
R1055 B.n118 B.n117 585
R1056 B.n116 B.n115 585
R1057 B.n817 B.n48 585
R1058 B.n821 B.n48 585
R1059 B.n816 B.n47 585
R1060 B.n822 B.n47 585
R1061 B.n815 B.n814 585
R1062 B.n814 B.n43 585
R1063 B.n813 B.n42 585
R1064 B.n828 B.n42 585
R1065 B.n812 B.n41 585
R1066 B.n829 B.n41 585
R1067 B.n811 B.n40 585
R1068 B.n830 B.n40 585
R1069 B.n810 B.n809 585
R1070 B.n809 B.n36 585
R1071 B.n808 B.n35 585
R1072 B.n836 B.n35 585
R1073 B.n807 B.n34 585
R1074 B.n837 B.n34 585
R1075 B.n806 B.n33 585
R1076 B.n838 B.n33 585
R1077 B.n805 B.n804 585
R1078 B.n804 B.n32 585
R1079 B.n803 B.n28 585
R1080 B.n844 B.n28 585
R1081 B.n802 B.n27 585
R1082 B.n845 B.n27 585
R1083 B.n801 B.n26 585
R1084 B.n846 B.n26 585
R1085 B.n800 B.n799 585
R1086 B.n799 B.n22 585
R1087 B.n798 B.n21 585
R1088 B.n852 B.n21 585
R1089 B.n797 B.n20 585
R1090 B.n853 B.n20 585
R1091 B.n796 B.n19 585
R1092 B.n854 B.n19 585
R1093 B.n795 B.n794 585
R1094 B.n794 B.n15 585
R1095 B.n793 B.n14 585
R1096 B.n860 B.n14 585
R1097 B.n792 B.n13 585
R1098 B.n861 B.n13 585
R1099 B.n791 B.n12 585
R1100 B.n862 B.n12 585
R1101 B.n790 B.n789 585
R1102 B.n789 B.n8 585
R1103 B.n788 B.n7 585
R1104 B.n868 B.n7 585
R1105 B.n787 B.n6 585
R1106 B.n869 B.n6 585
R1107 B.n786 B.n5 585
R1108 B.n870 B.n5 585
R1109 B.n785 B.n784 585
R1110 B.n784 B.n4 585
R1111 B.n783 B.n355 585
R1112 B.n783 B.n782 585
R1113 B.n773 B.n356 585
R1114 B.n357 B.n356 585
R1115 B.n775 B.n774 585
R1116 B.n776 B.n775 585
R1117 B.n772 B.n362 585
R1118 B.n362 B.n361 585
R1119 B.n771 B.n770 585
R1120 B.n770 B.n769 585
R1121 B.n364 B.n363 585
R1122 B.n365 B.n364 585
R1123 B.n762 B.n761 585
R1124 B.n763 B.n762 585
R1125 B.n760 B.n369 585
R1126 B.n373 B.n369 585
R1127 B.n759 B.n758 585
R1128 B.n758 B.n757 585
R1129 B.n371 B.n370 585
R1130 B.n372 B.n371 585
R1131 B.n750 B.n749 585
R1132 B.n751 B.n750 585
R1133 B.n748 B.n378 585
R1134 B.n378 B.n377 585
R1135 B.n747 B.n746 585
R1136 B.n746 B.n745 585
R1137 B.n380 B.n379 585
R1138 B.n738 B.n380 585
R1139 B.n737 B.n736 585
R1140 B.n739 B.n737 585
R1141 B.n735 B.n385 585
R1142 B.n385 B.n384 585
R1143 B.n734 B.n733 585
R1144 B.n733 B.n732 585
R1145 B.n387 B.n386 585
R1146 B.n388 B.n387 585
R1147 B.n725 B.n724 585
R1148 B.n726 B.n725 585
R1149 B.n723 B.n392 585
R1150 B.n396 B.n392 585
R1151 B.n722 B.n721 585
R1152 B.n721 B.n720 585
R1153 B.n394 B.n393 585
R1154 B.n395 B.n394 585
R1155 B.n713 B.n712 585
R1156 B.n714 B.n713 585
R1157 B.n711 B.n401 585
R1158 B.n401 B.n400 585
R1159 B.n705 B.n704 585
R1160 B.n703 B.n463 585
R1161 B.n702 B.n462 585
R1162 B.n707 B.n462 585
R1163 B.n701 B.n700 585
R1164 B.n699 B.n698 585
R1165 B.n697 B.n696 585
R1166 B.n695 B.n694 585
R1167 B.n693 B.n692 585
R1168 B.n691 B.n690 585
R1169 B.n689 B.n688 585
R1170 B.n687 B.n686 585
R1171 B.n685 B.n684 585
R1172 B.n683 B.n682 585
R1173 B.n681 B.n680 585
R1174 B.n679 B.n678 585
R1175 B.n677 B.n676 585
R1176 B.n675 B.n674 585
R1177 B.n673 B.n672 585
R1178 B.n671 B.n670 585
R1179 B.n669 B.n668 585
R1180 B.n667 B.n666 585
R1181 B.n665 B.n664 585
R1182 B.n663 B.n662 585
R1183 B.n661 B.n660 585
R1184 B.n659 B.n658 585
R1185 B.n657 B.n656 585
R1186 B.n655 B.n654 585
R1187 B.n653 B.n652 585
R1188 B.n651 B.n650 585
R1189 B.n649 B.n648 585
R1190 B.n647 B.n646 585
R1191 B.n645 B.n644 585
R1192 B.n643 B.n642 585
R1193 B.n641 B.n640 585
R1194 B.n639 B.n638 585
R1195 B.n637 B.n636 585
R1196 B.n635 B.n634 585
R1197 B.n633 B.n632 585
R1198 B.n631 B.n630 585
R1199 B.n629 B.n628 585
R1200 B.n627 B.n626 585
R1201 B.n625 B.n624 585
R1202 B.n623 B.n622 585
R1203 B.n621 B.n620 585
R1204 B.n619 B.n618 585
R1205 B.n617 B.n616 585
R1206 B.n615 B.n614 585
R1207 B.n613 B.n612 585
R1208 B.n611 B.n610 585
R1209 B.n609 B.n608 585
R1210 B.n607 B.n606 585
R1211 B.n605 B.n604 585
R1212 B.n603 B.n602 585
R1213 B.n601 B.n600 585
R1214 B.n599 B.n598 585
R1215 B.n597 B.n596 585
R1216 B.n594 B.n593 585
R1217 B.n592 B.n591 585
R1218 B.n590 B.n589 585
R1219 B.n588 B.n587 585
R1220 B.n586 B.n585 585
R1221 B.n584 B.n583 585
R1222 B.n582 B.n581 585
R1223 B.n580 B.n579 585
R1224 B.n578 B.n577 585
R1225 B.n576 B.n575 585
R1226 B.n574 B.n573 585
R1227 B.n572 B.n571 585
R1228 B.n570 B.n569 585
R1229 B.n568 B.n567 585
R1230 B.n566 B.n565 585
R1231 B.n564 B.n563 585
R1232 B.n562 B.n561 585
R1233 B.n560 B.n559 585
R1234 B.n558 B.n557 585
R1235 B.n556 B.n555 585
R1236 B.n554 B.n553 585
R1237 B.n552 B.n551 585
R1238 B.n550 B.n549 585
R1239 B.n548 B.n547 585
R1240 B.n546 B.n545 585
R1241 B.n544 B.n543 585
R1242 B.n542 B.n541 585
R1243 B.n540 B.n539 585
R1244 B.n538 B.n537 585
R1245 B.n536 B.n535 585
R1246 B.n534 B.n533 585
R1247 B.n532 B.n531 585
R1248 B.n530 B.n529 585
R1249 B.n528 B.n527 585
R1250 B.n526 B.n525 585
R1251 B.n524 B.n523 585
R1252 B.n522 B.n521 585
R1253 B.n520 B.n519 585
R1254 B.n518 B.n517 585
R1255 B.n516 B.n515 585
R1256 B.n514 B.n513 585
R1257 B.n512 B.n511 585
R1258 B.n510 B.n509 585
R1259 B.n508 B.n507 585
R1260 B.n506 B.n505 585
R1261 B.n504 B.n503 585
R1262 B.n502 B.n501 585
R1263 B.n500 B.n499 585
R1264 B.n498 B.n497 585
R1265 B.n496 B.n495 585
R1266 B.n494 B.n493 585
R1267 B.n492 B.n491 585
R1268 B.n490 B.n489 585
R1269 B.n488 B.n487 585
R1270 B.n486 B.n485 585
R1271 B.n484 B.n483 585
R1272 B.n482 B.n481 585
R1273 B.n480 B.n479 585
R1274 B.n478 B.n477 585
R1275 B.n476 B.n475 585
R1276 B.n474 B.n473 585
R1277 B.n472 B.n471 585
R1278 B.n470 B.n469 585
R1279 B.n403 B.n402 585
R1280 B.n710 B.n709 585
R1281 B.n399 B.n398 585
R1282 B.n400 B.n399 585
R1283 B.n716 B.n715 585
R1284 B.n715 B.n714 585
R1285 B.n717 B.n397 585
R1286 B.n397 B.n395 585
R1287 B.n719 B.n718 585
R1288 B.n720 B.n719 585
R1289 B.n391 B.n390 585
R1290 B.n396 B.n391 585
R1291 B.n728 B.n727 585
R1292 B.n727 B.n726 585
R1293 B.n729 B.n389 585
R1294 B.n389 B.n388 585
R1295 B.n731 B.n730 585
R1296 B.n732 B.n731 585
R1297 B.n383 B.n382 585
R1298 B.n384 B.n383 585
R1299 B.n741 B.n740 585
R1300 B.n740 B.n739 585
R1301 B.n742 B.n381 585
R1302 B.n738 B.n381 585
R1303 B.n744 B.n743 585
R1304 B.n745 B.n744 585
R1305 B.n376 B.n375 585
R1306 B.n377 B.n376 585
R1307 B.n753 B.n752 585
R1308 B.n752 B.n751 585
R1309 B.n754 B.n374 585
R1310 B.n374 B.n372 585
R1311 B.n756 B.n755 585
R1312 B.n757 B.n756 585
R1313 B.n368 B.n367 585
R1314 B.n373 B.n368 585
R1315 B.n765 B.n764 585
R1316 B.n764 B.n763 585
R1317 B.n766 B.n366 585
R1318 B.n366 B.n365 585
R1319 B.n768 B.n767 585
R1320 B.n769 B.n768 585
R1321 B.n360 B.n359 585
R1322 B.n361 B.n360 585
R1323 B.n778 B.n777 585
R1324 B.n777 B.n776 585
R1325 B.n779 B.n358 585
R1326 B.n358 B.n357 585
R1327 B.n781 B.n780 585
R1328 B.n782 B.n781 585
R1329 B.n2 B.n0 585
R1330 B.n4 B.n2 585
R1331 B.n3 B.n1 585
R1332 B.n869 B.n3 585
R1333 B.n867 B.n866 585
R1334 B.n868 B.n867 585
R1335 B.n865 B.n9 585
R1336 B.n9 B.n8 585
R1337 B.n864 B.n863 585
R1338 B.n863 B.n862 585
R1339 B.n11 B.n10 585
R1340 B.n861 B.n11 585
R1341 B.n859 B.n858 585
R1342 B.n860 B.n859 585
R1343 B.n857 B.n16 585
R1344 B.n16 B.n15 585
R1345 B.n856 B.n855 585
R1346 B.n855 B.n854 585
R1347 B.n18 B.n17 585
R1348 B.n853 B.n18 585
R1349 B.n851 B.n850 585
R1350 B.n852 B.n851 585
R1351 B.n849 B.n23 585
R1352 B.n23 B.n22 585
R1353 B.n848 B.n847 585
R1354 B.n847 B.n846 585
R1355 B.n25 B.n24 585
R1356 B.n845 B.n25 585
R1357 B.n843 B.n842 585
R1358 B.n844 B.n843 585
R1359 B.n841 B.n29 585
R1360 B.n32 B.n29 585
R1361 B.n840 B.n839 585
R1362 B.n839 B.n838 585
R1363 B.n31 B.n30 585
R1364 B.n837 B.n31 585
R1365 B.n835 B.n834 585
R1366 B.n836 B.n835 585
R1367 B.n833 B.n37 585
R1368 B.n37 B.n36 585
R1369 B.n832 B.n831 585
R1370 B.n831 B.n830 585
R1371 B.n39 B.n38 585
R1372 B.n829 B.n39 585
R1373 B.n827 B.n826 585
R1374 B.n828 B.n827 585
R1375 B.n825 B.n44 585
R1376 B.n44 B.n43 585
R1377 B.n824 B.n823 585
R1378 B.n823 B.n822 585
R1379 B.n46 B.n45 585
R1380 B.n821 B.n46 585
R1381 B.n872 B.n871 585
R1382 B.n871 B.n870 585
R1383 B.n705 B.n399 550.159
R1384 B.n115 B.n46 550.159
R1385 B.n709 B.n401 550.159
R1386 B.n819 B.n48 550.159
R1387 B.n466 B.t20 383.971
R1388 B.n110 B.t12 383.971
R1389 B.n464 B.t23 383.971
R1390 B.n112 B.t15 383.971
R1391 B.n467 B.t19 365.159
R1392 B.n111 B.t13 365.159
R1393 B.n465 B.t22 365.159
R1394 B.n113 B.t16 365.159
R1395 B.n820 B.n108 256.663
R1396 B.n820 B.n107 256.663
R1397 B.n820 B.n106 256.663
R1398 B.n820 B.n105 256.663
R1399 B.n820 B.n104 256.663
R1400 B.n820 B.n103 256.663
R1401 B.n820 B.n102 256.663
R1402 B.n820 B.n101 256.663
R1403 B.n820 B.n100 256.663
R1404 B.n820 B.n99 256.663
R1405 B.n820 B.n98 256.663
R1406 B.n820 B.n97 256.663
R1407 B.n820 B.n96 256.663
R1408 B.n820 B.n95 256.663
R1409 B.n820 B.n94 256.663
R1410 B.n820 B.n93 256.663
R1411 B.n820 B.n92 256.663
R1412 B.n820 B.n91 256.663
R1413 B.n820 B.n90 256.663
R1414 B.n820 B.n89 256.663
R1415 B.n820 B.n88 256.663
R1416 B.n820 B.n87 256.663
R1417 B.n820 B.n86 256.663
R1418 B.n820 B.n85 256.663
R1419 B.n820 B.n84 256.663
R1420 B.n820 B.n83 256.663
R1421 B.n820 B.n82 256.663
R1422 B.n820 B.n81 256.663
R1423 B.n820 B.n80 256.663
R1424 B.n820 B.n79 256.663
R1425 B.n820 B.n78 256.663
R1426 B.n820 B.n77 256.663
R1427 B.n820 B.n76 256.663
R1428 B.n820 B.n75 256.663
R1429 B.n820 B.n74 256.663
R1430 B.n820 B.n73 256.663
R1431 B.n820 B.n72 256.663
R1432 B.n820 B.n71 256.663
R1433 B.n820 B.n70 256.663
R1434 B.n820 B.n69 256.663
R1435 B.n820 B.n68 256.663
R1436 B.n820 B.n67 256.663
R1437 B.n820 B.n66 256.663
R1438 B.n820 B.n65 256.663
R1439 B.n820 B.n64 256.663
R1440 B.n820 B.n63 256.663
R1441 B.n820 B.n62 256.663
R1442 B.n820 B.n61 256.663
R1443 B.n820 B.n60 256.663
R1444 B.n820 B.n59 256.663
R1445 B.n820 B.n58 256.663
R1446 B.n820 B.n57 256.663
R1447 B.n820 B.n56 256.663
R1448 B.n820 B.n55 256.663
R1449 B.n820 B.n54 256.663
R1450 B.n820 B.n53 256.663
R1451 B.n820 B.n52 256.663
R1452 B.n820 B.n51 256.663
R1453 B.n820 B.n50 256.663
R1454 B.n820 B.n49 256.663
R1455 B.n707 B.n706 256.663
R1456 B.n707 B.n404 256.663
R1457 B.n707 B.n405 256.663
R1458 B.n707 B.n406 256.663
R1459 B.n707 B.n407 256.663
R1460 B.n707 B.n408 256.663
R1461 B.n707 B.n409 256.663
R1462 B.n707 B.n410 256.663
R1463 B.n707 B.n411 256.663
R1464 B.n707 B.n412 256.663
R1465 B.n707 B.n413 256.663
R1466 B.n707 B.n414 256.663
R1467 B.n707 B.n415 256.663
R1468 B.n707 B.n416 256.663
R1469 B.n707 B.n417 256.663
R1470 B.n707 B.n418 256.663
R1471 B.n707 B.n419 256.663
R1472 B.n707 B.n420 256.663
R1473 B.n707 B.n421 256.663
R1474 B.n707 B.n422 256.663
R1475 B.n707 B.n423 256.663
R1476 B.n707 B.n424 256.663
R1477 B.n707 B.n425 256.663
R1478 B.n707 B.n426 256.663
R1479 B.n707 B.n427 256.663
R1480 B.n707 B.n428 256.663
R1481 B.n707 B.n429 256.663
R1482 B.n707 B.n430 256.663
R1483 B.n707 B.n431 256.663
R1484 B.n707 B.n432 256.663
R1485 B.n707 B.n433 256.663
R1486 B.n707 B.n434 256.663
R1487 B.n707 B.n435 256.663
R1488 B.n707 B.n436 256.663
R1489 B.n707 B.n437 256.663
R1490 B.n707 B.n438 256.663
R1491 B.n707 B.n439 256.663
R1492 B.n707 B.n440 256.663
R1493 B.n707 B.n441 256.663
R1494 B.n707 B.n442 256.663
R1495 B.n707 B.n443 256.663
R1496 B.n707 B.n444 256.663
R1497 B.n707 B.n445 256.663
R1498 B.n707 B.n446 256.663
R1499 B.n707 B.n447 256.663
R1500 B.n707 B.n448 256.663
R1501 B.n707 B.n449 256.663
R1502 B.n707 B.n450 256.663
R1503 B.n707 B.n451 256.663
R1504 B.n707 B.n452 256.663
R1505 B.n707 B.n453 256.663
R1506 B.n707 B.n454 256.663
R1507 B.n707 B.n455 256.663
R1508 B.n707 B.n456 256.663
R1509 B.n707 B.n457 256.663
R1510 B.n707 B.n458 256.663
R1511 B.n707 B.n459 256.663
R1512 B.n707 B.n460 256.663
R1513 B.n707 B.n461 256.663
R1514 B.n708 B.n707 256.663
R1515 B.n715 B.n399 163.367
R1516 B.n715 B.n397 163.367
R1517 B.n719 B.n397 163.367
R1518 B.n719 B.n391 163.367
R1519 B.n727 B.n391 163.367
R1520 B.n727 B.n389 163.367
R1521 B.n731 B.n389 163.367
R1522 B.n731 B.n383 163.367
R1523 B.n740 B.n383 163.367
R1524 B.n740 B.n381 163.367
R1525 B.n744 B.n381 163.367
R1526 B.n744 B.n376 163.367
R1527 B.n752 B.n376 163.367
R1528 B.n752 B.n374 163.367
R1529 B.n756 B.n374 163.367
R1530 B.n756 B.n368 163.367
R1531 B.n764 B.n368 163.367
R1532 B.n764 B.n366 163.367
R1533 B.n768 B.n366 163.367
R1534 B.n768 B.n360 163.367
R1535 B.n777 B.n360 163.367
R1536 B.n777 B.n358 163.367
R1537 B.n781 B.n358 163.367
R1538 B.n781 B.n2 163.367
R1539 B.n871 B.n2 163.367
R1540 B.n871 B.n3 163.367
R1541 B.n867 B.n3 163.367
R1542 B.n867 B.n9 163.367
R1543 B.n863 B.n9 163.367
R1544 B.n863 B.n11 163.367
R1545 B.n859 B.n11 163.367
R1546 B.n859 B.n16 163.367
R1547 B.n855 B.n16 163.367
R1548 B.n855 B.n18 163.367
R1549 B.n851 B.n18 163.367
R1550 B.n851 B.n23 163.367
R1551 B.n847 B.n23 163.367
R1552 B.n847 B.n25 163.367
R1553 B.n843 B.n25 163.367
R1554 B.n843 B.n29 163.367
R1555 B.n839 B.n29 163.367
R1556 B.n839 B.n31 163.367
R1557 B.n835 B.n31 163.367
R1558 B.n835 B.n37 163.367
R1559 B.n831 B.n37 163.367
R1560 B.n831 B.n39 163.367
R1561 B.n827 B.n39 163.367
R1562 B.n827 B.n44 163.367
R1563 B.n823 B.n44 163.367
R1564 B.n823 B.n46 163.367
R1565 B.n463 B.n462 163.367
R1566 B.n700 B.n462 163.367
R1567 B.n698 B.n697 163.367
R1568 B.n694 B.n693 163.367
R1569 B.n690 B.n689 163.367
R1570 B.n686 B.n685 163.367
R1571 B.n682 B.n681 163.367
R1572 B.n678 B.n677 163.367
R1573 B.n674 B.n673 163.367
R1574 B.n670 B.n669 163.367
R1575 B.n666 B.n665 163.367
R1576 B.n662 B.n661 163.367
R1577 B.n658 B.n657 163.367
R1578 B.n654 B.n653 163.367
R1579 B.n650 B.n649 163.367
R1580 B.n646 B.n645 163.367
R1581 B.n642 B.n641 163.367
R1582 B.n638 B.n637 163.367
R1583 B.n634 B.n633 163.367
R1584 B.n630 B.n629 163.367
R1585 B.n626 B.n625 163.367
R1586 B.n622 B.n621 163.367
R1587 B.n618 B.n617 163.367
R1588 B.n614 B.n613 163.367
R1589 B.n610 B.n609 163.367
R1590 B.n606 B.n605 163.367
R1591 B.n602 B.n601 163.367
R1592 B.n598 B.n597 163.367
R1593 B.n593 B.n592 163.367
R1594 B.n589 B.n588 163.367
R1595 B.n585 B.n584 163.367
R1596 B.n581 B.n580 163.367
R1597 B.n577 B.n576 163.367
R1598 B.n573 B.n572 163.367
R1599 B.n569 B.n568 163.367
R1600 B.n565 B.n564 163.367
R1601 B.n561 B.n560 163.367
R1602 B.n557 B.n556 163.367
R1603 B.n553 B.n552 163.367
R1604 B.n549 B.n548 163.367
R1605 B.n545 B.n544 163.367
R1606 B.n541 B.n540 163.367
R1607 B.n537 B.n536 163.367
R1608 B.n533 B.n532 163.367
R1609 B.n529 B.n528 163.367
R1610 B.n525 B.n524 163.367
R1611 B.n521 B.n520 163.367
R1612 B.n517 B.n516 163.367
R1613 B.n513 B.n512 163.367
R1614 B.n509 B.n508 163.367
R1615 B.n505 B.n504 163.367
R1616 B.n501 B.n500 163.367
R1617 B.n497 B.n496 163.367
R1618 B.n493 B.n492 163.367
R1619 B.n489 B.n488 163.367
R1620 B.n485 B.n484 163.367
R1621 B.n481 B.n480 163.367
R1622 B.n477 B.n476 163.367
R1623 B.n473 B.n472 163.367
R1624 B.n469 B.n403 163.367
R1625 B.n713 B.n401 163.367
R1626 B.n713 B.n394 163.367
R1627 B.n721 B.n394 163.367
R1628 B.n721 B.n392 163.367
R1629 B.n725 B.n392 163.367
R1630 B.n725 B.n387 163.367
R1631 B.n733 B.n387 163.367
R1632 B.n733 B.n385 163.367
R1633 B.n737 B.n385 163.367
R1634 B.n737 B.n380 163.367
R1635 B.n746 B.n380 163.367
R1636 B.n746 B.n378 163.367
R1637 B.n750 B.n378 163.367
R1638 B.n750 B.n371 163.367
R1639 B.n758 B.n371 163.367
R1640 B.n758 B.n369 163.367
R1641 B.n762 B.n369 163.367
R1642 B.n762 B.n364 163.367
R1643 B.n770 B.n364 163.367
R1644 B.n770 B.n362 163.367
R1645 B.n775 B.n362 163.367
R1646 B.n775 B.n356 163.367
R1647 B.n783 B.n356 163.367
R1648 B.n784 B.n783 163.367
R1649 B.n784 B.n5 163.367
R1650 B.n6 B.n5 163.367
R1651 B.n7 B.n6 163.367
R1652 B.n789 B.n7 163.367
R1653 B.n789 B.n12 163.367
R1654 B.n13 B.n12 163.367
R1655 B.n14 B.n13 163.367
R1656 B.n794 B.n14 163.367
R1657 B.n794 B.n19 163.367
R1658 B.n20 B.n19 163.367
R1659 B.n21 B.n20 163.367
R1660 B.n799 B.n21 163.367
R1661 B.n799 B.n26 163.367
R1662 B.n27 B.n26 163.367
R1663 B.n28 B.n27 163.367
R1664 B.n804 B.n28 163.367
R1665 B.n804 B.n33 163.367
R1666 B.n34 B.n33 163.367
R1667 B.n35 B.n34 163.367
R1668 B.n809 B.n35 163.367
R1669 B.n809 B.n40 163.367
R1670 B.n41 B.n40 163.367
R1671 B.n42 B.n41 163.367
R1672 B.n814 B.n42 163.367
R1673 B.n814 B.n47 163.367
R1674 B.n48 B.n47 163.367
R1675 B.n119 B.n118 163.367
R1676 B.n123 B.n122 163.367
R1677 B.n127 B.n126 163.367
R1678 B.n131 B.n130 163.367
R1679 B.n135 B.n134 163.367
R1680 B.n139 B.n138 163.367
R1681 B.n143 B.n142 163.367
R1682 B.n147 B.n146 163.367
R1683 B.n151 B.n150 163.367
R1684 B.n155 B.n154 163.367
R1685 B.n159 B.n158 163.367
R1686 B.n163 B.n162 163.367
R1687 B.n167 B.n166 163.367
R1688 B.n171 B.n170 163.367
R1689 B.n175 B.n174 163.367
R1690 B.n179 B.n178 163.367
R1691 B.n183 B.n182 163.367
R1692 B.n187 B.n186 163.367
R1693 B.n191 B.n190 163.367
R1694 B.n195 B.n194 163.367
R1695 B.n199 B.n198 163.367
R1696 B.n203 B.n202 163.367
R1697 B.n207 B.n206 163.367
R1698 B.n211 B.n210 163.367
R1699 B.n215 B.n214 163.367
R1700 B.n219 B.n218 163.367
R1701 B.n223 B.n222 163.367
R1702 B.n227 B.n226 163.367
R1703 B.n231 B.n230 163.367
R1704 B.n235 B.n234 163.367
R1705 B.n239 B.n238 163.367
R1706 B.n243 B.n242 163.367
R1707 B.n248 B.n247 163.367
R1708 B.n252 B.n251 163.367
R1709 B.n256 B.n255 163.367
R1710 B.n260 B.n259 163.367
R1711 B.n264 B.n263 163.367
R1712 B.n268 B.n267 163.367
R1713 B.n272 B.n271 163.367
R1714 B.n276 B.n275 163.367
R1715 B.n280 B.n279 163.367
R1716 B.n284 B.n283 163.367
R1717 B.n288 B.n287 163.367
R1718 B.n292 B.n291 163.367
R1719 B.n296 B.n295 163.367
R1720 B.n300 B.n299 163.367
R1721 B.n304 B.n303 163.367
R1722 B.n308 B.n307 163.367
R1723 B.n312 B.n311 163.367
R1724 B.n316 B.n315 163.367
R1725 B.n320 B.n319 163.367
R1726 B.n324 B.n323 163.367
R1727 B.n328 B.n327 163.367
R1728 B.n332 B.n331 163.367
R1729 B.n336 B.n335 163.367
R1730 B.n340 B.n339 163.367
R1731 B.n344 B.n343 163.367
R1732 B.n348 B.n347 163.367
R1733 B.n352 B.n351 163.367
R1734 B.n819 B.n109 163.367
R1735 B.n706 B.n705 71.676
R1736 B.n700 B.n404 71.676
R1737 B.n697 B.n405 71.676
R1738 B.n693 B.n406 71.676
R1739 B.n689 B.n407 71.676
R1740 B.n685 B.n408 71.676
R1741 B.n681 B.n409 71.676
R1742 B.n677 B.n410 71.676
R1743 B.n673 B.n411 71.676
R1744 B.n669 B.n412 71.676
R1745 B.n665 B.n413 71.676
R1746 B.n661 B.n414 71.676
R1747 B.n657 B.n415 71.676
R1748 B.n653 B.n416 71.676
R1749 B.n649 B.n417 71.676
R1750 B.n645 B.n418 71.676
R1751 B.n641 B.n419 71.676
R1752 B.n637 B.n420 71.676
R1753 B.n633 B.n421 71.676
R1754 B.n629 B.n422 71.676
R1755 B.n625 B.n423 71.676
R1756 B.n621 B.n424 71.676
R1757 B.n617 B.n425 71.676
R1758 B.n613 B.n426 71.676
R1759 B.n609 B.n427 71.676
R1760 B.n605 B.n428 71.676
R1761 B.n601 B.n429 71.676
R1762 B.n597 B.n430 71.676
R1763 B.n592 B.n431 71.676
R1764 B.n588 B.n432 71.676
R1765 B.n584 B.n433 71.676
R1766 B.n580 B.n434 71.676
R1767 B.n576 B.n435 71.676
R1768 B.n572 B.n436 71.676
R1769 B.n568 B.n437 71.676
R1770 B.n564 B.n438 71.676
R1771 B.n560 B.n439 71.676
R1772 B.n556 B.n440 71.676
R1773 B.n552 B.n441 71.676
R1774 B.n548 B.n442 71.676
R1775 B.n544 B.n443 71.676
R1776 B.n540 B.n444 71.676
R1777 B.n536 B.n445 71.676
R1778 B.n532 B.n446 71.676
R1779 B.n528 B.n447 71.676
R1780 B.n524 B.n448 71.676
R1781 B.n520 B.n449 71.676
R1782 B.n516 B.n450 71.676
R1783 B.n512 B.n451 71.676
R1784 B.n508 B.n452 71.676
R1785 B.n504 B.n453 71.676
R1786 B.n500 B.n454 71.676
R1787 B.n496 B.n455 71.676
R1788 B.n492 B.n456 71.676
R1789 B.n488 B.n457 71.676
R1790 B.n484 B.n458 71.676
R1791 B.n480 B.n459 71.676
R1792 B.n476 B.n460 71.676
R1793 B.n472 B.n461 71.676
R1794 B.n708 B.n403 71.676
R1795 B.n115 B.n49 71.676
R1796 B.n119 B.n50 71.676
R1797 B.n123 B.n51 71.676
R1798 B.n127 B.n52 71.676
R1799 B.n131 B.n53 71.676
R1800 B.n135 B.n54 71.676
R1801 B.n139 B.n55 71.676
R1802 B.n143 B.n56 71.676
R1803 B.n147 B.n57 71.676
R1804 B.n151 B.n58 71.676
R1805 B.n155 B.n59 71.676
R1806 B.n159 B.n60 71.676
R1807 B.n163 B.n61 71.676
R1808 B.n167 B.n62 71.676
R1809 B.n171 B.n63 71.676
R1810 B.n175 B.n64 71.676
R1811 B.n179 B.n65 71.676
R1812 B.n183 B.n66 71.676
R1813 B.n187 B.n67 71.676
R1814 B.n191 B.n68 71.676
R1815 B.n195 B.n69 71.676
R1816 B.n199 B.n70 71.676
R1817 B.n203 B.n71 71.676
R1818 B.n207 B.n72 71.676
R1819 B.n211 B.n73 71.676
R1820 B.n215 B.n74 71.676
R1821 B.n219 B.n75 71.676
R1822 B.n223 B.n76 71.676
R1823 B.n227 B.n77 71.676
R1824 B.n231 B.n78 71.676
R1825 B.n235 B.n79 71.676
R1826 B.n239 B.n80 71.676
R1827 B.n243 B.n81 71.676
R1828 B.n248 B.n82 71.676
R1829 B.n252 B.n83 71.676
R1830 B.n256 B.n84 71.676
R1831 B.n260 B.n85 71.676
R1832 B.n264 B.n86 71.676
R1833 B.n268 B.n87 71.676
R1834 B.n272 B.n88 71.676
R1835 B.n276 B.n89 71.676
R1836 B.n280 B.n90 71.676
R1837 B.n284 B.n91 71.676
R1838 B.n288 B.n92 71.676
R1839 B.n292 B.n93 71.676
R1840 B.n296 B.n94 71.676
R1841 B.n300 B.n95 71.676
R1842 B.n304 B.n96 71.676
R1843 B.n308 B.n97 71.676
R1844 B.n312 B.n98 71.676
R1845 B.n316 B.n99 71.676
R1846 B.n320 B.n100 71.676
R1847 B.n324 B.n101 71.676
R1848 B.n328 B.n102 71.676
R1849 B.n332 B.n103 71.676
R1850 B.n336 B.n104 71.676
R1851 B.n340 B.n105 71.676
R1852 B.n344 B.n106 71.676
R1853 B.n348 B.n107 71.676
R1854 B.n352 B.n108 71.676
R1855 B.n109 B.n108 71.676
R1856 B.n351 B.n107 71.676
R1857 B.n347 B.n106 71.676
R1858 B.n343 B.n105 71.676
R1859 B.n339 B.n104 71.676
R1860 B.n335 B.n103 71.676
R1861 B.n331 B.n102 71.676
R1862 B.n327 B.n101 71.676
R1863 B.n323 B.n100 71.676
R1864 B.n319 B.n99 71.676
R1865 B.n315 B.n98 71.676
R1866 B.n311 B.n97 71.676
R1867 B.n307 B.n96 71.676
R1868 B.n303 B.n95 71.676
R1869 B.n299 B.n94 71.676
R1870 B.n295 B.n93 71.676
R1871 B.n291 B.n92 71.676
R1872 B.n287 B.n91 71.676
R1873 B.n283 B.n90 71.676
R1874 B.n279 B.n89 71.676
R1875 B.n275 B.n88 71.676
R1876 B.n271 B.n87 71.676
R1877 B.n267 B.n86 71.676
R1878 B.n263 B.n85 71.676
R1879 B.n259 B.n84 71.676
R1880 B.n255 B.n83 71.676
R1881 B.n251 B.n82 71.676
R1882 B.n247 B.n81 71.676
R1883 B.n242 B.n80 71.676
R1884 B.n238 B.n79 71.676
R1885 B.n234 B.n78 71.676
R1886 B.n230 B.n77 71.676
R1887 B.n226 B.n76 71.676
R1888 B.n222 B.n75 71.676
R1889 B.n218 B.n74 71.676
R1890 B.n214 B.n73 71.676
R1891 B.n210 B.n72 71.676
R1892 B.n206 B.n71 71.676
R1893 B.n202 B.n70 71.676
R1894 B.n198 B.n69 71.676
R1895 B.n194 B.n68 71.676
R1896 B.n190 B.n67 71.676
R1897 B.n186 B.n66 71.676
R1898 B.n182 B.n65 71.676
R1899 B.n178 B.n64 71.676
R1900 B.n174 B.n63 71.676
R1901 B.n170 B.n62 71.676
R1902 B.n166 B.n61 71.676
R1903 B.n162 B.n60 71.676
R1904 B.n158 B.n59 71.676
R1905 B.n154 B.n58 71.676
R1906 B.n150 B.n57 71.676
R1907 B.n146 B.n56 71.676
R1908 B.n142 B.n55 71.676
R1909 B.n138 B.n54 71.676
R1910 B.n134 B.n53 71.676
R1911 B.n130 B.n52 71.676
R1912 B.n126 B.n51 71.676
R1913 B.n122 B.n50 71.676
R1914 B.n118 B.n49 71.676
R1915 B.n706 B.n463 71.676
R1916 B.n698 B.n404 71.676
R1917 B.n694 B.n405 71.676
R1918 B.n690 B.n406 71.676
R1919 B.n686 B.n407 71.676
R1920 B.n682 B.n408 71.676
R1921 B.n678 B.n409 71.676
R1922 B.n674 B.n410 71.676
R1923 B.n670 B.n411 71.676
R1924 B.n666 B.n412 71.676
R1925 B.n662 B.n413 71.676
R1926 B.n658 B.n414 71.676
R1927 B.n654 B.n415 71.676
R1928 B.n650 B.n416 71.676
R1929 B.n646 B.n417 71.676
R1930 B.n642 B.n418 71.676
R1931 B.n638 B.n419 71.676
R1932 B.n634 B.n420 71.676
R1933 B.n630 B.n421 71.676
R1934 B.n626 B.n422 71.676
R1935 B.n622 B.n423 71.676
R1936 B.n618 B.n424 71.676
R1937 B.n614 B.n425 71.676
R1938 B.n610 B.n426 71.676
R1939 B.n606 B.n427 71.676
R1940 B.n602 B.n428 71.676
R1941 B.n598 B.n429 71.676
R1942 B.n593 B.n430 71.676
R1943 B.n589 B.n431 71.676
R1944 B.n585 B.n432 71.676
R1945 B.n581 B.n433 71.676
R1946 B.n577 B.n434 71.676
R1947 B.n573 B.n435 71.676
R1948 B.n569 B.n436 71.676
R1949 B.n565 B.n437 71.676
R1950 B.n561 B.n438 71.676
R1951 B.n557 B.n439 71.676
R1952 B.n553 B.n440 71.676
R1953 B.n549 B.n441 71.676
R1954 B.n545 B.n442 71.676
R1955 B.n541 B.n443 71.676
R1956 B.n537 B.n444 71.676
R1957 B.n533 B.n445 71.676
R1958 B.n529 B.n446 71.676
R1959 B.n525 B.n447 71.676
R1960 B.n521 B.n448 71.676
R1961 B.n517 B.n449 71.676
R1962 B.n513 B.n450 71.676
R1963 B.n509 B.n451 71.676
R1964 B.n505 B.n452 71.676
R1965 B.n501 B.n453 71.676
R1966 B.n497 B.n454 71.676
R1967 B.n493 B.n455 71.676
R1968 B.n489 B.n456 71.676
R1969 B.n485 B.n457 71.676
R1970 B.n481 B.n458 71.676
R1971 B.n477 B.n459 71.676
R1972 B.n473 B.n460 71.676
R1973 B.n469 B.n461 71.676
R1974 B.n709 B.n708 71.676
R1975 B.n707 B.n400 69.2017
R1976 B.n821 B.n820 69.2017
R1977 B.n468 B.n467 59.5399
R1978 B.n595 B.n465 59.5399
R1979 B.n114 B.n113 59.5399
R1980 B.n245 B.n111 59.5399
R1981 B.n818 B.n817 35.7468
R1982 B.n116 B.n45 35.7468
R1983 B.n711 B.n710 35.7468
R1984 B.n704 B.n398 35.7468
R1985 B.n714 B.n400 33.8543
R1986 B.n714 B.n395 33.8543
R1987 B.n720 B.n395 33.8543
R1988 B.n720 B.n396 33.8543
R1989 B.n726 B.n388 33.8543
R1990 B.n732 B.n388 33.8543
R1991 B.n732 B.n384 33.8543
R1992 B.n739 B.n384 33.8543
R1993 B.n739 B.n738 33.8543
R1994 B.n745 B.n377 33.8543
R1995 B.n751 B.n377 33.8543
R1996 B.n757 B.n372 33.8543
R1997 B.n757 B.n373 33.8543
R1998 B.n763 B.n365 33.8543
R1999 B.n769 B.n365 33.8543
R2000 B.n776 B.n361 33.8543
R2001 B.n782 B.n357 33.8543
R2002 B.n782 B.n4 33.8543
R2003 B.n870 B.n4 33.8543
R2004 B.n870 B.n869 33.8543
R2005 B.n869 B.n868 33.8543
R2006 B.n868 B.n8 33.8543
R2007 B.n862 B.n861 33.8543
R2008 B.n860 B.n15 33.8543
R2009 B.n854 B.n15 33.8543
R2010 B.n853 B.n852 33.8543
R2011 B.n852 B.n22 33.8543
R2012 B.n846 B.n845 33.8543
R2013 B.n845 B.n844 33.8543
R2014 B.n838 B.n32 33.8543
R2015 B.n838 B.n837 33.8543
R2016 B.n837 B.n836 33.8543
R2017 B.n836 B.n36 33.8543
R2018 B.n830 B.n36 33.8543
R2019 B.n829 B.n828 33.8543
R2020 B.n828 B.n43 33.8543
R2021 B.n822 B.n43 33.8543
R2022 B.n822 B.n821 33.8543
R2023 B.n776 B.t7 32.8586
R2024 B.n862 B.t1 32.8586
R2025 B.t9 B.n361 29.8715
R2026 B.n861 B.t4 29.8715
R2027 B.n763 B.t5 24.893
R2028 B.n854 B.t0 24.893
R2029 B.t2 B.n372 19.9145
R2030 B.t3 B.n22 19.9145
R2031 B.n738 B.t8 18.9188
R2032 B.n32 B.t6 18.9188
R2033 B.n467 B.n466 18.8126
R2034 B.n465 B.n464 18.8126
R2035 B.n113 B.n112 18.8126
R2036 B.n111 B.n110 18.8126
R2037 B B.n872 18.0485
R2038 B.n396 B.t18 16.9274
R2039 B.n726 B.t18 16.9274
R2040 B.n830 B.t11 16.9274
R2041 B.t11 B.n829 16.9274
R2042 B.n745 B.t8 14.936
R2043 B.n844 B.t6 14.936
R2044 B.n751 B.t2 13.9403
R2045 B.n846 B.t3 13.9403
R2046 B.n117 B.n116 10.6151
R2047 B.n120 B.n117 10.6151
R2048 B.n121 B.n120 10.6151
R2049 B.n124 B.n121 10.6151
R2050 B.n125 B.n124 10.6151
R2051 B.n128 B.n125 10.6151
R2052 B.n129 B.n128 10.6151
R2053 B.n132 B.n129 10.6151
R2054 B.n133 B.n132 10.6151
R2055 B.n136 B.n133 10.6151
R2056 B.n137 B.n136 10.6151
R2057 B.n140 B.n137 10.6151
R2058 B.n141 B.n140 10.6151
R2059 B.n144 B.n141 10.6151
R2060 B.n145 B.n144 10.6151
R2061 B.n148 B.n145 10.6151
R2062 B.n149 B.n148 10.6151
R2063 B.n152 B.n149 10.6151
R2064 B.n153 B.n152 10.6151
R2065 B.n156 B.n153 10.6151
R2066 B.n157 B.n156 10.6151
R2067 B.n160 B.n157 10.6151
R2068 B.n161 B.n160 10.6151
R2069 B.n164 B.n161 10.6151
R2070 B.n165 B.n164 10.6151
R2071 B.n168 B.n165 10.6151
R2072 B.n169 B.n168 10.6151
R2073 B.n172 B.n169 10.6151
R2074 B.n173 B.n172 10.6151
R2075 B.n176 B.n173 10.6151
R2076 B.n177 B.n176 10.6151
R2077 B.n180 B.n177 10.6151
R2078 B.n181 B.n180 10.6151
R2079 B.n184 B.n181 10.6151
R2080 B.n185 B.n184 10.6151
R2081 B.n188 B.n185 10.6151
R2082 B.n189 B.n188 10.6151
R2083 B.n192 B.n189 10.6151
R2084 B.n193 B.n192 10.6151
R2085 B.n196 B.n193 10.6151
R2086 B.n197 B.n196 10.6151
R2087 B.n200 B.n197 10.6151
R2088 B.n201 B.n200 10.6151
R2089 B.n204 B.n201 10.6151
R2090 B.n205 B.n204 10.6151
R2091 B.n208 B.n205 10.6151
R2092 B.n209 B.n208 10.6151
R2093 B.n212 B.n209 10.6151
R2094 B.n213 B.n212 10.6151
R2095 B.n216 B.n213 10.6151
R2096 B.n217 B.n216 10.6151
R2097 B.n220 B.n217 10.6151
R2098 B.n221 B.n220 10.6151
R2099 B.n224 B.n221 10.6151
R2100 B.n225 B.n224 10.6151
R2101 B.n229 B.n228 10.6151
R2102 B.n232 B.n229 10.6151
R2103 B.n233 B.n232 10.6151
R2104 B.n236 B.n233 10.6151
R2105 B.n237 B.n236 10.6151
R2106 B.n240 B.n237 10.6151
R2107 B.n241 B.n240 10.6151
R2108 B.n244 B.n241 10.6151
R2109 B.n249 B.n246 10.6151
R2110 B.n250 B.n249 10.6151
R2111 B.n253 B.n250 10.6151
R2112 B.n254 B.n253 10.6151
R2113 B.n257 B.n254 10.6151
R2114 B.n258 B.n257 10.6151
R2115 B.n261 B.n258 10.6151
R2116 B.n262 B.n261 10.6151
R2117 B.n265 B.n262 10.6151
R2118 B.n266 B.n265 10.6151
R2119 B.n269 B.n266 10.6151
R2120 B.n270 B.n269 10.6151
R2121 B.n273 B.n270 10.6151
R2122 B.n274 B.n273 10.6151
R2123 B.n277 B.n274 10.6151
R2124 B.n278 B.n277 10.6151
R2125 B.n281 B.n278 10.6151
R2126 B.n282 B.n281 10.6151
R2127 B.n285 B.n282 10.6151
R2128 B.n286 B.n285 10.6151
R2129 B.n289 B.n286 10.6151
R2130 B.n290 B.n289 10.6151
R2131 B.n293 B.n290 10.6151
R2132 B.n294 B.n293 10.6151
R2133 B.n297 B.n294 10.6151
R2134 B.n298 B.n297 10.6151
R2135 B.n301 B.n298 10.6151
R2136 B.n302 B.n301 10.6151
R2137 B.n305 B.n302 10.6151
R2138 B.n306 B.n305 10.6151
R2139 B.n309 B.n306 10.6151
R2140 B.n310 B.n309 10.6151
R2141 B.n313 B.n310 10.6151
R2142 B.n314 B.n313 10.6151
R2143 B.n317 B.n314 10.6151
R2144 B.n318 B.n317 10.6151
R2145 B.n321 B.n318 10.6151
R2146 B.n322 B.n321 10.6151
R2147 B.n325 B.n322 10.6151
R2148 B.n326 B.n325 10.6151
R2149 B.n329 B.n326 10.6151
R2150 B.n330 B.n329 10.6151
R2151 B.n333 B.n330 10.6151
R2152 B.n334 B.n333 10.6151
R2153 B.n337 B.n334 10.6151
R2154 B.n338 B.n337 10.6151
R2155 B.n341 B.n338 10.6151
R2156 B.n342 B.n341 10.6151
R2157 B.n345 B.n342 10.6151
R2158 B.n346 B.n345 10.6151
R2159 B.n349 B.n346 10.6151
R2160 B.n350 B.n349 10.6151
R2161 B.n353 B.n350 10.6151
R2162 B.n354 B.n353 10.6151
R2163 B.n818 B.n354 10.6151
R2164 B.n712 B.n711 10.6151
R2165 B.n712 B.n393 10.6151
R2166 B.n722 B.n393 10.6151
R2167 B.n723 B.n722 10.6151
R2168 B.n724 B.n723 10.6151
R2169 B.n724 B.n386 10.6151
R2170 B.n734 B.n386 10.6151
R2171 B.n735 B.n734 10.6151
R2172 B.n736 B.n735 10.6151
R2173 B.n736 B.n379 10.6151
R2174 B.n747 B.n379 10.6151
R2175 B.n748 B.n747 10.6151
R2176 B.n749 B.n748 10.6151
R2177 B.n749 B.n370 10.6151
R2178 B.n759 B.n370 10.6151
R2179 B.n760 B.n759 10.6151
R2180 B.n761 B.n760 10.6151
R2181 B.n761 B.n363 10.6151
R2182 B.n771 B.n363 10.6151
R2183 B.n772 B.n771 10.6151
R2184 B.n774 B.n772 10.6151
R2185 B.n774 B.n773 10.6151
R2186 B.n773 B.n355 10.6151
R2187 B.n785 B.n355 10.6151
R2188 B.n786 B.n785 10.6151
R2189 B.n787 B.n786 10.6151
R2190 B.n788 B.n787 10.6151
R2191 B.n790 B.n788 10.6151
R2192 B.n791 B.n790 10.6151
R2193 B.n792 B.n791 10.6151
R2194 B.n793 B.n792 10.6151
R2195 B.n795 B.n793 10.6151
R2196 B.n796 B.n795 10.6151
R2197 B.n797 B.n796 10.6151
R2198 B.n798 B.n797 10.6151
R2199 B.n800 B.n798 10.6151
R2200 B.n801 B.n800 10.6151
R2201 B.n802 B.n801 10.6151
R2202 B.n803 B.n802 10.6151
R2203 B.n805 B.n803 10.6151
R2204 B.n806 B.n805 10.6151
R2205 B.n807 B.n806 10.6151
R2206 B.n808 B.n807 10.6151
R2207 B.n810 B.n808 10.6151
R2208 B.n811 B.n810 10.6151
R2209 B.n812 B.n811 10.6151
R2210 B.n813 B.n812 10.6151
R2211 B.n815 B.n813 10.6151
R2212 B.n816 B.n815 10.6151
R2213 B.n817 B.n816 10.6151
R2214 B.n704 B.n703 10.6151
R2215 B.n703 B.n702 10.6151
R2216 B.n702 B.n701 10.6151
R2217 B.n701 B.n699 10.6151
R2218 B.n699 B.n696 10.6151
R2219 B.n696 B.n695 10.6151
R2220 B.n695 B.n692 10.6151
R2221 B.n692 B.n691 10.6151
R2222 B.n691 B.n688 10.6151
R2223 B.n688 B.n687 10.6151
R2224 B.n687 B.n684 10.6151
R2225 B.n684 B.n683 10.6151
R2226 B.n683 B.n680 10.6151
R2227 B.n680 B.n679 10.6151
R2228 B.n679 B.n676 10.6151
R2229 B.n676 B.n675 10.6151
R2230 B.n675 B.n672 10.6151
R2231 B.n672 B.n671 10.6151
R2232 B.n671 B.n668 10.6151
R2233 B.n668 B.n667 10.6151
R2234 B.n667 B.n664 10.6151
R2235 B.n664 B.n663 10.6151
R2236 B.n663 B.n660 10.6151
R2237 B.n660 B.n659 10.6151
R2238 B.n659 B.n656 10.6151
R2239 B.n656 B.n655 10.6151
R2240 B.n655 B.n652 10.6151
R2241 B.n652 B.n651 10.6151
R2242 B.n651 B.n648 10.6151
R2243 B.n648 B.n647 10.6151
R2244 B.n647 B.n644 10.6151
R2245 B.n644 B.n643 10.6151
R2246 B.n643 B.n640 10.6151
R2247 B.n640 B.n639 10.6151
R2248 B.n639 B.n636 10.6151
R2249 B.n636 B.n635 10.6151
R2250 B.n635 B.n632 10.6151
R2251 B.n632 B.n631 10.6151
R2252 B.n631 B.n628 10.6151
R2253 B.n628 B.n627 10.6151
R2254 B.n627 B.n624 10.6151
R2255 B.n624 B.n623 10.6151
R2256 B.n623 B.n620 10.6151
R2257 B.n620 B.n619 10.6151
R2258 B.n619 B.n616 10.6151
R2259 B.n616 B.n615 10.6151
R2260 B.n615 B.n612 10.6151
R2261 B.n612 B.n611 10.6151
R2262 B.n611 B.n608 10.6151
R2263 B.n608 B.n607 10.6151
R2264 B.n607 B.n604 10.6151
R2265 B.n604 B.n603 10.6151
R2266 B.n603 B.n600 10.6151
R2267 B.n600 B.n599 10.6151
R2268 B.n599 B.n596 10.6151
R2269 B.n594 B.n591 10.6151
R2270 B.n591 B.n590 10.6151
R2271 B.n590 B.n587 10.6151
R2272 B.n587 B.n586 10.6151
R2273 B.n586 B.n583 10.6151
R2274 B.n583 B.n582 10.6151
R2275 B.n582 B.n579 10.6151
R2276 B.n579 B.n578 10.6151
R2277 B.n575 B.n574 10.6151
R2278 B.n574 B.n571 10.6151
R2279 B.n571 B.n570 10.6151
R2280 B.n570 B.n567 10.6151
R2281 B.n567 B.n566 10.6151
R2282 B.n566 B.n563 10.6151
R2283 B.n563 B.n562 10.6151
R2284 B.n562 B.n559 10.6151
R2285 B.n559 B.n558 10.6151
R2286 B.n558 B.n555 10.6151
R2287 B.n555 B.n554 10.6151
R2288 B.n554 B.n551 10.6151
R2289 B.n551 B.n550 10.6151
R2290 B.n550 B.n547 10.6151
R2291 B.n547 B.n546 10.6151
R2292 B.n546 B.n543 10.6151
R2293 B.n543 B.n542 10.6151
R2294 B.n542 B.n539 10.6151
R2295 B.n539 B.n538 10.6151
R2296 B.n538 B.n535 10.6151
R2297 B.n535 B.n534 10.6151
R2298 B.n534 B.n531 10.6151
R2299 B.n531 B.n530 10.6151
R2300 B.n530 B.n527 10.6151
R2301 B.n527 B.n526 10.6151
R2302 B.n526 B.n523 10.6151
R2303 B.n523 B.n522 10.6151
R2304 B.n522 B.n519 10.6151
R2305 B.n519 B.n518 10.6151
R2306 B.n518 B.n515 10.6151
R2307 B.n515 B.n514 10.6151
R2308 B.n514 B.n511 10.6151
R2309 B.n511 B.n510 10.6151
R2310 B.n510 B.n507 10.6151
R2311 B.n507 B.n506 10.6151
R2312 B.n506 B.n503 10.6151
R2313 B.n503 B.n502 10.6151
R2314 B.n502 B.n499 10.6151
R2315 B.n499 B.n498 10.6151
R2316 B.n498 B.n495 10.6151
R2317 B.n495 B.n494 10.6151
R2318 B.n494 B.n491 10.6151
R2319 B.n491 B.n490 10.6151
R2320 B.n490 B.n487 10.6151
R2321 B.n487 B.n486 10.6151
R2322 B.n486 B.n483 10.6151
R2323 B.n483 B.n482 10.6151
R2324 B.n482 B.n479 10.6151
R2325 B.n479 B.n478 10.6151
R2326 B.n478 B.n475 10.6151
R2327 B.n475 B.n474 10.6151
R2328 B.n474 B.n471 10.6151
R2329 B.n471 B.n470 10.6151
R2330 B.n470 B.n402 10.6151
R2331 B.n710 B.n402 10.6151
R2332 B.n716 B.n398 10.6151
R2333 B.n717 B.n716 10.6151
R2334 B.n718 B.n717 10.6151
R2335 B.n718 B.n390 10.6151
R2336 B.n728 B.n390 10.6151
R2337 B.n729 B.n728 10.6151
R2338 B.n730 B.n729 10.6151
R2339 B.n730 B.n382 10.6151
R2340 B.n741 B.n382 10.6151
R2341 B.n742 B.n741 10.6151
R2342 B.n743 B.n742 10.6151
R2343 B.n743 B.n375 10.6151
R2344 B.n753 B.n375 10.6151
R2345 B.n754 B.n753 10.6151
R2346 B.n755 B.n754 10.6151
R2347 B.n755 B.n367 10.6151
R2348 B.n765 B.n367 10.6151
R2349 B.n766 B.n765 10.6151
R2350 B.n767 B.n766 10.6151
R2351 B.n767 B.n359 10.6151
R2352 B.n778 B.n359 10.6151
R2353 B.n779 B.n778 10.6151
R2354 B.n780 B.n779 10.6151
R2355 B.n780 B.n0 10.6151
R2356 B.n866 B.n1 10.6151
R2357 B.n866 B.n865 10.6151
R2358 B.n865 B.n864 10.6151
R2359 B.n864 B.n10 10.6151
R2360 B.n858 B.n10 10.6151
R2361 B.n858 B.n857 10.6151
R2362 B.n857 B.n856 10.6151
R2363 B.n856 B.n17 10.6151
R2364 B.n850 B.n17 10.6151
R2365 B.n850 B.n849 10.6151
R2366 B.n849 B.n848 10.6151
R2367 B.n848 B.n24 10.6151
R2368 B.n842 B.n24 10.6151
R2369 B.n842 B.n841 10.6151
R2370 B.n841 B.n840 10.6151
R2371 B.n840 B.n30 10.6151
R2372 B.n834 B.n30 10.6151
R2373 B.n834 B.n833 10.6151
R2374 B.n833 B.n832 10.6151
R2375 B.n832 B.n38 10.6151
R2376 B.n826 B.n38 10.6151
R2377 B.n826 B.n825 10.6151
R2378 B.n825 B.n824 10.6151
R2379 B.n824 B.n45 10.6151
R2380 B.n373 B.t5 8.9618
R2381 B.t0 B.n853 8.9618
R2382 B.n228 B.n114 6.5566
R2383 B.n245 B.n244 6.5566
R2384 B.n595 B.n594 6.5566
R2385 B.n578 B.n468 6.5566
R2386 B.n225 B.n114 4.05904
R2387 B.n246 B.n245 4.05904
R2388 B.n596 B.n595 4.05904
R2389 B.n575 B.n468 4.05904
R2390 B.n769 B.t9 3.9833
R2391 B.t4 B.n860 3.9833
R2392 B.n872 B.n0 2.81026
R2393 B.n872 B.n1 2.81026
R2394 B.t7 B.n357 0.9962
R2395 B.t1 B.n8 0.9962
R2396 VP.n4 VP.t1 721.58
R2397 VP.n10 VP.t9 694.759
R2398 VP.n1 VP.t0 694.759
R2399 VP.n14 VP.t3 694.759
R2400 VP.n15 VP.t6 694.759
R2401 VP.n16 VP.t7 694.759
R2402 VP.n8 VP.t4 694.759
R2403 VP.n7 VP.t2 694.759
R2404 VP.n6 VP.t8 694.759
R2405 VP.n5 VP.t5 694.759
R2406 VP.n17 VP.n16 161.3
R2407 VP.n9 VP.n8 161.3
R2408 VP.n11 VP.n10 161.3
R2409 VP.n6 VP.n3 80.6037
R2410 VP.n7 VP.n2 80.6037
R2411 VP.n15 VP.n0 80.6037
R2412 VP.n14 VP.n13 80.6037
R2413 VP.n12 VP.n1 80.6037
R2414 VP.n10 VP.n1 48.2005
R2415 VP.n14 VP.n1 48.2005
R2416 VP.n15 VP.n14 48.2005
R2417 VP.n16 VP.n15 48.2005
R2418 VP.n8 VP.n7 48.2005
R2419 VP.n7 VP.n6 48.2005
R2420 VP.n6 VP.n5 48.2005
R2421 VP.n11 VP.n9 46.1937
R2422 VP.n4 VP.n3 45.2318
R2423 VP.n5 VP.n4 13.3799
R2424 VP.n3 VP.n2 0.380177
R2425 VP.n13 VP.n12 0.380177
R2426 VP.n13 VP.n0 0.380177
R2427 VP.n9 VP.n2 0.285035
R2428 VP.n12 VP.n11 0.285035
R2429 VP.n17 VP.n0 0.285035
R2430 VP VP.n17 0.0516364
R2431 VDD1.n88 VDD1.n0 289.615
R2432 VDD1.n183 VDD1.n95 289.615
R2433 VDD1.n89 VDD1.n88 185
R2434 VDD1.n87 VDD1.n86 185
R2435 VDD1.n4 VDD1.n3 185
R2436 VDD1.n81 VDD1.n80 185
R2437 VDD1.n79 VDD1.n78 185
R2438 VDD1.n77 VDD1.n7 185
R2439 VDD1.n11 VDD1.n8 185
R2440 VDD1.n72 VDD1.n71 185
R2441 VDD1.n70 VDD1.n69 185
R2442 VDD1.n13 VDD1.n12 185
R2443 VDD1.n64 VDD1.n63 185
R2444 VDD1.n62 VDD1.n61 185
R2445 VDD1.n17 VDD1.n16 185
R2446 VDD1.n56 VDD1.n55 185
R2447 VDD1.n54 VDD1.n53 185
R2448 VDD1.n21 VDD1.n20 185
R2449 VDD1.n48 VDD1.n47 185
R2450 VDD1.n46 VDD1.n45 185
R2451 VDD1.n25 VDD1.n24 185
R2452 VDD1.n40 VDD1.n39 185
R2453 VDD1.n38 VDD1.n37 185
R2454 VDD1.n29 VDD1.n28 185
R2455 VDD1.n32 VDD1.n31 185
R2456 VDD1.n126 VDD1.n125 185
R2457 VDD1.n123 VDD1.n122 185
R2458 VDD1.n132 VDD1.n131 185
R2459 VDD1.n134 VDD1.n133 185
R2460 VDD1.n119 VDD1.n118 185
R2461 VDD1.n140 VDD1.n139 185
R2462 VDD1.n142 VDD1.n141 185
R2463 VDD1.n115 VDD1.n114 185
R2464 VDD1.n148 VDD1.n147 185
R2465 VDD1.n150 VDD1.n149 185
R2466 VDD1.n111 VDD1.n110 185
R2467 VDD1.n156 VDD1.n155 185
R2468 VDD1.n158 VDD1.n157 185
R2469 VDD1.n107 VDD1.n106 185
R2470 VDD1.n164 VDD1.n163 185
R2471 VDD1.n167 VDD1.n166 185
R2472 VDD1.n165 VDD1.n103 185
R2473 VDD1.n172 VDD1.n102 185
R2474 VDD1.n174 VDD1.n173 185
R2475 VDD1.n176 VDD1.n175 185
R2476 VDD1.n99 VDD1.n98 185
R2477 VDD1.n182 VDD1.n181 185
R2478 VDD1.n184 VDD1.n183 185
R2479 VDD1.t8 VDD1.n30 147.659
R2480 VDD1.t0 VDD1.n124 147.659
R2481 VDD1.n88 VDD1.n87 104.615
R2482 VDD1.n87 VDD1.n3 104.615
R2483 VDD1.n80 VDD1.n3 104.615
R2484 VDD1.n80 VDD1.n79 104.615
R2485 VDD1.n79 VDD1.n7 104.615
R2486 VDD1.n11 VDD1.n7 104.615
R2487 VDD1.n71 VDD1.n11 104.615
R2488 VDD1.n71 VDD1.n70 104.615
R2489 VDD1.n70 VDD1.n12 104.615
R2490 VDD1.n63 VDD1.n12 104.615
R2491 VDD1.n63 VDD1.n62 104.615
R2492 VDD1.n62 VDD1.n16 104.615
R2493 VDD1.n55 VDD1.n16 104.615
R2494 VDD1.n55 VDD1.n54 104.615
R2495 VDD1.n54 VDD1.n20 104.615
R2496 VDD1.n47 VDD1.n20 104.615
R2497 VDD1.n47 VDD1.n46 104.615
R2498 VDD1.n46 VDD1.n24 104.615
R2499 VDD1.n39 VDD1.n24 104.615
R2500 VDD1.n39 VDD1.n38 104.615
R2501 VDD1.n38 VDD1.n28 104.615
R2502 VDD1.n31 VDD1.n28 104.615
R2503 VDD1.n125 VDD1.n122 104.615
R2504 VDD1.n132 VDD1.n122 104.615
R2505 VDD1.n133 VDD1.n132 104.615
R2506 VDD1.n133 VDD1.n118 104.615
R2507 VDD1.n140 VDD1.n118 104.615
R2508 VDD1.n141 VDD1.n140 104.615
R2509 VDD1.n141 VDD1.n114 104.615
R2510 VDD1.n148 VDD1.n114 104.615
R2511 VDD1.n149 VDD1.n148 104.615
R2512 VDD1.n149 VDD1.n110 104.615
R2513 VDD1.n156 VDD1.n110 104.615
R2514 VDD1.n157 VDD1.n156 104.615
R2515 VDD1.n157 VDD1.n106 104.615
R2516 VDD1.n164 VDD1.n106 104.615
R2517 VDD1.n166 VDD1.n164 104.615
R2518 VDD1.n166 VDD1.n165 104.615
R2519 VDD1.n165 VDD1.n102 104.615
R2520 VDD1.n174 VDD1.n102 104.615
R2521 VDD1.n175 VDD1.n174 104.615
R2522 VDD1.n175 VDD1.n98 104.615
R2523 VDD1.n182 VDD1.n98 104.615
R2524 VDD1.n183 VDD1.n182 104.615
R2525 VDD1.n191 VDD1.n190 61.6843
R2526 VDD1.n94 VDD1.n93 61.1127
R2527 VDD1.n193 VDD1.n192 61.1125
R2528 VDD1.n189 VDD1.n188 61.1125
R2529 VDD1.n31 VDD1.t8 52.3082
R2530 VDD1.n125 VDD1.t0 52.3082
R2531 VDD1.n94 VDD1.n92 50.0882
R2532 VDD1.n189 VDD1.n187 50.0882
R2533 VDD1.n193 VDD1.n191 43.1884
R2534 VDD1.n32 VDD1.n30 15.6677
R2535 VDD1.n126 VDD1.n124 15.6677
R2536 VDD1.n78 VDD1.n77 13.1884
R2537 VDD1.n173 VDD1.n172 13.1884
R2538 VDD1.n81 VDD1.n6 12.8005
R2539 VDD1.n76 VDD1.n8 12.8005
R2540 VDD1.n33 VDD1.n29 12.8005
R2541 VDD1.n127 VDD1.n123 12.8005
R2542 VDD1.n171 VDD1.n103 12.8005
R2543 VDD1.n176 VDD1.n101 12.8005
R2544 VDD1.n82 VDD1.n4 12.0247
R2545 VDD1.n73 VDD1.n72 12.0247
R2546 VDD1.n37 VDD1.n36 12.0247
R2547 VDD1.n131 VDD1.n130 12.0247
R2548 VDD1.n168 VDD1.n167 12.0247
R2549 VDD1.n177 VDD1.n99 12.0247
R2550 VDD1.n86 VDD1.n85 11.249
R2551 VDD1.n69 VDD1.n10 11.249
R2552 VDD1.n40 VDD1.n27 11.249
R2553 VDD1.n134 VDD1.n121 11.249
R2554 VDD1.n163 VDD1.n105 11.249
R2555 VDD1.n181 VDD1.n180 11.249
R2556 VDD1.n89 VDD1.n2 10.4732
R2557 VDD1.n68 VDD1.n13 10.4732
R2558 VDD1.n41 VDD1.n25 10.4732
R2559 VDD1.n135 VDD1.n119 10.4732
R2560 VDD1.n162 VDD1.n107 10.4732
R2561 VDD1.n184 VDD1.n97 10.4732
R2562 VDD1.n90 VDD1.n0 9.69747
R2563 VDD1.n65 VDD1.n64 9.69747
R2564 VDD1.n45 VDD1.n44 9.69747
R2565 VDD1.n139 VDD1.n138 9.69747
R2566 VDD1.n159 VDD1.n158 9.69747
R2567 VDD1.n185 VDD1.n95 9.69747
R2568 VDD1.n92 VDD1.n91 9.45567
R2569 VDD1.n187 VDD1.n186 9.45567
R2570 VDD1.n58 VDD1.n57 9.3005
R2571 VDD1.n60 VDD1.n59 9.3005
R2572 VDD1.n15 VDD1.n14 9.3005
R2573 VDD1.n66 VDD1.n65 9.3005
R2574 VDD1.n68 VDD1.n67 9.3005
R2575 VDD1.n10 VDD1.n9 9.3005
R2576 VDD1.n74 VDD1.n73 9.3005
R2577 VDD1.n76 VDD1.n75 9.3005
R2578 VDD1.n91 VDD1.n90 9.3005
R2579 VDD1.n2 VDD1.n1 9.3005
R2580 VDD1.n85 VDD1.n84 9.3005
R2581 VDD1.n83 VDD1.n82 9.3005
R2582 VDD1.n6 VDD1.n5 9.3005
R2583 VDD1.n19 VDD1.n18 9.3005
R2584 VDD1.n52 VDD1.n51 9.3005
R2585 VDD1.n50 VDD1.n49 9.3005
R2586 VDD1.n23 VDD1.n22 9.3005
R2587 VDD1.n44 VDD1.n43 9.3005
R2588 VDD1.n42 VDD1.n41 9.3005
R2589 VDD1.n27 VDD1.n26 9.3005
R2590 VDD1.n36 VDD1.n35 9.3005
R2591 VDD1.n34 VDD1.n33 9.3005
R2592 VDD1.n186 VDD1.n185 9.3005
R2593 VDD1.n97 VDD1.n96 9.3005
R2594 VDD1.n180 VDD1.n179 9.3005
R2595 VDD1.n178 VDD1.n177 9.3005
R2596 VDD1.n101 VDD1.n100 9.3005
R2597 VDD1.n146 VDD1.n145 9.3005
R2598 VDD1.n144 VDD1.n143 9.3005
R2599 VDD1.n117 VDD1.n116 9.3005
R2600 VDD1.n138 VDD1.n137 9.3005
R2601 VDD1.n136 VDD1.n135 9.3005
R2602 VDD1.n121 VDD1.n120 9.3005
R2603 VDD1.n130 VDD1.n129 9.3005
R2604 VDD1.n128 VDD1.n127 9.3005
R2605 VDD1.n113 VDD1.n112 9.3005
R2606 VDD1.n152 VDD1.n151 9.3005
R2607 VDD1.n154 VDD1.n153 9.3005
R2608 VDD1.n109 VDD1.n108 9.3005
R2609 VDD1.n160 VDD1.n159 9.3005
R2610 VDD1.n162 VDD1.n161 9.3005
R2611 VDD1.n105 VDD1.n104 9.3005
R2612 VDD1.n169 VDD1.n168 9.3005
R2613 VDD1.n171 VDD1.n170 9.3005
R2614 VDD1.n61 VDD1.n15 8.92171
R2615 VDD1.n48 VDD1.n23 8.92171
R2616 VDD1.n142 VDD1.n117 8.92171
R2617 VDD1.n155 VDD1.n109 8.92171
R2618 VDD1.n60 VDD1.n17 8.14595
R2619 VDD1.n49 VDD1.n21 8.14595
R2620 VDD1.n143 VDD1.n115 8.14595
R2621 VDD1.n154 VDD1.n111 8.14595
R2622 VDD1.n57 VDD1.n56 7.3702
R2623 VDD1.n53 VDD1.n52 7.3702
R2624 VDD1.n147 VDD1.n146 7.3702
R2625 VDD1.n151 VDD1.n150 7.3702
R2626 VDD1.n56 VDD1.n19 6.59444
R2627 VDD1.n53 VDD1.n19 6.59444
R2628 VDD1.n147 VDD1.n113 6.59444
R2629 VDD1.n150 VDD1.n113 6.59444
R2630 VDD1.n57 VDD1.n17 5.81868
R2631 VDD1.n52 VDD1.n21 5.81868
R2632 VDD1.n146 VDD1.n115 5.81868
R2633 VDD1.n151 VDD1.n111 5.81868
R2634 VDD1.n61 VDD1.n60 5.04292
R2635 VDD1.n49 VDD1.n48 5.04292
R2636 VDD1.n143 VDD1.n142 5.04292
R2637 VDD1.n155 VDD1.n154 5.04292
R2638 VDD1.n34 VDD1.n30 4.38563
R2639 VDD1.n128 VDD1.n124 4.38563
R2640 VDD1.n92 VDD1.n0 4.26717
R2641 VDD1.n64 VDD1.n15 4.26717
R2642 VDD1.n45 VDD1.n23 4.26717
R2643 VDD1.n139 VDD1.n117 4.26717
R2644 VDD1.n158 VDD1.n109 4.26717
R2645 VDD1.n187 VDD1.n95 4.26717
R2646 VDD1.n90 VDD1.n89 3.49141
R2647 VDD1.n65 VDD1.n13 3.49141
R2648 VDD1.n44 VDD1.n25 3.49141
R2649 VDD1.n138 VDD1.n119 3.49141
R2650 VDD1.n159 VDD1.n107 3.49141
R2651 VDD1.n185 VDD1.n184 3.49141
R2652 VDD1.n86 VDD1.n2 2.71565
R2653 VDD1.n69 VDD1.n68 2.71565
R2654 VDD1.n41 VDD1.n40 2.71565
R2655 VDD1.n135 VDD1.n134 2.71565
R2656 VDD1.n163 VDD1.n162 2.71565
R2657 VDD1.n181 VDD1.n97 2.71565
R2658 VDD1.n85 VDD1.n4 1.93989
R2659 VDD1.n72 VDD1.n10 1.93989
R2660 VDD1.n37 VDD1.n27 1.93989
R2661 VDD1.n131 VDD1.n121 1.93989
R2662 VDD1.n167 VDD1.n105 1.93989
R2663 VDD1.n180 VDD1.n99 1.93989
R2664 VDD1.n192 VDD1.t7 1.17767
R2665 VDD1.n192 VDD1.t5 1.17767
R2666 VDD1.n93 VDD1.t4 1.17767
R2667 VDD1.n93 VDD1.t1 1.17767
R2668 VDD1.n190 VDD1.t3 1.17767
R2669 VDD1.n190 VDD1.t2 1.17767
R2670 VDD1.n188 VDD1.t9 1.17767
R2671 VDD1.n188 VDD1.t6 1.17767
R2672 VDD1.n82 VDD1.n81 1.16414
R2673 VDD1.n73 VDD1.n8 1.16414
R2674 VDD1.n36 VDD1.n29 1.16414
R2675 VDD1.n130 VDD1.n123 1.16414
R2676 VDD1.n168 VDD1.n103 1.16414
R2677 VDD1.n177 VDD1.n176 1.16414
R2678 VDD1 VDD1.n193 0.569465
R2679 VDD1.n78 VDD1.n6 0.388379
R2680 VDD1.n77 VDD1.n76 0.388379
R2681 VDD1.n33 VDD1.n32 0.388379
R2682 VDD1.n127 VDD1.n126 0.388379
R2683 VDD1.n172 VDD1.n171 0.388379
R2684 VDD1.n173 VDD1.n101 0.388379
R2685 VDD1 VDD1.n94 0.267741
R2686 VDD1.n91 VDD1.n1 0.155672
R2687 VDD1.n84 VDD1.n1 0.155672
R2688 VDD1.n84 VDD1.n83 0.155672
R2689 VDD1.n83 VDD1.n5 0.155672
R2690 VDD1.n75 VDD1.n5 0.155672
R2691 VDD1.n75 VDD1.n74 0.155672
R2692 VDD1.n74 VDD1.n9 0.155672
R2693 VDD1.n67 VDD1.n9 0.155672
R2694 VDD1.n67 VDD1.n66 0.155672
R2695 VDD1.n66 VDD1.n14 0.155672
R2696 VDD1.n59 VDD1.n14 0.155672
R2697 VDD1.n59 VDD1.n58 0.155672
R2698 VDD1.n58 VDD1.n18 0.155672
R2699 VDD1.n51 VDD1.n18 0.155672
R2700 VDD1.n51 VDD1.n50 0.155672
R2701 VDD1.n50 VDD1.n22 0.155672
R2702 VDD1.n43 VDD1.n22 0.155672
R2703 VDD1.n43 VDD1.n42 0.155672
R2704 VDD1.n42 VDD1.n26 0.155672
R2705 VDD1.n35 VDD1.n26 0.155672
R2706 VDD1.n35 VDD1.n34 0.155672
R2707 VDD1.n129 VDD1.n128 0.155672
R2708 VDD1.n129 VDD1.n120 0.155672
R2709 VDD1.n136 VDD1.n120 0.155672
R2710 VDD1.n137 VDD1.n136 0.155672
R2711 VDD1.n137 VDD1.n116 0.155672
R2712 VDD1.n144 VDD1.n116 0.155672
R2713 VDD1.n145 VDD1.n144 0.155672
R2714 VDD1.n145 VDD1.n112 0.155672
R2715 VDD1.n152 VDD1.n112 0.155672
R2716 VDD1.n153 VDD1.n152 0.155672
R2717 VDD1.n153 VDD1.n108 0.155672
R2718 VDD1.n160 VDD1.n108 0.155672
R2719 VDD1.n161 VDD1.n160 0.155672
R2720 VDD1.n161 VDD1.n104 0.155672
R2721 VDD1.n169 VDD1.n104 0.155672
R2722 VDD1.n170 VDD1.n169 0.155672
R2723 VDD1.n170 VDD1.n100 0.155672
R2724 VDD1.n178 VDD1.n100 0.155672
R2725 VDD1.n179 VDD1.n178 0.155672
R2726 VDD1.n179 VDD1.n96 0.155672
R2727 VDD1.n186 VDD1.n96 0.155672
R2728 VDD1.n191 VDD1.n189 0.154206
C0 VDD2 VN 8.75648f
C1 VDD2 VTAIL 19.7701f
C2 VDD1 VN 0.149339f
C3 VDD1 VTAIL 19.739302f
C4 VP VN 6.39551f
C5 VP VTAIL 8.389299f
C6 VDD1 VDD2 0.937327f
C7 VDD2 VP 0.335163f
C8 VN VTAIL 8.374459f
C9 VDD1 VP 8.93583f
C10 VDD2 B 5.769479f
C11 VDD1 B 5.686763f
C12 VTAIL B 8.189137f
C13 VN B 9.775981f
C14 VP B 7.52789f
C15 VDD1.n0 B 0.033906f
C16 VDD1.n1 B 0.024837f
C17 VDD1.n2 B 0.013347f
C18 VDD1.n3 B 0.031546f
C19 VDD1.n4 B 0.014132f
C20 VDD1.n5 B 0.024837f
C21 VDD1.n6 B 0.013347f
C22 VDD1.n7 B 0.031546f
C23 VDD1.n8 B 0.014132f
C24 VDD1.n9 B 0.024837f
C25 VDD1.n10 B 0.013347f
C26 VDD1.n11 B 0.031546f
C27 VDD1.n12 B 0.031546f
C28 VDD1.n13 B 0.014132f
C29 VDD1.n14 B 0.024837f
C30 VDD1.n15 B 0.013347f
C31 VDD1.n16 B 0.031546f
C32 VDD1.n17 B 0.014132f
C33 VDD1.n18 B 0.024837f
C34 VDD1.n19 B 0.013347f
C35 VDD1.n20 B 0.031546f
C36 VDD1.n21 B 0.014132f
C37 VDD1.n22 B 0.024837f
C38 VDD1.n23 B 0.013347f
C39 VDD1.n24 B 0.031546f
C40 VDD1.n25 B 0.014132f
C41 VDD1.n26 B 0.024837f
C42 VDD1.n27 B 0.013347f
C43 VDD1.n28 B 0.031546f
C44 VDD1.n29 B 0.014132f
C45 VDD1.n30 B 0.173328f
C46 VDD1.t8 B 0.052171f
C47 VDD1.n31 B 0.02366f
C48 VDD1.n32 B 0.018635f
C49 VDD1.n33 B 0.013347f
C50 VDD1.n34 B 1.82312f
C51 VDD1.n35 B 0.024837f
C52 VDD1.n36 B 0.013347f
C53 VDD1.n37 B 0.014132f
C54 VDD1.n38 B 0.031546f
C55 VDD1.n39 B 0.031546f
C56 VDD1.n40 B 0.014132f
C57 VDD1.n41 B 0.013347f
C58 VDD1.n42 B 0.024837f
C59 VDD1.n43 B 0.024837f
C60 VDD1.n44 B 0.013347f
C61 VDD1.n45 B 0.014132f
C62 VDD1.n46 B 0.031546f
C63 VDD1.n47 B 0.031546f
C64 VDD1.n48 B 0.014132f
C65 VDD1.n49 B 0.013347f
C66 VDD1.n50 B 0.024837f
C67 VDD1.n51 B 0.024837f
C68 VDD1.n52 B 0.013347f
C69 VDD1.n53 B 0.014132f
C70 VDD1.n54 B 0.031546f
C71 VDD1.n55 B 0.031546f
C72 VDD1.n56 B 0.014132f
C73 VDD1.n57 B 0.013347f
C74 VDD1.n58 B 0.024837f
C75 VDD1.n59 B 0.024837f
C76 VDD1.n60 B 0.013347f
C77 VDD1.n61 B 0.014132f
C78 VDD1.n62 B 0.031546f
C79 VDD1.n63 B 0.031546f
C80 VDD1.n64 B 0.014132f
C81 VDD1.n65 B 0.013347f
C82 VDD1.n66 B 0.024837f
C83 VDD1.n67 B 0.024837f
C84 VDD1.n68 B 0.013347f
C85 VDD1.n69 B 0.014132f
C86 VDD1.n70 B 0.031546f
C87 VDD1.n71 B 0.031546f
C88 VDD1.n72 B 0.014132f
C89 VDD1.n73 B 0.013347f
C90 VDD1.n74 B 0.024837f
C91 VDD1.n75 B 0.024837f
C92 VDD1.n76 B 0.013347f
C93 VDD1.n77 B 0.013739f
C94 VDD1.n78 B 0.013739f
C95 VDD1.n79 B 0.031546f
C96 VDD1.n80 B 0.031546f
C97 VDD1.n81 B 0.014132f
C98 VDD1.n82 B 0.013347f
C99 VDD1.n83 B 0.024837f
C100 VDD1.n84 B 0.024837f
C101 VDD1.n85 B 0.013347f
C102 VDD1.n86 B 0.014132f
C103 VDD1.n87 B 0.031546f
C104 VDD1.n88 B 0.066514f
C105 VDD1.n89 B 0.014132f
C106 VDD1.n90 B 0.013347f
C107 VDD1.n91 B 0.058089f
C108 VDD1.n92 B 0.056122f
C109 VDD1.t4 B 0.330129f
C110 VDD1.t1 B 0.330129f
C111 VDD1.n93 B 2.99947f
C112 VDD1.n94 B 0.406491f
C113 VDD1.n95 B 0.033906f
C114 VDD1.n96 B 0.024837f
C115 VDD1.n97 B 0.013347f
C116 VDD1.n98 B 0.031546f
C117 VDD1.n99 B 0.014132f
C118 VDD1.n100 B 0.024837f
C119 VDD1.n101 B 0.013347f
C120 VDD1.n102 B 0.031546f
C121 VDD1.n103 B 0.014132f
C122 VDD1.n104 B 0.024837f
C123 VDD1.n105 B 0.013347f
C124 VDD1.n106 B 0.031546f
C125 VDD1.n107 B 0.014132f
C126 VDD1.n108 B 0.024837f
C127 VDD1.n109 B 0.013347f
C128 VDD1.n110 B 0.031546f
C129 VDD1.n111 B 0.014132f
C130 VDD1.n112 B 0.024837f
C131 VDD1.n113 B 0.013347f
C132 VDD1.n114 B 0.031546f
C133 VDD1.n115 B 0.014132f
C134 VDD1.n116 B 0.024837f
C135 VDD1.n117 B 0.013347f
C136 VDD1.n118 B 0.031546f
C137 VDD1.n119 B 0.014132f
C138 VDD1.n120 B 0.024837f
C139 VDD1.n121 B 0.013347f
C140 VDD1.n122 B 0.031546f
C141 VDD1.n123 B 0.014132f
C142 VDD1.n124 B 0.173328f
C143 VDD1.t0 B 0.052171f
C144 VDD1.n125 B 0.02366f
C145 VDD1.n126 B 0.018635f
C146 VDD1.n127 B 0.013347f
C147 VDD1.n128 B 1.82312f
C148 VDD1.n129 B 0.024837f
C149 VDD1.n130 B 0.013347f
C150 VDD1.n131 B 0.014132f
C151 VDD1.n132 B 0.031546f
C152 VDD1.n133 B 0.031546f
C153 VDD1.n134 B 0.014132f
C154 VDD1.n135 B 0.013347f
C155 VDD1.n136 B 0.024837f
C156 VDD1.n137 B 0.024837f
C157 VDD1.n138 B 0.013347f
C158 VDD1.n139 B 0.014132f
C159 VDD1.n140 B 0.031546f
C160 VDD1.n141 B 0.031546f
C161 VDD1.n142 B 0.014132f
C162 VDD1.n143 B 0.013347f
C163 VDD1.n144 B 0.024837f
C164 VDD1.n145 B 0.024837f
C165 VDD1.n146 B 0.013347f
C166 VDD1.n147 B 0.014132f
C167 VDD1.n148 B 0.031546f
C168 VDD1.n149 B 0.031546f
C169 VDD1.n150 B 0.014132f
C170 VDD1.n151 B 0.013347f
C171 VDD1.n152 B 0.024837f
C172 VDD1.n153 B 0.024837f
C173 VDD1.n154 B 0.013347f
C174 VDD1.n155 B 0.014132f
C175 VDD1.n156 B 0.031546f
C176 VDD1.n157 B 0.031546f
C177 VDD1.n158 B 0.014132f
C178 VDD1.n159 B 0.013347f
C179 VDD1.n160 B 0.024837f
C180 VDD1.n161 B 0.024837f
C181 VDD1.n162 B 0.013347f
C182 VDD1.n163 B 0.014132f
C183 VDD1.n164 B 0.031546f
C184 VDD1.n165 B 0.031546f
C185 VDD1.n166 B 0.031546f
C186 VDD1.n167 B 0.014132f
C187 VDD1.n168 B 0.013347f
C188 VDD1.n169 B 0.024837f
C189 VDD1.n170 B 0.024837f
C190 VDD1.n171 B 0.013347f
C191 VDD1.n172 B 0.013739f
C192 VDD1.n173 B 0.013739f
C193 VDD1.n174 B 0.031546f
C194 VDD1.n175 B 0.031546f
C195 VDD1.n176 B 0.014132f
C196 VDD1.n177 B 0.013347f
C197 VDD1.n178 B 0.024837f
C198 VDD1.n179 B 0.024837f
C199 VDD1.n180 B 0.013347f
C200 VDD1.n181 B 0.014132f
C201 VDD1.n182 B 0.031546f
C202 VDD1.n183 B 0.066514f
C203 VDD1.n184 B 0.014132f
C204 VDD1.n185 B 0.013347f
C205 VDD1.n186 B 0.058089f
C206 VDD1.n187 B 0.056122f
C207 VDD1.t9 B 0.330129f
C208 VDD1.t6 B 0.330129f
C209 VDD1.n188 B 2.99946f
C210 VDD1.n189 B 0.401161f
C211 VDD1.t3 B 0.330129f
C212 VDD1.t2 B 0.330129f
C213 VDD1.n190 B 3.0025f
C214 VDD1.n191 B 2.23091f
C215 VDD1.t7 B 0.330129f
C216 VDD1.t5 B 0.330129f
C217 VDD1.n192 B 2.99946f
C218 VDD1.n193 B 2.71561f
C219 VP.n0 B 0.073781f
C220 VP.t0 B 1.35302f
C221 VP.n1 B 0.526195f
C222 VP.n2 B 0.073781f
C223 VP.t4 B 1.35302f
C224 VP.t2 B 1.35302f
C225 VP.t8 B 1.35302f
C226 VP.n3 B 0.234321f
C227 VP.t5 B 1.35302f
C228 VP.t1 B 1.37221f
C229 VP.n4 B 0.498316f
C230 VP.n5 B 0.526195f
C231 VP.n6 B 0.526195f
C232 VP.n7 B 0.526195f
C233 VP.n8 B 0.516144f
C234 VP.n9 B 2.14727f
C235 VP.t9 B 1.35302f
C236 VP.n10 B 0.516144f
C237 VP.n11 B 2.18184f
C238 VP.n12 B 0.073781f
C239 VP.n13 B 0.088593f
C240 VP.t3 B 1.35302f
C241 VP.n14 B 0.526195f
C242 VP.t6 B 1.35302f
C243 VP.n15 B 0.526195f
C244 VP.t7 B 1.35302f
C245 VP.n16 B 0.516144f
C246 VP.n17 B 0.04914f
C247 VTAIL.t14 B 0.339914f
C248 VTAIL.t8 B 0.339914f
C249 VTAIL.n0 B 3.01096f
C250 VTAIL.n1 B 0.383328f
C251 VTAIL.n2 B 0.034911f
C252 VTAIL.n3 B 0.025573f
C253 VTAIL.n4 B 0.013742f
C254 VTAIL.n5 B 0.032481f
C255 VTAIL.n6 B 0.01455f
C256 VTAIL.n7 B 0.025573f
C257 VTAIL.n8 B 0.013742f
C258 VTAIL.n9 B 0.032481f
C259 VTAIL.n10 B 0.01455f
C260 VTAIL.n11 B 0.025573f
C261 VTAIL.n12 B 0.013742f
C262 VTAIL.n13 B 0.032481f
C263 VTAIL.n14 B 0.01455f
C264 VTAIL.n15 B 0.025573f
C265 VTAIL.n16 B 0.013742f
C266 VTAIL.n17 B 0.032481f
C267 VTAIL.n18 B 0.01455f
C268 VTAIL.n19 B 0.025573f
C269 VTAIL.n20 B 0.013742f
C270 VTAIL.n21 B 0.032481f
C271 VTAIL.n22 B 0.01455f
C272 VTAIL.n23 B 0.025573f
C273 VTAIL.n24 B 0.013742f
C274 VTAIL.n25 B 0.032481f
C275 VTAIL.n26 B 0.01455f
C276 VTAIL.n27 B 0.025573f
C277 VTAIL.n28 B 0.013742f
C278 VTAIL.n29 B 0.032481f
C279 VTAIL.n30 B 0.01455f
C280 VTAIL.n31 B 0.178465f
C281 VTAIL.t16 B 0.053717f
C282 VTAIL.n32 B 0.024361f
C283 VTAIL.n33 B 0.019188f
C284 VTAIL.n34 B 0.013742f
C285 VTAIL.n35 B 1.87715f
C286 VTAIL.n36 B 0.025573f
C287 VTAIL.n37 B 0.013742f
C288 VTAIL.n38 B 0.01455f
C289 VTAIL.n39 B 0.032481f
C290 VTAIL.n40 B 0.032481f
C291 VTAIL.n41 B 0.01455f
C292 VTAIL.n42 B 0.013742f
C293 VTAIL.n43 B 0.025573f
C294 VTAIL.n44 B 0.025573f
C295 VTAIL.n45 B 0.013742f
C296 VTAIL.n46 B 0.01455f
C297 VTAIL.n47 B 0.032481f
C298 VTAIL.n48 B 0.032481f
C299 VTAIL.n49 B 0.01455f
C300 VTAIL.n50 B 0.013742f
C301 VTAIL.n51 B 0.025573f
C302 VTAIL.n52 B 0.025573f
C303 VTAIL.n53 B 0.013742f
C304 VTAIL.n54 B 0.01455f
C305 VTAIL.n55 B 0.032481f
C306 VTAIL.n56 B 0.032481f
C307 VTAIL.n57 B 0.01455f
C308 VTAIL.n58 B 0.013742f
C309 VTAIL.n59 B 0.025573f
C310 VTAIL.n60 B 0.025573f
C311 VTAIL.n61 B 0.013742f
C312 VTAIL.n62 B 0.01455f
C313 VTAIL.n63 B 0.032481f
C314 VTAIL.n64 B 0.032481f
C315 VTAIL.n65 B 0.01455f
C316 VTAIL.n66 B 0.013742f
C317 VTAIL.n67 B 0.025573f
C318 VTAIL.n68 B 0.025573f
C319 VTAIL.n69 B 0.013742f
C320 VTAIL.n70 B 0.01455f
C321 VTAIL.n71 B 0.032481f
C322 VTAIL.n72 B 0.032481f
C323 VTAIL.n73 B 0.032481f
C324 VTAIL.n74 B 0.01455f
C325 VTAIL.n75 B 0.013742f
C326 VTAIL.n76 B 0.025573f
C327 VTAIL.n77 B 0.025573f
C328 VTAIL.n78 B 0.013742f
C329 VTAIL.n79 B 0.014146f
C330 VTAIL.n80 B 0.014146f
C331 VTAIL.n81 B 0.032481f
C332 VTAIL.n82 B 0.032481f
C333 VTAIL.n83 B 0.01455f
C334 VTAIL.n84 B 0.013742f
C335 VTAIL.n85 B 0.025573f
C336 VTAIL.n86 B 0.025573f
C337 VTAIL.n87 B 0.013742f
C338 VTAIL.n88 B 0.01455f
C339 VTAIL.n89 B 0.032481f
C340 VTAIL.n90 B 0.068486f
C341 VTAIL.n91 B 0.01455f
C342 VTAIL.n92 B 0.013742f
C343 VTAIL.n93 B 0.05981f
C344 VTAIL.n94 B 0.038154f
C345 VTAIL.n95 B 0.164311f
C346 VTAIL.t5 B 0.339914f
C347 VTAIL.t18 B 0.339914f
C348 VTAIL.n96 B 3.01096f
C349 VTAIL.n97 B 0.391497f
C350 VTAIL.t19 B 0.339914f
C351 VTAIL.t2 B 0.339914f
C352 VTAIL.n98 B 3.01096f
C353 VTAIL.n99 B 2.00264f
C354 VTAIL.t13 B 0.339914f
C355 VTAIL.t7 B 0.339914f
C356 VTAIL.n100 B 3.01097f
C357 VTAIL.n101 B 2.00262f
C358 VTAIL.t11 B 0.339914f
C359 VTAIL.t15 B 0.339914f
C360 VTAIL.n102 B 3.01097f
C361 VTAIL.n103 B 0.391483f
C362 VTAIL.n104 B 0.034911f
C363 VTAIL.n105 B 0.025573f
C364 VTAIL.n106 B 0.013742f
C365 VTAIL.n107 B 0.032481f
C366 VTAIL.n108 B 0.01455f
C367 VTAIL.n109 B 0.025573f
C368 VTAIL.n110 B 0.013742f
C369 VTAIL.n111 B 0.032481f
C370 VTAIL.n112 B 0.01455f
C371 VTAIL.n113 B 0.025573f
C372 VTAIL.n114 B 0.013742f
C373 VTAIL.n115 B 0.032481f
C374 VTAIL.n116 B 0.032481f
C375 VTAIL.n117 B 0.01455f
C376 VTAIL.n118 B 0.025573f
C377 VTAIL.n119 B 0.013742f
C378 VTAIL.n120 B 0.032481f
C379 VTAIL.n121 B 0.01455f
C380 VTAIL.n122 B 0.025573f
C381 VTAIL.n123 B 0.013742f
C382 VTAIL.n124 B 0.032481f
C383 VTAIL.n125 B 0.01455f
C384 VTAIL.n126 B 0.025573f
C385 VTAIL.n127 B 0.013742f
C386 VTAIL.n128 B 0.032481f
C387 VTAIL.n129 B 0.01455f
C388 VTAIL.n130 B 0.025573f
C389 VTAIL.n131 B 0.013742f
C390 VTAIL.n132 B 0.032481f
C391 VTAIL.n133 B 0.01455f
C392 VTAIL.n134 B 0.178465f
C393 VTAIL.t9 B 0.053717f
C394 VTAIL.n135 B 0.024361f
C395 VTAIL.n136 B 0.019188f
C396 VTAIL.n137 B 0.013742f
C397 VTAIL.n138 B 1.87715f
C398 VTAIL.n139 B 0.025573f
C399 VTAIL.n140 B 0.013742f
C400 VTAIL.n141 B 0.01455f
C401 VTAIL.n142 B 0.032481f
C402 VTAIL.n143 B 0.032481f
C403 VTAIL.n144 B 0.01455f
C404 VTAIL.n145 B 0.013742f
C405 VTAIL.n146 B 0.025573f
C406 VTAIL.n147 B 0.025573f
C407 VTAIL.n148 B 0.013742f
C408 VTAIL.n149 B 0.01455f
C409 VTAIL.n150 B 0.032481f
C410 VTAIL.n151 B 0.032481f
C411 VTAIL.n152 B 0.01455f
C412 VTAIL.n153 B 0.013742f
C413 VTAIL.n154 B 0.025573f
C414 VTAIL.n155 B 0.025573f
C415 VTAIL.n156 B 0.013742f
C416 VTAIL.n157 B 0.01455f
C417 VTAIL.n158 B 0.032481f
C418 VTAIL.n159 B 0.032481f
C419 VTAIL.n160 B 0.01455f
C420 VTAIL.n161 B 0.013742f
C421 VTAIL.n162 B 0.025573f
C422 VTAIL.n163 B 0.025573f
C423 VTAIL.n164 B 0.013742f
C424 VTAIL.n165 B 0.01455f
C425 VTAIL.n166 B 0.032481f
C426 VTAIL.n167 B 0.032481f
C427 VTAIL.n168 B 0.01455f
C428 VTAIL.n169 B 0.013742f
C429 VTAIL.n170 B 0.025573f
C430 VTAIL.n171 B 0.025573f
C431 VTAIL.n172 B 0.013742f
C432 VTAIL.n173 B 0.01455f
C433 VTAIL.n174 B 0.032481f
C434 VTAIL.n175 B 0.032481f
C435 VTAIL.n176 B 0.01455f
C436 VTAIL.n177 B 0.013742f
C437 VTAIL.n178 B 0.025573f
C438 VTAIL.n179 B 0.025573f
C439 VTAIL.n180 B 0.013742f
C440 VTAIL.n181 B 0.014146f
C441 VTAIL.n182 B 0.014146f
C442 VTAIL.n183 B 0.032481f
C443 VTAIL.n184 B 0.032481f
C444 VTAIL.n185 B 0.01455f
C445 VTAIL.n186 B 0.013742f
C446 VTAIL.n187 B 0.025573f
C447 VTAIL.n188 B 0.025573f
C448 VTAIL.n189 B 0.013742f
C449 VTAIL.n190 B 0.01455f
C450 VTAIL.n191 B 0.032481f
C451 VTAIL.n192 B 0.068486f
C452 VTAIL.n193 B 0.01455f
C453 VTAIL.n194 B 0.013742f
C454 VTAIL.n195 B 0.05981f
C455 VTAIL.n196 B 0.038154f
C456 VTAIL.n197 B 0.164311f
C457 VTAIL.t1 B 0.339914f
C458 VTAIL.t4 B 0.339914f
C459 VTAIL.n198 B 3.01097f
C460 VTAIL.n199 B 0.395745f
C461 VTAIL.t0 B 0.339914f
C462 VTAIL.t3 B 0.339914f
C463 VTAIL.n200 B 3.01097f
C464 VTAIL.n201 B 0.391483f
C465 VTAIL.n202 B 0.034911f
C466 VTAIL.n203 B 0.025573f
C467 VTAIL.n204 B 0.013742f
C468 VTAIL.n205 B 0.032481f
C469 VTAIL.n206 B 0.01455f
C470 VTAIL.n207 B 0.025573f
C471 VTAIL.n208 B 0.013742f
C472 VTAIL.n209 B 0.032481f
C473 VTAIL.n210 B 0.01455f
C474 VTAIL.n211 B 0.025573f
C475 VTAIL.n212 B 0.013742f
C476 VTAIL.n213 B 0.032481f
C477 VTAIL.n214 B 0.032481f
C478 VTAIL.n215 B 0.01455f
C479 VTAIL.n216 B 0.025573f
C480 VTAIL.n217 B 0.013742f
C481 VTAIL.n218 B 0.032481f
C482 VTAIL.n219 B 0.01455f
C483 VTAIL.n220 B 0.025573f
C484 VTAIL.n221 B 0.013742f
C485 VTAIL.n222 B 0.032481f
C486 VTAIL.n223 B 0.01455f
C487 VTAIL.n224 B 0.025573f
C488 VTAIL.n225 B 0.013742f
C489 VTAIL.n226 B 0.032481f
C490 VTAIL.n227 B 0.01455f
C491 VTAIL.n228 B 0.025573f
C492 VTAIL.n229 B 0.013742f
C493 VTAIL.n230 B 0.032481f
C494 VTAIL.n231 B 0.01455f
C495 VTAIL.n232 B 0.178465f
C496 VTAIL.t17 B 0.053717f
C497 VTAIL.n233 B 0.024361f
C498 VTAIL.n234 B 0.019188f
C499 VTAIL.n235 B 0.013742f
C500 VTAIL.n236 B 1.87715f
C501 VTAIL.n237 B 0.025573f
C502 VTAIL.n238 B 0.013742f
C503 VTAIL.n239 B 0.01455f
C504 VTAIL.n240 B 0.032481f
C505 VTAIL.n241 B 0.032481f
C506 VTAIL.n242 B 0.01455f
C507 VTAIL.n243 B 0.013742f
C508 VTAIL.n244 B 0.025573f
C509 VTAIL.n245 B 0.025573f
C510 VTAIL.n246 B 0.013742f
C511 VTAIL.n247 B 0.01455f
C512 VTAIL.n248 B 0.032481f
C513 VTAIL.n249 B 0.032481f
C514 VTAIL.n250 B 0.01455f
C515 VTAIL.n251 B 0.013742f
C516 VTAIL.n252 B 0.025573f
C517 VTAIL.n253 B 0.025573f
C518 VTAIL.n254 B 0.013742f
C519 VTAIL.n255 B 0.01455f
C520 VTAIL.n256 B 0.032481f
C521 VTAIL.n257 B 0.032481f
C522 VTAIL.n258 B 0.01455f
C523 VTAIL.n259 B 0.013742f
C524 VTAIL.n260 B 0.025573f
C525 VTAIL.n261 B 0.025573f
C526 VTAIL.n262 B 0.013742f
C527 VTAIL.n263 B 0.01455f
C528 VTAIL.n264 B 0.032481f
C529 VTAIL.n265 B 0.032481f
C530 VTAIL.n266 B 0.01455f
C531 VTAIL.n267 B 0.013742f
C532 VTAIL.n268 B 0.025573f
C533 VTAIL.n269 B 0.025573f
C534 VTAIL.n270 B 0.013742f
C535 VTAIL.n271 B 0.01455f
C536 VTAIL.n272 B 0.032481f
C537 VTAIL.n273 B 0.032481f
C538 VTAIL.n274 B 0.01455f
C539 VTAIL.n275 B 0.013742f
C540 VTAIL.n276 B 0.025573f
C541 VTAIL.n277 B 0.025573f
C542 VTAIL.n278 B 0.013742f
C543 VTAIL.n279 B 0.014146f
C544 VTAIL.n280 B 0.014146f
C545 VTAIL.n281 B 0.032481f
C546 VTAIL.n282 B 0.032481f
C547 VTAIL.n283 B 0.01455f
C548 VTAIL.n284 B 0.013742f
C549 VTAIL.n285 B 0.025573f
C550 VTAIL.n286 B 0.025573f
C551 VTAIL.n287 B 0.013742f
C552 VTAIL.n288 B 0.01455f
C553 VTAIL.n289 B 0.032481f
C554 VTAIL.n290 B 0.068486f
C555 VTAIL.n291 B 0.01455f
C556 VTAIL.n292 B 0.013742f
C557 VTAIL.n293 B 0.05981f
C558 VTAIL.n294 B 0.038154f
C559 VTAIL.n295 B 1.70228f
C560 VTAIL.n296 B 0.034911f
C561 VTAIL.n297 B 0.025573f
C562 VTAIL.n298 B 0.013742f
C563 VTAIL.n299 B 0.032481f
C564 VTAIL.n300 B 0.01455f
C565 VTAIL.n301 B 0.025573f
C566 VTAIL.n302 B 0.013742f
C567 VTAIL.n303 B 0.032481f
C568 VTAIL.n304 B 0.01455f
C569 VTAIL.n305 B 0.025573f
C570 VTAIL.n306 B 0.013742f
C571 VTAIL.n307 B 0.032481f
C572 VTAIL.n308 B 0.01455f
C573 VTAIL.n309 B 0.025573f
C574 VTAIL.n310 B 0.013742f
C575 VTAIL.n311 B 0.032481f
C576 VTAIL.n312 B 0.01455f
C577 VTAIL.n313 B 0.025573f
C578 VTAIL.n314 B 0.013742f
C579 VTAIL.n315 B 0.032481f
C580 VTAIL.n316 B 0.01455f
C581 VTAIL.n317 B 0.025573f
C582 VTAIL.n318 B 0.013742f
C583 VTAIL.n319 B 0.032481f
C584 VTAIL.n320 B 0.01455f
C585 VTAIL.n321 B 0.025573f
C586 VTAIL.n322 B 0.013742f
C587 VTAIL.n323 B 0.032481f
C588 VTAIL.n324 B 0.01455f
C589 VTAIL.n325 B 0.178465f
C590 VTAIL.t6 B 0.053717f
C591 VTAIL.n326 B 0.024361f
C592 VTAIL.n327 B 0.019188f
C593 VTAIL.n328 B 0.013742f
C594 VTAIL.n329 B 1.87715f
C595 VTAIL.n330 B 0.025573f
C596 VTAIL.n331 B 0.013742f
C597 VTAIL.n332 B 0.01455f
C598 VTAIL.n333 B 0.032481f
C599 VTAIL.n334 B 0.032481f
C600 VTAIL.n335 B 0.01455f
C601 VTAIL.n336 B 0.013742f
C602 VTAIL.n337 B 0.025573f
C603 VTAIL.n338 B 0.025573f
C604 VTAIL.n339 B 0.013742f
C605 VTAIL.n340 B 0.01455f
C606 VTAIL.n341 B 0.032481f
C607 VTAIL.n342 B 0.032481f
C608 VTAIL.n343 B 0.01455f
C609 VTAIL.n344 B 0.013742f
C610 VTAIL.n345 B 0.025573f
C611 VTAIL.n346 B 0.025573f
C612 VTAIL.n347 B 0.013742f
C613 VTAIL.n348 B 0.01455f
C614 VTAIL.n349 B 0.032481f
C615 VTAIL.n350 B 0.032481f
C616 VTAIL.n351 B 0.01455f
C617 VTAIL.n352 B 0.013742f
C618 VTAIL.n353 B 0.025573f
C619 VTAIL.n354 B 0.025573f
C620 VTAIL.n355 B 0.013742f
C621 VTAIL.n356 B 0.01455f
C622 VTAIL.n357 B 0.032481f
C623 VTAIL.n358 B 0.032481f
C624 VTAIL.n359 B 0.01455f
C625 VTAIL.n360 B 0.013742f
C626 VTAIL.n361 B 0.025573f
C627 VTAIL.n362 B 0.025573f
C628 VTAIL.n363 B 0.013742f
C629 VTAIL.n364 B 0.01455f
C630 VTAIL.n365 B 0.032481f
C631 VTAIL.n366 B 0.032481f
C632 VTAIL.n367 B 0.032481f
C633 VTAIL.n368 B 0.01455f
C634 VTAIL.n369 B 0.013742f
C635 VTAIL.n370 B 0.025573f
C636 VTAIL.n371 B 0.025573f
C637 VTAIL.n372 B 0.013742f
C638 VTAIL.n373 B 0.014146f
C639 VTAIL.n374 B 0.014146f
C640 VTAIL.n375 B 0.032481f
C641 VTAIL.n376 B 0.032481f
C642 VTAIL.n377 B 0.01455f
C643 VTAIL.n378 B 0.013742f
C644 VTAIL.n379 B 0.025573f
C645 VTAIL.n380 B 0.025573f
C646 VTAIL.n381 B 0.013742f
C647 VTAIL.n382 B 0.01455f
C648 VTAIL.n383 B 0.032481f
C649 VTAIL.n384 B 0.068486f
C650 VTAIL.n385 B 0.01455f
C651 VTAIL.n386 B 0.013742f
C652 VTAIL.n387 B 0.05981f
C653 VTAIL.n388 B 0.038154f
C654 VTAIL.n389 B 1.70228f
C655 VTAIL.t10 B 0.339914f
C656 VTAIL.t12 B 0.339914f
C657 VTAIL.n390 B 3.01096f
C658 VTAIL.n391 B 0.335023f
C659 VDD2.n0 B 0.034015f
C660 VDD2.n1 B 0.024917f
C661 VDD2.n2 B 0.013389f
C662 VDD2.n3 B 0.031648f
C663 VDD2.n4 B 0.014177f
C664 VDD2.n5 B 0.024917f
C665 VDD2.n6 B 0.013389f
C666 VDD2.n7 B 0.031648f
C667 VDD2.n8 B 0.014177f
C668 VDD2.n9 B 0.024917f
C669 VDD2.n10 B 0.013389f
C670 VDD2.n11 B 0.031648f
C671 VDD2.n12 B 0.014177f
C672 VDD2.n13 B 0.024917f
C673 VDD2.n14 B 0.013389f
C674 VDD2.n15 B 0.031648f
C675 VDD2.n16 B 0.014177f
C676 VDD2.n17 B 0.024917f
C677 VDD2.n18 B 0.013389f
C678 VDD2.n19 B 0.031648f
C679 VDD2.n20 B 0.014177f
C680 VDD2.n21 B 0.024917f
C681 VDD2.n22 B 0.013389f
C682 VDD2.n23 B 0.031648f
C683 VDD2.n24 B 0.014177f
C684 VDD2.n25 B 0.024917f
C685 VDD2.n26 B 0.013389f
C686 VDD2.n27 B 0.031648f
C687 VDD2.n28 B 0.014177f
C688 VDD2.n29 B 0.173886f
C689 VDD2.t6 B 0.052339f
C690 VDD2.n30 B 0.023736f
C691 VDD2.n31 B 0.018695f
C692 VDD2.n32 B 0.013389f
C693 VDD2.n33 B 1.82899f
C694 VDD2.n34 B 0.024917f
C695 VDD2.n35 B 0.013389f
C696 VDD2.n36 B 0.014177f
C697 VDD2.n37 B 0.031648f
C698 VDD2.n38 B 0.031648f
C699 VDD2.n39 B 0.014177f
C700 VDD2.n40 B 0.013389f
C701 VDD2.n41 B 0.024917f
C702 VDD2.n42 B 0.024917f
C703 VDD2.n43 B 0.013389f
C704 VDD2.n44 B 0.014177f
C705 VDD2.n45 B 0.031648f
C706 VDD2.n46 B 0.031648f
C707 VDD2.n47 B 0.014177f
C708 VDD2.n48 B 0.013389f
C709 VDD2.n49 B 0.024917f
C710 VDD2.n50 B 0.024917f
C711 VDD2.n51 B 0.013389f
C712 VDD2.n52 B 0.014177f
C713 VDD2.n53 B 0.031648f
C714 VDD2.n54 B 0.031648f
C715 VDD2.n55 B 0.014177f
C716 VDD2.n56 B 0.013389f
C717 VDD2.n57 B 0.024917f
C718 VDD2.n58 B 0.024917f
C719 VDD2.n59 B 0.013389f
C720 VDD2.n60 B 0.014177f
C721 VDD2.n61 B 0.031648f
C722 VDD2.n62 B 0.031648f
C723 VDD2.n63 B 0.014177f
C724 VDD2.n64 B 0.013389f
C725 VDD2.n65 B 0.024917f
C726 VDD2.n66 B 0.024917f
C727 VDD2.n67 B 0.013389f
C728 VDD2.n68 B 0.014177f
C729 VDD2.n69 B 0.031648f
C730 VDD2.n70 B 0.031648f
C731 VDD2.n71 B 0.031648f
C732 VDD2.n72 B 0.014177f
C733 VDD2.n73 B 0.013389f
C734 VDD2.n74 B 0.024917f
C735 VDD2.n75 B 0.024917f
C736 VDD2.n76 B 0.013389f
C737 VDD2.n77 B 0.013783f
C738 VDD2.n78 B 0.013783f
C739 VDD2.n79 B 0.031648f
C740 VDD2.n80 B 0.031648f
C741 VDD2.n81 B 0.014177f
C742 VDD2.n82 B 0.013389f
C743 VDD2.n83 B 0.024917f
C744 VDD2.n84 B 0.024917f
C745 VDD2.n85 B 0.013389f
C746 VDD2.n86 B 0.014177f
C747 VDD2.n87 B 0.031648f
C748 VDD2.n88 B 0.066728f
C749 VDD2.n89 B 0.014177f
C750 VDD2.n90 B 0.013389f
C751 VDD2.n91 B 0.058276f
C752 VDD2.n92 B 0.056302f
C753 VDD2.t0 B 0.331192f
C754 VDD2.t2 B 0.331192f
C755 VDD2.n93 B 3.00911f
C756 VDD2.n94 B 0.402452f
C757 VDD2.t8 B 0.331192f
C758 VDD2.t4 B 0.331192f
C759 VDD2.n95 B 3.01216f
C760 VDD2.n96 B 2.16155f
C761 VDD2.n97 B 0.034015f
C762 VDD2.n98 B 0.024917f
C763 VDD2.n99 B 0.013389f
C764 VDD2.n100 B 0.031648f
C765 VDD2.n101 B 0.014177f
C766 VDD2.n102 B 0.024917f
C767 VDD2.n103 B 0.013389f
C768 VDD2.n104 B 0.031648f
C769 VDD2.n105 B 0.014177f
C770 VDD2.n106 B 0.024917f
C771 VDD2.n107 B 0.013389f
C772 VDD2.n108 B 0.031648f
C773 VDD2.n109 B 0.031648f
C774 VDD2.n110 B 0.014177f
C775 VDD2.n111 B 0.024917f
C776 VDD2.n112 B 0.013389f
C777 VDD2.n113 B 0.031648f
C778 VDD2.n114 B 0.014177f
C779 VDD2.n115 B 0.024917f
C780 VDD2.n116 B 0.013389f
C781 VDD2.n117 B 0.031648f
C782 VDD2.n118 B 0.014177f
C783 VDD2.n119 B 0.024917f
C784 VDD2.n120 B 0.013389f
C785 VDD2.n121 B 0.031648f
C786 VDD2.n122 B 0.014177f
C787 VDD2.n123 B 0.024917f
C788 VDD2.n124 B 0.013389f
C789 VDD2.n125 B 0.031648f
C790 VDD2.n126 B 0.014177f
C791 VDD2.n127 B 0.173886f
C792 VDD2.t9 B 0.052339f
C793 VDD2.n128 B 0.023736f
C794 VDD2.n129 B 0.018695f
C795 VDD2.n130 B 0.013389f
C796 VDD2.n131 B 1.82899f
C797 VDD2.n132 B 0.024917f
C798 VDD2.n133 B 0.013389f
C799 VDD2.n134 B 0.014177f
C800 VDD2.n135 B 0.031648f
C801 VDD2.n136 B 0.031648f
C802 VDD2.n137 B 0.014177f
C803 VDD2.n138 B 0.013389f
C804 VDD2.n139 B 0.024917f
C805 VDD2.n140 B 0.024917f
C806 VDD2.n141 B 0.013389f
C807 VDD2.n142 B 0.014177f
C808 VDD2.n143 B 0.031648f
C809 VDD2.n144 B 0.031648f
C810 VDD2.n145 B 0.014177f
C811 VDD2.n146 B 0.013389f
C812 VDD2.n147 B 0.024917f
C813 VDD2.n148 B 0.024917f
C814 VDD2.n149 B 0.013389f
C815 VDD2.n150 B 0.014177f
C816 VDD2.n151 B 0.031648f
C817 VDD2.n152 B 0.031648f
C818 VDD2.n153 B 0.014177f
C819 VDD2.n154 B 0.013389f
C820 VDD2.n155 B 0.024917f
C821 VDD2.n156 B 0.024917f
C822 VDD2.n157 B 0.013389f
C823 VDD2.n158 B 0.014177f
C824 VDD2.n159 B 0.031648f
C825 VDD2.n160 B 0.031648f
C826 VDD2.n161 B 0.014177f
C827 VDD2.n162 B 0.013389f
C828 VDD2.n163 B 0.024917f
C829 VDD2.n164 B 0.024917f
C830 VDD2.n165 B 0.013389f
C831 VDD2.n166 B 0.014177f
C832 VDD2.n167 B 0.031648f
C833 VDD2.n168 B 0.031648f
C834 VDD2.n169 B 0.014177f
C835 VDD2.n170 B 0.013389f
C836 VDD2.n171 B 0.024917f
C837 VDD2.n172 B 0.024917f
C838 VDD2.n173 B 0.013389f
C839 VDD2.n174 B 0.013783f
C840 VDD2.n175 B 0.013783f
C841 VDD2.n176 B 0.031648f
C842 VDD2.n177 B 0.031648f
C843 VDD2.n178 B 0.014177f
C844 VDD2.n179 B 0.013389f
C845 VDD2.n180 B 0.024917f
C846 VDD2.n181 B 0.024917f
C847 VDD2.n182 B 0.013389f
C848 VDD2.n183 B 0.014177f
C849 VDD2.n184 B 0.031648f
C850 VDD2.n185 B 0.066728f
C851 VDD2.n186 B 0.014177f
C852 VDD2.n187 B 0.013389f
C853 VDD2.n188 B 0.058276f
C854 VDD2.n189 B 0.054374f
C855 VDD2.n190 B 2.49588f
C856 VDD2.t5 B 0.331192f
C857 VDD2.t3 B 0.331192f
C858 VDD2.n191 B 3.00912f
C859 VDD2.n192 B 0.29422f
C860 VDD2.t7 B 0.331192f
C861 VDD2.t1 B 0.331192f
C862 VDD2.n193 B 3.01214f
C863 VN.n0 B 0.073277f
C864 VN.t7 B 1.34378f
C865 VN.n1 B 0.522602f
C866 VN.t1 B 1.36284f
C867 VN.n2 B 0.494914f
C868 VN.n3 B 0.232721f
C869 VN.t5 B 1.34378f
C870 VN.n4 B 0.522602f
C871 VN.t3 B 1.34378f
C872 VN.n5 B 0.522602f
C873 VN.t9 B 1.34378f
C874 VN.n6 B 0.512619f
C875 VN.n7 B 0.048804f
C876 VN.n8 B 0.073277f
C877 VN.t0 B 1.34378f
C878 VN.n9 B 0.522602f
C879 VN.t4 B 1.34378f
C880 VN.t6 B 1.36284f
C881 VN.n10 B 0.494914f
C882 VN.n11 B 0.232721f
C883 VN.n12 B 0.522602f
C884 VN.t8 B 1.34378f
C885 VN.n13 B 0.522602f
C886 VN.t2 B 1.34378f
C887 VN.n14 B 0.512619f
C888 VN.n15 B 2.16133f
.ends

