* NGSPICE file created from diff_pair_sample_1642.ext - technology: sky130A

.subckt diff_pair_sample_1642 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=2.78355 ps=17.2 w=16.87 l=2.22
X1 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X2 VTAIL.t17 VP.t1 VDD1.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X3 VTAIL.t18 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X4 VDD2.t8 VN.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=2.78355 ps=17.2 w=16.87 l=2.22
X5 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X6 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X7 VDD1.t6 VP.t3 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=2.78355 ps=17.2 w=16.87 l=2.22
X8 VDD1.t5 VP.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=6.5793 ps=34.52 w=16.87 l=2.22
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=0 ps=0 w=16.87 l=2.22
X10 VTAIL.t1 VN.t4 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X11 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=2.78355 ps=17.2 w=16.87 l=2.22
X12 VTAIL.t3 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X13 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=0 ps=0 w=16.87 l=2.22
X14 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=6.5793 ps=34.52 w=16.87 l=2.22
X15 VDD2.t1 VN.t8 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=6.5793 ps=34.52 w=16.87 l=2.22
X16 VTAIL.t14 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X17 VDD1.t3 VP.t6 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=0 ps=0 w=16.87 l=2.22
X19 VTAIL.t12 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X20 VDD1.t1 VP.t8 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X21 VTAIL.t7 VN.t9 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=2.78355 ps=17.2 w=16.87 l=2.22
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5793 pd=34.52 as=0 ps=0 w=16.87 l=2.22
X23 VDD1.t0 VP.t9 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.78355 pd=17.2 as=6.5793 ps=34.52 w=16.87 l=2.22
R0 VP.n19 VP.t0 216.532
R1 VP.n48 VP.t3 183.138
R2 VP.n56 VP.t1 183.138
R3 VP.n5 VP.t8 183.138
R4 VP.n73 VP.t7 183.138
R5 VP.n81 VP.t4 183.138
R6 VP.n45 VP.t9 183.138
R7 VP.n37 VP.t5 183.138
R8 VP.n16 VP.t6 183.138
R9 VP.n20 VP.t2 183.138
R10 VP.n22 VP.n21 161.3
R11 VP.n23 VP.n18 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n26 VP.n17 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n30 VP.n29 161.3
R16 VP.n31 VP.n15 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n34 VP.n14 161.3
R19 VP.n36 VP.n35 161.3
R20 VP.n38 VP.n13 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n41 VP.n12 161.3
R23 VP.n43 VP.n42 161.3
R24 VP.n44 VP.n11 161.3
R25 VP.n80 VP.n0 161.3
R26 VP.n79 VP.n78 161.3
R27 VP.n77 VP.n1 161.3
R28 VP.n76 VP.n75 161.3
R29 VP.n74 VP.n2 161.3
R30 VP.n72 VP.n71 161.3
R31 VP.n70 VP.n3 161.3
R32 VP.n69 VP.n68 161.3
R33 VP.n67 VP.n4 161.3
R34 VP.n66 VP.n65 161.3
R35 VP.n64 VP.n63 161.3
R36 VP.n62 VP.n6 161.3
R37 VP.n61 VP.n60 161.3
R38 VP.n59 VP.n7 161.3
R39 VP.n58 VP.n57 161.3
R40 VP.n55 VP.n8 161.3
R41 VP.n54 VP.n53 161.3
R42 VP.n52 VP.n9 161.3
R43 VP.n51 VP.n50 161.3
R44 VP.n49 VP.n10 161.3
R45 VP.n48 VP.n47 93.6295
R46 VP.n82 VP.n81 93.6295
R47 VP.n46 VP.n45 93.6295
R48 VP.n20 VP.n19 56.5548
R49 VP.n47 VP.n46 54.7761
R50 VP.n50 VP.n9 47.7779
R51 VP.n79 VP.n1 47.7779
R52 VP.n43 VP.n12 47.7779
R53 VP.n61 VP.n7 42.9216
R54 VP.n68 VP.n3 42.9216
R55 VP.n32 VP.n14 42.9216
R56 VP.n25 VP.n18 42.9216
R57 VP.n62 VP.n61 38.0652
R58 VP.n68 VP.n67 38.0652
R59 VP.n32 VP.n31 38.0652
R60 VP.n26 VP.n25 38.0652
R61 VP.n54 VP.n9 33.2089
R62 VP.n75 VP.n1 33.2089
R63 VP.n39 VP.n12 33.2089
R64 VP.n50 VP.n49 24.4675
R65 VP.n55 VP.n54 24.4675
R66 VP.n57 VP.n7 24.4675
R67 VP.n63 VP.n62 24.4675
R68 VP.n67 VP.n66 24.4675
R69 VP.n72 VP.n3 24.4675
R70 VP.n75 VP.n74 24.4675
R71 VP.n80 VP.n79 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n36 VP.n14 24.4675
R74 VP.n39 VP.n38 24.4675
R75 VP.n27 VP.n26 24.4675
R76 VP.n31 VP.n30 24.4675
R77 VP.n21 VP.n18 24.4675
R78 VP.n49 VP.n48 17.1274
R79 VP.n81 VP.n80 17.1274
R80 VP.n45 VP.n44 17.1274
R81 VP.n57 VP.n56 14.6807
R82 VP.n73 VP.n72 14.6807
R83 VP.n37 VP.n36 14.6807
R84 VP.n21 VP.n20 14.6807
R85 VP.n63 VP.n5 12.234
R86 VP.n66 VP.n5 12.234
R87 VP.n27 VP.n16 12.234
R88 VP.n30 VP.n16 12.234
R89 VP.n56 VP.n55 9.7873
R90 VP.n74 VP.n73 9.7873
R91 VP.n38 VP.n37 9.7873
R92 VP.n22 VP.n19 9.24318
R93 VP.n46 VP.n11 0.278367
R94 VP.n47 VP.n10 0.278367
R95 VP.n82 VP.n0 0.278367
R96 VP.n23 VP.n22 0.189894
R97 VP.n24 VP.n23 0.189894
R98 VP.n24 VP.n17 0.189894
R99 VP.n28 VP.n17 0.189894
R100 VP.n29 VP.n28 0.189894
R101 VP.n29 VP.n15 0.189894
R102 VP.n33 VP.n15 0.189894
R103 VP.n34 VP.n33 0.189894
R104 VP.n35 VP.n34 0.189894
R105 VP.n35 VP.n13 0.189894
R106 VP.n40 VP.n13 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n11 0.189894
R110 VP.n51 VP.n10 0.189894
R111 VP.n52 VP.n51 0.189894
R112 VP.n53 VP.n52 0.189894
R113 VP.n53 VP.n8 0.189894
R114 VP.n58 VP.n8 0.189894
R115 VP.n59 VP.n58 0.189894
R116 VP.n60 VP.n59 0.189894
R117 VP.n60 VP.n6 0.189894
R118 VP.n64 VP.n6 0.189894
R119 VP.n65 VP.n64 0.189894
R120 VP.n65 VP.n4 0.189894
R121 VP.n69 VP.n4 0.189894
R122 VP.n70 VP.n69 0.189894
R123 VP.n71 VP.n70 0.189894
R124 VP.n71 VP.n2 0.189894
R125 VP.n76 VP.n2 0.189894
R126 VP.n77 VP.n76 0.189894
R127 VP.n78 VP.n77 0.189894
R128 VP.n78 VP.n0 0.189894
R129 VP VP.n82 0.153454
R130 VTAIL.n384 VTAIL.n296 289.615
R131 VTAIL.n90 VTAIL.n2 289.615
R132 VTAIL.n290 VTAIL.n202 289.615
R133 VTAIL.n192 VTAIL.n104 289.615
R134 VTAIL.n327 VTAIL.n326 185
R135 VTAIL.n324 VTAIL.n323 185
R136 VTAIL.n333 VTAIL.n332 185
R137 VTAIL.n335 VTAIL.n334 185
R138 VTAIL.n320 VTAIL.n319 185
R139 VTAIL.n341 VTAIL.n340 185
R140 VTAIL.n343 VTAIL.n342 185
R141 VTAIL.n316 VTAIL.n315 185
R142 VTAIL.n349 VTAIL.n348 185
R143 VTAIL.n351 VTAIL.n350 185
R144 VTAIL.n312 VTAIL.n311 185
R145 VTAIL.n357 VTAIL.n356 185
R146 VTAIL.n359 VTAIL.n358 185
R147 VTAIL.n308 VTAIL.n307 185
R148 VTAIL.n365 VTAIL.n364 185
R149 VTAIL.n368 VTAIL.n367 185
R150 VTAIL.n366 VTAIL.n304 185
R151 VTAIL.n373 VTAIL.n303 185
R152 VTAIL.n375 VTAIL.n374 185
R153 VTAIL.n377 VTAIL.n376 185
R154 VTAIL.n300 VTAIL.n299 185
R155 VTAIL.n383 VTAIL.n382 185
R156 VTAIL.n385 VTAIL.n384 185
R157 VTAIL.n33 VTAIL.n32 185
R158 VTAIL.n30 VTAIL.n29 185
R159 VTAIL.n39 VTAIL.n38 185
R160 VTAIL.n41 VTAIL.n40 185
R161 VTAIL.n26 VTAIL.n25 185
R162 VTAIL.n47 VTAIL.n46 185
R163 VTAIL.n49 VTAIL.n48 185
R164 VTAIL.n22 VTAIL.n21 185
R165 VTAIL.n55 VTAIL.n54 185
R166 VTAIL.n57 VTAIL.n56 185
R167 VTAIL.n18 VTAIL.n17 185
R168 VTAIL.n63 VTAIL.n62 185
R169 VTAIL.n65 VTAIL.n64 185
R170 VTAIL.n14 VTAIL.n13 185
R171 VTAIL.n71 VTAIL.n70 185
R172 VTAIL.n74 VTAIL.n73 185
R173 VTAIL.n72 VTAIL.n10 185
R174 VTAIL.n79 VTAIL.n9 185
R175 VTAIL.n81 VTAIL.n80 185
R176 VTAIL.n83 VTAIL.n82 185
R177 VTAIL.n6 VTAIL.n5 185
R178 VTAIL.n89 VTAIL.n88 185
R179 VTAIL.n91 VTAIL.n90 185
R180 VTAIL.n291 VTAIL.n290 185
R181 VTAIL.n289 VTAIL.n288 185
R182 VTAIL.n206 VTAIL.n205 185
R183 VTAIL.n283 VTAIL.n282 185
R184 VTAIL.n281 VTAIL.n280 185
R185 VTAIL.n279 VTAIL.n209 185
R186 VTAIL.n213 VTAIL.n210 185
R187 VTAIL.n274 VTAIL.n273 185
R188 VTAIL.n272 VTAIL.n271 185
R189 VTAIL.n215 VTAIL.n214 185
R190 VTAIL.n266 VTAIL.n265 185
R191 VTAIL.n264 VTAIL.n263 185
R192 VTAIL.n219 VTAIL.n218 185
R193 VTAIL.n258 VTAIL.n257 185
R194 VTAIL.n256 VTAIL.n255 185
R195 VTAIL.n223 VTAIL.n222 185
R196 VTAIL.n250 VTAIL.n249 185
R197 VTAIL.n248 VTAIL.n247 185
R198 VTAIL.n227 VTAIL.n226 185
R199 VTAIL.n242 VTAIL.n241 185
R200 VTAIL.n240 VTAIL.n239 185
R201 VTAIL.n231 VTAIL.n230 185
R202 VTAIL.n234 VTAIL.n233 185
R203 VTAIL.n193 VTAIL.n192 185
R204 VTAIL.n191 VTAIL.n190 185
R205 VTAIL.n108 VTAIL.n107 185
R206 VTAIL.n185 VTAIL.n184 185
R207 VTAIL.n183 VTAIL.n182 185
R208 VTAIL.n181 VTAIL.n111 185
R209 VTAIL.n115 VTAIL.n112 185
R210 VTAIL.n176 VTAIL.n175 185
R211 VTAIL.n174 VTAIL.n173 185
R212 VTAIL.n117 VTAIL.n116 185
R213 VTAIL.n168 VTAIL.n167 185
R214 VTAIL.n166 VTAIL.n165 185
R215 VTAIL.n121 VTAIL.n120 185
R216 VTAIL.n160 VTAIL.n159 185
R217 VTAIL.n158 VTAIL.n157 185
R218 VTAIL.n125 VTAIL.n124 185
R219 VTAIL.n152 VTAIL.n151 185
R220 VTAIL.n150 VTAIL.n149 185
R221 VTAIL.n129 VTAIL.n128 185
R222 VTAIL.n144 VTAIL.n143 185
R223 VTAIL.n142 VTAIL.n141 185
R224 VTAIL.n133 VTAIL.n132 185
R225 VTAIL.n136 VTAIL.n135 185
R226 VTAIL.t13 VTAIL.n232 147.659
R227 VTAIL.t19 VTAIL.n134 147.659
R228 VTAIL.t5 VTAIL.n325 147.659
R229 VTAIL.t15 VTAIL.n31 147.659
R230 VTAIL.n326 VTAIL.n323 104.615
R231 VTAIL.n333 VTAIL.n323 104.615
R232 VTAIL.n334 VTAIL.n333 104.615
R233 VTAIL.n334 VTAIL.n319 104.615
R234 VTAIL.n341 VTAIL.n319 104.615
R235 VTAIL.n342 VTAIL.n341 104.615
R236 VTAIL.n342 VTAIL.n315 104.615
R237 VTAIL.n349 VTAIL.n315 104.615
R238 VTAIL.n350 VTAIL.n349 104.615
R239 VTAIL.n350 VTAIL.n311 104.615
R240 VTAIL.n357 VTAIL.n311 104.615
R241 VTAIL.n358 VTAIL.n357 104.615
R242 VTAIL.n358 VTAIL.n307 104.615
R243 VTAIL.n365 VTAIL.n307 104.615
R244 VTAIL.n367 VTAIL.n365 104.615
R245 VTAIL.n367 VTAIL.n366 104.615
R246 VTAIL.n366 VTAIL.n303 104.615
R247 VTAIL.n375 VTAIL.n303 104.615
R248 VTAIL.n376 VTAIL.n375 104.615
R249 VTAIL.n376 VTAIL.n299 104.615
R250 VTAIL.n383 VTAIL.n299 104.615
R251 VTAIL.n384 VTAIL.n383 104.615
R252 VTAIL.n32 VTAIL.n29 104.615
R253 VTAIL.n39 VTAIL.n29 104.615
R254 VTAIL.n40 VTAIL.n39 104.615
R255 VTAIL.n40 VTAIL.n25 104.615
R256 VTAIL.n47 VTAIL.n25 104.615
R257 VTAIL.n48 VTAIL.n47 104.615
R258 VTAIL.n48 VTAIL.n21 104.615
R259 VTAIL.n55 VTAIL.n21 104.615
R260 VTAIL.n56 VTAIL.n55 104.615
R261 VTAIL.n56 VTAIL.n17 104.615
R262 VTAIL.n63 VTAIL.n17 104.615
R263 VTAIL.n64 VTAIL.n63 104.615
R264 VTAIL.n64 VTAIL.n13 104.615
R265 VTAIL.n71 VTAIL.n13 104.615
R266 VTAIL.n73 VTAIL.n71 104.615
R267 VTAIL.n73 VTAIL.n72 104.615
R268 VTAIL.n72 VTAIL.n9 104.615
R269 VTAIL.n81 VTAIL.n9 104.615
R270 VTAIL.n82 VTAIL.n81 104.615
R271 VTAIL.n82 VTAIL.n5 104.615
R272 VTAIL.n89 VTAIL.n5 104.615
R273 VTAIL.n90 VTAIL.n89 104.615
R274 VTAIL.n290 VTAIL.n289 104.615
R275 VTAIL.n289 VTAIL.n205 104.615
R276 VTAIL.n282 VTAIL.n205 104.615
R277 VTAIL.n282 VTAIL.n281 104.615
R278 VTAIL.n281 VTAIL.n209 104.615
R279 VTAIL.n213 VTAIL.n209 104.615
R280 VTAIL.n273 VTAIL.n213 104.615
R281 VTAIL.n273 VTAIL.n272 104.615
R282 VTAIL.n272 VTAIL.n214 104.615
R283 VTAIL.n265 VTAIL.n214 104.615
R284 VTAIL.n265 VTAIL.n264 104.615
R285 VTAIL.n264 VTAIL.n218 104.615
R286 VTAIL.n257 VTAIL.n218 104.615
R287 VTAIL.n257 VTAIL.n256 104.615
R288 VTAIL.n256 VTAIL.n222 104.615
R289 VTAIL.n249 VTAIL.n222 104.615
R290 VTAIL.n249 VTAIL.n248 104.615
R291 VTAIL.n248 VTAIL.n226 104.615
R292 VTAIL.n241 VTAIL.n226 104.615
R293 VTAIL.n241 VTAIL.n240 104.615
R294 VTAIL.n240 VTAIL.n230 104.615
R295 VTAIL.n233 VTAIL.n230 104.615
R296 VTAIL.n192 VTAIL.n191 104.615
R297 VTAIL.n191 VTAIL.n107 104.615
R298 VTAIL.n184 VTAIL.n107 104.615
R299 VTAIL.n184 VTAIL.n183 104.615
R300 VTAIL.n183 VTAIL.n111 104.615
R301 VTAIL.n115 VTAIL.n111 104.615
R302 VTAIL.n175 VTAIL.n115 104.615
R303 VTAIL.n175 VTAIL.n174 104.615
R304 VTAIL.n174 VTAIL.n116 104.615
R305 VTAIL.n167 VTAIL.n116 104.615
R306 VTAIL.n167 VTAIL.n166 104.615
R307 VTAIL.n166 VTAIL.n120 104.615
R308 VTAIL.n159 VTAIL.n120 104.615
R309 VTAIL.n159 VTAIL.n158 104.615
R310 VTAIL.n158 VTAIL.n124 104.615
R311 VTAIL.n151 VTAIL.n124 104.615
R312 VTAIL.n151 VTAIL.n150 104.615
R313 VTAIL.n150 VTAIL.n128 104.615
R314 VTAIL.n143 VTAIL.n128 104.615
R315 VTAIL.n143 VTAIL.n142 104.615
R316 VTAIL.n142 VTAIL.n132 104.615
R317 VTAIL.n135 VTAIL.n132 104.615
R318 VTAIL.n326 VTAIL.t5 52.3082
R319 VTAIL.n32 VTAIL.t15 52.3082
R320 VTAIL.n233 VTAIL.t13 52.3082
R321 VTAIL.n135 VTAIL.t19 52.3082
R322 VTAIL.n201 VTAIL.n200 45.4036
R323 VTAIL.n199 VTAIL.n198 45.4036
R324 VTAIL.n103 VTAIL.n102 45.4036
R325 VTAIL.n101 VTAIL.n100 45.4036
R326 VTAIL.n391 VTAIL.n390 45.4034
R327 VTAIL.n1 VTAIL.n0 45.4034
R328 VTAIL.n97 VTAIL.n96 45.4034
R329 VTAIL.n99 VTAIL.n98 45.4034
R330 VTAIL.n389 VTAIL.n388 33.5429
R331 VTAIL.n95 VTAIL.n94 33.5429
R332 VTAIL.n295 VTAIL.n294 33.5429
R333 VTAIL.n197 VTAIL.n196 33.5429
R334 VTAIL.n101 VTAIL.n99 31.3065
R335 VTAIL.n389 VTAIL.n295 29.1083
R336 VTAIL.n327 VTAIL.n325 15.6677
R337 VTAIL.n33 VTAIL.n31 15.6677
R338 VTAIL.n234 VTAIL.n232 15.6677
R339 VTAIL.n136 VTAIL.n134 15.6677
R340 VTAIL.n374 VTAIL.n373 13.1884
R341 VTAIL.n80 VTAIL.n79 13.1884
R342 VTAIL.n280 VTAIL.n279 13.1884
R343 VTAIL.n182 VTAIL.n181 13.1884
R344 VTAIL.n328 VTAIL.n324 12.8005
R345 VTAIL.n372 VTAIL.n304 12.8005
R346 VTAIL.n377 VTAIL.n302 12.8005
R347 VTAIL.n34 VTAIL.n30 12.8005
R348 VTAIL.n78 VTAIL.n10 12.8005
R349 VTAIL.n83 VTAIL.n8 12.8005
R350 VTAIL.n283 VTAIL.n208 12.8005
R351 VTAIL.n278 VTAIL.n210 12.8005
R352 VTAIL.n235 VTAIL.n231 12.8005
R353 VTAIL.n185 VTAIL.n110 12.8005
R354 VTAIL.n180 VTAIL.n112 12.8005
R355 VTAIL.n137 VTAIL.n133 12.8005
R356 VTAIL.n332 VTAIL.n331 12.0247
R357 VTAIL.n369 VTAIL.n368 12.0247
R358 VTAIL.n378 VTAIL.n300 12.0247
R359 VTAIL.n38 VTAIL.n37 12.0247
R360 VTAIL.n75 VTAIL.n74 12.0247
R361 VTAIL.n84 VTAIL.n6 12.0247
R362 VTAIL.n284 VTAIL.n206 12.0247
R363 VTAIL.n275 VTAIL.n274 12.0247
R364 VTAIL.n239 VTAIL.n238 12.0247
R365 VTAIL.n186 VTAIL.n108 12.0247
R366 VTAIL.n177 VTAIL.n176 12.0247
R367 VTAIL.n141 VTAIL.n140 12.0247
R368 VTAIL.n335 VTAIL.n322 11.249
R369 VTAIL.n364 VTAIL.n306 11.249
R370 VTAIL.n382 VTAIL.n381 11.249
R371 VTAIL.n41 VTAIL.n28 11.249
R372 VTAIL.n70 VTAIL.n12 11.249
R373 VTAIL.n88 VTAIL.n87 11.249
R374 VTAIL.n288 VTAIL.n287 11.249
R375 VTAIL.n271 VTAIL.n212 11.249
R376 VTAIL.n242 VTAIL.n229 11.249
R377 VTAIL.n190 VTAIL.n189 11.249
R378 VTAIL.n173 VTAIL.n114 11.249
R379 VTAIL.n144 VTAIL.n131 11.249
R380 VTAIL.n336 VTAIL.n320 10.4732
R381 VTAIL.n363 VTAIL.n308 10.4732
R382 VTAIL.n385 VTAIL.n298 10.4732
R383 VTAIL.n42 VTAIL.n26 10.4732
R384 VTAIL.n69 VTAIL.n14 10.4732
R385 VTAIL.n91 VTAIL.n4 10.4732
R386 VTAIL.n291 VTAIL.n204 10.4732
R387 VTAIL.n270 VTAIL.n215 10.4732
R388 VTAIL.n243 VTAIL.n227 10.4732
R389 VTAIL.n193 VTAIL.n106 10.4732
R390 VTAIL.n172 VTAIL.n117 10.4732
R391 VTAIL.n145 VTAIL.n129 10.4732
R392 VTAIL.n340 VTAIL.n339 9.69747
R393 VTAIL.n360 VTAIL.n359 9.69747
R394 VTAIL.n386 VTAIL.n296 9.69747
R395 VTAIL.n46 VTAIL.n45 9.69747
R396 VTAIL.n66 VTAIL.n65 9.69747
R397 VTAIL.n92 VTAIL.n2 9.69747
R398 VTAIL.n292 VTAIL.n202 9.69747
R399 VTAIL.n267 VTAIL.n266 9.69747
R400 VTAIL.n247 VTAIL.n246 9.69747
R401 VTAIL.n194 VTAIL.n104 9.69747
R402 VTAIL.n169 VTAIL.n168 9.69747
R403 VTAIL.n149 VTAIL.n148 9.69747
R404 VTAIL.n388 VTAIL.n387 9.45567
R405 VTAIL.n94 VTAIL.n93 9.45567
R406 VTAIL.n294 VTAIL.n293 9.45567
R407 VTAIL.n196 VTAIL.n195 9.45567
R408 VTAIL.n387 VTAIL.n386 9.3005
R409 VTAIL.n298 VTAIL.n297 9.3005
R410 VTAIL.n381 VTAIL.n380 9.3005
R411 VTAIL.n379 VTAIL.n378 9.3005
R412 VTAIL.n302 VTAIL.n301 9.3005
R413 VTAIL.n347 VTAIL.n346 9.3005
R414 VTAIL.n345 VTAIL.n344 9.3005
R415 VTAIL.n318 VTAIL.n317 9.3005
R416 VTAIL.n339 VTAIL.n338 9.3005
R417 VTAIL.n337 VTAIL.n336 9.3005
R418 VTAIL.n322 VTAIL.n321 9.3005
R419 VTAIL.n331 VTAIL.n330 9.3005
R420 VTAIL.n329 VTAIL.n328 9.3005
R421 VTAIL.n314 VTAIL.n313 9.3005
R422 VTAIL.n353 VTAIL.n352 9.3005
R423 VTAIL.n355 VTAIL.n354 9.3005
R424 VTAIL.n310 VTAIL.n309 9.3005
R425 VTAIL.n361 VTAIL.n360 9.3005
R426 VTAIL.n363 VTAIL.n362 9.3005
R427 VTAIL.n306 VTAIL.n305 9.3005
R428 VTAIL.n370 VTAIL.n369 9.3005
R429 VTAIL.n372 VTAIL.n371 9.3005
R430 VTAIL.n93 VTAIL.n92 9.3005
R431 VTAIL.n4 VTAIL.n3 9.3005
R432 VTAIL.n87 VTAIL.n86 9.3005
R433 VTAIL.n85 VTAIL.n84 9.3005
R434 VTAIL.n8 VTAIL.n7 9.3005
R435 VTAIL.n53 VTAIL.n52 9.3005
R436 VTAIL.n51 VTAIL.n50 9.3005
R437 VTAIL.n24 VTAIL.n23 9.3005
R438 VTAIL.n45 VTAIL.n44 9.3005
R439 VTAIL.n43 VTAIL.n42 9.3005
R440 VTAIL.n28 VTAIL.n27 9.3005
R441 VTAIL.n37 VTAIL.n36 9.3005
R442 VTAIL.n35 VTAIL.n34 9.3005
R443 VTAIL.n20 VTAIL.n19 9.3005
R444 VTAIL.n59 VTAIL.n58 9.3005
R445 VTAIL.n61 VTAIL.n60 9.3005
R446 VTAIL.n16 VTAIL.n15 9.3005
R447 VTAIL.n67 VTAIL.n66 9.3005
R448 VTAIL.n69 VTAIL.n68 9.3005
R449 VTAIL.n12 VTAIL.n11 9.3005
R450 VTAIL.n76 VTAIL.n75 9.3005
R451 VTAIL.n78 VTAIL.n77 9.3005
R452 VTAIL.n260 VTAIL.n259 9.3005
R453 VTAIL.n262 VTAIL.n261 9.3005
R454 VTAIL.n217 VTAIL.n216 9.3005
R455 VTAIL.n268 VTAIL.n267 9.3005
R456 VTAIL.n270 VTAIL.n269 9.3005
R457 VTAIL.n212 VTAIL.n211 9.3005
R458 VTAIL.n276 VTAIL.n275 9.3005
R459 VTAIL.n278 VTAIL.n277 9.3005
R460 VTAIL.n293 VTAIL.n292 9.3005
R461 VTAIL.n204 VTAIL.n203 9.3005
R462 VTAIL.n287 VTAIL.n286 9.3005
R463 VTAIL.n285 VTAIL.n284 9.3005
R464 VTAIL.n208 VTAIL.n207 9.3005
R465 VTAIL.n221 VTAIL.n220 9.3005
R466 VTAIL.n254 VTAIL.n253 9.3005
R467 VTAIL.n252 VTAIL.n251 9.3005
R468 VTAIL.n225 VTAIL.n224 9.3005
R469 VTAIL.n246 VTAIL.n245 9.3005
R470 VTAIL.n244 VTAIL.n243 9.3005
R471 VTAIL.n229 VTAIL.n228 9.3005
R472 VTAIL.n238 VTAIL.n237 9.3005
R473 VTAIL.n236 VTAIL.n235 9.3005
R474 VTAIL.n162 VTAIL.n161 9.3005
R475 VTAIL.n164 VTAIL.n163 9.3005
R476 VTAIL.n119 VTAIL.n118 9.3005
R477 VTAIL.n170 VTAIL.n169 9.3005
R478 VTAIL.n172 VTAIL.n171 9.3005
R479 VTAIL.n114 VTAIL.n113 9.3005
R480 VTAIL.n178 VTAIL.n177 9.3005
R481 VTAIL.n180 VTAIL.n179 9.3005
R482 VTAIL.n195 VTAIL.n194 9.3005
R483 VTAIL.n106 VTAIL.n105 9.3005
R484 VTAIL.n189 VTAIL.n188 9.3005
R485 VTAIL.n187 VTAIL.n186 9.3005
R486 VTAIL.n110 VTAIL.n109 9.3005
R487 VTAIL.n123 VTAIL.n122 9.3005
R488 VTAIL.n156 VTAIL.n155 9.3005
R489 VTAIL.n154 VTAIL.n153 9.3005
R490 VTAIL.n127 VTAIL.n126 9.3005
R491 VTAIL.n148 VTAIL.n147 9.3005
R492 VTAIL.n146 VTAIL.n145 9.3005
R493 VTAIL.n131 VTAIL.n130 9.3005
R494 VTAIL.n140 VTAIL.n139 9.3005
R495 VTAIL.n138 VTAIL.n137 9.3005
R496 VTAIL.n343 VTAIL.n318 8.92171
R497 VTAIL.n356 VTAIL.n310 8.92171
R498 VTAIL.n49 VTAIL.n24 8.92171
R499 VTAIL.n62 VTAIL.n16 8.92171
R500 VTAIL.n263 VTAIL.n217 8.92171
R501 VTAIL.n250 VTAIL.n225 8.92171
R502 VTAIL.n165 VTAIL.n119 8.92171
R503 VTAIL.n152 VTAIL.n127 8.92171
R504 VTAIL.n344 VTAIL.n316 8.14595
R505 VTAIL.n355 VTAIL.n312 8.14595
R506 VTAIL.n50 VTAIL.n22 8.14595
R507 VTAIL.n61 VTAIL.n18 8.14595
R508 VTAIL.n262 VTAIL.n219 8.14595
R509 VTAIL.n251 VTAIL.n223 8.14595
R510 VTAIL.n164 VTAIL.n121 8.14595
R511 VTAIL.n153 VTAIL.n125 8.14595
R512 VTAIL.n348 VTAIL.n347 7.3702
R513 VTAIL.n352 VTAIL.n351 7.3702
R514 VTAIL.n54 VTAIL.n53 7.3702
R515 VTAIL.n58 VTAIL.n57 7.3702
R516 VTAIL.n259 VTAIL.n258 7.3702
R517 VTAIL.n255 VTAIL.n254 7.3702
R518 VTAIL.n161 VTAIL.n160 7.3702
R519 VTAIL.n157 VTAIL.n156 7.3702
R520 VTAIL.n348 VTAIL.n314 6.59444
R521 VTAIL.n351 VTAIL.n314 6.59444
R522 VTAIL.n54 VTAIL.n20 6.59444
R523 VTAIL.n57 VTAIL.n20 6.59444
R524 VTAIL.n258 VTAIL.n221 6.59444
R525 VTAIL.n255 VTAIL.n221 6.59444
R526 VTAIL.n160 VTAIL.n123 6.59444
R527 VTAIL.n157 VTAIL.n123 6.59444
R528 VTAIL.n347 VTAIL.n316 5.81868
R529 VTAIL.n352 VTAIL.n312 5.81868
R530 VTAIL.n53 VTAIL.n22 5.81868
R531 VTAIL.n58 VTAIL.n18 5.81868
R532 VTAIL.n259 VTAIL.n219 5.81868
R533 VTAIL.n254 VTAIL.n223 5.81868
R534 VTAIL.n161 VTAIL.n121 5.81868
R535 VTAIL.n156 VTAIL.n125 5.81868
R536 VTAIL.n344 VTAIL.n343 5.04292
R537 VTAIL.n356 VTAIL.n355 5.04292
R538 VTAIL.n50 VTAIL.n49 5.04292
R539 VTAIL.n62 VTAIL.n61 5.04292
R540 VTAIL.n263 VTAIL.n262 5.04292
R541 VTAIL.n251 VTAIL.n250 5.04292
R542 VTAIL.n165 VTAIL.n164 5.04292
R543 VTAIL.n153 VTAIL.n152 5.04292
R544 VTAIL.n236 VTAIL.n232 4.38563
R545 VTAIL.n138 VTAIL.n134 4.38563
R546 VTAIL.n329 VTAIL.n325 4.38563
R547 VTAIL.n35 VTAIL.n31 4.38563
R548 VTAIL.n340 VTAIL.n318 4.26717
R549 VTAIL.n359 VTAIL.n310 4.26717
R550 VTAIL.n388 VTAIL.n296 4.26717
R551 VTAIL.n46 VTAIL.n24 4.26717
R552 VTAIL.n65 VTAIL.n16 4.26717
R553 VTAIL.n94 VTAIL.n2 4.26717
R554 VTAIL.n294 VTAIL.n202 4.26717
R555 VTAIL.n266 VTAIL.n217 4.26717
R556 VTAIL.n247 VTAIL.n225 4.26717
R557 VTAIL.n196 VTAIL.n104 4.26717
R558 VTAIL.n168 VTAIL.n119 4.26717
R559 VTAIL.n149 VTAIL.n127 4.26717
R560 VTAIL.n339 VTAIL.n320 3.49141
R561 VTAIL.n360 VTAIL.n308 3.49141
R562 VTAIL.n386 VTAIL.n385 3.49141
R563 VTAIL.n45 VTAIL.n26 3.49141
R564 VTAIL.n66 VTAIL.n14 3.49141
R565 VTAIL.n92 VTAIL.n91 3.49141
R566 VTAIL.n292 VTAIL.n291 3.49141
R567 VTAIL.n267 VTAIL.n215 3.49141
R568 VTAIL.n246 VTAIL.n227 3.49141
R569 VTAIL.n194 VTAIL.n193 3.49141
R570 VTAIL.n169 VTAIL.n117 3.49141
R571 VTAIL.n148 VTAIL.n129 3.49141
R572 VTAIL.n336 VTAIL.n335 2.71565
R573 VTAIL.n364 VTAIL.n363 2.71565
R574 VTAIL.n382 VTAIL.n298 2.71565
R575 VTAIL.n42 VTAIL.n41 2.71565
R576 VTAIL.n70 VTAIL.n69 2.71565
R577 VTAIL.n88 VTAIL.n4 2.71565
R578 VTAIL.n288 VTAIL.n204 2.71565
R579 VTAIL.n271 VTAIL.n270 2.71565
R580 VTAIL.n243 VTAIL.n242 2.71565
R581 VTAIL.n190 VTAIL.n106 2.71565
R582 VTAIL.n173 VTAIL.n172 2.71565
R583 VTAIL.n145 VTAIL.n144 2.71565
R584 VTAIL.n103 VTAIL.n101 2.19878
R585 VTAIL.n197 VTAIL.n103 2.19878
R586 VTAIL.n201 VTAIL.n199 2.19878
R587 VTAIL.n295 VTAIL.n201 2.19878
R588 VTAIL.n99 VTAIL.n97 2.19878
R589 VTAIL.n97 VTAIL.n95 2.19878
R590 VTAIL.n391 VTAIL.n389 2.19878
R591 VTAIL.n332 VTAIL.n322 1.93989
R592 VTAIL.n368 VTAIL.n306 1.93989
R593 VTAIL.n381 VTAIL.n300 1.93989
R594 VTAIL.n38 VTAIL.n28 1.93989
R595 VTAIL.n74 VTAIL.n12 1.93989
R596 VTAIL.n87 VTAIL.n6 1.93989
R597 VTAIL.n287 VTAIL.n206 1.93989
R598 VTAIL.n274 VTAIL.n212 1.93989
R599 VTAIL.n239 VTAIL.n229 1.93989
R600 VTAIL.n189 VTAIL.n108 1.93989
R601 VTAIL.n176 VTAIL.n114 1.93989
R602 VTAIL.n141 VTAIL.n131 1.93989
R603 VTAIL VTAIL.n1 1.7074
R604 VTAIL.n199 VTAIL.n197 1.56947
R605 VTAIL.n95 VTAIL.n1 1.56947
R606 VTAIL.n390 VTAIL.t0 1.17418
R607 VTAIL.n390 VTAIL.t2 1.17418
R608 VTAIL.n0 VTAIL.t8 1.17418
R609 VTAIL.n0 VTAIL.t3 1.17418
R610 VTAIL.n96 VTAIL.t9 1.17418
R611 VTAIL.n96 VTAIL.t12 1.17418
R612 VTAIL.n98 VTAIL.t16 1.17418
R613 VTAIL.n98 VTAIL.t17 1.17418
R614 VTAIL.n200 VTAIL.t11 1.17418
R615 VTAIL.n200 VTAIL.t14 1.17418
R616 VTAIL.n198 VTAIL.t10 1.17418
R617 VTAIL.n198 VTAIL.t18 1.17418
R618 VTAIL.n102 VTAIL.t6 1.17418
R619 VTAIL.n102 VTAIL.t7 1.17418
R620 VTAIL.n100 VTAIL.t4 1.17418
R621 VTAIL.n100 VTAIL.t1 1.17418
R622 VTAIL.n331 VTAIL.n324 1.16414
R623 VTAIL.n369 VTAIL.n304 1.16414
R624 VTAIL.n378 VTAIL.n377 1.16414
R625 VTAIL.n37 VTAIL.n30 1.16414
R626 VTAIL.n75 VTAIL.n10 1.16414
R627 VTAIL.n84 VTAIL.n83 1.16414
R628 VTAIL.n284 VTAIL.n283 1.16414
R629 VTAIL.n275 VTAIL.n210 1.16414
R630 VTAIL.n238 VTAIL.n231 1.16414
R631 VTAIL.n186 VTAIL.n185 1.16414
R632 VTAIL.n177 VTAIL.n112 1.16414
R633 VTAIL.n140 VTAIL.n133 1.16414
R634 VTAIL VTAIL.n391 0.491879
R635 VTAIL.n328 VTAIL.n327 0.388379
R636 VTAIL.n373 VTAIL.n372 0.388379
R637 VTAIL.n374 VTAIL.n302 0.388379
R638 VTAIL.n34 VTAIL.n33 0.388379
R639 VTAIL.n79 VTAIL.n78 0.388379
R640 VTAIL.n80 VTAIL.n8 0.388379
R641 VTAIL.n280 VTAIL.n208 0.388379
R642 VTAIL.n279 VTAIL.n278 0.388379
R643 VTAIL.n235 VTAIL.n234 0.388379
R644 VTAIL.n182 VTAIL.n110 0.388379
R645 VTAIL.n181 VTAIL.n180 0.388379
R646 VTAIL.n137 VTAIL.n136 0.388379
R647 VTAIL.n330 VTAIL.n329 0.155672
R648 VTAIL.n330 VTAIL.n321 0.155672
R649 VTAIL.n337 VTAIL.n321 0.155672
R650 VTAIL.n338 VTAIL.n337 0.155672
R651 VTAIL.n338 VTAIL.n317 0.155672
R652 VTAIL.n345 VTAIL.n317 0.155672
R653 VTAIL.n346 VTAIL.n345 0.155672
R654 VTAIL.n346 VTAIL.n313 0.155672
R655 VTAIL.n353 VTAIL.n313 0.155672
R656 VTAIL.n354 VTAIL.n353 0.155672
R657 VTAIL.n354 VTAIL.n309 0.155672
R658 VTAIL.n361 VTAIL.n309 0.155672
R659 VTAIL.n362 VTAIL.n361 0.155672
R660 VTAIL.n362 VTAIL.n305 0.155672
R661 VTAIL.n370 VTAIL.n305 0.155672
R662 VTAIL.n371 VTAIL.n370 0.155672
R663 VTAIL.n371 VTAIL.n301 0.155672
R664 VTAIL.n379 VTAIL.n301 0.155672
R665 VTAIL.n380 VTAIL.n379 0.155672
R666 VTAIL.n380 VTAIL.n297 0.155672
R667 VTAIL.n387 VTAIL.n297 0.155672
R668 VTAIL.n36 VTAIL.n35 0.155672
R669 VTAIL.n36 VTAIL.n27 0.155672
R670 VTAIL.n43 VTAIL.n27 0.155672
R671 VTAIL.n44 VTAIL.n43 0.155672
R672 VTAIL.n44 VTAIL.n23 0.155672
R673 VTAIL.n51 VTAIL.n23 0.155672
R674 VTAIL.n52 VTAIL.n51 0.155672
R675 VTAIL.n52 VTAIL.n19 0.155672
R676 VTAIL.n59 VTAIL.n19 0.155672
R677 VTAIL.n60 VTAIL.n59 0.155672
R678 VTAIL.n60 VTAIL.n15 0.155672
R679 VTAIL.n67 VTAIL.n15 0.155672
R680 VTAIL.n68 VTAIL.n67 0.155672
R681 VTAIL.n68 VTAIL.n11 0.155672
R682 VTAIL.n76 VTAIL.n11 0.155672
R683 VTAIL.n77 VTAIL.n76 0.155672
R684 VTAIL.n77 VTAIL.n7 0.155672
R685 VTAIL.n85 VTAIL.n7 0.155672
R686 VTAIL.n86 VTAIL.n85 0.155672
R687 VTAIL.n86 VTAIL.n3 0.155672
R688 VTAIL.n93 VTAIL.n3 0.155672
R689 VTAIL.n293 VTAIL.n203 0.155672
R690 VTAIL.n286 VTAIL.n203 0.155672
R691 VTAIL.n286 VTAIL.n285 0.155672
R692 VTAIL.n285 VTAIL.n207 0.155672
R693 VTAIL.n277 VTAIL.n207 0.155672
R694 VTAIL.n277 VTAIL.n276 0.155672
R695 VTAIL.n276 VTAIL.n211 0.155672
R696 VTAIL.n269 VTAIL.n211 0.155672
R697 VTAIL.n269 VTAIL.n268 0.155672
R698 VTAIL.n268 VTAIL.n216 0.155672
R699 VTAIL.n261 VTAIL.n216 0.155672
R700 VTAIL.n261 VTAIL.n260 0.155672
R701 VTAIL.n260 VTAIL.n220 0.155672
R702 VTAIL.n253 VTAIL.n220 0.155672
R703 VTAIL.n253 VTAIL.n252 0.155672
R704 VTAIL.n252 VTAIL.n224 0.155672
R705 VTAIL.n245 VTAIL.n224 0.155672
R706 VTAIL.n245 VTAIL.n244 0.155672
R707 VTAIL.n244 VTAIL.n228 0.155672
R708 VTAIL.n237 VTAIL.n228 0.155672
R709 VTAIL.n237 VTAIL.n236 0.155672
R710 VTAIL.n195 VTAIL.n105 0.155672
R711 VTAIL.n188 VTAIL.n105 0.155672
R712 VTAIL.n188 VTAIL.n187 0.155672
R713 VTAIL.n187 VTAIL.n109 0.155672
R714 VTAIL.n179 VTAIL.n109 0.155672
R715 VTAIL.n179 VTAIL.n178 0.155672
R716 VTAIL.n178 VTAIL.n113 0.155672
R717 VTAIL.n171 VTAIL.n113 0.155672
R718 VTAIL.n171 VTAIL.n170 0.155672
R719 VTAIL.n170 VTAIL.n118 0.155672
R720 VTAIL.n163 VTAIL.n118 0.155672
R721 VTAIL.n163 VTAIL.n162 0.155672
R722 VTAIL.n162 VTAIL.n122 0.155672
R723 VTAIL.n155 VTAIL.n122 0.155672
R724 VTAIL.n155 VTAIL.n154 0.155672
R725 VTAIL.n154 VTAIL.n126 0.155672
R726 VTAIL.n147 VTAIL.n126 0.155672
R727 VTAIL.n147 VTAIL.n146 0.155672
R728 VTAIL.n146 VTAIL.n130 0.155672
R729 VTAIL.n139 VTAIL.n130 0.155672
R730 VTAIL.n139 VTAIL.n138 0.155672
R731 VDD1.n88 VDD1.n0 289.615
R732 VDD1.n183 VDD1.n95 289.615
R733 VDD1.n89 VDD1.n88 185
R734 VDD1.n87 VDD1.n86 185
R735 VDD1.n4 VDD1.n3 185
R736 VDD1.n81 VDD1.n80 185
R737 VDD1.n79 VDD1.n78 185
R738 VDD1.n77 VDD1.n7 185
R739 VDD1.n11 VDD1.n8 185
R740 VDD1.n72 VDD1.n71 185
R741 VDD1.n70 VDD1.n69 185
R742 VDD1.n13 VDD1.n12 185
R743 VDD1.n64 VDD1.n63 185
R744 VDD1.n62 VDD1.n61 185
R745 VDD1.n17 VDD1.n16 185
R746 VDD1.n56 VDD1.n55 185
R747 VDD1.n54 VDD1.n53 185
R748 VDD1.n21 VDD1.n20 185
R749 VDD1.n48 VDD1.n47 185
R750 VDD1.n46 VDD1.n45 185
R751 VDD1.n25 VDD1.n24 185
R752 VDD1.n40 VDD1.n39 185
R753 VDD1.n38 VDD1.n37 185
R754 VDD1.n29 VDD1.n28 185
R755 VDD1.n32 VDD1.n31 185
R756 VDD1.n126 VDD1.n125 185
R757 VDD1.n123 VDD1.n122 185
R758 VDD1.n132 VDD1.n131 185
R759 VDD1.n134 VDD1.n133 185
R760 VDD1.n119 VDD1.n118 185
R761 VDD1.n140 VDD1.n139 185
R762 VDD1.n142 VDD1.n141 185
R763 VDD1.n115 VDD1.n114 185
R764 VDD1.n148 VDD1.n147 185
R765 VDD1.n150 VDD1.n149 185
R766 VDD1.n111 VDD1.n110 185
R767 VDD1.n156 VDD1.n155 185
R768 VDD1.n158 VDD1.n157 185
R769 VDD1.n107 VDD1.n106 185
R770 VDD1.n164 VDD1.n163 185
R771 VDD1.n167 VDD1.n166 185
R772 VDD1.n165 VDD1.n103 185
R773 VDD1.n172 VDD1.n102 185
R774 VDD1.n174 VDD1.n173 185
R775 VDD1.n176 VDD1.n175 185
R776 VDD1.n99 VDD1.n98 185
R777 VDD1.n182 VDD1.n181 185
R778 VDD1.n184 VDD1.n183 185
R779 VDD1.t9 VDD1.n30 147.659
R780 VDD1.t6 VDD1.n124 147.659
R781 VDD1.n88 VDD1.n87 104.615
R782 VDD1.n87 VDD1.n3 104.615
R783 VDD1.n80 VDD1.n3 104.615
R784 VDD1.n80 VDD1.n79 104.615
R785 VDD1.n79 VDD1.n7 104.615
R786 VDD1.n11 VDD1.n7 104.615
R787 VDD1.n71 VDD1.n11 104.615
R788 VDD1.n71 VDD1.n70 104.615
R789 VDD1.n70 VDD1.n12 104.615
R790 VDD1.n63 VDD1.n12 104.615
R791 VDD1.n63 VDD1.n62 104.615
R792 VDD1.n62 VDD1.n16 104.615
R793 VDD1.n55 VDD1.n16 104.615
R794 VDD1.n55 VDD1.n54 104.615
R795 VDD1.n54 VDD1.n20 104.615
R796 VDD1.n47 VDD1.n20 104.615
R797 VDD1.n47 VDD1.n46 104.615
R798 VDD1.n46 VDD1.n24 104.615
R799 VDD1.n39 VDD1.n24 104.615
R800 VDD1.n39 VDD1.n38 104.615
R801 VDD1.n38 VDD1.n28 104.615
R802 VDD1.n31 VDD1.n28 104.615
R803 VDD1.n125 VDD1.n122 104.615
R804 VDD1.n132 VDD1.n122 104.615
R805 VDD1.n133 VDD1.n132 104.615
R806 VDD1.n133 VDD1.n118 104.615
R807 VDD1.n140 VDD1.n118 104.615
R808 VDD1.n141 VDD1.n140 104.615
R809 VDD1.n141 VDD1.n114 104.615
R810 VDD1.n148 VDD1.n114 104.615
R811 VDD1.n149 VDD1.n148 104.615
R812 VDD1.n149 VDD1.n110 104.615
R813 VDD1.n156 VDD1.n110 104.615
R814 VDD1.n157 VDD1.n156 104.615
R815 VDD1.n157 VDD1.n106 104.615
R816 VDD1.n164 VDD1.n106 104.615
R817 VDD1.n166 VDD1.n164 104.615
R818 VDD1.n166 VDD1.n165 104.615
R819 VDD1.n165 VDD1.n102 104.615
R820 VDD1.n174 VDD1.n102 104.615
R821 VDD1.n175 VDD1.n174 104.615
R822 VDD1.n175 VDD1.n98 104.615
R823 VDD1.n182 VDD1.n98 104.615
R824 VDD1.n183 VDD1.n182 104.615
R825 VDD1.n191 VDD1.n190 63.6756
R826 VDD1.n94 VDD1.n93 62.0824
R827 VDD1.n193 VDD1.n192 62.0822
R828 VDD1.n189 VDD1.n188 62.0822
R829 VDD1.n94 VDD1.n92 52.42
R830 VDD1.n189 VDD1.n187 52.42
R831 VDD1.n31 VDD1.t9 52.3082
R832 VDD1.n125 VDD1.t6 52.3082
R833 VDD1.n193 VDD1.n191 50.3824
R834 VDD1.n32 VDD1.n30 15.6677
R835 VDD1.n126 VDD1.n124 15.6677
R836 VDD1.n78 VDD1.n77 13.1884
R837 VDD1.n173 VDD1.n172 13.1884
R838 VDD1.n81 VDD1.n6 12.8005
R839 VDD1.n76 VDD1.n8 12.8005
R840 VDD1.n33 VDD1.n29 12.8005
R841 VDD1.n127 VDD1.n123 12.8005
R842 VDD1.n171 VDD1.n103 12.8005
R843 VDD1.n176 VDD1.n101 12.8005
R844 VDD1.n82 VDD1.n4 12.0247
R845 VDD1.n73 VDD1.n72 12.0247
R846 VDD1.n37 VDD1.n36 12.0247
R847 VDD1.n131 VDD1.n130 12.0247
R848 VDD1.n168 VDD1.n167 12.0247
R849 VDD1.n177 VDD1.n99 12.0247
R850 VDD1.n86 VDD1.n85 11.249
R851 VDD1.n69 VDD1.n10 11.249
R852 VDD1.n40 VDD1.n27 11.249
R853 VDD1.n134 VDD1.n121 11.249
R854 VDD1.n163 VDD1.n105 11.249
R855 VDD1.n181 VDD1.n180 11.249
R856 VDD1.n89 VDD1.n2 10.4732
R857 VDD1.n68 VDD1.n13 10.4732
R858 VDD1.n41 VDD1.n25 10.4732
R859 VDD1.n135 VDD1.n119 10.4732
R860 VDD1.n162 VDD1.n107 10.4732
R861 VDD1.n184 VDD1.n97 10.4732
R862 VDD1.n90 VDD1.n0 9.69747
R863 VDD1.n65 VDD1.n64 9.69747
R864 VDD1.n45 VDD1.n44 9.69747
R865 VDD1.n139 VDD1.n138 9.69747
R866 VDD1.n159 VDD1.n158 9.69747
R867 VDD1.n185 VDD1.n95 9.69747
R868 VDD1.n92 VDD1.n91 9.45567
R869 VDD1.n187 VDD1.n186 9.45567
R870 VDD1.n58 VDD1.n57 9.3005
R871 VDD1.n60 VDD1.n59 9.3005
R872 VDD1.n15 VDD1.n14 9.3005
R873 VDD1.n66 VDD1.n65 9.3005
R874 VDD1.n68 VDD1.n67 9.3005
R875 VDD1.n10 VDD1.n9 9.3005
R876 VDD1.n74 VDD1.n73 9.3005
R877 VDD1.n76 VDD1.n75 9.3005
R878 VDD1.n91 VDD1.n90 9.3005
R879 VDD1.n2 VDD1.n1 9.3005
R880 VDD1.n85 VDD1.n84 9.3005
R881 VDD1.n83 VDD1.n82 9.3005
R882 VDD1.n6 VDD1.n5 9.3005
R883 VDD1.n19 VDD1.n18 9.3005
R884 VDD1.n52 VDD1.n51 9.3005
R885 VDD1.n50 VDD1.n49 9.3005
R886 VDD1.n23 VDD1.n22 9.3005
R887 VDD1.n44 VDD1.n43 9.3005
R888 VDD1.n42 VDD1.n41 9.3005
R889 VDD1.n27 VDD1.n26 9.3005
R890 VDD1.n36 VDD1.n35 9.3005
R891 VDD1.n34 VDD1.n33 9.3005
R892 VDD1.n186 VDD1.n185 9.3005
R893 VDD1.n97 VDD1.n96 9.3005
R894 VDD1.n180 VDD1.n179 9.3005
R895 VDD1.n178 VDD1.n177 9.3005
R896 VDD1.n101 VDD1.n100 9.3005
R897 VDD1.n146 VDD1.n145 9.3005
R898 VDD1.n144 VDD1.n143 9.3005
R899 VDD1.n117 VDD1.n116 9.3005
R900 VDD1.n138 VDD1.n137 9.3005
R901 VDD1.n136 VDD1.n135 9.3005
R902 VDD1.n121 VDD1.n120 9.3005
R903 VDD1.n130 VDD1.n129 9.3005
R904 VDD1.n128 VDD1.n127 9.3005
R905 VDD1.n113 VDD1.n112 9.3005
R906 VDD1.n152 VDD1.n151 9.3005
R907 VDD1.n154 VDD1.n153 9.3005
R908 VDD1.n109 VDD1.n108 9.3005
R909 VDD1.n160 VDD1.n159 9.3005
R910 VDD1.n162 VDD1.n161 9.3005
R911 VDD1.n105 VDD1.n104 9.3005
R912 VDD1.n169 VDD1.n168 9.3005
R913 VDD1.n171 VDD1.n170 9.3005
R914 VDD1.n61 VDD1.n15 8.92171
R915 VDD1.n48 VDD1.n23 8.92171
R916 VDD1.n142 VDD1.n117 8.92171
R917 VDD1.n155 VDD1.n109 8.92171
R918 VDD1.n60 VDD1.n17 8.14595
R919 VDD1.n49 VDD1.n21 8.14595
R920 VDD1.n143 VDD1.n115 8.14595
R921 VDD1.n154 VDD1.n111 8.14595
R922 VDD1.n57 VDD1.n56 7.3702
R923 VDD1.n53 VDD1.n52 7.3702
R924 VDD1.n147 VDD1.n146 7.3702
R925 VDD1.n151 VDD1.n150 7.3702
R926 VDD1.n56 VDD1.n19 6.59444
R927 VDD1.n53 VDD1.n19 6.59444
R928 VDD1.n147 VDD1.n113 6.59444
R929 VDD1.n150 VDD1.n113 6.59444
R930 VDD1.n57 VDD1.n17 5.81868
R931 VDD1.n52 VDD1.n21 5.81868
R932 VDD1.n146 VDD1.n115 5.81868
R933 VDD1.n151 VDD1.n111 5.81868
R934 VDD1.n61 VDD1.n60 5.04292
R935 VDD1.n49 VDD1.n48 5.04292
R936 VDD1.n143 VDD1.n142 5.04292
R937 VDD1.n155 VDD1.n154 5.04292
R938 VDD1.n34 VDD1.n30 4.38563
R939 VDD1.n128 VDD1.n124 4.38563
R940 VDD1.n92 VDD1.n0 4.26717
R941 VDD1.n64 VDD1.n15 4.26717
R942 VDD1.n45 VDD1.n23 4.26717
R943 VDD1.n139 VDD1.n117 4.26717
R944 VDD1.n158 VDD1.n109 4.26717
R945 VDD1.n187 VDD1.n95 4.26717
R946 VDD1.n90 VDD1.n89 3.49141
R947 VDD1.n65 VDD1.n13 3.49141
R948 VDD1.n44 VDD1.n25 3.49141
R949 VDD1.n138 VDD1.n119 3.49141
R950 VDD1.n159 VDD1.n107 3.49141
R951 VDD1.n185 VDD1.n184 3.49141
R952 VDD1.n86 VDD1.n2 2.71565
R953 VDD1.n69 VDD1.n68 2.71565
R954 VDD1.n41 VDD1.n40 2.71565
R955 VDD1.n135 VDD1.n134 2.71565
R956 VDD1.n163 VDD1.n162 2.71565
R957 VDD1.n181 VDD1.n97 2.71565
R958 VDD1.n85 VDD1.n4 1.93989
R959 VDD1.n72 VDD1.n10 1.93989
R960 VDD1.n37 VDD1.n27 1.93989
R961 VDD1.n131 VDD1.n121 1.93989
R962 VDD1.n167 VDD1.n105 1.93989
R963 VDD1.n180 VDD1.n99 1.93989
R964 VDD1 VDD1.n193 1.59102
R965 VDD1.n192 VDD1.t4 1.17418
R966 VDD1.n192 VDD1.t0 1.17418
R967 VDD1.n93 VDD1.t7 1.17418
R968 VDD1.n93 VDD1.t3 1.17418
R969 VDD1.n190 VDD1.t2 1.17418
R970 VDD1.n190 VDD1.t5 1.17418
R971 VDD1.n188 VDD1.t8 1.17418
R972 VDD1.n188 VDD1.t1 1.17418
R973 VDD1.n82 VDD1.n81 1.16414
R974 VDD1.n73 VDD1.n8 1.16414
R975 VDD1.n36 VDD1.n29 1.16414
R976 VDD1.n130 VDD1.n123 1.16414
R977 VDD1.n168 VDD1.n103 1.16414
R978 VDD1.n177 VDD1.n176 1.16414
R979 VDD1 VDD1.n94 0.608259
R980 VDD1.n191 VDD1.n189 0.494723
R981 VDD1.n78 VDD1.n6 0.388379
R982 VDD1.n77 VDD1.n76 0.388379
R983 VDD1.n33 VDD1.n32 0.388379
R984 VDD1.n127 VDD1.n126 0.388379
R985 VDD1.n172 VDD1.n171 0.388379
R986 VDD1.n173 VDD1.n101 0.388379
R987 VDD1.n91 VDD1.n1 0.155672
R988 VDD1.n84 VDD1.n1 0.155672
R989 VDD1.n84 VDD1.n83 0.155672
R990 VDD1.n83 VDD1.n5 0.155672
R991 VDD1.n75 VDD1.n5 0.155672
R992 VDD1.n75 VDD1.n74 0.155672
R993 VDD1.n74 VDD1.n9 0.155672
R994 VDD1.n67 VDD1.n9 0.155672
R995 VDD1.n67 VDD1.n66 0.155672
R996 VDD1.n66 VDD1.n14 0.155672
R997 VDD1.n59 VDD1.n14 0.155672
R998 VDD1.n59 VDD1.n58 0.155672
R999 VDD1.n58 VDD1.n18 0.155672
R1000 VDD1.n51 VDD1.n18 0.155672
R1001 VDD1.n51 VDD1.n50 0.155672
R1002 VDD1.n50 VDD1.n22 0.155672
R1003 VDD1.n43 VDD1.n22 0.155672
R1004 VDD1.n43 VDD1.n42 0.155672
R1005 VDD1.n42 VDD1.n26 0.155672
R1006 VDD1.n35 VDD1.n26 0.155672
R1007 VDD1.n35 VDD1.n34 0.155672
R1008 VDD1.n129 VDD1.n128 0.155672
R1009 VDD1.n129 VDD1.n120 0.155672
R1010 VDD1.n136 VDD1.n120 0.155672
R1011 VDD1.n137 VDD1.n136 0.155672
R1012 VDD1.n137 VDD1.n116 0.155672
R1013 VDD1.n144 VDD1.n116 0.155672
R1014 VDD1.n145 VDD1.n144 0.155672
R1015 VDD1.n145 VDD1.n112 0.155672
R1016 VDD1.n152 VDD1.n112 0.155672
R1017 VDD1.n153 VDD1.n152 0.155672
R1018 VDD1.n153 VDD1.n108 0.155672
R1019 VDD1.n160 VDD1.n108 0.155672
R1020 VDD1.n161 VDD1.n160 0.155672
R1021 VDD1.n161 VDD1.n104 0.155672
R1022 VDD1.n169 VDD1.n104 0.155672
R1023 VDD1.n170 VDD1.n169 0.155672
R1024 VDD1.n170 VDD1.n100 0.155672
R1025 VDD1.n178 VDD1.n100 0.155672
R1026 VDD1.n179 VDD1.n178 0.155672
R1027 VDD1.n179 VDD1.n96 0.155672
R1028 VDD1.n186 VDD1.n96 0.155672
R1029 B.n1043 B.n1042 585
R1030 B.n1044 B.n1043 585
R1031 B.n403 B.n158 585
R1032 B.n402 B.n401 585
R1033 B.n400 B.n399 585
R1034 B.n398 B.n397 585
R1035 B.n396 B.n395 585
R1036 B.n394 B.n393 585
R1037 B.n392 B.n391 585
R1038 B.n390 B.n389 585
R1039 B.n388 B.n387 585
R1040 B.n386 B.n385 585
R1041 B.n384 B.n383 585
R1042 B.n382 B.n381 585
R1043 B.n380 B.n379 585
R1044 B.n378 B.n377 585
R1045 B.n376 B.n375 585
R1046 B.n374 B.n373 585
R1047 B.n372 B.n371 585
R1048 B.n370 B.n369 585
R1049 B.n368 B.n367 585
R1050 B.n366 B.n365 585
R1051 B.n364 B.n363 585
R1052 B.n362 B.n361 585
R1053 B.n360 B.n359 585
R1054 B.n358 B.n357 585
R1055 B.n356 B.n355 585
R1056 B.n354 B.n353 585
R1057 B.n352 B.n351 585
R1058 B.n350 B.n349 585
R1059 B.n348 B.n347 585
R1060 B.n346 B.n345 585
R1061 B.n344 B.n343 585
R1062 B.n342 B.n341 585
R1063 B.n340 B.n339 585
R1064 B.n338 B.n337 585
R1065 B.n336 B.n335 585
R1066 B.n334 B.n333 585
R1067 B.n332 B.n331 585
R1068 B.n330 B.n329 585
R1069 B.n328 B.n327 585
R1070 B.n326 B.n325 585
R1071 B.n324 B.n323 585
R1072 B.n322 B.n321 585
R1073 B.n320 B.n319 585
R1074 B.n318 B.n317 585
R1075 B.n316 B.n315 585
R1076 B.n314 B.n313 585
R1077 B.n312 B.n311 585
R1078 B.n310 B.n309 585
R1079 B.n308 B.n307 585
R1080 B.n306 B.n305 585
R1081 B.n304 B.n303 585
R1082 B.n302 B.n301 585
R1083 B.n300 B.n299 585
R1084 B.n298 B.n297 585
R1085 B.n296 B.n295 585
R1086 B.n293 B.n292 585
R1087 B.n291 B.n290 585
R1088 B.n289 B.n288 585
R1089 B.n287 B.n286 585
R1090 B.n285 B.n284 585
R1091 B.n283 B.n282 585
R1092 B.n281 B.n280 585
R1093 B.n279 B.n278 585
R1094 B.n277 B.n276 585
R1095 B.n275 B.n274 585
R1096 B.n273 B.n272 585
R1097 B.n271 B.n270 585
R1098 B.n269 B.n268 585
R1099 B.n267 B.n266 585
R1100 B.n265 B.n264 585
R1101 B.n263 B.n262 585
R1102 B.n261 B.n260 585
R1103 B.n259 B.n258 585
R1104 B.n257 B.n256 585
R1105 B.n255 B.n254 585
R1106 B.n253 B.n252 585
R1107 B.n251 B.n250 585
R1108 B.n249 B.n248 585
R1109 B.n247 B.n246 585
R1110 B.n245 B.n244 585
R1111 B.n243 B.n242 585
R1112 B.n241 B.n240 585
R1113 B.n239 B.n238 585
R1114 B.n237 B.n236 585
R1115 B.n235 B.n234 585
R1116 B.n233 B.n232 585
R1117 B.n231 B.n230 585
R1118 B.n229 B.n228 585
R1119 B.n227 B.n226 585
R1120 B.n225 B.n224 585
R1121 B.n223 B.n222 585
R1122 B.n221 B.n220 585
R1123 B.n219 B.n218 585
R1124 B.n217 B.n216 585
R1125 B.n215 B.n214 585
R1126 B.n213 B.n212 585
R1127 B.n211 B.n210 585
R1128 B.n209 B.n208 585
R1129 B.n207 B.n206 585
R1130 B.n205 B.n204 585
R1131 B.n203 B.n202 585
R1132 B.n201 B.n200 585
R1133 B.n199 B.n198 585
R1134 B.n197 B.n196 585
R1135 B.n195 B.n194 585
R1136 B.n193 B.n192 585
R1137 B.n191 B.n190 585
R1138 B.n189 B.n188 585
R1139 B.n187 B.n186 585
R1140 B.n185 B.n184 585
R1141 B.n183 B.n182 585
R1142 B.n181 B.n180 585
R1143 B.n179 B.n178 585
R1144 B.n177 B.n176 585
R1145 B.n175 B.n174 585
R1146 B.n173 B.n172 585
R1147 B.n171 B.n170 585
R1148 B.n169 B.n168 585
R1149 B.n167 B.n166 585
R1150 B.n165 B.n164 585
R1151 B.n1041 B.n97 585
R1152 B.n1045 B.n97 585
R1153 B.n1040 B.n96 585
R1154 B.n1046 B.n96 585
R1155 B.n1039 B.n1038 585
R1156 B.n1038 B.n92 585
R1157 B.n1037 B.n91 585
R1158 B.n1052 B.n91 585
R1159 B.n1036 B.n90 585
R1160 B.n1053 B.n90 585
R1161 B.n1035 B.n89 585
R1162 B.n1054 B.n89 585
R1163 B.n1034 B.n1033 585
R1164 B.n1033 B.n88 585
R1165 B.n1032 B.n84 585
R1166 B.n1060 B.n84 585
R1167 B.n1031 B.n83 585
R1168 B.n1061 B.n83 585
R1169 B.n1030 B.n82 585
R1170 B.n1062 B.n82 585
R1171 B.n1029 B.n1028 585
R1172 B.n1028 B.n78 585
R1173 B.n1027 B.n77 585
R1174 B.n1068 B.n77 585
R1175 B.n1026 B.n76 585
R1176 B.n1069 B.n76 585
R1177 B.n1025 B.n75 585
R1178 B.n1070 B.n75 585
R1179 B.n1024 B.n1023 585
R1180 B.n1023 B.n71 585
R1181 B.n1022 B.n70 585
R1182 B.n1076 B.n70 585
R1183 B.n1021 B.n69 585
R1184 B.n1077 B.n69 585
R1185 B.n1020 B.n68 585
R1186 B.n1078 B.n68 585
R1187 B.n1019 B.n1018 585
R1188 B.n1018 B.n64 585
R1189 B.n1017 B.n63 585
R1190 B.n1084 B.n63 585
R1191 B.n1016 B.n62 585
R1192 B.n1085 B.n62 585
R1193 B.n1015 B.n61 585
R1194 B.n1086 B.n61 585
R1195 B.n1014 B.n1013 585
R1196 B.n1013 B.n57 585
R1197 B.n1012 B.n56 585
R1198 B.n1092 B.n56 585
R1199 B.n1011 B.n55 585
R1200 B.n1093 B.n55 585
R1201 B.n1010 B.n54 585
R1202 B.n1094 B.n54 585
R1203 B.n1009 B.n1008 585
R1204 B.n1008 B.n50 585
R1205 B.n1007 B.n49 585
R1206 B.n1100 B.n49 585
R1207 B.n1006 B.n48 585
R1208 B.n1101 B.n48 585
R1209 B.n1005 B.n47 585
R1210 B.n1102 B.n47 585
R1211 B.n1004 B.n1003 585
R1212 B.n1003 B.n43 585
R1213 B.n1002 B.n42 585
R1214 B.n1108 B.n42 585
R1215 B.n1001 B.n41 585
R1216 B.n1109 B.n41 585
R1217 B.n1000 B.n40 585
R1218 B.n1110 B.n40 585
R1219 B.n999 B.n998 585
R1220 B.n998 B.n36 585
R1221 B.n997 B.n35 585
R1222 B.n1116 B.n35 585
R1223 B.n996 B.n34 585
R1224 B.n1117 B.n34 585
R1225 B.n995 B.n33 585
R1226 B.n1118 B.n33 585
R1227 B.n994 B.n993 585
R1228 B.n993 B.n29 585
R1229 B.n992 B.n28 585
R1230 B.n1124 B.n28 585
R1231 B.n991 B.n27 585
R1232 B.n1125 B.n27 585
R1233 B.n990 B.n26 585
R1234 B.n1126 B.n26 585
R1235 B.n989 B.n988 585
R1236 B.n988 B.n22 585
R1237 B.n987 B.n21 585
R1238 B.n1132 B.n21 585
R1239 B.n986 B.n20 585
R1240 B.n1133 B.n20 585
R1241 B.n985 B.n19 585
R1242 B.n1134 B.n19 585
R1243 B.n984 B.n983 585
R1244 B.n983 B.n15 585
R1245 B.n982 B.n14 585
R1246 B.n1140 B.n14 585
R1247 B.n981 B.n13 585
R1248 B.n1141 B.n13 585
R1249 B.n980 B.n12 585
R1250 B.n1142 B.n12 585
R1251 B.n979 B.n978 585
R1252 B.n978 B.n8 585
R1253 B.n977 B.n7 585
R1254 B.n1148 B.n7 585
R1255 B.n976 B.n6 585
R1256 B.n1149 B.n6 585
R1257 B.n975 B.n5 585
R1258 B.n1150 B.n5 585
R1259 B.n974 B.n973 585
R1260 B.n973 B.n4 585
R1261 B.n972 B.n404 585
R1262 B.n972 B.n971 585
R1263 B.n962 B.n405 585
R1264 B.n406 B.n405 585
R1265 B.n964 B.n963 585
R1266 B.n965 B.n964 585
R1267 B.n961 B.n411 585
R1268 B.n411 B.n410 585
R1269 B.n960 B.n959 585
R1270 B.n959 B.n958 585
R1271 B.n413 B.n412 585
R1272 B.n414 B.n413 585
R1273 B.n951 B.n950 585
R1274 B.n952 B.n951 585
R1275 B.n949 B.n419 585
R1276 B.n419 B.n418 585
R1277 B.n948 B.n947 585
R1278 B.n947 B.n946 585
R1279 B.n421 B.n420 585
R1280 B.n422 B.n421 585
R1281 B.n939 B.n938 585
R1282 B.n940 B.n939 585
R1283 B.n937 B.n426 585
R1284 B.n430 B.n426 585
R1285 B.n936 B.n935 585
R1286 B.n935 B.n934 585
R1287 B.n428 B.n427 585
R1288 B.n429 B.n428 585
R1289 B.n927 B.n926 585
R1290 B.n928 B.n927 585
R1291 B.n925 B.n435 585
R1292 B.n435 B.n434 585
R1293 B.n924 B.n923 585
R1294 B.n923 B.n922 585
R1295 B.n437 B.n436 585
R1296 B.n438 B.n437 585
R1297 B.n915 B.n914 585
R1298 B.n916 B.n915 585
R1299 B.n913 B.n442 585
R1300 B.n446 B.n442 585
R1301 B.n912 B.n911 585
R1302 B.n911 B.n910 585
R1303 B.n444 B.n443 585
R1304 B.n445 B.n444 585
R1305 B.n903 B.n902 585
R1306 B.n904 B.n903 585
R1307 B.n901 B.n451 585
R1308 B.n451 B.n450 585
R1309 B.n900 B.n899 585
R1310 B.n899 B.n898 585
R1311 B.n453 B.n452 585
R1312 B.n454 B.n453 585
R1313 B.n891 B.n890 585
R1314 B.n892 B.n891 585
R1315 B.n889 B.n459 585
R1316 B.n459 B.n458 585
R1317 B.n888 B.n887 585
R1318 B.n887 B.n886 585
R1319 B.n461 B.n460 585
R1320 B.n462 B.n461 585
R1321 B.n879 B.n878 585
R1322 B.n880 B.n879 585
R1323 B.n877 B.n467 585
R1324 B.n467 B.n466 585
R1325 B.n876 B.n875 585
R1326 B.n875 B.n874 585
R1327 B.n469 B.n468 585
R1328 B.n470 B.n469 585
R1329 B.n867 B.n866 585
R1330 B.n868 B.n867 585
R1331 B.n865 B.n475 585
R1332 B.n475 B.n474 585
R1333 B.n864 B.n863 585
R1334 B.n863 B.n862 585
R1335 B.n477 B.n476 585
R1336 B.n478 B.n477 585
R1337 B.n855 B.n854 585
R1338 B.n856 B.n855 585
R1339 B.n853 B.n483 585
R1340 B.n483 B.n482 585
R1341 B.n852 B.n851 585
R1342 B.n851 B.n850 585
R1343 B.n485 B.n484 585
R1344 B.n486 B.n485 585
R1345 B.n843 B.n842 585
R1346 B.n844 B.n843 585
R1347 B.n841 B.n491 585
R1348 B.n491 B.n490 585
R1349 B.n840 B.n839 585
R1350 B.n839 B.n838 585
R1351 B.n493 B.n492 585
R1352 B.n831 B.n493 585
R1353 B.n830 B.n829 585
R1354 B.n832 B.n830 585
R1355 B.n828 B.n498 585
R1356 B.n498 B.n497 585
R1357 B.n827 B.n826 585
R1358 B.n826 B.n825 585
R1359 B.n500 B.n499 585
R1360 B.n501 B.n500 585
R1361 B.n818 B.n817 585
R1362 B.n819 B.n818 585
R1363 B.n816 B.n506 585
R1364 B.n506 B.n505 585
R1365 B.n810 B.n809 585
R1366 B.n808 B.n568 585
R1367 B.n807 B.n567 585
R1368 B.n812 B.n567 585
R1369 B.n806 B.n805 585
R1370 B.n804 B.n803 585
R1371 B.n802 B.n801 585
R1372 B.n800 B.n799 585
R1373 B.n798 B.n797 585
R1374 B.n796 B.n795 585
R1375 B.n794 B.n793 585
R1376 B.n792 B.n791 585
R1377 B.n790 B.n789 585
R1378 B.n788 B.n787 585
R1379 B.n786 B.n785 585
R1380 B.n784 B.n783 585
R1381 B.n782 B.n781 585
R1382 B.n780 B.n779 585
R1383 B.n778 B.n777 585
R1384 B.n776 B.n775 585
R1385 B.n774 B.n773 585
R1386 B.n772 B.n771 585
R1387 B.n770 B.n769 585
R1388 B.n768 B.n767 585
R1389 B.n766 B.n765 585
R1390 B.n764 B.n763 585
R1391 B.n762 B.n761 585
R1392 B.n760 B.n759 585
R1393 B.n758 B.n757 585
R1394 B.n756 B.n755 585
R1395 B.n754 B.n753 585
R1396 B.n752 B.n751 585
R1397 B.n750 B.n749 585
R1398 B.n748 B.n747 585
R1399 B.n746 B.n745 585
R1400 B.n744 B.n743 585
R1401 B.n742 B.n741 585
R1402 B.n740 B.n739 585
R1403 B.n738 B.n737 585
R1404 B.n736 B.n735 585
R1405 B.n734 B.n733 585
R1406 B.n732 B.n731 585
R1407 B.n730 B.n729 585
R1408 B.n728 B.n727 585
R1409 B.n726 B.n725 585
R1410 B.n724 B.n723 585
R1411 B.n722 B.n721 585
R1412 B.n720 B.n719 585
R1413 B.n718 B.n717 585
R1414 B.n716 B.n715 585
R1415 B.n714 B.n713 585
R1416 B.n712 B.n711 585
R1417 B.n710 B.n709 585
R1418 B.n708 B.n707 585
R1419 B.n706 B.n705 585
R1420 B.n704 B.n703 585
R1421 B.n702 B.n701 585
R1422 B.n699 B.n698 585
R1423 B.n697 B.n696 585
R1424 B.n695 B.n694 585
R1425 B.n693 B.n692 585
R1426 B.n691 B.n690 585
R1427 B.n689 B.n688 585
R1428 B.n687 B.n686 585
R1429 B.n685 B.n684 585
R1430 B.n683 B.n682 585
R1431 B.n681 B.n680 585
R1432 B.n679 B.n678 585
R1433 B.n677 B.n676 585
R1434 B.n675 B.n674 585
R1435 B.n673 B.n672 585
R1436 B.n671 B.n670 585
R1437 B.n669 B.n668 585
R1438 B.n667 B.n666 585
R1439 B.n665 B.n664 585
R1440 B.n663 B.n662 585
R1441 B.n661 B.n660 585
R1442 B.n659 B.n658 585
R1443 B.n657 B.n656 585
R1444 B.n655 B.n654 585
R1445 B.n653 B.n652 585
R1446 B.n651 B.n650 585
R1447 B.n649 B.n648 585
R1448 B.n647 B.n646 585
R1449 B.n645 B.n644 585
R1450 B.n643 B.n642 585
R1451 B.n641 B.n640 585
R1452 B.n639 B.n638 585
R1453 B.n637 B.n636 585
R1454 B.n635 B.n634 585
R1455 B.n633 B.n632 585
R1456 B.n631 B.n630 585
R1457 B.n629 B.n628 585
R1458 B.n627 B.n626 585
R1459 B.n625 B.n624 585
R1460 B.n623 B.n622 585
R1461 B.n621 B.n620 585
R1462 B.n619 B.n618 585
R1463 B.n617 B.n616 585
R1464 B.n615 B.n614 585
R1465 B.n613 B.n612 585
R1466 B.n611 B.n610 585
R1467 B.n609 B.n608 585
R1468 B.n607 B.n606 585
R1469 B.n605 B.n604 585
R1470 B.n603 B.n602 585
R1471 B.n601 B.n600 585
R1472 B.n599 B.n598 585
R1473 B.n597 B.n596 585
R1474 B.n595 B.n594 585
R1475 B.n593 B.n592 585
R1476 B.n591 B.n590 585
R1477 B.n589 B.n588 585
R1478 B.n587 B.n586 585
R1479 B.n585 B.n584 585
R1480 B.n583 B.n582 585
R1481 B.n581 B.n580 585
R1482 B.n579 B.n578 585
R1483 B.n577 B.n576 585
R1484 B.n575 B.n574 585
R1485 B.n508 B.n507 585
R1486 B.n815 B.n814 585
R1487 B.n504 B.n503 585
R1488 B.n505 B.n504 585
R1489 B.n821 B.n820 585
R1490 B.n820 B.n819 585
R1491 B.n822 B.n502 585
R1492 B.n502 B.n501 585
R1493 B.n824 B.n823 585
R1494 B.n825 B.n824 585
R1495 B.n496 B.n495 585
R1496 B.n497 B.n496 585
R1497 B.n834 B.n833 585
R1498 B.n833 B.n832 585
R1499 B.n835 B.n494 585
R1500 B.n831 B.n494 585
R1501 B.n837 B.n836 585
R1502 B.n838 B.n837 585
R1503 B.n489 B.n488 585
R1504 B.n490 B.n489 585
R1505 B.n846 B.n845 585
R1506 B.n845 B.n844 585
R1507 B.n847 B.n487 585
R1508 B.n487 B.n486 585
R1509 B.n849 B.n848 585
R1510 B.n850 B.n849 585
R1511 B.n481 B.n480 585
R1512 B.n482 B.n481 585
R1513 B.n858 B.n857 585
R1514 B.n857 B.n856 585
R1515 B.n859 B.n479 585
R1516 B.n479 B.n478 585
R1517 B.n861 B.n860 585
R1518 B.n862 B.n861 585
R1519 B.n473 B.n472 585
R1520 B.n474 B.n473 585
R1521 B.n870 B.n869 585
R1522 B.n869 B.n868 585
R1523 B.n871 B.n471 585
R1524 B.n471 B.n470 585
R1525 B.n873 B.n872 585
R1526 B.n874 B.n873 585
R1527 B.n465 B.n464 585
R1528 B.n466 B.n465 585
R1529 B.n882 B.n881 585
R1530 B.n881 B.n880 585
R1531 B.n883 B.n463 585
R1532 B.n463 B.n462 585
R1533 B.n885 B.n884 585
R1534 B.n886 B.n885 585
R1535 B.n457 B.n456 585
R1536 B.n458 B.n457 585
R1537 B.n894 B.n893 585
R1538 B.n893 B.n892 585
R1539 B.n895 B.n455 585
R1540 B.n455 B.n454 585
R1541 B.n897 B.n896 585
R1542 B.n898 B.n897 585
R1543 B.n449 B.n448 585
R1544 B.n450 B.n449 585
R1545 B.n906 B.n905 585
R1546 B.n905 B.n904 585
R1547 B.n907 B.n447 585
R1548 B.n447 B.n445 585
R1549 B.n909 B.n908 585
R1550 B.n910 B.n909 585
R1551 B.n441 B.n440 585
R1552 B.n446 B.n441 585
R1553 B.n918 B.n917 585
R1554 B.n917 B.n916 585
R1555 B.n919 B.n439 585
R1556 B.n439 B.n438 585
R1557 B.n921 B.n920 585
R1558 B.n922 B.n921 585
R1559 B.n433 B.n432 585
R1560 B.n434 B.n433 585
R1561 B.n930 B.n929 585
R1562 B.n929 B.n928 585
R1563 B.n931 B.n431 585
R1564 B.n431 B.n429 585
R1565 B.n933 B.n932 585
R1566 B.n934 B.n933 585
R1567 B.n425 B.n424 585
R1568 B.n430 B.n425 585
R1569 B.n942 B.n941 585
R1570 B.n941 B.n940 585
R1571 B.n943 B.n423 585
R1572 B.n423 B.n422 585
R1573 B.n945 B.n944 585
R1574 B.n946 B.n945 585
R1575 B.n417 B.n416 585
R1576 B.n418 B.n417 585
R1577 B.n954 B.n953 585
R1578 B.n953 B.n952 585
R1579 B.n955 B.n415 585
R1580 B.n415 B.n414 585
R1581 B.n957 B.n956 585
R1582 B.n958 B.n957 585
R1583 B.n409 B.n408 585
R1584 B.n410 B.n409 585
R1585 B.n967 B.n966 585
R1586 B.n966 B.n965 585
R1587 B.n968 B.n407 585
R1588 B.n407 B.n406 585
R1589 B.n970 B.n969 585
R1590 B.n971 B.n970 585
R1591 B.n2 B.n0 585
R1592 B.n4 B.n2 585
R1593 B.n3 B.n1 585
R1594 B.n1149 B.n3 585
R1595 B.n1147 B.n1146 585
R1596 B.n1148 B.n1147 585
R1597 B.n1145 B.n9 585
R1598 B.n9 B.n8 585
R1599 B.n1144 B.n1143 585
R1600 B.n1143 B.n1142 585
R1601 B.n11 B.n10 585
R1602 B.n1141 B.n11 585
R1603 B.n1139 B.n1138 585
R1604 B.n1140 B.n1139 585
R1605 B.n1137 B.n16 585
R1606 B.n16 B.n15 585
R1607 B.n1136 B.n1135 585
R1608 B.n1135 B.n1134 585
R1609 B.n18 B.n17 585
R1610 B.n1133 B.n18 585
R1611 B.n1131 B.n1130 585
R1612 B.n1132 B.n1131 585
R1613 B.n1129 B.n23 585
R1614 B.n23 B.n22 585
R1615 B.n1128 B.n1127 585
R1616 B.n1127 B.n1126 585
R1617 B.n25 B.n24 585
R1618 B.n1125 B.n25 585
R1619 B.n1123 B.n1122 585
R1620 B.n1124 B.n1123 585
R1621 B.n1121 B.n30 585
R1622 B.n30 B.n29 585
R1623 B.n1120 B.n1119 585
R1624 B.n1119 B.n1118 585
R1625 B.n32 B.n31 585
R1626 B.n1117 B.n32 585
R1627 B.n1115 B.n1114 585
R1628 B.n1116 B.n1115 585
R1629 B.n1113 B.n37 585
R1630 B.n37 B.n36 585
R1631 B.n1112 B.n1111 585
R1632 B.n1111 B.n1110 585
R1633 B.n39 B.n38 585
R1634 B.n1109 B.n39 585
R1635 B.n1107 B.n1106 585
R1636 B.n1108 B.n1107 585
R1637 B.n1105 B.n44 585
R1638 B.n44 B.n43 585
R1639 B.n1104 B.n1103 585
R1640 B.n1103 B.n1102 585
R1641 B.n46 B.n45 585
R1642 B.n1101 B.n46 585
R1643 B.n1099 B.n1098 585
R1644 B.n1100 B.n1099 585
R1645 B.n1097 B.n51 585
R1646 B.n51 B.n50 585
R1647 B.n1096 B.n1095 585
R1648 B.n1095 B.n1094 585
R1649 B.n53 B.n52 585
R1650 B.n1093 B.n53 585
R1651 B.n1091 B.n1090 585
R1652 B.n1092 B.n1091 585
R1653 B.n1089 B.n58 585
R1654 B.n58 B.n57 585
R1655 B.n1088 B.n1087 585
R1656 B.n1087 B.n1086 585
R1657 B.n60 B.n59 585
R1658 B.n1085 B.n60 585
R1659 B.n1083 B.n1082 585
R1660 B.n1084 B.n1083 585
R1661 B.n1081 B.n65 585
R1662 B.n65 B.n64 585
R1663 B.n1080 B.n1079 585
R1664 B.n1079 B.n1078 585
R1665 B.n67 B.n66 585
R1666 B.n1077 B.n67 585
R1667 B.n1075 B.n1074 585
R1668 B.n1076 B.n1075 585
R1669 B.n1073 B.n72 585
R1670 B.n72 B.n71 585
R1671 B.n1072 B.n1071 585
R1672 B.n1071 B.n1070 585
R1673 B.n74 B.n73 585
R1674 B.n1069 B.n74 585
R1675 B.n1067 B.n1066 585
R1676 B.n1068 B.n1067 585
R1677 B.n1065 B.n79 585
R1678 B.n79 B.n78 585
R1679 B.n1064 B.n1063 585
R1680 B.n1063 B.n1062 585
R1681 B.n81 B.n80 585
R1682 B.n1061 B.n81 585
R1683 B.n1059 B.n1058 585
R1684 B.n1060 B.n1059 585
R1685 B.n1057 B.n85 585
R1686 B.n88 B.n85 585
R1687 B.n1056 B.n1055 585
R1688 B.n1055 B.n1054 585
R1689 B.n87 B.n86 585
R1690 B.n1053 B.n87 585
R1691 B.n1051 B.n1050 585
R1692 B.n1052 B.n1051 585
R1693 B.n1049 B.n93 585
R1694 B.n93 B.n92 585
R1695 B.n1048 B.n1047 585
R1696 B.n1047 B.n1046 585
R1697 B.n95 B.n94 585
R1698 B.n1045 B.n95 585
R1699 B.n1152 B.n1151 585
R1700 B.n1151 B.n1150 585
R1701 B.n810 B.n504 554.963
R1702 B.n164 B.n95 554.963
R1703 B.n814 B.n506 554.963
R1704 B.n1043 B.n97 554.963
R1705 B.n571 B.t13 415.582
R1706 B.n159 B.t16 415.582
R1707 B.n569 B.t20 415.582
R1708 B.n161 B.t22 415.582
R1709 B.n571 B.t10 390.529
R1710 B.n569 B.t18 390.529
R1711 B.n161 B.t21 390.529
R1712 B.n159 B.t14 390.529
R1713 B.n572 B.t12 366.128
R1714 B.n160 B.t17 366.128
R1715 B.n570 B.t19 366.128
R1716 B.n162 B.t23 366.128
R1717 B.n1044 B.n157 256.663
R1718 B.n1044 B.n156 256.663
R1719 B.n1044 B.n155 256.663
R1720 B.n1044 B.n154 256.663
R1721 B.n1044 B.n153 256.663
R1722 B.n1044 B.n152 256.663
R1723 B.n1044 B.n151 256.663
R1724 B.n1044 B.n150 256.663
R1725 B.n1044 B.n149 256.663
R1726 B.n1044 B.n148 256.663
R1727 B.n1044 B.n147 256.663
R1728 B.n1044 B.n146 256.663
R1729 B.n1044 B.n145 256.663
R1730 B.n1044 B.n144 256.663
R1731 B.n1044 B.n143 256.663
R1732 B.n1044 B.n142 256.663
R1733 B.n1044 B.n141 256.663
R1734 B.n1044 B.n140 256.663
R1735 B.n1044 B.n139 256.663
R1736 B.n1044 B.n138 256.663
R1737 B.n1044 B.n137 256.663
R1738 B.n1044 B.n136 256.663
R1739 B.n1044 B.n135 256.663
R1740 B.n1044 B.n134 256.663
R1741 B.n1044 B.n133 256.663
R1742 B.n1044 B.n132 256.663
R1743 B.n1044 B.n131 256.663
R1744 B.n1044 B.n130 256.663
R1745 B.n1044 B.n129 256.663
R1746 B.n1044 B.n128 256.663
R1747 B.n1044 B.n127 256.663
R1748 B.n1044 B.n126 256.663
R1749 B.n1044 B.n125 256.663
R1750 B.n1044 B.n124 256.663
R1751 B.n1044 B.n123 256.663
R1752 B.n1044 B.n122 256.663
R1753 B.n1044 B.n121 256.663
R1754 B.n1044 B.n120 256.663
R1755 B.n1044 B.n119 256.663
R1756 B.n1044 B.n118 256.663
R1757 B.n1044 B.n117 256.663
R1758 B.n1044 B.n116 256.663
R1759 B.n1044 B.n115 256.663
R1760 B.n1044 B.n114 256.663
R1761 B.n1044 B.n113 256.663
R1762 B.n1044 B.n112 256.663
R1763 B.n1044 B.n111 256.663
R1764 B.n1044 B.n110 256.663
R1765 B.n1044 B.n109 256.663
R1766 B.n1044 B.n108 256.663
R1767 B.n1044 B.n107 256.663
R1768 B.n1044 B.n106 256.663
R1769 B.n1044 B.n105 256.663
R1770 B.n1044 B.n104 256.663
R1771 B.n1044 B.n103 256.663
R1772 B.n1044 B.n102 256.663
R1773 B.n1044 B.n101 256.663
R1774 B.n1044 B.n100 256.663
R1775 B.n1044 B.n99 256.663
R1776 B.n1044 B.n98 256.663
R1777 B.n812 B.n811 256.663
R1778 B.n812 B.n509 256.663
R1779 B.n812 B.n510 256.663
R1780 B.n812 B.n511 256.663
R1781 B.n812 B.n512 256.663
R1782 B.n812 B.n513 256.663
R1783 B.n812 B.n514 256.663
R1784 B.n812 B.n515 256.663
R1785 B.n812 B.n516 256.663
R1786 B.n812 B.n517 256.663
R1787 B.n812 B.n518 256.663
R1788 B.n812 B.n519 256.663
R1789 B.n812 B.n520 256.663
R1790 B.n812 B.n521 256.663
R1791 B.n812 B.n522 256.663
R1792 B.n812 B.n523 256.663
R1793 B.n812 B.n524 256.663
R1794 B.n812 B.n525 256.663
R1795 B.n812 B.n526 256.663
R1796 B.n812 B.n527 256.663
R1797 B.n812 B.n528 256.663
R1798 B.n812 B.n529 256.663
R1799 B.n812 B.n530 256.663
R1800 B.n812 B.n531 256.663
R1801 B.n812 B.n532 256.663
R1802 B.n812 B.n533 256.663
R1803 B.n812 B.n534 256.663
R1804 B.n812 B.n535 256.663
R1805 B.n812 B.n536 256.663
R1806 B.n812 B.n537 256.663
R1807 B.n812 B.n538 256.663
R1808 B.n812 B.n539 256.663
R1809 B.n812 B.n540 256.663
R1810 B.n812 B.n541 256.663
R1811 B.n812 B.n542 256.663
R1812 B.n812 B.n543 256.663
R1813 B.n812 B.n544 256.663
R1814 B.n812 B.n545 256.663
R1815 B.n812 B.n546 256.663
R1816 B.n812 B.n547 256.663
R1817 B.n812 B.n548 256.663
R1818 B.n812 B.n549 256.663
R1819 B.n812 B.n550 256.663
R1820 B.n812 B.n551 256.663
R1821 B.n812 B.n552 256.663
R1822 B.n812 B.n553 256.663
R1823 B.n812 B.n554 256.663
R1824 B.n812 B.n555 256.663
R1825 B.n812 B.n556 256.663
R1826 B.n812 B.n557 256.663
R1827 B.n812 B.n558 256.663
R1828 B.n812 B.n559 256.663
R1829 B.n812 B.n560 256.663
R1830 B.n812 B.n561 256.663
R1831 B.n812 B.n562 256.663
R1832 B.n812 B.n563 256.663
R1833 B.n812 B.n564 256.663
R1834 B.n812 B.n565 256.663
R1835 B.n812 B.n566 256.663
R1836 B.n813 B.n812 256.663
R1837 B.n820 B.n504 163.367
R1838 B.n820 B.n502 163.367
R1839 B.n824 B.n502 163.367
R1840 B.n824 B.n496 163.367
R1841 B.n833 B.n496 163.367
R1842 B.n833 B.n494 163.367
R1843 B.n837 B.n494 163.367
R1844 B.n837 B.n489 163.367
R1845 B.n845 B.n489 163.367
R1846 B.n845 B.n487 163.367
R1847 B.n849 B.n487 163.367
R1848 B.n849 B.n481 163.367
R1849 B.n857 B.n481 163.367
R1850 B.n857 B.n479 163.367
R1851 B.n861 B.n479 163.367
R1852 B.n861 B.n473 163.367
R1853 B.n869 B.n473 163.367
R1854 B.n869 B.n471 163.367
R1855 B.n873 B.n471 163.367
R1856 B.n873 B.n465 163.367
R1857 B.n881 B.n465 163.367
R1858 B.n881 B.n463 163.367
R1859 B.n885 B.n463 163.367
R1860 B.n885 B.n457 163.367
R1861 B.n893 B.n457 163.367
R1862 B.n893 B.n455 163.367
R1863 B.n897 B.n455 163.367
R1864 B.n897 B.n449 163.367
R1865 B.n905 B.n449 163.367
R1866 B.n905 B.n447 163.367
R1867 B.n909 B.n447 163.367
R1868 B.n909 B.n441 163.367
R1869 B.n917 B.n441 163.367
R1870 B.n917 B.n439 163.367
R1871 B.n921 B.n439 163.367
R1872 B.n921 B.n433 163.367
R1873 B.n929 B.n433 163.367
R1874 B.n929 B.n431 163.367
R1875 B.n933 B.n431 163.367
R1876 B.n933 B.n425 163.367
R1877 B.n941 B.n425 163.367
R1878 B.n941 B.n423 163.367
R1879 B.n945 B.n423 163.367
R1880 B.n945 B.n417 163.367
R1881 B.n953 B.n417 163.367
R1882 B.n953 B.n415 163.367
R1883 B.n957 B.n415 163.367
R1884 B.n957 B.n409 163.367
R1885 B.n966 B.n409 163.367
R1886 B.n966 B.n407 163.367
R1887 B.n970 B.n407 163.367
R1888 B.n970 B.n2 163.367
R1889 B.n1151 B.n2 163.367
R1890 B.n1151 B.n3 163.367
R1891 B.n1147 B.n3 163.367
R1892 B.n1147 B.n9 163.367
R1893 B.n1143 B.n9 163.367
R1894 B.n1143 B.n11 163.367
R1895 B.n1139 B.n11 163.367
R1896 B.n1139 B.n16 163.367
R1897 B.n1135 B.n16 163.367
R1898 B.n1135 B.n18 163.367
R1899 B.n1131 B.n18 163.367
R1900 B.n1131 B.n23 163.367
R1901 B.n1127 B.n23 163.367
R1902 B.n1127 B.n25 163.367
R1903 B.n1123 B.n25 163.367
R1904 B.n1123 B.n30 163.367
R1905 B.n1119 B.n30 163.367
R1906 B.n1119 B.n32 163.367
R1907 B.n1115 B.n32 163.367
R1908 B.n1115 B.n37 163.367
R1909 B.n1111 B.n37 163.367
R1910 B.n1111 B.n39 163.367
R1911 B.n1107 B.n39 163.367
R1912 B.n1107 B.n44 163.367
R1913 B.n1103 B.n44 163.367
R1914 B.n1103 B.n46 163.367
R1915 B.n1099 B.n46 163.367
R1916 B.n1099 B.n51 163.367
R1917 B.n1095 B.n51 163.367
R1918 B.n1095 B.n53 163.367
R1919 B.n1091 B.n53 163.367
R1920 B.n1091 B.n58 163.367
R1921 B.n1087 B.n58 163.367
R1922 B.n1087 B.n60 163.367
R1923 B.n1083 B.n60 163.367
R1924 B.n1083 B.n65 163.367
R1925 B.n1079 B.n65 163.367
R1926 B.n1079 B.n67 163.367
R1927 B.n1075 B.n67 163.367
R1928 B.n1075 B.n72 163.367
R1929 B.n1071 B.n72 163.367
R1930 B.n1071 B.n74 163.367
R1931 B.n1067 B.n74 163.367
R1932 B.n1067 B.n79 163.367
R1933 B.n1063 B.n79 163.367
R1934 B.n1063 B.n81 163.367
R1935 B.n1059 B.n81 163.367
R1936 B.n1059 B.n85 163.367
R1937 B.n1055 B.n85 163.367
R1938 B.n1055 B.n87 163.367
R1939 B.n1051 B.n87 163.367
R1940 B.n1051 B.n93 163.367
R1941 B.n1047 B.n93 163.367
R1942 B.n1047 B.n95 163.367
R1943 B.n568 B.n567 163.367
R1944 B.n805 B.n567 163.367
R1945 B.n803 B.n802 163.367
R1946 B.n799 B.n798 163.367
R1947 B.n795 B.n794 163.367
R1948 B.n791 B.n790 163.367
R1949 B.n787 B.n786 163.367
R1950 B.n783 B.n782 163.367
R1951 B.n779 B.n778 163.367
R1952 B.n775 B.n774 163.367
R1953 B.n771 B.n770 163.367
R1954 B.n767 B.n766 163.367
R1955 B.n763 B.n762 163.367
R1956 B.n759 B.n758 163.367
R1957 B.n755 B.n754 163.367
R1958 B.n751 B.n750 163.367
R1959 B.n747 B.n746 163.367
R1960 B.n743 B.n742 163.367
R1961 B.n739 B.n738 163.367
R1962 B.n735 B.n734 163.367
R1963 B.n731 B.n730 163.367
R1964 B.n727 B.n726 163.367
R1965 B.n723 B.n722 163.367
R1966 B.n719 B.n718 163.367
R1967 B.n715 B.n714 163.367
R1968 B.n711 B.n710 163.367
R1969 B.n707 B.n706 163.367
R1970 B.n703 B.n702 163.367
R1971 B.n698 B.n697 163.367
R1972 B.n694 B.n693 163.367
R1973 B.n690 B.n689 163.367
R1974 B.n686 B.n685 163.367
R1975 B.n682 B.n681 163.367
R1976 B.n678 B.n677 163.367
R1977 B.n674 B.n673 163.367
R1978 B.n670 B.n669 163.367
R1979 B.n666 B.n665 163.367
R1980 B.n662 B.n661 163.367
R1981 B.n658 B.n657 163.367
R1982 B.n654 B.n653 163.367
R1983 B.n650 B.n649 163.367
R1984 B.n646 B.n645 163.367
R1985 B.n642 B.n641 163.367
R1986 B.n638 B.n637 163.367
R1987 B.n634 B.n633 163.367
R1988 B.n630 B.n629 163.367
R1989 B.n626 B.n625 163.367
R1990 B.n622 B.n621 163.367
R1991 B.n618 B.n617 163.367
R1992 B.n614 B.n613 163.367
R1993 B.n610 B.n609 163.367
R1994 B.n606 B.n605 163.367
R1995 B.n602 B.n601 163.367
R1996 B.n598 B.n597 163.367
R1997 B.n594 B.n593 163.367
R1998 B.n590 B.n589 163.367
R1999 B.n586 B.n585 163.367
R2000 B.n582 B.n581 163.367
R2001 B.n578 B.n577 163.367
R2002 B.n574 B.n508 163.367
R2003 B.n818 B.n506 163.367
R2004 B.n818 B.n500 163.367
R2005 B.n826 B.n500 163.367
R2006 B.n826 B.n498 163.367
R2007 B.n830 B.n498 163.367
R2008 B.n830 B.n493 163.367
R2009 B.n839 B.n493 163.367
R2010 B.n839 B.n491 163.367
R2011 B.n843 B.n491 163.367
R2012 B.n843 B.n485 163.367
R2013 B.n851 B.n485 163.367
R2014 B.n851 B.n483 163.367
R2015 B.n855 B.n483 163.367
R2016 B.n855 B.n477 163.367
R2017 B.n863 B.n477 163.367
R2018 B.n863 B.n475 163.367
R2019 B.n867 B.n475 163.367
R2020 B.n867 B.n469 163.367
R2021 B.n875 B.n469 163.367
R2022 B.n875 B.n467 163.367
R2023 B.n879 B.n467 163.367
R2024 B.n879 B.n461 163.367
R2025 B.n887 B.n461 163.367
R2026 B.n887 B.n459 163.367
R2027 B.n891 B.n459 163.367
R2028 B.n891 B.n453 163.367
R2029 B.n899 B.n453 163.367
R2030 B.n899 B.n451 163.367
R2031 B.n903 B.n451 163.367
R2032 B.n903 B.n444 163.367
R2033 B.n911 B.n444 163.367
R2034 B.n911 B.n442 163.367
R2035 B.n915 B.n442 163.367
R2036 B.n915 B.n437 163.367
R2037 B.n923 B.n437 163.367
R2038 B.n923 B.n435 163.367
R2039 B.n927 B.n435 163.367
R2040 B.n927 B.n428 163.367
R2041 B.n935 B.n428 163.367
R2042 B.n935 B.n426 163.367
R2043 B.n939 B.n426 163.367
R2044 B.n939 B.n421 163.367
R2045 B.n947 B.n421 163.367
R2046 B.n947 B.n419 163.367
R2047 B.n951 B.n419 163.367
R2048 B.n951 B.n413 163.367
R2049 B.n959 B.n413 163.367
R2050 B.n959 B.n411 163.367
R2051 B.n964 B.n411 163.367
R2052 B.n964 B.n405 163.367
R2053 B.n972 B.n405 163.367
R2054 B.n973 B.n972 163.367
R2055 B.n973 B.n5 163.367
R2056 B.n6 B.n5 163.367
R2057 B.n7 B.n6 163.367
R2058 B.n978 B.n7 163.367
R2059 B.n978 B.n12 163.367
R2060 B.n13 B.n12 163.367
R2061 B.n14 B.n13 163.367
R2062 B.n983 B.n14 163.367
R2063 B.n983 B.n19 163.367
R2064 B.n20 B.n19 163.367
R2065 B.n21 B.n20 163.367
R2066 B.n988 B.n21 163.367
R2067 B.n988 B.n26 163.367
R2068 B.n27 B.n26 163.367
R2069 B.n28 B.n27 163.367
R2070 B.n993 B.n28 163.367
R2071 B.n993 B.n33 163.367
R2072 B.n34 B.n33 163.367
R2073 B.n35 B.n34 163.367
R2074 B.n998 B.n35 163.367
R2075 B.n998 B.n40 163.367
R2076 B.n41 B.n40 163.367
R2077 B.n42 B.n41 163.367
R2078 B.n1003 B.n42 163.367
R2079 B.n1003 B.n47 163.367
R2080 B.n48 B.n47 163.367
R2081 B.n49 B.n48 163.367
R2082 B.n1008 B.n49 163.367
R2083 B.n1008 B.n54 163.367
R2084 B.n55 B.n54 163.367
R2085 B.n56 B.n55 163.367
R2086 B.n1013 B.n56 163.367
R2087 B.n1013 B.n61 163.367
R2088 B.n62 B.n61 163.367
R2089 B.n63 B.n62 163.367
R2090 B.n1018 B.n63 163.367
R2091 B.n1018 B.n68 163.367
R2092 B.n69 B.n68 163.367
R2093 B.n70 B.n69 163.367
R2094 B.n1023 B.n70 163.367
R2095 B.n1023 B.n75 163.367
R2096 B.n76 B.n75 163.367
R2097 B.n77 B.n76 163.367
R2098 B.n1028 B.n77 163.367
R2099 B.n1028 B.n82 163.367
R2100 B.n83 B.n82 163.367
R2101 B.n84 B.n83 163.367
R2102 B.n1033 B.n84 163.367
R2103 B.n1033 B.n89 163.367
R2104 B.n90 B.n89 163.367
R2105 B.n91 B.n90 163.367
R2106 B.n1038 B.n91 163.367
R2107 B.n1038 B.n96 163.367
R2108 B.n97 B.n96 163.367
R2109 B.n168 B.n167 163.367
R2110 B.n172 B.n171 163.367
R2111 B.n176 B.n175 163.367
R2112 B.n180 B.n179 163.367
R2113 B.n184 B.n183 163.367
R2114 B.n188 B.n187 163.367
R2115 B.n192 B.n191 163.367
R2116 B.n196 B.n195 163.367
R2117 B.n200 B.n199 163.367
R2118 B.n204 B.n203 163.367
R2119 B.n208 B.n207 163.367
R2120 B.n212 B.n211 163.367
R2121 B.n216 B.n215 163.367
R2122 B.n220 B.n219 163.367
R2123 B.n224 B.n223 163.367
R2124 B.n228 B.n227 163.367
R2125 B.n232 B.n231 163.367
R2126 B.n236 B.n235 163.367
R2127 B.n240 B.n239 163.367
R2128 B.n244 B.n243 163.367
R2129 B.n248 B.n247 163.367
R2130 B.n252 B.n251 163.367
R2131 B.n256 B.n255 163.367
R2132 B.n260 B.n259 163.367
R2133 B.n264 B.n263 163.367
R2134 B.n268 B.n267 163.367
R2135 B.n272 B.n271 163.367
R2136 B.n276 B.n275 163.367
R2137 B.n280 B.n279 163.367
R2138 B.n284 B.n283 163.367
R2139 B.n288 B.n287 163.367
R2140 B.n292 B.n291 163.367
R2141 B.n297 B.n296 163.367
R2142 B.n301 B.n300 163.367
R2143 B.n305 B.n304 163.367
R2144 B.n309 B.n308 163.367
R2145 B.n313 B.n312 163.367
R2146 B.n317 B.n316 163.367
R2147 B.n321 B.n320 163.367
R2148 B.n325 B.n324 163.367
R2149 B.n329 B.n328 163.367
R2150 B.n333 B.n332 163.367
R2151 B.n337 B.n336 163.367
R2152 B.n341 B.n340 163.367
R2153 B.n345 B.n344 163.367
R2154 B.n349 B.n348 163.367
R2155 B.n353 B.n352 163.367
R2156 B.n357 B.n356 163.367
R2157 B.n361 B.n360 163.367
R2158 B.n365 B.n364 163.367
R2159 B.n369 B.n368 163.367
R2160 B.n373 B.n372 163.367
R2161 B.n377 B.n376 163.367
R2162 B.n381 B.n380 163.367
R2163 B.n385 B.n384 163.367
R2164 B.n389 B.n388 163.367
R2165 B.n393 B.n392 163.367
R2166 B.n397 B.n396 163.367
R2167 B.n401 B.n400 163.367
R2168 B.n1043 B.n158 163.367
R2169 B.n811 B.n810 71.676
R2170 B.n805 B.n509 71.676
R2171 B.n802 B.n510 71.676
R2172 B.n798 B.n511 71.676
R2173 B.n794 B.n512 71.676
R2174 B.n790 B.n513 71.676
R2175 B.n786 B.n514 71.676
R2176 B.n782 B.n515 71.676
R2177 B.n778 B.n516 71.676
R2178 B.n774 B.n517 71.676
R2179 B.n770 B.n518 71.676
R2180 B.n766 B.n519 71.676
R2181 B.n762 B.n520 71.676
R2182 B.n758 B.n521 71.676
R2183 B.n754 B.n522 71.676
R2184 B.n750 B.n523 71.676
R2185 B.n746 B.n524 71.676
R2186 B.n742 B.n525 71.676
R2187 B.n738 B.n526 71.676
R2188 B.n734 B.n527 71.676
R2189 B.n730 B.n528 71.676
R2190 B.n726 B.n529 71.676
R2191 B.n722 B.n530 71.676
R2192 B.n718 B.n531 71.676
R2193 B.n714 B.n532 71.676
R2194 B.n710 B.n533 71.676
R2195 B.n706 B.n534 71.676
R2196 B.n702 B.n535 71.676
R2197 B.n697 B.n536 71.676
R2198 B.n693 B.n537 71.676
R2199 B.n689 B.n538 71.676
R2200 B.n685 B.n539 71.676
R2201 B.n681 B.n540 71.676
R2202 B.n677 B.n541 71.676
R2203 B.n673 B.n542 71.676
R2204 B.n669 B.n543 71.676
R2205 B.n665 B.n544 71.676
R2206 B.n661 B.n545 71.676
R2207 B.n657 B.n546 71.676
R2208 B.n653 B.n547 71.676
R2209 B.n649 B.n548 71.676
R2210 B.n645 B.n549 71.676
R2211 B.n641 B.n550 71.676
R2212 B.n637 B.n551 71.676
R2213 B.n633 B.n552 71.676
R2214 B.n629 B.n553 71.676
R2215 B.n625 B.n554 71.676
R2216 B.n621 B.n555 71.676
R2217 B.n617 B.n556 71.676
R2218 B.n613 B.n557 71.676
R2219 B.n609 B.n558 71.676
R2220 B.n605 B.n559 71.676
R2221 B.n601 B.n560 71.676
R2222 B.n597 B.n561 71.676
R2223 B.n593 B.n562 71.676
R2224 B.n589 B.n563 71.676
R2225 B.n585 B.n564 71.676
R2226 B.n581 B.n565 71.676
R2227 B.n577 B.n566 71.676
R2228 B.n813 B.n508 71.676
R2229 B.n164 B.n98 71.676
R2230 B.n168 B.n99 71.676
R2231 B.n172 B.n100 71.676
R2232 B.n176 B.n101 71.676
R2233 B.n180 B.n102 71.676
R2234 B.n184 B.n103 71.676
R2235 B.n188 B.n104 71.676
R2236 B.n192 B.n105 71.676
R2237 B.n196 B.n106 71.676
R2238 B.n200 B.n107 71.676
R2239 B.n204 B.n108 71.676
R2240 B.n208 B.n109 71.676
R2241 B.n212 B.n110 71.676
R2242 B.n216 B.n111 71.676
R2243 B.n220 B.n112 71.676
R2244 B.n224 B.n113 71.676
R2245 B.n228 B.n114 71.676
R2246 B.n232 B.n115 71.676
R2247 B.n236 B.n116 71.676
R2248 B.n240 B.n117 71.676
R2249 B.n244 B.n118 71.676
R2250 B.n248 B.n119 71.676
R2251 B.n252 B.n120 71.676
R2252 B.n256 B.n121 71.676
R2253 B.n260 B.n122 71.676
R2254 B.n264 B.n123 71.676
R2255 B.n268 B.n124 71.676
R2256 B.n272 B.n125 71.676
R2257 B.n276 B.n126 71.676
R2258 B.n280 B.n127 71.676
R2259 B.n284 B.n128 71.676
R2260 B.n288 B.n129 71.676
R2261 B.n292 B.n130 71.676
R2262 B.n297 B.n131 71.676
R2263 B.n301 B.n132 71.676
R2264 B.n305 B.n133 71.676
R2265 B.n309 B.n134 71.676
R2266 B.n313 B.n135 71.676
R2267 B.n317 B.n136 71.676
R2268 B.n321 B.n137 71.676
R2269 B.n325 B.n138 71.676
R2270 B.n329 B.n139 71.676
R2271 B.n333 B.n140 71.676
R2272 B.n337 B.n141 71.676
R2273 B.n341 B.n142 71.676
R2274 B.n345 B.n143 71.676
R2275 B.n349 B.n144 71.676
R2276 B.n353 B.n145 71.676
R2277 B.n357 B.n146 71.676
R2278 B.n361 B.n147 71.676
R2279 B.n365 B.n148 71.676
R2280 B.n369 B.n149 71.676
R2281 B.n373 B.n150 71.676
R2282 B.n377 B.n151 71.676
R2283 B.n381 B.n152 71.676
R2284 B.n385 B.n153 71.676
R2285 B.n389 B.n154 71.676
R2286 B.n393 B.n155 71.676
R2287 B.n397 B.n156 71.676
R2288 B.n401 B.n157 71.676
R2289 B.n158 B.n157 71.676
R2290 B.n400 B.n156 71.676
R2291 B.n396 B.n155 71.676
R2292 B.n392 B.n154 71.676
R2293 B.n388 B.n153 71.676
R2294 B.n384 B.n152 71.676
R2295 B.n380 B.n151 71.676
R2296 B.n376 B.n150 71.676
R2297 B.n372 B.n149 71.676
R2298 B.n368 B.n148 71.676
R2299 B.n364 B.n147 71.676
R2300 B.n360 B.n146 71.676
R2301 B.n356 B.n145 71.676
R2302 B.n352 B.n144 71.676
R2303 B.n348 B.n143 71.676
R2304 B.n344 B.n142 71.676
R2305 B.n340 B.n141 71.676
R2306 B.n336 B.n140 71.676
R2307 B.n332 B.n139 71.676
R2308 B.n328 B.n138 71.676
R2309 B.n324 B.n137 71.676
R2310 B.n320 B.n136 71.676
R2311 B.n316 B.n135 71.676
R2312 B.n312 B.n134 71.676
R2313 B.n308 B.n133 71.676
R2314 B.n304 B.n132 71.676
R2315 B.n300 B.n131 71.676
R2316 B.n296 B.n130 71.676
R2317 B.n291 B.n129 71.676
R2318 B.n287 B.n128 71.676
R2319 B.n283 B.n127 71.676
R2320 B.n279 B.n126 71.676
R2321 B.n275 B.n125 71.676
R2322 B.n271 B.n124 71.676
R2323 B.n267 B.n123 71.676
R2324 B.n263 B.n122 71.676
R2325 B.n259 B.n121 71.676
R2326 B.n255 B.n120 71.676
R2327 B.n251 B.n119 71.676
R2328 B.n247 B.n118 71.676
R2329 B.n243 B.n117 71.676
R2330 B.n239 B.n116 71.676
R2331 B.n235 B.n115 71.676
R2332 B.n231 B.n114 71.676
R2333 B.n227 B.n113 71.676
R2334 B.n223 B.n112 71.676
R2335 B.n219 B.n111 71.676
R2336 B.n215 B.n110 71.676
R2337 B.n211 B.n109 71.676
R2338 B.n207 B.n108 71.676
R2339 B.n203 B.n107 71.676
R2340 B.n199 B.n106 71.676
R2341 B.n195 B.n105 71.676
R2342 B.n191 B.n104 71.676
R2343 B.n187 B.n103 71.676
R2344 B.n183 B.n102 71.676
R2345 B.n179 B.n101 71.676
R2346 B.n175 B.n100 71.676
R2347 B.n171 B.n99 71.676
R2348 B.n167 B.n98 71.676
R2349 B.n811 B.n568 71.676
R2350 B.n803 B.n509 71.676
R2351 B.n799 B.n510 71.676
R2352 B.n795 B.n511 71.676
R2353 B.n791 B.n512 71.676
R2354 B.n787 B.n513 71.676
R2355 B.n783 B.n514 71.676
R2356 B.n779 B.n515 71.676
R2357 B.n775 B.n516 71.676
R2358 B.n771 B.n517 71.676
R2359 B.n767 B.n518 71.676
R2360 B.n763 B.n519 71.676
R2361 B.n759 B.n520 71.676
R2362 B.n755 B.n521 71.676
R2363 B.n751 B.n522 71.676
R2364 B.n747 B.n523 71.676
R2365 B.n743 B.n524 71.676
R2366 B.n739 B.n525 71.676
R2367 B.n735 B.n526 71.676
R2368 B.n731 B.n527 71.676
R2369 B.n727 B.n528 71.676
R2370 B.n723 B.n529 71.676
R2371 B.n719 B.n530 71.676
R2372 B.n715 B.n531 71.676
R2373 B.n711 B.n532 71.676
R2374 B.n707 B.n533 71.676
R2375 B.n703 B.n534 71.676
R2376 B.n698 B.n535 71.676
R2377 B.n694 B.n536 71.676
R2378 B.n690 B.n537 71.676
R2379 B.n686 B.n538 71.676
R2380 B.n682 B.n539 71.676
R2381 B.n678 B.n540 71.676
R2382 B.n674 B.n541 71.676
R2383 B.n670 B.n542 71.676
R2384 B.n666 B.n543 71.676
R2385 B.n662 B.n544 71.676
R2386 B.n658 B.n545 71.676
R2387 B.n654 B.n546 71.676
R2388 B.n650 B.n547 71.676
R2389 B.n646 B.n548 71.676
R2390 B.n642 B.n549 71.676
R2391 B.n638 B.n550 71.676
R2392 B.n634 B.n551 71.676
R2393 B.n630 B.n552 71.676
R2394 B.n626 B.n553 71.676
R2395 B.n622 B.n554 71.676
R2396 B.n618 B.n555 71.676
R2397 B.n614 B.n556 71.676
R2398 B.n610 B.n557 71.676
R2399 B.n606 B.n558 71.676
R2400 B.n602 B.n559 71.676
R2401 B.n598 B.n560 71.676
R2402 B.n594 B.n561 71.676
R2403 B.n590 B.n562 71.676
R2404 B.n586 B.n563 71.676
R2405 B.n582 B.n564 71.676
R2406 B.n578 B.n565 71.676
R2407 B.n574 B.n566 71.676
R2408 B.n814 B.n813 71.676
R2409 B.n812 B.n505 65.0716
R2410 B.n1045 B.n1044 65.0716
R2411 B.n573 B.n572 59.5399
R2412 B.n700 B.n570 59.5399
R2413 B.n163 B.n162 59.5399
R2414 B.n294 B.n160 59.5399
R2415 B.n572 B.n571 49.455
R2416 B.n570 B.n569 49.455
R2417 B.n162 B.n161 49.455
R2418 B.n160 B.n159 49.455
R2419 B.n165 B.n94 36.059
R2420 B.n816 B.n815 36.059
R2421 B.n809 B.n503 36.059
R2422 B.n1042 B.n1041 36.059
R2423 B.n819 B.n505 33.7779
R2424 B.n819 B.n501 33.7779
R2425 B.n825 B.n501 33.7779
R2426 B.n825 B.n497 33.7779
R2427 B.n832 B.n497 33.7779
R2428 B.n832 B.n831 33.7779
R2429 B.n838 B.n490 33.7779
R2430 B.n844 B.n490 33.7779
R2431 B.n844 B.n486 33.7779
R2432 B.n850 B.n486 33.7779
R2433 B.n850 B.n482 33.7779
R2434 B.n856 B.n482 33.7779
R2435 B.n856 B.n478 33.7779
R2436 B.n862 B.n478 33.7779
R2437 B.n862 B.n474 33.7779
R2438 B.n868 B.n474 33.7779
R2439 B.n874 B.n470 33.7779
R2440 B.n874 B.n466 33.7779
R2441 B.n880 B.n466 33.7779
R2442 B.n880 B.n462 33.7779
R2443 B.n886 B.n462 33.7779
R2444 B.n886 B.n458 33.7779
R2445 B.n892 B.n458 33.7779
R2446 B.n898 B.n454 33.7779
R2447 B.n898 B.n450 33.7779
R2448 B.n904 B.n450 33.7779
R2449 B.n904 B.n445 33.7779
R2450 B.n910 B.n445 33.7779
R2451 B.n910 B.n446 33.7779
R2452 B.n916 B.n438 33.7779
R2453 B.n922 B.n438 33.7779
R2454 B.n922 B.n434 33.7779
R2455 B.n928 B.n434 33.7779
R2456 B.n928 B.n429 33.7779
R2457 B.n934 B.n429 33.7779
R2458 B.n934 B.n430 33.7779
R2459 B.n940 B.n422 33.7779
R2460 B.n946 B.n422 33.7779
R2461 B.n946 B.n418 33.7779
R2462 B.n952 B.n418 33.7779
R2463 B.n952 B.n414 33.7779
R2464 B.n958 B.n414 33.7779
R2465 B.n965 B.n410 33.7779
R2466 B.n965 B.n406 33.7779
R2467 B.n971 B.n406 33.7779
R2468 B.n971 B.n4 33.7779
R2469 B.n1150 B.n4 33.7779
R2470 B.n1150 B.n1149 33.7779
R2471 B.n1149 B.n1148 33.7779
R2472 B.n1148 B.n8 33.7779
R2473 B.n1142 B.n8 33.7779
R2474 B.n1142 B.n1141 33.7779
R2475 B.n1140 B.n15 33.7779
R2476 B.n1134 B.n15 33.7779
R2477 B.n1134 B.n1133 33.7779
R2478 B.n1133 B.n1132 33.7779
R2479 B.n1132 B.n22 33.7779
R2480 B.n1126 B.n22 33.7779
R2481 B.n1125 B.n1124 33.7779
R2482 B.n1124 B.n29 33.7779
R2483 B.n1118 B.n29 33.7779
R2484 B.n1118 B.n1117 33.7779
R2485 B.n1117 B.n1116 33.7779
R2486 B.n1116 B.n36 33.7779
R2487 B.n1110 B.n36 33.7779
R2488 B.n1109 B.n1108 33.7779
R2489 B.n1108 B.n43 33.7779
R2490 B.n1102 B.n43 33.7779
R2491 B.n1102 B.n1101 33.7779
R2492 B.n1101 B.n1100 33.7779
R2493 B.n1100 B.n50 33.7779
R2494 B.n1094 B.n1093 33.7779
R2495 B.n1093 B.n1092 33.7779
R2496 B.n1092 B.n57 33.7779
R2497 B.n1086 B.n57 33.7779
R2498 B.n1086 B.n1085 33.7779
R2499 B.n1085 B.n1084 33.7779
R2500 B.n1084 B.n64 33.7779
R2501 B.n1078 B.n1077 33.7779
R2502 B.n1077 B.n1076 33.7779
R2503 B.n1076 B.n71 33.7779
R2504 B.n1070 B.n71 33.7779
R2505 B.n1070 B.n1069 33.7779
R2506 B.n1069 B.n1068 33.7779
R2507 B.n1068 B.n78 33.7779
R2508 B.n1062 B.n78 33.7779
R2509 B.n1062 B.n1061 33.7779
R2510 B.n1061 B.n1060 33.7779
R2511 B.n1054 B.n88 33.7779
R2512 B.n1054 B.n1053 33.7779
R2513 B.n1053 B.n1052 33.7779
R2514 B.n1052 B.n92 33.7779
R2515 B.n1046 B.n92 33.7779
R2516 B.n1046 B.n1045 33.7779
R2517 B.n831 B.t11 31.791
R2518 B.n88 B.t15 31.791
R2519 B.t1 B.n454 28.8106
R2520 B.n940 B.t7 28.8106
R2521 B.n1126 B.t3 28.8106
R2522 B.t2 B.n50 28.8106
R2523 B.n868 B.t4 21.8564
R2524 B.n446 B.t6 21.8564
R2525 B.n958 B.t9 21.8564
R2526 B.t8 B.n1140 21.8564
R2527 B.t0 B.n1109 21.8564
R2528 B.n1078 B.t5 21.8564
R2529 B B.n1152 18.0485
R2530 B.t4 B.n470 11.9219
R2531 B.n916 B.t6 11.9219
R2532 B.t9 B.n410 11.9219
R2533 B.n1141 B.t8 11.9219
R2534 B.n1110 B.t0 11.9219
R2535 B.t5 B.n64 11.9219
R2536 B.n166 B.n165 10.6151
R2537 B.n169 B.n166 10.6151
R2538 B.n170 B.n169 10.6151
R2539 B.n173 B.n170 10.6151
R2540 B.n174 B.n173 10.6151
R2541 B.n177 B.n174 10.6151
R2542 B.n178 B.n177 10.6151
R2543 B.n181 B.n178 10.6151
R2544 B.n182 B.n181 10.6151
R2545 B.n185 B.n182 10.6151
R2546 B.n186 B.n185 10.6151
R2547 B.n189 B.n186 10.6151
R2548 B.n190 B.n189 10.6151
R2549 B.n193 B.n190 10.6151
R2550 B.n194 B.n193 10.6151
R2551 B.n197 B.n194 10.6151
R2552 B.n198 B.n197 10.6151
R2553 B.n201 B.n198 10.6151
R2554 B.n202 B.n201 10.6151
R2555 B.n205 B.n202 10.6151
R2556 B.n206 B.n205 10.6151
R2557 B.n209 B.n206 10.6151
R2558 B.n210 B.n209 10.6151
R2559 B.n213 B.n210 10.6151
R2560 B.n214 B.n213 10.6151
R2561 B.n217 B.n214 10.6151
R2562 B.n218 B.n217 10.6151
R2563 B.n221 B.n218 10.6151
R2564 B.n222 B.n221 10.6151
R2565 B.n225 B.n222 10.6151
R2566 B.n226 B.n225 10.6151
R2567 B.n229 B.n226 10.6151
R2568 B.n230 B.n229 10.6151
R2569 B.n233 B.n230 10.6151
R2570 B.n234 B.n233 10.6151
R2571 B.n237 B.n234 10.6151
R2572 B.n238 B.n237 10.6151
R2573 B.n241 B.n238 10.6151
R2574 B.n242 B.n241 10.6151
R2575 B.n245 B.n242 10.6151
R2576 B.n246 B.n245 10.6151
R2577 B.n249 B.n246 10.6151
R2578 B.n250 B.n249 10.6151
R2579 B.n253 B.n250 10.6151
R2580 B.n254 B.n253 10.6151
R2581 B.n257 B.n254 10.6151
R2582 B.n258 B.n257 10.6151
R2583 B.n261 B.n258 10.6151
R2584 B.n262 B.n261 10.6151
R2585 B.n265 B.n262 10.6151
R2586 B.n266 B.n265 10.6151
R2587 B.n269 B.n266 10.6151
R2588 B.n270 B.n269 10.6151
R2589 B.n273 B.n270 10.6151
R2590 B.n274 B.n273 10.6151
R2591 B.n278 B.n277 10.6151
R2592 B.n281 B.n278 10.6151
R2593 B.n282 B.n281 10.6151
R2594 B.n285 B.n282 10.6151
R2595 B.n286 B.n285 10.6151
R2596 B.n289 B.n286 10.6151
R2597 B.n290 B.n289 10.6151
R2598 B.n293 B.n290 10.6151
R2599 B.n298 B.n295 10.6151
R2600 B.n299 B.n298 10.6151
R2601 B.n302 B.n299 10.6151
R2602 B.n303 B.n302 10.6151
R2603 B.n306 B.n303 10.6151
R2604 B.n307 B.n306 10.6151
R2605 B.n310 B.n307 10.6151
R2606 B.n311 B.n310 10.6151
R2607 B.n314 B.n311 10.6151
R2608 B.n315 B.n314 10.6151
R2609 B.n318 B.n315 10.6151
R2610 B.n319 B.n318 10.6151
R2611 B.n322 B.n319 10.6151
R2612 B.n323 B.n322 10.6151
R2613 B.n326 B.n323 10.6151
R2614 B.n327 B.n326 10.6151
R2615 B.n330 B.n327 10.6151
R2616 B.n331 B.n330 10.6151
R2617 B.n334 B.n331 10.6151
R2618 B.n335 B.n334 10.6151
R2619 B.n338 B.n335 10.6151
R2620 B.n339 B.n338 10.6151
R2621 B.n342 B.n339 10.6151
R2622 B.n343 B.n342 10.6151
R2623 B.n346 B.n343 10.6151
R2624 B.n347 B.n346 10.6151
R2625 B.n350 B.n347 10.6151
R2626 B.n351 B.n350 10.6151
R2627 B.n354 B.n351 10.6151
R2628 B.n355 B.n354 10.6151
R2629 B.n358 B.n355 10.6151
R2630 B.n359 B.n358 10.6151
R2631 B.n362 B.n359 10.6151
R2632 B.n363 B.n362 10.6151
R2633 B.n366 B.n363 10.6151
R2634 B.n367 B.n366 10.6151
R2635 B.n370 B.n367 10.6151
R2636 B.n371 B.n370 10.6151
R2637 B.n374 B.n371 10.6151
R2638 B.n375 B.n374 10.6151
R2639 B.n378 B.n375 10.6151
R2640 B.n379 B.n378 10.6151
R2641 B.n382 B.n379 10.6151
R2642 B.n383 B.n382 10.6151
R2643 B.n386 B.n383 10.6151
R2644 B.n387 B.n386 10.6151
R2645 B.n390 B.n387 10.6151
R2646 B.n391 B.n390 10.6151
R2647 B.n394 B.n391 10.6151
R2648 B.n395 B.n394 10.6151
R2649 B.n398 B.n395 10.6151
R2650 B.n399 B.n398 10.6151
R2651 B.n402 B.n399 10.6151
R2652 B.n403 B.n402 10.6151
R2653 B.n1042 B.n403 10.6151
R2654 B.n817 B.n816 10.6151
R2655 B.n817 B.n499 10.6151
R2656 B.n827 B.n499 10.6151
R2657 B.n828 B.n827 10.6151
R2658 B.n829 B.n828 10.6151
R2659 B.n829 B.n492 10.6151
R2660 B.n840 B.n492 10.6151
R2661 B.n841 B.n840 10.6151
R2662 B.n842 B.n841 10.6151
R2663 B.n842 B.n484 10.6151
R2664 B.n852 B.n484 10.6151
R2665 B.n853 B.n852 10.6151
R2666 B.n854 B.n853 10.6151
R2667 B.n854 B.n476 10.6151
R2668 B.n864 B.n476 10.6151
R2669 B.n865 B.n864 10.6151
R2670 B.n866 B.n865 10.6151
R2671 B.n866 B.n468 10.6151
R2672 B.n876 B.n468 10.6151
R2673 B.n877 B.n876 10.6151
R2674 B.n878 B.n877 10.6151
R2675 B.n878 B.n460 10.6151
R2676 B.n888 B.n460 10.6151
R2677 B.n889 B.n888 10.6151
R2678 B.n890 B.n889 10.6151
R2679 B.n890 B.n452 10.6151
R2680 B.n900 B.n452 10.6151
R2681 B.n901 B.n900 10.6151
R2682 B.n902 B.n901 10.6151
R2683 B.n902 B.n443 10.6151
R2684 B.n912 B.n443 10.6151
R2685 B.n913 B.n912 10.6151
R2686 B.n914 B.n913 10.6151
R2687 B.n914 B.n436 10.6151
R2688 B.n924 B.n436 10.6151
R2689 B.n925 B.n924 10.6151
R2690 B.n926 B.n925 10.6151
R2691 B.n926 B.n427 10.6151
R2692 B.n936 B.n427 10.6151
R2693 B.n937 B.n936 10.6151
R2694 B.n938 B.n937 10.6151
R2695 B.n938 B.n420 10.6151
R2696 B.n948 B.n420 10.6151
R2697 B.n949 B.n948 10.6151
R2698 B.n950 B.n949 10.6151
R2699 B.n950 B.n412 10.6151
R2700 B.n960 B.n412 10.6151
R2701 B.n961 B.n960 10.6151
R2702 B.n963 B.n961 10.6151
R2703 B.n963 B.n962 10.6151
R2704 B.n962 B.n404 10.6151
R2705 B.n974 B.n404 10.6151
R2706 B.n975 B.n974 10.6151
R2707 B.n976 B.n975 10.6151
R2708 B.n977 B.n976 10.6151
R2709 B.n979 B.n977 10.6151
R2710 B.n980 B.n979 10.6151
R2711 B.n981 B.n980 10.6151
R2712 B.n982 B.n981 10.6151
R2713 B.n984 B.n982 10.6151
R2714 B.n985 B.n984 10.6151
R2715 B.n986 B.n985 10.6151
R2716 B.n987 B.n986 10.6151
R2717 B.n989 B.n987 10.6151
R2718 B.n990 B.n989 10.6151
R2719 B.n991 B.n990 10.6151
R2720 B.n992 B.n991 10.6151
R2721 B.n994 B.n992 10.6151
R2722 B.n995 B.n994 10.6151
R2723 B.n996 B.n995 10.6151
R2724 B.n997 B.n996 10.6151
R2725 B.n999 B.n997 10.6151
R2726 B.n1000 B.n999 10.6151
R2727 B.n1001 B.n1000 10.6151
R2728 B.n1002 B.n1001 10.6151
R2729 B.n1004 B.n1002 10.6151
R2730 B.n1005 B.n1004 10.6151
R2731 B.n1006 B.n1005 10.6151
R2732 B.n1007 B.n1006 10.6151
R2733 B.n1009 B.n1007 10.6151
R2734 B.n1010 B.n1009 10.6151
R2735 B.n1011 B.n1010 10.6151
R2736 B.n1012 B.n1011 10.6151
R2737 B.n1014 B.n1012 10.6151
R2738 B.n1015 B.n1014 10.6151
R2739 B.n1016 B.n1015 10.6151
R2740 B.n1017 B.n1016 10.6151
R2741 B.n1019 B.n1017 10.6151
R2742 B.n1020 B.n1019 10.6151
R2743 B.n1021 B.n1020 10.6151
R2744 B.n1022 B.n1021 10.6151
R2745 B.n1024 B.n1022 10.6151
R2746 B.n1025 B.n1024 10.6151
R2747 B.n1026 B.n1025 10.6151
R2748 B.n1027 B.n1026 10.6151
R2749 B.n1029 B.n1027 10.6151
R2750 B.n1030 B.n1029 10.6151
R2751 B.n1031 B.n1030 10.6151
R2752 B.n1032 B.n1031 10.6151
R2753 B.n1034 B.n1032 10.6151
R2754 B.n1035 B.n1034 10.6151
R2755 B.n1036 B.n1035 10.6151
R2756 B.n1037 B.n1036 10.6151
R2757 B.n1039 B.n1037 10.6151
R2758 B.n1040 B.n1039 10.6151
R2759 B.n1041 B.n1040 10.6151
R2760 B.n809 B.n808 10.6151
R2761 B.n808 B.n807 10.6151
R2762 B.n807 B.n806 10.6151
R2763 B.n806 B.n804 10.6151
R2764 B.n804 B.n801 10.6151
R2765 B.n801 B.n800 10.6151
R2766 B.n800 B.n797 10.6151
R2767 B.n797 B.n796 10.6151
R2768 B.n796 B.n793 10.6151
R2769 B.n793 B.n792 10.6151
R2770 B.n792 B.n789 10.6151
R2771 B.n789 B.n788 10.6151
R2772 B.n788 B.n785 10.6151
R2773 B.n785 B.n784 10.6151
R2774 B.n784 B.n781 10.6151
R2775 B.n781 B.n780 10.6151
R2776 B.n780 B.n777 10.6151
R2777 B.n777 B.n776 10.6151
R2778 B.n776 B.n773 10.6151
R2779 B.n773 B.n772 10.6151
R2780 B.n772 B.n769 10.6151
R2781 B.n769 B.n768 10.6151
R2782 B.n768 B.n765 10.6151
R2783 B.n765 B.n764 10.6151
R2784 B.n764 B.n761 10.6151
R2785 B.n761 B.n760 10.6151
R2786 B.n760 B.n757 10.6151
R2787 B.n757 B.n756 10.6151
R2788 B.n756 B.n753 10.6151
R2789 B.n753 B.n752 10.6151
R2790 B.n752 B.n749 10.6151
R2791 B.n749 B.n748 10.6151
R2792 B.n748 B.n745 10.6151
R2793 B.n745 B.n744 10.6151
R2794 B.n744 B.n741 10.6151
R2795 B.n741 B.n740 10.6151
R2796 B.n740 B.n737 10.6151
R2797 B.n737 B.n736 10.6151
R2798 B.n736 B.n733 10.6151
R2799 B.n733 B.n732 10.6151
R2800 B.n732 B.n729 10.6151
R2801 B.n729 B.n728 10.6151
R2802 B.n728 B.n725 10.6151
R2803 B.n725 B.n724 10.6151
R2804 B.n724 B.n721 10.6151
R2805 B.n721 B.n720 10.6151
R2806 B.n720 B.n717 10.6151
R2807 B.n717 B.n716 10.6151
R2808 B.n716 B.n713 10.6151
R2809 B.n713 B.n712 10.6151
R2810 B.n712 B.n709 10.6151
R2811 B.n709 B.n708 10.6151
R2812 B.n708 B.n705 10.6151
R2813 B.n705 B.n704 10.6151
R2814 B.n704 B.n701 10.6151
R2815 B.n699 B.n696 10.6151
R2816 B.n696 B.n695 10.6151
R2817 B.n695 B.n692 10.6151
R2818 B.n692 B.n691 10.6151
R2819 B.n691 B.n688 10.6151
R2820 B.n688 B.n687 10.6151
R2821 B.n687 B.n684 10.6151
R2822 B.n684 B.n683 10.6151
R2823 B.n680 B.n679 10.6151
R2824 B.n679 B.n676 10.6151
R2825 B.n676 B.n675 10.6151
R2826 B.n675 B.n672 10.6151
R2827 B.n672 B.n671 10.6151
R2828 B.n671 B.n668 10.6151
R2829 B.n668 B.n667 10.6151
R2830 B.n667 B.n664 10.6151
R2831 B.n664 B.n663 10.6151
R2832 B.n663 B.n660 10.6151
R2833 B.n660 B.n659 10.6151
R2834 B.n659 B.n656 10.6151
R2835 B.n656 B.n655 10.6151
R2836 B.n655 B.n652 10.6151
R2837 B.n652 B.n651 10.6151
R2838 B.n651 B.n648 10.6151
R2839 B.n648 B.n647 10.6151
R2840 B.n647 B.n644 10.6151
R2841 B.n644 B.n643 10.6151
R2842 B.n643 B.n640 10.6151
R2843 B.n640 B.n639 10.6151
R2844 B.n639 B.n636 10.6151
R2845 B.n636 B.n635 10.6151
R2846 B.n635 B.n632 10.6151
R2847 B.n632 B.n631 10.6151
R2848 B.n631 B.n628 10.6151
R2849 B.n628 B.n627 10.6151
R2850 B.n627 B.n624 10.6151
R2851 B.n624 B.n623 10.6151
R2852 B.n623 B.n620 10.6151
R2853 B.n620 B.n619 10.6151
R2854 B.n619 B.n616 10.6151
R2855 B.n616 B.n615 10.6151
R2856 B.n615 B.n612 10.6151
R2857 B.n612 B.n611 10.6151
R2858 B.n611 B.n608 10.6151
R2859 B.n608 B.n607 10.6151
R2860 B.n607 B.n604 10.6151
R2861 B.n604 B.n603 10.6151
R2862 B.n603 B.n600 10.6151
R2863 B.n600 B.n599 10.6151
R2864 B.n599 B.n596 10.6151
R2865 B.n596 B.n595 10.6151
R2866 B.n595 B.n592 10.6151
R2867 B.n592 B.n591 10.6151
R2868 B.n591 B.n588 10.6151
R2869 B.n588 B.n587 10.6151
R2870 B.n587 B.n584 10.6151
R2871 B.n584 B.n583 10.6151
R2872 B.n583 B.n580 10.6151
R2873 B.n580 B.n579 10.6151
R2874 B.n579 B.n576 10.6151
R2875 B.n576 B.n575 10.6151
R2876 B.n575 B.n507 10.6151
R2877 B.n815 B.n507 10.6151
R2878 B.n821 B.n503 10.6151
R2879 B.n822 B.n821 10.6151
R2880 B.n823 B.n822 10.6151
R2881 B.n823 B.n495 10.6151
R2882 B.n834 B.n495 10.6151
R2883 B.n835 B.n834 10.6151
R2884 B.n836 B.n835 10.6151
R2885 B.n836 B.n488 10.6151
R2886 B.n846 B.n488 10.6151
R2887 B.n847 B.n846 10.6151
R2888 B.n848 B.n847 10.6151
R2889 B.n848 B.n480 10.6151
R2890 B.n858 B.n480 10.6151
R2891 B.n859 B.n858 10.6151
R2892 B.n860 B.n859 10.6151
R2893 B.n860 B.n472 10.6151
R2894 B.n870 B.n472 10.6151
R2895 B.n871 B.n870 10.6151
R2896 B.n872 B.n871 10.6151
R2897 B.n872 B.n464 10.6151
R2898 B.n882 B.n464 10.6151
R2899 B.n883 B.n882 10.6151
R2900 B.n884 B.n883 10.6151
R2901 B.n884 B.n456 10.6151
R2902 B.n894 B.n456 10.6151
R2903 B.n895 B.n894 10.6151
R2904 B.n896 B.n895 10.6151
R2905 B.n896 B.n448 10.6151
R2906 B.n906 B.n448 10.6151
R2907 B.n907 B.n906 10.6151
R2908 B.n908 B.n907 10.6151
R2909 B.n908 B.n440 10.6151
R2910 B.n918 B.n440 10.6151
R2911 B.n919 B.n918 10.6151
R2912 B.n920 B.n919 10.6151
R2913 B.n920 B.n432 10.6151
R2914 B.n930 B.n432 10.6151
R2915 B.n931 B.n930 10.6151
R2916 B.n932 B.n931 10.6151
R2917 B.n932 B.n424 10.6151
R2918 B.n942 B.n424 10.6151
R2919 B.n943 B.n942 10.6151
R2920 B.n944 B.n943 10.6151
R2921 B.n944 B.n416 10.6151
R2922 B.n954 B.n416 10.6151
R2923 B.n955 B.n954 10.6151
R2924 B.n956 B.n955 10.6151
R2925 B.n956 B.n408 10.6151
R2926 B.n967 B.n408 10.6151
R2927 B.n968 B.n967 10.6151
R2928 B.n969 B.n968 10.6151
R2929 B.n969 B.n0 10.6151
R2930 B.n1146 B.n1 10.6151
R2931 B.n1146 B.n1145 10.6151
R2932 B.n1145 B.n1144 10.6151
R2933 B.n1144 B.n10 10.6151
R2934 B.n1138 B.n10 10.6151
R2935 B.n1138 B.n1137 10.6151
R2936 B.n1137 B.n1136 10.6151
R2937 B.n1136 B.n17 10.6151
R2938 B.n1130 B.n17 10.6151
R2939 B.n1130 B.n1129 10.6151
R2940 B.n1129 B.n1128 10.6151
R2941 B.n1128 B.n24 10.6151
R2942 B.n1122 B.n24 10.6151
R2943 B.n1122 B.n1121 10.6151
R2944 B.n1121 B.n1120 10.6151
R2945 B.n1120 B.n31 10.6151
R2946 B.n1114 B.n31 10.6151
R2947 B.n1114 B.n1113 10.6151
R2948 B.n1113 B.n1112 10.6151
R2949 B.n1112 B.n38 10.6151
R2950 B.n1106 B.n38 10.6151
R2951 B.n1106 B.n1105 10.6151
R2952 B.n1105 B.n1104 10.6151
R2953 B.n1104 B.n45 10.6151
R2954 B.n1098 B.n45 10.6151
R2955 B.n1098 B.n1097 10.6151
R2956 B.n1097 B.n1096 10.6151
R2957 B.n1096 B.n52 10.6151
R2958 B.n1090 B.n52 10.6151
R2959 B.n1090 B.n1089 10.6151
R2960 B.n1089 B.n1088 10.6151
R2961 B.n1088 B.n59 10.6151
R2962 B.n1082 B.n59 10.6151
R2963 B.n1082 B.n1081 10.6151
R2964 B.n1081 B.n1080 10.6151
R2965 B.n1080 B.n66 10.6151
R2966 B.n1074 B.n66 10.6151
R2967 B.n1074 B.n1073 10.6151
R2968 B.n1073 B.n1072 10.6151
R2969 B.n1072 B.n73 10.6151
R2970 B.n1066 B.n73 10.6151
R2971 B.n1066 B.n1065 10.6151
R2972 B.n1065 B.n1064 10.6151
R2973 B.n1064 B.n80 10.6151
R2974 B.n1058 B.n80 10.6151
R2975 B.n1058 B.n1057 10.6151
R2976 B.n1057 B.n1056 10.6151
R2977 B.n1056 B.n86 10.6151
R2978 B.n1050 B.n86 10.6151
R2979 B.n1050 B.n1049 10.6151
R2980 B.n1049 B.n1048 10.6151
R2981 B.n1048 B.n94 10.6151
R2982 B.n277 B.n163 6.5566
R2983 B.n294 B.n293 6.5566
R2984 B.n700 B.n699 6.5566
R2985 B.n683 B.n573 6.5566
R2986 B.n892 B.t1 4.96776
R2987 B.n430 B.t7 4.96776
R2988 B.t3 B.n1125 4.96776
R2989 B.n1094 B.t2 4.96776
R2990 B.n274 B.n163 4.05904
R2991 B.n295 B.n294 4.05904
R2992 B.n701 B.n700 4.05904
R2993 B.n680 B.n573 4.05904
R2994 B.n1152 B.n0 2.81026
R2995 B.n1152 B.n1 2.81026
R2996 B.n838 B.t11 1.9874
R2997 B.n1060 B.t15 1.9874
R2998 VN.n8 VN.t1 216.532
R2999 VN.n44 VN.t8 216.532
R3000 VN.n9 VN.t6 183.138
R3001 VN.n5 VN.t0 183.138
R3002 VN.n26 VN.t3 183.138
R3003 VN.n34 VN.t7 183.138
R3004 VN.n45 VN.t9 183.138
R3005 VN.n41 VN.t2 183.138
R3006 VN.n62 VN.t4 183.138
R3007 VN.n70 VN.t5 183.138
R3008 VN.n69 VN.n36 161.3
R3009 VN.n68 VN.n67 161.3
R3010 VN.n66 VN.n37 161.3
R3011 VN.n65 VN.n64 161.3
R3012 VN.n63 VN.n38 161.3
R3013 VN.n61 VN.n60 161.3
R3014 VN.n59 VN.n39 161.3
R3015 VN.n58 VN.n57 161.3
R3016 VN.n56 VN.n40 161.3
R3017 VN.n55 VN.n54 161.3
R3018 VN.n53 VN.n52 161.3
R3019 VN.n51 VN.n42 161.3
R3020 VN.n50 VN.n49 161.3
R3021 VN.n48 VN.n43 161.3
R3022 VN.n47 VN.n46 161.3
R3023 VN.n33 VN.n0 161.3
R3024 VN.n32 VN.n31 161.3
R3025 VN.n30 VN.n1 161.3
R3026 VN.n29 VN.n28 161.3
R3027 VN.n27 VN.n2 161.3
R3028 VN.n25 VN.n24 161.3
R3029 VN.n23 VN.n3 161.3
R3030 VN.n22 VN.n21 161.3
R3031 VN.n20 VN.n4 161.3
R3032 VN.n19 VN.n18 161.3
R3033 VN.n17 VN.n16 161.3
R3034 VN.n15 VN.n6 161.3
R3035 VN.n14 VN.n13 161.3
R3036 VN.n12 VN.n7 161.3
R3037 VN.n11 VN.n10 161.3
R3038 VN.n35 VN.n34 93.6295
R3039 VN.n71 VN.n70 93.6295
R3040 VN.n9 VN.n8 56.5548
R3041 VN.n45 VN.n44 56.5548
R3042 VN VN.n71 55.055
R3043 VN.n32 VN.n1 47.7779
R3044 VN.n68 VN.n37 47.7779
R3045 VN.n14 VN.n7 42.9216
R3046 VN.n21 VN.n3 42.9216
R3047 VN.n50 VN.n43 42.9216
R3048 VN.n57 VN.n39 42.9216
R3049 VN.n15 VN.n14 38.0652
R3050 VN.n21 VN.n20 38.0652
R3051 VN.n51 VN.n50 38.0652
R3052 VN.n57 VN.n56 38.0652
R3053 VN.n28 VN.n1 33.2089
R3054 VN.n64 VN.n37 33.2089
R3055 VN.n10 VN.n7 24.4675
R3056 VN.n16 VN.n15 24.4675
R3057 VN.n20 VN.n19 24.4675
R3058 VN.n25 VN.n3 24.4675
R3059 VN.n28 VN.n27 24.4675
R3060 VN.n33 VN.n32 24.4675
R3061 VN.n46 VN.n43 24.4675
R3062 VN.n56 VN.n55 24.4675
R3063 VN.n52 VN.n51 24.4675
R3064 VN.n64 VN.n63 24.4675
R3065 VN.n61 VN.n39 24.4675
R3066 VN.n69 VN.n68 24.4675
R3067 VN.n34 VN.n33 17.1274
R3068 VN.n70 VN.n69 17.1274
R3069 VN.n10 VN.n9 14.6807
R3070 VN.n26 VN.n25 14.6807
R3071 VN.n46 VN.n45 14.6807
R3072 VN.n62 VN.n61 14.6807
R3073 VN.n16 VN.n5 12.234
R3074 VN.n19 VN.n5 12.234
R3075 VN.n55 VN.n41 12.234
R3076 VN.n52 VN.n41 12.234
R3077 VN.n27 VN.n26 9.7873
R3078 VN.n63 VN.n62 9.7873
R3079 VN.n47 VN.n44 9.24318
R3080 VN.n11 VN.n8 9.24318
R3081 VN.n71 VN.n36 0.278367
R3082 VN.n35 VN.n0 0.278367
R3083 VN.n67 VN.n36 0.189894
R3084 VN.n67 VN.n66 0.189894
R3085 VN.n66 VN.n65 0.189894
R3086 VN.n65 VN.n38 0.189894
R3087 VN.n60 VN.n38 0.189894
R3088 VN.n60 VN.n59 0.189894
R3089 VN.n59 VN.n58 0.189894
R3090 VN.n58 VN.n40 0.189894
R3091 VN.n54 VN.n40 0.189894
R3092 VN.n54 VN.n53 0.189894
R3093 VN.n53 VN.n42 0.189894
R3094 VN.n49 VN.n42 0.189894
R3095 VN.n49 VN.n48 0.189894
R3096 VN.n48 VN.n47 0.189894
R3097 VN.n12 VN.n11 0.189894
R3098 VN.n13 VN.n12 0.189894
R3099 VN.n13 VN.n6 0.189894
R3100 VN.n17 VN.n6 0.189894
R3101 VN.n18 VN.n17 0.189894
R3102 VN.n18 VN.n4 0.189894
R3103 VN.n22 VN.n4 0.189894
R3104 VN.n23 VN.n22 0.189894
R3105 VN.n24 VN.n23 0.189894
R3106 VN.n24 VN.n2 0.189894
R3107 VN.n29 VN.n2 0.189894
R3108 VN.n30 VN.n29 0.189894
R3109 VN.n31 VN.n30 0.189894
R3110 VN.n31 VN.n0 0.189894
R3111 VN VN.n35 0.153454
R3112 VDD2.n185 VDD2.n97 289.615
R3113 VDD2.n88 VDD2.n0 289.615
R3114 VDD2.n186 VDD2.n185 185
R3115 VDD2.n184 VDD2.n183 185
R3116 VDD2.n101 VDD2.n100 185
R3117 VDD2.n178 VDD2.n177 185
R3118 VDD2.n176 VDD2.n175 185
R3119 VDD2.n174 VDD2.n104 185
R3120 VDD2.n108 VDD2.n105 185
R3121 VDD2.n169 VDD2.n168 185
R3122 VDD2.n167 VDD2.n166 185
R3123 VDD2.n110 VDD2.n109 185
R3124 VDD2.n161 VDD2.n160 185
R3125 VDD2.n159 VDD2.n158 185
R3126 VDD2.n114 VDD2.n113 185
R3127 VDD2.n153 VDD2.n152 185
R3128 VDD2.n151 VDD2.n150 185
R3129 VDD2.n118 VDD2.n117 185
R3130 VDD2.n145 VDD2.n144 185
R3131 VDD2.n143 VDD2.n142 185
R3132 VDD2.n122 VDD2.n121 185
R3133 VDD2.n137 VDD2.n136 185
R3134 VDD2.n135 VDD2.n134 185
R3135 VDD2.n126 VDD2.n125 185
R3136 VDD2.n129 VDD2.n128 185
R3137 VDD2.n31 VDD2.n30 185
R3138 VDD2.n28 VDD2.n27 185
R3139 VDD2.n37 VDD2.n36 185
R3140 VDD2.n39 VDD2.n38 185
R3141 VDD2.n24 VDD2.n23 185
R3142 VDD2.n45 VDD2.n44 185
R3143 VDD2.n47 VDD2.n46 185
R3144 VDD2.n20 VDD2.n19 185
R3145 VDD2.n53 VDD2.n52 185
R3146 VDD2.n55 VDD2.n54 185
R3147 VDD2.n16 VDD2.n15 185
R3148 VDD2.n61 VDD2.n60 185
R3149 VDD2.n63 VDD2.n62 185
R3150 VDD2.n12 VDD2.n11 185
R3151 VDD2.n69 VDD2.n68 185
R3152 VDD2.n72 VDD2.n71 185
R3153 VDD2.n70 VDD2.n8 185
R3154 VDD2.n77 VDD2.n7 185
R3155 VDD2.n79 VDD2.n78 185
R3156 VDD2.n81 VDD2.n80 185
R3157 VDD2.n4 VDD2.n3 185
R3158 VDD2.n87 VDD2.n86 185
R3159 VDD2.n89 VDD2.n88 185
R3160 VDD2.t4 VDD2.n127 147.659
R3161 VDD2.t8 VDD2.n29 147.659
R3162 VDD2.n185 VDD2.n184 104.615
R3163 VDD2.n184 VDD2.n100 104.615
R3164 VDD2.n177 VDD2.n100 104.615
R3165 VDD2.n177 VDD2.n176 104.615
R3166 VDD2.n176 VDD2.n104 104.615
R3167 VDD2.n108 VDD2.n104 104.615
R3168 VDD2.n168 VDD2.n108 104.615
R3169 VDD2.n168 VDD2.n167 104.615
R3170 VDD2.n167 VDD2.n109 104.615
R3171 VDD2.n160 VDD2.n109 104.615
R3172 VDD2.n160 VDD2.n159 104.615
R3173 VDD2.n159 VDD2.n113 104.615
R3174 VDD2.n152 VDD2.n113 104.615
R3175 VDD2.n152 VDD2.n151 104.615
R3176 VDD2.n151 VDD2.n117 104.615
R3177 VDD2.n144 VDD2.n117 104.615
R3178 VDD2.n144 VDD2.n143 104.615
R3179 VDD2.n143 VDD2.n121 104.615
R3180 VDD2.n136 VDD2.n121 104.615
R3181 VDD2.n136 VDD2.n135 104.615
R3182 VDD2.n135 VDD2.n125 104.615
R3183 VDD2.n128 VDD2.n125 104.615
R3184 VDD2.n30 VDD2.n27 104.615
R3185 VDD2.n37 VDD2.n27 104.615
R3186 VDD2.n38 VDD2.n37 104.615
R3187 VDD2.n38 VDD2.n23 104.615
R3188 VDD2.n45 VDD2.n23 104.615
R3189 VDD2.n46 VDD2.n45 104.615
R3190 VDD2.n46 VDD2.n19 104.615
R3191 VDD2.n53 VDD2.n19 104.615
R3192 VDD2.n54 VDD2.n53 104.615
R3193 VDD2.n54 VDD2.n15 104.615
R3194 VDD2.n61 VDD2.n15 104.615
R3195 VDD2.n62 VDD2.n61 104.615
R3196 VDD2.n62 VDD2.n11 104.615
R3197 VDD2.n69 VDD2.n11 104.615
R3198 VDD2.n71 VDD2.n69 104.615
R3199 VDD2.n71 VDD2.n70 104.615
R3200 VDD2.n70 VDD2.n7 104.615
R3201 VDD2.n79 VDD2.n7 104.615
R3202 VDD2.n80 VDD2.n79 104.615
R3203 VDD2.n80 VDD2.n3 104.615
R3204 VDD2.n87 VDD2.n3 104.615
R3205 VDD2.n88 VDD2.n87 104.615
R3206 VDD2.n96 VDD2.n95 63.6756
R3207 VDD2 VDD2.n193 63.6727
R3208 VDD2.n192 VDD2.n191 62.0824
R3209 VDD2.n94 VDD2.n93 62.0822
R3210 VDD2.n94 VDD2.n92 52.42
R3211 VDD2.n128 VDD2.t4 52.3082
R3212 VDD2.n30 VDD2.t8 52.3082
R3213 VDD2.n190 VDD2.n189 50.2217
R3214 VDD2.n190 VDD2.n96 48.7002
R3215 VDD2.n129 VDD2.n127 15.6677
R3216 VDD2.n31 VDD2.n29 15.6677
R3217 VDD2.n175 VDD2.n174 13.1884
R3218 VDD2.n78 VDD2.n77 13.1884
R3219 VDD2.n178 VDD2.n103 12.8005
R3220 VDD2.n173 VDD2.n105 12.8005
R3221 VDD2.n130 VDD2.n126 12.8005
R3222 VDD2.n32 VDD2.n28 12.8005
R3223 VDD2.n76 VDD2.n8 12.8005
R3224 VDD2.n81 VDD2.n6 12.8005
R3225 VDD2.n179 VDD2.n101 12.0247
R3226 VDD2.n170 VDD2.n169 12.0247
R3227 VDD2.n134 VDD2.n133 12.0247
R3228 VDD2.n36 VDD2.n35 12.0247
R3229 VDD2.n73 VDD2.n72 12.0247
R3230 VDD2.n82 VDD2.n4 12.0247
R3231 VDD2.n183 VDD2.n182 11.249
R3232 VDD2.n166 VDD2.n107 11.249
R3233 VDD2.n137 VDD2.n124 11.249
R3234 VDD2.n39 VDD2.n26 11.249
R3235 VDD2.n68 VDD2.n10 11.249
R3236 VDD2.n86 VDD2.n85 11.249
R3237 VDD2.n186 VDD2.n99 10.4732
R3238 VDD2.n165 VDD2.n110 10.4732
R3239 VDD2.n138 VDD2.n122 10.4732
R3240 VDD2.n40 VDD2.n24 10.4732
R3241 VDD2.n67 VDD2.n12 10.4732
R3242 VDD2.n89 VDD2.n2 10.4732
R3243 VDD2.n187 VDD2.n97 9.69747
R3244 VDD2.n162 VDD2.n161 9.69747
R3245 VDD2.n142 VDD2.n141 9.69747
R3246 VDD2.n44 VDD2.n43 9.69747
R3247 VDD2.n64 VDD2.n63 9.69747
R3248 VDD2.n90 VDD2.n0 9.69747
R3249 VDD2.n189 VDD2.n188 9.45567
R3250 VDD2.n92 VDD2.n91 9.45567
R3251 VDD2.n155 VDD2.n154 9.3005
R3252 VDD2.n157 VDD2.n156 9.3005
R3253 VDD2.n112 VDD2.n111 9.3005
R3254 VDD2.n163 VDD2.n162 9.3005
R3255 VDD2.n165 VDD2.n164 9.3005
R3256 VDD2.n107 VDD2.n106 9.3005
R3257 VDD2.n171 VDD2.n170 9.3005
R3258 VDD2.n173 VDD2.n172 9.3005
R3259 VDD2.n188 VDD2.n187 9.3005
R3260 VDD2.n99 VDD2.n98 9.3005
R3261 VDD2.n182 VDD2.n181 9.3005
R3262 VDD2.n180 VDD2.n179 9.3005
R3263 VDD2.n103 VDD2.n102 9.3005
R3264 VDD2.n116 VDD2.n115 9.3005
R3265 VDD2.n149 VDD2.n148 9.3005
R3266 VDD2.n147 VDD2.n146 9.3005
R3267 VDD2.n120 VDD2.n119 9.3005
R3268 VDD2.n141 VDD2.n140 9.3005
R3269 VDD2.n139 VDD2.n138 9.3005
R3270 VDD2.n124 VDD2.n123 9.3005
R3271 VDD2.n133 VDD2.n132 9.3005
R3272 VDD2.n131 VDD2.n130 9.3005
R3273 VDD2.n91 VDD2.n90 9.3005
R3274 VDD2.n2 VDD2.n1 9.3005
R3275 VDD2.n85 VDD2.n84 9.3005
R3276 VDD2.n83 VDD2.n82 9.3005
R3277 VDD2.n6 VDD2.n5 9.3005
R3278 VDD2.n51 VDD2.n50 9.3005
R3279 VDD2.n49 VDD2.n48 9.3005
R3280 VDD2.n22 VDD2.n21 9.3005
R3281 VDD2.n43 VDD2.n42 9.3005
R3282 VDD2.n41 VDD2.n40 9.3005
R3283 VDD2.n26 VDD2.n25 9.3005
R3284 VDD2.n35 VDD2.n34 9.3005
R3285 VDD2.n33 VDD2.n32 9.3005
R3286 VDD2.n18 VDD2.n17 9.3005
R3287 VDD2.n57 VDD2.n56 9.3005
R3288 VDD2.n59 VDD2.n58 9.3005
R3289 VDD2.n14 VDD2.n13 9.3005
R3290 VDD2.n65 VDD2.n64 9.3005
R3291 VDD2.n67 VDD2.n66 9.3005
R3292 VDD2.n10 VDD2.n9 9.3005
R3293 VDD2.n74 VDD2.n73 9.3005
R3294 VDD2.n76 VDD2.n75 9.3005
R3295 VDD2.n158 VDD2.n112 8.92171
R3296 VDD2.n145 VDD2.n120 8.92171
R3297 VDD2.n47 VDD2.n22 8.92171
R3298 VDD2.n60 VDD2.n14 8.92171
R3299 VDD2.n157 VDD2.n114 8.14595
R3300 VDD2.n146 VDD2.n118 8.14595
R3301 VDD2.n48 VDD2.n20 8.14595
R3302 VDD2.n59 VDD2.n16 8.14595
R3303 VDD2.n154 VDD2.n153 7.3702
R3304 VDD2.n150 VDD2.n149 7.3702
R3305 VDD2.n52 VDD2.n51 7.3702
R3306 VDD2.n56 VDD2.n55 7.3702
R3307 VDD2.n153 VDD2.n116 6.59444
R3308 VDD2.n150 VDD2.n116 6.59444
R3309 VDD2.n52 VDD2.n18 6.59444
R3310 VDD2.n55 VDD2.n18 6.59444
R3311 VDD2.n154 VDD2.n114 5.81868
R3312 VDD2.n149 VDD2.n118 5.81868
R3313 VDD2.n51 VDD2.n20 5.81868
R3314 VDD2.n56 VDD2.n16 5.81868
R3315 VDD2.n158 VDD2.n157 5.04292
R3316 VDD2.n146 VDD2.n145 5.04292
R3317 VDD2.n48 VDD2.n47 5.04292
R3318 VDD2.n60 VDD2.n59 5.04292
R3319 VDD2.n131 VDD2.n127 4.38563
R3320 VDD2.n33 VDD2.n29 4.38563
R3321 VDD2.n189 VDD2.n97 4.26717
R3322 VDD2.n161 VDD2.n112 4.26717
R3323 VDD2.n142 VDD2.n120 4.26717
R3324 VDD2.n44 VDD2.n22 4.26717
R3325 VDD2.n63 VDD2.n14 4.26717
R3326 VDD2.n92 VDD2.n0 4.26717
R3327 VDD2.n187 VDD2.n186 3.49141
R3328 VDD2.n162 VDD2.n110 3.49141
R3329 VDD2.n141 VDD2.n122 3.49141
R3330 VDD2.n43 VDD2.n24 3.49141
R3331 VDD2.n64 VDD2.n12 3.49141
R3332 VDD2.n90 VDD2.n89 3.49141
R3333 VDD2.n183 VDD2.n99 2.71565
R3334 VDD2.n166 VDD2.n165 2.71565
R3335 VDD2.n138 VDD2.n137 2.71565
R3336 VDD2.n40 VDD2.n39 2.71565
R3337 VDD2.n68 VDD2.n67 2.71565
R3338 VDD2.n86 VDD2.n2 2.71565
R3339 VDD2.n192 VDD2.n190 2.19878
R3340 VDD2.n182 VDD2.n101 1.93989
R3341 VDD2.n169 VDD2.n107 1.93989
R3342 VDD2.n134 VDD2.n124 1.93989
R3343 VDD2.n36 VDD2.n26 1.93989
R3344 VDD2.n72 VDD2.n10 1.93989
R3345 VDD2.n85 VDD2.n4 1.93989
R3346 VDD2.n193 VDD2.t0 1.17418
R3347 VDD2.n193 VDD2.t1 1.17418
R3348 VDD2.n191 VDD2.t5 1.17418
R3349 VDD2.n191 VDD2.t7 1.17418
R3350 VDD2.n95 VDD2.t6 1.17418
R3351 VDD2.n95 VDD2.t2 1.17418
R3352 VDD2.n93 VDD2.t3 1.17418
R3353 VDD2.n93 VDD2.t9 1.17418
R3354 VDD2.n179 VDD2.n178 1.16414
R3355 VDD2.n170 VDD2.n105 1.16414
R3356 VDD2.n133 VDD2.n126 1.16414
R3357 VDD2.n35 VDD2.n28 1.16414
R3358 VDD2.n73 VDD2.n8 1.16414
R3359 VDD2.n82 VDD2.n81 1.16414
R3360 VDD2 VDD2.n192 0.608259
R3361 VDD2.n96 VDD2.n94 0.494723
R3362 VDD2.n175 VDD2.n103 0.388379
R3363 VDD2.n174 VDD2.n173 0.388379
R3364 VDD2.n130 VDD2.n129 0.388379
R3365 VDD2.n32 VDD2.n31 0.388379
R3366 VDD2.n77 VDD2.n76 0.388379
R3367 VDD2.n78 VDD2.n6 0.388379
R3368 VDD2.n188 VDD2.n98 0.155672
R3369 VDD2.n181 VDD2.n98 0.155672
R3370 VDD2.n181 VDD2.n180 0.155672
R3371 VDD2.n180 VDD2.n102 0.155672
R3372 VDD2.n172 VDD2.n102 0.155672
R3373 VDD2.n172 VDD2.n171 0.155672
R3374 VDD2.n171 VDD2.n106 0.155672
R3375 VDD2.n164 VDD2.n106 0.155672
R3376 VDD2.n164 VDD2.n163 0.155672
R3377 VDD2.n163 VDD2.n111 0.155672
R3378 VDD2.n156 VDD2.n111 0.155672
R3379 VDD2.n156 VDD2.n155 0.155672
R3380 VDD2.n155 VDD2.n115 0.155672
R3381 VDD2.n148 VDD2.n115 0.155672
R3382 VDD2.n148 VDD2.n147 0.155672
R3383 VDD2.n147 VDD2.n119 0.155672
R3384 VDD2.n140 VDD2.n119 0.155672
R3385 VDD2.n140 VDD2.n139 0.155672
R3386 VDD2.n139 VDD2.n123 0.155672
R3387 VDD2.n132 VDD2.n123 0.155672
R3388 VDD2.n132 VDD2.n131 0.155672
R3389 VDD2.n34 VDD2.n33 0.155672
R3390 VDD2.n34 VDD2.n25 0.155672
R3391 VDD2.n41 VDD2.n25 0.155672
R3392 VDD2.n42 VDD2.n41 0.155672
R3393 VDD2.n42 VDD2.n21 0.155672
R3394 VDD2.n49 VDD2.n21 0.155672
R3395 VDD2.n50 VDD2.n49 0.155672
R3396 VDD2.n50 VDD2.n17 0.155672
R3397 VDD2.n57 VDD2.n17 0.155672
R3398 VDD2.n58 VDD2.n57 0.155672
R3399 VDD2.n58 VDD2.n13 0.155672
R3400 VDD2.n65 VDD2.n13 0.155672
R3401 VDD2.n66 VDD2.n65 0.155672
R3402 VDD2.n66 VDD2.n9 0.155672
R3403 VDD2.n74 VDD2.n9 0.155672
R3404 VDD2.n75 VDD2.n74 0.155672
R3405 VDD2.n75 VDD2.n5 0.155672
R3406 VDD2.n83 VDD2.n5 0.155672
R3407 VDD2.n84 VDD2.n83 0.155672
R3408 VDD2.n84 VDD2.n1 0.155672
R3409 VDD2.n91 VDD2.n1 0.155672
C0 VDD1 VDD2 1.9259f
C1 VTAIL VDD1 12.8137f
C2 VP VDD2 0.535284f
C3 VP VTAIL 14.585599f
C4 VN VDD2 14.298599f
C5 VP VDD1 14.676901f
C6 VN VTAIL 14.571199f
C7 VN VDD1 0.152219f
C8 VP VN 8.74014f
C9 VTAIL VDD2 12.8604f
C10 VDD2 B 7.587809f
C11 VDD1 B 7.587282f
C12 VTAIL B 9.820148f
C13 VN B 16.77873f
C14 VP B 15.171201f
C15 VDD2.n0 B 0.030772f
C16 VDD2.n1 B 0.021999f
C17 VDD2.n2 B 0.011821f
C18 VDD2.n3 B 0.027941f
C19 VDD2.n4 B 0.012516f
C20 VDD2.n5 B 0.021999f
C21 VDD2.n6 B 0.011821f
C22 VDD2.n7 B 0.027941f
C23 VDD2.n8 B 0.012516f
C24 VDD2.n9 B 0.021999f
C25 VDD2.n10 B 0.011821f
C26 VDD2.n11 B 0.027941f
C27 VDD2.n12 B 0.012516f
C28 VDD2.n13 B 0.021999f
C29 VDD2.n14 B 0.011821f
C30 VDD2.n15 B 0.027941f
C31 VDD2.n16 B 0.012516f
C32 VDD2.n17 B 0.021999f
C33 VDD2.n18 B 0.011821f
C34 VDD2.n19 B 0.027941f
C35 VDD2.n20 B 0.012516f
C36 VDD2.n21 B 0.021999f
C37 VDD2.n22 B 0.011821f
C38 VDD2.n23 B 0.027941f
C39 VDD2.n24 B 0.012516f
C40 VDD2.n25 B 0.021999f
C41 VDD2.n26 B 0.011821f
C42 VDD2.n27 B 0.027941f
C43 VDD2.n28 B 0.012516f
C44 VDD2.n29 B 0.153793f
C45 VDD2.t8 B 0.046212f
C46 VDD2.n30 B 0.020955f
C47 VDD2.n31 B 0.016505f
C48 VDD2.n32 B 0.011821f
C49 VDD2.n33 B 1.61979f
C50 VDD2.n34 B 0.021999f
C51 VDD2.n35 B 0.011821f
C52 VDD2.n36 B 0.012516f
C53 VDD2.n37 B 0.027941f
C54 VDD2.n38 B 0.027941f
C55 VDD2.n39 B 0.012516f
C56 VDD2.n40 B 0.011821f
C57 VDD2.n41 B 0.021999f
C58 VDD2.n42 B 0.021999f
C59 VDD2.n43 B 0.011821f
C60 VDD2.n44 B 0.012516f
C61 VDD2.n45 B 0.027941f
C62 VDD2.n46 B 0.027941f
C63 VDD2.n47 B 0.012516f
C64 VDD2.n48 B 0.011821f
C65 VDD2.n49 B 0.021999f
C66 VDD2.n50 B 0.021999f
C67 VDD2.n51 B 0.011821f
C68 VDD2.n52 B 0.012516f
C69 VDD2.n53 B 0.027941f
C70 VDD2.n54 B 0.027941f
C71 VDD2.n55 B 0.012516f
C72 VDD2.n56 B 0.011821f
C73 VDD2.n57 B 0.021999f
C74 VDD2.n58 B 0.021999f
C75 VDD2.n59 B 0.011821f
C76 VDD2.n60 B 0.012516f
C77 VDD2.n61 B 0.027941f
C78 VDD2.n62 B 0.027941f
C79 VDD2.n63 B 0.012516f
C80 VDD2.n64 B 0.011821f
C81 VDD2.n65 B 0.021999f
C82 VDD2.n66 B 0.021999f
C83 VDD2.n67 B 0.011821f
C84 VDD2.n68 B 0.012516f
C85 VDD2.n69 B 0.027941f
C86 VDD2.n70 B 0.027941f
C87 VDD2.n71 B 0.027941f
C88 VDD2.n72 B 0.012516f
C89 VDD2.n73 B 0.011821f
C90 VDD2.n74 B 0.021999f
C91 VDD2.n75 B 0.021999f
C92 VDD2.n76 B 0.011821f
C93 VDD2.n77 B 0.012169f
C94 VDD2.n78 B 0.012169f
C95 VDD2.n79 B 0.027941f
C96 VDD2.n80 B 0.027941f
C97 VDD2.n81 B 0.012516f
C98 VDD2.n82 B 0.011821f
C99 VDD2.n83 B 0.021999f
C100 VDD2.n84 B 0.021999f
C101 VDD2.n85 B 0.011821f
C102 VDD2.n86 B 0.012516f
C103 VDD2.n87 B 0.027941f
C104 VDD2.n88 B 0.060224f
C105 VDD2.n89 B 0.012516f
C106 VDD2.n90 B 0.011821f
C107 VDD2.n91 B 0.052952f
C108 VDD2.n92 B 0.057269f
C109 VDD2.t3 B 0.293266f
C110 VDD2.t9 B 0.293266f
C111 VDD2.n93 B 2.66588f
C112 VDD2.n94 B 0.563482f
C113 VDD2.t6 B 0.293266f
C114 VDD2.t2 B 0.293266f
C115 VDD2.n95 B 2.67735f
C116 VDD2.n96 B 2.64823f
C117 VDD2.n97 B 0.030772f
C118 VDD2.n98 B 0.021999f
C119 VDD2.n99 B 0.011821f
C120 VDD2.n100 B 0.027941f
C121 VDD2.n101 B 0.012516f
C122 VDD2.n102 B 0.021999f
C123 VDD2.n103 B 0.011821f
C124 VDD2.n104 B 0.027941f
C125 VDD2.n105 B 0.012516f
C126 VDD2.n106 B 0.021999f
C127 VDD2.n107 B 0.011821f
C128 VDD2.n108 B 0.027941f
C129 VDD2.n109 B 0.027941f
C130 VDD2.n110 B 0.012516f
C131 VDD2.n111 B 0.021999f
C132 VDD2.n112 B 0.011821f
C133 VDD2.n113 B 0.027941f
C134 VDD2.n114 B 0.012516f
C135 VDD2.n115 B 0.021999f
C136 VDD2.n116 B 0.011821f
C137 VDD2.n117 B 0.027941f
C138 VDD2.n118 B 0.012516f
C139 VDD2.n119 B 0.021999f
C140 VDD2.n120 B 0.011821f
C141 VDD2.n121 B 0.027941f
C142 VDD2.n122 B 0.012516f
C143 VDD2.n123 B 0.021999f
C144 VDD2.n124 B 0.011821f
C145 VDD2.n125 B 0.027941f
C146 VDD2.n126 B 0.012516f
C147 VDD2.n127 B 0.153793f
C148 VDD2.t4 B 0.046212f
C149 VDD2.n128 B 0.020955f
C150 VDD2.n129 B 0.016505f
C151 VDD2.n130 B 0.011821f
C152 VDD2.n131 B 1.61979f
C153 VDD2.n132 B 0.021999f
C154 VDD2.n133 B 0.011821f
C155 VDD2.n134 B 0.012516f
C156 VDD2.n135 B 0.027941f
C157 VDD2.n136 B 0.027941f
C158 VDD2.n137 B 0.012516f
C159 VDD2.n138 B 0.011821f
C160 VDD2.n139 B 0.021999f
C161 VDD2.n140 B 0.021999f
C162 VDD2.n141 B 0.011821f
C163 VDD2.n142 B 0.012516f
C164 VDD2.n143 B 0.027941f
C165 VDD2.n144 B 0.027941f
C166 VDD2.n145 B 0.012516f
C167 VDD2.n146 B 0.011821f
C168 VDD2.n147 B 0.021999f
C169 VDD2.n148 B 0.021999f
C170 VDD2.n149 B 0.011821f
C171 VDD2.n150 B 0.012516f
C172 VDD2.n151 B 0.027941f
C173 VDD2.n152 B 0.027941f
C174 VDD2.n153 B 0.012516f
C175 VDD2.n154 B 0.011821f
C176 VDD2.n155 B 0.021999f
C177 VDD2.n156 B 0.021999f
C178 VDD2.n157 B 0.011821f
C179 VDD2.n158 B 0.012516f
C180 VDD2.n159 B 0.027941f
C181 VDD2.n160 B 0.027941f
C182 VDD2.n161 B 0.012516f
C183 VDD2.n162 B 0.011821f
C184 VDD2.n163 B 0.021999f
C185 VDD2.n164 B 0.021999f
C186 VDD2.n165 B 0.011821f
C187 VDD2.n166 B 0.012516f
C188 VDD2.n167 B 0.027941f
C189 VDD2.n168 B 0.027941f
C190 VDD2.n169 B 0.012516f
C191 VDD2.n170 B 0.011821f
C192 VDD2.n171 B 0.021999f
C193 VDD2.n172 B 0.021999f
C194 VDD2.n173 B 0.011821f
C195 VDD2.n174 B 0.012169f
C196 VDD2.n175 B 0.012169f
C197 VDD2.n176 B 0.027941f
C198 VDD2.n177 B 0.027941f
C199 VDD2.n178 B 0.012516f
C200 VDD2.n179 B 0.011821f
C201 VDD2.n180 B 0.021999f
C202 VDD2.n181 B 0.021999f
C203 VDD2.n182 B 0.011821f
C204 VDD2.n183 B 0.012516f
C205 VDD2.n184 B 0.027941f
C206 VDD2.n185 B 0.060224f
C207 VDD2.n186 B 0.012516f
C208 VDD2.n187 B 0.011821f
C209 VDD2.n188 B 0.052952f
C210 VDD2.n189 B 0.048908f
C211 VDD2.n190 B 2.74241f
C212 VDD2.t5 B 0.293266f
C213 VDD2.t7 B 0.293266f
C214 VDD2.n191 B 2.66588f
C215 VDD2.n192 B 0.379464f
C216 VDD2.t0 B 0.293266f
C217 VDD2.t1 B 0.293266f
C218 VDD2.n193 B 2.67732f
C219 VN.n0 B 0.030282f
C220 VN.t7 B 2.36305f
C221 VN.n1 B 0.020284f
C222 VN.n2 B 0.022968f
C223 VN.t3 B 2.36305f
C224 VN.n3 B 0.044988f
C225 VN.n4 B 0.022968f
C226 VN.t0 B 2.36305f
C227 VN.n5 B 0.824694f
C228 VN.n6 B 0.022968f
C229 VN.n7 B 0.044988f
C230 VN.t1 B 2.50976f
C231 VN.n8 B 0.875179f
C232 VN.t6 B 2.36305f
C233 VN.n9 B 0.886215f
C234 VN.n10 B 0.034354f
C235 VN.n11 B 0.196014f
C236 VN.n12 B 0.022968f
C237 VN.n13 B 0.022968f
C238 VN.n14 B 0.018754f
C239 VN.n15 B 0.046129f
C240 VN.n16 B 0.03224f
C241 VN.n17 B 0.022968f
C242 VN.n18 B 0.022968f
C243 VN.n19 B 0.03224f
C244 VN.n20 B 0.046129f
C245 VN.n21 B 0.018754f
C246 VN.n22 B 0.022968f
C247 VN.n23 B 0.022968f
C248 VN.n24 B 0.022968f
C249 VN.n25 B 0.034354f
C250 VN.n26 B 0.824694f
C251 VN.n27 B 0.030127f
C252 VN.n28 B 0.046368f
C253 VN.n29 B 0.022968f
C254 VN.n30 B 0.022968f
C255 VN.n31 B 0.022968f
C256 VN.n32 B 0.04322f
C257 VN.n33 B 0.036467f
C258 VN.n34 B 0.898973f
C259 VN.n35 B 0.030591f
C260 VN.n36 B 0.030282f
C261 VN.t5 B 2.36305f
C262 VN.n37 B 0.020284f
C263 VN.n38 B 0.022968f
C264 VN.t4 B 2.36305f
C265 VN.n39 B 0.044988f
C266 VN.n40 B 0.022968f
C267 VN.t2 B 2.36305f
C268 VN.n41 B 0.824694f
C269 VN.n42 B 0.022968f
C270 VN.n43 B 0.044988f
C271 VN.t8 B 2.50976f
C272 VN.n44 B 0.875179f
C273 VN.t9 B 2.36305f
C274 VN.n45 B 0.886215f
C275 VN.n46 B 0.034354f
C276 VN.n47 B 0.196014f
C277 VN.n48 B 0.022968f
C278 VN.n49 B 0.022968f
C279 VN.n50 B 0.018754f
C280 VN.n51 B 0.046129f
C281 VN.n52 B 0.03224f
C282 VN.n53 B 0.022968f
C283 VN.n54 B 0.022968f
C284 VN.n55 B 0.03224f
C285 VN.n56 B 0.046129f
C286 VN.n57 B 0.018754f
C287 VN.n58 B 0.022968f
C288 VN.n59 B 0.022968f
C289 VN.n60 B 0.022968f
C290 VN.n61 B 0.034354f
C291 VN.n62 B 0.824694f
C292 VN.n63 B 0.030127f
C293 VN.n64 B 0.046368f
C294 VN.n65 B 0.022968f
C295 VN.n66 B 0.022968f
C296 VN.n67 B 0.022968f
C297 VN.n68 B 0.04322f
C298 VN.n69 B 0.036467f
C299 VN.n70 B 0.898973f
C300 VN.n71 B 1.4625f
C301 VDD1.n0 B 0.031019f
C302 VDD1.n1 B 0.022175f
C303 VDD1.n2 B 0.011916f
C304 VDD1.n3 B 0.028165f
C305 VDD1.n4 B 0.012617f
C306 VDD1.n5 B 0.022175f
C307 VDD1.n6 B 0.011916f
C308 VDD1.n7 B 0.028165f
C309 VDD1.n8 B 0.012617f
C310 VDD1.n9 B 0.022175f
C311 VDD1.n10 B 0.011916f
C312 VDD1.n11 B 0.028165f
C313 VDD1.n12 B 0.028165f
C314 VDD1.n13 B 0.012617f
C315 VDD1.n14 B 0.022175f
C316 VDD1.n15 B 0.011916f
C317 VDD1.n16 B 0.028165f
C318 VDD1.n17 B 0.012617f
C319 VDD1.n18 B 0.022175f
C320 VDD1.n19 B 0.011916f
C321 VDD1.n20 B 0.028165f
C322 VDD1.n21 B 0.012617f
C323 VDD1.n22 B 0.022175f
C324 VDD1.n23 B 0.011916f
C325 VDD1.n24 B 0.028165f
C326 VDD1.n25 B 0.012617f
C327 VDD1.n26 B 0.022175f
C328 VDD1.n27 B 0.011916f
C329 VDD1.n28 B 0.028165f
C330 VDD1.n29 B 0.012617f
C331 VDD1.n30 B 0.155026f
C332 VDD1.t9 B 0.046582f
C333 VDD1.n31 B 0.021124f
C334 VDD1.n32 B 0.016638f
C335 VDD1.n33 B 0.011916f
C336 VDD1.n34 B 1.63277f
C337 VDD1.n35 B 0.022175f
C338 VDD1.n36 B 0.011916f
C339 VDD1.n37 B 0.012617f
C340 VDD1.n38 B 0.028165f
C341 VDD1.n39 B 0.028165f
C342 VDD1.n40 B 0.012617f
C343 VDD1.n41 B 0.011916f
C344 VDD1.n42 B 0.022175f
C345 VDD1.n43 B 0.022175f
C346 VDD1.n44 B 0.011916f
C347 VDD1.n45 B 0.012617f
C348 VDD1.n46 B 0.028165f
C349 VDD1.n47 B 0.028165f
C350 VDD1.n48 B 0.012617f
C351 VDD1.n49 B 0.011916f
C352 VDD1.n50 B 0.022175f
C353 VDD1.n51 B 0.022175f
C354 VDD1.n52 B 0.011916f
C355 VDD1.n53 B 0.012617f
C356 VDD1.n54 B 0.028165f
C357 VDD1.n55 B 0.028165f
C358 VDD1.n56 B 0.012617f
C359 VDD1.n57 B 0.011916f
C360 VDD1.n58 B 0.022175f
C361 VDD1.n59 B 0.022175f
C362 VDD1.n60 B 0.011916f
C363 VDD1.n61 B 0.012617f
C364 VDD1.n62 B 0.028165f
C365 VDD1.n63 B 0.028165f
C366 VDD1.n64 B 0.012617f
C367 VDD1.n65 B 0.011916f
C368 VDD1.n66 B 0.022175f
C369 VDD1.n67 B 0.022175f
C370 VDD1.n68 B 0.011916f
C371 VDD1.n69 B 0.012617f
C372 VDD1.n70 B 0.028165f
C373 VDD1.n71 B 0.028165f
C374 VDD1.n72 B 0.012617f
C375 VDD1.n73 B 0.011916f
C376 VDD1.n74 B 0.022175f
C377 VDD1.n75 B 0.022175f
C378 VDD1.n76 B 0.011916f
C379 VDD1.n77 B 0.012266f
C380 VDD1.n78 B 0.012266f
C381 VDD1.n79 B 0.028165f
C382 VDD1.n80 B 0.028165f
C383 VDD1.n81 B 0.012617f
C384 VDD1.n82 B 0.011916f
C385 VDD1.n83 B 0.022175f
C386 VDD1.n84 B 0.022175f
C387 VDD1.n85 B 0.011916f
C388 VDD1.n86 B 0.012617f
C389 VDD1.n87 B 0.028165f
C390 VDD1.n88 B 0.060707f
C391 VDD1.n89 B 0.012617f
C392 VDD1.n90 B 0.011916f
C393 VDD1.n91 B 0.053377f
C394 VDD1.n92 B 0.057729f
C395 VDD1.t7 B 0.295617f
C396 VDD1.t3 B 0.295617f
C397 VDD1.n93 B 2.68726f
C398 VDD1.n94 B 0.575064f
C399 VDD1.n95 B 0.031019f
C400 VDD1.n96 B 0.022175f
C401 VDD1.n97 B 0.011916f
C402 VDD1.n98 B 0.028165f
C403 VDD1.n99 B 0.012617f
C404 VDD1.n100 B 0.022175f
C405 VDD1.n101 B 0.011916f
C406 VDD1.n102 B 0.028165f
C407 VDD1.n103 B 0.012617f
C408 VDD1.n104 B 0.022175f
C409 VDD1.n105 B 0.011916f
C410 VDD1.n106 B 0.028165f
C411 VDD1.n107 B 0.012617f
C412 VDD1.n108 B 0.022175f
C413 VDD1.n109 B 0.011916f
C414 VDD1.n110 B 0.028165f
C415 VDD1.n111 B 0.012617f
C416 VDD1.n112 B 0.022175f
C417 VDD1.n113 B 0.011916f
C418 VDD1.n114 B 0.028165f
C419 VDD1.n115 B 0.012617f
C420 VDD1.n116 B 0.022175f
C421 VDD1.n117 B 0.011916f
C422 VDD1.n118 B 0.028165f
C423 VDD1.n119 B 0.012617f
C424 VDD1.n120 B 0.022175f
C425 VDD1.n121 B 0.011916f
C426 VDD1.n122 B 0.028165f
C427 VDD1.n123 B 0.012617f
C428 VDD1.n124 B 0.155026f
C429 VDD1.t6 B 0.046582f
C430 VDD1.n125 B 0.021124f
C431 VDD1.n126 B 0.016638f
C432 VDD1.n127 B 0.011916f
C433 VDD1.n128 B 1.63277f
C434 VDD1.n129 B 0.022175f
C435 VDD1.n130 B 0.011916f
C436 VDD1.n131 B 0.012617f
C437 VDD1.n132 B 0.028165f
C438 VDD1.n133 B 0.028165f
C439 VDD1.n134 B 0.012617f
C440 VDD1.n135 B 0.011916f
C441 VDD1.n136 B 0.022175f
C442 VDD1.n137 B 0.022175f
C443 VDD1.n138 B 0.011916f
C444 VDD1.n139 B 0.012617f
C445 VDD1.n140 B 0.028165f
C446 VDD1.n141 B 0.028165f
C447 VDD1.n142 B 0.012617f
C448 VDD1.n143 B 0.011916f
C449 VDD1.n144 B 0.022175f
C450 VDD1.n145 B 0.022175f
C451 VDD1.n146 B 0.011916f
C452 VDD1.n147 B 0.012617f
C453 VDD1.n148 B 0.028165f
C454 VDD1.n149 B 0.028165f
C455 VDD1.n150 B 0.012617f
C456 VDD1.n151 B 0.011916f
C457 VDD1.n152 B 0.022175f
C458 VDD1.n153 B 0.022175f
C459 VDD1.n154 B 0.011916f
C460 VDD1.n155 B 0.012617f
C461 VDD1.n156 B 0.028165f
C462 VDD1.n157 B 0.028165f
C463 VDD1.n158 B 0.012617f
C464 VDD1.n159 B 0.011916f
C465 VDD1.n160 B 0.022175f
C466 VDD1.n161 B 0.022175f
C467 VDD1.n162 B 0.011916f
C468 VDD1.n163 B 0.012617f
C469 VDD1.n164 B 0.028165f
C470 VDD1.n165 B 0.028165f
C471 VDD1.n166 B 0.028165f
C472 VDD1.n167 B 0.012617f
C473 VDD1.n168 B 0.011916f
C474 VDD1.n169 B 0.022175f
C475 VDD1.n170 B 0.022175f
C476 VDD1.n171 B 0.011916f
C477 VDD1.n172 B 0.012266f
C478 VDD1.n173 B 0.012266f
C479 VDD1.n174 B 0.028165f
C480 VDD1.n175 B 0.028165f
C481 VDD1.n176 B 0.012617f
C482 VDD1.n177 B 0.011916f
C483 VDD1.n178 B 0.022175f
C484 VDD1.n179 B 0.022175f
C485 VDD1.n180 B 0.011916f
C486 VDD1.n181 B 0.012617f
C487 VDD1.n182 B 0.028165f
C488 VDD1.n183 B 0.060707f
C489 VDD1.n184 B 0.012617f
C490 VDD1.n185 B 0.011916f
C491 VDD1.n186 B 0.053377f
C492 VDD1.n187 B 0.057729f
C493 VDD1.t8 B 0.295617f
C494 VDD1.t1 B 0.295617f
C495 VDD1.n188 B 2.68725f
C496 VDD1.n189 B 0.568f
C497 VDD1.t2 B 0.295617f
C498 VDD1.t5 B 0.295617f
C499 VDD1.n190 B 2.69882f
C500 VDD1.n191 B 2.77386f
C501 VDD1.t4 B 0.295617f
C502 VDD1.t0 B 0.295617f
C503 VDD1.n192 B 2.68725f
C504 VDD1.n193 B 3.00258f
C505 VTAIL.t8 B 0.316425f
C506 VTAIL.t3 B 0.316425f
C507 VTAIL.n0 B 2.80649f
C508 VTAIL.n1 B 0.483023f
C509 VTAIL.n2 B 0.033202f
C510 VTAIL.n3 B 0.023736f
C511 VTAIL.n4 B 0.012755f
C512 VTAIL.n5 B 0.030147f
C513 VTAIL.n6 B 0.013505f
C514 VTAIL.n7 B 0.023736f
C515 VTAIL.n8 B 0.012755f
C516 VTAIL.n9 B 0.030147f
C517 VTAIL.n10 B 0.013505f
C518 VTAIL.n11 B 0.023736f
C519 VTAIL.n12 B 0.012755f
C520 VTAIL.n13 B 0.030147f
C521 VTAIL.n14 B 0.013505f
C522 VTAIL.n15 B 0.023736f
C523 VTAIL.n16 B 0.012755f
C524 VTAIL.n17 B 0.030147f
C525 VTAIL.n18 B 0.013505f
C526 VTAIL.n19 B 0.023736f
C527 VTAIL.n20 B 0.012755f
C528 VTAIL.n21 B 0.030147f
C529 VTAIL.n22 B 0.013505f
C530 VTAIL.n23 B 0.023736f
C531 VTAIL.n24 B 0.012755f
C532 VTAIL.n25 B 0.030147f
C533 VTAIL.n26 B 0.013505f
C534 VTAIL.n27 B 0.023736f
C535 VTAIL.n28 B 0.012755f
C536 VTAIL.n29 B 0.030147f
C537 VTAIL.n30 B 0.013505f
C538 VTAIL.n31 B 0.165938f
C539 VTAIL.t15 B 0.049861f
C540 VTAIL.n32 B 0.02261f
C541 VTAIL.n33 B 0.017809f
C542 VTAIL.n34 B 0.012755f
C543 VTAIL.n35 B 1.7477f
C544 VTAIL.n36 B 0.023736f
C545 VTAIL.n37 B 0.012755f
C546 VTAIL.n38 B 0.013505f
C547 VTAIL.n39 B 0.030147f
C548 VTAIL.n40 B 0.030147f
C549 VTAIL.n41 B 0.013505f
C550 VTAIL.n42 B 0.012755f
C551 VTAIL.n43 B 0.023736f
C552 VTAIL.n44 B 0.023736f
C553 VTAIL.n45 B 0.012755f
C554 VTAIL.n46 B 0.013505f
C555 VTAIL.n47 B 0.030147f
C556 VTAIL.n48 B 0.030147f
C557 VTAIL.n49 B 0.013505f
C558 VTAIL.n50 B 0.012755f
C559 VTAIL.n51 B 0.023736f
C560 VTAIL.n52 B 0.023736f
C561 VTAIL.n53 B 0.012755f
C562 VTAIL.n54 B 0.013505f
C563 VTAIL.n55 B 0.030147f
C564 VTAIL.n56 B 0.030147f
C565 VTAIL.n57 B 0.013505f
C566 VTAIL.n58 B 0.012755f
C567 VTAIL.n59 B 0.023736f
C568 VTAIL.n60 B 0.023736f
C569 VTAIL.n61 B 0.012755f
C570 VTAIL.n62 B 0.013505f
C571 VTAIL.n63 B 0.030147f
C572 VTAIL.n64 B 0.030147f
C573 VTAIL.n65 B 0.013505f
C574 VTAIL.n66 B 0.012755f
C575 VTAIL.n67 B 0.023736f
C576 VTAIL.n68 B 0.023736f
C577 VTAIL.n69 B 0.012755f
C578 VTAIL.n70 B 0.013505f
C579 VTAIL.n71 B 0.030147f
C580 VTAIL.n72 B 0.030147f
C581 VTAIL.n73 B 0.030147f
C582 VTAIL.n74 B 0.013505f
C583 VTAIL.n75 B 0.012755f
C584 VTAIL.n76 B 0.023736f
C585 VTAIL.n77 B 0.023736f
C586 VTAIL.n78 B 0.012755f
C587 VTAIL.n79 B 0.01313f
C588 VTAIL.n80 B 0.01313f
C589 VTAIL.n81 B 0.030147f
C590 VTAIL.n82 B 0.030147f
C591 VTAIL.n83 B 0.013505f
C592 VTAIL.n84 B 0.012755f
C593 VTAIL.n85 B 0.023736f
C594 VTAIL.n86 B 0.023736f
C595 VTAIL.n87 B 0.012755f
C596 VTAIL.n88 B 0.013505f
C597 VTAIL.n89 B 0.030147f
C598 VTAIL.n90 B 0.06498f
C599 VTAIL.n91 B 0.013505f
C600 VTAIL.n92 B 0.012755f
C601 VTAIL.n93 B 0.057134f
C602 VTAIL.n94 B 0.036398f
C603 VTAIL.n95 B 0.30968f
C604 VTAIL.t9 B 0.316425f
C605 VTAIL.t12 B 0.316425f
C606 VTAIL.n96 B 2.80649f
C607 VTAIL.n97 B 0.568735f
C608 VTAIL.t16 B 0.316425f
C609 VTAIL.t17 B 0.316425f
C610 VTAIL.n98 B 2.80649f
C611 VTAIL.n99 B 2.17157f
C612 VTAIL.t4 B 0.316425f
C613 VTAIL.t1 B 0.316425f
C614 VTAIL.n100 B 2.8065f
C615 VTAIL.n101 B 2.17156f
C616 VTAIL.t6 B 0.316425f
C617 VTAIL.t7 B 0.316425f
C618 VTAIL.n102 B 2.8065f
C619 VTAIL.n103 B 0.568722f
C620 VTAIL.n104 B 0.033202f
C621 VTAIL.n105 B 0.023736f
C622 VTAIL.n106 B 0.012755f
C623 VTAIL.n107 B 0.030147f
C624 VTAIL.n108 B 0.013505f
C625 VTAIL.n109 B 0.023736f
C626 VTAIL.n110 B 0.012755f
C627 VTAIL.n111 B 0.030147f
C628 VTAIL.n112 B 0.013505f
C629 VTAIL.n113 B 0.023736f
C630 VTAIL.n114 B 0.012755f
C631 VTAIL.n115 B 0.030147f
C632 VTAIL.n116 B 0.030147f
C633 VTAIL.n117 B 0.013505f
C634 VTAIL.n118 B 0.023736f
C635 VTAIL.n119 B 0.012755f
C636 VTAIL.n120 B 0.030147f
C637 VTAIL.n121 B 0.013505f
C638 VTAIL.n122 B 0.023736f
C639 VTAIL.n123 B 0.012755f
C640 VTAIL.n124 B 0.030147f
C641 VTAIL.n125 B 0.013505f
C642 VTAIL.n126 B 0.023736f
C643 VTAIL.n127 B 0.012755f
C644 VTAIL.n128 B 0.030147f
C645 VTAIL.n129 B 0.013505f
C646 VTAIL.n130 B 0.023736f
C647 VTAIL.n131 B 0.012755f
C648 VTAIL.n132 B 0.030147f
C649 VTAIL.n133 B 0.013505f
C650 VTAIL.n134 B 0.165938f
C651 VTAIL.t19 B 0.049861f
C652 VTAIL.n135 B 0.02261f
C653 VTAIL.n136 B 0.017809f
C654 VTAIL.n137 B 0.012755f
C655 VTAIL.n138 B 1.7477f
C656 VTAIL.n139 B 0.023736f
C657 VTAIL.n140 B 0.012755f
C658 VTAIL.n141 B 0.013505f
C659 VTAIL.n142 B 0.030147f
C660 VTAIL.n143 B 0.030147f
C661 VTAIL.n144 B 0.013505f
C662 VTAIL.n145 B 0.012755f
C663 VTAIL.n146 B 0.023736f
C664 VTAIL.n147 B 0.023736f
C665 VTAIL.n148 B 0.012755f
C666 VTAIL.n149 B 0.013505f
C667 VTAIL.n150 B 0.030147f
C668 VTAIL.n151 B 0.030147f
C669 VTAIL.n152 B 0.013505f
C670 VTAIL.n153 B 0.012755f
C671 VTAIL.n154 B 0.023736f
C672 VTAIL.n155 B 0.023736f
C673 VTAIL.n156 B 0.012755f
C674 VTAIL.n157 B 0.013505f
C675 VTAIL.n158 B 0.030147f
C676 VTAIL.n159 B 0.030147f
C677 VTAIL.n160 B 0.013505f
C678 VTAIL.n161 B 0.012755f
C679 VTAIL.n162 B 0.023736f
C680 VTAIL.n163 B 0.023736f
C681 VTAIL.n164 B 0.012755f
C682 VTAIL.n165 B 0.013505f
C683 VTAIL.n166 B 0.030147f
C684 VTAIL.n167 B 0.030147f
C685 VTAIL.n168 B 0.013505f
C686 VTAIL.n169 B 0.012755f
C687 VTAIL.n170 B 0.023736f
C688 VTAIL.n171 B 0.023736f
C689 VTAIL.n172 B 0.012755f
C690 VTAIL.n173 B 0.013505f
C691 VTAIL.n174 B 0.030147f
C692 VTAIL.n175 B 0.030147f
C693 VTAIL.n176 B 0.013505f
C694 VTAIL.n177 B 0.012755f
C695 VTAIL.n178 B 0.023736f
C696 VTAIL.n179 B 0.023736f
C697 VTAIL.n180 B 0.012755f
C698 VTAIL.n181 B 0.01313f
C699 VTAIL.n182 B 0.01313f
C700 VTAIL.n183 B 0.030147f
C701 VTAIL.n184 B 0.030147f
C702 VTAIL.n185 B 0.013505f
C703 VTAIL.n186 B 0.012755f
C704 VTAIL.n187 B 0.023736f
C705 VTAIL.n188 B 0.023736f
C706 VTAIL.n189 B 0.012755f
C707 VTAIL.n190 B 0.013505f
C708 VTAIL.n191 B 0.030147f
C709 VTAIL.n192 B 0.06498f
C710 VTAIL.n193 B 0.013505f
C711 VTAIL.n194 B 0.012755f
C712 VTAIL.n195 B 0.057134f
C713 VTAIL.n196 B 0.036398f
C714 VTAIL.n197 B 0.30968f
C715 VTAIL.t10 B 0.316425f
C716 VTAIL.t18 B 0.316425f
C717 VTAIL.n198 B 2.8065f
C718 VTAIL.n199 B 0.520591f
C719 VTAIL.t11 B 0.316425f
C720 VTAIL.t14 B 0.316425f
C721 VTAIL.n200 B 2.8065f
C722 VTAIL.n201 B 0.568722f
C723 VTAIL.n202 B 0.033202f
C724 VTAIL.n203 B 0.023736f
C725 VTAIL.n204 B 0.012755f
C726 VTAIL.n205 B 0.030147f
C727 VTAIL.n206 B 0.013505f
C728 VTAIL.n207 B 0.023736f
C729 VTAIL.n208 B 0.012755f
C730 VTAIL.n209 B 0.030147f
C731 VTAIL.n210 B 0.013505f
C732 VTAIL.n211 B 0.023736f
C733 VTAIL.n212 B 0.012755f
C734 VTAIL.n213 B 0.030147f
C735 VTAIL.n214 B 0.030147f
C736 VTAIL.n215 B 0.013505f
C737 VTAIL.n216 B 0.023736f
C738 VTAIL.n217 B 0.012755f
C739 VTAIL.n218 B 0.030147f
C740 VTAIL.n219 B 0.013505f
C741 VTAIL.n220 B 0.023736f
C742 VTAIL.n221 B 0.012755f
C743 VTAIL.n222 B 0.030147f
C744 VTAIL.n223 B 0.013505f
C745 VTAIL.n224 B 0.023736f
C746 VTAIL.n225 B 0.012755f
C747 VTAIL.n226 B 0.030147f
C748 VTAIL.n227 B 0.013505f
C749 VTAIL.n228 B 0.023736f
C750 VTAIL.n229 B 0.012755f
C751 VTAIL.n230 B 0.030147f
C752 VTAIL.n231 B 0.013505f
C753 VTAIL.n232 B 0.165938f
C754 VTAIL.t13 B 0.049861f
C755 VTAIL.n233 B 0.02261f
C756 VTAIL.n234 B 0.017809f
C757 VTAIL.n235 B 0.012755f
C758 VTAIL.n236 B 1.7477f
C759 VTAIL.n237 B 0.023736f
C760 VTAIL.n238 B 0.012755f
C761 VTAIL.n239 B 0.013505f
C762 VTAIL.n240 B 0.030147f
C763 VTAIL.n241 B 0.030147f
C764 VTAIL.n242 B 0.013505f
C765 VTAIL.n243 B 0.012755f
C766 VTAIL.n244 B 0.023736f
C767 VTAIL.n245 B 0.023736f
C768 VTAIL.n246 B 0.012755f
C769 VTAIL.n247 B 0.013505f
C770 VTAIL.n248 B 0.030147f
C771 VTAIL.n249 B 0.030147f
C772 VTAIL.n250 B 0.013505f
C773 VTAIL.n251 B 0.012755f
C774 VTAIL.n252 B 0.023736f
C775 VTAIL.n253 B 0.023736f
C776 VTAIL.n254 B 0.012755f
C777 VTAIL.n255 B 0.013505f
C778 VTAIL.n256 B 0.030147f
C779 VTAIL.n257 B 0.030147f
C780 VTAIL.n258 B 0.013505f
C781 VTAIL.n259 B 0.012755f
C782 VTAIL.n260 B 0.023736f
C783 VTAIL.n261 B 0.023736f
C784 VTAIL.n262 B 0.012755f
C785 VTAIL.n263 B 0.013505f
C786 VTAIL.n264 B 0.030147f
C787 VTAIL.n265 B 0.030147f
C788 VTAIL.n266 B 0.013505f
C789 VTAIL.n267 B 0.012755f
C790 VTAIL.n268 B 0.023736f
C791 VTAIL.n269 B 0.023736f
C792 VTAIL.n270 B 0.012755f
C793 VTAIL.n271 B 0.013505f
C794 VTAIL.n272 B 0.030147f
C795 VTAIL.n273 B 0.030147f
C796 VTAIL.n274 B 0.013505f
C797 VTAIL.n275 B 0.012755f
C798 VTAIL.n276 B 0.023736f
C799 VTAIL.n277 B 0.023736f
C800 VTAIL.n278 B 0.012755f
C801 VTAIL.n279 B 0.01313f
C802 VTAIL.n280 B 0.01313f
C803 VTAIL.n281 B 0.030147f
C804 VTAIL.n282 B 0.030147f
C805 VTAIL.n283 B 0.013505f
C806 VTAIL.n284 B 0.012755f
C807 VTAIL.n285 B 0.023736f
C808 VTAIL.n286 B 0.023736f
C809 VTAIL.n287 B 0.012755f
C810 VTAIL.n288 B 0.013505f
C811 VTAIL.n289 B 0.030147f
C812 VTAIL.n290 B 0.06498f
C813 VTAIL.n291 B 0.013505f
C814 VTAIL.n292 B 0.012755f
C815 VTAIL.n293 B 0.057134f
C816 VTAIL.n294 B 0.036398f
C817 VTAIL.n295 B 1.79252f
C818 VTAIL.n296 B 0.033202f
C819 VTAIL.n297 B 0.023736f
C820 VTAIL.n298 B 0.012755f
C821 VTAIL.n299 B 0.030147f
C822 VTAIL.n300 B 0.013505f
C823 VTAIL.n301 B 0.023736f
C824 VTAIL.n302 B 0.012755f
C825 VTAIL.n303 B 0.030147f
C826 VTAIL.n304 B 0.013505f
C827 VTAIL.n305 B 0.023736f
C828 VTAIL.n306 B 0.012755f
C829 VTAIL.n307 B 0.030147f
C830 VTAIL.n308 B 0.013505f
C831 VTAIL.n309 B 0.023736f
C832 VTAIL.n310 B 0.012755f
C833 VTAIL.n311 B 0.030147f
C834 VTAIL.n312 B 0.013505f
C835 VTAIL.n313 B 0.023736f
C836 VTAIL.n314 B 0.012755f
C837 VTAIL.n315 B 0.030147f
C838 VTAIL.n316 B 0.013505f
C839 VTAIL.n317 B 0.023736f
C840 VTAIL.n318 B 0.012755f
C841 VTAIL.n319 B 0.030147f
C842 VTAIL.n320 B 0.013505f
C843 VTAIL.n321 B 0.023736f
C844 VTAIL.n322 B 0.012755f
C845 VTAIL.n323 B 0.030147f
C846 VTAIL.n324 B 0.013505f
C847 VTAIL.n325 B 0.165938f
C848 VTAIL.t5 B 0.049861f
C849 VTAIL.n326 B 0.02261f
C850 VTAIL.n327 B 0.017809f
C851 VTAIL.n328 B 0.012755f
C852 VTAIL.n329 B 1.7477f
C853 VTAIL.n330 B 0.023736f
C854 VTAIL.n331 B 0.012755f
C855 VTAIL.n332 B 0.013505f
C856 VTAIL.n333 B 0.030147f
C857 VTAIL.n334 B 0.030147f
C858 VTAIL.n335 B 0.013505f
C859 VTAIL.n336 B 0.012755f
C860 VTAIL.n337 B 0.023736f
C861 VTAIL.n338 B 0.023736f
C862 VTAIL.n339 B 0.012755f
C863 VTAIL.n340 B 0.013505f
C864 VTAIL.n341 B 0.030147f
C865 VTAIL.n342 B 0.030147f
C866 VTAIL.n343 B 0.013505f
C867 VTAIL.n344 B 0.012755f
C868 VTAIL.n345 B 0.023736f
C869 VTAIL.n346 B 0.023736f
C870 VTAIL.n347 B 0.012755f
C871 VTAIL.n348 B 0.013505f
C872 VTAIL.n349 B 0.030147f
C873 VTAIL.n350 B 0.030147f
C874 VTAIL.n351 B 0.013505f
C875 VTAIL.n352 B 0.012755f
C876 VTAIL.n353 B 0.023736f
C877 VTAIL.n354 B 0.023736f
C878 VTAIL.n355 B 0.012755f
C879 VTAIL.n356 B 0.013505f
C880 VTAIL.n357 B 0.030147f
C881 VTAIL.n358 B 0.030147f
C882 VTAIL.n359 B 0.013505f
C883 VTAIL.n360 B 0.012755f
C884 VTAIL.n361 B 0.023736f
C885 VTAIL.n362 B 0.023736f
C886 VTAIL.n363 B 0.012755f
C887 VTAIL.n364 B 0.013505f
C888 VTAIL.n365 B 0.030147f
C889 VTAIL.n366 B 0.030147f
C890 VTAIL.n367 B 0.030147f
C891 VTAIL.n368 B 0.013505f
C892 VTAIL.n369 B 0.012755f
C893 VTAIL.n370 B 0.023736f
C894 VTAIL.n371 B 0.023736f
C895 VTAIL.n372 B 0.012755f
C896 VTAIL.n373 B 0.01313f
C897 VTAIL.n374 B 0.01313f
C898 VTAIL.n375 B 0.030147f
C899 VTAIL.n376 B 0.030147f
C900 VTAIL.n377 B 0.013505f
C901 VTAIL.n378 B 0.012755f
C902 VTAIL.n379 B 0.023736f
C903 VTAIL.n380 B 0.023736f
C904 VTAIL.n381 B 0.012755f
C905 VTAIL.n382 B 0.013505f
C906 VTAIL.n383 B 0.030147f
C907 VTAIL.n384 B 0.06498f
C908 VTAIL.n385 B 0.013505f
C909 VTAIL.n386 B 0.012755f
C910 VTAIL.n387 B 0.057134f
C911 VTAIL.n388 B 0.036398f
C912 VTAIL.n389 B 1.79252f
C913 VTAIL.t0 B 0.316425f
C914 VTAIL.t2 B 0.316425f
C915 VTAIL.n390 B 2.80649f
C916 VTAIL.n391 B 0.438189f
C917 VP.n0 B 0.03063f
C918 VP.t4 B 2.39024f
C919 VP.n1 B 0.020517f
C920 VP.n2 B 0.023233f
C921 VP.t7 B 2.39024f
C922 VP.n3 B 0.045506f
C923 VP.n4 B 0.023233f
C924 VP.t8 B 2.39024f
C925 VP.n5 B 0.834184f
C926 VP.n6 B 0.023233f
C927 VP.n7 B 0.045506f
C928 VP.n8 B 0.023233f
C929 VP.t1 B 2.39024f
C930 VP.n9 B 0.020517f
C931 VP.n10 B 0.03063f
C932 VP.t3 B 2.39024f
C933 VP.n11 B 0.03063f
C934 VP.t9 B 2.39024f
C935 VP.n12 B 0.020517f
C936 VP.n13 B 0.023233f
C937 VP.t5 B 2.39024f
C938 VP.n14 B 0.045506f
C939 VP.n15 B 0.023233f
C940 VP.t6 B 2.39024f
C941 VP.n16 B 0.834184f
C942 VP.n17 B 0.023233f
C943 VP.n18 B 0.045506f
C944 VP.t0 B 2.53864f
C945 VP.n19 B 0.88525f
C946 VP.t2 B 2.39024f
C947 VP.n20 B 0.896413f
C948 VP.n21 B 0.034749f
C949 VP.n22 B 0.19827f
C950 VP.n23 B 0.023233f
C951 VP.n24 B 0.023233f
C952 VP.n25 B 0.01897f
C953 VP.n26 B 0.04666f
C954 VP.n27 B 0.032611f
C955 VP.n28 B 0.023233f
C956 VP.n29 B 0.023233f
C957 VP.n30 B 0.032611f
C958 VP.n31 B 0.04666f
C959 VP.n32 B 0.01897f
C960 VP.n33 B 0.023233f
C961 VP.n34 B 0.023233f
C962 VP.n35 B 0.023233f
C963 VP.n36 B 0.034749f
C964 VP.n37 B 0.834184f
C965 VP.n38 B 0.030473f
C966 VP.n39 B 0.046901f
C967 VP.n40 B 0.023233f
C968 VP.n41 B 0.023233f
C969 VP.n42 B 0.023233f
C970 VP.n43 B 0.043717f
C971 VP.n44 B 0.036887f
C972 VP.n45 B 0.909318f
C973 VP.n46 B 1.46702f
C974 VP.n47 B 1.48227f
C975 VP.n48 B 0.909318f
C976 VP.n49 B 0.036887f
C977 VP.n50 B 0.043717f
C978 VP.n51 B 0.023233f
C979 VP.n52 B 0.023233f
C980 VP.n53 B 0.023233f
C981 VP.n54 B 0.046901f
C982 VP.n55 B 0.030473f
C983 VP.n56 B 0.834184f
C984 VP.n57 B 0.034749f
C985 VP.n58 B 0.023233f
C986 VP.n59 B 0.023233f
C987 VP.n60 B 0.023233f
C988 VP.n61 B 0.01897f
C989 VP.n62 B 0.04666f
C990 VP.n63 B 0.032611f
C991 VP.n64 B 0.023233f
C992 VP.n65 B 0.023233f
C993 VP.n66 B 0.032611f
C994 VP.n67 B 0.04666f
C995 VP.n68 B 0.01897f
C996 VP.n69 B 0.023233f
C997 VP.n70 B 0.023233f
C998 VP.n71 B 0.023233f
C999 VP.n72 B 0.034749f
C1000 VP.n73 B 0.834184f
C1001 VP.n74 B 0.030473f
C1002 VP.n75 B 0.046901f
C1003 VP.n76 B 0.023233f
C1004 VP.n77 B 0.023233f
C1005 VP.n78 B 0.023233f
C1006 VP.n79 B 0.043717f
C1007 VP.n80 B 0.036887f
C1008 VP.n81 B 0.909318f
C1009 VP.n82 B 0.030943f
.ends

