* NGSPICE file created from diff_pair_sample_1724.ext - technology: sky130A

.subckt diff_pair_sample_1724 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=2.78685 ps=17.22 w=16.89 l=3.68
X1 B.t20 B.t18 B.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=0 ps=0 w=16.89 l=3.68
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=0 ps=0 w=16.89 l=3.68
X3 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X4 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=0 ps=0 w=16.89 l=3.68
X5 VTAIL.t7 VN.t1 VDD2.t8 B.t23 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X6 VTAIL.t9 VN.t2 VDD2.t7 B.t22 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X7 VTAIL.t6 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X8 VTAIL.t17 VP.t2 VDD1.t7 B.t23 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X9 VTAIL.t12 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X10 VTAIL.t8 VN.t4 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X11 VTAIL.t4 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X12 VDD2.t4 VN.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=6.5871 ps=34.56 w=16.89 l=3.68
X13 VDD2.t3 VN.t6 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X14 VDD1.t5 VP.t4 VTAIL.t19 B.t21 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=6.5871 ps=34.56 w=16.89 l=3.68
X15 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=2.78685 ps=17.22 w=16.89 l=3.68
X16 VDD1.t3 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=6.5871 ps=34.56 w=16.89 l=3.68
X17 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=0 ps=0 w=16.89 l=3.68
X18 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=2.78685 ps=17.22 w=16.89 l=3.68
X19 VDD2.t2 VN.t7 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X20 VDD2.t1 VN.t8 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5871 pd=34.56 as=2.78685 ps=17.22 w=16.89 l=3.68
X21 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X22 VTAIL.t18 VP.t9 VDD1.t0 B.t22 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=2.78685 ps=17.22 w=16.89 l=3.68
X23 VDD2.t0 VN.t9 VTAIL.t16 B.t21 sky130_fd_pr__nfet_01v8 ad=2.78685 pd=17.22 as=6.5871 ps=34.56 w=16.89 l=3.68
R0 VN.n108 VN.n107 161.3
R1 VN.n106 VN.n56 161.3
R2 VN.n105 VN.n104 161.3
R3 VN.n103 VN.n57 161.3
R4 VN.n102 VN.n101 161.3
R5 VN.n100 VN.n58 161.3
R6 VN.n99 VN.n98 161.3
R7 VN.n97 VN.n59 161.3
R8 VN.n96 VN.n95 161.3
R9 VN.n94 VN.n60 161.3
R10 VN.n93 VN.n92 161.3
R11 VN.n91 VN.n62 161.3
R12 VN.n90 VN.n89 161.3
R13 VN.n88 VN.n63 161.3
R14 VN.n87 VN.n86 161.3
R15 VN.n85 VN.n64 161.3
R16 VN.n84 VN.n83 161.3
R17 VN.n82 VN.n65 161.3
R18 VN.n81 VN.n80 161.3
R19 VN.n79 VN.n66 161.3
R20 VN.n78 VN.n77 161.3
R21 VN.n76 VN.n67 161.3
R22 VN.n75 VN.n74 161.3
R23 VN.n73 VN.n68 161.3
R24 VN.n72 VN.n71 161.3
R25 VN.n53 VN.n52 161.3
R26 VN.n51 VN.n1 161.3
R27 VN.n50 VN.n49 161.3
R28 VN.n48 VN.n2 161.3
R29 VN.n47 VN.n46 161.3
R30 VN.n45 VN.n3 161.3
R31 VN.n44 VN.n43 161.3
R32 VN.n42 VN.n4 161.3
R33 VN.n41 VN.n40 161.3
R34 VN.n38 VN.n5 161.3
R35 VN.n37 VN.n36 161.3
R36 VN.n35 VN.n6 161.3
R37 VN.n34 VN.n33 161.3
R38 VN.n32 VN.n7 161.3
R39 VN.n31 VN.n30 161.3
R40 VN.n29 VN.n8 161.3
R41 VN.n28 VN.n27 161.3
R42 VN.n26 VN.n9 161.3
R43 VN.n25 VN.n24 161.3
R44 VN.n23 VN.n10 161.3
R45 VN.n22 VN.n21 161.3
R46 VN.n20 VN.n11 161.3
R47 VN.n19 VN.n18 161.3
R48 VN.n17 VN.n12 161.3
R49 VN.n16 VN.n15 161.3
R50 VN.n69 VN.t5 141.933
R51 VN.n13 VN.t8 141.933
R52 VN.n27 VN.t7 110.612
R53 VN.n14 VN.t3 110.612
R54 VN.n39 VN.t2 110.612
R55 VN.n0 VN.t9 110.612
R56 VN.n83 VN.t6 110.612
R57 VN.n70 VN.t4 110.612
R58 VN.n61 VN.t1 110.612
R59 VN.n55 VN.t0 110.612
R60 VN.n54 VN.n0 89.0887
R61 VN.n109 VN.n55 89.0887
R62 VN.n14 VN.n13 74.5304
R63 VN.n70 VN.n69 74.5304
R64 VN VN.n109 62.8503
R65 VN.n46 VN.n2 41.9503
R66 VN.n101 VN.n57 41.9503
R67 VN.n21 VN.n20 40.979
R68 VN.n33 VN.n6 40.979
R69 VN.n77 VN.n76 40.979
R70 VN.n89 VN.n62 40.979
R71 VN.n21 VN.n10 40.0078
R72 VN.n33 VN.n32 40.0078
R73 VN.n77 VN.n66 40.0078
R74 VN.n89 VN.n88 40.0078
R75 VN.n46 VN.n45 39.0365
R76 VN.n101 VN.n100 39.0365
R77 VN.n15 VN.n12 24.4675
R78 VN.n19 VN.n12 24.4675
R79 VN.n20 VN.n19 24.4675
R80 VN.n25 VN.n10 24.4675
R81 VN.n26 VN.n25 24.4675
R82 VN.n27 VN.n26 24.4675
R83 VN.n27 VN.n8 24.4675
R84 VN.n31 VN.n8 24.4675
R85 VN.n32 VN.n31 24.4675
R86 VN.n37 VN.n6 24.4675
R87 VN.n38 VN.n37 24.4675
R88 VN.n40 VN.n38 24.4675
R89 VN.n44 VN.n4 24.4675
R90 VN.n45 VN.n44 24.4675
R91 VN.n50 VN.n2 24.4675
R92 VN.n51 VN.n50 24.4675
R93 VN.n52 VN.n51 24.4675
R94 VN.n76 VN.n75 24.4675
R95 VN.n75 VN.n68 24.4675
R96 VN.n71 VN.n68 24.4675
R97 VN.n88 VN.n87 24.4675
R98 VN.n87 VN.n64 24.4675
R99 VN.n83 VN.n64 24.4675
R100 VN.n83 VN.n82 24.4675
R101 VN.n82 VN.n81 24.4675
R102 VN.n81 VN.n66 24.4675
R103 VN.n100 VN.n99 24.4675
R104 VN.n99 VN.n59 24.4675
R105 VN.n95 VN.n94 24.4675
R106 VN.n94 VN.n93 24.4675
R107 VN.n93 VN.n62 24.4675
R108 VN.n107 VN.n106 24.4675
R109 VN.n106 VN.n105 24.4675
R110 VN.n105 VN.n57 24.4675
R111 VN.n39 VN.n4 23.9782
R112 VN.n61 VN.n59 23.9782
R113 VN.n16 VN.n13 3.44123
R114 VN.n72 VN.n69 3.44123
R115 VN.n52 VN.n0 0.97918
R116 VN.n107 VN.n55 0.97918
R117 VN.n15 VN.n14 0.48984
R118 VN.n40 VN.n39 0.48984
R119 VN.n71 VN.n70 0.48984
R120 VN.n95 VN.n61 0.48984
R121 VN.n109 VN.n108 0.354971
R122 VN.n54 VN.n53 0.354971
R123 VN VN.n54 0.26696
R124 VN.n108 VN.n56 0.189894
R125 VN.n104 VN.n56 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n102 0.189894
R128 VN.n102 VN.n58 0.189894
R129 VN.n98 VN.n58 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n96 0.189894
R132 VN.n96 VN.n60 0.189894
R133 VN.n92 VN.n60 0.189894
R134 VN.n92 VN.n91 0.189894
R135 VN.n91 VN.n90 0.189894
R136 VN.n90 VN.n63 0.189894
R137 VN.n86 VN.n63 0.189894
R138 VN.n86 VN.n85 0.189894
R139 VN.n85 VN.n84 0.189894
R140 VN.n84 VN.n65 0.189894
R141 VN.n80 VN.n65 0.189894
R142 VN.n80 VN.n79 0.189894
R143 VN.n79 VN.n78 0.189894
R144 VN.n78 VN.n67 0.189894
R145 VN.n74 VN.n67 0.189894
R146 VN.n74 VN.n73 0.189894
R147 VN.n73 VN.n72 0.189894
R148 VN.n17 VN.n16 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n18 VN.n11 0.189894
R151 VN.n22 VN.n11 0.189894
R152 VN.n23 VN.n22 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n24 VN.n9 0.189894
R155 VN.n28 VN.n9 0.189894
R156 VN.n29 VN.n28 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n30 VN.n7 0.189894
R159 VN.n34 VN.n7 0.189894
R160 VN.n35 VN.n34 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n36 VN.n5 0.189894
R163 VN.n41 VN.n5 0.189894
R164 VN.n42 VN.n41 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n43 VN.n3 0.189894
R167 VN.n47 VN.n3 0.189894
R168 VN.n48 VN.n47 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n49 VN.n1 0.189894
R171 VN.n53 VN.n1 0.189894
R172 VTAIL.n384 VTAIL.n296 289.615
R173 VTAIL.n90 VTAIL.n2 289.615
R174 VTAIL.n290 VTAIL.n202 289.615
R175 VTAIL.n192 VTAIL.n104 289.615
R176 VTAIL.n327 VTAIL.n326 185
R177 VTAIL.n324 VTAIL.n323 185
R178 VTAIL.n333 VTAIL.n332 185
R179 VTAIL.n335 VTAIL.n334 185
R180 VTAIL.n320 VTAIL.n319 185
R181 VTAIL.n341 VTAIL.n340 185
R182 VTAIL.n343 VTAIL.n342 185
R183 VTAIL.n316 VTAIL.n315 185
R184 VTAIL.n349 VTAIL.n348 185
R185 VTAIL.n351 VTAIL.n350 185
R186 VTAIL.n312 VTAIL.n311 185
R187 VTAIL.n357 VTAIL.n356 185
R188 VTAIL.n359 VTAIL.n358 185
R189 VTAIL.n308 VTAIL.n307 185
R190 VTAIL.n365 VTAIL.n364 185
R191 VTAIL.n368 VTAIL.n367 185
R192 VTAIL.n366 VTAIL.n304 185
R193 VTAIL.n373 VTAIL.n303 185
R194 VTAIL.n375 VTAIL.n374 185
R195 VTAIL.n377 VTAIL.n376 185
R196 VTAIL.n300 VTAIL.n299 185
R197 VTAIL.n383 VTAIL.n382 185
R198 VTAIL.n385 VTAIL.n384 185
R199 VTAIL.n33 VTAIL.n32 185
R200 VTAIL.n30 VTAIL.n29 185
R201 VTAIL.n39 VTAIL.n38 185
R202 VTAIL.n41 VTAIL.n40 185
R203 VTAIL.n26 VTAIL.n25 185
R204 VTAIL.n47 VTAIL.n46 185
R205 VTAIL.n49 VTAIL.n48 185
R206 VTAIL.n22 VTAIL.n21 185
R207 VTAIL.n55 VTAIL.n54 185
R208 VTAIL.n57 VTAIL.n56 185
R209 VTAIL.n18 VTAIL.n17 185
R210 VTAIL.n63 VTAIL.n62 185
R211 VTAIL.n65 VTAIL.n64 185
R212 VTAIL.n14 VTAIL.n13 185
R213 VTAIL.n71 VTAIL.n70 185
R214 VTAIL.n74 VTAIL.n73 185
R215 VTAIL.n72 VTAIL.n10 185
R216 VTAIL.n79 VTAIL.n9 185
R217 VTAIL.n81 VTAIL.n80 185
R218 VTAIL.n83 VTAIL.n82 185
R219 VTAIL.n6 VTAIL.n5 185
R220 VTAIL.n89 VTAIL.n88 185
R221 VTAIL.n91 VTAIL.n90 185
R222 VTAIL.n291 VTAIL.n290 185
R223 VTAIL.n289 VTAIL.n288 185
R224 VTAIL.n206 VTAIL.n205 185
R225 VTAIL.n283 VTAIL.n282 185
R226 VTAIL.n281 VTAIL.n280 185
R227 VTAIL.n279 VTAIL.n209 185
R228 VTAIL.n213 VTAIL.n210 185
R229 VTAIL.n274 VTAIL.n273 185
R230 VTAIL.n272 VTAIL.n271 185
R231 VTAIL.n215 VTAIL.n214 185
R232 VTAIL.n266 VTAIL.n265 185
R233 VTAIL.n264 VTAIL.n263 185
R234 VTAIL.n219 VTAIL.n218 185
R235 VTAIL.n258 VTAIL.n257 185
R236 VTAIL.n256 VTAIL.n255 185
R237 VTAIL.n223 VTAIL.n222 185
R238 VTAIL.n250 VTAIL.n249 185
R239 VTAIL.n248 VTAIL.n247 185
R240 VTAIL.n227 VTAIL.n226 185
R241 VTAIL.n242 VTAIL.n241 185
R242 VTAIL.n240 VTAIL.n239 185
R243 VTAIL.n231 VTAIL.n230 185
R244 VTAIL.n234 VTAIL.n233 185
R245 VTAIL.n193 VTAIL.n192 185
R246 VTAIL.n191 VTAIL.n190 185
R247 VTAIL.n108 VTAIL.n107 185
R248 VTAIL.n185 VTAIL.n184 185
R249 VTAIL.n183 VTAIL.n182 185
R250 VTAIL.n181 VTAIL.n111 185
R251 VTAIL.n115 VTAIL.n112 185
R252 VTAIL.n176 VTAIL.n175 185
R253 VTAIL.n174 VTAIL.n173 185
R254 VTAIL.n117 VTAIL.n116 185
R255 VTAIL.n168 VTAIL.n167 185
R256 VTAIL.n166 VTAIL.n165 185
R257 VTAIL.n121 VTAIL.n120 185
R258 VTAIL.n160 VTAIL.n159 185
R259 VTAIL.n158 VTAIL.n157 185
R260 VTAIL.n125 VTAIL.n124 185
R261 VTAIL.n152 VTAIL.n151 185
R262 VTAIL.n150 VTAIL.n149 185
R263 VTAIL.n129 VTAIL.n128 185
R264 VTAIL.n144 VTAIL.n143 185
R265 VTAIL.n142 VTAIL.n141 185
R266 VTAIL.n133 VTAIL.n132 185
R267 VTAIL.n136 VTAIL.n135 185
R268 VTAIL.t19 VTAIL.n232 147.659
R269 VTAIL.t10 VTAIL.n134 147.659
R270 VTAIL.t16 VTAIL.n325 147.659
R271 VTAIL.t1 VTAIL.n31 147.659
R272 VTAIL.n326 VTAIL.n323 104.615
R273 VTAIL.n333 VTAIL.n323 104.615
R274 VTAIL.n334 VTAIL.n333 104.615
R275 VTAIL.n334 VTAIL.n319 104.615
R276 VTAIL.n341 VTAIL.n319 104.615
R277 VTAIL.n342 VTAIL.n341 104.615
R278 VTAIL.n342 VTAIL.n315 104.615
R279 VTAIL.n349 VTAIL.n315 104.615
R280 VTAIL.n350 VTAIL.n349 104.615
R281 VTAIL.n350 VTAIL.n311 104.615
R282 VTAIL.n357 VTAIL.n311 104.615
R283 VTAIL.n358 VTAIL.n357 104.615
R284 VTAIL.n358 VTAIL.n307 104.615
R285 VTAIL.n365 VTAIL.n307 104.615
R286 VTAIL.n367 VTAIL.n365 104.615
R287 VTAIL.n367 VTAIL.n366 104.615
R288 VTAIL.n366 VTAIL.n303 104.615
R289 VTAIL.n375 VTAIL.n303 104.615
R290 VTAIL.n376 VTAIL.n375 104.615
R291 VTAIL.n376 VTAIL.n299 104.615
R292 VTAIL.n383 VTAIL.n299 104.615
R293 VTAIL.n384 VTAIL.n383 104.615
R294 VTAIL.n32 VTAIL.n29 104.615
R295 VTAIL.n39 VTAIL.n29 104.615
R296 VTAIL.n40 VTAIL.n39 104.615
R297 VTAIL.n40 VTAIL.n25 104.615
R298 VTAIL.n47 VTAIL.n25 104.615
R299 VTAIL.n48 VTAIL.n47 104.615
R300 VTAIL.n48 VTAIL.n21 104.615
R301 VTAIL.n55 VTAIL.n21 104.615
R302 VTAIL.n56 VTAIL.n55 104.615
R303 VTAIL.n56 VTAIL.n17 104.615
R304 VTAIL.n63 VTAIL.n17 104.615
R305 VTAIL.n64 VTAIL.n63 104.615
R306 VTAIL.n64 VTAIL.n13 104.615
R307 VTAIL.n71 VTAIL.n13 104.615
R308 VTAIL.n73 VTAIL.n71 104.615
R309 VTAIL.n73 VTAIL.n72 104.615
R310 VTAIL.n72 VTAIL.n9 104.615
R311 VTAIL.n81 VTAIL.n9 104.615
R312 VTAIL.n82 VTAIL.n81 104.615
R313 VTAIL.n82 VTAIL.n5 104.615
R314 VTAIL.n89 VTAIL.n5 104.615
R315 VTAIL.n90 VTAIL.n89 104.615
R316 VTAIL.n290 VTAIL.n289 104.615
R317 VTAIL.n289 VTAIL.n205 104.615
R318 VTAIL.n282 VTAIL.n205 104.615
R319 VTAIL.n282 VTAIL.n281 104.615
R320 VTAIL.n281 VTAIL.n209 104.615
R321 VTAIL.n213 VTAIL.n209 104.615
R322 VTAIL.n273 VTAIL.n213 104.615
R323 VTAIL.n273 VTAIL.n272 104.615
R324 VTAIL.n272 VTAIL.n214 104.615
R325 VTAIL.n265 VTAIL.n214 104.615
R326 VTAIL.n265 VTAIL.n264 104.615
R327 VTAIL.n264 VTAIL.n218 104.615
R328 VTAIL.n257 VTAIL.n218 104.615
R329 VTAIL.n257 VTAIL.n256 104.615
R330 VTAIL.n256 VTAIL.n222 104.615
R331 VTAIL.n249 VTAIL.n222 104.615
R332 VTAIL.n249 VTAIL.n248 104.615
R333 VTAIL.n248 VTAIL.n226 104.615
R334 VTAIL.n241 VTAIL.n226 104.615
R335 VTAIL.n241 VTAIL.n240 104.615
R336 VTAIL.n240 VTAIL.n230 104.615
R337 VTAIL.n233 VTAIL.n230 104.615
R338 VTAIL.n192 VTAIL.n191 104.615
R339 VTAIL.n191 VTAIL.n107 104.615
R340 VTAIL.n184 VTAIL.n107 104.615
R341 VTAIL.n184 VTAIL.n183 104.615
R342 VTAIL.n183 VTAIL.n111 104.615
R343 VTAIL.n115 VTAIL.n111 104.615
R344 VTAIL.n175 VTAIL.n115 104.615
R345 VTAIL.n175 VTAIL.n174 104.615
R346 VTAIL.n174 VTAIL.n116 104.615
R347 VTAIL.n167 VTAIL.n116 104.615
R348 VTAIL.n167 VTAIL.n166 104.615
R349 VTAIL.n166 VTAIL.n120 104.615
R350 VTAIL.n159 VTAIL.n120 104.615
R351 VTAIL.n159 VTAIL.n158 104.615
R352 VTAIL.n158 VTAIL.n124 104.615
R353 VTAIL.n151 VTAIL.n124 104.615
R354 VTAIL.n151 VTAIL.n150 104.615
R355 VTAIL.n150 VTAIL.n128 104.615
R356 VTAIL.n143 VTAIL.n128 104.615
R357 VTAIL.n143 VTAIL.n142 104.615
R358 VTAIL.n142 VTAIL.n132 104.615
R359 VTAIL.n135 VTAIL.n132 104.615
R360 VTAIL.n326 VTAIL.t16 52.3082
R361 VTAIL.n32 VTAIL.t1 52.3082
R362 VTAIL.n233 VTAIL.t19 52.3082
R363 VTAIL.n135 VTAIL.t10 52.3082
R364 VTAIL.n201 VTAIL.n200 45.7915
R365 VTAIL.n199 VTAIL.n198 45.7915
R366 VTAIL.n103 VTAIL.n102 45.7915
R367 VTAIL.n101 VTAIL.n100 45.7915
R368 VTAIL.n391 VTAIL.n390 45.7913
R369 VTAIL.n1 VTAIL.n0 45.7913
R370 VTAIL.n97 VTAIL.n96 45.7913
R371 VTAIL.n99 VTAIL.n98 45.7913
R372 VTAIL.n389 VTAIL.n388 33.9308
R373 VTAIL.n95 VTAIL.n94 33.9308
R374 VTAIL.n295 VTAIL.n294 33.9308
R375 VTAIL.n197 VTAIL.n196 33.9308
R376 VTAIL.n101 VTAIL.n99 33.841
R377 VTAIL.n389 VTAIL.n295 30.3841
R378 VTAIL.n327 VTAIL.n325 15.6677
R379 VTAIL.n33 VTAIL.n31 15.6677
R380 VTAIL.n234 VTAIL.n232 15.6677
R381 VTAIL.n136 VTAIL.n134 15.6677
R382 VTAIL.n374 VTAIL.n373 13.1884
R383 VTAIL.n80 VTAIL.n79 13.1884
R384 VTAIL.n280 VTAIL.n279 13.1884
R385 VTAIL.n182 VTAIL.n181 13.1884
R386 VTAIL.n328 VTAIL.n324 12.8005
R387 VTAIL.n372 VTAIL.n304 12.8005
R388 VTAIL.n377 VTAIL.n302 12.8005
R389 VTAIL.n34 VTAIL.n30 12.8005
R390 VTAIL.n78 VTAIL.n10 12.8005
R391 VTAIL.n83 VTAIL.n8 12.8005
R392 VTAIL.n283 VTAIL.n208 12.8005
R393 VTAIL.n278 VTAIL.n210 12.8005
R394 VTAIL.n235 VTAIL.n231 12.8005
R395 VTAIL.n185 VTAIL.n110 12.8005
R396 VTAIL.n180 VTAIL.n112 12.8005
R397 VTAIL.n137 VTAIL.n133 12.8005
R398 VTAIL.n332 VTAIL.n331 12.0247
R399 VTAIL.n369 VTAIL.n368 12.0247
R400 VTAIL.n378 VTAIL.n300 12.0247
R401 VTAIL.n38 VTAIL.n37 12.0247
R402 VTAIL.n75 VTAIL.n74 12.0247
R403 VTAIL.n84 VTAIL.n6 12.0247
R404 VTAIL.n284 VTAIL.n206 12.0247
R405 VTAIL.n275 VTAIL.n274 12.0247
R406 VTAIL.n239 VTAIL.n238 12.0247
R407 VTAIL.n186 VTAIL.n108 12.0247
R408 VTAIL.n177 VTAIL.n176 12.0247
R409 VTAIL.n141 VTAIL.n140 12.0247
R410 VTAIL.n335 VTAIL.n322 11.249
R411 VTAIL.n364 VTAIL.n306 11.249
R412 VTAIL.n382 VTAIL.n381 11.249
R413 VTAIL.n41 VTAIL.n28 11.249
R414 VTAIL.n70 VTAIL.n12 11.249
R415 VTAIL.n88 VTAIL.n87 11.249
R416 VTAIL.n288 VTAIL.n287 11.249
R417 VTAIL.n271 VTAIL.n212 11.249
R418 VTAIL.n242 VTAIL.n229 11.249
R419 VTAIL.n190 VTAIL.n189 11.249
R420 VTAIL.n173 VTAIL.n114 11.249
R421 VTAIL.n144 VTAIL.n131 11.249
R422 VTAIL.n336 VTAIL.n320 10.4732
R423 VTAIL.n363 VTAIL.n308 10.4732
R424 VTAIL.n385 VTAIL.n298 10.4732
R425 VTAIL.n42 VTAIL.n26 10.4732
R426 VTAIL.n69 VTAIL.n14 10.4732
R427 VTAIL.n91 VTAIL.n4 10.4732
R428 VTAIL.n291 VTAIL.n204 10.4732
R429 VTAIL.n270 VTAIL.n215 10.4732
R430 VTAIL.n243 VTAIL.n227 10.4732
R431 VTAIL.n193 VTAIL.n106 10.4732
R432 VTAIL.n172 VTAIL.n117 10.4732
R433 VTAIL.n145 VTAIL.n129 10.4732
R434 VTAIL.n340 VTAIL.n339 9.69747
R435 VTAIL.n360 VTAIL.n359 9.69747
R436 VTAIL.n386 VTAIL.n296 9.69747
R437 VTAIL.n46 VTAIL.n45 9.69747
R438 VTAIL.n66 VTAIL.n65 9.69747
R439 VTAIL.n92 VTAIL.n2 9.69747
R440 VTAIL.n292 VTAIL.n202 9.69747
R441 VTAIL.n267 VTAIL.n266 9.69747
R442 VTAIL.n247 VTAIL.n246 9.69747
R443 VTAIL.n194 VTAIL.n104 9.69747
R444 VTAIL.n169 VTAIL.n168 9.69747
R445 VTAIL.n149 VTAIL.n148 9.69747
R446 VTAIL.n388 VTAIL.n387 9.45567
R447 VTAIL.n94 VTAIL.n93 9.45567
R448 VTAIL.n294 VTAIL.n293 9.45567
R449 VTAIL.n196 VTAIL.n195 9.45567
R450 VTAIL.n387 VTAIL.n386 9.3005
R451 VTAIL.n298 VTAIL.n297 9.3005
R452 VTAIL.n381 VTAIL.n380 9.3005
R453 VTAIL.n379 VTAIL.n378 9.3005
R454 VTAIL.n302 VTAIL.n301 9.3005
R455 VTAIL.n347 VTAIL.n346 9.3005
R456 VTAIL.n345 VTAIL.n344 9.3005
R457 VTAIL.n318 VTAIL.n317 9.3005
R458 VTAIL.n339 VTAIL.n338 9.3005
R459 VTAIL.n337 VTAIL.n336 9.3005
R460 VTAIL.n322 VTAIL.n321 9.3005
R461 VTAIL.n331 VTAIL.n330 9.3005
R462 VTAIL.n329 VTAIL.n328 9.3005
R463 VTAIL.n314 VTAIL.n313 9.3005
R464 VTAIL.n353 VTAIL.n352 9.3005
R465 VTAIL.n355 VTAIL.n354 9.3005
R466 VTAIL.n310 VTAIL.n309 9.3005
R467 VTAIL.n361 VTAIL.n360 9.3005
R468 VTAIL.n363 VTAIL.n362 9.3005
R469 VTAIL.n306 VTAIL.n305 9.3005
R470 VTAIL.n370 VTAIL.n369 9.3005
R471 VTAIL.n372 VTAIL.n371 9.3005
R472 VTAIL.n93 VTAIL.n92 9.3005
R473 VTAIL.n4 VTAIL.n3 9.3005
R474 VTAIL.n87 VTAIL.n86 9.3005
R475 VTAIL.n85 VTAIL.n84 9.3005
R476 VTAIL.n8 VTAIL.n7 9.3005
R477 VTAIL.n53 VTAIL.n52 9.3005
R478 VTAIL.n51 VTAIL.n50 9.3005
R479 VTAIL.n24 VTAIL.n23 9.3005
R480 VTAIL.n45 VTAIL.n44 9.3005
R481 VTAIL.n43 VTAIL.n42 9.3005
R482 VTAIL.n28 VTAIL.n27 9.3005
R483 VTAIL.n37 VTAIL.n36 9.3005
R484 VTAIL.n35 VTAIL.n34 9.3005
R485 VTAIL.n20 VTAIL.n19 9.3005
R486 VTAIL.n59 VTAIL.n58 9.3005
R487 VTAIL.n61 VTAIL.n60 9.3005
R488 VTAIL.n16 VTAIL.n15 9.3005
R489 VTAIL.n67 VTAIL.n66 9.3005
R490 VTAIL.n69 VTAIL.n68 9.3005
R491 VTAIL.n12 VTAIL.n11 9.3005
R492 VTAIL.n76 VTAIL.n75 9.3005
R493 VTAIL.n78 VTAIL.n77 9.3005
R494 VTAIL.n260 VTAIL.n259 9.3005
R495 VTAIL.n262 VTAIL.n261 9.3005
R496 VTAIL.n217 VTAIL.n216 9.3005
R497 VTAIL.n268 VTAIL.n267 9.3005
R498 VTAIL.n270 VTAIL.n269 9.3005
R499 VTAIL.n212 VTAIL.n211 9.3005
R500 VTAIL.n276 VTAIL.n275 9.3005
R501 VTAIL.n278 VTAIL.n277 9.3005
R502 VTAIL.n293 VTAIL.n292 9.3005
R503 VTAIL.n204 VTAIL.n203 9.3005
R504 VTAIL.n287 VTAIL.n286 9.3005
R505 VTAIL.n285 VTAIL.n284 9.3005
R506 VTAIL.n208 VTAIL.n207 9.3005
R507 VTAIL.n221 VTAIL.n220 9.3005
R508 VTAIL.n254 VTAIL.n253 9.3005
R509 VTAIL.n252 VTAIL.n251 9.3005
R510 VTAIL.n225 VTAIL.n224 9.3005
R511 VTAIL.n246 VTAIL.n245 9.3005
R512 VTAIL.n244 VTAIL.n243 9.3005
R513 VTAIL.n229 VTAIL.n228 9.3005
R514 VTAIL.n238 VTAIL.n237 9.3005
R515 VTAIL.n236 VTAIL.n235 9.3005
R516 VTAIL.n162 VTAIL.n161 9.3005
R517 VTAIL.n164 VTAIL.n163 9.3005
R518 VTAIL.n119 VTAIL.n118 9.3005
R519 VTAIL.n170 VTAIL.n169 9.3005
R520 VTAIL.n172 VTAIL.n171 9.3005
R521 VTAIL.n114 VTAIL.n113 9.3005
R522 VTAIL.n178 VTAIL.n177 9.3005
R523 VTAIL.n180 VTAIL.n179 9.3005
R524 VTAIL.n195 VTAIL.n194 9.3005
R525 VTAIL.n106 VTAIL.n105 9.3005
R526 VTAIL.n189 VTAIL.n188 9.3005
R527 VTAIL.n187 VTAIL.n186 9.3005
R528 VTAIL.n110 VTAIL.n109 9.3005
R529 VTAIL.n123 VTAIL.n122 9.3005
R530 VTAIL.n156 VTAIL.n155 9.3005
R531 VTAIL.n154 VTAIL.n153 9.3005
R532 VTAIL.n127 VTAIL.n126 9.3005
R533 VTAIL.n148 VTAIL.n147 9.3005
R534 VTAIL.n146 VTAIL.n145 9.3005
R535 VTAIL.n131 VTAIL.n130 9.3005
R536 VTAIL.n140 VTAIL.n139 9.3005
R537 VTAIL.n138 VTAIL.n137 9.3005
R538 VTAIL.n343 VTAIL.n318 8.92171
R539 VTAIL.n356 VTAIL.n310 8.92171
R540 VTAIL.n49 VTAIL.n24 8.92171
R541 VTAIL.n62 VTAIL.n16 8.92171
R542 VTAIL.n263 VTAIL.n217 8.92171
R543 VTAIL.n250 VTAIL.n225 8.92171
R544 VTAIL.n165 VTAIL.n119 8.92171
R545 VTAIL.n152 VTAIL.n127 8.92171
R546 VTAIL.n344 VTAIL.n316 8.14595
R547 VTAIL.n355 VTAIL.n312 8.14595
R548 VTAIL.n50 VTAIL.n22 8.14595
R549 VTAIL.n61 VTAIL.n18 8.14595
R550 VTAIL.n262 VTAIL.n219 8.14595
R551 VTAIL.n251 VTAIL.n223 8.14595
R552 VTAIL.n164 VTAIL.n121 8.14595
R553 VTAIL.n153 VTAIL.n125 8.14595
R554 VTAIL.n348 VTAIL.n347 7.3702
R555 VTAIL.n352 VTAIL.n351 7.3702
R556 VTAIL.n54 VTAIL.n53 7.3702
R557 VTAIL.n58 VTAIL.n57 7.3702
R558 VTAIL.n259 VTAIL.n258 7.3702
R559 VTAIL.n255 VTAIL.n254 7.3702
R560 VTAIL.n161 VTAIL.n160 7.3702
R561 VTAIL.n157 VTAIL.n156 7.3702
R562 VTAIL.n348 VTAIL.n314 6.59444
R563 VTAIL.n351 VTAIL.n314 6.59444
R564 VTAIL.n54 VTAIL.n20 6.59444
R565 VTAIL.n57 VTAIL.n20 6.59444
R566 VTAIL.n258 VTAIL.n221 6.59444
R567 VTAIL.n255 VTAIL.n221 6.59444
R568 VTAIL.n160 VTAIL.n123 6.59444
R569 VTAIL.n157 VTAIL.n123 6.59444
R570 VTAIL.n347 VTAIL.n316 5.81868
R571 VTAIL.n352 VTAIL.n312 5.81868
R572 VTAIL.n53 VTAIL.n22 5.81868
R573 VTAIL.n58 VTAIL.n18 5.81868
R574 VTAIL.n259 VTAIL.n219 5.81868
R575 VTAIL.n254 VTAIL.n223 5.81868
R576 VTAIL.n161 VTAIL.n121 5.81868
R577 VTAIL.n156 VTAIL.n125 5.81868
R578 VTAIL.n344 VTAIL.n343 5.04292
R579 VTAIL.n356 VTAIL.n355 5.04292
R580 VTAIL.n50 VTAIL.n49 5.04292
R581 VTAIL.n62 VTAIL.n61 5.04292
R582 VTAIL.n263 VTAIL.n262 5.04292
R583 VTAIL.n251 VTAIL.n250 5.04292
R584 VTAIL.n165 VTAIL.n164 5.04292
R585 VTAIL.n153 VTAIL.n152 5.04292
R586 VTAIL.n236 VTAIL.n232 4.38563
R587 VTAIL.n138 VTAIL.n134 4.38563
R588 VTAIL.n329 VTAIL.n325 4.38563
R589 VTAIL.n35 VTAIL.n31 4.38563
R590 VTAIL.n340 VTAIL.n318 4.26717
R591 VTAIL.n359 VTAIL.n310 4.26717
R592 VTAIL.n388 VTAIL.n296 4.26717
R593 VTAIL.n46 VTAIL.n24 4.26717
R594 VTAIL.n65 VTAIL.n16 4.26717
R595 VTAIL.n94 VTAIL.n2 4.26717
R596 VTAIL.n294 VTAIL.n202 4.26717
R597 VTAIL.n266 VTAIL.n217 4.26717
R598 VTAIL.n247 VTAIL.n225 4.26717
R599 VTAIL.n196 VTAIL.n104 4.26717
R600 VTAIL.n168 VTAIL.n119 4.26717
R601 VTAIL.n149 VTAIL.n127 4.26717
R602 VTAIL.n339 VTAIL.n320 3.49141
R603 VTAIL.n360 VTAIL.n308 3.49141
R604 VTAIL.n386 VTAIL.n385 3.49141
R605 VTAIL.n45 VTAIL.n26 3.49141
R606 VTAIL.n66 VTAIL.n14 3.49141
R607 VTAIL.n92 VTAIL.n91 3.49141
R608 VTAIL.n292 VTAIL.n291 3.49141
R609 VTAIL.n267 VTAIL.n215 3.49141
R610 VTAIL.n246 VTAIL.n227 3.49141
R611 VTAIL.n194 VTAIL.n193 3.49141
R612 VTAIL.n169 VTAIL.n117 3.49141
R613 VTAIL.n148 VTAIL.n129 3.49141
R614 VTAIL.n103 VTAIL.n101 3.4574
R615 VTAIL.n197 VTAIL.n103 3.4574
R616 VTAIL.n201 VTAIL.n199 3.4574
R617 VTAIL.n295 VTAIL.n201 3.4574
R618 VTAIL.n99 VTAIL.n97 3.4574
R619 VTAIL.n97 VTAIL.n95 3.4574
R620 VTAIL.n391 VTAIL.n389 3.4574
R621 VTAIL.n336 VTAIL.n335 2.71565
R622 VTAIL.n364 VTAIL.n363 2.71565
R623 VTAIL.n382 VTAIL.n298 2.71565
R624 VTAIL.n42 VTAIL.n41 2.71565
R625 VTAIL.n70 VTAIL.n69 2.71565
R626 VTAIL.n88 VTAIL.n4 2.71565
R627 VTAIL.n288 VTAIL.n204 2.71565
R628 VTAIL.n271 VTAIL.n270 2.71565
R629 VTAIL.n243 VTAIL.n242 2.71565
R630 VTAIL.n190 VTAIL.n106 2.71565
R631 VTAIL.n173 VTAIL.n172 2.71565
R632 VTAIL.n145 VTAIL.n144 2.71565
R633 VTAIL VTAIL.n1 2.65136
R634 VTAIL.n199 VTAIL.n197 2.19878
R635 VTAIL.n95 VTAIL.n1 2.19878
R636 VTAIL.n332 VTAIL.n322 1.93989
R637 VTAIL.n368 VTAIL.n306 1.93989
R638 VTAIL.n381 VTAIL.n300 1.93989
R639 VTAIL.n38 VTAIL.n28 1.93989
R640 VTAIL.n74 VTAIL.n12 1.93989
R641 VTAIL.n87 VTAIL.n6 1.93989
R642 VTAIL.n287 VTAIL.n206 1.93989
R643 VTAIL.n274 VTAIL.n212 1.93989
R644 VTAIL.n239 VTAIL.n229 1.93989
R645 VTAIL.n189 VTAIL.n108 1.93989
R646 VTAIL.n176 VTAIL.n114 1.93989
R647 VTAIL.n141 VTAIL.n131 1.93989
R648 VTAIL.n390 VTAIL.t14 1.17279
R649 VTAIL.n390 VTAIL.t9 1.17279
R650 VTAIL.n0 VTAIL.t13 1.17279
R651 VTAIL.n0 VTAIL.t12 1.17279
R652 VTAIL.n96 VTAIL.t5 1.17279
R653 VTAIL.n96 VTAIL.t6 1.17279
R654 VTAIL.n98 VTAIL.t0 1.17279
R655 VTAIL.n98 VTAIL.t17 1.17279
R656 VTAIL.n200 VTAIL.t3 1.17279
R657 VTAIL.n200 VTAIL.t18 1.17279
R658 VTAIL.n198 VTAIL.t2 1.17279
R659 VTAIL.n198 VTAIL.t4 1.17279
R660 VTAIL.n102 VTAIL.t15 1.17279
R661 VTAIL.n102 VTAIL.t8 1.17279
R662 VTAIL.n100 VTAIL.t11 1.17279
R663 VTAIL.n100 VTAIL.t7 1.17279
R664 VTAIL.n331 VTAIL.n324 1.16414
R665 VTAIL.n369 VTAIL.n304 1.16414
R666 VTAIL.n378 VTAIL.n377 1.16414
R667 VTAIL.n37 VTAIL.n30 1.16414
R668 VTAIL.n75 VTAIL.n10 1.16414
R669 VTAIL.n84 VTAIL.n83 1.16414
R670 VTAIL.n284 VTAIL.n283 1.16414
R671 VTAIL.n275 VTAIL.n210 1.16414
R672 VTAIL.n238 VTAIL.n231 1.16414
R673 VTAIL.n186 VTAIL.n185 1.16414
R674 VTAIL.n177 VTAIL.n112 1.16414
R675 VTAIL.n140 VTAIL.n133 1.16414
R676 VTAIL VTAIL.n391 0.806535
R677 VTAIL.n328 VTAIL.n327 0.388379
R678 VTAIL.n373 VTAIL.n372 0.388379
R679 VTAIL.n374 VTAIL.n302 0.388379
R680 VTAIL.n34 VTAIL.n33 0.388379
R681 VTAIL.n79 VTAIL.n78 0.388379
R682 VTAIL.n80 VTAIL.n8 0.388379
R683 VTAIL.n280 VTAIL.n208 0.388379
R684 VTAIL.n279 VTAIL.n278 0.388379
R685 VTAIL.n235 VTAIL.n234 0.388379
R686 VTAIL.n182 VTAIL.n110 0.388379
R687 VTAIL.n181 VTAIL.n180 0.388379
R688 VTAIL.n137 VTAIL.n136 0.388379
R689 VTAIL.n330 VTAIL.n329 0.155672
R690 VTAIL.n330 VTAIL.n321 0.155672
R691 VTAIL.n337 VTAIL.n321 0.155672
R692 VTAIL.n338 VTAIL.n337 0.155672
R693 VTAIL.n338 VTAIL.n317 0.155672
R694 VTAIL.n345 VTAIL.n317 0.155672
R695 VTAIL.n346 VTAIL.n345 0.155672
R696 VTAIL.n346 VTAIL.n313 0.155672
R697 VTAIL.n353 VTAIL.n313 0.155672
R698 VTAIL.n354 VTAIL.n353 0.155672
R699 VTAIL.n354 VTAIL.n309 0.155672
R700 VTAIL.n361 VTAIL.n309 0.155672
R701 VTAIL.n362 VTAIL.n361 0.155672
R702 VTAIL.n362 VTAIL.n305 0.155672
R703 VTAIL.n370 VTAIL.n305 0.155672
R704 VTAIL.n371 VTAIL.n370 0.155672
R705 VTAIL.n371 VTAIL.n301 0.155672
R706 VTAIL.n379 VTAIL.n301 0.155672
R707 VTAIL.n380 VTAIL.n379 0.155672
R708 VTAIL.n380 VTAIL.n297 0.155672
R709 VTAIL.n387 VTAIL.n297 0.155672
R710 VTAIL.n36 VTAIL.n35 0.155672
R711 VTAIL.n36 VTAIL.n27 0.155672
R712 VTAIL.n43 VTAIL.n27 0.155672
R713 VTAIL.n44 VTAIL.n43 0.155672
R714 VTAIL.n44 VTAIL.n23 0.155672
R715 VTAIL.n51 VTAIL.n23 0.155672
R716 VTAIL.n52 VTAIL.n51 0.155672
R717 VTAIL.n52 VTAIL.n19 0.155672
R718 VTAIL.n59 VTAIL.n19 0.155672
R719 VTAIL.n60 VTAIL.n59 0.155672
R720 VTAIL.n60 VTAIL.n15 0.155672
R721 VTAIL.n67 VTAIL.n15 0.155672
R722 VTAIL.n68 VTAIL.n67 0.155672
R723 VTAIL.n68 VTAIL.n11 0.155672
R724 VTAIL.n76 VTAIL.n11 0.155672
R725 VTAIL.n77 VTAIL.n76 0.155672
R726 VTAIL.n77 VTAIL.n7 0.155672
R727 VTAIL.n85 VTAIL.n7 0.155672
R728 VTAIL.n86 VTAIL.n85 0.155672
R729 VTAIL.n86 VTAIL.n3 0.155672
R730 VTAIL.n93 VTAIL.n3 0.155672
R731 VTAIL.n293 VTAIL.n203 0.155672
R732 VTAIL.n286 VTAIL.n203 0.155672
R733 VTAIL.n286 VTAIL.n285 0.155672
R734 VTAIL.n285 VTAIL.n207 0.155672
R735 VTAIL.n277 VTAIL.n207 0.155672
R736 VTAIL.n277 VTAIL.n276 0.155672
R737 VTAIL.n276 VTAIL.n211 0.155672
R738 VTAIL.n269 VTAIL.n211 0.155672
R739 VTAIL.n269 VTAIL.n268 0.155672
R740 VTAIL.n268 VTAIL.n216 0.155672
R741 VTAIL.n261 VTAIL.n216 0.155672
R742 VTAIL.n261 VTAIL.n260 0.155672
R743 VTAIL.n260 VTAIL.n220 0.155672
R744 VTAIL.n253 VTAIL.n220 0.155672
R745 VTAIL.n253 VTAIL.n252 0.155672
R746 VTAIL.n252 VTAIL.n224 0.155672
R747 VTAIL.n245 VTAIL.n224 0.155672
R748 VTAIL.n245 VTAIL.n244 0.155672
R749 VTAIL.n244 VTAIL.n228 0.155672
R750 VTAIL.n237 VTAIL.n228 0.155672
R751 VTAIL.n237 VTAIL.n236 0.155672
R752 VTAIL.n195 VTAIL.n105 0.155672
R753 VTAIL.n188 VTAIL.n105 0.155672
R754 VTAIL.n188 VTAIL.n187 0.155672
R755 VTAIL.n187 VTAIL.n109 0.155672
R756 VTAIL.n179 VTAIL.n109 0.155672
R757 VTAIL.n179 VTAIL.n178 0.155672
R758 VTAIL.n178 VTAIL.n113 0.155672
R759 VTAIL.n171 VTAIL.n113 0.155672
R760 VTAIL.n171 VTAIL.n170 0.155672
R761 VTAIL.n170 VTAIL.n118 0.155672
R762 VTAIL.n163 VTAIL.n118 0.155672
R763 VTAIL.n163 VTAIL.n162 0.155672
R764 VTAIL.n162 VTAIL.n122 0.155672
R765 VTAIL.n155 VTAIL.n122 0.155672
R766 VTAIL.n155 VTAIL.n154 0.155672
R767 VTAIL.n154 VTAIL.n126 0.155672
R768 VTAIL.n147 VTAIL.n126 0.155672
R769 VTAIL.n147 VTAIL.n146 0.155672
R770 VTAIL.n146 VTAIL.n130 0.155672
R771 VTAIL.n139 VTAIL.n130 0.155672
R772 VTAIL.n139 VTAIL.n138 0.155672
R773 VDD2.n185 VDD2.n97 289.615
R774 VDD2.n88 VDD2.n0 289.615
R775 VDD2.n186 VDD2.n185 185
R776 VDD2.n184 VDD2.n183 185
R777 VDD2.n101 VDD2.n100 185
R778 VDD2.n178 VDD2.n177 185
R779 VDD2.n176 VDD2.n175 185
R780 VDD2.n174 VDD2.n104 185
R781 VDD2.n108 VDD2.n105 185
R782 VDD2.n169 VDD2.n168 185
R783 VDD2.n167 VDD2.n166 185
R784 VDD2.n110 VDD2.n109 185
R785 VDD2.n161 VDD2.n160 185
R786 VDD2.n159 VDD2.n158 185
R787 VDD2.n114 VDD2.n113 185
R788 VDD2.n153 VDD2.n152 185
R789 VDD2.n151 VDD2.n150 185
R790 VDD2.n118 VDD2.n117 185
R791 VDD2.n145 VDD2.n144 185
R792 VDD2.n143 VDD2.n142 185
R793 VDD2.n122 VDD2.n121 185
R794 VDD2.n137 VDD2.n136 185
R795 VDD2.n135 VDD2.n134 185
R796 VDD2.n126 VDD2.n125 185
R797 VDD2.n129 VDD2.n128 185
R798 VDD2.n31 VDD2.n30 185
R799 VDD2.n28 VDD2.n27 185
R800 VDD2.n37 VDD2.n36 185
R801 VDD2.n39 VDD2.n38 185
R802 VDD2.n24 VDD2.n23 185
R803 VDD2.n45 VDD2.n44 185
R804 VDD2.n47 VDD2.n46 185
R805 VDD2.n20 VDD2.n19 185
R806 VDD2.n53 VDD2.n52 185
R807 VDD2.n55 VDD2.n54 185
R808 VDD2.n16 VDD2.n15 185
R809 VDD2.n61 VDD2.n60 185
R810 VDD2.n63 VDD2.n62 185
R811 VDD2.n12 VDD2.n11 185
R812 VDD2.n69 VDD2.n68 185
R813 VDD2.n72 VDD2.n71 185
R814 VDD2.n70 VDD2.n8 185
R815 VDD2.n77 VDD2.n7 185
R816 VDD2.n79 VDD2.n78 185
R817 VDD2.n81 VDD2.n80 185
R818 VDD2.n4 VDD2.n3 185
R819 VDD2.n87 VDD2.n86 185
R820 VDD2.n89 VDD2.n88 185
R821 VDD2.t9 VDD2.n127 147.659
R822 VDD2.t1 VDD2.n29 147.659
R823 VDD2.n185 VDD2.n184 104.615
R824 VDD2.n184 VDD2.n100 104.615
R825 VDD2.n177 VDD2.n100 104.615
R826 VDD2.n177 VDD2.n176 104.615
R827 VDD2.n176 VDD2.n104 104.615
R828 VDD2.n108 VDD2.n104 104.615
R829 VDD2.n168 VDD2.n108 104.615
R830 VDD2.n168 VDD2.n167 104.615
R831 VDD2.n167 VDD2.n109 104.615
R832 VDD2.n160 VDD2.n109 104.615
R833 VDD2.n160 VDD2.n159 104.615
R834 VDD2.n159 VDD2.n113 104.615
R835 VDD2.n152 VDD2.n113 104.615
R836 VDD2.n152 VDD2.n151 104.615
R837 VDD2.n151 VDD2.n117 104.615
R838 VDD2.n144 VDD2.n117 104.615
R839 VDD2.n144 VDD2.n143 104.615
R840 VDD2.n143 VDD2.n121 104.615
R841 VDD2.n136 VDD2.n121 104.615
R842 VDD2.n136 VDD2.n135 104.615
R843 VDD2.n135 VDD2.n125 104.615
R844 VDD2.n128 VDD2.n125 104.615
R845 VDD2.n30 VDD2.n27 104.615
R846 VDD2.n37 VDD2.n27 104.615
R847 VDD2.n38 VDD2.n37 104.615
R848 VDD2.n38 VDD2.n23 104.615
R849 VDD2.n45 VDD2.n23 104.615
R850 VDD2.n46 VDD2.n45 104.615
R851 VDD2.n46 VDD2.n19 104.615
R852 VDD2.n53 VDD2.n19 104.615
R853 VDD2.n54 VDD2.n53 104.615
R854 VDD2.n54 VDD2.n15 104.615
R855 VDD2.n61 VDD2.n15 104.615
R856 VDD2.n62 VDD2.n61 104.615
R857 VDD2.n62 VDD2.n11 104.615
R858 VDD2.n69 VDD2.n11 104.615
R859 VDD2.n71 VDD2.n69 104.615
R860 VDD2.n71 VDD2.n70 104.615
R861 VDD2.n70 VDD2.n7 104.615
R862 VDD2.n79 VDD2.n7 104.615
R863 VDD2.n80 VDD2.n79 104.615
R864 VDD2.n80 VDD2.n3 104.615
R865 VDD2.n87 VDD2.n3 104.615
R866 VDD2.n88 VDD2.n87 104.615
R867 VDD2.n96 VDD2.n95 65.0074
R868 VDD2 VDD2.n193 65.0046
R869 VDD2.n192 VDD2.n191 62.4703
R870 VDD2.n94 VDD2.n93 62.4701
R871 VDD2.n190 VDD2.n96 54.6959
R872 VDD2.n94 VDD2.n92 54.0665
R873 VDD2.n128 VDD2.t9 52.3082
R874 VDD2.n30 VDD2.t1 52.3082
R875 VDD2.n190 VDD2.n189 50.6096
R876 VDD2.n129 VDD2.n127 15.6677
R877 VDD2.n31 VDD2.n29 15.6677
R878 VDD2.n175 VDD2.n174 13.1884
R879 VDD2.n78 VDD2.n77 13.1884
R880 VDD2.n178 VDD2.n103 12.8005
R881 VDD2.n173 VDD2.n105 12.8005
R882 VDD2.n130 VDD2.n126 12.8005
R883 VDD2.n32 VDD2.n28 12.8005
R884 VDD2.n76 VDD2.n8 12.8005
R885 VDD2.n81 VDD2.n6 12.8005
R886 VDD2.n179 VDD2.n101 12.0247
R887 VDD2.n170 VDD2.n169 12.0247
R888 VDD2.n134 VDD2.n133 12.0247
R889 VDD2.n36 VDD2.n35 12.0247
R890 VDD2.n73 VDD2.n72 12.0247
R891 VDD2.n82 VDD2.n4 12.0247
R892 VDD2.n183 VDD2.n182 11.249
R893 VDD2.n166 VDD2.n107 11.249
R894 VDD2.n137 VDD2.n124 11.249
R895 VDD2.n39 VDD2.n26 11.249
R896 VDD2.n68 VDD2.n10 11.249
R897 VDD2.n86 VDD2.n85 11.249
R898 VDD2.n186 VDD2.n99 10.4732
R899 VDD2.n165 VDD2.n110 10.4732
R900 VDD2.n138 VDD2.n122 10.4732
R901 VDD2.n40 VDD2.n24 10.4732
R902 VDD2.n67 VDD2.n12 10.4732
R903 VDD2.n89 VDD2.n2 10.4732
R904 VDD2.n187 VDD2.n97 9.69747
R905 VDD2.n162 VDD2.n161 9.69747
R906 VDD2.n142 VDD2.n141 9.69747
R907 VDD2.n44 VDD2.n43 9.69747
R908 VDD2.n64 VDD2.n63 9.69747
R909 VDD2.n90 VDD2.n0 9.69747
R910 VDD2.n189 VDD2.n188 9.45567
R911 VDD2.n92 VDD2.n91 9.45567
R912 VDD2.n155 VDD2.n154 9.3005
R913 VDD2.n157 VDD2.n156 9.3005
R914 VDD2.n112 VDD2.n111 9.3005
R915 VDD2.n163 VDD2.n162 9.3005
R916 VDD2.n165 VDD2.n164 9.3005
R917 VDD2.n107 VDD2.n106 9.3005
R918 VDD2.n171 VDD2.n170 9.3005
R919 VDD2.n173 VDD2.n172 9.3005
R920 VDD2.n188 VDD2.n187 9.3005
R921 VDD2.n99 VDD2.n98 9.3005
R922 VDD2.n182 VDD2.n181 9.3005
R923 VDD2.n180 VDD2.n179 9.3005
R924 VDD2.n103 VDD2.n102 9.3005
R925 VDD2.n116 VDD2.n115 9.3005
R926 VDD2.n149 VDD2.n148 9.3005
R927 VDD2.n147 VDD2.n146 9.3005
R928 VDD2.n120 VDD2.n119 9.3005
R929 VDD2.n141 VDD2.n140 9.3005
R930 VDD2.n139 VDD2.n138 9.3005
R931 VDD2.n124 VDD2.n123 9.3005
R932 VDD2.n133 VDD2.n132 9.3005
R933 VDD2.n131 VDD2.n130 9.3005
R934 VDD2.n91 VDD2.n90 9.3005
R935 VDD2.n2 VDD2.n1 9.3005
R936 VDD2.n85 VDD2.n84 9.3005
R937 VDD2.n83 VDD2.n82 9.3005
R938 VDD2.n6 VDD2.n5 9.3005
R939 VDD2.n51 VDD2.n50 9.3005
R940 VDD2.n49 VDD2.n48 9.3005
R941 VDD2.n22 VDD2.n21 9.3005
R942 VDD2.n43 VDD2.n42 9.3005
R943 VDD2.n41 VDD2.n40 9.3005
R944 VDD2.n26 VDD2.n25 9.3005
R945 VDD2.n35 VDD2.n34 9.3005
R946 VDD2.n33 VDD2.n32 9.3005
R947 VDD2.n18 VDD2.n17 9.3005
R948 VDD2.n57 VDD2.n56 9.3005
R949 VDD2.n59 VDD2.n58 9.3005
R950 VDD2.n14 VDD2.n13 9.3005
R951 VDD2.n65 VDD2.n64 9.3005
R952 VDD2.n67 VDD2.n66 9.3005
R953 VDD2.n10 VDD2.n9 9.3005
R954 VDD2.n74 VDD2.n73 9.3005
R955 VDD2.n76 VDD2.n75 9.3005
R956 VDD2.n158 VDD2.n112 8.92171
R957 VDD2.n145 VDD2.n120 8.92171
R958 VDD2.n47 VDD2.n22 8.92171
R959 VDD2.n60 VDD2.n14 8.92171
R960 VDD2.n157 VDD2.n114 8.14595
R961 VDD2.n146 VDD2.n118 8.14595
R962 VDD2.n48 VDD2.n20 8.14595
R963 VDD2.n59 VDD2.n16 8.14595
R964 VDD2.n154 VDD2.n153 7.3702
R965 VDD2.n150 VDD2.n149 7.3702
R966 VDD2.n52 VDD2.n51 7.3702
R967 VDD2.n56 VDD2.n55 7.3702
R968 VDD2.n153 VDD2.n116 6.59444
R969 VDD2.n150 VDD2.n116 6.59444
R970 VDD2.n52 VDD2.n18 6.59444
R971 VDD2.n55 VDD2.n18 6.59444
R972 VDD2.n154 VDD2.n114 5.81868
R973 VDD2.n149 VDD2.n118 5.81868
R974 VDD2.n51 VDD2.n20 5.81868
R975 VDD2.n56 VDD2.n16 5.81868
R976 VDD2.n158 VDD2.n157 5.04292
R977 VDD2.n146 VDD2.n145 5.04292
R978 VDD2.n48 VDD2.n47 5.04292
R979 VDD2.n60 VDD2.n59 5.04292
R980 VDD2.n131 VDD2.n127 4.38563
R981 VDD2.n33 VDD2.n29 4.38563
R982 VDD2.n189 VDD2.n97 4.26717
R983 VDD2.n161 VDD2.n112 4.26717
R984 VDD2.n142 VDD2.n120 4.26717
R985 VDD2.n44 VDD2.n22 4.26717
R986 VDD2.n63 VDD2.n14 4.26717
R987 VDD2.n92 VDD2.n0 4.26717
R988 VDD2.n187 VDD2.n186 3.49141
R989 VDD2.n162 VDD2.n110 3.49141
R990 VDD2.n141 VDD2.n122 3.49141
R991 VDD2.n43 VDD2.n24 3.49141
R992 VDD2.n64 VDD2.n12 3.49141
R993 VDD2.n90 VDD2.n89 3.49141
R994 VDD2.n192 VDD2.n190 3.4574
R995 VDD2.n183 VDD2.n99 2.71565
R996 VDD2.n166 VDD2.n165 2.71565
R997 VDD2.n138 VDD2.n137 2.71565
R998 VDD2.n40 VDD2.n39 2.71565
R999 VDD2.n68 VDD2.n67 2.71565
R1000 VDD2.n86 VDD2.n2 2.71565
R1001 VDD2.n182 VDD2.n101 1.93989
R1002 VDD2.n169 VDD2.n107 1.93989
R1003 VDD2.n134 VDD2.n124 1.93989
R1004 VDD2.n36 VDD2.n26 1.93989
R1005 VDD2.n72 VDD2.n10 1.93989
R1006 VDD2.n85 VDD2.n4 1.93989
R1007 VDD2.n193 VDD2.t5 1.17279
R1008 VDD2.n193 VDD2.t4 1.17279
R1009 VDD2.n191 VDD2.t8 1.17279
R1010 VDD2.n191 VDD2.t3 1.17279
R1011 VDD2.n95 VDD2.t7 1.17279
R1012 VDD2.n95 VDD2.t0 1.17279
R1013 VDD2.n93 VDD2.t6 1.17279
R1014 VDD2.n93 VDD2.t2 1.17279
R1015 VDD2.n179 VDD2.n178 1.16414
R1016 VDD2.n170 VDD2.n105 1.16414
R1017 VDD2.n133 VDD2.n126 1.16414
R1018 VDD2.n35 VDD2.n28 1.16414
R1019 VDD2.n73 VDD2.n8 1.16414
R1020 VDD2.n82 VDD2.n81 1.16414
R1021 VDD2 VDD2.n192 0.922914
R1022 VDD2.n96 VDD2.n94 0.809378
R1023 VDD2.n175 VDD2.n103 0.388379
R1024 VDD2.n174 VDD2.n173 0.388379
R1025 VDD2.n130 VDD2.n129 0.388379
R1026 VDD2.n32 VDD2.n31 0.388379
R1027 VDD2.n77 VDD2.n76 0.388379
R1028 VDD2.n78 VDD2.n6 0.388379
R1029 VDD2.n188 VDD2.n98 0.155672
R1030 VDD2.n181 VDD2.n98 0.155672
R1031 VDD2.n181 VDD2.n180 0.155672
R1032 VDD2.n180 VDD2.n102 0.155672
R1033 VDD2.n172 VDD2.n102 0.155672
R1034 VDD2.n172 VDD2.n171 0.155672
R1035 VDD2.n171 VDD2.n106 0.155672
R1036 VDD2.n164 VDD2.n106 0.155672
R1037 VDD2.n164 VDD2.n163 0.155672
R1038 VDD2.n163 VDD2.n111 0.155672
R1039 VDD2.n156 VDD2.n111 0.155672
R1040 VDD2.n156 VDD2.n155 0.155672
R1041 VDD2.n155 VDD2.n115 0.155672
R1042 VDD2.n148 VDD2.n115 0.155672
R1043 VDD2.n148 VDD2.n147 0.155672
R1044 VDD2.n147 VDD2.n119 0.155672
R1045 VDD2.n140 VDD2.n119 0.155672
R1046 VDD2.n140 VDD2.n139 0.155672
R1047 VDD2.n139 VDD2.n123 0.155672
R1048 VDD2.n132 VDD2.n123 0.155672
R1049 VDD2.n132 VDD2.n131 0.155672
R1050 VDD2.n34 VDD2.n33 0.155672
R1051 VDD2.n34 VDD2.n25 0.155672
R1052 VDD2.n41 VDD2.n25 0.155672
R1053 VDD2.n42 VDD2.n41 0.155672
R1054 VDD2.n42 VDD2.n21 0.155672
R1055 VDD2.n49 VDD2.n21 0.155672
R1056 VDD2.n50 VDD2.n49 0.155672
R1057 VDD2.n50 VDD2.n17 0.155672
R1058 VDD2.n57 VDD2.n17 0.155672
R1059 VDD2.n58 VDD2.n57 0.155672
R1060 VDD2.n58 VDD2.n13 0.155672
R1061 VDD2.n65 VDD2.n13 0.155672
R1062 VDD2.n66 VDD2.n65 0.155672
R1063 VDD2.n66 VDD2.n9 0.155672
R1064 VDD2.n74 VDD2.n9 0.155672
R1065 VDD2.n75 VDD2.n74 0.155672
R1066 VDD2.n75 VDD2.n5 0.155672
R1067 VDD2.n83 VDD2.n5 0.155672
R1068 VDD2.n84 VDD2.n83 0.155672
R1069 VDD2.n84 VDD2.n1 0.155672
R1070 VDD2.n91 VDD2.n1 0.155672
R1071 B.n1252 B.n1251 585
R1072 B.n448 B.n204 585
R1073 B.n447 B.n446 585
R1074 B.n445 B.n444 585
R1075 B.n443 B.n442 585
R1076 B.n441 B.n440 585
R1077 B.n439 B.n438 585
R1078 B.n437 B.n436 585
R1079 B.n435 B.n434 585
R1080 B.n433 B.n432 585
R1081 B.n431 B.n430 585
R1082 B.n429 B.n428 585
R1083 B.n427 B.n426 585
R1084 B.n425 B.n424 585
R1085 B.n423 B.n422 585
R1086 B.n421 B.n420 585
R1087 B.n419 B.n418 585
R1088 B.n417 B.n416 585
R1089 B.n415 B.n414 585
R1090 B.n413 B.n412 585
R1091 B.n411 B.n410 585
R1092 B.n409 B.n408 585
R1093 B.n407 B.n406 585
R1094 B.n405 B.n404 585
R1095 B.n403 B.n402 585
R1096 B.n401 B.n400 585
R1097 B.n399 B.n398 585
R1098 B.n397 B.n396 585
R1099 B.n395 B.n394 585
R1100 B.n393 B.n392 585
R1101 B.n391 B.n390 585
R1102 B.n389 B.n388 585
R1103 B.n387 B.n386 585
R1104 B.n385 B.n384 585
R1105 B.n383 B.n382 585
R1106 B.n381 B.n380 585
R1107 B.n379 B.n378 585
R1108 B.n377 B.n376 585
R1109 B.n375 B.n374 585
R1110 B.n373 B.n372 585
R1111 B.n371 B.n370 585
R1112 B.n369 B.n368 585
R1113 B.n367 B.n366 585
R1114 B.n365 B.n364 585
R1115 B.n363 B.n362 585
R1116 B.n361 B.n360 585
R1117 B.n359 B.n358 585
R1118 B.n357 B.n356 585
R1119 B.n355 B.n354 585
R1120 B.n353 B.n352 585
R1121 B.n351 B.n350 585
R1122 B.n349 B.n348 585
R1123 B.n347 B.n346 585
R1124 B.n345 B.n344 585
R1125 B.n343 B.n342 585
R1126 B.n341 B.n340 585
R1127 B.n339 B.n338 585
R1128 B.n337 B.n336 585
R1129 B.n335 B.n334 585
R1130 B.n333 B.n332 585
R1131 B.n331 B.n330 585
R1132 B.n329 B.n328 585
R1133 B.n327 B.n326 585
R1134 B.n325 B.n324 585
R1135 B.n323 B.n322 585
R1136 B.n321 B.n320 585
R1137 B.n319 B.n318 585
R1138 B.n317 B.n316 585
R1139 B.n315 B.n314 585
R1140 B.n313 B.n312 585
R1141 B.n311 B.n310 585
R1142 B.n309 B.n308 585
R1143 B.n307 B.n306 585
R1144 B.n305 B.n304 585
R1145 B.n303 B.n302 585
R1146 B.n301 B.n300 585
R1147 B.n299 B.n298 585
R1148 B.n297 B.n296 585
R1149 B.n295 B.n294 585
R1150 B.n293 B.n292 585
R1151 B.n291 B.n290 585
R1152 B.n289 B.n288 585
R1153 B.n287 B.n286 585
R1154 B.n285 B.n284 585
R1155 B.n283 B.n282 585
R1156 B.n281 B.n280 585
R1157 B.n279 B.n278 585
R1158 B.n277 B.n276 585
R1159 B.n275 B.n274 585
R1160 B.n273 B.n272 585
R1161 B.n271 B.n270 585
R1162 B.n269 B.n268 585
R1163 B.n267 B.n266 585
R1164 B.n265 B.n264 585
R1165 B.n263 B.n262 585
R1166 B.n261 B.n260 585
R1167 B.n259 B.n258 585
R1168 B.n257 B.n256 585
R1169 B.n255 B.n254 585
R1170 B.n253 B.n252 585
R1171 B.n251 B.n250 585
R1172 B.n249 B.n248 585
R1173 B.n247 B.n246 585
R1174 B.n245 B.n244 585
R1175 B.n243 B.n242 585
R1176 B.n241 B.n240 585
R1177 B.n239 B.n238 585
R1178 B.n237 B.n236 585
R1179 B.n235 B.n234 585
R1180 B.n233 B.n232 585
R1181 B.n231 B.n230 585
R1182 B.n229 B.n228 585
R1183 B.n227 B.n226 585
R1184 B.n225 B.n224 585
R1185 B.n223 B.n222 585
R1186 B.n221 B.n220 585
R1187 B.n219 B.n218 585
R1188 B.n217 B.n216 585
R1189 B.n215 B.n214 585
R1190 B.n213 B.n212 585
R1191 B.n144 B.n143 585
R1192 B.n1257 B.n1256 585
R1193 B.n1250 B.n205 585
R1194 B.n205 B.n141 585
R1195 B.n1249 B.n140 585
R1196 B.n1261 B.n140 585
R1197 B.n1248 B.n139 585
R1198 B.n1262 B.n139 585
R1199 B.n1247 B.n138 585
R1200 B.n1263 B.n138 585
R1201 B.n1246 B.n1245 585
R1202 B.n1245 B.n134 585
R1203 B.n1244 B.n133 585
R1204 B.n1269 B.n133 585
R1205 B.n1243 B.n132 585
R1206 B.n1270 B.n132 585
R1207 B.n1242 B.n131 585
R1208 B.n1271 B.n131 585
R1209 B.n1241 B.n1240 585
R1210 B.n1240 B.n127 585
R1211 B.n1239 B.n126 585
R1212 B.n1277 B.n126 585
R1213 B.n1238 B.n125 585
R1214 B.n1278 B.n125 585
R1215 B.n1237 B.n124 585
R1216 B.n1279 B.n124 585
R1217 B.n1236 B.n1235 585
R1218 B.n1235 B.n120 585
R1219 B.n1234 B.n119 585
R1220 B.n1285 B.n119 585
R1221 B.n1233 B.n118 585
R1222 B.n1286 B.n118 585
R1223 B.n1232 B.n117 585
R1224 B.n1287 B.n117 585
R1225 B.n1231 B.n1230 585
R1226 B.n1230 B.n113 585
R1227 B.n1229 B.n112 585
R1228 B.n1293 B.n112 585
R1229 B.n1228 B.n111 585
R1230 B.n1294 B.n111 585
R1231 B.n1227 B.n110 585
R1232 B.n1295 B.n110 585
R1233 B.n1226 B.n1225 585
R1234 B.n1225 B.n106 585
R1235 B.n1224 B.n105 585
R1236 B.n1301 B.n105 585
R1237 B.n1223 B.n104 585
R1238 B.n1302 B.n104 585
R1239 B.n1222 B.n103 585
R1240 B.n1303 B.n103 585
R1241 B.n1221 B.n1220 585
R1242 B.n1220 B.n102 585
R1243 B.n1219 B.n98 585
R1244 B.n1309 B.n98 585
R1245 B.n1218 B.n97 585
R1246 B.n1310 B.n97 585
R1247 B.n1217 B.n96 585
R1248 B.n1311 B.n96 585
R1249 B.n1216 B.n1215 585
R1250 B.n1215 B.n92 585
R1251 B.n1214 B.n91 585
R1252 B.n1317 B.n91 585
R1253 B.n1213 B.n90 585
R1254 B.n1318 B.n90 585
R1255 B.n1212 B.n89 585
R1256 B.n1319 B.n89 585
R1257 B.n1211 B.n1210 585
R1258 B.n1210 B.n85 585
R1259 B.n1209 B.n84 585
R1260 B.n1325 B.n84 585
R1261 B.n1208 B.n83 585
R1262 B.n1326 B.n83 585
R1263 B.n1207 B.n82 585
R1264 B.n1327 B.n82 585
R1265 B.n1206 B.n1205 585
R1266 B.n1205 B.n81 585
R1267 B.n1204 B.n77 585
R1268 B.n1333 B.n77 585
R1269 B.n1203 B.n76 585
R1270 B.n1334 B.n76 585
R1271 B.n1202 B.n75 585
R1272 B.n1335 B.n75 585
R1273 B.n1201 B.n1200 585
R1274 B.n1200 B.n71 585
R1275 B.n1199 B.n70 585
R1276 B.n1341 B.n70 585
R1277 B.n1198 B.n69 585
R1278 B.n1342 B.n69 585
R1279 B.n1197 B.n68 585
R1280 B.n1343 B.n68 585
R1281 B.n1196 B.n1195 585
R1282 B.n1195 B.n64 585
R1283 B.n1194 B.n63 585
R1284 B.n1349 B.n63 585
R1285 B.n1193 B.n62 585
R1286 B.n1350 B.n62 585
R1287 B.n1192 B.n61 585
R1288 B.n1351 B.n61 585
R1289 B.n1191 B.n1190 585
R1290 B.n1190 B.n57 585
R1291 B.n1189 B.n56 585
R1292 B.n1357 B.n56 585
R1293 B.n1188 B.n55 585
R1294 B.n1358 B.n55 585
R1295 B.n1187 B.n54 585
R1296 B.n1359 B.n54 585
R1297 B.n1186 B.n1185 585
R1298 B.n1185 B.n50 585
R1299 B.n1184 B.n49 585
R1300 B.n1365 B.n49 585
R1301 B.n1183 B.n48 585
R1302 B.n1366 B.n48 585
R1303 B.n1182 B.n47 585
R1304 B.n1367 B.n47 585
R1305 B.n1181 B.n1180 585
R1306 B.n1180 B.n43 585
R1307 B.n1179 B.n42 585
R1308 B.n1373 B.n42 585
R1309 B.n1178 B.n41 585
R1310 B.n1374 B.n41 585
R1311 B.n1177 B.n40 585
R1312 B.n1375 B.n40 585
R1313 B.n1176 B.n1175 585
R1314 B.n1175 B.n36 585
R1315 B.n1174 B.n35 585
R1316 B.n1381 B.n35 585
R1317 B.n1173 B.n34 585
R1318 B.n1382 B.n34 585
R1319 B.n1172 B.n33 585
R1320 B.n1383 B.n33 585
R1321 B.n1171 B.n1170 585
R1322 B.n1170 B.n29 585
R1323 B.n1169 B.n28 585
R1324 B.n1389 B.n28 585
R1325 B.n1168 B.n27 585
R1326 B.n1390 B.n27 585
R1327 B.n1167 B.n26 585
R1328 B.n1391 B.n26 585
R1329 B.n1166 B.n1165 585
R1330 B.n1165 B.n22 585
R1331 B.n1164 B.n21 585
R1332 B.n1397 B.n21 585
R1333 B.n1163 B.n20 585
R1334 B.n1398 B.n20 585
R1335 B.n1162 B.n19 585
R1336 B.n1399 B.n19 585
R1337 B.n1161 B.n1160 585
R1338 B.n1160 B.n15 585
R1339 B.n1159 B.n14 585
R1340 B.n1405 B.n14 585
R1341 B.n1158 B.n13 585
R1342 B.n1406 B.n13 585
R1343 B.n1157 B.n12 585
R1344 B.n1407 B.n12 585
R1345 B.n1156 B.n1155 585
R1346 B.n1155 B.n8 585
R1347 B.n1154 B.n7 585
R1348 B.n1413 B.n7 585
R1349 B.n1153 B.n6 585
R1350 B.n1414 B.n6 585
R1351 B.n1152 B.n5 585
R1352 B.n1415 B.n5 585
R1353 B.n1151 B.n1150 585
R1354 B.n1150 B.n4 585
R1355 B.n1149 B.n449 585
R1356 B.n1149 B.n1148 585
R1357 B.n1139 B.n450 585
R1358 B.n451 B.n450 585
R1359 B.n1141 B.n1140 585
R1360 B.n1142 B.n1141 585
R1361 B.n1138 B.n456 585
R1362 B.n456 B.n455 585
R1363 B.n1137 B.n1136 585
R1364 B.n1136 B.n1135 585
R1365 B.n458 B.n457 585
R1366 B.n459 B.n458 585
R1367 B.n1128 B.n1127 585
R1368 B.n1129 B.n1128 585
R1369 B.n1126 B.n464 585
R1370 B.n464 B.n463 585
R1371 B.n1125 B.n1124 585
R1372 B.n1124 B.n1123 585
R1373 B.n466 B.n465 585
R1374 B.n467 B.n466 585
R1375 B.n1116 B.n1115 585
R1376 B.n1117 B.n1116 585
R1377 B.n1114 B.n472 585
R1378 B.n472 B.n471 585
R1379 B.n1113 B.n1112 585
R1380 B.n1112 B.n1111 585
R1381 B.n474 B.n473 585
R1382 B.n475 B.n474 585
R1383 B.n1104 B.n1103 585
R1384 B.n1105 B.n1104 585
R1385 B.n1102 B.n480 585
R1386 B.n480 B.n479 585
R1387 B.n1101 B.n1100 585
R1388 B.n1100 B.n1099 585
R1389 B.n482 B.n481 585
R1390 B.n483 B.n482 585
R1391 B.n1092 B.n1091 585
R1392 B.n1093 B.n1092 585
R1393 B.n1090 B.n488 585
R1394 B.n488 B.n487 585
R1395 B.n1089 B.n1088 585
R1396 B.n1088 B.n1087 585
R1397 B.n490 B.n489 585
R1398 B.n491 B.n490 585
R1399 B.n1080 B.n1079 585
R1400 B.n1081 B.n1080 585
R1401 B.n1078 B.n496 585
R1402 B.n496 B.n495 585
R1403 B.n1077 B.n1076 585
R1404 B.n1076 B.n1075 585
R1405 B.n498 B.n497 585
R1406 B.n499 B.n498 585
R1407 B.n1068 B.n1067 585
R1408 B.n1069 B.n1068 585
R1409 B.n1066 B.n504 585
R1410 B.n504 B.n503 585
R1411 B.n1065 B.n1064 585
R1412 B.n1064 B.n1063 585
R1413 B.n506 B.n505 585
R1414 B.n507 B.n506 585
R1415 B.n1056 B.n1055 585
R1416 B.n1057 B.n1056 585
R1417 B.n1054 B.n512 585
R1418 B.n512 B.n511 585
R1419 B.n1053 B.n1052 585
R1420 B.n1052 B.n1051 585
R1421 B.n514 B.n513 585
R1422 B.n515 B.n514 585
R1423 B.n1044 B.n1043 585
R1424 B.n1045 B.n1044 585
R1425 B.n1042 B.n520 585
R1426 B.n520 B.n519 585
R1427 B.n1041 B.n1040 585
R1428 B.n1040 B.n1039 585
R1429 B.n522 B.n521 585
R1430 B.n523 B.n522 585
R1431 B.n1032 B.n1031 585
R1432 B.n1033 B.n1032 585
R1433 B.n1030 B.n528 585
R1434 B.n528 B.n527 585
R1435 B.n1029 B.n1028 585
R1436 B.n1028 B.n1027 585
R1437 B.n530 B.n529 585
R1438 B.n1020 B.n530 585
R1439 B.n1019 B.n1018 585
R1440 B.n1021 B.n1019 585
R1441 B.n1017 B.n535 585
R1442 B.n535 B.n534 585
R1443 B.n1016 B.n1015 585
R1444 B.n1015 B.n1014 585
R1445 B.n537 B.n536 585
R1446 B.n538 B.n537 585
R1447 B.n1007 B.n1006 585
R1448 B.n1008 B.n1007 585
R1449 B.n1005 B.n543 585
R1450 B.n543 B.n542 585
R1451 B.n1004 B.n1003 585
R1452 B.n1003 B.n1002 585
R1453 B.n545 B.n544 585
R1454 B.n546 B.n545 585
R1455 B.n995 B.n994 585
R1456 B.n996 B.n995 585
R1457 B.n993 B.n551 585
R1458 B.n551 B.n550 585
R1459 B.n992 B.n991 585
R1460 B.n991 B.n990 585
R1461 B.n553 B.n552 585
R1462 B.n983 B.n553 585
R1463 B.n982 B.n981 585
R1464 B.n984 B.n982 585
R1465 B.n980 B.n558 585
R1466 B.n558 B.n557 585
R1467 B.n979 B.n978 585
R1468 B.n978 B.n977 585
R1469 B.n560 B.n559 585
R1470 B.n561 B.n560 585
R1471 B.n970 B.n969 585
R1472 B.n971 B.n970 585
R1473 B.n968 B.n566 585
R1474 B.n566 B.n565 585
R1475 B.n967 B.n966 585
R1476 B.n966 B.n965 585
R1477 B.n568 B.n567 585
R1478 B.n569 B.n568 585
R1479 B.n958 B.n957 585
R1480 B.n959 B.n958 585
R1481 B.n956 B.n574 585
R1482 B.n574 B.n573 585
R1483 B.n955 B.n954 585
R1484 B.n954 B.n953 585
R1485 B.n576 B.n575 585
R1486 B.n577 B.n576 585
R1487 B.n946 B.n945 585
R1488 B.n947 B.n946 585
R1489 B.n944 B.n582 585
R1490 B.n582 B.n581 585
R1491 B.n943 B.n942 585
R1492 B.n942 B.n941 585
R1493 B.n584 B.n583 585
R1494 B.n585 B.n584 585
R1495 B.n934 B.n933 585
R1496 B.n935 B.n934 585
R1497 B.n932 B.n590 585
R1498 B.n590 B.n589 585
R1499 B.n931 B.n930 585
R1500 B.n930 B.n929 585
R1501 B.n592 B.n591 585
R1502 B.n593 B.n592 585
R1503 B.n922 B.n921 585
R1504 B.n923 B.n922 585
R1505 B.n920 B.n598 585
R1506 B.n598 B.n597 585
R1507 B.n919 B.n918 585
R1508 B.n918 B.n917 585
R1509 B.n600 B.n599 585
R1510 B.n601 B.n600 585
R1511 B.n913 B.n912 585
R1512 B.n604 B.n603 585
R1513 B.n909 B.n908 585
R1514 B.n910 B.n909 585
R1515 B.n907 B.n665 585
R1516 B.n906 B.n905 585
R1517 B.n904 B.n903 585
R1518 B.n902 B.n901 585
R1519 B.n900 B.n899 585
R1520 B.n898 B.n897 585
R1521 B.n896 B.n895 585
R1522 B.n894 B.n893 585
R1523 B.n892 B.n891 585
R1524 B.n890 B.n889 585
R1525 B.n888 B.n887 585
R1526 B.n886 B.n885 585
R1527 B.n884 B.n883 585
R1528 B.n882 B.n881 585
R1529 B.n880 B.n879 585
R1530 B.n878 B.n877 585
R1531 B.n876 B.n875 585
R1532 B.n874 B.n873 585
R1533 B.n872 B.n871 585
R1534 B.n870 B.n869 585
R1535 B.n868 B.n867 585
R1536 B.n866 B.n865 585
R1537 B.n864 B.n863 585
R1538 B.n862 B.n861 585
R1539 B.n860 B.n859 585
R1540 B.n858 B.n857 585
R1541 B.n856 B.n855 585
R1542 B.n854 B.n853 585
R1543 B.n852 B.n851 585
R1544 B.n850 B.n849 585
R1545 B.n848 B.n847 585
R1546 B.n846 B.n845 585
R1547 B.n844 B.n843 585
R1548 B.n842 B.n841 585
R1549 B.n840 B.n839 585
R1550 B.n838 B.n837 585
R1551 B.n836 B.n835 585
R1552 B.n834 B.n833 585
R1553 B.n832 B.n831 585
R1554 B.n830 B.n829 585
R1555 B.n828 B.n827 585
R1556 B.n826 B.n825 585
R1557 B.n824 B.n823 585
R1558 B.n822 B.n821 585
R1559 B.n820 B.n819 585
R1560 B.n818 B.n817 585
R1561 B.n816 B.n815 585
R1562 B.n814 B.n813 585
R1563 B.n812 B.n811 585
R1564 B.n810 B.n809 585
R1565 B.n808 B.n807 585
R1566 B.n806 B.n805 585
R1567 B.n804 B.n803 585
R1568 B.n801 B.n800 585
R1569 B.n799 B.n798 585
R1570 B.n797 B.n796 585
R1571 B.n795 B.n794 585
R1572 B.n793 B.n792 585
R1573 B.n791 B.n790 585
R1574 B.n789 B.n788 585
R1575 B.n787 B.n786 585
R1576 B.n785 B.n784 585
R1577 B.n783 B.n782 585
R1578 B.n780 B.n779 585
R1579 B.n778 B.n777 585
R1580 B.n776 B.n775 585
R1581 B.n774 B.n773 585
R1582 B.n772 B.n771 585
R1583 B.n770 B.n769 585
R1584 B.n768 B.n767 585
R1585 B.n766 B.n765 585
R1586 B.n764 B.n763 585
R1587 B.n762 B.n761 585
R1588 B.n760 B.n759 585
R1589 B.n758 B.n757 585
R1590 B.n756 B.n755 585
R1591 B.n754 B.n753 585
R1592 B.n752 B.n751 585
R1593 B.n750 B.n749 585
R1594 B.n748 B.n747 585
R1595 B.n746 B.n745 585
R1596 B.n744 B.n743 585
R1597 B.n742 B.n741 585
R1598 B.n740 B.n739 585
R1599 B.n738 B.n737 585
R1600 B.n736 B.n735 585
R1601 B.n734 B.n733 585
R1602 B.n732 B.n731 585
R1603 B.n730 B.n729 585
R1604 B.n728 B.n727 585
R1605 B.n726 B.n725 585
R1606 B.n724 B.n723 585
R1607 B.n722 B.n721 585
R1608 B.n720 B.n719 585
R1609 B.n718 B.n717 585
R1610 B.n716 B.n715 585
R1611 B.n714 B.n713 585
R1612 B.n712 B.n711 585
R1613 B.n710 B.n709 585
R1614 B.n708 B.n707 585
R1615 B.n706 B.n705 585
R1616 B.n704 B.n703 585
R1617 B.n702 B.n701 585
R1618 B.n700 B.n699 585
R1619 B.n698 B.n697 585
R1620 B.n696 B.n695 585
R1621 B.n694 B.n693 585
R1622 B.n692 B.n691 585
R1623 B.n690 B.n689 585
R1624 B.n688 B.n687 585
R1625 B.n686 B.n685 585
R1626 B.n684 B.n683 585
R1627 B.n682 B.n681 585
R1628 B.n680 B.n679 585
R1629 B.n678 B.n677 585
R1630 B.n676 B.n675 585
R1631 B.n674 B.n673 585
R1632 B.n672 B.n671 585
R1633 B.n670 B.n664 585
R1634 B.n910 B.n664 585
R1635 B.n914 B.n602 585
R1636 B.n602 B.n601 585
R1637 B.n916 B.n915 585
R1638 B.n917 B.n916 585
R1639 B.n596 B.n595 585
R1640 B.n597 B.n596 585
R1641 B.n925 B.n924 585
R1642 B.n924 B.n923 585
R1643 B.n926 B.n594 585
R1644 B.n594 B.n593 585
R1645 B.n928 B.n927 585
R1646 B.n929 B.n928 585
R1647 B.n588 B.n587 585
R1648 B.n589 B.n588 585
R1649 B.n937 B.n936 585
R1650 B.n936 B.n935 585
R1651 B.n938 B.n586 585
R1652 B.n586 B.n585 585
R1653 B.n940 B.n939 585
R1654 B.n941 B.n940 585
R1655 B.n580 B.n579 585
R1656 B.n581 B.n580 585
R1657 B.n949 B.n948 585
R1658 B.n948 B.n947 585
R1659 B.n950 B.n578 585
R1660 B.n578 B.n577 585
R1661 B.n952 B.n951 585
R1662 B.n953 B.n952 585
R1663 B.n572 B.n571 585
R1664 B.n573 B.n572 585
R1665 B.n961 B.n960 585
R1666 B.n960 B.n959 585
R1667 B.n962 B.n570 585
R1668 B.n570 B.n569 585
R1669 B.n964 B.n963 585
R1670 B.n965 B.n964 585
R1671 B.n564 B.n563 585
R1672 B.n565 B.n564 585
R1673 B.n973 B.n972 585
R1674 B.n972 B.n971 585
R1675 B.n974 B.n562 585
R1676 B.n562 B.n561 585
R1677 B.n976 B.n975 585
R1678 B.n977 B.n976 585
R1679 B.n556 B.n555 585
R1680 B.n557 B.n556 585
R1681 B.n986 B.n985 585
R1682 B.n985 B.n984 585
R1683 B.n987 B.n554 585
R1684 B.n983 B.n554 585
R1685 B.n989 B.n988 585
R1686 B.n990 B.n989 585
R1687 B.n549 B.n548 585
R1688 B.n550 B.n549 585
R1689 B.n998 B.n997 585
R1690 B.n997 B.n996 585
R1691 B.n999 B.n547 585
R1692 B.n547 B.n546 585
R1693 B.n1001 B.n1000 585
R1694 B.n1002 B.n1001 585
R1695 B.n541 B.n540 585
R1696 B.n542 B.n541 585
R1697 B.n1010 B.n1009 585
R1698 B.n1009 B.n1008 585
R1699 B.n1011 B.n539 585
R1700 B.n539 B.n538 585
R1701 B.n1013 B.n1012 585
R1702 B.n1014 B.n1013 585
R1703 B.n533 B.n532 585
R1704 B.n534 B.n533 585
R1705 B.n1023 B.n1022 585
R1706 B.n1022 B.n1021 585
R1707 B.n1024 B.n531 585
R1708 B.n1020 B.n531 585
R1709 B.n1026 B.n1025 585
R1710 B.n1027 B.n1026 585
R1711 B.n526 B.n525 585
R1712 B.n527 B.n526 585
R1713 B.n1035 B.n1034 585
R1714 B.n1034 B.n1033 585
R1715 B.n1036 B.n524 585
R1716 B.n524 B.n523 585
R1717 B.n1038 B.n1037 585
R1718 B.n1039 B.n1038 585
R1719 B.n518 B.n517 585
R1720 B.n519 B.n518 585
R1721 B.n1047 B.n1046 585
R1722 B.n1046 B.n1045 585
R1723 B.n1048 B.n516 585
R1724 B.n516 B.n515 585
R1725 B.n1050 B.n1049 585
R1726 B.n1051 B.n1050 585
R1727 B.n510 B.n509 585
R1728 B.n511 B.n510 585
R1729 B.n1059 B.n1058 585
R1730 B.n1058 B.n1057 585
R1731 B.n1060 B.n508 585
R1732 B.n508 B.n507 585
R1733 B.n1062 B.n1061 585
R1734 B.n1063 B.n1062 585
R1735 B.n502 B.n501 585
R1736 B.n503 B.n502 585
R1737 B.n1071 B.n1070 585
R1738 B.n1070 B.n1069 585
R1739 B.n1072 B.n500 585
R1740 B.n500 B.n499 585
R1741 B.n1074 B.n1073 585
R1742 B.n1075 B.n1074 585
R1743 B.n494 B.n493 585
R1744 B.n495 B.n494 585
R1745 B.n1083 B.n1082 585
R1746 B.n1082 B.n1081 585
R1747 B.n1084 B.n492 585
R1748 B.n492 B.n491 585
R1749 B.n1086 B.n1085 585
R1750 B.n1087 B.n1086 585
R1751 B.n486 B.n485 585
R1752 B.n487 B.n486 585
R1753 B.n1095 B.n1094 585
R1754 B.n1094 B.n1093 585
R1755 B.n1096 B.n484 585
R1756 B.n484 B.n483 585
R1757 B.n1098 B.n1097 585
R1758 B.n1099 B.n1098 585
R1759 B.n478 B.n477 585
R1760 B.n479 B.n478 585
R1761 B.n1107 B.n1106 585
R1762 B.n1106 B.n1105 585
R1763 B.n1108 B.n476 585
R1764 B.n476 B.n475 585
R1765 B.n1110 B.n1109 585
R1766 B.n1111 B.n1110 585
R1767 B.n470 B.n469 585
R1768 B.n471 B.n470 585
R1769 B.n1119 B.n1118 585
R1770 B.n1118 B.n1117 585
R1771 B.n1120 B.n468 585
R1772 B.n468 B.n467 585
R1773 B.n1122 B.n1121 585
R1774 B.n1123 B.n1122 585
R1775 B.n462 B.n461 585
R1776 B.n463 B.n462 585
R1777 B.n1131 B.n1130 585
R1778 B.n1130 B.n1129 585
R1779 B.n1132 B.n460 585
R1780 B.n460 B.n459 585
R1781 B.n1134 B.n1133 585
R1782 B.n1135 B.n1134 585
R1783 B.n454 B.n453 585
R1784 B.n455 B.n454 585
R1785 B.n1144 B.n1143 585
R1786 B.n1143 B.n1142 585
R1787 B.n1145 B.n452 585
R1788 B.n452 B.n451 585
R1789 B.n1147 B.n1146 585
R1790 B.n1148 B.n1147 585
R1791 B.n2 B.n0 585
R1792 B.n4 B.n2 585
R1793 B.n3 B.n1 585
R1794 B.n1414 B.n3 585
R1795 B.n1412 B.n1411 585
R1796 B.n1413 B.n1412 585
R1797 B.n1410 B.n9 585
R1798 B.n9 B.n8 585
R1799 B.n1409 B.n1408 585
R1800 B.n1408 B.n1407 585
R1801 B.n11 B.n10 585
R1802 B.n1406 B.n11 585
R1803 B.n1404 B.n1403 585
R1804 B.n1405 B.n1404 585
R1805 B.n1402 B.n16 585
R1806 B.n16 B.n15 585
R1807 B.n1401 B.n1400 585
R1808 B.n1400 B.n1399 585
R1809 B.n18 B.n17 585
R1810 B.n1398 B.n18 585
R1811 B.n1396 B.n1395 585
R1812 B.n1397 B.n1396 585
R1813 B.n1394 B.n23 585
R1814 B.n23 B.n22 585
R1815 B.n1393 B.n1392 585
R1816 B.n1392 B.n1391 585
R1817 B.n25 B.n24 585
R1818 B.n1390 B.n25 585
R1819 B.n1388 B.n1387 585
R1820 B.n1389 B.n1388 585
R1821 B.n1386 B.n30 585
R1822 B.n30 B.n29 585
R1823 B.n1385 B.n1384 585
R1824 B.n1384 B.n1383 585
R1825 B.n32 B.n31 585
R1826 B.n1382 B.n32 585
R1827 B.n1380 B.n1379 585
R1828 B.n1381 B.n1380 585
R1829 B.n1378 B.n37 585
R1830 B.n37 B.n36 585
R1831 B.n1377 B.n1376 585
R1832 B.n1376 B.n1375 585
R1833 B.n39 B.n38 585
R1834 B.n1374 B.n39 585
R1835 B.n1372 B.n1371 585
R1836 B.n1373 B.n1372 585
R1837 B.n1370 B.n44 585
R1838 B.n44 B.n43 585
R1839 B.n1369 B.n1368 585
R1840 B.n1368 B.n1367 585
R1841 B.n46 B.n45 585
R1842 B.n1366 B.n46 585
R1843 B.n1364 B.n1363 585
R1844 B.n1365 B.n1364 585
R1845 B.n1362 B.n51 585
R1846 B.n51 B.n50 585
R1847 B.n1361 B.n1360 585
R1848 B.n1360 B.n1359 585
R1849 B.n53 B.n52 585
R1850 B.n1358 B.n53 585
R1851 B.n1356 B.n1355 585
R1852 B.n1357 B.n1356 585
R1853 B.n1354 B.n58 585
R1854 B.n58 B.n57 585
R1855 B.n1353 B.n1352 585
R1856 B.n1352 B.n1351 585
R1857 B.n60 B.n59 585
R1858 B.n1350 B.n60 585
R1859 B.n1348 B.n1347 585
R1860 B.n1349 B.n1348 585
R1861 B.n1346 B.n65 585
R1862 B.n65 B.n64 585
R1863 B.n1345 B.n1344 585
R1864 B.n1344 B.n1343 585
R1865 B.n67 B.n66 585
R1866 B.n1342 B.n67 585
R1867 B.n1340 B.n1339 585
R1868 B.n1341 B.n1340 585
R1869 B.n1338 B.n72 585
R1870 B.n72 B.n71 585
R1871 B.n1337 B.n1336 585
R1872 B.n1336 B.n1335 585
R1873 B.n74 B.n73 585
R1874 B.n1334 B.n74 585
R1875 B.n1332 B.n1331 585
R1876 B.n1333 B.n1332 585
R1877 B.n1330 B.n78 585
R1878 B.n81 B.n78 585
R1879 B.n1329 B.n1328 585
R1880 B.n1328 B.n1327 585
R1881 B.n80 B.n79 585
R1882 B.n1326 B.n80 585
R1883 B.n1324 B.n1323 585
R1884 B.n1325 B.n1324 585
R1885 B.n1322 B.n86 585
R1886 B.n86 B.n85 585
R1887 B.n1321 B.n1320 585
R1888 B.n1320 B.n1319 585
R1889 B.n88 B.n87 585
R1890 B.n1318 B.n88 585
R1891 B.n1316 B.n1315 585
R1892 B.n1317 B.n1316 585
R1893 B.n1314 B.n93 585
R1894 B.n93 B.n92 585
R1895 B.n1313 B.n1312 585
R1896 B.n1312 B.n1311 585
R1897 B.n95 B.n94 585
R1898 B.n1310 B.n95 585
R1899 B.n1308 B.n1307 585
R1900 B.n1309 B.n1308 585
R1901 B.n1306 B.n99 585
R1902 B.n102 B.n99 585
R1903 B.n1305 B.n1304 585
R1904 B.n1304 B.n1303 585
R1905 B.n101 B.n100 585
R1906 B.n1302 B.n101 585
R1907 B.n1300 B.n1299 585
R1908 B.n1301 B.n1300 585
R1909 B.n1298 B.n107 585
R1910 B.n107 B.n106 585
R1911 B.n1297 B.n1296 585
R1912 B.n1296 B.n1295 585
R1913 B.n109 B.n108 585
R1914 B.n1294 B.n109 585
R1915 B.n1292 B.n1291 585
R1916 B.n1293 B.n1292 585
R1917 B.n1290 B.n114 585
R1918 B.n114 B.n113 585
R1919 B.n1289 B.n1288 585
R1920 B.n1288 B.n1287 585
R1921 B.n116 B.n115 585
R1922 B.n1286 B.n116 585
R1923 B.n1284 B.n1283 585
R1924 B.n1285 B.n1284 585
R1925 B.n1282 B.n121 585
R1926 B.n121 B.n120 585
R1927 B.n1281 B.n1280 585
R1928 B.n1280 B.n1279 585
R1929 B.n123 B.n122 585
R1930 B.n1278 B.n123 585
R1931 B.n1276 B.n1275 585
R1932 B.n1277 B.n1276 585
R1933 B.n1274 B.n128 585
R1934 B.n128 B.n127 585
R1935 B.n1273 B.n1272 585
R1936 B.n1272 B.n1271 585
R1937 B.n130 B.n129 585
R1938 B.n1270 B.n130 585
R1939 B.n1268 B.n1267 585
R1940 B.n1269 B.n1268 585
R1941 B.n1266 B.n135 585
R1942 B.n135 B.n134 585
R1943 B.n1265 B.n1264 585
R1944 B.n1264 B.n1263 585
R1945 B.n137 B.n136 585
R1946 B.n1262 B.n137 585
R1947 B.n1260 B.n1259 585
R1948 B.n1261 B.n1260 585
R1949 B.n1258 B.n142 585
R1950 B.n142 B.n141 585
R1951 B.n1417 B.n1416 585
R1952 B.n1416 B.n1415 585
R1953 B.n912 B.n602 444.452
R1954 B.n1256 B.n142 444.452
R1955 B.n664 B.n600 444.452
R1956 B.n1252 B.n205 444.452
R1957 B.n668 B.t14 444.286
R1958 B.n666 B.t17 444.286
R1959 B.n209 B.t19 444.286
R1960 B.n206 B.t9 444.286
R1961 B.n669 B.t13 366.517
R1962 B.n207 B.t10 366.517
R1963 B.n667 B.t16 366.517
R1964 B.n210 B.t20 366.517
R1965 B.n668 B.t11 319.86
R1966 B.n666 B.t15 319.86
R1967 B.n209 B.t18 319.86
R1968 B.n206 B.t7 319.86
R1969 B.n1254 B.n1253 256.663
R1970 B.n1254 B.n203 256.663
R1971 B.n1254 B.n202 256.663
R1972 B.n1254 B.n201 256.663
R1973 B.n1254 B.n200 256.663
R1974 B.n1254 B.n199 256.663
R1975 B.n1254 B.n198 256.663
R1976 B.n1254 B.n197 256.663
R1977 B.n1254 B.n196 256.663
R1978 B.n1254 B.n195 256.663
R1979 B.n1254 B.n194 256.663
R1980 B.n1254 B.n193 256.663
R1981 B.n1254 B.n192 256.663
R1982 B.n1254 B.n191 256.663
R1983 B.n1254 B.n190 256.663
R1984 B.n1254 B.n189 256.663
R1985 B.n1254 B.n188 256.663
R1986 B.n1254 B.n187 256.663
R1987 B.n1254 B.n186 256.663
R1988 B.n1254 B.n185 256.663
R1989 B.n1254 B.n184 256.663
R1990 B.n1254 B.n183 256.663
R1991 B.n1254 B.n182 256.663
R1992 B.n1254 B.n181 256.663
R1993 B.n1254 B.n180 256.663
R1994 B.n1254 B.n179 256.663
R1995 B.n1254 B.n178 256.663
R1996 B.n1254 B.n177 256.663
R1997 B.n1254 B.n176 256.663
R1998 B.n1254 B.n175 256.663
R1999 B.n1254 B.n174 256.663
R2000 B.n1254 B.n173 256.663
R2001 B.n1254 B.n172 256.663
R2002 B.n1254 B.n171 256.663
R2003 B.n1254 B.n170 256.663
R2004 B.n1254 B.n169 256.663
R2005 B.n1254 B.n168 256.663
R2006 B.n1254 B.n167 256.663
R2007 B.n1254 B.n166 256.663
R2008 B.n1254 B.n165 256.663
R2009 B.n1254 B.n164 256.663
R2010 B.n1254 B.n163 256.663
R2011 B.n1254 B.n162 256.663
R2012 B.n1254 B.n161 256.663
R2013 B.n1254 B.n160 256.663
R2014 B.n1254 B.n159 256.663
R2015 B.n1254 B.n158 256.663
R2016 B.n1254 B.n157 256.663
R2017 B.n1254 B.n156 256.663
R2018 B.n1254 B.n155 256.663
R2019 B.n1254 B.n154 256.663
R2020 B.n1254 B.n153 256.663
R2021 B.n1254 B.n152 256.663
R2022 B.n1254 B.n151 256.663
R2023 B.n1254 B.n150 256.663
R2024 B.n1254 B.n149 256.663
R2025 B.n1254 B.n148 256.663
R2026 B.n1254 B.n147 256.663
R2027 B.n1254 B.n146 256.663
R2028 B.n1254 B.n145 256.663
R2029 B.n1255 B.n1254 256.663
R2030 B.n911 B.n910 256.663
R2031 B.n910 B.n605 256.663
R2032 B.n910 B.n606 256.663
R2033 B.n910 B.n607 256.663
R2034 B.n910 B.n608 256.663
R2035 B.n910 B.n609 256.663
R2036 B.n910 B.n610 256.663
R2037 B.n910 B.n611 256.663
R2038 B.n910 B.n612 256.663
R2039 B.n910 B.n613 256.663
R2040 B.n910 B.n614 256.663
R2041 B.n910 B.n615 256.663
R2042 B.n910 B.n616 256.663
R2043 B.n910 B.n617 256.663
R2044 B.n910 B.n618 256.663
R2045 B.n910 B.n619 256.663
R2046 B.n910 B.n620 256.663
R2047 B.n910 B.n621 256.663
R2048 B.n910 B.n622 256.663
R2049 B.n910 B.n623 256.663
R2050 B.n910 B.n624 256.663
R2051 B.n910 B.n625 256.663
R2052 B.n910 B.n626 256.663
R2053 B.n910 B.n627 256.663
R2054 B.n910 B.n628 256.663
R2055 B.n910 B.n629 256.663
R2056 B.n910 B.n630 256.663
R2057 B.n910 B.n631 256.663
R2058 B.n910 B.n632 256.663
R2059 B.n910 B.n633 256.663
R2060 B.n910 B.n634 256.663
R2061 B.n910 B.n635 256.663
R2062 B.n910 B.n636 256.663
R2063 B.n910 B.n637 256.663
R2064 B.n910 B.n638 256.663
R2065 B.n910 B.n639 256.663
R2066 B.n910 B.n640 256.663
R2067 B.n910 B.n641 256.663
R2068 B.n910 B.n642 256.663
R2069 B.n910 B.n643 256.663
R2070 B.n910 B.n644 256.663
R2071 B.n910 B.n645 256.663
R2072 B.n910 B.n646 256.663
R2073 B.n910 B.n647 256.663
R2074 B.n910 B.n648 256.663
R2075 B.n910 B.n649 256.663
R2076 B.n910 B.n650 256.663
R2077 B.n910 B.n651 256.663
R2078 B.n910 B.n652 256.663
R2079 B.n910 B.n653 256.663
R2080 B.n910 B.n654 256.663
R2081 B.n910 B.n655 256.663
R2082 B.n910 B.n656 256.663
R2083 B.n910 B.n657 256.663
R2084 B.n910 B.n658 256.663
R2085 B.n910 B.n659 256.663
R2086 B.n910 B.n660 256.663
R2087 B.n910 B.n661 256.663
R2088 B.n910 B.n662 256.663
R2089 B.n910 B.n663 256.663
R2090 B.n916 B.n602 163.367
R2091 B.n916 B.n596 163.367
R2092 B.n924 B.n596 163.367
R2093 B.n924 B.n594 163.367
R2094 B.n928 B.n594 163.367
R2095 B.n928 B.n588 163.367
R2096 B.n936 B.n588 163.367
R2097 B.n936 B.n586 163.367
R2098 B.n940 B.n586 163.367
R2099 B.n940 B.n580 163.367
R2100 B.n948 B.n580 163.367
R2101 B.n948 B.n578 163.367
R2102 B.n952 B.n578 163.367
R2103 B.n952 B.n572 163.367
R2104 B.n960 B.n572 163.367
R2105 B.n960 B.n570 163.367
R2106 B.n964 B.n570 163.367
R2107 B.n964 B.n564 163.367
R2108 B.n972 B.n564 163.367
R2109 B.n972 B.n562 163.367
R2110 B.n976 B.n562 163.367
R2111 B.n976 B.n556 163.367
R2112 B.n985 B.n556 163.367
R2113 B.n985 B.n554 163.367
R2114 B.n989 B.n554 163.367
R2115 B.n989 B.n549 163.367
R2116 B.n997 B.n549 163.367
R2117 B.n997 B.n547 163.367
R2118 B.n1001 B.n547 163.367
R2119 B.n1001 B.n541 163.367
R2120 B.n1009 B.n541 163.367
R2121 B.n1009 B.n539 163.367
R2122 B.n1013 B.n539 163.367
R2123 B.n1013 B.n533 163.367
R2124 B.n1022 B.n533 163.367
R2125 B.n1022 B.n531 163.367
R2126 B.n1026 B.n531 163.367
R2127 B.n1026 B.n526 163.367
R2128 B.n1034 B.n526 163.367
R2129 B.n1034 B.n524 163.367
R2130 B.n1038 B.n524 163.367
R2131 B.n1038 B.n518 163.367
R2132 B.n1046 B.n518 163.367
R2133 B.n1046 B.n516 163.367
R2134 B.n1050 B.n516 163.367
R2135 B.n1050 B.n510 163.367
R2136 B.n1058 B.n510 163.367
R2137 B.n1058 B.n508 163.367
R2138 B.n1062 B.n508 163.367
R2139 B.n1062 B.n502 163.367
R2140 B.n1070 B.n502 163.367
R2141 B.n1070 B.n500 163.367
R2142 B.n1074 B.n500 163.367
R2143 B.n1074 B.n494 163.367
R2144 B.n1082 B.n494 163.367
R2145 B.n1082 B.n492 163.367
R2146 B.n1086 B.n492 163.367
R2147 B.n1086 B.n486 163.367
R2148 B.n1094 B.n486 163.367
R2149 B.n1094 B.n484 163.367
R2150 B.n1098 B.n484 163.367
R2151 B.n1098 B.n478 163.367
R2152 B.n1106 B.n478 163.367
R2153 B.n1106 B.n476 163.367
R2154 B.n1110 B.n476 163.367
R2155 B.n1110 B.n470 163.367
R2156 B.n1118 B.n470 163.367
R2157 B.n1118 B.n468 163.367
R2158 B.n1122 B.n468 163.367
R2159 B.n1122 B.n462 163.367
R2160 B.n1130 B.n462 163.367
R2161 B.n1130 B.n460 163.367
R2162 B.n1134 B.n460 163.367
R2163 B.n1134 B.n454 163.367
R2164 B.n1143 B.n454 163.367
R2165 B.n1143 B.n452 163.367
R2166 B.n1147 B.n452 163.367
R2167 B.n1147 B.n2 163.367
R2168 B.n1416 B.n2 163.367
R2169 B.n1416 B.n3 163.367
R2170 B.n1412 B.n3 163.367
R2171 B.n1412 B.n9 163.367
R2172 B.n1408 B.n9 163.367
R2173 B.n1408 B.n11 163.367
R2174 B.n1404 B.n11 163.367
R2175 B.n1404 B.n16 163.367
R2176 B.n1400 B.n16 163.367
R2177 B.n1400 B.n18 163.367
R2178 B.n1396 B.n18 163.367
R2179 B.n1396 B.n23 163.367
R2180 B.n1392 B.n23 163.367
R2181 B.n1392 B.n25 163.367
R2182 B.n1388 B.n25 163.367
R2183 B.n1388 B.n30 163.367
R2184 B.n1384 B.n30 163.367
R2185 B.n1384 B.n32 163.367
R2186 B.n1380 B.n32 163.367
R2187 B.n1380 B.n37 163.367
R2188 B.n1376 B.n37 163.367
R2189 B.n1376 B.n39 163.367
R2190 B.n1372 B.n39 163.367
R2191 B.n1372 B.n44 163.367
R2192 B.n1368 B.n44 163.367
R2193 B.n1368 B.n46 163.367
R2194 B.n1364 B.n46 163.367
R2195 B.n1364 B.n51 163.367
R2196 B.n1360 B.n51 163.367
R2197 B.n1360 B.n53 163.367
R2198 B.n1356 B.n53 163.367
R2199 B.n1356 B.n58 163.367
R2200 B.n1352 B.n58 163.367
R2201 B.n1352 B.n60 163.367
R2202 B.n1348 B.n60 163.367
R2203 B.n1348 B.n65 163.367
R2204 B.n1344 B.n65 163.367
R2205 B.n1344 B.n67 163.367
R2206 B.n1340 B.n67 163.367
R2207 B.n1340 B.n72 163.367
R2208 B.n1336 B.n72 163.367
R2209 B.n1336 B.n74 163.367
R2210 B.n1332 B.n74 163.367
R2211 B.n1332 B.n78 163.367
R2212 B.n1328 B.n78 163.367
R2213 B.n1328 B.n80 163.367
R2214 B.n1324 B.n80 163.367
R2215 B.n1324 B.n86 163.367
R2216 B.n1320 B.n86 163.367
R2217 B.n1320 B.n88 163.367
R2218 B.n1316 B.n88 163.367
R2219 B.n1316 B.n93 163.367
R2220 B.n1312 B.n93 163.367
R2221 B.n1312 B.n95 163.367
R2222 B.n1308 B.n95 163.367
R2223 B.n1308 B.n99 163.367
R2224 B.n1304 B.n99 163.367
R2225 B.n1304 B.n101 163.367
R2226 B.n1300 B.n101 163.367
R2227 B.n1300 B.n107 163.367
R2228 B.n1296 B.n107 163.367
R2229 B.n1296 B.n109 163.367
R2230 B.n1292 B.n109 163.367
R2231 B.n1292 B.n114 163.367
R2232 B.n1288 B.n114 163.367
R2233 B.n1288 B.n116 163.367
R2234 B.n1284 B.n116 163.367
R2235 B.n1284 B.n121 163.367
R2236 B.n1280 B.n121 163.367
R2237 B.n1280 B.n123 163.367
R2238 B.n1276 B.n123 163.367
R2239 B.n1276 B.n128 163.367
R2240 B.n1272 B.n128 163.367
R2241 B.n1272 B.n130 163.367
R2242 B.n1268 B.n130 163.367
R2243 B.n1268 B.n135 163.367
R2244 B.n1264 B.n135 163.367
R2245 B.n1264 B.n137 163.367
R2246 B.n1260 B.n137 163.367
R2247 B.n1260 B.n142 163.367
R2248 B.n909 B.n604 163.367
R2249 B.n909 B.n665 163.367
R2250 B.n905 B.n904 163.367
R2251 B.n901 B.n900 163.367
R2252 B.n897 B.n896 163.367
R2253 B.n893 B.n892 163.367
R2254 B.n889 B.n888 163.367
R2255 B.n885 B.n884 163.367
R2256 B.n881 B.n880 163.367
R2257 B.n877 B.n876 163.367
R2258 B.n873 B.n872 163.367
R2259 B.n869 B.n868 163.367
R2260 B.n865 B.n864 163.367
R2261 B.n861 B.n860 163.367
R2262 B.n857 B.n856 163.367
R2263 B.n853 B.n852 163.367
R2264 B.n849 B.n848 163.367
R2265 B.n845 B.n844 163.367
R2266 B.n841 B.n840 163.367
R2267 B.n837 B.n836 163.367
R2268 B.n833 B.n832 163.367
R2269 B.n829 B.n828 163.367
R2270 B.n825 B.n824 163.367
R2271 B.n821 B.n820 163.367
R2272 B.n817 B.n816 163.367
R2273 B.n813 B.n812 163.367
R2274 B.n809 B.n808 163.367
R2275 B.n805 B.n804 163.367
R2276 B.n800 B.n799 163.367
R2277 B.n796 B.n795 163.367
R2278 B.n792 B.n791 163.367
R2279 B.n788 B.n787 163.367
R2280 B.n784 B.n783 163.367
R2281 B.n779 B.n778 163.367
R2282 B.n775 B.n774 163.367
R2283 B.n771 B.n770 163.367
R2284 B.n767 B.n766 163.367
R2285 B.n763 B.n762 163.367
R2286 B.n759 B.n758 163.367
R2287 B.n755 B.n754 163.367
R2288 B.n751 B.n750 163.367
R2289 B.n747 B.n746 163.367
R2290 B.n743 B.n742 163.367
R2291 B.n739 B.n738 163.367
R2292 B.n735 B.n734 163.367
R2293 B.n731 B.n730 163.367
R2294 B.n727 B.n726 163.367
R2295 B.n723 B.n722 163.367
R2296 B.n719 B.n718 163.367
R2297 B.n715 B.n714 163.367
R2298 B.n711 B.n710 163.367
R2299 B.n707 B.n706 163.367
R2300 B.n703 B.n702 163.367
R2301 B.n699 B.n698 163.367
R2302 B.n695 B.n694 163.367
R2303 B.n691 B.n690 163.367
R2304 B.n687 B.n686 163.367
R2305 B.n683 B.n682 163.367
R2306 B.n679 B.n678 163.367
R2307 B.n675 B.n674 163.367
R2308 B.n671 B.n664 163.367
R2309 B.n918 B.n600 163.367
R2310 B.n918 B.n598 163.367
R2311 B.n922 B.n598 163.367
R2312 B.n922 B.n592 163.367
R2313 B.n930 B.n592 163.367
R2314 B.n930 B.n590 163.367
R2315 B.n934 B.n590 163.367
R2316 B.n934 B.n584 163.367
R2317 B.n942 B.n584 163.367
R2318 B.n942 B.n582 163.367
R2319 B.n946 B.n582 163.367
R2320 B.n946 B.n576 163.367
R2321 B.n954 B.n576 163.367
R2322 B.n954 B.n574 163.367
R2323 B.n958 B.n574 163.367
R2324 B.n958 B.n568 163.367
R2325 B.n966 B.n568 163.367
R2326 B.n966 B.n566 163.367
R2327 B.n970 B.n566 163.367
R2328 B.n970 B.n560 163.367
R2329 B.n978 B.n560 163.367
R2330 B.n978 B.n558 163.367
R2331 B.n982 B.n558 163.367
R2332 B.n982 B.n553 163.367
R2333 B.n991 B.n553 163.367
R2334 B.n991 B.n551 163.367
R2335 B.n995 B.n551 163.367
R2336 B.n995 B.n545 163.367
R2337 B.n1003 B.n545 163.367
R2338 B.n1003 B.n543 163.367
R2339 B.n1007 B.n543 163.367
R2340 B.n1007 B.n537 163.367
R2341 B.n1015 B.n537 163.367
R2342 B.n1015 B.n535 163.367
R2343 B.n1019 B.n535 163.367
R2344 B.n1019 B.n530 163.367
R2345 B.n1028 B.n530 163.367
R2346 B.n1028 B.n528 163.367
R2347 B.n1032 B.n528 163.367
R2348 B.n1032 B.n522 163.367
R2349 B.n1040 B.n522 163.367
R2350 B.n1040 B.n520 163.367
R2351 B.n1044 B.n520 163.367
R2352 B.n1044 B.n514 163.367
R2353 B.n1052 B.n514 163.367
R2354 B.n1052 B.n512 163.367
R2355 B.n1056 B.n512 163.367
R2356 B.n1056 B.n506 163.367
R2357 B.n1064 B.n506 163.367
R2358 B.n1064 B.n504 163.367
R2359 B.n1068 B.n504 163.367
R2360 B.n1068 B.n498 163.367
R2361 B.n1076 B.n498 163.367
R2362 B.n1076 B.n496 163.367
R2363 B.n1080 B.n496 163.367
R2364 B.n1080 B.n490 163.367
R2365 B.n1088 B.n490 163.367
R2366 B.n1088 B.n488 163.367
R2367 B.n1092 B.n488 163.367
R2368 B.n1092 B.n482 163.367
R2369 B.n1100 B.n482 163.367
R2370 B.n1100 B.n480 163.367
R2371 B.n1104 B.n480 163.367
R2372 B.n1104 B.n474 163.367
R2373 B.n1112 B.n474 163.367
R2374 B.n1112 B.n472 163.367
R2375 B.n1116 B.n472 163.367
R2376 B.n1116 B.n466 163.367
R2377 B.n1124 B.n466 163.367
R2378 B.n1124 B.n464 163.367
R2379 B.n1128 B.n464 163.367
R2380 B.n1128 B.n458 163.367
R2381 B.n1136 B.n458 163.367
R2382 B.n1136 B.n456 163.367
R2383 B.n1141 B.n456 163.367
R2384 B.n1141 B.n450 163.367
R2385 B.n1149 B.n450 163.367
R2386 B.n1150 B.n1149 163.367
R2387 B.n1150 B.n5 163.367
R2388 B.n6 B.n5 163.367
R2389 B.n7 B.n6 163.367
R2390 B.n1155 B.n7 163.367
R2391 B.n1155 B.n12 163.367
R2392 B.n13 B.n12 163.367
R2393 B.n14 B.n13 163.367
R2394 B.n1160 B.n14 163.367
R2395 B.n1160 B.n19 163.367
R2396 B.n20 B.n19 163.367
R2397 B.n21 B.n20 163.367
R2398 B.n1165 B.n21 163.367
R2399 B.n1165 B.n26 163.367
R2400 B.n27 B.n26 163.367
R2401 B.n28 B.n27 163.367
R2402 B.n1170 B.n28 163.367
R2403 B.n1170 B.n33 163.367
R2404 B.n34 B.n33 163.367
R2405 B.n35 B.n34 163.367
R2406 B.n1175 B.n35 163.367
R2407 B.n1175 B.n40 163.367
R2408 B.n41 B.n40 163.367
R2409 B.n42 B.n41 163.367
R2410 B.n1180 B.n42 163.367
R2411 B.n1180 B.n47 163.367
R2412 B.n48 B.n47 163.367
R2413 B.n49 B.n48 163.367
R2414 B.n1185 B.n49 163.367
R2415 B.n1185 B.n54 163.367
R2416 B.n55 B.n54 163.367
R2417 B.n56 B.n55 163.367
R2418 B.n1190 B.n56 163.367
R2419 B.n1190 B.n61 163.367
R2420 B.n62 B.n61 163.367
R2421 B.n63 B.n62 163.367
R2422 B.n1195 B.n63 163.367
R2423 B.n1195 B.n68 163.367
R2424 B.n69 B.n68 163.367
R2425 B.n70 B.n69 163.367
R2426 B.n1200 B.n70 163.367
R2427 B.n1200 B.n75 163.367
R2428 B.n76 B.n75 163.367
R2429 B.n77 B.n76 163.367
R2430 B.n1205 B.n77 163.367
R2431 B.n1205 B.n82 163.367
R2432 B.n83 B.n82 163.367
R2433 B.n84 B.n83 163.367
R2434 B.n1210 B.n84 163.367
R2435 B.n1210 B.n89 163.367
R2436 B.n90 B.n89 163.367
R2437 B.n91 B.n90 163.367
R2438 B.n1215 B.n91 163.367
R2439 B.n1215 B.n96 163.367
R2440 B.n97 B.n96 163.367
R2441 B.n98 B.n97 163.367
R2442 B.n1220 B.n98 163.367
R2443 B.n1220 B.n103 163.367
R2444 B.n104 B.n103 163.367
R2445 B.n105 B.n104 163.367
R2446 B.n1225 B.n105 163.367
R2447 B.n1225 B.n110 163.367
R2448 B.n111 B.n110 163.367
R2449 B.n112 B.n111 163.367
R2450 B.n1230 B.n112 163.367
R2451 B.n1230 B.n117 163.367
R2452 B.n118 B.n117 163.367
R2453 B.n119 B.n118 163.367
R2454 B.n1235 B.n119 163.367
R2455 B.n1235 B.n124 163.367
R2456 B.n125 B.n124 163.367
R2457 B.n126 B.n125 163.367
R2458 B.n1240 B.n126 163.367
R2459 B.n1240 B.n131 163.367
R2460 B.n132 B.n131 163.367
R2461 B.n133 B.n132 163.367
R2462 B.n1245 B.n133 163.367
R2463 B.n1245 B.n138 163.367
R2464 B.n139 B.n138 163.367
R2465 B.n140 B.n139 163.367
R2466 B.n205 B.n140 163.367
R2467 B.n212 B.n144 163.367
R2468 B.n216 B.n215 163.367
R2469 B.n220 B.n219 163.367
R2470 B.n224 B.n223 163.367
R2471 B.n228 B.n227 163.367
R2472 B.n232 B.n231 163.367
R2473 B.n236 B.n235 163.367
R2474 B.n240 B.n239 163.367
R2475 B.n244 B.n243 163.367
R2476 B.n248 B.n247 163.367
R2477 B.n252 B.n251 163.367
R2478 B.n256 B.n255 163.367
R2479 B.n260 B.n259 163.367
R2480 B.n264 B.n263 163.367
R2481 B.n268 B.n267 163.367
R2482 B.n272 B.n271 163.367
R2483 B.n276 B.n275 163.367
R2484 B.n280 B.n279 163.367
R2485 B.n284 B.n283 163.367
R2486 B.n288 B.n287 163.367
R2487 B.n292 B.n291 163.367
R2488 B.n296 B.n295 163.367
R2489 B.n300 B.n299 163.367
R2490 B.n304 B.n303 163.367
R2491 B.n308 B.n307 163.367
R2492 B.n312 B.n311 163.367
R2493 B.n316 B.n315 163.367
R2494 B.n320 B.n319 163.367
R2495 B.n324 B.n323 163.367
R2496 B.n328 B.n327 163.367
R2497 B.n332 B.n331 163.367
R2498 B.n336 B.n335 163.367
R2499 B.n340 B.n339 163.367
R2500 B.n344 B.n343 163.367
R2501 B.n348 B.n347 163.367
R2502 B.n352 B.n351 163.367
R2503 B.n356 B.n355 163.367
R2504 B.n360 B.n359 163.367
R2505 B.n364 B.n363 163.367
R2506 B.n368 B.n367 163.367
R2507 B.n372 B.n371 163.367
R2508 B.n376 B.n375 163.367
R2509 B.n380 B.n379 163.367
R2510 B.n384 B.n383 163.367
R2511 B.n388 B.n387 163.367
R2512 B.n392 B.n391 163.367
R2513 B.n396 B.n395 163.367
R2514 B.n400 B.n399 163.367
R2515 B.n404 B.n403 163.367
R2516 B.n408 B.n407 163.367
R2517 B.n412 B.n411 163.367
R2518 B.n416 B.n415 163.367
R2519 B.n420 B.n419 163.367
R2520 B.n424 B.n423 163.367
R2521 B.n428 B.n427 163.367
R2522 B.n432 B.n431 163.367
R2523 B.n436 B.n435 163.367
R2524 B.n440 B.n439 163.367
R2525 B.n444 B.n443 163.367
R2526 B.n446 B.n204 163.367
R2527 B.n669 B.n668 77.7702
R2528 B.n667 B.n666 77.7702
R2529 B.n210 B.n209 77.7702
R2530 B.n207 B.n206 77.7702
R2531 B.n912 B.n911 71.676
R2532 B.n665 B.n605 71.676
R2533 B.n904 B.n606 71.676
R2534 B.n900 B.n607 71.676
R2535 B.n896 B.n608 71.676
R2536 B.n892 B.n609 71.676
R2537 B.n888 B.n610 71.676
R2538 B.n884 B.n611 71.676
R2539 B.n880 B.n612 71.676
R2540 B.n876 B.n613 71.676
R2541 B.n872 B.n614 71.676
R2542 B.n868 B.n615 71.676
R2543 B.n864 B.n616 71.676
R2544 B.n860 B.n617 71.676
R2545 B.n856 B.n618 71.676
R2546 B.n852 B.n619 71.676
R2547 B.n848 B.n620 71.676
R2548 B.n844 B.n621 71.676
R2549 B.n840 B.n622 71.676
R2550 B.n836 B.n623 71.676
R2551 B.n832 B.n624 71.676
R2552 B.n828 B.n625 71.676
R2553 B.n824 B.n626 71.676
R2554 B.n820 B.n627 71.676
R2555 B.n816 B.n628 71.676
R2556 B.n812 B.n629 71.676
R2557 B.n808 B.n630 71.676
R2558 B.n804 B.n631 71.676
R2559 B.n799 B.n632 71.676
R2560 B.n795 B.n633 71.676
R2561 B.n791 B.n634 71.676
R2562 B.n787 B.n635 71.676
R2563 B.n783 B.n636 71.676
R2564 B.n778 B.n637 71.676
R2565 B.n774 B.n638 71.676
R2566 B.n770 B.n639 71.676
R2567 B.n766 B.n640 71.676
R2568 B.n762 B.n641 71.676
R2569 B.n758 B.n642 71.676
R2570 B.n754 B.n643 71.676
R2571 B.n750 B.n644 71.676
R2572 B.n746 B.n645 71.676
R2573 B.n742 B.n646 71.676
R2574 B.n738 B.n647 71.676
R2575 B.n734 B.n648 71.676
R2576 B.n730 B.n649 71.676
R2577 B.n726 B.n650 71.676
R2578 B.n722 B.n651 71.676
R2579 B.n718 B.n652 71.676
R2580 B.n714 B.n653 71.676
R2581 B.n710 B.n654 71.676
R2582 B.n706 B.n655 71.676
R2583 B.n702 B.n656 71.676
R2584 B.n698 B.n657 71.676
R2585 B.n694 B.n658 71.676
R2586 B.n690 B.n659 71.676
R2587 B.n686 B.n660 71.676
R2588 B.n682 B.n661 71.676
R2589 B.n678 B.n662 71.676
R2590 B.n674 B.n663 71.676
R2591 B.n1256 B.n1255 71.676
R2592 B.n212 B.n145 71.676
R2593 B.n216 B.n146 71.676
R2594 B.n220 B.n147 71.676
R2595 B.n224 B.n148 71.676
R2596 B.n228 B.n149 71.676
R2597 B.n232 B.n150 71.676
R2598 B.n236 B.n151 71.676
R2599 B.n240 B.n152 71.676
R2600 B.n244 B.n153 71.676
R2601 B.n248 B.n154 71.676
R2602 B.n252 B.n155 71.676
R2603 B.n256 B.n156 71.676
R2604 B.n260 B.n157 71.676
R2605 B.n264 B.n158 71.676
R2606 B.n268 B.n159 71.676
R2607 B.n272 B.n160 71.676
R2608 B.n276 B.n161 71.676
R2609 B.n280 B.n162 71.676
R2610 B.n284 B.n163 71.676
R2611 B.n288 B.n164 71.676
R2612 B.n292 B.n165 71.676
R2613 B.n296 B.n166 71.676
R2614 B.n300 B.n167 71.676
R2615 B.n304 B.n168 71.676
R2616 B.n308 B.n169 71.676
R2617 B.n312 B.n170 71.676
R2618 B.n316 B.n171 71.676
R2619 B.n320 B.n172 71.676
R2620 B.n324 B.n173 71.676
R2621 B.n328 B.n174 71.676
R2622 B.n332 B.n175 71.676
R2623 B.n336 B.n176 71.676
R2624 B.n340 B.n177 71.676
R2625 B.n344 B.n178 71.676
R2626 B.n348 B.n179 71.676
R2627 B.n352 B.n180 71.676
R2628 B.n356 B.n181 71.676
R2629 B.n360 B.n182 71.676
R2630 B.n364 B.n183 71.676
R2631 B.n368 B.n184 71.676
R2632 B.n372 B.n185 71.676
R2633 B.n376 B.n186 71.676
R2634 B.n380 B.n187 71.676
R2635 B.n384 B.n188 71.676
R2636 B.n388 B.n189 71.676
R2637 B.n392 B.n190 71.676
R2638 B.n396 B.n191 71.676
R2639 B.n400 B.n192 71.676
R2640 B.n404 B.n193 71.676
R2641 B.n408 B.n194 71.676
R2642 B.n412 B.n195 71.676
R2643 B.n416 B.n196 71.676
R2644 B.n420 B.n197 71.676
R2645 B.n424 B.n198 71.676
R2646 B.n428 B.n199 71.676
R2647 B.n432 B.n200 71.676
R2648 B.n436 B.n201 71.676
R2649 B.n440 B.n202 71.676
R2650 B.n444 B.n203 71.676
R2651 B.n1253 B.n204 71.676
R2652 B.n1253 B.n1252 71.676
R2653 B.n446 B.n203 71.676
R2654 B.n443 B.n202 71.676
R2655 B.n439 B.n201 71.676
R2656 B.n435 B.n200 71.676
R2657 B.n431 B.n199 71.676
R2658 B.n427 B.n198 71.676
R2659 B.n423 B.n197 71.676
R2660 B.n419 B.n196 71.676
R2661 B.n415 B.n195 71.676
R2662 B.n411 B.n194 71.676
R2663 B.n407 B.n193 71.676
R2664 B.n403 B.n192 71.676
R2665 B.n399 B.n191 71.676
R2666 B.n395 B.n190 71.676
R2667 B.n391 B.n189 71.676
R2668 B.n387 B.n188 71.676
R2669 B.n383 B.n187 71.676
R2670 B.n379 B.n186 71.676
R2671 B.n375 B.n185 71.676
R2672 B.n371 B.n184 71.676
R2673 B.n367 B.n183 71.676
R2674 B.n363 B.n182 71.676
R2675 B.n359 B.n181 71.676
R2676 B.n355 B.n180 71.676
R2677 B.n351 B.n179 71.676
R2678 B.n347 B.n178 71.676
R2679 B.n343 B.n177 71.676
R2680 B.n339 B.n176 71.676
R2681 B.n335 B.n175 71.676
R2682 B.n331 B.n174 71.676
R2683 B.n327 B.n173 71.676
R2684 B.n323 B.n172 71.676
R2685 B.n319 B.n171 71.676
R2686 B.n315 B.n170 71.676
R2687 B.n311 B.n169 71.676
R2688 B.n307 B.n168 71.676
R2689 B.n303 B.n167 71.676
R2690 B.n299 B.n166 71.676
R2691 B.n295 B.n165 71.676
R2692 B.n291 B.n164 71.676
R2693 B.n287 B.n163 71.676
R2694 B.n283 B.n162 71.676
R2695 B.n279 B.n161 71.676
R2696 B.n275 B.n160 71.676
R2697 B.n271 B.n159 71.676
R2698 B.n267 B.n158 71.676
R2699 B.n263 B.n157 71.676
R2700 B.n259 B.n156 71.676
R2701 B.n255 B.n155 71.676
R2702 B.n251 B.n154 71.676
R2703 B.n247 B.n153 71.676
R2704 B.n243 B.n152 71.676
R2705 B.n239 B.n151 71.676
R2706 B.n235 B.n150 71.676
R2707 B.n231 B.n149 71.676
R2708 B.n227 B.n148 71.676
R2709 B.n223 B.n147 71.676
R2710 B.n219 B.n146 71.676
R2711 B.n215 B.n145 71.676
R2712 B.n1255 B.n144 71.676
R2713 B.n911 B.n604 71.676
R2714 B.n905 B.n605 71.676
R2715 B.n901 B.n606 71.676
R2716 B.n897 B.n607 71.676
R2717 B.n893 B.n608 71.676
R2718 B.n889 B.n609 71.676
R2719 B.n885 B.n610 71.676
R2720 B.n881 B.n611 71.676
R2721 B.n877 B.n612 71.676
R2722 B.n873 B.n613 71.676
R2723 B.n869 B.n614 71.676
R2724 B.n865 B.n615 71.676
R2725 B.n861 B.n616 71.676
R2726 B.n857 B.n617 71.676
R2727 B.n853 B.n618 71.676
R2728 B.n849 B.n619 71.676
R2729 B.n845 B.n620 71.676
R2730 B.n841 B.n621 71.676
R2731 B.n837 B.n622 71.676
R2732 B.n833 B.n623 71.676
R2733 B.n829 B.n624 71.676
R2734 B.n825 B.n625 71.676
R2735 B.n821 B.n626 71.676
R2736 B.n817 B.n627 71.676
R2737 B.n813 B.n628 71.676
R2738 B.n809 B.n629 71.676
R2739 B.n805 B.n630 71.676
R2740 B.n800 B.n631 71.676
R2741 B.n796 B.n632 71.676
R2742 B.n792 B.n633 71.676
R2743 B.n788 B.n634 71.676
R2744 B.n784 B.n635 71.676
R2745 B.n779 B.n636 71.676
R2746 B.n775 B.n637 71.676
R2747 B.n771 B.n638 71.676
R2748 B.n767 B.n639 71.676
R2749 B.n763 B.n640 71.676
R2750 B.n759 B.n641 71.676
R2751 B.n755 B.n642 71.676
R2752 B.n751 B.n643 71.676
R2753 B.n747 B.n644 71.676
R2754 B.n743 B.n645 71.676
R2755 B.n739 B.n646 71.676
R2756 B.n735 B.n647 71.676
R2757 B.n731 B.n648 71.676
R2758 B.n727 B.n649 71.676
R2759 B.n723 B.n650 71.676
R2760 B.n719 B.n651 71.676
R2761 B.n715 B.n652 71.676
R2762 B.n711 B.n653 71.676
R2763 B.n707 B.n654 71.676
R2764 B.n703 B.n655 71.676
R2765 B.n699 B.n656 71.676
R2766 B.n695 B.n657 71.676
R2767 B.n691 B.n658 71.676
R2768 B.n687 B.n659 71.676
R2769 B.n683 B.n660 71.676
R2770 B.n679 B.n661 71.676
R2771 B.n675 B.n662 71.676
R2772 B.n671 B.n663 71.676
R2773 B.n781 B.n669 59.5399
R2774 B.n802 B.n667 59.5399
R2775 B.n211 B.n210 59.5399
R2776 B.n208 B.n207 59.5399
R2777 B.n910 B.n601 57.0725
R2778 B.n1254 B.n141 57.0725
R2779 B.n917 B.n601 33.7474
R2780 B.n917 B.n597 33.7474
R2781 B.n923 B.n597 33.7474
R2782 B.n923 B.n593 33.7474
R2783 B.n929 B.n593 33.7474
R2784 B.n929 B.n589 33.7474
R2785 B.n935 B.n589 33.7474
R2786 B.n935 B.n585 33.7474
R2787 B.n941 B.n585 33.7474
R2788 B.n947 B.n581 33.7474
R2789 B.n947 B.n577 33.7474
R2790 B.n953 B.n577 33.7474
R2791 B.n953 B.n573 33.7474
R2792 B.n959 B.n573 33.7474
R2793 B.n959 B.n569 33.7474
R2794 B.n965 B.n569 33.7474
R2795 B.n965 B.n565 33.7474
R2796 B.n971 B.n565 33.7474
R2797 B.n971 B.n561 33.7474
R2798 B.n977 B.n561 33.7474
R2799 B.n977 B.n557 33.7474
R2800 B.n984 B.n557 33.7474
R2801 B.n984 B.n983 33.7474
R2802 B.n990 B.n550 33.7474
R2803 B.n996 B.n550 33.7474
R2804 B.n996 B.n546 33.7474
R2805 B.n1002 B.n546 33.7474
R2806 B.n1002 B.n542 33.7474
R2807 B.n1008 B.n542 33.7474
R2808 B.n1008 B.n538 33.7474
R2809 B.n1014 B.n538 33.7474
R2810 B.n1014 B.n534 33.7474
R2811 B.n1021 B.n534 33.7474
R2812 B.n1021 B.n1020 33.7474
R2813 B.n1027 B.n527 33.7474
R2814 B.n1033 B.n527 33.7474
R2815 B.n1033 B.n523 33.7474
R2816 B.n1039 B.n523 33.7474
R2817 B.n1039 B.n519 33.7474
R2818 B.n1045 B.n519 33.7474
R2819 B.n1045 B.n515 33.7474
R2820 B.n1051 B.n515 33.7474
R2821 B.n1051 B.n511 33.7474
R2822 B.n1057 B.n511 33.7474
R2823 B.n1063 B.n507 33.7474
R2824 B.n1063 B.n503 33.7474
R2825 B.n1069 B.n503 33.7474
R2826 B.n1069 B.n499 33.7474
R2827 B.n1075 B.n499 33.7474
R2828 B.n1075 B.n495 33.7474
R2829 B.n1081 B.n495 33.7474
R2830 B.n1081 B.n491 33.7474
R2831 B.n1087 B.n491 33.7474
R2832 B.n1087 B.n487 33.7474
R2833 B.n1093 B.n487 33.7474
R2834 B.n1099 B.n483 33.7474
R2835 B.n1099 B.n479 33.7474
R2836 B.n1105 B.n479 33.7474
R2837 B.n1105 B.n475 33.7474
R2838 B.n1111 B.n475 33.7474
R2839 B.n1111 B.n471 33.7474
R2840 B.n1117 B.n471 33.7474
R2841 B.n1117 B.n467 33.7474
R2842 B.n1123 B.n467 33.7474
R2843 B.n1123 B.n463 33.7474
R2844 B.n1129 B.n463 33.7474
R2845 B.n1135 B.n459 33.7474
R2846 B.n1135 B.n455 33.7474
R2847 B.n1142 B.n455 33.7474
R2848 B.n1142 B.n451 33.7474
R2849 B.n1148 B.n451 33.7474
R2850 B.n1148 B.n4 33.7474
R2851 B.n1415 B.n4 33.7474
R2852 B.n1415 B.n1414 33.7474
R2853 B.n1414 B.n1413 33.7474
R2854 B.n1413 B.n8 33.7474
R2855 B.n1407 B.n8 33.7474
R2856 B.n1407 B.n1406 33.7474
R2857 B.n1406 B.n1405 33.7474
R2858 B.n1405 B.n15 33.7474
R2859 B.n1399 B.n1398 33.7474
R2860 B.n1398 B.n1397 33.7474
R2861 B.n1397 B.n22 33.7474
R2862 B.n1391 B.n22 33.7474
R2863 B.n1391 B.n1390 33.7474
R2864 B.n1390 B.n1389 33.7474
R2865 B.n1389 B.n29 33.7474
R2866 B.n1383 B.n29 33.7474
R2867 B.n1383 B.n1382 33.7474
R2868 B.n1382 B.n1381 33.7474
R2869 B.n1381 B.n36 33.7474
R2870 B.n1375 B.n1374 33.7474
R2871 B.n1374 B.n1373 33.7474
R2872 B.n1373 B.n43 33.7474
R2873 B.n1367 B.n43 33.7474
R2874 B.n1367 B.n1366 33.7474
R2875 B.n1366 B.n1365 33.7474
R2876 B.n1365 B.n50 33.7474
R2877 B.n1359 B.n50 33.7474
R2878 B.n1359 B.n1358 33.7474
R2879 B.n1358 B.n1357 33.7474
R2880 B.n1357 B.n57 33.7474
R2881 B.n1351 B.n1350 33.7474
R2882 B.n1350 B.n1349 33.7474
R2883 B.n1349 B.n64 33.7474
R2884 B.n1343 B.n64 33.7474
R2885 B.n1343 B.n1342 33.7474
R2886 B.n1342 B.n1341 33.7474
R2887 B.n1341 B.n71 33.7474
R2888 B.n1335 B.n71 33.7474
R2889 B.n1335 B.n1334 33.7474
R2890 B.n1334 B.n1333 33.7474
R2891 B.n1327 B.n81 33.7474
R2892 B.n1327 B.n1326 33.7474
R2893 B.n1326 B.n1325 33.7474
R2894 B.n1325 B.n85 33.7474
R2895 B.n1319 B.n85 33.7474
R2896 B.n1319 B.n1318 33.7474
R2897 B.n1318 B.n1317 33.7474
R2898 B.n1317 B.n92 33.7474
R2899 B.n1311 B.n92 33.7474
R2900 B.n1311 B.n1310 33.7474
R2901 B.n1310 B.n1309 33.7474
R2902 B.n1303 B.n102 33.7474
R2903 B.n1303 B.n1302 33.7474
R2904 B.n1302 B.n1301 33.7474
R2905 B.n1301 B.n106 33.7474
R2906 B.n1295 B.n106 33.7474
R2907 B.n1295 B.n1294 33.7474
R2908 B.n1294 B.n1293 33.7474
R2909 B.n1293 B.n113 33.7474
R2910 B.n1287 B.n113 33.7474
R2911 B.n1287 B.n1286 33.7474
R2912 B.n1286 B.n1285 33.7474
R2913 B.n1285 B.n120 33.7474
R2914 B.n1279 B.n120 33.7474
R2915 B.n1279 B.n1278 33.7474
R2916 B.n1277 B.n127 33.7474
R2917 B.n1271 B.n127 33.7474
R2918 B.n1271 B.n1270 33.7474
R2919 B.n1270 B.n1269 33.7474
R2920 B.n1269 B.n134 33.7474
R2921 B.n1263 B.n134 33.7474
R2922 B.n1263 B.n1262 33.7474
R2923 B.n1262 B.n1261 33.7474
R2924 B.n1261 B.n141 33.7474
R2925 B.n1057 B.t5 30.7697
R2926 B.n1351 B.t3 30.7697
R2927 B.n1027 B.t23 29.7772
R2928 B.n1333 B.t22 29.7772
R2929 B.n1251 B.n1250 28.8785
R2930 B.n1258 B.n1257 28.8785
R2931 B.n670 B.n599 28.8785
R2932 B.n914 B.n913 28.8785
R2933 B.n1093 B.t6 23.8218
R2934 B.n1375 B.t4 23.8218
R2935 B.t12 B.n581 22.8293
R2936 B.n990 B.t0 22.8293
R2937 B.n1309 B.t21 22.8293
R2938 B.n1278 B.t8 22.8293
R2939 B B.n1417 18.0485
R2940 B.n1129 B.t1 16.8739
R2941 B.t1 B.n459 16.8739
R2942 B.t2 B.n15 16.8739
R2943 B.n1399 B.t2 16.8739
R2944 B.n941 B.t12 10.9186
R2945 B.n983 B.t0 10.9186
R2946 B.n102 B.t21 10.9186
R2947 B.t8 B.n1277 10.9186
R2948 B.n1257 B.n143 10.6151
R2949 B.n213 B.n143 10.6151
R2950 B.n214 B.n213 10.6151
R2951 B.n217 B.n214 10.6151
R2952 B.n218 B.n217 10.6151
R2953 B.n221 B.n218 10.6151
R2954 B.n222 B.n221 10.6151
R2955 B.n225 B.n222 10.6151
R2956 B.n226 B.n225 10.6151
R2957 B.n229 B.n226 10.6151
R2958 B.n230 B.n229 10.6151
R2959 B.n233 B.n230 10.6151
R2960 B.n234 B.n233 10.6151
R2961 B.n237 B.n234 10.6151
R2962 B.n238 B.n237 10.6151
R2963 B.n241 B.n238 10.6151
R2964 B.n242 B.n241 10.6151
R2965 B.n245 B.n242 10.6151
R2966 B.n246 B.n245 10.6151
R2967 B.n249 B.n246 10.6151
R2968 B.n250 B.n249 10.6151
R2969 B.n253 B.n250 10.6151
R2970 B.n254 B.n253 10.6151
R2971 B.n257 B.n254 10.6151
R2972 B.n258 B.n257 10.6151
R2973 B.n261 B.n258 10.6151
R2974 B.n262 B.n261 10.6151
R2975 B.n265 B.n262 10.6151
R2976 B.n266 B.n265 10.6151
R2977 B.n269 B.n266 10.6151
R2978 B.n270 B.n269 10.6151
R2979 B.n273 B.n270 10.6151
R2980 B.n274 B.n273 10.6151
R2981 B.n277 B.n274 10.6151
R2982 B.n278 B.n277 10.6151
R2983 B.n281 B.n278 10.6151
R2984 B.n282 B.n281 10.6151
R2985 B.n285 B.n282 10.6151
R2986 B.n286 B.n285 10.6151
R2987 B.n289 B.n286 10.6151
R2988 B.n290 B.n289 10.6151
R2989 B.n293 B.n290 10.6151
R2990 B.n294 B.n293 10.6151
R2991 B.n297 B.n294 10.6151
R2992 B.n298 B.n297 10.6151
R2993 B.n301 B.n298 10.6151
R2994 B.n302 B.n301 10.6151
R2995 B.n305 B.n302 10.6151
R2996 B.n306 B.n305 10.6151
R2997 B.n309 B.n306 10.6151
R2998 B.n310 B.n309 10.6151
R2999 B.n313 B.n310 10.6151
R3000 B.n314 B.n313 10.6151
R3001 B.n317 B.n314 10.6151
R3002 B.n318 B.n317 10.6151
R3003 B.n322 B.n321 10.6151
R3004 B.n325 B.n322 10.6151
R3005 B.n326 B.n325 10.6151
R3006 B.n329 B.n326 10.6151
R3007 B.n330 B.n329 10.6151
R3008 B.n333 B.n330 10.6151
R3009 B.n334 B.n333 10.6151
R3010 B.n337 B.n334 10.6151
R3011 B.n338 B.n337 10.6151
R3012 B.n342 B.n341 10.6151
R3013 B.n345 B.n342 10.6151
R3014 B.n346 B.n345 10.6151
R3015 B.n349 B.n346 10.6151
R3016 B.n350 B.n349 10.6151
R3017 B.n353 B.n350 10.6151
R3018 B.n354 B.n353 10.6151
R3019 B.n357 B.n354 10.6151
R3020 B.n358 B.n357 10.6151
R3021 B.n361 B.n358 10.6151
R3022 B.n362 B.n361 10.6151
R3023 B.n365 B.n362 10.6151
R3024 B.n366 B.n365 10.6151
R3025 B.n369 B.n366 10.6151
R3026 B.n370 B.n369 10.6151
R3027 B.n373 B.n370 10.6151
R3028 B.n374 B.n373 10.6151
R3029 B.n377 B.n374 10.6151
R3030 B.n378 B.n377 10.6151
R3031 B.n381 B.n378 10.6151
R3032 B.n382 B.n381 10.6151
R3033 B.n385 B.n382 10.6151
R3034 B.n386 B.n385 10.6151
R3035 B.n389 B.n386 10.6151
R3036 B.n390 B.n389 10.6151
R3037 B.n393 B.n390 10.6151
R3038 B.n394 B.n393 10.6151
R3039 B.n397 B.n394 10.6151
R3040 B.n398 B.n397 10.6151
R3041 B.n401 B.n398 10.6151
R3042 B.n402 B.n401 10.6151
R3043 B.n405 B.n402 10.6151
R3044 B.n406 B.n405 10.6151
R3045 B.n409 B.n406 10.6151
R3046 B.n410 B.n409 10.6151
R3047 B.n413 B.n410 10.6151
R3048 B.n414 B.n413 10.6151
R3049 B.n417 B.n414 10.6151
R3050 B.n418 B.n417 10.6151
R3051 B.n421 B.n418 10.6151
R3052 B.n422 B.n421 10.6151
R3053 B.n425 B.n422 10.6151
R3054 B.n426 B.n425 10.6151
R3055 B.n429 B.n426 10.6151
R3056 B.n430 B.n429 10.6151
R3057 B.n433 B.n430 10.6151
R3058 B.n434 B.n433 10.6151
R3059 B.n437 B.n434 10.6151
R3060 B.n438 B.n437 10.6151
R3061 B.n441 B.n438 10.6151
R3062 B.n442 B.n441 10.6151
R3063 B.n445 B.n442 10.6151
R3064 B.n447 B.n445 10.6151
R3065 B.n448 B.n447 10.6151
R3066 B.n1251 B.n448 10.6151
R3067 B.n919 B.n599 10.6151
R3068 B.n920 B.n919 10.6151
R3069 B.n921 B.n920 10.6151
R3070 B.n921 B.n591 10.6151
R3071 B.n931 B.n591 10.6151
R3072 B.n932 B.n931 10.6151
R3073 B.n933 B.n932 10.6151
R3074 B.n933 B.n583 10.6151
R3075 B.n943 B.n583 10.6151
R3076 B.n944 B.n943 10.6151
R3077 B.n945 B.n944 10.6151
R3078 B.n945 B.n575 10.6151
R3079 B.n955 B.n575 10.6151
R3080 B.n956 B.n955 10.6151
R3081 B.n957 B.n956 10.6151
R3082 B.n957 B.n567 10.6151
R3083 B.n967 B.n567 10.6151
R3084 B.n968 B.n967 10.6151
R3085 B.n969 B.n968 10.6151
R3086 B.n969 B.n559 10.6151
R3087 B.n979 B.n559 10.6151
R3088 B.n980 B.n979 10.6151
R3089 B.n981 B.n980 10.6151
R3090 B.n981 B.n552 10.6151
R3091 B.n992 B.n552 10.6151
R3092 B.n993 B.n992 10.6151
R3093 B.n994 B.n993 10.6151
R3094 B.n994 B.n544 10.6151
R3095 B.n1004 B.n544 10.6151
R3096 B.n1005 B.n1004 10.6151
R3097 B.n1006 B.n1005 10.6151
R3098 B.n1006 B.n536 10.6151
R3099 B.n1016 B.n536 10.6151
R3100 B.n1017 B.n1016 10.6151
R3101 B.n1018 B.n1017 10.6151
R3102 B.n1018 B.n529 10.6151
R3103 B.n1029 B.n529 10.6151
R3104 B.n1030 B.n1029 10.6151
R3105 B.n1031 B.n1030 10.6151
R3106 B.n1031 B.n521 10.6151
R3107 B.n1041 B.n521 10.6151
R3108 B.n1042 B.n1041 10.6151
R3109 B.n1043 B.n1042 10.6151
R3110 B.n1043 B.n513 10.6151
R3111 B.n1053 B.n513 10.6151
R3112 B.n1054 B.n1053 10.6151
R3113 B.n1055 B.n1054 10.6151
R3114 B.n1055 B.n505 10.6151
R3115 B.n1065 B.n505 10.6151
R3116 B.n1066 B.n1065 10.6151
R3117 B.n1067 B.n1066 10.6151
R3118 B.n1067 B.n497 10.6151
R3119 B.n1077 B.n497 10.6151
R3120 B.n1078 B.n1077 10.6151
R3121 B.n1079 B.n1078 10.6151
R3122 B.n1079 B.n489 10.6151
R3123 B.n1089 B.n489 10.6151
R3124 B.n1090 B.n1089 10.6151
R3125 B.n1091 B.n1090 10.6151
R3126 B.n1091 B.n481 10.6151
R3127 B.n1101 B.n481 10.6151
R3128 B.n1102 B.n1101 10.6151
R3129 B.n1103 B.n1102 10.6151
R3130 B.n1103 B.n473 10.6151
R3131 B.n1113 B.n473 10.6151
R3132 B.n1114 B.n1113 10.6151
R3133 B.n1115 B.n1114 10.6151
R3134 B.n1115 B.n465 10.6151
R3135 B.n1125 B.n465 10.6151
R3136 B.n1126 B.n1125 10.6151
R3137 B.n1127 B.n1126 10.6151
R3138 B.n1127 B.n457 10.6151
R3139 B.n1137 B.n457 10.6151
R3140 B.n1138 B.n1137 10.6151
R3141 B.n1140 B.n1138 10.6151
R3142 B.n1140 B.n1139 10.6151
R3143 B.n1139 B.n449 10.6151
R3144 B.n1151 B.n449 10.6151
R3145 B.n1152 B.n1151 10.6151
R3146 B.n1153 B.n1152 10.6151
R3147 B.n1154 B.n1153 10.6151
R3148 B.n1156 B.n1154 10.6151
R3149 B.n1157 B.n1156 10.6151
R3150 B.n1158 B.n1157 10.6151
R3151 B.n1159 B.n1158 10.6151
R3152 B.n1161 B.n1159 10.6151
R3153 B.n1162 B.n1161 10.6151
R3154 B.n1163 B.n1162 10.6151
R3155 B.n1164 B.n1163 10.6151
R3156 B.n1166 B.n1164 10.6151
R3157 B.n1167 B.n1166 10.6151
R3158 B.n1168 B.n1167 10.6151
R3159 B.n1169 B.n1168 10.6151
R3160 B.n1171 B.n1169 10.6151
R3161 B.n1172 B.n1171 10.6151
R3162 B.n1173 B.n1172 10.6151
R3163 B.n1174 B.n1173 10.6151
R3164 B.n1176 B.n1174 10.6151
R3165 B.n1177 B.n1176 10.6151
R3166 B.n1178 B.n1177 10.6151
R3167 B.n1179 B.n1178 10.6151
R3168 B.n1181 B.n1179 10.6151
R3169 B.n1182 B.n1181 10.6151
R3170 B.n1183 B.n1182 10.6151
R3171 B.n1184 B.n1183 10.6151
R3172 B.n1186 B.n1184 10.6151
R3173 B.n1187 B.n1186 10.6151
R3174 B.n1188 B.n1187 10.6151
R3175 B.n1189 B.n1188 10.6151
R3176 B.n1191 B.n1189 10.6151
R3177 B.n1192 B.n1191 10.6151
R3178 B.n1193 B.n1192 10.6151
R3179 B.n1194 B.n1193 10.6151
R3180 B.n1196 B.n1194 10.6151
R3181 B.n1197 B.n1196 10.6151
R3182 B.n1198 B.n1197 10.6151
R3183 B.n1199 B.n1198 10.6151
R3184 B.n1201 B.n1199 10.6151
R3185 B.n1202 B.n1201 10.6151
R3186 B.n1203 B.n1202 10.6151
R3187 B.n1204 B.n1203 10.6151
R3188 B.n1206 B.n1204 10.6151
R3189 B.n1207 B.n1206 10.6151
R3190 B.n1208 B.n1207 10.6151
R3191 B.n1209 B.n1208 10.6151
R3192 B.n1211 B.n1209 10.6151
R3193 B.n1212 B.n1211 10.6151
R3194 B.n1213 B.n1212 10.6151
R3195 B.n1214 B.n1213 10.6151
R3196 B.n1216 B.n1214 10.6151
R3197 B.n1217 B.n1216 10.6151
R3198 B.n1218 B.n1217 10.6151
R3199 B.n1219 B.n1218 10.6151
R3200 B.n1221 B.n1219 10.6151
R3201 B.n1222 B.n1221 10.6151
R3202 B.n1223 B.n1222 10.6151
R3203 B.n1224 B.n1223 10.6151
R3204 B.n1226 B.n1224 10.6151
R3205 B.n1227 B.n1226 10.6151
R3206 B.n1228 B.n1227 10.6151
R3207 B.n1229 B.n1228 10.6151
R3208 B.n1231 B.n1229 10.6151
R3209 B.n1232 B.n1231 10.6151
R3210 B.n1233 B.n1232 10.6151
R3211 B.n1234 B.n1233 10.6151
R3212 B.n1236 B.n1234 10.6151
R3213 B.n1237 B.n1236 10.6151
R3214 B.n1238 B.n1237 10.6151
R3215 B.n1239 B.n1238 10.6151
R3216 B.n1241 B.n1239 10.6151
R3217 B.n1242 B.n1241 10.6151
R3218 B.n1243 B.n1242 10.6151
R3219 B.n1244 B.n1243 10.6151
R3220 B.n1246 B.n1244 10.6151
R3221 B.n1247 B.n1246 10.6151
R3222 B.n1248 B.n1247 10.6151
R3223 B.n1249 B.n1248 10.6151
R3224 B.n1250 B.n1249 10.6151
R3225 B.n913 B.n603 10.6151
R3226 B.n908 B.n603 10.6151
R3227 B.n908 B.n907 10.6151
R3228 B.n907 B.n906 10.6151
R3229 B.n906 B.n903 10.6151
R3230 B.n903 B.n902 10.6151
R3231 B.n902 B.n899 10.6151
R3232 B.n899 B.n898 10.6151
R3233 B.n898 B.n895 10.6151
R3234 B.n895 B.n894 10.6151
R3235 B.n894 B.n891 10.6151
R3236 B.n891 B.n890 10.6151
R3237 B.n890 B.n887 10.6151
R3238 B.n887 B.n886 10.6151
R3239 B.n886 B.n883 10.6151
R3240 B.n883 B.n882 10.6151
R3241 B.n882 B.n879 10.6151
R3242 B.n879 B.n878 10.6151
R3243 B.n878 B.n875 10.6151
R3244 B.n875 B.n874 10.6151
R3245 B.n874 B.n871 10.6151
R3246 B.n871 B.n870 10.6151
R3247 B.n870 B.n867 10.6151
R3248 B.n867 B.n866 10.6151
R3249 B.n866 B.n863 10.6151
R3250 B.n863 B.n862 10.6151
R3251 B.n862 B.n859 10.6151
R3252 B.n859 B.n858 10.6151
R3253 B.n858 B.n855 10.6151
R3254 B.n855 B.n854 10.6151
R3255 B.n854 B.n851 10.6151
R3256 B.n851 B.n850 10.6151
R3257 B.n850 B.n847 10.6151
R3258 B.n847 B.n846 10.6151
R3259 B.n846 B.n843 10.6151
R3260 B.n843 B.n842 10.6151
R3261 B.n842 B.n839 10.6151
R3262 B.n839 B.n838 10.6151
R3263 B.n838 B.n835 10.6151
R3264 B.n835 B.n834 10.6151
R3265 B.n834 B.n831 10.6151
R3266 B.n831 B.n830 10.6151
R3267 B.n830 B.n827 10.6151
R3268 B.n827 B.n826 10.6151
R3269 B.n826 B.n823 10.6151
R3270 B.n823 B.n822 10.6151
R3271 B.n822 B.n819 10.6151
R3272 B.n819 B.n818 10.6151
R3273 B.n818 B.n815 10.6151
R3274 B.n815 B.n814 10.6151
R3275 B.n814 B.n811 10.6151
R3276 B.n811 B.n810 10.6151
R3277 B.n810 B.n807 10.6151
R3278 B.n807 B.n806 10.6151
R3279 B.n806 B.n803 10.6151
R3280 B.n801 B.n798 10.6151
R3281 B.n798 B.n797 10.6151
R3282 B.n797 B.n794 10.6151
R3283 B.n794 B.n793 10.6151
R3284 B.n793 B.n790 10.6151
R3285 B.n790 B.n789 10.6151
R3286 B.n789 B.n786 10.6151
R3287 B.n786 B.n785 10.6151
R3288 B.n785 B.n782 10.6151
R3289 B.n780 B.n777 10.6151
R3290 B.n777 B.n776 10.6151
R3291 B.n776 B.n773 10.6151
R3292 B.n773 B.n772 10.6151
R3293 B.n772 B.n769 10.6151
R3294 B.n769 B.n768 10.6151
R3295 B.n768 B.n765 10.6151
R3296 B.n765 B.n764 10.6151
R3297 B.n764 B.n761 10.6151
R3298 B.n761 B.n760 10.6151
R3299 B.n760 B.n757 10.6151
R3300 B.n757 B.n756 10.6151
R3301 B.n756 B.n753 10.6151
R3302 B.n753 B.n752 10.6151
R3303 B.n752 B.n749 10.6151
R3304 B.n749 B.n748 10.6151
R3305 B.n748 B.n745 10.6151
R3306 B.n745 B.n744 10.6151
R3307 B.n744 B.n741 10.6151
R3308 B.n741 B.n740 10.6151
R3309 B.n740 B.n737 10.6151
R3310 B.n737 B.n736 10.6151
R3311 B.n736 B.n733 10.6151
R3312 B.n733 B.n732 10.6151
R3313 B.n732 B.n729 10.6151
R3314 B.n729 B.n728 10.6151
R3315 B.n728 B.n725 10.6151
R3316 B.n725 B.n724 10.6151
R3317 B.n724 B.n721 10.6151
R3318 B.n721 B.n720 10.6151
R3319 B.n720 B.n717 10.6151
R3320 B.n717 B.n716 10.6151
R3321 B.n716 B.n713 10.6151
R3322 B.n713 B.n712 10.6151
R3323 B.n712 B.n709 10.6151
R3324 B.n709 B.n708 10.6151
R3325 B.n708 B.n705 10.6151
R3326 B.n705 B.n704 10.6151
R3327 B.n704 B.n701 10.6151
R3328 B.n701 B.n700 10.6151
R3329 B.n700 B.n697 10.6151
R3330 B.n697 B.n696 10.6151
R3331 B.n696 B.n693 10.6151
R3332 B.n693 B.n692 10.6151
R3333 B.n692 B.n689 10.6151
R3334 B.n689 B.n688 10.6151
R3335 B.n688 B.n685 10.6151
R3336 B.n685 B.n684 10.6151
R3337 B.n684 B.n681 10.6151
R3338 B.n681 B.n680 10.6151
R3339 B.n680 B.n677 10.6151
R3340 B.n677 B.n676 10.6151
R3341 B.n676 B.n673 10.6151
R3342 B.n673 B.n672 10.6151
R3343 B.n672 B.n670 10.6151
R3344 B.n915 B.n914 10.6151
R3345 B.n915 B.n595 10.6151
R3346 B.n925 B.n595 10.6151
R3347 B.n926 B.n925 10.6151
R3348 B.n927 B.n926 10.6151
R3349 B.n927 B.n587 10.6151
R3350 B.n937 B.n587 10.6151
R3351 B.n938 B.n937 10.6151
R3352 B.n939 B.n938 10.6151
R3353 B.n939 B.n579 10.6151
R3354 B.n949 B.n579 10.6151
R3355 B.n950 B.n949 10.6151
R3356 B.n951 B.n950 10.6151
R3357 B.n951 B.n571 10.6151
R3358 B.n961 B.n571 10.6151
R3359 B.n962 B.n961 10.6151
R3360 B.n963 B.n962 10.6151
R3361 B.n963 B.n563 10.6151
R3362 B.n973 B.n563 10.6151
R3363 B.n974 B.n973 10.6151
R3364 B.n975 B.n974 10.6151
R3365 B.n975 B.n555 10.6151
R3366 B.n986 B.n555 10.6151
R3367 B.n987 B.n986 10.6151
R3368 B.n988 B.n987 10.6151
R3369 B.n988 B.n548 10.6151
R3370 B.n998 B.n548 10.6151
R3371 B.n999 B.n998 10.6151
R3372 B.n1000 B.n999 10.6151
R3373 B.n1000 B.n540 10.6151
R3374 B.n1010 B.n540 10.6151
R3375 B.n1011 B.n1010 10.6151
R3376 B.n1012 B.n1011 10.6151
R3377 B.n1012 B.n532 10.6151
R3378 B.n1023 B.n532 10.6151
R3379 B.n1024 B.n1023 10.6151
R3380 B.n1025 B.n1024 10.6151
R3381 B.n1025 B.n525 10.6151
R3382 B.n1035 B.n525 10.6151
R3383 B.n1036 B.n1035 10.6151
R3384 B.n1037 B.n1036 10.6151
R3385 B.n1037 B.n517 10.6151
R3386 B.n1047 B.n517 10.6151
R3387 B.n1048 B.n1047 10.6151
R3388 B.n1049 B.n1048 10.6151
R3389 B.n1049 B.n509 10.6151
R3390 B.n1059 B.n509 10.6151
R3391 B.n1060 B.n1059 10.6151
R3392 B.n1061 B.n1060 10.6151
R3393 B.n1061 B.n501 10.6151
R3394 B.n1071 B.n501 10.6151
R3395 B.n1072 B.n1071 10.6151
R3396 B.n1073 B.n1072 10.6151
R3397 B.n1073 B.n493 10.6151
R3398 B.n1083 B.n493 10.6151
R3399 B.n1084 B.n1083 10.6151
R3400 B.n1085 B.n1084 10.6151
R3401 B.n1085 B.n485 10.6151
R3402 B.n1095 B.n485 10.6151
R3403 B.n1096 B.n1095 10.6151
R3404 B.n1097 B.n1096 10.6151
R3405 B.n1097 B.n477 10.6151
R3406 B.n1107 B.n477 10.6151
R3407 B.n1108 B.n1107 10.6151
R3408 B.n1109 B.n1108 10.6151
R3409 B.n1109 B.n469 10.6151
R3410 B.n1119 B.n469 10.6151
R3411 B.n1120 B.n1119 10.6151
R3412 B.n1121 B.n1120 10.6151
R3413 B.n1121 B.n461 10.6151
R3414 B.n1131 B.n461 10.6151
R3415 B.n1132 B.n1131 10.6151
R3416 B.n1133 B.n1132 10.6151
R3417 B.n1133 B.n453 10.6151
R3418 B.n1144 B.n453 10.6151
R3419 B.n1145 B.n1144 10.6151
R3420 B.n1146 B.n1145 10.6151
R3421 B.n1146 B.n0 10.6151
R3422 B.n1411 B.n1 10.6151
R3423 B.n1411 B.n1410 10.6151
R3424 B.n1410 B.n1409 10.6151
R3425 B.n1409 B.n10 10.6151
R3426 B.n1403 B.n10 10.6151
R3427 B.n1403 B.n1402 10.6151
R3428 B.n1402 B.n1401 10.6151
R3429 B.n1401 B.n17 10.6151
R3430 B.n1395 B.n17 10.6151
R3431 B.n1395 B.n1394 10.6151
R3432 B.n1394 B.n1393 10.6151
R3433 B.n1393 B.n24 10.6151
R3434 B.n1387 B.n24 10.6151
R3435 B.n1387 B.n1386 10.6151
R3436 B.n1386 B.n1385 10.6151
R3437 B.n1385 B.n31 10.6151
R3438 B.n1379 B.n31 10.6151
R3439 B.n1379 B.n1378 10.6151
R3440 B.n1378 B.n1377 10.6151
R3441 B.n1377 B.n38 10.6151
R3442 B.n1371 B.n38 10.6151
R3443 B.n1371 B.n1370 10.6151
R3444 B.n1370 B.n1369 10.6151
R3445 B.n1369 B.n45 10.6151
R3446 B.n1363 B.n45 10.6151
R3447 B.n1363 B.n1362 10.6151
R3448 B.n1362 B.n1361 10.6151
R3449 B.n1361 B.n52 10.6151
R3450 B.n1355 B.n52 10.6151
R3451 B.n1355 B.n1354 10.6151
R3452 B.n1354 B.n1353 10.6151
R3453 B.n1353 B.n59 10.6151
R3454 B.n1347 B.n59 10.6151
R3455 B.n1347 B.n1346 10.6151
R3456 B.n1346 B.n1345 10.6151
R3457 B.n1345 B.n66 10.6151
R3458 B.n1339 B.n66 10.6151
R3459 B.n1339 B.n1338 10.6151
R3460 B.n1338 B.n1337 10.6151
R3461 B.n1337 B.n73 10.6151
R3462 B.n1331 B.n73 10.6151
R3463 B.n1331 B.n1330 10.6151
R3464 B.n1330 B.n1329 10.6151
R3465 B.n1329 B.n79 10.6151
R3466 B.n1323 B.n79 10.6151
R3467 B.n1323 B.n1322 10.6151
R3468 B.n1322 B.n1321 10.6151
R3469 B.n1321 B.n87 10.6151
R3470 B.n1315 B.n87 10.6151
R3471 B.n1315 B.n1314 10.6151
R3472 B.n1314 B.n1313 10.6151
R3473 B.n1313 B.n94 10.6151
R3474 B.n1307 B.n94 10.6151
R3475 B.n1307 B.n1306 10.6151
R3476 B.n1306 B.n1305 10.6151
R3477 B.n1305 B.n100 10.6151
R3478 B.n1299 B.n100 10.6151
R3479 B.n1299 B.n1298 10.6151
R3480 B.n1298 B.n1297 10.6151
R3481 B.n1297 B.n108 10.6151
R3482 B.n1291 B.n108 10.6151
R3483 B.n1291 B.n1290 10.6151
R3484 B.n1290 B.n1289 10.6151
R3485 B.n1289 B.n115 10.6151
R3486 B.n1283 B.n115 10.6151
R3487 B.n1283 B.n1282 10.6151
R3488 B.n1282 B.n1281 10.6151
R3489 B.n1281 B.n122 10.6151
R3490 B.n1275 B.n122 10.6151
R3491 B.n1275 B.n1274 10.6151
R3492 B.n1274 B.n1273 10.6151
R3493 B.n1273 B.n129 10.6151
R3494 B.n1267 B.n129 10.6151
R3495 B.n1267 B.n1266 10.6151
R3496 B.n1266 B.n1265 10.6151
R3497 B.n1265 B.n136 10.6151
R3498 B.n1259 B.n136 10.6151
R3499 B.n1259 B.n1258 10.6151
R3500 B.t6 B.n483 9.92606
R3501 B.t4 B.n36 9.92606
R3502 B.n318 B.n211 9.36635
R3503 B.n341 B.n208 9.36635
R3504 B.n803 B.n802 9.36635
R3505 B.n781 B.n780 9.36635
R3506 B.n1020 B.t23 3.97072
R3507 B.n81 B.t22 3.97072
R3508 B.t5 B.n507 2.97817
R3509 B.t3 B.n57 2.97817
R3510 B.n1417 B.n0 2.81026
R3511 B.n1417 B.n1 2.81026
R3512 B.n321 B.n211 1.24928
R3513 B.n338 B.n208 1.24928
R3514 B.n802 B.n801 1.24928
R3515 B.n782 B.n781 1.24928
R3516 VP.n33 VP.n32 161.3
R3517 VP.n34 VP.n29 161.3
R3518 VP.n36 VP.n35 161.3
R3519 VP.n37 VP.n28 161.3
R3520 VP.n39 VP.n38 161.3
R3521 VP.n40 VP.n27 161.3
R3522 VP.n42 VP.n41 161.3
R3523 VP.n43 VP.n26 161.3
R3524 VP.n45 VP.n44 161.3
R3525 VP.n46 VP.n25 161.3
R3526 VP.n48 VP.n47 161.3
R3527 VP.n49 VP.n24 161.3
R3528 VP.n51 VP.n50 161.3
R3529 VP.n52 VP.n23 161.3
R3530 VP.n54 VP.n53 161.3
R3531 VP.n55 VP.n22 161.3
R3532 VP.n58 VP.n57 161.3
R3533 VP.n59 VP.n21 161.3
R3534 VP.n61 VP.n60 161.3
R3535 VP.n62 VP.n20 161.3
R3536 VP.n64 VP.n63 161.3
R3537 VP.n65 VP.n19 161.3
R3538 VP.n67 VP.n66 161.3
R3539 VP.n68 VP.n18 161.3
R3540 VP.n70 VP.n69 161.3
R3541 VP.n125 VP.n124 161.3
R3542 VP.n123 VP.n1 161.3
R3543 VP.n122 VP.n121 161.3
R3544 VP.n120 VP.n2 161.3
R3545 VP.n119 VP.n118 161.3
R3546 VP.n117 VP.n3 161.3
R3547 VP.n116 VP.n115 161.3
R3548 VP.n114 VP.n4 161.3
R3549 VP.n113 VP.n112 161.3
R3550 VP.n110 VP.n5 161.3
R3551 VP.n109 VP.n108 161.3
R3552 VP.n107 VP.n6 161.3
R3553 VP.n106 VP.n105 161.3
R3554 VP.n104 VP.n7 161.3
R3555 VP.n103 VP.n102 161.3
R3556 VP.n101 VP.n8 161.3
R3557 VP.n100 VP.n99 161.3
R3558 VP.n98 VP.n9 161.3
R3559 VP.n97 VP.n96 161.3
R3560 VP.n95 VP.n10 161.3
R3561 VP.n94 VP.n93 161.3
R3562 VP.n92 VP.n11 161.3
R3563 VP.n91 VP.n90 161.3
R3564 VP.n89 VP.n12 161.3
R3565 VP.n88 VP.n87 161.3
R3566 VP.n85 VP.n13 161.3
R3567 VP.n84 VP.n83 161.3
R3568 VP.n82 VP.n14 161.3
R3569 VP.n81 VP.n80 161.3
R3570 VP.n79 VP.n15 161.3
R3571 VP.n78 VP.n77 161.3
R3572 VP.n76 VP.n16 161.3
R3573 VP.n75 VP.n74 161.3
R3574 VP.n30 VP.t5 141.931
R3575 VP.n99 VP.t8 110.612
R3576 VP.n73 VP.t7 110.612
R3577 VP.n86 VP.t2 110.612
R3578 VP.n111 VP.t1 110.612
R3579 VP.n0 VP.t6 110.612
R3580 VP.n44 VP.t0 110.612
R3581 VP.n17 VP.t4 110.612
R3582 VP.n56 VP.t9 110.612
R3583 VP.n31 VP.t3 110.612
R3584 VP.n73 VP.n72 89.0887
R3585 VP.n126 VP.n0 89.0887
R3586 VP.n71 VP.n17 89.0887
R3587 VP.n31 VP.n30 74.5304
R3588 VP.n72 VP.n71 62.6849
R3589 VP.n80 VP.n79 41.9503
R3590 VP.n118 VP.n2 41.9503
R3591 VP.n63 VP.n19 41.9503
R3592 VP.n93 VP.n92 40.979
R3593 VP.n105 VP.n6 40.979
R3594 VP.n50 VP.n23 40.979
R3595 VP.n38 VP.n37 40.979
R3596 VP.n93 VP.n10 40.0078
R3597 VP.n105 VP.n104 40.0078
R3598 VP.n50 VP.n49 40.0078
R3599 VP.n38 VP.n27 40.0078
R3600 VP.n80 VP.n14 39.0365
R3601 VP.n118 VP.n117 39.0365
R3602 VP.n63 VP.n62 39.0365
R3603 VP.n74 VP.n16 24.4675
R3604 VP.n78 VP.n16 24.4675
R3605 VP.n79 VP.n78 24.4675
R3606 VP.n84 VP.n14 24.4675
R3607 VP.n85 VP.n84 24.4675
R3608 VP.n87 VP.n12 24.4675
R3609 VP.n91 VP.n12 24.4675
R3610 VP.n92 VP.n91 24.4675
R3611 VP.n97 VP.n10 24.4675
R3612 VP.n98 VP.n97 24.4675
R3613 VP.n99 VP.n98 24.4675
R3614 VP.n99 VP.n8 24.4675
R3615 VP.n103 VP.n8 24.4675
R3616 VP.n104 VP.n103 24.4675
R3617 VP.n109 VP.n6 24.4675
R3618 VP.n110 VP.n109 24.4675
R3619 VP.n112 VP.n110 24.4675
R3620 VP.n116 VP.n4 24.4675
R3621 VP.n117 VP.n116 24.4675
R3622 VP.n122 VP.n2 24.4675
R3623 VP.n123 VP.n122 24.4675
R3624 VP.n124 VP.n123 24.4675
R3625 VP.n67 VP.n19 24.4675
R3626 VP.n68 VP.n67 24.4675
R3627 VP.n69 VP.n68 24.4675
R3628 VP.n54 VP.n23 24.4675
R3629 VP.n55 VP.n54 24.4675
R3630 VP.n57 VP.n55 24.4675
R3631 VP.n61 VP.n21 24.4675
R3632 VP.n62 VP.n61 24.4675
R3633 VP.n42 VP.n27 24.4675
R3634 VP.n43 VP.n42 24.4675
R3635 VP.n44 VP.n43 24.4675
R3636 VP.n44 VP.n25 24.4675
R3637 VP.n48 VP.n25 24.4675
R3638 VP.n49 VP.n48 24.4675
R3639 VP.n32 VP.n29 24.4675
R3640 VP.n36 VP.n29 24.4675
R3641 VP.n37 VP.n36 24.4675
R3642 VP.n86 VP.n85 23.9782
R3643 VP.n111 VP.n4 23.9782
R3644 VP.n56 VP.n21 23.9782
R3645 VP.n33 VP.n30 3.44122
R3646 VP.n74 VP.n73 0.97918
R3647 VP.n124 VP.n0 0.97918
R3648 VP.n69 VP.n17 0.97918
R3649 VP.n87 VP.n86 0.48984
R3650 VP.n112 VP.n111 0.48984
R3651 VP.n57 VP.n56 0.48984
R3652 VP.n32 VP.n31 0.48984
R3653 VP.n71 VP.n70 0.354971
R3654 VP.n75 VP.n72 0.354971
R3655 VP.n126 VP.n125 0.354971
R3656 VP VP.n126 0.26696
R3657 VP.n34 VP.n33 0.189894
R3658 VP.n35 VP.n34 0.189894
R3659 VP.n35 VP.n28 0.189894
R3660 VP.n39 VP.n28 0.189894
R3661 VP.n40 VP.n39 0.189894
R3662 VP.n41 VP.n40 0.189894
R3663 VP.n41 VP.n26 0.189894
R3664 VP.n45 VP.n26 0.189894
R3665 VP.n46 VP.n45 0.189894
R3666 VP.n47 VP.n46 0.189894
R3667 VP.n47 VP.n24 0.189894
R3668 VP.n51 VP.n24 0.189894
R3669 VP.n52 VP.n51 0.189894
R3670 VP.n53 VP.n52 0.189894
R3671 VP.n53 VP.n22 0.189894
R3672 VP.n58 VP.n22 0.189894
R3673 VP.n59 VP.n58 0.189894
R3674 VP.n60 VP.n59 0.189894
R3675 VP.n60 VP.n20 0.189894
R3676 VP.n64 VP.n20 0.189894
R3677 VP.n65 VP.n64 0.189894
R3678 VP.n66 VP.n65 0.189894
R3679 VP.n66 VP.n18 0.189894
R3680 VP.n70 VP.n18 0.189894
R3681 VP.n76 VP.n75 0.189894
R3682 VP.n77 VP.n76 0.189894
R3683 VP.n77 VP.n15 0.189894
R3684 VP.n81 VP.n15 0.189894
R3685 VP.n82 VP.n81 0.189894
R3686 VP.n83 VP.n82 0.189894
R3687 VP.n83 VP.n13 0.189894
R3688 VP.n88 VP.n13 0.189894
R3689 VP.n89 VP.n88 0.189894
R3690 VP.n90 VP.n89 0.189894
R3691 VP.n90 VP.n11 0.189894
R3692 VP.n94 VP.n11 0.189894
R3693 VP.n95 VP.n94 0.189894
R3694 VP.n96 VP.n95 0.189894
R3695 VP.n96 VP.n9 0.189894
R3696 VP.n100 VP.n9 0.189894
R3697 VP.n101 VP.n100 0.189894
R3698 VP.n102 VP.n101 0.189894
R3699 VP.n102 VP.n7 0.189894
R3700 VP.n106 VP.n7 0.189894
R3701 VP.n107 VP.n106 0.189894
R3702 VP.n108 VP.n107 0.189894
R3703 VP.n108 VP.n5 0.189894
R3704 VP.n113 VP.n5 0.189894
R3705 VP.n114 VP.n113 0.189894
R3706 VP.n115 VP.n114 0.189894
R3707 VP.n115 VP.n3 0.189894
R3708 VP.n119 VP.n3 0.189894
R3709 VP.n120 VP.n119 0.189894
R3710 VP.n121 VP.n120 0.189894
R3711 VP.n121 VP.n1 0.189894
R3712 VP.n125 VP.n1 0.189894
R3713 VDD1.n88 VDD1.n0 289.615
R3714 VDD1.n183 VDD1.n95 289.615
R3715 VDD1.n89 VDD1.n88 185
R3716 VDD1.n87 VDD1.n86 185
R3717 VDD1.n4 VDD1.n3 185
R3718 VDD1.n81 VDD1.n80 185
R3719 VDD1.n79 VDD1.n78 185
R3720 VDD1.n77 VDD1.n7 185
R3721 VDD1.n11 VDD1.n8 185
R3722 VDD1.n72 VDD1.n71 185
R3723 VDD1.n70 VDD1.n69 185
R3724 VDD1.n13 VDD1.n12 185
R3725 VDD1.n64 VDD1.n63 185
R3726 VDD1.n62 VDD1.n61 185
R3727 VDD1.n17 VDD1.n16 185
R3728 VDD1.n56 VDD1.n55 185
R3729 VDD1.n54 VDD1.n53 185
R3730 VDD1.n21 VDD1.n20 185
R3731 VDD1.n48 VDD1.n47 185
R3732 VDD1.n46 VDD1.n45 185
R3733 VDD1.n25 VDD1.n24 185
R3734 VDD1.n40 VDD1.n39 185
R3735 VDD1.n38 VDD1.n37 185
R3736 VDD1.n29 VDD1.n28 185
R3737 VDD1.n32 VDD1.n31 185
R3738 VDD1.n126 VDD1.n125 185
R3739 VDD1.n123 VDD1.n122 185
R3740 VDD1.n132 VDD1.n131 185
R3741 VDD1.n134 VDD1.n133 185
R3742 VDD1.n119 VDD1.n118 185
R3743 VDD1.n140 VDD1.n139 185
R3744 VDD1.n142 VDD1.n141 185
R3745 VDD1.n115 VDD1.n114 185
R3746 VDD1.n148 VDD1.n147 185
R3747 VDD1.n150 VDD1.n149 185
R3748 VDD1.n111 VDD1.n110 185
R3749 VDD1.n156 VDD1.n155 185
R3750 VDD1.n158 VDD1.n157 185
R3751 VDD1.n107 VDD1.n106 185
R3752 VDD1.n164 VDD1.n163 185
R3753 VDD1.n167 VDD1.n166 185
R3754 VDD1.n165 VDD1.n103 185
R3755 VDD1.n172 VDD1.n102 185
R3756 VDD1.n174 VDD1.n173 185
R3757 VDD1.n176 VDD1.n175 185
R3758 VDD1.n99 VDD1.n98 185
R3759 VDD1.n182 VDD1.n181 185
R3760 VDD1.n184 VDD1.n183 185
R3761 VDD1.t4 VDD1.n30 147.659
R3762 VDD1.t2 VDD1.n124 147.659
R3763 VDD1.n88 VDD1.n87 104.615
R3764 VDD1.n87 VDD1.n3 104.615
R3765 VDD1.n80 VDD1.n3 104.615
R3766 VDD1.n80 VDD1.n79 104.615
R3767 VDD1.n79 VDD1.n7 104.615
R3768 VDD1.n11 VDD1.n7 104.615
R3769 VDD1.n71 VDD1.n11 104.615
R3770 VDD1.n71 VDD1.n70 104.615
R3771 VDD1.n70 VDD1.n12 104.615
R3772 VDD1.n63 VDD1.n12 104.615
R3773 VDD1.n63 VDD1.n62 104.615
R3774 VDD1.n62 VDD1.n16 104.615
R3775 VDD1.n55 VDD1.n16 104.615
R3776 VDD1.n55 VDD1.n54 104.615
R3777 VDD1.n54 VDD1.n20 104.615
R3778 VDD1.n47 VDD1.n20 104.615
R3779 VDD1.n47 VDD1.n46 104.615
R3780 VDD1.n46 VDD1.n24 104.615
R3781 VDD1.n39 VDD1.n24 104.615
R3782 VDD1.n39 VDD1.n38 104.615
R3783 VDD1.n38 VDD1.n28 104.615
R3784 VDD1.n31 VDD1.n28 104.615
R3785 VDD1.n125 VDD1.n122 104.615
R3786 VDD1.n132 VDD1.n122 104.615
R3787 VDD1.n133 VDD1.n132 104.615
R3788 VDD1.n133 VDD1.n118 104.615
R3789 VDD1.n140 VDD1.n118 104.615
R3790 VDD1.n141 VDD1.n140 104.615
R3791 VDD1.n141 VDD1.n114 104.615
R3792 VDD1.n148 VDD1.n114 104.615
R3793 VDD1.n149 VDD1.n148 104.615
R3794 VDD1.n149 VDD1.n110 104.615
R3795 VDD1.n156 VDD1.n110 104.615
R3796 VDD1.n157 VDD1.n156 104.615
R3797 VDD1.n157 VDD1.n106 104.615
R3798 VDD1.n164 VDD1.n106 104.615
R3799 VDD1.n166 VDD1.n164 104.615
R3800 VDD1.n166 VDD1.n165 104.615
R3801 VDD1.n165 VDD1.n102 104.615
R3802 VDD1.n174 VDD1.n102 104.615
R3803 VDD1.n175 VDD1.n174 104.615
R3804 VDD1.n175 VDD1.n98 104.615
R3805 VDD1.n182 VDD1.n98 104.615
R3806 VDD1.n183 VDD1.n182 104.615
R3807 VDD1.n191 VDD1.n190 65.0074
R3808 VDD1.n94 VDD1.n93 62.4703
R3809 VDD1.n193 VDD1.n192 62.4701
R3810 VDD1.n189 VDD1.n188 62.4701
R3811 VDD1.n193 VDD1.n191 57.0074
R3812 VDD1.n94 VDD1.n92 54.0665
R3813 VDD1.n189 VDD1.n187 54.0665
R3814 VDD1.n31 VDD1.t4 52.3082
R3815 VDD1.n125 VDD1.t2 52.3082
R3816 VDD1.n32 VDD1.n30 15.6677
R3817 VDD1.n126 VDD1.n124 15.6677
R3818 VDD1.n78 VDD1.n77 13.1884
R3819 VDD1.n173 VDD1.n172 13.1884
R3820 VDD1.n81 VDD1.n6 12.8005
R3821 VDD1.n76 VDD1.n8 12.8005
R3822 VDD1.n33 VDD1.n29 12.8005
R3823 VDD1.n127 VDD1.n123 12.8005
R3824 VDD1.n171 VDD1.n103 12.8005
R3825 VDD1.n176 VDD1.n101 12.8005
R3826 VDD1.n82 VDD1.n4 12.0247
R3827 VDD1.n73 VDD1.n72 12.0247
R3828 VDD1.n37 VDD1.n36 12.0247
R3829 VDD1.n131 VDD1.n130 12.0247
R3830 VDD1.n168 VDD1.n167 12.0247
R3831 VDD1.n177 VDD1.n99 12.0247
R3832 VDD1.n86 VDD1.n85 11.249
R3833 VDD1.n69 VDD1.n10 11.249
R3834 VDD1.n40 VDD1.n27 11.249
R3835 VDD1.n134 VDD1.n121 11.249
R3836 VDD1.n163 VDD1.n105 11.249
R3837 VDD1.n181 VDD1.n180 11.249
R3838 VDD1.n89 VDD1.n2 10.4732
R3839 VDD1.n68 VDD1.n13 10.4732
R3840 VDD1.n41 VDD1.n25 10.4732
R3841 VDD1.n135 VDD1.n119 10.4732
R3842 VDD1.n162 VDD1.n107 10.4732
R3843 VDD1.n184 VDD1.n97 10.4732
R3844 VDD1.n90 VDD1.n0 9.69747
R3845 VDD1.n65 VDD1.n64 9.69747
R3846 VDD1.n45 VDD1.n44 9.69747
R3847 VDD1.n139 VDD1.n138 9.69747
R3848 VDD1.n159 VDD1.n158 9.69747
R3849 VDD1.n185 VDD1.n95 9.69747
R3850 VDD1.n92 VDD1.n91 9.45567
R3851 VDD1.n187 VDD1.n186 9.45567
R3852 VDD1.n58 VDD1.n57 9.3005
R3853 VDD1.n60 VDD1.n59 9.3005
R3854 VDD1.n15 VDD1.n14 9.3005
R3855 VDD1.n66 VDD1.n65 9.3005
R3856 VDD1.n68 VDD1.n67 9.3005
R3857 VDD1.n10 VDD1.n9 9.3005
R3858 VDD1.n74 VDD1.n73 9.3005
R3859 VDD1.n76 VDD1.n75 9.3005
R3860 VDD1.n91 VDD1.n90 9.3005
R3861 VDD1.n2 VDD1.n1 9.3005
R3862 VDD1.n85 VDD1.n84 9.3005
R3863 VDD1.n83 VDD1.n82 9.3005
R3864 VDD1.n6 VDD1.n5 9.3005
R3865 VDD1.n19 VDD1.n18 9.3005
R3866 VDD1.n52 VDD1.n51 9.3005
R3867 VDD1.n50 VDD1.n49 9.3005
R3868 VDD1.n23 VDD1.n22 9.3005
R3869 VDD1.n44 VDD1.n43 9.3005
R3870 VDD1.n42 VDD1.n41 9.3005
R3871 VDD1.n27 VDD1.n26 9.3005
R3872 VDD1.n36 VDD1.n35 9.3005
R3873 VDD1.n34 VDD1.n33 9.3005
R3874 VDD1.n186 VDD1.n185 9.3005
R3875 VDD1.n97 VDD1.n96 9.3005
R3876 VDD1.n180 VDD1.n179 9.3005
R3877 VDD1.n178 VDD1.n177 9.3005
R3878 VDD1.n101 VDD1.n100 9.3005
R3879 VDD1.n146 VDD1.n145 9.3005
R3880 VDD1.n144 VDD1.n143 9.3005
R3881 VDD1.n117 VDD1.n116 9.3005
R3882 VDD1.n138 VDD1.n137 9.3005
R3883 VDD1.n136 VDD1.n135 9.3005
R3884 VDD1.n121 VDD1.n120 9.3005
R3885 VDD1.n130 VDD1.n129 9.3005
R3886 VDD1.n128 VDD1.n127 9.3005
R3887 VDD1.n113 VDD1.n112 9.3005
R3888 VDD1.n152 VDD1.n151 9.3005
R3889 VDD1.n154 VDD1.n153 9.3005
R3890 VDD1.n109 VDD1.n108 9.3005
R3891 VDD1.n160 VDD1.n159 9.3005
R3892 VDD1.n162 VDD1.n161 9.3005
R3893 VDD1.n105 VDD1.n104 9.3005
R3894 VDD1.n169 VDD1.n168 9.3005
R3895 VDD1.n171 VDD1.n170 9.3005
R3896 VDD1.n61 VDD1.n15 8.92171
R3897 VDD1.n48 VDD1.n23 8.92171
R3898 VDD1.n142 VDD1.n117 8.92171
R3899 VDD1.n155 VDD1.n109 8.92171
R3900 VDD1.n60 VDD1.n17 8.14595
R3901 VDD1.n49 VDD1.n21 8.14595
R3902 VDD1.n143 VDD1.n115 8.14595
R3903 VDD1.n154 VDD1.n111 8.14595
R3904 VDD1.n57 VDD1.n56 7.3702
R3905 VDD1.n53 VDD1.n52 7.3702
R3906 VDD1.n147 VDD1.n146 7.3702
R3907 VDD1.n151 VDD1.n150 7.3702
R3908 VDD1.n56 VDD1.n19 6.59444
R3909 VDD1.n53 VDD1.n19 6.59444
R3910 VDD1.n147 VDD1.n113 6.59444
R3911 VDD1.n150 VDD1.n113 6.59444
R3912 VDD1.n57 VDD1.n17 5.81868
R3913 VDD1.n52 VDD1.n21 5.81868
R3914 VDD1.n146 VDD1.n115 5.81868
R3915 VDD1.n151 VDD1.n111 5.81868
R3916 VDD1.n61 VDD1.n60 5.04292
R3917 VDD1.n49 VDD1.n48 5.04292
R3918 VDD1.n143 VDD1.n142 5.04292
R3919 VDD1.n155 VDD1.n154 5.04292
R3920 VDD1.n34 VDD1.n30 4.38563
R3921 VDD1.n128 VDD1.n124 4.38563
R3922 VDD1.n92 VDD1.n0 4.26717
R3923 VDD1.n64 VDD1.n15 4.26717
R3924 VDD1.n45 VDD1.n23 4.26717
R3925 VDD1.n139 VDD1.n117 4.26717
R3926 VDD1.n158 VDD1.n109 4.26717
R3927 VDD1.n187 VDD1.n95 4.26717
R3928 VDD1.n90 VDD1.n89 3.49141
R3929 VDD1.n65 VDD1.n13 3.49141
R3930 VDD1.n44 VDD1.n25 3.49141
R3931 VDD1.n138 VDD1.n119 3.49141
R3932 VDD1.n159 VDD1.n107 3.49141
R3933 VDD1.n185 VDD1.n184 3.49141
R3934 VDD1.n86 VDD1.n2 2.71565
R3935 VDD1.n69 VDD1.n68 2.71565
R3936 VDD1.n41 VDD1.n40 2.71565
R3937 VDD1.n135 VDD1.n134 2.71565
R3938 VDD1.n163 VDD1.n162 2.71565
R3939 VDD1.n181 VDD1.n97 2.71565
R3940 VDD1 VDD1.n193 2.53498
R3941 VDD1.n85 VDD1.n4 1.93989
R3942 VDD1.n72 VDD1.n10 1.93989
R3943 VDD1.n37 VDD1.n27 1.93989
R3944 VDD1.n131 VDD1.n121 1.93989
R3945 VDD1.n167 VDD1.n105 1.93989
R3946 VDD1.n180 VDD1.n99 1.93989
R3947 VDD1.n192 VDD1.t0 1.17279
R3948 VDD1.n192 VDD1.t5 1.17279
R3949 VDD1.n93 VDD1.t6 1.17279
R3950 VDD1.n93 VDD1.t9 1.17279
R3951 VDD1.n190 VDD1.t8 1.17279
R3952 VDD1.n190 VDD1.t3 1.17279
R3953 VDD1.n188 VDD1.t7 1.17279
R3954 VDD1.n188 VDD1.t1 1.17279
R3955 VDD1.n82 VDD1.n81 1.16414
R3956 VDD1.n73 VDD1.n8 1.16414
R3957 VDD1.n36 VDD1.n29 1.16414
R3958 VDD1.n130 VDD1.n123 1.16414
R3959 VDD1.n168 VDD1.n103 1.16414
R3960 VDD1.n177 VDD1.n176 1.16414
R3961 VDD1 VDD1.n94 0.922914
R3962 VDD1.n191 VDD1.n189 0.809378
R3963 VDD1.n78 VDD1.n6 0.388379
R3964 VDD1.n77 VDD1.n76 0.388379
R3965 VDD1.n33 VDD1.n32 0.388379
R3966 VDD1.n127 VDD1.n126 0.388379
R3967 VDD1.n172 VDD1.n171 0.388379
R3968 VDD1.n173 VDD1.n101 0.388379
R3969 VDD1.n91 VDD1.n1 0.155672
R3970 VDD1.n84 VDD1.n1 0.155672
R3971 VDD1.n84 VDD1.n83 0.155672
R3972 VDD1.n83 VDD1.n5 0.155672
R3973 VDD1.n75 VDD1.n5 0.155672
R3974 VDD1.n75 VDD1.n74 0.155672
R3975 VDD1.n74 VDD1.n9 0.155672
R3976 VDD1.n67 VDD1.n9 0.155672
R3977 VDD1.n67 VDD1.n66 0.155672
R3978 VDD1.n66 VDD1.n14 0.155672
R3979 VDD1.n59 VDD1.n14 0.155672
R3980 VDD1.n59 VDD1.n58 0.155672
R3981 VDD1.n58 VDD1.n18 0.155672
R3982 VDD1.n51 VDD1.n18 0.155672
R3983 VDD1.n51 VDD1.n50 0.155672
R3984 VDD1.n50 VDD1.n22 0.155672
R3985 VDD1.n43 VDD1.n22 0.155672
R3986 VDD1.n43 VDD1.n42 0.155672
R3987 VDD1.n42 VDD1.n26 0.155672
R3988 VDD1.n35 VDD1.n26 0.155672
R3989 VDD1.n35 VDD1.n34 0.155672
R3990 VDD1.n129 VDD1.n128 0.155672
R3991 VDD1.n129 VDD1.n120 0.155672
R3992 VDD1.n136 VDD1.n120 0.155672
R3993 VDD1.n137 VDD1.n136 0.155672
R3994 VDD1.n137 VDD1.n116 0.155672
R3995 VDD1.n144 VDD1.n116 0.155672
R3996 VDD1.n145 VDD1.n144 0.155672
R3997 VDD1.n145 VDD1.n112 0.155672
R3998 VDD1.n152 VDD1.n112 0.155672
R3999 VDD1.n153 VDD1.n152 0.155672
R4000 VDD1.n153 VDD1.n108 0.155672
R4001 VDD1.n160 VDD1.n108 0.155672
R4002 VDD1.n161 VDD1.n160 0.155672
R4003 VDD1.n161 VDD1.n104 0.155672
R4004 VDD1.n169 VDD1.n104 0.155672
R4005 VDD1.n170 VDD1.n169 0.155672
R4006 VDD1.n170 VDD1.n100 0.155672
R4007 VDD1.n178 VDD1.n100 0.155672
R4008 VDD1.n179 VDD1.n178 0.155672
R4009 VDD1.n179 VDD1.n96 0.155672
R4010 VDD1.n186 VDD1.n96 0.155672
C0 VTAIL VDD2 12.9028f
C1 VP VN 10.9005f
C2 VDD1 VP 16.283f
C3 VDD2 VP 0.720937f
C4 VDD1 VN 0.155441f
C5 VDD2 VN 15.721801f
C6 VTAIL VP 16.6079f
C7 VDD1 VDD2 2.87569f
C8 VTAIL VN 16.593199f
C9 VTAIL VDD1 12.8445f
C10 VDD2 B 9.295241f
C11 VDD1 B 9.288852f
C12 VTAIL B 10.995021f
C13 VN B 23.68013f
C14 VP B 22.226114f
C15 VDD1.n0 B 0.034227f
C16 VDD1.n1 B 0.024234f
C17 VDD1.n2 B 0.013022f
C18 VDD1.n3 B 0.03078f
C19 VDD1.n4 B 0.013788f
C20 VDD1.n5 B 0.024234f
C21 VDD1.n6 B 0.013022f
C22 VDD1.n7 B 0.03078f
C23 VDD1.n8 B 0.013788f
C24 VDD1.n9 B 0.024234f
C25 VDD1.n10 B 0.013022f
C26 VDD1.n11 B 0.03078f
C27 VDD1.n12 B 0.03078f
C28 VDD1.n13 B 0.013788f
C29 VDD1.n14 B 0.024234f
C30 VDD1.n15 B 0.013022f
C31 VDD1.n16 B 0.03078f
C32 VDD1.n17 B 0.013788f
C33 VDD1.n18 B 0.024234f
C34 VDD1.n19 B 0.013022f
C35 VDD1.n20 B 0.03078f
C36 VDD1.n21 B 0.013788f
C37 VDD1.n22 B 0.024234f
C38 VDD1.n23 B 0.013022f
C39 VDD1.n24 B 0.03078f
C40 VDD1.n25 B 0.013788f
C41 VDD1.n26 B 0.024234f
C42 VDD1.n27 B 0.013022f
C43 VDD1.n28 B 0.03078f
C44 VDD1.n29 B 0.013788f
C45 VDD1.n30 B 0.169544f
C46 VDD1.t4 B 0.05091f
C47 VDD1.n31 B 0.023085f
C48 VDD1.n32 B 0.018183f
C49 VDD1.n33 B 0.013022f
C50 VDD1.n34 B 1.78662f
C51 VDD1.n35 B 0.024234f
C52 VDD1.n36 B 0.013022f
C53 VDD1.n37 B 0.013788f
C54 VDD1.n38 B 0.03078f
C55 VDD1.n39 B 0.03078f
C56 VDD1.n40 B 0.013788f
C57 VDD1.n41 B 0.013022f
C58 VDD1.n42 B 0.024234f
C59 VDD1.n43 B 0.024234f
C60 VDD1.n44 B 0.013022f
C61 VDD1.n45 B 0.013788f
C62 VDD1.n46 B 0.03078f
C63 VDD1.n47 B 0.03078f
C64 VDD1.n48 B 0.013788f
C65 VDD1.n49 B 0.013022f
C66 VDD1.n50 B 0.024234f
C67 VDD1.n51 B 0.024234f
C68 VDD1.n52 B 0.013022f
C69 VDD1.n53 B 0.013788f
C70 VDD1.n54 B 0.03078f
C71 VDD1.n55 B 0.03078f
C72 VDD1.n56 B 0.013788f
C73 VDD1.n57 B 0.013022f
C74 VDD1.n58 B 0.024234f
C75 VDD1.n59 B 0.024234f
C76 VDD1.n60 B 0.013022f
C77 VDD1.n61 B 0.013788f
C78 VDD1.n62 B 0.03078f
C79 VDD1.n63 B 0.03078f
C80 VDD1.n64 B 0.013788f
C81 VDD1.n65 B 0.013022f
C82 VDD1.n66 B 0.024234f
C83 VDD1.n67 B 0.024234f
C84 VDD1.n68 B 0.013022f
C85 VDD1.n69 B 0.013788f
C86 VDD1.n70 B 0.03078f
C87 VDD1.n71 B 0.03078f
C88 VDD1.n72 B 0.013788f
C89 VDD1.n73 B 0.013022f
C90 VDD1.n74 B 0.024234f
C91 VDD1.n75 B 0.024234f
C92 VDD1.n76 B 0.013022f
C93 VDD1.n77 B 0.013405f
C94 VDD1.n78 B 0.013405f
C95 VDD1.n79 B 0.03078f
C96 VDD1.n80 B 0.03078f
C97 VDD1.n81 B 0.013788f
C98 VDD1.n82 B 0.013022f
C99 VDD1.n83 B 0.024234f
C100 VDD1.n84 B 0.024234f
C101 VDD1.n85 B 0.013022f
C102 VDD1.n86 B 0.013788f
C103 VDD1.n87 B 0.03078f
C104 VDD1.n88 B 0.066923f
C105 VDD1.n89 B 0.013788f
C106 VDD1.n90 B 0.013022f
C107 VDD1.n91 B 0.058996f
C108 VDD1.n92 B 0.074629f
C109 VDD1.t6 B 0.323453f
C110 VDD1.t9 B 0.323453f
C111 VDD1.n93 B 2.94087f
C112 VDD1.n94 B 0.838429f
C113 VDD1.n95 B 0.034227f
C114 VDD1.n96 B 0.024234f
C115 VDD1.n97 B 0.013022f
C116 VDD1.n98 B 0.03078f
C117 VDD1.n99 B 0.013788f
C118 VDD1.n100 B 0.024234f
C119 VDD1.n101 B 0.013022f
C120 VDD1.n102 B 0.03078f
C121 VDD1.n103 B 0.013788f
C122 VDD1.n104 B 0.024234f
C123 VDD1.n105 B 0.013022f
C124 VDD1.n106 B 0.03078f
C125 VDD1.n107 B 0.013788f
C126 VDD1.n108 B 0.024234f
C127 VDD1.n109 B 0.013022f
C128 VDD1.n110 B 0.03078f
C129 VDD1.n111 B 0.013788f
C130 VDD1.n112 B 0.024234f
C131 VDD1.n113 B 0.013022f
C132 VDD1.n114 B 0.03078f
C133 VDD1.n115 B 0.013788f
C134 VDD1.n116 B 0.024234f
C135 VDD1.n117 B 0.013022f
C136 VDD1.n118 B 0.03078f
C137 VDD1.n119 B 0.013788f
C138 VDD1.n120 B 0.024234f
C139 VDD1.n121 B 0.013022f
C140 VDD1.n122 B 0.03078f
C141 VDD1.n123 B 0.013788f
C142 VDD1.n124 B 0.169544f
C143 VDD1.t2 B 0.05091f
C144 VDD1.n125 B 0.023085f
C145 VDD1.n126 B 0.018183f
C146 VDD1.n127 B 0.013022f
C147 VDD1.n128 B 1.78662f
C148 VDD1.n129 B 0.024234f
C149 VDD1.n130 B 0.013022f
C150 VDD1.n131 B 0.013788f
C151 VDD1.n132 B 0.03078f
C152 VDD1.n133 B 0.03078f
C153 VDD1.n134 B 0.013788f
C154 VDD1.n135 B 0.013022f
C155 VDD1.n136 B 0.024234f
C156 VDD1.n137 B 0.024234f
C157 VDD1.n138 B 0.013022f
C158 VDD1.n139 B 0.013788f
C159 VDD1.n140 B 0.03078f
C160 VDD1.n141 B 0.03078f
C161 VDD1.n142 B 0.013788f
C162 VDD1.n143 B 0.013022f
C163 VDD1.n144 B 0.024234f
C164 VDD1.n145 B 0.024234f
C165 VDD1.n146 B 0.013022f
C166 VDD1.n147 B 0.013788f
C167 VDD1.n148 B 0.03078f
C168 VDD1.n149 B 0.03078f
C169 VDD1.n150 B 0.013788f
C170 VDD1.n151 B 0.013022f
C171 VDD1.n152 B 0.024234f
C172 VDD1.n153 B 0.024234f
C173 VDD1.n154 B 0.013022f
C174 VDD1.n155 B 0.013788f
C175 VDD1.n156 B 0.03078f
C176 VDD1.n157 B 0.03078f
C177 VDD1.n158 B 0.013788f
C178 VDD1.n159 B 0.013022f
C179 VDD1.n160 B 0.024234f
C180 VDD1.n161 B 0.024234f
C181 VDD1.n162 B 0.013022f
C182 VDD1.n163 B 0.013788f
C183 VDD1.n164 B 0.03078f
C184 VDD1.n165 B 0.03078f
C185 VDD1.n166 B 0.03078f
C186 VDD1.n167 B 0.013788f
C187 VDD1.n168 B 0.013022f
C188 VDD1.n169 B 0.024234f
C189 VDD1.n170 B 0.024234f
C190 VDD1.n171 B 0.013022f
C191 VDD1.n172 B 0.013405f
C192 VDD1.n173 B 0.013405f
C193 VDD1.n174 B 0.03078f
C194 VDD1.n175 B 0.03078f
C195 VDD1.n176 B 0.013788f
C196 VDD1.n177 B 0.013022f
C197 VDD1.n178 B 0.024234f
C198 VDD1.n179 B 0.024234f
C199 VDD1.n180 B 0.013022f
C200 VDD1.n181 B 0.013788f
C201 VDD1.n182 B 0.03078f
C202 VDD1.n183 B 0.066923f
C203 VDD1.n184 B 0.013788f
C204 VDD1.n185 B 0.013022f
C205 VDD1.n186 B 0.058996f
C206 VDD1.n187 B 0.074629f
C207 VDD1.t7 B 0.323453f
C208 VDD1.t1 B 0.323453f
C209 VDD1.n188 B 2.94086f
C210 VDD1.n189 B 0.830267f
C211 VDD1.t8 B 0.323453f
C212 VDD1.t3 B 0.323453f
C213 VDD1.n190 B 2.96727f
C214 VDD1.n191 B 3.81155f
C215 VDD1.t0 B 0.323453f
C216 VDD1.t5 B 0.323453f
C217 VDD1.n192 B 2.94086f
C218 VDD1.n193 B 3.86583f
C219 VP.t6 B 2.81766f
C220 VP.n0 B 1.03181f
C221 VP.n1 B 0.016502f
C222 VP.n2 B 0.032527f
C223 VP.n3 B 0.016502f
C224 VP.n4 B 0.030451f
C225 VP.n5 B 0.016502f
C226 VP.n6 B 0.032713f
C227 VP.n7 B 0.016502f
C228 VP.n8 B 0.030755f
C229 VP.n9 B 0.016502f
C230 VP.t8 B 2.81766f
C231 VP.n10 B 0.032878f
C232 VP.n11 B 0.016502f
C233 VP.n12 B 0.030755f
C234 VP.n13 B 0.016502f
C235 VP.t2 B 2.81766f
C236 VP.n14 B 0.033022f
C237 VP.n15 B 0.016502f
C238 VP.n16 B 0.030755f
C239 VP.t4 B 2.81766f
C240 VP.n17 B 1.03181f
C241 VP.n18 B 0.016502f
C242 VP.n19 B 0.032527f
C243 VP.n20 B 0.016502f
C244 VP.n21 B 0.030451f
C245 VP.n22 B 0.016502f
C246 VP.n23 B 0.032713f
C247 VP.n24 B 0.016502f
C248 VP.n25 B 0.030755f
C249 VP.n26 B 0.016502f
C250 VP.t0 B 2.81766f
C251 VP.n27 B 0.032878f
C252 VP.n28 B 0.016502f
C253 VP.n29 B 0.030755f
C254 VP.t5 B 3.06001f
C255 VP.n30 B 0.985776f
C256 VP.t3 B 2.81766f
C257 VP.n31 B 1.02535f
C258 VP.n32 B 0.015875f
C259 VP.n33 B 0.209586f
C260 VP.n34 B 0.016502f
C261 VP.n35 B 0.016502f
C262 VP.n36 B 0.030755f
C263 VP.n37 B 0.032713f
C264 VP.n38 B 0.013346f
C265 VP.n39 B 0.016502f
C266 VP.n40 B 0.016502f
C267 VP.n41 B 0.016502f
C268 VP.n42 B 0.030755f
C269 VP.n43 B 0.030755f
C270 VP.n44 B 0.988886f
C271 VP.n45 B 0.016502f
C272 VP.n46 B 0.016502f
C273 VP.n47 B 0.016502f
C274 VP.n48 B 0.030755f
C275 VP.n49 B 0.032878f
C276 VP.n50 B 0.013346f
C277 VP.n51 B 0.016502f
C278 VP.n52 B 0.016502f
C279 VP.n53 B 0.016502f
C280 VP.n54 B 0.030755f
C281 VP.n55 B 0.030755f
C282 VP.t9 B 2.81766f
C283 VP.n56 B 0.973315f
C284 VP.n57 B 0.015875f
C285 VP.n58 B 0.016502f
C286 VP.n59 B 0.016502f
C287 VP.n60 B 0.016502f
C288 VP.n61 B 0.030755f
C289 VP.n62 B 0.033022f
C290 VP.n63 B 0.013388f
C291 VP.n64 B 0.016502f
C292 VP.n65 B 0.016502f
C293 VP.n66 B 0.016502f
C294 VP.n67 B 0.030755f
C295 VP.n68 B 0.030755f
C296 VP.n69 B 0.016178f
C297 VP.n70 B 0.026633f
C298 VP.n71 B 1.2902f
C299 VP.n72 B 1.29967f
C300 VP.t7 B 2.81766f
C301 VP.n73 B 1.03181f
C302 VP.n74 B 0.016178f
C303 VP.n75 B 0.026633f
C304 VP.n76 B 0.016502f
C305 VP.n77 B 0.016502f
C306 VP.n78 B 0.030755f
C307 VP.n79 B 0.032527f
C308 VP.n80 B 0.013388f
C309 VP.n81 B 0.016502f
C310 VP.n82 B 0.016502f
C311 VP.n83 B 0.016502f
C312 VP.n84 B 0.030755f
C313 VP.n85 B 0.030451f
C314 VP.n86 B 0.973315f
C315 VP.n87 B 0.015875f
C316 VP.n88 B 0.016502f
C317 VP.n89 B 0.016502f
C318 VP.n90 B 0.016502f
C319 VP.n91 B 0.030755f
C320 VP.n92 B 0.032713f
C321 VP.n93 B 0.013346f
C322 VP.n94 B 0.016502f
C323 VP.n95 B 0.016502f
C324 VP.n96 B 0.016502f
C325 VP.n97 B 0.030755f
C326 VP.n98 B 0.030755f
C327 VP.n99 B 0.988886f
C328 VP.n100 B 0.016502f
C329 VP.n101 B 0.016502f
C330 VP.n102 B 0.016502f
C331 VP.n103 B 0.030755f
C332 VP.n104 B 0.032878f
C333 VP.n105 B 0.013346f
C334 VP.n106 B 0.016502f
C335 VP.n107 B 0.016502f
C336 VP.n108 B 0.016502f
C337 VP.n109 B 0.030755f
C338 VP.n110 B 0.030755f
C339 VP.t1 B 2.81766f
C340 VP.n111 B 0.973315f
C341 VP.n112 B 0.015875f
C342 VP.n113 B 0.016502f
C343 VP.n114 B 0.016502f
C344 VP.n115 B 0.016502f
C345 VP.n116 B 0.030755f
C346 VP.n117 B 0.033022f
C347 VP.n118 B 0.013388f
C348 VP.n119 B 0.016502f
C349 VP.n120 B 0.016502f
C350 VP.n121 B 0.016502f
C351 VP.n122 B 0.030755f
C352 VP.n123 B 0.030755f
C353 VP.n124 B 0.016178f
C354 VP.n125 B 0.026633f
C355 VP.n126 B 0.050445f
C356 VDD2.n0 B 0.033786f
C357 VDD2.n1 B 0.023922f
C358 VDD2.n2 B 0.012855f
C359 VDD2.n3 B 0.030384f
C360 VDD2.n4 B 0.013611f
C361 VDD2.n5 B 0.023922f
C362 VDD2.n6 B 0.012855f
C363 VDD2.n7 B 0.030384f
C364 VDD2.n8 B 0.013611f
C365 VDD2.n9 B 0.023922f
C366 VDD2.n10 B 0.012855f
C367 VDD2.n11 B 0.030384f
C368 VDD2.n12 B 0.013611f
C369 VDD2.n13 B 0.023922f
C370 VDD2.n14 B 0.012855f
C371 VDD2.n15 B 0.030384f
C372 VDD2.n16 B 0.013611f
C373 VDD2.n17 B 0.023922f
C374 VDD2.n18 B 0.012855f
C375 VDD2.n19 B 0.030384f
C376 VDD2.n20 B 0.013611f
C377 VDD2.n21 B 0.023922f
C378 VDD2.n22 B 0.012855f
C379 VDD2.n23 B 0.030384f
C380 VDD2.n24 B 0.013611f
C381 VDD2.n25 B 0.023922f
C382 VDD2.n26 B 0.012855f
C383 VDD2.n27 B 0.030384f
C384 VDD2.n28 B 0.013611f
C385 VDD2.n29 B 0.167363f
C386 VDD2.t1 B 0.050255f
C387 VDD2.n30 B 0.022788f
C388 VDD2.n31 B 0.017949f
C389 VDD2.n32 B 0.012855f
C390 VDD2.n33 B 1.76364f
C391 VDD2.n34 B 0.023922f
C392 VDD2.n35 B 0.012855f
C393 VDD2.n36 B 0.013611f
C394 VDD2.n37 B 0.030384f
C395 VDD2.n38 B 0.030384f
C396 VDD2.n39 B 0.013611f
C397 VDD2.n40 B 0.012855f
C398 VDD2.n41 B 0.023922f
C399 VDD2.n42 B 0.023922f
C400 VDD2.n43 B 0.012855f
C401 VDD2.n44 B 0.013611f
C402 VDD2.n45 B 0.030384f
C403 VDD2.n46 B 0.030384f
C404 VDD2.n47 B 0.013611f
C405 VDD2.n48 B 0.012855f
C406 VDD2.n49 B 0.023922f
C407 VDD2.n50 B 0.023922f
C408 VDD2.n51 B 0.012855f
C409 VDD2.n52 B 0.013611f
C410 VDD2.n53 B 0.030384f
C411 VDD2.n54 B 0.030384f
C412 VDD2.n55 B 0.013611f
C413 VDD2.n56 B 0.012855f
C414 VDD2.n57 B 0.023922f
C415 VDD2.n58 B 0.023922f
C416 VDD2.n59 B 0.012855f
C417 VDD2.n60 B 0.013611f
C418 VDD2.n61 B 0.030384f
C419 VDD2.n62 B 0.030384f
C420 VDD2.n63 B 0.013611f
C421 VDD2.n64 B 0.012855f
C422 VDD2.n65 B 0.023922f
C423 VDD2.n66 B 0.023922f
C424 VDD2.n67 B 0.012855f
C425 VDD2.n68 B 0.013611f
C426 VDD2.n69 B 0.030384f
C427 VDD2.n70 B 0.030384f
C428 VDD2.n71 B 0.030384f
C429 VDD2.n72 B 0.013611f
C430 VDD2.n73 B 0.012855f
C431 VDD2.n74 B 0.023922f
C432 VDD2.n75 B 0.023922f
C433 VDD2.n76 B 0.012855f
C434 VDD2.n77 B 0.013233f
C435 VDD2.n78 B 0.013233f
C436 VDD2.n79 B 0.030384f
C437 VDD2.n80 B 0.030384f
C438 VDD2.n81 B 0.013611f
C439 VDD2.n82 B 0.012855f
C440 VDD2.n83 B 0.023922f
C441 VDD2.n84 B 0.023922f
C442 VDD2.n85 B 0.012855f
C443 VDD2.n86 B 0.013611f
C444 VDD2.n87 B 0.030384f
C445 VDD2.n88 B 0.066062f
C446 VDD2.n89 B 0.013611f
C447 VDD2.n90 B 0.012855f
C448 VDD2.n91 B 0.058237f
C449 VDD2.n92 B 0.073668f
C450 VDD2.t6 B 0.319292f
C451 VDD2.t2 B 0.319292f
C452 VDD2.n93 B 2.90303f
C453 VDD2.n94 B 0.819587f
C454 VDD2.t7 B 0.319292f
C455 VDD2.t0 B 0.319292f
C456 VDD2.n95 B 2.9291f
C457 VDD2.n96 B 3.61103f
C458 VDD2.n97 B 0.033786f
C459 VDD2.n98 B 0.023922f
C460 VDD2.n99 B 0.012855f
C461 VDD2.n100 B 0.030384f
C462 VDD2.n101 B 0.013611f
C463 VDD2.n102 B 0.023922f
C464 VDD2.n103 B 0.012855f
C465 VDD2.n104 B 0.030384f
C466 VDD2.n105 B 0.013611f
C467 VDD2.n106 B 0.023922f
C468 VDD2.n107 B 0.012855f
C469 VDD2.n108 B 0.030384f
C470 VDD2.n109 B 0.030384f
C471 VDD2.n110 B 0.013611f
C472 VDD2.n111 B 0.023922f
C473 VDD2.n112 B 0.012855f
C474 VDD2.n113 B 0.030384f
C475 VDD2.n114 B 0.013611f
C476 VDD2.n115 B 0.023922f
C477 VDD2.n116 B 0.012855f
C478 VDD2.n117 B 0.030384f
C479 VDD2.n118 B 0.013611f
C480 VDD2.n119 B 0.023922f
C481 VDD2.n120 B 0.012855f
C482 VDD2.n121 B 0.030384f
C483 VDD2.n122 B 0.013611f
C484 VDD2.n123 B 0.023922f
C485 VDD2.n124 B 0.012855f
C486 VDD2.n125 B 0.030384f
C487 VDD2.n126 B 0.013611f
C488 VDD2.n127 B 0.167363f
C489 VDD2.t9 B 0.050255f
C490 VDD2.n128 B 0.022788f
C491 VDD2.n129 B 0.017949f
C492 VDD2.n130 B 0.012855f
C493 VDD2.n131 B 1.76364f
C494 VDD2.n132 B 0.023922f
C495 VDD2.n133 B 0.012855f
C496 VDD2.n134 B 0.013611f
C497 VDD2.n135 B 0.030384f
C498 VDD2.n136 B 0.030384f
C499 VDD2.n137 B 0.013611f
C500 VDD2.n138 B 0.012855f
C501 VDD2.n139 B 0.023922f
C502 VDD2.n140 B 0.023922f
C503 VDD2.n141 B 0.012855f
C504 VDD2.n142 B 0.013611f
C505 VDD2.n143 B 0.030384f
C506 VDD2.n144 B 0.030384f
C507 VDD2.n145 B 0.013611f
C508 VDD2.n146 B 0.012855f
C509 VDD2.n147 B 0.023922f
C510 VDD2.n148 B 0.023922f
C511 VDD2.n149 B 0.012855f
C512 VDD2.n150 B 0.013611f
C513 VDD2.n151 B 0.030384f
C514 VDD2.n152 B 0.030384f
C515 VDD2.n153 B 0.013611f
C516 VDD2.n154 B 0.012855f
C517 VDD2.n155 B 0.023922f
C518 VDD2.n156 B 0.023922f
C519 VDD2.n157 B 0.012855f
C520 VDD2.n158 B 0.013611f
C521 VDD2.n159 B 0.030384f
C522 VDD2.n160 B 0.030384f
C523 VDD2.n161 B 0.013611f
C524 VDD2.n162 B 0.012855f
C525 VDD2.n163 B 0.023922f
C526 VDD2.n164 B 0.023922f
C527 VDD2.n165 B 0.012855f
C528 VDD2.n166 B 0.013611f
C529 VDD2.n167 B 0.030384f
C530 VDD2.n168 B 0.030384f
C531 VDD2.n169 B 0.013611f
C532 VDD2.n170 B 0.012855f
C533 VDD2.n171 B 0.023922f
C534 VDD2.n172 B 0.023922f
C535 VDD2.n173 B 0.012855f
C536 VDD2.n174 B 0.013233f
C537 VDD2.n175 B 0.013233f
C538 VDD2.n176 B 0.030384f
C539 VDD2.n177 B 0.030384f
C540 VDD2.n178 B 0.013611f
C541 VDD2.n179 B 0.012855f
C542 VDD2.n180 B 0.023922f
C543 VDD2.n181 B 0.023922f
C544 VDD2.n182 B 0.012855f
C545 VDD2.n183 B 0.013611f
C546 VDD2.n184 B 0.030384f
C547 VDD2.n185 B 0.066062f
C548 VDD2.n186 B 0.013611f
C549 VDD2.n187 B 0.012855f
C550 VDD2.n188 B 0.058237f
C551 VDD2.n189 B 0.053578f
C552 VDD2.n190 B 3.52602f
C553 VDD2.t8 B 0.319292f
C554 VDD2.t3 B 0.319292f
C555 VDD2.n191 B 2.90304f
C556 VDD2.n192 B 0.533517f
C557 VDD2.t5 B 0.319292f
C558 VDD2.t4 B 0.319292f
C559 VDD2.n193 B 2.92905f
C560 VTAIL.t13 B 0.325826f
C561 VTAIL.t12 B 0.325826f
C562 VTAIL.n0 B 2.89129f
C563 VTAIL.n1 B 0.619362f
C564 VTAIL.n2 B 0.034478f
C565 VTAIL.n3 B 0.024412f
C566 VTAIL.n4 B 0.013118f
C567 VTAIL.n5 B 0.031006f
C568 VTAIL.n6 B 0.01389f
C569 VTAIL.n7 B 0.024412f
C570 VTAIL.n8 B 0.013118f
C571 VTAIL.n9 B 0.031006f
C572 VTAIL.n10 B 0.01389f
C573 VTAIL.n11 B 0.024412f
C574 VTAIL.n12 B 0.013118f
C575 VTAIL.n13 B 0.031006f
C576 VTAIL.n14 B 0.01389f
C577 VTAIL.n15 B 0.024412f
C578 VTAIL.n16 B 0.013118f
C579 VTAIL.n17 B 0.031006f
C580 VTAIL.n18 B 0.01389f
C581 VTAIL.n19 B 0.024412f
C582 VTAIL.n20 B 0.013118f
C583 VTAIL.n21 B 0.031006f
C584 VTAIL.n22 B 0.01389f
C585 VTAIL.n23 B 0.024412f
C586 VTAIL.n24 B 0.013118f
C587 VTAIL.n25 B 0.031006f
C588 VTAIL.n26 B 0.01389f
C589 VTAIL.n27 B 0.024412f
C590 VTAIL.n28 B 0.013118f
C591 VTAIL.n29 B 0.031006f
C592 VTAIL.n30 B 0.01389f
C593 VTAIL.n31 B 0.170788f
C594 VTAIL.t1 B 0.051283f
C595 VTAIL.n32 B 0.023254f
C596 VTAIL.n33 B 0.018316f
C597 VTAIL.n34 B 0.013118f
C598 VTAIL.n35 B 1.79973f
C599 VTAIL.n36 B 0.024412f
C600 VTAIL.n37 B 0.013118f
C601 VTAIL.n38 B 0.01389f
C602 VTAIL.n39 B 0.031006f
C603 VTAIL.n40 B 0.031006f
C604 VTAIL.n41 B 0.01389f
C605 VTAIL.n42 B 0.013118f
C606 VTAIL.n43 B 0.024412f
C607 VTAIL.n44 B 0.024412f
C608 VTAIL.n45 B 0.013118f
C609 VTAIL.n46 B 0.01389f
C610 VTAIL.n47 B 0.031006f
C611 VTAIL.n48 B 0.031006f
C612 VTAIL.n49 B 0.01389f
C613 VTAIL.n50 B 0.013118f
C614 VTAIL.n51 B 0.024412f
C615 VTAIL.n52 B 0.024412f
C616 VTAIL.n53 B 0.013118f
C617 VTAIL.n54 B 0.01389f
C618 VTAIL.n55 B 0.031006f
C619 VTAIL.n56 B 0.031006f
C620 VTAIL.n57 B 0.01389f
C621 VTAIL.n58 B 0.013118f
C622 VTAIL.n59 B 0.024412f
C623 VTAIL.n60 B 0.024412f
C624 VTAIL.n61 B 0.013118f
C625 VTAIL.n62 B 0.01389f
C626 VTAIL.n63 B 0.031006f
C627 VTAIL.n64 B 0.031006f
C628 VTAIL.n65 B 0.01389f
C629 VTAIL.n66 B 0.013118f
C630 VTAIL.n67 B 0.024412f
C631 VTAIL.n68 B 0.024412f
C632 VTAIL.n69 B 0.013118f
C633 VTAIL.n70 B 0.01389f
C634 VTAIL.n71 B 0.031006f
C635 VTAIL.n72 B 0.031006f
C636 VTAIL.n73 B 0.031006f
C637 VTAIL.n74 B 0.01389f
C638 VTAIL.n75 B 0.013118f
C639 VTAIL.n76 B 0.024412f
C640 VTAIL.n77 B 0.024412f
C641 VTAIL.n78 B 0.013118f
C642 VTAIL.n79 B 0.013504f
C643 VTAIL.n80 B 0.013504f
C644 VTAIL.n81 B 0.031006f
C645 VTAIL.n82 B 0.031006f
C646 VTAIL.n83 B 0.01389f
C647 VTAIL.n84 B 0.013118f
C648 VTAIL.n85 B 0.024412f
C649 VTAIL.n86 B 0.024412f
C650 VTAIL.n87 B 0.013118f
C651 VTAIL.n88 B 0.01389f
C652 VTAIL.n89 B 0.031006f
C653 VTAIL.n90 B 0.067414f
C654 VTAIL.n91 B 0.01389f
C655 VTAIL.n92 B 0.013118f
C656 VTAIL.n93 B 0.059428f
C657 VTAIL.n94 B 0.037841f
C658 VTAIL.n95 B 0.467386f
C659 VTAIL.t5 B 0.325826f
C660 VTAIL.t6 B 0.325826f
C661 VTAIL.n96 B 2.89129f
C662 VTAIL.n97 B 0.781769f
C663 VTAIL.t0 B 0.325826f
C664 VTAIL.t17 B 0.325826f
C665 VTAIL.n98 B 2.89129f
C666 VTAIL.n99 B 2.53063f
C667 VTAIL.t11 B 0.325826f
C668 VTAIL.t7 B 0.325826f
C669 VTAIL.n100 B 2.89131f
C670 VTAIL.n101 B 2.53061f
C671 VTAIL.t15 B 0.325826f
C672 VTAIL.t8 B 0.325826f
C673 VTAIL.n102 B 2.89131f
C674 VTAIL.n103 B 0.781756f
C675 VTAIL.n104 B 0.034478f
C676 VTAIL.n105 B 0.024412f
C677 VTAIL.n106 B 0.013118f
C678 VTAIL.n107 B 0.031006f
C679 VTAIL.n108 B 0.01389f
C680 VTAIL.n109 B 0.024412f
C681 VTAIL.n110 B 0.013118f
C682 VTAIL.n111 B 0.031006f
C683 VTAIL.n112 B 0.01389f
C684 VTAIL.n113 B 0.024412f
C685 VTAIL.n114 B 0.013118f
C686 VTAIL.n115 B 0.031006f
C687 VTAIL.n116 B 0.031006f
C688 VTAIL.n117 B 0.01389f
C689 VTAIL.n118 B 0.024412f
C690 VTAIL.n119 B 0.013118f
C691 VTAIL.n120 B 0.031006f
C692 VTAIL.n121 B 0.01389f
C693 VTAIL.n122 B 0.024412f
C694 VTAIL.n123 B 0.013118f
C695 VTAIL.n124 B 0.031006f
C696 VTAIL.n125 B 0.01389f
C697 VTAIL.n126 B 0.024412f
C698 VTAIL.n127 B 0.013118f
C699 VTAIL.n128 B 0.031006f
C700 VTAIL.n129 B 0.01389f
C701 VTAIL.n130 B 0.024412f
C702 VTAIL.n131 B 0.013118f
C703 VTAIL.n132 B 0.031006f
C704 VTAIL.n133 B 0.01389f
C705 VTAIL.n134 B 0.170788f
C706 VTAIL.t10 B 0.051283f
C707 VTAIL.n135 B 0.023254f
C708 VTAIL.n136 B 0.018316f
C709 VTAIL.n137 B 0.013118f
C710 VTAIL.n138 B 1.79973f
C711 VTAIL.n139 B 0.024412f
C712 VTAIL.n140 B 0.013118f
C713 VTAIL.n141 B 0.01389f
C714 VTAIL.n142 B 0.031006f
C715 VTAIL.n143 B 0.031006f
C716 VTAIL.n144 B 0.01389f
C717 VTAIL.n145 B 0.013118f
C718 VTAIL.n146 B 0.024412f
C719 VTAIL.n147 B 0.024412f
C720 VTAIL.n148 B 0.013118f
C721 VTAIL.n149 B 0.01389f
C722 VTAIL.n150 B 0.031006f
C723 VTAIL.n151 B 0.031006f
C724 VTAIL.n152 B 0.01389f
C725 VTAIL.n153 B 0.013118f
C726 VTAIL.n154 B 0.024412f
C727 VTAIL.n155 B 0.024412f
C728 VTAIL.n156 B 0.013118f
C729 VTAIL.n157 B 0.01389f
C730 VTAIL.n158 B 0.031006f
C731 VTAIL.n159 B 0.031006f
C732 VTAIL.n160 B 0.01389f
C733 VTAIL.n161 B 0.013118f
C734 VTAIL.n162 B 0.024412f
C735 VTAIL.n163 B 0.024412f
C736 VTAIL.n164 B 0.013118f
C737 VTAIL.n165 B 0.01389f
C738 VTAIL.n166 B 0.031006f
C739 VTAIL.n167 B 0.031006f
C740 VTAIL.n168 B 0.01389f
C741 VTAIL.n169 B 0.013118f
C742 VTAIL.n170 B 0.024412f
C743 VTAIL.n171 B 0.024412f
C744 VTAIL.n172 B 0.013118f
C745 VTAIL.n173 B 0.01389f
C746 VTAIL.n174 B 0.031006f
C747 VTAIL.n175 B 0.031006f
C748 VTAIL.n176 B 0.01389f
C749 VTAIL.n177 B 0.013118f
C750 VTAIL.n178 B 0.024412f
C751 VTAIL.n179 B 0.024412f
C752 VTAIL.n180 B 0.013118f
C753 VTAIL.n181 B 0.013504f
C754 VTAIL.n182 B 0.013504f
C755 VTAIL.n183 B 0.031006f
C756 VTAIL.n184 B 0.031006f
C757 VTAIL.n185 B 0.01389f
C758 VTAIL.n186 B 0.013118f
C759 VTAIL.n187 B 0.024412f
C760 VTAIL.n188 B 0.024412f
C761 VTAIL.n189 B 0.013118f
C762 VTAIL.n190 B 0.01389f
C763 VTAIL.n191 B 0.031006f
C764 VTAIL.n192 B 0.067414f
C765 VTAIL.n193 B 0.01389f
C766 VTAIL.n194 B 0.013118f
C767 VTAIL.n195 B 0.059428f
C768 VTAIL.n196 B 0.037841f
C769 VTAIL.n197 B 0.467386f
C770 VTAIL.t2 B 0.325826f
C771 VTAIL.t4 B 0.325826f
C772 VTAIL.n198 B 2.89131f
C773 VTAIL.n199 B 0.682752f
C774 VTAIL.t3 B 0.325826f
C775 VTAIL.t18 B 0.325826f
C776 VTAIL.n200 B 2.89131f
C777 VTAIL.n201 B 0.781756f
C778 VTAIL.n202 B 0.034478f
C779 VTAIL.n203 B 0.024412f
C780 VTAIL.n204 B 0.013118f
C781 VTAIL.n205 B 0.031006f
C782 VTAIL.n206 B 0.01389f
C783 VTAIL.n207 B 0.024412f
C784 VTAIL.n208 B 0.013118f
C785 VTAIL.n209 B 0.031006f
C786 VTAIL.n210 B 0.01389f
C787 VTAIL.n211 B 0.024412f
C788 VTAIL.n212 B 0.013118f
C789 VTAIL.n213 B 0.031006f
C790 VTAIL.n214 B 0.031006f
C791 VTAIL.n215 B 0.01389f
C792 VTAIL.n216 B 0.024412f
C793 VTAIL.n217 B 0.013118f
C794 VTAIL.n218 B 0.031006f
C795 VTAIL.n219 B 0.01389f
C796 VTAIL.n220 B 0.024412f
C797 VTAIL.n221 B 0.013118f
C798 VTAIL.n222 B 0.031006f
C799 VTAIL.n223 B 0.01389f
C800 VTAIL.n224 B 0.024412f
C801 VTAIL.n225 B 0.013118f
C802 VTAIL.n226 B 0.031006f
C803 VTAIL.n227 B 0.01389f
C804 VTAIL.n228 B 0.024412f
C805 VTAIL.n229 B 0.013118f
C806 VTAIL.n230 B 0.031006f
C807 VTAIL.n231 B 0.01389f
C808 VTAIL.n232 B 0.170788f
C809 VTAIL.t19 B 0.051283f
C810 VTAIL.n233 B 0.023254f
C811 VTAIL.n234 B 0.018316f
C812 VTAIL.n235 B 0.013118f
C813 VTAIL.n236 B 1.79973f
C814 VTAIL.n237 B 0.024412f
C815 VTAIL.n238 B 0.013118f
C816 VTAIL.n239 B 0.01389f
C817 VTAIL.n240 B 0.031006f
C818 VTAIL.n241 B 0.031006f
C819 VTAIL.n242 B 0.01389f
C820 VTAIL.n243 B 0.013118f
C821 VTAIL.n244 B 0.024412f
C822 VTAIL.n245 B 0.024412f
C823 VTAIL.n246 B 0.013118f
C824 VTAIL.n247 B 0.01389f
C825 VTAIL.n248 B 0.031006f
C826 VTAIL.n249 B 0.031006f
C827 VTAIL.n250 B 0.01389f
C828 VTAIL.n251 B 0.013118f
C829 VTAIL.n252 B 0.024412f
C830 VTAIL.n253 B 0.024412f
C831 VTAIL.n254 B 0.013118f
C832 VTAIL.n255 B 0.01389f
C833 VTAIL.n256 B 0.031006f
C834 VTAIL.n257 B 0.031006f
C835 VTAIL.n258 B 0.01389f
C836 VTAIL.n259 B 0.013118f
C837 VTAIL.n260 B 0.024412f
C838 VTAIL.n261 B 0.024412f
C839 VTAIL.n262 B 0.013118f
C840 VTAIL.n263 B 0.01389f
C841 VTAIL.n264 B 0.031006f
C842 VTAIL.n265 B 0.031006f
C843 VTAIL.n266 B 0.01389f
C844 VTAIL.n267 B 0.013118f
C845 VTAIL.n268 B 0.024412f
C846 VTAIL.n269 B 0.024412f
C847 VTAIL.n270 B 0.013118f
C848 VTAIL.n271 B 0.01389f
C849 VTAIL.n272 B 0.031006f
C850 VTAIL.n273 B 0.031006f
C851 VTAIL.n274 B 0.01389f
C852 VTAIL.n275 B 0.013118f
C853 VTAIL.n276 B 0.024412f
C854 VTAIL.n277 B 0.024412f
C855 VTAIL.n278 B 0.013118f
C856 VTAIL.n279 B 0.013504f
C857 VTAIL.n280 B 0.013504f
C858 VTAIL.n281 B 0.031006f
C859 VTAIL.n282 B 0.031006f
C860 VTAIL.n283 B 0.01389f
C861 VTAIL.n284 B 0.013118f
C862 VTAIL.n285 B 0.024412f
C863 VTAIL.n286 B 0.024412f
C864 VTAIL.n287 B 0.013118f
C865 VTAIL.n288 B 0.01389f
C866 VTAIL.n289 B 0.031006f
C867 VTAIL.n290 B 0.067414f
C868 VTAIL.n291 B 0.01389f
C869 VTAIL.n292 B 0.013118f
C870 VTAIL.n293 B 0.059428f
C871 VTAIL.n294 B 0.037841f
C872 VTAIL.n295 B 2.04332f
C873 VTAIL.n296 B 0.034478f
C874 VTAIL.n297 B 0.024412f
C875 VTAIL.n298 B 0.013118f
C876 VTAIL.n299 B 0.031006f
C877 VTAIL.n300 B 0.01389f
C878 VTAIL.n301 B 0.024412f
C879 VTAIL.n302 B 0.013118f
C880 VTAIL.n303 B 0.031006f
C881 VTAIL.n304 B 0.01389f
C882 VTAIL.n305 B 0.024412f
C883 VTAIL.n306 B 0.013118f
C884 VTAIL.n307 B 0.031006f
C885 VTAIL.n308 B 0.01389f
C886 VTAIL.n309 B 0.024412f
C887 VTAIL.n310 B 0.013118f
C888 VTAIL.n311 B 0.031006f
C889 VTAIL.n312 B 0.01389f
C890 VTAIL.n313 B 0.024412f
C891 VTAIL.n314 B 0.013118f
C892 VTAIL.n315 B 0.031006f
C893 VTAIL.n316 B 0.01389f
C894 VTAIL.n317 B 0.024412f
C895 VTAIL.n318 B 0.013118f
C896 VTAIL.n319 B 0.031006f
C897 VTAIL.n320 B 0.01389f
C898 VTAIL.n321 B 0.024412f
C899 VTAIL.n322 B 0.013118f
C900 VTAIL.n323 B 0.031006f
C901 VTAIL.n324 B 0.01389f
C902 VTAIL.n325 B 0.170788f
C903 VTAIL.t16 B 0.051283f
C904 VTAIL.n326 B 0.023254f
C905 VTAIL.n327 B 0.018316f
C906 VTAIL.n328 B 0.013118f
C907 VTAIL.n329 B 1.79973f
C908 VTAIL.n330 B 0.024412f
C909 VTAIL.n331 B 0.013118f
C910 VTAIL.n332 B 0.01389f
C911 VTAIL.n333 B 0.031006f
C912 VTAIL.n334 B 0.031006f
C913 VTAIL.n335 B 0.01389f
C914 VTAIL.n336 B 0.013118f
C915 VTAIL.n337 B 0.024412f
C916 VTAIL.n338 B 0.024412f
C917 VTAIL.n339 B 0.013118f
C918 VTAIL.n340 B 0.01389f
C919 VTAIL.n341 B 0.031006f
C920 VTAIL.n342 B 0.031006f
C921 VTAIL.n343 B 0.01389f
C922 VTAIL.n344 B 0.013118f
C923 VTAIL.n345 B 0.024412f
C924 VTAIL.n346 B 0.024412f
C925 VTAIL.n347 B 0.013118f
C926 VTAIL.n348 B 0.01389f
C927 VTAIL.n349 B 0.031006f
C928 VTAIL.n350 B 0.031006f
C929 VTAIL.n351 B 0.01389f
C930 VTAIL.n352 B 0.013118f
C931 VTAIL.n353 B 0.024412f
C932 VTAIL.n354 B 0.024412f
C933 VTAIL.n355 B 0.013118f
C934 VTAIL.n356 B 0.01389f
C935 VTAIL.n357 B 0.031006f
C936 VTAIL.n358 B 0.031006f
C937 VTAIL.n359 B 0.01389f
C938 VTAIL.n360 B 0.013118f
C939 VTAIL.n361 B 0.024412f
C940 VTAIL.n362 B 0.024412f
C941 VTAIL.n363 B 0.013118f
C942 VTAIL.n364 B 0.01389f
C943 VTAIL.n365 B 0.031006f
C944 VTAIL.n366 B 0.031006f
C945 VTAIL.n367 B 0.031006f
C946 VTAIL.n368 B 0.01389f
C947 VTAIL.n369 B 0.013118f
C948 VTAIL.n370 B 0.024412f
C949 VTAIL.n371 B 0.024412f
C950 VTAIL.n372 B 0.013118f
C951 VTAIL.n373 B 0.013504f
C952 VTAIL.n374 B 0.013504f
C953 VTAIL.n375 B 0.031006f
C954 VTAIL.n376 B 0.031006f
C955 VTAIL.n377 B 0.01389f
C956 VTAIL.n378 B 0.013118f
C957 VTAIL.n379 B 0.024412f
C958 VTAIL.n380 B 0.024412f
C959 VTAIL.n381 B 0.013118f
C960 VTAIL.n382 B 0.01389f
C961 VTAIL.n383 B 0.031006f
C962 VTAIL.n384 B 0.067414f
C963 VTAIL.n385 B 0.01389f
C964 VTAIL.n386 B 0.013118f
C965 VTAIL.n387 B 0.059428f
C966 VTAIL.n388 B 0.037841f
C967 VTAIL.n389 B 2.04332f
C968 VTAIL.t14 B 0.325826f
C969 VTAIL.t9 B 0.325826f
C970 VTAIL.n390 B 2.89129f
C971 VTAIL.n391 B 0.57325f
C972 VN.t9 B 2.7776f
C973 VN.n0 B 1.01713f
C974 VN.n1 B 0.016267f
C975 VN.n2 B 0.032064f
C976 VN.n3 B 0.016267f
C977 VN.n4 B 0.030018f
C978 VN.n5 B 0.016267f
C979 VN.n6 B 0.032248f
C980 VN.n7 B 0.016267f
C981 VN.n8 B 0.030318f
C982 VN.n9 B 0.016267f
C983 VN.t7 B 2.7776f
C984 VN.n10 B 0.032411f
C985 VN.n11 B 0.016267f
C986 VN.n12 B 0.030318f
C987 VN.t8 B 3.0165f
C988 VN.n13 B 0.971757f
C989 VN.t3 B 2.7776f
C990 VN.n14 B 1.01077f
C991 VN.n15 B 0.015649f
C992 VN.n16 B 0.206605f
C993 VN.n17 B 0.016267f
C994 VN.n18 B 0.016267f
C995 VN.n19 B 0.030318f
C996 VN.n20 B 0.032248f
C997 VN.n21 B 0.013156f
C998 VN.n22 B 0.016267f
C999 VN.n23 B 0.016267f
C1000 VN.n24 B 0.016267f
C1001 VN.n25 B 0.030318f
C1002 VN.n26 B 0.030318f
C1003 VN.n27 B 0.974823f
C1004 VN.n28 B 0.016267f
C1005 VN.n29 B 0.016267f
C1006 VN.n30 B 0.016267f
C1007 VN.n31 B 0.030318f
C1008 VN.n32 B 0.032411f
C1009 VN.n33 B 0.013156f
C1010 VN.n34 B 0.016267f
C1011 VN.n35 B 0.016267f
C1012 VN.n36 B 0.016267f
C1013 VN.n37 B 0.030318f
C1014 VN.n38 B 0.030318f
C1015 VN.t2 B 2.7776f
C1016 VN.n39 B 0.959474f
C1017 VN.n40 B 0.015649f
C1018 VN.n41 B 0.016267f
C1019 VN.n42 B 0.016267f
C1020 VN.n43 B 0.016267f
C1021 VN.n44 B 0.030318f
C1022 VN.n45 B 0.032552f
C1023 VN.n46 B 0.013198f
C1024 VN.n47 B 0.016267f
C1025 VN.n48 B 0.016267f
C1026 VN.n49 B 0.016267f
C1027 VN.n50 B 0.030318f
C1028 VN.n51 B 0.030318f
C1029 VN.n52 B 0.015948f
C1030 VN.n53 B 0.026255f
C1031 VN.n54 B 0.049728f
C1032 VN.t0 B 2.7776f
C1033 VN.n55 B 1.01713f
C1034 VN.n56 B 0.016267f
C1035 VN.n57 B 0.032064f
C1036 VN.n58 B 0.016267f
C1037 VN.n59 B 0.030018f
C1038 VN.n60 B 0.016267f
C1039 VN.t1 B 2.7776f
C1040 VN.n61 B 0.959474f
C1041 VN.n62 B 0.032248f
C1042 VN.n63 B 0.016267f
C1043 VN.n64 B 0.030318f
C1044 VN.n65 B 0.016267f
C1045 VN.t6 B 2.7776f
C1046 VN.n66 B 0.032411f
C1047 VN.n67 B 0.016267f
C1048 VN.n68 B 0.030318f
C1049 VN.t5 B 3.0165f
C1050 VN.n69 B 0.971757f
C1051 VN.t4 B 2.7776f
C1052 VN.n70 B 1.01077f
C1053 VN.n71 B 0.015649f
C1054 VN.n72 B 0.206605f
C1055 VN.n73 B 0.016267f
C1056 VN.n74 B 0.016267f
C1057 VN.n75 B 0.030318f
C1058 VN.n76 B 0.032248f
C1059 VN.n77 B 0.013156f
C1060 VN.n78 B 0.016267f
C1061 VN.n79 B 0.016267f
C1062 VN.n80 B 0.016267f
C1063 VN.n81 B 0.030318f
C1064 VN.n82 B 0.030318f
C1065 VN.n83 B 0.974823f
C1066 VN.n84 B 0.016267f
C1067 VN.n85 B 0.016267f
C1068 VN.n86 B 0.016267f
C1069 VN.n87 B 0.030318f
C1070 VN.n88 B 0.032411f
C1071 VN.n89 B 0.013156f
C1072 VN.n90 B 0.016267f
C1073 VN.n91 B 0.016267f
C1074 VN.n92 B 0.016267f
C1075 VN.n93 B 0.030318f
C1076 VN.n94 B 0.030318f
C1077 VN.n95 B 0.015649f
C1078 VN.n96 B 0.016267f
C1079 VN.n97 B 0.016267f
C1080 VN.n98 B 0.016267f
C1081 VN.n99 B 0.030318f
C1082 VN.n100 B 0.032552f
C1083 VN.n101 B 0.013198f
C1084 VN.n102 B 0.016267f
C1085 VN.n103 B 0.016267f
C1086 VN.n104 B 0.016267f
C1087 VN.n105 B 0.030318f
C1088 VN.n106 B 0.030318f
C1089 VN.n107 B 0.015948f
C1090 VN.n108 B 0.026255f
C1091 VN.n109 B 1.27805f
.ends

