* NGSPICE file created from diff_pair_sample_1704.ext - technology: sky130A

.subckt diff_pair_sample_1704 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X1 VTAIL.t14 VN.t1 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=1.11375 ps=7.08 w=6.75 l=1.18
X2 VTAIL.t13 VN.t2 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X3 VTAIL.t12 VN.t3 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=1.11375 ps=7.08 w=6.75 l=1.18
X4 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=0 ps=0 w=6.75 l=1.18
X5 VTAIL.t0 VP.t0 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X6 VDD2.t6 VN.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=2.6325 ps=14.28 w=6.75 l=1.18
X7 VDD2.t4 VN.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X8 VTAIL.t1 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=1.11375 ps=7.08 w=6.75 l=1.18
X9 VDD1.t5 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=2.6325 ps=14.28 w=6.75 l=1.18
X10 VDD1.t4 VP.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=2.6325 ps=14.28 w=6.75 l=1.18
X11 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=0 ps=0 w=6.75 l=1.18
X12 VDD2.t3 VN.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X13 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X14 VDD2.t2 VN.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=2.6325 ps=14.28 w=6.75 l=1.18
X15 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=1.11375 ps=7.08 w=6.75 l=1.18
X16 VDD1.t1 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X17 VDD1.t0 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.11375 pd=7.08 as=1.11375 ps=7.08 w=6.75 l=1.18
X18 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=0 ps=0 w=6.75 l=1.18
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6325 pd=14.28 as=0 ps=0 w=6.75 l=1.18
R0 VN.n16 VN.n15 172.799
R1 VN.n33 VN.n32 172.799
R2 VN.n4 VN.t1 168.466
R3 VN.n22 VN.t7 168.466
R4 VN.n31 VN.n17 161.3
R5 VN.n30 VN.n29 161.3
R6 VN.n28 VN.n18 161.3
R7 VN.n27 VN.n26 161.3
R8 VN.n25 VN.n19 161.3
R9 VN.n24 VN.n23 161.3
R10 VN.n14 VN.n0 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n11 VN.n1 161.3
R13 VN.n10 VN.n9 161.3
R14 VN.n7 VN.n2 161.3
R15 VN.n6 VN.n5 161.3
R16 VN.n3 VN.t5 137.861
R17 VN.n8 VN.t0 137.861
R18 VN.n15 VN.t4 137.861
R19 VN.n21 VN.t2 137.861
R20 VN.n20 VN.t6 137.861
R21 VN.n32 VN.t3 137.861
R22 VN.n4 VN.n3 51.0708
R23 VN.n22 VN.n21 51.0708
R24 VN.n14 VN.n13 41.4647
R25 VN.n31 VN.n30 41.4647
R26 VN VN.n33 40.5478
R27 VN.n7 VN.n6 40.4934
R28 VN.n9 VN.n7 40.4934
R29 VN.n25 VN.n24 40.4934
R30 VN.n26 VN.n25 40.4934
R31 VN.n13 VN.n1 39.5221
R32 VN.n30 VN.n18 39.5221
R33 VN.n23 VN.n22 26.8925
R34 VN.n5 VN.n4 26.8925
R35 VN.n15 VN.n14 12.968
R36 VN.n32 VN.n31 12.968
R37 VN.n6 VN.n3 12.4787
R38 VN.n9 VN.n8 12.4787
R39 VN.n24 VN.n21 12.4787
R40 VN.n26 VN.n20 12.4787
R41 VN.n8 VN.n1 11.9893
R42 VN.n20 VN.n18 11.9893
R43 VN.n33 VN.n17 0.189894
R44 VN.n29 VN.n17 0.189894
R45 VN.n29 VN.n28 0.189894
R46 VN.n28 VN.n27 0.189894
R47 VN.n27 VN.n19 0.189894
R48 VN.n23 VN.n19 0.189894
R49 VN.n5 VN.n2 0.189894
R50 VN.n10 VN.n2 0.189894
R51 VN.n11 VN.n10 0.189894
R52 VN.n12 VN.n11 0.189894
R53 VN.n12 VN.n0 0.189894
R54 VN.n16 VN.n0 0.189894
R55 VN VN.n16 0.0516364
R56 VDD2.n2 VDD2.n1 67.2513
R57 VDD2.n2 VDD2.n0 67.2513
R58 VDD2 VDD2.n5 67.2484
R59 VDD2.n4 VDD2.n3 66.6559
R60 VDD2.n4 VDD2.n2 35.392
R61 VDD2.n5 VDD2.t1 2.93383
R62 VDD2.n5 VDD2.t2 2.93383
R63 VDD2.n3 VDD2.t5 2.93383
R64 VDD2.n3 VDD2.t3 2.93383
R65 VDD2.n1 VDD2.t0 2.93383
R66 VDD2.n1 VDD2.t6 2.93383
R67 VDD2.n0 VDD2.t7 2.93383
R68 VDD2.n0 VDD2.t4 2.93383
R69 VDD2 VDD2.n4 0.709552
R70 VTAIL.n290 VTAIL.n260 289.615
R71 VTAIL.n32 VTAIL.n2 289.615
R72 VTAIL.n68 VTAIL.n38 289.615
R73 VTAIL.n106 VTAIL.n76 289.615
R74 VTAIL.n254 VTAIL.n224 289.615
R75 VTAIL.n216 VTAIL.n186 289.615
R76 VTAIL.n180 VTAIL.n150 289.615
R77 VTAIL.n142 VTAIL.n112 289.615
R78 VTAIL.n273 VTAIL.n272 185
R79 VTAIL.n275 VTAIL.n274 185
R80 VTAIL.n268 VTAIL.n267 185
R81 VTAIL.n281 VTAIL.n280 185
R82 VTAIL.n283 VTAIL.n282 185
R83 VTAIL.n264 VTAIL.n263 185
R84 VTAIL.n289 VTAIL.n288 185
R85 VTAIL.n291 VTAIL.n290 185
R86 VTAIL.n15 VTAIL.n14 185
R87 VTAIL.n17 VTAIL.n16 185
R88 VTAIL.n10 VTAIL.n9 185
R89 VTAIL.n23 VTAIL.n22 185
R90 VTAIL.n25 VTAIL.n24 185
R91 VTAIL.n6 VTAIL.n5 185
R92 VTAIL.n31 VTAIL.n30 185
R93 VTAIL.n33 VTAIL.n32 185
R94 VTAIL.n51 VTAIL.n50 185
R95 VTAIL.n53 VTAIL.n52 185
R96 VTAIL.n46 VTAIL.n45 185
R97 VTAIL.n59 VTAIL.n58 185
R98 VTAIL.n61 VTAIL.n60 185
R99 VTAIL.n42 VTAIL.n41 185
R100 VTAIL.n67 VTAIL.n66 185
R101 VTAIL.n69 VTAIL.n68 185
R102 VTAIL.n89 VTAIL.n88 185
R103 VTAIL.n91 VTAIL.n90 185
R104 VTAIL.n84 VTAIL.n83 185
R105 VTAIL.n97 VTAIL.n96 185
R106 VTAIL.n99 VTAIL.n98 185
R107 VTAIL.n80 VTAIL.n79 185
R108 VTAIL.n105 VTAIL.n104 185
R109 VTAIL.n107 VTAIL.n106 185
R110 VTAIL.n255 VTAIL.n254 185
R111 VTAIL.n253 VTAIL.n252 185
R112 VTAIL.n228 VTAIL.n227 185
R113 VTAIL.n247 VTAIL.n246 185
R114 VTAIL.n245 VTAIL.n244 185
R115 VTAIL.n232 VTAIL.n231 185
R116 VTAIL.n239 VTAIL.n238 185
R117 VTAIL.n237 VTAIL.n236 185
R118 VTAIL.n217 VTAIL.n216 185
R119 VTAIL.n215 VTAIL.n214 185
R120 VTAIL.n190 VTAIL.n189 185
R121 VTAIL.n209 VTAIL.n208 185
R122 VTAIL.n207 VTAIL.n206 185
R123 VTAIL.n194 VTAIL.n193 185
R124 VTAIL.n201 VTAIL.n200 185
R125 VTAIL.n199 VTAIL.n198 185
R126 VTAIL.n181 VTAIL.n180 185
R127 VTAIL.n179 VTAIL.n178 185
R128 VTAIL.n154 VTAIL.n153 185
R129 VTAIL.n173 VTAIL.n172 185
R130 VTAIL.n171 VTAIL.n170 185
R131 VTAIL.n158 VTAIL.n157 185
R132 VTAIL.n165 VTAIL.n164 185
R133 VTAIL.n163 VTAIL.n162 185
R134 VTAIL.n143 VTAIL.n142 185
R135 VTAIL.n141 VTAIL.n140 185
R136 VTAIL.n116 VTAIL.n115 185
R137 VTAIL.n135 VTAIL.n134 185
R138 VTAIL.n133 VTAIL.n132 185
R139 VTAIL.n120 VTAIL.n119 185
R140 VTAIL.n127 VTAIL.n126 185
R141 VTAIL.n125 VTAIL.n124 185
R142 VTAIL.n271 VTAIL.t11 147.659
R143 VTAIL.n13 VTAIL.t14 147.659
R144 VTAIL.n49 VTAIL.t5 147.659
R145 VTAIL.n87 VTAIL.t4 147.659
R146 VTAIL.n235 VTAIL.t7 147.659
R147 VTAIL.n197 VTAIL.t1 147.659
R148 VTAIL.n161 VTAIL.t8 147.659
R149 VTAIL.n123 VTAIL.t12 147.659
R150 VTAIL.n274 VTAIL.n273 104.615
R151 VTAIL.n274 VTAIL.n267 104.615
R152 VTAIL.n281 VTAIL.n267 104.615
R153 VTAIL.n282 VTAIL.n281 104.615
R154 VTAIL.n282 VTAIL.n263 104.615
R155 VTAIL.n289 VTAIL.n263 104.615
R156 VTAIL.n290 VTAIL.n289 104.615
R157 VTAIL.n16 VTAIL.n15 104.615
R158 VTAIL.n16 VTAIL.n9 104.615
R159 VTAIL.n23 VTAIL.n9 104.615
R160 VTAIL.n24 VTAIL.n23 104.615
R161 VTAIL.n24 VTAIL.n5 104.615
R162 VTAIL.n31 VTAIL.n5 104.615
R163 VTAIL.n32 VTAIL.n31 104.615
R164 VTAIL.n52 VTAIL.n51 104.615
R165 VTAIL.n52 VTAIL.n45 104.615
R166 VTAIL.n59 VTAIL.n45 104.615
R167 VTAIL.n60 VTAIL.n59 104.615
R168 VTAIL.n60 VTAIL.n41 104.615
R169 VTAIL.n67 VTAIL.n41 104.615
R170 VTAIL.n68 VTAIL.n67 104.615
R171 VTAIL.n90 VTAIL.n89 104.615
R172 VTAIL.n90 VTAIL.n83 104.615
R173 VTAIL.n97 VTAIL.n83 104.615
R174 VTAIL.n98 VTAIL.n97 104.615
R175 VTAIL.n98 VTAIL.n79 104.615
R176 VTAIL.n105 VTAIL.n79 104.615
R177 VTAIL.n106 VTAIL.n105 104.615
R178 VTAIL.n254 VTAIL.n253 104.615
R179 VTAIL.n253 VTAIL.n227 104.615
R180 VTAIL.n246 VTAIL.n227 104.615
R181 VTAIL.n246 VTAIL.n245 104.615
R182 VTAIL.n245 VTAIL.n231 104.615
R183 VTAIL.n238 VTAIL.n231 104.615
R184 VTAIL.n238 VTAIL.n237 104.615
R185 VTAIL.n216 VTAIL.n215 104.615
R186 VTAIL.n215 VTAIL.n189 104.615
R187 VTAIL.n208 VTAIL.n189 104.615
R188 VTAIL.n208 VTAIL.n207 104.615
R189 VTAIL.n207 VTAIL.n193 104.615
R190 VTAIL.n200 VTAIL.n193 104.615
R191 VTAIL.n200 VTAIL.n199 104.615
R192 VTAIL.n180 VTAIL.n179 104.615
R193 VTAIL.n179 VTAIL.n153 104.615
R194 VTAIL.n172 VTAIL.n153 104.615
R195 VTAIL.n172 VTAIL.n171 104.615
R196 VTAIL.n171 VTAIL.n157 104.615
R197 VTAIL.n164 VTAIL.n157 104.615
R198 VTAIL.n164 VTAIL.n163 104.615
R199 VTAIL.n142 VTAIL.n141 104.615
R200 VTAIL.n141 VTAIL.n115 104.615
R201 VTAIL.n134 VTAIL.n115 104.615
R202 VTAIL.n134 VTAIL.n133 104.615
R203 VTAIL.n133 VTAIL.n119 104.615
R204 VTAIL.n126 VTAIL.n119 104.615
R205 VTAIL.n126 VTAIL.n125 104.615
R206 VTAIL.n273 VTAIL.t11 52.3082
R207 VTAIL.n15 VTAIL.t14 52.3082
R208 VTAIL.n51 VTAIL.t5 52.3082
R209 VTAIL.n89 VTAIL.t4 52.3082
R210 VTAIL.n237 VTAIL.t7 52.3082
R211 VTAIL.n199 VTAIL.t1 52.3082
R212 VTAIL.n163 VTAIL.t8 52.3082
R213 VTAIL.n125 VTAIL.t12 52.3082
R214 VTAIL.n223 VTAIL.n222 49.9772
R215 VTAIL.n149 VTAIL.n148 49.9772
R216 VTAIL.n1 VTAIL.n0 49.977
R217 VTAIL.n75 VTAIL.n74 49.977
R218 VTAIL.n295 VTAIL.n294 32.7672
R219 VTAIL.n37 VTAIL.n36 32.7672
R220 VTAIL.n73 VTAIL.n72 32.7672
R221 VTAIL.n111 VTAIL.n110 32.7672
R222 VTAIL.n259 VTAIL.n258 32.7672
R223 VTAIL.n221 VTAIL.n220 32.7672
R224 VTAIL.n185 VTAIL.n184 32.7672
R225 VTAIL.n147 VTAIL.n146 32.7672
R226 VTAIL.n295 VTAIL.n259 19.4876
R227 VTAIL.n147 VTAIL.n111 19.4876
R228 VTAIL.n272 VTAIL.n271 15.6676
R229 VTAIL.n14 VTAIL.n13 15.6676
R230 VTAIL.n50 VTAIL.n49 15.6676
R231 VTAIL.n88 VTAIL.n87 15.6676
R232 VTAIL.n236 VTAIL.n235 15.6676
R233 VTAIL.n198 VTAIL.n197 15.6676
R234 VTAIL.n162 VTAIL.n161 15.6676
R235 VTAIL.n124 VTAIL.n123 15.6676
R236 VTAIL.n275 VTAIL.n270 12.8005
R237 VTAIL.n17 VTAIL.n12 12.8005
R238 VTAIL.n53 VTAIL.n48 12.8005
R239 VTAIL.n91 VTAIL.n86 12.8005
R240 VTAIL.n239 VTAIL.n234 12.8005
R241 VTAIL.n201 VTAIL.n196 12.8005
R242 VTAIL.n165 VTAIL.n160 12.8005
R243 VTAIL.n127 VTAIL.n122 12.8005
R244 VTAIL.n276 VTAIL.n268 12.0247
R245 VTAIL.n18 VTAIL.n10 12.0247
R246 VTAIL.n54 VTAIL.n46 12.0247
R247 VTAIL.n92 VTAIL.n84 12.0247
R248 VTAIL.n240 VTAIL.n232 12.0247
R249 VTAIL.n202 VTAIL.n194 12.0247
R250 VTAIL.n166 VTAIL.n158 12.0247
R251 VTAIL.n128 VTAIL.n120 12.0247
R252 VTAIL.n280 VTAIL.n279 11.249
R253 VTAIL.n22 VTAIL.n21 11.249
R254 VTAIL.n58 VTAIL.n57 11.249
R255 VTAIL.n96 VTAIL.n95 11.249
R256 VTAIL.n244 VTAIL.n243 11.249
R257 VTAIL.n206 VTAIL.n205 11.249
R258 VTAIL.n170 VTAIL.n169 11.249
R259 VTAIL.n132 VTAIL.n131 11.249
R260 VTAIL.n283 VTAIL.n266 10.4732
R261 VTAIL.n25 VTAIL.n8 10.4732
R262 VTAIL.n61 VTAIL.n44 10.4732
R263 VTAIL.n99 VTAIL.n82 10.4732
R264 VTAIL.n247 VTAIL.n230 10.4732
R265 VTAIL.n209 VTAIL.n192 10.4732
R266 VTAIL.n173 VTAIL.n156 10.4732
R267 VTAIL.n135 VTAIL.n118 10.4732
R268 VTAIL.n284 VTAIL.n264 9.69747
R269 VTAIL.n26 VTAIL.n6 9.69747
R270 VTAIL.n62 VTAIL.n42 9.69747
R271 VTAIL.n100 VTAIL.n80 9.69747
R272 VTAIL.n248 VTAIL.n228 9.69747
R273 VTAIL.n210 VTAIL.n190 9.69747
R274 VTAIL.n174 VTAIL.n154 9.69747
R275 VTAIL.n136 VTAIL.n116 9.69747
R276 VTAIL.n294 VTAIL.n293 9.45567
R277 VTAIL.n36 VTAIL.n35 9.45567
R278 VTAIL.n72 VTAIL.n71 9.45567
R279 VTAIL.n110 VTAIL.n109 9.45567
R280 VTAIL.n258 VTAIL.n257 9.45567
R281 VTAIL.n220 VTAIL.n219 9.45567
R282 VTAIL.n184 VTAIL.n183 9.45567
R283 VTAIL.n146 VTAIL.n145 9.45567
R284 VTAIL.n262 VTAIL.n261 9.3005
R285 VTAIL.n287 VTAIL.n286 9.3005
R286 VTAIL.n285 VTAIL.n284 9.3005
R287 VTAIL.n266 VTAIL.n265 9.3005
R288 VTAIL.n279 VTAIL.n278 9.3005
R289 VTAIL.n277 VTAIL.n276 9.3005
R290 VTAIL.n270 VTAIL.n269 9.3005
R291 VTAIL.n293 VTAIL.n292 9.3005
R292 VTAIL.n4 VTAIL.n3 9.3005
R293 VTAIL.n29 VTAIL.n28 9.3005
R294 VTAIL.n27 VTAIL.n26 9.3005
R295 VTAIL.n8 VTAIL.n7 9.3005
R296 VTAIL.n21 VTAIL.n20 9.3005
R297 VTAIL.n19 VTAIL.n18 9.3005
R298 VTAIL.n12 VTAIL.n11 9.3005
R299 VTAIL.n35 VTAIL.n34 9.3005
R300 VTAIL.n40 VTAIL.n39 9.3005
R301 VTAIL.n65 VTAIL.n64 9.3005
R302 VTAIL.n63 VTAIL.n62 9.3005
R303 VTAIL.n44 VTAIL.n43 9.3005
R304 VTAIL.n57 VTAIL.n56 9.3005
R305 VTAIL.n55 VTAIL.n54 9.3005
R306 VTAIL.n48 VTAIL.n47 9.3005
R307 VTAIL.n71 VTAIL.n70 9.3005
R308 VTAIL.n78 VTAIL.n77 9.3005
R309 VTAIL.n103 VTAIL.n102 9.3005
R310 VTAIL.n101 VTAIL.n100 9.3005
R311 VTAIL.n82 VTAIL.n81 9.3005
R312 VTAIL.n95 VTAIL.n94 9.3005
R313 VTAIL.n93 VTAIL.n92 9.3005
R314 VTAIL.n86 VTAIL.n85 9.3005
R315 VTAIL.n109 VTAIL.n108 9.3005
R316 VTAIL.n257 VTAIL.n256 9.3005
R317 VTAIL.n226 VTAIL.n225 9.3005
R318 VTAIL.n251 VTAIL.n250 9.3005
R319 VTAIL.n249 VTAIL.n248 9.3005
R320 VTAIL.n230 VTAIL.n229 9.3005
R321 VTAIL.n243 VTAIL.n242 9.3005
R322 VTAIL.n241 VTAIL.n240 9.3005
R323 VTAIL.n234 VTAIL.n233 9.3005
R324 VTAIL.n219 VTAIL.n218 9.3005
R325 VTAIL.n188 VTAIL.n187 9.3005
R326 VTAIL.n213 VTAIL.n212 9.3005
R327 VTAIL.n211 VTAIL.n210 9.3005
R328 VTAIL.n192 VTAIL.n191 9.3005
R329 VTAIL.n205 VTAIL.n204 9.3005
R330 VTAIL.n203 VTAIL.n202 9.3005
R331 VTAIL.n196 VTAIL.n195 9.3005
R332 VTAIL.n183 VTAIL.n182 9.3005
R333 VTAIL.n152 VTAIL.n151 9.3005
R334 VTAIL.n177 VTAIL.n176 9.3005
R335 VTAIL.n175 VTAIL.n174 9.3005
R336 VTAIL.n156 VTAIL.n155 9.3005
R337 VTAIL.n169 VTAIL.n168 9.3005
R338 VTAIL.n167 VTAIL.n166 9.3005
R339 VTAIL.n160 VTAIL.n159 9.3005
R340 VTAIL.n145 VTAIL.n144 9.3005
R341 VTAIL.n114 VTAIL.n113 9.3005
R342 VTAIL.n139 VTAIL.n138 9.3005
R343 VTAIL.n137 VTAIL.n136 9.3005
R344 VTAIL.n118 VTAIL.n117 9.3005
R345 VTAIL.n131 VTAIL.n130 9.3005
R346 VTAIL.n129 VTAIL.n128 9.3005
R347 VTAIL.n122 VTAIL.n121 9.3005
R348 VTAIL.n288 VTAIL.n287 8.92171
R349 VTAIL.n30 VTAIL.n29 8.92171
R350 VTAIL.n66 VTAIL.n65 8.92171
R351 VTAIL.n104 VTAIL.n103 8.92171
R352 VTAIL.n252 VTAIL.n251 8.92171
R353 VTAIL.n214 VTAIL.n213 8.92171
R354 VTAIL.n178 VTAIL.n177 8.92171
R355 VTAIL.n140 VTAIL.n139 8.92171
R356 VTAIL.n291 VTAIL.n262 8.14595
R357 VTAIL.n33 VTAIL.n4 8.14595
R358 VTAIL.n69 VTAIL.n40 8.14595
R359 VTAIL.n107 VTAIL.n78 8.14595
R360 VTAIL.n255 VTAIL.n226 8.14595
R361 VTAIL.n217 VTAIL.n188 8.14595
R362 VTAIL.n181 VTAIL.n152 8.14595
R363 VTAIL.n143 VTAIL.n114 8.14595
R364 VTAIL.n292 VTAIL.n260 7.3702
R365 VTAIL.n34 VTAIL.n2 7.3702
R366 VTAIL.n70 VTAIL.n38 7.3702
R367 VTAIL.n108 VTAIL.n76 7.3702
R368 VTAIL.n256 VTAIL.n224 7.3702
R369 VTAIL.n218 VTAIL.n186 7.3702
R370 VTAIL.n182 VTAIL.n150 7.3702
R371 VTAIL.n144 VTAIL.n112 7.3702
R372 VTAIL.n294 VTAIL.n260 6.59444
R373 VTAIL.n36 VTAIL.n2 6.59444
R374 VTAIL.n72 VTAIL.n38 6.59444
R375 VTAIL.n110 VTAIL.n76 6.59444
R376 VTAIL.n258 VTAIL.n224 6.59444
R377 VTAIL.n220 VTAIL.n186 6.59444
R378 VTAIL.n184 VTAIL.n150 6.59444
R379 VTAIL.n146 VTAIL.n112 6.59444
R380 VTAIL.n292 VTAIL.n291 5.81868
R381 VTAIL.n34 VTAIL.n33 5.81868
R382 VTAIL.n70 VTAIL.n69 5.81868
R383 VTAIL.n108 VTAIL.n107 5.81868
R384 VTAIL.n256 VTAIL.n255 5.81868
R385 VTAIL.n218 VTAIL.n217 5.81868
R386 VTAIL.n182 VTAIL.n181 5.81868
R387 VTAIL.n144 VTAIL.n143 5.81868
R388 VTAIL.n288 VTAIL.n262 5.04292
R389 VTAIL.n30 VTAIL.n4 5.04292
R390 VTAIL.n66 VTAIL.n40 5.04292
R391 VTAIL.n104 VTAIL.n78 5.04292
R392 VTAIL.n252 VTAIL.n226 5.04292
R393 VTAIL.n214 VTAIL.n188 5.04292
R394 VTAIL.n178 VTAIL.n152 5.04292
R395 VTAIL.n140 VTAIL.n114 5.04292
R396 VTAIL.n271 VTAIL.n269 4.38571
R397 VTAIL.n13 VTAIL.n11 4.38571
R398 VTAIL.n49 VTAIL.n47 4.38571
R399 VTAIL.n87 VTAIL.n85 4.38571
R400 VTAIL.n235 VTAIL.n233 4.38571
R401 VTAIL.n197 VTAIL.n195 4.38571
R402 VTAIL.n161 VTAIL.n159 4.38571
R403 VTAIL.n123 VTAIL.n121 4.38571
R404 VTAIL.n287 VTAIL.n264 4.26717
R405 VTAIL.n29 VTAIL.n6 4.26717
R406 VTAIL.n65 VTAIL.n42 4.26717
R407 VTAIL.n103 VTAIL.n80 4.26717
R408 VTAIL.n251 VTAIL.n228 4.26717
R409 VTAIL.n213 VTAIL.n190 4.26717
R410 VTAIL.n177 VTAIL.n154 4.26717
R411 VTAIL.n139 VTAIL.n116 4.26717
R412 VTAIL.n284 VTAIL.n283 3.49141
R413 VTAIL.n26 VTAIL.n25 3.49141
R414 VTAIL.n62 VTAIL.n61 3.49141
R415 VTAIL.n100 VTAIL.n99 3.49141
R416 VTAIL.n248 VTAIL.n247 3.49141
R417 VTAIL.n210 VTAIL.n209 3.49141
R418 VTAIL.n174 VTAIL.n173 3.49141
R419 VTAIL.n136 VTAIL.n135 3.49141
R420 VTAIL.n0 VTAIL.t10 2.93383
R421 VTAIL.n0 VTAIL.t15 2.93383
R422 VTAIL.n74 VTAIL.t2 2.93383
R423 VTAIL.n74 VTAIL.t6 2.93383
R424 VTAIL.n222 VTAIL.t3 2.93383
R425 VTAIL.n222 VTAIL.t0 2.93383
R426 VTAIL.n148 VTAIL.t9 2.93383
R427 VTAIL.n148 VTAIL.t13 2.93383
R428 VTAIL.n280 VTAIL.n266 2.71565
R429 VTAIL.n22 VTAIL.n8 2.71565
R430 VTAIL.n58 VTAIL.n44 2.71565
R431 VTAIL.n96 VTAIL.n82 2.71565
R432 VTAIL.n244 VTAIL.n230 2.71565
R433 VTAIL.n206 VTAIL.n192 2.71565
R434 VTAIL.n170 VTAIL.n156 2.71565
R435 VTAIL.n132 VTAIL.n118 2.71565
R436 VTAIL.n279 VTAIL.n268 1.93989
R437 VTAIL.n21 VTAIL.n10 1.93989
R438 VTAIL.n57 VTAIL.n46 1.93989
R439 VTAIL.n95 VTAIL.n84 1.93989
R440 VTAIL.n243 VTAIL.n232 1.93989
R441 VTAIL.n205 VTAIL.n194 1.93989
R442 VTAIL.n169 VTAIL.n158 1.93989
R443 VTAIL.n131 VTAIL.n120 1.93989
R444 VTAIL.n149 VTAIL.n147 1.30222
R445 VTAIL.n185 VTAIL.n149 1.30222
R446 VTAIL.n223 VTAIL.n221 1.30222
R447 VTAIL.n259 VTAIL.n223 1.30222
R448 VTAIL.n111 VTAIL.n75 1.30222
R449 VTAIL.n75 VTAIL.n73 1.30222
R450 VTAIL.n37 VTAIL.n1 1.30222
R451 VTAIL VTAIL.n295 1.24403
R452 VTAIL.n276 VTAIL.n275 1.16414
R453 VTAIL.n18 VTAIL.n17 1.16414
R454 VTAIL.n54 VTAIL.n53 1.16414
R455 VTAIL.n92 VTAIL.n91 1.16414
R456 VTAIL.n240 VTAIL.n239 1.16414
R457 VTAIL.n202 VTAIL.n201 1.16414
R458 VTAIL.n166 VTAIL.n165 1.16414
R459 VTAIL.n128 VTAIL.n127 1.16414
R460 VTAIL.n221 VTAIL.n185 0.470328
R461 VTAIL.n73 VTAIL.n37 0.470328
R462 VTAIL.n272 VTAIL.n270 0.388379
R463 VTAIL.n14 VTAIL.n12 0.388379
R464 VTAIL.n50 VTAIL.n48 0.388379
R465 VTAIL.n88 VTAIL.n86 0.388379
R466 VTAIL.n236 VTAIL.n234 0.388379
R467 VTAIL.n198 VTAIL.n196 0.388379
R468 VTAIL.n162 VTAIL.n160 0.388379
R469 VTAIL.n124 VTAIL.n122 0.388379
R470 VTAIL.n277 VTAIL.n269 0.155672
R471 VTAIL.n278 VTAIL.n277 0.155672
R472 VTAIL.n278 VTAIL.n265 0.155672
R473 VTAIL.n285 VTAIL.n265 0.155672
R474 VTAIL.n286 VTAIL.n285 0.155672
R475 VTAIL.n286 VTAIL.n261 0.155672
R476 VTAIL.n293 VTAIL.n261 0.155672
R477 VTAIL.n19 VTAIL.n11 0.155672
R478 VTAIL.n20 VTAIL.n19 0.155672
R479 VTAIL.n20 VTAIL.n7 0.155672
R480 VTAIL.n27 VTAIL.n7 0.155672
R481 VTAIL.n28 VTAIL.n27 0.155672
R482 VTAIL.n28 VTAIL.n3 0.155672
R483 VTAIL.n35 VTAIL.n3 0.155672
R484 VTAIL.n55 VTAIL.n47 0.155672
R485 VTAIL.n56 VTAIL.n55 0.155672
R486 VTAIL.n56 VTAIL.n43 0.155672
R487 VTAIL.n63 VTAIL.n43 0.155672
R488 VTAIL.n64 VTAIL.n63 0.155672
R489 VTAIL.n64 VTAIL.n39 0.155672
R490 VTAIL.n71 VTAIL.n39 0.155672
R491 VTAIL.n93 VTAIL.n85 0.155672
R492 VTAIL.n94 VTAIL.n93 0.155672
R493 VTAIL.n94 VTAIL.n81 0.155672
R494 VTAIL.n101 VTAIL.n81 0.155672
R495 VTAIL.n102 VTAIL.n101 0.155672
R496 VTAIL.n102 VTAIL.n77 0.155672
R497 VTAIL.n109 VTAIL.n77 0.155672
R498 VTAIL.n257 VTAIL.n225 0.155672
R499 VTAIL.n250 VTAIL.n225 0.155672
R500 VTAIL.n250 VTAIL.n249 0.155672
R501 VTAIL.n249 VTAIL.n229 0.155672
R502 VTAIL.n242 VTAIL.n229 0.155672
R503 VTAIL.n242 VTAIL.n241 0.155672
R504 VTAIL.n241 VTAIL.n233 0.155672
R505 VTAIL.n219 VTAIL.n187 0.155672
R506 VTAIL.n212 VTAIL.n187 0.155672
R507 VTAIL.n212 VTAIL.n211 0.155672
R508 VTAIL.n211 VTAIL.n191 0.155672
R509 VTAIL.n204 VTAIL.n191 0.155672
R510 VTAIL.n204 VTAIL.n203 0.155672
R511 VTAIL.n203 VTAIL.n195 0.155672
R512 VTAIL.n183 VTAIL.n151 0.155672
R513 VTAIL.n176 VTAIL.n151 0.155672
R514 VTAIL.n176 VTAIL.n175 0.155672
R515 VTAIL.n175 VTAIL.n155 0.155672
R516 VTAIL.n168 VTAIL.n155 0.155672
R517 VTAIL.n168 VTAIL.n167 0.155672
R518 VTAIL.n167 VTAIL.n159 0.155672
R519 VTAIL.n145 VTAIL.n113 0.155672
R520 VTAIL.n138 VTAIL.n113 0.155672
R521 VTAIL.n138 VTAIL.n137 0.155672
R522 VTAIL.n137 VTAIL.n117 0.155672
R523 VTAIL.n130 VTAIL.n117 0.155672
R524 VTAIL.n130 VTAIL.n129 0.155672
R525 VTAIL.n129 VTAIL.n121 0.155672
R526 VTAIL VTAIL.n1 0.0586897
R527 B.n446 B.n445 585
R528 B.n447 B.n94 585
R529 B.n449 B.n448 585
R530 B.n451 B.n93 585
R531 B.n454 B.n453 585
R532 B.n455 B.n92 585
R533 B.n457 B.n456 585
R534 B.n459 B.n91 585
R535 B.n462 B.n461 585
R536 B.n463 B.n90 585
R537 B.n465 B.n464 585
R538 B.n467 B.n89 585
R539 B.n470 B.n469 585
R540 B.n471 B.n88 585
R541 B.n473 B.n472 585
R542 B.n475 B.n87 585
R543 B.n478 B.n477 585
R544 B.n479 B.n86 585
R545 B.n481 B.n480 585
R546 B.n483 B.n85 585
R547 B.n486 B.n485 585
R548 B.n487 B.n84 585
R549 B.n489 B.n488 585
R550 B.n491 B.n83 585
R551 B.n493 B.n492 585
R552 B.n495 B.n494 585
R553 B.n498 B.n497 585
R554 B.n499 B.n78 585
R555 B.n501 B.n500 585
R556 B.n503 B.n77 585
R557 B.n506 B.n505 585
R558 B.n507 B.n76 585
R559 B.n509 B.n508 585
R560 B.n511 B.n75 585
R561 B.n513 B.n512 585
R562 B.n515 B.n514 585
R563 B.n518 B.n517 585
R564 B.n519 B.n70 585
R565 B.n521 B.n520 585
R566 B.n523 B.n69 585
R567 B.n526 B.n525 585
R568 B.n527 B.n68 585
R569 B.n529 B.n528 585
R570 B.n531 B.n67 585
R571 B.n534 B.n533 585
R572 B.n535 B.n66 585
R573 B.n537 B.n536 585
R574 B.n539 B.n65 585
R575 B.n542 B.n541 585
R576 B.n543 B.n64 585
R577 B.n545 B.n544 585
R578 B.n547 B.n63 585
R579 B.n550 B.n549 585
R580 B.n551 B.n62 585
R581 B.n553 B.n552 585
R582 B.n555 B.n61 585
R583 B.n558 B.n557 585
R584 B.n559 B.n60 585
R585 B.n561 B.n560 585
R586 B.n563 B.n59 585
R587 B.n566 B.n565 585
R588 B.n567 B.n58 585
R589 B.n443 B.n56 585
R590 B.n570 B.n56 585
R591 B.n442 B.n55 585
R592 B.n571 B.n55 585
R593 B.n441 B.n54 585
R594 B.n572 B.n54 585
R595 B.n440 B.n439 585
R596 B.n439 B.n50 585
R597 B.n438 B.n49 585
R598 B.n578 B.n49 585
R599 B.n437 B.n48 585
R600 B.n579 B.n48 585
R601 B.n436 B.n47 585
R602 B.n580 B.n47 585
R603 B.n435 B.n434 585
R604 B.n434 B.n43 585
R605 B.n433 B.n42 585
R606 B.n586 B.n42 585
R607 B.n432 B.n41 585
R608 B.n587 B.n41 585
R609 B.n431 B.n40 585
R610 B.n588 B.n40 585
R611 B.n430 B.n429 585
R612 B.n429 B.n36 585
R613 B.n428 B.n35 585
R614 B.n594 B.n35 585
R615 B.n427 B.n34 585
R616 B.n595 B.n34 585
R617 B.n426 B.n33 585
R618 B.n596 B.n33 585
R619 B.n425 B.n424 585
R620 B.n424 B.n29 585
R621 B.n423 B.n28 585
R622 B.n602 B.n28 585
R623 B.n422 B.n27 585
R624 B.n603 B.n27 585
R625 B.n421 B.n26 585
R626 B.n604 B.n26 585
R627 B.n420 B.n419 585
R628 B.n419 B.n22 585
R629 B.n418 B.n21 585
R630 B.n610 B.n21 585
R631 B.n417 B.n20 585
R632 B.n611 B.n20 585
R633 B.n416 B.n19 585
R634 B.n612 B.n19 585
R635 B.n415 B.n414 585
R636 B.n414 B.n15 585
R637 B.n413 B.n14 585
R638 B.n618 B.n14 585
R639 B.n412 B.n13 585
R640 B.n619 B.n13 585
R641 B.n411 B.n12 585
R642 B.n620 B.n12 585
R643 B.n410 B.n409 585
R644 B.n409 B.n408 585
R645 B.n407 B.n406 585
R646 B.n407 B.n8 585
R647 B.n405 B.n7 585
R648 B.n627 B.n7 585
R649 B.n404 B.n6 585
R650 B.n628 B.n6 585
R651 B.n403 B.n5 585
R652 B.n629 B.n5 585
R653 B.n402 B.n401 585
R654 B.n401 B.n4 585
R655 B.n400 B.n95 585
R656 B.n400 B.n399 585
R657 B.n390 B.n96 585
R658 B.n97 B.n96 585
R659 B.n392 B.n391 585
R660 B.n393 B.n392 585
R661 B.n389 B.n102 585
R662 B.n102 B.n101 585
R663 B.n388 B.n387 585
R664 B.n387 B.n386 585
R665 B.n104 B.n103 585
R666 B.n105 B.n104 585
R667 B.n379 B.n378 585
R668 B.n380 B.n379 585
R669 B.n377 B.n110 585
R670 B.n110 B.n109 585
R671 B.n376 B.n375 585
R672 B.n375 B.n374 585
R673 B.n112 B.n111 585
R674 B.n113 B.n112 585
R675 B.n367 B.n366 585
R676 B.n368 B.n367 585
R677 B.n365 B.n117 585
R678 B.n121 B.n117 585
R679 B.n364 B.n363 585
R680 B.n363 B.n362 585
R681 B.n119 B.n118 585
R682 B.n120 B.n119 585
R683 B.n355 B.n354 585
R684 B.n356 B.n355 585
R685 B.n353 B.n125 585
R686 B.n129 B.n125 585
R687 B.n352 B.n351 585
R688 B.n351 B.n350 585
R689 B.n127 B.n126 585
R690 B.n128 B.n127 585
R691 B.n343 B.n342 585
R692 B.n344 B.n343 585
R693 B.n341 B.n134 585
R694 B.n134 B.n133 585
R695 B.n340 B.n339 585
R696 B.n339 B.n338 585
R697 B.n136 B.n135 585
R698 B.n137 B.n136 585
R699 B.n331 B.n330 585
R700 B.n332 B.n331 585
R701 B.n329 B.n141 585
R702 B.n145 B.n141 585
R703 B.n328 B.n327 585
R704 B.n327 B.n326 585
R705 B.n143 B.n142 585
R706 B.n144 B.n143 585
R707 B.n319 B.n318 585
R708 B.n320 B.n319 585
R709 B.n317 B.n150 585
R710 B.n150 B.n149 585
R711 B.n316 B.n315 585
R712 B.n315 B.n314 585
R713 B.n311 B.n154 585
R714 B.n310 B.n309 585
R715 B.n307 B.n155 585
R716 B.n307 B.n153 585
R717 B.n306 B.n305 585
R718 B.n304 B.n303 585
R719 B.n302 B.n157 585
R720 B.n300 B.n299 585
R721 B.n298 B.n158 585
R722 B.n297 B.n296 585
R723 B.n294 B.n159 585
R724 B.n292 B.n291 585
R725 B.n290 B.n160 585
R726 B.n289 B.n288 585
R727 B.n286 B.n161 585
R728 B.n284 B.n283 585
R729 B.n282 B.n162 585
R730 B.n281 B.n280 585
R731 B.n278 B.n163 585
R732 B.n276 B.n275 585
R733 B.n274 B.n164 585
R734 B.n273 B.n272 585
R735 B.n270 B.n165 585
R736 B.n268 B.n267 585
R737 B.n266 B.n166 585
R738 B.n265 B.n264 585
R739 B.n262 B.n167 585
R740 B.n260 B.n259 585
R741 B.n258 B.n168 585
R742 B.n257 B.n256 585
R743 B.n254 B.n172 585
R744 B.n252 B.n251 585
R745 B.n250 B.n173 585
R746 B.n249 B.n248 585
R747 B.n246 B.n174 585
R748 B.n244 B.n243 585
R749 B.n242 B.n175 585
R750 B.n240 B.n239 585
R751 B.n237 B.n178 585
R752 B.n235 B.n234 585
R753 B.n233 B.n179 585
R754 B.n232 B.n231 585
R755 B.n229 B.n180 585
R756 B.n227 B.n226 585
R757 B.n225 B.n181 585
R758 B.n224 B.n223 585
R759 B.n221 B.n182 585
R760 B.n219 B.n218 585
R761 B.n217 B.n183 585
R762 B.n216 B.n215 585
R763 B.n213 B.n184 585
R764 B.n211 B.n210 585
R765 B.n209 B.n185 585
R766 B.n208 B.n207 585
R767 B.n205 B.n186 585
R768 B.n203 B.n202 585
R769 B.n201 B.n187 585
R770 B.n200 B.n199 585
R771 B.n197 B.n188 585
R772 B.n195 B.n194 585
R773 B.n193 B.n189 585
R774 B.n192 B.n191 585
R775 B.n152 B.n151 585
R776 B.n153 B.n152 585
R777 B.n313 B.n312 585
R778 B.n314 B.n313 585
R779 B.n148 B.n147 585
R780 B.n149 B.n148 585
R781 B.n322 B.n321 585
R782 B.n321 B.n320 585
R783 B.n323 B.n146 585
R784 B.n146 B.n144 585
R785 B.n325 B.n324 585
R786 B.n326 B.n325 585
R787 B.n140 B.n139 585
R788 B.n145 B.n140 585
R789 B.n334 B.n333 585
R790 B.n333 B.n332 585
R791 B.n335 B.n138 585
R792 B.n138 B.n137 585
R793 B.n337 B.n336 585
R794 B.n338 B.n337 585
R795 B.n132 B.n131 585
R796 B.n133 B.n132 585
R797 B.n346 B.n345 585
R798 B.n345 B.n344 585
R799 B.n347 B.n130 585
R800 B.n130 B.n128 585
R801 B.n349 B.n348 585
R802 B.n350 B.n349 585
R803 B.n124 B.n123 585
R804 B.n129 B.n124 585
R805 B.n358 B.n357 585
R806 B.n357 B.n356 585
R807 B.n359 B.n122 585
R808 B.n122 B.n120 585
R809 B.n361 B.n360 585
R810 B.n362 B.n361 585
R811 B.n116 B.n115 585
R812 B.n121 B.n116 585
R813 B.n370 B.n369 585
R814 B.n369 B.n368 585
R815 B.n371 B.n114 585
R816 B.n114 B.n113 585
R817 B.n373 B.n372 585
R818 B.n374 B.n373 585
R819 B.n108 B.n107 585
R820 B.n109 B.n108 585
R821 B.n382 B.n381 585
R822 B.n381 B.n380 585
R823 B.n383 B.n106 585
R824 B.n106 B.n105 585
R825 B.n385 B.n384 585
R826 B.n386 B.n385 585
R827 B.n100 B.n99 585
R828 B.n101 B.n100 585
R829 B.n395 B.n394 585
R830 B.n394 B.n393 585
R831 B.n396 B.n98 585
R832 B.n98 B.n97 585
R833 B.n398 B.n397 585
R834 B.n399 B.n398 585
R835 B.n3 B.n0 585
R836 B.n4 B.n3 585
R837 B.n626 B.n1 585
R838 B.n627 B.n626 585
R839 B.n625 B.n624 585
R840 B.n625 B.n8 585
R841 B.n623 B.n9 585
R842 B.n408 B.n9 585
R843 B.n622 B.n621 585
R844 B.n621 B.n620 585
R845 B.n11 B.n10 585
R846 B.n619 B.n11 585
R847 B.n617 B.n616 585
R848 B.n618 B.n617 585
R849 B.n615 B.n16 585
R850 B.n16 B.n15 585
R851 B.n614 B.n613 585
R852 B.n613 B.n612 585
R853 B.n18 B.n17 585
R854 B.n611 B.n18 585
R855 B.n609 B.n608 585
R856 B.n610 B.n609 585
R857 B.n607 B.n23 585
R858 B.n23 B.n22 585
R859 B.n606 B.n605 585
R860 B.n605 B.n604 585
R861 B.n25 B.n24 585
R862 B.n603 B.n25 585
R863 B.n601 B.n600 585
R864 B.n602 B.n601 585
R865 B.n599 B.n30 585
R866 B.n30 B.n29 585
R867 B.n598 B.n597 585
R868 B.n597 B.n596 585
R869 B.n32 B.n31 585
R870 B.n595 B.n32 585
R871 B.n593 B.n592 585
R872 B.n594 B.n593 585
R873 B.n591 B.n37 585
R874 B.n37 B.n36 585
R875 B.n590 B.n589 585
R876 B.n589 B.n588 585
R877 B.n39 B.n38 585
R878 B.n587 B.n39 585
R879 B.n585 B.n584 585
R880 B.n586 B.n585 585
R881 B.n583 B.n44 585
R882 B.n44 B.n43 585
R883 B.n582 B.n581 585
R884 B.n581 B.n580 585
R885 B.n46 B.n45 585
R886 B.n579 B.n46 585
R887 B.n577 B.n576 585
R888 B.n578 B.n577 585
R889 B.n575 B.n51 585
R890 B.n51 B.n50 585
R891 B.n574 B.n573 585
R892 B.n573 B.n572 585
R893 B.n53 B.n52 585
R894 B.n571 B.n53 585
R895 B.n569 B.n568 585
R896 B.n570 B.n569 585
R897 B.n630 B.n629 585
R898 B.n628 B.n2 585
R899 B.n569 B.n58 463.671
R900 B.n445 B.n56 463.671
R901 B.n315 B.n152 463.671
R902 B.n313 B.n154 463.671
R903 B.n71 B.t8 341.872
R904 B.n79 B.t16 341.872
R905 B.n176 B.t12 341.872
R906 B.n169 B.t19 341.872
R907 B.n444 B.n57 256.663
R908 B.n450 B.n57 256.663
R909 B.n452 B.n57 256.663
R910 B.n458 B.n57 256.663
R911 B.n460 B.n57 256.663
R912 B.n466 B.n57 256.663
R913 B.n468 B.n57 256.663
R914 B.n474 B.n57 256.663
R915 B.n476 B.n57 256.663
R916 B.n482 B.n57 256.663
R917 B.n484 B.n57 256.663
R918 B.n490 B.n57 256.663
R919 B.n82 B.n57 256.663
R920 B.n496 B.n57 256.663
R921 B.n502 B.n57 256.663
R922 B.n504 B.n57 256.663
R923 B.n510 B.n57 256.663
R924 B.n74 B.n57 256.663
R925 B.n516 B.n57 256.663
R926 B.n522 B.n57 256.663
R927 B.n524 B.n57 256.663
R928 B.n530 B.n57 256.663
R929 B.n532 B.n57 256.663
R930 B.n538 B.n57 256.663
R931 B.n540 B.n57 256.663
R932 B.n546 B.n57 256.663
R933 B.n548 B.n57 256.663
R934 B.n554 B.n57 256.663
R935 B.n556 B.n57 256.663
R936 B.n562 B.n57 256.663
R937 B.n564 B.n57 256.663
R938 B.n308 B.n153 256.663
R939 B.n156 B.n153 256.663
R940 B.n301 B.n153 256.663
R941 B.n295 B.n153 256.663
R942 B.n293 B.n153 256.663
R943 B.n287 B.n153 256.663
R944 B.n285 B.n153 256.663
R945 B.n279 B.n153 256.663
R946 B.n277 B.n153 256.663
R947 B.n271 B.n153 256.663
R948 B.n269 B.n153 256.663
R949 B.n263 B.n153 256.663
R950 B.n261 B.n153 256.663
R951 B.n255 B.n153 256.663
R952 B.n253 B.n153 256.663
R953 B.n247 B.n153 256.663
R954 B.n245 B.n153 256.663
R955 B.n238 B.n153 256.663
R956 B.n236 B.n153 256.663
R957 B.n230 B.n153 256.663
R958 B.n228 B.n153 256.663
R959 B.n222 B.n153 256.663
R960 B.n220 B.n153 256.663
R961 B.n214 B.n153 256.663
R962 B.n212 B.n153 256.663
R963 B.n206 B.n153 256.663
R964 B.n204 B.n153 256.663
R965 B.n198 B.n153 256.663
R966 B.n196 B.n153 256.663
R967 B.n190 B.n153 256.663
R968 B.n632 B.n631 256.663
R969 B.n79 B.t17 221.308
R970 B.n176 B.t15 221.308
R971 B.n71 B.t10 221.308
R972 B.n169 B.t21 221.308
R973 B.n80 B.t18 192.023
R974 B.n177 B.t14 192.023
R975 B.n72 B.t11 192.023
R976 B.n170 B.t20 192.023
R977 B.n565 B.n563 163.367
R978 B.n561 B.n60 163.367
R979 B.n557 B.n555 163.367
R980 B.n553 B.n62 163.367
R981 B.n549 B.n547 163.367
R982 B.n545 B.n64 163.367
R983 B.n541 B.n539 163.367
R984 B.n537 B.n66 163.367
R985 B.n533 B.n531 163.367
R986 B.n529 B.n68 163.367
R987 B.n525 B.n523 163.367
R988 B.n521 B.n70 163.367
R989 B.n517 B.n515 163.367
R990 B.n512 B.n511 163.367
R991 B.n509 B.n76 163.367
R992 B.n505 B.n503 163.367
R993 B.n501 B.n78 163.367
R994 B.n497 B.n495 163.367
R995 B.n492 B.n491 163.367
R996 B.n489 B.n84 163.367
R997 B.n485 B.n483 163.367
R998 B.n481 B.n86 163.367
R999 B.n477 B.n475 163.367
R1000 B.n473 B.n88 163.367
R1001 B.n469 B.n467 163.367
R1002 B.n465 B.n90 163.367
R1003 B.n461 B.n459 163.367
R1004 B.n457 B.n92 163.367
R1005 B.n453 B.n451 163.367
R1006 B.n449 B.n94 163.367
R1007 B.n315 B.n150 163.367
R1008 B.n319 B.n150 163.367
R1009 B.n319 B.n143 163.367
R1010 B.n327 B.n143 163.367
R1011 B.n327 B.n141 163.367
R1012 B.n331 B.n141 163.367
R1013 B.n331 B.n136 163.367
R1014 B.n339 B.n136 163.367
R1015 B.n339 B.n134 163.367
R1016 B.n343 B.n134 163.367
R1017 B.n343 B.n127 163.367
R1018 B.n351 B.n127 163.367
R1019 B.n351 B.n125 163.367
R1020 B.n355 B.n125 163.367
R1021 B.n355 B.n119 163.367
R1022 B.n363 B.n119 163.367
R1023 B.n363 B.n117 163.367
R1024 B.n367 B.n117 163.367
R1025 B.n367 B.n112 163.367
R1026 B.n375 B.n112 163.367
R1027 B.n375 B.n110 163.367
R1028 B.n379 B.n110 163.367
R1029 B.n379 B.n104 163.367
R1030 B.n387 B.n104 163.367
R1031 B.n387 B.n102 163.367
R1032 B.n392 B.n102 163.367
R1033 B.n392 B.n96 163.367
R1034 B.n400 B.n96 163.367
R1035 B.n401 B.n400 163.367
R1036 B.n401 B.n5 163.367
R1037 B.n6 B.n5 163.367
R1038 B.n7 B.n6 163.367
R1039 B.n407 B.n7 163.367
R1040 B.n409 B.n407 163.367
R1041 B.n409 B.n12 163.367
R1042 B.n13 B.n12 163.367
R1043 B.n14 B.n13 163.367
R1044 B.n414 B.n14 163.367
R1045 B.n414 B.n19 163.367
R1046 B.n20 B.n19 163.367
R1047 B.n21 B.n20 163.367
R1048 B.n419 B.n21 163.367
R1049 B.n419 B.n26 163.367
R1050 B.n27 B.n26 163.367
R1051 B.n28 B.n27 163.367
R1052 B.n424 B.n28 163.367
R1053 B.n424 B.n33 163.367
R1054 B.n34 B.n33 163.367
R1055 B.n35 B.n34 163.367
R1056 B.n429 B.n35 163.367
R1057 B.n429 B.n40 163.367
R1058 B.n41 B.n40 163.367
R1059 B.n42 B.n41 163.367
R1060 B.n434 B.n42 163.367
R1061 B.n434 B.n47 163.367
R1062 B.n48 B.n47 163.367
R1063 B.n49 B.n48 163.367
R1064 B.n439 B.n49 163.367
R1065 B.n439 B.n54 163.367
R1066 B.n55 B.n54 163.367
R1067 B.n56 B.n55 163.367
R1068 B.n309 B.n307 163.367
R1069 B.n307 B.n306 163.367
R1070 B.n303 B.n302 163.367
R1071 B.n300 B.n158 163.367
R1072 B.n296 B.n294 163.367
R1073 B.n292 B.n160 163.367
R1074 B.n288 B.n286 163.367
R1075 B.n284 B.n162 163.367
R1076 B.n280 B.n278 163.367
R1077 B.n276 B.n164 163.367
R1078 B.n272 B.n270 163.367
R1079 B.n268 B.n166 163.367
R1080 B.n264 B.n262 163.367
R1081 B.n260 B.n168 163.367
R1082 B.n256 B.n254 163.367
R1083 B.n252 B.n173 163.367
R1084 B.n248 B.n246 163.367
R1085 B.n244 B.n175 163.367
R1086 B.n239 B.n237 163.367
R1087 B.n235 B.n179 163.367
R1088 B.n231 B.n229 163.367
R1089 B.n227 B.n181 163.367
R1090 B.n223 B.n221 163.367
R1091 B.n219 B.n183 163.367
R1092 B.n215 B.n213 163.367
R1093 B.n211 B.n185 163.367
R1094 B.n207 B.n205 163.367
R1095 B.n203 B.n187 163.367
R1096 B.n199 B.n197 163.367
R1097 B.n195 B.n189 163.367
R1098 B.n191 B.n152 163.367
R1099 B.n313 B.n148 163.367
R1100 B.n321 B.n148 163.367
R1101 B.n321 B.n146 163.367
R1102 B.n325 B.n146 163.367
R1103 B.n325 B.n140 163.367
R1104 B.n333 B.n140 163.367
R1105 B.n333 B.n138 163.367
R1106 B.n337 B.n138 163.367
R1107 B.n337 B.n132 163.367
R1108 B.n345 B.n132 163.367
R1109 B.n345 B.n130 163.367
R1110 B.n349 B.n130 163.367
R1111 B.n349 B.n124 163.367
R1112 B.n357 B.n124 163.367
R1113 B.n357 B.n122 163.367
R1114 B.n361 B.n122 163.367
R1115 B.n361 B.n116 163.367
R1116 B.n369 B.n116 163.367
R1117 B.n369 B.n114 163.367
R1118 B.n373 B.n114 163.367
R1119 B.n373 B.n108 163.367
R1120 B.n381 B.n108 163.367
R1121 B.n381 B.n106 163.367
R1122 B.n385 B.n106 163.367
R1123 B.n385 B.n100 163.367
R1124 B.n394 B.n100 163.367
R1125 B.n394 B.n98 163.367
R1126 B.n398 B.n98 163.367
R1127 B.n398 B.n3 163.367
R1128 B.n630 B.n3 163.367
R1129 B.n626 B.n2 163.367
R1130 B.n626 B.n625 163.367
R1131 B.n625 B.n9 163.367
R1132 B.n621 B.n9 163.367
R1133 B.n621 B.n11 163.367
R1134 B.n617 B.n11 163.367
R1135 B.n617 B.n16 163.367
R1136 B.n613 B.n16 163.367
R1137 B.n613 B.n18 163.367
R1138 B.n609 B.n18 163.367
R1139 B.n609 B.n23 163.367
R1140 B.n605 B.n23 163.367
R1141 B.n605 B.n25 163.367
R1142 B.n601 B.n25 163.367
R1143 B.n601 B.n30 163.367
R1144 B.n597 B.n30 163.367
R1145 B.n597 B.n32 163.367
R1146 B.n593 B.n32 163.367
R1147 B.n593 B.n37 163.367
R1148 B.n589 B.n37 163.367
R1149 B.n589 B.n39 163.367
R1150 B.n585 B.n39 163.367
R1151 B.n585 B.n44 163.367
R1152 B.n581 B.n44 163.367
R1153 B.n581 B.n46 163.367
R1154 B.n577 B.n46 163.367
R1155 B.n577 B.n51 163.367
R1156 B.n573 B.n51 163.367
R1157 B.n573 B.n53 163.367
R1158 B.n569 B.n53 163.367
R1159 B.n314 B.n153 101.538
R1160 B.n570 B.n57 101.538
R1161 B.n564 B.n58 71.676
R1162 B.n563 B.n562 71.676
R1163 B.n556 B.n60 71.676
R1164 B.n555 B.n554 71.676
R1165 B.n548 B.n62 71.676
R1166 B.n547 B.n546 71.676
R1167 B.n540 B.n64 71.676
R1168 B.n539 B.n538 71.676
R1169 B.n532 B.n66 71.676
R1170 B.n531 B.n530 71.676
R1171 B.n524 B.n68 71.676
R1172 B.n523 B.n522 71.676
R1173 B.n516 B.n70 71.676
R1174 B.n515 B.n74 71.676
R1175 B.n511 B.n510 71.676
R1176 B.n504 B.n76 71.676
R1177 B.n503 B.n502 71.676
R1178 B.n496 B.n78 71.676
R1179 B.n495 B.n82 71.676
R1180 B.n491 B.n490 71.676
R1181 B.n484 B.n84 71.676
R1182 B.n483 B.n482 71.676
R1183 B.n476 B.n86 71.676
R1184 B.n475 B.n474 71.676
R1185 B.n468 B.n88 71.676
R1186 B.n467 B.n466 71.676
R1187 B.n460 B.n90 71.676
R1188 B.n459 B.n458 71.676
R1189 B.n452 B.n92 71.676
R1190 B.n451 B.n450 71.676
R1191 B.n444 B.n94 71.676
R1192 B.n445 B.n444 71.676
R1193 B.n450 B.n449 71.676
R1194 B.n453 B.n452 71.676
R1195 B.n458 B.n457 71.676
R1196 B.n461 B.n460 71.676
R1197 B.n466 B.n465 71.676
R1198 B.n469 B.n468 71.676
R1199 B.n474 B.n473 71.676
R1200 B.n477 B.n476 71.676
R1201 B.n482 B.n481 71.676
R1202 B.n485 B.n484 71.676
R1203 B.n490 B.n489 71.676
R1204 B.n492 B.n82 71.676
R1205 B.n497 B.n496 71.676
R1206 B.n502 B.n501 71.676
R1207 B.n505 B.n504 71.676
R1208 B.n510 B.n509 71.676
R1209 B.n512 B.n74 71.676
R1210 B.n517 B.n516 71.676
R1211 B.n522 B.n521 71.676
R1212 B.n525 B.n524 71.676
R1213 B.n530 B.n529 71.676
R1214 B.n533 B.n532 71.676
R1215 B.n538 B.n537 71.676
R1216 B.n541 B.n540 71.676
R1217 B.n546 B.n545 71.676
R1218 B.n549 B.n548 71.676
R1219 B.n554 B.n553 71.676
R1220 B.n557 B.n556 71.676
R1221 B.n562 B.n561 71.676
R1222 B.n565 B.n564 71.676
R1223 B.n308 B.n154 71.676
R1224 B.n306 B.n156 71.676
R1225 B.n302 B.n301 71.676
R1226 B.n295 B.n158 71.676
R1227 B.n294 B.n293 71.676
R1228 B.n287 B.n160 71.676
R1229 B.n286 B.n285 71.676
R1230 B.n279 B.n162 71.676
R1231 B.n278 B.n277 71.676
R1232 B.n271 B.n164 71.676
R1233 B.n270 B.n269 71.676
R1234 B.n263 B.n166 71.676
R1235 B.n262 B.n261 71.676
R1236 B.n255 B.n168 71.676
R1237 B.n254 B.n253 71.676
R1238 B.n247 B.n173 71.676
R1239 B.n246 B.n245 71.676
R1240 B.n238 B.n175 71.676
R1241 B.n237 B.n236 71.676
R1242 B.n230 B.n179 71.676
R1243 B.n229 B.n228 71.676
R1244 B.n222 B.n181 71.676
R1245 B.n221 B.n220 71.676
R1246 B.n214 B.n183 71.676
R1247 B.n213 B.n212 71.676
R1248 B.n206 B.n185 71.676
R1249 B.n205 B.n204 71.676
R1250 B.n198 B.n187 71.676
R1251 B.n197 B.n196 71.676
R1252 B.n190 B.n189 71.676
R1253 B.n309 B.n308 71.676
R1254 B.n303 B.n156 71.676
R1255 B.n301 B.n300 71.676
R1256 B.n296 B.n295 71.676
R1257 B.n293 B.n292 71.676
R1258 B.n288 B.n287 71.676
R1259 B.n285 B.n284 71.676
R1260 B.n280 B.n279 71.676
R1261 B.n277 B.n276 71.676
R1262 B.n272 B.n271 71.676
R1263 B.n269 B.n268 71.676
R1264 B.n264 B.n263 71.676
R1265 B.n261 B.n260 71.676
R1266 B.n256 B.n255 71.676
R1267 B.n253 B.n252 71.676
R1268 B.n248 B.n247 71.676
R1269 B.n245 B.n244 71.676
R1270 B.n239 B.n238 71.676
R1271 B.n236 B.n235 71.676
R1272 B.n231 B.n230 71.676
R1273 B.n228 B.n227 71.676
R1274 B.n223 B.n222 71.676
R1275 B.n220 B.n219 71.676
R1276 B.n215 B.n214 71.676
R1277 B.n212 B.n211 71.676
R1278 B.n207 B.n206 71.676
R1279 B.n204 B.n203 71.676
R1280 B.n199 B.n198 71.676
R1281 B.n196 B.n195 71.676
R1282 B.n191 B.n190 71.676
R1283 B.n631 B.n630 71.676
R1284 B.n631 B.n2 71.676
R1285 B.n314 B.n149 62.2042
R1286 B.n320 B.n149 62.2042
R1287 B.n320 B.n144 62.2042
R1288 B.n326 B.n144 62.2042
R1289 B.n326 B.n145 62.2042
R1290 B.n332 B.n137 62.2042
R1291 B.n338 B.n137 62.2042
R1292 B.n338 B.n133 62.2042
R1293 B.n344 B.n133 62.2042
R1294 B.n344 B.n128 62.2042
R1295 B.n350 B.n128 62.2042
R1296 B.n350 B.n129 62.2042
R1297 B.n356 B.n120 62.2042
R1298 B.n362 B.n120 62.2042
R1299 B.n362 B.n121 62.2042
R1300 B.n368 B.n113 62.2042
R1301 B.n374 B.n113 62.2042
R1302 B.n374 B.n109 62.2042
R1303 B.n380 B.n109 62.2042
R1304 B.n386 B.n105 62.2042
R1305 B.n386 B.n101 62.2042
R1306 B.n393 B.n101 62.2042
R1307 B.n399 B.n97 62.2042
R1308 B.n399 B.n4 62.2042
R1309 B.n629 B.n4 62.2042
R1310 B.n629 B.n628 62.2042
R1311 B.n628 B.n627 62.2042
R1312 B.n627 B.n8 62.2042
R1313 B.n408 B.n8 62.2042
R1314 B.n620 B.n619 62.2042
R1315 B.n619 B.n618 62.2042
R1316 B.n618 B.n15 62.2042
R1317 B.n612 B.n611 62.2042
R1318 B.n611 B.n610 62.2042
R1319 B.n610 B.n22 62.2042
R1320 B.n604 B.n22 62.2042
R1321 B.n603 B.n602 62.2042
R1322 B.n602 B.n29 62.2042
R1323 B.n596 B.n29 62.2042
R1324 B.n595 B.n594 62.2042
R1325 B.n594 B.n36 62.2042
R1326 B.n588 B.n36 62.2042
R1327 B.n588 B.n587 62.2042
R1328 B.n587 B.n586 62.2042
R1329 B.n586 B.n43 62.2042
R1330 B.n580 B.n43 62.2042
R1331 B.n579 B.n578 62.2042
R1332 B.n578 B.n50 62.2042
R1333 B.n572 B.n50 62.2042
R1334 B.n572 B.n571 62.2042
R1335 B.n571 B.n570 62.2042
R1336 B.n73 B.n72 59.5399
R1337 B.n81 B.n80 59.5399
R1338 B.n241 B.n177 59.5399
R1339 B.n171 B.n170 59.5399
R1340 B.n121 B.t2 49.3976
R1341 B.t0 B.n603 49.3976
R1342 B.t6 B.n105 47.5681
R1343 B.t3 B.n15 47.5681
R1344 B.n145 B.t13 43.909
R1345 B.t9 B.n579 43.909
R1346 B.n393 B.t5 42.0795
R1347 B.n620 B.t1 42.0795
R1348 B.n356 B.t4 40.25
R1349 B.n596 B.t7 40.25
R1350 B.n312 B.n311 30.1273
R1351 B.n316 B.n151 30.1273
R1352 B.n568 B.n567 30.1273
R1353 B.n446 B.n443 30.1273
R1354 B.n72 B.n71 29.2853
R1355 B.n80 B.n79 29.2853
R1356 B.n177 B.n176 29.2853
R1357 B.n170 B.n169 29.2853
R1358 B.n129 B.t4 21.9548
R1359 B.t7 B.n595 21.9548
R1360 B.t5 B.n97 20.1252
R1361 B.n408 B.t1 20.1252
R1362 B.n332 B.t13 18.2957
R1363 B.n580 B.t9 18.2957
R1364 B B.n632 18.0485
R1365 B.n380 B.t6 14.6367
R1366 B.n612 B.t3 14.6367
R1367 B.n368 B.t2 12.8072
R1368 B.n604 B.t0 12.8072
R1369 B.n312 B.n147 10.6151
R1370 B.n322 B.n147 10.6151
R1371 B.n323 B.n322 10.6151
R1372 B.n324 B.n323 10.6151
R1373 B.n324 B.n139 10.6151
R1374 B.n334 B.n139 10.6151
R1375 B.n335 B.n334 10.6151
R1376 B.n336 B.n335 10.6151
R1377 B.n336 B.n131 10.6151
R1378 B.n346 B.n131 10.6151
R1379 B.n347 B.n346 10.6151
R1380 B.n348 B.n347 10.6151
R1381 B.n348 B.n123 10.6151
R1382 B.n358 B.n123 10.6151
R1383 B.n359 B.n358 10.6151
R1384 B.n360 B.n359 10.6151
R1385 B.n360 B.n115 10.6151
R1386 B.n370 B.n115 10.6151
R1387 B.n371 B.n370 10.6151
R1388 B.n372 B.n371 10.6151
R1389 B.n372 B.n107 10.6151
R1390 B.n382 B.n107 10.6151
R1391 B.n383 B.n382 10.6151
R1392 B.n384 B.n383 10.6151
R1393 B.n384 B.n99 10.6151
R1394 B.n395 B.n99 10.6151
R1395 B.n396 B.n395 10.6151
R1396 B.n397 B.n396 10.6151
R1397 B.n397 B.n0 10.6151
R1398 B.n311 B.n310 10.6151
R1399 B.n310 B.n155 10.6151
R1400 B.n305 B.n155 10.6151
R1401 B.n305 B.n304 10.6151
R1402 B.n304 B.n157 10.6151
R1403 B.n299 B.n157 10.6151
R1404 B.n299 B.n298 10.6151
R1405 B.n298 B.n297 10.6151
R1406 B.n297 B.n159 10.6151
R1407 B.n291 B.n159 10.6151
R1408 B.n291 B.n290 10.6151
R1409 B.n290 B.n289 10.6151
R1410 B.n289 B.n161 10.6151
R1411 B.n283 B.n161 10.6151
R1412 B.n283 B.n282 10.6151
R1413 B.n282 B.n281 10.6151
R1414 B.n281 B.n163 10.6151
R1415 B.n275 B.n163 10.6151
R1416 B.n275 B.n274 10.6151
R1417 B.n274 B.n273 10.6151
R1418 B.n273 B.n165 10.6151
R1419 B.n267 B.n165 10.6151
R1420 B.n267 B.n266 10.6151
R1421 B.n266 B.n265 10.6151
R1422 B.n265 B.n167 10.6151
R1423 B.n259 B.n258 10.6151
R1424 B.n258 B.n257 10.6151
R1425 B.n257 B.n172 10.6151
R1426 B.n251 B.n172 10.6151
R1427 B.n251 B.n250 10.6151
R1428 B.n250 B.n249 10.6151
R1429 B.n249 B.n174 10.6151
R1430 B.n243 B.n174 10.6151
R1431 B.n243 B.n242 10.6151
R1432 B.n240 B.n178 10.6151
R1433 B.n234 B.n178 10.6151
R1434 B.n234 B.n233 10.6151
R1435 B.n233 B.n232 10.6151
R1436 B.n232 B.n180 10.6151
R1437 B.n226 B.n180 10.6151
R1438 B.n226 B.n225 10.6151
R1439 B.n225 B.n224 10.6151
R1440 B.n224 B.n182 10.6151
R1441 B.n218 B.n182 10.6151
R1442 B.n218 B.n217 10.6151
R1443 B.n217 B.n216 10.6151
R1444 B.n216 B.n184 10.6151
R1445 B.n210 B.n184 10.6151
R1446 B.n210 B.n209 10.6151
R1447 B.n209 B.n208 10.6151
R1448 B.n208 B.n186 10.6151
R1449 B.n202 B.n186 10.6151
R1450 B.n202 B.n201 10.6151
R1451 B.n201 B.n200 10.6151
R1452 B.n200 B.n188 10.6151
R1453 B.n194 B.n188 10.6151
R1454 B.n194 B.n193 10.6151
R1455 B.n193 B.n192 10.6151
R1456 B.n192 B.n151 10.6151
R1457 B.n317 B.n316 10.6151
R1458 B.n318 B.n317 10.6151
R1459 B.n318 B.n142 10.6151
R1460 B.n328 B.n142 10.6151
R1461 B.n329 B.n328 10.6151
R1462 B.n330 B.n329 10.6151
R1463 B.n330 B.n135 10.6151
R1464 B.n340 B.n135 10.6151
R1465 B.n341 B.n340 10.6151
R1466 B.n342 B.n341 10.6151
R1467 B.n342 B.n126 10.6151
R1468 B.n352 B.n126 10.6151
R1469 B.n353 B.n352 10.6151
R1470 B.n354 B.n353 10.6151
R1471 B.n354 B.n118 10.6151
R1472 B.n364 B.n118 10.6151
R1473 B.n365 B.n364 10.6151
R1474 B.n366 B.n365 10.6151
R1475 B.n366 B.n111 10.6151
R1476 B.n376 B.n111 10.6151
R1477 B.n377 B.n376 10.6151
R1478 B.n378 B.n377 10.6151
R1479 B.n378 B.n103 10.6151
R1480 B.n388 B.n103 10.6151
R1481 B.n389 B.n388 10.6151
R1482 B.n391 B.n389 10.6151
R1483 B.n391 B.n390 10.6151
R1484 B.n390 B.n95 10.6151
R1485 B.n402 B.n95 10.6151
R1486 B.n403 B.n402 10.6151
R1487 B.n404 B.n403 10.6151
R1488 B.n405 B.n404 10.6151
R1489 B.n406 B.n405 10.6151
R1490 B.n410 B.n406 10.6151
R1491 B.n411 B.n410 10.6151
R1492 B.n412 B.n411 10.6151
R1493 B.n413 B.n412 10.6151
R1494 B.n415 B.n413 10.6151
R1495 B.n416 B.n415 10.6151
R1496 B.n417 B.n416 10.6151
R1497 B.n418 B.n417 10.6151
R1498 B.n420 B.n418 10.6151
R1499 B.n421 B.n420 10.6151
R1500 B.n422 B.n421 10.6151
R1501 B.n423 B.n422 10.6151
R1502 B.n425 B.n423 10.6151
R1503 B.n426 B.n425 10.6151
R1504 B.n427 B.n426 10.6151
R1505 B.n428 B.n427 10.6151
R1506 B.n430 B.n428 10.6151
R1507 B.n431 B.n430 10.6151
R1508 B.n432 B.n431 10.6151
R1509 B.n433 B.n432 10.6151
R1510 B.n435 B.n433 10.6151
R1511 B.n436 B.n435 10.6151
R1512 B.n437 B.n436 10.6151
R1513 B.n438 B.n437 10.6151
R1514 B.n440 B.n438 10.6151
R1515 B.n441 B.n440 10.6151
R1516 B.n442 B.n441 10.6151
R1517 B.n443 B.n442 10.6151
R1518 B.n624 B.n1 10.6151
R1519 B.n624 B.n623 10.6151
R1520 B.n623 B.n622 10.6151
R1521 B.n622 B.n10 10.6151
R1522 B.n616 B.n10 10.6151
R1523 B.n616 B.n615 10.6151
R1524 B.n615 B.n614 10.6151
R1525 B.n614 B.n17 10.6151
R1526 B.n608 B.n17 10.6151
R1527 B.n608 B.n607 10.6151
R1528 B.n607 B.n606 10.6151
R1529 B.n606 B.n24 10.6151
R1530 B.n600 B.n24 10.6151
R1531 B.n600 B.n599 10.6151
R1532 B.n599 B.n598 10.6151
R1533 B.n598 B.n31 10.6151
R1534 B.n592 B.n31 10.6151
R1535 B.n592 B.n591 10.6151
R1536 B.n591 B.n590 10.6151
R1537 B.n590 B.n38 10.6151
R1538 B.n584 B.n38 10.6151
R1539 B.n584 B.n583 10.6151
R1540 B.n583 B.n582 10.6151
R1541 B.n582 B.n45 10.6151
R1542 B.n576 B.n45 10.6151
R1543 B.n576 B.n575 10.6151
R1544 B.n575 B.n574 10.6151
R1545 B.n574 B.n52 10.6151
R1546 B.n568 B.n52 10.6151
R1547 B.n567 B.n566 10.6151
R1548 B.n566 B.n59 10.6151
R1549 B.n560 B.n59 10.6151
R1550 B.n560 B.n559 10.6151
R1551 B.n559 B.n558 10.6151
R1552 B.n558 B.n61 10.6151
R1553 B.n552 B.n61 10.6151
R1554 B.n552 B.n551 10.6151
R1555 B.n551 B.n550 10.6151
R1556 B.n550 B.n63 10.6151
R1557 B.n544 B.n63 10.6151
R1558 B.n544 B.n543 10.6151
R1559 B.n543 B.n542 10.6151
R1560 B.n542 B.n65 10.6151
R1561 B.n536 B.n65 10.6151
R1562 B.n536 B.n535 10.6151
R1563 B.n535 B.n534 10.6151
R1564 B.n534 B.n67 10.6151
R1565 B.n528 B.n67 10.6151
R1566 B.n528 B.n527 10.6151
R1567 B.n527 B.n526 10.6151
R1568 B.n526 B.n69 10.6151
R1569 B.n520 B.n69 10.6151
R1570 B.n520 B.n519 10.6151
R1571 B.n519 B.n518 10.6151
R1572 B.n514 B.n513 10.6151
R1573 B.n513 B.n75 10.6151
R1574 B.n508 B.n75 10.6151
R1575 B.n508 B.n507 10.6151
R1576 B.n507 B.n506 10.6151
R1577 B.n506 B.n77 10.6151
R1578 B.n500 B.n77 10.6151
R1579 B.n500 B.n499 10.6151
R1580 B.n499 B.n498 10.6151
R1581 B.n494 B.n493 10.6151
R1582 B.n493 B.n83 10.6151
R1583 B.n488 B.n83 10.6151
R1584 B.n488 B.n487 10.6151
R1585 B.n487 B.n486 10.6151
R1586 B.n486 B.n85 10.6151
R1587 B.n480 B.n85 10.6151
R1588 B.n480 B.n479 10.6151
R1589 B.n479 B.n478 10.6151
R1590 B.n478 B.n87 10.6151
R1591 B.n472 B.n87 10.6151
R1592 B.n472 B.n471 10.6151
R1593 B.n471 B.n470 10.6151
R1594 B.n470 B.n89 10.6151
R1595 B.n464 B.n89 10.6151
R1596 B.n464 B.n463 10.6151
R1597 B.n463 B.n462 10.6151
R1598 B.n462 B.n91 10.6151
R1599 B.n456 B.n91 10.6151
R1600 B.n456 B.n455 10.6151
R1601 B.n455 B.n454 10.6151
R1602 B.n454 B.n93 10.6151
R1603 B.n448 B.n93 10.6151
R1604 B.n448 B.n447 10.6151
R1605 B.n447 B.n446 10.6151
R1606 B.n171 B.n167 9.36635
R1607 B.n241 B.n240 9.36635
R1608 B.n518 B.n73 9.36635
R1609 B.n494 B.n81 9.36635
R1610 B.n632 B.n0 8.11757
R1611 B.n632 B.n1 8.11757
R1612 B.n259 B.n171 1.24928
R1613 B.n242 B.n241 1.24928
R1614 B.n514 B.n73 1.24928
R1615 B.n498 B.n81 1.24928
R1616 VP.n23 VP.n5 172.799
R1617 VP.n40 VP.n39 172.799
R1618 VP.n22 VP.n21 172.799
R1619 VP.n10 VP.t1 168.466
R1620 VP.n12 VP.n11 161.3
R1621 VP.n13 VP.n8 161.3
R1622 VP.n16 VP.n15 161.3
R1623 VP.n17 VP.n7 161.3
R1624 VP.n19 VP.n18 161.3
R1625 VP.n20 VP.n6 161.3
R1626 VP.n38 VP.n0 161.3
R1627 VP.n37 VP.n36 161.3
R1628 VP.n35 VP.n1 161.3
R1629 VP.n34 VP.n33 161.3
R1630 VP.n31 VP.n2 161.3
R1631 VP.n30 VP.n29 161.3
R1632 VP.n28 VP.n27 161.3
R1633 VP.n26 VP.n4 161.3
R1634 VP.n25 VP.n24 161.3
R1635 VP.n5 VP.t5 137.861
R1636 VP.n3 VP.t7 137.861
R1637 VP.n32 VP.t4 137.861
R1638 VP.n39 VP.t2 137.861
R1639 VP.n21 VP.t3 137.861
R1640 VP.n14 VP.t0 137.861
R1641 VP.n9 VP.t6 137.861
R1642 VP.n10 VP.n9 51.0709
R1643 VP.n26 VP.n25 41.4647
R1644 VP.n38 VP.n37 41.4647
R1645 VP.n20 VP.n19 41.4647
R1646 VP.n31 VP.n30 40.4934
R1647 VP.n33 VP.n31 40.4934
R1648 VP.n15 VP.n13 40.4934
R1649 VP.n13 VP.n12 40.4934
R1650 VP.n23 VP.n22 40.1672
R1651 VP.n27 VP.n26 39.5221
R1652 VP.n37 VP.n1 39.5221
R1653 VP.n19 VP.n7 39.5221
R1654 VP.n11 VP.n10 26.8925
R1655 VP.n25 VP.n5 12.968
R1656 VP.n39 VP.n38 12.968
R1657 VP.n21 VP.n20 12.968
R1658 VP.n30 VP.n3 12.4787
R1659 VP.n33 VP.n32 12.4787
R1660 VP.n15 VP.n14 12.4787
R1661 VP.n12 VP.n9 12.4787
R1662 VP.n27 VP.n3 11.9893
R1663 VP.n32 VP.n1 11.9893
R1664 VP.n14 VP.n7 11.9893
R1665 VP.n11 VP.n8 0.189894
R1666 VP.n16 VP.n8 0.189894
R1667 VP.n17 VP.n16 0.189894
R1668 VP.n18 VP.n17 0.189894
R1669 VP.n18 VP.n6 0.189894
R1670 VP.n22 VP.n6 0.189894
R1671 VP.n24 VP.n23 0.189894
R1672 VP.n24 VP.n4 0.189894
R1673 VP.n28 VP.n4 0.189894
R1674 VP.n29 VP.n28 0.189894
R1675 VP.n29 VP.n2 0.189894
R1676 VP.n34 VP.n2 0.189894
R1677 VP.n35 VP.n34 0.189894
R1678 VP.n36 VP.n35 0.189894
R1679 VP.n36 VP.n0 0.189894
R1680 VP.n40 VP.n0 0.189894
R1681 VP VP.n40 0.0516364
R1682 VDD1 VDD1.n0 67.365
R1683 VDD1.n3 VDD1.n2 67.2513
R1684 VDD1.n3 VDD1.n1 67.2513
R1685 VDD1.n5 VDD1.n4 66.6558
R1686 VDD1.n5 VDD1.n3 35.975
R1687 VDD1.n4 VDD1.t7 2.93383
R1688 VDD1.n4 VDD1.t4 2.93383
R1689 VDD1.n0 VDD1.t6 2.93383
R1690 VDD1.n0 VDD1.t1 2.93383
R1691 VDD1.n2 VDD1.t3 2.93383
R1692 VDD1.n2 VDD1.t5 2.93383
R1693 VDD1.n1 VDD1.t2 2.93383
R1694 VDD1.n1 VDD1.t0 2.93383
R1695 VDD1 VDD1.n5 0.593172
C0 VDD2 VP 0.36806f
C1 VTAIL VN 4.32696f
C2 VTAIL VDD1 6.22096f
C3 VDD1 VN 0.148653f
C4 VTAIL VP 4.34106f
C5 VP VN 4.956491f
C6 VP VDD1 4.32263f
C7 VDD2 VTAIL 6.26586f
C8 VDD2 VN 4.1039f
C9 VDD2 VDD1 1.06294f
C10 VDD2 B 3.53502f
C11 VDD1 B 3.817887f
C12 VTAIL B 6.148151f
C13 VN B 9.609029f
C14 VP B 8.057651f
C15 VDD1.t6 B 0.135595f
C16 VDD1.t1 B 0.135595f
C17 VDD1.n0 B 1.15064f
C18 VDD1.t2 B 0.135595f
C19 VDD1.t0 B 0.135595f
C20 VDD1.n1 B 1.14992f
C21 VDD1.t3 B 0.135595f
C22 VDD1.t5 B 0.135595f
C23 VDD1.n2 B 1.14992f
C24 VDD1.n3 B 2.22292f
C25 VDD1.t7 B 0.135595f
C26 VDD1.t4 B 0.135595f
C27 VDD1.n4 B 1.1466f
C28 VDD1.n5 B 2.10944f
C29 VP.n0 B 0.037293f
C30 VP.t2 B 0.79133f
C31 VP.n1 B 0.056967f
C32 VP.n2 B 0.037293f
C33 VP.t7 B 0.79133f
C34 VP.n3 B 0.311791f
C35 VP.n4 B 0.037293f
C36 VP.t5 B 0.79133f
C37 VP.n5 B 0.373145f
C38 VP.n6 B 0.037293f
C39 VP.t3 B 0.79133f
C40 VP.n7 B 0.056967f
C41 VP.n8 B 0.037293f
C42 VP.t6 B 0.79133f
C43 VP.n9 B 0.366897f
C44 VP.t1 B 0.867856f
C45 VP.n10 B 0.388133f
C46 VP.n11 B 0.193801f
C47 VP.n12 B 0.057303f
C48 VP.n13 B 0.030148f
C49 VP.t0 B 0.79133f
C50 VP.n14 B 0.311791f
C51 VP.n15 B 0.057303f
C52 VP.n16 B 0.037293f
C53 VP.n17 B 0.037293f
C54 VP.n18 B 0.037293f
C55 VP.n19 B 0.030196f
C56 VP.n20 B 0.057592f
C57 VP.n21 B 0.373145f
C58 VP.n22 B 1.43173f
C59 VP.n23 B 1.4651f
C60 VP.n24 B 0.037293f
C61 VP.n25 B 0.057592f
C62 VP.n26 B 0.030196f
C63 VP.n27 B 0.056967f
C64 VP.n28 B 0.037293f
C65 VP.n29 B 0.037293f
C66 VP.n30 B 0.057303f
C67 VP.n31 B 0.030148f
C68 VP.t4 B 0.79133f
C69 VP.n32 B 0.311791f
C70 VP.n33 B 0.057303f
C71 VP.n34 B 0.037293f
C72 VP.n35 B 0.037293f
C73 VP.n36 B 0.037293f
C74 VP.n37 B 0.030196f
C75 VP.n38 B 0.057592f
C76 VP.n39 B 0.373145f
C77 VP.n40 B 0.033275f
C78 VTAIL.t10 B 0.112368f
C79 VTAIL.t15 B 0.112368f
C80 VTAIL.n0 B 0.893925f
C81 VTAIL.n1 B 0.292554f
C82 VTAIL.n2 B 0.030605f
C83 VTAIL.n3 B 0.021066f
C84 VTAIL.n4 B 0.01132f
C85 VTAIL.n5 B 0.026756f
C86 VTAIL.n6 B 0.011986f
C87 VTAIL.n7 B 0.021066f
C88 VTAIL.n8 B 0.01132f
C89 VTAIL.n9 B 0.026756f
C90 VTAIL.n10 B 0.011986f
C91 VTAIL.n11 B 0.573842f
C92 VTAIL.n12 B 0.01132f
C93 VTAIL.t14 B 0.043601f
C94 VTAIL.n13 B 0.093987f
C95 VTAIL.n14 B 0.015806f
C96 VTAIL.n15 B 0.020067f
C97 VTAIL.n16 B 0.026756f
C98 VTAIL.n17 B 0.011986f
C99 VTAIL.n18 B 0.01132f
C100 VTAIL.n19 B 0.021066f
C101 VTAIL.n20 B 0.021066f
C102 VTAIL.n21 B 0.01132f
C103 VTAIL.n22 B 0.011986f
C104 VTAIL.n23 B 0.026756f
C105 VTAIL.n24 B 0.026756f
C106 VTAIL.n25 B 0.011986f
C107 VTAIL.n26 B 0.01132f
C108 VTAIL.n27 B 0.021066f
C109 VTAIL.n28 B 0.021066f
C110 VTAIL.n29 B 0.01132f
C111 VTAIL.n30 B 0.011986f
C112 VTAIL.n31 B 0.026756f
C113 VTAIL.n32 B 0.059682f
C114 VTAIL.n33 B 0.011986f
C115 VTAIL.n34 B 0.01132f
C116 VTAIL.n35 B 0.049557f
C117 VTAIL.n36 B 0.033602f
C118 VTAIL.n37 B 0.138732f
C119 VTAIL.n38 B 0.030605f
C120 VTAIL.n39 B 0.021066f
C121 VTAIL.n40 B 0.01132f
C122 VTAIL.n41 B 0.026756f
C123 VTAIL.n42 B 0.011986f
C124 VTAIL.n43 B 0.021066f
C125 VTAIL.n44 B 0.01132f
C126 VTAIL.n45 B 0.026756f
C127 VTAIL.n46 B 0.011986f
C128 VTAIL.n47 B 0.573842f
C129 VTAIL.n48 B 0.01132f
C130 VTAIL.t5 B 0.043601f
C131 VTAIL.n49 B 0.093987f
C132 VTAIL.n50 B 0.015806f
C133 VTAIL.n51 B 0.020067f
C134 VTAIL.n52 B 0.026756f
C135 VTAIL.n53 B 0.011986f
C136 VTAIL.n54 B 0.01132f
C137 VTAIL.n55 B 0.021066f
C138 VTAIL.n56 B 0.021066f
C139 VTAIL.n57 B 0.01132f
C140 VTAIL.n58 B 0.011986f
C141 VTAIL.n59 B 0.026756f
C142 VTAIL.n60 B 0.026756f
C143 VTAIL.n61 B 0.011986f
C144 VTAIL.n62 B 0.01132f
C145 VTAIL.n63 B 0.021066f
C146 VTAIL.n64 B 0.021066f
C147 VTAIL.n65 B 0.01132f
C148 VTAIL.n66 B 0.011986f
C149 VTAIL.n67 B 0.026756f
C150 VTAIL.n68 B 0.059682f
C151 VTAIL.n69 B 0.011986f
C152 VTAIL.n70 B 0.01132f
C153 VTAIL.n71 B 0.049557f
C154 VTAIL.n72 B 0.033602f
C155 VTAIL.n73 B 0.138732f
C156 VTAIL.t2 B 0.112368f
C157 VTAIL.t6 B 0.112368f
C158 VTAIL.n74 B 0.893925f
C159 VTAIL.n75 B 0.376965f
C160 VTAIL.n76 B 0.030605f
C161 VTAIL.n77 B 0.021066f
C162 VTAIL.n78 B 0.01132f
C163 VTAIL.n79 B 0.026756f
C164 VTAIL.n80 B 0.011986f
C165 VTAIL.n81 B 0.021066f
C166 VTAIL.n82 B 0.01132f
C167 VTAIL.n83 B 0.026756f
C168 VTAIL.n84 B 0.011986f
C169 VTAIL.n85 B 0.573842f
C170 VTAIL.n86 B 0.01132f
C171 VTAIL.t4 B 0.043601f
C172 VTAIL.n87 B 0.093987f
C173 VTAIL.n88 B 0.015806f
C174 VTAIL.n89 B 0.020067f
C175 VTAIL.n90 B 0.026756f
C176 VTAIL.n91 B 0.011986f
C177 VTAIL.n92 B 0.01132f
C178 VTAIL.n93 B 0.021066f
C179 VTAIL.n94 B 0.021066f
C180 VTAIL.n95 B 0.01132f
C181 VTAIL.n96 B 0.011986f
C182 VTAIL.n97 B 0.026756f
C183 VTAIL.n98 B 0.026756f
C184 VTAIL.n99 B 0.011986f
C185 VTAIL.n100 B 0.01132f
C186 VTAIL.n101 B 0.021066f
C187 VTAIL.n102 B 0.021066f
C188 VTAIL.n103 B 0.01132f
C189 VTAIL.n104 B 0.011986f
C190 VTAIL.n105 B 0.026756f
C191 VTAIL.n106 B 0.059682f
C192 VTAIL.n107 B 0.011986f
C193 VTAIL.n108 B 0.01132f
C194 VTAIL.n109 B 0.049557f
C195 VTAIL.n110 B 0.033602f
C196 VTAIL.n111 B 0.87635f
C197 VTAIL.n112 B 0.030605f
C198 VTAIL.n113 B 0.021066f
C199 VTAIL.n114 B 0.01132f
C200 VTAIL.n115 B 0.026756f
C201 VTAIL.n116 B 0.011986f
C202 VTAIL.n117 B 0.021066f
C203 VTAIL.n118 B 0.01132f
C204 VTAIL.n119 B 0.026756f
C205 VTAIL.n120 B 0.011986f
C206 VTAIL.n121 B 0.573842f
C207 VTAIL.n122 B 0.01132f
C208 VTAIL.t12 B 0.043601f
C209 VTAIL.n123 B 0.093987f
C210 VTAIL.n124 B 0.015806f
C211 VTAIL.n125 B 0.020067f
C212 VTAIL.n126 B 0.026756f
C213 VTAIL.n127 B 0.011986f
C214 VTAIL.n128 B 0.01132f
C215 VTAIL.n129 B 0.021066f
C216 VTAIL.n130 B 0.021066f
C217 VTAIL.n131 B 0.01132f
C218 VTAIL.n132 B 0.011986f
C219 VTAIL.n133 B 0.026756f
C220 VTAIL.n134 B 0.026756f
C221 VTAIL.n135 B 0.011986f
C222 VTAIL.n136 B 0.01132f
C223 VTAIL.n137 B 0.021066f
C224 VTAIL.n138 B 0.021066f
C225 VTAIL.n139 B 0.01132f
C226 VTAIL.n140 B 0.011986f
C227 VTAIL.n141 B 0.026756f
C228 VTAIL.n142 B 0.059682f
C229 VTAIL.n143 B 0.011986f
C230 VTAIL.n144 B 0.01132f
C231 VTAIL.n145 B 0.049557f
C232 VTAIL.n146 B 0.033602f
C233 VTAIL.n147 B 0.87635f
C234 VTAIL.t9 B 0.112368f
C235 VTAIL.t13 B 0.112368f
C236 VTAIL.n148 B 0.893931f
C237 VTAIL.n149 B 0.376959f
C238 VTAIL.n150 B 0.030605f
C239 VTAIL.n151 B 0.021066f
C240 VTAIL.n152 B 0.01132f
C241 VTAIL.n153 B 0.026756f
C242 VTAIL.n154 B 0.011986f
C243 VTAIL.n155 B 0.021066f
C244 VTAIL.n156 B 0.01132f
C245 VTAIL.n157 B 0.026756f
C246 VTAIL.n158 B 0.011986f
C247 VTAIL.n159 B 0.573842f
C248 VTAIL.n160 B 0.01132f
C249 VTAIL.t8 B 0.043601f
C250 VTAIL.n161 B 0.093987f
C251 VTAIL.n162 B 0.015806f
C252 VTAIL.n163 B 0.020067f
C253 VTAIL.n164 B 0.026756f
C254 VTAIL.n165 B 0.011986f
C255 VTAIL.n166 B 0.01132f
C256 VTAIL.n167 B 0.021066f
C257 VTAIL.n168 B 0.021066f
C258 VTAIL.n169 B 0.01132f
C259 VTAIL.n170 B 0.011986f
C260 VTAIL.n171 B 0.026756f
C261 VTAIL.n172 B 0.026756f
C262 VTAIL.n173 B 0.011986f
C263 VTAIL.n174 B 0.01132f
C264 VTAIL.n175 B 0.021066f
C265 VTAIL.n176 B 0.021066f
C266 VTAIL.n177 B 0.01132f
C267 VTAIL.n178 B 0.011986f
C268 VTAIL.n179 B 0.026756f
C269 VTAIL.n180 B 0.059682f
C270 VTAIL.n181 B 0.011986f
C271 VTAIL.n182 B 0.01132f
C272 VTAIL.n183 B 0.049557f
C273 VTAIL.n184 B 0.033602f
C274 VTAIL.n185 B 0.138732f
C275 VTAIL.n186 B 0.030605f
C276 VTAIL.n187 B 0.021066f
C277 VTAIL.n188 B 0.01132f
C278 VTAIL.n189 B 0.026756f
C279 VTAIL.n190 B 0.011986f
C280 VTAIL.n191 B 0.021066f
C281 VTAIL.n192 B 0.01132f
C282 VTAIL.n193 B 0.026756f
C283 VTAIL.n194 B 0.011986f
C284 VTAIL.n195 B 0.573842f
C285 VTAIL.n196 B 0.01132f
C286 VTAIL.t1 B 0.043601f
C287 VTAIL.n197 B 0.093987f
C288 VTAIL.n198 B 0.015806f
C289 VTAIL.n199 B 0.020067f
C290 VTAIL.n200 B 0.026756f
C291 VTAIL.n201 B 0.011986f
C292 VTAIL.n202 B 0.01132f
C293 VTAIL.n203 B 0.021066f
C294 VTAIL.n204 B 0.021066f
C295 VTAIL.n205 B 0.01132f
C296 VTAIL.n206 B 0.011986f
C297 VTAIL.n207 B 0.026756f
C298 VTAIL.n208 B 0.026756f
C299 VTAIL.n209 B 0.011986f
C300 VTAIL.n210 B 0.01132f
C301 VTAIL.n211 B 0.021066f
C302 VTAIL.n212 B 0.021066f
C303 VTAIL.n213 B 0.01132f
C304 VTAIL.n214 B 0.011986f
C305 VTAIL.n215 B 0.026756f
C306 VTAIL.n216 B 0.059682f
C307 VTAIL.n217 B 0.011986f
C308 VTAIL.n218 B 0.01132f
C309 VTAIL.n219 B 0.049557f
C310 VTAIL.n220 B 0.033602f
C311 VTAIL.n221 B 0.138732f
C312 VTAIL.t3 B 0.112368f
C313 VTAIL.t0 B 0.112368f
C314 VTAIL.n222 B 0.893931f
C315 VTAIL.n223 B 0.376959f
C316 VTAIL.n224 B 0.030605f
C317 VTAIL.n225 B 0.021066f
C318 VTAIL.n226 B 0.01132f
C319 VTAIL.n227 B 0.026756f
C320 VTAIL.n228 B 0.011986f
C321 VTAIL.n229 B 0.021066f
C322 VTAIL.n230 B 0.01132f
C323 VTAIL.n231 B 0.026756f
C324 VTAIL.n232 B 0.011986f
C325 VTAIL.n233 B 0.573842f
C326 VTAIL.n234 B 0.01132f
C327 VTAIL.t7 B 0.043601f
C328 VTAIL.n235 B 0.093987f
C329 VTAIL.n236 B 0.015806f
C330 VTAIL.n237 B 0.020067f
C331 VTAIL.n238 B 0.026756f
C332 VTAIL.n239 B 0.011986f
C333 VTAIL.n240 B 0.01132f
C334 VTAIL.n241 B 0.021066f
C335 VTAIL.n242 B 0.021066f
C336 VTAIL.n243 B 0.01132f
C337 VTAIL.n244 B 0.011986f
C338 VTAIL.n245 B 0.026756f
C339 VTAIL.n246 B 0.026756f
C340 VTAIL.n247 B 0.011986f
C341 VTAIL.n248 B 0.01132f
C342 VTAIL.n249 B 0.021066f
C343 VTAIL.n250 B 0.021066f
C344 VTAIL.n251 B 0.01132f
C345 VTAIL.n252 B 0.011986f
C346 VTAIL.n253 B 0.026756f
C347 VTAIL.n254 B 0.059682f
C348 VTAIL.n255 B 0.011986f
C349 VTAIL.n256 B 0.01132f
C350 VTAIL.n257 B 0.049557f
C351 VTAIL.n258 B 0.033602f
C352 VTAIL.n259 B 0.87635f
C353 VTAIL.n260 B 0.030605f
C354 VTAIL.n261 B 0.021066f
C355 VTAIL.n262 B 0.01132f
C356 VTAIL.n263 B 0.026756f
C357 VTAIL.n264 B 0.011986f
C358 VTAIL.n265 B 0.021066f
C359 VTAIL.n266 B 0.01132f
C360 VTAIL.n267 B 0.026756f
C361 VTAIL.n268 B 0.011986f
C362 VTAIL.n269 B 0.573842f
C363 VTAIL.n270 B 0.01132f
C364 VTAIL.t11 B 0.043601f
C365 VTAIL.n271 B 0.093987f
C366 VTAIL.n272 B 0.015806f
C367 VTAIL.n273 B 0.020067f
C368 VTAIL.n274 B 0.026756f
C369 VTAIL.n275 B 0.011986f
C370 VTAIL.n276 B 0.01132f
C371 VTAIL.n277 B 0.021066f
C372 VTAIL.n278 B 0.021066f
C373 VTAIL.n279 B 0.01132f
C374 VTAIL.n280 B 0.011986f
C375 VTAIL.n281 B 0.026756f
C376 VTAIL.n282 B 0.026756f
C377 VTAIL.n283 B 0.011986f
C378 VTAIL.n284 B 0.01132f
C379 VTAIL.n285 B 0.021066f
C380 VTAIL.n286 B 0.021066f
C381 VTAIL.n287 B 0.01132f
C382 VTAIL.n288 B 0.011986f
C383 VTAIL.n289 B 0.026756f
C384 VTAIL.n290 B 0.059682f
C385 VTAIL.n291 B 0.011986f
C386 VTAIL.n292 B 0.01132f
C387 VTAIL.n293 B 0.049557f
C388 VTAIL.n294 B 0.033602f
C389 VTAIL.n295 B 0.8724f
C390 VDD2.t7 B 0.135515f
C391 VDD2.t4 B 0.135515f
C392 VDD2.n0 B 1.14924f
C393 VDD2.t0 B 0.135515f
C394 VDD2.t6 B 0.135515f
C395 VDD2.n1 B 1.14924f
C396 VDD2.n2 B 2.16757f
C397 VDD2.t5 B 0.135515f
C398 VDD2.t3 B 0.135515f
C399 VDD2.n3 B 1.14593f
C400 VDD2.n4 B 2.07793f
C401 VDD2.t1 B 0.135515f
C402 VDD2.t2 B 0.135515f
C403 VDD2.n5 B 1.14922f
C404 VN.n0 B 0.036603f
C405 VN.t4 B 0.776699f
C406 VN.n1 B 0.055913f
C407 VN.n2 B 0.036603f
C408 VN.t5 B 0.776699f
C409 VN.n3 B 0.360113f
C410 VN.t1 B 0.85181f
C411 VN.n4 B 0.380957f
C412 VN.n5 B 0.190218f
C413 VN.n6 B 0.056244f
C414 VN.n7 B 0.02959f
C415 VN.t0 B 0.776699f
C416 VN.n8 B 0.306026f
C417 VN.n9 B 0.056244f
C418 VN.n10 B 0.036603f
C419 VN.n11 B 0.036603f
C420 VN.n12 B 0.036603f
C421 VN.n13 B 0.029637f
C422 VN.n14 B 0.056527f
C423 VN.n15 B 0.366246f
C424 VN.n16 B 0.032659f
C425 VN.n17 B 0.036603f
C426 VN.t3 B 0.776699f
C427 VN.n18 B 0.055913f
C428 VN.n19 B 0.036603f
C429 VN.t6 B 0.776699f
C430 VN.n20 B 0.306026f
C431 VN.t2 B 0.776699f
C432 VN.n21 B 0.360113f
C433 VN.t7 B 0.85181f
C434 VN.n22 B 0.380957f
C435 VN.n23 B 0.190218f
C436 VN.n24 B 0.056244f
C437 VN.n25 B 0.02959f
C438 VN.n26 B 0.056244f
C439 VN.n27 B 0.036603f
C440 VN.n28 B 0.036603f
C441 VN.n29 B 0.036603f
C442 VN.n30 B 0.029637f
C443 VN.n31 B 0.056527f
C444 VN.n32 B 0.366246f
C445 VN.n33 B 1.42935f
.ends

