* NGSPICE file created from diff_pair_sample_1260.ext - technology: sky130A

.subckt diff_pair_sample_1260 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=0 ps=0 w=7.14 l=0.56
X1 VDD1.t9 VP.t0 VTAIL.t10 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=1.1781 ps=7.47 w=7.14 l=0.56
X2 B.t8 B.t6 B.t7 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=0 ps=0 w=7.14 l=0.56
X3 VDD1.t8 VP.t1 VTAIL.t15 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=2.7846 ps=15.06 w=7.14 l=0.56
X4 VTAIL.t4 VN.t0 VDD2.t9 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X5 VDD2.t8 VN.t1 VTAIL.t3 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=1.1781 ps=7.47 w=7.14 l=0.56
X6 VDD1.t7 VP.t2 VTAIL.t19 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X7 VDD2.t7 VN.t2 VTAIL.t8 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X8 VDD2.t6 VN.t3 VTAIL.t0 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X9 VDD1.t6 VP.t3 VTAIL.t17 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=1.1781 ps=7.47 w=7.14 l=0.56
X10 VDD2.t5 VN.t4 VTAIL.t9 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=2.7846 ps=15.06 w=7.14 l=0.56
X11 VDD2.t4 VN.t5 VTAIL.t2 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=1.1781 ps=7.47 w=7.14 l=0.56
X12 VTAIL.t11 VP.t4 VDD1.t5 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X13 B.t5 B.t3 B.t4 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=0 ps=0 w=7.14 l=0.56
X14 VTAIL.t18 VP.t5 VDD1.t4 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X15 VDD1.t3 VP.t6 VTAIL.t12 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X16 B.t2 B.t0 B.t1 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=2.7846 pd=15.06 as=0 ps=0 w=7.14 l=0.56
X17 VTAIL.t14 VP.t7 VDD1.t2 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X18 VDD2.t3 VN.t6 VTAIL.t1 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=2.7846 ps=15.06 w=7.14 l=0.56
X19 VTAIL.t13 VP.t8 VDD1.t1 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X20 VTAIL.t5 VN.t7 VDD2.t2 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X21 VDD1.t0 VP.t9 VTAIL.t16 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=2.7846 ps=15.06 w=7.14 l=0.56
X22 VTAIL.t6 VN.t8 VDD2.t1 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
X23 VTAIL.t7 VN.t9 VDD2.t0 w_n2038_n2396# sky130_fd_pr__pfet_01v8 ad=1.1781 pd=7.47 as=1.1781 ps=7.47 w=7.14 l=0.56
R0 B.n330 B.n329 585
R1 B.n331 B.n50 585
R2 B.n333 B.n332 585
R3 B.n334 B.n49 585
R4 B.n336 B.n335 585
R5 B.n337 B.n48 585
R6 B.n339 B.n338 585
R7 B.n340 B.n47 585
R8 B.n342 B.n341 585
R9 B.n343 B.n46 585
R10 B.n345 B.n344 585
R11 B.n346 B.n45 585
R12 B.n348 B.n347 585
R13 B.n349 B.n44 585
R14 B.n351 B.n350 585
R15 B.n352 B.n43 585
R16 B.n354 B.n353 585
R17 B.n355 B.n42 585
R18 B.n357 B.n356 585
R19 B.n358 B.n41 585
R20 B.n360 B.n359 585
R21 B.n361 B.n40 585
R22 B.n363 B.n362 585
R23 B.n364 B.n39 585
R24 B.n366 B.n365 585
R25 B.n367 B.n35 585
R26 B.n369 B.n368 585
R27 B.n370 B.n34 585
R28 B.n372 B.n371 585
R29 B.n373 B.n33 585
R30 B.n375 B.n374 585
R31 B.n376 B.n32 585
R32 B.n378 B.n377 585
R33 B.n379 B.n31 585
R34 B.n381 B.n380 585
R35 B.n382 B.n30 585
R36 B.n384 B.n383 585
R37 B.n386 B.n27 585
R38 B.n388 B.n387 585
R39 B.n389 B.n26 585
R40 B.n391 B.n390 585
R41 B.n392 B.n25 585
R42 B.n394 B.n393 585
R43 B.n395 B.n24 585
R44 B.n397 B.n396 585
R45 B.n398 B.n23 585
R46 B.n400 B.n399 585
R47 B.n401 B.n22 585
R48 B.n403 B.n402 585
R49 B.n404 B.n21 585
R50 B.n406 B.n405 585
R51 B.n407 B.n20 585
R52 B.n409 B.n408 585
R53 B.n410 B.n19 585
R54 B.n412 B.n411 585
R55 B.n413 B.n18 585
R56 B.n415 B.n414 585
R57 B.n416 B.n17 585
R58 B.n418 B.n417 585
R59 B.n419 B.n16 585
R60 B.n421 B.n420 585
R61 B.n422 B.n15 585
R62 B.n424 B.n423 585
R63 B.n425 B.n14 585
R64 B.n328 B.n51 585
R65 B.n327 B.n326 585
R66 B.n325 B.n52 585
R67 B.n324 B.n323 585
R68 B.n322 B.n53 585
R69 B.n321 B.n320 585
R70 B.n319 B.n54 585
R71 B.n318 B.n317 585
R72 B.n316 B.n55 585
R73 B.n315 B.n314 585
R74 B.n313 B.n56 585
R75 B.n312 B.n311 585
R76 B.n310 B.n57 585
R77 B.n309 B.n308 585
R78 B.n307 B.n58 585
R79 B.n306 B.n305 585
R80 B.n304 B.n59 585
R81 B.n303 B.n302 585
R82 B.n301 B.n60 585
R83 B.n300 B.n299 585
R84 B.n298 B.n61 585
R85 B.n297 B.n296 585
R86 B.n295 B.n62 585
R87 B.n294 B.n293 585
R88 B.n292 B.n63 585
R89 B.n291 B.n290 585
R90 B.n289 B.n64 585
R91 B.n288 B.n287 585
R92 B.n286 B.n65 585
R93 B.n285 B.n284 585
R94 B.n283 B.n66 585
R95 B.n282 B.n281 585
R96 B.n280 B.n67 585
R97 B.n279 B.n278 585
R98 B.n277 B.n68 585
R99 B.n276 B.n275 585
R100 B.n274 B.n69 585
R101 B.n273 B.n272 585
R102 B.n271 B.n70 585
R103 B.n270 B.n269 585
R104 B.n268 B.n71 585
R105 B.n267 B.n266 585
R106 B.n265 B.n72 585
R107 B.n264 B.n263 585
R108 B.n262 B.n73 585
R109 B.n261 B.n260 585
R110 B.n259 B.n74 585
R111 B.n258 B.n257 585
R112 B.n256 B.n75 585
R113 B.n159 B.n158 585
R114 B.n160 B.n111 585
R115 B.n162 B.n161 585
R116 B.n163 B.n110 585
R117 B.n165 B.n164 585
R118 B.n166 B.n109 585
R119 B.n168 B.n167 585
R120 B.n169 B.n108 585
R121 B.n171 B.n170 585
R122 B.n172 B.n107 585
R123 B.n174 B.n173 585
R124 B.n175 B.n106 585
R125 B.n177 B.n176 585
R126 B.n178 B.n105 585
R127 B.n180 B.n179 585
R128 B.n181 B.n104 585
R129 B.n183 B.n182 585
R130 B.n184 B.n103 585
R131 B.n186 B.n185 585
R132 B.n187 B.n102 585
R133 B.n189 B.n188 585
R134 B.n190 B.n101 585
R135 B.n192 B.n191 585
R136 B.n193 B.n100 585
R137 B.n195 B.n194 585
R138 B.n196 B.n99 585
R139 B.n198 B.n197 585
R140 B.n200 B.n96 585
R141 B.n202 B.n201 585
R142 B.n203 B.n95 585
R143 B.n205 B.n204 585
R144 B.n206 B.n94 585
R145 B.n208 B.n207 585
R146 B.n209 B.n93 585
R147 B.n211 B.n210 585
R148 B.n212 B.n92 585
R149 B.n214 B.n213 585
R150 B.n216 B.n215 585
R151 B.n217 B.n88 585
R152 B.n219 B.n218 585
R153 B.n220 B.n87 585
R154 B.n222 B.n221 585
R155 B.n223 B.n86 585
R156 B.n225 B.n224 585
R157 B.n226 B.n85 585
R158 B.n228 B.n227 585
R159 B.n229 B.n84 585
R160 B.n231 B.n230 585
R161 B.n232 B.n83 585
R162 B.n234 B.n233 585
R163 B.n235 B.n82 585
R164 B.n237 B.n236 585
R165 B.n238 B.n81 585
R166 B.n240 B.n239 585
R167 B.n241 B.n80 585
R168 B.n243 B.n242 585
R169 B.n244 B.n79 585
R170 B.n246 B.n245 585
R171 B.n247 B.n78 585
R172 B.n249 B.n248 585
R173 B.n250 B.n77 585
R174 B.n252 B.n251 585
R175 B.n253 B.n76 585
R176 B.n255 B.n254 585
R177 B.n157 B.n112 585
R178 B.n156 B.n155 585
R179 B.n154 B.n113 585
R180 B.n153 B.n152 585
R181 B.n151 B.n114 585
R182 B.n150 B.n149 585
R183 B.n148 B.n115 585
R184 B.n147 B.n146 585
R185 B.n145 B.n116 585
R186 B.n144 B.n143 585
R187 B.n142 B.n117 585
R188 B.n141 B.n140 585
R189 B.n139 B.n118 585
R190 B.n138 B.n137 585
R191 B.n136 B.n119 585
R192 B.n135 B.n134 585
R193 B.n133 B.n120 585
R194 B.n132 B.n131 585
R195 B.n130 B.n121 585
R196 B.n129 B.n128 585
R197 B.n127 B.n122 585
R198 B.n126 B.n125 585
R199 B.n124 B.n123 585
R200 B.n2 B.n0 585
R201 B.n461 B.n1 585
R202 B.n460 B.n459 585
R203 B.n458 B.n3 585
R204 B.n457 B.n456 585
R205 B.n455 B.n4 585
R206 B.n454 B.n453 585
R207 B.n452 B.n5 585
R208 B.n451 B.n450 585
R209 B.n449 B.n6 585
R210 B.n448 B.n447 585
R211 B.n446 B.n7 585
R212 B.n445 B.n444 585
R213 B.n443 B.n8 585
R214 B.n442 B.n441 585
R215 B.n440 B.n9 585
R216 B.n439 B.n438 585
R217 B.n437 B.n10 585
R218 B.n436 B.n435 585
R219 B.n434 B.n11 585
R220 B.n433 B.n432 585
R221 B.n431 B.n12 585
R222 B.n430 B.n429 585
R223 B.n428 B.n13 585
R224 B.n427 B.n426 585
R225 B.n463 B.n462 585
R226 B.n89 B.t9 512.391
R227 B.n97 B.t0 512.391
R228 B.n28 B.t6 512.391
R229 B.n36 B.t3 512.391
R230 B.n159 B.n112 487.695
R231 B.n426 B.n425 487.695
R232 B.n256 B.n255 487.695
R233 B.n329 B.n328 487.695
R234 B.n155 B.n112 163.367
R235 B.n155 B.n154 163.367
R236 B.n154 B.n153 163.367
R237 B.n153 B.n114 163.367
R238 B.n149 B.n114 163.367
R239 B.n149 B.n148 163.367
R240 B.n148 B.n147 163.367
R241 B.n147 B.n116 163.367
R242 B.n143 B.n116 163.367
R243 B.n143 B.n142 163.367
R244 B.n142 B.n141 163.367
R245 B.n141 B.n118 163.367
R246 B.n137 B.n118 163.367
R247 B.n137 B.n136 163.367
R248 B.n136 B.n135 163.367
R249 B.n135 B.n120 163.367
R250 B.n131 B.n120 163.367
R251 B.n131 B.n130 163.367
R252 B.n130 B.n129 163.367
R253 B.n129 B.n122 163.367
R254 B.n125 B.n122 163.367
R255 B.n125 B.n124 163.367
R256 B.n124 B.n2 163.367
R257 B.n462 B.n2 163.367
R258 B.n462 B.n461 163.367
R259 B.n461 B.n460 163.367
R260 B.n460 B.n3 163.367
R261 B.n456 B.n3 163.367
R262 B.n456 B.n455 163.367
R263 B.n455 B.n454 163.367
R264 B.n454 B.n5 163.367
R265 B.n450 B.n5 163.367
R266 B.n450 B.n449 163.367
R267 B.n449 B.n448 163.367
R268 B.n448 B.n7 163.367
R269 B.n444 B.n7 163.367
R270 B.n444 B.n443 163.367
R271 B.n443 B.n442 163.367
R272 B.n442 B.n9 163.367
R273 B.n438 B.n9 163.367
R274 B.n438 B.n437 163.367
R275 B.n437 B.n436 163.367
R276 B.n436 B.n11 163.367
R277 B.n432 B.n11 163.367
R278 B.n432 B.n431 163.367
R279 B.n431 B.n430 163.367
R280 B.n430 B.n13 163.367
R281 B.n426 B.n13 163.367
R282 B.n160 B.n159 163.367
R283 B.n161 B.n160 163.367
R284 B.n161 B.n110 163.367
R285 B.n165 B.n110 163.367
R286 B.n166 B.n165 163.367
R287 B.n167 B.n166 163.367
R288 B.n167 B.n108 163.367
R289 B.n171 B.n108 163.367
R290 B.n172 B.n171 163.367
R291 B.n173 B.n172 163.367
R292 B.n173 B.n106 163.367
R293 B.n177 B.n106 163.367
R294 B.n178 B.n177 163.367
R295 B.n179 B.n178 163.367
R296 B.n179 B.n104 163.367
R297 B.n183 B.n104 163.367
R298 B.n184 B.n183 163.367
R299 B.n185 B.n184 163.367
R300 B.n185 B.n102 163.367
R301 B.n189 B.n102 163.367
R302 B.n190 B.n189 163.367
R303 B.n191 B.n190 163.367
R304 B.n191 B.n100 163.367
R305 B.n195 B.n100 163.367
R306 B.n196 B.n195 163.367
R307 B.n197 B.n196 163.367
R308 B.n197 B.n96 163.367
R309 B.n202 B.n96 163.367
R310 B.n203 B.n202 163.367
R311 B.n204 B.n203 163.367
R312 B.n204 B.n94 163.367
R313 B.n208 B.n94 163.367
R314 B.n209 B.n208 163.367
R315 B.n210 B.n209 163.367
R316 B.n210 B.n92 163.367
R317 B.n214 B.n92 163.367
R318 B.n215 B.n214 163.367
R319 B.n215 B.n88 163.367
R320 B.n219 B.n88 163.367
R321 B.n220 B.n219 163.367
R322 B.n221 B.n220 163.367
R323 B.n221 B.n86 163.367
R324 B.n225 B.n86 163.367
R325 B.n226 B.n225 163.367
R326 B.n227 B.n226 163.367
R327 B.n227 B.n84 163.367
R328 B.n231 B.n84 163.367
R329 B.n232 B.n231 163.367
R330 B.n233 B.n232 163.367
R331 B.n233 B.n82 163.367
R332 B.n237 B.n82 163.367
R333 B.n238 B.n237 163.367
R334 B.n239 B.n238 163.367
R335 B.n239 B.n80 163.367
R336 B.n243 B.n80 163.367
R337 B.n244 B.n243 163.367
R338 B.n245 B.n244 163.367
R339 B.n245 B.n78 163.367
R340 B.n249 B.n78 163.367
R341 B.n250 B.n249 163.367
R342 B.n251 B.n250 163.367
R343 B.n251 B.n76 163.367
R344 B.n255 B.n76 163.367
R345 B.n257 B.n256 163.367
R346 B.n257 B.n74 163.367
R347 B.n261 B.n74 163.367
R348 B.n262 B.n261 163.367
R349 B.n263 B.n262 163.367
R350 B.n263 B.n72 163.367
R351 B.n267 B.n72 163.367
R352 B.n268 B.n267 163.367
R353 B.n269 B.n268 163.367
R354 B.n269 B.n70 163.367
R355 B.n273 B.n70 163.367
R356 B.n274 B.n273 163.367
R357 B.n275 B.n274 163.367
R358 B.n275 B.n68 163.367
R359 B.n279 B.n68 163.367
R360 B.n280 B.n279 163.367
R361 B.n281 B.n280 163.367
R362 B.n281 B.n66 163.367
R363 B.n285 B.n66 163.367
R364 B.n286 B.n285 163.367
R365 B.n287 B.n286 163.367
R366 B.n287 B.n64 163.367
R367 B.n291 B.n64 163.367
R368 B.n292 B.n291 163.367
R369 B.n293 B.n292 163.367
R370 B.n293 B.n62 163.367
R371 B.n297 B.n62 163.367
R372 B.n298 B.n297 163.367
R373 B.n299 B.n298 163.367
R374 B.n299 B.n60 163.367
R375 B.n303 B.n60 163.367
R376 B.n304 B.n303 163.367
R377 B.n305 B.n304 163.367
R378 B.n305 B.n58 163.367
R379 B.n309 B.n58 163.367
R380 B.n310 B.n309 163.367
R381 B.n311 B.n310 163.367
R382 B.n311 B.n56 163.367
R383 B.n315 B.n56 163.367
R384 B.n316 B.n315 163.367
R385 B.n317 B.n316 163.367
R386 B.n317 B.n54 163.367
R387 B.n321 B.n54 163.367
R388 B.n322 B.n321 163.367
R389 B.n323 B.n322 163.367
R390 B.n323 B.n52 163.367
R391 B.n327 B.n52 163.367
R392 B.n328 B.n327 163.367
R393 B.n425 B.n424 163.367
R394 B.n424 B.n15 163.367
R395 B.n420 B.n15 163.367
R396 B.n420 B.n419 163.367
R397 B.n419 B.n418 163.367
R398 B.n418 B.n17 163.367
R399 B.n414 B.n17 163.367
R400 B.n414 B.n413 163.367
R401 B.n413 B.n412 163.367
R402 B.n412 B.n19 163.367
R403 B.n408 B.n19 163.367
R404 B.n408 B.n407 163.367
R405 B.n407 B.n406 163.367
R406 B.n406 B.n21 163.367
R407 B.n402 B.n21 163.367
R408 B.n402 B.n401 163.367
R409 B.n401 B.n400 163.367
R410 B.n400 B.n23 163.367
R411 B.n396 B.n23 163.367
R412 B.n396 B.n395 163.367
R413 B.n395 B.n394 163.367
R414 B.n394 B.n25 163.367
R415 B.n390 B.n25 163.367
R416 B.n390 B.n389 163.367
R417 B.n389 B.n388 163.367
R418 B.n388 B.n27 163.367
R419 B.n383 B.n27 163.367
R420 B.n383 B.n382 163.367
R421 B.n382 B.n381 163.367
R422 B.n381 B.n31 163.367
R423 B.n377 B.n31 163.367
R424 B.n377 B.n376 163.367
R425 B.n376 B.n375 163.367
R426 B.n375 B.n33 163.367
R427 B.n371 B.n33 163.367
R428 B.n371 B.n370 163.367
R429 B.n370 B.n369 163.367
R430 B.n369 B.n35 163.367
R431 B.n365 B.n35 163.367
R432 B.n365 B.n364 163.367
R433 B.n364 B.n363 163.367
R434 B.n363 B.n40 163.367
R435 B.n359 B.n40 163.367
R436 B.n359 B.n358 163.367
R437 B.n358 B.n357 163.367
R438 B.n357 B.n42 163.367
R439 B.n353 B.n42 163.367
R440 B.n353 B.n352 163.367
R441 B.n352 B.n351 163.367
R442 B.n351 B.n44 163.367
R443 B.n347 B.n44 163.367
R444 B.n347 B.n346 163.367
R445 B.n346 B.n345 163.367
R446 B.n345 B.n46 163.367
R447 B.n341 B.n46 163.367
R448 B.n341 B.n340 163.367
R449 B.n340 B.n339 163.367
R450 B.n339 B.n48 163.367
R451 B.n335 B.n48 163.367
R452 B.n335 B.n334 163.367
R453 B.n334 B.n333 163.367
R454 B.n333 B.n50 163.367
R455 B.n329 B.n50 163.367
R456 B.n89 B.t11 133.381
R457 B.n36 B.t4 133.381
R458 B.n97 B.t2 133.374
R459 B.n28 B.t7 133.374
R460 B.n90 B.t10 116.12
R461 B.n37 B.t5 116.12
R462 B.n98 B.t1 116.112
R463 B.n29 B.t8 116.112
R464 B.n91 B.n90 59.5399
R465 B.n199 B.n98 59.5399
R466 B.n385 B.n29 59.5399
R467 B.n38 B.n37 59.5399
R468 B.n427 B.n14 31.6883
R469 B.n330 B.n51 31.6883
R470 B.n254 B.n75 31.6883
R471 B.n158 B.n157 31.6883
R472 B B.n463 18.0485
R473 B.n90 B.n89 17.2611
R474 B.n98 B.n97 17.2611
R475 B.n29 B.n28 17.2611
R476 B.n37 B.n36 17.2611
R477 B.n423 B.n14 10.6151
R478 B.n423 B.n422 10.6151
R479 B.n422 B.n421 10.6151
R480 B.n421 B.n16 10.6151
R481 B.n417 B.n16 10.6151
R482 B.n417 B.n416 10.6151
R483 B.n416 B.n415 10.6151
R484 B.n415 B.n18 10.6151
R485 B.n411 B.n18 10.6151
R486 B.n411 B.n410 10.6151
R487 B.n410 B.n409 10.6151
R488 B.n409 B.n20 10.6151
R489 B.n405 B.n20 10.6151
R490 B.n405 B.n404 10.6151
R491 B.n404 B.n403 10.6151
R492 B.n403 B.n22 10.6151
R493 B.n399 B.n22 10.6151
R494 B.n399 B.n398 10.6151
R495 B.n398 B.n397 10.6151
R496 B.n397 B.n24 10.6151
R497 B.n393 B.n24 10.6151
R498 B.n393 B.n392 10.6151
R499 B.n392 B.n391 10.6151
R500 B.n391 B.n26 10.6151
R501 B.n387 B.n26 10.6151
R502 B.n387 B.n386 10.6151
R503 B.n384 B.n30 10.6151
R504 B.n380 B.n30 10.6151
R505 B.n380 B.n379 10.6151
R506 B.n379 B.n378 10.6151
R507 B.n378 B.n32 10.6151
R508 B.n374 B.n32 10.6151
R509 B.n374 B.n373 10.6151
R510 B.n373 B.n372 10.6151
R511 B.n372 B.n34 10.6151
R512 B.n368 B.n367 10.6151
R513 B.n367 B.n366 10.6151
R514 B.n366 B.n39 10.6151
R515 B.n362 B.n39 10.6151
R516 B.n362 B.n361 10.6151
R517 B.n361 B.n360 10.6151
R518 B.n360 B.n41 10.6151
R519 B.n356 B.n41 10.6151
R520 B.n356 B.n355 10.6151
R521 B.n355 B.n354 10.6151
R522 B.n354 B.n43 10.6151
R523 B.n350 B.n43 10.6151
R524 B.n350 B.n349 10.6151
R525 B.n349 B.n348 10.6151
R526 B.n348 B.n45 10.6151
R527 B.n344 B.n45 10.6151
R528 B.n344 B.n343 10.6151
R529 B.n343 B.n342 10.6151
R530 B.n342 B.n47 10.6151
R531 B.n338 B.n47 10.6151
R532 B.n338 B.n337 10.6151
R533 B.n337 B.n336 10.6151
R534 B.n336 B.n49 10.6151
R535 B.n332 B.n49 10.6151
R536 B.n332 B.n331 10.6151
R537 B.n331 B.n330 10.6151
R538 B.n258 B.n75 10.6151
R539 B.n259 B.n258 10.6151
R540 B.n260 B.n259 10.6151
R541 B.n260 B.n73 10.6151
R542 B.n264 B.n73 10.6151
R543 B.n265 B.n264 10.6151
R544 B.n266 B.n265 10.6151
R545 B.n266 B.n71 10.6151
R546 B.n270 B.n71 10.6151
R547 B.n271 B.n270 10.6151
R548 B.n272 B.n271 10.6151
R549 B.n272 B.n69 10.6151
R550 B.n276 B.n69 10.6151
R551 B.n277 B.n276 10.6151
R552 B.n278 B.n277 10.6151
R553 B.n278 B.n67 10.6151
R554 B.n282 B.n67 10.6151
R555 B.n283 B.n282 10.6151
R556 B.n284 B.n283 10.6151
R557 B.n284 B.n65 10.6151
R558 B.n288 B.n65 10.6151
R559 B.n289 B.n288 10.6151
R560 B.n290 B.n289 10.6151
R561 B.n290 B.n63 10.6151
R562 B.n294 B.n63 10.6151
R563 B.n295 B.n294 10.6151
R564 B.n296 B.n295 10.6151
R565 B.n296 B.n61 10.6151
R566 B.n300 B.n61 10.6151
R567 B.n301 B.n300 10.6151
R568 B.n302 B.n301 10.6151
R569 B.n302 B.n59 10.6151
R570 B.n306 B.n59 10.6151
R571 B.n307 B.n306 10.6151
R572 B.n308 B.n307 10.6151
R573 B.n308 B.n57 10.6151
R574 B.n312 B.n57 10.6151
R575 B.n313 B.n312 10.6151
R576 B.n314 B.n313 10.6151
R577 B.n314 B.n55 10.6151
R578 B.n318 B.n55 10.6151
R579 B.n319 B.n318 10.6151
R580 B.n320 B.n319 10.6151
R581 B.n320 B.n53 10.6151
R582 B.n324 B.n53 10.6151
R583 B.n325 B.n324 10.6151
R584 B.n326 B.n325 10.6151
R585 B.n326 B.n51 10.6151
R586 B.n158 B.n111 10.6151
R587 B.n162 B.n111 10.6151
R588 B.n163 B.n162 10.6151
R589 B.n164 B.n163 10.6151
R590 B.n164 B.n109 10.6151
R591 B.n168 B.n109 10.6151
R592 B.n169 B.n168 10.6151
R593 B.n170 B.n169 10.6151
R594 B.n170 B.n107 10.6151
R595 B.n174 B.n107 10.6151
R596 B.n175 B.n174 10.6151
R597 B.n176 B.n175 10.6151
R598 B.n176 B.n105 10.6151
R599 B.n180 B.n105 10.6151
R600 B.n181 B.n180 10.6151
R601 B.n182 B.n181 10.6151
R602 B.n182 B.n103 10.6151
R603 B.n186 B.n103 10.6151
R604 B.n187 B.n186 10.6151
R605 B.n188 B.n187 10.6151
R606 B.n188 B.n101 10.6151
R607 B.n192 B.n101 10.6151
R608 B.n193 B.n192 10.6151
R609 B.n194 B.n193 10.6151
R610 B.n194 B.n99 10.6151
R611 B.n198 B.n99 10.6151
R612 B.n201 B.n200 10.6151
R613 B.n201 B.n95 10.6151
R614 B.n205 B.n95 10.6151
R615 B.n206 B.n205 10.6151
R616 B.n207 B.n206 10.6151
R617 B.n207 B.n93 10.6151
R618 B.n211 B.n93 10.6151
R619 B.n212 B.n211 10.6151
R620 B.n213 B.n212 10.6151
R621 B.n217 B.n216 10.6151
R622 B.n218 B.n217 10.6151
R623 B.n218 B.n87 10.6151
R624 B.n222 B.n87 10.6151
R625 B.n223 B.n222 10.6151
R626 B.n224 B.n223 10.6151
R627 B.n224 B.n85 10.6151
R628 B.n228 B.n85 10.6151
R629 B.n229 B.n228 10.6151
R630 B.n230 B.n229 10.6151
R631 B.n230 B.n83 10.6151
R632 B.n234 B.n83 10.6151
R633 B.n235 B.n234 10.6151
R634 B.n236 B.n235 10.6151
R635 B.n236 B.n81 10.6151
R636 B.n240 B.n81 10.6151
R637 B.n241 B.n240 10.6151
R638 B.n242 B.n241 10.6151
R639 B.n242 B.n79 10.6151
R640 B.n246 B.n79 10.6151
R641 B.n247 B.n246 10.6151
R642 B.n248 B.n247 10.6151
R643 B.n248 B.n77 10.6151
R644 B.n252 B.n77 10.6151
R645 B.n253 B.n252 10.6151
R646 B.n254 B.n253 10.6151
R647 B.n157 B.n156 10.6151
R648 B.n156 B.n113 10.6151
R649 B.n152 B.n113 10.6151
R650 B.n152 B.n151 10.6151
R651 B.n151 B.n150 10.6151
R652 B.n150 B.n115 10.6151
R653 B.n146 B.n115 10.6151
R654 B.n146 B.n145 10.6151
R655 B.n145 B.n144 10.6151
R656 B.n144 B.n117 10.6151
R657 B.n140 B.n117 10.6151
R658 B.n140 B.n139 10.6151
R659 B.n139 B.n138 10.6151
R660 B.n138 B.n119 10.6151
R661 B.n134 B.n119 10.6151
R662 B.n134 B.n133 10.6151
R663 B.n133 B.n132 10.6151
R664 B.n132 B.n121 10.6151
R665 B.n128 B.n121 10.6151
R666 B.n128 B.n127 10.6151
R667 B.n127 B.n126 10.6151
R668 B.n126 B.n123 10.6151
R669 B.n123 B.n0 10.6151
R670 B.n459 B.n1 10.6151
R671 B.n459 B.n458 10.6151
R672 B.n458 B.n457 10.6151
R673 B.n457 B.n4 10.6151
R674 B.n453 B.n4 10.6151
R675 B.n453 B.n452 10.6151
R676 B.n452 B.n451 10.6151
R677 B.n451 B.n6 10.6151
R678 B.n447 B.n6 10.6151
R679 B.n447 B.n446 10.6151
R680 B.n446 B.n445 10.6151
R681 B.n445 B.n8 10.6151
R682 B.n441 B.n8 10.6151
R683 B.n441 B.n440 10.6151
R684 B.n440 B.n439 10.6151
R685 B.n439 B.n10 10.6151
R686 B.n435 B.n10 10.6151
R687 B.n435 B.n434 10.6151
R688 B.n434 B.n433 10.6151
R689 B.n433 B.n12 10.6151
R690 B.n429 B.n12 10.6151
R691 B.n429 B.n428 10.6151
R692 B.n428 B.n427 10.6151
R693 B.n386 B.n385 9.36635
R694 B.n368 B.n38 9.36635
R695 B.n199 B.n198 9.36635
R696 B.n216 B.n91 9.36635
R697 B.n463 B.n0 2.81026
R698 B.n463 B.n1 2.81026
R699 B.n385 B.n384 1.24928
R700 B.n38 B.n34 1.24928
R701 B.n200 B.n199 1.24928
R702 B.n213 B.n91 1.24928
R703 VP.n6 VP.t0 401.625
R704 VP.n14 VP.t3 377.423
R705 VP.n16 VP.t4 377.423
R706 VP.n1 VP.t6 377.423
R707 VP.n20 VP.t8 377.423
R708 VP.n22 VP.t9 377.423
R709 VP.n11 VP.t1 377.423
R710 VP.n9 VP.t5 377.423
R711 VP.n8 VP.t2 377.423
R712 VP.n7 VP.t7 377.423
R713 VP.n23 VP.n22 161.3
R714 VP.n9 VP.n4 161.3
R715 VP.n10 VP.n3 161.3
R716 VP.n12 VP.n11 161.3
R717 VP.n21 VP.n0 161.3
R718 VP.n20 VP.n19 161.3
R719 VP.n17 VP.n16 161.3
R720 VP.n15 VP.n2 161.3
R721 VP.n14 VP.n13 161.3
R722 VP.n8 VP.n5 80.6037
R723 VP.n18 VP.n1 80.6037
R724 VP.n16 VP.n1 48.2005
R725 VP.n20 VP.n1 48.2005
R726 VP.n9 VP.n8 48.2005
R727 VP.n8 VP.n7 48.2005
R728 VP.n6 VP.n5 45.0238
R729 VP.n13 VP.n12 38.2846
R730 VP.n15 VP.n14 36.5157
R731 VP.n22 VP.n21 36.5157
R732 VP.n11 VP.n10 36.5157
R733 VP.n7 VP.n6 17.2829
R734 VP.n16 VP.n15 11.6853
R735 VP.n21 VP.n20 11.6853
R736 VP.n10 VP.n9 11.6853
R737 VP.n5 VP.n4 0.285035
R738 VP.n18 VP.n17 0.285035
R739 VP.n19 VP.n18 0.285035
R740 VP.n4 VP.n3 0.189894
R741 VP.n12 VP.n3 0.189894
R742 VP.n13 VP.n2 0.189894
R743 VP.n17 VP.n2 0.189894
R744 VP.n19 VP.n0 0.189894
R745 VP.n23 VP.n0 0.189894
R746 VP VP.n23 0.0516364
R747 VTAIL.n11 VTAIL.t9 75.8035
R748 VTAIL.n16 VTAIL.t15 75.8033
R749 VTAIL.n17 VTAIL.t1 75.8033
R750 VTAIL.n2 VTAIL.t16 75.8033
R751 VTAIL.n15 VTAIL.n14 71.251
R752 VTAIL.n13 VTAIL.n12 71.251
R753 VTAIL.n10 VTAIL.n9 71.251
R754 VTAIL.n8 VTAIL.n7 71.251
R755 VTAIL.n19 VTAIL.n18 71.2509
R756 VTAIL.n1 VTAIL.n0 71.2509
R757 VTAIL.n4 VTAIL.n3 71.2509
R758 VTAIL.n6 VTAIL.n5 71.2509
R759 VTAIL.n8 VTAIL.n6 20.0565
R760 VTAIL.n17 VTAIL.n16 19.2893
R761 VTAIL.n18 VTAIL.t8 4.55302
R762 VTAIL.n18 VTAIL.t5 4.55302
R763 VTAIL.n0 VTAIL.t3 4.55302
R764 VTAIL.n0 VTAIL.t4 4.55302
R765 VTAIL.n3 VTAIL.t12 4.55302
R766 VTAIL.n3 VTAIL.t13 4.55302
R767 VTAIL.n5 VTAIL.t17 4.55302
R768 VTAIL.n5 VTAIL.t11 4.55302
R769 VTAIL.n14 VTAIL.t19 4.55302
R770 VTAIL.n14 VTAIL.t18 4.55302
R771 VTAIL.n12 VTAIL.t10 4.55302
R772 VTAIL.n12 VTAIL.t14 4.55302
R773 VTAIL.n9 VTAIL.t0 4.55302
R774 VTAIL.n9 VTAIL.t7 4.55302
R775 VTAIL.n7 VTAIL.t2 4.55302
R776 VTAIL.n7 VTAIL.t6 4.55302
R777 VTAIL.n13 VTAIL.n11 0.853948
R778 VTAIL.n2 VTAIL.n1 0.853948
R779 VTAIL.n10 VTAIL.n8 0.767741
R780 VTAIL.n11 VTAIL.n10 0.767741
R781 VTAIL.n15 VTAIL.n13 0.767741
R782 VTAIL.n16 VTAIL.n15 0.767741
R783 VTAIL.n6 VTAIL.n4 0.767741
R784 VTAIL.n4 VTAIL.n2 0.767741
R785 VTAIL.n19 VTAIL.n17 0.767741
R786 VTAIL VTAIL.n1 0.634121
R787 VTAIL VTAIL.n19 0.134121
R788 VDD1.n1 VDD1.t9 93.2495
R789 VDD1.n3 VDD1.t6 93.2493
R790 VDD1.n5 VDD1.n4 88.4498
R791 VDD1.n1 VDD1.n0 87.9298
R792 VDD1.n3 VDD1.n2 87.9297
R793 VDD1.n7 VDD1.n6 87.9296
R794 VDD1.n7 VDD1.n5 34.4815
R795 VDD1.n6 VDD1.t4 4.55302
R796 VDD1.n6 VDD1.t8 4.55302
R797 VDD1.n0 VDD1.t2 4.55302
R798 VDD1.n0 VDD1.t7 4.55302
R799 VDD1.n4 VDD1.t1 4.55302
R800 VDD1.n4 VDD1.t0 4.55302
R801 VDD1.n2 VDD1.t5 4.55302
R802 VDD1.n2 VDD1.t3 4.55302
R803 VDD1 VDD1.n7 0.517741
R804 VDD1 VDD1.n1 0.2505
R805 VDD1.n5 VDD1.n3 0.136964
R806 VN.n3 VN.t1 401.625
R807 VN.n13 VN.t4 401.625
R808 VN.n2 VN.t0 377.423
R809 VN.n1 VN.t2 377.423
R810 VN.n6 VN.t7 377.423
R811 VN.n8 VN.t6 377.423
R812 VN.n12 VN.t9 377.423
R813 VN.n11 VN.t3 377.423
R814 VN.n16 VN.t8 377.423
R815 VN.n18 VN.t5 377.423
R816 VN.n9 VN.n8 161.3
R817 VN.n19 VN.n18 161.3
R818 VN.n17 VN.n10 161.3
R819 VN.n16 VN.n15 161.3
R820 VN.n7 VN.n0 161.3
R821 VN.n6 VN.n5 161.3
R822 VN.n14 VN.n11 80.6037
R823 VN.n4 VN.n1 80.6037
R824 VN.n2 VN.n1 48.2005
R825 VN.n6 VN.n1 48.2005
R826 VN.n12 VN.n11 48.2005
R827 VN.n16 VN.n11 48.2005
R828 VN.n14 VN.n13 45.0238
R829 VN.n4 VN.n3 45.0238
R830 VN VN.n19 38.6653
R831 VN.n8 VN.n7 36.5157
R832 VN.n18 VN.n17 36.5157
R833 VN.n3 VN.n2 17.2829
R834 VN.n13 VN.n12 17.2829
R835 VN.n7 VN.n6 11.6853
R836 VN.n17 VN.n16 11.6853
R837 VN.n15 VN.n14 0.285035
R838 VN.n5 VN.n4 0.285035
R839 VN.n19 VN.n10 0.189894
R840 VN.n15 VN.n10 0.189894
R841 VN.n5 VN.n0 0.189894
R842 VN.n9 VN.n0 0.189894
R843 VN VN.n9 0.0516364
R844 VDD2.n1 VDD2.t8 93.2493
R845 VDD2.n4 VDD2.t4 92.4823
R846 VDD2.n3 VDD2.n2 88.4498
R847 VDD2 VDD2.n7 88.4468
R848 VDD2.n6 VDD2.n5 87.9298
R849 VDD2.n1 VDD2.n0 87.9297
R850 VDD2.n4 VDD2.n3 33.5149
R851 VDD2.n7 VDD2.t0 4.55302
R852 VDD2.n7 VDD2.t5 4.55302
R853 VDD2.n5 VDD2.t1 4.55302
R854 VDD2.n5 VDD2.t6 4.55302
R855 VDD2.n2 VDD2.t2 4.55302
R856 VDD2.n2 VDD2.t3 4.55302
R857 VDD2.n0 VDD2.t9 4.55302
R858 VDD2.n0 VDD2.t7 4.55302
R859 VDD2.n6 VDD2.n4 0.767741
R860 VDD2 VDD2.n6 0.2505
R861 VDD2.n3 VDD2.n1 0.136964
C0 B VTAIL 1.79385f
C1 VTAIL VN 3.69406f
C2 w_n2038_n2396# VDD1 1.61736f
C3 VP B 1.13137f
C4 w_n2038_n2396# VTAIL 2.26548f
C5 VP VN 4.49161f
C6 VP w_n2038_n2396# 3.91053f
C7 VTAIL VDD1 10.3009f
C8 B VDD2 1.33111f
C9 VDD2 VN 3.68213f
C10 VP VDD1 3.85335f
C11 VP VTAIL 3.70849f
C12 w_n2038_n2396# VDD2 1.65487f
C13 B VN 0.707032f
C14 w_n2038_n2396# B 5.75817f
C15 VDD2 VDD1 0.883714f
C16 w_n2038_n2396# VN 3.65149f
C17 VDD2 VTAIL 10.3365f
C18 VP VDD2 0.323314f
C19 B VDD1 1.29219f
C20 VDD1 VN 0.149005f
C21 VDD2 VSUBS 1.188597f
C22 VDD1 VSUBS 0.952821f
C23 VTAIL VSUBS 0.44689f
C24 VN VSUBS 4.37862f
C25 VP VSUBS 1.389303f
C26 B VSUBS 2.42447f
C27 w_n2038_n2396# VSUBS 60.724197f
C28 VDD2.t8 VSUBS 1.33328f
C29 VDD2.t9 VSUBS 0.143606f
C30 VDD2.t7 VSUBS 0.143606f
C31 VDD2.n0 VSUBS 0.998314f
C32 VDD2.n1 VSUBS 1.07406f
C33 VDD2.t2 VSUBS 0.143606f
C34 VDD2.t3 VSUBS 0.143606f
C35 VDD2.n2 VSUBS 1.00155f
C36 VDD2.n3 VSUBS 1.7887f
C37 VDD2.t4 VSUBS 1.32862f
C38 VDD2.n4 VSUBS 2.20229f
C39 VDD2.t1 VSUBS 0.143606f
C40 VDD2.t6 VSUBS 0.143606f
C41 VDD2.n5 VSUBS 0.998317f
C42 VDD2.n6 VSUBS 0.516305f
C43 VDD2.t0 VSUBS 0.143606f
C44 VDD2.t5 VSUBS 0.143606f
C45 VDD2.n7 VSUBS 1.00152f
C46 VN.n0 VSUBS 0.061133f
C47 VN.t2 VSUBS 0.705171f
C48 VN.n1 VSUBS 0.329322f
C49 VN.t1 VSUBS 0.72412f
C50 VN.t0 VSUBS 0.705171f
C51 VN.n2 VSUBS 0.326564f
C52 VN.n3 VSUBS 0.300979f
C53 VN.n4 VSUBS 0.288027f
C54 VN.n5 VSUBS 0.081575f
C55 VN.t7 VSUBS 0.705171f
C56 VN.n6 VSUBS 0.318464f
C57 VN.n7 VSUBS 0.013872f
C58 VN.t6 VSUBS 0.705171f
C59 VN.n8 VSUBS 0.312434f
C60 VN.n9 VSUBS 0.047376f
C61 VN.n10 VSUBS 0.061133f
C62 VN.t3 VSUBS 0.705171f
C63 VN.n11 VSUBS 0.329322f
C64 VN.t8 VSUBS 0.705171f
C65 VN.t4 VSUBS 0.72412f
C66 VN.t9 VSUBS 0.705171f
C67 VN.n12 VSUBS 0.326564f
C68 VN.n13 VSUBS 0.300979f
C69 VN.n14 VSUBS 0.288027f
C70 VN.n15 VSUBS 0.081575f
C71 VN.n16 VSUBS 0.318464f
C72 VN.n17 VSUBS 0.013872f
C73 VN.t5 VSUBS 0.705171f
C74 VN.n18 VSUBS 0.312434f
C75 VN.n19 VSUBS 2.19145f
C76 VDD1.t9 VSUBS 1.34331f
C77 VDD1.t2 VSUBS 0.144686f
C78 VDD1.t7 VSUBS 0.144686f
C79 VDD1.n0 VSUBS 1.00583f
C80 VDD1.n1 VSUBS 1.08716f
C81 VDD1.t6 VSUBS 1.34331f
C82 VDD1.t5 VSUBS 0.144686f
C83 VDD1.t3 VSUBS 0.144686f
C84 VDD1.n2 VSUBS 1.00582f
C85 VDD1.n3 VSUBS 1.08214f
C86 VDD1.t1 VSUBS 0.144686f
C87 VDD1.t0 VSUBS 0.144686f
C88 VDD1.n4 VSUBS 1.00908f
C89 VDD1.n5 VSUBS 1.87611f
C90 VDD1.t4 VSUBS 0.144686f
C91 VDD1.t8 VSUBS 0.144686f
C92 VDD1.n6 VSUBS 1.00582f
C93 VDD1.n7 VSUBS 2.22054f
C94 VTAIL.t3 VSUBS 0.169376f
C95 VTAIL.t4 VSUBS 0.169376f
C96 VTAIL.n0 VSUBS 1.05928f
C97 VTAIL.n1 VSUBS 0.731782f
C98 VTAIL.t16 VSUBS 1.44003f
C99 VTAIL.n2 VSUBS 0.825897f
C100 VTAIL.t12 VSUBS 0.169376f
C101 VTAIL.t13 VSUBS 0.169376f
C102 VTAIL.n3 VSUBS 1.05928f
C103 VTAIL.n4 VSUBS 0.736369f
C104 VTAIL.t17 VSUBS 0.169376f
C105 VTAIL.t11 VSUBS 0.169376f
C106 VTAIL.n5 VSUBS 1.05928f
C107 VTAIL.n6 VSUBS 1.81374f
C108 VTAIL.t2 VSUBS 0.169376f
C109 VTAIL.t6 VSUBS 0.169376f
C110 VTAIL.n7 VSUBS 1.05929f
C111 VTAIL.n8 VSUBS 1.81374f
C112 VTAIL.t0 VSUBS 0.169376f
C113 VTAIL.t7 VSUBS 0.169376f
C114 VTAIL.n9 VSUBS 1.05929f
C115 VTAIL.n10 VSUBS 0.736364f
C116 VTAIL.t9 VSUBS 1.44003f
C117 VTAIL.n11 VSUBS 0.825891f
C118 VTAIL.t10 VSUBS 0.169376f
C119 VTAIL.t14 VSUBS 0.169376f
C120 VTAIL.n12 VSUBS 1.05929f
C121 VTAIL.n13 VSUBS 0.744703f
C122 VTAIL.t19 VSUBS 0.169376f
C123 VTAIL.t18 VSUBS 0.169376f
C124 VTAIL.n14 VSUBS 1.05929f
C125 VTAIL.n15 VSUBS 0.736364f
C126 VTAIL.t15 VSUBS 1.44003f
C127 VTAIL.n16 VSUBS 1.82072f
C128 VTAIL.t1 VSUBS 1.44003f
C129 VTAIL.n17 VSUBS 1.82072f
C130 VTAIL.t8 VSUBS 0.169376f
C131 VTAIL.t5 VSUBS 0.169376f
C132 VTAIL.n18 VSUBS 1.05928f
C133 VTAIL.n19 VSUBS 0.675079f
C134 VP.n0 VSUBS 0.063048f
C135 VP.t6 VSUBS 0.727259f
C136 VP.n1 VSUBS 0.339637f
C137 VP.n2 VSUBS 0.063048f
C138 VP.n3 VSUBS 0.063048f
C139 VP.t1 VSUBS 0.727259f
C140 VP.t5 VSUBS 0.727259f
C141 VP.n4 VSUBS 0.08413f
C142 VP.t2 VSUBS 0.727259f
C143 VP.n5 VSUBS 0.297049f
C144 VP.t7 VSUBS 0.727259f
C145 VP.t0 VSUBS 0.746802f
C146 VP.n6 VSUBS 0.310407f
C147 VP.n7 VSUBS 0.336792f
C148 VP.n8 VSUBS 0.339637f
C149 VP.n9 VSUBS 0.328439f
C150 VP.n10 VSUBS 0.014307f
C151 VP.n11 VSUBS 0.32222f
C152 VP.n12 VSUBS 2.21845f
C153 VP.n13 VSUBS 2.27782f
C154 VP.t3 VSUBS 0.727259f
C155 VP.n14 VSUBS 0.32222f
C156 VP.n15 VSUBS 0.014307f
C157 VP.t4 VSUBS 0.727259f
C158 VP.n16 VSUBS 0.328439f
C159 VP.n17 VSUBS 0.08413f
C160 VP.n18 VSUBS 0.083933f
C161 VP.n19 VSUBS 0.08413f
C162 VP.t8 VSUBS 0.727259f
C163 VP.n20 VSUBS 0.328439f
C164 VP.n21 VSUBS 0.014307f
C165 VP.t9 VSUBS 0.727259f
C166 VP.n22 VSUBS 0.32222f
C167 VP.n23 VSUBS 0.04886f
C168 B.n0 VSUBS 0.004001f
C169 B.n1 VSUBS 0.004001f
C170 B.n2 VSUBS 0.006327f
C171 B.n3 VSUBS 0.006327f
C172 B.n4 VSUBS 0.006327f
C173 B.n5 VSUBS 0.006327f
C174 B.n6 VSUBS 0.006327f
C175 B.n7 VSUBS 0.006327f
C176 B.n8 VSUBS 0.006327f
C177 B.n9 VSUBS 0.006327f
C178 B.n10 VSUBS 0.006327f
C179 B.n11 VSUBS 0.006327f
C180 B.n12 VSUBS 0.006327f
C181 B.n13 VSUBS 0.006327f
C182 B.n14 VSUBS 0.014694f
C183 B.n15 VSUBS 0.006327f
C184 B.n16 VSUBS 0.006327f
C185 B.n17 VSUBS 0.006327f
C186 B.n18 VSUBS 0.006327f
C187 B.n19 VSUBS 0.006327f
C188 B.n20 VSUBS 0.006327f
C189 B.n21 VSUBS 0.006327f
C190 B.n22 VSUBS 0.006327f
C191 B.n23 VSUBS 0.006327f
C192 B.n24 VSUBS 0.006327f
C193 B.n25 VSUBS 0.006327f
C194 B.n26 VSUBS 0.006327f
C195 B.n27 VSUBS 0.006327f
C196 B.t8 VSUBS 0.195042f
C197 B.t7 VSUBS 0.201235f
C198 B.t6 VSUBS 0.15186f
C199 B.n28 VSUBS 0.082895f
C200 B.n29 VSUBS 0.056877f
C201 B.n30 VSUBS 0.006327f
C202 B.n31 VSUBS 0.006327f
C203 B.n32 VSUBS 0.006327f
C204 B.n33 VSUBS 0.006327f
C205 B.n34 VSUBS 0.003536f
C206 B.n35 VSUBS 0.006327f
C207 B.t5 VSUBS 0.195041f
C208 B.t4 VSUBS 0.201234f
C209 B.t3 VSUBS 0.15186f
C210 B.n36 VSUBS 0.082897f
C211 B.n37 VSUBS 0.056878f
C212 B.n38 VSUBS 0.01466f
C213 B.n39 VSUBS 0.006327f
C214 B.n40 VSUBS 0.006327f
C215 B.n41 VSUBS 0.006327f
C216 B.n42 VSUBS 0.006327f
C217 B.n43 VSUBS 0.006327f
C218 B.n44 VSUBS 0.006327f
C219 B.n45 VSUBS 0.006327f
C220 B.n46 VSUBS 0.006327f
C221 B.n47 VSUBS 0.006327f
C222 B.n48 VSUBS 0.006327f
C223 B.n49 VSUBS 0.006327f
C224 B.n50 VSUBS 0.006327f
C225 B.n51 VSUBS 0.015108f
C226 B.n52 VSUBS 0.006327f
C227 B.n53 VSUBS 0.006327f
C228 B.n54 VSUBS 0.006327f
C229 B.n55 VSUBS 0.006327f
C230 B.n56 VSUBS 0.006327f
C231 B.n57 VSUBS 0.006327f
C232 B.n58 VSUBS 0.006327f
C233 B.n59 VSUBS 0.006327f
C234 B.n60 VSUBS 0.006327f
C235 B.n61 VSUBS 0.006327f
C236 B.n62 VSUBS 0.006327f
C237 B.n63 VSUBS 0.006327f
C238 B.n64 VSUBS 0.006327f
C239 B.n65 VSUBS 0.006327f
C240 B.n66 VSUBS 0.006327f
C241 B.n67 VSUBS 0.006327f
C242 B.n68 VSUBS 0.006327f
C243 B.n69 VSUBS 0.006327f
C244 B.n70 VSUBS 0.006327f
C245 B.n71 VSUBS 0.006327f
C246 B.n72 VSUBS 0.006327f
C247 B.n73 VSUBS 0.006327f
C248 B.n74 VSUBS 0.006327f
C249 B.n75 VSUBS 0.014337f
C250 B.n76 VSUBS 0.006327f
C251 B.n77 VSUBS 0.006327f
C252 B.n78 VSUBS 0.006327f
C253 B.n79 VSUBS 0.006327f
C254 B.n80 VSUBS 0.006327f
C255 B.n81 VSUBS 0.006327f
C256 B.n82 VSUBS 0.006327f
C257 B.n83 VSUBS 0.006327f
C258 B.n84 VSUBS 0.006327f
C259 B.n85 VSUBS 0.006327f
C260 B.n86 VSUBS 0.006327f
C261 B.n87 VSUBS 0.006327f
C262 B.n88 VSUBS 0.006327f
C263 B.t10 VSUBS 0.195041f
C264 B.t11 VSUBS 0.201234f
C265 B.t9 VSUBS 0.15186f
C266 B.n89 VSUBS 0.082897f
C267 B.n90 VSUBS 0.056878f
C268 B.n91 VSUBS 0.01466f
C269 B.n92 VSUBS 0.006327f
C270 B.n93 VSUBS 0.006327f
C271 B.n94 VSUBS 0.006327f
C272 B.n95 VSUBS 0.006327f
C273 B.n96 VSUBS 0.006327f
C274 B.t1 VSUBS 0.195042f
C275 B.t2 VSUBS 0.201235f
C276 B.t0 VSUBS 0.15186f
C277 B.n97 VSUBS 0.082895f
C278 B.n98 VSUBS 0.056877f
C279 B.n99 VSUBS 0.006327f
C280 B.n100 VSUBS 0.006327f
C281 B.n101 VSUBS 0.006327f
C282 B.n102 VSUBS 0.006327f
C283 B.n103 VSUBS 0.006327f
C284 B.n104 VSUBS 0.006327f
C285 B.n105 VSUBS 0.006327f
C286 B.n106 VSUBS 0.006327f
C287 B.n107 VSUBS 0.006327f
C288 B.n108 VSUBS 0.006327f
C289 B.n109 VSUBS 0.006327f
C290 B.n110 VSUBS 0.006327f
C291 B.n111 VSUBS 0.006327f
C292 B.n112 VSUBS 0.014337f
C293 B.n113 VSUBS 0.006327f
C294 B.n114 VSUBS 0.006327f
C295 B.n115 VSUBS 0.006327f
C296 B.n116 VSUBS 0.006327f
C297 B.n117 VSUBS 0.006327f
C298 B.n118 VSUBS 0.006327f
C299 B.n119 VSUBS 0.006327f
C300 B.n120 VSUBS 0.006327f
C301 B.n121 VSUBS 0.006327f
C302 B.n122 VSUBS 0.006327f
C303 B.n123 VSUBS 0.006327f
C304 B.n124 VSUBS 0.006327f
C305 B.n125 VSUBS 0.006327f
C306 B.n126 VSUBS 0.006327f
C307 B.n127 VSUBS 0.006327f
C308 B.n128 VSUBS 0.006327f
C309 B.n129 VSUBS 0.006327f
C310 B.n130 VSUBS 0.006327f
C311 B.n131 VSUBS 0.006327f
C312 B.n132 VSUBS 0.006327f
C313 B.n133 VSUBS 0.006327f
C314 B.n134 VSUBS 0.006327f
C315 B.n135 VSUBS 0.006327f
C316 B.n136 VSUBS 0.006327f
C317 B.n137 VSUBS 0.006327f
C318 B.n138 VSUBS 0.006327f
C319 B.n139 VSUBS 0.006327f
C320 B.n140 VSUBS 0.006327f
C321 B.n141 VSUBS 0.006327f
C322 B.n142 VSUBS 0.006327f
C323 B.n143 VSUBS 0.006327f
C324 B.n144 VSUBS 0.006327f
C325 B.n145 VSUBS 0.006327f
C326 B.n146 VSUBS 0.006327f
C327 B.n147 VSUBS 0.006327f
C328 B.n148 VSUBS 0.006327f
C329 B.n149 VSUBS 0.006327f
C330 B.n150 VSUBS 0.006327f
C331 B.n151 VSUBS 0.006327f
C332 B.n152 VSUBS 0.006327f
C333 B.n153 VSUBS 0.006327f
C334 B.n154 VSUBS 0.006327f
C335 B.n155 VSUBS 0.006327f
C336 B.n156 VSUBS 0.006327f
C337 B.n157 VSUBS 0.014337f
C338 B.n158 VSUBS 0.014694f
C339 B.n159 VSUBS 0.014694f
C340 B.n160 VSUBS 0.006327f
C341 B.n161 VSUBS 0.006327f
C342 B.n162 VSUBS 0.006327f
C343 B.n163 VSUBS 0.006327f
C344 B.n164 VSUBS 0.006327f
C345 B.n165 VSUBS 0.006327f
C346 B.n166 VSUBS 0.006327f
C347 B.n167 VSUBS 0.006327f
C348 B.n168 VSUBS 0.006327f
C349 B.n169 VSUBS 0.006327f
C350 B.n170 VSUBS 0.006327f
C351 B.n171 VSUBS 0.006327f
C352 B.n172 VSUBS 0.006327f
C353 B.n173 VSUBS 0.006327f
C354 B.n174 VSUBS 0.006327f
C355 B.n175 VSUBS 0.006327f
C356 B.n176 VSUBS 0.006327f
C357 B.n177 VSUBS 0.006327f
C358 B.n178 VSUBS 0.006327f
C359 B.n179 VSUBS 0.006327f
C360 B.n180 VSUBS 0.006327f
C361 B.n181 VSUBS 0.006327f
C362 B.n182 VSUBS 0.006327f
C363 B.n183 VSUBS 0.006327f
C364 B.n184 VSUBS 0.006327f
C365 B.n185 VSUBS 0.006327f
C366 B.n186 VSUBS 0.006327f
C367 B.n187 VSUBS 0.006327f
C368 B.n188 VSUBS 0.006327f
C369 B.n189 VSUBS 0.006327f
C370 B.n190 VSUBS 0.006327f
C371 B.n191 VSUBS 0.006327f
C372 B.n192 VSUBS 0.006327f
C373 B.n193 VSUBS 0.006327f
C374 B.n194 VSUBS 0.006327f
C375 B.n195 VSUBS 0.006327f
C376 B.n196 VSUBS 0.006327f
C377 B.n197 VSUBS 0.006327f
C378 B.n198 VSUBS 0.005955f
C379 B.n199 VSUBS 0.01466f
C380 B.n200 VSUBS 0.003536f
C381 B.n201 VSUBS 0.006327f
C382 B.n202 VSUBS 0.006327f
C383 B.n203 VSUBS 0.006327f
C384 B.n204 VSUBS 0.006327f
C385 B.n205 VSUBS 0.006327f
C386 B.n206 VSUBS 0.006327f
C387 B.n207 VSUBS 0.006327f
C388 B.n208 VSUBS 0.006327f
C389 B.n209 VSUBS 0.006327f
C390 B.n210 VSUBS 0.006327f
C391 B.n211 VSUBS 0.006327f
C392 B.n212 VSUBS 0.006327f
C393 B.n213 VSUBS 0.003536f
C394 B.n214 VSUBS 0.006327f
C395 B.n215 VSUBS 0.006327f
C396 B.n216 VSUBS 0.005955f
C397 B.n217 VSUBS 0.006327f
C398 B.n218 VSUBS 0.006327f
C399 B.n219 VSUBS 0.006327f
C400 B.n220 VSUBS 0.006327f
C401 B.n221 VSUBS 0.006327f
C402 B.n222 VSUBS 0.006327f
C403 B.n223 VSUBS 0.006327f
C404 B.n224 VSUBS 0.006327f
C405 B.n225 VSUBS 0.006327f
C406 B.n226 VSUBS 0.006327f
C407 B.n227 VSUBS 0.006327f
C408 B.n228 VSUBS 0.006327f
C409 B.n229 VSUBS 0.006327f
C410 B.n230 VSUBS 0.006327f
C411 B.n231 VSUBS 0.006327f
C412 B.n232 VSUBS 0.006327f
C413 B.n233 VSUBS 0.006327f
C414 B.n234 VSUBS 0.006327f
C415 B.n235 VSUBS 0.006327f
C416 B.n236 VSUBS 0.006327f
C417 B.n237 VSUBS 0.006327f
C418 B.n238 VSUBS 0.006327f
C419 B.n239 VSUBS 0.006327f
C420 B.n240 VSUBS 0.006327f
C421 B.n241 VSUBS 0.006327f
C422 B.n242 VSUBS 0.006327f
C423 B.n243 VSUBS 0.006327f
C424 B.n244 VSUBS 0.006327f
C425 B.n245 VSUBS 0.006327f
C426 B.n246 VSUBS 0.006327f
C427 B.n247 VSUBS 0.006327f
C428 B.n248 VSUBS 0.006327f
C429 B.n249 VSUBS 0.006327f
C430 B.n250 VSUBS 0.006327f
C431 B.n251 VSUBS 0.006327f
C432 B.n252 VSUBS 0.006327f
C433 B.n253 VSUBS 0.006327f
C434 B.n254 VSUBS 0.014694f
C435 B.n255 VSUBS 0.014694f
C436 B.n256 VSUBS 0.014337f
C437 B.n257 VSUBS 0.006327f
C438 B.n258 VSUBS 0.006327f
C439 B.n259 VSUBS 0.006327f
C440 B.n260 VSUBS 0.006327f
C441 B.n261 VSUBS 0.006327f
C442 B.n262 VSUBS 0.006327f
C443 B.n263 VSUBS 0.006327f
C444 B.n264 VSUBS 0.006327f
C445 B.n265 VSUBS 0.006327f
C446 B.n266 VSUBS 0.006327f
C447 B.n267 VSUBS 0.006327f
C448 B.n268 VSUBS 0.006327f
C449 B.n269 VSUBS 0.006327f
C450 B.n270 VSUBS 0.006327f
C451 B.n271 VSUBS 0.006327f
C452 B.n272 VSUBS 0.006327f
C453 B.n273 VSUBS 0.006327f
C454 B.n274 VSUBS 0.006327f
C455 B.n275 VSUBS 0.006327f
C456 B.n276 VSUBS 0.006327f
C457 B.n277 VSUBS 0.006327f
C458 B.n278 VSUBS 0.006327f
C459 B.n279 VSUBS 0.006327f
C460 B.n280 VSUBS 0.006327f
C461 B.n281 VSUBS 0.006327f
C462 B.n282 VSUBS 0.006327f
C463 B.n283 VSUBS 0.006327f
C464 B.n284 VSUBS 0.006327f
C465 B.n285 VSUBS 0.006327f
C466 B.n286 VSUBS 0.006327f
C467 B.n287 VSUBS 0.006327f
C468 B.n288 VSUBS 0.006327f
C469 B.n289 VSUBS 0.006327f
C470 B.n290 VSUBS 0.006327f
C471 B.n291 VSUBS 0.006327f
C472 B.n292 VSUBS 0.006327f
C473 B.n293 VSUBS 0.006327f
C474 B.n294 VSUBS 0.006327f
C475 B.n295 VSUBS 0.006327f
C476 B.n296 VSUBS 0.006327f
C477 B.n297 VSUBS 0.006327f
C478 B.n298 VSUBS 0.006327f
C479 B.n299 VSUBS 0.006327f
C480 B.n300 VSUBS 0.006327f
C481 B.n301 VSUBS 0.006327f
C482 B.n302 VSUBS 0.006327f
C483 B.n303 VSUBS 0.006327f
C484 B.n304 VSUBS 0.006327f
C485 B.n305 VSUBS 0.006327f
C486 B.n306 VSUBS 0.006327f
C487 B.n307 VSUBS 0.006327f
C488 B.n308 VSUBS 0.006327f
C489 B.n309 VSUBS 0.006327f
C490 B.n310 VSUBS 0.006327f
C491 B.n311 VSUBS 0.006327f
C492 B.n312 VSUBS 0.006327f
C493 B.n313 VSUBS 0.006327f
C494 B.n314 VSUBS 0.006327f
C495 B.n315 VSUBS 0.006327f
C496 B.n316 VSUBS 0.006327f
C497 B.n317 VSUBS 0.006327f
C498 B.n318 VSUBS 0.006327f
C499 B.n319 VSUBS 0.006327f
C500 B.n320 VSUBS 0.006327f
C501 B.n321 VSUBS 0.006327f
C502 B.n322 VSUBS 0.006327f
C503 B.n323 VSUBS 0.006327f
C504 B.n324 VSUBS 0.006327f
C505 B.n325 VSUBS 0.006327f
C506 B.n326 VSUBS 0.006327f
C507 B.n327 VSUBS 0.006327f
C508 B.n328 VSUBS 0.014337f
C509 B.n329 VSUBS 0.014694f
C510 B.n330 VSUBS 0.013924f
C511 B.n331 VSUBS 0.006327f
C512 B.n332 VSUBS 0.006327f
C513 B.n333 VSUBS 0.006327f
C514 B.n334 VSUBS 0.006327f
C515 B.n335 VSUBS 0.006327f
C516 B.n336 VSUBS 0.006327f
C517 B.n337 VSUBS 0.006327f
C518 B.n338 VSUBS 0.006327f
C519 B.n339 VSUBS 0.006327f
C520 B.n340 VSUBS 0.006327f
C521 B.n341 VSUBS 0.006327f
C522 B.n342 VSUBS 0.006327f
C523 B.n343 VSUBS 0.006327f
C524 B.n344 VSUBS 0.006327f
C525 B.n345 VSUBS 0.006327f
C526 B.n346 VSUBS 0.006327f
C527 B.n347 VSUBS 0.006327f
C528 B.n348 VSUBS 0.006327f
C529 B.n349 VSUBS 0.006327f
C530 B.n350 VSUBS 0.006327f
C531 B.n351 VSUBS 0.006327f
C532 B.n352 VSUBS 0.006327f
C533 B.n353 VSUBS 0.006327f
C534 B.n354 VSUBS 0.006327f
C535 B.n355 VSUBS 0.006327f
C536 B.n356 VSUBS 0.006327f
C537 B.n357 VSUBS 0.006327f
C538 B.n358 VSUBS 0.006327f
C539 B.n359 VSUBS 0.006327f
C540 B.n360 VSUBS 0.006327f
C541 B.n361 VSUBS 0.006327f
C542 B.n362 VSUBS 0.006327f
C543 B.n363 VSUBS 0.006327f
C544 B.n364 VSUBS 0.006327f
C545 B.n365 VSUBS 0.006327f
C546 B.n366 VSUBS 0.006327f
C547 B.n367 VSUBS 0.006327f
C548 B.n368 VSUBS 0.005955f
C549 B.n369 VSUBS 0.006327f
C550 B.n370 VSUBS 0.006327f
C551 B.n371 VSUBS 0.006327f
C552 B.n372 VSUBS 0.006327f
C553 B.n373 VSUBS 0.006327f
C554 B.n374 VSUBS 0.006327f
C555 B.n375 VSUBS 0.006327f
C556 B.n376 VSUBS 0.006327f
C557 B.n377 VSUBS 0.006327f
C558 B.n378 VSUBS 0.006327f
C559 B.n379 VSUBS 0.006327f
C560 B.n380 VSUBS 0.006327f
C561 B.n381 VSUBS 0.006327f
C562 B.n382 VSUBS 0.006327f
C563 B.n383 VSUBS 0.006327f
C564 B.n384 VSUBS 0.003536f
C565 B.n385 VSUBS 0.01466f
C566 B.n386 VSUBS 0.005955f
C567 B.n387 VSUBS 0.006327f
C568 B.n388 VSUBS 0.006327f
C569 B.n389 VSUBS 0.006327f
C570 B.n390 VSUBS 0.006327f
C571 B.n391 VSUBS 0.006327f
C572 B.n392 VSUBS 0.006327f
C573 B.n393 VSUBS 0.006327f
C574 B.n394 VSUBS 0.006327f
C575 B.n395 VSUBS 0.006327f
C576 B.n396 VSUBS 0.006327f
C577 B.n397 VSUBS 0.006327f
C578 B.n398 VSUBS 0.006327f
C579 B.n399 VSUBS 0.006327f
C580 B.n400 VSUBS 0.006327f
C581 B.n401 VSUBS 0.006327f
C582 B.n402 VSUBS 0.006327f
C583 B.n403 VSUBS 0.006327f
C584 B.n404 VSUBS 0.006327f
C585 B.n405 VSUBS 0.006327f
C586 B.n406 VSUBS 0.006327f
C587 B.n407 VSUBS 0.006327f
C588 B.n408 VSUBS 0.006327f
C589 B.n409 VSUBS 0.006327f
C590 B.n410 VSUBS 0.006327f
C591 B.n411 VSUBS 0.006327f
C592 B.n412 VSUBS 0.006327f
C593 B.n413 VSUBS 0.006327f
C594 B.n414 VSUBS 0.006327f
C595 B.n415 VSUBS 0.006327f
C596 B.n416 VSUBS 0.006327f
C597 B.n417 VSUBS 0.006327f
C598 B.n418 VSUBS 0.006327f
C599 B.n419 VSUBS 0.006327f
C600 B.n420 VSUBS 0.006327f
C601 B.n421 VSUBS 0.006327f
C602 B.n422 VSUBS 0.006327f
C603 B.n423 VSUBS 0.006327f
C604 B.n424 VSUBS 0.006327f
C605 B.n425 VSUBS 0.014694f
C606 B.n426 VSUBS 0.014337f
C607 B.n427 VSUBS 0.014337f
C608 B.n428 VSUBS 0.006327f
C609 B.n429 VSUBS 0.006327f
C610 B.n430 VSUBS 0.006327f
C611 B.n431 VSUBS 0.006327f
C612 B.n432 VSUBS 0.006327f
C613 B.n433 VSUBS 0.006327f
C614 B.n434 VSUBS 0.006327f
C615 B.n435 VSUBS 0.006327f
C616 B.n436 VSUBS 0.006327f
C617 B.n437 VSUBS 0.006327f
C618 B.n438 VSUBS 0.006327f
C619 B.n439 VSUBS 0.006327f
C620 B.n440 VSUBS 0.006327f
C621 B.n441 VSUBS 0.006327f
C622 B.n442 VSUBS 0.006327f
C623 B.n443 VSUBS 0.006327f
C624 B.n444 VSUBS 0.006327f
C625 B.n445 VSUBS 0.006327f
C626 B.n446 VSUBS 0.006327f
C627 B.n447 VSUBS 0.006327f
C628 B.n448 VSUBS 0.006327f
C629 B.n449 VSUBS 0.006327f
C630 B.n450 VSUBS 0.006327f
C631 B.n451 VSUBS 0.006327f
C632 B.n452 VSUBS 0.006327f
C633 B.n453 VSUBS 0.006327f
C634 B.n454 VSUBS 0.006327f
C635 B.n455 VSUBS 0.006327f
C636 B.n456 VSUBS 0.006327f
C637 B.n457 VSUBS 0.006327f
C638 B.n458 VSUBS 0.006327f
C639 B.n459 VSUBS 0.006327f
C640 B.n460 VSUBS 0.006327f
C641 B.n461 VSUBS 0.006327f
C642 B.n462 VSUBS 0.006327f
C643 B.n463 VSUBS 0.014328f
.ends

