* NGSPICE file created from diff_pair_sample_0244.ext - technology: sky130A

.subckt diff_pair_sample_0244 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=0 ps=0 w=9.3 l=2.52
X1 VTAIL.t7 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=1.5345 ps=9.63 w=9.3 l=2.52
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=0 ps=0 w=9.3 l=2.52
X3 VDD2.t2 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5345 pd=9.63 as=3.627 ps=19.38 w=9.3 l=2.52
X4 VTAIL.t5 VN.t2 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=1.5345 ps=9.63 w=9.3 l=2.52
X5 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5345 pd=9.63 as=3.627 ps=19.38 w=9.3 l=2.52
X6 VDD2.t1 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5345 pd=9.63 as=3.627 ps=19.38 w=9.3 l=2.52
X7 VDD1.t2 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5345 pd=9.63 as=3.627 ps=19.38 w=9.3 l=2.52
X8 VTAIL.t1 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=1.5345 ps=9.63 w=9.3 l=2.52
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=0 ps=0 w=9.3 l=2.52
X10 VTAIL.t0 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=1.5345 ps=9.63 w=9.3 l=2.52
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.627 pd=19.38 as=0 ps=0 w=9.3 l=2.52
R0 B.n663 B.n662 585
R1 B.n664 B.n663 585
R2 B.n258 B.n101 585
R3 B.n257 B.n256 585
R4 B.n255 B.n254 585
R5 B.n253 B.n252 585
R6 B.n251 B.n250 585
R7 B.n249 B.n248 585
R8 B.n247 B.n246 585
R9 B.n245 B.n244 585
R10 B.n243 B.n242 585
R11 B.n241 B.n240 585
R12 B.n239 B.n238 585
R13 B.n237 B.n236 585
R14 B.n235 B.n234 585
R15 B.n233 B.n232 585
R16 B.n231 B.n230 585
R17 B.n229 B.n228 585
R18 B.n227 B.n226 585
R19 B.n225 B.n224 585
R20 B.n223 B.n222 585
R21 B.n221 B.n220 585
R22 B.n219 B.n218 585
R23 B.n217 B.n216 585
R24 B.n215 B.n214 585
R25 B.n213 B.n212 585
R26 B.n211 B.n210 585
R27 B.n209 B.n208 585
R28 B.n207 B.n206 585
R29 B.n205 B.n204 585
R30 B.n203 B.n202 585
R31 B.n201 B.n200 585
R32 B.n199 B.n198 585
R33 B.n197 B.n196 585
R34 B.n195 B.n194 585
R35 B.n192 B.n191 585
R36 B.n190 B.n189 585
R37 B.n188 B.n187 585
R38 B.n186 B.n185 585
R39 B.n184 B.n183 585
R40 B.n182 B.n181 585
R41 B.n180 B.n179 585
R42 B.n178 B.n177 585
R43 B.n176 B.n175 585
R44 B.n174 B.n173 585
R45 B.n172 B.n171 585
R46 B.n170 B.n169 585
R47 B.n168 B.n167 585
R48 B.n166 B.n165 585
R49 B.n164 B.n163 585
R50 B.n162 B.n161 585
R51 B.n160 B.n159 585
R52 B.n158 B.n157 585
R53 B.n156 B.n155 585
R54 B.n154 B.n153 585
R55 B.n152 B.n151 585
R56 B.n150 B.n149 585
R57 B.n148 B.n147 585
R58 B.n146 B.n145 585
R59 B.n144 B.n143 585
R60 B.n142 B.n141 585
R61 B.n140 B.n139 585
R62 B.n138 B.n137 585
R63 B.n136 B.n135 585
R64 B.n134 B.n133 585
R65 B.n132 B.n131 585
R66 B.n130 B.n129 585
R67 B.n128 B.n127 585
R68 B.n126 B.n125 585
R69 B.n124 B.n123 585
R70 B.n122 B.n121 585
R71 B.n120 B.n119 585
R72 B.n118 B.n117 585
R73 B.n116 B.n115 585
R74 B.n114 B.n113 585
R75 B.n112 B.n111 585
R76 B.n110 B.n109 585
R77 B.n108 B.n107 585
R78 B.n661 B.n62 585
R79 B.n665 B.n62 585
R80 B.n660 B.n61 585
R81 B.n666 B.n61 585
R82 B.n659 B.n658 585
R83 B.n658 B.n57 585
R84 B.n657 B.n56 585
R85 B.n672 B.n56 585
R86 B.n656 B.n55 585
R87 B.n673 B.n55 585
R88 B.n655 B.n54 585
R89 B.n674 B.n54 585
R90 B.n654 B.n653 585
R91 B.n653 B.n50 585
R92 B.n652 B.n49 585
R93 B.n680 B.n49 585
R94 B.n651 B.n48 585
R95 B.n681 B.n48 585
R96 B.n650 B.n47 585
R97 B.n682 B.n47 585
R98 B.n649 B.n648 585
R99 B.n648 B.n43 585
R100 B.n647 B.n42 585
R101 B.n688 B.n42 585
R102 B.n646 B.n41 585
R103 B.n689 B.n41 585
R104 B.n645 B.n40 585
R105 B.n690 B.n40 585
R106 B.n644 B.n643 585
R107 B.n643 B.n36 585
R108 B.n642 B.n35 585
R109 B.n696 B.n35 585
R110 B.n641 B.n34 585
R111 B.n697 B.n34 585
R112 B.n640 B.n33 585
R113 B.n698 B.n33 585
R114 B.n639 B.n638 585
R115 B.n638 B.n32 585
R116 B.n637 B.n28 585
R117 B.n704 B.n28 585
R118 B.n636 B.n27 585
R119 B.n705 B.n27 585
R120 B.n635 B.n26 585
R121 B.n706 B.n26 585
R122 B.n634 B.n633 585
R123 B.n633 B.n22 585
R124 B.n632 B.n21 585
R125 B.n712 B.n21 585
R126 B.n631 B.n20 585
R127 B.n713 B.n20 585
R128 B.n630 B.n19 585
R129 B.n714 B.n19 585
R130 B.n629 B.n628 585
R131 B.n628 B.n15 585
R132 B.n627 B.n14 585
R133 B.n720 B.n14 585
R134 B.n626 B.n13 585
R135 B.n721 B.n13 585
R136 B.n625 B.n12 585
R137 B.n722 B.n12 585
R138 B.n624 B.n623 585
R139 B.n623 B.n8 585
R140 B.n622 B.n7 585
R141 B.n728 B.n7 585
R142 B.n621 B.n6 585
R143 B.n729 B.n6 585
R144 B.n620 B.n5 585
R145 B.n730 B.n5 585
R146 B.n619 B.n618 585
R147 B.n618 B.n4 585
R148 B.n617 B.n259 585
R149 B.n617 B.n616 585
R150 B.n607 B.n260 585
R151 B.n261 B.n260 585
R152 B.n609 B.n608 585
R153 B.n610 B.n609 585
R154 B.n606 B.n266 585
R155 B.n266 B.n265 585
R156 B.n605 B.n604 585
R157 B.n604 B.n603 585
R158 B.n268 B.n267 585
R159 B.n269 B.n268 585
R160 B.n596 B.n595 585
R161 B.n597 B.n596 585
R162 B.n594 B.n274 585
R163 B.n274 B.n273 585
R164 B.n593 B.n592 585
R165 B.n592 B.n591 585
R166 B.n276 B.n275 585
R167 B.n277 B.n276 585
R168 B.n584 B.n583 585
R169 B.n585 B.n584 585
R170 B.n582 B.n282 585
R171 B.n282 B.n281 585
R172 B.n581 B.n580 585
R173 B.n580 B.n579 585
R174 B.n284 B.n283 585
R175 B.n572 B.n284 585
R176 B.n571 B.n570 585
R177 B.n573 B.n571 585
R178 B.n569 B.n289 585
R179 B.n289 B.n288 585
R180 B.n568 B.n567 585
R181 B.n567 B.n566 585
R182 B.n291 B.n290 585
R183 B.n292 B.n291 585
R184 B.n559 B.n558 585
R185 B.n560 B.n559 585
R186 B.n557 B.n297 585
R187 B.n297 B.n296 585
R188 B.n556 B.n555 585
R189 B.n555 B.n554 585
R190 B.n299 B.n298 585
R191 B.n300 B.n299 585
R192 B.n547 B.n546 585
R193 B.n548 B.n547 585
R194 B.n545 B.n305 585
R195 B.n305 B.n304 585
R196 B.n544 B.n543 585
R197 B.n543 B.n542 585
R198 B.n307 B.n306 585
R199 B.n308 B.n307 585
R200 B.n535 B.n534 585
R201 B.n536 B.n535 585
R202 B.n533 B.n313 585
R203 B.n313 B.n312 585
R204 B.n532 B.n531 585
R205 B.n531 B.n530 585
R206 B.n315 B.n314 585
R207 B.n316 B.n315 585
R208 B.n523 B.n522 585
R209 B.n524 B.n523 585
R210 B.n521 B.n321 585
R211 B.n321 B.n320 585
R212 B.n515 B.n514 585
R213 B.n513 B.n361 585
R214 B.n512 B.n360 585
R215 B.n517 B.n360 585
R216 B.n511 B.n510 585
R217 B.n509 B.n508 585
R218 B.n507 B.n506 585
R219 B.n505 B.n504 585
R220 B.n503 B.n502 585
R221 B.n501 B.n500 585
R222 B.n499 B.n498 585
R223 B.n497 B.n496 585
R224 B.n495 B.n494 585
R225 B.n493 B.n492 585
R226 B.n491 B.n490 585
R227 B.n489 B.n488 585
R228 B.n487 B.n486 585
R229 B.n485 B.n484 585
R230 B.n483 B.n482 585
R231 B.n481 B.n480 585
R232 B.n479 B.n478 585
R233 B.n477 B.n476 585
R234 B.n475 B.n474 585
R235 B.n473 B.n472 585
R236 B.n471 B.n470 585
R237 B.n469 B.n468 585
R238 B.n467 B.n466 585
R239 B.n465 B.n464 585
R240 B.n463 B.n462 585
R241 B.n461 B.n460 585
R242 B.n459 B.n458 585
R243 B.n457 B.n456 585
R244 B.n455 B.n454 585
R245 B.n453 B.n452 585
R246 B.n451 B.n450 585
R247 B.n448 B.n447 585
R248 B.n446 B.n445 585
R249 B.n444 B.n443 585
R250 B.n442 B.n441 585
R251 B.n440 B.n439 585
R252 B.n438 B.n437 585
R253 B.n436 B.n435 585
R254 B.n434 B.n433 585
R255 B.n432 B.n431 585
R256 B.n430 B.n429 585
R257 B.n428 B.n427 585
R258 B.n426 B.n425 585
R259 B.n424 B.n423 585
R260 B.n422 B.n421 585
R261 B.n420 B.n419 585
R262 B.n418 B.n417 585
R263 B.n416 B.n415 585
R264 B.n414 B.n413 585
R265 B.n412 B.n411 585
R266 B.n410 B.n409 585
R267 B.n408 B.n407 585
R268 B.n406 B.n405 585
R269 B.n404 B.n403 585
R270 B.n402 B.n401 585
R271 B.n400 B.n399 585
R272 B.n398 B.n397 585
R273 B.n396 B.n395 585
R274 B.n394 B.n393 585
R275 B.n392 B.n391 585
R276 B.n390 B.n389 585
R277 B.n388 B.n387 585
R278 B.n386 B.n385 585
R279 B.n384 B.n383 585
R280 B.n382 B.n381 585
R281 B.n380 B.n379 585
R282 B.n378 B.n377 585
R283 B.n376 B.n375 585
R284 B.n374 B.n373 585
R285 B.n372 B.n371 585
R286 B.n370 B.n369 585
R287 B.n368 B.n367 585
R288 B.n323 B.n322 585
R289 B.n520 B.n519 585
R290 B.n319 B.n318 585
R291 B.n320 B.n319 585
R292 B.n526 B.n525 585
R293 B.n525 B.n524 585
R294 B.n527 B.n317 585
R295 B.n317 B.n316 585
R296 B.n529 B.n528 585
R297 B.n530 B.n529 585
R298 B.n311 B.n310 585
R299 B.n312 B.n311 585
R300 B.n538 B.n537 585
R301 B.n537 B.n536 585
R302 B.n539 B.n309 585
R303 B.n309 B.n308 585
R304 B.n541 B.n540 585
R305 B.n542 B.n541 585
R306 B.n303 B.n302 585
R307 B.n304 B.n303 585
R308 B.n550 B.n549 585
R309 B.n549 B.n548 585
R310 B.n551 B.n301 585
R311 B.n301 B.n300 585
R312 B.n553 B.n552 585
R313 B.n554 B.n553 585
R314 B.n295 B.n294 585
R315 B.n296 B.n295 585
R316 B.n562 B.n561 585
R317 B.n561 B.n560 585
R318 B.n563 B.n293 585
R319 B.n293 B.n292 585
R320 B.n565 B.n564 585
R321 B.n566 B.n565 585
R322 B.n287 B.n286 585
R323 B.n288 B.n287 585
R324 B.n575 B.n574 585
R325 B.n574 B.n573 585
R326 B.n576 B.n285 585
R327 B.n572 B.n285 585
R328 B.n578 B.n577 585
R329 B.n579 B.n578 585
R330 B.n280 B.n279 585
R331 B.n281 B.n280 585
R332 B.n587 B.n586 585
R333 B.n586 B.n585 585
R334 B.n588 B.n278 585
R335 B.n278 B.n277 585
R336 B.n590 B.n589 585
R337 B.n591 B.n590 585
R338 B.n272 B.n271 585
R339 B.n273 B.n272 585
R340 B.n599 B.n598 585
R341 B.n598 B.n597 585
R342 B.n600 B.n270 585
R343 B.n270 B.n269 585
R344 B.n602 B.n601 585
R345 B.n603 B.n602 585
R346 B.n264 B.n263 585
R347 B.n265 B.n264 585
R348 B.n612 B.n611 585
R349 B.n611 B.n610 585
R350 B.n613 B.n262 585
R351 B.n262 B.n261 585
R352 B.n615 B.n614 585
R353 B.n616 B.n615 585
R354 B.n2 B.n0 585
R355 B.n4 B.n2 585
R356 B.n3 B.n1 585
R357 B.n729 B.n3 585
R358 B.n727 B.n726 585
R359 B.n728 B.n727 585
R360 B.n725 B.n9 585
R361 B.n9 B.n8 585
R362 B.n724 B.n723 585
R363 B.n723 B.n722 585
R364 B.n11 B.n10 585
R365 B.n721 B.n11 585
R366 B.n719 B.n718 585
R367 B.n720 B.n719 585
R368 B.n717 B.n16 585
R369 B.n16 B.n15 585
R370 B.n716 B.n715 585
R371 B.n715 B.n714 585
R372 B.n18 B.n17 585
R373 B.n713 B.n18 585
R374 B.n711 B.n710 585
R375 B.n712 B.n711 585
R376 B.n709 B.n23 585
R377 B.n23 B.n22 585
R378 B.n708 B.n707 585
R379 B.n707 B.n706 585
R380 B.n25 B.n24 585
R381 B.n705 B.n25 585
R382 B.n703 B.n702 585
R383 B.n704 B.n703 585
R384 B.n701 B.n29 585
R385 B.n32 B.n29 585
R386 B.n700 B.n699 585
R387 B.n699 B.n698 585
R388 B.n31 B.n30 585
R389 B.n697 B.n31 585
R390 B.n695 B.n694 585
R391 B.n696 B.n695 585
R392 B.n693 B.n37 585
R393 B.n37 B.n36 585
R394 B.n692 B.n691 585
R395 B.n691 B.n690 585
R396 B.n39 B.n38 585
R397 B.n689 B.n39 585
R398 B.n687 B.n686 585
R399 B.n688 B.n687 585
R400 B.n685 B.n44 585
R401 B.n44 B.n43 585
R402 B.n684 B.n683 585
R403 B.n683 B.n682 585
R404 B.n46 B.n45 585
R405 B.n681 B.n46 585
R406 B.n679 B.n678 585
R407 B.n680 B.n679 585
R408 B.n677 B.n51 585
R409 B.n51 B.n50 585
R410 B.n676 B.n675 585
R411 B.n675 B.n674 585
R412 B.n53 B.n52 585
R413 B.n673 B.n53 585
R414 B.n671 B.n670 585
R415 B.n672 B.n671 585
R416 B.n669 B.n58 585
R417 B.n58 B.n57 585
R418 B.n668 B.n667 585
R419 B.n667 B.n666 585
R420 B.n60 B.n59 585
R421 B.n665 B.n60 585
R422 B.n732 B.n731 585
R423 B.n731 B.n730 585
R424 B.n515 B.n319 535.745
R425 B.n107 B.n60 535.745
R426 B.n519 B.n321 535.745
R427 B.n663 B.n62 535.745
R428 B.n364 B.t8 296.863
R429 B.n362 B.t15 296.863
R430 B.n104 B.t4 296.863
R431 B.n102 B.t12 296.863
R432 B.n364 B.t11 290.82
R433 B.n102 B.t13 290.82
R434 B.n362 B.t17 290.82
R435 B.n104 B.t6 290.82
R436 B.n664 B.n100 256.663
R437 B.n664 B.n99 256.663
R438 B.n664 B.n98 256.663
R439 B.n664 B.n97 256.663
R440 B.n664 B.n96 256.663
R441 B.n664 B.n95 256.663
R442 B.n664 B.n94 256.663
R443 B.n664 B.n93 256.663
R444 B.n664 B.n92 256.663
R445 B.n664 B.n91 256.663
R446 B.n664 B.n90 256.663
R447 B.n664 B.n89 256.663
R448 B.n664 B.n88 256.663
R449 B.n664 B.n87 256.663
R450 B.n664 B.n86 256.663
R451 B.n664 B.n85 256.663
R452 B.n664 B.n84 256.663
R453 B.n664 B.n83 256.663
R454 B.n664 B.n82 256.663
R455 B.n664 B.n81 256.663
R456 B.n664 B.n80 256.663
R457 B.n664 B.n79 256.663
R458 B.n664 B.n78 256.663
R459 B.n664 B.n77 256.663
R460 B.n664 B.n76 256.663
R461 B.n664 B.n75 256.663
R462 B.n664 B.n74 256.663
R463 B.n664 B.n73 256.663
R464 B.n664 B.n72 256.663
R465 B.n664 B.n71 256.663
R466 B.n664 B.n70 256.663
R467 B.n664 B.n69 256.663
R468 B.n664 B.n68 256.663
R469 B.n664 B.n67 256.663
R470 B.n664 B.n66 256.663
R471 B.n664 B.n65 256.663
R472 B.n664 B.n64 256.663
R473 B.n664 B.n63 256.663
R474 B.n517 B.n516 256.663
R475 B.n517 B.n324 256.663
R476 B.n517 B.n325 256.663
R477 B.n517 B.n326 256.663
R478 B.n517 B.n327 256.663
R479 B.n517 B.n328 256.663
R480 B.n517 B.n329 256.663
R481 B.n517 B.n330 256.663
R482 B.n517 B.n331 256.663
R483 B.n517 B.n332 256.663
R484 B.n517 B.n333 256.663
R485 B.n517 B.n334 256.663
R486 B.n517 B.n335 256.663
R487 B.n517 B.n336 256.663
R488 B.n517 B.n337 256.663
R489 B.n517 B.n338 256.663
R490 B.n517 B.n339 256.663
R491 B.n517 B.n340 256.663
R492 B.n517 B.n341 256.663
R493 B.n517 B.n342 256.663
R494 B.n517 B.n343 256.663
R495 B.n517 B.n344 256.663
R496 B.n517 B.n345 256.663
R497 B.n517 B.n346 256.663
R498 B.n517 B.n347 256.663
R499 B.n517 B.n348 256.663
R500 B.n517 B.n349 256.663
R501 B.n517 B.n350 256.663
R502 B.n517 B.n351 256.663
R503 B.n517 B.n352 256.663
R504 B.n517 B.n353 256.663
R505 B.n517 B.n354 256.663
R506 B.n517 B.n355 256.663
R507 B.n517 B.n356 256.663
R508 B.n517 B.n357 256.663
R509 B.n517 B.n358 256.663
R510 B.n517 B.n359 256.663
R511 B.n518 B.n517 256.663
R512 B.n365 B.t10 235.548
R513 B.n103 B.t14 235.548
R514 B.n363 B.t16 235.548
R515 B.n105 B.t7 235.548
R516 B.n525 B.n319 163.367
R517 B.n525 B.n317 163.367
R518 B.n529 B.n317 163.367
R519 B.n529 B.n311 163.367
R520 B.n537 B.n311 163.367
R521 B.n537 B.n309 163.367
R522 B.n541 B.n309 163.367
R523 B.n541 B.n303 163.367
R524 B.n549 B.n303 163.367
R525 B.n549 B.n301 163.367
R526 B.n553 B.n301 163.367
R527 B.n553 B.n295 163.367
R528 B.n561 B.n295 163.367
R529 B.n561 B.n293 163.367
R530 B.n565 B.n293 163.367
R531 B.n565 B.n287 163.367
R532 B.n574 B.n287 163.367
R533 B.n574 B.n285 163.367
R534 B.n578 B.n285 163.367
R535 B.n578 B.n280 163.367
R536 B.n586 B.n280 163.367
R537 B.n586 B.n278 163.367
R538 B.n590 B.n278 163.367
R539 B.n590 B.n272 163.367
R540 B.n598 B.n272 163.367
R541 B.n598 B.n270 163.367
R542 B.n602 B.n270 163.367
R543 B.n602 B.n264 163.367
R544 B.n611 B.n264 163.367
R545 B.n611 B.n262 163.367
R546 B.n615 B.n262 163.367
R547 B.n615 B.n2 163.367
R548 B.n731 B.n2 163.367
R549 B.n731 B.n3 163.367
R550 B.n727 B.n3 163.367
R551 B.n727 B.n9 163.367
R552 B.n723 B.n9 163.367
R553 B.n723 B.n11 163.367
R554 B.n719 B.n11 163.367
R555 B.n719 B.n16 163.367
R556 B.n715 B.n16 163.367
R557 B.n715 B.n18 163.367
R558 B.n711 B.n18 163.367
R559 B.n711 B.n23 163.367
R560 B.n707 B.n23 163.367
R561 B.n707 B.n25 163.367
R562 B.n703 B.n25 163.367
R563 B.n703 B.n29 163.367
R564 B.n699 B.n29 163.367
R565 B.n699 B.n31 163.367
R566 B.n695 B.n31 163.367
R567 B.n695 B.n37 163.367
R568 B.n691 B.n37 163.367
R569 B.n691 B.n39 163.367
R570 B.n687 B.n39 163.367
R571 B.n687 B.n44 163.367
R572 B.n683 B.n44 163.367
R573 B.n683 B.n46 163.367
R574 B.n679 B.n46 163.367
R575 B.n679 B.n51 163.367
R576 B.n675 B.n51 163.367
R577 B.n675 B.n53 163.367
R578 B.n671 B.n53 163.367
R579 B.n671 B.n58 163.367
R580 B.n667 B.n58 163.367
R581 B.n667 B.n60 163.367
R582 B.n361 B.n360 163.367
R583 B.n510 B.n360 163.367
R584 B.n508 B.n507 163.367
R585 B.n504 B.n503 163.367
R586 B.n500 B.n499 163.367
R587 B.n496 B.n495 163.367
R588 B.n492 B.n491 163.367
R589 B.n488 B.n487 163.367
R590 B.n484 B.n483 163.367
R591 B.n480 B.n479 163.367
R592 B.n476 B.n475 163.367
R593 B.n472 B.n471 163.367
R594 B.n468 B.n467 163.367
R595 B.n464 B.n463 163.367
R596 B.n460 B.n459 163.367
R597 B.n456 B.n455 163.367
R598 B.n452 B.n451 163.367
R599 B.n447 B.n446 163.367
R600 B.n443 B.n442 163.367
R601 B.n439 B.n438 163.367
R602 B.n435 B.n434 163.367
R603 B.n431 B.n430 163.367
R604 B.n427 B.n426 163.367
R605 B.n423 B.n422 163.367
R606 B.n419 B.n418 163.367
R607 B.n415 B.n414 163.367
R608 B.n411 B.n410 163.367
R609 B.n407 B.n406 163.367
R610 B.n403 B.n402 163.367
R611 B.n399 B.n398 163.367
R612 B.n395 B.n394 163.367
R613 B.n391 B.n390 163.367
R614 B.n387 B.n386 163.367
R615 B.n383 B.n382 163.367
R616 B.n379 B.n378 163.367
R617 B.n375 B.n374 163.367
R618 B.n371 B.n370 163.367
R619 B.n367 B.n323 163.367
R620 B.n523 B.n321 163.367
R621 B.n523 B.n315 163.367
R622 B.n531 B.n315 163.367
R623 B.n531 B.n313 163.367
R624 B.n535 B.n313 163.367
R625 B.n535 B.n307 163.367
R626 B.n543 B.n307 163.367
R627 B.n543 B.n305 163.367
R628 B.n547 B.n305 163.367
R629 B.n547 B.n299 163.367
R630 B.n555 B.n299 163.367
R631 B.n555 B.n297 163.367
R632 B.n559 B.n297 163.367
R633 B.n559 B.n291 163.367
R634 B.n567 B.n291 163.367
R635 B.n567 B.n289 163.367
R636 B.n571 B.n289 163.367
R637 B.n571 B.n284 163.367
R638 B.n580 B.n284 163.367
R639 B.n580 B.n282 163.367
R640 B.n584 B.n282 163.367
R641 B.n584 B.n276 163.367
R642 B.n592 B.n276 163.367
R643 B.n592 B.n274 163.367
R644 B.n596 B.n274 163.367
R645 B.n596 B.n268 163.367
R646 B.n604 B.n268 163.367
R647 B.n604 B.n266 163.367
R648 B.n609 B.n266 163.367
R649 B.n609 B.n260 163.367
R650 B.n617 B.n260 163.367
R651 B.n618 B.n617 163.367
R652 B.n618 B.n5 163.367
R653 B.n6 B.n5 163.367
R654 B.n7 B.n6 163.367
R655 B.n623 B.n7 163.367
R656 B.n623 B.n12 163.367
R657 B.n13 B.n12 163.367
R658 B.n14 B.n13 163.367
R659 B.n628 B.n14 163.367
R660 B.n628 B.n19 163.367
R661 B.n20 B.n19 163.367
R662 B.n21 B.n20 163.367
R663 B.n633 B.n21 163.367
R664 B.n633 B.n26 163.367
R665 B.n27 B.n26 163.367
R666 B.n28 B.n27 163.367
R667 B.n638 B.n28 163.367
R668 B.n638 B.n33 163.367
R669 B.n34 B.n33 163.367
R670 B.n35 B.n34 163.367
R671 B.n643 B.n35 163.367
R672 B.n643 B.n40 163.367
R673 B.n41 B.n40 163.367
R674 B.n42 B.n41 163.367
R675 B.n648 B.n42 163.367
R676 B.n648 B.n47 163.367
R677 B.n48 B.n47 163.367
R678 B.n49 B.n48 163.367
R679 B.n653 B.n49 163.367
R680 B.n653 B.n54 163.367
R681 B.n55 B.n54 163.367
R682 B.n56 B.n55 163.367
R683 B.n658 B.n56 163.367
R684 B.n658 B.n61 163.367
R685 B.n62 B.n61 163.367
R686 B.n111 B.n110 163.367
R687 B.n115 B.n114 163.367
R688 B.n119 B.n118 163.367
R689 B.n123 B.n122 163.367
R690 B.n127 B.n126 163.367
R691 B.n131 B.n130 163.367
R692 B.n135 B.n134 163.367
R693 B.n139 B.n138 163.367
R694 B.n143 B.n142 163.367
R695 B.n147 B.n146 163.367
R696 B.n151 B.n150 163.367
R697 B.n155 B.n154 163.367
R698 B.n159 B.n158 163.367
R699 B.n163 B.n162 163.367
R700 B.n167 B.n166 163.367
R701 B.n171 B.n170 163.367
R702 B.n175 B.n174 163.367
R703 B.n179 B.n178 163.367
R704 B.n183 B.n182 163.367
R705 B.n187 B.n186 163.367
R706 B.n191 B.n190 163.367
R707 B.n196 B.n195 163.367
R708 B.n200 B.n199 163.367
R709 B.n204 B.n203 163.367
R710 B.n208 B.n207 163.367
R711 B.n212 B.n211 163.367
R712 B.n216 B.n215 163.367
R713 B.n220 B.n219 163.367
R714 B.n224 B.n223 163.367
R715 B.n228 B.n227 163.367
R716 B.n232 B.n231 163.367
R717 B.n236 B.n235 163.367
R718 B.n240 B.n239 163.367
R719 B.n244 B.n243 163.367
R720 B.n248 B.n247 163.367
R721 B.n252 B.n251 163.367
R722 B.n256 B.n255 163.367
R723 B.n663 B.n101 163.367
R724 B.n517 B.n320 106.415
R725 B.n665 B.n664 106.415
R726 B.n516 B.n515 71.676
R727 B.n510 B.n324 71.676
R728 B.n507 B.n325 71.676
R729 B.n503 B.n326 71.676
R730 B.n499 B.n327 71.676
R731 B.n495 B.n328 71.676
R732 B.n491 B.n329 71.676
R733 B.n487 B.n330 71.676
R734 B.n483 B.n331 71.676
R735 B.n479 B.n332 71.676
R736 B.n475 B.n333 71.676
R737 B.n471 B.n334 71.676
R738 B.n467 B.n335 71.676
R739 B.n463 B.n336 71.676
R740 B.n459 B.n337 71.676
R741 B.n455 B.n338 71.676
R742 B.n451 B.n339 71.676
R743 B.n446 B.n340 71.676
R744 B.n442 B.n341 71.676
R745 B.n438 B.n342 71.676
R746 B.n434 B.n343 71.676
R747 B.n430 B.n344 71.676
R748 B.n426 B.n345 71.676
R749 B.n422 B.n346 71.676
R750 B.n418 B.n347 71.676
R751 B.n414 B.n348 71.676
R752 B.n410 B.n349 71.676
R753 B.n406 B.n350 71.676
R754 B.n402 B.n351 71.676
R755 B.n398 B.n352 71.676
R756 B.n394 B.n353 71.676
R757 B.n390 B.n354 71.676
R758 B.n386 B.n355 71.676
R759 B.n382 B.n356 71.676
R760 B.n378 B.n357 71.676
R761 B.n374 B.n358 71.676
R762 B.n370 B.n359 71.676
R763 B.n518 B.n323 71.676
R764 B.n107 B.n63 71.676
R765 B.n111 B.n64 71.676
R766 B.n115 B.n65 71.676
R767 B.n119 B.n66 71.676
R768 B.n123 B.n67 71.676
R769 B.n127 B.n68 71.676
R770 B.n131 B.n69 71.676
R771 B.n135 B.n70 71.676
R772 B.n139 B.n71 71.676
R773 B.n143 B.n72 71.676
R774 B.n147 B.n73 71.676
R775 B.n151 B.n74 71.676
R776 B.n155 B.n75 71.676
R777 B.n159 B.n76 71.676
R778 B.n163 B.n77 71.676
R779 B.n167 B.n78 71.676
R780 B.n171 B.n79 71.676
R781 B.n175 B.n80 71.676
R782 B.n179 B.n81 71.676
R783 B.n183 B.n82 71.676
R784 B.n187 B.n83 71.676
R785 B.n191 B.n84 71.676
R786 B.n196 B.n85 71.676
R787 B.n200 B.n86 71.676
R788 B.n204 B.n87 71.676
R789 B.n208 B.n88 71.676
R790 B.n212 B.n89 71.676
R791 B.n216 B.n90 71.676
R792 B.n220 B.n91 71.676
R793 B.n224 B.n92 71.676
R794 B.n228 B.n93 71.676
R795 B.n232 B.n94 71.676
R796 B.n236 B.n95 71.676
R797 B.n240 B.n96 71.676
R798 B.n244 B.n97 71.676
R799 B.n248 B.n98 71.676
R800 B.n252 B.n99 71.676
R801 B.n256 B.n100 71.676
R802 B.n101 B.n100 71.676
R803 B.n255 B.n99 71.676
R804 B.n251 B.n98 71.676
R805 B.n247 B.n97 71.676
R806 B.n243 B.n96 71.676
R807 B.n239 B.n95 71.676
R808 B.n235 B.n94 71.676
R809 B.n231 B.n93 71.676
R810 B.n227 B.n92 71.676
R811 B.n223 B.n91 71.676
R812 B.n219 B.n90 71.676
R813 B.n215 B.n89 71.676
R814 B.n211 B.n88 71.676
R815 B.n207 B.n87 71.676
R816 B.n203 B.n86 71.676
R817 B.n199 B.n85 71.676
R818 B.n195 B.n84 71.676
R819 B.n190 B.n83 71.676
R820 B.n186 B.n82 71.676
R821 B.n182 B.n81 71.676
R822 B.n178 B.n80 71.676
R823 B.n174 B.n79 71.676
R824 B.n170 B.n78 71.676
R825 B.n166 B.n77 71.676
R826 B.n162 B.n76 71.676
R827 B.n158 B.n75 71.676
R828 B.n154 B.n74 71.676
R829 B.n150 B.n73 71.676
R830 B.n146 B.n72 71.676
R831 B.n142 B.n71 71.676
R832 B.n138 B.n70 71.676
R833 B.n134 B.n69 71.676
R834 B.n130 B.n68 71.676
R835 B.n126 B.n67 71.676
R836 B.n122 B.n66 71.676
R837 B.n118 B.n65 71.676
R838 B.n114 B.n64 71.676
R839 B.n110 B.n63 71.676
R840 B.n516 B.n361 71.676
R841 B.n508 B.n324 71.676
R842 B.n504 B.n325 71.676
R843 B.n500 B.n326 71.676
R844 B.n496 B.n327 71.676
R845 B.n492 B.n328 71.676
R846 B.n488 B.n329 71.676
R847 B.n484 B.n330 71.676
R848 B.n480 B.n331 71.676
R849 B.n476 B.n332 71.676
R850 B.n472 B.n333 71.676
R851 B.n468 B.n334 71.676
R852 B.n464 B.n335 71.676
R853 B.n460 B.n336 71.676
R854 B.n456 B.n337 71.676
R855 B.n452 B.n338 71.676
R856 B.n447 B.n339 71.676
R857 B.n443 B.n340 71.676
R858 B.n439 B.n341 71.676
R859 B.n435 B.n342 71.676
R860 B.n431 B.n343 71.676
R861 B.n427 B.n344 71.676
R862 B.n423 B.n345 71.676
R863 B.n419 B.n346 71.676
R864 B.n415 B.n347 71.676
R865 B.n411 B.n348 71.676
R866 B.n407 B.n349 71.676
R867 B.n403 B.n350 71.676
R868 B.n399 B.n351 71.676
R869 B.n395 B.n352 71.676
R870 B.n391 B.n353 71.676
R871 B.n387 B.n354 71.676
R872 B.n383 B.n355 71.676
R873 B.n379 B.n356 71.676
R874 B.n375 B.n357 71.676
R875 B.n371 B.n358 71.676
R876 B.n367 B.n359 71.676
R877 B.n519 B.n518 71.676
R878 B.n366 B.n365 59.5399
R879 B.n449 B.n363 59.5399
R880 B.n106 B.n105 59.5399
R881 B.n193 B.n103 59.5399
R882 B.n365 B.n364 55.2732
R883 B.n363 B.n362 55.2732
R884 B.n105 B.n104 55.2732
R885 B.n103 B.n102 55.2732
R886 B.n524 B.n320 51.3213
R887 B.n524 B.n316 51.3213
R888 B.n530 B.n316 51.3213
R889 B.n530 B.n312 51.3213
R890 B.n536 B.n312 51.3213
R891 B.n536 B.n308 51.3213
R892 B.n542 B.n308 51.3213
R893 B.n548 B.n304 51.3213
R894 B.n548 B.n300 51.3213
R895 B.n554 B.n300 51.3213
R896 B.n554 B.n296 51.3213
R897 B.n560 B.n296 51.3213
R898 B.n560 B.n292 51.3213
R899 B.n566 B.n292 51.3213
R900 B.n566 B.n288 51.3213
R901 B.n573 B.n288 51.3213
R902 B.n573 B.n572 51.3213
R903 B.n579 B.n281 51.3213
R904 B.n585 B.n281 51.3213
R905 B.n585 B.n277 51.3213
R906 B.n591 B.n277 51.3213
R907 B.n591 B.n273 51.3213
R908 B.n597 B.n273 51.3213
R909 B.n597 B.n269 51.3213
R910 B.n603 B.n269 51.3213
R911 B.n610 B.n265 51.3213
R912 B.n610 B.n261 51.3213
R913 B.n616 B.n261 51.3213
R914 B.n616 B.n4 51.3213
R915 B.n730 B.n4 51.3213
R916 B.n730 B.n729 51.3213
R917 B.n729 B.n728 51.3213
R918 B.n728 B.n8 51.3213
R919 B.n722 B.n8 51.3213
R920 B.n722 B.n721 51.3213
R921 B.n720 B.n15 51.3213
R922 B.n714 B.n15 51.3213
R923 B.n714 B.n713 51.3213
R924 B.n713 B.n712 51.3213
R925 B.n712 B.n22 51.3213
R926 B.n706 B.n22 51.3213
R927 B.n706 B.n705 51.3213
R928 B.n705 B.n704 51.3213
R929 B.n698 B.n32 51.3213
R930 B.n698 B.n697 51.3213
R931 B.n697 B.n696 51.3213
R932 B.n696 B.n36 51.3213
R933 B.n690 B.n36 51.3213
R934 B.n690 B.n689 51.3213
R935 B.n689 B.n688 51.3213
R936 B.n688 B.n43 51.3213
R937 B.n682 B.n43 51.3213
R938 B.n682 B.n681 51.3213
R939 B.n680 B.n50 51.3213
R940 B.n674 B.n50 51.3213
R941 B.n674 B.n673 51.3213
R942 B.n673 B.n672 51.3213
R943 B.n672 B.n57 51.3213
R944 B.n666 B.n57 51.3213
R945 B.n666 B.n665 51.3213
R946 B.n572 B.t1 42.2647
R947 B.n32 B.t3 42.2647
R948 B.t0 B.n265 40.7552
R949 B.n721 B.t2 40.7552
R950 B.t9 B.n304 39.2458
R951 B.n681 B.t5 39.2458
R952 B.n108 B.n59 34.8103
R953 B.n662 B.n661 34.8103
R954 B.n521 B.n520 34.8103
R955 B.n514 B.n318 34.8103
R956 B B.n732 18.0485
R957 B.n542 B.t9 12.076
R958 B.t5 B.n680 12.076
R959 B.n109 B.n108 10.6151
R960 B.n112 B.n109 10.6151
R961 B.n113 B.n112 10.6151
R962 B.n116 B.n113 10.6151
R963 B.n117 B.n116 10.6151
R964 B.n120 B.n117 10.6151
R965 B.n121 B.n120 10.6151
R966 B.n124 B.n121 10.6151
R967 B.n125 B.n124 10.6151
R968 B.n128 B.n125 10.6151
R969 B.n129 B.n128 10.6151
R970 B.n132 B.n129 10.6151
R971 B.n133 B.n132 10.6151
R972 B.n136 B.n133 10.6151
R973 B.n137 B.n136 10.6151
R974 B.n140 B.n137 10.6151
R975 B.n141 B.n140 10.6151
R976 B.n144 B.n141 10.6151
R977 B.n145 B.n144 10.6151
R978 B.n148 B.n145 10.6151
R979 B.n149 B.n148 10.6151
R980 B.n152 B.n149 10.6151
R981 B.n153 B.n152 10.6151
R982 B.n156 B.n153 10.6151
R983 B.n157 B.n156 10.6151
R984 B.n160 B.n157 10.6151
R985 B.n161 B.n160 10.6151
R986 B.n164 B.n161 10.6151
R987 B.n165 B.n164 10.6151
R988 B.n168 B.n165 10.6151
R989 B.n169 B.n168 10.6151
R990 B.n172 B.n169 10.6151
R991 B.n173 B.n172 10.6151
R992 B.n177 B.n176 10.6151
R993 B.n180 B.n177 10.6151
R994 B.n181 B.n180 10.6151
R995 B.n184 B.n181 10.6151
R996 B.n185 B.n184 10.6151
R997 B.n188 B.n185 10.6151
R998 B.n189 B.n188 10.6151
R999 B.n192 B.n189 10.6151
R1000 B.n197 B.n194 10.6151
R1001 B.n198 B.n197 10.6151
R1002 B.n201 B.n198 10.6151
R1003 B.n202 B.n201 10.6151
R1004 B.n205 B.n202 10.6151
R1005 B.n206 B.n205 10.6151
R1006 B.n209 B.n206 10.6151
R1007 B.n210 B.n209 10.6151
R1008 B.n213 B.n210 10.6151
R1009 B.n214 B.n213 10.6151
R1010 B.n217 B.n214 10.6151
R1011 B.n218 B.n217 10.6151
R1012 B.n221 B.n218 10.6151
R1013 B.n222 B.n221 10.6151
R1014 B.n225 B.n222 10.6151
R1015 B.n226 B.n225 10.6151
R1016 B.n229 B.n226 10.6151
R1017 B.n230 B.n229 10.6151
R1018 B.n233 B.n230 10.6151
R1019 B.n234 B.n233 10.6151
R1020 B.n237 B.n234 10.6151
R1021 B.n238 B.n237 10.6151
R1022 B.n241 B.n238 10.6151
R1023 B.n242 B.n241 10.6151
R1024 B.n245 B.n242 10.6151
R1025 B.n246 B.n245 10.6151
R1026 B.n249 B.n246 10.6151
R1027 B.n250 B.n249 10.6151
R1028 B.n253 B.n250 10.6151
R1029 B.n254 B.n253 10.6151
R1030 B.n257 B.n254 10.6151
R1031 B.n258 B.n257 10.6151
R1032 B.n662 B.n258 10.6151
R1033 B.n522 B.n521 10.6151
R1034 B.n522 B.n314 10.6151
R1035 B.n532 B.n314 10.6151
R1036 B.n533 B.n532 10.6151
R1037 B.n534 B.n533 10.6151
R1038 B.n534 B.n306 10.6151
R1039 B.n544 B.n306 10.6151
R1040 B.n545 B.n544 10.6151
R1041 B.n546 B.n545 10.6151
R1042 B.n546 B.n298 10.6151
R1043 B.n556 B.n298 10.6151
R1044 B.n557 B.n556 10.6151
R1045 B.n558 B.n557 10.6151
R1046 B.n558 B.n290 10.6151
R1047 B.n568 B.n290 10.6151
R1048 B.n569 B.n568 10.6151
R1049 B.n570 B.n569 10.6151
R1050 B.n570 B.n283 10.6151
R1051 B.n581 B.n283 10.6151
R1052 B.n582 B.n581 10.6151
R1053 B.n583 B.n582 10.6151
R1054 B.n583 B.n275 10.6151
R1055 B.n593 B.n275 10.6151
R1056 B.n594 B.n593 10.6151
R1057 B.n595 B.n594 10.6151
R1058 B.n595 B.n267 10.6151
R1059 B.n605 B.n267 10.6151
R1060 B.n606 B.n605 10.6151
R1061 B.n608 B.n606 10.6151
R1062 B.n608 B.n607 10.6151
R1063 B.n607 B.n259 10.6151
R1064 B.n619 B.n259 10.6151
R1065 B.n620 B.n619 10.6151
R1066 B.n621 B.n620 10.6151
R1067 B.n622 B.n621 10.6151
R1068 B.n624 B.n622 10.6151
R1069 B.n625 B.n624 10.6151
R1070 B.n626 B.n625 10.6151
R1071 B.n627 B.n626 10.6151
R1072 B.n629 B.n627 10.6151
R1073 B.n630 B.n629 10.6151
R1074 B.n631 B.n630 10.6151
R1075 B.n632 B.n631 10.6151
R1076 B.n634 B.n632 10.6151
R1077 B.n635 B.n634 10.6151
R1078 B.n636 B.n635 10.6151
R1079 B.n637 B.n636 10.6151
R1080 B.n639 B.n637 10.6151
R1081 B.n640 B.n639 10.6151
R1082 B.n641 B.n640 10.6151
R1083 B.n642 B.n641 10.6151
R1084 B.n644 B.n642 10.6151
R1085 B.n645 B.n644 10.6151
R1086 B.n646 B.n645 10.6151
R1087 B.n647 B.n646 10.6151
R1088 B.n649 B.n647 10.6151
R1089 B.n650 B.n649 10.6151
R1090 B.n651 B.n650 10.6151
R1091 B.n652 B.n651 10.6151
R1092 B.n654 B.n652 10.6151
R1093 B.n655 B.n654 10.6151
R1094 B.n656 B.n655 10.6151
R1095 B.n657 B.n656 10.6151
R1096 B.n659 B.n657 10.6151
R1097 B.n660 B.n659 10.6151
R1098 B.n661 B.n660 10.6151
R1099 B.n514 B.n513 10.6151
R1100 B.n513 B.n512 10.6151
R1101 B.n512 B.n511 10.6151
R1102 B.n511 B.n509 10.6151
R1103 B.n509 B.n506 10.6151
R1104 B.n506 B.n505 10.6151
R1105 B.n505 B.n502 10.6151
R1106 B.n502 B.n501 10.6151
R1107 B.n501 B.n498 10.6151
R1108 B.n498 B.n497 10.6151
R1109 B.n497 B.n494 10.6151
R1110 B.n494 B.n493 10.6151
R1111 B.n493 B.n490 10.6151
R1112 B.n490 B.n489 10.6151
R1113 B.n489 B.n486 10.6151
R1114 B.n486 B.n485 10.6151
R1115 B.n485 B.n482 10.6151
R1116 B.n482 B.n481 10.6151
R1117 B.n481 B.n478 10.6151
R1118 B.n478 B.n477 10.6151
R1119 B.n477 B.n474 10.6151
R1120 B.n474 B.n473 10.6151
R1121 B.n473 B.n470 10.6151
R1122 B.n470 B.n469 10.6151
R1123 B.n469 B.n466 10.6151
R1124 B.n466 B.n465 10.6151
R1125 B.n465 B.n462 10.6151
R1126 B.n462 B.n461 10.6151
R1127 B.n461 B.n458 10.6151
R1128 B.n458 B.n457 10.6151
R1129 B.n457 B.n454 10.6151
R1130 B.n454 B.n453 10.6151
R1131 B.n453 B.n450 10.6151
R1132 B.n448 B.n445 10.6151
R1133 B.n445 B.n444 10.6151
R1134 B.n444 B.n441 10.6151
R1135 B.n441 B.n440 10.6151
R1136 B.n440 B.n437 10.6151
R1137 B.n437 B.n436 10.6151
R1138 B.n436 B.n433 10.6151
R1139 B.n433 B.n432 10.6151
R1140 B.n429 B.n428 10.6151
R1141 B.n428 B.n425 10.6151
R1142 B.n425 B.n424 10.6151
R1143 B.n424 B.n421 10.6151
R1144 B.n421 B.n420 10.6151
R1145 B.n420 B.n417 10.6151
R1146 B.n417 B.n416 10.6151
R1147 B.n416 B.n413 10.6151
R1148 B.n413 B.n412 10.6151
R1149 B.n412 B.n409 10.6151
R1150 B.n409 B.n408 10.6151
R1151 B.n408 B.n405 10.6151
R1152 B.n405 B.n404 10.6151
R1153 B.n404 B.n401 10.6151
R1154 B.n401 B.n400 10.6151
R1155 B.n400 B.n397 10.6151
R1156 B.n397 B.n396 10.6151
R1157 B.n396 B.n393 10.6151
R1158 B.n393 B.n392 10.6151
R1159 B.n392 B.n389 10.6151
R1160 B.n389 B.n388 10.6151
R1161 B.n388 B.n385 10.6151
R1162 B.n385 B.n384 10.6151
R1163 B.n384 B.n381 10.6151
R1164 B.n381 B.n380 10.6151
R1165 B.n380 B.n377 10.6151
R1166 B.n377 B.n376 10.6151
R1167 B.n376 B.n373 10.6151
R1168 B.n373 B.n372 10.6151
R1169 B.n372 B.n369 10.6151
R1170 B.n369 B.n368 10.6151
R1171 B.n368 B.n322 10.6151
R1172 B.n520 B.n322 10.6151
R1173 B.n526 B.n318 10.6151
R1174 B.n527 B.n526 10.6151
R1175 B.n528 B.n527 10.6151
R1176 B.n528 B.n310 10.6151
R1177 B.n538 B.n310 10.6151
R1178 B.n539 B.n538 10.6151
R1179 B.n540 B.n539 10.6151
R1180 B.n540 B.n302 10.6151
R1181 B.n550 B.n302 10.6151
R1182 B.n551 B.n550 10.6151
R1183 B.n552 B.n551 10.6151
R1184 B.n552 B.n294 10.6151
R1185 B.n562 B.n294 10.6151
R1186 B.n563 B.n562 10.6151
R1187 B.n564 B.n563 10.6151
R1188 B.n564 B.n286 10.6151
R1189 B.n575 B.n286 10.6151
R1190 B.n576 B.n575 10.6151
R1191 B.n577 B.n576 10.6151
R1192 B.n577 B.n279 10.6151
R1193 B.n587 B.n279 10.6151
R1194 B.n588 B.n587 10.6151
R1195 B.n589 B.n588 10.6151
R1196 B.n589 B.n271 10.6151
R1197 B.n599 B.n271 10.6151
R1198 B.n600 B.n599 10.6151
R1199 B.n601 B.n600 10.6151
R1200 B.n601 B.n263 10.6151
R1201 B.n612 B.n263 10.6151
R1202 B.n613 B.n612 10.6151
R1203 B.n614 B.n613 10.6151
R1204 B.n614 B.n0 10.6151
R1205 B.n726 B.n1 10.6151
R1206 B.n726 B.n725 10.6151
R1207 B.n725 B.n724 10.6151
R1208 B.n724 B.n10 10.6151
R1209 B.n718 B.n10 10.6151
R1210 B.n718 B.n717 10.6151
R1211 B.n717 B.n716 10.6151
R1212 B.n716 B.n17 10.6151
R1213 B.n710 B.n17 10.6151
R1214 B.n710 B.n709 10.6151
R1215 B.n709 B.n708 10.6151
R1216 B.n708 B.n24 10.6151
R1217 B.n702 B.n24 10.6151
R1218 B.n702 B.n701 10.6151
R1219 B.n701 B.n700 10.6151
R1220 B.n700 B.n30 10.6151
R1221 B.n694 B.n30 10.6151
R1222 B.n694 B.n693 10.6151
R1223 B.n693 B.n692 10.6151
R1224 B.n692 B.n38 10.6151
R1225 B.n686 B.n38 10.6151
R1226 B.n686 B.n685 10.6151
R1227 B.n685 B.n684 10.6151
R1228 B.n684 B.n45 10.6151
R1229 B.n678 B.n45 10.6151
R1230 B.n678 B.n677 10.6151
R1231 B.n677 B.n676 10.6151
R1232 B.n676 B.n52 10.6151
R1233 B.n670 B.n52 10.6151
R1234 B.n670 B.n669 10.6151
R1235 B.n669 B.n668 10.6151
R1236 B.n668 B.n59 10.6151
R1237 B.n603 B.t0 10.5665
R1238 B.t2 B.n720 10.5665
R1239 B.n579 B.t1 9.0571
R1240 B.n704 B.t3 9.0571
R1241 B.n176 B.n106 6.5566
R1242 B.n193 B.n192 6.5566
R1243 B.n449 B.n448 6.5566
R1244 B.n432 B.n366 6.5566
R1245 B.n173 B.n106 4.05904
R1246 B.n194 B.n193 4.05904
R1247 B.n450 B.n449 4.05904
R1248 B.n429 B.n366 4.05904
R1249 B.n732 B.n0 2.81026
R1250 B.n732 B.n1 2.81026
R1251 VN.n0 VN.t0 124.448
R1252 VN.n1 VN.t3 124.448
R1253 VN.n0 VN.t1 123.688
R1254 VN.n1 VN.t2 123.688
R1255 VN VN.n1 48.764
R1256 VN VN.n0 4.50265
R1257 VDD2.n2 VDD2.n0 103.269
R1258 VDD2.n2 VDD2.n1 64.1655
R1259 VDD2.n1 VDD2.t0 2.12953
R1260 VDD2.n1 VDD2.t1 2.12953
R1261 VDD2.n0 VDD2.t3 2.12953
R1262 VDD2.n0 VDD2.t2 2.12953
R1263 VDD2 VDD2.n2 0.0586897
R1264 VTAIL.n394 VTAIL.n350 289.615
R1265 VTAIL.n44 VTAIL.n0 289.615
R1266 VTAIL.n94 VTAIL.n50 289.615
R1267 VTAIL.n144 VTAIL.n100 289.615
R1268 VTAIL.n344 VTAIL.n300 289.615
R1269 VTAIL.n294 VTAIL.n250 289.615
R1270 VTAIL.n244 VTAIL.n200 289.615
R1271 VTAIL.n194 VTAIL.n150 289.615
R1272 VTAIL.n367 VTAIL.n366 185
R1273 VTAIL.n369 VTAIL.n368 185
R1274 VTAIL.n362 VTAIL.n361 185
R1275 VTAIL.n375 VTAIL.n374 185
R1276 VTAIL.n377 VTAIL.n376 185
R1277 VTAIL.n358 VTAIL.n357 185
R1278 VTAIL.n384 VTAIL.n383 185
R1279 VTAIL.n385 VTAIL.n356 185
R1280 VTAIL.n387 VTAIL.n386 185
R1281 VTAIL.n354 VTAIL.n353 185
R1282 VTAIL.n393 VTAIL.n392 185
R1283 VTAIL.n395 VTAIL.n394 185
R1284 VTAIL.n17 VTAIL.n16 185
R1285 VTAIL.n19 VTAIL.n18 185
R1286 VTAIL.n12 VTAIL.n11 185
R1287 VTAIL.n25 VTAIL.n24 185
R1288 VTAIL.n27 VTAIL.n26 185
R1289 VTAIL.n8 VTAIL.n7 185
R1290 VTAIL.n34 VTAIL.n33 185
R1291 VTAIL.n35 VTAIL.n6 185
R1292 VTAIL.n37 VTAIL.n36 185
R1293 VTAIL.n4 VTAIL.n3 185
R1294 VTAIL.n43 VTAIL.n42 185
R1295 VTAIL.n45 VTAIL.n44 185
R1296 VTAIL.n67 VTAIL.n66 185
R1297 VTAIL.n69 VTAIL.n68 185
R1298 VTAIL.n62 VTAIL.n61 185
R1299 VTAIL.n75 VTAIL.n74 185
R1300 VTAIL.n77 VTAIL.n76 185
R1301 VTAIL.n58 VTAIL.n57 185
R1302 VTAIL.n84 VTAIL.n83 185
R1303 VTAIL.n85 VTAIL.n56 185
R1304 VTAIL.n87 VTAIL.n86 185
R1305 VTAIL.n54 VTAIL.n53 185
R1306 VTAIL.n93 VTAIL.n92 185
R1307 VTAIL.n95 VTAIL.n94 185
R1308 VTAIL.n117 VTAIL.n116 185
R1309 VTAIL.n119 VTAIL.n118 185
R1310 VTAIL.n112 VTAIL.n111 185
R1311 VTAIL.n125 VTAIL.n124 185
R1312 VTAIL.n127 VTAIL.n126 185
R1313 VTAIL.n108 VTAIL.n107 185
R1314 VTAIL.n134 VTAIL.n133 185
R1315 VTAIL.n135 VTAIL.n106 185
R1316 VTAIL.n137 VTAIL.n136 185
R1317 VTAIL.n104 VTAIL.n103 185
R1318 VTAIL.n143 VTAIL.n142 185
R1319 VTAIL.n145 VTAIL.n144 185
R1320 VTAIL.n345 VTAIL.n344 185
R1321 VTAIL.n343 VTAIL.n342 185
R1322 VTAIL.n304 VTAIL.n303 185
R1323 VTAIL.n308 VTAIL.n306 185
R1324 VTAIL.n337 VTAIL.n336 185
R1325 VTAIL.n335 VTAIL.n334 185
R1326 VTAIL.n310 VTAIL.n309 185
R1327 VTAIL.n329 VTAIL.n328 185
R1328 VTAIL.n327 VTAIL.n326 185
R1329 VTAIL.n314 VTAIL.n313 185
R1330 VTAIL.n321 VTAIL.n320 185
R1331 VTAIL.n319 VTAIL.n318 185
R1332 VTAIL.n295 VTAIL.n294 185
R1333 VTAIL.n293 VTAIL.n292 185
R1334 VTAIL.n254 VTAIL.n253 185
R1335 VTAIL.n258 VTAIL.n256 185
R1336 VTAIL.n287 VTAIL.n286 185
R1337 VTAIL.n285 VTAIL.n284 185
R1338 VTAIL.n260 VTAIL.n259 185
R1339 VTAIL.n279 VTAIL.n278 185
R1340 VTAIL.n277 VTAIL.n276 185
R1341 VTAIL.n264 VTAIL.n263 185
R1342 VTAIL.n271 VTAIL.n270 185
R1343 VTAIL.n269 VTAIL.n268 185
R1344 VTAIL.n245 VTAIL.n244 185
R1345 VTAIL.n243 VTAIL.n242 185
R1346 VTAIL.n204 VTAIL.n203 185
R1347 VTAIL.n208 VTAIL.n206 185
R1348 VTAIL.n237 VTAIL.n236 185
R1349 VTAIL.n235 VTAIL.n234 185
R1350 VTAIL.n210 VTAIL.n209 185
R1351 VTAIL.n229 VTAIL.n228 185
R1352 VTAIL.n227 VTAIL.n226 185
R1353 VTAIL.n214 VTAIL.n213 185
R1354 VTAIL.n221 VTAIL.n220 185
R1355 VTAIL.n219 VTAIL.n218 185
R1356 VTAIL.n195 VTAIL.n194 185
R1357 VTAIL.n193 VTAIL.n192 185
R1358 VTAIL.n154 VTAIL.n153 185
R1359 VTAIL.n158 VTAIL.n156 185
R1360 VTAIL.n187 VTAIL.n186 185
R1361 VTAIL.n185 VTAIL.n184 185
R1362 VTAIL.n160 VTAIL.n159 185
R1363 VTAIL.n179 VTAIL.n178 185
R1364 VTAIL.n177 VTAIL.n176 185
R1365 VTAIL.n164 VTAIL.n163 185
R1366 VTAIL.n171 VTAIL.n170 185
R1367 VTAIL.n169 VTAIL.n168 185
R1368 VTAIL.n365 VTAIL.t6 149.524
R1369 VTAIL.n15 VTAIL.t7 149.524
R1370 VTAIL.n65 VTAIL.t2 149.524
R1371 VTAIL.n115 VTAIL.t0 149.524
R1372 VTAIL.n317 VTAIL.t3 149.524
R1373 VTAIL.n267 VTAIL.t1 149.524
R1374 VTAIL.n217 VTAIL.t4 149.524
R1375 VTAIL.n167 VTAIL.t5 149.524
R1376 VTAIL.n368 VTAIL.n367 104.615
R1377 VTAIL.n368 VTAIL.n361 104.615
R1378 VTAIL.n375 VTAIL.n361 104.615
R1379 VTAIL.n376 VTAIL.n375 104.615
R1380 VTAIL.n376 VTAIL.n357 104.615
R1381 VTAIL.n384 VTAIL.n357 104.615
R1382 VTAIL.n385 VTAIL.n384 104.615
R1383 VTAIL.n386 VTAIL.n385 104.615
R1384 VTAIL.n386 VTAIL.n353 104.615
R1385 VTAIL.n393 VTAIL.n353 104.615
R1386 VTAIL.n394 VTAIL.n393 104.615
R1387 VTAIL.n18 VTAIL.n17 104.615
R1388 VTAIL.n18 VTAIL.n11 104.615
R1389 VTAIL.n25 VTAIL.n11 104.615
R1390 VTAIL.n26 VTAIL.n25 104.615
R1391 VTAIL.n26 VTAIL.n7 104.615
R1392 VTAIL.n34 VTAIL.n7 104.615
R1393 VTAIL.n35 VTAIL.n34 104.615
R1394 VTAIL.n36 VTAIL.n35 104.615
R1395 VTAIL.n36 VTAIL.n3 104.615
R1396 VTAIL.n43 VTAIL.n3 104.615
R1397 VTAIL.n44 VTAIL.n43 104.615
R1398 VTAIL.n68 VTAIL.n67 104.615
R1399 VTAIL.n68 VTAIL.n61 104.615
R1400 VTAIL.n75 VTAIL.n61 104.615
R1401 VTAIL.n76 VTAIL.n75 104.615
R1402 VTAIL.n76 VTAIL.n57 104.615
R1403 VTAIL.n84 VTAIL.n57 104.615
R1404 VTAIL.n85 VTAIL.n84 104.615
R1405 VTAIL.n86 VTAIL.n85 104.615
R1406 VTAIL.n86 VTAIL.n53 104.615
R1407 VTAIL.n93 VTAIL.n53 104.615
R1408 VTAIL.n94 VTAIL.n93 104.615
R1409 VTAIL.n118 VTAIL.n117 104.615
R1410 VTAIL.n118 VTAIL.n111 104.615
R1411 VTAIL.n125 VTAIL.n111 104.615
R1412 VTAIL.n126 VTAIL.n125 104.615
R1413 VTAIL.n126 VTAIL.n107 104.615
R1414 VTAIL.n134 VTAIL.n107 104.615
R1415 VTAIL.n135 VTAIL.n134 104.615
R1416 VTAIL.n136 VTAIL.n135 104.615
R1417 VTAIL.n136 VTAIL.n103 104.615
R1418 VTAIL.n143 VTAIL.n103 104.615
R1419 VTAIL.n144 VTAIL.n143 104.615
R1420 VTAIL.n344 VTAIL.n343 104.615
R1421 VTAIL.n343 VTAIL.n303 104.615
R1422 VTAIL.n308 VTAIL.n303 104.615
R1423 VTAIL.n336 VTAIL.n308 104.615
R1424 VTAIL.n336 VTAIL.n335 104.615
R1425 VTAIL.n335 VTAIL.n309 104.615
R1426 VTAIL.n328 VTAIL.n309 104.615
R1427 VTAIL.n328 VTAIL.n327 104.615
R1428 VTAIL.n327 VTAIL.n313 104.615
R1429 VTAIL.n320 VTAIL.n313 104.615
R1430 VTAIL.n320 VTAIL.n319 104.615
R1431 VTAIL.n294 VTAIL.n293 104.615
R1432 VTAIL.n293 VTAIL.n253 104.615
R1433 VTAIL.n258 VTAIL.n253 104.615
R1434 VTAIL.n286 VTAIL.n258 104.615
R1435 VTAIL.n286 VTAIL.n285 104.615
R1436 VTAIL.n285 VTAIL.n259 104.615
R1437 VTAIL.n278 VTAIL.n259 104.615
R1438 VTAIL.n278 VTAIL.n277 104.615
R1439 VTAIL.n277 VTAIL.n263 104.615
R1440 VTAIL.n270 VTAIL.n263 104.615
R1441 VTAIL.n270 VTAIL.n269 104.615
R1442 VTAIL.n244 VTAIL.n243 104.615
R1443 VTAIL.n243 VTAIL.n203 104.615
R1444 VTAIL.n208 VTAIL.n203 104.615
R1445 VTAIL.n236 VTAIL.n208 104.615
R1446 VTAIL.n236 VTAIL.n235 104.615
R1447 VTAIL.n235 VTAIL.n209 104.615
R1448 VTAIL.n228 VTAIL.n209 104.615
R1449 VTAIL.n228 VTAIL.n227 104.615
R1450 VTAIL.n227 VTAIL.n213 104.615
R1451 VTAIL.n220 VTAIL.n213 104.615
R1452 VTAIL.n220 VTAIL.n219 104.615
R1453 VTAIL.n194 VTAIL.n193 104.615
R1454 VTAIL.n193 VTAIL.n153 104.615
R1455 VTAIL.n158 VTAIL.n153 104.615
R1456 VTAIL.n186 VTAIL.n158 104.615
R1457 VTAIL.n186 VTAIL.n185 104.615
R1458 VTAIL.n185 VTAIL.n159 104.615
R1459 VTAIL.n178 VTAIL.n159 104.615
R1460 VTAIL.n178 VTAIL.n177 104.615
R1461 VTAIL.n177 VTAIL.n163 104.615
R1462 VTAIL.n170 VTAIL.n163 104.615
R1463 VTAIL.n170 VTAIL.n169 104.615
R1464 VTAIL.n367 VTAIL.t6 52.3082
R1465 VTAIL.n17 VTAIL.t7 52.3082
R1466 VTAIL.n67 VTAIL.t2 52.3082
R1467 VTAIL.n117 VTAIL.t0 52.3082
R1468 VTAIL.n319 VTAIL.t3 52.3082
R1469 VTAIL.n269 VTAIL.t1 52.3082
R1470 VTAIL.n219 VTAIL.t4 52.3082
R1471 VTAIL.n169 VTAIL.t5 52.3082
R1472 VTAIL.n399 VTAIL.n398 33.349
R1473 VTAIL.n49 VTAIL.n48 33.349
R1474 VTAIL.n99 VTAIL.n98 33.349
R1475 VTAIL.n149 VTAIL.n148 33.349
R1476 VTAIL.n349 VTAIL.n348 33.349
R1477 VTAIL.n299 VTAIL.n298 33.349
R1478 VTAIL.n249 VTAIL.n248 33.349
R1479 VTAIL.n199 VTAIL.n198 33.349
R1480 VTAIL.n399 VTAIL.n349 22.841
R1481 VTAIL.n199 VTAIL.n149 22.841
R1482 VTAIL.n387 VTAIL.n354 13.1884
R1483 VTAIL.n37 VTAIL.n4 13.1884
R1484 VTAIL.n87 VTAIL.n54 13.1884
R1485 VTAIL.n137 VTAIL.n104 13.1884
R1486 VTAIL.n306 VTAIL.n304 13.1884
R1487 VTAIL.n256 VTAIL.n254 13.1884
R1488 VTAIL.n206 VTAIL.n204 13.1884
R1489 VTAIL.n156 VTAIL.n154 13.1884
R1490 VTAIL.n388 VTAIL.n356 12.8005
R1491 VTAIL.n392 VTAIL.n391 12.8005
R1492 VTAIL.n38 VTAIL.n6 12.8005
R1493 VTAIL.n42 VTAIL.n41 12.8005
R1494 VTAIL.n88 VTAIL.n56 12.8005
R1495 VTAIL.n92 VTAIL.n91 12.8005
R1496 VTAIL.n138 VTAIL.n106 12.8005
R1497 VTAIL.n142 VTAIL.n141 12.8005
R1498 VTAIL.n342 VTAIL.n341 12.8005
R1499 VTAIL.n338 VTAIL.n337 12.8005
R1500 VTAIL.n292 VTAIL.n291 12.8005
R1501 VTAIL.n288 VTAIL.n287 12.8005
R1502 VTAIL.n242 VTAIL.n241 12.8005
R1503 VTAIL.n238 VTAIL.n237 12.8005
R1504 VTAIL.n192 VTAIL.n191 12.8005
R1505 VTAIL.n188 VTAIL.n187 12.8005
R1506 VTAIL.n383 VTAIL.n382 12.0247
R1507 VTAIL.n395 VTAIL.n352 12.0247
R1508 VTAIL.n33 VTAIL.n32 12.0247
R1509 VTAIL.n45 VTAIL.n2 12.0247
R1510 VTAIL.n83 VTAIL.n82 12.0247
R1511 VTAIL.n95 VTAIL.n52 12.0247
R1512 VTAIL.n133 VTAIL.n132 12.0247
R1513 VTAIL.n145 VTAIL.n102 12.0247
R1514 VTAIL.n345 VTAIL.n302 12.0247
R1515 VTAIL.n334 VTAIL.n307 12.0247
R1516 VTAIL.n295 VTAIL.n252 12.0247
R1517 VTAIL.n284 VTAIL.n257 12.0247
R1518 VTAIL.n245 VTAIL.n202 12.0247
R1519 VTAIL.n234 VTAIL.n207 12.0247
R1520 VTAIL.n195 VTAIL.n152 12.0247
R1521 VTAIL.n184 VTAIL.n157 12.0247
R1522 VTAIL.n381 VTAIL.n358 11.249
R1523 VTAIL.n396 VTAIL.n350 11.249
R1524 VTAIL.n31 VTAIL.n8 11.249
R1525 VTAIL.n46 VTAIL.n0 11.249
R1526 VTAIL.n81 VTAIL.n58 11.249
R1527 VTAIL.n96 VTAIL.n50 11.249
R1528 VTAIL.n131 VTAIL.n108 11.249
R1529 VTAIL.n146 VTAIL.n100 11.249
R1530 VTAIL.n346 VTAIL.n300 11.249
R1531 VTAIL.n333 VTAIL.n310 11.249
R1532 VTAIL.n296 VTAIL.n250 11.249
R1533 VTAIL.n283 VTAIL.n260 11.249
R1534 VTAIL.n246 VTAIL.n200 11.249
R1535 VTAIL.n233 VTAIL.n210 11.249
R1536 VTAIL.n196 VTAIL.n150 11.249
R1537 VTAIL.n183 VTAIL.n160 11.249
R1538 VTAIL.n378 VTAIL.n377 10.4732
R1539 VTAIL.n28 VTAIL.n27 10.4732
R1540 VTAIL.n78 VTAIL.n77 10.4732
R1541 VTAIL.n128 VTAIL.n127 10.4732
R1542 VTAIL.n330 VTAIL.n329 10.4732
R1543 VTAIL.n280 VTAIL.n279 10.4732
R1544 VTAIL.n230 VTAIL.n229 10.4732
R1545 VTAIL.n180 VTAIL.n179 10.4732
R1546 VTAIL.n366 VTAIL.n365 10.2747
R1547 VTAIL.n16 VTAIL.n15 10.2747
R1548 VTAIL.n66 VTAIL.n65 10.2747
R1549 VTAIL.n116 VTAIL.n115 10.2747
R1550 VTAIL.n318 VTAIL.n317 10.2747
R1551 VTAIL.n268 VTAIL.n267 10.2747
R1552 VTAIL.n218 VTAIL.n217 10.2747
R1553 VTAIL.n168 VTAIL.n167 10.2747
R1554 VTAIL.n374 VTAIL.n360 9.69747
R1555 VTAIL.n24 VTAIL.n10 9.69747
R1556 VTAIL.n74 VTAIL.n60 9.69747
R1557 VTAIL.n124 VTAIL.n110 9.69747
R1558 VTAIL.n326 VTAIL.n312 9.69747
R1559 VTAIL.n276 VTAIL.n262 9.69747
R1560 VTAIL.n226 VTAIL.n212 9.69747
R1561 VTAIL.n176 VTAIL.n162 9.69747
R1562 VTAIL.n398 VTAIL.n397 9.45567
R1563 VTAIL.n48 VTAIL.n47 9.45567
R1564 VTAIL.n98 VTAIL.n97 9.45567
R1565 VTAIL.n148 VTAIL.n147 9.45567
R1566 VTAIL.n348 VTAIL.n347 9.45567
R1567 VTAIL.n298 VTAIL.n297 9.45567
R1568 VTAIL.n248 VTAIL.n247 9.45567
R1569 VTAIL.n198 VTAIL.n197 9.45567
R1570 VTAIL.n397 VTAIL.n396 9.3005
R1571 VTAIL.n352 VTAIL.n351 9.3005
R1572 VTAIL.n391 VTAIL.n390 9.3005
R1573 VTAIL.n364 VTAIL.n363 9.3005
R1574 VTAIL.n371 VTAIL.n370 9.3005
R1575 VTAIL.n373 VTAIL.n372 9.3005
R1576 VTAIL.n360 VTAIL.n359 9.3005
R1577 VTAIL.n379 VTAIL.n378 9.3005
R1578 VTAIL.n381 VTAIL.n380 9.3005
R1579 VTAIL.n382 VTAIL.n355 9.3005
R1580 VTAIL.n389 VTAIL.n388 9.3005
R1581 VTAIL.n47 VTAIL.n46 9.3005
R1582 VTAIL.n2 VTAIL.n1 9.3005
R1583 VTAIL.n41 VTAIL.n40 9.3005
R1584 VTAIL.n14 VTAIL.n13 9.3005
R1585 VTAIL.n21 VTAIL.n20 9.3005
R1586 VTAIL.n23 VTAIL.n22 9.3005
R1587 VTAIL.n10 VTAIL.n9 9.3005
R1588 VTAIL.n29 VTAIL.n28 9.3005
R1589 VTAIL.n31 VTAIL.n30 9.3005
R1590 VTAIL.n32 VTAIL.n5 9.3005
R1591 VTAIL.n39 VTAIL.n38 9.3005
R1592 VTAIL.n97 VTAIL.n96 9.3005
R1593 VTAIL.n52 VTAIL.n51 9.3005
R1594 VTAIL.n91 VTAIL.n90 9.3005
R1595 VTAIL.n64 VTAIL.n63 9.3005
R1596 VTAIL.n71 VTAIL.n70 9.3005
R1597 VTAIL.n73 VTAIL.n72 9.3005
R1598 VTAIL.n60 VTAIL.n59 9.3005
R1599 VTAIL.n79 VTAIL.n78 9.3005
R1600 VTAIL.n81 VTAIL.n80 9.3005
R1601 VTAIL.n82 VTAIL.n55 9.3005
R1602 VTAIL.n89 VTAIL.n88 9.3005
R1603 VTAIL.n147 VTAIL.n146 9.3005
R1604 VTAIL.n102 VTAIL.n101 9.3005
R1605 VTAIL.n141 VTAIL.n140 9.3005
R1606 VTAIL.n114 VTAIL.n113 9.3005
R1607 VTAIL.n121 VTAIL.n120 9.3005
R1608 VTAIL.n123 VTAIL.n122 9.3005
R1609 VTAIL.n110 VTAIL.n109 9.3005
R1610 VTAIL.n129 VTAIL.n128 9.3005
R1611 VTAIL.n131 VTAIL.n130 9.3005
R1612 VTAIL.n132 VTAIL.n105 9.3005
R1613 VTAIL.n139 VTAIL.n138 9.3005
R1614 VTAIL.n316 VTAIL.n315 9.3005
R1615 VTAIL.n323 VTAIL.n322 9.3005
R1616 VTAIL.n325 VTAIL.n324 9.3005
R1617 VTAIL.n312 VTAIL.n311 9.3005
R1618 VTAIL.n331 VTAIL.n330 9.3005
R1619 VTAIL.n333 VTAIL.n332 9.3005
R1620 VTAIL.n307 VTAIL.n305 9.3005
R1621 VTAIL.n339 VTAIL.n338 9.3005
R1622 VTAIL.n347 VTAIL.n346 9.3005
R1623 VTAIL.n302 VTAIL.n301 9.3005
R1624 VTAIL.n341 VTAIL.n340 9.3005
R1625 VTAIL.n266 VTAIL.n265 9.3005
R1626 VTAIL.n273 VTAIL.n272 9.3005
R1627 VTAIL.n275 VTAIL.n274 9.3005
R1628 VTAIL.n262 VTAIL.n261 9.3005
R1629 VTAIL.n281 VTAIL.n280 9.3005
R1630 VTAIL.n283 VTAIL.n282 9.3005
R1631 VTAIL.n257 VTAIL.n255 9.3005
R1632 VTAIL.n289 VTAIL.n288 9.3005
R1633 VTAIL.n297 VTAIL.n296 9.3005
R1634 VTAIL.n252 VTAIL.n251 9.3005
R1635 VTAIL.n291 VTAIL.n290 9.3005
R1636 VTAIL.n216 VTAIL.n215 9.3005
R1637 VTAIL.n223 VTAIL.n222 9.3005
R1638 VTAIL.n225 VTAIL.n224 9.3005
R1639 VTAIL.n212 VTAIL.n211 9.3005
R1640 VTAIL.n231 VTAIL.n230 9.3005
R1641 VTAIL.n233 VTAIL.n232 9.3005
R1642 VTAIL.n207 VTAIL.n205 9.3005
R1643 VTAIL.n239 VTAIL.n238 9.3005
R1644 VTAIL.n247 VTAIL.n246 9.3005
R1645 VTAIL.n202 VTAIL.n201 9.3005
R1646 VTAIL.n241 VTAIL.n240 9.3005
R1647 VTAIL.n166 VTAIL.n165 9.3005
R1648 VTAIL.n173 VTAIL.n172 9.3005
R1649 VTAIL.n175 VTAIL.n174 9.3005
R1650 VTAIL.n162 VTAIL.n161 9.3005
R1651 VTAIL.n181 VTAIL.n180 9.3005
R1652 VTAIL.n183 VTAIL.n182 9.3005
R1653 VTAIL.n157 VTAIL.n155 9.3005
R1654 VTAIL.n189 VTAIL.n188 9.3005
R1655 VTAIL.n197 VTAIL.n196 9.3005
R1656 VTAIL.n152 VTAIL.n151 9.3005
R1657 VTAIL.n191 VTAIL.n190 9.3005
R1658 VTAIL.n373 VTAIL.n362 8.92171
R1659 VTAIL.n23 VTAIL.n12 8.92171
R1660 VTAIL.n73 VTAIL.n62 8.92171
R1661 VTAIL.n123 VTAIL.n112 8.92171
R1662 VTAIL.n325 VTAIL.n314 8.92171
R1663 VTAIL.n275 VTAIL.n264 8.92171
R1664 VTAIL.n225 VTAIL.n214 8.92171
R1665 VTAIL.n175 VTAIL.n164 8.92171
R1666 VTAIL.n370 VTAIL.n369 8.14595
R1667 VTAIL.n20 VTAIL.n19 8.14595
R1668 VTAIL.n70 VTAIL.n69 8.14595
R1669 VTAIL.n120 VTAIL.n119 8.14595
R1670 VTAIL.n322 VTAIL.n321 8.14595
R1671 VTAIL.n272 VTAIL.n271 8.14595
R1672 VTAIL.n222 VTAIL.n221 8.14595
R1673 VTAIL.n172 VTAIL.n171 8.14595
R1674 VTAIL.n366 VTAIL.n364 7.3702
R1675 VTAIL.n16 VTAIL.n14 7.3702
R1676 VTAIL.n66 VTAIL.n64 7.3702
R1677 VTAIL.n116 VTAIL.n114 7.3702
R1678 VTAIL.n318 VTAIL.n316 7.3702
R1679 VTAIL.n268 VTAIL.n266 7.3702
R1680 VTAIL.n218 VTAIL.n216 7.3702
R1681 VTAIL.n168 VTAIL.n166 7.3702
R1682 VTAIL.n369 VTAIL.n364 5.81868
R1683 VTAIL.n19 VTAIL.n14 5.81868
R1684 VTAIL.n69 VTAIL.n64 5.81868
R1685 VTAIL.n119 VTAIL.n114 5.81868
R1686 VTAIL.n321 VTAIL.n316 5.81868
R1687 VTAIL.n271 VTAIL.n266 5.81868
R1688 VTAIL.n221 VTAIL.n216 5.81868
R1689 VTAIL.n171 VTAIL.n166 5.81868
R1690 VTAIL.n370 VTAIL.n362 5.04292
R1691 VTAIL.n20 VTAIL.n12 5.04292
R1692 VTAIL.n70 VTAIL.n62 5.04292
R1693 VTAIL.n120 VTAIL.n112 5.04292
R1694 VTAIL.n322 VTAIL.n314 5.04292
R1695 VTAIL.n272 VTAIL.n264 5.04292
R1696 VTAIL.n222 VTAIL.n214 5.04292
R1697 VTAIL.n172 VTAIL.n164 5.04292
R1698 VTAIL.n374 VTAIL.n373 4.26717
R1699 VTAIL.n24 VTAIL.n23 4.26717
R1700 VTAIL.n74 VTAIL.n73 4.26717
R1701 VTAIL.n124 VTAIL.n123 4.26717
R1702 VTAIL.n326 VTAIL.n325 4.26717
R1703 VTAIL.n276 VTAIL.n275 4.26717
R1704 VTAIL.n226 VTAIL.n225 4.26717
R1705 VTAIL.n176 VTAIL.n175 4.26717
R1706 VTAIL.n377 VTAIL.n360 3.49141
R1707 VTAIL.n27 VTAIL.n10 3.49141
R1708 VTAIL.n77 VTAIL.n60 3.49141
R1709 VTAIL.n127 VTAIL.n110 3.49141
R1710 VTAIL.n329 VTAIL.n312 3.49141
R1711 VTAIL.n279 VTAIL.n262 3.49141
R1712 VTAIL.n229 VTAIL.n212 3.49141
R1713 VTAIL.n179 VTAIL.n162 3.49141
R1714 VTAIL.n365 VTAIL.n363 2.84303
R1715 VTAIL.n15 VTAIL.n13 2.84303
R1716 VTAIL.n65 VTAIL.n63 2.84303
R1717 VTAIL.n115 VTAIL.n113 2.84303
R1718 VTAIL.n317 VTAIL.n315 2.84303
R1719 VTAIL.n267 VTAIL.n265 2.84303
R1720 VTAIL.n217 VTAIL.n215 2.84303
R1721 VTAIL.n167 VTAIL.n165 2.84303
R1722 VTAIL.n378 VTAIL.n358 2.71565
R1723 VTAIL.n398 VTAIL.n350 2.71565
R1724 VTAIL.n28 VTAIL.n8 2.71565
R1725 VTAIL.n48 VTAIL.n0 2.71565
R1726 VTAIL.n78 VTAIL.n58 2.71565
R1727 VTAIL.n98 VTAIL.n50 2.71565
R1728 VTAIL.n128 VTAIL.n108 2.71565
R1729 VTAIL.n148 VTAIL.n100 2.71565
R1730 VTAIL.n348 VTAIL.n300 2.71565
R1731 VTAIL.n330 VTAIL.n310 2.71565
R1732 VTAIL.n298 VTAIL.n250 2.71565
R1733 VTAIL.n280 VTAIL.n260 2.71565
R1734 VTAIL.n248 VTAIL.n200 2.71565
R1735 VTAIL.n230 VTAIL.n210 2.71565
R1736 VTAIL.n198 VTAIL.n150 2.71565
R1737 VTAIL.n180 VTAIL.n160 2.71565
R1738 VTAIL.n249 VTAIL.n199 2.4574
R1739 VTAIL.n349 VTAIL.n299 2.4574
R1740 VTAIL.n149 VTAIL.n99 2.4574
R1741 VTAIL.n383 VTAIL.n381 1.93989
R1742 VTAIL.n396 VTAIL.n395 1.93989
R1743 VTAIL.n33 VTAIL.n31 1.93989
R1744 VTAIL.n46 VTAIL.n45 1.93989
R1745 VTAIL.n83 VTAIL.n81 1.93989
R1746 VTAIL.n96 VTAIL.n95 1.93989
R1747 VTAIL.n133 VTAIL.n131 1.93989
R1748 VTAIL.n146 VTAIL.n145 1.93989
R1749 VTAIL.n346 VTAIL.n345 1.93989
R1750 VTAIL.n334 VTAIL.n333 1.93989
R1751 VTAIL.n296 VTAIL.n295 1.93989
R1752 VTAIL.n284 VTAIL.n283 1.93989
R1753 VTAIL.n246 VTAIL.n245 1.93989
R1754 VTAIL.n234 VTAIL.n233 1.93989
R1755 VTAIL.n196 VTAIL.n195 1.93989
R1756 VTAIL.n184 VTAIL.n183 1.93989
R1757 VTAIL VTAIL.n49 1.28714
R1758 VTAIL VTAIL.n399 1.17076
R1759 VTAIL.n382 VTAIL.n356 1.16414
R1760 VTAIL.n392 VTAIL.n352 1.16414
R1761 VTAIL.n32 VTAIL.n6 1.16414
R1762 VTAIL.n42 VTAIL.n2 1.16414
R1763 VTAIL.n82 VTAIL.n56 1.16414
R1764 VTAIL.n92 VTAIL.n52 1.16414
R1765 VTAIL.n132 VTAIL.n106 1.16414
R1766 VTAIL.n142 VTAIL.n102 1.16414
R1767 VTAIL.n342 VTAIL.n302 1.16414
R1768 VTAIL.n337 VTAIL.n307 1.16414
R1769 VTAIL.n292 VTAIL.n252 1.16414
R1770 VTAIL.n287 VTAIL.n257 1.16414
R1771 VTAIL.n242 VTAIL.n202 1.16414
R1772 VTAIL.n237 VTAIL.n207 1.16414
R1773 VTAIL.n192 VTAIL.n152 1.16414
R1774 VTAIL.n187 VTAIL.n157 1.16414
R1775 VTAIL.n299 VTAIL.n249 0.470328
R1776 VTAIL.n99 VTAIL.n49 0.470328
R1777 VTAIL.n388 VTAIL.n387 0.388379
R1778 VTAIL.n391 VTAIL.n354 0.388379
R1779 VTAIL.n38 VTAIL.n37 0.388379
R1780 VTAIL.n41 VTAIL.n4 0.388379
R1781 VTAIL.n88 VTAIL.n87 0.388379
R1782 VTAIL.n91 VTAIL.n54 0.388379
R1783 VTAIL.n138 VTAIL.n137 0.388379
R1784 VTAIL.n141 VTAIL.n104 0.388379
R1785 VTAIL.n341 VTAIL.n304 0.388379
R1786 VTAIL.n338 VTAIL.n306 0.388379
R1787 VTAIL.n291 VTAIL.n254 0.388379
R1788 VTAIL.n288 VTAIL.n256 0.388379
R1789 VTAIL.n241 VTAIL.n204 0.388379
R1790 VTAIL.n238 VTAIL.n206 0.388379
R1791 VTAIL.n191 VTAIL.n154 0.388379
R1792 VTAIL.n188 VTAIL.n156 0.388379
R1793 VTAIL.n371 VTAIL.n363 0.155672
R1794 VTAIL.n372 VTAIL.n371 0.155672
R1795 VTAIL.n372 VTAIL.n359 0.155672
R1796 VTAIL.n379 VTAIL.n359 0.155672
R1797 VTAIL.n380 VTAIL.n379 0.155672
R1798 VTAIL.n380 VTAIL.n355 0.155672
R1799 VTAIL.n389 VTAIL.n355 0.155672
R1800 VTAIL.n390 VTAIL.n389 0.155672
R1801 VTAIL.n390 VTAIL.n351 0.155672
R1802 VTAIL.n397 VTAIL.n351 0.155672
R1803 VTAIL.n21 VTAIL.n13 0.155672
R1804 VTAIL.n22 VTAIL.n21 0.155672
R1805 VTAIL.n22 VTAIL.n9 0.155672
R1806 VTAIL.n29 VTAIL.n9 0.155672
R1807 VTAIL.n30 VTAIL.n29 0.155672
R1808 VTAIL.n30 VTAIL.n5 0.155672
R1809 VTAIL.n39 VTAIL.n5 0.155672
R1810 VTAIL.n40 VTAIL.n39 0.155672
R1811 VTAIL.n40 VTAIL.n1 0.155672
R1812 VTAIL.n47 VTAIL.n1 0.155672
R1813 VTAIL.n71 VTAIL.n63 0.155672
R1814 VTAIL.n72 VTAIL.n71 0.155672
R1815 VTAIL.n72 VTAIL.n59 0.155672
R1816 VTAIL.n79 VTAIL.n59 0.155672
R1817 VTAIL.n80 VTAIL.n79 0.155672
R1818 VTAIL.n80 VTAIL.n55 0.155672
R1819 VTAIL.n89 VTAIL.n55 0.155672
R1820 VTAIL.n90 VTAIL.n89 0.155672
R1821 VTAIL.n90 VTAIL.n51 0.155672
R1822 VTAIL.n97 VTAIL.n51 0.155672
R1823 VTAIL.n121 VTAIL.n113 0.155672
R1824 VTAIL.n122 VTAIL.n121 0.155672
R1825 VTAIL.n122 VTAIL.n109 0.155672
R1826 VTAIL.n129 VTAIL.n109 0.155672
R1827 VTAIL.n130 VTAIL.n129 0.155672
R1828 VTAIL.n130 VTAIL.n105 0.155672
R1829 VTAIL.n139 VTAIL.n105 0.155672
R1830 VTAIL.n140 VTAIL.n139 0.155672
R1831 VTAIL.n140 VTAIL.n101 0.155672
R1832 VTAIL.n147 VTAIL.n101 0.155672
R1833 VTAIL.n347 VTAIL.n301 0.155672
R1834 VTAIL.n340 VTAIL.n301 0.155672
R1835 VTAIL.n340 VTAIL.n339 0.155672
R1836 VTAIL.n339 VTAIL.n305 0.155672
R1837 VTAIL.n332 VTAIL.n305 0.155672
R1838 VTAIL.n332 VTAIL.n331 0.155672
R1839 VTAIL.n331 VTAIL.n311 0.155672
R1840 VTAIL.n324 VTAIL.n311 0.155672
R1841 VTAIL.n324 VTAIL.n323 0.155672
R1842 VTAIL.n323 VTAIL.n315 0.155672
R1843 VTAIL.n297 VTAIL.n251 0.155672
R1844 VTAIL.n290 VTAIL.n251 0.155672
R1845 VTAIL.n290 VTAIL.n289 0.155672
R1846 VTAIL.n289 VTAIL.n255 0.155672
R1847 VTAIL.n282 VTAIL.n255 0.155672
R1848 VTAIL.n282 VTAIL.n281 0.155672
R1849 VTAIL.n281 VTAIL.n261 0.155672
R1850 VTAIL.n274 VTAIL.n261 0.155672
R1851 VTAIL.n274 VTAIL.n273 0.155672
R1852 VTAIL.n273 VTAIL.n265 0.155672
R1853 VTAIL.n247 VTAIL.n201 0.155672
R1854 VTAIL.n240 VTAIL.n201 0.155672
R1855 VTAIL.n240 VTAIL.n239 0.155672
R1856 VTAIL.n239 VTAIL.n205 0.155672
R1857 VTAIL.n232 VTAIL.n205 0.155672
R1858 VTAIL.n232 VTAIL.n231 0.155672
R1859 VTAIL.n231 VTAIL.n211 0.155672
R1860 VTAIL.n224 VTAIL.n211 0.155672
R1861 VTAIL.n224 VTAIL.n223 0.155672
R1862 VTAIL.n223 VTAIL.n215 0.155672
R1863 VTAIL.n197 VTAIL.n151 0.155672
R1864 VTAIL.n190 VTAIL.n151 0.155672
R1865 VTAIL.n190 VTAIL.n189 0.155672
R1866 VTAIL.n189 VTAIL.n155 0.155672
R1867 VTAIL.n182 VTAIL.n155 0.155672
R1868 VTAIL.n182 VTAIL.n181 0.155672
R1869 VTAIL.n181 VTAIL.n161 0.155672
R1870 VTAIL.n174 VTAIL.n161 0.155672
R1871 VTAIL.n174 VTAIL.n173 0.155672
R1872 VTAIL.n173 VTAIL.n165 0.155672
R1873 VP.n14 VP.n0 161.3
R1874 VP.n13 VP.n12 161.3
R1875 VP.n11 VP.n1 161.3
R1876 VP.n10 VP.n9 161.3
R1877 VP.n8 VP.n2 161.3
R1878 VP.n7 VP.n6 161.3
R1879 VP.n4 VP.t2 124.448
R1880 VP.n4 VP.t0 123.688
R1881 VP.n5 VP.n3 102.085
R1882 VP.n16 VP.n15 102.085
R1883 VP.n3 VP.t3 88.941
R1884 VP.n15 VP.t1 88.941
R1885 VP.n9 VP.n1 56.4773
R1886 VP.n5 VP.n4 48.4851
R1887 VP.n8 VP.n7 24.3439
R1888 VP.n9 VP.n8 24.3439
R1889 VP.n13 VP.n1 24.3439
R1890 VP.n14 VP.n13 24.3439
R1891 VP.n7 VP.n3 8.5207
R1892 VP.n15 VP.n14 8.5207
R1893 VP.n6 VP.n5 0.278398
R1894 VP.n16 VP.n0 0.278398
R1895 VP.n6 VP.n2 0.189894
R1896 VP.n10 VP.n2 0.189894
R1897 VP.n11 VP.n10 0.189894
R1898 VP.n12 VP.n11 0.189894
R1899 VP.n12 VP.n0 0.189894
R1900 VP VP.n16 0.153422
R1901 VDD1 VDD1.n1 103.793
R1902 VDD1 VDD1.n0 64.2237
R1903 VDD1.n0 VDD1.t1 2.12953
R1904 VDD1.n0 VDD1.t3 2.12953
R1905 VDD1.n1 VDD1.t0 2.12953
R1906 VDD1.n1 VDD1.t2 2.12953
C0 VP VN 5.6382f
C1 VN VDD1 0.148728f
C2 VP VTAIL 3.76174f
C3 VDD1 VTAIL 4.74569f
C4 VP VDD1 3.96703f
C5 VDD2 VN 3.72746f
C6 VDD2 VTAIL 4.79936f
C7 VN VTAIL 3.74763f
C8 VP VDD2 0.389015f
C9 VDD2 VDD1 1.01457f
C10 VDD2 B 3.5066f
C11 VDD1 B 7.34513f
C12 VTAIL B 8.41236f
C13 VN B 10.31276f
C14 VP B 8.583734f
C15 VDD1.t1 B 0.200467f
C16 VDD1.t3 B 0.200467f
C17 VDD1.n0 B 1.75727f
C18 VDD1.t0 B 0.200467f
C19 VDD1.t2 B 0.200467f
C20 VDD1.n1 B 2.35347f
C21 VP.n0 B 0.036234f
C22 VP.t1 B 1.74027f
C23 VP.n1 B 0.040293f
C24 VP.n2 B 0.027482f
C25 VP.t3 B 1.74027f
C26 VP.n3 B 0.71465f
C27 VP.t0 B 1.96413f
C28 VP.t2 B 1.96893f
C29 VP.n4 B 2.62062f
C30 VP.n5 B 1.42289f
C31 VP.n6 B 0.036234f
C32 VP.n7 B 0.034956f
C33 VP.n8 B 0.051476f
C34 VP.n9 B 0.040293f
C35 VP.n10 B 0.027482f
C36 VP.n11 B 0.027482f
C37 VP.n12 B 0.027482f
C38 VP.n13 B 0.051476f
C39 VP.n14 B 0.034956f
C40 VP.n15 B 0.71465f
C41 VP.n16 B 0.044998f
C42 VTAIL.n0 B 0.023025f
C43 VTAIL.n1 B 0.017207f
C44 VTAIL.n2 B 0.009246f
C45 VTAIL.n3 B 0.021855f
C46 VTAIL.n4 B 0.009518f
C47 VTAIL.n5 B 0.017207f
C48 VTAIL.n6 B 0.00979f
C49 VTAIL.n7 B 0.021855f
C50 VTAIL.n8 B 0.00979f
C51 VTAIL.n9 B 0.017207f
C52 VTAIL.n10 B 0.009246f
C53 VTAIL.n11 B 0.021855f
C54 VTAIL.n12 B 0.00979f
C55 VTAIL.n13 B 0.661408f
C56 VTAIL.n14 B 0.009246f
C57 VTAIL.t7 B 0.036664f
C58 VTAIL.n15 B 0.106228f
C59 VTAIL.n16 B 0.01545f
C60 VTAIL.n17 B 0.016391f
C61 VTAIL.n18 B 0.021855f
C62 VTAIL.n19 B 0.00979f
C63 VTAIL.n20 B 0.009246f
C64 VTAIL.n21 B 0.017207f
C65 VTAIL.n22 B 0.017207f
C66 VTAIL.n23 B 0.009246f
C67 VTAIL.n24 B 0.00979f
C68 VTAIL.n25 B 0.021855f
C69 VTAIL.n26 B 0.021855f
C70 VTAIL.n27 B 0.00979f
C71 VTAIL.n28 B 0.009246f
C72 VTAIL.n29 B 0.017207f
C73 VTAIL.n30 B 0.017207f
C74 VTAIL.n31 B 0.009246f
C75 VTAIL.n32 B 0.009246f
C76 VTAIL.n33 B 0.00979f
C77 VTAIL.n34 B 0.021855f
C78 VTAIL.n35 B 0.021855f
C79 VTAIL.n36 B 0.021855f
C80 VTAIL.n37 B 0.009518f
C81 VTAIL.n38 B 0.009246f
C82 VTAIL.n39 B 0.017207f
C83 VTAIL.n40 B 0.017207f
C84 VTAIL.n41 B 0.009246f
C85 VTAIL.n42 B 0.00979f
C86 VTAIL.n43 B 0.021855f
C87 VTAIL.n44 B 0.045259f
C88 VTAIL.n45 B 0.00979f
C89 VTAIL.n46 B 0.009246f
C90 VTAIL.n47 B 0.041183f
C91 VTAIL.n48 B 0.025156f
C92 VTAIL.n49 B 0.112879f
C93 VTAIL.n50 B 0.023025f
C94 VTAIL.n51 B 0.017207f
C95 VTAIL.n52 B 0.009246f
C96 VTAIL.n53 B 0.021855f
C97 VTAIL.n54 B 0.009518f
C98 VTAIL.n55 B 0.017207f
C99 VTAIL.n56 B 0.00979f
C100 VTAIL.n57 B 0.021855f
C101 VTAIL.n58 B 0.00979f
C102 VTAIL.n59 B 0.017207f
C103 VTAIL.n60 B 0.009246f
C104 VTAIL.n61 B 0.021855f
C105 VTAIL.n62 B 0.00979f
C106 VTAIL.n63 B 0.661408f
C107 VTAIL.n64 B 0.009246f
C108 VTAIL.t2 B 0.036664f
C109 VTAIL.n65 B 0.106228f
C110 VTAIL.n66 B 0.01545f
C111 VTAIL.n67 B 0.016391f
C112 VTAIL.n68 B 0.021855f
C113 VTAIL.n69 B 0.00979f
C114 VTAIL.n70 B 0.009246f
C115 VTAIL.n71 B 0.017207f
C116 VTAIL.n72 B 0.017207f
C117 VTAIL.n73 B 0.009246f
C118 VTAIL.n74 B 0.00979f
C119 VTAIL.n75 B 0.021855f
C120 VTAIL.n76 B 0.021855f
C121 VTAIL.n77 B 0.00979f
C122 VTAIL.n78 B 0.009246f
C123 VTAIL.n79 B 0.017207f
C124 VTAIL.n80 B 0.017207f
C125 VTAIL.n81 B 0.009246f
C126 VTAIL.n82 B 0.009246f
C127 VTAIL.n83 B 0.00979f
C128 VTAIL.n84 B 0.021855f
C129 VTAIL.n85 B 0.021855f
C130 VTAIL.n86 B 0.021855f
C131 VTAIL.n87 B 0.009518f
C132 VTAIL.n88 B 0.009246f
C133 VTAIL.n89 B 0.017207f
C134 VTAIL.n90 B 0.017207f
C135 VTAIL.n91 B 0.009246f
C136 VTAIL.n92 B 0.00979f
C137 VTAIL.n93 B 0.021855f
C138 VTAIL.n94 B 0.045259f
C139 VTAIL.n95 B 0.00979f
C140 VTAIL.n96 B 0.009246f
C141 VTAIL.n97 B 0.041183f
C142 VTAIL.n98 B 0.025156f
C143 VTAIL.n99 B 0.177763f
C144 VTAIL.n100 B 0.023025f
C145 VTAIL.n101 B 0.017207f
C146 VTAIL.n102 B 0.009246f
C147 VTAIL.n103 B 0.021855f
C148 VTAIL.n104 B 0.009518f
C149 VTAIL.n105 B 0.017207f
C150 VTAIL.n106 B 0.00979f
C151 VTAIL.n107 B 0.021855f
C152 VTAIL.n108 B 0.00979f
C153 VTAIL.n109 B 0.017207f
C154 VTAIL.n110 B 0.009246f
C155 VTAIL.n111 B 0.021855f
C156 VTAIL.n112 B 0.00979f
C157 VTAIL.n113 B 0.661408f
C158 VTAIL.n114 B 0.009246f
C159 VTAIL.t0 B 0.036664f
C160 VTAIL.n115 B 0.106228f
C161 VTAIL.n116 B 0.01545f
C162 VTAIL.n117 B 0.016391f
C163 VTAIL.n118 B 0.021855f
C164 VTAIL.n119 B 0.00979f
C165 VTAIL.n120 B 0.009246f
C166 VTAIL.n121 B 0.017207f
C167 VTAIL.n122 B 0.017207f
C168 VTAIL.n123 B 0.009246f
C169 VTAIL.n124 B 0.00979f
C170 VTAIL.n125 B 0.021855f
C171 VTAIL.n126 B 0.021855f
C172 VTAIL.n127 B 0.00979f
C173 VTAIL.n128 B 0.009246f
C174 VTAIL.n129 B 0.017207f
C175 VTAIL.n130 B 0.017207f
C176 VTAIL.n131 B 0.009246f
C177 VTAIL.n132 B 0.009246f
C178 VTAIL.n133 B 0.00979f
C179 VTAIL.n134 B 0.021855f
C180 VTAIL.n135 B 0.021855f
C181 VTAIL.n136 B 0.021855f
C182 VTAIL.n137 B 0.009518f
C183 VTAIL.n138 B 0.009246f
C184 VTAIL.n139 B 0.017207f
C185 VTAIL.n140 B 0.017207f
C186 VTAIL.n141 B 0.009246f
C187 VTAIL.n142 B 0.00979f
C188 VTAIL.n143 B 0.021855f
C189 VTAIL.n144 B 0.045259f
C190 VTAIL.n145 B 0.00979f
C191 VTAIL.n146 B 0.009246f
C192 VTAIL.n147 B 0.041183f
C193 VTAIL.n148 B 0.025156f
C194 VTAIL.n149 B 0.966181f
C195 VTAIL.n150 B 0.023025f
C196 VTAIL.n151 B 0.017207f
C197 VTAIL.n152 B 0.009246f
C198 VTAIL.n153 B 0.021855f
C199 VTAIL.n154 B 0.009518f
C200 VTAIL.n155 B 0.017207f
C201 VTAIL.n156 B 0.009518f
C202 VTAIL.n157 B 0.009246f
C203 VTAIL.n158 B 0.021855f
C204 VTAIL.n159 B 0.021855f
C205 VTAIL.n160 B 0.00979f
C206 VTAIL.n161 B 0.017207f
C207 VTAIL.n162 B 0.009246f
C208 VTAIL.n163 B 0.021855f
C209 VTAIL.n164 B 0.00979f
C210 VTAIL.n165 B 0.661408f
C211 VTAIL.n166 B 0.009246f
C212 VTAIL.t5 B 0.036664f
C213 VTAIL.n167 B 0.106228f
C214 VTAIL.n168 B 0.01545f
C215 VTAIL.n169 B 0.016391f
C216 VTAIL.n170 B 0.021855f
C217 VTAIL.n171 B 0.00979f
C218 VTAIL.n172 B 0.009246f
C219 VTAIL.n173 B 0.017207f
C220 VTAIL.n174 B 0.017207f
C221 VTAIL.n175 B 0.009246f
C222 VTAIL.n176 B 0.00979f
C223 VTAIL.n177 B 0.021855f
C224 VTAIL.n178 B 0.021855f
C225 VTAIL.n179 B 0.00979f
C226 VTAIL.n180 B 0.009246f
C227 VTAIL.n181 B 0.017207f
C228 VTAIL.n182 B 0.017207f
C229 VTAIL.n183 B 0.009246f
C230 VTAIL.n184 B 0.00979f
C231 VTAIL.n185 B 0.021855f
C232 VTAIL.n186 B 0.021855f
C233 VTAIL.n187 B 0.00979f
C234 VTAIL.n188 B 0.009246f
C235 VTAIL.n189 B 0.017207f
C236 VTAIL.n190 B 0.017207f
C237 VTAIL.n191 B 0.009246f
C238 VTAIL.n192 B 0.00979f
C239 VTAIL.n193 B 0.021855f
C240 VTAIL.n194 B 0.045259f
C241 VTAIL.n195 B 0.00979f
C242 VTAIL.n196 B 0.009246f
C243 VTAIL.n197 B 0.041183f
C244 VTAIL.n198 B 0.025156f
C245 VTAIL.n199 B 0.966181f
C246 VTAIL.n200 B 0.023025f
C247 VTAIL.n201 B 0.017207f
C248 VTAIL.n202 B 0.009246f
C249 VTAIL.n203 B 0.021855f
C250 VTAIL.n204 B 0.009518f
C251 VTAIL.n205 B 0.017207f
C252 VTAIL.n206 B 0.009518f
C253 VTAIL.n207 B 0.009246f
C254 VTAIL.n208 B 0.021855f
C255 VTAIL.n209 B 0.021855f
C256 VTAIL.n210 B 0.00979f
C257 VTAIL.n211 B 0.017207f
C258 VTAIL.n212 B 0.009246f
C259 VTAIL.n213 B 0.021855f
C260 VTAIL.n214 B 0.00979f
C261 VTAIL.n215 B 0.661408f
C262 VTAIL.n216 B 0.009246f
C263 VTAIL.t4 B 0.036664f
C264 VTAIL.n217 B 0.106228f
C265 VTAIL.n218 B 0.01545f
C266 VTAIL.n219 B 0.016391f
C267 VTAIL.n220 B 0.021855f
C268 VTAIL.n221 B 0.00979f
C269 VTAIL.n222 B 0.009246f
C270 VTAIL.n223 B 0.017207f
C271 VTAIL.n224 B 0.017207f
C272 VTAIL.n225 B 0.009246f
C273 VTAIL.n226 B 0.00979f
C274 VTAIL.n227 B 0.021855f
C275 VTAIL.n228 B 0.021855f
C276 VTAIL.n229 B 0.00979f
C277 VTAIL.n230 B 0.009246f
C278 VTAIL.n231 B 0.017207f
C279 VTAIL.n232 B 0.017207f
C280 VTAIL.n233 B 0.009246f
C281 VTAIL.n234 B 0.00979f
C282 VTAIL.n235 B 0.021855f
C283 VTAIL.n236 B 0.021855f
C284 VTAIL.n237 B 0.00979f
C285 VTAIL.n238 B 0.009246f
C286 VTAIL.n239 B 0.017207f
C287 VTAIL.n240 B 0.017207f
C288 VTAIL.n241 B 0.009246f
C289 VTAIL.n242 B 0.00979f
C290 VTAIL.n243 B 0.021855f
C291 VTAIL.n244 B 0.045259f
C292 VTAIL.n245 B 0.00979f
C293 VTAIL.n246 B 0.009246f
C294 VTAIL.n247 B 0.041183f
C295 VTAIL.n248 B 0.025156f
C296 VTAIL.n249 B 0.177763f
C297 VTAIL.n250 B 0.023025f
C298 VTAIL.n251 B 0.017207f
C299 VTAIL.n252 B 0.009246f
C300 VTAIL.n253 B 0.021855f
C301 VTAIL.n254 B 0.009518f
C302 VTAIL.n255 B 0.017207f
C303 VTAIL.n256 B 0.009518f
C304 VTAIL.n257 B 0.009246f
C305 VTAIL.n258 B 0.021855f
C306 VTAIL.n259 B 0.021855f
C307 VTAIL.n260 B 0.00979f
C308 VTAIL.n261 B 0.017207f
C309 VTAIL.n262 B 0.009246f
C310 VTAIL.n263 B 0.021855f
C311 VTAIL.n264 B 0.00979f
C312 VTAIL.n265 B 0.661408f
C313 VTAIL.n266 B 0.009246f
C314 VTAIL.t1 B 0.036664f
C315 VTAIL.n267 B 0.106228f
C316 VTAIL.n268 B 0.01545f
C317 VTAIL.n269 B 0.016391f
C318 VTAIL.n270 B 0.021855f
C319 VTAIL.n271 B 0.00979f
C320 VTAIL.n272 B 0.009246f
C321 VTAIL.n273 B 0.017207f
C322 VTAIL.n274 B 0.017207f
C323 VTAIL.n275 B 0.009246f
C324 VTAIL.n276 B 0.00979f
C325 VTAIL.n277 B 0.021855f
C326 VTAIL.n278 B 0.021855f
C327 VTAIL.n279 B 0.00979f
C328 VTAIL.n280 B 0.009246f
C329 VTAIL.n281 B 0.017207f
C330 VTAIL.n282 B 0.017207f
C331 VTAIL.n283 B 0.009246f
C332 VTAIL.n284 B 0.00979f
C333 VTAIL.n285 B 0.021855f
C334 VTAIL.n286 B 0.021855f
C335 VTAIL.n287 B 0.00979f
C336 VTAIL.n288 B 0.009246f
C337 VTAIL.n289 B 0.017207f
C338 VTAIL.n290 B 0.017207f
C339 VTAIL.n291 B 0.009246f
C340 VTAIL.n292 B 0.00979f
C341 VTAIL.n293 B 0.021855f
C342 VTAIL.n294 B 0.045259f
C343 VTAIL.n295 B 0.00979f
C344 VTAIL.n296 B 0.009246f
C345 VTAIL.n297 B 0.041183f
C346 VTAIL.n298 B 0.025156f
C347 VTAIL.n299 B 0.177763f
C348 VTAIL.n300 B 0.023025f
C349 VTAIL.n301 B 0.017207f
C350 VTAIL.n302 B 0.009246f
C351 VTAIL.n303 B 0.021855f
C352 VTAIL.n304 B 0.009518f
C353 VTAIL.n305 B 0.017207f
C354 VTAIL.n306 B 0.009518f
C355 VTAIL.n307 B 0.009246f
C356 VTAIL.n308 B 0.021855f
C357 VTAIL.n309 B 0.021855f
C358 VTAIL.n310 B 0.00979f
C359 VTAIL.n311 B 0.017207f
C360 VTAIL.n312 B 0.009246f
C361 VTAIL.n313 B 0.021855f
C362 VTAIL.n314 B 0.00979f
C363 VTAIL.n315 B 0.661408f
C364 VTAIL.n316 B 0.009246f
C365 VTAIL.t3 B 0.036664f
C366 VTAIL.n317 B 0.106228f
C367 VTAIL.n318 B 0.01545f
C368 VTAIL.n319 B 0.016391f
C369 VTAIL.n320 B 0.021855f
C370 VTAIL.n321 B 0.00979f
C371 VTAIL.n322 B 0.009246f
C372 VTAIL.n323 B 0.017207f
C373 VTAIL.n324 B 0.017207f
C374 VTAIL.n325 B 0.009246f
C375 VTAIL.n326 B 0.00979f
C376 VTAIL.n327 B 0.021855f
C377 VTAIL.n328 B 0.021855f
C378 VTAIL.n329 B 0.00979f
C379 VTAIL.n330 B 0.009246f
C380 VTAIL.n331 B 0.017207f
C381 VTAIL.n332 B 0.017207f
C382 VTAIL.n333 B 0.009246f
C383 VTAIL.n334 B 0.00979f
C384 VTAIL.n335 B 0.021855f
C385 VTAIL.n336 B 0.021855f
C386 VTAIL.n337 B 0.00979f
C387 VTAIL.n338 B 0.009246f
C388 VTAIL.n339 B 0.017207f
C389 VTAIL.n340 B 0.017207f
C390 VTAIL.n341 B 0.009246f
C391 VTAIL.n342 B 0.00979f
C392 VTAIL.n343 B 0.021855f
C393 VTAIL.n344 B 0.045259f
C394 VTAIL.n345 B 0.00979f
C395 VTAIL.n346 B 0.009246f
C396 VTAIL.n347 B 0.041183f
C397 VTAIL.n348 B 0.025156f
C398 VTAIL.n349 B 0.966181f
C399 VTAIL.n350 B 0.023025f
C400 VTAIL.n351 B 0.017207f
C401 VTAIL.n352 B 0.009246f
C402 VTAIL.n353 B 0.021855f
C403 VTAIL.n354 B 0.009518f
C404 VTAIL.n355 B 0.017207f
C405 VTAIL.n356 B 0.00979f
C406 VTAIL.n357 B 0.021855f
C407 VTAIL.n358 B 0.00979f
C408 VTAIL.n359 B 0.017207f
C409 VTAIL.n360 B 0.009246f
C410 VTAIL.n361 B 0.021855f
C411 VTAIL.n362 B 0.00979f
C412 VTAIL.n363 B 0.661408f
C413 VTAIL.n364 B 0.009246f
C414 VTAIL.t6 B 0.036664f
C415 VTAIL.n365 B 0.106228f
C416 VTAIL.n366 B 0.01545f
C417 VTAIL.n367 B 0.016391f
C418 VTAIL.n368 B 0.021855f
C419 VTAIL.n369 B 0.00979f
C420 VTAIL.n370 B 0.009246f
C421 VTAIL.n371 B 0.017207f
C422 VTAIL.n372 B 0.017207f
C423 VTAIL.n373 B 0.009246f
C424 VTAIL.n374 B 0.00979f
C425 VTAIL.n375 B 0.021855f
C426 VTAIL.n376 B 0.021855f
C427 VTAIL.n377 B 0.00979f
C428 VTAIL.n378 B 0.009246f
C429 VTAIL.n379 B 0.017207f
C430 VTAIL.n380 B 0.017207f
C431 VTAIL.n381 B 0.009246f
C432 VTAIL.n382 B 0.009246f
C433 VTAIL.n383 B 0.00979f
C434 VTAIL.n384 B 0.021855f
C435 VTAIL.n385 B 0.021855f
C436 VTAIL.n386 B 0.021855f
C437 VTAIL.n387 B 0.009518f
C438 VTAIL.n388 B 0.009246f
C439 VTAIL.n389 B 0.017207f
C440 VTAIL.n390 B 0.017207f
C441 VTAIL.n391 B 0.009246f
C442 VTAIL.n392 B 0.00979f
C443 VTAIL.n393 B 0.021855f
C444 VTAIL.n394 B 0.045259f
C445 VTAIL.n395 B 0.00979f
C446 VTAIL.n396 B 0.009246f
C447 VTAIL.n397 B 0.041183f
C448 VTAIL.n398 B 0.025156f
C449 VTAIL.n399 B 0.894844f
C450 VDD2.t3 B 0.198153f
C451 VDD2.t2 B 0.198153f
C452 VDD2.n0 B 2.30102f
C453 VDD2.t0 B 0.198153f
C454 VDD2.t1 B 0.198153f
C455 VDD2.n1 B 1.73658f
C456 VDD2.n2 B 3.45053f
C457 VN.t0 B 1.90466f
C458 VN.t1 B 1.90002f
C459 VN.n0 B 1.21763f
C460 VN.t3 B 1.90466f
C461 VN.t2 B 1.90002f
C462 VN.n1 B 2.54911f
.ends

