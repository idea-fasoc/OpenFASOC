* NGSPICE file created from diff_pair_sample_0923.ext - technology: sky130A

.subckt diff_pair_sample_0923 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=1.68795 ps=10.56 w=10.23 l=1.14
X1 VDD1.t7 VP.t0 VTAIL.t0 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X2 B.t11 B.t9 B.t10 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=0 ps=0 w=10.23 l=1.14
X3 B.t8 B.t6 B.t7 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=0 ps=0 w=10.23 l=1.14
X4 VTAIL.t14 VN.t1 VDD2.t5 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X5 B.t5 B.t3 B.t4 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=0 ps=0 w=10.23 l=1.14
X6 VDD2.t2 VN.t2 VTAIL.t13 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=3.9897 ps=21.24 w=10.23 l=1.14
X7 VTAIL.t12 VN.t3 VDD2.t6 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X8 B.t2 B.t0 B.t1 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=0 ps=0 w=10.23 l=1.14
X9 VDD2.t3 VN.t4 VTAIL.t11 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X10 VDD2.t7 VN.t5 VTAIL.t10 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X11 VTAIL.t5 VP.t1 VDD1.t6 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X12 VTAIL.t6 VP.t2 VDD1.t5 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=1.68795 ps=10.56 w=10.23 l=1.14
X13 VTAIL.t4 VP.t3 VDD1.t4 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=1.68795 ps=10.56 w=10.23 l=1.14
X14 VDD1.t3 VP.t4 VTAIL.t7 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X15 VDD1.t2 VP.t5 VTAIL.t3 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=3.9897 ps=21.24 w=10.23 l=1.14
X16 VTAIL.t9 VN.t6 VDD2.t4 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=3.9897 pd=21.24 as=1.68795 ps=10.56 w=10.23 l=1.14
X17 VTAIL.t2 VP.t6 VDD1.t1 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=1.68795 ps=10.56 w=10.23 l=1.14
X18 VDD1.t0 VP.t7 VTAIL.t1 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=3.9897 ps=21.24 w=10.23 l=1.14
X19 VDD2.t1 VN.t7 VTAIL.t8 w_n2440_n3014# sky130_fd_pr__pfet_01v8 ad=1.68795 pd=10.56 as=3.9897 ps=21.24 w=10.23 l=1.14
R0 VN.n3 VN.t0 274.06
R1 VN.n16 VN.t2 274.06
R2 VN.n11 VN.t7 250.936
R3 VN.n24 VN.t6 250.936
R4 VN.n4 VN.t4 216.267
R5 VN.n1 VN.t1 216.267
R6 VN.n17 VN.t3 216.267
R7 VN.n14 VN.t5 216.267
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN.n11 VN.n10 50.8919
R21 VN.n24 VN.n23 50.8919
R22 VN VN.n25 43.2263
R23 VN.n4 VN.n3 33.4814
R24 VN.n17 VN.n16 33.4814
R25 VN.n16 VN.n15 28.089
R26 VN.n3 VN.n2 28.089
R27 VN.n10 VN.n9 24.4675
R28 VN.n23 VN.n22 24.4675
R29 VN.n5 VN.n4 23.7335
R30 VN.n6 VN.n1 23.7335
R31 VN.n18 VN.n17 23.7335
R32 VN.n19 VN.n14 23.7335
R33 VN.n9 VN.n1 0.73451
R34 VN.n22 VN.n14 0.73451
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 75.3013
R45 VDD2.n2 VDD2.n0 75.3013
R46 VDD2 VDD2.n5 75.2985
R47 VDD2.n4 VDD2.n3 74.7232
R48 VDD2.n4 VDD2.n2 38.2368
R49 VDD2.n5 VDD2.t6 3.17792
R50 VDD2.n5 VDD2.t2 3.17792
R51 VDD2.n3 VDD2.t4 3.17792
R52 VDD2.n3 VDD2.t7 3.17792
R53 VDD2.n1 VDD2.t5 3.17792
R54 VDD2.n1 VDD2.t1 3.17792
R55 VDD2.n0 VDD2.t0 3.17792
R56 VDD2.n0 VDD2.t3 3.17792
R57 VDD2 VDD2.n4 0.69231
R58 VTAIL.n11 VTAIL.t6 61.2219
R59 VTAIL.n10 VTAIL.t13 61.2219
R60 VTAIL.n7 VTAIL.t9 61.2219
R61 VTAIL.n14 VTAIL.t3 61.2216
R62 VTAIL.n15 VTAIL.t8 61.2216
R63 VTAIL.n2 VTAIL.t15 61.2216
R64 VTAIL.n3 VTAIL.t1 61.2216
R65 VTAIL.n6 VTAIL.t4 61.2216
R66 VTAIL.n13 VTAIL.n12 58.0445
R67 VTAIL.n9 VTAIL.n8 58.0445
R68 VTAIL.n1 VTAIL.n0 58.0442
R69 VTAIL.n5 VTAIL.n4 58.0442
R70 VTAIL.n15 VTAIL.n14 22.4531
R71 VTAIL.n7 VTAIL.n6 22.4531
R72 VTAIL.n0 VTAIL.t11 3.17792
R73 VTAIL.n0 VTAIL.t14 3.17792
R74 VTAIL.n4 VTAIL.t0 3.17792
R75 VTAIL.n4 VTAIL.t5 3.17792
R76 VTAIL.n12 VTAIL.t7 3.17792
R77 VTAIL.n12 VTAIL.t2 3.17792
R78 VTAIL.n8 VTAIL.t10 3.17792
R79 VTAIL.n8 VTAIL.t12 3.17792
R80 VTAIL.n9 VTAIL.n7 1.26774
R81 VTAIL.n10 VTAIL.n9 1.26774
R82 VTAIL.n13 VTAIL.n11 1.26774
R83 VTAIL.n14 VTAIL.n13 1.26774
R84 VTAIL.n6 VTAIL.n5 1.26774
R85 VTAIL.n5 VTAIL.n3 1.26774
R86 VTAIL.n2 VTAIL.n1 1.26774
R87 VTAIL VTAIL.n15 1.20955
R88 VTAIL.n11 VTAIL.n10 0.470328
R89 VTAIL.n3 VTAIL.n2 0.470328
R90 VTAIL VTAIL.n1 0.0586897
R91 VP.n7 VP.t2 274.06
R92 VP.n17 VP.t3 250.936
R93 VP.n29 VP.t7 250.936
R94 VP.n15 VP.t5 250.936
R95 VP.n22 VP.t0 216.267
R96 VP.n1 VP.t1 216.267
R97 VP.n5 VP.t6 216.267
R98 VP.n8 VP.t4 216.267
R99 VP.n9 VP.n6 161.3
R100 VP.n11 VP.n10 161.3
R101 VP.n13 VP.n12 161.3
R102 VP.n14 VP.n4 161.3
R103 VP.n28 VP.n0 161.3
R104 VP.n27 VP.n26 161.3
R105 VP.n25 VP.n24 161.3
R106 VP.n23 VP.n2 161.3
R107 VP.n21 VP.n20 161.3
R108 VP.n19 VP.n3 161.3
R109 VP.n16 VP.n15 80.6037
R110 VP.n30 VP.n29 80.6037
R111 VP.n18 VP.n17 80.6037
R112 VP.n24 VP.n23 56.5193
R113 VP.n10 VP.n9 56.5193
R114 VP.n17 VP.n3 50.8919
R115 VP.n29 VP.n28 50.8919
R116 VP.n15 VP.n14 50.8919
R117 VP.n18 VP.n16 42.9408
R118 VP.n8 VP.n7 33.4814
R119 VP.n7 VP.n6 28.089
R120 VP.n21 VP.n3 24.4675
R121 VP.n28 VP.n27 24.4675
R122 VP.n14 VP.n13 24.4675
R123 VP.n23 VP.n22 23.7335
R124 VP.n24 VP.n1 23.7335
R125 VP.n10 VP.n5 23.7335
R126 VP.n9 VP.n8 23.7335
R127 VP.n22 VP.n21 0.73451
R128 VP.n27 VP.n1 0.73451
R129 VP.n13 VP.n5 0.73451
R130 VP.n16 VP.n4 0.285035
R131 VP.n19 VP.n18 0.285035
R132 VP.n30 VP.n0 0.285035
R133 VP.n11 VP.n6 0.189894
R134 VP.n12 VP.n11 0.189894
R135 VP.n12 VP.n4 0.189894
R136 VP.n20 VP.n19 0.189894
R137 VP.n20 VP.n2 0.189894
R138 VP.n25 VP.n2 0.189894
R139 VP.n26 VP.n25 0.189894
R140 VP.n26 VP.n0 0.189894
R141 VP VP.n30 0.146778
R142 VDD1 VDD1.n0 75.4151
R143 VDD1.n3 VDD1.n2 75.3013
R144 VDD1.n3 VDD1.n1 75.3013
R145 VDD1.n5 VDD1.n4 74.7231
R146 VDD1.n5 VDD1.n3 38.8199
R147 VDD1.n4 VDD1.t1 3.17792
R148 VDD1.n4 VDD1.t2 3.17792
R149 VDD1.n0 VDD1.t5 3.17792
R150 VDD1.n0 VDD1.t3 3.17792
R151 VDD1.n2 VDD1.t6 3.17792
R152 VDD1.n2 VDD1.t0 3.17792
R153 VDD1.n1 VDD1.t4 3.17792
R154 VDD1.n1 VDD1.t7 3.17792
R155 VDD1 VDD1.n5 0.575931
R156 B.n318 B.n317 585
R157 B.n316 B.n93 585
R158 B.n315 B.n314 585
R159 B.n313 B.n94 585
R160 B.n312 B.n311 585
R161 B.n310 B.n95 585
R162 B.n309 B.n308 585
R163 B.n307 B.n96 585
R164 B.n306 B.n305 585
R165 B.n304 B.n97 585
R166 B.n303 B.n302 585
R167 B.n301 B.n98 585
R168 B.n300 B.n299 585
R169 B.n298 B.n99 585
R170 B.n297 B.n296 585
R171 B.n295 B.n100 585
R172 B.n294 B.n293 585
R173 B.n292 B.n101 585
R174 B.n291 B.n290 585
R175 B.n289 B.n102 585
R176 B.n288 B.n287 585
R177 B.n286 B.n103 585
R178 B.n285 B.n284 585
R179 B.n283 B.n104 585
R180 B.n282 B.n281 585
R181 B.n280 B.n105 585
R182 B.n279 B.n278 585
R183 B.n277 B.n106 585
R184 B.n276 B.n275 585
R185 B.n274 B.n107 585
R186 B.n273 B.n272 585
R187 B.n271 B.n108 585
R188 B.n270 B.n269 585
R189 B.n268 B.n109 585
R190 B.n267 B.n266 585
R191 B.n265 B.n110 585
R192 B.n263 B.n262 585
R193 B.n261 B.n113 585
R194 B.n260 B.n259 585
R195 B.n258 B.n114 585
R196 B.n257 B.n256 585
R197 B.n255 B.n115 585
R198 B.n254 B.n253 585
R199 B.n252 B.n116 585
R200 B.n251 B.n250 585
R201 B.n249 B.n117 585
R202 B.n248 B.n247 585
R203 B.n243 B.n118 585
R204 B.n242 B.n241 585
R205 B.n240 B.n119 585
R206 B.n239 B.n238 585
R207 B.n237 B.n120 585
R208 B.n236 B.n235 585
R209 B.n234 B.n121 585
R210 B.n233 B.n232 585
R211 B.n231 B.n122 585
R212 B.n230 B.n229 585
R213 B.n228 B.n123 585
R214 B.n227 B.n226 585
R215 B.n225 B.n124 585
R216 B.n224 B.n223 585
R217 B.n222 B.n125 585
R218 B.n221 B.n220 585
R219 B.n219 B.n126 585
R220 B.n218 B.n217 585
R221 B.n216 B.n127 585
R222 B.n215 B.n214 585
R223 B.n213 B.n128 585
R224 B.n212 B.n211 585
R225 B.n210 B.n129 585
R226 B.n209 B.n208 585
R227 B.n207 B.n130 585
R228 B.n206 B.n205 585
R229 B.n204 B.n131 585
R230 B.n203 B.n202 585
R231 B.n201 B.n132 585
R232 B.n200 B.n199 585
R233 B.n198 B.n133 585
R234 B.n197 B.n196 585
R235 B.n195 B.n134 585
R236 B.n194 B.n193 585
R237 B.n192 B.n135 585
R238 B.n319 B.n92 585
R239 B.n321 B.n320 585
R240 B.n322 B.n91 585
R241 B.n324 B.n323 585
R242 B.n325 B.n90 585
R243 B.n327 B.n326 585
R244 B.n328 B.n89 585
R245 B.n330 B.n329 585
R246 B.n331 B.n88 585
R247 B.n333 B.n332 585
R248 B.n334 B.n87 585
R249 B.n336 B.n335 585
R250 B.n337 B.n86 585
R251 B.n339 B.n338 585
R252 B.n340 B.n85 585
R253 B.n342 B.n341 585
R254 B.n343 B.n84 585
R255 B.n345 B.n344 585
R256 B.n346 B.n83 585
R257 B.n348 B.n347 585
R258 B.n349 B.n82 585
R259 B.n351 B.n350 585
R260 B.n352 B.n81 585
R261 B.n354 B.n353 585
R262 B.n355 B.n80 585
R263 B.n357 B.n356 585
R264 B.n358 B.n79 585
R265 B.n360 B.n359 585
R266 B.n361 B.n78 585
R267 B.n363 B.n362 585
R268 B.n364 B.n77 585
R269 B.n366 B.n365 585
R270 B.n367 B.n76 585
R271 B.n369 B.n368 585
R272 B.n370 B.n75 585
R273 B.n372 B.n371 585
R274 B.n373 B.n74 585
R275 B.n375 B.n374 585
R276 B.n376 B.n73 585
R277 B.n378 B.n377 585
R278 B.n379 B.n72 585
R279 B.n381 B.n380 585
R280 B.n382 B.n71 585
R281 B.n384 B.n383 585
R282 B.n385 B.n70 585
R283 B.n387 B.n386 585
R284 B.n388 B.n69 585
R285 B.n390 B.n389 585
R286 B.n391 B.n68 585
R287 B.n393 B.n392 585
R288 B.n394 B.n67 585
R289 B.n396 B.n395 585
R290 B.n397 B.n66 585
R291 B.n399 B.n398 585
R292 B.n400 B.n65 585
R293 B.n402 B.n401 585
R294 B.n403 B.n64 585
R295 B.n405 B.n404 585
R296 B.n406 B.n63 585
R297 B.n408 B.n407 585
R298 B.n532 B.n531 585
R299 B.n530 B.n17 585
R300 B.n529 B.n528 585
R301 B.n527 B.n18 585
R302 B.n526 B.n525 585
R303 B.n524 B.n19 585
R304 B.n523 B.n522 585
R305 B.n521 B.n20 585
R306 B.n520 B.n519 585
R307 B.n518 B.n21 585
R308 B.n517 B.n516 585
R309 B.n515 B.n22 585
R310 B.n514 B.n513 585
R311 B.n512 B.n23 585
R312 B.n511 B.n510 585
R313 B.n509 B.n24 585
R314 B.n508 B.n507 585
R315 B.n506 B.n25 585
R316 B.n505 B.n504 585
R317 B.n503 B.n26 585
R318 B.n502 B.n501 585
R319 B.n500 B.n27 585
R320 B.n499 B.n498 585
R321 B.n497 B.n28 585
R322 B.n496 B.n495 585
R323 B.n494 B.n29 585
R324 B.n493 B.n492 585
R325 B.n491 B.n30 585
R326 B.n490 B.n489 585
R327 B.n488 B.n31 585
R328 B.n487 B.n486 585
R329 B.n485 B.n32 585
R330 B.n484 B.n483 585
R331 B.n482 B.n33 585
R332 B.n481 B.n480 585
R333 B.n479 B.n34 585
R334 B.n478 B.n477 585
R335 B.n476 B.n35 585
R336 B.n475 B.n474 585
R337 B.n473 B.n39 585
R338 B.n472 B.n471 585
R339 B.n470 B.n40 585
R340 B.n469 B.n468 585
R341 B.n467 B.n41 585
R342 B.n466 B.n465 585
R343 B.n464 B.n42 585
R344 B.n462 B.n461 585
R345 B.n460 B.n45 585
R346 B.n459 B.n458 585
R347 B.n457 B.n46 585
R348 B.n456 B.n455 585
R349 B.n454 B.n47 585
R350 B.n453 B.n452 585
R351 B.n451 B.n48 585
R352 B.n450 B.n449 585
R353 B.n448 B.n49 585
R354 B.n447 B.n446 585
R355 B.n445 B.n50 585
R356 B.n444 B.n443 585
R357 B.n442 B.n51 585
R358 B.n441 B.n440 585
R359 B.n439 B.n52 585
R360 B.n438 B.n437 585
R361 B.n436 B.n53 585
R362 B.n435 B.n434 585
R363 B.n433 B.n54 585
R364 B.n432 B.n431 585
R365 B.n430 B.n55 585
R366 B.n429 B.n428 585
R367 B.n427 B.n56 585
R368 B.n426 B.n425 585
R369 B.n424 B.n57 585
R370 B.n423 B.n422 585
R371 B.n421 B.n58 585
R372 B.n420 B.n419 585
R373 B.n418 B.n59 585
R374 B.n417 B.n416 585
R375 B.n415 B.n60 585
R376 B.n414 B.n413 585
R377 B.n412 B.n61 585
R378 B.n411 B.n410 585
R379 B.n409 B.n62 585
R380 B.n533 B.n16 585
R381 B.n535 B.n534 585
R382 B.n536 B.n15 585
R383 B.n538 B.n537 585
R384 B.n539 B.n14 585
R385 B.n541 B.n540 585
R386 B.n542 B.n13 585
R387 B.n544 B.n543 585
R388 B.n545 B.n12 585
R389 B.n547 B.n546 585
R390 B.n548 B.n11 585
R391 B.n550 B.n549 585
R392 B.n551 B.n10 585
R393 B.n553 B.n552 585
R394 B.n554 B.n9 585
R395 B.n556 B.n555 585
R396 B.n557 B.n8 585
R397 B.n559 B.n558 585
R398 B.n560 B.n7 585
R399 B.n562 B.n561 585
R400 B.n563 B.n6 585
R401 B.n565 B.n564 585
R402 B.n566 B.n5 585
R403 B.n568 B.n567 585
R404 B.n569 B.n4 585
R405 B.n571 B.n570 585
R406 B.n572 B.n3 585
R407 B.n574 B.n573 585
R408 B.n575 B.n0 585
R409 B.n2 B.n1 585
R410 B.n150 B.n149 585
R411 B.n152 B.n151 585
R412 B.n153 B.n148 585
R413 B.n155 B.n154 585
R414 B.n156 B.n147 585
R415 B.n158 B.n157 585
R416 B.n159 B.n146 585
R417 B.n161 B.n160 585
R418 B.n162 B.n145 585
R419 B.n164 B.n163 585
R420 B.n165 B.n144 585
R421 B.n167 B.n166 585
R422 B.n168 B.n143 585
R423 B.n170 B.n169 585
R424 B.n171 B.n142 585
R425 B.n173 B.n172 585
R426 B.n174 B.n141 585
R427 B.n176 B.n175 585
R428 B.n177 B.n140 585
R429 B.n179 B.n178 585
R430 B.n180 B.n139 585
R431 B.n182 B.n181 585
R432 B.n183 B.n138 585
R433 B.n185 B.n184 585
R434 B.n186 B.n137 585
R435 B.n188 B.n187 585
R436 B.n189 B.n136 585
R437 B.n191 B.n190 585
R438 B.n192 B.n191 569.379
R439 B.n317 B.n92 569.379
R440 B.n407 B.n62 569.379
R441 B.n533 B.n532 569.379
R442 B.n244 B.t9 420.058
R443 B.n111 B.t0 420.058
R444 B.n43 B.t3 420.058
R445 B.n36 B.t6 420.058
R446 B.n577 B.n576 256.663
R447 B.n576 B.n575 235.042
R448 B.n576 B.n2 235.042
R449 B.n193 B.n192 163.367
R450 B.n193 B.n134 163.367
R451 B.n197 B.n134 163.367
R452 B.n198 B.n197 163.367
R453 B.n199 B.n198 163.367
R454 B.n199 B.n132 163.367
R455 B.n203 B.n132 163.367
R456 B.n204 B.n203 163.367
R457 B.n205 B.n204 163.367
R458 B.n205 B.n130 163.367
R459 B.n209 B.n130 163.367
R460 B.n210 B.n209 163.367
R461 B.n211 B.n210 163.367
R462 B.n211 B.n128 163.367
R463 B.n215 B.n128 163.367
R464 B.n216 B.n215 163.367
R465 B.n217 B.n216 163.367
R466 B.n217 B.n126 163.367
R467 B.n221 B.n126 163.367
R468 B.n222 B.n221 163.367
R469 B.n223 B.n222 163.367
R470 B.n223 B.n124 163.367
R471 B.n227 B.n124 163.367
R472 B.n228 B.n227 163.367
R473 B.n229 B.n228 163.367
R474 B.n229 B.n122 163.367
R475 B.n233 B.n122 163.367
R476 B.n234 B.n233 163.367
R477 B.n235 B.n234 163.367
R478 B.n235 B.n120 163.367
R479 B.n239 B.n120 163.367
R480 B.n240 B.n239 163.367
R481 B.n241 B.n240 163.367
R482 B.n241 B.n118 163.367
R483 B.n248 B.n118 163.367
R484 B.n249 B.n248 163.367
R485 B.n250 B.n249 163.367
R486 B.n250 B.n116 163.367
R487 B.n254 B.n116 163.367
R488 B.n255 B.n254 163.367
R489 B.n256 B.n255 163.367
R490 B.n256 B.n114 163.367
R491 B.n260 B.n114 163.367
R492 B.n261 B.n260 163.367
R493 B.n262 B.n261 163.367
R494 B.n262 B.n110 163.367
R495 B.n267 B.n110 163.367
R496 B.n268 B.n267 163.367
R497 B.n269 B.n268 163.367
R498 B.n269 B.n108 163.367
R499 B.n273 B.n108 163.367
R500 B.n274 B.n273 163.367
R501 B.n275 B.n274 163.367
R502 B.n275 B.n106 163.367
R503 B.n279 B.n106 163.367
R504 B.n280 B.n279 163.367
R505 B.n281 B.n280 163.367
R506 B.n281 B.n104 163.367
R507 B.n285 B.n104 163.367
R508 B.n286 B.n285 163.367
R509 B.n287 B.n286 163.367
R510 B.n287 B.n102 163.367
R511 B.n291 B.n102 163.367
R512 B.n292 B.n291 163.367
R513 B.n293 B.n292 163.367
R514 B.n293 B.n100 163.367
R515 B.n297 B.n100 163.367
R516 B.n298 B.n297 163.367
R517 B.n299 B.n298 163.367
R518 B.n299 B.n98 163.367
R519 B.n303 B.n98 163.367
R520 B.n304 B.n303 163.367
R521 B.n305 B.n304 163.367
R522 B.n305 B.n96 163.367
R523 B.n309 B.n96 163.367
R524 B.n310 B.n309 163.367
R525 B.n311 B.n310 163.367
R526 B.n311 B.n94 163.367
R527 B.n315 B.n94 163.367
R528 B.n316 B.n315 163.367
R529 B.n317 B.n316 163.367
R530 B.n407 B.n406 163.367
R531 B.n406 B.n405 163.367
R532 B.n405 B.n64 163.367
R533 B.n401 B.n64 163.367
R534 B.n401 B.n400 163.367
R535 B.n400 B.n399 163.367
R536 B.n399 B.n66 163.367
R537 B.n395 B.n66 163.367
R538 B.n395 B.n394 163.367
R539 B.n394 B.n393 163.367
R540 B.n393 B.n68 163.367
R541 B.n389 B.n68 163.367
R542 B.n389 B.n388 163.367
R543 B.n388 B.n387 163.367
R544 B.n387 B.n70 163.367
R545 B.n383 B.n70 163.367
R546 B.n383 B.n382 163.367
R547 B.n382 B.n381 163.367
R548 B.n381 B.n72 163.367
R549 B.n377 B.n72 163.367
R550 B.n377 B.n376 163.367
R551 B.n376 B.n375 163.367
R552 B.n375 B.n74 163.367
R553 B.n371 B.n74 163.367
R554 B.n371 B.n370 163.367
R555 B.n370 B.n369 163.367
R556 B.n369 B.n76 163.367
R557 B.n365 B.n76 163.367
R558 B.n365 B.n364 163.367
R559 B.n364 B.n363 163.367
R560 B.n363 B.n78 163.367
R561 B.n359 B.n78 163.367
R562 B.n359 B.n358 163.367
R563 B.n358 B.n357 163.367
R564 B.n357 B.n80 163.367
R565 B.n353 B.n80 163.367
R566 B.n353 B.n352 163.367
R567 B.n352 B.n351 163.367
R568 B.n351 B.n82 163.367
R569 B.n347 B.n82 163.367
R570 B.n347 B.n346 163.367
R571 B.n346 B.n345 163.367
R572 B.n345 B.n84 163.367
R573 B.n341 B.n84 163.367
R574 B.n341 B.n340 163.367
R575 B.n340 B.n339 163.367
R576 B.n339 B.n86 163.367
R577 B.n335 B.n86 163.367
R578 B.n335 B.n334 163.367
R579 B.n334 B.n333 163.367
R580 B.n333 B.n88 163.367
R581 B.n329 B.n88 163.367
R582 B.n329 B.n328 163.367
R583 B.n328 B.n327 163.367
R584 B.n327 B.n90 163.367
R585 B.n323 B.n90 163.367
R586 B.n323 B.n322 163.367
R587 B.n322 B.n321 163.367
R588 B.n321 B.n92 163.367
R589 B.n532 B.n17 163.367
R590 B.n528 B.n17 163.367
R591 B.n528 B.n527 163.367
R592 B.n527 B.n526 163.367
R593 B.n526 B.n19 163.367
R594 B.n522 B.n19 163.367
R595 B.n522 B.n521 163.367
R596 B.n521 B.n520 163.367
R597 B.n520 B.n21 163.367
R598 B.n516 B.n21 163.367
R599 B.n516 B.n515 163.367
R600 B.n515 B.n514 163.367
R601 B.n514 B.n23 163.367
R602 B.n510 B.n23 163.367
R603 B.n510 B.n509 163.367
R604 B.n509 B.n508 163.367
R605 B.n508 B.n25 163.367
R606 B.n504 B.n25 163.367
R607 B.n504 B.n503 163.367
R608 B.n503 B.n502 163.367
R609 B.n502 B.n27 163.367
R610 B.n498 B.n27 163.367
R611 B.n498 B.n497 163.367
R612 B.n497 B.n496 163.367
R613 B.n496 B.n29 163.367
R614 B.n492 B.n29 163.367
R615 B.n492 B.n491 163.367
R616 B.n491 B.n490 163.367
R617 B.n490 B.n31 163.367
R618 B.n486 B.n31 163.367
R619 B.n486 B.n485 163.367
R620 B.n485 B.n484 163.367
R621 B.n484 B.n33 163.367
R622 B.n480 B.n33 163.367
R623 B.n480 B.n479 163.367
R624 B.n479 B.n478 163.367
R625 B.n478 B.n35 163.367
R626 B.n474 B.n35 163.367
R627 B.n474 B.n473 163.367
R628 B.n473 B.n472 163.367
R629 B.n472 B.n40 163.367
R630 B.n468 B.n40 163.367
R631 B.n468 B.n467 163.367
R632 B.n467 B.n466 163.367
R633 B.n466 B.n42 163.367
R634 B.n461 B.n42 163.367
R635 B.n461 B.n460 163.367
R636 B.n460 B.n459 163.367
R637 B.n459 B.n46 163.367
R638 B.n455 B.n46 163.367
R639 B.n455 B.n454 163.367
R640 B.n454 B.n453 163.367
R641 B.n453 B.n48 163.367
R642 B.n449 B.n48 163.367
R643 B.n449 B.n448 163.367
R644 B.n448 B.n447 163.367
R645 B.n447 B.n50 163.367
R646 B.n443 B.n50 163.367
R647 B.n443 B.n442 163.367
R648 B.n442 B.n441 163.367
R649 B.n441 B.n52 163.367
R650 B.n437 B.n52 163.367
R651 B.n437 B.n436 163.367
R652 B.n436 B.n435 163.367
R653 B.n435 B.n54 163.367
R654 B.n431 B.n54 163.367
R655 B.n431 B.n430 163.367
R656 B.n430 B.n429 163.367
R657 B.n429 B.n56 163.367
R658 B.n425 B.n56 163.367
R659 B.n425 B.n424 163.367
R660 B.n424 B.n423 163.367
R661 B.n423 B.n58 163.367
R662 B.n419 B.n58 163.367
R663 B.n419 B.n418 163.367
R664 B.n418 B.n417 163.367
R665 B.n417 B.n60 163.367
R666 B.n413 B.n60 163.367
R667 B.n413 B.n412 163.367
R668 B.n412 B.n411 163.367
R669 B.n411 B.n62 163.367
R670 B.n534 B.n533 163.367
R671 B.n534 B.n15 163.367
R672 B.n538 B.n15 163.367
R673 B.n539 B.n538 163.367
R674 B.n540 B.n539 163.367
R675 B.n540 B.n13 163.367
R676 B.n544 B.n13 163.367
R677 B.n545 B.n544 163.367
R678 B.n546 B.n545 163.367
R679 B.n546 B.n11 163.367
R680 B.n550 B.n11 163.367
R681 B.n551 B.n550 163.367
R682 B.n552 B.n551 163.367
R683 B.n552 B.n9 163.367
R684 B.n556 B.n9 163.367
R685 B.n557 B.n556 163.367
R686 B.n558 B.n557 163.367
R687 B.n558 B.n7 163.367
R688 B.n562 B.n7 163.367
R689 B.n563 B.n562 163.367
R690 B.n564 B.n563 163.367
R691 B.n564 B.n5 163.367
R692 B.n568 B.n5 163.367
R693 B.n569 B.n568 163.367
R694 B.n570 B.n569 163.367
R695 B.n570 B.n3 163.367
R696 B.n574 B.n3 163.367
R697 B.n575 B.n574 163.367
R698 B.n150 B.n2 163.367
R699 B.n151 B.n150 163.367
R700 B.n151 B.n148 163.367
R701 B.n155 B.n148 163.367
R702 B.n156 B.n155 163.367
R703 B.n157 B.n156 163.367
R704 B.n157 B.n146 163.367
R705 B.n161 B.n146 163.367
R706 B.n162 B.n161 163.367
R707 B.n163 B.n162 163.367
R708 B.n163 B.n144 163.367
R709 B.n167 B.n144 163.367
R710 B.n168 B.n167 163.367
R711 B.n169 B.n168 163.367
R712 B.n169 B.n142 163.367
R713 B.n173 B.n142 163.367
R714 B.n174 B.n173 163.367
R715 B.n175 B.n174 163.367
R716 B.n175 B.n140 163.367
R717 B.n179 B.n140 163.367
R718 B.n180 B.n179 163.367
R719 B.n181 B.n180 163.367
R720 B.n181 B.n138 163.367
R721 B.n185 B.n138 163.367
R722 B.n186 B.n185 163.367
R723 B.n187 B.n186 163.367
R724 B.n187 B.n136 163.367
R725 B.n191 B.n136 163.367
R726 B.n111 B.t1 136.685
R727 B.n43 B.t5 136.685
R728 B.n244 B.t10 136.673
R729 B.n36 B.t8 136.673
R730 B.n112 B.t2 108.175
R731 B.n44 B.t4 108.175
R732 B.n245 B.t11 108.163
R733 B.n37 B.t7 108.163
R734 B.n246 B.n245 59.5399
R735 B.n264 B.n112 59.5399
R736 B.n463 B.n44 59.5399
R737 B.n38 B.n37 59.5399
R738 B.n531 B.n16 36.9956
R739 B.n409 B.n408 36.9956
R740 B.n319 B.n318 36.9956
R741 B.n190 B.n135 36.9956
R742 B.n245 B.n244 28.5096
R743 B.n112 B.n111 28.5096
R744 B.n44 B.n43 28.5096
R745 B.n37 B.n36 28.5096
R746 B B.n577 18.0485
R747 B.n535 B.n16 10.6151
R748 B.n536 B.n535 10.6151
R749 B.n537 B.n536 10.6151
R750 B.n537 B.n14 10.6151
R751 B.n541 B.n14 10.6151
R752 B.n542 B.n541 10.6151
R753 B.n543 B.n542 10.6151
R754 B.n543 B.n12 10.6151
R755 B.n547 B.n12 10.6151
R756 B.n548 B.n547 10.6151
R757 B.n549 B.n548 10.6151
R758 B.n549 B.n10 10.6151
R759 B.n553 B.n10 10.6151
R760 B.n554 B.n553 10.6151
R761 B.n555 B.n554 10.6151
R762 B.n555 B.n8 10.6151
R763 B.n559 B.n8 10.6151
R764 B.n560 B.n559 10.6151
R765 B.n561 B.n560 10.6151
R766 B.n561 B.n6 10.6151
R767 B.n565 B.n6 10.6151
R768 B.n566 B.n565 10.6151
R769 B.n567 B.n566 10.6151
R770 B.n567 B.n4 10.6151
R771 B.n571 B.n4 10.6151
R772 B.n572 B.n571 10.6151
R773 B.n573 B.n572 10.6151
R774 B.n573 B.n0 10.6151
R775 B.n531 B.n530 10.6151
R776 B.n530 B.n529 10.6151
R777 B.n529 B.n18 10.6151
R778 B.n525 B.n18 10.6151
R779 B.n525 B.n524 10.6151
R780 B.n524 B.n523 10.6151
R781 B.n523 B.n20 10.6151
R782 B.n519 B.n20 10.6151
R783 B.n519 B.n518 10.6151
R784 B.n518 B.n517 10.6151
R785 B.n517 B.n22 10.6151
R786 B.n513 B.n22 10.6151
R787 B.n513 B.n512 10.6151
R788 B.n512 B.n511 10.6151
R789 B.n511 B.n24 10.6151
R790 B.n507 B.n24 10.6151
R791 B.n507 B.n506 10.6151
R792 B.n506 B.n505 10.6151
R793 B.n505 B.n26 10.6151
R794 B.n501 B.n26 10.6151
R795 B.n501 B.n500 10.6151
R796 B.n500 B.n499 10.6151
R797 B.n499 B.n28 10.6151
R798 B.n495 B.n28 10.6151
R799 B.n495 B.n494 10.6151
R800 B.n494 B.n493 10.6151
R801 B.n493 B.n30 10.6151
R802 B.n489 B.n30 10.6151
R803 B.n489 B.n488 10.6151
R804 B.n488 B.n487 10.6151
R805 B.n487 B.n32 10.6151
R806 B.n483 B.n32 10.6151
R807 B.n483 B.n482 10.6151
R808 B.n482 B.n481 10.6151
R809 B.n481 B.n34 10.6151
R810 B.n477 B.n476 10.6151
R811 B.n476 B.n475 10.6151
R812 B.n475 B.n39 10.6151
R813 B.n471 B.n39 10.6151
R814 B.n471 B.n470 10.6151
R815 B.n470 B.n469 10.6151
R816 B.n469 B.n41 10.6151
R817 B.n465 B.n41 10.6151
R818 B.n465 B.n464 10.6151
R819 B.n462 B.n45 10.6151
R820 B.n458 B.n45 10.6151
R821 B.n458 B.n457 10.6151
R822 B.n457 B.n456 10.6151
R823 B.n456 B.n47 10.6151
R824 B.n452 B.n47 10.6151
R825 B.n452 B.n451 10.6151
R826 B.n451 B.n450 10.6151
R827 B.n450 B.n49 10.6151
R828 B.n446 B.n49 10.6151
R829 B.n446 B.n445 10.6151
R830 B.n445 B.n444 10.6151
R831 B.n444 B.n51 10.6151
R832 B.n440 B.n51 10.6151
R833 B.n440 B.n439 10.6151
R834 B.n439 B.n438 10.6151
R835 B.n438 B.n53 10.6151
R836 B.n434 B.n53 10.6151
R837 B.n434 B.n433 10.6151
R838 B.n433 B.n432 10.6151
R839 B.n432 B.n55 10.6151
R840 B.n428 B.n55 10.6151
R841 B.n428 B.n427 10.6151
R842 B.n427 B.n426 10.6151
R843 B.n426 B.n57 10.6151
R844 B.n422 B.n57 10.6151
R845 B.n422 B.n421 10.6151
R846 B.n421 B.n420 10.6151
R847 B.n420 B.n59 10.6151
R848 B.n416 B.n59 10.6151
R849 B.n416 B.n415 10.6151
R850 B.n415 B.n414 10.6151
R851 B.n414 B.n61 10.6151
R852 B.n410 B.n61 10.6151
R853 B.n410 B.n409 10.6151
R854 B.n408 B.n63 10.6151
R855 B.n404 B.n63 10.6151
R856 B.n404 B.n403 10.6151
R857 B.n403 B.n402 10.6151
R858 B.n402 B.n65 10.6151
R859 B.n398 B.n65 10.6151
R860 B.n398 B.n397 10.6151
R861 B.n397 B.n396 10.6151
R862 B.n396 B.n67 10.6151
R863 B.n392 B.n67 10.6151
R864 B.n392 B.n391 10.6151
R865 B.n391 B.n390 10.6151
R866 B.n390 B.n69 10.6151
R867 B.n386 B.n69 10.6151
R868 B.n386 B.n385 10.6151
R869 B.n385 B.n384 10.6151
R870 B.n384 B.n71 10.6151
R871 B.n380 B.n71 10.6151
R872 B.n380 B.n379 10.6151
R873 B.n379 B.n378 10.6151
R874 B.n378 B.n73 10.6151
R875 B.n374 B.n73 10.6151
R876 B.n374 B.n373 10.6151
R877 B.n373 B.n372 10.6151
R878 B.n372 B.n75 10.6151
R879 B.n368 B.n75 10.6151
R880 B.n368 B.n367 10.6151
R881 B.n367 B.n366 10.6151
R882 B.n366 B.n77 10.6151
R883 B.n362 B.n77 10.6151
R884 B.n362 B.n361 10.6151
R885 B.n361 B.n360 10.6151
R886 B.n360 B.n79 10.6151
R887 B.n356 B.n79 10.6151
R888 B.n356 B.n355 10.6151
R889 B.n355 B.n354 10.6151
R890 B.n354 B.n81 10.6151
R891 B.n350 B.n81 10.6151
R892 B.n350 B.n349 10.6151
R893 B.n349 B.n348 10.6151
R894 B.n348 B.n83 10.6151
R895 B.n344 B.n83 10.6151
R896 B.n344 B.n343 10.6151
R897 B.n343 B.n342 10.6151
R898 B.n342 B.n85 10.6151
R899 B.n338 B.n85 10.6151
R900 B.n338 B.n337 10.6151
R901 B.n337 B.n336 10.6151
R902 B.n336 B.n87 10.6151
R903 B.n332 B.n87 10.6151
R904 B.n332 B.n331 10.6151
R905 B.n331 B.n330 10.6151
R906 B.n330 B.n89 10.6151
R907 B.n326 B.n89 10.6151
R908 B.n326 B.n325 10.6151
R909 B.n325 B.n324 10.6151
R910 B.n324 B.n91 10.6151
R911 B.n320 B.n91 10.6151
R912 B.n320 B.n319 10.6151
R913 B.n149 B.n1 10.6151
R914 B.n152 B.n149 10.6151
R915 B.n153 B.n152 10.6151
R916 B.n154 B.n153 10.6151
R917 B.n154 B.n147 10.6151
R918 B.n158 B.n147 10.6151
R919 B.n159 B.n158 10.6151
R920 B.n160 B.n159 10.6151
R921 B.n160 B.n145 10.6151
R922 B.n164 B.n145 10.6151
R923 B.n165 B.n164 10.6151
R924 B.n166 B.n165 10.6151
R925 B.n166 B.n143 10.6151
R926 B.n170 B.n143 10.6151
R927 B.n171 B.n170 10.6151
R928 B.n172 B.n171 10.6151
R929 B.n172 B.n141 10.6151
R930 B.n176 B.n141 10.6151
R931 B.n177 B.n176 10.6151
R932 B.n178 B.n177 10.6151
R933 B.n178 B.n139 10.6151
R934 B.n182 B.n139 10.6151
R935 B.n183 B.n182 10.6151
R936 B.n184 B.n183 10.6151
R937 B.n184 B.n137 10.6151
R938 B.n188 B.n137 10.6151
R939 B.n189 B.n188 10.6151
R940 B.n190 B.n189 10.6151
R941 B.n194 B.n135 10.6151
R942 B.n195 B.n194 10.6151
R943 B.n196 B.n195 10.6151
R944 B.n196 B.n133 10.6151
R945 B.n200 B.n133 10.6151
R946 B.n201 B.n200 10.6151
R947 B.n202 B.n201 10.6151
R948 B.n202 B.n131 10.6151
R949 B.n206 B.n131 10.6151
R950 B.n207 B.n206 10.6151
R951 B.n208 B.n207 10.6151
R952 B.n208 B.n129 10.6151
R953 B.n212 B.n129 10.6151
R954 B.n213 B.n212 10.6151
R955 B.n214 B.n213 10.6151
R956 B.n214 B.n127 10.6151
R957 B.n218 B.n127 10.6151
R958 B.n219 B.n218 10.6151
R959 B.n220 B.n219 10.6151
R960 B.n220 B.n125 10.6151
R961 B.n224 B.n125 10.6151
R962 B.n225 B.n224 10.6151
R963 B.n226 B.n225 10.6151
R964 B.n226 B.n123 10.6151
R965 B.n230 B.n123 10.6151
R966 B.n231 B.n230 10.6151
R967 B.n232 B.n231 10.6151
R968 B.n232 B.n121 10.6151
R969 B.n236 B.n121 10.6151
R970 B.n237 B.n236 10.6151
R971 B.n238 B.n237 10.6151
R972 B.n238 B.n119 10.6151
R973 B.n242 B.n119 10.6151
R974 B.n243 B.n242 10.6151
R975 B.n247 B.n243 10.6151
R976 B.n251 B.n117 10.6151
R977 B.n252 B.n251 10.6151
R978 B.n253 B.n252 10.6151
R979 B.n253 B.n115 10.6151
R980 B.n257 B.n115 10.6151
R981 B.n258 B.n257 10.6151
R982 B.n259 B.n258 10.6151
R983 B.n259 B.n113 10.6151
R984 B.n263 B.n113 10.6151
R985 B.n266 B.n265 10.6151
R986 B.n266 B.n109 10.6151
R987 B.n270 B.n109 10.6151
R988 B.n271 B.n270 10.6151
R989 B.n272 B.n271 10.6151
R990 B.n272 B.n107 10.6151
R991 B.n276 B.n107 10.6151
R992 B.n277 B.n276 10.6151
R993 B.n278 B.n277 10.6151
R994 B.n278 B.n105 10.6151
R995 B.n282 B.n105 10.6151
R996 B.n283 B.n282 10.6151
R997 B.n284 B.n283 10.6151
R998 B.n284 B.n103 10.6151
R999 B.n288 B.n103 10.6151
R1000 B.n289 B.n288 10.6151
R1001 B.n290 B.n289 10.6151
R1002 B.n290 B.n101 10.6151
R1003 B.n294 B.n101 10.6151
R1004 B.n295 B.n294 10.6151
R1005 B.n296 B.n295 10.6151
R1006 B.n296 B.n99 10.6151
R1007 B.n300 B.n99 10.6151
R1008 B.n301 B.n300 10.6151
R1009 B.n302 B.n301 10.6151
R1010 B.n302 B.n97 10.6151
R1011 B.n306 B.n97 10.6151
R1012 B.n307 B.n306 10.6151
R1013 B.n308 B.n307 10.6151
R1014 B.n308 B.n95 10.6151
R1015 B.n312 B.n95 10.6151
R1016 B.n313 B.n312 10.6151
R1017 B.n314 B.n313 10.6151
R1018 B.n314 B.n93 10.6151
R1019 B.n318 B.n93 10.6151
R1020 B.n38 B.n34 9.36635
R1021 B.n463 B.n462 9.36635
R1022 B.n247 B.n246 9.36635
R1023 B.n265 B.n264 9.36635
R1024 B.n577 B.n0 8.11757
R1025 B.n577 B.n1 8.11757
R1026 B.n477 B.n38 1.24928
R1027 B.n464 B.n463 1.24928
R1028 B.n246 B.n117 1.24928
R1029 B.n264 B.n263 1.24928
C0 B VN 0.863983f
C1 B VP 1.37999f
C2 VDD2 VN 5.90952f
C3 VDD2 VP 0.364368f
C4 VTAIL VN 5.90332f
C5 B VDD2 1.20709f
C6 VP VTAIL 5.91743f
C7 B VTAIL 3.65848f
C8 VDD2 VTAIL 8.21562f
C9 w_n2440_n3014# VN 4.5136f
C10 w_n2440_n3014# VP 4.82606f
C11 VN VDD1 0.149145f
C12 VP VDD1 6.12409f
C13 B w_n2440_n3014# 7.384359f
C14 w_n2440_n3014# VDD2 1.47207f
C15 B VDD1 1.1568f
C16 VDD2 VDD1 1.04669f
C17 w_n2440_n3014# VTAIL 3.73473f
C18 VTAIL VDD1 8.170991f
C19 VP VN 5.54636f
C20 w_n2440_n3014# VDD1 1.41877f
C21 VDD2 VSUBS 1.356899f
C22 VDD1 VSUBS 1.744157f
C23 VTAIL VSUBS 0.962098f
C24 VN VSUBS 4.94391f
C25 VP VSUBS 2.049992f
C26 B VSUBS 3.226238f
C27 w_n2440_n3014# VSUBS 90.797295f
C28 B.n0 VSUBS 0.007048f
C29 B.n1 VSUBS 0.007048f
C30 B.n2 VSUBS 0.010423f
C31 B.n3 VSUBS 0.007987f
C32 B.n4 VSUBS 0.007987f
C33 B.n5 VSUBS 0.007987f
C34 B.n6 VSUBS 0.007987f
C35 B.n7 VSUBS 0.007987f
C36 B.n8 VSUBS 0.007987f
C37 B.n9 VSUBS 0.007987f
C38 B.n10 VSUBS 0.007987f
C39 B.n11 VSUBS 0.007987f
C40 B.n12 VSUBS 0.007987f
C41 B.n13 VSUBS 0.007987f
C42 B.n14 VSUBS 0.007987f
C43 B.n15 VSUBS 0.007987f
C44 B.n16 VSUBS 0.019904f
C45 B.n17 VSUBS 0.007987f
C46 B.n18 VSUBS 0.007987f
C47 B.n19 VSUBS 0.007987f
C48 B.n20 VSUBS 0.007987f
C49 B.n21 VSUBS 0.007987f
C50 B.n22 VSUBS 0.007987f
C51 B.n23 VSUBS 0.007987f
C52 B.n24 VSUBS 0.007987f
C53 B.n25 VSUBS 0.007987f
C54 B.n26 VSUBS 0.007987f
C55 B.n27 VSUBS 0.007987f
C56 B.n28 VSUBS 0.007987f
C57 B.n29 VSUBS 0.007987f
C58 B.n30 VSUBS 0.007987f
C59 B.n31 VSUBS 0.007987f
C60 B.n32 VSUBS 0.007987f
C61 B.n33 VSUBS 0.007987f
C62 B.n34 VSUBS 0.007517f
C63 B.n35 VSUBS 0.007987f
C64 B.t7 VSUBS 0.373356f
C65 B.t8 VSUBS 0.386595f
C66 B.t6 VSUBS 0.575948f
C67 B.n36 VSUBS 0.162629f
C68 B.n37 VSUBS 0.07486f
C69 B.n38 VSUBS 0.018506f
C70 B.n39 VSUBS 0.007987f
C71 B.n40 VSUBS 0.007987f
C72 B.n41 VSUBS 0.007987f
C73 B.n42 VSUBS 0.007987f
C74 B.t4 VSUBS 0.37335f
C75 B.t5 VSUBS 0.386589f
C76 B.t3 VSUBS 0.575948f
C77 B.n43 VSUBS 0.162634f
C78 B.n44 VSUBS 0.074865f
C79 B.n45 VSUBS 0.007987f
C80 B.n46 VSUBS 0.007987f
C81 B.n47 VSUBS 0.007987f
C82 B.n48 VSUBS 0.007987f
C83 B.n49 VSUBS 0.007987f
C84 B.n50 VSUBS 0.007987f
C85 B.n51 VSUBS 0.007987f
C86 B.n52 VSUBS 0.007987f
C87 B.n53 VSUBS 0.007987f
C88 B.n54 VSUBS 0.007987f
C89 B.n55 VSUBS 0.007987f
C90 B.n56 VSUBS 0.007987f
C91 B.n57 VSUBS 0.007987f
C92 B.n58 VSUBS 0.007987f
C93 B.n59 VSUBS 0.007987f
C94 B.n60 VSUBS 0.007987f
C95 B.n61 VSUBS 0.007987f
C96 B.n62 VSUBS 0.020737f
C97 B.n63 VSUBS 0.007987f
C98 B.n64 VSUBS 0.007987f
C99 B.n65 VSUBS 0.007987f
C100 B.n66 VSUBS 0.007987f
C101 B.n67 VSUBS 0.007987f
C102 B.n68 VSUBS 0.007987f
C103 B.n69 VSUBS 0.007987f
C104 B.n70 VSUBS 0.007987f
C105 B.n71 VSUBS 0.007987f
C106 B.n72 VSUBS 0.007987f
C107 B.n73 VSUBS 0.007987f
C108 B.n74 VSUBS 0.007987f
C109 B.n75 VSUBS 0.007987f
C110 B.n76 VSUBS 0.007987f
C111 B.n77 VSUBS 0.007987f
C112 B.n78 VSUBS 0.007987f
C113 B.n79 VSUBS 0.007987f
C114 B.n80 VSUBS 0.007987f
C115 B.n81 VSUBS 0.007987f
C116 B.n82 VSUBS 0.007987f
C117 B.n83 VSUBS 0.007987f
C118 B.n84 VSUBS 0.007987f
C119 B.n85 VSUBS 0.007987f
C120 B.n86 VSUBS 0.007987f
C121 B.n87 VSUBS 0.007987f
C122 B.n88 VSUBS 0.007987f
C123 B.n89 VSUBS 0.007987f
C124 B.n90 VSUBS 0.007987f
C125 B.n91 VSUBS 0.007987f
C126 B.n92 VSUBS 0.019904f
C127 B.n93 VSUBS 0.007987f
C128 B.n94 VSUBS 0.007987f
C129 B.n95 VSUBS 0.007987f
C130 B.n96 VSUBS 0.007987f
C131 B.n97 VSUBS 0.007987f
C132 B.n98 VSUBS 0.007987f
C133 B.n99 VSUBS 0.007987f
C134 B.n100 VSUBS 0.007987f
C135 B.n101 VSUBS 0.007987f
C136 B.n102 VSUBS 0.007987f
C137 B.n103 VSUBS 0.007987f
C138 B.n104 VSUBS 0.007987f
C139 B.n105 VSUBS 0.007987f
C140 B.n106 VSUBS 0.007987f
C141 B.n107 VSUBS 0.007987f
C142 B.n108 VSUBS 0.007987f
C143 B.n109 VSUBS 0.007987f
C144 B.n110 VSUBS 0.007987f
C145 B.t2 VSUBS 0.37335f
C146 B.t1 VSUBS 0.386589f
C147 B.t0 VSUBS 0.575948f
C148 B.n111 VSUBS 0.162634f
C149 B.n112 VSUBS 0.074865f
C150 B.n113 VSUBS 0.007987f
C151 B.n114 VSUBS 0.007987f
C152 B.n115 VSUBS 0.007987f
C153 B.n116 VSUBS 0.007987f
C154 B.n117 VSUBS 0.004463f
C155 B.n118 VSUBS 0.007987f
C156 B.n119 VSUBS 0.007987f
C157 B.n120 VSUBS 0.007987f
C158 B.n121 VSUBS 0.007987f
C159 B.n122 VSUBS 0.007987f
C160 B.n123 VSUBS 0.007987f
C161 B.n124 VSUBS 0.007987f
C162 B.n125 VSUBS 0.007987f
C163 B.n126 VSUBS 0.007987f
C164 B.n127 VSUBS 0.007987f
C165 B.n128 VSUBS 0.007987f
C166 B.n129 VSUBS 0.007987f
C167 B.n130 VSUBS 0.007987f
C168 B.n131 VSUBS 0.007987f
C169 B.n132 VSUBS 0.007987f
C170 B.n133 VSUBS 0.007987f
C171 B.n134 VSUBS 0.007987f
C172 B.n135 VSUBS 0.020737f
C173 B.n136 VSUBS 0.007987f
C174 B.n137 VSUBS 0.007987f
C175 B.n138 VSUBS 0.007987f
C176 B.n139 VSUBS 0.007987f
C177 B.n140 VSUBS 0.007987f
C178 B.n141 VSUBS 0.007987f
C179 B.n142 VSUBS 0.007987f
C180 B.n143 VSUBS 0.007987f
C181 B.n144 VSUBS 0.007987f
C182 B.n145 VSUBS 0.007987f
C183 B.n146 VSUBS 0.007987f
C184 B.n147 VSUBS 0.007987f
C185 B.n148 VSUBS 0.007987f
C186 B.n149 VSUBS 0.007987f
C187 B.n150 VSUBS 0.007987f
C188 B.n151 VSUBS 0.007987f
C189 B.n152 VSUBS 0.007987f
C190 B.n153 VSUBS 0.007987f
C191 B.n154 VSUBS 0.007987f
C192 B.n155 VSUBS 0.007987f
C193 B.n156 VSUBS 0.007987f
C194 B.n157 VSUBS 0.007987f
C195 B.n158 VSUBS 0.007987f
C196 B.n159 VSUBS 0.007987f
C197 B.n160 VSUBS 0.007987f
C198 B.n161 VSUBS 0.007987f
C199 B.n162 VSUBS 0.007987f
C200 B.n163 VSUBS 0.007987f
C201 B.n164 VSUBS 0.007987f
C202 B.n165 VSUBS 0.007987f
C203 B.n166 VSUBS 0.007987f
C204 B.n167 VSUBS 0.007987f
C205 B.n168 VSUBS 0.007987f
C206 B.n169 VSUBS 0.007987f
C207 B.n170 VSUBS 0.007987f
C208 B.n171 VSUBS 0.007987f
C209 B.n172 VSUBS 0.007987f
C210 B.n173 VSUBS 0.007987f
C211 B.n174 VSUBS 0.007987f
C212 B.n175 VSUBS 0.007987f
C213 B.n176 VSUBS 0.007987f
C214 B.n177 VSUBS 0.007987f
C215 B.n178 VSUBS 0.007987f
C216 B.n179 VSUBS 0.007987f
C217 B.n180 VSUBS 0.007987f
C218 B.n181 VSUBS 0.007987f
C219 B.n182 VSUBS 0.007987f
C220 B.n183 VSUBS 0.007987f
C221 B.n184 VSUBS 0.007987f
C222 B.n185 VSUBS 0.007987f
C223 B.n186 VSUBS 0.007987f
C224 B.n187 VSUBS 0.007987f
C225 B.n188 VSUBS 0.007987f
C226 B.n189 VSUBS 0.007987f
C227 B.n190 VSUBS 0.019904f
C228 B.n191 VSUBS 0.019904f
C229 B.n192 VSUBS 0.020737f
C230 B.n193 VSUBS 0.007987f
C231 B.n194 VSUBS 0.007987f
C232 B.n195 VSUBS 0.007987f
C233 B.n196 VSUBS 0.007987f
C234 B.n197 VSUBS 0.007987f
C235 B.n198 VSUBS 0.007987f
C236 B.n199 VSUBS 0.007987f
C237 B.n200 VSUBS 0.007987f
C238 B.n201 VSUBS 0.007987f
C239 B.n202 VSUBS 0.007987f
C240 B.n203 VSUBS 0.007987f
C241 B.n204 VSUBS 0.007987f
C242 B.n205 VSUBS 0.007987f
C243 B.n206 VSUBS 0.007987f
C244 B.n207 VSUBS 0.007987f
C245 B.n208 VSUBS 0.007987f
C246 B.n209 VSUBS 0.007987f
C247 B.n210 VSUBS 0.007987f
C248 B.n211 VSUBS 0.007987f
C249 B.n212 VSUBS 0.007987f
C250 B.n213 VSUBS 0.007987f
C251 B.n214 VSUBS 0.007987f
C252 B.n215 VSUBS 0.007987f
C253 B.n216 VSUBS 0.007987f
C254 B.n217 VSUBS 0.007987f
C255 B.n218 VSUBS 0.007987f
C256 B.n219 VSUBS 0.007987f
C257 B.n220 VSUBS 0.007987f
C258 B.n221 VSUBS 0.007987f
C259 B.n222 VSUBS 0.007987f
C260 B.n223 VSUBS 0.007987f
C261 B.n224 VSUBS 0.007987f
C262 B.n225 VSUBS 0.007987f
C263 B.n226 VSUBS 0.007987f
C264 B.n227 VSUBS 0.007987f
C265 B.n228 VSUBS 0.007987f
C266 B.n229 VSUBS 0.007987f
C267 B.n230 VSUBS 0.007987f
C268 B.n231 VSUBS 0.007987f
C269 B.n232 VSUBS 0.007987f
C270 B.n233 VSUBS 0.007987f
C271 B.n234 VSUBS 0.007987f
C272 B.n235 VSUBS 0.007987f
C273 B.n236 VSUBS 0.007987f
C274 B.n237 VSUBS 0.007987f
C275 B.n238 VSUBS 0.007987f
C276 B.n239 VSUBS 0.007987f
C277 B.n240 VSUBS 0.007987f
C278 B.n241 VSUBS 0.007987f
C279 B.n242 VSUBS 0.007987f
C280 B.n243 VSUBS 0.007987f
C281 B.t11 VSUBS 0.373356f
C282 B.t10 VSUBS 0.386595f
C283 B.t9 VSUBS 0.575948f
C284 B.n244 VSUBS 0.162629f
C285 B.n245 VSUBS 0.07486f
C286 B.n246 VSUBS 0.018506f
C287 B.n247 VSUBS 0.007517f
C288 B.n248 VSUBS 0.007987f
C289 B.n249 VSUBS 0.007987f
C290 B.n250 VSUBS 0.007987f
C291 B.n251 VSUBS 0.007987f
C292 B.n252 VSUBS 0.007987f
C293 B.n253 VSUBS 0.007987f
C294 B.n254 VSUBS 0.007987f
C295 B.n255 VSUBS 0.007987f
C296 B.n256 VSUBS 0.007987f
C297 B.n257 VSUBS 0.007987f
C298 B.n258 VSUBS 0.007987f
C299 B.n259 VSUBS 0.007987f
C300 B.n260 VSUBS 0.007987f
C301 B.n261 VSUBS 0.007987f
C302 B.n262 VSUBS 0.007987f
C303 B.n263 VSUBS 0.004463f
C304 B.n264 VSUBS 0.018506f
C305 B.n265 VSUBS 0.007517f
C306 B.n266 VSUBS 0.007987f
C307 B.n267 VSUBS 0.007987f
C308 B.n268 VSUBS 0.007987f
C309 B.n269 VSUBS 0.007987f
C310 B.n270 VSUBS 0.007987f
C311 B.n271 VSUBS 0.007987f
C312 B.n272 VSUBS 0.007987f
C313 B.n273 VSUBS 0.007987f
C314 B.n274 VSUBS 0.007987f
C315 B.n275 VSUBS 0.007987f
C316 B.n276 VSUBS 0.007987f
C317 B.n277 VSUBS 0.007987f
C318 B.n278 VSUBS 0.007987f
C319 B.n279 VSUBS 0.007987f
C320 B.n280 VSUBS 0.007987f
C321 B.n281 VSUBS 0.007987f
C322 B.n282 VSUBS 0.007987f
C323 B.n283 VSUBS 0.007987f
C324 B.n284 VSUBS 0.007987f
C325 B.n285 VSUBS 0.007987f
C326 B.n286 VSUBS 0.007987f
C327 B.n287 VSUBS 0.007987f
C328 B.n288 VSUBS 0.007987f
C329 B.n289 VSUBS 0.007987f
C330 B.n290 VSUBS 0.007987f
C331 B.n291 VSUBS 0.007987f
C332 B.n292 VSUBS 0.007987f
C333 B.n293 VSUBS 0.007987f
C334 B.n294 VSUBS 0.007987f
C335 B.n295 VSUBS 0.007987f
C336 B.n296 VSUBS 0.007987f
C337 B.n297 VSUBS 0.007987f
C338 B.n298 VSUBS 0.007987f
C339 B.n299 VSUBS 0.007987f
C340 B.n300 VSUBS 0.007987f
C341 B.n301 VSUBS 0.007987f
C342 B.n302 VSUBS 0.007987f
C343 B.n303 VSUBS 0.007987f
C344 B.n304 VSUBS 0.007987f
C345 B.n305 VSUBS 0.007987f
C346 B.n306 VSUBS 0.007987f
C347 B.n307 VSUBS 0.007987f
C348 B.n308 VSUBS 0.007987f
C349 B.n309 VSUBS 0.007987f
C350 B.n310 VSUBS 0.007987f
C351 B.n311 VSUBS 0.007987f
C352 B.n312 VSUBS 0.007987f
C353 B.n313 VSUBS 0.007987f
C354 B.n314 VSUBS 0.007987f
C355 B.n315 VSUBS 0.007987f
C356 B.n316 VSUBS 0.007987f
C357 B.n317 VSUBS 0.020737f
C358 B.n318 VSUBS 0.019904f
C359 B.n319 VSUBS 0.020737f
C360 B.n320 VSUBS 0.007987f
C361 B.n321 VSUBS 0.007987f
C362 B.n322 VSUBS 0.007987f
C363 B.n323 VSUBS 0.007987f
C364 B.n324 VSUBS 0.007987f
C365 B.n325 VSUBS 0.007987f
C366 B.n326 VSUBS 0.007987f
C367 B.n327 VSUBS 0.007987f
C368 B.n328 VSUBS 0.007987f
C369 B.n329 VSUBS 0.007987f
C370 B.n330 VSUBS 0.007987f
C371 B.n331 VSUBS 0.007987f
C372 B.n332 VSUBS 0.007987f
C373 B.n333 VSUBS 0.007987f
C374 B.n334 VSUBS 0.007987f
C375 B.n335 VSUBS 0.007987f
C376 B.n336 VSUBS 0.007987f
C377 B.n337 VSUBS 0.007987f
C378 B.n338 VSUBS 0.007987f
C379 B.n339 VSUBS 0.007987f
C380 B.n340 VSUBS 0.007987f
C381 B.n341 VSUBS 0.007987f
C382 B.n342 VSUBS 0.007987f
C383 B.n343 VSUBS 0.007987f
C384 B.n344 VSUBS 0.007987f
C385 B.n345 VSUBS 0.007987f
C386 B.n346 VSUBS 0.007987f
C387 B.n347 VSUBS 0.007987f
C388 B.n348 VSUBS 0.007987f
C389 B.n349 VSUBS 0.007987f
C390 B.n350 VSUBS 0.007987f
C391 B.n351 VSUBS 0.007987f
C392 B.n352 VSUBS 0.007987f
C393 B.n353 VSUBS 0.007987f
C394 B.n354 VSUBS 0.007987f
C395 B.n355 VSUBS 0.007987f
C396 B.n356 VSUBS 0.007987f
C397 B.n357 VSUBS 0.007987f
C398 B.n358 VSUBS 0.007987f
C399 B.n359 VSUBS 0.007987f
C400 B.n360 VSUBS 0.007987f
C401 B.n361 VSUBS 0.007987f
C402 B.n362 VSUBS 0.007987f
C403 B.n363 VSUBS 0.007987f
C404 B.n364 VSUBS 0.007987f
C405 B.n365 VSUBS 0.007987f
C406 B.n366 VSUBS 0.007987f
C407 B.n367 VSUBS 0.007987f
C408 B.n368 VSUBS 0.007987f
C409 B.n369 VSUBS 0.007987f
C410 B.n370 VSUBS 0.007987f
C411 B.n371 VSUBS 0.007987f
C412 B.n372 VSUBS 0.007987f
C413 B.n373 VSUBS 0.007987f
C414 B.n374 VSUBS 0.007987f
C415 B.n375 VSUBS 0.007987f
C416 B.n376 VSUBS 0.007987f
C417 B.n377 VSUBS 0.007987f
C418 B.n378 VSUBS 0.007987f
C419 B.n379 VSUBS 0.007987f
C420 B.n380 VSUBS 0.007987f
C421 B.n381 VSUBS 0.007987f
C422 B.n382 VSUBS 0.007987f
C423 B.n383 VSUBS 0.007987f
C424 B.n384 VSUBS 0.007987f
C425 B.n385 VSUBS 0.007987f
C426 B.n386 VSUBS 0.007987f
C427 B.n387 VSUBS 0.007987f
C428 B.n388 VSUBS 0.007987f
C429 B.n389 VSUBS 0.007987f
C430 B.n390 VSUBS 0.007987f
C431 B.n391 VSUBS 0.007987f
C432 B.n392 VSUBS 0.007987f
C433 B.n393 VSUBS 0.007987f
C434 B.n394 VSUBS 0.007987f
C435 B.n395 VSUBS 0.007987f
C436 B.n396 VSUBS 0.007987f
C437 B.n397 VSUBS 0.007987f
C438 B.n398 VSUBS 0.007987f
C439 B.n399 VSUBS 0.007987f
C440 B.n400 VSUBS 0.007987f
C441 B.n401 VSUBS 0.007987f
C442 B.n402 VSUBS 0.007987f
C443 B.n403 VSUBS 0.007987f
C444 B.n404 VSUBS 0.007987f
C445 B.n405 VSUBS 0.007987f
C446 B.n406 VSUBS 0.007987f
C447 B.n407 VSUBS 0.019904f
C448 B.n408 VSUBS 0.019904f
C449 B.n409 VSUBS 0.020737f
C450 B.n410 VSUBS 0.007987f
C451 B.n411 VSUBS 0.007987f
C452 B.n412 VSUBS 0.007987f
C453 B.n413 VSUBS 0.007987f
C454 B.n414 VSUBS 0.007987f
C455 B.n415 VSUBS 0.007987f
C456 B.n416 VSUBS 0.007987f
C457 B.n417 VSUBS 0.007987f
C458 B.n418 VSUBS 0.007987f
C459 B.n419 VSUBS 0.007987f
C460 B.n420 VSUBS 0.007987f
C461 B.n421 VSUBS 0.007987f
C462 B.n422 VSUBS 0.007987f
C463 B.n423 VSUBS 0.007987f
C464 B.n424 VSUBS 0.007987f
C465 B.n425 VSUBS 0.007987f
C466 B.n426 VSUBS 0.007987f
C467 B.n427 VSUBS 0.007987f
C468 B.n428 VSUBS 0.007987f
C469 B.n429 VSUBS 0.007987f
C470 B.n430 VSUBS 0.007987f
C471 B.n431 VSUBS 0.007987f
C472 B.n432 VSUBS 0.007987f
C473 B.n433 VSUBS 0.007987f
C474 B.n434 VSUBS 0.007987f
C475 B.n435 VSUBS 0.007987f
C476 B.n436 VSUBS 0.007987f
C477 B.n437 VSUBS 0.007987f
C478 B.n438 VSUBS 0.007987f
C479 B.n439 VSUBS 0.007987f
C480 B.n440 VSUBS 0.007987f
C481 B.n441 VSUBS 0.007987f
C482 B.n442 VSUBS 0.007987f
C483 B.n443 VSUBS 0.007987f
C484 B.n444 VSUBS 0.007987f
C485 B.n445 VSUBS 0.007987f
C486 B.n446 VSUBS 0.007987f
C487 B.n447 VSUBS 0.007987f
C488 B.n448 VSUBS 0.007987f
C489 B.n449 VSUBS 0.007987f
C490 B.n450 VSUBS 0.007987f
C491 B.n451 VSUBS 0.007987f
C492 B.n452 VSUBS 0.007987f
C493 B.n453 VSUBS 0.007987f
C494 B.n454 VSUBS 0.007987f
C495 B.n455 VSUBS 0.007987f
C496 B.n456 VSUBS 0.007987f
C497 B.n457 VSUBS 0.007987f
C498 B.n458 VSUBS 0.007987f
C499 B.n459 VSUBS 0.007987f
C500 B.n460 VSUBS 0.007987f
C501 B.n461 VSUBS 0.007987f
C502 B.n462 VSUBS 0.007517f
C503 B.n463 VSUBS 0.018506f
C504 B.n464 VSUBS 0.004463f
C505 B.n465 VSUBS 0.007987f
C506 B.n466 VSUBS 0.007987f
C507 B.n467 VSUBS 0.007987f
C508 B.n468 VSUBS 0.007987f
C509 B.n469 VSUBS 0.007987f
C510 B.n470 VSUBS 0.007987f
C511 B.n471 VSUBS 0.007987f
C512 B.n472 VSUBS 0.007987f
C513 B.n473 VSUBS 0.007987f
C514 B.n474 VSUBS 0.007987f
C515 B.n475 VSUBS 0.007987f
C516 B.n476 VSUBS 0.007987f
C517 B.n477 VSUBS 0.004463f
C518 B.n478 VSUBS 0.007987f
C519 B.n479 VSUBS 0.007987f
C520 B.n480 VSUBS 0.007987f
C521 B.n481 VSUBS 0.007987f
C522 B.n482 VSUBS 0.007987f
C523 B.n483 VSUBS 0.007987f
C524 B.n484 VSUBS 0.007987f
C525 B.n485 VSUBS 0.007987f
C526 B.n486 VSUBS 0.007987f
C527 B.n487 VSUBS 0.007987f
C528 B.n488 VSUBS 0.007987f
C529 B.n489 VSUBS 0.007987f
C530 B.n490 VSUBS 0.007987f
C531 B.n491 VSUBS 0.007987f
C532 B.n492 VSUBS 0.007987f
C533 B.n493 VSUBS 0.007987f
C534 B.n494 VSUBS 0.007987f
C535 B.n495 VSUBS 0.007987f
C536 B.n496 VSUBS 0.007987f
C537 B.n497 VSUBS 0.007987f
C538 B.n498 VSUBS 0.007987f
C539 B.n499 VSUBS 0.007987f
C540 B.n500 VSUBS 0.007987f
C541 B.n501 VSUBS 0.007987f
C542 B.n502 VSUBS 0.007987f
C543 B.n503 VSUBS 0.007987f
C544 B.n504 VSUBS 0.007987f
C545 B.n505 VSUBS 0.007987f
C546 B.n506 VSUBS 0.007987f
C547 B.n507 VSUBS 0.007987f
C548 B.n508 VSUBS 0.007987f
C549 B.n509 VSUBS 0.007987f
C550 B.n510 VSUBS 0.007987f
C551 B.n511 VSUBS 0.007987f
C552 B.n512 VSUBS 0.007987f
C553 B.n513 VSUBS 0.007987f
C554 B.n514 VSUBS 0.007987f
C555 B.n515 VSUBS 0.007987f
C556 B.n516 VSUBS 0.007987f
C557 B.n517 VSUBS 0.007987f
C558 B.n518 VSUBS 0.007987f
C559 B.n519 VSUBS 0.007987f
C560 B.n520 VSUBS 0.007987f
C561 B.n521 VSUBS 0.007987f
C562 B.n522 VSUBS 0.007987f
C563 B.n523 VSUBS 0.007987f
C564 B.n524 VSUBS 0.007987f
C565 B.n525 VSUBS 0.007987f
C566 B.n526 VSUBS 0.007987f
C567 B.n527 VSUBS 0.007987f
C568 B.n528 VSUBS 0.007987f
C569 B.n529 VSUBS 0.007987f
C570 B.n530 VSUBS 0.007987f
C571 B.n531 VSUBS 0.020737f
C572 B.n532 VSUBS 0.020737f
C573 B.n533 VSUBS 0.019904f
C574 B.n534 VSUBS 0.007987f
C575 B.n535 VSUBS 0.007987f
C576 B.n536 VSUBS 0.007987f
C577 B.n537 VSUBS 0.007987f
C578 B.n538 VSUBS 0.007987f
C579 B.n539 VSUBS 0.007987f
C580 B.n540 VSUBS 0.007987f
C581 B.n541 VSUBS 0.007987f
C582 B.n542 VSUBS 0.007987f
C583 B.n543 VSUBS 0.007987f
C584 B.n544 VSUBS 0.007987f
C585 B.n545 VSUBS 0.007987f
C586 B.n546 VSUBS 0.007987f
C587 B.n547 VSUBS 0.007987f
C588 B.n548 VSUBS 0.007987f
C589 B.n549 VSUBS 0.007987f
C590 B.n550 VSUBS 0.007987f
C591 B.n551 VSUBS 0.007987f
C592 B.n552 VSUBS 0.007987f
C593 B.n553 VSUBS 0.007987f
C594 B.n554 VSUBS 0.007987f
C595 B.n555 VSUBS 0.007987f
C596 B.n556 VSUBS 0.007987f
C597 B.n557 VSUBS 0.007987f
C598 B.n558 VSUBS 0.007987f
C599 B.n559 VSUBS 0.007987f
C600 B.n560 VSUBS 0.007987f
C601 B.n561 VSUBS 0.007987f
C602 B.n562 VSUBS 0.007987f
C603 B.n563 VSUBS 0.007987f
C604 B.n564 VSUBS 0.007987f
C605 B.n565 VSUBS 0.007987f
C606 B.n566 VSUBS 0.007987f
C607 B.n567 VSUBS 0.007987f
C608 B.n568 VSUBS 0.007987f
C609 B.n569 VSUBS 0.007987f
C610 B.n570 VSUBS 0.007987f
C611 B.n571 VSUBS 0.007987f
C612 B.n572 VSUBS 0.007987f
C613 B.n573 VSUBS 0.007987f
C614 B.n574 VSUBS 0.007987f
C615 B.n575 VSUBS 0.010423f
C616 B.n576 VSUBS 0.011103f
C617 B.n577 VSUBS 0.022079f
C618 VDD1.t5 VSUBS 0.207442f
C619 VDD1.t3 VSUBS 0.207442f
C620 VDD1.n0 VSUBS 1.57307f
C621 VDD1.t4 VSUBS 0.207442f
C622 VDD1.t7 VSUBS 0.207442f
C623 VDD1.n1 VSUBS 1.57204f
C624 VDD1.t6 VSUBS 0.207442f
C625 VDD1.t0 VSUBS 0.207442f
C626 VDD1.n2 VSUBS 1.57204f
C627 VDD1.n3 VSUBS 2.95507f
C628 VDD1.t1 VSUBS 0.207442f
C629 VDD1.t2 VSUBS 0.207442f
C630 VDD1.n4 VSUBS 1.56715f
C631 VDD1.n5 VSUBS 2.65793f
C632 VP.n0 VSUBS 0.06185f
C633 VP.t1 VSUBS 1.46554f
C634 VP.n1 VSUBS 0.547614f
C635 VP.n2 VSUBS 0.046352f
C636 VP.t0 VSUBS 1.46554f
C637 VP.n3 VSUBS 0.0618f
C638 VP.n4 VSUBS 0.06185f
C639 VP.t5 VSUBS 1.5465f
C640 VP.t6 VSUBS 1.46554f
C641 VP.n5 VSUBS 0.547614f
C642 VP.n6 VSUBS 0.245145f
C643 VP.t4 VSUBS 1.46554f
C644 VP.t2 VSUBS 1.60073f
C645 VP.n7 VSUBS 0.609477f
C646 VP.n8 VSUBS 0.623905f
C647 VP.n9 VSUBS 0.066383f
C648 VP.n10 VSUBS 0.066383f
C649 VP.n11 VSUBS 0.046352f
C650 VP.n12 VSUBS 0.046352f
C651 VP.n13 VSUBS 0.045015f
C652 VP.n14 VSUBS 0.0618f
C653 VP.n15 VSUBS 0.630852f
C654 VP.n16 VSUBS 2.00116f
C655 VP.t3 VSUBS 1.5465f
C656 VP.n17 VSUBS 0.630852f
C657 VP.n18 VSUBS 2.03996f
C658 VP.n19 VSUBS 0.06185f
C659 VP.n20 VSUBS 0.046352f
C660 VP.n21 VSUBS 0.045015f
C661 VP.n22 VSUBS 0.547614f
C662 VP.n23 VSUBS 0.066383f
C663 VP.n24 VSUBS 0.066383f
C664 VP.n25 VSUBS 0.046352f
C665 VP.n26 VSUBS 0.046352f
C666 VP.n27 VSUBS 0.045015f
C667 VP.n28 VSUBS 0.0618f
C668 VP.t7 VSUBS 1.5465f
C669 VP.n29 VSUBS 0.630852f
C670 VP.n30 VSUBS 0.04341f
C671 VTAIL.t11 VSUBS 0.200685f
C672 VTAIL.t14 VSUBS 0.200685f
C673 VTAIL.n0 VSUBS 1.38626f
C674 VTAIL.n1 VSUBS 0.658737f
C675 VTAIL.t15 VSUBS 1.84364f
C676 VTAIL.n2 VSUBS 0.781602f
C677 VTAIL.t1 VSUBS 1.84364f
C678 VTAIL.n3 VSUBS 0.781602f
C679 VTAIL.t0 VSUBS 0.200685f
C680 VTAIL.t5 VSUBS 0.200685f
C681 VTAIL.n4 VSUBS 1.38626f
C682 VTAIL.n5 VSUBS 0.75545f
C683 VTAIL.t4 VSUBS 1.84364f
C684 VTAIL.n6 VSUBS 1.88804f
C685 VTAIL.t9 VSUBS 1.84365f
C686 VTAIL.n7 VSUBS 1.88803f
C687 VTAIL.t10 VSUBS 0.200685f
C688 VTAIL.t12 VSUBS 0.200685f
C689 VTAIL.n8 VSUBS 1.38626f
C690 VTAIL.n9 VSUBS 0.755444f
C691 VTAIL.t13 VSUBS 1.84365f
C692 VTAIL.n10 VSUBS 0.781596f
C693 VTAIL.t6 VSUBS 1.84365f
C694 VTAIL.n11 VSUBS 0.781596f
C695 VTAIL.t7 VSUBS 0.200685f
C696 VTAIL.t2 VSUBS 0.200685f
C697 VTAIL.n12 VSUBS 1.38626f
C698 VTAIL.n13 VSUBS 0.755444f
C699 VTAIL.t3 VSUBS 1.84364f
C700 VTAIL.n14 VSUBS 1.88804f
C701 VTAIL.t8 VSUBS 1.84364f
C702 VTAIL.n15 VSUBS 1.88339f
C703 VDD2.t0 VSUBS 0.205905f
C704 VDD2.t3 VSUBS 0.205905f
C705 VDD2.n0 VSUBS 1.56039f
C706 VDD2.t5 VSUBS 0.205905f
C707 VDD2.t1 VSUBS 0.205905f
C708 VDD2.n1 VSUBS 1.56039f
C709 VDD2.n2 VSUBS 2.87909f
C710 VDD2.t4 VSUBS 0.205905f
C711 VDD2.t7 VSUBS 0.205905f
C712 VDD2.n3 VSUBS 1.55555f
C713 VDD2.n4 VSUBS 2.60781f
C714 VDD2.t6 VSUBS 0.205905f
C715 VDD2.t2 VSUBS 0.205905f
C716 VDD2.n5 VSUBS 1.56036f
C717 VN.n0 VSUBS 0.060287f
C718 VN.t1 VSUBS 1.42851f
C719 VN.n1 VSUBS 0.533776f
C720 VN.n2 VSUBS 0.23895f
C721 VN.t4 VSUBS 1.42851f
C722 VN.t0 VSUBS 1.56028f
C723 VN.n3 VSUBS 0.594076f
C724 VN.n4 VSUBS 0.608139f
C725 VN.n5 VSUBS 0.064706f
C726 VN.n6 VSUBS 0.064706f
C727 VN.n7 VSUBS 0.04518f
C728 VN.n8 VSUBS 0.04518f
C729 VN.n9 VSUBS 0.043877f
C730 VN.n10 VSUBS 0.060239f
C731 VN.t7 VSUBS 1.50742f
C732 VN.n11 VSUBS 0.614911f
C733 VN.n12 VSUBS 0.042313f
C734 VN.n13 VSUBS 0.060287f
C735 VN.t5 VSUBS 1.42851f
C736 VN.n14 VSUBS 0.533776f
C737 VN.n15 VSUBS 0.23895f
C738 VN.t3 VSUBS 1.42851f
C739 VN.t2 VSUBS 1.56028f
C740 VN.n16 VSUBS 0.594076f
C741 VN.n17 VSUBS 0.608139f
C742 VN.n18 VSUBS 0.064706f
C743 VN.n19 VSUBS 0.064706f
C744 VN.n20 VSUBS 0.04518f
C745 VN.n21 VSUBS 0.04518f
C746 VN.n22 VSUBS 0.043877f
C747 VN.n23 VSUBS 0.060239f
C748 VN.t6 VSUBS 1.50742f
C749 VN.n24 VSUBS 0.614911f
C750 VN.n25 VSUBS 1.97584f
.ends

