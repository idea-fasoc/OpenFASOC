* NGSPICE file created from diff_pair_sample_0371.ext - technology: sky130A

.subckt diff_pair_sample_0371 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=2.13675 ps=13.28 w=12.95 l=1.19
X1 VDD1.t0 VP.t1 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.13675 pd=13.28 as=5.0505 ps=26.68 w=12.95 l=1.19
X2 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=2.13675 ps=13.28 w=12.95 l=1.19
X3 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=2.13675 ps=13.28 w=12.95 l=1.19
X4 VDD1.t1 VP.t2 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.13675 pd=13.28 as=5.0505 ps=26.68 w=12.95 l=1.19
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=0 ps=0 w=12.95 l=1.19
X6 VTAIL.t3 VP.t3 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=2.13675 ps=13.28 w=12.95 l=1.19
X7 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=0 ps=0 w=12.95 l=1.19
X8 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.13675 pd=13.28 as=5.0505 ps=26.68 w=12.95 l=1.19
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=0 ps=0 w=12.95 l=1.19
X10 VDD2.t0 VN.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.13675 pd=13.28 as=5.0505 ps=26.68 w=12.95 l=1.19
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.0505 pd=26.68 as=0 ps=0 w=12.95 l=1.19
R0 VP.n2 VP.t3 298.18
R1 VP.n2 VP.t1 297.961
R2 VP.n3 VP.t0 262.265
R3 VP.n9 VP.t2 262.265
R4 VP.n4 VP.n3 173.044
R5 VP.n10 VP.n9 173.044
R6 VP.n8 VP.n0 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n5 VP.n1 161.3
R9 VP.n4 VP.n2 61.1175
R10 VP.n7 VP.n1 40.4934
R11 VP.n8 VP.n7 40.4934
R12 VP.n3 VP.n1 12.7233
R13 VP.n9 VP.n8 12.7233
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 102.644
R20 VDD1 VDD1.n0 63.3673
R21 VDD1.n0 VDD1.t3 1.52946
R22 VDD1.n0 VDD1.t0 1.52946
R23 VDD1.n1 VDD1.t2 1.52946
R24 VDD1.n1 VDD1.t1 1.52946
R25 VTAIL.n5 VTAIL.t3 48.1604
R26 VTAIL.n4 VTAIL.t0 48.1604
R27 VTAIL.n3 VTAIL.t2 48.1604
R28 VTAIL.n7 VTAIL.t7 48.1593
R29 VTAIL.n0 VTAIL.t1 48.1593
R30 VTAIL.n1 VTAIL.t4 48.1593
R31 VTAIL.n2 VTAIL.t6 48.1593
R32 VTAIL.n6 VTAIL.t5 48.1593
R33 VTAIL.n7 VTAIL.n6 24.841
R34 VTAIL.n3 VTAIL.n2 24.841
R35 VTAIL.n4 VTAIL.n3 1.31084
R36 VTAIL.n6 VTAIL.n5 1.31084
R37 VTAIL.n2 VTAIL.n1 1.31084
R38 VTAIL VTAIL.n0 0.713862
R39 VTAIL VTAIL.n7 0.597483
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 B.n674 B.n673 585
R43 B.n289 B.n90 585
R44 B.n288 B.n287 585
R45 B.n286 B.n285 585
R46 B.n284 B.n283 585
R47 B.n282 B.n281 585
R48 B.n280 B.n279 585
R49 B.n278 B.n277 585
R50 B.n276 B.n275 585
R51 B.n274 B.n273 585
R52 B.n272 B.n271 585
R53 B.n270 B.n269 585
R54 B.n268 B.n267 585
R55 B.n266 B.n265 585
R56 B.n264 B.n263 585
R57 B.n262 B.n261 585
R58 B.n260 B.n259 585
R59 B.n258 B.n257 585
R60 B.n256 B.n255 585
R61 B.n254 B.n253 585
R62 B.n252 B.n251 585
R63 B.n250 B.n249 585
R64 B.n248 B.n247 585
R65 B.n246 B.n245 585
R66 B.n244 B.n243 585
R67 B.n242 B.n241 585
R68 B.n240 B.n239 585
R69 B.n238 B.n237 585
R70 B.n236 B.n235 585
R71 B.n234 B.n233 585
R72 B.n232 B.n231 585
R73 B.n230 B.n229 585
R74 B.n228 B.n227 585
R75 B.n226 B.n225 585
R76 B.n224 B.n223 585
R77 B.n222 B.n221 585
R78 B.n220 B.n219 585
R79 B.n218 B.n217 585
R80 B.n216 B.n215 585
R81 B.n214 B.n213 585
R82 B.n212 B.n211 585
R83 B.n210 B.n209 585
R84 B.n208 B.n207 585
R85 B.n206 B.n205 585
R86 B.n204 B.n203 585
R87 B.n202 B.n201 585
R88 B.n200 B.n199 585
R89 B.n198 B.n197 585
R90 B.n196 B.n195 585
R91 B.n194 B.n193 585
R92 B.n192 B.n191 585
R93 B.n190 B.n189 585
R94 B.n188 B.n187 585
R95 B.n186 B.n185 585
R96 B.n184 B.n183 585
R97 B.n182 B.n181 585
R98 B.n180 B.n179 585
R99 B.n178 B.n177 585
R100 B.n176 B.n175 585
R101 B.n174 B.n173 585
R102 B.n172 B.n171 585
R103 B.n170 B.n169 585
R104 B.n168 B.n167 585
R105 B.n166 B.n165 585
R106 B.n164 B.n163 585
R107 B.n162 B.n161 585
R108 B.n160 B.n159 585
R109 B.n158 B.n157 585
R110 B.n156 B.n155 585
R111 B.n154 B.n153 585
R112 B.n152 B.n151 585
R113 B.n150 B.n149 585
R114 B.n148 B.n147 585
R115 B.n146 B.n145 585
R116 B.n144 B.n143 585
R117 B.n142 B.n141 585
R118 B.n140 B.n139 585
R119 B.n138 B.n137 585
R120 B.n136 B.n135 585
R121 B.n134 B.n133 585
R122 B.n132 B.n131 585
R123 B.n130 B.n129 585
R124 B.n128 B.n127 585
R125 B.n126 B.n125 585
R126 B.n124 B.n123 585
R127 B.n122 B.n121 585
R128 B.n120 B.n119 585
R129 B.n118 B.n117 585
R130 B.n116 B.n115 585
R131 B.n114 B.n113 585
R132 B.n112 B.n111 585
R133 B.n110 B.n109 585
R134 B.n108 B.n107 585
R135 B.n106 B.n105 585
R136 B.n104 B.n103 585
R137 B.n102 B.n101 585
R138 B.n100 B.n99 585
R139 B.n98 B.n97 585
R140 B.n672 B.n41 585
R141 B.n677 B.n41 585
R142 B.n671 B.n40 585
R143 B.n678 B.n40 585
R144 B.n670 B.n669 585
R145 B.n669 B.n36 585
R146 B.n668 B.n35 585
R147 B.n684 B.n35 585
R148 B.n667 B.n34 585
R149 B.n685 B.n34 585
R150 B.n666 B.n33 585
R151 B.n686 B.n33 585
R152 B.n665 B.n664 585
R153 B.n664 B.n29 585
R154 B.n663 B.n28 585
R155 B.n692 B.n28 585
R156 B.n662 B.n27 585
R157 B.n693 B.n27 585
R158 B.n661 B.n26 585
R159 B.n694 B.n26 585
R160 B.n660 B.n659 585
R161 B.n659 B.n22 585
R162 B.n658 B.n21 585
R163 B.n700 B.n21 585
R164 B.n657 B.n20 585
R165 B.n701 B.n20 585
R166 B.n656 B.n19 585
R167 B.n702 B.n19 585
R168 B.n655 B.n654 585
R169 B.n654 B.n15 585
R170 B.n653 B.n14 585
R171 B.n708 B.n14 585
R172 B.n652 B.n13 585
R173 B.n709 B.n13 585
R174 B.n651 B.n12 585
R175 B.n710 B.n12 585
R176 B.n650 B.n649 585
R177 B.n649 B.n648 585
R178 B.n647 B.n646 585
R179 B.n647 B.n8 585
R180 B.n645 B.n7 585
R181 B.n717 B.n7 585
R182 B.n644 B.n6 585
R183 B.n718 B.n6 585
R184 B.n643 B.n5 585
R185 B.n719 B.n5 585
R186 B.n642 B.n641 585
R187 B.n641 B.n4 585
R188 B.n640 B.n290 585
R189 B.n640 B.n639 585
R190 B.n630 B.n291 585
R191 B.n292 B.n291 585
R192 B.n632 B.n631 585
R193 B.n633 B.n632 585
R194 B.n629 B.n297 585
R195 B.n297 B.n296 585
R196 B.n628 B.n627 585
R197 B.n627 B.n626 585
R198 B.n299 B.n298 585
R199 B.n300 B.n299 585
R200 B.n619 B.n618 585
R201 B.n620 B.n619 585
R202 B.n617 B.n305 585
R203 B.n305 B.n304 585
R204 B.n616 B.n615 585
R205 B.n615 B.n614 585
R206 B.n307 B.n306 585
R207 B.n308 B.n307 585
R208 B.n607 B.n606 585
R209 B.n608 B.n607 585
R210 B.n605 B.n313 585
R211 B.n313 B.n312 585
R212 B.n604 B.n603 585
R213 B.n603 B.n602 585
R214 B.n315 B.n314 585
R215 B.n316 B.n315 585
R216 B.n595 B.n594 585
R217 B.n596 B.n595 585
R218 B.n593 B.n321 585
R219 B.n321 B.n320 585
R220 B.n592 B.n591 585
R221 B.n591 B.n590 585
R222 B.n323 B.n322 585
R223 B.n324 B.n323 585
R224 B.n583 B.n582 585
R225 B.n584 B.n583 585
R226 B.n581 B.n329 585
R227 B.n329 B.n328 585
R228 B.n576 B.n575 585
R229 B.n574 B.n380 585
R230 B.n573 B.n379 585
R231 B.n578 B.n379 585
R232 B.n572 B.n571 585
R233 B.n570 B.n569 585
R234 B.n568 B.n567 585
R235 B.n566 B.n565 585
R236 B.n564 B.n563 585
R237 B.n562 B.n561 585
R238 B.n560 B.n559 585
R239 B.n558 B.n557 585
R240 B.n556 B.n555 585
R241 B.n554 B.n553 585
R242 B.n552 B.n551 585
R243 B.n550 B.n549 585
R244 B.n548 B.n547 585
R245 B.n546 B.n545 585
R246 B.n544 B.n543 585
R247 B.n542 B.n541 585
R248 B.n540 B.n539 585
R249 B.n538 B.n537 585
R250 B.n536 B.n535 585
R251 B.n534 B.n533 585
R252 B.n532 B.n531 585
R253 B.n530 B.n529 585
R254 B.n528 B.n527 585
R255 B.n526 B.n525 585
R256 B.n524 B.n523 585
R257 B.n522 B.n521 585
R258 B.n520 B.n519 585
R259 B.n518 B.n517 585
R260 B.n516 B.n515 585
R261 B.n514 B.n513 585
R262 B.n512 B.n511 585
R263 B.n510 B.n509 585
R264 B.n508 B.n507 585
R265 B.n506 B.n505 585
R266 B.n504 B.n503 585
R267 B.n502 B.n501 585
R268 B.n500 B.n499 585
R269 B.n498 B.n497 585
R270 B.n496 B.n495 585
R271 B.n494 B.n493 585
R272 B.n492 B.n491 585
R273 B.n489 B.n488 585
R274 B.n487 B.n486 585
R275 B.n485 B.n484 585
R276 B.n483 B.n482 585
R277 B.n481 B.n480 585
R278 B.n479 B.n478 585
R279 B.n477 B.n476 585
R280 B.n475 B.n474 585
R281 B.n473 B.n472 585
R282 B.n471 B.n470 585
R283 B.n468 B.n467 585
R284 B.n466 B.n465 585
R285 B.n464 B.n463 585
R286 B.n462 B.n461 585
R287 B.n460 B.n459 585
R288 B.n458 B.n457 585
R289 B.n456 B.n455 585
R290 B.n454 B.n453 585
R291 B.n452 B.n451 585
R292 B.n450 B.n449 585
R293 B.n448 B.n447 585
R294 B.n446 B.n445 585
R295 B.n444 B.n443 585
R296 B.n442 B.n441 585
R297 B.n440 B.n439 585
R298 B.n438 B.n437 585
R299 B.n436 B.n435 585
R300 B.n434 B.n433 585
R301 B.n432 B.n431 585
R302 B.n430 B.n429 585
R303 B.n428 B.n427 585
R304 B.n426 B.n425 585
R305 B.n424 B.n423 585
R306 B.n422 B.n421 585
R307 B.n420 B.n419 585
R308 B.n418 B.n417 585
R309 B.n416 B.n415 585
R310 B.n414 B.n413 585
R311 B.n412 B.n411 585
R312 B.n410 B.n409 585
R313 B.n408 B.n407 585
R314 B.n406 B.n405 585
R315 B.n404 B.n403 585
R316 B.n402 B.n401 585
R317 B.n400 B.n399 585
R318 B.n398 B.n397 585
R319 B.n396 B.n395 585
R320 B.n394 B.n393 585
R321 B.n392 B.n391 585
R322 B.n390 B.n389 585
R323 B.n388 B.n387 585
R324 B.n386 B.n385 585
R325 B.n331 B.n330 585
R326 B.n580 B.n579 585
R327 B.n579 B.n578 585
R328 B.n327 B.n326 585
R329 B.n328 B.n327 585
R330 B.n586 B.n585 585
R331 B.n585 B.n584 585
R332 B.n587 B.n325 585
R333 B.n325 B.n324 585
R334 B.n589 B.n588 585
R335 B.n590 B.n589 585
R336 B.n319 B.n318 585
R337 B.n320 B.n319 585
R338 B.n598 B.n597 585
R339 B.n597 B.n596 585
R340 B.n599 B.n317 585
R341 B.n317 B.n316 585
R342 B.n601 B.n600 585
R343 B.n602 B.n601 585
R344 B.n311 B.n310 585
R345 B.n312 B.n311 585
R346 B.n610 B.n609 585
R347 B.n609 B.n608 585
R348 B.n611 B.n309 585
R349 B.n309 B.n308 585
R350 B.n613 B.n612 585
R351 B.n614 B.n613 585
R352 B.n303 B.n302 585
R353 B.n304 B.n303 585
R354 B.n622 B.n621 585
R355 B.n621 B.n620 585
R356 B.n623 B.n301 585
R357 B.n301 B.n300 585
R358 B.n625 B.n624 585
R359 B.n626 B.n625 585
R360 B.n295 B.n294 585
R361 B.n296 B.n295 585
R362 B.n635 B.n634 585
R363 B.n634 B.n633 585
R364 B.n636 B.n293 585
R365 B.n293 B.n292 585
R366 B.n638 B.n637 585
R367 B.n639 B.n638 585
R368 B.n3 B.n0 585
R369 B.n4 B.n3 585
R370 B.n716 B.n1 585
R371 B.n717 B.n716 585
R372 B.n715 B.n714 585
R373 B.n715 B.n8 585
R374 B.n713 B.n9 585
R375 B.n648 B.n9 585
R376 B.n712 B.n711 585
R377 B.n711 B.n710 585
R378 B.n11 B.n10 585
R379 B.n709 B.n11 585
R380 B.n707 B.n706 585
R381 B.n708 B.n707 585
R382 B.n705 B.n16 585
R383 B.n16 B.n15 585
R384 B.n704 B.n703 585
R385 B.n703 B.n702 585
R386 B.n18 B.n17 585
R387 B.n701 B.n18 585
R388 B.n699 B.n698 585
R389 B.n700 B.n699 585
R390 B.n697 B.n23 585
R391 B.n23 B.n22 585
R392 B.n696 B.n695 585
R393 B.n695 B.n694 585
R394 B.n25 B.n24 585
R395 B.n693 B.n25 585
R396 B.n691 B.n690 585
R397 B.n692 B.n691 585
R398 B.n689 B.n30 585
R399 B.n30 B.n29 585
R400 B.n688 B.n687 585
R401 B.n687 B.n686 585
R402 B.n32 B.n31 585
R403 B.n685 B.n32 585
R404 B.n683 B.n682 585
R405 B.n684 B.n683 585
R406 B.n681 B.n37 585
R407 B.n37 B.n36 585
R408 B.n680 B.n679 585
R409 B.n679 B.n678 585
R410 B.n39 B.n38 585
R411 B.n677 B.n39 585
R412 B.n720 B.n719 585
R413 B.n718 B.n2 585
R414 B.n97 B.n39 535.745
R415 B.n674 B.n41 535.745
R416 B.n579 B.n329 535.745
R417 B.n576 B.n327 535.745
R418 B.n94 B.t4 466.329
R419 B.n91 B.t12 466.329
R420 B.n383 B.t15 466.329
R421 B.n381 B.t8 466.329
R422 B.n676 B.n675 256.663
R423 B.n676 B.n89 256.663
R424 B.n676 B.n88 256.663
R425 B.n676 B.n87 256.663
R426 B.n676 B.n86 256.663
R427 B.n676 B.n85 256.663
R428 B.n676 B.n84 256.663
R429 B.n676 B.n83 256.663
R430 B.n676 B.n82 256.663
R431 B.n676 B.n81 256.663
R432 B.n676 B.n80 256.663
R433 B.n676 B.n79 256.663
R434 B.n676 B.n78 256.663
R435 B.n676 B.n77 256.663
R436 B.n676 B.n76 256.663
R437 B.n676 B.n75 256.663
R438 B.n676 B.n74 256.663
R439 B.n676 B.n73 256.663
R440 B.n676 B.n72 256.663
R441 B.n676 B.n71 256.663
R442 B.n676 B.n70 256.663
R443 B.n676 B.n69 256.663
R444 B.n676 B.n68 256.663
R445 B.n676 B.n67 256.663
R446 B.n676 B.n66 256.663
R447 B.n676 B.n65 256.663
R448 B.n676 B.n64 256.663
R449 B.n676 B.n63 256.663
R450 B.n676 B.n62 256.663
R451 B.n676 B.n61 256.663
R452 B.n676 B.n60 256.663
R453 B.n676 B.n59 256.663
R454 B.n676 B.n58 256.663
R455 B.n676 B.n57 256.663
R456 B.n676 B.n56 256.663
R457 B.n676 B.n55 256.663
R458 B.n676 B.n54 256.663
R459 B.n676 B.n53 256.663
R460 B.n676 B.n52 256.663
R461 B.n676 B.n51 256.663
R462 B.n676 B.n50 256.663
R463 B.n676 B.n49 256.663
R464 B.n676 B.n48 256.663
R465 B.n676 B.n47 256.663
R466 B.n676 B.n46 256.663
R467 B.n676 B.n45 256.663
R468 B.n676 B.n44 256.663
R469 B.n676 B.n43 256.663
R470 B.n676 B.n42 256.663
R471 B.n578 B.n577 256.663
R472 B.n578 B.n332 256.663
R473 B.n578 B.n333 256.663
R474 B.n578 B.n334 256.663
R475 B.n578 B.n335 256.663
R476 B.n578 B.n336 256.663
R477 B.n578 B.n337 256.663
R478 B.n578 B.n338 256.663
R479 B.n578 B.n339 256.663
R480 B.n578 B.n340 256.663
R481 B.n578 B.n341 256.663
R482 B.n578 B.n342 256.663
R483 B.n578 B.n343 256.663
R484 B.n578 B.n344 256.663
R485 B.n578 B.n345 256.663
R486 B.n578 B.n346 256.663
R487 B.n578 B.n347 256.663
R488 B.n578 B.n348 256.663
R489 B.n578 B.n349 256.663
R490 B.n578 B.n350 256.663
R491 B.n578 B.n351 256.663
R492 B.n578 B.n352 256.663
R493 B.n578 B.n353 256.663
R494 B.n578 B.n354 256.663
R495 B.n578 B.n355 256.663
R496 B.n578 B.n356 256.663
R497 B.n578 B.n357 256.663
R498 B.n578 B.n358 256.663
R499 B.n578 B.n359 256.663
R500 B.n578 B.n360 256.663
R501 B.n578 B.n361 256.663
R502 B.n578 B.n362 256.663
R503 B.n578 B.n363 256.663
R504 B.n578 B.n364 256.663
R505 B.n578 B.n365 256.663
R506 B.n578 B.n366 256.663
R507 B.n578 B.n367 256.663
R508 B.n578 B.n368 256.663
R509 B.n578 B.n369 256.663
R510 B.n578 B.n370 256.663
R511 B.n578 B.n371 256.663
R512 B.n578 B.n372 256.663
R513 B.n578 B.n373 256.663
R514 B.n578 B.n374 256.663
R515 B.n578 B.n375 256.663
R516 B.n578 B.n376 256.663
R517 B.n578 B.n377 256.663
R518 B.n578 B.n378 256.663
R519 B.n722 B.n721 256.663
R520 B.n101 B.n100 163.367
R521 B.n105 B.n104 163.367
R522 B.n109 B.n108 163.367
R523 B.n113 B.n112 163.367
R524 B.n117 B.n116 163.367
R525 B.n121 B.n120 163.367
R526 B.n125 B.n124 163.367
R527 B.n129 B.n128 163.367
R528 B.n133 B.n132 163.367
R529 B.n137 B.n136 163.367
R530 B.n141 B.n140 163.367
R531 B.n145 B.n144 163.367
R532 B.n149 B.n148 163.367
R533 B.n153 B.n152 163.367
R534 B.n157 B.n156 163.367
R535 B.n161 B.n160 163.367
R536 B.n165 B.n164 163.367
R537 B.n169 B.n168 163.367
R538 B.n173 B.n172 163.367
R539 B.n177 B.n176 163.367
R540 B.n181 B.n180 163.367
R541 B.n185 B.n184 163.367
R542 B.n189 B.n188 163.367
R543 B.n193 B.n192 163.367
R544 B.n197 B.n196 163.367
R545 B.n201 B.n200 163.367
R546 B.n205 B.n204 163.367
R547 B.n209 B.n208 163.367
R548 B.n213 B.n212 163.367
R549 B.n217 B.n216 163.367
R550 B.n221 B.n220 163.367
R551 B.n225 B.n224 163.367
R552 B.n229 B.n228 163.367
R553 B.n233 B.n232 163.367
R554 B.n237 B.n236 163.367
R555 B.n241 B.n240 163.367
R556 B.n245 B.n244 163.367
R557 B.n249 B.n248 163.367
R558 B.n253 B.n252 163.367
R559 B.n257 B.n256 163.367
R560 B.n261 B.n260 163.367
R561 B.n265 B.n264 163.367
R562 B.n269 B.n268 163.367
R563 B.n273 B.n272 163.367
R564 B.n277 B.n276 163.367
R565 B.n281 B.n280 163.367
R566 B.n285 B.n284 163.367
R567 B.n287 B.n90 163.367
R568 B.n583 B.n329 163.367
R569 B.n583 B.n323 163.367
R570 B.n591 B.n323 163.367
R571 B.n591 B.n321 163.367
R572 B.n595 B.n321 163.367
R573 B.n595 B.n315 163.367
R574 B.n603 B.n315 163.367
R575 B.n603 B.n313 163.367
R576 B.n607 B.n313 163.367
R577 B.n607 B.n307 163.367
R578 B.n615 B.n307 163.367
R579 B.n615 B.n305 163.367
R580 B.n619 B.n305 163.367
R581 B.n619 B.n299 163.367
R582 B.n627 B.n299 163.367
R583 B.n627 B.n297 163.367
R584 B.n632 B.n297 163.367
R585 B.n632 B.n291 163.367
R586 B.n640 B.n291 163.367
R587 B.n641 B.n640 163.367
R588 B.n641 B.n5 163.367
R589 B.n6 B.n5 163.367
R590 B.n7 B.n6 163.367
R591 B.n647 B.n7 163.367
R592 B.n649 B.n647 163.367
R593 B.n649 B.n12 163.367
R594 B.n13 B.n12 163.367
R595 B.n14 B.n13 163.367
R596 B.n654 B.n14 163.367
R597 B.n654 B.n19 163.367
R598 B.n20 B.n19 163.367
R599 B.n21 B.n20 163.367
R600 B.n659 B.n21 163.367
R601 B.n659 B.n26 163.367
R602 B.n27 B.n26 163.367
R603 B.n28 B.n27 163.367
R604 B.n664 B.n28 163.367
R605 B.n664 B.n33 163.367
R606 B.n34 B.n33 163.367
R607 B.n35 B.n34 163.367
R608 B.n669 B.n35 163.367
R609 B.n669 B.n40 163.367
R610 B.n41 B.n40 163.367
R611 B.n380 B.n379 163.367
R612 B.n571 B.n379 163.367
R613 B.n569 B.n568 163.367
R614 B.n565 B.n564 163.367
R615 B.n561 B.n560 163.367
R616 B.n557 B.n556 163.367
R617 B.n553 B.n552 163.367
R618 B.n549 B.n548 163.367
R619 B.n545 B.n544 163.367
R620 B.n541 B.n540 163.367
R621 B.n537 B.n536 163.367
R622 B.n533 B.n532 163.367
R623 B.n529 B.n528 163.367
R624 B.n525 B.n524 163.367
R625 B.n521 B.n520 163.367
R626 B.n517 B.n516 163.367
R627 B.n513 B.n512 163.367
R628 B.n509 B.n508 163.367
R629 B.n505 B.n504 163.367
R630 B.n501 B.n500 163.367
R631 B.n497 B.n496 163.367
R632 B.n493 B.n492 163.367
R633 B.n488 B.n487 163.367
R634 B.n484 B.n483 163.367
R635 B.n480 B.n479 163.367
R636 B.n476 B.n475 163.367
R637 B.n472 B.n471 163.367
R638 B.n467 B.n466 163.367
R639 B.n463 B.n462 163.367
R640 B.n459 B.n458 163.367
R641 B.n455 B.n454 163.367
R642 B.n451 B.n450 163.367
R643 B.n447 B.n446 163.367
R644 B.n443 B.n442 163.367
R645 B.n439 B.n438 163.367
R646 B.n435 B.n434 163.367
R647 B.n431 B.n430 163.367
R648 B.n427 B.n426 163.367
R649 B.n423 B.n422 163.367
R650 B.n419 B.n418 163.367
R651 B.n415 B.n414 163.367
R652 B.n411 B.n410 163.367
R653 B.n407 B.n406 163.367
R654 B.n403 B.n402 163.367
R655 B.n399 B.n398 163.367
R656 B.n395 B.n394 163.367
R657 B.n391 B.n390 163.367
R658 B.n387 B.n386 163.367
R659 B.n579 B.n331 163.367
R660 B.n585 B.n327 163.367
R661 B.n585 B.n325 163.367
R662 B.n589 B.n325 163.367
R663 B.n589 B.n319 163.367
R664 B.n597 B.n319 163.367
R665 B.n597 B.n317 163.367
R666 B.n601 B.n317 163.367
R667 B.n601 B.n311 163.367
R668 B.n609 B.n311 163.367
R669 B.n609 B.n309 163.367
R670 B.n613 B.n309 163.367
R671 B.n613 B.n303 163.367
R672 B.n621 B.n303 163.367
R673 B.n621 B.n301 163.367
R674 B.n625 B.n301 163.367
R675 B.n625 B.n295 163.367
R676 B.n634 B.n295 163.367
R677 B.n634 B.n293 163.367
R678 B.n638 B.n293 163.367
R679 B.n638 B.n3 163.367
R680 B.n720 B.n3 163.367
R681 B.n716 B.n2 163.367
R682 B.n716 B.n715 163.367
R683 B.n715 B.n9 163.367
R684 B.n711 B.n9 163.367
R685 B.n711 B.n11 163.367
R686 B.n707 B.n11 163.367
R687 B.n707 B.n16 163.367
R688 B.n703 B.n16 163.367
R689 B.n703 B.n18 163.367
R690 B.n699 B.n18 163.367
R691 B.n699 B.n23 163.367
R692 B.n695 B.n23 163.367
R693 B.n695 B.n25 163.367
R694 B.n691 B.n25 163.367
R695 B.n691 B.n30 163.367
R696 B.n687 B.n30 163.367
R697 B.n687 B.n32 163.367
R698 B.n683 B.n32 163.367
R699 B.n683 B.n37 163.367
R700 B.n679 B.n37 163.367
R701 B.n679 B.n39 163.367
R702 B.n91 B.t13 97.731
R703 B.n383 B.t17 97.731
R704 B.n94 B.t6 97.7142
R705 B.n381 B.t11 97.7142
R706 B.n578 B.n328 75.4463
R707 B.n677 B.n676 75.4463
R708 B.n97 B.n42 71.676
R709 B.n101 B.n43 71.676
R710 B.n105 B.n44 71.676
R711 B.n109 B.n45 71.676
R712 B.n113 B.n46 71.676
R713 B.n117 B.n47 71.676
R714 B.n121 B.n48 71.676
R715 B.n125 B.n49 71.676
R716 B.n129 B.n50 71.676
R717 B.n133 B.n51 71.676
R718 B.n137 B.n52 71.676
R719 B.n141 B.n53 71.676
R720 B.n145 B.n54 71.676
R721 B.n149 B.n55 71.676
R722 B.n153 B.n56 71.676
R723 B.n157 B.n57 71.676
R724 B.n161 B.n58 71.676
R725 B.n165 B.n59 71.676
R726 B.n169 B.n60 71.676
R727 B.n173 B.n61 71.676
R728 B.n177 B.n62 71.676
R729 B.n181 B.n63 71.676
R730 B.n185 B.n64 71.676
R731 B.n189 B.n65 71.676
R732 B.n193 B.n66 71.676
R733 B.n197 B.n67 71.676
R734 B.n201 B.n68 71.676
R735 B.n205 B.n69 71.676
R736 B.n209 B.n70 71.676
R737 B.n213 B.n71 71.676
R738 B.n217 B.n72 71.676
R739 B.n221 B.n73 71.676
R740 B.n225 B.n74 71.676
R741 B.n229 B.n75 71.676
R742 B.n233 B.n76 71.676
R743 B.n237 B.n77 71.676
R744 B.n241 B.n78 71.676
R745 B.n245 B.n79 71.676
R746 B.n249 B.n80 71.676
R747 B.n253 B.n81 71.676
R748 B.n257 B.n82 71.676
R749 B.n261 B.n83 71.676
R750 B.n265 B.n84 71.676
R751 B.n269 B.n85 71.676
R752 B.n273 B.n86 71.676
R753 B.n277 B.n87 71.676
R754 B.n281 B.n88 71.676
R755 B.n285 B.n89 71.676
R756 B.n675 B.n90 71.676
R757 B.n675 B.n674 71.676
R758 B.n287 B.n89 71.676
R759 B.n284 B.n88 71.676
R760 B.n280 B.n87 71.676
R761 B.n276 B.n86 71.676
R762 B.n272 B.n85 71.676
R763 B.n268 B.n84 71.676
R764 B.n264 B.n83 71.676
R765 B.n260 B.n82 71.676
R766 B.n256 B.n81 71.676
R767 B.n252 B.n80 71.676
R768 B.n248 B.n79 71.676
R769 B.n244 B.n78 71.676
R770 B.n240 B.n77 71.676
R771 B.n236 B.n76 71.676
R772 B.n232 B.n75 71.676
R773 B.n228 B.n74 71.676
R774 B.n224 B.n73 71.676
R775 B.n220 B.n72 71.676
R776 B.n216 B.n71 71.676
R777 B.n212 B.n70 71.676
R778 B.n208 B.n69 71.676
R779 B.n204 B.n68 71.676
R780 B.n200 B.n67 71.676
R781 B.n196 B.n66 71.676
R782 B.n192 B.n65 71.676
R783 B.n188 B.n64 71.676
R784 B.n184 B.n63 71.676
R785 B.n180 B.n62 71.676
R786 B.n176 B.n61 71.676
R787 B.n172 B.n60 71.676
R788 B.n168 B.n59 71.676
R789 B.n164 B.n58 71.676
R790 B.n160 B.n57 71.676
R791 B.n156 B.n56 71.676
R792 B.n152 B.n55 71.676
R793 B.n148 B.n54 71.676
R794 B.n144 B.n53 71.676
R795 B.n140 B.n52 71.676
R796 B.n136 B.n51 71.676
R797 B.n132 B.n50 71.676
R798 B.n128 B.n49 71.676
R799 B.n124 B.n48 71.676
R800 B.n120 B.n47 71.676
R801 B.n116 B.n46 71.676
R802 B.n112 B.n45 71.676
R803 B.n108 B.n44 71.676
R804 B.n104 B.n43 71.676
R805 B.n100 B.n42 71.676
R806 B.n577 B.n576 71.676
R807 B.n571 B.n332 71.676
R808 B.n568 B.n333 71.676
R809 B.n564 B.n334 71.676
R810 B.n560 B.n335 71.676
R811 B.n556 B.n336 71.676
R812 B.n552 B.n337 71.676
R813 B.n548 B.n338 71.676
R814 B.n544 B.n339 71.676
R815 B.n540 B.n340 71.676
R816 B.n536 B.n341 71.676
R817 B.n532 B.n342 71.676
R818 B.n528 B.n343 71.676
R819 B.n524 B.n344 71.676
R820 B.n520 B.n345 71.676
R821 B.n516 B.n346 71.676
R822 B.n512 B.n347 71.676
R823 B.n508 B.n348 71.676
R824 B.n504 B.n349 71.676
R825 B.n500 B.n350 71.676
R826 B.n496 B.n351 71.676
R827 B.n492 B.n352 71.676
R828 B.n487 B.n353 71.676
R829 B.n483 B.n354 71.676
R830 B.n479 B.n355 71.676
R831 B.n475 B.n356 71.676
R832 B.n471 B.n357 71.676
R833 B.n466 B.n358 71.676
R834 B.n462 B.n359 71.676
R835 B.n458 B.n360 71.676
R836 B.n454 B.n361 71.676
R837 B.n450 B.n362 71.676
R838 B.n446 B.n363 71.676
R839 B.n442 B.n364 71.676
R840 B.n438 B.n365 71.676
R841 B.n434 B.n366 71.676
R842 B.n430 B.n367 71.676
R843 B.n426 B.n368 71.676
R844 B.n422 B.n369 71.676
R845 B.n418 B.n370 71.676
R846 B.n414 B.n371 71.676
R847 B.n410 B.n372 71.676
R848 B.n406 B.n373 71.676
R849 B.n402 B.n374 71.676
R850 B.n398 B.n375 71.676
R851 B.n394 B.n376 71.676
R852 B.n390 B.n377 71.676
R853 B.n386 B.n378 71.676
R854 B.n577 B.n380 71.676
R855 B.n569 B.n332 71.676
R856 B.n565 B.n333 71.676
R857 B.n561 B.n334 71.676
R858 B.n557 B.n335 71.676
R859 B.n553 B.n336 71.676
R860 B.n549 B.n337 71.676
R861 B.n545 B.n338 71.676
R862 B.n541 B.n339 71.676
R863 B.n537 B.n340 71.676
R864 B.n533 B.n341 71.676
R865 B.n529 B.n342 71.676
R866 B.n525 B.n343 71.676
R867 B.n521 B.n344 71.676
R868 B.n517 B.n345 71.676
R869 B.n513 B.n346 71.676
R870 B.n509 B.n347 71.676
R871 B.n505 B.n348 71.676
R872 B.n501 B.n349 71.676
R873 B.n497 B.n350 71.676
R874 B.n493 B.n351 71.676
R875 B.n488 B.n352 71.676
R876 B.n484 B.n353 71.676
R877 B.n480 B.n354 71.676
R878 B.n476 B.n355 71.676
R879 B.n472 B.n356 71.676
R880 B.n467 B.n357 71.676
R881 B.n463 B.n358 71.676
R882 B.n459 B.n359 71.676
R883 B.n455 B.n360 71.676
R884 B.n451 B.n361 71.676
R885 B.n447 B.n362 71.676
R886 B.n443 B.n363 71.676
R887 B.n439 B.n364 71.676
R888 B.n435 B.n365 71.676
R889 B.n431 B.n366 71.676
R890 B.n427 B.n367 71.676
R891 B.n423 B.n368 71.676
R892 B.n419 B.n369 71.676
R893 B.n415 B.n370 71.676
R894 B.n411 B.n371 71.676
R895 B.n407 B.n372 71.676
R896 B.n403 B.n373 71.676
R897 B.n399 B.n374 71.676
R898 B.n395 B.n375 71.676
R899 B.n391 B.n376 71.676
R900 B.n387 B.n377 71.676
R901 B.n378 B.n331 71.676
R902 B.n721 B.n720 71.676
R903 B.n721 B.n2 71.676
R904 B.n92 B.t14 68.2522
R905 B.n384 B.t16 68.2522
R906 B.n95 B.t7 68.2354
R907 B.n382 B.t10 68.2354
R908 B.n96 B.n95 59.5399
R909 B.n93 B.n92 59.5399
R910 B.n469 B.n384 59.5399
R911 B.n490 B.n382 59.5399
R912 B.n584 B.n328 41.043
R913 B.n584 B.n324 41.043
R914 B.n590 B.n324 41.043
R915 B.n590 B.n320 41.043
R916 B.n596 B.n320 41.043
R917 B.n602 B.n316 41.043
R918 B.n602 B.n312 41.043
R919 B.n608 B.n312 41.043
R920 B.n608 B.n308 41.043
R921 B.n614 B.n308 41.043
R922 B.n614 B.n304 41.043
R923 B.n620 B.n304 41.043
R924 B.n626 B.n300 41.043
R925 B.n626 B.n296 41.043
R926 B.n633 B.n296 41.043
R927 B.n639 B.n292 41.043
R928 B.n639 B.n4 41.043
R929 B.n719 B.n4 41.043
R930 B.n719 B.n718 41.043
R931 B.n718 B.n717 41.043
R932 B.n717 B.n8 41.043
R933 B.n648 B.n8 41.043
R934 B.n710 B.n709 41.043
R935 B.n709 B.n708 41.043
R936 B.n708 B.n15 41.043
R937 B.n702 B.n701 41.043
R938 B.n701 B.n700 41.043
R939 B.n700 B.n22 41.043
R940 B.n694 B.n22 41.043
R941 B.n694 B.n693 41.043
R942 B.n693 B.n692 41.043
R943 B.n692 B.n29 41.043
R944 B.n686 B.n685 41.043
R945 B.n685 B.n684 41.043
R946 B.n684 B.n36 41.043
R947 B.n678 B.n36 41.043
R948 B.n678 B.n677 41.043
R949 B.n575 B.n326 34.8103
R950 B.n581 B.n580 34.8103
R951 B.n673 B.n672 34.8103
R952 B.n98 B.n38 34.8103
R953 B.t2 B.n300 33.1967
R954 B.t3 B.n15 33.1967
R955 B.n95 B.n94 29.4793
R956 B.n92 B.n91 29.4793
R957 B.n384 B.n383 29.4793
R958 B.n382 B.n381 29.4793
R959 B.n633 B.t0 27.161
R960 B.n710 B.t1 27.161
R961 B.n596 B.t9 21.1253
R962 B.n686 B.t5 21.1253
R963 B.t9 B.n316 19.9182
R964 B.t5 B.n29 19.9182
R965 B B.n722 18.0485
R966 B.t0 B.n292 13.8825
R967 B.n648 B.t1 13.8825
R968 B.n586 B.n326 10.6151
R969 B.n587 B.n586 10.6151
R970 B.n588 B.n587 10.6151
R971 B.n588 B.n318 10.6151
R972 B.n598 B.n318 10.6151
R973 B.n599 B.n598 10.6151
R974 B.n600 B.n599 10.6151
R975 B.n600 B.n310 10.6151
R976 B.n610 B.n310 10.6151
R977 B.n611 B.n610 10.6151
R978 B.n612 B.n611 10.6151
R979 B.n612 B.n302 10.6151
R980 B.n622 B.n302 10.6151
R981 B.n623 B.n622 10.6151
R982 B.n624 B.n623 10.6151
R983 B.n624 B.n294 10.6151
R984 B.n635 B.n294 10.6151
R985 B.n636 B.n635 10.6151
R986 B.n637 B.n636 10.6151
R987 B.n637 B.n0 10.6151
R988 B.n575 B.n574 10.6151
R989 B.n574 B.n573 10.6151
R990 B.n573 B.n572 10.6151
R991 B.n572 B.n570 10.6151
R992 B.n570 B.n567 10.6151
R993 B.n567 B.n566 10.6151
R994 B.n566 B.n563 10.6151
R995 B.n563 B.n562 10.6151
R996 B.n562 B.n559 10.6151
R997 B.n559 B.n558 10.6151
R998 B.n558 B.n555 10.6151
R999 B.n555 B.n554 10.6151
R1000 B.n554 B.n551 10.6151
R1001 B.n551 B.n550 10.6151
R1002 B.n550 B.n547 10.6151
R1003 B.n547 B.n546 10.6151
R1004 B.n546 B.n543 10.6151
R1005 B.n543 B.n542 10.6151
R1006 B.n542 B.n539 10.6151
R1007 B.n539 B.n538 10.6151
R1008 B.n538 B.n535 10.6151
R1009 B.n535 B.n534 10.6151
R1010 B.n534 B.n531 10.6151
R1011 B.n531 B.n530 10.6151
R1012 B.n530 B.n527 10.6151
R1013 B.n527 B.n526 10.6151
R1014 B.n526 B.n523 10.6151
R1015 B.n523 B.n522 10.6151
R1016 B.n522 B.n519 10.6151
R1017 B.n519 B.n518 10.6151
R1018 B.n518 B.n515 10.6151
R1019 B.n515 B.n514 10.6151
R1020 B.n514 B.n511 10.6151
R1021 B.n511 B.n510 10.6151
R1022 B.n510 B.n507 10.6151
R1023 B.n507 B.n506 10.6151
R1024 B.n506 B.n503 10.6151
R1025 B.n503 B.n502 10.6151
R1026 B.n502 B.n499 10.6151
R1027 B.n499 B.n498 10.6151
R1028 B.n498 B.n495 10.6151
R1029 B.n495 B.n494 10.6151
R1030 B.n494 B.n491 10.6151
R1031 B.n489 B.n486 10.6151
R1032 B.n486 B.n485 10.6151
R1033 B.n485 B.n482 10.6151
R1034 B.n482 B.n481 10.6151
R1035 B.n481 B.n478 10.6151
R1036 B.n478 B.n477 10.6151
R1037 B.n477 B.n474 10.6151
R1038 B.n474 B.n473 10.6151
R1039 B.n473 B.n470 10.6151
R1040 B.n468 B.n465 10.6151
R1041 B.n465 B.n464 10.6151
R1042 B.n464 B.n461 10.6151
R1043 B.n461 B.n460 10.6151
R1044 B.n460 B.n457 10.6151
R1045 B.n457 B.n456 10.6151
R1046 B.n456 B.n453 10.6151
R1047 B.n453 B.n452 10.6151
R1048 B.n452 B.n449 10.6151
R1049 B.n449 B.n448 10.6151
R1050 B.n448 B.n445 10.6151
R1051 B.n445 B.n444 10.6151
R1052 B.n444 B.n441 10.6151
R1053 B.n441 B.n440 10.6151
R1054 B.n440 B.n437 10.6151
R1055 B.n437 B.n436 10.6151
R1056 B.n436 B.n433 10.6151
R1057 B.n433 B.n432 10.6151
R1058 B.n432 B.n429 10.6151
R1059 B.n429 B.n428 10.6151
R1060 B.n428 B.n425 10.6151
R1061 B.n425 B.n424 10.6151
R1062 B.n424 B.n421 10.6151
R1063 B.n421 B.n420 10.6151
R1064 B.n420 B.n417 10.6151
R1065 B.n417 B.n416 10.6151
R1066 B.n416 B.n413 10.6151
R1067 B.n413 B.n412 10.6151
R1068 B.n412 B.n409 10.6151
R1069 B.n409 B.n408 10.6151
R1070 B.n408 B.n405 10.6151
R1071 B.n405 B.n404 10.6151
R1072 B.n404 B.n401 10.6151
R1073 B.n401 B.n400 10.6151
R1074 B.n400 B.n397 10.6151
R1075 B.n397 B.n396 10.6151
R1076 B.n396 B.n393 10.6151
R1077 B.n393 B.n392 10.6151
R1078 B.n392 B.n389 10.6151
R1079 B.n389 B.n388 10.6151
R1080 B.n388 B.n385 10.6151
R1081 B.n385 B.n330 10.6151
R1082 B.n580 B.n330 10.6151
R1083 B.n582 B.n581 10.6151
R1084 B.n582 B.n322 10.6151
R1085 B.n592 B.n322 10.6151
R1086 B.n593 B.n592 10.6151
R1087 B.n594 B.n593 10.6151
R1088 B.n594 B.n314 10.6151
R1089 B.n604 B.n314 10.6151
R1090 B.n605 B.n604 10.6151
R1091 B.n606 B.n605 10.6151
R1092 B.n606 B.n306 10.6151
R1093 B.n616 B.n306 10.6151
R1094 B.n617 B.n616 10.6151
R1095 B.n618 B.n617 10.6151
R1096 B.n618 B.n298 10.6151
R1097 B.n628 B.n298 10.6151
R1098 B.n629 B.n628 10.6151
R1099 B.n631 B.n629 10.6151
R1100 B.n631 B.n630 10.6151
R1101 B.n630 B.n290 10.6151
R1102 B.n642 B.n290 10.6151
R1103 B.n643 B.n642 10.6151
R1104 B.n644 B.n643 10.6151
R1105 B.n645 B.n644 10.6151
R1106 B.n646 B.n645 10.6151
R1107 B.n650 B.n646 10.6151
R1108 B.n651 B.n650 10.6151
R1109 B.n652 B.n651 10.6151
R1110 B.n653 B.n652 10.6151
R1111 B.n655 B.n653 10.6151
R1112 B.n656 B.n655 10.6151
R1113 B.n657 B.n656 10.6151
R1114 B.n658 B.n657 10.6151
R1115 B.n660 B.n658 10.6151
R1116 B.n661 B.n660 10.6151
R1117 B.n662 B.n661 10.6151
R1118 B.n663 B.n662 10.6151
R1119 B.n665 B.n663 10.6151
R1120 B.n666 B.n665 10.6151
R1121 B.n667 B.n666 10.6151
R1122 B.n668 B.n667 10.6151
R1123 B.n670 B.n668 10.6151
R1124 B.n671 B.n670 10.6151
R1125 B.n672 B.n671 10.6151
R1126 B.n714 B.n1 10.6151
R1127 B.n714 B.n713 10.6151
R1128 B.n713 B.n712 10.6151
R1129 B.n712 B.n10 10.6151
R1130 B.n706 B.n10 10.6151
R1131 B.n706 B.n705 10.6151
R1132 B.n705 B.n704 10.6151
R1133 B.n704 B.n17 10.6151
R1134 B.n698 B.n17 10.6151
R1135 B.n698 B.n697 10.6151
R1136 B.n697 B.n696 10.6151
R1137 B.n696 B.n24 10.6151
R1138 B.n690 B.n24 10.6151
R1139 B.n690 B.n689 10.6151
R1140 B.n689 B.n688 10.6151
R1141 B.n688 B.n31 10.6151
R1142 B.n682 B.n31 10.6151
R1143 B.n682 B.n681 10.6151
R1144 B.n681 B.n680 10.6151
R1145 B.n680 B.n38 10.6151
R1146 B.n99 B.n98 10.6151
R1147 B.n102 B.n99 10.6151
R1148 B.n103 B.n102 10.6151
R1149 B.n106 B.n103 10.6151
R1150 B.n107 B.n106 10.6151
R1151 B.n110 B.n107 10.6151
R1152 B.n111 B.n110 10.6151
R1153 B.n114 B.n111 10.6151
R1154 B.n115 B.n114 10.6151
R1155 B.n118 B.n115 10.6151
R1156 B.n119 B.n118 10.6151
R1157 B.n122 B.n119 10.6151
R1158 B.n123 B.n122 10.6151
R1159 B.n126 B.n123 10.6151
R1160 B.n127 B.n126 10.6151
R1161 B.n130 B.n127 10.6151
R1162 B.n131 B.n130 10.6151
R1163 B.n134 B.n131 10.6151
R1164 B.n135 B.n134 10.6151
R1165 B.n138 B.n135 10.6151
R1166 B.n139 B.n138 10.6151
R1167 B.n142 B.n139 10.6151
R1168 B.n143 B.n142 10.6151
R1169 B.n146 B.n143 10.6151
R1170 B.n147 B.n146 10.6151
R1171 B.n150 B.n147 10.6151
R1172 B.n151 B.n150 10.6151
R1173 B.n154 B.n151 10.6151
R1174 B.n155 B.n154 10.6151
R1175 B.n158 B.n155 10.6151
R1176 B.n159 B.n158 10.6151
R1177 B.n162 B.n159 10.6151
R1178 B.n163 B.n162 10.6151
R1179 B.n166 B.n163 10.6151
R1180 B.n167 B.n166 10.6151
R1181 B.n170 B.n167 10.6151
R1182 B.n171 B.n170 10.6151
R1183 B.n174 B.n171 10.6151
R1184 B.n175 B.n174 10.6151
R1185 B.n178 B.n175 10.6151
R1186 B.n179 B.n178 10.6151
R1187 B.n182 B.n179 10.6151
R1188 B.n183 B.n182 10.6151
R1189 B.n187 B.n186 10.6151
R1190 B.n190 B.n187 10.6151
R1191 B.n191 B.n190 10.6151
R1192 B.n194 B.n191 10.6151
R1193 B.n195 B.n194 10.6151
R1194 B.n198 B.n195 10.6151
R1195 B.n199 B.n198 10.6151
R1196 B.n202 B.n199 10.6151
R1197 B.n203 B.n202 10.6151
R1198 B.n207 B.n206 10.6151
R1199 B.n210 B.n207 10.6151
R1200 B.n211 B.n210 10.6151
R1201 B.n214 B.n211 10.6151
R1202 B.n215 B.n214 10.6151
R1203 B.n218 B.n215 10.6151
R1204 B.n219 B.n218 10.6151
R1205 B.n222 B.n219 10.6151
R1206 B.n223 B.n222 10.6151
R1207 B.n226 B.n223 10.6151
R1208 B.n227 B.n226 10.6151
R1209 B.n230 B.n227 10.6151
R1210 B.n231 B.n230 10.6151
R1211 B.n234 B.n231 10.6151
R1212 B.n235 B.n234 10.6151
R1213 B.n238 B.n235 10.6151
R1214 B.n239 B.n238 10.6151
R1215 B.n242 B.n239 10.6151
R1216 B.n243 B.n242 10.6151
R1217 B.n246 B.n243 10.6151
R1218 B.n247 B.n246 10.6151
R1219 B.n250 B.n247 10.6151
R1220 B.n251 B.n250 10.6151
R1221 B.n254 B.n251 10.6151
R1222 B.n255 B.n254 10.6151
R1223 B.n258 B.n255 10.6151
R1224 B.n259 B.n258 10.6151
R1225 B.n262 B.n259 10.6151
R1226 B.n263 B.n262 10.6151
R1227 B.n266 B.n263 10.6151
R1228 B.n267 B.n266 10.6151
R1229 B.n270 B.n267 10.6151
R1230 B.n271 B.n270 10.6151
R1231 B.n274 B.n271 10.6151
R1232 B.n275 B.n274 10.6151
R1233 B.n278 B.n275 10.6151
R1234 B.n279 B.n278 10.6151
R1235 B.n282 B.n279 10.6151
R1236 B.n283 B.n282 10.6151
R1237 B.n286 B.n283 10.6151
R1238 B.n288 B.n286 10.6151
R1239 B.n289 B.n288 10.6151
R1240 B.n673 B.n289 10.6151
R1241 B.n491 B.n490 9.36635
R1242 B.n469 B.n468 9.36635
R1243 B.n183 B.n96 9.36635
R1244 B.n206 B.n93 9.36635
R1245 B.n722 B.n0 8.11757
R1246 B.n722 B.n1 8.11757
R1247 B.n620 B.t2 7.84686
R1248 B.n702 B.t3 7.84686
R1249 B.n490 B.n489 1.24928
R1250 B.n470 B.n469 1.24928
R1251 B.n186 B.n96 1.24928
R1252 B.n203 B.n93 1.24928
R1253 VN.n0 VN.t1 298.18
R1254 VN.n1 VN.t2 298.18
R1255 VN.n0 VN.t3 297.961
R1256 VN.n1 VN.t0 297.961
R1257 VN VN.n1 61.4982
R1258 VN VN.n0 18.5626
R1259 VDD2.n2 VDD2.n0 102.118
R1260 VDD2.n2 VDD2.n1 63.3091
R1261 VDD2.n1 VDD2.t3 1.52946
R1262 VDD2.n1 VDD2.t1 1.52946
R1263 VDD2.n0 VDD2.t2 1.52946
R1264 VDD2.n0 VDD2.t0 1.52946
R1265 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.147538f
C1 VN VTAIL 3.83426f
C2 VDD1 VP 4.34042f
C3 VN VDD2 4.18395f
C4 VTAIL VP 3.84837f
C5 VDD1 VTAIL 6.10601f
C6 VP VDD2 0.304397f
C7 VN VP 5.35361f
C8 VDD1 VDD2 0.681986f
C9 VTAIL VDD2 6.15077f
C10 VDD2 B 3.048965f
C11 VDD1 B 6.84165f
C12 VTAIL B 9.718522f
C13 VN B 8.56203f
C14 VP B 6.000906f
C15 VDD2.t2 B 0.277531f
C16 VDD2.t0 B 0.277531f
C17 VDD2.n0 B 3.12157f
C18 VDD2.t3 B 0.277531f
C19 VDD2.t1 B 0.277531f
C20 VDD2.n1 B 2.49296f
C21 VDD2.n2 B 3.555f
C22 VN.t1 B 1.74842f
C23 VN.t3 B 1.74786f
C24 VN.n0 B 1.32098f
C25 VN.t2 B 1.74842f
C26 VN.t0 B 1.74786f
C27 VN.n1 B 2.62391f
C28 VTAIL.t1 B 1.78548f
C29 VTAIL.n0 B 0.261257f
C30 VTAIL.t4 B 1.78548f
C31 VTAIL.n1 B 0.291477f
C32 VTAIL.t6 B 1.78548f
C33 VTAIL.n2 B 1.11256f
C34 VTAIL.t2 B 1.78549f
C35 VTAIL.n3 B 1.11255f
C36 VTAIL.t0 B 1.78549f
C37 VTAIL.n4 B 0.291467f
C38 VTAIL.t3 B 1.78549f
C39 VTAIL.n5 B 0.291467f
C40 VTAIL.t5 B 1.78548f
C41 VTAIL.n6 B 1.11256f
C42 VTAIL.t7 B 1.78548f
C43 VTAIL.n7 B 1.07645f
C44 VDD1.t3 B 0.274884f
C45 VDD1.t0 B 0.274884f
C46 VDD1.n0 B 2.46949f
C47 VDD1.t2 B 0.274884f
C48 VDD1.t1 B 0.274884f
C49 VDD1.n1 B 3.11771f
C50 VP.n0 B 0.039929f
C51 VP.t2 B 1.68006f
C52 VP.n1 B 0.061724f
C53 VP.t3 B 1.76879f
C54 VP.t1 B 1.76823f
C55 VP.n2 B 2.63269f
C56 VP.t0 B 1.68006f
C57 VP.n3 B 0.677499f
C58 VP.n4 B 2.28976f
C59 VP.n5 B 0.039929f
C60 VP.n6 B 0.039929f
C61 VP.n7 B 0.032279f
C62 VP.n8 B 0.061724f
C63 VP.n9 B 0.677499f
C64 VP.n10 B 0.035745f
.ends

