* NGSPICE file created from diff_pair_sample_1117.ext - technology: sky130A

.subckt diff_pair_sample_1117 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0.78705 ps=5.1 w=4.77 l=0.85
X1 VTAIL.t6 VN.t1 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0.78705 ps=5.1 w=4.77 l=0.85
X2 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.78705 pd=5.1 as=1.8603 ps=10.32 w=4.77 l=0.85
X3 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.78705 pd=5.1 as=1.8603 ps=10.32 w=4.77 l=0.85
X4 VDD2.t2 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.78705 pd=5.1 as=1.8603 ps=10.32 w=4.77 l=0.85
X5 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0.78705 ps=5.1 w=4.77 l=0.85
X6 VDD2.t1 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.78705 pd=5.1 as=1.8603 ps=10.32 w=4.77 l=0.85
X7 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0.78705 ps=5.1 w=4.77 l=0.85
X8 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0 ps=0 w=4.77 l=0.85
X9 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0 ps=0 w=4.77 l=0.85
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0 ps=0 w=4.77 l=0.85
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8603 pd=10.32 as=0 ps=0 w=4.77 l=0.85
R0 VN.n0 VN.t0 202.739
R1 VN.n1 VN.t3 202.739
R2 VN.n0 VN.t2 202.69
R3 VN.n1 VN.t1 202.69
R4 VN VN.n1 80.5428
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 103.409
R7 VDD2.n2 VDD2.n1 72.5315
R8 VDD2.n1 VDD2.t0 4.15144
R9 VDD2.n1 VDD2.t1 4.15144
R10 VDD2.n0 VDD2.t3 4.15144
R11 VDD2.n0 VDD2.t2 4.15144
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 60.0045
R14 VTAIL.n4 VTAIL.t4 60.0045
R15 VTAIL.n3 VTAIL.t6 60.0045
R16 VTAIL.n6 VTAIL.t3 60.0036
R17 VTAIL.n7 VTAIL.t5 60.0035
R18 VTAIL.n0 VTAIL.t7 60.0035
R19 VTAIL.n1 VTAIL.t2 60.0035
R20 VTAIL.n2 VTAIL.t0 60.0035
R21 VTAIL.n7 VTAIL.n6 17.4962
R22 VTAIL.n3 VTAIL.n2 17.4962
R23 VTAIL.n4 VTAIL.n3 1.01774
R24 VTAIL.n6 VTAIL.n5 1.01774
R25 VTAIL.n2 VTAIL.n1 1.01774
R26 VTAIL VTAIL.n0 0.56731
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.450931
R30 B.n312 B.n311 585
R31 B.n314 B.n67 585
R32 B.n317 B.n316 585
R33 B.n318 B.n66 585
R34 B.n320 B.n319 585
R35 B.n322 B.n65 585
R36 B.n325 B.n324 585
R37 B.n326 B.n64 585
R38 B.n328 B.n327 585
R39 B.n330 B.n63 585
R40 B.n333 B.n332 585
R41 B.n334 B.n62 585
R42 B.n336 B.n335 585
R43 B.n338 B.n61 585
R44 B.n341 B.n340 585
R45 B.n342 B.n60 585
R46 B.n344 B.n343 585
R47 B.n346 B.n59 585
R48 B.n348 B.n347 585
R49 B.n350 B.n349 585
R50 B.n353 B.n352 585
R51 B.n354 B.n54 585
R52 B.n356 B.n355 585
R53 B.n358 B.n53 585
R54 B.n361 B.n360 585
R55 B.n362 B.n52 585
R56 B.n364 B.n363 585
R57 B.n366 B.n51 585
R58 B.n369 B.n368 585
R59 B.n370 B.n48 585
R60 B.n373 B.n372 585
R61 B.n375 B.n47 585
R62 B.n378 B.n377 585
R63 B.n379 B.n46 585
R64 B.n381 B.n380 585
R65 B.n383 B.n45 585
R66 B.n386 B.n385 585
R67 B.n387 B.n44 585
R68 B.n389 B.n388 585
R69 B.n391 B.n43 585
R70 B.n394 B.n393 585
R71 B.n395 B.n42 585
R72 B.n397 B.n396 585
R73 B.n399 B.n41 585
R74 B.n402 B.n401 585
R75 B.n403 B.n40 585
R76 B.n405 B.n404 585
R77 B.n407 B.n39 585
R78 B.n410 B.n409 585
R79 B.n411 B.n38 585
R80 B.n310 B.n36 585
R81 B.n414 B.n36 585
R82 B.n309 B.n35 585
R83 B.n415 B.n35 585
R84 B.n308 B.n34 585
R85 B.n416 B.n34 585
R86 B.n307 B.n306 585
R87 B.n306 B.n30 585
R88 B.n305 B.n29 585
R89 B.n422 B.n29 585
R90 B.n304 B.n28 585
R91 B.n423 B.n28 585
R92 B.n303 B.n27 585
R93 B.n424 B.n27 585
R94 B.n302 B.n301 585
R95 B.n301 B.n23 585
R96 B.n300 B.n22 585
R97 B.n430 B.n22 585
R98 B.n299 B.n21 585
R99 B.n431 B.n21 585
R100 B.n298 B.n20 585
R101 B.n432 B.n20 585
R102 B.n297 B.n296 585
R103 B.n296 B.n19 585
R104 B.n295 B.n15 585
R105 B.n438 B.n15 585
R106 B.n294 B.n14 585
R107 B.n439 B.n14 585
R108 B.n293 B.n13 585
R109 B.n440 B.n13 585
R110 B.n292 B.n291 585
R111 B.n291 B.n12 585
R112 B.n290 B.n289 585
R113 B.n290 B.n8 585
R114 B.n288 B.n7 585
R115 B.n447 B.n7 585
R116 B.n287 B.n6 585
R117 B.n448 B.n6 585
R118 B.n286 B.n5 585
R119 B.n449 B.n5 585
R120 B.n285 B.n284 585
R121 B.n284 B.n4 585
R122 B.n283 B.n68 585
R123 B.n283 B.n282 585
R124 B.n272 B.n69 585
R125 B.n275 B.n69 585
R126 B.n274 B.n273 585
R127 B.n276 B.n274 585
R128 B.n271 B.n74 585
R129 B.n74 B.n73 585
R130 B.n270 B.n269 585
R131 B.n269 B.n268 585
R132 B.n76 B.n75 585
R133 B.n261 B.n76 585
R134 B.n260 B.n259 585
R135 B.n262 B.n260 585
R136 B.n258 B.n81 585
R137 B.n81 B.n80 585
R138 B.n257 B.n256 585
R139 B.n256 B.n255 585
R140 B.n83 B.n82 585
R141 B.n84 B.n83 585
R142 B.n248 B.n247 585
R143 B.n249 B.n248 585
R144 B.n246 B.n88 585
R145 B.n92 B.n88 585
R146 B.n245 B.n244 585
R147 B.n244 B.n243 585
R148 B.n90 B.n89 585
R149 B.n91 B.n90 585
R150 B.n236 B.n235 585
R151 B.n237 B.n236 585
R152 B.n234 B.n97 585
R153 B.n97 B.n96 585
R154 B.n233 B.n232 585
R155 B.n232 B.n231 585
R156 B.n228 B.n101 585
R157 B.n227 B.n226 585
R158 B.n224 B.n102 585
R159 B.n224 B.n100 585
R160 B.n223 B.n222 585
R161 B.n221 B.n220 585
R162 B.n219 B.n104 585
R163 B.n217 B.n216 585
R164 B.n215 B.n105 585
R165 B.n214 B.n213 585
R166 B.n211 B.n106 585
R167 B.n209 B.n208 585
R168 B.n207 B.n107 585
R169 B.n206 B.n205 585
R170 B.n203 B.n108 585
R171 B.n201 B.n200 585
R172 B.n199 B.n109 585
R173 B.n198 B.n197 585
R174 B.n195 B.n110 585
R175 B.n193 B.n192 585
R176 B.n191 B.n111 585
R177 B.n189 B.n188 585
R178 B.n186 B.n114 585
R179 B.n184 B.n183 585
R180 B.n182 B.n115 585
R181 B.n181 B.n180 585
R182 B.n178 B.n116 585
R183 B.n176 B.n175 585
R184 B.n174 B.n117 585
R185 B.n173 B.n172 585
R186 B.n170 B.n118 585
R187 B.n168 B.n167 585
R188 B.n166 B.n119 585
R189 B.n165 B.n164 585
R190 B.n162 B.n123 585
R191 B.n160 B.n159 585
R192 B.n158 B.n124 585
R193 B.n157 B.n156 585
R194 B.n154 B.n125 585
R195 B.n152 B.n151 585
R196 B.n150 B.n126 585
R197 B.n149 B.n148 585
R198 B.n146 B.n127 585
R199 B.n144 B.n143 585
R200 B.n142 B.n128 585
R201 B.n141 B.n140 585
R202 B.n138 B.n129 585
R203 B.n136 B.n135 585
R204 B.n134 B.n130 585
R205 B.n133 B.n132 585
R206 B.n99 B.n98 585
R207 B.n100 B.n99 585
R208 B.n230 B.n229 585
R209 B.n231 B.n230 585
R210 B.n95 B.n94 585
R211 B.n96 B.n95 585
R212 B.n239 B.n238 585
R213 B.n238 B.n237 585
R214 B.n240 B.n93 585
R215 B.n93 B.n91 585
R216 B.n242 B.n241 585
R217 B.n243 B.n242 585
R218 B.n87 B.n86 585
R219 B.n92 B.n87 585
R220 B.n251 B.n250 585
R221 B.n250 B.n249 585
R222 B.n252 B.n85 585
R223 B.n85 B.n84 585
R224 B.n254 B.n253 585
R225 B.n255 B.n254 585
R226 B.n79 B.n78 585
R227 B.n80 B.n79 585
R228 B.n264 B.n263 585
R229 B.n263 B.n262 585
R230 B.n265 B.n77 585
R231 B.n261 B.n77 585
R232 B.n267 B.n266 585
R233 B.n268 B.n267 585
R234 B.n72 B.n71 585
R235 B.n73 B.n72 585
R236 B.n278 B.n277 585
R237 B.n277 B.n276 585
R238 B.n279 B.n70 585
R239 B.n275 B.n70 585
R240 B.n281 B.n280 585
R241 B.n282 B.n281 585
R242 B.n3 B.n0 585
R243 B.n4 B.n3 585
R244 B.n446 B.n1 585
R245 B.n447 B.n446 585
R246 B.n445 B.n444 585
R247 B.n445 B.n8 585
R248 B.n443 B.n9 585
R249 B.n12 B.n9 585
R250 B.n442 B.n441 585
R251 B.n441 B.n440 585
R252 B.n11 B.n10 585
R253 B.n439 B.n11 585
R254 B.n437 B.n436 585
R255 B.n438 B.n437 585
R256 B.n435 B.n16 585
R257 B.n19 B.n16 585
R258 B.n434 B.n433 585
R259 B.n433 B.n432 585
R260 B.n18 B.n17 585
R261 B.n431 B.n18 585
R262 B.n429 B.n428 585
R263 B.n430 B.n429 585
R264 B.n427 B.n24 585
R265 B.n24 B.n23 585
R266 B.n426 B.n425 585
R267 B.n425 B.n424 585
R268 B.n26 B.n25 585
R269 B.n423 B.n26 585
R270 B.n421 B.n420 585
R271 B.n422 B.n421 585
R272 B.n419 B.n31 585
R273 B.n31 B.n30 585
R274 B.n418 B.n417 585
R275 B.n417 B.n416 585
R276 B.n33 B.n32 585
R277 B.n415 B.n33 585
R278 B.n413 B.n412 585
R279 B.n414 B.n413 585
R280 B.n450 B.n449 585
R281 B.n448 B.n2 585
R282 B.n413 B.n38 526.135
R283 B.n312 B.n36 526.135
R284 B.n232 B.n99 526.135
R285 B.n230 B.n101 526.135
R286 B.n49 B.t11 337.033
R287 B.n55 B.t15 337.033
R288 B.n120 B.t4 337.033
R289 B.n112 B.t8 337.033
R290 B.n313 B.n37 256.663
R291 B.n315 B.n37 256.663
R292 B.n321 B.n37 256.663
R293 B.n323 B.n37 256.663
R294 B.n329 B.n37 256.663
R295 B.n331 B.n37 256.663
R296 B.n337 B.n37 256.663
R297 B.n339 B.n37 256.663
R298 B.n345 B.n37 256.663
R299 B.n58 B.n37 256.663
R300 B.n351 B.n37 256.663
R301 B.n357 B.n37 256.663
R302 B.n359 B.n37 256.663
R303 B.n365 B.n37 256.663
R304 B.n367 B.n37 256.663
R305 B.n374 B.n37 256.663
R306 B.n376 B.n37 256.663
R307 B.n382 B.n37 256.663
R308 B.n384 B.n37 256.663
R309 B.n390 B.n37 256.663
R310 B.n392 B.n37 256.663
R311 B.n398 B.n37 256.663
R312 B.n400 B.n37 256.663
R313 B.n406 B.n37 256.663
R314 B.n408 B.n37 256.663
R315 B.n225 B.n100 256.663
R316 B.n103 B.n100 256.663
R317 B.n218 B.n100 256.663
R318 B.n212 B.n100 256.663
R319 B.n210 B.n100 256.663
R320 B.n204 B.n100 256.663
R321 B.n202 B.n100 256.663
R322 B.n196 B.n100 256.663
R323 B.n194 B.n100 256.663
R324 B.n187 B.n100 256.663
R325 B.n185 B.n100 256.663
R326 B.n179 B.n100 256.663
R327 B.n177 B.n100 256.663
R328 B.n171 B.n100 256.663
R329 B.n169 B.n100 256.663
R330 B.n163 B.n100 256.663
R331 B.n161 B.n100 256.663
R332 B.n155 B.n100 256.663
R333 B.n153 B.n100 256.663
R334 B.n147 B.n100 256.663
R335 B.n145 B.n100 256.663
R336 B.n139 B.n100 256.663
R337 B.n137 B.n100 256.663
R338 B.n131 B.n100 256.663
R339 B.n452 B.n451 256.663
R340 B.n409 B.n407 163.367
R341 B.n405 B.n40 163.367
R342 B.n401 B.n399 163.367
R343 B.n397 B.n42 163.367
R344 B.n393 B.n391 163.367
R345 B.n389 B.n44 163.367
R346 B.n385 B.n383 163.367
R347 B.n381 B.n46 163.367
R348 B.n377 B.n375 163.367
R349 B.n373 B.n48 163.367
R350 B.n368 B.n366 163.367
R351 B.n364 B.n52 163.367
R352 B.n360 B.n358 163.367
R353 B.n356 B.n54 163.367
R354 B.n352 B.n350 163.367
R355 B.n347 B.n346 163.367
R356 B.n344 B.n60 163.367
R357 B.n340 B.n338 163.367
R358 B.n336 B.n62 163.367
R359 B.n332 B.n330 163.367
R360 B.n328 B.n64 163.367
R361 B.n324 B.n322 163.367
R362 B.n320 B.n66 163.367
R363 B.n316 B.n314 163.367
R364 B.n232 B.n97 163.367
R365 B.n236 B.n97 163.367
R366 B.n236 B.n90 163.367
R367 B.n244 B.n90 163.367
R368 B.n244 B.n88 163.367
R369 B.n248 B.n88 163.367
R370 B.n248 B.n83 163.367
R371 B.n256 B.n83 163.367
R372 B.n256 B.n81 163.367
R373 B.n260 B.n81 163.367
R374 B.n260 B.n76 163.367
R375 B.n269 B.n76 163.367
R376 B.n269 B.n74 163.367
R377 B.n274 B.n74 163.367
R378 B.n274 B.n69 163.367
R379 B.n283 B.n69 163.367
R380 B.n284 B.n283 163.367
R381 B.n284 B.n5 163.367
R382 B.n6 B.n5 163.367
R383 B.n7 B.n6 163.367
R384 B.n290 B.n7 163.367
R385 B.n291 B.n290 163.367
R386 B.n291 B.n13 163.367
R387 B.n14 B.n13 163.367
R388 B.n15 B.n14 163.367
R389 B.n296 B.n15 163.367
R390 B.n296 B.n20 163.367
R391 B.n21 B.n20 163.367
R392 B.n22 B.n21 163.367
R393 B.n301 B.n22 163.367
R394 B.n301 B.n27 163.367
R395 B.n28 B.n27 163.367
R396 B.n29 B.n28 163.367
R397 B.n306 B.n29 163.367
R398 B.n306 B.n34 163.367
R399 B.n35 B.n34 163.367
R400 B.n36 B.n35 163.367
R401 B.n226 B.n224 163.367
R402 B.n224 B.n223 163.367
R403 B.n220 B.n219 163.367
R404 B.n217 B.n105 163.367
R405 B.n213 B.n211 163.367
R406 B.n209 B.n107 163.367
R407 B.n205 B.n203 163.367
R408 B.n201 B.n109 163.367
R409 B.n197 B.n195 163.367
R410 B.n193 B.n111 163.367
R411 B.n188 B.n186 163.367
R412 B.n184 B.n115 163.367
R413 B.n180 B.n178 163.367
R414 B.n176 B.n117 163.367
R415 B.n172 B.n170 163.367
R416 B.n168 B.n119 163.367
R417 B.n164 B.n162 163.367
R418 B.n160 B.n124 163.367
R419 B.n156 B.n154 163.367
R420 B.n152 B.n126 163.367
R421 B.n148 B.n146 163.367
R422 B.n144 B.n128 163.367
R423 B.n140 B.n138 163.367
R424 B.n136 B.n130 163.367
R425 B.n132 B.n99 163.367
R426 B.n230 B.n95 163.367
R427 B.n238 B.n95 163.367
R428 B.n238 B.n93 163.367
R429 B.n242 B.n93 163.367
R430 B.n242 B.n87 163.367
R431 B.n250 B.n87 163.367
R432 B.n250 B.n85 163.367
R433 B.n254 B.n85 163.367
R434 B.n254 B.n79 163.367
R435 B.n263 B.n79 163.367
R436 B.n263 B.n77 163.367
R437 B.n267 B.n77 163.367
R438 B.n267 B.n72 163.367
R439 B.n277 B.n72 163.367
R440 B.n277 B.n70 163.367
R441 B.n281 B.n70 163.367
R442 B.n281 B.n3 163.367
R443 B.n450 B.n3 163.367
R444 B.n446 B.n2 163.367
R445 B.n446 B.n445 163.367
R446 B.n445 B.n9 163.367
R447 B.n441 B.n9 163.367
R448 B.n441 B.n11 163.367
R449 B.n437 B.n11 163.367
R450 B.n437 B.n16 163.367
R451 B.n433 B.n16 163.367
R452 B.n433 B.n18 163.367
R453 B.n429 B.n18 163.367
R454 B.n429 B.n24 163.367
R455 B.n425 B.n24 163.367
R456 B.n425 B.n26 163.367
R457 B.n421 B.n26 163.367
R458 B.n421 B.n31 163.367
R459 B.n417 B.n31 163.367
R460 B.n417 B.n33 163.367
R461 B.n413 B.n33 163.367
R462 B.n231 B.n100 136.885
R463 B.n414 B.n37 136.885
R464 B.n55 B.t16 93.4576
R465 B.n120 B.t7 93.4576
R466 B.n49 B.t13 93.4528
R467 B.n112 B.t10 93.4528
R468 B.n231 B.n96 74.4654
R469 B.n237 B.n96 74.4654
R470 B.n237 B.n91 74.4654
R471 B.n243 B.n91 74.4654
R472 B.n243 B.n92 74.4654
R473 B.n249 B.n84 74.4654
R474 B.n255 B.n84 74.4654
R475 B.n255 B.n80 74.4654
R476 B.n262 B.n80 74.4654
R477 B.n262 B.n261 74.4654
R478 B.n268 B.n73 74.4654
R479 B.n276 B.n73 74.4654
R480 B.n276 B.n275 74.4654
R481 B.n282 B.n4 74.4654
R482 B.n449 B.n4 74.4654
R483 B.n449 B.n448 74.4654
R484 B.n448 B.n447 74.4654
R485 B.n447 B.n8 74.4654
R486 B.n440 B.n12 74.4654
R487 B.n440 B.n439 74.4654
R488 B.n439 B.n438 74.4654
R489 B.n432 B.n19 74.4654
R490 B.n432 B.n431 74.4654
R491 B.n431 B.n430 74.4654
R492 B.n430 B.n23 74.4654
R493 B.n424 B.n23 74.4654
R494 B.n423 B.n422 74.4654
R495 B.n422 B.n30 74.4654
R496 B.n416 B.n30 74.4654
R497 B.n416 B.n415 74.4654
R498 B.n415 B.n414 74.4654
R499 B.n249 B.t5 73.3703
R500 B.n424 B.t12 73.3703
R501 B.n408 B.n38 71.676
R502 B.n407 B.n406 71.676
R503 B.n400 B.n40 71.676
R504 B.n399 B.n398 71.676
R505 B.n392 B.n42 71.676
R506 B.n391 B.n390 71.676
R507 B.n384 B.n44 71.676
R508 B.n383 B.n382 71.676
R509 B.n376 B.n46 71.676
R510 B.n375 B.n374 71.676
R511 B.n367 B.n48 71.676
R512 B.n366 B.n365 71.676
R513 B.n359 B.n52 71.676
R514 B.n358 B.n357 71.676
R515 B.n351 B.n54 71.676
R516 B.n350 B.n58 71.676
R517 B.n346 B.n345 71.676
R518 B.n339 B.n60 71.676
R519 B.n338 B.n337 71.676
R520 B.n331 B.n62 71.676
R521 B.n330 B.n329 71.676
R522 B.n323 B.n64 71.676
R523 B.n322 B.n321 71.676
R524 B.n315 B.n66 71.676
R525 B.n314 B.n313 71.676
R526 B.n313 B.n312 71.676
R527 B.n316 B.n315 71.676
R528 B.n321 B.n320 71.676
R529 B.n324 B.n323 71.676
R530 B.n329 B.n328 71.676
R531 B.n332 B.n331 71.676
R532 B.n337 B.n336 71.676
R533 B.n340 B.n339 71.676
R534 B.n345 B.n344 71.676
R535 B.n347 B.n58 71.676
R536 B.n352 B.n351 71.676
R537 B.n357 B.n356 71.676
R538 B.n360 B.n359 71.676
R539 B.n365 B.n364 71.676
R540 B.n368 B.n367 71.676
R541 B.n374 B.n373 71.676
R542 B.n377 B.n376 71.676
R543 B.n382 B.n381 71.676
R544 B.n385 B.n384 71.676
R545 B.n390 B.n389 71.676
R546 B.n393 B.n392 71.676
R547 B.n398 B.n397 71.676
R548 B.n401 B.n400 71.676
R549 B.n406 B.n405 71.676
R550 B.n409 B.n408 71.676
R551 B.n225 B.n101 71.676
R552 B.n223 B.n103 71.676
R553 B.n219 B.n218 71.676
R554 B.n212 B.n105 71.676
R555 B.n211 B.n210 71.676
R556 B.n204 B.n107 71.676
R557 B.n203 B.n202 71.676
R558 B.n196 B.n109 71.676
R559 B.n195 B.n194 71.676
R560 B.n187 B.n111 71.676
R561 B.n186 B.n185 71.676
R562 B.n179 B.n115 71.676
R563 B.n178 B.n177 71.676
R564 B.n171 B.n117 71.676
R565 B.n170 B.n169 71.676
R566 B.n163 B.n119 71.676
R567 B.n162 B.n161 71.676
R568 B.n155 B.n124 71.676
R569 B.n154 B.n153 71.676
R570 B.n147 B.n126 71.676
R571 B.n146 B.n145 71.676
R572 B.n139 B.n128 71.676
R573 B.n138 B.n137 71.676
R574 B.n131 B.n130 71.676
R575 B.n226 B.n225 71.676
R576 B.n220 B.n103 71.676
R577 B.n218 B.n217 71.676
R578 B.n213 B.n212 71.676
R579 B.n210 B.n209 71.676
R580 B.n205 B.n204 71.676
R581 B.n202 B.n201 71.676
R582 B.n197 B.n196 71.676
R583 B.n194 B.n193 71.676
R584 B.n188 B.n187 71.676
R585 B.n185 B.n184 71.676
R586 B.n180 B.n179 71.676
R587 B.n177 B.n176 71.676
R588 B.n172 B.n171 71.676
R589 B.n169 B.n168 71.676
R590 B.n164 B.n163 71.676
R591 B.n161 B.n160 71.676
R592 B.n156 B.n155 71.676
R593 B.n153 B.n152 71.676
R594 B.n148 B.n147 71.676
R595 B.n145 B.n144 71.676
R596 B.n140 B.n139 71.676
R597 B.n137 B.n136 71.676
R598 B.n132 B.n131 71.676
R599 B.n451 B.n450 71.676
R600 B.n451 B.n2 71.676
R601 B.n56 B.t17 70.5728
R602 B.n121 B.t6 70.5728
R603 B.n50 B.t14 70.568
R604 B.n113 B.t9 70.568
R605 B.n282 B.t2 62.4196
R606 B.t1 B.n8 62.4196
R607 B.n371 B.n50 59.5399
R608 B.n57 B.n56 59.5399
R609 B.n122 B.n121 59.5399
R610 B.n190 B.n113 59.5399
R611 B.n261 B.t0 51.4689
R612 B.n19 B.t3 51.4689
R613 B.n229 B.n228 34.1859
R614 B.n233 B.n98 34.1859
R615 B.n311 B.n310 34.1859
R616 B.n412 B.n411 34.1859
R617 B.n268 B.t0 22.997
R618 B.n438 B.t3 22.997
R619 B.n50 B.n49 22.8853
R620 B.n56 B.n55 22.8853
R621 B.n121 B.n120 22.8853
R622 B.n113 B.n112 22.8853
R623 B B.n452 18.0485
R624 B.n275 B.t2 12.0463
R625 B.n12 B.t1 12.0463
R626 B.n229 B.n94 10.6151
R627 B.n239 B.n94 10.6151
R628 B.n240 B.n239 10.6151
R629 B.n241 B.n240 10.6151
R630 B.n241 B.n86 10.6151
R631 B.n251 B.n86 10.6151
R632 B.n252 B.n251 10.6151
R633 B.n253 B.n252 10.6151
R634 B.n253 B.n78 10.6151
R635 B.n264 B.n78 10.6151
R636 B.n265 B.n264 10.6151
R637 B.n266 B.n265 10.6151
R638 B.n266 B.n71 10.6151
R639 B.n278 B.n71 10.6151
R640 B.n279 B.n278 10.6151
R641 B.n280 B.n279 10.6151
R642 B.n280 B.n0 10.6151
R643 B.n228 B.n227 10.6151
R644 B.n227 B.n102 10.6151
R645 B.n222 B.n102 10.6151
R646 B.n222 B.n221 10.6151
R647 B.n221 B.n104 10.6151
R648 B.n216 B.n104 10.6151
R649 B.n216 B.n215 10.6151
R650 B.n215 B.n214 10.6151
R651 B.n214 B.n106 10.6151
R652 B.n208 B.n106 10.6151
R653 B.n208 B.n207 10.6151
R654 B.n207 B.n206 10.6151
R655 B.n206 B.n108 10.6151
R656 B.n200 B.n108 10.6151
R657 B.n200 B.n199 10.6151
R658 B.n199 B.n198 10.6151
R659 B.n198 B.n110 10.6151
R660 B.n192 B.n110 10.6151
R661 B.n192 B.n191 10.6151
R662 B.n189 B.n114 10.6151
R663 B.n183 B.n114 10.6151
R664 B.n183 B.n182 10.6151
R665 B.n182 B.n181 10.6151
R666 B.n181 B.n116 10.6151
R667 B.n175 B.n116 10.6151
R668 B.n175 B.n174 10.6151
R669 B.n174 B.n173 10.6151
R670 B.n173 B.n118 10.6151
R671 B.n167 B.n166 10.6151
R672 B.n166 B.n165 10.6151
R673 B.n165 B.n123 10.6151
R674 B.n159 B.n123 10.6151
R675 B.n159 B.n158 10.6151
R676 B.n158 B.n157 10.6151
R677 B.n157 B.n125 10.6151
R678 B.n151 B.n125 10.6151
R679 B.n151 B.n150 10.6151
R680 B.n150 B.n149 10.6151
R681 B.n149 B.n127 10.6151
R682 B.n143 B.n127 10.6151
R683 B.n143 B.n142 10.6151
R684 B.n142 B.n141 10.6151
R685 B.n141 B.n129 10.6151
R686 B.n135 B.n129 10.6151
R687 B.n135 B.n134 10.6151
R688 B.n134 B.n133 10.6151
R689 B.n133 B.n98 10.6151
R690 B.n234 B.n233 10.6151
R691 B.n235 B.n234 10.6151
R692 B.n235 B.n89 10.6151
R693 B.n245 B.n89 10.6151
R694 B.n246 B.n245 10.6151
R695 B.n247 B.n246 10.6151
R696 B.n247 B.n82 10.6151
R697 B.n257 B.n82 10.6151
R698 B.n258 B.n257 10.6151
R699 B.n259 B.n258 10.6151
R700 B.n259 B.n75 10.6151
R701 B.n270 B.n75 10.6151
R702 B.n271 B.n270 10.6151
R703 B.n273 B.n271 10.6151
R704 B.n273 B.n272 10.6151
R705 B.n272 B.n68 10.6151
R706 B.n285 B.n68 10.6151
R707 B.n286 B.n285 10.6151
R708 B.n287 B.n286 10.6151
R709 B.n288 B.n287 10.6151
R710 B.n289 B.n288 10.6151
R711 B.n292 B.n289 10.6151
R712 B.n293 B.n292 10.6151
R713 B.n294 B.n293 10.6151
R714 B.n295 B.n294 10.6151
R715 B.n297 B.n295 10.6151
R716 B.n298 B.n297 10.6151
R717 B.n299 B.n298 10.6151
R718 B.n300 B.n299 10.6151
R719 B.n302 B.n300 10.6151
R720 B.n303 B.n302 10.6151
R721 B.n304 B.n303 10.6151
R722 B.n305 B.n304 10.6151
R723 B.n307 B.n305 10.6151
R724 B.n308 B.n307 10.6151
R725 B.n309 B.n308 10.6151
R726 B.n310 B.n309 10.6151
R727 B.n444 B.n1 10.6151
R728 B.n444 B.n443 10.6151
R729 B.n443 B.n442 10.6151
R730 B.n442 B.n10 10.6151
R731 B.n436 B.n10 10.6151
R732 B.n436 B.n435 10.6151
R733 B.n435 B.n434 10.6151
R734 B.n434 B.n17 10.6151
R735 B.n428 B.n17 10.6151
R736 B.n428 B.n427 10.6151
R737 B.n427 B.n426 10.6151
R738 B.n426 B.n25 10.6151
R739 B.n420 B.n25 10.6151
R740 B.n420 B.n419 10.6151
R741 B.n419 B.n418 10.6151
R742 B.n418 B.n32 10.6151
R743 B.n412 B.n32 10.6151
R744 B.n411 B.n410 10.6151
R745 B.n410 B.n39 10.6151
R746 B.n404 B.n39 10.6151
R747 B.n404 B.n403 10.6151
R748 B.n403 B.n402 10.6151
R749 B.n402 B.n41 10.6151
R750 B.n396 B.n41 10.6151
R751 B.n396 B.n395 10.6151
R752 B.n395 B.n394 10.6151
R753 B.n394 B.n43 10.6151
R754 B.n388 B.n43 10.6151
R755 B.n388 B.n387 10.6151
R756 B.n387 B.n386 10.6151
R757 B.n386 B.n45 10.6151
R758 B.n380 B.n45 10.6151
R759 B.n380 B.n379 10.6151
R760 B.n379 B.n378 10.6151
R761 B.n378 B.n47 10.6151
R762 B.n372 B.n47 10.6151
R763 B.n370 B.n369 10.6151
R764 B.n369 B.n51 10.6151
R765 B.n363 B.n51 10.6151
R766 B.n363 B.n362 10.6151
R767 B.n362 B.n361 10.6151
R768 B.n361 B.n53 10.6151
R769 B.n355 B.n53 10.6151
R770 B.n355 B.n354 10.6151
R771 B.n354 B.n353 10.6151
R772 B.n349 B.n348 10.6151
R773 B.n348 B.n59 10.6151
R774 B.n343 B.n59 10.6151
R775 B.n343 B.n342 10.6151
R776 B.n342 B.n341 10.6151
R777 B.n341 B.n61 10.6151
R778 B.n335 B.n61 10.6151
R779 B.n335 B.n334 10.6151
R780 B.n334 B.n333 10.6151
R781 B.n333 B.n63 10.6151
R782 B.n327 B.n63 10.6151
R783 B.n327 B.n326 10.6151
R784 B.n326 B.n325 10.6151
R785 B.n325 B.n65 10.6151
R786 B.n319 B.n65 10.6151
R787 B.n319 B.n318 10.6151
R788 B.n318 B.n317 10.6151
R789 B.n317 B.n67 10.6151
R790 B.n311 B.n67 10.6151
R791 B.n191 B.n190 9.36635
R792 B.n167 B.n122 9.36635
R793 B.n372 B.n371 9.36635
R794 B.n349 B.n57 9.36635
R795 B.n452 B.n0 8.11757
R796 B.n452 B.n1 8.11757
R797 B.n190 B.n189 1.24928
R798 B.n122 B.n118 1.24928
R799 B.n371 B.n370 1.24928
R800 B.n353 B.n57 1.24928
R801 B.n92 B.t5 1.09557
R802 B.t12 B.n423 1.09557
R803 VP.n1 VP.t3 202.739
R804 VP.n1 VP.t1 202.69
R805 VP.n3 VP.t2 181.743
R806 VP.n5 VP.t0 181.743
R807 VP.n6 VP.n5 161.3
R808 VP.n4 VP.n0 161.3
R809 VP.n3 VP.n2 161.3
R810 VP.n2 VP.n1 80.1621
R811 VP.n4 VP.n3 24.1005
R812 VP.n5 VP.n4 24.1005
R813 VP.n2 VP.n0 0.189894
R814 VP.n6 VP.n0 0.189894
R815 VP VP.n6 0.0516364
R816 VDD1 VDD1.n1 103.934
R817 VDD1 VDD1.n0 72.5897
R818 VDD1.n0 VDD1.t0 4.15144
R819 VDD1.n0 VDD1.t2 4.15144
R820 VDD1.n1 VDD1.t1 4.15144
R821 VDD1.n1 VDD1.t3 4.15144
C0 VTAIL VP 1.54484f
C1 VP VN 3.58831f
C2 VDD1 VDD2 0.601115f
C3 VDD1 VTAIL 3.4606f
C4 VTAIL VDD2 3.50307f
C5 VDD1 VN 0.151088f
C6 VDD1 VP 1.68041f
C7 VDD2 VN 1.54519f
C8 VDD2 VP 0.286914f
C9 VTAIL VN 1.53073f
C10 VDD2 B 2.180634f
C11 VDD1 B 4.12043f
C12 VTAIL B 4.631189f
C13 VN B 6.09924f
C14 VP B 4.628176f
C15 VDD1.t0 B 0.070123f
C16 VDD1.t2 B 0.070123f
C17 VDD1.n0 B 0.575336f
C18 VDD1.t1 B 0.070123f
C19 VDD1.t3 B 0.070123f
C20 VDD1.n1 B 0.812079f
C21 VP.n0 B 0.026125f
C22 VP.t1 B 0.325815f
C23 VP.t3 B 0.325861f
C24 VP.n1 B 0.655656f
C25 VP.n2 B 1.30584f
C26 VP.t2 B 0.310126f
C27 VP.n3 B 0.149932f
C28 VP.n4 B 0.005928f
C29 VP.t0 B 0.310126f
C30 VP.n5 B 0.149932f
C31 VP.n6 B 0.020246f
C32 VTAIL.t7 B 0.481859f
C33 VTAIL.n0 B 0.185659f
C34 VTAIL.t2 B 0.481859f
C35 VTAIL.n1 B 0.204778f
C36 VTAIL.t0 B 0.481859f
C37 VTAIL.n2 B 0.581503f
C38 VTAIL.t6 B 0.48186f
C39 VTAIL.n3 B 0.581503f
C40 VTAIL.t4 B 0.48186f
C41 VTAIL.n4 B 0.204778f
C42 VTAIL.t1 B 0.48186f
C43 VTAIL.n5 B 0.204778f
C44 VTAIL.t3 B 0.481858f
C45 VTAIL.n6 B 0.581505f
C46 VTAIL.t5 B 0.481859f
C47 VTAIL.n7 B 0.557444f
C48 VDD2.t3 B 0.071527f
C49 VDD2.t2 B 0.071527f
C50 VDD2.n0 B 0.813857f
C51 VDD2.t0 B 0.071527f
C52 VDD2.t1 B 0.071527f
C53 VDD2.n1 B 0.586684f
C54 VDD2.n2 B 1.74707f
C55 VN.t0 B 0.32257f
C56 VN.t2 B 0.322525f
C57 VN.n0 B 0.271882f
C58 VN.t3 B 0.32257f
C59 VN.t1 B 0.322525f
C60 VN.n1 B 0.658927f
.ends

