* NGSPICE file created from diff_pair_sample_0819.ext - technology: sky130A

.subckt diff_pair_sample_0819 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t2 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=1.1187 ps=7.11 w=6.78 l=1.07
X1 VTAIL.t1 VN.t0 VDD2.t5 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=1.1187 ps=7.11 w=6.78 l=1.07
X2 VDD1.t4 VP.t1 VTAIL.t5 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=1.1187 ps=7.11 w=6.78 l=1.07
X3 VDD2.t4 VN.t1 VTAIL.t0 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=1.1187 ps=7.11 w=6.78 l=1.07
X4 VDD1.t3 VP.t2 VTAIL.t7 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=2.6442 ps=14.34 w=6.78 l=1.07
X5 VDD2.t3 VN.t2 VTAIL.t8 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=2.6442 ps=14.34 w=6.78 l=1.07
X6 VTAIL.t9 VN.t3 VDD2.t2 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=1.1187 ps=7.11 w=6.78 l=1.07
X7 B.t11 B.t9 B.t10 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=0 ps=0 w=6.78 l=1.07
X8 VDD1.t2 VP.t3 VTAIL.t3 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=2.6442 ps=14.34 w=6.78 l=1.07
X9 VDD2.t1 VN.t4 VTAIL.t10 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=1.1187 ps=7.11 w=6.78 l=1.07
X10 VDD2.t0 VN.t5 VTAIL.t11 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=2.6442 ps=14.34 w=6.78 l=1.07
X11 VTAIL.t4 VP.t4 VDD1.t1 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=1.1187 ps=7.11 w=6.78 l=1.07
X12 B.t8 B.t6 B.t7 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=0 ps=0 w=6.78 l=1.07
X13 VTAIL.t6 VP.t5 VDD1.t0 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=1.1187 pd=7.11 as=1.1187 ps=7.11 w=6.78 l=1.07
X14 B.t5 B.t3 B.t4 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=0 ps=0 w=6.78 l=1.07
X15 B.t2 B.t0 B.t1 w_n2090_n2324# sky130_fd_pr__pfet_01v8 ad=2.6442 pd=14.34 as=0 ps=0 w=6.78 l=1.07
R0 VP.n3 VP.t1 212.304
R1 VP.n8 VP.t0 189.422
R2 VP.n14 VP.t3 189.422
R3 VP.n6 VP.t2 189.422
R4 VP.n5 VP.n2 161.3
R5 VP.n13 VP.n0 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n1 161.3
R8 VP.n12 VP.t5 152.708
R9 VP.n4 VP.t4 152.708
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 49.9219
R14 VP.n14 VP.n13 49.9219
R15 VP.n6 VP.n5 49.9219
R16 VP.n9 VP.n7 38.8802
R17 VP.n4 VP.n3 32.5705
R18 VP.n3 VP.n2 28.1996
R19 VP.n12 VP.n1 24.5923
R20 VP.n13 VP.n12 24.5923
R21 VP.n5 VP.n4 24.5923
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n146 VTAIL.n116 756.745
R29 VTAIL.n32 VTAIL.n2 756.745
R30 VTAIL.n110 VTAIL.n80 756.745
R31 VTAIL.n72 VTAIL.n42 756.745
R32 VTAIL.n129 VTAIL.n128 585
R33 VTAIL.n131 VTAIL.n130 585
R34 VTAIL.n124 VTAIL.n123 585
R35 VTAIL.n137 VTAIL.n136 585
R36 VTAIL.n139 VTAIL.n138 585
R37 VTAIL.n120 VTAIL.n119 585
R38 VTAIL.n145 VTAIL.n144 585
R39 VTAIL.n147 VTAIL.n146 585
R40 VTAIL.n15 VTAIL.n14 585
R41 VTAIL.n17 VTAIL.n16 585
R42 VTAIL.n10 VTAIL.n9 585
R43 VTAIL.n23 VTAIL.n22 585
R44 VTAIL.n25 VTAIL.n24 585
R45 VTAIL.n6 VTAIL.n5 585
R46 VTAIL.n31 VTAIL.n30 585
R47 VTAIL.n33 VTAIL.n32 585
R48 VTAIL.n111 VTAIL.n110 585
R49 VTAIL.n109 VTAIL.n108 585
R50 VTAIL.n84 VTAIL.n83 585
R51 VTAIL.n103 VTAIL.n102 585
R52 VTAIL.n101 VTAIL.n100 585
R53 VTAIL.n88 VTAIL.n87 585
R54 VTAIL.n95 VTAIL.n94 585
R55 VTAIL.n93 VTAIL.n92 585
R56 VTAIL.n73 VTAIL.n72 585
R57 VTAIL.n71 VTAIL.n70 585
R58 VTAIL.n46 VTAIL.n45 585
R59 VTAIL.n65 VTAIL.n64 585
R60 VTAIL.n63 VTAIL.n62 585
R61 VTAIL.n50 VTAIL.n49 585
R62 VTAIL.n57 VTAIL.n56 585
R63 VTAIL.n55 VTAIL.n54 585
R64 VTAIL.n127 VTAIL.t11 327.514
R65 VTAIL.n13 VTAIL.t3 327.514
R66 VTAIL.n91 VTAIL.t7 327.514
R67 VTAIL.n53 VTAIL.t8 327.514
R68 VTAIL.n130 VTAIL.n129 171.744
R69 VTAIL.n130 VTAIL.n123 171.744
R70 VTAIL.n137 VTAIL.n123 171.744
R71 VTAIL.n138 VTAIL.n137 171.744
R72 VTAIL.n138 VTAIL.n119 171.744
R73 VTAIL.n145 VTAIL.n119 171.744
R74 VTAIL.n146 VTAIL.n145 171.744
R75 VTAIL.n16 VTAIL.n15 171.744
R76 VTAIL.n16 VTAIL.n9 171.744
R77 VTAIL.n23 VTAIL.n9 171.744
R78 VTAIL.n24 VTAIL.n23 171.744
R79 VTAIL.n24 VTAIL.n5 171.744
R80 VTAIL.n31 VTAIL.n5 171.744
R81 VTAIL.n32 VTAIL.n31 171.744
R82 VTAIL.n110 VTAIL.n109 171.744
R83 VTAIL.n109 VTAIL.n83 171.744
R84 VTAIL.n102 VTAIL.n83 171.744
R85 VTAIL.n102 VTAIL.n101 171.744
R86 VTAIL.n101 VTAIL.n87 171.744
R87 VTAIL.n94 VTAIL.n87 171.744
R88 VTAIL.n94 VTAIL.n93 171.744
R89 VTAIL.n72 VTAIL.n71 171.744
R90 VTAIL.n71 VTAIL.n45 171.744
R91 VTAIL.n64 VTAIL.n45 171.744
R92 VTAIL.n64 VTAIL.n63 171.744
R93 VTAIL.n63 VTAIL.n49 171.744
R94 VTAIL.n56 VTAIL.n49 171.744
R95 VTAIL.n56 VTAIL.n55 171.744
R96 VTAIL.n129 VTAIL.t11 85.8723
R97 VTAIL.n15 VTAIL.t3 85.8723
R98 VTAIL.n93 VTAIL.t7 85.8723
R99 VTAIL.n55 VTAIL.t8 85.8723
R100 VTAIL.n79 VTAIL.n78 72.8838
R101 VTAIL.n41 VTAIL.n40 72.8838
R102 VTAIL.n1 VTAIL.n0 72.8836
R103 VTAIL.n39 VTAIL.n38 72.8836
R104 VTAIL.n151 VTAIL.n150 33.349
R105 VTAIL.n37 VTAIL.n36 33.349
R106 VTAIL.n115 VTAIL.n114 33.349
R107 VTAIL.n77 VTAIL.n76 33.349
R108 VTAIL.n41 VTAIL.n39 20.6255
R109 VTAIL.n151 VTAIL.n115 19.4186
R110 VTAIL.n128 VTAIL.n127 16.3884
R111 VTAIL.n14 VTAIL.n13 16.3884
R112 VTAIL.n92 VTAIL.n91 16.3884
R113 VTAIL.n54 VTAIL.n53 16.3884
R114 VTAIL.n131 VTAIL.n126 12.8005
R115 VTAIL.n17 VTAIL.n12 12.8005
R116 VTAIL.n95 VTAIL.n90 12.8005
R117 VTAIL.n57 VTAIL.n52 12.8005
R118 VTAIL.n132 VTAIL.n124 12.0247
R119 VTAIL.n18 VTAIL.n10 12.0247
R120 VTAIL.n96 VTAIL.n88 12.0247
R121 VTAIL.n58 VTAIL.n50 12.0247
R122 VTAIL.n136 VTAIL.n135 11.249
R123 VTAIL.n22 VTAIL.n21 11.249
R124 VTAIL.n100 VTAIL.n99 11.249
R125 VTAIL.n62 VTAIL.n61 11.249
R126 VTAIL.n139 VTAIL.n122 10.4732
R127 VTAIL.n25 VTAIL.n8 10.4732
R128 VTAIL.n103 VTAIL.n86 10.4732
R129 VTAIL.n65 VTAIL.n48 10.4732
R130 VTAIL.n140 VTAIL.n120 9.69747
R131 VTAIL.n26 VTAIL.n6 9.69747
R132 VTAIL.n104 VTAIL.n84 9.69747
R133 VTAIL.n66 VTAIL.n46 9.69747
R134 VTAIL.n150 VTAIL.n149 9.45567
R135 VTAIL.n36 VTAIL.n35 9.45567
R136 VTAIL.n114 VTAIL.n113 9.45567
R137 VTAIL.n76 VTAIL.n75 9.45567
R138 VTAIL.n118 VTAIL.n117 9.3005
R139 VTAIL.n143 VTAIL.n142 9.3005
R140 VTAIL.n141 VTAIL.n140 9.3005
R141 VTAIL.n122 VTAIL.n121 9.3005
R142 VTAIL.n135 VTAIL.n134 9.3005
R143 VTAIL.n133 VTAIL.n132 9.3005
R144 VTAIL.n126 VTAIL.n125 9.3005
R145 VTAIL.n149 VTAIL.n148 9.3005
R146 VTAIL.n4 VTAIL.n3 9.3005
R147 VTAIL.n29 VTAIL.n28 9.3005
R148 VTAIL.n27 VTAIL.n26 9.3005
R149 VTAIL.n8 VTAIL.n7 9.3005
R150 VTAIL.n21 VTAIL.n20 9.3005
R151 VTAIL.n19 VTAIL.n18 9.3005
R152 VTAIL.n12 VTAIL.n11 9.3005
R153 VTAIL.n35 VTAIL.n34 9.3005
R154 VTAIL.n113 VTAIL.n112 9.3005
R155 VTAIL.n82 VTAIL.n81 9.3005
R156 VTAIL.n107 VTAIL.n106 9.3005
R157 VTAIL.n105 VTAIL.n104 9.3005
R158 VTAIL.n86 VTAIL.n85 9.3005
R159 VTAIL.n99 VTAIL.n98 9.3005
R160 VTAIL.n97 VTAIL.n96 9.3005
R161 VTAIL.n90 VTAIL.n89 9.3005
R162 VTAIL.n75 VTAIL.n74 9.3005
R163 VTAIL.n44 VTAIL.n43 9.3005
R164 VTAIL.n69 VTAIL.n68 9.3005
R165 VTAIL.n67 VTAIL.n66 9.3005
R166 VTAIL.n48 VTAIL.n47 9.3005
R167 VTAIL.n61 VTAIL.n60 9.3005
R168 VTAIL.n59 VTAIL.n58 9.3005
R169 VTAIL.n52 VTAIL.n51 9.3005
R170 VTAIL.n144 VTAIL.n143 8.92171
R171 VTAIL.n30 VTAIL.n29 8.92171
R172 VTAIL.n108 VTAIL.n107 8.92171
R173 VTAIL.n70 VTAIL.n69 8.92171
R174 VTAIL.n147 VTAIL.n118 8.14595
R175 VTAIL.n33 VTAIL.n4 8.14595
R176 VTAIL.n111 VTAIL.n82 8.14595
R177 VTAIL.n73 VTAIL.n44 8.14595
R178 VTAIL.n148 VTAIL.n116 7.3702
R179 VTAIL.n34 VTAIL.n2 7.3702
R180 VTAIL.n112 VTAIL.n80 7.3702
R181 VTAIL.n74 VTAIL.n42 7.3702
R182 VTAIL.n150 VTAIL.n116 6.59444
R183 VTAIL.n36 VTAIL.n2 6.59444
R184 VTAIL.n114 VTAIL.n80 6.59444
R185 VTAIL.n76 VTAIL.n42 6.59444
R186 VTAIL.n148 VTAIL.n147 5.81868
R187 VTAIL.n34 VTAIL.n33 5.81868
R188 VTAIL.n112 VTAIL.n111 5.81868
R189 VTAIL.n74 VTAIL.n73 5.81868
R190 VTAIL.n144 VTAIL.n118 5.04292
R191 VTAIL.n30 VTAIL.n4 5.04292
R192 VTAIL.n108 VTAIL.n82 5.04292
R193 VTAIL.n70 VTAIL.n44 5.04292
R194 VTAIL.n0 VTAIL.t0 4.79475
R195 VTAIL.n0 VTAIL.t9 4.79475
R196 VTAIL.n38 VTAIL.t2 4.79475
R197 VTAIL.n38 VTAIL.t6 4.79475
R198 VTAIL.n78 VTAIL.t5 4.79475
R199 VTAIL.n78 VTAIL.t4 4.79475
R200 VTAIL.n40 VTAIL.t10 4.79475
R201 VTAIL.n40 VTAIL.t1 4.79475
R202 VTAIL.n143 VTAIL.n120 4.26717
R203 VTAIL.n29 VTAIL.n6 4.26717
R204 VTAIL.n107 VTAIL.n84 4.26717
R205 VTAIL.n69 VTAIL.n46 4.26717
R206 VTAIL.n127 VTAIL.n125 3.71088
R207 VTAIL.n13 VTAIL.n11 3.71088
R208 VTAIL.n91 VTAIL.n89 3.71088
R209 VTAIL.n53 VTAIL.n51 3.71088
R210 VTAIL.n140 VTAIL.n139 3.49141
R211 VTAIL.n26 VTAIL.n25 3.49141
R212 VTAIL.n104 VTAIL.n103 3.49141
R213 VTAIL.n66 VTAIL.n65 3.49141
R214 VTAIL.n136 VTAIL.n122 2.71565
R215 VTAIL.n22 VTAIL.n8 2.71565
R216 VTAIL.n100 VTAIL.n86 2.71565
R217 VTAIL.n62 VTAIL.n48 2.71565
R218 VTAIL.n135 VTAIL.n124 1.93989
R219 VTAIL.n21 VTAIL.n10 1.93989
R220 VTAIL.n99 VTAIL.n88 1.93989
R221 VTAIL.n61 VTAIL.n50 1.93989
R222 VTAIL.n77 VTAIL.n41 1.2074
R223 VTAIL.n115 VTAIL.n79 1.2074
R224 VTAIL.n39 VTAIL.n37 1.2074
R225 VTAIL.n132 VTAIL.n131 1.16414
R226 VTAIL.n18 VTAIL.n17 1.16414
R227 VTAIL.n96 VTAIL.n95 1.16414
R228 VTAIL.n58 VTAIL.n57 1.16414
R229 VTAIL.n79 VTAIL.n77 1.07378
R230 VTAIL.n37 VTAIL.n1 1.07378
R231 VTAIL VTAIL.n151 0.847483
R232 VTAIL.n128 VTAIL.n126 0.388379
R233 VTAIL.n14 VTAIL.n12 0.388379
R234 VTAIL.n92 VTAIL.n90 0.388379
R235 VTAIL.n54 VTAIL.n52 0.388379
R236 VTAIL VTAIL.n1 0.360414
R237 VTAIL.n133 VTAIL.n125 0.155672
R238 VTAIL.n134 VTAIL.n133 0.155672
R239 VTAIL.n134 VTAIL.n121 0.155672
R240 VTAIL.n141 VTAIL.n121 0.155672
R241 VTAIL.n142 VTAIL.n141 0.155672
R242 VTAIL.n142 VTAIL.n117 0.155672
R243 VTAIL.n149 VTAIL.n117 0.155672
R244 VTAIL.n19 VTAIL.n11 0.155672
R245 VTAIL.n20 VTAIL.n19 0.155672
R246 VTAIL.n20 VTAIL.n7 0.155672
R247 VTAIL.n27 VTAIL.n7 0.155672
R248 VTAIL.n28 VTAIL.n27 0.155672
R249 VTAIL.n28 VTAIL.n3 0.155672
R250 VTAIL.n35 VTAIL.n3 0.155672
R251 VTAIL.n113 VTAIL.n81 0.155672
R252 VTAIL.n106 VTAIL.n81 0.155672
R253 VTAIL.n106 VTAIL.n105 0.155672
R254 VTAIL.n105 VTAIL.n85 0.155672
R255 VTAIL.n98 VTAIL.n85 0.155672
R256 VTAIL.n98 VTAIL.n97 0.155672
R257 VTAIL.n97 VTAIL.n89 0.155672
R258 VTAIL.n75 VTAIL.n43 0.155672
R259 VTAIL.n68 VTAIL.n43 0.155672
R260 VTAIL.n68 VTAIL.n67 0.155672
R261 VTAIL.n67 VTAIL.n47 0.155672
R262 VTAIL.n60 VTAIL.n47 0.155672
R263 VTAIL.n60 VTAIL.n59 0.155672
R264 VTAIL.n59 VTAIL.n51 0.155672
R265 VDD1.n30 VDD1.n0 756.745
R266 VDD1.n65 VDD1.n35 756.745
R267 VDD1.n31 VDD1.n30 585
R268 VDD1.n29 VDD1.n28 585
R269 VDD1.n4 VDD1.n3 585
R270 VDD1.n23 VDD1.n22 585
R271 VDD1.n21 VDD1.n20 585
R272 VDD1.n8 VDD1.n7 585
R273 VDD1.n15 VDD1.n14 585
R274 VDD1.n13 VDD1.n12 585
R275 VDD1.n48 VDD1.n47 585
R276 VDD1.n50 VDD1.n49 585
R277 VDD1.n43 VDD1.n42 585
R278 VDD1.n56 VDD1.n55 585
R279 VDD1.n58 VDD1.n57 585
R280 VDD1.n39 VDD1.n38 585
R281 VDD1.n64 VDD1.n63 585
R282 VDD1.n66 VDD1.n65 585
R283 VDD1.n11 VDD1.t4 327.514
R284 VDD1.n46 VDD1.t5 327.514
R285 VDD1.n30 VDD1.n29 171.744
R286 VDD1.n29 VDD1.n3 171.744
R287 VDD1.n22 VDD1.n3 171.744
R288 VDD1.n22 VDD1.n21 171.744
R289 VDD1.n21 VDD1.n7 171.744
R290 VDD1.n14 VDD1.n7 171.744
R291 VDD1.n14 VDD1.n13 171.744
R292 VDD1.n49 VDD1.n48 171.744
R293 VDD1.n49 VDD1.n42 171.744
R294 VDD1.n56 VDD1.n42 171.744
R295 VDD1.n57 VDD1.n56 171.744
R296 VDD1.n57 VDD1.n38 171.744
R297 VDD1.n64 VDD1.n38 171.744
R298 VDD1.n65 VDD1.n64 171.744
R299 VDD1.n71 VDD1.n70 89.8088
R300 VDD1.n73 VDD1.n72 89.5624
R301 VDD1.n13 VDD1.t4 85.8723
R302 VDD1.n48 VDD1.t5 85.8723
R303 VDD1 VDD1.n34 50.9911
R304 VDD1.n71 VDD1.n69 50.8776
R305 VDD1.n73 VDD1.n71 34.669
R306 VDD1.n47 VDD1.n46 16.3884
R307 VDD1.n12 VDD1.n11 16.3884
R308 VDD1.n15 VDD1.n10 12.8005
R309 VDD1.n50 VDD1.n45 12.8005
R310 VDD1.n16 VDD1.n8 12.0247
R311 VDD1.n51 VDD1.n43 12.0247
R312 VDD1.n20 VDD1.n19 11.249
R313 VDD1.n55 VDD1.n54 11.249
R314 VDD1.n23 VDD1.n6 10.4732
R315 VDD1.n58 VDD1.n41 10.4732
R316 VDD1.n24 VDD1.n4 9.69747
R317 VDD1.n59 VDD1.n39 9.69747
R318 VDD1.n34 VDD1.n33 9.45567
R319 VDD1.n69 VDD1.n68 9.45567
R320 VDD1.n33 VDD1.n32 9.3005
R321 VDD1.n2 VDD1.n1 9.3005
R322 VDD1.n27 VDD1.n26 9.3005
R323 VDD1.n25 VDD1.n24 9.3005
R324 VDD1.n6 VDD1.n5 9.3005
R325 VDD1.n19 VDD1.n18 9.3005
R326 VDD1.n17 VDD1.n16 9.3005
R327 VDD1.n10 VDD1.n9 9.3005
R328 VDD1.n37 VDD1.n36 9.3005
R329 VDD1.n62 VDD1.n61 9.3005
R330 VDD1.n60 VDD1.n59 9.3005
R331 VDD1.n41 VDD1.n40 9.3005
R332 VDD1.n54 VDD1.n53 9.3005
R333 VDD1.n52 VDD1.n51 9.3005
R334 VDD1.n45 VDD1.n44 9.3005
R335 VDD1.n68 VDD1.n67 9.3005
R336 VDD1.n28 VDD1.n27 8.92171
R337 VDD1.n63 VDD1.n62 8.92171
R338 VDD1.n31 VDD1.n2 8.14595
R339 VDD1.n66 VDD1.n37 8.14595
R340 VDD1.n32 VDD1.n0 7.3702
R341 VDD1.n67 VDD1.n35 7.3702
R342 VDD1.n34 VDD1.n0 6.59444
R343 VDD1.n69 VDD1.n35 6.59444
R344 VDD1.n32 VDD1.n31 5.81868
R345 VDD1.n67 VDD1.n66 5.81868
R346 VDD1.n28 VDD1.n2 5.04292
R347 VDD1.n63 VDD1.n37 5.04292
R348 VDD1.n72 VDD1.t1 4.79475
R349 VDD1.n72 VDD1.t3 4.79475
R350 VDD1.n70 VDD1.t0 4.79475
R351 VDD1.n70 VDD1.t2 4.79475
R352 VDD1.n27 VDD1.n4 4.26717
R353 VDD1.n62 VDD1.n39 4.26717
R354 VDD1.n11 VDD1.n9 3.71088
R355 VDD1.n46 VDD1.n44 3.71088
R356 VDD1.n24 VDD1.n23 3.49141
R357 VDD1.n59 VDD1.n58 3.49141
R358 VDD1.n20 VDD1.n6 2.71565
R359 VDD1.n55 VDD1.n41 2.71565
R360 VDD1.n19 VDD1.n8 1.93989
R361 VDD1.n54 VDD1.n43 1.93989
R362 VDD1.n16 VDD1.n15 1.16414
R363 VDD1.n51 VDD1.n50 1.16414
R364 VDD1.n12 VDD1.n10 0.388379
R365 VDD1.n47 VDD1.n45 0.388379
R366 VDD1 VDD1.n73 0.244034
R367 VDD1.n33 VDD1.n1 0.155672
R368 VDD1.n26 VDD1.n1 0.155672
R369 VDD1.n26 VDD1.n25 0.155672
R370 VDD1.n25 VDD1.n5 0.155672
R371 VDD1.n18 VDD1.n5 0.155672
R372 VDD1.n18 VDD1.n17 0.155672
R373 VDD1.n17 VDD1.n9 0.155672
R374 VDD1.n52 VDD1.n44 0.155672
R375 VDD1.n53 VDD1.n52 0.155672
R376 VDD1.n53 VDD1.n40 0.155672
R377 VDD1.n60 VDD1.n40 0.155672
R378 VDD1.n61 VDD1.n60 0.155672
R379 VDD1.n61 VDD1.n36 0.155672
R380 VDD1.n68 VDD1.n36 0.155672
R381 VN.n1 VN.t1 212.304
R382 VN.n7 VN.t2 212.304
R383 VN.n4 VN.t5 189.422
R384 VN.n10 VN.t4 189.422
R385 VN.n9 VN.n6 161.3
R386 VN.n3 VN.n0 161.3
R387 VN.n2 VN.t3 152.708
R388 VN.n8 VN.t0 152.708
R389 VN.n11 VN.n10 80.6037
R390 VN.n5 VN.n4 80.6037
R391 VN.n4 VN.n3 49.9219
R392 VN.n10 VN.n9 49.9219
R393 VN VN.n11 39.1657
R394 VN.n2 VN.n1 32.5705
R395 VN.n8 VN.n7 32.5705
R396 VN.n7 VN.n6 28.1996
R397 VN.n1 VN.n0 28.1996
R398 VN.n3 VN.n2 24.5923
R399 VN.n9 VN.n8 24.5923
R400 VN.n11 VN.n6 0.285035
R401 VN.n5 VN.n0 0.285035
R402 VN VN.n5 0.146778
R403 VDD2.n67 VDD2.n37 756.745
R404 VDD2.n30 VDD2.n0 756.745
R405 VDD2.n68 VDD2.n67 585
R406 VDD2.n66 VDD2.n65 585
R407 VDD2.n41 VDD2.n40 585
R408 VDD2.n60 VDD2.n59 585
R409 VDD2.n58 VDD2.n57 585
R410 VDD2.n45 VDD2.n44 585
R411 VDD2.n52 VDD2.n51 585
R412 VDD2.n50 VDD2.n49 585
R413 VDD2.n13 VDD2.n12 585
R414 VDD2.n15 VDD2.n14 585
R415 VDD2.n8 VDD2.n7 585
R416 VDD2.n21 VDD2.n20 585
R417 VDD2.n23 VDD2.n22 585
R418 VDD2.n4 VDD2.n3 585
R419 VDD2.n29 VDD2.n28 585
R420 VDD2.n31 VDD2.n30 585
R421 VDD2.n48 VDD2.t1 327.514
R422 VDD2.n11 VDD2.t4 327.514
R423 VDD2.n67 VDD2.n66 171.744
R424 VDD2.n66 VDD2.n40 171.744
R425 VDD2.n59 VDD2.n40 171.744
R426 VDD2.n59 VDD2.n58 171.744
R427 VDD2.n58 VDD2.n44 171.744
R428 VDD2.n51 VDD2.n44 171.744
R429 VDD2.n51 VDD2.n50 171.744
R430 VDD2.n14 VDD2.n13 171.744
R431 VDD2.n14 VDD2.n7 171.744
R432 VDD2.n21 VDD2.n7 171.744
R433 VDD2.n22 VDD2.n21 171.744
R434 VDD2.n22 VDD2.n3 171.744
R435 VDD2.n29 VDD2.n3 171.744
R436 VDD2.n30 VDD2.n29 171.744
R437 VDD2.n36 VDD2.n35 89.8088
R438 VDD2 VDD2.n73 89.806
R439 VDD2.n50 VDD2.t1 85.8723
R440 VDD2.n13 VDD2.t4 85.8723
R441 VDD2.n36 VDD2.n34 50.8776
R442 VDD2.n72 VDD2.n71 50.0278
R443 VDD2.n72 VDD2.n36 33.4825
R444 VDD2.n12 VDD2.n11 16.3884
R445 VDD2.n49 VDD2.n48 16.3884
R446 VDD2.n52 VDD2.n47 12.8005
R447 VDD2.n15 VDD2.n10 12.8005
R448 VDD2.n53 VDD2.n45 12.0247
R449 VDD2.n16 VDD2.n8 12.0247
R450 VDD2.n57 VDD2.n56 11.249
R451 VDD2.n20 VDD2.n19 11.249
R452 VDD2.n60 VDD2.n43 10.4732
R453 VDD2.n23 VDD2.n6 10.4732
R454 VDD2.n61 VDD2.n41 9.69747
R455 VDD2.n24 VDD2.n4 9.69747
R456 VDD2.n71 VDD2.n70 9.45567
R457 VDD2.n34 VDD2.n33 9.45567
R458 VDD2.n70 VDD2.n69 9.3005
R459 VDD2.n39 VDD2.n38 9.3005
R460 VDD2.n64 VDD2.n63 9.3005
R461 VDD2.n62 VDD2.n61 9.3005
R462 VDD2.n43 VDD2.n42 9.3005
R463 VDD2.n56 VDD2.n55 9.3005
R464 VDD2.n54 VDD2.n53 9.3005
R465 VDD2.n47 VDD2.n46 9.3005
R466 VDD2.n2 VDD2.n1 9.3005
R467 VDD2.n27 VDD2.n26 9.3005
R468 VDD2.n25 VDD2.n24 9.3005
R469 VDD2.n6 VDD2.n5 9.3005
R470 VDD2.n19 VDD2.n18 9.3005
R471 VDD2.n17 VDD2.n16 9.3005
R472 VDD2.n10 VDD2.n9 9.3005
R473 VDD2.n33 VDD2.n32 9.3005
R474 VDD2.n65 VDD2.n64 8.92171
R475 VDD2.n28 VDD2.n27 8.92171
R476 VDD2.n68 VDD2.n39 8.14595
R477 VDD2.n31 VDD2.n2 8.14595
R478 VDD2.n69 VDD2.n37 7.3702
R479 VDD2.n32 VDD2.n0 7.3702
R480 VDD2.n71 VDD2.n37 6.59444
R481 VDD2.n34 VDD2.n0 6.59444
R482 VDD2.n69 VDD2.n68 5.81868
R483 VDD2.n32 VDD2.n31 5.81868
R484 VDD2.n65 VDD2.n39 5.04292
R485 VDD2.n28 VDD2.n2 5.04292
R486 VDD2.n73 VDD2.t5 4.79475
R487 VDD2.n73 VDD2.t3 4.79475
R488 VDD2.n35 VDD2.t2 4.79475
R489 VDD2.n35 VDD2.t0 4.79475
R490 VDD2.n64 VDD2.n41 4.26717
R491 VDD2.n27 VDD2.n4 4.26717
R492 VDD2.n48 VDD2.n46 3.71088
R493 VDD2.n11 VDD2.n9 3.71088
R494 VDD2.n61 VDD2.n60 3.49141
R495 VDD2.n24 VDD2.n23 3.49141
R496 VDD2.n57 VDD2.n43 2.71565
R497 VDD2.n20 VDD2.n6 2.71565
R498 VDD2.n56 VDD2.n45 1.93989
R499 VDD2.n19 VDD2.n8 1.93989
R500 VDD2.n53 VDD2.n52 1.16414
R501 VDD2.n16 VDD2.n15 1.16414
R502 VDD2 VDD2.n72 0.963862
R503 VDD2.n49 VDD2.n47 0.388379
R504 VDD2.n12 VDD2.n10 0.388379
R505 VDD2.n70 VDD2.n38 0.155672
R506 VDD2.n63 VDD2.n38 0.155672
R507 VDD2.n63 VDD2.n62 0.155672
R508 VDD2.n62 VDD2.n42 0.155672
R509 VDD2.n55 VDD2.n42 0.155672
R510 VDD2.n55 VDD2.n54 0.155672
R511 VDD2.n54 VDD2.n46 0.155672
R512 VDD2.n17 VDD2.n9 0.155672
R513 VDD2.n18 VDD2.n17 0.155672
R514 VDD2.n18 VDD2.n5 0.155672
R515 VDD2.n25 VDD2.n5 0.155672
R516 VDD2.n26 VDD2.n25 0.155672
R517 VDD2.n26 VDD2.n1 0.155672
R518 VDD2.n33 VDD2.n1 0.155672
R519 B.n250 B.n249 585
R520 B.n248 B.n75 585
R521 B.n247 B.n246 585
R522 B.n245 B.n76 585
R523 B.n244 B.n243 585
R524 B.n242 B.n77 585
R525 B.n241 B.n240 585
R526 B.n239 B.n78 585
R527 B.n238 B.n237 585
R528 B.n236 B.n79 585
R529 B.n235 B.n234 585
R530 B.n233 B.n80 585
R531 B.n232 B.n231 585
R532 B.n230 B.n81 585
R533 B.n229 B.n228 585
R534 B.n227 B.n82 585
R535 B.n226 B.n225 585
R536 B.n224 B.n83 585
R537 B.n223 B.n222 585
R538 B.n221 B.n84 585
R539 B.n220 B.n219 585
R540 B.n218 B.n85 585
R541 B.n217 B.n216 585
R542 B.n215 B.n86 585
R543 B.n214 B.n213 585
R544 B.n212 B.n87 585
R545 B.n210 B.n209 585
R546 B.n208 B.n90 585
R547 B.n207 B.n206 585
R548 B.n205 B.n91 585
R549 B.n204 B.n203 585
R550 B.n202 B.n92 585
R551 B.n201 B.n200 585
R552 B.n199 B.n93 585
R553 B.n198 B.n197 585
R554 B.n196 B.n94 585
R555 B.n195 B.n194 585
R556 B.n190 B.n95 585
R557 B.n189 B.n188 585
R558 B.n187 B.n96 585
R559 B.n186 B.n185 585
R560 B.n184 B.n97 585
R561 B.n183 B.n182 585
R562 B.n181 B.n98 585
R563 B.n180 B.n179 585
R564 B.n178 B.n99 585
R565 B.n177 B.n176 585
R566 B.n175 B.n100 585
R567 B.n174 B.n173 585
R568 B.n172 B.n101 585
R569 B.n171 B.n170 585
R570 B.n169 B.n102 585
R571 B.n168 B.n167 585
R572 B.n166 B.n103 585
R573 B.n165 B.n164 585
R574 B.n163 B.n104 585
R575 B.n162 B.n161 585
R576 B.n160 B.n105 585
R577 B.n159 B.n158 585
R578 B.n157 B.n106 585
R579 B.n156 B.n155 585
R580 B.n154 B.n107 585
R581 B.n251 B.n74 585
R582 B.n253 B.n252 585
R583 B.n254 B.n73 585
R584 B.n256 B.n255 585
R585 B.n257 B.n72 585
R586 B.n259 B.n258 585
R587 B.n260 B.n71 585
R588 B.n262 B.n261 585
R589 B.n263 B.n70 585
R590 B.n265 B.n264 585
R591 B.n266 B.n69 585
R592 B.n268 B.n267 585
R593 B.n269 B.n68 585
R594 B.n271 B.n270 585
R595 B.n272 B.n67 585
R596 B.n274 B.n273 585
R597 B.n275 B.n66 585
R598 B.n277 B.n276 585
R599 B.n278 B.n65 585
R600 B.n280 B.n279 585
R601 B.n281 B.n64 585
R602 B.n283 B.n282 585
R603 B.n284 B.n63 585
R604 B.n286 B.n285 585
R605 B.n287 B.n62 585
R606 B.n289 B.n288 585
R607 B.n290 B.n61 585
R608 B.n292 B.n291 585
R609 B.n293 B.n60 585
R610 B.n295 B.n294 585
R611 B.n296 B.n59 585
R612 B.n298 B.n297 585
R613 B.n299 B.n58 585
R614 B.n301 B.n300 585
R615 B.n302 B.n57 585
R616 B.n304 B.n303 585
R617 B.n305 B.n56 585
R618 B.n307 B.n306 585
R619 B.n308 B.n55 585
R620 B.n310 B.n309 585
R621 B.n311 B.n54 585
R622 B.n313 B.n312 585
R623 B.n314 B.n53 585
R624 B.n316 B.n315 585
R625 B.n317 B.n52 585
R626 B.n319 B.n318 585
R627 B.n320 B.n51 585
R628 B.n322 B.n321 585
R629 B.n323 B.n50 585
R630 B.n325 B.n324 585
R631 B.n419 B.n14 585
R632 B.n418 B.n417 585
R633 B.n416 B.n15 585
R634 B.n415 B.n414 585
R635 B.n413 B.n16 585
R636 B.n412 B.n411 585
R637 B.n410 B.n17 585
R638 B.n409 B.n408 585
R639 B.n407 B.n18 585
R640 B.n406 B.n405 585
R641 B.n404 B.n19 585
R642 B.n403 B.n402 585
R643 B.n401 B.n20 585
R644 B.n400 B.n399 585
R645 B.n398 B.n21 585
R646 B.n397 B.n396 585
R647 B.n395 B.n22 585
R648 B.n394 B.n393 585
R649 B.n392 B.n23 585
R650 B.n391 B.n390 585
R651 B.n389 B.n24 585
R652 B.n388 B.n387 585
R653 B.n386 B.n25 585
R654 B.n385 B.n384 585
R655 B.n383 B.n26 585
R656 B.n382 B.n381 585
R657 B.n379 B.n27 585
R658 B.n378 B.n377 585
R659 B.n376 B.n30 585
R660 B.n375 B.n374 585
R661 B.n373 B.n31 585
R662 B.n372 B.n371 585
R663 B.n370 B.n32 585
R664 B.n369 B.n368 585
R665 B.n367 B.n33 585
R666 B.n366 B.n365 585
R667 B.n364 B.n363 585
R668 B.n362 B.n37 585
R669 B.n361 B.n360 585
R670 B.n359 B.n38 585
R671 B.n358 B.n357 585
R672 B.n356 B.n39 585
R673 B.n355 B.n354 585
R674 B.n353 B.n40 585
R675 B.n352 B.n351 585
R676 B.n350 B.n41 585
R677 B.n349 B.n348 585
R678 B.n347 B.n42 585
R679 B.n346 B.n345 585
R680 B.n344 B.n43 585
R681 B.n343 B.n342 585
R682 B.n341 B.n44 585
R683 B.n340 B.n339 585
R684 B.n338 B.n45 585
R685 B.n337 B.n336 585
R686 B.n335 B.n46 585
R687 B.n334 B.n333 585
R688 B.n332 B.n47 585
R689 B.n331 B.n330 585
R690 B.n329 B.n48 585
R691 B.n328 B.n327 585
R692 B.n326 B.n49 585
R693 B.n421 B.n420 585
R694 B.n422 B.n13 585
R695 B.n424 B.n423 585
R696 B.n425 B.n12 585
R697 B.n427 B.n426 585
R698 B.n428 B.n11 585
R699 B.n430 B.n429 585
R700 B.n431 B.n10 585
R701 B.n433 B.n432 585
R702 B.n434 B.n9 585
R703 B.n436 B.n435 585
R704 B.n437 B.n8 585
R705 B.n439 B.n438 585
R706 B.n440 B.n7 585
R707 B.n442 B.n441 585
R708 B.n443 B.n6 585
R709 B.n445 B.n444 585
R710 B.n446 B.n5 585
R711 B.n448 B.n447 585
R712 B.n449 B.n4 585
R713 B.n451 B.n450 585
R714 B.n452 B.n3 585
R715 B.n454 B.n453 585
R716 B.n455 B.n0 585
R717 B.n2 B.n1 585
R718 B.n120 B.n119 585
R719 B.n121 B.n118 585
R720 B.n123 B.n122 585
R721 B.n124 B.n117 585
R722 B.n126 B.n125 585
R723 B.n127 B.n116 585
R724 B.n129 B.n128 585
R725 B.n130 B.n115 585
R726 B.n132 B.n131 585
R727 B.n133 B.n114 585
R728 B.n135 B.n134 585
R729 B.n136 B.n113 585
R730 B.n138 B.n137 585
R731 B.n139 B.n112 585
R732 B.n141 B.n140 585
R733 B.n142 B.n111 585
R734 B.n144 B.n143 585
R735 B.n145 B.n110 585
R736 B.n147 B.n146 585
R737 B.n148 B.n109 585
R738 B.n150 B.n149 585
R739 B.n151 B.n108 585
R740 B.n153 B.n152 585
R741 B.n152 B.n107 521.33
R742 B.n251 B.n250 521.33
R743 B.n324 B.n49 521.33
R744 B.n420 B.n419 521.33
R745 B.n191 B.t9 356.089
R746 B.n88 B.t6 356.089
R747 B.n34 B.t0 356.089
R748 B.n28 B.t3 356.089
R749 B.n88 B.t7 309.277
R750 B.n34 B.t2 309.277
R751 B.n191 B.t10 309.277
R752 B.n28 B.t5 309.277
R753 B.n89 B.t8 282.125
R754 B.n35 B.t1 282.125
R755 B.n192 B.t11 282.125
R756 B.n29 B.t4 282.125
R757 B.n457 B.n456 256.663
R758 B.n456 B.n455 235.042
R759 B.n456 B.n2 235.042
R760 B.n156 B.n107 163.367
R761 B.n157 B.n156 163.367
R762 B.n158 B.n157 163.367
R763 B.n158 B.n105 163.367
R764 B.n162 B.n105 163.367
R765 B.n163 B.n162 163.367
R766 B.n164 B.n163 163.367
R767 B.n164 B.n103 163.367
R768 B.n168 B.n103 163.367
R769 B.n169 B.n168 163.367
R770 B.n170 B.n169 163.367
R771 B.n170 B.n101 163.367
R772 B.n174 B.n101 163.367
R773 B.n175 B.n174 163.367
R774 B.n176 B.n175 163.367
R775 B.n176 B.n99 163.367
R776 B.n180 B.n99 163.367
R777 B.n181 B.n180 163.367
R778 B.n182 B.n181 163.367
R779 B.n182 B.n97 163.367
R780 B.n186 B.n97 163.367
R781 B.n187 B.n186 163.367
R782 B.n188 B.n187 163.367
R783 B.n188 B.n95 163.367
R784 B.n195 B.n95 163.367
R785 B.n196 B.n195 163.367
R786 B.n197 B.n196 163.367
R787 B.n197 B.n93 163.367
R788 B.n201 B.n93 163.367
R789 B.n202 B.n201 163.367
R790 B.n203 B.n202 163.367
R791 B.n203 B.n91 163.367
R792 B.n207 B.n91 163.367
R793 B.n208 B.n207 163.367
R794 B.n209 B.n208 163.367
R795 B.n209 B.n87 163.367
R796 B.n214 B.n87 163.367
R797 B.n215 B.n214 163.367
R798 B.n216 B.n215 163.367
R799 B.n216 B.n85 163.367
R800 B.n220 B.n85 163.367
R801 B.n221 B.n220 163.367
R802 B.n222 B.n221 163.367
R803 B.n222 B.n83 163.367
R804 B.n226 B.n83 163.367
R805 B.n227 B.n226 163.367
R806 B.n228 B.n227 163.367
R807 B.n228 B.n81 163.367
R808 B.n232 B.n81 163.367
R809 B.n233 B.n232 163.367
R810 B.n234 B.n233 163.367
R811 B.n234 B.n79 163.367
R812 B.n238 B.n79 163.367
R813 B.n239 B.n238 163.367
R814 B.n240 B.n239 163.367
R815 B.n240 B.n77 163.367
R816 B.n244 B.n77 163.367
R817 B.n245 B.n244 163.367
R818 B.n246 B.n245 163.367
R819 B.n246 B.n75 163.367
R820 B.n250 B.n75 163.367
R821 B.n324 B.n323 163.367
R822 B.n323 B.n322 163.367
R823 B.n322 B.n51 163.367
R824 B.n318 B.n51 163.367
R825 B.n318 B.n317 163.367
R826 B.n317 B.n316 163.367
R827 B.n316 B.n53 163.367
R828 B.n312 B.n53 163.367
R829 B.n312 B.n311 163.367
R830 B.n311 B.n310 163.367
R831 B.n310 B.n55 163.367
R832 B.n306 B.n55 163.367
R833 B.n306 B.n305 163.367
R834 B.n305 B.n304 163.367
R835 B.n304 B.n57 163.367
R836 B.n300 B.n57 163.367
R837 B.n300 B.n299 163.367
R838 B.n299 B.n298 163.367
R839 B.n298 B.n59 163.367
R840 B.n294 B.n59 163.367
R841 B.n294 B.n293 163.367
R842 B.n293 B.n292 163.367
R843 B.n292 B.n61 163.367
R844 B.n288 B.n61 163.367
R845 B.n288 B.n287 163.367
R846 B.n287 B.n286 163.367
R847 B.n286 B.n63 163.367
R848 B.n282 B.n63 163.367
R849 B.n282 B.n281 163.367
R850 B.n281 B.n280 163.367
R851 B.n280 B.n65 163.367
R852 B.n276 B.n65 163.367
R853 B.n276 B.n275 163.367
R854 B.n275 B.n274 163.367
R855 B.n274 B.n67 163.367
R856 B.n270 B.n67 163.367
R857 B.n270 B.n269 163.367
R858 B.n269 B.n268 163.367
R859 B.n268 B.n69 163.367
R860 B.n264 B.n69 163.367
R861 B.n264 B.n263 163.367
R862 B.n263 B.n262 163.367
R863 B.n262 B.n71 163.367
R864 B.n258 B.n71 163.367
R865 B.n258 B.n257 163.367
R866 B.n257 B.n256 163.367
R867 B.n256 B.n73 163.367
R868 B.n252 B.n73 163.367
R869 B.n252 B.n251 163.367
R870 B.n419 B.n418 163.367
R871 B.n418 B.n15 163.367
R872 B.n414 B.n15 163.367
R873 B.n414 B.n413 163.367
R874 B.n413 B.n412 163.367
R875 B.n412 B.n17 163.367
R876 B.n408 B.n17 163.367
R877 B.n408 B.n407 163.367
R878 B.n407 B.n406 163.367
R879 B.n406 B.n19 163.367
R880 B.n402 B.n19 163.367
R881 B.n402 B.n401 163.367
R882 B.n401 B.n400 163.367
R883 B.n400 B.n21 163.367
R884 B.n396 B.n21 163.367
R885 B.n396 B.n395 163.367
R886 B.n395 B.n394 163.367
R887 B.n394 B.n23 163.367
R888 B.n390 B.n23 163.367
R889 B.n390 B.n389 163.367
R890 B.n389 B.n388 163.367
R891 B.n388 B.n25 163.367
R892 B.n384 B.n25 163.367
R893 B.n384 B.n383 163.367
R894 B.n383 B.n382 163.367
R895 B.n382 B.n27 163.367
R896 B.n377 B.n27 163.367
R897 B.n377 B.n376 163.367
R898 B.n376 B.n375 163.367
R899 B.n375 B.n31 163.367
R900 B.n371 B.n31 163.367
R901 B.n371 B.n370 163.367
R902 B.n370 B.n369 163.367
R903 B.n369 B.n33 163.367
R904 B.n365 B.n33 163.367
R905 B.n365 B.n364 163.367
R906 B.n364 B.n37 163.367
R907 B.n360 B.n37 163.367
R908 B.n360 B.n359 163.367
R909 B.n359 B.n358 163.367
R910 B.n358 B.n39 163.367
R911 B.n354 B.n39 163.367
R912 B.n354 B.n353 163.367
R913 B.n353 B.n352 163.367
R914 B.n352 B.n41 163.367
R915 B.n348 B.n41 163.367
R916 B.n348 B.n347 163.367
R917 B.n347 B.n346 163.367
R918 B.n346 B.n43 163.367
R919 B.n342 B.n43 163.367
R920 B.n342 B.n341 163.367
R921 B.n341 B.n340 163.367
R922 B.n340 B.n45 163.367
R923 B.n336 B.n45 163.367
R924 B.n336 B.n335 163.367
R925 B.n335 B.n334 163.367
R926 B.n334 B.n47 163.367
R927 B.n330 B.n47 163.367
R928 B.n330 B.n329 163.367
R929 B.n329 B.n328 163.367
R930 B.n328 B.n49 163.367
R931 B.n420 B.n13 163.367
R932 B.n424 B.n13 163.367
R933 B.n425 B.n424 163.367
R934 B.n426 B.n425 163.367
R935 B.n426 B.n11 163.367
R936 B.n430 B.n11 163.367
R937 B.n431 B.n430 163.367
R938 B.n432 B.n431 163.367
R939 B.n432 B.n9 163.367
R940 B.n436 B.n9 163.367
R941 B.n437 B.n436 163.367
R942 B.n438 B.n437 163.367
R943 B.n438 B.n7 163.367
R944 B.n442 B.n7 163.367
R945 B.n443 B.n442 163.367
R946 B.n444 B.n443 163.367
R947 B.n444 B.n5 163.367
R948 B.n448 B.n5 163.367
R949 B.n449 B.n448 163.367
R950 B.n450 B.n449 163.367
R951 B.n450 B.n3 163.367
R952 B.n454 B.n3 163.367
R953 B.n455 B.n454 163.367
R954 B.n120 B.n2 163.367
R955 B.n121 B.n120 163.367
R956 B.n122 B.n121 163.367
R957 B.n122 B.n117 163.367
R958 B.n126 B.n117 163.367
R959 B.n127 B.n126 163.367
R960 B.n128 B.n127 163.367
R961 B.n128 B.n115 163.367
R962 B.n132 B.n115 163.367
R963 B.n133 B.n132 163.367
R964 B.n134 B.n133 163.367
R965 B.n134 B.n113 163.367
R966 B.n138 B.n113 163.367
R967 B.n139 B.n138 163.367
R968 B.n140 B.n139 163.367
R969 B.n140 B.n111 163.367
R970 B.n144 B.n111 163.367
R971 B.n145 B.n144 163.367
R972 B.n146 B.n145 163.367
R973 B.n146 B.n109 163.367
R974 B.n150 B.n109 163.367
R975 B.n151 B.n150 163.367
R976 B.n152 B.n151 163.367
R977 B.n193 B.n192 59.5399
R978 B.n211 B.n89 59.5399
R979 B.n36 B.n35 59.5399
R980 B.n380 B.n29 59.5399
R981 B.n421 B.n14 33.8737
R982 B.n326 B.n325 33.8737
R983 B.n249 B.n74 33.8737
R984 B.n154 B.n153 33.8737
R985 B.n192 B.n191 27.152
R986 B.n89 B.n88 27.152
R987 B.n35 B.n34 27.152
R988 B.n29 B.n28 27.152
R989 B B.n457 18.0485
R990 B.n422 B.n421 10.6151
R991 B.n423 B.n422 10.6151
R992 B.n423 B.n12 10.6151
R993 B.n427 B.n12 10.6151
R994 B.n428 B.n427 10.6151
R995 B.n429 B.n428 10.6151
R996 B.n429 B.n10 10.6151
R997 B.n433 B.n10 10.6151
R998 B.n434 B.n433 10.6151
R999 B.n435 B.n434 10.6151
R1000 B.n435 B.n8 10.6151
R1001 B.n439 B.n8 10.6151
R1002 B.n440 B.n439 10.6151
R1003 B.n441 B.n440 10.6151
R1004 B.n441 B.n6 10.6151
R1005 B.n445 B.n6 10.6151
R1006 B.n446 B.n445 10.6151
R1007 B.n447 B.n446 10.6151
R1008 B.n447 B.n4 10.6151
R1009 B.n451 B.n4 10.6151
R1010 B.n452 B.n451 10.6151
R1011 B.n453 B.n452 10.6151
R1012 B.n453 B.n0 10.6151
R1013 B.n417 B.n14 10.6151
R1014 B.n417 B.n416 10.6151
R1015 B.n416 B.n415 10.6151
R1016 B.n415 B.n16 10.6151
R1017 B.n411 B.n16 10.6151
R1018 B.n411 B.n410 10.6151
R1019 B.n410 B.n409 10.6151
R1020 B.n409 B.n18 10.6151
R1021 B.n405 B.n18 10.6151
R1022 B.n405 B.n404 10.6151
R1023 B.n404 B.n403 10.6151
R1024 B.n403 B.n20 10.6151
R1025 B.n399 B.n20 10.6151
R1026 B.n399 B.n398 10.6151
R1027 B.n398 B.n397 10.6151
R1028 B.n397 B.n22 10.6151
R1029 B.n393 B.n22 10.6151
R1030 B.n393 B.n392 10.6151
R1031 B.n392 B.n391 10.6151
R1032 B.n391 B.n24 10.6151
R1033 B.n387 B.n24 10.6151
R1034 B.n387 B.n386 10.6151
R1035 B.n386 B.n385 10.6151
R1036 B.n385 B.n26 10.6151
R1037 B.n381 B.n26 10.6151
R1038 B.n379 B.n378 10.6151
R1039 B.n378 B.n30 10.6151
R1040 B.n374 B.n30 10.6151
R1041 B.n374 B.n373 10.6151
R1042 B.n373 B.n372 10.6151
R1043 B.n372 B.n32 10.6151
R1044 B.n368 B.n32 10.6151
R1045 B.n368 B.n367 10.6151
R1046 B.n367 B.n366 10.6151
R1047 B.n363 B.n362 10.6151
R1048 B.n362 B.n361 10.6151
R1049 B.n361 B.n38 10.6151
R1050 B.n357 B.n38 10.6151
R1051 B.n357 B.n356 10.6151
R1052 B.n356 B.n355 10.6151
R1053 B.n355 B.n40 10.6151
R1054 B.n351 B.n40 10.6151
R1055 B.n351 B.n350 10.6151
R1056 B.n350 B.n349 10.6151
R1057 B.n349 B.n42 10.6151
R1058 B.n345 B.n42 10.6151
R1059 B.n345 B.n344 10.6151
R1060 B.n344 B.n343 10.6151
R1061 B.n343 B.n44 10.6151
R1062 B.n339 B.n44 10.6151
R1063 B.n339 B.n338 10.6151
R1064 B.n338 B.n337 10.6151
R1065 B.n337 B.n46 10.6151
R1066 B.n333 B.n46 10.6151
R1067 B.n333 B.n332 10.6151
R1068 B.n332 B.n331 10.6151
R1069 B.n331 B.n48 10.6151
R1070 B.n327 B.n48 10.6151
R1071 B.n327 B.n326 10.6151
R1072 B.n325 B.n50 10.6151
R1073 B.n321 B.n50 10.6151
R1074 B.n321 B.n320 10.6151
R1075 B.n320 B.n319 10.6151
R1076 B.n319 B.n52 10.6151
R1077 B.n315 B.n52 10.6151
R1078 B.n315 B.n314 10.6151
R1079 B.n314 B.n313 10.6151
R1080 B.n313 B.n54 10.6151
R1081 B.n309 B.n54 10.6151
R1082 B.n309 B.n308 10.6151
R1083 B.n308 B.n307 10.6151
R1084 B.n307 B.n56 10.6151
R1085 B.n303 B.n56 10.6151
R1086 B.n303 B.n302 10.6151
R1087 B.n302 B.n301 10.6151
R1088 B.n301 B.n58 10.6151
R1089 B.n297 B.n58 10.6151
R1090 B.n297 B.n296 10.6151
R1091 B.n296 B.n295 10.6151
R1092 B.n295 B.n60 10.6151
R1093 B.n291 B.n60 10.6151
R1094 B.n291 B.n290 10.6151
R1095 B.n290 B.n289 10.6151
R1096 B.n289 B.n62 10.6151
R1097 B.n285 B.n62 10.6151
R1098 B.n285 B.n284 10.6151
R1099 B.n284 B.n283 10.6151
R1100 B.n283 B.n64 10.6151
R1101 B.n279 B.n64 10.6151
R1102 B.n279 B.n278 10.6151
R1103 B.n278 B.n277 10.6151
R1104 B.n277 B.n66 10.6151
R1105 B.n273 B.n66 10.6151
R1106 B.n273 B.n272 10.6151
R1107 B.n272 B.n271 10.6151
R1108 B.n271 B.n68 10.6151
R1109 B.n267 B.n68 10.6151
R1110 B.n267 B.n266 10.6151
R1111 B.n266 B.n265 10.6151
R1112 B.n265 B.n70 10.6151
R1113 B.n261 B.n70 10.6151
R1114 B.n261 B.n260 10.6151
R1115 B.n260 B.n259 10.6151
R1116 B.n259 B.n72 10.6151
R1117 B.n255 B.n72 10.6151
R1118 B.n255 B.n254 10.6151
R1119 B.n254 B.n253 10.6151
R1120 B.n253 B.n74 10.6151
R1121 B.n119 B.n1 10.6151
R1122 B.n119 B.n118 10.6151
R1123 B.n123 B.n118 10.6151
R1124 B.n124 B.n123 10.6151
R1125 B.n125 B.n124 10.6151
R1126 B.n125 B.n116 10.6151
R1127 B.n129 B.n116 10.6151
R1128 B.n130 B.n129 10.6151
R1129 B.n131 B.n130 10.6151
R1130 B.n131 B.n114 10.6151
R1131 B.n135 B.n114 10.6151
R1132 B.n136 B.n135 10.6151
R1133 B.n137 B.n136 10.6151
R1134 B.n137 B.n112 10.6151
R1135 B.n141 B.n112 10.6151
R1136 B.n142 B.n141 10.6151
R1137 B.n143 B.n142 10.6151
R1138 B.n143 B.n110 10.6151
R1139 B.n147 B.n110 10.6151
R1140 B.n148 B.n147 10.6151
R1141 B.n149 B.n148 10.6151
R1142 B.n149 B.n108 10.6151
R1143 B.n153 B.n108 10.6151
R1144 B.n155 B.n154 10.6151
R1145 B.n155 B.n106 10.6151
R1146 B.n159 B.n106 10.6151
R1147 B.n160 B.n159 10.6151
R1148 B.n161 B.n160 10.6151
R1149 B.n161 B.n104 10.6151
R1150 B.n165 B.n104 10.6151
R1151 B.n166 B.n165 10.6151
R1152 B.n167 B.n166 10.6151
R1153 B.n167 B.n102 10.6151
R1154 B.n171 B.n102 10.6151
R1155 B.n172 B.n171 10.6151
R1156 B.n173 B.n172 10.6151
R1157 B.n173 B.n100 10.6151
R1158 B.n177 B.n100 10.6151
R1159 B.n178 B.n177 10.6151
R1160 B.n179 B.n178 10.6151
R1161 B.n179 B.n98 10.6151
R1162 B.n183 B.n98 10.6151
R1163 B.n184 B.n183 10.6151
R1164 B.n185 B.n184 10.6151
R1165 B.n185 B.n96 10.6151
R1166 B.n189 B.n96 10.6151
R1167 B.n190 B.n189 10.6151
R1168 B.n194 B.n190 10.6151
R1169 B.n198 B.n94 10.6151
R1170 B.n199 B.n198 10.6151
R1171 B.n200 B.n199 10.6151
R1172 B.n200 B.n92 10.6151
R1173 B.n204 B.n92 10.6151
R1174 B.n205 B.n204 10.6151
R1175 B.n206 B.n205 10.6151
R1176 B.n206 B.n90 10.6151
R1177 B.n210 B.n90 10.6151
R1178 B.n213 B.n212 10.6151
R1179 B.n213 B.n86 10.6151
R1180 B.n217 B.n86 10.6151
R1181 B.n218 B.n217 10.6151
R1182 B.n219 B.n218 10.6151
R1183 B.n219 B.n84 10.6151
R1184 B.n223 B.n84 10.6151
R1185 B.n224 B.n223 10.6151
R1186 B.n225 B.n224 10.6151
R1187 B.n225 B.n82 10.6151
R1188 B.n229 B.n82 10.6151
R1189 B.n230 B.n229 10.6151
R1190 B.n231 B.n230 10.6151
R1191 B.n231 B.n80 10.6151
R1192 B.n235 B.n80 10.6151
R1193 B.n236 B.n235 10.6151
R1194 B.n237 B.n236 10.6151
R1195 B.n237 B.n78 10.6151
R1196 B.n241 B.n78 10.6151
R1197 B.n242 B.n241 10.6151
R1198 B.n243 B.n242 10.6151
R1199 B.n243 B.n76 10.6151
R1200 B.n247 B.n76 10.6151
R1201 B.n248 B.n247 10.6151
R1202 B.n249 B.n248 10.6151
R1203 B.n381 B.n380 9.36635
R1204 B.n363 B.n36 9.36635
R1205 B.n194 B.n193 9.36635
R1206 B.n212 B.n211 9.36635
R1207 B.n457 B.n0 8.11757
R1208 B.n457 B.n1 8.11757
R1209 B.n380 B.n379 1.24928
R1210 B.n366 B.n36 1.24928
R1211 B.n193 B.n94 1.24928
R1212 B.n211 B.n210 1.24928
C0 VTAIL B 1.94704f
C1 VN w_n2090_n2324# 3.48521f
C2 VDD1 VP 3.27859f
C3 VDD2 w_n2090_n2324# 1.56804f
C4 VDD1 B 1.28185f
C5 VN VP 4.47013f
C6 VDD1 VTAIL 5.81775f
C7 VDD2 VP 0.328552f
C8 VN B 0.78362f
C9 VDD2 B 1.31952f
C10 VN VTAIL 3.17446f
C11 VDD2 VTAIL 5.85794f
C12 VP w_n2090_n2324# 3.75116f
C13 w_n2090_n2324# B 6.10215f
C14 VN VDD1 0.149042f
C15 VDD2 VDD1 0.845561f
C16 VTAIL w_n2090_n2324# 2.12516f
C17 VP B 1.21994f
C18 VN VDD2 3.10161f
C19 VTAIL VP 3.1888f
C20 VDD1 w_n2090_n2324# 1.53222f
C21 VDD2 VSUBS 1.15537f
C22 VDD1 VSUBS 1.079434f
C23 VTAIL VSUBS 0.522334f
C24 VN VSUBS 4.26057f
C25 VP VSUBS 1.503638f
C26 B VSUBS 2.68318f
C27 w_n2090_n2324# VSUBS 60.4679f
C28 B.n0 VSUBS 0.005395f
C29 B.n1 VSUBS 0.005395f
C30 B.n2 VSUBS 0.007979f
C31 B.n3 VSUBS 0.006114f
C32 B.n4 VSUBS 0.006114f
C33 B.n5 VSUBS 0.006114f
C34 B.n6 VSUBS 0.006114f
C35 B.n7 VSUBS 0.006114f
C36 B.n8 VSUBS 0.006114f
C37 B.n9 VSUBS 0.006114f
C38 B.n10 VSUBS 0.006114f
C39 B.n11 VSUBS 0.006114f
C40 B.n12 VSUBS 0.006114f
C41 B.n13 VSUBS 0.006114f
C42 B.n14 VSUBS 0.015004f
C43 B.n15 VSUBS 0.006114f
C44 B.n16 VSUBS 0.006114f
C45 B.n17 VSUBS 0.006114f
C46 B.n18 VSUBS 0.006114f
C47 B.n19 VSUBS 0.006114f
C48 B.n20 VSUBS 0.006114f
C49 B.n21 VSUBS 0.006114f
C50 B.n22 VSUBS 0.006114f
C51 B.n23 VSUBS 0.006114f
C52 B.n24 VSUBS 0.006114f
C53 B.n25 VSUBS 0.006114f
C54 B.n26 VSUBS 0.006114f
C55 B.n27 VSUBS 0.006114f
C56 B.t4 VSUBS 0.090553f
C57 B.t5 VSUBS 0.102372f
C58 B.t3 VSUBS 0.281001f
C59 B.n28 VSUBS 0.174913f
C60 B.n29 VSUBS 0.143352f
C61 B.n30 VSUBS 0.006114f
C62 B.n31 VSUBS 0.006114f
C63 B.n32 VSUBS 0.006114f
C64 B.n33 VSUBS 0.006114f
C65 B.t1 VSUBS 0.090555f
C66 B.t2 VSUBS 0.102374f
C67 B.t0 VSUBS 0.281001f
C68 B.n34 VSUBS 0.174911f
C69 B.n35 VSUBS 0.14335f
C70 B.n36 VSUBS 0.014166f
C71 B.n37 VSUBS 0.006114f
C72 B.n38 VSUBS 0.006114f
C73 B.n39 VSUBS 0.006114f
C74 B.n40 VSUBS 0.006114f
C75 B.n41 VSUBS 0.006114f
C76 B.n42 VSUBS 0.006114f
C77 B.n43 VSUBS 0.006114f
C78 B.n44 VSUBS 0.006114f
C79 B.n45 VSUBS 0.006114f
C80 B.n46 VSUBS 0.006114f
C81 B.n47 VSUBS 0.006114f
C82 B.n48 VSUBS 0.006114f
C83 B.n49 VSUBS 0.015004f
C84 B.n50 VSUBS 0.006114f
C85 B.n51 VSUBS 0.006114f
C86 B.n52 VSUBS 0.006114f
C87 B.n53 VSUBS 0.006114f
C88 B.n54 VSUBS 0.006114f
C89 B.n55 VSUBS 0.006114f
C90 B.n56 VSUBS 0.006114f
C91 B.n57 VSUBS 0.006114f
C92 B.n58 VSUBS 0.006114f
C93 B.n59 VSUBS 0.006114f
C94 B.n60 VSUBS 0.006114f
C95 B.n61 VSUBS 0.006114f
C96 B.n62 VSUBS 0.006114f
C97 B.n63 VSUBS 0.006114f
C98 B.n64 VSUBS 0.006114f
C99 B.n65 VSUBS 0.006114f
C100 B.n66 VSUBS 0.006114f
C101 B.n67 VSUBS 0.006114f
C102 B.n68 VSUBS 0.006114f
C103 B.n69 VSUBS 0.006114f
C104 B.n70 VSUBS 0.006114f
C105 B.n71 VSUBS 0.006114f
C106 B.n72 VSUBS 0.006114f
C107 B.n73 VSUBS 0.006114f
C108 B.n74 VSUBS 0.015004f
C109 B.n75 VSUBS 0.006114f
C110 B.n76 VSUBS 0.006114f
C111 B.n77 VSUBS 0.006114f
C112 B.n78 VSUBS 0.006114f
C113 B.n79 VSUBS 0.006114f
C114 B.n80 VSUBS 0.006114f
C115 B.n81 VSUBS 0.006114f
C116 B.n82 VSUBS 0.006114f
C117 B.n83 VSUBS 0.006114f
C118 B.n84 VSUBS 0.006114f
C119 B.n85 VSUBS 0.006114f
C120 B.n86 VSUBS 0.006114f
C121 B.n87 VSUBS 0.006114f
C122 B.t8 VSUBS 0.090555f
C123 B.t7 VSUBS 0.102374f
C124 B.t6 VSUBS 0.281001f
C125 B.n88 VSUBS 0.174911f
C126 B.n89 VSUBS 0.14335f
C127 B.n90 VSUBS 0.006114f
C128 B.n91 VSUBS 0.006114f
C129 B.n92 VSUBS 0.006114f
C130 B.n93 VSUBS 0.006114f
C131 B.n94 VSUBS 0.003417f
C132 B.n95 VSUBS 0.006114f
C133 B.n96 VSUBS 0.006114f
C134 B.n97 VSUBS 0.006114f
C135 B.n98 VSUBS 0.006114f
C136 B.n99 VSUBS 0.006114f
C137 B.n100 VSUBS 0.006114f
C138 B.n101 VSUBS 0.006114f
C139 B.n102 VSUBS 0.006114f
C140 B.n103 VSUBS 0.006114f
C141 B.n104 VSUBS 0.006114f
C142 B.n105 VSUBS 0.006114f
C143 B.n106 VSUBS 0.006114f
C144 B.n107 VSUBS 0.015004f
C145 B.n108 VSUBS 0.006114f
C146 B.n109 VSUBS 0.006114f
C147 B.n110 VSUBS 0.006114f
C148 B.n111 VSUBS 0.006114f
C149 B.n112 VSUBS 0.006114f
C150 B.n113 VSUBS 0.006114f
C151 B.n114 VSUBS 0.006114f
C152 B.n115 VSUBS 0.006114f
C153 B.n116 VSUBS 0.006114f
C154 B.n117 VSUBS 0.006114f
C155 B.n118 VSUBS 0.006114f
C156 B.n119 VSUBS 0.006114f
C157 B.n120 VSUBS 0.006114f
C158 B.n121 VSUBS 0.006114f
C159 B.n122 VSUBS 0.006114f
C160 B.n123 VSUBS 0.006114f
C161 B.n124 VSUBS 0.006114f
C162 B.n125 VSUBS 0.006114f
C163 B.n126 VSUBS 0.006114f
C164 B.n127 VSUBS 0.006114f
C165 B.n128 VSUBS 0.006114f
C166 B.n129 VSUBS 0.006114f
C167 B.n130 VSUBS 0.006114f
C168 B.n131 VSUBS 0.006114f
C169 B.n132 VSUBS 0.006114f
C170 B.n133 VSUBS 0.006114f
C171 B.n134 VSUBS 0.006114f
C172 B.n135 VSUBS 0.006114f
C173 B.n136 VSUBS 0.006114f
C174 B.n137 VSUBS 0.006114f
C175 B.n138 VSUBS 0.006114f
C176 B.n139 VSUBS 0.006114f
C177 B.n140 VSUBS 0.006114f
C178 B.n141 VSUBS 0.006114f
C179 B.n142 VSUBS 0.006114f
C180 B.n143 VSUBS 0.006114f
C181 B.n144 VSUBS 0.006114f
C182 B.n145 VSUBS 0.006114f
C183 B.n146 VSUBS 0.006114f
C184 B.n147 VSUBS 0.006114f
C185 B.n148 VSUBS 0.006114f
C186 B.n149 VSUBS 0.006114f
C187 B.n150 VSUBS 0.006114f
C188 B.n151 VSUBS 0.006114f
C189 B.n152 VSUBS 0.014308f
C190 B.n153 VSUBS 0.014308f
C191 B.n154 VSUBS 0.015004f
C192 B.n155 VSUBS 0.006114f
C193 B.n156 VSUBS 0.006114f
C194 B.n157 VSUBS 0.006114f
C195 B.n158 VSUBS 0.006114f
C196 B.n159 VSUBS 0.006114f
C197 B.n160 VSUBS 0.006114f
C198 B.n161 VSUBS 0.006114f
C199 B.n162 VSUBS 0.006114f
C200 B.n163 VSUBS 0.006114f
C201 B.n164 VSUBS 0.006114f
C202 B.n165 VSUBS 0.006114f
C203 B.n166 VSUBS 0.006114f
C204 B.n167 VSUBS 0.006114f
C205 B.n168 VSUBS 0.006114f
C206 B.n169 VSUBS 0.006114f
C207 B.n170 VSUBS 0.006114f
C208 B.n171 VSUBS 0.006114f
C209 B.n172 VSUBS 0.006114f
C210 B.n173 VSUBS 0.006114f
C211 B.n174 VSUBS 0.006114f
C212 B.n175 VSUBS 0.006114f
C213 B.n176 VSUBS 0.006114f
C214 B.n177 VSUBS 0.006114f
C215 B.n178 VSUBS 0.006114f
C216 B.n179 VSUBS 0.006114f
C217 B.n180 VSUBS 0.006114f
C218 B.n181 VSUBS 0.006114f
C219 B.n182 VSUBS 0.006114f
C220 B.n183 VSUBS 0.006114f
C221 B.n184 VSUBS 0.006114f
C222 B.n185 VSUBS 0.006114f
C223 B.n186 VSUBS 0.006114f
C224 B.n187 VSUBS 0.006114f
C225 B.n188 VSUBS 0.006114f
C226 B.n189 VSUBS 0.006114f
C227 B.n190 VSUBS 0.006114f
C228 B.t11 VSUBS 0.090553f
C229 B.t10 VSUBS 0.102372f
C230 B.t9 VSUBS 0.281001f
C231 B.n191 VSUBS 0.174913f
C232 B.n192 VSUBS 0.143352f
C233 B.n193 VSUBS 0.014166f
C234 B.n194 VSUBS 0.005755f
C235 B.n195 VSUBS 0.006114f
C236 B.n196 VSUBS 0.006114f
C237 B.n197 VSUBS 0.006114f
C238 B.n198 VSUBS 0.006114f
C239 B.n199 VSUBS 0.006114f
C240 B.n200 VSUBS 0.006114f
C241 B.n201 VSUBS 0.006114f
C242 B.n202 VSUBS 0.006114f
C243 B.n203 VSUBS 0.006114f
C244 B.n204 VSUBS 0.006114f
C245 B.n205 VSUBS 0.006114f
C246 B.n206 VSUBS 0.006114f
C247 B.n207 VSUBS 0.006114f
C248 B.n208 VSUBS 0.006114f
C249 B.n209 VSUBS 0.006114f
C250 B.n210 VSUBS 0.003417f
C251 B.n211 VSUBS 0.014166f
C252 B.n212 VSUBS 0.005755f
C253 B.n213 VSUBS 0.006114f
C254 B.n214 VSUBS 0.006114f
C255 B.n215 VSUBS 0.006114f
C256 B.n216 VSUBS 0.006114f
C257 B.n217 VSUBS 0.006114f
C258 B.n218 VSUBS 0.006114f
C259 B.n219 VSUBS 0.006114f
C260 B.n220 VSUBS 0.006114f
C261 B.n221 VSUBS 0.006114f
C262 B.n222 VSUBS 0.006114f
C263 B.n223 VSUBS 0.006114f
C264 B.n224 VSUBS 0.006114f
C265 B.n225 VSUBS 0.006114f
C266 B.n226 VSUBS 0.006114f
C267 B.n227 VSUBS 0.006114f
C268 B.n228 VSUBS 0.006114f
C269 B.n229 VSUBS 0.006114f
C270 B.n230 VSUBS 0.006114f
C271 B.n231 VSUBS 0.006114f
C272 B.n232 VSUBS 0.006114f
C273 B.n233 VSUBS 0.006114f
C274 B.n234 VSUBS 0.006114f
C275 B.n235 VSUBS 0.006114f
C276 B.n236 VSUBS 0.006114f
C277 B.n237 VSUBS 0.006114f
C278 B.n238 VSUBS 0.006114f
C279 B.n239 VSUBS 0.006114f
C280 B.n240 VSUBS 0.006114f
C281 B.n241 VSUBS 0.006114f
C282 B.n242 VSUBS 0.006114f
C283 B.n243 VSUBS 0.006114f
C284 B.n244 VSUBS 0.006114f
C285 B.n245 VSUBS 0.006114f
C286 B.n246 VSUBS 0.006114f
C287 B.n247 VSUBS 0.006114f
C288 B.n248 VSUBS 0.006114f
C289 B.n249 VSUBS 0.014308f
C290 B.n250 VSUBS 0.015004f
C291 B.n251 VSUBS 0.014308f
C292 B.n252 VSUBS 0.006114f
C293 B.n253 VSUBS 0.006114f
C294 B.n254 VSUBS 0.006114f
C295 B.n255 VSUBS 0.006114f
C296 B.n256 VSUBS 0.006114f
C297 B.n257 VSUBS 0.006114f
C298 B.n258 VSUBS 0.006114f
C299 B.n259 VSUBS 0.006114f
C300 B.n260 VSUBS 0.006114f
C301 B.n261 VSUBS 0.006114f
C302 B.n262 VSUBS 0.006114f
C303 B.n263 VSUBS 0.006114f
C304 B.n264 VSUBS 0.006114f
C305 B.n265 VSUBS 0.006114f
C306 B.n266 VSUBS 0.006114f
C307 B.n267 VSUBS 0.006114f
C308 B.n268 VSUBS 0.006114f
C309 B.n269 VSUBS 0.006114f
C310 B.n270 VSUBS 0.006114f
C311 B.n271 VSUBS 0.006114f
C312 B.n272 VSUBS 0.006114f
C313 B.n273 VSUBS 0.006114f
C314 B.n274 VSUBS 0.006114f
C315 B.n275 VSUBS 0.006114f
C316 B.n276 VSUBS 0.006114f
C317 B.n277 VSUBS 0.006114f
C318 B.n278 VSUBS 0.006114f
C319 B.n279 VSUBS 0.006114f
C320 B.n280 VSUBS 0.006114f
C321 B.n281 VSUBS 0.006114f
C322 B.n282 VSUBS 0.006114f
C323 B.n283 VSUBS 0.006114f
C324 B.n284 VSUBS 0.006114f
C325 B.n285 VSUBS 0.006114f
C326 B.n286 VSUBS 0.006114f
C327 B.n287 VSUBS 0.006114f
C328 B.n288 VSUBS 0.006114f
C329 B.n289 VSUBS 0.006114f
C330 B.n290 VSUBS 0.006114f
C331 B.n291 VSUBS 0.006114f
C332 B.n292 VSUBS 0.006114f
C333 B.n293 VSUBS 0.006114f
C334 B.n294 VSUBS 0.006114f
C335 B.n295 VSUBS 0.006114f
C336 B.n296 VSUBS 0.006114f
C337 B.n297 VSUBS 0.006114f
C338 B.n298 VSUBS 0.006114f
C339 B.n299 VSUBS 0.006114f
C340 B.n300 VSUBS 0.006114f
C341 B.n301 VSUBS 0.006114f
C342 B.n302 VSUBS 0.006114f
C343 B.n303 VSUBS 0.006114f
C344 B.n304 VSUBS 0.006114f
C345 B.n305 VSUBS 0.006114f
C346 B.n306 VSUBS 0.006114f
C347 B.n307 VSUBS 0.006114f
C348 B.n308 VSUBS 0.006114f
C349 B.n309 VSUBS 0.006114f
C350 B.n310 VSUBS 0.006114f
C351 B.n311 VSUBS 0.006114f
C352 B.n312 VSUBS 0.006114f
C353 B.n313 VSUBS 0.006114f
C354 B.n314 VSUBS 0.006114f
C355 B.n315 VSUBS 0.006114f
C356 B.n316 VSUBS 0.006114f
C357 B.n317 VSUBS 0.006114f
C358 B.n318 VSUBS 0.006114f
C359 B.n319 VSUBS 0.006114f
C360 B.n320 VSUBS 0.006114f
C361 B.n321 VSUBS 0.006114f
C362 B.n322 VSUBS 0.006114f
C363 B.n323 VSUBS 0.006114f
C364 B.n324 VSUBS 0.014308f
C365 B.n325 VSUBS 0.014308f
C366 B.n326 VSUBS 0.015004f
C367 B.n327 VSUBS 0.006114f
C368 B.n328 VSUBS 0.006114f
C369 B.n329 VSUBS 0.006114f
C370 B.n330 VSUBS 0.006114f
C371 B.n331 VSUBS 0.006114f
C372 B.n332 VSUBS 0.006114f
C373 B.n333 VSUBS 0.006114f
C374 B.n334 VSUBS 0.006114f
C375 B.n335 VSUBS 0.006114f
C376 B.n336 VSUBS 0.006114f
C377 B.n337 VSUBS 0.006114f
C378 B.n338 VSUBS 0.006114f
C379 B.n339 VSUBS 0.006114f
C380 B.n340 VSUBS 0.006114f
C381 B.n341 VSUBS 0.006114f
C382 B.n342 VSUBS 0.006114f
C383 B.n343 VSUBS 0.006114f
C384 B.n344 VSUBS 0.006114f
C385 B.n345 VSUBS 0.006114f
C386 B.n346 VSUBS 0.006114f
C387 B.n347 VSUBS 0.006114f
C388 B.n348 VSUBS 0.006114f
C389 B.n349 VSUBS 0.006114f
C390 B.n350 VSUBS 0.006114f
C391 B.n351 VSUBS 0.006114f
C392 B.n352 VSUBS 0.006114f
C393 B.n353 VSUBS 0.006114f
C394 B.n354 VSUBS 0.006114f
C395 B.n355 VSUBS 0.006114f
C396 B.n356 VSUBS 0.006114f
C397 B.n357 VSUBS 0.006114f
C398 B.n358 VSUBS 0.006114f
C399 B.n359 VSUBS 0.006114f
C400 B.n360 VSUBS 0.006114f
C401 B.n361 VSUBS 0.006114f
C402 B.n362 VSUBS 0.006114f
C403 B.n363 VSUBS 0.005755f
C404 B.n364 VSUBS 0.006114f
C405 B.n365 VSUBS 0.006114f
C406 B.n366 VSUBS 0.003417f
C407 B.n367 VSUBS 0.006114f
C408 B.n368 VSUBS 0.006114f
C409 B.n369 VSUBS 0.006114f
C410 B.n370 VSUBS 0.006114f
C411 B.n371 VSUBS 0.006114f
C412 B.n372 VSUBS 0.006114f
C413 B.n373 VSUBS 0.006114f
C414 B.n374 VSUBS 0.006114f
C415 B.n375 VSUBS 0.006114f
C416 B.n376 VSUBS 0.006114f
C417 B.n377 VSUBS 0.006114f
C418 B.n378 VSUBS 0.006114f
C419 B.n379 VSUBS 0.003417f
C420 B.n380 VSUBS 0.014166f
C421 B.n381 VSUBS 0.005755f
C422 B.n382 VSUBS 0.006114f
C423 B.n383 VSUBS 0.006114f
C424 B.n384 VSUBS 0.006114f
C425 B.n385 VSUBS 0.006114f
C426 B.n386 VSUBS 0.006114f
C427 B.n387 VSUBS 0.006114f
C428 B.n388 VSUBS 0.006114f
C429 B.n389 VSUBS 0.006114f
C430 B.n390 VSUBS 0.006114f
C431 B.n391 VSUBS 0.006114f
C432 B.n392 VSUBS 0.006114f
C433 B.n393 VSUBS 0.006114f
C434 B.n394 VSUBS 0.006114f
C435 B.n395 VSUBS 0.006114f
C436 B.n396 VSUBS 0.006114f
C437 B.n397 VSUBS 0.006114f
C438 B.n398 VSUBS 0.006114f
C439 B.n399 VSUBS 0.006114f
C440 B.n400 VSUBS 0.006114f
C441 B.n401 VSUBS 0.006114f
C442 B.n402 VSUBS 0.006114f
C443 B.n403 VSUBS 0.006114f
C444 B.n404 VSUBS 0.006114f
C445 B.n405 VSUBS 0.006114f
C446 B.n406 VSUBS 0.006114f
C447 B.n407 VSUBS 0.006114f
C448 B.n408 VSUBS 0.006114f
C449 B.n409 VSUBS 0.006114f
C450 B.n410 VSUBS 0.006114f
C451 B.n411 VSUBS 0.006114f
C452 B.n412 VSUBS 0.006114f
C453 B.n413 VSUBS 0.006114f
C454 B.n414 VSUBS 0.006114f
C455 B.n415 VSUBS 0.006114f
C456 B.n416 VSUBS 0.006114f
C457 B.n417 VSUBS 0.006114f
C458 B.n418 VSUBS 0.006114f
C459 B.n419 VSUBS 0.015004f
C460 B.n420 VSUBS 0.014308f
C461 B.n421 VSUBS 0.014308f
C462 B.n422 VSUBS 0.006114f
C463 B.n423 VSUBS 0.006114f
C464 B.n424 VSUBS 0.006114f
C465 B.n425 VSUBS 0.006114f
C466 B.n426 VSUBS 0.006114f
C467 B.n427 VSUBS 0.006114f
C468 B.n428 VSUBS 0.006114f
C469 B.n429 VSUBS 0.006114f
C470 B.n430 VSUBS 0.006114f
C471 B.n431 VSUBS 0.006114f
C472 B.n432 VSUBS 0.006114f
C473 B.n433 VSUBS 0.006114f
C474 B.n434 VSUBS 0.006114f
C475 B.n435 VSUBS 0.006114f
C476 B.n436 VSUBS 0.006114f
C477 B.n437 VSUBS 0.006114f
C478 B.n438 VSUBS 0.006114f
C479 B.n439 VSUBS 0.006114f
C480 B.n440 VSUBS 0.006114f
C481 B.n441 VSUBS 0.006114f
C482 B.n442 VSUBS 0.006114f
C483 B.n443 VSUBS 0.006114f
C484 B.n444 VSUBS 0.006114f
C485 B.n445 VSUBS 0.006114f
C486 B.n446 VSUBS 0.006114f
C487 B.n447 VSUBS 0.006114f
C488 B.n448 VSUBS 0.006114f
C489 B.n449 VSUBS 0.006114f
C490 B.n450 VSUBS 0.006114f
C491 B.n451 VSUBS 0.006114f
C492 B.n452 VSUBS 0.006114f
C493 B.n453 VSUBS 0.006114f
C494 B.n454 VSUBS 0.006114f
C495 B.n455 VSUBS 0.007979f
C496 B.n456 VSUBS 0.008499f
C497 B.n457 VSUBS 0.016902f
C498 VDD2.n0 VSUBS 0.025588f
C499 VDD2.n1 VSUBS 0.022505f
C500 VDD2.n2 VSUBS 0.012093f
C501 VDD2.n3 VSUBS 0.028584f
C502 VDD2.n4 VSUBS 0.012805f
C503 VDD2.n5 VSUBS 0.022505f
C504 VDD2.n6 VSUBS 0.012093f
C505 VDD2.n7 VSUBS 0.028584f
C506 VDD2.n8 VSUBS 0.012805f
C507 VDD2.n9 VSUBS 0.596287f
C508 VDD2.n10 VSUBS 0.012093f
C509 VDD2.t4 VSUBS 0.061189f
C510 VDD2.n11 VSUBS 0.104519f
C511 VDD2.n12 VSUBS 0.01818f
C512 VDD2.n13 VSUBS 0.021438f
C513 VDD2.n14 VSUBS 0.028584f
C514 VDD2.n15 VSUBS 0.012805f
C515 VDD2.n16 VSUBS 0.012093f
C516 VDD2.n17 VSUBS 0.022505f
C517 VDD2.n18 VSUBS 0.022505f
C518 VDD2.n19 VSUBS 0.012093f
C519 VDD2.n20 VSUBS 0.012805f
C520 VDD2.n21 VSUBS 0.028584f
C521 VDD2.n22 VSUBS 0.028584f
C522 VDD2.n23 VSUBS 0.012805f
C523 VDD2.n24 VSUBS 0.012093f
C524 VDD2.n25 VSUBS 0.022505f
C525 VDD2.n26 VSUBS 0.022505f
C526 VDD2.n27 VSUBS 0.012093f
C527 VDD2.n28 VSUBS 0.012805f
C528 VDD2.n29 VSUBS 0.028584f
C529 VDD2.n30 VSUBS 0.072128f
C530 VDD2.n31 VSUBS 0.012805f
C531 VDD2.n32 VSUBS 0.012093f
C532 VDD2.n33 VSUBS 0.053864f
C533 VDD2.n34 VSUBS 0.053764f
C534 VDD2.t2 VSUBS 0.120577f
C535 VDD2.t0 VSUBS 0.120577f
C536 VDD2.n35 VSUBS 0.828485f
C537 VDD2.n36 VSUBS 1.72493f
C538 VDD2.n37 VSUBS 0.025588f
C539 VDD2.n38 VSUBS 0.022505f
C540 VDD2.n39 VSUBS 0.012093f
C541 VDD2.n40 VSUBS 0.028584f
C542 VDD2.n41 VSUBS 0.012805f
C543 VDD2.n42 VSUBS 0.022505f
C544 VDD2.n43 VSUBS 0.012093f
C545 VDD2.n44 VSUBS 0.028584f
C546 VDD2.n45 VSUBS 0.012805f
C547 VDD2.n46 VSUBS 0.596287f
C548 VDD2.n47 VSUBS 0.012093f
C549 VDD2.t1 VSUBS 0.061189f
C550 VDD2.n48 VSUBS 0.104519f
C551 VDD2.n49 VSUBS 0.01818f
C552 VDD2.n50 VSUBS 0.021438f
C553 VDD2.n51 VSUBS 0.028584f
C554 VDD2.n52 VSUBS 0.012805f
C555 VDD2.n53 VSUBS 0.012093f
C556 VDD2.n54 VSUBS 0.022505f
C557 VDD2.n55 VSUBS 0.022505f
C558 VDD2.n56 VSUBS 0.012093f
C559 VDD2.n57 VSUBS 0.012805f
C560 VDD2.n58 VSUBS 0.028584f
C561 VDD2.n59 VSUBS 0.028584f
C562 VDD2.n60 VSUBS 0.012805f
C563 VDD2.n61 VSUBS 0.012093f
C564 VDD2.n62 VSUBS 0.022505f
C565 VDD2.n63 VSUBS 0.022505f
C566 VDD2.n64 VSUBS 0.012093f
C567 VDD2.n65 VSUBS 0.012805f
C568 VDD2.n66 VSUBS 0.028584f
C569 VDD2.n67 VSUBS 0.072128f
C570 VDD2.n68 VSUBS 0.012805f
C571 VDD2.n69 VSUBS 0.012093f
C572 VDD2.n70 VSUBS 0.053864f
C573 VDD2.n71 VSUBS 0.051983f
C574 VDD2.n72 VSUBS 1.55998f
C575 VDD2.t5 VSUBS 0.120577f
C576 VDD2.t3 VSUBS 0.120577f
C577 VDD2.n73 VSUBS 0.828463f
C578 VN.n0 VSUBS 0.293547f
C579 VN.t3 VSUBS 1.02914f
C580 VN.t1 VSUBS 1.1708f
C581 VN.n1 VSUBS 0.475776f
C582 VN.n2 VSUBS 0.494995f
C583 VN.n3 VSUBS 0.067149f
C584 VN.t5 VSUBS 1.11587f
C585 VN.n4 VSUBS 0.496461f
C586 VN.n5 VSUBS 0.049858f
C587 VN.n6 VSUBS 0.293547f
C588 VN.t0 VSUBS 1.02914f
C589 VN.t2 VSUBS 1.1708f
C590 VN.n7 VSUBS 0.475776f
C591 VN.n8 VSUBS 0.494995f
C592 VN.n9 VSUBS 0.067149f
C593 VN.t4 VSUBS 1.11587f
C594 VN.n10 VSUBS 0.496461f
C595 VN.n11 VSUBS 1.97445f
C596 VDD1.n0 VSUBS 0.025636f
C597 VDD1.n1 VSUBS 0.022547f
C598 VDD1.n2 VSUBS 0.012116f
C599 VDD1.n3 VSUBS 0.028637f
C600 VDD1.n4 VSUBS 0.012828f
C601 VDD1.n5 VSUBS 0.022547f
C602 VDD1.n6 VSUBS 0.012116f
C603 VDD1.n7 VSUBS 0.028637f
C604 VDD1.n8 VSUBS 0.012828f
C605 VDD1.n9 VSUBS 0.597395f
C606 VDD1.n10 VSUBS 0.012116f
C607 VDD1.t4 VSUBS 0.061303f
C608 VDD1.n11 VSUBS 0.104713f
C609 VDD1.n12 VSUBS 0.018214f
C610 VDD1.n13 VSUBS 0.021478f
C611 VDD1.n14 VSUBS 0.028637f
C612 VDD1.n15 VSUBS 0.012828f
C613 VDD1.n16 VSUBS 0.012116f
C614 VDD1.n17 VSUBS 0.022547f
C615 VDD1.n18 VSUBS 0.022547f
C616 VDD1.n19 VSUBS 0.012116f
C617 VDD1.n20 VSUBS 0.012828f
C618 VDD1.n21 VSUBS 0.028637f
C619 VDD1.n22 VSUBS 0.028637f
C620 VDD1.n23 VSUBS 0.012828f
C621 VDD1.n24 VSUBS 0.012116f
C622 VDD1.n25 VSUBS 0.022547f
C623 VDD1.n26 VSUBS 0.022547f
C624 VDD1.n27 VSUBS 0.012116f
C625 VDD1.n28 VSUBS 0.012828f
C626 VDD1.n29 VSUBS 0.028637f
C627 VDD1.n30 VSUBS 0.072262f
C628 VDD1.n31 VSUBS 0.012828f
C629 VDD1.n32 VSUBS 0.012116f
C630 VDD1.n33 VSUBS 0.053964f
C631 VDD1.n34 VSUBS 0.054242f
C632 VDD1.n35 VSUBS 0.025636f
C633 VDD1.n36 VSUBS 0.022547f
C634 VDD1.n37 VSUBS 0.012116f
C635 VDD1.n38 VSUBS 0.028637f
C636 VDD1.n39 VSUBS 0.012828f
C637 VDD1.n40 VSUBS 0.022547f
C638 VDD1.n41 VSUBS 0.012116f
C639 VDD1.n42 VSUBS 0.028637f
C640 VDD1.n43 VSUBS 0.012828f
C641 VDD1.n44 VSUBS 0.597395f
C642 VDD1.n45 VSUBS 0.012116f
C643 VDD1.t5 VSUBS 0.061303f
C644 VDD1.n46 VSUBS 0.104713f
C645 VDD1.n47 VSUBS 0.018214f
C646 VDD1.n48 VSUBS 0.021478f
C647 VDD1.n49 VSUBS 0.028637f
C648 VDD1.n50 VSUBS 0.012828f
C649 VDD1.n51 VSUBS 0.012116f
C650 VDD1.n52 VSUBS 0.022547f
C651 VDD1.n53 VSUBS 0.022547f
C652 VDD1.n54 VSUBS 0.012116f
C653 VDD1.n55 VSUBS 0.012828f
C654 VDD1.n56 VSUBS 0.028637f
C655 VDD1.n57 VSUBS 0.028637f
C656 VDD1.n58 VSUBS 0.012828f
C657 VDD1.n59 VSUBS 0.012116f
C658 VDD1.n60 VSUBS 0.022547f
C659 VDD1.n61 VSUBS 0.022547f
C660 VDD1.n62 VSUBS 0.012116f
C661 VDD1.n63 VSUBS 0.012828f
C662 VDD1.n64 VSUBS 0.028637f
C663 VDD1.n65 VSUBS 0.072262f
C664 VDD1.n66 VSUBS 0.012828f
C665 VDD1.n67 VSUBS 0.012116f
C666 VDD1.n68 VSUBS 0.053964f
C667 VDD1.n69 VSUBS 0.053864f
C668 VDD1.t0 VSUBS 0.120801f
C669 VDD1.t2 VSUBS 0.120801f
C670 VDD1.n70 VSUBS 0.830025f
C671 VDD1.n71 VSUBS 1.80304f
C672 VDD1.t1 VSUBS 0.120801f
C673 VDD1.t3 VSUBS 0.120801f
C674 VDD1.n72 VSUBS 0.828667f
C675 VDD1.n73 VSUBS 1.94939f
C676 VTAIL.t0 VSUBS 0.151033f
C677 VTAIL.t9 VSUBS 0.151033f
C678 VTAIL.n0 VSUBS 0.929088f
C679 VTAIL.n1 VSUBS 0.671605f
C680 VTAIL.n2 VSUBS 0.032051f
C681 VTAIL.n3 VSUBS 0.02819f
C682 VTAIL.n4 VSUBS 0.015148f
C683 VTAIL.n5 VSUBS 0.035804f
C684 VTAIL.n6 VSUBS 0.016039f
C685 VTAIL.n7 VSUBS 0.02819f
C686 VTAIL.n8 VSUBS 0.015148f
C687 VTAIL.n9 VSUBS 0.035804f
C688 VTAIL.n10 VSUBS 0.016039f
C689 VTAIL.n11 VSUBS 0.746901f
C690 VTAIL.n12 VSUBS 0.015148f
C691 VTAIL.t3 VSUBS 0.076644f
C692 VTAIL.n13 VSUBS 0.130919f
C693 VTAIL.n14 VSUBS 0.022772f
C694 VTAIL.n15 VSUBS 0.026853f
C695 VTAIL.n16 VSUBS 0.035804f
C696 VTAIL.n17 VSUBS 0.016039f
C697 VTAIL.n18 VSUBS 0.015148f
C698 VTAIL.n19 VSUBS 0.02819f
C699 VTAIL.n20 VSUBS 0.02819f
C700 VTAIL.n21 VSUBS 0.015148f
C701 VTAIL.n22 VSUBS 0.016039f
C702 VTAIL.n23 VSUBS 0.035804f
C703 VTAIL.n24 VSUBS 0.035804f
C704 VTAIL.n25 VSUBS 0.016039f
C705 VTAIL.n26 VSUBS 0.015148f
C706 VTAIL.n27 VSUBS 0.02819f
C707 VTAIL.n28 VSUBS 0.02819f
C708 VTAIL.n29 VSUBS 0.015148f
C709 VTAIL.n30 VSUBS 0.016039f
C710 VTAIL.n31 VSUBS 0.035804f
C711 VTAIL.n32 VSUBS 0.090346f
C712 VTAIL.n33 VSUBS 0.016039f
C713 VTAIL.n34 VSUBS 0.015148f
C714 VTAIL.n35 VSUBS 0.067469f
C715 VTAIL.n36 VSUBS 0.045667f
C716 VTAIL.n37 VSUBS 0.232496f
C717 VTAIL.t2 VSUBS 0.151033f
C718 VTAIL.t6 VSUBS 0.151033f
C719 VTAIL.n38 VSUBS 0.929088f
C720 VTAIL.n39 VSUBS 1.78413f
C721 VTAIL.t10 VSUBS 0.151033f
C722 VTAIL.t1 VSUBS 0.151033f
C723 VTAIL.n40 VSUBS 0.929094f
C724 VTAIL.n41 VSUBS 1.78412f
C725 VTAIL.n42 VSUBS 0.032051f
C726 VTAIL.n43 VSUBS 0.02819f
C727 VTAIL.n44 VSUBS 0.015148f
C728 VTAIL.n45 VSUBS 0.035804f
C729 VTAIL.n46 VSUBS 0.016039f
C730 VTAIL.n47 VSUBS 0.02819f
C731 VTAIL.n48 VSUBS 0.015148f
C732 VTAIL.n49 VSUBS 0.035804f
C733 VTAIL.n50 VSUBS 0.016039f
C734 VTAIL.n51 VSUBS 0.746901f
C735 VTAIL.n52 VSUBS 0.015148f
C736 VTAIL.t8 VSUBS 0.076644f
C737 VTAIL.n53 VSUBS 0.130919f
C738 VTAIL.n54 VSUBS 0.022772f
C739 VTAIL.n55 VSUBS 0.026853f
C740 VTAIL.n56 VSUBS 0.035804f
C741 VTAIL.n57 VSUBS 0.016039f
C742 VTAIL.n58 VSUBS 0.015148f
C743 VTAIL.n59 VSUBS 0.02819f
C744 VTAIL.n60 VSUBS 0.02819f
C745 VTAIL.n61 VSUBS 0.015148f
C746 VTAIL.n62 VSUBS 0.016039f
C747 VTAIL.n63 VSUBS 0.035804f
C748 VTAIL.n64 VSUBS 0.035804f
C749 VTAIL.n65 VSUBS 0.016039f
C750 VTAIL.n66 VSUBS 0.015148f
C751 VTAIL.n67 VSUBS 0.02819f
C752 VTAIL.n68 VSUBS 0.02819f
C753 VTAIL.n69 VSUBS 0.015148f
C754 VTAIL.n70 VSUBS 0.016039f
C755 VTAIL.n71 VSUBS 0.035804f
C756 VTAIL.n72 VSUBS 0.090346f
C757 VTAIL.n73 VSUBS 0.016039f
C758 VTAIL.n74 VSUBS 0.015148f
C759 VTAIL.n75 VSUBS 0.067469f
C760 VTAIL.n76 VSUBS 0.045667f
C761 VTAIL.n77 VSUBS 0.232496f
C762 VTAIL.t5 VSUBS 0.151033f
C763 VTAIL.t4 VSUBS 0.151033f
C764 VTAIL.n78 VSUBS 0.929094f
C765 VTAIL.n79 VSUBS 0.748533f
C766 VTAIL.n80 VSUBS 0.032051f
C767 VTAIL.n81 VSUBS 0.02819f
C768 VTAIL.n82 VSUBS 0.015148f
C769 VTAIL.n83 VSUBS 0.035804f
C770 VTAIL.n84 VSUBS 0.016039f
C771 VTAIL.n85 VSUBS 0.02819f
C772 VTAIL.n86 VSUBS 0.015148f
C773 VTAIL.n87 VSUBS 0.035804f
C774 VTAIL.n88 VSUBS 0.016039f
C775 VTAIL.n89 VSUBS 0.746901f
C776 VTAIL.n90 VSUBS 0.015148f
C777 VTAIL.t7 VSUBS 0.076644f
C778 VTAIL.n91 VSUBS 0.130919f
C779 VTAIL.n92 VSUBS 0.022772f
C780 VTAIL.n93 VSUBS 0.026853f
C781 VTAIL.n94 VSUBS 0.035804f
C782 VTAIL.n95 VSUBS 0.016039f
C783 VTAIL.n96 VSUBS 0.015148f
C784 VTAIL.n97 VSUBS 0.02819f
C785 VTAIL.n98 VSUBS 0.02819f
C786 VTAIL.n99 VSUBS 0.015148f
C787 VTAIL.n100 VSUBS 0.016039f
C788 VTAIL.n101 VSUBS 0.035804f
C789 VTAIL.n102 VSUBS 0.035804f
C790 VTAIL.n103 VSUBS 0.016039f
C791 VTAIL.n104 VSUBS 0.015148f
C792 VTAIL.n105 VSUBS 0.02819f
C793 VTAIL.n106 VSUBS 0.02819f
C794 VTAIL.n107 VSUBS 0.015148f
C795 VTAIL.n108 VSUBS 0.016039f
C796 VTAIL.n109 VSUBS 0.035804f
C797 VTAIL.n110 VSUBS 0.090346f
C798 VTAIL.n111 VSUBS 0.016039f
C799 VTAIL.n112 VSUBS 0.015148f
C800 VTAIL.n113 VSUBS 0.067469f
C801 VTAIL.n114 VSUBS 0.045667f
C802 VTAIL.n115 VSUBS 1.15846f
C803 VTAIL.n116 VSUBS 0.032051f
C804 VTAIL.n117 VSUBS 0.02819f
C805 VTAIL.n118 VSUBS 0.015148f
C806 VTAIL.n119 VSUBS 0.035804f
C807 VTAIL.n120 VSUBS 0.016039f
C808 VTAIL.n121 VSUBS 0.02819f
C809 VTAIL.n122 VSUBS 0.015148f
C810 VTAIL.n123 VSUBS 0.035804f
C811 VTAIL.n124 VSUBS 0.016039f
C812 VTAIL.n125 VSUBS 0.746901f
C813 VTAIL.n126 VSUBS 0.015148f
C814 VTAIL.t11 VSUBS 0.076644f
C815 VTAIL.n127 VSUBS 0.130919f
C816 VTAIL.n128 VSUBS 0.022772f
C817 VTAIL.n129 VSUBS 0.026853f
C818 VTAIL.n130 VSUBS 0.035804f
C819 VTAIL.n131 VSUBS 0.016039f
C820 VTAIL.n132 VSUBS 0.015148f
C821 VTAIL.n133 VSUBS 0.02819f
C822 VTAIL.n134 VSUBS 0.02819f
C823 VTAIL.n135 VSUBS 0.015148f
C824 VTAIL.n136 VSUBS 0.016039f
C825 VTAIL.n137 VSUBS 0.035804f
C826 VTAIL.n138 VSUBS 0.035804f
C827 VTAIL.n139 VSUBS 0.016039f
C828 VTAIL.n140 VSUBS 0.015148f
C829 VTAIL.n141 VSUBS 0.02819f
C830 VTAIL.n142 VSUBS 0.02819f
C831 VTAIL.n143 VSUBS 0.015148f
C832 VTAIL.n144 VSUBS 0.016039f
C833 VTAIL.n145 VSUBS 0.035804f
C834 VTAIL.n146 VSUBS 0.090346f
C835 VTAIL.n147 VSUBS 0.016039f
C836 VTAIL.n148 VSUBS 0.015148f
C837 VTAIL.n149 VSUBS 0.067469f
C838 VTAIL.n150 VSUBS 0.045667f
C839 VTAIL.n151 VSUBS 1.12576f
C840 VP.n0 VSUBS 0.073909f
C841 VP.t5 VSUBS 1.07072f
C842 VP.n1 VSUBS 0.069863f
C843 VP.n2 VSUBS 0.305409f
C844 VP.t2 VSUBS 1.16096f
C845 VP.t4 VSUBS 1.07072f
C846 VP.t1 VSUBS 1.21811f
C847 VP.n3 VSUBS 0.495002f
C848 VP.n4 VSUBS 0.514998f
C849 VP.n5 VSUBS 0.069863f
C850 VP.n6 VSUBS 0.516523f
C851 VP.n7 VSUBS 2.02273f
C852 VP.t0 VSUBS 1.16096f
C853 VP.n8 VSUBS 0.516523f
C854 VP.n9 VSUBS 2.07408f
C855 VP.n10 VSUBS 0.073909f
C856 VP.n11 VSUBS 0.055388f
C857 VP.n12 VSUBS 0.478074f
C858 VP.n13 VSUBS 0.069863f
C859 VP.t3 VSUBS 1.16096f
C860 VP.n14 VSUBS 0.516523f
C861 VP.n15 VSUBS 0.051873f
.ends

