* NGSPICE file created from diff_pair_sample_1741.ext - technology: sky130A

.subckt diff_pair_sample_1741 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1.12
X1 VTAIL.t9 VN.t1 VDD2.t4 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1.12
X2 VDD2.t3 VN.t2 VTAIL.t8 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1.12
X3 B.t11 B.t9 B.t10 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1.12
X4 VDD2.t2 VN.t3 VTAIL.t11 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1.12
X5 VTAIL.t0 VP.t0 VDD1.t5 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1.12
X6 B.t8 B.t6 B.t7 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1.12
X7 VDD2.t1 VN.t4 VTAIL.t6 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1.12
X8 B.t5 B.t3 B.t4 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1.12
X9 VDD1.t4 VP.t1 VTAIL.t1 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1.12
X10 VDD1.t3 VP.t2 VTAIL.t4 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1.12
X11 VTAIL.t5 VP.t3 VDD1.t2 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1.12
X12 VDD1.t1 VP.t4 VTAIL.t2 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1.12
X13 VTAIL.t7 VN.t5 VDD2.t0 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1.12
X14 VDD1.t0 VP.t5 VTAIL.t3 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1.12
X15 B.t2 B.t0 B.t1 w_n2130_n2368# sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1.12
R0 VN.n1 VN.t3 208.909
R1 VN.n7 VN.t4 208.909
R2 VN.n4 VN.t0 185.7
R3 VN.n10 VN.t2 185.7
R4 VN.n9 VN.n6 161.3
R5 VN.n3 VN.n0 161.3
R6 VN.n2 VN.t1 150.625
R7 VN.n8 VN.t5 150.625
R8 VN.n11 VN.n10 80.6037
R9 VN.n5 VN.n4 80.6037
R10 VN.n4 VN.n3 51.1515
R11 VN.n10 VN.n9 51.1515
R12 VN VN.n11 39.5786
R13 VN.n2 VN.n1 32.8731
R14 VN.n8 VN.n7 32.8731
R15 VN.n7 VN.n6 28.0424
R16 VN.n1 VN.n0 28.0424
R17 VN.n3 VN.n2 24.5923
R18 VN.n9 VN.n8 24.5923
R19 VN.n11 VN.n6 0.285035
R20 VN.n5 VN.n0 0.285035
R21 VN VN.n5 0.146778
R22 VTAIL.n7 VTAIL.t6 73.1794
R23 VTAIL.n11 VTAIL.t10 73.1792
R24 VTAIL.n2 VTAIL.t2 73.1792
R25 VTAIL.n10 VTAIL.t1 73.1792
R26 VTAIL.n9 VTAIL.n8 68.5358
R27 VTAIL.n6 VTAIL.n5 68.5358
R28 VTAIL.n1 VTAIL.n0 68.5358
R29 VTAIL.n4 VTAIL.n3 68.5358
R30 VTAIL.n6 VTAIL.n4 20.9014
R31 VTAIL.n11 VTAIL.n10 19.6514
R32 VTAIL.n0 VTAIL.t11 4.64407
R33 VTAIL.n0 VTAIL.t9 4.64407
R34 VTAIL.n3 VTAIL.t4 4.64407
R35 VTAIL.n3 VTAIL.t5 4.64407
R36 VTAIL.n8 VTAIL.t3 4.64407
R37 VTAIL.n8 VTAIL.t0 4.64407
R38 VTAIL.n5 VTAIL.t8 4.64407
R39 VTAIL.n5 VTAIL.t7 4.64407
R40 VTAIL.n7 VTAIL.n6 1.2505
R41 VTAIL.n10 VTAIL.n9 1.2505
R42 VTAIL.n4 VTAIL.n2 1.2505
R43 VTAIL.n9 VTAIL.n7 1.09533
R44 VTAIL.n2 VTAIL.n1 1.09533
R45 VTAIL VTAIL.n11 0.87981
R46 VTAIL VTAIL.n1 0.37119
R47 VDD2.n1 VDD2.t2 90.7401
R48 VDD2.n2 VDD2.t3 89.8582
R49 VDD2.n1 VDD2.n0 85.4717
R50 VDD2 VDD2.n3 85.4687
R51 VDD2.n2 VDD2.n1 33.8123
R52 VDD2.n3 VDD2.t0 4.64407
R53 VDD2.n3 VDD2.t1 4.64407
R54 VDD2.n0 VDD2.t4 4.64407
R55 VDD2.n0 VDD2.t5 4.64407
R56 VDD2 VDD2.n2 0.99619
R57 B.n333 B.n50 585
R58 B.n335 B.n334 585
R59 B.n336 B.n49 585
R60 B.n338 B.n337 585
R61 B.n339 B.n48 585
R62 B.n341 B.n340 585
R63 B.n342 B.n47 585
R64 B.n344 B.n343 585
R65 B.n345 B.n46 585
R66 B.n347 B.n346 585
R67 B.n348 B.n45 585
R68 B.n350 B.n349 585
R69 B.n351 B.n44 585
R70 B.n353 B.n352 585
R71 B.n354 B.n43 585
R72 B.n356 B.n355 585
R73 B.n357 B.n42 585
R74 B.n359 B.n358 585
R75 B.n360 B.n41 585
R76 B.n362 B.n361 585
R77 B.n363 B.n40 585
R78 B.n365 B.n364 585
R79 B.n366 B.n39 585
R80 B.n368 B.n367 585
R81 B.n369 B.n38 585
R82 B.n371 B.n370 585
R83 B.n372 B.n35 585
R84 B.n375 B.n374 585
R85 B.n376 B.n34 585
R86 B.n378 B.n377 585
R87 B.n379 B.n33 585
R88 B.n381 B.n380 585
R89 B.n382 B.n32 585
R90 B.n384 B.n383 585
R91 B.n385 B.n31 585
R92 B.n387 B.n386 585
R93 B.n389 B.n388 585
R94 B.n390 B.n27 585
R95 B.n392 B.n391 585
R96 B.n393 B.n26 585
R97 B.n395 B.n394 585
R98 B.n396 B.n25 585
R99 B.n398 B.n397 585
R100 B.n399 B.n24 585
R101 B.n401 B.n400 585
R102 B.n402 B.n23 585
R103 B.n404 B.n403 585
R104 B.n405 B.n22 585
R105 B.n407 B.n406 585
R106 B.n408 B.n21 585
R107 B.n410 B.n409 585
R108 B.n411 B.n20 585
R109 B.n413 B.n412 585
R110 B.n414 B.n19 585
R111 B.n416 B.n415 585
R112 B.n417 B.n18 585
R113 B.n419 B.n418 585
R114 B.n420 B.n17 585
R115 B.n422 B.n421 585
R116 B.n423 B.n16 585
R117 B.n425 B.n424 585
R118 B.n426 B.n15 585
R119 B.n428 B.n427 585
R120 B.n332 B.n331 585
R121 B.n330 B.n51 585
R122 B.n329 B.n328 585
R123 B.n327 B.n52 585
R124 B.n326 B.n325 585
R125 B.n324 B.n53 585
R126 B.n323 B.n322 585
R127 B.n321 B.n54 585
R128 B.n320 B.n319 585
R129 B.n318 B.n55 585
R130 B.n317 B.n316 585
R131 B.n315 B.n56 585
R132 B.n314 B.n313 585
R133 B.n312 B.n57 585
R134 B.n311 B.n310 585
R135 B.n309 B.n58 585
R136 B.n308 B.n307 585
R137 B.n306 B.n59 585
R138 B.n305 B.n304 585
R139 B.n303 B.n60 585
R140 B.n302 B.n301 585
R141 B.n300 B.n61 585
R142 B.n299 B.n298 585
R143 B.n297 B.n62 585
R144 B.n296 B.n295 585
R145 B.n294 B.n63 585
R146 B.n293 B.n292 585
R147 B.n291 B.n64 585
R148 B.n290 B.n289 585
R149 B.n288 B.n65 585
R150 B.n287 B.n286 585
R151 B.n285 B.n66 585
R152 B.n284 B.n283 585
R153 B.n282 B.n67 585
R154 B.n281 B.n280 585
R155 B.n279 B.n68 585
R156 B.n278 B.n277 585
R157 B.n276 B.n69 585
R158 B.n275 B.n274 585
R159 B.n273 B.n70 585
R160 B.n272 B.n271 585
R161 B.n270 B.n71 585
R162 B.n269 B.n268 585
R163 B.n267 B.n72 585
R164 B.n266 B.n265 585
R165 B.n264 B.n73 585
R166 B.n263 B.n262 585
R167 B.n261 B.n74 585
R168 B.n260 B.n259 585
R169 B.n258 B.n75 585
R170 B.n257 B.n256 585
R171 B.n161 B.n160 585
R172 B.n162 B.n111 585
R173 B.n164 B.n163 585
R174 B.n165 B.n110 585
R175 B.n167 B.n166 585
R176 B.n168 B.n109 585
R177 B.n170 B.n169 585
R178 B.n171 B.n108 585
R179 B.n173 B.n172 585
R180 B.n174 B.n107 585
R181 B.n176 B.n175 585
R182 B.n177 B.n106 585
R183 B.n179 B.n178 585
R184 B.n180 B.n105 585
R185 B.n182 B.n181 585
R186 B.n183 B.n104 585
R187 B.n185 B.n184 585
R188 B.n186 B.n103 585
R189 B.n188 B.n187 585
R190 B.n189 B.n102 585
R191 B.n191 B.n190 585
R192 B.n192 B.n101 585
R193 B.n194 B.n193 585
R194 B.n195 B.n100 585
R195 B.n197 B.n196 585
R196 B.n198 B.n99 585
R197 B.n200 B.n199 585
R198 B.n202 B.n201 585
R199 B.n203 B.n95 585
R200 B.n205 B.n204 585
R201 B.n206 B.n94 585
R202 B.n208 B.n207 585
R203 B.n209 B.n93 585
R204 B.n211 B.n210 585
R205 B.n212 B.n92 585
R206 B.n214 B.n213 585
R207 B.n216 B.n89 585
R208 B.n218 B.n217 585
R209 B.n219 B.n88 585
R210 B.n221 B.n220 585
R211 B.n222 B.n87 585
R212 B.n224 B.n223 585
R213 B.n225 B.n86 585
R214 B.n227 B.n226 585
R215 B.n228 B.n85 585
R216 B.n230 B.n229 585
R217 B.n231 B.n84 585
R218 B.n233 B.n232 585
R219 B.n234 B.n83 585
R220 B.n236 B.n235 585
R221 B.n237 B.n82 585
R222 B.n239 B.n238 585
R223 B.n240 B.n81 585
R224 B.n242 B.n241 585
R225 B.n243 B.n80 585
R226 B.n245 B.n244 585
R227 B.n246 B.n79 585
R228 B.n248 B.n247 585
R229 B.n249 B.n78 585
R230 B.n251 B.n250 585
R231 B.n252 B.n77 585
R232 B.n254 B.n253 585
R233 B.n255 B.n76 585
R234 B.n159 B.n112 585
R235 B.n158 B.n157 585
R236 B.n156 B.n113 585
R237 B.n155 B.n154 585
R238 B.n153 B.n114 585
R239 B.n152 B.n151 585
R240 B.n150 B.n115 585
R241 B.n149 B.n148 585
R242 B.n147 B.n116 585
R243 B.n146 B.n145 585
R244 B.n144 B.n117 585
R245 B.n143 B.n142 585
R246 B.n141 B.n118 585
R247 B.n140 B.n139 585
R248 B.n138 B.n119 585
R249 B.n137 B.n136 585
R250 B.n135 B.n120 585
R251 B.n134 B.n133 585
R252 B.n132 B.n121 585
R253 B.n131 B.n130 585
R254 B.n129 B.n122 585
R255 B.n128 B.n127 585
R256 B.n126 B.n123 585
R257 B.n125 B.n124 585
R258 B.n2 B.n0 585
R259 B.n465 B.n1 585
R260 B.n464 B.n463 585
R261 B.n462 B.n3 585
R262 B.n461 B.n460 585
R263 B.n459 B.n4 585
R264 B.n458 B.n457 585
R265 B.n456 B.n5 585
R266 B.n455 B.n454 585
R267 B.n453 B.n6 585
R268 B.n452 B.n451 585
R269 B.n450 B.n7 585
R270 B.n449 B.n448 585
R271 B.n447 B.n8 585
R272 B.n446 B.n445 585
R273 B.n444 B.n9 585
R274 B.n443 B.n442 585
R275 B.n441 B.n10 585
R276 B.n440 B.n439 585
R277 B.n438 B.n11 585
R278 B.n437 B.n436 585
R279 B.n435 B.n12 585
R280 B.n434 B.n433 585
R281 B.n432 B.n13 585
R282 B.n431 B.n430 585
R283 B.n429 B.n14 585
R284 B.n467 B.n466 585
R285 B.n160 B.n159 559.769
R286 B.n429 B.n428 559.769
R287 B.n256 B.n255 559.769
R288 B.n333 B.n332 559.769
R289 B.n90 B.t6 354.303
R290 B.n96 B.t9 354.303
R291 B.n28 B.t3 354.303
R292 B.n36 B.t0 354.303
R293 B.n159 B.n158 163.367
R294 B.n158 B.n113 163.367
R295 B.n154 B.n113 163.367
R296 B.n154 B.n153 163.367
R297 B.n153 B.n152 163.367
R298 B.n152 B.n115 163.367
R299 B.n148 B.n115 163.367
R300 B.n148 B.n147 163.367
R301 B.n147 B.n146 163.367
R302 B.n146 B.n117 163.367
R303 B.n142 B.n117 163.367
R304 B.n142 B.n141 163.367
R305 B.n141 B.n140 163.367
R306 B.n140 B.n119 163.367
R307 B.n136 B.n119 163.367
R308 B.n136 B.n135 163.367
R309 B.n135 B.n134 163.367
R310 B.n134 B.n121 163.367
R311 B.n130 B.n121 163.367
R312 B.n130 B.n129 163.367
R313 B.n129 B.n128 163.367
R314 B.n128 B.n123 163.367
R315 B.n124 B.n123 163.367
R316 B.n124 B.n2 163.367
R317 B.n466 B.n2 163.367
R318 B.n466 B.n465 163.367
R319 B.n465 B.n464 163.367
R320 B.n464 B.n3 163.367
R321 B.n460 B.n3 163.367
R322 B.n460 B.n459 163.367
R323 B.n459 B.n458 163.367
R324 B.n458 B.n5 163.367
R325 B.n454 B.n5 163.367
R326 B.n454 B.n453 163.367
R327 B.n453 B.n452 163.367
R328 B.n452 B.n7 163.367
R329 B.n448 B.n7 163.367
R330 B.n448 B.n447 163.367
R331 B.n447 B.n446 163.367
R332 B.n446 B.n9 163.367
R333 B.n442 B.n9 163.367
R334 B.n442 B.n441 163.367
R335 B.n441 B.n440 163.367
R336 B.n440 B.n11 163.367
R337 B.n436 B.n11 163.367
R338 B.n436 B.n435 163.367
R339 B.n435 B.n434 163.367
R340 B.n434 B.n13 163.367
R341 B.n430 B.n13 163.367
R342 B.n430 B.n429 163.367
R343 B.n160 B.n111 163.367
R344 B.n164 B.n111 163.367
R345 B.n165 B.n164 163.367
R346 B.n166 B.n165 163.367
R347 B.n166 B.n109 163.367
R348 B.n170 B.n109 163.367
R349 B.n171 B.n170 163.367
R350 B.n172 B.n171 163.367
R351 B.n172 B.n107 163.367
R352 B.n176 B.n107 163.367
R353 B.n177 B.n176 163.367
R354 B.n178 B.n177 163.367
R355 B.n178 B.n105 163.367
R356 B.n182 B.n105 163.367
R357 B.n183 B.n182 163.367
R358 B.n184 B.n183 163.367
R359 B.n184 B.n103 163.367
R360 B.n188 B.n103 163.367
R361 B.n189 B.n188 163.367
R362 B.n190 B.n189 163.367
R363 B.n190 B.n101 163.367
R364 B.n194 B.n101 163.367
R365 B.n195 B.n194 163.367
R366 B.n196 B.n195 163.367
R367 B.n196 B.n99 163.367
R368 B.n200 B.n99 163.367
R369 B.n201 B.n200 163.367
R370 B.n201 B.n95 163.367
R371 B.n205 B.n95 163.367
R372 B.n206 B.n205 163.367
R373 B.n207 B.n206 163.367
R374 B.n207 B.n93 163.367
R375 B.n211 B.n93 163.367
R376 B.n212 B.n211 163.367
R377 B.n213 B.n212 163.367
R378 B.n213 B.n89 163.367
R379 B.n218 B.n89 163.367
R380 B.n219 B.n218 163.367
R381 B.n220 B.n219 163.367
R382 B.n220 B.n87 163.367
R383 B.n224 B.n87 163.367
R384 B.n225 B.n224 163.367
R385 B.n226 B.n225 163.367
R386 B.n226 B.n85 163.367
R387 B.n230 B.n85 163.367
R388 B.n231 B.n230 163.367
R389 B.n232 B.n231 163.367
R390 B.n232 B.n83 163.367
R391 B.n236 B.n83 163.367
R392 B.n237 B.n236 163.367
R393 B.n238 B.n237 163.367
R394 B.n238 B.n81 163.367
R395 B.n242 B.n81 163.367
R396 B.n243 B.n242 163.367
R397 B.n244 B.n243 163.367
R398 B.n244 B.n79 163.367
R399 B.n248 B.n79 163.367
R400 B.n249 B.n248 163.367
R401 B.n250 B.n249 163.367
R402 B.n250 B.n77 163.367
R403 B.n254 B.n77 163.367
R404 B.n255 B.n254 163.367
R405 B.n256 B.n75 163.367
R406 B.n260 B.n75 163.367
R407 B.n261 B.n260 163.367
R408 B.n262 B.n261 163.367
R409 B.n262 B.n73 163.367
R410 B.n266 B.n73 163.367
R411 B.n267 B.n266 163.367
R412 B.n268 B.n267 163.367
R413 B.n268 B.n71 163.367
R414 B.n272 B.n71 163.367
R415 B.n273 B.n272 163.367
R416 B.n274 B.n273 163.367
R417 B.n274 B.n69 163.367
R418 B.n278 B.n69 163.367
R419 B.n279 B.n278 163.367
R420 B.n280 B.n279 163.367
R421 B.n280 B.n67 163.367
R422 B.n284 B.n67 163.367
R423 B.n285 B.n284 163.367
R424 B.n286 B.n285 163.367
R425 B.n286 B.n65 163.367
R426 B.n290 B.n65 163.367
R427 B.n291 B.n290 163.367
R428 B.n292 B.n291 163.367
R429 B.n292 B.n63 163.367
R430 B.n296 B.n63 163.367
R431 B.n297 B.n296 163.367
R432 B.n298 B.n297 163.367
R433 B.n298 B.n61 163.367
R434 B.n302 B.n61 163.367
R435 B.n303 B.n302 163.367
R436 B.n304 B.n303 163.367
R437 B.n304 B.n59 163.367
R438 B.n308 B.n59 163.367
R439 B.n309 B.n308 163.367
R440 B.n310 B.n309 163.367
R441 B.n310 B.n57 163.367
R442 B.n314 B.n57 163.367
R443 B.n315 B.n314 163.367
R444 B.n316 B.n315 163.367
R445 B.n316 B.n55 163.367
R446 B.n320 B.n55 163.367
R447 B.n321 B.n320 163.367
R448 B.n322 B.n321 163.367
R449 B.n322 B.n53 163.367
R450 B.n326 B.n53 163.367
R451 B.n327 B.n326 163.367
R452 B.n328 B.n327 163.367
R453 B.n328 B.n51 163.367
R454 B.n332 B.n51 163.367
R455 B.n428 B.n15 163.367
R456 B.n424 B.n15 163.367
R457 B.n424 B.n423 163.367
R458 B.n423 B.n422 163.367
R459 B.n422 B.n17 163.367
R460 B.n418 B.n17 163.367
R461 B.n418 B.n417 163.367
R462 B.n417 B.n416 163.367
R463 B.n416 B.n19 163.367
R464 B.n412 B.n19 163.367
R465 B.n412 B.n411 163.367
R466 B.n411 B.n410 163.367
R467 B.n410 B.n21 163.367
R468 B.n406 B.n21 163.367
R469 B.n406 B.n405 163.367
R470 B.n405 B.n404 163.367
R471 B.n404 B.n23 163.367
R472 B.n400 B.n23 163.367
R473 B.n400 B.n399 163.367
R474 B.n399 B.n398 163.367
R475 B.n398 B.n25 163.367
R476 B.n394 B.n25 163.367
R477 B.n394 B.n393 163.367
R478 B.n393 B.n392 163.367
R479 B.n392 B.n27 163.367
R480 B.n388 B.n27 163.367
R481 B.n388 B.n387 163.367
R482 B.n387 B.n31 163.367
R483 B.n383 B.n31 163.367
R484 B.n383 B.n382 163.367
R485 B.n382 B.n381 163.367
R486 B.n381 B.n33 163.367
R487 B.n377 B.n33 163.367
R488 B.n377 B.n376 163.367
R489 B.n376 B.n375 163.367
R490 B.n375 B.n35 163.367
R491 B.n370 B.n35 163.367
R492 B.n370 B.n369 163.367
R493 B.n369 B.n368 163.367
R494 B.n368 B.n39 163.367
R495 B.n364 B.n39 163.367
R496 B.n364 B.n363 163.367
R497 B.n363 B.n362 163.367
R498 B.n362 B.n41 163.367
R499 B.n358 B.n41 163.367
R500 B.n358 B.n357 163.367
R501 B.n357 B.n356 163.367
R502 B.n356 B.n43 163.367
R503 B.n352 B.n43 163.367
R504 B.n352 B.n351 163.367
R505 B.n351 B.n350 163.367
R506 B.n350 B.n45 163.367
R507 B.n346 B.n45 163.367
R508 B.n346 B.n345 163.367
R509 B.n345 B.n344 163.367
R510 B.n344 B.n47 163.367
R511 B.n340 B.n47 163.367
R512 B.n340 B.n339 163.367
R513 B.n339 B.n338 163.367
R514 B.n338 B.n49 163.367
R515 B.n334 B.n49 163.367
R516 B.n334 B.n333 163.367
R517 B.n90 B.t8 141.618
R518 B.n36 B.t1 141.618
R519 B.n96 B.t11 141.609
R520 B.n28 B.t4 141.609
R521 B.n91 B.t7 113.496
R522 B.n37 B.t2 113.496
R523 B.n97 B.t10 113.489
R524 B.n29 B.t5 113.489
R525 B.n215 B.n91 59.5399
R526 B.n98 B.n97 59.5399
R527 B.n30 B.n29 59.5399
R528 B.n373 B.n37 59.5399
R529 B.n427 B.n14 36.3712
R530 B.n331 B.n50 36.3712
R531 B.n257 B.n76 36.3712
R532 B.n161 B.n112 36.3712
R533 B.n91 B.n90 28.1217
R534 B.n97 B.n96 28.1217
R535 B.n29 B.n28 28.1217
R536 B.n37 B.n36 28.1217
R537 B B.n467 18.0485
R538 B.n427 B.n426 10.6151
R539 B.n426 B.n425 10.6151
R540 B.n425 B.n16 10.6151
R541 B.n421 B.n16 10.6151
R542 B.n421 B.n420 10.6151
R543 B.n420 B.n419 10.6151
R544 B.n419 B.n18 10.6151
R545 B.n415 B.n18 10.6151
R546 B.n415 B.n414 10.6151
R547 B.n414 B.n413 10.6151
R548 B.n413 B.n20 10.6151
R549 B.n409 B.n20 10.6151
R550 B.n409 B.n408 10.6151
R551 B.n408 B.n407 10.6151
R552 B.n407 B.n22 10.6151
R553 B.n403 B.n22 10.6151
R554 B.n403 B.n402 10.6151
R555 B.n402 B.n401 10.6151
R556 B.n401 B.n24 10.6151
R557 B.n397 B.n24 10.6151
R558 B.n397 B.n396 10.6151
R559 B.n396 B.n395 10.6151
R560 B.n395 B.n26 10.6151
R561 B.n391 B.n26 10.6151
R562 B.n391 B.n390 10.6151
R563 B.n390 B.n389 10.6151
R564 B.n386 B.n385 10.6151
R565 B.n385 B.n384 10.6151
R566 B.n384 B.n32 10.6151
R567 B.n380 B.n32 10.6151
R568 B.n380 B.n379 10.6151
R569 B.n379 B.n378 10.6151
R570 B.n378 B.n34 10.6151
R571 B.n374 B.n34 10.6151
R572 B.n372 B.n371 10.6151
R573 B.n371 B.n38 10.6151
R574 B.n367 B.n38 10.6151
R575 B.n367 B.n366 10.6151
R576 B.n366 B.n365 10.6151
R577 B.n365 B.n40 10.6151
R578 B.n361 B.n40 10.6151
R579 B.n361 B.n360 10.6151
R580 B.n360 B.n359 10.6151
R581 B.n359 B.n42 10.6151
R582 B.n355 B.n42 10.6151
R583 B.n355 B.n354 10.6151
R584 B.n354 B.n353 10.6151
R585 B.n353 B.n44 10.6151
R586 B.n349 B.n44 10.6151
R587 B.n349 B.n348 10.6151
R588 B.n348 B.n347 10.6151
R589 B.n347 B.n46 10.6151
R590 B.n343 B.n46 10.6151
R591 B.n343 B.n342 10.6151
R592 B.n342 B.n341 10.6151
R593 B.n341 B.n48 10.6151
R594 B.n337 B.n48 10.6151
R595 B.n337 B.n336 10.6151
R596 B.n336 B.n335 10.6151
R597 B.n335 B.n50 10.6151
R598 B.n258 B.n257 10.6151
R599 B.n259 B.n258 10.6151
R600 B.n259 B.n74 10.6151
R601 B.n263 B.n74 10.6151
R602 B.n264 B.n263 10.6151
R603 B.n265 B.n264 10.6151
R604 B.n265 B.n72 10.6151
R605 B.n269 B.n72 10.6151
R606 B.n270 B.n269 10.6151
R607 B.n271 B.n270 10.6151
R608 B.n271 B.n70 10.6151
R609 B.n275 B.n70 10.6151
R610 B.n276 B.n275 10.6151
R611 B.n277 B.n276 10.6151
R612 B.n277 B.n68 10.6151
R613 B.n281 B.n68 10.6151
R614 B.n282 B.n281 10.6151
R615 B.n283 B.n282 10.6151
R616 B.n283 B.n66 10.6151
R617 B.n287 B.n66 10.6151
R618 B.n288 B.n287 10.6151
R619 B.n289 B.n288 10.6151
R620 B.n289 B.n64 10.6151
R621 B.n293 B.n64 10.6151
R622 B.n294 B.n293 10.6151
R623 B.n295 B.n294 10.6151
R624 B.n295 B.n62 10.6151
R625 B.n299 B.n62 10.6151
R626 B.n300 B.n299 10.6151
R627 B.n301 B.n300 10.6151
R628 B.n301 B.n60 10.6151
R629 B.n305 B.n60 10.6151
R630 B.n306 B.n305 10.6151
R631 B.n307 B.n306 10.6151
R632 B.n307 B.n58 10.6151
R633 B.n311 B.n58 10.6151
R634 B.n312 B.n311 10.6151
R635 B.n313 B.n312 10.6151
R636 B.n313 B.n56 10.6151
R637 B.n317 B.n56 10.6151
R638 B.n318 B.n317 10.6151
R639 B.n319 B.n318 10.6151
R640 B.n319 B.n54 10.6151
R641 B.n323 B.n54 10.6151
R642 B.n324 B.n323 10.6151
R643 B.n325 B.n324 10.6151
R644 B.n325 B.n52 10.6151
R645 B.n329 B.n52 10.6151
R646 B.n330 B.n329 10.6151
R647 B.n331 B.n330 10.6151
R648 B.n162 B.n161 10.6151
R649 B.n163 B.n162 10.6151
R650 B.n163 B.n110 10.6151
R651 B.n167 B.n110 10.6151
R652 B.n168 B.n167 10.6151
R653 B.n169 B.n168 10.6151
R654 B.n169 B.n108 10.6151
R655 B.n173 B.n108 10.6151
R656 B.n174 B.n173 10.6151
R657 B.n175 B.n174 10.6151
R658 B.n175 B.n106 10.6151
R659 B.n179 B.n106 10.6151
R660 B.n180 B.n179 10.6151
R661 B.n181 B.n180 10.6151
R662 B.n181 B.n104 10.6151
R663 B.n185 B.n104 10.6151
R664 B.n186 B.n185 10.6151
R665 B.n187 B.n186 10.6151
R666 B.n187 B.n102 10.6151
R667 B.n191 B.n102 10.6151
R668 B.n192 B.n191 10.6151
R669 B.n193 B.n192 10.6151
R670 B.n193 B.n100 10.6151
R671 B.n197 B.n100 10.6151
R672 B.n198 B.n197 10.6151
R673 B.n199 B.n198 10.6151
R674 B.n203 B.n202 10.6151
R675 B.n204 B.n203 10.6151
R676 B.n204 B.n94 10.6151
R677 B.n208 B.n94 10.6151
R678 B.n209 B.n208 10.6151
R679 B.n210 B.n209 10.6151
R680 B.n210 B.n92 10.6151
R681 B.n214 B.n92 10.6151
R682 B.n217 B.n216 10.6151
R683 B.n217 B.n88 10.6151
R684 B.n221 B.n88 10.6151
R685 B.n222 B.n221 10.6151
R686 B.n223 B.n222 10.6151
R687 B.n223 B.n86 10.6151
R688 B.n227 B.n86 10.6151
R689 B.n228 B.n227 10.6151
R690 B.n229 B.n228 10.6151
R691 B.n229 B.n84 10.6151
R692 B.n233 B.n84 10.6151
R693 B.n234 B.n233 10.6151
R694 B.n235 B.n234 10.6151
R695 B.n235 B.n82 10.6151
R696 B.n239 B.n82 10.6151
R697 B.n240 B.n239 10.6151
R698 B.n241 B.n240 10.6151
R699 B.n241 B.n80 10.6151
R700 B.n245 B.n80 10.6151
R701 B.n246 B.n245 10.6151
R702 B.n247 B.n246 10.6151
R703 B.n247 B.n78 10.6151
R704 B.n251 B.n78 10.6151
R705 B.n252 B.n251 10.6151
R706 B.n253 B.n252 10.6151
R707 B.n253 B.n76 10.6151
R708 B.n157 B.n112 10.6151
R709 B.n157 B.n156 10.6151
R710 B.n156 B.n155 10.6151
R711 B.n155 B.n114 10.6151
R712 B.n151 B.n114 10.6151
R713 B.n151 B.n150 10.6151
R714 B.n150 B.n149 10.6151
R715 B.n149 B.n116 10.6151
R716 B.n145 B.n116 10.6151
R717 B.n145 B.n144 10.6151
R718 B.n144 B.n143 10.6151
R719 B.n143 B.n118 10.6151
R720 B.n139 B.n118 10.6151
R721 B.n139 B.n138 10.6151
R722 B.n138 B.n137 10.6151
R723 B.n137 B.n120 10.6151
R724 B.n133 B.n120 10.6151
R725 B.n133 B.n132 10.6151
R726 B.n132 B.n131 10.6151
R727 B.n131 B.n122 10.6151
R728 B.n127 B.n122 10.6151
R729 B.n127 B.n126 10.6151
R730 B.n126 B.n125 10.6151
R731 B.n125 B.n0 10.6151
R732 B.n463 B.n1 10.6151
R733 B.n463 B.n462 10.6151
R734 B.n462 B.n461 10.6151
R735 B.n461 B.n4 10.6151
R736 B.n457 B.n4 10.6151
R737 B.n457 B.n456 10.6151
R738 B.n456 B.n455 10.6151
R739 B.n455 B.n6 10.6151
R740 B.n451 B.n6 10.6151
R741 B.n451 B.n450 10.6151
R742 B.n450 B.n449 10.6151
R743 B.n449 B.n8 10.6151
R744 B.n445 B.n8 10.6151
R745 B.n445 B.n444 10.6151
R746 B.n444 B.n443 10.6151
R747 B.n443 B.n10 10.6151
R748 B.n439 B.n10 10.6151
R749 B.n439 B.n438 10.6151
R750 B.n438 B.n437 10.6151
R751 B.n437 B.n12 10.6151
R752 B.n433 B.n12 10.6151
R753 B.n433 B.n432 10.6151
R754 B.n432 B.n431 10.6151
R755 B.n431 B.n14 10.6151
R756 B.n386 B.n30 6.5566
R757 B.n374 B.n373 6.5566
R758 B.n202 B.n98 6.5566
R759 B.n215 B.n214 6.5566
R760 B.n389 B.n30 4.05904
R761 B.n373 B.n372 4.05904
R762 B.n199 B.n98 4.05904
R763 B.n216 B.n215 4.05904
R764 B.n467 B.n0 2.81026
R765 B.n467 B.n1 2.81026
R766 VP.n3 VP.t5 208.909
R767 VP.n8 VP.t2 185.7
R768 VP.n14 VP.t4 185.7
R769 VP.n6 VP.t1 185.7
R770 VP.n5 VP.n2 161.3
R771 VP.n13 VP.n0 161.3
R772 VP.n12 VP.n11 161.3
R773 VP.n10 VP.n1 161.3
R774 VP.n12 VP.t3 150.625
R775 VP.n4 VP.t0 150.625
R776 VP.n7 VP.n6 80.6037
R777 VP.n15 VP.n14 80.6037
R778 VP.n9 VP.n8 80.6037
R779 VP.n8 VP.n1 51.1515
R780 VP.n14 VP.n13 51.1515
R781 VP.n6 VP.n5 51.1515
R782 VP.n9 VP.n7 39.2931
R783 VP.n4 VP.n3 32.8731
R784 VP.n3 VP.n2 28.0424
R785 VP.n12 VP.n1 24.5923
R786 VP.n13 VP.n12 24.5923
R787 VP.n5 VP.n4 24.5923
R788 VP.n7 VP.n2 0.285035
R789 VP.n10 VP.n9 0.285035
R790 VP.n15 VP.n0 0.285035
R791 VP.n11 VP.n10 0.189894
R792 VP.n11 VP.n0 0.189894
R793 VP VP.n15 0.146778
R794 VDD1 VDD1.t0 90.8539
R795 VDD1.n1 VDD1.t3 90.7401
R796 VDD1.n1 VDD1.n0 85.4717
R797 VDD1.n3 VDD1.n2 85.2144
R798 VDD1.n3 VDD1.n1 35.0203
R799 VDD1.n2 VDD1.t5 4.64407
R800 VDD1.n2 VDD1.t4 4.64407
R801 VDD1.n0 VDD1.t2 4.64407
R802 VDD1.n0 VDD1.t1 4.64407
R803 VDD1 VDD1.n3 0.25481
C0 VN B 0.79724f
C1 VN VDD1 0.149111f
C2 VTAIL B 2.01197f
C3 VN w_n2130_n2368# 3.57078f
C4 VP B 1.24268f
C5 VDD1 VTAIL 5.8903f
C6 VDD2 B 1.35064f
C7 w_n2130_n2368# VTAIL 2.15643f
C8 VP VDD1 3.42677f
C9 VP w_n2130_n2368# 3.84203f
C10 VDD2 VDD1 0.864179f
C11 VDD2 w_n2130_n2368# 1.59951f
C12 VN VTAIL 3.32552f
C13 VN VP 4.55694f
C14 VDD1 B 1.31179f
C15 VN VDD2 3.24564f
C16 VP VTAIL 3.33986f
C17 w_n2130_n2368# B 6.23228f
C18 VDD2 VTAIL 5.93081f
C19 VDD1 w_n2130_n2368# 1.56215f
C20 VDD2 VP 0.332816f
C21 VDD2 VSUBS 1.170654f
C22 VDD1 VSUBS 1.50102f
C23 VTAIL VSUBS 0.544974f
C24 VN VSUBS 4.29817f
C25 VP VSUBS 1.549702f
C26 B VSUBS 2.753368f
C27 w_n2130_n2368# VSUBS 62.7498f
C28 VDD1.t0 VSUBS 1.14203f
C29 VDD1.t3 VSUBS 1.1413f
C30 VDD1.t2 VSUBS 0.124014f
C31 VDD1.t1 VSUBS 0.124014f
C32 VDD1.n0 VSUBS 0.854783f
C33 VDD1.n1 VSUBS 2.23329f
C34 VDD1.t5 VSUBS 0.124014f
C35 VDD1.t4 VSUBS 0.124014f
C36 VDD1.n2 VSUBS 0.853266f
C37 VDD1.n3 VSUBS 1.97476f
C38 VP.n0 VSUBS 0.07128f
C39 VP.t3 VSUBS 1.11777f
C40 VP.n1 VSUBS 0.071795f
C41 VP.n2 VSUBS 0.299402f
C42 VP.t1 VSUBS 1.20887f
C43 VP.t0 VSUBS 1.11777f
C44 VP.t5 VSUBS 1.26968f
C45 VP.n3 VSUBS 0.508903f
C46 VP.n4 VSUBS 0.528585f
C47 VP.n5 VSUBS 0.071795f
C48 VP.n6 VSUBS 0.533547f
C49 VP.n7 VSUBS 1.98693f
C50 VP.t2 VSUBS 1.20887f
C51 VP.n8 VSUBS 0.533547f
C52 VP.n9 VSUBS 2.03594f
C53 VP.n10 VSUBS 0.07128f
C54 VP.n11 VSUBS 0.053418f
C55 VP.n12 VSUBS 0.49028f
C56 VP.n13 VSUBS 0.071795f
C57 VP.t4 VSUBS 1.20887f
C58 VP.n14 VSUBS 0.533547f
C59 VP.n15 VSUBS 0.050028f
C60 B.n0 VSUBS 0.005015f
C61 B.n1 VSUBS 0.005015f
C62 B.n2 VSUBS 0.007931f
C63 B.n3 VSUBS 0.007931f
C64 B.n4 VSUBS 0.007931f
C65 B.n5 VSUBS 0.007931f
C66 B.n6 VSUBS 0.007931f
C67 B.n7 VSUBS 0.007931f
C68 B.n8 VSUBS 0.007931f
C69 B.n9 VSUBS 0.007931f
C70 B.n10 VSUBS 0.007931f
C71 B.n11 VSUBS 0.007931f
C72 B.n12 VSUBS 0.007931f
C73 B.n13 VSUBS 0.007931f
C74 B.n14 VSUBS 0.019564f
C75 B.n15 VSUBS 0.007931f
C76 B.n16 VSUBS 0.007931f
C77 B.n17 VSUBS 0.007931f
C78 B.n18 VSUBS 0.007931f
C79 B.n19 VSUBS 0.007931f
C80 B.n20 VSUBS 0.007931f
C81 B.n21 VSUBS 0.007931f
C82 B.n22 VSUBS 0.007931f
C83 B.n23 VSUBS 0.007931f
C84 B.n24 VSUBS 0.007931f
C85 B.n25 VSUBS 0.007931f
C86 B.n26 VSUBS 0.007931f
C87 B.n27 VSUBS 0.007931f
C88 B.t5 VSUBS 0.238907f
C89 B.t4 VSUBS 0.251306f
C90 B.t3 VSUBS 0.394404f
C91 B.n28 VSUBS 0.121487f
C92 B.n29 VSUBS 0.073747f
C93 B.n30 VSUBS 0.018375f
C94 B.n31 VSUBS 0.007931f
C95 B.n32 VSUBS 0.007931f
C96 B.n33 VSUBS 0.007931f
C97 B.n34 VSUBS 0.007931f
C98 B.n35 VSUBS 0.007931f
C99 B.t2 VSUBS 0.238906f
C100 B.t1 VSUBS 0.251304f
C101 B.t0 VSUBS 0.394404f
C102 B.n36 VSUBS 0.121489f
C103 B.n37 VSUBS 0.073748f
C104 B.n38 VSUBS 0.007931f
C105 B.n39 VSUBS 0.007931f
C106 B.n40 VSUBS 0.007931f
C107 B.n41 VSUBS 0.007931f
C108 B.n42 VSUBS 0.007931f
C109 B.n43 VSUBS 0.007931f
C110 B.n44 VSUBS 0.007931f
C111 B.n45 VSUBS 0.007931f
C112 B.n46 VSUBS 0.007931f
C113 B.n47 VSUBS 0.007931f
C114 B.n48 VSUBS 0.007931f
C115 B.n49 VSUBS 0.007931f
C116 B.n50 VSUBS 0.019482f
C117 B.n51 VSUBS 0.007931f
C118 B.n52 VSUBS 0.007931f
C119 B.n53 VSUBS 0.007931f
C120 B.n54 VSUBS 0.007931f
C121 B.n55 VSUBS 0.007931f
C122 B.n56 VSUBS 0.007931f
C123 B.n57 VSUBS 0.007931f
C124 B.n58 VSUBS 0.007931f
C125 B.n59 VSUBS 0.007931f
C126 B.n60 VSUBS 0.007931f
C127 B.n61 VSUBS 0.007931f
C128 B.n62 VSUBS 0.007931f
C129 B.n63 VSUBS 0.007931f
C130 B.n64 VSUBS 0.007931f
C131 B.n65 VSUBS 0.007931f
C132 B.n66 VSUBS 0.007931f
C133 B.n67 VSUBS 0.007931f
C134 B.n68 VSUBS 0.007931f
C135 B.n69 VSUBS 0.007931f
C136 B.n70 VSUBS 0.007931f
C137 B.n71 VSUBS 0.007931f
C138 B.n72 VSUBS 0.007931f
C139 B.n73 VSUBS 0.007931f
C140 B.n74 VSUBS 0.007931f
C141 B.n75 VSUBS 0.007931f
C142 B.n76 VSUBS 0.020324f
C143 B.n77 VSUBS 0.007931f
C144 B.n78 VSUBS 0.007931f
C145 B.n79 VSUBS 0.007931f
C146 B.n80 VSUBS 0.007931f
C147 B.n81 VSUBS 0.007931f
C148 B.n82 VSUBS 0.007931f
C149 B.n83 VSUBS 0.007931f
C150 B.n84 VSUBS 0.007931f
C151 B.n85 VSUBS 0.007931f
C152 B.n86 VSUBS 0.007931f
C153 B.n87 VSUBS 0.007931f
C154 B.n88 VSUBS 0.007931f
C155 B.n89 VSUBS 0.007931f
C156 B.t7 VSUBS 0.238906f
C157 B.t8 VSUBS 0.251304f
C158 B.t6 VSUBS 0.394404f
C159 B.n90 VSUBS 0.121489f
C160 B.n91 VSUBS 0.073748f
C161 B.n92 VSUBS 0.007931f
C162 B.n93 VSUBS 0.007931f
C163 B.n94 VSUBS 0.007931f
C164 B.n95 VSUBS 0.007931f
C165 B.t10 VSUBS 0.238907f
C166 B.t11 VSUBS 0.251306f
C167 B.t9 VSUBS 0.394404f
C168 B.n96 VSUBS 0.121487f
C169 B.n97 VSUBS 0.073747f
C170 B.n98 VSUBS 0.018375f
C171 B.n99 VSUBS 0.007931f
C172 B.n100 VSUBS 0.007931f
C173 B.n101 VSUBS 0.007931f
C174 B.n102 VSUBS 0.007931f
C175 B.n103 VSUBS 0.007931f
C176 B.n104 VSUBS 0.007931f
C177 B.n105 VSUBS 0.007931f
C178 B.n106 VSUBS 0.007931f
C179 B.n107 VSUBS 0.007931f
C180 B.n108 VSUBS 0.007931f
C181 B.n109 VSUBS 0.007931f
C182 B.n110 VSUBS 0.007931f
C183 B.n111 VSUBS 0.007931f
C184 B.n112 VSUBS 0.019564f
C185 B.n113 VSUBS 0.007931f
C186 B.n114 VSUBS 0.007931f
C187 B.n115 VSUBS 0.007931f
C188 B.n116 VSUBS 0.007931f
C189 B.n117 VSUBS 0.007931f
C190 B.n118 VSUBS 0.007931f
C191 B.n119 VSUBS 0.007931f
C192 B.n120 VSUBS 0.007931f
C193 B.n121 VSUBS 0.007931f
C194 B.n122 VSUBS 0.007931f
C195 B.n123 VSUBS 0.007931f
C196 B.n124 VSUBS 0.007931f
C197 B.n125 VSUBS 0.007931f
C198 B.n126 VSUBS 0.007931f
C199 B.n127 VSUBS 0.007931f
C200 B.n128 VSUBS 0.007931f
C201 B.n129 VSUBS 0.007931f
C202 B.n130 VSUBS 0.007931f
C203 B.n131 VSUBS 0.007931f
C204 B.n132 VSUBS 0.007931f
C205 B.n133 VSUBS 0.007931f
C206 B.n134 VSUBS 0.007931f
C207 B.n135 VSUBS 0.007931f
C208 B.n136 VSUBS 0.007931f
C209 B.n137 VSUBS 0.007931f
C210 B.n138 VSUBS 0.007931f
C211 B.n139 VSUBS 0.007931f
C212 B.n140 VSUBS 0.007931f
C213 B.n141 VSUBS 0.007931f
C214 B.n142 VSUBS 0.007931f
C215 B.n143 VSUBS 0.007931f
C216 B.n144 VSUBS 0.007931f
C217 B.n145 VSUBS 0.007931f
C218 B.n146 VSUBS 0.007931f
C219 B.n147 VSUBS 0.007931f
C220 B.n148 VSUBS 0.007931f
C221 B.n149 VSUBS 0.007931f
C222 B.n150 VSUBS 0.007931f
C223 B.n151 VSUBS 0.007931f
C224 B.n152 VSUBS 0.007931f
C225 B.n153 VSUBS 0.007931f
C226 B.n154 VSUBS 0.007931f
C227 B.n155 VSUBS 0.007931f
C228 B.n156 VSUBS 0.007931f
C229 B.n157 VSUBS 0.007931f
C230 B.n158 VSUBS 0.007931f
C231 B.n159 VSUBS 0.019564f
C232 B.n160 VSUBS 0.020324f
C233 B.n161 VSUBS 0.020324f
C234 B.n162 VSUBS 0.007931f
C235 B.n163 VSUBS 0.007931f
C236 B.n164 VSUBS 0.007931f
C237 B.n165 VSUBS 0.007931f
C238 B.n166 VSUBS 0.007931f
C239 B.n167 VSUBS 0.007931f
C240 B.n168 VSUBS 0.007931f
C241 B.n169 VSUBS 0.007931f
C242 B.n170 VSUBS 0.007931f
C243 B.n171 VSUBS 0.007931f
C244 B.n172 VSUBS 0.007931f
C245 B.n173 VSUBS 0.007931f
C246 B.n174 VSUBS 0.007931f
C247 B.n175 VSUBS 0.007931f
C248 B.n176 VSUBS 0.007931f
C249 B.n177 VSUBS 0.007931f
C250 B.n178 VSUBS 0.007931f
C251 B.n179 VSUBS 0.007931f
C252 B.n180 VSUBS 0.007931f
C253 B.n181 VSUBS 0.007931f
C254 B.n182 VSUBS 0.007931f
C255 B.n183 VSUBS 0.007931f
C256 B.n184 VSUBS 0.007931f
C257 B.n185 VSUBS 0.007931f
C258 B.n186 VSUBS 0.007931f
C259 B.n187 VSUBS 0.007931f
C260 B.n188 VSUBS 0.007931f
C261 B.n189 VSUBS 0.007931f
C262 B.n190 VSUBS 0.007931f
C263 B.n191 VSUBS 0.007931f
C264 B.n192 VSUBS 0.007931f
C265 B.n193 VSUBS 0.007931f
C266 B.n194 VSUBS 0.007931f
C267 B.n195 VSUBS 0.007931f
C268 B.n196 VSUBS 0.007931f
C269 B.n197 VSUBS 0.007931f
C270 B.n198 VSUBS 0.007931f
C271 B.n199 VSUBS 0.005482f
C272 B.n200 VSUBS 0.007931f
C273 B.n201 VSUBS 0.007931f
C274 B.n202 VSUBS 0.006415f
C275 B.n203 VSUBS 0.007931f
C276 B.n204 VSUBS 0.007931f
C277 B.n205 VSUBS 0.007931f
C278 B.n206 VSUBS 0.007931f
C279 B.n207 VSUBS 0.007931f
C280 B.n208 VSUBS 0.007931f
C281 B.n209 VSUBS 0.007931f
C282 B.n210 VSUBS 0.007931f
C283 B.n211 VSUBS 0.007931f
C284 B.n212 VSUBS 0.007931f
C285 B.n213 VSUBS 0.007931f
C286 B.n214 VSUBS 0.006415f
C287 B.n215 VSUBS 0.018375f
C288 B.n216 VSUBS 0.005482f
C289 B.n217 VSUBS 0.007931f
C290 B.n218 VSUBS 0.007931f
C291 B.n219 VSUBS 0.007931f
C292 B.n220 VSUBS 0.007931f
C293 B.n221 VSUBS 0.007931f
C294 B.n222 VSUBS 0.007931f
C295 B.n223 VSUBS 0.007931f
C296 B.n224 VSUBS 0.007931f
C297 B.n225 VSUBS 0.007931f
C298 B.n226 VSUBS 0.007931f
C299 B.n227 VSUBS 0.007931f
C300 B.n228 VSUBS 0.007931f
C301 B.n229 VSUBS 0.007931f
C302 B.n230 VSUBS 0.007931f
C303 B.n231 VSUBS 0.007931f
C304 B.n232 VSUBS 0.007931f
C305 B.n233 VSUBS 0.007931f
C306 B.n234 VSUBS 0.007931f
C307 B.n235 VSUBS 0.007931f
C308 B.n236 VSUBS 0.007931f
C309 B.n237 VSUBS 0.007931f
C310 B.n238 VSUBS 0.007931f
C311 B.n239 VSUBS 0.007931f
C312 B.n240 VSUBS 0.007931f
C313 B.n241 VSUBS 0.007931f
C314 B.n242 VSUBS 0.007931f
C315 B.n243 VSUBS 0.007931f
C316 B.n244 VSUBS 0.007931f
C317 B.n245 VSUBS 0.007931f
C318 B.n246 VSUBS 0.007931f
C319 B.n247 VSUBS 0.007931f
C320 B.n248 VSUBS 0.007931f
C321 B.n249 VSUBS 0.007931f
C322 B.n250 VSUBS 0.007931f
C323 B.n251 VSUBS 0.007931f
C324 B.n252 VSUBS 0.007931f
C325 B.n253 VSUBS 0.007931f
C326 B.n254 VSUBS 0.007931f
C327 B.n255 VSUBS 0.020324f
C328 B.n256 VSUBS 0.019564f
C329 B.n257 VSUBS 0.019564f
C330 B.n258 VSUBS 0.007931f
C331 B.n259 VSUBS 0.007931f
C332 B.n260 VSUBS 0.007931f
C333 B.n261 VSUBS 0.007931f
C334 B.n262 VSUBS 0.007931f
C335 B.n263 VSUBS 0.007931f
C336 B.n264 VSUBS 0.007931f
C337 B.n265 VSUBS 0.007931f
C338 B.n266 VSUBS 0.007931f
C339 B.n267 VSUBS 0.007931f
C340 B.n268 VSUBS 0.007931f
C341 B.n269 VSUBS 0.007931f
C342 B.n270 VSUBS 0.007931f
C343 B.n271 VSUBS 0.007931f
C344 B.n272 VSUBS 0.007931f
C345 B.n273 VSUBS 0.007931f
C346 B.n274 VSUBS 0.007931f
C347 B.n275 VSUBS 0.007931f
C348 B.n276 VSUBS 0.007931f
C349 B.n277 VSUBS 0.007931f
C350 B.n278 VSUBS 0.007931f
C351 B.n279 VSUBS 0.007931f
C352 B.n280 VSUBS 0.007931f
C353 B.n281 VSUBS 0.007931f
C354 B.n282 VSUBS 0.007931f
C355 B.n283 VSUBS 0.007931f
C356 B.n284 VSUBS 0.007931f
C357 B.n285 VSUBS 0.007931f
C358 B.n286 VSUBS 0.007931f
C359 B.n287 VSUBS 0.007931f
C360 B.n288 VSUBS 0.007931f
C361 B.n289 VSUBS 0.007931f
C362 B.n290 VSUBS 0.007931f
C363 B.n291 VSUBS 0.007931f
C364 B.n292 VSUBS 0.007931f
C365 B.n293 VSUBS 0.007931f
C366 B.n294 VSUBS 0.007931f
C367 B.n295 VSUBS 0.007931f
C368 B.n296 VSUBS 0.007931f
C369 B.n297 VSUBS 0.007931f
C370 B.n298 VSUBS 0.007931f
C371 B.n299 VSUBS 0.007931f
C372 B.n300 VSUBS 0.007931f
C373 B.n301 VSUBS 0.007931f
C374 B.n302 VSUBS 0.007931f
C375 B.n303 VSUBS 0.007931f
C376 B.n304 VSUBS 0.007931f
C377 B.n305 VSUBS 0.007931f
C378 B.n306 VSUBS 0.007931f
C379 B.n307 VSUBS 0.007931f
C380 B.n308 VSUBS 0.007931f
C381 B.n309 VSUBS 0.007931f
C382 B.n310 VSUBS 0.007931f
C383 B.n311 VSUBS 0.007931f
C384 B.n312 VSUBS 0.007931f
C385 B.n313 VSUBS 0.007931f
C386 B.n314 VSUBS 0.007931f
C387 B.n315 VSUBS 0.007931f
C388 B.n316 VSUBS 0.007931f
C389 B.n317 VSUBS 0.007931f
C390 B.n318 VSUBS 0.007931f
C391 B.n319 VSUBS 0.007931f
C392 B.n320 VSUBS 0.007931f
C393 B.n321 VSUBS 0.007931f
C394 B.n322 VSUBS 0.007931f
C395 B.n323 VSUBS 0.007931f
C396 B.n324 VSUBS 0.007931f
C397 B.n325 VSUBS 0.007931f
C398 B.n326 VSUBS 0.007931f
C399 B.n327 VSUBS 0.007931f
C400 B.n328 VSUBS 0.007931f
C401 B.n329 VSUBS 0.007931f
C402 B.n330 VSUBS 0.007931f
C403 B.n331 VSUBS 0.020406f
C404 B.n332 VSUBS 0.019564f
C405 B.n333 VSUBS 0.020324f
C406 B.n334 VSUBS 0.007931f
C407 B.n335 VSUBS 0.007931f
C408 B.n336 VSUBS 0.007931f
C409 B.n337 VSUBS 0.007931f
C410 B.n338 VSUBS 0.007931f
C411 B.n339 VSUBS 0.007931f
C412 B.n340 VSUBS 0.007931f
C413 B.n341 VSUBS 0.007931f
C414 B.n342 VSUBS 0.007931f
C415 B.n343 VSUBS 0.007931f
C416 B.n344 VSUBS 0.007931f
C417 B.n345 VSUBS 0.007931f
C418 B.n346 VSUBS 0.007931f
C419 B.n347 VSUBS 0.007931f
C420 B.n348 VSUBS 0.007931f
C421 B.n349 VSUBS 0.007931f
C422 B.n350 VSUBS 0.007931f
C423 B.n351 VSUBS 0.007931f
C424 B.n352 VSUBS 0.007931f
C425 B.n353 VSUBS 0.007931f
C426 B.n354 VSUBS 0.007931f
C427 B.n355 VSUBS 0.007931f
C428 B.n356 VSUBS 0.007931f
C429 B.n357 VSUBS 0.007931f
C430 B.n358 VSUBS 0.007931f
C431 B.n359 VSUBS 0.007931f
C432 B.n360 VSUBS 0.007931f
C433 B.n361 VSUBS 0.007931f
C434 B.n362 VSUBS 0.007931f
C435 B.n363 VSUBS 0.007931f
C436 B.n364 VSUBS 0.007931f
C437 B.n365 VSUBS 0.007931f
C438 B.n366 VSUBS 0.007931f
C439 B.n367 VSUBS 0.007931f
C440 B.n368 VSUBS 0.007931f
C441 B.n369 VSUBS 0.007931f
C442 B.n370 VSUBS 0.007931f
C443 B.n371 VSUBS 0.007931f
C444 B.n372 VSUBS 0.005482f
C445 B.n373 VSUBS 0.018375f
C446 B.n374 VSUBS 0.006415f
C447 B.n375 VSUBS 0.007931f
C448 B.n376 VSUBS 0.007931f
C449 B.n377 VSUBS 0.007931f
C450 B.n378 VSUBS 0.007931f
C451 B.n379 VSUBS 0.007931f
C452 B.n380 VSUBS 0.007931f
C453 B.n381 VSUBS 0.007931f
C454 B.n382 VSUBS 0.007931f
C455 B.n383 VSUBS 0.007931f
C456 B.n384 VSUBS 0.007931f
C457 B.n385 VSUBS 0.007931f
C458 B.n386 VSUBS 0.006415f
C459 B.n387 VSUBS 0.007931f
C460 B.n388 VSUBS 0.007931f
C461 B.n389 VSUBS 0.005482f
C462 B.n390 VSUBS 0.007931f
C463 B.n391 VSUBS 0.007931f
C464 B.n392 VSUBS 0.007931f
C465 B.n393 VSUBS 0.007931f
C466 B.n394 VSUBS 0.007931f
C467 B.n395 VSUBS 0.007931f
C468 B.n396 VSUBS 0.007931f
C469 B.n397 VSUBS 0.007931f
C470 B.n398 VSUBS 0.007931f
C471 B.n399 VSUBS 0.007931f
C472 B.n400 VSUBS 0.007931f
C473 B.n401 VSUBS 0.007931f
C474 B.n402 VSUBS 0.007931f
C475 B.n403 VSUBS 0.007931f
C476 B.n404 VSUBS 0.007931f
C477 B.n405 VSUBS 0.007931f
C478 B.n406 VSUBS 0.007931f
C479 B.n407 VSUBS 0.007931f
C480 B.n408 VSUBS 0.007931f
C481 B.n409 VSUBS 0.007931f
C482 B.n410 VSUBS 0.007931f
C483 B.n411 VSUBS 0.007931f
C484 B.n412 VSUBS 0.007931f
C485 B.n413 VSUBS 0.007931f
C486 B.n414 VSUBS 0.007931f
C487 B.n415 VSUBS 0.007931f
C488 B.n416 VSUBS 0.007931f
C489 B.n417 VSUBS 0.007931f
C490 B.n418 VSUBS 0.007931f
C491 B.n419 VSUBS 0.007931f
C492 B.n420 VSUBS 0.007931f
C493 B.n421 VSUBS 0.007931f
C494 B.n422 VSUBS 0.007931f
C495 B.n423 VSUBS 0.007931f
C496 B.n424 VSUBS 0.007931f
C497 B.n425 VSUBS 0.007931f
C498 B.n426 VSUBS 0.007931f
C499 B.n427 VSUBS 0.020324f
C500 B.n428 VSUBS 0.020324f
C501 B.n429 VSUBS 0.019564f
C502 B.n430 VSUBS 0.007931f
C503 B.n431 VSUBS 0.007931f
C504 B.n432 VSUBS 0.007931f
C505 B.n433 VSUBS 0.007931f
C506 B.n434 VSUBS 0.007931f
C507 B.n435 VSUBS 0.007931f
C508 B.n436 VSUBS 0.007931f
C509 B.n437 VSUBS 0.007931f
C510 B.n438 VSUBS 0.007931f
C511 B.n439 VSUBS 0.007931f
C512 B.n440 VSUBS 0.007931f
C513 B.n441 VSUBS 0.007931f
C514 B.n442 VSUBS 0.007931f
C515 B.n443 VSUBS 0.007931f
C516 B.n444 VSUBS 0.007931f
C517 B.n445 VSUBS 0.007931f
C518 B.n446 VSUBS 0.007931f
C519 B.n447 VSUBS 0.007931f
C520 B.n448 VSUBS 0.007931f
C521 B.n449 VSUBS 0.007931f
C522 B.n450 VSUBS 0.007931f
C523 B.n451 VSUBS 0.007931f
C524 B.n452 VSUBS 0.007931f
C525 B.n453 VSUBS 0.007931f
C526 B.n454 VSUBS 0.007931f
C527 B.n455 VSUBS 0.007931f
C528 B.n456 VSUBS 0.007931f
C529 B.n457 VSUBS 0.007931f
C530 B.n458 VSUBS 0.007931f
C531 B.n459 VSUBS 0.007931f
C532 B.n460 VSUBS 0.007931f
C533 B.n461 VSUBS 0.007931f
C534 B.n462 VSUBS 0.007931f
C535 B.n463 VSUBS 0.007931f
C536 B.n464 VSUBS 0.007931f
C537 B.n465 VSUBS 0.007931f
C538 B.n466 VSUBS 0.007931f
C539 B.n467 VSUBS 0.017958f
C540 VDD2.t2 VSUBS 1.12679f
C541 VDD2.t4 VSUBS 0.122438f
C542 VDD2.t5 VSUBS 0.122438f
C543 VDD2.n0 VSUBS 0.843915f
C544 VDD2.n1 VSUBS 2.13025f
C545 VDD2.t3 VSUBS 1.12188f
C546 VDD2.n2 VSUBS 1.96073f
C547 VDD2.t0 VSUBS 0.122438f
C548 VDD2.t1 VSUBS 0.122438f
C549 VDD2.n3 VSUBS 0.84389f
C550 VTAIL.t11 VSUBS 0.16945f
C551 VTAIL.t9 VSUBS 0.16945f
C552 VTAIL.n0 VSUBS 1.03968f
C553 VTAIL.n1 VSUBS 0.753627f
C554 VTAIL.t2 VSUBS 1.41727f
C555 VTAIL.n2 VSUBS 0.924968f
C556 VTAIL.t4 VSUBS 0.16945f
C557 VTAIL.t5 VSUBS 0.16945f
C558 VTAIL.n3 VSUBS 1.03968f
C559 VTAIL.n4 VSUBS 1.99087f
C560 VTAIL.t8 VSUBS 0.16945f
C561 VTAIL.t7 VSUBS 0.16945f
C562 VTAIL.n5 VSUBS 1.03968f
C563 VTAIL.n6 VSUBS 1.99087f
C564 VTAIL.t6 VSUBS 1.41728f
C565 VTAIL.n7 VSUBS 0.924961f
C566 VTAIL.t3 VSUBS 0.16945f
C567 VTAIL.t0 VSUBS 0.16945f
C568 VTAIL.n8 VSUBS 1.03968f
C569 VTAIL.n9 VSUBS 0.840416f
C570 VTAIL.t1 VSUBS 1.41727f
C571 VTAIL.n10 VSUBS 1.95204f
C572 VTAIL.t10 VSUBS 1.41727f
C573 VTAIL.n11 VSUBS 1.91545f
C574 VN.n0 VSUBS 0.290029f
C575 VN.t1 VSUBS 1.08278f
C576 VN.t3 VSUBS 1.22993f
C577 VN.n1 VSUBS 0.492971f
C578 VN.n2 VSUBS 0.512036f
C579 VN.n3 VSUBS 0.069548f
C580 VN.t0 VSUBS 1.17103f
C581 VN.n4 VSUBS 0.516843f
C582 VN.n5 VSUBS 0.048462f
C583 VN.n6 VSUBS 0.290029f
C584 VN.t5 VSUBS 1.08278f
C585 VN.t4 VSUBS 1.22993f
C586 VN.n7 VSUBS 0.492971f
C587 VN.n8 VSUBS 0.512036f
C588 VN.n9 VSUBS 0.069548f
C589 VN.t2 VSUBS 1.17103f
C590 VN.n10 VSUBS 0.516843f
C591 VN.n11 VSUBS 1.95411f
.ends

