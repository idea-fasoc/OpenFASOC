* NGSPICE file created from diff_pair_sample_1297.ext - technology: sky130A

.subckt diff_pair_sample_1297 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=1.63
X1 VDD2.t4 VN.t1 VTAIL.t11 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=1.63
X2 B.t11 B.t9 B.t10 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=1.63
X3 VTAIL.t0 VP.t0 VDD1.t5 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=2.57565 ps=15.94 w=15.61 l=1.63
X4 VTAIL.t9 VN.t2 VDD2.t3 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=2.57565 ps=15.94 w=15.61 l=1.63
X5 VDD1.t4 VP.t1 VTAIL.t5 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=1.63
X6 VDD2.t2 VN.t3 VTAIL.t7 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=1.63
X7 VDD2.t1 VN.t4 VTAIL.t10 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=1.63
X8 B.t8 B.t6 B.t7 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=1.63
X9 B.t5 B.t3 B.t4 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=1.63
X10 VTAIL.t3 VP.t2 VDD1.t3 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=2.57565 ps=15.94 w=15.61 l=1.63
X11 VDD1.t2 VP.t3 VTAIL.t2 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=1.63
X12 VTAIL.t8 VN.t5 VDD2.t0 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=2.57565 ps=15.94 w=15.61 l=1.63
X13 VDD1.t1 VP.t4 VTAIL.t1 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=1.63
X14 VDD1.t0 VP.t5 VTAIL.t4 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=1.63
X15 B.t2 B.t0 B.t1 w_n2538_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=1.63
R0 VN.n2 VN.t0 264.673
R1 VN.n14 VN.t3 264.673
R2 VN.n3 VN.t2 230.798
R3 VN.n10 VN.t4 230.798
R4 VN.n15 VN.t5 230.798
R5 VN.n22 VN.t1 230.798
R6 VN.n11 VN.n10 175.492
R7 VN.n23 VN.n22 175.492
R8 VN.n21 VN.n12 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n13 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n9 VN.n0 161.3
R13 VN.n8 VN.n7 161.3
R14 VN.n6 VN.n1 161.3
R15 VN.n5 VN.n4 161.3
R16 VN.n8 VN.n1 56.5193
R17 VN.n20 VN.n13 56.5193
R18 VN.n3 VN.n2 54.1657
R19 VN.n15 VN.n14 54.1657
R20 VN VN.n23 47.9494
R21 VN.n4 VN.n1 24.4675
R22 VN.n9 VN.n8 24.4675
R23 VN.n16 VN.n13 24.4675
R24 VN.n21 VN.n20 24.4675
R25 VN.n17 VN.n14 17.7577
R26 VN.n5 VN.n2 17.7577
R27 VN.n4 VN.n3 12.234
R28 VN.n16 VN.n15 12.234
R29 VN.n10 VN.n9 10.2766
R30 VN.n22 VN.n21 10.2766
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n346 VTAIL.n266 756.745
R41 VTAIL.n82 VTAIL.n2 756.745
R42 VTAIL.n260 VTAIL.n180 756.745
R43 VTAIL.n172 VTAIL.n92 756.745
R44 VTAIL.n295 VTAIL.n294 585
R45 VTAIL.n297 VTAIL.n296 585
R46 VTAIL.n290 VTAIL.n289 585
R47 VTAIL.n303 VTAIL.n302 585
R48 VTAIL.n305 VTAIL.n304 585
R49 VTAIL.n286 VTAIL.n285 585
R50 VTAIL.n312 VTAIL.n311 585
R51 VTAIL.n313 VTAIL.n284 585
R52 VTAIL.n315 VTAIL.n314 585
R53 VTAIL.n282 VTAIL.n281 585
R54 VTAIL.n321 VTAIL.n320 585
R55 VTAIL.n323 VTAIL.n322 585
R56 VTAIL.n278 VTAIL.n277 585
R57 VTAIL.n329 VTAIL.n328 585
R58 VTAIL.n331 VTAIL.n330 585
R59 VTAIL.n274 VTAIL.n273 585
R60 VTAIL.n337 VTAIL.n336 585
R61 VTAIL.n339 VTAIL.n338 585
R62 VTAIL.n270 VTAIL.n269 585
R63 VTAIL.n345 VTAIL.n344 585
R64 VTAIL.n347 VTAIL.n346 585
R65 VTAIL.n31 VTAIL.n30 585
R66 VTAIL.n33 VTAIL.n32 585
R67 VTAIL.n26 VTAIL.n25 585
R68 VTAIL.n39 VTAIL.n38 585
R69 VTAIL.n41 VTAIL.n40 585
R70 VTAIL.n22 VTAIL.n21 585
R71 VTAIL.n48 VTAIL.n47 585
R72 VTAIL.n49 VTAIL.n20 585
R73 VTAIL.n51 VTAIL.n50 585
R74 VTAIL.n18 VTAIL.n17 585
R75 VTAIL.n57 VTAIL.n56 585
R76 VTAIL.n59 VTAIL.n58 585
R77 VTAIL.n14 VTAIL.n13 585
R78 VTAIL.n65 VTAIL.n64 585
R79 VTAIL.n67 VTAIL.n66 585
R80 VTAIL.n10 VTAIL.n9 585
R81 VTAIL.n73 VTAIL.n72 585
R82 VTAIL.n75 VTAIL.n74 585
R83 VTAIL.n6 VTAIL.n5 585
R84 VTAIL.n81 VTAIL.n80 585
R85 VTAIL.n83 VTAIL.n82 585
R86 VTAIL.n261 VTAIL.n260 585
R87 VTAIL.n259 VTAIL.n258 585
R88 VTAIL.n184 VTAIL.n183 585
R89 VTAIL.n253 VTAIL.n252 585
R90 VTAIL.n251 VTAIL.n250 585
R91 VTAIL.n188 VTAIL.n187 585
R92 VTAIL.n245 VTAIL.n244 585
R93 VTAIL.n243 VTAIL.n242 585
R94 VTAIL.n192 VTAIL.n191 585
R95 VTAIL.n237 VTAIL.n236 585
R96 VTAIL.n235 VTAIL.n234 585
R97 VTAIL.n196 VTAIL.n195 585
R98 VTAIL.n200 VTAIL.n198 585
R99 VTAIL.n229 VTAIL.n228 585
R100 VTAIL.n227 VTAIL.n226 585
R101 VTAIL.n202 VTAIL.n201 585
R102 VTAIL.n221 VTAIL.n220 585
R103 VTAIL.n219 VTAIL.n218 585
R104 VTAIL.n206 VTAIL.n205 585
R105 VTAIL.n213 VTAIL.n212 585
R106 VTAIL.n211 VTAIL.n210 585
R107 VTAIL.n173 VTAIL.n172 585
R108 VTAIL.n171 VTAIL.n170 585
R109 VTAIL.n96 VTAIL.n95 585
R110 VTAIL.n165 VTAIL.n164 585
R111 VTAIL.n163 VTAIL.n162 585
R112 VTAIL.n100 VTAIL.n99 585
R113 VTAIL.n157 VTAIL.n156 585
R114 VTAIL.n155 VTAIL.n154 585
R115 VTAIL.n104 VTAIL.n103 585
R116 VTAIL.n149 VTAIL.n148 585
R117 VTAIL.n147 VTAIL.n146 585
R118 VTAIL.n108 VTAIL.n107 585
R119 VTAIL.n112 VTAIL.n110 585
R120 VTAIL.n141 VTAIL.n140 585
R121 VTAIL.n139 VTAIL.n138 585
R122 VTAIL.n114 VTAIL.n113 585
R123 VTAIL.n133 VTAIL.n132 585
R124 VTAIL.n131 VTAIL.n130 585
R125 VTAIL.n118 VTAIL.n117 585
R126 VTAIL.n125 VTAIL.n124 585
R127 VTAIL.n123 VTAIL.n122 585
R128 VTAIL.n293 VTAIL.t10 329.036
R129 VTAIL.n29 VTAIL.t5 329.036
R130 VTAIL.n209 VTAIL.t2 329.036
R131 VTAIL.n121 VTAIL.t7 329.036
R132 VTAIL.n296 VTAIL.n295 171.744
R133 VTAIL.n296 VTAIL.n289 171.744
R134 VTAIL.n303 VTAIL.n289 171.744
R135 VTAIL.n304 VTAIL.n303 171.744
R136 VTAIL.n304 VTAIL.n285 171.744
R137 VTAIL.n312 VTAIL.n285 171.744
R138 VTAIL.n313 VTAIL.n312 171.744
R139 VTAIL.n314 VTAIL.n313 171.744
R140 VTAIL.n314 VTAIL.n281 171.744
R141 VTAIL.n321 VTAIL.n281 171.744
R142 VTAIL.n322 VTAIL.n321 171.744
R143 VTAIL.n322 VTAIL.n277 171.744
R144 VTAIL.n329 VTAIL.n277 171.744
R145 VTAIL.n330 VTAIL.n329 171.744
R146 VTAIL.n330 VTAIL.n273 171.744
R147 VTAIL.n337 VTAIL.n273 171.744
R148 VTAIL.n338 VTAIL.n337 171.744
R149 VTAIL.n338 VTAIL.n269 171.744
R150 VTAIL.n345 VTAIL.n269 171.744
R151 VTAIL.n346 VTAIL.n345 171.744
R152 VTAIL.n32 VTAIL.n31 171.744
R153 VTAIL.n32 VTAIL.n25 171.744
R154 VTAIL.n39 VTAIL.n25 171.744
R155 VTAIL.n40 VTAIL.n39 171.744
R156 VTAIL.n40 VTAIL.n21 171.744
R157 VTAIL.n48 VTAIL.n21 171.744
R158 VTAIL.n49 VTAIL.n48 171.744
R159 VTAIL.n50 VTAIL.n49 171.744
R160 VTAIL.n50 VTAIL.n17 171.744
R161 VTAIL.n57 VTAIL.n17 171.744
R162 VTAIL.n58 VTAIL.n57 171.744
R163 VTAIL.n58 VTAIL.n13 171.744
R164 VTAIL.n65 VTAIL.n13 171.744
R165 VTAIL.n66 VTAIL.n65 171.744
R166 VTAIL.n66 VTAIL.n9 171.744
R167 VTAIL.n73 VTAIL.n9 171.744
R168 VTAIL.n74 VTAIL.n73 171.744
R169 VTAIL.n74 VTAIL.n5 171.744
R170 VTAIL.n81 VTAIL.n5 171.744
R171 VTAIL.n82 VTAIL.n81 171.744
R172 VTAIL.n260 VTAIL.n259 171.744
R173 VTAIL.n259 VTAIL.n183 171.744
R174 VTAIL.n252 VTAIL.n183 171.744
R175 VTAIL.n252 VTAIL.n251 171.744
R176 VTAIL.n251 VTAIL.n187 171.744
R177 VTAIL.n244 VTAIL.n187 171.744
R178 VTAIL.n244 VTAIL.n243 171.744
R179 VTAIL.n243 VTAIL.n191 171.744
R180 VTAIL.n236 VTAIL.n191 171.744
R181 VTAIL.n236 VTAIL.n235 171.744
R182 VTAIL.n235 VTAIL.n195 171.744
R183 VTAIL.n200 VTAIL.n195 171.744
R184 VTAIL.n228 VTAIL.n200 171.744
R185 VTAIL.n228 VTAIL.n227 171.744
R186 VTAIL.n227 VTAIL.n201 171.744
R187 VTAIL.n220 VTAIL.n201 171.744
R188 VTAIL.n220 VTAIL.n219 171.744
R189 VTAIL.n219 VTAIL.n205 171.744
R190 VTAIL.n212 VTAIL.n205 171.744
R191 VTAIL.n212 VTAIL.n211 171.744
R192 VTAIL.n172 VTAIL.n171 171.744
R193 VTAIL.n171 VTAIL.n95 171.744
R194 VTAIL.n164 VTAIL.n95 171.744
R195 VTAIL.n164 VTAIL.n163 171.744
R196 VTAIL.n163 VTAIL.n99 171.744
R197 VTAIL.n156 VTAIL.n99 171.744
R198 VTAIL.n156 VTAIL.n155 171.744
R199 VTAIL.n155 VTAIL.n103 171.744
R200 VTAIL.n148 VTAIL.n103 171.744
R201 VTAIL.n148 VTAIL.n147 171.744
R202 VTAIL.n147 VTAIL.n107 171.744
R203 VTAIL.n112 VTAIL.n107 171.744
R204 VTAIL.n140 VTAIL.n112 171.744
R205 VTAIL.n140 VTAIL.n139 171.744
R206 VTAIL.n139 VTAIL.n113 171.744
R207 VTAIL.n132 VTAIL.n113 171.744
R208 VTAIL.n132 VTAIL.n131 171.744
R209 VTAIL.n131 VTAIL.n117 171.744
R210 VTAIL.n124 VTAIL.n117 171.744
R211 VTAIL.n124 VTAIL.n123 171.744
R212 VTAIL.n295 VTAIL.t10 85.8723
R213 VTAIL.n31 VTAIL.t5 85.8723
R214 VTAIL.n211 VTAIL.t2 85.8723
R215 VTAIL.n123 VTAIL.t7 85.8723
R216 VTAIL.n1 VTAIL.n0 51.727
R217 VTAIL.n89 VTAIL.n88 51.727
R218 VTAIL.n179 VTAIL.n178 51.727
R219 VTAIL.n91 VTAIL.n90 51.727
R220 VTAIL.n351 VTAIL.n350 30.052
R221 VTAIL.n87 VTAIL.n86 30.052
R222 VTAIL.n265 VTAIL.n264 30.052
R223 VTAIL.n177 VTAIL.n176 30.052
R224 VTAIL.n91 VTAIL.n89 29.2031
R225 VTAIL.n351 VTAIL.n265 27.5134
R226 VTAIL.n315 VTAIL.n282 13.1884
R227 VTAIL.n51 VTAIL.n18 13.1884
R228 VTAIL.n198 VTAIL.n196 13.1884
R229 VTAIL.n110 VTAIL.n108 13.1884
R230 VTAIL.n316 VTAIL.n284 12.8005
R231 VTAIL.n320 VTAIL.n319 12.8005
R232 VTAIL.n52 VTAIL.n20 12.8005
R233 VTAIL.n56 VTAIL.n55 12.8005
R234 VTAIL.n234 VTAIL.n233 12.8005
R235 VTAIL.n230 VTAIL.n229 12.8005
R236 VTAIL.n146 VTAIL.n145 12.8005
R237 VTAIL.n142 VTAIL.n141 12.8005
R238 VTAIL.n311 VTAIL.n310 12.0247
R239 VTAIL.n323 VTAIL.n280 12.0247
R240 VTAIL.n47 VTAIL.n46 12.0247
R241 VTAIL.n59 VTAIL.n16 12.0247
R242 VTAIL.n237 VTAIL.n194 12.0247
R243 VTAIL.n226 VTAIL.n199 12.0247
R244 VTAIL.n149 VTAIL.n106 12.0247
R245 VTAIL.n138 VTAIL.n111 12.0247
R246 VTAIL.n309 VTAIL.n286 11.249
R247 VTAIL.n324 VTAIL.n278 11.249
R248 VTAIL.n45 VTAIL.n22 11.249
R249 VTAIL.n60 VTAIL.n14 11.249
R250 VTAIL.n238 VTAIL.n192 11.249
R251 VTAIL.n225 VTAIL.n202 11.249
R252 VTAIL.n150 VTAIL.n104 11.249
R253 VTAIL.n137 VTAIL.n114 11.249
R254 VTAIL.n294 VTAIL.n293 10.7239
R255 VTAIL.n30 VTAIL.n29 10.7239
R256 VTAIL.n210 VTAIL.n209 10.7239
R257 VTAIL.n122 VTAIL.n121 10.7239
R258 VTAIL.n306 VTAIL.n305 10.4732
R259 VTAIL.n328 VTAIL.n327 10.4732
R260 VTAIL.n42 VTAIL.n41 10.4732
R261 VTAIL.n64 VTAIL.n63 10.4732
R262 VTAIL.n242 VTAIL.n241 10.4732
R263 VTAIL.n222 VTAIL.n221 10.4732
R264 VTAIL.n154 VTAIL.n153 10.4732
R265 VTAIL.n134 VTAIL.n133 10.4732
R266 VTAIL.n302 VTAIL.n288 9.69747
R267 VTAIL.n331 VTAIL.n276 9.69747
R268 VTAIL.n350 VTAIL.n266 9.69747
R269 VTAIL.n38 VTAIL.n24 9.69747
R270 VTAIL.n67 VTAIL.n12 9.69747
R271 VTAIL.n86 VTAIL.n2 9.69747
R272 VTAIL.n264 VTAIL.n180 9.69747
R273 VTAIL.n245 VTAIL.n190 9.69747
R274 VTAIL.n218 VTAIL.n204 9.69747
R275 VTAIL.n176 VTAIL.n92 9.69747
R276 VTAIL.n157 VTAIL.n102 9.69747
R277 VTAIL.n130 VTAIL.n116 9.69747
R278 VTAIL.n350 VTAIL.n349 9.45567
R279 VTAIL.n86 VTAIL.n85 9.45567
R280 VTAIL.n264 VTAIL.n263 9.45567
R281 VTAIL.n176 VTAIL.n175 9.45567
R282 VTAIL.n341 VTAIL.n340 9.3005
R283 VTAIL.n343 VTAIL.n342 9.3005
R284 VTAIL.n268 VTAIL.n267 9.3005
R285 VTAIL.n349 VTAIL.n348 9.3005
R286 VTAIL.n335 VTAIL.n334 9.3005
R287 VTAIL.n333 VTAIL.n332 9.3005
R288 VTAIL.n276 VTAIL.n275 9.3005
R289 VTAIL.n327 VTAIL.n326 9.3005
R290 VTAIL.n325 VTAIL.n324 9.3005
R291 VTAIL.n280 VTAIL.n279 9.3005
R292 VTAIL.n319 VTAIL.n318 9.3005
R293 VTAIL.n292 VTAIL.n291 9.3005
R294 VTAIL.n299 VTAIL.n298 9.3005
R295 VTAIL.n301 VTAIL.n300 9.3005
R296 VTAIL.n288 VTAIL.n287 9.3005
R297 VTAIL.n307 VTAIL.n306 9.3005
R298 VTAIL.n309 VTAIL.n308 9.3005
R299 VTAIL.n310 VTAIL.n283 9.3005
R300 VTAIL.n317 VTAIL.n316 9.3005
R301 VTAIL.n272 VTAIL.n271 9.3005
R302 VTAIL.n77 VTAIL.n76 9.3005
R303 VTAIL.n79 VTAIL.n78 9.3005
R304 VTAIL.n4 VTAIL.n3 9.3005
R305 VTAIL.n85 VTAIL.n84 9.3005
R306 VTAIL.n71 VTAIL.n70 9.3005
R307 VTAIL.n69 VTAIL.n68 9.3005
R308 VTAIL.n12 VTAIL.n11 9.3005
R309 VTAIL.n63 VTAIL.n62 9.3005
R310 VTAIL.n61 VTAIL.n60 9.3005
R311 VTAIL.n16 VTAIL.n15 9.3005
R312 VTAIL.n55 VTAIL.n54 9.3005
R313 VTAIL.n28 VTAIL.n27 9.3005
R314 VTAIL.n35 VTAIL.n34 9.3005
R315 VTAIL.n37 VTAIL.n36 9.3005
R316 VTAIL.n24 VTAIL.n23 9.3005
R317 VTAIL.n43 VTAIL.n42 9.3005
R318 VTAIL.n45 VTAIL.n44 9.3005
R319 VTAIL.n46 VTAIL.n19 9.3005
R320 VTAIL.n53 VTAIL.n52 9.3005
R321 VTAIL.n8 VTAIL.n7 9.3005
R322 VTAIL.n182 VTAIL.n181 9.3005
R323 VTAIL.n257 VTAIL.n256 9.3005
R324 VTAIL.n255 VTAIL.n254 9.3005
R325 VTAIL.n186 VTAIL.n185 9.3005
R326 VTAIL.n249 VTAIL.n248 9.3005
R327 VTAIL.n247 VTAIL.n246 9.3005
R328 VTAIL.n190 VTAIL.n189 9.3005
R329 VTAIL.n241 VTAIL.n240 9.3005
R330 VTAIL.n239 VTAIL.n238 9.3005
R331 VTAIL.n194 VTAIL.n193 9.3005
R332 VTAIL.n233 VTAIL.n232 9.3005
R333 VTAIL.n231 VTAIL.n230 9.3005
R334 VTAIL.n199 VTAIL.n197 9.3005
R335 VTAIL.n225 VTAIL.n224 9.3005
R336 VTAIL.n223 VTAIL.n222 9.3005
R337 VTAIL.n204 VTAIL.n203 9.3005
R338 VTAIL.n217 VTAIL.n216 9.3005
R339 VTAIL.n215 VTAIL.n214 9.3005
R340 VTAIL.n208 VTAIL.n207 9.3005
R341 VTAIL.n263 VTAIL.n262 9.3005
R342 VTAIL.n120 VTAIL.n119 9.3005
R343 VTAIL.n127 VTAIL.n126 9.3005
R344 VTAIL.n129 VTAIL.n128 9.3005
R345 VTAIL.n116 VTAIL.n115 9.3005
R346 VTAIL.n135 VTAIL.n134 9.3005
R347 VTAIL.n137 VTAIL.n136 9.3005
R348 VTAIL.n111 VTAIL.n109 9.3005
R349 VTAIL.n143 VTAIL.n142 9.3005
R350 VTAIL.n169 VTAIL.n168 9.3005
R351 VTAIL.n94 VTAIL.n93 9.3005
R352 VTAIL.n175 VTAIL.n174 9.3005
R353 VTAIL.n167 VTAIL.n166 9.3005
R354 VTAIL.n98 VTAIL.n97 9.3005
R355 VTAIL.n161 VTAIL.n160 9.3005
R356 VTAIL.n159 VTAIL.n158 9.3005
R357 VTAIL.n102 VTAIL.n101 9.3005
R358 VTAIL.n153 VTAIL.n152 9.3005
R359 VTAIL.n151 VTAIL.n150 9.3005
R360 VTAIL.n106 VTAIL.n105 9.3005
R361 VTAIL.n145 VTAIL.n144 9.3005
R362 VTAIL.n301 VTAIL.n290 8.92171
R363 VTAIL.n332 VTAIL.n274 8.92171
R364 VTAIL.n348 VTAIL.n347 8.92171
R365 VTAIL.n37 VTAIL.n26 8.92171
R366 VTAIL.n68 VTAIL.n10 8.92171
R367 VTAIL.n84 VTAIL.n83 8.92171
R368 VTAIL.n262 VTAIL.n261 8.92171
R369 VTAIL.n246 VTAIL.n188 8.92171
R370 VTAIL.n217 VTAIL.n206 8.92171
R371 VTAIL.n174 VTAIL.n173 8.92171
R372 VTAIL.n158 VTAIL.n100 8.92171
R373 VTAIL.n129 VTAIL.n118 8.92171
R374 VTAIL.n298 VTAIL.n297 8.14595
R375 VTAIL.n336 VTAIL.n335 8.14595
R376 VTAIL.n344 VTAIL.n268 8.14595
R377 VTAIL.n34 VTAIL.n33 8.14595
R378 VTAIL.n72 VTAIL.n71 8.14595
R379 VTAIL.n80 VTAIL.n4 8.14595
R380 VTAIL.n258 VTAIL.n182 8.14595
R381 VTAIL.n250 VTAIL.n249 8.14595
R382 VTAIL.n214 VTAIL.n213 8.14595
R383 VTAIL.n170 VTAIL.n94 8.14595
R384 VTAIL.n162 VTAIL.n161 8.14595
R385 VTAIL.n126 VTAIL.n125 8.14595
R386 VTAIL.n294 VTAIL.n292 7.3702
R387 VTAIL.n339 VTAIL.n272 7.3702
R388 VTAIL.n343 VTAIL.n270 7.3702
R389 VTAIL.n30 VTAIL.n28 7.3702
R390 VTAIL.n75 VTAIL.n8 7.3702
R391 VTAIL.n79 VTAIL.n6 7.3702
R392 VTAIL.n257 VTAIL.n184 7.3702
R393 VTAIL.n253 VTAIL.n186 7.3702
R394 VTAIL.n210 VTAIL.n208 7.3702
R395 VTAIL.n169 VTAIL.n96 7.3702
R396 VTAIL.n165 VTAIL.n98 7.3702
R397 VTAIL.n122 VTAIL.n120 7.3702
R398 VTAIL.n340 VTAIL.n339 6.59444
R399 VTAIL.n340 VTAIL.n270 6.59444
R400 VTAIL.n76 VTAIL.n75 6.59444
R401 VTAIL.n76 VTAIL.n6 6.59444
R402 VTAIL.n254 VTAIL.n184 6.59444
R403 VTAIL.n254 VTAIL.n253 6.59444
R404 VTAIL.n166 VTAIL.n96 6.59444
R405 VTAIL.n166 VTAIL.n165 6.59444
R406 VTAIL.n297 VTAIL.n292 5.81868
R407 VTAIL.n336 VTAIL.n272 5.81868
R408 VTAIL.n344 VTAIL.n343 5.81868
R409 VTAIL.n33 VTAIL.n28 5.81868
R410 VTAIL.n72 VTAIL.n8 5.81868
R411 VTAIL.n80 VTAIL.n79 5.81868
R412 VTAIL.n258 VTAIL.n257 5.81868
R413 VTAIL.n250 VTAIL.n186 5.81868
R414 VTAIL.n213 VTAIL.n208 5.81868
R415 VTAIL.n170 VTAIL.n169 5.81868
R416 VTAIL.n162 VTAIL.n98 5.81868
R417 VTAIL.n125 VTAIL.n120 5.81868
R418 VTAIL.n298 VTAIL.n290 5.04292
R419 VTAIL.n335 VTAIL.n274 5.04292
R420 VTAIL.n347 VTAIL.n268 5.04292
R421 VTAIL.n34 VTAIL.n26 5.04292
R422 VTAIL.n71 VTAIL.n10 5.04292
R423 VTAIL.n83 VTAIL.n4 5.04292
R424 VTAIL.n261 VTAIL.n182 5.04292
R425 VTAIL.n249 VTAIL.n188 5.04292
R426 VTAIL.n214 VTAIL.n206 5.04292
R427 VTAIL.n173 VTAIL.n94 5.04292
R428 VTAIL.n161 VTAIL.n100 5.04292
R429 VTAIL.n126 VTAIL.n118 5.04292
R430 VTAIL.n302 VTAIL.n301 4.26717
R431 VTAIL.n332 VTAIL.n331 4.26717
R432 VTAIL.n348 VTAIL.n266 4.26717
R433 VTAIL.n38 VTAIL.n37 4.26717
R434 VTAIL.n68 VTAIL.n67 4.26717
R435 VTAIL.n84 VTAIL.n2 4.26717
R436 VTAIL.n262 VTAIL.n180 4.26717
R437 VTAIL.n246 VTAIL.n245 4.26717
R438 VTAIL.n218 VTAIL.n217 4.26717
R439 VTAIL.n174 VTAIL.n92 4.26717
R440 VTAIL.n158 VTAIL.n157 4.26717
R441 VTAIL.n130 VTAIL.n129 4.26717
R442 VTAIL.n305 VTAIL.n288 3.49141
R443 VTAIL.n328 VTAIL.n276 3.49141
R444 VTAIL.n41 VTAIL.n24 3.49141
R445 VTAIL.n64 VTAIL.n12 3.49141
R446 VTAIL.n242 VTAIL.n190 3.49141
R447 VTAIL.n221 VTAIL.n204 3.49141
R448 VTAIL.n154 VTAIL.n102 3.49141
R449 VTAIL.n133 VTAIL.n116 3.49141
R450 VTAIL.n306 VTAIL.n286 2.71565
R451 VTAIL.n327 VTAIL.n278 2.71565
R452 VTAIL.n42 VTAIL.n22 2.71565
R453 VTAIL.n63 VTAIL.n14 2.71565
R454 VTAIL.n241 VTAIL.n192 2.71565
R455 VTAIL.n222 VTAIL.n202 2.71565
R456 VTAIL.n153 VTAIL.n104 2.71565
R457 VTAIL.n134 VTAIL.n114 2.71565
R458 VTAIL.n293 VTAIL.n291 2.41282
R459 VTAIL.n29 VTAIL.n27 2.41282
R460 VTAIL.n209 VTAIL.n207 2.41282
R461 VTAIL.n121 VTAIL.n119 2.41282
R462 VTAIL.n0 VTAIL.t6 2.08282
R463 VTAIL.n0 VTAIL.t9 2.08282
R464 VTAIL.n88 VTAIL.t1 2.08282
R465 VTAIL.n88 VTAIL.t3 2.08282
R466 VTAIL.n178 VTAIL.t4 2.08282
R467 VTAIL.n178 VTAIL.t0 2.08282
R468 VTAIL.n90 VTAIL.t11 2.08282
R469 VTAIL.n90 VTAIL.t8 2.08282
R470 VTAIL.n311 VTAIL.n309 1.93989
R471 VTAIL.n324 VTAIL.n323 1.93989
R472 VTAIL.n47 VTAIL.n45 1.93989
R473 VTAIL.n60 VTAIL.n59 1.93989
R474 VTAIL.n238 VTAIL.n237 1.93989
R475 VTAIL.n226 VTAIL.n225 1.93989
R476 VTAIL.n150 VTAIL.n149 1.93989
R477 VTAIL.n138 VTAIL.n137 1.93989
R478 VTAIL.n177 VTAIL.n91 1.69016
R479 VTAIL.n265 VTAIL.n179 1.69016
R480 VTAIL.n89 VTAIL.n87 1.69016
R481 VTAIL.n179 VTAIL.n177 1.31516
R482 VTAIL.n87 VTAIL.n1 1.31516
R483 VTAIL VTAIL.n351 1.20955
R484 VTAIL.n310 VTAIL.n284 1.16414
R485 VTAIL.n320 VTAIL.n280 1.16414
R486 VTAIL.n46 VTAIL.n20 1.16414
R487 VTAIL.n56 VTAIL.n16 1.16414
R488 VTAIL.n234 VTAIL.n194 1.16414
R489 VTAIL.n229 VTAIL.n199 1.16414
R490 VTAIL.n146 VTAIL.n106 1.16414
R491 VTAIL.n141 VTAIL.n111 1.16414
R492 VTAIL VTAIL.n1 0.481103
R493 VTAIL.n316 VTAIL.n315 0.388379
R494 VTAIL.n319 VTAIL.n282 0.388379
R495 VTAIL.n52 VTAIL.n51 0.388379
R496 VTAIL.n55 VTAIL.n18 0.388379
R497 VTAIL.n233 VTAIL.n196 0.388379
R498 VTAIL.n230 VTAIL.n198 0.388379
R499 VTAIL.n145 VTAIL.n108 0.388379
R500 VTAIL.n142 VTAIL.n110 0.388379
R501 VTAIL.n299 VTAIL.n291 0.155672
R502 VTAIL.n300 VTAIL.n299 0.155672
R503 VTAIL.n300 VTAIL.n287 0.155672
R504 VTAIL.n307 VTAIL.n287 0.155672
R505 VTAIL.n308 VTAIL.n307 0.155672
R506 VTAIL.n308 VTAIL.n283 0.155672
R507 VTAIL.n317 VTAIL.n283 0.155672
R508 VTAIL.n318 VTAIL.n317 0.155672
R509 VTAIL.n318 VTAIL.n279 0.155672
R510 VTAIL.n325 VTAIL.n279 0.155672
R511 VTAIL.n326 VTAIL.n325 0.155672
R512 VTAIL.n326 VTAIL.n275 0.155672
R513 VTAIL.n333 VTAIL.n275 0.155672
R514 VTAIL.n334 VTAIL.n333 0.155672
R515 VTAIL.n334 VTAIL.n271 0.155672
R516 VTAIL.n341 VTAIL.n271 0.155672
R517 VTAIL.n342 VTAIL.n341 0.155672
R518 VTAIL.n342 VTAIL.n267 0.155672
R519 VTAIL.n349 VTAIL.n267 0.155672
R520 VTAIL.n35 VTAIL.n27 0.155672
R521 VTAIL.n36 VTAIL.n35 0.155672
R522 VTAIL.n36 VTAIL.n23 0.155672
R523 VTAIL.n43 VTAIL.n23 0.155672
R524 VTAIL.n44 VTAIL.n43 0.155672
R525 VTAIL.n44 VTAIL.n19 0.155672
R526 VTAIL.n53 VTAIL.n19 0.155672
R527 VTAIL.n54 VTAIL.n53 0.155672
R528 VTAIL.n54 VTAIL.n15 0.155672
R529 VTAIL.n61 VTAIL.n15 0.155672
R530 VTAIL.n62 VTAIL.n61 0.155672
R531 VTAIL.n62 VTAIL.n11 0.155672
R532 VTAIL.n69 VTAIL.n11 0.155672
R533 VTAIL.n70 VTAIL.n69 0.155672
R534 VTAIL.n70 VTAIL.n7 0.155672
R535 VTAIL.n77 VTAIL.n7 0.155672
R536 VTAIL.n78 VTAIL.n77 0.155672
R537 VTAIL.n78 VTAIL.n3 0.155672
R538 VTAIL.n85 VTAIL.n3 0.155672
R539 VTAIL.n263 VTAIL.n181 0.155672
R540 VTAIL.n256 VTAIL.n181 0.155672
R541 VTAIL.n256 VTAIL.n255 0.155672
R542 VTAIL.n255 VTAIL.n185 0.155672
R543 VTAIL.n248 VTAIL.n185 0.155672
R544 VTAIL.n248 VTAIL.n247 0.155672
R545 VTAIL.n247 VTAIL.n189 0.155672
R546 VTAIL.n240 VTAIL.n189 0.155672
R547 VTAIL.n240 VTAIL.n239 0.155672
R548 VTAIL.n239 VTAIL.n193 0.155672
R549 VTAIL.n232 VTAIL.n193 0.155672
R550 VTAIL.n232 VTAIL.n231 0.155672
R551 VTAIL.n231 VTAIL.n197 0.155672
R552 VTAIL.n224 VTAIL.n197 0.155672
R553 VTAIL.n224 VTAIL.n223 0.155672
R554 VTAIL.n223 VTAIL.n203 0.155672
R555 VTAIL.n216 VTAIL.n203 0.155672
R556 VTAIL.n216 VTAIL.n215 0.155672
R557 VTAIL.n215 VTAIL.n207 0.155672
R558 VTAIL.n175 VTAIL.n93 0.155672
R559 VTAIL.n168 VTAIL.n93 0.155672
R560 VTAIL.n168 VTAIL.n167 0.155672
R561 VTAIL.n167 VTAIL.n97 0.155672
R562 VTAIL.n160 VTAIL.n97 0.155672
R563 VTAIL.n160 VTAIL.n159 0.155672
R564 VTAIL.n159 VTAIL.n101 0.155672
R565 VTAIL.n152 VTAIL.n101 0.155672
R566 VTAIL.n152 VTAIL.n151 0.155672
R567 VTAIL.n151 VTAIL.n105 0.155672
R568 VTAIL.n144 VTAIL.n105 0.155672
R569 VTAIL.n144 VTAIL.n143 0.155672
R570 VTAIL.n143 VTAIL.n109 0.155672
R571 VTAIL.n136 VTAIL.n109 0.155672
R572 VTAIL.n136 VTAIL.n135 0.155672
R573 VTAIL.n135 VTAIL.n115 0.155672
R574 VTAIL.n128 VTAIL.n115 0.155672
R575 VTAIL.n128 VTAIL.n127 0.155672
R576 VTAIL.n127 VTAIL.n119 0.155672
R577 VDD2.n167 VDD2.n87 756.745
R578 VDD2.n80 VDD2.n0 756.745
R579 VDD2.n168 VDD2.n167 585
R580 VDD2.n166 VDD2.n165 585
R581 VDD2.n91 VDD2.n90 585
R582 VDD2.n160 VDD2.n159 585
R583 VDD2.n158 VDD2.n157 585
R584 VDD2.n95 VDD2.n94 585
R585 VDD2.n152 VDD2.n151 585
R586 VDD2.n150 VDD2.n149 585
R587 VDD2.n99 VDD2.n98 585
R588 VDD2.n144 VDD2.n143 585
R589 VDD2.n142 VDD2.n141 585
R590 VDD2.n103 VDD2.n102 585
R591 VDD2.n107 VDD2.n105 585
R592 VDD2.n136 VDD2.n135 585
R593 VDD2.n134 VDD2.n133 585
R594 VDD2.n109 VDD2.n108 585
R595 VDD2.n128 VDD2.n127 585
R596 VDD2.n126 VDD2.n125 585
R597 VDD2.n113 VDD2.n112 585
R598 VDD2.n120 VDD2.n119 585
R599 VDD2.n118 VDD2.n117 585
R600 VDD2.n29 VDD2.n28 585
R601 VDD2.n31 VDD2.n30 585
R602 VDD2.n24 VDD2.n23 585
R603 VDD2.n37 VDD2.n36 585
R604 VDD2.n39 VDD2.n38 585
R605 VDD2.n20 VDD2.n19 585
R606 VDD2.n46 VDD2.n45 585
R607 VDD2.n47 VDD2.n18 585
R608 VDD2.n49 VDD2.n48 585
R609 VDD2.n16 VDD2.n15 585
R610 VDD2.n55 VDD2.n54 585
R611 VDD2.n57 VDD2.n56 585
R612 VDD2.n12 VDD2.n11 585
R613 VDD2.n63 VDD2.n62 585
R614 VDD2.n65 VDD2.n64 585
R615 VDD2.n8 VDD2.n7 585
R616 VDD2.n71 VDD2.n70 585
R617 VDD2.n73 VDD2.n72 585
R618 VDD2.n4 VDD2.n3 585
R619 VDD2.n79 VDD2.n78 585
R620 VDD2.n81 VDD2.n80 585
R621 VDD2.n116 VDD2.t4 329.036
R622 VDD2.n27 VDD2.t5 329.036
R623 VDD2.n167 VDD2.n166 171.744
R624 VDD2.n166 VDD2.n90 171.744
R625 VDD2.n159 VDD2.n90 171.744
R626 VDD2.n159 VDD2.n158 171.744
R627 VDD2.n158 VDD2.n94 171.744
R628 VDD2.n151 VDD2.n94 171.744
R629 VDD2.n151 VDD2.n150 171.744
R630 VDD2.n150 VDD2.n98 171.744
R631 VDD2.n143 VDD2.n98 171.744
R632 VDD2.n143 VDD2.n142 171.744
R633 VDD2.n142 VDD2.n102 171.744
R634 VDD2.n107 VDD2.n102 171.744
R635 VDD2.n135 VDD2.n107 171.744
R636 VDD2.n135 VDD2.n134 171.744
R637 VDD2.n134 VDD2.n108 171.744
R638 VDD2.n127 VDD2.n108 171.744
R639 VDD2.n127 VDD2.n126 171.744
R640 VDD2.n126 VDD2.n112 171.744
R641 VDD2.n119 VDD2.n112 171.744
R642 VDD2.n119 VDD2.n118 171.744
R643 VDD2.n30 VDD2.n29 171.744
R644 VDD2.n30 VDD2.n23 171.744
R645 VDD2.n37 VDD2.n23 171.744
R646 VDD2.n38 VDD2.n37 171.744
R647 VDD2.n38 VDD2.n19 171.744
R648 VDD2.n46 VDD2.n19 171.744
R649 VDD2.n47 VDD2.n46 171.744
R650 VDD2.n48 VDD2.n47 171.744
R651 VDD2.n48 VDD2.n15 171.744
R652 VDD2.n55 VDD2.n15 171.744
R653 VDD2.n56 VDD2.n55 171.744
R654 VDD2.n56 VDD2.n11 171.744
R655 VDD2.n63 VDD2.n11 171.744
R656 VDD2.n64 VDD2.n63 171.744
R657 VDD2.n64 VDD2.n7 171.744
R658 VDD2.n71 VDD2.n7 171.744
R659 VDD2.n72 VDD2.n71 171.744
R660 VDD2.n72 VDD2.n3 171.744
R661 VDD2.n79 VDD2.n3 171.744
R662 VDD2.n80 VDD2.n79 171.744
R663 VDD2.n118 VDD2.t4 85.8723
R664 VDD2.n29 VDD2.t5 85.8723
R665 VDD2.n86 VDD2.n85 68.7728
R666 VDD2 VDD2.n173 68.77
R667 VDD2.n86 VDD2.n84 47.9427
R668 VDD2.n172 VDD2.n171 46.7308
R669 VDD2.n172 VDD2.n86 42.6636
R670 VDD2.n105 VDD2.n103 13.1884
R671 VDD2.n49 VDD2.n16 13.1884
R672 VDD2.n141 VDD2.n140 12.8005
R673 VDD2.n137 VDD2.n136 12.8005
R674 VDD2.n50 VDD2.n18 12.8005
R675 VDD2.n54 VDD2.n53 12.8005
R676 VDD2.n144 VDD2.n101 12.0247
R677 VDD2.n133 VDD2.n106 12.0247
R678 VDD2.n45 VDD2.n44 12.0247
R679 VDD2.n57 VDD2.n14 12.0247
R680 VDD2.n145 VDD2.n99 11.249
R681 VDD2.n132 VDD2.n109 11.249
R682 VDD2.n43 VDD2.n20 11.249
R683 VDD2.n58 VDD2.n12 11.249
R684 VDD2.n117 VDD2.n116 10.7239
R685 VDD2.n28 VDD2.n27 10.7239
R686 VDD2.n149 VDD2.n148 10.4732
R687 VDD2.n129 VDD2.n128 10.4732
R688 VDD2.n40 VDD2.n39 10.4732
R689 VDD2.n62 VDD2.n61 10.4732
R690 VDD2.n171 VDD2.n87 9.69747
R691 VDD2.n152 VDD2.n97 9.69747
R692 VDD2.n125 VDD2.n111 9.69747
R693 VDD2.n36 VDD2.n22 9.69747
R694 VDD2.n65 VDD2.n10 9.69747
R695 VDD2.n84 VDD2.n0 9.69747
R696 VDD2.n171 VDD2.n170 9.45567
R697 VDD2.n84 VDD2.n83 9.45567
R698 VDD2.n115 VDD2.n114 9.3005
R699 VDD2.n122 VDD2.n121 9.3005
R700 VDD2.n124 VDD2.n123 9.3005
R701 VDD2.n111 VDD2.n110 9.3005
R702 VDD2.n130 VDD2.n129 9.3005
R703 VDD2.n132 VDD2.n131 9.3005
R704 VDD2.n106 VDD2.n104 9.3005
R705 VDD2.n138 VDD2.n137 9.3005
R706 VDD2.n164 VDD2.n163 9.3005
R707 VDD2.n89 VDD2.n88 9.3005
R708 VDD2.n170 VDD2.n169 9.3005
R709 VDD2.n162 VDD2.n161 9.3005
R710 VDD2.n93 VDD2.n92 9.3005
R711 VDD2.n156 VDD2.n155 9.3005
R712 VDD2.n154 VDD2.n153 9.3005
R713 VDD2.n97 VDD2.n96 9.3005
R714 VDD2.n148 VDD2.n147 9.3005
R715 VDD2.n146 VDD2.n145 9.3005
R716 VDD2.n101 VDD2.n100 9.3005
R717 VDD2.n140 VDD2.n139 9.3005
R718 VDD2.n75 VDD2.n74 9.3005
R719 VDD2.n77 VDD2.n76 9.3005
R720 VDD2.n2 VDD2.n1 9.3005
R721 VDD2.n83 VDD2.n82 9.3005
R722 VDD2.n69 VDD2.n68 9.3005
R723 VDD2.n67 VDD2.n66 9.3005
R724 VDD2.n10 VDD2.n9 9.3005
R725 VDD2.n61 VDD2.n60 9.3005
R726 VDD2.n59 VDD2.n58 9.3005
R727 VDD2.n14 VDD2.n13 9.3005
R728 VDD2.n53 VDD2.n52 9.3005
R729 VDD2.n26 VDD2.n25 9.3005
R730 VDD2.n33 VDD2.n32 9.3005
R731 VDD2.n35 VDD2.n34 9.3005
R732 VDD2.n22 VDD2.n21 9.3005
R733 VDD2.n41 VDD2.n40 9.3005
R734 VDD2.n43 VDD2.n42 9.3005
R735 VDD2.n44 VDD2.n17 9.3005
R736 VDD2.n51 VDD2.n50 9.3005
R737 VDD2.n6 VDD2.n5 9.3005
R738 VDD2.n169 VDD2.n168 8.92171
R739 VDD2.n153 VDD2.n95 8.92171
R740 VDD2.n124 VDD2.n113 8.92171
R741 VDD2.n35 VDD2.n24 8.92171
R742 VDD2.n66 VDD2.n8 8.92171
R743 VDD2.n82 VDD2.n81 8.92171
R744 VDD2.n165 VDD2.n89 8.14595
R745 VDD2.n157 VDD2.n156 8.14595
R746 VDD2.n121 VDD2.n120 8.14595
R747 VDD2.n32 VDD2.n31 8.14595
R748 VDD2.n70 VDD2.n69 8.14595
R749 VDD2.n78 VDD2.n2 8.14595
R750 VDD2.n164 VDD2.n91 7.3702
R751 VDD2.n160 VDD2.n93 7.3702
R752 VDD2.n117 VDD2.n115 7.3702
R753 VDD2.n28 VDD2.n26 7.3702
R754 VDD2.n73 VDD2.n6 7.3702
R755 VDD2.n77 VDD2.n4 7.3702
R756 VDD2.n161 VDD2.n91 6.59444
R757 VDD2.n161 VDD2.n160 6.59444
R758 VDD2.n74 VDD2.n73 6.59444
R759 VDD2.n74 VDD2.n4 6.59444
R760 VDD2.n165 VDD2.n164 5.81868
R761 VDD2.n157 VDD2.n93 5.81868
R762 VDD2.n120 VDD2.n115 5.81868
R763 VDD2.n31 VDD2.n26 5.81868
R764 VDD2.n70 VDD2.n6 5.81868
R765 VDD2.n78 VDD2.n77 5.81868
R766 VDD2.n168 VDD2.n89 5.04292
R767 VDD2.n156 VDD2.n95 5.04292
R768 VDD2.n121 VDD2.n113 5.04292
R769 VDD2.n32 VDD2.n24 5.04292
R770 VDD2.n69 VDD2.n8 5.04292
R771 VDD2.n81 VDD2.n2 5.04292
R772 VDD2.n169 VDD2.n87 4.26717
R773 VDD2.n153 VDD2.n152 4.26717
R774 VDD2.n125 VDD2.n124 4.26717
R775 VDD2.n36 VDD2.n35 4.26717
R776 VDD2.n66 VDD2.n65 4.26717
R777 VDD2.n82 VDD2.n0 4.26717
R778 VDD2.n149 VDD2.n97 3.49141
R779 VDD2.n128 VDD2.n111 3.49141
R780 VDD2.n39 VDD2.n22 3.49141
R781 VDD2.n62 VDD2.n10 3.49141
R782 VDD2.n148 VDD2.n99 2.71565
R783 VDD2.n129 VDD2.n109 2.71565
R784 VDD2.n40 VDD2.n20 2.71565
R785 VDD2.n61 VDD2.n12 2.71565
R786 VDD2.n116 VDD2.n114 2.41282
R787 VDD2.n27 VDD2.n25 2.41282
R788 VDD2.n173 VDD2.t0 2.08282
R789 VDD2.n173 VDD2.t2 2.08282
R790 VDD2.n85 VDD2.t3 2.08282
R791 VDD2.n85 VDD2.t1 2.08282
R792 VDD2.n145 VDD2.n144 1.93989
R793 VDD2.n133 VDD2.n132 1.93989
R794 VDD2.n45 VDD2.n43 1.93989
R795 VDD2.n58 VDD2.n57 1.93989
R796 VDD2 VDD2.n172 1.32593
R797 VDD2.n141 VDD2.n101 1.16414
R798 VDD2.n136 VDD2.n106 1.16414
R799 VDD2.n44 VDD2.n18 1.16414
R800 VDD2.n54 VDD2.n14 1.16414
R801 VDD2.n140 VDD2.n103 0.388379
R802 VDD2.n137 VDD2.n105 0.388379
R803 VDD2.n50 VDD2.n49 0.388379
R804 VDD2.n53 VDD2.n16 0.388379
R805 VDD2.n170 VDD2.n88 0.155672
R806 VDD2.n163 VDD2.n88 0.155672
R807 VDD2.n163 VDD2.n162 0.155672
R808 VDD2.n162 VDD2.n92 0.155672
R809 VDD2.n155 VDD2.n92 0.155672
R810 VDD2.n155 VDD2.n154 0.155672
R811 VDD2.n154 VDD2.n96 0.155672
R812 VDD2.n147 VDD2.n96 0.155672
R813 VDD2.n147 VDD2.n146 0.155672
R814 VDD2.n146 VDD2.n100 0.155672
R815 VDD2.n139 VDD2.n100 0.155672
R816 VDD2.n139 VDD2.n138 0.155672
R817 VDD2.n138 VDD2.n104 0.155672
R818 VDD2.n131 VDD2.n104 0.155672
R819 VDD2.n131 VDD2.n130 0.155672
R820 VDD2.n130 VDD2.n110 0.155672
R821 VDD2.n123 VDD2.n110 0.155672
R822 VDD2.n123 VDD2.n122 0.155672
R823 VDD2.n122 VDD2.n114 0.155672
R824 VDD2.n33 VDD2.n25 0.155672
R825 VDD2.n34 VDD2.n33 0.155672
R826 VDD2.n34 VDD2.n21 0.155672
R827 VDD2.n41 VDD2.n21 0.155672
R828 VDD2.n42 VDD2.n41 0.155672
R829 VDD2.n42 VDD2.n17 0.155672
R830 VDD2.n51 VDD2.n17 0.155672
R831 VDD2.n52 VDD2.n51 0.155672
R832 VDD2.n52 VDD2.n13 0.155672
R833 VDD2.n59 VDD2.n13 0.155672
R834 VDD2.n60 VDD2.n59 0.155672
R835 VDD2.n60 VDD2.n9 0.155672
R836 VDD2.n67 VDD2.n9 0.155672
R837 VDD2.n68 VDD2.n67 0.155672
R838 VDD2.n68 VDD2.n5 0.155672
R839 VDD2.n75 VDD2.n5 0.155672
R840 VDD2.n76 VDD2.n75 0.155672
R841 VDD2.n76 VDD2.n1 0.155672
R842 VDD2.n83 VDD2.n1 0.155672
R843 B.n500 B.n79 585
R844 B.n502 B.n501 585
R845 B.n503 B.n78 585
R846 B.n505 B.n504 585
R847 B.n506 B.n77 585
R848 B.n508 B.n507 585
R849 B.n509 B.n76 585
R850 B.n511 B.n510 585
R851 B.n512 B.n75 585
R852 B.n514 B.n513 585
R853 B.n515 B.n74 585
R854 B.n517 B.n516 585
R855 B.n518 B.n73 585
R856 B.n520 B.n519 585
R857 B.n521 B.n72 585
R858 B.n523 B.n522 585
R859 B.n524 B.n71 585
R860 B.n526 B.n525 585
R861 B.n527 B.n70 585
R862 B.n529 B.n528 585
R863 B.n530 B.n69 585
R864 B.n532 B.n531 585
R865 B.n533 B.n68 585
R866 B.n535 B.n534 585
R867 B.n536 B.n67 585
R868 B.n538 B.n537 585
R869 B.n539 B.n66 585
R870 B.n541 B.n540 585
R871 B.n542 B.n65 585
R872 B.n544 B.n543 585
R873 B.n545 B.n64 585
R874 B.n547 B.n546 585
R875 B.n548 B.n63 585
R876 B.n550 B.n549 585
R877 B.n551 B.n62 585
R878 B.n553 B.n552 585
R879 B.n554 B.n61 585
R880 B.n556 B.n555 585
R881 B.n557 B.n60 585
R882 B.n559 B.n558 585
R883 B.n560 B.n59 585
R884 B.n562 B.n561 585
R885 B.n563 B.n58 585
R886 B.n565 B.n564 585
R887 B.n566 B.n57 585
R888 B.n568 B.n567 585
R889 B.n569 B.n56 585
R890 B.n571 B.n570 585
R891 B.n572 B.n55 585
R892 B.n574 B.n573 585
R893 B.n575 B.n51 585
R894 B.n577 B.n576 585
R895 B.n578 B.n50 585
R896 B.n580 B.n579 585
R897 B.n581 B.n49 585
R898 B.n583 B.n582 585
R899 B.n584 B.n48 585
R900 B.n586 B.n585 585
R901 B.n587 B.n47 585
R902 B.n589 B.n588 585
R903 B.n590 B.n46 585
R904 B.n592 B.n591 585
R905 B.n594 B.n43 585
R906 B.n596 B.n595 585
R907 B.n597 B.n42 585
R908 B.n599 B.n598 585
R909 B.n600 B.n41 585
R910 B.n602 B.n601 585
R911 B.n603 B.n40 585
R912 B.n605 B.n604 585
R913 B.n606 B.n39 585
R914 B.n608 B.n607 585
R915 B.n609 B.n38 585
R916 B.n611 B.n610 585
R917 B.n612 B.n37 585
R918 B.n614 B.n613 585
R919 B.n615 B.n36 585
R920 B.n617 B.n616 585
R921 B.n618 B.n35 585
R922 B.n620 B.n619 585
R923 B.n621 B.n34 585
R924 B.n623 B.n622 585
R925 B.n624 B.n33 585
R926 B.n626 B.n625 585
R927 B.n627 B.n32 585
R928 B.n629 B.n628 585
R929 B.n630 B.n31 585
R930 B.n632 B.n631 585
R931 B.n633 B.n30 585
R932 B.n635 B.n634 585
R933 B.n636 B.n29 585
R934 B.n638 B.n637 585
R935 B.n639 B.n28 585
R936 B.n641 B.n640 585
R937 B.n642 B.n27 585
R938 B.n644 B.n643 585
R939 B.n645 B.n26 585
R940 B.n647 B.n646 585
R941 B.n648 B.n25 585
R942 B.n650 B.n649 585
R943 B.n651 B.n24 585
R944 B.n653 B.n652 585
R945 B.n654 B.n23 585
R946 B.n656 B.n655 585
R947 B.n657 B.n22 585
R948 B.n659 B.n658 585
R949 B.n660 B.n21 585
R950 B.n662 B.n661 585
R951 B.n663 B.n20 585
R952 B.n665 B.n664 585
R953 B.n666 B.n19 585
R954 B.n668 B.n667 585
R955 B.n669 B.n18 585
R956 B.n671 B.n670 585
R957 B.n499 B.n498 585
R958 B.n497 B.n80 585
R959 B.n496 B.n495 585
R960 B.n494 B.n81 585
R961 B.n493 B.n492 585
R962 B.n491 B.n82 585
R963 B.n490 B.n489 585
R964 B.n488 B.n83 585
R965 B.n487 B.n486 585
R966 B.n485 B.n84 585
R967 B.n484 B.n483 585
R968 B.n482 B.n85 585
R969 B.n481 B.n480 585
R970 B.n479 B.n86 585
R971 B.n478 B.n477 585
R972 B.n476 B.n87 585
R973 B.n475 B.n474 585
R974 B.n473 B.n88 585
R975 B.n472 B.n471 585
R976 B.n470 B.n89 585
R977 B.n469 B.n468 585
R978 B.n467 B.n90 585
R979 B.n466 B.n465 585
R980 B.n464 B.n91 585
R981 B.n463 B.n462 585
R982 B.n461 B.n92 585
R983 B.n460 B.n459 585
R984 B.n458 B.n93 585
R985 B.n457 B.n456 585
R986 B.n455 B.n94 585
R987 B.n454 B.n453 585
R988 B.n452 B.n95 585
R989 B.n451 B.n450 585
R990 B.n449 B.n96 585
R991 B.n448 B.n447 585
R992 B.n446 B.n97 585
R993 B.n445 B.n444 585
R994 B.n443 B.n98 585
R995 B.n442 B.n441 585
R996 B.n440 B.n99 585
R997 B.n439 B.n438 585
R998 B.n437 B.n100 585
R999 B.n436 B.n435 585
R1000 B.n434 B.n101 585
R1001 B.n433 B.n432 585
R1002 B.n431 B.n102 585
R1003 B.n430 B.n429 585
R1004 B.n428 B.n103 585
R1005 B.n427 B.n426 585
R1006 B.n425 B.n104 585
R1007 B.n424 B.n423 585
R1008 B.n422 B.n105 585
R1009 B.n421 B.n420 585
R1010 B.n419 B.n106 585
R1011 B.n418 B.n417 585
R1012 B.n416 B.n107 585
R1013 B.n415 B.n414 585
R1014 B.n413 B.n108 585
R1015 B.n412 B.n411 585
R1016 B.n410 B.n109 585
R1017 B.n409 B.n408 585
R1018 B.n407 B.n110 585
R1019 B.n406 B.n405 585
R1020 B.n233 B.n172 585
R1021 B.n235 B.n234 585
R1022 B.n236 B.n171 585
R1023 B.n238 B.n237 585
R1024 B.n239 B.n170 585
R1025 B.n241 B.n240 585
R1026 B.n242 B.n169 585
R1027 B.n244 B.n243 585
R1028 B.n245 B.n168 585
R1029 B.n247 B.n246 585
R1030 B.n248 B.n167 585
R1031 B.n250 B.n249 585
R1032 B.n251 B.n166 585
R1033 B.n253 B.n252 585
R1034 B.n254 B.n165 585
R1035 B.n256 B.n255 585
R1036 B.n257 B.n164 585
R1037 B.n259 B.n258 585
R1038 B.n260 B.n163 585
R1039 B.n262 B.n261 585
R1040 B.n263 B.n162 585
R1041 B.n265 B.n264 585
R1042 B.n266 B.n161 585
R1043 B.n268 B.n267 585
R1044 B.n269 B.n160 585
R1045 B.n271 B.n270 585
R1046 B.n272 B.n159 585
R1047 B.n274 B.n273 585
R1048 B.n275 B.n158 585
R1049 B.n277 B.n276 585
R1050 B.n278 B.n157 585
R1051 B.n280 B.n279 585
R1052 B.n281 B.n156 585
R1053 B.n283 B.n282 585
R1054 B.n284 B.n155 585
R1055 B.n286 B.n285 585
R1056 B.n287 B.n154 585
R1057 B.n289 B.n288 585
R1058 B.n290 B.n153 585
R1059 B.n292 B.n291 585
R1060 B.n293 B.n152 585
R1061 B.n295 B.n294 585
R1062 B.n296 B.n151 585
R1063 B.n298 B.n297 585
R1064 B.n299 B.n150 585
R1065 B.n301 B.n300 585
R1066 B.n302 B.n149 585
R1067 B.n304 B.n303 585
R1068 B.n305 B.n148 585
R1069 B.n307 B.n306 585
R1070 B.n308 B.n147 585
R1071 B.n310 B.n309 585
R1072 B.n312 B.n144 585
R1073 B.n314 B.n313 585
R1074 B.n315 B.n143 585
R1075 B.n317 B.n316 585
R1076 B.n318 B.n142 585
R1077 B.n320 B.n319 585
R1078 B.n321 B.n141 585
R1079 B.n323 B.n322 585
R1080 B.n324 B.n140 585
R1081 B.n326 B.n325 585
R1082 B.n328 B.n327 585
R1083 B.n329 B.n136 585
R1084 B.n331 B.n330 585
R1085 B.n332 B.n135 585
R1086 B.n334 B.n333 585
R1087 B.n335 B.n134 585
R1088 B.n337 B.n336 585
R1089 B.n338 B.n133 585
R1090 B.n340 B.n339 585
R1091 B.n341 B.n132 585
R1092 B.n343 B.n342 585
R1093 B.n344 B.n131 585
R1094 B.n346 B.n345 585
R1095 B.n347 B.n130 585
R1096 B.n349 B.n348 585
R1097 B.n350 B.n129 585
R1098 B.n352 B.n351 585
R1099 B.n353 B.n128 585
R1100 B.n355 B.n354 585
R1101 B.n356 B.n127 585
R1102 B.n358 B.n357 585
R1103 B.n359 B.n126 585
R1104 B.n361 B.n360 585
R1105 B.n362 B.n125 585
R1106 B.n364 B.n363 585
R1107 B.n365 B.n124 585
R1108 B.n367 B.n366 585
R1109 B.n368 B.n123 585
R1110 B.n370 B.n369 585
R1111 B.n371 B.n122 585
R1112 B.n373 B.n372 585
R1113 B.n374 B.n121 585
R1114 B.n376 B.n375 585
R1115 B.n377 B.n120 585
R1116 B.n379 B.n378 585
R1117 B.n380 B.n119 585
R1118 B.n382 B.n381 585
R1119 B.n383 B.n118 585
R1120 B.n385 B.n384 585
R1121 B.n386 B.n117 585
R1122 B.n388 B.n387 585
R1123 B.n389 B.n116 585
R1124 B.n391 B.n390 585
R1125 B.n392 B.n115 585
R1126 B.n394 B.n393 585
R1127 B.n395 B.n114 585
R1128 B.n397 B.n396 585
R1129 B.n398 B.n113 585
R1130 B.n400 B.n399 585
R1131 B.n401 B.n112 585
R1132 B.n403 B.n402 585
R1133 B.n404 B.n111 585
R1134 B.n232 B.n231 585
R1135 B.n230 B.n173 585
R1136 B.n229 B.n228 585
R1137 B.n227 B.n174 585
R1138 B.n226 B.n225 585
R1139 B.n224 B.n175 585
R1140 B.n223 B.n222 585
R1141 B.n221 B.n176 585
R1142 B.n220 B.n219 585
R1143 B.n218 B.n177 585
R1144 B.n217 B.n216 585
R1145 B.n215 B.n178 585
R1146 B.n214 B.n213 585
R1147 B.n212 B.n179 585
R1148 B.n211 B.n210 585
R1149 B.n209 B.n180 585
R1150 B.n208 B.n207 585
R1151 B.n206 B.n181 585
R1152 B.n205 B.n204 585
R1153 B.n203 B.n182 585
R1154 B.n202 B.n201 585
R1155 B.n200 B.n183 585
R1156 B.n199 B.n198 585
R1157 B.n197 B.n184 585
R1158 B.n196 B.n195 585
R1159 B.n194 B.n185 585
R1160 B.n193 B.n192 585
R1161 B.n191 B.n186 585
R1162 B.n190 B.n189 585
R1163 B.n188 B.n187 585
R1164 B.n2 B.n0 585
R1165 B.n717 B.n1 585
R1166 B.n716 B.n715 585
R1167 B.n714 B.n3 585
R1168 B.n713 B.n712 585
R1169 B.n711 B.n4 585
R1170 B.n710 B.n709 585
R1171 B.n708 B.n5 585
R1172 B.n707 B.n706 585
R1173 B.n705 B.n6 585
R1174 B.n704 B.n703 585
R1175 B.n702 B.n7 585
R1176 B.n701 B.n700 585
R1177 B.n699 B.n8 585
R1178 B.n698 B.n697 585
R1179 B.n696 B.n9 585
R1180 B.n695 B.n694 585
R1181 B.n693 B.n10 585
R1182 B.n692 B.n691 585
R1183 B.n690 B.n11 585
R1184 B.n689 B.n688 585
R1185 B.n687 B.n12 585
R1186 B.n686 B.n685 585
R1187 B.n684 B.n13 585
R1188 B.n683 B.n682 585
R1189 B.n681 B.n14 585
R1190 B.n680 B.n679 585
R1191 B.n678 B.n15 585
R1192 B.n677 B.n676 585
R1193 B.n675 B.n16 585
R1194 B.n674 B.n673 585
R1195 B.n672 B.n17 585
R1196 B.n719 B.n718 585
R1197 B.n231 B.n172 530.939
R1198 B.n670 B.n17 530.939
R1199 B.n405 B.n404 530.939
R1200 B.n500 B.n499 530.939
R1201 B.n137 B.t2 478.853
R1202 B.n52 B.t7 478.853
R1203 B.n145 B.t11 478.853
R1204 B.n44 B.t4 478.853
R1205 B.n138 B.t1 440.841
R1206 B.n53 B.t8 440.841
R1207 B.n146 B.t10 440.841
R1208 B.n45 B.t5 440.841
R1209 B.n137 B.t0 436.692
R1210 B.n145 B.t9 436.692
R1211 B.n44 B.t3 436.692
R1212 B.n52 B.t6 436.692
R1213 B.n231 B.n230 163.367
R1214 B.n230 B.n229 163.367
R1215 B.n229 B.n174 163.367
R1216 B.n225 B.n174 163.367
R1217 B.n225 B.n224 163.367
R1218 B.n224 B.n223 163.367
R1219 B.n223 B.n176 163.367
R1220 B.n219 B.n176 163.367
R1221 B.n219 B.n218 163.367
R1222 B.n218 B.n217 163.367
R1223 B.n217 B.n178 163.367
R1224 B.n213 B.n178 163.367
R1225 B.n213 B.n212 163.367
R1226 B.n212 B.n211 163.367
R1227 B.n211 B.n180 163.367
R1228 B.n207 B.n180 163.367
R1229 B.n207 B.n206 163.367
R1230 B.n206 B.n205 163.367
R1231 B.n205 B.n182 163.367
R1232 B.n201 B.n182 163.367
R1233 B.n201 B.n200 163.367
R1234 B.n200 B.n199 163.367
R1235 B.n199 B.n184 163.367
R1236 B.n195 B.n184 163.367
R1237 B.n195 B.n194 163.367
R1238 B.n194 B.n193 163.367
R1239 B.n193 B.n186 163.367
R1240 B.n189 B.n186 163.367
R1241 B.n189 B.n188 163.367
R1242 B.n188 B.n2 163.367
R1243 B.n718 B.n2 163.367
R1244 B.n718 B.n717 163.367
R1245 B.n717 B.n716 163.367
R1246 B.n716 B.n3 163.367
R1247 B.n712 B.n3 163.367
R1248 B.n712 B.n711 163.367
R1249 B.n711 B.n710 163.367
R1250 B.n710 B.n5 163.367
R1251 B.n706 B.n5 163.367
R1252 B.n706 B.n705 163.367
R1253 B.n705 B.n704 163.367
R1254 B.n704 B.n7 163.367
R1255 B.n700 B.n7 163.367
R1256 B.n700 B.n699 163.367
R1257 B.n699 B.n698 163.367
R1258 B.n698 B.n9 163.367
R1259 B.n694 B.n9 163.367
R1260 B.n694 B.n693 163.367
R1261 B.n693 B.n692 163.367
R1262 B.n692 B.n11 163.367
R1263 B.n688 B.n11 163.367
R1264 B.n688 B.n687 163.367
R1265 B.n687 B.n686 163.367
R1266 B.n686 B.n13 163.367
R1267 B.n682 B.n13 163.367
R1268 B.n682 B.n681 163.367
R1269 B.n681 B.n680 163.367
R1270 B.n680 B.n15 163.367
R1271 B.n676 B.n15 163.367
R1272 B.n676 B.n675 163.367
R1273 B.n675 B.n674 163.367
R1274 B.n674 B.n17 163.367
R1275 B.n235 B.n172 163.367
R1276 B.n236 B.n235 163.367
R1277 B.n237 B.n236 163.367
R1278 B.n237 B.n170 163.367
R1279 B.n241 B.n170 163.367
R1280 B.n242 B.n241 163.367
R1281 B.n243 B.n242 163.367
R1282 B.n243 B.n168 163.367
R1283 B.n247 B.n168 163.367
R1284 B.n248 B.n247 163.367
R1285 B.n249 B.n248 163.367
R1286 B.n249 B.n166 163.367
R1287 B.n253 B.n166 163.367
R1288 B.n254 B.n253 163.367
R1289 B.n255 B.n254 163.367
R1290 B.n255 B.n164 163.367
R1291 B.n259 B.n164 163.367
R1292 B.n260 B.n259 163.367
R1293 B.n261 B.n260 163.367
R1294 B.n261 B.n162 163.367
R1295 B.n265 B.n162 163.367
R1296 B.n266 B.n265 163.367
R1297 B.n267 B.n266 163.367
R1298 B.n267 B.n160 163.367
R1299 B.n271 B.n160 163.367
R1300 B.n272 B.n271 163.367
R1301 B.n273 B.n272 163.367
R1302 B.n273 B.n158 163.367
R1303 B.n277 B.n158 163.367
R1304 B.n278 B.n277 163.367
R1305 B.n279 B.n278 163.367
R1306 B.n279 B.n156 163.367
R1307 B.n283 B.n156 163.367
R1308 B.n284 B.n283 163.367
R1309 B.n285 B.n284 163.367
R1310 B.n285 B.n154 163.367
R1311 B.n289 B.n154 163.367
R1312 B.n290 B.n289 163.367
R1313 B.n291 B.n290 163.367
R1314 B.n291 B.n152 163.367
R1315 B.n295 B.n152 163.367
R1316 B.n296 B.n295 163.367
R1317 B.n297 B.n296 163.367
R1318 B.n297 B.n150 163.367
R1319 B.n301 B.n150 163.367
R1320 B.n302 B.n301 163.367
R1321 B.n303 B.n302 163.367
R1322 B.n303 B.n148 163.367
R1323 B.n307 B.n148 163.367
R1324 B.n308 B.n307 163.367
R1325 B.n309 B.n308 163.367
R1326 B.n309 B.n144 163.367
R1327 B.n314 B.n144 163.367
R1328 B.n315 B.n314 163.367
R1329 B.n316 B.n315 163.367
R1330 B.n316 B.n142 163.367
R1331 B.n320 B.n142 163.367
R1332 B.n321 B.n320 163.367
R1333 B.n322 B.n321 163.367
R1334 B.n322 B.n140 163.367
R1335 B.n326 B.n140 163.367
R1336 B.n327 B.n326 163.367
R1337 B.n327 B.n136 163.367
R1338 B.n331 B.n136 163.367
R1339 B.n332 B.n331 163.367
R1340 B.n333 B.n332 163.367
R1341 B.n333 B.n134 163.367
R1342 B.n337 B.n134 163.367
R1343 B.n338 B.n337 163.367
R1344 B.n339 B.n338 163.367
R1345 B.n339 B.n132 163.367
R1346 B.n343 B.n132 163.367
R1347 B.n344 B.n343 163.367
R1348 B.n345 B.n344 163.367
R1349 B.n345 B.n130 163.367
R1350 B.n349 B.n130 163.367
R1351 B.n350 B.n349 163.367
R1352 B.n351 B.n350 163.367
R1353 B.n351 B.n128 163.367
R1354 B.n355 B.n128 163.367
R1355 B.n356 B.n355 163.367
R1356 B.n357 B.n356 163.367
R1357 B.n357 B.n126 163.367
R1358 B.n361 B.n126 163.367
R1359 B.n362 B.n361 163.367
R1360 B.n363 B.n362 163.367
R1361 B.n363 B.n124 163.367
R1362 B.n367 B.n124 163.367
R1363 B.n368 B.n367 163.367
R1364 B.n369 B.n368 163.367
R1365 B.n369 B.n122 163.367
R1366 B.n373 B.n122 163.367
R1367 B.n374 B.n373 163.367
R1368 B.n375 B.n374 163.367
R1369 B.n375 B.n120 163.367
R1370 B.n379 B.n120 163.367
R1371 B.n380 B.n379 163.367
R1372 B.n381 B.n380 163.367
R1373 B.n381 B.n118 163.367
R1374 B.n385 B.n118 163.367
R1375 B.n386 B.n385 163.367
R1376 B.n387 B.n386 163.367
R1377 B.n387 B.n116 163.367
R1378 B.n391 B.n116 163.367
R1379 B.n392 B.n391 163.367
R1380 B.n393 B.n392 163.367
R1381 B.n393 B.n114 163.367
R1382 B.n397 B.n114 163.367
R1383 B.n398 B.n397 163.367
R1384 B.n399 B.n398 163.367
R1385 B.n399 B.n112 163.367
R1386 B.n403 B.n112 163.367
R1387 B.n404 B.n403 163.367
R1388 B.n405 B.n110 163.367
R1389 B.n409 B.n110 163.367
R1390 B.n410 B.n409 163.367
R1391 B.n411 B.n410 163.367
R1392 B.n411 B.n108 163.367
R1393 B.n415 B.n108 163.367
R1394 B.n416 B.n415 163.367
R1395 B.n417 B.n416 163.367
R1396 B.n417 B.n106 163.367
R1397 B.n421 B.n106 163.367
R1398 B.n422 B.n421 163.367
R1399 B.n423 B.n422 163.367
R1400 B.n423 B.n104 163.367
R1401 B.n427 B.n104 163.367
R1402 B.n428 B.n427 163.367
R1403 B.n429 B.n428 163.367
R1404 B.n429 B.n102 163.367
R1405 B.n433 B.n102 163.367
R1406 B.n434 B.n433 163.367
R1407 B.n435 B.n434 163.367
R1408 B.n435 B.n100 163.367
R1409 B.n439 B.n100 163.367
R1410 B.n440 B.n439 163.367
R1411 B.n441 B.n440 163.367
R1412 B.n441 B.n98 163.367
R1413 B.n445 B.n98 163.367
R1414 B.n446 B.n445 163.367
R1415 B.n447 B.n446 163.367
R1416 B.n447 B.n96 163.367
R1417 B.n451 B.n96 163.367
R1418 B.n452 B.n451 163.367
R1419 B.n453 B.n452 163.367
R1420 B.n453 B.n94 163.367
R1421 B.n457 B.n94 163.367
R1422 B.n458 B.n457 163.367
R1423 B.n459 B.n458 163.367
R1424 B.n459 B.n92 163.367
R1425 B.n463 B.n92 163.367
R1426 B.n464 B.n463 163.367
R1427 B.n465 B.n464 163.367
R1428 B.n465 B.n90 163.367
R1429 B.n469 B.n90 163.367
R1430 B.n470 B.n469 163.367
R1431 B.n471 B.n470 163.367
R1432 B.n471 B.n88 163.367
R1433 B.n475 B.n88 163.367
R1434 B.n476 B.n475 163.367
R1435 B.n477 B.n476 163.367
R1436 B.n477 B.n86 163.367
R1437 B.n481 B.n86 163.367
R1438 B.n482 B.n481 163.367
R1439 B.n483 B.n482 163.367
R1440 B.n483 B.n84 163.367
R1441 B.n487 B.n84 163.367
R1442 B.n488 B.n487 163.367
R1443 B.n489 B.n488 163.367
R1444 B.n489 B.n82 163.367
R1445 B.n493 B.n82 163.367
R1446 B.n494 B.n493 163.367
R1447 B.n495 B.n494 163.367
R1448 B.n495 B.n80 163.367
R1449 B.n499 B.n80 163.367
R1450 B.n670 B.n669 163.367
R1451 B.n669 B.n668 163.367
R1452 B.n668 B.n19 163.367
R1453 B.n664 B.n19 163.367
R1454 B.n664 B.n663 163.367
R1455 B.n663 B.n662 163.367
R1456 B.n662 B.n21 163.367
R1457 B.n658 B.n21 163.367
R1458 B.n658 B.n657 163.367
R1459 B.n657 B.n656 163.367
R1460 B.n656 B.n23 163.367
R1461 B.n652 B.n23 163.367
R1462 B.n652 B.n651 163.367
R1463 B.n651 B.n650 163.367
R1464 B.n650 B.n25 163.367
R1465 B.n646 B.n25 163.367
R1466 B.n646 B.n645 163.367
R1467 B.n645 B.n644 163.367
R1468 B.n644 B.n27 163.367
R1469 B.n640 B.n27 163.367
R1470 B.n640 B.n639 163.367
R1471 B.n639 B.n638 163.367
R1472 B.n638 B.n29 163.367
R1473 B.n634 B.n29 163.367
R1474 B.n634 B.n633 163.367
R1475 B.n633 B.n632 163.367
R1476 B.n632 B.n31 163.367
R1477 B.n628 B.n31 163.367
R1478 B.n628 B.n627 163.367
R1479 B.n627 B.n626 163.367
R1480 B.n626 B.n33 163.367
R1481 B.n622 B.n33 163.367
R1482 B.n622 B.n621 163.367
R1483 B.n621 B.n620 163.367
R1484 B.n620 B.n35 163.367
R1485 B.n616 B.n35 163.367
R1486 B.n616 B.n615 163.367
R1487 B.n615 B.n614 163.367
R1488 B.n614 B.n37 163.367
R1489 B.n610 B.n37 163.367
R1490 B.n610 B.n609 163.367
R1491 B.n609 B.n608 163.367
R1492 B.n608 B.n39 163.367
R1493 B.n604 B.n39 163.367
R1494 B.n604 B.n603 163.367
R1495 B.n603 B.n602 163.367
R1496 B.n602 B.n41 163.367
R1497 B.n598 B.n41 163.367
R1498 B.n598 B.n597 163.367
R1499 B.n597 B.n596 163.367
R1500 B.n596 B.n43 163.367
R1501 B.n591 B.n43 163.367
R1502 B.n591 B.n590 163.367
R1503 B.n590 B.n589 163.367
R1504 B.n589 B.n47 163.367
R1505 B.n585 B.n47 163.367
R1506 B.n585 B.n584 163.367
R1507 B.n584 B.n583 163.367
R1508 B.n583 B.n49 163.367
R1509 B.n579 B.n49 163.367
R1510 B.n579 B.n578 163.367
R1511 B.n578 B.n577 163.367
R1512 B.n577 B.n51 163.367
R1513 B.n573 B.n51 163.367
R1514 B.n573 B.n572 163.367
R1515 B.n572 B.n571 163.367
R1516 B.n571 B.n56 163.367
R1517 B.n567 B.n56 163.367
R1518 B.n567 B.n566 163.367
R1519 B.n566 B.n565 163.367
R1520 B.n565 B.n58 163.367
R1521 B.n561 B.n58 163.367
R1522 B.n561 B.n560 163.367
R1523 B.n560 B.n559 163.367
R1524 B.n559 B.n60 163.367
R1525 B.n555 B.n60 163.367
R1526 B.n555 B.n554 163.367
R1527 B.n554 B.n553 163.367
R1528 B.n553 B.n62 163.367
R1529 B.n549 B.n62 163.367
R1530 B.n549 B.n548 163.367
R1531 B.n548 B.n547 163.367
R1532 B.n547 B.n64 163.367
R1533 B.n543 B.n64 163.367
R1534 B.n543 B.n542 163.367
R1535 B.n542 B.n541 163.367
R1536 B.n541 B.n66 163.367
R1537 B.n537 B.n66 163.367
R1538 B.n537 B.n536 163.367
R1539 B.n536 B.n535 163.367
R1540 B.n535 B.n68 163.367
R1541 B.n531 B.n68 163.367
R1542 B.n531 B.n530 163.367
R1543 B.n530 B.n529 163.367
R1544 B.n529 B.n70 163.367
R1545 B.n525 B.n70 163.367
R1546 B.n525 B.n524 163.367
R1547 B.n524 B.n523 163.367
R1548 B.n523 B.n72 163.367
R1549 B.n519 B.n72 163.367
R1550 B.n519 B.n518 163.367
R1551 B.n518 B.n517 163.367
R1552 B.n517 B.n74 163.367
R1553 B.n513 B.n74 163.367
R1554 B.n513 B.n512 163.367
R1555 B.n512 B.n511 163.367
R1556 B.n511 B.n76 163.367
R1557 B.n507 B.n76 163.367
R1558 B.n507 B.n506 163.367
R1559 B.n506 B.n505 163.367
R1560 B.n505 B.n78 163.367
R1561 B.n501 B.n78 163.367
R1562 B.n501 B.n500 163.367
R1563 B.n139 B.n138 59.5399
R1564 B.n311 B.n146 59.5399
R1565 B.n593 B.n45 59.5399
R1566 B.n54 B.n53 59.5399
R1567 B.n138 B.n137 38.0126
R1568 B.n146 B.n145 38.0126
R1569 B.n45 B.n44 38.0126
R1570 B.n53 B.n52 38.0126
R1571 B.n672 B.n671 34.4981
R1572 B.n498 B.n79 34.4981
R1573 B.n406 B.n111 34.4981
R1574 B.n233 B.n232 34.4981
R1575 B B.n719 18.0485
R1576 B.n671 B.n18 10.6151
R1577 B.n667 B.n18 10.6151
R1578 B.n667 B.n666 10.6151
R1579 B.n666 B.n665 10.6151
R1580 B.n665 B.n20 10.6151
R1581 B.n661 B.n20 10.6151
R1582 B.n661 B.n660 10.6151
R1583 B.n660 B.n659 10.6151
R1584 B.n659 B.n22 10.6151
R1585 B.n655 B.n22 10.6151
R1586 B.n655 B.n654 10.6151
R1587 B.n654 B.n653 10.6151
R1588 B.n653 B.n24 10.6151
R1589 B.n649 B.n24 10.6151
R1590 B.n649 B.n648 10.6151
R1591 B.n648 B.n647 10.6151
R1592 B.n647 B.n26 10.6151
R1593 B.n643 B.n26 10.6151
R1594 B.n643 B.n642 10.6151
R1595 B.n642 B.n641 10.6151
R1596 B.n641 B.n28 10.6151
R1597 B.n637 B.n28 10.6151
R1598 B.n637 B.n636 10.6151
R1599 B.n636 B.n635 10.6151
R1600 B.n635 B.n30 10.6151
R1601 B.n631 B.n30 10.6151
R1602 B.n631 B.n630 10.6151
R1603 B.n630 B.n629 10.6151
R1604 B.n629 B.n32 10.6151
R1605 B.n625 B.n32 10.6151
R1606 B.n625 B.n624 10.6151
R1607 B.n624 B.n623 10.6151
R1608 B.n623 B.n34 10.6151
R1609 B.n619 B.n34 10.6151
R1610 B.n619 B.n618 10.6151
R1611 B.n618 B.n617 10.6151
R1612 B.n617 B.n36 10.6151
R1613 B.n613 B.n36 10.6151
R1614 B.n613 B.n612 10.6151
R1615 B.n612 B.n611 10.6151
R1616 B.n611 B.n38 10.6151
R1617 B.n607 B.n38 10.6151
R1618 B.n607 B.n606 10.6151
R1619 B.n606 B.n605 10.6151
R1620 B.n605 B.n40 10.6151
R1621 B.n601 B.n40 10.6151
R1622 B.n601 B.n600 10.6151
R1623 B.n600 B.n599 10.6151
R1624 B.n599 B.n42 10.6151
R1625 B.n595 B.n42 10.6151
R1626 B.n595 B.n594 10.6151
R1627 B.n592 B.n46 10.6151
R1628 B.n588 B.n46 10.6151
R1629 B.n588 B.n587 10.6151
R1630 B.n587 B.n586 10.6151
R1631 B.n586 B.n48 10.6151
R1632 B.n582 B.n48 10.6151
R1633 B.n582 B.n581 10.6151
R1634 B.n581 B.n580 10.6151
R1635 B.n580 B.n50 10.6151
R1636 B.n576 B.n575 10.6151
R1637 B.n575 B.n574 10.6151
R1638 B.n574 B.n55 10.6151
R1639 B.n570 B.n55 10.6151
R1640 B.n570 B.n569 10.6151
R1641 B.n569 B.n568 10.6151
R1642 B.n568 B.n57 10.6151
R1643 B.n564 B.n57 10.6151
R1644 B.n564 B.n563 10.6151
R1645 B.n563 B.n562 10.6151
R1646 B.n562 B.n59 10.6151
R1647 B.n558 B.n59 10.6151
R1648 B.n558 B.n557 10.6151
R1649 B.n557 B.n556 10.6151
R1650 B.n556 B.n61 10.6151
R1651 B.n552 B.n61 10.6151
R1652 B.n552 B.n551 10.6151
R1653 B.n551 B.n550 10.6151
R1654 B.n550 B.n63 10.6151
R1655 B.n546 B.n63 10.6151
R1656 B.n546 B.n545 10.6151
R1657 B.n545 B.n544 10.6151
R1658 B.n544 B.n65 10.6151
R1659 B.n540 B.n65 10.6151
R1660 B.n540 B.n539 10.6151
R1661 B.n539 B.n538 10.6151
R1662 B.n538 B.n67 10.6151
R1663 B.n534 B.n67 10.6151
R1664 B.n534 B.n533 10.6151
R1665 B.n533 B.n532 10.6151
R1666 B.n532 B.n69 10.6151
R1667 B.n528 B.n69 10.6151
R1668 B.n528 B.n527 10.6151
R1669 B.n527 B.n526 10.6151
R1670 B.n526 B.n71 10.6151
R1671 B.n522 B.n71 10.6151
R1672 B.n522 B.n521 10.6151
R1673 B.n521 B.n520 10.6151
R1674 B.n520 B.n73 10.6151
R1675 B.n516 B.n73 10.6151
R1676 B.n516 B.n515 10.6151
R1677 B.n515 B.n514 10.6151
R1678 B.n514 B.n75 10.6151
R1679 B.n510 B.n75 10.6151
R1680 B.n510 B.n509 10.6151
R1681 B.n509 B.n508 10.6151
R1682 B.n508 B.n77 10.6151
R1683 B.n504 B.n77 10.6151
R1684 B.n504 B.n503 10.6151
R1685 B.n503 B.n502 10.6151
R1686 B.n502 B.n79 10.6151
R1687 B.n407 B.n406 10.6151
R1688 B.n408 B.n407 10.6151
R1689 B.n408 B.n109 10.6151
R1690 B.n412 B.n109 10.6151
R1691 B.n413 B.n412 10.6151
R1692 B.n414 B.n413 10.6151
R1693 B.n414 B.n107 10.6151
R1694 B.n418 B.n107 10.6151
R1695 B.n419 B.n418 10.6151
R1696 B.n420 B.n419 10.6151
R1697 B.n420 B.n105 10.6151
R1698 B.n424 B.n105 10.6151
R1699 B.n425 B.n424 10.6151
R1700 B.n426 B.n425 10.6151
R1701 B.n426 B.n103 10.6151
R1702 B.n430 B.n103 10.6151
R1703 B.n431 B.n430 10.6151
R1704 B.n432 B.n431 10.6151
R1705 B.n432 B.n101 10.6151
R1706 B.n436 B.n101 10.6151
R1707 B.n437 B.n436 10.6151
R1708 B.n438 B.n437 10.6151
R1709 B.n438 B.n99 10.6151
R1710 B.n442 B.n99 10.6151
R1711 B.n443 B.n442 10.6151
R1712 B.n444 B.n443 10.6151
R1713 B.n444 B.n97 10.6151
R1714 B.n448 B.n97 10.6151
R1715 B.n449 B.n448 10.6151
R1716 B.n450 B.n449 10.6151
R1717 B.n450 B.n95 10.6151
R1718 B.n454 B.n95 10.6151
R1719 B.n455 B.n454 10.6151
R1720 B.n456 B.n455 10.6151
R1721 B.n456 B.n93 10.6151
R1722 B.n460 B.n93 10.6151
R1723 B.n461 B.n460 10.6151
R1724 B.n462 B.n461 10.6151
R1725 B.n462 B.n91 10.6151
R1726 B.n466 B.n91 10.6151
R1727 B.n467 B.n466 10.6151
R1728 B.n468 B.n467 10.6151
R1729 B.n468 B.n89 10.6151
R1730 B.n472 B.n89 10.6151
R1731 B.n473 B.n472 10.6151
R1732 B.n474 B.n473 10.6151
R1733 B.n474 B.n87 10.6151
R1734 B.n478 B.n87 10.6151
R1735 B.n479 B.n478 10.6151
R1736 B.n480 B.n479 10.6151
R1737 B.n480 B.n85 10.6151
R1738 B.n484 B.n85 10.6151
R1739 B.n485 B.n484 10.6151
R1740 B.n486 B.n485 10.6151
R1741 B.n486 B.n83 10.6151
R1742 B.n490 B.n83 10.6151
R1743 B.n491 B.n490 10.6151
R1744 B.n492 B.n491 10.6151
R1745 B.n492 B.n81 10.6151
R1746 B.n496 B.n81 10.6151
R1747 B.n497 B.n496 10.6151
R1748 B.n498 B.n497 10.6151
R1749 B.n234 B.n233 10.6151
R1750 B.n234 B.n171 10.6151
R1751 B.n238 B.n171 10.6151
R1752 B.n239 B.n238 10.6151
R1753 B.n240 B.n239 10.6151
R1754 B.n240 B.n169 10.6151
R1755 B.n244 B.n169 10.6151
R1756 B.n245 B.n244 10.6151
R1757 B.n246 B.n245 10.6151
R1758 B.n246 B.n167 10.6151
R1759 B.n250 B.n167 10.6151
R1760 B.n251 B.n250 10.6151
R1761 B.n252 B.n251 10.6151
R1762 B.n252 B.n165 10.6151
R1763 B.n256 B.n165 10.6151
R1764 B.n257 B.n256 10.6151
R1765 B.n258 B.n257 10.6151
R1766 B.n258 B.n163 10.6151
R1767 B.n262 B.n163 10.6151
R1768 B.n263 B.n262 10.6151
R1769 B.n264 B.n263 10.6151
R1770 B.n264 B.n161 10.6151
R1771 B.n268 B.n161 10.6151
R1772 B.n269 B.n268 10.6151
R1773 B.n270 B.n269 10.6151
R1774 B.n270 B.n159 10.6151
R1775 B.n274 B.n159 10.6151
R1776 B.n275 B.n274 10.6151
R1777 B.n276 B.n275 10.6151
R1778 B.n276 B.n157 10.6151
R1779 B.n280 B.n157 10.6151
R1780 B.n281 B.n280 10.6151
R1781 B.n282 B.n281 10.6151
R1782 B.n282 B.n155 10.6151
R1783 B.n286 B.n155 10.6151
R1784 B.n287 B.n286 10.6151
R1785 B.n288 B.n287 10.6151
R1786 B.n288 B.n153 10.6151
R1787 B.n292 B.n153 10.6151
R1788 B.n293 B.n292 10.6151
R1789 B.n294 B.n293 10.6151
R1790 B.n294 B.n151 10.6151
R1791 B.n298 B.n151 10.6151
R1792 B.n299 B.n298 10.6151
R1793 B.n300 B.n299 10.6151
R1794 B.n300 B.n149 10.6151
R1795 B.n304 B.n149 10.6151
R1796 B.n305 B.n304 10.6151
R1797 B.n306 B.n305 10.6151
R1798 B.n306 B.n147 10.6151
R1799 B.n310 B.n147 10.6151
R1800 B.n313 B.n312 10.6151
R1801 B.n313 B.n143 10.6151
R1802 B.n317 B.n143 10.6151
R1803 B.n318 B.n317 10.6151
R1804 B.n319 B.n318 10.6151
R1805 B.n319 B.n141 10.6151
R1806 B.n323 B.n141 10.6151
R1807 B.n324 B.n323 10.6151
R1808 B.n325 B.n324 10.6151
R1809 B.n329 B.n328 10.6151
R1810 B.n330 B.n329 10.6151
R1811 B.n330 B.n135 10.6151
R1812 B.n334 B.n135 10.6151
R1813 B.n335 B.n334 10.6151
R1814 B.n336 B.n335 10.6151
R1815 B.n336 B.n133 10.6151
R1816 B.n340 B.n133 10.6151
R1817 B.n341 B.n340 10.6151
R1818 B.n342 B.n341 10.6151
R1819 B.n342 B.n131 10.6151
R1820 B.n346 B.n131 10.6151
R1821 B.n347 B.n346 10.6151
R1822 B.n348 B.n347 10.6151
R1823 B.n348 B.n129 10.6151
R1824 B.n352 B.n129 10.6151
R1825 B.n353 B.n352 10.6151
R1826 B.n354 B.n353 10.6151
R1827 B.n354 B.n127 10.6151
R1828 B.n358 B.n127 10.6151
R1829 B.n359 B.n358 10.6151
R1830 B.n360 B.n359 10.6151
R1831 B.n360 B.n125 10.6151
R1832 B.n364 B.n125 10.6151
R1833 B.n365 B.n364 10.6151
R1834 B.n366 B.n365 10.6151
R1835 B.n366 B.n123 10.6151
R1836 B.n370 B.n123 10.6151
R1837 B.n371 B.n370 10.6151
R1838 B.n372 B.n371 10.6151
R1839 B.n372 B.n121 10.6151
R1840 B.n376 B.n121 10.6151
R1841 B.n377 B.n376 10.6151
R1842 B.n378 B.n377 10.6151
R1843 B.n378 B.n119 10.6151
R1844 B.n382 B.n119 10.6151
R1845 B.n383 B.n382 10.6151
R1846 B.n384 B.n383 10.6151
R1847 B.n384 B.n117 10.6151
R1848 B.n388 B.n117 10.6151
R1849 B.n389 B.n388 10.6151
R1850 B.n390 B.n389 10.6151
R1851 B.n390 B.n115 10.6151
R1852 B.n394 B.n115 10.6151
R1853 B.n395 B.n394 10.6151
R1854 B.n396 B.n395 10.6151
R1855 B.n396 B.n113 10.6151
R1856 B.n400 B.n113 10.6151
R1857 B.n401 B.n400 10.6151
R1858 B.n402 B.n401 10.6151
R1859 B.n402 B.n111 10.6151
R1860 B.n232 B.n173 10.6151
R1861 B.n228 B.n173 10.6151
R1862 B.n228 B.n227 10.6151
R1863 B.n227 B.n226 10.6151
R1864 B.n226 B.n175 10.6151
R1865 B.n222 B.n175 10.6151
R1866 B.n222 B.n221 10.6151
R1867 B.n221 B.n220 10.6151
R1868 B.n220 B.n177 10.6151
R1869 B.n216 B.n177 10.6151
R1870 B.n216 B.n215 10.6151
R1871 B.n215 B.n214 10.6151
R1872 B.n214 B.n179 10.6151
R1873 B.n210 B.n179 10.6151
R1874 B.n210 B.n209 10.6151
R1875 B.n209 B.n208 10.6151
R1876 B.n208 B.n181 10.6151
R1877 B.n204 B.n181 10.6151
R1878 B.n204 B.n203 10.6151
R1879 B.n203 B.n202 10.6151
R1880 B.n202 B.n183 10.6151
R1881 B.n198 B.n183 10.6151
R1882 B.n198 B.n197 10.6151
R1883 B.n197 B.n196 10.6151
R1884 B.n196 B.n185 10.6151
R1885 B.n192 B.n185 10.6151
R1886 B.n192 B.n191 10.6151
R1887 B.n191 B.n190 10.6151
R1888 B.n190 B.n187 10.6151
R1889 B.n187 B.n0 10.6151
R1890 B.n715 B.n1 10.6151
R1891 B.n715 B.n714 10.6151
R1892 B.n714 B.n713 10.6151
R1893 B.n713 B.n4 10.6151
R1894 B.n709 B.n4 10.6151
R1895 B.n709 B.n708 10.6151
R1896 B.n708 B.n707 10.6151
R1897 B.n707 B.n6 10.6151
R1898 B.n703 B.n6 10.6151
R1899 B.n703 B.n702 10.6151
R1900 B.n702 B.n701 10.6151
R1901 B.n701 B.n8 10.6151
R1902 B.n697 B.n8 10.6151
R1903 B.n697 B.n696 10.6151
R1904 B.n696 B.n695 10.6151
R1905 B.n695 B.n10 10.6151
R1906 B.n691 B.n10 10.6151
R1907 B.n691 B.n690 10.6151
R1908 B.n690 B.n689 10.6151
R1909 B.n689 B.n12 10.6151
R1910 B.n685 B.n12 10.6151
R1911 B.n685 B.n684 10.6151
R1912 B.n684 B.n683 10.6151
R1913 B.n683 B.n14 10.6151
R1914 B.n679 B.n14 10.6151
R1915 B.n679 B.n678 10.6151
R1916 B.n678 B.n677 10.6151
R1917 B.n677 B.n16 10.6151
R1918 B.n673 B.n16 10.6151
R1919 B.n673 B.n672 10.6151
R1920 B.n594 B.n593 9.36635
R1921 B.n576 B.n54 9.36635
R1922 B.n311 B.n310 9.36635
R1923 B.n328 B.n139 9.36635
R1924 B.n719 B.n0 2.81026
R1925 B.n719 B.n1 2.81026
R1926 B.n593 B.n592 1.24928
R1927 B.n54 B.n50 1.24928
R1928 B.n312 B.n311 1.24928
R1929 B.n325 B.n139 1.24928
R1930 VP.n6 VP.t5 264.673
R1931 VP.n17 VP.t4 230.798
R1932 VP.n24 VP.t2 230.798
R1933 VP.n31 VP.t1 230.798
R1934 VP.n14 VP.t3 230.798
R1935 VP.n7 VP.t0 230.798
R1936 VP.n17 VP.n16 175.492
R1937 VP.n32 VP.n31 175.492
R1938 VP.n15 VP.n14 175.492
R1939 VP.n9 VP.n8 161.3
R1940 VP.n10 VP.n5 161.3
R1941 VP.n12 VP.n11 161.3
R1942 VP.n13 VP.n4 161.3
R1943 VP.n30 VP.n0 161.3
R1944 VP.n29 VP.n28 161.3
R1945 VP.n27 VP.n1 161.3
R1946 VP.n26 VP.n25 161.3
R1947 VP.n23 VP.n2 161.3
R1948 VP.n22 VP.n21 161.3
R1949 VP.n20 VP.n3 161.3
R1950 VP.n19 VP.n18 161.3
R1951 VP.n22 VP.n3 56.5193
R1952 VP.n29 VP.n1 56.5193
R1953 VP.n12 VP.n5 56.5193
R1954 VP.n7 VP.n6 54.1657
R1955 VP.n16 VP.n15 47.5687
R1956 VP.n18 VP.n3 24.4675
R1957 VP.n23 VP.n22 24.4675
R1958 VP.n25 VP.n1 24.4675
R1959 VP.n30 VP.n29 24.4675
R1960 VP.n13 VP.n12 24.4675
R1961 VP.n8 VP.n5 24.4675
R1962 VP.n9 VP.n6 17.7577
R1963 VP.n24 VP.n23 12.234
R1964 VP.n25 VP.n24 12.234
R1965 VP.n8 VP.n7 12.234
R1966 VP.n18 VP.n17 10.2766
R1967 VP.n31 VP.n30 10.2766
R1968 VP.n14 VP.n13 10.2766
R1969 VP.n10 VP.n9 0.189894
R1970 VP.n11 VP.n10 0.189894
R1971 VP.n11 VP.n4 0.189894
R1972 VP.n15 VP.n4 0.189894
R1973 VP.n19 VP.n16 0.189894
R1974 VP.n20 VP.n19 0.189894
R1975 VP.n21 VP.n20 0.189894
R1976 VP.n21 VP.n2 0.189894
R1977 VP.n26 VP.n2 0.189894
R1978 VP.n27 VP.n26 0.189894
R1979 VP.n28 VP.n27 0.189894
R1980 VP.n28 VP.n0 0.189894
R1981 VP.n32 VP.n0 0.189894
R1982 VP VP.n32 0.0516364
R1983 VDD1.n80 VDD1.n0 756.745
R1984 VDD1.n165 VDD1.n85 756.745
R1985 VDD1.n81 VDD1.n80 585
R1986 VDD1.n79 VDD1.n78 585
R1987 VDD1.n4 VDD1.n3 585
R1988 VDD1.n73 VDD1.n72 585
R1989 VDD1.n71 VDD1.n70 585
R1990 VDD1.n8 VDD1.n7 585
R1991 VDD1.n65 VDD1.n64 585
R1992 VDD1.n63 VDD1.n62 585
R1993 VDD1.n12 VDD1.n11 585
R1994 VDD1.n57 VDD1.n56 585
R1995 VDD1.n55 VDD1.n54 585
R1996 VDD1.n16 VDD1.n15 585
R1997 VDD1.n20 VDD1.n18 585
R1998 VDD1.n49 VDD1.n48 585
R1999 VDD1.n47 VDD1.n46 585
R2000 VDD1.n22 VDD1.n21 585
R2001 VDD1.n41 VDD1.n40 585
R2002 VDD1.n39 VDD1.n38 585
R2003 VDD1.n26 VDD1.n25 585
R2004 VDD1.n33 VDD1.n32 585
R2005 VDD1.n31 VDD1.n30 585
R2006 VDD1.n114 VDD1.n113 585
R2007 VDD1.n116 VDD1.n115 585
R2008 VDD1.n109 VDD1.n108 585
R2009 VDD1.n122 VDD1.n121 585
R2010 VDD1.n124 VDD1.n123 585
R2011 VDD1.n105 VDD1.n104 585
R2012 VDD1.n131 VDD1.n130 585
R2013 VDD1.n132 VDD1.n103 585
R2014 VDD1.n134 VDD1.n133 585
R2015 VDD1.n101 VDD1.n100 585
R2016 VDD1.n140 VDD1.n139 585
R2017 VDD1.n142 VDD1.n141 585
R2018 VDD1.n97 VDD1.n96 585
R2019 VDD1.n148 VDD1.n147 585
R2020 VDD1.n150 VDD1.n149 585
R2021 VDD1.n93 VDD1.n92 585
R2022 VDD1.n156 VDD1.n155 585
R2023 VDD1.n158 VDD1.n157 585
R2024 VDD1.n89 VDD1.n88 585
R2025 VDD1.n164 VDD1.n163 585
R2026 VDD1.n166 VDD1.n165 585
R2027 VDD1.n29 VDD1.t0 329.036
R2028 VDD1.n112 VDD1.t1 329.036
R2029 VDD1.n80 VDD1.n79 171.744
R2030 VDD1.n79 VDD1.n3 171.744
R2031 VDD1.n72 VDD1.n3 171.744
R2032 VDD1.n72 VDD1.n71 171.744
R2033 VDD1.n71 VDD1.n7 171.744
R2034 VDD1.n64 VDD1.n7 171.744
R2035 VDD1.n64 VDD1.n63 171.744
R2036 VDD1.n63 VDD1.n11 171.744
R2037 VDD1.n56 VDD1.n11 171.744
R2038 VDD1.n56 VDD1.n55 171.744
R2039 VDD1.n55 VDD1.n15 171.744
R2040 VDD1.n20 VDD1.n15 171.744
R2041 VDD1.n48 VDD1.n20 171.744
R2042 VDD1.n48 VDD1.n47 171.744
R2043 VDD1.n47 VDD1.n21 171.744
R2044 VDD1.n40 VDD1.n21 171.744
R2045 VDD1.n40 VDD1.n39 171.744
R2046 VDD1.n39 VDD1.n25 171.744
R2047 VDD1.n32 VDD1.n25 171.744
R2048 VDD1.n32 VDD1.n31 171.744
R2049 VDD1.n115 VDD1.n114 171.744
R2050 VDD1.n115 VDD1.n108 171.744
R2051 VDD1.n122 VDD1.n108 171.744
R2052 VDD1.n123 VDD1.n122 171.744
R2053 VDD1.n123 VDD1.n104 171.744
R2054 VDD1.n131 VDD1.n104 171.744
R2055 VDD1.n132 VDD1.n131 171.744
R2056 VDD1.n133 VDD1.n132 171.744
R2057 VDD1.n133 VDD1.n100 171.744
R2058 VDD1.n140 VDD1.n100 171.744
R2059 VDD1.n141 VDD1.n140 171.744
R2060 VDD1.n141 VDD1.n96 171.744
R2061 VDD1.n148 VDD1.n96 171.744
R2062 VDD1.n149 VDD1.n148 171.744
R2063 VDD1.n149 VDD1.n92 171.744
R2064 VDD1.n156 VDD1.n92 171.744
R2065 VDD1.n157 VDD1.n156 171.744
R2066 VDD1.n157 VDD1.n88 171.744
R2067 VDD1.n164 VDD1.n88 171.744
R2068 VDD1.n165 VDD1.n164 171.744
R2069 VDD1.n31 VDD1.t0 85.8723
R2070 VDD1.n114 VDD1.t1 85.8723
R2071 VDD1.n171 VDD1.n170 68.7728
R2072 VDD1.n173 VDD1.n172 68.4058
R2073 VDD1 VDD1.n84 48.0562
R2074 VDD1.n171 VDD1.n169 47.9427
R2075 VDD1.n173 VDD1.n171 44.0914
R2076 VDD1.n18 VDD1.n16 13.1884
R2077 VDD1.n134 VDD1.n101 13.1884
R2078 VDD1.n54 VDD1.n53 12.8005
R2079 VDD1.n50 VDD1.n49 12.8005
R2080 VDD1.n135 VDD1.n103 12.8005
R2081 VDD1.n139 VDD1.n138 12.8005
R2082 VDD1.n57 VDD1.n14 12.0247
R2083 VDD1.n46 VDD1.n19 12.0247
R2084 VDD1.n130 VDD1.n129 12.0247
R2085 VDD1.n142 VDD1.n99 12.0247
R2086 VDD1.n58 VDD1.n12 11.249
R2087 VDD1.n45 VDD1.n22 11.249
R2088 VDD1.n128 VDD1.n105 11.249
R2089 VDD1.n143 VDD1.n97 11.249
R2090 VDD1.n30 VDD1.n29 10.7239
R2091 VDD1.n113 VDD1.n112 10.7239
R2092 VDD1.n62 VDD1.n61 10.4732
R2093 VDD1.n42 VDD1.n41 10.4732
R2094 VDD1.n125 VDD1.n124 10.4732
R2095 VDD1.n147 VDD1.n146 10.4732
R2096 VDD1.n84 VDD1.n0 9.69747
R2097 VDD1.n65 VDD1.n10 9.69747
R2098 VDD1.n38 VDD1.n24 9.69747
R2099 VDD1.n121 VDD1.n107 9.69747
R2100 VDD1.n150 VDD1.n95 9.69747
R2101 VDD1.n169 VDD1.n85 9.69747
R2102 VDD1.n84 VDD1.n83 9.45567
R2103 VDD1.n169 VDD1.n168 9.45567
R2104 VDD1.n28 VDD1.n27 9.3005
R2105 VDD1.n35 VDD1.n34 9.3005
R2106 VDD1.n37 VDD1.n36 9.3005
R2107 VDD1.n24 VDD1.n23 9.3005
R2108 VDD1.n43 VDD1.n42 9.3005
R2109 VDD1.n45 VDD1.n44 9.3005
R2110 VDD1.n19 VDD1.n17 9.3005
R2111 VDD1.n51 VDD1.n50 9.3005
R2112 VDD1.n77 VDD1.n76 9.3005
R2113 VDD1.n2 VDD1.n1 9.3005
R2114 VDD1.n83 VDD1.n82 9.3005
R2115 VDD1.n75 VDD1.n74 9.3005
R2116 VDD1.n6 VDD1.n5 9.3005
R2117 VDD1.n69 VDD1.n68 9.3005
R2118 VDD1.n67 VDD1.n66 9.3005
R2119 VDD1.n10 VDD1.n9 9.3005
R2120 VDD1.n61 VDD1.n60 9.3005
R2121 VDD1.n59 VDD1.n58 9.3005
R2122 VDD1.n14 VDD1.n13 9.3005
R2123 VDD1.n53 VDD1.n52 9.3005
R2124 VDD1.n160 VDD1.n159 9.3005
R2125 VDD1.n162 VDD1.n161 9.3005
R2126 VDD1.n87 VDD1.n86 9.3005
R2127 VDD1.n168 VDD1.n167 9.3005
R2128 VDD1.n154 VDD1.n153 9.3005
R2129 VDD1.n152 VDD1.n151 9.3005
R2130 VDD1.n95 VDD1.n94 9.3005
R2131 VDD1.n146 VDD1.n145 9.3005
R2132 VDD1.n144 VDD1.n143 9.3005
R2133 VDD1.n99 VDD1.n98 9.3005
R2134 VDD1.n138 VDD1.n137 9.3005
R2135 VDD1.n111 VDD1.n110 9.3005
R2136 VDD1.n118 VDD1.n117 9.3005
R2137 VDD1.n120 VDD1.n119 9.3005
R2138 VDD1.n107 VDD1.n106 9.3005
R2139 VDD1.n126 VDD1.n125 9.3005
R2140 VDD1.n128 VDD1.n127 9.3005
R2141 VDD1.n129 VDD1.n102 9.3005
R2142 VDD1.n136 VDD1.n135 9.3005
R2143 VDD1.n91 VDD1.n90 9.3005
R2144 VDD1.n82 VDD1.n81 8.92171
R2145 VDD1.n66 VDD1.n8 8.92171
R2146 VDD1.n37 VDD1.n26 8.92171
R2147 VDD1.n120 VDD1.n109 8.92171
R2148 VDD1.n151 VDD1.n93 8.92171
R2149 VDD1.n167 VDD1.n166 8.92171
R2150 VDD1.n78 VDD1.n2 8.14595
R2151 VDD1.n70 VDD1.n69 8.14595
R2152 VDD1.n34 VDD1.n33 8.14595
R2153 VDD1.n117 VDD1.n116 8.14595
R2154 VDD1.n155 VDD1.n154 8.14595
R2155 VDD1.n163 VDD1.n87 8.14595
R2156 VDD1.n77 VDD1.n4 7.3702
R2157 VDD1.n73 VDD1.n6 7.3702
R2158 VDD1.n30 VDD1.n28 7.3702
R2159 VDD1.n113 VDD1.n111 7.3702
R2160 VDD1.n158 VDD1.n91 7.3702
R2161 VDD1.n162 VDD1.n89 7.3702
R2162 VDD1.n74 VDD1.n4 6.59444
R2163 VDD1.n74 VDD1.n73 6.59444
R2164 VDD1.n159 VDD1.n158 6.59444
R2165 VDD1.n159 VDD1.n89 6.59444
R2166 VDD1.n78 VDD1.n77 5.81868
R2167 VDD1.n70 VDD1.n6 5.81868
R2168 VDD1.n33 VDD1.n28 5.81868
R2169 VDD1.n116 VDD1.n111 5.81868
R2170 VDD1.n155 VDD1.n91 5.81868
R2171 VDD1.n163 VDD1.n162 5.81868
R2172 VDD1.n81 VDD1.n2 5.04292
R2173 VDD1.n69 VDD1.n8 5.04292
R2174 VDD1.n34 VDD1.n26 5.04292
R2175 VDD1.n117 VDD1.n109 5.04292
R2176 VDD1.n154 VDD1.n93 5.04292
R2177 VDD1.n166 VDD1.n87 5.04292
R2178 VDD1.n82 VDD1.n0 4.26717
R2179 VDD1.n66 VDD1.n65 4.26717
R2180 VDD1.n38 VDD1.n37 4.26717
R2181 VDD1.n121 VDD1.n120 4.26717
R2182 VDD1.n151 VDD1.n150 4.26717
R2183 VDD1.n167 VDD1.n85 4.26717
R2184 VDD1.n62 VDD1.n10 3.49141
R2185 VDD1.n41 VDD1.n24 3.49141
R2186 VDD1.n124 VDD1.n107 3.49141
R2187 VDD1.n147 VDD1.n95 3.49141
R2188 VDD1.n61 VDD1.n12 2.71565
R2189 VDD1.n42 VDD1.n22 2.71565
R2190 VDD1.n125 VDD1.n105 2.71565
R2191 VDD1.n146 VDD1.n97 2.71565
R2192 VDD1.n29 VDD1.n27 2.41282
R2193 VDD1.n112 VDD1.n110 2.41282
R2194 VDD1.n172 VDD1.t5 2.08282
R2195 VDD1.n172 VDD1.t2 2.08282
R2196 VDD1.n170 VDD1.t3 2.08282
R2197 VDD1.n170 VDD1.t4 2.08282
R2198 VDD1.n58 VDD1.n57 1.93989
R2199 VDD1.n46 VDD1.n45 1.93989
R2200 VDD1.n130 VDD1.n128 1.93989
R2201 VDD1.n143 VDD1.n142 1.93989
R2202 VDD1.n54 VDD1.n14 1.16414
R2203 VDD1.n49 VDD1.n19 1.16414
R2204 VDD1.n129 VDD1.n103 1.16414
R2205 VDD1.n139 VDD1.n99 1.16414
R2206 VDD1.n53 VDD1.n16 0.388379
R2207 VDD1.n50 VDD1.n18 0.388379
R2208 VDD1.n135 VDD1.n134 0.388379
R2209 VDD1.n138 VDD1.n101 0.388379
R2210 VDD1 VDD1.n173 0.364724
R2211 VDD1.n83 VDD1.n1 0.155672
R2212 VDD1.n76 VDD1.n1 0.155672
R2213 VDD1.n76 VDD1.n75 0.155672
R2214 VDD1.n75 VDD1.n5 0.155672
R2215 VDD1.n68 VDD1.n5 0.155672
R2216 VDD1.n68 VDD1.n67 0.155672
R2217 VDD1.n67 VDD1.n9 0.155672
R2218 VDD1.n60 VDD1.n9 0.155672
R2219 VDD1.n60 VDD1.n59 0.155672
R2220 VDD1.n59 VDD1.n13 0.155672
R2221 VDD1.n52 VDD1.n13 0.155672
R2222 VDD1.n52 VDD1.n51 0.155672
R2223 VDD1.n51 VDD1.n17 0.155672
R2224 VDD1.n44 VDD1.n17 0.155672
R2225 VDD1.n44 VDD1.n43 0.155672
R2226 VDD1.n43 VDD1.n23 0.155672
R2227 VDD1.n36 VDD1.n23 0.155672
R2228 VDD1.n36 VDD1.n35 0.155672
R2229 VDD1.n35 VDD1.n27 0.155672
R2230 VDD1.n118 VDD1.n110 0.155672
R2231 VDD1.n119 VDD1.n118 0.155672
R2232 VDD1.n119 VDD1.n106 0.155672
R2233 VDD1.n126 VDD1.n106 0.155672
R2234 VDD1.n127 VDD1.n126 0.155672
R2235 VDD1.n127 VDD1.n102 0.155672
R2236 VDD1.n136 VDD1.n102 0.155672
R2237 VDD1.n137 VDD1.n136 0.155672
R2238 VDD1.n137 VDD1.n98 0.155672
R2239 VDD1.n144 VDD1.n98 0.155672
R2240 VDD1.n145 VDD1.n144 0.155672
R2241 VDD1.n145 VDD1.n94 0.155672
R2242 VDD1.n152 VDD1.n94 0.155672
R2243 VDD1.n153 VDD1.n152 0.155672
R2244 VDD1.n153 VDD1.n90 0.155672
R2245 VDD1.n160 VDD1.n90 0.155672
R2246 VDD1.n161 VDD1.n160 0.155672
R2247 VDD1.n161 VDD1.n86 0.155672
R2248 VDD1.n168 VDD1.n86 0.155672
C0 VDD1 VDD2 1.05733f
C1 VDD1 w_n2538_n4090# 2.31111f
C2 VDD1 VTAIL 9.48214f
C3 VDD2 w_n2538_n4090# 2.36506f
C4 VDD1 B 2.10807f
C5 VDD2 VTAIL 9.523809f
C6 w_n2538_n4090# VTAIL 3.44082f
C7 VDD1 VN 0.149481f
C8 VDD1 VP 7.94738f
C9 VDD2 B 2.15898f
C10 w_n2538_n4090# B 9.348821f
C11 VDD2 VN 7.7247f
C12 w_n2538_n4090# VN 4.63176f
C13 B VTAIL 3.99428f
C14 VDD2 VP 0.376637f
C15 w_n2538_n4090# VP 4.957181f
C16 VN VTAIL 7.50863f
C17 VP VTAIL 7.52312f
C18 B VN 1.00437f
C19 B VP 1.54282f
C20 VP VN 6.65007f
C21 VDD2 VSUBS 1.774958f
C22 VDD1 VSUBS 1.577748f
C23 VTAIL VSUBS 1.12442f
C24 VN VSUBS 5.16394f
C25 VP VSUBS 2.308644f
C26 B VSUBS 3.984979f
C27 w_n2538_n4090# VSUBS 0.127215p
C28 VDD1.n0 VSUBS 0.030727f
C29 VDD1.n1 VSUBS 0.027126f
C30 VDD1.n2 VSUBS 0.014576f
C31 VDD1.n3 VSUBS 0.034453f
C32 VDD1.n4 VSUBS 0.015434f
C33 VDD1.n5 VSUBS 0.027126f
C34 VDD1.n6 VSUBS 0.014576f
C35 VDD1.n7 VSUBS 0.034453f
C36 VDD1.n8 VSUBS 0.015434f
C37 VDD1.n9 VSUBS 0.027126f
C38 VDD1.n10 VSUBS 0.014576f
C39 VDD1.n11 VSUBS 0.034453f
C40 VDD1.n12 VSUBS 0.015434f
C41 VDD1.n13 VSUBS 0.027126f
C42 VDD1.n14 VSUBS 0.014576f
C43 VDD1.n15 VSUBS 0.034453f
C44 VDD1.n16 VSUBS 0.015005f
C45 VDD1.n17 VSUBS 0.027126f
C46 VDD1.n18 VSUBS 0.015005f
C47 VDD1.n19 VSUBS 0.014576f
C48 VDD1.n20 VSUBS 0.034453f
C49 VDD1.n21 VSUBS 0.034453f
C50 VDD1.n22 VSUBS 0.015434f
C51 VDD1.n23 VSUBS 0.027126f
C52 VDD1.n24 VSUBS 0.014576f
C53 VDD1.n25 VSUBS 0.034453f
C54 VDD1.n26 VSUBS 0.015434f
C55 VDD1.n27 VSUBS 1.76187f
C56 VDD1.n28 VSUBS 0.014576f
C57 VDD1.t0 VSUBS 0.074571f
C58 VDD1.n29 VSUBS 0.25791f
C59 VDD1.n30 VSUBS 0.025918f
C60 VDD1.n31 VSUBS 0.02584f
C61 VDD1.n32 VSUBS 0.034453f
C62 VDD1.n33 VSUBS 0.015434f
C63 VDD1.n34 VSUBS 0.014576f
C64 VDD1.n35 VSUBS 0.027126f
C65 VDD1.n36 VSUBS 0.027126f
C66 VDD1.n37 VSUBS 0.014576f
C67 VDD1.n38 VSUBS 0.015434f
C68 VDD1.n39 VSUBS 0.034453f
C69 VDD1.n40 VSUBS 0.034453f
C70 VDD1.n41 VSUBS 0.015434f
C71 VDD1.n42 VSUBS 0.014576f
C72 VDD1.n43 VSUBS 0.027126f
C73 VDD1.n44 VSUBS 0.027126f
C74 VDD1.n45 VSUBS 0.014576f
C75 VDD1.n46 VSUBS 0.015434f
C76 VDD1.n47 VSUBS 0.034453f
C77 VDD1.n48 VSUBS 0.034453f
C78 VDD1.n49 VSUBS 0.015434f
C79 VDD1.n50 VSUBS 0.014576f
C80 VDD1.n51 VSUBS 0.027126f
C81 VDD1.n52 VSUBS 0.027126f
C82 VDD1.n53 VSUBS 0.014576f
C83 VDD1.n54 VSUBS 0.015434f
C84 VDD1.n55 VSUBS 0.034453f
C85 VDD1.n56 VSUBS 0.034453f
C86 VDD1.n57 VSUBS 0.015434f
C87 VDD1.n58 VSUBS 0.014576f
C88 VDD1.n59 VSUBS 0.027126f
C89 VDD1.n60 VSUBS 0.027126f
C90 VDD1.n61 VSUBS 0.014576f
C91 VDD1.n62 VSUBS 0.015434f
C92 VDD1.n63 VSUBS 0.034453f
C93 VDD1.n64 VSUBS 0.034453f
C94 VDD1.n65 VSUBS 0.015434f
C95 VDD1.n66 VSUBS 0.014576f
C96 VDD1.n67 VSUBS 0.027126f
C97 VDD1.n68 VSUBS 0.027126f
C98 VDD1.n69 VSUBS 0.014576f
C99 VDD1.n70 VSUBS 0.015434f
C100 VDD1.n71 VSUBS 0.034453f
C101 VDD1.n72 VSUBS 0.034453f
C102 VDD1.n73 VSUBS 0.015434f
C103 VDD1.n74 VSUBS 0.014576f
C104 VDD1.n75 VSUBS 0.027126f
C105 VDD1.n76 VSUBS 0.027126f
C106 VDD1.n77 VSUBS 0.014576f
C107 VDD1.n78 VSUBS 0.015434f
C108 VDD1.n79 VSUBS 0.034453f
C109 VDD1.n80 VSUBS 0.086547f
C110 VDD1.n81 VSUBS 0.015434f
C111 VDD1.n82 VSUBS 0.014576f
C112 VDD1.n83 VSUBS 0.058625f
C113 VDD1.n84 VSUBS 0.06687f
C114 VDD1.n85 VSUBS 0.030727f
C115 VDD1.n86 VSUBS 0.027126f
C116 VDD1.n87 VSUBS 0.014576f
C117 VDD1.n88 VSUBS 0.034453f
C118 VDD1.n89 VSUBS 0.015434f
C119 VDD1.n90 VSUBS 0.027126f
C120 VDD1.n91 VSUBS 0.014576f
C121 VDD1.n92 VSUBS 0.034453f
C122 VDD1.n93 VSUBS 0.015434f
C123 VDD1.n94 VSUBS 0.027126f
C124 VDD1.n95 VSUBS 0.014576f
C125 VDD1.n96 VSUBS 0.034453f
C126 VDD1.n97 VSUBS 0.015434f
C127 VDD1.n98 VSUBS 0.027126f
C128 VDD1.n99 VSUBS 0.014576f
C129 VDD1.n100 VSUBS 0.034453f
C130 VDD1.n101 VSUBS 0.015005f
C131 VDD1.n102 VSUBS 0.027126f
C132 VDD1.n103 VSUBS 0.015434f
C133 VDD1.n104 VSUBS 0.034453f
C134 VDD1.n105 VSUBS 0.015434f
C135 VDD1.n106 VSUBS 0.027126f
C136 VDD1.n107 VSUBS 0.014576f
C137 VDD1.n108 VSUBS 0.034453f
C138 VDD1.n109 VSUBS 0.015434f
C139 VDD1.n110 VSUBS 1.76187f
C140 VDD1.n111 VSUBS 0.014576f
C141 VDD1.t1 VSUBS 0.074571f
C142 VDD1.n112 VSUBS 0.25791f
C143 VDD1.n113 VSUBS 0.025918f
C144 VDD1.n114 VSUBS 0.02584f
C145 VDD1.n115 VSUBS 0.034453f
C146 VDD1.n116 VSUBS 0.015434f
C147 VDD1.n117 VSUBS 0.014576f
C148 VDD1.n118 VSUBS 0.027126f
C149 VDD1.n119 VSUBS 0.027126f
C150 VDD1.n120 VSUBS 0.014576f
C151 VDD1.n121 VSUBS 0.015434f
C152 VDD1.n122 VSUBS 0.034453f
C153 VDD1.n123 VSUBS 0.034453f
C154 VDD1.n124 VSUBS 0.015434f
C155 VDD1.n125 VSUBS 0.014576f
C156 VDD1.n126 VSUBS 0.027126f
C157 VDD1.n127 VSUBS 0.027126f
C158 VDD1.n128 VSUBS 0.014576f
C159 VDD1.n129 VSUBS 0.014576f
C160 VDD1.n130 VSUBS 0.015434f
C161 VDD1.n131 VSUBS 0.034453f
C162 VDD1.n132 VSUBS 0.034453f
C163 VDD1.n133 VSUBS 0.034453f
C164 VDD1.n134 VSUBS 0.015005f
C165 VDD1.n135 VSUBS 0.014576f
C166 VDD1.n136 VSUBS 0.027126f
C167 VDD1.n137 VSUBS 0.027126f
C168 VDD1.n138 VSUBS 0.014576f
C169 VDD1.n139 VSUBS 0.015434f
C170 VDD1.n140 VSUBS 0.034453f
C171 VDD1.n141 VSUBS 0.034453f
C172 VDD1.n142 VSUBS 0.015434f
C173 VDD1.n143 VSUBS 0.014576f
C174 VDD1.n144 VSUBS 0.027126f
C175 VDD1.n145 VSUBS 0.027126f
C176 VDD1.n146 VSUBS 0.014576f
C177 VDD1.n147 VSUBS 0.015434f
C178 VDD1.n148 VSUBS 0.034453f
C179 VDD1.n149 VSUBS 0.034453f
C180 VDD1.n150 VSUBS 0.015434f
C181 VDD1.n151 VSUBS 0.014576f
C182 VDD1.n152 VSUBS 0.027126f
C183 VDD1.n153 VSUBS 0.027126f
C184 VDD1.n154 VSUBS 0.014576f
C185 VDD1.n155 VSUBS 0.015434f
C186 VDD1.n156 VSUBS 0.034453f
C187 VDD1.n157 VSUBS 0.034453f
C188 VDD1.n158 VSUBS 0.015434f
C189 VDD1.n159 VSUBS 0.014576f
C190 VDD1.n160 VSUBS 0.027126f
C191 VDD1.n161 VSUBS 0.027126f
C192 VDD1.n162 VSUBS 0.014576f
C193 VDD1.n163 VSUBS 0.015434f
C194 VDD1.n164 VSUBS 0.034453f
C195 VDD1.n165 VSUBS 0.086547f
C196 VDD1.n166 VSUBS 0.015434f
C197 VDD1.n167 VSUBS 0.014576f
C198 VDD1.n168 VSUBS 0.058625f
C199 VDD1.n169 VSUBS 0.066251f
C200 VDD1.t3 VSUBS 0.334615f
C201 VDD1.t4 VSUBS 0.334615f
C202 VDD1.n170 VSUBS 2.7122f
C203 VDD1.n171 VSUBS 3.11917f
C204 VDD1.t5 VSUBS 0.334615f
C205 VDD1.t2 VSUBS 0.334615f
C206 VDD1.n172 VSUBS 2.70828f
C207 VDD1.n173 VSUBS 3.3514f
C208 VP.n0 VSUBS 0.037658f
C209 VP.t1 VSUBS 2.62796f
C210 VP.n1 VSUBS 0.052876f
C211 VP.n2 VSUBS 0.037658f
C212 VP.t2 VSUBS 2.62796f
C213 VP.n3 VSUBS 0.057073f
C214 VP.n4 VSUBS 0.037658f
C215 VP.t3 VSUBS 2.62796f
C216 VP.n5 VSUBS 0.052876f
C217 VP.t5 VSUBS 2.76707f
C218 VP.n6 VSUBS 1.01961f
C219 VP.t0 VSUBS 2.62796f
C220 VP.n7 VSUBS 1.00402f
C221 VP.n8 VSUBS 0.05286f
C222 VP.n9 VSUBS 0.242137f
C223 VP.n10 VSUBS 0.037658f
C224 VP.n11 VSUBS 0.037658f
C225 VP.n12 VSUBS 0.057073f
C226 VP.n13 VSUBS 0.050088f
C227 VP.n14 VSUBS 1.01592f
C228 VP.n15 VSUBS 1.90523f
C229 VP.n16 VSUBS 1.93368f
C230 VP.t4 VSUBS 2.62796f
C231 VP.n17 VSUBS 1.01592f
C232 VP.n18 VSUBS 0.050088f
C233 VP.n19 VSUBS 0.037658f
C234 VP.n20 VSUBS 0.037658f
C235 VP.n21 VSUBS 0.037658f
C236 VP.n22 VSUBS 0.052876f
C237 VP.n23 VSUBS 0.05286f
C238 VP.n24 VSUBS 0.929752f
C239 VP.n25 VSUBS 0.05286f
C240 VP.n26 VSUBS 0.037658f
C241 VP.n27 VSUBS 0.037658f
C242 VP.n28 VSUBS 0.037658f
C243 VP.n29 VSUBS 0.057073f
C244 VP.n30 VSUBS 0.050088f
C245 VP.n31 VSUBS 1.01592f
C246 VP.n32 VSUBS 0.036765f
C247 B.n0 VSUBS 0.005176f
C248 B.n1 VSUBS 0.005176f
C249 B.n2 VSUBS 0.008185f
C250 B.n3 VSUBS 0.008185f
C251 B.n4 VSUBS 0.008185f
C252 B.n5 VSUBS 0.008185f
C253 B.n6 VSUBS 0.008185f
C254 B.n7 VSUBS 0.008185f
C255 B.n8 VSUBS 0.008185f
C256 B.n9 VSUBS 0.008185f
C257 B.n10 VSUBS 0.008185f
C258 B.n11 VSUBS 0.008185f
C259 B.n12 VSUBS 0.008185f
C260 B.n13 VSUBS 0.008185f
C261 B.n14 VSUBS 0.008185f
C262 B.n15 VSUBS 0.008185f
C263 B.n16 VSUBS 0.008185f
C264 B.n17 VSUBS 0.019314f
C265 B.n18 VSUBS 0.008185f
C266 B.n19 VSUBS 0.008185f
C267 B.n20 VSUBS 0.008185f
C268 B.n21 VSUBS 0.008185f
C269 B.n22 VSUBS 0.008185f
C270 B.n23 VSUBS 0.008185f
C271 B.n24 VSUBS 0.008185f
C272 B.n25 VSUBS 0.008185f
C273 B.n26 VSUBS 0.008185f
C274 B.n27 VSUBS 0.008185f
C275 B.n28 VSUBS 0.008185f
C276 B.n29 VSUBS 0.008185f
C277 B.n30 VSUBS 0.008185f
C278 B.n31 VSUBS 0.008185f
C279 B.n32 VSUBS 0.008185f
C280 B.n33 VSUBS 0.008185f
C281 B.n34 VSUBS 0.008185f
C282 B.n35 VSUBS 0.008185f
C283 B.n36 VSUBS 0.008185f
C284 B.n37 VSUBS 0.008185f
C285 B.n38 VSUBS 0.008185f
C286 B.n39 VSUBS 0.008185f
C287 B.n40 VSUBS 0.008185f
C288 B.n41 VSUBS 0.008185f
C289 B.n42 VSUBS 0.008185f
C290 B.n43 VSUBS 0.008185f
C291 B.t5 VSUBS 0.343968f
C292 B.t4 VSUBS 0.370441f
C293 B.t3 VSUBS 1.286f
C294 B.n44 VSUBS 0.540412f
C295 B.n45 VSUBS 0.345171f
C296 B.n46 VSUBS 0.008185f
C297 B.n47 VSUBS 0.008185f
C298 B.n48 VSUBS 0.008185f
C299 B.n49 VSUBS 0.008185f
C300 B.n50 VSUBS 0.004574f
C301 B.n51 VSUBS 0.008185f
C302 B.t8 VSUBS 0.343972f
C303 B.t7 VSUBS 0.370445f
C304 B.t6 VSUBS 1.286f
C305 B.n52 VSUBS 0.540409f
C306 B.n53 VSUBS 0.345167f
C307 B.n54 VSUBS 0.018964f
C308 B.n55 VSUBS 0.008185f
C309 B.n56 VSUBS 0.008185f
C310 B.n57 VSUBS 0.008185f
C311 B.n58 VSUBS 0.008185f
C312 B.n59 VSUBS 0.008185f
C313 B.n60 VSUBS 0.008185f
C314 B.n61 VSUBS 0.008185f
C315 B.n62 VSUBS 0.008185f
C316 B.n63 VSUBS 0.008185f
C317 B.n64 VSUBS 0.008185f
C318 B.n65 VSUBS 0.008185f
C319 B.n66 VSUBS 0.008185f
C320 B.n67 VSUBS 0.008185f
C321 B.n68 VSUBS 0.008185f
C322 B.n69 VSUBS 0.008185f
C323 B.n70 VSUBS 0.008185f
C324 B.n71 VSUBS 0.008185f
C325 B.n72 VSUBS 0.008185f
C326 B.n73 VSUBS 0.008185f
C327 B.n74 VSUBS 0.008185f
C328 B.n75 VSUBS 0.008185f
C329 B.n76 VSUBS 0.008185f
C330 B.n77 VSUBS 0.008185f
C331 B.n78 VSUBS 0.008185f
C332 B.n79 VSUBS 0.019492f
C333 B.n80 VSUBS 0.008185f
C334 B.n81 VSUBS 0.008185f
C335 B.n82 VSUBS 0.008185f
C336 B.n83 VSUBS 0.008185f
C337 B.n84 VSUBS 0.008185f
C338 B.n85 VSUBS 0.008185f
C339 B.n86 VSUBS 0.008185f
C340 B.n87 VSUBS 0.008185f
C341 B.n88 VSUBS 0.008185f
C342 B.n89 VSUBS 0.008185f
C343 B.n90 VSUBS 0.008185f
C344 B.n91 VSUBS 0.008185f
C345 B.n92 VSUBS 0.008185f
C346 B.n93 VSUBS 0.008185f
C347 B.n94 VSUBS 0.008185f
C348 B.n95 VSUBS 0.008185f
C349 B.n96 VSUBS 0.008185f
C350 B.n97 VSUBS 0.008185f
C351 B.n98 VSUBS 0.008185f
C352 B.n99 VSUBS 0.008185f
C353 B.n100 VSUBS 0.008185f
C354 B.n101 VSUBS 0.008185f
C355 B.n102 VSUBS 0.008185f
C356 B.n103 VSUBS 0.008185f
C357 B.n104 VSUBS 0.008185f
C358 B.n105 VSUBS 0.008185f
C359 B.n106 VSUBS 0.008185f
C360 B.n107 VSUBS 0.008185f
C361 B.n108 VSUBS 0.008185f
C362 B.n109 VSUBS 0.008185f
C363 B.n110 VSUBS 0.008185f
C364 B.n111 VSUBS 0.020408f
C365 B.n112 VSUBS 0.008185f
C366 B.n113 VSUBS 0.008185f
C367 B.n114 VSUBS 0.008185f
C368 B.n115 VSUBS 0.008185f
C369 B.n116 VSUBS 0.008185f
C370 B.n117 VSUBS 0.008185f
C371 B.n118 VSUBS 0.008185f
C372 B.n119 VSUBS 0.008185f
C373 B.n120 VSUBS 0.008185f
C374 B.n121 VSUBS 0.008185f
C375 B.n122 VSUBS 0.008185f
C376 B.n123 VSUBS 0.008185f
C377 B.n124 VSUBS 0.008185f
C378 B.n125 VSUBS 0.008185f
C379 B.n126 VSUBS 0.008185f
C380 B.n127 VSUBS 0.008185f
C381 B.n128 VSUBS 0.008185f
C382 B.n129 VSUBS 0.008185f
C383 B.n130 VSUBS 0.008185f
C384 B.n131 VSUBS 0.008185f
C385 B.n132 VSUBS 0.008185f
C386 B.n133 VSUBS 0.008185f
C387 B.n134 VSUBS 0.008185f
C388 B.n135 VSUBS 0.008185f
C389 B.n136 VSUBS 0.008185f
C390 B.t1 VSUBS 0.343972f
C391 B.t2 VSUBS 0.370445f
C392 B.t0 VSUBS 1.286f
C393 B.n137 VSUBS 0.540409f
C394 B.n138 VSUBS 0.345167f
C395 B.n139 VSUBS 0.018964f
C396 B.n140 VSUBS 0.008185f
C397 B.n141 VSUBS 0.008185f
C398 B.n142 VSUBS 0.008185f
C399 B.n143 VSUBS 0.008185f
C400 B.n144 VSUBS 0.008185f
C401 B.t10 VSUBS 0.343968f
C402 B.t11 VSUBS 0.370441f
C403 B.t9 VSUBS 1.286f
C404 B.n145 VSUBS 0.540412f
C405 B.n146 VSUBS 0.345171f
C406 B.n147 VSUBS 0.008185f
C407 B.n148 VSUBS 0.008185f
C408 B.n149 VSUBS 0.008185f
C409 B.n150 VSUBS 0.008185f
C410 B.n151 VSUBS 0.008185f
C411 B.n152 VSUBS 0.008185f
C412 B.n153 VSUBS 0.008185f
C413 B.n154 VSUBS 0.008185f
C414 B.n155 VSUBS 0.008185f
C415 B.n156 VSUBS 0.008185f
C416 B.n157 VSUBS 0.008185f
C417 B.n158 VSUBS 0.008185f
C418 B.n159 VSUBS 0.008185f
C419 B.n160 VSUBS 0.008185f
C420 B.n161 VSUBS 0.008185f
C421 B.n162 VSUBS 0.008185f
C422 B.n163 VSUBS 0.008185f
C423 B.n164 VSUBS 0.008185f
C424 B.n165 VSUBS 0.008185f
C425 B.n166 VSUBS 0.008185f
C426 B.n167 VSUBS 0.008185f
C427 B.n168 VSUBS 0.008185f
C428 B.n169 VSUBS 0.008185f
C429 B.n170 VSUBS 0.008185f
C430 B.n171 VSUBS 0.008185f
C431 B.n172 VSUBS 0.020408f
C432 B.n173 VSUBS 0.008185f
C433 B.n174 VSUBS 0.008185f
C434 B.n175 VSUBS 0.008185f
C435 B.n176 VSUBS 0.008185f
C436 B.n177 VSUBS 0.008185f
C437 B.n178 VSUBS 0.008185f
C438 B.n179 VSUBS 0.008185f
C439 B.n180 VSUBS 0.008185f
C440 B.n181 VSUBS 0.008185f
C441 B.n182 VSUBS 0.008185f
C442 B.n183 VSUBS 0.008185f
C443 B.n184 VSUBS 0.008185f
C444 B.n185 VSUBS 0.008185f
C445 B.n186 VSUBS 0.008185f
C446 B.n187 VSUBS 0.008185f
C447 B.n188 VSUBS 0.008185f
C448 B.n189 VSUBS 0.008185f
C449 B.n190 VSUBS 0.008185f
C450 B.n191 VSUBS 0.008185f
C451 B.n192 VSUBS 0.008185f
C452 B.n193 VSUBS 0.008185f
C453 B.n194 VSUBS 0.008185f
C454 B.n195 VSUBS 0.008185f
C455 B.n196 VSUBS 0.008185f
C456 B.n197 VSUBS 0.008185f
C457 B.n198 VSUBS 0.008185f
C458 B.n199 VSUBS 0.008185f
C459 B.n200 VSUBS 0.008185f
C460 B.n201 VSUBS 0.008185f
C461 B.n202 VSUBS 0.008185f
C462 B.n203 VSUBS 0.008185f
C463 B.n204 VSUBS 0.008185f
C464 B.n205 VSUBS 0.008185f
C465 B.n206 VSUBS 0.008185f
C466 B.n207 VSUBS 0.008185f
C467 B.n208 VSUBS 0.008185f
C468 B.n209 VSUBS 0.008185f
C469 B.n210 VSUBS 0.008185f
C470 B.n211 VSUBS 0.008185f
C471 B.n212 VSUBS 0.008185f
C472 B.n213 VSUBS 0.008185f
C473 B.n214 VSUBS 0.008185f
C474 B.n215 VSUBS 0.008185f
C475 B.n216 VSUBS 0.008185f
C476 B.n217 VSUBS 0.008185f
C477 B.n218 VSUBS 0.008185f
C478 B.n219 VSUBS 0.008185f
C479 B.n220 VSUBS 0.008185f
C480 B.n221 VSUBS 0.008185f
C481 B.n222 VSUBS 0.008185f
C482 B.n223 VSUBS 0.008185f
C483 B.n224 VSUBS 0.008185f
C484 B.n225 VSUBS 0.008185f
C485 B.n226 VSUBS 0.008185f
C486 B.n227 VSUBS 0.008185f
C487 B.n228 VSUBS 0.008185f
C488 B.n229 VSUBS 0.008185f
C489 B.n230 VSUBS 0.008185f
C490 B.n231 VSUBS 0.019314f
C491 B.n232 VSUBS 0.019314f
C492 B.n233 VSUBS 0.020408f
C493 B.n234 VSUBS 0.008185f
C494 B.n235 VSUBS 0.008185f
C495 B.n236 VSUBS 0.008185f
C496 B.n237 VSUBS 0.008185f
C497 B.n238 VSUBS 0.008185f
C498 B.n239 VSUBS 0.008185f
C499 B.n240 VSUBS 0.008185f
C500 B.n241 VSUBS 0.008185f
C501 B.n242 VSUBS 0.008185f
C502 B.n243 VSUBS 0.008185f
C503 B.n244 VSUBS 0.008185f
C504 B.n245 VSUBS 0.008185f
C505 B.n246 VSUBS 0.008185f
C506 B.n247 VSUBS 0.008185f
C507 B.n248 VSUBS 0.008185f
C508 B.n249 VSUBS 0.008185f
C509 B.n250 VSUBS 0.008185f
C510 B.n251 VSUBS 0.008185f
C511 B.n252 VSUBS 0.008185f
C512 B.n253 VSUBS 0.008185f
C513 B.n254 VSUBS 0.008185f
C514 B.n255 VSUBS 0.008185f
C515 B.n256 VSUBS 0.008185f
C516 B.n257 VSUBS 0.008185f
C517 B.n258 VSUBS 0.008185f
C518 B.n259 VSUBS 0.008185f
C519 B.n260 VSUBS 0.008185f
C520 B.n261 VSUBS 0.008185f
C521 B.n262 VSUBS 0.008185f
C522 B.n263 VSUBS 0.008185f
C523 B.n264 VSUBS 0.008185f
C524 B.n265 VSUBS 0.008185f
C525 B.n266 VSUBS 0.008185f
C526 B.n267 VSUBS 0.008185f
C527 B.n268 VSUBS 0.008185f
C528 B.n269 VSUBS 0.008185f
C529 B.n270 VSUBS 0.008185f
C530 B.n271 VSUBS 0.008185f
C531 B.n272 VSUBS 0.008185f
C532 B.n273 VSUBS 0.008185f
C533 B.n274 VSUBS 0.008185f
C534 B.n275 VSUBS 0.008185f
C535 B.n276 VSUBS 0.008185f
C536 B.n277 VSUBS 0.008185f
C537 B.n278 VSUBS 0.008185f
C538 B.n279 VSUBS 0.008185f
C539 B.n280 VSUBS 0.008185f
C540 B.n281 VSUBS 0.008185f
C541 B.n282 VSUBS 0.008185f
C542 B.n283 VSUBS 0.008185f
C543 B.n284 VSUBS 0.008185f
C544 B.n285 VSUBS 0.008185f
C545 B.n286 VSUBS 0.008185f
C546 B.n287 VSUBS 0.008185f
C547 B.n288 VSUBS 0.008185f
C548 B.n289 VSUBS 0.008185f
C549 B.n290 VSUBS 0.008185f
C550 B.n291 VSUBS 0.008185f
C551 B.n292 VSUBS 0.008185f
C552 B.n293 VSUBS 0.008185f
C553 B.n294 VSUBS 0.008185f
C554 B.n295 VSUBS 0.008185f
C555 B.n296 VSUBS 0.008185f
C556 B.n297 VSUBS 0.008185f
C557 B.n298 VSUBS 0.008185f
C558 B.n299 VSUBS 0.008185f
C559 B.n300 VSUBS 0.008185f
C560 B.n301 VSUBS 0.008185f
C561 B.n302 VSUBS 0.008185f
C562 B.n303 VSUBS 0.008185f
C563 B.n304 VSUBS 0.008185f
C564 B.n305 VSUBS 0.008185f
C565 B.n306 VSUBS 0.008185f
C566 B.n307 VSUBS 0.008185f
C567 B.n308 VSUBS 0.008185f
C568 B.n309 VSUBS 0.008185f
C569 B.n310 VSUBS 0.007704f
C570 B.n311 VSUBS 0.018964f
C571 B.n312 VSUBS 0.004574f
C572 B.n313 VSUBS 0.008185f
C573 B.n314 VSUBS 0.008185f
C574 B.n315 VSUBS 0.008185f
C575 B.n316 VSUBS 0.008185f
C576 B.n317 VSUBS 0.008185f
C577 B.n318 VSUBS 0.008185f
C578 B.n319 VSUBS 0.008185f
C579 B.n320 VSUBS 0.008185f
C580 B.n321 VSUBS 0.008185f
C581 B.n322 VSUBS 0.008185f
C582 B.n323 VSUBS 0.008185f
C583 B.n324 VSUBS 0.008185f
C584 B.n325 VSUBS 0.004574f
C585 B.n326 VSUBS 0.008185f
C586 B.n327 VSUBS 0.008185f
C587 B.n328 VSUBS 0.007704f
C588 B.n329 VSUBS 0.008185f
C589 B.n330 VSUBS 0.008185f
C590 B.n331 VSUBS 0.008185f
C591 B.n332 VSUBS 0.008185f
C592 B.n333 VSUBS 0.008185f
C593 B.n334 VSUBS 0.008185f
C594 B.n335 VSUBS 0.008185f
C595 B.n336 VSUBS 0.008185f
C596 B.n337 VSUBS 0.008185f
C597 B.n338 VSUBS 0.008185f
C598 B.n339 VSUBS 0.008185f
C599 B.n340 VSUBS 0.008185f
C600 B.n341 VSUBS 0.008185f
C601 B.n342 VSUBS 0.008185f
C602 B.n343 VSUBS 0.008185f
C603 B.n344 VSUBS 0.008185f
C604 B.n345 VSUBS 0.008185f
C605 B.n346 VSUBS 0.008185f
C606 B.n347 VSUBS 0.008185f
C607 B.n348 VSUBS 0.008185f
C608 B.n349 VSUBS 0.008185f
C609 B.n350 VSUBS 0.008185f
C610 B.n351 VSUBS 0.008185f
C611 B.n352 VSUBS 0.008185f
C612 B.n353 VSUBS 0.008185f
C613 B.n354 VSUBS 0.008185f
C614 B.n355 VSUBS 0.008185f
C615 B.n356 VSUBS 0.008185f
C616 B.n357 VSUBS 0.008185f
C617 B.n358 VSUBS 0.008185f
C618 B.n359 VSUBS 0.008185f
C619 B.n360 VSUBS 0.008185f
C620 B.n361 VSUBS 0.008185f
C621 B.n362 VSUBS 0.008185f
C622 B.n363 VSUBS 0.008185f
C623 B.n364 VSUBS 0.008185f
C624 B.n365 VSUBS 0.008185f
C625 B.n366 VSUBS 0.008185f
C626 B.n367 VSUBS 0.008185f
C627 B.n368 VSUBS 0.008185f
C628 B.n369 VSUBS 0.008185f
C629 B.n370 VSUBS 0.008185f
C630 B.n371 VSUBS 0.008185f
C631 B.n372 VSUBS 0.008185f
C632 B.n373 VSUBS 0.008185f
C633 B.n374 VSUBS 0.008185f
C634 B.n375 VSUBS 0.008185f
C635 B.n376 VSUBS 0.008185f
C636 B.n377 VSUBS 0.008185f
C637 B.n378 VSUBS 0.008185f
C638 B.n379 VSUBS 0.008185f
C639 B.n380 VSUBS 0.008185f
C640 B.n381 VSUBS 0.008185f
C641 B.n382 VSUBS 0.008185f
C642 B.n383 VSUBS 0.008185f
C643 B.n384 VSUBS 0.008185f
C644 B.n385 VSUBS 0.008185f
C645 B.n386 VSUBS 0.008185f
C646 B.n387 VSUBS 0.008185f
C647 B.n388 VSUBS 0.008185f
C648 B.n389 VSUBS 0.008185f
C649 B.n390 VSUBS 0.008185f
C650 B.n391 VSUBS 0.008185f
C651 B.n392 VSUBS 0.008185f
C652 B.n393 VSUBS 0.008185f
C653 B.n394 VSUBS 0.008185f
C654 B.n395 VSUBS 0.008185f
C655 B.n396 VSUBS 0.008185f
C656 B.n397 VSUBS 0.008185f
C657 B.n398 VSUBS 0.008185f
C658 B.n399 VSUBS 0.008185f
C659 B.n400 VSUBS 0.008185f
C660 B.n401 VSUBS 0.008185f
C661 B.n402 VSUBS 0.008185f
C662 B.n403 VSUBS 0.008185f
C663 B.n404 VSUBS 0.020408f
C664 B.n405 VSUBS 0.019314f
C665 B.n406 VSUBS 0.019314f
C666 B.n407 VSUBS 0.008185f
C667 B.n408 VSUBS 0.008185f
C668 B.n409 VSUBS 0.008185f
C669 B.n410 VSUBS 0.008185f
C670 B.n411 VSUBS 0.008185f
C671 B.n412 VSUBS 0.008185f
C672 B.n413 VSUBS 0.008185f
C673 B.n414 VSUBS 0.008185f
C674 B.n415 VSUBS 0.008185f
C675 B.n416 VSUBS 0.008185f
C676 B.n417 VSUBS 0.008185f
C677 B.n418 VSUBS 0.008185f
C678 B.n419 VSUBS 0.008185f
C679 B.n420 VSUBS 0.008185f
C680 B.n421 VSUBS 0.008185f
C681 B.n422 VSUBS 0.008185f
C682 B.n423 VSUBS 0.008185f
C683 B.n424 VSUBS 0.008185f
C684 B.n425 VSUBS 0.008185f
C685 B.n426 VSUBS 0.008185f
C686 B.n427 VSUBS 0.008185f
C687 B.n428 VSUBS 0.008185f
C688 B.n429 VSUBS 0.008185f
C689 B.n430 VSUBS 0.008185f
C690 B.n431 VSUBS 0.008185f
C691 B.n432 VSUBS 0.008185f
C692 B.n433 VSUBS 0.008185f
C693 B.n434 VSUBS 0.008185f
C694 B.n435 VSUBS 0.008185f
C695 B.n436 VSUBS 0.008185f
C696 B.n437 VSUBS 0.008185f
C697 B.n438 VSUBS 0.008185f
C698 B.n439 VSUBS 0.008185f
C699 B.n440 VSUBS 0.008185f
C700 B.n441 VSUBS 0.008185f
C701 B.n442 VSUBS 0.008185f
C702 B.n443 VSUBS 0.008185f
C703 B.n444 VSUBS 0.008185f
C704 B.n445 VSUBS 0.008185f
C705 B.n446 VSUBS 0.008185f
C706 B.n447 VSUBS 0.008185f
C707 B.n448 VSUBS 0.008185f
C708 B.n449 VSUBS 0.008185f
C709 B.n450 VSUBS 0.008185f
C710 B.n451 VSUBS 0.008185f
C711 B.n452 VSUBS 0.008185f
C712 B.n453 VSUBS 0.008185f
C713 B.n454 VSUBS 0.008185f
C714 B.n455 VSUBS 0.008185f
C715 B.n456 VSUBS 0.008185f
C716 B.n457 VSUBS 0.008185f
C717 B.n458 VSUBS 0.008185f
C718 B.n459 VSUBS 0.008185f
C719 B.n460 VSUBS 0.008185f
C720 B.n461 VSUBS 0.008185f
C721 B.n462 VSUBS 0.008185f
C722 B.n463 VSUBS 0.008185f
C723 B.n464 VSUBS 0.008185f
C724 B.n465 VSUBS 0.008185f
C725 B.n466 VSUBS 0.008185f
C726 B.n467 VSUBS 0.008185f
C727 B.n468 VSUBS 0.008185f
C728 B.n469 VSUBS 0.008185f
C729 B.n470 VSUBS 0.008185f
C730 B.n471 VSUBS 0.008185f
C731 B.n472 VSUBS 0.008185f
C732 B.n473 VSUBS 0.008185f
C733 B.n474 VSUBS 0.008185f
C734 B.n475 VSUBS 0.008185f
C735 B.n476 VSUBS 0.008185f
C736 B.n477 VSUBS 0.008185f
C737 B.n478 VSUBS 0.008185f
C738 B.n479 VSUBS 0.008185f
C739 B.n480 VSUBS 0.008185f
C740 B.n481 VSUBS 0.008185f
C741 B.n482 VSUBS 0.008185f
C742 B.n483 VSUBS 0.008185f
C743 B.n484 VSUBS 0.008185f
C744 B.n485 VSUBS 0.008185f
C745 B.n486 VSUBS 0.008185f
C746 B.n487 VSUBS 0.008185f
C747 B.n488 VSUBS 0.008185f
C748 B.n489 VSUBS 0.008185f
C749 B.n490 VSUBS 0.008185f
C750 B.n491 VSUBS 0.008185f
C751 B.n492 VSUBS 0.008185f
C752 B.n493 VSUBS 0.008185f
C753 B.n494 VSUBS 0.008185f
C754 B.n495 VSUBS 0.008185f
C755 B.n496 VSUBS 0.008185f
C756 B.n497 VSUBS 0.008185f
C757 B.n498 VSUBS 0.020229f
C758 B.n499 VSUBS 0.019314f
C759 B.n500 VSUBS 0.020408f
C760 B.n501 VSUBS 0.008185f
C761 B.n502 VSUBS 0.008185f
C762 B.n503 VSUBS 0.008185f
C763 B.n504 VSUBS 0.008185f
C764 B.n505 VSUBS 0.008185f
C765 B.n506 VSUBS 0.008185f
C766 B.n507 VSUBS 0.008185f
C767 B.n508 VSUBS 0.008185f
C768 B.n509 VSUBS 0.008185f
C769 B.n510 VSUBS 0.008185f
C770 B.n511 VSUBS 0.008185f
C771 B.n512 VSUBS 0.008185f
C772 B.n513 VSUBS 0.008185f
C773 B.n514 VSUBS 0.008185f
C774 B.n515 VSUBS 0.008185f
C775 B.n516 VSUBS 0.008185f
C776 B.n517 VSUBS 0.008185f
C777 B.n518 VSUBS 0.008185f
C778 B.n519 VSUBS 0.008185f
C779 B.n520 VSUBS 0.008185f
C780 B.n521 VSUBS 0.008185f
C781 B.n522 VSUBS 0.008185f
C782 B.n523 VSUBS 0.008185f
C783 B.n524 VSUBS 0.008185f
C784 B.n525 VSUBS 0.008185f
C785 B.n526 VSUBS 0.008185f
C786 B.n527 VSUBS 0.008185f
C787 B.n528 VSUBS 0.008185f
C788 B.n529 VSUBS 0.008185f
C789 B.n530 VSUBS 0.008185f
C790 B.n531 VSUBS 0.008185f
C791 B.n532 VSUBS 0.008185f
C792 B.n533 VSUBS 0.008185f
C793 B.n534 VSUBS 0.008185f
C794 B.n535 VSUBS 0.008185f
C795 B.n536 VSUBS 0.008185f
C796 B.n537 VSUBS 0.008185f
C797 B.n538 VSUBS 0.008185f
C798 B.n539 VSUBS 0.008185f
C799 B.n540 VSUBS 0.008185f
C800 B.n541 VSUBS 0.008185f
C801 B.n542 VSUBS 0.008185f
C802 B.n543 VSUBS 0.008185f
C803 B.n544 VSUBS 0.008185f
C804 B.n545 VSUBS 0.008185f
C805 B.n546 VSUBS 0.008185f
C806 B.n547 VSUBS 0.008185f
C807 B.n548 VSUBS 0.008185f
C808 B.n549 VSUBS 0.008185f
C809 B.n550 VSUBS 0.008185f
C810 B.n551 VSUBS 0.008185f
C811 B.n552 VSUBS 0.008185f
C812 B.n553 VSUBS 0.008185f
C813 B.n554 VSUBS 0.008185f
C814 B.n555 VSUBS 0.008185f
C815 B.n556 VSUBS 0.008185f
C816 B.n557 VSUBS 0.008185f
C817 B.n558 VSUBS 0.008185f
C818 B.n559 VSUBS 0.008185f
C819 B.n560 VSUBS 0.008185f
C820 B.n561 VSUBS 0.008185f
C821 B.n562 VSUBS 0.008185f
C822 B.n563 VSUBS 0.008185f
C823 B.n564 VSUBS 0.008185f
C824 B.n565 VSUBS 0.008185f
C825 B.n566 VSUBS 0.008185f
C826 B.n567 VSUBS 0.008185f
C827 B.n568 VSUBS 0.008185f
C828 B.n569 VSUBS 0.008185f
C829 B.n570 VSUBS 0.008185f
C830 B.n571 VSUBS 0.008185f
C831 B.n572 VSUBS 0.008185f
C832 B.n573 VSUBS 0.008185f
C833 B.n574 VSUBS 0.008185f
C834 B.n575 VSUBS 0.008185f
C835 B.n576 VSUBS 0.007704f
C836 B.n577 VSUBS 0.008185f
C837 B.n578 VSUBS 0.008185f
C838 B.n579 VSUBS 0.008185f
C839 B.n580 VSUBS 0.008185f
C840 B.n581 VSUBS 0.008185f
C841 B.n582 VSUBS 0.008185f
C842 B.n583 VSUBS 0.008185f
C843 B.n584 VSUBS 0.008185f
C844 B.n585 VSUBS 0.008185f
C845 B.n586 VSUBS 0.008185f
C846 B.n587 VSUBS 0.008185f
C847 B.n588 VSUBS 0.008185f
C848 B.n589 VSUBS 0.008185f
C849 B.n590 VSUBS 0.008185f
C850 B.n591 VSUBS 0.008185f
C851 B.n592 VSUBS 0.004574f
C852 B.n593 VSUBS 0.018964f
C853 B.n594 VSUBS 0.007704f
C854 B.n595 VSUBS 0.008185f
C855 B.n596 VSUBS 0.008185f
C856 B.n597 VSUBS 0.008185f
C857 B.n598 VSUBS 0.008185f
C858 B.n599 VSUBS 0.008185f
C859 B.n600 VSUBS 0.008185f
C860 B.n601 VSUBS 0.008185f
C861 B.n602 VSUBS 0.008185f
C862 B.n603 VSUBS 0.008185f
C863 B.n604 VSUBS 0.008185f
C864 B.n605 VSUBS 0.008185f
C865 B.n606 VSUBS 0.008185f
C866 B.n607 VSUBS 0.008185f
C867 B.n608 VSUBS 0.008185f
C868 B.n609 VSUBS 0.008185f
C869 B.n610 VSUBS 0.008185f
C870 B.n611 VSUBS 0.008185f
C871 B.n612 VSUBS 0.008185f
C872 B.n613 VSUBS 0.008185f
C873 B.n614 VSUBS 0.008185f
C874 B.n615 VSUBS 0.008185f
C875 B.n616 VSUBS 0.008185f
C876 B.n617 VSUBS 0.008185f
C877 B.n618 VSUBS 0.008185f
C878 B.n619 VSUBS 0.008185f
C879 B.n620 VSUBS 0.008185f
C880 B.n621 VSUBS 0.008185f
C881 B.n622 VSUBS 0.008185f
C882 B.n623 VSUBS 0.008185f
C883 B.n624 VSUBS 0.008185f
C884 B.n625 VSUBS 0.008185f
C885 B.n626 VSUBS 0.008185f
C886 B.n627 VSUBS 0.008185f
C887 B.n628 VSUBS 0.008185f
C888 B.n629 VSUBS 0.008185f
C889 B.n630 VSUBS 0.008185f
C890 B.n631 VSUBS 0.008185f
C891 B.n632 VSUBS 0.008185f
C892 B.n633 VSUBS 0.008185f
C893 B.n634 VSUBS 0.008185f
C894 B.n635 VSUBS 0.008185f
C895 B.n636 VSUBS 0.008185f
C896 B.n637 VSUBS 0.008185f
C897 B.n638 VSUBS 0.008185f
C898 B.n639 VSUBS 0.008185f
C899 B.n640 VSUBS 0.008185f
C900 B.n641 VSUBS 0.008185f
C901 B.n642 VSUBS 0.008185f
C902 B.n643 VSUBS 0.008185f
C903 B.n644 VSUBS 0.008185f
C904 B.n645 VSUBS 0.008185f
C905 B.n646 VSUBS 0.008185f
C906 B.n647 VSUBS 0.008185f
C907 B.n648 VSUBS 0.008185f
C908 B.n649 VSUBS 0.008185f
C909 B.n650 VSUBS 0.008185f
C910 B.n651 VSUBS 0.008185f
C911 B.n652 VSUBS 0.008185f
C912 B.n653 VSUBS 0.008185f
C913 B.n654 VSUBS 0.008185f
C914 B.n655 VSUBS 0.008185f
C915 B.n656 VSUBS 0.008185f
C916 B.n657 VSUBS 0.008185f
C917 B.n658 VSUBS 0.008185f
C918 B.n659 VSUBS 0.008185f
C919 B.n660 VSUBS 0.008185f
C920 B.n661 VSUBS 0.008185f
C921 B.n662 VSUBS 0.008185f
C922 B.n663 VSUBS 0.008185f
C923 B.n664 VSUBS 0.008185f
C924 B.n665 VSUBS 0.008185f
C925 B.n666 VSUBS 0.008185f
C926 B.n667 VSUBS 0.008185f
C927 B.n668 VSUBS 0.008185f
C928 B.n669 VSUBS 0.008185f
C929 B.n670 VSUBS 0.020408f
C930 B.n671 VSUBS 0.020408f
C931 B.n672 VSUBS 0.019314f
C932 B.n673 VSUBS 0.008185f
C933 B.n674 VSUBS 0.008185f
C934 B.n675 VSUBS 0.008185f
C935 B.n676 VSUBS 0.008185f
C936 B.n677 VSUBS 0.008185f
C937 B.n678 VSUBS 0.008185f
C938 B.n679 VSUBS 0.008185f
C939 B.n680 VSUBS 0.008185f
C940 B.n681 VSUBS 0.008185f
C941 B.n682 VSUBS 0.008185f
C942 B.n683 VSUBS 0.008185f
C943 B.n684 VSUBS 0.008185f
C944 B.n685 VSUBS 0.008185f
C945 B.n686 VSUBS 0.008185f
C946 B.n687 VSUBS 0.008185f
C947 B.n688 VSUBS 0.008185f
C948 B.n689 VSUBS 0.008185f
C949 B.n690 VSUBS 0.008185f
C950 B.n691 VSUBS 0.008185f
C951 B.n692 VSUBS 0.008185f
C952 B.n693 VSUBS 0.008185f
C953 B.n694 VSUBS 0.008185f
C954 B.n695 VSUBS 0.008185f
C955 B.n696 VSUBS 0.008185f
C956 B.n697 VSUBS 0.008185f
C957 B.n698 VSUBS 0.008185f
C958 B.n699 VSUBS 0.008185f
C959 B.n700 VSUBS 0.008185f
C960 B.n701 VSUBS 0.008185f
C961 B.n702 VSUBS 0.008185f
C962 B.n703 VSUBS 0.008185f
C963 B.n704 VSUBS 0.008185f
C964 B.n705 VSUBS 0.008185f
C965 B.n706 VSUBS 0.008185f
C966 B.n707 VSUBS 0.008185f
C967 B.n708 VSUBS 0.008185f
C968 B.n709 VSUBS 0.008185f
C969 B.n710 VSUBS 0.008185f
C970 B.n711 VSUBS 0.008185f
C971 B.n712 VSUBS 0.008185f
C972 B.n713 VSUBS 0.008185f
C973 B.n714 VSUBS 0.008185f
C974 B.n715 VSUBS 0.008185f
C975 B.n716 VSUBS 0.008185f
C976 B.n717 VSUBS 0.008185f
C977 B.n718 VSUBS 0.008185f
C978 B.n719 VSUBS 0.018534f
C979 VDD2.n0 VSUBS 0.030869f
C980 VDD2.n1 VSUBS 0.027251f
C981 VDD2.n2 VSUBS 0.014644f
C982 VDD2.n3 VSUBS 0.034612f
C983 VDD2.n4 VSUBS 0.015505f
C984 VDD2.n5 VSUBS 0.027251f
C985 VDD2.n6 VSUBS 0.014644f
C986 VDD2.n7 VSUBS 0.034612f
C987 VDD2.n8 VSUBS 0.015505f
C988 VDD2.n9 VSUBS 0.027251f
C989 VDD2.n10 VSUBS 0.014644f
C990 VDD2.n11 VSUBS 0.034612f
C991 VDD2.n12 VSUBS 0.015505f
C992 VDD2.n13 VSUBS 0.027251f
C993 VDD2.n14 VSUBS 0.014644f
C994 VDD2.n15 VSUBS 0.034612f
C995 VDD2.n16 VSUBS 0.015074f
C996 VDD2.n17 VSUBS 0.027251f
C997 VDD2.n18 VSUBS 0.015505f
C998 VDD2.n19 VSUBS 0.034612f
C999 VDD2.n20 VSUBS 0.015505f
C1000 VDD2.n21 VSUBS 0.027251f
C1001 VDD2.n22 VSUBS 0.014644f
C1002 VDD2.n23 VSUBS 0.034612f
C1003 VDD2.n24 VSUBS 0.015505f
C1004 VDD2.n25 VSUBS 1.77001f
C1005 VDD2.n26 VSUBS 0.014644f
C1006 VDD2.t5 VSUBS 0.074915f
C1007 VDD2.n27 VSUBS 0.259101f
C1008 VDD2.n28 VSUBS 0.026037f
C1009 VDD2.n29 VSUBS 0.025959f
C1010 VDD2.n30 VSUBS 0.034612f
C1011 VDD2.n31 VSUBS 0.015505f
C1012 VDD2.n32 VSUBS 0.014644f
C1013 VDD2.n33 VSUBS 0.027251f
C1014 VDD2.n34 VSUBS 0.027251f
C1015 VDD2.n35 VSUBS 0.014644f
C1016 VDD2.n36 VSUBS 0.015505f
C1017 VDD2.n37 VSUBS 0.034612f
C1018 VDD2.n38 VSUBS 0.034612f
C1019 VDD2.n39 VSUBS 0.015505f
C1020 VDD2.n40 VSUBS 0.014644f
C1021 VDD2.n41 VSUBS 0.027251f
C1022 VDD2.n42 VSUBS 0.027251f
C1023 VDD2.n43 VSUBS 0.014644f
C1024 VDD2.n44 VSUBS 0.014644f
C1025 VDD2.n45 VSUBS 0.015505f
C1026 VDD2.n46 VSUBS 0.034612f
C1027 VDD2.n47 VSUBS 0.034612f
C1028 VDD2.n48 VSUBS 0.034612f
C1029 VDD2.n49 VSUBS 0.015074f
C1030 VDD2.n50 VSUBS 0.014644f
C1031 VDD2.n51 VSUBS 0.027251f
C1032 VDD2.n52 VSUBS 0.027251f
C1033 VDD2.n53 VSUBS 0.014644f
C1034 VDD2.n54 VSUBS 0.015505f
C1035 VDD2.n55 VSUBS 0.034612f
C1036 VDD2.n56 VSUBS 0.034612f
C1037 VDD2.n57 VSUBS 0.015505f
C1038 VDD2.n58 VSUBS 0.014644f
C1039 VDD2.n59 VSUBS 0.027251f
C1040 VDD2.n60 VSUBS 0.027251f
C1041 VDD2.n61 VSUBS 0.014644f
C1042 VDD2.n62 VSUBS 0.015505f
C1043 VDD2.n63 VSUBS 0.034612f
C1044 VDD2.n64 VSUBS 0.034612f
C1045 VDD2.n65 VSUBS 0.015505f
C1046 VDD2.n66 VSUBS 0.014644f
C1047 VDD2.n67 VSUBS 0.027251f
C1048 VDD2.n68 VSUBS 0.027251f
C1049 VDD2.n69 VSUBS 0.014644f
C1050 VDD2.n70 VSUBS 0.015505f
C1051 VDD2.n71 VSUBS 0.034612f
C1052 VDD2.n72 VSUBS 0.034612f
C1053 VDD2.n73 VSUBS 0.015505f
C1054 VDD2.n74 VSUBS 0.014644f
C1055 VDD2.n75 VSUBS 0.027251f
C1056 VDD2.n76 VSUBS 0.027251f
C1057 VDD2.n77 VSUBS 0.014644f
C1058 VDD2.n78 VSUBS 0.015505f
C1059 VDD2.n79 VSUBS 0.034612f
C1060 VDD2.n80 VSUBS 0.086946f
C1061 VDD2.n81 VSUBS 0.015505f
C1062 VDD2.n82 VSUBS 0.014644f
C1063 VDD2.n83 VSUBS 0.058895f
C1064 VDD2.n84 VSUBS 0.066557f
C1065 VDD2.t3 VSUBS 0.33616f
C1066 VDD2.t1 VSUBS 0.33616f
C1067 VDD2.n85 VSUBS 2.72472f
C1068 VDD2.n86 VSUBS 3.02312f
C1069 VDD2.n87 VSUBS 0.030869f
C1070 VDD2.n88 VSUBS 0.027251f
C1071 VDD2.n89 VSUBS 0.014644f
C1072 VDD2.n90 VSUBS 0.034612f
C1073 VDD2.n91 VSUBS 0.015505f
C1074 VDD2.n92 VSUBS 0.027251f
C1075 VDD2.n93 VSUBS 0.014644f
C1076 VDD2.n94 VSUBS 0.034612f
C1077 VDD2.n95 VSUBS 0.015505f
C1078 VDD2.n96 VSUBS 0.027251f
C1079 VDD2.n97 VSUBS 0.014644f
C1080 VDD2.n98 VSUBS 0.034612f
C1081 VDD2.n99 VSUBS 0.015505f
C1082 VDD2.n100 VSUBS 0.027251f
C1083 VDD2.n101 VSUBS 0.014644f
C1084 VDD2.n102 VSUBS 0.034612f
C1085 VDD2.n103 VSUBS 0.015074f
C1086 VDD2.n104 VSUBS 0.027251f
C1087 VDD2.n105 VSUBS 0.015074f
C1088 VDD2.n106 VSUBS 0.014644f
C1089 VDD2.n107 VSUBS 0.034612f
C1090 VDD2.n108 VSUBS 0.034612f
C1091 VDD2.n109 VSUBS 0.015505f
C1092 VDD2.n110 VSUBS 0.027251f
C1093 VDD2.n111 VSUBS 0.014644f
C1094 VDD2.n112 VSUBS 0.034612f
C1095 VDD2.n113 VSUBS 0.015505f
C1096 VDD2.n114 VSUBS 1.77001f
C1097 VDD2.n115 VSUBS 0.014644f
C1098 VDD2.t4 VSUBS 0.074915f
C1099 VDD2.n116 VSUBS 0.259101f
C1100 VDD2.n117 VSUBS 0.026037f
C1101 VDD2.n118 VSUBS 0.025959f
C1102 VDD2.n119 VSUBS 0.034612f
C1103 VDD2.n120 VSUBS 0.015505f
C1104 VDD2.n121 VSUBS 0.014644f
C1105 VDD2.n122 VSUBS 0.027251f
C1106 VDD2.n123 VSUBS 0.027251f
C1107 VDD2.n124 VSUBS 0.014644f
C1108 VDD2.n125 VSUBS 0.015505f
C1109 VDD2.n126 VSUBS 0.034612f
C1110 VDD2.n127 VSUBS 0.034612f
C1111 VDD2.n128 VSUBS 0.015505f
C1112 VDD2.n129 VSUBS 0.014644f
C1113 VDD2.n130 VSUBS 0.027251f
C1114 VDD2.n131 VSUBS 0.027251f
C1115 VDD2.n132 VSUBS 0.014644f
C1116 VDD2.n133 VSUBS 0.015505f
C1117 VDD2.n134 VSUBS 0.034612f
C1118 VDD2.n135 VSUBS 0.034612f
C1119 VDD2.n136 VSUBS 0.015505f
C1120 VDD2.n137 VSUBS 0.014644f
C1121 VDD2.n138 VSUBS 0.027251f
C1122 VDD2.n139 VSUBS 0.027251f
C1123 VDD2.n140 VSUBS 0.014644f
C1124 VDD2.n141 VSUBS 0.015505f
C1125 VDD2.n142 VSUBS 0.034612f
C1126 VDD2.n143 VSUBS 0.034612f
C1127 VDD2.n144 VSUBS 0.015505f
C1128 VDD2.n145 VSUBS 0.014644f
C1129 VDD2.n146 VSUBS 0.027251f
C1130 VDD2.n147 VSUBS 0.027251f
C1131 VDD2.n148 VSUBS 0.014644f
C1132 VDD2.n149 VSUBS 0.015505f
C1133 VDD2.n150 VSUBS 0.034612f
C1134 VDD2.n151 VSUBS 0.034612f
C1135 VDD2.n152 VSUBS 0.015505f
C1136 VDD2.n153 VSUBS 0.014644f
C1137 VDD2.n154 VSUBS 0.027251f
C1138 VDD2.n155 VSUBS 0.027251f
C1139 VDD2.n156 VSUBS 0.014644f
C1140 VDD2.n157 VSUBS 0.015505f
C1141 VDD2.n158 VSUBS 0.034612f
C1142 VDD2.n159 VSUBS 0.034612f
C1143 VDD2.n160 VSUBS 0.015505f
C1144 VDD2.n161 VSUBS 0.014644f
C1145 VDD2.n162 VSUBS 0.027251f
C1146 VDD2.n163 VSUBS 0.027251f
C1147 VDD2.n164 VSUBS 0.014644f
C1148 VDD2.n165 VSUBS 0.015505f
C1149 VDD2.n166 VSUBS 0.034612f
C1150 VDD2.n167 VSUBS 0.086946f
C1151 VDD2.n168 VSUBS 0.015505f
C1152 VDD2.n169 VSUBS 0.014644f
C1153 VDD2.n170 VSUBS 0.058895f
C1154 VDD2.n171 VSUBS 0.062586f
C1155 VDD2.n172 VSUBS 2.8047f
C1156 VDD2.t0 VSUBS 0.33616f
C1157 VDD2.t2 VSUBS 0.33616f
C1158 VDD2.n173 VSUBS 2.72469f
C1159 VTAIL.t6 VSUBS 0.339854f
C1160 VTAIL.t9 VSUBS 0.339854f
C1161 VTAIL.n0 VSUBS 2.57399f
C1162 VTAIL.n1 VSUBS 0.851802f
C1163 VTAIL.n2 VSUBS 0.031208f
C1164 VTAIL.n3 VSUBS 0.027551f
C1165 VTAIL.n4 VSUBS 0.014805f
C1166 VTAIL.n5 VSUBS 0.034993f
C1167 VTAIL.n6 VSUBS 0.015676f
C1168 VTAIL.n7 VSUBS 0.027551f
C1169 VTAIL.n8 VSUBS 0.014805f
C1170 VTAIL.n9 VSUBS 0.034993f
C1171 VTAIL.n10 VSUBS 0.015676f
C1172 VTAIL.n11 VSUBS 0.027551f
C1173 VTAIL.n12 VSUBS 0.014805f
C1174 VTAIL.n13 VSUBS 0.034993f
C1175 VTAIL.n14 VSUBS 0.015676f
C1176 VTAIL.n15 VSUBS 0.027551f
C1177 VTAIL.n16 VSUBS 0.014805f
C1178 VTAIL.n17 VSUBS 0.034993f
C1179 VTAIL.n18 VSUBS 0.01524f
C1180 VTAIL.n19 VSUBS 0.027551f
C1181 VTAIL.n20 VSUBS 0.015676f
C1182 VTAIL.n21 VSUBS 0.034993f
C1183 VTAIL.n22 VSUBS 0.015676f
C1184 VTAIL.n23 VSUBS 0.027551f
C1185 VTAIL.n24 VSUBS 0.014805f
C1186 VTAIL.n25 VSUBS 0.034993f
C1187 VTAIL.n26 VSUBS 0.015676f
C1188 VTAIL.n27 VSUBS 1.78946f
C1189 VTAIL.n28 VSUBS 0.014805f
C1190 VTAIL.t5 VSUBS 0.075739f
C1191 VTAIL.n29 VSUBS 0.261948f
C1192 VTAIL.n30 VSUBS 0.026323f
C1193 VTAIL.n31 VSUBS 0.026245f
C1194 VTAIL.n32 VSUBS 0.034993f
C1195 VTAIL.n33 VSUBS 0.015676f
C1196 VTAIL.n34 VSUBS 0.014805f
C1197 VTAIL.n35 VSUBS 0.027551f
C1198 VTAIL.n36 VSUBS 0.027551f
C1199 VTAIL.n37 VSUBS 0.014805f
C1200 VTAIL.n38 VSUBS 0.015676f
C1201 VTAIL.n39 VSUBS 0.034993f
C1202 VTAIL.n40 VSUBS 0.034993f
C1203 VTAIL.n41 VSUBS 0.015676f
C1204 VTAIL.n42 VSUBS 0.014805f
C1205 VTAIL.n43 VSUBS 0.027551f
C1206 VTAIL.n44 VSUBS 0.027551f
C1207 VTAIL.n45 VSUBS 0.014805f
C1208 VTAIL.n46 VSUBS 0.014805f
C1209 VTAIL.n47 VSUBS 0.015676f
C1210 VTAIL.n48 VSUBS 0.034993f
C1211 VTAIL.n49 VSUBS 0.034993f
C1212 VTAIL.n50 VSUBS 0.034993f
C1213 VTAIL.n51 VSUBS 0.01524f
C1214 VTAIL.n52 VSUBS 0.014805f
C1215 VTAIL.n53 VSUBS 0.027551f
C1216 VTAIL.n54 VSUBS 0.027551f
C1217 VTAIL.n55 VSUBS 0.014805f
C1218 VTAIL.n56 VSUBS 0.015676f
C1219 VTAIL.n57 VSUBS 0.034993f
C1220 VTAIL.n58 VSUBS 0.034993f
C1221 VTAIL.n59 VSUBS 0.015676f
C1222 VTAIL.n60 VSUBS 0.014805f
C1223 VTAIL.n61 VSUBS 0.027551f
C1224 VTAIL.n62 VSUBS 0.027551f
C1225 VTAIL.n63 VSUBS 0.014805f
C1226 VTAIL.n64 VSUBS 0.015676f
C1227 VTAIL.n65 VSUBS 0.034993f
C1228 VTAIL.n66 VSUBS 0.034993f
C1229 VTAIL.n67 VSUBS 0.015676f
C1230 VTAIL.n68 VSUBS 0.014805f
C1231 VTAIL.n69 VSUBS 0.027551f
C1232 VTAIL.n70 VSUBS 0.027551f
C1233 VTAIL.n71 VSUBS 0.014805f
C1234 VTAIL.n72 VSUBS 0.015676f
C1235 VTAIL.n73 VSUBS 0.034993f
C1236 VTAIL.n74 VSUBS 0.034993f
C1237 VTAIL.n75 VSUBS 0.015676f
C1238 VTAIL.n76 VSUBS 0.014805f
C1239 VTAIL.n77 VSUBS 0.027551f
C1240 VTAIL.n78 VSUBS 0.027551f
C1241 VTAIL.n79 VSUBS 0.014805f
C1242 VTAIL.n80 VSUBS 0.015676f
C1243 VTAIL.n81 VSUBS 0.034993f
C1244 VTAIL.n82 VSUBS 0.087902f
C1245 VTAIL.n83 VSUBS 0.015676f
C1246 VTAIL.n84 VSUBS 0.014805f
C1247 VTAIL.n85 VSUBS 0.059542f
C1248 VTAIL.n86 VSUBS 0.044215f
C1249 VTAIL.n87 VSUBS 0.287906f
C1250 VTAIL.t1 VSUBS 0.339854f
C1251 VTAIL.t3 VSUBS 0.339854f
C1252 VTAIL.n88 VSUBS 2.57399f
C1253 VTAIL.n89 VSUBS 2.71131f
C1254 VTAIL.t11 VSUBS 0.339854f
C1255 VTAIL.t8 VSUBS 0.339854f
C1256 VTAIL.n90 VSUBS 2.574f
C1257 VTAIL.n91 VSUBS 2.7113f
C1258 VTAIL.n92 VSUBS 0.031208f
C1259 VTAIL.n93 VSUBS 0.027551f
C1260 VTAIL.n94 VSUBS 0.014805f
C1261 VTAIL.n95 VSUBS 0.034993f
C1262 VTAIL.n96 VSUBS 0.015676f
C1263 VTAIL.n97 VSUBS 0.027551f
C1264 VTAIL.n98 VSUBS 0.014805f
C1265 VTAIL.n99 VSUBS 0.034993f
C1266 VTAIL.n100 VSUBS 0.015676f
C1267 VTAIL.n101 VSUBS 0.027551f
C1268 VTAIL.n102 VSUBS 0.014805f
C1269 VTAIL.n103 VSUBS 0.034993f
C1270 VTAIL.n104 VSUBS 0.015676f
C1271 VTAIL.n105 VSUBS 0.027551f
C1272 VTAIL.n106 VSUBS 0.014805f
C1273 VTAIL.n107 VSUBS 0.034993f
C1274 VTAIL.n108 VSUBS 0.01524f
C1275 VTAIL.n109 VSUBS 0.027551f
C1276 VTAIL.n110 VSUBS 0.01524f
C1277 VTAIL.n111 VSUBS 0.014805f
C1278 VTAIL.n112 VSUBS 0.034993f
C1279 VTAIL.n113 VSUBS 0.034993f
C1280 VTAIL.n114 VSUBS 0.015676f
C1281 VTAIL.n115 VSUBS 0.027551f
C1282 VTAIL.n116 VSUBS 0.014805f
C1283 VTAIL.n117 VSUBS 0.034993f
C1284 VTAIL.n118 VSUBS 0.015676f
C1285 VTAIL.n119 VSUBS 1.78946f
C1286 VTAIL.n120 VSUBS 0.014805f
C1287 VTAIL.t7 VSUBS 0.075739f
C1288 VTAIL.n121 VSUBS 0.261948f
C1289 VTAIL.n122 VSUBS 0.026323f
C1290 VTAIL.n123 VSUBS 0.026245f
C1291 VTAIL.n124 VSUBS 0.034993f
C1292 VTAIL.n125 VSUBS 0.015676f
C1293 VTAIL.n126 VSUBS 0.014805f
C1294 VTAIL.n127 VSUBS 0.027551f
C1295 VTAIL.n128 VSUBS 0.027551f
C1296 VTAIL.n129 VSUBS 0.014805f
C1297 VTAIL.n130 VSUBS 0.015676f
C1298 VTAIL.n131 VSUBS 0.034993f
C1299 VTAIL.n132 VSUBS 0.034993f
C1300 VTAIL.n133 VSUBS 0.015676f
C1301 VTAIL.n134 VSUBS 0.014805f
C1302 VTAIL.n135 VSUBS 0.027551f
C1303 VTAIL.n136 VSUBS 0.027551f
C1304 VTAIL.n137 VSUBS 0.014805f
C1305 VTAIL.n138 VSUBS 0.015676f
C1306 VTAIL.n139 VSUBS 0.034993f
C1307 VTAIL.n140 VSUBS 0.034993f
C1308 VTAIL.n141 VSUBS 0.015676f
C1309 VTAIL.n142 VSUBS 0.014805f
C1310 VTAIL.n143 VSUBS 0.027551f
C1311 VTAIL.n144 VSUBS 0.027551f
C1312 VTAIL.n145 VSUBS 0.014805f
C1313 VTAIL.n146 VSUBS 0.015676f
C1314 VTAIL.n147 VSUBS 0.034993f
C1315 VTAIL.n148 VSUBS 0.034993f
C1316 VTAIL.n149 VSUBS 0.015676f
C1317 VTAIL.n150 VSUBS 0.014805f
C1318 VTAIL.n151 VSUBS 0.027551f
C1319 VTAIL.n152 VSUBS 0.027551f
C1320 VTAIL.n153 VSUBS 0.014805f
C1321 VTAIL.n154 VSUBS 0.015676f
C1322 VTAIL.n155 VSUBS 0.034993f
C1323 VTAIL.n156 VSUBS 0.034993f
C1324 VTAIL.n157 VSUBS 0.015676f
C1325 VTAIL.n158 VSUBS 0.014805f
C1326 VTAIL.n159 VSUBS 0.027551f
C1327 VTAIL.n160 VSUBS 0.027551f
C1328 VTAIL.n161 VSUBS 0.014805f
C1329 VTAIL.n162 VSUBS 0.015676f
C1330 VTAIL.n163 VSUBS 0.034993f
C1331 VTAIL.n164 VSUBS 0.034993f
C1332 VTAIL.n165 VSUBS 0.015676f
C1333 VTAIL.n166 VSUBS 0.014805f
C1334 VTAIL.n167 VSUBS 0.027551f
C1335 VTAIL.n168 VSUBS 0.027551f
C1336 VTAIL.n169 VSUBS 0.014805f
C1337 VTAIL.n170 VSUBS 0.015676f
C1338 VTAIL.n171 VSUBS 0.034993f
C1339 VTAIL.n172 VSUBS 0.087902f
C1340 VTAIL.n173 VSUBS 0.015676f
C1341 VTAIL.n174 VSUBS 0.014805f
C1342 VTAIL.n175 VSUBS 0.059542f
C1343 VTAIL.n176 VSUBS 0.044215f
C1344 VTAIL.n177 VSUBS 0.287906f
C1345 VTAIL.t4 VSUBS 0.339854f
C1346 VTAIL.t0 VSUBS 0.339854f
C1347 VTAIL.n178 VSUBS 2.574f
C1348 VTAIL.n179 VSUBS 0.959123f
C1349 VTAIL.n180 VSUBS 0.031208f
C1350 VTAIL.n181 VSUBS 0.027551f
C1351 VTAIL.n182 VSUBS 0.014805f
C1352 VTAIL.n183 VSUBS 0.034993f
C1353 VTAIL.n184 VSUBS 0.015676f
C1354 VTAIL.n185 VSUBS 0.027551f
C1355 VTAIL.n186 VSUBS 0.014805f
C1356 VTAIL.n187 VSUBS 0.034993f
C1357 VTAIL.n188 VSUBS 0.015676f
C1358 VTAIL.n189 VSUBS 0.027551f
C1359 VTAIL.n190 VSUBS 0.014805f
C1360 VTAIL.n191 VSUBS 0.034993f
C1361 VTAIL.n192 VSUBS 0.015676f
C1362 VTAIL.n193 VSUBS 0.027551f
C1363 VTAIL.n194 VSUBS 0.014805f
C1364 VTAIL.n195 VSUBS 0.034993f
C1365 VTAIL.n196 VSUBS 0.01524f
C1366 VTAIL.n197 VSUBS 0.027551f
C1367 VTAIL.n198 VSUBS 0.01524f
C1368 VTAIL.n199 VSUBS 0.014805f
C1369 VTAIL.n200 VSUBS 0.034993f
C1370 VTAIL.n201 VSUBS 0.034993f
C1371 VTAIL.n202 VSUBS 0.015676f
C1372 VTAIL.n203 VSUBS 0.027551f
C1373 VTAIL.n204 VSUBS 0.014805f
C1374 VTAIL.n205 VSUBS 0.034993f
C1375 VTAIL.n206 VSUBS 0.015676f
C1376 VTAIL.n207 VSUBS 1.78946f
C1377 VTAIL.n208 VSUBS 0.014805f
C1378 VTAIL.t2 VSUBS 0.075739f
C1379 VTAIL.n209 VSUBS 0.261948f
C1380 VTAIL.n210 VSUBS 0.026323f
C1381 VTAIL.n211 VSUBS 0.026245f
C1382 VTAIL.n212 VSUBS 0.034993f
C1383 VTAIL.n213 VSUBS 0.015676f
C1384 VTAIL.n214 VSUBS 0.014805f
C1385 VTAIL.n215 VSUBS 0.027551f
C1386 VTAIL.n216 VSUBS 0.027551f
C1387 VTAIL.n217 VSUBS 0.014805f
C1388 VTAIL.n218 VSUBS 0.015676f
C1389 VTAIL.n219 VSUBS 0.034993f
C1390 VTAIL.n220 VSUBS 0.034993f
C1391 VTAIL.n221 VSUBS 0.015676f
C1392 VTAIL.n222 VSUBS 0.014805f
C1393 VTAIL.n223 VSUBS 0.027551f
C1394 VTAIL.n224 VSUBS 0.027551f
C1395 VTAIL.n225 VSUBS 0.014805f
C1396 VTAIL.n226 VSUBS 0.015676f
C1397 VTAIL.n227 VSUBS 0.034993f
C1398 VTAIL.n228 VSUBS 0.034993f
C1399 VTAIL.n229 VSUBS 0.015676f
C1400 VTAIL.n230 VSUBS 0.014805f
C1401 VTAIL.n231 VSUBS 0.027551f
C1402 VTAIL.n232 VSUBS 0.027551f
C1403 VTAIL.n233 VSUBS 0.014805f
C1404 VTAIL.n234 VSUBS 0.015676f
C1405 VTAIL.n235 VSUBS 0.034993f
C1406 VTAIL.n236 VSUBS 0.034993f
C1407 VTAIL.n237 VSUBS 0.015676f
C1408 VTAIL.n238 VSUBS 0.014805f
C1409 VTAIL.n239 VSUBS 0.027551f
C1410 VTAIL.n240 VSUBS 0.027551f
C1411 VTAIL.n241 VSUBS 0.014805f
C1412 VTAIL.n242 VSUBS 0.015676f
C1413 VTAIL.n243 VSUBS 0.034993f
C1414 VTAIL.n244 VSUBS 0.034993f
C1415 VTAIL.n245 VSUBS 0.015676f
C1416 VTAIL.n246 VSUBS 0.014805f
C1417 VTAIL.n247 VSUBS 0.027551f
C1418 VTAIL.n248 VSUBS 0.027551f
C1419 VTAIL.n249 VSUBS 0.014805f
C1420 VTAIL.n250 VSUBS 0.015676f
C1421 VTAIL.n251 VSUBS 0.034993f
C1422 VTAIL.n252 VSUBS 0.034993f
C1423 VTAIL.n253 VSUBS 0.015676f
C1424 VTAIL.n254 VSUBS 0.014805f
C1425 VTAIL.n255 VSUBS 0.027551f
C1426 VTAIL.n256 VSUBS 0.027551f
C1427 VTAIL.n257 VSUBS 0.014805f
C1428 VTAIL.n258 VSUBS 0.015676f
C1429 VTAIL.n259 VSUBS 0.034993f
C1430 VTAIL.n260 VSUBS 0.087902f
C1431 VTAIL.n261 VSUBS 0.015676f
C1432 VTAIL.n262 VSUBS 0.014805f
C1433 VTAIL.n263 VSUBS 0.059542f
C1434 VTAIL.n264 VSUBS 0.044215f
C1435 VTAIL.n265 VSUBS 1.89008f
C1436 VTAIL.n266 VSUBS 0.031208f
C1437 VTAIL.n267 VSUBS 0.027551f
C1438 VTAIL.n268 VSUBS 0.014805f
C1439 VTAIL.n269 VSUBS 0.034993f
C1440 VTAIL.n270 VSUBS 0.015676f
C1441 VTAIL.n271 VSUBS 0.027551f
C1442 VTAIL.n272 VSUBS 0.014805f
C1443 VTAIL.n273 VSUBS 0.034993f
C1444 VTAIL.n274 VSUBS 0.015676f
C1445 VTAIL.n275 VSUBS 0.027551f
C1446 VTAIL.n276 VSUBS 0.014805f
C1447 VTAIL.n277 VSUBS 0.034993f
C1448 VTAIL.n278 VSUBS 0.015676f
C1449 VTAIL.n279 VSUBS 0.027551f
C1450 VTAIL.n280 VSUBS 0.014805f
C1451 VTAIL.n281 VSUBS 0.034993f
C1452 VTAIL.n282 VSUBS 0.01524f
C1453 VTAIL.n283 VSUBS 0.027551f
C1454 VTAIL.n284 VSUBS 0.015676f
C1455 VTAIL.n285 VSUBS 0.034993f
C1456 VTAIL.n286 VSUBS 0.015676f
C1457 VTAIL.n287 VSUBS 0.027551f
C1458 VTAIL.n288 VSUBS 0.014805f
C1459 VTAIL.n289 VSUBS 0.034993f
C1460 VTAIL.n290 VSUBS 0.015676f
C1461 VTAIL.n291 VSUBS 1.78946f
C1462 VTAIL.n292 VSUBS 0.014805f
C1463 VTAIL.t10 VSUBS 0.075739f
C1464 VTAIL.n293 VSUBS 0.261948f
C1465 VTAIL.n294 VSUBS 0.026323f
C1466 VTAIL.n295 VSUBS 0.026245f
C1467 VTAIL.n296 VSUBS 0.034993f
C1468 VTAIL.n297 VSUBS 0.015676f
C1469 VTAIL.n298 VSUBS 0.014805f
C1470 VTAIL.n299 VSUBS 0.027551f
C1471 VTAIL.n300 VSUBS 0.027551f
C1472 VTAIL.n301 VSUBS 0.014805f
C1473 VTAIL.n302 VSUBS 0.015676f
C1474 VTAIL.n303 VSUBS 0.034993f
C1475 VTAIL.n304 VSUBS 0.034993f
C1476 VTAIL.n305 VSUBS 0.015676f
C1477 VTAIL.n306 VSUBS 0.014805f
C1478 VTAIL.n307 VSUBS 0.027551f
C1479 VTAIL.n308 VSUBS 0.027551f
C1480 VTAIL.n309 VSUBS 0.014805f
C1481 VTAIL.n310 VSUBS 0.014805f
C1482 VTAIL.n311 VSUBS 0.015676f
C1483 VTAIL.n312 VSUBS 0.034993f
C1484 VTAIL.n313 VSUBS 0.034993f
C1485 VTAIL.n314 VSUBS 0.034993f
C1486 VTAIL.n315 VSUBS 0.01524f
C1487 VTAIL.n316 VSUBS 0.014805f
C1488 VTAIL.n317 VSUBS 0.027551f
C1489 VTAIL.n318 VSUBS 0.027551f
C1490 VTAIL.n319 VSUBS 0.014805f
C1491 VTAIL.n320 VSUBS 0.015676f
C1492 VTAIL.n321 VSUBS 0.034993f
C1493 VTAIL.n322 VSUBS 0.034993f
C1494 VTAIL.n323 VSUBS 0.015676f
C1495 VTAIL.n324 VSUBS 0.014805f
C1496 VTAIL.n325 VSUBS 0.027551f
C1497 VTAIL.n326 VSUBS 0.027551f
C1498 VTAIL.n327 VSUBS 0.014805f
C1499 VTAIL.n328 VSUBS 0.015676f
C1500 VTAIL.n329 VSUBS 0.034993f
C1501 VTAIL.n330 VSUBS 0.034993f
C1502 VTAIL.n331 VSUBS 0.015676f
C1503 VTAIL.n332 VSUBS 0.014805f
C1504 VTAIL.n333 VSUBS 0.027551f
C1505 VTAIL.n334 VSUBS 0.027551f
C1506 VTAIL.n335 VSUBS 0.014805f
C1507 VTAIL.n336 VSUBS 0.015676f
C1508 VTAIL.n337 VSUBS 0.034993f
C1509 VTAIL.n338 VSUBS 0.034993f
C1510 VTAIL.n339 VSUBS 0.015676f
C1511 VTAIL.n340 VSUBS 0.014805f
C1512 VTAIL.n341 VSUBS 0.027551f
C1513 VTAIL.n342 VSUBS 0.027551f
C1514 VTAIL.n343 VSUBS 0.014805f
C1515 VTAIL.n344 VSUBS 0.015676f
C1516 VTAIL.n345 VSUBS 0.034993f
C1517 VTAIL.n346 VSUBS 0.087902f
C1518 VTAIL.n347 VSUBS 0.015676f
C1519 VTAIL.n348 VSUBS 0.014805f
C1520 VTAIL.n349 VSUBS 0.059542f
C1521 VTAIL.n350 VSUBS 0.044215f
C1522 VTAIL.n351 VSUBS 1.84741f
C1523 VN.n0 VSUBS 0.036753f
C1524 VN.t4 VSUBS 2.56477f
C1525 VN.n1 VSUBS 0.051604f
C1526 VN.t0 VSUBS 2.70053f
C1527 VN.n2 VSUBS 0.995093f
C1528 VN.t2 VSUBS 2.56477f
C1529 VN.n3 VSUBS 0.979874f
C1530 VN.n4 VSUBS 0.051589f
C1531 VN.n5 VSUBS 0.236314f
C1532 VN.n6 VSUBS 0.036753f
C1533 VN.n7 VSUBS 0.036753f
C1534 VN.n8 VSUBS 0.055701f
C1535 VN.n9 VSUBS 0.048884f
C1536 VN.n10 VSUBS 0.99149f
C1537 VN.n11 VSUBS 0.035881f
C1538 VN.n12 VSUBS 0.036753f
C1539 VN.t1 VSUBS 2.56477f
C1540 VN.n13 VSUBS 0.051604f
C1541 VN.t3 VSUBS 2.70053f
C1542 VN.n14 VSUBS 0.995093f
C1543 VN.t5 VSUBS 2.56477f
C1544 VN.n15 VSUBS 0.979874f
C1545 VN.n16 VSUBS 0.051589f
C1546 VN.n17 VSUBS 0.236314f
C1547 VN.n18 VSUBS 0.036753f
C1548 VN.n19 VSUBS 0.036753f
C1549 VN.n20 VSUBS 0.055701f
C1550 VN.n21 VSUBS 0.048884f
C1551 VN.n22 VSUBS 0.99149f
C1552 VN.n23 VSUBS 1.88337f
.ends

