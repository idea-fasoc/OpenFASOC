* NGSPICE file created from diff_pair_sample_0563.ext - technology: sky130A

.subckt diff_pair_sample_0563 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=3.0195 ps=18.63 w=18.3 l=0.73
X1 VDD1.t8 VP.t1 VTAIL.t13 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=7.137 ps=37.38 w=18.3 l=0.73
X2 B.t11 B.t9 B.t10 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=0 ps=0 w=18.3 l=0.73
X3 VDD1.t7 VP.t2 VTAIL.t17 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X4 B.t8 B.t6 B.t7 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=0 ps=0 w=18.3 l=0.73
X5 VDD2.t9 VN.t0 VTAIL.t4 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=7.137 ps=37.38 w=18.3 l=0.73
X6 VTAIL.t1 VN.t1 VDD2.t8 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X7 VDD2.t7 VN.t2 VTAIL.t18 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=7.137 ps=37.38 w=18.3 l=0.73
X8 VDD2.t6 VN.t3 VTAIL.t3 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=3.0195 ps=18.63 w=18.3 l=0.73
X9 VDD2.t5 VN.t4 VTAIL.t0 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=3.0195 ps=18.63 w=18.3 l=0.73
X10 VDD2.t4 VN.t5 VTAIL.t19 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X11 VTAIL.t2 VN.t6 VDD2.t3 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X12 VDD2.t2 VN.t7 VTAIL.t6 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X13 VTAIL.t15 VP.t3 VDD1.t6 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X14 VDD1.t5 VP.t4 VTAIL.t16 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=3.0195 ps=18.63 w=18.3 l=0.73
X15 B.t5 B.t3 B.t4 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=0 ps=0 w=18.3 l=0.73
X16 VTAIL.t12 VP.t5 VDD1.t4 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X17 B.t2 B.t0 B.t1 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=7.137 pd=37.38 as=0 ps=0 w=18.3 l=0.73
X18 VTAIL.t10 VP.t6 VDD1.t3 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X19 VTAIL.t5 VN.t8 VDD2.t1 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X20 VTAIL.t7 VN.t9 VDD2.t0 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X21 VTAIL.t14 VP.t7 VDD1.t2 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X22 VDD1.t1 VP.t8 VTAIL.t8 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=3.0195 ps=18.63 w=18.3 l=0.73
X23 VDD1.t0 VP.t9 VTAIL.t9 w_n2242_n4628# sky130_fd_pr__pfet_01v8 ad=3.0195 pd=18.63 as=7.137 ps=37.38 w=18.3 l=0.73
R0 VP.n7 VP.t0 682.338
R1 VP.n18 VP.t4 657.963
R2 VP.n22 VP.t6 657.963
R3 VP.n24 VP.t8 657.963
R4 VP.n28 VP.t7 657.963
R5 VP.n30 VP.t9 657.963
R6 VP.n16 VP.t1 657.963
R7 VP.n14 VP.t5 657.963
R8 VP.n6 VP.t2 657.963
R9 VP.n8 VP.t3 657.963
R10 VP.n31 VP.n30 161.3
R11 VP.n10 VP.n9 161.3
R12 VP.n11 VP.n6 161.3
R13 VP.n13 VP.n12 161.3
R14 VP.n14 VP.n5 161.3
R15 VP.n15 VP.n4 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n29 VP.n0 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.n1 161.3
R20 VP.n25 VP.n24 161.3
R21 VP.n23 VP.n2 161.3
R22 VP.n22 VP.n21 161.3
R23 VP.n20 VP.n3 161.3
R24 VP.n19 VP.n18 161.3
R25 VP.n19 VP.n17 47.7732
R26 VP.n10 VP.n7 44.9377
R27 VP.n18 VP.n3 37.246
R28 VP.n30 VP.n29 37.246
R29 VP.n16 VP.n15 37.246
R30 VP.n23 VP.n22 28.4823
R31 VP.n28 VP.n1 28.4823
R32 VP.n14 VP.n13 28.4823
R33 VP.n9 VP.n8 28.4823
R34 VP.n24 VP.n23 19.7187
R35 VP.n24 VP.n1 19.7187
R36 VP.n13 VP.n6 19.7187
R37 VP.n9 VP.n6 19.7187
R38 VP.n8 VP.n7 17.0522
R39 VP.n22 VP.n3 10.955
R40 VP.n29 VP.n28 10.955
R41 VP.n15 VP.n14 10.955
R42 VP.n11 VP.n10 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n5 0.189894
R45 VP.n5 VP.n4 0.189894
R46 VP.n17 VP.n4 0.189894
R47 VP.n20 VP.n19 0.189894
R48 VP.n21 VP.n20 0.189894
R49 VP.n21 VP.n2 0.189894
R50 VP.n25 VP.n2 0.189894
R51 VP.n26 VP.n25 0.189894
R52 VP.n27 VP.n26 0.189894
R53 VP.n27 VP.n0 0.189894
R54 VP.n31 VP.n0 0.189894
R55 VP VP.n31 0.0516364
R56 VTAIL.n416 VTAIL.n320 756.745
R57 VTAIL.n98 VTAIL.n2 756.745
R58 VTAIL.n314 VTAIL.n218 756.745
R59 VTAIL.n208 VTAIL.n112 756.745
R60 VTAIL.n352 VTAIL.n351 585
R61 VTAIL.n357 VTAIL.n356 585
R62 VTAIL.n359 VTAIL.n358 585
R63 VTAIL.n348 VTAIL.n347 585
R64 VTAIL.n365 VTAIL.n364 585
R65 VTAIL.n367 VTAIL.n366 585
R66 VTAIL.n344 VTAIL.n343 585
R67 VTAIL.n373 VTAIL.n372 585
R68 VTAIL.n375 VTAIL.n374 585
R69 VTAIL.n340 VTAIL.n339 585
R70 VTAIL.n381 VTAIL.n380 585
R71 VTAIL.n383 VTAIL.n382 585
R72 VTAIL.n336 VTAIL.n335 585
R73 VTAIL.n389 VTAIL.n388 585
R74 VTAIL.n391 VTAIL.n390 585
R75 VTAIL.n332 VTAIL.n331 585
R76 VTAIL.n398 VTAIL.n397 585
R77 VTAIL.n399 VTAIL.n330 585
R78 VTAIL.n401 VTAIL.n400 585
R79 VTAIL.n328 VTAIL.n327 585
R80 VTAIL.n407 VTAIL.n406 585
R81 VTAIL.n409 VTAIL.n408 585
R82 VTAIL.n324 VTAIL.n323 585
R83 VTAIL.n415 VTAIL.n414 585
R84 VTAIL.n417 VTAIL.n416 585
R85 VTAIL.n34 VTAIL.n33 585
R86 VTAIL.n39 VTAIL.n38 585
R87 VTAIL.n41 VTAIL.n40 585
R88 VTAIL.n30 VTAIL.n29 585
R89 VTAIL.n47 VTAIL.n46 585
R90 VTAIL.n49 VTAIL.n48 585
R91 VTAIL.n26 VTAIL.n25 585
R92 VTAIL.n55 VTAIL.n54 585
R93 VTAIL.n57 VTAIL.n56 585
R94 VTAIL.n22 VTAIL.n21 585
R95 VTAIL.n63 VTAIL.n62 585
R96 VTAIL.n65 VTAIL.n64 585
R97 VTAIL.n18 VTAIL.n17 585
R98 VTAIL.n71 VTAIL.n70 585
R99 VTAIL.n73 VTAIL.n72 585
R100 VTAIL.n14 VTAIL.n13 585
R101 VTAIL.n80 VTAIL.n79 585
R102 VTAIL.n81 VTAIL.n12 585
R103 VTAIL.n83 VTAIL.n82 585
R104 VTAIL.n10 VTAIL.n9 585
R105 VTAIL.n89 VTAIL.n88 585
R106 VTAIL.n91 VTAIL.n90 585
R107 VTAIL.n6 VTAIL.n5 585
R108 VTAIL.n97 VTAIL.n96 585
R109 VTAIL.n99 VTAIL.n98 585
R110 VTAIL.n315 VTAIL.n314 585
R111 VTAIL.n313 VTAIL.n312 585
R112 VTAIL.n222 VTAIL.n221 585
R113 VTAIL.n307 VTAIL.n306 585
R114 VTAIL.n305 VTAIL.n304 585
R115 VTAIL.n226 VTAIL.n225 585
R116 VTAIL.n299 VTAIL.n298 585
R117 VTAIL.n297 VTAIL.n228 585
R118 VTAIL.n296 VTAIL.n295 585
R119 VTAIL.n231 VTAIL.n229 585
R120 VTAIL.n290 VTAIL.n289 585
R121 VTAIL.n288 VTAIL.n287 585
R122 VTAIL.n235 VTAIL.n234 585
R123 VTAIL.n282 VTAIL.n281 585
R124 VTAIL.n280 VTAIL.n279 585
R125 VTAIL.n239 VTAIL.n238 585
R126 VTAIL.n274 VTAIL.n273 585
R127 VTAIL.n272 VTAIL.n271 585
R128 VTAIL.n243 VTAIL.n242 585
R129 VTAIL.n266 VTAIL.n265 585
R130 VTAIL.n264 VTAIL.n263 585
R131 VTAIL.n247 VTAIL.n246 585
R132 VTAIL.n258 VTAIL.n257 585
R133 VTAIL.n256 VTAIL.n255 585
R134 VTAIL.n251 VTAIL.n250 585
R135 VTAIL.n209 VTAIL.n208 585
R136 VTAIL.n207 VTAIL.n206 585
R137 VTAIL.n116 VTAIL.n115 585
R138 VTAIL.n201 VTAIL.n200 585
R139 VTAIL.n199 VTAIL.n198 585
R140 VTAIL.n120 VTAIL.n119 585
R141 VTAIL.n193 VTAIL.n192 585
R142 VTAIL.n191 VTAIL.n122 585
R143 VTAIL.n190 VTAIL.n189 585
R144 VTAIL.n125 VTAIL.n123 585
R145 VTAIL.n184 VTAIL.n183 585
R146 VTAIL.n182 VTAIL.n181 585
R147 VTAIL.n129 VTAIL.n128 585
R148 VTAIL.n176 VTAIL.n175 585
R149 VTAIL.n174 VTAIL.n173 585
R150 VTAIL.n133 VTAIL.n132 585
R151 VTAIL.n168 VTAIL.n167 585
R152 VTAIL.n166 VTAIL.n165 585
R153 VTAIL.n137 VTAIL.n136 585
R154 VTAIL.n160 VTAIL.n159 585
R155 VTAIL.n158 VTAIL.n157 585
R156 VTAIL.n141 VTAIL.n140 585
R157 VTAIL.n152 VTAIL.n151 585
R158 VTAIL.n150 VTAIL.n149 585
R159 VTAIL.n145 VTAIL.n144 585
R160 VTAIL.n353 VTAIL.t4 327.466
R161 VTAIL.n35 VTAIL.t9 327.466
R162 VTAIL.n252 VTAIL.t13 327.466
R163 VTAIL.n146 VTAIL.t18 327.466
R164 VTAIL.n357 VTAIL.n351 171.744
R165 VTAIL.n358 VTAIL.n357 171.744
R166 VTAIL.n358 VTAIL.n347 171.744
R167 VTAIL.n365 VTAIL.n347 171.744
R168 VTAIL.n366 VTAIL.n365 171.744
R169 VTAIL.n366 VTAIL.n343 171.744
R170 VTAIL.n373 VTAIL.n343 171.744
R171 VTAIL.n374 VTAIL.n373 171.744
R172 VTAIL.n374 VTAIL.n339 171.744
R173 VTAIL.n381 VTAIL.n339 171.744
R174 VTAIL.n382 VTAIL.n381 171.744
R175 VTAIL.n382 VTAIL.n335 171.744
R176 VTAIL.n389 VTAIL.n335 171.744
R177 VTAIL.n390 VTAIL.n389 171.744
R178 VTAIL.n390 VTAIL.n331 171.744
R179 VTAIL.n398 VTAIL.n331 171.744
R180 VTAIL.n399 VTAIL.n398 171.744
R181 VTAIL.n400 VTAIL.n399 171.744
R182 VTAIL.n400 VTAIL.n327 171.744
R183 VTAIL.n407 VTAIL.n327 171.744
R184 VTAIL.n408 VTAIL.n407 171.744
R185 VTAIL.n408 VTAIL.n323 171.744
R186 VTAIL.n415 VTAIL.n323 171.744
R187 VTAIL.n416 VTAIL.n415 171.744
R188 VTAIL.n39 VTAIL.n33 171.744
R189 VTAIL.n40 VTAIL.n39 171.744
R190 VTAIL.n40 VTAIL.n29 171.744
R191 VTAIL.n47 VTAIL.n29 171.744
R192 VTAIL.n48 VTAIL.n47 171.744
R193 VTAIL.n48 VTAIL.n25 171.744
R194 VTAIL.n55 VTAIL.n25 171.744
R195 VTAIL.n56 VTAIL.n55 171.744
R196 VTAIL.n56 VTAIL.n21 171.744
R197 VTAIL.n63 VTAIL.n21 171.744
R198 VTAIL.n64 VTAIL.n63 171.744
R199 VTAIL.n64 VTAIL.n17 171.744
R200 VTAIL.n71 VTAIL.n17 171.744
R201 VTAIL.n72 VTAIL.n71 171.744
R202 VTAIL.n72 VTAIL.n13 171.744
R203 VTAIL.n80 VTAIL.n13 171.744
R204 VTAIL.n81 VTAIL.n80 171.744
R205 VTAIL.n82 VTAIL.n81 171.744
R206 VTAIL.n82 VTAIL.n9 171.744
R207 VTAIL.n89 VTAIL.n9 171.744
R208 VTAIL.n90 VTAIL.n89 171.744
R209 VTAIL.n90 VTAIL.n5 171.744
R210 VTAIL.n97 VTAIL.n5 171.744
R211 VTAIL.n98 VTAIL.n97 171.744
R212 VTAIL.n314 VTAIL.n313 171.744
R213 VTAIL.n313 VTAIL.n221 171.744
R214 VTAIL.n306 VTAIL.n221 171.744
R215 VTAIL.n306 VTAIL.n305 171.744
R216 VTAIL.n305 VTAIL.n225 171.744
R217 VTAIL.n298 VTAIL.n225 171.744
R218 VTAIL.n298 VTAIL.n297 171.744
R219 VTAIL.n297 VTAIL.n296 171.744
R220 VTAIL.n296 VTAIL.n229 171.744
R221 VTAIL.n289 VTAIL.n229 171.744
R222 VTAIL.n289 VTAIL.n288 171.744
R223 VTAIL.n288 VTAIL.n234 171.744
R224 VTAIL.n281 VTAIL.n234 171.744
R225 VTAIL.n281 VTAIL.n280 171.744
R226 VTAIL.n280 VTAIL.n238 171.744
R227 VTAIL.n273 VTAIL.n238 171.744
R228 VTAIL.n273 VTAIL.n272 171.744
R229 VTAIL.n272 VTAIL.n242 171.744
R230 VTAIL.n265 VTAIL.n242 171.744
R231 VTAIL.n265 VTAIL.n264 171.744
R232 VTAIL.n264 VTAIL.n246 171.744
R233 VTAIL.n257 VTAIL.n246 171.744
R234 VTAIL.n257 VTAIL.n256 171.744
R235 VTAIL.n256 VTAIL.n250 171.744
R236 VTAIL.n208 VTAIL.n207 171.744
R237 VTAIL.n207 VTAIL.n115 171.744
R238 VTAIL.n200 VTAIL.n115 171.744
R239 VTAIL.n200 VTAIL.n199 171.744
R240 VTAIL.n199 VTAIL.n119 171.744
R241 VTAIL.n192 VTAIL.n119 171.744
R242 VTAIL.n192 VTAIL.n191 171.744
R243 VTAIL.n191 VTAIL.n190 171.744
R244 VTAIL.n190 VTAIL.n123 171.744
R245 VTAIL.n183 VTAIL.n123 171.744
R246 VTAIL.n183 VTAIL.n182 171.744
R247 VTAIL.n182 VTAIL.n128 171.744
R248 VTAIL.n175 VTAIL.n128 171.744
R249 VTAIL.n175 VTAIL.n174 171.744
R250 VTAIL.n174 VTAIL.n132 171.744
R251 VTAIL.n167 VTAIL.n132 171.744
R252 VTAIL.n167 VTAIL.n166 171.744
R253 VTAIL.n166 VTAIL.n136 171.744
R254 VTAIL.n159 VTAIL.n136 171.744
R255 VTAIL.n159 VTAIL.n158 171.744
R256 VTAIL.n158 VTAIL.n140 171.744
R257 VTAIL.n151 VTAIL.n140 171.744
R258 VTAIL.n151 VTAIL.n150 171.744
R259 VTAIL.n150 VTAIL.n144 171.744
R260 VTAIL.t4 VTAIL.n351 85.8723
R261 VTAIL.t9 VTAIL.n33 85.8723
R262 VTAIL.t13 VTAIL.n250 85.8723
R263 VTAIL.t18 VTAIL.n144 85.8723
R264 VTAIL.n217 VTAIL.n216 53.1727
R265 VTAIL.n215 VTAIL.n214 53.1727
R266 VTAIL.n111 VTAIL.n110 53.1727
R267 VTAIL.n109 VTAIL.n108 53.1727
R268 VTAIL.n423 VTAIL.n422 53.1726
R269 VTAIL.n1 VTAIL.n0 53.1726
R270 VTAIL.n105 VTAIL.n104 53.1726
R271 VTAIL.n107 VTAIL.n106 53.1726
R272 VTAIL.n421 VTAIL.n420 33.349
R273 VTAIL.n103 VTAIL.n102 33.349
R274 VTAIL.n319 VTAIL.n318 33.349
R275 VTAIL.n213 VTAIL.n212 33.349
R276 VTAIL.n109 VTAIL.n107 29.9703
R277 VTAIL.n421 VTAIL.n319 29.0565
R278 VTAIL.n353 VTAIL.n352 16.3895
R279 VTAIL.n35 VTAIL.n34 16.3895
R280 VTAIL.n252 VTAIL.n251 16.3895
R281 VTAIL.n146 VTAIL.n145 16.3895
R282 VTAIL.n401 VTAIL.n330 13.1884
R283 VTAIL.n83 VTAIL.n12 13.1884
R284 VTAIL.n299 VTAIL.n228 13.1884
R285 VTAIL.n193 VTAIL.n122 13.1884
R286 VTAIL.n356 VTAIL.n355 12.8005
R287 VTAIL.n397 VTAIL.n396 12.8005
R288 VTAIL.n402 VTAIL.n328 12.8005
R289 VTAIL.n38 VTAIL.n37 12.8005
R290 VTAIL.n79 VTAIL.n78 12.8005
R291 VTAIL.n84 VTAIL.n10 12.8005
R292 VTAIL.n300 VTAIL.n226 12.8005
R293 VTAIL.n295 VTAIL.n230 12.8005
R294 VTAIL.n255 VTAIL.n254 12.8005
R295 VTAIL.n194 VTAIL.n120 12.8005
R296 VTAIL.n189 VTAIL.n124 12.8005
R297 VTAIL.n149 VTAIL.n148 12.8005
R298 VTAIL.n359 VTAIL.n350 12.0247
R299 VTAIL.n395 VTAIL.n332 12.0247
R300 VTAIL.n406 VTAIL.n405 12.0247
R301 VTAIL.n41 VTAIL.n32 12.0247
R302 VTAIL.n77 VTAIL.n14 12.0247
R303 VTAIL.n88 VTAIL.n87 12.0247
R304 VTAIL.n304 VTAIL.n303 12.0247
R305 VTAIL.n294 VTAIL.n231 12.0247
R306 VTAIL.n258 VTAIL.n249 12.0247
R307 VTAIL.n198 VTAIL.n197 12.0247
R308 VTAIL.n188 VTAIL.n125 12.0247
R309 VTAIL.n152 VTAIL.n143 12.0247
R310 VTAIL.n360 VTAIL.n348 11.249
R311 VTAIL.n392 VTAIL.n391 11.249
R312 VTAIL.n409 VTAIL.n326 11.249
R313 VTAIL.n42 VTAIL.n30 11.249
R314 VTAIL.n74 VTAIL.n73 11.249
R315 VTAIL.n91 VTAIL.n8 11.249
R316 VTAIL.n307 VTAIL.n224 11.249
R317 VTAIL.n291 VTAIL.n290 11.249
R318 VTAIL.n259 VTAIL.n247 11.249
R319 VTAIL.n201 VTAIL.n118 11.249
R320 VTAIL.n185 VTAIL.n184 11.249
R321 VTAIL.n153 VTAIL.n141 11.249
R322 VTAIL.n364 VTAIL.n363 10.4732
R323 VTAIL.n388 VTAIL.n334 10.4732
R324 VTAIL.n410 VTAIL.n324 10.4732
R325 VTAIL.n46 VTAIL.n45 10.4732
R326 VTAIL.n70 VTAIL.n16 10.4732
R327 VTAIL.n92 VTAIL.n6 10.4732
R328 VTAIL.n308 VTAIL.n222 10.4732
R329 VTAIL.n287 VTAIL.n233 10.4732
R330 VTAIL.n263 VTAIL.n262 10.4732
R331 VTAIL.n202 VTAIL.n116 10.4732
R332 VTAIL.n181 VTAIL.n127 10.4732
R333 VTAIL.n157 VTAIL.n156 10.4732
R334 VTAIL.n367 VTAIL.n346 9.69747
R335 VTAIL.n387 VTAIL.n336 9.69747
R336 VTAIL.n414 VTAIL.n413 9.69747
R337 VTAIL.n49 VTAIL.n28 9.69747
R338 VTAIL.n69 VTAIL.n18 9.69747
R339 VTAIL.n96 VTAIL.n95 9.69747
R340 VTAIL.n312 VTAIL.n311 9.69747
R341 VTAIL.n286 VTAIL.n235 9.69747
R342 VTAIL.n266 VTAIL.n245 9.69747
R343 VTAIL.n206 VTAIL.n205 9.69747
R344 VTAIL.n180 VTAIL.n129 9.69747
R345 VTAIL.n160 VTAIL.n139 9.69747
R346 VTAIL.n420 VTAIL.n419 9.45567
R347 VTAIL.n102 VTAIL.n101 9.45567
R348 VTAIL.n318 VTAIL.n317 9.45567
R349 VTAIL.n212 VTAIL.n211 9.45567
R350 VTAIL.n419 VTAIL.n418 9.3005
R351 VTAIL.n322 VTAIL.n321 9.3005
R352 VTAIL.n413 VTAIL.n412 9.3005
R353 VTAIL.n411 VTAIL.n410 9.3005
R354 VTAIL.n326 VTAIL.n325 9.3005
R355 VTAIL.n405 VTAIL.n404 9.3005
R356 VTAIL.n403 VTAIL.n402 9.3005
R357 VTAIL.n342 VTAIL.n341 9.3005
R358 VTAIL.n371 VTAIL.n370 9.3005
R359 VTAIL.n369 VTAIL.n368 9.3005
R360 VTAIL.n346 VTAIL.n345 9.3005
R361 VTAIL.n363 VTAIL.n362 9.3005
R362 VTAIL.n361 VTAIL.n360 9.3005
R363 VTAIL.n350 VTAIL.n349 9.3005
R364 VTAIL.n355 VTAIL.n354 9.3005
R365 VTAIL.n377 VTAIL.n376 9.3005
R366 VTAIL.n379 VTAIL.n378 9.3005
R367 VTAIL.n338 VTAIL.n337 9.3005
R368 VTAIL.n385 VTAIL.n384 9.3005
R369 VTAIL.n387 VTAIL.n386 9.3005
R370 VTAIL.n334 VTAIL.n333 9.3005
R371 VTAIL.n393 VTAIL.n392 9.3005
R372 VTAIL.n395 VTAIL.n394 9.3005
R373 VTAIL.n396 VTAIL.n329 9.3005
R374 VTAIL.n101 VTAIL.n100 9.3005
R375 VTAIL.n4 VTAIL.n3 9.3005
R376 VTAIL.n95 VTAIL.n94 9.3005
R377 VTAIL.n93 VTAIL.n92 9.3005
R378 VTAIL.n8 VTAIL.n7 9.3005
R379 VTAIL.n87 VTAIL.n86 9.3005
R380 VTAIL.n85 VTAIL.n84 9.3005
R381 VTAIL.n24 VTAIL.n23 9.3005
R382 VTAIL.n53 VTAIL.n52 9.3005
R383 VTAIL.n51 VTAIL.n50 9.3005
R384 VTAIL.n28 VTAIL.n27 9.3005
R385 VTAIL.n45 VTAIL.n44 9.3005
R386 VTAIL.n43 VTAIL.n42 9.3005
R387 VTAIL.n32 VTAIL.n31 9.3005
R388 VTAIL.n37 VTAIL.n36 9.3005
R389 VTAIL.n59 VTAIL.n58 9.3005
R390 VTAIL.n61 VTAIL.n60 9.3005
R391 VTAIL.n20 VTAIL.n19 9.3005
R392 VTAIL.n67 VTAIL.n66 9.3005
R393 VTAIL.n69 VTAIL.n68 9.3005
R394 VTAIL.n16 VTAIL.n15 9.3005
R395 VTAIL.n75 VTAIL.n74 9.3005
R396 VTAIL.n77 VTAIL.n76 9.3005
R397 VTAIL.n78 VTAIL.n11 9.3005
R398 VTAIL.n278 VTAIL.n277 9.3005
R399 VTAIL.n237 VTAIL.n236 9.3005
R400 VTAIL.n284 VTAIL.n283 9.3005
R401 VTAIL.n286 VTAIL.n285 9.3005
R402 VTAIL.n233 VTAIL.n232 9.3005
R403 VTAIL.n292 VTAIL.n291 9.3005
R404 VTAIL.n294 VTAIL.n293 9.3005
R405 VTAIL.n230 VTAIL.n227 9.3005
R406 VTAIL.n317 VTAIL.n316 9.3005
R407 VTAIL.n220 VTAIL.n219 9.3005
R408 VTAIL.n311 VTAIL.n310 9.3005
R409 VTAIL.n309 VTAIL.n308 9.3005
R410 VTAIL.n224 VTAIL.n223 9.3005
R411 VTAIL.n303 VTAIL.n302 9.3005
R412 VTAIL.n301 VTAIL.n300 9.3005
R413 VTAIL.n276 VTAIL.n275 9.3005
R414 VTAIL.n241 VTAIL.n240 9.3005
R415 VTAIL.n270 VTAIL.n269 9.3005
R416 VTAIL.n268 VTAIL.n267 9.3005
R417 VTAIL.n245 VTAIL.n244 9.3005
R418 VTAIL.n262 VTAIL.n261 9.3005
R419 VTAIL.n260 VTAIL.n259 9.3005
R420 VTAIL.n249 VTAIL.n248 9.3005
R421 VTAIL.n254 VTAIL.n253 9.3005
R422 VTAIL.n172 VTAIL.n171 9.3005
R423 VTAIL.n131 VTAIL.n130 9.3005
R424 VTAIL.n178 VTAIL.n177 9.3005
R425 VTAIL.n180 VTAIL.n179 9.3005
R426 VTAIL.n127 VTAIL.n126 9.3005
R427 VTAIL.n186 VTAIL.n185 9.3005
R428 VTAIL.n188 VTAIL.n187 9.3005
R429 VTAIL.n124 VTAIL.n121 9.3005
R430 VTAIL.n211 VTAIL.n210 9.3005
R431 VTAIL.n114 VTAIL.n113 9.3005
R432 VTAIL.n205 VTAIL.n204 9.3005
R433 VTAIL.n203 VTAIL.n202 9.3005
R434 VTAIL.n118 VTAIL.n117 9.3005
R435 VTAIL.n197 VTAIL.n196 9.3005
R436 VTAIL.n195 VTAIL.n194 9.3005
R437 VTAIL.n170 VTAIL.n169 9.3005
R438 VTAIL.n135 VTAIL.n134 9.3005
R439 VTAIL.n164 VTAIL.n163 9.3005
R440 VTAIL.n162 VTAIL.n161 9.3005
R441 VTAIL.n139 VTAIL.n138 9.3005
R442 VTAIL.n156 VTAIL.n155 9.3005
R443 VTAIL.n154 VTAIL.n153 9.3005
R444 VTAIL.n143 VTAIL.n142 9.3005
R445 VTAIL.n148 VTAIL.n147 9.3005
R446 VTAIL.n368 VTAIL.n344 8.92171
R447 VTAIL.n384 VTAIL.n383 8.92171
R448 VTAIL.n417 VTAIL.n322 8.92171
R449 VTAIL.n50 VTAIL.n26 8.92171
R450 VTAIL.n66 VTAIL.n65 8.92171
R451 VTAIL.n99 VTAIL.n4 8.92171
R452 VTAIL.n315 VTAIL.n220 8.92171
R453 VTAIL.n283 VTAIL.n282 8.92171
R454 VTAIL.n267 VTAIL.n243 8.92171
R455 VTAIL.n209 VTAIL.n114 8.92171
R456 VTAIL.n177 VTAIL.n176 8.92171
R457 VTAIL.n161 VTAIL.n137 8.92171
R458 VTAIL.n372 VTAIL.n371 8.14595
R459 VTAIL.n380 VTAIL.n338 8.14595
R460 VTAIL.n418 VTAIL.n320 8.14595
R461 VTAIL.n54 VTAIL.n53 8.14595
R462 VTAIL.n62 VTAIL.n20 8.14595
R463 VTAIL.n100 VTAIL.n2 8.14595
R464 VTAIL.n316 VTAIL.n218 8.14595
R465 VTAIL.n279 VTAIL.n237 8.14595
R466 VTAIL.n271 VTAIL.n270 8.14595
R467 VTAIL.n210 VTAIL.n112 8.14595
R468 VTAIL.n173 VTAIL.n131 8.14595
R469 VTAIL.n165 VTAIL.n164 8.14595
R470 VTAIL.n375 VTAIL.n342 7.3702
R471 VTAIL.n379 VTAIL.n340 7.3702
R472 VTAIL.n57 VTAIL.n24 7.3702
R473 VTAIL.n61 VTAIL.n22 7.3702
R474 VTAIL.n278 VTAIL.n239 7.3702
R475 VTAIL.n274 VTAIL.n241 7.3702
R476 VTAIL.n172 VTAIL.n133 7.3702
R477 VTAIL.n168 VTAIL.n135 7.3702
R478 VTAIL.n376 VTAIL.n375 6.59444
R479 VTAIL.n376 VTAIL.n340 6.59444
R480 VTAIL.n58 VTAIL.n57 6.59444
R481 VTAIL.n58 VTAIL.n22 6.59444
R482 VTAIL.n275 VTAIL.n239 6.59444
R483 VTAIL.n275 VTAIL.n274 6.59444
R484 VTAIL.n169 VTAIL.n133 6.59444
R485 VTAIL.n169 VTAIL.n168 6.59444
R486 VTAIL.n372 VTAIL.n342 5.81868
R487 VTAIL.n380 VTAIL.n379 5.81868
R488 VTAIL.n420 VTAIL.n320 5.81868
R489 VTAIL.n54 VTAIL.n24 5.81868
R490 VTAIL.n62 VTAIL.n61 5.81868
R491 VTAIL.n102 VTAIL.n2 5.81868
R492 VTAIL.n318 VTAIL.n218 5.81868
R493 VTAIL.n279 VTAIL.n278 5.81868
R494 VTAIL.n271 VTAIL.n241 5.81868
R495 VTAIL.n212 VTAIL.n112 5.81868
R496 VTAIL.n173 VTAIL.n172 5.81868
R497 VTAIL.n165 VTAIL.n135 5.81868
R498 VTAIL.n371 VTAIL.n344 5.04292
R499 VTAIL.n383 VTAIL.n338 5.04292
R500 VTAIL.n418 VTAIL.n417 5.04292
R501 VTAIL.n53 VTAIL.n26 5.04292
R502 VTAIL.n65 VTAIL.n20 5.04292
R503 VTAIL.n100 VTAIL.n99 5.04292
R504 VTAIL.n316 VTAIL.n315 5.04292
R505 VTAIL.n282 VTAIL.n237 5.04292
R506 VTAIL.n270 VTAIL.n243 5.04292
R507 VTAIL.n210 VTAIL.n209 5.04292
R508 VTAIL.n176 VTAIL.n131 5.04292
R509 VTAIL.n164 VTAIL.n137 5.04292
R510 VTAIL.n368 VTAIL.n367 4.26717
R511 VTAIL.n384 VTAIL.n336 4.26717
R512 VTAIL.n414 VTAIL.n322 4.26717
R513 VTAIL.n50 VTAIL.n49 4.26717
R514 VTAIL.n66 VTAIL.n18 4.26717
R515 VTAIL.n96 VTAIL.n4 4.26717
R516 VTAIL.n312 VTAIL.n220 4.26717
R517 VTAIL.n283 VTAIL.n235 4.26717
R518 VTAIL.n267 VTAIL.n266 4.26717
R519 VTAIL.n206 VTAIL.n114 4.26717
R520 VTAIL.n177 VTAIL.n129 4.26717
R521 VTAIL.n161 VTAIL.n160 4.26717
R522 VTAIL.n354 VTAIL.n353 3.70982
R523 VTAIL.n36 VTAIL.n35 3.70982
R524 VTAIL.n253 VTAIL.n252 3.70982
R525 VTAIL.n147 VTAIL.n146 3.70982
R526 VTAIL.n364 VTAIL.n346 3.49141
R527 VTAIL.n388 VTAIL.n387 3.49141
R528 VTAIL.n413 VTAIL.n324 3.49141
R529 VTAIL.n46 VTAIL.n28 3.49141
R530 VTAIL.n70 VTAIL.n69 3.49141
R531 VTAIL.n95 VTAIL.n6 3.49141
R532 VTAIL.n311 VTAIL.n222 3.49141
R533 VTAIL.n287 VTAIL.n286 3.49141
R534 VTAIL.n263 VTAIL.n245 3.49141
R535 VTAIL.n205 VTAIL.n116 3.49141
R536 VTAIL.n181 VTAIL.n180 3.49141
R537 VTAIL.n157 VTAIL.n139 3.49141
R538 VTAIL.n363 VTAIL.n348 2.71565
R539 VTAIL.n391 VTAIL.n334 2.71565
R540 VTAIL.n410 VTAIL.n409 2.71565
R541 VTAIL.n45 VTAIL.n30 2.71565
R542 VTAIL.n73 VTAIL.n16 2.71565
R543 VTAIL.n92 VTAIL.n91 2.71565
R544 VTAIL.n308 VTAIL.n307 2.71565
R545 VTAIL.n290 VTAIL.n233 2.71565
R546 VTAIL.n262 VTAIL.n247 2.71565
R547 VTAIL.n202 VTAIL.n201 2.71565
R548 VTAIL.n184 VTAIL.n127 2.71565
R549 VTAIL.n156 VTAIL.n141 2.71565
R550 VTAIL.n360 VTAIL.n359 1.93989
R551 VTAIL.n392 VTAIL.n332 1.93989
R552 VTAIL.n406 VTAIL.n326 1.93989
R553 VTAIL.n42 VTAIL.n41 1.93989
R554 VTAIL.n74 VTAIL.n14 1.93989
R555 VTAIL.n88 VTAIL.n8 1.93989
R556 VTAIL.n304 VTAIL.n224 1.93989
R557 VTAIL.n291 VTAIL.n231 1.93989
R558 VTAIL.n259 VTAIL.n258 1.93989
R559 VTAIL.n198 VTAIL.n118 1.93989
R560 VTAIL.n185 VTAIL.n125 1.93989
R561 VTAIL.n153 VTAIL.n152 1.93989
R562 VTAIL.n422 VTAIL.t6 1.77673
R563 VTAIL.n422 VTAIL.t2 1.77673
R564 VTAIL.n0 VTAIL.t0 1.77673
R565 VTAIL.n0 VTAIL.t1 1.77673
R566 VTAIL.n104 VTAIL.t8 1.77673
R567 VTAIL.n104 VTAIL.t14 1.77673
R568 VTAIL.n106 VTAIL.t16 1.77673
R569 VTAIL.n106 VTAIL.t10 1.77673
R570 VTAIL.n216 VTAIL.t17 1.77673
R571 VTAIL.n216 VTAIL.t12 1.77673
R572 VTAIL.n214 VTAIL.t11 1.77673
R573 VTAIL.n214 VTAIL.t15 1.77673
R574 VTAIL.n110 VTAIL.t19 1.77673
R575 VTAIL.n110 VTAIL.t5 1.77673
R576 VTAIL.n108 VTAIL.t3 1.77673
R577 VTAIL.n108 VTAIL.t7 1.77673
R578 VTAIL.n356 VTAIL.n350 1.16414
R579 VTAIL.n397 VTAIL.n395 1.16414
R580 VTAIL.n405 VTAIL.n328 1.16414
R581 VTAIL.n38 VTAIL.n32 1.16414
R582 VTAIL.n79 VTAIL.n77 1.16414
R583 VTAIL.n87 VTAIL.n10 1.16414
R584 VTAIL.n303 VTAIL.n226 1.16414
R585 VTAIL.n295 VTAIL.n294 1.16414
R586 VTAIL.n255 VTAIL.n249 1.16414
R587 VTAIL.n197 VTAIL.n120 1.16414
R588 VTAIL.n189 VTAIL.n188 1.16414
R589 VTAIL.n149 VTAIL.n143 1.16414
R590 VTAIL.n215 VTAIL.n213 0.927224
R591 VTAIL.n103 VTAIL.n1 0.927224
R592 VTAIL.n111 VTAIL.n109 0.914293
R593 VTAIL.n213 VTAIL.n111 0.914293
R594 VTAIL.n217 VTAIL.n215 0.914293
R595 VTAIL.n319 VTAIL.n217 0.914293
R596 VTAIL.n107 VTAIL.n105 0.914293
R597 VTAIL.n105 VTAIL.n103 0.914293
R598 VTAIL.n423 VTAIL.n421 0.914293
R599 VTAIL VTAIL.n1 0.744035
R600 VTAIL.n355 VTAIL.n352 0.388379
R601 VTAIL.n396 VTAIL.n330 0.388379
R602 VTAIL.n402 VTAIL.n401 0.388379
R603 VTAIL.n37 VTAIL.n34 0.388379
R604 VTAIL.n78 VTAIL.n12 0.388379
R605 VTAIL.n84 VTAIL.n83 0.388379
R606 VTAIL.n300 VTAIL.n299 0.388379
R607 VTAIL.n230 VTAIL.n228 0.388379
R608 VTAIL.n254 VTAIL.n251 0.388379
R609 VTAIL.n194 VTAIL.n193 0.388379
R610 VTAIL.n124 VTAIL.n122 0.388379
R611 VTAIL.n148 VTAIL.n145 0.388379
R612 VTAIL VTAIL.n423 0.170759
R613 VTAIL.n354 VTAIL.n349 0.155672
R614 VTAIL.n361 VTAIL.n349 0.155672
R615 VTAIL.n362 VTAIL.n361 0.155672
R616 VTAIL.n362 VTAIL.n345 0.155672
R617 VTAIL.n369 VTAIL.n345 0.155672
R618 VTAIL.n370 VTAIL.n369 0.155672
R619 VTAIL.n370 VTAIL.n341 0.155672
R620 VTAIL.n377 VTAIL.n341 0.155672
R621 VTAIL.n378 VTAIL.n377 0.155672
R622 VTAIL.n378 VTAIL.n337 0.155672
R623 VTAIL.n385 VTAIL.n337 0.155672
R624 VTAIL.n386 VTAIL.n385 0.155672
R625 VTAIL.n386 VTAIL.n333 0.155672
R626 VTAIL.n393 VTAIL.n333 0.155672
R627 VTAIL.n394 VTAIL.n393 0.155672
R628 VTAIL.n394 VTAIL.n329 0.155672
R629 VTAIL.n403 VTAIL.n329 0.155672
R630 VTAIL.n404 VTAIL.n403 0.155672
R631 VTAIL.n404 VTAIL.n325 0.155672
R632 VTAIL.n411 VTAIL.n325 0.155672
R633 VTAIL.n412 VTAIL.n411 0.155672
R634 VTAIL.n412 VTAIL.n321 0.155672
R635 VTAIL.n419 VTAIL.n321 0.155672
R636 VTAIL.n36 VTAIL.n31 0.155672
R637 VTAIL.n43 VTAIL.n31 0.155672
R638 VTAIL.n44 VTAIL.n43 0.155672
R639 VTAIL.n44 VTAIL.n27 0.155672
R640 VTAIL.n51 VTAIL.n27 0.155672
R641 VTAIL.n52 VTAIL.n51 0.155672
R642 VTAIL.n52 VTAIL.n23 0.155672
R643 VTAIL.n59 VTAIL.n23 0.155672
R644 VTAIL.n60 VTAIL.n59 0.155672
R645 VTAIL.n60 VTAIL.n19 0.155672
R646 VTAIL.n67 VTAIL.n19 0.155672
R647 VTAIL.n68 VTAIL.n67 0.155672
R648 VTAIL.n68 VTAIL.n15 0.155672
R649 VTAIL.n75 VTAIL.n15 0.155672
R650 VTAIL.n76 VTAIL.n75 0.155672
R651 VTAIL.n76 VTAIL.n11 0.155672
R652 VTAIL.n85 VTAIL.n11 0.155672
R653 VTAIL.n86 VTAIL.n85 0.155672
R654 VTAIL.n86 VTAIL.n7 0.155672
R655 VTAIL.n93 VTAIL.n7 0.155672
R656 VTAIL.n94 VTAIL.n93 0.155672
R657 VTAIL.n94 VTAIL.n3 0.155672
R658 VTAIL.n101 VTAIL.n3 0.155672
R659 VTAIL.n317 VTAIL.n219 0.155672
R660 VTAIL.n310 VTAIL.n219 0.155672
R661 VTAIL.n310 VTAIL.n309 0.155672
R662 VTAIL.n309 VTAIL.n223 0.155672
R663 VTAIL.n302 VTAIL.n223 0.155672
R664 VTAIL.n302 VTAIL.n301 0.155672
R665 VTAIL.n301 VTAIL.n227 0.155672
R666 VTAIL.n293 VTAIL.n227 0.155672
R667 VTAIL.n293 VTAIL.n292 0.155672
R668 VTAIL.n292 VTAIL.n232 0.155672
R669 VTAIL.n285 VTAIL.n232 0.155672
R670 VTAIL.n285 VTAIL.n284 0.155672
R671 VTAIL.n284 VTAIL.n236 0.155672
R672 VTAIL.n277 VTAIL.n236 0.155672
R673 VTAIL.n277 VTAIL.n276 0.155672
R674 VTAIL.n276 VTAIL.n240 0.155672
R675 VTAIL.n269 VTAIL.n240 0.155672
R676 VTAIL.n269 VTAIL.n268 0.155672
R677 VTAIL.n268 VTAIL.n244 0.155672
R678 VTAIL.n261 VTAIL.n244 0.155672
R679 VTAIL.n261 VTAIL.n260 0.155672
R680 VTAIL.n260 VTAIL.n248 0.155672
R681 VTAIL.n253 VTAIL.n248 0.155672
R682 VTAIL.n211 VTAIL.n113 0.155672
R683 VTAIL.n204 VTAIL.n113 0.155672
R684 VTAIL.n204 VTAIL.n203 0.155672
R685 VTAIL.n203 VTAIL.n117 0.155672
R686 VTAIL.n196 VTAIL.n117 0.155672
R687 VTAIL.n196 VTAIL.n195 0.155672
R688 VTAIL.n195 VTAIL.n121 0.155672
R689 VTAIL.n187 VTAIL.n121 0.155672
R690 VTAIL.n187 VTAIL.n186 0.155672
R691 VTAIL.n186 VTAIL.n126 0.155672
R692 VTAIL.n179 VTAIL.n126 0.155672
R693 VTAIL.n179 VTAIL.n178 0.155672
R694 VTAIL.n178 VTAIL.n130 0.155672
R695 VTAIL.n171 VTAIL.n130 0.155672
R696 VTAIL.n171 VTAIL.n170 0.155672
R697 VTAIL.n170 VTAIL.n134 0.155672
R698 VTAIL.n163 VTAIL.n134 0.155672
R699 VTAIL.n163 VTAIL.n162 0.155672
R700 VTAIL.n162 VTAIL.n138 0.155672
R701 VTAIL.n155 VTAIL.n138 0.155672
R702 VTAIL.n155 VTAIL.n154 0.155672
R703 VTAIL.n154 VTAIL.n142 0.155672
R704 VTAIL.n147 VTAIL.n142 0.155672
R705 VDD1.n96 VDD1.n0 756.745
R706 VDD1.n199 VDD1.n103 756.745
R707 VDD1.n97 VDD1.n96 585
R708 VDD1.n95 VDD1.n94 585
R709 VDD1.n4 VDD1.n3 585
R710 VDD1.n89 VDD1.n88 585
R711 VDD1.n87 VDD1.n86 585
R712 VDD1.n8 VDD1.n7 585
R713 VDD1.n81 VDD1.n80 585
R714 VDD1.n79 VDD1.n10 585
R715 VDD1.n78 VDD1.n77 585
R716 VDD1.n13 VDD1.n11 585
R717 VDD1.n72 VDD1.n71 585
R718 VDD1.n70 VDD1.n69 585
R719 VDD1.n17 VDD1.n16 585
R720 VDD1.n64 VDD1.n63 585
R721 VDD1.n62 VDD1.n61 585
R722 VDD1.n21 VDD1.n20 585
R723 VDD1.n56 VDD1.n55 585
R724 VDD1.n54 VDD1.n53 585
R725 VDD1.n25 VDD1.n24 585
R726 VDD1.n48 VDD1.n47 585
R727 VDD1.n46 VDD1.n45 585
R728 VDD1.n29 VDD1.n28 585
R729 VDD1.n40 VDD1.n39 585
R730 VDD1.n38 VDD1.n37 585
R731 VDD1.n33 VDD1.n32 585
R732 VDD1.n135 VDD1.n134 585
R733 VDD1.n140 VDD1.n139 585
R734 VDD1.n142 VDD1.n141 585
R735 VDD1.n131 VDD1.n130 585
R736 VDD1.n148 VDD1.n147 585
R737 VDD1.n150 VDD1.n149 585
R738 VDD1.n127 VDD1.n126 585
R739 VDD1.n156 VDD1.n155 585
R740 VDD1.n158 VDD1.n157 585
R741 VDD1.n123 VDD1.n122 585
R742 VDD1.n164 VDD1.n163 585
R743 VDD1.n166 VDD1.n165 585
R744 VDD1.n119 VDD1.n118 585
R745 VDD1.n172 VDD1.n171 585
R746 VDD1.n174 VDD1.n173 585
R747 VDD1.n115 VDD1.n114 585
R748 VDD1.n181 VDD1.n180 585
R749 VDD1.n182 VDD1.n113 585
R750 VDD1.n184 VDD1.n183 585
R751 VDD1.n111 VDD1.n110 585
R752 VDD1.n190 VDD1.n189 585
R753 VDD1.n192 VDD1.n191 585
R754 VDD1.n107 VDD1.n106 585
R755 VDD1.n198 VDD1.n197 585
R756 VDD1.n200 VDD1.n199 585
R757 VDD1.n34 VDD1.t9 327.466
R758 VDD1.n136 VDD1.t5 327.466
R759 VDD1.n96 VDD1.n95 171.744
R760 VDD1.n95 VDD1.n3 171.744
R761 VDD1.n88 VDD1.n3 171.744
R762 VDD1.n88 VDD1.n87 171.744
R763 VDD1.n87 VDD1.n7 171.744
R764 VDD1.n80 VDD1.n7 171.744
R765 VDD1.n80 VDD1.n79 171.744
R766 VDD1.n79 VDD1.n78 171.744
R767 VDD1.n78 VDD1.n11 171.744
R768 VDD1.n71 VDD1.n11 171.744
R769 VDD1.n71 VDD1.n70 171.744
R770 VDD1.n70 VDD1.n16 171.744
R771 VDD1.n63 VDD1.n16 171.744
R772 VDD1.n63 VDD1.n62 171.744
R773 VDD1.n62 VDD1.n20 171.744
R774 VDD1.n55 VDD1.n20 171.744
R775 VDD1.n55 VDD1.n54 171.744
R776 VDD1.n54 VDD1.n24 171.744
R777 VDD1.n47 VDD1.n24 171.744
R778 VDD1.n47 VDD1.n46 171.744
R779 VDD1.n46 VDD1.n28 171.744
R780 VDD1.n39 VDD1.n28 171.744
R781 VDD1.n39 VDD1.n38 171.744
R782 VDD1.n38 VDD1.n32 171.744
R783 VDD1.n140 VDD1.n134 171.744
R784 VDD1.n141 VDD1.n140 171.744
R785 VDD1.n141 VDD1.n130 171.744
R786 VDD1.n148 VDD1.n130 171.744
R787 VDD1.n149 VDD1.n148 171.744
R788 VDD1.n149 VDD1.n126 171.744
R789 VDD1.n156 VDD1.n126 171.744
R790 VDD1.n157 VDD1.n156 171.744
R791 VDD1.n157 VDD1.n122 171.744
R792 VDD1.n164 VDD1.n122 171.744
R793 VDD1.n165 VDD1.n164 171.744
R794 VDD1.n165 VDD1.n118 171.744
R795 VDD1.n172 VDD1.n118 171.744
R796 VDD1.n173 VDD1.n172 171.744
R797 VDD1.n173 VDD1.n114 171.744
R798 VDD1.n181 VDD1.n114 171.744
R799 VDD1.n182 VDD1.n181 171.744
R800 VDD1.n183 VDD1.n182 171.744
R801 VDD1.n183 VDD1.n110 171.744
R802 VDD1.n190 VDD1.n110 171.744
R803 VDD1.n191 VDD1.n190 171.744
R804 VDD1.n191 VDD1.n106 171.744
R805 VDD1.n198 VDD1.n106 171.744
R806 VDD1.n199 VDD1.n198 171.744
R807 VDD1.t9 VDD1.n32 85.8723
R808 VDD1.t5 VDD1.n134 85.8723
R809 VDD1.n207 VDD1.n206 70.4813
R810 VDD1.n102 VDD1.n101 69.8515
R811 VDD1.n209 VDD1.n208 69.8513
R812 VDD1.n205 VDD1.n204 69.8513
R813 VDD1.n102 VDD1.n100 50.9416
R814 VDD1.n205 VDD1.n203 50.9416
R815 VDD1.n209 VDD1.n207 44.8716
R816 VDD1.n34 VDD1.n33 16.3895
R817 VDD1.n136 VDD1.n135 16.3895
R818 VDD1.n81 VDD1.n10 13.1884
R819 VDD1.n184 VDD1.n113 13.1884
R820 VDD1.n82 VDD1.n8 12.8005
R821 VDD1.n77 VDD1.n12 12.8005
R822 VDD1.n37 VDD1.n36 12.8005
R823 VDD1.n139 VDD1.n138 12.8005
R824 VDD1.n180 VDD1.n179 12.8005
R825 VDD1.n185 VDD1.n111 12.8005
R826 VDD1.n86 VDD1.n85 12.0247
R827 VDD1.n76 VDD1.n13 12.0247
R828 VDD1.n40 VDD1.n31 12.0247
R829 VDD1.n142 VDD1.n133 12.0247
R830 VDD1.n178 VDD1.n115 12.0247
R831 VDD1.n189 VDD1.n188 12.0247
R832 VDD1.n89 VDD1.n6 11.249
R833 VDD1.n73 VDD1.n72 11.249
R834 VDD1.n41 VDD1.n29 11.249
R835 VDD1.n143 VDD1.n131 11.249
R836 VDD1.n175 VDD1.n174 11.249
R837 VDD1.n192 VDD1.n109 11.249
R838 VDD1.n90 VDD1.n4 10.4732
R839 VDD1.n69 VDD1.n15 10.4732
R840 VDD1.n45 VDD1.n44 10.4732
R841 VDD1.n147 VDD1.n146 10.4732
R842 VDD1.n171 VDD1.n117 10.4732
R843 VDD1.n193 VDD1.n107 10.4732
R844 VDD1.n94 VDD1.n93 9.69747
R845 VDD1.n68 VDD1.n17 9.69747
R846 VDD1.n48 VDD1.n27 9.69747
R847 VDD1.n150 VDD1.n129 9.69747
R848 VDD1.n170 VDD1.n119 9.69747
R849 VDD1.n197 VDD1.n196 9.69747
R850 VDD1.n100 VDD1.n99 9.45567
R851 VDD1.n203 VDD1.n202 9.45567
R852 VDD1.n60 VDD1.n59 9.3005
R853 VDD1.n19 VDD1.n18 9.3005
R854 VDD1.n66 VDD1.n65 9.3005
R855 VDD1.n68 VDD1.n67 9.3005
R856 VDD1.n15 VDD1.n14 9.3005
R857 VDD1.n74 VDD1.n73 9.3005
R858 VDD1.n76 VDD1.n75 9.3005
R859 VDD1.n12 VDD1.n9 9.3005
R860 VDD1.n99 VDD1.n98 9.3005
R861 VDD1.n2 VDD1.n1 9.3005
R862 VDD1.n93 VDD1.n92 9.3005
R863 VDD1.n91 VDD1.n90 9.3005
R864 VDD1.n6 VDD1.n5 9.3005
R865 VDD1.n85 VDD1.n84 9.3005
R866 VDD1.n83 VDD1.n82 9.3005
R867 VDD1.n58 VDD1.n57 9.3005
R868 VDD1.n23 VDD1.n22 9.3005
R869 VDD1.n52 VDD1.n51 9.3005
R870 VDD1.n50 VDD1.n49 9.3005
R871 VDD1.n27 VDD1.n26 9.3005
R872 VDD1.n44 VDD1.n43 9.3005
R873 VDD1.n42 VDD1.n41 9.3005
R874 VDD1.n31 VDD1.n30 9.3005
R875 VDD1.n36 VDD1.n35 9.3005
R876 VDD1.n202 VDD1.n201 9.3005
R877 VDD1.n105 VDD1.n104 9.3005
R878 VDD1.n196 VDD1.n195 9.3005
R879 VDD1.n194 VDD1.n193 9.3005
R880 VDD1.n109 VDD1.n108 9.3005
R881 VDD1.n188 VDD1.n187 9.3005
R882 VDD1.n186 VDD1.n185 9.3005
R883 VDD1.n125 VDD1.n124 9.3005
R884 VDD1.n154 VDD1.n153 9.3005
R885 VDD1.n152 VDD1.n151 9.3005
R886 VDD1.n129 VDD1.n128 9.3005
R887 VDD1.n146 VDD1.n145 9.3005
R888 VDD1.n144 VDD1.n143 9.3005
R889 VDD1.n133 VDD1.n132 9.3005
R890 VDD1.n138 VDD1.n137 9.3005
R891 VDD1.n160 VDD1.n159 9.3005
R892 VDD1.n162 VDD1.n161 9.3005
R893 VDD1.n121 VDD1.n120 9.3005
R894 VDD1.n168 VDD1.n167 9.3005
R895 VDD1.n170 VDD1.n169 9.3005
R896 VDD1.n117 VDD1.n116 9.3005
R897 VDD1.n176 VDD1.n175 9.3005
R898 VDD1.n178 VDD1.n177 9.3005
R899 VDD1.n179 VDD1.n112 9.3005
R900 VDD1.n97 VDD1.n2 8.92171
R901 VDD1.n65 VDD1.n64 8.92171
R902 VDD1.n49 VDD1.n25 8.92171
R903 VDD1.n151 VDD1.n127 8.92171
R904 VDD1.n167 VDD1.n166 8.92171
R905 VDD1.n200 VDD1.n105 8.92171
R906 VDD1.n98 VDD1.n0 8.14595
R907 VDD1.n61 VDD1.n19 8.14595
R908 VDD1.n53 VDD1.n52 8.14595
R909 VDD1.n155 VDD1.n154 8.14595
R910 VDD1.n163 VDD1.n121 8.14595
R911 VDD1.n201 VDD1.n103 8.14595
R912 VDD1.n60 VDD1.n21 7.3702
R913 VDD1.n56 VDD1.n23 7.3702
R914 VDD1.n158 VDD1.n125 7.3702
R915 VDD1.n162 VDD1.n123 7.3702
R916 VDD1.n57 VDD1.n21 6.59444
R917 VDD1.n57 VDD1.n56 6.59444
R918 VDD1.n159 VDD1.n158 6.59444
R919 VDD1.n159 VDD1.n123 6.59444
R920 VDD1.n100 VDD1.n0 5.81868
R921 VDD1.n61 VDD1.n60 5.81868
R922 VDD1.n53 VDD1.n23 5.81868
R923 VDD1.n155 VDD1.n125 5.81868
R924 VDD1.n163 VDD1.n162 5.81868
R925 VDD1.n203 VDD1.n103 5.81868
R926 VDD1.n98 VDD1.n97 5.04292
R927 VDD1.n64 VDD1.n19 5.04292
R928 VDD1.n52 VDD1.n25 5.04292
R929 VDD1.n154 VDD1.n127 5.04292
R930 VDD1.n166 VDD1.n121 5.04292
R931 VDD1.n201 VDD1.n200 5.04292
R932 VDD1.n94 VDD1.n2 4.26717
R933 VDD1.n65 VDD1.n17 4.26717
R934 VDD1.n49 VDD1.n48 4.26717
R935 VDD1.n151 VDD1.n150 4.26717
R936 VDD1.n167 VDD1.n119 4.26717
R937 VDD1.n197 VDD1.n105 4.26717
R938 VDD1.n35 VDD1.n34 3.70982
R939 VDD1.n137 VDD1.n136 3.70982
R940 VDD1.n93 VDD1.n4 3.49141
R941 VDD1.n69 VDD1.n68 3.49141
R942 VDD1.n45 VDD1.n27 3.49141
R943 VDD1.n147 VDD1.n129 3.49141
R944 VDD1.n171 VDD1.n170 3.49141
R945 VDD1.n196 VDD1.n107 3.49141
R946 VDD1.n90 VDD1.n89 2.71565
R947 VDD1.n72 VDD1.n15 2.71565
R948 VDD1.n44 VDD1.n29 2.71565
R949 VDD1.n146 VDD1.n131 2.71565
R950 VDD1.n174 VDD1.n117 2.71565
R951 VDD1.n193 VDD1.n192 2.71565
R952 VDD1.n86 VDD1.n6 1.93989
R953 VDD1.n73 VDD1.n13 1.93989
R954 VDD1.n41 VDD1.n40 1.93989
R955 VDD1.n143 VDD1.n142 1.93989
R956 VDD1.n175 VDD1.n115 1.93989
R957 VDD1.n189 VDD1.n109 1.93989
R958 VDD1.n208 VDD1.t4 1.77673
R959 VDD1.n208 VDD1.t8 1.77673
R960 VDD1.n101 VDD1.t6 1.77673
R961 VDD1.n101 VDD1.t7 1.77673
R962 VDD1.n206 VDD1.t2 1.77673
R963 VDD1.n206 VDD1.t0 1.77673
R964 VDD1.n204 VDD1.t3 1.77673
R965 VDD1.n204 VDD1.t1 1.77673
R966 VDD1.n85 VDD1.n8 1.16414
R967 VDD1.n77 VDD1.n76 1.16414
R968 VDD1.n37 VDD1.n31 1.16414
R969 VDD1.n139 VDD1.n133 1.16414
R970 VDD1.n180 VDD1.n178 1.16414
R971 VDD1.n188 VDD1.n111 1.16414
R972 VDD1 VDD1.n209 0.627655
R973 VDD1.n82 VDD1.n81 0.388379
R974 VDD1.n12 VDD1.n10 0.388379
R975 VDD1.n36 VDD1.n33 0.388379
R976 VDD1.n138 VDD1.n135 0.388379
R977 VDD1.n179 VDD1.n113 0.388379
R978 VDD1.n185 VDD1.n184 0.388379
R979 VDD1 VDD1.n102 0.287138
R980 VDD1.n207 VDD1.n205 0.173602
R981 VDD1.n99 VDD1.n1 0.155672
R982 VDD1.n92 VDD1.n1 0.155672
R983 VDD1.n92 VDD1.n91 0.155672
R984 VDD1.n91 VDD1.n5 0.155672
R985 VDD1.n84 VDD1.n5 0.155672
R986 VDD1.n84 VDD1.n83 0.155672
R987 VDD1.n83 VDD1.n9 0.155672
R988 VDD1.n75 VDD1.n9 0.155672
R989 VDD1.n75 VDD1.n74 0.155672
R990 VDD1.n74 VDD1.n14 0.155672
R991 VDD1.n67 VDD1.n14 0.155672
R992 VDD1.n67 VDD1.n66 0.155672
R993 VDD1.n66 VDD1.n18 0.155672
R994 VDD1.n59 VDD1.n18 0.155672
R995 VDD1.n59 VDD1.n58 0.155672
R996 VDD1.n58 VDD1.n22 0.155672
R997 VDD1.n51 VDD1.n22 0.155672
R998 VDD1.n51 VDD1.n50 0.155672
R999 VDD1.n50 VDD1.n26 0.155672
R1000 VDD1.n43 VDD1.n26 0.155672
R1001 VDD1.n43 VDD1.n42 0.155672
R1002 VDD1.n42 VDD1.n30 0.155672
R1003 VDD1.n35 VDD1.n30 0.155672
R1004 VDD1.n137 VDD1.n132 0.155672
R1005 VDD1.n144 VDD1.n132 0.155672
R1006 VDD1.n145 VDD1.n144 0.155672
R1007 VDD1.n145 VDD1.n128 0.155672
R1008 VDD1.n152 VDD1.n128 0.155672
R1009 VDD1.n153 VDD1.n152 0.155672
R1010 VDD1.n153 VDD1.n124 0.155672
R1011 VDD1.n160 VDD1.n124 0.155672
R1012 VDD1.n161 VDD1.n160 0.155672
R1013 VDD1.n161 VDD1.n120 0.155672
R1014 VDD1.n168 VDD1.n120 0.155672
R1015 VDD1.n169 VDD1.n168 0.155672
R1016 VDD1.n169 VDD1.n116 0.155672
R1017 VDD1.n176 VDD1.n116 0.155672
R1018 VDD1.n177 VDD1.n176 0.155672
R1019 VDD1.n177 VDD1.n112 0.155672
R1020 VDD1.n186 VDD1.n112 0.155672
R1021 VDD1.n187 VDD1.n186 0.155672
R1022 VDD1.n187 VDD1.n108 0.155672
R1023 VDD1.n194 VDD1.n108 0.155672
R1024 VDD1.n195 VDD1.n194 0.155672
R1025 VDD1.n195 VDD1.n104 0.155672
R1026 VDD1.n202 VDD1.n104 0.155672
R1027 B.n143 B.t3 806.763
R1028 B.n151 B.t0 806.763
R1029 B.n46 B.t9 806.763
R1030 B.n54 B.t6 806.763
R1031 B.n514 B.n85 585
R1032 B.n516 B.n515 585
R1033 B.n517 B.n84 585
R1034 B.n519 B.n518 585
R1035 B.n520 B.n83 585
R1036 B.n522 B.n521 585
R1037 B.n523 B.n82 585
R1038 B.n525 B.n524 585
R1039 B.n526 B.n81 585
R1040 B.n528 B.n527 585
R1041 B.n529 B.n80 585
R1042 B.n531 B.n530 585
R1043 B.n532 B.n79 585
R1044 B.n534 B.n533 585
R1045 B.n535 B.n78 585
R1046 B.n537 B.n536 585
R1047 B.n538 B.n77 585
R1048 B.n540 B.n539 585
R1049 B.n541 B.n76 585
R1050 B.n543 B.n542 585
R1051 B.n544 B.n75 585
R1052 B.n546 B.n545 585
R1053 B.n547 B.n74 585
R1054 B.n549 B.n548 585
R1055 B.n550 B.n73 585
R1056 B.n552 B.n551 585
R1057 B.n553 B.n72 585
R1058 B.n555 B.n554 585
R1059 B.n556 B.n71 585
R1060 B.n558 B.n557 585
R1061 B.n559 B.n70 585
R1062 B.n561 B.n560 585
R1063 B.n562 B.n69 585
R1064 B.n564 B.n563 585
R1065 B.n565 B.n68 585
R1066 B.n567 B.n566 585
R1067 B.n568 B.n67 585
R1068 B.n570 B.n569 585
R1069 B.n571 B.n66 585
R1070 B.n573 B.n572 585
R1071 B.n574 B.n65 585
R1072 B.n576 B.n575 585
R1073 B.n577 B.n64 585
R1074 B.n579 B.n578 585
R1075 B.n580 B.n63 585
R1076 B.n582 B.n581 585
R1077 B.n583 B.n62 585
R1078 B.n585 B.n584 585
R1079 B.n586 B.n61 585
R1080 B.n588 B.n587 585
R1081 B.n589 B.n60 585
R1082 B.n591 B.n590 585
R1083 B.n592 B.n59 585
R1084 B.n594 B.n593 585
R1085 B.n595 B.n58 585
R1086 B.n597 B.n596 585
R1087 B.n598 B.n57 585
R1088 B.n600 B.n599 585
R1089 B.n601 B.n53 585
R1090 B.n603 B.n602 585
R1091 B.n604 B.n52 585
R1092 B.n606 B.n605 585
R1093 B.n607 B.n51 585
R1094 B.n609 B.n608 585
R1095 B.n610 B.n50 585
R1096 B.n612 B.n611 585
R1097 B.n613 B.n49 585
R1098 B.n615 B.n614 585
R1099 B.n616 B.n48 585
R1100 B.n618 B.n617 585
R1101 B.n620 B.n45 585
R1102 B.n622 B.n621 585
R1103 B.n623 B.n44 585
R1104 B.n625 B.n624 585
R1105 B.n626 B.n43 585
R1106 B.n628 B.n627 585
R1107 B.n629 B.n42 585
R1108 B.n631 B.n630 585
R1109 B.n632 B.n41 585
R1110 B.n634 B.n633 585
R1111 B.n635 B.n40 585
R1112 B.n637 B.n636 585
R1113 B.n638 B.n39 585
R1114 B.n640 B.n639 585
R1115 B.n641 B.n38 585
R1116 B.n643 B.n642 585
R1117 B.n644 B.n37 585
R1118 B.n646 B.n645 585
R1119 B.n647 B.n36 585
R1120 B.n649 B.n648 585
R1121 B.n650 B.n35 585
R1122 B.n652 B.n651 585
R1123 B.n653 B.n34 585
R1124 B.n655 B.n654 585
R1125 B.n656 B.n33 585
R1126 B.n658 B.n657 585
R1127 B.n659 B.n32 585
R1128 B.n661 B.n660 585
R1129 B.n662 B.n31 585
R1130 B.n664 B.n663 585
R1131 B.n665 B.n30 585
R1132 B.n667 B.n666 585
R1133 B.n668 B.n29 585
R1134 B.n670 B.n669 585
R1135 B.n671 B.n28 585
R1136 B.n673 B.n672 585
R1137 B.n674 B.n27 585
R1138 B.n676 B.n675 585
R1139 B.n677 B.n26 585
R1140 B.n679 B.n678 585
R1141 B.n680 B.n25 585
R1142 B.n682 B.n681 585
R1143 B.n683 B.n24 585
R1144 B.n685 B.n684 585
R1145 B.n686 B.n23 585
R1146 B.n688 B.n687 585
R1147 B.n689 B.n22 585
R1148 B.n691 B.n690 585
R1149 B.n692 B.n21 585
R1150 B.n694 B.n693 585
R1151 B.n695 B.n20 585
R1152 B.n697 B.n696 585
R1153 B.n698 B.n19 585
R1154 B.n700 B.n699 585
R1155 B.n701 B.n18 585
R1156 B.n703 B.n702 585
R1157 B.n704 B.n17 585
R1158 B.n706 B.n705 585
R1159 B.n707 B.n16 585
R1160 B.n709 B.n708 585
R1161 B.n513 B.n512 585
R1162 B.n511 B.n86 585
R1163 B.n510 B.n509 585
R1164 B.n508 B.n87 585
R1165 B.n507 B.n506 585
R1166 B.n505 B.n88 585
R1167 B.n504 B.n503 585
R1168 B.n502 B.n89 585
R1169 B.n501 B.n500 585
R1170 B.n499 B.n90 585
R1171 B.n498 B.n497 585
R1172 B.n496 B.n91 585
R1173 B.n495 B.n494 585
R1174 B.n493 B.n92 585
R1175 B.n492 B.n491 585
R1176 B.n490 B.n93 585
R1177 B.n489 B.n488 585
R1178 B.n487 B.n94 585
R1179 B.n486 B.n485 585
R1180 B.n484 B.n95 585
R1181 B.n483 B.n482 585
R1182 B.n481 B.n96 585
R1183 B.n480 B.n479 585
R1184 B.n478 B.n97 585
R1185 B.n477 B.n476 585
R1186 B.n475 B.n98 585
R1187 B.n474 B.n473 585
R1188 B.n472 B.n99 585
R1189 B.n471 B.n470 585
R1190 B.n469 B.n100 585
R1191 B.n468 B.n467 585
R1192 B.n466 B.n101 585
R1193 B.n465 B.n464 585
R1194 B.n463 B.n102 585
R1195 B.n462 B.n461 585
R1196 B.n460 B.n103 585
R1197 B.n459 B.n458 585
R1198 B.n457 B.n104 585
R1199 B.n456 B.n455 585
R1200 B.n454 B.n105 585
R1201 B.n453 B.n452 585
R1202 B.n451 B.n106 585
R1203 B.n450 B.n449 585
R1204 B.n448 B.n107 585
R1205 B.n447 B.n446 585
R1206 B.n445 B.n108 585
R1207 B.n444 B.n443 585
R1208 B.n442 B.n109 585
R1209 B.n441 B.n440 585
R1210 B.n439 B.n110 585
R1211 B.n438 B.n437 585
R1212 B.n436 B.n111 585
R1213 B.n435 B.n434 585
R1214 B.n433 B.n112 585
R1215 B.n432 B.n431 585
R1216 B.n235 B.n182 585
R1217 B.n237 B.n236 585
R1218 B.n238 B.n181 585
R1219 B.n240 B.n239 585
R1220 B.n241 B.n180 585
R1221 B.n243 B.n242 585
R1222 B.n244 B.n179 585
R1223 B.n246 B.n245 585
R1224 B.n247 B.n178 585
R1225 B.n249 B.n248 585
R1226 B.n250 B.n177 585
R1227 B.n252 B.n251 585
R1228 B.n253 B.n176 585
R1229 B.n255 B.n254 585
R1230 B.n256 B.n175 585
R1231 B.n258 B.n257 585
R1232 B.n259 B.n174 585
R1233 B.n261 B.n260 585
R1234 B.n262 B.n173 585
R1235 B.n264 B.n263 585
R1236 B.n265 B.n172 585
R1237 B.n267 B.n266 585
R1238 B.n268 B.n171 585
R1239 B.n270 B.n269 585
R1240 B.n271 B.n170 585
R1241 B.n273 B.n272 585
R1242 B.n274 B.n169 585
R1243 B.n276 B.n275 585
R1244 B.n277 B.n168 585
R1245 B.n279 B.n278 585
R1246 B.n280 B.n167 585
R1247 B.n282 B.n281 585
R1248 B.n283 B.n166 585
R1249 B.n285 B.n284 585
R1250 B.n286 B.n165 585
R1251 B.n288 B.n287 585
R1252 B.n289 B.n164 585
R1253 B.n291 B.n290 585
R1254 B.n292 B.n163 585
R1255 B.n294 B.n293 585
R1256 B.n295 B.n162 585
R1257 B.n297 B.n296 585
R1258 B.n298 B.n161 585
R1259 B.n300 B.n299 585
R1260 B.n301 B.n160 585
R1261 B.n303 B.n302 585
R1262 B.n304 B.n159 585
R1263 B.n306 B.n305 585
R1264 B.n307 B.n158 585
R1265 B.n309 B.n308 585
R1266 B.n310 B.n157 585
R1267 B.n312 B.n311 585
R1268 B.n313 B.n156 585
R1269 B.n315 B.n314 585
R1270 B.n316 B.n155 585
R1271 B.n318 B.n317 585
R1272 B.n319 B.n154 585
R1273 B.n321 B.n320 585
R1274 B.n322 B.n153 585
R1275 B.n324 B.n323 585
R1276 B.n326 B.n150 585
R1277 B.n328 B.n327 585
R1278 B.n329 B.n149 585
R1279 B.n331 B.n330 585
R1280 B.n332 B.n148 585
R1281 B.n334 B.n333 585
R1282 B.n335 B.n147 585
R1283 B.n337 B.n336 585
R1284 B.n338 B.n146 585
R1285 B.n340 B.n339 585
R1286 B.n342 B.n341 585
R1287 B.n343 B.n142 585
R1288 B.n345 B.n344 585
R1289 B.n346 B.n141 585
R1290 B.n348 B.n347 585
R1291 B.n349 B.n140 585
R1292 B.n351 B.n350 585
R1293 B.n352 B.n139 585
R1294 B.n354 B.n353 585
R1295 B.n355 B.n138 585
R1296 B.n357 B.n356 585
R1297 B.n358 B.n137 585
R1298 B.n360 B.n359 585
R1299 B.n361 B.n136 585
R1300 B.n363 B.n362 585
R1301 B.n364 B.n135 585
R1302 B.n366 B.n365 585
R1303 B.n367 B.n134 585
R1304 B.n369 B.n368 585
R1305 B.n370 B.n133 585
R1306 B.n372 B.n371 585
R1307 B.n373 B.n132 585
R1308 B.n375 B.n374 585
R1309 B.n376 B.n131 585
R1310 B.n378 B.n377 585
R1311 B.n379 B.n130 585
R1312 B.n381 B.n380 585
R1313 B.n382 B.n129 585
R1314 B.n384 B.n383 585
R1315 B.n385 B.n128 585
R1316 B.n387 B.n386 585
R1317 B.n388 B.n127 585
R1318 B.n390 B.n389 585
R1319 B.n391 B.n126 585
R1320 B.n393 B.n392 585
R1321 B.n394 B.n125 585
R1322 B.n396 B.n395 585
R1323 B.n397 B.n124 585
R1324 B.n399 B.n398 585
R1325 B.n400 B.n123 585
R1326 B.n402 B.n401 585
R1327 B.n403 B.n122 585
R1328 B.n405 B.n404 585
R1329 B.n406 B.n121 585
R1330 B.n408 B.n407 585
R1331 B.n409 B.n120 585
R1332 B.n411 B.n410 585
R1333 B.n412 B.n119 585
R1334 B.n414 B.n413 585
R1335 B.n415 B.n118 585
R1336 B.n417 B.n416 585
R1337 B.n418 B.n117 585
R1338 B.n420 B.n419 585
R1339 B.n421 B.n116 585
R1340 B.n423 B.n422 585
R1341 B.n424 B.n115 585
R1342 B.n426 B.n425 585
R1343 B.n427 B.n114 585
R1344 B.n429 B.n428 585
R1345 B.n430 B.n113 585
R1346 B.n234 B.n233 585
R1347 B.n232 B.n183 585
R1348 B.n231 B.n230 585
R1349 B.n229 B.n184 585
R1350 B.n228 B.n227 585
R1351 B.n226 B.n185 585
R1352 B.n225 B.n224 585
R1353 B.n223 B.n186 585
R1354 B.n222 B.n221 585
R1355 B.n220 B.n187 585
R1356 B.n219 B.n218 585
R1357 B.n217 B.n188 585
R1358 B.n216 B.n215 585
R1359 B.n214 B.n189 585
R1360 B.n213 B.n212 585
R1361 B.n211 B.n190 585
R1362 B.n210 B.n209 585
R1363 B.n208 B.n191 585
R1364 B.n207 B.n206 585
R1365 B.n205 B.n192 585
R1366 B.n204 B.n203 585
R1367 B.n202 B.n193 585
R1368 B.n201 B.n200 585
R1369 B.n199 B.n194 585
R1370 B.n198 B.n197 585
R1371 B.n196 B.n195 585
R1372 B.n2 B.n0 585
R1373 B.n749 B.n1 585
R1374 B.n748 B.n747 585
R1375 B.n746 B.n3 585
R1376 B.n745 B.n744 585
R1377 B.n743 B.n4 585
R1378 B.n742 B.n741 585
R1379 B.n740 B.n5 585
R1380 B.n739 B.n738 585
R1381 B.n737 B.n6 585
R1382 B.n736 B.n735 585
R1383 B.n734 B.n7 585
R1384 B.n733 B.n732 585
R1385 B.n731 B.n8 585
R1386 B.n730 B.n729 585
R1387 B.n728 B.n9 585
R1388 B.n727 B.n726 585
R1389 B.n725 B.n10 585
R1390 B.n724 B.n723 585
R1391 B.n722 B.n11 585
R1392 B.n721 B.n720 585
R1393 B.n719 B.n12 585
R1394 B.n718 B.n717 585
R1395 B.n716 B.n13 585
R1396 B.n715 B.n714 585
R1397 B.n713 B.n14 585
R1398 B.n712 B.n711 585
R1399 B.n710 B.n15 585
R1400 B.n751 B.n750 585
R1401 B.n143 B.t5 509.81
R1402 B.n54 B.t7 509.81
R1403 B.n151 B.t2 509.81
R1404 B.n46 B.t10 509.81
R1405 B.n144 B.t4 489.252
R1406 B.n55 B.t8 489.252
R1407 B.n152 B.t1 489.252
R1408 B.n47 B.t11 489.252
R1409 B.n233 B.n182 458.866
R1410 B.n708 B.n15 458.866
R1411 B.n431 B.n430 458.866
R1412 B.n514 B.n513 458.866
R1413 B.n233 B.n232 163.367
R1414 B.n232 B.n231 163.367
R1415 B.n231 B.n184 163.367
R1416 B.n227 B.n184 163.367
R1417 B.n227 B.n226 163.367
R1418 B.n226 B.n225 163.367
R1419 B.n225 B.n186 163.367
R1420 B.n221 B.n186 163.367
R1421 B.n221 B.n220 163.367
R1422 B.n220 B.n219 163.367
R1423 B.n219 B.n188 163.367
R1424 B.n215 B.n188 163.367
R1425 B.n215 B.n214 163.367
R1426 B.n214 B.n213 163.367
R1427 B.n213 B.n190 163.367
R1428 B.n209 B.n190 163.367
R1429 B.n209 B.n208 163.367
R1430 B.n208 B.n207 163.367
R1431 B.n207 B.n192 163.367
R1432 B.n203 B.n192 163.367
R1433 B.n203 B.n202 163.367
R1434 B.n202 B.n201 163.367
R1435 B.n201 B.n194 163.367
R1436 B.n197 B.n194 163.367
R1437 B.n197 B.n196 163.367
R1438 B.n196 B.n2 163.367
R1439 B.n750 B.n2 163.367
R1440 B.n750 B.n749 163.367
R1441 B.n749 B.n748 163.367
R1442 B.n748 B.n3 163.367
R1443 B.n744 B.n3 163.367
R1444 B.n744 B.n743 163.367
R1445 B.n743 B.n742 163.367
R1446 B.n742 B.n5 163.367
R1447 B.n738 B.n5 163.367
R1448 B.n738 B.n737 163.367
R1449 B.n737 B.n736 163.367
R1450 B.n736 B.n7 163.367
R1451 B.n732 B.n7 163.367
R1452 B.n732 B.n731 163.367
R1453 B.n731 B.n730 163.367
R1454 B.n730 B.n9 163.367
R1455 B.n726 B.n9 163.367
R1456 B.n726 B.n725 163.367
R1457 B.n725 B.n724 163.367
R1458 B.n724 B.n11 163.367
R1459 B.n720 B.n11 163.367
R1460 B.n720 B.n719 163.367
R1461 B.n719 B.n718 163.367
R1462 B.n718 B.n13 163.367
R1463 B.n714 B.n13 163.367
R1464 B.n714 B.n713 163.367
R1465 B.n713 B.n712 163.367
R1466 B.n712 B.n15 163.367
R1467 B.n237 B.n182 163.367
R1468 B.n238 B.n237 163.367
R1469 B.n239 B.n238 163.367
R1470 B.n239 B.n180 163.367
R1471 B.n243 B.n180 163.367
R1472 B.n244 B.n243 163.367
R1473 B.n245 B.n244 163.367
R1474 B.n245 B.n178 163.367
R1475 B.n249 B.n178 163.367
R1476 B.n250 B.n249 163.367
R1477 B.n251 B.n250 163.367
R1478 B.n251 B.n176 163.367
R1479 B.n255 B.n176 163.367
R1480 B.n256 B.n255 163.367
R1481 B.n257 B.n256 163.367
R1482 B.n257 B.n174 163.367
R1483 B.n261 B.n174 163.367
R1484 B.n262 B.n261 163.367
R1485 B.n263 B.n262 163.367
R1486 B.n263 B.n172 163.367
R1487 B.n267 B.n172 163.367
R1488 B.n268 B.n267 163.367
R1489 B.n269 B.n268 163.367
R1490 B.n269 B.n170 163.367
R1491 B.n273 B.n170 163.367
R1492 B.n274 B.n273 163.367
R1493 B.n275 B.n274 163.367
R1494 B.n275 B.n168 163.367
R1495 B.n279 B.n168 163.367
R1496 B.n280 B.n279 163.367
R1497 B.n281 B.n280 163.367
R1498 B.n281 B.n166 163.367
R1499 B.n285 B.n166 163.367
R1500 B.n286 B.n285 163.367
R1501 B.n287 B.n286 163.367
R1502 B.n287 B.n164 163.367
R1503 B.n291 B.n164 163.367
R1504 B.n292 B.n291 163.367
R1505 B.n293 B.n292 163.367
R1506 B.n293 B.n162 163.367
R1507 B.n297 B.n162 163.367
R1508 B.n298 B.n297 163.367
R1509 B.n299 B.n298 163.367
R1510 B.n299 B.n160 163.367
R1511 B.n303 B.n160 163.367
R1512 B.n304 B.n303 163.367
R1513 B.n305 B.n304 163.367
R1514 B.n305 B.n158 163.367
R1515 B.n309 B.n158 163.367
R1516 B.n310 B.n309 163.367
R1517 B.n311 B.n310 163.367
R1518 B.n311 B.n156 163.367
R1519 B.n315 B.n156 163.367
R1520 B.n316 B.n315 163.367
R1521 B.n317 B.n316 163.367
R1522 B.n317 B.n154 163.367
R1523 B.n321 B.n154 163.367
R1524 B.n322 B.n321 163.367
R1525 B.n323 B.n322 163.367
R1526 B.n323 B.n150 163.367
R1527 B.n328 B.n150 163.367
R1528 B.n329 B.n328 163.367
R1529 B.n330 B.n329 163.367
R1530 B.n330 B.n148 163.367
R1531 B.n334 B.n148 163.367
R1532 B.n335 B.n334 163.367
R1533 B.n336 B.n335 163.367
R1534 B.n336 B.n146 163.367
R1535 B.n340 B.n146 163.367
R1536 B.n341 B.n340 163.367
R1537 B.n341 B.n142 163.367
R1538 B.n345 B.n142 163.367
R1539 B.n346 B.n345 163.367
R1540 B.n347 B.n346 163.367
R1541 B.n347 B.n140 163.367
R1542 B.n351 B.n140 163.367
R1543 B.n352 B.n351 163.367
R1544 B.n353 B.n352 163.367
R1545 B.n353 B.n138 163.367
R1546 B.n357 B.n138 163.367
R1547 B.n358 B.n357 163.367
R1548 B.n359 B.n358 163.367
R1549 B.n359 B.n136 163.367
R1550 B.n363 B.n136 163.367
R1551 B.n364 B.n363 163.367
R1552 B.n365 B.n364 163.367
R1553 B.n365 B.n134 163.367
R1554 B.n369 B.n134 163.367
R1555 B.n370 B.n369 163.367
R1556 B.n371 B.n370 163.367
R1557 B.n371 B.n132 163.367
R1558 B.n375 B.n132 163.367
R1559 B.n376 B.n375 163.367
R1560 B.n377 B.n376 163.367
R1561 B.n377 B.n130 163.367
R1562 B.n381 B.n130 163.367
R1563 B.n382 B.n381 163.367
R1564 B.n383 B.n382 163.367
R1565 B.n383 B.n128 163.367
R1566 B.n387 B.n128 163.367
R1567 B.n388 B.n387 163.367
R1568 B.n389 B.n388 163.367
R1569 B.n389 B.n126 163.367
R1570 B.n393 B.n126 163.367
R1571 B.n394 B.n393 163.367
R1572 B.n395 B.n394 163.367
R1573 B.n395 B.n124 163.367
R1574 B.n399 B.n124 163.367
R1575 B.n400 B.n399 163.367
R1576 B.n401 B.n400 163.367
R1577 B.n401 B.n122 163.367
R1578 B.n405 B.n122 163.367
R1579 B.n406 B.n405 163.367
R1580 B.n407 B.n406 163.367
R1581 B.n407 B.n120 163.367
R1582 B.n411 B.n120 163.367
R1583 B.n412 B.n411 163.367
R1584 B.n413 B.n412 163.367
R1585 B.n413 B.n118 163.367
R1586 B.n417 B.n118 163.367
R1587 B.n418 B.n417 163.367
R1588 B.n419 B.n418 163.367
R1589 B.n419 B.n116 163.367
R1590 B.n423 B.n116 163.367
R1591 B.n424 B.n423 163.367
R1592 B.n425 B.n424 163.367
R1593 B.n425 B.n114 163.367
R1594 B.n429 B.n114 163.367
R1595 B.n430 B.n429 163.367
R1596 B.n431 B.n112 163.367
R1597 B.n435 B.n112 163.367
R1598 B.n436 B.n435 163.367
R1599 B.n437 B.n436 163.367
R1600 B.n437 B.n110 163.367
R1601 B.n441 B.n110 163.367
R1602 B.n442 B.n441 163.367
R1603 B.n443 B.n442 163.367
R1604 B.n443 B.n108 163.367
R1605 B.n447 B.n108 163.367
R1606 B.n448 B.n447 163.367
R1607 B.n449 B.n448 163.367
R1608 B.n449 B.n106 163.367
R1609 B.n453 B.n106 163.367
R1610 B.n454 B.n453 163.367
R1611 B.n455 B.n454 163.367
R1612 B.n455 B.n104 163.367
R1613 B.n459 B.n104 163.367
R1614 B.n460 B.n459 163.367
R1615 B.n461 B.n460 163.367
R1616 B.n461 B.n102 163.367
R1617 B.n465 B.n102 163.367
R1618 B.n466 B.n465 163.367
R1619 B.n467 B.n466 163.367
R1620 B.n467 B.n100 163.367
R1621 B.n471 B.n100 163.367
R1622 B.n472 B.n471 163.367
R1623 B.n473 B.n472 163.367
R1624 B.n473 B.n98 163.367
R1625 B.n477 B.n98 163.367
R1626 B.n478 B.n477 163.367
R1627 B.n479 B.n478 163.367
R1628 B.n479 B.n96 163.367
R1629 B.n483 B.n96 163.367
R1630 B.n484 B.n483 163.367
R1631 B.n485 B.n484 163.367
R1632 B.n485 B.n94 163.367
R1633 B.n489 B.n94 163.367
R1634 B.n490 B.n489 163.367
R1635 B.n491 B.n490 163.367
R1636 B.n491 B.n92 163.367
R1637 B.n495 B.n92 163.367
R1638 B.n496 B.n495 163.367
R1639 B.n497 B.n496 163.367
R1640 B.n497 B.n90 163.367
R1641 B.n501 B.n90 163.367
R1642 B.n502 B.n501 163.367
R1643 B.n503 B.n502 163.367
R1644 B.n503 B.n88 163.367
R1645 B.n507 B.n88 163.367
R1646 B.n508 B.n507 163.367
R1647 B.n509 B.n508 163.367
R1648 B.n509 B.n86 163.367
R1649 B.n513 B.n86 163.367
R1650 B.n708 B.n707 163.367
R1651 B.n707 B.n706 163.367
R1652 B.n706 B.n17 163.367
R1653 B.n702 B.n17 163.367
R1654 B.n702 B.n701 163.367
R1655 B.n701 B.n700 163.367
R1656 B.n700 B.n19 163.367
R1657 B.n696 B.n19 163.367
R1658 B.n696 B.n695 163.367
R1659 B.n695 B.n694 163.367
R1660 B.n694 B.n21 163.367
R1661 B.n690 B.n21 163.367
R1662 B.n690 B.n689 163.367
R1663 B.n689 B.n688 163.367
R1664 B.n688 B.n23 163.367
R1665 B.n684 B.n23 163.367
R1666 B.n684 B.n683 163.367
R1667 B.n683 B.n682 163.367
R1668 B.n682 B.n25 163.367
R1669 B.n678 B.n25 163.367
R1670 B.n678 B.n677 163.367
R1671 B.n677 B.n676 163.367
R1672 B.n676 B.n27 163.367
R1673 B.n672 B.n27 163.367
R1674 B.n672 B.n671 163.367
R1675 B.n671 B.n670 163.367
R1676 B.n670 B.n29 163.367
R1677 B.n666 B.n29 163.367
R1678 B.n666 B.n665 163.367
R1679 B.n665 B.n664 163.367
R1680 B.n664 B.n31 163.367
R1681 B.n660 B.n31 163.367
R1682 B.n660 B.n659 163.367
R1683 B.n659 B.n658 163.367
R1684 B.n658 B.n33 163.367
R1685 B.n654 B.n33 163.367
R1686 B.n654 B.n653 163.367
R1687 B.n653 B.n652 163.367
R1688 B.n652 B.n35 163.367
R1689 B.n648 B.n35 163.367
R1690 B.n648 B.n647 163.367
R1691 B.n647 B.n646 163.367
R1692 B.n646 B.n37 163.367
R1693 B.n642 B.n37 163.367
R1694 B.n642 B.n641 163.367
R1695 B.n641 B.n640 163.367
R1696 B.n640 B.n39 163.367
R1697 B.n636 B.n39 163.367
R1698 B.n636 B.n635 163.367
R1699 B.n635 B.n634 163.367
R1700 B.n634 B.n41 163.367
R1701 B.n630 B.n41 163.367
R1702 B.n630 B.n629 163.367
R1703 B.n629 B.n628 163.367
R1704 B.n628 B.n43 163.367
R1705 B.n624 B.n43 163.367
R1706 B.n624 B.n623 163.367
R1707 B.n623 B.n622 163.367
R1708 B.n622 B.n45 163.367
R1709 B.n617 B.n45 163.367
R1710 B.n617 B.n616 163.367
R1711 B.n616 B.n615 163.367
R1712 B.n615 B.n49 163.367
R1713 B.n611 B.n49 163.367
R1714 B.n611 B.n610 163.367
R1715 B.n610 B.n609 163.367
R1716 B.n609 B.n51 163.367
R1717 B.n605 B.n51 163.367
R1718 B.n605 B.n604 163.367
R1719 B.n604 B.n603 163.367
R1720 B.n603 B.n53 163.367
R1721 B.n599 B.n53 163.367
R1722 B.n599 B.n598 163.367
R1723 B.n598 B.n597 163.367
R1724 B.n597 B.n58 163.367
R1725 B.n593 B.n58 163.367
R1726 B.n593 B.n592 163.367
R1727 B.n592 B.n591 163.367
R1728 B.n591 B.n60 163.367
R1729 B.n587 B.n60 163.367
R1730 B.n587 B.n586 163.367
R1731 B.n586 B.n585 163.367
R1732 B.n585 B.n62 163.367
R1733 B.n581 B.n62 163.367
R1734 B.n581 B.n580 163.367
R1735 B.n580 B.n579 163.367
R1736 B.n579 B.n64 163.367
R1737 B.n575 B.n64 163.367
R1738 B.n575 B.n574 163.367
R1739 B.n574 B.n573 163.367
R1740 B.n573 B.n66 163.367
R1741 B.n569 B.n66 163.367
R1742 B.n569 B.n568 163.367
R1743 B.n568 B.n567 163.367
R1744 B.n567 B.n68 163.367
R1745 B.n563 B.n68 163.367
R1746 B.n563 B.n562 163.367
R1747 B.n562 B.n561 163.367
R1748 B.n561 B.n70 163.367
R1749 B.n557 B.n70 163.367
R1750 B.n557 B.n556 163.367
R1751 B.n556 B.n555 163.367
R1752 B.n555 B.n72 163.367
R1753 B.n551 B.n72 163.367
R1754 B.n551 B.n550 163.367
R1755 B.n550 B.n549 163.367
R1756 B.n549 B.n74 163.367
R1757 B.n545 B.n74 163.367
R1758 B.n545 B.n544 163.367
R1759 B.n544 B.n543 163.367
R1760 B.n543 B.n76 163.367
R1761 B.n539 B.n76 163.367
R1762 B.n539 B.n538 163.367
R1763 B.n538 B.n537 163.367
R1764 B.n537 B.n78 163.367
R1765 B.n533 B.n78 163.367
R1766 B.n533 B.n532 163.367
R1767 B.n532 B.n531 163.367
R1768 B.n531 B.n80 163.367
R1769 B.n527 B.n80 163.367
R1770 B.n527 B.n526 163.367
R1771 B.n526 B.n525 163.367
R1772 B.n525 B.n82 163.367
R1773 B.n521 B.n82 163.367
R1774 B.n521 B.n520 163.367
R1775 B.n520 B.n519 163.367
R1776 B.n519 B.n84 163.367
R1777 B.n515 B.n84 163.367
R1778 B.n515 B.n514 163.367
R1779 B.n145 B.n144 59.5399
R1780 B.n325 B.n152 59.5399
R1781 B.n619 B.n47 59.5399
R1782 B.n56 B.n55 59.5399
R1783 B.n710 B.n709 29.8151
R1784 B.n432 B.n113 29.8151
R1785 B.n235 B.n234 29.8151
R1786 B.n512 B.n85 29.8151
R1787 B.n144 B.n143 20.5581
R1788 B.n152 B.n151 20.5581
R1789 B.n47 B.n46 20.5581
R1790 B.n55 B.n54 20.5581
R1791 B B.n751 18.0485
R1792 B.n709 B.n16 10.6151
R1793 B.n705 B.n16 10.6151
R1794 B.n705 B.n704 10.6151
R1795 B.n704 B.n703 10.6151
R1796 B.n703 B.n18 10.6151
R1797 B.n699 B.n18 10.6151
R1798 B.n699 B.n698 10.6151
R1799 B.n698 B.n697 10.6151
R1800 B.n697 B.n20 10.6151
R1801 B.n693 B.n20 10.6151
R1802 B.n693 B.n692 10.6151
R1803 B.n692 B.n691 10.6151
R1804 B.n691 B.n22 10.6151
R1805 B.n687 B.n22 10.6151
R1806 B.n687 B.n686 10.6151
R1807 B.n686 B.n685 10.6151
R1808 B.n685 B.n24 10.6151
R1809 B.n681 B.n24 10.6151
R1810 B.n681 B.n680 10.6151
R1811 B.n680 B.n679 10.6151
R1812 B.n679 B.n26 10.6151
R1813 B.n675 B.n26 10.6151
R1814 B.n675 B.n674 10.6151
R1815 B.n674 B.n673 10.6151
R1816 B.n673 B.n28 10.6151
R1817 B.n669 B.n28 10.6151
R1818 B.n669 B.n668 10.6151
R1819 B.n668 B.n667 10.6151
R1820 B.n667 B.n30 10.6151
R1821 B.n663 B.n30 10.6151
R1822 B.n663 B.n662 10.6151
R1823 B.n662 B.n661 10.6151
R1824 B.n661 B.n32 10.6151
R1825 B.n657 B.n32 10.6151
R1826 B.n657 B.n656 10.6151
R1827 B.n656 B.n655 10.6151
R1828 B.n655 B.n34 10.6151
R1829 B.n651 B.n34 10.6151
R1830 B.n651 B.n650 10.6151
R1831 B.n650 B.n649 10.6151
R1832 B.n649 B.n36 10.6151
R1833 B.n645 B.n36 10.6151
R1834 B.n645 B.n644 10.6151
R1835 B.n644 B.n643 10.6151
R1836 B.n643 B.n38 10.6151
R1837 B.n639 B.n38 10.6151
R1838 B.n639 B.n638 10.6151
R1839 B.n638 B.n637 10.6151
R1840 B.n637 B.n40 10.6151
R1841 B.n633 B.n40 10.6151
R1842 B.n633 B.n632 10.6151
R1843 B.n632 B.n631 10.6151
R1844 B.n631 B.n42 10.6151
R1845 B.n627 B.n42 10.6151
R1846 B.n627 B.n626 10.6151
R1847 B.n626 B.n625 10.6151
R1848 B.n625 B.n44 10.6151
R1849 B.n621 B.n44 10.6151
R1850 B.n621 B.n620 10.6151
R1851 B.n618 B.n48 10.6151
R1852 B.n614 B.n48 10.6151
R1853 B.n614 B.n613 10.6151
R1854 B.n613 B.n612 10.6151
R1855 B.n612 B.n50 10.6151
R1856 B.n608 B.n50 10.6151
R1857 B.n608 B.n607 10.6151
R1858 B.n607 B.n606 10.6151
R1859 B.n606 B.n52 10.6151
R1860 B.n602 B.n601 10.6151
R1861 B.n601 B.n600 10.6151
R1862 B.n600 B.n57 10.6151
R1863 B.n596 B.n57 10.6151
R1864 B.n596 B.n595 10.6151
R1865 B.n595 B.n594 10.6151
R1866 B.n594 B.n59 10.6151
R1867 B.n590 B.n59 10.6151
R1868 B.n590 B.n589 10.6151
R1869 B.n589 B.n588 10.6151
R1870 B.n588 B.n61 10.6151
R1871 B.n584 B.n61 10.6151
R1872 B.n584 B.n583 10.6151
R1873 B.n583 B.n582 10.6151
R1874 B.n582 B.n63 10.6151
R1875 B.n578 B.n63 10.6151
R1876 B.n578 B.n577 10.6151
R1877 B.n577 B.n576 10.6151
R1878 B.n576 B.n65 10.6151
R1879 B.n572 B.n65 10.6151
R1880 B.n572 B.n571 10.6151
R1881 B.n571 B.n570 10.6151
R1882 B.n570 B.n67 10.6151
R1883 B.n566 B.n67 10.6151
R1884 B.n566 B.n565 10.6151
R1885 B.n565 B.n564 10.6151
R1886 B.n564 B.n69 10.6151
R1887 B.n560 B.n69 10.6151
R1888 B.n560 B.n559 10.6151
R1889 B.n559 B.n558 10.6151
R1890 B.n558 B.n71 10.6151
R1891 B.n554 B.n71 10.6151
R1892 B.n554 B.n553 10.6151
R1893 B.n553 B.n552 10.6151
R1894 B.n552 B.n73 10.6151
R1895 B.n548 B.n73 10.6151
R1896 B.n548 B.n547 10.6151
R1897 B.n547 B.n546 10.6151
R1898 B.n546 B.n75 10.6151
R1899 B.n542 B.n75 10.6151
R1900 B.n542 B.n541 10.6151
R1901 B.n541 B.n540 10.6151
R1902 B.n540 B.n77 10.6151
R1903 B.n536 B.n77 10.6151
R1904 B.n536 B.n535 10.6151
R1905 B.n535 B.n534 10.6151
R1906 B.n534 B.n79 10.6151
R1907 B.n530 B.n79 10.6151
R1908 B.n530 B.n529 10.6151
R1909 B.n529 B.n528 10.6151
R1910 B.n528 B.n81 10.6151
R1911 B.n524 B.n81 10.6151
R1912 B.n524 B.n523 10.6151
R1913 B.n523 B.n522 10.6151
R1914 B.n522 B.n83 10.6151
R1915 B.n518 B.n83 10.6151
R1916 B.n518 B.n517 10.6151
R1917 B.n517 B.n516 10.6151
R1918 B.n516 B.n85 10.6151
R1919 B.n433 B.n432 10.6151
R1920 B.n434 B.n433 10.6151
R1921 B.n434 B.n111 10.6151
R1922 B.n438 B.n111 10.6151
R1923 B.n439 B.n438 10.6151
R1924 B.n440 B.n439 10.6151
R1925 B.n440 B.n109 10.6151
R1926 B.n444 B.n109 10.6151
R1927 B.n445 B.n444 10.6151
R1928 B.n446 B.n445 10.6151
R1929 B.n446 B.n107 10.6151
R1930 B.n450 B.n107 10.6151
R1931 B.n451 B.n450 10.6151
R1932 B.n452 B.n451 10.6151
R1933 B.n452 B.n105 10.6151
R1934 B.n456 B.n105 10.6151
R1935 B.n457 B.n456 10.6151
R1936 B.n458 B.n457 10.6151
R1937 B.n458 B.n103 10.6151
R1938 B.n462 B.n103 10.6151
R1939 B.n463 B.n462 10.6151
R1940 B.n464 B.n463 10.6151
R1941 B.n464 B.n101 10.6151
R1942 B.n468 B.n101 10.6151
R1943 B.n469 B.n468 10.6151
R1944 B.n470 B.n469 10.6151
R1945 B.n470 B.n99 10.6151
R1946 B.n474 B.n99 10.6151
R1947 B.n475 B.n474 10.6151
R1948 B.n476 B.n475 10.6151
R1949 B.n476 B.n97 10.6151
R1950 B.n480 B.n97 10.6151
R1951 B.n481 B.n480 10.6151
R1952 B.n482 B.n481 10.6151
R1953 B.n482 B.n95 10.6151
R1954 B.n486 B.n95 10.6151
R1955 B.n487 B.n486 10.6151
R1956 B.n488 B.n487 10.6151
R1957 B.n488 B.n93 10.6151
R1958 B.n492 B.n93 10.6151
R1959 B.n493 B.n492 10.6151
R1960 B.n494 B.n493 10.6151
R1961 B.n494 B.n91 10.6151
R1962 B.n498 B.n91 10.6151
R1963 B.n499 B.n498 10.6151
R1964 B.n500 B.n499 10.6151
R1965 B.n500 B.n89 10.6151
R1966 B.n504 B.n89 10.6151
R1967 B.n505 B.n504 10.6151
R1968 B.n506 B.n505 10.6151
R1969 B.n506 B.n87 10.6151
R1970 B.n510 B.n87 10.6151
R1971 B.n511 B.n510 10.6151
R1972 B.n512 B.n511 10.6151
R1973 B.n236 B.n235 10.6151
R1974 B.n236 B.n181 10.6151
R1975 B.n240 B.n181 10.6151
R1976 B.n241 B.n240 10.6151
R1977 B.n242 B.n241 10.6151
R1978 B.n242 B.n179 10.6151
R1979 B.n246 B.n179 10.6151
R1980 B.n247 B.n246 10.6151
R1981 B.n248 B.n247 10.6151
R1982 B.n248 B.n177 10.6151
R1983 B.n252 B.n177 10.6151
R1984 B.n253 B.n252 10.6151
R1985 B.n254 B.n253 10.6151
R1986 B.n254 B.n175 10.6151
R1987 B.n258 B.n175 10.6151
R1988 B.n259 B.n258 10.6151
R1989 B.n260 B.n259 10.6151
R1990 B.n260 B.n173 10.6151
R1991 B.n264 B.n173 10.6151
R1992 B.n265 B.n264 10.6151
R1993 B.n266 B.n265 10.6151
R1994 B.n266 B.n171 10.6151
R1995 B.n270 B.n171 10.6151
R1996 B.n271 B.n270 10.6151
R1997 B.n272 B.n271 10.6151
R1998 B.n272 B.n169 10.6151
R1999 B.n276 B.n169 10.6151
R2000 B.n277 B.n276 10.6151
R2001 B.n278 B.n277 10.6151
R2002 B.n278 B.n167 10.6151
R2003 B.n282 B.n167 10.6151
R2004 B.n283 B.n282 10.6151
R2005 B.n284 B.n283 10.6151
R2006 B.n284 B.n165 10.6151
R2007 B.n288 B.n165 10.6151
R2008 B.n289 B.n288 10.6151
R2009 B.n290 B.n289 10.6151
R2010 B.n290 B.n163 10.6151
R2011 B.n294 B.n163 10.6151
R2012 B.n295 B.n294 10.6151
R2013 B.n296 B.n295 10.6151
R2014 B.n296 B.n161 10.6151
R2015 B.n300 B.n161 10.6151
R2016 B.n301 B.n300 10.6151
R2017 B.n302 B.n301 10.6151
R2018 B.n302 B.n159 10.6151
R2019 B.n306 B.n159 10.6151
R2020 B.n307 B.n306 10.6151
R2021 B.n308 B.n307 10.6151
R2022 B.n308 B.n157 10.6151
R2023 B.n312 B.n157 10.6151
R2024 B.n313 B.n312 10.6151
R2025 B.n314 B.n313 10.6151
R2026 B.n314 B.n155 10.6151
R2027 B.n318 B.n155 10.6151
R2028 B.n319 B.n318 10.6151
R2029 B.n320 B.n319 10.6151
R2030 B.n320 B.n153 10.6151
R2031 B.n324 B.n153 10.6151
R2032 B.n327 B.n326 10.6151
R2033 B.n327 B.n149 10.6151
R2034 B.n331 B.n149 10.6151
R2035 B.n332 B.n331 10.6151
R2036 B.n333 B.n332 10.6151
R2037 B.n333 B.n147 10.6151
R2038 B.n337 B.n147 10.6151
R2039 B.n338 B.n337 10.6151
R2040 B.n339 B.n338 10.6151
R2041 B.n343 B.n342 10.6151
R2042 B.n344 B.n343 10.6151
R2043 B.n344 B.n141 10.6151
R2044 B.n348 B.n141 10.6151
R2045 B.n349 B.n348 10.6151
R2046 B.n350 B.n349 10.6151
R2047 B.n350 B.n139 10.6151
R2048 B.n354 B.n139 10.6151
R2049 B.n355 B.n354 10.6151
R2050 B.n356 B.n355 10.6151
R2051 B.n356 B.n137 10.6151
R2052 B.n360 B.n137 10.6151
R2053 B.n361 B.n360 10.6151
R2054 B.n362 B.n361 10.6151
R2055 B.n362 B.n135 10.6151
R2056 B.n366 B.n135 10.6151
R2057 B.n367 B.n366 10.6151
R2058 B.n368 B.n367 10.6151
R2059 B.n368 B.n133 10.6151
R2060 B.n372 B.n133 10.6151
R2061 B.n373 B.n372 10.6151
R2062 B.n374 B.n373 10.6151
R2063 B.n374 B.n131 10.6151
R2064 B.n378 B.n131 10.6151
R2065 B.n379 B.n378 10.6151
R2066 B.n380 B.n379 10.6151
R2067 B.n380 B.n129 10.6151
R2068 B.n384 B.n129 10.6151
R2069 B.n385 B.n384 10.6151
R2070 B.n386 B.n385 10.6151
R2071 B.n386 B.n127 10.6151
R2072 B.n390 B.n127 10.6151
R2073 B.n391 B.n390 10.6151
R2074 B.n392 B.n391 10.6151
R2075 B.n392 B.n125 10.6151
R2076 B.n396 B.n125 10.6151
R2077 B.n397 B.n396 10.6151
R2078 B.n398 B.n397 10.6151
R2079 B.n398 B.n123 10.6151
R2080 B.n402 B.n123 10.6151
R2081 B.n403 B.n402 10.6151
R2082 B.n404 B.n403 10.6151
R2083 B.n404 B.n121 10.6151
R2084 B.n408 B.n121 10.6151
R2085 B.n409 B.n408 10.6151
R2086 B.n410 B.n409 10.6151
R2087 B.n410 B.n119 10.6151
R2088 B.n414 B.n119 10.6151
R2089 B.n415 B.n414 10.6151
R2090 B.n416 B.n415 10.6151
R2091 B.n416 B.n117 10.6151
R2092 B.n420 B.n117 10.6151
R2093 B.n421 B.n420 10.6151
R2094 B.n422 B.n421 10.6151
R2095 B.n422 B.n115 10.6151
R2096 B.n426 B.n115 10.6151
R2097 B.n427 B.n426 10.6151
R2098 B.n428 B.n427 10.6151
R2099 B.n428 B.n113 10.6151
R2100 B.n234 B.n183 10.6151
R2101 B.n230 B.n183 10.6151
R2102 B.n230 B.n229 10.6151
R2103 B.n229 B.n228 10.6151
R2104 B.n228 B.n185 10.6151
R2105 B.n224 B.n185 10.6151
R2106 B.n224 B.n223 10.6151
R2107 B.n223 B.n222 10.6151
R2108 B.n222 B.n187 10.6151
R2109 B.n218 B.n187 10.6151
R2110 B.n218 B.n217 10.6151
R2111 B.n217 B.n216 10.6151
R2112 B.n216 B.n189 10.6151
R2113 B.n212 B.n189 10.6151
R2114 B.n212 B.n211 10.6151
R2115 B.n211 B.n210 10.6151
R2116 B.n210 B.n191 10.6151
R2117 B.n206 B.n191 10.6151
R2118 B.n206 B.n205 10.6151
R2119 B.n205 B.n204 10.6151
R2120 B.n204 B.n193 10.6151
R2121 B.n200 B.n193 10.6151
R2122 B.n200 B.n199 10.6151
R2123 B.n199 B.n198 10.6151
R2124 B.n198 B.n195 10.6151
R2125 B.n195 B.n0 10.6151
R2126 B.n747 B.n1 10.6151
R2127 B.n747 B.n746 10.6151
R2128 B.n746 B.n745 10.6151
R2129 B.n745 B.n4 10.6151
R2130 B.n741 B.n4 10.6151
R2131 B.n741 B.n740 10.6151
R2132 B.n740 B.n739 10.6151
R2133 B.n739 B.n6 10.6151
R2134 B.n735 B.n6 10.6151
R2135 B.n735 B.n734 10.6151
R2136 B.n734 B.n733 10.6151
R2137 B.n733 B.n8 10.6151
R2138 B.n729 B.n8 10.6151
R2139 B.n729 B.n728 10.6151
R2140 B.n728 B.n727 10.6151
R2141 B.n727 B.n10 10.6151
R2142 B.n723 B.n10 10.6151
R2143 B.n723 B.n722 10.6151
R2144 B.n722 B.n721 10.6151
R2145 B.n721 B.n12 10.6151
R2146 B.n717 B.n12 10.6151
R2147 B.n717 B.n716 10.6151
R2148 B.n716 B.n715 10.6151
R2149 B.n715 B.n14 10.6151
R2150 B.n711 B.n14 10.6151
R2151 B.n711 B.n710 10.6151
R2152 B.n620 B.n619 9.36635
R2153 B.n602 B.n56 9.36635
R2154 B.n325 B.n324 9.36635
R2155 B.n342 B.n145 9.36635
R2156 B.n751 B.n0 2.81026
R2157 B.n751 B.n1 2.81026
R2158 B.n619 B.n618 1.24928
R2159 B.n56 B.n52 1.24928
R2160 B.n326 B.n325 1.24928
R2161 B.n339 B.n145 1.24928
R2162 VN.n3 VN.t4 682.338
R2163 VN.n17 VN.t2 682.338
R2164 VN.n4 VN.t1 657.963
R2165 VN.n6 VN.t7 657.963
R2166 VN.n10 VN.t6 657.963
R2167 VN.n12 VN.t0 657.963
R2168 VN.n18 VN.t8 657.963
R2169 VN.n20 VN.t5 657.963
R2170 VN.n24 VN.t9 657.963
R2171 VN.n26 VN.t3 657.963
R2172 VN.n13 VN.n12 161.3
R2173 VN.n27 VN.n26 161.3
R2174 VN.n25 VN.n14 161.3
R2175 VN.n24 VN.n23 161.3
R2176 VN.n22 VN.n15 161.3
R2177 VN.n21 VN.n20 161.3
R2178 VN.n19 VN.n16 161.3
R2179 VN.n11 VN.n0 161.3
R2180 VN.n10 VN.n9 161.3
R2181 VN.n8 VN.n1 161.3
R2182 VN.n7 VN.n6 161.3
R2183 VN.n5 VN.n2 161.3
R2184 VN VN.n27 48.1539
R2185 VN.n17 VN.n16 44.9377
R2186 VN.n3 VN.n2 44.9377
R2187 VN.n12 VN.n11 37.246
R2188 VN.n26 VN.n25 37.246
R2189 VN.n5 VN.n4 28.4823
R2190 VN.n10 VN.n1 28.4823
R2191 VN.n19 VN.n18 28.4823
R2192 VN.n24 VN.n15 28.4823
R2193 VN.n6 VN.n5 19.7187
R2194 VN.n6 VN.n1 19.7187
R2195 VN.n20 VN.n19 19.7187
R2196 VN.n20 VN.n15 19.7187
R2197 VN.n4 VN.n3 17.0522
R2198 VN.n18 VN.n17 17.0522
R2199 VN.n11 VN.n10 10.955
R2200 VN.n25 VN.n24 10.955
R2201 VN.n27 VN.n14 0.189894
R2202 VN.n23 VN.n14 0.189894
R2203 VN.n23 VN.n22 0.189894
R2204 VN.n22 VN.n21 0.189894
R2205 VN.n21 VN.n16 0.189894
R2206 VN.n7 VN.n2 0.189894
R2207 VN.n8 VN.n7 0.189894
R2208 VN.n9 VN.n8 0.189894
R2209 VN.n9 VN.n0 0.189894
R2210 VN.n13 VN.n0 0.189894
R2211 VN VN.n13 0.0516364
R2212 VDD2.n201 VDD2.n105 756.745
R2213 VDD2.n96 VDD2.n0 756.745
R2214 VDD2.n202 VDD2.n201 585
R2215 VDD2.n200 VDD2.n199 585
R2216 VDD2.n109 VDD2.n108 585
R2217 VDD2.n194 VDD2.n193 585
R2218 VDD2.n192 VDD2.n191 585
R2219 VDD2.n113 VDD2.n112 585
R2220 VDD2.n186 VDD2.n185 585
R2221 VDD2.n184 VDD2.n115 585
R2222 VDD2.n183 VDD2.n182 585
R2223 VDD2.n118 VDD2.n116 585
R2224 VDD2.n177 VDD2.n176 585
R2225 VDD2.n175 VDD2.n174 585
R2226 VDD2.n122 VDD2.n121 585
R2227 VDD2.n169 VDD2.n168 585
R2228 VDD2.n167 VDD2.n166 585
R2229 VDD2.n126 VDD2.n125 585
R2230 VDD2.n161 VDD2.n160 585
R2231 VDD2.n159 VDD2.n158 585
R2232 VDD2.n130 VDD2.n129 585
R2233 VDD2.n153 VDD2.n152 585
R2234 VDD2.n151 VDD2.n150 585
R2235 VDD2.n134 VDD2.n133 585
R2236 VDD2.n145 VDD2.n144 585
R2237 VDD2.n143 VDD2.n142 585
R2238 VDD2.n138 VDD2.n137 585
R2239 VDD2.n32 VDD2.n31 585
R2240 VDD2.n37 VDD2.n36 585
R2241 VDD2.n39 VDD2.n38 585
R2242 VDD2.n28 VDD2.n27 585
R2243 VDD2.n45 VDD2.n44 585
R2244 VDD2.n47 VDD2.n46 585
R2245 VDD2.n24 VDD2.n23 585
R2246 VDD2.n53 VDD2.n52 585
R2247 VDD2.n55 VDD2.n54 585
R2248 VDD2.n20 VDD2.n19 585
R2249 VDD2.n61 VDD2.n60 585
R2250 VDD2.n63 VDD2.n62 585
R2251 VDD2.n16 VDD2.n15 585
R2252 VDD2.n69 VDD2.n68 585
R2253 VDD2.n71 VDD2.n70 585
R2254 VDD2.n12 VDD2.n11 585
R2255 VDD2.n78 VDD2.n77 585
R2256 VDD2.n79 VDD2.n10 585
R2257 VDD2.n81 VDD2.n80 585
R2258 VDD2.n8 VDD2.n7 585
R2259 VDD2.n87 VDD2.n86 585
R2260 VDD2.n89 VDD2.n88 585
R2261 VDD2.n4 VDD2.n3 585
R2262 VDD2.n95 VDD2.n94 585
R2263 VDD2.n97 VDD2.n96 585
R2264 VDD2.n139 VDD2.t6 327.466
R2265 VDD2.n33 VDD2.t5 327.466
R2266 VDD2.n201 VDD2.n200 171.744
R2267 VDD2.n200 VDD2.n108 171.744
R2268 VDD2.n193 VDD2.n108 171.744
R2269 VDD2.n193 VDD2.n192 171.744
R2270 VDD2.n192 VDD2.n112 171.744
R2271 VDD2.n185 VDD2.n112 171.744
R2272 VDD2.n185 VDD2.n184 171.744
R2273 VDD2.n184 VDD2.n183 171.744
R2274 VDD2.n183 VDD2.n116 171.744
R2275 VDD2.n176 VDD2.n116 171.744
R2276 VDD2.n176 VDD2.n175 171.744
R2277 VDD2.n175 VDD2.n121 171.744
R2278 VDD2.n168 VDD2.n121 171.744
R2279 VDD2.n168 VDD2.n167 171.744
R2280 VDD2.n167 VDD2.n125 171.744
R2281 VDD2.n160 VDD2.n125 171.744
R2282 VDD2.n160 VDD2.n159 171.744
R2283 VDD2.n159 VDD2.n129 171.744
R2284 VDD2.n152 VDD2.n129 171.744
R2285 VDD2.n152 VDD2.n151 171.744
R2286 VDD2.n151 VDD2.n133 171.744
R2287 VDD2.n144 VDD2.n133 171.744
R2288 VDD2.n144 VDD2.n143 171.744
R2289 VDD2.n143 VDD2.n137 171.744
R2290 VDD2.n37 VDD2.n31 171.744
R2291 VDD2.n38 VDD2.n37 171.744
R2292 VDD2.n38 VDD2.n27 171.744
R2293 VDD2.n45 VDD2.n27 171.744
R2294 VDD2.n46 VDD2.n45 171.744
R2295 VDD2.n46 VDD2.n23 171.744
R2296 VDD2.n53 VDD2.n23 171.744
R2297 VDD2.n54 VDD2.n53 171.744
R2298 VDD2.n54 VDD2.n19 171.744
R2299 VDD2.n61 VDD2.n19 171.744
R2300 VDD2.n62 VDD2.n61 171.744
R2301 VDD2.n62 VDD2.n15 171.744
R2302 VDD2.n69 VDD2.n15 171.744
R2303 VDD2.n70 VDD2.n69 171.744
R2304 VDD2.n70 VDD2.n11 171.744
R2305 VDD2.n78 VDD2.n11 171.744
R2306 VDD2.n79 VDD2.n78 171.744
R2307 VDD2.n80 VDD2.n79 171.744
R2308 VDD2.n80 VDD2.n7 171.744
R2309 VDD2.n87 VDD2.n7 171.744
R2310 VDD2.n88 VDD2.n87 171.744
R2311 VDD2.n88 VDD2.n3 171.744
R2312 VDD2.n95 VDD2.n3 171.744
R2313 VDD2.n96 VDD2.n95 171.744
R2314 VDD2.t6 VDD2.n137 85.8723
R2315 VDD2.t5 VDD2.n31 85.8723
R2316 VDD2.n104 VDD2.n103 70.4813
R2317 VDD2 VDD2.n209 70.4785
R2318 VDD2.n208 VDD2.n207 69.8515
R2319 VDD2.n102 VDD2.n101 69.8513
R2320 VDD2.n102 VDD2.n100 50.9416
R2321 VDD2.n206 VDD2.n205 50.0278
R2322 VDD2.n206 VDD2.n104 43.8317
R2323 VDD2.n139 VDD2.n138 16.3895
R2324 VDD2.n33 VDD2.n32 16.3895
R2325 VDD2.n186 VDD2.n115 13.1884
R2326 VDD2.n81 VDD2.n10 13.1884
R2327 VDD2.n187 VDD2.n113 12.8005
R2328 VDD2.n182 VDD2.n117 12.8005
R2329 VDD2.n142 VDD2.n141 12.8005
R2330 VDD2.n36 VDD2.n35 12.8005
R2331 VDD2.n77 VDD2.n76 12.8005
R2332 VDD2.n82 VDD2.n8 12.8005
R2333 VDD2.n191 VDD2.n190 12.0247
R2334 VDD2.n181 VDD2.n118 12.0247
R2335 VDD2.n145 VDD2.n136 12.0247
R2336 VDD2.n39 VDD2.n30 12.0247
R2337 VDD2.n75 VDD2.n12 12.0247
R2338 VDD2.n86 VDD2.n85 12.0247
R2339 VDD2.n194 VDD2.n111 11.249
R2340 VDD2.n178 VDD2.n177 11.249
R2341 VDD2.n146 VDD2.n134 11.249
R2342 VDD2.n40 VDD2.n28 11.249
R2343 VDD2.n72 VDD2.n71 11.249
R2344 VDD2.n89 VDD2.n6 11.249
R2345 VDD2.n195 VDD2.n109 10.4732
R2346 VDD2.n174 VDD2.n120 10.4732
R2347 VDD2.n150 VDD2.n149 10.4732
R2348 VDD2.n44 VDD2.n43 10.4732
R2349 VDD2.n68 VDD2.n14 10.4732
R2350 VDD2.n90 VDD2.n4 10.4732
R2351 VDD2.n199 VDD2.n198 9.69747
R2352 VDD2.n173 VDD2.n122 9.69747
R2353 VDD2.n153 VDD2.n132 9.69747
R2354 VDD2.n47 VDD2.n26 9.69747
R2355 VDD2.n67 VDD2.n16 9.69747
R2356 VDD2.n94 VDD2.n93 9.69747
R2357 VDD2.n205 VDD2.n204 9.45567
R2358 VDD2.n100 VDD2.n99 9.45567
R2359 VDD2.n165 VDD2.n164 9.3005
R2360 VDD2.n124 VDD2.n123 9.3005
R2361 VDD2.n171 VDD2.n170 9.3005
R2362 VDD2.n173 VDD2.n172 9.3005
R2363 VDD2.n120 VDD2.n119 9.3005
R2364 VDD2.n179 VDD2.n178 9.3005
R2365 VDD2.n181 VDD2.n180 9.3005
R2366 VDD2.n117 VDD2.n114 9.3005
R2367 VDD2.n204 VDD2.n203 9.3005
R2368 VDD2.n107 VDD2.n106 9.3005
R2369 VDD2.n198 VDD2.n197 9.3005
R2370 VDD2.n196 VDD2.n195 9.3005
R2371 VDD2.n111 VDD2.n110 9.3005
R2372 VDD2.n190 VDD2.n189 9.3005
R2373 VDD2.n188 VDD2.n187 9.3005
R2374 VDD2.n163 VDD2.n162 9.3005
R2375 VDD2.n128 VDD2.n127 9.3005
R2376 VDD2.n157 VDD2.n156 9.3005
R2377 VDD2.n155 VDD2.n154 9.3005
R2378 VDD2.n132 VDD2.n131 9.3005
R2379 VDD2.n149 VDD2.n148 9.3005
R2380 VDD2.n147 VDD2.n146 9.3005
R2381 VDD2.n136 VDD2.n135 9.3005
R2382 VDD2.n141 VDD2.n140 9.3005
R2383 VDD2.n99 VDD2.n98 9.3005
R2384 VDD2.n2 VDD2.n1 9.3005
R2385 VDD2.n93 VDD2.n92 9.3005
R2386 VDD2.n91 VDD2.n90 9.3005
R2387 VDD2.n6 VDD2.n5 9.3005
R2388 VDD2.n85 VDD2.n84 9.3005
R2389 VDD2.n83 VDD2.n82 9.3005
R2390 VDD2.n22 VDD2.n21 9.3005
R2391 VDD2.n51 VDD2.n50 9.3005
R2392 VDD2.n49 VDD2.n48 9.3005
R2393 VDD2.n26 VDD2.n25 9.3005
R2394 VDD2.n43 VDD2.n42 9.3005
R2395 VDD2.n41 VDD2.n40 9.3005
R2396 VDD2.n30 VDD2.n29 9.3005
R2397 VDD2.n35 VDD2.n34 9.3005
R2398 VDD2.n57 VDD2.n56 9.3005
R2399 VDD2.n59 VDD2.n58 9.3005
R2400 VDD2.n18 VDD2.n17 9.3005
R2401 VDD2.n65 VDD2.n64 9.3005
R2402 VDD2.n67 VDD2.n66 9.3005
R2403 VDD2.n14 VDD2.n13 9.3005
R2404 VDD2.n73 VDD2.n72 9.3005
R2405 VDD2.n75 VDD2.n74 9.3005
R2406 VDD2.n76 VDD2.n9 9.3005
R2407 VDD2.n202 VDD2.n107 8.92171
R2408 VDD2.n170 VDD2.n169 8.92171
R2409 VDD2.n154 VDD2.n130 8.92171
R2410 VDD2.n48 VDD2.n24 8.92171
R2411 VDD2.n64 VDD2.n63 8.92171
R2412 VDD2.n97 VDD2.n2 8.92171
R2413 VDD2.n203 VDD2.n105 8.14595
R2414 VDD2.n166 VDD2.n124 8.14595
R2415 VDD2.n158 VDD2.n157 8.14595
R2416 VDD2.n52 VDD2.n51 8.14595
R2417 VDD2.n60 VDD2.n18 8.14595
R2418 VDD2.n98 VDD2.n0 8.14595
R2419 VDD2.n165 VDD2.n126 7.3702
R2420 VDD2.n161 VDD2.n128 7.3702
R2421 VDD2.n55 VDD2.n22 7.3702
R2422 VDD2.n59 VDD2.n20 7.3702
R2423 VDD2.n162 VDD2.n126 6.59444
R2424 VDD2.n162 VDD2.n161 6.59444
R2425 VDD2.n56 VDD2.n55 6.59444
R2426 VDD2.n56 VDD2.n20 6.59444
R2427 VDD2.n205 VDD2.n105 5.81868
R2428 VDD2.n166 VDD2.n165 5.81868
R2429 VDD2.n158 VDD2.n128 5.81868
R2430 VDD2.n52 VDD2.n22 5.81868
R2431 VDD2.n60 VDD2.n59 5.81868
R2432 VDD2.n100 VDD2.n0 5.81868
R2433 VDD2.n203 VDD2.n202 5.04292
R2434 VDD2.n169 VDD2.n124 5.04292
R2435 VDD2.n157 VDD2.n130 5.04292
R2436 VDD2.n51 VDD2.n24 5.04292
R2437 VDD2.n63 VDD2.n18 5.04292
R2438 VDD2.n98 VDD2.n97 5.04292
R2439 VDD2.n199 VDD2.n107 4.26717
R2440 VDD2.n170 VDD2.n122 4.26717
R2441 VDD2.n154 VDD2.n153 4.26717
R2442 VDD2.n48 VDD2.n47 4.26717
R2443 VDD2.n64 VDD2.n16 4.26717
R2444 VDD2.n94 VDD2.n2 4.26717
R2445 VDD2.n140 VDD2.n139 3.70982
R2446 VDD2.n34 VDD2.n33 3.70982
R2447 VDD2.n198 VDD2.n109 3.49141
R2448 VDD2.n174 VDD2.n173 3.49141
R2449 VDD2.n150 VDD2.n132 3.49141
R2450 VDD2.n44 VDD2.n26 3.49141
R2451 VDD2.n68 VDD2.n67 3.49141
R2452 VDD2.n93 VDD2.n4 3.49141
R2453 VDD2.n195 VDD2.n194 2.71565
R2454 VDD2.n177 VDD2.n120 2.71565
R2455 VDD2.n149 VDD2.n134 2.71565
R2456 VDD2.n43 VDD2.n28 2.71565
R2457 VDD2.n71 VDD2.n14 2.71565
R2458 VDD2.n90 VDD2.n89 2.71565
R2459 VDD2.n191 VDD2.n111 1.93989
R2460 VDD2.n178 VDD2.n118 1.93989
R2461 VDD2.n146 VDD2.n145 1.93989
R2462 VDD2.n40 VDD2.n39 1.93989
R2463 VDD2.n72 VDD2.n12 1.93989
R2464 VDD2.n86 VDD2.n6 1.93989
R2465 VDD2.n209 VDD2.t1 1.77673
R2466 VDD2.n209 VDD2.t7 1.77673
R2467 VDD2.n207 VDD2.t0 1.77673
R2468 VDD2.n207 VDD2.t4 1.77673
R2469 VDD2.n103 VDD2.t3 1.77673
R2470 VDD2.n103 VDD2.t9 1.77673
R2471 VDD2.n101 VDD2.t8 1.77673
R2472 VDD2.n101 VDD2.t2 1.77673
R2473 VDD2.n190 VDD2.n113 1.16414
R2474 VDD2.n182 VDD2.n181 1.16414
R2475 VDD2.n142 VDD2.n136 1.16414
R2476 VDD2.n36 VDD2.n30 1.16414
R2477 VDD2.n77 VDD2.n75 1.16414
R2478 VDD2.n85 VDD2.n8 1.16414
R2479 VDD2.n208 VDD2.n206 0.914293
R2480 VDD2.n187 VDD2.n186 0.388379
R2481 VDD2.n117 VDD2.n115 0.388379
R2482 VDD2.n141 VDD2.n138 0.388379
R2483 VDD2.n35 VDD2.n32 0.388379
R2484 VDD2.n76 VDD2.n10 0.388379
R2485 VDD2.n82 VDD2.n81 0.388379
R2486 VDD2 VDD2.n208 0.287138
R2487 VDD2.n104 VDD2.n102 0.173602
R2488 VDD2.n204 VDD2.n106 0.155672
R2489 VDD2.n197 VDD2.n106 0.155672
R2490 VDD2.n197 VDD2.n196 0.155672
R2491 VDD2.n196 VDD2.n110 0.155672
R2492 VDD2.n189 VDD2.n110 0.155672
R2493 VDD2.n189 VDD2.n188 0.155672
R2494 VDD2.n188 VDD2.n114 0.155672
R2495 VDD2.n180 VDD2.n114 0.155672
R2496 VDD2.n180 VDD2.n179 0.155672
R2497 VDD2.n179 VDD2.n119 0.155672
R2498 VDD2.n172 VDD2.n119 0.155672
R2499 VDD2.n172 VDD2.n171 0.155672
R2500 VDD2.n171 VDD2.n123 0.155672
R2501 VDD2.n164 VDD2.n123 0.155672
R2502 VDD2.n164 VDD2.n163 0.155672
R2503 VDD2.n163 VDD2.n127 0.155672
R2504 VDD2.n156 VDD2.n127 0.155672
R2505 VDD2.n156 VDD2.n155 0.155672
R2506 VDD2.n155 VDD2.n131 0.155672
R2507 VDD2.n148 VDD2.n131 0.155672
R2508 VDD2.n148 VDD2.n147 0.155672
R2509 VDD2.n147 VDD2.n135 0.155672
R2510 VDD2.n140 VDD2.n135 0.155672
R2511 VDD2.n34 VDD2.n29 0.155672
R2512 VDD2.n41 VDD2.n29 0.155672
R2513 VDD2.n42 VDD2.n41 0.155672
R2514 VDD2.n42 VDD2.n25 0.155672
R2515 VDD2.n49 VDD2.n25 0.155672
R2516 VDD2.n50 VDD2.n49 0.155672
R2517 VDD2.n50 VDD2.n21 0.155672
R2518 VDD2.n57 VDD2.n21 0.155672
R2519 VDD2.n58 VDD2.n57 0.155672
R2520 VDD2.n58 VDD2.n17 0.155672
R2521 VDD2.n65 VDD2.n17 0.155672
R2522 VDD2.n66 VDD2.n65 0.155672
R2523 VDD2.n66 VDD2.n13 0.155672
R2524 VDD2.n73 VDD2.n13 0.155672
R2525 VDD2.n74 VDD2.n73 0.155672
R2526 VDD2.n74 VDD2.n9 0.155672
R2527 VDD2.n83 VDD2.n9 0.155672
R2528 VDD2.n84 VDD2.n83 0.155672
R2529 VDD2.n84 VDD2.n5 0.155672
R2530 VDD2.n91 VDD2.n5 0.155672
R2531 VDD2.n92 VDD2.n91 0.155672
R2532 VDD2.n92 VDD2.n1 0.155672
R2533 VDD2.n99 VDD2.n1 0.155672
C0 B VP 1.35319f
C1 VDD2 VN 10.2058f
C2 VDD2 w_n2242_n4628# 2.56024f
C3 VTAIL VDD1 19.9433f
C4 B VN 0.882367f
C5 w_n2242_n4628# B 9.170759f
C6 VP VDD1 10.3962f
C7 VN VDD1 0.149158f
C8 VP VTAIL 9.83488f
C9 w_n2242_n4628# VDD1 2.51409f
C10 VN VTAIL 9.82003f
C11 w_n2242_n4628# VTAIL 3.9758f
C12 VP VN 6.80299f
C13 w_n2242_n4628# VP 4.62534f
C14 w_n2242_n4628# VN 4.33922f
C15 VDD2 B 2.22138f
C16 VDD2 VDD1 0.991158f
C17 B VDD1 2.17595f
C18 VDD2 VTAIL 19.974401f
C19 VDD2 VP 0.34641f
C20 B VTAIL 3.88167f
C21 VDD2 VSUBS 1.726496f
C22 VDD1 VSUBS 1.375886f
C23 VTAIL VSUBS 0.969134f
C24 VN VSUBS 5.43891f
C25 VP VSUBS 2.093827f
C26 B VSUBS 3.582797f
C27 w_n2242_n4628# VSUBS 0.126852p
C28 VDD2.n0 VSUBS 0.031528f
C29 VDD2.n1 VSUBS 0.028149f
C30 VDD2.n2 VSUBS 0.015126f
C31 VDD2.n3 VSUBS 0.035752f
C32 VDD2.n4 VSUBS 0.016016f
C33 VDD2.n5 VSUBS 0.028149f
C34 VDD2.n6 VSUBS 0.015126f
C35 VDD2.n7 VSUBS 0.035752f
C36 VDD2.n8 VSUBS 0.016016f
C37 VDD2.n9 VSUBS 0.028149f
C38 VDD2.n10 VSUBS 0.015571f
C39 VDD2.n11 VSUBS 0.035752f
C40 VDD2.n12 VSUBS 0.016016f
C41 VDD2.n13 VSUBS 0.028149f
C42 VDD2.n14 VSUBS 0.015126f
C43 VDD2.n15 VSUBS 0.035752f
C44 VDD2.n16 VSUBS 0.016016f
C45 VDD2.n17 VSUBS 0.028149f
C46 VDD2.n18 VSUBS 0.015126f
C47 VDD2.n19 VSUBS 0.035752f
C48 VDD2.n20 VSUBS 0.016016f
C49 VDD2.n21 VSUBS 0.028149f
C50 VDD2.n22 VSUBS 0.015126f
C51 VDD2.n23 VSUBS 0.035752f
C52 VDD2.n24 VSUBS 0.016016f
C53 VDD2.n25 VSUBS 0.028149f
C54 VDD2.n26 VSUBS 0.015126f
C55 VDD2.n27 VSUBS 0.035752f
C56 VDD2.n28 VSUBS 0.016016f
C57 VDD2.n29 VSUBS 0.028149f
C58 VDD2.n30 VSUBS 0.015126f
C59 VDD2.n31 VSUBS 0.026814f
C60 VDD2.n32 VSUBS 0.022744f
C61 VDD2.t5 VSUBS 0.076769f
C62 VDD2.n33 VSUBS 0.225822f
C63 VDD2.n34 VSUBS 2.21904f
C64 VDD2.n35 VSUBS 0.015126f
C65 VDD2.n36 VSUBS 0.016016f
C66 VDD2.n37 VSUBS 0.035752f
C67 VDD2.n38 VSUBS 0.035752f
C68 VDD2.n39 VSUBS 0.016016f
C69 VDD2.n40 VSUBS 0.015126f
C70 VDD2.n41 VSUBS 0.028149f
C71 VDD2.n42 VSUBS 0.028149f
C72 VDD2.n43 VSUBS 0.015126f
C73 VDD2.n44 VSUBS 0.016016f
C74 VDD2.n45 VSUBS 0.035752f
C75 VDD2.n46 VSUBS 0.035752f
C76 VDD2.n47 VSUBS 0.016016f
C77 VDD2.n48 VSUBS 0.015126f
C78 VDD2.n49 VSUBS 0.028149f
C79 VDD2.n50 VSUBS 0.028149f
C80 VDD2.n51 VSUBS 0.015126f
C81 VDD2.n52 VSUBS 0.016016f
C82 VDD2.n53 VSUBS 0.035752f
C83 VDD2.n54 VSUBS 0.035752f
C84 VDD2.n55 VSUBS 0.016016f
C85 VDD2.n56 VSUBS 0.015126f
C86 VDD2.n57 VSUBS 0.028149f
C87 VDD2.n58 VSUBS 0.028149f
C88 VDD2.n59 VSUBS 0.015126f
C89 VDD2.n60 VSUBS 0.016016f
C90 VDD2.n61 VSUBS 0.035752f
C91 VDD2.n62 VSUBS 0.035752f
C92 VDD2.n63 VSUBS 0.016016f
C93 VDD2.n64 VSUBS 0.015126f
C94 VDD2.n65 VSUBS 0.028149f
C95 VDD2.n66 VSUBS 0.028149f
C96 VDD2.n67 VSUBS 0.015126f
C97 VDD2.n68 VSUBS 0.016016f
C98 VDD2.n69 VSUBS 0.035752f
C99 VDD2.n70 VSUBS 0.035752f
C100 VDD2.n71 VSUBS 0.016016f
C101 VDD2.n72 VSUBS 0.015126f
C102 VDD2.n73 VSUBS 0.028149f
C103 VDD2.n74 VSUBS 0.028149f
C104 VDD2.n75 VSUBS 0.015126f
C105 VDD2.n76 VSUBS 0.015126f
C106 VDD2.n77 VSUBS 0.016016f
C107 VDD2.n78 VSUBS 0.035752f
C108 VDD2.n79 VSUBS 0.035752f
C109 VDD2.n80 VSUBS 0.035752f
C110 VDD2.n81 VSUBS 0.015571f
C111 VDD2.n82 VSUBS 0.015126f
C112 VDD2.n83 VSUBS 0.028149f
C113 VDD2.n84 VSUBS 0.028149f
C114 VDD2.n85 VSUBS 0.015126f
C115 VDD2.n86 VSUBS 0.016016f
C116 VDD2.n87 VSUBS 0.035752f
C117 VDD2.n88 VSUBS 0.035752f
C118 VDD2.n89 VSUBS 0.016016f
C119 VDD2.n90 VSUBS 0.015126f
C120 VDD2.n91 VSUBS 0.028149f
C121 VDD2.n92 VSUBS 0.028149f
C122 VDD2.n93 VSUBS 0.015126f
C123 VDD2.n94 VSUBS 0.016016f
C124 VDD2.n95 VSUBS 0.035752f
C125 VDD2.n96 VSUBS 0.088589f
C126 VDD2.n97 VSUBS 0.016016f
C127 VDD2.n98 VSUBS 0.015126f
C128 VDD2.n99 VSUBS 0.067371f
C129 VDD2.n100 VSUBS 0.066612f
C130 VDD2.t8 VSUBS 0.407062f
C131 VDD2.t2 VSUBS 0.407062f
C132 VDD2.n101 VSUBS 3.39335f
C133 VDD2.n102 VSUBS 0.789805f
C134 VDD2.t3 VSUBS 0.407062f
C135 VDD2.t9 VSUBS 0.407062f
C136 VDD2.n103 VSUBS 3.39965f
C137 VDD2.n104 VSUBS 2.91763f
C138 VDD2.n105 VSUBS 0.031528f
C139 VDD2.n106 VSUBS 0.028149f
C140 VDD2.n107 VSUBS 0.015126f
C141 VDD2.n108 VSUBS 0.035752f
C142 VDD2.n109 VSUBS 0.016016f
C143 VDD2.n110 VSUBS 0.028149f
C144 VDD2.n111 VSUBS 0.015126f
C145 VDD2.n112 VSUBS 0.035752f
C146 VDD2.n113 VSUBS 0.016016f
C147 VDD2.n114 VSUBS 0.028149f
C148 VDD2.n115 VSUBS 0.015571f
C149 VDD2.n116 VSUBS 0.035752f
C150 VDD2.n117 VSUBS 0.015126f
C151 VDD2.n118 VSUBS 0.016016f
C152 VDD2.n119 VSUBS 0.028149f
C153 VDD2.n120 VSUBS 0.015126f
C154 VDD2.n121 VSUBS 0.035752f
C155 VDD2.n122 VSUBS 0.016016f
C156 VDD2.n123 VSUBS 0.028149f
C157 VDD2.n124 VSUBS 0.015126f
C158 VDD2.n125 VSUBS 0.035752f
C159 VDD2.n126 VSUBS 0.016016f
C160 VDD2.n127 VSUBS 0.028149f
C161 VDD2.n128 VSUBS 0.015126f
C162 VDD2.n129 VSUBS 0.035752f
C163 VDD2.n130 VSUBS 0.016016f
C164 VDD2.n131 VSUBS 0.028149f
C165 VDD2.n132 VSUBS 0.015126f
C166 VDD2.n133 VSUBS 0.035752f
C167 VDD2.n134 VSUBS 0.016016f
C168 VDD2.n135 VSUBS 0.028149f
C169 VDD2.n136 VSUBS 0.015126f
C170 VDD2.n137 VSUBS 0.026814f
C171 VDD2.n138 VSUBS 0.022744f
C172 VDD2.t6 VSUBS 0.076769f
C173 VDD2.n139 VSUBS 0.225822f
C174 VDD2.n140 VSUBS 2.21904f
C175 VDD2.n141 VSUBS 0.015126f
C176 VDD2.n142 VSUBS 0.016016f
C177 VDD2.n143 VSUBS 0.035752f
C178 VDD2.n144 VSUBS 0.035752f
C179 VDD2.n145 VSUBS 0.016016f
C180 VDD2.n146 VSUBS 0.015126f
C181 VDD2.n147 VSUBS 0.028149f
C182 VDD2.n148 VSUBS 0.028149f
C183 VDD2.n149 VSUBS 0.015126f
C184 VDD2.n150 VSUBS 0.016016f
C185 VDD2.n151 VSUBS 0.035752f
C186 VDD2.n152 VSUBS 0.035752f
C187 VDD2.n153 VSUBS 0.016016f
C188 VDD2.n154 VSUBS 0.015126f
C189 VDD2.n155 VSUBS 0.028149f
C190 VDD2.n156 VSUBS 0.028149f
C191 VDD2.n157 VSUBS 0.015126f
C192 VDD2.n158 VSUBS 0.016016f
C193 VDD2.n159 VSUBS 0.035752f
C194 VDD2.n160 VSUBS 0.035752f
C195 VDD2.n161 VSUBS 0.016016f
C196 VDD2.n162 VSUBS 0.015126f
C197 VDD2.n163 VSUBS 0.028149f
C198 VDD2.n164 VSUBS 0.028149f
C199 VDD2.n165 VSUBS 0.015126f
C200 VDD2.n166 VSUBS 0.016016f
C201 VDD2.n167 VSUBS 0.035752f
C202 VDD2.n168 VSUBS 0.035752f
C203 VDD2.n169 VSUBS 0.016016f
C204 VDD2.n170 VSUBS 0.015126f
C205 VDD2.n171 VSUBS 0.028149f
C206 VDD2.n172 VSUBS 0.028149f
C207 VDD2.n173 VSUBS 0.015126f
C208 VDD2.n174 VSUBS 0.016016f
C209 VDD2.n175 VSUBS 0.035752f
C210 VDD2.n176 VSUBS 0.035752f
C211 VDD2.n177 VSUBS 0.016016f
C212 VDD2.n178 VSUBS 0.015126f
C213 VDD2.n179 VSUBS 0.028149f
C214 VDD2.n180 VSUBS 0.028149f
C215 VDD2.n181 VSUBS 0.015126f
C216 VDD2.n182 VSUBS 0.016016f
C217 VDD2.n183 VSUBS 0.035752f
C218 VDD2.n184 VSUBS 0.035752f
C219 VDD2.n185 VSUBS 0.035752f
C220 VDD2.n186 VSUBS 0.015571f
C221 VDD2.n187 VSUBS 0.015126f
C222 VDD2.n188 VSUBS 0.028149f
C223 VDD2.n189 VSUBS 0.028149f
C224 VDD2.n190 VSUBS 0.015126f
C225 VDD2.n191 VSUBS 0.016016f
C226 VDD2.n192 VSUBS 0.035752f
C227 VDD2.n193 VSUBS 0.035752f
C228 VDD2.n194 VSUBS 0.016016f
C229 VDD2.n195 VSUBS 0.015126f
C230 VDD2.n196 VSUBS 0.028149f
C231 VDD2.n197 VSUBS 0.028149f
C232 VDD2.n198 VSUBS 0.015126f
C233 VDD2.n199 VSUBS 0.016016f
C234 VDD2.n200 VSUBS 0.035752f
C235 VDD2.n201 VSUBS 0.088589f
C236 VDD2.n202 VSUBS 0.016016f
C237 VDD2.n203 VSUBS 0.015126f
C238 VDD2.n204 VSUBS 0.067371f
C239 VDD2.n205 VSUBS 0.064129f
C240 VDD2.n206 VSUBS 2.98621f
C241 VDD2.t0 VSUBS 0.407062f
C242 VDD2.t4 VSUBS 0.407062f
C243 VDD2.n207 VSUBS 3.39337f
C244 VDD2.n208 VSUBS 0.660397f
C245 VDD2.t1 VSUBS 0.407062f
C246 VDD2.t7 VSUBS 0.407062f
C247 VDD2.n209 VSUBS 3.39961f
C248 VN.n0 VSUBS 0.04837f
C249 VN.n1 VSUBS 0.010976f
C250 VN.n2 VSUBS 0.206467f
C251 VN.t4 VSUBS 1.85631f
C252 VN.n3 VSUBS 0.668662f
C253 VN.t1 VSUBS 1.83168f
C254 VN.n4 VSUBS 0.694984f
C255 VN.n5 VSUBS 0.010976f
C256 VN.t7 VSUBS 1.83168f
C257 VN.n6 VSUBS 0.688357f
C258 VN.n7 VSUBS 0.04837f
C259 VN.n8 VSUBS 0.04837f
C260 VN.n9 VSUBS 0.04837f
C261 VN.t6 VSUBS 1.83168f
C262 VN.n10 VSUBS 0.688357f
C263 VN.n11 VSUBS 0.010976f
C264 VN.t0 VSUBS 1.83168f
C265 VN.n12 VSUBS 0.68791f
C266 VN.n13 VSUBS 0.037485f
C267 VN.n14 VSUBS 0.04837f
C268 VN.n15 VSUBS 0.010976f
C269 VN.t9 VSUBS 1.83168f
C270 VN.n16 VSUBS 0.206467f
C271 VN.t2 VSUBS 1.85631f
C272 VN.n17 VSUBS 0.668662f
C273 VN.t8 VSUBS 1.83168f
C274 VN.n18 VSUBS 0.694984f
C275 VN.n19 VSUBS 0.010976f
C276 VN.t5 VSUBS 1.83168f
C277 VN.n20 VSUBS 0.688357f
C278 VN.n21 VSUBS 0.04837f
C279 VN.n22 VSUBS 0.04837f
C280 VN.n23 VSUBS 0.04837f
C281 VN.n24 VSUBS 0.688357f
C282 VN.n25 VSUBS 0.010976f
C283 VN.t3 VSUBS 1.83168f
C284 VN.n26 VSUBS 0.68791f
C285 VN.n27 VSUBS 2.48509f
C286 B.n0 VSUBS 0.00572f
C287 B.n1 VSUBS 0.00572f
C288 B.n2 VSUBS 0.009046f
C289 B.n3 VSUBS 0.009046f
C290 B.n4 VSUBS 0.009046f
C291 B.n5 VSUBS 0.009046f
C292 B.n6 VSUBS 0.009046f
C293 B.n7 VSUBS 0.009046f
C294 B.n8 VSUBS 0.009046f
C295 B.n9 VSUBS 0.009046f
C296 B.n10 VSUBS 0.009046f
C297 B.n11 VSUBS 0.009046f
C298 B.n12 VSUBS 0.009046f
C299 B.n13 VSUBS 0.009046f
C300 B.n14 VSUBS 0.009046f
C301 B.n15 VSUBS 0.019512f
C302 B.n16 VSUBS 0.009046f
C303 B.n17 VSUBS 0.009046f
C304 B.n18 VSUBS 0.009046f
C305 B.n19 VSUBS 0.009046f
C306 B.n20 VSUBS 0.009046f
C307 B.n21 VSUBS 0.009046f
C308 B.n22 VSUBS 0.009046f
C309 B.n23 VSUBS 0.009046f
C310 B.n24 VSUBS 0.009046f
C311 B.n25 VSUBS 0.009046f
C312 B.n26 VSUBS 0.009046f
C313 B.n27 VSUBS 0.009046f
C314 B.n28 VSUBS 0.009046f
C315 B.n29 VSUBS 0.009046f
C316 B.n30 VSUBS 0.009046f
C317 B.n31 VSUBS 0.009046f
C318 B.n32 VSUBS 0.009046f
C319 B.n33 VSUBS 0.009046f
C320 B.n34 VSUBS 0.009046f
C321 B.n35 VSUBS 0.009046f
C322 B.n36 VSUBS 0.009046f
C323 B.n37 VSUBS 0.009046f
C324 B.n38 VSUBS 0.009046f
C325 B.n39 VSUBS 0.009046f
C326 B.n40 VSUBS 0.009046f
C327 B.n41 VSUBS 0.009046f
C328 B.n42 VSUBS 0.009046f
C329 B.n43 VSUBS 0.009046f
C330 B.n44 VSUBS 0.009046f
C331 B.n45 VSUBS 0.009046f
C332 B.t11 VSUBS 0.463279f
C333 B.t10 VSUBS 0.479662f
C334 B.t9 VSUBS 0.696993f
C335 B.n46 VSUBS 0.578235f
C336 B.n47 VSUBS 0.419204f
C337 B.n48 VSUBS 0.009046f
C338 B.n49 VSUBS 0.009046f
C339 B.n50 VSUBS 0.009046f
C340 B.n51 VSUBS 0.009046f
C341 B.n52 VSUBS 0.005055f
C342 B.n53 VSUBS 0.009046f
C343 B.t8 VSUBS 0.463283f
C344 B.t7 VSUBS 0.479667f
C345 B.t6 VSUBS 0.696993f
C346 B.n54 VSUBS 0.578231f
C347 B.n55 VSUBS 0.419199f
C348 B.n56 VSUBS 0.020958f
C349 B.n57 VSUBS 0.009046f
C350 B.n58 VSUBS 0.009046f
C351 B.n59 VSUBS 0.009046f
C352 B.n60 VSUBS 0.009046f
C353 B.n61 VSUBS 0.009046f
C354 B.n62 VSUBS 0.009046f
C355 B.n63 VSUBS 0.009046f
C356 B.n64 VSUBS 0.009046f
C357 B.n65 VSUBS 0.009046f
C358 B.n66 VSUBS 0.009046f
C359 B.n67 VSUBS 0.009046f
C360 B.n68 VSUBS 0.009046f
C361 B.n69 VSUBS 0.009046f
C362 B.n70 VSUBS 0.009046f
C363 B.n71 VSUBS 0.009046f
C364 B.n72 VSUBS 0.009046f
C365 B.n73 VSUBS 0.009046f
C366 B.n74 VSUBS 0.009046f
C367 B.n75 VSUBS 0.009046f
C368 B.n76 VSUBS 0.009046f
C369 B.n77 VSUBS 0.009046f
C370 B.n78 VSUBS 0.009046f
C371 B.n79 VSUBS 0.009046f
C372 B.n80 VSUBS 0.009046f
C373 B.n81 VSUBS 0.009046f
C374 B.n82 VSUBS 0.009046f
C375 B.n83 VSUBS 0.009046f
C376 B.n84 VSUBS 0.009046f
C377 B.n85 VSUBS 0.019226f
C378 B.n86 VSUBS 0.009046f
C379 B.n87 VSUBS 0.009046f
C380 B.n88 VSUBS 0.009046f
C381 B.n89 VSUBS 0.009046f
C382 B.n90 VSUBS 0.009046f
C383 B.n91 VSUBS 0.009046f
C384 B.n92 VSUBS 0.009046f
C385 B.n93 VSUBS 0.009046f
C386 B.n94 VSUBS 0.009046f
C387 B.n95 VSUBS 0.009046f
C388 B.n96 VSUBS 0.009046f
C389 B.n97 VSUBS 0.009046f
C390 B.n98 VSUBS 0.009046f
C391 B.n99 VSUBS 0.009046f
C392 B.n100 VSUBS 0.009046f
C393 B.n101 VSUBS 0.009046f
C394 B.n102 VSUBS 0.009046f
C395 B.n103 VSUBS 0.009046f
C396 B.n104 VSUBS 0.009046f
C397 B.n105 VSUBS 0.009046f
C398 B.n106 VSUBS 0.009046f
C399 B.n107 VSUBS 0.009046f
C400 B.n108 VSUBS 0.009046f
C401 B.n109 VSUBS 0.009046f
C402 B.n110 VSUBS 0.009046f
C403 B.n111 VSUBS 0.009046f
C404 B.n112 VSUBS 0.009046f
C405 B.n113 VSUBS 0.020397f
C406 B.n114 VSUBS 0.009046f
C407 B.n115 VSUBS 0.009046f
C408 B.n116 VSUBS 0.009046f
C409 B.n117 VSUBS 0.009046f
C410 B.n118 VSUBS 0.009046f
C411 B.n119 VSUBS 0.009046f
C412 B.n120 VSUBS 0.009046f
C413 B.n121 VSUBS 0.009046f
C414 B.n122 VSUBS 0.009046f
C415 B.n123 VSUBS 0.009046f
C416 B.n124 VSUBS 0.009046f
C417 B.n125 VSUBS 0.009046f
C418 B.n126 VSUBS 0.009046f
C419 B.n127 VSUBS 0.009046f
C420 B.n128 VSUBS 0.009046f
C421 B.n129 VSUBS 0.009046f
C422 B.n130 VSUBS 0.009046f
C423 B.n131 VSUBS 0.009046f
C424 B.n132 VSUBS 0.009046f
C425 B.n133 VSUBS 0.009046f
C426 B.n134 VSUBS 0.009046f
C427 B.n135 VSUBS 0.009046f
C428 B.n136 VSUBS 0.009046f
C429 B.n137 VSUBS 0.009046f
C430 B.n138 VSUBS 0.009046f
C431 B.n139 VSUBS 0.009046f
C432 B.n140 VSUBS 0.009046f
C433 B.n141 VSUBS 0.009046f
C434 B.n142 VSUBS 0.009046f
C435 B.t4 VSUBS 0.463283f
C436 B.t5 VSUBS 0.479667f
C437 B.t3 VSUBS 0.696993f
C438 B.n143 VSUBS 0.578231f
C439 B.n144 VSUBS 0.419199f
C440 B.n145 VSUBS 0.020958f
C441 B.n146 VSUBS 0.009046f
C442 B.n147 VSUBS 0.009046f
C443 B.n148 VSUBS 0.009046f
C444 B.n149 VSUBS 0.009046f
C445 B.n150 VSUBS 0.009046f
C446 B.t1 VSUBS 0.463279f
C447 B.t2 VSUBS 0.479662f
C448 B.t0 VSUBS 0.696993f
C449 B.n151 VSUBS 0.578235f
C450 B.n152 VSUBS 0.419204f
C451 B.n153 VSUBS 0.009046f
C452 B.n154 VSUBS 0.009046f
C453 B.n155 VSUBS 0.009046f
C454 B.n156 VSUBS 0.009046f
C455 B.n157 VSUBS 0.009046f
C456 B.n158 VSUBS 0.009046f
C457 B.n159 VSUBS 0.009046f
C458 B.n160 VSUBS 0.009046f
C459 B.n161 VSUBS 0.009046f
C460 B.n162 VSUBS 0.009046f
C461 B.n163 VSUBS 0.009046f
C462 B.n164 VSUBS 0.009046f
C463 B.n165 VSUBS 0.009046f
C464 B.n166 VSUBS 0.009046f
C465 B.n167 VSUBS 0.009046f
C466 B.n168 VSUBS 0.009046f
C467 B.n169 VSUBS 0.009046f
C468 B.n170 VSUBS 0.009046f
C469 B.n171 VSUBS 0.009046f
C470 B.n172 VSUBS 0.009046f
C471 B.n173 VSUBS 0.009046f
C472 B.n174 VSUBS 0.009046f
C473 B.n175 VSUBS 0.009046f
C474 B.n176 VSUBS 0.009046f
C475 B.n177 VSUBS 0.009046f
C476 B.n178 VSUBS 0.009046f
C477 B.n179 VSUBS 0.009046f
C478 B.n180 VSUBS 0.009046f
C479 B.n181 VSUBS 0.009046f
C480 B.n182 VSUBS 0.020397f
C481 B.n183 VSUBS 0.009046f
C482 B.n184 VSUBS 0.009046f
C483 B.n185 VSUBS 0.009046f
C484 B.n186 VSUBS 0.009046f
C485 B.n187 VSUBS 0.009046f
C486 B.n188 VSUBS 0.009046f
C487 B.n189 VSUBS 0.009046f
C488 B.n190 VSUBS 0.009046f
C489 B.n191 VSUBS 0.009046f
C490 B.n192 VSUBS 0.009046f
C491 B.n193 VSUBS 0.009046f
C492 B.n194 VSUBS 0.009046f
C493 B.n195 VSUBS 0.009046f
C494 B.n196 VSUBS 0.009046f
C495 B.n197 VSUBS 0.009046f
C496 B.n198 VSUBS 0.009046f
C497 B.n199 VSUBS 0.009046f
C498 B.n200 VSUBS 0.009046f
C499 B.n201 VSUBS 0.009046f
C500 B.n202 VSUBS 0.009046f
C501 B.n203 VSUBS 0.009046f
C502 B.n204 VSUBS 0.009046f
C503 B.n205 VSUBS 0.009046f
C504 B.n206 VSUBS 0.009046f
C505 B.n207 VSUBS 0.009046f
C506 B.n208 VSUBS 0.009046f
C507 B.n209 VSUBS 0.009046f
C508 B.n210 VSUBS 0.009046f
C509 B.n211 VSUBS 0.009046f
C510 B.n212 VSUBS 0.009046f
C511 B.n213 VSUBS 0.009046f
C512 B.n214 VSUBS 0.009046f
C513 B.n215 VSUBS 0.009046f
C514 B.n216 VSUBS 0.009046f
C515 B.n217 VSUBS 0.009046f
C516 B.n218 VSUBS 0.009046f
C517 B.n219 VSUBS 0.009046f
C518 B.n220 VSUBS 0.009046f
C519 B.n221 VSUBS 0.009046f
C520 B.n222 VSUBS 0.009046f
C521 B.n223 VSUBS 0.009046f
C522 B.n224 VSUBS 0.009046f
C523 B.n225 VSUBS 0.009046f
C524 B.n226 VSUBS 0.009046f
C525 B.n227 VSUBS 0.009046f
C526 B.n228 VSUBS 0.009046f
C527 B.n229 VSUBS 0.009046f
C528 B.n230 VSUBS 0.009046f
C529 B.n231 VSUBS 0.009046f
C530 B.n232 VSUBS 0.009046f
C531 B.n233 VSUBS 0.019512f
C532 B.n234 VSUBS 0.019512f
C533 B.n235 VSUBS 0.020397f
C534 B.n236 VSUBS 0.009046f
C535 B.n237 VSUBS 0.009046f
C536 B.n238 VSUBS 0.009046f
C537 B.n239 VSUBS 0.009046f
C538 B.n240 VSUBS 0.009046f
C539 B.n241 VSUBS 0.009046f
C540 B.n242 VSUBS 0.009046f
C541 B.n243 VSUBS 0.009046f
C542 B.n244 VSUBS 0.009046f
C543 B.n245 VSUBS 0.009046f
C544 B.n246 VSUBS 0.009046f
C545 B.n247 VSUBS 0.009046f
C546 B.n248 VSUBS 0.009046f
C547 B.n249 VSUBS 0.009046f
C548 B.n250 VSUBS 0.009046f
C549 B.n251 VSUBS 0.009046f
C550 B.n252 VSUBS 0.009046f
C551 B.n253 VSUBS 0.009046f
C552 B.n254 VSUBS 0.009046f
C553 B.n255 VSUBS 0.009046f
C554 B.n256 VSUBS 0.009046f
C555 B.n257 VSUBS 0.009046f
C556 B.n258 VSUBS 0.009046f
C557 B.n259 VSUBS 0.009046f
C558 B.n260 VSUBS 0.009046f
C559 B.n261 VSUBS 0.009046f
C560 B.n262 VSUBS 0.009046f
C561 B.n263 VSUBS 0.009046f
C562 B.n264 VSUBS 0.009046f
C563 B.n265 VSUBS 0.009046f
C564 B.n266 VSUBS 0.009046f
C565 B.n267 VSUBS 0.009046f
C566 B.n268 VSUBS 0.009046f
C567 B.n269 VSUBS 0.009046f
C568 B.n270 VSUBS 0.009046f
C569 B.n271 VSUBS 0.009046f
C570 B.n272 VSUBS 0.009046f
C571 B.n273 VSUBS 0.009046f
C572 B.n274 VSUBS 0.009046f
C573 B.n275 VSUBS 0.009046f
C574 B.n276 VSUBS 0.009046f
C575 B.n277 VSUBS 0.009046f
C576 B.n278 VSUBS 0.009046f
C577 B.n279 VSUBS 0.009046f
C578 B.n280 VSUBS 0.009046f
C579 B.n281 VSUBS 0.009046f
C580 B.n282 VSUBS 0.009046f
C581 B.n283 VSUBS 0.009046f
C582 B.n284 VSUBS 0.009046f
C583 B.n285 VSUBS 0.009046f
C584 B.n286 VSUBS 0.009046f
C585 B.n287 VSUBS 0.009046f
C586 B.n288 VSUBS 0.009046f
C587 B.n289 VSUBS 0.009046f
C588 B.n290 VSUBS 0.009046f
C589 B.n291 VSUBS 0.009046f
C590 B.n292 VSUBS 0.009046f
C591 B.n293 VSUBS 0.009046f
C592 B.n294 VSUBS 0.009046f
C593 B.n295 VSUBS 0.009046f
C594 B.n296 VSUBS 0.009046f
C595 B.n297 VSUBS 0.009046f
C596 B.n298 VSUBS 0.009046f
C597 B.n299 VSUBS 0.009046f
C598 B.n300 VSUBS 0.009046f
C599 B.n301 VSUBS 0.009046f
C600 B.n302 VSUBS 0.009046f
C601 B.n303 VSUBS 0.009046f
C602 B.n304 VSUBS 0.009046f
C603 B.n305 VSUBS 0.009046f
C604 B.n306 VSUBS 0.009046f
C605 B.n307 VSUBS 0.009046f
C606 B.n308 VSUBS 0.009046f
C607 B.n309 VSUBS 0.009046f
C608 B.n310 VSUBS 0.009046f
C609 B.n311 VSUBS 0.009046f
C610 B.n312 VSUBS 0.009046f
C611 B.n313 VSUBS 0.009046f
C612 B.n314 VSUBS 0.009046f
C613 B.n315 VSUBS 0.009046f
C614 B.n316 VSUBS 0.009046f
C615 B.n317 VSUBS 0.009046f
C616 B.n318 VSUBS 0.009046f
C617 B.n319 VSUBS 0.009046f
C618 B.n320 VSUBS 0.009046f
C619 B.n321 VSUBS 0.009046f
C620 B.n322 VSUBS 0.009046f
C621 B.n323 VSUBS 0.009046f
C622 B.n324 VSUBS 0.008514f
C623 B.n325 VSUBS 0.020958f
C624 B.n326 VSUBS 0.005055f
C625 B.n327 VSUBS 0.009046f
C626 B.n328 VSUBS 0.009046f
C627 B.n329 VSUBS 0.009046f
C628 B.n330 VSUBS 0.009046f
C629 B.n331 VSUBS 0.009046f
C630 B.n332 VSUBS 0.009046f
C631 B.n333 VSUBS 0.009046f
C632 B.n334 VSUBS 0.009046f
C633 B.n335 VSUBS 0.009046f
C634 B.n336 VSUBS 0.009046f
C635 B.n337 VSUBS 0.009046f
C636 B.n338 VSUBS 0.009046f
C637 B.n339 VSUBS 0.005055f
C638 B.n340 VSUBS 0.009046f
C639 B.n341 VSUBS 0.009046f
C640 B.n342 VSUBS 0.008514f
C641 B.n343 VSUBS 0.009046f
C642 B.n344 VSUBS 0.009046f
C643 B.n345 VSUBS 0.009046f
C644 B.n346 VSUBS 0.009046f
C645 B.n347 VSUBS 0.009046f
C646 B.n348 VSUBS 0.009046f
C647 B.n349 VSUBS 0.009046f
C648 B.n350 VSUBS 0.009046f
C649 B.n351 VSUBS 0.009046f
C650 B.n352 VSUBS 0.009046f
C651 B.n353 VSUBS 0.009046f
C652 B.n354 VSUBS 0.009046f
C653 B.n355 VSUBS 0.009046f
C654 B.n356 VSUBS 0.009046f
C655 B.n357 VSUBS 0.009046f
C656 B.n358 VSUBS 0.009046f
C657 B.n359 VSUBS 0.009046f
C658 B.n360 VSUBS 0.009046f
C659 B.n361 VSUBS 0.009046f
C660 B.n362 VSUBS 0.009046f
C661 B.n363 VSUBS 0.009046f
C662 B.n364 VSUBS 0.009046f
C663 B.n365 VSUBS 0.009046f
C664 B.n366 VSUBS 0.009046f
C665 B.n367 VSUBS 0.009046f
C666 B.n368 VSUBS 0.009046f
C667 B.n369 VSUBS 0.009046f
C668 B.n370 VSUBS 0.009046f
C669 B.n371 VSUBS 0.009046f
C670 B.n372 VSUBS 0.009046f
C671 B.n373 VSUBS 0.009046f
C672 B.n374 VSUBS 0.009046f
C673 B.n375 VSUBS 0.009046f
C674 B.n376 VSUBS 0.009046f
C675 B.n377 VSUBS 0.009046f
C676 B.n378 VSUBS 0.009046f
C677 B.n379 VSUBS 0.009046f
C678 B.n380 VSUBS 0.009046f
C679 B.n381 VSUBS 0.009046f
C680 B.n382 VSUBS 0.009046f
C681 B.n383 VSUBS 0.009046f
C682 B.n384 VSUBS 0.009046f
C683 B.n385 VSUBS 0.009046f
C684 B.n386 VSUBS 0.009046f
C685 B.n387 VSUBS 0.009046f
C686 B.n388 VSUBS 0.009046f
C687 B.n389 VSUBS 0.009046f
C688 B.n390 VSUBS 0.009046f
C689 B.n391 VSUBS 0.009046f
C690 B.n392 VSUBS 0.009046f
C691 B.n393 VSUBS 0.009046f
C692 B.n394 VSUBS 0.009046f
C693 B.n395 VSUBS 0.009046f
C694 B.n396 VSUBS 0.009046f
C695 B.n397 VSUBS 0.009046f
C696 B.n398 VSUBS 0.009046f
C697 B.n399 VSUBS 0.009046f
C698 B.n400 VSUBS 0.009046f
C699 B.n401 VSUBS 0.009046f
C700 B.n402 VSUBS 0.009046f
C701 B.n403 VSUBS 0.009046f
C702 B.n404 VSUBS 0.009046f
C703 B.n405 VSUBS 0.009046f
C704 B.n406 VSUBS 0.009046f
C705 B.n407 VSUBS 0.009046f
C706 B.n408 VSUBS 0.009046f
C707 B.n409 VSUBS 0.009046f
C708 B.n410 VSUBS 0.009046f
C709 B.n411 VSUBS 0.009046f
C710 B.n412 VSUBS 0.009046f
C711 B.n413 VSUBS 0.009046f
C712 B.n414 VSUBS 0.009046f
C713 B.n415 VSUBS 0.009046f
C714 B.n416 VSUBS 0.009046f
C715 B.n417 VSUBS 0.009046f
C716 B.n418 VSUBS 0.009046f
C717 B.n419 VSUBS 0.009046f
C718 B.n420 VSUBS 0.009046f
C719 B.n421 VSUBS 0.009046f
C720 B.n422 VSUBS 0.009046f
C721 B.n423 VSUBS 0.009046f
C722 B.n424 VSUBS 0.009046f
C723 B.n425 VSUBS 0.009046f
C724 B.n426 VSUBS 0.009046f
C725 B.n427 VSUBS 0.009046f
C726 B.n428 VSUBS 0.009046f
C727 B.n429 VSUBS 0.009046f
C728 B.n430 VSUBS 0.020397f
C729 B.n431 VSUBS 0.019512f
C730 B.n432 VSUBS 0.019512f
C731 B.n433 VSUBS 0.009046f
C732 B.n434 VSUBS 0.009046f
C733 B.n435 VSUBS 0.009046f
C734 B.n436 VSUBS 0.009046f
C735 B.n437 VSUBS 0.009046f
C736 B.n438 VSUBS 0.009046f
C737 B.n439 VSUBS 0.009046f
C738 B.n440 VSUBS 0.009046f
C739 B.n441 VSUBS 0.009046f
C740 B.n442 VSUBS 0.009046f
C741 B.n443 VSUBS 0.009046f
C742 B.n444 VSUBS 0.009046f
C743 B.n445 VSUBS 0.009046f
C744 B.n446 VSUBS 0.009046f
C745 B.n447 VSUBS 0.009046f
C746 B.n448 VSUBS 0.009046f
C747 B.n449 VSUBS 0.009046f
C748 B.n450 VSUBS 0.009046f
C749 B.n451 VSUBS 0.009046f
C750 B.n452 VSUBS 0.009046f
C751 B.n453 VSUBS 0.009046f
C752 B.n454 VSUBS 0.009046f
C753 B.n455 VSUBS 0.009046f
C754 B.n456 VSUBS 0.009046f
C755 B.n457 VSUBS 0.009046f
C756 B.n458 VSUBS 0.009046f
C757 B.n459 VSUBS 0.009046f
C758 B.n460 VSUBS 0.009046f
C759 B.n461 VSUBS 0.009046f
C760 B.n462 VSUBS 0.009046f
C761 B.n463 VSUBS 0.009046f
C762 B.n464 VSUBS 0.009046f
C763 B.n465 VSUBS 0.009046f
C764 B.n466 VSUBS 0.009046f
C765 B.n467 VSUBS 0.009046f
C766 B.n468 VSUBS 0.009046f
C767 B.n469 VSUBS 0.009046f
C768 B.n470 VSUBS 0.009046f
C769 B.n471 VSUBS 0.009046f
C770 B.n472 VSUBS 0.009046f
C771 B.n473 VSUBS 0.009046f
C772 B.n474 VSUBS 0.009046f
C773 B.n475 VSUBS 0.009046f
C774 B.n476 VSUBS 0.009046f
C775 B.n477 VSUBS 0.009046f
C776 B.n478 VSUBS 0.009046f
C777 B.n479 VSUBS 0.009046f
C778 B.n480 VSUBS 0.009046f
C779 B.n481 VSUBS 0.009046f
C780 B.n482 VSUBS 0.009046f
C781 B.n483 VSUBS 0.009046f
C782 B.n484 VSUBS 0.009046f
C783 B.n485 VSUBS 0.009046f
C784 B.n486 VSUBS 0.009046f
C785 B.n487 VSUBS 0.009046f
C786 B.n488 VSUBS 0.009046f
C787 B.n489 VSUBS 0.009046f
C788 B.n490 VSUBS 0.009046f
C789 B.n491 VSUBS 0.009046f
C790 B.n492 VSUBS 0.009046f
C791 B.n493 VSUBS 0.009046f
C792 B.n494 VSUBS 0.009046f
C793 B.n495 VSUBS 0.009046f
C794 B.n496 VSUBS 0.009046f
C795 B.n497 VSUBS 0.009046f
C796 B.n498 VSUBS 0.009046f
C797 B.n499 VSUBS 0.009046f
C798 B.n500 VSUBS 0.009046f
C799 B.n501 VSUBS 0.009046f
C800 B.n502 VSUBS 0.009046f
C801 B.n503 VSUBS 0.009046f
C802 B.n504 VSUBS 0.009046f
C803 B.n505 VSUBS 0.009046f
C804 B.n506 VSUBS 0.009046f
C805 B.n507 VSUBS 0.009046f
C806 B.n508 VSUBS 0.009046f
C807 B.n509 VSUBS 0.009046f
C808 B.n510 VSUBS 0.009046f
C809 B.n511 VSUBS 0.009046f
C810 B.n512 VSUBS 0.020683f
C811 B.n513 VSUBS 0.019512f
C812 B.n514 VSUBS 0.020397f
C813 B.n515 VSUBS 0.009046f
C814 B.n516 VSUBS 0.009046f
C815 B.n517 VSUBS 0.009046f
C816 B.n518 VSUBS 0.009046f
C817 B.n519 VSUBS 0.009046f
C818 B.n520 VSUBS 0.009046f
C819 B.n521 VSUBS 0.009046f
C820 B.n522 VSUBS 0.009046f
C821 B.n523 VSUBS 0.009046f
C822 B.n524 VSUBS 0.009046f
C823 B.n525 VSUBS 0.009046f
C824 B.n526 VSUBS 0.009046f
C825 B.n527 VSUBS 0.009046f
C826 B.n528 VSUBS 0.009046f
C827 B.n529 VSUBS 0.009046f
C828 B.n530 VSUBS 0.009046f
C829 B.n531 VSUBS 0.009046f
C830 B.n532 VSUBS 0.009046f
C831 B.n533 VSUBS 0.009046f
C832 B.n534 VSUBS 0.009046f
C833 B.n535 VSUBS 0.009046f
C834 B.n536 VSUBS 0.009046f
C835 B.n537 VSUBS 0.009046f
C836 B.n538 VSUBS 0.009046f
C837 B.n539 VSUBS 0.009046f
C838 B.n540 VSUBS 0.009046f
C839 B.n541 VSUBS 0.009046f
C840 B.n542 VSUBS 0.009046f
C841 B.n543 VSUBS 0.009046f
C842 B.n544 VSUBS 0.009046f
C843 B.n545 VSUBS 0.009046f
C844 B.n546 VSUBS 0.009046f
C845 B.n547 VSUBS 0.009046f
C846 B.n548 VSUBS 0.009046f
C847 B.n549 VSUBS 0.009046f
C848 B.n550 VSUBS 0.009046f
C849 B.n551 VSUBS 0.009046f
C850 B.n552 VSUBS 0.009046f
C851 B.n553 VSUBS 0.009046f
C852 B.n554 VSUBS 0.009046f
C853 B.n555 VSUBS 0.009046f
C854 B.n556 VSUBS 0.009046f
C855 B.n557 VSUBS 0.009046f
C856 B.n558 VSUBS 0.009046f
C857 B.n559 VSUBS 0.009046f
C858 B.n560 VSUBS 0.009046f
C859 B.n561 VSUBS 0.009046f
C860 B.n562 VSUBS 0.009046f
C861 B.n563 VSUBS 0.009046f
C862 B.n564 VSUBS 0.009046f
C863 B.n565 VSUBS 0.009046f
C864 B.n566 VSUBS 0.009046f
C865 B.n567 VSUBS 0.009046f
C866 B.n568 VSUBS 0.009046f
C867 B.n569 VSUBS 0.009046f
C868 B.n570 VSUBS 0.009046f
C869 B.n571 VSUBS 0.009046f
C870 B.n572 VSUBS 0.009046f
C871 B.n573 VSUBS 0.009046f
C872 B.n574 VSUBS 0.009046f
C873 B.n575 VSUBS 0.009046f
C874 B.n576 VSUBS 0.009046f
C875 B.n577 VSUBS 0.009046f
C876 B.n578 VSUBS 0.009046f
C877 B.n579 VSUBS 0.009046f
C878 B.n580 VSUBS 0.009046f
C879 B.n581 VSUBS 0.009046f
C880 B.n582 VSUBS 0.009046f
C881 B.n583 VSUBS 0.009046f
C882 B.n584 VSUBS 0.009046f
C883 B.n585 VSUBS 0.009046f
C884 B.n586 VSUBS 0.009046f
C885 B.n587 VSUBS 0.009046f
C886 B.n588 VSUBS 0.009046f
C887 B.n589 VSUBS 0.009046f
C888 B.n590 VSUBS 0.009046f
C889 B.n591 VSUBS 0.009046f
C890 B.n592 VSUBS 0.009046f
C891 B.n593 VSUBS 0.009046f
C892 B.n594 VSUBS 0.009046f
C893 B.n595 VSUBS 0.009046f
C894 B.n596 VSUBS 0.009046f
C895 B.n597 VSUBS 0.009046f
C896 B.n598 VSUBS 0.009046f
C897 B.n599 VSUBS 0.009046f
C898 B.n600 VSUBS 0.009046f
C899 B.n601 VSUBS 0.009046f
C900 B.n602 VSUBS 0.008514f
C901 B.n603 VSUBS 0.009046f
C902 B.n604 VSUBS 0.009046f
C903 B.n605 VSUBS 0.009046f
C904 B.n606 VSUBS 0.009046f
C905 B.n607 VSUBS 0.009046f
C906 B.n608 VSUBS 0.009046f
C907 B.n609 VSUBS 0.009046f
C908 B.n610 VSUBS 0.009046f
C909 B.n611 VSUBS 0.009046f
C910 B.n612 VSUBS 0.009046f
C911 B.n613 VSUBS 0.009046f
C912 B.n614 VSUBS 0.009046f
C913 B.n615 VSUBS 0.009046f
C914 B.n616 VSUBS 0.009046f
C915 B.n617 VSUBS 0.009046f
C916 B.n618 VSUBS 0.005055f
C917 B.n619 VSUBS 0.020958f
C918 B.n620 VSUBS 0.008514f
C919 B.n621 VSUBS 0.009046f
C920 B.n622 VSUBS 0.009046f
C921 B.n623 VSUBS 0.009046f
C922 B.n624 VSUBS 0.009046f
C923 B.n625 VSUBS 0.009046f
C924 B.n626 VSUBS 0.009046f
C925 B.n627 VSUBS 0.009046f
C926 B.n628 VSUBS 0.009046f
C927 B.n629 VSUBS 0.009046f
C928 B.n630 VSUBS 0.009046f
C929 B.n631 VSUBS 0.009046f
C930 B.n632 VSUBS 0.009046f
C931 B.n633 VSUBS 0.009046f
C932 B.n634 VSUBS 0.009046f
C933 B.n635 VSUBS 0.009046f
C934 B.n636 VSUBS 0.009046f
C935 B.n637 VSUBS 0.009046f
C936 B.n638 VSUBS 0.009046f
C937 B.n639 VSUBS 0.009046f
C938 B.n640 VSUBS 0.009046f
C939 B.n641 VSUBS 0.009046f
C940 B.n642 VSUBS 0.009046f
C941 B.n643 VSUBS 0.009046f
C942 B.n644 VSUBS 0.009046f
C943 B.n645 VSUBS 0.009046f
C944 B.n646 VSUBS 0.009046f
C945 B.n647 VSUBS 0.009046f
C946 B.n648 VSUBS 0.009046f
C947 B.n649 VSUBS 0.009046f
C948 B.n650 VSUBS 0.009046f
C949 B.n651 VSUBS 0.009046f
C950 B.n652 VSUBS 0.009046f
C951 B.n653 VSUBS 0.009046f
C952 B.n654 VSUBS 0.009046f
C953 B.n655 VSUBS 0.009046f
C954 B.n656 VSUBS 0.009046f
C955 B.n657 VSUBS 0.009046f
C956 B.n658 VSUBS 0.009046f
C957 B.n659 VSUBS 0.009046f
C958 B.n660 VSUBS 0.009046f
C959 B.n661 VSUBS 0.009046f
C960 B.n662 VSUBS 0.009046f
C961 B.n663 VSUBS 0.009046f
C962 B.n664 VSUBS 0.009046f
C963 B.n665 VSUBS 0.009046f
C964 B.n666 VSUBS 0.009046f
C965 B.n667 VSUBS 0.009046f
C966 B.n668 VSUBS 0.009046f
C967 B.n669 VSUBS 0.009046f
C968 B.n670 VSUBS 0.009046f
C969 B.n671 VSUBS 0.009046f
C970 B.n672 VSUBS 0.009046f
C971 B.n673 VSUBS 0.009046f
C972 B.n674 VSUBS 0.009046f
C973 B.n675 VSUBS 0.009046f
C974 B.n676 VSUBS 0.009046f
C975 B.n677 VSUBS 0.009046f
C976 B.n678 VSUBS 0.009046f
C977 B.n679 VSUBS 0.009046f
C978 B.n680 VSUBS 0.009046f
C979 B.n681 VSUBS 0.009046f
C980 B.n682 VSUBS 0.009046f
C981 B.n683 VSUBS 0.009046f
C982 B.n684 VSUBS 0.009046f
C983 B.n685 VSUBS 0.009046f
C984 B.n686 VSUBS 0.009046f
C985 B.n687 VSUBS 0.009046f
C986 B.n688 VSUBS 0.009046f
C987 B.n689 VSUBS 0.009046f
C988 B.n690 VSUBS 0.009046f
C989 B.n691 VSUBS 0.009046f
C990 B.n692 VSUBS 0.009046f
C991 B.n693 VSUBS 0.009046f
C992 B.n694 VSUBS 0.009046f
C993 B.n695 VSUBS 0.009046f
C994 B.n696 VSUBS 0.009046f
C995 B.n697 VSUBS 0.009046f
C996 B.n698 VSUBS 0.009046f
C997 B.n699 VSUBS 0.009046f
C998 B.n700 VSUBS 0.009046f
C999 B.n701 VSUBS 0.009046f
C1000 B.n702 VSUBS 0.009046f
C1001 B.n703 VSUBS 0.009046f
C1002 B.n704 VSUBS 0.009046f
C1003 B.n705 VSUBS 0.009046f
C1004 B.n706 VSUBS 0.009046f
C1005 B.n707 VSUBS 0.009046f
C1006 B.n708 VSUBS 0.020397f
C1007 B.n709 VSUBS 0.020397f
C1008 B.n710 VSUBS 0.019512f
C1009 B.n711 VSUBS 0.009046f
C1010 B.n712 VSUBS 0.009046f
C1011 B.n713 VSUBS 0.009046f
C1012 B.n714 VSUBS 0.009046f
C1013 B.n715 VSUBS 0.009046f
C1014 B.n716 VSUBS 0.009046f
C1015 B.n717 VSUBS 0.009046f
C1016 B.n718 VSUBS 0.009046f
C1017 B.n719 VSUBS 0.009046f
C1018 B.n720 VSUBS 0.009046f
C1019 B.n721 VSUBS 0.009046f
C1020 B.n722 VSUBS 0.009046f
C1021 B.n723 VSUBS 0.009046f
C1022 B.n724 VSUBS 0.009046f
C1023 B.n725 VSUBS 0.009046f
C1024 B.n726 VSUBS 0.009046f
C1025 B.n727 VSUBS 0.009046f
C1026 B.n728 VSUBS 0.009046f
C1027 B.n729 VSUBS 0.009046f
C1028 B.n730 VSUBS 0.009046f
C1029 B.n731 VSUBS 0.009046f
C1030 B.n732 VSUBS 0.009046f
C1031 B.n733 VSUBS 0.009046f
C1032 B.n734 VSUBS 0.009046f
C1033 B.n735 VSUBS 0.009046f
C1034 B.n736 VSUBS 0.009046f
C1035 B.n737 VSUBS 0.009046f
C1036 B.n738 VSUBS 0.009046f
C1037 B.n739 VSUBS 0.009046f
C1038 B.n740 VSUBS 0.009046f
C1039 B.n741 VSUBS 0.009046f
C1040 B.n742 VSUBS 0.009046f
C1041 B.n743 VSUBS 0.009046f
C1042 B.n744 VSUBS 0.009046f
C1043 B.n745 VSUBS 0.009046f
C1044 B.n746 VSUBS 0.009046f
C1045 B.n747 VSUBS 0.009046f
C1046 B.n748 VSUBS 0.009046f
C1047 B.n749 VSUBS 0.009046f
C1048 B.n750 VSUBS 0.009046f
C1049 B.n751 VSUBS 0.020483f
C1050 VDD1.n0 VSUBS 0.031434f
C1051 VDD1.n1 VSUBS 0.028065f
C1052 VDD1.n2 VSUBS 0.015081f
C1053 VDD1.n3 VSUBS 0.035646f
C1054 VDD1.n4 VSUBS 0.015968f
C1055 VDD1.n5 VSUBS 0.028065f
C1056 VDD1.n6 VSUBS 0.015081f
C1057 VDD1.n7 VSUBS 0.035646f
C1058 VDD1.n8 VSUBS 0.015968f
C1059 VDD1.n9 VSUBS 0.028065f
C1060 VDD1.n10 VSUBS 0.015525f
C1061 VDD1.n11 VSUBS 0.035646f
C1062 VDD1.n12 VSUBS 0.015081f
C1063 VDD1.n13 VSUBS 0.015968f
C1064 VDD1.n14 VSUBS 0.028065f
C1065 VDD1.n15 VSUBS 0.015081f
C1066 VDD1.n16 VSUBS 0.035646f
C1067 VDD1.n17 VSUBS 0.015968f
C1068 VDD1.n18 VSUBS 0.028065f
C1069 VDD1.n19 VSUBS 0.015081f
C1070 VDD1.n20 VSUBS 0.035646f
C1071 VDD1.n21 VSUBS 0.015968f
C1072 VDD1.n22 VSUBS 0.028065f
C1073 VDD1.n23 VSUBS 0.015081f
C1074 VDD1.n24 VSUBS 0.035646f
C1075 VDD1.n25 VSUBS 0.015968f
C1076 VDD1.n26 VSUBS 0.028065f
C1077 VDD1.n27 VSUBS 0.015081f
C1078 VDD1.n28 VSUBS 0.035646f
C1079 VDD1.n29 VSUBS 0.015968f
C1080 VDD1.n30 VSUBS 0.028065f
C1081 VDD1.n31 VSUBS 0.015081f
C1082 VDD1.n32 VSUBS 0.026735f
C1083 VDD1.n33 VSUBS 0.022676f
C1084 VDD1.t9 VSUBS 0.076541f
C1085 VDD1.n34 VSUBS 0.225153f
C1086 VDD1.n35 VSUBS 2.21247f
C1087 VDD1.n36 VSUBS 0.015081f
C1088 VDD1.n37 VSUBS 0.015968f
C1089 VDD1.n38 VSUBS 0.035646f
C1090 VDD1.n39 VSUBS 0.035646f
C1091 VDD1.n40 VSUBS 0.015968f
C1092 VDD1.n41 VSUBS 0.015081f
C1093 VDD1.n42 VSUBS 0.028065f
C1094 VDD1.n43 VSUBS 0.028065f
C1095 VDD1.n44 VSUBS 0.015081f
C1096 VDD1.n45 VSUBS 0.015968f
C1097 VDD1.n46 VSUBS 0.035646f
C1098 VDD1.n47 VSUBS 0.035646f
C1099 VDD1.n48 VSUBS 0.015968f
C1100 VDD1.n49 VSUBS 0.015081f
C1101 VDD1.n50 VSUBS 0.028065f
C1102 VDD1.n51 VSUBS 0.028065f
C1103 VDD1.n52 VSUBS 0.015081f
C1104 VDD1.n53 VSUBS 0.015968f
C1105 VDD1.n54 VSUBS 0.035646f
C1106 VDD1.n55 VSUBS 0.035646f
C1107 VDD1.n56 VSUBS 0.015968f
C1108 VDD1.n57 VSUBS 0.015081f
C1109 VDD1.n58 VSUBS 0.028065f
C1110 VDD1.n59 VSUBS 0.028065f
C1111 VDD1.n60 VSUBS 0.015081f
C1112 VDD1.n61 VSUBS 0.015968f
C1113 VDD1.n62 VSUBS 0.035646f
C1114 VDD1.n63 VSUBS 0.035646f
C1115 VDD1.n64 VSUBS 0.015968f
C1116 VDD1.n65 VSUBS 0.015081f
C1117 VDD1.n66 VSUBS 0.028065f
C1118 VDD1.n67 VSUBS 0.028065f
C1119 VDD1.n68 VSUBS 0.015081f
C1120 VDD1.n69 VSUBS 0.015968f
C1121 VDD1.n70 VSUBS 0.035646f
C1122 VDD1.n71 VSUBS 0.035646f
C1123 VDD1.n72 VSUBS 0.015968f
C1124 VDD1.n73 VSUBS 0.015081f
C1125 VDD1.n74 VSUBS 0.028065f
C1126 VDD1.n75 VSUBS 0.028065f
C1127 VDD1.n76 VSUBS 0.015081f
C1128 VDD1.n77 VSUBS 0.015968f
C1129 VDD1.n78 VSUBS 0.035646f
C1130 VDD1.n79 VSUBS 0.035646f
C1131 VDD1.n80 VSUBS 0.035646f
C1132 VDD1.n81 VSUBS 0.015525f
C1133 VDD1.n82 VSUBS 0.015081f
C1134 VDD1.n83 VSUBS 0.028065f
C1135 VDD1.n84 VSUBS 0.028065f
C1136 VDD1.n85 VSUBS 0.015081f
C1137 VDD1.n86 VSUBS 0.015968f
C1138 VDD1.n87 VSUBS 0.035646f
C1139 VDD1.n88 VSUBS 0.035646f
C1140 VDD1.n89 VSUBS 0.015968f
C1141 VDD1.n90 VSUBS 0.015081f
C1142 VDD1.n91 VSUBS 0.028065f
C1143 VDD1.n92 VSUBS 0.028065f
C1144 VDD1.n93 VSUBS 0.015081f
C1145 VDD1.n94 VSUBS 0.015968f
C1146 VDD1.n95 VSUBS 0.035646f
C1147 VDD1.n96 VSUBS 0.088327f
C1148 VDD1.n97 VSUBS 0.015968f
C1149 VDD1.n98 VSUBS 0.015081f
C1150 VDD1.n99 VSUBS 0.067172f
C1151 VDD1.n100 VSUBS 0.066415f
C1152 VDD1.t6 VSUBS 0.405857f
C1153 VDD1.t7 VSUBS 0.405857f
C1154 VDD1.n101 VSUBS 3.38332f
C1155 VDD1.n102 VSUBS 0.79396f
C1156 VDD1.n103 VSUBS 0.031434f
C1157 VDD1.n104 VSUBS 0.028065f
C1158 VDD1.n105 VSUBS 0.015081f
C1159 VDD1.n106 VSUBS 0.035646f
C1160 VDD1.n107 VSUBS 0.015968f
C1161 VDD1.n108 VSUBS 0.028065f
C1162 VDD1.n109 VSUBS 0.015081f
C1163 VDD1.n110 VSUBS 0.035646f
C1164 VDD1.n111 VSUBS 0.015968f
C1165 VDD1.n112 VSUBS 0.028065f
C1166 VDD1.n113 VSUBS 0.015525f
C1167 VDD1.n114 VSUBS 0.035646f
C1168 VDD1.n115 VSUBS 0.015968f
C1169 VDD1.n116 VSUBS 0.028065f
C1170 VDD1.n117 VSUBS 0.015081f
C1171 VDD1.n118 VSUBS 0.035646f
C1172 VDD1.n119 VSUBS 0.015968f
C1173 VDD1.n120 VSUBS 0.028065f
C1174 VDD1.n121 VSUBS 0.015081f
C1175 VDD1.n122 VSUBS 0.035646f
C1176 VDD1.n123 VSUBS 0.015968f
C1177 VDD1.n124 VSUBS 0.028065f
C1178 VDD1.n125 VSUBS 0.015081f
C1179 VDD1.n126 VSUBS 0.035646f
C1180 VDD1.n127 VSUBS 0.015968f
C1181 VDD1.n128 VSUBS 0.028065f
C1182 VDD1.n129 VSUBS 0.015081f
C1183 VDD1.n130 VSUBS 0.035646f
C1184 VDD1.n131 VSUBS 0.015968f
C1185 VDD1.n132 VSUBS 0.028065f
C1186 VDD1.n133 VSUBS 0.015081f
C1187 VDD1.n134 VSUBS 0.026735f
C1188 VDD1.n135 VSUBS 0.022676f
C1189 VDD1.t5 VSUBS 0.076541f
C1190 VDD1.n136 VSUBS 0.225153f
C1191 VDD1.n137 VSUBS 2.21247f
C1192 VDD1.n138 VSUBS 0.015081f
C1193 VDD1.n139 VSUBS 0.015968f
C1194 VDD1.n140 VSUBS 0.035646f
C1195 VDD1.n141 VSUBS 0.035646f
C1196 VDD1.n142 VSUBS 0.015968f
C1197 VDD1.n143 VSUBS 0.015081f
C1198 VDD1.n144 VSUBS 0.028065f
C1199 VDD1.n145 VSUBS 0.028065f
C1200 VDD1.n146 VSUBS 0.015081f
C1201 VDD1.n147 VSUBS 0.015968f
C1202 VDD1.n148 VSUBS 0.035646f
C1203 VDD1.n149 VSUBS 0.035646f
C1204 VDD1.n150 VSUBS 0.015968f
C1205 VDD1.n151 VSUBS 0.015081f
C1206 VDD1.n152 VSUBS 0.028065f
C1207 VDD1.n153 VSUBS 0.028065f
C1208 VDD1.n154 VSUBS 0.015081f
C1209 VDD1.n155 VSUBS 0.015968f
C1210 VDD1.n156 VSUBS 0.035646f
C1211 VDD1.n157 VSUBS 0.035646f
C1212 VDD1.n158 VSUBS 0.015968f
C1213 VDD1.n159 VSUBS 0.015081f
C1214 VDD1.n160 VSUBS 0.028065f
C1215 VDD1.n161 VSUBS 0.028065f
C1216 VDD1.n162 VSUBS 0.015081f
C1217 VDD1.n163 VSUBS 0.015968f
C1218 VDD1.n164 VSUBS 0.035646f
C1219 VDD1.n165 VSUBS 0.035646f
C1220 VDD1.n166 VSUBS 0.015968f
C1221 VDD1.n167 VSUBS 0.015081f
C1222 VDD1.n168 VSUBS 0.028065f
C1223 VDD1.n169 VSUBS 0.028065f
C1224 VDD1.n170 VSUBS 0.015081f
C1225 VDD1.n171 VSUBS 0.015968f
C1226 VDD1.n172 VSUBS 0.035646f
C1227 VDD1.n173 VSUBS 0.035646f
C1228 VDD1.n174 VSUBS 0.015968f
C1229 VDD1.n175 VSUBS 0.015081f
C1230 VDD1.n176 VSUBS 0.028065f
C1231 VDD1.n177 VSUBS 0.028065f
C1232 VDD1.n178 VSUBS 0.015081f
C1233 VDD1.n179 VSUBS 0.015081f
C1234 VDD1.n180 VSUBS 0.015968f
C1235 VDD1.n181 VSUBS 0.035646f
C1236 VDD1.n182 VSUBS 0.035646f
C1237 VDD1.n183 VSUBS 0.035646f
C1238 VDD1.n184 VSUBS 0.015525f
C1239 VDD1.n185 VSUBS 0.015081f
C1240 VDD1.n186 VSUBS 0.028065f
C1241 VDD1.n187 VSUBS 0.028065f
C1242 VDD1.n188 VSUBS 0.015081f
C1243 VDD1.n189 VSUBS 0.015968f
C1244 VDD1.n190 VSUBS 0.035646f
C1245 VDD1.n191 VSUBS 0.035646f
C1246 VDD1.n192 VSUBS 0.015968f
C1247 VDD1.n193 VSUBS 0.015081f
C1248 VDD1.n194 VSUBS 0.028065f
C1249 VDD1.n195 VSUBS 0.028065f
C1250 VDD1.n196 VSUBS 0.015081f
C1251 VDD1.n197 VSUBS 0.015968f
C1252 VDD1.n198 VSUBS 0.035646f
C1253 VDD1.n199 VSUBS 0.088327f
C1254 VDD1.n200 VSUBS 0.015968f
C1255 VDD1.n201 VSUBS 0.015081f
C1256 VDD1.n202 VSUBS 0.067172f
C1257 VDD1.n203 VSUBS 0.066415f
C1258 VDD1.t3 VSUBS 0.405857f
C1259 VDD1.t1 VSUBS 0.405857f
C1260 VDD1.n204 VSUBS 3.3833f
C1261 VDD1.n205 VSUBS 0.787466f
C1262 VDD1.t2 VSUBS 0.405857f
C1263 VDD1.t0 VSUBS 0.405857f
C1264 VDD1.n206 VSUBS 3.38958f
C1265 VDD1.n207 VSUBS 2.99805f
C1266 VDD1.t4 VSUBS 0.405857f
C1267 VDD1.t8 VSUBS 0.405857f
C1268 VDD1.n208 VSUBS 3.38331f
C1269 VDD1.n209 VSUBS 3.55452f
C1270 VTAIL.t0 VSUBS 0.407996f
C1271 VTAIL.t1 VSUBS 0.407996f
C1272 VTAIL.n0 VSUBS 3.22942f
C1273 VTAIL.n1 VSUBS 0.838002f
C1274 VTAIL.n2 VSUBS 0.0316f
C1275 VTAIL.n3 VSUBS 0.028213f
C1276 VTAIL.n4 VSUBS 0.015161f
C1277 VTAIL.n5 VSUBS 0.035834f
C1278 VTAIL.n6 VSUBS 0.016052f
C1279 VTAIL.n7 VSUBS 0.028213f
C1280 VTAIL.n8 VSUBS 0.015161f
C1281 VTAIL.n9 VSUBS 0.035834f
C1282 VTAIL.n10 VSUBS 0.016052f
C1283 VTAIL.n11 VSUBS 0.028213f
C1284 VTAIL.n12 VSUBS 0.015606f
C1285 VTAIL.n13 VSUBS 0.035834f
C1286 VTAIL.n14 VSUBS 0.016052f
C1287 VTAIL.n15 VSUBS 0.028213f
C1288 VTAIL.n16 VSUBS 0.015161f
C1289 VTAIL.n17 VSUBS 0.035834f
C1290 VTAIL.n18 VSUBS 0.016052f
C1291 VTAIL.n19 VSUBS 0.028213f
C1292 VTAIL.n20 VSUBS 0.015161f
C1293 VTAIL.n21 VSUBS 0.035834f
C1294 VTAIL.n22 VSUBS 0.016052f
C1295 VTAIL.n23 VSUBS 0.028213f
C1296 VTAIL.n24 VSUBS 0.015161f
C1297 VTAIL.n25 VSUBS 0.035834f
C1298 VTAIL.n26 VSUBS 0.016052f
C1299 VTAIL.n27 VSUBS 0.028213f
C1300 VTAIL.n28 VSUBS 0.015161f
C1301 VTAIL.n29 VSUBS 0.035834f
C1302 VTAIL.n30 VSUBS 0.016052f
C1303 VTAIL.n31 VSUBS 0.028213f
C1304 VTAIL.n32 VSUBS 0.015161f
C1305 VTAIL.n33 VSUBS 0.026875f
C1306 VTAIL.n34 VSUBS 0.022796f
C1307 VTAIL.t9 VSUBS 0.076945f
C1308 VTAIL.n35 VSUBS 0.226339f
C1309 VTAIL.n36 VSUBS 2.22413f
C1310 VTAIL.n37 VSUBS 0.015161f
C1311 VTAIL.n38 VSUBS 0.016052f
C1312 VTAIL.n39 VSUBS 0.035834f
C1313 VTAIL.n40 VSUBS 0.035834f
C1314 VTAIL.n41 VSUBS 0.016052f
C1315 VTAIL.n42 VSUBS 0.015161f
C1316 VTAIL.n43 VSUBS 0.028213f
C1317 VTAIL.n44 VSUBS 0.028213f
C1318 VTAIL.n45 VSUBS 0.015161f
C1319 VTAIL.n46 VSUBS 0.016052f
C1320 VTAIL.n47 VSUBS 0.035834f
C1321 VTAIL.n48 VSUBS 0.035834f
C1322 VTAIL.n49 VSUBS 0.016052f
C1323 VTAIL.n50 VSUBS 0.015161f
C1324 VTAIL.n51 VSUBS 0.028213f
C1325 VTAIL.n52 VSUBS 0.028213f
C1326 VTAIL.n53 VSUBS 0.015161f
C1327 VTAIL.n54 VSUBS 0.016052f
C1328 VTAIL.n55 VSUBS 0.035834f
C1329 VTAIL.n56 VSUBS 0.035834f
C1330 VTAIL.n57 VSUBS 0.016052f
C1331 VTAIL.n58 VSUBS 0.015161f
C1332 VTAIL.n59 VSUBS 0.028213f
C1333 VTAIL.n60 VSUBS 0.028213f
C1334 VTAIL.n61 VSUBS 0.015161f
C1335 VTAIL.n62 VSUBS 0.016052f
C1336 VTAIL.n63 VSUBS 0.035834f
C1337 VTAIL.n64 VSUBS 0.035834f
C1338 VTAIL.n65 VSUBS 0.016052f
C1339 VTAIL.n66 VSUBS 0.015161f
C1340 VTAIL.n67 VSUBS 0.028213f
C1341 VTAIL.n68 VSUBS 0.028213f
C1342 VTAIL.n69 VSUBS 0.015161f
C1343 VTAIL.n70 VSUBS 0.016052f
C1344 VTAIL.n71 VSUBS 0.035834f
C1345 VTAIL.n72 VSUBS 0.035834f
C1346 VTAIL.n73 VSUBS 0.016052f
C1347 VTAIL.n74 VSUBS 0.015161f
C1348 VTAIL.n75 VSUBS 0.028213f
C1349 VTAIL.n76 VSUBS 0.028213f
C1350 VTAIL.n77 VSUBS 0.015161f
C1351 VTAIL.n78 VSUBS 0.015161f
C1352 VTAIL.n79 VSUBS 0.016052f
C1353 VTAIL.n80 VSUBS 0.035834f
C1354 VTAIL.n81 VSUBS 0.035834f
C1355 VTAIL.n82 VSUBS 0.035834f
C1356 VTAIL.n83 VSUBS 0.015606f
C1357 VTAIL.n84 VSUBS 0.015161f
C1358 VTAIL.n85 VSUBS 0.028213f
C1359 VTAIL.n86 VSUBS 0.028213f
C1360 VTAIL.n87 VSUBS 0.015161f
C1361 VTAIL.n88 VSUBS 0.016052f
C1362 VTAIL.n89 VSUBS 0.035834f
C1363 VTAIL.n90 VSUBS 0.035834f
C1364 VTAIL.n91 VSUBS 0.016052f
C1365 VTAIL.n92 VSUBS 0.015161f
C1366 VTAIL.n93 VSUBS 0.028213f
C1367 VTAIL.n94 VSUBS 0.028213f
C1368 VTAIL.n95 VSUBS 0.015161f
C1369 VTAIL.n96 VSUBS 0.016052f
C1370 VTAIL.n97 VSUBS 0.035834f
C1371 VTAIL.n98 VSUBS 0.088792f
C1372 VTAIL.n99 VSUBS 0.016052f
C1373 VTAIL.n100 VSUBS 0.015161f
C1374 VTAIL.n101 VSUBS 0.067526f
C1375 VTAIL.n102 VSUBS 0.044814f
C1376 VTAIL.n103 VSUBS 0.192722f
C1377 VTAIL.t8 VSUBS 0.407996f
C1378 VTAIL.t14 VSUBS 0.407996f
C1379 VTAIL.n104 VSUBS 3.22942f
C1380 VTAIL.n105 VSUBS 0.852305f
C1381 VTAIL.t16 VSUBS 0.407996f
C1382 VTAIL.t10 VSUBS 0.407996f
C1383 VTAIL.n106 VSUBS 3.22942f
C1384 VTAIL.n107 VSUBS 2.75279f
C1385 VTAIL.t3 VSUBS 0.407996f
C1386 VTAIL.t7 VSUBS 0.407996f
C1387 VTAIL.n108 VSUBS 3.22944f
C1388 VTAIL.n109 VSUBS 2.75277f
C1389 VTAIL.t19 VSUBS 0.407996f
C1390 VTAIL.t5 VSUBS 0.407996f
C1391 VTAIL.n110 VSUBS 3.22944f
C1392 VTAIL.n111 VSUBS 0.852286f
C1393 VTAIL.n112 VSUBS 0.0316f
C1394 VTAIL.n113 VSUBS 0.028213f
C1395 VTAIL.n114 VSUBS 0.015161f
C1396 VTAIL.n115 VSUBS 0.035834f
C1397 VTAIL.n116 VSUBS 0.016052f
C1398 VTAIL.n117 VSUBS 0.028213f
C1399 VTAIL.n118 VSUBS 0.015161f
C1400 VTAIL.n119 VSUBS 0.035834f
C1401 VTAIL.n120 VSUBS 0.016052f
C1402 VTAIL.n121 VSUBS 0.028213f
C1403 VTAIL.n122 VSUBS 0.015606f
C1404 VTAIL.n123 VSUBS 0.035834f
C1405 VTAIL.n124 VSUBS 0.015161f
C1406 VTAIL.n125 VSUBS 0.016052f
C1407 VTAIL.n126 VSUBS 0.028213f
C1408 VTAIL.n127 VSUBS 0.015161f
C1409 VTAIL.n128 VSUBS 0.035834f
C1410 VTAIL.n129 VSUBS 0.016052f
C1411 VTAIL.n130 VSUBS 0.028213f
C1412 VTAIL.n131 VSUBS 0.015161f
C1413 VTAIL.n132 VSUBS 0.035834f
C1414 VTAIL.n133 VSUBS 0.016052f
C1415 VTAIL.n134 VSUBS 0.028213f
C1416 VTAIL.n135 VSUBS 0.015161f
C1417 VTAIL.n136 VSUBS 0.035834f
C1418 VTAIL.n137 VSUBS 0.016052f
C1419 VTAIL.n138 VSUBS 0.028213f
C1420 VTAIL.n139 VSUBS 0.015161f
C1421 VTAIL.n140 VSUBS 0.035834f
C1422 VTAIL.n141 VSUBS 0.016052f
C1423 VTAIL.n142 VSUBS 0.028213f
C1424 VTAIL.n143 VSUBS 0.015161f
C1425 VTAIL.n144 VSUBS 0.026875f
C1426 VTAIL.n145 VSUBS 0.022796f
C1427 VTAIL.t18 VSUBS 0.076945f
C1428 VTAIL.n146 VSUBS 0.226339f
C1429 VTAIL.n147 VSUBS 2.22413f
C1430 VTAIL.n148 VSUBS 0.015161f
C1431 VTAIL.n149 VSUBS 0.016052f
C1432 VTAIL.n150 VSUBS 0.035834f
C1433 VTAIL.n151 VSUBS 0.035834f
C1434 VTAIL.n152 VSUBS 0.016052f
C1435 VTAIL.n153 VSUBS 0.015161f
C1436 VTAIL.n154 VSUBS 0.028213f
C1437 VTAIL.n155 VSUBS 0.028213f
C1438 VTAIL.n156 VSUBS 0.015161f
C1439 VTAIL.n157 VSUBS 0.016052f
C1440 VTAIL.n158 VSUBS 0.035834f
C1441 VTAIL.n159 VSUBS 0.035834f
C1442 VTAIL.n160 VSUBS 0.016052f
C1443 VTAIL.n161 VSUBS 0.015161f
C1444 VTAIL.n162 VSUBS 0.028213f
C1445 VTAIL.n163 VSUBS 0.028213f
C1446 VTAIL.n164 VSUBS 0.015161f
C1447 VTAIL.n165 VSUBS 0.016052f
C1448 VTAIL.n166 VSUBS 0.035834f
C1449 VTAIL.n167 VSUBS 0.035834f
C1450 VTAIL.n168 VSUBS 0.016052f
C1451 VTAIL.n169 VSUBS 0.015161f
C1452 VTAIL.n170 VSUBS 0.028213f
C1453 VTAIL.n171 VSUBS 0.028213f
C1454 VTAIL.n172 VSUBS 0.015161f
C1455 VTAIL.n173 VSUBS 0.016052f
C1456 VTAIL.n174 VSUBS 0.035834f
C1457 VTAIL.n175 VSUBS 0.035834f
C1458 VTAIL.n176 VSUBS 0.016052f
C1459 VTAIL.n177 VSUBS 0.015161f
C1460 VTAIL.n178 VSUBS 0.028213f
C1461 VTAIL.n179 VSUBS 0.028213f
C1462 VTAIL.n180 VSUBS 0.015161f
C1463 VTAIL.n181 VSUBS 0.016052f
C1464 VTAIL.n182 VSUBS 0.035834f
C1465 VTAIL.n183 VSUBS 0.035834f
C1466 VTAIL.n184 VSUBS 0.016052f
C1467 VTAIL.n185 VSUBS 0.015161f
C1468 VTAIL.n186 VSUBS 0.028213f
C1469 VTAIL.n187 VSUBS 0.028213f
C1470 VTAIL.n188 VSUBS 0.015161f
C1471 VTAIL.n189 VSUBS 0.016052f
C1472 VTAIL.n190 VSUBS 0.035834f
C1473 VTAIL.n191 VSUBS 0.035834f
C1474 VTAIL.n192 VSUBS 0.035834f
C1475 VTAIL.n193 VSUBS 0.015606f
C1476 VTAIL.n194 VSUBS 0.015161f
C1477 VTAIL.n195 VSUBS 0.028213f
C1478 VTAIL.n196 VSUBS 0.028213f
C1479 VTAIL.n197 VSUBS 0.015161f
C1480 VTAIL.n198 VSUBS 0.016052f
C1481 VTAIL.n199 VSUBS 0.035834f
C1482 VTAIL.n200 VSUBS 0.035834f
C1483 VTAIL.n201 VSUBS 0.016052f
C1484 VTAIL.n202 VSUBS 0.015161f
C1485 VTAIL.n203 VSUBS 0.028213f
C1486 VTAIL.n204 VSUBS 0.028213f
C1487 VTAIL.n205 VSUBS 0.015161f
C1488 VTAIL.n206 VSUBS 0.016052f
C1489 VTAIL.n207 VSUBS 0.035834f
C1490 VTAIL.n208 VSUBS 0.088792f
C1491 VTAIL.n209 VSUBS 0.016052f
C1492 VTAIL.n210 VSUBS 0.015161f
C1493 VTAIL.n211 VSUBS 0.067526f
C1494 VTAIL.n212 VSUBS 0.044814f
C1495 VTAIL.n213 VSUBS 0.192722f
C1496 VTAIL.t11 VSUBS 0.407996f
C1497 VTAIL.t15 VSUBS 0.407996f
C1498 VTAIL.n214 VSUBS 3.22944f
C1499 VTAIL.n215 VSUBS 0.853462f
C1500 VTAIL.t17 VSUBS 0.407996f
C1501 VTAIL.t12 VSUBS 0.407996f
C1502 VTAIL.n216 VSUBS 3.22944f
C1503 VTAIL.n217 VSUBS 0.852286f
C1504 VTAIL.n218 VSUBS 0.0316f
C1505 VTAIL.n219 VSUBS 0.028213f
C1506 VTAIL.n220 VSUBS 0.015161f
C1507 VTAIL.n221 VSUBS 0.035834f
C1508 VTAIL.n222 VSUBS 0.016052f
C1509 VTAIL.n223 VSUBS 0.028213f
C1510 VTAIL.n224 VSUBS 0.015161f
C1511 VTAIL.n225 VSUBS 0.035834f
C1512 VTAIL.n226 VSUBS 0.016052f
C1513 VTAIL.n227 VSUBS 0.028213f
C1514 VTAIL.n228 VSUBS 0.015606f
C1515 VTAIL.n229 VSUBS 0.035834f
C1516 VTAIL.n230 VSUBS 0.015161f
C1517 VTAIL.n231 VSUBS 0.016052f
C1518 VTAIL.n232 VSUBS 0.028213f
C1519 VTAIL.n233 VSUBS 0.015161f
C1520 VTAIL.n234 VSUBS 0.035834f
C1521 VTAIL.n235 VSUBS 0.016052f
C1522 VTAIL.n236 VSUBS 0.028213f
C1523 VTAIL.n237 VSUBS 0.015161f
C1524 VTAIL.n238 VSUBS 0.035834f
C1525 VTAIL.n239 VSUBS 0.016052f
C1526 VTAIL.n240 VSUBS 0.028213f
C1527 VTAIL.n241 VSUBS 0.015161f
C1528 VTAIL.n242 VSUBS 0.035834f
C1529 VTAIL.n243 VSUBS 0.016052f
C1530 VTAIL.n244 VSUBS 0.028213f
C1531 VTAIL.n245 VSUBS 0.015161f
C1532 VTAIL.n246 VSUBS 0.035834f
C1533 VTAIL.n247 VSUBS 0.016052f
C1534 VTAIL.n248 VSUBS 0.028213f
C1535 VTAIL.n249 VSUBS 0.015161f
C1536 VTAIL.n250 VSUBS 0.026875f
C1537 VTAIL.n251 VSUBS 0.022796f
C1538 VTAIL.t13 VSUBS 0.076945f
C1539 VTAIL.n252 VSUBS 0.226339f
C1540 VTAIL.n253 VSUBS 2.22413f
C1541 VTAIL.n254 VSUBS 0.015161f
C1542 VTAIL.n255 VSUBS 0.016052f
C1543 VTAIL.n256 VSUBS 0.035834f
C1544 VTAIL.n257 VSUBS 0.035834f
C1545 VTAIL.n258 VSUBS 0.016052f
C1546 VTAIL.n259 VSUBS 0.015161f
C1547 VTAIL.n260 VSUBS 0.028213f
C1548 VTAIL.n261 VSUBS 0.028213f
C1549 VTAIL.n262 VSUBS 0.015161f
C1550 VTAIL.n263 VSUBS 0.016052f
C1551 VTAIL.n264 VSUBS 0.035834f
C1552 VTAIL.n265 VSUBS 0.035834f
C1553 VTAIL.n266 VSUBS 0.016052f
C1554 VTAIL.n267 VSUBS 0.015161f
C1555 VTAIL.n268 VSUBS 0.028213f
C1556 VTAIL.n269 VSUBS 0.028213f
C1557 VTAIL.n270 VSUBS 0.015161f
C1558 VTAIL.n271 VSUBS 0.016052f
C1559 VTAIL.n272 VSUBS 0.035834f
C1560 VTAIL.n273 VSUBS 0.035834f
C1561 VTAIL.n274 VSUBS 0.016052f
C1562 VTAIL.n275 VSUBS 0.015161f
C1563 VTAIL.n276 VSUBS 0.028213f
C1564 VTAIL.n277 VSUBS 0.028213f
C1565 VTAIL.n278 VSUBS 0.015161f
C1566 VTAIL.n279 VSUBS 0.016052f
C1567 VTAIL.n280 VSUBS 0.035834f
C1568 VTAIL.n281 VSUBS 0.035834f
C1569 VTAIL.n282 VSUBS 0.016052f
C1570 VTAIL.n283 VSUBS 0.015161f
C1571 VTAIL.n284 VSUBS 0.028213f
C1572 VTAIL.n285 VSUBS 0.028213f
C1573 VTAIL.n286 VSUBS 0.015161f
C1574 VTAIL.n287 VSUBS 0.016052f
C1575 VTAIL.n288 VSUBS 0.035834f
C1576 VTAIL.n289 VSUBS 0.035834f
C1577 VTAIL.n290 VSUBS 0.016052f
C1578 VTAIL.n291 VSUBS 0.015161f
C1579 VTAIL.n292 VSUBS 0.028213f
C1580 VTAIL.n293 VSUBS 0.028213f
C1581 VTAIL.n294 VSUBS 0.015161f
C1582 VTAIL.n295 VSUBS 0.016052f
C1583 VTAIL.n296 VSUBS 0.035834f
C1584 VTAIL.n297 VSUBS 0.035834f
C1585 VTAIL.n298 VSUBS 0.035834f
C1586 VTAIL.n299 VSUBS 0.015606f
C1587 VTAIL.n300 VSUBS 0.015161f
C1588 VTAIL.n301 VSUBS 0.028213f
C1589 VTAIL.n302 VSUBS 0.028213f
C1590 VTAIL.n303 VSUBS 0.015161f
C1591 VTAIL.n304 VSUBS 0.016052f
C1592 VTAIL.n305 VSUBS 0.035834f
C1593 VTAIL.n306 VSUBS 0.035834f
C1594 VTAIL.n307 VSUBS 0.016052f
C1595 VTAIL.n308 VSUBS 0.015161f
C1596 VTAIL.n309 VSUBS 0.028213f
C1597 VTAIL.n310 VSUBS 0.028213f
C1598 VTAIL.n311 VSUBS 0.015161f
C1599 VTAIL.n312 VSUBS 0.016052f
C1600 VTAIL.n313 VSUBS 0.035834f
C1601 VTAIL.n314 VSUBS 0.088792f
C1602 VTAIL.n315 VSUBS 0.016052f
C1603 VTAIL.n316 VSUBS 0.015161f
C1604 VTAIL.n317 VSUBS 0.067526f
C1605 VTAIL.n318 VSUBS 0.044814f
C1606 VTAIL.n319 VSUBS 2.00895f
C1607 VTAIL.n320 VSUBS 0.0316f
C1608 VTAIL.n321 VSUBS 0.028213f
C1609 VTAIL.n322 VSUBS 0.015161f
C1610 VTAIL.n323 VSUBS 0.035834f
C1611 VTAIL.n324 VSUBS 0.016052f
C1612 VTAIL.n325 VSUBS 0.028213f
C1613 VTAIL.n326 VSUBS 0.015161f
C1614 VTAIL.n327 VSUBS 0.035834f
C1615 VTAIL.n328 VSUBS 0.016052f
C1616 VTAIL.n329 VSUBS 0.028213f
C1617 VTAIL.n330 VSUBS 0.015606f
C1618 VTAIL.n331 VSUBS 0.035834f
C1619 VTAIL.n332 VSUBS 0.016052f
C1620 VTAIL.n333 VSUBS 0.028213f
C1621 VTAIL.n334 VSUBS 0.015161f
C1622 VTAIL.n335 VSUBS 0.035834f
C1623 VTAIL.n336 VSUBS 0.016052f
C1624 VTAIL.n337 VSUBS 0.028213f
C1625 VTAIL.n338 VSUBS 0.015161f
C1626 VTAIL.n339 VSUBS 0.035834f
C1627 VTAIL.n340 VSUBS 0.016052f
C1628 VTAIL.n341 VSUBS 0.028213f
C1629 VTAIL.n342 VSUBS 0.015161f
C1630 VTAIL.n343 VSUBS 0.035834f
C1631 VTAIL.n344 VSUBS 0.016052f
C1632 VTAIL.n345 VSUBS 0.028213f
C1633 VTAIL.n346 VSUBS 0.015161f
C1634 VTAIL.n347 VSUBS 0.035834f
C1635 VTAIL.n348 VSUBS 0.016052f
C1636 VTAIL.n349 VSUBS 0.028213f
C1637 VTAIL.n350 VSUBS 0.015161f
C1638 VTAIL.n351 VSUBS 0.026875f
C1639 VTAIL.n352 VSUBS 0.022796f
C1640 VTAIL.t4 VSUBS 0.076945f
C1641 VTAIL.n353 VSUBS 0.226339f
C1642 VTAIL.n354 VSUBS 2.22413f
C1643 VTAIL.n355 VSUBS 0.015161f
C1644 VTAIL.n356 VSUBS 0.016052f
C1645 VTAIL.n357 VSUBS 0.035834f
C1646 VTAIL.n358 VSUBS 0.035834f
C1647 VTAIL.n359 VSUBS 0.016052f
C1648 VTAIL.n360 VSUBS 0.015161f
C1649 VTAIL.n361 VSUBS 0.028213f
C1650 VTAIL.n362 VSUBS 0.028213f
C1651 VTAIL.n363 VSUBS 0.015161f
C1652 VTAIL.n364 VSUBS 0.016052f
C1653 VTAIL.n365 VSUBS 0.035834f
C1654 VTAIL.n366 VSUBS 0.035834f
C1655 VTAIL.n367 VSUBS 0.016052f
C1656 VTAIL.n368 VSUBS 0.015161f
C1657 VTAIL.n369 VSUBS 0.028213f
C1658 VTAIL.n370 VSUBS 0.028213f
C1659 VTAIL.n371 VSUBS 0.015161f
C1660 VTAIL.n372 VSUBS 0.016052f
C1661 VTAIL.n373 VSUBS 0.035834f
C1662 VTAIL.n374 VSUBS 0.035834f
C1663 VTAIL.n375 VSUBS 0.016052f
C1664 VTAIL.n376 VSUBS 0.015161f
C1665 VTAIL.n377 VSUBS 0.028213f
C1666 VTAIL.n378 VSUBS 0.028213f
C1667 VTAIL.n379 VSUBS 0.015161f
C1668 VTAIL.n380 VSUBS 0.016052f
C1669 VTAIL.n381 VSUBS 0.035834f
C1670 VTAIL.n382 VSUBS 0.035834f
C1671 VTAIL.n383 VSUBS 0.016052f
C1672 VTAIL.n384 VSUBS 0.015161f
C1673 VTAIL.n385 VSUBS 0.028213f
C1674 VTAIL.n386 VSUBS 0.028213f
C1675 VTAIL.n387 VSUBS 0.015161f
C1676 VTAIL.n388 VSUBS 0.016052f
C1677 VTAIL.n389 VSUBS 0.035834f
C1678 VTAIL.n390 VSUBS 0.035834f
C1679 VTAIL.n391 VSUBS 0.016052f
C1680 VTAIL.n392 VSUBS 0.015161f
C1681 VTAIL.n393 VSUBS 0.028213f
C1682 VTAIL.n394 VSUBS 0.028213f
C1683 VTAIL.n395 VSUBS 0.015161f
C1684 VTAIL.n396 VSUBS 0.015161f
C1685 VTAIL.n397 VSUBS 0.016052f
C1686 VTAIL.n398 VSUBS 0.035834f
C1687 VTAIL.n399 VSUBS 0.035834f
C1688 VTAIL.n400 VSUBS 0.035834f
C1689 VTAIL.n401 VSUBS 0.015606f
C1690 VTAIL.n402 VSUBS 0.015161f
C1691 VTAIL.n403 VSUBS 0.028213f
C1692 VTAIL.n404 VSUBS 0.028213f
C1693 VTAIL.n405 VSUBS 0.015161f
C1694 VTAIL.n406 VSUBS 0.016052f
C1695 VTAIL.n407 VSUBS 0.035834f
C1696 VTAIL.n408 VSUBS 0.035834f
C1697 VTAIL.n409 VSUBS 0.016052f
C1698 VTAIL.n410 VSUBS 0.015161f
C1699 VTAIL.n411 VSUBS 0.028213f
C1700 VTAIL.n412 VSUBS 0.028213f
C1701 VTAIL.n413 VSUBS 0.015161f
C1702 VTAIL.n414 VSUBS 0.016052f
C1703 VTAIL.n415 VSUBS 0.035834f
C1704 VTAIL.n416 VSUBS 0.088792f
C1705 VTAIL.n417 VSUBS 0.016052f
C1706 VTAIL.n418 VSUBS 0.015161f
C1707 VTAIL.n419 VSUBS 0.067526f
C1708 VTAIL.n420 VSUBS 0.044814f
C1709 VTAIL.n421 VSUBS 2.00895f
C1710 VTAIL.t6 VSUBS 0.407996f
C1711 VTAIL.t2 VSUBS 0.407996f
C1712 VTAIL.n422 VSUBS 3.22942f
C1713 VTAIL.n423 VSUBS 0.784711f
C1714 VP.n0 VSUBS 0.049256f
C1715 VP.n1 VSUBS 0.011177f
C1716 VP.n2 VSUBS 0.049256f
C1717 VP.n3 VSUBS 0.011177f
C1718 VP.n4 VSUBS 0.049256f
C1719 VP.t1 VSUBS 1.86521f
C1720 VP.t5 VSUBS 1.86521f
C1721 VP.n5 VSUBS 0.049256f
C1722 VP.t2 VSUBS 1.86521f
C1723 VP.n6 VSUBS 0.700957f
C1724 VP.t0 VSUBS 1.89029f
C1725 VP.n7 VSUBS 0.680901f
C1726 VP.t3 VSUBS 1.86521f
C1727 VP.n8 VSUBS 0.707704f
C1728 VP.n9 VSUBS 0.011177f
C1729 VP.n10 VSUBS 0.210246f
C1730 VP.n11 VSUBS 0.049256f
C1731 VP.n12 VSUBS 0.049256f
C1732 VP.n13 VSUBS 0.011177f
C1733 VP.n14 VSUBS 0.700957f
C1734 VP.n15 VSUBS 0.011177f
C1735 VP.n16 VSUBS 0.700501f
C1736 VP.n17 VSUBS 2.49847f
C1737 VP.t4 VSUBS 1.86521f
C1738 VP.n18 VSUBS 0.700501f
C1739 VP.n19 VSUBS 2.53564f
C1740 VP.n20 VSUBS 0.049256f
C1741 VP.n21 VSUBS 0.049256f
C1742 VP.t6 VSUBS 1.86521f
C1743 VP.n22 VSUBS 0.700957f
C1744 VP.n23 VSUBS 0.011177f
C1745 VP.t8 VSUBS 1.86521f
C1746 VP.n24 VSUBS 0.700957f
C1747 VP.n25 VSUBS 0.049256f
C1748 VP.n26 VSUBS 0.049256f
C1749 VP.n27 VSUBS 0.049256f
C1750 VP.t7 VSUBS 1.86521f
C1751 VP.n28 VSUBS 0.700957f
C1752 VP.n29 VSUBS 0.011177f
C1753 VP.t9 VSUBS 1.86521f
C1754 VP.n30 VSUBS 0.700501f
C1755 VP.n31 VSUBS 0.038171f
.ends

