* NGSPICE file created from diff_pair_sample_1372.ext - technology: sky130A

.subckt diff_pair_sample_1372 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=1.2
X1 B.t11 B.t9 B.t10 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=1.2
X2 VDD1.t4 VP.t1 VTAIL.t9 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=1.2
X3 VDD2.t5 VN.t0 VTAIL.t4 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=1.2
X4 VDD2.t4 VN.t1 VTAIL.t3 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=1.2
X5 B.t8 B.t6 B.t7 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=1.2
X6 VTAIL.t11 VN.t2 VDD2.t3 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=1.2
X7 VDD1.t3 VP.t2 VTAIL.t6 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=1.2
X8 B.t5 B.t3 B.t4 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=1.2
X9 VTAIL.t10 VP.t3 VDD1.t2 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=1.2
X10 VDD2.t2 VN.t3 VTAIL.t0 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=1.2
X11 VDD1.t1 VP.t4 VTAIL.t7 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=1.2
X12 VTAIL.t1 VN.t4 VDD2.t1 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=1.2
X13 VTAIL.t5 VP.t5 VDD1.t0 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=1.2
X14 B.t2 B.t0 B.t1 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=1.2
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n2194_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=1.2
R0 VP.n7 VP.t2 272.635
R1 VP.n3 VP.t1 241.602
R2 VP.n18 VP.t3 241.602
R3 VP.n25 VP.t4 241.602
R4 VP.n12 VP.t0 241.602
R5 VP.n6 VP.t5 241.602
R6 VP.n14 VP.n3 172.065
R7 VP.n26 VP.n25 172.065
R8 VP.n13 VP.n12 172.065
R9 VP.n8 VP.n5 161.3
R10 VP.n10 VP.n9 161.3
R11 VP.n11 VP.n4 161.3
R12 VP.n24 VP.n0 161.3
R13 VP.n23 VP.n22 161.3
R14 VP.n21 VP.n1 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n17 VP.n2 161.3
R17 VP.n16 VP.n15 161.3
R18 VP.n7 VP.n6 51.3222
R19 VP.n14 VP.n13 43.1179
R20 VP.n17 VP.n16 41.9503
R21 VP.n24 VP.n23 41.9503
R22 VP.n11 VP.n10 41.9503
R23 VP.n19 VP.n17 39.0365
R24 VP.n23 VP.n1 39.0365
R25 VP.n10 VP.n5 39.0365
R26 VP.n8 VP.n7 26.7683
R27 VP.n16 VP.n3 13.702
R28 VP.n25 VP.n24 13.702
R29 VP.n12 VP.n11 13.702
R30 VP.n19 VP.n18 12.234
R31 VP.n18 VP.n1 12.234
R32 VP.n6 VP.n5 12.234
R33 VP.n9 VP.n8 0.189894
R34 VP.n9 VP.n4 0.189894
R35 VP.n13 VP.n4 0.189894
R36 VP.n15 VP.n14 0.189894
R37 VP.n15 VP.n2 0.189894
R38 VP.n20 VP.n2 0.189894
R39 VP.n21 VP.n20 0.189894
R40 VP.n22 VP.n21 0.189894
R41 VP.n22 VP.n0 0.189894
R42 VP.n26 VP.n0 0.189894
R43 VP VP.n26 0.0516364
R44 VTAIL.n266 VTAIL.n206 756.745
R45 VTAIL.n62 VTAIL.n2 756.745
R46 VTAIL.n200 VTAIL.n140 756.745
R47 VTAIL.n132 VTAIL.n72 756.745
R48 VTAIL.n226 VTAIL.n225 585
R49 VTAIL.n231 VTAIL.n230 585
R50 VTAIL.n233 VTAIL.n232 585
R51 VTAIL.n222 VTAIL.n221 585
R52 VTAIL.n239 VTAIL.n238 585
R53 VTAIL.n241 VTAIL.n240 585
R54 VTAIL.n218 VTAIL.n217 585
R55 VTAIL.n248 VTAIL.n247 585
R56 VTAIL.n249 VTAIL.n216 585
R57 VTAIL.n251 VTAIL.n250 585
R58 VTAIL.n214 VTAIL.n213 585
R59 VTAIL.n257 VTAIL.n256 585
R60 VTAIL.n259 VTAIL.n258 585
R61 VTAIL.n210 VTAIL.n209 585
R62 VTAIL.n265 VTAIL.n264 585
R63 VTAIL.n267 VTAIL.n266 585
R64 VTAIL.n22 VTAIL.n21 585
R65 VTAIL.n27 VTAIL.n26 585
R66 VTAIL.n29 VTAIL.n28 585
R67 VTAIL.n18 VTAIL.n17 585
R68 VTAIL.n35 VTAIL.n34 585
R69 VTAIL.n37 VTAIL.n36 585
R70 VTAIL.n14 VTAIL.n13 585
R71 VTAIL.n44 VTAIL.n43 585
R72 VTAIL.n45 VTAIL.n12 585
R73 VTAIL.n47 VTAIL.n46 585
R74 VTAIL.n10 VTAIL.n9 585
R75 VTAIL.n53 VTAIL.n52 585
R76 VTAIL.n55 VTAIL.n54 585
R77 VTAIL.n6 VTAIL.n5 585
R78 VTAIL.n61 VTAIL.n60 585
R79 VTAIL.n63 VTAIL.n62 585
R80 VTAIL.n201 VTAIL.n200 585
R81 VTAIL.n199 VTAIL.n198 585
R82 VTAIL.n144 VTAIL.n143 585
R83 VTAIL.n193 VTAIL.n192 585
R84 VTAIL.n191 VTAIL.n190 585
R85 VTAIL.n148 VTAIL.n147 585
R86 VTAIL.n185 VTAIL.n184 585
R87 VTAIL.n183 VTAIL.n150 585
R88 VTAIL.n182 VTAIL.n181 585
R89 VTAIL.n153 VTAIL.n151 585
R90 VTAIL.n176 VTAIL.n175 585
R91 VTAIL.n174 VTAIL.n173 585
R92 VTAIL.n157 VTAIL.n156 585
R93 VTAIL.n168 VTAIL.n167 585
R94 VTAIL.n166 VTAIL.n165 585
R95 VTAIL.n161 VTAIL.n160 585
R96 VTAIL.n133 VTAIL.n132 585
R97 VTAIL.n131 VTAIL.n130 585
R98 VTAIL.n76 VTAIL.n75 585
R99 VTAIL.n125 VTAIL.n124 585
R100 VTAIL.n123 VTAIL.n122 585
R101 VTAIL.n80 VTAIL.n79 585
R102 VTAIL.n117 VTAIL.n116 585
R103 VTAIL.n115 VTAIL.n82 585
R104 VTAIL.n114 VTAIL.n113 585
R105 VTAIL.n85 VTAIL.n83 585
R106 VTAIL.n108 VTAIL.n107 585
R107 VTAIL.n106 VTAIL.n105 585
R108 VTAIL.n89 VTAIL.n88 585
R109 VTAIL.n100 VTAIL.n99 585
R110 VTAIL.n98 VTAIL.n97 585
R111 VTAIL.n93 VTAIL.n92 585
R112 VTAIL.n227 VTAIL.t3 329.036
R113 VTAIL.n23 VTAIL.t7 329.036
R114 VTAIL.n162 VTAIL.t8 329.036
R115 VTAIL.n94 VTAIL.t4 329.036
R116 VTAIL.n231 VTAIL.n225 171.744
R117 VTAIL.n232 VTAIL.n231 171.744
R118 VTAIL.n232 VTAIL.n221 171.744
R119 VTAIL.n239 VTAIL.n221 171.744
R120 VTAIL.n240 VTAIL.n239 171.744
R121 VTAIL.n240 VTAIL.n217 171.744
R122 VTAIL.n248 VTAIL.n217 171.744
R123 VTAIL.n249 VTAIL.n248 171.744
R124 VTAIL.n250 VTAIL.n249 171.744
R125 VTAIL.n250 VTAIL.n213 171.744
R126 VTAIL.n257 VTAIL.n213 171.744
R127 VTAIL.n258 VTAIL.n257 171.744
R128 VTAIL.n258 VTAIL.n209 171.744
R129 VTAIL.n265 VTAIL.n209 171.744
R130 VTAIL.n266 VTAIL.n265 171.744
R131 VTAIL.n27 VTAIL.n21 171.744
R132 VTAIL.n28 VTAIL.n27 171.744
R133 VTAIL.n28 VTAIL.n17 171.744
R134 VTAIL.n35 VTAIL.n17 171.744
R135 VTAIL.n36 VTAIL.n35 171.744
R136 VTAIL.n36 VTAIL.n13 171.744
R137 VTAIL.n44 VTAIL.n13 171.744
R138 VTAIL.n45 VTAIL.n44 171.744
R139 VTAIL.n46 VTAIL.n45 171.744
R140 VTAIL.n46 VTAIL.n9 171.744
R141 VTAIL.n53 VTAIL.n9 171.744
R142 VTAIL.n54 VTAIL.n53 171.744
R143 VTAIL.n54 VTAIL.n5 171.744
R144 VTAIL.n61 VTAIL.n5 171.744
R145 VTAIL.n62 VTAIL.n61 171.744
R146 VTAIL.n200 VTAIL.n199 171.744
R147 VTAIL.n199 VTAIL.n143 171.744
R148 VTAIL.n192 VTAIL.n143 171.744
R149 VTAIL.n192 VTAIL.n191 171.744
R150 VTAIL.n191 VTAIL.n147 171.744
R151 VTAIL.n184 VTAIL.n147 171.744
R152 VTAIL.n184 VTAIL.n183 171.744
R153 VTAIL.n183 VTAIL.n182 171.744
R154 VTAIL.n182 VTAIL.n151 171.744
R155 VTAIL.n175 VTAIL.n151 171.744
R156 VTAIL.n175 VTAIL.n174 171.744
R157 VTAIL.n174 VTAIL.n156 171.744
R158 VTAIL.n167 VTAIL.n156 171.744
R159 VTAIL.n167 VTAIL.n166 171.744
R160 VTAIL.n166 VTAIL.n160 171.744
R161 VTAIL.n132 VTAIL.n131 171.744
R162 VTAIL.n131 VTAIL.n75 171.744
R163 VTAIL.n124 VTAIL.n75 171.744
R164 VTAIL.n124 VTAIL.n123 171.744
R165 VTAIL.n123 VTAIL.n79 171.744
R166 VTAIL.n116 VTAIL.n79 171.744
R167 VTAIL.n116 VTAIL.n115 171.744
R168 VTAIL.n115 VTAIL.n114 171.744
R169 VTAIL.n114 VTAIL.n83 171.744
R170 VTAIL.n107 VTAIL.n83 171.744
R171 VTAIL.n107 VTAIL.n106 171.744
R172 VTAIL.n106 VTAIL.n88 171.744
R173 VTAIL.n99 VTAIL.n88 171.744
R174 VTAIL.n99 VTAIL.n98 171.744
R175 VTAIL.n98 VTAIL.n92 171.744
R176 VTAIL.t3 VTAIL.n225 85.8723
R177 VTAIL.t7 VTAIL.n21 85.8723
R178 VTAIL.t8 VTAIL.n160 85.8723
R179 VTAIL.t4 VTAIL.n92 85.8723
R180 VTAIL.n139 VTAIL.n138 55.415
R181 VTAIL.n71 VTAIL.n70 55.415
R182 VTAIL.n1 VTAIL.n0 55.4148
R183 VTAIL.n69 VTAIL.n68 55.4148
R184 VTAIL.n271 VTAIL.n270 30.4399
R185 VTAIL.n67 VTAIL.n66 30.4399
R186 VTAIL.n205 VTAIL.n204 30.4399
R187 VTAIL.n137 VTAIL.n136 30.4399
R188 VTAIL.n71 VTAIL.n69 25.3755
R189 VTAIL.n271 VTAIL.n205 24.0565
R190 VTAIL.n251 VTAIL.n216 13.1884
R191 VTAIL.n47 VTAIL.n12 13.1884
R192 VTAIL.n185 VTAIL.n150 13.1884
R193 VTAIL.n117 VTAIL.n82 13.1884
R194 VTAIL.n247 VTAIL.n246 12.8005
R195 VTAIL.n252 VTAIL.n214 12.8005
R196 VTAIL.n43 VTAIL.n42 12.8005
R197 VTAIL.n48 VTAIL.n10 12.8005
R198 VTAIL.n186 VTAIL.n148 12.8005
R199 VTAIL.n181 VTAIL.n152 12.8005
R200 VTAIL.n118 VTAIL.n80 12.8005
R201 VTAIL.n113 VTAIL.n84 12.8005
R202 VTAIL.n245 VTAIL.n218 12.0247
R203 VTAIL.n256 VTAIL.n255 12.0247
R204 VTAIL.n41 VTAIL.n14 12.0247
R205 VTAIL.n52 VTAIL.n51 12.0247
R206 VTAIL.n190 VTAIL.n189 12.0247
R207 VTAIL.n180 VTAIL.n153 12.0247
R208 VTAIL.n122 VTAIL.n121 12.0247
R209 VTAIL.n112 VTAIL.n85 12.0247
R210 VTAIL.n242 VTAIL.n241 11.249
R211 VTAIL.n259 VTAIL.n212 11.249
R212 VTAIL.n38 VTAIL.n37 11.249
R213 VTAIL.n55 VTAIL.n8 11.249
R214 VTAIL.n193 VTAIL.n146 11.249
R215 VTAIL.n177 VTAIL.n176 11.249
R216 VTAIL.n125 VTAIL.n78 11.249
R217 VTAIL.n109 VTAIL.n108 11.249
R218 VTAIL.n227 VTAIL.n226 10.7239
R219 VTAIL.n23 VTAIL.n22 10.7239
R220 VTAIL.n162 VTAIL.n161 10.7239
R221 VTAIL.n94 VTAIL.n93 10.7239
R222 VTAIL.n238 VTAIL.n220 10.4732
R223 VTAIL.n260 VTAIL.n210 10.4732
R224 VTAIL.n34 VTAIL.n16 10.4732
R225 VTAIL.n56 VTAIL.n6 10.4732
R226 VTAIL.n194 VTAIL.n144 10.4732
R227 VTAIL.n173 VTAIL.n155 10.4732
R228 VTAIL.n126 VTAIL.n76 10.4732
R229 VTAIL.n105 VTAIL.n87 10.4732
R230 VTAIL.n237 VTAIL.n222 9.69747
R231 VTAIL.n264 VTAIL.n263 9.69747
R232 VTAIL.n33 VTAIL.n18 9.69747
R233 VTAIL.n60 VTAIL.n59 9.69747
R234 VTAIL.n198 VTAIL.n197 9.69747
R235 VTAIL.n172 VTAIL.n157 9.69747
R236 VTAIL.n130 VTAIL.n129 9.69747
R237 VTAIL.n104 VTAIL.n89 9.69747
R238 VTAIL.n270 VTAIL.n269 9.45567
R239 VTAIL.n66 VTAIL.n65 9.45567
R240 VTAIL.n204 VTAIL.n203 9.45567
R241 VTAIL.n136 VTAIL.n135 9.45567
R242 VTAIL.n269 VTAIL.n268 9.3005
R243 VTAIL.n208 VTAIL.n207 9.3005
R244 VTAIL.n263 VTAIL.n262 9.3005
R245 VTAIL.n261 VTAIL.n260 9.3005
R246 VTAIL.n212 VTAIL.n211 9.3005
R247 VTAIL.n255 VTAIL.n254 9.3005
R248 VTAIL.n253 VTAIL.n252 9.3005
R249 VTAIL.n229 VTAIL.n228 9.3005
R250 VTAIL.n224 VTAIL.n223 9.3005
R251 VTAIL.n235 VTAIL.n234 9.3005
R252 VTAIL.n237 VTAIL.n236 9.3005
R253 VTAIL.n220 VTAIL.n219 9.3005
R254 VTAIL.n243 VTAIL.n242 9.3005
R255 VTAIL.n245 VTAIL.n244 9.3005
R256 VTAIL.n246 VTAIL.n215 9.3005
R257 VTAIL.n65 VTAIL.n64 9.3005
R258 VTAIL.n4 VTAIL.n3 9.3005
R259 VTAIL.n59 VTAIL.n58 9.3005
R260 VTAIL.n57 VTAIL.n56 9.3005
R261 VTAIL.n8 VTAIL.n7 9.3005
R262 VTAIL.n51 VTAIL.n50 9.3005
R263 VTAIL.n49 VTAIL.n48 9.3005
R264 VTAIL.n25 VTAIL.n24 9.3005
R265 VTAIL.n20 VTAIL.n19 9.3005
R266 VTAIL.n31 VTAIL.n30 9.3005
R267 VTAIL.n33 VTAIL.n32 9.3005
R268 VTAIL.n16 VTAIL.n15 9.3005
R269 VTAIL.n39 VTAIL.n38 9.3005
R270 VTAIL.n41 VTAIL.n40 9.3005
R271 VTAIL.n42 VTAIL.n11 9.3005
R272 VTAIL.n164 VTAIL.n163 9.3005
R273 VTAIL.n159 VTAIL.n158 9.3005
R274 VTAIL.n170 VTAIL.n169 9.3005
R275 VTAIL.n172 VTAIL.n171 9.3005
R276 VTAIL.n155 VTAIL.n154 9.3005
R277 VTAIL.n178 VTAIL.n177 9.3005
R278 VTAIL.n180 VTAIL.n179 9.3005
R279 VTAIL.n152 VTAIL.n149 9.3005
R280 VTAIL.n203 VTAIL.n202 9.3005
R281 VTAIL.n142 VTAIL.n141 9.3005
R282 VTAIL.n197 VTAIL.n196 9.3005
R283 VTAIL.n195 VTAIL.n194 9.3005
R284 VTAIL.n146 VTAIL.n145 9.3005
R285 VTAIL.n189 VTAIL.n188 9.3005
R286 VTAIL.n187 VTAIL.n186 9.3005
R287 VTAIL.n96 VTAIL.n95 9.3005
R288 VTAIL.n91 VTAIL.n90 9.3005
R289 VTAIL.n102 VTAIL.n101 9.3005
R290 VTAIL.n104 VTAIL.n103 9.3005
R291 VTAIL.n87 VTAIL.n86 9.3005
R292 VTAIL.n110 VTAIL.n109 9.3005
R293 VTAIL.n112 VTAIL.n111 9.3005
R294 VTAIL.n84 VTAIL.n81 9.3005
R295 VTAIL.n135 VTAIL.n134 9.3005
R296 VTAIL.n74 VTAIL.n73 9.3005
R297 VTAIL.n129 VTAIL.n128 9.3005
R298 VTAIL.n127 VTAIL.n126 9.3005
R299 VTAIL.n78 VTAIL.n77 9.3005
R300 VTAIL.n121 VTAIL.n120 9.3005
R301 VTAIL.n119 VTAIL.n118 9.3005
R302 VTAIL.n234 VTAIL.n233 8.92171
R303 VTAIL.n267 VTAIL.n208 8.92171
R304 VTAIL.n30 VTAIL.n29 8.92171
R305 VTAIL.n63 VTAIL.n4 8.92171
R306 VTAIL.n201 VTAIL.n142 8.92171
R307 VTAIL.n169 VTAIL.n168 8.92171
R308 VTAIL.n133 VTAIL.n74 8.92171
R309 VTAIL.n101 VTAIL.n100 8.92171
R310 VTAIL.n230 VTAIL.n224 8.14595
R311 VTAIL.n268 VTAIL.n206 8.14595
R312 VTAIL.n26 VTAIL.n20 8.14595
R313 VTAIL.n64 VTAIL.n2 8.14595
R314 VTAIL.n202 VTAIL.n140 8.14595
R315 VTAIL.n165 VTAIL.n159 8.14595
R316 VTAIL.n134 VTAIL.n72 8.14595
R317 VTAIL.n97 VTAIL.n91 8.14595
R318 VTAIL.n229 VTAIL.n226 7.3702
R319 VTAIL.n25 VTAIL.n22 7.3702
R320 VTAIL.n164 VTAIL.n161 7.3702
R321 VTAIL.n96 VTAIL.n93 7.3702
R322 VTAIL.n230 VTAIL.n229 5.81868
R323 VTAIL.n270 VTAIL.n206 5.81868
R324 VTAIL.n26 VTAIL.n25 5.81868
R325 VTAIL.n66 VTAIL.n2 5.81868
R326 VTAIL.n204 VTAIL.n140 5.81868
R327 VTAIL.n165 VTAIL.n164 5.81868
R328 VTAIL.n136 VTAIL.n72 5.81868
R329 VTAIL.n97 VTAIL.n96 5.81868
R330 VTAIL.n233 VTAIL.n224 5.04292
R331 VTAIL.n268 VTAIL.n267 5.04292
R332 VTAIL.n29 VTAIL.n20 5.04292
R333 VTAIL.n64 VTAIL.n63 5.04292
R334 VTAIL.n202 VTAIL.n201 5.04292
R335 VTAIL.n168 VTAIL.n159 5.04292
R336 VTAIL.n134 VTAIL.n133 5.04292
R337 VTAIL.n100 VTAIL.n91 5.04292
R338 VTAIL.n234 VTAIL.n222 4.26717
R339 VTAIL.n264 VTAIL.n208 4.26717
R340 VTAIL.n30 VTAIL.n18 4.26717
R341 VTAIL.n60 VTAIL.n4 4.26717
R342 VTAIL.n198 VTAIL.n142 4.26717
R343 VTAIL.n169 VTAIL.n157 4.26717
R344 VTAIL.n130 VTAIL.n74 4.26717
R345 VTAIL.n101 VTAIL.n89 4.26717
R346 VTAIL.n238 VTAIL.n237 3.49141
R347 VTAIL.n263 VTAIL.n210 3.49141
R348 VTAIL.n34 VTAIL.n33 3.49141
R349 VTAIL.n59 VTAIL.n6 3.49141
R350 VTAIL.n197 VTAIL.n144 3.49141
R351 VTAIL.n173 VTAIL.n172 3.49141
R352 VTAIL.n129 VTAIL.n76 3.49141
R353 VTAIL.n105 VTAIL.n104 3.49141
R354 VTAIL.n241 VTAIL.n220 2.71565
R355 VTAIL.n260 VTAIL.n259 2.71565
R356 VTAIL.n37 VTAIL.n16 2.71565
R357 VTAIL.n56 VTAIL.n55 2.71565
R358 VTAIL.n194 VTAIL.n193 2.71565
R359 VTAIL.n176 VTAIL.n155 2.71565
R360 VTAIL.n126 VTAIL.n125 2.71565
R361 VTAIL.n108 VTAIL.n87 2.71565
R362 VTAIL.n0 VTAIL.t2 2.7025
R363 VTAIL.n0 VTAIL.t1 2.7025
R364 VTAIL.n68 VTAIL.t9 2.7025
R365 VTAIL.n68 VTAIL.t10 2.7025
R366 VTAIL.n138 VTAIL.t6 2.7025
R367 VTAIL.n138 VTAIL.t5 2.7025
R368 VTAIL.n70 VTAIL.t0 2.7025
R369 VTAIL.n70 VTAIL.t11 2.7025
R370 VTAIL.n163 VTAIL.n162 2.41282
R371 VTAIL.n95 VTAIL.n94 2.41282
R372 VTAIL.n228 VTAIL.n227 2.41282
R373 VTAIL.n24 VTAIL.n23 2.41282
R374 VTAIL.n242 VTAIL.n218 1.93989
R375 VTAIL.n256 VTAIL.n212 1.93989
R376 VTAIL.n38 VTAIL.n14 1.93989
R377 VTAIL.n52 VTAIL.n8 1.93989
R378 VTAIL.n190 VTAIL.n146 1.93989
R379 VTAIL.n177 VTAIL.n153 1.93989
R380 VTAIL.n122 VTAIL.n78 1.93989
R381 VTAIL.n109 VTAIL.n85 1.93989
R382 VTAIL.n137 VTAIL.n71 1.31947
R383 VTAIL.n205 VTAIL.n139 1.31947
R384 VTAIL.n69 VTAIL.n67 1.31947
R385 VTAIL.n247 VTAIL.n245 1.16414
R386 VTAIL.n255 VTAIL.n214 1.16414
R387 VTAIL.n43 VTAIL.n41 1.16414
R388 VTAIL.n51 VTAIL.n10 1.16414
R389 VTAIL.n189 VTAIL.n148 1.16414
R390 VTAIL.n181 VTAIL.n180 1.16414
R391 VTAIL.n121 VTAIL.n80 1.16414
R392 VTAIL.n113 VTAIL.n112 1.16414
R393 VTAIL.n139 VTAIL.n137 1.12981
R394 VTAIL.n67 VTAIL.n1 1.12981
R395 VTAIL VTAIL.n271 0.931535
R396 VTAIL VTAIL.n1 0.388431
R397 VTAIL.n246 VTAIL.n216 0.388379
R398 VTAIL.n252 VTAIL.n251 0.388379
R399 VTAIL.n42 VTAIL.n12 0.388379
R400 VTAIL.n48 VTAIL.n47 0.388379
R401 VTAIL.n186 VTAIL.n185 0.388379
R402 VTAIL.n152 VTAIL.n150 0.388379
R403 VTAIL.n118 VTAIL.n117 0.388379
R404 VTAIL.n84 VTAIL.n82 0.388379
R405 VTAIL.n228 VTAIL.n223 0.155672
R406 VTAIL.n235 VTAIL.n223 0.155672
R407 VTAIL.n236 VTAIL.n235 0.155672
R408 VTAIL.n236 VTAIL.n219 0.155672
R409 VTAIL.n243 VTAIL.n219 0.155672
R410 VTAIL.n244 VTAIL.n243 0.155672
R411 VTAIL.n244 VTAIL.n215 0.155672
R412 VTAIL.n253 VTAIL.n215 0.155672
R413 VTAIL.n254 VTAIL.n253 0.155672
R414 VTAIL.n254 VTAIL.n211 0.155672
R415 VTAIL.n261 VTAIL.n211 0.155672
R416 VTAIL.n262 VTAIL.n261 0.155672
R417 VTAIL.n262 VTAIL.n207 0.155672
R418 VTAIL.n269 VTAIL.n207 0.155672
R419 VTAIL.n24 VTAIL.n19 0.155672
R420 VTAIL.n31 VTAIL.n19 0.155672
R421 VTAIL.n32 VTAIL.n31 0.155672
R422 VTAIL.n32 VTAIL.n15 0.155672
R423 VTAIL.n39 VTAIL.n15 0.155672
R424 VTAIL.n40 VTAIL.n39 0.155672
R425 VTAIL.n40 VTAIL.n11 0.155672
R426 VTAIL.n49 VTAIL.n11 0.155672
R427 VTAIL.n50 VTAIL.n49 0.155672
R428 VTAIL.n50 VTAIL.n7 0.155672
R429 VTAIL.n57 VTAIL.n7 0.155672
R430 VTAIL.n58 VTAIL.n57 0.155672
R431 VTAIL.n58 VTAIL.n3 0.155672
R432 VTAIL.n65 VTAIL.n3 0.155672
R433 VTAIL.n203 VTAIL.n141 0.155672
R434 VTAIL.n196 VTAIL.n141 0.155672
R435 VTAIL.n196 VTAIL.n195 0.155672
R436 VTAIL.n195 VTAIL.n145 0.155672
R437 VTAIL.n188 VTAIL.n145 0.155672
R438 VTAIL.n188 VTAIL.n187 0.155672
R439 VTAIL.n187 VTAIL.n149 0.155672
R440 VTAIL.n179 VTAIL.n149 0.155672
R441 VTAIL.n179 VTAIL.n178 0.155672
R442 VTAIL.n178 VTAIL.n154 0.155672
R443 VTAIL.n171 VTAIL.n154 0.155672
R444 VTAIL.n171 VTAIL.n170 0.155672
R445 VTAIL.n170 VTAIL.n158 0.155672
R446 VTAIL.n163 VTAIL.n158 0.155672
R447 VTAIL.n135 VTAIL.n73 0.155672
R448 VTAIL.n128 VTAIL.n73 0.155672
R449 VTAIL.n128 VTAIL.n127 0.155672
R450 VTAIL.n127 VTAIL.n77 0.155672
R451 VTAIL.n120 VTAIL.n77 0.155672
R452 VTAIL.n120 VTAIL.n119 0.155672
R453 VTAIL.n119 VTAIL.n81 0.155672
R454 VTAIL.n111 VTAIL.n81 0.155672
R455 VTAIL.n111 VTAIL.n110 0.155672
R456 VTAIL.n110 VTAIL.n86 0.155672
R457 VTAIL.n103 VTAIL.n86 0.155672
R458 VTAIL.n103 VTAIL.n102 0.155672
R459 VTAIL.n102 VTAIL.n90 0.155672
R460 VTAIL.n95 VTAIL.n90 0.155672
R461 VDD1.n60 VDD1.n0 756.745
R462 VDD1.n125 VDD1.n65 756.745
R463 VDD1.n61 VDD1.n60 585
R464 VDD1.n59 VDD1.n58 585
R465 VDD1.n4 VDD1.n3 585
R466 VDD1.n53 VDD1.n52 585
R467 VDD1.n51 VDD1.n50 585
R468 VDD1.n8 VDD1.n7 585
R469 VDD1.n45 VDD1.n44 585
R470 VDD1.n43 VDD1.n10 585
R471 VDD1.n42 VDD1.n41 585
R472 VDD1.n13 VDD1.n11 585
R473 VDD1.n36 VDD1.n35 585
R474 VDD1.n34 VDD1.n33 585
R475 VDD1.n17 VDD1.n16 585
R476 VDD1.n28 VDD1.n27 585
R477 VDD1.n26 VDD1.n25 585
R478 VDD1.n21 VDD1.n20 585
R479 VDD1.n85 VDD1.n84 585
R480 VDD1.n90 VDD1.n89 585
R481 VDD1.n92 VDD1.n91 585
R482 VDD1.n81 VDD1.n80 585
R483 VDD1.n98 VDD1.n97 585
R484 VDD1.n100 VDD1.n99 585
R485 VDD1.n77 VDD1.n76 585
R486 VDD1.n107 VDD1.n106 585
R487 VDD1.n108 VDD1.n75 585
R488 VDD1.n110 VDD1.n109 585
R489 VDD1.n73 VDD1.n72 585
R490 VDD1.n116 VDD1.n115 585
R491 VDD1.n118 VDD1.n117 585
R492 VDD1.n69 VDD1.n68 585
R493 VDD1.n124 VDD1.n123 585
R494 VDD1.n126 VDD1.n125 585
R495 VDD1.n22 VDD1.t3 329.036
R496 VDD1.n86 VDD1.t4 329.036
R497 VDD1.n60 VDD1.n59 171.744
R498 VDD1.n59 VDD1.n3 171.744
R499 VDD1.n52 VDD1.n3 171.744
R500 VDD1.n52 VDD1.n51 171.744
R501 VDD1.n51 VDD1.n7 171.744
R502 VDD1.n44 VDD1.n7 171.744
R503 VDD1.n44 VDD1.n43 171.744
R504 VDD1.n43 VDD1.n42 171.744
R505 VDD1.n42 VDD1.n11 171.744
R506 VDD1.n35 VDD1.n11 171.744
R507 VDD1.n35 VDD1.n34 171.744
R508 VDD1.n34 VDD1.n16 171.744
R509 VDD1.n27 VDD1.n16 171.744
R510 VDD1.n27 VDD1.n26 171.744
R511 VDD1.n26 VDD1.n20 171.744
R512 VDD1.n90 VDD1.n84 171.744
R513 VDD1.n91 VDD1.n90 171.744
R514 VDD1.n91 VDD1.n80 171.744
R515 VDD1.n98 VDD1.n80 171.744
R516 VDD1.n99 VDD1.n98 171.744
R517 VDD1.n99 VDD1.n76 171.744
R518 VDD1.n107 VDD1.n76 171.744
R519 VDD1.n108 VDD1.n107 171.744
R520 VDD1.n109 VDD1.n108 171.744
R521 VDD1.n109 VDD1.n72 171.744
R522 VDD1.n116 VDD1.n72 171.744
R523 VDD1.n117 VDD1.n116 171.744
R524 VDD1.n117 VDD1.n68 171.744
R525 VDD1.n124 VDD1.n68 171.744
R526 VDD1.n125 VDD1.n124 171.744
R527 VDD1.t3 VDD1.n20 85.8723
R528 VDD1.t4 VDD1.n84 85.8723
R529 VDD1.n131 VDD1.n130 72.368
R530 VDD1.n133 VDD1.n132 72.0936
R531 VDD1 VDD1.n64 48.1661
R532 VDD1.n131 VDD1.n129 48.0526
R533 VDD1.n133 VDD1.n131 39.6151
R534 VDD1.n45 VDD1.n10 13.1884
R535 VDD1.n110 VDD1.n75 13.1884
R536 VDD1.n46 VDD1.n8 12.8005
R537 VDD1.n41 VDD1.n12 12.8005
R538 VDD1.n106 VDD1.n105 12.8005
R539 VDD1.n111 VDD1.n73 12.8005
R540 VDD1.n50 VDD1.n49 12.0247
R541 VDD1.n40 VDD1.n13 12.0247
R542 VDD1.n104 VDD1.n77 12.0247
R543 VDD1.n115 VDD1.n114 12.0247
R544 VDD1.n53 VDD1.n6 11.249
R545 VDD1.n37 VDD1.n36 11.249
R546 VDD1.n101 VDD1.n100 11.249
R547 VDD1.n118 VDD1.n71 11.249
R548 VDD1.n22 VDD1.n21 10.7239
R549 VDD1.n86 VDD1.n85 10.7239
R550 VDD1.n54 VDD1.n4 10.4732
R551 VDD1.n33 VDD1.n15 10.4732
R552 VDD1.n97 VDD1.n79 10.4732
R553 VDD1.n119 VDD1.n69 10.4732
R554 VDD1.n58 VDD1.n57 9.69747
R555 VDD1.n32 VDD1.n17 9.69747
R556 VDD1.n96 VDD1.n81 9.69747
R557 VDD1.n123 VDD1.n122 9.69747
R558 VDD1.n64 VDD1.n63 9.45567
R559 VDD1.n129 VDD1.n128 9.45567
R560 VDD1.n24 VDD1.n23 9.3005
R561 VDD1.n19 VDD1.n18 9.3005
R562 VDD1.n30 VDD1.n29 9.3005
R563 VDD1.n32 VDD1.n31 9.3005
R564 VDD1.n15 VDD1.n14 9.3005
R565 VDD1.n38 VDD1.n37 9.3005
R566 VDD1.n40 VDD1.n39 9.3005
R567 VDD1.n12 VDD1.n9 9.3005
R568 VDD1.n63 VDD1.n62 9.3005
R569 VDD1.n2 VDD1.n1 9.3005
R570 VDD1.n57 VDD1.n56 9.3005
R571 VDD1.n55 VDD1.n54 9.3005
R572 VDD1.n6 VDD1.n5 9.3005
R573 VDD1.n49 VDD1.n48 9.3005
R574 VDD1.n47 VDD1.n46 9.3005
R575 VDD1.n128 VDD1.n127 9.3005
R576 VDD1.n67 VDD1.n66 9.3005
R577 VDD1.n122 VDD1.n121 9.3005
R578 VDD1.n120 VDD1.n119 9.3005
R579 VDD1.n71 VDD1.n70 9.3005
R580 VDD1.n114 VDD1.n113 9.3005
R581 VDD1.n112 VDD1.n111 9.3005
R582 VDD1.n88 VDD1.n87 9.3005
R583 VDD1.n83 VDD1.n82 9.3005
R584 VDD1.n94 VDD1.n93 9.3005
R585 VDD1.n96 VDD1.n95 9.3005
R586 VDD1.n79 VDD1.n78 9.3005
R587 VDD1.n102 VDD1.n101 9.3005
R588 VDD1.n104 VDD1.n103 9.3005
R589 VDD1.n105 VDD1.n74 9.3005
R590 VDD1.n61 VDD1.n2 8.92171
R591 VDD1.n29 VDD1.n28 8.92171
R592 VDD1.n93 VDD1.n92 8.92171
R593 VDD1.n126 VDD1.n67 8.92171
R594 VDD1.n62 VDD1.n0 8.14595
R595 VDD1.n25 VDD1.n19 8.14595
R596 VDD1.n89 VDD1.n83 8.14595
R597 VDD1.n127 VDD1.n65 8.14595
R598 VDD1.n24 VDD1.n21 7.3702
R599 VDD1.n88 VDD1.n85 7.3702
R600 VDD1.n64 VDD1.n0 5.81868
R601 VDD1.n25 VDD1.n24 5.81868
R602 VDD1.n89 VDD1.n88 5.81868
R603 VDD1.n129 VDD1.n65 5.81868
R604 VDD1.n62 VDD1.n61 5.04292
R605 VDD1.n28 VDD1.n19 5.04292
R606 VDD1.n92 VDD1.n83 5.04292
R607 VDD1.n127 VDD1.n126 5.04292
R608 VDD1.n58 VDD1.n2 4.26717
R609 VDD1.n29 VDD1.n17 4.26717
R610 VDD1.n93 VDD1.n81 4.26717
R611 VDD1.n123 VDD1.n67 4.26717
R612 VDD1.n57 VDD1.n4 3.49141
R613 VDD1.n33 VDD1.n32 3.49141
R614 VDD1.n97 VDD1.n96 3.49141
R615 VDD1.n122 VDD1.n69 3.49141
R616 VDD1.n54 VDD1.n53 2.71565
R617 VDD1.n36 VDD1.n15 2.71565
R618 VDD1.n100 VDD1.n79 2.71565
R619 VDD1.n119 VDD1.n118 2.71565
R620 VDD1.n132 VDD1.t0 2.7025
R621 VDD1.n132 VDD1.t5 2.7025
R622 VDD1.n130 VDD1.t2 2.7025
R623 VDD1.n130 VDD1.t1 2.7025
R624 VDD1.n23 VDD1.n22 2.41282
R625 VDD1.n87 VDD1.n86 2.41282
R626 VDD1.n50 VDD1.n6 1.93989
R627 VDD1.n37 VDD1.n13 1.93989
R628 VDD1.n101 VDD1.n77 1.93989
R629 VDD1.n115 VDD1.n71 1.93989
R630 VDD1.n49 VDD1.n8 1.16414
R631 VDD1.n41 VDD1.n40 1.16414
R632 VDD1.n106 VDD1.n104 1.16414
R633 VDD1.n114 VDD1.n73 1.16414
R634 VDD1.n46 VDD1.n45 0.388379
R635 VDD1.n12 VDD1.n10 0.388379
R636 VDD1.n105 VDD1.n75 0.388379
R637 VDD1.n111 VDD1.n110 0.388379
R638 VDD1 VDD1.n133 0.272052
R639 VDD1.n63 VDD1.n1 0.155672
R640 VDD1.n56 VDD1.n1 0.155672
R641 VDD1.n56 VDD1.n55 0.155672
R642 VDD1.n55 VDD1.n5 0.155672
R643 VDD1.n48 VDD1.n5 0.155672
R644 VDD1.n48 VDD1.n47 0.155672
R645 VDD1.n47 VDD1.n9 0.155672
R646 VDD1.n39 VDD1.n9 0.155672
R647 VDD1.n39 VDD1.n38 0.155672
R648 VDD1.n38 VDD1.n14 0.155672
R649 VDD1.n31 VDD1.n14 0.155672
R650 VDD1.n31 VDD1.n30 0.155672
R651 VDD1.n30 VDD1.n18 0.155672
R652 VDD1.n23 VDD1.n18 0.155672
R653 VDD1.n87 VDD1.n82 0.155672
R654 VDD1.n94 VDD1.n82 0.155672
R655 VDD1.n95 VDD1.n94 0.155672
R656 VDD1.n95 VDD1.n78 0.155672
R657 VDD1.n102 VDD1.n78 0.155672
R658 VDD1.n103 VDD1.n102 0.155672
R659 VDD1.n103 VDD1.n74 0.155672
R660 VDD1.n112 VDD1.n74 0.155672
R661 VDD1.n113 VDD1.n112 0.155672
R662 VDD1.n113 VDD1.n70 0.155672
R663 VDD1.n120 VDD1.n70 0.155672
R664 VDD1.n121 VDD1.n120 0.155672
R665 VDD1.n121 VDD1.n66 0.155672
R666 VDD1.n128 VDD1.n66 0.155672
R667 B.n415 B.n414 585
R668 B.n416 B.n65 585
R669 B.n418 B.n417 585
R670 B.n419 B.n64 585
R671 B.n421 B.n420 585
R672 B.n422 B.n63 585
R673 B.n424 B.n423 585
R674 B.n425 B.n62 585
R675 B.n427 B.n426 585
R676 B.n428 B.n61 585
R677 B.n430 B.n429 585
R678 B.n431 B.n60 585
R679 B.n433 B.n432 585
R680 B.n434 B.n59 585
R681 B.n436 B.n435 585
R682 B.n437 B.n58 585
R683 B.n439 B.n438 585
R684 B.n440 B.n57 585
R685 B.n442 B.n441 585
R686 B.n443 B.n56 585
R687 B.n445 B.n444 585
R688 B.n446 B.n55 585
R689 B.n448 B.n447 585
R690 B.n449 B.n54 585
R691 B.n451 B.n450 585
R692 B.n452 B.n53 585
R693 B.n454 B.n453 585
R694 B.n455 B.n52 585
R695 B.n457 B.n456 585
R696 B.n458 B.n51 585
R697 B.n460 B.n459 585
R698 B.n461 B.n50 585
R699 B.n463 B.n462 585
R700 B.n464 B.n49 585
R701 B.n466 B.n465 585
R702 B.n467 B.n48 585
R703 B.n469 B.n468 585
R704 B.n470 B.n47 585
R705 B.n472 B.n471 585
R706 B.n473 B.n46 585
R707 B.n475 B.n474 585
R708 B.n476 B.n43 585
R709 B.n479 B.n478 585
R710 B.n480 B.n42 585
R711 B.n482 B.n481 585
R712 B.n483 B.n41 585
R713 B.n485 B.n484 585
R714 B.n486 B.n40 585
R715 B.n488 B.n487 585
R716 B.n489 B.n39 585
R717 B.n491 B.n490 585
R718 B.n493 B.n492 585
R719 B.n494 B.n35 585
R720 B.n496 B.n495 585
R721 B.n497 B.n34 585
R722 B.n499 B.n498 585
R723 B.n500 B.n33 585
R724 B.n502 B.n501 585
R725 B.n503 B.n32 585
R726 B.n505 B.n504 585
R727 B.n506 B.n31 585
R728 B.n508 B.n507 585
R729 B.n509 B.n30 585
R730 B.n511 B.n510 585
R731 B.n512 B.n29 585
R732 B.n514 B.n513 585
R733 B.n515 B.n28 585
R734 B.n517 B.n516 585
R735 B.n518 B.n27 585
R736 B.n520 B.n519 585
R737 B.n521 B.n26 585
R738 B.n523 B.n522 585
R739 B.n524 B.n25 585
R740 B.n526 B.n525 585
R741 B.n527 B.n24 585
R742 B.n529 B.n528 585
R743 B.n530 B.n23 585
R744 B.n532 B.n531 585
R745 B.n533 B.n22 585
R746 B.n535 B.n534 585
R747 B.n536 B.n21 585
R748 B.n538 B.n537 585
R749 B.n539 B.n20 585
R750 B.n541 B.n540 585
R751 B.n542 B.n19 585
R752 B.n544 B.n543 585
R753 B.n545 B.n18 585
R754 B.n547 B.n546 585
R755 B.n548 B.n17 585
R756 B.n550 B.n549 585
R757 B.n551 B.n16 585
R758 B.n553 B.n552 585
R759 B.n554 B.n15 585
R760 B.n413 B.n66 585
R761 B.n412 B.n411 585
R762 B.n410 B.n67 585
R763 B.n409 B.n408 585
R764 B.n407 B.n68 585
R765 B.n406 B.n405 585
R766 B.n404 B.n69 585
R767 B.n403 B.n402 585
R768 B.n401 B.n70 585
R769 B.n400 B.n399 585
R770 B.n398 B.n71 585
R771 B.n397 B.n396 585
R772 B.n395 B.n72 585
R773 B.n394 B.n393 585
R774 B.n392 B.n73 585
R775 B.n391 B.n390 585
R776 B.n389 B.n74 585
R777 B.n388 B.n387 585
R778 B.n386 B.n75 585
R779 B.n385 B.n384 585
R780 B.n383 B.n76 585
R781 B.n382 B.n381 585
R782 B.n380 B.n77 585
R783 B.n379 B.n378 585
R784 B.n377 B.n78 585
R785 B.n376 B.n375 585
R786 B.n374 B.n79 585
R787 B.n373 B.n372 585
R788 B.n371 B.n80 585
R789 B.n370 B.n369 585
R790 B.n368 B.n81 585
R791 B.n367 B.n366 585
R792 B.n365 B.n82 585
R793 B.n364 B.n363 585
R794 B.n362 B.n83 585
R795 B.n361 B.n360 585
R796 B.n359 B.n84 585
R797 B.n358 B.n357 585
R798 B.n356 B.n85 585
R799 B.n355 B.n354 585
R800 B.n353 B.n86 585
R801 B.n352 B.n351 585
R802 B.n350 B.n87 585
R803 B.n349 B.n348 585
R804 B.n347 B.n88 585
R805 B.n346 B.n345 585
R806 B.n344 B.n89 585
R807 B.n343 B.n342 585
R808 B.n341 B.n90 585
R809 B.n340 B.n339 585
R810 B.n338 B.n91 585
R811 B.n337 B.n336 585
R812 B.n335 B.n92 585
R813 B.n194 B.n143 585
R814 B.n196 B.n195 585
R815 B.n197 B.n142 585
R816 B.n199 B.n198 585
R817 B.n200 B.n141 585
R818 B.n202 B.n201 585
R819 B.n203 B.n140 585
R820 B.n205 B.n204 585
R821 B.n206 B.n139 585
R822 B.n208 B.n207 585
R823 B.n209 B.n138 585
R824 B.n211 B.n210 585
R825 B.n212 B.n137 585
R826 B.n214 B.n213 585
R827 B.n215 B.n136 585
R828 B.n217 B.n216 585
R829 B.n218 B.n135 585
R830 B.n220 B.n219 585
R831 B.n221 B.n134 585
R832 B.n223 B.n222 585
R833 B.n224 B.n133 585
R834 B.n226 B.n225 585
R835 B.n227 B.n132 585
R836 B.n229 B.n228 585
R837 B.n230 B.n131 585
R838 B.n232 B.n231 585
R839 B.n233 B.n130 585
R840 B.n235 B.n234 585
R841 B.n236 B.n129 585
R842 B.n238 B.n237 585
R843 B.n239 B.n128 585
R844 B.n241 B.n240 585
R845 B.n242 B.n127 585
R846 B.n244 B.n243 585
R847 B.n245 B.n126 585
R848 B.n247 B.n246 585
R849 B.n248 B.n125 585
R850 B.n250 B.n249 585
R851 B.n251 B.n124 585
R852 B.n253 B.n252 585
R853 B.n254 B.n123 585
R854 B.n256 B.n255 585
R855 B.n258 B.n257 585
R856 B.n259 B.n119 585
R857 B.n261 B.n260 585
R858 B.n262 B.n118 585
R859 B.n264 B.n263 585
R860 B.n265 B.n117 585
R861 B.n267 B.n266 585
R862 B.n268 B.n116 585
R863 B.n270 B.n269 585
R864 B.n272 B.n113 585
R865 B.n274 B.n273 585
R866 B.n275 B.n112 585
R867 B.n277 B.n276 585
R868 B.n278 B.n111 585
R869 B.n280 B.n279 585
R870 B.n281 B.n110 585
R871 B.n283 B.n282 585
R872 B.n284 B.n109 585
R873 B.n286 B.n285 585
R874 B.n287 B.n108 585
R875 B.n289 B.n288 585
R876 B.n290 B.n107 585
R877 B.n292 B.n291 585
R878 B.n293 B.n106 585
R879 B.n295 B.n294 585
R880 B.n296 B.n105 585
R881 B.n298 B.n297 585
R882 B.n299 B.n104 585
R883 B.n301 B.n300 585
R884 B.n302 B.n103 585
R885 B.n304 B.n303 585
R886 B.n305 B.n102 585
R887 B.n307 B.n306 585
R888 B.n308 B.n101 585
R889 B.n310 B.n309 585
R890 B.n311 B.n100 585
R891 B.n313 B.n312 585
R892 B.n314 B.n99 585
R893 B.n316 B.n315 585
R894 B.n317 B.n98 585
R895 B.n319 B.n318 585
R896 B.n320 B.n97 585
R897 B.n322 B.n321 585
R898 B.n323 B.n96 585
R899 B.n325 B.n324 585
R900 B.n326 B.n95 585
R901 B.n328 B.n327 585
R902 B.n329 B.n94 585
R903 B.n331 B.n330 585
R904 B.n332 B.n93 585
R905 B.n334 B.n333 585
R906 B.n193 B.n192 585
R907 B.n191 B.n144 585
R908 B.n190 B.n189 585
R909 B.n188 B.n145 585
R910 B.n187 B.n186 585
R911 B.n185 B.n146 585
R912 B.n184 B.n183 585
R913 B.n182 B.n147 585
R914 B.n181 B.n180 585
R915 B.n179 B.n148 585
R916 B.n178 B.n177 585
R917 B.n176 B.n149 585
R918 B.n175 B.n174 585
R919 B.n173 B.n150 585
R920 B.n172 B.n171 585
R921 B.n170 B.n151 585
R922 B.n169 B.n168 585
R923 B.n167 B.n152 585
R924 B.n166 B.n165 585
R925 B.n164 B.n153 585
R926 B.n163 B.n162 585
R927 B.n161 B.n154 585
R928 B.n160 B.n159 585
R929 B.n158 B.n155 585
R930 B.n157 B.n156 585
R931 B.n2 B.n0 585
R932 B.n593 B.n1 585
R933 B.n592 B.n591 585
R934 B.n590 B.n3 585
R935 B.n589 B.n588 585
R936 B.n587 B.n4 585
R937 B.n586 B.n585 585
R938 B.n584 B.n5 585
R939 B.n583 B.n582 585
R940 B.n581 B.n6 585
R941 B.n580 B.n579 585
R942 B.n578 B.n7 585
R943 B.n577 B.n576 585
R944 B.n575 B.n8 585
R945 B.n574 B.n573 585
R946 B.n572 B.n9 585
R947 B.n571 B.n570 585
R948 B.n569 B.n10 585
R949 B.n568 B.n567 585
R950 B.n566 B.n11 585
R951 B.n565 B.n564 585
R952 B.n563 B.n12 585
R953 B.n562 B.n561 585
R954 B.n560 B.n13 585
R955 B.n559 B.n558 585
R956 B.n557 B.n14 585
R957 B.n556 B.n555 585
R958 B.n595 B.n594 585
R959 B.n192 B.n143 516.524
R960 B.n556 B.n15 516.524
R961 B.n335 B.n334 516.524
R962 B.n414 B.n413 516.524
R963 B.n114 B.t9 445.719
R964 B.n120 B.t6 445.719
R965 B.n36 B.t0 445.719
R966 B.n44 B.t3 445.719
R967 B.n114 B.t11 405.784
R968 B.n44 B.t4 405.784
R969 B.n120 B.t8 405.784
R970 B.n36 B.t1 405.784
R971 B.n115 B.t10 376.111
R972 B.n45 B.t5 376.111
R973 B.n121 B.t7 376.111
R974 B.n37 B.t2 376.111
R975 B.n192 B.n191 163.367
R976 B.n191 B.n190 163.367
R977 B.n190 B.n145 163.367
R978 B.n186 B.n145 163.367
R979 B.n186 B.n185 163.367
R980 B.n185 B.n184 163.367
R981 B.n184 B.n147 163.367
R982 B.n180 B.n147 163.367
R983 B.n180 B.n179 163.367
R984 B.n179 B.n178 163.367
R985 B.n178 B.n149 163.367
R986 B.n174 B.n149 163.367
R987 B.n174 B.n173 163.367
R988 B.n173 B.n172 163.367
R989 B.n172 B.n151 163.367
R990 B.n168 B.n151 163.367
R991 B.n168 B.n167 163.367
R992 B.n167 B.n166 163.367
R993 B.n166 B.n153 163.367
R994 B.n162 B.n153 163.367
R995 B.n162 B.n161 163.367
R996 B.n161 B.n160 163.367
R997 B.n160 B.n155 163.367
R998 B.n156 B.n155 163.367
R999 B.n156 B.n2 163.367
R1000 B.n594 B.n2 163.367
R1001 B.n594 B.n593 163.367
R1002 B.n593 B.n592 163.367
R1003 B.n592 B.n3 163.367
R1004 B.n588 B.n3 163.367
R1005 B.n588 B.n587 163.367
R1006 B.n587 B.n586 163.367
R1007 B.n586 B.n5 163.367
R1008 B.n582 B.n5 163.367
R1009 B.n582 B.n581 163.367
R1010 B.n581 B.n580 163.367
R1011 B.n580 B.n7 163.367
R1012 B.n576 B.n7 163.367
R1013 B.n576 B.n575 163.367
R1014 B.n575 B.n574 163.367
R1015 B.n574 B.n9 163.367
R1016 B.n570 B.n9 163.367
R1017 B.n570 B.n569 163.367
R1018 B.n569 B.n568 163.367
R1019 B.n568 B.n11 163.367
R1020 B.n564 B.n11 163.367
R1021 B.n564 B.n563 163.367
R1022 B.n563 B.n562 163.367
R1023 B.n562 B.n13 163.367
R1024 B.n558 B.n13 163.367
R1025 B.n558 B.n557 163.367
R1026 B.n557 B.n556 163.367
R1027 B.n196 B.n143 163.367
R1028 B.n197 B.n196 163.367
R1029 B.n198 B.n197 163.367
R1030 B.n198 B.n141 163.367
R1031 B.n202 B.n141 163.367
R1032 B.n203 B.n202 163.367
R1033 B.n204 B.n203 163.367
R1034 B.n204 B.n139 163.367
R1035 B.n208 B.n139 163.367
R1036 B.n209 B.n208 163.367
R1037 B.n210 B.n209 163.367
R1038 B.n210 B.n137 163.367
R1039 B.n214 B.n137 163.367
R1040 B.n215 B.n214 163.367
R1041 B.n216 B.n215 163.367
R1042 B.n216 B.n135 163.367
R1043 B.n220 B.n135 163.367
R1044 B.n221 B.n220 163.367
R1045 B.n222 B.n221 163.367
R1046 B.n222 B.n133 163.367
R1047 B.n226 B.n133 163.367
R1048 B.n227 B.n226 163.367
R1049 B.n228 B.n227 163.367
R1050 B.n228 B.n131 163.367
R1051 B.n232 B.n131 163.367
R1052 B.n233 B.n232 163.367
R1053 B.n234 B.n233 163.367
R1054 B.n234 B.n129 163.367
R1055 B.n238 B.n129 163.367
R1056 B.n239 B.n238 163.367
R1057 B.n240 B.n239 163.367
R1058 B.n240 B.n127 163.367
R1059 B.n244 B.n127 163.367
R1060 B.n245 B.n244 163.367
R1061 B.n246 B.n245 163.367
R1062 B.n246 B.n125 163.367
R1063 B.n250 B.n125 163.367
R1064 B.n251 B.n250 163.367
R1065 B.n252 B.n251 163.367
R1066 B.n252 B.n123 163.367
R1067 B.n256 B.n123 163.367
R1068 B.n257 B.n256 163.367
R1069 B.n257 B.n119 163.367
R1070 B.n261 B.n119 163.367
R1071 B.n262 B.n261 163.367
R1072 B.n263 B.n262 163.367
R1073 B.n263 B.n117 163.367
R1074 B.n267 B.n117 163.367
R1075 B.n268 B.n267 163.367
R1076 B.n269 B.n268 163.367
R1077 B.n269 B.n113 163.367
R1078 B.n274 B.n113 163.367
R1079 B.n275 B.n274 163.367
R1080 B.n276 B.n275 163.367
R1081 B.n276 B.n111 163.367
R1082 B.n280 B.n111 163.367
R1083 B.n281 B.n280 163.367
R1084 B.n282 B.n281 163.367
R1085 B.n282 B.n109 163.367
R1086 B.n286 B.n109 163.367
R1087 B.n287 B.n286 163.367
R1088 B.n288 B.n287 163.367
R1089 B.n288 B.n107 163.367
R1090 B.n292 B.n107 163.367
R1091 B.n293 B.n292 163.367
R1092 B.n294 B.n293 163.367
R1093 B.n294 B.n105 163.367
R1094 B.n298 B.n105 163.367
R1095 B.n299 B.n298 163.367
R1096 B.n300 B.n299 163.367
R1097 B.n300 B.n103 163.367
R1098 B.n304 B.n103 163.367
R1099 B.n305 B.n304 163.367
R1100 B.n306 B.n305 163.367
R1101 B.n306 B.n101 163.367
R1102 B.n310 B.n101 163.367
R1103 B.n311 B.n310 163.367
R1104 B.n312 B.n311 163.367
R1105 B.n312 B.n99 163.367
R1106 B.n316 B.n99 163.367
R1107 B.n317 B.n316 163.367
R1108 B.n318 B.n317 163.367
R1109 B.n318 B.n97 163.367
R1110 B.n322 B.n97 163.367
R1111 B.n323 B.n322 163.367
R1112 B.n324 B.n323 163.367
R1113 B.n324 B.n95 163.367
R1114 B.n328 B.n95 163.367
R1115 B.n329 B.n328 163.367
R1116 B.n330 B.n329 163.367
R1117 B.n330 B.n93 163.367
R1118 B.n334 B.n93 163.367
R1119 B.n336 B.n335 163.367
R1120 B.n336 B.n91 163.367
R1121 B.n340 B.n91 163.367
R1122 B.n341 B.n340 163.367
R1123 B.n342 B.n341 163.367
R1124 B.n342 B.n89 163.367
R1125 B.n346 B.n89 163.367
R1126 B.n347 B.n346 163.367
R1127 B.n348 B.n347 163.367
R1128 B.n348 B.n87 163.367
R1129 B.n352 B.n87 163.367
R1130 B.n353 B.n352 163.367
R1131 B.n354 B.n353 163.367
R1132 B.n354 B.n85 163.367
R1133 B.n358 B.n85 163.367
R1134 B.n359 B.n358 163.367
R1135 B.n360 B.n359 163.367
R1136 B.n360 B.n83 163.367
R1137 B.n364 B.n83 163.367
R1138 B.n365 B.n364 163.367
R1139 B.n366 B.n365 163.367
R1140 B.n366 B.n81 163.367
R1141 B.n370 B.n81 163.367
R1142 B.n371 B.n370 163.367
R1143 B.n372 B.n371 163.367
R1144 B.n372 B.n79 163.367
R1145 B.n376 B.n79 163.367
R1146 B.n377 B.n376 163.367
R1147 B.n378 B.n377 163.367
R1148 B.n378 B.n77 163.367
R1149 B.n382 B.n77 163.367
R1150 B.n383 B.n382 163.367
R1151 B.n384 B.n383 163.367
R1152 B.n384 B.n75 163.367
R1153 B.n388 B.n75 163.367
R1154 B.n389 B.n388 163.367
R1155 B.n390 B.n389 163.367
R1156 B.n390 B.n73 163.367
R1157 B.n394 B.n73 163.367
R1158 B.n395 B.n394 163.367
R1159 B.n396 B.n395 163.367
R1160 B.n396 B.n71 163.367
R1161 B.n400 B.n71 163.367
R1162 B.n401 B.n400 163.367
R1163 B.n402 B.n401 163.367
R1164 B.n402 B.n69 163.367
R1165 B.n406 B.n69 163.367
R1166 B.n407 B.n406 163.367
R1167 B.n408 B.n407 163.367
R1168 B.n408 B.n67 163.367
R1169 B.n412 B.n67 163.367
R1170 B.n413 B.n412 163.367
R1171 B.n552 B.n15 163.367
R1172 B.n552 B.n551 163.367
R1173 B.n551 B.n550 163.367
R1174 B.n550 B.n17 163.367
R1175 B.n546 B.n17 163.367
R1176 B.n546 B.n545 163.367
R1177 B.n545 B.n544 163.367
R1178 B.n544 B.n19 163.367
R1179 B.n540 B.n19 163.367
R1180 B.n540 B.n539 163.367
R1181 B.n539 B.n538 163.367
R1182 B.n538 B.n21 163.367
R1183 B.n534 B.n21 163.367
R1184 B.n534 B.n533 163.367
R1185 B.n533 B.n532 163.367
R1186 B.n532 B.n23 163.367
R1187 B.n528 B.n23 163.367
R1188 B.n528 B.n527 163.367
R1189 B.n527 B.n526 163.367
R1190 B.n526 B.n25 163.367
R1191 B.n522 B.n25 163.367
R1192 B.n522 B.n521 163.367
R1193 B.n521 B.n520 163.367
R1194 B.n520 B.n27 163.367
R1195 B.n516 B.n27 163.367
R1196 B.n516 B.n515 163.367
R1197 B.n515 B.n514 163.367
R1198 B.n514 B.n29 163.367
R1199 B.n510 B.n29 163.367
R1200 B.n510 B.n509 163.367
R1201 B.n509 B.n508 163.367
R1202 B.n508 B.n31 163.367
R1203 B.n504 B.n31 163.367
R1204 B.n504 B.n503 163.367
R1205 B.n503 B.n502 163.367
R1206 B.n502 B.n33 163.367
R1207 B.n498 B.n33 163.367
R1208 B.n498 B.n497 163.367
R1209 B.n497 B.n496 163.367
R1210 B.n496 B.n35 163.367
R1211 B.n492 B.n35 163.367
R1212 B.n492 B.n491 163.367
R1213 B.n491 B.n39 163.367
R1214 B.n487 B.n39 163.367
R1215 B.n487 B.n486 163.367
R1216 B.n486 B.n485 163.367
R1217 B.n485 B.n41 163.367
R1218 B.n481 B.n41 163.367
R1219 B.n481 B.n480 163.367
R1220 B.n480 B.n479 163.367
R1221 B.n479 B.n43 163.367
R1222 B.n474 B.n43 163.367
R1223 B.n474 B.n473 163.367
R1224 B.n473 B.n472 163.367
R1225 B.n472 B.n47 163.367
R1226 B.n468 B.n47 163.367
R1227 B.n468 B.n467 163.367
R1228 B.n467 B.n466 163.367
R1229 B.n466 B.n49 163.367
R1230 B.n462 B.n49 163.367
R1231 B.n462 B.n461 163.367
R1232 B.n461 B.n460 163.367
R1233 B.n460 B.n51 163.367
R1234 B.n456 B.n51 163.367
R1235 B.n456 B.n455 163.367
R1236 B.n455 B.n454 163.367
R1237 B.n454 B.n53 163.367
R1238 B.n450 B.n53 163.367
R1239 B.n450 B.n449 163.367
R1240 B.n449 B.n448 163.367
R1241 B.n448 B.n55 163.367
R1242 B.n444 B.n55 163.367
R1243 B.n444 B.n443 163.367
R1244 B.n443 B.n442 163.367
R1245 B.n442 B.n57 163.367
R1246 B.n438 B.n57 163.367
R1247 B.n438 B.n437 163.367
R1248 B.n437 B.n436 163.367
R1249 B.n436 B.n59 163.367
R1250 B.n432 B.n59 163.367
R1251 B.n432 B.n431 163.367
R1252 B.n431 B.n430 163.367
R1253 B.n430 B.n61 163.367
R1254 B.n426 B.n61 163.367
R1255 B.n426 B.n425 163.367
R1256 B.n425 B.n424 163.367
R1257 B.n424 B.n63 163.367
R1258 B.n420 B.n63 163.367
R1259 B.n420 B.n419 163.367
R1260 B.n419 B.n418 163.367
R1261 B.n418 B.n65 163.367
R1262 B.n414 B.n65 163.367
R1263 B.n271 B.n115 59.5399
R1264 B.n122 B.n121 59.5399
R1265 B.n38 B.n37 59.5399
R1266 B.n477 B.n45 59.5399
R1267 B.n555 B.n554 33.5615
R1268 B.n415 B.n66 33.5615
R1269 B.n333 B.n92 33.5615
R1270 B.n194 B.n193 33.5615
R1271 B.n115 B.n114 29.6732
R1272 B.n121 B.n120 29.6732
R1273 B.n37 B.n36 29.6732
R1274 B.n45 B.n44 29.6732
R1275 B B.n595 18.0485
R1276 B.n554 B.n553 10.6151
R1277 B.n553 B.n16 10.6151
R1278 B.n549 B.n16 10.6151
R1279 B.n549 B.n548 10.6151
R1280 B.n548 B.n547 10.6151
R1281 B.n547 B.n18 10.6151
R1282 B.n543 B.n18 10.6151
R1283 B.n543 B.n542 10.6151
R1284 B.n542 B.n541 10.6151
R1285 B.n541 B.n20 10.6151
R1286 B.n537 B.n20 10.6151
R1287 B.n537 B.n536 10.6151
R1288 B.n536 B.n535 10.6151
R1289 B.n535 B.n22 10.6151
R1290 B.n531 B.n22 10.6151
R1291 B.n531 B.n530 10.6151
R1292 B.n530 B.n529 10.6151
R1293 B.n529 B.n24 10.6151
R1294 B.n525 B.n24 10.6151
R1295 B.n525 B.n524 10.6151
R1296 B.n524 B.n523 10.6151
R1297 B.n523 B.n26 10.6151
R1298 B.n519 B.n26 10.6151
R1299 B.n519 B.n518 10.6151
R1300 B.n518 B.n517 10.6151
R1301 B.n517 B.n28 10.6151
R1302 B.n513 B.n28 10.6151
R1303 B.n513 B.n512 10.6151
R1304 B.n512 B.n511 10.6151
R1305 B.n511 B.n30 10.6151
R1306 B.n507 B.n30 10.6151
R1307 B.n507 B.n506 10.6151
R1308 B.n506 B.n505 10.6151
R1309 B.n505 B.n32 10.6151
R1310 B.n501 B.n32 10.6151
R1311 B.n501 B.n500 10.6151
R1312 B.n500 B.n499 10.6151
R1313 B.n499 B.n34 10.6151
R1314 B.n495 B.n34 10.6151
R1315 B.n495 B.n494 10.6151
R1316 B.n494 B.n493 10.6151
R1317 B.n490 B.n489 10.6151
R1318 B.n489 B.n488 10.6151
R1319 B.n488 B.n40 10.6151
R1320 B.n484 B.n40 10.6151
R1321 B.n484 B.n483 10.6151
R1322 B.n483 B.n482 10.6151
R1323 B.n482 B.n42 10.6151
R1324 B.n478 B.n42 10.6151
R1325 B.n476 B.n475 10.6151
R1326 B.n475 B.n46 10.6151
R1327 B.n471 B.n46 10.6151
R1328 B.n471 B.n470 10.6151
R1329 B.n470 B.n469 10.6151
R1330 B.n469 B.n48 10.6151
R1331 B.n465 B.n48 10.6151
R1332 B.n465 B.n464 10.6151
R1333 B.n464 B.n463 10.6151
R1334 B.n463 B.n50 10.6151
R1335 B.n459 B.n50 10.6151
R1336 B.n459 B.n458 10.6151
R1337 B.n458 B.n457 10.6151
R1338 B.n457 B.n52 10.6151
R1339 B.n453 B.n52 10.6151
R1340 B.n453 B.n452 10.6151
R1341 B.n452 B.n451 10.6151
R1342 B.n451 B.n54 10.6151
R1343 B.n447 B.n54 10.6151
R1344 B.n447 B.n446 10.6151
R1345 B.n446 B.n445 10.6151
R1346 B.n445 B.n56 10.6151
R1347 B.n441 B.n56 10.6151
R1348 B.n441 B.n440 10.6151
R1349 B.n440 B.n439 10.6151
R1350 B.n439 B.n58 10.6151
R1351 B.n435 B.n58 10.6151
R1352 B.n435 B.n434 10.6151
R1353 B.n434 B.n433 10.6151
R1354 B.n433 B.n60 10.6151
R1355 B.n429 B.n60 10.6151
R1356 B.n429 B.n428 10.6151
R1357 B.n428 B.n427 10.6151
R1358 B.n427 B.n62 10.6151
R1359 B.n423 B.n62 10.6151
R1360 B.n423 B.n422 10.6151
R1361 B.n422 B.n421 10.6151
R1362 B.n421 B.n64 10.6151
R1363 B.n417 B.n64 10.6151
R1364 B.n417 B.n416 10.6151
R1365 B.n416 B.n415 10.6151
R1366 B.n337 B.n92 10.6151
R1367 B.n338 B.n337 10.6151
R1368 B.n339 B.n338 10.6151
R1369 B.n339 B.n90 10.6151
R1370 B.n343 B.n90 10.6151
R1371 B.n344 B.n343 10.6151
R1372 B.n345 B.n344 10.6151
R1373 B.n345 B.n88 10.6151
R1374 B.n349 B.n88 10.6151
R1375 B.n350 B.n349 10.6151
R1376 B.n351 B.n350 10.6151
R1377 B.n351 B.n86 10.6151
R1378 B.n355 B.n86 10.6151
R1379 B.n356 B.n355 10.6151
R1380 B.n357 B.n356 10.6151
R1381 B.n357 B.n84 10.6151
R1382 B.n361 B.n84 10.6151
R1383 B.n362 B.n361 10.6151
R1384 B.n363 B.n362 10.6151
R1385 B.n363 B.n82 10.6151
R1386 B.n367 B.n82 10.6151
R1387 B.n368 B.n367 10.6151
R1388 B.n369 B.n368 10.6151
R1389 B.n369 B.n80 10.6151
R1390 B.n373 B.n80 10.6151
R1391 B.n374 B.n373 10.6151
R1392 B.n375 B.n374 10.6151
R1393 B.n375 B.n78 10.6151
R1394 B.n379 B.n78 10.6151
R1395 B.n380 B.n379 10.6151
R1396 B.n381 B.n380 10.6151
R1397 B.n381 B.n76 10.6151
R1398 B.n385 B.n76 10.6151
R1399 B.n386 B.n385 10.6151
R1400 B.n387 B.n386 10.6151
R1401 B.n387 B.n74 10.6151
R1402 B.n391 B.n74 10.6151
R1403 B.n392 B.n391 10.6151
R1404 B.n393 B.n392 10.6151
R1405 B.n393 B.n72 10.6151
R1406 B.n397 B.n72 10.6151
R1407 B.n398 B.n397 10.6151
R1408 B.n399 B.n398 10.6151
R1409 B.n399 B.n70 10.6151
R1410 B.n403 B.n70 10.6151
R1411 B.n404 B.n403 10.6151
R1412 B.n405 B.n404 10.6151
R1413 B.n405 B.n68 10.6151
R1414 B.n409 B.n68 10.6151
R1415 B.n410 B.n409 10.6151
R1416 B.n411 B.n410 10.6151
R1417 B.n411 B.n66 10.6151
R1418 B.n195 B.n194 10.6151
R1419 B.n195 B.n142 10.6151
R1420 B.n199 B.n142 10.6151
R1421 B.n200 B.n199 10.6151
R1422 B.n201 B.n200 10.6151
R1423 B.n201 B.n140 10.6151
R1424 B.n205 B.n140 10.6151
R1425 B.n206 B.n205 10.6151
R1426 B.n207 B.n206 10.6151
R1427 B.n207 B.n138 10.6151
R1428 B.n211 B.n138 10.6151
R1429 B.n212 B.n211 10.6151
R1430 B.n213 B.n212 10.6151
R1431 B.n213 B.n136 10.6151
R1432 B.n217 B.n136 10.6151
R1433 B.n218 B.n217 10.6151
R1434 B.n219 B.n218 10.6151
R1435 B.n219 B.n134 10.6151
R1436 B.n223 B.n134 10.6151
R1437 B.n224 B.n223 10.6151
R1438 B.n225 B.n224 10.6151
R1439 B.n225 B.n132 10.6151
R1440 B.n229 B.n132 10.6151
R1441 B.n230 B.n229 10.6151
R1442 B.n231 B.n230 10.6151
R1443 B.n231 B.n130 10.6151
R1444 B.n235 B.n130 10.6151
R1445 B.n236 B.n235 10.6151
R1446 B.n237 B.n236 10.6151
R1447 B.n237 B.n128 10.6151
R1448 B.n241 B.n128 10.6151
R1449 B.n242 B.n241 10.6151
R1450 B.n243 B.n242 10.6151
R1451 B.n243 B.n126 10.6151
R1452 B.n247 B.n126 10.6151
R1453 B.n248 B.n247 10.6151
R1454 B.n249 B.n248 10.6151
R1455 B.n249 B.n124 10.6151
R1456 B.n253 B.n124 10.6151
R1457 B.n254 B.n253 10.6151
R1458 B.n255 B.n254 10.6151
R1459 B.n259 B.n258 10.6151
R1460 B.n260 B.n259 10.6151
R1461 B.n260 B.n118 10.6151
R1462 B.n264 B.n118 10.6151
R1463 B.n265 B.n264 10.6151
R1464 B.n266 B.n265 10.6151
R1465 B.n266 B.n116 10.6151
R1466 B.n270 B.n116 10.6151
R1467 B.n273 B.n272 10.6151
R1468 B.n273 B.n112 10.6151
R1469 B.n277 B.n112 10.6151
R1470 B.n278 B.n277 10.6151
R1471 B.n279 B.n278 10.6151
R1472 B.n279 B.n110 10.6151
R1473 B.n283 B.n110 10.6151
R1474 B.n284 B.n283 10.6151
R1475 B.n285 B.n284 10.6151
R1476 B.n285 B.n108 10.6151
R1477 B.n289 B.n108 10.6151
R1478 B.n290 B.n289 10.6151
R1479 B.n291 B.n290 10.6151
R1480 B.n291 B.n106 10.6151
R1481 B.n295 B.n106 10.6151
R1482 B.n296 B.n295 10.6151
R1483 B.n297 B.n296 10.6151
R1484 B.n297 B.n104 10.6151
R1485 B.n301 B.n104 10.6151
R1486 B.n302 B.n301 10.6151
R1487 B.n303 B.n302 10.6151
R1488 B.n303 B.n102 10.6151
R1489 B.n307 B.n102 10.6151
R1490 B.n308 B.n307 10.6151
R1491 B.n309 B.n308 10.6151
R1492 B.n309 B.n100 10.6151
R1493 B.n313 B.n100 10.6151
R1494 B.n314 B.n313 10.6151
R1495 B.n315 B.n314 10.6151
R1496 B.n315 B.n98 10.6151
R1497 B.n319 B.n98 10.6151
R1498 B.n320 B.n319 10.6151
R1499 B.n321 B.n320 10.6151
R1500 B.n321 B.n96 10.6151
R1501 B.n325 B.n96 10.6151
R1502 B.n326 B.n325 10.6151
R1503 B.n327 B.n326 10.6151
R1504 B.n327 B.n94 10.6151
R1505 B.n331 B.n94 10.6151
R1506 B.n332 B.n331 10.6151
R1507 B.n333 B.n332 10.6151
R1508 B.n193 B.n144 10.6151
R1509 B.n189 B.n144 10.6151
R1510 B.n189 B.n188 10.6151
R1511 B.n188 B.n187 10.6151
R1512 B.n187 B.n146 10.6151
R1513 B.n183 B.n146 10.6151
R1514 B.n183 B.n182 10.6151
R1515 B.n182 B.n181 10.6151
R1516 B.n181 B.n148 10.6151
R1517 B.n177 B.n148 10.6151
R1518 B.n177 B.n176 10.6151
R1519 B.n176 B.n175 10.6151
R1520 B.n175 B.n150 10.6151
R1521 B.n171 B.n150 10.6151
R1522 B.n171 B.n170 10.6151
R1523 B.n170 B.n169 10.6151
R1524 B.n169 B.n152 10.6151
R1525 B.n165 B.n152 10.6151
R1526 B.n165 B.n164 10.6151
R1527 B.n164 B.n163 10.6151
R1528 B.n163 B.n154 10.6151
R1529 B.n159 B.n154 10.6151
R1530 B.n159 B.n158 10.6151
R1531 B.n158 B.n157 10.6151
R1532 B.n157 B.n0 10.6151
R1533 B.n591 B.n1 10.6151
R1534 B.n591 B.n590 10.6151
R1535 B.n590 B.n589 10.6151
R1536 B.n589 B.n4 10.6151
R1537 B.n585 B.n4 10.6151
R1538 B.n585 B.n584 10.6151
R1539 B.n584 B.n583 10.6151
R1540 B.n583 B.n6 10.6151
R1541 B.n579 B.n6 10.6151
R1542 B.n579 B.n578 10.6151
R1543 B.n578 B.n577 10.6151
R1544 B.n577 B.n8 10.6151
R1545 B.n573 B.n8 10.6151
R1546 B.n573 B.n572 10.6151
R1547 B.n572 B.n571 10.6151
R1548 B.n571 B.n10 10.6151
R1549 B.n567 B.n10 10.6151
R1550 B.n567 B.n566 10.6151
R1551 B.n566 B.n565 10.6151
R1552 B.n565 B.n12 10.6151
R1553 B.n561 B.n12 10.6151
R1554 B.n561 B.n560 10.6151
R1555 B.n560 B.n559 10.6151
R1556 B.n559 B.n14 10.6151
R1557 B.n555 B.n14 10.6151
R1558 B.n490 B.n38 6.5566
R1559 B.n478 B.n477 6.5566
R1560 B.n258 B.n122 6.5566
R1561 B.n271 B.n270 6.5566
R1562 B.n493 B.n38 4.05904
R1563 B.n477 B.n476 4.05904
R1564 B.n255 B.n122 4.05904
R1565 B.n272 B.n271 4.05904
R1566 B.n595 B.n0 2.81026
R1567 B.n595 B.n1 2.81026
R1568 VN.n3 VN.t5 272.635
R1569 VN.n13 VN.t0 272.635
R1570 VN.n2 VN.t4 241.602
R1571 VN.n8 VN.t1 241.602
R1572 VN.n12 VN.t2 241.602
R1573 VN.n18 VN.t3 241.602
R1574 VN.n9 VN.n8 172.065
R1575 VN.n19 VN.n18 172.065
R1576 VN.n17 VN.n10 161.3
R1577 VN.n16 VN.n15 161.3
R1578 VN.n14 VN.n11 161.3
R1579 VN.n7 VN.n0 161.3
R1580 VN.n6 VN.n5 161.3
R1581 VN.n4 VN.n1 161.3
R1582 VN.n3 VN.n2 51.3222
R1583 VN.n13 VN.n12 51.3222
R1584 VN VN.n19 43.4986
R1585 VN.n7 VN.n6 41.9503
R1586 VN.n17 VN.n16 41.9503
R1587 VN.n6 VN.n1 39.0365
R1588 VN.n16 VN.n11 39.0365
R1589 VN.n14 VN.n13 26.7683
R1590 VN.n4 VN.n3 26.7683
R1591 VN.n8 VN.n7 13.702
R1592 VN.n18 VN.n17 13.702
R1593 VN.n2 VN.n1 12.234
R1594 VN.n12 VN.n11 12.234
R1595 VN.n19 VN.n10 0.189894
R1596 VN.n15 VN.n10 0.189894
R1597 VN.n15 VN.n14 0.189894
R1598 VN.n5 VN.n4 0.189894
R1599 VN.n5 VN.n0 0.189894
R1600 VN.n9 VN.n0 0.189894
R1601 VN VN.n9 0.0516364
R1602 VDD2.n127 VDD2.n67 756.745
R1603 VDD2.n60 VDD2.n0 756.745
R1604 VDD2.n128 VDD2.n127 585
R1605 VDD2.n126 VDD2.n125 585
R1606 VDD2.n71 VDD2.n70 585
R1607 VDD2.n120 VDD2.n119 585
R1608 VDD2.n118 VDD2.n117 585
R1609 VDD2.n75 VDD2.n74 585
R1610 VDD2.n112 VDD2.n111 585
R1611 VDD2.n110 VDD2.n77 585
R1612 VDD2.n109 VDD2.n108 585
R1613 VDD2.n80 VDD2.n78 585
R1614 VDD2.n103 VDD2.n102 585
R1615 VDD2.n101 VDD2.n100 585
R1616 VDD2.n84 VDD2.n83 585
R1617 VDD2.n95 VDD2.n94 585
R1618 VDD2.n93 VDD2.n92 585
R1619 VDD2.n88 VDD2.n87 585
R1620 VDD2.n20 VDD2.n19 585
R1621 VDD2.n25 VDD2.n24 585
R1622 VDD2.n27 VDD2.n26 585
R1623 VDD2.n16 VDD2.n15 585
R1624 VDD2.n33 VDD2.n32 585
R1625 VDD2.n35 VDD2.n34 585
R1626 VDD2.n12 VDD2.n11 585
R1627 VDD2.n42 VDD2.n41 585
R1628 VDD2.n43 VDD2.n10 585
R1629 VDD2.n45 VDD2.n44 585
R1630 VDD2.n8 VDD2.n7 585
R1631 VDD2.n51 VDD2.n50 585
R1632 VDD2.n53 VDD2.n52 585
R1633 VDD2.n4 VDD2.n3 585
R1634 VDD2.n59 VDD2.n58 585
R1635 VDD2.n61 VDD2.n60 585
R1636 VDD2.n89 VDD2.t2 329.036
R1637 VDD2.n21 VDD2.t0 329.036
R1638 VDD2.n127 VDD2.n126 171.744
R1639 VDD2.n126 VDD2.n70 171.744
R1640 VDD2.n119 VDD2.n70 171.744
R1641 VDD2.n119 VDD2.n118 171.744
R1642 VDD2.n118 VDD2.n74 171.744
R1643 VDD2.n111 VDD2.n74 171.744
R1644 VDD2.n111 VDD2.n110 171.744
R1645 VDD2.n110 VDD2.n109 171.744
R1646 VDD2.n109 VDD2.n78 171.744
R1647 VDD2.n102 VDD2.n78 171.744
R1648 VDD2.n102 VDD2.n101 171.744
R1649 VDD2.n101 VDD2.n83 171.744
R1650 VDD2.n94 VDD2.n83 171.744
R1651 VDD2.n94 VDD2.n93 171.744
R1652 VDD2.n93 VDD2.n87 171.744
R1653 VDD2.n25 VDD2.n19 171.744
R1654 VDD2.n26 VDD2.n25 171.744
R1655 VDD2.n26 VDD2.n15 171.744
R1656 VDD2.n33 VDD2.n15 171.744
R1657 VDD2.n34 VDD2.n33 171.744
R1658 VDD2.n34 VDD2.n11 171.744
R1659 VDD2.n42 VDD2.n11 171.744
R1660 VDD2.n43 VDD2.n42 171.744
R1661 VDD2.n44 VDD2.n43 171.744
R1662 VDD2.n44 VDD2.n7 171.744
R1663 VDD2.n51 VDD2.n7 171.744
R1664 VDD2.n52 VDD2.n51 171.744
R1665 VDD2.n52 VDD2.n3 171.744
R1666 VDD2.n59 VDD2.n3 171.744
R1667 VDD2.n60 VDD2.n59 171.744
R1668 VDD2.t2 VDD2.n87 85.8723
R1669 VDD2.t0 VDD2.n19 85.8723
R1670 VDD2.n66 VDD2.n65 72.368
R1671 VDD2 VDD2.n133 72.3651
R1672 VDD2.n66 VDD2.n64 48.0526
R1673 VDD2.n132 VDD2.n131 47.1187
R1674 VDD2.n132 VDD2.n66 38.3726
R1675 VDD2.n112 VDD2.n77 13.1884
R1676 VDD2.n45 VDD2.n10 13.1884
R1677 VDD2.n113 VDD2.n75 12.8005
R1678 VDD2.n108 VDD2.n79 12.8005
R1679 VDD2.n41 VDD2.n40 12.8005
R1680 VDD2.n46 VDD2.n8 12.8005
R1681 VDD2.n117 VDD2.n116 12.0247
R1682 VDD2.n107 VDD2.n80 12.0247
R1683 VDD2.n39 VDD2.n12 12.0247
R1684 VDD2.n50 VDD2.n49 12.0247
R1685 VDD2.n120 VDD2.n73 11.249
R1686 VDD2.n104 VDD2.n103 11.249
R1687 VDD2.n36 VDD2.n35 11.249
R1688 VDD2.n53 VDD2.n6 11.249
R1689 VDD2.n89 VDD2.n88 10.7239
R1690 VDD2.n21 VDD2.n20 10.7239
R1691 VDD2.n121 VDD2.n71 10.4732
R1692 VDD2.n100 VDD2.n82 10.4732
R1693 VDD2.n32 VDD2.n14 10.4732
R1694 VDD2.n54 VDD2.n4 10.4732
R1695 VDD2.n125 VDD2.n124 9.69747
R1696 VDD2.n99 VDD2.n84 9.69747
R1697 VDD2.n31 VDD2.n16 9.69747
R1698 VDD2.n58 VDD2.n57 9.69747
R1699 VDD2.n131 VDD2.n130 9.45567
R1700 VDD2.n64 VDD2.n63 9.45567
R1701 VDD2.n91 VDD2.n90 9.3005
R1702 VDD2.n86 VDD2.n85 9.3005
R1703 VDD2.n97 VDD2.n96 9.3005
R1704 VDD2.n99 VDD2.n98 9.3005
R1705 VDD2.n82 VDD2.n81 9.3005
R1706 VDD2.n105 VDD2.n104 9.3005
R1707 VDD2.n107 VDD2.n106 9.3005
R1708 VDD2.n79 VDD2.n76 9.3005
R1709 VDD2.n130 VDD2.n129 9.3005
R1710 VDD2.n69 VDD2.n68 9.3005
R1711 VDD2.n124 VDD2.n123 9.3005
R1712 VDD2.n122 VDD2.n121 9.3005
R1713 VDD2.n73 VDD2.n72 9.3005
R1714 VDD2.n116 VDD2.n115 9.3005
R1715 VDD2.n114 VDD2.n113 9.3005
R1716 VDD2.n63 VDD2.n62 9.3005
R1717 VDD2.n2 VDD2.n1 9.3005
R1718 VDD2.n57 VDD2.n56 9.3005
R1719 VDD2.n55 VDD2.n54 9.3005
R1720 VDD2.n6 VDD2.n5 9.3005
R1721 VDD2.n49 VDD2.n48 9.3005
R1722 VDD2.n47 VDD2.n46 9.3005
R1723 VDD2.n23 VDD2.n22 9.3005
R1724 VDD2.n18 VDD2.n17 9.3005
R1725 VDD2.n29 VDD2.n28 9.3005
R1726 VDD2.n31 VDD2.n30 9.3005
R1727 VDD2.n14 VDD2.n13 9.3005
R1728 VDD2.n37 VDD2.n36 9.3005
R1729 VDD2.n39 VDD2.n38 9.3005
R1730 VDD2.n40 VDD2.n9 9.3005
R1731 VDD2.n128 VDD2.n69 8.92171
R1732 VDD2.n96 VDD2.n95 8.92171
R1733 VDD2.n28 VDD2.n27 8.92171
R1734 VDD2.n61 VDD2.n2 8.92171
R1735 VDD2.n129 VDD2.n67 8.14595
R1736 VDD2.n92 VDD2.n86 8.14595
R1737 VDD2.n24 VDD2.n18 8.14595
R1738 VDD2.n62 VDD2.n0 8.14595
R1739 VDD2.n91 VDD2.n88 7.3702
R1740 VDD2.n23 VDD2.n20 7.3702
R1741 VDD2.n131 VDD2.n67 5.81868
R1742 VDD2.n92 VDD2.n91 5.81868
R1743 VDD2.n24 VDD2.n23 5.81868
R1744 VDD2.n64 VDD2.n0 5.81868
R1745 VDD2.n129 VDD2.n128 5.04292
R1746 VDD2.n95 VDD2.n86 5.04292
R1747 VDD2.n27 VDD2.n18 5.04292
R1748 VDD2.n62 VDD2.n61 5.04292
R1749 VDD2.n125 VDD2.n69 4.26717
R1750 VDD2.n96 VDD2.n84 4.26717
R1751 VDD2.n28 VDD2.n16 4.26717
R1752 VDD2.n58 VDD2.n2 4.26717
R1753 VDD2.n124 VDD2.n71 3.49141
R1754 VDD2.n100 VDD2.n99 3.49141
R1755 VDD2.n32 VDD2.n31 3.49141
R1756 VDD2.n57 VDD2.n4 3.49141
R1757 VDD2.n121 VDD2.n120 2.71565
R1758 VDD2.n103 VDD2.n82 2.71565
R1759 VDD2.n35 VDD2.n14 2.71565
R1760 VDD2.n54 VDD2.n53 2.71565
R1761 VDD2.n133 VDD2.t3 2.7025
R1762 VDD2.n133 VDD2.t5 2.7025
R1763 VDD2.n65 VDD2.t1 2.7025
R1764 VDD2.n65 VDD2.t4 2.7025
R1765 VDD2.n90 VDD2.n89 2.41282
R1766 VDD2.n22 VDD2.n21 2.41282
R1767 VDD2.n117 VDD2.n73 1.93989
R1768 VDD2.n104 VDD2.n80 1.93989
R1769 VDD2.n36 VDD2.n12 1.93989
R1770 VDD2.n50 VDD2.n6 1.93989
R1771 VDD2.n116 VDD2.n75 1.16414
R1772 VDD2.n108 VDD2.n107 1.16414
R1773 VDD2.n41 VDD2.n39 1.16414
R1774 VDD2.n49 VDD2.n8 1.16414
R1775 VDD2 VDD2.n132 1.04791
R1776 VDD2.n113 VDD2.n112 0.388379
R1777 VDD2.n79 VDD2.n77 0.388379
R1778 VDD2.n40 VDD2.n10 0.388379
R1779 VDD2.n46 VDD2.n45 0.388379
R1780 VDD2.n130 VDD2.n68 0.155672
R1781 VDD2.n123 VDD2.n68 0.155672
R1782 VDD2.n123 VDD2.n122 0.155672
R1783 VDD2.n122 VDD2.n72 0.155672
R1784 VDD2.n115 VDD2.n72 0.155672
R1785 VDD2.n115 VDD2.n114 0.155672
R1786 VDD2.n114 VDD2.n76 0.155672
R1787 VDD2.n106 VDD2.n76 0.155672
R1788 VDD2.n106 VDD2.n105 0.155672
R1789 VDD2.n105 VDD2.n81 0.155672
R1790 VDD2.n98 VDD2.n81 0.155672
R1791 VDD2.n98 VDD2.n97 0.155672
R1792 VDD2.n97 VDD2.n85 0.155672
R1793 VDD2.n90 VDD2.n85 0.155672
R1794 VDD2.n22 VDD2.n17 0.155672
R1795 VDD2.n29 VDD2.n17 0.155672
R1796 VDD2.n30 VDD2.n29 0.155672
R1797 VDD2.n30 VDD2.n13 0.155672
R1798 VDD2.n37 VDD2.n13 0.155672
R1799 VDD2.n38 VDD2.n37 0.155672
R1800 VDD2.n38 VDD2.n9 0.155672
R1801 VDD2.n47 VDD2.n9 0.155672
R1802 VDD2.n48 VDD2.n47 0.155672
R1803 VDD2.n48 VDD2.n5 0.155672
R1804 VDD2.n55 VDD2.n5 0.155672
R1805 VDD2.n56 VDD2.n55 0.155672
R1806 VDD2.n56 VDD2.n1 0.155672
R1807 VDD2.n63 VDD2.n1 0.155672
C0 VDD1 VP 5.6618f
C1 VTAIL VDD1 8.39307f
C2 VTAIL VP 5.31953f
C3 w_n2194_n3374# VDD2 1.98253f
C4 VDD2 B 1.75201f
C5 VDD2 VN 5.47475f
C6 w_n2194_n3374# B 7.751161f
C7 w_n2194_n3374# VN 3.82804f
C8 VDD1 VDD2 0.893151f
C9 B VN 0.871253f
C10 VDD2 VP 0.339618f
C11 w_n2194_n3374# VDD1 1.94264f
C12 VTAIL VDD2 8.432111f
C13 w_n2194_n3374# VP 4.10779f
C14 VDD1 B 1.71127f
C15 B VP 1.33128f
C16 w_n2194_n3374# VTAIL 2.89547f
C17 VDD1 VN 0.148614f
C18 VTAIL B 3.02505f
C19 VN VP 5.57378f
C20 VTAIL VN 5.30505f
C21 VDD2 VSUBS 1.386734f
C22 VDD1 VSUBS 1.280644f
C23 VTAIL VSUBS 0.896828f
C24 VN VSUBS 4.6667f
C25 VP VSUBS 1.842733f
C26 B VSUBS 3.256646f
C27 w_n2194_n3374# VSUBS 91.1212f
C28 VDD2.n0 VSUBS 0.023283f
C29 VDD2.n1 VSUBS 0.022038f
C30 VDD2.n2 VSUBS 0.011843f
C31 VDD2.n3 VSUBS 0.027991f
C32 VDD2.n4 VSUBS 0.012539f
C33 VDD2.n5 VSUBS 0.022038f
C34 VDD2.n6 VSUBS 0.011843f
C35 VDD2.n7 VSUBS 0.027991f
C36 VDD2.n8 VSUBS 0.012539f
C37 VDD2.n9 VSUBS 0.022038f
C38 VDD2.n10 VSUBS 0.012191f
C39 VDD2.n11 VSUBS 0.027991f
C40 VDD2.n12 VSUBS 0.012539f
C41 VDD2.n13 VSUBS 0.022038f
C42 VDD2.n14 VSUBS 0.011843f
C43 VDD2.n15 VSUBS 0.027991f
C44 VDD2.n16 VSUBS 0.012539f
C45 VDD2.n17 VSUBS 0.022038f
C46 VDD2.n18 VSUBS 0.011843f
C47 VDD2.n19 VSUBS 0.020993f
C48 VDD2.n20 VSUBS 0.021057f
C49 VDD2.t0 VSUBS 0.06032f
C50 VDD2.n21 VSUBS 0.173864f
C51 VDD2.n22 VSUBS 1.08572f
C52 VDD2.n23 VSUBS 0.011843f
C53 VDD2.n24 VSUBS 0.012539f
C54 VDD2.n25 VSUBS 0.027991f
C55 VDD2.n26 VSUBS 0.027991f
C56 VDD2.n27 VSUBS 0.012539f
C57 VDD2.n28 VSUBS 0.011843f
C58 VDD2.n29 VSUBS 0.022038f
C59 VDD2.n30 VSUBS 0.022038f
C60 VDD2.n31 VSUBS 0.011843f
C61 VDD2.n32 VSUBS 0.012539f
C62 VDD2.n33 VSUBS 0.027991f
C63 VDD2.n34 VSUBS 0.027991f
C64 VDD2.n35 VSUBS 0.012539f
C65 VDD2.n36 VSUBS 0.011843f
C66 VDD2.n37 VSUBS 0.022038f
C67 VDD2.n38 VSUBS 0.022038f
C68 VDD2.n39 VSUBS 0.011843f
C69 VDD2.n40 VSUBS 0.011843f
C70 VDD2.n41 VSUBS 0.012539f
C71 VDD2.n42 VSUBS 0.027991f
C72 VDD2.n43 VSUBS 0.027991f
C73 VDD2.n44 VSUBS 0.027991f
C74 VDD2.n45 VSUBS 0.012191f
C75 VDD2.n46 VSUBS 0.011843f
C76 VDD2.n47 VSUBS 0.022038f
C77 VDD2.n48 VSUBS 0.022038f
C78 VDD2.n49 VSUBS 0.011843f
C79 VDD2.n50 VSUBS 0.012539f
C80 VDD2.n51 VSUBS 0.027991f
C81 VDD2.n52 VSUBS 0.027991f
C82 VDD2.n53 VSUBS 0.012539f
C83 VDD2.n54 VSUBS 0.011843f
C84 VDD2.n55 VSUBS 0.022038f
C85 VDD2.n56 VSUBS 0.022038f
C86 VDD2.n57 VSUBS 0.011843f
C87 VDD2.n58 VSUBS 0.012539f
C88 VDD2.n59 VSUBS 0.027991f
C89 VDD2.n60 VSUBS 0.064586f
C90 VDD2.n61 VSUBS 0.012539f
C91 VDD2.n62 VSUBS 0.011843f
C92 VDD2.n63 VSUBS 0.048231f
C93 VDD2.n64 VSUBS 0.049587f
C94 VDD2.t1 VSUBS 0.209507f
C95 VDD2.t4 VSUBS 0.209507f
C96 VDD2.n65 VSUBS 1.63153f
C97 VDD2.n66 VSUBS 2.06323f
C98 VDD2.n67 VSUBS 0.023283f
C99 VDD2.n68 VSUBS 0.022038f
C100 VDD2.n69 VSUBS 0.011843f
C101 VDD2.n70 VSUBS 0.027991f
C102 VDD2.n71 VSUBS 0.012539f
C103 VDD2.n72 VSUBS 0.022038f
C104 VDD2.n73 VSUBS 0.011843f
C105 VDD2.n74 VSUBS 0.027991f
C106 VDD2.n75 VSUBS 0.012539f
C107 VDD2.n76 VSUBS 0.022038f
C108 VDD2.n77 VSUBS 0.012191f
C109 VDD2.n78 VSUBS 0.027991f
C110 VDD2.n79 VSUBS 0.011843f
C111 VDD2.n80 VSUBS 0.012539f
C112 VDD2.n81 VSUBS 0.022038f
C113 VDD2.n82 VSUBS 0.011843f
C114 VDD2.n83 VSUBS 0.027991f
C115 VDD2.n84 VSUBS 0.012539f
C116 VDD2.n85 VSUBS 0.022038f
C117 VDD2.n86 VSUBS 0.011843f
C118 VDD2.n87 VSUBS 0.020993f
C119 VDD2.n88 VSUBS 0.021057f
C120 VDD2.t2 VSUBS 0.06032f
C121 VDD2.n89 VSUBS 0.173864f
C122 VDD2.n90 VSUBS 1.08572f
C123 VDD2.n91 VSUBS 0.011843f
C124 VDD2.n92 VSUBS 0.012539f
C125 VDD2.n93 VSUBS 0.027991f
C126 VDD2.n94 VSUBS 0.027991f
C127 VDD2.n95 VSUBS 0.012539f
C128 VDD2.n96 VSUBS 0.011843f
C129 VDD2.n97 VSUBS 0.022038f
C130 VDD2.n98 VSUBS 0.022038f
C131 VDD2.n99 VSUBS 0.011843f
C132 VDD2.n100 VSUBS 0.012539f
C133 VDD2.n101 VSUBS 0.027991f
C134 VDD2.n102 VSUBS 0.027991f
C135 VDD2.n103 VSUBS 0.012539f
C136 VDD2.n104 VSUBS 0.011843f
C137 VDD2.n105 VSUBS 0.022038f
C138 VDD2.n106 VSUBS 0.022038f
C139 VDD2.n107 VSUBS 0.011843f
C140 VDD2.n108 VSUBS 0.012539f
C141 VDD2.n109 VSUBS 0.027991f
C142 VDD2.n110 VSUBS 0.027991f
C143 VDD2.n111 VSUBS 0.027991f
C144 VDD2.n112 VSUBS 0.012191f
C145 VDD2.n113 VSUBS 0.011843f
C146 VDD2.n114 VSUBS 0.022038f
C147 VDD2.n115 VSUBS 0.022038f
C148 VDD2.n116 VSUBS 0.011843f
C149 VDD2.n117 VSUBS 0.012539f
C150 VDD2.n118 VSUBS 0.027991f
C151 VDD2.n119 VSUBS 0.027991f
C152 VDD2.n120 VSUBS 0.012539f
C153 VDD2.n121 VSUBS 0.011843f
C154 VDD2.n122 VSUBS 0.022038f
C155 VDD2.n123 VSUBS 0.022038f
C156 VDD2.n124 VSUBS 0.011843f
C157 VDD2.n125 VSUBS 0.012539f
C158 VDD2.n126 VSUBS 0.027991f
C159 VDD2.n127 VSUBS 0.064586f
C160 VDD2.n128 VSUBS 0.012539f
C161 VDD2.n129 VSUBS 0.011843f
C162 VDD2.n130 VSUBS 0.048231f
C163 VDD2.n131 VSUBS 0.047493f
C164 VDD2.n132 VSUBS 1.92216f
C165 VDD2.t3 VSUBS 0.209507f
C166 VDD2.t5 VSUBS 0.209507f
C167 VDD2.n133 VSUBS 1.6315f
C168 VN.n0 VSUBS 0.045069f
C169 VN.t1 VSUBS 1.7728f
C170 VN.n1 VSUBS 0.069453f
C171 VN.t5 VSUBS 1.86207f
C172 VN.t4 VSUBS 1.7728f
C173 VN.n2 VSUBS 0.716389f
C174 VN.n3 VSUBS 0.74891f
C175 VN.n4 VSUBS 0.235436f
C176 VN.n5 VSUBS 0.045069f
C177 VN.n6 VSUBS 0.036566f
C178 VN.n7 VSUBS 0.070589f
C179 VN.n8 VSUBS 0.72643f
C180 VN.n9 VSUBS 0.040078f
C181 VN.n10 VSUBS 0.045069f
C182 VN.t3 VSUBS 1.7728f
C183 VN.n11 VSUBS 0.069453f
C184 VN.t0 VSUBS 1.86207f
C185 VN.t2 VSUBS 1.7728f
C186 VN.n12 VSUBS 0.716389f
C187 VN.n13 VSUBS 0.74891f
C188 VN.n14 VSUBS 0.235436f
C189 VN.n15 VSUBS 0.045069f
C190 VN.n16 VSUBS 0.036566f
C191 VN.n17 VSUBS 0.070589f
C192 VN.n18 VSUBS 0.72643f
C193 VN.n19 VSUBS 1.9775f
C194 B.n0 VSUBS 0.004384f
C195 B.n1 VSUBS 0.004384f
C196 B.n2 VSUBS 0.006933f
C197 B.n3 VSUBS 0.006933f
C198 B.n4 VSUBS 0.006933f
C199 B.n5 VSUBS 0.006933f
C200 B.n6 VSUBS 0.006933f
C201 B.n7 VSUBS 0.006933f
C202 B.n8 VSUBS 0.006933f
C203 B.n9 VSUBS 0.006933f
C204 B.n10 VSUBS 0.006933f
C205 B.n11 VSUBS 0.006933f
C206 B.n12 VSUBS 0.006933f
C207 B.n13 VSUBS 0.006933f
C208 B.n14 VSUBS 0.006933f
C209 B.n15 VSUBS 0.016975f
C210 B.n16 VSUBS 0.006933f
C211 B.n17 VSUBS 0.006933f
C212 B.n18 VSUBS 0.006933f
C213 B.n19 VSUBS 0.006933f
C214 B.n20 VSUBS 0.006933f
C215 B.n21 VSUBS 0.006933f
C216 B.n22 VSUBS 0.006933f
C217 B.n23 VSUBS 0.006933f
C218 B.n24 VSUBS 0.006933f
C219 B.n25 VSUBS 0.006933f
C220 B.n26 VSUBS 0.006933f
C221 B.n27 VSUBS 0.006933f
C222 B.n28 VSUBS 0.006933f
C223 B.n29 VSUBS 0.006933f
C224 B.n30 VSUBS 0.006933f
C225 B.n31 VSUBS 0.006933f
C226 B.n32 VSUBS 0.006933f
C227 B.n33 VSUBS 0.006933f
C228 B.n34 VSUBS 0.006933f
C229 B.n35 VSUBS 0.006933f
C230 B.t2 VSUBS 0.209608f
C231 B.t1 VSUBS 0.22674f
C232 B.t0 VSUBS 0.614378f
C233 B.n36 VSUBS 0.338767f
C234 B.n37 VSUBS 0.24418f
C235 B.n38 VSUBS 0.016064f
C236 B.n39 VSUBS 0.006933f
C237 B.n40 VSUBS 0.006933f
C238 B.n41 VSUBS 0.006933f
C239 B.n42 VSUBS 0.006933f
C240 B.n43 VSUBS 0.006933f
C241 B.t5 VSUBS 0.209611f
C242 B.t4 VSUBS 0.226743f
C243 B.t3 VSUBS 0.614378f
C244 B.n44 VSUBS 0.338765f
C245 B.n45 VSUBS 0.244177f
C246 B.n46 VSUBS 0.006933f
C247 B.n47 VSUBS 0.006933f
C248 B.n48 VSUBS 0.006933f
C249 B.n49 VSUBS 0.006933f
C250 B.n50 VSUBS 0.006933f
C251 B.n51 VSUBS 0.006933f
C252 B.n52 VSUBS 0.006933f
C253 B.n53 VSUBS 0.006933f
C254 B.n54 VSUBS 0.006933f
C255 B.n55 VSUBS 0.006933f
C256 B.n56 VSUBS 0.006933f
C257 B.n57 VSUBS 0.006933f
C258 B.n58 VSUBS 0.006933f
C259 B.n59 VSUBS 0.006933f
C260 B.n60 VSUBS 0.006933f
C261 B.n61 VSUBS 0.006933f
C262 B.n62 VSUBS 0.006933f
C263 B.n63 VSUBS 0.006933f
C264 B.n64 VSUBS 0.006933f
C265 B.n65 VSUBS 0.006933f
C266 B.n66 VSUBS 0.016858f
C267 B.n67 VSUBS 0.006933f
C268 B.n68 VSUBS 0.006933f
C269 B.n69 VSUBS 0.006933f
C270 B.n70 VSUBS 0.006933f
C271 B.n71 VSUBS 0.006933f
C272 B.n72 VSUBS 0.006933f
C273 B.n73 VSUBS 0.006933f
C274 B.n74 VSUBS 0.006933f
C275 B.n75 VSUBS 0.006933f
C276 B.n76 VSUBS 0.006933f
C277 B.n77 VSUBS 0.006933f
C278 B.n78 VSUBS 0.006933f
C279 B.n79 VSUBS 0.006933f
C280 B.n80 VSUBS 0.006933f
C281 B.n81 VSUBS 0.006933f
C282 B.n82 VSUBS 0.006933f
C283 B.n83 VSUBS 0.006933f
C284 B.n84 VSUBS 0.006933f
C285 B.n85 VSUBS 0.006933f
C286 B.n86 VSUBS 0.006933f
C287 B.n87 VSUBS 0.006933f
C288 B.n88 VSUBS 0.006933f
C289 B.n89 VSUBS 0.006933f
C290 B.n90 VSUBS 0.006933f
C291 B.n91 VSUBS 0.006933f
C292 B.n92 VSUBS 0.016061f
C293 B.n93 VSUBS 0.006933f
C294 B.n94 VSUBS 0.006933f
C295 B.n95 VSUBS 0.006933f
C296 B.n96 VSUBS 0.006933f
C297 B.n97 VSUBS 0.006933f
C298 B.n98 VSUBS 0.006933f
C299 B.n99 VSUBS 0.006933f
C300 B.n100 VSUBS 0.006933f
C301 B.n101 VSUBS 0.006933f
C302 B.n102 VSUBS 0.006933f
C303 B.n103 VSUBS 0.006933f
C304 B.n104 VSUBS 0.006933f
C305 B.n105 VSUBS 0.006933f
C306 B.n106 VSUBS 0.006933f
C307 B.n107 VSUBS 0.006933f
C308 B.n108 VSUBS 0.006933f
C309 B.n109 VSUBS 0.006933f
C310 B.n110 VSUBS 0.006933f
C311 B.n111 VSUBS 0.006933f
C312 B.n112 VSUBS 0.006933f
C313 B.n113 VSUBS 0.006933f
C314 B.t10 VSUBS 0.209611f
C315 B.t11 VSUBS 0.226743f
C316 B.t9 VSUBS 0.614378f
C317 B.n114 VSUBS 0.338765f
C318 B.n115 VSUBS 0.244177f
C319 B.n116 VSUBS 0.006933f
C320 B.n117 VSUBS 0.006933f
C321 B.n118 VSUBS 0.006933f
C322 B.n119 VSUBS 0.006933f
C323 B.t7 VSUBS 0.209608f
C324 B.t8 VSUBS 0.22674f
C325 B.t6 VSUBS 0.614378f
C326 B.n120 VSUBS 0.338767f
C327 B.n121 VSUBS 0.24418f
C328 B.n122 VSUBS 0.016064f
C329 B.n123 VSUBS 0.006933f
C330 B.n124 VSUBS 0.006933f
C331 B.n125 VSUBS 0.006933f
C332 B.n126 VSUBS 0.006933f
C333 B.n127 VSUBS 0.006933f
C334 B.n128 VSUBS 0.006933f
C335 B.n129 VSUBS 0.006933f
C336 B.n130 VSUBS 0.006933f
C337 B.n131 VSUBS 0.006933f
C338 B.n132 VSUBS 0.006933f
C339 B.n133 VSUBS 0.006933f
C340 B.n134 VSUBS 0.006933f
C341 B.n135 VSUBS 0.006933f
C342 B.n136 VSUBS 0.006933f
C343 B.n137 VSUBS 0.006933f
C344 B.n138 VSUBS 0.006933f
C345 B.n139 VSUBS 0.006933f
C346 B.n140 VSUBS 0.006933f
C347 B.n141 VSUBS 0.006933f
C348 B.n142 VSUBS 0.006933f
C349 B.n143 VSUBS 0.016975f
C350 B.n144 VSUBS 0.006933f
C351 B.n145 VSUBS 0.006933f
C352 B.n146 VSUBS 0.006933f
C353 B.n147 VSUBS 0.006933f
C354 B.n148 VSUBS 0.006933f
C355 B.n149 VSUBS 0.006933f
C356 B.n150 VSUBS 0.006933f
C357 B.n151 VSUBS 0.006933f
C358 B.n152 VSUBS 0.006933f
C359 B.n153 VSUBS 0.006933f
C360 B.n154 VSUBS 0.006933f
C361 B.n155 VSUBS 0.006933f
C362 B.n156 VSUBS 0.006933f
C363 B.n157 VSUBS 0.006933f
C364 B.n158 VSUBS 0.006933f
C365 B.n159 VSUBS 0.006933f
C366 B.n160 VSUBS 0.006933f
C367 B.n161 VSUBS 0.006933f
C368 B.n162 VSUBS 0.006933f
C369 B.n163 VSUBS 0.006933f
C370 B.n164 VSUBS 0.006933f
C371 B.n165 VSUBS 0.006933f
C372 B.n166 VSUBS 0.006933f
C373 B.n167 VSUBS 0.006933f
C374 B.n168 VSUBS 0.006933f
C375 B.n169 VSUBS 0.006933f
C376 B.n170 VSUBS 0.006933f
C377 B.n171 VSUBS 0.006933f
C378 B.n172 VSUBS 0.006933f
C379 B.n173 VSUBS 0.006933f
C380 B.n174 VSUBS 0.006933f
C381 B.n175 VSUBS 0.006933f
C382 B.n176 VSUBS 0.006933f
C383 B.n177 VSUBS 0.006933f
C384 B.n178 VSUBS 0.006933f
C385 B.n179 VSUBS 0.006933f
C386 B.n180 VSUBS 0.006933f
C387 B.n181 VSUBS 0.006933f
C388 B.n182 VSUBS 0.006933f
C389 B.n183 VSUBS 0.006933f
C390 B.n184 VSUBS 0.006933f
C391 B.n185 VSUBS 0.006933f
C392 B.n186 VSUBS 0.006933f
C393 B.n187 VSUBS 0.006933f
C394 B.n188 VSUBS 0.006933f
C395 B.n189 VSUBS 0.006933f
C396 B.n190 VSUBS 0.006933f
C397 B.n191 VSUBS 0.006933f
C398 B.n192 VSUBS 0.016061f
C399 B.n193 VSUBS 0.016061f
C400 B.n194 VSUBS 0.016975f
C401 B.n195 VSUBS 0.006933f
C402 B.n196 VSUBS 0.006933f
C403 B.n197 VSUBS 0.006933f
C404 B.n198 VSUBS 0.006933f
C405 B.n199 VSUBS 0.006933f
C406 B.n200 VSUBS 0.006933f
C407 B.n201 VSUBS 0.006933f
C408 B.n202 VSUBS 0.006933f
C409 B.n203 VSUBS 0.006933f
C410 B.n204 VSUBS 0.006933f
C411 B.n205 VSUBS 0.006933f
C412 B.n206 VSUBS 0.006933f
C413 B.n207 VSUBS 0.006933f
C414 B.n208 VSUBS 0.006933f
C415 B.n209 VSUBS 0.006933f
C416 B.n210 VSUBS 0.006933f
C417 B.n211 VSUBS 0.006933f
C418 B.n212 VSUBS 0.006933f
C419 B.n213 VSUBS 0.006933f
C420 B.n214 VSUBS 0.006933f
C421 B.n215 VSUBS 0.006933f
C422 B.n216 VSUBS 0.006933f
C423 B.n217 VSUBS 0.006933f
C424 B.n218 VSUBS 0.006933f
C425 B.n219 VSUBS 0.006933f
C426 B.n220 VSUBS 0.006933f
C427 B.n221 VSUBS 0.006933f
C428 B.n222 VSUBS 0.006933f
C429 B.n223 VSUBS 0.006933f
C430 B.n224 VSUBS 0.006933f
C431 B.n225 VSUBS 0.006933f
C432 B.n226 VSUBS 0.006933f
C433 B.n227 VSUBS 0.006933f
C434 B.n228 VSUBS 0.006933f
C435 B.n229 VSUBS 0.006933f
C436 B.n230 VSUBS 0.006933f
C437 B.n231 VSUBS 0.006933f
C438 B.n232 VSUBS 0.006933f
C439 B.n233 VSUBS 0.006933f
C440 B.n234 VSUBS 0.006933f
C441 B.n235 VSUBS 0.006933f
C442 B.n236 VSUBS 0.006933f
C443 B.n237 VSUBS 0.006933f
C444 B.n238 VSUBS 0.006933f
C445 B.n239 VSUBS 0.006933f
C446 B.n240 VSUBS 0.006933f
C447 B.n241 VSUBS 0.006933f
C448 B.n242 VSUBS 0.006933f
C449 B.n243 VSUBS 0.006933f
C450 B.n244 VSUBS 0.006933f
C451 B.n245 VSUBS 0.006933f
C452 B.n246 VSUBS 0.006933f
C453 B.n247 VSUBS 0.006933f
C454 B.n248 VSUBS 0.006933f
C455 B.n249 VSUBS 0.006933f
C456 B.n250 VSUBS 0.006933f
C457 B.n251 VSUBS 0.006933f
C458 B.n252 VSUBS 0.006933f
C459 B.n253 VSUBS 0.006933f
C460 B.n254 VSUBS 0.006933f
C461 B.n255 VSUBS 0.004792f
C462 B.n256 VSUBS 0.006933f
C463 B.n257 VSUBS 0.006933f
C464 B.n258 VSUBS 0.005608f
C465 B.n259 VSUBS 0.006933f
C466 B.n260 VSUBS 0.006933f
C467 B.n261 VSUBS 0.006933f
C468 B.n262 VSUBS 0.006933f
C469 B.n263 VSUBS 0.006933f
C470 B.n264 VSUBS 0.006933f
C471 B.n265 VSUBS 0.006933f
C472 B.n266 VSUBS 0.006933f
C473 B.n267 VSUBS 0.006933f
C474 B.n268 VSUBS 0.006933f
C475 B.n269 VSUBS 0.006933f
C476 B.n270 VSUBS 0.005608f
C477 B.n271 VSUBS 0.016064f
C478 B.n272 VSUBS 0.004792f
C479 B.n273 VSUBS 0.006933f
C480 B.n274 VSUBS 0.006933f
C481 B.n275 VSUBS 0.006933f
C482 B.n276 VSUBS 0.006933f
C483 B.n277 VSUBS 0.006933f
C484 B.n278 VSUBS 0.006933f
C485 B.n279 VSUBS 0.006933f
C486 B.n280 VSUBS 0.006933f
C487 B.n281 VSUBS 0.006933f
C488 B.n282 VSUBS 0.006933f
C489 B.n283 VSUBS 0.006933f
C490 B.n284 VSUBS 0.006933f
C491 B.n285 VSUBS 0.006933f
C492 B.n286 VSUBS 0.006933f
C493 B.n287 VSUBS 0.006933f
C494 B.n288 VSUBS 0.006933f
C495 B.n289 VSUBS 0.006933f
C496 B.n290 VSUBS 0.006933f
C497 B.n291 VSUBS 0.006933f
C498 B.n292 VSUBS 0.006933f
C499 B.n293 VSUBS 0.006933f
C500 B.n294 VSUBS 0.006933f
C501 B.n295 VSUBS 0.006933f
C502 B.n296 VSUBS 0.006933f
C503 B.n297 VSUBS 0.006933f
C504 B.n298 VSUBS 0.006933f
C505 B.n299 VSUBS 0.006933f
C506 B.n300 VSUBS 0.006933f
C507 B.n301 VSUBS 0.006933f
C508 B.n302 VSUBS 0.006933f
C509 B.n303 VSUBS 0.006933f
C510 B.n304 VSUBS 0.006933f
C511 B.n305 VSUBS 0.006933f
C512 B.n306 VSUBS 0.006933f
C513 B.n307 VSUBS 0.006933f
C514 B.n308 VSUBS 0.006933f
C515 B.n309 VSUBS 0.006933f
C516 B.n310 VSUBS 0.006933f
C517 B.n311 VSUBS 0.006933f
C518 B.n312 VSUBS 0.006933f
C519 B.n313 VSUBS 0.006933f
C520 B.n314 VSUBS 0.006933f
C521 B.n315 VSUBS 0.006933f
C522 B.n316 VSUBS 0.006933f
C523 B.n317 VSUBS 0.006933f
C524 B.n318 VSUBS 0.006933f
C525 B.n319 VSUBS 0.006933f
C526 B.n320 VSUBS 0.006933f
C527 B.n321 VSUBS 0.006933f
C528 B.n322 VSUBS 0.006933f
C529 B.n323 VSUBS 0.006933f
C530 B.n324 VSUBS 0.006933f
C531 B.n325 VSUBS 0.006933f
C532 B.n326 VSUBS 0.006933f
C533 B.n327 VSUBS 0.006933f
C534 B.n328 VSUBS 0.006933f
C535 B.n329 VSUBS 0.006933f
C536 B.n330 VSUBS 0.006933f
C537 B.n331 VSUBS 0.006933f
C538 B.n332 VSUBS 0.006933f
C539 B.n333 VSUBS 0.016975f
C540 B.n334 VSUBS 0.016975f
C541 B.n335 VSUBS 0.016061f
C542 B.n336 VSUBS 0.006933f
C543 B.n337 VSUBS 0.006933f
C544 B.n338 VSUBS 0.006933f
C545 B.n339 VSUBS 0.006933f
C546 B.n340 VSUBS 0.006933f
C547 B.n341 VSUBS 0.006933f
C548 B.n342 VSUBS 0.006933f
C549 B.n343 VSUBS 0.006933f
C550 B.n344 VSUBS 0.006933f
C551 B.n345 VSUBS 0.006933f
C552 B.n346 VSUBS 0.006933f
C553 B.n347 VSUBS 0.006933f
C554 B.n348 VSUBS 0.006933f
C555 B.n349 VSUBS 0.006933f
C556 B.n350 VSUBS 0.006933f
C557 B.n351 VSUBS 0.006933f
C558 B.n352 VSUBS 0.006933f
C559 B.n353 VSUBS 0.006933f
C560 B.n354 VSUBS 0.006933f
C561 B.n355 VSUBS 0.006933f
C562 B.n356 VSUBS 0.006933f
C563 B.n357 VSUBS 0.006933f
C564 B.n358 VSUBS 0.006933f
C565 B.n359 VSUBS 0.006933f
C566 B.n360 VSUBS 0.006933f
C567 B.n361 VSUBS 0.006933f
C568 B.n362 VSUBS 0.006933f
C569 B.n363 VSUBS 0.006933f
C570 B.n364 VSUBS 0.006933f
C571 B.n365 VSUBS 0.006933f
C572 B.n366 VSUBS 0.006933f
C573 B.n367 VSUBS 0.006933f
C574 B.n368 VSUBS 0.006933f
C575 B.n369 VSUBS 0.006933f
C576 B.n370 VSUBS 0.006933f
C577 B.n371 VSUBS 0.006933f
C578 B.n372 VSUBS 0.006933f
C579 B.n373 VSUBS 0.006933f
C580 B.n374 VSUBS 0.006933f
C581 B.n375 VSUBS 0.006933f
C582 B.n376 VSUBS 0.006933f
C583 B.n377 VSUBS 0.006933f
C584 B.n378 VSUBS 0.006933f
C585 B.n379 VSUBS 0.006933f
C586 B.n380 VSUBS 0.006933f
C587 B.n381 VSUBS 0.006933f
C588 B.n382 VSUBS 0.006933f
C589 B.n383 VSUBS 0.006933f
C590 B.n384 VSUBS 0.006933f
C591 B.n385 VSUBS 0.006933f
C592 B.n386 VSUBS 0.006933f
C593 B.n387 VSUBS 0.006933f
C594 B.n388 VSUBS 0.006933f
C595 B.n389 VSUBS 0.006933f
C596 B.n390 VSUBS 0.006933f
C597 B.n391 VSUBS 0.006933f
C598 B.n392 VSUBS 0.006933f
C599 B.n393 VSUBS 0.006933f
C600 B.n394 VSUBS 0.006933f
C601 B.n395 VSUBS 0.006933f
C602 B.n396 VSUBS 0.006933f
C603 B.n397 VSUBS 0.006933f
C604 B.n398 VSUBS 0.006933f
C605 B.n399 VSUBS 0.006933f
C606 B.n400 VSUBS 0.006933f
C607 B.n401 VSUBS 0.006933f
C608 B.n402 VSUBS 0.006933f
C609 B.n403 VSUBS 0.006933f
C610 B.n404 VSUBS 0.006933f
C611 B.n405 VSUBS 0.006933f
C612 B.n406 VSUBS 0.006933f
C613 B.n407 VSUBS 0.006933f
C614 B.n408 VSUBS 0.006933f
C615 B.n409 VSUBS 0.006933f
C616 B.n410 VSUBS 0.006933f
C617 B.n411 VSUBS 0.006933f
C618 B.n412 VSUBS 0.006933f
C619 B.n413 VSUBS 0.016061f
C620 B.n414 VSUBS 0.016975f
C621 B.n415 VSUBS 0.016178f
C622 B.n416 VSUBS 0.006933f
C623 B.n417 VSUBS 0.006933f
C624 B.n418 VSUBS 0.006933f
C625 B.n419 VSUBS 0.006933f
C626 B.n420 VSUBS 0.006933f
C627 B.n421 VSUBS 0.006933f
C628 B.n422 VSUBS 0.006933f
C629 B.n423 VSUBS 0.006933f
C630 B.n424 VSUBS 0.006933f
C631 B.n425 VSUBS 0.006933f
C632 B.n426 VSUBS 0.006933f
C633 B.n427 VSUBS 0.006933f
C634 B.n428 VSUBS 0.006933f
C635 B.n429 VSUBS 0.006933f
C636 B.n430 VSUBS 0.006933f
C637 B.n431 VSUBS 0.006933f
C638 B.n432 VSUBS 0.006933f
C639 B.n433 VSUBS 0.006933f
C640 B.n434 VSUBS 0.006933f
C641 B.n435 VSUBS 0.006933f
C642 B.n436 VSUBS 0.006933f
C643 B.n437 VSUBS 0.006933f
C644 B.n438 VSUBS 0.006933f
C645 B.n439 VSUBS 0.006933f
C646 B.n440 VSUBS 0.006933f
C647 B.n441 VSUBS 0.006933f
C648 B.n442 VSUBS 0.006933f
C649 B.n443 VSUBS 0.006933f
C650 B.n444 VSUBS 0.006933f
C651 B.n445 VSUBS 0.006933f
C652 B.n446 VSUBS 0.006933f
C653 B.n447 VSUBS 0.006933f
C654 B.n448 VSUBS 0.006933f
C655 B.n449 VSUBS 0.006933f
C656 B.n450 VSUBS 0.006933f
C657 B.n451 VSUBS 0.006933f
C658 B.n452 VSUBS 0.006933f
C659 B.n453 VSUBS 0.006933f
C660 B.n454 VSUBS 0.006933f
C661 B.n455 VSUBS 0.006933f
C662 B.n456 VSUBS 0.006933f
C663 B.n457 VSUBS 0.006933f
C664 B.n458 VSUBS 0.006933f
C665 B.n459 VSUBS 0.006933f
C666 B.n460 VSUBS 0.006933f
C667 B.n461 VSUBS 0.006933f
C668 B.n462 VSUBS 0.006933f
C669 B.n463 VSUBS 0.006933f
C670 B.n464 VSUBS 0.006933f
C671 B.n465 VSUBS 0.006933f
C672 B.n466 VSUBS 0.006933f
C673 B.n467 VSUBS 0.006933f
C674 B.n468 VSUBS 0.006933f
C675 B.n469 VSUBS 0.006933f
C676 B.n470 VSUBS 0.006933f
C677 B.n471 VSUBS 0.006933f
C678 B.n472 VSUBS 0.006933f
C679 B.n473 VSUBS 0.006933f
C680 B.n474 VSUBS 0.006933f
C681 B.n475 VSUBS 0.006933f
C682 B.n476 VSUBS 0.004792f
C683 B.n477 VSUBS 0.016064f
C684 B.n478 VSUBS 0.005608f
C685 B.n479 VSUBS 0.006933f
C686 B.n480 VSUBS 0.006933f
C687 B.n481 VSUBS 0.006933f
C688 B.n482 VSUBS 0.006933f
C689 B.n483 VSUBS 0.006933f
C690 B.n484 VSUBS 0.006933f
C691 B.n485 VSUBS 0.006933f
C692 B.n486 VSUBS 0.006933f
C693 B.n487 VSUBS 0.006933f
C694 B.n488 VSUBS 0.006933f
C695 B.n489 VSUBS 0.006933f
C696 B.n490 VSUBS 0.005608f
C697 B.n491 VSUBS 0.006933f
C698 B.n492 VSUBS 0.006933f
C699 B.n493 VSUBS 0.004792f
C700 B.n494 VSUBS 0.006933f
C701 B.n495 VSUBS 0.006933f
C702 B.n496 VSUBS 0.006933f
C703 B.n497 VSUBS 0.006933f
C704 B.n498 VSUBS 0.006933f
C705 B.n499 VSUBS 0.006933f
C706 B.n500 VSUBS 0.006933f
C707 B.n501 VSUBS 0.006933f
C708 B.n502 VSUBS 0.006933f
C709 B.n503 VSUBS 0.006933f
C710 B.n504 VSUBS 0.006933f
C711 B.n505 VSUBS 0.006933f
C712 B.n506 VSUBS 0.006933f
C713 B.n507 VSUBS 0.006933f
C714 B.n508 VSUBS 0.006933f
C715 B.n509 VSUBS 0.006933f
C716 B.n510 VSUBS 0.006933f
C717 B.n511 VSUBS 0.006933f
C718 B.n512 VSUBS 0.006933f
C719 B.n513 VSUBS 0.006933f
C720 B.n514 VSUBS 0.006933f
C721 B.n515 VSUBS 0.006933f
C722 B.n516 VSUBS 0.006933f
C723 B.n517 VSUBS 0.006933f
C724 B.n518 VSUBS 0.006933f
C725 B.n519 VSUBS 0.006933f
C726 B.n520 VSUBS 0.006933f
C727 B.n521 VSUBS 0.006933f
C728 B.n522 VSUBS 0.006933f
C729 B.n523 VSUBS 0.006933f
C730 B.n524 VSUBS 0.006933f
C731 B.n525 VSUBS 0.006933f
C732 B.n526 VSUBS 0.006933f
C733 B.n527 VSUBS 0.006933f
C734 B.n528 VSUBS 0.006933f
C735 B.n529 VSUBS 0.006933f
C736 B.n530 VSUBS 0.006933f
C737 B.n531 VSUBS 0.006933f
C738 B.n532 VSUBS 0.006933f
C739 B.n533 VSUBS 0.006933f
C740 B.n534 VSUBS 0.006933f
C741 B.n535 VSUBS 0.006933f
C742 B.n536 VSUBS 0.006933f
C743 B.n537 VSUBS 0.006933f
C744 B.n538 VSUBS 0.006933f
C745 B.n539 VSUBS 0.006933f
C746 B.n540 VSUBS 0.006933f
C747 B.n541 VSUBS 0.006933f
C748 B.n542 VSUBS 0.006933f
C749 B.n543 VSUBS 0.006933f
C750 B.n544 VSUBS 0.006933f
C751 B.n545 VSUBS 0.006933f
C752 B.n546 VSUBS 0.006933f
C753 B.n547 VSUBS 0.006933f
C754 B.n548 VSUBS 0.006933f
C755 B.n549 VSUBS 0.006933f
C756 B.n550 VSUBS 0.006933f
C757 B.n551 VSUBS 0.006933f
C758 B.n552 VSUBS 0.006933f
C759 B.n553 VSUBS 0.006933f
C760 B.n554 VSUBS 0.016975f
C761 B.n555 VSUBS 0.016061f
C762 B.n556 VSUBS 0.016061f
C763 B.n557 VSUBS 0.006933f
C764 B.n558 VSUBS 0.006933f
C765 B.n559 VSUBS 0.006933f
C766 B.n560 VSUBS 0.006933f
C767 B.n561 VSUBS 0.006933f
C768 B.n562 VSUBS 0.006933f
C769 B.n563 VSUBS 0.006933f
C770 B.n564 VSUBS 0.006933f
C771 B.n565 VSUBS 0.006933f
C772 B.n566 VSUBS 0.006933f
C773 B.n567 VSUBS 0.006933f
C774 B.n568 VSUBS 0.006933f
C775 B.n569 VSUBS 0.006933f
C776 B.n570 VSUBS 0.006933f
C777 B.n571 VSUBS 0.006933f
C778 B.n572 VSUBS 0.006933f
C779 B.n573 VSUBS 0.006933f
C780 B.n574 VSUBS 0.006933f
C781 B.n575 VSUBS 0.006933f
C782 B.n576 VSUBS 0.006933f
C783 B.n577 VSUBS 0.006933f
C784 B.n578 VSUBS 0.006933f
C785 B.n579 VSUBS 0.006933f
C786 B.n580 VSUBS 0.006933f
C787 B.n581 VSUBS 0.006933f
C788 B.n582 VSUBS 0.006933f
C789 B.n583 VSUBS 0.006933f
C790 B.n584 VSUBS 0.006933f
C791 B.n585 VSUBS 0.006933f
C792 B.n586 VSUBS 0.006933f
C793 B.n587 VSUBS 0.006933f
C794 B.n588 VSUBS 0.006933f
C795 B.n589 VSUBS 0.006933f
C796 B.n590 VSUBS 0.006933f
C797 B.n591 VSUBS 0.006933f
C798 B.n592 VSUBS 0.006933f
C799 B.n593 VSUBS 0.006933f
C800 B.n594 VSUBS 0.006933f
C801 B.n595 VSUBS 0.0157f
C802 VDD1.n0 VSUBS 0.02348f
C803 VDD1.n1 VSUBS 0.022225f
C804 VDD1.n2 VSUBS 0.011943f
C805 VDD1.n3 VSUBS 0.028229f
C806 VDD1.n4 VSUBS 0.012646f
C807 VDD1.n5 VSUBS 0.022225f
C808 VDD1.n6 VSUBS 0.011943f
C809 VDD1.n7 VSUBS 0.028229f
C810 VDD1.n8 VSUBS 0.012646f
C811 VDD1.n9 VSUBS 0.022225f
C812 VDD1.n10 VSUBS 0.012294f
C813 VDD1.n11 VSUBS 0.028229f
C814 VDD1.n12 VSUBS 0.011943f
C815 VDD1.n13 VSUBS 0.012646f
C816 VDD1.n14 VSUBS 0.022225f
C817 VDD1.n15 VSUBS 0.011943f
C818 VDD1.n16 VSUBS 0.028229f
C819 VDD1.n17 VSUBS 0.012646f
C820 VDD1.n18 VSUBS 0.022225f
C821 VDD1.n19 VSUBS 0.011943f
C822 VDD1.n20 VSUBS 0.021172f
C823 VDD1.n21 VSUBS 0.021235f
C824 VDD1.t3 VSUBS 0.060831f
C825 VDD1.n22 VSUBS 0.175338f
C826 VDD1.n23 VSUBS 1.09492f
C827 VDD1.n24 VSUBS 0.011943f
C828 VDD1.n25 VSUBS 0.012646f
C829 VDD1.n26 VSUBS 0.028229f
C830 VDD1.n27 VSUBS 0.028229f
C831 VDD1.n28 VSUBS 0.012646f
C832 VDD1.n29 VSUBS 0.011943f
C833 VDD1.n30 VSUBS 0.022225f
C834 VDD1.n31 VSUBS 0.022225f
C835 VDD1.n32 VSUBS 0.011943f
C836 VDD1.n33 VSUBS 0.012646f
C837 VDD1.n34 VSUBS 0.028229f
C838 VDD1.n35 VSUBS 0.028229f
C839 VDD1.n36 VSUBS 0.012646f
C840 VDD1.n37 VSUBS 0.011943f
C841 VDD1.n38 VSUBS 0.022225f
C842 VDD1.n39 VSUBS 0.022225f
C843 VDD1.n40 VSUBS 0.011943f
C844 VDD1.n41 VSUBS 0.012646f
C845 VDD1.n42 VSUBS 0.028229f
C846 VDD1.n43 VSUBS 0.028229f
C847 VDD1.n44 VSUBS 0.028229f
C848 VDD1.n45 VSUBS 0.012294f
C849 VDD1.n46 VSUBS 0.011943f
C850 VDD1.n47 VSUBS 0.022225f
C851 VDD1.n48 VSUBS 0.022225f
C852 VDD1.n49 VSUBS 0.011943f
C853 VDD1.n50 VSUBS 0.012646f
C854 VDD1.n51 VSUBS 0.028229f
C855 VDD1.n52 VSUBS 0.028229f
C856 VDD1.n53 VSUBS 0.012646f
C857 VDD1.n54 VSUBS 0.011943f
C858 VDD1.n55 VSUBS 0.022225f
C859 VDD1.n56 VSUBS 0.022225f
C860 VDD1.n57 VSUBS 0.011943f
C861 VDD1.n58 VSUBS 0.012646f
C862 VDD1.n59 VSUBS 0.028229f
C863 VDD1.n60 VSUBS 0.065134f
C864 VDD1.n61 VSUBS 0.012646f
C865 VDD1.n62 VSUBS 0.011943f
C866 VDD1.n63 VSUBS 0.04864f
C867 VDD1.n64 VSUBS 0.050424f
C868 VDD1.n65 VSUBS 0.02348f
C869 VDD1.n66 VSUBS 0.022225f
C870 VDD1.n67 VSUBS 0.011943f
C871 VDD1.n68 VSUBS 0.028229f
C872 VDD1.n69 VSUBS 0.012646f
C873 VDD1.n70 VSUBS 0.022225f
C874 VDD1.n71 VSUBS 0.011943f
C875 VDD1.n72 VSUBS 0.028229f
C876 VDD1.n73 VSUBS 0.012646f
C877 VDD1.n74 VSUBS 0.022225f
C878 VDD1.n75 VSUBS 0.012294f
C879 VDD1.n76 VSUBS 0.028229f
C880 VDD1.n77 VSUBS 0.012646f
C881 VDD1.n78 VSUBS 0.022225f
C882 VDD1.n79 VSUBS 0.011943f
C883 VDD1.n80 VSUBS 0.028229f
C884 VDD1.n81 VSUBS 0.012646f
C885 VDD1.n82 VSUBS 0.022225f
C886 VDD1.n83 VSUBS 0.011943f
C887 VDD1.n84 VSUBS 0.021172f
C888 VDD1.n85 VSUBS 0.021235f
C889 VDD1.t4 VSUBS 0.060831f
C890 VDD1.n86 VSUBS 0.175339f
C891 VDD1.n87 VSUBS 1.09493f
C892 VDD1.n88 VSUBS 0.011943f
C893 VDD1.n89 VSUBS 0.012646f
C894 VDD1.n90 VSUBS 0.028229f
C895 VDD1.n91 VSUBS 0.028229f
C896 VDD1.n92 VSUBS 0.012646f
C897 VDD1.n93 VSUBS 0.011943f
C898 VDD1.n94 VSUBS 0.022225f
C899 VDD1.n95 VSUBS 0.022225f
C900 VDD1.n96 VSUBS 0.011943f
C901 VDD1.n97 VSUBS 0.012646f
C902 VDD1.n98 VSUBS 0.028229f
C903 VDD1.n99 VSUBS 0.028229f
C904 VDD1.n100 VSUBS 0.012646f
C905 VDD1.n101 VSUBS 0.011943f
C906 VDD1.n102 VSUBS 0.022225f
C907 VDD1.n103 VSUBS 0.022225f
C908 VDD1.n104 VSUBS 0.011943f
C909 VDD1.n105 VSUBS 0.011943f
C910 VDD1.n106 VSUBS 0.012646f
C911 VDD1.n107 VSUBS 0.028229f
C912 VDD1.n108 VSUBS 0.028229f
C913 VDD1.n109 VSUBS 0.028229f
C914 VDD1.n110 VSUBS 0.012294f
C915 VDD1.n111 VSUBS 0.011943f
C916 VDD1.n112 VSUBS 0.022225f
C917 VDD1.n113 VSUBS 0.022225f
C918 VDD1.n114 VSUBS 0.011943f
C919 VDD1.n115 VSUBS 0.012646f
C920 VDD1.n116 VSUBS 0.028229f
C921 VDD1.n117 VSUBS 0.028229f
C922 VDD1.n118 VSUBS 0.012646f
C923 VDD1.n119 VSUBS 0.011943f
C924 VDD1.n120 VSUBS 0.022225f
C925 VDD1.n121 VSUBS 0.022225f
C926 VDD1.n122 VSUBS 0.011943f
C927 VDD1.n123 VSUBS 0.012646f
C928 VDD1.n124 VSUBS 0.028229f
C929 VDD1.n125 VSUBS 0.065134f
C930 VDD1.n126 VSUBS 0.012646f
C931 VDD1.n127 VSUBS 0.011943f
C932 VDD1.n128 VSUBS 0.04864f
C933 VDD1.n129 VSUBS 0.050008f
C934 VDD1.t2 VSUBS 0.211285f
C935 VDD1.t1 VSUBS 0.211285f
C936 VDD1.n130 VSUBS 1.64537f
C937 VDD1.n131 VSUBS 2.15983f
C938 VDD1.t0 VSUBS 0.211285f
C939 VDD1.t5 VSUBS 0.211285f
C940 VDD1.n132 VSUBS 1.64329f
C941 VDD1.n133 VSUBS 2.37175f
C942 VTAIL.t2 VSUBS 0.26943f
C943 VTAIL.t1 VSUBS 0.26943f
C944 VTAIL.n0 VSUBS 1.93454f
C945 VTAIL.n1 VSUBS 0.801289f
C946 VTAIL.n2 VSUBS 0.029942f
C947 VTAIL.n3 VSUBS 0.028342f
C948 VTAIL.n4 VSUBS 0.01523f
C949 VTAIL.n5 VSUBS 0.035997f
C950 VTAIL.n6 VSUBS 0.016125f
C951 VTAIL.n7 VSUBS 0.028342f
C952 VTAIL.n8 VSUBS 0.01523f
C953 VTAIL.n9 VSUBS 0.035997f
C954 VTAIL.n10 VSUBS 0.016125f
C955 VTAIL.n11 VSUBS 0.028342f
C956 VTAIL.n12 VSUBS 0.015678f
C957 VTAIL.n13 VSUBS 0.035997f
C958 VTAIL.n14 VSUBS 0.016125f
C959 VTAIL.n15 VSUBS 0.028342f
C960 VTAIL.n16 VSUBS 0.01523f
C961 VTAIL.n17 VSUBS 0.035997f
C962 VTAIL.n18 VSUBS 0.016125f
C963 VTAIL.n19 VSUBS 0.028342f
C964 VTAIL.n20 VSUBS 0.01523f
C965 VTAIL.n21 VSUBS 0.026998f
C966 VTAIL.n22 VSUBS 0.027079f
C967 VTAIL.t7 VSUBS 0.077572f
C968 VTAIL.n23 VSUBS 0.223592f
C969 VTAIL.n24 VSUBS 1.39625f
C970 VTAIL.n25 VSUBS 0.01523f
C971 VTAIL.n26 VSUBS 0.016125f
C972 VTAIL.n27 VSUBS 0.035997f
C973 VTAIL.n28 VSUBS 0.035997f
C974 VTAIL.n29 VSUBS 0.016125f
C975 VTAIL.n30 VSUBS 0.01523f
C976 VTAIL.n31 VSUBS 0.028342f
C977 VTAIL.n32 VSUBS 0.028342f
C978 VTAIL.n33 VSUBS 0.01523f
C979 VTAIL.n34 VSUBS 0.016125f
C980 VTAIL.n35 VSUBS 0.035997f
C981 VTAIL.n36 VSUBS 0.035997f
C982 VTAIL.n37 VSUBS 0.016125f
C983 VTAIL.n38 VSUBS 0.01523f
C984 VTAIL.n39 VSUBS 0.028342f
C985 VTAIL.n40 VSUBS 0.028342f
C986 VTAIL.n41 VSUBS 0.01523f
C987 VTAIL.n42 VSUBS 0.01523f
C988 VTAIL.n43 VSUBS 0.016125f
C989 VTAIL.n44 VSUBS 0.035997f
C990 VTAIL.n45 VSUBS 0.035997f
C991 VTAIL.n46 VSUBS 0.035997f
C992 VTAIL.n47 VSUBS 0.015678f
C993 VTAIL.n48 VSUBS 0.01523f
C994 VTAIL.n49 VSUBS 0.028342f
C995 VTAIL.n50 VSUBS 0.028342f
C996 VTAIL.n51 VSUBS 0.01523f
C997 VTAIL.n52 VSUBS 0.016125f
C998 VTAIL.n53 VSUBS 0.035997f
C999 VTAIL.n54 VSUBS 0.035997f
C1000 VTAIL.n55 VSUBS 0.016125f
C1001 VTAIL.n56 VSUBS 0.01523f
C1002 VTAIL.n57 VSUBS 0.028342f
C1003 VTAIL.n58 VSUBS 0.028342f
C1004 VTAIL.n59 VSUBS 0.01523f
C1005 VTAIL.n60 VSUBS 0.016125f
C1006 VTAIL.n61 VSUBS 0.035997f
C1007 VTAIL.n62 VSUBS 0.083059f
C1008 VTAIL.n63 VSUBS 0.016125f
C1009 VTAIL.n64 VSUBS 0.01523f
C1010 VTAIL.n65 VSUBS 0.062026f
C1011 VTAIL.n66 VSUBS 0.041478f
C1012 VTAIL.n67 VSUBS 0.245827f
C1013 VTAIL.t9 VSUBS 0.26943f
C1014 VTAIL.t10 VSUBS 0.26943f
C1015 VTAIL.n68 VSUBS 1.93454f
C1016 VTAIL.n69 VSUBS 2.35617f
C1017 VTAIL.t0 VSUBS 0.26943f
C1018 VTAIL.t11 VSUBS 0.26943f
C1019 VTAIL.n70 VSUBS 1.93455f
C1020 VTAIL.n71 VSUBS 2.35615f
C1021 VTAIL.n72 VSUBS 0.029942f
C1022 VTAIL.n73 VSUBS 0.028342f
C1023 VTAIL.n74 VSUBS 0.01523f
C1024 VTAIL.n75 VSUBS 0.035997f
C1025 VTAIL.n76 VSUBS 0.016125f
C1026 VTAIL.n77 VSUBS 0.028342f
C1027 VTAIL.n78 VSUBS 0.01523f
C1028 VTAIL.n79 VSUBS 0.035997f
C1029 VTAIL.n80 VSUBS 0.016125f
C1030 VTAIL.n81 VSUBS 0.028342f
C1031 VTAIL.n82 VSUBS 0.015678f
C1032 VTAIL.n83 VSUBS 0.035997f
C1033 VTAIL.n84 VSUBS 0.01523f
C1034 VTAIL.n85 VSUBS 0.016125f
C1035 VTAIL.n86 VSUBS 0.028342f
C1036 VTAIL.n87 VSUBS 0.01523f
C1037 VTAIL.n88 VSUBS 0.035997f
C1038 VTAIL.n89 VSUBS 0.016125f
C1039 VTAIL.n90 VSUBS 0.028342f
C1040 VTAIL.n91 VSUBS 0.01523f
C1041 VTAIL.n92 VSUBS 0.026998f
C1042 VTAIL.n93 VSUBS 0.027079f
C1043 VTAIL.t4 VSUBS 0.077572f
C1044 VTAIL.n94 VSUBS 0.223592f
C1045 VTAIL.n95 VSUBS 1.39625f
C1046 VTAIL.n96 VSUBS 0.01523f
C1047 VTAIL.n97 VSUBS 0.016125f
C1048 VTAIL.n98 VSUBS 0.035997f
C1049 VTAIL.n99 VSUBS 0.035997f
C1050 VTAIL.n100 VSUBS 0.016125f
C1051 VTAIL.n101 VSUBS 0.01523f
C1052 VTAIL.n102 VSUBS 0.028342f
C1053 VTAIL.n103 VSUBS 0.028342f
C1054 VTAIL.n104 VSUBS 0.01523f
C1055 VTAIL.n105 VSUBS 0.016125f
C1056 VTAIL.n106 VSUBS 0.035997f
C1057 VTAIL.n107 VSUBS 0.035997f
C1058 VTAIL.n108 VSUBS 0.016125f
C1059 VTAIL.n109 VSUBS 0.01523f
C1060 VTAIL.n110 VSUBS 0.028342f
C1061 VTAIL.n111 VSUBS 0.028342f
C1062 VTAIL.n112 VSUBS 0.01523f
C1063 VTAIL.n113 VSUBS 0.016125f
C1064 VTAIL.n114 VSUBS 0.035997f
C1065 VTAIL.n115 VSUBS 0.035997f
C1066 VTAIL.n116 VSUBS 0.035997f
C1067 VTAIL.n117 VSUBS 0.015678f
C1068 VTAIL.n118 VSUBS 0.01523f
C1069 VTAIL.n119 VSUBS 0.028342f
C1070 VTAIL.n120 VSUBS 0.028342f
C1071 VTAIL.n121 VSUBS 0.01523f
C1072 VTAIL.n122 VSUBS 0.016125f
C1073 VTAIL.n123 VSUBS 0.035997f
C1074 VTAIL.n124 VSUBS 0.035997f
C1075 VTAIL.n125 VSUBS 0.016125f
C1076 VTAIL.n126 VSUBS 0.01523f
C1077 VTAIL.n127 VSUBS 0.028342f
C1078 VTAIL.n128 VSUBS 0.028342f
C1079 VTAIL.n129 VSUBS 0.01523f
C1080 VTAIL.n130 VSUBS 0.016125f
C1081 VTAIL.n131 VSUBS 0.035997f
C1082 VTAIL.n132 VSUBS 0.083059f
C1083 VTAIL.n133 VSUBS 0.016125f
C1084 VTAIL.n134 VSUBS 0.01523f
C1085 VTAIL.n135 VSUBS 0.062026f
C1086 VTAIL.n136 VSUBS 0.041478f
C1087 VTAIL.n137 VSUBS 0.245827f
C1088 VTAIL.t6 VSUBS 0.26943f
C1089 VTAIL.t5 VSUBS 0.26943f
C1090 VTAIL.n138 VSUBS 1.93455f
C1091 VTAIL.n139 VSUBS 0.8863f
C1092 VTAIL.n140 VSUBS 0.029942f
C1093 VTAIL.n141 VSUBS 0.028342f
C1094 VTAIL.n142 VSUBS 0.01523f
C1095 VTAIL.n143 VSUBS 0.035997f
C1096 VTAIL.n144 VSUBS 0.016125f
C1097 VTAIL.n145 VSUBS 0.028342f
C1098 VTAIL.n146 VSUBS 0.01523f
C1099 VTAIL.n147 VSUBS 0.035997f
C1100 VTAIL.n148 VSUBS 0.016125f
C1101 VTAIL.n149 VSUBS 0.028342f
C1102 VTAIL.n150 VSUBS 0.015678f
C1103 VTAIL.n151 VSUBS 0.035997f
C1104 VTAIL.n152 VSUBS 0.01523f
C1105 VTAIL.n153 VSUBS 0.016125f
C1106 VTAIL.n154 VSUBS 0.028342f
C1107 VTAIL.n155 VSUBS 0.01523f
C1108 VTAIL.n156 VSUBS 0.035997f
C1109 VTAIL.n157 VSUBS 0.016125f
C1110 VTAIL.n158 VSUBS 0.028342f
C1111 VTAIL.n159 VSUBS 0.01523f
C1112 VTAIL.n160 VSUBS 0.026998f
C1113 VTAIL.n161 VSUBS 0.027079f
C1114 VTAIL.t8 VSUBS 0.077572f
C1115 VTAIL.n162 VSUBS 0.223592f
C1116 VTAIL.n163 VSUBS 1.39625f
C1117 VTAIL.n164 VSUBS 0.01523f
C1118 VTAIL.n165 VSUBS 0.016125f
C1119 VTAIL.n166 VSUBS 0.035997f
C1120 VTAIL.n167 VSUBS 0.035997f
C1121 VTAIL.n168 VSUBS 0.016125f
C1122 VTAIL.n169 VSUBS 0.01523f
C1123 VTAIL.n170 VSUBS 0.028342f
C1124 VTAIL.n171 VSUBS 0.028342f
C1125 VTAIL.n172 VSUBS 0.01523f
C1126 VTAIL.n173 VSUBS 0.016125f
C1127 VTAIL.n174 VSUBS 0.035997f
C1128 VTAIL.n175 VSUBS 0.035997f
C1129 VTAIL.n176 VSUBS 0.016125f
C1130 VTAIL.n177 VSUBS 0.01523f
C1131 VTAIL.n178 VSUBS 0.028342f
C1132 VTAIL.n179 VSUBS 0.028342f
C1133 VTAIL.n180 VSUBS 0.01523f
C1134 VTAIL.n181 VSUBS 0.016125f
C1135 VTAIL.n182 VSUBS 0.035997f
C1136 VTAIL.n183 VSUBS 0.035997f
C1137 VTAIL.n184 VSUBS 0.035997f
C1138 VTAIL.n185 VSUBS 0.015678f
C1139 VTAIL.n186 VSUBS 0.01523f
C1140 VTAIL.n187 VSUBS 0.028342f
C1141 VTAIL.n188 VSUBS 0.028342f
C1142 VTAIL.n189 VSUBS 0.01523f
C1143 VTAIL.n190 VSUBS 0.016125f
C1144 VTAIL.n191 VSUBS 0.035997f
C1145 VTAIL.n192 VSUBS 0.035997f
C1146 VTAIL.n193 VSUBS 0.016125f
C1147 VTAIL.n194 VSUBS 0.01523f
C1148 VTAIL.n195 VSUBS 0.028342f
C1149 VTAIL.n196 VSUBS 0.028342f
C1150 VTAIL.n197 VSUBS 0.01523f
C1151 VTAIL.n198 VSUBS 0.016125f
C1152 VTAIL.n199 VSUBS 0.035997f
C1153 VTAIL.n200 VSUBS 0.083059f
C1154 VTAIL.n201 VSUBS 0.016125f
C1155 VTAIL.n202 VSUBS 0.01523f
C1156 VTAIL.n203 VSUBS 0.062026f
C1157 VTAIL.n204 VSUBS 0.041478f
C1158 VTAIL.n205 VSUBS 1.59523f
C1159 VTAIL.n206 VSUBS 0.029942f
C1160 VTAIL.n207 VSUBS 0.028342f
C1161 VTAIL.n208 VSUBS 0.01523f
C1162 VTAIL.n209 VSUBS 0.035997f
C1163 VTAIL.n210 VSUBS 0.016125f
C1164 VTAIL.n211 VSUBS 0.028342f
C1165 VTAIL.n212 VSUBS 0.01523f
C1166 VTAIL.n213 VSUBS 0.035997f
C1167 VTAIL.n214 VSUBS 0.016125f
C1168 VTAIL.n215 VSUBS 0.028342f
C1169 VTAIL.n216 VSUBS 0.015678f
C1170 VTAIL.n217 VSUBS 0.035997f
C1171 VTAIL.n218 VSUBS 0.016125f
C1172 VTAIL.n219 VSUBS 0.028342f
C1173 VTAIL.n220 VSUBS 0.01523f
C1174 VTAIL.n221 VSUBS 0.035997f
C1175 VTAIL.n222 VSUBS 0.016125f
C1176 VTAIL.n223 VSUBS 0.028342f
C1177 VTAIL.n224 VSUBS 0.01523f
C1178 VTAIL.n225 VSUBS 0.026998f
C1179 VTAIL.n226 VSUBS 0.027079f
C1180 VTAIL.t3 VSUBS 0.077572f
C1181 VTAIL.n227 VSUBS 0.223592f
C1182 VTAIL.n228 VSUBS 1.39625f
C1183 VTAIL.n229 VSUBS 0.01523f
C1184 VTAIL.n230 VSUBS 0.016125f
C1185 VTAIL.n231 VSUBS 0.035997f
C1186 VTAIL.n232 VSUBS 0.035997f
C1187 VTAIL.n233 VSUBS 0.016125f
C1188 VTAIL.n234 VSUBS 0.01523f
C1189 VTAIL.n235 VSUBS 0.028342f
C1190 VTAIL.n236 VSUBS 0.028342f
C1191 VTAIL.n237 VSUBS 0.01523f
C1192 VTAIL.n238 VSUBS 0.016125f
C1193 VTAIL.n239 VSUBS 0.035997f
C1194 VTAIL.n240 VSUBS 0.035997f
C1195 VTAIL.n241 VSUBS 0.016125f
C1196 VTAIL.n242 VSUBS 0.01523f
C1197 VTAIL.n243 VSUBS 0.028342f
C1198 VTAIL.n244 VSUBS 0.028342f
C1199 VTAIL.n245 VSUBS 0.01523f
C1200 VTAIL.n246 VSUBS 0.01523f
C1201 VTAIL.n247 VSUBS 0.016125f
C1202 VTAIL.n248 VSUBS 0.035997f
C1203 VTAIL.n249 VSUBS 0.035997f
C1204 VTAIL.n250 VSUBS 0.035997f
C1205 VTAIL.n251 VSUBS 0.015678f
C1206 VTAIL.n252 VSUBS 0.01523f
C1207 VTAIL.n253 VSUBS 0.028342f
C1208 VTAIL.n254 VSUBS 0.028342f
C1209 VTAIL.n255 VSUBS 0.01523f
C1210 VTAIL.n256 VSUBS 0.016125f
C1211 VTAIL.n257 VSUBS 0.035997f
C1212 VTAIL.n258 VSUBS 0.035997f
C1213 VTAIL.n259 VSUBS 0.016125f
C1214 VTAIL.n260 VSUBS 0.01523f
C1215 VTAIL.n261 VSUBS 0.028342f
C1216 VTAIL.n262 VSUBS 0.028342f
C1217 VTAIL.n263 VSUBS 0.01523f
C1218 VTAIL.n264 VSUBS 0.016125f
C1219 VTAIL.n265 VSUBS 0.035997f
C1220 VTAIL.n266 VSUBS 0.083059f
C1221 VTAIL.n267 VSUBS 0.016125f
C1222 VTAIL.n268 VSUBS 0.01523f
C1223 VTAIL.n269 VSUBS 0.062026f
C1224 VTAIL.n270 VSUBS 0.041478f
C1225 VTAIL.n271 VSUBS 1.5598f
C1226 VP.n0 VSUBS 0.04633f
C1227 VP.t4 VSUBS 1.8224f
C1228 VP.n1 VSUBS 0.071396f
C1229 VP.n2 VSUBS 0.04633f
C1230 VP.t1 VSUBS 1.8224f
C1231 VP.n3 VSUBS 0.746753f
C1232 VP.n4 VSUBS 0.04633f
C1233 VP.t0 VSUBS 1.8224f
C1234 VP.n5 VSUBS 0.071396f
C1235 VP.t2 VSUBS 1.91416f
C1236 VP.t5 VSUBS 1.8224f
C1237 VP.n6 VSUBS 0.736432f
C1238 VP.n7 VSUBS 0.769862f
C1239 VP.n8 VSUBS 0.242023f
C1240 VP.n9 VSUBS 0.04633f
C1241 VP.n10 VSUBS 0.037589f
C1242 VP.n11 VSUBS 0.072564f
C1243 VP.n12 VSUBS 0.746753f
C1244 VP.n13 VSUBS 2.00246f
C1245 VP.n14 VSUBS 2.04108f
C1246 VP.n15 VSUBS 0.04633f
C1247 VP.n16 VSUBS 0.072564f
C1248 VP.n17 VSUBS 0.037589f
C1249 VP.t3 VSUBS 1.8224f
C1250 VP.n18 VSUBS 0.667407f
C1251 VP.n19 VSUBS 0.071396f
C1252 VP.n20 VSUBS 0.04633f
C1253 VP.n21 VSUBS 0.04633f
C1254 VP.n22 VSUBS 0.04633f
C1255 VP.n23 VSUBS 0.037589f
C1256 VP.n24 VSUBS 0.072564f
C1257 VP.n25 VSUBS 0.746753f
C1258 VP.n26 VSUBS 0.041199f
.ends

