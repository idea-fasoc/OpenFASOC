* NGSPICE file created from diff_pair_sample_0150.ext - technology: sky130A

.subckt diff_pair_sample_0150 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t9 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X1 VDD2.t9 VN.t0 VTAIL.t5 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=4.1106 ps=21.86 w=10.54 l=3.57
X2 VTAIL.t18 VP.t1 VDD1.t8 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X3 VTAIL.t17 VP.t2 VDD1.t2 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X4 VDD2.t8 VN.t1 VTAIL.t9 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=1.7391 ps=10.87 w=10.54 l=3.57
X5 B.t11 B.t9 B.t10 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=0 ps=0 w=10.54 l=3.57
X6 VTAIL.t2 VN.t2 VDD2.t7 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X7 VDD1.t1 VP.t3 VTAIL.t16 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=4.1106 ps=21.86 w=10.54 l=3.57
X8 VTAIL.t0 VN.t3 VDD2.t6 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X9 VTAIL.t8 VN.t4 VDD2.t5 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X10 VDD1.t0 VP.t4 VTAIL.t15 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=4.1106 ps=21.86 w=10.54 l=3.57
X11 VDD2.t4 VN.t5 VTAIL.t3 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=4.1106 ps=21.86 w=10.54 l=3.57
X12 VTAIL.t4 VN.t6 VDD2.t3 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X13 VDD2.t2 VN.t7 VTAIL.t1 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=1.7391 ps=10.87 w=10.54 l=3.57
X14 VDD1.t7 VP.t5 VTAIL.t14 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X15 B.t8 B.t6 B.t7 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=0 ps=0 w=10.54 l=3.57
X16 B.t5 B.t3 B.t4 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=0 ps=0 w=10.54 l=3.57
X17 VDD1.t6 VP.t6 VTAIL.t13 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=1.7391 ps=10.87 w=10.54 l=3.57
X18 VDD1.t5 VP.t7 VTAIL.t12 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=1.7391 ps=10.87 w=10.54 l=3.57
X19 VDD1.t3 VP.t8 VTAIL.t11 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X20 B.t2 B.t0 B.t1 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=4.1106 pd=21.86 as=0 ps=0 w=10.54 l=3.57
X21 VTAIL.t10 VP.t9 VDD1.t4 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X22 VDD2.t1 VN.t8 VTAIL.t6 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
X23 VDD2.t0 VN.t9 VTAIL.t7 w_n5650_n3076# sky130_fd_pr__pfet_01v8 ad=1.7391 pd=10.87 as=1.7391 ps=10.87 w=10.54 l=3.57
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n31 VP.t7 103.013
R57 VP.n72 VP.n71 87.7864
R58 VP.n124 VP.n0 87.7864
R59 VP.n70 VP.n17 87.7864
R60 VP.n71 VP.t6 71.1529
R61 VP.n83 VP.t0 71.1529
R62 VP.n96 VP.t8 71.1529
R63 VP.n109 VP.t1 71.1529
R64 VP.n0 VP.t4 71.1529
R65 VP.n17 VP.t3 71.1529
R66 VP.n55 VP.t2 71.1529
R67 VP.n42 VP.t5 71.1529
R68 VP.n30 VP.t9 71.1529
R69 VP.n31 VP.n30 67.5381
R70 VP.n72 VP.n70 57.2723
R71 VP.n90 VP.n10 56.5617
R72 VP.n103 VP.n6 56.5617
R73 VP.n49 VP.n23 56.5617
R74 VP.n36 VP.n27 56.5617
R75 VP.n77 VP.n14 50.2647
R76 VP.n116 VP.n2 50.2647
R77 VP.n62 VP.n19 50.2647
R78 VP.n81 VP.n14 30.8893
R79 VP.n116 VP.n115 30.8893
R80 VP.n62 VP.n61 30.8893
R81 VP.n75 VP.n16 24.5923
R82 VP.n76 VP.n75 24.5923
R83 VP.n77 VP.n76 24.5923
R84 VP.n82 VP.n81 24.5923
R85 VP.n84 VP.n82 24.5923
R86 VP.n88 VP.n12 24.5923
R87 VP.n89 VP.n88 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n94 VP.n10 24.5923
R90 VP.n95 VP.n94 24.5923
R91 VP.n97 VP.n95 24.5923
R92 VP.n101 VP.n8 24.5923
R93 VP.n102 VP.n101 24.5923
R94 VP.n103 VP.n102 24.5923
R95 VP.n107 VP.n6 24.5923
R96 VP.n108 VP.n107 24.5923
R97 VP.n110 VP.n108 24.5923
R98 VP.n114 VP.n4 24.5923
R99 VP.n115 VP.n114 24.5923
R100 VP.n120 VP.n2 24.5923
R101 VP.n121 VP.n120 24.5923
R102 VP.n122 VP.n121 24.5923
R103 VP.n66 VP.n19 24.5923
R104 VP.n67 VP.n66 24.5923
R105 VP.n68 VP.n67 24.5923
R106 VP.n53 VP.n23 24.5923
R107 VP.n54 VP.n53 24.5923
R108 VP.n56 VP.n54 24.5923
R109 VP.n60 VP.n21 24.5923
R110 VP.n61 VP.n60 24.5923
R111 VP.n40 VP.n27 24.5923
R112 VP.n41 VP.n40 24.5923
R113 VP.n43 VP.n41 24.5923
R114 VP.n47 VP.n25 24.5923
R115 VP.n48 VP.n47 24.5923
R116 VP.n49 VP.n48 24.5923
R117 VP.n34 VP.n29 24.5923
R118 VP.n35 VP.n34 24.5923
R119 VP.n36 VP.n35 24.5923
R120 VP.n84 VP.n83 17.2148
R121 VP.n109 VP.n4 17.2148
R122 VP.n55 VP.n21 17.2148
R123 VP.n97 VP.n96 12.2964
R124 VP.n96 VP.n8 12.2964
R125 VP.n43 VP.n42 12.2964
R126 VP.n42 VP.n25 12.2964
R127 VP.n83 VP.n12 7.37805
R128 VP.n110 VP.n109 7.37805
R129 VP.n56 VP.n55 7.37805
R130 VP.n30 VP.n29 7.37805
R131 VP.n32 VP.n31 3.3822
R132 VP.n71 VP.n16 2.45968
R133 VP.n122 VP.n0 2.45968
R134 VP.n68 VP.n17 2.45968
R135 VP.n70 VP.n69 0.354861
R136 VP.n73 VP.n72 0.354861
R137 VP.n124 VP.n123 0.354861
R138 VP VP.n124 0.267071
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VDD1.n1 VDD1.t5 87.1814
R194 VDD1.n3 VDD1.t6 87.1811
R195 VDD1.n5 VDD1.n4 83.2013
R196 VDD1.n1 VDD1.n0 80.7354
R197 VDD1.n7 VDD1.n6 80.7352
R198 VDD1.n3 VDD1.n2 80.7351
R199 VDD1.n7 VDD1.n5 51.0354
R200 VDD1.n6 VDD1.t2 3.08447
R201 VDD1.n6 VDD1.t1 3.08447
R202 VDD1.n0 VDD1.t4 3.08447
R203 VDD1.n0 VDD1.t7 3.08447
R204 VDD1.n4 VDD1.t8 3.08447
R205 VDD1.n4 VDD1.t0 3.08447
R206 VDD1.n2 VDD1.t9 3.08447
R207 VDD1.n2 VDD1.t3 3.08447
R208 VDD1 VDD1.n7 2.46386
R209 VDD1 VDD1.n1 0.899207
R210 VDD1.n5 VDD1.n3 0.785671
R211 VTAIL.n11 VTAIL.t3 67.1405
R212 VTAIL.n16 VTAIL.t16 67.1403
R213 VTAIL.n17 VTAIL.t5 67.1403
R214 VTAIL.n2 VTAIL.t15 67.1403
R215 VTAIL.n15 VTAIL.n14 64.0566
R216 VTAIL.n13 VTAIL.n12 64.0566
R217 VTAIL.n10 VTAIL.n9 64.0566
R218 VTAIL.n8 VTAIL.n7 64.0566
R219 VTAIL.n19 VTAIL.n18 64.0563
R220 VTAIL.n1 VTAIL.n0 64.0563
R221 VTAIL.n4 VTAIL.n3 64.0563
R222 VTAIL.n6 VTAIL.n5 64.0563
R223 VTAIL.n8 VTAIL.n6 28.1772
R224 VTAIL.n17 VTAIL.n16 24.8152
R225 VTAIL.n10 VTAIL.n8 3.36257
R226 VTAIL.n11 VTAIL.n10 3.36257
R227 VTAIL.n15 VTAIL.n13 3.36257
R228 VTAIL.n16 VTAIL.n15 3.36257
R229 VTAIL.n6 VTAIL.n4 3.36257
R230 VTAIL.n4 VTAIL.n2 3.36257
R231 VTAIL.n19 VTAIL.n17 3.36257
R232 VTAIL.n18 VTAIL.t7 3.08447
R233 VTAIL.n18 VTAIL.t2 3.08447
R234 VTAIL.n0 VTAIL.t1 3.08447
R235 VTAIL.n0 VTAIL.t0 3.08447
R236 VTAIL.n3 VTAIL.t11 3.08447
R237 VTAIL.n3 VTAIL.t18 3.08447
R238 VTAIL.n5 VTAIL.t13 3.08447
R239 VTAIL.n5 VTAIL.t19 3.08447
R240 VTAIL.n14 VTAIL.t14 3.08447
R241 VTAIL.n14 VTAIL.t17 3.08447
R242 VTAIL.n12 VTAIL.t12 3.08447
R243 VTAIL.n12 VTAIL.t10 3.08447
R244 VTAIL.n9 VTAIL.t6 3.08447
R245 VTAIL.n9 VTAIL.t4 3.08447
R246 VTAIL.n7 VTAIL.t9 3.08447
R247 VTAIL.n7 VTAIL.t8 3.08447
R248 VTAIL VTAIL.n1 2.58024
R249 VTAIL.n13 VTAIL.n11 2.15136
R250 VTAIL.n2 VTAIL.n1 2.15136
R251 VTAIL VTAIL.n19 0.782828
R252 VN.n106 VN.n105 161.3
R253 VN.n104 VN.n55 161.3
R254 VN.n103 VN.n102 161.3
R255 VN.n101 VN.n56 161.3
R256 VN.n100 VN.n99 161.3
R257 VN.n98 VN.n57 161.3
R258 VN.n97 VN.n96 161.3
R259 VN.n95 VN.n58 161.3
R260 VN.n94 VN.n93 161.3
R261 VN.n92 VN.n59 161.3
R262 VN.n91 VN.n90 161.3
R263 VN.n89 VN.n61 161.3
R264 VN.n88 VN.n87 161.3
R265 VN.n86 VN.n62 161.3
R266 VN.n85 VN.n84 161.3
R267 VN.n83 VN.n63 161.3
R268 VN.n82 VN.n81 161.3
R269 VN.n80 VN.n64 161.3
R270 VN.n79 VN.n78 161.3
R271 VN.n77 VN.n66 161.3
R272 VN.n76 VN.n75 161.3
R273 VN.n74 VN.n67 161.3
R274 VN.n73 VN.n72 161.3
R275 VN.n71 VN.n68 161.3
R276 VN.n52 VN.n51 161.3
R277 VN.n50 VN.n1 161.3
R278 VN.n49 VN.n48 161.3
R279 VN.n47 VN.n2 161.3
R280 VN.n46 VN.n45 161.3
R281 VN.n44 VN.n3 161.3
R282 VN.n43 VN.n42 161.3
R283 VN.n41 VN.n4 161.3
R284 VN.n40 VN.n39 161.3
R285 VN.n37 VN.n5 161.3
R286 VN.n36 VN.n35 161.3
R287 VN.n34 VN.n6 161.3
R288 VN.n33 VN.n32 161.3
R289 VN.n31 VN.n7 161.3
R290 VN.n30 VN.n29 161.3
R291 VN.n28 VN.n8 161.3
R292 VN.n27 VN.n26 161.3
R293 VN.n24 VN.n9 161.3
R294 VN.n23 VN.n22 161.3
R295 VN.n21 VN.n10 161.3
R296 VN.n20 VN.n19 161.3
R297 VN.n18 VN.n11 161.3
R298 VN.n17 VN.n16 161.3
R299 VN.n15 VN.n12 161.3
R300 VN.n70 VN.t5 103.013
R301 VN.n14 VN.t7 103.013
R302 VN.n53 VN.n0 87.7864
R303 VN.n107 VN.n54 87.7864
R304 VN.n13 VN.t3 71.1529
R305 VN.n25 VN.t9 71.1529
R306 VN.n38 VN.t2 71.1529
R307 VN.n0 VN.t0 71.1529
R308 VN.n69 VN.t6 71.1529
R309 VN.n65 VN.t8 71.1529
R310 VN.n60 VN.t4 71.1529
R311 VN.n54 VN.t1 71.1529
R312 VN.n14 VN.n13 67.5381
R313 VN.n70 VN.n69 67.5381
R314 VN VN.n107 57.4375
R315 VN.n19 VN.n10 56.5617
R316 VN.n32 VN.n6 56.5617
R317 VN.n75 VN.n66 56.5617
R318 VN.n87 VN.n61 56.5617
R319 VN.n45 VN.n2 50.2647
R320 VN.n99 VN.n56 50.2647
R321 VN.n45 VN.n44 30.8893
R322 VN.n99 VN.n98 30.8893
R323 VN.n17 VN.n12 24.5923
R324 VN.n18 VN.n17 24.5923
R325 VN.n19 VN.n18 24.5923
R326 VN.n23 VN.n10 24.5923
R327 VN.n24 VN.n23 24.5923
R328 VN.n26 VN.n24 24.5923
R329 VN.n30 VN.n8 24.5923
R330 VN.n31 VN.n30 24.5923
R331 VN.n32 VN.n31 24.5923
R332 VN.n36 VN.n6 24.5923
R333 VN.n37 VN.n36 24.5923
R334 VN.n39 VN.n37 24.5923
R335 VN.n43 VN.n4 24.5923
R336 VN.n44 VN.n43 24.5923
R337 VN.n49 VN.n2 24.5923
R338 VN.n50 VN.n49 24.5923
R339 VN.n51 VN.n50 24.5923
R340 VN.n75 VN.n74 24.5923
R341 VN.n74 VN.n73 24.5923
R342 VN.n73 VN.n68 24.5923
R343 VN.n87 VN.n86 24.5923
R344 VN.n86 VN.n85 24.5923
R345 VN.n85 VN.n63 24.5923
R346 VN.n81 VN.n80 24.5923
R347 VN.n80 VN.n79 24.5923
R348 VN.n79 VN.n66 24.5923
R349 VN.n98 VN.n97 24.5923
R350 VN.n97 VN.n58 24.5923
R351 VN.n93 VN.n92 24.5923
R352 VN.n92 VN.n91 24.5923
R353 VN.n91 VN.n61 24.5923
R354 VN.n105 VN.n104 24.5923
R355 VN.n104 VN.n103 24.5923
R356 VN.n103 VN.n56 24.5923
R357 VN.n38 VN.n4 17.2148
R358 VN.n60 VN.n58 17.2148
R359 VN.n26 VN.n25 12.2964
R360 VN.n25 VN.n8 12.2964
R361 VN.n65 VN.n63 12.2964
R362 VN.n81 VN.n65 12.2964
R363 VN.n13 VN.n12 7.37805
R364 VN.n39 VN.n38 7.37805
R365 VN.n69 VN.n68 7.37805
R366 VN.n93 VN.n60 7.37805
R367 VN.n71 VN.n70 3.38222
R368 VN.n15 VN.n14 3.38222
R369 VN.n51 VN.n0 2.45968
R370 VN.n105 VN.n54 2.45968
R371 VN.n107 VN.n106 0.354861
R372 VN.n53 VN.n52 0.354861
R373 VN VN.n53 0.267071
R374 VN.n106 VN.n55 0.189894
R375 VN.n102 VN.n55 0.189894
R376 VN.n102 VN.n101 0.189894
R377 VN.n101 VN.n100 0.189894
R378 VN.n100 VN.n57 0.189894
R379 VN.n96 VN.n57 0.189894
R380 VN.n96 VN.n95 0.189894
R381 VN.n95 VN.n94 0.189894
R382 VN.n94 VN.n59 0.189894
R383 VN.n90 VN.n59 0.189894
R384 VN.n90 VN.n89 0.189894
R385 VN.n89 VN.n88 0.189894
R386 VN.n88 VN.n62 0.189894
R387 VN.n84 VN.n62 0.189894
R388 VN.n84 VN.n83 0.189894
R389 VN.n83 VN.n82 0.189894
R390 VN.n82 VN.n64 0.189894
R391 VN.n78 VN.n64 0.189894
R392 VN.n78 VN.n77 0.189894
R393 VN.n77 VN.n76 0.189894
R394 VN.n76 VN.n67 0.189894
R395 VN.n72 VN.n67 0.189894
R396 VN.n72 VN.n71 0.189894
R397 VN.n16 VN.n15 0.189894
R398 VN.n16 VN.n11 0.189894
R399 VN.n20 VN.n11 0.189894
R400 VN.n21 VN.n20 0.189894
R401 VN.n22 VN.n21 0.189894
R402 VN.n22 VN.n9 0.189894
R403 VN.n27 VN.n9 0.189894
R404 VN.n28 VN.n27 0.189894
R405 VN.n29 VN.n28 0.189894
R406 VN.n29 VN.n7 0.189894
R407 VN.n33 VN.n7 0.189894
R408 VN.n34 VN.n33 0.189894
R409 VN.n35 VN.n34 0.189894
R410 VN.n35 VN.n5 0.189894
R411 VN.n40 VN.n5 0.189894
R412 VN.n41 VN.n40 0.189894
R413 VN.n42 VN.n41 0.189894
R414 VN.n42 VN.n3 0.189894
R415 VN.n46 VN.n3 0.189894
R416 VN.n47 VN.n46 0.189894
R417 VN.n48 VN.n47 0.189894
R418 VN.n48 VN.n1 0.189894
R419 VN.n52 VN.n1 0.189894
R420 VDD2.n1 VDD2.t2 87.1811
R421 VDD2.n4 VDD2.t8 83.8193
R422 VDD2.n3 VDD2.n2 83.2013
R423 VDD2 VDD2.n7 83.1985
R424 VDD2.n6 VDD2.n5 80.7354
R425 VDD2.n1 VDD2.n0 80.7351
R426 VDD2.n4 VDD2.n3 48.7713
R427 VDD2.n6 VDD2.n4 3.36257
R428 VDD2.n7 VDD2.t3 3.08447
R429 VDD2.n7 VDD2.t4 3.08447
R430 VDD2.n5 VDD2.t5 3.08447
R431 VDD2.n5 VDD2.t1 3.08447
R432 VDD2.n2 VDD2.t7 3.08447
R433 VDD2.n2 VDD2.t9 3.08447
R434 VDD2.n0 VDD2.t6 3.08447
R435 VDD2.n0 VDD2.t0 3.08447
R436 VDD2 VDD2.n6 0.899207
R437 VDD2.n3 VDD2.n1 0.785671
R438 B.n724 B.n723 585
R439 B.n725 B.n86 585
R440 B.n727 B.n726 585
R441 B.n728 B.n85 585
R442 B.n730 B.n729 585
R443 B.n731 B.n84 585
R444 B.n733 B.n732 585
R445 B.n734 B.n83 585
R446 B.n736 B.n735 585
R447 B.n737 B.n82 585
R448 B.n739 B.n738 585
R449 B.n740 B.n81 585
R450 B.n742 B.n741 585
R451 B.n743 B.n80 585
R452 B.n745 B.n744 585
R453 B.n746 B.n79 585
R454 B.n748 B.n747 585
R455 B.n749 B.n78 585
R456 B.n751 B.n750 585
R457 B.n752 B.n77 585
R458 B.n754 B.n753 585
R459 B.n755 B.n76 585
R460 B.n757 B.n756 585
R461 B.n758 B.n75 585
R462 B.n760 B.n759 585
R463 B.n761 B.n74 585
R464 B.n763 B.n762 585
R465 B.n764 B.n73 585
R466 B.n766 B.n765 585
R467 B.n767 B.n72 585
R468 B.n769 B.n768 585
R469 B.n770 B.n71 585
R470 B.n772 B.n771 585
R471 B.n773 B.n70 585
R472 B.n775 B.n774 585
R473 B.n776 B.n69 585
R474 B.n778 B.n777 585
R475 B.n780 B.n779 585
R476 B.n781 B.n65 585
R477 B.n783 B.n782 585
R478 B.n784 B.n64 585
R479 B.n786 B.n785 585
R480 B.n787 B.n63 585
R481 B.n789 B.n788 585
R482 B.n790 B.n62 585
R483 B.n792 B.n791 585
R484 B.n793 B.n59 585
R485 B.n796 B.n795 585
R486 B.n797 B.n58 585
R487 B.n799 B.n798 585
R488 B.n800 B.n57 585
R489 B.n802 B.n801 585
R490 B.n803 B.n56 585
R491 B.n805 B.n804 585
R492 B.n806 B.n55 585
R493 B.n808 B.n807 585
R494 B.n809 B.n54 585
R495 B.n811 B.n810 585
R496 B.n812 B.n53 585
R497 B.n814 B.n813 585
R498 B.n815 B.n52 585
R499 B.n817 B.n816 585
R500 B.n818 B.n51 585
R501 B.n820 B.n819 585
R502 B.n821 B.n50 585
R503 B.n823 B.n822 585
R504 B.n824 B.n49 585
R505 B.n826 B.n825 585
R506 B.n827 B.n48 585
R507 B.n829 B.n828 585
R508 B.n830 B.n47 585
R509 B.n832 B.n831 585
R510 B.n833 B.n46 585
R511 B.n835 B.n834 585
R512 B.n836 B.n45 585
R513 B.n838 B.n837 585
R514 B.n839 B.n44 585
R515 B.n841 B.n840 585
R516 B.n842 B.n43 585
R517 B.n844 B.n843 585
R518 B.n845 B.n42 585
R519 B.n847 B.n846 585
R520 B.n848 B.n41 585
R521 B.n850 B.n849 585
R522 B.n722 B.n87 585
R523 B.n721 B.n720 585
R524 B.n719 B.n88 585
R525 B.n718 B.n717 585
R526 B.n716 B.n89 585
R527 B.n715 B.n714 585
R528 B.n713 B.n90 585
R529 B.n712 B.n711 585
R530 B.n710 B.n91 585
R531 B.n709 B.n708 585
R532 B.n707 B.n92 585
R533 B.n706 B.n705 585
R534 B.n704 B.n93 585
R535 B.n703 B.n702 585
R536 B.n701 B.n94 585
R537 B.n700 B.n699 585
R538 B.n698 B.n95 585
R539 B.n697 B.n696 585
R540 B.n695 B.n96 585
R541 B.n694 B.n693 585
R542 B.n692 B.n97 585
R543 B.n691 B.n690 585
R544 B.n689 B.n98 585
R545 B.n688 B.n687 585
R546 B.n686 B.n99 585
R547 B.n685 B.n684 585
R548 B.n683 B.n100 585
R549 B.n682 B.n681 585
R550 B.n680 B.n101 585
R551 B.n679 B.n678 585
R552 B.n677 B.n102 585
R553 B.n676 B.n675 585
R554 B.n674 B.n103 585
R555 B.n673 B.n672 585
R556 B.n671 B.n104 585
R557 B.n670 B.n669 585
R558 B.n668 B.n105 585
R559 B.n667 B.n666 585
R560 B.n665 B.n106 585
R561 B.n664 B.n663 585
R562 B.n662 B.n107 585
R563 B.n661 B.n660 585
R564 B.n659 B.n108 585
R565 B.n658 B.n657 585
R566 B.n656 B.n109 585
R567 B.n655 B.n654 585
R568 B.n653 B.n110 585
R569 B.n652 B.n651 585
R570 B.n650 B.n111 585
R571 B.n649 B.n648 585
R572 B.n647 B.n112 585
R573 B.n646 B.n645 585
R574 B.n644 B.n113 585
R575 B.n643 B.n642 585
R576 B.n641 B.n114 585
R577 B.n640 B.n639 585
R578 B.n638 B.n115 585
R579 B.n637 B.n636 585
R580 B.n635 B.n116 585
R581 B.n634 B.n633 585
R582 B.n632 B.n117 585
R583 B.n631 B.n630 585
R584 B.n629 B.n118 585
R585 B.n628 B.n627 585
R586 B.n626 B.n119 585
R587 B.n625 B.n624 585
R588 B.n623 B.n120 585
R589 B.n622 B.n621 585
R590 B.n620 B.n121 585
R591 B.n619 B.n618 585
R592 B.n617 B.n122 585
R593 B.n616 B.n615 585
R594 B.n614 B.n123 585
R595 B.n613 B.n612 585
R596 B.n611 B.n124 585
R597 B.n610 B.n609 585
R598 B.n608 B.n125 585
R599 B.n607 B.n606 585
R600 B.n605 B.n126 585
R601 B.n604 B.n603 585
R602 B.n602 B.n127 585
R603 B.n601 B.n600 585
R604 B.n599 B.n128 585
R605 B.n598 B.n597 585
R606 B.n596 B.n129 585
R607 B.n595 B.n594 585
R608 B.n593 B.n130 585
R609 B.n592 B.n591 585
R610 B.n590 B.n131 585
R611 B.n589 B.n588 585
R612 B.n587 B.n132 585
R613 B.n586 B.n585 585
R614 B.n584 B.n133 585
R615 B.n583 B.n582 585
R616 B.n581 B.n134 585
R617 B.n580 B.n579 585
R618 B.n578 B.n135 585
R619 B.n577 B.n576 585
R620 B.n575 B.n136 585
R621 B.n574 B.n573 585
R622 B.n572 B.n137 585
R623 B.n571 B.n570 585
R624 B.n569 B.n138 585
R625 B.n568 B.n567 585
R626 B.n566 B.n139 585
R627 B.n565 B.n564 585
R628 B.n563 B.n140 585
R629 B.n562 B.n561 585
R630 B.n560 B.n141 585
R631 B.n559 B.n558 585
R632 B.n557 B.n142 585
R633 B.n556 B.n555 585
R634 B.n554 B.n143 585
R635 B.n553 B.n552 585
R636 B.n551 B.n144 585
R637 B.n550 B.n549 585
R638 B.n548 B.n145 585
R639 B.n547 B.n546 585
R640 B.n545 B.n146 585
R641 B.n544 B.n543 585
R642 B.n542 B.n147 585
R643 B.n541 B.n540 585
R644 B.n539 B.n148 585
R645 B.n538 B.n537 585
R646 B.n536 B.n149 585
R647 B.n535 B.n534 585
R648 B.n533 B.n150 585
R649 B.n532 B.n531 585
R650 B.n530 B.n151 585
R651 B.n529 B.n528 585
R652 B.n527 B.n152 585
R653 B.n526 B.n525 585
R654 B.n524 B.n153 585
R655 B.n523 B.n522 585
R656 B.n521 B.n154 585
R657 B.n520 B.n519 585
R658 B.n518 B.n155 585
R659 B.n517 B.n516 585
R660 B.n515 B.n156 585
R661 B.n514 B.n513 585
R662 B.n512 B.n157 585
R663 B.n511 B.n510 585
R664 B.n509 B.n158 585
R665 B.n508 B.n507 585
R666 B.n506 B.n159 585
R667 B.n505 B.n504 585
R668 B.n503 B.n160 585
R669 B.n502 B.n501 585
R670 B.n500 B.n161 585
R671 B.n499 B.n498 585
R672 B.n497 B.n162 585
R673 B.n496 B.n495 585
R674 B.n494 B.n163 585
R675 B.n493 B.n492 585
R676 B.n491 B.n164 585
R677 B.n364 B.n363 585
R678 B.n365 B.n210 585
R679 B.n367 B.n366 585
R680 B.n368 B.n209 585
R681 B.n370 B.n369 585
R682 B.n371 B.n208 585
R683 B.n373 B.n372 585
R684 B.n374 B.n207 585
R685 B.n376 B.n375 585
R686 B.n377 B.n206 585
R687 B.n379 B.n378 585
R688 B.n380 B.n205 585
R689 B.n382 B.n381 585
R690 B.n383 B.n204 585
R691 B.n385 B.n384 585
R692 B.n386 B.n203 585
R693 B.n388 B.n387 585
R694 B.n389 B.n202 585
R695 B.n391 B.n390 585
R696 B.n392 B.n201 585
R697 B.n394 B.n393 585
R698 B.n395 B.n200 585
R699 B.n397 B.n396 585
R700 B.n398 B.n199 585
R701 B.n400 B.n399 585
R702 B.n401 B.n198 585
R703 B.n403 B.n402 585
R704 B.n404 B.n197 585
R705 B.n406 B.n405 585
R706 B.n407 B.n196 585
R707 B.n409 B.n408 585
R708 B.n410 B.n195 585
R709 B.n412 B.n411 585
R710 B.n413 B.n194 585
R711 B.n415 B.n414 585
R712 B.n416 B.n193 585
R713 B.n418 B.n417 585
R714 B.n420 B.n419 585
R715 B.n421 B.n189 585
R716 B.n423 B.n422 585
R717 B.n424 B.n188 585
R718 B.n426 B.n425 585
R719 B.n427 B.n187 585
R720 B.n429 B.n428 585
R721 B.n430 B.n186 585
R722 B.n432 B.n431 585
R723 B.n433 B.n183 585
R724 B.n436 B.n435 585
R725 B.n437 B.n182 585
R726 B.n439 B.n438 585
R727 B.n440 B.n181 585
R728 B.n442 B.n441 585
R729 B.n443 B.n180 585
R730 B.n445 B.n444 585
R731 B.n446 B.n179 585
R732 B.n448 B.n447 585
R733 B.n449 B.n178 585
R734 B.n451 B.n450 585
R735 B.n452 B.n177 585
R736 B.n454 B.n453 585
R737 B.n455 B.n176 585
R738 B.n457 B.n456 585
R739 B.n458 B.n175 585
R740 B.n460 B.n459 585
R741 B.n461 B.n174 585
R742 B.n463 B.n462 585
R743 B.n464 B.n173 585
R744 B.n466 B.n465 585
R745 B.n467 B.n172 585
R746 B.n469 B.n468 585
R747 B.n470 B.n171 585
R748 B.n472 B.n471 585
R749 B.n473 B.n170 585
R750 B.n475 B.n474 585
R751 B.n476 B.n169 585
R752 B.n478 B.n477 585
R753 B.n479 B.n168 585
R754 B.n481 B.n480 585
R755 B.n482 B.n167 585
R756 B.n484 B.n483 585
R757 B.n485 B.n166 585
R758 B.n487 B.n486 585
R759 B.n488 B.n165 585
R760 B.n490 B.n489 585
R761 B.n362 B.n211 585
R762 B.n361 B.n360 585
R763 B.n359 B.n212 585
R764 B.n358 B.n357 585
R765 B.n356 B.n213 585
R766 B.n355 B.n354 585
R767 B.n353 B.n214 585
R768 B.n352 B.n351 585
R769 B.n350 B.n215 585
R770 B.n349 B.n348 585
R771 B.n347 B.n216 585
R772 B.n346 B.n345 585
R773 B.n344 B.n217 585
R774 B.n343 B.n342 585
R775 B.n341 B.n218 585
R776 B.n340 B.n339 585
R777 B.n338 B.n219 585
R778 B.n337 B.n336 585
R779 B.n335 B.n220 585
R780 B.n334 B.n333 585
R781 B.n332 B.n221 585
R782 B.n331 B.n330 585
R783 B.n329 B.n222 585
R784 B.n328 B.n327 585
R785 B.n326 B.n223 585
R786 B.n325 B.n324 585
R787 B.n323 B.n224 585
R788 B.n322 B.n321 585
R789 B.n320 B.n225 585
R790 B.n319 B.n318 585
R791 B.n317 B.n226 585
R792 B.n316 B.n315 585
R793 B.n314 B.n227 585
R794 B.n313 B.n312 585
R795 B.n311 B.n228 585
R796 B.n310 B.n309 585
R797 B.n308 B.n229 585
R798 B.n307 B.n306 585
R799 B.n305 B.n230 585
R800 B.n304 B.n303 585
R801 B.n302 B.n231 585
R802 B.n301 B.n300 585
R803 B.n299 B.n232 585
R804 B.n298 B.n297 585
R805 B.n296 B.n233 585
R806 B.n295 B.n294 585
R807 B.n293 B.n234 585
R808 B.n292 B.n291 585
R809 B.n290 B.n235 585
R810 B.n289 B.n288 585
R811 B.n287 B.n236 585
R812 B.n286 B.n285 585
R813 B.n284 B.n237 585
R814 B.n283 B.n282 585
R815 B.n281 B.n238 585
R816 B.n280 B.n279 585
R817 B.n278 B.n239 585
R818 B.n277 B.n276 585
R819 B.n275 B.n240 585
R820 B.n274 B.n273 585
R821 B.n272 B.n241 585
R822 B.n271 B.n270 585
R823 B.n269 B.n242 585
R824 B.n268 B.n267 585
R825 B.n266 B.n243 585
R826 B.n265 B.n264 585
R827 B.n263 B.n244 585
R828 B.n262 B.n261 585
R829 B.n260 B.n245 585
R830 B.n259 B.n258 585
R831 B.n257 B.n246 585
R832 B.n256 B.n255 585
R833 B.n254 B.n247 585
R834 B.n253 B.n252 585
R835 B.n251 B.n248 585
R836 B.n250 B.n249 585
R837 B.n2 B.n0 585
R838 B.n965 B.n1 585
R839 B.n964 B.n963 585
R840 B.n962 B.n3 585
R841 B.n961 B.n960 585
R842 B.n959 B.n4 585
R843 B.n958 B.n957 585
R844 B.n956 B.n5 585
R845 B.n955 B.n954 585
R846 B.n953 B.n6 585
R847 B.n952 B.n951 585
R848 B.n950 B.n7 585
R849 B.n949 B.n948 585
R850 B.n947 B.n8 585
R851 B.n946 B.n945 585
R852 B.n944 B.n9 585
R853 B.n943 B.n942 585
R854 B.n941 B.n10 585
R855 B.n940 B.n939 585
R856 B.n938 B.n11 585
R857 B.n937 B.n936 585
R858 B.n935 B.n12 585
R859 B.n934 B.n933 585
R860 B.n932 B.n13 585
R861 B.n931 B.n930 585
R862 B.n929 B.n14 585
R863 B.n928 B.n927 585
R864 B.n926 B.n15 585
R865 B.n925 B.n924 585
R866 B.n923 B.n16 585
R867 B.n922 B.n921 585
R868 B.n920 B.n17 585
R869 B.n919 B.n918 585
R870 B.n917 B.n18 585
R871 B.n916 B.n915 585
R872 B.n914 B.n19 585
R873 B.n913 B.n912 585
R874 B.n911 B.n20 585
R875 B.n910 B.n909 585
R876 B.n908 B.n21 585
R877 B.n907 B.n906 585
R878 B.n905 B.n22 585
R879 B.n904 B.n903 585
R880 B.n902 B.n23 585
R881 B.n901 B.n900 585
R882 B.n899 B.n24 585
R883 B.n898 B.n897 585
R884 B.n896 B.n25 585
R885 B.n895 B.n894 585
R886 B.n893 B.n26 585
R887 B.n892 B.n891 585
R888 B.n890 B.n27 585
R889 B.n889 B.n888 585
R890 B.n887 B.n28 585
R891 B.n886 B.n885 585
R892 B.n884 B.n29 585
R893 B.n883 B.n882 585
R894 B.n881 B.n30 585
R895 B.n880 B.n879 585
R896 B.n878 B.n31 585
R897 B.n877 B.n876 585
R898 B.n875 B.n32 585
R899 B.n874 B.n873 585
R900 B.n872 B.n33 585
R901 B.n871 B.n870 585
R902 B.n869 B.n34 585
R903 B.n868 B.n867 585
R904 B.n866 B.n35 585
R905 B.n865 B.n864 585
R906 B.n863 B.n36 585
R907 B.n862 B.n861 585
R908 B.n860 B.n37 585
R909 B.n859 B.n858 585
R910 B.n857 B.n38 585
R911 B.n856 B.n855 585
R912 B.n854 B.n39 585
R913 B.n853 B.n852 585
R914 B.n851 B.n40 585
R915 B.n967 B.n966 585
R916 B.n364 B.n211 506.916
R917 B.n851 B.n850 506.916
R918 B.n491 B.n490 506.916
R919 B.n724 B.n87 506.916
R920 B.n184 B.t9 280.308
R921 B.n190 B.t3 280.308
R922 B.n60 B.t0 280.308
R923 B.n66 B.t6 280.308
R924 B.n184 B.t11 189.731
R925 B.n66 B.t7 189.731
R926 B.n190 B.t5 189.719
R927 B.n60 B.t1 189.719
R928 B.n360 B.n211 163.367
R929 B.n360 B.n359 163.367
R930 B.n359 B.n358 163.367
R931 B.n358 B.n213 163.367
R932 B.n354 B.n213 163.367
R933 B.n354 B.n353 163.367
R934 B.n353 B.n352 163.367
R935 B.n352 B.n215 163.367
R936 B.n348 B.n215 163.367
R937 B.n348 B.n347 163.367
R938 B.n347 B.n346 163.367
R939 B.n346 B.n217 163.367
R940 B.n342 B.n217 163.367
R941 B.n342 B.n341 163.367
R942 B.n341 B.n340 163.367
R943 B.n340 B.n219 163.367
R944 B.n336 B.n219 163.367
R945 B.n336 B.n335 163.367
R946 B.n335 B.n334 163.367
R947 B.n334 B.n221 163.367
R948 B.n330 B.n221 163.367
R949 B.n330 B.n329 163.367
R950 B.n329 B.n328 163.367
R951 B.n328 B.n223 163.367
R952 B.n324 B.n223 163.367
R953 B.n324 B.n323 163.367
R954 B.n323 B.n322 163.367
R955 B.n322 B.n225 163.367
R956 B.n318 B.n225 163.367
R957 B.n318 B.n317 163.367
R958 B.n317 B.n316 163.367
R959 B.n316 B.n227 163.367
R960 B.n312 B.n227 163.367
R961 B.n312 B.n311 163.367
R962 B.n311 B.n310 163.367
R963 B.n310 B.n229 163.367
R964 B.n306 B.n229 163.367
R965 B.n306 B.n305 163.367
R966 B.n305 B.n304 163.367
R967 B.n304 B.n231 163.367
R968 B.n300 B.n231 163.367
R969 B.n300 B.n299 163.367
R970 B.n299 B.n298 163.367
R971 B.n298 B.n233 163.367
R972 B.n294 B.n233 163.367
R973 B.n294 B.n293 163.367
R974 B.n293 B.n292 163.367
R975 B.n292 B.n235 163.367
R976 B.n288 B.n235 163.367
R977 B.n288 B.n287 163.367
R978 B.n287 B.n286 163.367
R979 B.n286 B.n237 163.367
R980 B.n282 B.n237 163.367
R981 B.n282 B.n281 163.367
R982 B.n281 B.n280 163.367
R983 B.n280 B.n239 163.367
R984 B.n276 B.n239 163.367
R985 B.n276 B.n275 163.367
R986 B.n275 B.n274 163.367
R987 B.n274 B.n241 163.367
R988 B.n270 B.n241 163.367
R989 B.n270 B.n269 163.367
R990 B.n269 B.n268 163.367
R991 B.n268 B.n243 163.367
R992 B.n264 B.n243 163.367
R993 B.n264 B.n263 163.367
R994 B.n263 B.n262 163.367
R995 B.n262 B.n245 163.367
R996 B.n258 B.n245 163.367
R997 B.n258 B.n257 163.367
R998 B.n257 B.n256 163.367
R999 B.n256 B.n247 163.367
R1000 B.n252 B.n247 163.367
R1001 B.n252 B.n251 163.367
R1002 B.n251 B.n250 163.367
R1003 B.n250 B.n2 163.367
R1004 B.n966 B.n2 163.367
R1005 B.n966 B.n965 163.367
R1006 B.n965 B.n964 163.367
R1007 B.n964 B.n3 163.367
R1008 B.n960 B.n3 163.367
R1009 B.n960 B.n959 163.367
R1010 B.n959 B.n958 163.367
R1011 B.n958 B.n5 163.367
R1012 B.n954 B.n5 163.367
R1013 B.n954 B.n953 163.367
R1014 B.n953 B.n952 163.367
R1015 B.n952 B.n7 163.367
R1016 B.n948 B.n7 163.367
R1017 B.n948 B.n947 163.367
R1018 B.n947 B.n946 163.367
R1019 B.n946 B.n9 163.367
R1020 B.n942 B.n9 163.367
R1021 B.n942 B.n941 163.367
R1022 B.n941 B.n940 163.367
R1023 B.n940 B.n11 163.367
R1024 B.n936 B.n11 163.367
R1025 B.n936 B.n935 163.367
R1026 B.n935 B.n934 163.367
R1027 B.n934 B.n13 163.367
R1028 B.n930 B.n13 163.367
R1029 B.n930 B.n929 163.367
R1030 B.n929 B.n928 163.367
R1031 B.n928 B.n15 163.367
R1032 B.n924 B.n15 163.367
R1033 B.n924 B.n923 163.367
R1034 B.n923 B.n922 163.367
R1035 B.n922 B.n17 163.367
R1036 B.n918 B.n17 163.367
R1037 B.n918 B.n917 163.367
R1038 B.n917 B.n916 163.367
R1039 B.n916 B.n19 163.367
R1040 B.n912 B.n19 163.367
R1041 B.n912 B.n911 163.367
R1042 B.n911 B.n910 163.367
R1043 B.n910 B.n21 163.367
R1044 B.n906 B.n21 163.367
R1045 B.n906 B.n905 163.367
R1046 B.n905 B.n904 163.367
R1047 B.n904 B.n23 163.367
R1048 B.n900 B.n23 163.367
R1049 B.n900 B.n899 163.367
R1050 B.n899 B.n898 163.367
R1051 B.n898 B.n25 163.367
R1052 B.n894 B.n25 163.367
R1053 B.n894 B.n893 163.367
R1054 B.n893 B.n892 163.367
R1055 B.n892 B.n27 163.367
R1056 B.n888 B.n27 163.367
R1057 B.n888 B.n887 163.367
R1058 B.n887 B.n886 163.367
R1059 B.n886 B.n29 163.367
R1060 B.n882 B.n29 163.367
R1061 B.n882 B.n881 163.367
R1062 B.n881 B.n880 163.367
R1063 B.n880 B.n31 163.367
R1064 B.n876 B.n31 163.367
R1065 B.n876 B.n875 163.367
R1066 B.n875 B.n874 163.367
R1067 B.n874 B.n33 163.367
R1068 B.n870 B.n33 163.367
R1069 B.n870 B.n869 163.367
R1070 B.n869 B.n868 163.367
R1071 B.n868 B.n35 163.367
R1072 B.n864 B.n35 163.367
R1073 B.n864 B.n863 163.367
R1074 B.n863 B.n862 163.367
R1075 B.n862 B.n37 163.367
R1076 B.n858 B.n37 163.367
R1077 B.n858 B.n857 163.367
R1078 B.n857 B.n856 163.367
R1079 B.n856 B.n39 163.367
R1080 B.n852 B.n39 163.367
R1081 B.n852 B.n851 163.367
R1082 B.n365 B.n364 163.367
R1083 B.n366 B.n365 163.367
R1084 B.n366 B.n209 163.367
R1085 B.n370 B.n209 163.367
R1086 B.n371 B.n370 163.367
R1087 B.n372 B.n371 163.367
R1088 B.n372 B.n207 163.367
R1089 B.n376 B.n207 163.367
R1090 B.n377 B.n376 163.367
R1091 B.n378 B.n377 163.367
R1092 B.n378 B.n205 163.367
R1093 B.n382 B.n205 163.367
R1094 B.n383 B.n382 163.367
R1095 B.n384 B.n383 163.367
R1096 B.n384 B.n203 163.367
R1097 B.n388 B.n203 163.367
R1098 B.n389 B.n388 163.367
R1099 B.n390 B.n389 163.367
R1100 B.n390 B.n201 163.367
R1101 B.n394 B.n201 163.367
R1102 B.n395 B.n394 163.367
R1103 B.n396 B.n395 163.367
R1104 B.n396 B.n199 163.367
R1105 B.n400 B.n199 163.367
R1106 B.n401 B.n400 163.367
R1107 B.n402 B.n401 163.367
R1108 B.n402 B.n197 163.367
R1109 B.n406 B.n197 163.367
R1110 B.n407 B.n406 163.367
R1111 B.n408 B.n407 163.367
R1112 B.n408 B.n195 163.367
R1113 B.n412 B.n195 163.367
R1114 B.n413 B.n412 163.367
R1115 B.n414 B.n413 163.367
R1116 B.n414 B.n193 163.367
R1117 B.n418 B.n193 163.367
R1118 B.n419 B.n418 163.367
R1119 B.n419 B.n189 163.367
R1120 B.n423 B.n189 163.367
R1121 B.n424 B.n423 163.367
R1122 B.n425 B.n424 163.367
R1123 B.n425 B.n187 163.367
R1124 B.n429 B.n187 163.367
R1125 B.n430 B.n429 163.367
R1126 B.n431 B.n430 163.367
R1127 B.n431 B.n183 163.367
R1128 B.n436 B.n183 163.367
R1129 B.n437 B.n436 163.367
R1130 B.n438 B.n437 163.367
R1131 B.n438 B.n181 163.367
R1132 B.n442 B.n181 163.367
R1133 B.n443 B.n442 163.367
R1134 B.n444 B.n443 163.367
R1135 B.n444 B.n179 163.367
R1136 B.n448 B.n179 163.367
R1137 B.n449 B.n448 163.367
R1138 B.n450 B.n449 163.367
R1139 B.n450 B.n177 163.367
R1140 B.n454 B.n177 163.367
R1141 B.n455 B.n454 163.367
R1142 B.n456 B.n455 163.367
R1143 B.n456 B.n175 163.367
R1144 B.n460 B.n175 163.367
R1145 B.n461 B.n460 163.367
R1146 B.n462 B.n461 163.367
R1147 B.n462 B.n173 163.367
R1148 B.n466 B.n173 163.367
R1149 B.n467 B.n466 163.367
R1150 B.n468 B.n467 163.367
R1151 B.n468 B.n171 163.367
R1152 B.n472 B.n171 163.367
R1153 B.n473 B.n472 163.367
R1154 B.n474 B.n473 163.367
R1155 B.n474 B.n169 163.367
R1156 B.n478 B.n169 163.367
R1157 B.n479 B.n478 163.367
R1158 B.n480 B.n479 163.367
R1159 B.n480 B.n167 163.367
R1160 B.n484 B.n167 163.367
R1161 B.n485 B.n484 163.367
R1162 B.n486 B.n485 163.367
R1163 B.n486 B.n165 163.367
R1164 B.n490 B.n165 163.367
R1165 B.n492 B.n491 163.367
R1166 B.n492 B.n163 163.367
R1167 B.n496 B.n163 163.367
R1168 B.n497 B.n496 163.367
R1169 B.n498 B.n497 163.367
R1170 B.n498 B.n161 163.367
R1171 B.n502 B.n161 163.367
R1172 B.n503 B.n502 163.367
R1173 B.n504 B.n503 163.367
R1174 B.n504 B.n159 163.367
R1175 B.n508 B.n159 163.367
R1176 B.n509 B.n508 163.367
R1177 B.n510 B.n509 163.367
R1178 B.n510 B.n157 163.367
R1179 B.n514 B.n157 163.367
R1180 B.n515 B.n514 163.367
R1181 B.n516 B.n515 163.367
R1182 B.n516 B.n155 163.367
R1183 B.n520 B.n155 163.367
R1184 B.n521 B.n520 163.367
R1185 B.n522 B.n521 163.367
R1186 B.n522 B.n153 163.367
R1187 B.n526 B.n153 163.367
R1188 B.n527 B.n526 163.367
R1189 B.n528 B.n527 163.367
R1190 B.n528 B.n151 163.367
R1191 B.n532 B.n151 163.367
R1192 B.n533 B.n532 163.367
R1193 B.n534 B.n533 163.367
R1194 B.n534 B.n149 163.367
R1195 B.n538 B.n149 163.367
R1196 B.n539 B.n538 163.367
R1197 B.n540 B.n539 163.367
R1198 B.n540 B.n147 163.367
R1199 B.n544 B.n147 163.367
R1200 B.n545 B.n544 163.367
R1201 B.n546 B.n545 163.367
R1202 B.n546 B.n145 163.367
R1203 B.n550 B.n145 163.367
R1204 B.n551 B.n550 163.367
R1205 B.n552 B.n551 163.367
R1206 B.n552 B.n143 163.367
R1207 B.n556 B.n143 163.367
R1208 B.n557 B.n556 163.367
R1209 B.n558 B.n557 163.367
R1210 B.n558 B.n141 163.367
R1211 B.n562 B.n141 163.367
R1212 B.n563 B.n562 163.367
R1213 B.n564 B.n563 163.367
R1214 B.n564 B.n139 163.367
R1215 B.n568 B.n139 163.367
R1216 B.n569 B.n568 163.367
R1217 B.n570 B.n569 163.367
R1218 B.n570 B.n137 163.367
R1219 B.n574 B.n137 163.367
R1220 B.n575 B.n574 163.367
R1221 B.n576 B.n575 163.367
R1222 B.n576 B.n135 163.367
R1223 B.n580 B.n135 163.367
R1224 B.n581 B.n580 163.367
R1225 B.n582 B.n581 163.367
R1226 B.n582 B.n133 163.367
R1227 B.n586 B.n133 163.367
R1228 B.n587 B.n586 163.367
R1229 B.n588 B.n587 163.367
R1230 B.n588 B.n131 163.367
R1231 B.n592 B.n131 163.367
R1232 B.n593 B.n592 163.367
R1233 B.n594 B.n593 163.367
R1234 B.n594 B.n129 163.367
R1235 B.n598 B.n129 163.367
R1236 B.n599 B.n598 163.367
R1237 B.n600 B.n599 163.367
R1238 B.n600 B.n127 163.367
R1239 B.n604 B.n127 163.367
R1240 B.n605 B.n604 163.367
R1241 B.n606 B.n605 163.367
R1242 B.n606 B.n125 163.367
R1243 B.n610 B.n125 163.367
R1244 B.n611 B.n610 163.367
R1245 B.n612 B.n611 163.367
R1246 B.n612 B.n123 163.367
R1247 B.n616 B.n123 163.367
R1248 B.n617 B.n616 163.367
R1249 B.n618 B.n617 163.367
R1250 B.n618 B.n121 163.367
R1251 B.n622 B.n121 163.367
R1252 B.n623 B.n622 163.367
R1253 B.n624 B.n623 163.367
R1254 B.n624 B.n119 163.367
R1255 B.n628 B.n119 163.367
R1256 B.n629 B.n628 163.367
R1257 B.n630 B.n629 163.367
R1258 B.n630 B.n117 163.367
R1259 B.n634 B.n117 163.367
R1260 B.n635 B.n634 163.367
R1261 B.n636 B.n635 163.367
R1262 B.n636 B.n115 163.367
R1263 B.n640 B.n115 163.367
R1264 B.n641 B.n640 163.367
R1265 B.n642 B.n641 163.367
R1266 B.n642 B.n113 163.367
R1267 B.n646 B.n113 163.367
R1268 B.n647 B.n646 163.367
R1269 B.n648 B.n647 163.367
R1270 B.n648 B.n111 163.367
R1271 B.n652 B.n111 163.367
R1272 B.n653 B.n652 163.367
R1273 B.n654 B.n653 163.367
R1274 B.n654 B.n109 163.367
R1275 B.n658 B.n109 163.367
R1276 B.n659 B.n658 163.367
R1277 B.n660 B.n659 163.367
R1278 B.n660 B.n107 163.367
R1279 B.n664 B.n107 163.367
R1280 B.n665 B.n664 163.367
R1281 B.n666 B.n665 163.367
R1282 B.n666 B.n105 163.367
R1283 B.n670 B.n105 163.367
R1284 B.n671 B.n670 163.367
R1285 B.n672 B.n671 163.367
R1286 B.n672 B.n103 163.367
R1287 B.n676 B.n103 163.367
R1288 B.n677 B.n676 163.367
R1289 B.n678 B.n677 163.367
R1290 B.n678 B.n101 163.367
R1291 B.n682 B.n101 163.367
R1292 B.n683 B.n682 163.367
R1293 B.n684 B.n683 163.367
R1294 B.n684 B.n99 163.367
R1295 B.n688 B.n99 163.367
R1296 B.n689 B.n688 163.367
R1297 B.n690 B.n689 163.367
R1298 B.n690 B.n97 163.367
R1299 B.n694 B.n97 163.367
R1300 B.n695 B.n694 163.367
R1301 B.n696 B.n695 163.367
R1302 B.n696 B.n95 163.367
R1303 B.n700 B.n95 163.367
R1304 B.n701 B.n700 163.367
R1305 B.n702 B.n701 163.367
R1306 B.n702 B.n93 163.367
R1307 B.n706 B.n93 163.367
R1308 B.n707 B.n706 163.367
R1309 B.n708 B.n707 163.367
R1310 B.n708 B.n91 163.367
R1311 B.n712 B.n91 163.367
R1312 B.n713 B.n712 163.367
R1313 B.n714 B.n713 163.367
R1314 B.n714 B.n89 163.367
R1315 B.n718 B.n89 163.367
R1316 B.n719 B.n718 163.367
R1317 B.n720 B.n719 163.367
R1318 B.n720 B.n87 163.367
R1319 B.n850 B.n41 163.367
R1320 B.n846 B.n41 163.367
R1321 B.n846 B.n845 163.367
R1322 B.n845 B.n844 163.367
R1323 B.n844 B.n43 163.367
R1324 B.n840 B.n43 163.367
R1325 B.n840 B.n839 163.367
R1326 B.n839 B.n838 163.367
R1327 B.n838 B.n45 163.367
R1328 B.n834 B.n45 163.367
R1329 B.n834 B.n833 163.367
R1330 B.n833 B.n832 163.367
R1331 B.n832 B.n47 163.367
R1332 B.n828 B.n47 163.367
R1333 B.n828 B.n827 163.367
R1334 B.n827 B.n826 163.367
R1335 B.n826 B.n49 163.367
R1336 B.n822 B.n49 163.367
R1337 B.n822 B.n821 163.367
R1338 B.n821 B.n820 163.367
R1339 B.n820 B.n51 163.367
R1340 B.n816 B.n51 163.367
R1341 B.n816 B.n815 163.367
R1342 B.n815 B.n814 163.367
R1343 B.n814 B.n53 163.367
R1344 B.n810 B.n53 163.367
R1345 B.n810 B.n809 163.367
R1346 B.n809 B.n808 163.367
R1347 B.n808 B.n55 163.367
R1348 B.n804 B.n55 163.367
R1349 B.n804 B.n803 163.367
R1350 B.n803 B.n802 163.367
R1351 B.n802 B.n57 163.367
R1352 B.n798 B.n57 163.367
R1353 B.n798 B.n797 163.367
R1354 B.n797 B.n796 163.367
R1355 B.n796 B.n59 163.367
R1356 B.n791 B.n59 163.367
R1357 B.n791 B.n790 163.367
R1358 B.n790 B.n789 163.367
R1359 B.n789 B.n63 163.367
R1360 B.n785 B.n63 163.367
R1361 B.n785 B.n784 163.367
R1362 B.n784 B.n783 163.367
R1363 B.n783 B.n65 163.367
R1364 B.n779 B.n65 163.367
R1365 B.n779 B.n778 163.367
R1366 B.n778 B.n69 163.367
R1367 B.n774 B.n69 163.367
R1368 B.n774 B.n773 163.367
R1369 B.n773 B.n772 163.367
R1370 B.n772 B.n71 163.367
R1371 B.n768 B.n71 163.367
R1372 B.n768 B.n767 163.367
R1373 B.n767 B.n766 163.367
R1374 B.n766 B.n73 163.367
R1375 B.n762 B.n73 163.367
R1376 B.n762 B.n761 163.367
R1377 B.n761 B.n760 163.367
R1378 B.n760 B.n75 163.367
R1379 B.n756 B.n75 163.367
R1380 B.n756 B.n755 163.367
R1381 B.n755 B.n754 163.367
R1382 B.n754 B.n77 163.367
R1383 B.n750 B.n77 163.367
R1384 B.n750 B.n749 163.367
R1385 B.n749 B.n748 163.367
R1386 B.n748 B.n79 163.367
R1387 B.n744 B.n79 163.367
R1388 B.n744 B.n743 163.367
R1389 B.n743 B.n742 163.367
R1390 B.n742 B.n81 163.367
R1391 B.n738 B.n81 163.367
R1392 B.n738 B.n737 163.367
R1393 B.n737 B.n736 163.367
R1394 B.n736 B.n83 163.367
R1395 B.n732 B.n83 163.367
R1396 B.n732 B.n731 163.367
R1397 B.n731 B.n730 163.367
R1398 B.n730 B.n85 163.367
R1399 B.n726 B.n85 163.367
R1400 B.n726 B.n725 163.367
R1401 B.n725 B.n724 163.367
R1402 B.n185 B.t10 114.094
R1403 B.n67 B.t8 114.094
R1404 B.n191 B.t4 114.082
R1405 B.n61 B.t2 114.082
R1406 B.n185 B.n184 75.6369
R1407 B.n191 B.n190 75.6369
R1408 B.n61 B.n60 75.6369
R1409 B.n67 B.n66 75.6369
R1410 B.n434 B.n185 59.5399
R1411 B.n192 B.n191 59.5399
R1412 B.n794 B.n61 59.5399
R1413 B.n68 B.n67 59.5399
R1414 B.n849 B.n40 32.9371
R1415 B.n723 B.n722 32.9371
R1416 B.n489 B.n164 32.9371
R1417 B.n363 B.n362 32.9371
R1418 B B.n967 18.0485
R1419 B.n849 B.n848 10.6151
R1420 B.n848 B.n847 10.6151
R1421 B.n847 B.n42 10.6151
R1422 B.n843 B.n42 10.6151
R1423 B.n843 B.n842 10.6151
R1424 B.n842 B.n841 10.6151
R1425 B.n841 B.n44 10.6151
R1426 B.n837 B.n44 10.6151
R1427 B.n837 B.n836 10.6151
R1428 B.n836 B.n835 10.6151
R1429 B.n835 B.n46 10.6151
R1430 B.n831 B.n46 10.6151
R1431 B.n831 B.n830 10.6151
R1432 B.n830 B.n829 10.6151
R1433 B.n829 B.n48 10.6151
R1434 B.n825 B.n48 10.6151
R1435 B.n825 B.n824 10.6151
R1436 B.n824 B.n823 10.6151
R1437 B.n823 B.n50 10.6151
R1438 B.n819 B.n50 10.6151
R1439 B.n819 B.n818 10.6151
R1440 B.n818 B.n817 10.6151
R1441 B.n817 B.n52 10.6151
R1442 B.n813 B.n52 10.6151
R1443 B.n813 B.n812 10.6151
R1444 B.n812 B.n811 10.6151
R1445 B.n811 B.n54 10.6151
R1446 B.n807 B.n54 10.6151
R1447 B.n807 B.n806 10.6151
R1448 B.n806 B.n805 10.6151
R1449 B.n805 B.n56 10.6151
R1450 B.n801 B.n56 10.6151
R1451 B.n801 B.n800 10.6151
R1452 B.n800 B.n799 10.6151
R1453 B.n799 B.n58 10.6151
R1454 B.n795 B.n58 10.6151
R1455 B.n793 B.n792 10.6151
R1456 B.n792 B.n62 10.6151
R1457 B.n788 B.n62 10.6151
R1458 B.n788 B.n787 10.6151
R1459 B.n787 B.n786 10.6151
R1460 B.n786 B.n64 10.6151
R1461 B.n782 B.n64 10.6151
R1462 B.n782 B.n781 10.6151
R1463 B.n781 B.n780 10.6151
R1464 B.n777 B.n776 10.6151
R1465 B.n776 B.n775 10.6151
R1466 B.n775 B.n70 10.6151
R1467 B.n771 B.n70 10.6151
R1468 B.n771 B.n770 10.6151
R1469 B.n770 B.n769 10.6151
R1470 B.n769 B.n72 10.6151
R1471 B.n765 B.n72 10.6151
R1472 B.n765 B.n764 10.6151
R1473 B.n764 B.n763 10.6151
R1474 B.n763 B.n74 10.6151
R1475 B.n759 B.n74 10.6151
R1476 B.n759 B.n758 10.6151
R1477 B.n758 B.n757 10.6151
R1478 B.n757 B.n76 10.6151
R1479 B.n753 B.n76 10.6151
R1480 B.n753 B.n752 10.6151
R1481 B.n752 B.n751 10.6151
R1482 B.n751 B.n78 10.6151
R1483 B.n747 B.n78 10.6151
R1484 B.n747 B.n746 10.6151
R1485 B.n746 B.n745 10.6151
R1486 B.n745 B.n80 10.6151
R1487 B.n741 B.n80 10.6151
R1488 B.n741 B.n740 10.6151
R1489 B.n740 B.n739 10.6151
R1490 B.n739 B.n82 10.6151
R1491 B.n735 B.n82 10.6151
R1492 B.n735 B.n734 10.6151
R1493 B.n734 B.n733 10.6151
R1494 B.n733 B.n84 10.6151
R1495 B.n729 B.n84 10.6151
R1496 B.n729 B.n728 10.6151
R1497 B.n728 B.n727 10.6151
R1498 B.n727 B.n86 10.6151
R1499 B.n723 B.n86 10.6151
R1500 B.n493 B.n164 10.6151
R1501 B.n494 B.n493 10.6151
R1502 B.n495 B.n494 10.6151
R1503 B.n495 B.n162 10.6151
R1504 B.n499 B.n162 10.6151
R1505 B.n500 B.n499 10.6151
R1506 B.n501 B.n500 10.6151
R1507 B.n501 B.n160 10.6151
R1508 B.n505 B.n160 10.6151
R1509 B.n506 B.n505 10.6151
R1510 B.n507 B.n506 10.6151
R1511 B.n507 B.n158 10.6151
R1512 B.n511 B.n158 10.6151
R1513 B.n512 B.n511 10.6151
R1514 B.n513 B.n512 10.6151
R1515 B.n513 B.n156 10.6151
R1516 B.n517 B.n156 10.6151
R1517 B.n518 B.n517 10.6151
R1518 B.n519 B.n518 10.6151
R1519 B.n519 B.n154 10.6151
R1520 B.n523 B.n154 10.6151
R1521 B.n524 B.n523 10.6151
R1522 B.n525 B.n524 10.6151
R1523 B.n525 B.n152 10.6151
R1524 B.n529 B.n152 10.6151
R1525 B.n530 B.n529 10.6151
R1526 B.n531 B.n530 10.6151
R1527 B.n531 B.n150 10.6151
R1528 B.n535 B.n150 10.6151
R1529 B.n536 B.n535 10.6151
R1530 B.n537 B.n536 10.6151
R1531 B.n537 B.n148 10.6151
R1532 B.n541 B.n148 10.6151
R1533 B.n542 B.n541 10.6151
R1534 B.n543 B.n542 10.6151
R1535 B.n543 B.n146 10.6151
R1536 B.n547 B.n146 10.6151
R1537 B.n548 B.n547 10.6151
R1538 B.n549 B.n548 10.6151
R1539 B.n549 B.n144 10.6151
R1540 B.n553 B.n144 10.6151
R1541 B.n554 B.n553 10.6151
R1542 B.n555 B.n554 10.6151
R1543 B.n555 B.n142 10.6151
R1544 B.n559 B.n142 10.6151
R1545 B.n560 B.n559 10.6151
R1546 B.n561 B.n560 10.6151
R1547 B.n561 B.n140 10.6151
R1548 B.n565 B.n140 10.6151
R1549 B.n566 B.n565 10.6151
R1550 B.n567 B.n566 10.6151
R1551 B.n567 B.n138 10.6151
R1552 B.n571 B.n138 10.6151
R1553 B.n572 B.n571 10.6151
R1554 B.n573 B.n572 10.6151
R1555 B.n573 B.n136 10.6151
R1556 B.n577 B.n136 10.6151
R1557 B.n578 B.n577 10.6151
R1558 B.n579 B.n578 10.6151
R1559 B.n579 B.n134 10.6151
R1560 B.n583 B.n134 10.6151
R1561 B.n584 B.n583 10.6151
R1562 B.n585 B.n584 10.6151
R1563 B.n585 B.n132 10.6151
R1564 B.n589 B.n132 10.6151
R1565 B.n590 B.n589 10.6151
R1566 B.n591 B.n590 10.6151
R1567 B.n591 B.n130 10.6151
R1568 B.n595 B.n130 10.6151
R1569 B.n596 B.n595 10.6151
R1570 B.n597 B.n596 10.6151
R1571 B.n597 B.n128 10.6151
R1572 B.n601 B.n128 10.6151
R1573 B.n602 B.n601 10.6151
R1574 B.n603 B.n602 10.6151
R1575 B.n603 B.n126 10.6151
R1576 B.n607 B.n126 10.6151
R1577 B.n608 B.n607 10.6151
R1578 B.n609 B.n608 10.6151
R1579 B.n609 B.n124 10.6151
R1580 B.n613 B.n124 10.6151
R1581 B.n614 B.n613 10.6151
R1582 B.n615 B.n614 10.6151
R1583 B.n615 B.n122 10.6151
R1584 B.n619 B.n122 10.6151
R1585 B.n620 B.n619 10.6151
R1586 B.n621 B.n620 10.6151
R1587 B.n621 B.n120 10.6151
R1588 B.n625 B.n120 10.6151
R1589 B.n626 B.n625 10.6151
R1590 B.n627 B.n626 10.6151
R1591 B.n627 B.n118 10.6151
R1592 B.n631 B.n118 10.6151
R1593 B.n632 B.n631 10.6151
R1594 B.n633 B.n632 10.6151
R1595 B.n633 B.n116 10.6151
R1596 B.n637 B.n116 10.6151
R1597 B.n638 B.n637 10.6151
R1598 B.n639 B.n638 10.6151
R1599 B.n639 B.n114 10.6151
R1600 B.n643 B.n114 10.6151
R1601 B.n644 B.n643 10.6151
R1602 B.n645 B.n644 10.6151
R1603 B.n645 B.n112 10.6151
R1604 B.n649 B.n112 10.6151
R1605 B.n650 B.n649 10.6151
R1606 B.n651 B.n650 10.6151
R1607 B.n651 B.n110 10.6151
R1608 B.n655 B.n110 10.6151
R1609 B.n656 B.n655 10.6151
R1610 B.n657 B.n656 10.6151
R1611 B.n657 B.n108 10.6151
R1612 B.n661 B.n108 10.6151
R1613 B.n662 B.n661 10.6151
R1614 B.n663 B.n662 10.6151
R1615 B.n663 B.n106 10.6151
R1616 B.n667 B.n106 10.6151
R1617 B.n668 B.n667 10.6151
R1618 B.n669 B.n668 10.6151
R1619 B.n669 B.n104 10.6151
R1620 B.n673 B.n104 10.6151
R1621 B.n674 B.n673 10.6151
R1622 B.n675 B.n674 10.6151
R1623 B.n675 B.n102 10.6151
R1624 B.n679 B.n102 10.6151
R1625 B.n680 B.n679 10.6151
R1626 B.n681 B.n680 10.6151
R1627 B.n681 B.n100 10.6151
R1628 B.n685 B.n100 10.6151
R1629 B.n686 B.n685 10.6151
R1630 B.n687 B.n686 10.6151
R1631 B.n687 B.n98 10.6151
R1632 B.n691 B.n98 10.6151
R1633 B.n692 B.n691 10.6151
R1634 B.n693 B.n692 10.6151
R1635 B.n693 B.n96 10.6151
R1636 B.n697 B.n96 10.6151
R1637 B.n698 B.n697 10.6151
R1638 B.n699 B.n698 10.6151
R1639 B.n699 B.n94 10.6151
R1640 B.n703 B.n94 10.6151
R1641 B.n704 B.n703 10.6151
R1642 B.n705 B.n704 10.6151
R1643 B.n705 B.n92 10.6151
R1644 B.n709 B.n92 10.6151
R1645 B.n710 B.n709 10.6151
R1646 B.n711 B.n710 10.6151
R1647 B.n711 B.n90 10.6151
R1648 B.n715 B.n90 10.6151
R1649 B.n716 B.n715 10.6151
R1650 B.n717 B.n716 10.6151
R1651 B.n717 B.n88 10.6151
R1652 B.n721 B.n88 10.6151
R1653 B.n722 B.n721 10.6151
R1654 B.n363 B.n210 10.6151
R1655 B.n367 B.n210 10.6151
R1656 B.n368 B.n367 10.6151
R1657 B.n369 B.n368 10.6151
R1658 B.n369 B.n208 10.6151
R1659 B.n373 B.n208 10.6151
R1660 B.n374 B.n373 10.6151
R1661 B.n375 B.n374 10.6151
R1662 B.n375 B.n206 10.6151
R1663 B.n379 B.n206 10.6151
R1664 B.n380 B.n379 10.6151
R1665 B.n381 B.n380 10.6151
R1666 B.n381 B.n204 10.6151
R1667 B.n385 B.n204 10.6151
R1668 B.n386 B.n385 10.6151
R1669 B.n387 B.n386 10.6151
R1670 B.n387 B.n202 10.6151
R1671 B.n391 B.n202 10.6151
R1672 B.n392 B.n391 10.6151
R1673 B.n393 B.n392 10.6151
R1674 B.n393 B.n200 10.6151
R1675 B.n397 B.n200 10.6151
R1676 B.n398 B.n397 10.6151
R1677 B.n399 B.n398 10.6151
R1678 B.n399 B.n198 10.6151
R1679 B.n403 B.n198 10.6151
R1680 B.n404 B.n403 10.6151
R1681 B.n405 B.n404 10.6151
R1682 B.n405 B.n196 10.6151
R1683 B.n409 B.n196 10.6151
R1684 B.n410 B.n409 10.6151
R1685 B.n411 B.n410 10.6151
R1686 B.n411 B.n194 10.6151
R1687 B.n415 B.n194 10.6151
R1688 B.n416 B.n415 10.6151
R1689 B.n417 B.n416 10.6151
R1690 B.n421 B.n420 10.6151
R1691 B.n422 B.n421 10.6151
R1692 B.n422 B.n188 10.6151
R1693 B.n426 B.n188 10.6151
R1694 B.n427 B.n426 10.6151
R1695 B.n428 B.n427 10.6151
R1696 B.n428 B.n186 10.6151
R1697 B.n432 B.n186 10.6151
R1698 B.n433 B.n432 10.6151
R1699 B.n435 B.n182 10.6151
R1700 B.n439 B.n182 10.6151
R1701 B.n440 B.n439 10.6151
R1702 B.n441 B.n440 10.6151
R1703 B.n441 B.n180 10.6151
R1704 B.n445 B.n180 10.6151
R1705 B.n446 B.n445 10.6151
R1706 B.n447 B.n446 10.6151
R1707 B.n447 B.n178 10.6151
R1708 B.n451 B.n178 10.6151
R1709 B.n452 B.n451 10.6151
R1710 B.n453 B.n452 10.6151
R1711 B.n453 B.n176 10.6151
R1712 B.n457 B.n176 10.6151
R1713 B.n458 B.n457 10.6151
R1714 B.n459 B.n458 10.6151
R1715 B.n459 B.n174 10.6151
R1716 B.n463 B.n174 10.6151
R1717 B.n464 B.n463 10.6151
R1718 B.n465 B.n464 10.6151
R1719 B.n465 B.n172 10.6151
R1720 B.n469 B.n172 10.6151
R1721 B.n470 B.n469 10.6151
R1722 B.n471 B.n470 10.6151
R1723 B.n471 B.n170 10.6151
R1724 B.n475 B.n170 10.6151
R1725 B.n476 B.n475 10.6151
R1726 B.n477 B.n476 10.6151
R1727 B.n477 B.n168 10.6151
R1728 B.n481 B.n168 10.6151
R1729 B.n482 B.n481 10.6151
R1730 B.n483 B.n482 10.6151
R1731 B.n483 B.n166 10.6151
R1732 B.n487 B.n166 10.6151
R1733 B.n488 B.n487 10.6151
R1734 B.n489 B.n488 10.6151
R1735 B.n362 B.n361 10.6151
R1736 B.n361 B.n212 10.6151
R1737 B.n357 B.n212 10.6151
R1738 B.n357 B.n356 10.6151
R1739 B.n356 B.n355 10.6151
R1740 B.n355 B.n214 10.6151
R1741 B.n351 B.n214 10.6151
R1742 B.n351 B.n350 10.6151
R1743 B.n350 B.n349 10.6151
R1744 B.n349 B.n216 10.6151
R1745 B.n345 B.n216 10.6151
R1746 B.n345 B.n344 10.6151
R1747 B.n344 B.n343 10.6151
R1748 B.n343 B.n218 10.6151
R1749 B.n339 B.n218 10.6151
R1750 B.n339 B.n338 10.6151
R1751 B.n338 B.n337 10.6151
R1752 B.n337 B.n220 10.6151
R1753 B.n333 B.n220 10.6151
R1754 B.n333 B.n332 10.6151
R1755 B.n332 B.n331 10.6151
R1756 B.n331 B.n222 10.6151
R1757 B.n327 B.n222 10.6151
R1758 B.n327 B.n326 10.6151
R1759 B.n326 B.n325 10.6151
R1760 B.n325 B.n224 10.6151
R1761 B.n321 B.n224 10.6151
R1762 B.n321 B.n320 10.6151
R1763 B.n320 B.n319 10.6151
R1764 B.n319 B.n226 10.6151
R1765 B.n315 B.n226 10.6151
R1766 B.n315 B.n314 10.6151
R1767 B.n314 B.n313 10.6151
R1768 B.n313 B.n228 10.6151
R1769 B.n309 B.n228 10.6151
R1770 B.n309 B.n308 10.6151
R1771 B.n308 B.n307 10.6151
R1772 B.n307 B.n230 10.6151
R1773 B.n303 B.n230 10.6151
R1774 B.n303 B.n302 10.6151
R1775 B.n302 B.n301 10.6151
R1776 B.n301 B.n232 10.6151
R1777 B.n297 B.n232 10.6151
R1778 B.n297 B.n296 10.6151
R1779 B.n296 B.n295 10.6151
R1780 B.n295 B.n234 10.6151
R1781 B.n291 B.n234 10.6151
R1782 B.n291 B.n290 10.6151
R1783 B.n290 B.n289 10.6151
R1784 B.n289 B.n236 10.6151
R1785 B.n285 B.n236 10.6151
R1786 B.n285 B.n284 10.6151
R1787 B.n284 B.n283 10.6151
R1788 B.n283 B.n238 10.6151
R1789 B.n279 B.n238 10.6151
R1790 B.n279 B.n278 10.6151
R1791 B.n278 B.n277 10.6151
R1792 B.n277 B.n240 10.6151
R1793 B.n273 B.n240 10.6151
R1794 B.n273 B.n272 10.6151
R1795 B.n272 B.n271 10.6151
R1796 B.n271 B.n242 10.6151
R1797 B.n267 B.n242 10.6151
R1798 B.n267 B.n266 10.6151
R1799 B.n266 B.n265 10.6151
R1800 B.n265 B.n244 10.6151
R1801 B.n261 B.n244 10.6151
R1802 B.n261 B.n260 10.6151
R1803 B.n260 B.n259 10.6151
R1804 B.n259 B.n246 10.6151
R1805 B.n255 B.n246 10.6151
R1806 B.n255 B.n254 10.6151
R1807 B.n254 B.n253 10.6151
R1808 B.n253 B.n248 10.6151
R1809 B.n249 B.n248 10.6151
R1810 B.n249 B.n0 10.6151
R1811 B.n963 B.n1 10.6151
R1812 B.n963 B.n962 10.6151
R1813 B.n962 B.n961 10.6151
R1814 B.n961 B.n4 10.6151
R1815 B.n957 B.n4 10.6151
R1816 B.n957 B.n956 10.6151
R1817 B.n956 B.n955 10.6151
R1818 B.n955 B.n6 10.6151
R1819 B.n951 B.n6 10.6151
R1820 B.n951 B.n950 10.6151
R1821 B.n950 B.n949 10.6151
R1822 B.n949 B.n8 10.6151
R1823 B.n945 B.n8 10.6151
R1824 B.n945 B.n944 10.6151
R1825 B.n944 B.n943 10.6151
R1826 B.n943 B.n10 10.6151
R1827 B.n939 B.n10 10.6151
R1828 B.n939 B.n938 10.6151
R1829 B.n938 B.n937 10.6151
R1830 B.n937 B.n12 10.6151
R1831 B.n933 B.n12 10.6151
R1832 B.n933 B.n932 10.6151
R1833 B.n932 B.n931 10.6151
R1834 B.n931 B.n14 10.6151
R1835 B.n927 B.n14 10.6151
R1836 B.n927 B.n926 10.6151
R1837 B.n926 B.n925 10.6151
R1838 B.n925 B.n16 10.6151
R1839 B.n921 B.n16 10.6151
R1840 B.n921 B.n920 10.6151
R1841 B.n920 B.n919 10.6151
R1842 B.n919 B.n18 10.6151
R1843 B.n915 B.n18 10.6151
R1844 B.n915 B.n914 10.6151
R1845 B.n914 B.n913 10.6151
R1846 B.n913 B.n20 10.6151
R1847 B.n909 B.n20 10.6151
R1848 B.n909 B.n908 10.6151
R1849 B.n908 B.n907 10.6151
R1850 B.n907 B.n22 10.6151
R1851 B.n903 B.n22 10.6151
R1852 B.n903 B.n902 10.6151
R1853 B.n902 B.n901 10.6151
R1854 B.n901 B.n24 10.6151
R1855 B.n897 B.n24 10.6151
R1856 B.n897 B.n896 10.6151
R1857 B.n896 B.n895 10.6151
R1858 B.n895 B.n26 10.6151
R1859 B.n891 B.n26 10.6151
R1860 B.n891 B.n890 10.6151
R1861 B.n890 B.n889 10.6151
R1862 B.n889 B.n28 10.6151
R1863 B.n885 B.n28 10.6151
R1864 B.n885 B.n884 10.6151
R1865 B.n884 B.n883 10.6151
R1866 B.n883 B.n30 10.6151
R1867 B.n879 B.n30 10.6151
R1868 B.n879 B.n878 10.6151
R1869 B.n878 B.n877 10.6151
R1870 B.n877 B.n32 10.6151
R1871 B.n873 B.n32 10.6151
R1872 B.n873 B.n872 10.6151
R1873 B.n872 B.n871 10.6151
R1874 B.n871 B.n34 10.6151
R1875 B.n867 B.n34 10.6151
R1876 B.n867 B.n866 10.6151
R1877 B.n866 B.n865 10.6151
R1878 B.n865 B.n36 10.6151
R1879 B.n861 B.n36 10.6151
R1880 B.n861 B.n860 10.6151
R1881 B.n860 B.n859 10.6151
R1882 B.n859 B.n38 10.6151
R1883 B.n855 B.n38 10.6151
R1884 B.n855 B.n854 10.6151
R1885 B.n854 B.n853 10.6151
R1886 B.n853 B.n40 10.6151
R1887 B.n795 B.n794 9.36635
R1888 B.n777 B.n68 9.36635
R1889 B.n417 B.n192 9.36635
R1890 B.n435 B.n434 9.36635
R1891 B.n967 B.n0 2.81026
R1892 B.n967 B.n1 2.81026
R1893 B.n794 B.n793 1.24928
R1894 B.n780 B.n68 1.24928
R1895 B.n420 B.n192 1.24928
R1896 B.n434 B.n433 1.24928
C0 VDD2 VN 9.963731f
C1 w_n5650_n3076# B 11.768201f
C2 VDD1 VTAIL 10.268099f
C3 VTAIL VP 11.1053f
C4 VN VTAIL 11.091001f
C5 w_n5650_n3076# VDD2 3.25143f
C6 VDD1 VP 10.5116f
C7 VN VDD1 0.155963f
C8 VN VP 9.554481f
C9 VDD2 B 2.89564f
C10 w_n5650_n3076# VTAIL 3.15483f
C11 VTAIL B 3.7562f
C12 w_n5650_n3076# VDD1 3.05746f
C13 w_n5650_n3076# VP 13.0841f
C14 w_n5650_n3076# VN 12.3455f
C15 VDD2 VTAIL 10.3266f
C16 VDD1 B 2.73995f
C17 B VP 2.76491f
C18 VN B 1.51757f
C19 VDD2 VDD1 2.80656f
C20 VDD2 VP 0.707626f
C21 VDD2 VSUBS 2.50192f
C22 VDD1 VSUBS 2.328182f
C23 VTAIL VSUBS 1.488997f
C24 VN VSUBS 9.28988f
C25 VP VSUBS 5.419412f
C26 B VSUBS 6.445994f
C27 w_n5650_n3076# VSUBS 0.214451p
C28 B.n0 VSUBS 0.005939f
C29 B.n1 VSUBS 0.005939f
C30 B.n2 VSUBS 0.009391f
C31 B.n3 VSUBS 0.009391f
C32 B.n4 VSUBS 0.009391f
C33 B.n5 VSUBS 0.009391f
C34 B.n6 VSUBS 0.009391f
C35 B.n7 VSUBS 0.009391f
C36 B.n8 VSUBS 0.009391f
C37 B.n9 VSUBS 0.009391f
C38 B.n10 VSUBS 0.009391f
C39 B.n11 VSUBS 0.009391f
C40 B.n12 VSUBS 0.009391f
C41 B.n13 VSUBS 0.009391f
C42 B.n14 VSUBS 0.009391f
C43 B.n15 VSUBS 0.009391f
C44 B.n16 VSUBS 0.009391f
C45 B.n17 VSUBS 0.009391f
C46 B.n18 VSUBS 0.009391f
C47 B.n19 VSUBS 0.009391f
C48 B.n20 VSUBS 0.009391f
C49 B.n21 VSUBS 0.009391f
C50 B.n22 VSUBS 0.009391f
C51 B.n23 VSUBS 0.009391f
C52 B.n24 VSUBS 0.009391f
C53 B.n25 VSUBS 0.009391f
C54 B.n26 VSUBS 0.009391f
C55 B.n27 VSUBS 0.009391f
C56 B.n28 VSUBS 0.009391f
C57 B.n29 VSUBS 0.009391f
C58 B.n30 VSUBS 0.009391f
C59 B.n31 VSUBS 0.009391f
C60 B.n32 VSUBS 0.009391f
C61 B.n33 VSUBS 0.009391f
C62 B.n34 VSUBS 0.009391f
C63 B.n35 VSUBS 0.009391f
C64 B.n36 VSUBS 0.009391f
C65 B.n37 VSUBS 0.009391f
C66 B.n38 VSUBS 0.009391f
C67 B.n39 VSUBS 0.009391f
C68 B.n40 VSUBS 0.021735f
C69 B.n41 VSUBS 0.009391f
C70 B.n42 VSUBS 0.009391f
C71 B.n43 VSUBS 0.009391f
C72 B.n44 VSUBS 0.009391f
C73 B.n45 VSUBS 0.009391f
C74 B.n46 VSUBS 0.009391f
C75 B.n47 VSUBS 0.009391f
C76 B.n48 VSUBS 0.009391f
C77 B.n49 VSUBS 0.009391f
C78 B.n50 VSUBS 0.009391f
C79 B.n51 VSUBS 0.009391f
C80 B.n52 VSUBS 0.009391f
C81 B.n53 VSUBS 0.009391f
C82 B.n54 VSUBS 0.009391f
C83 B.n55 VSUBS 0.009391f
C84 B.n56 VSUBS 0.009391f
C85 B.n57 VSUBS 0.009391f
C86 B.n58 VSUBS 0.009391f
C87 B.n59 VSUBS 0.009391f
C88 B.t2 VSUBS 0.453958f
C89 B.t1 VSUBS 0.489121f
C90 B.t0 VSUBS 2.36195f
C91 B.n60 VSUBS 0.27675f
C92 B.n61 VSUBS 0.101595f
C93 B.n62 VSUBS 0.009391f
C94 B.n63 VSUBS 0.009391f
C95 B.n64 VSUBS 0.009391f
C96 B.n65 VSUBS 0.009391f
C97 B.t8 VSUBS 0.453951f
C98 B.t7 VSUBS 0.489115f
C99 B.t6 VSUBS 2.36195f
C100 B.n66 VSUBS 0.276756f
C101 B.n67 VSUBS 0.101601f
C102 B.n68 VSUBS 0.021759f
C103 B.n69 VSUBS 0.009391f
C104 B.n70 VSUBS 0.009391f
C105 B.n71 VSUBS 0.009391f
C106 B.n72 VSUBS 0.009391f
C107 B.n73 VSUBS 0.009391f
C108 B.n74 VSUBS 0.009391f
C109 B.n75 VSUBS 0.009391f
C110 B.n76 VSUBS 0.009391f
C111 B.n77 VSUBS 0.009391f
C112 B.n78 VSUBS 0.009391f
C113 B.n79 VSUBS 0.009391f
C114 B.n80 VSUBS 0.009391f
C115 B.n81 VSUBS 0.009391f
C116 B.n82 VSUBS 0.009391f
C117 B.n83 VSUBS 0.009391f
C118 B.n84 VSUBS 0.009391f
C119 B.n85 VSUBS 0.009391f
C120 B.n86 VSUBS 0.009391f
C121 B.n87 VSUBS 0.021735f
C122 B.n88 VSUBS 0.009391f
C123 B.n89 VSUBS 0.009391f
C124 B.n90 VSUBS 0.009391f
C125 B.n91 VSUBS 0.009391f
C126 B.n92 VSUBS 0.009391f
C127 B.n93 VSUBS 0.009391f
C128 B.n94 VSUBS 0.009391f
C129 B.n95 VSUBS 0.009391f
C130 B.n96 VSUBS 0.009391f
C131 B.n97 VSUBS 0.009391f
C132 B.n98 VSUBS 0.009391f
C133 B.n99 VSUBS 0.009391f
C134 B.n100 VSUBS 0.009391f
C135 B.n101 VSUBS 0.009391f
C136 B.n102 VSUBS 0.009391f
C137 B.n103 VSUBS 0.009391f
C138 B.n104 VSUBS 0.009391f
C139 B.n105 VSUBS 0.009391f
C140 B.n106 VSUBS 0.009391f
C141 B.n107 VSUBS 0.009391f
C142 B.n108 VSUBS 0.009391f
C143 B.n109 VSUBS 0.009391f
C144 B.n110 VSUBS 0.009391f
C145 B.n111 VSUBS 0.009391f
C146 B.n112 VSUBS 0.009391f
C147 B.n113 VSUBS 0.009391f
C148 B.n114 VSUBS 0.009391f
C149 B.n115 VSUBS 0.009391f
C150 B.n116 VSUBS 0.009391f
C151 B.n117 VSUBS 0.009391f
C152 B.n118 VSUBS 0.009391f
C153 B.n119 VSUBS 0.009391f
C154 B.n120 VSUBS 0.009391f
C155 B.n121 VSUBS 0.009391f
C156 B.n122 VSUBS 0.009391f
C157 B.n123 VSUBS 0.009391f
C158 B.n124 VSUBS 0.009391f
C159 B.n125 VSUBS 0.009391f
C160 B.n126 VSUBS 0.009391f
C161 B.n127 VSUBS 0.009391f
C162 B.n128 VSUBS 0.009391f
C163 B.n129 VSUBS 0.009391f
C164 B.n130 VSUBS 0.009391f
C165 B.n131 VSUBS 0.009391f
C166 B.n132 VSUBS 0.009391f
C167 B.n133 VSUBS 0.009391f
C168 B.n134 VSUBS 0.009391f
C169 B.n135 VSUBS 0.009391f
C170 B.n136 VSUBS 0.009391f
C171 B.n137 VSUBS 0.009391f
C172 B.n138 VSUBS 0.009391f
C173 B.n139 VSUBS 0.009391f
C174 B.n140 VSUBS 0.009391f
C175 B.n141 VSUBS 0.009391f
C176 B.n142 VSUBS 0.009391f
C177 B.n143 VSUBS 0.009391f
C178 B.n144 VSUBS 0.009391f
C179 B.n145 VSUBS 0.009391f
C180 B.n146 VSUBS 0.009391f
C181 B.n147 VSUBS 0.009391f
C182 B.n148 VSUBS 0.009391f
C183 B.n149 VSUBS 0.009391f
C184 B.n150 VSUBS 0.009391f
C185 B.n151 VSUBS 0.009391f
C186 B.n152 VSUBS 0.009391f
C187 B.n153 VSUBS 0.009391f
C188 B.n154 VSUBS 0.009391f
C189 B.n155 VSUBS 0.009391f
C190 B.n156 VSUBS 0.009391f
C191 B.n157 VSUBS 0.009391f
C192 B.n158 VSUBS 0.009391f
C193 B.n159 VSUBS 0.009391f
C194 B.n160 VSUBS 0.009391f
C195 B.n161 VSUBS 0.009391f
C196 B.n162 VSUBS 0.009391f
C197 B.n163 VSUBS 0.009391f
C198 B.n164 VSUBS 0.021735f
C199 B.n165 VSUBS 0.009391f
C200 B.n166 VSUBS 0.009391f
C201 B.n167 VSUBS 0.009391f
C202 B.n168 VSUBS 0.009391f
C203 B.n169 VSUBS 0.009391f
C204 B.n170 VSUBS 0.009391f
C205 B.n171 VSUBS 0.009391f
C206 B.n172 VSUBS 0.009391f
C207 B.n173 VSUBS 0.009391f
C208 B.n174 VSUBS 0.009391f
C209 B.n175 VSUBS 0.009391f
C210 B.n176 VSUBS 0.009391f
C211 B.n177 VSUBS 0.009391f
C212 B.n178 VSUBS 0.009391f
C213 B.n179 VSUBS 0.009391f
C214 B.n180 VSUBS 0.009391f
C215 B.n181 VSUBS 0.009391f
C216 B.n182 VSUBS 0.009391f
C217 B.n183 VSUBS 0.009391f
C218 B.t10 VSUBS 0.453951f
C219 B.t11 VSUBS 0.489115f
C220 B.t9 VSUBS 2.36195f
C221 B.n184 VSUBS 0.276756f
C222 B.n185 VSUBS 0.101601f
C223 B.n186 VSUBS 0.009391f
C224 B.n187 VSUBS 0.009391f
C225 B.n188 VSUBS 0.009391f
C226 B.n189 VSUBS 0.009391f
C227 B.t4 VSUBS 0.453958f
C228 B.t5 VSUBS 0.489121f
C229 B.t3 VSUBS 2.36195f
C230 B.n190 VSUBS 0.27675f
C231 B.n191 VSUBS 0.101595f
C232 B.n192 VSUBS 0.021759f
C233 B.n193 VSUBS 0.009391f
C234 B.n194 VSUBS 0.009391f
C235 B.n195 VSUBS 0.009391f
C236 B.n196 VSUBS 0.009391f
C237 B.n197 VSUBS 0.009391f
C238 B.n198 VSUBS 0.009391f
C239 B.n199 VSUBS 0.009391f
C240 B.n200 VSUBS 0.009391f
C241 B.n201 VSUBS 0.009391f
C242 B.n202 VSUBS 0.009391f
C243 B.n203 VSUBS 0.009391f
C244 B.n204 VSUBS 0.009391f
C245 B.n205 VSUBS 0.009391f
C246 B.n206 VSUBS 0.009391f
C247 B.n207 VSUBS 0.009391f
C248 B.n208 VSUBS 0.009391f
C249 B.n209 VSUBS 0.009391f
C250 B.n210 VSUBS 0.009391f
C251 B.n211 VSUBS 0.021735f
C252 B.n212 VSUBS 0.009391f
C253 B.n213 VSUBS 0.009391f
C254 B.n214 VSUBS 0.009391f
C255 B.n215 VSUBS 0.009391f
C256 B.n216 VSUBS 0.009391f
C257 B.n217 VSUBS 0.009391f
C258 B.n218 VSUBS 0.009391f
C259 B.n219 VSUBS 0.009391f
C260 B.n220 VSUBS 0.009391f
C261 B.n221 VSUBS 0.009391f
C262 B.n222 VSUBS 0.009391f
C263 B.n223 VSUBS 0.009391f
C264 B.n224 VSUBS 0.009391f
C265 B.n225 VSUBS 0.009391f
C266 B.n226 VSUBS 0.009391f
C267 B.n227 VSUBS 0.009391f
C268 B.n228 VSUBS 0.009391f
C269 B.n229 VSUBS 0.009391f
C270 B.n230 VSUBS 0.009391f
C271 B.n231 VSUBS 0.009391f
C272 B.n232 VSUBS 0.009391f
C273 B.n233 VSUBS 0.009391f
C274 B.n234 VSUBS 0.009391f
C275 B.n235 VSUBS 0.009391f
C276 B.n236 VSUBS 0.009391f
C277 B.n237 VSUBS 0.009391f
C278 B.n238 VSUBS 0.009391f
C279 B.n239 VSUBS 0.009391f
C280 B.n240 VSUBS 0.009391f
C281 B.n241 VSUBS 0.009391f
C282 B.n242 VSUBS 0.009391f
C283 B.n243 VSUBS 0.009391f
C284 B.n244 VSUBS 0.009391f
C285 B.n245 VSUBS 0.009391f
C286 B.n246 VSUBS 0.009391f
C287 B.n247 VSUBS 0.009391f
C288 B.n248 VSUBS 0.009391f
C289 B.n249 VSUBS 0.009391f
C290 B.n250 VSUBS 0.009391f
C291 B.n251 VSUBS 0.009391f
C292 B.n252 VSUBS 0.009391f
C293 B.n253 VSUBS 0.009391f
C294 B.n254 VSUBS 0.009391f
C295 B.n255 VSUBS 0.009391f
C296 B.n256 VSUBS 0.009391f
C297 B.n257 VSUBS 0.009391f
C298 B.n258 VSUBS 0.009391f
C299 B.n259 VSUBS 0.009391f
C300 B.n260 VSUBS 0.009391f
C301 B.n261 VSUBS 0.009391f
C302 B.n262 VSUBS 0.009391f
C303 B.n263 VSUBS 0.009391f
C304 B.n264 VSUBS 0.009391f
C305 B.n265 VSUBS 0.009391f
C306 B.n266 VSUBS 0.009391f
C307 B.n267 VSUBS 0.009391f
C308 B.n268 VSUBS 0.009391f
C309 B.n269 VSUBS 0.009391f
C310 B.n270 VSUBS 0.009391f
C311 B.n271 VSUBS 0.009391f
C312 B.n272 VSUBS 0.009391f
C313 B.n273 VSUBS 0.009391f
C314 B.n274 VSUBS 0.009391f
C315 B.n275 VSUBS 0.009391f
C316 B.n276 VSUBS 0.009391f
C317 B.n277 VSUBS 0.009391f
C318 B.n278 VSUBS 0.009391f
C319 B.n279 VSUBS 0.009391f
C320 B.n280 VSUBS 0.009391f
C321 B.n281 VSUBS 0.009391f
C322 B.n282 VSUBS 0.009391f
C323 B.n283 VSUBS 0.009391f
C324 B.n284 VSUBS 0.009391f
C325 B.n285 VSUBS 0.009391f
C326 B.n286 VSUBS 0.009391f
C327 B.n287 VSUBS 0.009391f
C328 B.n288 VSUBS 0.009391f
C329 B.n289 VSUBS 0.009391f
C330 B.n290 VSUBS 0.009391f
C331 B.n291 VSUBS 0.009391f
C332 B.n292 VSUBS 0.009391f
C333 B.n293 VSUBS 0.009391f
C334 B.n294 VSUBS 0.009391f
C335 B.n295 VSUBS 0.009391f
C336 B.n296 VSUBS 0.009391f
C337 B.n297 VSUBS 0.009391f
C338 B.n298 VSUBS 0.009391f
C339 B.n299 VSUBS 0.009391f
C340 B.n300 VSUBS 0.009391f
C341 B.n301 VSUBS 0.009391f
C342 B.n302 VSUBS 0.009391f
C343 B.n303 VSUBS 0.009391f
C344 B.n304 VSUBS 0.009391f
C345 B.n305 VSUBS 0.009391f
C346 B.n306 VSUBS 0.009391f
C347 B.n307 VSUBS 0.009391f
C348 B.n308 VSUBS 0.009391f
C349 B.n309 VSUBS 0.009391f
C350 B.n310 VSUBS 0.009391f
C351 B.n311 VSUBS 0.009391f
C352 B.n312 VSUBS 0.009391f
C353 B.n313 VSUBS 0.009391f
C354 B.n314 VSUBS 0.009391f
C355 B.n315 VSUBS 0.009391f
C356 B.n316 VSUBS 0.009391f
C357 B.n317 VSUBS 0.009391f
C358 B.n318 VSUBS 0.009391f
C359 B.n319 VSUBS 0.009391f
C360 B.n320 VSUBS 0.009391f
C361 B.n321 VSUBS 0.009391f
C362 B.n322 VSUBS 0.009391f
C363 B.n323 VSUBS 0.009391f
C364 B.n324 VSUBS 0.009391f
C365 B.n325 VSUBS 0.009391f
C366 B.n326 VSUBS 0.009391f
C367 B.n327 VSUBS 0.009391f
C368 B.n328 VSUBS 0.009391f
C369 B.n329 VSUBS 0.009391f
C370 B.n330 VSUBS 0.009391f
C371 B.n331 VSUBS 0.009391f
C372 B.n332 VSUBS 0.009391f
C373 B.n333 VSUBS 0.009391f
C374 B.n334 VSUBS 0.009391f
C375 B.n335 VSUBS 0.009391f
C376 B.n336 VSUBS 0.009391f
C377 B.n337 VSUBS 0.009391f
C378 B.n338 VSUBS 0.009391f
C379 B.n339 VSUBS 0.009391f
C380 B.n340 VSUBS 0.009391f
C381 B.n341 VSUBS 0.009391f
C382 B.n342 VSUBS 0.009391f
C383 B.n343 VSUBS 0.009391f
C384 B.n344 VSUBS 0.009391f
C385 B.n345 VSUBS 0.009391f
C386 B.n346 VSUBS 0.009391f
C387 B.n347 VSUBS 0.009391f
C388 B.n348 VSUBS 0.009391f
C389 B.n349 VSUBS 0.009391f
C390 B.n350 VSUBS 0.009391f
C391 B.n351 VSUBS 0.009391f
C392 B.n352 VSUBS 0.009391f
C393 B.n353 VSUBS 0.009391f
C394 B.n354 VSUBS 0.009391f
C395 B.n355 VSUBS 0.009391f
C396 B.n356 VSUBS 0.009391f
C397 B.n357 VSUBS 0.009391f
C398 B.n358 VSUBS 0.009391f
C399 B.n359 VSUBS 0.009391f
C400 B.n360 VSUBS 0.009391f
C401 B.n361 VSUBS 0.009391f
C402 B.n362 VSUBS 0.021735f
C403 B.n363 VSUBS 0.022459f
C404 B.n364 VSUBS 0.02246f
C405 B.n365 VSUBS 0.009391f
C406 B.n366 VSUBS 0.009391f
C407 B.n367 VSUBS 0.009391f
C408 B.n368 VSUBS 0.009391f
C409 B.n369 VSUBS 0.009391f
C410 B.n370 VSUBS 0.009391f
C411 B.n371 VSUBS 0.009391f
C412 B.n372 VSUBS 0.009391f
C413 B.n373 VSUBS 0.009391f
C414 B.n374 VSUBS 0.009391f
C415 B.n375 VSUBS 0.009391f
C416 B.n376 VSUBS 0.009391f
C417 B.n377 VSUBS 0.009391f
C418 B.n378 VSUBS 0.009391f
C419 B.n379 VSUBS 0.009391f
C420 B.n380 VSUBS 0.009391f
C421 B.n381 VSUBS 0.009391f
C422 B.n382 VSUBS 0.009391f
C423 B.n383 VSUBS 0.009391f
C424 B.n384 VSUBS 0.009391f
C425 B.n385 VSUBS 0.009391f
C426 B.n386 VSUBS 0.009391f
C427 B.n387 VSUBS 0.009391f
C428 B.n388 VSUBS 0.009391f
C429 B.n389 VSUBS 0.009391f
C430 B.n390 VSUBS 0.009391f
C431 B.n391 VSUBS 0.009391f
C432 B.n392 VSUBS 0.009391f
C433 B.n393 VSUBS 0.009391f
C434 B.n394 VSUBS 0.009391f
C435 B.n395 VSUBS 0.009391f
C436 B.n396 VSUBS 0.009391f
C437 B.n397 VSUBS 0.009391f
C438 B.n398 VSUBS 0.009391f
C439 B.n399 VSUBS 0.009391f
C440 B.n400 VSUBS 0.009391f
C441 B.n401 VSUBS 0.009391f
C442 B.n402 VSUBS 0.009391f
C443 B.n403 VSUBS 0.009391f
C444 B.n404 VSUBS 0.009391f
C445 B.n405 VSUBS 0.009391f
C446 B.n406 VSUBS 0.009391f
C447 B.n407 VSUBS 0.009391f
C448 B.n408 VSUBS 0.009391f
C449 B.n409 VSUBS 0.009391f
C450 B.n410 VSUBS 0.009391f
C451 B.n411 VSUBS 0.009391f
C452 B.n412 VSUBS 0.009391f
C453 B.n413 VSUBS 0.009391f
C454 B.n414 VSUBS 0.009391f
C455 B.n415 VSUBS 0.009391f
C456 B.n416 VSUBS 0.009391f
C457 B.n417 VSUBS 0.008839f
C458 B.n418 VSUBS 0.009391f
C459 B.n419 VSUBS 0.009391f
C460 B.n420 VSUBS 0.005248f
C461 B.n421 VSUBS 0.009391f
C462 B.n422 VSUBS 0.009391f
C463 B.n423 VSUBS 0.009391f
C464 B.n424 VSUBS 0.009391f
C465 B.n425 VSUBS 0.009391f
C466 B.n426 VSUBS 0.009391f
C467 B.n427 VSUBS 0.009391f
C468 B.n428 VSUBS 0.009391f
C469 B.n429 VSUBS 0.009391f
C470 B.n430 VSUBS 0.009391f
C471 B.n431 VSUBS 0.009391f
C472 B.n432 VSUBS 0.009391f
C473 B.n433 VSUBS 0.005248f
C474 B.n434 VSUBS 0.021759f
C475 B.n435 VSUBS 0.008839f
C476 B.n436 VSUBS 0.009391f
C477 B.n437 VSUBS 0.009391f
C478 B.n438 VSUBS 0.009391f
C479 B.n439 VSUBS 0.009391f
C480 B.n440 VSUBS 0.009391f
C481 B.n441 VSUBS 0.009391f
C482 B.n442 VSUBS 0.009391f
C483 B.n443 VSUBS 0.009391f
C484 B.n444 VSUBS 0.009391f
C485 B.n445 VSUBS 0.009391f
C486 B.n446 VSUBS 0.009391f
C487 B.n447 VSUBS 0.009391f
C488 B.n448 VSUBS 0.009391f
C489 B.n449 VSUBS 0.009391f
C490 B.n450 VSUBS 0.009391f
C491 B.n451 VSUBS 0.009391f
C492 B.n452 VSUBS 0.009391f
C493 B.n453 VSUBS 0.009391f
C494 B.n454 VSUBS 0.009391f
C495 B.n455 VSUBS 0.009391f
C496 B.n456 VSUBS 0.009391f
C497 B.n457 VSUBS 0.009391f
C498 B.n458 VSUBS 0.009391f
C499 B.n459 VSUBS 0.009391f
C500 B.n460 VSUBS 0.009391f
C501 B.n461 VSUBS 0.009391f
C502 B.n462 VSUBS 0.009391f
C503 B.n463 VSUBS 0.009391f
C504 B.n464 VSUBS 0.009391f
C505 B.n465 VSUBS 0.009391f
C506 B.n466 VSUBS 0.009391f
C507 B.n467 VSUBS 0.009391f
C508 B.n468 VSUBS 0.009391f
C509 B.n469 VSUBS 0.009391f
C510 B.n470 VSUBS 0.009391f
C511 B.n471 VSUBS 0.009391f
C512 B.n472 VSUBS 0.009391f
C513 B.n473 VSUBS 0.009391f
C514 B.n474 VSUBS 0.009391f
C515 B.n475 VSUBS 0.009391f
C516 B.n476 VSUBS 0.009391f
C517 B.n477 VSUBS 0.009391f
C518 B.n478 VSUBS 0.009391f
C519 B.n479 VSUBS 0.009391f
C520 B.n480 VSUBS 0.009391f
C521 B.n481 VSUBS 0.009391f
C522 B.n482 VSUBS 0.009391f
C523 B.n483 VSUBS 0.009391f
C524 B.n484 VSUBS 0.009391f
C525 B.n485 VSUBS 0.009391f
C526 B.n486 VSUBS 0.009391f
C527 B.n487 VSUBS 0.009391f
C528 B.n488 VSUBS 0.009391f
C529 B.n489 VSUBS 0.022459f
C530 B.n490 VSUBS 0.02246f
C531 B.n491 VSUBS 0.021735f
C532 B.n492 VSUBS 0.009391f
C533 B.n493 VSUBS 0.009391f
C534 B.n494 VSUBS 0.009391f
C535 B.n495 VSUBS 0.009391f
C536 B.n496 VSUBS 0.009391f
C537 B.n497 VSUBS 0.009391f
C538 B.n498 VSUBS 0.009391f
C539 B.n499 VSUBS 0.009391f
C540 B.n500 VSUBS 0.009391f
C541 B.n501 VSUBS 0.009391f
C542 B.n502 VSUBS 0.009391f
C543 B.n503 VSUBS 0.009391f
C544 B.n504 VSUBS 0.009391f
C545 B.n505 VSUBS 0.009391f
C546 B.n506 VSUBS 0.009391f
C547 B.n507 VSUBS 0.009391f
C548 B.n508 VSUBS 0.009391f
C549 B.n509 VSUBS 0.009391f
C550 B.n510 VSUBS 0.009391f
C551 B.n511 VSUBS 0.009391f
C552 B.n512 VSUBS 0.009391f
C553 B.n513 VSUBS 0.009391f
C554 B.n514 VSUBS 0.009391f
C555 B.n515 VSUBS 0.009391f
C556 B.n516 VSUBS 0.009391f
C557 B.n517 VSUBS 0.009391f
C558 B.n518 VSUBS 0.009391f
C559 B.n519 VSUBS 0.009391f
C560 B.n520 VSUBS 0.009391f
C561 B.n521 VSUBS 0.009391f
C562 B.n522 VSUBS 0.009391f
C563 B.n523 VSUBS 0.009391f
C564 B.n524 VSUBS 0.009391f
C565 B.n525 VSUBS 0.009391f
C566 B.n526 VSUBS 0.009391f
C567 B.n527 VSUBS 0.009391f
C568 B.n528 VSUBS 0.009391f
C569 B.n529 VSUBS 0.009391f
C570 B.n530 VSUBS 0.009391f
C571 B.n531 VSUBS 0.009391f
C572 B.n532 VSUBS 0.009391f
C573 B.n533 VSUBS 0.009391f
C574 B.n534 VSUBS 0.009391f
C575 B.n535 VSUBS 0.009391f
C576 B.n536 VSUBS 0.009391f
C577 B.n537 VSUBS 0.009391f
C578 B.n538 VSUBS 0.009391f
C579 B.n539 VSUBS 0.009391f
C580 B.n540 VSUBS 0.009391f
C581 B.n541 VSUBS 0.009391f
C582 B.n542 VSUBS 0.009391f
C583 B.n543 VSUBS 0.009391f
C584 B.n544 VSUBS 0.009391f
C585 B.n545 VSUBS 0.009391f
C586 B.n546 VSUBS 0.009391f
C587 B.n547 VSUBS 0.009391f
C588 B.n548 VSUBS 0.009391f
C589 B.n549 VSUBS 0.009391f
C590 B.n550 VSUBS 0.009391f
C591 B.n551 VSUBS 0.009391f
C592 B.n552 VSUBS 0.009391f
C593 B.n553 VSUBS 0.009391f
C594 B.n554 VSUBS 0.009391f
C595 B.n555 VSUBS 0.009391f
C596 B.n556 VSUBS 0.009391f
C597 B.n557 VSUBS 0.009391f
C598 B.n558 VSUBS 0.009391f
C599 B.n559 VSUBS 0.009391f
C600 B.n560 VSUBS 0.009391f
C601 B.n561 VSUBS 0.009391f
C602 B.n562 VSUBS 0.009391f
C603 B.n563 VSUBS 0.009391f
C604 B.n564 VSUBS 0.009391f
C605 B.n565 VSUBS 0.009391f
C606 B.n566 VSUBS 0.009391f
C607 B.n567 VSUBS 0.009391f
C608 B.n568 VSUBS 0.009391f
C609 B.n569 VSUBS 0.009391f
C610 B.n570 VSUBS 0.009391f
C611 B.n571 VSUBS 0.009391f
C612 B.n572 VSUBS 0.009391f
C613 B.n573 VSUBS 0.009391f
C614 B.n574 VSUBS 0.009391f
C615 B.n575 VSUBS 0.009391f
C616 B.n576 VSUBS 0.009391f
C617 B.n577 VSUBS 0.009391f
C618 B.n578 VSUBS 0.009391f
C619 B.n579 VSUBS 0.009391f
C620 B.n580 VSUBS 0.009391f
C621 B.n581 VSUBS 0.009391f
C622 B.n582 VSUBS 0.009391f
C623 B.n583 VSUBS 0.009391f
C624 B.n584 VSUBS 0.009391f
C625 B.n585 VSUBS 0.009391f
C626 B.n586 VSUBS 0.009391f
C627 B.n587 VSUBS 0.009391f
C628 B.n588 VSUBS 0.009391f
C629 B.n589 VSUBS 0.009391f
C630 B.n590 VSUBS 0.009391f
C631 B.n591 VSUBS 0.009391f
C632 B.n592 VSUBS 0.009391f
C633 B.n593 VSUBS 0.009391f
C634 B.n594 VSUBS 0.009391f
C635 B.n595 VSUBS 0.009391f
C636 B.n596 VSUBS 0.009391f
C637 B.n597 VSUBS 0.009391f
C638 B.n598 VSUBS 0.009391f
C639 B.n599 VSUBS 0.009391f
C640 B.n600 VSUBS 0.009391f
C641 B.n601 VSUBS 0.009391f
C642 B.n602 VSUBS 0.009391f
C643 B.n603 VSUBS 0.009391f
C644 B.n604 VSUBS 0.009391f
C645 B.n605 VSUBS 0.009391f
C646 B.n606 VSUBS 0.009391f
C647 B.n607 VSUBS 0.009391f
C648 B.n608 VSUBS 0.009391f
C649 B.n609 VSUBS 0.009391f
C650 B.n610 VSUBS 0.009391f
C651 B.n611 VSUBS 0.009391f
C652 B.n612 VSUBS 0.009391f
C653 B.n613 VSUBS 0.009391f
C654 B.n614 VSUBS 0.009391f
C655 B.n615 VSUBS 0.009391f
C656 B.n616 VSUBS 0.009391f
C657 B.n617 VSUBS 0.009391f
C658 B.n618 VSUBS 0.009391f
C659 B.n619 VSUBS 0.009391f
C660 B.n620 VSUBS 0.009391f
C661 B.n621 VSUBS 0.009391f
C662 B.n622 VSUBS 0.009391f
C663 B.n623 VSUBS 0.009391f
C664 B.n624 VSUBS 0.009391f
C665 B.n625 VSUBS 0.009391f
C666 B.n626 VSUBS 0.009391f
C667 B.n627 VSUBS 0.009391f
C668 B.n628 VSUBS 0.009391f
C669 B.n629 VSUBS 0.009391f
C670 B.n630 VSUBS 0.009391f
C671 B.n631 VSUBS 0.009391f
C672 B.n632 VSUBS 0.009391f
C673 B.n633 VSUBS 0.009391f
C674 B.n634 VSUBS 0.009391f
C675 B.n635 VSUBS 0.009391f
C676 B.n636 VSUBS 0.009391f
C677 B.n637 VSUBS 0.009391f
C678 B.n638 VSUBS 0.009391f
C679 B.n639 VSUBS 0.009391f
C680 B.n640 VSUBS 0.009391f
C681 B.n641 VSUBS 0.009391f
C682 B.n642 VSUBS 0.009391f
C683 B.n643 VSUBS 0.009391f
C684 B.n644 VSUBS 0.009391f
C685 B.n645 VSUBS 0.009391f
C686 B.n646 VSUBS 0.009391f
C687 B.n647 VSUBS 0.009391f
C688 B.n648 VSUBS 0.009391f
C689 B.n649 VSUBS 0.009391f
C690 B.n650 VSUBS 0.009391f
C691 B.n651 VSUBS 0.009391f
C692 B.n652 VSUBS 0.009391f
C693 B.n653 VSUBS 0.009391f
C694 B.n654 VSUBS 0.009391f
C695 B.n655 VSUBS 0.009391f
C696 B.n656 VSUBS 0.009391f
C697 B.n657 VSUBS 0.009391f
C698 B.n658 VSUBS 0.009391f
C699 B.n659 VSUBS 0.009391f
C700 B.n660 VSUBS 0.009391f
C701 B.n661 VSUBS 0.009391f
C702 B.n662 VSUBS 0.009391f
C703 B.n663 VSUBS 0.009391f
C704 B.n664 VSUBS 0.009391f
C705 B.n665 VSUBS 0.009391f
C706 B.n666 VSUBS 0.009391f
C707 B.n667 VSUBS 0.009391f
C708 B.n668 VSUBS 0.009391f
C709 B.n669 VSUBS 0.009391f
C710 B.n670 VSUBS 0.009391f
C711 B.n671 VSUBS 0.009391f
C712 B.n672 VSUBS 0.009391f
C713 B.n673 VSUBS 0.009391f
C714 B.n674 VSUBS 0.009391f
C715 B.n675 VSUBS 0.009391f
C716 B.n676 VSUBS 0.009391f
C717 B.n677 VSUBS 0.009391f
C718 B.n678 VSUBS 0.009391f
C719 B.n679 VSUBS 0.009391f
C720 B.n680 VSUBS 0.009391f
C721 B.n681 VSUBS 0.009391f
C722 B.n682 VSUBS 0.009391f
C723 B.n683 VSUBS 0.009391f
C724 B.n684 VSUBS 0.009391f
C725 B.n685 VSUBS 0.009391f
C726 B.n686 VSUBS 0.009391f
C727 B.n687 VSUBS 0.009391f
C728 B.n688 VSUBS 0.009391f
C729 B.n689 VSUBS 0.009391f
C730 B.n690 VSUBS 0.009391f
C731 B.n691 VSUBS 0.009391f
C732 B.n692 VSUBS 0.009391f
C733 B.n693 VSUBS 0.009391f
C734 B.n694 VSUBS 0.009391f
C735 B.n695 VSUBS 0.009391f
C736 B.n696 VSUBS 0.009391f
C737 B.n697 VSUBS 0.009391f
C738 B.n698 VSUBS 0.009391f
C739 B.n699 VSUBS 0.009391f
C740 B.n700 VSUBS 0.009391f
C741 B.n701 VSUBS 0.009391f
C742 B.n702 VSUBS 0.009391f
C743 B.n703 VSUBS 0.009391f
C744 B.n704 VSUBS 0.009391f
C745 B.n705 VSUBS 0.009391f
C746 B.n706 VSUBS 0.009391f
C747 B.n707 VSUBS 0.009391f
C748 B.n708 VSUBS 0.009391f
C749 B.n709 VSUBS 0.009391f
C750 B.n710 VSUBS 0.009391f
C751 B.n711 VSUBS 0.009391f
C752 B.n712 VSUBS 0.009391f
C753 B.n713 VSUBS 0.009391f
C754 B.n714 VSUBS 0.009391f
C755 B.n715 VSUBS 0.009391f
C756 B.n716 VSUBS 0.009391f
C757 B.n717 VSUBS 0.009391f
C758 B.n718 VSUBS 0.009391f
C759 B.n719 VSUBS 0.009391f
C760 B.n720 VSUBS 0.009391f
C761 B.n721 VSUBS 0.009391f
C762 B.n722 VSUBS 0.022835f
C763 B.n723 VSUBS 0.021359f
C764 B.n724 VSUBS 0.02246f
C765 B.n725 VSUBS 0.009391f
C766 B.n726 VSUBS 0.009391f
C767 B.n727 VSUBS 0.009391f
C768 B.n728 VSUBS 0.009391f
C769 B.n729 VSUBS 0.009391f
C770 B.n730 VSUBS 0.009391f
C771 B.n731 VSUBS 0.009391f
C772 B.n732 VSUBS 0.009391f
C773 B.n733 VSUBS 0.009391f
C774 B.n734 VSUBS 0.009391f
C775 B.n735 VSUBS 0.009391f
C776 B.n736 VSUBS 0.009391f
C777 B.n737 VSUBS 0.009391f
C778 B.n738 VSUBS 0.009391f
C779 B.n739 VSUBS 0.009391f
C780 B.n740 VSUBS 0.009391f
C781 B.n741 VSUBS 0.009391f
C782 B.n742 VSUBS 0.009391f
C783 B.n743 VSUBS 0.009391f
C784 B.n744 VSUBS 0.009391f
C785 B.n745 VSUBS 0.009391f
C786 B.n746 VSUBS 0.009391f
C787 B.n747 VSUBS 0.009391f
C788 B.n748 VSUBS 0.009391f
C789 B.n749 VSUBS 0.009391f
C790 B.n750 VSUBS 0.009391f
C791 B.n751 VSUBS 0.009391f
C792 B.n752 VSUBS 0.009391f
C793 B.n753 VSUBS 0.009391f
C794 B.n754 VSUBS 0.009391f
C795 B.n755 VSUBS 0.009391f
C796 B.n756 VSUBS 0.009391f
C797 B.n757 VSUBS 0.009391f
C798 B.n758 VSUBS 0.009391f
C799 B.n759 VSUBS 0.009391f
C800 B.n760 VSUBS 0.009391f
C801 B.n761 VSUBS 0.009391f
C802 B.n762 VSUBS 0.009391f
C803 B.n763 VSUBS 0.009391f
C804 B.n764 VSUBS 0.009391f
C805 B.n765 VSUBS 0.009391f
C806 B.n766 VSUBS 0.009391f
C807 B.n767 VSUBS 0.009391f
C808 B.n768 VSUBS 0.009391f
C809 B.n769 VSUBS 0.009391f
C810 B.n770 VSUBS 0.009391f
C811 B.n771 VSUBS 0.009391f
C812 B.n772 VSUBS 0.009391f
C813 B.n773 VSUBS 0.009391f
C814 B.n774 VSUBS 0.009391f
C815 B.n775 VSUBS 0.009391f
C816 B.n776 VSUBS 0.009391f
C817 B.n777 VSUBS 0.008839f
C818 B.n778 VSUBS 0.009391f
C819 B.n779 VSUBS 0.009391f
C820 B.n780 VSUBS 0.005248f
C821 B.n781 VSUBS 0.009391f
C822 B.n782 VSUBS 0.009391f
C823 B.n783 VSUBS 0.009391f
C824 B.n784 VSUBS 0.009391f
C825 B.n785 VSUBS 0.009391f
C826 B.n786 VSUBS 0.009391f
C827 B.n787 VSUBS 0.009391f
C828 B.n788 VSUBS 0.009391f
C829 B.n789 VSUBS 0.009391f
C830 B.n790 VSUBS 0.009391f
C831 B.n791 VSUBS 0.009391f
C832 B.n792 VSUBS 0.009391f
C833 B.n793 VSUBS 0.005248f
C834 B.n794 VSUBS 0.021759f
C835 B.n795 VSUBS 0.008839f
C836 B.n796 VSUBS 0.009391f
C837 B.n797 VSUBS 0.009391f
C838 B.n798 VSUBS 0.009391f
C839 B.n799 VSUBS 0.009391f
C840 B.n800 VSUBS 0.009391f
C841 B.n801 VSUBS 0.009391f
C842 B.n802 VSUBS 0.009391f
C843 B.n803 VSUBS 0.009391f
C844 B.n804 VSUBS 0.009391f
C845 B.n805 VSUBS 0.009391f
C846 B.n806 VSUBS 0.009391f
C847 B.n807 VSUBS 0.009391f
C848 B.n808 VSUBS 0.009391f
C849 B.n809 VSUBS 0.009391f
C850 B.n810 VSUBS 0.009391f
C851 B.n811 VSUBS 0.009391f
C852 B.n812 VSUBS 0.009391f
C853 B.n813 VSUBS 0.009391f
C854 B.n814 VSUBS 0.009391f
C855 B.n815 VSUBS 0.009391f
C856 B.n816 VSUBS 0.009391f
C857 B.n817 VSUBS 0.009391f
C858 B.n818 VSUBS 0.009391f
C859 B.n819 VSUBS 0.009391f
C860 B.n820 VSUBS 0.009391f
C861 B.n821 VSUBS 0.009391f
C862 B.n822 VSUBS 0.009391f
C863 B.n823 VSUBS 0.009391f
C864 B.n824 VSUBS 0.009391f
C865 B.n825 VSUBS 0.009391f
C866 B.n826 VSUBS 0.009391f
C867 B.n827 VSUBS 0.009391f
C868 B.n828 VSUBS 0.009391f
C869 B.n829 VSUBS 0.009391f
C870 B.n830 VSUBS 0.009391f
C871 B.n831 VSUBS 0.009391f
C872 B.n832 VSUBS 0.009391f
C873 B.n833 VSUBS 0.009391f
C874 B.n834 VSUBS 0.009391f
C875 B.n835 VSUBS 0.009391f
C876 B.n836 VSUBS 0.009391f
C877 B.n837 VSUBS 0.009391f
C878 B.n838 VSUBS 0.009391f
C879 B.n839 VSUBS 0.009391f
C880 B.n840 VSUBS 0.009391f
C881 B.n841 VSUBS 0.009391f
C882 B.n842 VSUBS 0.009391f
C883 B.n843 VSUBS 0.009391f
C884 B.n844 VSUBS 0.009391f
C885 B.n845 VSUBS 0.009391f
C886 B.n846 VSUBS 0.009391f
C887 B.n847 VSUBS 0.009391f
C888 B.n848 VSUBS 0.009391f
C889 B.n849 VSUBS 0.022459f
C890 B.n850 VSUBS 0.02246f
C891 B.n851 VSUBS 0.021735f
C892 B.n852 VSUBS 0.009391f
C893 B.n853 VSUBS 0.009391f
C894 B.n854 VSUBS 0.009391f
C895 B.n855 VSUBS 0.009391f
C896 B.n856 VSUBS 0.009391f
C897 B.n857 VSUBS 0.009391f
C898 B.n858 VSUBS 0.009391f
C899 B.n859 VSUBS 0.009391f
C900 B.n860 VSUBS 0.009391f
C901 B.n861 VSUBS 0.009391f
C902 B.n862 VSUBS 0.009391f
C903 B.n863 VSUBS 0.009391f
C904 B.n864 VSUBS 0.009391f
C905 B.n865 VSUBS 0.009391f
C906 B.n866 VSUBS 0.009391f
C907 B.n867 VSUBS 0.009391f
C908 B.n868 VSUBS 0.009391f
C909 B.n869 VSUBS 0.009391f
C910 B.n870 VSUBS 0.009391f
C911 B.n871 VSUBS 0.009391f
C912 B.n872 VSUBS 0.009391f
C913 B.n873 VSUBS 0.009391f
C914 B.n874 VSUBS 0.009391f
C915 B.n875 VSUBS 0.009391f
C916 B.n876 VSUBS 0.009391f
C917 B.n877 VSUBS 0.009391f
C918 B.n878 VSUBS 0.009391f
C919 B.n879 VSUBS 0.009391f
C920 B.n880 VSUBS 0.009391f
C921 B.n881 VSUBS 0.009391f
C922 B.n882 VSUBS 0.009391f
C923 B.n883 VSUBS 0.009391f
C924 B.n884 VSUBS 0.009391f
C925 B.n885 VSUBS 0.009391f
C926 B.n886 VSUBS 0.009391f
C927 B.n887 VSUBS 0.009391f
C928 B.n888 VSUBS 0.009391f
C929 B.n889 VSUBS 0.009391f
C930 B.n890 VSUBS 0.009391f
C931 B.n891 VSUBS 0.009391f
C932 B.n892 VSUBS 0.009391f
C933 B.n893 VSUBS 0.009391f
C934 B.n894 VSUBS 0.009391f
C935 B.n895 VSUBS 0.009391f
C936 B.n896 VSUBS 0.009391f
C937 B.n897 VSUBS 0.009391f
C938 B.n898 VSUBS 0.009391f
C939 B.n899 VSUBS 0.009391f
C940 B.n900 VSUBS 0.009391f
C941 B.n901 VSUBS 0.009391f
C942 B.n902 VSUBS 0.009391f
C943 B.n903 VSUBS 0.009391f
C944 B.n904 VSUBS 0.009391f
C945 B.n905 VSUBS 0.009391f
C946 B.n906 VSUBS 0.009391f
C947 B.n907 VSUBS 0.009391f
C948 B.n908 VSUBS 0.009391f
C949 B.n909 VSUBS 0.009391f
C950 B.n910 VSUBS 0.009391f
C951 B.n911 VSUBS 0.009391f
C952 B.n912 VSUBS 0.009391f
C953 B.n913 VSUBS 0.009391f
C954 B.n914 VSUBS 0.009391f
C955 B.n915 VSUBS 0.009391f
C956 B.n916 VSUBS 0.009391f
C957 B.n917 VSUBS 0.009391f
C958 B.n918 VSUBS 0.009391f
C959 B.n919 VSUBS 0.009391f
C960 B.n920 VSUBS 0.009391f
C961 B.n921 VSUBS 0.009391f
C962 B.n922 VSUBS 0.009391f
C963 B.n923 VSUBS 0.009391f
C964 B.n924 VSUBS 0.009391f
C965 B.n925 VSUBS 0.009391f
C966 B.n926 VSUBS 0.009391f
C967 B.n927 VSUBS 0.009391f
C968 B.n928 VSUBS 0.009391f
C969 B.n929 VSUBS 0.009391f
C970 B.n930 VSUBS 0.009391f
C971 B.n931 VSUBS 0.009391f
C972 B.n932 VSUBS 0.009391f
C973 B.n933 VSUBS 0.009391f
C974 B.n934 VSUBS 0.009391f
C975 B.n935 VSUBS 0.009391f
C976 B.n936 VSUBS 0.009391f
C977 B.n937 VSUBS 0.009391f
C978 B.n938 VSUBS 0.009391f
C979 B.n939 VSUBS 0.009391f
C980 B.n940 VSUBS 0.009391f
C981 B.n941 VSUBS 0.009391f
C982 B.n942 VSUBS 0.009391f
C983 B.n943 VSUBS 0.009391f
C984 B.n944 VSUBS 0.009391f
C985 B.n945 VSUBS 0.009391f
C986 B.n946 VSUBS 0.009391f
C987 B.n947 VSUBS 0.009391f
C988 B.n948 VSUBS 0.009391f
C989 B.n949 VSUBS 0.009391f
C990 B.n950 VSUBS 0.009391f
C991 B.n951 VSUBS 0.009391f
C992 B.n952 VSUBS 0.009391f
C993 B.n953 VSUBS 0.009391f
C994 B.n954 VSUBS 0.009391f
C995 B.n955 VSUBS 0.009391f
C996 B.n956 VSUBS 0.009391f
C997 B.n957 VSUBS 0.009391f
C998 B.n958 VSUBS 0.009391f
C999 B.n959 VSUBS 0.009391f
C1000 B.n960 VSUBS 0.009391f
C1001 B.n961 VSUBS 0.009391f
C1002 B.n962 VSUBS 0.009391f
C1003 B.n963 VSUBS 0.009391f
C1004 B.n964 VSUBS 0.009391f
C1005 B.n965 VSUBS 0.009391f
C1006 B.n966 VSUBS 0.009391f
C1007 B.n967 VSUBS 0.021265f
C1008 VDD2.t2 VSUBS 2.70456f
C1009 VDD2.t6 VSUBS 0.264822f
C1010 VDD2.t0 VSUBS 0.264822f
C1011 VDD2.n0 VSUBS 2.03488f
C1012 VDD2.n1 VSUBS 1.96733f
C1013 VDD2.t7 VSUBS 0.264822f
C1014 VDD2.t9 VSUBS 0.264822f
C1015 VDD2.n2 VSUBS 2.06974f
C1016 VDD2.n3 VSUBS 4.52392f
C1017 VDD2.t8 VSUBS 2.66543f
C1018 VDD2.n4 VSUBS 4.62353f
C1019 VDD2.t5 VSUBS 0.264822f
C1020 VDD2.t1 VSUBS 0.264822f
C1021 VDD2.n5 VSUBS 2.03489f
C1022 VDD2.n6 VSUBS 1.00236f
C1023 VDD2.t3 VSUBS 0.264822f
C1024 VDD2.t4 VSUBS 0.264822f
C1025 VDD2.n7 VSUBS 2.06968f
C1026 VN.t0 VSUBS 2.55919f
C1027 VN.n0 VSUBS 0.991371f
C1028 VN.n1 VSUBS 0.025062f
C1029 VN.n2 VSUBS 0.045771f
C1030 VN.n3 VSUBS 0.025062f
C1031 VN.n4 VSUBS 0.039592f
C1032 VN.n5 VSUBS 0.025062f
C1033 VN.n6 VSUBS 0.039898f
C1034 VN.n7 VSUBS 0.025062f
C1035 VN.n8 VSUBS 0.035003f
C1036 VN.n9 VSUBS 0.025062f
C1037 VN.n10 VSUBS 0.032964f
C1038 VN.n11 VSUBS 0.025062f
C1039 VN.n12 VSUBS 0.030414f
C1040 VN.t3 VSUBS 2.55919f
C1041 VN.n13 VSUBS 0.986056f
C1042 VN.t7 VSUBS 2.8962f
C1043 VN.n14 VSUBS 0.943094f
C1044 VN.n15 VSUBS 0.314052f
C1045 VN.n16 VSUBS 0.025062f
C1046 VN.n17 VSUBS 0.046475f
C1047 VN.n18 VSUBS 0.046475f
C1048 VN.n19 VSUBS 0.039898f
C1049 VN.n20 VSUBS 0.025062f
C1050 VN.n21 VSUBS 0.025062f
C1051 VN.n22 VSUBS 0.025062f
C1052 VN.n23 VSUBS 0.046475f
C1053 VN.n24 VSUBS 0.046475f
C1054 VN.t9 VSUBS 2.55919f
C1055 VN.n25 VSUBS 0.903867f
C1056 VN.n26 VSUBS 0.035003f
C1057 VN.n27 VSUBS 0.025062f
C1058 VN.n28 VSUBS 0.025062f
C1059 VN.n29 VSUBS 0.025062f
C1060 VN.n30 VSUBS 0.046475f
C1061 VN.n31 VSUBS 0.046475f
C1062 VN.n32 VSUBS 0.032964f
C1063 VN.n33 VSUBS 0.025062f
C1064 VN.n34 VSUBS 0.025062f
C1065 VN.n35 VSUBS 0.025062f
C1066 VN.n36 VSUBS 0.046475f
C1067 VN.n37 VSUBS 0.046475f
C1068 VN.t2 VSUBS 2.55919f
C1069 VN.n38 VSUBS 0.903867f
C1070 VN.n39 VSUBS 0.030414f
C1071 VN.n40 VSUBS 0.025062f
C1072 VN.n41 VSUBS 0.025062f
C1073 VN.n42 VSUBS 0.025062f
C1074 VN.n43 VSUBS 0.046475f
C1075 VN.n44 VSUBS 0.049936f
C1076 VN.n45 VSUBS 0.023629f
C1077 VN.n46 VSUBS 0.025062f
C1078 VN.n47 VSUBS 0.025062f
C1079 VN.n48 VSUBS 0.025062f
C1080 VN.n49 VSUBS 0.046475f
C1081 VN.n50 VSUBS 0.046475f
C1082 VN.n51 VSUBS 0.025826f
C1083 VN.n52 VSUBS 0.040443f
C1084 VN.n53 VSUBS 0.073972f
C1085 VN.t1 VSUBS 2.55919f
C1086 VN.n54 VSUBS 0.991371f
C1087 VN.n55 VSUBS 0.025062f
C1088 VN.n56 VSUBS 0.045771f
C1089 VN.n57 VSUBS 0.025062f
C1090 VN.n58 VSUBS 0.039592f
C1091 VN.n59 VSUBS 0.025062f
C1092 VN.t4 VSUBS 2.55919f
C1093 VN.n60 VSUBS 0.903867f
C1094 VN.n61 VSUBS 0.039898f
C1095 VN.n62 VSUBS 0.025062f
C1096 VN.n63 VSUBS 0.035003f
C1097 VN.n64 VSUBS 0.025062f
C1098 VN.t8 VSUBS 2.55919f
C1099 VN.n65 VSUBS 0.903867f
C1100 VN.n66 VSUBS 0.032964f
C1101 VN.n67 VSUBS 0.025062f
C1102 VN.n68 VSUBS 0.030414f
C1103 VN.t5 VSUBS 2.8962f
C1104 VN.t6 VSUBS 2.55919f
C1105 VN.n69 VSUBS 0.986056f
C1106 VN.n70 VSUBS 0.943094f
C1107 VN.n71 VSUBS 0.314052f
C1108 VN.n72 VSUBS 0.025062f
C1109 VN.n73 VSUBS 0.046475f
C1110 VN.n74 VSUBS 0.046475f
C1111 VN.n75 VSUBS 0.039898f
C1112 VN.n76 VSUBS 0.025062f
C1113 VN.n77 VSUBS 0.025062f
C1114 VN.n78 VSUBS 0.025062f
C1115 VN.n79 VSUBS 0.046475f
C1116 VN.n80 VSUBS 0.046475f
C1117 VN.n81 VSUBS 0.035003f
C1118 VN.n82 VSUBS 0.025062f
C1119 VN.n83 VSUBS 0.025062f
C1120 VN.n84 VSUBS 0.025062f
C1121 VN.n85 VSUBS 0.046475f
C1122 VN.n86 VSUBS 0.046475f
C1123 VN.n87 VSUBS 0.032964f
C1124 VN.n88 VSUBS 0.025062f
C1125 VN.n89 VSUBS 0.025062f
C1126 VN.n90 VSUBS 0.025062f
C1127 VN.n91 VSUBS 0.046475f
C1128 VN.n92 VSUBS 0.046475f
C1129 VN.n93 VSUBS 0.030414f
C1130 VN.n94 VSUBS 0.025062f
C1131 VN.n95 VSUBS 0.025062f
C1132 VN.n96 VSUBS 0.025062f
C1133 VN.n97 VSUBS 0.046475f
C1134 VN.n98 VSUBS 0.049936f
C1135 VN.n99 VSUBS 0.023629f
C1136 VN.n100 VSUBS 0.025062f
C1137 VN.n101 VSUBS 0.025062f
C1138 VN.n102 VSUBS 0.025062f
C1139 VN.n103 VSUBS 0.046475f
C1140 VN.n104 VSUBS 0.046475f
C1141 VN.n105 VSUBS 0.025826f
C1142 VN.n106 VSUBS 0.040443f
C1143 VN.n107 VSUBS 1.7447f
C1144 VTAIL.t1 VSUBS 0.254958f
C1145 VTAIL.t0 VSUBS 0.254958f
C1146 VTAIL.n0 VSUBS 1.81876f
C1147 VTAIL.n1 VSUBS 1.11009f
C1148 VTAIL.t15 VSUBS 2.41033f
C1149 VTAIL.n2 VSUBS 1.29103f
C1150 VTAIL.t11 VSUBS 0.254958f
C1151 VTAIL.t18 VSUBS 0.254958f
C1152 VTAIL.n3 VSUBS 1.81876f
C1153 VTAIL.n4 VSUBS 1.30672f
C1154 VTAIL.t13 VSUBS 0.254958f
C1155 VTAIL.t19 VSUBS 0.254958f
C1156 VTAIL.n5 VSUBS 1.81876f
C1157 VTAIL.n6 VSUBS 2.95037f
C1158 VTAIL.t9 VSUBS 0.254958f
C1159 VTAIL.t8 VSUBS 0.254958f
C1160 VTAIL.n7 VSUBS 1.81877f
C1161 VTAIL.n8 VSUBS 2.95036f
C1162 VTAIL.t6 VSUBS 0.254958f
C1163 VTAIL.t4 VSUBS 0.254958f
C1164 VTAIL.n9 VSUBS 1.81877f
C1165 VTAIL.n10 VSUBS 1.30672f
C1166 VTAIL.t3 VSUBS 2.41034f
C1167 VTAIL.n11 VSUBS 1.29102f
C1168 VTAIL.t12 VSUBS 0.254958f
C1169 VTAIL.t10 VSUBS 0.254958f
C1170 VTAIL.n12 VSUBS 1.81877f
C1171 VTAIL.n13 VSUBS 1.18725f
C1172 VTAIL.t14 VSUBS 0.254958f
C1173 VTAIL.t17 VSUBS 0.254958f
C1174 VTAIL.n14 VSUBS 1.81877f
C1175 VTAIL.n15 VSUBS 1.30672f
C1176 VTAIL.t16 VSUBS 2.41033f
C1177 VTAIL.n16 VSUBS 2.72252f
C1178 VTAIL.t5 VSUBS 2.41033f
C1179 VTAIL.n17 VSUBS 2.72252f
C1180 VTAIL.t7 VSUBS 0.254958f
C1181 VTAIL.t2 VSUBS 0.254958f
C1182 VTAIL.n18 VSUBS 1.81876f
C1183 VTAIL.n19 VSUBS 1.05227f
C1184 VDD1.t5 VSUBS 2.70296f
C1185 VDD1.t4 VSUBS 0.264665f
C1186 VDD1.t7 VSUBS 0.264665f
C1187 VDD1.n0 VSUBS 2.03368f
C1188 VDD1.n1 VSUBS 1.97684f
C1189 VDD1.t6 VSUBS 2.70295f
C1190 VDD1.t9 VSUBS 0.264665f
C1191 VDD1.t3 VSUBS 0.264665f
C1192 VDD1.n2 VSUBS 2.03368f
C1193 VDD1.n3 VSUBS 1.96616f
C1194 VDD1.t8 VSUBS 0.264665f
C1195 VDD1.t0 VSUBS 0.264665f
C1196 VDD1.n4 VSUBS 2.06851f
C1197 VDD1.n5 VSUBS 4.71257f
C1198 VDD1.t2 VSUBS 0.264665f
C1199 VDD1.t1 VSUBS 0.264665f
C1200 VDD1.n6 VSUBS 2.03367f
C1201 VDD1.n7 VSUBS 4.70741f
C1202 VP.t4 VSUBS 2.80551f
C1203 VP.n0 VSUBS 1.08679f
C1204 VP.n1 VSUBS 0.027474f
C1205 VP.n2 VSUBS 0.050177f
C1206 VP.n3 VSUBS 0.027474f
C1207 VP.n4 VSUBS 0.043402f
C1208 VP.n5 VSUBS 0.027474f
C1209 VP.n6 VSUBS 0.043738f
C1210 VP.n7 VSUBS 0.027474f
C1211 VP.n8 VSUBS 0.038372f
C1212 VP.n9 VSUBS 0.027474f
C1213 VP.n10 VSUBS 0.036137f
C1214 VP.n11 VSUBS 0.027474f
C1215 VP.n12 VSUBS 0.033342f
C1216 VP.n13 VSUBS 0.027474f
C1217 VP.n14 VSUBS 0.025904f
C1218 VP.n15 VSUBS 0.027474f
C1219 VP.n16 VSUBS 0.028311f
C1220 VP.t3 VSUBS 2.80551f
C1221 VP.n17 VSUBS 1.08679f
C1222 VP.n18 VSUBS 0.027474f
C1223 VP.n19 VSUBS 0.050177f
C1224 VP.n20 VSUBS 0.027474f
C1225 VP.n21 VSUBS 0.043402f
C1226 VP.n22 VSUBS 0.027474f
C1227 VP.n23 VSUBS 0.043738f
C1228 VP.n24 VSUBS 0.027474f
C1229 VP.n25 VSUBS 0.038372f
C1230 VP.n26 VSUBS 0.027474f
C1231 VP.n27 VSUBS 0.036137f
C1232 VP.n28 VSUBS 0.027474f
C1233 VP.n29 VSUBS 0.033342f
C1234 VP.t7 VSUBS 3.17495f
C1235 VP.t9 VSUBS 2.80551f
C1236 VP.n30 VSUBS 1.08096f
C1237 VP.n31 VSUBS 1.03386f
C1238 VP.n32 VSUBS 0.344279f
C1239 VP.n33 VSUBS 0.027474f
C1240 VP.n34 VSUBS 0.050948f
C1241 VP.n35 VSUBS 0.050948f
C1242 VP.n36 VSUBS 0.043738f
C1243 VP.n37 VSUBS 0.027474f
C1244 VP.n38 VSUBS 0.027474f
C1245 VP.n39 VSUBS 0.027474f
C1246 VP.n40 VSUBS 0.050948f
C1247 VP.n41 VSUBS 0.050948f
C1248 VP.t5 VSUBS 2.80551f
C1249 VP.n42 VSUBS 0.990862f
C1250 VP.n43 VSUBS 0.038372f
C1251 VP.n44 VSUBS 0.027474f
C1252 VP.n45 VSUBS 0.027474f
C1253 VP.n46 VSUBS 0.027474f
C1254 VP.n47 VSUBS 0.050948f
C1255 VP.n48 VSUBS 0.050948f
C1256 VP.n49 VSUBS 0.036137f
C1257 VP.n50 VSUBS 0.027474f
C1258 VP.n51 VSUBS 0.027474f
C1259 VP.n52 VSUBS 0.027474f
C1260 VP.n53 VSUBS 0.050948f
C1261 VP.n54 VSUBS 0.050948f
C1262 VP.t2 VSUBS 2.80551f
C1263 VP.n55 VSUBS 0.990862f
C1264 VP.n56 VSUBS 0.033342f
C1265 VP.n57 VSUBS 0.027474f
C1266 VP.n58 VSUBS 0.027474f
C1267 VP.n59 VSUBS 0.027474f
C1268 VP.n60 VSUBS 0.050948f
C1269 VP.n61 VSUBS 0.054742f
C1270 VP.n62 VSUBS 0.025904f
C1271 VP.n63 VSUBS 0.027474f
C1272 VP.n64 VSUBS 0.027474f
C1273 VP.n65 VSUBS 0.027474f
C1274 VP.n66 VSUBS 0.050948f
C1275 VP.n67 VSUBS 0.050948f
C1276 VP.n68 VSUBS 0.028311f
C1277 VP.n69 VSUBS 0.044335f
C1278 VP.n70 VSUBS 1.90187f
C1279 VP.t6 VSUBS 2.80551f
C1280 VP.n71 VSUBS 1.08679f
C1281 VP.n72 VSUBS 1.91916f
C1282 VP.n73 VSUBS 0.044335f
C1283 VP.n74 VSUBS 0.027474f
C1284 VP.n75 VSUBS 0.050948f
C1285 VP.n76 VSUBS 0.050948f
C1286 VP.n77 VSUBS 0.050177f
C1287 VP.n78 VSUBS 0.027474f
C1288 VP.n79 VSUBS 0.027474f
C1289 VP.n80 VSUBS 0.027474f
C1290 VP.n81 VSUBS 0.054742f
C1291 VP.n82 VSUBS 0.050948f
C1292 VP.t0 VSUBS 2.80551f
C1293 VP.n83 VSUBS 0.990862f
C1294 VP.n84 VSUBS 0.043402f
C1295 VP.n85 VSUBS 0.027474f
C1296 VP.n86 VSUBS 0.027474f
C1297 VP.n87 VSUBS 0.027474f
C1298 VP.n88 VSUBS 0.050948f
C1299 VP.n89 VSUBS 0.050948f
C1300 VP.n90 VSUBS 0.043738f
C1301 VP.n91 VSUBS 0.027474f
C1302 VP.n92 VSUBS 0.027474f
C1303 VP.n93 VSUBS 0.027474f
C1304 VP.n94 VSUBS 0.050948f
C1305 VP.n95 VSUBS 0.050948f
C1306 VP.t8 VSUBS 2.80551f
C1307 VP.n96 VSUBS 0.990862f
C1308 VP.n97 VSUBS 0.038372f
C1309 VP.n98 VSUBS 0.027474f
C1310 VP.n99 VSUBS 0.027474f
C1311 VP.n100 VSUBS 0.027474f
C1312 VP.n101 VSUBS 0.050948f
C1313 VP.n102 VSUBS 0.050948f
C1314 VP.n103 VSUBS 0.036137f
C1315 VP.n104 VSUBS 0.027474f
C1316 VP.n105 VSUBS 0.027474f
C1317 VP.n106 VSUBS 0.027474f
C1318 VP.n107 VSUBS 0.050948f
C1319 VP.n108 VSUBS 0.050948f
C1320 VP.t1 VSUBS 2.80551f
C1321 VP.n109 VSUBS 0.990862f
C1322 VP.n110 VSUBS 0.033342f
C1323 VP.n111 VSUBS 0.027474f
C1324 VP.n112 VSUBS 0.027474f
C1325 VP.n113 VSUBS 0.027474f
C1326 VP.n114 VSUBS 0.050948f
C1327 VP.n115 VSUBS 0.054742f
C1328 VP.n116 VSUBS 0.025904f
C1329 VP.n117 VSUBS 0.027474f
C1330 VP.n118 VSUBS 0.027474f
C1331 VP.n119 VSUBS 0.027474f
C1332 VP.n120 VSUBS 0.050948f
C1333 VP.n121 VSUBS 0.050948f
C1334 VP.n122 VSUBS 0.028311f
C1335 VP.n123 VSUBS 0.044335f
C1336 VP.n124 VSUBS 0.081091f
.ends

