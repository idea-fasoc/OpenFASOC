* NGSPICE file created from diff_pair_sample_0344.ext - technology: sky130A

.subckt diff_pair_sample_0344 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=2.23
X1 VTAIL.t11 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=2.23
X2 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=2.23
X3 VDD2.t0 VN.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=2.23
X4 VTAIL.t5 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=2.23
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=2.23
X6 VTAIL.t9 VN.t2 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=2.23
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=2.23
X8 VDD2.t4 VN.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=2.23
X9 VDD1.t3 VP.t2 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=2.23
X10 VDD1.t2 VP.t3 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=2.23
X11 VTAIL.t1 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=2.23
X12 VDD2.t5 VN.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=2.23
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=2.23
X14 VDD2.t2 VN.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=2.23
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=2.23
R0 B.n729 B.n144 585
R1 B.n144 B.n71 585
R2 B.n731 B.n730 585
R3 B.n733 B.n143 585
R4 B.n736 B.n735 585
R5 B.n737 B.n142 585
R6 B.n739 B.n738 585
R7 B.n741 B.n141 585
R8 B.n744 B.n743 585
R9 B.n745 B.n140 585
R10 B.n747 B.n746 585
R11 B.n749 B.n139 585
R12 B.n752 B.n751 585
R13 B.n753 B.n138 585
R14 B.n755 B.n754 585
R15 B.n757 B.n137 585
R16 B.n760 B.n759 585
R17 B.n761 B.n136 585
R18 B.n763 B.n762 585
R19 B.n765 B.n135 585
R20 B.n768 B.n767 585
R21 B.n769 B.n134 585
R22 B.n771 B.n770 585
R23 B.n773 B.n133 585
R24 B.n776 B.n775 585
R25 B.n777 B.n132 585
R26 B.n779 B.n778 585
R27 B.n781 B.n131 585
R28 B.n784 B.n783 585
R29 B.n785 B.n130 585
R30 B.n787 B.n786 585
R31 B.n789 B.n129 585
R32 B.n792 B.n791 585
R33 B.n793 B.n128 585
R34 B.n795 B.n794 585
R35 B.n797 B.n127 585
R36 B.n800 B.n799 585
R37 B.n801 B.n126 585
R38 B.n803 B.n802 585
R39 B.n805 B.n125 585
R40 B.n808 B.n807 585
R41 B.n809 B.n124 585
R42 B.n811 B.n810 585
R43 B.n813 B.n123 585
R44 B.n816 B.n815 585
R45 B.n817 B.n122 585
R46 B.n819 B.n818 585
R47 B.n821 B.n121 585
R48 B.n824 B.n823 585
R49 B.n825 B.n120 585
R50 B.n827 B.n826 585
R51 B.n829 B.n119 585
R52 B.n832 B.n831 585
R53 B.n833 B.n118 585
R54 B.n835 B.n834 585
R55 B.n837 B.n117 585
R56 B.n840 B.n839 585
R57 B.n841 B.n116 585
R58 B.n843 B.n842 585
R59 B.n845 B.n115 585
R60 B.n848 B.n847 585
R61 B.n849 B.n114 585
R62 B.n851 B.n850 585
R63 B.n853 B.n113 585
R64 B.n856 B.n855 585
R65 B.n858 B.n110 585
R66 B.n860 B.n859 585
R67 B.n862 B.n109 585
R68 B.n865 B.n864 585
R69 B.n866 B.n108 585
R70 B.n868 B.n867 585
R71 B.n870 B.n107 585
R72 B.n873 B.n872 585
R73 B.n874 B.n104 585
R74 B.n877 B.n876 585
R75 B.n879 B.n103 585
R76 B.n882 B.n881 585
R77 B.n883 B.n102 585
R78 B.n885 B.n884 585
R79 B.n887 B.n101 585
R80 B.n890 B.n889 585
R81 B.n891 B.n100 585
R82 B.n893 B.n892 585
R83 B.n895 B.n99 585
R84 B.n898 B.n897 585
R85 B.n899 B.n98 585
R86 B.n901 B.n900 585
R87 B.n903 B.n97 585
R88 B.n906 B.n905 585
R89 B.n907 B.n96 585
R90 B.n909 B.n908 585
R91 B.n911 B.n95 585
R92 B.n914 B.n913 585
R93 B.n915 B.n94 585
R94 B.n917 B.n916 585
R95 B.n919 B.n93 585
R96 B.n922 B.n921 585
R97 B.n923 B.n92 585
R98 B.n925 B.n924 585
R99 B.n927 B.n91 585
R100 B.n930 B.n929 585
R101 B.n931 B.n90 585
R102 B.n933 B.n932 585
R103 B.n935 B.n89 585
R104 B.n938 B.n937 585
R105 B.n939 B.n88 585
R106 B.n941 B.n940 585
R107 B.n943 B.n87 585
R108 B.n946 B.n945 585
R109 B.n947 B.n86 585
R110 B.n949 B.n948 585
R111 B.n951 B.n85 585
R112 B.n954 B.n953 585
R113 B.n955 B.n84 585
R114 B.n957 B.n956 585
R115 B.n959 B.n83 585
R116 B.n962 B.n961 585
R117 B.n963 B.n82 585
R118 B.n965 B.n964 585
R119 B.n967 B.n81 585
R120 B.n970 B.n969 585
R121 B.n971 B.n80 585
R122 B.n973 B.n972 585
R123 B.n975 B.n79 585
R124 B.n978 B.n977 585
R125 B.n979 B.n78 585
R126 B.n981 B.n980 585
R127 B.n983 B.n77 585
R128 B.n986 B.n985 585
R129 B.n987 B.n76 585
R130 B.n989 B.n988 585
R131 B.n991 B.n75 585
R132 B.n994 B.n993 585
R133 B.n995 B.n74 585
R134 B.n997 B.n996 585
R135 B.n999 B.n73 585
R136 B.n1002 B.n1001 585
R137 B.n1003 B.n72 585
R138 B.n728 B.n70 585
R139 B.n1006 B.n70 585
R140 B.n727 B.n69 585
R141 B.n1007 B.n69 585
R142 B.n726 B.n68 585
R143 B.n1008 B.n68 585
R144 B.n725 B.n724 585
R145 B.n724 B.n64 585
R146 B.n723 B.n63 585
R147 B.n1014 B.n63 585
R148 B.n722 B.n62 585
R149 B.n1015 B.n62 585
R150 B.n721 B.n61 585
R151 B.n1016 B.n61 585
R152 B.n720 B.n719 585
R153 B.n719 B.n57 585
R154 B.n718 B.n56 585
R155 B.n1022 B.n56 585
R156 B.n717 B.n55 585
R157 B.n1023 B.n55 585
R158 B.n716 B.n54 585
R159 B.n1024 B.n54 585
R160 B.n715 B.n714 585
R161 B.n714 B.n50 585
R162 B.n713 B.n49 585
R163 B.n1030 B.n49 585
R164 B.n712 B.n48 585
R165 B.n1031 B.n48 585
R166 B.n711 B.n47 585
R167 B.n1032 B.n47 585
R168 B.n710 B.n709 585
R169 B.n709 B.n43 585
R170 B.n708 B.n42 585
R171 B.n1038 B.n42 585
R172 B.n707 B.n41 585
R173 B.n1039 B.n41 585
R174 B.n706 B.n40 585
R175 B.n1040 B.n40 585
R176 B.n705 B.n704 585
R177 B.n704 B.n36 585
R178 B.n703 B.n35 585
R179 B.n1046 B.n35 585
R180 B.n702 B.n34 585
R181 B.n1047 B.n34 585
R182 B.n701 B.n33 585
R183 B.n1048 B.n33 585
R184 B.n700 B.n699 585
R185 B.n699 B.n29 585
R186 B.n698 B.n28 585
R187 B.n1054 B.n28 585
R188 B.n697 B.n27 585
R189 B.n1055 B.n27 585
R190 B.n696 B.n26 585
R191 B.n1056 B.n26 585
R192 B.n695 B.n694 585
R193 B.n694 B.n22 585
R194 B.n693 B.n21 585
R195 B.n1062 B.n21 585
R196 B.n692 B.n20 585
R197 B.n1063 B.n20 585
R198 B.n691 B.n19 585
R199 B.n1064 B.n19 585
R200 B.n690 B.n689 585
R201 B.n689 B.n15 585
R202 B.n688 B.n14 585
R203 B.n1070 B.n14 585
R204 B.n687 B.n13 585
R205 B.n1071 B.n13 585
R206 B.n686 B.n12 585
R207 B.n1072 B.n12 585
R208 B.n685 B.n684 585
R209 B.n684 B.n8 585
R210 B.n683 B.n7 585
R211 B.n1078 B.n7 585
R212 B.n682 B.n6 585
R213 B.n1079 B.n6 585
R214 B.n681 B.n5 585
R215 B.n1080 B.n5 585
R216 B.n680 B.n679 585
R217 B.n679 B.n4 585
R218 B.n678 B.n145 585
R219 B.n678 B.n677 585
R220 B.n668 B.n146 585
R221 B.n147 B.n146 585
R222 B.n670 B.n669 585
R223 B.n671 B.n670 585
R224 B.n667 B.n152 585
R225 B.n152 B.n151 585
R226 B.n666 B.n665 585
R227 B.n665 B.n664 585
R228 B.n154 B.n153 585
R229 B.n155 B.n154 585
R230 B.n657 B.n656 585
R231 B.n658 B.n657 585
R232 B.n655 B.n160 585
R233 B.n160 B.n159 585
R234 B.n654 B.n653 585
R235 B.n653 B.n652 585
R236 B.n162 B.n161 585
R237 B.n163 B.n162 585
R238 B.n645 B.n644 585
R239 B.n646 B.n645 585
R240 B.n643 B.n167 585
R241 B.n171 B.n167 585
R242 B.n642 B.n641 585
R243 B.n641 B.n640 585
R244 B.n169 B.n168 585
R245 B.n170 B.n169 585
R246 B.n633 B.n632 585
R247 B.n634 B.n633 585
R248 B.n631 B.n176 585
R249 B.n176 B.n175 585
R250 B.n630 B.n629 585
R251 B.n629 B.n628 585
R252 B.n178 B.n177 585
R253 B.n179 B.n178 585
R254 B.n621 B.n620 585
R255 B.n622 B.n621 585
R256 B.n619 B.n183 585
R257 B.n187 B.n183 585
R258 B.n618 B.n617 585
R259 B.n617 B.n616 585
R260 B.n185 B.n184 585
R261 B.n186 B.n185 585
R262 B.n609 B.n608 585
R263 B.n610 B.n609 585
R264 B.n607 B.n192 585
R265 B.n192 B.n191 585
R266 B.n606 B.n605 585
R267 B.n605 B.n604 585
R268 B.n194 B.n193 585
R269 B.n195 B.n194 585
R270 B.n597 B.n596 585
R271 B.n598 B.n597 585
R272 B.n595 B.n200 585
R273 B.n200 B.n199 585
R274 B.n594 B.n593 585
R275 B.n593 B.n592 585
R276 B.n202 B.n201 585
R277 B.n203 B.n202 585
R278 B.n585 B.n584 585
R279 B.n586 B.n585 585
R280 B.n583 B.n208 585
R281 B.n208 B.n207 585
R282 B.n582 B.n581 585
R283 B.n581 B.n580 585
R284 B.n210 B.n209 585
R285 B.n211 B.n210 585
R286 B.n573 B.n572 585
R287 B.n574 B.n573 585
R288 B.n571 B.n216 585
R289 B.n216 B.n215 585
R290 B.n570 B.n569 585
R291 B.n569 B.n568 585
R292 B.n565 B.n220 585
R293 B.n564 B.n563 585
R294 B.n561 B.n221 585
R295 B.n561 B.n219 585
R296 B.n560 B.n559 585
R297 B.n558 B.n557 585
R298 B.n556 B.n223 585
R299 B.n554 B.n553 585
R300 B.n552 B.n224 585
R301 B.n551 B.n550 585
R302 B.n548 B.n225 585
R303 B.n546 B.n545 585
R304 B.n544 B.n226 585
R305 B.n543 B.n542 585
R306 B.n540 B.n227 585
R307 B.n538 B.n537 585
R308 B.n536 B.n228 585
R309 B.n535 B.n534 585
R310 B.n532 B.n229 585
R311 B.n530 B.n529 585
R312 B.n528 B.n230 585
R313 B.n527 B.n526 585
R314 B.n524 B.n231 585
R315 B.n522 B.n521 585
R316 B.n520 B.n232 585
R317 B.n519 B.n518 585
R318 B.n516 B.n233 585
R319 B.n514 B.n513 585
R320 B.n512 B.n234 585
R321 B.n511 B.n510 585
R322 B.n508 B.n235 585
R323 B.n506 B.n505 585
R324 B.n504 B.n236 585
R325 B.n503 B.n502 585
R326 B.n500 B.n237 585
R327 B.n498 B.n497 585
R328 B.n496 B.n238 585
R329 B.n495 B.n494 585
R330 B.n492 B.n239 585
R331 B.n490 B.n489 585
R332 B.n488 B.n240 585
R333 B.n487 B.n486 585
R334 B.n484 B.n241 585
R335 B.n482 B.n481 585
R336 B.n480 B.n242 585
R337 B.n479 B.n478 585
R338 B.n476 B.n243 585
R339 B.n474 B.n473 585
R340 B.n472 B.n244 585
R341 B.n471 B.n470 585
R342 B.n468 B.n245 585
R343 B.n466 B.n465 585
R344 B.n464 B.n246 585
R345 B.n463 B.n462 585
R346 B.n460 B.n247 585
R347 B.n458 B.n457 585
R348 B.n456 B.n248 585
R349 B.n455 B.n454 585
R350 B.n452 B.n249 585
R351 B.n450 B.n449 585
R352 B.n448 B.n250 585
R353 B.n447 B.n446 585
R354 B.n444 B.n251 585
R355 B.n442 B.n441 585
R356 B.n440 B.n252 585
R357 B.n438 B.n437 585
R358 B.n435 B.n255 585
R359 B.n433 B.n432 585
R360 B.n431 B.n256 585
R361 B.n430 B.n429 585
R362 B.n427 B.n257 585
R363 B.n425 B.n424 585
R364 B.n423 B.n258 585
R365 B.n422 B.n421 585
R366 B.n419 B.n418 585
R367 B.n417 B.n416 585
R368 B.n415 B.n263 585
R369 B.n413 B.n412 585
R370 B.n411 B.n264 585
R371 B.n410 B.n409 585
R372 B.n407 B.n265 585
R373 B.n405 B.n404 585
R374 B.n403 B.n266 585
R375 B.n402 B.n401 585
R376 B.n399 B.n267 585
R377 B.n397 B.n396 585
R378 B.n395 B.n268 585
R379 B.n394 B.n393 585
R380 B.n391 B.n269 585
R381 B.n389 B.n388 585
R382 B.n387 B.n270 585
R383 B.n386 B.n385 585
R384 B.n383 B.n271 585
R385 B.n381 B.n380 585
R386 B.n379 B.n272 585
R387 B.n378 B.n377 585
R388 B.n375 B.n273 585
R389 B.n373 B.n372 585
R390 B.n371 B.n274 585
R391 B.n370 B.n369 585
R392 B.n367 B.n275 585
R393 B.n365 B.n364 585
R394 B.n363 B.n276 585
R395 B.n362 B.n361 585
R396 B.n359 B.n277 585
R397 B.n357 B.n356 585
R398 B.n355 B.n278 585
R399 B.n354 B.n353 585
R400 B.n351 B.n279 585
R401 B.n349 B.n348 585
R402 B.n347 B.n280 585
R403 B.n346 B.n345 585
R404 B.n343 B.n281 585
R405 B.n341 B.n340 585
R406 B.n339 B.n282 585
R407 B.n338 B.n337 585
R408 B.n335 B.n283 585
R409 B.n333 B.n332 585
R410 B.n331 B.n284 585
R411 B.n330 B.n329 585
R412 B.n327 B.n285 585
R413 B.n325 B.n324 585
R414 B.n323 B.n286 585
R415 B.n322 B.n321 585
R416 B.n319 B.n287 585
R417 B.n317 B.n316 585
R418 B.n315 B.n288 585
R419 B.n314 B.n313 585
R420 B.n311 B.n289 585
R421 B.n309 B.n308 585
R422 B.n307 B.n290 585
R423 B.n306 B.n305 585
R424 B.n303 B.n291 585
R425 B.n301 B.n300 585
R426 B.n299 B.n292 585
R427 B.n298 B.n297 585
R428 B.n295 B.n293 585
R429 B.n218 B.n217 585
R430 B.n567 B.n566 585
R431 B.n568 B.n567 585
R432 B.n214 B.n213 585
R433 B.n215 B.n214 585
R434 B.n576 B.n575 585
R435 B.n575 B.n574 585
R436 B.n577 B.n212 585
R437 B.n212 B.n211 585
R438 B.n579 B.n578 585
R439 B.n580 B.n579 585
R440 B.n206 B.n205 585
R441 B.n207 B.n206 585
R442 B.n588 B.n587 585
R443 B.n587 B.n586 585
R444 B.n589 B.n204 585
R445 B.n204 B.n203 585
R446 B.n591 B.n590 585
R447 B.n592 B.n591 585
R448 B.n198 B.n197 585
R449 B.n199 B.n198 585
R450 B.n600 B.n599 585
R451 B.n599 B.n598 585
R452 B.n601 B.n196 585
R453 B.n196 B.n195 585
R454 B.n603 B.n602 585
R455 B.n604 B.n603 585
R456 B.n190 B.n189 585
R457 B.n191 B.n190 585
R458 B.n612 B.n611 585
R459 B.n611 B.n610 585
R460 B.n613 B.n188 585
R461 B.n188 B.n186 585
R462 B.n615 B.n614 585
R463 B.n616 B.n615 585
R464 B.n182 B.n181 585
R465 B.n187 B.n182 585
R466 B.n624 B.n623 585
R467 B.n623 B.n622 585
R468 B.n625 B.n180 585
R469 B.n180 B.n179 585
R470 B.n627 B.n626 585
R471 B.n628 B.n627 585
R472 B.n174 B.n173 585
R473 B.n175 B.n174 585
R474 B.n636 B.n635 585
R475 B.n635 B.n634 585
R476 B.n637 B.n172 585
R477 B.n172 B.n170 585
R478 B.n639 B.n638 585
R479 B.n640 B.n639 585
R480 B.n166 B.n165 585
R481 B.n171 B.n166 585
R482 B.n648 B.n647 585
R483 B.n647 B.n646 585
R484 B.n649 B.n164 585
R485 B.n164 B.n163 585
R486 B.n651 B.n650 585
R487 B.n652 B.n651 585
R488 B.n158 B.n157 585
R489 B.n159 B.n158 585
R490 B.n660 B.n659 585
R491 B.n659 B.n658 585
R492 B.n661 B.n156 585
R493 B.n156 B.n155 585
R494 B.n663 B.n662 585
R495 B.n664 B.n663 585
R496 B.n150 B.n149 585
R497 B.n151 B.n150 585
R498 B.n673 B.n672 585
R499 B.n672 B.n671 585
R500 B.n674 B.n148 585
R501 B.n148 B.n147 585
R502 B.n676 B.n675 585
R503 B.n677 B.n676 585
R504 B.n2 B.n0 585
R505 B.n4 B.n2 585
R506 B.n3 B.n1 585
R507 B.n1079 B.n3 585
R508 B.n1077 B.n1076 585
R509 B.n1078 B.n1077 585
R510 B.n1075 B.n9 585
R511 B.n9 B.n8 585
R512 B.n1074 B.n1073 585
R513 B.n1073 B.n1072 585
R514 B.n11 B.n10 585
R515 B.n1071 B.n11 585
R516 B.n1069 B.n1068 585
R517 B.n1070 B.n1069 585
R518 B.n1067 B.n16 585
R519 B.n16 B.n15 585
R520 B.n1066 B.n1065 585
R521 B.n1065 B.n1064 585
R522 B.n18 B.n17 585
R523 B.n1063 B.n18 585
R524 B.n1061 B.n1060 585
R525 B.n1062 B.n1061 585
R526 B.n1059 B.n23 585
R527 B.n23 B.n22 585
R528 B.n1058 B.n1057 585
R529 B.n1057 B.n1056 585
R530 B.n25 B.n24 585
R531 B.n1055 B.n25 585
R532 B.n1053 B.n1052 585
R533 B.n1054 B.n1053 585
R534 B.n1051 B.n30 585
R535 B.n30 B.n29 585
R536 B.n1050 B.n1049 585
R537 B.n1049 B.n1048 585
R538 B.n32 B.n31 585
R539 B.n1047 B.n32 585
R540 B.n1045 B.n1044 585
R541 B.n1046 B.n1045 585
R542 B.n1043 B.n37 585
R543 B.n37 B.n36 585
R544 B.n1042 B.n1041 585
R545 B.n1041 B.n1040 585
R546 B.n39 B.n38 585
R547 B.n1039 B.n39 585
R548 B.n1037 B.n1036 585
R549 B.n1038 B.n1037 585
R550 B.n1035 B.n44 585
R551 B.n44 B.n43 585
R552 B.n1034 B.n1033 585
R553 B.n1033 B.n1032 585
R554 B.n46 B.n45 585
R555 B.n1031 B.n46 585
R556 B.n1029 B.n1028 585
R557 B.n1030 B.n1029 585
R558 B.n1027 B.n51 585
R559 B.n51 B.n50 585
R560 B.n1026 B.n1025 585
R561 B.n1025 B.n1024 585
R562 B.n53 B.n52 585
R563 B.n1023 B.n53 585
R564 B.n1021 B.n1020 585
R565 B.n1022 B.n1021 585
R566 B.n1019 B.n58 585
R567 B.n58 B.n57 585
R568 B.n1018 B.n1017 585
R569 B.n1017 B.n1016 585
R570 B.n60 B.n59 585
R571 B.n1015 B.n60 585
R572 B.n1013 B.n1012 585
R573 B.n1014 B.n1013 585
R574 B.n1011 B.n65 585
R575 B.n65 B.n64 585
R576 B.n1010 B.n1009 585
R577 B.n1009 B.n1008 585
R578 B.n67 B.n66 585
R579 B.n1007 B.n67 585
R580 B.n1005 B.n1004 585
R581 B.n1006 B.n1005 585
R582 B.n1082 B.n1081 585
R583 B.n1081 B.n1080 585
R584 B.n567 B.n220 540.549
R585 B.n1005 B.n72 540.549
R586 B.n569 B.n218 540.549
R587 B.n144 B.n70 540.549
R588 B.n259 B.t13 461.269
R589 B.n111 B.t8 461.269
R590 B.n253 B.t19 461.269
R591 B.n105 B.t15 461.269
R592 B.n259 B.t10 418.368
R593 B.n253 B.t17 418.368
R594 B.n105 B.t14 418.368
R595 B.n111 B.t6 418.368
R596 B.n260 B.t12 411.62
R597 B.n112 B.t9 411.62
R598 B.n254 B.t18 411.62
R599 B.n106 B.t16 411.62
R600 B.n732 B.n71 256.663
R601 B.n734 B.n71 256.663
R602 B.n740 B.n71 256.663
R603 B.n742 B.n71 256.663
R604 B.n748 B.n71 256.663
R605 B.n750 B.n71 256.663
R606 B.n756 B.n71 256.663
R607 B.n758 B.n71 256.663
R608 B.n764 B.n71 256.663
R609 B.n766 B.n71 256.663
R610 B.n772 B.n71 256.663
R611 B.n774 B.n71 256.663
R612 B.n780 B.n71 256.663
R613 B.n782 B.n71 256.663
R614 B.n788 B.n71 256.663
R615 B.n790 B.n71 256.663
R616 B.n796 B.n71 256.663
R617 B.n798 B.n71 256.663
R618 B.n804 B.n71 256.663
R619 B.n806 B.n71 256.663
R620 B.n812 B.n71 256.663
R621 B.n814 B.n71 256.663
R622 B.n820 B.n71 256.663
R623 B.n822 B.n71 256.663
R624 B.n828 B.n71 256.663
R625 B.n830 B.n71 256.663
R626 B.n836 B.n71 256.663
R627 B.n838 B.n71 256.663
R628 B.n844 B.n71 256.663
R629 B.n846 B.n71 256.663
R630 B.n852 B.n71 256.663
R631 B.n854 B.n71 256.663
R632 B.n861 B.n71 256.663
R633 B.n863 B.n71 256.663
R634 B.n869 B.n71 256.663
R635 B.n871 B.n71 256.663
R636 B.n878 B.n71 256.663
R637 B.n880 B.n71 256.663
R638 B.n886 B.n71 256.663
R639 B.n888 B.n71 256.663
R640 B.n894 B.n71 256.663
R641 B.n896 B.n71 256.663
R642 B.n902 B.n71 256.663
R643 B.n904 B.n71 256.663
R644 B.n910 B.n71 256.663
R645 B.n912 B.n71 256.663
R646 B.n918 B.n71 256.663
R647 B.n920 B.n71 256.663
R648 B.n926 B.n71 256.663
R649 B.n928 B.n71 256.663
R650 B.n934 B.n71 256.663
R651 B.n936 B.n71 256.663
R652 B.n942 B.n71 256.663
R653 B.n944 B.n71 256.663
R654 B.n950 B.n71 256.663
R655 B.n952 B.n71 256.663
R656 B.n958 B.n71 256.663
R657 B.n960 B.n71 256.663
R658 B.n966 B.n71 256.663
R659 B.n968 B.n71 256.663
R660 B.n974 B.n71 256.663
R661 B.n976 B.n71 256.663
R662 B.n982 B.n71 256.663
R663 B.n984 B.n71 256.663
R664 B.n990 B.n71 256.663
R665 B.n992 B.n71 256.663
R666 B.n998 B.n71 256.663
R667 B.n1000 B.n71 256.663
R668 B.n562 B.n219 256.663
R669 B.n222 B.n219 256.663
R670 B.n555 B.n219 256.663
R671 B.n549 B.n219 256.663
R672 B.n547 B.n219 256.663
R673 B.n541 B.n219 256.663
R674 B.n539 B.n219 256.663
R675 B.n533 B.n219 256.663
R676 B.n531 B.n219 256.663
R677 B.n525 B.n219 256.663
R678 B.n523 B.n219 256.663
R679 B.n517 B.n219 256.663
R680 B.n515 B.n219 256.663
R681 B.n509 B.n219 256.663
R682 B.n507 B.n219 256.663
R683 B.n501 B.n219 256.663
R684 B.n499 B.n219 256.663
R685 B.n493 B.n219 256.663
R686 B.n491 B.n219 256.663
R687 B.n485 B.n219 256.663
R688 B.n483 B.n219 256.663
R689 B.n477 B.n219 256.663
R690 B.n475 B.n219 256.663
R691 B.n469 B.n219 256.663
R692 B.n467 B.n219 256.663
R693 B.n461 B.n219 256.663
R694 B.n459 B.n219 256.663
R695 B.n453 B.n219 256.663
R696 B.n451 B.n219 256.663
R697 B.n445 B.n219 256.663
R698 B.n443 B.n219 256.663
R699 B.n436 B.n219 256.663
R700 B.n434 B.n219 256.663
R701 B.n428 B.n219 256.663
R702 B.n426 B.n219 256.663
R703 B.n420 B.n219 256.663
R704 B.n262 B.n219 256.663
R705 B.n414 B.n219 256.663
R706 B.n408 B.n219 256.663
R707 B.n406 B.n219 256.663
R708 B.n400 B.n219 256.663
R709 B.n398 B.n219 256.663
R710 B.n392 B.n219 256.663
R711 B.n390 B.n219 256.663
R712 B.n384 B.n219 256.663
R713 B.n382 B.n219 256.663
R714 B.n376 B.n219 256.663
R715 B.n374 B.n219 256.663
R716 B.n368 B.n219 256.663
R717 B.n366 B.n219 256.663
R718 B.n360 B.n219 256.663
R719 B.n358 B.n219 256.663
R720 B.n352 B.n219 256.663
R721 B.n350 B.n219 256.663
R722 B.n344 B.n219 256.663
R723 B.n342 B.n219 256.663
R724 B.n336 B.n219 256.663
R725 B.n334 B.n219 256.663
R726 B.n328 B.n219 256.663
R727 B.n326 B.n219 256.663
R728 B.n320 B.n219 256.663
R729 B.n318 B.n219 256.663
R730 B.n312 B.n219 256.663
R731 B.n310 B.n219 256.663
R732 B.n304 B.n219 256.663
R733 B.n302 B.n219 256.663
R734 B.n296 B.n219 256.663
R735 B.n294 B.n219 256.663
R736 B.n567 B.n214 163.367
R737 B.n575 B.n214 163.367
R738 B.n575 B.n212 163.367
R739 B.n579 B.n212 163.367
R740 B.n579 B.n206 163.367
R741 B.n587 B.n206 163.367
R742 B.n587 B.n204 163.367
R743 B.n591 B.n204 163.367
R744 B.n591 B.n198 163.367
R745 B.n599 B.n198 163.367
R746 B.n599 B.n196 163.367
R747 B.n603 B.n196 163.367
R748 B.n603 B.n190 163.367
R749 B.n611 B.n190 163.367
R750 B.n611 B.n188 163.367
R751 B.n615 B.n188 163.367
R752 B.n615 B.n182 163.367
R753 B.n623 B.n182 163.367
R754 B.n623 B.n180 163.367
R755 B.n627 B.n180 163.367
R756 B.n627 B.n174 163.367
R757 B.n635 B.n174 163.367
R758 B.n635 B.n172 163.367
R759 B.n639 B.n172 163.367
R760 B.n639 B.n166 163.367
R761 B.n647 B.n166 163.367
R762 B.n647 B.n164 163.367
R763 B.n651 B.n164 163.367
R764 B.n651 B.n158 163.367
R765 B.n659 B.n158 163.367
R766 B.n659 B.n156 163.367
R767 B.n663 B.n156 163.367
R768 B.n663 B.n150 163.367
R769 B.n672 B.n150 163.367
R770 B.n672 B.n148 163.367
R771 B.n676 B.n148 163.367
R772 B.n676 B.n2 163.367
R773 B.n1081 B.n2 163.367
R774 B.n1081 B.n3 163.367
R775 B.n1077 B.n3 163.367
R776 B.n1077 B.n9 163.367
R777 B.n1073 B.n9 163.367
R778 B.n1073 B.n11 163.367
R779 B.n1069 B.n11 163.367
R780 B.n1069 B.n16 163.367
R781 B.n1065 B.n16 163.367
R782 B.n1065 B.n18 163.367
R783 B.n1061 B.n18 163.367
R784 B.n1061 B.n23 163.367
R785 B.n1057 B.n23 163.367
R786 B.n1057 B.n25 163.367
R787 B.n1053 B.n25 163.367
R788 B.n1053 B.n30 163.367
R789 B.n1049 B.n30 163.367
R790 B.n1049 B.n32 163.367
R791 B.n1045 B.n32 163.367
R792 B.n1045 B.n37 163.367
R793 B.n1041 B.n37 163.367
R794 B.n1041 B.n39 163.367
R795 B.n1037 B.n39 163.367
R796 B.n1037 B.n44 163.367
R797 B.n1033 B.n44 163.367
R798 B.n1033 B.n46 163.367
R799 B.n1029 B.n46 163.367
R800 B.n1029 B.n51 163.367
R801 B.n1025 B.n51 163.367
R802 B.n1025 B.n53 163.367
R803 B.n1021 B.n53 163.367
R804 B.n1021 B.n58 163.367
R805 B.n1017 B.n58 163.367
R806 B.n1017 B.n60 163.367
R807 B.n1013 B.n60 163.367
R808 B.n1013 B.n65 163.367
R809 B.n1009 B.n65 163.367
R810 B.n1009 B.n67 163.367
R811 B.n1005 B.n67 163.367
R812 B.n563 B.n561 163.367
R813 B.n561 B.n560 163.367
R814 B.n557 B.n556 163.367
R815 B.n554 B.n224 163.367
R816 B.n550 B.n548 163.367
R817 B.n546 B.n226 163.367
R818 B.n542 B.n540 163.367
R819 B.n538 B.n228 163.367
R820 B.n534 B.n532 163.367
R821 B.n530 B.n230 163.367
R822 B.n526 B.n524 163.367
R823 B.n522 B.n232 163.367
R824 B.n518 B.n516 163.367
R825 B.n514 B.n234 163.367
R826 B.n510 B.n508 163.367
R827 B.n506 B.n236 163.367
R828 B.n502 B.n500 163.367
R829 B.n498 B.n238 163.367
R830 B.n494 B.n492 163.367
R831 B.n490 B.n240 163.367
R832 B.n486 B.n484 163.367
R833 B.n482 B.n242 163.367
R834 B.n478 B.n476 163.367
R835 B.n474 B.n244 163.367
R836 B.n470 B.n468 163.367
R837 B.n466 B.n246 163.367
R838 B.n462 B.n460 163.367
R839 B.n458 B.n248 163.367
R840 B.n454 B.n452 163.367
R841 B.n450 B.n250 163.367
R842 B.n446 B.n444 163.367
R843 B.n442 B.n252 163.367
R844 B.n437 B.n435 163.367
R845 B.n433 B.n256 163.367
R846 B.n429 B.n427 163.367
R847 B.n425 B.n258 163.367
R848 B.n421 B.n419 163.367
R849 B.n416 B.n415 163.367
R850 B.n413 B.n264 163.367
R851 B.n409 B.n407 163.367
R852 B.n405 B.n266 163.367
R853 B.n401 B.n399 163.367
R854 B.n397 B.n268 163.367
R855 B.n393 B.n391 163.367
R856 B.n389 B.n270 163.367
R857 B.n385 B.n383 163.367
R858 B.n381 B.n272 163.367
R859 B.n377 B.n375 163.367
R860 B.n373 B.n274 163.367
R861 B.n369 B.n367 163.367
R862 B.n365 B.n276 163.367
R863 B.n361 B.n359 163.367
R864 B.n357 B.n278 163.367
R865 B.n353 B.n351 163.367
R866 B.n349 B.n280 163.367
R867 B.n345 B.n343 163.367
R868 B.n341 B.n282 163.367
R869 B.n337 B.n335 163.367
R870 B.n333 B.n284 163.367
R871 B.n329 B.n327 163.367
R872 B.n325 B.n286 163.367
R873 B.n321 B.n319 163.367
R874 B.n317 B.n288 163.367
R875 B.n313 B.n311 163.367
R876 B.n309 B.n290 163.367
R877 B.n305 B.n303 163.367
R878 B.n301 B.n292 163.367
R879 B.n297 B.n295 163.367
R880 B.n569 B.n216 163.367
R881 B.n573 B.n216 163.367
R882 B.n573 B.n210 163.367
R883 B.n581 B.n210 163.367
R884 B.n581 B.n208 163.367
R885 B.n585 B.n208 163.367
R886 B.n585 B.n202 163.367
R887 B.n593 B.n202 163.367
R888 B.n593 B.n200 163.367
R889 B.n597 B.n200 163.367
R890 B.n597 B.n194 163.367
R891 B.n605 B.n194 163.367
R892 B.n605 B.n192 163.367
R893 B.n609 B.n192 163.367
R894 B.n609 B.n185 163.367
R895 B.n617 B.n185 163.367
R896 B.n617 B.n183 163.367
R897 B.n621 B.n183 163.367
R898 B.n621 B.n178 163.367
R899 B.n629 B.n178 163.367
R900 B.n629 B.n176 163.367
R901 B.n633 B.n176 163.367
R902 B.n633 B.n169 163.367
R903 B.n641 B.n169 163.367
R904 B.n641 B.n167 163.367
R905 B.n645 B.n167 163.367
R906 B.n645 B.n162 163.367
R907 B.n653 B.n162 163.367
R908 B.n653 B.n160 163.367
R909 B.n657 B.n160 163.367
R910 B.n657 B.n154 163.367
R911 B.n665 B.n154 163.367
R912 B.n665 B.n152 163.367
R913 B.n670 B.n152 163.367
R914 B.n670 B.n146 163.367
R915 B.n678 B.n146 163.367
R916 B.n679 B.n678 163.367
R917 B.n679 B.n5 163.367
R918 B.n6 B.n5 163.367
R919 B.n7 B.n6 163.367
R920 B.n684 B.n7 163.367
R921 B.n684 B.n12 163.367
R922 B.n13 B.n12 163.367
R923 B.n14 B.n13 163.367
R924 B.n689 B.n14 163.367
R925 B.n689 B.n19 163.367
R926 B.n20 B.n19 163.367
R927 B.n21 B.n20 163.367
R928 B.n694 B.n21 163.367
R929 B.n694 B.n26 163.367
R930 B.n27 B.n26 163.367
R931 B.n28 B.n27 163.367
R932 B.n699 B.n28 163.367
R933 B.n699 B.n33 163.367
R934 B.n34 B.n33 163.367
R935 B.n35 B.n34 163.367
R936 B.n704 B.n35 163.367
R937 B.n704 B.n40 163.367
R938 B.n41 B.n40 163.367
R939 B.n42 B.n41 163.367
R940 B.n709 B.n42 163.367
R941 B.n709 B.n47 163.367
R942 B.n48 B.n47 163.367
R943 B.n49 B.n48 163.367
R944 B.n714 B.n49 163.367
R945 B.n714 B.n54 163.367
R946 B.n55 B.n54 163.367
R947 B.n56 B.n55 163.367
R948 B.n719 B.n56 163.367
R949 B.n719 B.n61 163.367
R950 B.n62 B.n61 163.367
R951 B.n63 B.n62 163.367
R952 B.n724 B.n63 163.367
R953 B.n724 B.n68 163.367
R954 B.n69 B.n68 163.367
R955 B.n70 B.n69 163.367
R956 B.n1001 B.n999 163.367
R957 B.n997 B.n74 163.367
R958 B.n993 B.n991 163.367
R959 B.n989 B.n76 163.367
R960 B.n985 B.n983 163.367
R961 B.n981 B.n78 163.367
R962 B.n977 B.n975 163.367
R963 B.n973 B.n80 163.367
R964 B.n969 B.n967 163.367
R965 B.n965 B.n82 163.367
R966 B.n961 B.n959 163.367
R967 B.n957 B.n84 163.367
R968 B.n953 B.n951 163.367
R969 B.n949 B.n86 163.367
R970 B.n945 B.n943 163.367
R971 B.n941 B.n88 163.367
R972 B.n937 B.n935 163.367
R973 B.n933 B.n90 163.367
R974 B.n929 B.n927 163.367
R975 B.n925 B.n92 163.367
R976 B.n921 B.n919 163.367
R977 B.n917 B.n94 163.367
R978 B.n913 B.n911 163.367
R979 B.n909 B.n96 163.367
R980 B.n905 B.n903 163.367
R981 B.n901 B.n98 163.367
R982 B.n897 B.n895 163.367
R983 B.n893 B.n100 163.367
R984 B.n889 B.n887 163.367
R985 B.n885 B.n102 163.367
R986 B.n881 B.n879 163.367
R987 B.n877 B.n104 163.367
R988 B.n872 B.n870 163.367
R989 B.n868 B.n108 163.367
R990 B.n864 B.n862 163.367
R991 B.n860 B.n110 163.367
R992 B.n855 B.n853 163.367
R993 B.n851 B.n114 163.367
R994 B.n847 B.n845 163.367
R995 B.n843 B.n116 163.367
R996 B.n839 B.n837 163.367
R997 B.n835 B.n118 163.367
R998 B.n831 B.n829 163.367
R999 B.n827 B.n120 163.367
R1000 B.n823 B.n821 163.367
R1001 B.n819 B.n122 163.367
R1002 B.n815 B.n813 163.367
R1003 B.n811 B.n124 163.367
R1004 B.n807 B.n805 163.367
R1005 B.n803 B.n126 163.367
R1006 B.n799 B.n797 163.367
R1007 B.n795 B.n128 163.367
R1008 B.n791 B.n789 163.367
R1009 B.n787 B.n130 163.367
R1010 B.n783 B.n781 163.367
R1011 B.n779 B.n132 163.367
R1012 B.n775 B.n773 163.367
R1013 B.n771 B.n134 163.367
R1014 B.n767 B.n765 163.367
R1015 B.n763 B.n136 163.367
R1016 B.n759 B.n757 163.367
R1017 B.n755 B.n138 163.367
R1018 B.n751 B.n749 163.367
R1019 B.n747 B.n140 163.367
R1020 B.n743 B.n741 163.367
R1021 B.n739 B.n142 163.367
R1022 B.n735 B.n733 163.367
R1023 B.n731 B.n144 163.367
R1024 B.n562 B.n220 71.676
R1025 B.n560 B.n222 71.676
R1026 B.n556 B.n555 71.676
R1027 B.n549 B.n224 71.676
R1028 B.n548 B.n547 71.676
R1029 B.n541 B.n226 71.676
R1030 B.n540 B.n539 71.676
R1031 B.n533 B.n228 71.676
R1032 B.n532 B.n531 71.676
R1033 B.n525 B.n230 71.676
R1034 B.n524 B.n523 71.676
R1035 B.n517 B.n232 71.676
R1036 B.n516 B.n515 71.676
R1037 B.n509 B.n234 71.676
R1038 B.n508 B.n507 71.676
R1039 B.n501 B.n236 71.676
R1040 B.n500 B.n499 71.676
R1041 B.n493 B.n238 71.676
R1042 B.n492 B.n491 71.676
R1043 B.n485 B.n240 71.676
R1044 B.n484 B.n483 71.676
R1045 B.n477 B.n242 71.676
R1046 B.n476 B.n475 71.676
R1047 B.n469 B.n244 71.676
R1048 B.n468 B.n467 71.676
R1049 B.n461 B.n246 71.676
R1050 B.n460 B.n459 71.676
R1051 B.n453 B.n248 71.676
R1052 B.n452 B.n451 71.676
R1053 B.n445 B.n250 71.676
R1054 B.n444 B.n443 71.676
R1055 B.n436 B.n252 71.676
R1056 B.n435 B.n434 71.676
R1057 B.n428 B.n256 71.676
R1058 B.n427 B.n426 71.676
R1059 B.n420 B.n258 71.676
R1060 B.n419 B.n262 71.676
R1061 B.n415 B.n414 71.676
R1062 B.n408 B.n264 71.676
R1063 B.n407 B.n406 71.676
R1064 B.n400 B.n266 71.676
R1065 B.n399 B.n398 71.676
R1066 B.n392 B.n268 71.676
R1067 B.n391 B.n390 71.676
R1068 B.n384 B.n270 71.676
R1069 B.n383 B.n382 71.676
R1070 B.n376 B.n272 71.676
R1071 B.n375 B.n374 71.676
R1072 B.n368 B.n274 71.676
R1073 B.n367 B.n366 71.676
R1074 B.n360 B.n276 71.676
R1075 B.n359 B.n358 71.676
R1076 B.n352 B.n278 71.676
R1077 B.n351 B.n350 71.676
R1078 B.n344 B.n280 71.676
R1079 B.n343 B.n342 71.676
R1080 B.n336 B.n282 71.676
R1081 B.n335 B.n334 71.676
R1082 B.n328 B.n284 71.676
R1083 B.n327 B.n326 71.676
R1084 B.n320 B.n286 71.676
R1085 B.n319 B.n318 71.676
R1086 B.n312 B.n288 71.676
R1087 B.n311 B.n310 71.676
R1088 B.n304 B.n290 71.676
R1089 B.n303 B.n302 71.676
R1090 B.n296 B.n292 71.676
R1091 B.n295 B.n294 71.676
R1092 B.n1000 B.n72 71.676
R1093 B.n999 B.n998 71.676
R1094 B.n992 B.n74 71.676
R1095 B.n991 B.n990 71.676
R1096 B.n984 B.n76 71.676
R1097 B.n983 B.n982 71.676
R1098 B.n976 B.n78 71.676
R1099 B.n975 B.n974 71.676
R1100 B.n968 B.n80 71.676
R1101 B.n967 B.n966 71.676
R1102 B.n960 B.n82 71.676
R1103 B.n959 B.n958 71.676
R1104 B.n952 B.n84 71.676
R1105 B.n951 B.n950 71.676
R1106 B.n944 B.n86 71.676
R1107 B.n943 B.n942 71.676
R1108 B.n936 B.n88 71.676
R1109 B.n935 B.n934 71.676
R1110 B.n928 B.n90 71.676
R1111 B.n927 B.n926 71.676
R1112 B.n920 B.n92 71.676
R1113 B.n919 B.n918 71.676
R1114 B.n912 B.n94 71.676
R1115 B.n911 B.n910 71.676
R1116 B.n904 B.n96 71.676
R1117 B.n903 B.n902 71.676
R1118 B.n896 B.n98 71.676
R1119 B.n895 B.n894 71.676
R1120 B.n888 B.n100 71.676
R1121 B.n887 B.n886 71.676
R1122 B.n880 B.n102 71.676
R1123 B.n879 B.n878 71.676
R1124 B.n871 B.n104 71.676
R1125 B.n870 B.n869 71.676
R1126 B.n863 B.n108 71.676
R1127 B.n862 B.n861 71.676
R1128 B.n854 B.n110 71.676
R1129 B.n853 B.n852 71.676
R1130 B.n846 B.n114 71.676
R1131 B.n845 B.n844 71.676
R1132 B.n838 B.n116 71.676
R1133 B.n837 B.n836 71.676
R1134 B.n830 B.n118 71.676
R1135 B.n829 B.n828 71.676
R1136 B.n822 B.n120 71.676
R1137 B.n821 B.n820 71.676
R1138 B.n814 B.n122 71.676
R1139 B.n813 B.n812 71.676
R1140 B.n806 B.n124 71.676
R1141 B.n805 B.n804 71.676
R1142 B.n798 B.n126 71.676
R1143 B.n797 B.n796 71.676
R1144 B.n790 B.n128 71.676
R1145 B.n789 B.n788 71.676
R1146 B.n782 B.n130 71.676
R1147 B.n781 B.n780 71.676
R1148 B.n774 B.n132 71.676
R1149 B.n773 B.n772 71.676
R1150 B.n766 B.n134 71.676
R1151 B.n765 B.n764 71.676
R1152 B.n758 B.n136 71.676
R1153 B.n757 B.n756 71.676
R1154 B.n750 B.n138 71.676
R1155 B.n749 B.n748 71.676
R1156 B.n742 B.n140 71.676
R1157 B.n741 B.n740 71.676
R1158 B.n734 B.n142 71.676
R1159 B.n733 B.n732 71.676
R1160 B.n732 B.n731 71.676
R1161 B.n735 B.n734 71.676
R1162 B.n740 B.n739 71.676
R1163 B.n743 B.n742 71.676
R1164 B.n748 B.n747 71.676
R1165 B.n751 B.n750 71.676
R1166 B.n756 B.n755 71.676
R1167 B.n759 B.n758 71.676
R1168 B.n764 B.n763 71.676
R1169 B.n767 B.n766 71.676
R1170 B.n772 B.n771 71.676
R1171 B.n775 B.n774 71.676
R1172 B.n780 B.n779 71.676
R1173 B.n783 B.n782 71.676
R1174 B.n788 B.n787 71.676
R1175 B.n791 B.n790 71.676
R1176 B.n796 B.n795 71.676
R1177 B.n799 B.n798 71.676
R1178 B.n804 B.n803 71.676
R1179 B.n807 B.n806 71.676
R1180 B.n812 B.n811 71.676
R1181 B.n815 B.n814 71.676
R1182 B.n820 B.n819 71.676
R1183 B.n823 B.n822 71.676
R1184 B.n828 B.n827 71.676
R1185 B.n831 B.n830 71.676
R1186 B.n836 B.n835 71.676
R1187 B.n839 B.n838 71.676
R1188 B.n844 B.n843 71.676
R1189 B.n847 B.n846 71.676
R1190 B.n852 B.n851 71.676
R1191 B.n855 B.n854 71.676
R1192 B.n861 B.n860 71.676
R1193 B.n864 B.n863 71.676
R1194 B.n869 B.n868 71.676
R1195 B.n872 B.n871 71.676
R1196 B.n878 B.n877 71.676
R1197 B.n881 B.n880 71.676
R1198 B.n886 B.n885 71.676
R1199 B.n889 B.n888 71.676
R1200 B.n894 B.n893 71.676
R1201 B.n897 B.n896 71.676
R1202 B.n902 B.n901 71.676
R1203 B.n905 B.n904 71.676
R1204 B.n910 B.n909 71.676
R1205 B.n913 B.n912 71.676
R1206 B.n918 B.n917 71.676
R1207 B.n921 B.n920 71.676
R1208 B.n926 B.n925 71.676
R1209 B.n929 B.n928 71.676
R1210 B.n934 B.n933 71.676
R1211 B.n937 B.n936 71.676
R1212 B.n942 B.n941 71.676
R1213 B.n945 B.n944 71.676
R1214 B.n950 B.n949 71.676
R1215 B.n953 B.n952 71.676
R1216 B.n958 B.n957 71.676
R1217 B.n961 B.n960 71.676
R1218 B.n966 B.n965 71.676
R1219 B.n969 B.n968 71.676
R1220 B.n974 B.n973 71.676
R1221 B.n977 B.n976 71.676
R1222 B.n982 B.n981 71.676
R1223 B.n985 B.n984 71.676
R1224 B.n990 B.n989 71.676
R1225 B.n993 B.n992 71.676
R1226 B.n998 B.n997 71.676
R1227 B.n1001 B.n1000 71.676
R1228 B.n563 B.n562 71.676
R1229 B.n557 B.n222 71.676
R1230 B.n555 B.n554 71.676
R1231 B.n550 B.n549 71.676
R1232 B.n547 B.n546 71.676
R1233 B.n542 B.n541 71.676
R1234 B.n539 B.n538 71.676
R1235 B.n534 B.n533 71.676
R1236 B.n531 B.n530 71.676
R1237 B.n526 B.n525 71.676
R1238 B.n523 B.n522 71.676
R1239 B.n518 B.n517 71.676
R1240 B.n515 B.n514 71.676
R1241 B.n510 B.n509 71.676
R1242 B.n507 B.n506 71.676
R1243 B.n502 B.n501 71.676
R1244 B.n499 B.n498 71.676
R1245 B.n494 B.n493 71.676
R1246 B.n491 B.n490 71.676
R1247 B.n486 B.n485 71.676
R1248 B.n483 B.n482 71.676
R1249 B.n478 B.n477 71.676
R1250 B.n475 B.n474 71.676
R1251 B.n470 B.n469 71.676
R1252 B.n467 B.n466 71.676
R1253 B.n462 B.n461 71.676
R1254 B.n459 B.n458 71.676
R1255 B.n454 B.n453 71.676
R1256 B.n451 B.n450 71.676
R1257 B.n446 B.n445 71.676
R1258 B.n443 B.n442 71.676
R1259 B.n437 B.n436 71.676
R1260 B.n434 B.n433 71.676
R1261 B.n429 B.n428 71.676
R1262 B.n426 B.n425 71.676
R1263 B.n421 B.n420 71.676
R1264 B.n416 B.n262 71.676
R1265 B.n414 B.n413 71.676
R1266 B.n409 B.n408 71.676
R1267 B.n406 B.n405 71.676
R1268 B.n401 B.n400 71.676
R1269 B.n398 B.n397 71.676
R1270 B.n393 B.n392 71.676
R1271 B.n390 B.n389 71.676
R1272 B.n385 B.n384 71.676
R1273 B.n382 B.n381 71.676
R1274 B.n377 B.n376 71.676
R1275 B.n374 B.n373 71.676
R1276 B.n369 B.n368 71.676
R1277 B.n366 B.n365 71.676
R1278 B.n361 B.n360 71.676
R1279 B.n358 B.n357 71.676
R1280 B.n353 B.n352 71.676
R1281 B.n350 B.n349 71.676
R1282 B.n345 B.n344 71.676
R1283 B.n342 B.n341 71.676
R1284 B.n337 B.n336 71.676
R1285 B.n334 B.n333 71.676
R1286 B.n329 B.n328 71.676
R1287 B.n326 B.n325 71.676
R1288 B.n321 B.n320 71.676
R1289 B.n318 B.n317 71.676
R1290 B.n313 B.n312 71.676
R1291 B.n310 B.n309 71.676
R1292 B.n305 B.n304 71.676
R1293 B.n302 B.n301 71.676
R1294 B.n297 B.n296 71.676
R1295 B.n294 B.n218 71.676
R1296 B.n568 B.n219 61.6662
R1297 B.n1006 B.n71 61.6662
R1298 B.n261 B.n260 59.5399
R1299 B.n439 B.n254 59.5399
R1300 B.n875 B.n106 59.5399
R1301 B.n857 B.n112 59.5399
R1302 B.n260 B.n259 49.649
R1303 B.n254 B.n253 49.649
R1304 B.n106 B.n105 49.649
R1305 B.n112 B.n111 49.649
R1306 B.n1004 B.n1003 35.1225
R1307 B.n729 B.n728 35.1225
R1308 B.n570 B.n217 35.1225
R1309 B.n566 B.n565 35.1225
R1310 B.n568 B.n215 30.1679
R1311 B.n574 B.n215 30.1679
R1312 B.n574 B.n211 30.1679
R1313 B.n580 B.n211 30.1679
R1314 B.n580 B.n207 30.1679
R1315 B.n586 B.n207 30.1679
R1316 B.n592 B.n203 30.1679
R1317 B.n592 B.n199 30.1679
R1318 B.n598 B.n199 30.1679
R1319 B.n598 B.n195 30.1679
R1320 B.n604 B.n195 30.1679
R1321 B.n604 B.n191 30.1679
R1322 B.n610 B.n191 30.1679
R1323 B.n610 B.n186 30.1679
R1324 B.n616 B.n186 30.1679
R1325 B.n616 B.n187 30.1679
R1326 B.n622 B.n179 30.1679
R1327 B.n628 B.n179 30.1679
R1328 B.n628 B.n175 30.1679
R1329 B.n634 B.n175 30.1679
R1330 B.n634 B.n170 30.1679
R1331 B.n640 B.n170 30.1679
R1332 B.n640 B.n171 30.1679
R1333 B.n646 B.n163 30.1679
R1334 B.n652 B.n163 30.1679
R1335 B.n652 B.n159 30.1679
R1336 B.n658 B.n159 30.1679
R1337 B.n658 B.n155 30.1679
R1338 B.n664 B.n155 30.1679
R1339 B.n671 B.n151 30.1679
R1340 B.n671 B.n147 30.1679
R1341 B.n677 B.n147 30.1679
R1342 B.n677 B.n4 30.1679
R1343 B.n1080 B.n4 30.1679
R1344 B.n1080 B.n1079 30.1679
R1345 B.n1079 B.n1078 30.1679
R1346 B.n1078 B.n8 30.1679
R1347 B.n1072 B.n8 30.1679
R1348 B.n1072 B.n1071 30.1679
R1349 B.n1070 B.n15 30.1679
R1350 B.n1064 B.n15 30.1679
R1351 B.n1064 B.n1063 30.1679
R1352 B.n1063 B.n1062 30.1679
R1353 B.n1062 B.n22 30.1679
R1354 B.n1056 B.n22 30.1679
R1355 B.n1055 B.n1054 30.1679
R1356 B.n1054 B.n29 30.1679
R1357 B.n1048 B.n29 30.1679
R1358 B.n1048 B.n1047 30.1679
R1359 B.n1047 B.n1046 30.1679
R1360 B.n1046 B.n36 30.1679
R1361 B.n1040 B.n36 30.1679
R1362 B.n1039 B.n1038 30.1679
R1363 B.n1038 B.n43 30.1679
R1364 B.n1032 B.n43 30.1679
R1365 B.n1032 B.n1031 30.1679
R1366 B.n1031 B.n1030 30.1679
R1367 B.n1030 B.n50 30.1679
R1368 B.n1024 B.n50 30.1679
R1369 B.n1024 B.n1023 30.1679
R1370 B.n1023 B.n1022 30.1679
R1371 B.n1022 B.n57 30.1679
R1372 B.n1016 B.n1015 30.1679
R1373 B.n1015 B.n1014 30.1679
R1374 B.n1014 B.n64 30.1679
R1375 B.n1008 B.n64 30.1679
R1376 B.n1008 B.n1007 30.1679
R1377 B.n1007 B.n1006 30.1679
R1378 B.n646 B.t0 27.0624
R1379 B.n1056 B.t4 27.0624
R1380 B.n586 B.t11 25.2879
R1381 B.n1016 B.t7 25.2879
R1382 B.n664 B.t1 19.0769
R1383 B.t2 B.n1070 19.0769
R1384 B B.n1082 18.0485
R1385 B.n187 B.t5 17.3024
R1386 B.t3 B.n1039 17.3024
R1387 B.n622 B.t5 12.866
R1388 B.n1040 B.t3 12.866
R1389 B.t1 B.n151 11.0914
R1390 B.n1071 B.t2 11.0914
R1391 B.n1003 B.n1002 10.6151
R1392 B.n1002 B.n73 10.6151
R1393 B.n996 B.n73 10.6151
R1394 B.n996 B.n995 10.6151
R1395 B.n995 B.n994 10.6151
R1396 B.n994 B.n75 10.6151
R1397 B.n988 B.n75 10.6151
R1398 B.n988 B.n987 10.6151
R1399 B.n987 B.n986 10.6151
R1400 B.n986 B.n77 10.6151
R1401 B.n980 B.n77 10.6151
R1402 B.n980 B.n979 10.6151
R1403 B.n979 B.n978 10.6151
R1404 B.n978 B.n79 10.6151
R1405 B.n972 B.n79 10.6151
R1406 B.n972 B.n971 10.6151
R1407 B.n971 B.n970 10.6151
R1408 B.n970 B.n81 10.6151
R1409 B.n964 B.n81 10.6151
R1410 B.n964 B.n963 10.6151
R1411 B.n963 B.n962 10.6151
R1412 B.n962 B.n83 10.6151
R1413 B.n956 B.n83 10.6151
R1414 B.n956 B.n955 10.6151
R1415 B.n955 B.n954 10.6151
R1416 B.n954 B.n85 10.6151
R1417 B.n948 B.n85 10.6151
R1418 B.n948 B.n947 10.6151
R1419 B.n947 B.n946 10.6151
R1420 B.n946 B.n87 10.6151
R1421 B.n940 B.n87 10.6151
R1422 B.n940 B.n939 10.6151
R1423 B.n939 B.n938 10.6151
R1424 B.n938 B.n89 10.6151
R1425 B.n932 B.n89 10.6151
R1426 B.n932 B.n931 10.6151
R1427 B.n931 B.n930 10.6151
R1428 B.n930 B.n91 10.6151
R1429 B.n924 B.n91 10.6151
R1430 B.n924 B.n923 10.6151
R1431 B.n923 B.n922 10.6151
R1432 B.n922 B.n93 10.6151
R1433 B.n916 B.n93 10.6151
R1434 B.n916 B.n915 10.6151
R1435 B.n915 B.n914 10.6151
R1436 B.n914 B.n95 10.6151
R1437 B.n908 B.n95 10.6151
R1438 B.n908 B.n907 10.6151
R1439 B.n907 B.n906 10.6151
R1440 B.n906 B.n97 10.6151
R1441 B.n900 B.n97 10.6151
R1442 B.n900 B.n899 10.6151
R1443 B.n899 B.n898 10.6151
R1444 B.n898 B.n99 10.6151
R1445 B.n892 B.n99 10.6151
R1446 B.n892 B.n891 10.6151
R1447 B.n891 B.n890 10.6151
R1448 B.n890 B.n101 10.6151
R1449 B.n884 B.n101 10.6151
R1450 B.n884 B.n883 10.6151
R1451 B.n883 B.n882 10.6151
R1452 B.n882 B.n103 10.6151
R1453 B.n876 B.n103 10.6151
R1454 B.n874 B.n873 10.6151
R1455 B.n873 B.n107 10.6151
R1456 B.n867 B.n107 10.6151
R1457 B.n867 B.n866 10.6151
R1458 B.n866 B.n865 10.6151
R1459 B.n865 B.n109 10.6151
R1460 B.n859 B.n109 10.6151
R1461 B.n859 B.n858 10.6151
R1462 B.n856 B.n113 10.6151
R1463 B.n850 B.n113 10.6151
R1464 B.n850 B.n849 10.6151
R1465 B.n849 B.n848 10.6151
R1466 B.n848 B.n115 10.6151
R1467 B.n842 B.n115 10.6151
R1468 B.n842 B.n841 10.6151
R1469 B.n841 B.n840 10.6151
R1470 B.n840 B.n117 10.6151
R1471 B.n834 B.n117 10.6151
R1472 B.n834 B.n833 10.6151
R1473 B.n833 B.n832 10.6151
R1474 B.n832 B.n119 10.6151
R1475 B.n826 B.n119 10.6151
R1476 B.n826 B.n825 10.6151
R1477 B.n825 B.n824 10.6151
R1478 B.n824 B.n121 10.6151
R1479 B.n818 B.n121 10.6151
R1480 B.n818 B.n817 10.6151
R1481 B.n817 B.n816 10.6151
R1482 B.n816 B.n123 10.6151
R1483 B.n810 B.n123 10.6151
R1484 B.n810 B.n809 10.6151
R1485 B.n809 B.n808 10.6151
R1486 B.n808 B.n125 10.6151
R1487 B.n802 B.n125 10.6151
R1488 B.n802 B.n801 10.6151
R1489 B.n801 B.n800 10.6151
R1490 B.n800 B.n127 10.6151
R1491 B.n794 B.n127 10.6151
R1492 B.n794 B.n793 10.6151
R1493 B.n793 B.n792 10.6151
R1494 B.n792 B.n129 10.6151
R1495 B.n786 B.n129 10.6151
R1496 B.n786 B.n785 10.6151
R1497 B.n785 B.n784 10.6151
R1498 B.n784 B.n131 10.6151
R1499 B.n778 B.n131 10.6151
R1500 B.n778 B.n777 10.6151
R1501 B.n777 B.n776 10.6151
R1502 B.n776 B.n133 10.6151
R1503 B.n770 B.n133 10.6151
R1504 B.n770 B.n769 10.6151
R1505 B.n769 B.n768 10.6151
R1506 B.n768 B.n135 10.6151
R1507 B.n762 B.n135 10.6151
R1508 B.n762 B.n761 10.6151
R1509 B.n761 B.n760 10.6151
R1510 B.n760 B.n137 10.6151
R1511 B.n754 B.n137 10.6151
R1512 B.n754 B.n753 10.6151
R1513 B.n753 B.n752 10.6151
R1514 B.n752 B.n139 10.6151
R1515 B.n746 B.n139 10.6151
R1516 B.n746 B.n745 10.6151
R1517 B.n745 B.n744 10.6151
R1518 B.n744 B.n141 10.6151
R1519 B.n738 B.n141 10.6151
R1520 B.n738 B.n737 10.6151
R1521 B.n737 B.n736 10.6151
R1522 B.n736 B.n143 10.6151
R1523 B.n730 B.n143 10.6151
R1524 B.n730 B.n729 10.6151
R1525 B.n571 B.n570 10.6151
R1526 B.n572 B.n571 10.6151
R1527 B.n572 B.n209 10.6151
R1528 B.n582 B.n209 10.6151
R1529 B.n583 B.n582 10.6151
R1530 B.n584 B.n583 10.6151
R1531 B.n584 B.n201 10.6151
R1532 B.n594 B.n201 10.6151
R1533 B.n595 B.n594 10.6151
R1534 B.n596 B.n595 10.6151
R1535 B.n596 B.n193 10.6151
R1536 B.n606 B.n193 10.6151
R1537 B.n607 B.n606 10.6151
R1538 B.n608 B.n607 10.6151
R1539 B.n608 B.n184 10.6151
R1540 B.n618 B.n184 10.6151
R1541 B.n619 B.n618 10.6151
R1542 B.n620 B.n619 10.6151
R1543 B.n620 B.n177 10.6151
R1544 B.n630 B.n177 10.6151
R1545 B.n631 B.n630 10.6151
R1546 B.n632 B.n631 10.6151
R1547 B.n632 B.n168 10.6151
R1548 B.n642 B.n168 10.6151
R1549 B.n643 B.n642 10.6151
R1550 B.n644 B.n643 10.6151
R1551 B.n644 B.n161 10.6151
R1552 B.n654 B.n161 10.6151
R1553 B.n655 B.n654 10.6151
R1554 B.n656 B.n655 10.6151
R1555 B.n656 B.n153 10.6151
R1556 B.n666 B.n153 10.6151
R1557 B.n667 B.n666 10.6151
R1558 B.n669 B.n667 10.6151
R1559 B.n669 B.n668 10.6151
R1560 B.n668 B.n145 10.6151
R1561 B.n680 B.n145 10.6151
R1562 B.n681 B.n680 10.6151
R1563 B.n682 B.n681 10.6151
R1564 B.n683 B.n682 10.6151
R1565 B.n685 B.n683 10.6151
R1566 B.n686 B.n685 10.6151
R1567 B.n687 B.n686 10.6151
R1568 B.n688 B.n687 10.6151
R1569 B.n690 B.n688 10.6151
R1570 B.n691 B.n690 10.6151
R1571 B.n692 B.n691 10.6151
R1572 B.n693 B.n692 10.6151
R1573 B.n695 B.n693 10.6151
R1574 B.n696 B.n695 10.6151
R1575 B.n697 B.n696 10.6151
R1576 B.n698 B.n697 10.6151
R1577 B.n700 B.n698 10.6151
R1578 B.n701 B.n700 10.6151
R1579 B.n702 B.n701 10.6151
R1580 B.n703 B.n702 10.6151
R1581 B.n705 B.n703 10.6151
R1582 B.n706 B.n705 10.6151
R1583 B.n707 B.n706 10.6151
R1584 B.n708 B.n707 10.6151
R1585 B.n710 B.n708 10.6151
R1586 B.n711 B.n710 10.6151
R1587 B.n712 B.n711 10.6151
R1588 B.n713 B.n712 10.6151
R1589 B.n715 B.n713 10.6151
R1590 B.n716 B.n715 10.6151
R1591 B.n717 B.n716 10.6151
R1592 B.n718 B.n717 10.6151
R1593 B.n720 B.n718 10.6151
R1594 B.n721 B.n720 10.6151
R1595 B.n722 B.n721 10.6151
R1596 B.n723 B.n722 10.6151
R1597 B.n725 B.n723 10.6151
R1598 B.n726 B.n725 10.6151
R1599 B.n727 B.n726 10.6151
R1600 B.n728 B.n727 10.6151
R1601 B.n565 B.n564 10.6151
R1602 B.n564 B.n221 10.6151
R1603 B.n559 B.n221 10.6151
R1604 B.n559 B.n558 10.6151
R1605 B.n558 B.n223 10.6151
R1606 B.n553 B.n223 10.6151
R1607 B.n553 B.n552 10.6151
R1608 B.n552 B.n551 10.6151
R1609 B.n551 B.n225 10.6151
R1610 B.n545 B.n225 10.6151
R1611 B.n545 B.n544 10.6151
R1612 B.n544 B.n543 10.6151
R1613 B.n543 B.n227 10.6151
R1614 B.n537 B.n227 10.6151
R1615 B.n537 B.n536 10.6151
R1616 B.n536 B.n535 10.6151
R1617 B.n535 B.n229 10.6151
R1618 B.n529 B.n229 10.6151
R1619 B.n529 B.n528 10.6151
R1620 B.n528 B.n527 10.6151
R1621 B.n527 B.n231 10.6151
R1622 B.n521 B.n231 10.6151
R1623 B.n521 B.n520 10.6151
R1624 B.n520 B.n519 10.6151
R1625 B.n519 B.n233 10.6151
R1626 B.n513 B.n233 10.6151
R1627 B.n513 B.n512 10.6151
R1628 B.n512 B.n511 10.6151
R1629 B.n511 B.n235 10.6151
R1630 B.n505 B.n235 10.6151
R1631 B.n505 B.n504 10.6151
R1632 B.n504 B.n503 10.6151
R1633 B.n503 B.n237 10.6151
R1634 B.n497 B.n237 10.6151
R1635 B.n497 B.n496 10.6151
R1636 B.n496 B.n495 10.6151
R1637 B.n495 B.n239 10.6151
R1638 B.n489 B.n239 10.6151
R1639 B.n489 B.n488 10.6151
R1640 B.n488 B.n487 10.6151
R1641 B.n487 B.n241 10.6151
R1642 B.n481 B.n241 10.6151
R1643 B.n481 B.n480 10.6151
R1644 B.n480 B.n479 10.6151
R1645 B.n479 B.n243 10.6151
R1646 B.n473 B.n243 10.6151
R1647 B.n473 B.n472 10.6151
R1648 B.n472 B.n471 10.6151
R1649 B.n471 B.n245 10.6151
R1650 B.n465 B.n245 10.6151
R1651 B.n465 B.n464 10.6151
R1652 B.n464 B.n463 10.6151
R1653 B.n463 B.n247 10.6151
R1654 B.n457 B.n247 10.6151
R1655 B.n457 B.n456 10.6151
R1656 B.n456 B.n455 10.6151
R1657 B.n455 B.n249 10.6151
R1658 B.n449 B.n249 10.6151
R1659 B.n449 B.n448 10.6151
R1660 B.n448 B.n447 10.6151
R1661 B.n447 B.n251 10.6151
R1662 B.n441 B.n251 10.6151
R1663 B.n441 B.n440 10.6151
R1664 B.n438 B.n255 10.6151
R1665 B.n432 B.n255 10.6151
R1666 B.n432 B.n431 10.6151
R1667 B.n431 B.n430 10.6151
R1668 B.n430 B.n257 10.6151
R1669 B.n424 B.n257 10.6151
R1670 B.n424 B.n423 10.6151
R1671 B.n423 B.n422 10.6151
R1672 B.n418 B.n417 10.6151
R1673 B.n417 B.n263 10.6151
R1674 B.n412 B.n263 10.6151
R1675 B.n412 B.n411 10.6151
R1676 B.n411 B.n410 10.6151
R1677 B.n410 B.n265 10.6151
R1678 B.n404 B.n265 10.6151
R1679 B.n404 B.n403 10.6151
R1680 B.n403 B.n402 10.6151
R1681 B.n402 B.n267 10.6151
R1682 B.n396 B.n267 10.6151
R1683 B.n396 B.n395 10.6151
R1684 B.n395 B.n394 10.6151
R1685 B.n394 B.n269 10.6151
R1686 B.n388 B.n269 10.6151
R1687 B.n388 B.n387 10.6151
R1688 B.n387 B.n386 10.6151
R1689 B.n386 B.n271 10.6151
R1690 B.n380 B.n271 10.6151
R1691 B.n380 B.n379 10.6151
R1692 B.n379 B.n378 10.6151
R1693 B.n378 B.n273 10.6151
R1694 B.n372 B.n273 10.6151
R1695 B.n372 B.n371 10.6151
R1696 B.n371 B.n370 10.6151
R1697 B.n370 B.n275 10.6151
R1698 B.n364 B.n275 10.6151
R1699 B.n364 B.n363 10.6151
R1700 B.n363 B.n362 10.6151
R1701 B.n362 B.n277 10.6151
R1702 B.n356 B.n277 10.6151
R1703 B.n356 B.n355 10.6151
R1704 B.n355 B.n354 10.6151
R1705 B.n354 B.n279 10.6151
R1706 B.n348 B.n279 10.6151
R1707 B.n348 B.n347 10.6151
R1708 B.n347 B.n346 10.6151
R1709 B.n346 B.n281 10.6151
R1710 B.n340 B.n281 10.6151
R1711 B.n340 B.n339 10.6151
R1712 B.n339 B.n338 10.6151
R1713 B.n338 B.n283 10.6151
R1714 B.n332 B.n283 10.6151
R1715 B.n332 B.n331 10.6151
R1716 B.n331 B.n330 10.6151
R1717 B.n330 B.n285 10.6151
R1718 B.n324 B.n285 10.6151
R1719 B.n324 B.n323 10.6151
R1720 B.n323 B.n322 10.6151
R1721 B.n322 B.n287 10.6151
R1722 B.n316 B.n287 10.6151
R1723 B.n316 B.n315 10.6151
R1724 B.n315 B.n314 10.6151
R1725 B.n314 B.n289 10.6151
R1726 B.n308 B.n289 10.6151
R1727 B.n308 B.n307 10.6151
R1728 B.n307 B.n306 10.6151
R1729 B.n306 B.n291 10.6151
R1730 B.n300 B.n291 10.6151
R1731 B.n300 B.n299 10.6151
R1732 B.n299 B.n298 10.6151
R1733 B.n298 B.n293 10.6151
R1734 B.n293 B.n217 10.6151
R1735 B.n566 B.n213 10.6151
R1736 B.n576 B.n213 10.6151
R1737 B.n577 B.n576 10.6151
R1738 B.n578 B.n577 10.6151
R1739 B.n578 B.n205 10.6151
R1740 B.n588 B.n205 10.6151
R1741 B.n589 B.n588 10.6151
R1742 B.n590 B.n589 10.6151
R1743 B.n590 B.n197 10.6151
R1744 B.n600 B.n197 10.6151
R1745 B.n601 B.n600 10.6151
R1746 B.n602 B.n601 10.6151
R1747 B.n602 B.n189 10.6151
R1748 B.n612 B.n189 10.6151
R1749 B.n613 B.n612 10.6151
R1750 B.n614 B.n613 10.6151
R1751 B.n614 B.n181 10.6151
R1752 B.n624 B.n181 10.6151
R1753 B.n625 B.n624 10.6151
R1754 B.n626 B.n625 10.6151
R1755 B.n626 B.n173 10.6151
R1756 B.n636 B.n173 10.6151
R1757 B.n637 B.n636 10.6151
R1758 B.n638 B.n637 10.6151
R1759 B.n638 B.n165 10.6151
R1760 B.n648 B.n165 10.6151
R1761 B.n649 B.n648 10.6151
R1762 B.n650 B.n649 10.6151
R1763 B.n650 B.n157 10.6151
R1764 B.n660 B.n157 10.6151
R1765 B.n661 B.n660 10.6151
R1766 B.n662 B.n661 10.6151
R1767 B.n662 B.n149 10.6151
R1768 B.n673 B.n149 10.6151
R1769 B.n674 B.n673 10.6151
R1770 B.n675 B.n674 10.6151
R1771 B.n675 B.n0 10.6151
R1772 B.n1076 B.n1 10.6151
R1773 B.n1076 B.n1075 10.6151
R1774 B.n1075 B.n1074 10.6151
R1775 B.n1074 B.n10 10.6151
R1776 B.n1068 B.n10 10.6151
R1777 B.n1068 B.n1067 10.6151
R1778 B.n1067 B.n1066 10.6151
R1779 B.n1066 B.n17 10.6151
R1780 B.n1060 B.n17 10.6151
R1781 B.n1060 B.n1059 10.6151
R1782 B.n1059 B.n1058 10.6151
R1783 B.n1058 B.n24 10.6151
R1784 B.n1052 B.n24 10.6151
R1785 B.n1052 B.n1051 10.6151
R1786 B.n1051 B.n1050 10.6151
R1787 B.n1050 B.n31 10.6151
R1788 B.n1044 B.n31 10.6151
R1789 B.n1044 B.n1043 10.6151
R1790 B.n1043 B.n1042 10.6151
R1791 B.n1042 B.n38 10.6151
R1792 B.n1036 B.n38 10.6151
R1793 B.n1036 B.n1035 10.6151
R1794 B.n1035 B.n1034 10.6151
R1795 B.n1034 B.n45 10.6151
R1796 B.n1028 B.n45 10.6151
R1797 B.n1028 B.n1027 10.6151
R1798 B.n1027 B.n1026 10.6151
R1799 B.n1026 B.n52 10.6151
R1800 B.n1020 B.n52 10.6151
R1801 B.n1020 B.n1019 10.6151
R1802 B.n1019 B.n1018 10.6151
R1803 B.n1018 B.n59 10.6151
R1804 B.n1012 B.n59 10.6151
R1805 B.n1012 B.n1011 10.6151
R1806 B.n1011 B.n1010 10.6151
R1807 B.n1010 B.n66 10.6151
R1808 B.n1004 B.n66 10.6151
R1809 B.n875 B.n874 6.5566
R1810 B.n858 B.n857 6.5566
R1811 B.n439 B.n438 6.5566
R1812 B.n422 B.n261 6.5566
R1813 B.t11 B.n203 4.88052
R1814 B.t7 B.n57 4.88052
R1815 B.n876 B.n875 4.05904
R1816 B.n857 B.n856 4.05904
R1817 B.n440 B.n439 4.05904
R1818 B.n418 B.n261 4.05904
R1819 B.n171 B.t0 3.10596
R1820 B.t4 B.n1055 3.10596
R1821 B.n1082 B.n0 2.81026
R1822 B.n1082 B.n1 2.81026
R1823 VN.n3 VN.t5 243.868
R1824 VN.n17 VN.t3 243.868
R1825 VN.n4 VN.t2 210.957
R1826 VN.n12 VN.t1 210.957
R1827 VN.n18 VN.t0 210.957
R1828 VN.n26 VN.t4 210.957
R1829 VN.n25 VN.n14 161.3
R1830 VN.n24 VN.n23 161.3
R1831 VN.n22 VN.n15 161.3
R1832 VN.n21 VN.n20 161.3
R1833 VN.n19 VN.n16 161.3
R1834 VN.n11 VN.n0 161.3
R1835 VN.n10 VN.n9 161.3
R1836 VN.n8 VN.n1 161.3
R1837 VN.n7 VN.n6 161.3
R1838 VN.n5 VN.n2 161.3
R1839 VN.n13 VN.n12 95.6613
R1840 VN.n27 VN.n26 95.6613
R1841 VN.n4 VN.n3 59.417
R1842 VN.n18 VN.n17 59.417
R1843 VN VN.n27 53.2103
R1844 VN.n10 VN.n1 43.4833
R1845 VN.n24 VN.n15 43.4833
R1846 VN.n6 VN.n1 37.6707
R1847 VN.n20 VN.n15 37.6707
R1848 VN.n6 VN.n5 24.5923
R1849 VN.n11 VN.n10 24.5923
R1850 VN.n20 VN.n19 24.5923
R1851 VN.n25 VN.n24 24.5923
R1852 VN.n12 VN.n11 15.2474
R1853 VN.n26 VN.n25 15.2474
R1854 VN.n5 VN.n4 12.2964
R1855 VN.n19 VN.n18 12.2964
R1856 VN.n17 VN.n16 9.41768
R1857 VN.n3 VN.n2 9.41768
R1858 VN.n27 VN.n14 0.278335
R1859 VN.n13 VN.n0 0.278335
R1860 VN.n23 VN.n14 0.189894
R1861 VN.n23 VN.n22 0.189894
R1862 VN.n22 VN.n21 0.189894
R1863 VN.n21 VN.n16 0.189894
R1864 VN.n7 VN.n2 0.189894
R1865 VN.n8 VN.n7 0.189894
R1866 VN.n9 VN.n8 0.189894
R1867 VN.n9 VN.n0 0.189894
R1868 VN VN.n13 0.153485
R1869 VDD2.n207 VDD2.n107 214.453
R1870 VDD2.n100 VDD2.n0 214.453
R1871 VDD2.n208 VDD2.n207 185
R1872 VDD2.n206 VDD2.n205 185
R1873 VDD2.n111 VDD2.n110 185
R1874 VDD2.n200 VDD2.n199 185
R1875 VDD2.n198 VDD2.n197 185
R1876 VDD2.n115 VDD2.n114 185
R1877 VDD2.n192 VDD2.n191 185
R1878 VDD2.n190 VDD2.n189 185
R1879 VDD2.n119 VDD2.n118 185
R1880 VDD2.n184 VDD2.n183 185
R1881 VDD2.n182 VDD2.n181 185
R1882 VDD2.n123 VDD2.n122 185
R1883 VDD2.n176 VDD2.n175 185
R1884 VDD2.n174 VDD2.n173 185
R1885 VDD2.n127 VDD2.n126 185
R1886 VDD2.n168 VDD2.n167 185
R1887 VDD2.n166 VDD2.n165 185
R1888 VDD2.n164 VDD2.n130 185
R1889 VDD2.n134 VDD2.n131 185
R1890 VDD2.n159 VDD2.n158 185
R1891 VDD2.n157 VDD2.n156 185
R1892 VDD2.n136 VDD2.n135 185
R1893 VDD2.n151 VDD2.n150 185
R1894 VDD2.n149 VDD2.n148 185
R1895 VDD2.n140 VDD2.n139 185
R1896 VDD2.n143 VDD2.n142 185
R1897 VDD2.n35 VDD2.n34 185
R1898 VDD2.n32 VDD2.n31 185
R1899 VDD2.n41 VDD2.n40 185
R1900 VDD2.n43 VDD2.n42 185
R1901 VDD2.n28 VDD2.n27 185
R1902 VDD2.n49 VDD2.n48 185
R1903 VDD2.n52 VDD2.n51 185
R1904 VDD2.n50 VDD2.n24 185
R1905 VDD2.n57 VDD2.n23 185
R1906 VDD2.n59 VDD2.n58 185
R1907 VDD2.n61 VDD2.n60 185
R1908 VDD2.n20 VDD2.n19 185
R1909 VDD2.n67 VDD2.n66 185
R1910 VDD2.n69 VDD2.n68 185
R1911 VDD2.n16 VDD2.n15 185
R1912 VDD2.n75 VDD2.n74 185
R1913 VDD2.n77 VDD2.n76 185
R1914 VDD2.n12 VDD2.n11 185
R1915 VDD2.n83 VDD2.n82 185
R1916 VDD2.n85 VDD2.n84 185
R1917 VDD2.n8 VDD2.n7 185
R1918 VDD2.n91 VDD2.n90 185
R1919 VDD2.n93 VDD2.n92 185
R1920 VDD2.n4 VDD2.n3 185
R1921 VDD2.n99 VDD2.n98 185
R1922 VDD2.n101 VDD2.n100 185
R1923 VDD2.t5 VDD2.n141 149.524
R1924 VDD2.t2 VDD2.n33 149.524
R1925 VDD2.n207 VDD2.n206 104.615
R1926 VDD2.n206 VDD2.n110 104.615
R1927 VDD2.n199 VDD2.n110 104.615
R1928 VDD2.n199 VDD2.n198 104.615
R1929 VDD2.n198 VDD2.n114 104.615
R1930 VDD2.n191 VDD2.n114 104.615
R1931 VDD2.n191 VDD2.n190 104.615
R1932 VDD2.n190 VDD2.n118 104.615
R1933 VDD2.n183 VDD2.n118 104.615
R1934 VDD2.n183 VDD2.n182 104.615
R1935 VDD2.n182 VDD2.n122 104.615
R1936 VDD2.n175 VDD2.n122 104.615
R1937 VDD2.n175 VDD2.n174 104.615
R1938 VDD2.n174 VDD2.n126 104.615
R1939 VDD2.n167 VDD2.n126 104.615
R1940 VDD2.n167 VDD2.n166 104.615
R1941 VDD2.n166 VDD2.n130 104.615
R1942 VDD2.n134 VDD2.n130 104.615
R1943 VDD2.n158 VDD2.n134 104.615
R1944 VDD2.n158 VDD2.n157 104.615
R1945 VDD2.n157 VDD2.n135 104.615
R1946 VDD2.n150 VDD2.n135 104.615
R1947 VDD2.n150 VDD2.n149 104.615
R1948 VDD2.n149 VDD2.n139 104.615
R1949 VDD2.n142 VDD2.n139 104.615
R1950 VDD2.n34 VDD2.n31 104.615
R1951 VDD2.n41 VDD2.n31 104.615
R1952 VDD2.n42 VDD2.n41 104.615
R1953 VDD2.n42 VDD2.n27 104.615
R1954 VDD2.n49 VDD2.n27 104.615
R1955 VDD2.n51 VDD2.n49 104.615
R1956 VDD2.n51 VDD2.n50 104.615
R1957 VDD2.n50 VDD2.n23 104.615
R1958 VDD2.n59 VDD2.n23 104.615
R1959 VDD2.n60 VDD2.n59 104.615
R1960 VDD2.n60 VDD2.n19 104.615
R1961 VDD2.n67 VDD2.n19 104.615
R1962 VDD2.n68 VDD2.n67 104.615
R1963 VDD2.n68 VDD2.n15 104.615
R1964 VDD2.n75 VDD2.n15 104.615
R1965 VDD2.n76 VDD2.n75 104.615
R1966 VDD2.n76 VDD2.n11 104.615
R1967 VDD2.n83 VDD2.n11 104.615
R1968 VDD2.n84 VDD2.n83 104.615
R1969 VDD2.n84 VDD2.n7 104.615
R1970 VDD2.n91 VDD2.n7 104.615
R1971 VDD2.n92 VDD2.n91 104.615
R1972 VDD2.n92 VDD2.n3 104.615
R1973 VDD2.n99 VDD2.n3 104.615
R1974 VDD2.n100 VDD2.n99 104.615
R1975 VDD2.n106 VDD2.n105 64.5768
R1976 VDD2 VDD2.n213 64.574
R1977 VDD2.n106 VDD2.n104 54.3428
R1978 VDD2.n212 VDD2.n211 52.7429
R1979 VDD2.n142 VDD2.t5 52.3082
R1980 VDD2.n34 VDD2.t2 52.3082
R1981 VDD2.n212 VDD2.n106 47.7153
R1982 VDD2.n165 VDD2.n164 13.1884
R1983 VDD2.n58 VDD2.n57 13.1884
R1984 VDD2.n209 VDD2.n208 12.8005
R1985 VDD2.n168 VDD2.n129 12.8005
R1986 VDD2.n163 VDD2.n131 12.8005
R1987 VDD2.n56 VDD2.n24 12.8005
R1988 VDD2.n61 VDD2.n22 12.8005
R1989 VDD2.n102 VDD2.n101 12.8005
R1990 VDD2.n205 VDD2.n109 12.0247
R1991 VDD2.n169 VDD2.n127 12.0247
R1992 VDD2.n160 VDD2.n159 12.0247
R1993 VDD2.n53 VDD2.n52 12.0247
R1994 VDD2.n62 VDD2.n20 12.0247
R1995 VDD2.n98 VDD2.n2 12.0247
R1996 VDD2.n204 VDD2.n111 11.249
R1997 VDD2.n173 VDD2.n172 11.249
R1998 VDD2.n156 VDD2.n133 11.249
R1999 VDD2.n48 VDD2.n26 11.249
R2000 VDD2.n66 VDD2.n65 11.249
R2001 VDD2.n97 VDD2.n4 11.249
R2002 VDD2.n201 VDD2.n200 10.4732
R2003 VDD2.n176 VDD2.n125 10.4732
R2004 VDD2.n155 VDD2.n136 10.4732
R2005 VDD2.n47 VDD2.n28 10.4732
R2006 VDD2.n69 VDD2.n18 10.4732
R2007 VDD2.n94 VDD2.n93 10.4732
R2008 VDD2.n143 VDD2.n141 10.2747
R2009 VDD2.n35 VDD2.n33 10.2747
R2010 VDD2.n197 VDD2.n113 9.69747
R2011 VDD2.n177 VDD2.n123 9.69747
R2012 VDD2.n152 VDD2.n151 9.69747
R2013 VDD2.n44 VDD2.n43 9.69747
R2014 VDD2.n70 VDD2.n16 9.69747
R2015 VDD2.n90 VDD2.n6 9.69747
R2016 VDD2.n211 VDD2.n210 9.45567
R2017 VDD2.n104 VDD2.n103 9.45567
R2018 VDD2.n145 VDD2.n144 9.3005
R2019 VDD2.n147 VDD2.n146 9.3005
R2020 VDD2.n138 VDD2.n137 9.3005
R2021 VDD2.n153 VDD2.n152 9.3005
R2022 VDD2.n155 VDD2.n154 9.3005
R2023 VDD2.n133 VDD2.n132 9.3005
R2024 VDD2.n161 VDD2.n160 9.3005
R2025 VDD2.n163 VDD2.n162 9.3005
R2026 VDD2.n117 VDD2.n116 9.3005
R2027 VDD2.n194 VDD2.n193 9.3005
R2028 VDD2.n196 VDD2.n195 9.3005
R2029 VDD2.n113 VDD2.n112 9.3005
R2030 VDD2.n202 VDD2.n201 9.3005
R2031 VDD2.n204 VDD2.n203 9.3005
R2032 VDD2.n109 VDD2.n108 9.3005
R2033 VDD2.n210 VDD2.n209 9.3005
R2034 VDD2.n188 VDD2.n187 9.3005
R2035 VDD2.n186 VDD2.n185 9.3005
R2036 VDD2.n121 VDD2.n120 9.3005
R2037 VDD2.n180 VDD2.n179 9.3005
R2038 VDD2.n178 VDD2.n177 9.3005
R2039 VDD2.n125 VDD2.n124 9.3005
R2040 VDD2.n172 VDD2.n171 9.3005
R2041 VDD2.n170 VDD2.n169 9.3005
R2042 VDD2.n129 VDD2.n128 9.3005
R2043 VDD2.n79 VDD2.n78 9.3005
R2044 VDD2.n14 VDD2.n13 9.3005
R2045 VDD2.n73 VDD2.n72 9.3005
R2046 VDD2.n71 VDD2.n70 9.3005
R2047 VDD2.n18 VDD2.n17 9.3005
R2048 VDD2.n65 VDD2.n64 9.3005
R2049 VDD2.n63 VDD2.n62 9.3005
R2050 VDD2.n22 VDD2.n21 9.3005
R2051 VDD2.n37 VDD2.n36 9.3005
R2052 VDD2.n39 VDD2.n38 9.3005
R2053 VDD2.n30 VDD2.n29 9.3005
R2054 VDD2.n45 VDD2.n44 9.3005
R2055 VDD2.n47 VDD2.n46 9.3005
R2056 VDD2.n26 VDD2.n25 9.3005
R2057 VDD2.n54 VDD2.n53 9.3005
R2058 VDD2.n56 VDD2.n55 9.3005
R2059 VDD2.n81 VDD2.n80 9.3005
R2060 VDD2.n10 VDD2.n9 9.3005
R2061 VDD2.n87 VDD2.n86 9.3005
R2062 VDD2.n89 VDD2.n88 9.3005
R2063 VDD2.n6 VDD2.n5 9.3005
R2064 VDD2.n95 VDD2.n94 9.3005
R2065 VDD2.n97 VDD2.n96 9.3005
R2066 VDD2.n2 VDD2.n1 9.3005
R2067 VDD2.n103 VDD2.n102 9.3005
R2068 VDD2.n196 VDD2.n115 8.92171
R2069 VDD2.n181 VDD2.n180 8.92171
R2070 VDD2.n148 VDD2.n138 8.92171
R2071 VDD2.n40 VDD2.n30 8.92171
R2072 VDD2.n74 VDD2.n73 8.92171
R2073 VDD2.n89 VDD2.n8 8.92171
R2074 VDD2.n211 VDD2.n107 8.2187
R2075 VDD2.n104 VDD2.n0 8.2187
R2076 VDD2.n193 VDD2.n192 8.14595
R2077 VDD2.n184 VDD2.n121 8.14595
R2078 VDD2.n147 VDD2.n140 8.14595
R2079 VDD2.n39 VDD2.n32 8.14595
R2080 VDD2.n77 VDD2.n14 8.14595
R2081 VDD2.n86 VDD2.n85 8.14595
R2082 VDD2.n189 VDD2.n117 7.3702
R2083 VDD2.n185 VDD2.n119 7.3702
R2084 VDD2.n144 VDD2.n143 7.3702
R2085 VDD2.n36 VDD2.n35 7.3702
R2086 VDD2.n78 VDD2.n12 7.3702
R2087 VDD2.n82 VDD2.n10 7.3702
R2088 VDD2.n189 VDD2.n188 6.59444
R2089 VDD2.n188 VDD2.n119 6.59444
R2090 VDD2.n81 VDD2.n12 6.59444
R2091 VDD2.n82 VDD2.n81 6.59444
R2092 VDD2.n192 VDD2.n117 5.81868
R2093 VDD2.n185 VDD2.n184 5.81868
R2094 VDD2.n144 VDD2.n140 5.81868
R2095 VDD2.n36 VDD2.n32 5.81868
R2096 VDD2.n78 VDD2.n77 5.81868
R2097 VDD2.n85 VDD2.n10 5.81868
R2098 VDD2.n209 VDD2.n107 5.3904
R2099 VDD2.n102 VDD2.n0 5.3904
R2100 VDD2.n193 VDD2.n115 5.04292
R2101 VDD2.n181 VDD2.n121 5.04292
R2102 VDD2.n148 VDD2.n147 5.04292
R2103 VDD2.n40 VDD2.n39 5.04292
R2104 VDD2.n74 VDD2.n14 5.04292
R2105 VDD2.n86 VDD2.n8 5.04292
R2106 VDD2.n197 VDD2.n196 4.26717
R2107 VDD2.n180 VDD2.n123 4.26717
R2108 VDD2.n151 VDD2.n138 4.26717
R2109 VDD2.n43 VDD2.n30 4.26717
R2110 VDD2.n73 VDD2.n16 4.26717
R2111 VDD2.n90 VDD2.n89 4.26717
R2112 VDD2.n200 VDD2.n113 3.49141
R2113 VDD2.n177 VDD2.n176 3.49141
R2114 VDD2.n152 VDD2.n136 3.49141
R2115 VDD2.n44 VDD2.n28 3.49141
R2116 VDD2.n70 VDD2.n69 3.49141
R2117 VDD2.n93 VDD2.n6 3.49141
R2118 VDD2.n37 VDD2.n33 2.84303
R2119 VDD2.n145 VDD2.n141 2.84303
R2120 VDD2.n201 VDD2.n111 2.71565
R2121 VDD2.n173 VDD2.n125 2.71565
R2122 VDD2.n156 VDD2.n155 2.71565
R2123 VDD2.n48 VDD2.n47 2.71565
R2124 VDD2.n66 VDD2.n18 2.71565
R2125 VDD2.n94 VDD2.n4 2.71565
R2126 VDD2.n205 VDD2.n204 1.93989
R2127 VDD2.n172 VDD2.n127 1.93989
R2128 VDD2.n159 VDD2.n133 1.93989
R2129 VDD2.n52 VDD2.n26 1.93989
R2130 VDD2.n65 VDD2.n20 1.93989
R2131 VDD2.n98 VDD2.n97 1.93989
R2132 VDD2 VDD2.n212 1.71386
R2133 VDD2.n208 VDD2.n109 1.16414
R2134 VDD2.n169 VDD2.n168 1.16414
R2135 VDD2.n160 VDD2.n131 1.16414
R2136 VDD2.n53 VDD2.n24 1.16414
R2137 VDD2.n62 VDD2.n61 1.16414
R2138 VDD2.n101 VDD2.n2 1.16414
R2139 VDD2.n213 VDD2.t3 1.01484
R2140 VDD2.n213 VDD2.t4 1.01484
R2141 VDD2.n105 VDD2.t1 1.01484
R2142 VDD2.n105 VDD2.t0 1.01484
R2143 VDD2.n165 VDD2.n129 0.388379
R2144 VDD2.n164 VDD2.n163 0.388379
R2145 VDD2.n57 VDD2.n56 0.388379
R2146 VDD2.n58 VDD2.n22 0.388379
R2147 VDD2.n210 VDD2.n108 0.155672
R2148 VDD2.n203 VDD2.n108 0.155672
R2149 VDD2.n203 VDD2.n202 0.155672
R2150 VDD2.n202 VDD2.n112 0.155672
R2151 VDD2.n195 VDD2.n112 0.155672
R2152 VDD2.n195 VDD2.n194 0.155672
R2153 VDD2.n194 VDD2.n116 0.155672
R2154 VDD2.n187 VDD2.n116 0.155672
R2155 VDD2.n187 VDD2.n186 0.155672
R2156 VDD2.n186 VDD2.n120 0.155672
R2157 VDD2.n179 VDD2.n120 0.155672
R2158 VDD2.n179 VDD2.n178 0.155672
R2159 VDD2.n178 VDD2.n124 0.155672
R2160 VDD2.n171 VDD2.n124 0.155672
R2161 VDD2.n171 VDD2.n170 0.155672
R2162 VDD2.n170 VDD2.n128 0.155672
R2163 VDD2.n162 VDD2.n128 0.155672
R2164 VDD2.n162 VDD2.n161 0.155672
R2165 VDD2.n161 VDD2.n132 0.155672
R2166 VDD2.n154 VDD2.n132 0.155672
R2167 VDD2.n154 VDD2.n153 0.155672
R2168 VDD2.n153 VDD2.n137 0.155672
R2169 VDD2.n146 VDD2.n137 0.155672
R2170 VDD2.n146 VDD2.n145 0.155672
R2171 VDD2.n38 VDD2.n37 0.155672
R2172 VDD2.n38 VDD2.n29 0.155672
R2173 VDD2.n45 VDD2.n29 0.155672
R2174 VDD2.n46 VDD2.n45 0.155672
R2175 VDD2.n46 VDD2.n25 0.155672
R2176 VDD2.n54 VDD2.n25 0.155672
R2177 VDD2.n55 VDD2.n54 0.155672
R2178 VDD2.n55 VDD2.n21 0.155672
R2179 VDD2.n63 VDD2.n21 0.155672
R2180 VDD2.n64 VDD2.n63 0.155672
R2181 VDD2.n64 VDD2.n17 0.155672
R2182 VDD2.n71 VDD2.n17 0.155672
R2183 VDD2.n72 VDD2.n71 0.155672
R2184 VDD2.n72 VDD2.n13 0.155672
R2185 VDD2.n79 VDD2.n13 0.155672
R2186 VDD2.n80 VDD2.n79 0.155672
R2187 VDD2.n80 VDD2.n9 0.155672
R2188 VDD2.n87 VDD2.n9 0.155672
R2189 VDD2.n88 VDD2.n87 0.155672
R2190 VDD2.n88 VDD2.n5 0.155672
R2191 VDD2.n95 VDD2.n5 0.155672
R2192 VDD2.n96 VDD2.n95 0.155672
R2193 VDD2.n96 VDD2.n1 0.155672
R2194 VDD2.n103 VDD2.n1 0.155672
R2195 VTAIL.n426 VTAIL.n326 214.453
R2196 VTAIL.n102 VTAIL.n2 214.453
R2197 VTAIL.n320 VTAIL.n220 214.453
R2198 VTAIL.n212 VTAIL.n112 214.453
R2199 VTAIL.n361 VTAIL.n360 185
R2200 VTAIL.n358 VTAIL.n357 185
R2201 VTAIL.n367 VTAIL.n366 185
R2202 VTAIL.n369 VTAIL.n368 185
R2203 VTAIL.n354 VTAIL.n353 185
R2204 VTAIL.n375 VTAIL.n374 185
R2205 VTAIL.n378 VTAIL.n377 185
R2206 VTAIL.n376 VTAIL.n350 185
R2207 VTAIL.n383 VTAIL.n349 185
R2208 VTAIL.n385 VTAIL.n384 185
R2209 VTAIL.n387 VTAIL.n386 185
R2210 VTAIL.n346 VTAIL.n345 185
R2211 VTAIL.n393 VTAIL.n392 185
R2212 VTAIL.n395 VTAIL.n394 185
R2213 VTAIL.n342 VTAIL.n341 185
R2214 VTAIL.n401 VTAIL.n400 185
R2215 VTAIL.n403 VTAIL.n402 185
R2216 VTAIL.n338 VTAIL.n337 185
R2217 VTAIL.n409 VTAIL.n408 185
R2218 VTAIL.n411 VTAIL.n410 185
R2219 VTAIL.n334 VTAIL.n333 185
R2220 VTAIL.n417 VTAIL.n416 185
R2221 VTAIL.n419 VTAIL.n418 185
R2222 VTAIL.n330 VTAIL.n329 185
R2223 VTAIL.n425 VTAIL.n424 185
R2224 VTAIL.n427 VTAIL.n426 185
R2225 VTAIL.n37 VTAIL.n36 185
R2226 VTAIL.n34 VTAIL.n33 185
R2227 VTAIL.n43 VTAIL.n42 185
R2228 VTAIL.n45 VTAIL.n44 185
R2229 VTAIL.n30 VTAIL.n29 185
R2230 VTAIL.n51 VTAIL.n50 185
R2231 VTAIL.n54 VTAIL.n53 185
R2232 VTAIL.n52 VTAIL.n26 185
R2233 VTAIL.n59 VTAIL.n25 185
R2234 VTAIL.n61 VTAIL.n60 185
R2235 VTAIL.n63 VTAIL.n62 185
R2236 VTAIL.n22 VTAIL.n21 185
R2237 VTAIL.n69 VTAIL.n68 185
R2238 VTAIL.n71 VTAIL.n70 185
R2239 VTAIL.n18 VTAIL.n17 185
R2240 VTAIL.n77 VTAIL.n76 185
R2241 VTAIL.n79 VTAIL.n78 185
R2242 VTAIL.n14 VTAIL.n13 185
R2243 VTAIL.n85 VTAIL.n84 185
R2244 VTAIL.n87 VTAIL.n86 185
R2245 VTAIL.n10 VTAIL.n9 185
R2246 VTAIL.n93 VTAIL.n92 185
R2247 VTAIL.n95 VTAIL.n94 185
R2248 VTAIL.n6 VTAIL.n5 185
R2249 VTAIL.n101 VTAIL.n100 185
R2250 VTAIL.n103 VTAIL.n102 185
R2251 VTAIL.n321 VTAIL.n320 185
R2252 VTAIL.n319 VTAIL.n318 185
R2253 VTAIL.n224 VTAIL.n223 185
R2254 VTAIL.n313 VTAIL.n312 185
R2255 VTAIL.n311 VTAIL.n310 185
R2256 VTAIL.n228 VTAIL.n227 185
R2257 VTAIL.n305 VTAIL.n304 185
R2258 VTAIL.n303 VTAIL.n302 185
R2259 VTAIL.n232 VTAIL.n231 185
R2260 VTAIL.n297 VTAIL.n296 185
R2261 VTAIL.n295 VTAIL.n294 185
R2262 VTAIL.n236 VTAIL.n235 185
R2263 VTAIL.n289 VTAIL.n288 185
R2264 VTAIL.n287 VTAIL.n286 185
R2265 VTAIL.n240 VTAIL.n239 185
R2266 VTAIL.n281 VTAIL.n280 185
R2267 VTAIL.n279 VTAIL.n278 185
R2268 VTAIL.n277 VTAIL.n243 185
R2269 VTAIL.n247 VTAIL.n244 185
R2270 VTAIL.n272 VTAIL.n271 185
R2271 VTAIL.n270 VTAIL.n269 185
R2272 VTAIL.n249 VTAIL.n248 185
R2273 VTAIL.n264 VTAIL.n263 185
R2274 VTAIL.n262 VTAIL.n261 185
R2275 VTAIL.n253 VTAIL.n252 185
R2276 VTAIL.n256 VTAIL.n255 185
R2277 VTAIL.n213 VTAIL.n212 185
R2278 VTAIL.n211 VTAIL.n210 185
R2279 VTAIL.n116 VTAIL.n115 185
R2280 VTAIL.n205 VTAIL.n204 185
R2281 VTAIL.n203 VTAIL.n202 185
R2282 VTAIL.n120 VTAIL.n119 185
R2283 VTAIL.n197 VTAIL.n196 185
R2284 VTAIL.n195 VTAIL.n194 185
R2285 VTAIL.n124 VTAIL.n123 185
R2286 VTAIL.n189 VTAIL.n188 185
R2287 VTAIL.n187 VTAIL.n186 185
R2288 VTAIL.n128 VTAIL.n127 185
R2289 VTAIL.n181 VTAIL.n180 185
R2290 VTAIL.n179 VTAIL.n178 185
R2291 VTAIL.n132 VTAIL.n131 185
R2292 VTAIL.n173 VTAIL.n172 185
R2293 VTAIL.n171 VTAIL.n170 185
R2294 VTAIL.n169 VTAIL.n135 185
R2295 VTAIL.n139 VTAIL.n136 185
R2296 VTAIL.n164 VTAIL.n163 185
R2297 VTAIL.n162 VTAIL.n161 185
R2298 VTAIL.n141 VTAIL.n140 185
R2299 VTAIL.n156 VTAIL.n155 185
R2300 VTAIL.n154 VTAIL.n153 185
R2301 VTAIL.n145 VTAIL.n144 185
R2302 VTAIL.n148 VTAIL.n147 185
R2303 VTAIL.t10 VTAIL.n359 149.524
R2304 VTAIL.t3 VTAIL.n35 149.524
R2305 VTAIL.t4 VTAIL.n254 149.524
R2306 VTAIL.t8 VTAIL.n146 149.524
R2307 VTAIL.n360 VTAIL.n357 104.615
R2308 VTAIL.n367 VTAIL.n357 104.615
R2309 VTAIL.n368 VTAIL.n367 104.615
R2310 VTAIL.n368 VTAIL.n353 104.615
R2311 VTAIL.n375 VTAIL.n353 104.615
R2312 VTAIL.n377 VTAIL.n375 104.615
R2313 VTAIL.n377 VTAIL.n376 104.615
R2314 VTAIL.n376 VTAIL.n349 104.615
R2315 VTAIL.n385 VTAIL.n349 104.615
R2316 VTAIL.n386 VTAIL.n385 104.615
R2317 VTAIL.n386 VTAIL.n345 104.615
R2318 VTAIL.n393 VTAIL.n345 104.615
R2319 VTAIL.n394 VTAIL.n393 104.615
R2320 VTAIL.n394 VTAIL.n341 104.615
R2321 VTAIL.n401 VTAIL.n341 104.615
R2322 VTAIL.n402 VTAIL.n401 104.615
R2323 VTAIL.n402 VTAIL.n337 104.615
R2324 VTAIL.n409 VTAIL.n337 104.615
R2325 VTAIL.n410 VTAIL.n409 104.615
R2326 VTAIL.n410 VTAIL.n333 104.615
R2327 VTAIL.n417 VTAIL.n333 104.615
R2328 VTAIL.n418 VTAIL.n417 104.615
R2329 VTAIL.n418 VTAIL.n329 104.615
R2330 VTAIL.n425 VTAIL.n329 104.615
R2331 VTAIL.n426 VTAIL.n425 104.615
R2332 VTAIL.n36 VTAIL.n33 104.615
R2333 VTAIL.n43 VTAIL.n33 104.615
R2334 VTAIL.n44 VTAIL.n43 104.615
R2335 VTAIL.n44 VTAIL.n29 104.615
R2336 VTAIL.n51 VTAIL.n29 104.615
R2337 VTAIL.n53 VTAIL.n51 104.615
R2338 VTAIL.n53 VTAIL.n52 104.615
R2339 VTAIL.n52 VTAIL.n25 104.615
R2340 VTAIL.n61 VTAIL.n25 104.615
R2341 VTAIL.n62 VTAIL.n61 104.615
R2342 VTAIL.n62 VTAIL.n21 104.615
R2343 VTAIL.n69 VTAIL.n21 104.615
R2344 VTAIL.n70 VTAIL.n69 104.615
R2345 VTAIL.n70 VTAIL.n17 104.615
R2346 VTAIL.n77 VTAIL.n17 104.615
R2347 VTAIL.n78 VTAIL.n77 104.615
R2348 VTAIL.n78 VTAIL.n13 104.615
R2349 VTAIL.n85 VTAIL.n13 104.615
R2350 VTAIL.n86 VTAIL.n85 104.615
R2351 VTAIL.n86 VTAIL.n9 104.615
R2352 VTAIL.n93 VTAIL.n9 104.615
R2353 VTAIL.n94 VTAIL.n93 104.615
R2354 VTAIL.n94 VTAIL.n5 104.615
R2355 VTAIL.n101 VTAIL.n5 104.615
R2356 VTAIL.n102 VTAIL.n101 104.615
R2357 VTAIL.n320 VTAIL.n319 104.615
R2358 VTAIL.n319 VTAIL.n223 104.615
R2359 VTAIL.n312 VTAIL.n223 104.615
R2360 VTAIL.n312 VTAIL.n311 104.615
R2361 VTAIL.n311 VTAIL.n227 104.615
R2362 VTAIL.n304 VTAIL.n227 104.615
R2363 VTAIL.n304 VTAIL.n303 104.615
R2364 VTAIL.n303 VTAIL.n231 104.615
R2365 VTAIL.n296 VTAIL.n231 104.615
R2366 VTAIL.n296 VTAIL.n295 104.615
R2367 VTAIL.n295 VTAIL.n235 104.615
R2368 VTAIL.n288 VTAIL.n235 104.615
R2369 VTAIL.n288 VTAIL.n287 104.615
R2370 VTAIL.n287 VTAIL.n239 104.615
R2371 VTAIL.n280 VTAIL.n239 104.615
R2372 VTAIL.n280 VTAIL.n279 104.615
R2373 VTAIL.n279 VTAIL.n243 104.615
R2374 VTAIL.n247 VTAIL.n243 104.615
R2375 VTAIL.n271 VTAIL.n247 104.615
R2376 VTAIL.n271 VTAIL.n270 104.615
R2377 VTAIL.n270 VTAIL.n248 104.615
R2378 VTAIL.n263 VTAIL.n248 104.615
R2379 VTAIL.n263 VTAIL.n262 104.615
R2380 VTAIL.n262 VTAIL.n252 104.615
R2381 VTAIL.n255 VTAIL.n252 104.615
R2382 VTAIL.n212 VTAIL.n211 104.615
R2383 VTAIL.n211 VTAIL.n115 104.615
R2384 VTAIL.n204 VTAIL.n115 104.615
R2385 VTAIL.n204 VTAIL.n203 104.615
R2386 VTAIL.n203 VTAIL.n119 104.615
R2387 VTAIL.n196 VTAIL.n119 104.615
R2388 VTAIL.n196 VTAIL.n195 104.615
R2389 VTAIL.n195 VTAIL.n123 104.615
R2390 VTAIL.n188 VTAIL.n123 104.615
R2391 VTAIL.n188 VTAIL.n187 104.615
R2392 VTAIL.n187 VTAIL.n127 104.615
R2393 VTAIL.n180 VTAIL.n127 104.615
R2394 VTAIL.n180 VTAIL.n179 104.615
R2395 VTAIL.n179 VTAIL.n131 104.615
R2396 VTAIL.n172 VTAIL.n131 104.615
R2397 VTAIL.n172 VTAIL.n171 104.615
R2398 VTAIL.n171 VTAIL.n135 104.615
R2399 VTAIL.n139 VTAIL.n135 104.615
R2400 VTAIL.n163 VTAIL.n139 104.615
R2401 VTAIL.n163 VTAIL.n162 104.615
R2402 VTAIL.n162 VTAIL.n140 104.615
R2403 VTAIL.n155 VTAIL.n140 104.615
R2404 VTAIL.n155 VTAIL.n154 104.615
R2405 VTAIL.n154 VTAIL.n144 104.615
R2406 VTAIL.n147 VTAIL.n144 104.615
R2407 VTAIL.n360 VTAIL.t10 52.3082
R2408 VTAIL.n36 VTAIL.t3 52.3082
R2409 VTAIL.n255 VTAIL.t4 52.3082
R2410 VTAIL.n147 VTAIL.t8 52.3082
R2411 VTAIL.n219 VTAIL.n218 47.4018
R2412 VTAIL.n111 VTAIL.n110 47.4018
R2413 VTAIL.n1 VTAIL.n0 47.4016
R2414 VTAIL.n109 VTAIL.n108 47.4016
R2415 VTAIL.n431 VTAIL.n430 36.0641
R2416 VTAIL.n107 VTAIL.n106 36.0641
R2417 VTAIL.n325 VTAIL.n324 36.0641
R2418 VTAIL.n217 VTAIL.n216 36.0641
R2419 VTAIL.n111 VTAIL.n109 33.6083
R2420 VTAIL.n431 VTAIL.n325 31.4014
R2421 VTAIL.n384 VTAIL.n383 13.1884
R2422 VTAIL.n60 VTAIL.n59 13.1884
R2423 VTAIL.n278 VTAIL.n277 13.1884
R2424 VTAIL.n170 VTAIL.n169 13.1884
R2425 VTAIL.n382 VTAIL.n350 12.8005
R2426 VTAIL.n387 VTAIL.n348 12.8005
R2427 VTAIL.n428 VTAIL.n427 12.8005
R2428 VTAIL.n58 VTAIL.n26 12.8005
R2429 VTAIL.n63 VTAIL.n24 12.8005
R2430 VTAIL.n104 VTAIL.n103 12.8005
R2431 VTAIL.n322 VTAIL.n321 12.8005
R2432 VTAIL.n281 VTAIL.n242 12.8005
R2433 VTAIL.n276 VTAIL.n244 12.8005
R2434 VTAIL.n214 VTAIL.n213 12.8005
R2435 VTAIL.n173 VTAIL.n134 12.8005
R2436 VTAIL.n168 VTAIL.n136 12.8005
R2437 VTAIL.n379 VTAIL.n378 12.0247
R2438 VTAIL.n388 VTAIL.n346 12.0247
R2439 VTAIL.n424 VTAIL.n328 12.0247
R2440 VTAIL.n55 VTAIL.n54 12.0247
R2441 VTAIL.n64 VTAIL.n22 12.0247
R2442 VTAIL.n100 VTAIL.n4 12.0247
R2443 VTAIL.n318 VTAIL.n222 12.0247
R2444 VTAIL.n282 VTAIL.n240 12.0247
R2445 VTAIL.n273 VTAIL.n272 12.0247
R2446 VTAIL.n210 VTAIL.n114 12.0247
R2447 VTAIL.n174 VTAIL.n132 12.0247
R2448 VTAIL.n165 VTAIL.n164 12.0247
R2449 VTAIL.n374 VTAIL.n352 11.249
R2450 VTAIL.n392 VTAIL.n391 11.249
R2451 VTAIL.n423 VTAIL.n330 11.249
R2452 VTAIL.n50 VTAIL.n28 11.249
R2453 VTAIL.n68 VTAIL.n67 11.249
R2454 VTAIL.n99 VTAIL.n6 11.249
R2455 VTAIL.n317 VTAIL.n224 11.249
R2456 VTAIL.n286 VTAIL.n285 11.249
R2457 VTAIL.n269 VTAIL.n246 11.249
R2458 VTAIL.n209 VTAIL.n116 11.249
R2459 VTAIL.n178 VTAIL.n177 11.249
R2460 VTAIL.n161 VTAIL.n138 11.249
R2461 VTAIL.n373 VTAIL.n354 10.4732
R2462 VTAIL.n395 VTAIL.n344 10.4732
R2463 VTAIL.n420 VTAIL.n419 10.4732
R2464 VTAIL.n49 VTAIL.n30 10.4732
R2465 VTAIL.n71 VTAIL.n20 10.4732
R2466 VTAIL.n96 VTAIL.n95 10.4732
R2467 VTAIL.n314 VTAIL.n313 10.4732
R2468 VTAIL.n289 VTAIL.n238 10.4732
R2469 VTAIL.n268 VTAIL.n249 10.4732
R2470 VTAIL.n206 VTAIL.n205 10.4732
R2471 VTAIL.n181 VTAIL.n130 10.4732
R2472 VTAIL.n160 VTAIL.n141 10.4732
R2473 VTAIL.n361 VTAIL.n359 10.2747
R2474 VTAIL.n37 VTAIL.n35 10.2747
R2475 VTAIL.n256 VTAIL.n254 10.2747
R2476 VTAIL.n148 VTAIL.n146 10.2747
R2477 VTAIL.n370 VTAIL.n369 9.69747
R2478 VTAIL.n396 VTAIL.n342 9.69747
R2479 VTAIL.n416 VTAIL.n332 9.69747
R2480 VTAIL.n46 VTAIL.n45 9.69747
R2481 VTAIL.n72 VTAIL.n18 9.69747
R2482 VTAIL.n92 VTAIL.n8 9.69747
R2483 VTAIL.n310 VTAIL.n226 9.69747
R2484 VTAIL.n290 VTAIL.n236 9.69747
R2485 VTAIL.n265 VTAIL.n264 9.69747
R2486 VTAIL.n202 VTAIL.n118 9.69747
R2487 VTAIL.n182 VTAIL.n128 9.69747
R2488 VTAIL.n157 VTAIL.n156 9.69747
R2489 VTAIL.n430 VTAIL.n429 9.45567
R2490 VTAIL.n106 VTAIL.n105 9.45567
R2491 VTAIL.n324 VTAIL.n323 9.45567
R2492 VTAIL.n216 VTAIL.n215 9.45567
R2493 VTAIL.n405 VTAIL.n404 9.3005
R2494 VTAIL.n340 VTAIL.n339 9.3005
R2495 VTAIL.n399 VTAIL.n398 9.3005
R2496 VTAIL.n397 VTAIL.n396 9.3005
R2497 VTAIL.n344 VTAIL.n343 9.3005
R2498 VTAIL.n391 VTAIL.n390 9.3005
R2499 VTAIL.n389 VTAIL.n388 9.3005
R2500 VTAIL.n348 VTAIL.n347 9.3005
R2501 VTAIL.n363 VTAIL.n362 9.3005
R2502 VTAIL.n365 VTAIL.n364 9.3005
R2503 VTAIL.n356 VTAIL.n355 9.3005
R2504 VTAIL.n371 VTAIL.n370 9.3005
R2505 VTAIL.n373 VTAIL.n372 9.3005
R2506 VTAIL.n352 VTAIL.n351 9.3005
R2507 VTAIL.n380 VTAIL.n379 9.3005
R2508 VTAIL.n382 VTAIL.n381 9.3005
R2509 VTAIL.n407 VTAIL.n406 9.3005
R2510 VTAIL.n336 VTAIL.n335 9.3005
R2511 VTAIL.n413 VTAIL.n412 9.3005
R2512 VTAIL.n415 VTAIL.n414 9.3005
R2513 VTAIL.n332 VTAIL.n331 9.3005
R2514 VTAIL.n421 VTAIL.n420 9.3005
R2515 VTAIL.n423 VTAIL.n422 9.3005
R2516 VTAIL.n328 VTAIL.n327 9.3005
R2517 VTAIL.n429 VTAIL.n428 9.3005
R2518 VTAIL.n81 VTAIL.n80 9.3005
R2519 VTAIL.n16 VTAIL.n15 9.3005
R2520 VTAIL.n75 VTAIL.n74 9.3005
R2521 VTAIL.n73 VTAIL.n72 9.3005
R2522 VTAIL.n20 VTAIL.n19 9.3005
R2523 VTAIL.n67 VTAIL.n66 9.3005
R2524 VTAIL.n65 VTAIL.n64 9.3005
R2525 VTAIL.n24 VTAIL.n23 9.3005
R2526 VTAIL.n39 VTAIL.n38 9.3005
R2527 VTAIL.n41 VTAIL.n40 9.3005
R2528 VTAIL.n32 VTAIL.n31 9.3005
R2529 VTAIL.n47 VTAIL.n46 9.3005
R2530 VTAIL.n49 VTAIL.n48 9.3005
R2531 VTAIL.n28 VTAIL.n27 9.3005
R2532 VTAIL.n56 VTAIL.n55 9.3005
R2533 VTAIL.n58 VTAIL.n57 9.3005
R2534 VTAIL.n83 VTAIL.n82 9.3005
R2535 VTAIL.n12 VTAIL.n11 9.3005
R2536 VTAIL.n89 VTAIL.n88 9.3005
R2537 VTAIL.n91 VTAIL.n90 9.3005
R2538 VTAIL.n8 VTAIL.n7 9.3005
R2539 VTAIL.n97 VTAIL.n96 9.3005
R2540 VTAIL.n99 VTAIL.n98 9.3005
R2541 VTAIL.n4 VTAIL.n3 9.3005
R2542 VTAIL.n105 VTAIL.n104 9.3005
R2543 VTAIL.n258 VTAIL.n257 9.3005
R2544 VTAIL.n260 VTAIL.n259 9.3005
R2545 VTAIL.n251 VTAIL.n250 9.3005
R2546 VTAIL.n266 VTAIL.n265 9.3005
R2547 VTAIL.n268 VTAIL.n267 9.3005
R2548 VTAIL.n246 VTAIL.n245 9.3005
R2549 VTAIL.n274 VTAIL.n273 9.3005
R2550 VTAIL.n276 VTAIL.n275 9.3005
R2551 VTAIL.n230 VTAIL.n229 9.3005
R2552 VTAIL.n307 VTAIL.n306 9.3005
R2553 VTAIL.n309 VTAIL.n308 9.3005
R2554 VTAIL.n226 VTAIL.n225 9.3005
R2555 VTAIL.n315 VTAIL.n314 9.3005
R2556 VTAIL.n317 VTAIL.n316 9.3005
R2557 VTAIL.n222 VTAIL.n221 9.3005
R2558 VTAIL.n323 VTAIL.n322 9.3005
R2559 VTAIL.n301 VTAIL.n300 9.3005
R2560 VTAIL.n299 VTAIL.n298 9.3005
R2561 VTAIL.n234 VTAIL.n233 9.3005
R2562 VTAIL.n293 VTAIL.n292 9.3005
R2563 VTAIL.n291 VTAIL.n290 9.3005
R2564 VTAIL.n238 VTAIL.n237 9.3005
R2565 VTAIL.n285 VTAIL.n284 9.3005
R2566 VTAIL.n283 VTAIL.n282 9.3005
R2567 VTAIL.n242 VTAIL.n241 9.3005
R2568 VTAIL.n150 VTAIL.n149 9.3005
R2569 VTAIL.n152 VTAIL.n151 9.3005
R2570 VTAIL.n143 VTAIL.n142 9.3005
R2571 VTAIL.n158 VTAIL.n157 9.3005
R2572 VTAIL.n160 VTAIL.n159 9.3005
R2573 VTAIL.n138 VTAIL.n137 9.3005
R2574 VTAIL.n166 VTAIL.n165 9.3005
R2575 VTAIL.n168 VTAIL.n167 9.3005
R2576 VTAIL.n122 VTAIL.n121 9.3005
R2577 VTAIL.n199 VTAIL.n198 9.3005
R2578 VTAIL.n201 VTAIL.n200 9.3005
R2579 VTAIL.n118 VTAIL.n117 9.3005
R2580 VTAIL.n207 VTAIL.n206 9.3005
R2581 VTAIL.n209 VTAIL.n208 9.3005
R2582 VTAIL.n114 VTAIL.n113 9.3005
R2583 VTAIL.n215 VTAIL.n214 9.3005
R2584 VTAIL.n193 VTAIL.n192 9.3005
R2585 VTAIL.n191 VTAIL.n190 9.3005
R2586 VTAIL.n126 VTAIL.n125 9.3005
R2587 VTAIL.n185 VTAIL.n184 9.3005
R2588 VTAIL.n183 VTAIL.n182 9.3005
R2589 VTAIL.n130 VTAIL.n129 9.3005
R2590 VTAIL.n177 VTAIL.n176 9.3005
R2591 VTAIL.n175 VTAIL.n174 9.3005
R2592 VTAIL.n134 VTAIL.n133 9.3005
R2593 VTAIL.n366 VTAIL.n356 8.92171
R2594 VTAIL.n400 VTAIL.n399 8.92171
R2595 VTAIL.n415 VTAIL.n334 8.92171
R2596 VTAIL.n42 VTAIL.n32 8.92171
R2597 VTAIL.n76 VTAIL.n75 8.92171
R2598 VTAIL.n91 VTAIL.n10 8.92171
R2599 VTAIL.n309 VTAIL.n228 8.92171
R2600 VTAIL.n294 VTAIL.n293 8.92171
R2601 VTAIL.n261 VTAIL.n251 8.92171
R2602 VTAIL.n201 VTAIL.n120 8.92171
R2603 VTAIL.n186 VTAIL.n185 8.92171
R2604 VTAIL.n153 VTAIL.n143 8.92171
R2605 VTAIL.n430 VTAIL.n326 8.2187
R2606 VTAIL.n106 VTAIL.n2 8.2187
R2607 VTAIL.n324 VTAIL.n220 8.2187
R2608 VTAIL.n216 VTAIL.n112 8.2187
R2609 VTAIL.n365 VTAIL.n358 8.14595
R2610 VTAIL.n403 VTAIL.n340 8.14595
R2611 VTAIL.n412 VTAIL.n411 8.14595
R2612 VTAIL.n41 VTAIL.n34 8.14595
R2613 VTAIL.n79 VTAIL.n16 8.14595
R2614 VTAIL.n88 VTAIL.n87 8.14595
R2615 VTAIL.n306 VTAIL.n305 8.14595
R2616 VTAIL.n297 VTAIL.n234 8.14595
R2617 VTAIL.n260 VTAIL.n253 8.14595
R2618 VTAIL.n198 VTAIL.n197 8.14595
R2619 VTAIL.n189 VTAIL.n126 8.14595
R2620 VTAIL.n152 VTAIL.n145 8.14595
R2621 VTAIL.n362 VTAIL.n361 7.3702
R2622 VTAIL.n404 VTAIL.n338 7.3702
R2623 VTAIL.n408 VTAIL.n336 7.3702
R2624 VTAIL.n38 VTAIL.n37 7.3702
R2625 VTAIL.n80 VTAIL.n14 7.3702
R2626 VTAIL.n84 VTAIL.n12 7.3702
R2627 VTAIL.n302 VTAIL.n230 7.3702
R2628 VTAIL.n298 VTAIL.n232 7.3702
R2629 VTAIL.n257 VTAIL.n256 7.3702
R2630 VTAIL.n194 VTAIL.n122 7.3702
R2631 VTAIL.n190 VTAIL.n124 7.3702
R2632 VTAIL.n149 VTAIL.n148 7.3702
R2633 VTAIL.n407 VTAIL.n338 6.59444
R2634 VTAIL.n408 VTAIL.n407 6.59444
R2635 VTAIL.n83 VTAIL.n14 6.59444
R2636 VTAIL.n84 VTAIL.n83 6.59444
R2637 VTAIL.n302 VTAIL.n301 6.59444
R2638 VTAIL.n301 VTAIL.n232 6.59444
R2639 VTAIL.n194 VTAIL.n193 6.59444
R2640 VTAIL.n193 VTAIL.n124 6.59444
R2641 VTAIL.n362 VTAIL.n358 5.81868
R2642 VTAIL.n404 VTAIL.n403 5.81868
R2643 VTAIL.n411 VTAIL.n336 5.81868
R2644 VTAIL.n38 VTAIL.n34 5.81868
R2645 VTAIL.n80 VTAIL.n79 5.81868
R2646 VTAIL.n87 VTAIL.n12 5.81868
R2647 VTAIL.n305 VTAIL.n230 5.81868
R2648 VTAIL.n298 VTAIL.n297 5.81868
R2649 VTAIL.n257 VTAIL.n253 5.81868
R2650 VTAIL.n197 VTAIL.n122 5.81868
R2651 VTAIL.n190 VTAIL.n189 5.81868
R2652 VTAIL.n149 VTAIL.n145 5.81868
R2653 VTAIL.n428 VTAIL.n326 5.3904
R2654 VTAIL.n104 VTAIL.n2 5.3904
R2655 VTAIL.n322 VTAIL.n220 5.3904
R2656 VTAIL.n214 VTAIL.n112 5.3904
R2657 VTAIL.n366 VTAIL.n365 5.04292
R2658 VTAIL.n400 VTAIL.n340 5.04292
R2659 VTAIL.n412 VTAIL.n334 5.04292
R2660 VTAIL.n42 VTAIL.n41 5.04292
R2661 VTAIL.n76 VTAIL.n16 5.04292
R2662 VTAIL.n88 VTAIL.n10 5.04292
R2663 VTAIL.n306 VTAIL.n228 5.04292
R2664 VTAIL.n294 VTAIL.n234 5.04292
R2665 VTAIL.n261 VTAIL.n260 5.04292
R2666 VTAIL.n198 VTAIL.n120 5.04292
R2667 VTAIL.n186 VTAIL.n126 5.04292
R2668 VTAIL.n153 VTAIL.n152 5.04292
R2669 VTAIL.n369 VTAIL.n356 4.26717
R2670 VTAIL.n399 VTAIL.n342 4.26717
R2671 VTAIL.n416 VTAIL.n415 4.26717
R2672 VTAIL.n45 VTAIL.n32 4.26717
R2673 VTAIL.n75 VTAIL.n18 4.26717
R2674 VTAIL.n92 VTAIL.n91 4.26717
R2675 VTAIL.n310 VTAIL.n309 4.26717
R2676 VTAIL.n293 VTAIL.n236 4.26717
R2677 VTAIL.n264 VTAIL.n251 4.26717
R2678 VTAIL.n202 VTAIL.n201 4.26717
R2679 VTAIL.n185 VTAIL.n128 4.26717
R2680 VTAIL.n156 VTAIL.n143 4.26717
R2681 VTAIL.n370 VTAIL.n354 3.49141
R2682 VTAIL.n396 VTAIL.n395 3.49141
R2683 VTAIL.n419 VTAIL.n332 3.49141
R2684 VTAIL.n46 VTAIL.n30 3.49141
R2685 VTAIL.n72 VTAIL.n71 3.49141
R2686 VTAIL.n95 VTAIL.n8 3.49141
R2687 VTAIL.n313 VTAIL.n226 3.49141
R2688 VTAIL.n290 VTAIL.n289 3.49141
R2689 VTAIL.n265 VTAIL.n249 3.49141
R2690 VTAIL.n205 VTAIL.n118 3.49141
R2691 VTAIL.n182 VTAIL.n181 3.49141
R2692 VTAIL.n157 VTAIL.n141 3.49141
R2693 VTAIL.n363 VTAIL.n359 2.84303
R2694 VTAIL.n39 VTAIL.n35 2.84303
R2695 VTAIL.n258 VTAIL.n254 2.84303
R2696 VTAIL.n150 VTAIL.n146 2.84303
R2697 VTAIL.n374 VTAIL.n373 2.71565
R2698 VTAIL.n392 VTAIL.n344 2.71565
R2699 VTAIL.n420 VTAIL.n330 2.71565
R2700 VTAIL.n50 VTAIL.n49 2.71565
R2701 VTAIL.n68 VTAIL.n20 2.71565
R2702 VTAIL.n96 VTAIL.n6 2.71565
R2703 VTAIL.n314 VTAIL.n224 2.71565
R2704 VTAIL.n286 VTAIL.n238 2.71565
R2705 VTAIL.n269 VTAIL.n268 2.71565
R2706 VTAIL.n206 VTAIL.n116 2.71565
R2707 VTAIL.n178 VTAIL.n130 2.71565
R2708 VTAIL.n161 VTAIL.n160 2.71565
R2709 VTAIL.n217 VTAIL.n111 2.2074
R2710 VTAIL.n325 VTAIL.n219 2.2074
R2711 VTAIL.n109 VTAIL.n107 2.2074
R2712 VTAIL.n378 VTAIL.n352 1.93989
R2713 VTAIL.n391 VTAIL.n346 1.93989
R2714 VTAIL.n424 VTAIL.n423 1.93989
R2715 VTAIL.n54 VTAIL.n28 1.93989
R2716 VTAIL.n67 VTAIL.n22 1.93989
R2717 VTAIL.n100 VTAIL.n99 1.93989
R2718 VTAIL.n318 VTAIL.n317 1.93989
R2719 VTAIL.n285 VTAIL.n240 1.93989
R2720 VTAIL.n272 VTAIL.n246 1.93989
R2721 VTAIL.n210 VTAIL.n209 1.93989
R2722 VTAIL.n177 VTAIL.n132 1.93989
R2723 VTAIL.n164 VTAIL.n138 1.93989
R2724 VTAIL VTAIL.n431 1.59748
R2725 VTAIL.n219 VTAIL.n217 1.57378
R2726 VTAIL.n107 VTAIL.n1 1.57378
R2727 VTAIL.n379 VTAIL.n350 1.16414
R2728 VTAIL.n388 VTAIL.n387 1.16414
R2729 VTAIL.n427 VTAIL.n328 1.16414
R2730 VTAIL.n55 VTAIL.n26 1.16414
R2731 VTAIL.n64 VTAIL.n63 1.16414
R2732 VTAIL.n103 VTAIL.n4 1.16414
R2733 VTAIL.n321 VTAIL.n222 1.16414
R2734 VTAIL.n282 VTAIL.n281 1.16414
R2735 VTAIL.n273 VTAIL.n244 1.16414
R2736 VTAIL.n213 VTAIL.n114 1.16414
R2737 VTAIL.n174 VTAIL.n173 1.16414
R2738 VTAIL.n165 VTAIL.n136 1.16414
R2739 VTAIL.n0 VTAIL.t6 1.01484
R2740 VTAIL.n0 VTAIL.t9 1.01484
R2741 VTAIL.n108 VTAIL.t0 1.01484
R2742 VTAIL.n108 VTAIL.t5 1.01484
R2743 VTAIL.n218 VTAIL.t2 1.01484
R2744 VTAIL.n218 VTAIL.t1 1.01484
R2745 VTAIL.n110 VTAIL.t7 1.01484
R2746 VTAIL.n110 VTAIL.t11 1.01484
R2747 VTAIL VTAIL.n1 0.610414
R2748 VTAIL.n383 VTAIL.n382 0.388379
R2749 VTAIL.n384 VTAIL.n348 0.388379
R2750 VTAIL.n59 VTAIL.n58 0.388379
R2751 VTAIL.n60 VTAIL.n24 0.388379
R2752 VTAIL.n278 VTAIL.n242 0.388379
R2753 VTAIL.n277 VTAIL.n276 0.388379
R2754 VTAIL.n170 VTAIL.n134 0.388379
R2755 VTAIL.n169 VTAIL.n168 0.388379
R2756 VTAIL.n364 VTAIL.n363 0.155672
R2757 VTAIL.n364 VTAIL.n355 0.155672
R2758 VTAIL.n371 VTAIL.n355 0.155672
R2759 VTAIL.n372 VTAIL.n371 0.155672
R2760 VTAIL.n372 VTAIL.n351 0.155672
R2761 VTAIL.n380 VTAIL.n351 0.155672
R2762 VTAIL.n381 VTAIL.n380 0.155672
R2763 VTAIL.n381 VTAIL.n347 0.155672
R2764 VTAIL.n389 VTAIL.n347 0.155672
R2765 VTAIL.n390 VTAIL.n389 0.155672
R2766 VTAIL.n390 VTAIL.n343 0.155672
R2767 VTAIL.n397 VTAIL.n343 0.155672
R2768 VTAIL.n398 VTAIL.n397 0.155672
R2769 VTAIL.n398 VTAIL.n339 0.155672
R2770 VTAIL.n405 VTAIL.n339 0.155672
R2771 VTAIL.n406 VTAIL.n405 0.155672
R2772 VTAIL.n406 VTAIL.n335 0.155672
R2773 VTAIL.n413 VTAIL.n335 0.155672
R2774 VTAIL.n414 VTAIL.n413 0.155672
R2775 VTAIL.n414 VTAIL.n331 0.155672
R2776 VTAIL.n421 VTAIL.n331 0.155672
R2777 VTAIL.n422 VTAIL.n421 0.155672
R2778 VTAIL.n422 VTAIL.n327 0.155672
R2779 VTAIL.n429 VTAIL.n327 0.155672
R2780 VTAIL.n40 VTAIL.n39 0.155672
R2781 VTAIL.n40 VTAIL.n31 0.155672
R2782 VTAIL.n47 VTAIL.n31 0.155672
R2783 VTAIL.n48 VTAIL.n47 0.155672
R2784 VTAIL.n48 VTAIL.n27 0.155672
R2785 VTAIL.n56 VTAIL.n27 0.155672
R2786 VTAIL.n57 VTAIL.n56 0.155672
R2787 VTAIL.n57 VTAIL.n23 0.155672
R2788 VTAIL.n65 VTAIL.n23 0.155672
R2789 VTAIL.n66 VTAIL.n65 0.155672
R2790 VTAIL.n66 VTAIL.n19 0.155672
R2791 VTAIL.n73 VTAIL.n19 0.155672
R2792 VTAIL.n74 VTAIL.n73 0.155672
R2793 VTAIL.n74 VTAIL.n15 0.155672
R2794 VTAIL.n81 VTAIL.n15 0.155672
R2795 VTAIL.n82 VTAIL.n81 0.155672
R2796 VTAIL.n82 VTAIL.n11 0.155672
R2797 VTAIL.n89 VTAIL.n11 0.155672
R2798 VTAIL.n90 VTAIL.n89 0.155672
R2799 VTAIL.n90 VTAIL.n7 0.155672
R2800 VTAIL.n97 VTAIL.n7 0.155672
R2801 VTAIL.n98 VTAIL.n97 0.155672
R2802 VTAIL.n98 VTAIL.n3 0.155672
R2803 VTAIL.n105 VTAIL.n3 0.155672
R2804 VTAIL.n323 VTAIL.n221 0.155672
R2805 VTAIL.n316 VTAIL.n221 0.155672
R2806 VTAIL.n316 VTAIL.n315 0.155672
R2807 VTAIL.n315 VTAIL.n225 0.155672
R2808 VTAIL.n308 VTAIL.n225 0.155672
R2809 VTAIL.n308 VTAIL.n307 0.155672
R2810 VTAIL.n307 VTAIL.n229 0.155672
R2811 VTAIL.n300 VTAIL.n229 0.155672
R2812 VTAIL.n300 VTAIL.n299 0.155672
R2813 VTAIL.n299 VTAIL.n233 0.155672
R2814 VTAIL.n292 VTAIL.n233 0.155672
R2815 VTAIL.n292 VTAIL.n291 0.155672
R2816 VTAIL.n291 VTAIL.n237 0.155672
R2817 VTAIL.n284 VTAIL.n237 0.155672
R2818 VTAIL.n284 VTAIL.n283 0.155672
R2819 VTAIL.n283 VTAIL.n241 0.155672
R2820 VTAIL.n275 VTAIL.n241 0.155672
R2821 VTAIL.n275 VTAIL.n274 0.155672
R2822 VTAIL.n274 VTAIL.n245 0.155672
R2823 VTAIL.n267 VTAIL.n245 0.155672
R2824 VTAIL.n267 VTAIL.n266 0.155672
R2825 VTAIL.n266 VTAIL.n250 0.155672
R2826 VTAIL.n259 VTAIL.n250 0.155672
R2827 VTAIL.n259 VTAIL.n258 0.155672
R2828 VTAIL.n215 VTAIL.n113 0.155672
R2829 VTAIL.n208 VTAIL.n113 0.155672
R2830 VTAIL.n208 VTAIL.n207 0.155672
R2831 VTAIL.n207 VTAIL.n117 0.155672
R2832 VTAIL.n200 VTAIL.n117 0.155672
R2833 VTAIL.n200 VTAIL.n199 0.155672
R2834 VTAIL.n199 VTAIL.n121 0.155672
R2835 VTAIL.n192 VTAIL.n121 0.155672
R2836 VTAIL.n192 VTAIL.n191 0.155672
R2837 VTAIL.n191 VTAIL.n125 0.155672
R2838 VTAIL.n184 VTAIL.n125 0.155672
R2839 VTAIL.n184 VTAIL.n183 0.155672
R2840 VTAIL.n183 VTAIL.n129 0.155672
R2841 VTAIL.n176 VTAIL.n129 0.155672
R2842 VTAIL.n176 VTAIL.n175 0.155672
R2843 VTAIL.n175 VTAIL.n133 0.155672
R2844 VTAIL.n167 VTAIL.n133 0.155672
R2845 VTAIL.n167 VTAIL.n166 0.155672
R2846 VTAIL.n166 VTAIL.n137 0.155672
R2847 VTAIL.n159 VTAIL.n137 0.155672
R2848 VTAIL.n159 VTAIL.n158 0.155672
R2849 VTAIL.n158 VTAIL.n142 0.155672
R2850 VTAIL.n151 VTAIL.n142 0.155672
R2851 VTAIL.n151 VTAIL.n150 0.155672
R2852 VP.n9 VP.t0 243.868
R2853 VP.n5 VP.t5 210.957
R2854 VP.n29 VP.t1 210.957
R2855 VP.n37 VP.t3 210.957
R2856 VP.n18 VP.t2 210.957
R2857 VP.n10 VP.t4 210.957
R2858 VP.n11 VP.n8 161.3
R2859 VP.n13 VP.n12 161.3
R2860 VP.n14 VP.n7 161.3
R2861 VP.n16 VP.n15 161.3
R2862 VP.n17 VP.n6 161.3
R2863 VP.n36 VP.n0 161.3
R2864 VP.n35 VP.n34 161.3
R2865 VP.n33 VP.n1 161.3
R2866 VP.n32 VP.n31 161.3
R2867 VP.n30 VP.n2 161.3
R2868 VP.n28 VP.n27 161.3
R2869 VP.n26 VP.n3 161.3
R2870 VP.n25 VP.n24 161.3
R2871 VP.n23 VP.n4 161.3
R2872 VP.n22 VP.n21 161.3
R2873 VP.n20 VP.n5 95.6613
R2874 VP.n38 VP.n37 95.6613
R2875 VP.n19 VP.n18 95.6613
R2876 VP.n10 VP.n9 59.417
R2877 VP.n20 VP.n19 52.9315
R2878 VP.n24 VP.n23 43.4833
R2879 VP.n35 VP.n1 43.4833
R2880 VP.n16 VP.n7 43.4833
R2881 VP.n24 VP.n3 37.6707
R2882 VP.n31 VP.n1 37.6707
R2883 VP.n12 VP.n7 37.6707
R2884 VP.n23 VP.n22 24.5923
R2885 VP.n28 VP.n3 24.5923
R2886 VP.n31 VP.n30 24.5923
R2887 VP.n36 VP.n35 24.5923
R2888 VP.n17 VP.n16 24.5923
R2889 VP.n12 VP.n11 24.5923
R2890 VP.n22 VP.n5 15.2474
R2891 VP.n37 VP.n36 15.2474
R2892 VP.n18 VP.n17 15.2474
R2893 VP.n29 VP.n28 12.2964
R2894 VP.n30 VP.n29 12.2964
R2895 VP.n11 VP.n10 12.2964
R2896 VP.n9 VP.n8 9.41768
R2897 VP.n19 VP.n6 0.278335
R2898 VP.n21 VP.n20 0.278335
R2899 VP.n38 VP.n0 0.278335
R2900 VP.n13 VP.n8 0.189894
R2901 VP.n14 VP.n13 0.189894
R2902 VP.n15 VP.n14 0.189894
R2903 VP.n15 VP.n6 0.189894
R2904 VP.n21 VP.n4 0.189894
R2905 VP.n25 VP.n4 0.189894
R2906 VP.n26 VP.n25 0.189894
R2907 VP.n27 VP.n26 0.189894
R2908 VP.n27 VP.n2 0.189894
R2909 VP.n32 VP.n2 0.189894
R2910 VP.n33 VP.n32 0.189894
R2911 VP.n34 VP.n33 0.189894
R2912 VP.n34 VP.n0 0.189894
R2913 VP VP.n38 0.153485
R2914 VDD1.n100 VDD1.n0 214.453
R2915 VDD1.n205 VDD1.n105 214.453
R2916 VDD1.n101 VDD1.n100 185
R2917 VDD1.n99 VDD1.n98 185
R2918 VDD1.n4 VDD1.n3 185
R2919 VDD1.n93 VDD1.n92 185
R2920 VDD1.n91 VDD1.n90 185
R2921 VDD1.n8 VDD1.n7 185
R2922 VDD1.n85 VDD1.n84 185
R2923 VDD1.n83 VDD1.n82 185
R2924 VDD1.n12 VDD1.n11 185
R2925 VDD1.n77 VDD1.n76 185
R2926 VDD1.n75 VDD1.n74 185
R2927 VDD1.n16 VDD1.n15 185
R2928 VDD1.n69 VDD1.n68 185
R2929 VDD1.n67 VDD1.n66 185
R2930 VDD1.n20 VDD1.n19 185
R2931 VDD1.n61 VDD1.n60 185
R2932 VDD1.n59 VDD1.n58 185
R2933 VDD1.n57 VDD1.n23 185
R2934 VDD1.n27 VDD1.n24 185
R2935 VDD1.n52 VDD1.n51 185
R2936 VDD1.n50 VDD1.n49 185
R2937 VDD1.n29 VDD1.n28 185
R2938 VDD1.n44 VDD1.n43 185
R2939 VDD1.n42 VDD1.n41 185
R2940 VDD1.n33 VDD1.n32 185
R2941 VDD1.n36 VDD1.n35 185
R2942 VDD1.n140 VDD1.n139 185
R2943 VDD1.n137 VDD1.n136 185
R2944 VDD1.n146 VDD1.n145 185
R2945 VDD1.n148 VDD1.n147 185
R2946 VDD1.n133 VDD1.n132 185
R2947 VDD1.n154 VDD1.n153 185
R2948 VDD1.n157 VDD1.n156 185
R2949 VDD1.n155 VDD1.n129 185
R2950 VDD1.n162 VDD1.n128 185
R2951 VDD1.n164 VDD1.n163 185
R2952 VDD1.n166 VDD1.n165 185
R2953 VDD1.n125 VDD1.n124 185
R2954 VDD1.n172 VDD1.n171 185
R2955 VDD1.n174 VDD1.n173 185
R2956 VDD1.n121 VDD1.n120 185
R2957 VDD1.n180 VDD1.n179 185
R2958 VDD1.n182 VDD1.n181 185
R2959 VDD1.n117 VDD1.n116 185
R2960 VDD1.n188 VDD1.n187 185
R2961 VDD1.n190 VDD1.n189 185
R2962 VDD1.n113 VDD1.n112 185
R2963 VDD1.n196 VDD1.n195 185
R2964 VDD1.n198 VDD1.n197 185
R2965 VDD1.n109 VDD1.n108 185
R2966 VDD1.n204 VDD1.n203 185
R2967 VDD1.n206 VDD1.n205 185
R2968 VDD1.t5 VDD1.n34 149.524
R2969 VDD1.t0 VDD1.n138 149.524
R2970 VDD1.n100 VDD1.n99 104.615
R2971 VDD1.n99 VDD1.n3 104.615
R2972 VDD1.n92 VDD1.n3 104.615
R2973 VDD1.n92 VDD1.n91 104.615
R2974 VDD1.n91 VDD1.n7 104.615
R2975 VDD1.n84 VDD1.n7 104.615
R2976 VDD1.n84 VDD1.n83 104.615
R2977 VDD1.n83 VDD1.n11 104.615
R2978 VDD1.n76 VDD1.n11 104.615
R2979 VDD1.n76 VDD1.n75 104.615
R2980 VDD1.n75 VDD1.n15 104.615
R2981 VDD1.n68 VDD1.n15 104.615
R2982 VDD1.n68 VDD1.n67 104.615
R2983 VDD1.n67 VDD1.n19 104.615
R2984 VDD1.n60 VDD1.n19 104.615
R2985 VDD1.n60 VDD1.n59 104.615
R2986 VDD1.n59 VDD1.n23 104.615
R2987 VDD1.n27 VDD1.n23 104.615
R2988 VDD1.n51 VDD1.n27 104.615
R2989 VDD1.n51 VDD1.n50 104.615
R2990 VDD1.n50 VDD1.n28 104.615
R2991 VDD1.n43 VDD1.n28 104.615
R2992 VDD1.n43 VDD1.n42 104.615
R2993 VDD1.n42 VDD1.n32 104.615
R2994 VDD1.n35 VDD1.n32 104.615
R2995 VDD1.n139 VDD1.n136 104.615
R2996 VDD1.n146 VDD1.n136 104.615
R2997 VDD1.n147 VDD1.n146 104.615
R2998 VDD1.n147 VDD1.n132 104.615
R2999 VDD1.n154 VDD1.n132 104.615
R3000 VDD1.n156 VDD1.n154 104.615
R3001 VDD1.n156 VDD1.n155 104.615
R3002 VDD1.n155 VDD1.n128 104.615
R3003 VDD1.n164 VDD1.n128 104.615
R3004 VDD1.n165 VDD1.n164 104.615
R3005 VDD1.n165 VDD1.n124 104.615
R3006 VDD1.n172 VDD1.n124 104.615
R3007 VDD1.n173 VDD1.n172 104.615
R3008 VDD1.n173 VDD1.n120 104.615
R3009 VDD1.n180 VDD1.n120 104.615
R3010 VDD1.n181 VDD1.n180 104.615
R3011 VDD1.n181 VDD1.n116 104.615
R3012 VDD1.n188 VDD1.n116 104.615
R3013 VDD1.n189 VDD1.n188 104.615
R3014 VDD1.n189 VDD1.n112 104.615
R3015 VDD1.n196 VDD1.n112 104.615
R3016 VDD1.n197 VDD1.n196 104.615
R3017 VDD1.n197 VDD1.n108 104.615
R3018 VDD1.n204 VDD1.n108 104.615
R3019 VDD1.n205 VDD1.n204 104.615
R3020 VDD1.n211 VDD1.n210 64.5768
R3021 VDD1.n213 VDD1.n212 64.0804
R3022 VDD1 VDD1.n104 54.4563
R3023 VDD1.n211 VDD1.n209 54.3428
R3024 VDD1.n35 VDD1.t5 52.3082
R3025 VDD1.n139 VDD1.t0 52.3082
R3026 VDD1.n213 VDD1.n211 49.4018
R3027 VDD1.n58 VDD1.n57 13.1884
R3028 VDD1.n163 VDD1.n162 13.1884
R3029 VDD1.n102 VDD1.n101 12.8005
R3030 VDD1.n61 VDD1.n22 12.8005
R3031 VDD1.n56 VDD1.n24 12.8005
R3032 VDD1.n161 VDD1.n129 12.8005
R3033 VDD1.n166 VDD1.n127 12.8005
R3034 VDD1.n207 VDD1.n206 12.8005
R3035 VDD1.n98 VDD1.n2 12.0247
R3036 VDD1.n62 VDD1.n20 12.0247
R3037 VDD1.n53 VDD1.n52 12.0247
R3038 VDD1.n158 VDD1.n157 12.0247
R3039 VDD1.n167 VDD1.n125 12.0247
R3040 VDD1.n203 VDD1.n107 12.0247
R3041 VDD1.n97 VDD1.n4 11.249
R3042 VDD1.n66 VDD1.n65 11.249
R3043 VDD1.n49 VDD1.n26 11.249
R3044 VDD1.n153 VDD1.n131 11.249
R3045 VDD1.n171 VDD1.n170 11.249
R3046 VDD1.n202 VDD1.n109 11.249
R3047 VDD1.n94 VDD1.n93 10.4732
R3048 VDD1.n69 VDD1.n18 10.4732
R3049 VDD1.n48 VDD1.n29 10.4732
R3050 VDD1.n152 VDD1.n133 10.4732
R3051 VDD1.n174 VDD1.n123 10.4732
R3052 VDD1.n199 VDD1.n198 10.4732
R3053 VDD1.n36 VDD1.n34 10.2747
R3054 VDD1.n140 VDD1.n138 10.2747
R3055 VDD1.n90 VDD1.n6 9.69747
R3056 VDD1.n70 VDD1.n16 9.69747
R3057 VDD1.n45 VDD1.n44 9.69747
R3058 VDD1.n149 VDD1.n148 9.69747
R3059 VDD1.n175 VDD1.n121 9.69747
R3060 VDD1.n195 VDD1.n111 9.69747
R3061 VDD1.n104 VDD1.n103 9.45567
R3062 VDD1.n209 VDD1.n208 9.45567
R3063 VDD1.n38 VDD1.n37 9.3005
R3064 VDD1.n40 VDD1.n39 9.3005
R3065 VDD1.n31 VDD1.n30 9.3005
R3066 VDD1.n46 VDD1.n45 9.3005
R3067 VDD1.n48 VDD1.n47 9.3005
R3068 VDD1.n26 VDD1.n25 9.3005
R3069 VDD1.n54 VDD1.n53 9.3005
R3070 VDD1.n56 VDD1.n55 9.3005
R3071 VDD1.n10 VDD1.n9 9.3005
R3072 VDD1.n87 VDD1.n86 9.3005
R3073 VDD1.n89 VDD1.n88 9.3005
R3074 VDD1.n6 VDD1.n5 9.3005
R3075 VDD1.n95 VDD1.n94 9.3005
R3076 VDD1.n97 VDD1.n96 9.3005
R3077 VDD1.n2 VDD1.n1 9.3005
R3078 VDD1.n103 VDD1.n102 9.3005
R3079 VDD1.n81 VDD1.n80 9.3005
R3080 VDD1.n79 VDD1.n78 9.3005
R3081 VDD1.n14 VDD1.n13 9.3005
R3082 VDD1.n73 VDD1.n72 9.3005
R3083 VDD1.n71 VDD1.n70 9.3005
R3084 VDD1.n18 VDD1.n17 9.3005
R3085 VDD1.n65 VDD1.n64 9.3005
R3086 VDD1.n63 VDD1.n62 9.3005
R3087 VDD1.n22 VDD1.n21 9.3005
R3088 VDD1.n184 VDD1.n183 9.3005
R3089 VDD1.n119 VDD1.n118 9.3005
R3090 VDD1.n178 VDD1.n177 9.3005
R3091 VDD1.n176 VDD1.n175 9.3005
R3092 VDD1.n123 VDD1.n122 9.3005
R3093 VDD1.n170 VDD1.n169 9.3005
R3094 VDD1.n168 VDD1.n167 9.3005
R3095 VDD1.n127 VDD1.n126 9.3005
R3096 VDD1.n142 VDD1.n141 9.3005
R3097 VDD1.n144 VDD1.n143 9.3005
R3098 VDD1.n135 VDD1.n134 9.3005
R3099 VDD1.n150 VDD1.n149 9.3005
R3100 VDD1.n152 VDD1.n151 9.3005
R3101 VDD1.n131 VDD1.n130 9.3005
R3102 VDD1.n159 VDD1.n158 9.3005
R3103 VDD1.n161 VDD1.n160 9.3005
R3104 VDD1.n186 VDD1.n185 9.3005
R3105 VDD1.n115 VDD1.n114 9.3005
R3106 VDD1.n192 VDD1.n191 9.3005
R3107 VDD1.n194 VDD1.n193 9.3005
R3108 VDD1.n111 VDD1.n110 9.3005
R3109 VDD1.n200 VDD1.n199 9.3005
R3110 VDD1.n202 VDD1.n201 9.3005
R3111 VDD1.n107 VDD1.n106 9.3005
R3112 VDD1.n208 VDD1.n207 9.3005
R3113 VDD1.n89 VDD1.n8 8.92171
R3114 VDD1.n74 VDD1.n73 8.92171
R3115 VDD1.n41 VDD1.n31 8.92171
R3116 VDD1.n145 VDD1.n135 8.92171
R3117 VDD1.n179 VDD1.n178 8.92171
R3118 VDD1.n194 VDD1.n113 8.92171
R3119 VDD1.n104 VDD1.n0 8.2187
R3120 VDD1.n209 VDD1.n105 8.2187
R3121 VDD1.n86 VDD1.n85 8.14595
R3122 VDD1.n77 VDD1.n14 8.14595
R3123 VDD1.n40 VDD1.n33 8.14595
R3124 VDD1.n144 VDD1.n137 8.14595
R3125 VDD1.n182 VDD1.n119 8.14595
R3126 VDD1.n191 VDD1.n190 8.14595
R3127 VDD1.n82 VDD1.n10 7.3702
R3128 VDD1.n78 VDD1.n12 7.3702
R3129 VDD1.n37 VDD1.n36 7.3702
R3130 VDD1.n141 VDD1.n140 7.3702
R3131 VDD1.n183 VDD1.n117 7.3702
R3132 VDD1.n187 VDD1.n115 7.3702
R3133 VDD1.n82 VDD1.n81 6.59444
R3134 VDD1.n81 VDD1.n12 6.59444
R3135 VDD1.n186 VDD1.n117 6.59444
R3136 VDD1.n187 VDD1.n186 6.59444
R3137 VDD1.n85 VDD1.n10 5.81868
R3138 VDD1.n78 VDD1.n77 5.81868
R3139 VDD1.n37 VDD1.n33 5.81868
R3140 VDD1.n141 VDD1.n137 5.81868
R3141 VDD1.n183 VDD1.n182 5.81868
R3142 VDD1.n190 VDD1.n115 5.81868
R3143 VDD1.n102 VDD1.n0 5.3904
R3144 VDD1.n207 VDD1.n105 5.3904
R3145 VDD1.n86 VDD1.n8 5.04292
R3146 VDD1.n74 VDD1.n14 5.04292
R3147 VDD1.n41 VDD1.n40 5.04292
R3148 VDD1.n145 VDD1.n144 5.04292
R3149 VDD1.n179 VDD1.n119 5.04292
R3150 VDD1.n191 VDD1.n113 5.04292
R3151 VDD1.n90 VDD1.n89 4.26717
R3152 VDD1.n73 VDD1.n16 4.26717
R3153 VDD1.n44 VDD1.n31 4.26717
R3154 VDD1.n148 VDD1.n135 4.26717
R3155 VDD1.n178 VDD1.n121 4.26717
R3156 VDD1.n195 VDD1.n194 4.26717
R3157 VDD1.n93 VDD1.n6 3.49141
R3158 VDD1.n70 VDD1.n69 3.49141
R3159 VDD1.n45 VDD1.n29 3.49141
R3160 VDD1.n149 VDD1.n133 3.49141
R3161 VDD1.n175 VDD1.n174 3.49141
R3162 VDD1.n198 VDD1.n111 3.49141
R3163 VDD1.n142 VDD1.n138 2.84303
R3164 VDD1.n38 VDD1.n34 2.84303
R3165 VDD1.n94 VDD1.n4 2.71565
R3166 VDD1.n66 VDD1.n18 2.71565
R3167 VDD1.n49 VDD1.n48 2.71565
R3168 VDD1.n153 VDD1.n152 2.71565
R3169 VDD1.n171 VDD1.n123 2.71565
R3170 VDD1.n199 VDD1.n109 2.71565
R3171 VDD1.n98 VDD1.n97 1.93989
R3172 VDD1.n65 VDD1.n20 1.93989
R3173 VDD1.n52 VDD1.n26 1.93989
R3174 VDD1.n157 VDD1.n131 1.93989
R3175 VDD1.n170 VDD1.n125 1.93989
R3176 VDD1.n203 VDD1.n202 1.93989
R3177 VDD1.n101 VDD1.n2 1.16414
R3178 VDD1.n62 VDD1.n61 1.16414
R3179 VDD1.n53 VDD1.n24 1.16414
R3180 VDD1.n158 VDD1.n129 1.16414
R3181 VDD1.n167 VDD1.n166 1.16414
R3182 VDD1.n206 VDD1.n107 1.16414
R3183 VDD1.n212 VDD1.t1 1.01484
R3184 VDD1.n212 VDD1.t3 1.01484
R3185 VDD1.n210 VDD1.t4 1.01484
R3186 VDD1.n210 VDD1.t2 1.01484
R3187 VDD1 VDD1.n213 0.494034
R3188 VDD1.n58 VDD1.n22 0.388379
R3189 VDD1.n57 VDD1.n56 0.388379
R3190 VDD1.n162 VDD1.n161 0.388379
R3191 VDD1.n163 VDD1.n127 0.388379
R3192 VDD1.n103 VDD1.n1 0.155672
R3193 VDD1.n96 VDD1.n1 0.155672
R3194 VDD1.n96 VDD1.n95 0.155672
R3195 VDD1.n95 VDD1.n5 0.155672
R3196 VDD1.n88 VDD1.n5 0.155672
R3197 VDD1.n88 VDD1.n87 0.155672
R3198 VDD1.n87 VDD1.n9 0.155672
R3199 VDD1.n80 VDD1.n9 0.155672
R3200 VDD1.n80 VDD1.n79 0.155672
R3201 VDD1.n79 VDD1.n13 0.155672
R3202 VDD1.n72 VDD1.n13 0.155672
R3203 VDD1.n72 VDD1.n71 0.155672
R3204 VDD1.n71 VDD1.n17 0.155672
R3205 VDD1.n64 VDD1.n17 0.155672
R3206 VDD1.n64 VDD1.n63 0.155672
R3207 VDD1.n63 VDD1.n21 0.155672
R3208 VDD1.n55 VDD1.n21 0.155672
R3209 VDD1.n55 VDD1.n54 0.155672
R3210 VDD1.n54 VDD1.n25 0.155672
R3211 VDD1.n47 VDD1.n25 0.155672
R3212 VDD1.n47 VDD1.n46 0.155672
R3213 VDD1.n46 VDD1.n30 0.155672
R3214 VDD1.n39 VDD1.n30 0.155672
R3215 VDD1.n39 VDD1.n38 0.155672
R3216 VDD1.n143 VDD1.n142 0.155672
R3217 VDD1.n143 VDD1.n134 0.155672
R3218 VDD1.n150 VDD1.n134 0.155672
R3219 VDD1.n151 VDD1.n150 0.155672
R3220 VDD1.n151 VDD1.n130 0.155672
R3221 VDD1.n159 VDD1.n130 0.155672
R3222 VDD1.n160 VDD1.n159 0.155672
R3223 VDD1.n160 VDD1.n126 0.155672
R3224 VDD1.n168 VDD1.n126 0.155672
R3225 VDD1.n169 VDD1.n168 0.155672
R3226 VDD1.n169 VDD1.n122 0.155672
R3227 VDD1.n176 VDD1.n122 0.155672
R3228 VDD1.n177 VDD1.n176 0.155672
R3229 VDD1.n177 VDD1.n118 0.155672
R3230 VDD1.n184 VDD1.n118 0.155672
R3231 VDD1.n185 VDD1.n184 0.155672
R3232 VDD1.n185 VDD1.n114 0.155672
R3233 VDD1.n192 VDD1.n114 0.155672
R3234 VDD1.n193 VDD1.n192 0.155672
R3235 VDD1.n193 VDD1.n110 0.155672
R3236 VDD1.n200 VDD1.n110 0.155672
R3237 VDD1.n201 VDD1.n200 0.155672
R3238 VDD1.n201 VDD1.n106 0.155672
R3239 VDD1.n208 VDD1.n106 0.155672
C0 VTAIL VDD1 10.598401f
C1 VTAIL VDD2 10.6443f
C2 VDD1 VDD2 1.26272f
C3 VP VN 7.95639f
C4 VP VTAIL 10.1313f
C5 VN VTAIL 10.116799f
C6 VP VDD1 10.642799f
C7 VP VDD2 0.427803f
C8 VN VDD1 0.150396f
C9 VN VDD2 10.3701f
C10 VDD2 B 7.037685f
C11 VDD1 B 7.154613f
C12 VTAIL B 10.542236f
C13 VN B 12.50609f
C14 VP B 10.905023f
C15 VDD1.n0 B 0.029838f
C16 VDD1.n1 B 0.021349f
C17 VDD1.n2 B 0.011472f
C18 VDD1.n3 B 0.027116f
C19 VDD1.n4 B 0.012147f
C20 VDD1.n5 B 0.021349f
C21 VDD1.n6 B 0.011472f
C22 VDD1.n7 B 0.027116f
C23 VDD1.n8 B 0.012147f
C24 VDD1.n9 B 0.021349f
C25 VDD1.n10 B 0.011472f
C26 VDD1.n11 B 0.027116f
C27 VDD1.n12 B 0.012147f
C28 VDD1.n13 B 0.021349f
C29 VDD1.n14 B 0.011472f
C30 VDD1.n15 B 0.027116f
C31 VDD1.n16 B 0.012147f
C32 VDD1.n17 B 0.021349f
C33 VDD1.n18 B 0.011472f
C34 VDD1.n19 B 0.027116f
C35 VDD1.n20 B 0.012147f
C36 VDD1.n21 B 0.021349f
C37 VDD1.n22 B 0.011472f
C38 VDD1.n23 B 0.027116f
C39 VDD1.n24 B 0.012147f
C40 VDD1.n25 B 0.021349f
C41 VDD1.n26 B 0.011472f
C42 VDD1.n27 B 0.027116f
C43 VDD1.n28 B 0.027116f
C44 VDD1.n29 B 0.012147f
C45 VDD1.n30 B 0.021349f
C46 VDD1.n31 B 0.011472f
C47 VDD1.n32 B 0.027116f
C48 VDD1.n33 B 0.012147f
C49 VDD1.n34 B 0.21556f
C50 VDD1.t5 B 0.046661f
C51 VDD1.n35 B 0.020337f
C52 VDD1.n36 B 0.019169f
C53 VDD1.n37 B 0.011472f
C54 VDD1.n38 B 1.7911f
C55 VDD1.n39 B 0.021349f
C56 VDD1.n40 B 0.011472f
C57 VDD1.n41 B 0.012147f
C58 VDD1.n42 B 0.027116f
C59 VDD1.n43 B 0.027116f
C60 VDD1.n44 B 0.012147f
C61 VDD1.n45 B 0.011472f
C62 VDD1.n46 B 0.021349f
C63 VDD1.n47 B 0.021349f
C64 VDD1.n48 B 0.011472f
C65 VDD1.n49 B 0.012147f
C66 VDD1.n50 B 0.027116f
C67 VDD1.n51 B 0.027116f
C68 VDD1.n52 B 0.012147f
C69 VDD1.n53 B 0.011472f
C70 VDD1.n54 B 0.021349f
C71 VDD1.n55 B 0.021349f
C72 VDD1.n56 B 0.011472f
C73 VDD1.n57 B 0.011809f
C74 VDD1.n58 B 0.011809f
C75 VDD1.n59 B 0.027116f
C76 VDD1.n60 B 0.027116f
C77 VDD1.n61 B 0.012147f
C78 VDD1.n62 B 0.011472f
C79 VDD1.n63 B 0.021349f
C80 VDD1.n64 B 0.021349f
C81 VDD1.n65 B 0.011472f
C82 VDD1.n66 B 0.012147f
C83 VDD1.n67 B 0.027116f
C84 VDD1.n68 B 0.027116f
C85 VDD1.n69 B 0.012147f
C86 VDD1.n70 B 0.011472f
C87 VDD1.n71 B 0.021349f
C88 VDD1.n72 B 0.021349f
C89 VDD1.n73 B 0.011472f
C90 VDD1.n74 B 0.012147f
C91 VDD1.n75 B 0.027116f
C92 VDD1.n76 B 0.027116f
C93 VDD1.n77 B 0.012147f
C94 VDD1.n78 B 0.011472f
C95 VDD1.n79 B 0.021349f
C96 VDD1.n80 B 0.021349f
C97 VDD1.n81 B 0.011472f
C98 VDD1.n82 B 0.012147f
C99 VDD1.n83 B 0.027116f
C100 VDD1.n84 B 0.027116f
C101 VDD1.n85 B 0.012147f
C102 VDD1.n86 B 0.011472f
C103 VDD1.n87 B 0.021349f
C104 VDD1.n88 B 0.021349f
C105 VDD1.n89 B 0.011472f
C106 VDD1.n90 B 0.012147f
C107 VDD1.n91 B 0.027116f
C108 VDD1.n92 B 0.027116f
C109 VDD1.n93 B 0.012147f
C110 VDD1.n94 B 0.011472f
C111 VDD1.n95 B 0.021349f
C112 VDD1.n96 B 0.021349f
C113 VDD1.n97 B 0.011472f
C114 VDD1.n98 B 0.012147f
C115 VDD1.n99 B 0.027116f
C116 VDD1.n100 B 0.056137f
C117 VDD1.n101 B 0.012147f
C118 VDD1.n102 B 0.022432f
C119 VDD1.n103 B 0.05518f
C120 VDD1.n104 B 0.078646f
C121 VDD1.n105 B 0.029838f
C122 VDD1.n106 B 0.021349f
C123 VDD1.n107 B 0.011472f
C124 VDD1.n108 B 0.027116f
C125 VDD1.n109 B 0.012147f
C126 VDD1.n110 B 0.021349f
C127 VDD1.n111 B 0.011472f
C128 VDD1.n112 B 0.027116f
C129 VDD1.n113 B 0.012147f
C130 VDD1.n114 B 0.021349f
C131 VDD1.n115 B 0.011472f
C132 VDD1.n116 B 0.027116f
C133 VDD1.n117 B 0.012147f
C134 VDD1.n118 B 0.021349f
C135 VDD1.n119 B 0.011472f
C136 VDD1.n120 B 0.027116f
C137 VDD1.n121 B 0.012147f
C138 VDD1.n122 B 0.021349f
C139 VDD1.n123 B 0.011472f
C140 VDD1.n124 B 0.027116f
C141 VDD1.n125 B 0.012147f
C142 VDD1.n126 B 0.021349f
C143 VDD1.n127 B 0.011472f
C144 VDD1.n128 B 0.027116f
C145 VDD1.n129 B 0.012147f
C146 VDD1.n130 B 0.021349f
C147 VDD1.n131 B 0.011472f
C148 VDD1.n132 B 0.027116f
C149 VDD1.n133 B 0.012147f
C150 VDD1.n134 B 0.021349f
C151 VDD1.n135 B 0.011472f
C152 VDD1.n136 B 0.027116f
C153 VDD1.n137 B 0.012147f
C154 VDD1.n138 B 0.21556f
C155 VDD1.t0 B 0.046661f
C156 VDD1.n139 B 0.020337f
C157 VDD1.n140 B 0.019169f
C158 VDD1.n141 B 0.011472f
C159 VDD1.n142 B 1.7911f
C160 VDD1.n143 B 0.021349f
C161 VDD1.n144 B 0.011472f
C162 VDD1.n145 B 0.012147f
C163 VDD1.n146 B 0.027116f
C164 VDD1.n147 B 0.027116f
C165 VDD1.n148 B 0.012147f
C166 VDD1.n149 B 0.011472f
C167 VDD1.n150 B 0.021349f
C168 VDD1.n151 B 0.021349f
C169 VDD1.n152 B 0.011472f
C170 VDD1.n153 B 0.012147f
C171 VDD1.n154 B 0.027116f
C172 VDD1.n155 B 0.027116f
C173 VDD1.n156 B 0.027116f
C174 VDD1.n157 B 0.012147f
C175 VDD1.n158 B 0.011472f
C176 VDD1.n159 B 0.021349f
C177 VDD1.n160 B 0.021349f
C178 VDD1.n161 B 0.011472f
C179 VDD1.n162 B 0.011809f
C180 VDD1.n163 B 0.011809f
C181 VDD1.n164 B 0.027116f
C182 VDD1.n165 B 0.027116f
C183 VDD1.n166 B 0.012147f
C184 VDD1.n167 B 0.011472f
C185 VDD1.n168 B 0.021349f
C186 VDD1.n169 B 0.021349f
C187 VDD1.n170 B 0.011472f
C188 VDD1.n171 B 0.012147f
C189 VDD1.n172 B 0.027116f
C190 VDD1.n173 B 0.027116f
C191 VDD1.n174 B 0.012147f
C192 VDD1.n175 B 0.011472f
C193 VDD1.n176 B 0.021349f
C194 VDD1.n177 B 0.021349f
C195 VDD1.n178 B 0.011472f
C196 VDD1.n179 B 0.012147f
C197 VDD1.n180 B 0.027116f
C198 VDD1.n181 B 0.027116f
C199 VDD1.n182 B 0.012147f
C200 VDD1.n183 B 0.011472f
C201 VDD1.n184 B 0.021349f
C202 VDD1.n185 B 0.021349f
C203 VDD1.n186 B 0.011472f
C204 VDD1.n187 B 0.012147f
C205 VDD1.n188 B 0.027116f
C206 VDD1.n189 B 0.027116f
C207 VDD1.n190 B 0.012147f
C208 VDD1.n191 B 0.011472f
C209 VDD1.n192 B 0.021349f
C210 VDD1.n193 B 0.021349f
C211 VDD1.n194 B 0.011472f
C212 VDD1.n195 B 0.012147f
C213 VDD1.n196 B 0.027116f
C214 VDD1.n197 B 0.027116f
C215 VDD1.n198 B 0.012147f
C216 VDD1.n199 B 0.011472f
C217 VDD1.n200 B 0.021349f
C218 VDD1.n201 B 0.021349f
C219 VDD1.n202 B 0.011472f
C220 VDD1.n203 B 0.012147f
C221 VDD1.n204 B 0.027116f
C222 VDD1.n205 B 0.056137f
C223 VDD1.n206 B 0.012147f
C224 VDD1.n207 B 0.022432f
C225 VDD1.n208 B 0.05518f
C226 VDD1.n209 B 0.078097f
C227 VDD1.t4 B 0.329315f
C228 VDD1.t2 B 0.329315f
C229 VDD1.n210 B 3.02012f
C230 VDD1.n211 B 2.65204f
C231 VDD1.t1 B 0.329315f
C232 VDD1.t3 B 0.329315f
C233 VDD1.n212 B 3.0173f
C234 VDD1.n213 B 2.77442f
C235 VP.n0 B 0.032632f
C236 VP.t3 B 2.96803f
C237 VP.n1 B 0.020277f
C238 VP.n2 B 0.024753f
C239 VP.t1 B 2.96803f
C240 VP.n3 B 0.049521f
C241 VP.n4 B 0.024753f
C242 VP.t5 B 2.96803f
C243 VP.n5 B 1.10629f
C244 VP.n6 B 0.032632f
C245 VP.t2 B 2.96803f
C246 VP.n7 B 0.020277f
C247 VP.n8 B 0.211474f
C248 VP.t4 B 2.96803f
C249 VP.t0 B 3.12505f
C250 VP.n9 B 1.08341f
C251 VP.n10 B 1.09319f
C252 VP.n11 B 0.034571f
C253 VP.n12 B 0.049521f
C254 VP.n13 B 0.024753f
C255 VP.n14 B 0.024753f
C256 VP.n15 B 0.024753f
C257 VP.n16 B 0.048068f
C258 VP.n17 B 0.037291f
C259 VP.n18 B 1.10629f
C260 VP.n19 B 1.48949f
C261 VP.n20 B 1.50634f
C262 VP.n21 B 0.032632f
C263 VP.n22 B 0.037291f
C264 VP.n23 B 0.048068f
C265 VP.n24 B 0.020277f
C266 VP.n25 B 0.024753f
C267 VP.n26 B 0.024753f
C268 VP.n27 B 0.024753f
C269 VP.n28 B 0.034571f
C270 VP.n29 B 1.02919f
C271 VP.n30 B 0.034571f
C272 VP.n31 B 0.049521f
C273 VP.n32 B 0.024753f
C274 VP.n33 B 0.024753f
C275 VP.n34 B 0.024753f
C276 VP.n35 B 0.048068f
C277 VP.n36 B 0.037291f
C278 VP.n37 B 1.10629f
C279 VP.n38 B 0.034363f
C280 VTAIL.t6 B 0.342158f
C281 VTAIL.t9 B 0.342158f
C282 VTAIL.n0 B 3.07413f
C283 VTAIL.n1 B 0.36389f
C284 VTAIL.n2 B 0.031001f
C285 VTAIL.n3 B 0.022182f
C286 VTAIL.n4 B 0.011919f
C287 VTAIL.n5 B 0.028173f
C288 VTAIL.n6 B 0.012621f
C289 VTAIL.n7 B 0.022182f
C290 VTAIL.n8 B 0.011919f
C291 VTAIL.n9 B 0.028173f
C292 VTAIL.n10 B 0.012621f
C293 VTAIL.n11 B 0.022182f
C294 VTAIL.n12 B 0.011919f
C295 VTAIL.n13 B 0.028173f
C296 VTAIL.n14 B 0.012621f
C297 VTAIL.n15 B 0.022182f
C298 VTAIL.n16 B 0.011919f
C299 VTAIL.n17 B 0.028173f
C300 VTAIL.n18 B 0.012621f
C301 VTAIL.n19 B 0.022182f
C302 VTAIL.n20 B 0.011919f
C303 VTAIL.n21 B 0.028173f
C304 VTAIL.n22 B 0.012621f
C305 VTAIL.n23 B 0.022182f
C306 VTAIL.n24 B 0.011919f
C307 VTAIL.n25 B 0.028173f
C308 VTAIL.n26 B 0.012621f
C309 VTAIL.n27 B 0.022182f
C310 VTAIL.n28 B 0.011919f
C311 VTAIL.n29 B 0.028173f
C312 VTAIL.n30 B 0.012621f
C313 VTAIL.n31 B 0.022182f
C314 VTAIL.n32 B 0.011919f
C315 VTAIL.n33 B 0.028173f
C316 VTAIL.n34 B 0.012621f
C317 VTAIL.n35 B 0.223967f
C318 VTAIL.t3 B 0.048481f
C319 VTAIL.n36 B 0.02113f
C320 VTAIL.n37 B 0.019916f
C321 VTAIL.n38 B 0.011919f
C322 VTAIL.n39 B 1.86095f
C323 VTAIL.n40 B 0.022182f
C324 VTAIL.n41 B 0.011919f
C325 VTAIL.n42 B 0.012621f
C326 VTAIL.n43 B 0.028173f
C327 VTAIL.n44 B 0.028173f
C328 VTAIL.n45 B 0.012621f
C329 VTAIL.n46 B 0.011919f
C330 VTAIL.n47 B 0.022182f
C331 VTAIL.n48 B 0.022182f
C332 VTAIL.n49 B 0.011919f
C333 VTAIL.n50 B 0.012621f
C334 VTAIL.n51 B 0.028173f
C335 VTAIL.n52 B 0.028173f
C336 VTAIL.n53 B 0.028173f
C337 VTAIL.n54 B 0.012621f
C338 VTAIL.n55 B 0.011919f
C339 VTAIL.n56 B 0.022182f
C340 VTAIL.n57 B 0.022182f
C341 VTAIL.n58 B 0.011919f
C342 VTAIL.n59 B 0.01227f
C343 VTAIL.n60 B 0.01227f
C344 VTAIL.n61 B 0.028173f
C345 VTAIL.n62 B 0.028173f
C346 VTAIL.n63 B 0.012621f
C347 VTAIL.n64 B 0.011919f
C348 VTAIL.n65 B 0.022182f
C349 VTAIL.n66 B 0.022182f
C350 VTAIL.n67 B 0.011919f
C351 VTAIL.n68 B 0.012621f
C352 VTAIL.n69 B 0.028173f
C353 VTAIL.n70 B 0.028173f
C354 VTAIL.n71 B 0.012621f
C355 VTAIL.n72 B 0.011919f
C356 VTAIL.n73 B 0.022182f
C357 VTAIL.n74 B 0.022182f
C358 VTAIL.n75 B 0.011919f
C359 VTAIL.n76 B 0.012621f
C360 VTAIL.n77 B 0.028173f
C361 VTAIL.n78 B 0.028173f
C362 VTAIL.n79 B 0.012621f
C363 VTAIL.n80 B 0.011919f
C364 VTAIL.n81 B 0.022182f
C365 VTAIL.n82 B 0.022182f
C366 VTAIL.n83 B 0.011919f
C367 VTAIL.n84 B 0.012621f
C368 VTAIL.n85 B 0.028173f
C369 VTAIL.n86 B 0.028173f
C370 VTAIL.n87 B 0.012621f
C371 VTAIL.n88 B 0.011919f
C372 VTAIL.n89 B 0.022182f
C373 VTAIL.n90 B 0.022182f
C374 VTAIL.n91 B 0.011919f
C375 VTAIL.n92 B 0.012621f
C376 VTAIL.n93 B 0.028173f
C377 VTAIL.n94 B 0.028173f
C378 VTAIL.n95 B 0.012621f
C379 VTAIL.n96 B 0.011919f
C380 VTAIL.n97 B 0.022182f
C381 VTAIL.n98 B 0.022182f
C382 VTAIL.n99 B 0.011919f
C383 VTAIL.n100 B 0.012621f
C384 VTAIL.n101 B 0.028173f
C385 VTAIL.n102 B 0.058326f
C386 VTAIL.n103 B 0.012621f
C387 VTAIL.n104 B 0.023306f
C388 VTAIL.n105 B 0.057332f
C389 VTAIL.n106 B 0.061133f
C390 VTAIL.n107 B 0.292559f
C391 VTAIL.t0 B 0.342158f
C392 VTAIL.t5 B 0.342158f
C393 VTAIL.n108 B 3.07413f
C394 VTAIL.n109 B 2.1851f
C395 VTAIL.t7 B 0.342158f
C396 VTAIL.t11 B 0.342158f
C397 VTAIL.n110 B 3.07414f
C398 VTAIL.n111 B 2.18509f
C399 VTAIL.n112 B 0.031001f
C400 VTAIL.n113 B 0.022182f
C401 VTAIL.n114 B 0.011919f
C402 VTAIL.n115 B 0.028173f
C403 VTAIL.n116 B 0.012621f
C404 VTAIL.n117 B 0.022182f
C405 VTAIL.n118 B 0.011919f
C406 VTAIL.n119 B 0.028173f
C407 VTAIL.n120 B 0.012621f
C408 VTAIL.n121 B 0.022182f
C409 VTAIL.n122 B 0.011919f
C410 VTAIL.n123 B 0.028173f
C411 VTAIL.n124 B 0.012621f
C412 VTAIL.n125 B 0.022182f
C413 VTAIL.n126 B 0.011919f
C414 VTAIL.n127 B 0.028173f
C415 VTAIL.n128 B 0.012621f
C416 VTAIL.n129 B 0.022182f
C417 VTAIL.n130 B 0.011919f
C418 VTAIL.n131 B 0.028173f
C419 VTAIL.n132 B 0.012621f
C420 VTAIL.n133 B 0.022182f
C421 VTAIL.n134 B 0.011919f
C422 VTAIL.n135 B 0.028173f
C423 VTAIL.n136 B 0.012621f
C424 VTAIL.n137 B 0.022182f
C425 VTAIL.n138 B 0.011919f
C426 VTAIL.n139 B 0.028173f
C427 VTAIL.n140 B 0.028173f
C428 VTAIL.n141 B 0.012621f
C429 VTAIL.n142 B 0.022182f
C430 VTAIL.n143 B 0.011919f
C431 VTAIL.n144 B 0.028173f
C432 VTAIL.n145 B 0.012621f
C433 VTAIL.n146 B 0.223967f
C434 VTAIL.t8 B 0.048481f
C435 VTAIL.n147 B 0.02113f
C436 VTAIL.n148 B 0.019916f
C437 VTAIL.n149 B 0.011919f
C438 VTAIL.n150 B 1.86095f
C439 VTAIL.n151 B 0.022182f
C440 VTAIL.n152 B 0.011919f
C441 VTAIL.n153 B 0.012621f
C442 VTAIL.n154 B 0.028173f
C443 VTAIL.n155 B 0.028173f
C444 VTAIL.n156 B 0.012621f
C445 VTAIL.n157 B 0.011919f
C446 VTAIL.n158 B 0.022182f
C447 VTAIL.n159 B 0.022182f
C448 VTAIL.n160 B 0.011919f
C449 VTAIL.n161 B 0.012621f
C450 VTAIL.n162 B 0.028173f
C451 VTAIL.n163 B 0.028173f
C452 VTAIL.n164 B 0.012621f
C453 VTAIL.n165 B 0.011919f
C454 VTAIL.n166 B 0.022182f
C455 VTAIL.n167 B 0.022182f
C456 VTAIL.n168 B 0.011919f
C457 VTAIL.n169 B 0.01227f
C458 VTAIL.n170 B 0.01227f
C459 VTAIL.n171 B 0.028173f
C460 VTAIL.n172 B 0.028173f
C461 VTAIL.n173 B 0.012621f
C462 VTAIL.n174 B 0.011919f
C463 VTAIL.n175 B 0.022182f
C464 VTAIL.n176 B 0.022182f
C465 VTAIL.n177 B 0.011919f
C466 VTAIL.n178 B 0.012621f
C467 VTAIL.n179 B 0.028173f
C468 VTAIL.n180 B 0.028173f
C469 VTAIL.n181 B 0.012621f
C470 VTAIL.n182 B 0.011919f
C471 VTAIL.n183 B 0.022182f
C472 VTAIL.n184 B 0.022182f
C473 VTAIL.n185 B 0.011919f
C474 VTAIL.n186 B 0.012621f
C475 VTAIL.n187 B 0.028173f
C476 VTAIL.n188 B 0.028173f
C477 VTAIL.n189 B 0.012621f
C478 VTAIL.n190 B 0.011919f
C479 VTAIL.n191 B 0.022182f
C480 VTAIL.n192 B 0.022182f
C481 VTAIL.n193 B 0.011919f
C482 VTAIL.n194 B 0.012621f
C483 VTAIL.n195 B 0.028173f
C484 VTAIL.n196 B 0.028173f
C485 VTAIL.n197 B 0.012621f
C486 VTAIL.n198 B 0.011919f
C487 VTAIL.n199 B 0.022182f
C488 VTAIL.n200 B 0.022182f
C489 VTAIL.n201 B 0.011919f
C490 VTAIL.n202 B 0.012621f
C491 VTAIL.n203 B 0.028173f
C492 VTAIL.n204 B 0.028173f
C493 VTAIL.n205 B 0.012621f
C494 VTAIL.n206 B 0.011919f
C495 VTAIL.n207 B 0.022182f
C496 VTAIL.n208 B 0.022182f
C497 VTAIL.n209 B 0.011919f
C498 VTAIL.n210 B 0.012621f
C499 VTAIL.n211 B 0.028173f
C500 VTAIL.n212 B 0.058326f
C501 VTAIL.n213 B 0.012621f
C502 VTAIL.n214 B 0.023306f
C503 VTAIL.n215 B 0.057332f
C504 VTAIL.n216 B 0.061133f
C505 VTAIL.n217 B 0.292559f
C506 VTAIL.t2 B 0.342158f
C507 VTAIL.t1 B 0.342158f
C508 VTAIL.n218 B 3.07414f
C509 VTAIL.n219 B 0.47802f
C510 VTAIL.n220 B 0.031001f
C511 VTAIL.n221 B 0.022182f
C512 VTAIL.n222 B 0.011919f
C513 VTAIL.n223 B 0.028173f
C514 VTAIL.n224 B 0.012621f
C515 VTAIL.n225 B 0.022182f
C516 VTAIL.n226 B 0.011919f
C517 VTAIL.n227 B 0.028173f
C518 VTAIL.n228 B 0.012621f
C519 VTAIL.n229 B 0.022182f
C520 VTAIL.n230 B 0.011919f
C521 VTAIL.n231 B 0.028173f
C522 VTAIL.n232 B 0.012621f
C523 VTAIL.n233 B 0.022182f
C524 VTAIL.n234 B 0.011919f
C525 VTAIL.n235 B 0.028173f
C526 VTAIL.n236 B 0.012621f
C527 VTAIL.n237 B 0.022182f
C528 VTAIL.n238 B 0.011919f
C529 VTAIL.n239 B 0.028173f
C530 VTAIL.n240 B 0.012621f
C531 VTAIL.n241 B 0.022182f
C532 VTAIL.n242 B 0.011919f
C533 VTAIL.n243 B 0.028173f
C534 VTAIL.n244 B 0.012621f
C535 VTAIL.n245 B 0.022182f
C536 VTAIL.n246 B 0.011919f
C537 VTAIL.n247 B 0.028173f
C538 VTAIL.n248 B 0.028173f
C539 VTAIL.n249 B 0.012621f
C540 VTAIL.n250 B 0.022182f
C541 VTAIL.n251 B 0.011919f
C542 VTAIL.n252 B 0.028173f
C543 VTAIL.n253 B 0.012621f
C544 VTAIL.n254 B 0.223967f
C545 VTAIL.t4 B 0.048481f
C546 VTAIL.n255 B 0.02113f
C547 VTAIL.n256 B 0.019916f
C548 VTAIL.n257 B 0.011919f
C549 VTAIL.n258 B 1.86095f
C550 VTAIL.n259 B 0.022182f
C551 VTAIL.n260 B 0.011919f
C552 VTAIL.n261 B 0.012621f
C553 VTAIL.n262 B 0.028173f
C554 VTAIL.n263 B 0.028173f
C555 VTAIL.n264 B 0.012621f
C556 VTAIL.n265 B 0.011919f
C557 VTAIL.n266 B 0.022182f
C558 VTAIL.n267 B 0.022182f
C559 VTAIL.n268 B 0.011919f
C560 VTAIL.n269 B 0.012621f
C561 VTAIL.n270 B 0.028173f
C562 VTAIL.n271 B 0.028173f
C563 VTAIL.n272 B 0.012621f
C564 VTAIL.n273 B 0.011919f
C565 VTAIL.n274 B 0.022182f
C566 VTAIL.n275 B 0.022182f
C567 VTAIL.n276 B 0.011919f
C568 VTAIL.n277 B 0.01227f
C569 VTAIL.n278 B 0.01227f
C570 VTAIL.n279 B 0.028173f
C571 VTAIL.n280 B 0.028173f
C572 VTAIL.n281 B 0.012621f
C573 VTAIL.n282 B 0.011919f
C574 VTAIL.n283 B 0.022182f
C575 VTAIL.n284 B 0.022182f
C576 VTAIL.n285 B 0.011919f
C577 VTAIL.n286 B 0.012621f
C578 VTAIL.n287 B 0.028173f
C579 VTAIL.n288 B 0.028173f
C580 VTAIL.n289 B 0.012621f
C581 VTAIL.n290 B 0.011919f
C582 VTAIL.n291 B 0.022182f
C583 VTAIL.n292 B 0.022182f
C584 VTAIL.n293 B 0.011919f
C585 VTAIL.n294 B 0.012621f
C586 VTAIL.n295 B 0.028173f
C587 VTAIL.n296 B 0.028173f
C588 VTAIL.n297 B 0.012621f
C589 VTAIL.n298 B 0.011919f
C590 VTAIL.n299 B 0.022182f
C591 VTAIL.n300 B 0.022182f
C592 VTAIL.n301 B 0.011919f
C593 VTAIL.n302 B 0.012621f
C594 VTAIL.n303 B 0.028173f
C595 VTAIL.n304 B 0.028173f
C596 VTAIL.n305 B 0.012621f
C597 VTAIL.n306 B 0.011919f
C598 VTAIL.n307 B 0.022182f
C599 VTAIL.n308 B 0.022182f
C600 VTAIL.n309 B 0.011919f
C601 VTAIL.n310 B 0.012621f
C602 VTAIL.n311 B 0.028173f
C603 VTAIL.n312 B 0.028173f
C604 VTAIL.n313 B 0.012621f
C605 VTAIL.n314 B 0.011919f
C606 VTAIL.n315 B 0.022182f
C607 VTAIL.n316 B 0.022182f
C608 VTAIL.n317 B 0.011919f
C609 VTAIL.n318 B 0.012621f
C610 VTAIL.n319 B 0.028173f
C611 VTAIL.n320 B 0.058326f
C612 VTAIL.n321 B 0.012621f
C613 VTAIL.n322 B 0.023306f
C614 VTAIL.n323 B 0.057332f
C615 VTAIL.n324 B 0.061133f
C616 VTAIL.n325 B 1.84189f
C617 VTAIL.n326 B 0.031001f
C618 VTAIL.n327 B 0.022182f
C619 VTAIL.n328 B 0.011919f
C620 VTAIL.n329 B 0.028173f
C621 VTAIL.n330 B 0.012621f
C622 VTAIL.n331 B 0.022182f
C623 VTAIL.n332 B 0.011919f
C624 VTAIL.n333 B 0.028173f
C625 VTAIL.n334 B 0.012621f
C626 VTAIL.n335 B 0.022182f
C627 VTAIL.n336 B 0.011919f
C628 VTAIL.n337 B 0.028173f
C629 VTAIL.n338 B 0.012621f
C630 VTAIL.n339 B 0.022182f
C631 VTAIL.n340 B 0.011919f
C632 VTAIL.n341 B 0.028173f
C633 VTAIL.n342 B 0.012621f
C634 VTAIL.n343 B 0.022182f
C635 VTAIL.n344 B 0.011919f
C636 VTAIL.n345 B 0.028173f
C637 VTAIL.n346 B 0.012621f
C638 VTAIL.n347 B 0.022182f
C639 VTAIL.n348 B 0.011919f
C640 VTAIL.n349 B 0.028173f
C641 VTAIL.n350 B 0.012621f
C642 VTAIL.n351 B 0.022182f
C643 VTAIL.n352 B 0.011919f
C644 VTAIL.n353 B 0.028173f
C645 VTAIL.n354 B 0.012621f
C646 VTAIL.n355 B 0.022182f
C647 VTAIL.n356 B 0.011919f
C648 VTAIL.n357 B 0.028173f
C649 VTAIL.n358 B 0.012621f
C650 VTAIL.n359 B 0.223967f
C651 VTAIL.t10 B 0.048481f
C652 VTAIL.n360 B 0.02113f
C653 VTAIL.n361 B 0.019916f
C654 VTAIL.n362 B 0.011919f
C655 VTAIL.n363 B 1.86095f
C656 VTAIL.n364 B 0.022182f
C657 VTAIL.n365 B 0.011919f
C658 VTAIL.n366 B 0.012621f
C659 VTAIL.n367 B 0.028173f
C660 VTAIL.n368 B 0.028173f
C661 VTAIL.n369 B 0.012621f
C662 VTAIL.n370 B 0.011919f
C663 VTAIL.n371 B 0.022182f
C664 VTAIL.n372 B 0.022182f
C665 VTAIL.n373 B 0.011919f
C666 VTAIL.n374 B 0.012621f
C667 VTAIL.n375 B 0.028173f
C668 VTAIL.n376 B 0.028173f
C669 VTAIL.n377 B 0.028173f
C670 VTAIL.n378 B 0.012621f
C671 VTAIL.n379 B 0.011919f
C672 VTAIL.n380 B 0.022182f
C673 VTAIL.n381 B 0.022182f
C674 VTAIL.n382 B 0.011919f
C675 VTAIL.n383 B 0.01227f
C676 VTAIL.n384 B 0.01227f
C677 VTAIL.n385 B 0.028173f
C678 VTAIL.n386 B 0.028173f
C679 VTAIL.n387 B 0.012621f
C680 VTAIL.n388 B 0.011919f
C681 VTAIL.n389 B 0.022182f
C682 VTAIL.n390 B 0.022182f
C683 VTAIL.n391 B 0.011919f
C684 VTAIL.n392 B 0.012621f
C685 VTAIL.n393 B 0.028173f
C686 VTAIL.n394 B 0.028173f
C687 VTAIL.n395 B 0.012621f
C688 VTAIL.n396 B 0.011919f
C689 VTAIL.n397 B 0.022182f
C690 VTAIL.n398 B 0.022182f
C691 VTAIL.n399 B 0.011919f
C692 VTAIL.n400 B 0.012621f
C693 VTAIL.n401 B 0.028173f
C694 VTAIL.n402 B 0.028173f
C695 VTAIL.n403 B 0.012621f
C696 VTAIL.n404 B 0.011919f
C697 VTAIL.n405 B 0.022182f
C698 VTAIL.n406 B 0.022182f
C699 VTAIL.n407 B 0.011919f
C700 VTAIL.n408 B 0.012621f
C701 VTAIL.n409 B 0.028173f
C702 VTAIL.n410 B 0.028173f
C703 VTAIL.n411 B 0.012621f
C704 VTAIL.n412 B 0.011919f
C705 VTAIL.n413 B 0.022182f
C706 VTAIL.n414 B 0.022182f
C707 VTAIL.n415 B 0.011919f
C708 VTAIL.n416 B 0.012621f
C709 VTAIL.n417 B 0.028173f
C710 VTAIL.n418 B 0.028173f
C711 VTAIL.n419 B 0.012621f
C712 VTAIL.n420 B 0.011919f
C713 VTAIL.n421 B 0.022182f
C714 VTAIL.n422 B 0.022182f
C715 VTAIL.n423 B 0.011919f
C716 VTAIL.n424 B 0.012621f
C717 VTAIL.n425 B 0.028173f
C718 VTAIL.n426 B 0.058326f
C719 VTAIL.n427 B 0.012621f
C720 VTAIL.n428 B 0.023306f
C721 VTAIL.n429 B 0.057332f
C722 VTAIL.n430 B 0.061133f
C723 VTAIL.n431 B 1.7983f
C724 VDD2.n0 B 0.029666f
C725 VDD2.n1 B 0.021227f
C726 VDD2.n2 B 0.011406f
C727 VDD2.n3 B 0.02696f
C728 VDD2.n4 B 0.012077f
C729 VDD2.n5 B 0.021227f
C730 VDD2.n6 B 0.011406f
C731 VDD2.n7 B 0.02696f
C732 VDD2.n8 B 0.012077f
C733 VDD2.n9 B 0.021227f
C734 VDD2.n10 B 0.011406f
C735 VDD2.n11 B 0.02696f
C736 VDD2.n12 B 0.012077f
C737 VDD2.n13 B 0.021227f
C738 VDD2.n14 B 0.011406f
C739 VDD2.n15 B 0.02696f
C740 VDD2.n16 B 0.012077f
C741 VDD2.n17 B 0.021227f
C742 VDD2.n18 B 0.011406f
C743 VDD2.n19 B 0.02696f
C744 VDD2.n20 B 0.012077f
C745 VDD2.n21 B 0.021227f
C746 VDD2.n22 B 0.011406f
C747 VDD2.n23 B 0.02696f
C748 VDD2.n24 B 0.012077f
C749 VDD2.n25 B 0.021227f
C750 VDD2.n26 B 0.011406f
C751 VDD2.n27 B 0.02696f
C752 VDD2.n28 B 0.012077f
C753 VDD2.n29 B 0.021227f
C754 VDD2.n30 B 0.011406f
C755 VDD2.n31 B 0.02696f
C756 VDD2.n32 B 0.012077f
C757 VDD2.n33 B 0.214324f
C758 VDD2.t2 B 0.046394f
C759 VDD2.n34 B 0.02022f
C760 VDD2.n35 B 0.019059f
C761 VDD2.n36 B 0.011406f
C762 VDD2.n37 B 1.78083f
C763 VDD2.n38 B 0.021227f
C764 VDD2.n39 B 0.011406f
C765 VDD2.n40 B 0.012077f
C766 VDD2.n41 B 0.02696f
C767 VDD2.n42 B 0.02696f
C768 VDD2.n43 B 0.012077f
C769 VDD2.n44 B 0.011406f
C770 VDD2.n45 B 0.021227f
C771 VDD2.n46 B 0.021227f
C772 VDD2.n47 B 0.011406f
C773 VDD2.n48 B 0.012077f
C774 VDD2.n49 B 0.02696f
C775 VDD2.n50 B 0.02696f
C776 VDD2.n51 B 0.02696f
C777 VDD2.n52 B 0.012077f
C778 VDD2.n53 B 0.011406f
C779 VDD2.n54 B 0.021227f
C780 VDD2.n55 B 0.021227f
C781 VDD2.n56 B 0.011406f
C782 VDD2.n57 B 0.011742f
C783 VDD2.n58 B 0.011742f
C784 VDD2.n59 B 0.02696f
C785 VDD2.n60 B 0.02696f
C786 VDD2.n61 B 0.012077f
C787 VDD2.n62 B 0.011406f
C788 VDD2.n63 B 0.021227f
C789 VDD2.n64 B 0.021227f
C790 VDD2.n65 B 0.011406f
C791 VDD2.n66 B 0.012077f
C792 VDD2.n67 B 0.02696f
C793 VDD2.n68 B 0.02696f
C794 VDD2.n69 B 0.012077f
C795 VDD2.n70 B 0.011406f
C796 VDD2.n71 B 0.021227f
C797 VDD2.n72 B 0.021227f
C798 VDD2.n73 B 0.011406f
C799 VDD2.n74 B 0.012077f
C800 VDD2.n75 B 0.02696f
C801 VDD2.n76 B 0.02696f
C802 VDD2.n77 B 0.012077f
C803 VDD2.n78 B 0.011406f
C804 VDD2.n79 B 0.021227f
C805 VDD2.n80 B 0.021227f
C806 VDD2.n81 B 0.011406f
C807 VDD2.n82 B 0.012077f
C808 VDD2.n83 B 0.02696f
C809 VDD2.n84 B 0.02696f
C810 VDD2.n85 B 0.012077f
C811 VDD2.n86 B 0.011406f
C812 VDD2.n87 B 0.021227f
C813 VDD2.n88 B 0.021227f
C814 VDD2.n89 B 0.011406f
C815 VDD2.n90 B 0.012077f
C816 VDD2.n91 B 0.02696f
C817 VDD2.n92 B 0.02696f
C818 VDD2.n93 B 0.012077f
C819 VDD2.n94 B 0.011406f
C820 VDD2.n95 B 0.021227f
C821 VDD2.n96 B 0.021227f
C822 VDD2.n97 B 0.011406f
C823 VDD2.n98 B 0.012077f
C824 VDD2.n99 B 0.02696f
C825 VDD2.n100 B 0.055815f
C826 VDD2.n101 B 0.012077f
C827 VDD2.n102 B 0.022303f
C828 VDD2.n103 B 0.054864f
C829 VDD2.n104 B 0.077649f
C830 VDD2.t1 B 0.327426f
C831 VDD2.t0 B 0.327426f
C832 VDD2.n105 B 3.00279f
C833 VDD2.n106 B 2.53586f
C834 VDD2.n107 B 0.029666f
C835 VDD2.n108 B 0.021227f
C836 VDD2.n109 B 0.011406f
C837 VDD2.n110 B 0.02696f
C838 VDD2.n111 B 0.012077f
C839 VDD2.n112 B 0.021227f
C840 VDD2.n113 B 0.011406f
C841 VDD2.n114 B 0.02696f
C842 VDD2.n115 B 0.012077f
C843 VDD2.n116 B 0.021227f
C844 VDD2.n117 B 0.011406f
C845 VDD2.n118 B 0.02696f
C846 VDD2.n119 B 0.012077f
C847 VDD2.n120 B 0.021227f
C848 VDD2.n121 B 0.011406f
C849 VDD2.n122 B 0.02696f
C850 VDD2.n123 B 0.012077f
C851 VDD2.n124 B 0.021227f
C852 VDD2.n125 B 0.011406f
C853 VDD2.n126 B 0.02696f
C854 VDD2.n127 B 0.012077f
C855 VDD2.n128 B 0.021227f
C856 VDD2.n129 B 0.011406f
C857 VDD2.n130 B 0.02696f
C858 VDD2.n131 B 0.012077f
C859 VDD2.n132 B 0.021227f
C860 VDD2.n133 B 0.011406f
C861 VDD2.n134 B 0.02696f
C862 VDD2.n135 B 0.02696f
C863 VDD2.n136 B 0.012077f
C864 VDD2.n137 B 0.021227f
C865 VDD2.n138 B 0.011406f
C866 VDD2.n139 B 0.02696f
C867 VDD2.n140 B 0.012077f
C868 VDD2.n141 B 0.214324f
C869 VDD2.t5 B 0.046394f
C870 VDD2.n142 B 0.02022f
C871 VDD2.n143 B 0.019059f
C872 VDD2.n144 B 0.011406f
C873 VDD2.n145 B 1.78083f
C874 VDD2.n146 B 0.021227f
C875 VDD2.n147 B 0.011406f
C876 VDD2.n148 B 0.012077f
C877 VDD2.n149 B 0.02696f
C878 VDD2.n150 B 0.02696f
C879 VDD2.n151 B 0.012077f
C880 VDD2.n152 B 0.011406f
C881 VDD2.n153 B 0.021227f
C882 VDD2.n154 B 0.021227f
C883 VDD2.n155 B 0.011406f
C884 VDD2.n156 B 0.012077f
C885 VDD2.n157 B 0.02696f
C886 VDD2.n158 B 0.02696f
C887 VDD2.n159 B 0.012077f
C888 VDD2.n160 B 0.011406f
C889 VDD2.n161 B 0.021227f
C890 VDD2.n162 B 0.021227f
C891 VDD2.n163 B 0.011406f
C892 VDD2.n164 B 0.011742f
C893 VDD2.n165 B 0.011742f
C894 VDD2.n166 B 0.02696f
C895 VDD2.n167 B 0.02696f
C896 VDD2.n168 B 0.012077f
C897 VDD2.n169 B 0.011406f
C898 VDD2.n170 B 0.021227f
C899 VDD2.n171 B 0.021227f
C900 VDD2.n172 B 0.011406f
C901 VDD2.n173 B 0.012077f
C902 VDD2.n174 B 0.02696f
C903 VDD2.n175 B 0.02696f
C904 VDD2.n176 B 0.012077f
C905 VDD2.n177 B 0.011406f
C906 VDD2.n178 B 0.021227f
C907 VDD2.n179 B 0.021227f
C908 VDD2.n180 B 0.011406f
C909 VDD2.n181 B 0.012077f
C910 VDD2.n182 B 0.02696f
C911 VDD2.n183 B 0.02696f
C912 VDD2.n184 B 0.012077f
C913 VDD2.n185 B 0.011406f
C914 VDD2.n186 B 0.021227f
C915 VDD2.n187 B 0.021227f
C916 VDD2.n188 B 0.011406f
C917 VDD2.n189 B 0.012077f
C918 VDD2.n190 B 0.02696f
C919 VDD2.n191 B 0.02696f
C920 VDD2.n192 B 0.012077f
C921 VDD2.n193 B 0.011406f
C922 VDD2.n194 B 0.021227f
C923 VDD2.n195 B 0.021227f
C924 VDD2.n196 B 0.011406f
C925 VDD2.n197 B 0.012077f
C926 VDD2.n198 B 0.02696f
C927 VDD2.n199 B 0.02696f
C928 VDD2.n200 B 0.012077f
C929 VDD2.n201 B 0.011406f
C930 VDD2.n202 B 0.021227f
C931 VDD2.n203 B 0.021227f
C932 VDD2.n204 B 0.011406f
C933 VDD2.n205 B 0.012077f
C934 VDD2.n206 B 0.02696f
C935 VDD2.n207 B 0.055815f
C936 VDD2.n208 B 0.012077f
C937 VDD2.n209 B 0.022303f
C938 VDD2.n210 B 0.054864f
C939 VDD2.n211 B 0.073118f
C940 VDD2.n212 B 2.57968f
C941 VDD2.t3 B 0.327426f
C942 VDD2.t4 B 0.327426f
C943 VDD2.n213 B 3.00277f
C944 VN.n0 B 0.032365f
C945 VN.t1 B 2.94378f
C946 VN.n1 B 0.020112f
C947 VN.n2 B 0.209746f
C948 VN.t2 B 2.94378f
C949 VN.t5 B 3.09951f
C950 VN.n3 B 1.07456f
C951 VN.n4 B 1.08425f
C952 VN.n5 B 0.034289f
C953 VN.n6 B 0.049116f
C954 VN.n7 B 0.024551f
C955 VN.n8 B 0.024551f
C956 VN.n9 B 0.024551f
C957 VN.n10 B 0.047675f
C958 VN.n11 B 0.036986f
C959 VN.n12 B 1.09725f
C960 VN.n13 B 0.034083f
C961 VN.n14 B 0.032365f
C962 VN.t4 B 2.94378f
C963 VN.n15 B 0.020112f
C964 VN.n16 B 0.209746f
C965 VN.t0 B 2.94378f
C966 VN.t3 B 3.09951f
C967 VN.n17 B 1.07456f
C968 VN.n18 B 1.08425f
C969 VN.n19 B 0.034289f
C970 VN.n20 B 0.049116f
C971 VN.n21 B 0.024551f
C972 VN.n22 B 0.024551f
C973 VN.n23 B 0.024551f
C974 VN.n24 B 0.047675f
C975 VN.n25 B 0.036986f
C976 VN.n26 B 1.09725f
C977 VN.n27 B 1.49039f
.ends

