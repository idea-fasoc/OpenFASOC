* NGSPICE file created from diff_pair_sample_1094.ext - technology: sky130A

.subckt diff_pair_sample_1094 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VP.t0 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=1.2771 ps=8.07 w=7.74 l=1.14
X1 VDD1.t0 VP.t1 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=3.0186 ps=16.26 w=7.74 l=1.14
X2 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=3.0186 ps=16.26 w=7.74 l=1.14
X3 VTAIL.t14 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=1.2771 ps=8.07 w=7.74 l=1.14
X4 VDD1.t2 VP.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X5 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=0 ps=0 w=7.74 l=1.14
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=0 ps=0 w=7.74 l=1.14
X7 VDD2.t5 VN.t2 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=3.0186 ps=16.26 w=7.74 l=1.14
X8 VTAIL.t0 VN.t3 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X9 VTAIL.t13 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X10 VDD2.t2 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=0 ps=0 w=7.74 l=1.14
X12 VTAIL.t9 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=1.2771 ps=8.07 w=7.74 l=1.14
X13 VDD1.t3 VP.t4 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=0 ps=0 w=7.74 l=1.14
X15 VDD1.t7 VP.t5 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=3.0186 ps=16.26 w=7.74 l=1.14
X16 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0186 pd=16.26 as=1.2771 ps=8.07 w=7.74 l=1.14
X17 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X18 VTAIL.t6 VP.t6 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
X19 VTAIL.t5 VP.t7 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2771 pd=8.07 as=1.2771 ps=8.07 w=7.74 l=1.14
R0 VP.n7 VP.t3 221.611
R1 VP.n17 VP.t0 198.508
R2 VP.n29 VP.t1 198.508
R3 VP.n15 VP.t5 198.508
R4 VP.n22 VP.t2 163.626
R5 VP.n1 VP.t6 163.626
R6 VP.n5 VP.t7 163.626
R7 VP.n8 VP.t4 163.626
R8 VP.n9 VP.n6 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n4 161.3
R12 VP.n28 VP.n0 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n25 VP.n24 161.3
R15 VP.n23 VP.n2 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n19 VP.n3 161.3
R18 VP.n16 VP.n15 80.6037
R19 VP.n30 VP.n29 80.6037
R20 VP.n18 VP.n17 80.6037
R21 VP.n24 VP.n23 56.4773
R22 VP.n10 VP.n9 56.4773
R23 VP.n17 VP.n3 50.8783
R24 VP.n29 VP.n28 50.8783
R25 VP.n15 VP.n14 50.8783
R26 VP.n18 VP.n16 41.0544
R27 VP.n8 VP.n7 33.4129
R28 VP.n7 VP.n6 28.104
R29 VP.n21 VP.n3 24.3439
R30 VP.n28 VP.n27 24.3439
R31 VP.n14 VP.n13 24.3439
R32 VP.n23 VP.n22 23.6136
R33 VP.n24 VP.n1 23.6136
R34 VP.n10 VP.n5 23.6136
R35 VP.n9 VP.n8 23.6136
R36 VP.n22 VP.n21 0.730803
R37 VP.n27 VP.n1 0.730803
R38 VP.n13 VP.n5 0.730803
R39 VP.n16 VP.n4 0.285035
R40 VP.n19 VP.n18 0.285035
R41 VP.n30 VP.n0 0.285035
R42 VP.n11 VP.n6 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n20 VP.n2 0.189894
R47 VP.n25 VP.n2 0.189894
R48 VP.n26 VP.n25 0.189894
R49 VP.n26 VP.n0 0.189894
R50 VP VP.n30 0.146778
R51 VDD1 VDD1.n0 64.3608
R52 VDD1.n3 VDD1.n2 64.2472
R53 VDD1.n3 VDD1.n1 64.2472
R54 VDD1.n5 VDD1.n4 63.669
R55 VDD1.n5 VDD1.n3 36.6733
R56 VDD1.n4 VDD1.t5 2.55864
R57 VDD1.n4 VDD1.t7 2.55864
R58 VDD1.n0 VDD1.t4 2.55864
R59 VDD1.n0 VDD1.t3 2.55864
R60 VDD1.n2 VDD1.t6 2.55864
R61 VDD1.n2 VDD1.t0 2.55864
R62 VDD1.n1 VDD1.t1 2.55864
R63 VDD1.n1 VDD1.t2 2.55864
R64 VDD1 VDD1.n5 0.575931
R65 VTAIL.n14 VTAIL.t7 49.5483
R66 VTAIL.n11 VTAIL.t9 49.5483
R67 VTAIL.n10 VTAIL.t15 49.5483
R68 VTAIL.n7 VTAIL.t2 49.5483
R69 VTAIL.n15 VTAIL.t1 49.5482
R70 VTAIL.n2 VTAIL.t14 49.5482
R71 VTAIL.n3 VTAIL.t11 49.5482
R72 VTAIL.n6 VTAIL.t12 49.5482
R73 VTAIL.n13 VTAIL.n12 46.9902
R74 VTAIL.n9 VTAIL.n8 46.9902
R75 VTAIL.n1 VTAIL.n0 46.9902
R76 VTAIL.n5 VTAIL.n4 46.9902
R77 VTAIL.n15 VTAIL.n14 20.3065
R78 VTAIL.n7 VTAIL.n6 20.3065
R79 VTAIL.n0 VTAIL.t4 2.55864
R80 VTAIL.n0 VTAIL.t0 2.55864
R81 VTAIL.n4 VTAIL.t10 2.55864
R82 VTAIL.n4 VTAIL.t6 2.55864
R83 VTAIL.n12 VTAIL.t8 2.55864
R84 VTAIL.n12 VTAIL.t5 2.55864
R85 VTAIL.n8 VTAIL.t3 2.55864
R86 VTAIL.n8 VTAIL.t13 2.55864
R87 VTAIL.n9 VTAIL.n7 1.26774
R88 VTAIL.n10 VTAIL.n9 1.26774
R89 VTAIL.n13 VTAIL.n11 1.26774
R90 VTAIL.n14 VTAIL.n13 1.26774
R91 VTAIL.n6 VTAIL.n5 1.26774
R92 VTAIL.n5 VTAIL.n3 1.26774
R93 VTAIL.n2 VTAIL.n1 1.26774
R94 VTAIL VTAIL.n15 1.20955
R95 VTAIL.n11 VTAIL.n10 0.470328
R96 VTAIL.n3 VTAIL.n2 0.470328
R97 VTAIL VTAIL.n1 0.0586897
R98 B.n588 B.n587 585
R99 B.n228 B.n89 585
R100 B.n227 B.n226 585
R101 B.n225 B.n224 585
R102 B.n223 B.n222 585
R103 B.n221 B.n220 585
R104 B.n219 B.n218 585
R105 B.n217 B.n216 585
R106 B.n215 B.n214 585
R107 B.n213 B.n212 585
R108 B.n211 B.n210 585
R109 B.n209 B.n208 585
R110 B.n207 B.n206 585
R111 B.n205 B.n204 585
R112 B.n203 B.n202 585
R113 B.n201 B.n200 585
R114 B.n199 B.n198 585
R115 B.n197 B.n196 585
R116 B.n195 B.n194 585
R117 B.n193 B.n192 585
R118 B.n191 B.n190 585
R119 B.n189 B.n188 585
R120 B.n187 B.n186 585
R121 B.n185 B.n184 585
R122 B.n183 B.n182 585
R123 B.n181 B.n180 585
R124 B.n179 B.n178 585
R125 B.n177 B.n176 585
R126 B.n175 B.n174 585
R127 B.n172 B.n171 585
R128 B.n170 B.n169 585
R129 B.n168 B.n167 585
R130 B.n166 B.n165 585
R131 B.n164 B.n163 585
R132 B.n162 B.n161 585
R133 B.n160 B.n159 585
R134 B.n158 B.n157 585
R135 B.n156 B.n155 585
R136 B.n154 B.n153 585
R137 B.n151 B.n150 585
R138 B.n149 B.n148 585
R139 B.n147 B.n146 585
R140 B.n145 B.n144 585
R141 B.n143 B.n142 585
R142 B.n141 B.n140 585
R143 B.n139 B.n138 585
R144 B.n137 B.n136 585
R145 B.n135 B.n134 585
R146 B.n133 B.n132 585
R147 B.n131 B.n130 585
R148 B.n129 B.n128 585
R149 B.n127 B.n126 585
R150 B.n125 B.n124 585
R151 B.n123 B.n122 585
R152 B.n121 B.n120 585
R153 B.n119 B.n118 585
R154 B.n117 B.n116 585
R155 B.n115 B.n114 585
R156 B.n113 B.n112 585
R157 B.n111 B.n110 585
R158 B.n109 B.n108 585
R159 B.n107 B.n106 585
R160 B.n105 B.n104 585
R161 B.n103 B.n102 585
R162 B.n101 B.n100 585
R163 B.n99 B.n98 585
R164 B.n97 B.n96 585
R165 B.n95 B.n94 585
R166 B.n586 B.n55 585
R167 B.n591 B.n55 585
R168 B.n585 B.n54 585
R169 B.n592 B.n54 585
R170 B.n584 B.n583 585
R171 B.n583 B.n50 585
R172 B.n582 B.n49 585
R173 B.n598 B.n49 585
R174 B.n581 B.n48 585
R175 B.n599 B.n48 585
R176 B.n580 B.n47 585
R177 B.n600 B.n47 585
R178 B.n579 B.n578 585
R179 B.n578 B.n43 585
R180 B.n577 B.n42 585
R181 B.n606 B.n42 585
R182 B.n576 B.n41 585
R183 B.n607 B.n41 585
R184 B.n575 B.n40 585
R185 B.n608 B.n40 585
R186 B.n574 B.n573 585
R187 B.n573 B.n36 585
R188 B.n572 B.n35 585
R189 B.n614 B.n35 585
R190 B.n571 B.n34 585
R191 B.n615 B.n34 585
R192 B.n570 B.n33 585
R193 B.n616 B.n33 585
R194 B.n569 B.n568 585
R195 B.n568 B.n29 585
R196 B.n567 B.n28 585
R197 B.n622 B.n28 585
R198 B.n566 B.n27 585
R199 B.n623 B.n27 585
R200 B.n565 B.n26 585
R201 B.n624 B.n26 585
R202 B.n564 B.n563 585
R203 B.n563 B.n22 585
R204 B.n562 B.n21 585
R205 B.n630 B.n21 585
R206 B.n561 B.n20 585
R207 B.n631 B.n20 585
R208 B.n560 B.n19 585
R209 B.n632 B.n19 585
R210 B.n559 B.n558 585
R211 B.n558 B.n15 585
R212 B.n557 B.n14 585
R213 B.n638 B.n14 585
R214 B.n556 B.n13 585
R215 B.n639 B.n13 585
R216 B.n555 B.n12 585
R217 B.n640 B.n12 585
R218 B.n554 B.n553 585
R219 B.n553 B.n552 585
R220 B.n551 B.n550 585
R221 B.n551 B.n8 585
R222 B.n549 B.n7 585
R223 B.n647 B.n7 585
R224 B.n548 B.n6 585
R225 B.n648 B.n6 585
R226 B.n547 B.n5 585
R227 B.n649 B.n5 585
R228 B.n546 B.n545 585
R229 B.n545 B.n4 585
R230 B.n544 B.n229 585
R231 B.n544 B.n543 585
R232 B.n534 B.n230 585
R233 B.n231 B.n230 585
R234 B.n536 B.n535 585
R235 B.n537 B.n536 585
R236 B.n533 B.n236 585
R237 B.n236 B.n235 585
R238 B.n532 B.n531 585
R239 B.n531 B.n530 585
R240 B.n238 B.n237 585
R241 B.n239 B.n238 585
R242 B.n523 B.n522 585
R243 B.n524 B.n523 585
R244 B.n521 B.n244 585
R245 B.n244 B.n243 585
R246 B.n520 B.n519 585
R247 B.n519 B.n518 585
R248 B.n246 B.n245 585
R249 B.n247 B.n246 585
R250 B.n511 B.n510 585
R251 B.n512 B.n511 585
R252 B.n509 B.n252 585
R253 B.n252 B.n251 585
R254 B.n508 B.n507 585
R255 B.n507 B.n506 585
R256 B.n254 B.n253 585
R257 B.n255 B.n254 585
R258 B.n499 B.n498 585
R259 B.n500 B.n499 585
R260 B.n497 B.n259 585
R261 B.n263 B.n259 585
R262 B.n496 B.n495 585
R263 B.n495 B.n494 585
R264 B.n261 B.n260 585
R265 B.n262 B.n261 585
R266 B.n487 B.n486 585
R267 B.n488 B.n487 585
R268 B.n485 B.n268 585
R269 B.n268 B.n267 585
R270 B.n484 B.n483 585
R271 B.n483 B.n482 585
R272 B.n270 B.n269 585
R273 B.n271 B.n270 585
R274 B.n475 B.n474 585
R275 B.n476 B.n475 585
R276 B.n473 B.n276 585
R277 B.n276 B.n275 585
R278 B.n472 B.n471 585
R279 B.n471 B.n470 585
R280 B.n278 B.n277 585
R281 B.n279 B.n278 585
R282 B.n463 B.n462 585
R283 B.n464 B.n463 585
R284 B.n461 B.n284 585
R285 B.n284 B.n283 585
R286 B.n456 B.n455 585
R287 B.n454 B.n320 585
R288 B.n453 B.n319 585
R289 B.n458 B.n319 585
R290 B.n452 B.n451 585
R291 B.n450 B.n449 585
R292 B.n448 B.n447 585
R293 B.n446 B.n445 585
R294 B.n444 B.n443 585
R295 B.n442 B.n441 585
R296 B.n440 B.n439 585
R297 B.n438 B.n437 585
R298 B.n436 B.n435 585
R299 B.n434 B.n433 585
R300 B.n432 B.n431 585
R301 B.n430 B.n429 585
R302 B.n428 B.n427 585
R303 B.n426 B.n425 585
R304 B.n424 B.n423 585
R305 B.n422 B.n421 585
R306 B.n420 B.n419 585
R307 B.n418 B.n417 585
R308 B.n416 B.n415 585
R309 B.n414 B.n413 585
R310 B.n412 B.n411 585
R311 B.n410 B.n409 585
R312 B.n408 B.n407 585
R313 B.n406 B.n405 585
R314 B.n404 B.n403 585
R315 B.n402 B.n401 585
R316 B.n400 B.n399 585
R317 B.n398 B.n397 585
R318 B.n396 B.n395 585
R319 B.n394 B.n393 585
R320 B.n392 B.n391 585
R321 B.n390 B.n389 585
R322 B.n388 B.n387 585
R323 B.n386 B.n385 585
R324 B.n384 B.n383 585
R325 B.n382 B.n381 585
R326 B.n380 B.n379 585
R327 B.n378 B.n377 585
R328 B.n376 B.n375 585
R329 B.n374 B.n373 585
R330 B.n372 B.n371 585
R331 B.n370 B.n369 585
R332 B.n368 B.n367 585
R333 B.n366 B.n365 585
R334 B.n364 B.n363 585
R335 B.n362 B.n361 585
R336 B.n360 B.n359 585
R337 B.n358 B.n357 585
R338 B.n356 B.n355 585
R339 B.n354 B.n353 585
R340 B.n352 B.n351 585
R341 B.n350 B.n349 585
R342 B.n348 B.n347 585
R343 B.n346 B.n345 585
R344 B.n344 B.n343 585
R345 B.n342 B.n341 585
R346 B.n340 B.n339 585
R347 B.n338 B.n337 585
R348 B.n336 B.n335 585
R349 B.n334 B.n333 585
R350 B.n332 B.n331 585
R351 B.n330 B.n329 585
R352 B.n328 B.n327 585
R353 B.n286 B.n285 585
R354 B.n460 B.n459 585
R355 B.n459 B.n458 585
R356 B.n282 B.n281 585
R357 B.n283 B.n282 585
R358 B.n466 B.n465 585
R359 B.n465 B.n464 585
R360 B.n467 B.n280 585
R361 B.n280 B.n279 585
R362 B.n469 B.n468 585
R363 B.n470 B.n469 585
R364 B.n274 B.n273 585
R365 B.n275 B.n274 585
R366 B.n478 B.n477 585
R367 B.n477 B.n476 585
R368 B.n479 B.n272 585
R369 B.n272 B.n271 585
R370 B.n481 B.n480 585
R371 B.n482 B.n481 585
R372 B.n266 B.n265 585
R373 B.n267 B.n266 585
R374 B.n490 B.n489 585
R375 B.n489 B.n488 585
R376 B.n491 B.n264 585
R377 B.n264 B.n262 585
R378 B.n493 B.n492 585
R379 B.n494 B.n493 585
R380 B.n258 B.n257 585
R381 B.n263 B.n258 585
R382 B.n502 B.n501 585
R383 B.n501 B.n500 585
R384 B.n503 B.n256 585
R385 B.n256 B.n255 585
R386 B.n505 B.n504 585
R387 B.n506 B.n505 585
R388 B.n250 B.n249 585
R389 B.n251 B.n250 585
R390 B.n514 B.n513 585
R391 B.n513 B.n512 585
R392 B.n515 B.n248 585
R393 B.n248 B.n247 585
R394 B.n517 B.n516 585
R395 B.n518 B.n517 585
R396 B.n242 B.n241 585
R397 B.n243 B.n242 585
R398 B.n526 B.n525 585
R399 B.n525 B.n524 585
R400 B.n527 B.n240 585
R401 B.n240 B.n239 585
R402 B.n529 B.n528 585
R403 B.n530 B.n529 585
R404 B.n234 B.n233 585
R405 B.n235 B.n234 585
R406 B.n539 B.n538 585
R407 B.n538 B.n537 585
R408 B.n540 B.n232 585
R409 B.n232 B.n231 585
R410 B.n542 B.n541 585
R411 B.n543 B.n542 585
R412 B.n3 B.n0 585
R413 B.n4 B.n3 585
R414 B.n646 B.n1 585
R415 B.n647 B.n646 585
R416 B.n645 B.n644 585
R417 B.n645 B.n8 585
R418 B.n643 B.n9 585
R419 B.n552 B.n9 585
R420 B.n642 B.n641 585
R421 B.n641 B.n640 585
R422 B.n11 B.n10 585
R423 B.n639 B.n11 585
R424 B.n637 B.n636 585
R425 B.n638 B.n637 585
R426 B.n635 B.n16 585
R427 B.n16 B.n15 585
R428 B.n634 B.n633 585
R429 B.n633 B.n632 585
R430 B.n18 B.n17 585
R431 B.n631 B.n18 585
R432 B.n629 B.n628 585
R433 B.n630 B.n629 585
R434 B.n627 B.n23 585
R435 B.n23 B.n22 585
R436 B.n626 B.n625 585
R437 B.n625 B.n624 585
R438 B.n25 B.n24 585
R439 B.n623 B.n25 585
R440 B.n621 B.n620 585
R441 B.n622 B.n621 585
R442 B.n619 B.n30 585
R443 B.n30 B.n29 585
R444 B.n618 B.n617 585
R445 B.n617 B.n616 585
R446 B.n32 B.n31 585
R447 B.n615 B.n32 585
R448 B.n613 B.n612 585
R449 B.n614 B.n613 585
R450 B.n611 B.n37 585
R451 B.n37 B.n36 585
R452 B.n610 B.n609 585
R453 B.n609 B.n608 585
R454 B.n39 B.n38 585
R455 B.n607 B.n39 585
R456 B.n605 B.n604 585
R457 B.n606 B.n605 585
R458 B.n603 B.n44 585
R459 B.n44 B.n43 585
R460 B.n602 B.n601 585
R461 B.n601 B.n600 585
R462 B.n46 B.n45 585
R463 B.n599 B.n46 585
R464 B.n597 B.n596 585
R465 B.n598 B.n597 585
R466 B.n595 B.n51 585
R467 B.n51 B.n50 585
R468 B.n594 B.n593 585
R469 B.n593 B.n592 585
R470 B.n53 B.n52 585
R471 B.n591 B.n53 585
R472 B.n650 B.n649 585
R473 B.n648 B.n2 585
R474 B.n94 B.n53 516.524
R475 B.n588 B.n55 516.524
R476 B.n459 B.n284 516.524
R477 B.n456 B.n282 516.524
R478 B.n92 B.t16 367.418
R479 B.n90 B.t8 367.418
R480 B.n324 B.t12 367.418
R481 B.n321 B.t19 367.418
R482 B.n590 B.n589 256.663
R483 B.n590 B.n88 256.663
R484 B.n590 B.n87 256.663
R485 B.n590 B.n86 256.663
R486 B.n590 B.n85 256.663
R487 B.n590 B.n84 256.663
R488 B.n590 B.n83 256.663
R489 B.n590 B.n82 256.663
R490 B.n590 B.n81 256.663
R491 B.n590 B.n80 256.663
R492 B.n590 B.n79 256.663
R493 B.n590 B.n78 256.663
R494 B.n590 B.n77 256.663
R495 B.n590 B.n76 256.663
R496 B.n590 B.n75 256.663
R497 B.n590 B.n74 256.663
R498 B.n590 B.n73 256.663
R499 B.n590 B.n72 256.663
R500 B.n590 B.n71 256.663
R501 B.n590 B.n70 256.663
R502 B.n590 B.n69 256.663
R503 B.n590 B.n68 256.663
R504 B.n590 B.n67 256.663
R505 B.n590 B.n66 256.663
R506 B.n590 B.n65 256.663
R507 B.n590 B.n64 256.663
R508 B.n590 B.n63 256.663
R509 B.n590 B.n62 256.663
R510 B.n590 B.n61 256.663
R511 B.n590 B.n60 256.663
R512 B.n590 B.n59 256.663
R513 B.n590 B.n58 256.663
R514 B.n590 B.n57 256.663
R515 B.n590 B.n56 256.663
R516 B.n458 B.n457 256.663
R517 B.n458 B.n287 256.663
R518 B.n458 B.n288 256.663
R519 B.n458 B.n289 256.663
R520 B.n458 B.n290 256.663
R521 B.n458 B.n291 256.663
R522 B.n458 B.n292 256.663
R523 B.n458 B.n293 256.663
R524 B.n458 B.n294 256.663
R525 B.n458 B.n295 256.663
R526 B.n458 B.n296 256.663
R527 B.n458 B.n297 256.663
R528 B.n458 B.n298 256.663
R529 B.n458 B.n299 256.663
R530 B.n458 B.n300 256.663
R531 B.n458 B.n301 256.663
R532 B.n458 B.n302 256.663
R533 B.n458 B.n303 256.663
R534 B.n458 B.n304 256.663
R535 B.n458 B.n305 256.663
R536 B.n458 B.n306 256.663
R537 B.n458 B.n307 256.663
R538 B.n458 B.n308 256.663
R539 B.n458 B.n309 256.663
R540 B.n458 B.n310 256.663
R541 B.n458 B.n311 256.663
R542 B.n458 B.n312 256.663
R543 B.n458 B.n313 256.663
R544 B.n458 B.n314 256.663
R545 B.n458 B.n315 256.663
R546 B.n458 B.n316 256.663
R547 B.n458 B.n317 256.663
R548 B.n458 B.n318 256.663
R549 B.n652 B.n651 256.663
R550 B.n98 B.n97 163.367
R551 B.n102 B.n101 163.367
R552 B.n106 B.n105 163.367
R553 B.n110 B.n109 163.367
R554 B.n114 B.n113 163.367
R555 B.n118 B.n117 163.367
R556 B.n122 B.n121 163.367
R557 B.n126 B.n125 163.367
R558 B.n130 B.n129 163.367
R559 B.n134 B.n133 163.367
R560 B.n138 B.n137 163.367
R561 B.n142 B.n141 163.367
R562 B.n146 B.n145 163.367
R563 B.n150 B.n149 163.367
R564 B.n155 B.n154 163.367
R565 B.n159 B.n158 163.367
R566 B.n163 B.n162 163.367
R567 B.n167 B.n166 163.367
R568 B.n171 B.n170 163.367
R569 B.n176 B.n175 163.367
R570 B.n180 B.n179 163.367
R571 B.n184 B.n183 163.367
R572 B.n188 B.n187 163.367
R573 B.n192 B.n191 163.367
R574 B.n196 B.n195 163.367
R575 B.n200 B.n199 163.367
R576 B.n204 B.n203 163.367
R577 B.n208 B.n207 163.367
R578 B.n212 B.n211 163.367
R579 B.n216 B.n215 163.367
R580 B.n220 B.n219 163.367
R581 B.n224 B.n223 163.367
R582 B.n226 B.n89 163.367
R583 B.n463 B.n284 163.367
R584 B.n463 B.n278 163.367
R585 B.n471 B.n278 163.367
R586 B.n471 B.n276 163.367
R587 B.n475 B.n276 163.367
R588 B.n475 B.n270 163.367
R589 B.n483 B.n270 163.367
R590 B.n483 B.n268 163.367
R591 B.n487 B.n268 163.367
R592 B.n487 B.n261 163.367
R593 B.n495 B.n261 163.367
R594 B.n495 B.n259 163.367
R595 B.n499 B.n259 163.367
R596 B.n499 B.n254 163.367
R597 B.n507 B.n254 163.367
R598 B.n507 B.n252 163.367
R599 B.n511 B.n252 163.367
R600 B.n511 B.n246 163.367
R601 B.n519 B.n246 163.367
R602 B.n519 B.n244 163.367
R603 B.n523 B.n244 163.367
R604 B.n523 B.n238 163.367
R605 B.n531 B.n238 163.367
R606 B.n531 B.n236 163.367
R607 B.n536 B.n236 163.367
R608 B.n536 B.n230 163.367
R609 B.n544 B.n230 163.367
R610 B.n545 B.n544 163.367
R611 B.n545 B.n5 163.367
R612 B.n6 B.n5 163.367
R613 B.n7 B.n6 163.367
R614 B.n551 B.n7 163.367
R615 B.n553 B.n551 163.367
R616 B.n553 B.n12 163.367
R617 B.n13 B.n12 163.367
R618 B.n14 B.n13 163.367
R619 B.n558 B.n14 163.367
R620 B.n558 B.n19 163.367
R621 B.n20 B.n19 163.367
R622 B.n21 B.n20 163.367
R623 B.n563 B.n21 163.367
R624 B.n563 B.n26 163.367
R625 B.n27 B.n26 163.367
R626 B.n28 B.n27 163.367
R627 B.n568 B.n28 163.367
R628 B.n568 B.n33 163.367
R629 B.n34 B.n33 163.367
R630 B.n35 B.n34 163.367
R631 B.n573 B.n35 163.367
R632 B.n573 B.n40 163.367
R633 B.n41 B.n40 163.367
R634 B.n42 B.n41 163.367
R635 B.n578 B.n42 163.367
R636 B.n578 B.n47 163.367
R637 B.n48 B.n47 163.367
R638 B.n49 B.n48 163.367
R639 B.n583 B.n49 163.367
R640 B.n583 B.n54 163.367
R641 B.n55 B.n54 163.367
R642 B.n320 B.n319 163.367
R643 B.n451 B.n319 163.367
R644 B.n449 B.n448 163.367
R645 B.n445 B.n444 163.367
R646 B.n441 B.n440 163.367
R647 B.n437 B.n436 163.367
R648 B.n433 B.n432 163.367
R649 B.n429 B.n428 163.367
R650 B.n425 B.n424 163.367
R651 B.n421 B.n420 163.367
R652 B.n417 B.n416 163.367
R653 B.n413 B.n412 163.367
R654 B.n409 B.n408 163.367
R655 B.n405 B.n404 163.367
R656 B.n401 B.n400 163.367
R657 B.n397 B.n396 163.367
R658 B.n393 B.n392 163.367
R659 B.n389 B.n388 163.367
R660 B.n385 B.n384 163.367
R661 B.n381 B.n380 163.367
R662 B.n377 B.n376 163.367
R663 B.n373 B.n372 163.367
R664 B.n369 B.n368 163.367
R665 B.n365 B.n364 163.367
R666 B.n361 B.n360 163.367
R667 B.n357 B.n356 163.367
R668 B.n353 B.n352 163.367
R669 B.n349 B.n348 163.367
R670 B.n345 B.n344 163.367
R671 B.n341 B.n340 163.367
R672 B.n337 B.n336 163.367
R673 B.n333 B.n332 163.367
R674 B.n329 B.n328 163.367
R675 B.n459 B.n286 163.367
R676 B.n465 B.n282 163.367
R677 B.n465 B.n280 163.367
R678 B.n469 B.n280 163.367
R679 B.n469 B.n274 163.367
R680 B.n477 B.n274 163.367
R681 B.n477 B.n272 163.367
R682 B.n481 B.n272 163.367
R683 B.n481 B.n266 163.367
R684 B.n489 B.n266 163.367
R685 B.n489 B.n264 163.367
R686 B.n493 B.n264 163.367
R687 B.n493 B.n258 163.367
R688 B.n501 B.n258 163.367
R689 B.n501 B.n256 163.367
R690 B.n505 B.n256 163.367
R691 B.n505 B.n250 163.367
R692 B.n513 B.n250 163.367
R693 B.n513 B.n248 163.367
R694 B.n517 B.n248 163.367
R695 B.n517 B.n242 163.367
R696 B.n525 B.n242 163.367
R697 B.n525 B.n240 163.367
R698 B.n529 B.n240 163.367
R699 B.n529 B.n234 163.367
R700 B.n538 B.n234 163.367
R701 B.n538 B.n232 163.367
R702 B.n542 B.n232 163.367
R703 B.n542 B.n3 163.367
R704 B.n650 B.n3 163.367
R705 B.n646 B.n2 163.367
R706 B.n646 B.n645 163.367
R707 B.n645 B.n9 163.367
R708 B.n641 B.n9 163.367
R709 B.n641 B.n11 163.367
R710 B.n637 B.n11 163.367
R711 B.n637 B.n16 163.367
R712 B.n633 B.n16 163.367
R713 B.n633 B.n18 163.367
R714 B.n629 B.n18 163.367
R715 B.n629 B.n23 163.367
R716 B.n625 B.n23 163.367
R717 B.n625 B.n25 163.367
R718 B.n621 B.n25 163.367
R719 B.n621 B.n30 163.367
R720 B.n617 B.n30 163.367
R721 B.n617 B.n32 163.367
R722 B.n613 B.n32 163.367
R723 B.n613 B.n37 163.367
R724 B.n609 B.n37 163.367
R725 B.n609 B.n39 163.367
R726 B.n605 B.n39 163.367
R727 B.n605 B.n44 163.367
R728 B.n601 B.n44 163.367
R729 B.n601 B.n46 163.367
R730 B.n597 B.n46 163.367
R731 B.n597 B.n51 163.367
R732 B.n593 B.n51 163.367
R733 B.n593 B.n53 163.367
R734 B.n458 B.n283 117.481
R735 B.n591 B.n590 117.481
R736 B.n90 B.t10 102.245
R737 B.n324 B.t15 102.245
R738 B.n92 B.t17 102.236
R739 B.n321 B.t21 102.236
R740 B.n91 B.t11 73.7354
R741 B.n325 B.t14 73.7354
R742 B.n93 B.t18 73.7266
R743 B.n322 B.t20 73.7266
R744 B.n94 B.n56 71.676
R745 B.n98 B.n57 71.676
R746 B.n102 B.n58 71.676
R747 B.n106 B.n59 71.676
R748 B.n110 B.n60 71.676
R749 B.n114 B.n61 71.676
R750 B.n118 B.n62 71.676
R751 B.n122 B.n63 71.676
R752 B.n126 B.n64 71.676
R753 B.n130 B.n65 71.676
R754 B.n134 B.n66 71.676
R755 B.n138 B.n67 71.676
R756 B.n142 B.n68 71.676
R757 B.n146 B.n69 71.676
R758 B.n150 B.n70 71.676
R759 B.n155 B.n71 71.676
R760 B.n159 B.n72 71.676
R761 B.n163 B.n73 71.676
R762 B.n167 B.n74 71.676
R763 B.n171 B.n75 71.676
R764 B.n176 B.n76 71.676
R765 B.n180 B.n77 71.676
R766 B.n184 B.n78 71.676
R767 B.n188 B.n79 71.676
R768 B.n192 B.n80 71.676
R769 B.n196 B.n81 71.676
R770 B.n200 B.n82 71.676
R771 B.n204 B.n83 71.676
R772 B.n208 B.n84 71.676
R773 B.n212 B.n85 71.676
R774 B.n216 B.n86 71.676
R775 B.n220 B.n87 71.676
R776 B.n224 B.n88 71.676
R777 B.n589 B.n89 71.676
R778 B.n589 B.n588 71.676
R779 B.n226 B.n88 71.676
R780 B.n223 B.n87 71.676
R781 B.n219 B.n86 71.676
R782 B.n215 B.n85 71.676
R783 B.n211 B.n84 71.676
R784 B.n207 B.n83 71.676
R785 B.n203 B.n82 71.676
R786 B.n199 B.n81 71.676
R787 B.n195 B.n80 71.676
R788 B.n191 B.n79 71.676
R789 B.n187 B.n78 71.676
R790 B.n183 B.n77 71.676
R791 B.n179 B.n76 71.676
R792 B.n175 B.n75 71.676
R793 B.n170 B.n74 71.676
R794 B.n166 B.n73 71.676
R795 B.n162 B.n72 71.676
R796 B.n158 B.n71 71.676
R797 B.n154 B.n70 71.676
R798 B.n149 B.n69 71.676
R799 B.n145 B.n68 71.676
R800 B.n141 B.n67 71.676
R801 B.n137 B.n66 71.676
R802 B.n133 B.n65 71.676
R803 B.n129 B.n64 71.676
R804 B.n125 B.n63 71.676
R805 B.n121 B.n62 71.676
R806 B.n117 B.n61 71.676
R807 B.n113 B.n60 71.676
R808 B.n109 B.n59 71.676
R809 B.n105 B.n58 71.676
R810 B.n101 B.n57 71.676
R811 B.n97 B.n56 71.676
R812 B.n457 B.n456 71.676
R813 B.n451 B.n287 71.676
R814 B.n448 B.n288 71.676
R815 B.n444 B.n289 71.676
R816 B.n440 B.n290 71.676
R817 B.n436 B.n291 71.676
R818 B.n432 B.n292 71.676
R819 B.n428 B.n293 71.676
R820 B.n424 B.n294 71.676
R821 B.n420 B.n295 71.676
R822 B.n416 B.n296 71.676
R823 B.n412 B.n297 71.676
R824 B.n408 B.n298 71.676
R825 B.n404 B.n299 71.676
R826 B.n400 B.n300 71.676
R827 B.n396 B.n301 71.676
R828 B.n392 B.n302 71.676
R829 B.n388 B.n303 71.676
R830 B.n384 B.n304 71.676
R831 B.n380 B.n305 71.676
R832 B.n376 B.n306 71.676
R833 B.n372 B.n307 71.676
R834 B.n368 B.n308 71.676
R835 B.n364 B.n309 71.676
R836 B.n360 B.n310 71.676
R837 B.n356 B.n311 71.676
R838 B.n352 B.n312 71.676
R839 B.n348 B.n313 71.676
R840 B.n344 B.n314 71.676
R841 B.n340 B.n315 71.676
R842 B.n336 B.n316 71.676
R843 B.n332 B.n317 71.676
R844 B.n328 B.n318 71.676
R845 B.n457 B.n320 71.676
R846 B.n449 B.n287 71.676
R847 B.n445 B.n288 71.676
R848 B.n441 B.n289 71.676
R849 B.n437 B.n290 71.676
R850 B.n433 B.n291 71.676
R851 B.n429 B.n292 71.676
R852 B.n425 B.n293 71.676
R853 B.n421 B.n294 71.676
R854 B.n417 B.n295 71.676
R855 B.n413 B.n296 71.676
R856 B.n409 B.n297 71.676
R857 B.n405 B.n298 71.676
R858 B.n401 B.n299 71.676
R859 B.n397 B.n300 71.676
R860 B.n393 B.n301 71.676
R861 B.n389 B.n302 71.676
R862 B.n385 B.n303 71.676
R863 B.n381 B.n304 71.676
R864 B.n377 B.n305 71.676
R865 B.n373 B.n306 71.676
R866 B.n369 B.n307 71.676
R867 B.n365 B.n308 71.676
R868 B.n361 B.n309 71.676
R869 B.n357 B.n310 71.676
R870 B.n353 B.n311 71.676
R871 B.n349 B.n312 71.676
R872 B.n345 B.n313 71.676
R873 B.n341 B.n314 71.676
R874 B.n337 B.n315 71.676
R875 B.n333 B.n316 71.676
R876 B.n329 B.n317 71.676
R877 B.n318 B.n286 71.676
R878 B.n651 B.n650 71.676
R879 B.n651 B.n2 71.676
R880 B.n152 B.n93 59.5399
R881 B.n173 B.n91 59.5399
R882 B.n326 B.n325 59.5399
R883 B.n323 B.n322 59.5399
R884 B.n464 B.n283 57.4726
R885 B.n464 B.n279 57.4726
R886 B.n470 B.n279 57.4726
R887 B.n470 B.n275 57.4726
R888 B.n476 B.n275 57.4726
R889 B.n482 B.n271 57.4726
R890 B.n482 B.n267 57.4726
R891 B.n488 B.n267 57.4726
R892 B.n488 B.n262 57.4726
R893 B.n494 B.n262 57.4726
R894 B.n494 B.n263 57.4726
R895 B.n500 B.n255 57.4726
R896 B.n506 B.n255 57.4726
R897 B.n506 B.n251 57.4726
R898 B.n512 B.n251 57.4726
R899 B.n518 B.n247 57.4726
R900 B.n518 B.n243 57.4726
R901 B.n524 B.n243 57.4726
R902 B.n530 B.n239 57.4726
R903 B.n530 B.n235 57.4726
R904 B.n537 B.n235 57.4726
R905 B.n543 B.n231 57.4726
R906 B.n543 B.n4 57.4726
R907 B.n649 B.n4 57.4726
R908 B.n649 B.n648 57.4726
R909 B.n648 B.n647 57.4726
R910 B.n647 B.n8 57.4726
R911 B.n552 B.n8 57.4726
R912 B.n640 B.n639 57.4726
R913 B.n639 B.n638 57.4726
R914 B.n638 B.n15 57.4726
R915 B.n632 B.n631 57.4726
R916 B.n631 B.n630 57.4726
R917 B.n630 B.n22 57.4726
R918 B.n624 B.n623 57.4726
R919 B.n623 B.n622 57.4726
R920 B.n622 B.n29 57.4726
R921 B.n616 B.n29 57.4726
R922 B.n615 B.n614 57.4726
R923 B.n614 B.n36 57.4726
R924 B.n608 B.n36 57.4726
R925 B.n608 B.n607 57.4726
R926 B.n607 B.n606 57.4726
R927 B.n606 B.n43 57.4726
R928 B.n600 B.n599 57.4726
R929 B.n599 B.n598 57.4726
R930 B.n598 B.n50 57.4726
R931 B.n592 B.n50 57.4726
R932 B.n592 B.n591 57.4726
R933 B.t3 B.n247 52.4016
R934 B.t0 B.n22 52.4016
R935 B.t13 B.n271 43.9498
R936 B.n263 B.t2 43.9498
R937 B.t1 B.n615 43.9498
R938 B.t9 B.n43 43.9498
R939 B.n537 B.t7 42.2594
R940 B.n640 B.t6 42.2594
R941 B.t5 B.n239 33.8076
R942 B.t4 B.n15 33.8076
R943 B.n455 B.n281 33.5615
R944 B.n461 B.n460 33.5615
R945 B.n587 B.n586 33.5615
R946 B.n95 B.n52 33.5615
R947 B.n93 B.n92 28.5096
R948 B.n91 B.n90 28.5096
R949 B.n325 B.n324 28.5096
R950 B.n322 B.n321 28.5096
R951 B.n524 B.t5 23.6655
R952 B.n632 B.t4 23.6655
R953 B B.n652 18.0485
R954 B.t7 B.n231 15.2137
R955 B.n552 B.t6 15.2137
R956 B.n476 B.t13 13.5234
R957 B.n500 B.t2 13.5234
R958 B.n616 B.t1 13.5234
R959 B.n600 B.t9 13.5234
R960 B.n466 B.n281 10.6151
R961 B.n467 B.n466 10.6151
R962 B.n468 B.n467 10.6151
R963 B.n468 B.n273 10.6151
R964 B.n478 B.n273 10.6151
R965 B.n479 B.n478 10.6151
R966 B.n480 B.n479 10.6151
R967 B.n480 B.n265 10.6151
R968 B.n490 B.n265 10.6151
R969 B.n491 B.n490 10.6151
R970 B.n492 B.n491 10.6151
R971 B.n492 B.n257 10.6151
R972 B.n502 B.n257 10.6151
R973 B.n503 B.n502 10.6151
R974 B.n504 B.n503 10.6151
R975 B.n504 B.n249 10.6151
R976 B.n514 B.n249 10.6151
R977 B.n515 B.n514 10.6151
R978 B.n516 B.n515 10.6151
R979 B.n516 B.n241 10.6151
R980 B.n526 B.n241 10.6151
R981 B.n527 B.n526 10.6151
R982 B.n528 B.n527 10.6151
R983 B.n528 B.n233 10.6151
R984 B.n539 B.n233 10.6151
R985 B.n540 B.n539 10.6151
R986 B.n541 B.n540 10.6151
R987 B.n541 B.n0 10.6151
R988 B.n455 B.n454 10.6151
R989 B.n454 B.n453 10.6151
R990 B.n453 B.n452 10.6151
R991 B.n452 B.n450 10.6151
R992 B.n450 B.n447 10.6151
R993 B.n447 B.n446 10.6151
R994 B.n446 B.n443 10.6151
R995 B.n443 B.n442 10.6151
R996 B.n442 B.n439 10.6151
R997 B.n439 B.n438 10.6151
R998 B.n438 B.n435 10.6151
R999 B.n435 B.n434 10.6151
R1000 B.n434 B.n431 10.6151
R1001 B.n431 B.n430 10.6151
R1002 B.n430 B.n427 10.6151
R1003 B.n427 B.n426 10.6151
R1004 B.n426 B.n423 10.6151
R1005 B.n423 B.n422 10.6151
R1006 B.n422 B.n419 10.6151
R1007 B.n419 B.n418 10.6151
R1008 B.n418 B.n415 10.6151
R1009 B.n415 B.n414 10.6151
R1010 B.n414 B.n411 10.6151
R1011 B.n411 B.n410 10.6151
R1012 B.n410 B.n407 10.6151
R1013 B.n407 B.n406 10.6151
R1014 B.n406 B.n403 10.6151
R1015 B.n403 B.n402 10.6151
R1016 B.n399 B.n398 10.6151
R1017 B.n398 B.n395 10.6151
R1018 B.n395 B.n394 10.6151
R1019 B.n394 B.n391 10.6151
R1020 B.n391 B.n390 10.6151
R1021 B.n390 B.n387 10.6151
R1022 B.n387 B.n386 10.6151
R1023 B.n386 B.n383 10.6151
R1024 B.n383 B.n382 10.6151
R1025 B.n379 B.n378 10.6151
R1026 B.n378 B.n375 10.6151
R1027 B.n375 B.n374 10.6151
R1028 B.n374 B.n371 10.6151
R1029 B.n371 B.n370 10.6151
R1030 B.n370 B.n367 10.6151
R1031 B.n367 B.n366 10.6151
R1032 B.n366 B.n363 10.6151
R1033 B.n363 B.n362 10.6151
R1034 B.n362 B.n359 10.6151
R1035 B.n359 B.n358 10.6151
R1036 B.n358 B.n355 10.6151
R1037 B.n355 B.n354 10.6151
R1038 B.n354 B.n351 10.6151
R1039 B.n351 B.n350 10.6151
R1040 B.n350 B.n347 10.6151
R1041 B.n347 B.n346 10.6151
R1042 B.n346 B.n343 10.6151
R1043 B.n343 B.n342 10.6151
R1044 B.n342 B.n339 10.6151
R1045 B.n339 B.n338 10.6151
R1046 B.n338 B.n335 10.6151
R1047 B.n335 B.n334 10.6151
R1048 B.n334 B.n331 10.6151
R1049 B.n331 B.n330 10.6151
R1050 B.n330 B.n327 10.6151
R1051 B.n327 B.n285 10.6151
R1052 B.n460 B.n285 10.6151
R1053 B.n462 B.n461 10.6151
R1054 B.n462 B.n277 10.6151
R1055 B.n472 B.n277 10.6151
R1056 B.n473 B.n472 10.6151
R1057 B.n474 B.n473 10.6151
R1058 B.n474 B.n269 10.6151
R1059 B.n484 B.n269 10.6151
R1060 B.n485 B.n484 10.6151
R1061 B.n486 B.n485 10.6151
R1062 B.n486 B.n260 10.6151
R1063 B.n496 B.n260 10.6151
R1064 B.n497 B.n496 10.6151
R1065 B.n498 B.n497 10.6151
R1066 B.n498 B.n253 10.6151
R1067 B.n508 B.n253 10.6151
R1068 B.n509 B.n508 10.6151
R1069 B.n510 B.n509 10.6151
R1070 B.n510 B.n245 10.6151
R1071 B.n520 B.n245 10.6151
R1072 B.n521 B.n520 10.6151
R1073 B.n522 B.n521 10.6151
R1074 B.n522 B.n237 10.6151
R1075 B.n532 B.n237 10.6151
R1076 B.n533 B.n532 10.6151
R1077 B.n535 B.n533 10.6151
R1078 B.n535 B.n534 10.6151
R1079 B.n534 B.n229 10.6151
R1080 B.n546 B.n229 10.6151
R1081 B.n547 B.n546 10.6151
R1082 B.n548 B.n547 10.6151
R1083 B.n549 B.n548 10.6151
R1084 B.n550 B.n549 10.6151
R1085 B.n554 B.n550 10.6151
R1086 B.n555 B.n554 10.6151
R1087 B.n556 B.n555 10.6151
R1088 B.n557 B.n556 10.6151
R1089 B.n559 B.n557 10.6151
R1090 B.n560 B.n559 10.6151
R1091 B.n561 B.n560 10.6151
R1092 B.n562 B.n561 10.6151
R1093 B.n564 B.n562 10.6151
R1094 B.n565 B.n564 10.6151
R1095 B.n566 B.n565 10.6151
R1096 B.n567 B.n566 10.6151
R1097 B.n569 B.n567 10.6151
R1098 B.n570 B.n569 10.6151
R1099 B.n571 B.n570 10.6151
R1100 B.n572 B.n571 10.6151
R1101 B.n574 B.n572 10.6151
R1102 B.n575 B.n574 10.6151
R1103 B.n576 B.n575 10.6151
R1104 B.n577 B.n576 10.6151
R1105 B.n579 B.n577 10.6151
R1106 B.n580 B.n579 10.6151
R1107 B.n581 B.n580 10.6151
R1108 B.n582 B.n581 10.6151
R1109 B.n584 B.n582 10.6151
R1110 B.n585 B.n584 10.6151
R1111 B.n586 B.n585 10.6151
R1112 B.n644 B.n1 10.6151
R1113 B.n644 B.n643 10.6151
R1114 B.n643 B.n642 10.6151
R1115 B.n642 B.n10 10.6151
R1116 B.n636 B.n10 10.6151
R1117 B.n636 B.n635 10.6151
R1118 B.n635 B.n634 10.6151
R1119 B.n634 B.n17 10.6151
R1120 B.n628 B.n17 10.6151
R1121 B.n628 B.n627 10.6151
R1122 B.n627 B.n626 10.6151
R1123 B.n626 B.n24 10.6151
R1124 B.n620 B.n24 10.6151
R1125 B.n620 B.n619 10.6151
R1126 B.n619 B.n618 10.6151
R1127 B.n618 B.n31 10.6151
R1128 B.n612 B.n31 10.6151
R1129 B.n612 B.n611 10.6151
R1130 B.n611 B.n610 10.6151
R1131 B.n610 B.n38 10.6151
R1132 B.n604 B.n38 10.6151
R1133 B.n604 B.n603 10.6151
R1134 B.n603 B.n602 10.6151
R1135 B.n602 B.n45 10.6151
R1136 B.n596 B.n45 10.6151
R1137 B.n596 B.n595 10.6151
R1138 B.n595 B.n594 10.6151
R1139 B.n594 B.n52 10.6151
R1140 B.n96 B.n95 10.6151
R1141 B.n99 B.n96 10.6151
R1142 B.n100 B.n99 10.6151
R1143 B.n103 B.n100 10.6151
R1144 B.n104 B.n103 10.6151
R1145 B.n107 B.n104 10.6151
R1146 B.n108 B.n107 10.6151
R1147 B.n111 B.n108 10.6151
R1148 B.n112 B.n111 10.6151
R1149 B.n115 B.n112 10.6151
R1150 B.n116 B.n115 10.6151
R1151 B.n119 B.n116 10.6151
R1152 B.n120 B.n119 10.6151
R1153 B.n123 B.n120 10.6151
R1154 B.n124 B.n123 10.6151
R1155 B.n127 B.n124 10.6151
R1156 B.n128 B.n127 10.6151
R1157 B.n131 B.n128 10.6151
R1158 B.n132 B.n131 10.6151
R1159 B.n135 B.n132 10.6151
R1160 B.n136 B.n135 10.6151
R1161 B.n139 B.n136 10.6151
R1162 B.n140 B.n139 10.6151
R1163 B.n143 B.n140 10.6151
R1164 B.n144 B.n143 10.6151
R1165 B.n147 B.n144 10.6151
R1166 B.n148 B.n147 10.6151
R1167 B.n151 B.n148 10.6151
R1168 B.n156 B.n153 10.6151
R1169 B.n157 B.n156 10.6151
R1170 B.n160 B.n157 10.6151
R1171 B.n161 B.n160 10.6151
R1172 B.n164 B.n161 10.6151
R1173 B.n165 B.n164 10.6151
R1174 B.n168 B.n165 10.6151
R1175 B.n169 B.n168 10.6151
R1176 B.n172 B.n169 10.6151
R1177 B.n177 B.n174 10.6151
R1178 B.n178 B.n177 10.6151
R1179 B.n181 B.n178 10.6151
R1180 B.n182 B.n181 10.6151
R1181 B.n185 B.n182 10.6151
R1182 B.n186 B.n185 10.6151
R1183 B.n189 B.n186 10.6151
R1184 B.n190 B.n189 10.6151
R1185 B.n193 B.n190 10.6151
R1186 B.n194 B.n193 10.6151
R1187 B.n197 B.n194 10.6151
R1188 B.n198 B.n197 10.6151
R1189 B.n201 B.n198 10.6151
R1190 B.n202 B.n201 10.6151
R1191 B.n205 B.n202 10.6151
R1192 B.n206 B.n205 10.6151
R1193 B.n209 B.n206 10.6151
R1194 B.n210 B.n209 10.6151
R1195 B.n213 B.n210 10.6151
R1196 B.n214 B.n213 10.6151
R1197 B.n217 B.n214 10.6151
R1198 B.n218 B.n217 10.6151
R1199 B.n221 B.n218 10.6151
R1200 B.n222 B.n221 10.6151
R1201 B.n225 B.n222 10.6151
R1202 B.n227 B.n225 10.6151
R1203 B.n228 B.n227 10.6151
R1204 B.n587 B.n228 10.6151
R1205 B.n402 B.n323 9.36635
R1206 B.n379 B.n326 9.36635
R1207 B.n152 B.n151 9.36635
R1208 B.n174 B.n173 9.36635
R1209 B.n652 B.n0 8.11757
R1210 B.n652 B.n1 8.11757
R1211 B.n512 B.t3 5.07157
R1212 B.n624 B.t0 5.07157
R1213 B.n399 B.n323 1.24928
R1214 B.n382 B.n326 1.24928
R1215 B.n153 B.n152 1.24928
R1216 B.n173 B.n172 1.24928
R1217 VN.n3 VN.t1 221.611
R1218 VN.n16 VN.t2 221.611
R1219 VN.n11 VN.t0 198.508
R1220 VN.n24 VN.t6 198.508
R1221 VN.n4 VN.t7 163.626
R1222 VN.n1 VN.t3 163.626
R1223 VN.n17 VN.t4 163.626
R1224 VN.n14 VN.t5 163.626
R1225 VN.n23 VN.n13 161.3
R1226 VN.n22 VN.n21 161.3
R1227 VN.n20 VN.n19 161.3
R1228 VN.n18 VN.n15 161.3
R1229 VN.n10 VN.n0 161.3
R1230 VN.n9 VN.n8 161.3
R1231 VN.n7 VN.n6 161.3
R1232 VN.n5 VN.n2 161.3
R1233 VN.n25 VN.n24 80.6037
R1234 VN.n12 VN.n11 80.6037
R1235 VN.n6 VN.n5 56.4773
R1236 VN.n19 VN.n18 56.4773
R1237 VN.n11 VN.n10 50.8783
R1238 VN.n24 VN.n23 50.8783
R1239 VN VN.n25 41.34
R1240 VN.n4 VN.n3 33.4129
R1241 VN.n17 VN.n16 33.4129
R1242 VN.n16 VN.n15 28.104
R1243 VN.n3 VN.n2 28.104
R1244 VN.n10 VN.n9 24.3439
R1245 VN.n23 VN.n22 24.3439
R1246 VN.n5 VN.n4 23.6136
R1247 VN.n6 VN.n1 23.6136
R1248 VN.n18 VN.n17 23.6136
R1249 VN.n19 VN.n14 23.6136
R1250 VN.n9 VN.n1 0.730803
R1251 VN.n22 VN.n14 0.730803
R1252 VN.n25 VN.n13 0.285035
R1253 VN.n12 VN.n0 0.285035
R1254 VN.n21 VN.n13 0.189894
R1255 VN.n21 VN.n20 0.189894
R1256 VN.n20 VN.n15 0.189894
R1257 VN.n7 VN.n2 0.189894
R1258 VN.n8 VN.n7 0.189894
R1259 VN.n8 VN.n0 0.189894
R1260 VN VN.n12 0.146778
R1261 VDD2.n2 VDD2.n1 64.2472
R1262 VDD2.n2 VDD2.n0 64.2472
R1263 VDD2 VDD2.n5 64.2444
R1264 VDD2.n4 VDD2.n3 63.669
R1265 VDD2.n4 VDD2.n2 36.0903
R1266 VDD2.n5 VDD2.t3 2.55864
R1267 VDD2.n5 VDD2.t5 2.55864
R1268 VDD2.n3 VDD2.t1 2.55864
R1269 VDD2.n3 VDD2.t2 2.55864
R1270 VDD2.n1 VDD2.t4 2.55864
R1271 VDD2.n1 VDD2.t7 2.55864
R1272 VDD2.n0 VDD2.t6 2.55864
R1273 VDD2.n0 VDD2.t0 2.55864
R1274 VDD2 VDD2.n4 0.69231
C0 VP VN 5.08903f
C1 VDD2 VN 4.56709f
C2 VDD1 VN 0.148813f
C3 VTAIL VN 4.65754f
C4 VP VDD2 0.364036f
C5 VP VDD1 4.78166f
C6 VDD1 VDD2 1.04669f
C7 VTAIL VP 4.67165f
C8 VTAIL VDD2 6.84852f
C9 VTAIL VDD1 6.80389f
C10 VDD2 B 3.588057f
C11 VDD1 B 3.870937f
C12 VTAIL B 6.903407f
C13 VN B 9.67345f
C14 VP B 8.080469f
C15 VDD2.t6 B 0.155254f
C16 VDD2.t0 B 0.155254f
C17 VDD2.n0 B 1.33367f
C18 VDD2.t4 B 0.155254f
C19 VDD2.t7 B 0.155254f
C20 VDD2.n1 B 1.33367f
C21 VDD2.n2 B 2.20883f
C22 VDD2.t1 B 0.155254f
C23 VDD2.t2 B 0.155254f
C24 VDD2.n3 B 1.33031f
C25 VDD2.n4 B 2.14505f
C26 VDD2.t3 B 0.155254f
C27 VDD2.t5 B 0.155254f
C28 VDD2.n5 B 1.33365f
C29 VN.n0 B 0.049057f
C30 VN.t3 B 0.869942f
C31 VN.n1 B 0.337031f
C32 VN.n2 B 0.194438f
C33 VN.t7 B 0.869942f
C34 VN.t1 B 0.977565f
C35 VN.n3 B 0.386345f
C36 VN.n4 B 0.39789f
C37 VN.n5 B 0.052882f
C38 VN.n6 B 0.052882f
C39 VN.n7 B 0.036764f
C40 VN.n8 B 0.036764f
C41 VN.n9 B 0.035882f
C42 VN.n10 B 0.049232f
C43 VN.t0 B 0.934542f
C44 VN.n11 B 0.403266f
C45 VN.n12 B 0.034431f
C46 VN.n13 B 0.049057f
C47 VN.t5 B 0.869942f
C48 VN.n14 B 0.337031f
C49 VN.n15 B 0.194438f
C50 VN.t4 B 0.869942f
C51 VN.t2 B 0.977565f
C52 VN.n16 B 0.386345f
C53 VN.n17 B 0.39789f
C54 VN.n18 B 0.052882f
C55 VN.n19 B 0.052882f
C56 VN.n20 B 0.036764f
C57 VN.n21 B 0.036764f
C58 VN.n22 B 0.035882f
C59 VN.n23 B 0.049232f
C60 VN.t6 B 0.934542f
C61 VN.n24 B 0.403266f
C62 VN.n25 B 1.4944f
C63 VTAIL.t4 B 0.125264f
C64 VTAIL.t0 B 0.125264f
C65 VTAIL.n0 B 1.01414f
C66 VTAIL.n1 B 0.289506f
C67 VTAIL.t14 B 1.29224f
C68 VTAIL.n2 B 0.380206f
C69 VTAIL.t11 B 1.29224f
C70 VTAIL.n3 B 0.380206f
C71 VTAIL.t10 B 0.125264f
C72 VTAIL.t6 B 0.125264f
C73 VTAIL.n4 B 1.01414f
C74 VTAIL.n5 B 0.369293f
C75 VTAIL.t12 B 1.29224f
C76 VTAIL.n6 B 1.15135f
C77 VTAIL.t2 B 1.29225f
C78 VTAIL.n7 B 1.15134f
C79 VTAIL.t3 B 0.125264f
C80 VTAIL.t13 B 0.125264f
C81 VTAIL.n8 B 1.01415f
C82 VTAIL.n9 B 0.369291f
C83 VTAIL.t15 B 1.29225f
C84 VTAIL.n10 B 0.380198f
C85 VTAIL.t9 B 1.29225f
C86 VTAIL.n11 B 0.380198f
C87 VTAIL.t8 B 0.125264f
C88 VTAIL.t5 B 0.125264f
C89 VTAIL.n12 B 1.01415f
C90 VTAIL.n13 B 0.369291f
C91 VTAIL.t7 B 1.29225f
C92 VTAIL.n14 B 1.15134f
C93 VTAIL.t1 B 1.29224f
C94 VTAIL.n15 B 1.14751f
C95 VDD1.t4 B 0.156689f
C96 VDD1.t3 B 0.156689f
C97 VDD1.n0 B 1.34675f
C98 VDD1.t1 B 0.156689f
C99 VDD1.t2 B 0.156689f
C100 VDD1.n1 B 1.346f
C101 VDD1.t6 B 0.156689f
C102 VDD1.t0 B 0.156689f
C103 VDD1.n2 B 1.346f
C104 VDD1.n3 B 2.28375f
C105 VDD1.t5 B 0.156689f
C106 VDD1.t7 B 0.156689f
C107 VDD1.n4 B 1.34261f
C108 VDD1.n5 B 2.19539f
C109 VP.n0 B 0.049917f
C110 VP.t6 B 0.885201f
C111 VP.n1 B 0.342943f
C112 VP.n2 B 0.037409f
C113 VP.t2 B 0.885201f
C114 VP.n3 B 0.050095f
C115 VP.n4 B 0.049917f
C116 VP.t5 B 0.950934f
C117 VP.t7 B 0.885201f
C118 VP.n5 B 0.342943f
C119 VP.n6 B 0.197849f
C120 VP.t4 B 0.885201f
C121 VP.t3 B 0.994712f
C122 VP.n7 B 0.393122f
C123 VP.n8 B 0.404869f
C124 VP.n9 B 0.05381f
C125 VP.n10 B 0.05381f
C126 VP.n11 B 0.037409f
C127 VP.n12 B 0.037409f
C128 VP.n13 B 0.036512f
C129 VP.n14 B 0.050095f
C130 VP.n15 B 0.41034f
C131 VP.n16 B 1.49954f
C132 VP.t0 B 0.950934f
C133 VP.n17 B 0.41034f
C134 VP.n18 B 1.5322f
C135 VP.n19 B 0.049917f
C136 VP.n20 B 0.037409f
C137 VP.n21 B 0.036512f
C138 VP.n22 B 0.342943f
C139 VP.n23 B 0.05381f
C140 VP.n24 B 0.05381f
C141 VP.n25 B 0.037409f
C142 VP.n26 B 0.037409f
C143 VP.n27 B 0.036512f
C144 VP.n28 B 0.050095f
C145 VP.t1 B 0.950934f
C146 VP.n29 B 0.41034f
C147 VP.n30 B 0.035035f
.ends

