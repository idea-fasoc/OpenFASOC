* NGSPICE file created from diff_pair_sample_0345.ext - technology: sky130A

.subckt diff_pair_sample_0345 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t13 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X1 B.t11 B.t9 B.t10 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0 ps=0 w=3.41 l=3.82
X2 B.t8 B.t6 B.t7 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0 ps=0 w=3.41 l=3.82
X3 VTAIL.t7 VN.t0 VDD2.t9 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X4 VTAIL.t3 VN.t1 VDD2.t8 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X5 VDD1.t8 VP.t1 VTAIL.t19 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=1.3299 ps=7.6 w=3.41 l=3.82
X6 VTAIL.t1 VN.t2 VDD2.t7 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X7 VDD1.t7 VP.t2 VTAIL.t17 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0.56265 ps=3.74 w=3.41 l=3.82
X8 VDD1.t6 VP.t3 VTAIL.t11 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X9 VTAIL.t12 VP.t4 VDD1.t5 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X10 VDD2.t6 VN.t3 VTAIL.t2 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=1.3299 ps=7.6 w=3.41 l=3.82
X11 VDD1.t4 VP.t5 VTAIL.t18 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=1.3299 ps=7.6 w=3.41 l=3.82
X12 VDD2.t5 VN.t4 VTAIL.t6 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X13 VDD2.t4 VN.t5 VTAIL.t9 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X14 VDD2.t3 VN.t6 VTAIL.t0 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0.56265 ps=3.74 w=3.41 l=3.82
X15 B.t5 B.t3 B.t4 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0 ps=0 w=3.41 l=3.82
X16 VTAIL.t10 VP.t6 VDD1.t3 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X17 VDD2.t2 VN.t7 VTAIL.t8 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0.56265 ps=3.74 w=3.41 l=3.82
X18 VDD2.t1 VN.t8 VTAIL.t5 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=1.3299 ps=7.6 w=3.41 l=3.82
X19 VDD1.t2 VP.t7 VTAIL.t16 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0.56265 ps=3.74 w=3.41 l=3.82
X20 VTAIL.t15 VP.t8 VDD1.t1 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X21 VTAIL.t14 VP.t9 VDD1.t0 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X22 VTAIL.t4 VN.t9 VDD2.t0 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=0.56265 pd=3.74 as=0.56265 ps=3.74 w=3.41 l=3.82
X23 B.t2 B.t0 B.t1 w_n5950_n1650# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=7.6 as=0 ps=0 w=3.41 l=3.82
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n75 VP.n74 87.6207
R60 VP.n130 VP.n0 87.6207
R61 VP.n73 VP.n18 87.6207
R62 VP.n96 VP.n95 56.5193
R63 VP.n109 VP.n108 56.5193
R64 VP.n52 VP.n51 56.5193
R65 VP.n39 VP.n38 56.5193
R66 VP.n32 VP.n31 55.4712
R67 VP.n31 VP.t7 54.2692
R68 VP.n74 VP.n73 53.291
R69 VP.n83 VP.n82 42.9216
R70 VP.n122 VP.n121 42.9216
R71 VP.n65 VP.n64 42.9216
R72 VP.n82 VP.n81 38.0652
R73 VP.n122 VP.n2 38.0652
R74 VP.n65 VP.n20 38.0652
R75 VP.n77 VP.n76 24.4675
R76 VP.n77 VP.n16 24.4675
R77 VP.n81 VP.n16 24.4675
R78 VP.n83 VP.n14 24.4675
R79 VP.n87 VP.n14 24.4675
R80 VP.n88 VP.n87 24.4675
R81 VP.n90 VP.n12 24.4675
R82 VP.n94 VP.n12 24.4675
R83 VP.n95 VP.n94 24.4675
R84 VP.n96 VP.n10 24.4675
R85 VP.n100 VP.n10 24.4675
R86 VP.n101 VP.n100 24.4675
R87 VP.n103 VP.n8 24.4675
R88 VP.n107 VP.n8 24.4675
R89 VP.n108 VP.n107 24.4675
R90 VP.n109 VP.n6 24.4675
R91 VP.n113 VP.n6 24.4675
R92 VP.n114 VP.n113 24.4675
R93 VP.n116 VP.n4 24.4675
R94 VP.n120 VP.n4 24.4675
R95 VP.n121 VP.n120 24.4675
R96 VP.n126 VP.n2 24.4675
R97 VP.n127 VP.n126 24.4675
R98 VP.n128 VP.n127 24.4675
R99 VP.n69 VP.n20 24.4675
R100 VP.n70 VP.n69 24.4675
R101 VP.n71 VP.n70 24.4675
R102 VP.n52 VP.n24 24.4675
R103 VP.n56 VP.n24 24.4675
R104 VP.n57 VP.n56 24.4675
R105 VP.n59 VP.n22 24.4675
R106 VP.n63 VP.n22 24.4675
R107 VP.n64 VP.n63 24.4675
R108 VP.n39 VP.n28 24.4675
R109 VP.n43 VP.n28 24.4675
R110 VP.n44 VP.n43 24.4675
R111 VP.n46 VP.n26 24.4675
R112 VP.n50 VP.n26 24.4675
R113 VP.n51 VP.n50 24.4675
R114 VP.n33 VP.n30 24.4675
R115 VP.n37 VP.n30 24.4675
R116 VP.n38 VP.n37 24.4675
R117 VP.n75 VP.t2 21.5139
R118 VP.n89 VP.t9 21.5139
R119 VP.n102 VP.t3 21.5139
R120 VP.n115 VP.t8 21.5139
R121 VP.n0 VP.t1 21.5139
R122 VP.n18 VP.t5 21.5139
R123 VP.n58 VP.t6 21.5139
R124 VP.n45 VP.t0 21.5139
R125 VP.n32 VP.t4 21.5139
R126 VP.n90 VP.n89 19.5741
R127 VP.n115 VP.n114 19.5741
R128 VP.n58 VP.n57 19.5741
R129 VP.n33 VP.n32 19.5741
R130 VP.n102 VP.n101 12.234
R131 VP.n103 VP.n102 12.234
R132 VP.n45 VP.n44 12.234
R133 VP.n46 VP.n45 12.234
R134 VP.n89 VP.n88 4.8939
R135 VP.n116 VP.n115 4.8939
R136 VP.n59 VP.n58 4.8939
R137 VP.n34 VP.n31 2.47313
R138 VP.n76 VP.n75 2.4472
R139 VP.n128 VP.n0 2.4472
R140 VP.n71 VP.n18 2.4472
R141 VP.n73 VP.n72 0.354971
R142 VP.n74 VP.n17 0.354971
R143 VP.n130 VP.n129 0.354971
R144 VP VP.n130 0.26696
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n11 VTAIL.t2 111.404
R203 VTAIL.n17 VTAIL.t5 111.404
R204 VTAIL.n2 VTAIL.t19 111.404
R205 VTAIL.n16 VTAIL.t18 111.404
R206 VTAIL.n15 VTAIL.n14 101.871
R207 VTAIL.n13 VTAIL.n12 101.871
R208 VTAIL.n10 VTAIL.n9 101.871
R209 VTAIL.n8 VTAIL.n7 101.871
R210 VTAIL.n19 VTAIL.n18 101.871
R211 VTAIL.n1 VTAIL.n0 101.871
R212 VTAIL.n4 VTAIL.n3 101.871
R213 VTAIL.n6 VTAIL.n5 101.871
R214 VTAIL.n8 VTAIL.n6 22.4617
R215 VTAIL.n17 VTAIL.n16 18.8841
R216 VTAIL.n18 VTAIL.t9 9.53276
R217 VTAIL.n18 VTAIL.t4 9.53276
R218 VTAIL.n0 VTAIL.t0 9.53276
R219 VTAIL.n0 VTAIL.t7 9.53276
R220 VTAIL.n3 VTAIL.t11 9.53276
R221 VTAIL.n3 VTAIL.t15 9.53276
R222 VTAIL.n5 VTAIL.t17 9.53276
R223 VTAIL.n5 VTAIL.t14 9.53276
R224 VTAIL.n14 VTAIL.t13 9.53276
R225 VTAIL.n14 VTAIL.t10 9.53276
R226 VTAIL.n12 VTAIL.t16 9.53276
R227 VTAIL.n12 VTAIL.t12 9.53276
R228 VTAIL.n9 VTAIL.t6 9.53276
R229 VTAIL.n9 VTAIL.t1 9.53276
R230 VTAIL.n7 VTAIL.t8 9.53276
R231 VTAIL.n7 VTAIL.t3 9.53276
R232 VTAIL.n10 VTAIL.n8 3.57809
R233 VTAIL.n11 VTAIL.n10 3.57809
R234 VTAIL.n15 VTAIL.n13 3.57809
R235 VTAIL.n16 VTAIL.n15 3.57809
R236 VTAIL.n6 VTAIL.n4 3.57809
R237 VTAIL.n4 VTAIL.n2 3.57809
R238 VTAIL.n19 VTAIL.n17 3.57809
R239 VTAIL VTAIL.n1 2.74188
R240 VTAIL.n13 VTAIL.n11 2.25912
R241 VTAIL.n2 VTAIL.n1 2.25912
R242 VTAIL VTAIL.n19 0.836707
R243 VDD1.n1 VDD1.t2 131.661
R244 VDD1.n3 VDD1.t7 131.661
R245 VDD1.n5 VDD1.n4 121.178
R246 VDD1.n1 VDD1.n0 118.55
R247 VDD1.n7 VDD1.n6 118.55
R248 VDD1.n3 VDD1.n2 118.55
R249 VDD1.n7 VDD1.n5 46.0203
R250 VDD1.n6 VDD1.t3 9.53276
R251 VDD1.n6 VDD1.t4 9.53276
R252 VDD1.n0 VDD1.t5 9.53276
R253 VDD1.n0 VDD1.t9 9.53276
R254 VDD1.n4 VDD1.t1 9.53276
R255 VDD1.n4 VDD1.t8 9.53276
R256 VDD1.n2 VDD1.t0 9.53276
R257 VDD1.n2 VDD1.t6 9.53276
R258 VDD1 VDD1.n7 2.6255
R259 VDD1 VDD1.n1 0.953086
R260 VDD1.n5 VDD1.n3 0.839551
R261 B.n400 B.n399 585
R262 B.n398 B.n151 585
R263 B.n397 B.n396 585
R264 B.n395 B.n152 585
R265 B.n394 B.n393 585
R266 B.n392 B.n153 585
R267 B.n391 B.n390 585
R268 B.n389 B.n154 585
R269 B.n388 B.n387 585
R270 B.n386 B.n155 585
R271 B.n385 B.n384 585
R272 B.n383 B.n156 585
R273 B.n382 B.n381 585
R274 B.n380 B.n157 585
R275 B.n379 B.n378 585
R276 B.n377 B.n158 585
R277 B.n375 B.n374 585
R278 B.n373 B.n161 585
R279 B.n372 B.n371 585
R280 B.n370 B.n162 585
R281 B.n369 B.n368 585
R282 B.n367 B.n163 585
R283 B.n366 B.n365 585
R284 B.n364 B.n164 585
R285 B.n363 B.n362 585
R286 B.n361 B.n165 585
R287 B.n360 B.n359 585
R288 B.n355 B.n166 585
R289 B.n354 B.n353 585
R290 B.n352 B.n167 585
R291 B.n351 B.n350 585
R292 B.n349 B.n168 585
R293 B.n348 B.n347 585
R294 B.n346 B.n169 585
R295 B.n345 B.n344 585
R296 B.n343 B.n170 585
R297 B.n342 B.n341 585
R298 B.n340 B.n171 585
R299 B.n339 B.n338 585
R300 B.n337 B.n172 585
R301 B.n336 B.n335 585
R302 B.n334 B.n173 585
R303 B.n401 B.n150 585
R304 B.n403 B.n402 585
R305 B.n404 B.n149 585
R306 B.n406 B.n405 585
R307 B.n407 B.n148 585
R308 B.n409 B.n408 585
R309 B.n410 B.n147 585
R310 B.n412 B.n411 585
R311 B.n413 B.n146 585
R312 B.n415 B.n414 585
R313 B.n416 B.n145 585
R314 B.n418 B.n417 585
R315 B.n419 B.n144 585
R316 B.n421 B.n420 585
R317 B.n422 B.n143 585
R318 B.n424 B.n423 585
R319 B.n425 B.n142 585
R320 B.n427 B.n426 585
R321 B.n428 B.n141 585
R322 B.n430 B.n429 585
R323 B.n431 B.n140 585
R324 B.n433 B.n432 585
R325 B.n434 B.n139 585
R326 B.n436 B.n435 585
R327 B.n437 B.n138 585
R328 B.n439 B.n438 585
R329 B.n440 B.n137 585
R330 B.n442 B.n441 585
R331 B.n443 B.n136 585
R332 B.n445 B.n444 585
R333 B.n446 B.n135 585
R334 B.n448 B.n447 585
R335 B.n449 B.n134 585
R336 B.n451 B.n450 585
R337 B.n452 B.n133 585
R338 B.n454 B.n453 585
R339 B.n455 B.n132 585
R340 B.n457 B.n456 585
R341 B.n458 B.n131 585
R342 B.n460 B.n459 585
R343 B.n461 B.n130 585
R344 B.n463 B.n462 585
R345 B.n464 B.n129 585
R346 B.n466 B.n465 585
R347 B.n467 B.n128 585
R348 B.n469 B.n468 585
R349 B.n470 B.n127 585
R350 B.n472 B.n471 585
R351 B.n473 B.n126 585
R352 B.n475 B.n474 585
R353 B.n476 B.n125 585
R354 B.n478 B.n477 585
R355 B.n479 B.n124 585
R356 B.n481 B.n480 585
R357 B.n482 B.n123 585
R358 B.n484 B.n483 585
R359 B.n485 B.n122 585
R360 B.n487 B.n486 585
R361 B.n488 B.n121 585
R362 B.n490 B.n489 585
R363 B.n491 B.n120 585
R364 B.n493 B.n492 585
R365 B.n494 B.n119 585
R366 B.n496 B.n495 585
R367 B.n497 B.n118 585
R368 B.n499 B.n498 585
R369 B.n500 B.n117 585
R370 B.n502 B.n501 585
R371 B.n503 B.n116 585
R372 B.n505 B.n504 585
R373 B.n506 B.n115 585
R374 B.n508 B.n507 585
R375 B.n509 B.n114 585
R376 B.n511 B.n510 585
R377 B.n512 B.n113 585
R378 B.n514 B.n513 585
R379 B.n515 B.n112 585
R380 B.n517 B.n516 585
R381 B.n518 B.n111 585
R382 B.n520 B.n519 585
R383 B.n521 B.n110 585
R384 B.n523 B.n522 585
R385 B.n524 B.n109 585
R386 B.n526 B.n525 585
R387 B.n527 B.n108 585
R388 B.n529 B.n528 585
R389 B.n530 B.n107 585
R390 B.n532 B.n531 585
R391 B.n533 B.n106 585
R392 B.n535 B.n534 585
R393 B.n536 B.n105 585
R394 B.n538 B.n537 585
R395 B.n539 B.n104 585
R396 B.n541 B.n540 585
R397 B.n542 B.n103 585
R398 B.n544 B.n543 585
R399 B.n545 B.n102 585
R400 B.n547 B.n546 585
R401 B.n548 B.n101 585
R402 B.n550 B.n549 585
R403 B.n551 B.n100 585
R404 B.n553 B.n552 585
R405 B.n554 B.n99 585
R406 B.n556 B.n555 585
R407 B.n557 B.n98 585
R408 B.n559 B.n558 585
R409 B.n560 B.n97 585
R410 B.n562 B.n561 585
R411 B.n563 B.n96 585
R412 B.n565 B.n564 585
R413 B.n566 B.n95 585
R414 B.n568 B.n567 585
R415 B.n569 B.n94 585
R416 B.n571 B.n570 585
R417 B.n572 B.n93 585
R418 B.n574 B.n573 585
R419 B.n575 B.n92 585
R420 B.n577 B.n576 585
R421 B.n578 B.n91 585
R422 B.n580 B.n579 585
R423 B.n581 B.n90 585
R424 B.n583 B.n582 585
R425 B.n584 B.n89 585
R426 B.n586 B.n585 585
R427 B.n587 B.n88 585
R428 B.n589 B.n588 585
R429 B.n590 B.n87 585
R430 B.n592 B.n591 585
R431 B.n593 B.n86 585
R432 B.n595 B.n594 585
R433 B.n596 B.n85 585
R434 B.n598 B.n597 585
R435 B.n599 B.n84 585
R436 B.n601 B.n600 585
R437 B.n602 B.n83 585
R438 B.n604 B.n603 585
R439 B.n605 B.n82 585
R440 B.n607 B.n606 585
R441 B.n608 B.n81 585
R442 B.n610 B.n609 585
R443 B.n611 B.n80 585
R444 B.n613 B.n612 585
R445 B.n614 B.n79 585
R446 B.n616 B.n615 585
R447 B.n617 B.n78 585
R448 B.n619 B.n618 585
R449 B.n620 B.n77 585
R450 B.n622 B.n621 585
R451 B.n623 B.n76 585
R452 B.n625 B.n624 585
R453 B.n626 B.n75 585
R454 B.n628 B.n627 585
R455 B.n629 B.n74 585
R456 B.n631 B.n630 585
R457 B.n632 B.n73 585
R458 B.n634 B.n633 585
R459 B.n635 B.n72 585
R460 B.n637 B.n636 585
R461 B.n638 B.n71 585
R462 B.n640 B.n639 585
R463 B.n641 B.n70 585
R464 B.n643 B.n642 585
R465 B.n644 B.n69 585
R466 B.n646 B.n645 585
R467 B.n710 B.n709 585
R468 B.n708 B.n43 585
R469 B.n707 B.n706 585
R470 B.n705 B.n44 585
R471 B.n704 B.n703 585
R472 B.n702 B.n45 585
R473 B.n701 B.n700 585
R474 B.n699 B.n46 585
R475 B.n698 B.n697 585
R476 B.n696 B.n47 585
R477 B.n695 B.n694 585
R478 B.n693 B.n48 585
R479 B.n692 B.n691 585
R480 B.n690 B.n49 585
R481 B.n689 B.n688 585
R482 B.n687 B.n50 585
R483 B.n686 B.n685 585
R484 B.n684 B.n51 585
R485 B.n683 B.n682 585
R486 B.n681 B.n55 585
R487 B.n680 B.n679 585
R488 B.n678 B.n56 585
R489 B.n677 B.n676 585
R490 B.n675 B.n57 585
R491 B.n674 B.n673 585
R492 B.n672 B.n58 585
R493 B.n670 B.n669 585
R494 B.n668 B.n61 585
R495 B.n667 B.n666 585
R496 B.n665 B.n62 585
R497 B.n664 B.n663 585
R498 B.n662 B.n63 585
R499 B.n661 B.n660 585
R500 B.n659 B.n64 585
R501 B.n658 B.n657 585
R502 B.n656 B.n65 585
R503 B.n655 B.n654 585
R504 B.n653 B.n66 585
R505 B.n652 B.n651 585
R506 B.n650 B.n67 585
R507 B.n649 B.n648 585
R508 B.n647 B.n68 585
R509 B.n711 B.n42 585
R510 B.n713 B.n712 585
R511 B.n714 B.n41 585
R512 B.n716 B.n715 585
R513 B.n717 B.n40 585
R514 B.n719 B.n718 585
R515 B.n720 B.n39 585
R516 B.n722 B.n721 585
R517 B.n723 B.n38 585
R518 B.n725 B.n724 585
R519 B.n726 B.n37 585
R520 B.n728 B.n727 585
R521 B.n729 B.n36 585
R522 B.n731 B.n730 585
R523 B.n732 B.n35 585
R524 B.n734 B.n733 585
R525 B.n735 B.n34 585
R526 B.n737 B.n736 585
R527 B.n738 B.n33 585
R528 B.n740 B.n739 585
R529 B.n741 B.n32 585
R530 B.n743 B.n742 585
R531 B.n744 B.n31 585
R532 B.n746 B.n745 585
R533 B.n747 B.n30 585
R534 B.n749 B.n748 585
R535 B.n750 B.n29 585
R536 B.n752 B.n751 585
R537 B.n753 B.n28 585
R538 B.n755 B.n754 585
R539 B.n756 B.n27 585
R540 B.n758 B.n757 585
R541 B.n759 B.n26 585
R542 B.n761 B.n760 585
R543 B.n762 B.n25 585
R544 B.n764 B.n763 585
R545 B.n765 B.n24 585
R546 B.n767 B.n766 585
R547 B.n768 B.n23 585
R548 B.n770 B.n769 585
R549 B.n771 B.n22 585
R550 B.n773 B.n772 585
R551 B.n774 B.n21 585
R552 B.n776 B.n775 585
R553 B.n777 B.n20 585
R554 B.n779 B.n778 585
R555 B.n780 B.n19 585
R556 B.n782 B.n781 585
R557 B.n783 B.n18 585
R558 B.n785 B.n784 585
R559 B.n786 B.n17 585
R560 B.n788 B.n787 585
R561 B.n789 B.n16 585
R562 B.n791 B.n790 585
R563 B.n792 B.n15 585
R564 B.n794 B.n793 585
R565 B.n795 B.n14 585
R566 B.n797 B.n796 585
R567 B.n798 B.n13 585
R568 B.n800 B.n799 585
R569 B.n801 B.n12 585
R570 B.n803 B.n802 585
R571 B.n804 B.n11 585
R572 B.n806 B.n805 585
R573 B.n807 B.n10 585
R574 B.n809 B.n808 585
R575 B.n810 B.n9 585
R576 B.n812 B.n811 585
R577 B.n813 B.n8 585
R578 B.n815 B.n814 585
R579 B.n816 B.n7 585
R580 B.n818 B.n817 585
R581 B.n819 B.n6 585
R582 B.n821 B.n820 585
R583 B.n822 B.n5 585
R584 B.n824 B.n823 585
R585 B.n825 B.n4 585
R586 B.n827 B.n826 585
R587 B.n828 B.n3 585
R588 B.n830 B.n829 585
R589 B.n831 B.n0 585
R590 B.n2 B.n1 585
R591 B.n214 B.n213 585
R592 B.n216 B.n215 585
R593 B.n217 B.n212 585
R594 B.n219 B.n218 585
R595 B.n220 B.n211 585
R596 B.n222 B.n221 585
R597 B.n223 B.n210 585
R598 B.n225 B.n224 585
R599 B.n226 B.n209 585
R600 B.n228 B.n227 585
R601 B.n229 B.n208 585
R602 B.n231 B.n230 585
R603 B.n232 B.n207 585
R604 B.n234 B.n233 585
R605 B.n235 B.n206 585
R606 B.n237 B.n236 585
R607 B.n238 B.n205 585
R608 B.n240 B.n239 585
R609 B.n241 B.n204 585
R610 B.n243 B.n242 585
R611 B.n244 B.n203 585
R612 B.n246 B.n245 585
R613 B.n247 B.n202 585
R614 B.n249 B.n248 585
R615 B.n250 B.n201 585
R616 B.n252 B.n251 585
R617 B.n253 B.n200 585
R618 B.n255 B.n254 585
R619 B.n256 B.n199 585
R620 B.n258 B.n257 585
R621 B.n259 B.n198 585
R622 B.n261 B.n260 585
R623 B.n262 B.n197 585
R624 B.n264 B.n263 585
R625 B.n265 B.n196 585
R626 B.n267 B.n266 585
R627 B.n268 B.n195 585
R628 B.n270 B.n269 585
R629 B.n271 B.n194 585
R630 B.n273 B.n272 585
R631 B.n274 B.n193 585
R632 B.n276 B.n275 585
R633 B.n277 B.n192 585
R634 B.n279 B.n278 585
R635 B.n280 B.n191 585
R636 B.n282 B.n281 585
R637 B.n283 B.n190 585
R638 B.n285 B.n284 585
R639 B.n286 B.n189 585
R640 B.n288 B.n287 585
R641 B.n289 B.n188 585
R642 B.n291 B.n290 585
R643 B.n292 B.n187 585
R644 B.n294 B.n293 585
R645 B.n295 B.n186 585
R646 B.n297 B.n296 585
R647 B.n298 B.n185 585
R648 B.n300 B.n299 585
R649 B.n301 B.n184 585
R650 B.n303 B.n302 585
R651 B.n304 B.n183 585
R652 B.n306 B.n305 585
R653 B.n307 B.n182 585
R654 B.n309 B.n308 585
R655 B.n310 B.n181 585
R656 B.n312 B.n311 585
R657 B.n313 B.n180 585
R658 B.n315 B.n314 585
R659 B.n316 B.n179 585
R660 B.n318 B.n317 585
R661 B.n319 B.n178 585
R662 B.n321 B.n320 585
R663 B.n322 B.n177 585
R664 B.n324 B.n323 585
R665 B.n325 B.n176 585
R666 B.n327 B.n326 585
R667 B.n328 B.n175 585
R668 B.n330 B.n329 585
R669 B.n331 B.n174 585
R670 B.n333 B.n332 585
R671 B.n334 B.n333 497.305
R672 B.n399 B.n150 497.305
R673 B.n645 B.n68 497.305
R674 B.n711 B.n710 497.305
R675 B.n833 B.n832 256.663
R676 B.n832 B.n831 235.042
R677 B.n832 B.n2 235.042
R678 B.n356 B.t3 230.873
R679 B.n159 B.t6 230.873
R680 B.n59 B.t0 230.873
R681 B.n52 B.t9 230.873
R682 B.n159 B.t7 207.28
R683 B.n59 B.t2 207.28
R684 B.n356 B.t4 207.276
R685 B.n52 B.t11 207.276
R686 B.n335 B.n334 163.367
R687 B.n335 B.n172 163.367
R688 B.n339 B.n172 163.367
R689 B.n340 B.n339 163.367
R690 B.n341 B.n340 163.367
R691 B.n341 B.n170 163.367
R692 B.n345 B.n170 163.367
R693 B.n346 B.n345 163.367
R694 B.n347 B.n346 163.367
R695 B.n347 B.n168 163.367
R696 B.n351 B.n168 163.367
R697 B.n352 B.n351 163.367
R698 B.n353 B.n352 163.367
R699 B.n353 B.n166 163.367
R700 B.n360 B.n166 163.367
R701 B.n361 B.n360 163.367
R702 B.n362 B.n361 163.367
R703 B.n362 B.n164 163.367
R704 B.n366 B.n164 163.367
R705 B.n367 B.n366 163.367
R706 B.n368 B.n367 163.367
R707 B.n368 B.n162 163.367
R708 B.n372 B.n162 163.367
R709 B.n373 B.n372 163.367
R710 B.n374 B.n373 163.367
R711 B.n374 B.n158 163.367
R712 B.n379 B.n158 163.367
R713 B.n380 B.n379 163.367
R714 B.n381 B.n380 163.367
R715 B.n381 B.n156 163.367
R716 B.n385 B.n156 163.367
R717 B.n386 B.n385 163.367
R718 B.n387 B.n386 163.367
R719 B.n387 B.n154 163.367
R720 B.n391 B.n154 163.367
R721 B.n392 B.n391 163.367
R722 B.n393 B.n392 163.367
R723 B.n393 B.n152 163.367
R724 B.n397 B.n152 163.367
R725 B.n398 B.n397 163.367
R726 B.n399 B.n398 163.367
R727 B.n645 B.n644 163.367
R728 B.n644 B.n643 163.367
R729 B.n643 B.n70 163.367
R730 B.n639 B.n70 163.367
R731 B.n639 B.n638 163.367
R732 B.n638 B.n637 163.367
R733 B.n637 B.n72 163.367
R734 B.n633 B.n72 163.367
R735 B.n633 B.n632 163.367
R736 B.n632 B.n631 163.367
R737 B.n631 B.n74 163.367
R738 B.n627 B.n74 163.367
R739 B.n627 B.n626 163.367
R740 B.n626 B.n625 163.367
R741 B.n625 B.n76 163.367
R742 B.n621 B.n76 163.367
R743 B.n621 B.n620 163.367
R744 B.n620 B.n619 163.367
R745 B.n619 B.n78 163.367
R746 B.n615 B.n78 163.367
R747 B.n615 B.n614 163.367
R748 B.n614 B.n613 163.367
R749 B.n613 B.n80 163.367
R750 B.n609 B.n80 163.367
R751 B.n609 B.n608 163.367
R752 B.n608 B.n607 163.367
R753 B.n607 B.n82 163.367
R754 B.n603 B.n82 163.367
R755 B.n603 B.n602 163.367
R756 B.n602 B.n601 163.367
R757 B.n601 B.n84 163.367
R758 B.n597 B.n84 163.367
R759 B.n597 B.n596 163.367
R760 B.n596 B.n595 163.367
R761 B.n595 B.n86 163.367
R762 B.n591 B.n86 163.367
R763 B.n591 B.n590 163.367
R764 B.n590 B.n589 163.367
R765 B.n589 B.n88 163.367
R766 B.n585 B.n88 163.367
R767 B.n585 B.n584 163.367
R768 B.n584 B.n583 163.367
R769 B.n583 B.n90 163.367
R770 B.n579 B.n90 163.367
R771 B.n579 B.n578 163.367
R772 B.n578 B.n577 163.367
R773 B.n577 B.n92 163.367
R774 B.n573 B.n92 163.367
R775 B.n573 B.n572 163.367
R776 B.n572 B.n571 163.367
R777 B.n571 B.n94 163.367
R778 B.n567 B.n94 163.367
R779 B.n567 B.n566 163.367
R780 B.n566 B.n565 163.367
R781 B.n565 B.n96 163.367
R782 B.n561 B.n96 163.367
R783 B.n561 B.n560 163.367
R784 B.n560 B.n559 163.367
R785 B.n559 B.n98 163.367
R786 B.n555 B.n98 163.367
R787 B.n555 B.n554 163.367
R788 B.n554 B.n553 163.367
R789 B.n553 B.n100 163.367
R790 B.n549 B.n100 163.367
R791 B.n549 B.n548 163.367
R792 B.n548 B.n547 163.367
R793 B.n547 B.n102 163.367
R794 B.n543 B.n102 163.367
R795 B.n543 B.n542 163.367
R796 B.n542 B.n541 163.367
R797 B.n541 B.n104 163.367
R798 B.n537 B.n104 163.367
R799 B.n537 B.n536 163.367
R800 B.n536 B.n535 163.367
R801 B.n535 B.n106 163.367
R802 B.n531 B.n106 163.367
R803 B.n531 B.n530 163.367
R804 B.n530 B.n529 163.367
R805 B.n529 B.n108 163.367
R806 B.n525 B.n108 163.367
R807 B.n525 B.n524 163.367
R808 B.n524 B.n523 163.367
R809 B.n523 B.n110 163.367
R810 B.n519 B.n110 163.367
R811 B.n519 B.n518 163.367
R812 B.n518 B.n517 163.367
R813 B.n517 B.n112 163.367
R814 B.n513 B.n112 163.367
R815 B.n513 B.n512 163.367
R816 B.n512 B.n511 163.367
R817 B.n511 B.n114 163.367
R818 B.n507 B.n114 163.367
R819 B.n507 B.n506 163.367
R820 B.n506 B.n505 163.367
R821 B.n505 B.n116 163.367
R822 B.n501 B.n116 163.367
R823 B.n501 B.n500 163.367
R824 B.n500 B.n499 163.367
R825 B.n499 B.n118 163.367
R826 B.n495 B.n118 163.367
R827 B.n495 B.n494 163.367
R828 B.n494 B.n493 163.367
R829 B.n493 B.n120 163.367
R830 B.n489 B.n120 163.367
R831 B.n489 B.n488 163.367
R832 B.n488 B.n487 163.367
R833 B.n487 B.n122 163.367
R834 B.n483 B.n122 163.367
R835 B.n483 B.n482 163.367
R836 B.n482 B.n481 163.367
R837 B.n481 B.n124 163.367
R838 B.n477 B.n124 163.367
R839 B.n477 B.n476 163.367
R840 B.n476 B.n475 163.367
R841 B.n475 B.n126 163.367
R842 B.n471 B.n126 163.367
R843 B.n471 B.n470 163.367
R844 B.n470 B.n469 163.367
R845 B.n469 B.n128 163.367
R846 B.n465 B.n128 163.367
R847 B.n465 B.n464 163.367
R848 B.n464 B.n463 163.367
R849 B.n463 B.n130 163.367
R850 B.n459 B.n130 163.367
R851 B.n459 B.n458 163.367
R852 B.n458 B.n457 163.367
R853 B.n457 B.n132 163.367
R854 B.n453 B.n132 163.367
R855 B.n453 B.n452 163.367
R856 B.n452 B.n451 163.367
R857 B.n451 B.n134 163.367
R858 B.n447 B.n134 163.367
R859 B.n447 B.n446 163.367
R860 B.n446 B.n445 163.367
R861 B.n445 B.n136 163.367
R862 B.n441 B.n136 163.367
R863 B.n441 B.n440 163.367
R864 B.n440 B.n439 163.367
R865 B.n439 B.n138 163.367
R866 B.n435 B.n138 163.367
R867 B.n435 B.n434 163.367
R868 B.n434 B.n433 163.367
R869 B.n433 B.n140 163.367
R870 B.n429 B.n140 163.367
R871 B.n429 B.n428 163.367
R872 B.n428 B.n427 163.367
R873 B.n427 B.n142 163.367
R874 B.n423 B.n142 163.367
R875 B.n423 B.n422 163.367
R876 B.n422 B.n421 163.367
R877 B.n421 B.n144 163.367
R878 B.n417 B.n144 163.367
R879 B.n417 B.n416 163.367
R880 B.n416 B.n415 163.367
R881 B.n415 B.n146 163.367
R882 B.n411 B.n146 163.367
R883 B.n411 B.n410 163.367
R884 B.n410 B.n409 163.367
R885 B.n409 B.n148 163.367
R886 B.n405 B.n148 163.367
R887 B.n405 B.n404 163.367
R888 B.n404 B.n403 163.367
R889 B.n403 B.n150 163.367
R890 B.n710 B.n43 163.367
R891 B.n706 B.n43 163.367
R892 B.n706 B.n705 163.367
R893 B.n705 B.n704 163.367
R894 B.n704 B.n45 163.367
R895 B.n700 B.n45 163.367
R896 B.n700 B.n699 163.367
R897 B.n699 B.n698 163.367
R898 B.n698 B.n47 163.367
R899 B.n694 B.n47 163.367
R900 B.n694 B.n693 163.367
R901 B.n693 B.n692 163.367
R902 B.n692 B.n49 163.367
R903 B.n688 B.n49 163.367
R904 B.n688 B.n687 163.367
R905 B.n687 B.n686 163.367
R906 B.n686 B.n51 163.367
R907 B.n682 B.n51 163.367
R908 B.n682 B.n681 163.367
R909 B.n681 B.n680 163.367
R910 B.n680 B.n56 163.367
R911 B.n676 B.n56 163.367
R912 B.n676 B.n675 163.367
R913 B.n675 B.n674 163.367
R914 B.n674 B.n58 163.367
R915 B.n669 B.n58 163.367
R916 B.n669 B.n668 163.367
R917 B.n668 B.n667 163.367
R918 B.n667 B.n62 163.367
R919 B.n663 B.n62 163.367
R920 B.n663 B.n662 163.367
R921 B.n662 B.n661 163.367
R922 B.n661 B.n64 163.367
R923 B.n657 B.n64 163.367
R924 B.n657 B.n656 163.367
R925 B.n656 B.n655 163.367
R926 B.n655 B.n66 163.367
R927 B.n651 B.n66 163.367
R928 B.n651 B.n650 163.367
R929 B.n650 B.n649 163.367
R930 B.n649 B.n68 163.367
R931 B.n712 B.n711 163.367
R932 B.n712 B.n41 163.367
R933 B.n716 B.n41 163.367
R934 B.n717 B.n716 163.367
R935 B.n718 B.n717 163.367
R936 B.n718 B.n39 163.367
R937 B.n722 B.n39 163.367
R938 B.n723 B.n722 163.367
R939 B.n724 B.n723 163.367
R940 B.n724 B.n37 163.367
R941 B.n728 B.n37 163.367
R942 B.n729 B.n728 163.367
R943 B.n730 B.n729 163.367
R944 B.n730 B.n35 163.367
R945 B.n734 B.n35 163.367
R946 B.n735 B.n734 163.367
R947 B.n736 B.n735 163.367
R948 B.n736 B.n33 163.367
R949 B.n740 B.n33 163.367
R950 B.n741 B.n740 163.367
R951 B.n742 B.n741 163.367
R952 B.n742 B.n31 163.367
R953 B.n746 B.n31 163.367
R954 B.n747 B.n746 163.367
R955 B.n748 B.n747 163.367
R956 B.n748 B.n29 163.367
R957 B.n752 B.n29 163.367
R958 B.n753 B.n752 163.367
R959 B.n754 B.n753 163.367
R960 B.n754 B.n27 163.367
R961 B.n758 B.n27 163.367
R962 B.n759 B.n758 163.367
R963 B.n760 B.n759 163.367
R964 B.n760 B.n25 163.367
R965 B.n764 B.n25 163.367
R966 B.n765 B.n764 163.367
R967 B.n766 B.n765 163.367
R968 B.n766 B.n23 163.367
R969 B.n770 B.n23 163.367
R970 B.n771 B.n770 163.367
R971 B.n772 B.n771 163.367
R972 B.n772 B.n21 163.367
R973 B.n776 B.n21 163.367
R974 B.n777 B.n776 163.367
R975 B.n778 B.n777 163.367
R976 B.n778 B.n19 163.367
R977 B.n782 B.n19 163.367
R978 B.n783 B.n782 163.367
R979 B.n784 B.n783 163.367
R980 B.n784 B.n17 163.367
R981 B.n788 B.n17 163.367
R982 B.n789 B.n788 163.367
R983 B.n790 B.n789 163.367
R984 B.n790 B.n15 163.367
R985 B.n794 B.n15 163.367
R986 B.n795 B.n794 163.367
R987 B.n796 B.n795 163.367
R988 B.n796 B.n13 163.367
R989 B.n800 B.n13 163.367
R990 B.n801 B.n800 163.367
R991 B.n802 B.n801 163.367
R992 B.n802 B.n11 163.367
R993 B.n806 B.n11 163.367
R994 B.n807 B.n806 163.367
R995 B.n808 B.n807 163.367
R996 B.n808 B.n9 163.367
R997 B.n812 B.n9 163.367
R998 B.n813 B.n812 163.367
R999 B.n814 B.n813 163.367
R1000 B.n814 B.n7 163.367
R1001 B.n818 B.n7 163.367
R1002 B.n819 B.n818 163.367
R1003 B.n820 B.n819 163.367
R1004 B.n820 B.n5 163.367
R1005 B.n824 B.n5 163.367
R1006 B.n825 B.n824 163.367
R1007 B.n826 B.n825 163.367
R1008 B.n826 B.n3 163.367
R1009 B.n830 B.n3 163.367
R1010 B.n831 B.n830 163.367
R1011 B.n214 B.n2 163.367
R1012 B.n215 B.n214 163.367
R1013 B.n215 B.n212 163.367
R1014 B.n219 B.n212 163.367
R1015 B.n220 B.n219 163.367
R1016 B.n221 B.n220 163.367
R1017 B.n221 B.n210 163.367
R1018 B.n225 B.n210 163.367
R1019 B.n226 B.n225 163.367
R1020 B.n227 B.n226 163.367
R1021 B.n227 B.n208 163.367
R1022 B.n231 B.n208 163.367
R1023 B.n232 B.n231 163.367
R1024 B.n233 B.n232 163.367
R1025 B.n233 B.n206 163.367
R1026 B.n237 B.n206 163.367
R1027 B.n238 B.n237 163.367
R1028 B.n239 B.n238 163.367
R1029 B.n239 B.n204 163.367
R1030 B.n243 B.n204 163.367
R1031 B.n244 B.n243 163.367
R1032 B.n245 B.n244 163.367
R1033 B.n245 B.n202 163.367
R1034 B.n249 B.n202 163.367
R1035 B.n250 B.n249 163.367
R1036 B.n251 B.n250 163.367
R1037 B.n251 B.n200 163.367
R1038 B.n255 B.n200 163.367
R1039 B.n256 B.n255 163.367
R1040 B.n257 B.n256 163.367
R1041 B.n257 B.n198 163.367
R1042 B.n261 B.n198 163.367
R1043 B.n262 B.n261 163.367
R1044 B.n263 B.n262 163.367
R1045 B.n263 B.n196 163.367
R1046 B.n267 B.n196 163.367
R1047 B.n268 B.n267 163.367
R1048 B.n269 B.n268 163.367
R1049 B.n269 B.n194 163.367
R1050 B.n273 B.n194 163.367
R1051 B.n274 B.n273 163.367
R1052 B.n275 B.n274 163.367
R1053 B.n275 B.n192 163.367
R1054 B.n279 B.n192 163.367
R1055 B.n280 B.n279 163.367
R1056 B.n281 B.n280 163.367
R1057 B.n281 B.n190 163.367
R1058 B.n285 B.n190 163.367
R1059 B.n286 B.n285 163.367
R1060 B.n287 B.n286 163.367
R1061 B.n287 B.n188 163.367
R1062 B.n291 B.n188 163.367
R1063 B.n292 B.n291 163.367
R1064 B.n293 B.n292 163.367
R1065 B.n293 B.n186 163.367
R1066 B.n297 B.n186 163.367
R1067 B.n298 B.n297 163.367
R1068 B.n299 B.n298 163.367
R1069 B.n299 B.n184 163.367
R1070 B.n303 B.n184 163.367
R1071 B.n304 B.n303 163.367
R1072 B.n305 B.n304 163.367
R1073 B.n305 B.n182 163.367
R1074 B.n309 B.n182 163.367
R1075 B.n310 B.n309 163.367
R1076 B.n311 B.n310 163.367
R1077 B.n311 B.n180 163.367
R1078 B.n315 B.n180 163.367
R1079 B.n316 B.n315 163.367
R1080 B.n317 B.n316 163.367
R1081 B.n317 B.n178 163.367
R1082 B.n321 B.n178 163.367
R1083 B.n322 B.n321 163.367
R1084 B.n323 B.n322 163.367
R1085 B.n323 B.n176 163.367
R1086 B.n327 B.n176 163.367
R1087 B.n328 B.n327 163.367
R1088 B.n329 B.n328 163.367
R1089 B.n329 B.n174 163.367
R1090 B.n333 B.n174 163.367
R1091 B.n160 B.t8 126.794
R1092 B.n60 B.t1 126.794
R1093 B.n357 B.t5 126.793
R1094 B.n53 B.t10 126.793
R1095 B.n357 B.n356 80.4853
R1096 B.n160 B.n159 80.4853
R1097 B.n60 B.n59 80.4853
R1098 B.n53 B.n52 80.4853
R1099 B.n358 B.n357 59.5399
R1100 B.n376 B.n160 59.5399
R1101 B.n671 B.n60 59.5399
R1102 B.n54 B.n53 59.5399
R1103 B.n709 B.n42 32.3127
R1104 B.n647 B.n646 32.3127
R1105 B.n401 B.n400 32.3127
R1106 B.n332 B.n173 32.3127
R1107 B B.n833 18.0485
R1108 B.n713 B.n42 10.6151
R1109 B.n714 B.n713 10.6151
R1110 B.n715 B.n714 10.6151
R1111 B.n715 B.n40 10.6151
R1112 B.n719 B.n40 10.6151
R1113 B.n720 B.n719 10.6151
R1114 B.n721 B.n720 10.6151
R1115 B.n721 B.n38 10.6151
R1116 B.n725 B.n38 10.6151
R1117 B.n726 B.n725 10.6151
R1118 B.n727 B.n726 10.6151
R1119 B.n727 B.n36 10.6151
R1120 B.n731 B.n36 10.6151
R1121 B.n732 B.n731 10.6151
R1122 B.n733 B.n732 10.6151
R1123 B.n733 B.n34 10.6151
R1124 B.n737 B.n34 10.6151
R1125 B.n738 B.n737 10.6151
R1126 B.n739 B.n738 10.6151
R1127 B.n739 B.n32 10.6151
R1128 B.n743 B.n32 10.6151
R1129 B.n744 B.n743 10.6151
R1130 B.n745 B.n744 10.6151
R1131 B.n745 B.n30 10.6151
R1132 B.n749 B.n30 10.6151
R1133 B.n750 B.n749 10.6151
R1134 B.n751 B.n750 10.6151
R1135 B.n751 B.n28 10.6151
R1136 B.n755 B.n28 10.6151
R1137 B.n756 B.n755 10.6151
R1138 B.n757 B.n756 10.6151
R1139 B.n757 B.n26 10.6151
R1140 B.n761 B.n26 10.6151
R1141 B.n762 B.n761 10.6151
R1142 B.n763 B.n762 10.6151
R1143 B.n763 B.n24 10.6151
R1144 B.n767 B.n24 10.6151
R1145 B.n768 B.n767 10.6151
R1146 B.n769 B.n768 10.6151
R1147 B.n769 B.n22 10.6151
R1148 B.n773 B.n22 10.6151
R1149 B.n774 B.n773 10.6151
R1150 B.n775 B.n774 10.6151
R1151 B.n775 B.n20 10.6151
R1152 B.n779 B.n20 10.6151
R1153 B.n780 B.n779 10.6151
R1154 B.n781 B.n780 10.6151
R1155 B.n781 B.n18 10.6151
R1156 B.n785 B.n18 10.6151
R1157 B.n786 B.n785 10.6151
R1158 B.n787 B.n786 10.6151
R1159 B.n787 B.n16 10.6151
R1160 B.n791 B.n16 10.6151
R1161 B.n792 B.n791 10.6151
R1162 B.n793 B.n792 10.6151
R1163 B.n793 B.n14 10.6151
R1164 B.n797 B.n14 10.6151
R1165 B.n798 B.n797 10.6151
R1166 B.n799 B.n798 10.6151
R1167 B.n799 B.n12 10.6151
R1168 B.n803 B.n12 10.6151
R1169 B.n804 B.n803 10.6151
R1170 B.n805 B.n804 10.6151
R1171 B.n805 B.n10 10.6151
R1172 B.n809 B.n10 10.6151
R1173 B.n810 B.n809 10.6151
R1174 B.n811 B.n810 10.6151
R1175 B.n811 B.n8 10.6151
R1176 B.n815 B.n8 10.6151
R1177 B.n816 B.n815 10.6151
R1178 B.n817 B.n816 10.6151
R1179 B.n817 B.n6 10.6151
R1180 B.n821 B.n6 10.6151
R1181 B.n822 B.n821 10.6151
R1182 B.n823 B.n822 10.6151
R1183 B.n823 B.n4 10.6151
R1184 B.n827 B.n4 10.6151
R1185 B.n828 B.n827 10.6151
R1186 B.n829 B.n828 10.6151
R1187 B.n829 B.n0 10.6151
R1188 B.n709 B.n708 10.6151
R1189 B.n708 B.n707 10.6151
R1190 B.n707 B.n44 10.6151
R1191 B.n703 B.n44 10.6151
R1192 B.n703 B.n702 10.6151
R1193 B.n702 B.n701 10.6151
R1194 B.n701 B.n46 10.6151
R1195 B.n697 B.n46 10.6151
R1196 B.n697 B.n696 10.6151
R1197 B.n696 B.n695 10.6151
R1198 B.n695 B.n48 10.6151
R1199 B.n691 B.n48 10.6151
R1200 B.n691 B.n690 10.6151
R1201 B.n690 B.n689 10.6151
R1202 B.n689 B.n50 10.6151
R1203 B.n685 B.n684 10.6151
R1204 B.n684 B.n683 10.6151
R1205 B.n683 B.n55 10.6151
R1206 B.n679 B.n55 10.6151
R1207 B.n679 B.n678 10.6151
R1208 B.n678 B.n677 10.6151
R1209 B.n677 B.n57 10.6151
R1210 B.n673 B.n57 10.6151
R1211 B.n673 B.n672 10.6151
R1212 B.n670 B.n61 10.6151
R1213 B.n666 B.n61 10.6151
R1214 B.n666 B.n665 10.6151
R1215 B.n665 B.n664 10.6151
R1216 B.n664 B.n63 10.6151
R1217 B.n660 B.n63 10.6151
R1218 B.n660 B.n659 10.6151
R1219 B.n659 B.n658 10.6151
R1220 B.n658 B.n65 10.6151
R1221 B.n654 B.n65 10.6151
R1222 B.n654 B.n653 10.6151
R1223 B.n653 B.n652 10.6151
R1224 B.n652 B.n67 10.6151
R1225 B.n648 B.n67 10.6151
R1226 B.n648 B.n647 10.6151
R1227 B.n646 B.n69 10.6151
R1228 B.n642 B.n69 10.6151
R1229 B.n642 B.n641 10.6151
R1230 B.n641 B.n640 10.6151
R1231 B.n640 B.n71 10.6151
R1232 B.n636 B.n71 10.6151
R1233 B.n636 B.n635 10.6151
R1234 B.n635 B.n634 10.6151
R1235 B.n634 B.n73 10.6151
R1236 B.n630 B.n73 10.6151
R1237 B.n630 B.n629 10.6151
R1238 B.n629 B.n628 10.6151
R1239 B.n628 B.n75 10.6151
R1240 B.n624 B.n75 10.6151
R1241 B.n624 B.n623 10.6151
R1242 B.n623 B.n622 10.6151
R1243 B.n622 B.n77 10.6151
R1244 B.n618 B.n77 10.6151
R1245 B.n618 B.n617 10.6151
R1246 B.n617 B.n616 10.6151
R1247 B.n616 B.n79 10.6151
R1248 B.n612 B.n79 10.6151
R1249 B.n612 B.n611 10.6151
R1250 B.n611 B.n610 10.6151
R1251 B.n610 B.n81 10.6151
R1252 B.n606 B.n81 10.6151
R1253 B.n606 B.n605 10.6151
R1254 B.n605 B.n604 10.6151
R1255 B.n604 B.n83 10.6151
R1256 B.n600 B.n83 10.6151
R1257 B.n600 B.n599 10.6151
R1258 B.n599 B.n598 10.6151
R1259 B.n598 B.n85 10.6151
R1260 B.n594 B.n85 10.6151
R1261 B.n594 B.n593 10.6151
R1262 B.n593 B.n592 10.6151
R1263 B.n592 B.n87 10.6151
R1264 B.n588 B.n87 10.6151
R1265 B.n588 B.n587 10.6151
R1266 B.n587 B.n586 10.6151
R1267 B.n586 B.n89 10.6151
R1268 B.n582 B.n89 10.6151
R1269 B.n582 B.n581 10.6151
R1270 B.n581 B.n580 10.6151
R1271 B.n580 B.n91 10.6151
R1272 B.n576 B.n91 10.6151
R1273 B.n576 B.n575 10.6151
R1274 B.n575 B.n574 10.6151
R1275 B.n574 B.n93 10.6151
R1276 B.n570 B.n93 10.6151
R1277 B.n570 B.n569 10.6151
R1278 B.n569 B.n568 10.6151
R1279 B.n568 B.n95 10.6151
R1280 B.n564 B.n95 10.6151
R1281 B.n564 B.n563 10.6151
R1282 B.n563 B.n562 10.6151
R1283 B.n562 B.n97 10.6151
R1284 B.n558 B.n97 10.6151
R1285 B.n558 B.n557 10.6151
R1286 B.n557 B.n556 10.6151
R1287 B.n556 B.n99 10.6151
R1288 B.n552 B.n99 10.6151
R1289 B.n552 B.n551 10.6151
R1290 B.n551 B.n550 10.6151
R1291 B.n550 B.n101 10.6151
R1292 B.n546 B.n101 10.6151
R1293 B.n546 B.n545 10.6151
R1294 B.n545 B.n544 10.6151
R1295 B.n544 B.n103 10.6151
R1296 B.n540 B.n103 10.6151
R1297 B.n540 B.n539 10.6151
R1298 B.n539 B.n538 10.6151
R1299 B.n538 B.n105 10.6151
R1300 B.n534 B.n105 10.6151
R1301 B.n534 B.n533 10.6151
R1302 B.n533 B.n532 10.6151
R1303 B.n532 B.n107 10.6151
R1304 B.n528 B.n107 10.6151
R1305 B.n528 B.n527 10.6151
R1306 B.n527 B.n526 10.6151
R1307 B.n526 B.n109 10.6151
R1308 B.n522 B.n109 10.6151
R1309 B.n522 B.n521 10.6151
R1310 B.n521 B.n520 10.6151
R1311 B.n520 B.n111 10.6151
R1312 B.n516 B.n111 10.6151
R1313 B.n516 B.n515 10.6151
R1314 B.n515 B.n514 10.6151
R1315 B.n514 B.n113 10.6151
R1316 B.n510 B.n113 10.6151
R1317 B.n510 B.n509 10.6151
R1318 B.n509 B.n508 10.6151
R1319 B.n508 B.n115 10.6151
R1320 B.n504 B.n115 10.6151
R1321 B.n504 B.n503 10.6151
R1322 B.n503 B.n502 10.6151
R1323 B.n502 B.n117 10.6151
R1324 B.n498 B.n117 10.6151
R1325 B.n498 B.n497 10.6151
R1326 B.n497 B.n496 10.6151
R1327 B.n496 B.n119 10.6151
R1328 B.n492 B.n119 10.6151
R1329 B.n492 B.n491 10.6151
R1330 B.n491 B.n490 10.6151
R1331 B.n490 B.n121 10.6151
R1332 B.n486 B.n121 10.6151
R1333 B.n486 B.n485 10.6151
R1334 B.n485 B.n484 10.6151
R1335 B.n484 B.n123 10.6151
R1336 B.n480 B.n123 10.6151
R1337 B.n480 B.n479 10.6151
R1338 B.n479 B.n478 10.6151
R1339 B.n478 B.n125 10.6151
R1340 B.n474 B.n125 10.6151
R1341 B.n474 B.n473 10.6151
R1342 B.n473 B.n472 10.6151
R1343 B.n472 B.n127 10.6151
R1344 B.n468 B.n127 10.6151
R1345 B.n468 B.n467 10.6151
R1346 B.n467 B.n466 10.6151
R1347 B.n466 B.n129 10.6151
R1348 B.n462 B.n129 10.6151
R1349 B.n462 B.n461 10.6151
R1350 B.n461 B.n460 10.6151
R1351 B.n460 B.n131 10.6151
R1352 B.n456 B.n131 10.6151
R1353 B.n456 B.n455 10.6151
R1354 B.n455 B.n454 10.6151
R1355 B.n454 B.n133 10.6151
R1356 B.n450 B.n133 10.6151
R1357 B.n450 B.n449 10.6151
R1358 B.n449 B.n448 10.6151
R1359 B.n448 B.n135 10.6151
R1360 B.n444 B.n135 10.6151
R1361 B.n444 B.n443 10.6151
R1362 B.n443 B.n442 10.6151
R1363 B.n442 B.n137 10.6151
R1364 B.n438 B.n137 10.6151
R1365 B.n438 B.n437 10.6151
R1366 B.n437 B.n436 10.6151
R1367 B.n436 B.n139 10.6151
R1368 B.n432 B.n139 10.6151
R1369 B.n432 B.n431 10.6151
R1370 B.n431 B.n430 10.6151
R1371 B.n430 B.n141 10.6151
R1372 B.n426 B.n141 10.6151
R1373 B.n426 B.n425 10.6151
R1374 B.n425 B.n424 10.6151
R1375 B.n424 B.n143 10.6151
R1376 B.n420 B.n143 10.6151
R1377 B.n420 B.n419 10.6151
R1378 B.n419 B.n418 10.6151
R1379 B.n418 B.n145 10.6151
R1380 B.n414 B.n145 10.6151
R1381 B.n414 B.n413 10.6151
R1382 B.n413 B.n412 10.6151
R1383 B.n412 B.n147 10.6151
R1384 B.n408 B.n147 10.6151
R1385 B.n408 B.n407 10.6151
R1386 B.n407 B.n406 10.6151
R1387 B.n406 B.n149 10.6151
R1388 B.n402 B.n149 10.6151
R1389 B.n402 B.n401 10.6151
R1390 B.n213 B.n1 10.6151
R1391 B.n216 B.n213 10.6151
R1392 B.n217 B.n216 10.6151
R1393 B.n218 B.n217 10.6151
R1394 B.n218 B.n211 10.6151
R1395 B.n222 B.n211 10.6151
R1396 B.n223 B.n222 10.6151
R1397 B.n224 B.n223 10.6151
R1398 B.n224 B.n209 10.6151
R1399 B.n228 B.n209 10.6151
R1400 B.n229 B.n228 10.6151
R1401 B.n230 B.n229 10.6151
R1402 B.n230 B.n207 10.6151
R1403 B.n234 B.n207 10.6151
R1404 B.n235 B.n234 10.6151
R1405 B.n236 B.n235 10.6151
R1406 B.n236 B.n205 10.6151
R1407 B.n240 B.n205 10.6151
R1408 B.n241 B.n240 10.6151
R1409 B.n242 B.n241 10.6151
R1410 B.n242 B.n203 10.6151
R1411 B.n246 B.n203 10.6151
R1412 B.n247 B.n246 10.6151
R1413 B.n248 B.n247 10.6151
R1414 B.n248 B.n201 10.6151
R1415 B.n252 B.n201 10.6151
R1416 B.n253 B.n252 10.6151
R1417 B.n254 B.n253 10.6151
R1418 B.n254 B.n199 10.6151
R1419 B.n258 B.n199 10.6151
R1420 B.n259 B.n258 10.6151
R1421 B.n260 B.n259 10.6151
R1422 B.n260 B.n197 10.6151
R1423 B.n264 B.n197 10.6151
R1424 B.n265 B.n264 10.6151
R1425 B.n266 B.n265 10.6151
R1426 B.n266 B.n195 10.6151
R1427 B.n270 B.n195 10.6151
R1428 B.n271 B.n270 10.6151
R1429 B.n272 B.n271 10.6151
R1430 B.n272 B.n193 10.6151
R1431 B.n276 B.n193 10.6151
R1432 B.n277 B.n276 10.6151
R1433 B.n278 B.n277 10.6151
R1434 B.n278 B.n191 10.6151
R1435 B.n282 B.n191 10.6151
R1436 B.n283 B.n282 10.6151
R1437 B.n284 B.n283 10.6151
R1438 B.n284 B.n189 10.6151
R1439 B.n288 B.n189 10.6151
R1440 B.n289 B.n288 10.6151
R1441 B.n290 B.n289 10.6151
R1442 B.n290 B.n187 10.6151
R1443 B.n294 B.n187 10.6151
R1444 B.n295 B.n294 10.6151
R1445 B.n296 B.n295 10.6151
R1446 B.n296 B.n185 10.6151
R1447 B.n300 B.n185 10.6151
R1448 B.n301 B.n300 10.6151
R1449 B.n302 B.n301 10.6151
R1450 B.n302 B.n183 10.6151
R1451 B.n306 B.n183 10.6151
R1452 B.n307 B.n306 10.6151
R1453 B.n308 B.n307 10.6151
R1454 B.n308 B.n181 10.6151
R1455 B.n312 B.n181 10.6151
R1456 B.n313 B.n312 10.6151
R1457 B.n314 B.n313 10.6151
R1458 B.n314 B.n179 10.6151
R1459 B.n318 B.n179 10.6151
R1460 B.n319 B.n318 10.6151
R1461 B.n320 B.n319 10.6151
R1462 B.n320 B.n177 10.6151
R1463 B.n324 B.n177 10.6151
R1464 B.n325 B.n324 10.6151
R1465 B.n326 B.n325 10.6151
R1466 B.n326 B.n175 10.6151
R1467 B.n330 B.n175 10.6151
R1468 B.n331 B.n330 10.6151
R1469 B.n332 B.n331 10.6151
R1470 B.n336 B.n173 10.6151
R1471 B.n337 B.n336 10.6151
R1472 B.n338 B.n337 10.6151
R1473 B.n338 B.n171 10.6151
R1474 B.n342 B.n171 10.6151
R1475 B.n343 B.n342 10.6151
R1476 B.n344 B.n343 10.6151
R1477 B.n344 B.n169 10.6151
R1478 B.n348 B.n169 10.6151
R1479 B.n349 B.n348 10.6151
R1480 B.n350 B.n349 10.6151
R1481 B.n350 B.n167 10.6151
R1482 B.n354 B.n167 10.6151
R1483 B.n355 B.n354 10.6151
R1484 B.n359 B.n355 10.6151
R1485 B.n363 B.n165 10.6151
R1486 B.n364 B.n363 10.6151
R1487 B.n365 B.n364 10.6151
R1488 B.n365 B.n163 10.6151
R1489 B.n369 B.n163 10.6151
R1490 B.n370 B.n369 10.6151
R1491 B.n371 B.n370 10.6151
R1492 B.n371 B.n161 10.6151
R1493 B.n375 B.n161 10.6151
R1494 B.n378 B.n377 10.6151
R1495 B.n378 B.n157 10.6151
R1496 B.n382 B.n157 10.6151
R1497 B.n383 B.n382 10.6151
R1498 B.n384 B.n383 10.6151
R1499 B.n384 B.n155 10.6151
R1500 B.n388 B.n155 10.6151
R1501 B.n389 B.n388 10.6151
R1502 B.n390 B.n389 10.6151
R1503 B.n390 B.n153 10.6151
R1504 B.n394 B.n153 10.6151
R1505 B.n395 B.n394 10.6151
R1506 B.n396 B.n395 10.6151
R1507 B.n396 B.n151 10.6151
R1508 B.n400 B.n151 10.6151
R1509 B.n54 B.n50 9.36635
R1510 B.n671 B.n670 9.36635
R1511 B.n359 B.n358 9.36635
R1512 B.n377 B.n376 9.36635
R1513 B.n833 B.n0 8.11757
R1514 B.n833 B.n1 8.11757
R1515 B.n685 B.n54 1.24928
R1516 B.n672 B.n671 1.24928
R1517 B.n358 B.n165 1.24928
R1518 B.n376 B.n375 1.24928
R1519 VN.n110 VN.n109 161.3
R1520 VN.n108 VN.n57 161.3
R1521 VN.n107 VN.n106 161.3
R1522 VN.n105 VN.n58 161.3
R1523 VN.n104 VN.n103 161.3
R1524 VN.n102 VN.n59 161.3
R1525 VN.n101 VN.n100 161.3
R1526 VN.n99 VN.n60 161.3
R1527 VN.n98 VN.n97 161.3
R1528 VN.n95 VN.n61 161.3
R1529 VN.n94 VN.n93 161.3
R1530 VN.n92 VN.n62 161.3
R1531 VN.n91 VN.n90 161.3
R1532 VN.n89 VN.n63 161.3
R1533 VN.n88 VN.n87 161.3
R1534 VN.n86 VN.n64 161.3
R1535 VN.n85 VN.n84 161.3
R1536 VN.n82 VN.n65 161.3
R1537 VN.n81 VN.n80 161.3
R1538 VN.n79 VN.n66 161.3
R1539 VN.n78 VN.n77 161.3
R1540 VN.n76 VN.n67 161.3
R1541 VN.n75 VN.n74 161.3
R1542 VN.n73 VN.n68 161.3
R1543 VN.n72 VN.n71 161.3
R1544 VN.n54 VN.n53 161.3
R1545 VN.n52 VN.n1 161.3
R1546 VN.n51 VN.n50 161.3
R1547 VN.n49 VN.n2 161.3
R1548 VN.n48 VN.n47 161.3
R1549 VN.n46 VN.n3 161.3
R1550 VN.n45 VN.n44 161.3
R1551 VN.n43 VN.n4 161.3
R1552 VN.n42 VN.n41 161.3
R1553 VN.n39 VN.n5 161.3
R1554 VN.n38 VN.n37 161.3
R1555 VN.n36 VN.n6 161.3
R1556 VN.n35 VN.n34 161.3
R1557 VN.n33 VN.n7 161.3
R1558 VN.n32 VN.n31 161.3
R1559 VN.n30 VN.n8 161.3
R1560 VN.n29 VN.n28 161.3
R1561 VN.n26 VN.n9 161.3
R1562 VN.n25 VN.n24 161.3
R1563 VN.n23 VN.n10 161.3
R1564 VN.n22 VN.n21 161.3
R1565 VN.n20 VN.n11 161.3
R1566 VN.n19 VN.n18 161.3
R1567 VN.n17 VN.n12 161.3
R1568 VN.n16 VN.n15 161.3
R1569 VN.n55 VN.n0 87.6207
R1570 VN.n111 VN.n56 87.6207
R1571 VN.n21 VN.n20 56.5193
R1572 VN.n34 VN.n33 56.5193
R1573 VN.n77 VN.n76 56.5193
R1574 VN.n90 VN.n89 56.5193
R1575 VN.n14 VN.n13 55.4712
R1576 VN.n70 VN.n69 55.4712
R1577 VN.n69 VN.t3 54.2693
R1578 VN.n13 VN.t6 54.2693
R1579 VN VN.n111 53.4564
R1580 VN.n47 VN.n46 42.9216
R1581 VN.n103 VN.n102 42.9216
R1582 VN.n47 VN.n2 38.0652
R1583 VN.n103 VN.n58 38.0652
R1584 VN.n15 VN.n12 24.4675
R1585 VN.n19 VN.n12 24.4675
R1586 VN.n20 VN.n19 24.4675
R1587 VN.n21 VN.n10 24.4675
R1588 VN.n25 VN.n10 24.4675
R1589 VN.n26 VN.n25 24.4675
R1590 VN.n28 VN.n8 24.4675
R1591 VN.n32 VN.n8 24.4675
R1592 VN.n33 VN.n32 24.4675
R1593 VN.n34 VN.n6 24.4675
R1594 VN.n38 VN.n6 24.4675
R1595 VN.n39 VN.n38 24.4675
R1596 VN.n41 VN.n4 24.4675
R1597 VN.n45 VN.n4 24.4675
R1598 VN.n46 VN.n45 24.4675
R1599 VN.n51 VN.n2 24.4675
R1600 VN.n52 VN.n51 24.4675
R1601 VN.n53 VN.n52 24.4675
R1602 VN.n76 VN.n75 24.4675
R1603 VN.n75 VN.n68 24.4675
R1604 VN.n71 VN.n68 24.4675
R1605 VN.n89 VN.n88 24.4675
R1606 VN.n88 VN.n64 24.4675
R1607 VN.n84 VN.n64 24.4675
R1608 VN.n82 VN.n81 24.4675
R1609 VN.n81 VN.n66 24.4675
R1610 VN.n77 VN.n66 24.4675
R1611 VN.n102 VN.n101 24.4675
R1612 VN.n101 VN.n60 24.4675
R1613 VN.n97 VN.n60 24.4675
R1614 VN.n95 VN.n94 24.4675
R1615 VN.n94 VN.n62 24.4675
R1616 VN.n90 VN.n62 24.4675
R1617 VN.n109 VN.n108 24.4675
R1618 VN.n108 VN.n107 24.4675
R1619 VN.n107 VN.n58 24.4675
R1620 VN.n14 VN.t0 21.5139
R1621 VN.n27 VN.t5 21.5139
R1622 VN.n40 VN.t9 21.5139
R1623 VN.n0 VN.t8 21.5139
R1624 VN.n70 VN.t2 21.5139
R1625 VN.n83 VN.t4 21.5139
R1626 VN.n96 VN.t1 21.5139
R1627 VN.n56 VN.t7 21.5139
R1628 VN.n15 VN.n14 19.5741
R1629 VN.n40 VN.n39 19.5741
R1630 VN.n71 VN.n70 19.5741
R1631 VN.n96 VN.n95 19.5741
R1632 VN.n27 VN.n26 12.234
R1633 VN.n28 VN.n27 12.234
R1634 VN.n84 VN.n83 12.234
R1635 VN.n83 VN.n82 12.234
R1636 VN.n41 VN.n40 4.8939
R1637 VN.n97 VN.n96 4.8939
R1638 VN.n72 VN.n69 2.47314
R1639 VN.n16 VN.n13 2.47314
R1640 VN.n53 VN.n0 2.4472
R1641 VN.n109 VN.n56 2.4472
R1642 VN.n111 VN.n110 0.354971
R1643 VN.n55 VN.n54 0.354971
R1644 VN VN.n55 0.26696
R1645 VN.n110 VN.n57 0.189894
R1646 VN.n106 VN.n57 0.189894
R1647 VN.n106 VN.n105 0.189894
R1648 VN.n105 VN.n104 0.189894
R1649 VN.n104 VN.n59 0.189894
R1650 VN.n100 VN.n59 0.189894
R1651 VN.n100 VN.n99 0.189894
R1652 VN.n99 VN.n98 0.189894
R1653 VN.n98 VN.n61 0.189894
R1654 VN.n93 VN.n61 0.189894
R1655 VN.n93 VN.n92 0.189894
R1656 VN.n92 VN.n91 0.189894
R1657 VN.n91 VN.n63 0.189894
R1658 VN.n87 VN.n63 0.189894
R1659 VN.n87 VN.n86 0.189894
R1660 VN.n86 VN.n85 0.189894
R1661 VN.n85 VN.n65 0.189894
R1662 VN.n80 VN.n65 0.189894
R1663 VN.n80 VN.n79 0.189894
R1664 VN.n79 VN.n78 0.189894
R1665 VN.n78 VN.n67 0.189894
R1666 VN.n74 VN.n67 0.189894
R1667 VN.n74 VN.n73 0.189894
R1668 VN.n73 VN.n72 0.189894
R1669 VN.n17 VN.n16 0.189894
R1670 VN.n18 VN.n17 0.189894
R1671 VN.n18 VN.n11 0.189894
R1672 VN.n22 VN.n11 0.189894
R1673 VN.n23 VN.n22 0.189894
R1674 VN.n24 VN.n23 0.189894
R1675 VN.n24 VN.n9 0.189894
R1676 VN.n29 VN.n9 0.189894
R1677 VN.n30 VN.n29 0.189894
R1678 VN.n31 VN.n30 0.189894
R1679 VN.n31 VN.n7 0.189894
R1680 VN.n35 VN.n7 0.189894
R1681 VN.n36 VN.n35 0.189894
R1682 VN.n37 VN.n36 0.189894
R1683 VN.n37 VN.n5 0.189894
R1684 VN.n42 VN.n5 0.189894
R1685 VN.n43 VN.n42 0.189894
R1686 VN.n44 VN.n43 0.189894
R1687 VN.n44 VN.n3 0.189894
R1688 VN.n48 VN.n3 0.189894
R1689 VN.n49 VN.n48 0.189894
R1690 VN.n50 VN.n49 0.189894
R1691 VN.n50 VN.n1 0.189894
R1692 VN.n54 VN.n1 0.189894
R1693 VDD2.n1 VDD2.t3 131.661
R1694 VDD2.n4 VDD2.t2 128.083
R1695 VDD2.n3 VDD2.n2 121.178
R1696 VDD2 VDD2.n7 121.175
R1697 VDD2.n6 VDD2.n5 118.55
R1698 VDD2.n1 VDD2.n0 118.55
R1699 VDD2.n4 VDD2.n3 43.6485
R1700 VDD2.n7 VDD2.t7 9.53276
R1701 VDD2.n7 VDD2.t6 9.53276
R1702 VDD2.n5 VDD2.t8 9.53276
R1703 VDD2.n5 VDD2.t5 9.53276
R1704 VDD2.n2 VDD2.t0 9.53276
R1705 VDD2.n2 VDD2.t1 9.53276
R1706 VDD2.n0 VDD2.t9 9.53276
R1707 VDD2.n0 VDD2.t4 9.53276
R1708 VDD2.n6 VDD2.n4 3.57809
R1709 VDD2 VDD2.n6 0.953086
R1710 VDD2.n3 VDD2.n1 0.839551
C0 VN VTAIL 5.57025f
C1 VN w_n5950_n1650# 12.973701f
C2 VP VTAIL 5.58454f
C3 VP w_n5950_n1650# 13.7505f
C4 VTAIL w_n5950_n1650# 2.20571f
C5 B VDD1 2.25904f
C6 VDD1 VDD2 2.96809f
C7 B VDD2 2.42473f
C8 VN VDD1 0.160861f
C9 VP VDD1 4.21442f
C10 VN B 1.53912f
C11 VP B 2.85449f
C12 VTAIL VDD1 7.70595f
C13 VDD1 w_n5950_n1650# 2.66084f
C14 VN VDD2 3.63506f
C15 VP VDD2 0.744317f
C16 B VTAIL 2.06616f
C17 B w_n5950_n1650# 10.2416f
C18 VTAIL VDD2 7.76737f
C19 VDD2 w_n5950_n1650# 2.86736f
C20 VN VP 8.61357f
C21 VDD2 VSUBS 2.592382f
C22 VDD1 VSUBS 2.312575f
C23 VTAIL VSUBS 0.777844f
C24 VN VSUBS 9.703111f
C25 VP VSUBS 5.063719f
C26 B VSUBS 5.764848f
C27 w_n5950_n1650# VSUBS 0.124022p
C28 VDD2.t3 VSUBS 0.851644f
C29 VDD2.t9 VSUBS 0.106601f
C30 VDD2.t4 VSUBS 0.106601f
C31 VDD2.n0 VSUBS 0.589857f
C32 VDD2.n1 VSUBS 2.11526f
C33 VDD2.t0 VSUBS 0.106601f
C34 VDD2.t1 VSUBS 0.106601f
C35 VDD2.n2 VSUBS 0.618751f
C36 VDD2.n3 VSUBS 4.985f
C37 VDD2.t2 VSUBS 0.822988f
C38 VDD2.n4 VSUBS 4.79363f
C39 VDD2.t8 VSUBS 0.106601f
C40 VDD2.t5 VSUBS 0.106601f
C41 VDD2.n5 VSUBS 0.589859f
C42 VDD2.n6 VSUBS 1.10259f
C43 VDD2.t7 VSUBS 0.106601f
C44 VDD2.t6 VSUBS 0.106601f
C45 VDD2.n7 VSUBS 0.618705f
C46 VN.t8 VSUBS 1.27529f
C47 VN.n0 VSUBS 0.651937f
C48 VN.n1 VSUBS 0.038719f
C49 VN.n2 VSUBS 0.077762f
C50 VN.n3 VSUBS 0.038719f
C51 VN.n4 VSUBS 0.072163f
C52 VN.n5 VSUBS 0.038719f
C53 VN.t9 VSUBS 1.27529f
C54 VN.n6 VSUBS 0.072163f
C55 VN.n7 VSUBS 0.038719f
C56 VN.n8 VSUBS 0.072163f
C57 VN.n9 VSUBS 0.038719f
C58 VN.t5 VSUBS 1.27529f
C59 VN.n10 VSUBS 0.072163f
C60 VN.n11 VSUBS 0.038719f
C61 VN.n12 VSUBS 0.072163f
C62 VN.t6 VSUBS 1.76798f
C63 VN.n13 VSUBS 0.678096f
C64 VN.t0 VSUBS 1.27529f
C65 VN.n14 VSUBS 0.657571f
C66 VN.n15 VSUBS 0.065037f
C67 VN.n16 VSUBS 0.499054f
C68 VN.n17 VSUBS 0.038719f
C69 VN.n18 VSUBS 0.038719f
C70 VN.n19 VSUBS 0.072163f
C71 VN.n20 VSUBS 0.048435f
C72 VN.n21 VSUBS 0.064618f
C73 VN.n22 VSUBS 0.038719f
C74 VN.n23 VSUBS 0.038719f
C75 VN.n24 VSUBS 0.038719f
C76 VN.n25 VSUBS 0.072163f
C77 VN.n26 VSUBS 0.054349f
C78 VN.n27 VSUBS 0.506781f
C79 VN.n28 VSUBS 0.054349f
C80 VN.n29 VSUBS 0.038719f
C81 VN.n30 VSUBS 0.038719f
C82 VN.n31 VSUBS 0.038719f
C83 VN.n32 VSUBS 0.072163f
C84 VN.n33 VSUBS 0.064618f
C85 VN.n34 VSUBS 0.048435f
C86 VN.n35 VSUBS 0.038719f
C87 VN.n36 VSUBS 0.038719f
C88 VN.n37 VSUBS 0.038719f
C89 VN.n38 VSUBS 0.072163f
C90 VN.n39 VSUBS 0.065037f
C91 VN.n40 VSUBS 0.506781f
C92 VN.n41 VSUBS 0.043661f
C93 VN.n42 VSUBS 0.038719f
C94 VN.n43 VSUBS 0.038719f
C95 VN.n44 VSUBS 0.038719f
C96 VN.n45 VSUBS 0.072163f
C97 VN.n46 VSUBS 0.075839f
C98 VN.n47 VSUBS 0.031614f
C99 VN.n48 VSUBS 0.038719f
C100 VN.n49 VSUBS 0.038719f
C101 VN.n50 VSUBS 0.038719f
C102 VN.n51 VSUBS 0.072163f
C103 VN.n52 VSUBS 0.072163f
C104 VN.n53 VSUBS 0.040098f
C105 VN.n54 VSUBS 0.062492f
C106 VN.n55 VSUBS 0.119879f
C107 VN.t7 VSUBS 1.27529f
C108 VN.n56 VSUBS 0.651937f
C109 VN.n57 VSUBS 0.038719f
C110 VN.n58 VSUBS 0.077762f
C111 VN.n59 VSUBS 0.038719f
C112 VN.n60 VSUBS 0.072163f
C113 VN.n61 VSUBS 0.038719f
C114 VN.t1 VSUBS 1.27529f
C115 VN.n62 VSUBS 0.072163f
C116 VN.n63 VSUBS 0.038719f
C117 VN.n64 VSUBS 0.072163f
C118 VN.n65 VSUBS 0.038719f
C119 VN.t4 VSUBS 1.27529f
C120 VN.n66 VSUBS 0.072163f
C121 VN.n67 VSUBS 0.038719f
C122 VN.n68 VSUBS 0.072163f
C123 VN.t3 VSUBS 1.76798f
C124 VN.n69 VSUBS 0.678096f
C125 VN.t2 VSUBS 1.27529f
C126 VN.n70 VSUBS 0.657571f
C127 VN.n71 VSUBS 0.065037f
C128 VN.n72 VSUBS 0.499054f
C129 VN.n73 VSUBS 0.038719f
C130 VN.n74 VSUBS 0.038719f
C131 VN.n75 VSUBS 0.072163f
C132 VN.n76 VSUBS 0.048435f
C133 VN.n77 VSUBS 0.064618f
C134 VN.n78 VSUBS 0.038719f
C135 VN.n79 VSUBS 0.038719f
C136 VN.n80 VSUBS 0.038719f
C137 VN.n81 VSUBS 0.072163f
C138 VN.n82 VSUBS 0.054349f
C139 VN.n83 VSUBS 0.506781f
C140 VN.n84 VSUBS 0.054349f
C141 VN.n85 VSUBS 0.038719f
C142 VN.n86 VSUBS 0.038719f
C143 VN.n87 VSUBS 0.038719f
C144 VN.n88 VSUBS 0.072163f
C145 VN.n89 VSUBS 0.064618f
C146 VN.n90 VSUBS 0.048435f
C147 VN.n91 VSUBS 0.038719f
C148 VN.n92 VSUBS 0.038719f
C149 VN.n93 VSUBS 0.038719f
C150 VN.n94 VSUBS 0.072163f
C151 VN.n95 VSUBS 0.065037f
C152 VN.n96 VSUBS 0.506781f
C153 VN.n97 VSUBS 0.043661f
C154 VN.n98 VSUBS 0.038719f
C155 VN.n99 VSUBS 0.038719f
C156 VN.n100 VSUBS 0.038719f
C157 VN.n101 VSUBS 0.072163f
C158 VN.n102 VSUBS 0.075839f
C159 VN.n103 VSUBS 0.031614f
C160 VN.n104 VSUBS 0.038719f
C161 VN.n105 VSUBS 0.038719f
C162 VN.n106 VSUBS 0.038719f
C163 VN.n107 VSUBS 0.072163f
C164 VN.n108 VSUBS 0.072163f
C165 VN.n109 VSUBS 0.040098f
C166 VN.n110 VSUBS 0.062492f
C167 VN.n111 VSUBS 2.45302f
C168 B.n0 VSUBS 0.012323f
C169 B.n1 VSUBS 0.012323f
C170 B.n2 VSUBS 0.018225f
C171 B.n3 VSUBS 0.013966f
C172 B.n4 VSUBS 0.013966f
C173 B.n5 VSUBS 0.013966f
C174 B.n6 VSUBS 0.013966f
C175 B.n7 VSUBS 0.013966f
C176 B.n8 VSUBS 0.013966f
C177 B.n9 VSUBS 0.013966f
C178 B.n10 VSUBS 0.013966f
C179 B.n11 VSUBS 0.013966f
C180 B.n12 VSUBS 0.013966f
C181 B.n13 VSUBS 0.013966f
C182 B.n14 VSUBS 0.013966f
C183 B.n15 VSUBS 0.013966f
C184 B.n16 VSUBS 0.013966f
C185 B.n17 VSUBS 0.013966f
C186 B.n18 VSUBS 0.013966f
C187 B.n19 VSUBS 0.013966f
C188 B.n20 VSUBS 0.013966f
C189 B.n21 VSUBS 0.013966f
C190 B.n22 VSUBS 0.013966f
C191 B.n23 VSUBS 0.013966f
C192 B.n24 VSUBS 0.013966f
C193 B.n25 VSUBS 0.013966f
C194 B.n26 VSUBS 0.013966f
C195 B.n27 VSUBS 0.013966f
C196 B.n28 VSUBS 0.013966f
C197 B.n29 VSUBS 0.013966f
C198 B.n30 VSUBS 0.013966f
C199 B.n31 VSUBS 0.013966f
C200 B.n32 VSUBS 0.013966f
C201 B.n33 VSUBS 0.013966f
C202 B.n34 VSUBS 0.013966f
C203 B.n35 VSUBS 0.013966f
C204 B.n36 VSUBS 0.013966f
C205 B.n37 VSUBS 0.013966f
C206 B.n38 VSUBS 0.013966f
C207 B.n39 VSUBS 0.013966f
C208 B.n40 VSUBS 0.013966f
C209 B.n41 VSUBS 0.013966f
C210 B.n42 VSUBS 0.032064f
C211 B.n43 VSUBS 0.013966f
C212 B.n44 VSUBS 0.013966f
C213 B.n45 VSUBS 0.013966f
C214 B.n46 VSUBS 0.013966f
C215 B.n47 VSUBS 0.013966f
C216 B.n48 VSUBS 0.013966f
C217 B.n49 VSUBS 0.013966f
C218 B.n50 VSUBS 0.013144f
C219 B.n51 VSUBS 0.013966f
C220 B.t10 VSUBS 0.17092f
C221 B.t11 VSUBS 0.218711f
C222 B.t9 VSUBS 1.2712f
C223 B.n52 VSUBS 0.188634f
C224 B.n53 VSUBS 0.142996f
C225 B.n54 VSUBS 0.032357f
C226 B.n55 VSUBS 0.013966f
C227 B.n56 VSUBS 0.013966f
C228 B.n57 VSUBS 0.013966f
C229 B.n58 VSUBS 0.013966f
C230 B.t1 VSUBS 0.170921f
C231 B.t2 VSUBS 0.21871f
C232 B.t0 VSUBS 1.2712f
C233 B.n59 VSUBS 0.188635f
C234 B.n60 VSUBS 0.142995f
C235 B.n61 VSUBS 0.013966f
C236 B.n62 VSUBS 0.013966f
C237 B.n63 VSUBS 0.013966f
C238 B.n64 VSUBS 0.013966f
C239 B.n65 VSUBS 0.013966f
C240 B.n66 VSUBS 0.013966f
C241 B.n67 VSUBS 0.013966f
C242 B.n68 VSUBS 0.032837f
C243 B.n69 VSUBS 0.013966f
C244 B.n70 VSUBS 0.013966f
C245 B.n71 VSUBS 0.013966f
C246 B.n72 VSUBS 0.013966f
C247 B.n73 VSUBS 0.013966f
C248 B.n74 VSUBS 0.013966f
C249 B.n75 VSUBS 0.013966f
C250 B.n76 VSUBS 0.013966f
C251 B.n77 VSUBS 0.013966f
C252 B.n78 VSUBS 0.013966f
C253 B.n79 VSUBS 0.013966f
C254 B.n80 VSUBS 0.013966f
C255 B.n81 VSUBS 0.013966f
C256 B.n82 VSUBS 0.013966f
C257 B.n83 VSUBS 0.013966f
C258 B.n84 VSUBS 0.013966f
C259 B.n85 VSUBS 0.013966f
C260 B.n86 VSUBS 0.013966f
C261 B.n87 VSUBS 0.013966f
C262 B.n88 VSUBS 0.013966f
C263 B.n89 VSUBS 0.013966f
C264 B.n90 VSUBS 0.013966f
C265 B.n91 VSUBS 0.013966f
C266 B.n92 VSUBS 0.013966f
C267 B.n93 VSUBS 0.013966f
C268 B.n94 VSUBS 0.013966f
C269 B.n95 VSUBS 0.013966f
C270 B.n96 VSUBS 0.013966f
C271 B.n97 VSUBS 0.013966f
C272 B.n98 VSUBS 0.013966f
C273 B.n99 VSUBS 0.013966f
C274 B.n100 VSUBS 0.013966f
C275 B.n101 VSUBS 0.013966f
C276 B.n102 VSUBS 0.013966f
C277 B.n103 VSUBS 0.013966f
C278 B.n104 VSUBS 0.013966f
C279 B.n105 VSUBS 0.013966f
C280 B.n106 VSUBS 0.013966f
C281 B.n107 VSUBS 0.013966f
C282 B.n108 VSUBS 0.013966f
C283 B.n109 VSUBS 0.013966f
C284 B.n110 VSUBS 0.013966f
C285 B.n111 VSUBS 0.013966f
C286 B.n112 VSUBS 0.013966f
C287 B.n113 VSUBS 0.013966f
C288 B.n114 VSUBS 0.013966f
C289 B.n115 VSUBS 0.013966f
C290 B.n116 VSUBS 0.013966f
C291 B.n117 VSUBS 0.013966f
C292 B.n118 VSUBS 0.013966f
C293 B.n119 VSUBS 0.013966f
C294 B.n120 VSUBS 0.013966f
C295 B.n121 VSUBS 0.013966f
C296 B.n122 VSUBS 0.013966f
C297 B.n123 VSUBS 0.013966f
C298 B.n124 VSUBS 0.013966f
C299 B.n125 VSUBS 0.013966f
C300 B.n126 VSUBS 0.013966f
C301 B.n127 VSUBS 0.013966f
C302 B.n128 VSUBS 0.013966f
C303 B.n129 VSUBS 0.013966f
C304 B.n130 VSUBS 0.013966f
C305 B.n131 VSUBS 0.013966f
C306 B.n132 VSUBS 0.013966f
C307 B.n133 VSUBS 0.013966f
C308 B.n134 VSUBS 0.013966f
C309 B.n135 VSUBS 0.013966f
C310 B.n136 VSUBS 0.013966f
C311 B.n137 VSUBS 0.013966f
C312 B.n138 VSUBS 0.013966f
C313 B.n139 VSUBS 0.013966f
C314 B.n140 VSUBS 0.013966f
C315 B.n141 VSUBS 0.013966f
C316 B.n142 VSUBS 0.013966f
C317 B.n143 VSUBS 0.013966f
C318 B.n144 VSUBS 0.013966f
C319 B.n145 VSUBS 0.013966f
C320 B.n146 VSUBS 0.013966f
C321 B.n147 VSUBS 0.013966f
C322 B.n148 VSUBS 0.013966f
C323 B.n149 VSUBS 0.013966f
C324 B.n150 VSUBS 0.032064f
C325 B.n151 VSUBS 0.013966f
C326 B.n152 VSUBS 0.013966f
C327 B.n153 VSUBS 0.013966f
C328 B.n154 VSUBS 0.013966f
C329 B.n155 VSUBS 0.013966f
C330 B.n156 VSUBS 0.013966f
C331 B.n157 VSUBS 0.013966f
C332 B.n158 VSUBS 0.013966f
C333 B.t8 VSUBS 0.170921f
C334 B.t7 VSUBS 0.21871f
C335 B.t6 VSUBS 1.2712f
C336 B.n159 VSUBS 0.188635f
C337 B.n160 VSUBS 0.142995f
C338 B.n161 VSUBS 0.013966f
C339 B.n162 VSUBS 0.013966f
C340 B.n163 VSUBS 0.013966f
C341 B.n164 VSUBS 0.013966f
C342 B.n165 VSUBS 0.007804f
C343 B.n166 VSUBS 0.013966f
C344 B.n167 VSUBS 0.013966f
C345 B.n168 VSUBS 0.013966f
C346 B.n169 VSUBS 0.013966f
C347 B.n170 VSUBS 0.013966f
C348 B.n171 VSUBS 0.013966f
C349 B.n172 VSUBS 0.013966f
C350 B.n173 VSUBS 0.032837f
C351 B.n174 VSUBS 0.013966f
C352 B.n175 VSUBS 0.013966f
C353 B.n176 VSUBS 0.013966f
C354 B.n177 VSUBS 0.013966f
C355 B.n178 VSUBS 0.013966f
C356 B.n179 VSUBS 0.013966f
C357 B.n180 VSUBS 0.013966f
C358 B.n181 VSUBS 0.013966f
C359 B.n182 VSUBS 0.013966f
C360 B.n183 VSUBS 0.013966f
C361 B.n184 VSUBS 0.013966f
C362 B.n185 VSUBS 0.013966f
C363 B.n186 VSUBS 0.013966f
C364 B.n187 VSUBS 0.013966f
C365 B.n188 VSUBS 0.013966f
C366 B.n189 VSUBS 0.013966f
C367 B.n190 VSUBS 0.013966f
C368 B.n191 VSUBS 0.013966f
C369 B.n192 VSUBS 0.013966f
C370 B.n193 VSUBS 0.013966f
C371 B.n194 VSUBS 0.013966f
C372 B.n195 VSUBS 0.013966f
C373 B.n196 VSUBS 0.013966f
C374 B.n197 VSUBS 0.013966f
C375 B.n198 VSUBS 0.013966f
C376 B.n199 VSUBS 0.013966f
C377 B.n200 VSUBS 0.013966f
C378 B.n201 VSUBS 0.013966f
C379 B.n202 VSUBS 0.013966f
C380 B.n203 VSUBS 0.013966f
C381 B.n204 VSUBS 0.013966f
C382 B.n205 VSUBS 0.013966f
C383 B.n206 VSUBS 0.013966f
C384 B.n207 VSUBS 0.013966f
C385 B.n208 VSUBS 0.013966f
C386 B.n209 VSUBS 0.013966f
C387 B.n210 VSUBS 0.013966f
C388 B.n211 VSUBS 0.013966f
C389 B.n212 VSUBS 0.013966f
C390 B.n213 VSUBS 0.013966f
C391 B.n214 VSUBS 0.013966f
C392 B.n215 VSUBS 0.013966f
C393 B.n216 VSUBS 0.013966f
C394 B.n217 VSUBS 0.013966f
C395 B.n218 VSUBS 0.013966f
C396 B.n219 VSUBS 0.013966f
C397 B.n220 VSUBS 0.013966f
C398 B.n221 VSUBS 0.013966f
C399 B.n222 VSUBS 0.013966f
C400 B.n223 VSUBS 0.013966f
C401 B.n224 VSUBS 0.013966f
C402 B.n225 VSUBS 0.013966f
C403 B.n226 VSUBS 0.013966f
C404 B.n227 VSUBS 0.013966f
C405 B.n228 VSUBS 0.013966f
C406 B.n229 VSUBS 0.013966f
C407 B.n230 VSUBS 0.013966f
C408 B.n231 VSUBS 0.013966f
C409 B.n232 VSUBS 0.013966f
C410 B.n233 VSUBS 0.013966f
C411 B.n234 VSUBS 0.013966f
C412 B.n235 VSUBS 0.013966f
C413 B.n236 VSUBS 0.013966f
C414 B.n237 VSUBS 0.013966f
C415 B.n238 VSUBS 0.013966f
C416 B.n239 VSUBS 0.013966f
C417 B.n240 VSUBS 0.013966f
C418 B.n241 VSUBS 0.013966f
C419 B.n242 VSUBS 0.013966f
C420 B.n243 VSUBS 0.013966f
C421 B.n244 VSUBS 0.013966f
C422 B.n245 VSUBS 0.013966f
C423 B.n246 VSUBS 0.013966f
C424 B.n247 VSUBS 0.013966f
C425 B.n248 VSUBS 0.013966f
C426 B.n249 VSUBS 0.013966f
C427 B.n250 VSUBS 0.013966f
C428 B.n251 VSUBS 0.013966f
C429 B.n252 VSUBS 0.013966f
C430 B.n253 VSUBS 0.013966f
C431 B.n254 VSUBS 0.013966f
C432 B.n255 VSUBS 0.013966f
C433 B.n256 VSUBS 0.013966f
C434 B.n257 VSUBS 0.013966f
C435 B.n258 VSUBS 0.013966f
C436 B.n259 VSUBS 0.013966f
C437 B.n260 VSUBS 0.013966f
C438 B.n261 VSUBS 0.013966f
C439 B.n262 VSUBS 0.013966f
C440 B.n263 VSUBS 0.013966f
C441 B.n264 VSUBS 0.013966f
C442 B.n265 VSUBS 0.013966f
C443 B.n266 VSUBS 0.013966f
C444 B.n267 VSUBS 0.013966f
C445 B.n268 VSUBS 0.013966f
C446 B.n269 VSUBS 0.013966f
C447 B.n270 VSUBS 0.013966f
C448 B.n271 VSUBS 0.013966f
C449 B.n272 VSUBS 0.013966f
C450 B.n273 VSUBS 0.013966f
C451 B.n274 VSUBS 0.013966f
C452 B.n275 VSUBS 0.013966f
C453 B.n276 VSUBS 0.013966f
C454 B.n277 VSUBS 0.013966f
C455 B.n278 VSUBS 0.013966f
C456 B.n279 VSUBS 0.013966f
C457 B.n280 VSUBS 0.013966f
C458 B.n281 VSUBS 0.013966f
C459 B.n282 VSUBS 0.013966f
C460 B.n283 VSUBS 0.013966f
C461 B.n284 VSUBS 0.013966f
C462 B.n285 VSUBS 0.013966f
C463 B.n286 VSUBS 0.013966f
C464 B.n287 VSUBS 0.013966f
C465 B.n288 VSUBS 0.013966f
C466 B.n289 VSUBS 0.013966f
C467 B.n290 VSUBS 0.013966f
C468 B.n291 VSUBS 0.013966f
C469 B.n292 VSUBS 0.013966f
C470 B.n293 VSUBS 0.013966f
C471 B.n294 VSUBS 0.013966f
C472 B.n295 VSUBS 0.013966f
C473 B.n296 VSUBS 0.013966f
C474 B.n297 VSUBS 0.013966f
C475 B.n298 VSUBS 0.013966f
C476 B.n299 VSUBS 0.013966f
C477 B.n300 VSUBS 0.013966f
C478 B.n301 VSUBS 0.013966f
C479 B.n302 VSUBS 0.013966f
C480 B.n303 VSUBS 0.013966f
C481 B.n304 VSUBS 0.013966f
C482 B.n305 VSUBS 0.013966f
C483 B.n306 VSUBS 0.013966f
C484 B.n307 VSUBS 0.013966f
C485 B.n308 VSUBS 0.013966f
C486 B.n309 VSUBS 0.013966f
C487 B.n310 VSUBS 0.013966f
C488 B.n311 VSUBS 0.013966f
C489 B.n312 VSUBS 0.013966f
C490 B.n313 VSUBS 0.013966f
C491 B.n314 VSUBS 0.013966f
C492 B.n315 VSUBS 0.013966f
C493 B.n316 VSUBS 0.013966f
C494 B.n317 VSUBS 0.013966f
C495 B.n318 VSUBS 0.013966f
C496 B.n319 VSUBS 0.013966f
C497 B.n320 VSUBS 0.013966f
C498 B.n321 VSUBS 0.013966f
C499 B.n322 VSUBS 0.013966f
C500 B.n323 VSUBS 0.013966f
C501 B.n324 VSUBS 0.013966f
C502 B.n325 VSUBS 0.013966f
C503 B.n326 VSUBS 0.013966f
C504 B.n327 VSUBS 0.013966f
C505 B.n328 VSUBS 0.013966f
C506 B.n329 VSUBS 0.013966f
C507 B.n330 VSUBS 0.013966f
C508 B.n331 VSUBS 0.013966f
C509 B.n332 VSUBS 0.032064f
C510 B.n333 VSUBS 0.032064f
C511 B.n334 VSUBS 0.032837f
C512 B.n335 VSUBS 0.013966f
C513 B.n336 VSUBS 0.013966f
C514 B.n337 VSUBS 0.013966f
C515 B.n338 VSUBS 0.013966f
C516 B.n339 VSUBS 0.013966f
C517 B.n340 VSUBS 0.013966f
C518 B.n341 VSUBS 0.013966f
C519 B.n342 VSUBS 0.013966f
C520 B.n343 VSUBS 0.013966f
C521 B.n344 VSUBS 0.013966f
C522 B.n345 VSUBS 0.013966f
C523 B.n346 VSUBS 0.013966f
C524 B.n347 VSUBS 0.013966f
C525 B.n348 VSUBS 0.013966f
C526 B.n349 VSUBS 0.013966f
C527 B.n350 VSUBS 0.013966f
C528 B.n351 VSUBS 0.013966f
C529 B.n352 VSUBS 0.013966f
C530 B.n353 VSUBS 0.013966f
C531 B.n354 VSUBS 0.013966f
C532 B.n355 VSUBS 0.013966f
C533 B.t5 VSUBS 0.17092f
C534 B.t4 VSUBS 0.218711f
C535 B.t3 VSUBS 1.2712f
C536 B.n356 VSUBS 0.188634f
C537 B.n357 VSUBS 0.142996f
C538 B.n358 VSUBS 0.032357f
C539 B.n359 VSUBS 0.013144f
C540 B.n360 VSUBS 0.013966f
C541 B.n361 VSUBS 0.013966f
C542 B.n362 VSUBS 0.013966f
C543 B.n363 VSUBS 0.013966f
C544 B.n364 VSUBS 0.013966f
C545 B.n365 VSUBS 0.013966f
C546 B.n366 VSUBS 0.013966f
C547 B.n367 VSUBS 0.013966f
C548 B.n368 VSUBS 0.013966f
C549 B.n369 VSUBS 0.013966f
C550 B.n370 VSUBS 0.013966f
C551 B.n371 VSUBS 0.013966f
C552 B.n372 VSUBS 0.013966f
C553 B.n373 VSUBS 0.013966f
C554 B.n374 VSUBS 0.013966f
C555 B.n375 VSUBS 0.007804f
C556 B.n376 VSUBS 0.032357f
C557 B.n377 VSUBS 0.013144f
C558 B.n378 VSUBS 0.013966f
C559 B.n379 VSUBS 0.013966f
C560 B.n380 VSUBS 0.013966f
C561 B.n381 VSUBS 0.013966f
C562 B.n382 VSUBS 0.013966f
C563 B.n383 VSUBS 0.013966f
C564 B.n384 VSUBS 0.013966f
C565 B.n385 VSUBS 0.013966f
C566 B.n386 VSUBS 0.013966f
C567 B.n387 VSUBS 0.013966f
C568 B.n388 VSUBS 0.013966f
C569 B.n389 VSUBS 0.013966f
C570 B.n390 VSUBS 0.013966f
C571 B.n391 VSUBS 0.013966f
C572 B.n392 VSUBS 0.013966f
C573 B.n393 VSUBS 0.013966f
C574 B.n394 VSUBS 0.013966f
C575 B.n395 VSUBS 0.013966f
C576 B.n396 VSUBS 0.013966f
C577 B.n397 VSUBS 0.013966f
C578 B.n398 VSUBS 0.013966f
C579 B.n399 VSUBS 0.032837f
C580 B.n400 VSUBS 0.031169f
C581 B.n401 VSUBS 0.033731f
C582 B.n402 VSUBS 0.013966f
C583 B.n403 VSUBS 0.013966f
C584 B.n404 VSUBS 0.013966f
C585 B.n405 VSUBS 0.013966f
C586 B.n406 VSUBS 0.013966f
C587 B.n407 VSUBS 0.013966f
C588 B.n408 VSUBS 0.013966f
C589 B.n409 VSUBS 0.013966f
C590 B.n410 VSUBS 0.013966f
C591 B.n411 VSUBS 0.013966f
C592 B.n412 VSUBS 0.013966f
C593 B.n413 VSUBS 0.013966f
C594 B.n414 VSUBS 0.013966f
C595 B.n415 VSUBS 0.013966f
C596 B.n416 VSUBS 0.013966f
C597 B.n417 VSUBS 0.013966f
C598 B.n418 VSUBS 0.013966f
C599 B.n419 VSUBS 0.013966f
C600 B.n420 VSUBS 0.013966f
C601 B.n421 VSUBS 0.013966f
C602 B.n422 VSUBS 0.013966f
C603 B.n423 VSUBS 0.013966f
C604 B.n424 VSUBS 0.013966f
C605 B.n425 VSUBS 0.013966f
C606 B.n426 VSUBS 0.013966f
C607 B.n427 VSUBS 0.013966f
C608 B.n428 VSUBS 0.013966f
C609 B.n429 VSUBS 0.013966f
C610 B.n430 VSUBS 0.013966f
C611 B.n431 VSUBS 0.013966f
C612 B.n432 VSUBS 0.013966f
C613 B.n433 VSUBS 0.013966f
C614 B.n434 VSUBS 0.013966f
C615 B.n435 VSUBS 0.013966f
C616 B.n436 VSUBS 0.013966f
C617 B.n437 VSUBS 0.013966f
C618 B.n438 VSUBS 0.013966f
C619 B.n439 VSUBS 0.013966f
C620 B.n440 VSUBS 0.013966f
C621 B.n441 VSUBS 0.013966f
C622 B.n442 VSUBS 0.013966f
C623 B.n443 VSUBS 0.013966f
C624 B.n444 VSUBS 0.013966f
C625 B.n445 VSUBS 0.013966f
C626 B.n446 VSUBS 0.013966f
C627 B.n447 VSUBS 0.013966f
C628 B.n448 VSUBS 0.013966f
C629 B.n449 VSUBS 0.013966f
C630 B.n450 VSUBS 0.013966f
C631 B.n451 VSUBS 0.013966f
C632 B.n452 VSUBS 0.013966f
C633 B.n453 VSUBS 0.013966f
C634 B.n454 VSUBS 0.013966f
C635 B.n455 VSUBS 0.013966f
C636 B.n456 VSUBS 0.013966f
C637 B.n457 VSUBS 0.013966f
C638 B.n458 VSUBS 0.013966f
C639 B.n459 VSUBS 0.013966f
C640 B.n460 VSUBS 0.013966f
C641 B.n461 VSUBS 0.013966f
C642 B.n462 VSUBS 0.013966f
C643 B.n463 VSUBS 0.013966f
C644 B.n464 VSUBS 0.013966f
C645 B.n465 VSUBS 0.013966f
C646 B.n466 VSUBS 0.013966f
C647 B.n467 VSUBS 0.013966f
C648 B.n468 VSUBS 0.013966f
C649 B.n469 VSUBS 0.013966f
C650 B.n470 VSUBS 0.013966f
C651 B.n471 VSUBS 0.013966f
C652 B.n472 VSUBS 0.013966f
C653 B.n473 VSUBS 0.013966f
C654 B.n474 VSUBS 0.013966f
C655 B.n475 VSUBS 0.013966f
C656 B.n476 VSUBS 0.013966f
C657 B.n477 VSUBS 0.013966f
C658 B.n478 VSUBS 0.013966f
C659 B.n479 VSUBS 0.013966f
C660 B.n480 VSUBS 0.013966f
C661 B.n481 VSUBS 0.013966f
C662 B.n482 VSUBS 0.013966f
C663 B.n483 VSUBS 0.013966f
C664 B.n484 VSUBS 0.013966f
C665 B.n485 VSUBS 0.013966f
C666 B.n486 VSUBS 0.013966f
C667 B.n487 VSUBS 0.013966f
C668 B.n488 VSUBS 0.013966f
C669 B.n489 VSUBS 0.013966f
C670 B.n490 VSUBS 0.013966f
C671 B.n491 VSUBS 0.013966f
C672 B.n492 VSUBS 0.013966f
C673 B.n493 VSUBS 0.013966f
C674 B.n494 VSUBS 0.013966f
C675 B.n495 VSUBS 0.013966f
C676 B.n496 VSUBS 0.013966f
C677 B.n497 VSUBS 0.013966f
C678 B.n498 VSUBS 0.013966f
C679 B.n499 VSUBS 0.013966f
C680 B.n500 VSUBS 0.013966f
C681 B.n501 VSUBS 0.013966f
C682 B.n502 VSUBS 0.013966f
C683 B.n503 VSUBS 0.013966f
C684 B.n504 VSUBS 0.013966f
C685 B.n505 VSUBS 0.013966f
C686 B.n506 VSUBS 0.013966f
C687 B.n507 VSUBS 0.013966f
C688 B.n508 VSUBS 0.013966f
C689 B.n509 VSUBS 0.013966f
C690 B.n510 VSUBS 0.013966f
C691 B.n511 VSUBS 0.013966f
C692 B.n512 VSUBS 0.013966f
C693 B.n513 VSUBS 0.013966f
C694 B.n514 VSUBS 0.013966f
C695 B.n515 VSUBS 0.013966f
C696 B.n516 VSUBS 0.013966f
C697 B.n517 VSUBS 0.013966f
C698 B.n518 VSUBS 0.013966f
C699 B.n519 VSUBS 0.013966f
C700 B.n520 VSUBS 0.013966f
C701 B.n521 VSUBS 0.013966f
C702 B.n522 VSUBS 0.013966f
C703 B.n523 VSUBS 0.013966f
C704 B.n524 VSUBS 0.013966f
C705 B.n525 VSUBS 0.013966f
C706 B.n526 VSUBS 0.013966f
C707 B.n527 VSUBS 0.013966f
C708 B.n528 VSUBS 0.013966f
C709 B.n529 VSUBS 0.013966f
C710 B.n530 VSUBS 0.013966f
C711 B.n531 VSUBS 0.013966f
C712 B.n532 VSUBS 0.013966f
C713 B.n533 VSUBS 0.013966f
C714 B.n534 VSUBS 0.013966f
C715 B.n535 VSUBS 0.013966f
C716 B.n536 VSUBS 0.013966f
C717 B.n537 VSUBS 0.013966f
C718 B.n538 VSUBS 0.013966f
C719 B.n539 VSUBS 0.013966f
C720 B.n540 VSUBS 0.013966f
C721 B.n541 VSUBS 0.013966f
C722 B.n542 VSUBS 0.013966f
C723 B.n543 VSUBS 0.013966f
C724 B.n544 VSUBS 0.013966f
C725 B.n545 VSUBS 0.013966f
C726 B.n546 VSUBS 0.013966f
C727 B.n547 VSUBS 0.013966f
C728 B.n548 VSUBS 0.013966f
C729 B.n549 VSUBS 0.013966f
C730 B.n550 VSUBS 0.013966f
C731 B.n551 VSUBS 0.013966f
C732 B.n552 VSUBS 0.013966f
C733 B.n553 VSUBS 0.013966f
C734 B.n554 VSUBS 0.013966f
C735 B.n555 VSUBS 0.013966f
C736 B.n556 VSUBS 0.013966f
C737 B.n557 VSUBS 0.013966f
C738 B.n558 VSUBS 0.013966f
C739 B.n559 VSUBS 0.013966f
C740 B.n560 VSUBS 0.013966f
C741 B.n561 VSUBS 0.013966f
C742 B.n562 VSUBS 0.013966f
C743 B.n563 VSUBS 0.013966f
C744 B.n564 VSUBS 0.013966f
C745 B.n565 VSUBS 0.013966f
C746 B.n566 VSUBS 0.013966f
C747 B.n567 VSUBS 0.013966f
C748 B.n568 VSUBS 0.013966f
C749 B.n569 VSUBS 0.013966f
C750 B.n570 VSUBS 0.013966f
C751 B.n571 VSUBS 0.013966f
C752 B.n572 VSUBS 0.013966f
C753 B.n573 VSUBS 0.013966f
C754 B.n574 VSUBS 0.013966f
C755 B.n575 VSUBS 0.013966f
C756 B.n576 VSUBS 0.013966f
C757 B.n577 VSUBS 0.013966f
C758 B.n578 VSUBS 0.013966f
C759 B.n579 VSUBS 0.013966f
C760 B.n580 VSUBS 0.013966f
C761 B.n581 VSUBS 0.013966f
C762 B.n582 VSUBS 0.013966f
C763 B.n583 VSUBS 0.013966f
C764 B.n584 VSUBS 0.013966f
C765 B.n585 VSUBS 0.013966f
C766 B.n586 VSUBS 0.013966f
C767 B.n587 VSUBS 0.013966f
C768 B.n588 VSUBS 0.013966f
C769 B.n589 VSUBS 0.013966f
C770 B.n590 VSUBS 0.013966f
C771 B.n591 VSUBS 0.013966f
C772 B.n592 VSUBS 0.013966f
C773 B.n593 VSUBS 0.013966f
C774 B.n594 VSUBS 0.013966f
C775 B.n595 VSUBS 0.013966f
C776 B.n596 VSUBS 0.013966f
C777 B.n597 VSUBS 0.013966f
C778 B.n598 VSUBS 0.013966f
C779 B.n599 VSUBS 0.013966f
C780 B.n600 VSUBS 0.013966f
C781 B.n601 VSUBS 0.013966f
C782 B.n602 VSUBS 0.013966f
C783 B.n603 VSUBS 0.013966f
C784 B.n604 VSUBS 0.013966f
C785 B.n605 VSUBS 0.013966f
C786 B.n606 VSUBS 0.013966f
C787 B.n607 VSUBS 0.013966f
C788 B.n608 VSUBS 0.013966f
C789 B.n609 VSUBS 0.013966f
C790 B.n610 VSUBS 0.013966f
C791 B.n611 VSUBS 0.013966f
C792 B.n612 VSUBS 0.013966f
C793 B.n613 VSUBS 0.013966f
C794 B.n614 VSUBS 0.013966f
C795 B.n615 VSUBS 0.013966f
C796 B.n616 VSUBS 0.013966f
C797 B.n617 VSUBS 0.013966f
C798 B.n618 VSUBS 0.013966f
C799 B.n619 VSUBS 0.013966f
C800 B.n620 VSUBS 0.013966f
C801 B.n621 VSUBS 0.013966f
C802 B.n622 VSUBS 0.013966f
C803 B.n623 VSUBS 0.013966f
C804 B.n624 VSUBS 0.013966f
C805 B.n625 VSUBS 0.013966f
C806 B.n626 VSUBS 0.013966f
C807 B.n627 VSUBS 0.013966f
C808 B.n628 VSUBS 0.013966f
C809 B.n629 VSUBS 0.013966f
C810 B.n630 VSUBS 0.013966f
C811 B.n631 VSUBS 0.013966f
C812 B.n632 VSUBS 0.013966f
C813 B.n633 VSUBS 0.013966f
C814 B.n634 VSUBS 0.013966f
C815 B.n635 VSUBS 0.013966f
C816 B.n636 VSUBS 0.013966f
C817 B.n637 VSUBS 0.013966f
C818 B.n638 VSUBS 0.013966f
C819 B.n639 VSUBS 0.013966f
C820 B.n640 VSUBS 0.013966f
C821 B.n641 VSUBS 0.013966f
C822 B.n642 VSUBS 0.013966f
C823 B.n643 VSUBS 0.013966f
C824 B.n644 VSUBS 0.013966f
C825 B.n645 VSUBS 0.032064f
C826 B.n646 VSUBS 0.032064f
C827 B.n647 VSUBS 0.032837f
C828 B.n648 VSUBS 0.013966f
C829 B.n649 VSUBS 0.013966f
C830 B.n650 VSUBS 0.013966f
C831 B.n651 VSUBS 0.013966f
C832 B.n652 VSUBS 0.013966f
C833 B.n653 VSUBS 0.013966f
C834 B.n654 VSUBS 0.013966f
C835 B.n655 VSUBS 0.013966f
C836 B.n656 VSUBS 0.013966f
C837 B.n657 VSUBS 0.013966f
C838 B.n658 VSUBS 0.013966f
C839 B.n659 VSUBS 0.013966f
C840 B.n660 VSUBS 0.013966f
C841 B.n661 VSUBS 0.013966f
C842 B.n662 VSUBS 0.013966f
C843 B.n663 VSUBS 0.013966f
C844 B.n664 VSUBS 0.013966f
C845 B.n665 VSUBS 0.013966f
C846 B.n666 VSUBS 0.013966f
C847 B.n667 VSUBS 0.013966f
C848 B.n668 VSUBS 0.013966f
C849 B.n669 VSUBS 0.013966f
C850 B.n670 VSUBS 0.013144f
C851 B.n671 VSUBS 0.032357f
C852 B.n672 VSUBS 0.007804f
C853 B.n673 VSUBS 0.013966f
C854 B.n674 VSUBS 0.013966f
C855 B.n675 VSUBS 0.013966f
C856 B.n676 VSUBS 0.013966f
C857 B.n677 VSUBS 0.013966f
C858 B.n678 VSUBS 0.013966f
C859 B.n679 VSUBS 0.013966f
C860 B.n680 VSUBS 0.013966f
C861 B.n681 VSUBS 0.013966f
C862 B.n682 VSUBS 0.013966f
C863 B.n683 VSUBS 0.013966f
C864 B.n684 VSUBS 0.013966f
C865 B.n685 VSUBS 0.007804f
C866 B.n686 VSUBS 0.013966f
C867 B.n687 VSUBS 0.013966f
C868 B.n688 VSUBS 0.013966f
C869 B.n689 VSUBS 0.013966f
C870 B.n690 VSUBS 0.013966f
C871 B.n691 VSUBS 0.013966f
C872 B.n692 VSUBS 0.013966f
C873 B.n693 VSUBS 0.013966f
C874 B.n694 VSUBS 0.013966f
C875 B.n695 VSUBS 0.013966f
C876 B.n696 VSUBS 0.013966f
C877 B.n697 VSUBS 0.013966f
C878 B.n698 VSUBS 0.013966f
C879 B.n699 VSUBS 0.013966f
C880 B.n700 VSUBS 0.013966f
C881 B.n701 VSUBS 0.013966f
C882 B.n702 VSUBS 0.013966f
C883 B.n703 VSUBS 0.013966f
C884 B.n704 VSUBS 0.013966f
C885 B.n705 VSUBS 0.013966f
C886 B.n706 VSUBS 0.013966f
C887 B.n707 VSUBS 0.013966f
C888 B.n708 VSUBS 0.013966f
C889 B.n709 VSUBS 0.032837f
C890 B.n710 VSUBS 0.032837f
C891 B.n711 VSUBS 0.032064f
C892 B.n712 VSUBS 0.013966f
C893 B.n713 VSUBS 0.013966f
C894 B.n714 VSUBS 0.013966f
C895 B.n715 VSUBS 0.013966f
C896 B.n716 VSUBS 0.013966f
C897 B.n717 VSUBS 0.013966f
C898 B.n718 VSUBS 0.013966f
C899 B.n719 VSUBS 0.013966f
C900 B.n720 VSUBS 0.013966f
C901 B.n721 VSUBS 0.013966f
C902 B.n722 VSUBS 0.013966f
C903 B.n723 VSUBS 0.013966f
C904 B.n724 VSUBS 0.013966f
C905 B.n725 VSUBS 0.013966f
C906 B.n726 VSUBS 0.013966f
C907 B.n727 VSUBS 0.013966f
C908 B.n728 VSUBS 0.013966f
C909 B.n729 VSUBS 0.013966f
C910 B.n730 VSUBS 0.013966f
C911 B.n731 VSUBS 0.013966f
C912 B.n732 VSUBS 0.013966f
C913 B.n733 VSUBS 0.013966f
C914 B.n734 VSUBS 0.013966f
C915 B.n735 VSUBS 0.013966f
C916 B.n736 VSUBS 0.013966f
C917 B.n737 VSUBS 0.013966f
C918 B.n738 VSUBS 0.013966f
C919 B.n739 VSUBS 0.013966f
C920 B.n740 VSUBS 0.013966f
C921 B.n741 VSUBS 0.013966f
C922 B.n742 VSUBS 0.013966f
C923 B.n743 VSUBS 0.013966f
C924 B.n744 VSUBS 0.013966f
C925 B.n745 VSUBS 0.013966f
C926 B.n746 VSUBS 0.013966f
C927 B.n747 VSUBS 0.013966f
C928 B.n748 VSUBS 0.013966f
C929 B.n749 VSUBS 0.013966f
C930 B.n750 VSUBS 0.013966f
C931 B.n751 VSUBS 0.013966f
C932 B.n752 VSUBS 0.013966f
C933 B.n753 VSUBS 0.013966f
C934 B.n754 VSUBS 0.013966f
C935 B.n755 VSUBS 0.013966f
C936 B.n756 VSUBS 0.013966f
C937 B.n757 VSUBS 0.013966f
C938 B.n758 VSUBS 0.013966f
C939 B.n759 VSUBS 0.013966f
C940 B.n760 VSUBS 0.013966f
C941 B.n761 VSUBS 0.013966f
C942 B.n762 VSUBS 0.013966f
C943 B.n763 VSUBS 0.013966f
C944 B.n764 VSUBS 0.013966f
C945 B.n765 VSUBS 0.013966f
C946 B.n766 VSUBS 0.013966f
C947 B.n767 VSUBS 0.013966f
C948 B.n768 VSUBS 0.013966f
C949 B.n769 VSUBS 0.013966f
C950 B.n770 VSUBS 0.013966f
C951 B.n771 VSUBS 0.013966f
C952 B.n772 VSUBS 0.013966f
C953 B.n773 VSUBS 0.013966f
C954 B.n774 VSUBS 0.013966f
C955 B.n775 VSUBS 0.013966f
C956 B.n776 VSUBS 0.013966f
C957 B.n777 VSUBS 0.013966f
C958 B.n778 VSUBS 0.013966f
C959 B.n779 VSUBS 0.013966f
C960 B.n780 VSUBS 0.013966f
C961 B.n781 VSUBS 0.013966f
C962 B.n782 VSUBS 0.013966f
C963 B.n783 VSUBS 0.013966f
C964 B.n784 VSUBS 0.013966f
C965 B.n785 VSUBS 0.013966f
C966 B.n786 VSUBS 0.013966f
C967 B.n787 VSUBS 0.013966f
C968 B.n788 VSUBS 0.013966f
C969 B.n789 VSUBS 0.013966f
C970 B.n790 VSUBS 0.013966f
C971 B.n791 VSUBS 0.013966f
C972 B.n792 VSUBS 0.013966f
C973 B.n793 VSUBS 0.013966f
C974 B.n794 VSUBS 0.013966f
C975 B.n795 VSUBS 0.013966f
C976 B.n796 VSUBS 0.013966f
C977 B.n797 VSUBS 0.013966f
C978 B.n798 VSUBS 0.013966f
C979 B.n799 VSUBS 0.013966f
C980 B.n800 VSUBS 0.013966f
C981 B.n801 VSUBS 0.013966f
C982 B.n802 VSUBS 0.013966f
C983 B.n803 VSUBS 0.013966f
C984 B.n804 VSUBS 0.013966f
C985 B.n805 VSUBS 0.013966f
C986 B.n806 VSUBS 0.013966f
C987 B.n807 VSUBS 0.013966f
C988 B.n808 VSUBS 0.013966f
C989 B.n809 VSUBS 0.013966f
C990 B.n810 VSUBS 0.013966f
C991 B.n811 VSUBS 0.013966f
C992 B.n812 VSUBS 0.013966f
C993 B.n813 VSUBS 0.013966f
C994 B.n814 VSUBS 0.013966f
C995 B.n815 VSUBS 0.013966f
C996 B.n816 VSUBS 0.013966f
C997 B.n817 VSUBS 0.013966f
C998 B.n818 VSUBS 0.013966f
C999 B.n819 VSUBS 0.013966f
C1000 B.n820 VSUBS 0.013966f
C1001 B.n821 VSUBS 0.013966f
C1002 B.n822 VSUBS 0.013966f
C1003 B.n823 VSUBS 0.013966f
C1004 B.n824 VSUBS 0.013966f
C1005 B.n825 VSUBS 0.013966f
C1006 B.n826 VSUBS 0.013966f
C1007 B.n827 VSUBS 0.013966f
C1008 B.n828 VSUBS 0.013966f
C1009 B.n829 VSUBS 0.013966f
C1010 B.n830 VSUBS 0.013966f
C1011 B.n831 VSUBS 0.018225f
C1012 B.n832 VSUBS 0.019414f
C1013 B.n833 VSUBS 0.038606f
C1014 VDD1.t2 VSUBS 0.853959f
C1015 VDD1.t5 VSUBS 0.106891f
C1016 VDD1.t9 VSUBS 0.106891f
C1017 VDD1.n0 VSUBS 0.591461f
C1018 VDD1.n1 VSUBS 2.13441f
C1019 VDD1.t7 VSUBS 0.853956f
C1020 VDD1.t0 VSUBS 0.106891f
C1021 VDD1.t6 VSUBS 0.106891f
C1022 VDD1.n2 VSUBS 0.591458f
C1023 VDD1.n3 VSUBS 2.121f
C1024 VDD1.t1 VSUBS 0.106891f
C1025 VDD1.t8 VSUBS 0.106891f
C1026 VDD1.n4 VSUBS 0.620432f
C1027 VDD1.n5 VSUBS 5.23684f
C1028 VDD1.t3 VSUBS 0.106891f
C1029 VDD1.t4 VSUBS 0.106891f
C1030 VDD1.n6 VSUBS 0.591458f
C1031 VDD1.n7 VSUBS 4.99262f
C1032 VTAIL.t0 VSUBS 0.108577f
C1033 VTAIL.t7 VSUBS 0.108577f
C1034 VTAIL.n0 VSUBS 0.514474f
C1035 VTAIL.n1 VSUBS 1.21557f
C1036 VTAIL.t19 VSUBS 0.750524f
C1037 VTAIL.n2 VSUBS 1.38421f
C1038 VTAIL.t11 VSUBS 0.108577f
C1039 VTAIL.t15 VSUBS 0.108577f
C1040 VTAIL.n3 VSUBS 0.514474f
C1041 VTAIL.n4 VSUBS 1.49539f
C1042 VTAIL.t17 VSUBS 0.108577f
C1043 VTAIL.t14 VSUBS 0.108577f
C1044 VTAIL.n5 VSUBS 0.514474f
C1045 VTAIL.n6 VSUBS 2.88887f
C1046 VTAIL.t8 VSUBS 0.108577f
C1047 VTAIL.t3 VSUBS 0.108577f
C1048 VTAIL.n7 VSUBS 0.514477f
C1049 VTAIL.n8 VSUBS 2.88887f
C1050 VTAIL.t6 VSUBS 0.108577f
C1051 VTAIL.t1 VSUBS 0.108577f
C1052 VTAIL.n9 VSUBS 0.514477f
C1053 VTAIL.n10 VSUBS 1.49538f
C1054 VTAIL.t2 VSUBS 0.750528f
C1055 VTAIL.n11 VSUBS 1.38421f
C1056 VTAIL.t16 VSUBS 0.108577f
C1057 VTAIL.t12 VSUBS 0.108577f
C1058 VTAIL.n12 VSUBS 0.514477f
C1059 VTAIL.n13 VSUBS 1.32414f
C1060 VTAIL.t13 VSUBS 0.108577f
C1061 VTAIL.t10 VSUBS 0.108577f
C1062 VTAIL.n14 VSUBS 0.514477f
C1063 VTAIL.n15 VSUBS 1.49538f
C1064 VTAIL.t18 VSUBS 0.750524f
C1065 VTAIL.n16 VSUBS 2.48445f
C1066 VTAIL.t5 VSUBS 0.750524f
C1067 VTAIL.n17 VSUBS 2.48445f
C1068 VTAIL.t9 VSUBS 0.108577f
C1069 VTAIL.t4 VSUBS 0.108577f
C1070 VTAIL.n18 VSUBS 0.514474f
C1071 VTAIL.n19 VSUBS 1.13947f
C1072 VP.t1 VSUBS 1.45591f
C1073 VP.n0 VSUBS 0.74427f
C1074 VP.n1 VSUBS 0.044203f
C1075 VP.n2 VSUBS 0.088776f
C1076 VP.n3 VSUBS 0.044203f
C1077 VP.n4 VSUBS 0.082383f
C1078 VP.n5 VSUBS 0.044203f
C1079 VP.t8 VSUBS 1.45591f
C1080 VP.n6 VSUBS 0.082383f
C1081 VP.n7 VSUBS 0.044203f
C1082 VP.n8 VSUBS 0.082383f
C1083 VP.n9 VSUBS 0.044203f
C1084 VP.t3 VSUBS 1.45591f
C1085 VP.n10 VSUBS 0.082383f
C1086 VP.n11 VSUBS 0.044203f
C1087 VP.n12 VSUBS 0.082383f
C1088 VP.n13 VSUBS 0.044203f
C1089 VP.t9 VSUBS 1.45591f
C1090 VP.n14 VSUBS 0.082383f
C1091 VP.n15 VSUBS 0.044203f
C1092 VP.n16 VSUBS 0.082383f
C1093 VP.n17 VSUBS 0.071342f
C1094 VP.t2 VSUBS 1.45591f
C1095 VP.t5 VSUBS 1.45591f
C1096 VP.n18 VSUBS 0.74427f
C1097 VP.n19 VSUBS 0.044203f
C1098 VP.n20 VSUBS 0.088776f
C1099 VP.n21 VSUBS 0.044203f
C1100 VP.n22 VSUBS 0.082383f
C1101 VP.n23 VSUBS 0.044203f
C1102 VP.t6 VSUBS 1.45591f
C1103 VP.n24 VSUBS 0.082383f
C1104 VP.n25 VSUBS 0.044203f
C1105 VP.n26 VSUBS 0.082383f
C1106 VP.n27 VSUBS 0.044203f
C1107 VP.t0 VSUBS 1.45591f
C1108 VP.n28 VSUBS 0.082383f
C1109 VP.n29 VSUBS 0.044203f
C1110 VP.n30 VSUBS 0.082383f
C1111 VP.t7 VSUBS 2.01838f
C1112 VP.n31 VSUBS 0.774134f
C1113 VP.t4 VSUBS 1.45591f
C1114 VP.n32 VSUBS 0.750701f
C1115 VP.n33 VSUBS 0.074248f
C1116 VP.n34 VSUBS 0.569735f
C1117 VP.n35 VSUBS 0.044203f
C1118 VP.n36 VSUBS 0.044203f
C1119 VP.n37 VSUBS 0.082383f
C1120 VP.n38 VSUBS 0.055294f
C1121 VP.n39 VSUBS 0.07377f
C1122 VP.n40 VSUBS 0.044203f
C1123 VP.n41 VSUBS 0.044203f
C1124 VP.n42 VSUBS 0.044203f
C1125 VP.n43 VSUBS 0.082383f
C1126 VP.n44 VSUBS 0.062046f
C1127 VP.n45 VSUBS 0.578555f
C1128 VP.n46 VSUBS 0.062046f
C1129 VP.n47 VSUBS 0.044203f
C1130 VP.n48 VSUBS 0.044203f
C1131 VP.n49 VSUBS 0.044203f
C1132 VP.n50 VSUBS 0.082383f
C1133 VP.n51 VSUBS 0.07377f
C1134 VP.n52 VSUBS 0.055294f
C1135 VP.n53 VSUBS 0.044203f
C1136 VP.n54 VSUBS 0.044203f
C1137 VP.n55 VSUBS 0.044203f
C1138 VP.n56 VSUBS 0.082383f
C1139 VP.n57 VSUBS 0.074248f
C1140 VP.n58 VSUBS 0.578555f
C1141 VP.n59 VSUBS 0.049845f
C1142 VP.n60 VSUBS 0.044203f
C1143 VP.n61 VSUBS 0.044203f
C1144 VP.n62 VSUBS 0.044203f
C1145 VP.n63 VSUBS 0.082383f
C1146 VP.n64 VSUBS 0.08658f
C1147 VP.n65 VSUBS 0.036092f
C1148 VP.n66 VSUBS 0.044203f
C1149 VP.n67 VSUBS 0.044203f
C1150 VP.n68 VSUBS 0.044203f
C1151 VP.n69 VSUBS 0.082383f
C1152 VP.n70 VSUBS 0.082383f
C1153 VP.n71 VSUBS 0.045777f
C1154 VP.n72 VSUBS 0.071342f
C1155 VP.n73 VSUBS 2.78274f
C1156 VP.n74 VSUBS 2.81255f
C1157 VP.n75 VSUBS 0.74427f
C1158 VP.n76 VSUBS 0.045777f
C1159 VP.n77 VSUBS 0.082383f
C1160 VP.n78 VSUBS 0.044203f
C1161 VP.n79 VSUBS 0.044203f
C1162 VP.n80 VSUBS 0.044203f
C1163 VP.n81 VSUBS 0.088776f
C1164 VP.n82 VSUBS 0.036092f
C1165 VP.n83 VSUBS 0.08658f
C1166 VP.n84 VSUBS 0.044203f
C1167 VP.n85 VSUBS 0.044203f
C1168 VP.n86 VSUBS 0.044203f
C1169 VP.n87 VSUBS 0.082383f
C1170 VP.n88 VSUBS 0.049845f
C1171 VP.n89 VSUBS 0.578555f
C1172 VP.n90 VSUBS 0.074248f
C1173 VP.n91 VSUBS 0.044203f
C1174 VP.n92 VSUBS 0.044203f
C1175 VP.n93 VSUBS 0.044203f
C1176 VP.n94 VSUBS 0.082383f
C1177 VP.n95 VSUBS 0.055294f
C1178 VP.n96 VSUBS 0.07377f
C1179 VP.n97 VSUBS 0.044203f
C1180 VP.n98 VSUBS 0.044203f
C1181 VP.n99 VSUBS 0.044203f
C1182 VP.n100 VSUBS 0.082383f
C1183 VP.n101 VSUBS 0.062046f
C1184 VP.n102 VSUBS 0.578555f
C1185 VP.n103 VSUBS 0.062046f
C1186 VP.n104 VSUBS 0.044203f
C1187 VP.n105 VSUBS 0.044203f
C1188 VP.n106 VSUBS 0.044203f
C1189 VP.n107 VSUBS 0.082383f
C1190 VP.n108 VSUBS 0.07377f
C1191 VP.n109 VSUBS 0.055294f
C1192 VP.n110 VSUBS 0.044203f
C1193 VP.n111 VSUBS 0.044203f
C1194 VP.n112 VSUBS 0.044203f
C1195 VP.n113 VSUBS 0.082383f
C1196 VP.n114 VSUBS 0.074248f
C1197 VP.n115 VSUBS 0.578555f
C1198 VP.n116 VSUBS 0.049845f
C1199 VP.n117 VSUBS 0.044203f
C1200 VP.n118 VSUBS 0.044203f
C1201 VP.n119 VSUBS 0.044203f
C1202 VP.n120 VSUBS 0.082383f
C1203 VP.n121 VSUBS 0.08658f
C1204 VP.n122 VSUBS 0.036092f
C1205 VP.n123 VSUBS 0.044203f
C1206 VP.n124 VSUBS 0.044203f
C1207 VP.n125 VSUBS 0.044203f
C1208 VP.n126 VSUBS 0.082383f
C1209 VP.n127 VSUBS 0.082383f
C1210 VP.n128 VSUBS 0.045777f
C1211 VP.n129 VSUBS 0.071342f
C1212 VP.n130 VSUBS 0.136858f
.ends

