* NGSPICE file created from tg_sample_0005.ext - technology: sky130A

.subckt tg_sample_0005 VIN VGN VGP VSS VCC VOUT
X0 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=0.37
X1 VOUT.t3 VGN.t0 VIN.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=1.6665 pd=10.43 as=3.939 ps=20.98 w=10.1 l=2.14
X2 VSS.t9 VSS.t6 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=2.14
X3 VIN.t0 VGP.t0 VOUT.t0 VCC.t8 sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=1.96515 ps=12.24 w=11.91 l=0.37
X4 VSS.t5 VSS.t2 VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=3.939 pd=20.98 as=0 ps=0 w=10.1 l=2.14
X5 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=0.37
X6 VOUT.t1 VGP.t1 VIN.t1 VCC.t9 sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=4.6449 ps=24.6 w=11.91 l=0.37
X7 VIN.t3 VGN.t1 VOUT.t2 VSS.t0 sky130_fd_pr__nfet_01v8 ad=3.939 pd=20.98 as=1.6665 ps=10.43 w=10.1 l=2.14
R0 VCC.n192 VCC.t0 986.402
R1 VCC.n54 VCC.t4 986.402
R2 VCC.n279 VCC.n9 421.464
R3 VCC.n277 VCC.n12 421.464
R4 VCC.n138 VCC.n32 421.464
R5 VCC.n134 VCC.n28 421.464
R6 VCC.n192 VCC.t2 387.361
R7 VCC.n54 VCC.t7 387.361
R8 VCC.n193 VCC.t3 373.784
R9 VCC.n55 VCC.t6 373.784
R10 VCC.n277 VCC.n276 185
R11 VCC.n278 VCC.n277 185
R12 VCC.n13 VCC.n11 185
R13 VCC.n165 VCC.n11 185
R14 VCC.n169 VCC.n168 185
R15 VCC.n168 VCC.n167 185
R16 VCC.n16 VCC.n15 185
R17 VCC.n164 VCC.n16 185
R18 VCC.n162 VCC.n161 185
R19 VCC.n163 VCC.n162 185
R20 VCC.n18 VCC.n17 185
R21 VCC.n23 VCC.n17 185
R22 VCC.n157 VCC.n156 185
R23 VCC.n156 VCC.n155 185
R24 VCC.n21 VCC.n20 185
R25 VCC.n22 VCC.n21 185
R26 VCC.n144 VCC.n143 185
R27 VCC.n145 VCC.n144 185
R28 VCC.n30 VCC.n29 185
R29 VCC.n146 VCC.n29 185
R30 VCC.n139 VCC.n138 185
R31 VCC.n138 VCC.n137 185
R32 VCC.n28 VCC.n27 185
R33 VCC.n137 VCC.n28 185
R34 VCC.n148 VCC.n147 185
R35 VCC.n147 VCC.n146 185
R36 VCC.n25 VCC.n24 185
R37 VCC.n145 VCC.n24 185
R38 VCC.n153 VCC.n152 185
R39 VCC.n153 VCC.n22 185
R40 VCC.n154 VCC.n2 185
R41 VCC.n155 VCC.n154 185
R42 VCC.n287 VCC.n3 185
R43 VCC.n23 VCC.n3 185
R44 VCC.n286 VCC.n4 185
R45 VCC.n163 VCC.n4 185
R46 VCC.n285 VCC.n5 185
R47 VCC.n164 VCC.n5 185
R48 VCC.n166 VCC.n6 185
R49 VCC.n167 VCC.n166 185
R50 VCC.n281 VCC.n8 185
R51 VCC.n165 VCC.n8 185
R52 VCC.n280 VCC.n279 185
R53 VCC.n279 VCC.n278 185
R54 VCC.n274 VCC.n12 185
R55 VCC.n273 VCC.n272 185
R56 VCC.n270 VCC.n172 185
R57 VCC.n268 VCC.n267 185
R58 VCC.n266 VCC.n173 185
R59 VCC.n265 VCC.n264 185
R60 VCC.n262 VCC.n174 185
R61 VCC.n260 VCC.n259 185
R62 VCC.n258 VCC.n175 185
R63 VCC.n257 VCC.n256 185
R64 VCC.n254 VCC.n176 185
R65 VCC.n252 VCC.n251 185
R66 VCC.n250 VCC.n177 185
R67 VCC.n249 VCC.n248 185
R68 VCC.n246 VCC.n178 185
R69 VCC.n244 VCC.n243 185
R70 VCC.n242 VCC.n179 185
R71 VCC.n241 VCC.n240 185
R72 VCC.n238 VCC.n180 185
R73 VCC.n236 VCC.n235 185
R74 VCC.n234 VCC.n181 185
R75 VCC.n233 VCC.n232 185
R76 VCC.n230 VCC.n182 185
R77 VCC.n228 VCC.n227 185
R78 VCC.n226 VCC.n183 185
R79 VCC.n225 VCC.n224 185
R80 VCC.n222 VCC.n184 185
R81 VCC.n220 VCC.n219 185
R82 VCC.n218 VCC.n185 185
R83 VCC.n217 VCC.n216 185
R84 VCC.n214 VCC.n186 185
R85 VCC.n212 VCC.n211 185
R86 VCC.n210 VCC.n187 185
R87 VCC.n209 VCC.n208 185
R88 VCC.n206 VCC.n188 185
R89 VCC.n204 VCC.n203 185
R90 VCC.n202 VCC.n189 185
R91 VCC.n201 VCC.n200 185
R92 VCC.n198 VCC.n190 185
R93 VCC.n196 VCC.n195 185
R94 VCC.n191 VCC.n9 185
R95 VCC.n10 VCC.n9 185
R96 VCC.n134 VCC.n133 185
R97 VCC.n132 VCC.n53 185
R98 VCC.n130 VCC.n52 185
R99 VCC.n136 VCC.n52 185
R100 VCC.n129 VCC.n128 185
R101 VCC.n127 VCC.n126 185
R102 VCC.n125 VCC.n124 185
R103 VCC.n123 VCC.n122 185
R104 VCC.n121 VCC.n120 185
R105 VCC.n119 VCC.n118 185
R106 VCC.n117 VCC.n116 185
R107 VCC.n115 VCC.n114 185
R108 VCC.n113 VCC.n112 185
R109 VCC.n111 VCC.n110 185
R110 VCC.n109 VCC.n108 185
R111 VCC.n107 VCC.n106 185
R112 VCC.n105 VCC.n104 185
R113 VCC.n103 VCC.n102 185
R114 VCC.n101 VCC.n100 185
R115 VCC.n99 VCC.n98 185
R116 VCC.n97 VCC.n96 185
R117 VCC.n95 VCC.n94 185
R118 VCC.n93 VCC.n92 185
R119 VCC.n91 VCC.n90 185
R120 VCC.n89 VCC.n88 185
R121 VCC.n87 VCC.n86 185
R122 VCC.n85 VCC.n84 185
R123 VCC.n83 VCC.n82 185
R124 VCC.n81 VCC.n80 185
R125 VCC.n79 VCC.n78 185
R126 VCC.n77 VCC.n76 185
R127 VCC.n75 VCC.n74 185
R128 VCC.n73 VCC.n72 185
R129 VCC.n71 VCC.n70 185
R130 VCC.n69 VCC.n68 185
R131 VCC.n67 VCC.n66 185
R132 VCC.n65 VCC.n64 185
R133 VCC.n63 VCC.n62 185
R134 VCC.n61 VCC.n60 185
R135 VCC.n59 VCC.n58 185
R136 VCC.n57 VCC.n56 185
R137 VCC.n32 VCC.n31 185
R138 VCC.n138 VCC.n29 146.341
R139 VCC.n144 VCC.n29 146.341
R140 VCC.n144 VCC.n21 146.341
R141 VCC.n156 VCC.n21 146.341
R142 VCC.n156 VCC.n17 146.341
R143 VCC.n162 VCC.n17 146.341
R144 VCC.n162 VCC.n16 146.341
R145 VCC.n168 VCC.n16 146.341
R146 VCC.n168 VCC.n11 146.341
R147 VCC.n277 VCC.n11 146.341
R148 VCC.n147 VCC.n28 146.341
R149 VCC.n147 VCC.n24 146.341
R150 VCC.n153 VCC.n24 146.341
R151 VCC.n154 VCC.n153 146.341
R152 VCC.n154 VCC.n3 146.341
R153 VCC.n4 VCC.n3 146.341
R154 VCC.n5 VCC.n4 146.341
R155 VCC.n166 VCC.n5 146.341
R156 VCC.n166 VCC.n8 146.341
R157 VCC.n279 VCC.n8 146.341
R158 VCC.n196 VCC.n9 99.5127
R159 VCC.n200 VCC.n198 99.5127
R160 VCC.n204 VCC.n189 99.5127
R161 VCC.n208 VCC.n206 99.5127
R162 VCC.n212 VCC.n187 99.5127
R163 VCC.n216 VCC.n214 99.5127
R164 VCC.n220 VCC.n185 99.5127
R165 VCC.n224 VCC.n222 99.5127
R166 VCC.n228 VCC.n183 99.5127
R167 VCC.n232 VCC.n230 99.5127
R168 VCC.n236 VCC.n181 99.5127
R169 VCC.n240 VCC.n238 99.5127
R170 VCC.n244 VCC.n179 99.5127
R171 VCC.n248 VCC.n246 99.5127
R172 VCC.n252 VCC.n177 99.5127
R173 VCC.n256 VCC.n254 99.5127
R174 VCC.n260 VCC.n175 99.5127
R175 VCC.n264 VCC.n262 99.5127
R176 VCC.n268 VCC.n173 99.5127
R177 VCC.n272 VCC.n270 99.5127
R178 VCC.n53 VCC.n52 99.5127
R179 VCC.n128 VCC.n52 99.5127
R180 VCC.n126 VCC.n125 99.5127
R181 VCC.n122 VCC.n121 99.5127
R182 VCC.n118 VCC.n117 99.5127
R183 VCC.n114 VCC.n113 99.5127
R184 VCC.n110 VCC.n109 99.5127
R185 VCC.n106 VCC.n105 99.5127
R186 VCC.n102 VCC.n101 99.5127
R187 VCC.n98 VCC.n97 99.5127
R188 VCC.n94 VCC.n93 99.5127
R189 VCC.n90 VCC.n89 99.5127
R190 VCC.n86 VCC.n85 99.5127
R191 VCC.n82 VCC.n81 99.5127
R192 VCC.n78 VCC.n77 99.5127
R193 VCC.n74 VCC.n73 99.5127
R194 VCC.n70 VCC.n69 99.5127
R195 VCC.n66 VCC.n65 99.5127
R196 VCC.n62 VCC.n61 99.5127
R197 VCC.n58 VCC.n57 99.5127
R198 VCC.n271 VCC.n10 72.8958
R199 VCC.n269 VCC.n10 72.8958
R200 VCC.n263 VCC.n10 72.8958
R201 VCC.n261 VCC.n10 72.8958
R202 VCC.n255 VCC.n10 72.8958
R203 VCC.n253 VCC.n10 72.8958
R204 VCC.n247 VCC.n10 72.8958
R205 VCC.n245 VCC.n10 72.8958
R206 VCC.n239 VCC.n10 72.8958
R207 VCC.n237 VCC.n10 72.8958
R208 VCC.n231 VCC.n10 72.8958
R209 VCC.n229 VCC.n10 72.8958
R210 VCC.n223 VCC.n10 72.8958
R211 VCC.n221 VCC.n10 72.8958
R212 VCC.n215 VCC.n10 72.8958
R213 VCC.n213 VCC.n10 72.8958
R214 VCC.n207 VCC.n10 72.8958
R215 VCC.n205 VCC.n10 72.8958
R216 VCC.n199 VCC.n10 72.8958
R217 VCC.n197 VCC.n10 72.8958
R218 VCC.n136 VCC.n135 72.8958
R219 VCC.n136 VCC.n33 72.8958
R220 VCC.n136 VCC.n34 72.8958
R221 VCC.n136 VCC.n35 72.8958
R222 VCC.n136 VCC.n36 72.8958
R223 VCC.n136 VCC.n37 72.8958
R224 VCC.n136 VCC.n38 72.8958
R225 VCC.n136 VCC.n39 72.8958
R226 VCC.n136 VCC.n40 72.8958
R227 VCC.n136 VCC.n41 72.8958
R228 VCC.n136 VCC.n42 72.8958
R229 VCC.n136 VCC.n43 72.8958
R230 VCC.n136 VCC.n44 72.8958
R231 VCC.n136 VCC.n45 72.8958
R232 VCC.n136 VCC.n46 72.8958
R233 VCC.n136 VCC.n47 72.8958
R234 VCC.n136 VCC.n48 72.8958
R235 VCC.n136 VCC.n49 72.8958
R236 VCC.n136 VCC.n50 72.8958
R237 VCC.n136 VCC.n51 72.8958
R238 VCC.n137 VCC.n136 56.3363
R239 VCC.n278 VCC.n10 56.3363
R240 VCC.n198 VCC.n197 39.2114
R241 VCC.n199 VCC.n189 39.2114
R242 VCC.n206 VCC.n205 39.2114
R243 VCC.n207 VCC.n187 39.2114
R244 VCC.n214 VCC.n213 39.2114
R245 VCC.n215 VCC.n185 39.2114
R246 VCC.n222 VCC.n221 39.2114
R247 VCC.n223 VCC.n183 39.2114
R248 VCC.n230 VCC.n229 39.2114
R249 VCC.n231 VCC.n181 39.2114
R250 VCC.n238 VCC.n237 39.2114
R251 VCC.n239 VCC.n179 39.2114
R252 VCC.n246 VCC.n245 39.2114
R253 VCC.n247 VCC.n177 39.2114
R254 VCC.n254 VCC.n253 39.2114
R255 VCC.n255 VCC.n175 39.2114
R256 VCC.n262 VCC.n261 39.2114
R257 VCC.n263 VCC.n173 39.2114
R258 VCC.n270 VCC.n269 39.2114
R259 VCC.n271 VCC.n12 39.2114
R260 VCC.n135 VCC.n134 39.2114
R261 VCC.n128 VCC.n33 39.2114
R262 VCC.n125 VCC.n34 39.2114
R263 VCC.n121 VCC.n35 39.2114
R264 VCC.n117 VCC.n36 39.2114
R265 VCC.n113 VCC.n37 39.2114
R266 VCC.n109 VCC.n38 39.2114
R267 VCC.n105 VCC.n39 39.2114
R268 VCC.n101 VCC.n40 39.2114
R269 VCC.n97 VCC.n41 39.2114
R270 VCC.n93 VCC.n42 39.2114
R271 VCC.n89 VCC.n43 39.2114
R272 VCC.n85 VCC.n44 39.2114
R273 VCC.n81 VCC.n45 39.2114
R274 VCC.n77 VCC.n46 39.2114
R275 VCC.n73 VCC.n47 39.2114
R276 VCC.n69 VCC.n48 39.2114
R277 VCC.n65 VCC.n49 39.2114
R278 VCC.n61 VCC.n50 39.2114
R279 VCC.n57 VCC.n51 39.2114
R280 VCC.n272 VCC.n271 39.2114
R281 VCC.n269 VCC.n268 39.2114
R282 VCC.n264 VCC.n263 39.2114
R283 VCC.n261 VCC.n260 39.2114
R284 VCC.n256 VCC.n255 39.2114
R285 VCC.n253 VCC.n252 39.2114
R286 VCC.n248 VCC.n247 39.2114
R287 VCC.n245 VCC.n244 39.2114
R288 VCC.n240 VCC.n239 39.2114
R289 VCC.n237 VCC.n236 39.2114
R290 VCC.n232 VCC.n231 39.2114
R291 VCC.n229 VCC.n228 39.2114
R292 VCC.n224 VCC.n223 39.2114
R293 VCC.n221 VCC.n220 39.2114
R294 VCC.n216 VCC.n215 39.2114
R295 VCC.n213 VCC.n212 39.2114
R296 VCC.n208 VCC.n207 39.2114
R297 VCC.n205 VCC.n204 39.2114
R298 VCC.n200 VCC.n199 39.2114
R299 VCC.n197 VCC.n196 39.2114
R300 VCC.n135 VCC.n53 39.2114
R301 VCC.n126 VCC.n33 39.2114
R302 VCC.n122 VCC.n34 39.2114
R303 VCC.n118 VCC.n35 39.2114
R304 VCC.n114 VCC.n36 39.2114
R305 VCC.n110 VCC.n37 39.2114
R306 VCC.n106 VCC.n38 39.2114
R307 VCC.n102 VCC.n39 39.2114
R308 VCC.n98 VCC.n40 39.2114
R309 VCC.n94 VCC.n41 39.2114
R310 VCC.n90 VCC.n42 39.2114
R311 VCC.n86 VCC.n43 39.2114
R312 VCC.n82 VCC.n44 39.2114
R313 VCC.n78 VCC.n45 39.2114
R314 VCC.n74 VCC.n46 39.2114
R315 VCC.n70 VCC.n47 39.2114
R316 VCC.n66 VCC.n48 39.2114
R317 VCC.n62 VCC.n49 39.2114
R318 VCC.n58 VCC.n50 39.2114
R319 VCC.n51 VCC.n32 39.2114
R320 VCC.n191 VCC.n7 31.2877
R321 VCC.n275 VCC.n274 31.2877
R322 VCC.n133 VCC.n26 31.2877
R323 VCC.n140 VCC.n31 31.2877
R324 VCC.n146 VCC.n145 29.6509
R325 VCC.n145 VCC.n22 29.6509
R326 VCC.n155 VCC.n22 29.6509
R327 VCC.n164 VCC.n163 29.6509
R328 VCC.n167 VCC.n164 29.6509
R329 VCC.n167 VCC.n165 29.6509
R330 VCC.n194 VCC.n193 29.2853
R331 VCC.n131 VCC.n55 29.2853
R332 VCC.n137 VCC.t5 21.3488
R333 VCC.n278 VCC.t1 21.3488
R334 VCC.t8 VCC.n23 20.7558
R335 VCC.n23 VCC.t9 20.7558
R336 VCC.n139 VCC.n30 19.3944
R337 VCC.n143 VCC.n30 19.3944
R338 VCC.n143 VCC.n20 19.3944
R339 VCC.n157 VCC.n20 19.3944
R340 VCC.n157 VCC.n18 19.3944
R341 VCC.n161 VCC.n18 19.3944
R342 VCC.n161 VCC.n15 19.3944
R343 VCC.n169 VCC.n15 19.3944
R344 VCC.n169 VCC.n13 19.3944
R345 VCC.n276 VCC.n13 19.3944
R346 VCC.n148 VCC.n27 19.3944
R347 VCC.n148 VCC.n25 19.3944
R348 VCC.n152 VCC.n25 19.3944
R349 VCC.n152 VCC.n2 19.3944
R350 VCC.n287 VCC.n2 19.3944
R351 VCC.n287 VCC.n286 19.3944
R352 VCC.n286 VCC.n285 19.3944
R353 VCC.n285 VCC.n6 19.3944
R354 VCC.n281 VCC.n6 19.3944
R355 VCC.n281 VCC.n280 19.3944
R356 VCC.n193 VCC.n192 13.5763
R357 VCC.n55 VCC.n54 13.5763
R358 VCC.n195 VCC.n191 10.6151
R359 VCC.n201 VCC.n190 10.6151
R360 VCC.n202 VCC.n201 10.6151
R361 VCC.n203 VCC.n202 10.6151
R362 VCC.n203 VCC.n188 10.6151
R363 VCC.n209 VCC.n188 10.6151
R364 VCC.n210 VCC.n209 10.6151
R365 VCC.n211 VCC.n210 10.6151
R366 VCC.n211 VCC.n186 10.6151
R367 VCC.n217 VCC.n186 10.6151
R368 VCC.n218 VCC.n217 10.6151
R369 VCC.n219 VCC.n218 10.6151
R370 VCC.n219 VCC.n184 10.6151
R371 VCC.n225 VCC.n184 10.6151
R372 VCC.n226 VCC.n225 10.6151
R373 VCC.n227 VCC.n226 10.6151
R374 VCC.n227 VCC.n182 10.6151
R375 VCC.n233 VCC.n182 10.6151
R376 VCC.n234 VCC.n233 10.6151
R377 VCC.n235 VCC.n234 10.6151
R378 VCC.n235 VCC.n180 10.6151
R379 VCC.n241 VCC.n180 10.6151
R380 VCC.n242 VCC.n241 10.6151
R381 VCC.n243 VCC.n242 10.6151
R382 VCC.n243 VCC.n178 10.6151
R383 VCC.n249 VCC.n178 10.6151
R384 VCC.n250 VCC.n249 10.6151
R385 VCC.n251 VCC.n250 10.6151
R386 VCC.n251 VCC.n176 10.6151
R387 VCC.n257 VCC.n176 10.6151
R388 VCC.n258 VCC.n257 10.6151
R389 VCC.n259 VCC.n258 10.6151
R390 VCC.n259 VCC.n174 10.6151
R391 VCC.n265 VCC.n174 10.6151
R392 VCC.n266 VCC.n265 10.6151
R393 VCC.n267 VCC.n266 10.6151
R394 VCC.n267 VCC.n172 10.6151
R395 VCC.n273 VCC.n172 10.6151
R396 VCC.n274 VCC.n273 10.6151
R397 VCC.n133 VCC.n132 10.6151
R398 VCC.n130 VCC.n129 10.6151
R399 VCC.n129 VCC.n127 10.6151
R400 VCC.n127 VCC.n124 10.6151
R401 VCC.n124 VCC.n123 10.6151
R402 VCC.n123 VCC.n120 10.6151
R403 VCC.n120 VCC.n119 10.6151
R404 VCC.n119 VCC.n116 10.6151
R405 VCC.n116 VCC.n115 10.6151
R406 VCC.n115 VCC.n112 10.6151
R407 VCC.n112 VCC.n111 10.6151
R408 VCC.n111 VCC.n108 10.6151
R409 VCC.n108 VCC.n107 10.6151
R410 VCC.n107 VCC.n104 10.6151
R411 VCC.n104 VCC.n103 10.6151
R412 VCC.n103 VCC.n100 10.6151
R413 VCC.n100 VCC.n99 10.6151
R414 VCC.n99 VCC.n96 10.6151
R415 VCC.n96 VCC.n95 10.6151
R416 VCC.n95 VCC.n92 10.6151
R417 VCC.n92 VCC.n91 10.6151
R418 VCC.n91 VCC.n88 10.6151
R419 VCC.n88 VCC.n87 10.6151
R420 VCC.n87 VCC.n84 10.6151
R421 VCC.n84 VCC.n83 10.6151
R422 VCC.n83 VCC.n80 10.6151
R423 VCC.n80 VCC.n79 10.6151
R424 VCC.n79 VCC.n76 10.6151
R425 VCC.n76 VCC.n75 10.6151
R426 VCC.n75 VCC.n72 10.6151
R427 VCC.n72 VCC.n71 10.6151
R428 VCC.n71 VCC.n68 10.6151
R429 VCC.n68 VCC.n67 10.6151
R430 VCC.n67 VCC.n64 10.6151
R431 VCC.n64 VCC.n63 10.6151
R432 VCC.n63 VCC.n60 10.6151
R433 VCC.n60 VCC.n59 10.6151
R434 VCC.n59 VCC.n56 10.6151
R435 VCC.n56 VCC.n31 10.6151
R436 VCC.n286 VCC.n0 9.3005
R437 VCC.n285 VCC.n284 9.3005
R438 VCC.n283 VCC.n6 9.3005
R439 VCC.n282 VCC.n281 9.3005
R440 VCC.n280 VCC.n7 9.3005
R441 VCC.n141 VCC.n30 9.3005
R442 VCC.n143 VCC.n142 9.3005
R443 VCC.n20 VCC.n19 9.3005
R444 VCC.n158 VCC.n157 9.3005
R445 VCC.n159 VCC.n18 9.3005
R446 VCC.n161 VCC.n160 9.3005
R447 VCC.n15 VCC.n14 9.3005
R448 VCC.n170 VCC.n169 9.3005
R449 VCC.n171 VCC.n13 9.3005
R450 VCC.n276 VCC.n275 9.3005
R451 VCC.n140 VCC.n139 9.3005
R452 VCC.n27 VCC.n26 9.3005
R453 VCC.n149 VCC.n148 9.3005
R454 VCC.n150 VCC.n25 9.3005
R455 VCC.n152 VCC.n151 9.3005
R456 VCC.n2 VCC.n1 9.3005
R457 VCC.n288 VCC.n287 9.3005
R458 VCC.n155 VCC.t8 8.89563
R459 VCC.n163 VCC.t9 8.89563
R460 VCC.n146 VCC.t5 8.30262
R461 VCC.n165 VCC.t1 8.30262
R462 VCC.n194 VCC.n190 5.62001
R463 VCC.n131 VCC.n130 5.62001
R464 VCC.n195 VCC.n194 4.99562
R465 VCC.n132 VCC.n131 4.99562
R466 VCC.n284 VCC.n0 0.152939
R467 VCC.n284 VCC.n283 0.152939
R468 VCC.n283 VCC.n282 0.152939
R469 VCC.n282 VCC.n7 0.152939
R470 VCC.n141 VCC.n140 0.152939
R471 VCC.n142 VCC.n141 0.152939
R472 VCC.n142 VCC.n19 0.152939
R473 VCC.n158 VCC.n19 0.152939
R474 VCC.n159 VCC.n158 0.152939
R475 VCC.n160 VCC.n159 0.152939
R476 VCC.n160 VCC.n14 0.152939
R477 VCC.n170 VCC.n14 0.152939
R478 VCC.n171 VCC.n170 0.152939
R479 VCC.n275 VCC.n171 0.152939
R480 VCC.n149 VCC.n26 0.152939
R481 VCC.n150 VCC.n149 0.152939
R482 VCC.n151 VCC.n150 0.152939
R483 VCC.n151 VCC.n1 0.152939
R484 VCC.n288 VCC.n1 0.13922
R485 VCC VCC.n0 0.0767195
R486 VCC VCC.n288 0.063
R487 VGN.n0 VGN.t0 150.111
R488 VGN.n0 VGN.t1 149.555
R489 VGN VGN.n0 6.84834
R490 VIN.n64 VIN.n63 756.745
R491 VIN.n129 VIN.n128 756.745
R492 VIN.n23 VIN.n22 585
R493 VIN.n25 VIN.n24 585
R494 VIN.n18 VIN.n17 585
R495 VIN.n31 VIN.n30 585
R496 VIN.n33 VIN.n32 585
R497 VIN.n14 VIN.n13 585
R498 VIN.n39 VIN.n38 585
R499 VIN.n41 VIN.n40 585
R500 VIN.n10 VIN.n9 585
R501 VIN.n47 VIN.n46 585
R502 VIN.n49 VIN.n48 585
R503 VIN.n6 VIN.n5 585
R504 VIN.n55 VIN.n54 585
R505 VIN.n57 VIN.n56 585
R506 VIN.n2 VIN.n1 585
R507 VIN.n63 VIN.n62 585
R508 VIN.n88 VIN.n87 585
R509 VIN.n90 VIN.n89 585
R510 VIN.n83 VIN.n82 585
R511 VIN.n96 VIN.n95 585
R512 VIN.n98 VIN.n97 585
R513 VIN.n79 VIN.n78 585
R514 VIN.n104 VIN.n103 585
R515 VIN.n106 VIN.n105 585
R516 VIN.n75 VIN.n74 585
R517 VIN.n112 VIN.n111 585
R518 VIN.n114 VIN.n113 585
R519 VIN.n71 VIN.n70 585
R520 VIN.n120 VIN.n119 585
R521 VIN.n122 VIN.n121 585
R522 VIN.n67 VIN.n66 585
R523 VIN.n128 VIN.n127 585
R524 VIN.n21 VIN.t1 327.466
R525 VIN.n86 VIN.t0 327.466
R526 VIN.n179 VIN.n131 289.615
R527 VIN.n232 VIN.n184 289.615
R528 VIN.n180 VIN.n179 185
R529 VIN.n178 VIN.n177 185
R530 VIN.n135 VIN.n134 185
R531 VIN.n172 VIN.n171 185
R532 VIN.n170 VIN.n137 185
R533 VIN.n169 VIN.n168 185
R534 VIN.n140 VIN.n138 185
R535 VIN.n163 VIN.n162 185
R536 VIN.n161 VIN.n160 185
R537 VIN.n144 VIN.n143 185
R538 VIN.n155 VIN.n154 185
R539 VIN.n153 VIN.n152 185
R540 VIN.n148 VIN.n147 185
R541 VIN.n233 VIN.n232 185
R542 VIN.n231 VIN.n230 185
R543 VIN.n188 VIN.n187 185
R544 VIN.n225 VIN.n224 185
R545 VIN.n223 VIN.n190 185
R546 VIN.n222 VIN.n221 185
R547 VIN.n193 VIN.n191 185
R548 VIN.n216 VIN.n215 185
R549 VIN.n214 VIN.n213 185
R550 VIN.n197 VIN.n196 185
R551 VIN.n208 VIN.n207 185
R552 VIN.n206 VIN.n205 185
R553 VIN.n201 VIN.n200 185
R554 VIN.n24 VIN.n23 171.744
R555 VIN.n24 VIN.n17 171.744
R556 VIN.n31 VIN.n17 171.744
R557 VIN.n32 VIN.n31 171.744
R558 VIN.n32 VIN.n13 171.744
R559 VIN.n39 VIN.n13 171.744
R560 VIN.n40 VIN.n39 171.744
R561 VIN.n40 VIN.n9 171.744
R562 VIN.n47 VIN.n9 171.744
R563 VIN.n48 VIN.n47 171.744
R564 VIN.n48 VIN.n5 171.744
R565 VIN.n55 VIN.n5 171.744
R566 VIN.n56 VIN.n55 171.744
R567 VIN.n56 VIN.n1 171.744
R568 VIN.n63 VIN.n1 171.744
R569 VIN.n89 VIN.n88 171.744
R570 VIN.n89 VIN.n82 171.744
R571 VIN.n96 VIN.n82 171.744
R572 VIN.n97 VIN.n96 171.744
R573 VIN.n97 VIN.n78 171.744
R574 VIN.n104 VIN.n78 171.744
R575 VIN.n105 VIN.n104 171.744
R576 VIN.n105 VIN.n74 171.744
R577 VIN.n112 VIN.n74 171.744
R578 VIN.n113 VIN.n112 171.744
R579 VIN.n113 VIN.n70 171.744
R580 VIN.n120 VIN.n70 171.744
R581 VIN.n121 VIN.n120 171.744
R582 VIN.n121 VIN.n66 171.744
R583 VIN.n128 VIN.n66 171.744
R584 VIN.n149 VIN.t2 149.524
R585 VIN.n202 VIN.t3 149.524
R586 VIN.n179 VIN.n178 104.615
R587 VIN.n178 VIN.n134 104.615
R588 VIN.n171 VIN.n134 104.615
R589 VIN.n171 VIN.n170 104.615
R590 VIN.n170 VIN.n169 104.615
R591 VIN.n169 VIN.n138 104.615
R592 VIN.n162 VIN.n138 104.615
R593 VIN.n162 VIN.n161 104.615
R594 VIN.n161 VIN.n143 104.615
R595 VIN.n154 VIN.n143 104.615
R596 VIN.n154 VIN.n153 104.615
R597 VIN.n153 VIN.n147 104.615
R598 VIN.n232 VIN.n231 104.615
R599 VIN.n231 VIN.n187 104.615
R600 VIN.n224 VIN.n187 104.615
R601 VIN.n224 VIN.n223 104.615
R602 VIN.n223 VIN.n222 104.615
R603 VIN.n222 VIN.n191 104.615
R604 VIN.n215 VIN.n191 104.615
R605 VIN.n215 VIN.n214 104.615
R606 VIN.n214 VIN.n196 104.615
R607 VIN.n207 VIN.n196 104.615
R608 VIN.n207 VIN.n206 104.615
R609 VIN.n206 VIN.n200 104.615
R610 VIN.n23 VIN.t1 85.8723
R611 VIN.n88 VIN.t0 85.8723
R612 VIN.t2 VIN.n147 52.3082
R613 VIN.t3 VIN.n200 52.3082
R614 VIN.n237 VIN.n183 37.0298
R615 VIN.n237 VIN.n236 34.9005
R616 VIN.n130 VIN.n64 34.5342
R617 VIN.n130 VIN.n129 33.9308
R618 VIN.n22 VIN.n21 16.3895
R619 VIN.n87 VIN.n86 16.3895
R620 VIN.n172 VIN.n137 13.1884
R621 VIN.n225 VIN.n190 13.1884
R622 VIN.n173 VIN.n135 12.8005
R623 VIN.n168 VIN.n139 12.8005
R624 VIN.n226 VIN.n188 12.8005
R625 VIN.n221 VIN.n192 12.8005
R626 VIN.n25 VIN.n20 12.8005
R627 VIN.n90 VIN.n85 12.8005
R628 VIN VIN.n130 12.132
R629 VIN.n177 VIN.n176 12.0247
R630 VIN.n167 VIN.n140 12.0247
R631 VIN.n230 VIN.n229 12.0247
R632 VIN.n220 VIN.n193 12.0247
R633 VIN.n26 VIN.n18 12.0247
R634 VIN.n62 VIN.n0 12.0247
R635 VIN.n91 VIN.n83 12.0247
R636 VIN.n127 VIN.n65 12.0247
R637 VIN.n180 VIN.n133 11.249
R638 VIN.n164 VIN.n163 11.249
R639 VIN.n233 VIN.n186 11.249
R640 VIN.n217 VIN.n216 11.249
R641 VIN.n30 VIN.n29 11.249
R642 VIN.n61 VIN.n2 11.249
R643 VIN.n95 VIN.n94 11.249
R644 VIN.n126 VIN.n67 11.249
R645 VIN.n181 VIN.n131 10.4732
R646 VIN.n160 VIN.n142 10.4732
R647 VIN.n234 VIN.n184 10.4732
R648 VIN.n213 VIN.n195 10.4732
R649 VIN.n33 VIN.n16 10.4732
R650 VIN.n58 VIN.n57 10.4732
R651 VIN.n98 VIN.n81 10.4732
R652 VIN.n123 VIN.n122 10.4732
R653 VIN.n149 VIN.n148 10.2747
R654 VIN.n202 VIN.n201 10.2747
R655 VIN.n159 VIN.n144 9.69747
R656 VIN.n212 VIN.n197 9.69747
R657 VIN.n34 VIN.n14 9.69747
R658 VIN.n54 VIN.n4 9.69747
R659 VIN.n99 VIN.n79 9.69747
R660 VIN.n119 VIN.n69 9.69747
R661 VIN.n183 VIN.n182 9.45567
R662 VIN.n236 VIN.n235 9.45567
R663 VIN.n60 VIN.n0 9.45567
R664 VIN.n125 VIN.n65 9.45567
R665 VIN.n151 VIN.n150 9.3005
R666 VIN.n146 VIN.n145 9.3005
R667 VIN.n157 VIN.n156 9.3005
R668 VIN.n159 VIN.n158 9.3005
R669 VIN.n142 VIN.n141 9.3005
R670 VIN.n165 VIN.n164 9.3005
R671 VIN.n167 VIN.n166 9.3005
R672 VIN.n139 VIN.n136 9.3005
R673 VIN.n182 VIN.n181 9.3005
R674 VIN.n133 VIN.n132 9.3005
R675 VIN.n176 VIN.n175 9.3005
R676 VIN.n174 VIN.n173 9.3005
R677 VIN.n204 VIN.n203 9.3005
R678 VIN.n199 VIN.n198 9.3005
R679 VIN.n210 VIN.n209 9.3005
R680 VIN.n212 VIN.n211 9.3005
R681 VIN.n195 VIN.n194 9.3005
R682 VIN.n218 VIN.n217 9.3005
R683 VIN.n220 VIN.n219 9.3005
R684 VIN.n192 VIN.n189 9.3005
R685 VIN.n235 VIN.n234 9.3005
R686 VIN.n186 VIN.n185 9.3005
R687 VIN.n229 VIN.n228 9.3005
R688 VIN.n227 VIN.n226 9.3005
R689 VIN.n20 VIN.n19 9.3005
R690 VIN.n27 VIN.n26 9.3005
R691 VIN.n29 VIN.n28 9.3005
R692 VIN.n16 VIN.n15 9.3005
R693 VIN.n35 VIN.n34 9.3005
R694 VIN.n37 VIN.n36 9.3005
R695 VIN.n12 VIN.n11 9.3005
R696 VIN.n43 VIN.n42 9.3005
R697 VIN.n45 VIN.n44 9.3005
R698 VIN.n8 VIN.n7 9.3005
R699 VIN.n51 VIN.n50 9.3005
R700 VIN.n53 VIN.n52 9.3005
R701 VIN.n4 VIN.n3 9.3005
R702 VIN.n59 VIN.n58 9.3005
R703 VIN.n61 VIN.n60 9.3005
R704 VIN.n110 VIN.n109 9.3005
R705 VIN.n73 VIN.n72 9.3005
R706 VIN.n116 VIN.n115 9.3005
R707 VIN.n118 VIN.n117 9.3005
R708 VIN.n69 VIN.n68 9.3005
R709 VIN.n124 VIN.n123 9.3005
R710 VIN.n126 VIN.n125 9.3005
R711 VIN.n77 VIN.n76 9.3005
R712 VIN.n102 VIN.n101 9.3005
R713 VIN.n100 VIN.n99 9.3005
R714 VIN.n81 VIN.n80 9.3005
R715 VIN.n94 VIN.n93 9.3005
R716 VIN.n92 VIN.n91 9.3005
R717 VIN.n85 VIN.n84 9.3005
R718 VIN.n108 VIN.n107 9.3005
R719 VIN.n156 VIN.n155 8.92171
R720 VIN.n209 VIN.n208 8.92171
R721 VIN.n38 VIN.n37 8.92171
R722 VIN.n53 VIN.n6 8.92171
R723 VIN.n103 VIN.n102 8.92171
R724 VIN.n118 VIN.n71 8.92171
R725 VIN.n152 VIN.n146 8.14595
R726 VIN.n205 VIN.n199 8.14595
R727 VIN.n41 VIN.n12 8.14595
R728 VIN.n50 VIN.n49 8.14595
R729 VIN.n106 VIN.n77 8.14595
R730 VIN.n115 VIN.n114 8.14595
R731 VIN.n151 VIN.n148 7.3702
R732 VIN.n204 VIN.n201 7.3702
R733 VIN.n42 VIN.n10 7.3702
R734 VIN.n46 VIN.n8 7.3702
R735 VIN.n107 VIN.n75 7.3702
R736 VIN.n111 VIN.n73 7.3702
R737 VIN.n45 VIN.n10 6.59444
R738 VIN.n46 VIN.n45 6.59444
R739 VIN.n110 VIN.n75 6.59444
R740 VIN.n111 VIN.n110 6.59444
R741 VIN.n152 VIN.n151 5.81868
R742 VIN.n205 VIN.n204 5.81868
R743 VIN.n42 VIN.n41 5.81868
R744 VIN.n49 VIN.n8 5.81868
R745 VIN.n107 VIN.n106 5.81868
R746 VIN.n114 VIN.n73 5.81868
R747 VIN.n155 VIN.n146 5.04292
R748 VIN.n208 VIN.n199 5.04292
R749 VIN.n38 VIN.n12 5.04292
R750 VIN.n50 VIN.n6 5.04292
R751 VIN.n103 VIN.n77 5.04292
R752 VIN.n115 VIN.n71 5.04292
R753 VIN.n156 VIN.n144 4.26717
R754 VIN.n209 VIN.n197 4.26717
R755 VIN.n37 VIN.n14 4.26717
R756 VIN.n54 VIN.n53 4.26717
R757 VIN.n102 VIN.n79 4.26717
R758 VIN.n119 VIN.n118 4.26717
R759 VIN.n21 VIN.n19 3.70982
R760 VIN.n86 VIN.n84 3.70982
R761 VIN.n183 VIN.n131 3.49141
R762 VIN.n160 VIN.n159 3.49141
R763 VIN.n236 VIN.n184 3.49141
R764 VIN.n213 VIN.n212 3.49141
R765 VIN.n34 VIN.n33 3.49141
R766 VIN.n57 VIN.n4 3.49141
R767 VIN.n99 VIN.n98 3.49141
R768 VIN.n122 VIN.n69 3.49141
R769 VIN.n150 VIN.n149 2.84303
R770 VIN.n203 VIN.n202 2.84303
R771 VIN.n181 VIN.n180 2.71565
R772 VIN.n163 VIN.n142 2.71565
R773 VIN.n234 VIN.n233 2.71565
R774 VIN.n216 VIN.n195 2.71565
R775 VIN.n30 VIN.n16 2.71565
R776 VIN.n58 VIN.n2 2.71565
R777 VIN.n95 VIN.n81 2.71565
R778 VIN.n123 VIN.n67 2.71565
R779 VIN.n177 VIN.n133 1.93989
R780 VIN.n164 VIN.n140 1.93989
R781 VIN.n230 VIN.n186 1.93989
R782 VIN.n217 VIN.n193 1.93989
R783 VIN.n29 VIN.n18 1.93989
R784 VIN.n62 VIN.n61 1.93989
R785 VIN.n94 VIN.n83 1.93989
R786 VIN.n127 VIN.n126 1.93989
R787 VIN.n176 VIN.n135 1.16414
R788 VIN.n168 VIN.n167 1.16414
R789 VIN.n229 VIN.n188 1.16414
R790 VIN.n221 VIN.n220 1.16414
R791 VIN.n26 VIN.n25 1.16414
R792 VIN.n64 VIN.n0 1.16414
R793 VIN.n91 VIN.n90 1.16414
R794 VIN.n129 VIN.n65 1.16414
R795 VIN.n173 VIN.n172 0.388379
R796 VIN.n139 VIN.n137 0.388379
R797 VIN.n226 VIN.n225 0.388379
R798 VIN.n192 VIN.n190 0.388379
R799 VIN.n22 VIN.n20 0.388379
R800 VIN.n87 VIN.n85 0.388379
R801 VIN.n182 VIN.n132 0.155672
R802 VIN.n175 VIN.n132 0.155672
R803 VIN.n175 VIN.n174 0.155672
R804 VIN.n174 VIN.n136 0.155672
R805 VIN.n166 VIN.n136 0.155672
R806 VIN.n166 VIN.n165 0.155672
R807 VIN.n165 VIN.n141 0.155672
R808 VIN.n158 VIN.n141 0.155672
R809 VIN.n158 VIN.n157 0.155672
R810 VIN.n157 VIN.n145 0.155672
R811 VIN.n150 VIN.n145 0.155672
R812 VIN.n235 VIN.n185 0.155672
R813 VIN.n228 VIN.n185 0.155672
R814 VIN.n228 VIN.n227 0.155672
R815 VIN.n227 VIN.n189 0.155672
R816 VIN.n219 VIN.n189 0.155672
R817 VIN.n219 VIN.n218 0.155672
R818 VIN.n218 VIN.n194 0.155672
R819 VIN.n211 VIN.n194 0.155672
R820 VIN.n211 VIN.n210 0.155672
R821 VIN.n210 VIN.n198 0.155672
R822 VIN.n203 VIN.n198 0.155672
R823 VIN.n27 VIN.n19 0.155672
R824 VIN.n28 VIN.n27 0.155672
R825 VIN.n28 VIN.n15 0.155672
R826 VIN.n35 VIN.n15 0.155672
R827 VIN.n36 VIN.n35 0.155672
R828 VIN.n36 VIN.n11 0.155672
R829 VIN.n43 VIN.n11 0.155672
R830 VIN.n44 VIN.n43 0.155672
R831 VIN.n44 VIN.n7 0.155672
R832 VIN.n51 VIN.n7 0.155672
R833 VIN.n52 VIN.n51 0.155672
R834 VIN.n52 VIN.n3 0.155672
R835 VIN.n59 VIN.n3 0.155672
R836 VIN.n60 VIN.n59 0.155672
R837 VIN.n92 VIN.n84 0.155672
R838 VIN.n93 VIN.n92 0.155672
R839 VIN.n93 VIN.n80 0.155672
R840 VIN.n100 VIN.n80 0.155672
R841 VIN.n101 VIN.n100 0.155672
R842 VIN.n101 VIN.n76 0.155672
R843 VIN.n108 VIN.n76 0.155672
R844 VIN.n109 VIN.n108 0.155672
R845 VIN.n109 VIN.n72 0.155672
R846 VIN.n116 VIN.n72 0.155672
R847 VIN.n117 VIN.n116 0.155672
R848 VIN.n117 VIN.n68 0.155672
R849 VIN.n124 VIN.n68 0.155672
R850 VIN.n125 VIN.n124 0.155672
R851 VIN VIN.n237 0.00481034
R852 VOUT VOUT.n1 77.9438
R853 VOUT VOUT.n0 76.7474
R854 VOUT.n0 VOUT.t0 2.72972
R855 VOUT.n0 VOUT.t1 2.72972
R856 VOUT.n1 VOUT.t2 1.9609
R857 VOUT.n1 VOUT.t3 1.9609
R858 VSS.n176 VSS.n80 610.22
R859 VSS.n104 VSS.n77 610.22
R860 VSS.n351 VSS.n23 610.22
R861 VSS.n353 VSS.n19 610.22
R862 VSS.n81 VSS.n80 585
R863 VSS.n80 VSS.n78 585
R864 VSS.n181 VSS.n180 585
R865 VSS.n182 VSS.n181 585
R866 VSS.n72 VSS.n71 585
R867 VSS.n79 VSS.n72 585
R868 VSS.n192 VSS.n191 585
R869 VSS.n191 VSS.n190 585
R870 VSS.n69 VSS.n68 585
R871 VSS.n68 VSS.n67 585
R872 VSS.n197 VSS.n196 585
R873 VSS.n198 VSS.n197 585
R874 VSS.n60 VSS.n59 585
R875 VSS.n61 VSS.n60 585
R876 VSS.n208 VSS.n207 585
R877 VSS.n207 VSS.n206 585
R878 VSS.n57 VSS.n56 585
R879 VSS.n56 VSS.n54 585
R880 VSS.n213 VSS.n212 585
R881 VSS.n214 VSS.n213 585
R882 VSS.n47 VSS.n46 585
R883 VSS.n55 VSS.n47 585
R884 VSS.n224 VSS.n223 585
R885 VSS.n223 VSS.n222 585
R886 VSS.n44 VSS.n43 585
R887 VSS.n43 VSS.n42 585
R888 VSS.n229 VSS.n228 585
R889 VSS.n230 VSS.n229 585
R890 VSS.n41 VSS.n40 585
R891 VSS.n231 VSS.n41 585
R892 VSS.n234 VSS.n233 585
R893 VSS.n233 VSS.n232 585
R894 VSS.n38 VSS.n37 585
R895 VSS.n37 VSS.n36 585
R896 VSS.n239 VSS.n238 585
R897 VSS.n240 VSS.n239 585
R898 VSS.n34 VSS.n33 585
R899 VSS.n241 VSS.n34 585
R900 VSS.n244 VSS.n243 585
R901 VSS.n243 VSS.n242 585
R902 VSS.n31 VSS.n30 585
R903 VSS.n30 VSS.n29 585
R904 VSS.n249 VSS.n248 585
R905 VSS.n250 VSS.n249 585
R906 VSS.n27 VSS.n26 585
R907 VSS.n251 VSS.n27 585
R908 VSS.n254 VSS.n253 585
R909 VSS.n253 VSS.n252 585
R910 VSS.n24 VSS.n22 585
R911 VSS.n22 VSS.n20 585
R912 VSS.n351 VSS.n350 585
R913 VSS.n352 VSS.n351 585
R914 VSS.n354 VSS.n353 585
R915 VSS.n353 VSS.n352 585
R916 VSS.n18 VSS.n16 585
R917 VSS.n20 VSS.n18 585
R918 VSS.n358 VSS.n15 585
R919 VSS.n252 VSS.n15 585
R920 VSS.n359 VSS.n14 585
R921 VSS.n251 VSS.n14 585
R922 VSS.n360 VSS.n13 585
R923 VSS.n250 VSS.n13 585
R924 VSS.n28 VSS.n11 585
R925 VSS.n29 VSS.n28 585
R926 VSS.n364 VSS.n10 585
R927 VSS.n242 VSS.n10 585
R928 VSS.n365 VSS.n9 585
R929 VSS.n241 VSS.n9 585
R930 VSS.n366 VSS.n8 585
R931 VSS.n240 VSS.n8 585
R932 VSS.n35 VSS.n6 585
R933 VSS.n36 VSS.n35 585
R934 VSS.n370 VSS.n5 585
R935 VSS.n232 VSS.n5 585
R936 VSS.n371 VSS.n4 585
R937 VSS.n231 VSS.n4 585
R938 VSS.n372 VSS.n3 585
R939 VSS.n230 VSS.n3 585
R940 VSS.n49 VSS.n2 585
R941 VSS.n49 VSS.n42 585
R942 VSS.n221 VSS.n220 585
R943 VSS.n222 VSS.n221 585
R944 VSS.n50 VSS.n48 585
R945 VSS.n55 VSS.n48 585
R946 VSS.n216 VSS.n215 585
R947 VSS.n215 VSS.n214 585
R948 VSS.n53 VSS.n52 585
R949 VSS.n54 VSS.n53 585
R950 VSS.n205 VSS.n204 585
R951 VSS.n206 VSS.n205 585
R952 VSS.n63 VSS.n62 585
R953 VSS.n62 VSS.n61 585
R954 VSS.n200 VSS.n199 585
R955 VSS.n199 VSS.n198 585
R956 VSS.n66 VSS.n65 585
R957 VSS.n67 VSS.n66 585
R958 VSS.n189 VSS.n188 585
R959 VSS.n190 VSS.n189 585
R960 VSS.n74 VSS.n73 585
R961 VSS.n79 VSS.n73 585
R962 VSS.n184 VSS.n183 585
R963 VSS.n183 VSS.n182 585
R964 VSS.n77 VSS.n76 585
R965 VSS.n78 VSS.n77 585
R966 VSS.n19 VSS.n17 585
R967 VSS.n286 VSS.n283 585
R968 VSS.n288 VSS.n287 585
R969 VSS.n290 VSS.n280 585
R970 VSS.n292 VSS.n291 585
R971 VSS.n294 VSS.n278 585
R972 VSS.n296 VSS.n295 585
R973 VSS.n297 VSS.n277 585
R974 VSS.n299 VSS.n298 585
R975 VSS.n301 VSS.n275 585
R976 VSS.n303 VSS.n302 585
R977 VSS.n304 VSS.n274 585
R978 VSS.n306 VSS.n305 585
R979 VSS.n308 VSS.n272 585
R980 VSS.n310 VSS.n309 585
R981 VSS.n311 VSS.n271 585
R982 VSS.n313 VSS.n312 585
R983 VSS.n315 VSS.n269 585
R984 VSS.n317 VSS.n316 585
R985 VSS.n318 VSS.n268 585
R986 VSS.n320 VSS.n319 585
R987 VSS.n322 VSS.n266 585
R988 VSS.n324 VSS.n323 585
R989 VSS.n325 VSS.n265 585
R990 VSS.n327 VSS.n326 585
R991 VSS.n329 VSS.n263 585
R992 VSS.n331 VSS.n330 585
R993 VSS.n332 VSS.n262 585
R994 VSS.n334 VSS.n333 585
R995 VSS.n336 VSS.n260 585
R996 VSS.n338 VSS.n337 585
R997 VSS.n339 VSS.n259 585
R998 VSS.n341 VSS.n340 585
R999 VSS.n343 VSS.n258 585
R1000 VSS.n344 VSS.n257 585
R1001 VSS.n347 VSS.n346 585
R1002 VSS.n348 VSS.n23 585
R1003 VSS.n23 VSS.n21 585
R1004 VSS.n177 VSS.n176 585
R1005 VSS.n83 VSS.n82 585
R1006 VSS.n173 VSS.n172 585
R1007 VSS.n174 VSS.n173 585
R1008 VSS.n171 VSS.n101 585
R1009 VSS.n170 VSS.n169 585
R1010 VSS.n168 VSS.n167 585
R1011 VSS.n166 VSS.n165 585
R1012 VSS.n164 VSS.n163 585
R1013 VSS.n162 VSS.n161 585
R1014 VSS.n160 VSS.n159 585
R1015 VSS.n158 VSS.n157 585
R1016 VSS.n156 VSS.n155 585
R1017 VSS.n154 VSS.n153 585
R1018 VSS.n152 VSS.n151 585
R1019 VSS.n150 VSS.n149 585
R1020 VSS.n148 VSS.n147 585
R1021 VSS.n146 VSS.n145 585
R1022 VSS.n144 VSS.n143 585
R1023 VSS.n142 VSS.n141 585
R1024 VSS.n140 VSS.n139 585
R1025 VSS.n138 VSS.n137 585
R1026 VSS.n136 VSS.n135 585
R1027 VSS.n134 VSS.n133 585
R1028 VSS.n132 VSS.n131 585
R1029 VSS.n130 VSS.n129 585
R1030 VSS.n128 VSS.n127 585
R1031 VSS.n126 VSS.n125 585
R1032 VSS.n124 VSS.n123 585
R1033 VSS.n122 VSS.n121 585
R1034 VSS.n120 VSS.n119 585
R1035 VSS.n118 VSS.n117 585
R1036 VSS.n116 VSS.n115 585
R1037 VSS.n114 VSS.n113 585
R1038 VSS.n112 VSS.n111 585
R1039 VSS.n109 VSS.n108 585
R1040 VSS.n107 VSS.n106 585
R1041 VSS.n105 VSS.n104 585
R1042 VSS.n281 VSS.t6 320.971
R1043 VSS.n102 VSS.t2 320.971
R1044 VSS.n281 VSS.t8 297.49
R1045 VSS.n102 VSS.t5 297.49
R1046 VSS.n174 VSS.n78 260.409
R1047 VSS.n352 VSS.n21 260.409
R1048 VSS.n285 VSS.n21 256.663
R1049 VSS.n284 VSS.n21 256.663
R1050 VSS.n293 VSS.n21 256.663
R1051 VSS.n279 VSS.n21 256.663
R1052 VSS.n300 VSS.n21 256.663
R1053 VSS.n276 VSS.n21 256.663
R1054 VSS.n307 VSS.n21 256.663
R1055 VSS.n273 VSS.n21 256.663
R1056 VSS.n314 VSS.n21 256.663
R1057 VSS.n270 VSS.n21 256.663
R1058 VSS.n321 VSS.n21 256.663
R1059 VSS.n267 VSS.n21 256.663
R1060 VSS.n328 VSS.n21 256.663
R1061 VSS.n264 VSS.n21 256.663
R1062 VSS.n335 VSS.n21 256.663
R1063 VSS.n261 VSS.n21 256.663
R1064 VSS.n342 VSS.n21 256.663
R1065 VSS.n345 VSS.n21 256.663
R1066 VSS.n175 VSS.n174 256.663
R1067 VSS.n174 VSS.n84 256.663
R1068 VSS.n174 VSS.n85 256.663
R1069 VSS.n174 VSS.n86 256.663
R1070 VSS.n174 VSS.n87 256.663
R1071 VSS.n174 VSS.n88 256.663
R1072 VSS.n174 VSS.n89 256.663
R1073 VSS.n174 VSS.n90 256.663
R1074 VSS.n174 VSS.n91 256.663
R1075 VSS.n174 VSS.n92 256.663
R1076 VSS.n174 VSS.n93 256.663
R1077 VSS.n174 VSS.n94 256.663
R1078 VSS.n174 VSS.n95 256.663
R1079 VSS.n174 VSS.n96 256.663
R1080 VSS.n174 VSS.n97 256.663
R1081 VSS.n174 VSS.n98 256.663
R1082 VSS.n174 VSS.n99 256.663
R1083 VSS.n174 VSS.n100 256.663
R1084 VSS.n282 VSS.t9 249.587
R1085 VSS.n103 VSS.t4 249.587
R1086 VSS.n181 VSS.n80 240.244
R1087 VSS.n181 VSS.n72 240.244
R1088 VSS.n191 VSS.n72 240.244
R1089 VSS.n191 VSS.n68 240.244
R1090 VSS.n197 VSS.n68 240.244
R1091 VSS.n197 VSS.n60 240.244
R1092 VSS.n207 VSS.n60 240.244
R1093 VSS.n207 VSS.n56 240.244
R1094 VSS.n213 VSS.n56 240.244
R1095 VSS.n213 VSS.n47 240.244
R1096 VSS.n223 VSS.n47 240.244
R1097 VSS.n223 VSS.n43 240.244
R1098 VSS.n229 VSS.n43 240.244
R1099 VSS.n229 VSS.n41 240.244
R1100 VSS.n233 VSS.n41 240.244
R1101 VSS.n233 VSS.n37 240.244
R1102 VSS.n239 VSS.n37 240.244
R1103 VSS.n239 VSS.n34 240.244
R1104 VSS.n243 VSS.n34 240.244
R1105 VSS.n243 VSS.n30 240.244
R1106 VSS.n249 VSS.n30 240.244
R1107 VSS.n249 VSS.n27 240.244
R1108 VSS.n253 VSS.n27 240.244
R1109 VSS.n253 VSS.n22 240.244
R1110 VSS.n351 VSS.n22 240.244
R1111 VSS.n183 VSS.n77 240.244
R1112 VSS.n183 VSS.n73 240.244
R1113 VSS.n189 VSS.n73 240.244
R1114 VSS.n189 VSS.n66 240.244
R1115 VSS.n199 VSS.n66 240.244
R1116 VSS.n199 VSS.n62 240.244
R1117 VSS.n205 VSS.n62 240.244
R1118 VSS.n205 VSS.n53 240.244
R1119 VSS.n215 VSS.n53 240.244
R1120 VSS.n215 VSS.n48 240.244
R1121 VSS.n221 VSS.n48 240.244
R1122 VSS.n221 VSS.n49 240.244
R1123 VSS.n49 VSS.n3 240.244
R1124 VSS.n4 VSS.n3 240.244
R1125 VSS.n5 VSS.n4 240.244
R1126 VSS.n35 VSS.n5 240.244
R1127 VSS.n35 VSS.n8 240.244
R1128 VSS.n9 VSS.n8 240.244
R1129 VSS.n10 VSS.n9 240.244
R1130 VSS.n28 VSS.n10 240.244
R1131 VSS.n28 VSS.n13 240.244
R1132 VSS.n14 VSS.n13 240.244
R1133 VSS.n15 VSS.n14 240.244
R1134 VSS.n18 VSS.n15 240.244
R1135 VSS.n353 VSS.n18 240.244
R1136 VSS.n173 VSS.n83 163.367
R1137 VSS.n173 VSS.n101 163.367
R1138 VSS.n169 VSS.n168 163.367
R1139 VSS.n165 VSS.n164 163.367
R1140 VSS.n161 VSS.n160 163.367
R1141 VSS.n157 VSS.n156 163.367
R1142 VSS.n153 VSS.n152 163.367
R1143 VSS.n149 VSS.n148 163.367
R1144 VSS.n145 VSS.n144 163.367
R1145 VSS.n141 VSS.n140 163.367
R1146 VSS.n137 VSS.n136 163.367
R1147 VSS.n133 VSS.n132 163.367
R1148 VSS.n129 VSS.n128 163.367
R1149 VSS.n125 VSS.n124 163.367
R1150 VSS.n121 VSS.n120 163.367
R1151 VSS.n117 VSS.n116 163.367
R1152 VSS.n113 VSS.n112 163.367
R1153 VSS.n108 VSS.n107 163.367
R1154 VSS.n346 VSS.n23 163.367
R1155 VSS.n344 VSS.n343 163.367
R1156 VSS.n341 VSS.n259 163.367
R1157 VSS.n337 VSS.n336 163.367
R1158 VSS.n334 VSS.n262 163.367
R1159 VSS.n330 VSS.n329 163.367
R1160 VSS.n327 VSS.n265 163.367
R1161 VSS.n323 VSS.n322 163.367
R1162 VSS.n320 VSS.n268 163.367
R1163 VSS.n316 VSS.n315 163.367
R1164 VSS.n313 VSS.n271 163.367
R1165 VSS.n309 VSS.n308 163.367
R1166 VSS.n306 VSS.n274 163.367
R1167 VSS.n302 VSS.n301 163.367
R1168 VSS.n299 VSS.n277 163.367
R1169 VSS.n295 VSS.n294 163.367
R1170 VSS.n292 VSS.n280 163.367
R1171 VSS.n287 VSS.n286 163.367
R1172 VSS.n182 VSS.n79 149.661
R1173 VSS.n252 VSS.n20 149.661
R1174 VSS.n182 VSS.n78 149.661
R1175 VSS.n190 VSS.n67 149.661
R1176 VSS.n198 VSS.n67 149.661
R1177 VSS.n198 VSS.n61 149.661
R1178 VSS.n206 VSS.n61 149.661
R1179 VSS.n206 VSS.n54 149.661
R1180 VSS.n214 VSS.n54 149.661
R1181 VSS.n214 VSS.n55 149.661
R1182 VSS.n222 VSS.n42 149.661
R1183 VSS.n230 VSS.n42 149.661
R1184 VSS.n231 VSS.n230 149.661
R1185 VSS.n232 VSS.n36 149.661
R1186 VSS.n240 VSS.n36 149.661
R1187 VSS.n241 VSS.n240 149.661
R1188 VSS.n242 VSS.n241 149.661
R1189 VSS.n242 VSS.n29 149.661
R1190 VSS.n250 VSS.n29 149.661
R1191 VSS.n251 VSS.n250 149.661
R1192 VSS.n352 VSS.n20 149.661
R1193 VSS.n222 VSS.t0 145.171
R1194 VSS.t1 VSS.n231 145.171
R1195 VSS.n79 VSS.t3 136.19
R1196 VSS.n252 VSS.t7 136.19
R1197 VSS.n176 VSS.n175 71.676
R1198 VSS.n101 VSS.n84 71.676
R1199 VSS.n168 VSS.n85 71.676
R1200 VSS.n164 VSS.n86 71.676
R1201 VSS.n160 VSS.n87 71.676
R1202 VSS.n156 VSS.n88 71.676
R1203 VSS.n152 VSS.n89 71.676
R1204 VSS.n148 VSS.n90 71.676
R1205 VSS.n144 VSS.n91 71.676
R1206 VSS.n140 VSS.n92 71.676
R1207 VSS.n136 VSS.n93 71.676
R1208 VSS.n132 VSS.n94 71.676
R1209 VSS.n128 VSS.n95 71.676
R1210 VSS.n124 VSS.n96 71.676
R1211 VSS.n120 VSS.n97 71.676
R1212 VSS.n116 VSS.n98 71.676
R1213 VSS.n112 VSS.n99 71.676
R1214 VSS.n107 VSS.n100 71.676
R1215 VSS.n345 VSS.n344 71.676
R1216 VSS.n342 VSS.n341 71.676
R1217 VSS.n337 VSS.n261 71.676
R1218 VSS.n335 VSS.n334 71.676
R1219 VSS.n330 VSS.n264 71.676
R1220 VSS.n328 VSS.n327 71.676
R1221 VSS.n323 VSS.n267 71.676
R1222 VSS.n321 VSS.n320 71.676
R1223 VSS.n316 VSS.n270 71.676
R1224 VSS.n314 VSS.n313 71.676
R1225 VSS.n309 VSS.n273 71.676
R1226 VSS.n307 VSS.n306 71.676
R1227 VSS.n302 VSS.n276 71.676
R1228 VSS.n300 VSS.n299 71.676
R1229 VSS.n295 VSS.n279 71.676
R1230 VSS.n293 VSS.n292 71.676
R1231 VSS.n287 VSS.n284 71.676
R1232 VSS.n285 VSS.n19 71.676
R1233 VSS.n286 VSS.n285 71.676
R1234 VSS.n284 VSS.n280 71.676
R1235 VSS.n294 VSS.n293 71.676
R1236 VSS.n279 VSS.n277 71.676
R1237 VSS.n301 VSS.n300 71.676
R1238 VSS.n276 VSS.n274 71.676
R1239 VSS.n308 VSS.n307 71.676
R1240 VSS.n273 VSS.n271 71.676
R1241 VSS.n315 VSS.n314 71.676
R1242 VSS.n270 VSS.n268 71.676
R1243 VSS.n322 VSS.n321 71.676
R1244 VSS.n267 VSS.n265 71.676
R1245 VSS.n329 VSS.n328 71.676
R1246 VSS.n264 VSS.n262 71.676
R1247 VSS.n336 VSS.n335 71.676
R1248 VSS.n261 VSS.n259 71.676
R1249 VSS.n343 VSS.n342 71.676
R1250 VSS.n346 VSS.n345 71.676
R1251 VSS.n175 VSS.n83 71.676
R1252 VSS.n169 VSS.n84 71.676
R1253 VSS.n165 VSS.n85 71.676
R1254 VSS.n161 VSS.n86 71.676
R1255 VSS.n157 VSS.n87 71.676
R1256 VSS.n153 VSS.n88 71.676
R1257 VSS.n149 VSS.n89 71.676
R1258 VSS.n145 VSS.n90 71.676
R1259 VSS.n141 VSS.n91 71.676
R1260 VSS.n137 VSS.n92 71.676
R1261 VSS.n133 VSS.n93 71.676
R1262 VSS.n129 VSS.n94 71.676
R1263 VSS.n125 VSS.n95 71.676
R1264 VSS.n121 VSS.n96 71.676
R1265 VSS.n117 VSS.n97 71.676
R1266 VSS.n113 VSS.n98 71.676
R1267 VSS.n108 VSS.n99 71.676
R1268 VSS.n104 VSS.n100 71.676
R1269 VSS.n282 VSS.n281 47.9035
R1270 VSS.n103 VSS.n102 47.9035
R1271 VSS.n289 VSS.n282 34.3278
R1272 VSS.n110 VSS.n103 34.3278
R1273 VSS.n349 VSS.n348 28.4535
R1274 VSS.n355 VSS.n17 28.4535
R1275 VSS.n178 VSS.n177 28.4535
R1276 VSS.n105 VSS.n75 28.4535
R1277 VSS.n180 VSS.n81 19.3944
R1278 VSS.n180 VSS.n71 19.3944
R1279 VSS.n192 VSS.n71 19.3944
R1280 VSS.n192 VSS.n69 19.3944
R1281 VSS.n196 VSS.n69 19.3944
R1282 VSS.n196 VSS.n59 19.3944
R1283 VSS.n208 VSS.n59 19.3944
R1284 VSS.n208 VSS.n57 19.3944
R1285 VSS.n212 VSS.n57 19.3944
R1286 VSS.n212 VSS.n46 19.3944
R1287 VSS.n224 VSS.n46 19.3944
R1288 VSS.n224 VSS.n44 19.3944
R1289 VSS.n228 VSS.n44 19.3944
R1290 VSS.n228 VSS.n40 19.3944
R1291 VSS.n234 VSS.n40 19.3944
R1292 VSS.n234 VSS.n38 19.3944
R1293 VSS.n238 VSS.n38 19.3944
R1294 VSS.n238 VSS.n33 19.3944
R1295 VSS.n244 VSS.n33 19.3944
R1296 VSS.n244 VSS.n31 19.3944
R1297 VSS.n248 VSS.n31 19.3944
R1298 VSS.n248 VSS.n26 19.3944
R1299 VSS.n254 VSS.n26 19.3944
R1300 VSS.n254 VSS.n24 19.3944
R1301 VSS.n350 VSS.n24 19.3944
R1302 VSS.n184 VSS.n76 19.3944
R1303 VSS.n184 VSS.n74 19.3944
R1304 VSS.n188 VSS.n74 19.3944
R1305 VSS.n188 VSS.n65 19.3944
R1306 VSS.n200 VSS.n65 19.3944
R1307 VSS.n200 VSS.n63 19.3944
R1308 VSS.n204 VSS.n63 19.3944
R1309 VSS.n204 VSS.n52 19.3944
R1310 VSS.n216 VSS.n52 19.3944
R1311 VSS.n216 VSS.n50 19.3944
R1312 VSS.n220 VSS.n50 19.3944
R1313 VSS.n220 VSS.n2 19.3944
R1314 VSS.n372 VSS.n2 19.3944
R1315 VSS.n372 VSS.n371 19.3944
R1316 VSS.n371 VSS.n370 19.3944
R1317 VSS.n370 VSS.n6 19.3944
R1318 VSS.n366 VSS.n6 19.3944
R1319 VSS.n366 VSS.n365 19.3944
R1320 VSS.n365 VSS.n364 19.3944
R1321 VSS.n364 VSS.n11 19.3944
R1322 VSS.n360 VSS.n11 19.3944
R1323 VSS.n360 VSS.n359 19.3944
R1324 VSS.n359 VSS.n358 19.3944
R1325 VSS.n358 VSS.n16 19.3944
R1326 VSS.n354 VSS.n16 19.3944
R1327 VSS.n190 VSS.t3 13.4699
R1328 VSS.t7 VSS.n251 13.4699
R1329 VSS.n348 VSS.n347 10.6151
R1330 VSS.n347 VSS.n257 10.6151
R1331 VSS.n258 VSS.n257 10.6151
R1332 VSS.n340 VSS.n258 10.6151
R1333 VSS.n340 VSS.n339 10.6151
R1334 VSS.n339 VSS.n338 10.6151
R1335 VSS.n338 VSS.n260 10.6151
R1336 VSS.n333 VSS.n260 10.6151
R1337 VSS.n333 VSS.n332 10.6151
R1338 VSS.n332 VSS.n331 10.6151
R1339 VSS.n331 VSS.n263 10.6151
R1340 VSS.n326 VSS.n263 10.6151
R1341 VSS.n326 VSS.n325 10.6151
R1342 VSS.n325 VSS.n324 10.6151
R1343 VSS.n324 VSS.n266 10.6151
R1344 VSS.n319 VSS.n266 10.6151
R1345 VSS.n319 VSS.n318 10.6151
R1346 VSS.n318 VSS.n317 10.6151
R1347 VSS.n317 VSS.n269 10.6151
R1348 VSS.n312 VSS.n269 10.6151
R1349 VSS.n312 VSS.n311 10.6151
R1350 VSS.n311 VSS.n310 10.6151
R1351 VSS.n310 VSS.n272 10.6151
R1352 VSS.n305 VSS.n272 10.6151
R1353 VSS.n305 VSS.n304 10.6151
R1354 VSS.n304 VSS.n303 10.6151
R1355 VSS.n303 VSS.n275 10.6151
R1356 VSS.n298 VSS.n275 10.6151
R1357 VSS.n298 VSS.n297 10.6151
R1358 VSS.n297 VSS.n296 10.6151
R1359 VSS.n296 VSS.n278 10.6151
R1360 VSS.n291 VSS.n278 10.6151
R1361 VSS.n291 VSS.n290 10.6151
R1362 VSS.n288 VSS.n283 10.6151
R1363 VSS.n283 VSS.n17 10.6151
R1364 VSS.n177 VSS.n82 10.6151
R1365 VSS.n172 VSS.n82 10.6151
R1366 VSS.n172 VSS.n171 10.6151
R1367 VSS.n171 VSS.n170 10.6151
R1368 VSS.n170 VSS.n167 10.6151
R1369 VSS.n167 VSS.n166 10.6151
R1370 VSS.n166 VSS.n163 10.6151
R1371 VSS.n163 VSS.n162 10.6151
R1372 VSS.n162 VSS.n159 10.6151
R1373 VSS.n159 VSS.n158 10.6151
R1374 VSS.n158 VSS.n155 10.6151
R1375 VSS.n155 VSS.n154 10.6151
R1376 VSS.n154 VSS.n151 10.6151
R1377 VSS.n151 VSS.n150 10.6151
R1378 VSS.n150 VSS.n147 10.6151
R1379 VSS.n147 VSS.n146 10.6151
R1380 VSS.n146 VSS.n143 10.6151
R1381 VSS.n143 VSS.n142 10.6151
R1382 VSS.n142 VSS.n139 10.6151
R1383 VSS.n139 VSS.n138 10.6151
R1384 VSS.n138 VSS.n135 10.6151
R1385 VSS.n135 VSS.n134 10.6151
R1386 VSS.n134 VSS.n131 10.6151
R1387 VSS.n131 VSS.n130 10.6151
R1388 VSS.n130 VSS.n127 10.6151
R1389 VSS.n127 VSS.n126 10.6151
R1390 VSS.n126 VSS.n123 10.6151
R1391 VSS.n123 VSS.n122 10.6151
R1392 VSS.n122 VSS.n119 10.6151
R1393 VSS.n119 VSS.n118 10.6151
R1394 VSS.n118 VSS.n115 10.6151
R1395 VSS.n115 VSS.n114 10.6151
R1396 VSS.n114 VSS.n111 10.6151
R1397 VSS.n109 VSS.n106 10.6151
R1398 VSS.n106 VSS.n105 10.6151
R1399 VSS.n371 VSS.n0 9.3005
R1400 VSS.n370 VSS.n369 9.3005
R1401 VSS.n368 VSS.n6 9.3005
R1402 VSS.n367 VSS.n366 9.3005
R1403 VSS.n365 VSS.n7 9.3005
R1404 VSS.n364 VSS.n363 9.3005
R1405 VSS.n362 VSS.n11 9.3005
R1406 VSS.n361 VSS.n360 9.3005
R1407 VSS.n359 VSS.n12 9.3005
R1408 VSS.n358 VSS.n357 9.3005
R1409 VSS.n356 VSS.n16 9.3005
R1410 VSS.n355 VSS.n354 9.3005
R1411 VSS.n178 VSS.n81 9.3005
R1412 VSS.n180 VSS.n179 9.3005
R1413 VSS.n71 VSS.n70 9.3005
R1414 VSS.n193 VSS.n192 9.3005
R1415 VSS.n194 VSS.n69 9.3005
R1416 VSS.n196 VSS.n195 9.3005
R1417 VSS.n59 VSS.n58 9.3005
R1418 VSS.n209 VSS.n208 9.3005
R1419 VSS.n210 VSS.n57 9.3005
R1420 VSS.n212 VSS.n211 9.3005
R1421 VSS.n46 VSS.n45 9.3005
R1422 VSS.n225 VSS.n224 9.3005
R1423 VSS.n226 VSS.n44 9.3005
R1424 VSS.n228 VSS.n227 9.3005
R1425 VSS.n40 VSS.n39 9.3005
R1426 VSS.n235 VSS.n234 9.3005
R1427 VSS.n236 VSS.n38 9.3005
R1428 VSS.n238 VSS.n237 9.3005
R1429 VSS.n33 VSS.n32 9.3005
R1430 VSS.n245 VSS.n244 9.3005
R1431 VSS.n246 VSS.n31 9.3005
R1432 VSS.n248 VSS.n247 9.3005
R1433 VSS.n26 VSS.n25 9.3005
R1434 VSS.n255 VSS.n254 9.3005
R1435 VSS.n256 VSS.n24 9.3005
R1436 VSS.n350 VSS.n349 9.3005
R1437 VSS.n185 VSS.n184 9.3005
R1438 VSS.n186 VSS.n74 9.3005
R1439 VSS.n188 VSS.n187 9.3005
R1440 VSS.n65 VSS.n64 9.3005
R1441 VSS.n201 VSS.n200 9.3005
R1442 VSS.n202 VSS.n63 9.3005
R1443 VSS.n204 VSS.n203 9.3005
R1444 VSS.n52 VSS.n51 9.3005
R1445 VSS.n217 VSS.n216 9.3005
R1446 VSS.n218 VSS.n50 9.3005
R1447 VSS.n220 VSS.n219 9.3005
R1448 VSS.n2 VSS.n1 9.3005
R1449 VSS.n76 VSS.n75 9.3005
R1450 VSS VSS.n372 9.3005
R1451 VSS.n290 VSS.n289 9.21026
R1452 VSS.n111 VSS.n110 9.21026
R1453 VSS.n55 VSS.t0 4.4903
R1454 VSS.n232 VSS.t1 4.4903
R1455 VSS.n289 VSS.n288 1.40538
R1456 VSS.n110 VSS.n109 1.40538
R1457 VSS VSS.n0 0.152939
R1458 VSS.n369 VSS.n0 0.152939
R1459 VSS.n369 VSS.n368 0.152939
R1460 VSS.n368 VSS.n367 0.152939
R1461 VSS.n367 VSS.n7 0.152939
R1462 VSS.n363 VSS.n7 0.152939
R1463 VSS.n363 VSS.n362 0.152939
R1464 VSS.n362 VSS.n361 0.152939
R1465 VSS.n361 VSS.n12 0.152939
R1466 VSS.n357 VSS.n12 0.152939
R1467 VSS.n357 VSS.n356 0.152939
R1468 VSS.n356 VSS.n355 0.152939
R1469 VSS.n179 VSS.n178 0.152939
R1470 VSS.n179 VSS.n70 0.152939
R1471 VSS.n193 VSS.n70 0.152939
R1472 VSS.n194 VSS.n193 0.152939
R1473 VSS.n195 VSS.n194 0.152939
R1474 VSS.n195 VSS.n58 0.152939
R1475 VSS.n209 VSS.n58 0.152939
R1476 VSS.n210 VSS.n209 0.152939
R1477 VSS.n211 VSS.n210 0.152939
R1478 VSS.n211 VSS.n45 0.152939
R1479 VSS.n225 VSS.n45 0.152939
R1480 VSS.n226 VSS.n225 0.152939
R1481 VSS.n227 VSS.n226 0.152939
R1482 VSS.n227 VSS.n39 0.152939
R1483 VSS.n235 VSS.n39 0.152939
R1484 VSS.n236 VSS.n235 0.152939
R1485 VSS.n237 VSS.n236 0.152939
R1486 VSS.n237 VSS.n32 0.152939
R1487 VSS.n245 VSS.n32 0.152939
R1488 VSS.n246 VSS.n245 0.152939
R1489 VSS.n247 VSS.n246 0.152939
R1490 VSS.n247 VSS.n25 0.152939
R1491 VSS.n255 VSS.n25 0.152939
R1492 VSS.n256 VSS.n255 0.152939
R1493 VSS.n349 VSS.n256 0.152939
R1494 VSS.n185 VSS.n75 0.152939
R1495 VSS.n186 VSS.n185 0.152939
R1496 VSS.n187 VSS.n186 0.152939
R1497 VSS.n187 VSS.n64 0.152939
R1498 VSS.n201 VSS.n64 0.152939
R1499 VSS.n202 VSS.n201 0.152939
R1500 VSS.n203 VSS.n202 0.152939
R1501 VSS.n203 VSS.n51 0.152939
R1502 VSS.n217 VSS.n51 0.152939
R1503 VSS.n218 VSS.n217 0.152939
R1504 VSS.n219 VSS.n218 0.152939
R1505 VSS.n219 VSS.n1 0.152939
R1506 VSS VSS.n1 0.1255
R1507 VGP.n0 VGP.t1 906.682
R1508 VGP.n0 VGP.t0 906.682
R1509 VGP VGP.n0 161.452
C0 VGP VIN 0.762738f
C1 VCC VGP 0.580019f
C2 VCC VIN 2.21639f
C3 VOUT VGN 1.59386f
C4 VGN VGP 0.002956f
C5 VOUT VGP 0.74915f
C6 VGN VIN 1.78185f
C7 VOUT VIN 4.42483f
C8 VGN VCC 0.024367f
C9 VOUT VCC 0.710361f
C10 VGN VSS 2.34879f
C11 VOUT VSS 2.016706f
C12 VIN VSS 2.827107f
C13 VGP VSS 0.119165f
C14 VCC VSS 16.92188f
C15 VOUT.t0 VSS 0.168131f
C16 VOUT.t1 VSS 0.168131f
C17 VOUT.n0 VSS 1.32675f
C18 VOUT.t2 VSS 0.14258f
C19 VOUT.t3 VSS 0.14258f
C20 VOUT.n1 VSS 1.34595f
C21 VIN.n0 VSS 0.007823f
C22 VIN.n1 VSS 0.017659f
C23 VIN.n2 VSS 0.007911f
C24 VIN.n3 VSS 0.013903f
C25 VIN.n4 VSS 0.007471f
C26 VIN.n5 VSS 0.017659f
C27 VIN.n6 VSS 0.007911f
C28 VIN.n7 VSS 0.013903f
C29 VIN.n8 VSS 0.007471f
C30 VIN.n9 VSS 0.017659f
C31 VIN.n10 VSS 0.007911f
C32 VIN.n11 VSS 0.013903f
C33 VIN.n12 VSS 0.007471f
C34 VIN.n13 VSS 0.017659f
C35 VIN.n14 VSS 0.007911f
C36 VIN.n15 VSS 0.013903f
C37 VIN.n16 VSS 0.007471f
C38 VIN.n17 VSS 0.017659f
C39 VIN.n18 VSS 0.007911f
C40 VIN.n19 VSS 0.692724f
C41 VIN.n20 VSS 0.007471f
C42 VIN.t1 VSS 0.037699f
C43 VIN.n21 VSS 0.085337f
C44 VIN.n22 VSS 0.011234f
C45 VIN.n23 VSS 0.013244f
C46 VIN.n24 VSS 0.017659f
C47 VIN.n25 VSS 0.007911f
C48 VIN.n26 VSS 0.007471f
C49 VIN.n27 VSS 0.013903f
C50 VIN.n28 VSS 0.013903f
C51 VIN.n29 VSS 0.007471f
C52 VIN.n30 VSS 0.007911f
C53 VIN.n31 VSS 0.017659f
C54 VIN.n32 VSS 0.017659f
C55 VIN.n33 VSS 0.007911f
C56 VIN.n34 VSS 0.007471f
C57 VIN.n35 VSS 0.013903f
C58 VIN.n36 VSS 0.013903f
C59 VIN.n37 VSS 0.007471f
C60 VIN.n38 VSS 0.007911f
C61 VIN.n39 VSS 0.017659f
C62 VIN.n40 VSS 0.017659f
C63 VIN.n41 VSS 0.007911f
C64 VIN.n42 VSS 0.007471f
C65 VIN.n43 VSS 0.013903f
C66 VIN.n44 VSS 0.013903f
C67 VIN.n45 VSS 0.007471f
C68 VIN.n46 VSS 0.007911f
C69 VIN.n47 VSS 0.017659f
C70 VIN.n48 VSS 0.017659f
C71 VIN.n49 VSS 0.007911f
C72 VIN.n50 VSS 0.007471f
C73 VIN.n51 VSS 0.013903f
C74 VIN.n52 VSS 0.013903f
C75 VIN.n53 VSS 0.007471f
C76 VIN.n54 VSS 0.007911f
C77 VIN.n55 VSS 0.017659f
C78 VIN.n56 VSS 0.017659f
C79 VIN.n57 VSS 0.007911f
C80 VIN.n58 VSS 0.007471f
C81 VIN.n59 VSS 0.013903f
C82 VIN.n60 VSS 0.034986f
C83 VIN.n61 VSS 0.007471f
C84 VIN.n62 VSS 0.007911f
C85 VIN.n63 VSS 0.038337f
C86 VIN.n64 VSS 0.026326f
C87 VIN.n65 VSS 0.007823f
C88 VIN.n66 VSS 0.017659f
C89 VIN.n67 VSS 0.007911f
C90 VIN.n68 VSS 0.013903f
C91 VIN.n69 VSS 0.007471f
C92 VIN.n70 VSS 0.017659f
C93 VIN.n71 VSS 0.007911f
C94 VIN.n72 VSS 0.013903f
C95 VIN.n73 VSS 0.007471f
C96 VIN.n74 VSS 0.017659f
C97 VIN.n75 VSS 0.007911f
C98 VIN.n76 VSS 0.013903f
C99 VIN.n77 VSS 0.007471f
C100 VIN.n78 VSS 0.017659f
C101 VIN.n79 VSS 0.007911f
C102 VIN.n80 VSS 0.013903f
C103 VIN.n81 VSS 0.007471f
C104 VIN.n82 VSS 0.017659f
C105 VIN.n83 VSS 0.007911f
C106 VIN.n84 VSS 0.692724f
C107 VIN.n85 VSS 0.007471f
C108 VIN.t0 VSS 0.037699f
C109 VIN.n86 VSS 0.085337f
C110 VIN.n87 VSS 0.011234f
C111 VIN.n88 VSS 0.013244f
C112 VIN.n89 VSS 0.017659f
C113 VIN.n90 VSS 0.007911f
C114 VIN.n91 VSS 0.007471f
C115 VIN.n92 VSS 0.013903f
C116 VIN.n93 VSS 0.013903f
C117 VIN.n94 VSS 0.007471f
C118 VIN.n95 VSS 0.007911f
C119 VIN.n96 VSS 0.017659f
C120 VIN.n97 VSS 0.017659f
C121 VIN.n98 VSS 0.007911f
C122 VIN.n99 VSS 0.007471f
C123 VIN.n100 VSS 0.013903f
C124 VIN.n101 VSS 0.013903f
C125 VIN.n102 VSS 0.007471f
C126 VIN.n103 VSS 0.007911f
C127 VIN.n104 VSS 0.017659f
C128 VIN.n105 VSS 0.017659f
C129 VIN.n106 VSS 0.007911f
C130 VIN.n107 VSS 0.007471f
C131 VIN.n108 VSS 0.013903f
C132 VIN.n109 VSS 0.013903f
C133 VIN.n110 VSS 0.007471f
C134 VIN.n111 VSS 0.007911f
C135 VIN.n112 VSS 0.017659f
C136 VIN.n113 VSS 0.017659f
C137 VIN.n114 VSS 0.007911f
C138 VIN.n115 VSS 0.007471f
C139 VIN.n116 VSS 0.013903f
C140 VIN.n117 VSS 0.013903f
C141 VIN.n118 VSS 0.007471f
C142 VIN.n119 VSS 0.007911f
C143 VIN.n120 VSS 0.017659f
C144 VIN.n121 VSS 0.017659f
C145 VIN.n122 VSS 0.007911f
C146 VIN.n123 VSS 0.007471f
C147 VIN.n124 VSS 0.013903f
C148 VIN.n125 VSS 0.034986f
C149 VIN.n126 VSS 0.007471f
C150 VIN.n127 VSS 0.007911f
C151 VIN.n128 VSS 0.038337f
C152 VIN.n129 VSS 0.025531f
C153 VIN.n130 VSS 0.285986f
C154 VIN.n131 VSS 0.01973f
C155 VIN.n132 VSS 0.013903f
C156 VIN.n133 VSS 0.007471f
C157 VIN.n134 VSS 0.017659f
C158 VIN.n135 VSS 0.007911f
C159 VIN.n136 VSS 0.013903f
C160 VIN.n137 VSS 0.007691f
C161 VIN.n138 VSS 0.017659f
C162 VIN.n139 VSS 0.007471f
C163 VIN.n140 VSS 0.007911f
C164 VIN.n141 VSS 0.013903f
C165 VIN.n142 VSS 0.007471f
C166 VIN.n143 VSS 0.017659f
C167 VIN.n144 VSS 0.007911f
C168 VIN.n145 VSS 0.013903f
C169 VIN.n146 VSS 0.007471f
C170 VIN.n147 VSS 0.013244f
C171 VIN.n148 VSS 0.012483f
C172 VIN.t2 VSS 0.029684f
C173 VIN.n149 VSS 0.090103f
C174 VIN.n150 VSS 0.583903f
C175 VIN.n151 VSS 0.007471f
C176 VIN.n152 VSS 0.007911f
C177 VIN.n153 VSS 0.017659f
C178 VIN.n154 VSS 0.017659f
C179 VIN.n155 VSS 0.007911f
C180 VIN.n156 VSS 0.007471f
C181 VIN.n157 VSS 0.013903f
C182 VIN.n158 VSS 0.013903f
C183 VIN.n159 VSS 0.007471f
C184 VIN.n160 VSS 0.007911f
C185 VIN.n161 VSS 0.017659f
C186 VIN.n162 VSS 0.017659f
C187 VIN.n163 VSS 0.007911f
C188 VIN.n164 VSS 0.007471f
C189 VIN.n165 VSS 0.013903f
C190 VIN.n166 VSS 0.013903f
C191 VIN.n167 VSS 0.007471f
C192 VIN.n168 VSS 0.007911f
C193 VIN.n169 VSS 0.017659f
C194 VIN.n170 VSS 0.017659f
C195 VIN.n171 VSS 0.017659f
C196 VIN.n172 VSS 0.007691f
C197 VIN.n173 VSS 0.007471f
C198 VIN.n174 VSS 0.013903f
C199 VIN.n175 VSS 0.013903f
C200 VIN.n176 VSS 0.007471f
C201 VIN.n177 VSS 0.007911f
C202 VIN.n178 VSS 0.017659f
C203 VIN.n179 VSS 0.03856f
C204 VIN.n180 VSS 0.007911f
C205 VIN.n181 VSS 0.007471f
C206 VIN.n182 VSS 0.034796f
C207 VIN.n183 VSS 0.028266f
C208 VIN.n184 VSS 0.01973f
C209 VIN.n185 VSS 0.013903f
C210 VIN.n186 VSS 0.007471f
C211 VIN.n187 VSS 0.017659f
C212 VIN.n188 VSS 0.007911f
C213 VIN.n189 VSS 0.013903f
C214 VIN.n190 VSS 0.007691f
C215 VIN.n191 VSS 0.017659f
C216 VIN.n192 VSS 0.007471f
C217 VIN.n193 VSS 0.007911f
C218 VIN.n194 VSS 0.013903f
C219 VIN.n195 VSS 0.007471f
C220 VIN.n196 VSS 0.017659f
C221 VIN.n197 VSS 0.007911f
C222 VIN.n198 VSS 0.013903f
C223 VIN.n199 VSS 0.007471f
C224 VIN.n200 VSS 0.013244f
C225 VIN.n201 VSS 0.012483f
C226 VIN.t3 VSS 0.029684f
C227 VIN.n202 VSS 0.090103f
C228 VIN.n203 VSS 0.583903f
C229 VIN.n204 VSS 0.007471f
C230 VIN.n205 VSS 0.007911f
C231 VIN.n206 VSS 0.017659f
C232 VIN.n207 VSS 0.017659f
C233 VIN.n208 VSS 0.007911f
C234 VIN.n209 VSS 0.007471f
C235 VIN.n210 VSS 0.013903f
C236 VIN.n211 VSS 0.013903f
C237 VIN.n212 VSS 0.007471f
C238 VIN.n213 VSS 0.007911f
C239 VIN.n214 VSS 0.017659f
C240 VIN.n215 VSS 0.017659f
C241 VIN.n216 VSS 0.007911f
C242 VIN.n217 VSS 0.007471f
C243 VIN.n218 VSS 0.013903f
C244 VIN.n219 VSS 0.013903f
C245 VIN.n220 VSS 0.007471f
C246 VIN.n221 VSS 0.007911f
C247 VIN.n222 VSS 0.017659f
C248 VIN.n223 VSS 0.017659f
C249 VIN.n224 VSS 0.017659f
C250 VIN.n225 VSS 0.007691f
C251 VIN.n226 VSS 0.007471f
C252 VIN.n227 VSS 0.013903f
C253 VIN.n228 VSS 0.013903f
C254 VIN.n229 VSS 0.007471f
C255 VIN.n230 VSS 0.007911f
C256 VIN.n231 VSS 0.017659f
C257 VIN.n232 VSS 0.03856f
C258 VIN.n233 VSS 0.007911f
C259 VIN.n234 VSS 0.007471f
C260 VIN.n235 VSS 0.034796f
C261 VIN.n236 VSS 0.021689f
C262 VIN.n237 VSS 0.216759f
C263 VCC.n0 VSS 0.001596f
C264 VCC.n1 VSS 0.002128f
C265 VCC.n2 VSS 0.001713f
C266 VCC.n3 VSS 0.002128f
C267 VCC.n4 VSS 0.002128f
C268 VCC.n5 VSS 0.002128f
C269 VCC.n6 VSS 0.001713f
C270 VCC.n7 VSS 0.007585f
C271 VCC.n8 VSS 0.002128f
C272 VCC.n9 VSS 0.004364f
C273 VCC.t1 VSS 0.04158f
C274 VCC.n10 VSS 0.164657f
C275 VCC.n11 VSS 0.002128f
C276 VCC.n12 VSS 0.004364f
C277 VCC.n13 VSS 0.001713f
C278 VCC.n14 VSS 0.002128f
C279 VCC.n15 VSS 0.001713f
C280 VCC.n16 VSS 0.002128f
C281 VCC.t9 VSS 0.04158f
C282 VCC.n17 VSS 0.002128f
C283 VCC.n18 VSS 0.001713f
C284 VCC.n19 VSS 0.002128f
C285 VCC.n20 VSS 0.001713f
C286 VCC.n21 VSS 0.002128f
C287 VCC.n22 VSS 0.08316f
C288 VCC.n23 VSS 0.058212f
C289 VCC.t8 VSS 0.04158f
C290 VCC.n24 VSS 0.002128f
C291 VCC.n25 VSS 0.001713f
C292 VCC.n26 VSS 0.007585f
C293 VCC.n27 VSS 0.001422f
C294 VCC.n28 VSS 0.004426f
C295 VCC.t5 VSS 0.04158f
C296 VCC.n29 VSS 0.002128f
C297 VCC.n30 VSS 0.001713f
C298 VCC.n31 VSS 0.00295f
C299 VCC.n32 VSS 0.004364f
C300 VCC.n52 VSS 0.001447f
C301 VCC.n53 VSS 0.001447f
C302 VCC.t6 VSS 0.043163f
C303 VCC.t7 VSS 0.044841f
C304 VCC.t4 VSS 0.036165f
C305 VCC.n54 VSS 0.058123f
C306 VCC.n55 VSS 0.048615f
C307 VCC.n56 VSS 0.001447f
C308 VCC.n57 VSS 0.001447f
C309 VCC.n58 VSS 0.001447f
C310 VCC.n59 VSS 0.001447f
C311 VCC.n60 VSS 0.001447f
C312 VCC.n61 VSS 0.001447f
C313 VCC.n62 VSS 0.001447f
C314 VCC.n63 VSS 0.001447f
C315 VCC.n64 VSS 0.001447f
C316 VCC.n65 VSS 0.001447f
C317 VCC.n66 VSS 0.001447f
C318 VCC.n67 VSS 0.001447f
C319 VCC.n68 VSS 0.001447f
C320 VCC.n69 VSS 0.001447f
C321 VCC.n70 VSS 0.001447f
C322 VCC.n71 VSS 0.001447f
C323 VCC.n72 VSS 0.001447f
C324 VCC.n73 VSS 0.001447f
C325 VCC.n74 VSS 0.001447f
C326 VCC.n75 VSS 0.001447f
C327 VCC.n76 VSS 0.001447f
C328 VCC.n77 VSS 0.001447f
C329 VCC.n78 VSS 0.001447f
C330 VCC.n79 VSS 0.001447f
C331 VCC.n80 VSS 0.001447f
C332 VCC.n81 VSS 0.001447f
C333 VCC.n82 VSS 0.001447f
C334 VCC.n83 VSS 0.001447f
C335 VCC.n84 VSS 0.001447f
C336 VCC.n85 VSS 0.001447f
C337 VCC.n86 VSS 0.001447f
C338 VCC.n87 VSS 0.001447f
C339 VCC.n88 VSS 0.001447f
C340 VCC.n89 VSS 0.001447f
C341 VCC.n90 VSS 0.001447f
C342 VCC.n91 VSS 0.001447f
C343 VCC.n92 VSS 0.001447f
C344 VCC.n93 VSS 0.001447f
C345 VCC.n94 VSS 0.001447f
C346 VCC.n95 VSS 0.001447f
C347 VCC.n96 VSS 0.001447f
C348 VCC.n97 VSS 0.001447f
C349 VCC.n98 VSS 0.001447f
C350 VCC.n99 VSS 0.001447f
C351 VCC.n100 VSS 0.001447f
C352 VCC.n101 VSS 0.001447f
C353 VCC.n102 VSS 0.001447f
C354 VCC.n103 VSS 0.001447f
C355 VCC.n104 VSS 0.001447f
C356 VCC.n105 VSS 0.001447f
C357 VCC.n106 VSS 0.001447f
C358 VCC.n107 VSS 0.001447f
C359 VCC.n108 VSS 0.001447f
C360 VCC.n109 VSS 0.001447f
C361 VCC.n110 VSS 0.001447f
C362 VCC.n111 VSS 0.001447f
C363 VCC.n112 VSS 0.001447f
C364 VCC.n113 VSS 0.001447f
C365 VCC.n114 VSS 0.001447f
C366 VCC.n115 VSS 0.001447f
C367 VCC.n116 VSS 0.001447f
C368 VCC.n117 VSS 0.001447f
C369 VCC.n118 VSS 0.001447f
C370 VCC.n119 VSS 0.001447f
C371 VCC.n120 VSS 0.001447f
C372 VCC.n121 VSS 0.001447f
C373 VCC.n122 VSS 0.001447f
C374 VCC.n123 VSS 0.001447f
C375 VCC.n124 VSS 0.001447f
C376 VCC.n125 VSS 0.001447f
C377 VCC.n126 VSS 0.001447f
C378 VCC.n127 VSS 0.001447f
C379 VCC.n128 VSS 0.001447f
C380 VCC.n129 VSS 0.001447f
C381 VCC.n130 VSS 0.001107f
C382 VCC.n131 VSS 0.002017f
C383 VCC.n132 VSS 0.001064f
C384 VCC.n133 VSS 0.00295f
C385 VCC.n134 VSS 0.004364f
C386 VCC.n136 VSS 0.164657f
C387 VCC.n137 VSS 0.10894f
C388 VCC.n138 VSS 0.004426f
C389 VCC.n139 VSS 0.001422f
C390 VCC.n140 VSS 0.007585f
C391 VCC.n141 VSS 0.002128f
C392 VCC.n142 VSS 0.002128f
C393 VCC.n143 VSS 0.001713f
C394 VCC.n144 VSS 0.002128f
C395 VCC.n145 VSS 0.08316f
C396 VCC.n146 VSS 0.053222f
C397 VCC.n147 VSS 0.002128f
C398 VCC.n148 VSS 0.001713f
C399 VCC.n149 VSS 0.002128f
C400 VCC.n150 VSS 0.002128f
C401 VCC.n151 VSS 0.002128f
C402 VCC.n152 VSS 0.001713f
C403 VCC.n153 VSS 0.002128f
C404 VCC.n154 VSS 0.002128f
C405 VCC.n155 VSS 0.054054f
C406 VCC.n156 VSS 0.002128f
C407 VCC.n157 VSS 0.001713f
C408 VCC.n158 VSS 0.002128f
C409 VCC.n159 VSS 0.002128f
C410 VCC.n160 VSS 0.002128f
C411 VCC.n161 VSS 0.001713f
C412 VCC.n162 VSS 0.002128f
C413 VCC.n163 VSS 0.054054f
C414 VCC.n164 VSS 0.08316f
C415 VCC.n165 VSS 0.053222f
C416 VCC.n166 VSS 0.002128f
C417 VCC.n167 VSS 0.08316f
C418 VCC.n168 VSS 0.002128f
C419 VCC.n169 VSS 0.001713f
C420 VCC.n170 VSS 0.002128f
C421 VCC.n171 VSS 0.002128f
C422 VCC.n172 VSS 0.001447f
C423 VCC.n173 VSS 0.001447f
C424 VCC.n174 VSS 0.001447f
C425 VCC.n175 VSS 0.001447f
C426 VCC.n176 VSS 0.001447f
C427 VCC.n177 VSS 0.001447f
C428 VCC.n178 VSS 0.001447f
C429 VCC.n179 VSS 0.001447f
C430 VCC.n180 VSS 0.001447f
C431 VCC.n181 VSS 0.001447f
C432 VCC.n182 VSS 0.001447f
C433 VCC.n183 VSS 0.001447f
C434 VCC.n184 VSS 0.001447f
C435 VCC.n185 VSS 0.001447f
C436 VCC.n186 VSS 0.001447f
C437 VCC.n187 VSS 0.001447f
C438 VCC.n188 VSS 0.001447f
C439 VCC.n189 VSS 0.001447f
C440 VCC.n190 VSS 0.001107f
C441 VCC.n191 VSS 0.00295f
C442 VCC.t3 VSS 0.043163f
C443 VCC.t2 VSS 0.044841f
C444 VCC.t0 VSS 0.036165f
C445 VCC.n192 VSS 0.058123f
C446 VCC.n193 VSS 0.048615f
C447 VCC.n194 VSS 0.002017f
C448 VCC.n195 VSS 0.001064f
C449 VCC.n196 VSS 0.001447f
C450 VCC.n198 VSS 0.001447f
C451 VCC.n200 VSS 0.001447f
C452 VCC.n201 VSS 0.001447f
C453 VCC.n202 VSS 0.001447f
C454 VCC.n203 VSS 0.001447f
C455 VCC.n204 VSS 0.001447f
C456 VCC.n206 VSS 0.001447f
C457 VCC.n208 VSS 0.001447f
C458 VCC.n209 VSS 0.001447f
C459 VCC.n210 VSS 0.001447f
C460 VCC.n211 VSS 0.001447f
C461 VCC.n212 VSS 0.001447f
C462 VCC.n214 VSS 0.001447f
C463 VCC.n216 VSS 0.001447f
C464 VCC.n217 VSS 0.001447f
C465 VCC.n218 VSS 0.001447f
C466 VCC.n219 VSS 0.001447f
C467 VCC.n220 VSS 0.001447f
C468 VCC.n222 VSS 0.001447f
C469 VCC.n224 VSS 0.001447f
C470 VCC.n225 VSS 0.001447f
C471 VCC.n226 VSS 0.001447f
C472 VCC.n227 VSS 0.001447f
C473 VCC.n228 VSS 0.001447f
C474 VCC.n230 VSS 0.001447f
C475 VCC.n232 VSS 0.001447f
C476 VCC.n233 VSS 0.001447f
C477 VCC.n234 VSS 0.001447f
C478 VCC.n235 VSS 0.001447f
C479 VCC.n236 VSS 0.001447f
C480 VCC.n238 VSS 0.001447f
C481 VCC.n240 VSS 0.001447f
C482 VCC.n241 VSS 0.001447f
C483 VCC.n242 VSS 0.001447f
C484 VCC.n243 VSS 0.001447f
C485 VCC.n244 VSS 0.001447f
C486 VCC.n246 VSS 0.001447f
C487 VCC.n248 VSS 0.001447f
C488 VCC.n249 VSS 0.001447f
C489 VCC.n250 VSS 0.001447f
C490 VCC.n251 VSS 0.001447f
C491 VCC.n252 VSS 0.001447f
C492 VCC.n254 VSS 0.001447f
C493 VCC.n256 VSS 0.001447f
C494 VCC.n257 VSS 0.001447f
C495 VCC.n258 VSS 0.001447f
C496 VCC.n259 VSS 0.001447f
C497 VCC.n260 VSS 0.001447f
C498 VCC.n262 VSS 0.001447f
C499 VCC.n264 VSS 0.001447f
C500 VCC.n265 VSS 0.001447f
C501 VCC.n266 VSS 0.001447f
C502 VCC.n267 VSS 0.001447f
C503 VCC.n268 VSS 0.001447f
C504 VCC.n270 VSS 0.001447f
C505 VCC.n272 VSS 0.001447f
C506 VCC.n273 VSS 0.001447f
C507 VCC.n274 VSS 0.00295f
C508 VCC.n275 VSS 0.007585f
C509 VCC.n276 VSS 0.001422f
C510 VCC.n277 VSS 0.004426f
C511 VCC.n278 VSS 0.10894f
C512 VCC.n279 VSS 0.004426f
C513 VCC.n280 VSS 0.001422f
C514 VCC.n281 VSS 0.001713f
C515 VCC.n282 VSS 0.002128f
C516 VCC.n283 VSS 0.002128f
C517 VCC.n284 VSS 0.002128f
C518 VCC.n285 VSS 0.001713f
C519 VCC.n286 VSS 0.001713f
C520 VCC.n287 VSS 0.001713f
C521 VCC.n288 VSS 0.001947f
.ends

