* NGSPICE file created from diff_pair_sample_0853.ext - technology: sky130A

.subckt diff_pair_sample_0853 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=3.15
X1 VDD1.t6 VP.t1 VTAIL.t15 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=3.15
X2 VTAIL.t5 VN.t0 VDD2.t7 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=3.15
X3 VDD2.t6 VN.t1 VTAIL.t0 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=3.15
X4 VDD1.t5 VP.t2 VTAIL.t8 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X5 B.t11 B.t9 B.t10 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=3.15
X6 VDD2.t5 VN.t2 VTAIL.t6 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=4.2198 ps=22.42 w=10.82 l=3.15
X7 VTAIL.t3 VN.t3 VDD2.t4 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X8 B.t8 B.t6 B.t7 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=3.15
X9 B.t5 B.t3 B.t4 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=3.15
X10 B.t2 B.t0 B.t1 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=0 ps=0 w=10.82 l=3.15
X11 VTAIL.t2 VN.t4 VDD2.t3 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X12 VTAIL.t11 VP.t3 VDD1.t4 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=3.15
X13 VTAIL.t9 VP.t4 VDD1.t3 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=3.15
X14 VTAIL.t14 VP.t5 VDD1.t2 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X15 VTAIL.t4 VN.t5 VDD2.t2 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=4.2198 pd=22.42 as=1.7853 ps=11.15 w=10.82 l=3.15
X16 VDD1.t1 VP.t6 VTAIL.t10 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X17 VDD2.t1 VN.t6 VTAIL.t1 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X18 VDD2.t0 VN.t7 VTAIL.t7 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
X19 VTAIL.t13 VP.t7 VDD1.t0 w_n4450_n3132# sky130_fd_pr__pfet_01v8 ad=1.7853 pd=11.15 as=1.7853 ps=11.15 w=10.82 l=3.15
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n19 VP.t3 116.111
R34 VP.n43 VP.t4 82.7821
R35 VP.n55 VP.t2 82.7821
R36 VP.n4 VP.t7 82.7821
R37 VP.n0 VP.t1 82.7821
R38 VP.n11 VP.t0 82.7821
R39 VP.n15 VP.t5 82.7821
R40 VP.n20 VP.t6 82.7821
R41 VP.n43 VP.n42 67.0082
R42 VP.n76 VP.n0 67.0082
R43 VP.n41 VP.n11 67.0082
R44 VP.n49 VP.n48 56.4773
R45 VP.n37 VP.n13 56.4773
R46 VP.n61 VP.n6 56.4773
R47 VP.n72 VP.n2 56.4773
R48 VP.n26 VP.n17 56.4773
R49 VP.n42 VP.n41 52.7794
R50 VP.n20 VP.n19 49.9216
R51 VP.n44 VP.n10 24.3439
R52 VP.n48 VP.n10 24.3439
R53 VP.n50 VP.n49 24.3439
R54 VP.n50 VP.n8 24.3439
R55 VP.n54 VP.n8 24.3439
R56 VP.n57 VP.n56 24.3439
R57 VP.n57 VP.n6 24.3439
R58 VP.n62 VP.n61 24.3439
R59 VP.n63 VP.n62 24.3439
R60 VP.n67 VP.n66 24.3439
R61 VP.n68 VP.n67 24.3439
R62 VP.n68 VP.n2 24.3439
R63 VP.n73 VP.n72 24.3439
R64 VP.n74 VP.n73 24.3439
R65 VP.n38 VP.n37 24.3439
R66 VP.n39 VP.n38 24.3439
R67 VP.n27 VP.n26 24.3439
R68 VP.n28 VP.n27 24.3439
R69 VP.n32 VP.n31 24.3439
R70 VP.n33 VP.n32 24.3439
R71 VP.n33 VP.n13 24.3439
R72 VP.n22 VP.n21 24.3439
R73 VP.n22 VP.n17 24.3439
R74 VP.n56 VP.n55 23.8571
R75 VP.n63 VP.n4 23.8571
R76 VP.n28 VP.n15 23.8571
R77 VP.n21 VP.n20 23.8571
R78 VP.n44 VP.n43 22.8833
R79 VP.n74 VP.n0 22.8833
R80 VP.n39 VP.n11 22.8833
R81 VP.n19 VP.n18 3.785
R82 VP.n55 VP.n54 0.487369
R83 VP.n66 VP.n4 0.487369
R84 VP.n31 VP.n15 0.487369
R85 VP.n41 VP.n40 0.355081
R86 VP.n45 VP.n42 0.355081
R87 VP.n76 VP.n75 0.355081
R88 VP VP.n76 0.26685
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VTAIL.n466 VTAIL.n414 756.745
R121 VTAIL.n54 VTAIL.n2 756.745
R122 VTAIL.n112 VTAIL.n60 756.745
R123 VTAIL.n172 VTAIL.n120 756.745
R124 VTAIL.n408 VTAIL.n356 756.745
R125 VTAIL.n348 VTAIL.n296 756.745
R126 VTAIL.n290 VTAIL.n238 756.745
R127 VTAIL.n230 VTAIL.n178 756.745
R128 VTAIL.n433 VTAIL.n432 585
R129 VTAIL.n430 VTAIL.n429 585
R130 VTAIL.n439 VTAIL.n438 585
R131 VTAIL.n441 VTAIL.n440 585
R132 VTAIL.n426 VTAIL.n425 585
R133 VTAIL.n447 VTAIL.n446 585
R134 VTAIL.n450 VTAIL.n449 585
R135 VTAIL.n448 VTAIL.n422 585
R136 VTAIL.n455 VTAIL.n421 585
R137 VTAIL.n457 VTAIL.n456 585
R138 VTAIL.n459 VTAIL.n458 585
R139 VTAIL.n418 VTAIL.n417 585
R140 VTAIL.n465 VTAIL.n464 585
R141 VTAIL.n467 VTAIL.n466 585
R142 VTAIL.n21 VTAIL.n20 585
R143 VTAIL.n18 VTAIL.n17 585
R144 VTAIL.n27 VTAIL.n26 585
R145 VTAIL.n29 VTAIL.n28 585
R146 VTAIL.n14 VTAIL.n13 585
R147 VTAIL.n35 VTAIL.n34 585
R148 VTAIL.n38 VTAIL.n37 585
R149 VTAIL.n36 VTAIL.n10 585
R150 VTAIL.n43 VTAIL.n9 585
R151 VTAIL.n45 VTAIL.n44 585
R152 VTAIL.n47 VTAIL.n46 585
R153 VTAIL.n6 VTAIL.n5 585
R154 VTAIL.n53 VTAIL.n52 585
R155 VTAIL.n55 VTAIL.n54 585
R156 VTAIL.n79 VTAIL.n78 585
R157 VTAIL.n76 VTAIL.n75 585
R158 VTAIL.n85 VTAIL.n84 585
R159 VTAIL.n87 VTAIL.n86 585
R160 VTAIL.n72 VTAIL.n71 585
R161 VTAIL.n93 VTAIL.n92 585
R162 VTAIL.n96 VTAIL.n95 585
R163 VTAIL.n94 VTAIL.n68 585
R164 VTAIL.n101 VTAIL.n67 585
R165 VTAIL.n103 VTAIL.n102 585
R166 VTAIL.n105 VTAIL.n104 585
R167 VTAIL.n64 VTAIL.n63 585
R168 VTAIL.n111 VTAIL.n110 585
R169 VTAIL.n113 VTAIL.n112 585
R170 VTAIL.n139 VTAIL.n138 585
R171 VTAIL.n136 VTAIL.n135 585
R172 VTAIL.n145 VTAIL.n144 585
R173 VTAIL.n147 VTAIL.n146 585
R174 VTAIL.n132 VTAIL.n131 585
R175 VTAIL.n153 VTAIL.n152 585
R176 VTAIL.n156 VTAIL.n155 585
R177 VTAIL.n154 VTAIL.n128 585
R178 VTAIL.n161 VTAIL.n127 585
R179 VTAIL.n163 VTAIL.n162 585
R180 VTAIL.n165 VTAIL.n164 585
R181 VTAIL.n124 VTAIL.n123 585
R182 VTAIL.n171 VTAIL.n170 585
R183 VTAIL.n173 VTAIL.n172 585
R184 VTAIL.n409 VTAIL.n408 585
R185 VTAIL.n407 VTAIL.n406 585
R186 VTAIL.n360 VTAIL.n359 585
R187 VTAIL.n401 VTAIL.n400 585
R188 VTAIL.n399 VTAIL.n398 585
R189 VTAIL.n397 VTAIL.n363 585
R190 VTAIL.n367 VTAIL.n364 585
R191 VTAIL.n392 VTAIL.n391 585
R192 VTAIL.n390 VTAIL.n389 585
R193 VTAIL.n369 VTAIL.n368 585
R194 VTAIL.n384 VTAIL.n383 585
R195 VTAIL.n382 VTAIL.n381 585
R196 VTAIL.n373 VTAIL.n372 585
R197 VTAIL.n376 VTAIL.n375 585
R198 VTAIL.n349 VTAIL.n348 585
R199 VTAIL.n347 VTAIL.n346 585
R200 VTAIL.n300 VTAIL.n299 585
R201 VTAIL.n341 VTAIL.n340 585
R202 VTAIL.n339 VTAIL.n338 585
R203 VTAIL.n337 VTAIL.n303 585
R204 VTAIL.n307 VTAIL.n304 585
R205 VTAIL.n332 VTAIL.n331 585
R206 VTAIL.n330 VTAIL.n329 585
R207 VTAIL.n309 VTAIL.n308 585
R208 VTAIL.n324 VTAIL.n323 585
R209 VTAIL.n322 VTAIL.n321 585
R210 VTAIL.n313 VTAIL.n312 585
R211 VTAIL.n316 VTAIL.n315 585
R212 VTAIL.n291 VTAIL.n290 585
R213 VTAIL.n289 VTAIL.n288 585
R214 VTAIL.n242 VTAIL.n241 585
R215 VTAIL.n283 VTAIL.n282 585
R216 VTAIL.n281 VTAIL.n280 585
R217 VTAIL.n279 VTAIL.n245 585
R218 VTAIL.n249 VTAIL.n246 585
R219 VTAIL.n274 VTAIL.n273 585
R220 VTAIL.n272 VTAIL.n271 585
R221 VTAIL.n251 VTAIL.n250 585
R222 VTAIL.n266 VTAIL.n265 585
R223 VTAIL.n264 VTAIL.n263 585
R224 VTAIL.n255 VTAIL.n254 585
R225 VTAIL.n258 VTAIL.n257 585
R226 VTAIL.n231 VTAIL.n230 585
R227 VTAIL.n229 VTAIL.n228 585
R228 VTAIL.n182 VTAIL.n181 585
R229 VTAIL.n223 VTAIL.n222 585
R230 VTAIL.n221 VTAIL.n220 585
R231 VTAIL.n219 VTAIL.n185 585
R232 VTAIL.n189 VTAIL.n186 585
R233 VTAIL.n214 VTAIL.n213 585
R234 VTAIL.n212 VTAIL.n211 585
R235 VTAIL.n191 VTAIL.n190 585
R236 VTAIL.n206 VTAIL.n205 585
R237 VTAIL.n204 VTAIL.n203 585
R238 VTAIL.n195 VTAIL.n194 585
R239 VTAIL.n198 VTAIL.n197 585
R240 VTAIL.t12 VTAIL.n374 329.038
R241 VTAIL.t11 VTAIL.n314 329.038
R242 VTAIL.t6 VTAIL.n256 329.038
R243 VTAIL.t4 VTAIL.n196 329.038
R244 VTAIL.t0 VTAIL.n431 329.038
R245 VTAIL.t5 VTAIL.n19 329.038
R246 VTAIL.t15 VTAIL.n77 329.038
R247 VTAIL.t9 VTAIL.n137 329.038
R248 VTAIL.n432 VTAIL.n429 171.744
R249 VTAIL.n439 VTAIL.n429 171.744
R250 VTAIL.n440 VTAIL.n439 171.744
R251 VTAIL.n440 VTAIL.n425 171.744
R252 VTAIL.n447 VTAIL.n425 171.744
R253 VTAIL.n449 VTAIL.n447 171.744
R254 VTAIL.n449 VTAIL.n448 171.744
R255 VTAIL.n448 VTAIL.n421 171.744
R256 VTAIL.n457 VTAIL.n421 171.744
R257 VTAIL.n458 VTAIL.n457 171.744
R258 VTAIL.n458 VTAIL.n417 171.744
R259 VTAIL.n465 VTAIL.n417 171.744
R260 VTAIL.n466 VTAIL.n465 171.744
R261 VTAIL.n20 VTAIL.n17 171.744
R262 VTAIL.n27 VTAIL.n17 171.744
R263 VTAIL.n28 VTAIL.n27 171.744
R264 VTAIL.n28 VTAIL.n13 171.744
R265 VTAIL.n35 VTAIL.n13 171.744
R266 VTAIL.n37 VTAIL.n35 171.744
R267 VTAIL.n37 VTAIL.n36 171.744
R268 VTAIL.n36 VTAIL.n9 171.744
R269 VTAIL.n45 VTAIL.n9 171.744
R270 VTAIL.n46 VTAIL.n45 171.744
R271 VTAIL.n46 VTAIL.n5 171.744
R272 VTAIL.n53 VTAIL.n5 171.744
R273 VTAIL.n54 VTAIL.n53 171.744
R274 VTAIL.n78 VTAIL.n75 171.744
R275 VTAIL.n85 VTAIL.n75 171.744
R276 VTAIL.n86 VTAIL.n85 171.744
R277 VTAIL.n86 VTAIL.n71 171.744
R278 VTAIL.n93 VTAIL.n71 171.744
R279 VTAIL.n95 VTAIL.n93 171.744
R280 VTAIL.n95 VTAIL.n94 171.744
R281 VTAIL.n94 VTAIL.n67 171.744
R282 VTAIL.n103 VTAIL.n67 171.744
R283 VTAIL.n104 VTAIL.n103 171.744
R284 VTAIL.n104 VTAIL.n63 171.744
R285 VTAIL.n111 VTAIL.n63 171.744
R286 VTAIL.n112 VTAIL.n111 171.744
R287 VTAIL.n138 VTAIL.n135 171.744
R288 VTAIL.n145 VTAIL.n135 171.744
R289 VTAIL.n146 VTAIL.n145 171.744
R290 VTAIL.n146 VTAIL.n131 171.744
R291 VTAIL.n153 VTAIL.n131 171.744
R292 VTAIL.n155 VTAIL.n153 171.744
R293 VTAIL.n155 VTAIL.n154 171.744
R294 VTAIL.n154 VTAIL.n127 171.744
R295 VTAIL.n163 VTAIL.n127 171.744
R296 VTAIL.n164 VTAIL.n163 171.744
R297 VTAIL.n164 VTAIL.n123 171.744
R298 VTAIL.n171 VTAIL.n123 171.744
R299 VTAIL.n172 VTAIL.n171 171.744
R300 VTAIL.n408 VTAIL.n407 171.744
R301 VTAIL.n407 VTAIL.n359 171.744
R302 VTAIL.n400 VTAIL.n359 171.744
R303 VTAIL.n400 VTAIL.n399 171.744
R304 VTAIL.n399 VTAIL.n363 171.744
R305 VTAIL.n367 VTAIL.n363 171.744
R306 VTAIL.n391 VTAIL.n367 171.744
R307 VTAIL.n391 VTAIL.n390 171.744
R308 VTAIL.n390 VTAIL.n368 171.744
R309 VTAIL.n383 VTAIL.n368 171.744
R310 VTAIL.n383 VTAIL.n382 171.744
R311 VTAIL.n382 VTAIL.n372 171.744
R312 VTAIL.n375 VTAIL.n372 171.744
R313 VTAIL.n348 VTAIL.n347 171.744
R314 VTAIL.n347 VTAIL.n299 171.744
R315 VTAIL.n340 VTAIL.n299 171.744
R316 VTAIL.n340 VTAIL.n339 171.744
R317 VTAIL.n339 VTAIL.n303 171.744
R318 VTAIL.n307 VTAIL.n303 171.744
R319 VTAIL.n331 VTAIL.n307 171.744
R320 VTAIL.n331 VTAIL.n330 171.744
R321 VTAIL.n330 VTAIL.n308 171.744
R322 VTAIL.n323 VTAIL.n308 171.744
R323 VTAIL.n323 VTAIL.n322 171.744
R324 VTAIL.n322 VTAIL.n312 171.744
R325 VTAIL.n315 VTAIL.n312 171.744
R326 VTAIL.n290 VTAIL.n289 171.744
R327 VTAIL.n289 VTAIL.n241 171.744
R328 VTAIL.n282 VTAIL.n241 171.744
R329 VTAIL.n282 VTAIL.n281 171.744
R330 VTAIL.n281 VTAIL.n245 171.744
R331 VTAIL.n249 VTAIL.n245 171.744
R332 VTAIL.n273 VTAIL.n249 171.744
R333 VTAIL.n273 VTAIL.n272 171.744
R334 VTAIL.n272 VTAIL.n250 171.744
R335 VTAIL.n265 VTAIL.n250 171.744
R336 VTAIL.n265 VTAIL.n264 171.744
R337 VTAIL.n264 VTAIL.n254 171.744
R338 VTAIL.n257 VTAIL.n254 171.744
R339 VTAIL.n230 VTAIL.n229 171.744
R340 VTAIL.n229 VTAIL.n181 171.744
R341 VTAIL.n222 VTAIL.n181 171.744
R342 VTAIL.n222 VTAIL.n221 171.744
R343 VTAIL.n221 VTAIL.n185 171.744
R344 VTAIL.n189 VTAIL.n185 171.744
R345 VTAIL.n213 VTAIL.n189 171.744
R346 VTAIL.n213 VTAIL.n212 171.744
R347 VTAIL.n212 VTAIL.n190 171.744
R348 VTAIL.n205 VTAIL.n190 171.744
R349 VTAIL.n205 VTAIL.n204 171.744
R350 VTAIL.n204 VTAIL.n194 171.744
R351 VTAIL.n197 VTAIL.n194 171.744
R352 VTAIL.n432 VTAIL.t0 85.8723
R353 VTAIL.n20 VTAIL.t5 85.8723
R354 VTAIL.n78 VTAIL.t15 85.8723
R355 VTAIL.n138 VTAIL.t9 85.8723
R356 VTAIL.n375 VTAIL.t12 85.8723
R357 VTAIL.n315 VTAIL.t11 85.8723
R358 VTAIL.n257 VTAIL.t6 85.8723
R359 VTAIL.n197 VTAIL.t4 85.8723
R360 VTAIL.n355 VTAIL.n354 61.9025
R361 VTAIL.n237 VTAIL.n236 61.9025
R362 VTAIL.n1 VTAIL.n0 61.9023
R363 VTAIL.n119 VTAIL.n118 61.9023
R364 VTAIL.n471 VTAIL.n470 34.9005
R365 VTAIL.n59 VTAIL.n58 34.9005
R366 VTAIL.n117 VTAIL.n116 34.9005
R367 VTAIL.n177 VTAIL.n176 34.9005
R368 VTAIL.n413 VTAIL.n412 34.9005
R369 VTAIL.n353 VTAIL.n352 34.9005
R370 VTAIL.n295 VTAIL.n294 34.9005
R371 VTAIL.n235 VTAIL.n234 34.9005
R372 VTAIL.n471 VTAIL.n413 24.6945
R373 VTAIL.n235 VTAIL.n177 24.6945
R374 VTAIL.n456 VTAIL.n455 13.1884
R375 VTAIL.n44 VTAIL.n43 13.1884
R376 VTAIL.n102 VTAIL.n101 13.1884
R377 VTAIL.n162 VTAIL.n161 13.1884
R378 VTAIL.n398 VTAIL.n397 13.1884
R379 VTAIL.n338 VTAIL.n337 13.1884
R380 VTAIL.n280 VTAIL.n279 13.1884
R381 VTAIL.n220 VTAIL.n219 13.1884
R382 VTAIL.n454 VTAIL.n422 12.8005
R383 VTAIL.n459 VTAIL.n420 12.8005
R384 VTAIL.n42 VTAIL.n10 12.8005
R385 VTAIL.n47 VTAIL.n8 12.8005
R386 VTAIL.n100 VTAIL.n68 12.8005
R387 VTAIL.n105 VTAIL.n66 12.8005
R388 VTAIL.n160 VTAIL.n128 12.8005
R389 VTAIL.n165 VTAIL.n126 12.8005
R390 VTAIL.n401 VTAIL.n362 12.8005
R391 VTAIL.n396 VTAIL.n364 12.8005
R392 VTAIL.n341 VTAIL.n302 12.8005
R393 VTAIL.n336 VTAIL.n304 12.8005
R394 VTAIL.n283 VTAIL.n244 12.8005
R395 VTAIL.n278 VTAIL.n246 12.8005
R396 VTAIL.n223 VTAIL.n184 12.8005
R397 VTAIL.n218 VTAIL.n186 12.8005
R398 VTAIL.n451 VTAIL.n450 12.0247
R399 VTAIL.n460 VTAIL.n418 12.0247
R400 VTAIL.n39 VTAIL.n38 12.0247
R401 VTAIL.n48 VTAIL.n6 12.0247
R402 VTAIL.n97 VTAIL.n96 12.0247
R403 VTAIL.n106 VTAIL.n64 12.0247
R404 VTAIL.n157 VTAIL.n156 12.0247
R405 VTAIL.n166 VTAIL.n124 12.0247
R406 VTAIL.n402 VTAIL.n360 12.0247
R407 VTAIL.n393 VTAIL.n392 12.0247
R408 VTAIL.n342 VTAIL.n300 12.0247
R409 VTAIL.n333 VTAIL.n332 12.0247
R410 VTAIL.n284 VTAIL.n242 12.0247
R411 VTAIL.n275 VTAIL.n274 12.0247
R412 VTAIL.n224 VTAIL.n182 12.0247
R413 VTAIL.n215 VTAIL.n214 12.0247
R414 VTAIL.n446 VTAIL.n424 11.249
R415 VTAIL.n464 VTAIL.n463 11.249
R416 VTAIL.n34 VTAIL.n12 11.249
R417 VTAIL.n52 VTAIL.n51 11.249
R418 VTAIL.n92 VTAIL.n70 11.249
R419 VTAIL.n110 VTAIL.n109 11.249
R420 VTAIL.n152 VTAIL.n130 11.249
R421 VTAIL.n170 VTAIL.n169 11.249
R422 VTAIL.n406 VTAIL.n405 11.249
R423 VTAIL.n389 VTAIL.n366 11.249
R424 VTAIL.n346 VTAIL.n345 11.249
R425 VTAIL.n329 VTAIL.n306 11.249
R426 VTAIL.n288 VTAIL.n287 11.249
R427 VTAIL.n271 VTAIL.n248 11.249
R428 VTAIL.n228 VTAIL.n227 11.249
R429 VTAIL.n211 VTAIL.n188 11.249
R430 VTAIL.n433 VTAIL.n431 10.7239
R431 VTAIL.n21 VTAIL.n19 10.7239
R432 VTAIL.n79 VTAIL.n77 10.7239
R433 VTAIL.n139 VTAIL.n137 10.7239
R434 VTAIL.n376 VTAIL.n374 10.7239
R435 VTAIL.n316 VTAIL.n314 10.7239
R436 VTAIL.n258 VTAIL.n256 10.7239
R437 VTAIL.n198 VTAIL.n196 10.7239
R438 VTAIL.n445 VTAIL.n426 10.4732
R439 VTAIL.n467 VTAIL.n416 10.4732
R440 VTAIL.n33 VTAIL.n14 10.4732
R441 VTAIL.n55 VTAIL.n4 10.4732
R442 VTAIL.n91 VTAIL.n72 10.4732
R443 VTAIL.n113 VTAIL.n62 10.4732
R444 VTAIL.n151 VTAIL.n132 10.4732
R445 VTAIL.n173 VTAIL.n122 10.4732
R446 VTAIL.n409 VTAIL.n358 10.4732
R447 VTAIL.n388 VTAIL.n369 10.4732
R448 VTAIL.n349 VTAIL.n298 10.4732
R449 VTAIL.n328 VTAIL.n309 10.4732
R450 VTAIL.n291 VTAIL.n240 10.4732
R451 VTAIL.n270 VTAIL.n251 10.4732
R452 VTAIL.n231 VTAIL.n180 10.4732
R453 VTAIL.n210 VTAIL.n191 10.4732
R454 VTAIL.n442 VTAIL.n441 9.69747
R455 VTAIL.n468 VTAIL.n414 9.69747
R456 VTAIL.n30 VTAIL.n29 9.69747
R457 VTAIL.n56 VTAIL.n2 9.69747
R458 VTAIL.n88 VTAIL.n87 9.69747
R459 VTAIL.n114 VTAIL.n60 9.69747
R460 VTAIL.n148 VTAIL.n147 9.69747
R461 VTAIL.n174 VTAIL.n120 9.69747
R462 VTAIL.n410 VTAIL.n356 9.69747
R463 VTAIL.n385 VTAIL.n384 9.69747
R464 VTAIL.n350 VTAIL.n296 9.69747
R465 VTAIL.n325 VTAIL.n324 9.69747
R466 VTAIL.n292 VTAIL.n238 9.69747
R467 VTAIL.n267 VTAIL.n266 9.69747
R468 VTAIL.n232 VTAIL.n178 9.69747
R469 VTAIL.n207 VTAIL.n206 9.69747
R470 VTAIL.n470 VTAIL.n469 9.45567
R471 VTAIL.n58 VTAIL.n57 9.45567
R472 VTAIL.n116 VTAIL.n115 9.45567
R473 VTAIL.n176 VTAIL.n175 9.45567
R474 VTAIL.n412 VTAIL.n411 9.45567
R475 VTAIL.n352 VTAIL.n351 9.45567
R476 VTAIL.n294 VTAIL.n293 9.45567
R477 VTAIL.n234 VTAIL.n233 9.45567
R478 VTAIL.n469 VTAIL.n468 9.3005
R479 VTAIL.n416 VTAIL.n415 9.3005
R480 VTAIL.n463 VTAIL.n462 9.3005
R481 VTAIL.n461 VTAIL.n460 9.3005
R482 VTAIL.n420 VTAIL.n419 9.3005
R483 VTAIL.n435 VTAIL.n434 9.3005
R484 VTAIL.n437 VTAIL.n436 9.3005
R485 VTAIL.n428 VTAIL.n427 9.3005
R486 VTAIL.n443 VTAIL.n442 9.3005
R487 VTAIL.n445 VTAIL.n444 9.3005
R488 VTAIL.n424 VTAIL.n423 9.3005
R489 VTAIL.n452 VTAIL.n451 9.3005
R490 VTAIL.n454 VTAIL.n453 9.3005
R491 VTAIL.n57 VTAIL.n56 9.3005
R492 VTAIL.n4 VTAIL.n3 9.3005
R493 VTAIL.n51 VTAIL.n50 9.3005
R494 VTAIL.n49 VTAIL.n48 9.3005
R495 VTAIL.n8 VTAIL.n7 9.3005
R496 VTAIL.n23 VTAIL.n22 9.3005
R497 VTAIL.n25 VTAIL.n24 9.3005
R498 VTAIL.n16 VTAIL.n15 9.3005
R499 VTAIL.n31 VTAIL.n30 9.3005
R500 VTAIL.n33 VTAIL.n32 9.3005
R501 VTAIL.n12 VTAIL.n11 9.3005
R502 VTAIL.n40 VTAIL.n39 9.3005
R503 VTAIL.n42 VTAIL.n41 9.3005
R504 VTAIL.n115 VTAIL.n114 9.3005
R505 VTAIL.n62 VTAIL.n61 9.3005
R506 VTAIL.n109 VTAIL.n108 9.3005
R507 VTAIL.n107 VTAIL.n106 9.3005
R508 VTAIL.n66 VTAIL.n65 9.3005
R509 VTAIL.n81 VTAIL.n80 9.3005
R510 VTAIL.n83 VTAIL.n82 9.3005
R511 VTAIL.n74 VTAIL.n73 9.3005
R512 VTAIL.n89 VTAIL.n88 9.3005
R513 VTAIL.n91 VTAIL.n90 9.3005
R514 VTAIL.n70 VTAIL.n69 9.3005
R515 VTAIL.n98 VTAIL.n97 9.3005
R516 VTAIL.n100 VTAIL.n99 9.3005
R517 VTAIL.n175 VTAIL.n174 9.3005
R518 VTAIL.n122 VTAIL.n121 9.3005
R519 VTAIL.n169 VTAIL.n168 9.3005
R520 VTAIL.n167 VTAIL.n166 9.3005
R521 VTAIL.n126 VTAIL.n125 9.3005
R522 VTAIL.n141 VTAIL.n140 9.3005
R523 VTAIL.n143 VTAIL.n142 9.3005
R524 VTAIL.n134 VTAIL.n133 9.3005
R525 VTAIL.n149 VTAIL.n148 9.3005
R526 VTAIL.n151 VTAIL.n150 9.3005
R527 VTAIL.n130 VTAIL.n129 9.3005
R528 VTAIL.n158 VTAIL.n157 9.3005
R529 VTAIL.n160 VTAIL.n159 9.3005
R530 VTAIL.n378 VTAIL.n377 9.3005
R531 VTAIL.n380 VTAIL.n379 9.3005
R532 VTAIL.n371 VTAIL.n370 9.3005
R533 VTAIL.n386 VTAIL.n385 9.3005
R534 VTAIL.n388 VTAIL.n387 9.3005
R535 VTAIL.n366 VTAIL.n365 9.3005
R536 VTAIL.n394 VTAIL.n393 9.3005
R537 VTAIL.n396 VTAIL.n395 9.3005
R538 VTAIL.n411 VTAIL.n410 9.3005
R539 VTAIL.n358 VTAIL.n357 9.3005
R540 VTAIL.n405 VTAIL.n404 9.3005
R541 VTAIL.n403 VTAIL.n402 9.3005
R542 VTAIL.n362 VTAIL.n361 9.3005
R543 VTAIL.n318 VTAIL.n317 9.3005
R544 VTAIL.n320 VTAIL.n319 9.3005
R545 VTAIL.n311 VTAIL.n310 9.3005
R546 VTAIL.n326 VTAIL.n325 9.3005
R547 VTAIL.n328 VTAIL.n327 9.3005
R548 VTAIL.n306 VTAIL.n305 9.3005
R549 VTAIL.n334 VTAIL.n333 9.3005
R550 VTAIL.n336 VTAIL.n335 9.3005
R551 VTAIL.n351 VTAIL.n350 9.3005
R552 VTAIL.n298 VTAIL.n297 9.3005
R553 VTAIL.n345 VTAIL.n344 9.3005
R554 VTAIL.n343 VTAIL.n342 9.3005
R555 VTAIL.n302 VTAIL.n301 9.3005
R556 VTAIL.n260 VTAIL.n259 9.3005
R557 VTAIL.n262 VTAIL.n261 9.3005
R558 VTAIL.n253 VTAIL.n252 9.3005
R559 VTAIL.n268 VTAIL.n267 9.3005
R560 VTAIL.n270 VTAIL.n269 9.3005
R561 VTAIL.n248 VTAIL.n247 9.3005
R562 VTAIL.n276 VTAIL.n275 9.3005
R563 VTAIL.n278 VTAIL.n277 9.3005
R564 VTAIL.n293 VTAIL.n292 9.3005
R565 VTAIL.n240 VTAIL.n239 9.3005
R566 VTAIL.n287 VTAIL.n286 9.3005
R567 VTAIL.n285 VTAIL.n284 9.3005
R568 VTAIL.n244 VTAIL.n243 9.3005
R569 VTAIL.n200 VTAIL.n199 9.3005
R570 VTAIL.n202 VTAIL.n201 9.3005
R571 VTAIL.n193 VTAIL.n192 9.3005
R572 VTAIL.n208 VTAIL.n207 9.3005
R573 VTAIL.n210 VTAIL.n209 9.3005
R574 VTAIL.n188 VTAIL.n187 9.3005
R575 VTAIL.n216 VTAIL.n215 9.3005
R576 VTAIL.n218 VTAIL.n217 9.3005
R577 VTAIL.n233 VTAIL.n232 9.3005
R578 VTAIL.n180 VTAIL.n179 9.3005
R579 VTAIL.n227 VTAIL.n226 9.3005
R580 VTAIL.n225 VTAIL.n224 9.3005
R581 VTAIL.n184 VTAIL.n183 9.3005
R582 VTAIL.n438 VTAIL.n428 8.92171
R583 VTAIL.n26 VTAIL.n16 8.92171
R584 VTAIL.n84 VTAIL.n74 8.92171
R585 VTAIL.n144 VTAIL.n134 8.92171
R586 VTAIL.n381 VTAIL.n371 8.92171
R587 VTAIL.n321 VTAIL.n311 8.92171
R588 VTAIL.n263 VTAIL.n253 8.92171
R589 VTAIL.n203 VTAIL.n193 8.92171
R590 VTAIL.n437 VTAIL.n430 8.14595
R591 VTAIL.n25 VTAIL.n18 8.14595
R592 VTAIL.n83 VTAIL.n76 8.14595
R593 VTAIL.n143 VTAIL.n136 8.14595
R594 VTAIL.n380 VTAIL.n373 8.14595
R595 VTAIL.n320 VTAIL.n313 8.14595
R596 VTAIL.n262 VTAIL.n255 8.14595
R597 VTAIL.n202 VTAIL.n195 8.14595
R598 VTAIL.n434 VTAIL.n433 7.3702
R599 VTAIL.n22 VTAIL.n21 7.3702
R600 VTAIL.n80 VTAIL.n79 7.3702
R601 VTAIL.n140 VTAIL.n139 7.3702
R602 VTAIL.n377 VTAIL.n376 7.3702
R603 VTAIL.n317 VTAIL.n316 7.3702
R604 VTAIL.n259 VTAIL.n258 7.3702
R605 VTAIL.n199 VTAIL.n198 7.3702
R606 VTAIL.n434 VTAIL.n430 5.81868
R607 VTAIL.n22 VTAIL.n18 5.81868
R608 VTAIL.n80 VTAIL.n76 5.81868
R609 VTAIL.n140 VTAIL.n136 5.81868
R610 VTAIL.n377 VTAIL.n373 5.81868
R611 VTAIL.n317 VTAIL.n313 5.81868
R612 VTAIL.n259 VTAIL.n255 5.81868
R613 VTAIL.n199 VTAIL.n195 5.81868
R614 VTAIL.n438 VTAIL.n437 5.04292
R615 VTAIL.n26 VTAIL.n25 5.04292
R616 VTAIL.n84 VTAIL.n83 5.04292
R617 VTAIL.n144 VTAIL.n143 5.04292
R618 VTAIL.n381 VTAIL.n380 5.04292
R619 VTAIL.n321 VTAIL.n320 5.04292
R620 VTAIL.n263 VTAIL.n262 5.04292
R621 VTAIL.n203 VTAIL.n202 5.04292
R622 VTAIL.n441 VTAIL.n428 4.26717
R623 VTAIL.n470 VTAIL.n414 4.26717
R624 VTAIL.n29 VTAIL.n16 4.26717
R625 VTAIL.n58 VTAIL.n2 4.26717
R626 VTAIL.n87 VTAIL.n74 4.26717
R627 VTAIL.n116 VTAIL.n60 4.26717
R628 VTAIL.n147 VTAIL.n134 4.26717
R629 VTAIL.n176 VTAIL.n120 4.26717
R630 VTAIL.n412 VTAIL.n356 4.26717
R631 VTAIL.n384 VTAIL.n371 4.26717
R632 VTAIL.n352 VTAIL.n296 4.26717
R633 VTAIL.n324 VTAIL.n311 4.26717
R634 VTAIL.n294 VTAIL.n238 4.26717
R635 VTAIL.n266 VTAIL.n253 4.26717
R636 VTAIL.n234 VTAIL.n178 4.26717
R637 VTAIL.n206 VTAIL.n193 4.26717
R638 VTAIL.n442 VTAIL.n426 3.49141
R639 VTAIL.n468 VTAIL.n467 3.49141
R640 VTAIL.n30 VTAIL.n14 3.49141
R641 VTAIL.n56 VTAIL.n55 3.49141
R642 VTAIL.n88 VTAIL.n72 3.49141
R643 VTAIL.n114 VTAIL.n113 3.49141
R644 VTAIL.n148 VTAIL.n132 3.49141
R645 VTAIL.n174 VTAIL.n173 3.49141
R646 VTAIL.n410 VTAIL.n409 3.49141
R647 VTAIL.n385 VTAIL.n369 3.49141
R648 VTAIL.n350 VTAIL.n349 3.49141
R649 VTAIL.n325 VTAIL.n309 3.49141
R650 VTAIL.n292 VTAIL.n291 3.49141
R651 VTAIL.n267 VTAIL.n251 3.49141
R652 VTAIL.n232 VTAIL.n231 3.49141
R653 VTAIL.n207 VTAIL.n191 3.49141
R654 VTAIL.n0 VTAIL.t7 3.00466
R655 VTAIL.n0 VTAIL.t3 3.00466
R656 VTAIL.n118 VTAIL.t8 3.00466
R657 VTAIL.n118 VTAIL.t13 3.00466
R658 VTAIL.n354 VTAIL.t10 3.00466
R659 VTAIL.n354 VTAIL.t14 3.00466
R660 VTAIL.n236 VTAIL.t1 3.00466
R661 VTAIL.n236 VTAIL.t2 3.00466
R662 VTAIL.n237 VTAIL.n235 3.0005
R663 VTAIL.n295 VTAIL.n237 3.0005
R664 VTAIL.n355 VTAIL.n353 3.0005
R665 VTAIL.n413 VTAIL.n355 3.0005
R666 VTAIL.n177 VTAIL.n119 3.0005
R667 VTAIL.n119 VTAIL.n117 3.0005
R668 VTAIL.n59 VTAIL.n1 3.0005
R669 VTAIL VTAIL.n471 2.94231
R670 VTAIL.n446 VTAIL.n445 2.71565
R671 VTAIL.n464 VTAIL.n416 2.71565
R672 VTAIL.n34 VTAIL.n33 2.71565
R673 VTAIL.n52 VTAIL.n4 2.71565
R674 VTAIL.n92 VTAIL.n91 2.71565
R675 VTAIL.n110 VTAIL.n62 2.71565
R676 VTAIL.n152 VTAIL.n151 2.71565
R677 VTAIL.n170 VTAIL.n122 2.71565
R678 VTAIL.n406 VTAIL.n358 2.71565
R679 VTAIL.n389 VTAIL.n388 2.71565
R680 VTAIL.n346 VTAIL.n298 2.71565
R681 VTAIL.n329 VTAIL.n328 2.71565
R682 VTAIL.n288 VTAIL.n240 2.71565
R683 VTAIL.n271 VTAIL.n270 2.71565
R684 VTAIL.n228 VTAIL.n180 2.71565
R685 VTAIL.n211 VTAIL.n210 2.71565
R686 VTAIL.n435 VTAIL.n431 2.41282
R687 VTAIL.n23 VTAIL.n19 2.41282
R688 VTAIL.n81 VTAIL.n77 2.41282
R689 VTAIL.n141 VTAIL.n137 2.41282
R690 VTAIL.n378 VTAIL.n374 2.41282
R691 VTAIL.n318 VTAIL.n314 2.41282
R692 VTAIL.n260 VTAIL.n256 2.41282
R693 VTAIL.n200 VTAIL.n196 2.41282
R694 VTAIL.n450 VTAIL.n424 1.93989
R695 VTAIL.n463 VTAIL.n418 1.93989
R696 VTAIL.n38 VTAIL.n12 1.93989
R697 VTAIL.n51 VTAIL.n6 1.93989
R698 VTAIL.n96 VTAIL.n70 1.93989
R699 VTAIL.n109 VTAIL.n64 1.93989
R700 VTAIL.n156 VTAIL.n130 1.93989
R701 VTAIL.n169 VTAIL.n124 1.93989
R702 VTAIL.n405 VTAIL.n360 1.93989
R703 VTAIL.n392 VTAIL.n366 1.93989
R704 VTAIL.n345 VTAIL.n300 1.93989
R705 VTAIL.n332 VTAIL.n306 1.93989
R706 VTAIL.n287 VTAIL.n242 1.93989
R707 VTAIL.n274 VTAIL.n248 1.93989
R708 VTAIL.n227 VTAIL.n182 1.93989
R709 VTAIL.n214 VTAIL.n188 1.93989
R710 VTAIL.n451 VTAIL.n422 1.16414
R711 VTAIL.n460 VTAIL.n459 1.16414
R712 VTAIL.n39 VTAIL.n10 1.16414
R713 VTAIL.n48 VTAIL.n47 1.16414
R714 VTAIL.n97 VTAIL.n68 1.16414
R715 VTAIL.n106 VTAIL.n105 1.16414
R716 VTAIL.n157 VTAIL.n128 1.16414
R717 VTAIL.n166 VTAIL.n165 1.16414
R718 VTAIL.n402 VTAIL.n401 1.16414
R719 VTAIL.n393 VTAIL.n364 1.16414
R720 VTAIL.n342 VTAIL.n341 1.16414
R721 VTAIL.n333 VTAIL.n304 1.16414
R722 VTAIL.n284 VTAIL.n283 1.16414
R723 VTAIL.n275 VTAIL.n246 1.16414
R724 VTAIL.n224 VTAIL.n223 1.16414
R725 VTAIL.n215 VTAIL.n186 1.16414
R726 VTAIL.n353 VTAIL.n295 0.470328
R727 VTAIL.n117 VTAIL.n59 0.470328
R728 VTAIL.n455 VTAIL.n454 0.388379
R729 VTAIL.n456 VTAIL.n420 0.388379
R730 VTAIL.n43 VTAIL.n42 0.388379
R731 VTAIL.n44 VTAIL.n8 0.388379
R732 VTAIL.n101 VTAIL.n100 0.388379
R733 VTAIL.n102 VTAIL.n66 0.388379
R734 VTAIL.n161 VTAIL.n160 0.388379
R735 VTAIL.n162 VTAIL.n126 0.388379
R736 VTAIL.n398 VTAIL.n362 0.388379
R737 VTAIL.n397 VTAIL.n396 0.388379
R738 VTAIL.n338 VTAIL.n302 0.388379
R739 VTAIL.n337 VTAIL.n336 0.388379
R740 VTAIL.n280 VTAIL.n244 0.388379
R741 VTAIL.n279 VTAIL.n278 0.388379
R742 VTAIL.n220 VTAIL.n184 0.388379
R743 VTAIL.n219 VTAIL.n218 0.388379
R744 VTAIL.n436 VTAIL.n435 0.155672
R745 VTAIL.n436 VTAIL.n427 0.155672
R746 VTAIL.n443 VTAIL.n427 0.155672
R747 VTAIL.n444 VTAIL.n443 0.155672
R748 VTAIL.n444 VTAIL.n423 0.155672
R749 VTAIL.n452 VTAIL.n423 0.155672
R750 VTAIL.n453 VTAIL.n452 0.155672
R751 VTAIL.n453 VTAIL.n419 0.155672
R752 VTAIL.n461 VTAIL.n419 0.155672
R753 VTAIL.n462 VTAIL.n461 0.155672
R754 VTAIL.n462 VTAIL.n415 0.155672
R755 VTAIL.n469 VTAIL.n415 0.155672
R756 VTAIL.n24 VTAIL.n23 0.155672
R757 VTAIL.n24 VTAIL.n15 0.155672
R758 VTAIL.n31 VTAIL.n15 0.155672
R759 VTAIL.n32 VTAIL.n31 0.155672
R760 VTAIL.n32 VTAIL.n11 0.155672
R761 VTAIL.n40 VTAIL.n11 0.155672
R762 VTAIL.n41 VTAIL.n40 0.155672
R763 VTAIL.n41 VTAIL.n7 0.155672
R764 VTAIL.n49 VTAIL.n7 0.155672
R765 VTAIL.n50 VTAIL.n49 0.155672
R766 VTAIL.n50 VTAIL.n3 0.155672
R767 VTAIL.n57 VTAIL.n3 0.155672
R768 VTAIL.n82 VTAIL.n81 0.155672
R769 VTAIL.n82 VTAIL.n73 0.155672
R770 VTAIL.n89 VTAIL.n73 0.155672
R771 VTAIL.n90 VTAIL.n89 0.155672
R772 VTAIL.n90 VTAIL.n69 0.155672
R773 VTAIL.n98 VTAIL.n69 0.155672
R774 VTAIL.n99 VTAIL.n98 0.155672
R775 VTAIL.n99 VTAIL.n65 0.155672
R776 VTAIL.n107 VTAIL.n65 0.155672
R777 VTAIL.n108 VTAIL.n107 0.155672
R778 VTAIL.n108 VTAIL.n61 0.155672
R779 VTAIL.n115 VTAIL.n61 0.155672
R780 VTAIL.n142 VTAIL.n141 0.155672
R781 VTAIL.n142 VTAIL.n133 0.155672
R782 VTAIL.n149 VTAIL.n133 0.155672
R783 VTAIL.n150 VTAIL.n149 0.155672
R784 VTAIL.n150 VTAIL.n129 0.155672
R785 VTAIL.n158 VTAIL.n129 0.155672
R786 VTAIL.n159 VTAIL.n158 0.155672
R787 VTAIL.n159 VTAIL.n125 0.155672
R788 VTAIL.n167 VTAIL.n125 0.155672
R789 VTAIL.n168 VTAIL.n167 0.155672
R790 VTAIL.n168 VTAIL.n121 0.155672
R791 VTAIL.n175 VTAIL.n121 0.155672
R792 VTAIL.n411 VTAIL.n357 0.155672
R793 VTAIL.n404 VTAIL.n357 0.155672
R794 VTAIL.n404 VTAIL.n403 0.155672
R795 VTAIL.n403 VTAIL.n361 0.155672
R796 VTAIL.n395 VTAIL.n361 0.155672
R797 VTAIL.n395 VTAIL.n394 0.155672
R798 VTAIL.n394 VTAIL.n365 0.155672
R799 VTAIL.n387 VTAIL.n365 0.155672
R800 VTAIL.n387 VTAIL.n386 0.155672
R801 VTAIL.n386 VTAIL.n370 0.155672
R802 VTAIL.n379 VTAIL.n370 0.155672
R803 VTAIL.n379 VTAIL.n378 0.155672
R804 VTAIL.n351 VTAIL.n297 0.155672
R805 VTAIL.n344 VTAIL.n297 0.155672
R806 VTAIL.n344 VTAIL.n343 0.155672
R807 VTAIL.n343 VTAIL.n301 0.155672
R808 VTAIL.n335 VTAIL.n301 0.155672
R809 VTAIL.n335 VTAIL.n334 0.155672
R810 VTAIL.n334 VTAIL.n305 0.155672
R811 VTAIL.n327 VTAIL.n305 0.155672
R812 VTAIL.n327 VTAIL.n326 0.155672
R813 VTAIL.n326 VTAIL.n310 0.155672
R814 VTAIL.n319 VTAIL.n310 0.155672
R815 VTAIL.n319 VTAIL.n318 0.155672
R816 VTAIL.n293 VTAIL.n239 0.155672
R817 VTAIL.n286 VTAIL.n239 0.155672
R818 VTAIL.n286 VTAIL.n285 0.155672
R819 VTAIL.n285 VTAIL.n243 0.155672
R820 VTAIL.n277 VTAIL.n243 0.155672
R821 VTAIL.n277 VTAIL.n276 0.155672
R822 VTAIL.n276 VTAIL.n247 0.155672
R823 VTAIL.n269 VTAIL.n247 0.155672
R824 VTAIL.n269 VTAIL.n268 0.155672
R825 VTAIL.n268 VTAIL.n252 0.155672
R826 VTAIL.n261 VTAIL.n252 0.155672
R827 VTAIL.n261 VTAIL.n260 0.155672
R828 VTAIL.n233 VTAIL.n179 0.155672
R829 VTAIL.n226 VTAIL.n179 0.155672
R830 VTAIL.n226 VTAIL.n225 0.155672
R831 VTAIL.n225 VTAIL.n183 0.155672
R832 VTAIL.n217 VTAIL.n183 0.155672
R833 VTAIL.n217 VTAIL.n216 0.155672
R834 VTAIL.n216 VTAIL.n187 0.155672
R835 VTAIL.n209 VTAIL.n187 0.155672
R836 VTAIL.n209 VTAIL.n208 0.155672
R837 VTAIL.n208 VTAIL.n192 0.155672
R838 VTAIL.n201 VTAIL.n192 0.155672
R839 VTAIL.n201 VTAIL.n200 0.155672
R840 VTAIL VTAIL.n1 0.0586897
R841 VDD1 VDD1.n0 80.1395
R842 VDD1.n3 VDD1.n2 80.0258
R843 VDD1.n3 VDD1.n1 80.0258
R844 VDD1.n5 VDD1.n4 78.5811
R845 VDD1.n5 VDD1.n3 47.1259
R846 VDD1.n4 VDD1.t2 3.00466
R847 VDD1.n4 VDD1.t7 3.00466
R848 VDD1.n0 VDD1.t4 3.00466
R849 VDD1.n0 VDD1.t1 3.00466
R850 VDD1.n2 VDD1.t0 3.00466
R851 VDD1.n2 VDD1.t6 3.00466
R852 VDD1.n1 VDD1.t3 3.00466
R853 VDD1.n1 VDD1.t5 3.00466
R854 VDD1 VDD1.n5 1.44231
R855 VN.n60 VN.n59 161.3
R856 VN.n58 VN.n32 161.3
R857 VN.n57 VN.n56 161.3
R858 VN.n55 VN.n33 161.3
R859 VN.n54 VN.n53 161.3
R860 VN.n52 VN.n34 161.3
R861 VN.n51 VN.n50 161.3
R862 VN.n49 VN.n48 161.3
R863 VN.n47 VN.n36 161.3
R864 VN.n46 VN.n45 161.3
R865 VN.n44 VN.n37 161.3
R866 VN.n43 VN.n42 161.3
R867 VN.n41 VN.n38 161.3
R868 VN.n29 VN.n28 161.3
R869 VN.n27 VN.n1 161.3
R870 VN.n26 VN.n25 161.3
R871 VN.n24 VN.n2 161.3
R872 VN.n23 VN.n22 161.3
R873 VN.n21 VN.n3 161.3
R874 VN.n20 VN.n19 161.3
R875 VN.n18 VN.n17 161.3
R876 VN.n16 VN.n5 161.3
R877 VN.n15 VN.n14 161.3
R878 VN.n13 VN.n6 161.3
R879 VN.n12 VN.n11 161.3
R880 VN.n10 VN.n7 161.3
R881 VN.n8 VN.t0 116.111
R882 VN.n39 VN.t2 116.111
R883 VN.n9 VN.t7 82.7821
R884 VN.n4 VN.t3 82.7821
R885 VN.n0 VN.t1 82.7821
R886 VN.n40 VN.t4 82.7821
R887 VN.n35 VN.t6 82.7821
R888 VN.n31 VN.t5 82.7821
R889 VN.n30 VN.n0 67.0082
R890 VN.n61 VN.n31 67.0082
R891 VN.n15 VN.n6 56.4773
R892 VN.n26 VN.n2 56.4773
R893 VN.n46 VN.n37 56.4773
R894 VN.n57 VN.n33 56.4773
R895 VN VN.n61 52.9449
R896 VN.n9 VN.n8 49.9216
R897 VN.n40 VN.n39 49.9216
R898 VN.n11 VN.n10 24.3439
R899 VN.n11 VN.n6 24.3439
R900 VN.n16 VN.n15 24.3439
R901 VN.n17 VN.n16 24.3439
R902 VN.n21 VN.n20 24.3439
R903 VN.n22 VN.n21 24.3439
R904 VN.n22 VN.n2 24.3439
R905 VN.n27 VN.n26 24.3439
R906 VN.n28 VN.n27 24.3439
R907 VN.n42 VN.n37 24.3439
R908 VN.n42 VN.n41 24.3439
R909 VN.n53 VN.n33 24.3439
R910 VN.n53 VN.n52 24.3439
R911 VN.n52 VN.n51 24.3439
R912 VN.n48 VN.n47 24.3439
R913 VN.n47 VN.n46 24.3439
R914 VN.n59 VN.n58 24.3439
R915 VN.n58 VN.n57 24.3439
R916 VN.n10 VN.n9 23.8571
R917 VN.n17 VN.n4 23.8571
R918 VN.n41 VN.n40 23.8571
R919 VN.n48 VN.n35 23.8571
R920 VN.n28 VN.n0 22.8833
R921 VN.n59 VN.n31 22.8833
R922 VN.n39 VN.n38 3.78503
R923 VN.n8 VN.n7 3.78503
R924 VN.n20 VN.n4 0.487369
R925 VN.n51 VN.n35 0.487369
R926 VN.n61 VN.n60 0.355081
R927 VN.n30 VN.n29 0.355081
R928 VN VN.n30 0.26685
R929 VN.n60 VN.n32 0.189894
R930 VN.n56 VN.n32 0.189894
R931 VN.n56 VN.n55 0.189894
R932 VN.n55 VN.n54 0.189894
R933 VN.n54 VN.n34 0.189894
R934 VN.n50 VN.n34 0.189894
R935 VN.n50 VN.n49 0.189894
R936 VN.n49 VN.n36 0.189894
R937 VN.n45 VN.n36 0.189894
R938 VN.n45 VN.n44 0.189894
R939 VN.n44 VN.n43 0.189894
R940 VN.n43 VN.n38 0.189894
R941 VN.n12 VN.n7 0.189894
R942 VN.n13 VN.n12 0.189894
R943 VN.n14 VN.n13 0.189894
R944 VN.n14 VN.n5 0.189894
R945 VN.n18 VN.n5 0.189894
R946 VN.n19 VN.n18 0.189894
R947 VN.n19 VN.n3 0.189894
R948 VN.n23 VN.n3 0.189894
R949 VN.n24 VN.n23 0.189894
R950 VN.n25 VN.n24 0.189894
R951 VN.n25 VN.n1 0.189894
R952 VN.n29 VN.n1 0.189894
R953 VDD2.n2 VDD2.n1 80.0258
R954 VDD2.n2 VDD2.n0 80.0258
R955 VDD2 VDD2.n5 80.0229
R956 VDD2.n4 VDD2.n3 78.5813
R957 VDD2.n4 VDD2.n2 46.5429
R958 VDD2.n5 VDD2.t3 3.00466
R959 VDD2.n5 VDD2.t5 3.00466
R960 VDD2.n3 VDD2.t2 3.00466
R961 VDD2.n3 VDD2.t1 3.00466
R962 VDD2.n1 VDD2.t4 3.00466
R963 VDD2.n1 VDD2.t6 3.00466
R964 VDD2.n0 VDD2.t7 3.00466
R965 VDD2.n0 VDD2.t0 3.00466
R966 VDD2 VDD2.n4 1.55869
R967 B.n433 B.n432 585
R968 B.n431 B.n140 585
R969 B.n430 B.n429 585
R970 B.n428 B.n141 585
R971 B.n427 B.n426 585
R972 B.n425 B.n142 585
R973 B.n424 B.n423 585
R974 B.n422 B.n143 585
R975 B.n421 B.n420 585
R976 B.n419 B.n144 585
R977 B.n418 B.n417 585
R978 B.n416 B.n145 585
R979 B.n415 B.n414 585
R980 B.n413 B.n146 585
R981 B.n412 B.n411 585
R982 B.n410 B.n147 585
R983 B.n409 B.n408 585
R984 B.n407 B.n148 585
R985 B.n406 B.n405 585
R986 B.n404 B.n149 585
R987 B.n403 B.n402 585
R988 B.n401 B.n150 585
R989 B.n400 B.n399 585
R990 B.n398 B.n151 585
R991 B.n397 B.n396 585
R992 B.n395 B.n152 585
R993 B.n394 B.n393 585
R994 B.n392 B.n153 585
R995 B.n391 B.n390 585
R996 B.n389 B.n154 585
R997 B.n388 B.n387 585
R998 B.n386 B.n155 585
R999 B.n385 B.n384 585
R1000 B.n383 B.n156 585
R1001 B.n382 B.n381 585
R1002 B.n380 B.n157 585
R1003 B.n379 B.n378 585
R1004 B.n377 B.n158 585
R1005 B.n375 B.n374 585
R1006 B.n373 B.n161 585
R1007 B.n372 B.n371 585
R1008 B.n370 B.n162 585
R1009 B.n369 B.n368 585
R1010 B.n367 B.n163 585
R1011 B.n366 B.n365 585
R1012 B.n364 B.n164 585
R1013 B.n363 B.n362 585
R1014 B.n361 B.n165 585
R1015 B.n360 B.n359 585
R1016 B.n355 B.n166 585
R1017 B.n354 B.n353 585
R1018 B.n352 B.n167 585
R1019 B.n351 B.n350 585
R1020 B.n349 B.n168 585
R1021 B.n348 B.n347 585
R1022 B.n346 B.n169 585
R1023 B.n345 B.n344 585
R1024 B.n343 B.n170 585
R1025 B.n342 B.n341 585
R1026 B.n340 B.n171 585
R1027 B.n339 B.n338 585
R1028 B.n337 B.n172 585
R1029 B.n336 B.n335 585
R1030 B.n334 B.n173 585
R1031 B.n333 B.n332 585
R1032 B.n331 B.n174 585
R1033 B.n330 B.n329 585
R1034 B.n328 B.n175 585
R1035 B.n327 B.n326 585
R1036 B.n325 B.n176 585
R1037 B.n324 B.n323 585
R1038 B.n322 B.n177 585
R1039 B.n321 B.n320 585
R1040 B.n319 B.n178 585
R1041 B.n318 B.n317 585
R1042 B.n316 B.n179 585
R1043 B.n315 B.n314 585
R1044 B.n313 B.n180 585
R1045 B.n312 B.n311 585
R1046 B.n310 B.n181 585
R1047 B.n309 B.n308 585
R1048 B.n307 B.n182 585
R1049 B.n306 B.n305 585
R1050 B.n304 B.n183 585
R1051 B.n303 B.n302 585
R1052 B.n301 B.n184 585
R1053 B.n434 B.n139 585
R1054 B.n436 B.n435 585
R1055 B.n437 B.n138 585
R1056 B.n439 B.n438 585
R1057 B.n440 B.n137 585
R1058 B.n442 B.n441 585
R1059 B.n443 B.n136 585
R1060 B.n445 B.n444 585
R1061 B.n446 B.n135 585
R1062 B.n448 B.n447 585
R1063 B.n449 B.n134 585
R1064 B.n451 B.n450 585
R1065 B.n452 B.n133 585
R1066 B.n454 B.n453 585
R1067 B.n455 B.n132 585
R1068 B.n457 B.n456 585
R1069 B.n458 B.n131 585
R1070 B.n460 B.n459 585
R1071 B.n461 B.n130 585
R1072 B.n463 B.n462 585
R1073 B.n464 B.n129 585
R1074 B.n466 B.n465 585
R1075 B.n467 B.n128 585
R1076 B.n469 B.n468 585
R1077 B.n470 B.n127 585
R1078 B.n472 B.n471 585
R1079 B.n473 B.n126 585
R1080 B.n475 B.n474 585
R1081 B.n476 B.n125 585
R1082 B.n478 B.n477 585
R1083 B.n479 B.n124 585
R1084 B.n481 B.n480 585
R1085 B.n482 B.n123 585
R1086 B.n484 B.n483 585
R1087 B.n485 B.n122 585
R1088 B.n487 B.n486 585
R1089 B.n488 B.n121 585
R1090 B.n490 B.n489 585
R1091 B.n491 B.n120 585
R1092 B.n493 B.n492 585
R1093 B.n494 B.n119 585
R1094 B.n496 B.n495 585
R1095 B.n497 B.n118 585
R1096 B.n499 B.n498 585
R1097 B.n500 B.n117 585
R1098 B.n502 B.n501 585
R1099 B.n503 B.n116 585
R1100 B.n505 B.n504 585
R1101 B.n506 B.n115 585
R1102 B.n508 B.n507 585
R1103 B.n509 B.n114 585
R1104 B.n511 B.n510 585
R1105 B.n512 B.n113 585
R1106 B.n514 B.n513 585
R1107 B.n515 B.n112 585
R1108 B.n517 B.n516 585
R1109 B.n518 B.n111 585
R1110 B.n520 B.n519 585
R1111 B.n521 B.n110 585
R1112 B.n523 B.n522 585
R1113 B.n524 B.n109 585
R1114 B.n526 B.n525 585
R1115 B.n527 B.n108 585
R1116 B.n529 B.n528 585
R1117 B.n530 B.n107 585
R1118 B.n532 B.n531 585
R1119 B.n533 B.n106 585
R1120 B.n535 B.n534 585
R1121 B.n536 B.n105 585
R1122 B.n538 B.n537 585
R1123 B.n539 B.n104 585
R1124 B.n541 B.n540 585
R1125 B.n542 B.n103 585
R1126 B.n544 B.n543 585
R1127 B.n545 B.n102 585
R1128 B.n547 B.n546 585
R1129 B.n548 B.n101 585
R1130 B.n550 B.n549 585
R1131 B.n551 B.n100 585
R1132 B.n553 B.n552 585
R1133 B.n554 B.n99 585
R1134 B.n556 B.n555 585
R1135 B.n557 B.n98 585
R1136 B.n559 B.n558 585
R1137 B.n560 B.n97 585
R1138 B.n562 B.n561 585
R1139 B.n563 B.n96 585
R1140 B.n565 B.n564 585
R1141 B.n566 B.n95 585
R1142 B.n568 B.n567 585
R1143 B.n569 B.n94 585
R1144 B.n571 B.n570 585
R1145 B.n572 B.n93 585
R1146 B.n574 B.n573 585
R1147 B.n575 B.n92 585
R1148 B.n577 B.n576 585
R1149 B.n578 B.n91 585
R1150 B.n580 B.n579 585
R1151 B.n581 B.n90 585
R1152 B.n583 B.n582 585
R1153 B.n584 B.n89 585
R1154 B.n586 B.n585 585
R1155 B.n587 B.n88 585
R1156 B.n589 B.n588 585
R1157 B.n590 B.n87 585
R1158 B.n592 B.n591 585
R1159 B.n593 B.n86 585
R1160 B.n595 B.n594 585
R1161 B.n596 B.n85 585
R1162 B.n598 B.n597 585
R1163 B.n599 B.n84 585
R1164 B.n601 B.n600 585
R1165 B.n602 B.n83 585
R1166 B.n604 B.n603 585
R1167 B.n605 B.n82 585
R1168 B.n607 B.n606 585
R1169 B.n608 B.n81 585
R1170 B.n610 B.n609 585
R1171 B.n611 B.n80 585
R1172 B.n613 B.n612 585
R1173 B.n743 B.n742 585
R1174 B.n741 B.n32 585
R1175 B.n740 B.n739 585
R1176 B.n738 B.n33 585
R1177 B.n737 B.n736 585
R1178 B.n735 B.n34 585
R1179 B.n734 B.n733 585
R1180 B.n732 B.n35 585
R1181 B.n731 B.n730 585
R1182 B.n729 B.n36 585
R1183 B.n728 B.n727 585
R1184 B.n726 B.n37 585
R1185 B.n725 B.n724 585
R1186 B.n723 B.n38 585
R1187 B.n722 B.n721 585
R1188 B.n720 B.n39 585
R1189 B.n719 B.n718 585
R1190 B.n717 B.n40 585
R1191 B.n716 B.n715 585
R1192 B.n714 B.n41 585
R1193 B.n713 B.n712 585
R1194 B.n711 B.n42 585
R1195 B.n710 B.n709 585
R1196 B.n708 B.n43 585
R1197 B.n707 B.n706 585
R1198 B.n705 B.n44 585
R1199 B.n704 B.n703 585
R1200 B.n702 B.n45 585
R1201 B.n701 B.n700 585
R1202 B.n699 B.n46 585
R1203 B.n698 B.n697 585
R1204 B.n696 B.n47 585
R1205 B.n695 B.n694 585
R1206 B.n693 B.n48 585
R1207 B.n692 B.n691 585
R1208 B.n690 B.n49 585
R1209 B.n689 B.n688 585
R1210 B.n687 B.n50 585
R1211 B.n686 B.n685 585
R1212 B.n684 B.n51 585
R1213 B.n683 B.n682 585
R1214 B.n681 B.n55 585
R1215 B.n680 B.n679 585
R1216 B.n678 B.n56 585
R1217 B.n677 B.n676 585
R1218 B.n675 B.n57 585
R1219 B.n674 B.n673 585
R1220 B.n672 B.n58 585
R1221 B.n670 B.n669 585
R1222 B.n668 B.n61 585
R1223 B.n667 B.n666 585
R1224 B.n665 B.n62 585
R1225 B.n664 B.n663 585
R1226 B.n662 B.n63 585
R1227 B.n661 B.n660 585
R1228 B.n659 B.n64 585
R1229 B.n658 B.n657 585
R1230 B.n656 B.n65 585
R1231 B.n655 B.n654 585
R1232 B.n653 B.n66 585
R1233 B.n652 B.n651 585
R1234 B.n650 B.n67 585
R1235 B.n649 B.n648 585
R1236 B.n647 B.n68 585
R1237 B.n646 B.n645 585
R1238 B.n644 B.n69 585
R1239 B.n643 B.n642 585
R1240 B.n641 B.n70 585
R1241 B.n640 B.n639 585
R1242 B.n638 B.n71 585
R1243 B.n637 B.n636 585
R1244 B.n635 B.n72 585
R1245 B.n634 B.n633 585
R1246 B.n632 B.n73 585
R1247 B.n631 B.n630 585
R1248 B.n629 B.n74 585
R1249 B.n628 B.n627 585
R1250 B.n626 B.n75 585
R1251 B.n625 B.n624 585
R1252 B.n623 B.n76 585
R1253 B.n622 B.n621 585
R1254 B.n620 B.n77 585
R1255 B.n619 B.n618 585
R1256 B.n617 B.n78 585
R1257 B.n616 B.n615 585
R1258 B.n614 B.n79 585
R1259 B.n744 B.n31 585
R1260 B.n746 B.n745 585
R1261 B.n747 B.n30 585
R1262 B.n749 B.n748 585
R1263 B.n750 B.n29 585
R1264 B.n752 B.n751 585
R1265 B.n753 B.n28 585
R1266 B.n755 B.n754 585
R1267 B.n756 B.n27 585
R1268 B.n758 B.n757 585
R1269 B.n759 B.n26 585
R1270 B.n761 B.n760 585
R1271 B.n762 B.n25 585
R1272 B.n764 B.n763 585
R1273 B.n765 B.n24 585
R1274 B.n767 B.n766 585
R1275 B.n768 B.n23 585
R1276 B.n770 B.n769 585
R1277 B.n771 B.n22 585
R1278 B.n773 B.n772 585
R1279 B.n774 B.n21 585
R1280 B.n776 B.n775 585
R1281 B.n777 B.n20 585
R1282 B.n779 B.n778 585
R1283 B.n780 B.n19 585
R1284 B.n782 B.n781 585
R1285 B.n783 B.n18 585
R1286 B.n785 B.n784 585
R1287 B.n786 B.n17 585
R1288 B.n788 B.n787 585
R1289 B.n789 B.n16 585
R1290 B.n791 B.n790 585
R1291 B.n792 B.n15 585
R1292 B.n794 B.n793 585
R1293 B.n795 B.n14 585
R1294 B.n797 B.n796 585
R1295 B.n798 B.n13 585
R1296 B.n800 B.n799 585
R1297 B.n801 B.n12 585
R1298 B.n803 B.n802 585
R1299 B.n804 B.n11 585
R1300 B.n806 B.n805 585
R1301 B.n807 B.n10 585
R1302 B.n809 B.n808 585
R1303 B.n810 B.n9 585
R1304 B.n812 B.n811 585
R1305 B.n813 B.n8 585
R1306 B.n815 B.n814 585
R1307 B.n816 B.n7 585
R1308 B.n818 B.n817 585
R1309 B.n819 B.n6 585
R1310 B.n821 B.n820 585
R1311 B.n822 B.n5 585
R1312 B.n824 B.n823 585
R1313 B.n825 B.n4 585
R1314 B.n827 B.n826 585
R1315 B.n828 B.n3 585
R1316 B.n830 B.n829 585
R1317 B.n831 B.n0 585
R1318 B.n2 B.n1 585
R1319 B.n214 B.n213 585
R1320 B.n216 B.n215 585
R1321 B.n217 B.n212 585
R1322 B.n219 B.n218 585
R1323 B.n220 B.n211 585
R1324 B.n222 B.n221 585
R1325 B.n223 B.n210 585
R1326 B.n225 B.n224 585
R1327 B.n226 B.n209 585
R1328 B.n228 B.n227 585
R1329 B.n229 B.n208 585
R1330 B.n231 B.n230 585
R1331 B.n232 B.n207 585
R1332 B.n234 B.n233 585
R1333 B.n235 B.n206 585
R1334 B.n237 B.n236 585
R1335 B.n238 B.n205 585
R1336 B.n240 B.n239 585
R1337 B.n241 B.n204 585
R1338 B.n243 B.n242 585
R1339 B.n244 B.n203 585
R1340 B.n246 B.n245 585
R1341 B.n247 B.n202 585
R1342 B.n249 B.n248 585
R1343 B.n250 B.n201 585
R1344 B.n252 B.n251 585
R1345 B.n253 B.n200 585
R1346 B.n255 B.n254 585
R1347 B.n256 B.n199 585
R1348 B.n258 B.n257 585
R1349 B.n259 B.n198 585
R1350 B.n261 B.n260 585
R1351 B.n262 B.n197 585
R1352 B.n264 B.n263 585
R1353 B.n265 B.n196 585
R1354 B.n267 B.n266 585
R1355 B.n268 B.n195 585
R1356 B.n270 B.n269 585
R1357 B.n271 B.n194 585
R1358 B.n273 B.n272 585
R1359 B.n274 B.n193 585
R1360 B.n276 B.n275 585
R1361 B.n277 B.n192 585
R1362 B.n279 B.n278 585
R1363 B.n280 B.n191 585
R1364 B.n282 B.n281 585
R1365 B.n283 B.n190 585
R1366 B.n285 B.n284 585
R1367 B.n286 B.n189 585
R1368 B.n288 B.n287 585
R1369 B.n289 B.n188 585
R1370 B.n291 B.n290 585
R1371 B.n292 B.n187 585
R1372 B.n294 B.n293 585
R1373 B.n295 B.n186 585
R1374 B.n297 B.n296 585
R1375 B.n298 B.n185 585
R1376 B.n300 B.n299 585
R1377 B.n299 B.n184 454.062
R1378 B.n434 B.n433 454.062
R1379 B.n614 B.n613 454.062
R1380 B.n742 B.n31 454.062
R1381 B.n159 B.t1 422.022
R1382 B.n59 B.t8 422.022
R1383 B.n356 B.t4 422.022
R1384 B.n52 B.t11 422.022
R1385 B.n160 B.t2 354.531
R1386 B.n60 B.t7 354.531
R1387 B.n357 B.t5 354.531
R1388 B.n53 B.t10 354.531
R1389 B.n356 B.t3 291.531
R1390 B.n159 B.t0 291.531
R1391 B.n59 B.t6 291.531
R1392 B.n52 B.t9 291.531
R1393 B.n833 B.n832 256.663
R1394 B.n832 B.n831 235.042
R1395 B.n832 B.n2 235.042
R1396 B.n303 B.n184 163.367
R1397 B.n304 B.n303 163.367
R1398 B.n305 B.n304 163.367
R1399 B.n305 B.n182 163.367
R1400 B.n309 B.n182 163.367
R1401 B.n310 B.n309 163.367
R1402 B.n311 B.n310 163.367
R1403 B.n311 B.n180 163.367
R1404 B.n315 B.n180 163.367
R1405 B.n316 B.n315 163.367
R1406 B.n317 B.n316 163.367
R1407 B.n317 B.n178 163.367
R1408 B.n321 B.n178 163.367
R1409 B.n322 B.n321 163.367
R1410 B.n323 B.n322 163.367
R1411 B.n323 B.n176 163.367
R1412 B.n327 B.n176 163.367
R1413 B.n328 B.n327 163.367
R1414 B.n329 B.n328 163.367
R1415 B.n329 B.n174 163.367
R1416 B.n333 B.n174 163.367
R1417 B.n334 B.n333 163.367
R1418 B.n335 B.n334 163.367
R1419 B.n335 B.n172 163.367
R1420 B.n339 B.n172 163.367
R1421 B.n340 B.n339 163.367
R1422 B.n341 B.n340 163.367
R1423 B.n341 B.n170 163.367
R1424 B.n345 B.n170 163.367
R1425 B.n346 B.n345 163.367
R1426 B.n347 B.n346 163.367
R1427 B.n347 B.n168 163.367
R1428 B.n351 B.n168 163.367
R1429 B.n352 B.n351 163.367
R1430 B.n353 B.n352 163.367
R1431 B.n353 B.n166 163.367
R1432 B.n360 B.n166 163.367
R1433 B.n361 B.n360 163.367
R1434 B.n362 B.n361 163.367
R1435 B.n362 B.n164 163.367
R1436 B.n366 B.n164 163.367
R1437 B.n367 B.n366 163.367
R1438 B.n368 B.n367 163.367
R1439 B.n368 B.n162 163.367
R1440 B.n372 B.n162 163.367
R1441 B.n373 B.n372 163.367
R1442 B.n374 B.n373 163.367
R1443 B.n374 B.n158 163.367
R1444 B.n379 B.n158 163.367
R1445 B.n380 B.n379 163.367
R1446 B.n381 B.n380 163.367
R1447 B.n381 B.n156 163.367
R1448 B.n385 B.n156 163.367
R1449 B.n386 B.n385 163.367
R1450 B.n387 B.n386 163.367
R1451 B.n387 B.n154 163.367
R1452 B.n391 B.n154 163.367
R1453 B.n392 B.n391 163.367
R1454 B.n393 B.n392 163.367
R1455 B.n393 B.n152 163.367
R1456 B.n397 B.n152 163.367
R1457 B.n398 B.n397 163.367
R1458 B.n399 B.n398 163.367
R1459 B.n399 B.n150 163.367
R1460 B.n403 B.n150 163.367
R1461 B.n404 B.n403 163.367
R1462 B.n405 B.n404 163.367
R1463 B.n405 B.n148 163.367
R1464 B.n409 B.n148 163.367
R1465 B.n410 B.n409 163.367
R1466 B.n411 B.n410 163.367
R1467 B.n411 B.n146 163.367
R1468 B.n415 B.n146 163.367
R1469 B.n416 B.n415 163.367
R1470 B.n417 B.n416 163.367
R1471 B.n417 B.n144 163.367
R1472 B.n421 B.n144 163.367
R1473 B.n422 B.n421 163.367
R1474 B.n423 B.n422 163.367
R1475 B.n423 B.n142 163.367
R1476 B.n427 B.n142 163.367
R1477 B.n428 B.n427 163.367
R1478 B.n429 B.n428 163.367
R1479 B.n429 B.n140 163.367
R1480 B.n433 B.n140 163.367
R1481 B.n613 B.n80 163.367
R1482 B.n609 B.n80 163.367
R1483 B.n609 B.n608 163.367
R1484 B.n608 B.n607 163.367
R1485 B.n607 B.n82 163.367
R1486 B.n603 B.n82 163.367
R1487 B.n603 B.n602 163.367
R1488 B.n602 B.n601 163.367
R1489 B.n601 B.n84 163.367
R1490 B.n597 B.n84 163.367
R1491 B.n597 B.n596 163.367
R1492 B.n596 B.n595 163.367
R1493 B.n595 B.n86 163.367
R1494 B.n591 B.n86 163.367
R1495 B.n591 B.n590 163.367
R1496 B.n590 B.n589 163.367
R1497 B.n589 B.n88 163.367
R1498 B.n585 B.n88 163.367
R1499 B.n585 B.n584 163.367
R1500 B.n584 B.n583 163.367
R1501 B.n583 B.n90 163.367
R1502 B.n579 B.n90 163.367
R1503 B.n579 B.n578 163.367
R1504 B.n578 B.n577 163.367
R1505 B.n577 B.n92 163.367
R1506 B.n573 B.n92 163.367
R1507 B.n573 B.n572 163.367
R1508 B.n572 B.n571 163.367
R1509 B.n571 B.n94 163.367
R1510 B.n567 B.n94 163.367
R1511 B.n567 B.n566 163.367
R1512 B.n566 B.n565 163.367
R1513 B.n565 B.n96 163.367
R1514 B.n561 B.n96 163.367
R1515 B.n561 B.n560 163.367
R1516 B.n560 B.n559 163.367
R1517 B.n559 B.n98 163.367
R1518 B.n555 B.n98 163.367
R1519 B.n555 B.n554 163.367
R1520 B.n554 B.n553 163.367
R1521 B.n553 B.n100 163.367
R1522 B.n549 B.n100 163.367
R1523 B.n549 B.n548 163.367
R1524 B.n548 B.n547 163.367
R1525 B.n547 B.n102 163.367
R1526 B.n543 B.n102 163.367
R1527 B.n543 B.n542 163.367
R1528 B.n542 B.n541 163.367
R1529 B.n541 B.n104 163.367
R1530 B.n537 B.n104 163.367
R1531 B.n537 B.n536 163.367
R1532 B.n536 B.n535 163.367
R1533 B.n535 B.n106 163.367
R1534 B.n531 B.n106 163.367
R1535 B.n531 B.n530 163.367
R1536 B.n530 B.n529 163.367
R1537 B.n529 B.n108 163.367
R1538 B.n525 B.n108 163.367
R1539 B.n525 B.n524 163.367
R1540 B.n524 B.n523 163.367
R1541 B.n523 B.n110 163.367
R1542 B.n519 B.n110 163.367
R1543 B.n519 B.n518 163.367
R1544 B.n518 B.n517 163.367
R1545 B.n517 B.n112 163.367
R1546 B.n513 B.n112 163.367
R1547 B.n513 B.n512 163.367
R1548 B.n512 B.n511 163.367
R1549 B.n511 B.n114 163.367
R1550 B.n507 B.n114 163.367
R1551 B.n507 B.n506 163.367
R1552 B.n506 B.n505 163.367
R1553 B.n505 B.n116 163.367
R1554 B.n501 B.n116 163.367
R1555 B.n501 B.n500 163.367
R1556 B.n500 B.n499 163.367
R1557 B.n499 B.n118 163.367
R1558 B.n495 B.n118 163.367
R1559 B.n495 B.n494 163.367
R1560 B.n494 B.n493 163.367
R1561 B.n493 B.n120 163.367
R1562 B.n489 B.n120 163.367
R1563 B.n489 B.n488 163.367
R1564 B.n488 B.n487 163.367
R1565 B.n487 B.n122 163.367
R1566 B.n483 B.n122 163.367
R1567 B.n483 B.n482 163.367
R1568 B.n482 B.n481 163.367
R1569 B.n481 B.n124 163.367
R1570 B.n477 B.n124 163.367
R1571 B.n477 B.n476 163.367
R1572 B.n476 B.n475 163.367
R1573 B.n475 B.n126 163.367
R1574 B.n471 B.n126 163.367
R1575 B.n471 B.n470 163.367
R1576 B.n470 B.n469 163.367
R1577 B.n469 B.n128 163.367
R1578 B.n465 B.n128 163.367
R1579 B.n465 B.n464 163.367
R1580 B.n464 B.n463 163.367
R1581 B.n463 B.n130 163.367
R1582 B.n459 B.n130 163.367
R1583 B.n459 B.n458 163.367
R1584 B.n458 B.n457 163.367
R1585 B.n457 B.n132 163.367
R1586 B.n453 B.n132 163.367
R1587 B.n453 B.n452 163.367
R1588 B.n452 B.n451 163.367
R1589 B.n451 B.n134 163.367
R1590 B.n447 B.n134 163.367
R1591 B.n447 B.n446 163.367
R1592 B.n446 B.n445 163.367
R1593 B.n445 B.n136 163.367
R1594 B.n441 B.n136 163.367
R1595 B.n441 B.n440 163.367
R1596 B.n440 B.n439 163.367
R1597 B.n439 B.n138 163.367
R1598 B.n435 B.n138 163.367
R1599 B.n435 B.n434 163.367
R1600 B.n742 B.n741 163.367
R1601 B.n741 B.n740 163.367
R1602 B.n740 B.n33 163.367
R1603 B.n736 B.n33 163.367
R1604 B.n736 B.n735 163.367
R1605 B.n735 B.n734 163.367
R1606 B.n734 B.n35 163.367
R1607 B.n730 B.n35 163.367
R1608 B.n730 B.n729 163.367
R1609 B.n729 B.n728 163.367
R1610 B.n728 B.n37 163.367
R1611 B.n724 B.n37 163.367
R1612 B.n724 B.n723 163.367
R1613 B.n723 B.n722 163.367
R1614 B.n722 B.n39 163.367
R1615 B.n718 B.n39 163.367
R1616 B.n718 B.n717 163.367
R1617 B.n717 B.n716 163.367
R1618 B.n716 B.n41 163.367
R1619 B.n712 B.n41 163.367
R1620 B.n712 B.n711 163.367
R1621 B.n711 B.n710 163.367
R1622 B.n710 B.n43 163.367
R1623 B.n706 B.n43 163.367
R1624 B.n706 B.n705 163.367
R1625 B.n705 B.n704 163.367
R1626 B.n704 B.n45 163.367
R1627 B.n700 B.n45 163.367
R1628 B.n700 B.n699 163.367
R1629 B.n699 B.n698 163.367
R1630 B.n698 B.n47 163.367
R1631 B.n694 B.n47 163.367
R1632 B.n694 B.n693 163.367
R1633 B.n693 B.n692 163.367
R1634 B.n692 B.n49 163.367
R1635 B.n688 B.n49 163.367
R1636 B.n688 B.n687 163.367
R1637 B.n687 B.n686 163.367
R1638 B.n686 B.n51 163.367
R1639 B.n682 B.n51 163.367
R1640 B.n682 B.n681 163.367
R1641 B.n681 B.n680 163.367
R1642 B.n680 B.n56 163.367
R1643 B.n676 B.n56 163.367
R1644 B.n676 B.n675 163.367
R1645 B.n675 B.n674 163.367
R1646 B.n674 B.n58 163.367
R1647 B.n669 B.n58 163.367
R1648 B.n669 B.n668 163.367
R1649 B.n668 B.n667 163.367
R1650 B.n667 B.n62 163.367
R1651 B.n663 B.n62 163.367
R1652 B.n663 B.n662 163.367
R1653 B.n662 B.n661 163.367
R1654 B.n661 B.n64 163.367
R1655 B.n657 B.n64 163.367
R1656 B.n657 B.n656 163.367
R1657 B.n656 B.n655 163.367
R1658 B.n655 B.n66 163.367
R1659 B.n651 B.n66 163.367
R1660 B.n651 B.n650 163.367
R1661 B.n650 B.n649 163.367
R1662 B.n649 B.n68 163.367
R1663 B.n645 B.n68 163.367
R1664 B.n645 B.n644 163.367
R1665 B.n644 B.n643 163.367
R1666 B.n643 B.n70 163.367
R1667 B.n639 B.n70 163.367
R1668 B.n639 B.n638 163.367
R1669 B.n638 B.n637 163.367
R1670 B.n637 B.n72 163.367
R1671 B.n633 B.n72 163.367
R1672 B.n633 B.n632 163.367
R1673 B.n632 B.n631 163.367
R1674 B.n631 B.n74 163.367
R1675 B.n627 B.n74 163.367
R1676 B.n627 B.n626 163.367
R1677 B.n626 B.n625 163.367
R1678 B.n625 B.n76 163.367
R1679 B.n621 B.n76 163.367
R1680 B.n621 B.n620 163.367
R1681 B.n620 B.n619 163.367
R1682 B.n619 B.n78 163.367
R1683 B.n615 B.n78 163.367
R1684 B.n615 B.n614 163.367
R1685 B.n746 B.n31 163.367
R1686 B.n747 B.n746 163.367
R1687 B.n748 B.n747 163.367
R1688 B.n748 B.n29 163.367
R1689 B.n752 B.n29 163.367
R1690 B.n753 B.n752 163.367
R1691 B.n754 B.n753 163.367
R1692 B.n754 B.n27 163.367
R1693 B.n758 B.n27 163.367
R1694 B.n759 B.n758 163.367
R1695 B.n760 B.n759 163.367
R1696 B.n760 B.n25 163.367
R1697 B.n764 B.n25 163.367
R1698 B.n765 B.n764 163.367
R1699 B.n766 B.n765 163.367
R1700 B.n766 B.n23 163.367
R1701 B.n770 B.n23 163.367
R1702 B.n771 B.n770 163.367
R1703 B.n772 B.n771 163.367
R1704 B.n772 B.n21 163.367
R1705 B.n776 B.n21 163.367
R1706 B.n777 B.n776 163.367
R1707 B.n778 B.n777 163.367
R1708 B.n778 B.n19 163.367
R1709 B.n782 B.n19 163.367
R1710 B.n783 B.n782 163.367
R1711 B.n784 B.n783 163.367
R1712 B.n784 B.n17 163.367
R1713 B.n788 B.n17 163.367
R1714 B.n789 B.n788 163.367
R1715 B.n790 B.n789 163.367
R1716 B.n790 B.n15 163.367
R1717 B.n794 B.n15 163.367
R1718 B.n795 B.n794 163.367
R1719 B.n796 B.n795 163.367
R1720 B.n796 B.n13 163.367
R1721 B.n800 B.n13 163.367
R1722 B.n801 B.n800 163.367
R1723 B.n802 B.n801 163.367
R1724 B.n802 B.n11 163.367
R1725 B.n806 B.n11 163.367
R1726 B.n807 B.n806 163.367
R1727 B.n808 B.n807 163.367
R1728 B.n808 B.n9 163.367
R1729 B.n812 B.n9 163.367
R1730 B.n813 B.n812 163.367
R1731 B.n814 B.n813 163.367
R1732 B.n814 B.n7 163.367
R1733 B.n818 B.n7 163.367
R1734 B.n819 B.n818 163.367
R1735 B.n820 B.n819 163.367
R1736 B.n820 B.n5 163.367
R1737 B.n824 B.n5 163.367
R1738 B.n825 B.n824 163.367
R1739 B.n826 B.n825 163.367
R1740 B.n826 B.n3 163.367
R1741 B.n830 B.n3 163.367
R1742 B.n831 B.n830 163.367
R1743 B.n214 B.n2 163.367
R1744 B.n215 B.n214 163.367
R1745 B.n215 B.n212 163.367
R1746 B.n219 B.n212 163.367
R1747 B.n220 B.n219 163.367
R1748 B.n221 B.n220 163.367
R1749 B.n221 B.n210 163.367
R1750 B.n225 B.n210 163.367
R1751 B.n226 B.n225 163.367
R1752 B.n227 B.n226 163.367
R1753 B.n227 B.n208 163.367
R1754 B.n231 B.n208 163.367
R1755 B.n232 B.n231 163.367
R1756 B.n233 B.n232 163.367
R1757 B.n233 B.n206 163.367
R1758 B.n237 B.n206 163.367
R1759 B.n238 B.n237 163.367
R1760 B.n239 B.n238 163.367
R1761 B.n239 B.n204 163.367
R1762 B.n243 B.n204 163.367
R1763 B.n244 B.n243 163.367
R1764 B.n245 B.n244 163.367
R1765 B.n245 B.n202 163.367
R1766 B.n249 B.n202 163.367
R1767 B.n250 B.n249 163.367
R1768 B.n251 B.n250 163.367
R1769 B.n251 B.n200 163.367
R1770 B.n255 B.n200 163.367
R1771 B.n256 B.n255 163.367
R1772 B.n257 B.n256 163.367
R1773 B.n257 B.n198 163.367
R1774 B.n261 B.n198 163.367
R1775 B.n262 B.n261 163.367
R1776 B.n263 B.n262 163.367
R1777 B.n263 B.n196 163.367
R1778 B.n267 B.n196 163.367
R1779 B.n268 B.n267 163.367
R1780 B.n269 B.n268 163.367
R1781 B.n269 B.n194 163.367
R1782 B.n273 B.n194 163.367
R1783 B.n274 B.n273 163.367
R1784 B.n275 B.n274 163.367
R1785 B.n275 B.n192 163.367
R1786 B.n279 B.n192 163.367
R1787 B.n280 B.n279 163.367
R1788 B.n281 B.n280 163.367
R1789 B.n281 B.n190 163.367
R1790 B.n285 B.n190 163.367
R1791 B.n286 B.n285 163.367
R1792 B.n287 B.n286 163.367
R1793 B.n287 B.n188 163.367
R1794 B.n291 B.n188 163.367
R1795 B.n292 B.n291 163.367
R1796 B.n293 B.n292 163.367
R1797 B.n293 B.n186 163.367
R1798 B.n297 B.n186 163.367
R1799 B.n298 B.n297 163.367
R1800 B.n299 B.n298 163.367
R1801 B.n357 B.n356 67.4914
R1802 B.n160 B.n159 67.4914
R1803 B.n60 B.n59 67.4914
R1804 B.n53 B.n52 67.4914
R1805 B.n358 B.n357 59.5399
R1806 B.n376 B.n160 59.5399
R1807 B.n671 B.n60 59.5399
R1808 B.n54 B.n53 59.5399
R1809 B.n744 B.n743 29.5029
R1810 B.n612 B.n79 29.5029
R1811 B.n301 B.n300 29.5029
R1812 B.n432 B.n139 29.5029
R1813 B B.n833 18.0485
R1814 B.n745 B.n744 10.6151
R1815 B.n745 B.n30 10.6151
R1816 B.n749 B.n30 10.6151
R1817 B.n750 B.n749 10.6151
R1818 B.n751 B.n750 10.6151
R1819 B.n751 B.n28 10.6151
R1820 B.n755 B.n28 10.6151
R1821 B.n756 B.n755 10.6151
R1822 B.n757 B.n756 10.6151
R1823 B.n757 B.n26 10.6151
R1824 B.n761 B.n26 10.6151
R1825 B.n762 B.n761 10.6151
R1826 B.n763 B.n762 10.6151
R1827 B.n763 B.n24 10.6151
R1828 B.n767 B.n24 10.6151
R1829 B.n768 B.n767 10.6151
R1830 B.n769 B.n768 10.6151
R1831 B.n769 B.n22 10.6151
R1832 B.n773 B.n22 10.6151
R1833 B.n774 B.n773 10.6151
R1834 B.n775 B.n774 10.6151
R1835 B.n775 B.n20 10.6151
R1836 B.n779 B.n20 10.6151
R1837 B.n780 B.n779 10.6151
R1838 B.n781 B.n780 10.6151
R1839 B.n781 B.n18 10.6151
R1840 B.n785 B.n18 10.6151
R1841 B.n786 B.n785 10.6151
R1842 B.n787 B.n786 10.6151
R1843 B.n787 B.n16 10.6151
R1844 B.n791 B.n16 10.6151
R1845 B.n792 B.n791 10.6151
R1846 B.n793 B.n792 10.6151
R1847 B.n793 B.n14 10.6151
R1848 B.n797 B.n14 10.6151
R1849 B.n798 B.n797 10.6151
R1850 B.n799 B.n798 10.6151
R1851 B.n799 B.n12 10.6151
R1852 B.n803 B.n12 10.6151
R1853 B.n804 B.n803 10.6151
R1854 B.n805 B.n804 10.6151
R1855 B.n805 B.n10 10.6151
R1856 B.n809 B.n10 10.6151
R1857 B.n810 B.n809 10.6151
R1858 B.n811 B.n810 10.6151
R1859 B.n811 B.n8 10.6151
R1860 B.n815 B.n8 10.6151
R1861 B.n816 B.n815 10.6151
R1862 B.n817 B.n816 10.6151
R1863 B.n817 B.n6 10.6151
R1864 B.n821 B.n6 10.6151
R1865 B.n822 B.n821 10.6151
R1866 B.n823 B.n822 10.6151
R1867 B.n823 B.n4 10.6151
R1868 B.n827 B.n4 10.6151
R1869 B.n828 B.n827 10.6151
R1870 B.n829 B.n828 10.6151
R1871 B.n829 B.n0 10.6151
R1872 B.n743 B.n32 10.6151
R1873 B.n739 B.n32 10.6151
R1874 B.n739 B.n738 10.6151
R1875 B.n738 B.n737 10.6151
R1876 B.n737 B.n34 10.6151
R1877 B.n733 B.n34 10.6151
R1878 B.n733 B.n732 10.6151
R1879 B.n732 B.n731 10.6151
R1880 B.n731 B.n36 10.6151
R1881 B.n727 B.n36 10.6151
R1882 B.n727 B.n726 10.6151
R1883 B.n726 B.n725 10.6151
R1884 B.n725 B.n38 10.6151
R1885 B.n721 B.n38 10.6151
R1886 B.n721 B.n720 10.6151
R1887 B.n720 B.n719 10.6151
R1888 B.n719 B.n40 10.6151
R1889 B.n715 B.n40 10.6151
R1890 B.n715 B.n714 10.6151
R1891 B.n714 B.n713 10.6151
R1892 B.n713 B.n42 10.6151
R1893 B.n709 B.n42 10.6151
R1894 B.n709 B.n708 10.6151
R1895 B.n708 B.n707 10.6151
R1896 B.n707 B.n44 10.6151
R1897 B.n703 B.n44 10.6151
R1898 B.n703 B.n702 10.6151
R1899 B.n702 B.n701 10.6151
R1900 B.n701 B.n46 10.6151
R1901 B.n697 B.n46 10.6151
R1902 B.n697 B.n696 10.6151
R1903 B.n696 B.n695 10.6151
R1904 B.n695 B.n48 10.6151
R1905 B.n691 B.n48 10.6151
R1906 B.n691 B.n690 10.6151
R1907 B.n690 B.n689 10.6151
R1908 B.n689 B.n50 10.6151
R1909 B.n685 B.n684 10.6151
R1910 B.n684 B.n683 10.6151
R1911 B.n683 B.n55 10.6151
R1912 B.n679 B.n55 10.6151
R1913 B.n679 B.n678 10.6151
R1914 B.n678 B.n677 10.6151
R1915 B.n677 B.n57 10.6151
R1916 B.n673 B.n57 10.6151
R1917 B.n673 B.n672 10.6151
R1918 B.n670 B.n61 10.6151
R1919 B.n666 B.n61 10.6151
R1920 B.n666 B.n665 10.6151
R1921 B.n665 B.n664 10.6151
R1922 B.n664 B.n63 10.6151
R1923 B.n660 B.n63 10.6151
R1924 B.n660 B.n659 10.6151
R1925 B.n659 B.n658 10.6151
R1926 B.n658 B.n65 10.6151
R1927 B.n654 B.n65 10.6151
R1928 B.n654 B.n653 10.6151
R1929 B.n653 B.n652 10.6151
R1930 B.n652 B.n67 10.6151
R1931 B.n648 B.n67 10.6151
R1932 B.n648 B.n647 10.6151
R1933 B.n647 B.n646 10.6151
R1934 B.n646 B.n69 10.6151
R1935 B.n642 B.n69 10.6151
R1936 B.n642 B.n641 10.6151
R1937 B.n641 B.n640 10.6151
R1938 B.n640 B.n71 10.6151
R1939 B.n636 B.n71 10.6151
R1940 B.n636 B.n635 10.6151
R1941 B.n635 B.n634 10.6151
R1942 B.n634 B.n73 10.6151
R1943 B.n630 B.n73 10.6151
R1944 B.n630 B.n629 10.6151
R1945 B.n629 B.n628 10.6151
R1946 B.n628 B.n75 10.6151
R1947 B.n624 B.n75 10.6151
R1948 B.n624 B.n623 10.6151
R1949 B.n623 B.n622 10.6151
R1950 B.n622 B.n77 10.6151
R1951 B.n618 B.n77 10.6151
R1952 B.n618 B.n617 10.6151
R1953 B.n617 B.n616 10.6151
R1954 B.n616 B.n79 10.6151
R1955 B.n612 B.n611 10.6151
R1956 B.n611 B.n610 10.6151
R1957 B.n610 B.n81 10.6151
R1958 B.n606 B.n81 10.6151
R1959 B.n606 B.n605 10.6151
R1960 B.n605 B.n604 10.6151
R1961 B.n604 B.n83 10.6151
R1962 B.n600 B.n83 10.6151
R1963 B.n600 B.n599 10.6151
R1964 B.n599 B.n598 10.6151
R1965 B.n598 B.n85 10.6151
R1966 B.n594 B.n85 10.6151
R1967 B.n594 B.n593 10.6151
R1968 B.n593 B.n592 10.6151
R1969 B.n592 B.n87 10.6151
R1970 B.n588 B.n87 10.6151
R1971 B.n588 B.n587 10.6151
R1972 B.n587 B.n586 10.6151
R1973 B.n586 B.n89 10.6151
R1974 B.n582 B.n89 10.6151
R1975 B.n582 B.n581 10.6151
R1976 B.n581 B.n580 10.6151
R1977 B.n580 B.n91 10.6151
R1978 B.n576 B.n91 10.6151
R1979 B.n576 B.n575 10.6151
R1980 B.n575 B.n574 10.6151
R1981 B.n574 B.n93 10.6151
R1982 B.n570 B.n93 10.6151
R1983 B.n570 B.n569 10.6151
R1984 B.n569 B.n568 10.6151
R1985 B.n568 B.n95 10.6151
R1986 B.n564 B.n95 10.6151
R1987 B.n564 B.n563 10.6151
R1988 B.n563 B.n562 10.6151
R1989 B.n562 B.n97 10.6151
R1990 B.n558 B.n97 10.6151
R1991 B.n558 B.n557 10.6151
R1992 B.n557 B.n556 10.6151
R1993 B.n556 B.n99 10.6151
R1994 B.n552 B.n99 10.6151
R1995 B.n552 B.n551 10.6151
R1996 B.n551 B.n550 10.6151
R1997 B.n550 B.n101 10.6151
R1998 B.n546 B.n101 10.6151
R1999 B.n546 B.n545 10.6151
R2000 B.n545 B.n544 10.6151
R2001 B.n544 B.n103 10.6151
R2002 B.n540 B.n103 10.6151
R2003 B.n540 B.n539 10.6151
R2004 B.n539 B.n538 10.6151
R2005 B.n538 B.n105 10.6151
R2006 B.n534 B.n105 10.6151
R2007 B.n534 B.n533 10.6151
R2008 B.n533 B.n532 10.6151
R2009 B.n532 B.n107 10.6151
R2010 B.n528 B.n107 10.6151
R2011 B.n528 B.n527 10.6151
R2012 B.n527 B.n526 10.6151
R2013 B.n526 B.n109 10.6151
R2014 B.n522 B.n109 10.6151
R2015 B.n522 B.n521 10.6151
R2016 B.n521 B.n520 10.6151
R2017 B.n520 B.n111 10.6151
R2018 B.n516 B.n111 10.6151
R2019 B.n516 B.n515 10.6151
R2020 B.n515 B.n514 10.6151
R2021 B.n514 B.n113 10.6151
R2022 B.n510 B.n113 10.6151
R2023 B.n510 B.n509 10.6151
R2024 B.n509 B.n508 10.6151
R2025 B.n508 B.n115 10.6151
R2026 B.n504 B.n115 10.6151
R2027 B.n504 B.n503 10.6151
R2028 B.n503 B.n502 10.6151
R2029 B.n502 B.n117 10.6151
R2030 B.n498 B.n117 10.6151
R2031 B.n498 B.n497 10.6151
R2032 B.n497 B.n496 10.6151
R2033 B.n496 B.n119 10.6151
R2034 B.n492 B.n119 10.6151
R2035 B.n492 B.n491 10.6151
R2036 B.n491 B.n490 10.6151
R2037 B.n490 B.n121 10.6151
R2038 B.n486 B.n121 10.6151
R2039 B.n486 B.n485 10.6151
R2040 B.n485 B.n484 10.6151
R2041 B.n484 B.n123 10.6151
R2042 B.n480 B.n123 10.6151
R2043 B.n480 B.n479 10.6151
R2044 B.n479 B.n478 10.6151
R2045 B.n478 B.n125 10.6151
R2046 B.n474 B.n125 10.6151
R2047 B.n474 B.n473 10.6151
R2048 B.n473 B.n472 10.6151
R2049 B.n472 B.n127 10.6151
R2050 B.n468 B.n127 10.6151
R2051 B.n468 B.n467 10.6151
R2052 B.n467 B.n466 10.6151
R2053 B.n466 B.n129 10.6151
R2054 B.n462 B.n129 10.6151
R2055 B.n462 B.n461 10.6151
R2056 B.n461 B.n460 10.6151
R2057 B.n460 B.n131 10.6151
R2058 B.n456 B.n131 10.6151
R2059 B.n456 B.n455 10.6151
R2060 B.n455 B.n454 10.6151
R2061 B.n454 B.n133 10.6151
R2062 B.n450 B.n133 10.6151
R2063 B.n450 B.n449 10.6151
R2064 B.n449 B.n448 10.6151
R2065 B.n448 B.n135 10.6151
R2066 B.n444 B.n135 10.6151
R2067 B.n444 B.n443 10.6151
R2068 B.n443 B.n442 10.6151
R2069 B.n442 B.n137 10.6151
R2070 B.n438 B.n137 10.6151
R2071 B.n438 B.n437 10.6151
R2072 B.n437 B.n436 10.6151
R2073 B.n436 B.n139 10.6151
R2074 B.n213 B.n1 10.6151
R2075 B.n216 B.n213 10.6151
R2076 B.n217 B.n216 10.6151
R2077 B.n218 B.n217 10.6151
R2078 B.n218 B.n211 10.6151
R2079 B.n222 B.n211 10.6151
R2080 B.n223 B.n222 10.6151
R2081 B.n224 B.n223 10.6151
R2082 B.n224 B.n209 10.6151
R2083 B.n228 B.n209 10.6151
R2084 B.n229 B.n228 10.6151
R2085 B.n230 B.n229 10.6151
R2086 B.n230 B.n207 10.6151
R2087 B.n234 B.n207 10.6151
R2088 B.n235 B.n234 10.6151
R2089 B.n236 B.n235 10.6151
R2090 B.n236 B.n205 10.6151
R2091 B.n240 B.n205 10.6151
R2092 B.n241 B.n240 10.6151
R2093 B.n242 B.n241 10.6151
R2094 B.n242 B.n203 10.6151
R2095 B.n246 B.n203 10.6151
R2096 B.n247 B.n246 10.6151
R2097 B.n248 B.n247 10.6151
R2098 B.n248 B.n201 10.6151
R2099 B.n252 B.n201 10.6151
R2100 B.n253 B.n252 10.6151
R2101 B.n254 B.n253 10.6151
R2102 B.n254 B.n199 10.6151
R2103 B.n258 B.n199 10.6151
R2104 B.n259 B.n258 10.6151
R2105 B.n260 B.n259 10.6151
R2106 B.n260 B.n197 10.6151
R2107 B.n264 B.n197 10.6151
R2108 B.n265 B.n264 10.6151
R2109 B.n266 B.n265 10.6151
R2110 B.n266 B.n195 10.6151
R2111 B.n270 B.n195 10.6151
R2112 B.n271 B.n270 10.6151
R2113 B.n272 B.n271 10.6151
R2114 B.n272 B.n193 10.6151
R2115 B.n276 B.n193 10.6151
R2116 B.n277 B.n276 10.6151
R2117 B.n278 B.n277 10.6151
R2118 B.n278 B.n191 10.6151
R2119 B.n282 B.n191 10.6151
R2120 B.n283 B.n282 10.6151
R2121 B.n284 B.n283 10.6151
R2122 B.n284 B.n189 10.6151
R2123 B.n288 B.n189 10.6151
R2124 B.n289 B.n288 10.6151
R2125 B.n290 B.n289 10.6151
R2126 B.n290 B.n187 10.6151
R2127 B.n294 B.n187 10.6151
R2128 B.n295 B.n294 10.6151
R2129 B.n296 B.n295 10.6151
R2130 B.n296 B.n185 10.6151
R2131 B.n300 B.n185 10.6151
R2132 B.n302 B.n301 10.6151
R2133 B.n302 B.n183 10.6151
R2134 B.n306 B.n183 10.6151
R2135 B.n307 B.n306 10.6151
R2136 B.n308 B.n307 10.6151
R2137 B.n308 B.n181 10.6151
R2138 B.n312 B.n181 10.6151
R2139 B.n313 B.n312 10.6151
R2140 B.n314 B.n313 10.6151
R2141 B.n314 B.n179 10.6151
R2142 B.n318 B.n179 10.6151
R2143 B.n319 B.n318 10.6151
R2144 B.n320 B.n319 10.6151
R2145 B.n320 B.n177 10.6151
R2146 B.n324 B.n177 10.6151
R2147 B.n325 B.n324 10.6151
R2148 B.n326 B.n325 10.6151
R2149 B.n326 B.n175 10.6151
R2150 B.n330 B.n175 10.6151
R2151 B.n331 B.n330 10.6151
R2152 B.n332 B.n331 10.6151
R2153 B.n332 B.n173 10.6151
R2154 B.n336 B.n173 10.6151
R2155 B.n337 B.n336 10.6151
R2156 B.n338 B.n337 10.6151
R2157 B.n338 B.n171 10.6151
R2158 B.n342 B.n171 10.6151
R2159 B.n343 B.n342 10.6151
R2160 B.n344 B.n343 10.6151
R2161 B.n344 B.n169 10.6151
R2162 B.n348 B.n169 10.6151
R2163 B.n349 B.n348 10.6151
R2164 B.n350 B.n349 10.6151
R2165 B.n350 B.n167 10.6151
R2166 B.n354 B.n167 10.6151
R2167 B.n355 B.n354 10.6151
R2168 B.n359 B.n355 10.6151
R2169 B.n363 B.n165 10.6151
R2170 B.n364 B.n363 10.6151
R2171 B.n365 B.n364 10.6151
R2172 B.n365 B.n163 10.6151
R2173 B.n369 B.n163 10.6151
R2174 B.n370 B.n369 10.6151
R2175 B.n371 B.n370 10.6151
R2176 B.n371 B.n161 10.6151
R2177 B.n375 B.n161 10.6151
R2178 B.n378 B.n377 10.6151
R2179 B.n378 B.n157 10.6151
R2180 B.n382 B.n157 10.6151
R2181 B.n383 B.n382 10.6151
R2182 B.n384 B.n383 10.6151
R2183 B.n384 B.n155 10.6151
R2184 B.n388 B.n155 10.6151
R2185 B.n389 B.n388 10.6151
R2186 B.n390 B.n389 10.6151
R2187 B.n390 B.n153 10.6151
R2188 B.n394 B.n153 10.6151
R2189 B.n395 B.n394 10.6151
R2190 B.n396 B.n395 10.6151
R2191 B.n396 B.n151 10.6151
R2192 B.n400 B.n151 10.6151
R2193 B.n401 B.n400 10.6151
R2194 B.n402 B.n401 10.6151
R2195 B.n402 B.n149 10.6151
R2196 B.n406 B.n149 10.6151
R2197 B.n407 B.n406 10.6151
R2198 B.n408 B.n407 10.6151
R2199 B.n408 B.n147 10.6151
R2200 B.n412 B.n147 10.6151
R2201 B.n413 B.n412 10.6151
R2202 B.n414 B.n413 10.6151
R2203 B.n414 B.n145 10.6151
R2204 B.n418 B.n145 10.6151
R2205 B.n419 B.n418 10.6151
R2206 B.n420 B.n419 10.6151
R2207 B.n420 B.n143 10.6151
R2208 B.n424 B.n143 10.6151
R2209 B.n425 B.n424 10.6151
R2210 B.n426 B.n425 10.6151
R2211 B.n426 B.n141 10.6151
R2212 B.n430 B.n141 10.6151
R2213 B.n431 B.n430 10.6151
R2214 B.n432 B.n431 10.6151
R2215 B.n54 B.n50 9.36635
R2216 B.n671 B.n670 9.36635
R2217 B.n359 B.n358 9.36635
R2218 B.n377 B.n376 9.36635
R2219 B.n833 B.n0 8.11757
R2220 B.n833 B.n1 8.11757
R2221 B.n685 B.n54 1.24928
R2222 B.n672 B.n671 1.24928
R2223 B.n358 B.n165 1.24928
R2224 B.n376 B.n375 1.24928
C0 VTAIL w_n4450_n3132# 4.00042f
C1 VTAIL B 4.82243f
C2 B w_n4450_n3132# 10.6268f
C3 VN VTAIL 8.79099f
C4 VN w_n4450_n3132# 9.18821f
C5 VTAIL VP 8.805099f
C6 VP w_n4450_n3132# 9.76754f
C7 VTAIL VDD1 7.89639f
C8 VDD1 w_n4450_n3132# 2.10331f
C9 VN B 1.3351f
C10 B VP 2.30917f
C11 VDD1 B 1.785f
C12 VDD2 w_n4450_n3132# 2.24109f
C13 VTAIL VDD2 7.9545f
C14 VN VP 8.1213f
C15 VN VDD1 0.152515f
C16 VDD2 B 1.89833f
C17 VDD1 VP 8.577559f
C18 VN VDD2 8.153759f
C19 VDD2 VP 0.577989f
C20 VDD1 VDD2 2.0648f
C21 VDD2 VSUBS 2.151032f
C22 VDD1 VSUBS 2.89422f
C23 VTAIL VSUBS 1.385179f
C24 VN VSUBS 7.45745f
C25 VP VSUBS 4.124053f
C26 B VSUBS 5.517858f
C27 w_n4450_n3132# VSUBS 0.171895p
C28 B.n0 VSUBS 0.006712f
C29 B.n1 VSUBS 0.006712f
C30 B.n2 VSUBS 0.009927f
C31 B.n3 VSUBS 0.007607f
C32 B.n4 VSUBS 0.007607f
C33 B.n5 VSUBS 0.007607f
C34 B.n6 VSUBS 0.007607f
C35 B.n7 VSUBS 0.007607f
C36 B.n8 VSUBS 0.007607f
C37 B.n9 VSUBS 0.007607f
C38 B.n10 VSUBS 0.007607f
C39 B.n11 VSUBS 0.007607f
C40 B.n12 VSUBS 0.007607f
C41 B.n13 VSUBS 0.007607f
C42 B.n14 VSUBS 0.007607f
C43 B.n15 VSUBS 0.007607f
C44 B.n16 VSUBS 0.007607f
C45 B.n17 VSUBS 0.007607f
C46 B.n18 VSUBS 0.007607f
C47 B.n19 VSUBS 0.007607f
C48 B.n20 VSUBS 0.007607f
C49 B.n21 VSUBS 0.007607f
C50 B.n22 VSUBS 0.007607f
C51 B.n23 VSUBS 0.007607f
C52 B.n24 VSUBS 0.007607f
C53 B.n25 VSUBS 0.007607f
C54 B.n26 VSUBS 0.007607f
C55 B.n27 VSUBS 0.007607f
C56 B.n28 VSUBS 0.007607f
C57 B.n29 VSUBS 0.007607f
C58 B.n30 VSUBS 0.007607f
C59 B.n31 VSUBS 0.016316f
C60 B.n32 VSUBS 0.007607f
C61 B.n33 VSUBS 0.007607f
C62 B.n34 VSUBS 0.007607f
C63 B.n35 VSUBS 0.007607f
C64 B.n36 VSUBS 0.007607f
C65 B.n37 VSUBS 0.007607f
C66 B.n38 VSUBS 0.007607f
C67 B.n39 VSUBS 0.007607f
C68 B.n40 VSUBS 0.007607f
C69 B.n41 VSUBS 0.007607f
C70 B.n42 VSUBS 0.007607f
C71 B.n43 VSUBS 0.007607f
C72 B.n44 VSUBS 0.007607f
C73 B.n45 VSUBS 0.007607f
C74 B.n46 VSUBS 0.007607f
C75 B.n47 VSUBS 0.007607f
C76 B.n48 VSUBS 0.007607f
C77 B.n49 VSUBS 0.007607f
C78 B.n50 VSUBS 0.007159f
C79 B.n51 VSUBS 0.007607f
C80 B.t10 VSUBS 0.201344f
C81 B.t11 VSUBS 0.24083f
C82 B.t9 VSUBS 1.71815f
C83 B.n52 VSUBS 0.386422f
C84 B.n53 VSUBS 0.257759f
C85 B.n54 VSUBS 0.017624f
C86 B.n55 VSUBS 0.007607f
C87 B.n56 VSUBS 0.007607f
C88 B.n57 VSUBS 0.007607f
C89 B.n58 VSUBS 0.007607f
C90 B.t7 VSUBS 0.201347f
C91 B.t8 VSUBS 0.240833f
C92 B.t6 VSUBS 1.71815f
C93 B.n59 VSUBS 0.386419f
C94 B.n60 VSUBS 0.257756f
C95 B.n61 VSUBS 0.007607f
C96 B.n62 VSUBS 0.007607f
C97 B.n63 VSUBS 0.007607f
C98 B.n64 VSUBS 0.007607f
C99 B.n65 VSUBS 0.007607f
C100 B.n66 VSUBS 0.007607f
C101 B.n67 VSUBS 0.007607f
C102 B.n68 VSUBS 0.007607f
C103 B.n69 VSUBS 0.007607f
C104 B.n70 VSUBS 0.007607f
C105 B.n71 VSUBS 0.007607f
C106 B.n72 VSUBS 0.007607f
C107 B.n73 VSUBS 0.007607f
C108 B.n74 VSUBS 0.007607f
C109 B.n75 VSUBS 0.007607f
C110 B.n76 VSUBS 0.007607f
C111 B.n77 VSUBS 0.007607f
C112 B.n78 VSUBS 0.007607f
C113 B.n79 VSUBS 0.01702f
C114 B.n80 VSUBS 0.007607f
C115 B.n81 VSUBS 0.007607f
C116 B.n82 VSUBS 0.007607f
C117 B.n83 VSUBS 0.007607f
C118 B.n84 VSUBS 0.007607f
C119 B.n85 VSUBS 0.007607f
C120 B.n86 VSUBS 0.007607f
C121 B.n87 VSUBS 0.007607f
C122 B.n88 VSUBS 0.007607f
C123 B.n89 VSUBS 0.007607f
C124 B.n90 VSUBS 0.007607f
C125 B.n91 VSUBS 0.007607f
C126 B.n92 VSUBS 0.007607f
C127 B.n93 VSUBS 0.007607f
C128 B.n94 VSUBS 0.007607f
C129 B.n95 VSUBS 0.007607f
C130 B.n96 VSUBS 0.007607f
C131 B.n97 VSUBS 0.007607f
C132 B.n98 VSUBS 0.007607f
C133 B.n99 VSUBS 0.007607f
C134 B.n100 VSUBS 0.007607f
C135 B.n101 VSUBS 0.007607f
C136 B.n102 VSUBS 0.007607f
C137 B.n103 VSUBS 0.007607f
C138 B.n104 VSUBS 0.007607f
C139 B.n105 VSUBS 0.007607f
C140 B.n106 VSUBS 0.007607f
C141 B.n107 VSUBS 0.007607f
C142 B.n108 VSUBS 0.007607f
C143 B.n109 VSUBS 0.007607f
C144 B.n110 VSUBS 0.007607f
C145 B.n111 VSUBS 0.007607f
C146 B.n112 VSUBS 0.007607f
C147 B.n113 VSUBS 0.007607f
C148 B.n114 VSUBS 0.007607f
C149 B.n115 VSUBS 0.007607f
C150 B.n116 VSUBS 0.007607f
C151 B.n117 VSUBS 0.007607f
C152 B.n118 VSUBS 0.007607f
C153 B.n119 VSUBS 0.007607f
C154 B.n120 VSUBS 0.007607f
C155 B.n121 VSUBS 0.007607f
C156 B.n122 VSUBS 0.007607f
C157 B.n123 VSUBS 0.007607f
C158 B.n124 VSUBS 0.007607f
C159 B.n125 VSUBS 0.007607f
C160 B.n126 VSUBS 0.007607f
C161 B.n127 VSUBS 0.007607f
C162 B.n128 VSUBS 0.007607f
C163 B.n129 VSUBS 0.007607f
C164 B.n130 VSUBS 0.007607f
C165 B.n131 VSUBS 0.007607f
C166 B.n132 VSUBS 0.007607f
C167 B.n133 VSUBS 0.007607f
C168 B.n134 VSUBS 0.007607f
C169 B.n135 VSUBS 0.007607f
C170 B.n136 VSUBS 0.007607f
C171 B.n137 VSUBS 0.007607f
C172 B.n138 VSUBS 0.007607f
C173 B.n139 VSUBS 0.017311f
C174 B.n140 VSUBS 0.007607f
C175 B.n141 VSUBS 0.007607f
C176 B.n142 VSUBS 0.007607f
C177 B.n143 VSUBS 0.007607f
C178 B.n144 VSUBS 0.007607f
C179 B.n145 VSUBS 0.007607f
C180 B.n146 VSUBS 0.007607f
C181 B.n147 VSUBS 0.007607f
C182 B.n148 VSUBS 0.007607f
C183 B.n149 VSUBS 0.007607f
C184 B.n150 VSUBS 0.007607f
C185 B.n151 VSUBS 0.007607f
C186 B.n152 VSUBS 0.007607f
C187 B.n153 VSUBS 0.007607f
C188 B.n154 VSUBS 0.007607f
C189 B.n155 VSUBS 0.007607f
C190 B.n156 VSUBS 0.007607f
C191 B.n157 VSUBS 0.007607f
C192 B.n158 VSUBS 0.007607f
C193 B.t2 VSUBS 0.201347f
C194 B.t1 VSUBS 0.240833f
C195 B.t0 VSUBS 1.71815f
C196 B.n159 VSUBS 0.386419f
C197 B.n160 VSUBS 0.257756f
C198 B.n161 VSUBS 0.007607f
C199 B.n162 VSUBS 0.007607f
C200 B.n163 VSUBS 0.007607f
C201 B.n164 VSUBS 0.007607f
C202 B.n165 VSUBS 0.004251f
C203 B.n166 VSUBS 0.007607f
C204 B.n167 VSUBS 0.007607f
C205 B.n168 VSUBS 0.007607f
C206 B.n169 VSUBS 0.007607f
C207 B.n170 VSUBS 0.007607f
C208 B.n171 VSUBS 0.007607f
C209 B.n172 VSUBS 0.007607f
C210 B.n173 VSUBS 0.007607f
C211 B.n174 VSUBS 0.007607f
C212 B.n175 VSUBS 0.007607f
C213 B.n176 VSUBS 0.007607f
C214 B.n177 VSUBS 0.007607f
C215 B.n178 VSUBS 0.007607f
C216 B.n179 VSUBS 0.007607f
C217 B.n180 VSUBS 0.007607f
C218 B.n181 VSUBS 0.007607f
C219 B.n182 VSUBS 0.007607f
C220 B.n183 VSUBS 0.007607f
C221 B.n184 VSUBS 0.01702f
C222 B.n185 VSUBS 0.007607f
C223 B.n186 VSUBS 0.007607f
C224 B.n187 VSUBS 0.007607f
C225 B.n188 VSUBS 0.007607f
C226 B.n189 VSUBS 0.007607f
C227 B.n190 VSUBS 0.007607f
C228 B.n191 VSUBS 0.007607f
C229 B.n192 VSUBS 0.007607f
C230 B.n193 VSUBS 0.007607f
C231 B.n194 VSUBS 0.007607f
C232 B.n195 VSUBS 0.007607f
C233 B.n196 VSUBS 0.007607f
C234 B.n197 VSUBS 0.007607f
C235 B.n198 VSUBS 0.007607f
C236 B.n199 VSUBS 0.007607f
C237 B.n200 VSUBS 0.007607f
C238 B.n201 VSUBS 0.007607f
C239 B.n202 VSUBS 0.007607f
C240 B.n203 VSUBS 0.007607f
C241 B.n204 VSUBS 0.007607f
C242 B.n205 VSUBS 0.007607f
C243 B.n206 VSUBS 0.007607f
C244 B.n207 VSUBS 0.007607f
C245 B.n208 VSUBS 0.007607f
C246 B.n209 VSUBS 0.007607f
C247 B.n210 VSUBS 0.007607f
C248 B.n211 VSUBS 0.007607f
C249 B.n212 VSUBS 0.007607f
C250 B.n213 VSUBS 0.007607f
C251 B.n214 VSUBS 0.007607f
C252 B.n215 VSUBS 0.007607f
C253 B.n216 VSUBS 0.007607f
C254 B.n217 VSUBS 0.007607f
C255 B.n218 VSUBS 0.007607f
C256 B.n219 VSUBS 0.007607f
C257 B.n220 VSUBS 0.007607f
C258 B.n221 VSUBS 0.007607f
C259 B.n222 VSUBS 0.007607f
C260 B.n223 VSUBS 0.007607f
C261 B.n224 VSUBS 0.007607f
C262 B.n225 VSUBS 0.007607f
C263 B.n226 VSUBS 0.007607f
C264 B.n227 VSUBS 0.007607f
C265 B.n228 VSUBS 0.007607f
C266 B.n229 VSUBS 0.007607f
C267 B.n230 VSUBS 0.007607f
C268 B.n231 VSUBS 0.007607f
C269 B.n232 VSUBS 0.007607f
C270 B.n233 VSUBS 0.007607f
C271 B.n234 VSUBS 0.007607f
C272 B.n235 VSUBS 0.007607f
C273 B.n236 VSUBS 0.007607f
C274 B.n237 VSUBS 0.007607f
C275 B.n238 VSUBS 0.007607f
C276 B.n239 VSUBS 0.007607f
C277 B.n240 VSUBS 0.007607f
C278 B.n241 VSUBS 0.007607f
C279 B.n242 VSUBS 0.007607f
C280 B.n243 VSUBS 0.007607f
C281 B.n244 VSUBS 0.007607f
C282 B.n245 VSUBS 0.007607f
C283 B.n246 VSUBS 0.007607f
C284 B.n247 VSUBS 0.007607f
C285 B.n248 VSUBS 0.007607f
C286 B.n249 VSUBS 0.007607f
C287 B.n250 VSUBS 0.007607f
C288 B.n251 VSUBS 0.007607f
C289 B.n252 VSUBS 0.007607f
C290 B.n253 VSUBS 0.007607f
C291 B.n254 VSUBS 0.007607f
C292 B.n255 VSUBS 0.007607f
C293 B.n256 VSUBS 0.007607f
C294 B.n257 VSUBS 0.007607f
C295 B.n258 VSUBS 0.007607f
C296 B.n259 VSUBS 0.007607f
C297 B.n260 VSUBS 0.007607f
C298 B.n261 VSUBS 0.007607f
C299 B.n262 VSUBS 0.007607f
C300 B.n263 VSUBS 0.007607f
C301 B.n264 VSUBS 0.007607f
C302 B.n265 VSUBS 0.007607f
C303 B.n266 VSUBS 0.007607f
C304 B.n267 VSUBS 0.007607f
C305 B.n268 VSUBS 0.007607f
C306 B.n269 VSUBS 0.007607f
C307 B.n270 VSUBS 0.007607f
C308 B.n271 VSUBS 0.007607f
C309 B.n272 VSUBS 0.007607f
C310 B.n273 VSUBS 0.007607f
C311 B.n274 VSUBS 0.007607f
C312 B.n275 VSUBS 0.007607f
C313 B.n276 VSUBS 0.007607f
C314 B.n277 VSUBS 0.007607f
C315 B.n278 VSUBS 0.007607f
C316 B.n279 VSUBS 0.007607f
C317 B.n280 VSUBS 0.007607f
C318 B.n281 VSUBS 0.007607f
C319 B.n282 VSUBS 0.007607f
C320 B.n283 VSUBS 0.007607f
C321 B.n284 VSUBS 0.007607f
C322 B.n285 VSUBS 0.007607f
C323 B.n286 VSUBS 0.007607f
C324 B.n287 VSUBS 0.007607f
C325 B.n288 VSUBS 0.007607f
C326 B.n289 VSUBS 0.007607f
C327 B.n290 VSUBS 0.007607f
C328 B.n291 VSUBS 0.007607f
C329 B.n292 VSUBS 0.007607f
C330 B.n293 VSUBS 0.007607f
C331 B.n294 VSUBS 0.007607f
C332 B.n295 VSUBS 0.007607f
C333 B.n296 VSUBS 0.007607f
C334 B.n297 VSUBS 0.007607f
C335 B.n298 VSUBS 0.007607f
C336 B.n299 VSUBS 0.016316f
C337 B.n300 VSUBS 0.016316f
C338 B.n301 VSUBS 0.01702f
C339 B.n302 VSUBS 0.007607f
C340 B.n303 VSUBS 0.007607f
C341 B.n304 VSUBS 0.007607f
C342 B.n305 VSUBS 0.007607f
C343 B.n306 VSUBS 0.007607f
C344 B.n307 VSUBS 0.007607f
C345 B.n308 VSUBS 0.007607f
C346 B.n309 VSUBS 0.007607f
C347 B.n310 VSUBS 0.007607f
C348 B.n311 VSUBS 0.007607f
C349 B.n312 VSUBS 0.007607f
C350 B.n313 VSUBS 0.007607f
C351 B.n314 VSUBS 0.007607f
C352 B.n315 VSUBS 0.007607f
C353 B.n316 VSUBS 0.007607f
C354 B.n317 VSUBS 0.007607f
C355 B.n318 VSUBS 0.007607f
C356 B.n319 VSUBS 0.007607f
C357 B.n320 VSUBS 0.007607f
C358 B.n321 VSUBS 0.007607f
C359 B.n322 VSUBS 0.007607f
C360 B.n323 VSUBS 0.007607f
C361 B.n324 VSUBS 0.007607f
C362 B.n325 VSUBS 0.007607f
C363 B.n326 VSUBS 0.007607f
C364 B.n327 VSUBS 0.007607f
C365 B.n328 VSUBS 0.007607f
C366 B.n329 VSUBS 0.007607f
C367 B.n330 VSUBS 0.007607f
C368 B.n331 VSUBS 0.007607f
C369 B.n332 VSUBS 0.007607f
C370 B.n333 VSUBS 0.007607f
C371 B.n334 VSUBS 0.007607f
C372 B.n335 VSUBS 0.007607f
C373 B.n336 VSUBS 0.007607f
C374 B.n337 VSUBS 0.007607f
C375 B.n338 VSUBS 0.007607f
C376 B.n339 VSUBS 0.007607f
C377 B.n340 VSUBS 0.007607f
C378 B.n341 VSUBS 0.007607f
C379 B.n342 VSUBS 0.007607f
C380 B.n343 VSUBS 0.007607f
C381 B.n344 VSUBS 0.007607f
C382 B.n345 VSUBS 0.007607f
C383 B.n346 VSUBS 0.007607f
C384 B.n347 VSUBS 0.007607f
C385 B.n348 VSUBS 0.007607f
C386 B.n349 VSUBS 0.007607f
C387 B.n350 VSUBS 0.007607f
C388 B.n351 VSUBS 0.007607f
C389 B.n352 VSUBS 0.007607f
C390 B.n353 VSUBS 0.007607f
C391 B.n354 VSUBS 0.007607f
C392 B.n355 VSUBS 0.007607f
C393 B.t5 VSUBS 0.201344f
C394 B.t4 VSUBS 0.24083f
C395 B.t3 VSUBS 1.71815f
C396 B.n356 VSUBS 0.386422f
C397 B.n357 VSUBS 0.257759f
C398 B.n358 VSUBS 0.017624f
C399 B.n359 VSUBS 0.007159f
C400 B.n360 VSUBS 0.007607f
C401 B.n361 VSUBS 0.007607f
C402 B.n362 VSUBS 0.007607f
C403 B.n363 VSUBS 0.007607f
C404 B.n364 VSUBS 0.007607f
C405 B.n365 VSUBS 0.007607f
C406 B.n366 VSUBS 0.007607f
C407 B.n367 VSUBS 0.007607f
C408 B.n368 VSUBS 0.007607f
C409 B.n369 VSUBS 0.007607f
C410 B.n370 VSUBS 0.007607f
C411 B.n371 VSUBS 0.007607f
C412 B.n372 VSUBS 0.007607f
C413 B.n373 VSUBS 0.007607f
C414 B.n374 VSUBS 0.007607f
C415 B.n375 VSUBS 0.004251f
C416 B.n376 VSUBS 0.017624f
C417 B.n377 VSUBS 0.007159f
C418 B.n378 VSUBS 0.007607f
C419 B.n379 VSUBS 0.007607f
C420 B.n380 VSUBS 0.007607f
C421 B.n381 VSUBS 0.007607f
C422 B.n382 VSUBS 0.007607f
C423 B.n383 VSUBS 0.007607f
C424 B.n384 VSUBS 0.007607f
C425 B.n385 VSUBS 0.007607f
C426 B.n386 VSUBS 0.007607f
C427 B.n387 VSUBS 0.007607f
C428 B.n388 VSUBS 0.007607f
C429 B.n389 VSUBS 0.007607f
C430 B.n390 VSUBS 0.007607f
C431 B.n391 VSUBS 0.007607f
C432 B.n392 VSUBS 0.007607f
C433 B.n393 VSUBS 0.007607f
C434 B.n394 VSUBS 0.007607f
C435 B.n395 VSUBS 0.007607f
C436 B.n396 VSUBS 0.007607f
C437 B.n397 VSUBS 0.007607f
C438 B.n398 VSUBS 0.007607f
C439 B.n399 VSUBS 0.007607f
C440 B.n400 VSUBS 0.007607f
C441 B.n401 VSUBS 0.007607f
C442 B.n402 VSUBS 0.007607f
C443 B.n403 VSUBS 0.007607f
C444 B.n404 VSUBS 0.007607f
C445 B.n405 VSUBS 0.007607f
C446 B.n406 VSUBS 0.007607f
C447 B.n407 VSUBS 0.007607f
C448 B.n408 VSUBS 0.007607f
C449 B.n409 VSUBS 0.007607f
C450 B.n410 VSUBS 0.007607f
C451 B.n411 VSUBS 0.007607f
C452 B.n412 VSUBS 0.007607f
C453 B.n413 VSUBS 0.007607f
C454 B.n414 VSUBS 0.007607f
C455 B.n415 VSUBS 0.007607f
C456 B.n416 VSUBS 0.007607f
C457 B.n417 VSUBS 0.007607f
C458 B.n418 VSUBS 0.007607f
C459 B.n419 VSUBS 0.007607f
C460 B.n420 VSUBS 0.007607f
C461 B.n421 VSUBS 0.007607f
C462 B.n422 VSUBS 0.007607f
C463 B.n423 VSUBS 0.007607f
C464 B.n424 VSUBS 0.007607f
C465 B.n425 VSUBS 0.007607f
C466 B.n426 VSUBS 0.007607f
C467 B.n427 VSUBS 0.007607f
C468 B.n428 VSUBS 0.007607f
C469 B.n429 VSUBS 0.007607f
C470 B.n430 VSUBS 0.007607f
C471 B.n431 VSUBS 0.007607f
C472 B.n432 VSUBS 0.016025f
C473 B.n433 VSUBS 0.01702f
C474 B.n434 VSUBS 0.016316f
C475 B.n435 VSUBS 0.007607f
C476 B.n436 VSUBS 0.007607f
C477 B.n437 VSUBS 0.007607f
C478 B.n438 VSUBS 0.007607f
C479 B.n439 VSUBS 0.007607f
C480 B.n440 VSUBS 0.007607f
C481 B.n441 VSUBS 0.007607f
C482 B.n442 VSUBS 0.007607f
C483 B.n443 VSUBS 0.007607f
C484 B.n444 VSUBS 0.007607f
C485 B.n445 VSUBS 0.007607f
C486 B.n446 VSUBS 0.007607f
C487 B.n447 VSUBS 0.007607f
C488 B.n448 VSUBS 0.007607f
C489 B.n449 VSUBS 0.007607f
C490 B.n450 VSUBS 0.007607f
C491 B.n451 VSUBS 0.007607f
C492 B.n452 VSUBS 0.007607f
C493 B.n453 VSUBS 0.007607f
C494 B.n454 VSUBS 0.007607f
C495 B.n455 VSUBS 0.007607f
C496 B.n456 VSUBS 0.007607f
C497 B.n457 VSUBS 0.007607f
C498 B.n458 VSUBS 0.007607f
C499 B.n459 VSUBS 0.007607f
C500 B.n460 VSUBS 0.007607f
C501 B.n461 VSUBS 0.007607f
C502 B.n462 VSUBS 0.007607f
C503 B.n463 VSUBS 0.007607f
C504 B.n464 VSUBS 0.007607f
C505 B.n465 VSUBS 0.007607f
C506 B.n466 VSUBS 0.007607f
C507 B.n467 VSUBS 0.007607f
C508 B.n468 VSUBS 0.007607f
C509 B.n469 VSUBS 0.007607f
C510 B.n470 VSUBS 0.007607f
C511 B.n471 VSUBS 0.007607f
C512 B.n472 VSUBS 0.007607f
C513 B.n473 VSUBS 0.007607f
C514 B.n474 VSUBS 0.007607f
C515 B.n475 VSUBS 0.007607f
C516 B.n476 VSUBS 0.007607f
C517 B.n477 VSUBS 0.007607f
C518 B.n478 VSUBS 0.007607f
C519 B.n479 VSUBS 0.007607f
C520 B.n480 VSUBS 0.007607f
C521 B.n481 VSUBS 0.007607f
C522 B.n482 VSUBS 0.007607f
C523 B.n483 VSUBS 0.007607f
C524 B.n484 VSUBS 0.007607f
C525 B.n485 VSUBS 0.007607f
C526 B.n486 VSUBS 0.007607f
C527 B.n487 VSUBS 0.007607f
C528 B.n488 VSUBS 0.007607f
C529 B.n489 VSUBS 0.007607f
C530 B.n490 VSUBS 0.007607f
C531 B.n491 VSUBS 0.007607f
C532 B.n492 VSUBS 0.007607f
C533 B.n493 VSUBS 0.007607f
C534 B.n494 VSUBS 0.007607f
C535 B.n495 VSUBS 0.007607f
C536 B.n496 VSUBS 0.007607f
C537 B.n497 VSUBS 0.007607f
C538 B.n498 VSUBS 0.007607f
C539 B.n499 VSUBS 0.007607f
C540 B.n500 VSUBS 0.007607f
C541 B.n501 VSUBS 0.007607f
C542 B.n502 VSUBS 0.007607f
C543 B.n503 VSUBS 0.007607f
C544 B.n504 VSUBS 0.007607f
C545 B.n505 VSUBS 0.007607f
C546 B.n506 VSUBS 0.007607f
C547 B.n507 VSUBS 0.007607f
C548 B.n508 VSUBS 0.007607f
C549 B.n509 VSUBS 0.007607f
C550 B.n510 VSUBS 0.007607f
C551 B.n511 VSUBS 0.007607f
C552 B.n512 VSUBS 0.007607f
C553 B.n513 VSUBS 0.007607f
C554 B.n514 VSUBS 0.007607f
C555 B.n515 VSUBS 0.007607f
C556 B.n516 VSUBS 0.007607f
C557 B.n517 VSUBS 0.007607f
C558 B.n518 VSUBS 0.007607f
C559 B.n519 VSUBS 0.007607f
C560 B.n520 VSUBS 0.007607f
C561 B.n521 VSUBS 0.007607f
C562 B.n522 VSUBS 0.007607f
C563 B.n523 VSUBS 0.007607f
C564 B.n524 VSUBS 0.007607f
C565 B.n525 VSUBS 0.007607f
C566 B.n526 VSUBS 0.007607f
C567 B.n527 VSUBS 0.007607f
C568 B.n528 VSUBS 0.007607f
C569 B.n529 VSUBS 0.007607f
C570 B.n530 VSUBS 0.007607f
C571 B.n531 VSUBS 0.007607f
C572 B.n532 VSUBS 0.007607f
C573 B.n533 VSUBS 0.007607f
C574 B.n534 VSUBS 0.007607f
C575 B.n535 VSUBS 0.007607f
C576 B.n536 VSUBS 0.007607f
C577 B.n537 VSUBS 0.007607f
C578 B.n538 VSUBS 0.007607f
C579 B.n539 VSUBS 0.007607f
C580 B.n540 VSUBS 0.007607f
C581 B.n541 VSUBS 0.007607f
C582 B.n542 VSUBS 0.007607f
C583 B.n543 VSUBS 0.007607f
C584 B.n544 VSUBS 0.007607f
C585 B.n545 VSUBS 0.007607f
C586 B.n546 VSUBS 0.007607f
C587 B.n547 VSUBS 0.007607f
C588 B.n548 VSUBS 0.007607f
C589 B.n549 VSUBS 0.007607f
C590 B.n550 VSUBS 0.007607f
C591 B.n551 VSUBS 0.007607f
C592 B.n552 VSUBS 0.007607f
C593 B.n553 VSUBS 0.007607f
C594 B.n554 VSUBS 0.007607f
C595 B.n555 VSUBS 0.007607f
C596 B.n556 VSUBS 0.007607f
C597 B.n557 VSUBS 0.007607f
C598 B.n558 VSUBS 0.007607f
C599 B.n559 VSUBS 0.007607f
C600 B.n560 VSUBS 0.007607f
C601 B.n561 VSUBS 0.007607f
C602 B.n562 VSUBS 0.007607f
C603 B.n563 VSUBS 0.007607f
C604 B.n564 VSUBS 0.007607f
C605 B.n565 VSUBS 0.007607f
C606 B.n566 VSUBS 0.007607f
C607 B.n567 VSUBS 0.007607f
C608 B.n568 VSUBS 0.007607f
C609 B.n569 VSUBS 0.007607f
C610 B.n570 VSUBS 0.007607f
C611 B.n571 VSUBS 0.007607f
C612 B.n572 VSUBS 0.007607f
C613 B.n573 VSUBS 0.007607f
C614 B.n574 VSUBS 0.007607f
C615 B.n575 VSUBS 0.007607f
C616 B.n576 VSUBS 0.007607f
C617 B.n577 VSUBS 0.007607f
C618 B.n578 VSUBS 0.007607f
C619 B.n579 VSUBS 0.007607f
C620 B.n580 VSUBS 0.007607f
C621 B.n581 VSUBS 0.007607f
C622 B.n582 VSUBS 0.007607f
C623 B.n583 VSUBS 0.007607f
C624 B.n584 VSUBS 0.007607f
C625 B.n585 VSUBS 0.007607f
C626 B.n586 VSUBS 0.007607f
C627 B.n587 VSUBS 0.007607f
C628 B.n588 VSUBS 0.007607f
C629 B.n589 VSUBS 0.007607f
C630 B.n590 VSUBS 0.007607f
C631 B.n591 VSUBS 0.007607f
C632 B.n592 VSUBS 0.007607f
C633 B.n593 VSUBS 0.007607f
C634 B.n594 VSUBS 0.007607f
C635 B.n595 VSUBS 0.007607f
C636 B.n596 VSUBS 0.007607f
C637 B.n597 VSUBS 0.007607f
C638 B.n598 VSUBS 0.007607f
C639 B.n599 VSUBS 0.007607f
C640 B.n600 VSUBS 0.007607f
C641 B.n601 VSUBS 0.007607f
C642 B.n602 VSUBS 0.007607f
C643 B.n603 VSUBS 0.007607f
C644 B.n604 VSUBS 0.007607f
C645 B.n605 VSUBS 0.007607f
C646 B.n606 VSUBS 0.007607f
C647 B.n607 VSUBS 0.007607f
C648 B.n608 VSUBS 0.007607f
C649 B.n609 VSUBS 0.007607f
C650 B.n610 VSUBS 0.007607f
C651 B.n611 VSUBS 0.007607f
C652 B.n612 VSUBS 0.016316f
C653 B.n613 VSUBS 0.016316f
C654 B.n614 VSUBS 0.01702f
C655 B.n615 VSUBS 0.007607f
C656 B.n616 VSUBS 0.007607f
C657 B.n617 VSUBS 0.007607f
C658 B.n618 VSUBS 0.007607f
C659 B.n619 VSUBS 0.007607f
C660 B.n620 VSUBS 0.007607f
C661 B.n621 VSUBS 0.007607f
C662 B.n622 VSUBS 0.007607f
C663 B.n623 VSUBS 0.007607f
C664 B.n624 VSUBS 0.007607f
C665 B.n625 VSUBS 0.007607f
C666 B.n626 VSUBS 0.007607f
C667 B.n627 VSUBS 0.007607f
C668 B.n628 VSUBS 0.007607f
C669 B.n629 VSUBS 0.007607f
C670 B.n630 VSUBS 0.007607f
C671 B.n631 VSUBS 0.007607f
C672 B.n632 VSUBS 0.007607f
C673 B.n633 VSUBS 0.007607f
C674 B.n634 VSUBS 0.007607f
C675 B.n635 VSUBS 0.007607f
C676 B.n636 VSUBS 0.007607f
C677 B.n637 VSUBS 0.007607f
C678 B.n638 VSUBS 0.007607f
C679 B.n639 VSUBS 0.007607f
C680 B.n640 VSUBS 0.007607f
C681 B.n641 VSUBS 0.007607f
C682 B.n642 VSUBS 0.007607f
C683 B.n643 VSUBS 0.007607f
C684 B.n644 VSUBS 0.007607f
C685 B.n645 VSUBS 0.007607f
C686 B.n646 VSUBS 0.007607f
C687 B.n647 VSUBS 0.007607f
C688 B.n648 VSUBS 0.007607f
C689 B.n649 VSUBS 0.007607f
C690 B.n650 VSUBS 0.007607f
C691 B.n651 VSUBS 0.007607f
C692 B.n652 VSUBS 0.007607f
C693 B.n653 VSUBS 0.007607f
C694 B.n654 VSUBS 0.007607f
C695 B.n655 VSUBS 0.007607f
C696 B.n656 VSUBS 0.007607f
C697 B.n657 VSUBS 0.007607f
C698 B.n658 VSUBS 0.007607f
C699 B.n659 VSUBS 0.007607f
C700 B.n660 VSUBS 0.007607f
C701 B.n661 VSUBS 0.007607f
C702 B.n662 VSUBS 0.007607f
C703 B.n663 VSUBS 0.007607f
C704 B.n664 VSUBS 0.007607f
C705 B.n665 VSUBS 0.007607f
C706 B.n666 VSUBS 0.007607f
C707 B.n667 VSUBS 0.007607f
C708 B.n668 VSUBS 0.007607f
C709 B.n669 VSUBS 0.007607f
C710 B.n670 VSUBS 0.007159f
C711 B.n671 VSUBS 0.017624f
C712 B.n672 VSUBS 0.004251f
C713 B.n673 VSUBS 0.007607f
C714 B.n674 VSUBS 0.007607f
C715 B.n675 VSUBS 0.007607f
C716 B.n676 VSUBS 0.007607f
C717 B.n677 VSUBS 0.007607f
C718 B.n678 VSUBS 0.007607f
C719 B.n679 VSUBS 0.007607f
C720 B.n680 VSUBS 0.007607f
C721 B.n681 VSUBS 0.007607f
C722 B.n682 VSUBS 0.007607f
C723 B.n683 VSUBS 0.007607f
C724 B.n684 VSUBS 0.007607f
C725 B.n685 VSUBS 0.004251f
C726 B.n686 VSUBS 0.007607f
C727 B.n687 VSUBS 0.007607f
C728 B.n688 VSUBS 0.007607f
C729 B.n689 VSUBS 0.007607f
C730 B.n690 VSUBS 0.007607f
C731 B.n691 VSUBS 0.007607f
C732 B.n692 VSUBS 0.007607f
C733 B.n693 VSUBS 0.007607f
C734 B.n694 VSUBS 0.007607f
C735 B.n695 VSUBS 0.007607f
C736 B.n696 VSUBS 0.007607f
C737 B.n697 VSUBS 0.007607f
C738 B.n698 VSUBS 0.007607f
C739 B.n699 VSUBS 0.007607f
C740 B.n700 VSUBS 0.007607f
C741 B.n701 VSUBS 0.007607f
C742 B.n702 VSUBS 0.007607f
C743 B.n703 VSUBS 0.007607f
C744 B.n704 VSUBS 0.007607f
C745 B.n705 VSUBS 0.007607f
C746 B.n706 VSUBS 0.007607f
C747 B.n707 VSUBS 0.007607f
C748 B.n708 VSUBS 0.007607f
C749 B.n709 VSUBS 0.007607f
C750 B.n710 VSUBS 0.007607f
C751 B.n711 VSUBS 0.007607f
C752 B.n712 VSUBS 0.007607f
C753 B.n713 VSUBS 0.007607f
C754 B.n714 VSUBS 0.007607f
C755 B.n715 VSUBS 0.007607f
C756 B.n716 VSUBS 0.007607f
C757 B.n717 VSUBS 0.007607f
C758 B.n718 VSUBS 0.007607f
C759 B.n719 VSUBS 0.007607f
C760 B.n720 VSUBS 0.007607f
C761 B.n721 VSUBS 0.007607f
C762 B.n722 VSUBS 0.007607f
C763 B.n723 VSUBS 0.007607f
C764 B.n724 VSUBS 0.007607f
C765 B.n725 VSUBS 0.007607f
C766 B.n726 VSUBS 0.007607f
C767 B.n727 VSUBS 0.007607f
C768 B.n728 VSUBS 0.007607f
C769 B.n729 VSUBS 0.007607f
C770 B.n730 VSUBS 0.007607f
C771 B.n731 VSUBS 0.007607f
C772 B.n732 VSUBS 0.007607f
C773 B.n733 VSUBS 0.007607f
C774 B.n734 VSUBS 0.007607f
C775 B.n735 VSUBS 0.007607f
C776 B.n736 VSUBS 0.007607f
C777 B.n737 VSUBS 0.007607f
C778 B.n738 VSUBS 0.007607f
C779 B.n739 VSUBS 0.007607f
C780 B.n740 VSUBS 0.007607f
C781 B.n741 VSUBS 0.007607f
C782 B.n742 VSUBS 0.01702f
C783 B.n743 VSUBS 0.01702f
C784 B.n744 VSUBS 0.016316f
C785 B.n745 VSUBS 0.007607f
C786 B.n746 VSUBS 0.007607f
C787 B.n747 VSUBS 0.007607f
C788 B.n748 VSUBS 0.007607f
C789 B.n749 VSUBS 0.007607f
C790 B.n750 VSUBS 0.007607f
C791 B.n751 VSUBS 0.007607f
C792 B.n752 VSUBS 0.007607f
C793 B.n753 VSUBS 0.007607f
C794 B.n754 VSUBS 0.007607f
C795 B.n755 VSUBS 0.007607f
C796 B.n756 VSUBS 0.007607f
C797 B.n757 VSUBS 0.007607f
C798 B.n758 VSUBS 0.007607f
C799 B.n759 VSUBS 0.007607f
C800 B.n760 VSUBS 0.007607f
C801 B.n761 VSUBS 0.007607f
C802 B.n762 VSUBS 0.007607f
C803 B.n763 VSUBS 0.007607f
C804 B.n764 VSUBS 0.007607f
C805 B.n765 VSUBS 0.007607f
C806 B.n766 VSUBS 0.007607f
C807 B.n767 VSUBS 0.007607f
C808 B.n768 VSUBS 0.007607f
C809 B.n769 VSUBS 0.007607f
C810 B.n770 VSUBS 0.007607f
C811 B.n771 VSUBS 0.007607f
C812 B.n772 VSUBS 0.007607f
C813 B.n773 VSUBS 0.007607f
C814 B.n774 VSUBS 0.007607f
C815 B.n775 VSUBS 0.007607f
C816 B.n776 VSUBS 0.007607f
C817 B.n777 VSUBS 0.007607f
C818 B.n778 VSUBS 0.007607f
C819 B.n779 VSUBS 0.007607f
C820 B.n780 VSUBS 0.007607f
C821 B.n781 VSUBS 0.007607f
C822 B.n782 VSUBS 0.007607f
C823 B.n783 VSUBS 0.007607f
C824 B.n784 VSUBS 0.007607f
C825 B.n785 VSUBS 0.007607f
C826 B.n786 VSUBS 0.007607f
C827 B.n787 VSUBS 0.007607f
C828 B.n788 VSUBS 0.007607f
C829 B.n789 VSUBS 0.007607f
C830 B.n790 VSUBS 0.007607f
C831 B.n791 VSUBS 0.007607f
C832 B.n792 VSUBS 0.007607f
C833 B.n793 VSUBS 0.007607f
C834 B.n794 VSUBS 0.007607f
C835 B.n795 VSUBS 0.007607f
C836 B.n796 VSUBS 0.007607f
C837 B.n797 VSUBS 0.007607f
C838 B.n798 VSUBS 0.007607f
C839 B.n799 VSUBS 0.007607f
C840 B.n800 VSUBS 0.007607f
C841 B.n801 VSUBS 0.007607f
C842 B.n802 VSUBS 0.007607f
C843 B.n803 VSUBS 0.007607f
C844 B.n804 VSUBS 0.007607f
C845 B.n805 VSUBS 0.007607f
C846 B.n806 VSUBS 0.007607f
C847 B.n807 VSUBS 0.007607f
C848 B.n808 VSUBS 0.007607f
C849 B.n809 VSUBS 0.007607f
C850 B.n810 VSUBS 0.007607f
C851 B.n811 VSUBS 0.007607f
C852 B.n812 VSUBS 0.007607f
C853 B.n813 VSUBS 0.007607f
C854 B.n814 VSUBS 0.007607f
C855 B.n815 VSUBS 0.007607f
C856 B.n816 VSUBS 0.007607f
C857 B.n817 VSUBS 0.007607f
C858 B.n818 VSUBS 0.007607f
C859 B.n819 VSUBS 0.007607f
C860 B.n820 VSUBS 0.007607f
C861 B.n821 VSUBS 0.007607f
C862 B.n822 VSUBS 0.007607f
C863 B.n823 VSUBS 0.007607f
C864 B.n824 VSUBS 0.007607f
C865 B.n825 VSUBS 0.007607f
C866 B.n826 VSUBS 0.007607f
C867 B.n827 VSUBS 0.007607f
C868 B.n828 VSUBS 0.007607f
C869 B.n829 VSUBS 0.007607f
C870 B.n830 VSUBS 0.007607f
C871 B.n831 VSUBS 0.009927f
C872 B.n832 VSUBS 0.010574f
C873 B.n833 VSUBS 0.021028f
C874 VDD2.t7 VSUBS 0.262528f
C875 VDD2.t0 VSUBS 0.262528f
C876 VDD2.n0 VSUBS 2.03969f
C877 VDD2.t4 VSUBS 0.262528f
C878 VDD2.t6 VSUBS 0.262528f
C879 VDD2.n1 VSUBS 2.03969f
C880 VDD2.n2 VSUBS 4.92506f
C881 VDD2.t2 VSUBS 0.262528f
C882 VDD2.t1 VSUBS 0.262528f
C883 VDD2.n3 VSUBS 2.02152f
C884 VDD2.n4 VSUBS 4.04908f
C885 VDD2.t3 VSUBS 0.262528f
C886 VDD2.t5 VSUBS 0.262528f
C887 VDD2.n5 VSUBS 2.03964f
C888 VN.t1 VSUBS 2.51724f
C889 VN.n0 VSUBS 1.00988f
C890 VN.n1 VSUBS 0.027192f
C891 VN.n2 VSUBS 0.038341f
C892 VN.n3 VSUBS 0.027192f
C893 VN.t3 VSUBS 2.51724f
C894 VN.n4 VSUBS 0.890897f
C895 VN.n5 VSUBS 0.027192f
C896 VN.n6 VSUBS 0.039868f
C897 VN.n7 VSUBS 0.309485f
C898 VN.t7 VSUBS 2.51724f
C899 VN.t0 VSUBS 2.83058f
C900 VN.n8 VSUBS 0.941011f
C901 VN.n9 VSUBS 0.994026f
C902 VN.n10 VSUBS 0.050429f
C903 VN.n11 VSUBS 0.050932f
C904 VN.n12 VSUBS 0.027192f
C905 VN.n13 VSUBS 0.027192f
C906 VN.n14 VSUBS 0.027192f
C907 VN.n15 VSUBS 0.039868f
C908 VN.n16 VSUBS 0.050932f
C909 VN.n17 VSUBS 0.050429f
C910 VN.n18 VSUBS 0.027192f
C911 VN.n19 VSUBS 0.027192f
C912 VN.n20 VSUBS 0.026288f
C913 VN.n21 VSUBS 0.050932f
C914 VN.n22 VSUBS 0.050932f
C915 VN.n23 VSUBS 0.027192f
C916 VN.n24 VSUBS 0.027192f
C917 VN.n25 VSUBS 0.027192f
C918 VN.n26 VSUBS 0.041394f
C919 VN.n27 VSUBS 0.050932f
C920 VN.n28 VSUBS 0.049424f
C921 VN.n29 VSUBS 0.043894f
C922 VN.n30 VSUBS 0.053802f
C923 VN.t5 VSUBS 2.51724f
C924 VN.n31 VSUBS 1.00988f
C925 VN.n32 VSUBS 0.027192f
C926 VN.n33 VSUBS 0.038341f
C927 VN.n34 VSUBS 0.027192f
C928 VN.t6 VSUBS 2.51724f
C929 VN.n35 VSUBS 0.890897f
C930 VN.n36 VSUBS 0.027192f
C931 VN.n37 VSUBS 0.039868f
C932 VN.n38 VSUBS 0.309485f
C933 VN.t4 VSUBS 2.51724f
C934 VN.t2 VSUBS 2.83058f
C935 VN.n39 VSUBS 0.941011f
C936 VN.n40 VSUBS 0.994026f
C937 VN.n41 VSUBS 0.050429f
C938 VN.n42 VSUBS 0.050932f
C939 VN.n43 VSUBS 0.027192f
C940 VN.n44 VSUBS 0.027192f
C941 VN.n45 VSUBS 0.027192f
C942 VN.n46 VSUBS 0.039868f
C943 VN.n47 VSUBS 0.050932f
C944 VN.n48 VSUBS 0.050429f
C945 VN.n49 VSUBS 0.027192f
C946 VN.n50 VSUBS 0.027192f
C947 VN.n51 VSUBS 0.026288f
C948 VN.n52 VSUBS 0.050932f
C949 VN.n53 VSUBS 0.050932f
C950 VN.n54 VSUBS 0.027192f
C951 VN.n55 VSUBS 0.027192f
C952 VN.n56 VSUBS 0.027192f
C953 VN.n57 VSUBS 0.041394f
C954 VN.n58 VSUBS 0.050932f
C955 VN.n59 VSUBS 0.049424f
C956 VN.n60 VSUBS 0.043894f
C957 VN.n61 VSUBS 1.67127f
C958 VDD1.t4 VSUBS 0.26363f
C959 VDD1.t1 VSUBS 0.26363f
C960 VDD1.n0 VSUBS 2.04988f
C961 VDD1.t3 VSUBS 0.26363f
C962 VDD1.t5 VSUBS 0.26363f
C963 VDD1.n1 VSUBS 2.04826f
C964 VDD1.t0 VSUBS 0.26363f
C965 VDD1.t6 VSUBS 0.26363f
C966 VDD1.n2 VSUBS 2.04826f
C967 VDD1.n3 VSUBS 5.00965f
C968 VDD1.t2 VSUBS 0.26363f
C969 VDD1.t7 VSUBS 0.26363f
C970 VDD1.n4 VSUBS 2.03f
C971 VDD1.n5 VSUBS 4.10452f
C972 VTAIL.t7 VSUBS 0.223339f
C973 VTAIL.t3 VSUBS 0.223339f
C974 VTAIL.n0 VSUBS 1.59396f
C975 VTAIL.n1 VSUBS 0.819501f
C976 VTAIL.n2 VSUBS 0.029256f
C977 VTAIL.n3 VSUBS 0.026121f
C978 VTAIL.n4 VSUBS 0.014036f
C979 VTAIL.n5 VSUBS 0.033176f
C980 VTAIL.n6 VSUBS 0.014862f
C981 VTAIL.n7 VSUBS 0.026121f
C982 VTAIL.n8 VSUBS 0.014036f
C983 VTAIL.n9 VSUBS 0.033176f
C984 VTAIL.n10 VSUBS 0.014862f
C985 VTAIL.n11 VSUBS 0.026121f
C986 VTAIL.n12 VSUBS 0.014036f
C987 VTAIL.n13 VSUBS 0.033176f
C988 VTAIL.n14 VSUBS 0.014862f
C989 VTAIL.n15 VSUBS 0.026121f
C990 VTAIL.n16 VSUBS 0.014036f
C991 VTAIL.n17 VSUBS 0.033176f
C992 VTAIL.n18 VSUBS 0.014862f
C993 VTAIL.n19 VSUBS 0.19179f
C994 VTAIL.t5 VSUBS 0.0714f
C995 VTAIL.n20 VSUBS 0.024882f
C996 VTAIL.n21 VSUBS 0.024957f
C997 VTAIL.n22 VSUBS 0.014036f
C998 VTAIL.n23 VSUBS 1.14831f
C999 VTAIL.n24 VSUBS 0.026121f
C1000 VTAIL.n25 VSUBS 0.014036f
C1001 VTAIL.n26 VSUBS 0.014862f
C1002 VTAIL.n27 VSUBS 0.033176f
C1003 VTAIL.n28 VSUBS 0.033176f
C1004 VTAIL.n29 VSUBS 0.014862f
C1005 VTAIL.n30 VSUBS 0.014036f
C1006 VTAIL.n31 VSUBS 0.026121f
C1007 VTAIL.n32 VSUBS 0.026121f
C1008 VTAIL.n33 VSUBS 0.014036f
C1009 VTAIL.n34 VSUBS 0.014862f
C1010 VTAIL.n35 VSUBS 0.033176f
C1011 VTAIL.n36 VSUBS 0.033176f
C1012 VTAIL.n37 VSUBS 0.033176f
C1013 VTAIL.n38 VSUBS 0.014862f
C1014 VTAIL.n39 VSUBS 0.014036f
C1015 VTAIL.n40 VSUBS 0.026121f
C1016 VTAIL.n41 VSUBS 0.026121f
C1017 VTAIL.n42 VSUBS 0.014036f
C1018 VTAIL.n43 VSUBS 0.014449f
C1019 VTAIL.n44 VSUBS 0.014449f
C1020 VTAIL.n45 VSUBS 0.033176f
C1021 VTAIL.n46 VSUBS 0.033176f
C1022 VTAIL.n47 VSUBS 0.014862f
C1023 VTAIL.n48 VSUBS 0.014036f
C1024 VTAIL.n49 VSUBS 0.026121f
C1025 VTAIL.n50 VSUBS 0.026121f
C1026 VTAIL.n51 VSUBS 0.014036f
C1027 VTAIL.n52 VSUBS 0.014862f
C1028 VTAIL.n53 VSUBS 0.033176f
C1029 VTAIL.n54 VSUBS 0.082207f
C1030 VTAIL.n55 VSUBS 0.014862f
C1031 VTAIL.n56 VSUBS 0.014036f
C1032 VTAIL.n57 VSUBS 0.065372f
C1033 VTAIL.n58 VSUBS 0.041573f
C1034 VTAIL.n59 VSUBS 0.317177f
C1035 VTAIL.n60 VSUBS 0.029256f
C1036 VTAIL.n61 VSUBS 0.026121f
C1037 VTAIL.n62 VSUBS 0.014036f
C1038 VTAIL.n63 VSUBS 0.033176f
C1039 VTAIL.n64 VSUBS 0.014862f
C1040 VTAIL.n65 VSUBS 0.026121f
C1041 VTAIL.n66 VSUBS 0.014036f
C1042 VTAIL.n67 VSUBS 0.033176f
C1043 VTAIL.n68 VSUBS 0.014862f
C1044 VTAIL.n69 VSUBS 0.026121f
C1045 VTAIL.n70 VSUBS 0.014036f
C1046 VTAIL.n71 VSUBS 0.033176f
C1047 VTAIL.n72 VSUBS 0.014862f
C1048 VTAIL.n73 VSUBS 0.026121f
C1049 VTAIL.n74 VSUBS 0.014036f
C1050 VTAIL.n75 VSUBS 0.033176f
C1051 VTAIL.n76 VSUBS 0.014862f
C1052 VTAIL.n77 VSUBS 0.19179f
C1053 VTAIL.t15 VSUBS 0.0714f
C1054 VTAIL.n78 VSUBS 0.024882f
C1055 VTAIL.n79 VSUBS 0.024957f
C1056 VTAIL.n80 VSUBS 0.014036f
C1057 VTAIL.n81 VSUBS 1.14831f
C1058 VTAIL.n82 VSUBS 0.026121f
C1059 VTAIL.n83 VSUBS 0.014036f
C1060 VTAIL.n84 VSUBS 0.014862f
C1061 VTAIL.n85 VSUBS 0.033176f
C1062 VTAIL.n86 VSUBS 0.033176f
C1063 VTAIL.n87 VSUBS 0.014862f
C1064 VTAIL.n88 VSUBS 0.014036f
C1065 VTAIL.n89 VSUBS 0.026121f
C1066 VTAIL.n90 VSUBS 0.026121f
C1067 VTAIL.n91 VSUBS 0.014036f
C1068 VTAIL.n92 VSUBS 0.014862f
C1069 VTAIL.n93 VSUBS 0.033176f
C1070 VTAIL.n94 VSUBS 0.033176f
C1071 VTAIL.n95 VSUBS 0.033176f
C1072 VTAIL.n96 VSUBS 0.014862f
C1073 VTAIL.n97 VSUBS 0.014036f
C1074 VTAIL.n98 VSUBS 0.026121f
C1075 VTAIL.n99 VSUBS 0.026121f
C1076 VTAIL.n100 VSUBS 0.014036f
C1077 VTAIL.n101 VSUBS 0.014449f
C1078 VTAIL.n102 VSUBS 0.014449f
C1079 VTAIL.n103 VSUBS 0.033176f
C1080 VTAIL.n104 VSUBS 0.033176f
C1081 VTAIL.n105 VSUBS 0.014862f
C1082 VTAIL.n106 VSUBS 0.014036f
C1083 VTAIL.n107 VSUBS 0.026121f
C1084 VTAIL.n108 VSUBS 0.026121f
C1085 VTAIL.n109 VSUBS 0.014036f
C1086 VTAIL.n110 VSUBS 0.014862f
C1087 VTAIL.n111 VSUBS 0.033176f
C1088 VTAIL.n112 VSUBS 0.082207f
C1089 VTAIL.n113 VSUBS 0.014862f
C1090 VTAIL.n114 VSUBS 0.014036f
C1091 VTAIL.n115 VSUBS 0.065372f
C1092 VTAIL.n116 VSUBS 0.041573f
C1093 VTAIL.n117 VSUBS 0.317177f
C1094 VTAIL.t8 VSUBS 0.223339f
C1095 VTAIL.t13 VSUBS 0.223339f
C1096 VTAIL.n118 VSUBS 1.59396f
C1097 VTAIL.n119 VSUBS 1.0671f
C1098 VTAIL.n120 VSUBS 0.029256f
C1099 VTAIL.n121 VSUBS 0.026121f
C1100 VTAIL.n122 VSUBS 0.014036f
C1101 VTAIL.n123 VSUBS 0.033176f
C1102 VTAIL.n124 VSUBS 0.014862f
C1103 VTAIL.n125 VSUBS 0.026121f
C1104 VTAIL.n126 VSUBS 0.014036f
C1105 VTAIL.n127 VSUBS 0.033176f
C1106 VTAIL.n128 VSUBS 0.014862f
C1107 VTAIL.n129 VSUBS 0.026121f
C1108 VTAIL.n130 VSUBS 0.014036f
C1109 VTAIL.n131 VSUBS 0.033176f
C1110 VTAIL.n132 VSUBS 0.014862f
C1111 VTAIL.n133 VSUBS 0.026121f
C1112 VTAIL.n134 VSUBS 0.014036f
C1113 VTAIL.n135 VSUBS 0.033176f
C1114 VTAIL.n136 VSUBS 0.014862f
C1115 VTAIL.n137 VSUBS 0.19179f
C1116 VTAIL.t9 VSUBS 0.0714f
C1117 VTAIL.n138 VSUBS 0.024882f
C1118 VTAIL.n139 VSUBS 0.024957f
C1119 VTAIL.n140 VSUBS 0.014036f
C1120 VTAIL.n141 VSUBS 1.14831f
C1121 VTAIL.n142 VSUBS 0.026121f
C1122 VTAIL.n143 VSUBS 0.014036f
C1123 VTAIL.n144 VSUBS 0.014862f
C1124 VTAIL.n145 VSUBS 0.033176f
C1125 VTAIL.n146 VSUBS 0.033176f
C1126 VTAIL.n147 VSUBS 0.014862f
C1127 VTAIL.n148 VSUBS 0.014036f
C1128 VTAIL.n149 VSUBS 0.026121f
C1129 VTAIL.n150 VSUBS 0.026121f
C1130 VTAIL.n151 VSUBS 0.014036f
C1131 VTAIL.n152 VSUBS 0.014862f
C1132 VTAIL.n153 VSUBS 0.033176f
C1133 VTAIL.n154 VSUBS 0.033176f
C1134 VTAIL.n155 VSUBS 0.033176f
C1135 VTAIL.n156 VSUBS 0.014862f
C1136 VTAIL.n157 VSUBS 0.014036f
C1137 VTAIL.n158 VSUBS 0.026121f
C1138 VTAIL.n159 VSUBS 0.026121f
C1139 VTAIL.n160 VSUBS 0.014036f
C1140 VTAIL.n161 VSUBS 0.014449f
C1141 VTAIL.n162 VSUBS 0.014449f
C1142 VTAIL.n163 VSUBS 0.033176f
C1143 VTAIL.n164 VSUBS 0.033176f
C1144 VTAIL.n165 VSUBS 0.014862f
C1145 VTAIL.n166 VSUBS 0.014036f
C1146 VTAIL.n167 VSUBS 0.026121f
C1147 VTAIL.n168 VSUBS 0.026121f
C1148 VTAIL.n169 VSUBS 0.014036f
C1149 VTAIL.n170 VSUBS 0.014862f
C1150 VTAIL.n171 VSUBS 0.033176f
C1151 VTAIL.n172 VSUBS 0.082207f
C1152 VTAIL.n173 VSUBS 0.014862f
C1153 VTAIL.n174 VSUBS 0.014036f
C1154 VTAIL.n175 VSUBS 0.065372f
C1155 VTAIL.n176 VSUBS 0.041573f
C1156 VTAIL.n177 VSUBS 1.67002f
C1157 VTAIL.n178 VSUBS 0.029256f
C1158 VTAIL.n179 VSUBS 0.026121f
C1159 VTAIL.n180 VSUBS 0.014036f
C1160 VTAIL.n181 VSUBS 0.033176f
C1161 VTAIL.n182 VSUBS 0.014862f
C1162 VTAIL.n183 VSUBS 0.026121f
C1163 VTAIL.n184 VSUBS 0.014036f
C1164 VTAIL.n185 VSUBS 0.033176f
C1165 VTAIL.n186 VSUBS 0.014862f
C1166 VTAIL.n187 VSUBS 0.026121f
C1167 VTAIL.n188 VSUBS 0.014036f
C1168 VTAIL.n189 VSUBS 0.033176f
C1169 VTAIL.n190 VSUBS 0.033176f
C1170 VTAIL.n191 VSUBS 0.014862f
C1171 VTAIL.n192 VSUBS 0.026121f
C1172 VTAIL.n193 VSUBS 0.014036f
C1173 VTAIL.n194 VSUBS 0.033176f
C1174 VTAIL.n195 VSUBS 0.014862f
C1175 VTAIL.n196 VSUBS 0.19179f
C1176 VTAIL.t4 VSUBS 0.0714f
C1177 VTAIL.n197 VSUBS 0.024882f
C1178 VTAIL.n198 VSUBS 0.024957f
C1179 VTAIL.n199 VSUBS 0.014036f
C1180 VTAIL.n200 VSUBS 1.14831f
C1181 VTAIL.n201 VSUBS 0.026121f
C1182 VTAIL.n202 VSUBS 0.014036f
C1183 VTAIL.n203 VSUBS 0.014862f
C1184 VTAIL.n204 VSUBS 0.033176f
C1185 VTAIL.n205 VSUBS 0.033176f
C1186 VTAIL.n206 VSUBS 0.014862f
C1187 VTAIL.n207 VSUBS 0.014036f
C1188 VTAIL.n208 VSUBS 0.026121f
C1189 VTAIL.n209 VSUBS 0.026121f
C1190 VTAIL.n210 VSUBS 0.014036f
C1191 VTAIL.n211 VSUBS 0.014862f
C1192 VTAIL.n212 VSUBS 0.033176f
C1193 VTAIL.n213 VSUBS 0.033176f
C1194 VTAIL.n214 VSUBS 0.014862f
C1195 VTAIL.n215 VSUBS 0.014036f
C1196 VTAIL.n216 VSUBS 0.026121f
C1197 VTAIL.n217 VSUBS 0.026121f
C1198 VTAIL.n218 VSUBS 0.014036f
C1199 VTAIL.n219 VSUBS 0.014449f
C1200 VTAIL.n220 VSUBS 0.014449f
C1201 VTAIL.n221 VSUBS 0.033176f
C1202 VTAIL.n222 VSUBS 0.033176f
C1203 VTAIL.n223 VSUBS 0.014862f
C1204 VTAIL.n224 VSUBS 0.014036f
C1205 VTAIL.n225 VSUBS 0.026121f
C1206 VTAIL.n226 VSUBS 0.026121f
C1207 VTAIL.n227 VSUBS 0.014036f
C1208 VTAIL.n228 VSUBS 0.014862f
C1209 VTAIL.n229 VSUBS 0.033176f
C1210 VTAIL.n230 VSUBS 0.082207f
C1211 VTAIL.n231 VSUBS 0.014862f
C1212 VTAIL.n232 VSUBS 0.014036f
C1213 VTAIL.n233 VSUBS 0.065372f
C1214 VTAIL.n234 VSUBS 0.041573f
C1215 VTAIL.n235 VSUBS 1.67002f
C1216 VTAIL.t1 VSUBS 0.223339f
C1217 VTAIL.t2 VSUBS 0.223339f
C1218 VTAIL.n236 VSUBS 1.59397f
C1219 VTAIL.n237 VSUBS 1.06709f
C1220 VTAIL.n238 VSUBS 0.029256f
C1221 VTAIL.n239 VSUBS 0.026121f
C1222 VTAIL.n240 VSUBS 0.014036f
C1223 VTAIL.n241 VSUBS 0.033176f
C1224 VTAIL.n242 VSUBS 0.014862f
C1225 VTAIL.n243 VSUBS 0.026121f
C1226 VTAIL.n244 VSUBS 0.014036f
C1227 VTAIL.n245 VSUBS 0.033176f
C1228 VTAIL.n246 VSUBS 0.014862f
C1229 VTAIL.n247 VSUBS 0.026121f
C1230 VTAIL.n248 VSUBS 0.014036f
C1231 VTAIL.n249 VSUBS 0.033176f
C1232 VTAIL.n250 VSUBS 0.033176f
C1233 VTAIL.n251 VSUBS 0.014862f
C1234 VTAIL.n252 VSUBS 0.026121f
C1235 VTAIL.n253 VSUBS 0.014036f
C1236 VTAIL.n254 VSUBS 0.033176f
C1237 VTAIL.n255 VSUBS 0.014862f
C1238 VTAIL.n256 VSUBS 0.19179f
C1239 VTAIL.t6 VSUBS 0.0714f
C1240 VTAIL.n257 VSUBS 0.024882f
C1241 VTAIL.n258 VSUBS 0.024957f
C1242 VTAIL.n259 VSUBS 0.014036f
C1243 VTAIL.n260 VSUBS 1.14831f
C1244 VTAIL.n261 VSUBS 0.026121f
C1245 VTAIL.n262 VSUBS 0.014036f
C1246 VTAIL.n263 VSUBS 0.014862f
C1247 VTAIL.n264 VSUBS 0.033176f
C1248 VTAIL.n265 VSUBS 0.033176f
C1249 VTAIL.n266 VSUBS 0.014862f
C1250 VTAIL.n267 VSUBS 0.014036f
C1251 VTAIL.n268 VSUBS 0.026121f
C1252 VTAIL.n269 VSUBS 0.026121f
C1253 VTAIL.n270 VSUBS 0.014036f
C1254 VTAIL.n271 VSUBS 0.014862f
C1255 VTAIL.n272 VSUBS 0.033176f
C1256 VTAIL.n273 VSUBS 0.033176f
C1257 VTAIL.n274 VSUBS 0.014862f
C1258 VTAIL.n275 VSUBS 0.014036f
C1259 VTAIL.n276 VSUBS 0.026121f
C1260 VTAIL.n277 VSUBS 0.026121f
C1261 VTAIL.n278 VSUBS 0.014036f
C1262 VTAIL.n279 VSUBS 0.014449f
C1263 VTAIL.n280 VSUBS 0.014449f
C1264 VTAIL.n281 VSUBS 0.033176f
C1265 VTAIL.n282 VSUBS 0.033176f
C1266 VTAIL.n283 VSUBS 0.014862f
C1267 VTAIL.n284 VSUBS 0.014036f
C1268 VTAIL.n285 VSUBS 0.026121f
C1269 VTAIL.n286 VSUBS 0.026121f
C1270 VTAIL.n287 VSUBS 0.014036f
C1271 VTAIL.n288 VSUBS 0.014862f
C1272 VTAIL.n289 VSUBS 0.033176f
C1273 VTAIL.n290 VSUBS 0.082207f
C1274 VTAIL.n291 VSUBS 0.014862f
C1275 VTAIL.n292 VSUBS 0.014036f
C1276 VTAIL.n293 VSUBS 0.065372f
C1277 VTAIL.n294 VSUBS 0.041573f
C1278 VTAIL.n295 VSUBS 0.317177f
C1279 VTAIL.n296 VSUBS 0.029256f
C1280 VTAIL.n297 VSUBS 0.026121f
C1281 VTAIL.n298 VSUBS 0.014036f
C1282 VTAIL.n299 VSUBS 0.033176f
C1283 VTAIL.n300 VSUBS 0.014862f
C1284 VTAIL.n301 VSUBS 0.026121f
C1285 VTAIL.n302 VSUBS 0.014036f
C1286 VTAIL.n303 VSUBS 0.033176f
C1287 VTAIL.n304 VSUBS 0.014862f
C1288 VTAIL.n305 VSUBS 0.026121f
C1289 VTAIL.n306 VSUBS 0.014036f
C1290 VTAIL.n307 VSUBS 0.033176f
C1291 VTAIL.n308 VSUBS 0.033176f
C1292 VTAIL.n309 VSUBS 0.014862f
C1293 VTAIL.n310 VSUBS 0.026121f
C1294 VTAIL.n311 VSUBS 0.014036f
C1295 VTAIL.n312 VSUBS 0.033176f
C1296 VTAIL.n313 VSUBS 0.014862f
C1297 VTAIL.n314 VSUBS 0.19179f
C1298 VTAIL.t11 VSUBS 0.0714f
C1299 VTAIL.n315 VSUBS 0.024882f
C1300 VTAIL.n316 VSUBS 0.024957f
C1301 VTAIL.n317 VSUBS 0.014036f
C1302 VTAIL.n318 VSUBS 1.14831f
C1303 VTAIL.n319 VSUBS 0.026121f
C1304 VTAIL.n320 VSUBS 0.014036f
C1305 VTAIL.n321 VSUBS 0.014862f
C1306 VTAIL.n322 VSUBS 0.033176f
C1307 VTAIL.n323 VSUBS 0.033176f
C1308 VTAIL.n324 VSUBS 0.014862f
C1309 VTAIL.n325 VSUBS 0.014036f
C1310 VTAIL.n326 VSUBS 0.026121f
C1311 VTAIL.n327 VSUBS 0.026121f
C1312 VTAIL.n328 VSUBS 0.014036f
C1313 VTAIL.n329 VSUBS 0.014862f
C1314 VTAIL.n330 VSUBS 0.033176f
C1315 VTAIL.n331 VSUBS 0.033176f
C1316 VTAIL.n332 VSUBS 0.014862f
C1317 VTAIL.n333 VSUBS 0.014036f
C1318 VTAIL.n334 VSUBS 0.026121f
C1319 VTAIL.n335 VSUBS 0.026121f
C1320 VTAIL.n336 VSUBS 0.014036f
C1321 VTAIL.n337 VSUBS 0.014449f
C1322 VTAIL.n338 VSUBS 0.014449f
C1323 VTAIL.n339 VSUBS 0.033176f
C1324 VTAIL.n340 VSUBS 0.033176f
C1325 VTAIL.n341 VSUBS 0.014862f
C1326 VTAIL.n342 VSUBS 0.014036f
C1327 VTAIL.n343 VSUBS 0.026121f
C1328 VTAIL.n344 VSUBS 0.026121f
C1329 VTAIL.n345 VSUBS 0.014036f
C1330 VTAIL.n346 VSUBS 0.014862f
C1331 VTAIL.n347 VSUBS 0.033176f
C1332 VTAIL.n348 VSUBS 0.082207f
C1333 VTAIL.n349 VSUBS 0.014862f
C1334 VTAIL.n350 VSUBS 0.014036f
C1335 VTAIL.n351 VSUBS 0.065372f
C1336 VTAIL.n352 VSUBS 0.041573f
C1337 VTAIL.n353 VSUBS 0.317177f
C1338 VTAIL.t10 VSUBS 0.223339f
C1339 VTAIL.t14 VSUBS 0.223339f
C1340 VTAIL.n354 VSUBS 1.59397f
C1341 VTAIL.n355 VSUBS 1.06709f
C1342 VTAIL.n356 VSUBS 0.029256f
C1343 VTAIL.n357 VSUBS 0.026121f
C1344 VTAIL.n358 VSUBS 0.014036f
C1345 VTAIL.n359 VSUBS 0.033176f
C1346 VTAIL.n360 VSUBS 0.014862f
C1347 VTAIL.n361 VSUBS 0.026121f
C1348 VTAIL.n362 VSUBS 0.014036f
C1349 VTAIL.n363 VSUBS 0.033176f
C1350 VTAIL.n364 VSUBS 0.014862f
C1351 VTAIL.n365 VSUBS 0.026121f
C1352 VTAIL.n366 VSUBS 0.014036f
C1353 VTAIL.n367 VSUBS 0.033176f
C1354 VTAIL.n368 VSUBS 0.033176f
C1355 VTAIL.n369 VSUBS 0.014862f
C1356 VTAIL.n370 VSUBS 0.026121f
C1357 VTAIL.n371 VSUBS 0.014036f
C1358 VTAIL.n372 VSUBS 0.033176f
C1359 VTAIL.n373 VSUBS 0.014862f
C1360 VTAIL.n374 VSUBS 0.19179f
C1361 VTAIL.t12 VSUBS 0.0714f
C1362 VTAIL.n375 VSUBS 0.024882f
C1363 VTAIL.n376 VSUBS 0.024957f
C1364 VTAIL.n377 VSUBS 0.014036f
C1365 VTAIL.n378 VSUBS 1.14831f
C1366 VTAIL.n379 VSUBS 0.026121f
C1367 VTAIL.n380 VSUBS 0.014036f
C1368 VTAIL.n381 VSUBS 0.014862f
C1369 VTAIL.n382 VSUBS 0.033176f
C1370 VTAIL.n383 VSUBS 0.033176f
C1371 VTAIL.n384 VSUBS 0.014862f
C1372 VTAIL.n385 VSUBS 0.014036f
C1373 VTAIL.n386 VSUBS 0.026121f
C1374 VTAIL.n387 VSUBS 0.026121f
C1375 VTAIL.n388 VSUBS 0.014036f
C1376 VTAIL.n389 VSUBS 0.014862f
C1377 VTAIL.n390 VSUBS 0.033176f
C1378 VTAIL.n391 VSUBS 0.033176f
C1379 VTAIL.n392 VSUBS 0.014862f
C1380 VTAIL.n393 VSUBS 0.014036f
C1381 VTAIL.n394 VSUBS 0.026121f
C1382 VTAIL.n395 VSUBS 0.026121f
C1383 VTAIL.n396 VSUBS 0.014036f
C1384 VTAIL.n397 VSUBS 0.014449f
C1385 VTAIL.n398 VSUBS 0.014449f
C1386 VTAIL.n399 VSUBS 0.033176f
C1387 VTAIL.n400 VSUBS 0.033176f
C1388 VTAIL.n401 VSUBS 0.014862f
C1389 VTAIL.n402 VSUBS 0.014036f
C1390 VTAIL.n403 VSUBS 0.026121f
C1391 VTAIL.n404 VSUBS 0.026121f
C1392 VTAIL.n405 VSUBS 0.014036f
C1393 VTAIL.n406 VSUBS 0.014862f
C1394 VTAIL.n407 VSUBS 0.033176f
C1395 VTAIL.n408 VSUBS 0.082207f
C1396 VTAIL.n409 VSUBS 0.014862f
C1397 VTAIL.n410 VSUBS 0.014036f
C1398 VTAIL.n411 VSUBS 0.065372f
C1399 VTAIL.n412 VSUBS 0.041573f
C1400 VTAIL.n413 VSUBS 1.67002f
C1401 VTAIL.n414 VSUBS 0.029256f
C1402 VTAIL.n415 VSUBS 0.026121f
C1403 VTAIL.n416 VSUBS 0.014036f
C1404 VTAIL.n417 VSUBS 0.033176f
C1405 VTAIL.n418 VSUBS 0.014862f
C1406 VTAIL.n419 VSUBS 0.026121f
C1407 VTAIL.n420 VSUBS 0.014036f
C1408 VTAIL.n421 VSUBS 0.033176f
C1409 VTAIL.n422 VSUBS 0.014862f
C1410 VTAIL.n423 VSUBS 0.026121f
C1411 VTAIL.n424 VSUBS 0.014036f
C1412 VTAIL.n425 VSUBS 0.033176f
C1413 VTAIL.n426 VSUBS 0.014862f
C1414 VTAIL.n427 VSUBS 0.026121f
C1415 VTAIL.n428 VSUBS 0.014036f
C1416 VTAIL.n429 VSUBS 0.033176f
C1417 VTAIL.n430 VSUBS 0.014862f
C1418 VTAIL.n431 VSUBS 0.19179f
C1419 VTAIL.t0 VSUBS 0.0714f
C1420 VTAIL.n432 VSUBS 0.024882f
C1421 VTAIL.n433 VSUBS 0.024957f
C1422 VTAIL.n434 VSUBS 0.014036f
C1423 VTAIL.n435 VSUBS 1.14831f
C1424 VTAIL.n436 VSUBS 0.026121f
C1425 VTAIL.n437 VSUBS 0.014036f
C1426 VTAIL.n438 VSUBS 0.014862f
C1427 VTAIL.n439 VSUBS 0.033176f
C1428 VTAIL.n440 VSUBS 0.033176f
C1429 VTAIL.n441 VSUBS 0.014862f
C1430 VTAIL.n442 VSUBS 0.014036f
C1431 VTAIL.n443 VSUBS 0.026121f
C1432 VTAIL.n444 VSUBS 0.026121f
C1433 VTAIL.n445 VSUBS 0.014036f
C1434 VTAIL.n446 VSUBS 0.014862f
C1435 VTAIL.n447 VSUBS 0.033176f
C1436 VTAIL.n448 VSUBS 0.033176f
C1437 VTAIL.n449 VSUBS 0.033176f
C1438 VTAIL.n450 VSUBS 0.014862f
C1439 VTAIL.n451 VSUBS 0.014036f
C1440 VTAIL.n452 VSUBS 0.026121f
C1441 VTAIL.n453 VSUBS 0.026121f
C1442 VTAIL.n454 VSUBS 0.014036f
C1443 VTAIL.n455 VSUBS 0.014449f
C1444 VTAIL.n456 VSUBS 0.014449f
C1445 VTAIL.n457 VSUBS 0.033176f
C1446 VTAIL.n458 VSUBS 0.033176f
C1447 VTAIL.n459 VSUBS 0.014862f
C1448 VTAIL.n460 VSUBS 0.014036f
C1449 VTAIL.n461 VSUBS 0.026121f
C1450 VTAIL.n462 VSUBS 0.026121f
C1451 VTAIL.n463 VSUBS 0.014036f
C1452 VTAIL.n464 VSUBS 0.014862f
C1453 VTAIL.n465 VSUBS 0.033176f
C1454 VTAIL.n466 VSUBS 0.082207f
C1455 VTAIL.n467 VSUBS 0.014862f
C1456 VTAIL.n468 VSUBS 0.014036f
C1457 VTAIL.n469 VSUBS 0.065372f
C1458 VTAIL.n470 VSUBS 0.041573f
C1459 VTAIL.n471 VSUBS 1.66512f
C1460 VP.t1 VSUBS 2.7625f
C1461 VP.n0 VSUBS 1.10828f
C1462 VP.n1 VSUBS 0.029841f
C1463 VP.n2 VSUBS 0.042077f
C1464 VP.n3 VSUBS 0.029841f
C1465 VP.t7 VSUBS 2.7625f
C1466 VP.n4 VSUBS 0.9777f
C1467 VP.n5 VSUBS 0.029841f
C1468 VP.n6 VSUBS 0.043752f
C1469 VP.n7 VSUBS 0.029841f
C1470 VP.t2 VSUBS 2.7625f
C1471 VP.n8 VSUBS 0.055895f
C1472 VP.n9 VSUBS 0.029841f
C1473 VP.n10 VSUBS 0.055895f
C1474 VP.t0 VSUBS 2.7625f
C1475 VP.n11 VSUBS 1.10828f
C1476 VP.n12 VSUBS 0.029841f
C1477 VP.n13 VSUBS 0.042077f
C1478 VP.n14 VSUBS 0.029841f
C1479 VP.t5 VSUBS 2.7625f
C1480 VP.n15 VSUBS 0.9777f
C1481 VP.n16 VSUBS 0.029841f
C1482 VP.n17 VSUBS 0.043752f
C1483 VP.n18 VSUBS 0.33964f
C1484 VP.t6 VSUBS 2.7625f
C1485 VP.t3 VSUBS 3.10637f
C1486 VP.n19 VSUBS 1.0327f
C1487 VP.n20 VSUBS 1.09088f
C1488 VP.n21 VSUBS 0.055343f
C1489 VP.n22 VSUBS 0.055895f
C1490 VP.n23 VSUBS 0.029841f
C1491 VP.n24 VSUBS 0.029841f
C1492 VP.n25 VSUBS 0.029841f
C1493 VP.n26 VSUBS 0.043752f
C1494 VP.n27 VSUBS 0.055895f
C1495 VP.n28 VSUBS 0.055343f
C1496 VP.n29 VSUBS 0.029841f
C1497 VP.n30 VSUBS 0.029841f
C1498 VP.n31 VSUBS 0.028849f
C1499 VP.n32 VSUBS 0.055895f
C1500 VP.n33 VSUBS 0.055895f
C1501 VP.n34 VSUBS 0.029841f
C1502 VP.n35 VSUBS 0.029841f
C1503 VP.n36 VSUBS 0.029841f
C1504 VP.n37 VSUBS 0.045427f
C1505 VP.n38 VSUBS 0.055895f
C1506 VP.n39 VSUBS 0.054239f
C1507 VP.n40 VSUBS 0.04817f
C1508 VP.n41 VSUBS 1.82213f
C1509 VP.n42 VSUBS 1.84239f
C1510 VP.t4 VSUBS 2.7625f
C1511 VP.n43 VSUBS 1.10828f
C1512 VP.n44 VSUBS 0.054239f
C1513 VP.n45 VSUBS 0.04817f
C1514 VP.n46 VSUBS 0.029841f
C1515 VP.n47 VSUBS 0.029841f
C1516 VP.n48 VSUBS 0.045427f
C1517 VP.n49 VSUBS 0.042077f
C1518 VP.n50 VSUBS 0.055895f
C1519 VP.n51 VSUBS 0.029841f
C1520 VP.n52 VSUBS 0.029841f
C1521 VP.n53 VSUBS 0.029841f
C1522 VP.n54 VSUBS 0.028849f
C1523 VP.n55 VSUBS 0.9777f
C1524 VP.n56 VSUBS 0.055343f
C1525 VP.n57 VSUBS 0.055895f
C1526 VP.n58 VSUBS 0.029841f
C1527 VP.n59 VSUBS 0.029841f
C1528 VP.n60 VSUBS 0.029841f
C1529 VP.n61 VSUBS 0.043752f
C1530 VP.n62 VSUBS 0.055895f
C1531 VP.n63 VSUBS 0.055343f
C1532 VP.n64 VSUBS 0.029841f
C1533 VP.n65 VSUBS 0.029841f
C1534 VP.n66 VSUBS 0.028849f
C1535 VP.n67 VSUBS 0.055895f
C1536 VP.n68 VSUBS 0.055895f
C1537 VP.n69 VSUBS 0.029841f
C1538 VP.n70 VSUBS 0.029841f
C1539 VP.n71 VSUBS 0.029841f
C1540 VP.n72 VSUBS 0.045427f
C1541 VP.n73 VSUBS 0.055895f
C1542 VP.n74 VSUBS 0.054239f
C1543 VP.n75 VSUBS 0.04817f
C1544 VP.n76 VSUBS 0.059044f
.ends

