* NGSPICE file created from diff_pair_sample_0633.ext - technology: sky130A

.subckt diff_pair_sample_0633 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=5.7291 ps=30.16 w=14.69 l=1.81
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=5.7291 ps=30.16 w=14.69 l=1.81
X2 VDD2.t0 VN.t1 VTAIL.t1 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=5.7291 ps=30.16 w=14.69 l=1.81
X3 VDD1.t0 VP.t1 VTAIL.t2 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=5.7291 ps=30.16 w=14.69 l=1.81
X4 B.t11 B.t9 B.t10 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=0 ps=0 w=14.69 l=1.81
X5 B.t8 B.t6 B.t7 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=0 ps=0 w=14.69 l=1.81
X6 B.t5 B.t3 B.t4 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=0 ps=0 w=14.69 l=1.81
X7 B.t2 B.t0 B.t1 w_n1826_n3906# sky130_fd_pr__pfet_01v8 ad=5.7291 pd=30.16 as=0 ps=0 w=14.69 l=1.81
R0 VP.n0 VP.t1 299.057
R1 VP.n0 VP.t0 254.458
R2 VP VP.n0 0.241678
R3 VTAIL.n322 VTAIL.n246 756.745
R4 VTAIL.n76 VTAIL.n0 756.745
R5 VTAIL.n240 VTAIL.n164 756.745
R6 VTAIL.n158 VTAIL.n82 756.745
R7 VTAIL.n273 VTAIL.n272 585
R8 VTAIL.n270 VTAIL.n269 585
R9 VTAIL.n279 VTAIL.n278 585
R10 VTAIL.n281 VTAIL.n280 585
R11 VTAIL.n266 VTAIL.n265 585
R12 VTAIL.n287 VTAIL.n286 585
R13 VTAIL.n289 VTAIL.n288 585
R14 VTAIL.n262 VTAIL.n261 585
R15 VTAIL.n295 VTAIL.n294 585
R16 VTAIL.n297 VTAIL.n296 585
R17 VTAIL.n258 VTAIL.n257 585
R18 VTAIL.n303 VTAIL.n302 585
R19 VTAIL.n305 VTAIL.n304 585
R20 VTAIL.n254 VTAIL.n253 585
R21 VTAIL.n311 VTAIL.n310 585
R22 VTAIL.n314 VTAIL.n313 585
R23 VTAIL.n312 VTAIL.n250 585
R24 VTAIL.n319 VTAIL.n249 585
R25 VTAIL.n321 VTAIL.n320 585
R26 VTAIL.n323 VTAIL.n322 585
R27 VTAIL.n27 VTAIL.n26 585
R28 VTAIL.n24 VTAIL.n23 585
R29 VTAIL.n33 VTAIL.n32 585
R30 VTAIL.n35 VTAIL.n34 585
R31 VTAIL.n20 VTAIL.n19 585
R32 VTAIL.n41 VTAIL.n40 585
R33 VTAIL.n43 VTAIL.n42 585
R34 VTAIL.n16 VTAIL.n15 585
R35 VTAIL.n49 VTAIL.n48 585
R36 VTAIL.n51 VTAIL.n50 585
R37 VTAIL.n12 VTAIL.n11 585
R38 VTAIL.n57 VTAIL.n56 585
R39 VTAIL.n59 VTAIL.n58 585
R40 VTAIL.n8 VTAIL.n7 585
R41 VTAIL.n65 VTAIL.n64 585
R42 VTAIL.n68 VTAIL.n67 585
R43 VTAIL.n66 VTAIL.n4 585
R44 VTAIL.n73 VTAIL.n3 585
R45 VTAIL.n75 VTAIL.n74 585
R46 VTAIL.n77 VTAIL.n76 585
R47 VTAIL.n241 VTAIL.n240 585
R48 VTAIL.n239 VTAIL.n238 585
R49 VTAIL.n237 VTAIL.n167 585
R50 VTAIL.n171 VTAIL.n168 585
R51 VTAIL.n232 VTAIL.n231 585
R52 VTAIL.n230 VTAIL.n229 585
R53 VTAIL.n173 VTAIL.n172 585
R54 VTAIL.n224 VTAIL.n223 585
R55 VTAIL.n222 VTAIL.n221 585
R56 VTAIL.n177 VTAIL.n176 585
R57 VTAIL.n216 VTAIL.n215 585
R58 VTAIL.n214 VTAIL.n213 585
R59 VTAIL.n181 VTAIL.n180 585
R60 VTAIL.n208 VTAIL.n207 585
R61 VTAIL.n206 VTAIL.n205 585
R62 VTAIL.n185 VTAIL.n184 585
R63 VTAIL.n200 VTAIL.n199 585
R64 VTAIL.n198 VTAIL.n197 585
R65 VTAIL.n189 VTAIL.n188 585
R66 VTAIL.n192 VTAIL.n191 585
R67 VTAIL.n159 VTAIL.n158 585
R68 VTAIL.n157 VTAIL.n156 585
R69 VTAIL.n155 VTAIL.n85 585
R70 VTAIL.n89 VTAIL.n86 585
R71 VTAIL.n150 VTAIL.n149 585
R72 VTAIL.n148 VTAIL.n147 585
R73 VTAIL.n91 VTAIL.n90 585
R74 VTAIL.n142 VTAIL.n141 585
R75 VTAIL.n140 VTAIL.n139 585
R76 VTAIL.n95 VTAIL.n94 585
R77 VTAIL.n134 VTAIL.n133 585
R78 VTAIL.n132 VTAIL.n131 585
R79 VTAIL.n99 VTAIL.n98 585
R80 VTAIL.n126 VTAIL.n125 585
R81 VTAIL.n124 VTAIL.n123 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n118 VTAIL.n117 585
R84 VTAIL.n116 VTAIL.n115 585
R85 VTAIL.n107 VTAIL.n106 585
R86 VTAIL.n110 VTAIL.n109 585
R87 VTAIL.t2 VTAIL.n190 327.466
R88 VTAIL.t1 VTAIL.n108 327.466
R89 VTAIL.t0 VTAIL.n271 327.466
R90 VTAIL.t3 VTAIL.n25 327.466
R91 VTAIL.n272 VTAIL.n269 171.744
R92 VTAIL.n279 VTAIL.n269 171.744
R93 VTAIL.n280 VTAIL.n279 171.744
R94 VTAIL.n280 VTAIL.n265 171.744
R95 VTAIL.n287 VTAIL.n265 171.744
R96 VTAIL.n288 VTAIL.n287 171.744
R97 VTAIL.n288 VTAIL.n261 171.744
R98 VTAIL.n295 VTAIL.n261 171.744
R99 VTAIL.n296 VTAIL.n295 171.744
R100 VTAIL.n296 VTAIL.n257 171.744
R101 VTAIL.n303 VTAIL.n257 171.744
R102 VTAIL.n304 VTAIL.n303 171.744
R103 VTAIL.n304 VTAIL.n253 171.744
R104 VTAIL.n311 VTAIL.n253 171.744
R105 VTAIL.n313 VTAIL.n311 171.744
R106 VTAIL.n313 VTAIL.n312 171.744
R107 VTAIL.n312 VTAIL.n249 171.744
R108 VTAIL.n321 VTAIL.n249 171.744
R109 VTAIL.n322 VTAIL.n321 171.744
R110 VTAIL.n26 VTAIL.n23 171.744
R111 VTAIL.n33 VTAIL.n23 171.744
R112 VTAIL.n34 VTAIL.n33 171.744
R113 VTAIL.n34 VTAIL.n19 171.744
R114 VTAIL.n41 VTAIL.n19 171.744
R115 VTAIL.n42 VTAIL.n41 171.744
R116 VTAIL.n42 VTAIL.n15 171.744
R117 VTAIL.n49 VTAIL.n15 171.744
R118 VTAIL.n50 VTAIL.n49 171.744
R119 VTAIL.n50 VTAIL.n11 171.744
R120 VTAIL.n57 VTAIL.n11 171.744
R121 VTAIL.n58 VTAIL.n57 171.744
R122 VTAIL.n58 VTAIL.n7 171.744
R123 VTAIL.n65 VTAIL.n7 171.744
R124 VTAIL.n67 VTAIL.n65 171.744
R125 VTAIL.n67 VTAIL.n66 171.744
R126 VTAIL.n66 VTAIL.n3 171.744
R127 VTAIL.n75 VTAIL.n3 171.744
R128 VTAIL.n76 VTAIL.n75 171.744
R129 VTAIL.n240 VTAIL.n239 171.744
R130 VTAIL.n239 VTAIL.n167 171.744
R131 VTAIL.n171 VTAIL.n167 171.744
R132 VTAIL.n231 VTAIL.n171 171.744
R133 VTAIL.n231 VTAIL.n230 171.744
R134 VTAIL.n230 VTAIL.n172 171.744
R135 VTAIL.n223 VTAIL.n172 171.744
R136 VTAIL.n223 VTAIL.n222 171.744
R137 VTAIL.n222 VTAIL.n176 171.744
R138 VTAIL.n215 VTAIL.n176 171.744
R139 VTAIL.n215 VTAIL.n214 171.744
R140 VTAIL.n214 VTAIL.n180 171.744
R141 VTAIL.n207 VTAIL.n180 171.744
R142 VTAIL.n207 VTAIL.n206 171.744
R143 VTAIL.n206 VTAIL.n184 171.744
R144 VTAIL.n199 VTAIL.n184 171.744
R145 VTAIL.n199 VTAIL.n198 171.744
R146 VTAIL.n198 VTAIL.n188 171.744
R147 VTAIL.n191 VTAIL.n188 171.744
R148 VTAIL.n158 VTAIL.n157 171.744
R149 VTAIL.n157 VTAIL.n85 171.744
R150 VTAIL.n89 VTAIL.n85 171.744
R151 VTAIL.n149 VTAIL.n89 171.744
R152 VTAIL.n149 VTAIL.n148 171.744
R153 VTAIL.n148 VTAIL.n90 171.744
R154 VTAIL.n141 VTAIL.n90 171.744
R155 VTAIL.n141 VTAIL.n140 171.744
R156 VTAIL.n140 VTAIL.n94 171.744
R157 VTAIL.n133 VTAIL.n94 171.744
R158 VTAIL.n133 VTAIL.n132 171.744
R159 VTAIL.n132 VTAIL.n98 171.744
R160 VTAIL.n125 VTAIL.n98 171.744
R161 VTAIL.n125 VTAIL.n124 171.744
R162 VTAIL.n124 VTAIL.n102 171.744
R163 VTAIL.n117 VTAIL.n102 171.744
R164 VTAIL.n117 VTAIL.n116 171.744
R165 VTAIL.n116 VTAIL.n106 171.744
R166 VTAIL.n109 VTAIL.n106 171.744
R167 VTAIL.n272 VTAIL.t0 85.8723
R168 VTAIL.n26 VTAIL.t3 85.8723
R169 VTAIL.n191 VTAIL.t2 85.8723
R170 VTAIL.n109 VTAIL.t1 85.8723
R171 VTAIL.n327 VTAIL.n326 33.155
R172 VTAIL.n81 VTAIL.n80 33.155
R173 VTAIL.n245 VTAIL.n244 33.155
R174 VTAIL.n163 VTAIL.n162 33.155
R175 VTAIL.n163 VTAIL.n81 28.7203
R176 VTAIL.n327 VTAIL.n245 26.8755
R177 VTAIL.n273 VTAIL.n271 16.3895
R178 VTAIL.n27 VTAIL.n25 16.3895
R179 VTAIL.n192 VTAIL.n190 16.3895
R180 VTAIL.n110 VTAIL.n108 16.3895
R181 VTAIL.n320 VTAIL.n319 13.1884
R182 VTAIL.n74 VTAIL.n73 13.1884
R183 VTAIL.n238 VTAIL.n237 13.1884
R184 VTAIL.n156 VTAIL.n155 13.1884
R185 VTAIL.n274 VTAIL.n270 12.8005
R186 VTAIL.n318 VTAIL.n250 12.8005
R187 VTAIL.n323 VTAIL.n248 12.8005
R188 VTAIL.n28 VTAIL.n24 12.8005
R189 VTAIL.n72 VTAIL.n4 12.8005
R190 VTAIL.n77 VTAIL.n2 12.8005
R191 VTAIL.n241 VTAIL.n166 12.8005
R192 VTAIL.n236 VTAIL.n168 12.8005
R193 VTAIL.n193 VTAIL.n189 12.8005
R194 VTAIL.n159 VTAIL.n84 12.8005
R195 VTAIL.n154 VTAIL.n86 12.8005
R196 VTAIL.n111 VTAIL.n107 12.8005
R197 VTAIL.n278 VTAIL.n277 12.0247
R198 VTAIL.n315 VTAIL.n314 12.0247
R199 VTAIL.n324 VTAIL.n246 12.0247
R200 VTAIL.n32 VTAIL.n31 12.0247
R201 VTAIL.n69 VTAIL.n68 12.0247
R202 VTAIL.n78 VTAIL.n0 12.0247
R203 VTAIL.n242 VTAIL.n164 12.0247
R204 VTAIL.n233 VTAIL.n232 12.0247
R205 VTAIL.n197 VTAIL.n196 12.0247
R206 VTAIL.n160 VTAIL.n82 12.0247
R207 VTAIL.n151 VTAIL.n150 12.0247
R208 VTAIL.n115 VTAIL.n114 12.0247
R209 VTAIL.n281 VTAIL.n268 11.249
R210 VTAIL.n310 VTAIL.n252 11.249
R211 VTAIL.n35 VTAIL.n22 11.249
R212 VTAIL.n64 VTAIL.n6 11.249
R213 VTAIL.n229 VTAIL.n170 11.249
R214 VTAIL.n200 VTAIL.n187 11.249
R215 VTAIL.n147 VTAIL.n88 11.249
R216 VTAIL.n118 VTAIL.n105 11.249
R217 VTAIL.n282 VTAIL.n266 10.4732
R218 VTAIL.n309 VTAIL.n254 10.4732
R219 VTAIL.n36 VTAIL.n20 10.4732
R220 VTAIL.n63 VTAIL.n8 10.4732
R221 VTAIL.n228 VTAIL.n173 10.4732
R222 VTAIL.n201 VTAIL.n185 10.4732
R223 VTAIL.n146 VTAIL.n91 10.4732
R224 VTAIL.n119 VTAIL.n103 10.4732
R225 VTAIL.n286 VTAIL.n285 9.69747
R226 VTAIL.n306 VTAIL.n305 9.69747
R227 VTAIL.n40 VTAIL.n39 9.69747
R228 VTAIL.n60 VTAIL.n59 9.69747
R229 VTAIL.n225 VTAIL.n224 9.69747
R230 VTAIL.n205 VTAIL.n204 9.69747
R231 VTAIL.n143 VTAIL.n142 9.69747
R232 VTAIL.n123 VTAIL.n122 9.69747
R233 VTAIL.n326 VTAIL.n325 9.45567
R234 VTAIL.n80 VTAIL.n79 9.45567
R235 VTAIL.n244 VTAIL.n243 9.45567
R236 VTAIL.n162 VTAIL.n161 9.45567
R237 VTAIL.n325 VTAIL.n324 9.3005
R238 VTAIL.n248 VTAIL.n247 9.3005
R239 VTAIL.n293 VTAIL.n292 9.3005
R240 VTAIL.n291 VTAIL.n290 9.3005
R241 VTAIL.n264 VTAIL.n263 9.3005
R242 VTAIL.n285 VTAIL.n284 9.3005
R243 VTAIL.n283 VTAIL.n282 9.3005
R244 VTAIL.n268 VTAIL.n267 9.3005
R245 VTAIL.n277 VTAIL.n276 9.3005
R246 VTAIL.n275 VTAIL.n274 9.3005
R247 VTAIL.n260 VTAIL.n259 9.3005
R248 VTAIL.n299 VTAIL.n298 9.3005
R249 VTAIL.n301 VTAIL.n300 9.3005
R250 VTAIL.n256 VTAIL.n255 9.3005
R251 VTAIL.n307 VTAIL.n306 9.3005
R252 VTAIL.n309 VTAIL.n308 9.3005
R253 VTAIL.n252 VTAIL.n251 9.3005
R254 VTAIL.n316 VTAIL.n315 9.3005
R255 VTAIL.n318 VTAIL.n317 9.3005
R256 VTAIL.n79 VTAIL.n78 9.3005
R257 VTAIL.n2 VTAIL.n1 9.3005
R258 VTAIL.n47 VTAIL.n46 9.3005
R259 VTAIL.n45 VTAIL.n44 9.3005
R260 VTAIL.n18 VTAIL.n17 9.3005
R261 VTAIL.n39 VTAIL.n38 9.3005
R262 VTAIL.n37 VTAIL.n36 9.3005
R263 VTAIL.n22 VTAIL.n21 9.3005
R264 VTAIL.n31 VTAIL.n30 9.3005
R265 VTAIL.n29 VTAIL.n28 9.3005
R266 VTAIL.n14 VTAIL.n13 9.3005
R267 VTAIL.n53 VTAIL.n52 9.3005
R268 VTAIL.n55 VTAIL.n54 9.3005
R269 VTAIL.n10 VTAIL.n9 9.3005
R270 VTAIL.n61 VTAIL.n60 9.3005
R271 VTAIL.n63 VTAIL.n62 9.3005
R272 VTAIL.n6 VTAIL.n5 9.3005
R273 VTAIL.n70 VTAIL.n69 9.3005
R274 VTAIL.n72 VTAIL.n71 9.3005
R275 VTAIL.n218 VTAIL.n217 9.3005
R276 VTAIL.n220 VTAIL.n219 9.3005
R277 VTAIL.n175 VTAIL.n174 9.3005
R278 VTAIL.n226 VTAIL.n225 9.3005
R279 VTAIL.n228 VTAIL.n227 9.3005
R280 VTAIL.n170 VTAIL.n169 9.3005
R281 VTAIL.n234 VTAIL.n233 9.3005
R282 VTAIL.n236 VTAIL.n235 9.3005
R283 VTAIL.n243 VTAIL.n242 9.3005
R284 VTAIL.n166 VTAIL.n165 9.3005
R285 VTAIL.n179 VTAIL.n178 9.3005
R286 VTAIL.n212 VTAIL.n211 9.3005
R287 VTAIL.n210 VTAIL.n209 9.3005
R288 VTAIL.n183 VTAIL.n182 9.3005
R289 VTAIL.n204 VTAIL.n203 9.3005
R290 VTAIL.n202 VTAIL.n201 9.3005
R291 VTAIL.n187 VTAIL.n186 9.3005
R292 VTAIL.n196 VTAIL.n195 9.3005
R293 VTAIL.n194 VTAIL.n193 9.3005
R294 VTAIL.n136 VTAIL.n135 9.3005
R295 VTAIL.n138 VTAIL.n137 9.3005
R296 VTAIL.n93 VTAIL.n92 9.3005
R297 VTAIL.n144 VTAIL.n143 9.3005
R298 VTAIL.n146 VTAIL.n145 9.3005
R299 VTAIL.n88 VTAIL.n87 9.3005
R300 VTAIL.n152 VTAIL.n151 9.3005
R301 VTAIL.n154 VTAIL.n153 9.3005
R302 VTAIL.n161 VTAIL.n160 9.3005
R303 VTAIL.n84 VTAIL.n83 9.3005
R304 VTAIL.n97 VTAIL.n96 9.3005
R305 VTAIL.n130 VTAIL.n129 9.3005
R306 VTAIL.n128 VTAIL.n127 9.3005
R307 VTAIL.n101 VTAIL.n100 9.3005
R308 VTAIL.n122 VTAIL.n121 9.3005
R309 VTAIL.n120 VTAIL.n119 9.3005
R310 VTAIL.n105 VTAIL.n104 9.3005
R311 VTAIL.n114 VTAIL.n113 9.3005
R312 VTAIL.n112 VTAIL.n111 9.3005
R313 VTAIL.n289 VTAIL.n264 8.92171
R314 VTAIL.n302 VTAIL.n256 8.92171
R315 VTAIL.n43 VTAIL.n18 8.92171
R316 VTAIL.n56 VTAIL.n10 8.92171
R317 VTAIL.n221 VTAIL.n175 8.92171
R318 VTAIL.n208 VTAIL.n183 8.92171
R319 VTAIL.n139 VTAIL.n93 8.92171
R320 VTAIL.n126 VTAIL.n101 8.92171
R321 VTAIL.n290 VTAIL.n262 8.14595
R322 VTAIL.n301 VTAIL.n258 8.14595
R323 VTAIL.n44 VTAIL.n16 8.14595
R324 VTAIL.n55 VTAIL.n12 8.14595
R325 VTAIL.n220 VTAIL.n177 8.14595
R326 VTAIL.n209 VTAIL.n181 8.14595
R327 VTAIL.n138 VTAIL.n95 8.14595
R328 VTAIL.n127 VTAIL.n99 8.14595
R329 VTAIL.n294 VTAIL.n293 7.3702
R330 VTAIL.n298 VTAIL.n297 7.3702
R331 VTAIL.n48 VTAIL.n47 7.3702
R332 VTAIL.n52 VTAIL.n51 7.3702
R333 VTAIL.n217 VTAIL.n216 7.3702
R334 VTAIL.n213 VTAIL.n212 7.3702
R335 VTAIL.n135 VTAIL.n134 7.3702
R336 VTAIL.n131 VTAIL.n130 7.3702
R337 VTAIL.n294 VTAIL.n260 6.59444
R338 VTAIL.n297 VTAIL.n260 6.59444
R339 VTAIL.n48 VTAIL.n14 6.59444
R340 VTAIL.n51 VTAIL.n14 6.59444
R341 VTAIL.n216 VTAIL.n179 6.59444
R342 VTAIL.n213 VTAIL.n179 6.59444
R343 VTAIL.n134 VTAIL.n97 6.59444
R344 VTAIL.n131 VTAIL.n97 6.59444
R345 VTAIL.n293 VTAIL.n262 5.81868
R346 VTAIL.n298 VTAIL.n258 5.81868
R347 VTAIL.n47 VTAIL.n16 5.81868
R348 VTAIL.n52 VTAIL.n12 5.81868
R349 VTAIL.n217 VTAIL.n177 5.81868
R350 VTAIL.n212 VTAIL.n181 5.81868
R351 VTAIL.n135 VTAIL.n95 5.81868
R352 VTAIL.n130 VTAIL.n99 5.81868
R353 VTAIL.n290 VTAIL.n289 5.04292
R354 VTAIL.n302 VTAIL.n301 5.04292
R355 VTAIL.n44 VTAIL.n43 5.04292
R356 VTAIL.n56 VTAIL.n55 5.04292
R357 VTAIL.n221 VTAIL.n220 5.04292
R358 VTAIL.n209 VTAIL.n208 5.04292
R359 VTAIL.n139 VTAIL.n138 5.04292
R360 VTAIL.n127 VTAIL.n126 5.04292
R361 VTAIL.n286 VTAIL.n264 4.26717
R362 VTAIL.n305 VTAIL.n256 4.26717
R363 VTAIL.n40 VTAIL.n18 4.26717
R364 VTAIL.n59 VTAIL.n10 4.26717
R365 VTAIL.n224 VTAIL.n175 4.26717
R366 VTAIL.n205 VTAIL.n183 4.26717
R367 VTAIL.n142 VTAIL.n93 4.26717
R368 VTAIL.n123 VTAIL.n101 4.26717
R369 VTAIL.n275 VTAIL.n271 3.70982
R370 VTAIL.n29 VTAIL.n25 3.70982
R371 VTAIL.n194 VTAIL.n190 3.70982
R372 VTAIL.n112 VTAIL.n108 3.70982
R373 VTAIL.n285 VTAIL.n266 3.49141
R374 VTAIL.n306 VTAIL.n254 3.49141
R375 VTAIL.n39 VTAIL.n20 3.49141
R376 VTAIL.n60 VTAIL.n8 3.49141
R377 VTAIL.n225 VTAIL.n173 3.49141
R378 VTAIL.n204 VTAIL.n185 3.49141
R379 VTAIL.n143 VTAIL.n91 3.49141
R380 VTAIL.n122 VTAIL.n103 3.49141
R381 VTAIL.n282 VTAIL.n281 2.71565
R382 VTAIL.n310 VTAIL.n309 2.71565
R383 VTAIL.n36 VTAIL.n35 2.71565
R384 VTAIL.n64 VTAIL.n63 2.71565
R385 VTAIL.n229 VTAIL.n228 2.71565
R386 VTAIL.n201 VTAIL.n200 2.71565
R387 VTAIL.n147 VTAIL.n146 2.71565
R388 VTAIL.n119 VTAIL.n118 2.71565
R389 VTAIL.n278 VTAIL.n268 1.93989
R390 VTAIL.n314 VTAIL.n252 1.93989
R391 VTAIL.n326 VTAIL.n246 1.93989
R392 VTAIL.n32 VTAIL.n22 1.93989
R393 VTAIL.n68 VTAIL.n6 1.93989
R394 VTAIL.n80 VTAIL.n0 1.93989
R395 VTAIL.n244 VTAIL.n164 1.93989
R396 VTAIL.n232 VTAIL.n170 1.93989
R397 VTAIL.n197 VTAIL.n187 1.93989
R398 VTAIL.n162 VTAIL.n82 1.93989
R399 VTAIL.n150 VTAIL.n88 1.93989
R400 VTAIL.n115 VTAIL.n105 1.93989
R401 VTAIL.n245 VTAIL.n163 1.39274
R402 VTAIL.n277 VTAIL.n270 1.16414
R403 VTAIL.n315 VTAIL.n250 1.16414
R404 VTAIL.n324 VTAIL.n323 1.16414
R405 VTAIL.n31 VTAIL.n24 1.16414
R406 VTAIL.n69 VTAIL.n4 1.16414
R407 VTAIL.n78 VTAIL.n77 1.16414
R408 VTAIL.n242 VTAIL.n241 1.16414
R409 VTAIL.n233 VTAIL.n168 1.16414
R410 VTAIL.n196 VTAIL.n189 1.16414
R411 VTAIL.n160 VTAIL.n159 1.16414
R412 VTAIL.n151 VTAIL.n86 1.16414
R413 VTAIL.n114 VTAIL.n107 1.16414
R414 VTAIL VTAIL.n81 0.989724
R415 VTAIL VTAIL.n327 0.403517
R416 VTAIL.n274 VTAIL.n273 0.388379
R417 VTAIL.n319 VTAIL.n318 0.388379
R418 VTAIL.n320 VTAIL.n248 0.388379
R419 VTAIL.n28 VTAIL.n27 0.388379
R420 VTAIL.n73 VTAIL.n72 0.388379
R421 VTAIL.n74 VTAIL.n2 0.388379
R422 VTAIL.n238 VTAIL.n166 0.388379
R423 VTAIL.n237 VTAIL.n236 0.388379
R424 VTAIL.n193 VTAIL.n192 0.388379
R425 VTAIL.n156 VTAIL.n84 0.388379
R426 VTAIL.n155 VTAIL.n154 0.388379
R427 VTAIL.n111 VTAIL.n110 0.388379
R428 VTAIL.n276 VTAIL.n275 0.155672
R429 VTAIL.n276 VTAIL.n267 0.155672
R430 VTAIL.n283 VTAIL.n267 0.155672
R431 VTAIL.n284 VTAIL.n283 0.155672
R432 VTAIL.n284 VTAIL.n263 0.155672
R433 VTAIL.n291 VTAIL.n263 0.155672
R434 VTAIL.n292 VTAIL.n291 0.155672
R435 VTAIL.n292 VTAIL.n259 0.155672
R436 VTAIL.n299 VTAIL.n259 0.155672
R437 VTAIL.n300 VTAIL.n299 0.155672
R438 VTAIL.n300 VTAIL.n255 0.155672
R439 VTAIL.n307 VTAIL.n255 0.155672
R440 VTAIL.n308 VTAIL.n307 0.155672
R441 VTAIL.n308 VTAIL.n251 0.155672
R442 VTAIL.n316 VTAIL.n251 0.155672
R443 VTAIL.n317 VTAIL.n316 0.155672
R444 VTAIL.n317 VTAIL.n247 0.155672
R445 VTAIL.n325 VTAIL.n247 0.155672
R446 VTAIL.n30 VTAIL.n29 0.155672
R447 VTAIL.n30 VTAIL.n21 0.155672
R448 VTAIL.n37 VTAIL.n21 0.155672
R449 VTAIL.n38 VTAIL.n37 0.155672
R450 VTAIL.n38 VTAIL.n17 0.155672
R451 VTAIL.n45 VTAIL.n17 0.155672
R452 VTAIL.n46 VTAIL.n45 0.155672
R453 VTAIL.n46 VTAIL.n13 0.155672
R454 VTAIL.n53 VTAIL.n13 0.155672
R455 VTAIL.n54 VTAIL.n53 0.155672
R456 VTAIL.n54 VTAIL.n9 0.155672
R457 VTAIL.n61 VTAIL.n9 0.155672
R458 VTAIL.n62 VTAIL.n61 0.155672
R459 VTAIL.n62 VTAIL.n5 0.155672
R460 VTAIL.n70 VTAIL.n5 0.155672
R461 VTAIL.n71 VTAIL.n70 0.155672
R462 VTAIL.n71 VTAIL.n1 0.155672
R463 VTAIL.n79 VTAIL.n1 0.155672
R464 VTAIL.n243 VTAIL.n165 0.155672
R465 VTAIL.n235 VTAIL.n165 0.155672
R466 VTAIL.n235 VTAIL.n234 0.155672
R467 VTAIL.n234 VTAIL.n169 0.155672
R468 VTAIL.n227 VTAIL.n169 0.155672
R469 VTAIL.n227 VTAIL.n226 0.155672
R470 VTAIL.n226 VTAIL.n174 0.155672
R471 VTAIL.n219 VTAIL.n174 0.155672
R472 VTAIL.n219 VTAIL.n218 0.155672
R473 VTAIL.n218 VTAIL.n178 0.155672
R474 VTAIL.n211 VTAIL.n178 0.155672
R475 VTAIL.n211 VTAIL.n210 0.155672
R476 VTAIL.n210 VTAIL.n182 0.155672
R477 VTAIL.n203 VTAIL.n182 0.155672
R478 VTAIL.n203 VTAIL.n202 0.155672
R479 VTAIL.n202 VTAIL.n186 0.155672
R480 VTAIL.n195 VTAIL.n186 0.155672
R481 VTAIL.n195 VTAIL.n194 0.155672
R482 VTAIL.n161 VTAIL.n83 0.155672
R483 VTAIL.n153 VTAIL.n83 0.155672
R484 VTAIL.n153 VTAIL.n152 0.155672
R485 VTAIL.n152 VTAIL.n87 0.155672
R486 VTAIL.n145 VTAIL.n87 0.155672
R487 VTAIL.n145 VTAIL.n144 0.155672
R488 VTAIL.n144 VTAIL.n92 0.155672
R489 VTAIL.n137 VTAIL.n92 0.155672
R490 VTAIL.n137 VTAIL.n136 0.155672
R491 VTAIL.n136 VTAIL.n96 0.155672
R492 VTAIL.n129 VTAIL.n96 0.155672
R493 VTAIL.n129 VTAIL.n128 0.155672
R494 VTAIL.n128 VTAIL.n100 0.155672
R495 VTAIL.n121 VTAIL.n100 0.155672
R496 VTAIL.n121 VTAIL.n120 0.155672
R497 VTAIL.n120 VTAIL.n104 0.155672
R498 VTAIL.n113 VTAIL.n104 0.155672
R499 VTAIL.n113 VTAIL.n112 0.155672
R500 VDD1.n76 VDD1.n0 756.745
R501 VDD1.n157 VDD1.n81 756.745
R502 VDD1.n77 VDD1.n76 585
R503 VDD1.n75 VDD1.n74 585
R504 VDD1.n73 VDD1.n3 585
R505 VDD1.n7 VDD1.n4 585
R506 VDD1.n68 VDD1.n67 585
R507 VDD1.n66 VDD1.n65 585
R508 VDD1.n9 VDD1.n8 585
R509 VDD1.n60 VDD1.n59 585
R510 VDD1.n58 VDD1.n57 585
R511 VDD1.n13 VDD1.n12 585
R512 VDD1.n52 VDD1.n51 585
R513 VDD1.n50 VDD1.n49 585
R514 VDD1.n17 VDD1.n16 585
R515 VDD1.n44 VDD1.n43 585
R516 VDD1.n42 VDD1.n41 585
R517 VDD1.n21 VDD1.n20 585
R518 VDD1.n36 VDD1.n35 585
R519 VDD1.n34 VDD1.n33 585
R520 VDD1.n25 VDD1.n24 585
R521 VDD1.n28 VDD1.n27 585
R522 VDD1.n108 VDD1.n107 585
R523 VDD1.n105 VDD1.n104 585
R524 VDD1.n114 VDD1.n113 585
R525 VDD1.n116 VDD1.n115 585
R526 VDD1.n101 VDD1.n100 585
R527 VDD1.n122 VDD1.n121 585
R528 VDD1.n124 VDD1.n123 585
R529 VDD1.n97 VDD1.n96 585
R530 VDD1.n130 VDD1.n129 585
R531 VDD1.n132 VDD1.n131 585
R532 VDD1.n93 VDD1.n92 585
R533 VDD1.n138 VDD1.n137 585
R534 VDD1.n140 VDD1.n139 585
R535 VDD1.n89 VDD1.n88 585
R536 VDD1.n146 VDD1.n145 585
R537 VDD1.n149 VDD1.n148 585
R538 VDD1.n147 VDD1.n85 585
R539 VDD1.n154 VDD1.n84 585
R540 VDD1.n156 VDD1.n155 585
R541 VDD1.n158 VDD1.n157 585
R542 VDD1.t0 VDD1.n26 327.466
R543 VDD1.t1 VDD1.n106 327.466
R544 VDD1.n76 VDD1.n75 171.744
R545 VDD1.n75 VDD1.n3 171.744
R546 VDD1.n7 VDD1.n3 171.744
R547 VDD1.n67 VDD1.n7 171.744
R548 VDD1.n67 VDD1.n66 171.744
R549 VDD1.n66 VDD1.n8 171.744
R550 VDD1.n59 VDD1.n8 171.744
R551 VDD1.n59 VDD1.n58 171.744
R552 VDD1.n58 VDD1.n12 171.744
R553 VDD1.n51 VDD1.n12 171.744
R554 VDD1.n51 VDD1.n50 171.744
R555 VDD1.n50 VDD1.n16 171.744
R556 VDD1.n43 VDD1.n16 171.744
R557 VDD1.n43 VDD1.n42 171.744
R558 VDD1.n42 VDD1.n20 171.744
R559 VDD1.n35 VDD1.n20 171.744
R560 VDD1.n35 VDD1.n34 171.744
R561 VDD1.n34 VDD1.n24 171.744
R562 VDD1.n27 VDD1.n24 171.744
R563 VDD1.n107 VDD1.n104 171.744
R564 VDD1.n114 VDD1.n104 171.744
R565 VDD1.n115 VDD1.n114 171.744
R566 VDD1.n115 VDD1.n100 171.744
R567 VDD1.n122 VDD1.n100 171.744
R568 VDD1.n123 VDD1.n122 171.744
R569 VDD1.n123 VDD1.n96 171.744
R570 VDD1.n130 VDD1.n96 171.744
R571 VDD1.n131 VDD1.n130 171.744
R572 VDD1.n131 VDD1.n92 171.744
R573 VDD1.n138 VDD1.n92 171.744
R574 VDD1.n139 VDD1.n138 171.744
R575 VDD1.n139 VDD1.n88 171.744
R576 VDD1.n146 VDD1.n88 171.744
R577 VDD1.n148 VDD1.n146 171.744
R578 VDD1.n148 VDD1.n147 171.744
R579 VDD1.n147 VDD1.n84 171.744
R580 VDD1.n156 VDD1.n84 171.744
R581 VDD1.n157 VDD1.n156 171.744
R582 VDD1 VDD1.n161 90.8328
R583 VDD1.n27 VDD1.t0 85.8723
R584 VDD1.n107 VDD1.t1 85.8723
R585 VDD1 VDD1.n80 50.3532
R586 VDD1.n28 VDD1.n26 16.3895
R587 VDD1.n108 VDD1.n106 16.3895
R588 VDD1.n74 VDD1.n73 13.1884
R589 VDD1.n155 VDD1.n154 13.1884
R590 VDD1.n77 VDD1.n2 12.8005
R591 VDD1.n72 VDD1.n4 12.8005
R592 VDD1.n29 VDD1.n25 12.8005
R593 VDD1.n109 VDD1.n105 12.8005
R594 VDD1.n153 VDD1.n85 12.8005
R595 VDD1.n158 VDD1.n83 12.8005
R596 VDD1.n78 VDD1.n0 12.0247
R597 VDD1.n69 VDD1.n68 12.0247
R598 VDD1.n33 VDD1.n32 12.0247
R599 VDD1.n113 VDD1.n112 12.0247
R600 VDD1.n150 VDD1.n149 12.0247
R601 VDD1.n159 VDD1.n81 12.0247
R602 VDD1.n65 VDD1.n6 11.249
R603 VDD1.n36 VDD1.n23 11.249
R604 VDD1.n116 VDD1.n103 11.249
R605 VDD1.n145 VDD1.n87 11.249
R606 VDD1.n64 VDD1.n9 10.4732
R607 VDD1.n37 VDD1.n21 10.4732
R608 VDD1.n117 VDD1.n101 10.4732
R609 VDD1.n144 VDD1.n89 10.4732
R610 VDD1.n61 VDD1.n60 9.69747
R611 VDD1.n41 VDD1.n40 9.69747
R612 VDD1.n121 VDD1.n120 9.69747
R613 VDD1.n141 VDD1.n140 9.69747
R614 VDD1.n80 VDD1.n79 9.45567
R615 VDD1.n161 VDD1.n160 9.45567
R616 VDD1.n54 VDD1.n53 9.3005
R617 VDD1.n56 VDD1.n55 9.3005
R618 VDD1.n11 VDD1.n10 9.3005
R619 VDD1.n62 VDD1.n61 9.3005
R620 VDD1.n64 VDD1.n63 9.3005
R621 VDD1.n6 VDD1.n5 9.3005
R622 VDD1.n70 VDD1.n69 9.3005
R623 VDD1.n72 VDD1.n71 9.3005
R624 VDD1.n79 VDD1.n78 9.3005
R625 VDD1.n2 VDD1.n1 9.3005
R626 VDD1.n15 VDD1.n14 9.3005
R627 VDD1.n48 VDD1.n47 9.3005
R628 VDD1.n46 VDD1.n45 9.3005
R629 VDD1.n19 VDD1.n18 9.3005
R630 VDD1.n40 VDD1.n39 9.3005
R631 VDD1.n38 VDD1.n37 9.3005
R632 VDD1.n23 VDD1.n22 9.3005
R633 VDD1.n32 VDD1.n31 9.3005
R634 VDD1.n30 VDD1.n29 9.3005
R635 VDD1.n160 VDD1.n159 9.3005
R636 VDD1.n83 VDD1.n82 9.3005
R637 VDD1.n128 VDD1.n127 9.3005
R638 VDD1.n126 VDD1.n125 9.3005
R639 VDD1.n99 VDD1.n98 9.3005
R640 VDD1.n120 VDD1.n119 9.3005
R641 VDD1.n118 VDD1.n117 9.3005
R642 VDD1.n103 VDD1.n102 9.3005
R643 VDD1.n112 VDD1.n111 9.3005
R644 VDD1.n110 VDD1.n109 9.3005
R645 VDD1.n95 VDD1.n94 9.3005
R646 VDD1.n134 VDD1.n133 9.3005
R647 VDD1.n136 VDD1.n135 9.3005
R648 VDD1.n91 VDD1.n90 9.3005
R649 VDD1.n142 VDD1.n141 9.3005
R650 VDD1.n144 VDD1.n143 9.3005
R651 VDD1.n87 VDD1.n86 9.3005
R652 VDD1.n151 VDD1.n150 9.3005
R653 VDD1.n153 VDD1.n152 9.3005
R654 VDD1.n57 VDD1.n11 8.92171
R655 VDD1.n44 VDD1.n19 8.92171
R656 VDD1.n124 VDD1.n99 8.92171
R657 VDD1.n137 VDD1.n91 8.92171
R658 VDD1.n56 VDD1.n13 8.14595
R659 VDD1.n45 VDD1.n17 8.14595
R660 VDD1.n125 VDD1.n97 8.14595
R661 VDD1.n136 VDD1.n93 8.14595
R662 VDD1.n53 VDD1.n52 7.3702
R663 VDD1.n49 VDD1.n48 7.3702
R664 VDD1.n129 VDD1.n128 7.3702
R665 VDD1.n133 VDD1.n132 7.3702
R666 VDD1.n52 VDD1.n15 6.59444
R667 VDD1.n49 VDD1.n15 6.59444
R668 VDD1.n129 VDD1.n95 6.59444
R669 VDD1.n132 VDD1.n95 6.59444
R670 VDD1.n53 VDD1.n13 5.81868
R671 VDD1.n48 VDD1.n17 5.81868
R672 VDD1.n128 VDD1.n97 5.81868
R673 VDD1.n133 VDD1.n93 5.81868
R674 VDD1.n57 VDD1.n56 5.04292
R675 VDD1.n45 VDD1.n44 5.04292
R676 VDD1.n125 VDD1.n124 5.04292
R677 VDD1.n137 VDD1.n136 5.04292
R678 VDD1.n60 VDD1.n11 4.26717
R679 VDD1.n41 VDD1.n19 4.26717
R680 VDD1.n121 VDD1.n99 4.26717
R681 VDD1.n140 VDD1.n91 4.26717
R682 VDD1.n30 VDD1.n26 3.70982
R683 VDD1.n110 VDD1.n106 3.70982
R684 VDD1.n61 VDD1.n9 3.49141
R685 VDD1.n40 VDD1.n21 3.49141
R686 VDD1.n120 VDD1.n101 3.49141
R687 VDD1.n141 VDD1.n89 3.49141
R688 VDD1.n65 VDD1.n64 2.71565
R689 VDD1.n37 VDD1.n36 2.71565
R690 VDD1.n117 VDD1.n116 2.71565
R691 VDD1.n145 VDD1.n144 2.71565
R692 VDD1.n80 VDD1.n0 1.93989
R693 VDD1.n68 VDD1.n6 1.93989
R694 VDD1.n33 VDD1.n23 1.93989
R695 VDD1.n113 VDD1.n103 1.93989
R696 VDD1.n149 VDD1.n87 1.93989
R697 VDD1.n161 VDD1.n81 1.93989
R698 VDD1.n78 VDD1.n77 1.16414
R699 VDD1.n69 VDD1.n4 1.16414
R700 VDD1.n32 VDD1.n25 1.16414
R701 VDD1.n112 VDD1.n105 1.16414
R702 VDD1.n150 VDD1.n85 1.16414
R703 VDD1.n159 VDD1.n158 1.16414
R704 VDD1.n74 VDD1.n2 0.388379
R705 VDD1.n73 VDD1.n72 0.388379
R706 VDD1.n29 VDD1.n28 0.388379
R707 VDD1.n109 VDD1.n108 0.388379
R708 VDD1.n154 VDD1.n153 0.388379
R709 VDD1.n155 VDD1.n83 0.388379
R710 VDD1.n79 VDD1.n1 0.155672
R711 VDD1.n71 VDD1.n1 0.155672
R712 VDD1.n71 VDD1.n70 0.155672
R713 VDD1.n70 VDD1.n5 0.155672
R714 VDD1.n63 VDD1.n5 0.155672
R715 VDD1.n63 VDD1.n62 0.155672
R716 VDD1.n62 VDD1.n10 0.155672
R717 VDD1.n55 VDD1.n10 0.155672
R718 VDD1.n55 VDD1.n54 0.155672
R719 VDD1.n54 VDD1.n14 0.155672
R720 VDD1.n47 VDD1.n14 0.155672
R721 VDD1.n47 VDD1.n46 0.155672
R722 VDD1.n46 VDD1.n18 0.155672
R723 VDD1.n39 VDD1.n18 0.155672
R724 VDD1.n39 VDD1.n38 0.155672
R725 VDD1.n38 VDD1.n22 0.155672
R726 VDD1.n31 VDD1.n22 0.155672
R727 VDD1.n31 VDD1.n30 0.155672
R728 VDD1.n111 VDD1.n110 0.155672
R729 VDD1.n111 VDD1.n102 0.155672
R730 VDD1.n118 VDD1.n102 0.155672
R731 VDD1.n119 VDD1.n118 0.155672
R732 VDD1.n119 VDD1.n98 0.155672
R733 VDD1.n126 VDD1.n98 0.155672
R734 VDD1.n127 VDD1.n126 0.155672
R735 VDD1.n127 VDD1.n94 0.155672
R736 VDD1.n134 VDD1.n94 0.155672
R737 VDD1.n135 VDD1.n134 0.155672
R738 VDD1.n135 VDD1.n90 0.155672
R739 VDD1.n142 VDD1.n90 0.155672
R740 VDD1.n143 VDD1.n142 0.155672
R741 VDD1.n143 VDD1.n86 0.155672
R742 VDD1.n151 VDD1.n86 0.155672
R743 VDD1.n152 VDD1.n151 0.155672
R744 VDD1.n152 VDD1.n82 0.155672
R745 VDD1.n160 VDD1.n82 0.155672
R746 VN VN.t1 299.248
R747 VN VN.t0 254.698
R748 VDD2.n157 VDD2.n81 756.745
R749 VDD2.n76 VDD2.n0 756.745
R750 VDD2.n158 VDD2.n157 585
R751 VDD2.n156 VDD2.n155 585
R752 VDD2.n154 VDD2.n84 585
R753 VDD2.n88 VDD2.n85 585
R754 VDD2.n149 VDD2.n148 585
R755 VDD2.n147 VDD2.n146 585
R756 VDD2.n90 VDD2.n89 585
R757 VDD2.n141 VDD2.n140 585
R758 VDD2.n139 VDD2.n138 585
R759 VDD2.n94 VDD2.n93 585
R760 VDD2.n133 VDD2.n132 585
R761 VDD2.n131 VDD2.n130 585
R762 VDD2.n98 VDD2.n97 585
R763 VDD2.n125 VDD2.n124 585
R764 VDD2.n123 VDD2.n122 585
R765 VDD2.n102 VDD2.n101 585
R766 VDD2.n117 VDD2.n116 585
R767 VDD2.n115 VDD2.n114 585
R768 VDD2.n106 VDD2.n105 585
R769 VDD2.n109 VDD2.n108 585
R770 VDD2.n27 VDD2.n26 585
R771 VDD2.n24 VDD2.n23 585
R772 VDD2.n33 VDD2.n32 585
R773 VDD2.n35 VDD2.n34 585
R774 VDD2.n20 VDD2.n19 585
R775 VDD2.n41 VDD2.n40 585
R776 VDD2.n43 VDD2.n42 585
R777 VDD2.n16 VDD2.n15 585
R778 VDD2.n49 VDD2.n48 585
R779 VDD2.n51 VDD2.n50 585
R780 VDD2.n12 VDD2.n11 585
R781 VDD2.n57 VDD2.n56 585
R782 VDD2.n59 VDD2.n58 585
R783 VDD2.n8 VDD2.n7 585
R784 VDD2.n65 VDD2.n64 585
R785 VDD2.n68 VDD2.n67 585
R786 VDD2.n66 VDD2.n4 585
R787 VDD2.n73 VDD2.n3 585
R788 VDD2.n75 VDD2.n74 585
R789 VDD2.n77 VDD2.n76 585
R790 VDD2.t0 VDD2.n107 327.466
R791 VDD2.t1 VDD2.n25 327.466
R792 VDD2.n157 VDD2.n156 171.744
R793 VDD2.n156 VDD2.n84 171.744
R794 VDD2.n88 VDD2.n84 171.744
R795 VDD2.n148 VDD2.n88 171.744
R796 VDD2.n148 VDD2.n147 171.744
R797 VDD2.n147 VDD2.n89 171.744
R798 VDD2.n140 VDD2.n89 171.744
R799 VDD2.n140 VDD2.n139 171.744
R800 VDD2.n139 VDD2.n93 171.744
R801 VDD2.n132 VDD2.n93 171.744
R802 VDD2.n132 VDD2.n131 171.744
R803 VDD2.n131 VDD2.n97 171.744
R804 VDD2.n124 VDD2.n97 171.744
R805 VDD2.n124 VDD2.n123 171.744
R806 VDD2.n123 VDD2.n101 171.744
R807 VDD2.n116 VDD2.n101 171.744
R808 VDD2.n116 VDD2.n115 171.744
R809 VDD2.n115 VDD2.n105 171.744
R810 VDD2.n108 VDD2.n105 171.744
R811 VDD2.n26 VDD2.n23 171.744
R812 VDD2.n33 VDD2.n23 171.744
R813 VDD2.n34 VDD2.n33 171.744
R814 VDD2.n34 VDD2.n19 171.744
R815 VDD2.n41 VDD2.n19 171.744
R816 VDD2.n42 VDD2.n41 171.744
R817 VDD2.n42 VDD2.n15 171.744
R818 VDD2.n49 VDD2.n15 171.744
R819 VDD2.n50 VDD2.n49 171.744
R820 VDD2.n50 VDD2.n11 171.744
R821 VDD2.n57 VDD2.n11 171.744
R822 VDD2.n58 VDD2.n57 171.744
R823 VDD2.n58 VDD2.n7 171.744
R824 VDD2.n65 VDD2.n7 171.744
R825 VDD2.n67 VDD2.n65 171.744
R826 VDD2.n67 VDD2.n66 171.744
R827 VDD2.n66 VDD2.n3 171.744
R828 VDD2.n75 VDD2.n3 171.744
R829 VDD2.n76 VDD2.n75 171.744
R830 VDD2.n162 VDD2.n80 89.8467
R831 VDD2.n108 VDD2.t0 85.8723
R832 VDD2.n26 VDD2.t1 85.8723
R833 VDD2.n162 VDD2.n161 49.8338
R834 VDD2.n109 VDD2.n107 16.3895
R835 VDD2.n27 VDD2.n25 16.3895
R836 VDD2.n155 VDD2.n154 13.1884
R837 VDD2.n74 VDD2.n73 13.1884
R838 VDD2.n158 VDD2.n83 12.8005
R839 VDD2.n153 VDD2.n85 12.8005
R840 VDD2.n110 VDD2.n106 12.8005
R841 VDD2.n28 VDD2.n24 12.8005
R842 VDD2.n72 VDD2.n4 12.8005
R843 VDD2.n77 VDD2.n2 12.8005
R844 VDD2.n159 VDD2.n81 12.0247
R845 VDD2.n150 VDD2.n149 12.0247
R846 VDD2.n114 VDD2.n113 12.0247
R847 VDD2.n32 VDD2.n31 12.0247
R848 VDD2.n69 VDD2.n68 12.0247
R849 VDD2.n78 VDD2.n0 12.0247
R850 VDD2.n146 VDD2.n87 11.249
R851 VDD2.n117 VDD2.n104 11.249
R852 VDD2.n35 VDD2.n22 11.249
R853 VDD2.n64 VDD2.n6 11.249
R854 VDD2.n145 VDD2.n90 10.4732
R855 VDD2.n118 VDD2.n102 10.4732
R856 VDD2.n36 VDD2.n20 10.4732
R857 VDD2.n63 VDD2.n8 10.4732
R858 VDD2.n142 VDD2.n141 9.69747
R859 VDD2.n122 VDD2.n121 9.69747
R860 VDD2.n40 VDD2.n39 9.69747
R861 VDD2.n60 VDD2.n59 9.69747
R862 VDD2.n161 VDD2.n160 9.45567
R863 VDD2.n80 VDD2.n79 9.45567
R864 VDD2.n135 VDD2.n134 9.3005
R865 VDD2.n137 VDD2.n136 9.3005
R866 VDD2.n92 VDD2.n91 9.3005
R867 VDD2.n143 VDD2.n142 9.3005
R868 VDD2.n145 VDD2.n144 9.3005
R869 VDD2.n87 VDD2.n86 9.3005
R870 VDD2.n151 VDD2.n150 9.3005
R871 VDD2.n153 VDD2.n152 9.3005
R872 VDD2.n160 VDD2.n159 9.3005
R873 VDD2.n83 VDD2.n82 9.3005
R874 VDD2.n96 VDD2.n95 9.3005
R875 VDD2.n129 VDD2.n128 9.3005
R876 VDD2.n127 VDD2.n126 9.3005
R877 VDD2.n100 VDD2.n99 9.3005
R878 VDD2.n121 VDD2.n120 9.3005
R879 VDD2.n119 VDD2.n118 9.3005
R880 VDD2.n104 VDD2.n103 9.3005
R881 VDD2.n113 VDD2.n112 9.3005
R882 VDD2.n111 VDD2.n110 9.3005
R883 VDD2.n79 VDD2.n78 9.3005
R884 VDD2.n2 VDD2.n1 9.3005
R885 VDD2.n47 VDD2.n46 9.3005
R886 VDD2.n45 VDD2.n44 9.3005
R887 VDD2.n18 VDD2.n17 9.3005
R888 VDD2.n39 VDD2.n38 9.3005
R889 VDD2.n37 VDD2.n36 9.3005
R890 VDD2.n22 VDD2.n21 9.3005
R891 VDD2.n31 VDD2.n30 9.3005
R892 VDD2.n29 VDD2.n28 9.3005
R893 VDD2.n14 VDD2.n13 9.3005
R894 VDD2.n53 VDD2.n52 9.3005
R895 VDD2.n55 VDD2.n54 9.3005
R896 VDD2.n10 VDD2.n9 9.3005
R897 VDD2.n61 VDD2.n60 9.3005
R898 VDD2.n63 VDD2.n62 9.3005
R899 VDD2.n6 VDD2.n5 9.3005
R900 VDD2.n70 VDD2.n69 9.3005
R901 VDD2.n72 VDD2.n71 9.3005
R902 VDD2.n138 VDD2.n92 8.92171
R903 VDD2.n125 VDD2.n100 8.92171
R904 VDD2.n43 VDD2.n18 8.92171
R905 VDD2.n56 VDD2.n10 8.92171
R906 VDD2.n137 VDD2.n94 8.14595
R907 VDD2.n126 VDD2.n98 8.14595
R908 VDD2.n44 VDD2.n16 8.14595
R909 VDD2.n55 VDD2.n12 8.14595
R910 VDD2.n134 VDD2.n133 7.3702
R911 VDD2.n130 VDD2.n129 7.3702
R912 VDD2.n48 VDD2.n47 7.3702
R913 VDD2.n52 VDD2.n51 7.3702
R914 VDD2.n133 VDD2.n96 6.59444
R915 VDD2.n130 VDD2.n96 6.59444
R916 VDD2.n48 VDD2.n14 6.59444
R917 VDD2.n51 VDD2.n14 6.59444
R918 VDD2.n134 VDD2.n94 5.81868
R919 VDD2.n129 VDD2.n98 5.81868
R920 VDD2.n47 VDD2.n16 5.81868
R921 VDD2.n52 VDD2.n12 5.81868
R922 VDD2.n138 VDD2.n137 5.04292
R923 VDD2.n126 VDD2.n125 5.04292
R924 VDD2.n44 VDD2.n43 5.04292
R925 VDD2.n56 VDD2.n55 5.04292
R926 VDD2.n141 VDD2.n92 4.26717
R927 VDD2.n122 VDD2.n100 4.26717
R928 VDD2.n40 VDD2.n18 4.26717
R929 VDD2.n59 VDD2.n10 4.26717
R930 VDD2.n111 VDD2.n107 3.70982
R931 VDD2.n29 VDD2.n25 3.70982
R932 VDD2.n142 VDD2.n90 3.49141
R933 VDD2.n121 VDD2.n102 3.49141
R934 VDD2.n39 VDD2.n20 3.49141
R935 VDD2.n60 VDD2.n8 3.49141
R936 VDD2.n146 VDD2.n145 2.71565
R937 VDD2.n118 VDD2.n117 2.71565
R938 VDD2.n36 VDD2.n35 2.71565
R939 VDD2.n64 VDD2.n63 2.71565
R940 VDD2.n161 VDD2.n81 1.93989
R941 VDD2.n149 VDD2.n87 1.93989
R942 VDD2.n114 VDD2.n104 1.93989
R943 VDD2.n32 VDD2.n22 1.93989
R944 VDD2.n68 VDD2.n6 1.93989
R945 VDD2.n80 VDD2.n0 1.93989
R946 VDD2.n159 VDD2.n158 1.16414
R947 VDD2.n150 VDD2.n85 1.16414
R948 VDD2.n113 VDD2.n106 1.16414
R949 VDD2.n31 VDD2.n24 1.16414
R950 VDD2.n69 VDD2.n4 1.16414
R951 VDD2.n78 VDD2.n77 1.16414
R952 VDD2 VDD2.n162 0.519897
R953 VDD2.n155 VDD2.n83 0.388379
R954 VDD2.n154 VDD2.n153 0.388379
R955 VDD2.n110 VDD2.n109 0.388379
R956 VDD2.n28 VDD2.n27 0.388379
R957 VDD2.n73 VDD2.n72 0.388379
R958 VDD2.n74 VDD2.n2 0.388379
R959 VDD2.n160 VDD2.n82 0.155672
R960 VDD2.n152 VDD2.n82 0.155672
R961 VDD2.n152 VDD2.n151 0.155672
R962 VDD2.n151 VDD2.n86 0.155672
R963 VDD2.n144 VDD2.n86 0.155672
R964 VDD2.n144 VDD2.n143 0.155672
R965 VDD2.n143 VDD2.n91 0.155672
R966 VDD2.n136 VDD2.n91 0.155672
R967 VDD2.n136 VDD2.n135 0.155672
R968 VDD2.n135 VDD2.n95 0.155672
R969 VDD2.n128 VDD2.n95 0.155672
R970 VDD2.n128 VDD2.n127 0.155672
R971 VDD2.n127 VDD2.n99 0.155672
R972 VDD2.n120 VDD2.n99 0.155672
R973 VDD2.n120 VDD2.n119 0.155672
R974 VDD2.n119 VDD2.n103 0.155672
R975 VDD2.n112 VDD2.n103 0.155672
R976 VDD2.n112 VDD2.n111 0.155672
R977 VDD2.n30 VDD2.n29 0.155672
R978 VDD2.n30 VDD2.n21 0.155672
R979 VDD2.n37 VDD2.n21 0.155672
R980 VDD2.n38 VDD2.n37 0.155672
R981 VDD2.n38 VDD2.n17 0.155672
R982 VDD2.n45 VDD2.n17 0.155672
R983 VDD2.n46 VDD2.n45 0.155672
R984 VDD2.n46 VDD2.n13 0.155672
R985 VDD2.n53 VDD2.n13 0.155672
R986 VDD2.n54 VDD2.n53 0.155672
R987 VDD2.n54 VDD2.n9 0.155672
R988 VDD2.n61 VDD2.n9 0.155672
R989 VDD2.n62 VDD2.n61 0.155672
R990 VDD2.n62 VDD2.n5 0.155672
R991 VDD2.n70 VDD2.n5 0.155672
R992 VDD2.n71 VDD2.n70 0.155672
R993 VDD2.n71 VDD2.n1 0.155672
R994 VDD2.n79 VDD2.n1 0.155672
R995 B.n353 B.n352 585
R996 B.n351 B.n92 585
R997 B.n350 B.n349 585
R998 B.n348 B.n93 585
R999 B.n347 B.n346 585
R1000 B.n345 B.n94 585
R1001 B.n344 B.n343 585
R1002 B.n342 B.n95 585
R1003 B.n341 B.n340 585
R1004 B.n339 B.n96 585
R1005 B.n338 B.n337 585
R1006 B.n336 B.n97 585
R1007 B.n335 B.n334 585
R1008 B.n333 B.n98 585
R1009 B.n332 B.n331 585
R1010 B.n330 B.n99 585
R1011 B.n329 B.n328 585
R1012 B.n327 B.n100 585
R1013 B.n326 B.n325 585
R1014 B.n324 B.n101 585
R1015 B.n323 B.n322 585
R1016 B.n321 B.n102 585
R1017 B.n320 B.n319 585
R1018 B.n318 B.n103 585
R1019 B.n317 B.n316 585
R1020 B.n315 B.n104 585
R1021 B.n314 B.n313 585
R1022 B.n312 B.n105 585
R1023 B.n311 B.n310 585
R1024 B.n309 B.n106 585
R1025 B.n308 B.n307 585
R1026 B.n306 B.n107 585
R1027 B.n305 B.n304 585
R1028 B.n303 B.n108 585
R1029 B.n302 B.n301 585
R1030 B.n300 B.n109 585
R1031 B.n299 B.n298 585
R1032 B.n297 B.n110 585
R1033 B.n296 B.n295 585
R1034 B.n294 B.n111 585
R1035 B.n293 B.n292 585
R1036 B.n291 B.n112 585
R1037 B.n290 B.n289 585
R1038 B.n288 B.n113 585
R1039 B.n287 B.n286 585
R1040 B.n285 B.n114 585
R1041 B.n284 B.n283 585
R1042 B.n282 B.n115 585
R1043 B.n281 B.n280 585
R1044 B.n279 B.n116 585
R1045 B.n278 B.n277 585
R1046 B.n273 B.n117 585
R1047 B.n272 B.n271 585
R1048 B.n270 B.n118 585
R1049 B.n269 B.n268 585
R1050 B.n267 B.n119 585
R1051 B.n266 B.n265 585
R1052 B.n264 B.n120 585
R1053 B.n263 B.n262 585
R1054 B.n260 B.n121 585
R1055 B.n259 B.n258 585
R1056 B.n257 B.n124 585
R1057 B.n256 B.n255 585
R1058 B.n254 B.n125 585
R1059 B.n253 B.n252 585
R1060 B.n251 B.n126 585
R1061 B.n250 B.n249 585
R1062 B.n248 B.n127 585
R1063 B.n247 B.n246 585
R1064 B.n245 B.n128 585
R1065 B.n244 B.n243 585
R1066 B.n242 B.n129 585
R1067 B.n241 B.n240 585
R1068 B.n239 B.n130 585
R1069 B.n238 B.n237 585
R1070 B.n236 B.n131 585
R1071 B.n235 B.n234 585
R1072 B.n233 B.n132 585
R1073 B.n232 B.n231 585
R1074 B.n230 B.n133 585
R1075 B.n229 B.n228 585
R1076 B.n227 B.n134 585
R1077 B.n226 B.n225 585
R1078 B.n224 B.n135 585
R1079 B.n223 B.n222 585
R1080 B.n221 B.n136 585
R1081 B.n220 B.n219 585
R1082 B.n218 B.n137 585
R1083 B.n217 B.n216 585
R1084 B.n215 B.n138 585
R1085 B.n214 B.n213 585
R1086 B.n212 B.n139 585
R1087 B.n211 B.n210 585
R1088 B.n209 B.n140 585
R1089 B.n208 B.n207 585
R1090 B.n206 B.n141 585
R1091 B.n205 B.n204 585
R1092 B.n203 B.n142 585
R1093 B.n202 B.n201 585
R1094 B.n200 B.n143 585
R1095 B.n199 B.n198 585
R1096 B.n197 B.n144 585
R1097 B.n196 B.n195 585
R1098 B.n194 B.n145 585
R1099 B.n193 B.n192 585
R1100 B.n191 B.n146 585
R1101 B.n190 B.n189 585
R1102 B.n188 B.n147 585
R1103 B.n187 B.n186 585
R1104 B.n354 B.n91 585
R1105 B.n356 B.n355 585
R1106 B.n357 B.n90 585
R1107 B.n359 B.n358 585
R1108 B.n360 B.n89 585
R1109 B.n362 B.n361 585
R1110 B.n363 B.n88 585
R1111 B.n365 B.n364 585
R1112 B.n366 B.n87 585
R1113 B.n368 B.n367 585
R1114 B.n369 B.n86 585
R1115 B.n371 B.n370 585
R1116 B.n372 B.n85 585
R1117 B.n374 B.n373 585
R1118 B.n375 B.n84 585
R1119 B.n377 B.n376 585
R1120 B.n378 B.n83 585
R1121 B.n380 B.n379 585
R1122 B.n381 B.n82 585
R1123 B.n383 B.n382 585
R1124 B.n384 B.n81 585
R1125 B.n386 B.n385 585
R1126 B.n387 B.n80 585
R1127 B.n389 B.n388 585
R1128 B.n390 B.n79 585
R1129 B.n392 B.n391 585
R1130 B.n393 B.n78 585
R1131 B.n395 B.n394 585
R1132 B.n396 B.n77 585
R1133 B.n398 B.n397 585
R1134 B.n399 B.n76 585
R1135 B.n401 B.n400 585
R1136 B.n402 B.n75 585
R1137 B.n404 B.n403 585
R1138 B.n405 B.n74 585
R1139 B.n407 B.n406 585
R1140 B.n408 B.n73 585
R1141 B.n410 B.n409 585
R1142 B.n411 B.n72 585
R1143 B.n413 B.n412 585
R1144 B.n414 B.n71 585
R1145 B.n416 B.n415 585
R1146 B.n581 B.n12 585
R1147 B.n580 B.n579 585
R1148 B.n578 B.n13 585
R1149 B.n577 B.n576 585
R1150 B.n575 B.n14 585
R1151 B.n574 B.n573 585
R1152 B.n572 B.n15 585
R1153 B.n571 B.n570 585
R1154 B.n569 B.n16 585
R1155 B.n568 B.n567 585
R1156 B.n566 B.n17 585
R1157 B.n565 B.n564 585
R1158 B.n563 B.n18 585
R1159 B.n562 B.n561 585
R1160 B.n560 B.n19 585
R1161 B.n559 B.n558 585
R1162 B.n557 B.n20 585
R1163 B.n556 B.n555 585
R1164 B.n554 B.n21 585
R1165 B.n553 B.n552 585
R1166 B.n551 B.n22 585
R1167 B.n550 B.n549 585
R1168 B.n548 B.n23 585
R1169 B.n547 B.n546 585
R1170 B.n545 B.n24 585
R1171 B.n544 B.n543 585
R1172 B.n542 B.n25 585
R1173 B.n541 B.n540 585
R1174 B.n539 B.n26 585
R1175 B.n538 B.n537 585
R1176 B.n536 B.n27 585
R1177 B.n535 B.n534 585
R1178 B.n533 B.n28 585
R1179 B.n532 B.n531 585
R1180 B.n530 B.n29 585
R1181 B.n529 B.n528 585
R1182 B.n527 B.n30 585
R1183 B.n526 B.n525 585
R1184 B.n524 B.n31 585
R1185 B.n523 B.n522 585
R1186 B.n521 B.n32 585
R1187 B.n520 B.n519 585
R1188 B.n518 B.n33 585
R1189 B.n517 B.n516 585
R1190 B.n515 B.n34 585
R1191 B.n514 B.n513 585
R1192 B.n512 B.n35 585
R1193 B.n511 B.n510 585
R1194 B.n509 B.n36 585
R1195 B.n508 B.n507 585
R1196 B.n505 B.n37 585
R1197 B.n504 B.n503 585
R1198 B.n502 B.n40 585
R1199 B.n501 B.n500 585
R1200 B.n499 B.n41 585
R1201 B.n498 B.n497 585
R1202 B.n496 B.n42 585
R1203 B.n495 B.n494 585
R1204 B.n493 B.n43 585
R1205 B.n491 B.n490 585
R1206 B.n489 B.n46 585
R1207 B.n488 B.n487 585
R1208 B.n486 B.n47 585
R1209 B.n485 B.n484 585
R1210 B.n483 B.n48 585
R1211 B.n482 B.n481 585
R1212 B.n480 B.n49 585
R1213 B.n479 B.n478 585
R1214 B.n477 B.n50 585
R1215 B.n476 B.n475 585
R1216 B.n474 B.n51 585
R1217 B.n473 B.n472 585
R1218 B.n471 B.n52 585
R1219 B.n470 B.n469 585
R1220 B.n468 B.n53 585
R1221 B.n467 B.n466 585
R1222 B.n465 B.n54 585
R1223 B.n464 B.n463 585
R1224 B.n462 B.n55 585
R1225 B.n461 B.n460 585
R1226 B.n459 B.n56 585
R1227 B.n458 B.n457 585
R1228 B.n456 B.n57 585
R1229 B.n455 B.n454 585
R1230 B.n453 B.n58 585
R1231 B.n452 B.n451 585
R1232 B.n450 B.n59 585
R1233 B.n449 B.n448 585
R1234 B.n447 B.n60 585
R1235 B.n446 B.n445 585
R1236 B.n444 B.n61 585
R1237 B.n443 B.n442 585
R1238 B.n441 B.n62 585
R1239 B.n440 B.n439 585
R1240 B.n438 B.n63 585
R1241 B.n437 B.n436 585
R1242 B.n435 B.n64 585
R1243 B.n434 B.n433 585
R1244 B.n432 B.n65 585
R1245 B.n431 B.n430 585
R1246 B.n429 B.n66 585
R1247 B.n428 B.n427 585
R1248 B.n426 B.n67 585
R1249 B.n425 B.n424 585
R1250 B.n423 B.n68 585
R1251 B.n422 B.n421 585
R1252 B.n420 B.n69 585
R1253 B.n419 B.n418 585
R1254 B.n417 B.n70 585
R1255 B.n583 B.n582 585
R1256 B.n584 B.n11 585
R1257 B.n586 B.n585 585
R1258 B.n587 B.n10 585
R1259 B.n589 B.n588 585
R1260 B.n590 B.n9 585
R1261 B.n592 B.n591 585
R1262 B.n593 B.n8 585
R1263 B.n595 B.n594 585
R1264 B.n596 B.n7 585
R1265 B.n598 B.n597 585
R1266 B.n599 B.n6 585
R1267 B.n601 B.n600 585
R1268 B.n602 B.n5 585
R1269 B.n604 B.n603 585
R1270 B.n605 B.n4 585
R1271 B.n607 B.n606 585
R1272 B.n608 B.n3 585
R1273 B.n610 B.n609 585
R1274 B.n611 B.n0 585
R1275 B.n2 B.n1 585
R1276 B.n158 B.n157 585
R1277 B.n160 B.n159 585
R1278 B.n161 B.n156 585
R1279 B.n163 B.n162 585
R1280 B.n164 B.n155 585
R1281 B.n166 B.n165 585
R1282 B.n167 B.n154 585
R1283 B.n169 B.n168 585
R1284 B.n170 B.n153 585
R1285 B.n172 B.n171 585
R1286 B.n173 B.n152 585
R1287 B.n175 B.n174 585
R1288 B.n176 B.n151 585
R1289 B.n178 B.n177 585
R1290 B.n179 B.n150 585
R1291 B.n181 B.n180 585
R1292 B.n182 B.n149 585
R1293 B.n184 B.n183 585
R1294 B.n185 B.n148 585
R1295 B.n186 B.n185 502.111
R1296 B.n352 B.n91 502.111
R1297 B.n417 B.n416 502.111
R1298 B.n582 B.n581 502.111
R1299 B.n274 B.t1 465.442
R1300 B.n44 B.t5 465.442
R1301 B.n122 B.t10 465.442
R1302 B.n38 B.t8 465.442
R1303 B.n275 B.t2 423.938
R1304 B.n45 B.t4 423.938
R1305 B.n123 B.t11 423.938
R1306 B.n39 B.t7 423.938
R1307 B.n122 B.t9 402.031
R1308 B.n274 B.t0 402.031
R1309 B.n44 B.t3 402.031
R1310 B.n38 B.t6 402.031
R1311 B.n613 B.n612 256.663
R1312 B.n612 B.n611 235.042
R1313 B.n612 B.n2 235.042
R1314 B.n186 B.n147 163.367
R1315 B.n190 B.n147 163.367
R1316 B.n191 B.n190 163.367
R1317 B.n192 B.n191 163.367
R1318 B.n192 B.n145 163.367
R1319 B.n196 B.n145 163.367
R1320 B.n197 B.n196 163.367
R1321 B.n198 B.n197 163.367
R1322 B.n198 B.n143 163.367
R1323 B.n202 B.n143 163.367
R1324 B.n203 B.n202 163.367
R1325 B.n204 B.n203 163.367
R1326 B.n204 B.n141 163.367
R1327 B.n208 B.n141 163.367
R1328 B.n209 B.n208 163.367
R1329 B.n210 B.n209 163.367
R1330 B.n210 B.n139 163.367
R1331 B.n214 B.n139 163.367
R1332 B.n215 B.n214 163.367
R1333 B.n216 B.n215 163.367
R1334 B.n216 B.n137 163.367
R1335 B.n220 B.n137 163.367
R1336 B.n221 B.n220 163.367
R1337 B.n222 B.n221 163.367
R1338 B.n222 B.n135 163.367
R1339 B.n226 B.n135 163.367
R1340 B.n227 B.n226 163.367
R1341 B.n228 B.n227 163.367
R1342 B.n228 B.n133 163.367
R1343 B.n232 B.n133 163.367
R1344 B.n233 B.n232 163.367
R1345 B.n234 B.n233 163.367
R1346 B.n234 B.n131 163.367
R1347 B.n238 B.n131 163.367
R1348 B.n239 B.n238 163.367
R1349 B.n240 B.n239 163.367
R1350 B.n240 B.n129 163.367
R1351 B.n244 B.n129 163.367
R1352 B.n245 B.n244 163.367
R1353 B.n246 B.n245 163.367
R1354 B.n246 B.n127 163.367
R1355 B.n250 B.n127 163.367
R1356 B.n251 B.n250 163.367
R1357 B.n252 B.n251 163.367
R1358 B.n252 B.n125 163.367
R1359 B.n256 B.n125 163.367
R1360 B.n257 B.n256 163.367
R1361 B.n258 B.n257 163.367
R1362 B.n258 B.n121 163.367
R1363 B.n263 B.n121 163.367
R1364 B.n264 B.n263 163.367
R1365 B.n265 B.n264 163.367
R1366 B.n265 B.n119 163.367
R1367 B.n269 B.n119 163.367
R1368 B.n270 B.n269 163.367
R1369 B.n271 B.n270 163.367
R1370 B.n271 B.n117 163.367
R1371 B.n278 B.n117 163.367
R1372 B.n279 B.n278 163.367
R1373 B.n280 B.n279 163.367
R1374 B.n280 B.n115 163.367
R1375 B.n284 B.n115 163.367
R1376 B.n285 B.n284 163.367
R1377 B.n286 B.n285 163.367
R1378 B.n286 B.n113 163.367
R1379 B.n290 B.n113 163.367
R1380 B.n291 B.n290 163.367
R1381 B.n292 B.n291 163.367
R1382 B.n292 B.n111 163.367
R1383 B.n296 B.n111 163.367
R1384 B.n297 B.n296 163.367
R1385 B.n298 B.n297 163.367
R1386 B.n298 B.n109 163.367
R1387 B.n302 B.n109 163.367
R1388 B.n303 B.n302 163.367
R1389 B.n304 B.n303 163.367
R1390 B.n304 B.n107 163.367
R1391 B.n308 B.n107 163.367
R1392 B.n309 B.n308 163.367
R1393 B.n310 B.n309 163.367
R1394 B.n310 B.n105 163.367
R1395 B.n314 B.n105 163.367
R1396 B.n315 B.n314 163.367
R1397 B.n316 B.n315 163.367
R1398 B.n316 B.n103 163.367
R1399 B.n320 B.n103 163.367
R1400 B.n321 B.n320 163.367
R1401 B.n322 B.n321 163.367
R1402 B.n322 B.n101 163.367
R1403 B.n326 B.n101 163.367
R1404 B.n327 B.n326 163.367
R1405 B.n328 B.n327 163.367
R1406 B.n328 B.n99 163.367
R1407 B.n332 B.n99 163.367
R1408 B.n333 B.n332 163.367
R1409 B.n334 B.n333 163.367
R1410 B.n334 B.n97 163.367
R1411 B.n338 B.n97 163.367
R1412 B.n339 B.n338 163.367
R1413 B.n340 B.n339 163.367
R1414 B.n340 B.n95 163.367
R1415 B.n344 B.n95 163.367
R1416 B.n345 B.n344 163.367
R1417 B.n346 B.n345 163.367
R1418 B.n346 B.n93 163.367
R1419 B.n350 B.n93 163.367
R1420 B.n351 B.n350 163.367
R1421 B.n352 B.n351 163.367
R1422 B.n416 B.n71 163.367
R1423 B.n412 B.n71 163.367
R1424 B.n412 B.n411 163.367
R1425 B.n411 B.n410 163.367
R1426 B.n410 B.n73 163.367
R1427 B.n406 B.n73 163.367
R1428 B.n406 B.n405 163.367
R1429 B.n405 B.n404 163.367
R1430 B.n404 B.n75 163.367
R1431 B.n400 B.n75 163.367
R1432 B.n400 B.n399 163.367
R1433 B.n399 B.n398 163.367
R1434 B.n398 B.n77 163.367
R1435 B.n394 B.n77 163.367
R1436 B.n394 B.n393 163.367
R1437 B.n393 B.n392 163.367
R1438 B.n392 B.n79 163.367
R1439 B.n388 B.n79 163.367
R1440 B.n388 B.n387 163.367
R1441 B.n387 B.n386 163.367
R1442 B.n386 B.n81 163.367
R1443 B.n382 B.n81 163.367
R1444 B.n382 B.n381 163.367
R1445 B.n381 B.n380 163.367
R1446 B.n380 B.n83 163.367
R1447 B.n376 B.n83 163.367
R1448 B.n376 B.n375 163.367
R1449 B.n375 B.n374 163.367
R1450 B.n374 B.n85 163.367
R1451 B.n370 B.n85 163.367
R1452 B.n370 B.n369 163.367
R1453 B.n369 B.n368 163.367
R1454 B.n368 B.n87 163.367
R1455 B.n364 B.n87 163.367
R1456 B.n364 B.n363 163.367
R1457 B.n363 B.n362 163.367
R1458 B.n362 B.n89 163.367
R1459 B.n358 B.n89 163.367
R1460 B.n358 B.n357 163.367
R1461 B.n357 B.n356 163.367
R1462 B.n356 B.n91 163.367
R1463 B.n581 B.n580 163.367
R1464 B.n580 B.n13 163.367
R1465 B.n576 B.n13 163.367
R1466 B.n576 B.n575 163.367
R1467 B.n575 B.n574 163.367
R1468 B.n574 B.n15 163.367
R1469 B.n570 B.n15 163.367
R1470 B.n570 B.n569 163.367
R1471 B.n569 B.n568 163.367
R1472 B.n568 B.n17 163.367
R1473 B.n564 B.n17 163.367
R1474 B.n564 B.n563 163.367
R1475 B.n563 B.n562 163.367
R1476 B.n562 B.n19 163.367
R1477 B.n558 B.n19 163.367
R1478 B.n558 B.n557 163.367
R1479 B.n557 B.n556 163.367
R1480 B.n556 B.n21 163.367
R1481 B.n552 B.n21 163.367
R1482 B.n552 B.n551 163.367
R1483 B.n551 B.n550 163.367
R1484 B.n550 B.n23 163.367
R1485 B.n546 B.n23 163.367
R1486 B.n546 B.n545 163.367
R1487 B.n545 B.n544 163.367
R1488 B.n544 B.n25 163.367
R1489 B.n540 B.n25 163.367
R1490 B.n540 B.n539 163.367
R1491 B.n539 B.n538 163.367
R1492 B.n538 B.n27 163.367
R1493 B.n534 B.n27 163.367
R1494 B.n534 B.n533 163.367
R1495 B.n533 B.n532 163.367
R1496 B.n532 B.n29 163.367
R1497 B.n528 B.n29 163.367
R1498 B.n528 B.n527 163.367
R1499 B.n527 B.n526 163.367
R1500 B.n526 B.n31 163.367
R1501 B.n522 B.n31 163.367
R1502 B.n522 B.n521 163.367
R1503 B.n521 B.n520 163.367
R1504 B.n520 B.n33 163.367
R1505 B.n516 B.n33 163.367
R1506 B.n516 B.n515 163.367
R1507 B.n515 B.n514 163.367
R1508 B.n514 B.n35 163.367
R1509 B.n510 B.n35 163.367
R1510 B.n510 B.n509 163.367
R1511 B.n509 B.n508 163.367
R1512 B.n508 B.n37 163.367
R1513 B.n503 B.n37 163.367
R1514 B.n503 B.n502 163.367
R1515 B.n502 B.n501 163.367
R1516 B.n501 B.n41 163.367
R1517 B.n497 B.n41 163.367
R1518 B.n497 B.n496 163.367
R1519 B.n496 B.n495 163.367
R1520 B.n495 B.n43 163.367
R1521 B.n490 B.n43 163.367
R1522 B.n490 B.n489 163.367
R1523 B.n489 B.n488 163.367
R1524 B.n488 B.n47 163.367
R1525 B.n484 B.n47 163.367
R1526 B.n484 B.n483 163.367
R1527 B.n483 B.n482 163.367
R1528 B.n482 B.n49 163.367
R1529 B.n478 B.n49 163.367
R1530 B.n478 B.n477 163.367
R1531 B.n477 B.n476 163.367
R1532 B.n476 B.n51 163.367
R1533 B.n472 B.n51 163.367
R1534 B.n472 B.n471 163.367
R1535 B.n471 B.n470 163.367
R1536 B.n470 B.n53 163.367
R1537 B.n466 B.n53 163.367
R1538 B.n466 B.n465 163.367
R1539 B.n465 B.n464 163.367
R1540 B.n464 B.n55 163.367
R1541 B.n460 B.n55 163.367
R1542 B.n460 B.n459 163.367
R1543 B.n459 B.n458 163.367
R1544 B.n458 B.n57 163.367
R1545 B.n454 B.n57 163.367
R1546 B.n454 B.n453 163.367
R1547 B.n453 B.n452 163.367
R1548 B.n452 B.n59 163.367
R1549 B.n448 B.n59 163.367
R1550 B.n448 B.n447 163.367
R1551 B.n447 B.n446 163.367
R1552 B.n446 B.n61 163.367
R1553 B.n442 B.n61 163.367
R1554 B.n442 B.n441 163.367
R1555 B.n441 B.n440 163.367
R1556 B.n440 B.n63 163.367
R1557 B.n436 B.n63 163.367
R1558 B.n436 B.n435 163.367
R1559 B.n435 B.n434 163.367
R1560 B.n434 B.n65 163.367
R1561 B.n430 B.n65 163.367
R1562 B.n430 B.n429 163.367
R1563 B.n429 B.n428 163.367
R1564 B.n428 B.n67 163.367
R1565 B.n424 B.n67 163.367
R1566 B.n424 B.n423 163.367
R1567 B.n423 B.n422 163.367
R1568 B.n422 B.n69 163.367
R1569 B.n418 B.n69 163.367
R1570 B.n418 B.n417 163.367
R1571 B.n582 B.n11 163.367
R1572 B.n586 B.n11 163.367
R1573 B.n587 B.n586 163.367
R1574 B.n588 B.n587 163.367
R1575 B.n588 B.n9 163.367
R1576 B.n592 B.n9 163.367
R1577 B.n593 B.n592 163.367
R1578 B.n594 B.n593 163.367
R1579 B.n594 B.n7 163.367
R1580 B.n598 B.n7 163.367
R1581 B.n599 B.n598 163.367
R1582 B.n600 B.n599 163.367
R1583 B.n600 B.n5 163.367
R1584 B.n604 B.n5 163.367
R1585 B.n605 B.n604 163.367
R1586 B.n606 B.n605 163.367
R1587 B.n606 B.n3 163.367
R1588 B.n610 B.n3 163.367
R1589 B.n611 B.n610 163.367
R1590 B.n157 B.n2 163.367
R1591 B.n160 B.n157 163.367
R1592 B.n161 B.n160 163.367
R1593 B.n162 B.n161 163.367
R1594 B.n162 B.n155 163.367
R1595 B.n166 B.n155 163.367
R1596 B.n167 B.n166 163.367
R1597 B.n168 B.n167 163.367
R1598 B.n168 B.n153 163.367
R1599 B.n172 B.n153 163.367
R1600 B.n173 B.n172 163.367
R1601 B.n174 B.n173 163.367
R1602 B.n174 B.n151 163.367
R1603 B.n178 B.n151 163.367
R1604 B.n179 B.n178 163.367
R1605 B.n180 B.n179 163.367
R1606 B.n180 B.n149 163.367
R1607 B.n184 B.n149 163.367
R1608 B.n185 B.n184 163.367
R1609 B.n261 B.n123 59.5399
R1610 B.n276 B.n275 59.5399
R1611 B.n492 B.n45 59.5399
R1612 B.n506 B.n39 59.5399
R1613 B.n123 B.n122 41.5035
R1614 B.n275 B.n274 41.5035
R1615 B.n45 B.n44 41.5035
R1616 B.n39 B.n38 41.5035
R1617 B.n583 B.n12 32.6249
R1618 B.n415 B.n70 32.6249
R1619 B.n354 B.n353 32.6249
R1620 B.n187 B.n148 32.6249
R1621 B B.n613 18.0485
R1622 B.n584 B.n583 10.6151
R1623 B.n585 B.n584 10.6151
R1624 B.n585 B.n10 10.6151
R1625 B.n589 B.n10 10.6151
R1626 B.n590 B.n589 10.6151
R1627 B.n591 B.n590 10.6151
R1628 B.n591 B.n8 10.6151
R1629 B.n595 B.n8 10.6151
R1630 B.n596 B.n595 10.6151
R1631 B.n597 B.n596 10.6151
R1632 B.n597 B.n6 10.6151
R1633 B.n601 B.n6 10.6151
R1634 B.n602 B.n601 10.6151
R1635 B.n603 B.n602 10.6151
R1636 B.n603 B.n4 10.6151
R1637 B.n607 B.n4 10.6151
R1638 B.n608 B.n607 10.6151
R1639 B.n609 B.n608 10.6151
R1640 B.n609 B.n0 10.6151
R1641 B.n579 B.n12 10.6151
R1642 B.n579 B.n578 10.6151
R1643 B.n578 B.n577 10.6151
R1644 B.n577 B.n14 10.6151
R1645 B.n573 B.n14 10.6151
R1646 B.n573 B.n572 10.6151
R1647 B.n572 B.n571 10.6151
R1648 B.n571 B.n16 10.6151
R1649 B.n567 B.n16 10.6151
R1650 B.n567 B.n566 10.6151
R1651 B.n566 B.n565 10.6151
R1652 B.n565 B.n18 10.6151
R1653 B.n561 B.n18 10.6151
R1654 B.n561 B.n560 10.6151
R1655 B.n560 B.n559 10.6151
R1656 B.n559 B.n20 10.6151
R1657 B.n555 B.n20 10.6151
R1658 B.n555 B.n554 10.6151
R1659 B.n554 B.n553 10.6151
R1660 B.n553 B.n22 10.6151
R1661 B.n549 B.n22 10.6151
R1662 B.n549 B.n548 10.6151
R1663 B.n548 B.n547 10.6151
R1664 B.n547 B.n24 10.6151
R1665 B.n543 B.n24 10.6151
R1666 B.n543 B.n542 10.6151
R1667 B.n542 B.n541 10.6151
R1668 B.n541 B.n26 10.6151
R1669 B.n537 B.n26 10.6151
R1670 B.n537 B.n536 10.6151
R1671 B.n536 B.n535 10.6151
R1672 B.n535 B.n28 10.6151
R1673 B.n531 B.n28 10.6151
R1674 B.n531 B.n530 10.6151
R1675 B.n530 B.n529 10.6151
R1676 B.n529 B.n30 10.6151
R1677 B.n525 B.n30 10.6151
R1678 B.n525 B.n524 10.6151
R1679 B.n524 B.n523 10.6151
R1680 B.n523 B.n32 10.6151
R1681 B.n519 B.n32 10.6151
R1682 B.n519 B.n518 10.6151
R1683 B.n518 B.n517 10.6151
R1684 B.n517 B.n34 10.6151
R1685 B.n513 B.n34 10.6151
R1686 B.n513 B.n512 10.6151
R1687 B.n512 B.n511 10.6151
R1688 B.n511 B.n36 10.6151
R1689 B.n507 B.n36 10.6151
R1690 B.n505 B.n504 10.6151
R1691 B.n504 B.n40 10.6151
R1692 B.n500 B.n40 10.6151
R1693 B.n500 B.n499 10.6151
R1694 B.n499 B.n498 10.6151
R1695 B.n498 B.n42 10.6151
R1696 B.n494 B.n42 10.6151
R1697 B.n494 B.n493 10.6151
R1698 B.n491 B.n46 10.6151
R1699 B.n487 B.n46 10.6151
R1700 B.n487 B.n486 10.6151
R1701 B.n486 B.n485 10.6151
R1702 B.n485 B.n48 10.6151
R1703 B.n481 B.n48 10.6151
R1704 B.n481 B.n480 10.6151
R1705 B.n480 B.n479 10.6151
R1706 B.n479 B.n50 10.6151
R1707 B.n475 B.n50 10.6151
R1708 B.n475 B.n474 10.6151
R1709 B.n474 B.n473 10.6151
R1710 B.n473 B.n52 10.6151
R1711 B.n469 B.n52 10.6151
R1712 B.n469 B.n468 10.6151
R1713 B.n468 B.n467 10.6151
R1714 B.n467 B.n54 10.6151
R1715 B.n463 B.n54 10.6151
R1716 B.n463 B.n462 10.6151
R1717 B.n462 B.n461 10.6151
R1718 B.n461 B.n56 10.6151
R1719 B.n457 B.n56 10.6151
R1720 B.n457 B.n456 10.6151
R1721 B.n456 B.n455 10.6151
R1722 B.n455 B.n58 10.6151
R1723 B.n451 B.n58 10.6151
R1724 B.n451 B.n450 10.6151
R1725 B.n450 B.n449 10.6151
R1726 B.n449 B.n60 10.6151
R1727 B.n445 B.n60 10.6151
R1728 B.n445 B.n444 10.6151
R1729 B.n444 B.n443 10.6151
R1730 B.n443 B.n62 10.6151
R1731 B.n439 B.n62 10.6151
R1732 B.n439 B.n438 10.6151
R1733 B.n438 B.n437 10.6151
R1734 B.n437 B.n64 10.6151
R1735 B.n433 B.n64 10.6151
R1736 B.n433 B.n432 10.6151
R1737 B.n432 B.n431 10.6151
R1738 B.n431 B.n66 10.6151
R1739 B.n427 B.n66 10.6151
R1740 B.n427 B.n426 10.6151
R1741 B.n426 B.n425 10.6151
R1742 B.n425 B.n68 10.6151
R1743 B.n421 B.n68 10.6151
R1744 B.n421 B.n420 10.6151
R1745 B.n420 B.n419 10.6151
R1746 B.n419 B.n70 10.6151
R1747 B.n415 B.n414 10.6151
R1748 B.n414 B.n413 10.6151
R1749 B.n413 B.n72 10.6151
R1750 B.n409 B.n72 10.6151
R1751 B.n409 B.n408 10.6151
R1752 B.n408 B.n407 10.6151
R1753 B.n407 B.n74 10.6151
R1754 B.n403 B.n74 10.6151
R1755 B.n403 B.n402 10.6151
R1756 B.n402 B.n401 10.6151
R1757 B.n401 B.n76 10.6151
R1758 B.n397 B.n76 10.6151
R1759 B.n397 B.n396 10.6151
R1760 B.n396 B.n395 10.6151
R1761 B.n395 B.n78 10.6151
R1762 B.n391 B.n78 10.6151
R1763 B.n391 B.n390 10.6151
R1764 B.n390 B.n389 10.6151
R1765 B.n389 B.n80 10.6151
R1766 B.n385 B.n80 10.6151
R1767 B.n385 B.n384 10.6151
R1768 B.n384 B.n383 10.6151
R1769 B.n383 B.n82 10.6151
R1770 B.n379 B.n82 10.6151
R1771 B.n379 B.n378 10.6151
R1772 B.n378 B.n377 10.6151
R1773 B.n377 B.n84 10.6151
R1774 B.n373 B.n84 10.6151
R1775 B.n373 B.n372 10.6151
R1776 B.n372 B.n371 10.6151
R1777 B.n371 B.n86 10.6151
R1778 B.n367 B.n86 10.6151
R1779 B.n367 B.n366 10.6151
R1780 B.n366 B.n365 10.6151
R1781 B.n365 B.n88 10.6151
R1782 B.n361 B.n88 10.6151
R1783 B.n361 B.n360 10.6151
R1784 B.n360 B.n359 10.6151
R1785 B.n359 B.n90 10.6151
R1786 B.n355 B.n90 10.6151
R1787 B.n355 B.n354 10.6151
R1788 B.n158 B.n1 10.6151
R1789 B.n159 B.n158 10.6151
R1790 B.n159 B.n156 10.6151
R1791 B.n163 B.n156 10.6151
R1792 B.n164 B.n163 10.6151
R1793 B.n165 B.n164 10.6151
R1794 B.n165 B.n154 10.6151
R1795 B.n169 B.n154 10.6151
R1796 B.n170 B.n169 10.6151
R1797 B.n171 B.n170 10.6151
R1798 B.n171 B.n152 10.6151
R1799 B.n175 B.n152 10.6151
R1800 B.n176 B.n175 10.6151
R1801 B.n177 B.n176 10.6151
R1802 B.n177 B.n150 10.6151
R1803 B.n181 B.n150 10.6151
R1804 B.n182 B.n181 10.6151
R1805 B.n183 B.n182 10.6151
R1806 B.n183 B.n148 10.6151
R1807 B.n188 B.n187 10.6151
R1808 B.n189 B.n188 10.6151
R1809 B.n189 B.n146 10.6151
R1810 B.n193 B.n146 10.6151
R1811 B.n194 B.n193 10.6151
R1812 B.n195 B.n194 10.6151
R1813 B.n195 B.n144 10.6151
R1814 B.n199 B.n144 10.6151
R1815 B.n200 B.n199 10.6151
R1816 B.n201 B.n200 10.6151
R1817 B.n201 B.n142 10.6151
R1818 B.n205 B.n142 10.6151
R1819 B.n206 B.n205 10.6151
R1820 B.n207 B.n206 10.6151
R1821 B.n207 B.n140 10.6151
R1822 B.n211 B.n140 10.6151
R1823 B.n212 B.n211 10.6151
R1824 B.n213 B.n212 10.6151
R1825 B.n213 B.n138 10.6151
R1826 B.n217 B.n138 10.6151
R1827 B.n218 B.n217 10.6151
R1828 B.n219 B.n218 10.6151
R1829 B.n219 B.n136 10.6151
R1830 B.n223 B.n136 10.6151
R1831 B.n224 B.n223 10.6151
R1832 B.n225 B.n224 10.6151
R1833 B.n225 B.n134 10.6151
R1834 B.n229 B.n134 10.6151
R1835 B.n230 B.n229 10.6151
R1836 B.n231 B.n230 10.6151
R1837 B.n231 B.n132 10.6151
R1838 B.n235 B.n132 10.6151
R1839 B.n236 B.n235 10.6151
R1840 B.n237 B.n236 10.6151
R1841 B.n237 B.n130 10.6151
R1842 B.n241 B.n130 10.6151
R1843 B.n242 B.n241 10.6151
R1844 B.n243 B.n242 10.6151
R1845 B.n243 B.n128 10.6151
R1846 B.n247 B.n128 10.6151
R1847 B.n248 B.n247 10.6151
R1848 B.n249 B.n248 10.6151
R1849 B.n249 B.n126 10.6151
R1850 B.n253 B.n126 10.6151
R1851 B.n254 B.n253 10.6151
R1852 B.n255 B.n254 10.6151
R1853 B.n255 B.n124 10.6151
R1854 B.n259 B.n124 10.6151
R1855 B.n260 B.n259 10.6151
R1856 B.n262 B.n120 10.6151
R1857 B.n266 B.n120 10.6151
R1858 B.n267 B.n266 10.6151
R1859 B.n268 B.n267 10.6151
R1860 B.n268 B.n118 10.6151
R1861 B.n272 B.n118 10.6151
R1862 B.n273 B.n272 10.6151
R1863 B.n277 B.n273 10.6151
R1864 B.n281 B.n116 10.6151
R1865 B.n282 B.n281 10.6151
R1866 B.n283 B.n282 10.6151
R1867 B.n283 B.n114 10.6151
R1868 B.n287 B.n114 10.6151
R1869 B.n288 B.n287 10.6151
R1870 B.n289 B.n288 10.6151
R1871 B.n289 B.n112 10.6151
R1872 B.n293 B.n112 10.6151
R1873 B.n294 B.n293 10.6151
R1874 B.n295 B.n294 10.6151
R1875 B.n295 B.n110 10.6151
R1876 B.n299 B.n110 10.6151
R1877 B.n300 B.n299 10.6151
R1878 B.n301 B.n300 10.6151
R1879 B.n301 B.n108 10.6151
R1880 B.n305 B.n108 10.6151
R1881 B.n306 B.n305 10.6151
R1882 B.n307 B.n306 10.6151
R1883 B.n307 B.n106 10.6151
R1884 B.n311 B.n106 10.6151
R1885 B.n312 B.n311 10.6151
R1886 B.n313 B.n312 10.6151
R1887 B.n313 B.n104 10.6151
R1888 B.n317 B.n104 10.6151
R1889 B.n318 B.n317 10.6151
R1890 B.n319 B.n318 10.6151
R1891 B.n319 B.n102 10.6151
R1892 B.n323 B.n102 10.6151
R1893 B.n324 B.n323 10.6151
R1894 B.n325 B.n324 10.6151
R1895 B.n325 B.n100 10.6151
R1896 B.n329 B.n100 10.6151
R1897 B.n330 B.n329 10.6151
R1898 B.n331 B.n330 10.6151
R1899 B.n331 B.n98 10.6151
R1900 B.n335 B.n98 10.6151
R1901 B.n336 B.n335 10.6151
R1902 B.n337 B.n336 10.6151
R1903 B.n337 B.n96 10.6151
R1904 B.n341 B.n96 10.6151
R1905 B.n342 B.n341 10.6151
R1906 B.n343 B.n342 10.6151
R1907 B.n343 B.n94 10.6151
R1908 B.n347 B.n94 10.6151
R1909 B.n348 B.n347 10.6151
R1910 B.n349 B.n348 10.6151
R1911 B.n349 B.n92 10.6151
R1912 B.n353 B.n92 10.6151
R1913 B.n613 B.n0 8.11757
R1914 B.n613 B.n1 8.11757
R1915 B.n506 B.n505 6.5566
R1916 B.n493 B.n492 6.5566
R1917 B.n262 B.n261 6.5566
R1918 B.n277 B.n276 6.5566
R1919 B.n507 B.n506 4.05904
R1920 B.n492 B.n491 4.05904
R1921 B.n261 B.n260 4.05904
R1922 B.n276 B.n116 4.05904
C0 VP w_n1826_n3906# 2.73758f
C1 VDD2 VDD1 0.58179f
C2 VDD1 VTAIL 5.787529f
C3 VDD2 B 1.82585f
C4 VTAIL B 3.87479f
C5 VDD1 VN 0.14776f
C6 VP VDD2 0.300227f
C7 VP VTAIL 2.64089f
C8 VN B 0.947962f
C9 w_n1826_n3906# VDD2 1.89957f
C10 w_n1826_n3906# VTAIL 3.17726f
C11 VP VN 5.58392f
C12 VDD1 B 1.80276f
C13 w_n1826_n3906# VN 2.50669f
C14 VDD2 VTAIL 5.8309f
C15 VP VDD1 3.28343f
C16 VP B 1.32439f
C17 w_n1826_n3906# VDD1 1.8832f
C18 w_n1826_n3906# B 8.70964f
C19 VDD2 VN 3.13461f
C20 VN VTAIL 2.62645f
C21 VDD2 VSUBS 0.911017f
C22 VDD1 VSUBS 3.74428f
C23 VTAIL VSUBS 1.015633f
C24 VN VSUBS 8.279039f
C25 VP VSUBS 1.552968f
C26 B VSUBS 3.534734f
C27 w_n1826_n3906# VSUBS 87.4946f
C28 B.n0 VSUBS 0.005446f
C29 B.n1 VSUBS 0.005446f
C30 B.n2 VSUBS 0.008055f
C31 B.n3 VSUBS 0.006172f
C32 B.n4 VSUBS 0.006172f
C33 B.n5 VSUBS 0.006172f
C34 B.n6 VSUBS 0.006172f
C35 B.n7 VSUBS 0.006172f
C36 B.n8 VSUBS 0.006172f
C37 B.n9 VSUBS 0.006172f
C38 B.n10 VSUBS 0.006172f
C39 B.n11 VSUBS 0.006172f
C40 B.n12 VSUBS 0.015011f
C41 B.n13 VSUBS 0.006172f
C42 B.n14 VSUBS 0.006172f
C43 B.n15 VSUBS 0.006172f
C44 B.n16 VSUBS 0.006172f
C45 B.n17 VSUBS 0.006172f
C46 B.n18 VSUBS 0.006172f
C47 B.n19 VSUBS 0.006172f
C48 B.n20 VSUBS 0.006172f
C49 B.n21 VSUBS 0.006172f
C50 B.n22 VSUBS 0.006172f
C51 B.n23 VSUBS 0.006172f
C52 B.n24 VSUBS 0.006172f
C53 B.n25 VSUBS 0.006172f
C54 B.n26 VSUBS 0.006172f
C55 B.n27 VSUBS 0.006172f
C56 B.n28 VSUBS 0.006172f
C57 B.n29 VSUBS 0.006172f
C58 B.n30 VSUBS 0.006172f
C59 B.n31 VSUBS 0.006172f
C60 B.n32 VSUBS 0.006172f
C61 B.n33 VSUBS 0.006172f
C62 B.n34 VSUBS 0.006172f
C63 B.n35 VSUBS 0.006172f
C64 B.n36 VSUBS 0.006172f
C65 B.n37 VSUBS 0.006172f
C66 B.t7 VSUBS 0.24004f
C67 B.t8 VSUBS 0.261633f
C68 B.t6 VSUBS 1.026f
C69 B.n38 VSUBS 0.392316f
C70 B.n39 VSUBS 0.250962f
C71 B.n40 VSUBS 0.006172f
C72 B.n41 VSUBS 0.006172f
C73 B.n42 VSUBS 0.006172f
C74 B.n43 VSUBS 0.006172f
C75 B.t4 VSUBS 0.240043f
C76 B.t5 VSUBS 0.261636f
C77 B.t3 VSUBS 1.026f
C78 B.n44 VSUBS 0.392314f
C79 B.n45 VSUBS 0.250959f
C80 B.n46 VSUBS 0.006172f
C81 B.n47 VSUBS 0.006172f
C82 B.n48 VSUBS 0.006172f
C83 B.n49 VSUBS 0.006172f
C84 B.n50 VSUBS 0.006172f
C85 B.n51 VSUBS 0.006172f
C86 B.n52 VSUBS 0.006172f
C87 B.n53 VSUBS 0.006172f
C88 B.n54 VSUBS 0.006172f
C89 B.n55 VSUBS 0.006172f
C90 B.n56 VSUBS 0.006172f
C91 B.n57 VSUBS 0.006172f
C92 B.n58 VSUBS 0.006172f
C93 B.n59 VSUBS 0.006172f
C94 B.n60 VSUBS 0.006172f
C95 B.n61 VSUBS 0.006172f
C96 B.n62 VSUBS 0.006172f
C97 B.n63 VSUBS 0.006172f
C98 B.n64 VSUBS 0.006172f
C99 B.n65 VSUBS 0.006172f
C100 B.n66 VSUBS 0.006172f
C101 B.n67 VSUBS 0.006172f
C102 B.n68 VSUBS 0.006172f
C103 B.n69 VSUBS 0.006172f
C104 B.n70 VSUBS 0.015011f
C105 B.n71 VSUBS 0.006172f
C106 B.n72 VSUBS 0.006172f
C107 B.n73 VSUBS 0.006172f
C108 B.n74 VSUBS 0.006172f
C109 B.n75 VSUBS 0.006172f
C110 B.n76 VSUBS 0.006172f
C111 B.n77 VSUBS 0.006172f
C112 B.n78 VSUBS 0.006172f
C113 B.n79 VSUBS 0.006172f
C114 B.n80 VSUBS 0.006172f
C115 B.n81 VSUBS 0.006172f
C116 B.n82 VSUBS 0.006172f
C117 B.n83 VSUBS 0.006172f
C118 B.n84 VSUBS 0.006172f
C119 B.n85 VSUBS 0.006172f
C120 B.n86 VSUBS 0.006172f
C121 B.n87 VSUBS 0.006172f
C122 B.n88 VSUBS 0.006172f
C123 B.n89 VSUBS 0.006172f
C124 B.n90 VSUBS 0.006172f
C125 B.n91 VSUBS 0.013854f
C126 B.n92 VSUBS 0.006172f
C127 B.n93 VSUBS 0.006172f
C128 B.n94 VSUBS 0.006172f
C129 B.n95 VSUBS 0.006172f
C130 B.n96 VSUBS 0.006172f
C131 B.n97 VSUBS 0.006172f
C132 B.n98 VSUBS 0.006172f
C133 B.n99 VSUBS 0.006172f
C134 B.n100 VSUBS 0.006172f
C135 B.n101 VSUBS 0.006172f
C136 B.n102 VSUBS 0.006172f
C137 B.n103 VSUBS 0.006172f
C138 B.n104 VSUBS 0.006172f
C139 B.n105 VSUBS 0.006172f
C140 B.n106 VSUBS 0.006172f
C141 B.n107 VSUBS 0.006172f
C142 B.n108 VSUBS 0.006172f
C143 B.n109 VSUBS 0.006172f
C144 B.n110 VSUBS 0.006172f
C145 B.n111 VSUBS 0.006172f
C146 B.n112 VSUBS 0.006172f
C147 B.n113 VSUBS 0.006172f
C148 B.n114 VSUBS 0.006172f
C149 B.n115 VSUBS 0.006172f
C150 B.n116 VSUBS 0.004266f
C151 B.n117 VSUBS 0.006172f
C152 B.n118 VSUBS 0.006172f
C153 B.n119 VSUBS 0.006172f
C154 B.n120 VSUBS 0.006172f
C155 B.n121 VSUBS 0.006172f
C156 B.t11 VSUBS 0.24004f
C157 B.t10 VSUBS 0.261633f
C158 B.t9 VSUBS 1.026f
C159 B.n122 VSUBS 0.392316f
C160 B.n123 VSUBS 0.250962f
C161 B.n124 VSUBS 0.006172f
C162 B.n125 VSUBS 0.006172f
C163 B.n126 VSUBS 0.006172f
C164 B.n127 VSUBS 0.006172f
C165 B.n128 VSUBS 0.006172f
C166 B.n129 VSUBS 0.006172f
C167 B.n130 VSUBS 0.006172f
C168 B.n131 VSUBS 0.006172f
C169 B.n132 VSUBS 0.006172f
C170 B.n133 VSUBS 0.006172f
C171 B.n134 VSUBS 0.006172f
C172 B.n135 VSUBS 0.006172f
C173 B.n136 VSUBS 0.006172f
C174 B.n137 VSUBS 0.006172f
C175 B.n138 VSUBS 0.006172f
C176 B.n139 VSUBS 0.006172f
C177 B.n140 VSUBS 0.006172f
C178 B.n141 VSUBS 0.006172f
C179 B.n142 VSUBS 0.006172f
C180 B.n143 VSUBS 0.006172f
C181 B.n144 VSUBS 0.006172f
C182 B.n145 VSUBS 0.006172f
C183 B.n146 VSUBS 0.006172f
C184 B.n147 VSUBS 0.006172f
C185 B.n148 VSUBS 0.013854f
C186 B.n149 VSUBS 0.006172f
C187 B.n150 VSUBS 0.006172f
C188 B.n151 VSUBS 0.006172f
C189 B.n152 VSUBS 0.006172f
C190 B.n153 VSUBS 0.006172f
C191 B.n154 VSUBS 0.006172f
C192 B.n155 VSUBS 0.006172f
C193 B.n156 VSUBS 0.006172f
C194 B.n157 VSUBS 0.006172f
C195 B.n158 VSUBS 0.006172f
C196 B.n159 VSUBS 0.006172f
C197 B.n160 VSUBS 0.006172f
C198 B.n161 VSUBS 0.006172f
C199 B.n162 VSUBS 0.006172f
C200 B.n163 VSUBS 0.006172f
C201 B.n164 VSUBS 0.006172f
C202 B.n165 VSUBS 0.006172f
C203 B.n166 VSUBS 0.006172f
C204 B.n167 VSUBS 0.006172f
C205 B.n168 VSUBS 0.006172f
C206 B.n169 VSUBS 0.006172f
C207 B.n170 VSUBS 0.006172f
C208 B.n171 VSUBS 0.006172f
C209 B.n172 VSUBS 0.006172f
C210 B.n173 VSUBS 0.006172f
C211 B.n174 VSUBS 0.006172f
C212 B.n175 VSUBS 0.006172f
C213 B.n176 VSUBS 0.006172f
C214 B.n177 VSUBS 0.006172f
C215 B.n178 VSUBS 0.006172f
C216 B.n179 VSUBS 0.006172f
C217 B.n180 VSUBS 0.006172f
C218 B.n181 VSUBS 0.006172f
C219 B.n182 VSUBS 0.006172f
C220 B.n183 VSUBS 0.006172f
C221 B.n184 VSUBS 0.006172f
C222 B.n185 VSUBS 0.013854f
C223 B.n186 VSUBS 0.015011f
C224 B.n187 VSUBS 0.015011f
C225 B.n188 VSUBS 0.006172f
C226 B.n189 VSUBS 0.006172f
C227 B.n190 VSUBS 0.006172f
C228 B.n191 VSUBS 0.006172f
C229 B.n192 VSUBS 0.006172f
C230 B.n193 VSUBS 0.006172f
C231 B.n194 VSUBS 0.006172f
C232 B.n195 VSUBS 0.006172f
C233 B.n196 VSUBS 0.006172f
C234 B.n197 VSUBS 0.006172f
C235 B.n198 VSUBS 0.006172f
C236 B.n199 VSUBS 0.006172f
C237 B.n200 VSUBS 0.006172f
C238 B.n201 VSUBS 0.006172f
C239 B.n202 VSUBS 0.006172f
C240 B.n203 VSUBS 0.006172f
C241 B.n204 VSUBS 0.006172f
C242 B.n205 VSUBS 0.006172f
C243 B.n206 VSUBS 0.006172f
C244 B.n207 VSUBS 0.006172f
C245 B.n208 VSUBS 0.006172f
C246 B.n209 VSUBS 0.006172f
C247 B.n210 VSUBS 0.006172f
C248 B.n211 VSUBS 0.006172f
C249 B.n212 VSUBS 0.006172f
C250 B.n213 VSUBS 0.006172f
C251 B.n214 VSUBS 0.006172f
C252 B.n215 VSUBS 0.006172f
C253 B.n216 VSUBS 0.006172f
C254 B.n217 VSUBS 0.006172f
C255 B.n218 VSUBS 0.006172f
C256 B.n219 VSUBS 0.006172f
C257 B.n220 VSUBS 0.006172f
C258 B.n221 VSUBS 0.006172f
C259 B.n222 VSUBS 0.006172f
C260 B.n223 VSUBS 0.006172f
C261 B.n224 VSUBS 0.006172f
C262 B.n225 VSUBS 0.006172f
C263 B.n226 VSUBS 0.006172f
C264 B.n227 VSUBS 0.006172f
C265 B.n228 VSUBS 0.006172f
C266 B.n229 VSUBS 0.006172f
C267 B.n230 VSUBS 0.006172f
C268 B.n231 VSUBS 0.006172f
C269 B.n232 VSUBS 0.006172f
C270 B.n233 VSUBS 0.006172f
C271 B.n234 VSUBS 0.006172f
C272 B.n235 VSUBS 0.006172f
C273 B.n236 VSUBS 0.006172f
C274 B.n237 VSUBS 0.006172f
C275 B.n238 VSUBS 0.006172f
C276 B.n239 VSUBS 0.006172f
C277 B.n240 VSUBS 0.006172f
C278 B.n241 VSUBS 0.006172f
C279 B.n242 VSUBS 0.006172f
C280 B.n243 VSUBS 0.006172f
C281 B.n244 VSUBS 0.006172f
C282 B.n245 VSUBS 0.006172f
C283 B.n246 VSUBS 0.006172f
C284 B.n247 VSUBS 0.006172f
C285 B.n248 VSUBS 0.006172f
C286 B.n249 VSUBS 0.006172f
C287 B.n250 VSUBS 0.006172f
C288 B.n251 VSUBS 0.006172f
C289 B.n252 VSUBS 0.006172f
C290 B.n253 VSUBS 0.006172f
C291 B.n254 VSUBS 0.006172f
C292 B.n255 VSUBS 0.006172f
C293 B.n256 VSUBS 0.006172f
C294 B.n257 VSUBS 0.006172f
C295 B.n258 VSUBS 0.006172f
C296 B.n259 VSUBS 0.006172f
C297 B.n260 VSUBS 0.004266f
C298 B.n261 VSUBS 0.014301f
C299 B.n262 VSUBS 0.004992f
C300 B.n263 VSUBS 0.006172f
C301 B.n264 VSUBS 0.006172f
C302 B.n265 VSUBS 0.006172f
C303 B.n266 VSUBS 0.006172f
C304 B.n267 VSUBS 0.006172f
C305 B.n268 VSUBS 0.006172f
C306 B.n269 VSUBS 0.006172f
C307 B.n270 VSUBS 0.006172f
C308 B.n271 VSUBS 0.006172f
C309 B.n272 VSUBS 0.006172f
C310 B.n273 VSUBS 0.006172f
C311 B.t2 VSUBS 0.240043f
C312 B.t1 VSUBS 0.261636f
C313 B.t0 VSUBS 1.026f
C314 B.n274 VSUBS 0.392314f
C315 B.n275 VSUBS 0.250959f
C316 B.n276 VSUBS 0.014301f
C317 B.n277 VSUBS 0.004992f
C318 B.n278 VSUBS 0.006172f
C319 B.n279 VSUBS 0.006172f
C320 B.n280 VSUBS 0.006172f
C321 B.n281 VSUBS 0.006172f
C322 B.n282 VSUBS 0.006172f
C323 B.n283 VSUBS 0.006172f
C324 B.n284 VSUBS 0.006172f
C325 B.n285 VSUBS 0.006172f
C326 B.n286 VSUBS 0.006172f
C327 B.n287 VSUBS 0.006172f
C328 B.n288 VSUBS 0.006172f
C329 B.n289 VSUBS 0.006172f
C330 B.n290 VSUBS 0.006172f
C331 B.n291 VSUBS 0.006172f
C332 B.n292 VSUBS 0.006172f
C333 B.n293 VSUBS 0.006172f
C334 B.n294 VSUBS 0.006172f
C335 B.n295 VSUBS 0.006172f
C336 B.n296 VSUBS 0.006172f
C337 B.n297 VSUBS 0.006172f
C338 B.n298 VSUBS 0.006172f
C339 B.n299 VSUBS 0.006172f
C340 B.n300 VSUBS 0.006172f
C341 B.n301 VSUBS 0.006172f
C342 B.n302 VSUBS 0.006172f
C343 B.n303 VSUBS 0.006172f
C344 B.n304 VSUBS 0.006172f
C345 B.n305 VSUBS 0.006172f
C346 B.n306 VSUBS 0.006172f
C347 B.n307 VSUBS 0.006172f
C348 B.n308 VSUBS 0.006172f
C349 B.n309 VSUBS 0.006172f
C350 B.n310 VSUBS 0.006172f
C351 B.n311 VSUBS 0.006172f
C352 B.n312 VSUBS 0.006172f
C353 B.n313 VSUBS 0.006172f
C354 B.n314 VSUBS 0.006172f
C355 B.n315 VSUBS 0.006172f
C356 B.n316 VSUBS 0.006172f
C357 B.n317 VSUBS 0.006172f
C358 B.n318 VSUBS 0.006172f
C359 B.n319 VSUBS 0.006172f
C360 B.n320 VSUBS 0.006172f
C361 B.n321 VSUBS 0.006172f
C362 B.n322 VSUBS 0.006172f
C363 B.n323 VSUBS 0.006172f
C364 B.n324 VSUBS 0.006172f
C365 B.n325 VSUBS 0.006172f
C366 B.n326 VSUBS 0.006172f
C367 B.n327 VSUBS 0.006172f
C368 B.n328 VSUBS 0.006172f
C369 B.n329 VSUBS 0.006172f
C370 B.n330 VSUBS 0.006172f
C371 B.n331 VSUBS 0.006172f
C372 B.n332 VSUBS 0.006172f
C373 B.n333 VSUBS 0.006172f
C374 B.n334 VSUBS 0.006172f
C375 B.n335 VSUBS 0.006172f
C376 B.n336 VSUBS 0.006172f
C377 B.n337 VSUBS 0.006172f
C378 B.n338 VSUBS 0.006172f
C379 B.n339 VSUBS 0.006172f
C380 B.n340 VSUBS 0.006172f
C381 B.n341 VSUBS 0.006172f
C382 B.n342 VSUBS 0.006172f
C383 B.n343 VSUBS 0.006172f
C384 B.n344 VSUBS 0.006172f
C385 B.n345 VSUBS 0.006172f
C386 B.n346 VSUBS 0.006172f
C387 B.n347 VSUBS 0.006172f
C388 B.n348 VSUBS 0.006172f
C389 B.n349 VSUBS 0.006172f
C390 B.n350 VSUBS 0.006172f
C391 B.n351 VSUBS 0.006172f
C392 B.n352 VSUBS 0.015011f
C393 B.n353 VSUBS 0.014281f
C394 B.n354 VSUBS 0.014584f
C395 B.n355 VSUBS 0.006172f
C396 B.n356 VSUBS 0.006172f
C397 B.n357 VSUBS 0.006172f
C398 B.n358 VSUBS 0.006172f
C399 B.n359 VSUBS 0.006172f
C400 B.n360 VSUBS 0.006172f
C401 B.n361 VSUBS 0.006172f
C402 B.n362 VSUBS 0.006172f
C403 B.n363 VSUBS 0.006172f
C404 B.n364 VSUBS 0.006172f
C405 B.n365 VSUBS 0.006172f
C406 B.n366 VSUBS 0.006172f
C407 B.n367 VSUBS 0.006172f
C408 B.n368 VSUBS 0.006172f
C409 B.n369 VSUBS 0.006172f
C410 B.n370 VSUBS 0.006172f
C411 B.n371 VSUBS 0.006172f
C412 B.n372 VSUBS 0.006172f
C413 B.n373 VSUBS 0.006172f
C414 B.n374 VSUBS 0.006172f
C415 B.n375 VSUBS 0.006172f
C416 B.n376 VSUBS 0.006172f
C417 B.n377 VSUBS 0.006172f
C418 B.n378 VSUBS 0.006172f
C419 B.n379 VSUBS 0.006172f
C420 B.n380 VSUBS 0.006172f
C421 B.n381 VSUBS 0.006172f
C422 B.n382 VSUBS 0.006172f
C423 B.n383 VSUBS 0.006172f
C424 B.n384 VSUBS 0.006172f
C425 B.n385 VSUBS 0.006172f
C426 B.n386 VSUBS 0.006172f
C427 B.n387 VSUBS 0.006172f
C428 B.n388 VSUBS 0.006172f
C429 B.n389 VSUBS 0.006172f
C430 B.n390 VSUBS 0.006172f
C431 B.n391 VSUBS 0.006172f
C432 B.n392 VSUBS 0.006172f
C433 B.n393 VSUBS 0.006172f
C434 B.n394 VSUBS 0.006172f
C435 B.n395 VSUBS 0.006172f
C436 B.n396 VSUBS 0.006172f
C437 B.n397 VSUBS 0.006172f
C438 B.n398 VSUBS 0.006172f
C439 B.n399 VSUBS 0.006172f
C440 B.n400 VSUBS 0.006172f
C441 B.n401 VSUBS 0.006172f
C442 B.n402 VSUBS 0.006172f
C443 B.n403 VSUBS 0.006172f
C444 B.n404 VSUBS 0.006172f
C445 B.n405 VSUBS 0.006172f
C446 B.n406 VSUBS 0.006172f
C447 B.n407 VSUBS 0.006172f
C448 B.n408 VSUBS 0.006172f
C449 B.n409 VSUBS 0.006172f
C450 B.n410 VSUBS 0.006172f
C451 B.n411 VSUBS 0.006172f
C452 B.n412 VSUBS 0.006172f
C453 B.n413 VSUBS 0.006172f
C454 B.n414 VSUBS 0.006172f
C455 B.n415 VSUBS 0.013854f
C456 B.n416 VSUBS 0.013854f
C457 B.n417 VSUBS 0.015011f
C458 B.n418 VSUBS 0.006172f
C459 B.n419 VSUBS 0.006172f
C460 B.n420 VSUBS 0.006172f
C461 B.n421 VSUBS 0.006172f
C462 B.n422 VSUBS 0.006172f
C463 B.n423 VSUBS 0.006172f
C464 B.n424 VSUBS 0.006172f
C465 B.n425 VSUBS 0.006172f
C466 B.n426 VSUBS 0.006172f
C467 B.n427 VSUBS 0.006172f
C468 B.n428 VSUBS 0.006172f
C469 B.n429 VSUBS 0.006172f
C470 B.n430 VSUBS 0.006172f
C471 B.n431 VSUBS 0.006172f
C472 B.n432 VSUBS 0.006172f
C473 B.n433 VSUBS 0.006172f
C474 B.n434 VSUBS 0.006172f
C475 B.n435 VSUBS 0.006172f
C476 B.n436 VSUBS 0.006172f
C477 B.n437 VSUBS 0.006172f
C478 B.n438 VSUBS 0.006172f
C479 B.n439 VSUBS 0.006172f
C480 B.n440 VSUBS 0.006172f
C481 B.n441 VSUBS 0.006172f
C482 B.n442 VSUBS 0.006172f
C483 B.n443 VSUBS 0.006172f
C484 B.n444 VSUBS 0.006172f
C485 B.n445 VSUBS 0.006172f
C486 B.n446 VSUBS 0.006172f
C487 B.n447 VSUBS 0.006172f
C488 B.n448 VSUBS 0.006172f
C489 B.n449 VSUBS 0.006172f
C490 B.n450 VSUBS 0.006172f
C491 B.n451 VSUBS 0.006172f
C492 B.n452 VSUBS 0.006172f
C493 B.n453 VSUBS 0.006172f
C494 B.n454 VSUBS 0.006172f
C495 B.n455 VSUBS 0.006172f
C496 B.n456 VSUBS 0.006172f
C497 B.n457 VSUBS 0.006172f
C498 B.n458 VSUBS 0.006172f
C499 B.n459 VSUBS 0.006172f
C500 B.n460 VSUBS 0.006172f
C501 B.n461 VSUBS 0.006172f
C502 B.n462 VSUBS 0.006172f
C503 B.n463 VSUBS 0.006172f
C504 B.n464 VSUBS 0.006172f
C505 B.n465 VSUBS 0.006172f
C506 B.n466 VSUBS 0.006172f
C507 B.n467 VSUBS 0.006172f
C508 B.n468 VSUBS 0.006172f
C509 B.n469 VSUBS 0.006172f
C510 B.n470 VSUBS 0.006172f
C511 B.n471 VSUBS 0.006172f
C512 B.n472 VSUBS 0.006172f
C513 B.n473 VSUBS 0.006172f
C514 B.n474 VSUBS 0.006172f
C515 B.n475 VSUBS 0.006172f
C516 B.n476 VSUBS 0.006172f
C517 B.n477 VSUBS 0.006172f
C518 B.n478 VSUBS 0.006172f
C519 B.n479 VSUBS 0.006172f
C520 B.n480 VSUBS 0.006172f
C521 B.n481 VSUBS 0.006172f
C522 B.n482 VSUBS 0.006172f
C523 B.n483 VSUBS 0.006172f
C524 B.n484 VSUBS 0.006172f
C525 B.n485 VSUBS 0.006172f
C526 B.n486 VSUBS 0.006172f
C527 B.n487 VSUBS 0.006172f
C528 B.n488 VSUBS 0.006172f
C529 B.n489 VSUBS 0.006172f
C530 B.n490 VSUBS 0.006172f
C531 B.n491 VSUBS 0.004266f
C532 B.n492 VSUBS 0.014301f
C533 B.n493 VSUBS 0.004992f
C534 B.n494 VSUBS 0.006172f
C535 B.n495 VSUBS 0.006172f
C536 B.n496 VSUBS 0.006172f
C537 B.n497 VSUBS 0.006172f
C538 B.n498 VSUBS 0.006172f
C539 B.n499 VSUBS 0.006172f
C540 B.n500 VSUBS 0.006172f
C541 B.n501 VSUBS 0.006172f
C542 B.n502 VSUBS 0.006172f
C543 B.n503 VSUBS 0.006172f
C544 B.n504 VSUBS 0.006172f
C545 B.n505 VSUBS 0.004992f
C546 B.n506 VSUBS 0.014301f
C547 B.n507 VSUBS 0.004266f
C548 B.n508 VSUBS 0.006172f
C549 B.n509 VSUBS 0.006172f
C550 B.n510 VSUBS 0.006172f
C551 B.n511 VSUBS 0.006172f
C552 B.n512 VSUBS 0.006172f
C553 B.n513 VSUBS 0.006172f
C554 B.n514 VSUBS 0.006172f
C555 B.n515 VSUBS 0.006172f
C556 B.n516 VSUBS 0.006172f
C557 B.n517 VSUBS 0.006172f
C558 B.n518 VSUBS 0.006172f
C559 B.n519 VSUBS 0.006172f
C560 B.n520 VSUBS 0.006172f
C561 B.n521 VSUBS 0.006172f
C562 B.n522 VSUBS 0.006172f
C563 B.n523 VSUBS 0.006172f
C564 B.n524 VSUBS 0.006172f
C565 B.n525 VSUBS 0.006172f
C566 B.n526 VSUBS 0.006172f
C567 B.n527 VSUBS 0.006172f
C568 B.n528 VSUBS 0.006172f
C569 B.n529 VSUBS 0.006172f
C570 B.n530 VSUBS 0.006172f
C571 B.n531 VSUBS 0.006172f
C572 B.n532 VSUBS 0.006172f
C573 B.n533 VSUBS 0.006172f
C574 B.n534 VSUBS 0.006172f
C575 B.n535 VSUBS 0.006172f
C576 B.n536 VSUBS 0.006172f
C577 B.n537 VSUBS 0.006172f
C578 B.n538 VSUBS 0.006172f
C579 B.n539 VSUBS 0.006172f
C580 B.n540 VSUBS 0.006172f
C581 B.n541 VSUBS 0.006172f
C582 B.n542 VSUBS 0.006172f
C583 B.n543 VSUBS 0.006172f
C584 B.n544 VSUBS 0.006172f
C585 B.n545 VSUBS 0.006172f
C586 B.n546 VSUBS 0.006172f
C587 B.n547 VSUBS 0.006172f
C588 B.n548 VSUBS 0.006172f
C589 B.n549 VSUBS 0.006172f
C590 B.n550 VSUBS 0.006172f
C591 B.n551 VSUBS 0.006172f
C592 B.n552 VSUBS 0.006172f
C593 B.n553 VSUBS 0.006172f
C594 B.n554 VSUBS 0.006172f
C595 B.n555 VSUBS 0.006172f
C596 B.n556 VSUBS 0.006172f
C597 B.n557 VSUBS 0.006172f
C598 B.n558 VSUBS 0.006172f
C599 B.n559 VSUBS 0.006172f
C600 B.n560 VSUBS 0.006172f
C601 B.n561 VSUBS 0.006172f
C602 B.n562 VSUBS 0.006172f
C603 B.n563 VSUBS 0.006172f
C604 B.n564 VSUBS 0.006172f
C605 B.n565 VSUBS 0.006172f
C606 B.n566 VSUBS 0.006172f
C607 B.n567 VSUBS 0.006172f
C608 B.n568 VSUBS 0.006172f
C609 B.n569 VSUBS 0.006172f
C610 B.n570 VSUBS 0.006172f
C611 B.n571 VSUBS 0.006172f
C612 B.n572 VSUBS 0.006172f
C613 B.n573 VSUBS 0.006172f
C614 B.n574 VSUBS 0.006172f
C615 B.n575 VSUBS 0.006172f
C616 B.n576 VSUBS 0.006172f
C617 B.n577 VSUBS 0.006172f
C618 B.n578 VSUBS 0.006172f
C619 B.n579 VSUBS 0.006172f
C620 B.n580 VSUBS 0.006172f
C621 B.n581 VSUBS 0.015011f
C622 B.n582 VSUBS 0.013854f
C623 B.n583 VSUBS 0.013854f
C624 B.n584 VSUBS 0.006172f
C625 B.n585 VSUBS 0.006172f
C626 B.n586 VSUBS 0.006172f
C627 B.n587 VSUBS 0.006172f
C628 B.n588 VSUBS 0.006172f
C629 B.n589 VSUBS 0.006172f
C630 B.n590 VSUBS 0.006172f
C631 B.n591 VSUBS 0.006172f
C632 B.n592 VSUBS 0.006172f
C633 B.n593 VSUBS 0.006172f
C634 B.n594 VSUBS 0.006172f
C635 B.n595 VSUBS 0.006172f
C636 B.n596 VSUBS 0.006172f
C637 B.n597 VSUBS 0.006172f
C638 B.n598 VSUBS 0.006172f
C639 B.n599 VSUBS 0.006172f
C640 B.n600 VSUBS 0.006172f
C641 B.n601 VSUBS 0.006172f
C642 B.n602 VSUBS 0.006172f
C643 B.n603 VSUBS 0.006172f
C644 B.n604 VSUBS 0.006172f
C645 B.n605 VSUBS 0.006172f
C646 B.n606 VSUBS 0.006172f
C647 B.n607 VSUBS 0.006172f
C648 B.n608 VSUBS 0.006172f
C649 B.n609 VSUBS 0.006172f
C650 B.n610 VSUBS 0.006172f
C651 B.n611 VSUBS 0.008055f
C652 B.n612 VSUBS 0.00858f
C653 B.n613 VSUBS 0.017063f
C654 VDD2.n0 VSUBS 0.02053f
C655 VDD2.n1 VSUBS 0.019913f
C656 VDD2.n2 VSUBS 0.0107f
C657 VDD2.n3 VSUBS 0.025292f
C658 VDD2.n4 VSUBS 0.01133f
C659 VDD2.n5 VSUBS 0.019913f
C660 VDD2.n6 VSUBS 0.0107f
C661 VDD2.n7 VSUBS 0.025292f
C662 VDD2.n8 VSUBS 0.01133f
C663 VDD2.n9 VSUBS 0.019913f
C664 VDD2.n10 VSUBS 0.0107f
C665 VDD2.n11 VSUBS 0.025292f
C666 VDD2.n12 VSUBS 0.01133f
C667 VDD2.n13 VSUBS 0.019913f
C668 VDD2.n14 VSUBS 0.0107f
C669 VDD2.n15 VSUBS 0.025292f
C670 VDD2.n16 VSUBS 0.01133f
C671 VDD2.n17 VSUBS 0.019913f
C672 VDD2.n18 VSUBS 0.0107f
C673 VDD2.n19 VSUBS 0.025292f
C674 VDD2.n20 VSUBS 0.01133f
C675 VDD2.n21 VSUBS 0.019913f
C676 VDD2.n22 VSUBS 0.0107f
C677 VDD2.n23 VSUBS 0.025292f
C678 VDD2.n24 VSUBS 0.01133f
C679 VDD2.n25 VSUBS 0.138547f
C680 VDD2.t1 VSUBS 0.054129f
C681 VDD2.n26 VSUBS 0.018969f
C682 VDD2.n27 VSUBS 0.016089f
C683 VDD2.n28 VSUBS 0.0107f
C684 VDD2.n29 VSUBS 1.24344f
C685 VDD2.n30 VSUBS 0.019913f
C686 VDD2.n31 VSUBS 0.0107f
C687 VDD2.n32 VSUBS 0.01133f
C688 VDD2.n33 VSUBS 0.025292f
C689 VDD2.n34 VSUBS 0.025292f
C690 VDD2.n35 VSUBS 0.01133f
C691 VDD2.n36 VSUBS 0.0107f
C692 VDD2.n37 VSUBS 0.019913f
C693 VDD2.n38 VSUBS 0.019913f
C694 VDD2.n39 VSUBS 0.0107f
C695 VDD2.n40 VSUBS 0.01133f
C696 VDD2.n41 VSUBS 0.025292f
C697 VDD2.n42 VSUBS 0.025292f
C698 VDD2.n43 VSUBS 0.01133f
C699 VDD2.n44 VSUBS 0.0107f
C700 VDD2.n45 VSUBS 0.019913f
C701 VDD2.n46 VSUBS 0.019913f
C702 VDD2.n47 VSUBS 0.0107f
C703 VDD2.n48 VSUBS 0.01133f
C704 VDD2.n49 VSUBS 0.025292f
C705 VDD2.n50 VSUBS 0.025292f
C706 VDD2.n51 VSUBS 0.01133f
C707 VDD2.n52 VSUBS 0.0107f
C708 VDD2.n53 VSUBS 0.019913f
C709 VDD2.n54 VSUBS 0.019913f
C710 VDD2.n55 VSUBS 0.0107f
C711 VDD2.n56 VSUBS 0.01133f
C712 VDD2.n57 VSUBS 0.025292f
C713 VDD2.n58 VSUBS 0.025292f
C714 VDD2.n59 VSUBS 0.01133f
C715 VDD2.n60 VSUBS 0.0107f
C716 VDD2.n61 VSUBS 0.019913f
C717 VDD2.n62 VSUBS 0.019913f
C718 VDD2.n63 VSUBS 0.0107f
C719 VDD2.n64 VSUBS 0.01133f
C720 VDD2.n65 VSUBS 0.025292f
C721 VDD2.n66 VSUBS 0.025292f
C722 VDD2.n67 VSUBS 0.025292f
C723 VDD2.n68 VSUBS 0.01133f
C724 VDD2.n69 VSUBS 0.0107f
C725 VDD2.n70 VSUBS 0.019913f
C726 VDD2.n71 VSUBS 0.019913f
C727 VDD2.n72 VSUBS 0.0107f
C728 VDD2.n73 VSUBS 0.011015f
C729 VDD2.n74 VSUBS 0.011015f
C730 VDD2.n75 VSUBS 0.025292f
C731 VDD2.n76 VSUBS 0.056631f
C732 VDD2.n77 VSUBS 0.01133f
C733 VDD2.n78 VSUBS 0.0107f
C734 VDD2.n79 VSUBS 0.047387f
C735 VDD2.n80 VSUBS 0.612547f
C736 VDD2.n81 VSUBS 0.02053f
C737 VDD2.n82 VSUBS 0.019913f
C738 VDD2.n83 VSUBS 0.0107f
C739 VDD2.n84 VSUBS 0.025292f
C740 VDD2.n85 VSUBS 0.01133f
C741 VDD2.n86 VSUBS 0.019913f
C742 VDD2.n87 VSUBS 0.0107f
C743 VDD2.n88 VSUBS 0.025292f
C744 VDD2.n89 VSUBS 0.025292f
C745 VDD2.n90 VSUBS 0.01133f
C746 VDD2.n91 VSUBS 0.019913f
C747 VDD2.n92 VSUBS 0.0107f
C748 VDD2.n93 VSUBS 0.025292f
C749 VDD2.n94 VSUBS 0.01133f
C750 VDD2.n95 VSUBS 0.019913f
C751 VDD2.n96 VSUBS 0.0107f
C752 VDD2.n97 VSUBS 0.025292f
C753 VDD2.n98 VSUBS 0.01133f
C754 VDD2.n99 VSUBS 0.019913f
C755 VDD2.n100 VSUBS 0.0107f
C756 VDD2.n101 VSUBS 0.025292f
C757 VDD2.n102 VSUBS 0.01133f
C758 VDD2.n103 VSUBS 0.019913f
C759 VDD2.n104 VSUBS 0.0107f
C760 VDD2.n105 VSUBS 0.025292f
C761 VDD2.n106 VSUBS 0.01133f
C762 VDD2.n107 VSUBS 0.138547f
C763 VDD2.t0 VSUBS 0.054129f
C764 VDD2.n108 VSUBS 0.018969f
C765 VDD2.n109 VSUBS 0.016089f
C766 VDD2.n110 VSUBS 0.0107f
C767 VDD2.n111 VSUBS 1.24344f
C768 VDD2.n112 VSUBS 0.019913f
C769 VDD2.n113 VSUBS 0.0107f
C770 VDD2.n114 VSUBS 0.01133f
C771 VDD2.n115 VSUBS 0.025292f
C772 VDD2.n116 VSUBS 0.025292f
C773 VDD2.n117 VSUBS 0.01133f
C774 VDD2.n118 VSUBS 0.0107f
C775 VDD2.n119 VSUBS 0.019913f
C776 VDD2.n120 VSUBS 0.019913f
C777 VDD2.n121 VSUBS 0.0107f
C778 VDD2.n122 VSUBS 0.01133f
C779 VDD2.n123 VSUBS 0.025292f
C780 VDD2.n124 VSUBS 0.025292f
C781 VDD2.n125 VSUBS 0.01133f
C782 VDD2.n126 VSUBS 0.0107f
C783 VDD2.n127 VSUBS 0.019913f
C784 VDD2.n128 VSUBS 0.019913f
C785 VDD2.n129 VSUBS 0.0107f
C786 VDD2.n130 VSUBS 0.01133f
C787 VDD2.n131 VSUBS 0.025292f
C788 VDD2.n132 VSUBS 0.025292f
C789 VDD2.n133 VSUBS 0.01133f
C790 VDD2.n134 VSUBS 0.0107f
C791 VDD2.n135 VSUBS 0.019913f
C792 VDD2.n136 VSUBS 0.019913f
C793 VDD2.n137 VSUBS 0.0107f
C794 VDD2.n138 VSUBS 0.01133f
C795 VDD2.n139 VSUBS 0.025292f
C796 VDD2.n140 VSUBS 0.025292f
C797 VDD2.n141 VSUBS 0.01133f
C798 VDD2.n142 VSUBS 0.0107f
C799 VDD2.n143 VSUBS 0.019913f
C800 VDD2.n144 VSUBS 0.019913f
C801 VDD2.n145 VSUBS 0.0107f
C802 VDD2.n146 VSUBS 0.01133f
C803 VDD2.n147 VSUBS 0.025292f
C804 VDD2.n148 VSUBS 0.025292f
C805 VDD2.n149 VSUBS 0.01133f
C806 VDD2.n150 VSUBS 0.0107f
C807 VDD2.n151 VSUBS 0.019913f
C808 VDD2.n152 VSUBS 0.019913f
C809 VDD2.n153 VSUBS 0.0107f
C810 VDD2.n154 VSUBS 0.011015f
C811 VDD2.n155 VSUBS 0.011015f
C812 VDD2.n156 VSUBS 0.025292f
C813 VDD2.n157 VSUBS 0.056631f
C814 VDD2.n158 VSUBS 0.01133f
C815 VDD2.n159 VSUBS 0.0107f
C816 VDD2.n160 VSUBS 0.047387f
C817 VDD2.n161 VSUBS 0.042055f
C818 VDD2.n162 VSUBS 2.53748f
C819 VN.t0 VSUBS 3.61728f
C820 VN.t1 VSUBS 4.10327f
C821 VDD1.n0 VSUBS 0.02082f
C822 VDD1.n1 VSUBS 0.020193f
C823 VDD1.n2 VSUBS 0.010851f
C824 VDD1.n3 VSUBS 0.025648f
C825 VDD1.n4 VSUBS 0.011489f
C826 VDD1.n5 VSUBS 0.020193f
C827 VDD1.n6 VSUBS 0.010851f
C828 VDD1.n7 VSUBS 0.025648f
C829 VDD1.n8 VSUBS 0.025648f
C830 VDD1.n9 VSUBS 0.011489f
C831 VDD1.n10 VSUBS 0.020193f
C832 VDD1.n11 VSUBS 0.010851f
C833 VDD1.n12 VSUBS 0.025648f
C834 VDD1.n13 VSUBS 0.011489f
C835 VDD1.n14 VSUBS 0.020193f
C836 VDD1.n15 VSUBS 0.010851f
C837 VDD1.n16 VSUBS 0.025648f
C838 VDD1.n17 VSUBS 0.011489f
C839 VDD1.n18 VSUBS 0.020193f
C840 VDD1.n19 VSUBS 0.010851f
C841 VDD1.n20 VSUBS 0.025648f
C842 VDD1.n21 VSUBS 0.011489f
C843 VDD1.n22 VSUBS 0.020193f
C844 VDD1.n23 VSUBS 0.010851f
C845 VDD1.n24 VSUBS 0.025648f
C846 VDD1.n25 VSUBS 0.011489f
C847 VDD1.n26 VSUBS 0.140499f
C848 VDD1.t0 VSUBS 0.054891f
C849 VDD1.n27 VSUBS 0.019236f
C850 VDD1.n28 VSUBS 0.016316f
C851 VDD1.n29 VSUBS 0.010851f
C852 VDD1.n30 VSUBS 1.26097f
C853 VDD1.n31 VSUBS 0.020193f
C854 VDD1.n32 VSUBS 0.010851f
C855 VDD1.n33 VSUBS 0.011489f
C856 VDD1.n34 VSUBS 0.025648f
C857 VDD1.n35 VSUBS 0.025648f
C858 VDD1.n36 VSUBS 0.011489f
C859 VDD1.n37 VSUBS 0.010851f
C860 VDD1.n38 VSUBS 0.020193f
C861 VDD1.n39 VSUBS 0.020193f
C862 VDD1.n40 VSUBS 0.010851f
C863 VDD1.n41 VSUBS 0.011489f
C864 VDD1.n42 VSUBS 0.025648f
C865 VDD1.n43 VSUBS 0.025648f
C866 VDD1.n44 VSUBS 0.011489f
C867 VDD1.n45 VSUBS 0.010851f
C868 VDD1.n46 VSUBS 0.020193f
C869 VDD1.n47 VSUBS 0.020193f
C870 VDD1.n48 VSUBS 0.010851f
C871 VDD1.n49 VSUBS 0.011489f
C872 VDD1.n50 VSUBS 0.025648f
C873 VDD1.n51 VSUBS 0.025648f
C874 VDD1.n52 VSUBS 0.011489f
C875 VDD1.n53 VSUBS 0.010851f
C876 VDD1.n54 VSUBS 0.020193f
C877 VDD1.n55 VSUBS 0.020193f
C878 VDD1.n56 VSUBS 0.010851f
C879 VDD1.n57 VSUBS 0.011489f
C880 VDD1.n58 VSUBS 0.025648f
C881 VDD1.n59 VSUBS 0.025648f
C882 VDD1.n60 VSUBS 0.011489f
C883 VDD1.n61 VSUBS 0.010851f
C884 VDD1.n62 VSUBS 0.020193f
C885 VDD1.n63 VSUBS 0.020193f
C886 VDD1.n64 VSUBS 0.010851f
C887 VDD1.n65 VSUBS 0.011489f
C888 VDD1.n66 VSUBS 0.025648f
C889 VDD1.n67 VSUBS 0.025648f
C890 VDD1.n68 VSUBS 0.011489f
C891 VDD1.n69 VSUBS 0.010851f
C892 VDD1.n70 VSUBS 0.020193f
C893 VDD1.n71 VSUBS 0.020193f
C894 VDD1.n72 VSUBS 0.010851f
C895 VDD1.n73 VSUBS 0.01117f
C896 VDD1.n74 VSUBS 0.01117f
C897 VDD1.n75 VSUBS 0.025648f
C898 VDD1.n76 VSUBS 0.057429f
C899 VDD1.n77 VSUBS 0.011489f
C900 VDD1.n78 VSUBS 0.010851f
C901 VDD1.n79 VSUBS 0.048055f
C902 VDD1.n80 VSUBS 0.043406f
C903 VDD1.n81 VSUBS 0.02082f
C904 VDD1.n82 VSUBS 0.020193f
C905 VDD1.n83 VSUBS 0.010851f
C906 VDD1.n84 VSUBS 0.025648f
C907 VDD1.n85 VSUBS 0.011489f
C908 VDD1.n86 VSUBS 0.020193f
C909 VDD1.n87 VSUBS 0.010851f
C910 VDD1.n88 VSUBS 0.025648f
C911 VDD1.n89 VSUBS 0.011489f
C912 VDD1.n90 VSUBS 0.020193f
C913 VDD1.n91 VSUBS 0.010851f
C914 VDD1.n92 VSUBS 0.025648f
C915 VDD1.n93 VSUBS 0.011489f
C916 VDD1.n94 VSUBS 0.020193f
C917 VDD1.n95 VSUBS 0.010851f
C918 VDD1.n96 VSUBS 0.025648f
C919 VDD1.n97 VSUBS 0.011489f
C920 VDD1.n98 VSUBS 0.020193f
C921 VDD1.n99 VSUBS 0.010851f
C922 VDD1.n100 VSUBS 0.025648f
C923 VDD1.n101 VSUBS 0.011489f
C924 VDD1.n102 VSUBS 0.020193f
C925 VDD1.n103 VSUBS 0.010851f
C926 VDD1.n104 VSUBS 0.025648f
C927 VDD1.n105 VSUBS 0.011489f
C928 VDD1.n106 VSUBS 0.140499f
C929 VDD1.t1 VSUBS 0.054891f
C930 VDD1.n107 VSUBS 0.019236f
C931 VDD1.n108 VSUBS 0.016316f
C932 VDD1.n109 VSUBS 0.010851f
C933 VDD1.n110 VSUBS 1.26097f
C934 VDD1.n111 VSUBS 0.020193f
C935 VDD1.n112 VSUBS 0.010851f
C936 VDD1.n113 VSUBS 0.011489f
C937 VDD1.n114 VSUBS 0.025648f
C938 VDD1.n115 VSUBS 0.025648f
C939 VDD1.n116 VSUBS 0.011489f
C940 VDD1.n117 VSUBS 0.010851f
C941 VDD1.n118 VSUBS 0.020193f
C942 VDD1.n119 VSUBS 0.020193f
C943 VDD1.n120 VSUBS 0.010851f
C944 VDD1.n121 VSUBS 0.011489f
C945 VDD1.n122 VSUBS 0.025648f
C946 VDD1.n123 VSUBS 0.025648f
C947 VDD1.n124 VSUBS 0.011489f
C948 VDD1.n125 VSUBS 0.010851f
C949 VDD1.n126 VSUBS 0.020193f
C950 VDD1.n127 VSUBS 0.020193f
C951 VDD1.n128 VSUBS 0.010851f
C952 VDD1.n129 VSUBS 0.011489f
C953 VDD1.n130 VSUBS 0.025648f
C954 VDD1.n131 VSUBS 0.025648f
C955 VDD1.n132 VSUBS 0.011489f
C956 VDD1.n133 VSUBS 0.010851f
C957 VDD1.n134 VSUBS 0.020193f
C958 VDD1.n135 VSUBS 0.020193f
C959 VDD1.n136 VSUBS 0.010851f
C960 VDD1.n137 VSUBS 0.011489f
C961 VDD1.n138 VSUBS 0.025648f
C962 VDD1.n139 VSUBS 0.025648f
C963 VDD1.n140 VSUBS 0.011489f
C964 VDD1.n141 VSUBS 0.010851f
C965 VDD1.n142 VSUBS 0.020193f
C966 VDD1.n143 VSUBS 0.020193f
C967 VDD1.n144 VSUBS 0.010851f
C968 VDD1.n145 VSUBS 0.011489f
C969 VDD1.n146 VSUBS 0.025648f
C970 VDD1.n147 VSUBS 0.025648f
C971 VDD1.n148 VSUBS 0.025648f
C972 VDD1.n149 VSUBS 0.011489f
C973 VDD1.n150 VSUBS 0.010851f
C974 VDD1.n151 VSUBS 0.020193f
C975 VDD1.n152 VSUBS 0.020193f
C976 VDD1.n153 VSUBS 0.010851f
C977 VDD1.n154 VSUBS 0.01117f
C978 VDD1.n155 VSUBS 0.01117f
C979 VDD1.n156 VSUBS 0.025648f
C980 VDD1.n157 VSUBS 0.057429f
C981 VDD1.n158 VSUBS 0.011489f
C982 VDD1.n159 VSUBS 0.010851f
C983 VDD1.n160 VSUBS 0.048055f
C984 VDD1.n161 VSUBS 0.656561f
C985 VTAIL.n0 VSUBS 0.029183f
C986 VTAIL.n1 VSUBS 0.028305f
C987 VTAIL.n2 VSUBS 0.01521f
C988 VTAIL.n3 VSUBS 0.035951f
C989 VTAIL.n4 VSUBS 0.016105f
C990 VTAIL.n5 VSUBS 0.028305f
C991 VTAIL.n6 VSUBS 0.01521f
C992 VTAIL.n7 VSUBS 0.035951f
C993 VTAIL.n8 VSUBS 0.016105f
C994 VTAIL.n9 VSUBS 0.028305f
C995 VTAIL.n10 VSUBS 0.01521f
C996 VTAIL.n11 VSUBS 0.035951f
C997 VTAIL.n12 VSUBS 0.016105f
C998 VTAIL.n13 VSUBS 0.028305f
C999 VTAIL.n14 VSUBS 0.01521f
C1000 VTAIL.n15 VSUBS 0.035951f
C1001 VTAIL.n16 VSUBS 0.016105f
C1002 VTAIL.n17 VSUBS 0.028305f
C1003 VTAIL.n18 VSUBS 0.01521f
C1004 VTAIL.n19 VSUBS 0.035951f
C1005 VTAIL.n20 VSUBS 0.016105f
C1006 VTAIL.n21 VSUBS 0.028305f
C1007 VTAIL.n22 VSUBS 0.01521f
C1008 VTAIL.n23 VSUBS 0.035951f
C1009 VTAIL.n24 VSUBS 0.016105f
C1010 VTAIL.n25 VSUBS 0.196938f
C1011 VTAIL.t3 VSUBS 0.076941f
C1012 VTAIL.n26 VSUBS 0.026963f
C1013 VTAIL.n27 VSUBS 0.02287f
C1014 VTAIL.n28 VSUBS 0.01521f
C1015 VTAIL.n29 VSUBS 1.7675f
C1016 VTAIL.n30 VSUBS 0.028305f
C1017 VTAIL.n31 VSUBS 0.01521f
C1018 VTAIL.n32 VSUBS 0.016105f
C1019 VTAIL.n33 VSUBS 0.035951f
C1020 VTAIL.n34 VSUBS 0.035951f
C1021 VTAIL.n35 VSUBS 0.016105f
C1022 VTAIL.n36 VSUBS 0.01521f
C1023 VTAIL.n37 VSUBS 0.028305f
C1024 VTAIL.n38 VSUBS 0.028305f
C1025 VTAIL.n39 VSUBS 0.01521f
C1026 VTAIL.n40 VSUBS 0.016105f
C1027 VTAIL.n41 VSUBS 0.035951f
C1028 VTAIL.n42 VSUBS 0.035951f
C1029 VTAIL.n43 VSUBS 0.016105f
C1030 VTAIL.n44 VSUBS 0.01521f
C1031 VTAIL.n45 VSUBS 0.028305f
C1032 VTAIL.n46 VSUBS 0.028305f
C1033 VTAIL.n47 VSUBS 0.01521f
C1034 VTAIL.n48 VSUBS 0.016105f
C1035 VTAIL.n49 VSUBS 0.035951f
C1036 VTAIL.n50 VSUBS 0.035951f
C1037 VTAIL.n51 VSUBS 0.016105f
C1038 VTAIL.n52 VSUBS 0.01521f
C1039 VTAIL.n53 VSUBS 0.028305f
C1040 VTAIL.n54 VSUBS 0.028305f
C1041 VTAIL.n55 VSUBS 0.01521f
C1042 VTAIL.n56 VSUBS 0.016105f
C1043 VTAIL.n57 VSUBS 0.035951f
C1044 VTAIL.n58 VSUBS 0.035951f
C1045 VTAIL.n59 VSUBS 0.016105f
C1046 VTAIL.n60 VSUBS 0.01521f
C1047 VTAIL.n61 VSUBS 0.028305f
C1048 VTAIL.n62 VSUBS 0.028305f
C1049 VTAIL.n63 VSUBS 0.01521f
C1050 VTAIL.n64 VSUBS 0.016105f
C1051 VTAIL.n65 VSUBS 0.035951f
C1052 VTAIL.n66 VSUBS 0.035951f
C1053 VTAIL.n67 VSUBS 0.035951f
C1054 VTAIL.n68 VSUBS 0.016105f
C1055 VTAIL.n69 VSUBS 0.01521f
C1056 VTAIL.n70 VSUBS 0.028305f
C1057 VTAIL.n71 VSUBS 0.028305f
C1058 VTAIL.n72 VSUBS 0.01521f
C1059 VTAIL.n73 VSUBS 0.015657f
C1060 VTAIL.n74 VSUBS 0.015657f
C1061 VTAIL.n75 VSUBS 0.035951f
C1062 VTAIL.n76 VSUBS 0.080499f
C1063 VTAIL.n77 VSUBS 0.016105f
C1064 VTAIL.n78 VSUBS 0.01521f
C1065 VTAIL.n79 VSUBS 0.067359f
C1066 VTAIL.n80 VSUBS 0.040251f
C1067 VTAIL.n81 VSUBS 1.9915f
C1068 VTAIL.n82 VSUBS 0.029183f
C1069 VTAIL.n83 VSUBS 0.028305f
C1070 VTAIL.n84 VSUBS 0.01521f
C1071 VTAIL.n85 VSUBS 0.035951f
C1072 VTAIL.n86 VSUBS 0.016105f
C1073 VTAIL.n87 VSUBS 0.028305f
C1074 VTAIL.n88 VSUBS 0.01521f
C1075 VTAIL.n89 VSUBS 0.035951f
C1076 VTAIL.n90 VSUBS 0.035951f
C1077 VTAIL.n91 VSUBS 0.016105f
C1078 VTAIL.n92 VSUBS 0.028305f
C1079 VTAIL.n93 VSUBS 0.01521f
C1080 VTAIL.n94 VSUBS 0.035951f
C1081 VTAIL.n95 VSUBS 0.016105f
C1082 VTAIL.n96 VSUBS 0.028305f
C1083 VTAIL.n97 VSUBS 0.01521f
C1084 VTAIL.n98 VSUBS 0.035951f
C1085 VTAIL.n99 VSUBS 0.016105f
C1086 VTAIL.n100 VSUBS 0.028305f
C1087 VTAIL.n101 VSUBS 0.01521f
C1088 VTAIL.n102 VSUBS 0.035951f
C1089 VTAIL.n103 VSUBS 0.016105f
C1090 VTAIL.n104 VSUBS 0.028305f
C1091 VTAIL.n105 VSUBS 0.01521f
C1092 VTAIL.n106 VSUBS 0.035951f
C1093 VTAIL.n107 VSUBS 0.016105f
C1094 VTAIL.n108 VSUBS 0.196938f
C1095 VTAIL.t1 VSUBS 0.076941f
C1096 VTAIL.n109 VSUBS 0.026963f
C1097 VTAIL.n110 VSUBS 0.02287f
C1098 VTAIL.n111 VSUBS 0.01521f
C1099 VTAIL.n112 VSUBS 1.7675f
C1100 VTAIL.n113 VSUBS 0.028305f
C1101 VTAIL.n114 VSUBS 0.01521f
C1102 VTAIL.n115 VSUBS 0.016105f
C1103 VTAIL.n116 VSUBS 0.035951f
C1104 VTAIL.n117 VSUBS 0.035951f
C1105 VTAIL.n118 VSUBS 0.016105f
C1106 VTAIL.n119 VSUBS 0.01521f
C1107 VTAIL.n120 VSUBS 0.028305f
C1108 VTAIL.n121 VSUBS 0.028305f
C1109 VTAIL.n122 VSUBS 0.01521f
C1110 VTAIL.n123 VSUBS 0.016105f
C1111 VTAIL.n124 VSUBS 0.035951f
C1112 VTAIL.n125 VSUBS 0.035951f
C1113 VTAIL.n126 VSUBS 0.016105f
C1114 VTAIL.n127 VSUBS 0.01521f
C1115 VTAIL.n128 VSUBS 0.028305f
C1116 VTAIL.n129 VSUBS 0.028305f
C1117 VTAIL.n130 VSUBS 0.01521f
C1118 VTAIL.n131 VSUBS 0.016105f
C1119 VTAIL.n132 VSUBS 0.035951f
C1120 VTAIL.n133 VSUBS 0.035951f
C1121 VTAIL.n134 VSUBS 0.016105f
C1122 VTAIL.n135 VSUBS 0.01521f
C1123 VTAIL.n136 VSUBS 0.028305f
C1124 VTAIL.n137 VSUBS 0.028305f
C1125 VTAIL.n138 VSUBS 0.01521f
C1126 VTAIL.n139 VSUBS 0.016105f
C1127 VTAIL.n140 VSUBS 0.035951f
C1128 VTAIL.n141 VSUBS 0.035951f
C1129 VTAIL.n142 VSUBS 0.016105f
C1130 VTAIL.n143 VSUBS 0.01521f
C1131 VTAIL.n144 VSUBS 0.028305f
C1132 VTAIL.n145 VSUBS 0.028305f
C1133 VTAIL.n146 VSUBS 0.01521f
C1134 VTAIL.n147 VSUBS 0.016105f
C1135 VTAIL.n148 VSUBS 0.035951f
C1136 VTAIL.n149 VSUBS 0.035951f
C1137 VTAIL.n150 VSUBS 0.016105f
C1138 VTAIL.n151 VSUBS 0.01521f
C1139 VTAIL.n152 VSUBS 0.028305f
C1140 VTAIL.n153 VSUBS 0.028305f
C1141 VTAIL.n154 VSUBS 0.01521f
C1142 VTAIL.n155 VSUBS 0.015657f
C1143 VTAIL.n156 VSUBS 0.015657f
C1144 VTAIL.n157 VSUBS 0.035951f
C1145 VTAIL.n158 VSUBS 0.080499f
C1146 VTAIL.n159 VSUBS 0.016105f
C1147 VTAIL.n160 VSUBS 0.01521f
C1148 VTAIL.n161 VSUBS 0.067359f
C1149 VTAIL.n162 VSUBS 0.040251f
C1150 VTAIL.n163 VSUBS 2.02825f
C1151 VTAIL.n164 VSUBS 0.029183f
C1152 VTAIL.n165 VSUBS 0.028305f
C1153 VTAIL.n166 VSUBS 0.01521f
C1154 VTAIL.n167 VSUBS 0.035951f
C1155 VTAIL.n168 VSUBS 0.016105f
C1156 VTAIL.n169 VSUBS 0.028305f
C1157 VTAIL.n170 VSUBS 0.01521f
C1158 VTAIL.n171 VSUBS 0.035951f
C1159 VTAIL.n172 VSUBS 0.035951f
C1160 VTAIL.n173 VSUBS 0.016105f
C1161 VTAIL.n174 VSUBS 0.028305f
C1162 VTAIL.n175 VSUBS 0.01521f
C1163 VTAIL.n176 VSUBS 0.035951f
C1164 VTAIL.n177 VSUBS 0.016105f
C1165 VTAIL.n178 VSUBS 0.028305f
C1166 VTAIL.n179 VSUBS 0.01521f
C1167 VTAIL.n180 VSUBS 0.035951f
C1168 VTAIL.n181 VSUBS 0.016105f
C1169 VTAIL.n182 VSUBS 0.028305f
C1170 VTAIL.n183 VSUBS 0.01521f
C1171 VTAIL.n184 VSUBS 0.035951f
C1172 VTAIL.n185 VSUBS 0.016105f
C1173 VTAIL.n186 VSUBS 0.028305f
C1174 VTAIL.n187 VSUBS 0.01521f
C1175 VTAIL.n188 VSUBS 0.035951f
C1176 VTAIL.n189 VSUBS 0.016105f
C1177 VTAIL.n190 VSUBS 0.196938f
C1178 VTAIL.t2 VSUBS 0.076941f
C1179 VTAIL.n191 VSUBS 0.026963f
C1180 VTAIL.n192 VSUBS 0.02287f
C1181 VTAIL.n193 VSUBS 0.01521f
C1182 VTAIL.n194 VSUBS 1.7675f
C1183 VTAIL.n195 VSUBS 0.028305f
C1184 VTAIL.n196 VSUBS 0.01521f
C1185 VTAIL.n197 VSUBS 0.016105f
C1186 VTAIL.n198 VSUBS 0.035951f
C1187 VTAIL.n199 VSUBS 0.035951f
C1188 VTAIL.n200 VSUBS 0.016105f
C1189 VTAIL.n201 VSUBS 0.01521f
C1190 VTAIL.n202 VSUBS 0.028305f
C1191 VTAIL.n203 VSUBS 0.028305f
C1192 VTAIL.n204 VSUBS 0.01521f
C1193 VTAIL.n205 VSUBS 0.016105f
C1194 VTAIL.n206 VSUBS 0.035951f
C1195 VTAIL.n207 VSUBS 0.035951f
C1196 VTAIL.n208 VSUBS 0.016105f
C1197 VTAIL.n209 VSUBS 0.01521f
C1198 VTAIL.n210 VSUBS 0.028305f
C1199 VTAIL.n211 VSUBS 0.028305f
C1200 VTAIL.n212 VSUBS 0.01521f
C1201 VTAIL.n213 VSUBS 0.016105f
C1202 VTAIL.n214 VSUBS 0.035951f
C1203 VTAIL.n215 VSUBS 0.035951f
C1204 VTAIL.n216 VSUBS 0.016105f
C1205 VTAIL.n217 VSUBS 0.01521f
C1206 VTAIL.n218 VSUBS 0.028305f
C1207 VTAIL.n219 VSUBS 0.028305f
C1208 VTAIL.n220 VSUBS 0.01521f
C1209 VTAIL.n221 VSUBS 0.016105f
C1210 VTAIL.n222 VSUBS 0.035951f
C1211 VTAIL.n223 VSUBS 0.035951f
C1212 VTAIL.n224 VSUBS 0.016105f
C1213 VTAIL.n225 VSUBS 0.01521f
C1214 VTAIL.n226 VSUBS 0.028305f
C1215 VTAIL.n227 VSUBS 0.028305f
C1216 VTAIL.n228 VSUBS 0.01521f
C1217 VTAIL.n229 VSUBS 0.016105f
C1218 VTAIL.n230 VSUBS 0.035951f
C1219 VTAIL.n231 VSUBS 0.035951f
C1220 VTAIL.n232 VSUBS 0.016105f
C1221 VTAIL.n233 VSUBS 0.01521f
C1222 VTAIL.n234 VSUBS 0.028305f
C1223 VTAIL.n235 VSUBS 0.028305f
C1224 VTAIL.n236 VSUBS 0.01521f
C1225 VTAIL.n237 VSUBS 0.015657f
C1226 VTAIL.n238 VSUBS 0.015657f
C1227 VTAIL.n239 VSUBS 0.035951f
C1228 VTAIL.n240 VSUBS 0.080499f
C1229 VTAIL.n241 VSUBS 0.016105f
C1230 VTAIL.n242 VSUBS 0.01521f
C1231 VTAIL.n243 VSUBS 0.067359f
C1232 VTAIL.n244 VSUBS 0.040251f
C1233 VTAIL.n245 VSUBS 1.85999f
C1234 VTAIL.n246 VSUBS 0.029183f
C1235 VTAIL.n247 VSUBS 0.028305f
C1236 VTAIL.n248 VSUBS 0.01521f
C1237 VTAIL.n249 VSUBS 0.035951f
C1238 VTAIL.n250 VSUBS 0.016105f
C1239 VTAIL.n251 VSUBS 0.028305f
C1240 VTAIL.n252 VSUBS 0.01521f
C1241 VTAIL.n253 VSUBS 0.035951f
C1242 VTAIL.n254 VSUBS 0.016105f
C1243 VTAIL.n255 VSUBS 0.028305f
C1244 VTAIL.n256 VSUBS 0.01521f
C1245 VTAIL.n257 VSUBS 0.035951f
C1246 VTAIL.n258 VSUBS 0.016105f
C1247 VTAIL.n259 VSUBS 0.028305f
C1248 VTAIL.n260 VSUBS 0.01521f
C1249 VTAIL.n261 VSUBS 0.035951f
C1250 VTAIL.n262 VSUBS 0.016105f
C1251 VTAIL.n263 VSUBS 0.028305f
C1252 VTAIL.n264 VSUBS 0.01521f
C1253 VTAIL.n265 VSUBS 0.035951f
C1254 VTAIL.n266 VSUBS 0.016105f
C1255 VTAIL.n267 VSUBS 0.028305f
C1256 VTAIL.n268 VSUBS 0.01521f
C1257 VTAIL.n269 VSUBS 0.035951f
C1258 VTAIL.n270 VSUBS 0.016105f
C1259 VTAIL.n271 VSUBS 0.196938f
C1260 VTAIL.t0 VSUBS 0.076941f
C1261 VTAIL.n272 VSUBS 0.026963f
C1262 VTAIL.n273 VSUBS 0.02287f
C1263 VTAIL.n274 VSUBS 0.01521f
C1264 VTAIL.n275 VSUBS 1.7675f
C1265 VTAIL.n276 VSUBS 0.028305f
C1266 VTAIL.n277 VSUBS 0.01521f
C1267 VTAIL.n278 VSUBS 0.016105f
C1268 VTAIL.n279 VSUBS 0.035951f
C1269 VTAIL.n280 VSUBS 0.035951f
C1270 VTAIL.n281 VSUBS 0.016105f
C1271 VTAIL.n282 VSUBS 0.01521f
C1272 VTAIL.n283 VSUBS 0.028305f
C1273 VTAIL.n284 VSUBS 0.028305f
C1274 VTAIL.n285 VSUBS 0.01521f
C1275 VTAIL.n286 VSUBS 0.016105f
C1276 VTAIL.n287 VSUBS 0.035951f
C1277 VTAIL.n288 VSUBS 0.035951f
C1278 VTAIL.n289 VSUBS 0.016105f
C1279 VTAIL.n290 VSUBS 0.01521f
C1280 VTAIL.n291 VSUBS 0.028305f
C1281 VTAIL.n292 VSUBS 0.028305f
C1282 VTAIL.n293 VSUBS 0.01521f
C1283 VTAIL.n294 VSUBS 0.016105f
C1284 VTAIL.n295 VSUBS 0.035951f
C1285 VTAIL.n296 VSUBS 0.035951f
C1286 VTAIL.n297 VSUBS 0.016105f
C1287 VTAIL.n298 VSUBS 0.01521f
C1288 VTAIL.n299 VSUBS 0.028305f
C1289 VTAIL.n300 VSUBS 0.028305f
C1290 VTAIL.n301 VSUBS 0.01521f
C1291 VTAIL.n302 VSUBS 0.016105f
C1292 VTAIL.n303 VSUBS 0.035951f
C1293 VTAIL.n304 VSUBS 0.035951f
C1294 VTAIL.n305 VSUBS 0.016105f
C1295 VTAIL.n306 VSUBS 0.01521f
C1296 VTAIL.n307 VSUBS 0.028305f
C1297 VTAIL.n308 VSUBS 0.028305f
C1298 VTAIL.n309 VSUBS 0.01521f
C1299 VTAIL.n310 VSUBS 0.016105f
C1300 VTAIL.n311 VSUBS 0.035951f
C1301 VTAIL.n312 VSUBS 0.035951f
C1302 VTAIL.n313 VSUBS 0.035951f
C1303 VTAIL.n314 VSUBS 0.016105f
C1304 VTAIL.n315 VSUBS 0.01521f
C1305 VTAIL.n316 VSUBS 0.028305f
C1306 VTAIL.n317 VSUBS 0.028305f
C1307 VTAIL.n318 VSUBS 0.01521f
C1308 VTAIL.n319 VSUBS 0.015657f
C1309 VTAIL.n320 VSUBS 0.015657f
C1310 VTAIL.n321 VSUBS 0.035951f
C1311 VTAIL.n322 VSUBS 0.080499f
C1312 VTAIL.n323 VSUBS 0.016105f
C1313 VTAIL.n324 VSUBS 0.01521f
C1314 VTAIL.n325 VSUBS 0.067359f
C1315 VTAIL.n326 VSUBS 0.040251f
C1316 VTAIL.n327 VSUBS 1.76977f
C1317 VP.t1 VSUBS 4.23675f
C1318 VP.t0 VSUBS 3.73819f
C1319 VP.n0 VSUBS 6.15353f
.ends

