* NGSPICE file created from diff_pair_sample_1204.ext - technology: sky130A

.subckt diff_pair_sample_1204 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=1.1
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=1.1
X2 VDD1.t2 VP.t1 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=1.1
X3 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=1.1
X4 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=1.1
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=1.1
X6 VTAIL.t6 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=1.1
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=1.1
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3761 pd=8.67 as=3.2526 ps=17.46 w=8.34 l=1.1
X9 VTAIL.t5 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=1.1
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=0 ps=0 w=8.34 l=1.1
X11 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2526 pd=17.46 as=1.3761 ps=8.67 w=8.34 l=1.1
R0 VP.n0 VP.t2 237.042
R1 VP.n0 VP.t0 236.953
R2 VP.n2 VP.t3 218.435
R3 VP.n3 VP.t1 218.435
R4 VP.n4 VP.n3 80.6037
R5 VP.n2 VP.n1 80.6037
R6 VP.n1 VP.n0 70.2683
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VTAIL.n5 VTAIL.t6 52.8819
R11 VTAIL.n4 VTAIL.t2 52.8819
R12 VTAIL.n3 VTAIL.t1 52.8819
R13 VTAIL.n7 VTAIL.t3 52.8818
R14 VTAIL.n0 VTAIL.t0 52.8818
R15 VTAIL.n1 VTAIL.t7 52.8818
R16 VTAIL.n2 VTAIL.t5 52.8818
R17 VTAIL.n6 VTAIL.t4 52.8818
R18 VTAIL.n7 VTAIL.n6 20.7893
R19 VTAIL.n3 VTAIL.n2 20.7893
R20 VTAIL.n4 VTAIL.n3 1.23326
R21 VTAIL.n6 VTAIL.n5 1.23326
R22 VTAIL.n2 VTAIL.n1 1.23326
R23 VTAIL VTAIL.n0 0.675069
R24 VTAIL VTAIL.n7 0.55869
R25 VTAIL.n5 VTAIL.n4 0.470328
R26 VTAIL.n1 VTAIL.n0 0.470328
R27 VDD1 VDD1.n1 102.314
R28 VDD1 VDD1.n0 67.2447
R29 VDD1.n0 VDD1.t1 2.3746
R30 VDD1.n0 VDD1.t3 2.3746
R31 VDD1.n1 VDD1.t0 2.3746
R32 VDD1.n1 VDD1.t2 2.3746
R33 B.n531 B.n530 585
R34 B.n532 B.n531 585
R35 B.n219 B.n76 585
R36 B.n218 B.n217 585
R37 B.n216 B.n215 585
R38 B.n214 B.n213 585
R39 B.n212 B.n211 585
R40 B.n210 B.n209 585
R41 B.n208 B.n207 585
R42 B.n206 B.n205 585
R43 B.n204 B.n203 585
R44 B.n202 B.n201 585
R45 B.n200 B.n199 585
R46 B.n198 B.n197 585
R47 B.n196 B.n195 585
R48 B.n194 B.n193 585
R49 B.n192 B.n191 585
R50 B.n190 B.n189 585
R51 B.n188 B.n187 585
R52 B.n186 B.n185 585
R53 B.n184 B.n183 585
R54 B.n182 B.n181 585
R55 B.n180 B.n179 585
R56 B.n178 B.n177 585
R57 B.n176 B.n175 585
R58 B.n174 B.n173 585
R59 B.n172 B.n171 585
R60 B.n170 B.n169 585
R61 B.n168 B.n167 585
R62 B.n166 B.n165 585
R63 B.n164 B.n163 585
R64 B.n162 B.n161 585
R65 B.n160 B.n159 585
R66 B.n158 B.n157 585
R67 B.n156 B.n155 585
R68 B.n154 B.n153 585
R69 B.n152 B.n151 585
R70 B.n150 B.n149 585
R71 B.n148 B.n147 585
R72 B.n146 B.n145 585
R73 B.n144 B.n143 585
R74 B.n141 B.n140 585
R75 B.n139 B.n138 585
R76 B.n137 B.n136 585
R77 B.n135 B.n134 585
R78 B.n133 B.n132 585
R79 B.n131 B.n130 585
R80 B.n129 B.n128 585
R81 B.n127 B.n126 585
R82 B.n125 B.n124 585
R83 B.n123 B.n122 585
R84 B.n121 B.n120 585
R85 B.n119 B.n118 585
R86 B.n117 B.n116 585
R87 B.n115 B.n114 585
R88 B.n113 B.n112 585
R89 B.n111 B.n110 585
R90 B.n109 B.n108 585
R91 B.n107 B.n106 585
R92 B.n105 B.n104 585
R93 B.n103 B.n102 585
R94 B.n101 B.n100 585
R95 B.n99 B.n98 585
R96 B.n97 B.n96 585
R97 B.n95 B.n94 585
R98 B.n93 B.n92 585
R99 B.n91 B.n90 585
R100 B.n89 B.n88 585
R101 B.n87 B.n86 585
R102 B.n85 B.n84 585
R103 B.n83 B.n82 585
R104 B.n39 B.n38 585
R105 B.n529 B.n40 585
R106 B.n533 B.n40 585
R107 B.n528 B.n527 585
R108 B.n527 B.n36 585
R109 B.n526 B.n35 585
R110 B.n539 B.n35 585
R111 B.n525 B.n34 585
R112 B.n540 B.n34 585
R113 B.n524 B.n33 585
R114 B.n541 B.n33 585
R115 B.n523 B.n522 585
R116 B.n522 B.n32 585
R117 B.n521 B.n28 585
R118 B.n547 B.n28 585
R119 B.n520 B.n27 585
R120 B.n548 B.n27 585
R121 B.n519 B.n26 585
R122 B.n549 B.n26 585
R123 B.n518 B.n517 585
R124 B.n517 B.n22 585
R125 B.n516 B.n21 585
R126 B.n555 B.n21 585
R127 B.n515 B.n20 585
R128 B.n556 B.n20 585
R129 B.n514 B.n19 585
R130 B.n557 B.n19 585
R131 B.n513 B.n512 585
R132 B.n512 B.n15 585
R133 B.n511 B.n14 585
R134 B.n563 B.n14 585
R135 B.n510 B.n13 585
R136 B.n564 B.n13 585
R137 B.n509 B.n12 585
R138 B.n565 B.n12 585
R139 B.n508 B.n507 585
R140 B.n507 B.n506 585
R141 B.n505 B.n504 585
R142 B.n505 B.n8 585
R143 B.n503 B.n7 585
R144 B.n572 B.n7 585
R145 B.n502 B.n6 585
R146 B.n573 B.n6 585
R147 B.n501 B.n5 585
R148 B.n574 B.n5 585
R149 B.n500 B.n499 585
R150 B.n499 B.n4 585
R151 B.n498 B.n220 585
R152 B.n498 B.n497 585
R153 B.n488 B.n221 585
R154 B.n222 B.n221 585
R155 B.n490 B.n489 585
R156 B.n491 B.n490 585
R157 B.n487 B.n227 585
R158 B.n227 B.n226 585
R159 B.n486 B.n485 585
R160 B.n485 B.n484 585
R161 B.n229 B.n228 585
R162 B.n230 B.n229 585
R163 B.n477 B.n476 585
R164 B.n478 B.n477 585
R165 B.n475 B.n235 585
R166 B.n235 B.n234 585
R167 B.n474 B.n473 585
R168 B.n473 B.n472 585
R169 B.n237 B.n236 585
R170 B.n238 B.n237 585
R171 B.n465 B.n464 585
R172 B.n466 B.n465 585
R173 B.n463 B.n243 585
R174 B.n243 B.n242 585
R175 B.n462 B.n461 585
R176 B.n461 B.n460 585
R177 B.n245 B.n244 585
R178 B.n453 B.n245 585
R179 B.n452 B.n451 585
R180 B.n454 B.n452 585
R181 B.n450 B.n250 585
R182 B.n250 B.n249 585
R183 B.n449 B.n448 585
R184 B.n448 B.n447 585
R185 B.n252 B.n251 585
R186 B.n253 B.n252 585
R187 B.n440 B.n439 585
R188 B.n441 B.n440 585
R189 B.n256 B.n255 585
R190 B.n297 B.n296 585
R191 B.n298 B.n294 585
R192 B.n294 B.n257 585
R193 B.n300 B.n299 585
R194 B.n302 B.n293 585
R195 B.n305 B.n304 585
R196 B.n306 B.n292 585
R197 B.n308 B.n307 585
R198 B.n310 B.n291 585
R199 B.n313 B.n312 585
R200 B.n314 B.n290 585
R201 B.n316 B.n315 585
R202 B.n318 B.n289 585
R203 B.n321 B.n320 585
R204 B.n322 B.n288 585
R205 B.n324 B.n323 585
R206 B.n326 B.n287 585
R207 B.n329 B.n328 585
R208 B.n330 B.n286 585
R209 B.n332 B.n331 585
R210 B.n334 B.n285 585
R211 B.n337 B.n336 585
R212 B.n338 B.n284 585
R213 B.n340 B.n339 585
R214 B.n342 B.n283 585
R215 B.n345 B.n344 585
R216 B.n346 B.n282 585
R217 B.n348 B.n347 585
R218 B.n350 B.n281 585
R219 B.n353 B.n352 585
R220 B.n354 B.n278 585
R221 B.n357 B.n356 585
R222 B.n359 B.n277 585
R223 B.n362 B.n361 585
R224 B.n363 B.n276 585
R225 B.n365 B.n364 585
R226 B.n367 B.n275 585
R227 B.n370 B.n369 585
R228 B.n371 B.n274 585
R229 B.n376 B.n375 585
R230 B.n378 B.n273 585
R231 B.n381 B.n380 585
R232 B.n382 B.n272 585
R233 B.n384 B.n383 585
R234 B.n386 B.n271 585
R235 B.n389 B.n388 585
R236 B.n390 B.n270 585
R237 B.n392 B.n391 585
R238 B.n394 B.n269 585
R239 B.n397 B.n396 585
R240 B.n398 B.n268 585
R241 B.n400 B.n399 585
R242 B.n402 B.n267 585
R243 B.n405 B.n404 585
R244 B.n406 B.n266 585
R245 B.n408 B.n407 585
R246 B.n410 B.n265 585
R247 B.n413 B.n412 585
R248 B.n414 B.n264 585
R249 B.n416 B.n415 585
R250 B.n418 B.n263 585
R251 B.n421 B.n420 585
R252 B.n422 B.n262 585
R253 B.n424 B.n423 585
R254 B.n426 B.n261 585
R255 B.n429 B.n428 585
R256 B.n430 B.n260 585
R257 B.n432 B.n431 585
R258 B.n434 B.n259 585
R259 B.n437 B.n436 585
R260 B.n438 B.n258 585
R261 B.n443 B.n442 585
R262 B.n442 B.n441 585
R263 B.n444 B.n254 585
R264 B.n254 B.n253 585
R265 B.n446 B.n445 585
R266 B.n447 B.n446 585
R267 B.n248 B.n247 585
R268 B.n249 B.n248 585
R269 B.n456 B.n455 585
R270 B.n455 B.n454 585
R271 B.n457 B.n246 585
R272 B.n453 B.n246 585
R273 B.n459 B.n458 585
R274 B.n460 B.n459 585
R275 B.n241 B.n240 585
R276 B.n242 B.n241 585
R277 B.n468 B.n467 585
R278 B.n467 B.n466 585
R279 B.n469 B.n239 585
R280 B.n239 B.n238 585
R281 B.n471 B.n470 585
R282 B.n472 B.n471 585
R283 B.n233 B.n232 585
R284 B.n234 B.n233 585
R285 B.n480 B.n479 585
R286 B.n479 B.n478 585
R287 B.n481 B.n231 585
R288 B.n231 B.n230 585
R289 B.n483 B.n482 585
R290 B.n484 B.n483 585
R291 B.n225 B.n224 585
R292 B.n226 B.n225 585
R293 B.n493 B.n492 585
R294 B.n492 B.n491 585
R295 B.n494 B.n223 585
R296 B.n223 B.n222 585
R297 B.n496 B.n495 585
R298 B.n497 B.n496 585
R299 B.n3 B.n0 585
R300 B.n4 B.n3 585
R301 B.n571 B.n1 585
R302 B.n572 B.n571 585
R303 B.n570 B.n569 585
R304 B.n570 B.n8 585
R305 B.n568 B.n9 585
R306 B.n506 B.n9 585
R307 B.n567 B.n566 585
R308 B.n566 B.n565 585
R309 B.n11 B.n10 585
R310 B.n564 B.n11 585
R311 B.n562 B.n561 585
R312 B.n563 B.n562 585
R313 B.n560 B.n16 585
R314 B.n16 B.n15 585
R315 B.n559 B.n558 585
R316 B.n558 B.n557 585
R317 B.n18 B.n17 585
R318 B.n556 B.n18 585
R319 B.n554 B.n553 585
R320 B.n555 B.n554 585
R321 B.n552 B.n23 585
R322 B.n23 B.n22 585
R323 B.n551 B.n550 585
R324 B.n550 B.n549 585
R325 B.n25 B.n24 585
R326 B.n548 B.n25 585
R327 B.n546 B.n545 585
R328 B.n547 B.n546 585
R329 B.n544 B.n29 585
R330 B.n32 B.n29 585
R331 B.n543 B.n542 585
R332 B.n542 B.n541 585
R333 B.n31 B.n30 585
R334 B.n540 B.n31 585
R335 B.n538 B.n537 585
R336 B.n539 B.n538 585
R337 B.n536 B.n37 585
R338 B.n37 B.n36 585
R339 B.n535 B.n534 585
R340 B.n534 B.n533 585
R341 B.n575 B.n574 585
R342 B.n573 B.n2 585
R343 B.n534 B.n39 559.769
R344 B.n531 B.n40 559.769
R345 B.n440 B.n258 559.769
R346 B.n442 B.n256 559.769
R347 B.n80 B.t15 386.283
R348 B.n77 B.t11 386.283
R349 B.n372 B.t4 386.283
R350 B.n279 B.t8 386.283
R351 B.n532 B.n75 256.663
R352 B.n532 B.n74 256.663
R353 B.n532 B.n73 256.663
R354 B.n532 B.n72 256.663
R355 B.n532 B.n71 256.663
R356 B.n532 B.n70 256.663
R357 B.n532 B.n69 256.663
R358 B.n532 B.n68 256.663
R359 B.n532 B.n67 256.663
R360 B.n532 B.n66 256.663
R361 B.n532 B.n65 256.663
R362 B.n532 B.n64 256.663
R363 B.n532 B.n63 256.663
R364 B.n532 B.n62 256.663
R365 B.n532 B.n61 256.663
R366 B.n532 B.n60 256.663
R367 B.n532 B.n59 256.663
R368 B.n532 B.n58 256.663
R369 B.n532 B.n57 256.663
R370 B.n532 B.n56 256.663
R371 B.n532 B.n55 256.663
R372 B.n532 B.n54 256.663
R373 B.n532 B.n53 256.663
R374 B.n532 B.n52 256.663
R375 B.n532 B.n51 256.663
R376 B.n532 B.n50 256.663
R377 B.n532 B.n49 256.663
R378 B.n532 B.n48 256.663
R379 B.n532 B.n47 256.663
R380 B.n532 B.n46 256.663
R381 B.n532 B.n45 256.663
R382 B.n532 B.n44 256.663
R383 B.n532 B.n43 256.663
R384 B.n532 B.n42 256.663
R385 B.n532 B.n41 256.663
R386 B.n295 B.n257 256.663
R387 B.n301 B.n257 256.663
R388 B.n303 B.n257 256.663
R389 B.n309 B.n257 256.663
R390 B.n311 B.n257 256.663
R391 B.n317 B.n257 256.663
R392 B.n319 B.n257 256.663
R393 B.n325 B.n257 256.663
R394 B.n327 B.n257 256.663
R395 B.n333 B.n257 256.663
R396 B.n335 B.n257 256.663
R397 B.n341 B.n257 256.663
R398 B.n343 B.n257 256.663
R399 B.n349 B.n257 256.663
R400 B.n351 B.n257 256.663
R401 B.n358 B.n257 256.663
R402 B.n360 B.n257 256.663
R403 B.n366 B.n257 256.663
R404 B.n368 B.n257 256.663
R405 B.n377 B.n257 256.663
R406 B.n379 B.n257 256.663
R407 B.n385 B.n257 256.663
R408 B.n387 B.n257 256.663
R409 B.n393 B.n257 256.663
R410 B.n395 B.n257 256.663
R411 B.n401 B.n257 256.663
R412 B.n403 B.n257 256.663
R413 B.n409 B.n257 256.663
R414 B.n411 B.n257 256.663
R415 B.n417 B.n257 256.663
R416 B.n419 B.n257 256.663
R417 B.n425 B.n257 256.663
R418 B.n427 B.n257 256.663
R419 B.n433 B.n257 256.663
R420 B.n435 B.n257 256.663
R421 B.n577 B.n576 256.663
R422 B.n84 B.n83 163.367
R423 B.n88 B.n87 163.367
R424 B.n92 B.n91 163.367
R425 B.n96 B.n95 163.367
R426 B.n100 B.n99 163.367
R427 B.n104 B.n103 163.367
R428 B.n108 B.n107 163.367
R429 B.n112 B.n111 163.367
R430 B.n116 B.n115 163.367
R431 B.n120 B.n119 163.367
R432 B.n124 B.n123 163.367
R433 B.n128 B.n127 163.367
R434 B.n132 B.n131 163.367
R435 B.n136 B.n135 163.367
R436 B.n140 B.n139 163.367
R437 B.n145 B.n144 163.367
R438 B.n149 B.n148 163.367
R439 B.n153 B.n152 163.367
R440 B.n157 B.n156 163.367
R441 B.n161 B.n160 163.367
R442 B.n165 B.n164 163.367
R443 B.n169 B.n168 163.367
R444 B.n173 B.n172 163.367
R445 B.n177 B.n176 163.367
R446 B.n181 B.n180 163.367
R447 B.n185 B.n184 163.367
R448 B.n189 B.n188 163.367
R449 B.n193 B.n192 163.367
R450 B.n197 B.n196 163.367
R451 B.n201 B.n200 163.367
R452 B.n205 B.n204 163.367
R453 B.n209 B.n208 163.367
R454 B.n213 B.n212 163.367
R455 B.n217 B.n216 163.367
R456 B.n531 B.n76 163.367
R457 B.n440 B.n252 163.367
R458 B.n448 B.n252 163.367
R459 B.n448 B.n250 163.367
R460 B.n452 B.n250 163.367
R461 B.n452 B.n245 163.367
R462 B.n461 B.n245 163.367
R463 B.n461 B.n243 163.367
R464 B.n465 B.n243 163.367
R465 B.n465 B.n237 163.367
R466 B.n473 B.n237 163.367
R467 B.n473 B.n235 163.367
R468 B.n477 B.n235 163.367
R469 B.n477 B.n229 163.367
R470 B.n485 B.n229 163.367
R471 B.n485 B.n227 163.367
R472 B.n490 B.n227 163.367
R473 B.n490 B.n221 163.367
R474 B.n498 B.n221 163.367
R475 B.n499 B.n498 163.367
R476 B.n499 B.n5 163.367
R477 B.n6 B.n5 163.367
R478 B.n7 B.n6 163.367
R479 B.n505 B.n7 163.367
R480 B.n507 B.n505 163.367
R481 B.n507 B.n12 163.367
R482 B.n13 B.n12 163.367
R483 B.n14 B.n13 163.367
R484 B.n512 B.n14 163.367
R485 B.n512 B.n19 163.367
R486 B.n20 B.n19 163.367
R487 B.n21 B.n20 163.367
R488 B.n517 B.n21 163.367
R489 B.n517 B.n26 163.367
R490 B.n27 B.n26 163.367
R491 B.n28 B.n27 163.367
R492 B.n522 B.n28 163.367
R493 B.n522 B.n33 163.367
R494 B.n34 B.n33 163.367
R495 B.n35 B.n34 163.367
R496 B.n527 B.n35 163.367
R497 B.n527 B.n40 163.367
R498 B.n296 B.n294 163.367
R499 B.n300 B.n294 163.367
R500 B.n304 B.n302 163.367
R501 B.n308 B.n292 163.367
R502 B.n312 B.n310 163.367
R503 B.n316 B.n290 163.367
R504 B.n320 B.n318 163.367
R505 B.n324 B.n288 163.367
R506 B.n328 B.n326 163.367
R507 B.n332 B.n286 163.367
R508 B.n336 B.n334 163.367
R509 B.n340 B.n284 163.367
R510 B.n344 B.n342 163.367
R511 B.n348 B.n282 163.367
R512 B.n352 B.n350 163.367
R513 B.n357 B.n278 163.367
R514 B.n361 B.n359 163.367
R515 B.n365 B.n276 163.367
R516 B.n369 B.n367 163.367
R517 B.n376 B.n274 163.367
R518 B.n380 B.n378 163.367
R519 B.n384 B.n272 163.367
R520 B.n388 B.n386 163.367
R521 B.n392 B.n270 163.367
R522 B.n396 B.n394 163.367
R523 B.n400 B.n268 163.367
R524 B.n404 B.n402 163.367
R525 B.n408 B.n266 163.367
R526 B.n412 B.n410 163.367
R527 B.n416 B.n264 163.367
R528 B.n420 B.n418 163.367
R529 B.n424 B.n262 163.367
R530 B.n428 B.n426 163.367
R531 B.n432 B.n260 163.367
R532 B.n436 B.n434 163.367
R533 B.n442 B.n254 163.367
R534 B.n446 B.n254 163.367
R535 B.n446 B.n248 163.367
R536 B.n455 B.n248 163.367
R537 B.n455 B.n246 163.367
R538 B.n459 B.n246 163.367
R539 B.n459 B.n241 163.367
R540 B.n467 B.n241 163.367
R541 B.n467 B.n239 163.367
R542 B.n471 B.n239 163.367
R543 B.n471 B.n233 163.367
R544 B.n479 B.n233 163.367
R545 B.n479 B.n231 163.367
R546 B.n483 B.n231 163.367
R547 B.n483 B.n225 163.367
R548 B.n492 B.n225 163.367
R549 B.n492 B.n223 163.367
R550 B.n496 B.n223 163.367
R551 B.n496 B.n3 163.367
R552 B.n575 B.n3 163.367
R553 B.n571 B.n2 163.367
R554 B.n571 B.n570 163.367
R555 B.n570 B.n9 163.367
R556 B.n566 B.n9 163.367
R557 B.n566 B.n11 163.367
R558 B.n562 B.n11 163.367
R559 B.n562 B.n16 163.367
R560 B.n558 B.n16 163.367
R561 B.n558 B.n18 163.367
R562 B.n554 B.n18 163.367
R563 B.n554 B.n23 163.367
R564 B.n550 B.n23 163.367
R565 B.n550 B.n25 163.367
R566 B.n546 B.n25 163.367
R567 B.n546 B.n29 163.367
R568 B.n542 B.n29 163.367
R569 B.n542 B.n31 163.367
R570 B.n538 B.n31 163.367
R571 B.n538 B.n37 163.367
R572 B.n534 B.n37 163.367
R573 B.n441 B.n257 112.303
R574 B.n533 B.n532 112.303
R575 B.n77 B.t13 99.7332
R576 B.n372 B.t7 99.7332
R577 B.n80 B.t16 99.7235
R578 B.n279 B.t10 99.7235
R579 B.n78 B.t14 71.9999
R580 B.n373 B.t6 71.9999
R581 B.n81 B.t17 71.9901
R582 B.n280 B.t9 71.9901
R583 B.n41 B.n39 71.676
R584 B.n84 B.n42 71.676
R585 B.n88 B.n43 71.676
R586 B.n92 B.n44 71.676
R587 B.n96 B.n45 71.676
R588 B.n100 B.n46 71.676
R589 B.n104 B.n47 71.676
R590 B.n108 B.n48 71.676
R591 B.n112 B.n49 71.676
R592 B.n116 B.n50 71.676
R593 B.n120 B.n51 71.676
R594 B.n124 B.n52 71.676
R595 B.n128 B.n53 71.676
R596 B.n132 B.n54 71.676
R597 B.n136 B.n55 71.676
R598 B.n140 B.n56 71.676
R599 B.n145 B.n57 71.676
R600 B.n149 B.n58 71.676
R601 B.n153 B.n59 71.676
R602 B.n157 B.n60 71.676
R603 B.n161 B.n61 71.676
R604 B.n165 B.n62 71.676
R605 B.n169 B.n63 71.676
R606 B.n173 B.n64 71.676
R607 B.n177 B.n65 71.676
R608 B.n181 B.n66 71.676
R609 B.n185 B.n67 71.676
R610 B.n189 B.n68 71.676
R611 B.n193 B.n69 71.676
R612 B.n197 B.n70 71.676
R613 B.n201 B.n71 71.676
R614 B.n205 B.n72 71.676
R615 B.n209 B.n73 71.676
R616 B.n213 B.n74 71.676
R617 B.n217 B.n75 71.676
R618 B.n76 B.n75 71.676
R619 B.n216 B.n74 71.676
R620 B.n212 B.n73 71.676
R621 B.n208 B.n72 71.676
R622 B.n204 B.n71 71.676
R623 B.n200 B.n70 71.676
R624 B.n196 B.n69 71.676
R625 B.n192 B.n68 71.676
R626 B.n188 B.n67 71.676
R627 B.n184 B.n66 71.676
R628 B.n180 B.n65 71.676
R629 B.n176 B.n64 71.676
R630 B.n172 B.n63 71.676
R631 B.n168 B.n62 71.676
R632 B.n164 B.n61 71.676
R633 B.n160 B.n60 71.676
R634 B.n156 B.n59 71.676
R635 B.n152 B.n58 71.676
R636 B.n148 B.n57 71.676
R637 B.n144 B.n56 71.676
R638 B.n139 B.n55 71.676
R639 B.n135 B.n54 71.676
R640 B.n131 B.n53 71.676
R641 B.n127 B.n52 71.676
R642 B.n123 B.n51 71.676
R643 B.n119 B.n50 71.676
R644 B.n115 B.n49 71.676
R645 B.n111 B.n48 71.676
R646 B.n107 B.n47 71.676
R647 B.n103 B.n46 71.676
R648 B.n99 B.n45 71.676
R649 B.n95 B.n44 71.676
R650 B.n91 B.n43 71.676
R651 B.n87 B.n42 71.676
R652 B.n83 B.n41 71.676
R653 B.n295 B.n256 71.676
R654 B.n301 B.n300 71.676
R655 B.n304 B.n303 71.676
R656 B.n309 B.n308 71.676
R657 B.n312 B.n311 71.676
R658 B.n317 B.n316 71.676
R659 B.n320 B.n319 71.676
R660 B.n325 B.n324 71.676
R661 B.n328 B.n327 71.676
R662 B.n333 B.n332 71.676
R663 B.n336 B.n335 71.676
R664 B.n341 B.n340 71.676
R665 B.n344 B.n343 71.676
R666 B.n349 B.n348 71.676
R667 B.n352 B.n351 71.676
R668 B.n358 B.n357 71.676
R669 B.n361 B.n360 71.676
R670 B.n366 B.n365 71.676
R671 B.n369 B.n368 71.676
R672 B.n377 B.n376 71.676
R673 B.n380 B.n379 71.676
R674 B.n385 B.n384 71.676
R675 B.n388 B.n387 71.676
R676 B.n393 B.n392 71.676
R677 B.n396 B.n395 71.676
R678 B.n401 B.n400 71.676
R679 B.n404 B.n403 71.676
R680 B.n409 B.n408 71.676
R681 B.n412 B.n411 71.676
R682 B.n417 B.n416 71.676
R683 B.n420 B.n419 71.676
R684 B.n425 B.n424 71.676
R685 B.n428 B.n427 71.676
R686 B.n433 B.n432 71.676
R687 B.n436 B.n435 71.676
R688 B.n296 B.n295 71.676
R689 B.n302 B.n301 71.676
R690 B.n303 B.n292 71.676
R691 B.n310 B.n309 71.676
R692 B.n311 B.n290 71.676
R693 B.n318 B.n317 71.676
R694 B.n319 B.n288 71.676
R695 B.n326 B.n325 71.676
R696 B.n327 B.n286 71.676
R697 B.n334 B.n333 71.676
R698 B.n335 B.n284 71.676
R699 B.n342 B.n341 71.676
R700 B.n343 B.n282 71.676
R701 B.n350 B.n349 71.676
R702 B.n351 B.n278 71.676
R703 B.n359 B.n358 71.676
R704 B.n360 B.n276 71.676
R705 B.n367 B.n366 71.676
R706 B.n368 B.n274 71.676
R707 B.n378 B.n377 71.676
R708 B.n379 B.n272 71.676
R709 B.n386 B.n385 71.676
R710 B.n387 B.n270 71.676
R711 B.n394 B.n393 71.676
R712 B.n395 B.n268 71.676
R713 B.n402 B.n401 71.676
R714 B.n403 B.n266 71.676
R715 B.n410 B.n409 71.676
R716 B.n411 B.n264 71.676
R717 B.n418 B.n417 71.676
R718 B.n419 B.n262 71.676
R719 B.n426 B.n425 71.676
R720 B.n427 B.n260 71.676
R721 B.n434 B.n433 71.676
R722 B.n435 B.n258 71.676
R723 B.n576 B.n575 71.676
R724 B.n576 B.n2 71.676
R725 B.n142 B.n81 59.5399
R726 B.n79 B.n78 59.5399
R727 B.n374 B.n373 59.5399
R728 B.n355 B.n280 59.5399
R729 B.n441 B.n253 54.9399
R730 B.n447 B.n253 54.9399
R731 B.n447 B.n249 54.9399
R732 B.n454 B.n249 54.9399
R733 B.n454 B.n453 54.9399
R734 B.n460 B.n242 54.9399
R735 B.n466 B.n242 54.9399
R736 B.n466 B.n238 54.9399
R737 B.n472 B.n238 54.9399
R738 B.n472 B.n234 54.9399
R739 B.n478 B.n234 54.9399
R740 B.n484 B.n230 54.9399
R741 B.n484 B.n226 54.9399
R742 B.n491 B.n226 54.9399
R743 B.n497 B.n222 54.9399
R744 B.n497 B.n4 54.9399
R745 B.n574 B.n4 54.9399
R746 B.n574 B.n573 54.9399
R747 B.n573 B.n572 54.9399
R748 B.n572 B.n8 54.9399
R749 B.n506 B.n8 54.9399
R750 B.n565 B.n564 54.9399
R751 B.n564 B.n563 54.9399
R752 B.n563 B.n15 54.9399
R753 B.n557 B.n556 54.9399
R754 B.n556 B.n555 54.9399
R755 B.n555 B.n22 54.9399
R756 B.n549 B.n22 54.9399
R757 B.n549 B.n548 54.9399
R758 B.n548 B.n547 54.9399
R759 B.n541 B.n32 54.9399
R760 B.n541 B.n540 54.9399
R761 B.n540 B.n539 54.9399
R762 B.n539 B.n36 54.9399
R763 B.n533 B.n36 54.9399
R764 B.n460 B.t5 45.2447
R765 B.n547 B.t12 45.2447
R766 B.n491 B.t2 43.6289
R767 B.n565 B.t0 43.6289
R768 B.n443 B.n255 36.3712
R769 B.n439 B.n438 36.3712
R770 B.n530 B.n529 36.3712
R771 B.n535 B.n38 36.3712
R772 B.n478 B.t1 32.3178
R773 B.n557 B.t3 32.3178
R774 B.n81 B.n80 27.7338
R775 B.n78 B.n77 27.7338
R776 B.n373 B.n372 27.7338
R777 B.n280 B.n279 27.7338
R778 B.t1 B.n230 22.6226
R779 B.t3 B.n15 22.6226
R780 B B.n577 18.0485
R781 B.t2 B.n222 11.3116
R782 B.n506 B.t0 11.3116
R783 B.n444 B.n443 10.6151
R784 B.n445 B.n444 10.6151
R785 B.n445 B.n247 10.6151
R786 B.n456 B.n247 10.6151
R787 B.n457 B.n456 10.6151
R788 B.n458 B.n457 10.6151
R789 B.n458 B.n240 10.6151
R790 B.n468 B.n240 10.6151
R791 B.n469 B.n468 10.6151
R792 B.n470 B.n469 10.6151
R793 B.n470 B.n232 10.6151
R794 B.n480 B.n232 10.6151
R795 B.n481 B.n480 10.6151
R796 B.n482 B.n481 10.6151
R797 B.n482 B.n224 10.6151
R798 B.n493 B.n224 10.6151
R799 B.n494 B.n493 10.6151
R800 B.n495 B.n494 10.6151
R801 B.n495 B.n0 10.6151
R802 B.n297 B.n255 10.6151
R803 B.n298 B.n297 10.6151
R804 B.n299 B.n298 10.6151
R805 B.n299 B.n293 10.6151
R806 B.n305 B.n293 10.6151
R807 B.n306 B.n305 10.6151
R808 B.n307 B.n306 10.6151
R809 B.n307 B.n291 10.6151
R810 B.n313 B.n291 10.6151
R811 B.n314 B.n313 10.6151
R812 B.n315 B.n314 10.6151
R813 B.n315 B.n289 10.6151
R814 B.n321 B.n289 10.6151
R815 B.n322 B.n321 10.6151
R816 B.n323 B.n322 10.6151
R817 B.n323 B.n287 10.6151
R818 B.n329 B.n287 10.6151
R819 B.n330 B.n329 10.6151
R820 B.n331 B.n330 10.6151
R821 B.n331 B.n285 10.6151
R822 B.n337 B.n285 10.6151
R823 B.n338 B.n337 10.6151
R824 B.n339 B.n338 10.6151
R825 B.n339 B.n283 10.6151
R826 B.n345 B.n283 10.6151
R827 B.n346 B.n345 10.6151
R828 B.n347 B.n346 10.6151
R829 B.n347 B.n281 10.6151
R830 B.n353 B.n281 10.6151
R831 B.n354 B.n353 10.6151
R832 B.n356 B.n277 10.6151
R833 B.n362 B.n277 10.6151
R834 B.n363 B.n362 10.6151
R835 B.n364 B.n363 10.6151
R836 B.n364 B.n275 10.6151
R837 B.n370 B.n275 10.6151
R838 B.n371 B.n370 10.6151
R839 B.n375 B.n371 10.6151
R840 B.n381 B.n273 10.6151
R841 B.n382 B.n381 10.6151
R842 B.n383 B.n382 10.6151
R843 B.n383 B.n271 10.6151
R844 B.n389 B.n271 10.6151
R845 B.n390 B.n389 10.6151
R846 B.n391 B.n390 10.6151
R847 B.n391 B.n269 10.6151
R848 B.n397 B.n269 10.6151
R849 B.n398 B.n397 10.6151
R850 B.n399 B.n398 10.6151
R851 B.n399 B.n267 10.6151
R852 B.n405 B.n267 10.6151
R853 B.n406 B.n405 10.6151
R854 B.n407 B.n406 10.6151
R855 B.n407 B.n265 10.6151
R856 B.n413 B.n265 10.6151
R857 B.n414 B.n413 10.6151
R858 B.n415 B.n414 10.6151
R859 B.n415 B.n263 10.6151
R860 B.n421 B.n263 10.6151
R861 B.n422 B.n421 10.6151
R862 B.n423 B.n422 10.6151
R863 B.n423 B.n261 10.6151
R864 B.n429 B.n261 10.6151
R865 B.n430 B.n429 10.6151
R866 B.n431 B.n430 10.6151
R867 B.n431 B.n259 10.6151
R868 B.n437 B.n259 10.6151
R869 B.n438 B.n437 10.6151
R870 B.n439 B.n251 10.6151
R871 B.n449 B.n251 10.6151
R872 B.n450 B.n449 10.6151
R873 B.n451 B.n450 10.6151
R874 B.n451 B.n244 10.6151
R875 B.n462 B.n244 10.6151
R876 B.n463 B.n462 10.6151
R877 B.n464 B.n463 10.6151
R878 B.n464 B.n236 10.6151
R879 B.n474 B.n236 10.6151
R880 B.n475 B.n474 10.6151
R881 B.n476 B.n475 10.6151
R882 B.n476 B.n228 10.6151
R883 B.n486 B.n228 10.6151
R884 B.n487 B.n486 10.6151
R885 B.n489 B.n487 10.6151
R886 B.n489 B.n488 10.6151
R887 B.n488 B.n220 10.6151
R888 B.n500 B.n220 10.6151
R889 B.n501 B.n500 10.6151
R890 B.n502 B.n501 10.6151
R891 B.n503 B.n502 10.6151
R892 B.n504 B.n503 10.6151
R893 B.n508 B.n504 10.6151
R894 B.n509 B.n508 10.6151
R895 B.n510 B.n509 10.6151
R896 B.n511 B.n510 10.6151
R897 B.n513 B.n511 10.6151
R898 B.n514 B.n513 10.6151
R899 B.n515 B.n514 10.6151
R900 B.n516 B.n515 10.6151
R901 B.n518 B.n516 10.6151
R902 B.n519 B.n518 10.6151
R903 B.n520 B.n519 10.6151
R904 B.n521 B.n520 10.6151
R905 B.n523 B.n521 10.6151
R906 B.n524 B.n523 10.6151
R907 B.n525 B.n524 10.6151
R908 B.n526 B.n525 10.6151
R909 B.n528 B.n526 10.6151
R910 B.n529 B.n528 10.6151
R911 B.n569 B.n1 10.6151
R912 B.n569 B.n568 10.6151
R913 B.n568 B.n567 10.6151
R914 B.n567 B.n10 10.6151
R915 B.n561 B.n10 10.6151
R916 B.n561 B.n560 10.6151
R917 B.n560 B.n559 10.6151
R918 B.n559 B.n17 10.6151
R919 B.n553 B.n17 10.6151
R920 B.n553 B.n552 10.6151
R921 B.n552 B.n551 10.6151
R922 B.n551 B.n24 10.6151
R923 B.n545 B.n24 10.6151
R924 B.n545 B.n544 10.6151
R925 B.n544 B.n543 10.6151
R926 B.n543 B.n30 10.6151
R927 B.n537 B.n30 10.6151
R928 B.n537 B.n536 10.6151
R929 B.n536 B.n535 10.6151
R930 B.n82 B.n38 10.6151
R931 B.n85 B.n82 10.6151
R932 B.n86 B.n85 10.6151
R933 B.n89 B.n86 10.6151
R934 B.n90 B.n89 10.6151
R935 B.n93 B.n90 10.6151
R936 B.n94 B.n93 10.6151
R937 B.n97 B.n94 10.6151
R938 B.n98 B.n97 10.6151
R939 B.n101 B.n98 10.6151
R940 B.n102 B.n101 10.6151
R941 B.n105 B.n102 10.6151
R942 B.n106 B.n105 10.6151
R943 B.n109 B.n106 10.6151
R944 B.n110 B.n109 10.6151
R945 B.n113 B.n110 10.6151
R946 B.n114 B.n113 10.6151
R947 B.n117 B.n114 10.6151
R948 B.n118 B.n117 10.6151
R949 B.n121 B.n118 10.6151
R950 B.n122 B.n121 10.6151
R951 B.n125 B.n122 10.6151
R952 B.n126 B.n125 10.6151
R953 B.n129 B.n126 10.6151
R954 B.n130 B.n129 10.6151
R955 B.n133 B.n130 10.6151
R956 B.n134 B.n133 10.6151
R957 B.n137 B.n134 10.6151
R958 B.n138 B.n137 10.6151
R959 B.n141 B.n138 10.6151
R960 B.n146 B.n143 10.6151
R961 B.n147 B.n146 10.6151
R962 B.n150 B.n147 10.6151
R963 B.n151 B.n150 10.6151
R964 B.n154 B.n151 10.6151
R965 B.n155 B.n154 10.6151
R966 B.n158 B.n155 10.6151
R967 B.n159 B.n158 10.6151
R968 B.n163 B.n162 10.6151
R969 B.n166 B.n163 10.6151
R970 B.n167 B.n166 10.6151
R971 B.n170 B.n167 10.6151
R972 B.n171 B.n170 10.6151
R973 B.n174 B.n171 10.6151
R974 B.n175 B.n174 10.6151
R975 B.n178 B.n175 10.6151
R976 B.n179 B.n178 10.6151
R977 B.n182 B.n179 10.6151
R978 B.n183 B.n182 10.6151
R979 B.n186 B.n183 10.6151
R980 B.n187 B.n186 10.6151
R981 B.n190 B.n187 10.6151
R982 B.n191 B.n190 10.6151
R983 B.n194 B.n191 10.6151
R984 B.n195 B.n194 10.6151
R985 B.n198 B.n195 10.6151
R986 B.n199 B.n198 10.6151
R987 B.n202 B.n199 10.6151
R988 B.n203 B.n202 10.6151
R989 B.n206 B.n203 10.6151
R990 B.n207 B.n206 10.6151
R991 B.n210 B.n207 10.6151
R992 B.n211 B.n210 10.6151
R993 B.n214 B.n211 10.6151
R994 B.n215 B.n214 10.6151
R995 B.n218 B.n215 10.6151
R996 B.n219 B.n218 10.6151
R997 B.n530 B.n219 10.6151
R998 B.n453 B.t5 9.69569
R999 B.n32 B.t12 9.69569
R1000 B.n577 B.n0 8.11757
R1001 B.n577 B.n1 8.11757
R1002 B.n356 B.n355 6.5566
R1003 B.n375 B.n374 6.5566
R1004 B.n143 B.n142 6.5566
R1005 B.n159 B.n79 6.5566
R1006 B.n355 B.n354 4.05904
R1007 B.n374 B.n273 4.05904
R1008 B.n142 B.n141 4.05904
R1009 B.n162 B.n79 4.05904
R1010 VN.n0 VN.t3 237.042
R1011 VN.n1 VN.t2 237.042
R1012 VN.n1 VN.t1 236.953
R1013 VN.n0 VN.t0 236.953
R1014 VN VN.n1 70.5539
R1015 VN VN.n0 31.2622
R1016 VDD2.n2 VDD2.n0 101.79
R1017 VDD2.n2 VDD2.n1 67.1865
R1018 VDD2.n1 VDD2.t2 2.3746
R1019 VDD2.n1 VDD2.t1 2.3746
R1020 VDD2.n0 VDD2.t0 2.3746
R1021 VDD2.n0 VDD2.t3 2.3746
R1022 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 2.71938f
C1 VDD1 VDD2 0.66245f
C2 VP VTAIL 2.56554f
C3 VN VTAIL 2.55143f
C4 VP VN 4.42695f
C5 VDD1 VTAIL 4.6143f
C6 VDD1 VP 2.87024f
C7 VDD1 VN 0.14809f
C8 VDD2 VTAIL 4.658451f
C9 VP VDD2 0.299303f
C10 VDD2 B 2.643013f
C11 VDD1 B 5.9183f
C12 VTAIL B 6.992882f
C13 VN B 8.0495f
C14 VP B 5.510529f
C15 VDD2.t0 B 0.178826f
C16 VDD2.t3 B 0.178826f
C17 VDD2.n0 B 2.01175f
C18 VDD2.t2 B 0.178826f
C19 VDD2.t1 B 0.178826f
C20 VDD2.n1 B 1.55534f
C21 VDD2.n2 B 3.00397f
C22 VN.t3 B 1.14017f
C23 VN.t0 B 1.13997f
C24 VN.n0 B 0.863373f
C25 VN.t2 B 1.14017f
C26 VN.t1 B 1.13997f
C27 VN.n1 B 1.80303f
C28 VDD1.t1 B 0.178821f
C29 VDD1.t3 B 0.178821f
C30 VDD1.n0 B 1.55559f
C31 VDD1.t0 B 0.178821f
C32 VDD1.t2 B 0.178821f
C33 VDD1.n1 B 2.0352f
C34 VTAIL.t0 B 1.18228f
C35 VTAIL.n0 B 0.267537f
C36 VTAIL.t7 B 1.18228f
C37 VTAIL.n1 B 0.298016f
C38 VTAIL.t5 B 1.18228f
C39 VTAIL.n2 B 0.962434f
C40 VTAIL.t1 B 1.18228f
C41 VTAIL.n3 B 0.962425f
C42 VTAIL.t2 B 1.18228f
C43 VTAIL.n4 B 0.298008f
C44 VTAIL.t6 B 1.18228f
C45 VTAIL.n5 B 0.298008f
C46 VTAIL.t4 B 1.18228f
C47 VTAIL.n6 B 0.962434f
C48 VTAIL.t3 B 1.18228f
C49 VTAIL.n7 B 0.9256f
C50 VP.t0 B 1.17058f
C51 VP.t2 B 1.17078f
C52 VP.n0 B 1.83474f
C53 VP.n1 B 2.39717f
C54 VP.t3 B 1.13304f
C55 VP.n2 B 0.480322f
C56 VP.t1 B 1.13304f
C57 VP.n3 B 0.480322f
C58 VP.n4 B 0.054634f
.ends

