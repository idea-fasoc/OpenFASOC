* NGSPICE file created from diff_pair_sample_0383.ext - technology: sky130A

.subckt diff_pair_sample_0383 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t1 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=2.9865 ps=18.43 w=18.1 l=1.88
X1 VDD1.t3 VP.t0 VTAIL.t0 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=2.9865 pd=18.43 as=7.059 ps=36.98 w=18.1 l=1.88
X2 VDD2.t0 VN.t1 VTAIL.t5 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=2.9865 pd=18.43 as=7.059 ps=36.98 w=18.1 l=1.88
X3 VDD1.t2 VP.t1 VTAIL.t7 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=2.9865 pd=18.43 as=7.059 ps=36.98 w=18.1 l=1.88
X4 VTAIL.t2 VP.t2 VDD1.t1 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=2.9865 ps=18.43 w=18.1 l=1.88
X5 VDD2.t3 VN.t2 VTAIL.t4 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=2.9865 pd=18.43 as=7.059 ps=36.98 w=18.1 l=1.88
X6 B.t11 B.t9 B.t10 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=0 ps=0 w=18.1 l=1.88
X7 B.t8 B.t6 B.t7 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=0 ps=0 w=18.1 l=1.88
X8 VTAIL.t3 VN.t3 VDD2.t2 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=2.9865 ps=18.43 w=18.1 l=1.88
X9 B.t5 B.t3 B.t4 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=0 ps=0 w=18.1 l=1.88
X10 B.t2 B.t0 B.t1 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=0 ps=0 w=18.1 l=1.88
X11 VTAIL.t1 VP.t3 VDD1.t0 w_n2296_n4588# sky130_fd_pr__pfet_01v8 ad=7.059 pd=36.98 as=2.9865 ps=18.43 w=18.1 l=1.88
R0 VN.n0 VN.t0 269.659
R1 VN.n1 VN.t2 269.659
R2 VN.n0 VN.t1 269.221
R3 VN.n1 VN.t3 269.221
R4 VN VN.n1 58.2164
R5 VN VN.n0 9.14446
R6 VDD2.n2 VDD2.n0 117.639
R7 VDD2.n2 VDD2.n1 72.6043
R8 VDD2.n1 VDD2.t2 1.79636
R9 VDD2.n1 VDD2.t3 1.79636
R10 VDD2.n0 VDD2.t1 1.79636
R11 VDD2.n0 VDD2.t0 1.79636
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n798 VTAIL.n797 756.745
R14 VTAIL.n98 VTAIL.n97 756.745
R15 VTAIL.n198 VTAIL.n197 756.745
R16 VTAIL.n298 VTAIL.n297 756.745
R17 VTAIL.n698 VTAIL.n697 756.745
R18 VTAIL.n598 VTAIL.n597 756.745
R19 VTAIL.n498 VTAIL.n497 756.745
R20 VTAIL.n398 VTAIL.n397 756.745
R21 VTAIL.n733 VTAIL.n732 585
R22 VTAIL.n730 VTAIL.n729 585
R23 VTAIL.n739 VTAIL.n738 585
R24 VTAIL.n741 VTAIL.n740 585
R25 VTAIL.n726 VTAIL.n725 585
R26 VTAIL.n747 VTAIL.n746 585
R27 VTAIL.n750 VTAIL.n749 585
R28 VTAIL.n748 VTAIL.n722 585
R29 VTAIL.n755 VTAIL.n721 585
R30 VTAIL.n757 VTAIL.n756 585
R31 VTAIL.n759 VTAIL.n758 585
R32 VTAIL.n718 VTAIL.n717 585
R33 VTAIL.n765 VTAIL.n764 585
R34 VTAIL.n767 VTAIL.n766 585
R35 VTAIL.n714 VTAIL.n713 585
R36 VTAIL.n773 VTAIL.n772 585
R37 VTAIL.n775 VTAIL.n774 585
R38 VTAIL.n710 VTAIL.n709 585
R39 VTAIL.n781 VTAIL.n780 585
R40 VTAIL.n783 VTAIL.n782 585
R41 VTAIL.n706 VTAIL.n705 585
R42 VTAIL.n789 VTAIL.n788 585
R43 VTAIL.n791 VTAIL.n790 585
R44 VTAIL.n702 VTAIL.n701 585
R45 VTAIL.n797 VTAIL.n796 585
R46 VTAIL.n33 VTAIL.n32 585
R47 VTAIL.n30 VTAIL.n29 585
R48 VTAIL.n39 VTAIL.n38 585
R49 VTAIL.n41 VTAIL.n40 585
R50 VTAIL.n26 VTAIL.n25 585
R51 VTAIL.n47 VTAIL.n46 585
R52 VTAIL.n50 VTAIL.n49 585
R53 VTAIL.n48 VTAIL.n22 585
R54 VTAIL.n55 VTAIL.n21 585
R55 VTAIL.n57 VTAIL.n56 585
R56 VTAIL.n59 VTAIL.n58 585
R57 VTAIL.n18 VTAIL.n17 585
R58 VTAIL.n65 VTAIL.n64 585
R59 VTAIL.n67 VTAIL.n66 585
R60 VTAIL.n14 VTAIL.n13 585
R61 VTAIL.n73 VTAIL.n72 585
R62 VTAIL.n75 VTAIL.n74 585
R63 VTAIL.n10 VTAIL.n9 585
R64 VTAIL.n81 VTAIL.n80 585
R65 VTAIL.n83 VTAIL.n82 585
R66 VTAIL.n6 VTAIL.n5 585
R67 VTAIL.n89 VTAIL.n88 585
R68 VTAIL.n91 VTAIL.n90 585
R69 VTAIL.n2 VTAIL.n1 585
R70 VTAIL.n97 VTAIL.n96 585
R71 VTAIL.n133 VTAIL.n132 585
R72 VTAIL.n130 VTAIL.n129 585
R73 VTAIL.n139 VTAIL.n138 585
R74 VTAIL.n141 VTAIL.n140 585
R75 VTAIL.n126 VTAIL.n125 585
R76 VTAIL.n147 VTAIL.n146 585
R77 VTAIL.n150 VTAIL.n149 585
R78 VTAIL.n148 VTAIL.n122 585
R79 VTAIL.n155 VTAIL.n121 585
R80 VTAIL.n157 VTAIL.n156 585
R81 VTAIL.n159 VTAIL.n158 585
R82 VTAIL.n118 VTAIL.n117 585
R83 VTAIL.n165 VTAIL.n164 585
R84 VTAIL.n167 VTAIL.n166 585
R85 VTAIL.n114 VTAIL.n113 585
R86 VTAIL.n173 VTAIL.n172 585
R87 VTAIL.n175 VTAIL.n174 585
R88 VTAIL.n110 VTAIL.n109 585
R89 VTAIL.n181 VTAIL.n180 585
R90 VTAIL.n183 VTAIL.n182 585
R91 VTAIL.n106 VTAIL.n105 585
R92 VTAIL.n189 VTAIL.n188 585
R93 VTAIL.n191 VTAIL.n190 585
R94 VTAIL.n102 VTAIL.n101 585
R95 VTAIL.n197 VTAIL.n196 585
R96 VTAIL.n233 VTAIL.n232 585
R97 VTAIL.n230 VTAIL.n229 585
R98 VTAIL.n239 VTAIL.n238 585
R99 VTAIL.n241 VTAIL.n240 585
R100 VTAIL.n226 VTAIL.n225 585
R101 VTAIL.n247 VTAIL.n246 585
R102 VTAIL.n250 VTAIL.n249 585
R103 VTAIL.n248 VTAIL.n222 585
R104 VTAIL.n255 VTAIL.n221 585
R105 VTAIL.n257 VTAIL.n256 585
R106 VTAIL.n259 VTAIL.n258 585
R107 VTAIL.n218 VTAIL.n217 585
R108 VTAIL.n265 VTAIL.n264 585
R109 VTAIL.n267 VTAIL.n266 585
R110 VTAIL.n214 VTAIL.n213 585
R111 VTAIL.n273 VTAIL.n272 585
R112 VTAIL.n275 VTAIL.n274 585
R113 VTAIL.n210 VTAIL.n209 585
R114 VTAIL.n281 VTAIL.n280 585
R115 VTAIL.n283 VTAIL.n282 585
R116 VTAIL.n206 VTAIL.n205 585
R117 VTAIL.n289 VTAIL.n288 585
R118 VTAIL.n291 VTAIL.n290 585
R119 VTAIL.n202 VTAIL.n201 585
R120 VTAIL.n297 VTAIL.n296 585
R121 VTAIL.n697 VTAIL.n696 585
R122 VTAIL.n602 VTAIL.n601 585
R123 VTAIL.n691 VTAIL.n690 585
R124 VTAIL.n689 VTAIL.n688 585
R125 VTAIL.n606 VTAIL.n605 585
R126 VTAIL.n683 VTAIL.n682 585
R127 VTAIL.n681 VTAIL.n680 585
R128 VTAIL.n610 VTAIL.n609 585
R129 VTAIL.n675 VTAIL.n674 585
R130 VTAIL.n673 VTAIL.n672 585
R131 VTAIL.n614 VTAIL.n613 585
R132 VTAIL.n667 VTAIL.n666 585
R133 VTAIL.n665 VTAIL.n664 585
R134 VTAIL.n618 VTAIL.n617 585
R135 VTAIL.n659 VTAIL.n658 585
R136 VTAIL.n657 VTAIL.n656 585
R137 VTAIL.n655 VTAIL.n621 585
R138 VTAIL.n625 VTAIL.n622 585
R139 VTAIL.n650 VTAIL.n649 585
R140 VTAIL.n648 VTAIL.n647 585
R141 VTAIL.n627 VTAIL.n626 585
R142 VTAIL.n642 VTAIL.n641 585
R143 VTAIL.n640 VTAIL.n639 585
R144 VTAIL.n631 VTAIL.n630 585
R145 VTAIL.n634 VTAIL.n633 585
R146 VTAIL.n597 VTAIL.n596 585
R147 VTAIL.n502 VTAIL.n501 585
R148 VTAIL.n591 VTAIL.n590 585
R149 VTAIL.n589 VTAIL.n588 585
R150 VTAIL.n506 VTAIL.n505 585
R151 VTAIL.n583 VTAIL.n582 585
R152 VTAIL.n581 VTAIL.n580 585
R153 VTAIL.n510 VTAIL.n509 585
R154 VTAIL.n575 VTAIL.n574 585
R155 VTAIL.n573 VTAIL.n572 585
R156 VTAIL.n514 VTAIL.n513 585
R157 VTAIL.n567 VTAIL.n566 585
R158 VTAIL.n565 VTAIL.n564 585
R159 VTAIL.n518 VTAIL.n517 585
R160 VTAIL.n559 VTAIL.n558 585
R161 VTAIL.n557 VTAIL.n556 585
R162 VTAIL.n555 VTAIL.n521 585
R163 VTAIL.n525 VTAIL.n522 585
R164 VTAIL.n550 VTAIL.n549 585
R165 VTAIL.n548 VTAIL.n547 585
R166 VTAIL.n527 VTAIL.n526 585
R167 VTAIL.n542 VTAIL.n541 585
R168 VTAIL.n540 VTAIL.n539 585
R169 VTAIL.n531 VTAIL.n530 585
R170 VTAIL.n534 VTAIL.n533 585
R171 VTAIL.n497 VTAIL.n496 585
R172 VTAIL.n402 VTAIL.n401 585
R173 VTAIL.n491 VTAIL.n490 585
R174 VTAIL.n489 VTAIL.n488 585
R175 VTAIL.n406 VTAIL.n405 585
R176 VTAIL.n483 VTAIL.n482 585
R177 VTAIL.n481 VTAIL.n480 585
R178 VTAIL.n410 VTAIL.n409 585
R179 VTAIL.n475 VTAIL.n474 585
R180 VTAIL.n473 VTAIL.n472 585
R181 VTAIL.n414 VTAIL.n413 585
R182 VTAIL.n467 VTAIL.n466 585
R183 VTAIL.n465 VTAIL.n464 585
R184 VTAIL.n418 VTAIL.n417 585
R185 VTAIL.n459 VTAIL.n458 585
R186 VTAIL.n457 VTAIL.n456 585
R187 VTAIL.n455 VTAIL.n421 585
R188 VTAIL.n425 VTAIL.n422 585
R189 VTAIL.n450 VTAIL.n449 585
R190 VTAIL.n448 VTAIL.n447 585
R191 VTAIL.n427 VTAIL.n426 585
R192 VTAIL.n442 VTAIL.n441 585
R193 VTAIL.n440 VTAIL.n439 585
R194 VTAIL.n431 VTAIL.n430 585
R195 VTAIL.n434 VTAIL.n433 585
R196 VTAIL.n397 VTAIL.n396 585
R197 VTAIL.n302 VTAIL.n301 585
R198 VTAIL.n391 VTAIL.n390 585
R199 VTAIL.n389 VTAIL.n388 585
R200 VTAIL.n306 VTAIL.n305 585
R201 VTAIL.n383 VTAIL.n382 585
R202 VTAIL.n381 VTAIL.n380 585
R203 VTAIL.n310 VTAIL.n309 585
R204 VTAIL.n375 VTAIL.n374 585
R205 VTAIL.n373 VTAIL.n372 585
R206 VTAIL.n314 VTAIL.n313 585
R207 VTAIL.n367 VTAIL.n366 585
R208 VTAIL.n365 VTAIL.n364 585
R209 VTAIL.n318 VTAIL.n317 585
R210 VTAIL.n359 VTAIL.n358 585
R211 VTAIL.n357 VTAIL.n356 585
R212 VTAIL.n355 VTAIL.n321 585
R213 VTAIL.n325 VTAIL.n322 585
R214 VTAIL.n350 VTAIL.n349 585
R215 VTAIL.n348 VTAIL.n347 585
R216 VTAIL.n327 VTAIL.n326 585
R217 VTAIL.n342 VTAIL.n341 585
R218 VTAIL.n340 VTAIL.n339 585
R219 VTAIL.n331 VTAIL.n330 585
R220 VTAIL.n334 VTAIL.n333 585
R221 VTAIL.t5 VTAIL.n731 329.036
R222 VTAIL.t6 VTAIL.n31 329.036
R223 VTAIL.t7 VTAIL.n131 329.036
R224 VTAIL.t2 VTAIL.n231 329.036
R225 VTAIL.t1 VTAIL.n532 329.036
R226 VTAIL.t4 VTAIL.n432 329.036
R227 VTAIL.t3 VTAIL.n332 329.036
R228 VTAIL.t0 VTAIL.n632 329.036
R229 VTAIL.n732 VTAIL.n729 171.744
R230 VTAIL.n739 VTAIL.n729 171.744
R231 VTAIL.n740 VTAIL.n739 171.744
R232 VTAIL.n740 VTAIL.n725 171.744
R233 VTAIL.n747 VTAIL.n725 171.744
R234 VTAIL.n749 VTAIL.n747 171.744
R235 VTAIL.n749 VTAIL.n748 171.744
R236 VTAIL.n748 VTAIL.n721 171.744
R237 VTAIL.n757 VTAIL.n721 171.744
R238 VTAIL.n758 VTAIL.n757 171.744
R239 VTAIL.n758 VTAIL.n717 171.744
R240 VTAIL.n765 VTAIL.n717 171.744
R241 VTAIL.n766 VTAIL.n765 171.744
R242 VTAIL.n766 VTAIL.n713 171.744
R243 VTAIL.n773 VTAIL.n713 171.744
R244 VTAIL.n774 VTAIL.n773 171.744
R245 VTAIL.n774 VTAIL.n709 171.744
R246 VTAIL.n781 VTAIL.n709 171.744
R247 VTAIL.n782 VTAIL.n781 171.744
R248 VTAIL.n782 VTAIL.n705 171.744
R249 VTAIL.n789 VTAIL.n705 171.744
R250 VTAIL.n790 VTAIL.n789 171.744
R251 VTAIL.n790 VTAIL.n701 171.744
R252 VTAIL.n797 VTAIL.n701 171.744
R253 VTAIL.n32 VTAIL.n29 171.744
R254 VTAIL.n39 VTAIL.n29 171.744
R255 VTAIL.n40 VTAIL.n39 171.744
R256 VTAIL.n40 VTAIL.n25 171.744
R257 VTAIL.n47 VTAIL.n25 171.744
R258 VTAIL.n49 VTAIL.n47 171.744
R259 VTAIL.n49 VTAIL.n48 171.744
R260 VTAIL.n48 VTAIL.n21 171.744
R261 VTAIL.n57 VTAIL.n21 171.744
R262 VTAIL.n58 VTAIL.n57 171.744
R263 VTAIL.n58 VTAIL.n17 171.744
R264 VTAIL.n65 VTAIL.n17 171.744
R265 VTAIL.n66 VTAIL.n65 171.744
R266 VTAIL.n66 VTAIL.n13 171.744
R267 VTAIL.n73 VTAIL.n13 171.744
R268 VTAIL.n74 VTAIL.n73 171.744
R269 VTAIL.n74 VTAIL.n9 171.744
R270 VTAIL.n81 VTAIL.n9 171.744
R271 VTAIL.n82 VTAIL.n81 171.744
R272 VTAIL.n82 VTAIL.n5 171.744
R273 VTAIL.n89 VTAIL.n5 171.744
R274 VTAIL.n90 VTAIL.n89 171.744
R275 VTAIL.n90 VTAIL.n1 171.744
R276 VTAIL.n97 VTAIL.n1 171.744
R277 VTAIL.n132 VTAIL.n129 171.744
R278 VTAIL.n139 VTAIL.n129 171.744
R279 VTAIL.n140 VTAIL.n139 171.744
R280 VTAIL.n140 VTAIL.n125 171.744
R281 VTAIL.n147 VTAIL.n125 171.744
R282 VTAIL.n149 VTAIL.n147 171.744
R283 VTAIL.n149 VTAIL.n148 171.744
R284 VTAIL.n148 VTAIL.n121 171.744
R285 VTAIL.n157 VTAIL.n121 171.744
R286 VTAIL.n158 VTAIL.n157 171.744
R287 VTAIL.n158 VTAIL.n117 171.744
R288 VTAIL.n165 VTAIL.n117 171.744
R289 VTAIL.n166 VTAIL.n165 171.744
R290 VTAIL.n166 VTAIL.n113 171.744
R291 VTAIL.n173 VTAIL.n113 171.744
R292 VTAIL.n174 VTAIL.n173 171.744
R293 VTAIL.n174 VTAIL.n109 171.744
R294 VTAIL.n181 VTAIL.n109 171.744
R295 VTAIL.n182 VTAIL.n181 171.744
R296 VTAIL.n182 VTAIL.n105 171.744
R297 VTAIL.n189 VTAIL.n105 171.744
R298 VTAIL.n190 VTAIL.n189 171.744
R299 VTAIL.n190 VTAIL.n101 171.744
R300 VTAIL.n197 VTAIL.n101 171.744
R301 VTAIL.n232 VTAIL.n229 171.744
R302 VTAIL.n239 VTAIL.n229 171.744
R303 VTAIL.n240 VTAIL.n239 171.744
R304 VTAIL.n240 VTAIL.n225 171.744
R305 VTAIL.n247 VTAIL.n225 171.744
R306 VTAIL.n249 VTAIL.n247 171.744
R307 VTAIL.n249 VTAIL.n248 171.744
R308 VTAIL.n248 VTAIL.n221 171.744
R309 VTAIL.n257 VTAIL.n221 171.744
R310 VTAIL.n258 VTAIL.n257 171.744
R311 VTAIL.n258 VTAIL.n217 171.744
R312 VTAIL.n265 VTAIL.n217 171.744
R313 VTAIL.n266 VTAIL.n265 171.744
R314 VTAIL.n266 VTAIL.n213 171.744
R315 VTAIL.n273 VTAIL.n213 171.744
R316 VTAIL.n274 VTAIL.n273 171.744
R317 VTAIL.n274 VTAIL.n209 171.744
R318 VTAIL.n281 VTAIL.n209 171.744
R319 VTAIL.n282 VTAIL.n281 171.744
R320 VTAIL.n282 VTAIL.n205 171.744
R321 VTAIL.n289 VTAIL.n205 171.744
R322 VTAIL.n290 VTAIL.n289 171.744
R323 VTAIL.n290 VTAIL.n201 171.744
R324 VTAIL.n297 VTAIL.n201 171.744
R325 VTAIL.n697 VTAIL.n601 171.744
R326 VTAIL.n690 VTAIL.n601 171.744
R327 VTAIL.n690 VTAIL.n689 171.744
R328 VTAIL.n689 VTAIL.n605 171.744
R329 VTAIL.n682 VTAIL.n605 171.744
R330 VTAIL.n682 VTAIL.n681 171.744
R331 VTAIL.n681 VTAIL.n609 171.744
R332 VTAIL.n674 VTAIL.n609 171.744
R333 VTAIL.n674 VTAIL.n673 171.744
R334 VTAIL.n673 VTAIL.n613 171.744
R335 VTAIL.n666 VTAIL.n613 171.744
R336 VTAIL.n666 VTAIL.n665 171.744
R337 VTAIL.n665 VTAIL.n617 171.744
R338 VTAIL.n658 VTAIL.n617 171.744
R339 VTAIL.n658 VTAIL.n657 171.744
R340 VTAIL.n657 VTAIL.n621 171.744
R341 VTAIL.n625 VTAIL.n621 171.744
R342 VTAIL.n649 VTAIL.n625 171.744
R343 VTAIL.n649 VTAIL.n648 171.744
R344 VTAIL.n648 VTAIL.n626 171.744
R345 VTAIL.n641 VTAIL.n626 171.744
R346 VTAIL.n641 VTAIL.n640 171.744
R347 VTAIL.n640 VTAIL.n630 171.744
R348 VTAIL.n633 VTAIL.n630 171.744
R349 VTAIL.n597 VTAIL.n501 171.744
R350 VTAIL.n590 VTAIL.n501 171.744
R351 VTAIL.n590 VTAIL.n589 171.744
R352 VTAIL.n589 VTAIL.n505 171.744
R353 VTAIL.n582 VTAIL.n505 171.744
R354 VTAIL.n582 VTAIL.n581 171.744
R355 VTAIL.n581 VTAIL.n509 171.744
R356 VTAIL.n574 VTAIL.n509 171.744
R357 VTAIL.n574 VTAIL.n573 171.744
R358 VTAIL.n573 VTAIL.n513 171.744
R359 VTAIL.n566 VTAIL.n513 171.744
R360 VTAIL.n566 VTAIL.n565 171.744
R361 VTAIL.n565 VTAIL.n517 171.744
R362 VTAIL.n558 VTAIL.n517 171.744
R363 VTAIL.n558 VTAIL.n557 171.744
R364 VTAIL.n557 VTAIL.n521 171.744
R365 VTAIL.n525 VTAIL.n521 171.744
R366 VTAIL.n549 VTAIL.n525 171.744
R367 VTAIL.n549 VTAIL.n548 171.744
R368 VTAIL.n548 VTAIL.n526 171.744
R369 VTAIL.n541 VTAIL.n526 171.744
R370 VTAIL.n541 VTAIL.n540 171.744
R371 VTAIL.n540 VTAIL.n530 171.744
R372 VTAIL.n533 VTAIL.n530 171.744
R373 VTAIL.n497 VTAIL.n401 171.744
R374 VTAIL.n490 VTAIL.n401 171.744
R375 VTAIL.n490 VTAIL.n489 171.744
R376 VTAIL.n489 VTAIL.n405 171.744
R377 VTAIL.n482 VTAIL.n405 171.744
R378 VTAIL.n482 VTAIL.n481 171.744
R379 VTAIL.n481 VTAIL.n409 171.744
R380 VTAIL.n474 VTAIL.n409 171.744
R381 VTAIL.n474 VTAIL.n473 171.744
R382 VTAIL.n473 VTAIL.n413 171.744
R383 VTAIL.n466 VTAIL.n413 171.744
R384 VTAIL.n466 VTAIL.n465 171.744
R385 VTAIL.n465 VTAIL.n417 171.744
R386 VTAIL.n458 VTAIL.n417 171.744
R387 VTAIL.n458 VTAIL.n457 171.744
R388 VTAIL.n457 VTAIL.n421 171.744
R389 VTAIL.n425 VTAIL.n421 171.744
R390 VTAIL.n449 VTAIL.n425 171.744
R391 VTAIL.n449 VTAIL.n448 171.744
R392 VTAIL.n448 VTAIL.n426 171.744
R393 VTAIL.n441 VTAIL.n426 171.744
R394 VTAIL.n441 VTAIL.n440 171.744
R395 VTAIL.n440 VTAIL.n430 171.744
R396 VTAIL.n433 VTAIL.n430 171.744
R397 VTAIL.n397 VTAIL.n301 171.744
R398 VTAIL.n390 VTAIL.n301 171.744
R399 VTAIL.n390 VTAIL.n389 171.744
R400 VTAIL.n389 VTAIL.n305 171.744
R401 VTAIL.n382 VTAIL.n305 171.744
R402 VTAIL.n382 VTAIL.n381 171.744
R403 VTAIL.n381 VTAIL.n309 171.744
R404 VTAIL.n374 VTAIL.n309 171.744
R405 VTAIL.n374 VTAIL.n373 171.744
R406 VTAIL.n373 VTAIL.n313 171.744
R407 VTAIL.n366 VTAIL.n313 171.744
R408 VTAIL.n366 VTAIL.n365 171.744
R409 VTAIL.n365 VTAIL.n317 171.744
R410 VTAIL.n358 VTAIL.n317 171.744
R411 VTAIL.n358 VTAIL.n357 171.744
R412 VTAIL.n357 VTAIL.n321 171.744
R413 VTAIL.n325 VTAIL.n321 171.744
R414 VTAIL.n349 VTAIL.n325 171.744
R415 VTAIL.n349 VTAIL.n348 171.744
R416 VTAIL.n348 VTAIL.n326 171.744
R417 VTAIL.n341 VTAIL.n326 171.744
R418 VTAIL.n341 VTAIL.n340 171.744
R419 VTAIL.n340 VTAIL.n330 171.744
R420 VTAIL.n333 VTAIL.n330 171.744
R421 VTAIL.n732 VTAIL.t5 85.8723
R422 VTAIL.n32 VTAIL.t6 85.8723
R423 VTAIL.n132 VTAIL.t7 85.8723
R424 VTAIL.n232 VTAIL.t2 85.8723
R425 VTAIL.n633 VTAIL.t0 85.8723
R426 VTAIL.n533 VTAIL.t1 85.8723
R427 VTAIL.n433 VTAIL.t4 85.8723
R428 VTAIL.n333 VTAIL.t3 85.8723
R429 VTAIL.n799 VTAIL.n798 35.2884
R430 VTAIL.n99 VTAIL.n98 35.2884
R431 VTAIL.n199 VTAIL.n198 35.2884
R432 VTAIL.n299 VTAIL.n298 35.2884
R433 VTAIL.n699 VTAIL.n698 35.2884
R434 VTAIL.n599 VTAIL.n598 35.2884
R435 VTAIL.n499 VTAIL.n498 35.2884
R436 VTAIL.n399 VTAIL.n398 35.2884
R437 VTAIL.n799 VTAIL.n699 29.8755
R438 VTAIL.n399 VTAIL.n299 29.8755
R439 VTAIL.n756 VTAIL.n755 13.1884
R440 VTAIL.n56 VTAIL.n55 13.1884
R441 VTAIL.n156 VTAIL.n155 13.1884
R442 VTAIL.n256 VTAIL.n255 13.1884
R443 VTAIL.n656 VTAIL.n655 13.1884
R444 VTAIL.n556 VTAIL.n555 13.1884
R445 VTAIL.n456 VTAIL.n455 13.1884
R446 VTAIL.n356 VTAIL.n355 13.1884
R447 VTAIL.n754 VTAIL.n722 12.8005
R448 VTAIL.n759 VTAIL.n720 12.8005
R449 VTAIL.n54 VTAIL.n22 12.8005
R450 VTAIL.n59 VTAIL.n20 12.8005
R451 VTAIL.n154 VTAIL.n122 12.8005
R452 VTAIL.n159 VTAIL.n120 12.8005
R453 VTAIL.n254 VTAIL.n222 12.8005
R454 VTAIL.n259 VTAIL.n220 12.8005
R455 VTAIL.n659 VTAIL.n620 12.8005
R456 VTAIL.n654 VTAIL.n622 12.8005
R457 VTAIL.n559 VTAIL.n520 12.8005
R458 VTAIL.n554 VTAIL.n522 12.8005
R459 VTAIL.n459 VTAIL.n420 12.8005
R460 VTAIL.n454 VTAIL.n422 12.8005
R461 VTAIL.n359 VTAIL.n320 12.8005
R462 VTAIL.n354 VTAIL.n322 12.8005
R463 VTAIL.n751 VTAIL.n750 12.0247
R464 VTAIL.n760 VTAIL.n718 12.0247
R465 VTAIL.n796 VTAIL.n700 12.0247
R466 VTAIL.n51 VTAIL.n50 12.0247
R467 VTAIL.n60 VTAIL.n18 12.0247
R468 VTAIL.n96 VTAIL.n0 12.0247
R469 VTAIL.n151 VTAIL.n150 12.0247
R470 VTAIL.n160 VTAIL.n118 12.0247
R471 VTAIL.n196 VTAIL.n100 12.0247
R472 VTAIL.n251 VTAIL.n250 12.0247
R473 VTAIL.n260 VTAIL.n218 12.0247
R474 VTAIL.n296 VTAIL.n200 12.0247
R475 VTAIL.n696 VTAIL.n600 12.0247
R476 VTAIL.n660 VTAIL.n618 12.0247
R477 VTAIL.n651 VTAIL.n650 12.0247
R478 VTAIL.n596 VTAIL.n500 12.0247
R479 VTAIL.n560 VTAIL.n518 12.0247
R480 VTAIL.n551 VTAIL.n550 12.0247
R481 VTAIL.n496 VTAIL.n400 12.0247
R482 VTAIL.n460 VTAIL.n418 12.0247
R483 VTAIL.n451 VTAIL.n450 12.0247
R484 VTAIL.n396 VTAIL.n300 12.0247
R485 VTAIL.n360 VTAIL.n318 12.0247
R486 VTAIL.n351 VTAIL.n350 12.0247
R487 VTAIL.n746 VTAIL.n724 11.249
R488 VTAIL.n764 VTAIL.n763 11.249
R489 VTAIL.n795 VTAIL.n702 11.249
R490 VTAIL.n46 VTAIL.n24 11.249
R491 VTAIL.n64 VTAIL.n63 11.249
R492 VTAIL.n95 VTAIL.n2 11.249
R493 VTAIL.n146 VTAIL.n124 11.249
R494 VTAIL.n164 VTAIL.n163 11.249
R495 VTAIL.n195 VTAIL.n102 11.249
R496 VTAIL.n246 VTAIL.n224 11.249
R497 VTAIL.n264 VTAIL.n263 11.249
R498 VTAIL.n295 VTAIL.n202 11.249
R499 VTAIL.n695 VTAIL.n602 11.249
R500 VTAIL.n664 VTAIL.n663 11.249
R501 VTAIL.n647 VTAIL.n624 11.249
R502 VTAIL.n595 VTAIL.n502 11.249
R503 VTAIL.n564 VTAIL.n563 11.249
R504 VTAIL.n547 VTAIL.n524 11.249
R505 VTAIL.n495 VTAIL.n402 11.249
R506 VTAIL.n464 VTAIL.n463 11.249
R507 VTAIL.n447 VTAIL.n424 11.249
R508 VTAIL.n395 VTAIL.n302 11.249
R509 VTAIL.n364 VTAIL.n363 11.249
R510 VTAIL.n347 VTAIL.n324 11.249
R511 VTAIL.n733 VTAIL.n731 10.7239
R512 VTAIL.n33 VTAIL.n31 10.7239
R513 VTAIL.n133 VTAIL.n131 10.7239
R514 VTAIL.n233 VTAIL.n231 10.7239
R515 VTAIL.n634 VTAIL.n632 10.7239
R516 VTAIL.n534 VTAIL.n532 10.7239
R517 VTAIL.n434 VTAIL.n432 10.7239
R518 VTAIL.n334 VTAIL.n332 10.7239
R519 VTAIL.n745 VTAIL.n726 10.4732
R520 VTAIL.n767 VTAIL.n716 10.4732
R521 VTAIL.n792 VTAIL.n791 10.4732
R522 VTAIL.n45 VTAIL.n26 10.4732
R523 VTAIL.n67 VTAIL.n16 10.4732
R524 VTAIL.n92 VTAIL.n91 10.4732
R525 VTAIL.n145 VTAIL.n126 10.4732
R526 VTAIL.n167 VTAIL.n116 10.4732
R527 VTAIL.n192 VTAIL.n191 10.4732
R528 VTAIL.n245 VTAIL.n226 10.4732
R529 VTAIL.n267 VTAIL.n216 10.4732
R530 VTAIL.n292 VTAIL.n291 10.4732
R531 VTAIL.n692 VTAIL.n691 10.4732
R532 VTAIL.n667 VTAIL.n616 10.4732
R533 VTAIL.n646 VTAIL.n627 10.4732
R534 VTAIL.n592 VTAIL.n591 10.4732
R535 VTAIL.n567 VTAIL.n516 10.4732
R536 VTAIL.n546 VTAIL.n527 10.4732
R537 VTAIL.n492 VTAIL.n491 10.4732
R538 VTAIL.n467 VTAIL.n416 10.4732
R539 VTAIL.n446 VTAIL.n427 10.4732
R540 VTAIL.n392 VTAIL.n391 10.4732
R541 VTAIL.n367 VTAIL.n316 10.4732
R542 VTAIL.n346 VTAIL.n327 10.4732
R543 VTAIL.n742 VTAIL.n741 9.69747
R544 VTAIL.n768 VTAIL.n714 9.69747
R545 VTAIL.n788 VTAIL.n704 9.69747
R546 VTAIL.n42 VTAIL.n41 9.69747
R547 VTAIL.n68 VTAIL.n14 9.69747
R548 VTAIL.n88 VTAIL.n4 9.69747
R549 VTAIL.n142 VTAIL.n141 9.69747
R550 VTAIL.n168 VTAIL.n114 9.69747
R551 VTAIL.n188 VTAIL.n104 9.69747
R552 VTAIL.n242 VTAIL.n241 9.69747
R553 VTAIL.n268 VTAIL.n214 9.69747
R554 VTAIL.n288 VTAIL.n204 9.69747
R555 VTAIL.n688 VTAIL.n604 9.69747
R556 VTAIL.n668 VTAIL.n614 9.69747
R557 VTAIL.n643 VTAIL.n642 9.69747
R558 VTAIL.n588 VTAIL.n504 9.69747
R559 VTAIL.n568 VTAIL.n514 9.69747
R560 VTAIL.n543 VTAIL.n542 9.69747
R561 VTAIL.n488 VTAIL.n404 9.69747
R562 VTAIL.n468 VTAIL.n414 9.69747
R563 VTAIL.n443 VTAIL.n442 9.69747
R564 VTAIL.n388 VTAIL.n304 9.69747
R565 VTAIL.n368 VTAIL.n314 9.69747
R566 VTAIL.n343 VTAIL.n342 9.69747
R567 VTAIL.n794 VTAIL.n700 9.45567
R568 VTAIL.n94 VTAIL.n0 9.45567
R569 VTAIL.n194 VTAIL.n100 9.45567
R570 VTAIL.n294 VTAIL.n200 9.45567
R571 VTAIL.n694 VTAIL.n600 9.45567
R572 VTAIL.n594 VTAIL.n500 9.45567
R573 VTAIL.n494 VTAIL.n400 9.45567
R574 VTAIL.n394 VTAIL.n300 9.45567
R575 VTAIL.n779 VTAIL.n778 9.3005
R576 VTAIL.n708 VTAIL.n707 9.3005
R577 VTAIL.n785 VTAIL.n784 9.3005
R578 VTAIL.n787 VTAIL.n786 9.3005
R579 VTAIL.n704 VTAIL.n703 9.3005
R580 VTAIL.n793 VTAIL.n792 9.3005
R581 VTAIL.n795 VTAIL.n794 9.3005
R582 VTAIL.n712 VTAIL.n711 9.3005
R583 VTAIL.n771 VTAIL.n770 9.3005
R584 VTAIL.n769 VTAIL.n768 9.3005
R585 VTAIL.n716 VTAIL.n715 9.3005
R586 VTAIL.n763 VTAIL.n762 9.3005
R587 VTAIL.n761 VTAIL.n760 9.3005
R588 VTAIL.n720 VTAIL.n719 9.3005
R589 VTAIL.n735 VTAIL.n734 9.3005
R590 VTAIL.n737 VTAIL.n736 9.3005
R591 VTAIL.n728 VTAIL.n727 9.3005
R592 VTAIL.n743 VTAIL.n742 9.3005
R593 VTAIL.n745 VTAIL.n744 9.3005
R594 VTAIL.n724 VTAIL.n723 9.3005
R595 VTAIL.n752 VTAIL.n751 9.3005
R596 VTAIL.n754 VTAIL.n753 9.3005
R597 VTAIL.n777 VTAIL.n776 9.3005
R598 VTAIL.n79 VTAIL.n78 9.3005
R599 VTAIL.n8 VTAIL.n7 9.3005
R600 VTAIL.n85 VTAIL.n84 9.3005
R601 VTAIL.n87 VTAIL.n86 9.3005
R602 VTAIL.n4 VTAIL.n3 9.3005
R603 VTAIL.n93 VTAIL.n92 9.3005
R604 VTAIL.n95 VTAIL.n94 9.3005
R605 VTAIL.n12 VTAIL.n11 9.3005
R606 VTAIL.n71 VTAIL.n70 9.3005
R607 VTAIL.n69 VTAIL.n68 9.3005
R608 VTAIL.n16 VTAIL.n15 9.3005
R609 VTAIL.n63 VTAIL.n62 9.3005
R610 VTAIL.n61 VTAIL.n60 9.3005
R611 VTAIL.n20 VTAIL.n19 9.3005
R612 VTAIL.n35 VTAIL.n34 9.3005
R613 VTAIL.n37 VTAIL.n36 9.3005
R614 VTAIL.n28 VTAIL.n27 9.3005
R615 VTAIL.n43 VTAIL.n42 9.3005
R616 VTAIL.n45 VTAIL.n44 9.3005
R617 VTAIL.n24 VTAIL.n23 9.3005
R618 VTAIL.n52 VTAIL.n51 9.3005
R619 VTAIL.n54 VTAIL.n53 9.3005
R620 VTAIL.n77 VTAIL.n76 9.3005
R621 VTAIL.n179 VTAIL.n178 9.3005
R622 VTAIL.n108 VTAIL.n107 9.3005
R623 VTAIL.n185 VTAIL.n184 9.3005
R624 VTAIL.n187 VTAIL.n186 9.3005
R625 VTAIL.n104 VTAIL.n103 9.3005
R626 VTAIL.n193 VTAIL.n192 9.3005
R627 VTAIL.n195 VTAIL.n194 9.3005
R628 VTAIL.n112 VTAIL.n111 9.3005
R629 VTAIL.n171 VTAIL.n170 9.3005
R630 VTAIL.n169 VTAIL.n168 9.3005
R631 VTAIL.n116 VTAIL.n115 9.3005
R632 VTAIL.n163 VTAIL.n162 9.3005
R633 VTAIL.n161 VTAIL.n160 9.3005
R634 VTAIL.n120 VTAIL.n119 9.3005
R635 VTAIL.n135 VTAIL.n134 9.3005
R636 VTAIL.n137 VTAIL.n136 9.3005
R637 VTAIL.n128 VTAIL.n127 9.3005
R638 VTAIL.n143 VTAIL.n142 9.3005
R639 VTAIL.n145 VTAIL.n144 9.3005
R640 VTAIL.n124 VTAIL.n123 9.3005
R641 VTAIL.n152 VTAIL.n151 9.3005
R642 VTAIL.n154 VTAIL.n153 9.3005
R643 VTAIL.n177 VTAIL.n176 9.3005
R644 VTAIL.n279 VTAIL.n278 9.3005
R645 VTAIL.n208 VTAIL.n207 9.3005
R646 VTAIL.n285 VTAIL.n284 9.3005
R647 VTAIL.n287 VTAIL.n286 9.3005
R648 VTAIL.n204 VTAIL.n203 9.3005
R649 VTAIL.n293 VTAIL.n292 9.3005
R650 VTAIL.n295 VTAIL.n294 9.3005
R651 VTAIL.n212 VTAIL.n211 9.3005
R652 VTAIL.n271 VTAIL.n270 9.3005
R653 VTAIL.n269 VTAIL.n268 9.3005
R654 VTAIL.n216 VTAIL.n215 9.3005
R655 VTAIL.n263 VTAIL.n262 9.3005
R656 VTAIL.n261 VTAIL.n260 9.3005
R657 VTAIL.n220 VTAIL.n219 9.3005
R658 VTAIL.n235 VTAIL.n234 9.3005
R659 VTAIL.n237 VTAIL.n236 9.3005
R660 VTAIL.n228 VTAIL.n227 9.3005
R661 VTAIL.n243 VTAIL.n242 9.3005
R662 VTAIL.n245 VTAIL.n244 9.3005
R663 VTAIL.n224 VTAIL.n223 9.3005
R664 VTAIL.n252 VTAIL.n251 9.3005
R665 VTAIL.n254 VTAIL.n253 9.3005
R666 VTAIL.n277 VTAIL.n276 9.3005
R667 VTAIL.n695 VTAIL.n694 9.3005
R668 VTAIL.n693 VTAIL.n692 9.3005
R669 VTAIL.n604 VTAIL.n603 9.3005
R670 VTAIL.n687 VTAIL.n686 9.3005
R671 VTAIL.n685 VTAIL.n684 9.3005
R672 VTAIL.n608 VTAIL.n607 9.3005
R673 VTAIL.n679 VTAIL.n678 9.3005
R674 VTAIL.n677 VTAIL.n676 9.3005
R675 VTAIL.n612 VTAIL.n611 9.3005
R676 VTAIL.n671 VTAIL.n670 9.3005
R677 VTAIL.n669 VTAIL.n668 9.3005
R678 VTAIL.n616 VTAIL.n615 9.3005
R679 VTAIL.n663 VTAIL.n662 9.3005
R680 VTAIL.n661 VTAIL.n660 9.3005
R681 VTAIL.n620 VTAIL.n619 9.3005
R682 VTAIL.n654 VTAIL.n653 9.3005
R683 VTAIL.n652 VTAIL.n651 9.3005
R684 VTAIL.n624 VTAIL.n623 9.3005
R685 VTAIL.n646 VTAIL.n645 9.3005
R686 VTAIL.n644 VTAIL.n643 9.3005
R687 VTAIL.n629 VTAIL.n628 9.3005
R688 VTAIL.n638 VTAIL.n637 9.3005
R689 VTAIL.n636 VTAIL.n635 9.3005
R690 VTAIL.n536 VTAIL.n535 9.3005
R691 VTAIL.n538 VTAIL.n537 9.3005
R692 VTAIL.n529 VTAIL.n528 9.3005
R693 VTAIL.n544 VTAIL.n543 9.3005
R694 VTAIL.n546 VTAIL.n545 9.3005
R695 VTAIL.n524 VTAIL.n523 9.3005
R696 VTAIL.n552 VTAIL.n551 9.3005
R697 VTAIL.n554 VTAIL.n553 9.3005
R698 VTAIL.n508 VTAIL.n507 9.3005
R699 VTAIL.n585 VTAIL.n584 9.3005
R700 VTAIL.n587 VTAIL.n586 9.3005
R701 VTAIL.n504 VTAIL.n503 9.3005
R702 VTAIL.n593 VTAIL.n592 9.3005
R703 VTAIL.n595 VTAIL.n594 9.3005
R704 VTAIL.n579 VTAIL.n578 9.3005
R705 VTAIL.n577 VTAIL.n576 9.3005
R706 VTAIL.n512 VTAIL.n511 9.3005
R707 VTAIL.n571 VTAIL.n570 9.3005
R708 VTAIL.n569 VTAIL.n568 9.3005
R709 VTAIL.n516 VTAIL.n515 9.3005
R710 VTAIL.n563 VTAIL.n562 9.3005
R711 VTAIL.n561 VTAIL.n560 9.3005
R712 VTAIL.n520 VTAIL.n519 9.3005
R713 VTAIL.n436 VTAIL.n435 9.3005
R714 VTAIL.n438 VTAIL.n437 9.3005
R715 VTAIL.n429 VTAIL.n428 9.3005
R716 VTAIL.n444 VTAIL.n443 9.3005
R717 VTAIL.n446 VTAIL.n445 9.3005
R718 VTAIL.n424 VTAIL.n423 9.3005
R719 VTAIL.n452 VTAIL.n451 9.3005
R720 VTAIL.n454 VTAIL.n453 9.3005
R721 VTAIL.n408 VTAIL.n407 9.3005
R722 VTAIL.n485 VTAIL.n484 9.3005
R723 VTAIL.n487 VTAIL.n486 9.3005
R724 VTAIL.n404 VTAIL.n403 9.3005
R725 VTAIL.n493 VTAIL.n492 9.3005
R726 VTAIL.n495 VTAIL.n494 9.3005
R727 VTAIL.n479 VTAIL.n478 9.3005
R728 VTAIL.n477 VTAIL.n476 9.3005
R729 VTAIL.n412 VTAIL.n411 9.3005
R730 VTAIL.n471 VTAIL.n470 9.3005
R731 VTAIL.n469 VTAIL.n468 9.3005
R732 VTAIL.n416 VTAIL.n415 9.3005
R733 VTAIL.n463 VTAIL.n462 9.3005
R734 VTAIL.n461 VTAIL.n460 9.3005
R735 VTAIL.n420 VTAIL.n419 9.3005
R736 VTAIL.n336 VTAIL.n335 9.3005
R737 VTAIL.n338 VTAIL.n337 9.3005
R738 VTAIL.n329 VTAIL.n328 9.3005
R739 VTAIL.n344 VTAIL.n343 9.3005
R740 VTAIL.n346 VTAIL.n345 9.3005
R741 VTAIL.n324 VTAIL.n323 9.3005
R742 VTAIL.n352 VTAIL.n351 9.3005
R743 VTAIL.n354 VTAIL.n353 9.3005
R744 VTAIL.n308 VTAIL.n307 9.3005
R745 VTAIL.n385 VTAIL.n384 9.3005
R746 VTAIL.n387 VTAIL.n386 9.3005
R747 VTAIL.n304 VTAIL.n303 9.3005
R748 VTAIL.n393 VTAIL.n392 9.3005
R749 VTAIL.n395 VTAIL.n394 9.3005
R750 VTAIL.n379 VTAIL.n378 9.3005
R751 VTAIL.n377 VTAIL.n376 9.3005
R752 VTAIL.n312 VTAIL.n311 9.3005
R753 VTAIL.n371 VTAIL.n370 9.3005
R754 VTAIL.n369 VTAIL.n368 9.3005
R755 VTAIL.n316 VTAIL.n315 9.3005
R756 VTAIL.n363 VTAIL.n362 9.3005
R757 VTAIL.n361 VTAIL.n360 9.3005
R758 VTAIL.n320 VTAIL.n319 9.3005
R759 VTAIL.n738 VTAIL.n728 8.92171
R760 VTAIL.n772 VTAIL.n771 8.92171
R761 VTAIL.n787 VTAIL.n706 8.92171
R762 VTAIL.n38 VTAIL.n28 8.92171
R763 VTAIL.n72 VTAIL.n71 8.92171
R764 VTAIL.n87 VTAIL.n6 8.92171
R765 VTAIL.n138 VTAIL.n128 8.92171
R766 VTAIL.n172 VTAIL.n171 8.92171
R767 VTAIL.n187 VTAIL.n106 8.92171
R768 VTAIL.n238 VTAIL.n228 8.92171
R769 VTAIL.n272 VTAIL.n271 8.92171
R770 VTAIL.n287 VTAIL.n206 8.92171
R771 VTAIL.n687 VTAIL.n606 8.92171
R772 VTAIL.n672 VTAIL.n671 8.92171
R773 VTAIL.n639 VTAIL.n629 8.92171
R774 VTAIL.n587 VTAIL.n506 8.92171
R775 VTAIL.n572 VTAIL.n571 8.92171
R776 VTAIL.n539 VTAIL.n529 8.92171
R777 VTAIL.n487 VTAIL.n406 8.92171
R778 VTAIL.n472 VTAIL.n471 8.92171
R779 VTAIL.n439 VTAIL.n429 8.92171
R780 VTAIL.n387 VTAIL.n306 8.92171
R781 VTAIL.n372 VTAIL.n371 8.92171
R782 VTAIL.n339 VTAIL.n329 8.92171
R783 VTAIL.n737 VTAIL.n730 8.14595
R784 VTAIL.n775 VTAIL.n712 8.14595
R785 VTAIL.n784 VTAIL.n783 8.14595
R786 VTAIL.n37 VTAIL.n30 8.14595
R787 VTAIL.n75 VTAIL.n12 8.14595
R788 VTAIL.n84 VTAIL.n83 8.14595
R789 VTAIL.n137 VTAIL.n130 8.14595
R790 VTAIL.n175 VTAIL.n112 8.14595
R791 VTAIL.n184 VTAIL.n183 8.14595
R792 VTAIL.n237 VTAIL.n230 8.14595
R793 VTAIL.n275 VTAIL.n212 8.14595
R794 VTAIL.n284 VTAIL.n283 8.14595
R795 VTAIL.n684 VTAIL.n683 8.14595
R796 VTAIL.n675 VTAIL.n612 8.14595
R797 VTAIL.n638 VTAIL.n631 8.14595
R798 VTAIL.n584 VTAIL.n583 8.14595
R799 VTAIL.n575 VTAIL.n512 8.14595
R800 VTAIL.n538 VTAIL.n531 8.14595
R801 VTAIL.n484 VTAIL.n483 8.14595
R802 VTAIL.n475 VTAIL.n412 8.14595
R803 VTAIL.n438 VTAIL.n431 8.14595
R804 VTAIL.n384 VTAIL.n383 8.14595
R805 VTAIL.n375 VTAIL.n312 8.14595
R806 VTAIL.n338 VTAIL.n331 8.14595
R807 VTAIL.n734 VTAIL.n733 7.3702
R808 VTAIL.n776 VTAIL.n710 7.3702
R809 VTAIL.n780 VTAIL.n708 7.3702
R810 VTAIL.n34 VTAIL.n33 7.3702
R811 VTAIL.n76 VTAIL.n10 7.3702
R812 VTAIL.n80 VTAIL.n8 7.3702
R813 VTAIL.n134 VTAIL.n133 7.3702
R814 VTAIL.n176 VTAIL.n110 7.3702
R815 VTAIL.n180 VTAIL.n108 7.3702
R816 VTAIL.n234 VTAIL.n233 7.3702
R817 VTAIL.n276 VTAIL.n210 7.3702
R818 VTAIL.n280 VTAIL.n208 7.3702
R819 VTAIL.n680 VTAIL.n608 7.3702
R820 VTAIL.n676 VTAIL.n610 7.3702
R821 VTAIL.n635 VTAIL.n634 7.3702
R822 VTAIL.n580 VTAIL.n508 7.3702
R823 VTAIL.n576 VTAIL.n510 7.3702
R824 VTAIL.n535 VTAIL.n534 7.3702
R825 VTAIL.n480 VTAIL.n408 7.3702
R826 VTAIL.n476 VTAIL.n410 7.3702
R827 VTAIL.n435 VTAIL.n434 7.3702
R828 VTAIL.n380 VTAIL.n308 7.3702
R829 VTAIL.n376 VTAIL.n310 7.3702
R830 VTAIL.n335 VTAIL.n334 7.3702
R831 VTAIL.n779 VTAIL.n710 6.59444
R832 VTAIL.n780 VTAIL.n779 6.59444
R833 VTAIL.n79 VTAIL.n10 6.59444
R834 VTAIL.n80 VTAIL.n79 6.59444
R835 VTAIL.n179 VTAIL.n110 6.59444
R836 VTAIL.n180 VTAIL.n179 6.59444
R837 VTAIL.n279 VTAIL.n210 6.59444
R838 VTAIL.n280 VTAIL.n279 6.59444
R839 VTAIL.n680 VTAIL.n679 6.59444
R840 VTAIL.n679 VTAIL.n610 6.59444
R841 VTAIL.n580 VTAIL.n579 6.59444
R842 VTAIL.n579 VTAIL.n510 6.59444
R843 VTAIL.n480 VTAIL.n479 6.59444
R844 VTAIL.n479 VTAIL.n410 6.59444
R845 VTAIL.n380 VTAIL.n379 6.59444
R846 VTAIL.n379 VTAIL.n310 6.59444
R847 VTAIL.n734 VTAIL.n730 5.81868
R848 VTAIL.n776 VTAIL.n775 5.81868
R849 VTAIL.n783 VTAIL.n708 5.81868
R850 VTAIL.n34 VTAIL.n30 5.81868
R851 VTAIL.n76 VTAIL.n75 5.81868
R852 VTAIL.n83 VTAIL.n8 5.81868
R853 VTAIL.n134 VTAIL.n130 5.81868
R854 VTAIL.n176 VTAIL.n175 5.81868
R855 VTAIL.n183 VTAIL.n108 5.81868
R856 VTAIL.n234 VTAIL.n230 5.81868
R857 VTAIL.n276 VTAIL.n275 5.81868
R858 VTAIL.n283 VTAIL.n208 5.81868
R859 VTAIL.n683 VTAIL.n608 5.81868
R860 VTAIL.n676 VTAIL.n675 5.81868
R861 VTAIL.n635 VTAIL.n631 5.81868
R862 VTAIL.n583 VTAIL.n508 5.81868
R863 VTAIL.n576 VTAIL.n575 5.81868
R864 VTAIL.n535 VTAIL.n531 5.81868
R865 VTAIL.n483 VTAIL.n408 5.81868
R866 VTAIL.n476 VTAIL.n475 5.81868
R867 VTAIL.n435 VTAIL.n431 5.81868
R868 VTAIL.n383 VTAIL.n308 5.81868
R869 VTAIL.n376 VTAIL.n375 5.81868
R870 VTAIL.n335 VTAIL.n331 5.81868
R871 VTAIL.n738 VTAIL.n737 5.04292
R872 VTAIL.n772 VTAIL.n712 5.04292
R873 VTAIL.n784 VTAIL.n706 5.04292
R874 VTAIL.n38 VTAIL.n37 5.04292
R875 VTAIL.n72 VTAIL.n12 5.04292
R876 VTAIL.n84 VTAIL.n6 5.04292
R877 VTAIL.n138 VTAIL.n137 5.04292
R878 VTAIL.n172 VTAIL.n112 5.04292
R879 VTAIL.n184 VTAIL.n106 5.04292
R880 VTAIL.n238 VTAIL.n237 5.04292
R881 VTAIL.n272 VTAIL.n212 5.04292
R882 VTAIL.n284 VTAIL.n206 5.04292
R883 VTAIL.n684 VTAIL.n606 5.04292
R884 VTAIL.n672 VTAIL.n612 5.04292
R885 VTAIL.n639 VTAIL.n638 5.04292
R886 VTAIL.n584 VTAIL.n506 5.04292
R887 VTAIL.n572 VTAIL.n512 5.04292
R888 VTAIL.n539 VTAIL.n538 5.04292
R889 VTAIL.n484 VTAIL.n406 5.04292
R890 VTAIL.n472 VTAIL.n412 5.04292
R891 VTAIL.n439 VTAIL.n438 5.04292
R892 VTAIL.n384 VTAIL.n306 5.04292
R893 VTAIL.n372 VTAIL.n312 5.04292
R894 VTAIL.n339 VTAIL.n338 5.04292
R895 VTAIL.n741 VTAIL.n728 4.26717
R896 VTAIL.n771 VTAIL.n714 4.26717
R897 VTAIL.n788 VTAIL.n787 4.26717
R898 VTAIL.n41 VTAIL.n28 4.26717
R899 VTAIL.n71 VTAIL.n14 4.26717
R900 VTAIL.n88 VTAIL.n87 4.26717
R901 VTAIL.n141 VTAIL.n128 4.26717
R902 VTAIL.n171 VTAIL.n114 4.26717
R903 VTAIL.n188 VTAIL.n187 4.26717
R904 VTAIL.n241 VTAIL.n228 4.26717
R905 VTAIL.n271 VTAIL.n214 4.26717
R906 VTAIL.n288 VTAIL.n287 4.26717
R907 VTAIL.n688 VTAIL.n687 4.26717
R908 VTAIL.n671 VTAIL.n614 4.26717
R909 VTAIL.n642 VTAIL.n629 4.26717
R910 VTAIL.n588 VTAIL.n587 4.26717
R911 VTAIL.n571 VTAIL.n514 4.26717
R912 VTAIL.n542 VTAIL.n529 4.26717
R913 VTAIL.n488 VTAIL.n487 4.26717
R914 VTAIL.n471 VTAIL.n414 4.26717
R915 VTAIL.n442 VTAIL.n429 4.26717
R916 VTAIL.n388 VTAIL.n387 4.26717
R917 VTAIL.n371 VTAIL.n314 4.26717
R918 VTAIL.n342 VTAIL.n329 4.26717
R919 VTAIL.n742 VTAIL.n726 3.49141
R920 VTAIL.n768 VTAIL.n767 3.49141
R921 VTAIL.n791 VTAIL.n704 3.49141
R922 VTAIL.n42 VTAIL.n26 3.49141
R923 VTAIL.n68 VTAIL.n67 3.49141
R924 VTAIL.n91 VTAIL.n4 3.49141
R925 VTAIL.n142 VTAIL.n126 3.49141
R926 VTAIL.n168 VTAIL.n167 3.49141
R927 VTAIL.n191 VTAIL.n104 3.49141
R928 VTAIL.n242 VTAIL.n226 3.49141
R929 VTAIL.n268 VTAIL.n267 3.49141
R930 VTAIL.n291 VTAIL.n204 3.49141
R931 VTAIL.n691 VTAIL.n604 3.49141
R932 VTAIL.n668 VTAIL.n667 3.49141
R933 VTAIL.n643 VTAIL.n627 3.49141
R934 VTAIL.n591 VTAIL.n504 3.49141
R935 VTAIL.n568 VTAIL.n567 3.49141
R936 VTAIL.n543 VTAIL.n527 3.49141
R937 VTAIL.n491 VTAIL.n404 3.49141
R938 VTAIL.n468 VTAIL.n467 3.49141
R939 VTAIL.n443 VTAIL.n427 3.49141
R940 VTAIL.n391 VTAIL.n304 3.49141
R941 VTAIL.n368 VTAIL.n367 3.49141
R942 VTAIL.n343 VTAIL.n327 3.49141
R943 VTAIL.n746 VTAIL.n745 2.71565
R944 VTAIL.n764 VTAIL.n716 2.71565
R945 VTAIL.n792 VTAIL.n702 2.71565
R946 VTAIL.n46 VTAIL.n45 2.71565
R947 VTAIL.n64 VTAIL.n16 2.71565
R948 VTAIL.n92 VTAIL.n2 2.71565
R949 VTAIL.n146 VTAIL.n145 2.71565
R950 VTAIL.n164 VTAIL.n116 2.71565
R951 VTAIL.n192 VTAIL.n102 2.71565
R952 VTAIL.n246 VTAIL.n245 2.71565
R953 VTAIL.n264 VTAIL.n216 2.71565
R954 VTAIL.n292 VTAIL.n202 2.71565
R955 VTAIL.n692 VTAIL.n602 2.71565
R956 VTAIL.n664 VTAIL.n616 2.71565
R957 VTAIL.n647 VTAIL.n646 2.71565
R958 VTAIL.n592 VTAIL.n502 2.71565
R959 VTAIL.n564 VTAIL.n516 2.71565
R960 VTAIL.n547 VTAIL.n546 2.71565
R961 VTAIL.n492 VTAIL.n402 2.71565
R962 VTAIL.n464 VTAIL.n416 2.71565
R963 VTAIL.n447 VTAIL.n446 2.71565
R964 VTAIL.n392 VTAIL.n302 2.71565
R965 VTAIL.n364 VTAIL.n316 2.71565
R966 VTAIL.n347 VTAIL.n346 2.71565
R967 VTAIL.n735 VTAIL.n731 2.41282
R968 VTAIL.n35 VTAIL.n31 2.41282
R969 VTAIL.n135 VTAIL.n131 2.41282
R970 VTAIL.n235 VTAIL.n231 2.41282
R971 VTAIL.n636 VTAIL.n632 2.41282
R972 VTAIL.n536 VTAIL.n532 2.41282
R973 VTAIL.n436 VTAIL.n432 2.41282
R974 VTAIL.n336 VTAIL.n332 2.41282
R975 VTAIL.n750 VTAIL.n724 1.93989
R976 VTAIL.n763 VTAIL.n718 1.93989
R977 VTAIL.n796 VTAIL.n795 1.93989
R978 VTAIL.n50 VTAIL.n24 1.93989
R979 VTAIL.n63 VTAIL.n18 1.93989
R980 VTAIL.n96 VTAIL.n95 1.93989
R981 VTAIL.n150 VTAIL.n124 1.93989
R982 VTAIL.n163 VTAIL.n118 1.93989
R983 VTAIL.n196 VTAIL.n195 1.93989
R984 VTAIL.n250 VTAIL.n224 1.93989
R985 VTAIL.n263 VTAIL.n218 1.93989
R986 VTAIL.n296 VTAIL.n295 1.93989
R987 VTAIL.n696 VTAIL.n695 1.93989
R988 VTAIL.n663 VTAIL.n618 1.93989
R989 VTAIL.n650 VTAIL.n624 1.93989
R990 VTAIL.n596 VTAIL.n595 1.93989
R991 VTAIL.n563 VTAIL.n518 1.93989
R992 VTAIL.n550 VTAIL.n524 1.93989
R993 VTAIL.n496 VTAIL.n495 1.93989
R994 VTAIL.n463 VTAIL.n418 1.93989
R995 VTAIL.n450 VTAIL.n424 1.93989
R996 VTAIL.n396 VTAIL.n395 1.93989
R997 VTAIL.n363 VTAIL.n318 1.93989
R998 VTAIL.n350 VTAIL.n324 1.93989
R999 VTAIL.n499 VTAIL.n399 1.90567
R1000 VTAIL.n699 VTAIL.n599 1.90567
R1001 VTAIL.n299 VTAIL.n199 1.90567
R1002 VTAIL.n751 VTAIL.n722 1.16414
R1003 VTAIL.n760 VTAIL.n759 1.16414
R1004 VTAIL.n798 VTAIL.n700 1.16414
R1005 VTAIL.n51 VTAIL.n22 1.16414
R1006 VTAIL.n60 VTAIL.n59 1.16414
R1007 VTAIL.n98 VTAIL.n0 1.16414
R1008 VTAIL.n151 VTAIL.n122 1.16414
R1009 VTAIL.n160 VTAIL.n159 1.16414
R1010 VTAIL.n198 VTAIL.n100 1.16414
R1011 VTAIL.n251 VTAIL.n222 1.16414
R1012 VTAIL.n260 VTAIL.n259 1.16414
R1013 VTAIL.n298 VTAIL.n200 1.16414
R1014 VTAIL.n698 VTAIL.n600 1.16414
R1015 VTAIL.n660 VTAIL.n659 1.16414
R1016 VTAIL.n651 VTAIL.n622 1.16414
R1017 VTAIL.n598 VTAIL.n500 1.16414
R1018 VTAIL.n560 VTAIL.n559 1.16414
R1019 VTAIL.n551 VTAIL.n522 1.16414
R1020 VTAIL.n498 VTAIL.n400 1.16414
R1021 VTAIL.n460 VTAIL.n459 1.16414
R1022 VTAIL.n451 VTAIL.n422 1.16414
R1023 VTAIL.n398 VTAIL.n300 1.16414
R1024 VTAIL.n360 VTAIL.n359 1.16414
R1025 VTAIL.n351 VTAIL.n322 1.16414
R1026 VTAIL VTAIL.n99 1.01128
R1027 VTAIL VTAIL.n799 0.894897
R1028 VTAIL.n599 VTAIL.n499 0.470328
R1029 VTAIL.n199 VTAIL.n99 0.470328
R1030 VTAIL.n755 VTAIL.n754 0.388379
R1031 VTAIL.n756 VTAIL.n720 0.388379
R1032 VTAIL.n55 VTAIL.n54 0.388379
R1033 VTAIL.n56 VTAIL.n20 0.388379
R1034 VTAIL.n155 VTAIL.n154 0.388379
R1035 VTAIL.n156 VTAIL.n120 0.388379
R1036 VTAIL.n255 VTAIL.n254 0.388379
R1037 VTAIL.n256 VTAIL.n220 0.388379
R1038 VTAIL.n656 VTAIL.n620 0.388379
R1039 VTAIL.n655 VTAIL.n654 0.388379
R1040 VTAIL.n556 VTAIL.n520 0.388379
R1041 VTAIL.n555 VTAIL.n554 0.388379
R1042 VTAIL.n456 VTAIL.n420 0.388379
R1043 VTAIL.n455 VTAIL.n454 0.388379
R1044 VTAIL.n356 VTAIL.n320 0.388379
R1045 VTAIL.n355 VTAIL.n354 0.388379
R1046 VTAIL.n736 VTAIL.n735 0.155672
R1047 VTAIL.n736 VTAIL.n727 0.155672
R1048 VTAIL.n743 VTAIL.n727 0.155672
R1049 VTAIL.n744 VTAIL.n743 0.155672
R1050 VTAIL.n744 VTAIL.n723 0.155672
R1051 VTAIL.n752 VTAIL.n723 0.155672
R1052 VTAIL.n753 VTAIL.n752 0.155672
R1053 VTAIL.n753 VTAIL.n719 0.155672
R1054 VTAIL.n761 VTAIL.n719 0.155672
R1055 VTAIL.n762 VTAIL.n761 0.155672
R1056 VTAIL.n762 VTAIL.n715 0.155672
R1057 VTAIL.n769 VTAIL.n715 0.155672
R1058 VTAIL.n770 VTAIL.n769 0.155672
R1059 VTAIL.n770 VTAIL.n711 0.155672
R1060 VTAIL.n777 VTAIL.n711 0.155672
R1061 VTAIL.n778 VTAIL.n777 0.155672
R1062 VTAIL.n778 VTAIL.n707 0.155672
R1063 VTAIL.n785 VTAIL.n707 0.155672
R1064 VTAIL.n786 VTAIL.n785 0.155672
R1065 VTAIL.n786 VTAIL.n703 0.155672
R1066 VTAIL.n793 VTAIL.n703 0.155672
R1067 VTAIL.n794 VTAIL.n793 0.155672
R1068 VTAIL.n36 VTAIL.n35 0.155672
R1069 VTAIL.n36 VTAIL.n27 0.155672
R1070 VTAIL.n43 VTAIL.n27 0.155672
R1071 VTAIL.n44 VTAIL.n43 0.155672
R1072 VTAIL.n44 VTAIL.n23 0.155672
R1073 VTAIL.n52 VTAIL.n23 0.155672
R1074 VTAIL.n53 VTAIL.n52 0.155672
R1075 VTAIL.n53 VTAIL.n19 0.155672
R1076 VTAIL.n61 VTAIL.n19 0.155672
R1077 VTAIL.n62 VTAIL.n61 0.155672
R1078 VTAIL.n62 VTAIL.n15 0.155672
R1079 VTAIL.n69 VTAIL.n15 0.155672
R1080 VTAIL.n70 VTAIL.n69 0.155672
R1081 VTAIL.n70 VTAIL.n11 0.155672
R1082 VTAIL.n77 VTAIL.n11 0.155672
R1083 VTAIL.n78 VTAIL.n77 0.155672
R1084 VTAIL.n78 VTAIL.n7 0.155672
R1085 VTAIL.n85 VTAIL.n7 0.155672
R1086 VTAIL.n86 VTAIL.n85 0.155672
R1087 VTAIL.n86 VTAIL.n3 0.155672
R1088 VTAIL.n93 VTAIL.n3 0.155672
R1089 VTAIL.n94 VTAIL.n93 0.155672
R1090 VTAIL.n136 VTAIL.n135 0.155672
R1091 VTAIL.n136 VTAIL.n127 0.155672
R1092 VTAIL.n143 VTAIL.n127 0.155672
R1093 VTAIL.n144 VTAIL.n143 0.155672
R1094 VTAIL.n144 VTAIL.n123 0.155672
R1095 VTAIL.n152 VTAIL.n123 0.155672
R1096 VTAIL.n153 VTAIL.n152 0.155672
R1097 VTAIL.n153 VTAIL.n119 0.155672
R1098 VTAIL.n161 VTAIL.n119 0.155672
R1099 VTAIL.n162 VTAIL.n161 0.155672
R1100 VTAIL.n162 VTAIL.n115 0.155672
R1101 VTAIL.n169 VTAIL.n115 0.155672
R1102 VTAIL.n170 VTAIL.n169 0.155672
R1103 VTAIL.n170 VTAIL.n111 0.155672
R1104 VTAIL.n177 VTAIL.n111 0.155672
R1105 VTAIL.n178 VTAIL.n177 0.155672
R1106 VTAIL.n178 VTAIL.n107 0.155672
R1107 VTAIL.n185 VTAIL.n107 0.155672
R1108 VTAIL.n186 VTAIL.n185 0.155672
R1109 VTAIL.n186 VTAIL.n103 0.155672
R1110 VTAIL.n193 VTAIL.n103 0.155672
R1111 VTAIL.n194 VTAIL.n193 0.155672
R1112 VTAIL.n236 VTAIL.n235 0.155672
R1113 VTAIL.n236 VTAIL.n227 0.155672
R1114 VTAIL.n243 VTAIL.n227 0.155672
R1115 VTAIL.n244 VTAIL.n243 0.155672
R1116 VTAIL.n244 VTAIL.n223 0.155672
R1117 VTAIL.n252 VTAIL.n223 0.155672
R1118 VTAIL.n253 VTAIL.n252 0.155672
R1119 VTAIL.n253 VTAIL.n219 0.155672
R1120 VTAIL.n261 VTAIL.n219 0.155672
R1121 VTAIL.n262 VTAIL.n261 0.155672
R1122 VTAIL.n262 VTAIL.n215 0.155672
R1123 VTAIL.n269 VTAIL.n215 0.155672
R1124 VTAIL.n270 VTAIL.n269 0.155672
R1125 VTAIL.n270 VTAIL.n211 0.155672
R1126 VTAIL.n277 VTAIL.n211 0.155672
R1127 VTAIL.n278 VTAIL.n277 0.155672
R1128 VTAIL.n278 VTAIL.n207 0.155672
R1129 VTAIL.n285 VTAIL.n207 0.155672
R1130 VTAIL.n286 VTAIL.n285 0.155672
R1131 VTAIL.n286 VTAIL.n203 0.155672
R1132 VTAIL.n293 VTAIL.n203 0.155672
R1133 VTAIL.n294 VTAIL.n293 0.155672
R1134 VTAIL.n694 VTAIL.n693 0.155672
R1135 VTAIL.n693 VTAIL.n603 0.155672
R1136 VTAIL.n686 VTAIL.n603 0.155672
R1137 VTAIL.n686 VTAIL.n685 0.155672
R1138 VTAIL.n685 VTAIL.n607 0.155672
R1139 VTAIL.n678 VTAIL.n607 0.155672
R1140 VTAIL.n678 VTAIL.n677 0.155672
R1141 VTAIL.n677 VTAIL.n611 0.155672
R1142 VTAIL.n670 VTAIL.n611 0.155672
R1143 VTAIL.n670 VTAIL.n669 0.155672
R1144 VTAIL.n669 VTAIL.n615 0.155672
R1145 VTAIL.n662 VTAIL.n615 0.155672
R1146 VTAIL.n662 VTAIL.n661 0.155672
R1147 VTAIL.n661 VTAIL.n619 0.155672
R1148 VTAIL.n653 VTAIL.n619 0.155672
R1149 VTAIL.n653 VTAIL.n652 0.155672
R1150 VTAIL.n652 VTAIL.n623 0.155672
R1151 VTAIL.n645 VTAIL.n623 0.155672
R1152 VTAIL.n645 VTAIL.n644 0.155672
R1153 VTAIL.n644 VTAIL.n628 0.155672
R1154 VTAIL.n637 VTAIL.n628 0.155672
R1155 VTAIL.n637 VTAIL.n636 0.155672
R1156 VTAIL.n594 VTAIL.n593 0.155672
R1157 VTAIL.n593 VTAIL.n503 0.155672
R1158 VTAIL.n586 VTAIL.n503 0.155672
R1159 VTAIL.n586 VTAIL.n585 0.155672
R1160 VTAIL.n585 VTAIL.n507 0.155672
R1161 VTAIL.n578 VTAIL.n507 0.155672
R1162 VTAIL.n578 VTAIL.n577 0.155672
R1163 VTAIL.n577 VTAIL.n511 0.155672
R1164 VTAIL.n570 VTAIL.n511 0.155672
R1165 VTAIL.n570 VTAIL.n569 0.155672
R1166 VTAIL.n569 VTAIL.n515 0.155672
R1167 VTAIL.n562 VTAIL.n515 0.155672
R1168 VTAIL.n562 VTAIL.n561 0.155672
R1169 VTAIL.n561 VTAIL.n519 0.155672
R1170 VTAIL.n553 VTAIL.n519 0.155672
R1171 VTAIL.n553 VTAIL.n552 0.155672
R1172 VTAIL.n552 VTAIL.n523 0.155672
R1173 VTAIL.n545 VTAIL.n523 0.155672
R1174 VTAIL.n545 VTAIL.n544 0.155672
R1175 VTAIL.n544 VTAIL.n528 0.155672
R1176 VTAIL.n537 VTAIL.n528 0.155672
R1177 VTAIL.n537 VTAIL.n536 0.155672
R1178 VTAIL.n494 VTAIL.n493 0.155672
R1179 VTAIL.n493 VTAIL.n403 0.155672
R1180 VTAIL.n486 VTAIL.n403 0.155672
R1181 VTAIL.n486 VTAIL.n485 0.155672
R1182 VTAIL.n485 VTAIL.n407 0.155672
R1183 VTAIL.n478 VTAIL.n407 0.155672
R1184 VTAIL.n478 VTAIL.n477 0.155672
R1185 VTAIL.n477 VTAIL.n411 0.155672
R1186 VTAIL.n470 VTAIL.n411 0.155672
R1187 VTAIL.n470 VTAIL.n469 0.155672
R1188 VTAIL.n469 VTAIL.n415 0.155672
R1189 VTAIL.n462 VTAIL.n415 0.155672
R1190 VTAIL.n462 VTAIL.n461 0.155672
R1191 VTAIL.n461 VTAIL.n419 0.155672
R1192 VTAIL.n453 VTAIL.n419 0.155672
R1193 VTAIL.n453 VTAIL.n452 0.155672
R1194 VTAIL.n452 VTAIL.n423 0.155672
R1195 VTAIL.n445 VTAIL.n423 0.155672
R1196 VTAIL.n445 VTAIL.n444 0.155672
R1197 VTAIL.n444 VTAIL.n428 0.155672
R1198 VTAIL.n437 VTAIL.n428 0.155672
R1199 VTAIL.n437 VTAIL.n436 0.155672
R1200 VTAIL.n394 VTAIL.n393 0.155672
R1201 VTAIL.n393 VTAIL.n303 0.155672
R1202 VTAIL.n386 VTAIL.n303 0.155672
R1203 VTAIL.n386 VTAIL.n385 0.155672
R1204 VTAIL.n385 VTAIL.n307 0.155672
R1205 VTAIL.n378 VTAIL.n307 0.155672
R1206 VTAIL.n378 VTAIL.n377 0.155672
R1207 VTAIL.n377 VTAIL.n311 0.155672
R1208 VTAIL.n370 VTAIL.n311 0.155672
R1209 VTAIL.n370 VTAIL.n369 0.155672
R1210 VTAIL.n369 VTAIL.n315 0.155672
R1211 VTAIL.n362 VTAIL.n315 0.155672
R1212 VTAIL.n362 VTAIL.n361 0.155672
R1213 VTAIL.n361 VTAIL.n319 0.155672
R1214 VTAIL.n353 VTAIL.n319 0.155672
R1215 VTAIL.n353 VTAIL.n352 0.155672
R1216 VTAIL.n352 VTAIL.n323 0.155672
R1217 VTAIL.n345 VTAIL.n323 0.155672
R1218 VTAIL.n345 VTAIL.n344 0.155672
R1219 VTAIL.n344 VTAIL.n328 0.155672
R1220 VTAIL.n337 VTAIL.n328 0.155672
R1221 VTAIL.n337 VTAIL.n336 0.155672
R1222 VP.n3 VP.t3 269.659
R1223 VP.n3 VP.t0 269.221
R1224 VP.n5 VP.t2 232.028
R1225 VP.n13 VP.t1 232.028
R1226 VP.n5 VP.n4 180.531
R1227 VP.n14 VP.n13 180.531
R1228 VP.n12 VP.n0 161.3
R1229 VP.n11 VP.n10 161.3
R1230 VP.n9 VP.n1 161.3
R1231 VP.n8 VP.n7 161.3
R1232 VP.n6 VP.n2 161.3
R1233 VP.n4 VP.n3 57.8357
R1234 VP.n7 VP.n1 40.4106
R1235 VP.n11 VP.n1 40.4106
R1236 VP.n7 VP.n6 24.3439
R1237 VP.n12 VP.n11 24.3439
R1238 VP.n6 VP.n5 5.11262
R1239 VP.n13 VP.n12 5.11262
R1240 VP.n4 VP.n2 0.189894
R1241 VP.n8 VP.n2 0.189894
R1242 VP.n9 VP.n8 0.189894
R1243 VP.n10 VP.n9 0.189894
R1244 VP.n10 VP.n0 0.189894
R1245 VP.n14 VP.n0 0.189894
R1246 VP VP.n14 0.0516364
R1247 VDD1 VDD1.n1 118.163
R1248 VDD1 VDD1.n0 72.6625
R1249 VDD1.n0 VDD1.t0 1.79636
R1250 VDD1.n0 VDD1.t3 1.79636
R1251 VDD1.n1 VDD1.t1 1.79636
R1252 VDD1.n1 VDD1.t2 1.79636
R1253 B.n428 B.n427 585
R1254 B.n426 B.n113 585
R1255 B.n425 B.n424 585
R1256 B.n423 B.n114 585
R1257 B.n422 B.n421 585
R1258 B.n420 B.n115 585
R1259 B.n419 B.n418 585
R1260 B.n417 B.n116 585
R1261 B.n416 B.n415 585
R1262 B.n414 B.n117 585
R1263 B.n413 B.n412 585
R1264 B.n411 B.n118 585
R1265 B.n410 B.n409 585
R1266 B.n408 B.n119 585
R1267 B.n407 B.n406 585
R1268 B.n405 B.n120 585
R1269 B.n404 B.n403 585
R1270 B.n402 B.n121 585
R1271 B.n401 B.n400 585
R1272 B.n399 B.n122 585
R1273 B.n398 B.n397 585
R1274 B.n396 B.n123 585
R1275 B.n395 B.n394 585
R1276 B.n393 B.n124 585
R1277 B.n392 B.n391 585
R1278 B.n390 B.n125 585
R1279 B.n389 B.n388 585
R1280 B.n387 B.n126 585
R1281 B.n386 B.n385 585
R1282 B.n384 B.n127 585
R1283 B.n383 B.n382 585
R1284 B.n381 B.n128 585
R1285 B.n380 B.n379 585
R1286 B.n378 B.n129 585
R1287 B.n377 B.n376 585
R1288 B.n375 B.n130 585
R1289 B.n374 B.n373 585
R1290 B.n372 B.n131 585
R1291 B.n371 B.n370 585
R1292 B.n369 B.n132 585
R1293 B.n368 B.n367 585
R1294 B.n366 B.n133 585
R1295 B.n365 B.n364 585
R1296 B.n363 B.n134 585
R1297 B.n362 B.n361 585
R1298 B.n360 B.n135 585
R1299 B.n359 B.n358 585
R1300 B.n357 B.n136 585
R1301 B.n356 B.n355 585
R1302 B.n354 B.n137 585
R1303 B.n353 B.n352 585
R1304 B.n351 B.n138 585
R1305 B.n350 B.n349 585
R1306 B.n348 B.n139 585
R1307 B.n347 B.n346 585
R1308 B.n345 B.n140 585
R1309 B.n344 B.n343 585
R1310 B.n342 B.n141 585
R1311 B.n341 B.n340 585
R1312 B.n339 B.n142 585
R1313 B.n338 B.n337 585
R1314 B.n333 B.n143 585
R1315 B.n332 B.n331 585
R1316 B.n330 B.n144 585
R1317 B.n329 B.n328 585
R1318 B.n327 B.n145 585
R1319 B.n326 B.n325 585
R1320 B.n324 B.n146 585
R1321 B.n323 B.n322 585
R1322 B.n320 B.n147 585
R1323 B.n319 B.n318 585
R1324 B.n317 B.n150 585
R1325 B.n316 B.n315 585
R1326 B.n314 B.n151 585
R1327 B.n313 B.n312 585
R1328 B.n311 B.n152 585
R1329 B.n310 B.n309 585
R1330 B.n308 B.n153 585
R1331 B.n307 B.n306 585
R1332 B.n305 B.n154 585
R1333 B.n304 B.n303 585
R1334 B.n302 B.n155 585
R1335 B.n301 B.n300 585
R1336 B.n299 B.n156 585
R1337 B.n298 B.n297 585
R1338 B.n296 B.n157 585
R1339 B.n295 B.n294 585
R1340 B.n293 B.n158 585
R1341 B.n292 B.n291 585
R1342 B.n290 B.n159 585
R1343 B.n289 B.n288 585
R1344 B.n287 B.n160 585
R1345 B.n286 B.n285 585
R1346 B.n284 B.n161 585
R1347 B.n283 B.n282 585
R1348 B.n281 B.n162 585
R1349 B.n280 B.n279 585
R1350 B.n278 B.n163 585
R1351 B.n277 B.n276 585
R1352 B.n275 B.n164 585
R1353 B.n274 B.n273 585
R1354 B.n272 B.n165 585
R1355 B.n271 B.n270 585
R1356 B.n269 B.n166 585
R1357 B.n268 B.n267 585
R1358 B.n266 B.n167 585
R1359 B.n265 B.n264 585
R1360 B.n263 B.n168 585
R1361 B.n262 B.n261 585
R1362 B.n260 B.n169 585
R1363 B.n259 B.n258 585
R1364 B.n257 B.n170 585
R1365 B.n256 B.n255 585
R1366 B.n254 B.n171 585
R1367 B.n253 B.n252 585
R1368 B.n251 B.n172 585
R1369 B.n250 B.n249 585
R1370 B.n248 B.n173 585
R1371 B.n247 B.n246 585
R1372 B.n245 B.n174 585
R1373 B.n244 B.n243 585
R1374 B.n242 B.n175 585
R1375 B.n241 B.n240 585
R1376 B.n239 B.n176 585
R1377 B.n238 B.n237 585
R1378 B.n236 B.n177 585
R1379 B.n235 B.n234 585
R1380 B.n233 B.n178 585
R1381 B.n232 B.n231 585
R1382 B.n429 B.n112 585
R1383 B.n431 B.n430 585
R1384 B.n432 B.n111 585
R1385 B.n434 B.n433 585
R1386 B.n435 B.n110 585
R1387 B.n437 B.n436 585
R1388 B.n438 B.n109 585
R1389 B.n440 B.n439 585
R1390 B.n441 B.n108 585
R1391 B.n443 B.n442 585
R1392 B.n444 B.n107 585
R1393 B.n446 B.n445 585
R1394 B.n447 B.n106 585
R1395 B.n449 B.n448 585
R1396 B.n450 B.n105 585
R1397 B.n452 B.n451 585
R1398 B.n453 B.n104 585
R1399 B.n455 B.n454 585
R1400 B.n456 B.n103 585
R1401 B.n458 B.n457 585
R1402 B.n459 B.n102 585
R1403 B.n461 B.n460 585
R1404 B.n462 B.n101 585
R1405 B.n464 B.n463 585
R1406 B.n465 B.n100 585
R1407 B.n467 B.n466 585
R1408 B.n468 B.n99 585
R1409 B.n470 B.n469 585
R1410 B.n471 B.n98 585
R1411 B.n473 B.n472 585
R1412 B.n474 B.n97 585
R1413 B.n476 B.n475 585
R1414 B.n477 B.n96 585
R1415 B.n479 B.n478 585
R1416 B.n480 B.n95 585
R1417 B.n482 B.n481 585
R1418 B.n483 B.n94 585
R1419 B.n485 B.n484 585
R1420 B.n486 B.n93 585
R1421 B.n488 B.n487 585
R1422 B.n489 B.n92 585
R1423 B.n491 B.n490 585
R1424 B.n492 B.n91 585
R1425 B.n494 B.n493 585
R1426 B.n495 B.n90 585
R1427 B.n497 B.n496 585
R1428 B.n498 B.n89 585
R1429 B.n500 B.n499 585
R1430 B.n501 B.n88 585
R1431 B.n503 B.n502 585
R1432 B.n504 B.n87 585
R1433 B.n506 B.n505 585
R1434 B.n507 B.n86 585
R1435 B.n509 B.n508 585
R1436 B.n510 B.n85 585
R1437 B.n512 B.n511 585
R1438 B.n707 B.n706 585
R1439 B.n705 B.n16 585
R1440 B.n704 B.n703 585
R1441 B.n702 B.n17 585
R1442 B.n701 B.n700 585
R1443 B.n699 B.n18 585
R1444 B.n698 B.n697 585
R1445 B.n696 B.n19 585
R1446 B.n695 B.n694 585
R1447 B.n693 B.n20 585
R1448 B.n692 B.n691 585
R1449 B.n690 B.n21 585
R1450 B.n689 B.n688 585
R1451 B.n687 B.n22 585
R1452 B.n686 B.n685 585
R1453 B.n684 B.n23 585
R1454 B.n683 B.n682 585
R1455 B.n681 B.n24 585
R1456 B.n680 B.n679 585
R1457 B.n678 B.n25 585
R1458 B.n677 B.n676 585
R1459 B.n675 B.n26 585
R1460 B.n674 B.n673 585
R1461 B.n672 B.n27 585
R1462 B.n671 B.n670 585
R1463 B.n669 B.n28 585
R1464 B.n668 B.n667 585
R1465 B.n666 B.n29 585
R1466 B.n665 B.n664 585
R1467 B.n663 B.n30 585
R1468 B.n662 B.n661 585
R1469 B.n660 B.n31 585
R1470 B.n659 B.n658 585
R1471 B.n657 B.n32 585
R1472 B.n656 B.n655 585
R1473 B.n654 B.n33 585
R1474 B.n653 B.n652 585
R1475 B.n651 B.n34 585
R1476 B.n650 B.n649 585
R1477 B.n648 B.n35 585
R1478 B.n647 B.n646 585
R1479 B.n645 B.n36 585
R1480 B.n644 B.n643 585
R1481 B.n642 B.n37 585
R1482 B.n641 B.n640 585
R1483 B.n639 B.n38 585
R1484 B.n638 B.n637 585
R1485 B.n636 B.n39 585
R1486 B.n635 B.n634 585
R1487 B.n633 B.n40 585
R1488 B.n632 B.n631 585
R1489 B.n630 B.n41 585
R1490 B.n629 B.n628 585
R1491 B.n627 B.n42 585
R1492 B.n626 B.n625 585
R1493 B.n624 B.n43 585
R1494 B.n623 B.n622 585
R1495 B.n621 B.n44 585
R1496 B.n620 B.n619 585
R1497 B.n618 B.n45 585
R1498 B.n616 B.n615 585
R1499 B.n614 B.n48 585
R1500 B.n613 B.n612 585
R1501 B.n611 B.n49 585
R1502 B.n610 B.n609 585
R1503 B.n608 B.n50 585
R1504 B.n607 B.n606 585
R1505 B.n605 B.n51 585
R1506 B.n604 B.n603 585
R1507 B.n602 B.n601 585
R1508 B.n600 B.n55 585
R1509 B.n599 B.n598 585
R1510 B.n597 B.n56 585
R1511 B.n596 B.n595 585
R1512 B.n594 B.n57 585
R1513 B.n593 B.n592 585
R1514 B.n591 B.n58 585
R1515 B.n590 B.n589 585
R1516 B.n588 B.n59 585
R1517 B.n587 B.n586 585
R1518 B.n585 B.n60 585
R1519 B.n584 B.n583 585
R1520 B.n582 B.n61 585
R1521 B.n581 B.n580 585
R1522 B.n579 B.n62 585
R1523 B.n578 B.n577 585
R1524 B.n576 B.n63 585
R1525 B.n575 B.n574 585
R1526 B.n573 B.n64 585
R1527 B.n572 B.n571 585
R1528 B.n570 B.n65 585
R1529 B.n569 B.n568 585
R1530 B.n567 B.n66 585
R1531 B.n566 B.n565 585
R1532 B.n564 B.n67 585
R1533 B.n563 B.n562 585
R1534 B.n561 B.n68 585
R1535 B.n560 B.n559 585
R1536 B.n558 B.n69 585
R1537 B.n557 B.n556 585
R1538 B.n555 B.n70 585
R1539 B.n554 B.n553 585
R1540 B.n552 B.n71 585
R1541 B.n551 B.n550 585
R1542 B.n549 B.n72 585
R1543 B.n548 B.n547 585
R1544 B.n546 B.n73 585
R1545 B.n545 B.n544 585
R1546 B.n543 B.n74 585
R1547 B.n542 B.n541 585
R1548 B.n540 B.n75 585
R1549 B.n539 B.n538 585
R1550 B.n537 B.n76 585
R1551 B.n536 B.n535 585
R1552 B.n534 B.n77 585
R1553 B.n533 B.n532 585
R1554 B.n531 B.n78 585
R1555 B.n530 B.n529 585
R1556 B.n528 B.n79 585
R1557 B.n527 B.n526 585
R1558 B.n525 B.n80 585
R1559 B.n524 B.n523 585
R1560 B.n522 B.n81 585
R1561 B.n521 B.n520 585
R1562 B.n519 B.n82 585
R1563 B.n518 B.n517 585
R1564 B.n516 B.n83 585
R1565 B.n515 B.n514 585
R1566 B.n513 B.n84 585
R1567 B.n708 B.n15 585
R1568 B.n710 B.n709 585
R1569 B.n711 B.n14 585
R1570 B.n713 B.n712 585
R1571 B.n714 B.n13 585
R1572 B.n716 B.n715 585
R1573 B.n717 B.n12 585
R1574 B.n719 B.n718 585
R1575 B.n720 B.n11 585
R1576 B.n722 B.n721 585
R1577 B.n723 B.n10 585
R1578 B.n725 B.n724 585
R1579 B.n726 B.n9 585
R1580 B.n728 B.n727 585
R1581 B.n729 B.n8 585
R1582 B.n731 B.n730 585
R1583 B.n732 B.n7 585
R1584 B.n734 B.n733 585
R1585 B.n735 B.n6 585
R1586 B.n737 B.n736 585
R1587 B.n738 B.n5 585
R1588 B.n740 B.n739 585
R1589 B.n741 B.n4 585
R1590 B.n743 B.n742 585
R1591 B.n744 B.n3 585
R1592 B.n746 B.n745 585
R1593 B.n747 B.n0 585
R1594 B.n2 B.n1 585
R1595 B.n193 B.n192 585
R1596 B.n194 B.n191 585
R1597 B.n196 B.n195 585
R1598 B.n197 B.n190 585
R1599 B.n199 B.n198 585
R1600 B.n200 B.n189 585
R1601 B.n202 B.n201 585
R1602 B.n203 B.n188 585
R1603 B.n205 B.n204 585
R1604 B.n206 B.n187 585
R1605 B.n208 B.n207 585
R1606 B.n209 B.n186 585
R1607 B.n211 B.n210 585
R1608 B.n212 B.n185 585
R1609 B.n214 B.n213 585
R1610 B.n215 B.n184 585
R1611 B.n217 B.n216 585
R1612 B.n218 B.n183 585
R1613 B.n220 B.n219 585
R1614 B.n221 B.n182 585
R1615 B.n223 B.n222 585
R1616 B.n224 B.n181 585
R1617 B.n226 B.n225 585
R1618 B.n227 B.n180 585
R1619 B.n229 B.n228 585
R1620 B.n230 B.n179 585
R1621 B.n334 B.t7 528.235
R1622 B.n52 B.t11 528.235
R1623 B.n148 B.t1 528.235
R1624 B.n46 B.t5 528.235
R1625 B.n232 B.n179 492.5
R1626 B.n429 B.n428 492.5
R1627 B.n513 B.n512 492.5
R1628 B.n706 B.n15 492.5
R1629 B.n335 B.t8 485.373
R1630 B.n53 B.t10 485.373
R1631 B.n149 B.t2 485.373
R1632 B.n47 B.t4 485.373
R1633 B.n148 B.t0 438.649
R1634 B.n334 B.t6 438.649
R1635 B.n52 B.t9 438.649
R1636 B.n46 B.t3 438.649
R1637 B.n749 B.n748 256.663
R1638 B.n748 B.n747 235.042
R1639 B.n748 B.n2 235.042
R1640 B.n233 B.n232 163.367
R1641 B.n234 B.n233 163.367
R1642 B.n234 B.n177 163.367
R1643 B.n238 B.n177 163.367
R1644 B.n239 B.n238 163.367
R1645 B.n240 B.n239 163.367
R1646 B.n240 B.n175 163.367
R1647 B.n244 B.n175 163.367
R1648 B.n245 B.n244 163.367
R1649 B.n246 B.n245 163.367
R1650 B.n246 B.n173 163.367
R1651 B.n250 B.n173 163.367
R1652 B.n251 B.n250 163.367
R1653 B.n252 B.n251 163.367
R1654 B.n252 B.n171 163.367
R1655 B.n256 B.n171 163.367
R1656 B.n257 B.n256 163.367
R1657 B.n258 B.n257 163.367
R1658 B.n258 B.n169 163.367
R1659 B.n262 B.n169 163.367
R1660 B.n263 B.n262 163.367
R1661 B.n264 B.n263 163.367
R1662 B.n264 B.n167 163.367
R1663 B.n268 B.n167 163.367
R1664 B.n269 B.n268 163.367
R1665 B.n270 B.n269 163.367
R1666 B.n270 B.n165 163.367
R1667 B.n274 B.n165 163.367
R1668 B.n275 B.n274 163.367
R1669 B.n276 B.n275 163.367
R1670 B.n276 B.n163 163.367
R1671 B.n280 B.n163 163.367
R1672 B.n281 B.n280 163.367
R1673 B.n282 B.n281 163.367
R1674 B.n282 B.n161 163.367
R1675 B.n286 B.n161 163.367
R1676 B.n287 B.n286 163.367
R1677 B.n288 B.n287 163.367
R1678 B.n288 B.n159 163.367
R1679 B.n292 B.n159 163.367
R1680 B.n293 B.n292 163.367
R1681 B.n294 B.n293 163.367
R1682 B.n294 B.n157 163.367
R1683 B.n298 B.n157 163.367
R1684 B.n299 B.n298 163.367
R1685 B.n300 B.n299 163.367
R1686 B.n300 B.n155 163.367
R1687 B.n304 B.n155 163.367
R1688 B.n305 B.n304 163.367
R1689 B.n306 B.n305 163.367
R1690 B.n306 B.n153 163.367
R1691 B.n310 B.n153 163.367
R1692 B.n311 B.n310 163.367
R1693 B.n312 B.n311 163.367
R1694 B.n312 B.n151 163.367
R1695 B.n316 B.n151 163.367
R1696 B.n317 B.n316 163.367
R1697 B.n318 B.n317 163.367
R1698 B.n318 B.n147 163.367
R1699 B.n323 B.n147 163.367
R1700 B.n324 B.n323 163.367
R1701 B.n325 B.n324 163.367
R1702 B.n325 B.n145 163.367
R1703 B.n329 B.n145 163.367
R1704 B.n330 B.n329 163.367
R1705 B.n331 B.n330 163.367
R1706 B.n331 B.n143 163.367
R1707 B.n338 B.n143 163.367
R1708 B.n339 B.n338 163.367
R1709 B.n340 B.n339 163.367
R1710 B.n340 B.n141 163.367
R1711 B.n344 B.n141 163.367
R1712 B.n345 B.n344 163.367
R1713 B.n346 B.n345 163.367
R1714 B.n346 B.n139 163.367
R1715 B.n350 B.n139 163.367
R1716 B.n351 B.n350 163.367
R1717 B.n352 B.n351 163.367
R1718 B.n352 B.n137 163.367
R1719 B.n356 B.n137 163.367
R1720 B.n357 B.n356 163.367
R1721 B.n358 B.n357 163.367
R1722 B.n358 B.n135 163.367
R1723 B.n362 B.n135 163.367
R1724 B.n363 B.n362 163.367
R1725 B.n364 B.n363 163.367
R1726 B.n364 B.n133 163.367
R1727 B.n368 B.n133 163.367
R1728 B.n369 B.n368 163.367
R1729 B.n370 B.n369 163.367
R1730 B.n370 B.n131 163.367
R1731 B.n374 B.n131 163.367
R1732 B.n375 B.n374 163.367
R1733 B.n376 B.n375 163.367
R1734 B.n376 B.n129 163.367
R1735 B.n380 B.n129 163.367
R1736 B.n381 B.n380 163.367
R1737 B.n382 B.n381 163.367
R1738 B.n382 B.n127 163.367
R1739 B.n386 B.n127 163.367
R1740 B.n387 B.n386 163.367
R1741 B.n388 B.n387 163.367
R1742 B.n388 B.n125 163.367
R1743 B.n392 B.n125 163.367
R1744 B.n393 B.n392 163.367
R1745 B.n394 B.n393 163.367
R1746 B.n394 B.n123 163.367
R1747 B.n398 B.n123 163.367
R1748 B.n399 B.n398 163.367
R1749 B.n400 B.n399 163.367
R1750 B.n400 B.n121 163.367
R1751 B.n404 B.n121 163.367
R1752 B.n405 B.n404 163.367
R1753 B.n406 B.n405 163.367
R1754 B.n406 B.n119 163.367
R1755 B.n410 B.n119 163.367
R1756 B.n411 B.n410 163.367
R1757 B.n412 B.n411 163.367
R1758 B.n412 B.n117 163.367
R1759 B.n416 B.n117 163.367
R1760 B.n417 B.n416 163.367
R1761 B.n418 B.n417 163.367
R1762 B.n418 B.n115 163.367
R1763 B.n422 B.n115 163.367
R1764 B.n423 B.n422 163.367
R1765 B.n424 B.n423 163.367
R1766 B.n424 B.n113 163.367
R1767 B.n428 B.n113 163.367
R1768 B.n512 B.n85 163.367
R1769 B.n508 B.n85 163.367
R1770 B.n508 B.n507 163.367
R1771 B.n507 B.n506 163.367
R1772 B.n506 B.n87 163.367
R1773 B.n502 B.n87 163.367
R1774 B.n502 B.n501 163.367
R1775 B.n501 B.n500 163.367
R1776 B.n500 B.n89 163.367
R1777 B.n496 B.n89 163.367
R1778 B.n496 B.n495 163.367
R1779 B.n495 B.n494 163.367
R1780 B.n494 B.n91 163.367
R1781 B.n490 B.n91 163.367
R1782 B.n490 B.n489 163.367
R1783 B.n489 B.n488 163.367
R1784 B.n488 B.n93 163.367
R1785 B.n484 B.n93 163.367
R1786 B.n484 B.n483 163.367
R1787 B.n483 B.n482 163.367
R1788 B.n482 B.n95 163.367
R1789 B.n478 B.n95 163.367
R1790 B.n478 B.n477 163.367
R1791 B.n477 B.n476 163.367
R1792 B.n476 B.n97 163.367
R1793 B.n472 B.n97 163.367
R1794 B.n472 B.n471 163.367
R1795 B.n471 B.n470 163.367
R1796 B.n470 B.n99 163.367
R1797 B.n466 B.n99 163.367
R1798 B.n466 B.n465 163.367
R1799 B.n465 B.n464 163.367
R1800 B.n464 B.n101 163.367
R1801 B.n460 B.n101 163.367
R1802 B.n460 B.n459 163.367
R1803 B.n459 B.n458 163.367
R1804 B.n458 B.n103 163.367
R1805 B.n454 B.n103 163.367
R1806 B.n454 B.n453 163.367
R1807 B.n453 B.n452 163.367
R1808 B.n452 B.n105 163.367
R1809 B.n448 B.n105 163.367
R1810 B.n448 B.n447 163.367
R1811 B.n447 B.n446 163.367
R1812 B.n446 B.n107 163.367
R1813 B.n442 B.n107 163.367
R1814 B.n442 B.n441 163.367
R1815 B.n441 B.n440 163.367
R1816 B.n440 B.n109 163.367
R1817 B.n436 B.n109 163.367
R1818 B.n436 B.n435 163.367
R1819 B.n435 B.n434 163.367
R1820 B.n434 B.n111 163.367
R1821 B.n430 B.n111 163.367
R1822 B.n430 B.n429 163.367
R1823 B.n706 B.n705 163.367
R1824 B.n705 B.n704 163.367
R1825 B.n704 B.n17 163.367
R1826 B.n700 B.n17 163.367
R1827 B.n700 B.n699 163.367
R1828 B.n699 B.n698 163.367
R1829 B.n698 B.n19 163.367
R1830 B.n694 B.n19 163.367
R1831 B.n694 B.n693 163.367
R1832 B.n693 B.n692 163.367
R1833 B.n692 B.n21 163.367
R1834 B.n688 B.n21 163.367
R1835 B.n688 B.n687 163.367
R1836 B.n687 B.n686 163.367
R1837 B.n686 B.n23 163.367
R1838 B.n682 B.n23 163.367
R1839 B.n682 B.n681 163.367
R1840 B.n681 B.n680 163.367
R1841 B.n680 B.n25 163.367
R1842 B.n676 B.n25 163.367
R1843 B.n676 B.n675 163.367
R1844 B.n675 B.n674 163.367
R1845 B.n674 B.n27 163.367
R1846 B.n670 B.n27 163.367
R1847 B.n670 B.n669 163.367
R1848 B.n669 B.n668 163.367
R1849 B.n668 B.n29 163.367
R1850 B.n664 B.n29 163.367
R1851 B.n664 B.n663 163.367
R1852 B.n663 B.n662 163.367
R1853 B.n662 B.n31 163.367
R1854 B.n658 B.n31 163.367
R1855 B.n658 B.n657 163.367
R1856 B.n657 B.n656 163.367
R1857 B.n656 B.n33 163.367
R1858 B.n652 B.n33 163.367
R1859 B.n652 B.n651 163.367
R1860 B.n651 B.n650 163.367
R1861 B.n650 B.n35 163.367
R1862 B.n646 B.n35 163.367
R1863 B.n646 B.n645 163.367
R1864 B.n645 B.n644 163.367
R1865 B.n644 B.n37 163.367
R1866 B.n640 B.n37 163.367
R1867 B.n640 B.n639 163.367
R1868 B.n639 B.n638 163.367
R1869 B.n638 B.n39 163.367
R1870 B.n634 B.n39 163.367
R1871 B.n634 B.n633 163.367
R1872 B.n633 B.n632 163.367
R1873 B.n632 B.n41 163.367
R1874 B.n628 B.n41 163.367
R1875 B.n628 B.n627 163.367
R1876 B.n627 B.n626 163.367
R1877 B.n626 B.n43 163.367
R1878 B.n622 B.n43 163.367
R1879 B.n622 B.n621 163.367
R1880 B.n621 B.n620 163.367
R1881 B.n620 B.n45 163.367
R1882 B.n615 B.n45 163.367
R1883 B.n615 B.n614 163.367
R1884 B.n614 B.n613 163.367
R1885 B.n613 B.n49 163.367
R1886 B.n609 B.n49 163.367
R1887 B.n609 B.n608 163.367
R1888 B.n608 B.n607 163.367
R1889 B.n607 B.n51 163.367
R1890 B.n603 B.n51 163.367
R1891 B.n603 B.n602 163.367
R1892 B.n602 B.n55 163.367
R1893 B.n598 B.n55 163.367
R1894 B.n598 B.n597 163.367
R1895 B.n597 B.n596 163.367
R1896 B.n596 B.n57 163.367
R1897 B.n592 B.n57 163.367
R1898 B.n592 B.n591 163.367
R1899 B.n591 B.n590 163.367
R1900 B.n590 B.n59 163.367
R1901 B.n586 B.n59 163.367
R1902 B.n586 B.n585 163.367
R1903 B.n585 B.n584 163.367
R1904 B.n584 B.n61 163.367
R1905 B.n580 B.n61 163.367
R1906 B.n580 B.n579 163.367
R1907 B.n579 B.n578 163.367
R1908 B.n578 B.n63 163.367
R1909 B.n574 B.n63 163.367
R1910 B.n574 B.n573 163.367
R1911 B.n573 B.n572 163.367
R1912 B.n572 B.n65 163.367
R1913 B.n568 B.n65 163.367
R1914 B.n568 B.n567 163.367
R1915 B.n567 B.n566 163.367
R1916 B.n566 B.n67 163.367
R1917 B.n562 B.n67 163.367
R1918 B.n562 B.n561 163.367
R1919 B.n561 B.n560 163.367
R1920 B.n560 B.n69 163.367
R1921 B.n556 B.n69 163.367
R1922 B.n556 B.n555 163.367
R1923 B.n555 B.n554 163.367
R1924 B.n554 B.n71 163.367
R1925 B.n550 B.n71 163.367
R1926 B.n550 B.n549 163.367
R1927 B.n549 B.n548 163.367
R1928 B.n548 B.n73 163.367
R1929 B.n544 B.n73 163.367
R1930 B.n544 B.n543 163.367
R1931 B.n543 B.n542 163.367
R1932 B.n542 B.n75 163.367
R1933 B.n538 B.n75 163.367
R1934 B.n538 B.n537 163.367
R1935 B.n537 B.n536 163.367
R1936 B.n536 B.n77 163.367
R1937 B.n532 B.n77 163.367
R1938 B.n532 B.n531 163.367
R1939 B.n531 B.n530 163.367
R1940 B.n530 B.n79 163.367
R1941 B.n526 B.n79 163.367
R1942 B.n526 B.n525 163.367
R1943 B.n525 B.n524 163.367
R1944 B.n524 B.n81 163.367
R1945 B.n520 B.n81 163.367
R1946 B.n520 B.n519 163.367
R1947 B.n519 B.n518 163.367
R1948 B.n518 B.n83 163.367
R1949 B.n514 B.n83 163.367
R1950 B.n514 B.n513 163.367
R1951 B.n710 B.n15 163.367
R1952 B.n711 B.n710 163.367
R1953 B.n712 B.n711 163.367
R1954 B.n712 B.n13 163.367
R1955 B.n716 B.n13 163.367
R1956 B.n717 B.n716 163.367
R1957 B.n718 B.n717 163.367
R1958 B.n718 B.n11 163.367
R1959 B.n722 B.n11 163.367
R1960 B.n723 B.n722 163.367
R1961 B.n724 B.n723 163.367
R1962 B.n724 B.n9 163.367
R1963 B.n728 B.n9 163.367
R1964 B.n729 B.n728 163.367
R1965 B.n730 B.n729 163.367
R1966 B.n730 B.n7 163.367
R1967 B.n734 B.n7 163.367
R1968 B.n735 B.n734 163.367
R1969 B.n736 B.n735 163.367
R1970 B.n736 B.n5 163.367
R1971 B.n740 B.n5 163.367
R1972 B.n741 B.n740 163.367
R1973 B.n742 B.n741 163.367
R1974 B.n742 B.n3 163.367
R1975 B.n746 B.n3 163.367
R1976 B.n747 B.n746 163.367
R1977 B.n192 B.n2 163.367
R1978 B.n192 B.n191 163.367
R1979 B.n196 B.n191 163.367
R1980 B.n197 B.n196 163.367
R1981 B.n198 B.n197 163.367
R1982 B.n198 B.n189 163.367
R1983 B.n202 B.n189 163.367
R1984 B.n203 B.n202 163.367
R1985 B.n204 B.n203 163.367
R1986 B.n204 B.n187 163.367
R1987 B.n208 B.n187 163.367
R1988 B.n209 B.n208 163.367
R1989 B.n210 B.n209 163.367
R1990 B.n210 B.n185 163.367
R1991 B.n214 B.n185 163.367
R1992 B.n215 B.n214 163.367
R1993 B.n216 B.n215 163.367
R1994 B.n216 B.n183 163.367
R1995 B.n220 B.n183 163.367
R1996 B.n221 B.n220 163.367
R1997 B.n222 B.n221 163.367
R1998 B.n222 B.n181 163.367
R1999 B.n226 B.n181 163.367
R2000 B.n227 B.n226 163.367
R2001 B.n228 B.n227 163.367
R2002 B.n228 B.n179 163.367
R2003 B.n321 B.n149 59.5399
R2004 B.n336 B.n335 59.5399
R2005 B.n54 B.n53 59.5399
R2006 B.n617 B.n47 59.5399
R2007 B.n149 B.n148 42.8611
R2008 B.n335 B.n334 42.8611
R2009 B.n53 B.n52 42.8611
R2010 B.n47 B.n46 42.8611
R2011 B.n708 B.n707 32.0005
R2012 B.n511 B.n84 32.0005
R2013 B.n427 B.n112 32.0005
R2014 B.n231 B.n230 32.0005
R2015 B B.n749 18.0485
R2016 B.n709 B.n708 10.6151
R2017 B.n709 B.n14 10.6151
R2018 B.n713 B.n14 10.6151
R2019 B.n714 B.n713 10.6151
R2020 B.n715 B.n714 10.6151
R2021 B.n715 B.n12 10.6151
R2022 B.n719 B.n12 10.6151
R2023 B.n720 B.n719 10.6151
R2024 B.n721 B.n720 10.6151
R2025 B.n721 B.n10 10.6151
R2026 B.n725 B.n10 10.6151
R2027 B.n726 B.n725 10.6151
R2028 B.n727 B.n726 10.6151
R2029 B.n727 B.n8 10.6151
R2030 B.n731 B.n8 10.6151
R2031 B.n732 B.n731 10.6151
R2032 B.n733 B.n732 10.6151
R2033 B.n733 B.n6 10.6151
R2034 B.n737 B.n6 10.6151
R2035 B.n738 B.n737 10.6151
R2036 B.n739 B.n738 10.6151
R2037 B.n739 B.n4 10.6151
R2038 B.n743 B.n4 10.6151
R2039 B.n744 B.n743 10.6151
R2040 B.n745 B.n744 10.6151
R2041 B.n745 B.n0 10.6151
R2042 B.n707 B.n16 10.6151
R2043 B.n703 B.n16 10.6151
R2044 B.n703 B.n702 10.6151
R2045 B.n702 B.n701 10.6151
R2046 B.n701 B.n18 10.6151
R2047 B.n697 B.n18 10.6151
R2048 B.n697 B.n696 10.6151
R2049 B.n696 B.n695 10.6151
R2050 B.n695 B.n20 10.6151
R2051 B.n691 B.n20 10.6151
R2052 B.n691 B.n690 10.6151
R2053 B.n690 B.n689 10.6151
R2054 B.n689 B.n22 10.6151
R2055 B.n685 B.n22 10.6151
R2056 B.n685 B.n684 10.6151
R2057 B.n684 B.n683 10.6151
R2058 B.n683 B.n24 10.6151
R2059 B.n679 B.n24 10.6151
R2060 B.n679 B.n678 10.6151
R2061 B.n678 B.n677 10.6151
R2062 B.n677 B.n26 10.6151
R2063 B.n673 B.n26 10.6151
R2064 B.n673 B.n672 10.6151
R2065 B.n672 B.n671 10.6151
R2066 B.n671 B.n28 10.6151
R2067 B.n667 B.n28 10.6151
R2068 B.n667 B.n666 10.6151
R2069 B.n666 B.n665 10.6151
R2070 B.n665 B.n30 10.6151
R2071 B.n661 B.n30 10.6151
R2072 B.n661 B.n660 10.6151
R2073 B.n660 B.n659 10.6151
R2074 B.n659 B.n32 10.6151
R2075 B.n655 B.n32 10.6151
R2076 B.n655 B.n654 10.6151
R2077 B.n654 B.n653 10.6151
R2078 B.n653 B.n34 10.6151
R2079 B.n649 B.n34 10.6151
R2080 B.n649 B.n648 10.6151
R2081 B.n648 B.n647 10.6151
R2082 B.n647 B.n36 10.6151
R2083 B.n643 B.n36 10.6151
R2084 B.n643 B.n642 10.6151
R2085 B.n642 B.n641 10.6151
R2086 B.n641 B.n38 10.6151
R2087 B.n637 B.n38 10.6151
R2088 B.n637 B.n636 10.6151
R2089 B.n636 B.n635 10.6151
R2090 B.n635 B.n40 10.6151
R2091 B.n631 B.n40 10.6151
R2092 B.n631 B.n630 10.6151
R2093 B.n630 B.n629 10.6151
R2094 B.n629 B.n42 10.6151
R2095 B.n625 B.n42 10.6151
R2096 B.n625 B.n624 10.6151
R2097 B.n624 B.n623 10.6151
R2098 B.n623 B.n44 10.6151
R2099 B.n619 B.n44 10.6151
R2100 B.n619 B.n618 10.6151
R2101 B.n616 B.n48 10.6151
R2102 B.n612 B.n48 10.6151
R2103 B.n612 B.n611 10.6151
R2104 B.n611 B.n610 10.6151
R2105 B.n610 B.n50 10.6151
R2106 B.n606 B.n50 10.6151
R2107 B.n606 B.n605 10.6151
R2108 B.n605 B.n604 10.6151
R2109 B.n601 B.n600 10.6151
R2110 B.n600 B.n599 10.6151
R2111 B.n599 B.n56 10.6151
R2112 B.n595 B.n56 10.6151
R2113 B.n595 B.n594 10.6151
R2114 B.n594 B.n593 10.6151
R2115 B.n593 B.n58 10.6151
R2116 B.n589 B.n58 10.6151
R2117 B.n589 B.n588 10.6151
R2118 B.n588 B.n587 10.6151
R2119 B.n587 B.n60 10.6151
R2120 B.n583 B.n60 10.6151
R2121 B.n583 B.n582 10.6151
R2122 B.n582 B.n581 10.6151
R2123 B.n581 B.n62 10.6151
R2124 B.n577 B.n62 10.6151
R2125 B.n577 B.n576 10.6151
R2126 B.n576 B.n575 10.6151
R2127 B.n575 B.n64 10.6151
R2128 B.n571 B.n64 10.6151
R2129 B.n571 B.n570 10.6151
R2130 B.n570 B.n569 10.6151
R2131 B.n569 B.n66 10.6151
R2132 B.n565 B.n66 10.6151
R2133 B.n565 B.n564 10.6151
R2134 B.n564 B.n563 10.6151
R2135 B.n563 B.n68 10.6151
R2136 B.n559 B.n68 10.6151
R2137 B.n559 B.n558 10.6151
R2138 B.n558 B.n557 10.6151
R2139 B.n557 B.n70 10.6151
R2140 B.n553 B.n70 10.6151
R2141 B.n553 B.n552 10.6151
R2142 B.n552 B.n551 10.6151
R2143 B.n551 B.n72 10.6151
R2144 B.n547 B.n72 10.6151
R2145 B.n547 B.n546 10.6151
R2146 B.n546 B.n545 10.6151
R2147 B.n545 B.n74 10.6151
R2148 B.n541 B.n74 10.6151
R2149 B.n541 B.n540 10.6151
R2150 B.n540 B.n539 10.6151
R2151 B.n539 B.n76 10.6151
R2152 B.n535 B.n76 10.6151
R2153 B.n535 B.n534 10.6151
R2154 B.n534 B.n533 10.6151
R2155 B.n533 B.n78 10.6151
R2156 B.n529 B.n78 10.6151
R2157 B.n529 B.n528 10.6151
R2158 B.n528 B.n527 10.6151
R2159 B.n527 B.n80 10.6151
R2160 B.n523 B.n80 10.6151
R2161 B.n523 B.n522 10.6151
R2162 B.n522 B.n521 10.6151
R2163 B.n521 B.n82 10.6151
R2164 B.n517 B.n82 10.6151
R2165 B.n517 B.n516 10.6151
R2166 B.n516 B.n515 10.6151
R2167 B.n515 B.n84 10.6151
R2168 B.n511 B.n510 10.6151
R2169 B.n510 B.n509 10.6151
R2170 B.n509 B.n86 10.6151
R2171 B.n505 B.n86 10.6151
R2172 B.n505 B.n504 10.6151
R2173 B.n504 B.n503 10.6151
R2174 B.n503 B.n88 10.6151
R2175 B.n499 B.n88 10.6151
R2176 B.n499 B.n498 10.6151
R2177 B.n498 B.n497 10.6151
R2178 B.n497 B.n90 10.6151
R2179 B.n493 B.n90 10.6151
R2180 B.n493 B.n492 10.6151
R2181 B.n492 B.n491 10.6151
R2182 B.n491 B.n92 10.6151
R2183 B.n487 B.n92 10.6151
R2184 B.n487 B.n486 10.6151
R2185 B.n486 B.n485 10.6151
R2186 B.n485 B.n94 10.6151
R2187 B.n481 B.n94 10.6151
R2188 B.n481 B.n480 10.6151
R2189 B.n480 B.n479 10.6151
R2190 B.n479 B.n96 10.6151
R2191 B.n475 B.n96 10.6151
R2192 B.n475 B.n474 10.6151
R2193 B.n474 B.n473 10.6151
R2194 B.n473 B.n98 10.6151
R2195 B.n469 B.n98 10.6151
R2196 B.n469 B.n468 10.6151
R2197 B.n468 B.n467 10.6151
R2198 B.n467 B.n100 10.6151
R2199 B.n463 B.n100 10.6151
R2200 B.n463 B.n462 10.6151
R2201 B.n462 B.n461 10.6151
R2202 B.n461 B.n102 10.6151
R2203 B.n457 B.n102 10.6151
R2204 B.n457 B.n456 10.6151
R2205 B.n456 B.n455 10.6151
R2206 B.n455 B.n104 10.6151
R2207 B.n451 B.n104 10.6151
R2208 B.n451 B.n450 10.6151
R2209 B.n450 B.n449 10.6151
R2210 B.n449 B.n106 10.6151
R2211 B.n445 B.n106 10.6151
R2212 B.n445 B.n444 10.6151
R2213 B.n444 B.n443 10.6151
R2214 B.n443 B.n108 10.6151
R2215 B.n439 B.n108 10.6151
R2216 B.n439 B.n438 10.6151
R2217 B.n438 B.n437 10.6151
R2218 B.n437 B.n110 10.6151
R2219 B.n433 B.n110 10.6151
R2220 B.n433 B.n432 10.6151
R2221 B.n432 B.n431 10.6151
R2222 B.n431 B.n112 10.6151
R2223 B.n193 B.n1 10.6151
R2224 B.n194 B.n193 10.6151
R2225 B.n195 B.n194 10.6151
R2226 B.n195 B.n190 10.6151
R2227 B.n199 B.n190 10.6151
R2228 B.n200 B.n199 10.6151
R2229 B.n201 B.n200 10.6151
R2230 B.n201 B.n188 10.6151
R2231 B.n205 B.n188 10.6151
R2232 B.n206 B.n205 10.6151
R2233 B.n207 B.n206 10.6151
R2234 B.n207 B.n186 10.6151
R2235 B.n211 B.n186 10.6151
R2236 B.n212 B.n211 10.6151
R2237 B.n213 B.n212 10.6151
R2238 B.n213 B.n184 10.6151
R2239 B.n217 B.n184 10.6151
R2240 B.n218 B.n217 10.6151
R2241 B.n219 B.n218 10.6151
R2242 B.n219 B.n182 10.6151
R2243 B.n223 B.n182 10.6151
R2244 B.n224 B.n223 10.6151
R2245 B.n225 B.n224 10.6151
R2246 B.n225 B.n180 10.6151
R2247 B.n229 B.n180 10.6151
R2248 B.n230 B.n229 10.6151
R2249 B.n231 B.n178 10.6151
R2250 B.n235 B.n178 10.6151
R2251 B.n236 B.n235 10.6151
R2252 B.n237 B.n236 10.6151
R2253 B.n237 B.n176 10.6151
R2254 B.n241 B.n176 10.6151
R2255 B.n242 B.n241 10.6151
R2256 B.n243 B.n242 10.6151
R2257 B.n243 B.n174 10.6151
R2258 B.n247 B.n174 10.6151
R2259 B.n248 B.n247 10.6151
R2260 B.n249 B.n248 10.6151
R2261 B.n249 B.n172 10.6151
R2262 B.n253 B.n172 10.6151
R2263 B.n254 B.n253 10.6151
R2264 B.n255 B.n254 10.6151
R2265 B.n255 B.n170 10.6151
R2266 B.n259 B.n170 10.6151
R2267 B.n260 B.n259 10.6151
R2268 B.n261 B.n260 10.6151
R2269 B.n261 B.n168 10.6151
R2270 B.n265 B.n168 10.6151
R2271 B.n266 B.n265 10.6151
R2272 B.n267 B.n266 10.6151
R2273 B.n267 B.n166 10.6151
R2274 B.n271 B.n166 10.6151
R2275 B.n272 B.n271 10.6151
R2276 B.n273 B.n272 10.6151
R2277 B.n273 B.n164 10.6151
R2278 B.n277 B.n164 10.6151
R2279 B.n278 B.n277 10.6151
R2280 B.n279 B.n278 10.6151
R2281 B.n279 B.n162 10.6151
R2282 B.n283 B.n162 10.6151
R2283 B.n284 B.n283 10.6151
R2284 B.n285 B.n284 10.6151
R2285 B.n285 B.n160 10.6151
R2286 B.n289 B.n160 10.6151
R2287 B.n290 B.n289 10.6151
R2288 B.n291 B.n290 10.6151
R2289 B.n291 B.n158 10.6151
R2290 B.n295 B.n158 10.6151
R2291 B.n296 B.n295 10.6151
R2292 B.n297 B.n296 10.6151
R2293 B.n297 B.n156 10.6151
R2294 B.n301 B.n156 10.6151
R2295 B.n302 B.n301 10.6151
R2296 B.n303 B.n302 10.6151
R2297 B.n303 B.n154 10.6151
R2298 B.n307 B.n154 10.6151
R2299 B.n308 B.n307 10.6151
R2300 B.n309 B.n308 10.6151
R2301 B.n309 B.n152 10.6151
R2302 B.n313 B.n152 10.6151
R2303 B.n314 B.n313 10.6151
R2304 B.n315 B.n314 10.6151
R2305 B.n315 B.n150 10.6151
R2306 B.n319 B.n150 10.6151
R2307 B.n320 B.n319 10.6151
R2308 B.n322 B.n146 10.6151
R2309 B.n326 B.n146 10.6151
R2310 B.n327 B.n326 10.6151
R2311 B.n328 B.n327 10.6151
R2312 B.n328 B.n144 10.6151
R2313 B.n332 B.n144 10.6151
R2314 B.n333 B.n332 10.6151
R2315 B.n337 B.n333 10.6151
R2316 B.n341 B.n142 10.6151
R2317 B.n342 B.n341 10.6151
R2318 B.n343 B.n342 10.6151
R2319 B.n343 B.n140 10.6151
R2320 B.n347 B.n140 10.6151
R2321 B.n348 B.n347 10.6151
R2322 B.n349 B.n348 10.6151
R2323 B.n349 B.n138 10.6151
R2324 B.n353 B.n138 10.6151
R2325 B.n354 B.n353 10.6151
R2326 B.n355 B.n354 10.6151
R2327 B.n355 B.n136 10.6151
R2328 B.n359 B.n136 10.6151
R2329 B.n360 B.n359 10.6151
R2330 B.n361 B.n360 10.6151
R2331 B.n361 B.n134 10.6151
R2332 B.n365 B.n134 10.6151
R2333 B.n366 B.n365 10.6151
R2334 B.n367 B.n366 10.6151
R2335 B.n367 B.n132 10.6151
R2336 B.n371 B.n132 10.6151
R2337 B.n372 B.n371 10.6151
R2338 B.n373 B.n372 10.6151
R2339 B.n373 B.n130 10.6151
R2340 B.n377 B.n130 10.6151
R2341 B.n378 B.n377 10.6151
R2342 B.n379 B.n378 10.6151
R2343 B.n379 B.n128 10.6151
R2344 B.n383 B.n128 10.6151
R2345 B.n384 B.n383 10.6151
R2346 B.n385 B.n384 10.6151
R2347 B.n385 B.n126 10.6151
R2348 B.n389 B.n126 10.6151
R2349 B.n390 B.n389 10.6151
R2350 B.n391 B.n390 10.6151
R2351 B.n391 B.n124 10.6151
R2352 B.n395 B.n124 10.6151
R2353 B.n396 B.n395 10.6151
R2354 B.n397 B.n396 10.6151
R2355 B.n397 B.n122 10.6151
R2356 B.n401 B.n122 10.6151
R2357 B.n402 B.n401 10.6151
R2358 B.n403 B.n402 10.6151
R2359 B.n403 B.n120 10.6151
R2360 B.n407 B.n120 10.6151
R2361 B.n408 B.n407 10.6151
R2362 B.n409 B.n408 10.6151
R2363 B.n409 B.n118 10.6151
R2364 B.n413 B.n118 10.6151
R2365 B.n414 B.n413 10.6151
R2366 B.n415 B.n414 10.6151
R2367 B.n415 B.n116 10.6151
R2368 B.n419 B.n116 10.6151
R2369 B.n420 B.n419 10.6151
R2370 B.n421 B.n420 10.6151
R2371 B.n421 B.n114 10.6151
R2372 B.n425 B.n114 10.6151
R2373 B.n426 B.n425 10.6151
R2374 B.n427 B.n426 10.6151
R2375 B.n749 B.n0 8.11757
R2376 B.n749 B.n1 8.11757
R2377 B.n617 B.n616 6.5566
R2378 B.n604 B.n54 6.5566
R2379 B.n322 B.n321 6.5566
R2380 B.n337 B.n336 6.5566
R2381 B.n618 B.n617 4.05904
R2382 B.n601 B.n54 4.05904
R2383 B.n321 B.n320 4.05904
R2384 B.n336 B.n142 4.05904
C0 VN B 1.04058f
C1 VP VDD2 0.347979f
C2 VTAIL VDD2 7.10601f
C3 VDD1 w_n2296_n4588# 1.47317f
C4 VP VN 6.80205f
C5 VP B 1.52401f
C6 VN VTAIL 6.10386f
C7 VTAIL B 6.49452f
C8 VDD1 VDD2 0.851707f
C9 VN VDD1 0.147838f
C10 VDD1 B 1.29993f
C11 w_n2296_n4588# VDD2 1.51319f
C12 VP VTAIL 6.11797f
C13 VN w_n2296_n4588# 3.86798f
C14 w_n2296_n4588# B 10.070001f
C15 VP VDD1 6.74677f
C16 VTAIL VDD1 7.05663f
C17 VN VDD2 6.54719f
C18 B VDD2 1.34029f
C19 VP w_n2296_n4588# 4.16133f
C20 VTAIL w_n2296_n4588# 5.38465f
C21 VDD2 VSUBS 0.978104f
C22 VDD1 VSUBS 6.12255f
C23 VTAIL VSUBS 1.430611f
C24 VN VSUBS 5.50214f
C25 VP VSUBS 2.118095f
C26 B VSUBS 4.16697f
C27 w_n2296_n4588# VSUBS 0.128806p
C28 B.n0 VSUBS 0.005785f
C29 B.n1 VSUBS 0.005785f
C30 B.n2 VSUBS 0.008556f
C31 B.n3 VSUBS 0.006556f
C32 B.n4 VSUBS 0.006556f
C33 B.n5 VSUBS 0.006556f
C34 B.n6 VSUBS 0.006556f
C35 B.n7 VSUBS 0.006556f
C36 B.n8 VSUBS 0.006556f
C37 B.n9 VSUBS 0.006556f
C38 B.n10 VSUBS 0.006556f
C39 B.n11 VSUBS 0.006556f
C40 B.n12 VSUBS 0.006556f
C41 B.n13 VSUBS 0.006556f
C42 B.n14 VSUBS 0.006556f
C43 B.n15 VSUBS 0.014588f
C44 B.n16 VSUBS 0.006556f
C45 B.n17 VSUBS 0.006556f
C46 B.n18 VSUBS 0.006556f
C47 B.n19 VSUBS 0.006556f
C48 B.n20 VSUBS 0.006556f
C49 B.n21 VSUBS 0.006556f
C50 B.n22 VSUBS 0.006556f
C51 B.n23 VSUBS 0.006556f
C52 B.n24 VSUBS 0.006556f
C53 B.n25 VSUBS 0.006556f
C54 B.n26 VSUBS 0.006556f
C55 B.n27 VSUBS 0.006556f
C56 B.n28 VSUBS 0.006556f
C57 B.n29 VSUBS 0.006556f
C58 B.n30 VSUBS 0.006556f
C59 B.n31 VSUBS 0.006556f
C60 B.n32 VSUBS 0.006556f
C61 B.n33 VSUBS 0.006556f
C62 B.n34 VSUBS 0.006556f
C63 B.n35 VSUBS 0.006556f
C64 B.n36 VSUBS 0.006556f
C65 B.n37 VSUBS 0.006556f
C66 B.n38 VSUBS 0.006556f
C67 B.n39 VSUBS 0.006556f
C68 B.n40 VSUBS 0.006556f
C69 B.n41 VSUBS 0.006556f
C70 B.n42 VSUBS 0.006556f
C71 B.n43 VSUBS 0.006556f
C72 B.n44 VSUBS 0.006556f
C73 B.n45 VSUBS 0.006556f
C74 B.t4 VSUBS 0.330961f
C75 B.t5 VSUBS 0.355058f
C76 B.t3 VSUBS 1.37868f
C77 B.n46 VSUBS 0.516888f
C78 B.n47 VSUBS 0.306329f
C79 B.n48 VSUBS 0.006556f
C80 B.n49 VSUBS 0.006556f
C81 B.n50 VSUBS 0.006556f
C82 B.n51 VSUBS 0.006556f
C83 B.t10 VSUBS 0.330964f
C84 B.t11 VSUBS 0.355061f
C85 B.t9 VSUBS 1.37868f
C86 B.n52 VSUBS 0.516885f
C87 B.n53 VSUBS 0.306326f
C88 B.n54 VSUBS 0.01519f
C89 B.n55 VSUBS 0.006556f
C90 B.n56 VSUBS 0.006556f
C91 B.n57 VSUBS 0.006556f
C92 B.n58 VSUBS 0.006556f
C93 B.n59 VSUBS 0.006556f
C94 B.n60 VSUBS 0.006556f
C95 B.n61 VSUBS 0.006556f
C96 B.n62 VSUBS 0.006556f
C97 B.n63 VSUBS 0.006556f
C98 B.n64 VSUBS 0.006556f
C99 B.n65 VSUBS 0.006556f
C100 B.n66 VSUBS 0.006556f
C101 B.n67 VSUBS 0.006556f
C102 B.n68 VSUBS 0.006556f
C103 B.n69 VSUBS 0.006556f
C104 B.n70 VSUBS 0.006556f
C105 B.n71 VSUBS 0.006556f
C106 B.n72 VSUBS 0.006556f
C107 B.n73 VSUBS 0.006556f
C108 B.n74 VSUBS 0.006556f
C109 B.n75 VSUBS 0.006556f
C110 B.n76 VSUBS 0.006556f
C111 B.n77 VSUBS 0.006556f
C112 B.n78 VSUBS 0.006556f
C113 B.n79 VSUBS 0.006556f
C114 B.n80 VSUBS 0.006556f
C115 B.n81 VSUBS 0.006556f
C116 B.n82 VSUBS 0.006556f
C117 B.n83 VSUBS 0.006556f
C118 B.n84 VSUBS 0.015687f
C119 B.n85 VSUBS 0.006556f
C120 B.n86 VSUBS 0.006556f
C121 B.n87 VSUBS 0.006556f
C122 B.n88 VSUBS 0.006556f
C123 B.n89 VSUBS 0.006556f
C124 B.n90 VSUBS 0.006556f
C125 B.n91 VSUBS 0.006556f
C126 B.n92 VSUBS 0.006556f
C127 B.n93 VSUBS 0.006556f
C128 B.n94 VSUBS 0.006556f
C129 B.n95 VSUBS 0.006556f
C130 B.n96 VSUBS 0.006556f
C131 B.n97 VSUBS 0.006556f
C132 B.n98 VSUBS 0.006556f
C133 B.n99 VSUBS 0.006556f
C134 B.n100 VSUBS 0.006556f
C135 B.n101 VSUBS 0.006556f
C136 B.n102 VSUBS 0.006556f
C137 B.n103 VSUBS 0.006556f
C138 B.n104 VSUBS 0.006556f
C139 B.n105 VSUBS 0.006556f
C140 B.n106 VSUBS 0.006556f
C141 B.n107 VSUBS 0.006556f
C142 B.n108 VSUBS 0.006556f
C143 B.n109 VSUBS 0.006556f
C144 B.n110 VSUBS 0.006556f
C145 B.n111 VSUBS 0.006556f
C146 B.n112 VSUBS 0.015378f
C147 B.n113 VSUBS 0.006556f
C148 B.n114 VSUBS 0.006556f
C149 B.n115 VSUBS 0.006556f
C150 B.n116 VSUBS 0.006556f
C151 B.n117 VSUBS 0.006556f
C152 B.n118 VSUBS 0.006556f
C153 B.n119 VSUBS 0.006556f
C154 B.n120 VSUBS 0.006556f
C155 B.n121 VSUBS 0.006556f
C156 B.n122 VSUBS 0.006556f
C157 B.n123 VSUBS 0.006556f
C158 B.n124 VSUBS 0.006556f
C159 B.n125 VSUBS 0.006556f
C160 B.n126 VSUBS 0.006556f
C161 B.n127 VSUBS 0.006556f
C162 B.n128 VSUBS 0.006556f
C163 B.n129 VSUBS 0.006556f
C164 B.n130 VSUBS 0.006556f
C165 B.n131 VSUBS 0.006556f
C166 B.n132 VSUBS 0.006556f
C167 B.n133 VSUBS 0.006556f
C168 B.n134 VSUBS 0.006556f
C169 B.n135 VSUBS 0.006556f
C170 B.n136 VSUBS 0.006556f
C171 B.n137 VSUBS 0.006556f
C172 B.n138 VSUBS 0.006556f
C173 B.n139 VSUBS 0.006556f
C174 B.n140 VSUBS 0.006556f
C175 B.n141 VSUBS 0.006556f
C176 B.n142 VSUBS 0.004532f
C177 B.n143 VSUBS 0.006556f
C178 B.n144 VSUBS 0.006556f
C179 B.n145 VSUBS 0.006556f
C180 B.n146 VSUBS 0.006556f
C181 B.n147 VSUBS 0.006556f
C182 B.t2 VSUBS 0.330961f
C183 B.t1 VSUBS 0.355058f
C184 B.t0 VSUBS 1.37868f
C185 B.n148 VSUBS 0.516888f
C186 B.n149 VSUBS 0.306329f
C187 B.n150 VSUBS 0.006556f
C188 B.n151 VSUBS 0.006556f
C189 B.n152 VSUBS 0.006556f
C190 B.n153 VSUBS 0.006556f
C191 B.n154 VSUBS 0.006556f
C192 B.n155 VSUBS 0.006556f
C193 B.n156 VSUBS 0.006556f
C194 B.n157 VSUBS 0.006556f
C195 B.n158 VSUBS 0.006556f
C196 B.n159 VSUBS 0.006556f
C197 B.n160 VSUBS 0.006556f
C198 B.n161 VSUBS 0.006556f
C199 B.n162 VSUBS 0.006556f
C200 B.n163 VSUBS 0.006556f
C201 B.n164 VSUBS 0.006556f
C202 B.n165 VSUBS 0.006556f
C203 B.n166 VSUBS 0.006556f
C204 B.n167 VSUBS 0.006556f
C205 B.n168 VSUBS 0.006556f
C206 B.n169 VSUBS 0.006556f
C207 B.n170 VSUBS 0.006556f
C208 B.n171 VSUBS 0.006556f
C209 B.n172 VSUBS 0.006556f
C210 B.n173 VSUBS 0.006556f
C211 B.n174 VSUBS 0.006556f
C212 B.n175 VSUBS 0.006556f
C213 B.n176 VSUBS 0.006556f
C214 B.n177 VSUBS 0.006556f
C215 B.n178 VSUBS 0.006556f
C216 B.n179 VSUBS 0.014588f
C217 B.n180 VSUBS 0.006556f
C218 B.n181 VSUBS 0.006556f
C219 B.n182 VSUBS 0.006556f
C220 B.n183 VSUBS 0.006556f
C221 B.n184 VSUBS 0.006556f
C222 B.n185 VSUBS 0.006556f
C223 B.n186 VSUBS 0.006556f
C224 B.n187 VSUBS 0.006556f
C225 B.n188 VSUBS 0.006556f
C226 B.n189 VSUBS 0.006556f
C227 B.n190 VSUBS 0.006556f
C228 B.n191 VSUBS 0.006556f
C229 B.n192 VSUBS 0.006556f
C230 B.n193 VSUBS 0.006556f
C231 B.n194 VSUBS 0.006556f
C232 B.n195 VSUBS 0.006556f
C233 B.n196 VSUBS 0.006556f
C234 B.n197 VSUBS 0.006556f
C235 B.n198 VSUBS 0.006556f
C236 B.n199 VSUBS 0.006556f
C237 B.n200 VSUBS 0.006556f
C238 B.n201 VSUBS 0.006556f
C239 B.n202 VSUBS 0.006556f
C240 B.n203 VSUBS 0.006556f
C241 B.n204 VSUBS 0.006556f
C242 B.n205 VSUBS 0.006556f
C243 B.n206 VSUBS 0.006556f
C244 B.n207 VSUBS 0.006556f
C245 B.n208 VSUBS 0.006556f
C246 B.n209 VSUBS 0.006556f
C247 B.n210 VSUBS 0.006556f
C248 B.n211 VSUBS 0.006556f
C249 B.n212 VSUBS 0.006556f
C250 B.n213 VSUBS 0.006556f
C251 B.n214 VSUBS 0.006556f
C252 B.n215 VSUBS 0.006556f
C253 B.n216 VSUBS 0.006556f
C254 B.n217 VSUBS 0.006556f
C255 B.n218 VSUBS 0.006556f
C256 B.n219 VSUBS 0.006556f
C257 B.n220 VSUBS 0.006556f
C258 B.n221 VSUBS 0.006556f
C259 B.n222 VSUBS 0.006556f
C260 B.n223 VSUBS 0.006556f
C261 B.n224 VSUBS 0.006556f
C262 B.n225 VSUBS 0.006556f
C263 B.n226 VSUBS 0.006556f
C264 B.n227 VSUBS 0.006556f
C265 B.n228 VSUBS 0.006556f
C266 B.n229 VSUBS 0.006556f
C267 B.n230 VSUBS 0.014588f
C268 B.n231 VSUBS 0.015687f
C269 B.n232 VSUBS 0.015687f
C270 B.n233 VSUBS 0.006556f
C271 B.n234 VSUBS 0.006556f
C272 B.n235 VSUBS 0.006556f
C273 B.n236 VSUBS 0.006556f
C274 B.n237 VSUBS 0.006556f
C275 B.n238 VSUBS 0.006556f
C276 B.n239 VSUBS 0.006556f
C277 B.n240 VSUBS 0.006556f
C278 B.n241 VSUBS 0.006556f
C279 B.n242 VSUBS 0.006556f
C280 B.n243 VSUBS 0.006556f
C281 B.n244 VSUBS 0.006556f
C282 B.n245 VSUBS 0.006556f
C283 B.n246 VSUBS 0.006556f
C284 B.n247 VSUBS 0.006556f
C285 B.n248 VSUBS 0.006556f
C286 B.n249 VSUBS 0.006556f
C287 B.n250 VSUBS 0.006556f
C288 B.n251 VSUBS 0.006556f
C289 B.n252 VSUBS 0.006556f
C290 B.n253 VSUBS 0.006556f
C291 B.n254 VSUBS 0.006556f
C292 B.n255 VSUBS 0.006556f
C293 B.n256 VSUBS 0.006556f
C294 B.n257 VSUBS 0.006556f
C295 B.n258 VSUBS 0.006556f
C296 B.n259 VSUBS 0.006556f
C297 B.n260 VSUBS 0.006556f
C298 B.n261 VSUBS 0.006556f
C299 B.n262 VSUBS 0.006556f
C300 B.n263 VSUBS 0.006556f
C301 B.n264 VSUBS 0.006556f
C302 B.n265 VSUBS 0.006556f
C303 B.n266 VSUBS 0.006556f
C304 B.n267 VSUBS 0.006556f
C305 B.n268 VSUBS 0.006556f
C306 B.n269 VSUBS 0.006556f
C307 B.n270 VSUBS 0.006556f
C308 B.n271 VSUBS 0.006556f
C309 B.n272 VSUBS 0.006556f
C310 B.n273 VSUBS 0.006556f
C311 B.n274 VSUBS 0.006556f
C312 B.n275 VSUBS 0.006556f
C313 B.n276 VSUBS 0.006556f
C314 B.n277 VSUBS 0.006556f
C315 B.n278 VSUBS 0.006556f
C316 B.n279 VSUBS 0.006556f
C317 B.n280 VSUBS 0.006556f
C318 B.n281 VSUBS 0.006556f
C319 B.n282 VSUBS 0.006556f
C320 B.n283 VSUBS 0.006556f
C321 B.n284 VSUBS 0.006556f
C322 B.n285 VSUBS 0.006556f
C323 B.n286 VSUBS 0.006556f
C324 B.n287 VSUBS 0.006556f
C325 B.n288 VSUBS 0.006556f
C326 B.n289 VSUBS 0.006556f
C327 B.n290 VSUBS 0.006556f
C328 B.n291 VSUBS 0.006556f
C329 B.n292 VSUBS 0.006556f
C330 B.n293 VSUBS 0.006556f
C331 B.n294 VSUBS 0.006556f
C332 B.n295 VSUBS 0.006556f
C333 B.n296 VSUBS 0.006556f
C334 B.n297 VSUBS 0.006556f
C335 B.n298 VSUBS 0.006556f
C336 B.n299 VSUBS 0.006556f
C337 B.n300 VSUBS 0.006556f
C338 B.n301 VSUBS 0.006556f
C339 B.n302 VSUBS 0.006556f
C340 B.n303 VSUBS 0.006556f
C341 B.n304 VSUBS 0.006556f
C342 B.n305 VSUBS 0.006556f
C343 B.n306 VSUBS 0.006556f
C344 B.n307 VSUBS 0.006556f
C345 B.n308 VSUBS 0.006556f
C346 B.n309 VSUBS 0.006556f
C347 B.n310 VSUBS 0.006556f
C348 B.n311 VSUBS 0.006556f
C349 B.n312 VSUBS 0.006556f
C350 B.n313 VSUBS 0.006556f
C351 B.n314 VSUBS 0.006556f
C352 B.n315 VSUBS 0.006556f
C353 B.n316 VSUBS 0.006556f
C354 B.n317 VSUBS 0.006556f
C355 B.n318 VSUBS 0.006556f
C356 B.n319 VSUBS 0.006556f
C357 B.n320 VSUBS 0.004532f
C358 B.n321 VSUBS 0.01519f
C359 B.n322 VSUBS 0.005303f
C360 B.n323 VSUBS 0.006556f
C361 B.n324 VSUBS 0.006556f
C362 B.n325 VSUBS 0.006556f
C363 B.n326 VSUBS 0.006556f
C364 B.n327 VSUBS 0.006556f
C365 B.n328 VSUBS 0.006556f
C366 B.n329 VSUBS 0.006556f
C367 B.n330 VSUBS 0.006556f
C368 B.n331 VSUBS 0.006556f
C369 B.n332 VSUBS 0.006556f
C370 B.n333 VSUBS 0.006556f
C371 B.t8 VSUBS 0.330964f
C372 B.t7 VSUBS 0.355061f
C373 B.t6 VSUBS 1.37868f
C374 B.n334 VSUBS 0.516885f
C375 B.n335 VSUBS 0.306326f
C376 B.n336 VSUBS 0.01519f
C377 B.n337 VSUBS 0.005303f
C378 B.n338 VSUBS 0.006556f
C379 B.n339 VSUBS 0.006556f
C380 B.n340 VSUBS 0.006556f
C381 B.n341 VSUBS 0.006556f
C382 B.n342 VSUBS 0.006556f
C383 B.n343 VSUBS 0.006556f
C384 B.n344 VSUBS 0.006556f
C385 B.n345 VSUBS 0.006556f
C386 B.n346 VSUBS 0.006556f
C387 B.n347 VSUBS 0.006556f
C388 B.n348 VSUBS 0.006556f
C389 B.n349 VSUBS 0.006556f
C390 B.n350 VSUBS 0.006556f
C391 B.n351 VSUBS 0.006556f
C392 B.n352 VSUBS 0.006556f
C393 B.n353 VSUBS 0.006556f
C394 B.n354 VSUBS 0.006556f
C395 B.n355 VSUBS 0.006556f
C396 B.n356 VSUBS 0.006556f
C397 B.n357 VSUBS 0.006556f
C398 B.n358 VSUBS 0.006556f
C399 B.n359 VSUBS 0.006556f
C400 B.n360 VSUBS 0.006556f
C401 B.n361 VSUBS 0.006556f
C402 B.n362 VSUBS 0.006556f
C403 B.n363 VSUBS 0.006556f
C404 B.n364 VSUBS 0.006556f
C405 B.n365 VSUBS 0.006556f
C406 B.n366 VSUBS 0.006556f
C407 B.n367 VSUBS 0.006556f
C408 B.n368 VSUBS 0.006556f
C409 B.n369 VSUBS 0.006556f
C410 B.n370 VSUBS 0.006556f
C411 B.n371 VSUBS 0.006556f
C412 B.n372 VSUBS 0.006556f
C413 B.n373 VSUBS 0.006556f
C414 B.n374 VSUBS 0.006556f
C415 B.n375 VSUBS 0.006556f
C416 B.n376 VSUBS 0.006556f
C417 B.n377 VSUBS 0.006556f
C418 B.n378 VSUBS 0.006556f
C419 B.n379 VSUBS 0.006556f
C420 B.n380 VSUBS 0.006556f
C421 B.n381 VSUBS 0.006556f
C422 B.n382 VSUBS 0.006556f
C423 B.n383 VSUBS 0.006556f
C424 B.n384 VSUBS 0.006556f
C425 B.n385 VSUBS 0.006556f
C426 B.n386 VSUBS 0.006556f
C427 B.n387 VSUBS 0.006556f
C428 B.n388 VSUBS 0.006556f
C429 B.n389 VSUBS 0.006556f
C430 B.n390 VSUBS 0.006556f
C431 B.n391 VSUBS 0.006556f
C432 B.n392 VSUBS 0.006556f
C433 B.n393 VSUBS 0.006556f
C434 B.n394 VSUBS 0.006556f
C435 B.n395 VSUBS 0.006556f
C436 B.n396 VSUBS 0.006556f
C437 B.n397 VSUBS 0.006556f
C438 B.n398 VSUBS 0.006556f
C439 B.n399 VSUBS 0.006556f
C440 B.n400 VSUBS 0.006556f
C441 B.n401 VSUBS 0.006556f
C442 B.n402 VSUBS 0.006556f
C443 B.n403 VSUBS 0.006556f
C444 B.n404 VSUBS 0.006556f
C445 B.n405 VSUBS 0.006556f
C446 B.n406 VSUBS 0.006556f
C447 B.n407 VSUBS 0.006556f
C448 B.n408 VSUBS 0.006556f
C449 B.n409 VSUBS 0.006556f
C450 B.n410 VSUBS 0.006556f
C451 B.n411 VSUBS 0.006556f
C452 B.n412 VSUBS 0.006556f
C453 B.n413 VSUBS 0.006556f
C454 B.n414 VSUBS 0.006556f
C455 B.n415 VSUBS 0.006556f
C456 B.n416 VSUBS 0.006556f
C457 B.n417 VSUBS 0.006556f
C458 B.n418 VSUBS 0.006556f
C459 B.n419 VSUBS 0.006556f
C460 B.n420 VSUBS 0.006556f
C461 B.n421 VSUBS 0.006556f
C462 B.n422 VSUBS 0.006556f
C463 B.n423 VSUBS 0.006556f
C464 B.n424 VSUBS 0.006556f
C465 B.n425 VSUBS 0.006556f
C466 B.n426 VSUBS 0.006556f
C467 B.n427 VSUBS 0.014896f
C468 B.n428 VSUBS 0.015687f
C469 B.n429 VSUBS 0.014588f
C470 B.n430 VSUBS 0.006556f
C471 B.n431 VSUBS 0.006556f
C472 B.n432 VSUBS 0.006556f
C473 B.n433 VSUBS 0.006556f
C474 B.n434 VSUBS 0.006556f
C475 B.n435 VSUBS 0.006556f
C476 B.n436 VSUBS 0.006556f
C477 B.n437 VSUBS 0.006556f
C478 B.n438 VSUBS 0.006556f
C479 B.n439 VSUBS 0.006556f
C480 B.n440 VSUBS 0.006556f
C481 B.n441 VSUBS 0.006556f
C482 B.n442 VSUBS 0.006556f
C483 B.n443 VSUBS 0.006556f
C484 B.n444 VSUBS 0.006556f
C485 B.n445 VSUBS 0.006556f
C486 B.n446 VSUBS 0.006556f
C487 B.n447 VSUBS 0.006556f
C488 B.n448 VSUBS 0.006556f
C489 B.n449 VSUBS 0.006556f
C490 B.n450 VSUBS 0.006556f
C491 B.n451 VSUBS 0.006556f
C492 B.n452 VSUBS 0.006556f
C493 B.n453 VSUBS 0.006556f
C494 B.n454 VSUBS 0.006556f
C495 B.n455 VSUBS 0.006556f
C496 B.n456 VSUBS 0.006556f
C497 B.n457 VSUBS 0.006556f
C498 B.n458 VSUBS 0.006556f
C499 B.n459 VSUBS 0.006556f
C500 B.n460 VSUBS 0.006556f
C501 B.n461 VSUBS 0.006556f
C502 B.n462 VSUBS 0.006556f
C503 B.n463 VSUBS 0.006556f
C504 B.n464 VSUBS 0.006556f
C505 B.n465 VSUBS 0.006556f
C506 B.n466 VSUBS 0.006556f
C507 B.n467 VSUBS 0.006556f
C508 B.n468 VSUBS 0.006556f
C509 B.n469 VSUBS 0.006556f
C510 B.n470 VSUBS 0.006556f
C511 B.n471 VSUBS 0.006556f
C512 B.n472 VSUBS 0.006556f
C513 B.n473 VSUBS 0.006556f
C514 B.n474 VSUBS 0.006556f
C515 B.n475 VSUBS 0.006556f
C516 B.n476 VSUBS 0.006556f
C517 B.n477 VSUBS 0.006556f
C518 B.n478 VSUBS 0.006556f
C519 B.n479 VSUBS 0.006556f
C520 B.n480 VSUBS 0.006556f
C521 B.n481 VSUBS 0.006556f
C522 B.n482 VSUBS 0.006556f
C523 B.n483 VSUBS 0.006556f
C524 B.n484 VSUBS 0.006556f
C525 B.n485 VSUBS 0.006556f
C526 B.n486 VSUBS 0.006556f
C527 B.n487 VSUBS 0.006556f
C528 B.n488 VSUBS 0.006556f
C529 B.n489 VSUBS 0.006556f
C530 B.n490 VSUBS 0.006556f
C531 B.n491 VSUBS 0.006556f
C532 B.n492 VSUBS 0.006556f
C533 B.n493 VSUBS 0.006556f
C534 B.n494 VSUBS 0.006556f
C535 B.n495 VSUBS 0.006556f
C536 B.n496 VSUBS 0.006556f
C537 B.n497 VSUBS 0.006556f
C538 B.n498 VSUBS 0.006556f
C539 B.n499 VSUBS 0.006556f
C540 B.n500 VSUBS 0.006556f
C541 B.n501 VSUBS 0.006556f
C542 B.n502 VSUBS 0.006556f
C543 B.n503 VSUBS 0.006556f
C544 B.n504 VSUBS 0.006556f
C545 B.n505 VSUBS 0.006556f
C546 B.n506 VSUBS 0.006556f
C547 B.n507 VSUBS 0.006556f
C548 B.n508 VSUBS 0.006556f
C549 B.n509 VSUBS 0.006556f
C550 B.n510 VSUBS 0.006556f
C551 B.n511 VSUBS 0.014588f
C552 B.n512 VSUBS 0.014588f
C553 B.n513 VSUBS 0.015687f
C554 B.n514 VSUBS 0.006556f
C555 B.n515 VSUBS 0.006556f
C556 B.n516 VSUBS 0.006556f
C557 B.n517 VSUBS 0.006556f
C558 B.n518 VSUBS 0.006556f
C559 B.n519 VSUBS 0.006556f
C560 B.n520 VSUBS 0.006556f
C561 B.n521 VSUBS 0.006556f
C562 B.n522 VSUBS 0.006556f
C563 B.n523 VSUBS 0.006556f
C564 B.n524 VSUBS 0.006556f
C565 B.n525 VSUBS 0.006556f
C566 B.n526 VSUBS 0.006556f
C567 B.n527 VSUBS 0.006556f
C568 B.n528 VSUBS 0.006556f
C569 B.n529 VSUBS 0.006556f
C570 B.n530 VSUBS 0.006556f
C571 B.n531 VSUBS 0.006556f
C572 B.n532 VSUBS 0.006556f
C573 B.n533 VSUBS 0.006556f
C574 B.n534 VSUBS 0.006556f
C575 B.n535 VSUBS 0.006556f
C576 B.n536 VSUBS 0.006556f
C577 B.n537 VSUBS 0.006556f
C578 B.n538 VSUBS 0.006556f
C579 B.n539 VSUBS 0.006556f
C580 B.n540 VSUBS 0.006556f
C581 B.n541 VSUBS 0.006556f
C582 B.n542 VSUBS 0.006556f
C583 B.n543 VSUBS 0.006556f
C584 B.n544 VSUBS 0.006556f
C585 B.n545 VSUBS 0.006556f
C586 B.n546 VSUBS 0.006556f
C587 B.n547 VSUBS 0.006556f
C588 B.n548 VSUBS 0.006556f
C589 B.n549 VSUBS 0.006556f
C590 B.n550 VSUBS 0.006556f
C591 B.n551 VSUBS 0.006556f
C592 B.n552 VSUBS 0.006556f
C593 B.n553 VSUBS 0.006556f
C594 B.n554 VSUBS 0.006556f
C595 B.n555 VSUBS 0.006556f
C596 B.n556 VSUBS 0.006556f
C597 B.n557 VSUBS 0.006556f
C598 B.n558 VSUBS 0.006556f
C599 B.n559 VSUBS 0.006556f
C600 B.n560 VSUBS 0.006556f
C601 B.n561 VSUBS 0.006556f
C602 B.n562 VSUBS 0.006556f
C603 B.n563 VSUBS 0.006556f
C604 B.n564 VSUBS 0.006556f
C605 B.n565 VSUBS 0.006556f
C606 B.n566 VSUBS 0.006556f
C607 B.n567 VSUBS 0.006556f
C608 B.n568 VSUBS 0.006556f
C609 B.n569 VSUBS 0.006556f
C610 B.n570 VSUBS 0.006556f
C611 B.n571 VSUBS 0.006556f
C612 B.n572 VSUBS 0.006556f
C613 B.n573 VSUBS 0.006556f
C614 B.n574 VSUBS 0.006556f
C615 B.n575 VSUBS 0.006556f
C616 B.n576 VSUBS 0.006556f
C617 B.n577 VSUBS 0.006556f
C618 B.n578 VSUBS 0.006556f
C619 B.n579 VSUBS 0.006556f
C620 B.n580 VSUBS 0.006556f
C621 B.n581 VSUBS 0.006556f
C622 B.n582 VSUBS 0.006556f
C623 B.n583 VSUBS 0.006556f
C624 B.n584 VSUBS 0.006556f
C625 B.n585 VSUBS 0.006556f
C626 B.n586 VSUBS 0.006556f
C627 B.n587 VSUBS 0.006556f
C628 B.n588 VSUBS 0.006556f
C629 B.n589 VSUBS 0.006556f
C630 B.n590 VSUBS 0.006556f
C631 B.n591 VSUBS 0.006556f
C632 B.n592 VSUBS 0.006556f
C633 B.n593 VSUBS 0.006556f
C634 B.n594 VSUBS 0.006556f
C635 B.n595 VSUBS 0.006556f
C636 B.n596 VSUBS 0.006556f
C637 B.n597 VSUBS 0.006556f
C638 B.n598 VSUBS 0.006556f
C639 B.n599 VSUBS 0.006556f
C640 B.n600 VSUBS 0.006556f
C641 B.n601 VSUBS 0.004532f
C642 B.n602 VSUBS 0.006556f
C643 B.n603 VSUBS 0.006556f
C644 B.n604 VSUBS 0.005303f
C645 B.n605 VSUBS 0.006556f
C646 B.n606 VSUBS 0.006556f
C647 B.n607 VSUBS 0.006556f
C648 B.n608 VSUBS 0.006556f
C649 B.n609 VSUBS 0.006556f
C650 B.n610 VSUBS 0.006556f
C651 B.n611 VSUBS 0.006556f
C652 B.n612 VSUBS 0.006556f
C653 B.n613 VSUBS 0.006556f
C654 B.n614 VSUBS 0.006556f
C655 B.n615 VSUBS 0.006556f
C656 B.n616 VSUBS 0.005303f
C657 B.n617 VSUBS 0.01519f
C658 B.n618 VSUBS 0.004532f
C659 B.n619 VSUBS 0.006556f
C660 B.n620 VSUBS 0.006556f
C661 B.n621 VSUBS 0.006556f
C662 B.n622 VSUBS 0.006556f
C663 B.n623 VSUBS 0.006556f
C664 B.n624 VSUBS 0.006556f
C665 B.n625 VSUBS 0.006556f
C666 B.n626 VSUBS 0.006556f
C667 B.n627 VSUBS 0.006556f
C668 B.n628 VSUBS 0.006556f
C669 B.n629 VSUBS 0.006556f
C670 B.n630 VSUBS 0.006556f
C671 B.n631 VSUBS 0.006556f
C672 B.n632 VSUBS 0.006556f
C673 B.n633 VSUBS 0.006556f
C674 B.n634 VSUBS 0.006556f
C675 B.n635 VSUBS 0.006556f
C676 B.n636 VSUBS 0.006556f
C677 B.n637 VSUBS 0.006556f
C678 B.n638 VSUBS 0.006556f
C679 B.n639 VSUBS 0.006556f
C680 B.n640 VSUBS 0.006556f
C681 B.n641 VSUBS 0.006556f
C682 B.n642 VSUBS 0.006556f
C683 B.n643 VSUBS 0.006556f
C684 B.n644 VSUBS 0.006556f
C685 B.n645 VSUBS 0.006556f
C686 B.n646 VSUBS 0.006556f
C687 B.n647 VSUBS 0.006556f
C688 B.n648 VSUBS 0.006556f
C689 B.n649 VSUBS 0.006556f
C690 B.n650 VSUBS 0.006556f
C691 B.n651 VSUBS 0.006556f
C692 B.n652 VSUBS 0.006556f
C693 B.n653 VSUBS 0.006556f
C694 B.n654 VSUBS 0.006556f
C695 B.n655 VSUBS 0.006556f
C696 B.n656 VSUBS 0.006556f
C697 B.n657 VSUBS 0.006556f
C698 B.n658 VSUBS 0.006556f
C699 B.n659 VSUBS 0.006556f
C700 B.n660 VSUBS 0.006556f
C701 B.n661 VSUBS 0.006556f
C702 B.n662 VSUBS 0.006556f
C703 B.n663 VSUBS 0.006556f
C704 B.n664 VSUBS 0.006556f
C705 B.n665 VSUBS 0.006556f
C706 B.n666 VSUBS 0.006556f
C707 B.n667 VSUBS 0.006556f
C708 B.n668 VSUBS 0.006556f
C709 B.n669 VSUBS 0.006556f
C710 B.n670 VSUBS 0.006556f
C711 B.n671 VSUBS 0.006556f
C712 B.n672 VSUBS 0.006556f
C713 B.n673 VSUBS 0.006556f
C714 B.n674 VSUBS 0.006556f
C715 B.n675 VSUBS 0.006556f
C716 B.n676 VSUBS 0.006556f
C717 B.n677 VSUBS 0.006556f
C718 B.n678 VSUBS 0.006556f
C719 B.n679 VSUBS 0.006556f
C720 B.n680 VSUBS 0.006556f
C721 B.n681 VSUBS 0.006556f
C722 B.n682 VSUBS 0.006556f
C723 B.n683 VSUBS 0.006556f
C724 B.n684 VSUBS 0.006556f
C725 B.n685 VSUBS 0.006556f
C726 B.n686 VSUBS 0.006556f
C727 B.n687 VSUBS 0.006556f
C728 B.n688 VSUBS 0.006556f
C729 B.n689 VSUBS 0.006556f
C730 B.n690 VSUBS 0.006556f
C731 B.n691 VSUBS 0.006556f
C732 B.n692 VSUBS 0.006556f
C733 B.n693 VSUBS 0.006556f
C734 B.n694 VSUBS 0.006556f
C735 B.n695 VSUBS 0.006556f
C736 B.n696 VSUBS 0.006556f
C737 B.n697 VSUBS 0.006556f
C738 B.n698 VSUBS 0.006556f
C739 B.n699 VSUBS 0.006556f
C740 B.n700 VSUBS 0.006556f
C741 B.n701 VSUBS 0.006556f
C742 B.n702 VSUBS 0.006556f
C743 B.n703 VSUBS 0.006556f
C744 B.n704 VSUBS 0.006556f
C745 B.n705 VSUBS 0.006556f
C746 B.n706 VSUBS 0.015687f
C747 B.n707 VSUBS 0.015687f
C748 B.n708 VSUBS 0.014588f
C749 B.n709 VSUBS 0.006556f
C750 B.n710 VSUBS 0.006556f
C751 B.n711 VSUBS 0.006556f
C752 B.n712 VSUBS 0.006556f
C753 B.n713 VSUBS 0.006556f
C754 B.n714 VSUBS 0.006556f
C755 B.n715 VSUBS 0.006556f
C756 B.n716 VSUBS 0.006556f
C757 B.n717 VSUBS 0.006556f
C758 B.n718 VSUBS 0.006556f
C759 B.n719 VSUBS 0.006556f
C760 B.n720 VSUBS 0.006556f
C761 B.n721 VSUBS 0.006556f
C762 B.n722 VSUBS 0.006556f
C763 B.n723 VSUBS 0.006556f
C764 B.n724 VSUBS 0.006556f
C765 B.n725 VSUBS 0.006556f
C766 B.n726 VSUBS 0.006556f
C767 B.n727 VSUBS 0.006556f
C768 B.n728 VSUBS 0.006556f
C769 B.n729 VSUBS 0.006556f
C770 B.n730 VSUBS 0.006556f
C771 B.n731 VSUBS 0.006556f
C772 B.n732 VSUBS 0.006556f
C773 B.n733 VSUBS 0.006556f
C774 B.n734 VSUBS 0.006556f
C775 B.n735 VSUBS 0.006556f
C776 B.n736 VSUBS 0.006556f
C777 B.n737 VSUBS 0.006556f
C778 B.n738 VSUBS 0.006556f
C779 B.n739 VSUBS 0.006556f
C780 B.n740 VSUBS 0.006556f
C781 B.n741 VSUBS 0.006556f
C782 B.n742 VSUBS 0.006556f
C783 B.n743 VSUBS 0.006556f
C784 B.n744 VSUBS 0.006556f
C785 B.n745 VSUBS 0.006556f
C786 B.n746 VSUBS 0.006556f
C787 B.n747 VSUBS 0.008556f
C788 B.n748 VSUBS 0.009114f
C789 B.n749 VSUBS 0.018124f
C790 VDD1.t0 VSUBS 0.380245f
C791 VDD1.t3 VSUBS 0.380245f
C792 VDD1.n0 VSUBS 3.18939f
C793 VDD1.t1 VSUBS 0.380245f
C794 VDD1.t2 VSUBS 0.380245f
C795 VDD1.n1 VSUBS 4.09433f
C796 VP.n0 VSUBS 0.036693f
C797 VP.t1 VSUBS 3.4347f
C798 VP.n1 VSUBS 0.029693f
C799 VP.n2 VSUBS 0.036693f
C800 VP.t2 VSUBS 3.4347f
C801 VP.t3 VSUBS 3.62831f
C802 VP.t0 VSUBS 3.62607f
C803 VP.n3 VSUBS 4.29143f
C804 VP.n4 VSUBS 2.29801f
C805 VP.n5 VSUBS 1.29113f
C806 VP.n6 VSUBS 0.041921f
C807 VP.n7 VSUBS 0.073317f
C808 VP.n8 VSUBS 0.036693f
C809 VP.n9 VSUBS 0.036693f
C810 VP.n10 VSUBS 0.036693f
C811 VP.n11 VSUBS 0.073317f
C812 VP.n12 VSUBS 0.041921f
C813 VP.n13 VSUBS 1.29113f
C814 VP.n14 VSUBS 0.039264f
C815 VTAIL.n0 VSUBS 0.012381f
C816 VTAIL.n1 VSUBS 0.027869f
C817 VTAIL.n2 VSUBS 0.012484f
C818 VTAIL.n3 VSUBS 0.021942f
C819 VTAIL.n4 VSUBS 0.011791f
C820 VTAIL.n5 VSUBS 0.027869f
C821 VTAIL.n6 VSUBS 0.012484f
C822 VTAIL.n7 VSUBS 0.021942f
C823 VTAIL.n8 VSUBS 0.011791f
C824 VTAIL.n9 VSUBS 0.027869f
C825 VTAIL.n10 VSUBS 0.012484f
C826 VTAIL.n11 VSUBS 0.021942f
C827 VTAIL.n12 VSUBS 0.011791f
C828 VTAIL.n13 VSUBS 0.027869f
C829 VTAIL.n14 VSUBS 0.012484f
C830 VTAIL.n15 VSUBS 0.021942f
C831 VTAIL.n16 VSUBS 0.011791f
C832 VTAIL.n17 VSUBS 0.027869f
C833 VTAIL.n18 VSUBS 0.012484f
C834 VTAIL.n19 VSUBS 0.021942f
C835 VTAIL.n20 VSUBS 0.011791f
C836 VTAIL.n21 VSUBS 0.027869f
C837 VTAIL.n22 VSUBS 0.012484f
C838 VTAIL.n23 VSUBS 0.021942f
C839 VTAIL.n24 VSUBS 0.011791f
C840 VTAIL.n25 VSUBS 0.027869f
C841 VTAIL.n26 VSUBS 0.012484f
C842 VTAIL.n27 VSUBS 0.021942f
C843 VTAIL.n28 VSUBS 0.011791f
C844 VTAIL.n29 VSUBS 0.027869f
C845 VTAIL.n30 VSUBS 0.012484f
C846 VTAIL.n31 VSUBS 0.233327f
C847 VTAIL.t6 VSUBS 0.060506f
C848 VTAIL.n32 VSUBS 0.020902f
C849 VTAIL.n33 VSUBS 0.020965f
C850 VTAIL.n34 VSUBS 0.011791f
C851 VTAIL.n35 VSUBS 1.66456f
C852 VTAIL.n36 VSUBS 0.021942f
C853 VTAIL.n37 VSUBS 0.011791f
C854 VTAIL.n38 VSUBS 0.012484f
C855 VTAIL.n39 VSUBS 0.027869f
C856 VTAIL.n40 VSUBS 0.027869f
C857 VTAIL.n41 VSUBS 0.012484f
C858 VTAIL.n42 VSUBS 0.011791f
C859 VTAIL.n43 VSUBS 0.021942f
C860 VTAIL.n44 VSUBS 0.021942f
C861 VTAIL.n45 VSUBS 0.011791f
C862 VTAIL.n46 VSUBS 0.012484f
C863 VTAIL.n47 VSUBS 0.027869f
C864 VTAIL.n48 VSUBS 0.027869f
C865 VTAIL.n49 VSUBS 0.027869f
C866 VTAIL.n50 VSUBS 0.012484f
C867 VTAIL.n51 VSUBS 0.011791f
C868 VTAIL.n52 VSUBS 0.021942f
C869 VTAIL.n53 VSUBS 0.021942f
C870 VTAIL.n54 VSUBS 0.011791f
C871 VTAIL.n55 VSUBS 0.012138f
C872 VTAIL.n56 VSUBS 0.012138f
C873 VTAIL.n57 VSUBS 0.027869f
C874 VTAIL.n58 VSUBS 0.027869f
C875 VTAIL.n59 VSUBS 0.012484f
C876 VTAIL.n60 VSUBS 0.011791f
C877 VTAIL.n61 VSUBS 0.021942f
C878 VTAIL.n62 VSUBS 0.021942f
C879 VTAIL.n63 VSUBS 0.011791f
C880 VTAIL.n64 VSUBS 0.012484f
C881 VTAIL.n65 VSUBS 0.027869f
C882 VTAIL.n66 VSUBS 0.027869f
C883 VTAIL.n67 VSUBS 0.012484f
C884 VTAIL.n68 VSUBS 0.011791f
C885 VTAIL.n69 VSUBS 0.021942f
C886 VTAIL.n70 VSUBS 0.021942f
C887 VTAIL.n71 VSUBS 0.011791f
C888 VTAIL.n72 VSUBS 0.012484f
C889 VTAIL.n73 VSUBS 0.027869f
C890 VTAIL.n74 VSUBS 0.027869f
C891 VTAIL.n75 VSUBS 0.012484f
C892 VTAIL.n76 VSUBS 0.011791f
C893 VTAIL.n77 VSUBS 0.021942f
C894 VTAIL.n78 VSUBS 0.021942f
C895 VTAIL.n79 VSUBS 0.011791f
C896 VTAIL.n80 VSUBS 0.012484f
C897 VTAIL.n81 VSUBS 0.027869f
C898 VTAIL.n82 VSUBS 0.027869f
C899 VTAIL.n83 VSUBS 0.012484f
C900 VTAIL.n84 VSUBS 0.011791f
C901 VTAIL.n85 VSUBS 0.021942f
C902 VTAIL.n86 VSUBS 0.021942f
C903 VTAIL.n87 VSUBS 0.011791f
C904 VTAIL.n88 VSUBS 0.012484f
C905 VTAIL.n89 VSUBS 0.027869f
C906 VTAIL.n90 VSUBS 0.027869f
C907 VTAIL.n91 VSUBS 0.012484f
C908 VTAIL.n92 VSUBS 0.011791f
C909 VTAIL.n93 VSUBS 0.021942f
C910 VTAIL.n94 VSUBS 0.057313f
C911 VTAIL.n95 VSUBS 0.011791f
C912 VTAIL.n96 VSUBS 0.012484f
C913 VTAIL.n97 VSUBS 0.06272f
C914 VTAIL.n98 VSUBS 0.042184f
C915 VTAIL.n99 VSUBS 0.126136f
C916 VTAIL.n100 VSUBS 0.012381f
C917 VTAIL.n101 VSUBS 0.027869f
C918 VTAIL.n102 VSUBS 0.012484f
C919 VTAIL.n103 VSUBS 0.021942f
C920 VTAIL.n104 VSUBS 0.011791f
C921 VTAIL.n105 VSUBS 0.027869f
C922 VTAIL.n106 VSUBS 0.012484f
C923 VTAIL.n107 VSUBS 0.021942f
C924 VTAIL.n108 VSUBS 0.011791f
C925 VTAIL.n109 VSUBS 0.027869f
C926 VTAIL.n110 VSUBS 0.012484f
C927 VTAIL.n111 VSUBS 0.021942f
C928 VTAIL.n112 VSUBS 0.011791f
C929 VTAIL.n113 VSUBS 0.027869f
C930 VTAIL.n114 VSUBS 0.012484f
C931 VTAIL.n115 VSUBS 0.021942f
C932 VTAIL.n116 VSUBS 0.011791f
C933 VTAIL.n117 VSUBS 0.027869f
C934 VTAIL.n118 VSUBS 0.012484f
C935 VTAIL.n119 VSUBS 0.021942f
C936 VTAIL.n120 VSUBS 0.011791f
C937 VTAIL.n121 VSUBS 0.027869f
C938 VTAIL.n122 VSUBS 0.012484f
C939 VTAIL.n123 VSUBS 0.021942f
C940 VTAIL.n124 VSUBS 0.011791f
C941 VTAIL.n125 VSUBS 0.027869f
C942 VTAIL.n126 VSUBS 0.012484f
C943 VTAIL.n127 VSUBS 0.021942f
C944 VTAIL.n128 VSUBS 0.011791f
C945 VTAIL.n129 VSUBS 0.027869f
C946 VTAIL.n130 VSUBS 0.012484f
C947 VTAIL.n131 VSUBS 0.233327f
C948 VTAIL.t7 VSUBS 0.060506f
C949 VTAIL.n132 VSUBS 0.020902f
C950 VTAIL.n133 VSUBS 0.020965f
C951 VTAIL.n134 VSUBS 0.011791f
C952 VTAIL.n135 VSUBS 1.66456f
C953 VTAIL.n136 VSUBS 0.021942f
C954 VTAIL.n137 VSUBS 0.011791f
C955 VTAIL.n138 VSUBS 0.012484f
C956 VTAIL.n139 VSUBS 0.027869f
C957 VTAIL.n140 VSUBS 0.027869f
C958 VTAIL.n141 VSUBS 0.012484f
C959 VTAIL.n142 VSUBS 0.011791f
C960 VTAIL.n143 VSUBS 0.021942f
C961 VTAIL.n144 VSUBS 0.021942f
C962 VTAIL.n145 VSUBS 0.011791f
C963 VTAIL.n146 VSUBS 0.012484f
C964 VTAIL.n147 VSUBS 0.027869f
C965 VTAIL.n148 VSUBS 0.027869f
C966 VTAIL.n149 VSUBS 0.027869f
C967 VTAIL.n150 VSUBS 0.012484f
C968 VTAIL.n151 VSUBS 0.011791f
C969 VTAIL.n152 VSUBS 0.021942f
C970 VTAIL.n153 VSUBS 0.021942f
C971 VTAIL.n154 VSUBS 0.011791f
C972 VTAIL.n155 VSUBS 0.012138f
C973 VTAIL.n156 VSUBS 0.012138f
C974 VTAIL.n157 VSUBS 0.027869f
C975 VTAIL.n158 VSUBS 0.027869f
C976 VTAIL.n159 VSUBS 0.012484f
C977 VTAIL.n160 VSUBS 0.011791f
C978 VTAIL.n161 VSUBS 0.021942f
C979 VTAIL.n162 VSUBS 0.021942f
C980 VTAIL.n163 VSUBS 0.011791f
C981 VTAIL.n164 VSUBS 0.012484f
C982 VTAIL.n165 VSUBS 0.027869f
C983 VTAIL.n166 VSUBS 0.027869f
C984 VTAIL.n167 VSUBS 0.012484f
C985 VTAIL.n168 VSUBS 0.011791f
C986 VTAIL.n169 VSUBS 0.021942f
C987 VTAIL.n170 VSUBS 0.021942f
C988 VTAIL.n171 VSUBS 0.011791f
C989 VTAIL.n172 VSUBS 0.012484f
C990 VTAIL.n173 VSUBS 0.027869f
C991 VTAIL.n174 VSUBS 0.027869f
C992 VTAIL.n175 VSUBS 0.012484f
C993 VTAIL.n176 VSUBS 0.011791f
C994 VTAIL.n177 VSUBS 0.021942f
C995 VTAIL.n178 VSUBS 0.021942f
C996 VTAIL.n179 VSUBS 0.011791f
C997 VTAIL.n180 VSUBS 0.012484f
C998 VTAIL.n181 VSUBS 0.027869f
C999 VTAIL.n182 VSUBS 0.027869f
C1000 VTAIL.n183 VSUBS 0.012484f
C1001 VTAIL.n184 VSUBS 0.011791f
C1002 VTAIL.n185 VSUBS 0.021942f
C1003 VTAIL.n186 VSUBS 0.021942f
C1004 VTAIL.n187 VSUBS 0.011791f
C1005 VTAIL.n188 VSUBS 0.012484f
C1006 VTAIL.n189 VSUBS 0.027869f
C1007 VTAIL.n190 VSUBS 0.027869f
C1008 VTAIL.n191 VSUBS 0.012484f
C1009 VTAIL.n192 VSUBS 0.011791f
C1010 VTAIL.n193 VSUBS 0.021942f
C1011 VTAIL.n194 VSUBS 0.057313f
C1012 VTAIL.n195 VSUBS 0.011791f
C1013 VTAIL.n196 VSUBS 0.012484f
C1014 VTAIL.n197 VSUBS 0.06272f
C1015 VTAIL.n198 VSUBS 0.042184f
C1016 VTAIL.n199 VSUBS 0.189372f
C1017 VTAIL.n200 VSUBS 0.012381f
C1018 VTAIL.n201 VSUBS 0.027869f
C1019 VTAIL.n202 VSUBS 0.012484f
C1020 VTAIL.n203 VSUBS 0.021942f
C1021 VTAIL.n204 VSUBS 0.011791f
C1022 VTAIL.n205 VSUBS 0.027869f
C1023 VTAIL.n206 VSUBS 0.012484f
C1024 VTAIL.n207 VSUBS 0.021942f
C1025 VTAIL.n208 VSUBS 0.011791f
C1026 VTAIL.n209 VSUBS 0.027869f
C1027 VTAIL.n210 VSUBS 0.012484f
C1028 VTAIL.n211 VSUBS 0.021942f
C1029 VTAIL.n212 VSUBS 0.011791f
C1030 VTAIL.n213 VSUBS 0.027869f
C1031 VTAIL.n214 VSUBS 0.012484f
C1032 VTAIL.n215 VSUBS 0.021942f
C1033 VTAIL.n216 VSUBS 0.011791f
C1034 VTAIL.n217 VSUBS 0.027869f
C1035 VTAIL.n218 VSUBS 0.012484f
C1036 VTAIL.n219 VSUBS 0.021942f
C1037 VTAIL.n220 VSUBS 0.011791f
C1038 VTAIL.n221 VSUBS 0.027869f
C1039 VTAIL.n222 VSUBS 0.012484f
C1040 VTAIL.n223 VSUBS 0.021942f
C1041 VTAIL.n224 VSUBS 0.011791f
C1042 VTAIL.n225 VSUBS 0.027869f
C1043 VTAIL.n226 VSUBS 0.012484f
C1044 VTAIL.n227 VSUBS 0.021942f
C1045 VTAIL.n228 VSUBS 0.011791f
C1046 VTAIL.n229 VSUBS 0.027869f
C1047 VTAIL.n230 VSUBS 0.012484f
C1048 VTAIL.n231 VSUBS 0.233327f
C1049 VTAIL.t2 VSUBS 0.060506f
C1050 VTAIL.n232 VSUBS 0.020902f
C1051 VTAIL.n233 VSUBS 0.020965f
C1052 VTAIL.n234 VSUBS 0.011791f
C1053 VTAIL.n235 VSUBS 1.66456f
C1054 VTAIL.n236 VSUBS 0.021942f
C1055 VTAIL.n237 VSUBS 0.011791f
C1056 VTAIL.n238 VSUBS 0.012484f
C1057 VTAIL.n239 VSUBS 0.027869f
C1058 VTAIL.n240 VSUBS 0.027869f
C1059 VTAIL.n241 VSUBS 0.012484f
C1060 VTAIL.n242 VSUBS 0.011791f
C1061 VTAIL.n243 VSUBS 0.021942f
C1062 VTAIL.n244 VSUBS 0.021942f
C1063 VTAIL.n245 VSUBS 0.011791f
C1064 VTAIL.n246 VSUBS 0.012484f
C1065 VTAIL.n247 VSUBS 0.027869f
C1066 VTAIL.n248 VSUBS 0.027869f
C1067 VTAIL.n249 VSUBS 0.027869f
C1068 VTAIL.n250 VSUBS 0.012484f
C1069 VTAIL.n251 VSUBS 0.011791f
C1070 VTAIL.n252 VSUBS 0.021942f
C1071 VTAIL.n253 VSUBS 0.021942f
C1072 VTAIL.n254 VSUBS 0.011791f
C1073 VTAIL.n255 VSUBS 0.012138f
C1074 VTAIL.n256 VSUBS 0.012138f
C1075 VTAIL.n257 VSUBS 0.027869f
C1076 VTAIL.n258 VSUBS 0.027869f
C1077 VTAIL.n259 VSUBS 0.012484f
C1078 VTAIL.n260 VSUBS 0.011791f
C1079 VTAIL.n261 VSUBS 0.021942f
C1080 VTAIL.n262 VSUBS 0.021942f
C1081 VTAIL.n263 VSUBS 0.011791f
C1082 VTAIL.n264 VSUBS 0.012484f
C1083 VTAIL.n265 VSUBS 0.027869f
C1084 VTAIL.n266 VSUBS 0.027869f
C1085 VTAIL.n267 VSUBS 0.012484f
C1086 VTAIL.n268 VSUBS 0.011791f
C1087 VTAIL.n269 VSUBS 0.021942f
C1088 VTAIL.n270 VSUBS 0.021942f
C1089 VTAIL.n271 VSUBS 0.011791f
C1090 VTAIL.n272 VSUBS 0.012484f
C1091 VTAIL.n273 VSUBS 0.027869f
C1092 VTAIL.n274 VSUBS 0.027869f
C1093 VTAIL.n275 VSUBS 0.012484f
C1094 VTAIL.n276 VSUBS 0.011791f
C1095 VTAIL.n277 VSUBS 0.021942f
C1096 VTAIL.n278 VSUBS 0.021942f
C1097 VTAIL.n279 VSUBS 0.011791f
C1098 VTAIL.n280 VSUBS 0.012484f
C1099 VTAIL.n281 VSUBS 0.027869f
C1100 VTAIL.n282 VSUBS 0.027869f
C1101 VTAIL.n283 VSUBS 0.012484f
C1102 VTAIL.n284 VSUBS 0.011791f
C1103 VTAIL.n285 VSUBS 0.021942f
C1104 VTAIL.n286 VSUBS 0.021942f
C1105 VTAIL.n287 VSUBS 0.011791f
C1106 VTAIL.n288 VSUBS 0.012484f
C1107 VTAIL.n289 VSUBS 0.027869f
C1108 VTAIL.n290 VSUBS 0.027869f
C1109 VTAIL.n291 VSUBS 0.012484f
C1110 VTAIL.n292 VSUBS 0.011791f
C1111 VTAIL.n293 VSUBS 0.021942f
C1112 VTAIL.n294 VSUBS 0.057313f
C1113 VTAIL.n295 VSUBS 0.011791f
C1114 VTAIL.n296 VSUBS 0.012484f
C1115 VTAIL.n297 VSUBS 0.06272f
C1116 VTAIL.n298 VSUBS 0.042184f
C1117 VTAIL.n299 VSUBS 1.69212f
C1118 VTAIL.n300 VSUBS 0.012381f
C1119 VTAIL.n301 VSUBS 0.027869f
C1120 VTAIL.n302 VSUBS 0.012484f
C1121 VTAIL.n303 VSUBS 0.021942f
C1122 VTAIL.n304 VSUBS 0.011791f
C1123 VTAIL.n305 VSUBS 0.027869f
C1124 VTAIL.n306 VSUBS 0.012484f
C1125 VTAIL.n307 VSUBS 0.021942f
C1126 VTAIL.n308 VSUBS 0.011791f
C1127 VTAIL.n309 VSUBS 0.027869f
C1128 VTAIL.n310 VSUBS 0.012484f
C1129 VTAIL.n311 VSUBS 0.021942f
C1130 VTAIL.n312 VSUBS 0.011791f
C1131 VTAIL.n313 VSUBS 0.027869f
C1132 VTAIL.n314 VSUBS 0.012484f
C1133 VTAIL.n315 VSUBS 0.021942f
C1134 VTAIL.n316 VSUBS 0.011791f
C1135 VTAIL.n317 VSUBS 0.027869f
C1136 VTAIL.n318 VSUBS 0.012484f
C1137 VTAIL.n319 VSUBS 0.021942f
C1138 VTAIL.n320 VSUBS 0.011791f
C1139 VTAIL.n321 VSUBS 0.027869f
C1140 VTAIL.n322 VSUBS 0.012484f
C1141 VTAIL.n323 VSUBS 0.021942f
C1142 VTAIL.n324 VSUBS 0.011791f
C1143 VTAIL.n325 VSUBS 0.027869f
C1144 VTAIL.n326 VSUBS 0.027869f
C1145 VTAIL.n327 VSUBS 0.012484f
C1146 VTAIL.n328 VSUBS 0.021942f
C1147 VTAIL.n329 VSUBS 0.011791f
C1148 VTAIL.n330 VSUBS 0.027869f
C1149 VTAIL.n331 VSUBS 0.012484f
C1150 VTAIL.n332 VSUBS 0.233327f
C1151 VTAIL.t3 VSUBS 0.060506f
C1152 VTAIL.n333 VSUBS 0.020902f
C1153 VTAIL.n334 VSUBS 0.020965f
C1154 VTAIL.n335 VSUBS 0.011791f
C1155 VTAIL.n336 VSUBS 1.66456f
C1156 VTAIL.n337 VSUBS 0.021942f
C1157 VTAIL.n338 VSUBS 0.011791f
C1158 VTAIL.n339 VSUBS 0.012484f
C1159 VTAIL.n340 VSUBS 0.027869f
C1160 VTAIL.n341 VSUBS 0.027869f
C1161 VTAIL.n342 VSUBS 0.012484f
C1162 VTAIL.n343 VSUBS 0.011791f
C1163 VTAIL.n344 VSUBS 0.021942f
C1164 VTAIL.n345 VSUBS 0.021942f
C1165 VTAIL.n346 VSUBS 0.011791f
C1166 VTAIL.n347 VSUBS 0.012484f
C1167 VTAIL.n348 VSUBS 0.027869f
C1168 VTAIL.n349 VSUBS 0.027869f
C1169 VTAIL.n350 VSUBS 0.012484f
C1170 VTAIL.n351 VSUBS 0.011791f
C1171 VTAIL.n352 VSUBS 0.021942f
C1172 VTAIL.n353 VSUBS 0.021942f
C1173 VTAIL.n354 VSUBS 0.011791f
C1174 VTAIL.n355 VSUBS 0.012138f
C1175 VTAIL.n356 VSUBS 0.012138f
C1176 VTAIL.n357 VSUBS 0.027869f
C1177 VTAIL.n358 VSUBS 0.027869f
C1178 VTAIL.n359 VSUBS 0.012484f
C1179 VTAIL.n360 VSUBS 0.011791f
C1180 VTAIL.n361 VSUBS 0.021942f
C1181 VTAIL.n362 VSUBS 0.021942f
C1182 VTAIL.n363 VSUBS 0.011791f
C1183 VTAIL.n364 VSUBS 0.012484f
C1184 VTAIL.n365 VSUBS 0.027869f
C1185 VTAIL.n366 VSUBS 0.027869f
C1186 VTAIL.n367 VSUBS 0.012484f
C1187 VTAIL.n368 VSUBS 0.011791f
C1188 VTAIL.n369 VSUBS 0.021942f
C1189 VTAIL.n370 VSUBS 0.021942f
C1190 VTAIL.n371 VSUBS 0.011791f
C1191 VTAIL.n372 VSUBS 0.012484f
C1192 VTAIL.n373 VSUBS 0.027869f
C1193 VTAIL.n374 VSUBS 0.027869f
C1194 VTAIL.n375 VSUBS 0.012484f
C1195 VTAIL.n376 VSUBS 0.011791f
C1196 VTAIL.n377 VSUBS 0.021942f
C1197 VTAIL.n378 VSUBS 0.021942f
C1198 VTAIL.n379 VSUBS 0.011791f
C1199 VTAIL.n380 VSUBS 0.012484f
C1200 VTAIL.n381 VSUBS 0.027869f
C1201 VTAIL.n382 VSUBS 0.027869f
C1202 VTAIL.n383 VSUBS 0.012484f
C1203 VTAIL.n384 VSUBS 0.011791f
C1204 VTAIL.n385 VSUBS 0.021942f
C1205 VTAIL.n386 VSUBS 0.021942f
C1206 VTAIL.n387 VSUBS 0.011791f
C1207 VTAIL.n388 VSUBS 0.012484f
C1208 VTAIL.n389 VSUBS 0.027869f
C1209 VTAIL.n390 VSUBS 0.027869f
C1210 VTAIL.n391 VSUBS 0.012484f
C1211 VTAIL.n392 VSUBS 0.011791f
C1212 VTAIL.n393 VSUBS 0.021942f
C1213 VTAIL.n394 VSUBS 0.057313f
C1214 VTAIL.n395 VSUBS 0.011791f
C1215 VTAIL.n396 VSUBS 0.012484f
C1216 VTAIL.n397 VSUBS 0.06272f
C1217 VTAIL.n398 VSUBS 0.042184f
C1218 VTAIL.n399 VSUBS 1.69212f
C1219 VTAIL.n400 VSUBS 0.012381f
C1220 VTAIL.n401 VSUBS 0.027869f
C1221 VTAIL.n402 VSUBS 0.012484f
C1222 VTAIL.n403 VSUBS 0.021942f
C1223 VTAIL.n404 VSUBS 0.011791f
C1224 VTAIL.n405 VSUBS 0.027869f
C1225 VTAIL.n406 VSUBS 0.012484f
C1226 VTAIL.n407 VSUBS 0.021942f
C1227 VTAIL.n408 VSUBS 0.011791f
C1228 VTAIL.n409 VSUBS 0.027869f
C1229 VTAIL.n410 VSUBS 0.012484f
C1230 VTAIL.n411 VSUBS 0.021942f
C1231 VTAIL.n412 VSUBS 0.011791f
C1232 VTAIL.n413 VSUBS 0.027869f
C1233 VTAIL.n414 VSUBS 0.012484f
C1234 VTAIL.n415 VSUBS 0.021942f
C1235 VTAIL.n416 VSUBS 0.011791f
C1236 VTAIL.n417 VSUBS 0.027869f
C1237 VTAIL.n418 VSUBS 0.012484f
C1238 VTAIL.n419 VSUBS 0.021942f
C1239 VTAIL.n420 VSUBS 0.011791f
C1240 VTAIL.n421 VSUBS 0.027869f
C1241 VTAIL.n422 VSUBS 0.012484f
C1242 VTAIL.n423 VSUBS 0.021942f
C1243 VTAIL.n424 VSUBS 0.011791f
C1244 VTAIL.n425 VSUBS 0.027869f
C1245 VTAIL.n426 VSUBS 0.027869f
C1246 VTAIL.n427 VSUBS 0.012484f
C1247 VTAIL.n428 VSUBS 0.021942f
C1248 VTAIL.n429 VSUBS 0.011791f
C1249 VTAIL.n430 VSUBS 0.027869f
C1250 VTAIL.n431 VSUBS 0.012484f
C1251 VTAIL.n432 VSUBS 0.233327f
C1252 VTAIL.t4 VSUBS 0.060506f
C1253 VTAIL.n433 VSUBS 0.020902f
C1254 VTAIL.n434 VSUBS 0.020965f
C1255 VTAIL.n435 VSUBS 0.011791f
C1256 VTAIL.n436 VSUBS 1.66456f
C1257 VTAIL.n437 VSUBS 0.021942f
C1258 VTAIL.n438 VSUBS 0.011791f
C1259 VTAIL.n439 VSUBS 0.012484f
C1260 VTAIL.n440 VSUBS 0.027869f
C1261 VTAIL.n441 VSUBS 0.027869f
C1262 VTAIL.n442 VSUBS 0.012484f
C1263 VTAIL.n443 VSUBS 0.011791f
C1264 VTAIL.n444 VSUBS 0.021942f
C1265 VTAIL.n445 VSUBS 0.021942f
C1266 VTAIL.n446 VSUBS 0.011791f
C1267 VTAIL.n447 VSUBS 0.012484f
C1268 VTAIL.n448 VSUBS 0.027869f
C1269 VTAIL.n449 VSUBS 0.027869f
C1270 VTAIL.n450 VSUBS 0.012484f
C1271 VTAIL.n451 VSUBS 0.011791f
C1272 VTAIL.n452 VSUBS 0.021942f
C1273 VTAIL.n453 VSUBS 0.021942f
C1274 VTAIL.n454 VSUBS 0.011791f
C1275 VTAIL.n455 VSUBS 0.012138f
C1276 VTAIL.n456 VSUBS 0.012138f
C1277 VTAIL.n457 VSUBS 0.027869f
C1278 VTAIL.n458 VSUBS 0.027869f
C1279 VTAIL.n459 VSUBS 0.012484f
C1280 VTAIL.n460 VSUBS 0.011791f
C1281 VTAIL.n461 VSUBS 0.021942f
C1282 VTAIL.n462 VSUBS 0.021942f
C1283 VTAIL.n463 VSUBS 0.011791f
C1284 VTAIL.n464 VSUBS 0.012484f
C1285 VTAIL.n465 VSUBS 0.027869f
C1286 VTAIL.n466 VSUBS 0.027869f
C1287 VTAIL.n467 VSUBS 0.012484f
C1288 VTAIL.n468 VSUBS 0.011791f
C1289 VTAIL.n469 VSUBS 0.021942f
C1290 VTAIL.n470 VSUBS 0.021942f
C1291 VTAIL.n471 VSUBS 0.011791f
C1292 VTAIL.n472 VSUBS 0.012484f
C1293 VTAIL.n473 VSUBS 0.027869f
C1294 VTAIL.n474 VSUBS 0.027869f
C1295 VTAIL.n475 VSUBS 0.012484f
C1296 VTAIL.n476 VSUBS 0.011791f
C1297 VTAIL.n477 VSUBS 0.021942f
C1298 VTAIL.n478 VSUBS 0.021942f
C1299 VTAIL.n479 VSUBS 0.011791f
C1300 VTAIL.n480 VSUBS 0.012484f
C1301 VTAIL.n481 VSUBS 0.027869f
C1302 VTAIL.n482 VSUBS 0.027869f
C1303 VTAIL.n483 VSUBS 0.012484f
C1304 VTAIL.n484 VSUBS 0.011791f
C1305 VTAIL.n485 VSUBS 0.021942f
C1306 VTAIL.n486 VSUBS 0.021942f
C1307 VTAIL.n487 VSUBS 0.011791f
C1308 VTAIL.n488 VSUBS 0.012484f
C1309 VTAIL.n489 VSUBS 0.027869f
C1310 VTAIL.n490 VSUBS 0.027869f
C1311 VTAIL.n491 VSUBS 0.012484f
C1312 VTAIL.n492 VSUBS 0.011791f
C1313 VTAIL.n493 VSUBS 0.021942f
C1314 VTAIL.n494 VSUBS 0.057313f
C1315 VTAIL.n495 VSUBS 0.011791f
C1316 VTAIL.n496 VSUBS 0.012484f
C1317 VTAIL.n497 VSUBS 0.06272f
C1318 VTAIL.n498 VSUBS 0.042184f
C1319 VTAIL.n499 VSUBS 0.189372f
C1320 VTAIL.n500 VSUBS 0.012381f
C1321 VTAIL.n501 VSUBS 0.027869f
C1322 VTAIL.n502 VSUBS 0.012484f
C1323 VTAIL.n503 VSUBS 0.021942f
C1324 VTAIL.n504 VSUBS 0.011791f
C1325 VTAIL.n505 VSUBS 0.027869f
C1326 VTAIL.n506 VSUBS 0.012484f
C1327 VTAIL.n507 VSUBS 0.021942f
C1328 VTAIL.n508 VSUBS 0.011791f
C1329 VTAIL.n509 VSUBS 0.027869f
C1330 VTAIL.n510 VSUBS 0.012484f
C1331 VTAIL.n511 VSUBS 0.021942f
C1332 VTAIL.n512 VSUBS 0.011791f
C1333 VTAIL.n513 VSUBS 0.027869f
C1334 VTAIL.n514 VSUBS 0.012484f
C1335 VTAIL.n515 VSUBS 0.021942f
C1336 VTAIL.n516 VSUBS 0.011791f
C1337 VTAIL.n517 VSUBS 0.027869f
C1338 VTAIL.n518 VSUBS 0.012484f
C1339 VTAIL.n519 VSUBS 0.021942f
C1340 VTAIL.n520 VSUBS 0.011791f
C1341 VTAIL.n521 VSUBS 0.027869f
C1342 VTAIL.n522 VSUBS 0.012484f
C1343 VTAIL.n523 VSUBS 0.021942f
C1344 VTAIL.n524 VSUBS 0.011791f
C1345 VTAIL.n525 VSUBS 0.027869f
C1346 VTAIL.n526 VSUBS 0.027869f
C1347 VTAIL.n527 VSUBS 0.012484f
C1348 VTAIL.n528 VSUBS 0.021942f
C1349 VTAIL.n529 VSUBS 0.011791f
C1350 VTAIL.n530 VSUBS 0.027869f
C1351 VTAIL.n531 VSUBS 0.012484f
C1352 VTAIL.n532 VSUBS 0.233327f
C1353 VTAIL.t1 VSUBS 0.060506f
C1354 VTAIL.n533 VSUBS 0.020902f
C1355 VTAIL.n534 VSUBS 0.020965f
C1356 VTAIL.n535 VSUBS 0.011791f
C1357 VTAIL.n536 VSUBS 1.66456f
C1358 VTAIL.n537 VSUBS 0.021942f
C1359 VTAIL.n538 VSUBS 0.011791f
C1360 VTAIL.n539 VSUBS 0.012484f
C1361 VTAIL.n540 VSUBS 0.027869f
C1362 VTAIL.n541 VSUBS 0.027869f
C1363 VTAIL.n542 VSUBS 0.012484f
C1364 VTAIL.n543 VSUBS 0.011791f
C1365 VTAIL.n544 VSUBS 0.021942f
C1366 VTAIL.n545 VSUBS 0.021942f
C1367 VTAIL.n546 VSUBS 0.011791f
C1368 VTAIL.n547 VSUBS 0.012484f
C1369 VTAIL.n548 VSUBS 0.027869f
C1370 VTAIL.n549 VSUBS 0.027869f
C1371 VTAIL.n550 VSUBS 0.012484f
C1372 VTAIL.n551 VSUBS 0.011791f
C1373 VTAIL.n552 VSUBS 0.021942f
C1374 VTAIL.n553 VSUBS 0.021942f
C1375 VTAIL.n554 VSUBS 0.011791f
C1376 VTAIL.n555 VSUBS 0.012138f
C1377 VTAIL.n556 VSUBS 0.012138f
C1378 VTAIL.n557 VSUBS 0.027869f
C1379 VTAIL.n558 VSUBS 0.027869f
C1380 VTAIL.n559 VSUBS 0.012484f
C1381 VTAIL.n560 VSUBS 0.011791f
C1382 VTAIL.n561 VSUBS 0.021942f
C1383 VTAIL.n562 VSUBS 0.021942f
C1384 VTAIL.n563 VSUBS 0.011791f
C1385 VTAIL.n564 VSUBS 0.012484f
C1386 VTAIL.n565 VSUBS 0.027869f
C1387 VTAIL.n566 VSUBS 0.027869f
C1388 VTAIL.n567 VSUBS 0.012484f
C1389 VTAIL.n568 VSUBS 0.011791f
C1390 VTAIL.n569 VSUBS 0.021942f
C1391 VTAIL.n570 VSUBS 0.021942f
C1392 VTAIL.n571 VSUBS 0.011791f
C1393 VTAIL.n572 VSUBS 0.012484f
C1394 VTAIL.n573 VSUBS 0.027869f
C1395 VTAIL.n574 VSUBS 0.027869f
C1396 VTAIL.n575 VSUBS 0.012484f
C1397 VTAIL.n576 VSUBS 0.011791f
C1398 VTAIL.n577 VSUBS 0.021942f
C1399 VTAIL.n578 VSUBS 0.021942f
C1400 VTAIL.n579 VSUBS 0.011791f
C1401 VTAIL.n580 VSUBS 0.012484f
C1402 VTAIL.n581 VSUBS 0.027869f
C1403 VTAIL.n582 VSUBS 0.027869f
C1404 VTAIL.n583 VSUBS 0.012484f
C1405 VTAIL.n584 VSUBS 0.011791f
C1406 VTAIL.n585 VSUBS 0.021942f
C1407 VTAIL.n586 VSUBS 0.021942f
C1408 VTAIL.n587 VSUBS 0.011791f
C1409 VTAIL.n588 VSUBS 0.012484f
C1410 VTAIL.n589 VSUBS 0.027869f
C1411 VTAIL.n590 VSUBS 0.027869f
C1412 VTAIL.n591 VSUBS 0.012484f
C1413 VTAIL.n592 VSUBS 0.011791f
C1414 VTAIL.n593 VSUBS 0.021942f
C1415 VTAIL.n594 VSUBS 0.057313f
C1416 VTAIL.n595 VSUBS 0.011791f
C1417 VTAIL.n596 VSUBS 0.012484f
C1418 VTAIL.n597 VSUBS 0.06272f
C1419 VTAIL.n598 VSUBS 0.042184f
C1420 VTAIL.n599 VSUBS 0.189372f
C1421 VTAIL.n600 VSUBS 0.012381f
C1422 VTAIL.n601 VSUBS 0.027869f
C1423 VTAIL.n602 VSUBS 0.012484f
C1424 VTAIL.n603 VSUBS 0.021942f
C1425 VTAIL.n604 VSUBS 0.011791f
C1426 VTAIL.n605 VSUBS 0.027869f
C1427 VTAIL.n606 VSUBS 0.012484f
C1428 VTAIL.n607 VSUBS 0.021942f
C1429 VTAIL.n608 VSUBS 0.011791f
C1430 VTAIL.n609 VSUBS 0.027869f
C1431 VTAIL.n610 VSUBS 0.012484f
C1432 VTAIL.n611 VSUBS 0.021942f
C1433 VTAIL.n612 VSUBS 0.011791f
C1434 VTAIL.n613 VSUBS 0.027869f
C1435 VTAIL.n614 VSUBS 0.012484f
C1436 VTAIL.n615 VSUBS 0.021942f
C1437 VTAIL.n616 VSUBS 0.011791f
C1438 VTAIL.n617 VSUBS 0.027869f
C1439 VTAIL.n618 VSUBS 0.012484f
C1440 VTAIL.n619 VSUBS 0.021942f
C1441 VTAIL.n620 VSUBS 0.011791f
C1442 VTAIL.n621 VSUBS 0.027869f
C1443 VTAIL.n622 VSUBS 0.012484f
C1444 VTAIL.n623 VSUBS 0.021942f
C1445 VTAIL.n624 VSUBS 0.011791f
C1446 VTAIL.n625 VSUBS 0.027869f
C1447 VTAIL.n626 VSUBS 0.027869f
C1448 VTAIL.n627 VSUBS 0.012484f
C1449 VTAIL.n628 VSUBS 0.021942f
C1450 VTAIL.n629 VSUBS 0.011791f
C1451 VTAIL.n630 VSUBS 0.027869f
C1452 VTAIL.n631 VSUBS 0.012484f
C1453 VTAIL.n632 VSUBS 0.233327f
C1454 VTAIL.t0 VSUBS 0.060506f
C1455 VTAIL.n633 VSUBS 0.020902f
C1456 VTAIL.n634 VSUBS 0.020965f
C1457 VTAIL.n635 VSUBS 0.011791f
C1458 VTAIL.n636 VSUBS 1.66456f
C1459 VTAIL.n637 VSUBS 0.021942f
C1460 VTAIL.n638 VSUBS 0.011791f
C1461 VTAIL.n639 VSUBS 0.012484f
C1462 VTAIL.n640 VSUBS 0.027869f
C1463 VTAIL.n641 VSUBS 0.027869f
C1464 VTAIL.n642 VSUBS 0.012484f
C1465 VTAIL.n643 VSUBS 0.011791f
C1466 VTAIL.n644 VSUBS 0.021942f
C1467 VTAIL.n645 VSUBS 0.021942f
C1468 VTAIL.n646 VSUBS 0.011791f
C1469 VTAIL.n647 VSUBS 0.012484f
C1470 VTAIL.n648 VSUBS 0.027869f
C1471 VTAIL.n649 VSUBS 0.027869f
C1472 VTAIL.n650 VSUBS 0.012484f
C1473 VTAIL.n651 VSUBS 0.011791f
C1474 VTAIL.n652 VSUBS 0.021942f
C1475 VTAIL.n653 VSUBS 0.021942f
C1476 VTAIL.n654 VSUBS 0.011791f
C1477 VTAIL.n655 VSUBS 0.012138f
C1478 VTAIL.n656 VSUBS 0.012138f
C1479 VTAIL.n657 VSUBS 0.027869f
C1480 VTAIL.n658 VSUBS 0.027869f
C1481 VTAIL.n659 VSUBS 0.012484f
C1482 VTAIL.n660 VSUBS 0.011791f
C1483 VTAIL.n661 VSUBS 0.021942f
C1484 VTAIL.n662 VSUBS 0.021942f
C1485 VTAIL.n663 VSUBS 0.011791f
C1486 VTAIL.n664 VSUBS 0.012484f
C1487 VTAIL.n665 VSUBS 0.027869f
C1488 VTAIL.n666 VSUBS 0.027869f
C1489 VTAIL.n667 VSUBS 0.012484f
C1490 VTAIL.n668 VSUBS 0.011791f
C1491 VTAIL.n669 VSUBS 0.021942f
C1492 VTAIL.n670 VSUBS 0.021942f
C1493 VTAIL.n671 VSUBS 0.011791f
C1494 VTAIL.n672 VSUBS 0.012484f
C1495 VTAIL.n673 VSUBS 0.027869f
C1496 VTAIL.n674 VSUBS 0.027869f
C1497 VTAIL.n675 VSUBS 0.012484f
C1498 VTAIL.n676 VSUBS 0.011791f
C1499 VTAIL.n677 VSUBS 0.021942f
C1500 VTAIL.n678 VSUBS 0.021942f
C1501 VTAIL.n679 VSUBS 0.011791f
C1502 VTAIL.n680 VSUBS 0.012484f
C1503 VTAIL.n681 VSUBS 0.027869f
C1504 VTAIL.n682 VSUBS 0.027869f
C1505 VTAIL.n683 VSUBS 0.012484f
C1506 VTAIL.n684 VSUBS 0.011791f
C1507 VTAIL.n685 VSUBS 0.021942f
C1508 VTAIL.n686 VSUBS 0.021942f
C1509 VTAIL.n687 VSUBS 0.011791f
C1510 VTAIL.n688 VSUBS 0.012484f
C1511 VTAIL.n689 VSUBS 0.027869f
C1512 VTAIL.n690 VSUBS 0.027869f
C1513 VTAIL.n691 VSUBS 0.012484f
C1514 VTAIL.n692 VSUBS 0.011791f
C1515 VTAIL.n693 VSUBS 0.021942f
C1516 VTAIL.n694 VSUBS 0.057313f
C1517 VTAIL.n695 VSUBS 0.011791f
C1518 VTAIL.n696 VSUBS 0.012484f
C1519 VTAIL.n697 VSUBS 0.06272f
C1520 VTAIL.n698 VSUBS 0.042184f
C1521 VTAIL.n699 VSUBS 1.69212f
C1522 VTAIL.n700 VSUBS 0.012381f
C1523 VTAIL.n701 VSUBS 0.027869f
C1524 VTAIL.n702 VSUBS 0.012484f
C1525 VTAIL.n703 VSUBS 0.021942f
C1526 VTAIL.n704 VSUBS 0.011791f
C1527 VTAIL.n705 VSUBS 0.027869f
C1528 VTAIL.n706 VSUBS 0.012484f
C1529 VTAIL.n707 VSUBS 0.021942f
C1530 VTAIL.n708 VSUBS 0.011791f
C1531 VTAIL.n709 VSUBS 0.027869f
C1532 VTAIL.n710 VSUBS 0.012484f
C1533 VTAIL.n711 VSUBS 0.021942f
C1534 VTAIL.n712 VSUBS 0.011791f
C1535 VTAIL.n713 VSUBS 0.027869f
C1536 VTAIL.n714 VSUBS 0.012484f
C1537 VTAIL.n715 VSUBS 0.021942f
C1538 VTAIL.n716 VSUBS 0.011791f
C1539 VTAIL.n717 VSUBS 0.027869f
C1540 VTAIL.n718 VSUBS 0.012484f
C1541 VTAIL.n719 VSUBS 0.021942f
C1542 VTAIL.n720 VSUBS 0.011791f
C1543 VTAIL.n721 VSUBS 0.027869f
C1544 VTAIL.n722 VSUBS 0.012484f
C1545 VTAIL.n723 VSUBS 0.021942f
C1546 VTAIL.n724 VSUBS 0.011791f
C1547 VTAIL.n725 VSUBS 0.027869f
C1548 VTAIL.n726 VSUBS 0.012484f
C1549 VTAIL.n727 VSUBS 0.021942f
C1550 VTAIL.n728 VSUBS 0.011791f
C1551 VTAIL.n729 VSUBS 0.027869f
C1552 VTAIL.n730 VSUBS 0.012484f
C1553 VTAIL.n731 VSUBS 0.233327f
C1554 VTAIL.t5 VSUBS 0.060506f
C1555 VTAIL.n732 VSUBS 0.020902f
C1556 VTAIL.n733 VSUBS 0.020965f
C1557 VTAIL.n734 VSUBS 0.011791f
C1558 VTAIL.n735 VSUBS 1.66456f
C1559 VTAIL.n736 VSUBS 0.021942f
C1560 VTAIL.n737 VSUBS 0.011791f
C1561 VTAIL.n738 VSUBS 0.012484f
C1562 VTAIL.n739 VSUBS 0.027869f
C1563 VTAIL.n740 VSUBS 0.027869f
C1564 VTAIL.n741 VSUBS 0.012484f
C1565 VTAIL.n742 VSUBS 0.011791f
C1566 VTAIL.n743 VSUBS 0.021942f
C1567 VTAIL.n744 VSUBS 0.021942f
C1568 VTAIL.n745 VSUBS 0.011791f
C1569 VTAIL.n746 VSUBS 0.012484f
C1570 VTAIL.n747 VSUBS 0.027869f
C1571 VTAIL.n748 VSUBS 0.027869f
C1572 VTAIL.n749 VSUBS 0.027869f
C1573 VTAIL.n750 VSUBS 0.012484f
C1574 VTAIL.n751 VSUBS 0.011791f
C1575 VTAIL.n752 VSUBS 0.021942f
C1576 VTAIL.n753 VSUBS 0.021942f
C1577 VTAIL.n754 VSUBS 0.011791f
C1578 VTAIL.n755 VSUBS 0.012138f
C1579 VTAIL.n756 VSUBS 0.012138f
C1580 VTAIL.n757 VSUBS 0.027869f
C1581 VTAIL.n758 VSUBS 0.027869f
C1582 VTAIL.n759 VSUBS 0.012484f
C1583 VTAIL.n760 VSUBS 0.011791f
C1584 VTAIL.n761 VSUBS 0.021942f
C1585 VTAIL.n762 VSUBS 0.021942f
C1586 VTAIL.n763 VSUBS 0.011791f
C1587 VTAIL.n764 VSUBS 0.012484f
C1588 VTAIL.n765 VSUBS 0.027869f
C1589 VTAIL.n766 VSUBS 0.027869f
C1590 VTAIL.n767 VSUBS 0.012484f
C1591 VTAIL.n768 VSUBS 0.011791f
C1592 VTAIL.n769 VSUBS 0.021942f
C1593 VTAIL.n770 VSUBS 0.021942f
C1594 VTAIL.n771 VSUBS 0.011791f
C1595 VTAIL.n772 VSUBS 0.012484f
C1596 VTAIL.n773 VSUBS 0.027869f
C1597 VTAIL.n774 VSUBS 0.027869f
C1598 VTAIL.n775 VSUBS 0.012484f
C1599 VTAIL.n776 VSUBS 0.011791f
C1600 VTAIL.n777 VSUBS 0.021942f
C1601 VTAIL.n778 VSUBS 0.021942f
C1602 VTAIL.n779 VSUBS 0.011791f
C1603 VTAIL.n780 VSUBS 0.012484f
C1604 VTAIL.n781 VSUBS 0.027869f
C1605 VTAIL.n782 VSUBS 0.027869f
C1606 VTAIL.n783 VSUBS 0.012484f
C1607 VTAIL.n784 VSUBS 0.011791f
C1608 VTAIL.n785 VSUBS 0.021942f
C1609 VTAIL.n786 VSUBS 0.021942f
C1610 VTAIL.n787 VSUBS 0.011791f
C1611 VTAIL.n788 VSUBS 0.012484f
C1612 VTAIL.n789 VSUBS 0.027869f
C1613 VTAIL.n790 VSUBS 0.027869f
C1614 VTAIL.n791 VSUBS 0.012484f
C1615 VTAIL.n792 VSUBS 0.011791f
C1616 VTAIL.n793 VSUBS 0.021942f
C1617 VTAIL.n794 VSUBS 0.057313f
C1618 VTAIL.n795 VSUBS 0.011791f
C1619 VTAIL.n796 VSUBS 0.012484f
C1620 VTAIL.n797 VSUBS 0.06272f
C1621 VTAIL.n798 VSUBS 0.042184f
C1622 VTAIL.n799 VSUBS 1.62065f
C1623 VDD2.t1 VSUBS 0.37742f
C1624 VDD2.t0 VSUBS 0.37742f
C1625 VDD2.n0 VSUBS 4.03754f
C1626 VDD2.t2 VSUBS 0.37742f
C1627 VDD2.t3 VSUBS 0.37742f
C1628 VDD2.n1 VSUBS 3.16515f
C1629 VDD2.n2 VSUBS 4.71996f
C1630 VN.t0 VSUBS 3.54441f
C1631 VN.t1 VSUBS 3.54222f
C1632 VN.n0 VSUBS 2.40962f
C1633 VN.t2 VSUBS 3.54441f
C1634 VN.t3 VSUBS 3.54222f
C1635 VN.n1 VSUBS 4.21405f
.ends

