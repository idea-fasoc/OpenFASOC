* NGSPICE file created from diff_pair_sample_0294.ext - technology: sky130A

.subckt diff_pair_sample_0294 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=2.9094 ps=15.7 w=7.46 l=0.93
X1 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=2.9094 ps=15.7 w=7.46 l=0.93
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=2.9094 ps=15.7 w=7.46 l=0.93
X3 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=0 ps=0 w=7.46 l=0.93
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=0 ps=0 w=7.46 l=0.93
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=0 ps=0 w=7.46 l=0.93
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=2.9094 ps=15.7 w=7.46 l=0.93
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9094 pd=15.7 as=0 ps=0 w=7.46 l=0.93
R0 VN VN.t0 434.043
R1 VN VN.t1 396.909
R2 VTAIL.n154 VTAIL.n120 289.615
R3 VTAIL.n34 VTAIL.n0 289.615
R4 VTAIL.n114 VTAIL.n80 289.615
R5 VTAIL.n74 VTAIL.n40 289.615
R6 VTAIL.n132 VTAIL.n131 185
R7 VTAIL.n137 VTAIL.n136 185
R8 VTAIL.n139 VTAIL.n138 185
R9 VTAIL.n128 VTAIL.n127 185
R10 VTAIL.n145 VTAIL.n144 185
R11 VTAIL.n147 VTAIL.n146 185
R12 VTAIL.n124 VTAIL.n123 185
R13 VTAIL.n153 VTAIL.n152 185
R14 VTAIL.n155 VTAIL.n154 185
R15 VTAIL.n12 VTAIL.n11 185
R16 VTAIL.n17 VTAIL.n16 185
R17 VTAIL.n19 VTAIL.n18 185
R18 VTAIL.n8 VTAIL.n7 185
R19 VTAIL.n25 VTAIL.n24 185
R20 VTAIL.n27 VTAIL.n26 185
R21 VTAIL.n4 VTAIL.n3 185
R22 VTAIL.n33 VTAIL.n32 185
R23 VTAIL.n35 VTAIL.n34 185
R24 VTAIL.n115 VTAIL.n114 185
R25 VTAIL.n113 VTAIL.n112 185
R26 VTAIL.n84 VTAIL.n83 185
R27 VTAIL.n107 VTAIL.n106 185
R28 VTAIL.n105 VTAIL.n104 185
R29 VTAIL.n88 VTAIL.n87 185
R30 VTAIL.n99 VTAIL.n98 185
R31 VTAIL.n97 VTAIL.n96 185
R32 VTAIL.n92 VTAIL.n91 185
R33 VTAIL.n75 VTAIL.n74 185
R34 VTAIL.n73 VTAIL.n72 185
R35 VTAIL.n44 VTAIL.n43 185
R36 VTAIL.n67 VTAIL.n66 185
R37 VTAIL.n65 VTAIL.n64 185
R38 VTAIL.n48 VTAIL.n47 185
R39 VTAIL.n59 VTAIL.n58 185
R40 VTAIL.n57 VTAIL.n56 185
R41 VTAIL.n52 VTAIL.n51 185
R42 VTAIL.n133 VTAIL.t2 147.659
R43 VTAIL.n13 VTAIL.t1 147.659
R44 VTAIL.n93 VTAIL.t0 147.659
R45 VTAIL.n53 VTAIL.t3 147.659
R46 VTAIL.n137 VTAIL.n131 104.615
R47 VTAIL.n138 VTAIL.n137 104.615
R48 VTAIL.n138 VTAIL.n127 104.615
R49 VTAIL.n145 VTAIL.n127 104.615
R50 VTAIL.n146 VTAIL.n145 104.615
R51 VTAIL.n146 VTAIL.n123 104.615
R52 VTAIL.n153 VTAIL.n123 104.615
R53 VTAIL.n154 VTAIL.n153 104.615
R54 VTAIL.n17 VTAIL.n11 104.615
R55 VTAIL.n18 VTAIL.n17 104.615
R56 VTAIL.n18 VTAIL.n7 104.615
R57 VTAIL.n25 VTAIL.n7 104.615
R58 VTAIL.n26 VTAIL.n25 104.615
R59 VTAIL.n26 VTAIL.n3 104.615
R60 VTAIL.n33 VTAIL.n3 104.615
R61 VTAIL.n34 VTAIL.n33 104.615
R62 VTAIL.n114 VTAIL.n113 104.615
R63 VTAIL.n113 VTAIL.n83 104.615
R64 VTAIL.n106 VTAIL.n83 104.615
R65 VTAIL.n106 VTAIL.n105 104.615
R66 VTAIL.n105 VTAIL.n87 104.615
R67 VTAIL.n98 VTAIL.n87 104.615
R68 VTAIL.n98 VTAIL.n97 104.615
R69 VTAIL.n97 VTAIL.n91 104.615
R70 VTAIL.n74 VTAIL.n73 104.615
R71 VTAIL.n73 VTAIL.n43 104.615
R72 VTAIL.n66 VTAIL.n43 104.615
R73 VTAIL.n66 VTAIL.n65 104.615
R74 VTAIL.n65 VTAIL.n47 104.615
R75 VTAIL.n58 VTAIL.n47 104.615
R76 VTAIL.n58 VTAIL.n57 104.615
R77 VTAIL.n57 VTAIL.n51 104.615
R78 VTAIL.t2 VTAIL.n131 52.3082
R79 VTAIL.t1 VTAIL.n11 52.3082
R80 VTAIL.t0 VTAIL.n91 52.3082
R81 VTAIL.t3 VTAIL.n51 52.3082
R82 VTAIL.n159 VTAIL.n158 32.5732
R83 VTAIL.n39 VTAIL.n38 32.5732
R84 VTAIL.n119 VTAIL.n118 32.5732
R85 VTAIL.n79 VTAIL.n78 32.5732
R86 VTAIL.n79 VTAIL.n39 20.9876
R87 VTAIL.n159 VTAIL.n119 19.9014
R88 VTAIL.n133 VTAIL.n132 15.6677
R89 VTAIL.n13 VTAIL.n12 15.6677
R90 VTAIL.n93 VTAIL.n92 15.6677
R91 VTAIL.n53 VTAIL.n52 15.6677
R92 VTAIL.n136 VTAIL.n135 12.8005
R93 VTAIL.n16 VTAIL.n15 12.8005
R94 VTAIL.n96 VTAIL.n95 12.8005
R95 VTAIL.n56 VTAIL.n55 12.8005
R96 VTAIL.n139 VTAIL.n130 12.0247
R97 VTAIL.n19 VTAIL.n10 12.0247
R98 VTAIL.n99 VTAIL.n90 12.0247
R99 VTAIL.n59 VTAIL.n50 12.0247
R100 VTAIL.n140 VTAIL.n128 11.249
R101 VTAIL.n20 VTAIL.n8 11.249
R102 VTAIL.n100 VTAIL.n88 11.249
R103 VTAIL.n60 VTAIL.n48 11.249
R104 VTAIL.n144 VTAIL.n143 10.4732
R105 VTAIL.n24 VTAIL.n23 10.4732
R106 VTAIL.n104 VTAIL.n103 10.4732
R107 VTAIL.n64 VTAIL.n63 10.4732
R108 VTAIL.n147 VTAIL.n126 9.69747
R109 VTAIL.n27 VTAIL.n6 9.69747
R110 VTAIL.n107 VTAIL.n86 9.69747
R111 VTAIL.n67 VTAIL.n46 9.69747
R112 VTAIL.n158 VTAIL.n157 9.45567
R113 VTAIL.n38 VTAIL.n37 9.45567
R114 VTAIL.n118 VTAIL.n117 9.45567
R115 VTAIL.n78 VTAIL.n77 9.45567
R116 VTAIL.n157 VTAIL.n156 9.3005
R117 VTAIL.n151 VTAIL.n150 9.3005
R118 VTAIL.n149 VTAIL.n148 9.3005
R119 VTAIL.n126 VTAIL.n125 9.3005
R120 VTAIL.n143 VTAIL.n142 9.3005
R121 VTAIL.n141 VTAIL.n140 9.3005
R122 VTAIL.n130 VTAIL.n129 9.3005
R123 VTAIL.n135 VTAIL.n134 9.3005
R124 VTAIL.n122 VTAIL.n121 9.3005
R125 VTAIL.n37 VTAIL.n36 9.3005
R126 VTAIL.n31 VTAIL.n30 9.3005
R127 VTAIL.n29 VTAIL.n28 9.3005
R128 VTAIL.n6 VTAIL.n5 9.3005
R129 VTAIL.n23 VTAIL.n22 9.3005
R130 VTAIL.n21 VTAIL.n20 9.3005
R131 VTAIL.n10 VTAIL.n9 9.3005
R132 VTAIL.n15 VTAIL.n14 9.3005
R133 VTAIL.n2 VTAIL.n1 9.3005
R134 VTAIL.n117 VTAIL.n116 9.3005
R135 VTAIL.n82 VTAIL.n81 9.3005
R136 VTAIL.n111 VTAIL.n110 9.3005
R137 VTAIL.n109 VTAIL.n108 9.3005
R138 VTAIL.n86 VTAIL.n85 9.3005
R139 VTAIL.n103 VTAIL.n102 9.3005
R140 VTAIL.n101 VTAIL.n100 9.3005
R141 VTAIL.n90 VTAIL.n89 9.3005
R142 VTAIL.n95 VTAIL.n94 9.3005
R143 VTAIL.n77 VTAIL.n76 9.3005
R144 VTAIL.n42 VTAIL.n41 9.3005
R145 VTAIL.n71 VTAIL.n70 9.3005
R146 VTAIL.n69 VTAIL.n68 9.3005
R147 VTAIL.n46 VTAIL.n45 9.3005
R148 VTAIL.n63 VTAIL.n62 9.3005
R149 VTAIL.n61 VTAIL.n60 9.3005
R150 VTAIL.n50 VTAIL.n49 9.3005
R151 VTAIL.n55 VTAIL.n54 9.3005
R152 VTAIL.n148 VTAIL.n124 8.92171
R153 VTAIL.n28 VTAIL.n4 8.92171
R154 VTAIL.n108 VTAIL.n84 8.92171
R155 VTAIL.n68 VTAIL.n44 8.92171
R156 VTAIL.n152 VTAIL.n151 8.14595
R157 VTAIL.n32 VTAIL.n31 8.14595
R158 VTAIL.n112 VTAIL.n111 8.14595
R159 VTAIL.n72 VTAIL.n71 8.14595
R160 VTAIL.n155 VTAIL.n122 7.3702
R161 VTAIL.n158 VTAIL.n120 7.3702
R162 VTAIL.n35 VTAIL.n2 7.3702
R163 VTAIL.n38 VTAIL.n0 7.3702
R164 VTAIL.n118 VTAIL.n80 7.3702
R165 VTAIL.n115 VTAIL.n82 7.3702
R166 VTAIL.n78 VTAIL.n40 7.3702
R167 VTAIL.n75 VTAIL.n42 7.3702
R168 VTAIL.n156 VTAIL.n155 6.59444
R169 VTAIL.n156 VTAIL.n120 6.59444
R170 VTAIL.n36 VTAIL.n35 6.59444
R171 VTAIL.n36 VTAIL.n0 6.59444
R172 VTAIL.n116 VTAIL.n80 6.59444
R173 VTAIL.n116 VTAIL.n115 6.59444
R174 VTAIL.n76 VTAIL.n40 6.59444
R175 VTAIL.n76 VTAIL.n75 6.59444
R176 VTAIL.n152 VTAIL.n122 5.81868
R177 VTAIL.n32 VTAIL.n2 5.81868
R178 VTAIL.n112 VTAIL.n82 5.81868
R179 VTAIL.n72 VTAIL.n42 5.81868
R180 VTAIL.n151 VTAIL.n124 5.04292
R181 VTAIL.n31 VTAIL.n4 5.04292
R182 VTAIL.n111 VTAIL.n84 5.04292
R183 VTAIL.n71 VTAIL.n44 5.04292
R184 VTAIL.n94 VTAIL.n93 4.38565
R185 VTAIL.n54 VTAIL.n53 4.38565
R186 VTAIL.n134 VTAIL.n133 4.38565
R187 VTAIL.n14 VTAIL.n13 4.38565
R188 VTAIL.n148 VTAIL.n147 4.26717
R189 VTAIL.n28 VTAIL.n27 4.26717
R190 VTAIL.n108 VTAIL.n107 4.26717
R191 VTAIL.n68 VTAIL.n67 4.26717
R192 VTAIL.n144 VTAIL.n126 3.49141
R193 VTAIL.n24 VTAIL.n6 3.49141
R194 VTAIL.n104 VTAIL.n86 3.49141
R195 VTAIL.n64 VTAIL.n46 3.49141
R196 VTAIL.n143 VTAIL.n128 2.71565
R197 VTAIL.n23 VTAIL.n8 2.71565
R198 VTAIL.n103 VTAIL.n88 2.71565
R199 VTAIL.n63 VTAIL.n48 2.71565
R200 VTAIL.n140 VTAIL.n139 1.93989
R201 VTAIL.n20 VTAIL.n19 1.93989
R202 VTAIL.n100 VTAIL.n99 1.93989
R203 VTAIL.n60 VTAIL.n59 1.93989
R204 VTAIL.n136 VTAIL.n130 1.16414
R205 VTAIL.n16 VTAIL.n10 1.16414
R206 VTAIL.n96 VTAIL.n90 1.16414
R207 VTAIL.n56 VTAIL.n50 1.16414
R208 VTAIL.n119 VTAIL.n79 1.01343
R209 VTAIL VTAIL.n39 0.800069
R210 VTAIL.n135 VTAIL.n132 0.388379
R211 VTAIL.n15 VTAIL.n12 0.388379
R212 VTAIL.n95 VTAIL.n92 0.388379
R213 VTAIL.n55 VTAIL.n52 0.388379
R214 VTAIL VTAIL.n159 0.213862
R215 VTAIL.n134 VTAIL.n129 0.155672
R216 VTAIL.n141 VTAIL.n129 0.155672
R217 VTAIL.n142 VTAIL.n141 0.155672
R218 VTAIL.n142 VTAIL.n125 0.155672
R219 VTAIL.n149 VTAIL.n125 0.155672
R220 VTAIL.n150 VTAIL.n149 0.155672
R221 VTAIL.n150 VTAIL.n121 0.155672
R222 VTAIL.n157 VTAIL.n121 0.155672
R223 VTAIL.n14 VTAIL.n9 0.155672
R224 VTAIL.n21 VTAIL.n9 0.155672
R225 VTAIL.n22 VTAIL.n21 0.155672
R226 VTAIL.n22 VTAIL.n5 0.155672
R227 VTAIL.n29 VTAIL.n5 0.155672
R228 VTAIL.n30 VTAIL.n29 0.155672
R229 VTAIL.n30 VTAIL.n1 0.155672
R230 VTAIL.n37 VTAIL.n1 0.155672
R231 VTAIL.n117 VTAIL.n81 0.155672
R232 VTAIL.n110 VTAIL.n81 0.155672
R233 VTAIL.n110 VTAIL.n109 0.155672
R234 VTAIL.n109 VTAIL.n85 0.155672
R235 VTAIL.n102 VTAIL.n85 0.155672
R236 VTAIL.n102 VTAIL.n101 0.155672
R237 VTAIL.n101 VTAIL.n89 0.155672
R238 VTAIL.n94 VTAIL.n89 0.155672
R239 VTAIL.n77 VTAIL.n41 0.155672
R240 VTAIL.n70 VTAIL.n41 0.155672
R241 VTAIL.n70 VTAIL.n69 0.155672
R242 VTAIL.n69 VTAIL.n45 0.155672
R243 VTAIL.n62 VTAIL.n45 0.155672
R244 VTAIL.n62 VTAIL.n61 0.155672
R245 VTAIL.n61 VTAIL.n49 0.155672
R246 VTAIL.n54 VTAIL.n49 0.155672
R247 VDD2.n73 VDD2.n39 289.615
R248 VDD2.n34 VDD2.n0 289.615
R249 VDD2.n74 VDD2.n73 185
R250 VDD2.n72 VDD2.n71 185
R251 VDD2.n43 VDD2.n42 185
R252 VDD2.n66 VDD2.n65 185
R253 VDD2.n64 VDD2.n63 185
R254 VDD2.n47 VDD2.n46 185
R255 VDD2.n58 VDD2.n57 185
R256 VDD2.n56 VDD2.n55 185
R257 VDD2.n51 VDD2.n50 185
R258 VDD2.n12 VDD2.n11 185
R259 VDD2.n17 VDD2.n16 185
R260 VDD2.n19 VDD2.n18 185
R261 VDD2.n8 VDD2.n7 185
R262 VDD2.n25 VDD2.n24 185
R263 VDD2.n27 VDD2.n26 185
R264 VDD2.n4 VDD2.n3 185
R265 VDD2.n33 VDD2.n32 185
R266 VDD2.n35 VDD2.n34 185
R267 VDD2.n52 VDD2.t1 147.659
R268 VDD2.n13 VDD2.t0 147.659
R269 VDD2.n73 VDD2.n72 104.615
R270 VDD2.n72 VDD2.n42 104.615
R271 VDD2.n65 VDD2.n42 104.615
R272 VDD2.n65 VDD2.n64 104.615
R273 VDD2.n64 VDD2.n46 104.615
R274 VDD2.n57 VDD2.n46 104.615
R275 VDD2.n57 VDD2.n56 104.615
R276 VDD2.n56 VDD2.n50 104.615
R277 VDD2.n17 VDD2.n11 104.615
R278 VDD2.n18 VDD2.n17 104.615
R279 VDD2.n18 VDD2.n7 104.615
R280 VDD2.n25 VDD2.n7 104.615
R281 VDD2.n26 VDD2.n25 104.615
R282 VDD2.n26 VDD2.n3 104.615
R283 VDD2.n33 VDD2.n3 104.615
R284 VDD2.n34 VDD2.n33 104.615
R285 VDD2.n78 VDD2.n38 81.5322
R286 VDD2.t1 VDD2.n50 52.3082
R287 VDD2.t0 VDD2.n11 52.3082
R288 VDD2.n78 VDD2.n77 49.252
R289 VDD2.n52 VDD2.n51 15.6677
R290 VDD2.n13 VDD2.n12 15.6677
R291 VDD2.n55 VDD2.n54 12.8005
R292 VDD2.n16 VDD2.n15 12.8005
R293 VDD2.n58 VDD2.n49 12.0247
R294 VDD2.n19 VDD2.n10 12.0247
R295 VDD2.n59 VDD2.n47 11.249
R296 VDD2.n20 VDD2.n8 11.249
R297 VDD2.n63 VDD2.n62 10.4732
R298 VDD2.n24 VDD2.n23 10.4732
R299 VDD2.n66 VDD2.n45 9.69747
R300 VDD2.n27 VDD2.n6 9.69747
R301 VDD2.n77 VDD2.n76 9.45567
R302 VDD2.n38 VDD2.n37 9.45567
R303 VDD2.n76 VDD2.n75 9.3005
R304 VDD2.n41 VDD2.n40 9.3005
R305 VDD2.n70 VDD2.n69 9.3005
R306 VDD2.n68 VDD2.n67 9.3005
R307 VDD2.n45 VDD2.n44 9.3005
R308 VDD2.n62 VDD2.n61 9.3005
R309 VDD2.n60 VDD2.n59 9.3005
R310 VDD2.n49 VDD2.n48 9.3005
R311 VDD2.n54 VDD2.n53 9.3005
R312 VDD2.n37 VDD2.n36 9.3005
R313 VDD2.n31 VDD2.n30 9.3005
R314 VDD2.n29 VDD2.n28 9.3005
R315 VDD2.n6 VDD2.n5 9.3005
R316 VDD2.n23 VDD2.n22 9.3005
R317 VDD2.n21 VDD2.n20 9.3005
R318 VDD2.n10 VDD2.n9 9.3005
R319 VDD2.n15 VDD2.n14 9.3005
R320 VDD2.n2 VDD2.n1 9.3005
R321 VDD2.n67 VDD2.n43 8.92171
R322 VDD2.n28 VDD2.n4 8.92171
R323 VDD2.n71 VDD2.n70 8.14595
R324 VDD2.n32 VDD2.n31 8.14595
R325 VDD2.n77 VDD2.n39 7.3702
R326 VDD2.n74 VDD2.n41 7.3702
R327 VDD2.n35 VDD2.n2 7.3702
R328 VDD2.n38 VDD2.n0 7.3702
R329 VDD2.n75 VDD2.n39 6.59444
R330 VDD2.n75 VDD2.n74 6.59444
R331 VDD2.n36 VDD2.n35 6.59444
R332 VDD2.n36 VDD2.n0 6.59444
R333 VDD2.n71 VDD2.n41 5.81868
R334 VDD2.n32 VDD2.n2 5.81868
R335 VDD2.n70 VDD2.n43 5.04292
R336 VDD2.n31 VDD2.n4 5.04292
R337 VDD2.n53 VDD2.n52 4.38565
R338 VDD2.n14 VDD2.n13 4.38565
R339 VDD2.n67 VDD2.n66 4.26717
R340 VDD2.n28 VDD2.n27 4.26717
R341 VDD2.n63 VDD2.n45 3.49141
R342 VDD2.n24 VDD2.n6 3.49141
R343 VDD2.n62 VDD2.n47 2.71565
R344 VDD2.n23 VDD2.n8 2.71565
R345 VDD2.n59 VDD2.n58 1.93989
R346 VDD2.n20 VDD2.n19 1.93989
R347 VDD2.n55 VDD2.n49 1.16414
R348 VDD2.n16 VDD2.n10 1.16414
R349 VDD2.n54 VDD2.n51 0.388379
R350 VDD2.n15 VDD2.n12 0.388379
R351 VDD2 VDD2.n78 0.330241
R352 VDD2.n76 VDD2.n40 0.155672
R353 VDD2.n69 VDD2.n40 0.155672
R354 VDD2.n69 VDD2.n68 0.155672
R355 VDD2.n68 VDD2.n44 0.155672
R356 VDD2.n61 VDD2.n44 0.155672
R357 VDD2.n61 VDD2.n60 0.155672
R358 VDD2.n60 VDD2.n48 0.155672
R359 VDD2.n53 VDD2.n48 0.155672
R360 VDD2.n14 VDD2.n9 0.155672
R361 VDD2.n21 VDD2.n9 0.155672
R362 VDD2.n22 VDD2.n21 0.155672
R363 VDD2.n22 VDD2.n5 0.155672
R364 VDD2.n29 VDD2.n5 0.155672
R365 VDD2.n30 VDD2.n29 0.155672
R366 VDD2.n30 VDD2.n1 0.155672
R367 VDD2.n37 VDD2.n1 0.155672
R368 B.n463 B.n462 585
R369 B.n197 B.n65 585
R370 B.n196 B.n195 585
R371 B.n194 B.n193 585
R372 B.n192 B.n191 585
R373 B.n190 B.n189 585
R374 B.n188 B.n187 585
R375 B.n186 B.n185 585
R376 B.n184 B.n183 585
R377 B.n182 B.n181 585
R378 B.n180 B.n179 585
R379 B.n178 B.n177 585
R380 B.n176 B.n175 585
R381 B.n174 B.n173 585
R382 B.n172 B.n171 585
R383 B.n170 B.n169 585
R384 B.n168 B.n167 585
R385 B.n166 B.n165 585
R386 B.n164 B.n163 585
R387 B.n162 B.n161 585
R388 B.n160 B.n159 585
R389 B.n158 B.n157 585
R390 B.n156 B.n155 585
R391 B.n154 B.n153 585
R392 B.n152 B.n151 585
R393 B.n150 B.n149 585
R394 B.n148 B.n147 585
R395 B.n146 B.n145 585
R396 B.n144 B.n143 585
R397 B.n142 B.n141 585
R398 B.n140 B.n139 585
R399 B.n138 B.n137 585
R400 B.n136 B.n135 585
R401 B.n134 B.n133 585
R402 B.n132 B.n131 585
R403 B.n130 B.n129 585
R404 B.n128 B.n127 585
R405 B.n126 B.n125 585
R406 B.n124 B.n123 585
R407 B.n122 B.n121 585
R408 B.n120 B.n119 585
R409 B.n118 B.n117 585
R410 B.n116 B.n115 585
R411 B.n114 B.n113 585
R412 B.n112 B.n111 585
R413 B.n110 B.n109 585
R414 B.n108 B.n107 585
R415 B.n106 B.n105 585
R416 B.n104 B.n103 585
R417 B.n102 B.n101 585
R418 B.n100 B.n99 585
R419 B.n98 B.n97 585
R420 B.n96 B.n95 585
R421 B.n94 B.n93 585
R422 B.n92 B.n91 585
R423 B.n90 B.n89 585
R424 B.n88 B.n87 585
R425 B.n86 B.n85 585
R426 B.n84 B.n83 585
R427 B.n82 B.n81 585
R428 B.n80 B.n79 585
R429 B.n78 B.n77 585
R430 B.n76 B.n75 585
R431 B.n74 B.n73 585
R432 B.n33 B.n32 585
R433 B.n468 B.n467 585
R434 B.n461 B.n66 585
R435 B.n66 B.n30 585
R436 B.n460 B.n29 585
R437 B.n472 B.n29 585
R438 B.n459 B.n28 585
R439 B.n473 B.n28 585
R440 B.n458 B.n27 585
R441 B.n474 B.n27 585
R442 B.n457 B.n456 585
R443 B.n456 B.n23 585
R444 B.n455 B.n22 585
R445 B.n480 B.n22 585
R446 B.n454 B.n21 585
R447 B.n481 B.n21 585
R448 B.n453 B.n20 585
R449 B.n482 B.n20 585
R450 B.n452 B.n451 585
R451 B.n451 B.n16 585
R452 B.n450 B.n15 585
R453 B.n488 B.n15 585
R454 B.n449 B.n14 585
R455 B.n489 B.n14 585
R456 B.n448 B.n13 585
R457 B.n490 B.n13 585
R458 B.n447 B.n446 585
R459 B.n446 B.n12 585
R460 B.n445 B.n444 585
R461 B.n445 B.n8 585
R462 B.n443 B.n7 585
R463 B.n497 B.n7 585
R464 B.n442 B.n6 585
R465 B.n498 B.n6 585
R466 B.n441 B.n5 585
R467 B.n499 B.n5 585
R468 B.n440 B.n439 585
R469 B.n439 B.n4 585
R470 B.n438 B.n198 585
R471 B.n438 B.n437 585
R472 B.n427 B.n199 585
R473 B.n430 B.n199 585
R474 B.n429 B.n428 585
R475 B.n431 B.n429 585
R476 B.n426 B.n204 585
R477 B.n204 B.n203 585
R478 B.n425 B.n424 585
R479 B.n424 B.n423 585
R480 B.n206 B.n205 585
R481 B.n207 B.n206 585
R482 B.n416 B.n415 585
R483 B.n417 B.n416 585
R484 B.n414 B.n212 585
R485 B.n212 B.n211 585
R486 B.n413 B.n412 585
R487 B.n412 B.n411 585
R488 B.n214 B.n213 585
R489 B.n215 B.n214 585
R490 B.n404 B.n403 585
R491 B.n405 B.n404 585
R492 B.n402 B.n220 585
R493 B.n220 B.n219 585
R494 B.n401 B.n400 585
R495 B.n400 B.n399 585
R496 B.n222 B.n221 585
R497 B.n223 B.n222 585
R498 B.n395 B.n394 585
R499 B.n226 B.n225 585
R500 B.n391 B.n390 585
R501 B.n392 B.n391 585
R502 B.n389 B.n259 585
R503 B.n388 B.n387 585
R504 B.n386 B.n385 585
R505 B.n384 B.n383 585
R506 B.n382 B.n381 585
R507 B.n380 B.n379 585
R508 B.n378 B.n377 585
R509 B.n376 B.n375 585
R510 B.n374 B.n373 585
R511 B.n372 B.n371 585
R512 B.n370 B.n369 585
R513 B.n368 B.n367 585
R514 B.n366 B.n365 585
R515 B.n364 B.n363 585
R516 B.n362 B.n361 585
R517 B.n360 B.n359 585
R518 B.n358 B.n357 585
R519 B.n356 B.n355 585
R520 B.n354 B.n353 585
R521 B.n352 B.n351 585
R522 B.n350 B.n349 585
R523 B.n348 B.n347 585
R524 B.n346 B.n345 585
R525 B.n344 B.n343 585
R526 B.n342 B.n341 585
R527 B.n339 B.n338 585
R528 B.n337 B.n336 585
R529 B.n335 B.n334 585
R530 B.n333 B.n332 585
R531 B.n331 B.n330 585
R532 B.n329 B.n328 585
R533 B.n327 B.n326 585
R534 B.n325 B.n324 585
R535 B.n323 B.n322 585
R536 B.n321 B.n320 585
R537 B.n318 B.n317 585
R538 B.n316 B.n315 585
R539 B.n314 B.n313 585
R540 B.n312 B.n311 585
R541 B.n310 B.n309 585
R542 B.n308 B.n307 585
R543 B.n306 B.n305 585
R544 B.n304 B.n303 585
R545 B.n302 B.n301 585
R546 B.n300 B.n299 585
R547 B.n298 B.n297 585
R548 B.n296 B.n295 585
R549 B.n294 B.n293 585
R550 B.n292 B.n291 585
R551 B.n290 B.n289 585
R552 B.n288 B.n287 585
R553 B.n286 B.n285 585
R554 B.n284 B.n283 585
R555 B.n282 B.n281 585
R556 B.n280 B.n279 585
R557 B.n278 B.n277 585
R558 B.n276 B.n275 585
R559 B.n274 B.n273 585
R560 B.n272 B.n271 585
R561 B.n270 B.n269 585
R562 B.n268 B.n267 585
R563 B.n266 B.n265 585
R564 B.n264 B.n258 585
R565 B.n392 B.n258 585
R566 B.n396 B.n224 585
R567 B.n224 B.n223 585
R568 B.n398 B.n397 585
R569 B.n399 B.n398 585
R570 B.n218 B.n217 585
R571 B.n219 B.n218 585
R572 B.n407 B.n406 585
R573 B.n406 B.n405 585
R574 B.n408 B.n216 585
R575 B.n216 B.n215 585
R576 B.n410 B.n409 585
R577 B.n411 B.n410 585
R578 B.n210 B.n209 585
R579 B.n211 B.n210 585
R580 B.n419 B.n418 585
R581 B.n418 B.n417 585
R582 B.n420 B.n208 585
R583 B.n208 B.n207 585
R584 B.n422 B.n421 585
R585 B.n423 B.n422 585
R586 B.n202 B.n201 585
R587 B.n203 B.n202 585
R588 B.n433 B.n432 585
R589 B.n432 B.n431 585
R590 B.n434 B.n200 585
R591 B.n430 B.n200 585
R592 B.n436 B.n435 585
R593 B.n437 B.n436 585
R594 B.n3 B.n0 585
R595 B.n4 B.n3 585
R596 B.n496 B.n1 585
R597 B.n497 B.n496 585
R598 B.n495 B.n494 585
R599 B.n495 B.n8 585
R600 B.n493 B.n9 585
R601 B.n12 B.n9 585
R602 B.n492 B.n491 585
R603 B.n491 B.n490 585
R604 B.n11 B.n10 585
R605 B.n489 B.n11 585
R606 B.n487 B.n486 585
R607 B.n488 B.n487 585
R608 B.n485 B.n17 585
R609 B.n17 B.n16 585
R610 B.n484 B.n483 585
R611 B.n483 B.n482 585
R612 B.n19 B.n18 585
R613 B.n481 B.n19 585
R614 B.n479 B.n478 585
R615 B.n480 B.n479 585
R616 B.n477 B.n24 585
R617 B.n24 B.n23 585
R618 B.n476 B.n475 585
R619 B.n475 B.n474 585
R620 B.n26 B.n25 585
R621 B.n473 B.n26 585
R622 B.n471 B.n470 585
R623 B.n472 B.n471 585
R624 B.n469 B.n31 585
R625 B.n31 B.n30 585
R626 B.n500 B.n499 585
R627 B.n498 B.n2 585
R628 B.n467 B.n31 521.33
R629 B.n463 B.n66 521.33
R630 B.n258 B.n222 521.33
R631 B.n394 B.n224 521.33
R632 B.n70 B.t6 395.745
R633 B.n67 B.t2 395.745
R634 B.n262 B.t9 395.745
R635 B.n260 B.t13 395.745
R636 B.n465 B.n464 256.663
R637 B.n465 B.n64 256.663
R638 B.n465 B.n63 256.663
R639 B.n465 B.n62 256.663
R640 B.n465 B.n61 256.663
R641 B.n465 B.n60 256.663
R642 B.n465 B.n59 256.663
R643 B.n465 B.n58 256.663
R644 B.n465 B.n57 256.663
R645 B.n465 B.n56 256.663
R646 B.n465 B.n55 256.663
R647 B.n465 B.n54 256.663
R648 B.n465 B.n53 256.663
R649 B.n465 B.n52 256.663
R650 B.n465 B.n51 256.663
R651 B.n465 B.n50 256.663
R652 B.n465 B.n49 256.663
R653 B.n465 B.n48 256.663
R654 B.n465 B.n47 256.663
R655 B.n465 B.n46 256.663
R656 B.n465 B.n45 256.663
R657 B.n465 B.n44 256.663
R658 B.n465 B.n43 256.663
R659 B.n465 B.n42 256.663
R660 B.n465 B.n41 256.663
R661 B.n465 B.n40 256.663
R662 B.n465 B.n39 256.663
R663 B.n465 B.n38 256.663
R664 B.n465 B.n37 256.663
R665 B.n465 B.n36 256.663
R666 B.n465 B.n35 256.663
R667 B.n465 B.n34 256.663
R668 B.n466 B.n465 256.663
R669 B.n393 B.n392 256.663
R670 B.n392 B.n227 256.663
R671 B.n392 B.n228 256.663
R672 B.n392 B.n229 256.663
R673 B.n392 B.n230 256.663
R674 B.n392 B.n231 256.663
R675 B.n392 B.n232 256.663
R676 B.n392 B.n233 256.663
R677 B.n392 B.n234 256.663
R678 B.n392 B.n235 256.663
R679 B.n392 B.n236 256.663
R680 B.n392 B.n237 256.663
R681 B.n392 B.n238 256.663
R682 B.n392 B.n239 256.663
R683 B.n392 B.n240 256.663
R684 B.n392 B.n241 256.663
R685 B.n392 B.n242 256.663
R686 B.n392 B.n243 256.663
R687 B.n392 B.n244 256.663
R688 B.n392 B.n245 256.663
R689 B.n392 B.n246 256.663
R690 B.n392 B.n247 256.663
R691 B.n392 B.n248 256.663
R692 B.n392 B.n249 256.663
R693 B.n392 B.n250 256.663
R694 B.n392 B.n251 256.663
R695 B.n392 B.n252 256.663
R696 B.n392 B.n253 256.663
R697 B.n392 B.n254 256.663
R698 B.n392 B.n255 256.663
R699 B.n392 B.n256 256.663
R700 B.n392 B.n257 256.663
R701 B.n502 B.n501 256.663
R702 B.n67 B.t4 228.738
R703 B.n262 B.t12 228.738
R704 B.n70 B.t7 228.738
R705 B.n260 B.t15 228.738
R706 B.n68 B.t5 204.302
R707 B.n263 B.t11 204.302
R708 B.n71 B.t8 204.3
R709 B.n261 B.t14 204.3
R710 B.n73 B.n33 163.367
R711 B.n77 B.n76 163.367
R712 B.n81 B.n80 163.367
R713 B.n85 B.n84 163.367
R714 B.n89 B.n88 163.367
R715 B.n93 B.n92 163.367
R716 B.n97 B.n96 163.367
R717 B.n101 B.n100 163.367
R718 B.n105 B.n104 163.367
R719 B.n109 B.n108 163.367
R720 B.n113 B.n112 163.367
R721 B.n117 B.n116 163.367
R722 B.n121 B.n120 163.367
R723 B.n125 B.n124 163.367
R724 B.n129 B.n128 163.367
R725 B.n133 B.n132 163.367
R726 B.n137 B.n136 163.367
R727 B.n141 B.n140 163.367
R728 B.n145 B.n144 163.367
R729 B.n149 B.n148 163.367
R730 B.n153 B.n152 163.367
R731 B.n157 B.n156 163.367
R732 B.n161 B.n160 163.367
R733 B.n165 B.n164 163.367
R734 B.n169 B.n168 163.367
R735 B.n173 B.n172 163.367
R736 B.n177 B.n176 163.367
R737 B.n181 B.n180 163.367
R738 B.n185 B.n184 163.367
R739 B.n189 B.n188 163.367
R740 B.n193 B.n192 163.367
R741 B.n195 B.n65 163.367
R742 B.n400 B.n222 163.367
R743 B.n400 B.n220 163.367
R744 B.n404 B.n220 163.367
R745 B.n404 B.n214 163.367
R746 B.n412 B.n214 163.367
R747 B.n412 B.n212 163.367
R748 B.n416 B.n212 163.367
R749 B.n416 B.n206 163.367
R750 B.n424 B.n206 163.367
R751 B.n424 B.n204 163.367
R752 B.n429 B.n204 163.367
R753 B.n429 B.n199 163.367
R754 B.n438 B.n199 163.367
R755 B.n439 B.n438 163.367
R756 B.n439 B.n5 163.367
R757 B.n6 B.n5 163.367
R758 B.n7 B.n6 163.367
R759 B.n445 B.n7 163.367
R760 B.n446 B.n445 163.367
R761 B.n446 B.n13 163.367
R762 B.n14 B.n13 163.367
R763 B.n15 B.n14 163.367
R764 B.n451 B.n15 163.367
R765 B.n451 B.n20 163.367
R766 B.n21 B.n20 163.367
R767 B.n22 B.n21 163.367
R768 B.n456 B.n22 163.367
R769 B.n456 B.n27 163.367
R770 B.n28 B.n27 163.367
R771 B.n29 B.n28 163.367
R772 B.n66 B.n29 163.367
R773 B.n391 B.n226 163.367
R774 B.n391 B.n259 163.367
R775 B.n387 B.n386 163.367
R776 B.n383 B.n382 163.367
R777 B.n379 B.n378 163.367
R778 B.n375 B.n374 163.367
R779 B.n371 B.n370 163.367
R780 B.n367 B.n366 163.367
R781 B.n363 B.n362 163.367
R782 B.n359 B.n358 163.367
R783 B.n355 B.n354 163.367
R784 B.n351 B.n350 163.367
R785 B.n347 B.n346 163.367
R786 B.n343 B.n342 163.367
R787 B.n338 B.n337 163.367
R788 B.n334 B.n333 163.367
R789 B.n330 B.n329 163.367
R790 B.n326 B.n325 163.367
R791 B.n322 B.n321 163.367
R792 B.n317 B.n316 163.367
R793 B.n313 B.n312 163.367
R794 B.n309 B.n308 163.367
R795 B.n305 B.n304 163.367
R796 B.n301 B.n300 163.367
R797 B.n297 B.n296 163.367
R798 B.n293 B.n292 163.367
R799 B.n289 B.n288 163.367
R800 B.n285 B.n284 163.367
R801 B.n281 B.n280 163.367
R802 B.n277 B.n276 163.367
R803 B.n273 B.n272 163.367
R804 B.n269 B.n268 163.367
R805 B.n265 B.n258 163.367
R806 B.n398 B.n224 163.367
R807 B.n398 B.n218 163.367
R808 B.n406 B.n218 163.367
R809 B.n406 B.n216 163.367
R810 B.n410 B.n216 163.367
R811 B.n410 B.n210 163.367
R812 B.n418 B.n210 163.367
R813 B.n418 B.n208 163.367
R814 B.n422 B.n208 163.367
R815 B.n422 B.n202 163.367
R816 B.n432 B.n202 163.367
R817 B.n432 B.n200 163.367
R818 B.n436 B.n200 163.367
R819 B.n436 B.n3 163.367
R820 B.n500 B.n3 163.367
R821 B.n496 B.n2 163.367
R822 B.n496 B.n495 163.367
R823 B.n495 B.n9 163.367
R824 B.n491 B.n9 163.367
R825 B.n491 B.n11 163.367
R826 B.n487 B.n11 163.367
R827 B.n487 B.n17 163.367
R828 B.n483 B.n17 163.367
R829 B.n483 B.n19 163.367
R830 B.n479 B.n19 163.367
R831 B.n479 B.n24 163.367
R832 B.n475 B.n24 163.367
R833 B.n475 B.n26 163.367
R834 B.n471 B.n26 163.367
R835 B.n471 B.n31 163.367
R836 B.n392 B.n223 107.802
R837 B.n465 B.n30 107.802
R838 B.n467 B.n466 71.676
R839 B.n73 B.n34 71.676
R840 B.n77 B.n35 71.676
R841 B.n81 B.n36 71.676
R842 B.n85 B.n37 71.676
R843 B.n89 B.n38 71.676
R844 B.n93 B.n39 71.676
R845 B.n97 B.n40 71.676
R846 B.n101 B.n41 71.676
R847 B.n105 B.n42 71.676
R848 B.n109 B.n43 71.676
R849 B.n113 B.n44 71.676
R850 B.n117 B.n45 71.676
R851 B.n121 B.n46 71.676
R852 B.n125 B.n47 71.676
R853 B.n129 B.n48 71.676
R854 B.n133 B.n49 71.676
R855 B.n137 B.n50 71.676
R856 B.n141 B.n51 71.676
R857 B.n145 B.n52 71.676
R858 B.n149 B.n53 71.676
R859 B.n153 B.n54 71.676
R860 B.n157 B.n55 71.676
R861 B.n161 B.n56 71.676
R862 B.n165 B.n57 71.676
R863 B.n169 B.n58 71.676
R864 B.n173 B.n59 71.676
R865 B.n177 B.n60 71.676
R866 B.n181 B.n61 71.676
R867 B.n185 B.n62 71.676
R868 B.n189 B.n63 71.676
R869 B.n193 B.n64 71.676
R870 B.n464 B.n65 71.676
R871 B.n464 B.n463 71.676
R872 B.n195 B.n64 71.676
R873 B.n192 B.n63 71.676
R874 B.n188 B.n62 71.676
R875 B.n184 B.n61 71.676
R876 B.n180 B.n60 71.676
R877 B.n176 B.n59 71.676
R878 B.n172 B.n58 71.676
R879 B.n168 B.n57 71.676
R880 B.n164 B.n56 71.676
R881 B.n160 B.n55 71.676
R882 B.n156 B.n54 71.676
R883 B.n152 B.n53 71.676
R884 B.n148 B.n52 71.676
R885 B.n144 B.n51 71.676
R886 B.n140 B.n50 71.676
R887 B.n136 B.n49 71.676
R888 B.n132 B.n48 71.676
R889 B.n128 B.n47 71.676
R890 B.n124 B.n46 71.676
R891 B.n120 B.n45 71.676
R892 B.n116 B.n44 71.676
R893 B.n112 B.n43 71.676
R894 B.n108 B.n42 71.676
R895 B.n104 B.n41 71.676
R896 B.n100 B.n40 71.676
R897 B.n96 B.n39 71.676
R898 B.n92 B.n38 71.676
R899 B.n88 B.n37 71.676
R900 B.n84 B.n36 71.676
R901 B.n80 B.n35 71.676
R902 B.n76 B.n34 71.676
R903 B.n466 B.n33 71.676
R904 B.n394 B.n393 71.676
R905 B.n259 B.n227 71.676
R906 B.n386 B.n228 71.676
R907 B.n382 B.n229 71.676
R908 B.n378 B.n230 71.676
R909 B.n374 B.n231 71.676
R910 B.n370 B.n232 71.676
R911 B.n366 B.n233 71.676
R912 B.n362 B.n234 71.676
R913 B.n358 B.n235 71.676
R914 B.n354 B.n236 71.676
R915 B.n350 B.n237 71.676
R916 B.n346 B.n238 71.676
R917 B.n342 B.n239 71.676
R918 B.n337 B.n240 71.676
R919 B.n333 B.n241 71.676
R920 B.n329 B.n242 71.676
R921 B.n325 B.n243 71.676
R922 B.n321 B.n244 71.676
R923 B.n316 B.n245 71.676
R924 B.n312 B.n246 71.676
R925 B.n308 B.n247 71.676
R926 B.n304 B.n248 71.676
R927 B.n300 B.n249 71.676
R928 B.n296 B.n250 71.676
R929 B.n292 B.n251 71.676
R930 B.n288 B.n252 71.676
R931 B.n284 B.n253 71.676
R932 B.n280 B.n254 71.676
R933 B.n276 B.n255 71.676
R934 B.n272 B.n256 71.676
R935 B.n268 B.n257 71.676
R936 B.n393 B.n226 71.676
R937 B.n387 B.n227 71.676
R938 B.n383 B.n228 71.676
R939 B.n379 B.n229 71.676
R940 B.n375 B.n230 71.676
R941 B.n371 B.n231 71.676
R942 B.n367 B.n232 71.676
R943 B.n363 B.n233 71.676
R944 B.n359 B.n234 71.676
R945 B.n355 B.n235 71.676
R946 B.n351 B.n236 71.676
R947 B.n347 B.n237 71.676
R948 B.n343 B.n238 71.676
R949 B.n338 B.n239 71.676
R950 B.n334 B.n240 71.676
R951 B.n330 B.n241 71.676
R952 B.n326 B.n242 71.676
R953 B.n322 B.n243 71.676
R954 B.n317 B.n244 71.676
R955 B.n313 B.n245 71.676
R956 B.n309 B.n246 71.676
R957 B.n305 B.n247 71.676
R958 B.n301 B.n248 71.676
R959 B.n297 B.n249 71.676
R960 B.n293 B.n250 71.676
R961 B.n289 B.n251 71.676
R962 B.n285 B.n252 71.676
R963 B.n281 B.n253 71.676
R964 B.n277 B.n254 71.676
R965 B.n273 B.n255 71.676
R966 B.n269 B.n256 71.676
R967 B.n265 B.n257 71.676
R968 B.n501 B.n500 71.676
R969 B.n501 B.n2 71.676
R970 B.n72 B.n71 59.5399
R971 B.n69 B.n68 59.5399
R972 B.n319 B.n263 59.5399
R973 B.n340 B.n261 59.5399
R974 B.n399 B.n223 58.6442
R975 B.n399 B.n219 58.6442
R976 B.n405 B.n219 58.6442
R977 B.n405 B.n215 58.6442
R978 B.n411 B.n215 58.6442
R979 B.n417 B.n211 58.6442
R980 B.n417 B.n207 58.6442
R981 B.n423 B.n207 58.6442
R982 B.n423 B.n203 58.6442
R983 B.n431 B.n203 58.6442
R984 B.n431 B.n430 58.6442
R985 B.n437 B.n4 58.6442
R986 B.n499 B.n4 58.6442
R987 B.n499 B.n498 58.6442
R988 B.n498 B.n497 58.6442
R989 B.n497 B.n8 58.6442
R990 B.n490 B.n12 58.6442
R991 B.n490 B.n489 58.6442
R992 B.n489 B.n488 58.6442
R993 B.n488 B.n16 58.6442
R994 B.n482 B.n16 58.6442
R995 B.n482 B.n481 58.6442
R996 B.n480 B.n23 58.6442
R997 B.n474 B.n23 58.6442
R998 B.n474 B.n473 58.6442
R999 B.n473 B.n472 58.6442
R1000 B.n472 B.n30 58.6442
R1001 B.n437 B.t1 56.0569
R1002 B.t0 B.n8 56.0569
R1003 B.t10 B.n211 50.8825
R1004 B.n481 B.t3 50.8825
R1005 B.n396 B.n395 33.8737
R1006 B.n264 B.n221 33.8737
R1007 B.n462 B.n461 33.8737
R1008 B.n469 B.n468 33.8737
R1009 B.n71 B.n70 24.4369
R1010 B.n68 B.n67 24.4369
R1011 B.n263 B.n262 24.4369
R1012 B.n261 B.n260 24.4369
R1013 B B.n502 18.0485
R1014 B.n397 B.n396 10.6151
R1015 B.n397 B.n217 10.6151
R1016 B.n407 B.n217 10.6151
R1017 B.n408 B.n407 10.6151
R1018 B.n409 B.n408 10.6151
R1019 B.n409 B.n209 10.6151
R1020 B.n419 B.n209 10.6151
R1021 B.n420 B.n419 10.6151
R1022 B.n421 B.n420 10.6151
R1023 B.n421 B.n201 10.6151
R1024 B.n433 B.n201 10.6151
R1025 B.n434 B.n433 10.6151
R1026 B.n435 B.n434 10.6151
R1027 B.n435 B.n0 10.6151
R1028 B.n395 B.n225 10.6151
R1029 B.n390 B.n225 10.6151
R1030 B.n390 B.n389 10.6151
R1031 B.n389 B.n388 10.6151
R1032 B.n388 B.n385 10.6151
R1033 B.n385 B.n384 10.6151
R1034 B.n384 B.n381 10.6151
R1035 B.n381 B.n380 10.6151
R1036 B.n380 B.n377 10.6151
R1037 B.n377 B.n376 10.6151
R1038 B.n376 B.n373 10.6151
R1039 B.n373 B.n372 10.6151
R1040 B.n372 B.n369 10.6151
R1041 B.n369 B.n368 10.6151
R1042 B.n368 B.n365 10.6151
R1043 B.n365 B.n364 10.6151
R1044 B.n364 B.n361 10.6151
R1045 B.n361 B.n360 10.6151
R1046 B.n360 B.n357 10.6151
R1047 B.n357 B.n356 10.6151
R1048 B.n356 B.n353 10.6151
R1049 B.n353 B.n352 10.6151
R1050 B.n352 B.n349 10.6151
R1051 B.n349 B.n348 10.6151
R1052 B.n348 B.n345 10.6151
R1053 B.n345 B.n344 10.6151
R1054 B.n344 B.n341 10.6151
R1055 B.n339 B.n336 10.6151
R1056 B.n336 B.n335 10.6151
R1057 B.n335 B.n332 10.6151
R1058 B.n332 B.n331 10.6151
R1059 B.n331 B.n328 10.6151
R1060 B.n328 B.n327 10.6151
R1061 B.n327 B.n324 10.6151
R1062 B.n324 B.n323 10.6151
R1063 B.n323 B.n320 10.6151
R1064 B.n318 B.n315 10.6151
R1065 B.n315 B.n314 10.6151
R1066 B.n314 B.n311 10.6151
R1067 B.n311 B.n310 10.6151
R1068 B.n310 B.n307 10.6151
R1069 B.n307 B.n306 10.6151
R1070 B.n306 B.n303 10.6151
R1071 B.n303 B.n302 10.6151
R1072 B.n302 B.n299 10.6151
R1073 B.n299 B.n298 10.6151
R1074 B.n298 B.n295 10.6151
R1075 B.n295 B.n294 10.6151
R1076 B.n294 B.n291 10.6151
R1077 B.n291 B.n290 10.6151
R1078 B.n290 B.n287 10.6151
R1079 B.n287 B.n286 10.6151
R1080 B.n286 B.n283 10.6151
R1081 B.n283 B.n282 10.6151
R1082 B.n282 B.n279 10.6151
R1083 B.n279 B.n278 10.6151
R1084 B.n278 B.n275 10.6151
R1085 B.n275 B.n274 10.6151
R1086 B.n274 B.n271 10.6151
R1087 B.n271 B.n270 10.6151
R1088 B.n270 B.n267 10.6151
R1089 B.n267 B.n266 10.6151
R1090 B.n266 B.n264 10.6151
R1091 B.n401 B.n221 10.6151
R1092 B.n402 B.n401 10.6151
R1093 B.n403 B.n402 10.6151
R1094 B.n403 B.n213 10.6151
R1095 B.n413 B.n213 10.6151
R1096 B.n414 B.n413 10.6151
R1097 B.n415 B.n414 10.6151
R1098 B.n415 B.n205 10.6151
R1099 B.n425 B.n205 10.6151
R1100 B.n426 B.n425 10.6151
R1101 B.n428 B.n426 10.6151
R1102 B.n428 B.n427 10.6151
R1103 B.n427 B.n198 10.6151
R1104 B.n440 B.n198 10.6151
R1105 B.n441 B.n440 10.6151
R1106 B.n442 B.n441 10.6151
R1107 B.n443 B.n442 10.6151
R1108 B.n444 B.n443 10.6151
R1109 B.n447 B.n444 10.6151
R1110 B.n448 B.n447 10.6151
R1111 B.n449 B.n448 10.6151
R1112 B.n450 B.n449 10.6151
R1113 B.n452 B.n450 10.6151
R1114 B.n453 B.n452 10.6151
R1115 B.n454 B.n453 10.6151
R1116 B.n455 B.n454 10.6151
R1117 B.n457 B.n455 10.6151
R1118 B.n458 B.n457 10.6151
R1119 B.n459 B.n458 10.6151
R1120 B.n460 B.n459 10.6151
R1121 B.n461 B.n460 10.6151
R1122 B.n494 B.n1 10.6151
R1123 B.n494 B.n493 10.6151
R1124 B.n493 B.n492 10.6151
R1125 B.n492 B.n10 10.6151
R1126 B.n486 B.n10 10.6151
R1127 B.n486 B.n485 10.6151
R1128 B.n485 B.n484 10.6151
R1129 B.n484 B.n18 10.6151
R1130 B.n478 B.n18 10.6151
R1131 B.n478 B.n477 10.6151
R1132 B.n477 B.n476 10.6151
R1133 B.n476 B.n25 10.6151
R1134 B.n470 B.n25 10.6151
R1135 B.n470 B.n469 10.6151
R1136 B.n468 B.n32 10.6151
R1137 B.n74 B.n32 10.6151
R1138 B.n75 B.n74 10.6151
R1139 B.n78 B.n75 10.6151
R1140 B.n79 B.n78 10.6151
R1141 B.n82 B.n79 10.6151
R1142 B.n83 B.n82 10.6151
R1143 B.n86 B.n83 10.6151
R1144 B.n87 B.n86 10.6151
R1145 B.n90 B.n87 10.6151
R1146 B.n91 B.n90 10.6151
R1147 B.n94 B.n91 10.6151
R1148 B.n95 B.n94 10.6151
R1149 B.n98 B.n95 10.6151
R1150 B.n99 B.n98 10.6151
R1151 B.n102 B.n99 10.6151
R1152 B.n103 B.n102 10.6151
R1153 B.n106 B.n103 10.6151
R1154 B.n107 B.n106 10.6151
R1155 B.n110 B.n107 10.6151
R1156 B.n111 B.n110 10.6151
R1157 B.n114 B.n111 10.6151
R1158 B.n115 B.n114 10.6151
R1159 B.n118 B.n115 10.6151
R1160 B.n119 B.n118 10.6151
R1161 B.n122 B.n119 10.6151
R1162 B.n123 B.n122 10.6151
R1163 B.n127 B.n126 10.6151
R1164 B.n130 B.n127 10.6151
R1165 B.n131 B.n130 10.6151
R1166 B.n134 B.n131 10.6151
R1167 B.n135 B.n134 10.6151
R1168 B.n138 B.n135 10.6151
R1169 B.n139 B.n138 10.6151
R1170 B.n142 B.n139 10.6151
R1171 B.n143 B.n142 10.6151
R1172 B.n147 B.n146 10.6151
R1173 B.n150 B.n147 10.6151
R1174 B.n151 B.n150 10.6151
R1175 B.n154 B.n151 10.6151
R1176 B.n155 B.n154 10.6151
R1177 B.n158 B.n155 10.6151
R1178 B.n159 B.n158 10.6151
R1179 B.n162 B.n159 10.6151
R1180 B.n163 B.n162 10.6151
R1181 B.n166 B.n163 10.6151
R1182 B.n167 B.n166 10.6151
R1183 B.n170 B.n167 10.6151
R1184 B.n171 B.n170 10.6151
R1185 B.n174 B.n171 10.6151
R1186 B.n175 B.n174 10.6151
R1187 B.n178 B.n175 10.6151
R1188 B.n179 B.n178 10.6151
R1189 B.n182 B.n179 10.6151
R1190 B.n183 B.n182 10.6151
R1191 B.n186 B.n183 10.6151
R1192 B.n187 B.n186 10.6151
R1193 B.n190 B.n187 10.6151
R1194 B.n191 B.n190 10.6151
R1195 B.n194 B.n191 10.6151
R1196 B.n196 B.n194 10.6151
R1197 B.n197 B.n196 10.6151
R1198 B.n462 B.n197 10.6151
R1199 B.n341 B.n340 8.74196
R1200 B.n319 B.n318 8.74196
R1201 B.n123 B.n72 8.74196
R1202 B.n146 B.n69 8.74196
R1203 B.n502 B.n0 8.11757
R1204 B.n502 B.n1 8.11757
R1205 B.n411 B.t10 7.76216
R1206 B.t3 B.n480 7.76216
R1207 B.n430 B.t1 2.58772
R1208 B.n12 B.t0 2.58772
R1209 B.n340 B.n339 1.87367
R1210 B.n320 B.n319 1.87367
R1211 B.n126 B.n72 1.87367
R1212 B.n143 B.n69 1.87367
R1213 VP.n0 VP.t1 433.661
R1214 VP.n0 VP.t0 396.858
R1215 VP VP.n0 0.0516364
R1216 VDD1.n34 VDD1.n0 289.615
R1217 VDD1.n73 VDD1.n39 289.615
R1218 VDD1.n35 VDD1.n34 185
R1219 VDD1.n33 VDD1.n32 185
R1220 VDD1.n4 VDD1.n3 185
R1221 VDD1.n27 VDD1.n26 185
R1222 VDD1.n25 VDD1.n24 185
R1223 VDD1.n8 VDD1.n7 185
R1224 VDD1.n19 VDD1.n18 185
R1225 VDD1.n17 VDD1.n16 185
R1226 VDD1.n12 VDD1.n11 185
R1227 VDD1.n51 VDD1.n50 185
R1228 VDD1.n56 VDD1.n55 185
R1229 VDD1.n58 VDD1.n57 185
R1230 VDD1.n47 VDD1.n46 185
R1231 VDD1.n64 VDD1.n63 185
R1232 VDD1.n66 VDD1.n65 185
R1233 VDD1.n43 VDD1.n42 185
R1234 VDD1.n72 VDD1.n71 185
R1235 VDD1.n74 VDD1.n73 185
R1236 VDD1.n13 VDD1.t0 147.659
R1237 VDD1.n52 VDD1.t1 147.659
R1238 VDD1.n34 VDD1.n33 104.615
R1239 VDD1.n33 VDD1.n3 104.615
R1240 VDD1.n26 VDD1.n3 104.615
R1241 VDD1.n26 VDD1.n25 104.615
R1242 VDD1.n25 VDD1.n7 104.615
R1243 VDD1.n18 VDD1.n7 104.615
R1244 VDD1.n18 VDD1.n17 104.615
R1245 VDD1.n17 VDD1.n11 104.615
R1246 VDD1.n56 VDD1.n50 104.615
R1247 VDD1.n57 VDD1.n56 104.615
R1248 VDD1.n57 VDD1.n46 104.615
R1249 VDD1.n64 VDD1.n46 104.615
R1250 VDD1.n65 VDD1.n64 104.615
R1251 VDD1.n65 VDD1.n42 104.615
R1252 VDD1.n72 VDD1.n42 104.615
R1253 VDD1.n73 VDD1.n72 104.615
R1254 VDD1 VDD1.n77 82.3285
R1255 VDD1.t0 VDD1.n11 52.3082
R1256 VDD1.t1 VDD1.n50 52.3082
R1257 VDD1 VDD1.n38 49.5818
R1258 VDD1.n13 VDD1.n12 15.6677
R1259 VDD1.n52 VDD1.n51 15.6677
R1260 VDD1.n16 VDD1.n15 12.8005
R1261 VDD1.n55 VDD1.n54 12.8005
R1262 VDD1.n19 VDD1.n10 12.0247
R1263 VDD1.n58 VDD1.n49 12.0247
R1264 VDD1.n20 VDD1.n8 11.249
R1265 VDD1.n59 VDD1.n47 11.249
R1266 VDD1.n24 VDD1.n23 10.4732
R1267 VDD1.n63 VDD1.n62 10.4732
R1268 VDD1.n27 VDD1.n6 9.69747
R1269 VDD1.n66 VDD1.n45 9.69747
R1270 VDD1.n38 VDD1.n37 9.45567
R1271 VDD1.n77 VDD1.n76 9.45567
R1272 VDD1.n37 VDD1.n36 9.3005
R1273 VDD1.n2 VDD1.n1 9.3005
R1274 VDD1.n31 VDD1.n30 9.3005
R1275 VDD1.n29 VDD1.n28 9.3005
R1276 VDD1.n6 VDD1.n5 9.3005
R1277 VDD1.n23 VDD1.n22 9.3005
R1278 VDD1.n21 VDD1.n20 9.3005
R1279 VDD1.n10 VDD1.n9 9.3005
R1280 VDD1.n15 VDD1.n14 9.3005
R1281 VDD1.n76 VDD1.n75 9.3005
R1282 VDD1.n70 VDD1.n69 9.3005
R1283 VDD1.n68 VDD1.n67 9.3005
R1284 VDD1.n45 VDD1.n44 9.3005
R1285 VDD1.n62 VDD1.n61 9.3005
R1286 VDD1.n60 VDD1.n59 9.3005
R1287 VDD1.n49 VDD1.n48 9.3005
R1288 VDD1.n54 VDD1.n53 9.3005
R1289 VDD1.n41 VDD1.n40 9.3005
R1290 VDD1.n28 VDD1.n4 8.92171
R1291 VDD1.n67 VDD1.n43 8.92171
R1292 VDD1.n32 VDD1.n31 8.14595
R1293 VDD1.n71 VDD1.n70 8.14595
R1294 VDD1.n38 VDD1.n0 7.3702
R1295 VDD1.n35 VDD1.n2 7.3702
R1296 VDD1.n74 VDD1.n41 7.3702
R1297 VDD1.n77 VDD1.n39 7.3702
R1298 VDD1.n36 VDD1.n0 6.59444
R1299 VDD1.n36 VDD1.n35 6.59444
R1300 VDD1.n75 VDD1.n74 6.59444
R1301 VDD1.n75 VDD1.n39 6.59444
R1302 VDD1.n32 VDD1.n2 5.81868
R1303 VDD1.n71 VDD1.n41 5.81868
R1304 VDD1.n31 VDD1.n4 5.04292
R1305 VDD1.n70 VDD1.n43 5.04292
R1306 VDD1.n14 VDD1.n13 4.38565
R1307 VDD1.n53 VDD1.n52 4.38565
R1308 VDD1.n28 VDD1.n27 4.26717
R1309 VDD1.n67 VDD1.n66 4.26717
R1310 VDD1.n24 VDD1.n6 3.49141
R1311 VDD1.n63 VDD1.n45 3.49141
R1312 VDD1.n23 VDD1.n8 2.71565
R1313 VDD1.n62 VDD1.n47 2.71565
R1314 VDD1.n20 VDD1.n19 1.93989
R1315 VDD1.n59 VDD1.n58 1.93989
R1316 VDD1.n16 VDD1.n10 1.16414
R1317 VDD1.n55 VDD1.n49 1.16414
R1318 VDD1.n15 VDD1.n12 0.388379
R1319 VDD1.n54 VDD1.n51 0.388379
R1320 VDD1.n37 VDD1.n1 0.155672
R1321 VDD1.n30 VDD1.n1 0.155672
R1322 VDD1.n30 VDD1.n29 0.155672
R1323 VDD1.n29 VDD1.n5 0.155672
R1324 VDD1.n22 VDD1.n5 0.155672
R1325 VDD1.n22 VDD1.n21 0.155672
R1326 VDD1.n21 VDD1.n9 0.155672
R1327 VDD1.n14 VDD1.n9 0.155672
R1328 VDD1.n53 VDD1.n48 0.155672
R1329 VDD1.n60 VDD1.n48 0.155672
R1330 VDD1.n61 VDD1.n60 0.155672
R1331 VDD1.n61 VDD1.n44 0.155672
R1332 VDD1.n68 VDD1.n44 0.155672
R1333 VDD1.n69 VDD1.n68 0.155672
R1334 VDD1.n69 VDD1.n40 0.155672
R1335 VDD1.n76 VDD1.n40 0.155672
C0 VP VTAIL 1.18836f
C1 VDD1 VDD2 0.483798f
C2 VN VDD1 0.149027f
C3 VP VDD2 0.26426f
C4 VP VN 3.82271f
C5 VDD2 VTAIL 3.86773f
C6 VN VTAIL 1.17399f
C7 VP VDD1 1.55994f
C8 VDD1 VTAIL 3.82928f
C9 VN VDD2 1.44727f
C10 VDD2 B 3.006809f
C11 VDD1 B 4.49208f
C12 VTAIL B 4.744366f
C13 VN B 6.35704f
C14 VP B 3.993592f
C15 VDD1.n0 B 0.021554f
C16 VDD1.n1 B 0.014632f
C17 VDD1.n2 B 0.007863f
C18 VDD1.n3 B 0.018585f
C19 VDD1.n4 B 0.008325f
C20 VDD1.n5 B 0.014632f
C21 VDD1.n6 B 0.007863f
C22 VDD1.n7 B 0.018585f
C23 VDD1.n8 B 0.008325f
C24 VDD1.n9 B 0.014632f
C25 VDD1.n10 B 0.007863f
C26 VDD1.n11 B 0.013939f
C27 VDD1.n12 B 0.010979f
C28 VDD1.t0 B 0.030294f
C29 VDD1.n13 B 0.067834f
C30 VDD1.n14 B 0.446281f
C31 VDD1.n15 B 0.007863f
C32 VDD1.n16 B 0.008325f
C33 VDD1.n17 B 0.018585f
C34 VDD1.n18 B 0.018585f
C35 VDD1.n19 B 0.008325f
C36 VDD1.n20 B 0.007863f
C37 VDD1.n21 B 0.014632f
C38 VDD1.n22 B 0.014632f
C39 VDD1.n23 B 0.007863f
C40 VDD1.n24 B 0.008325f
C41 VDD1.n25 B 0.018585f
C42 VDD1.n26 B 0.018585f
C43 VDD1.n27 B 0.008325f
C44 VDD1.n28 B 0.007863f
C45 VDD1.n29 B 0.014632f
C46 VDD1.n30 B 0.014632f
C47 VDD1.n31 B 0.007863f
C48 VDD1.n32 B 0.008325f
C49 VDD1.n33 B 0.018585f
C50 VDD1.n34 B 0.041979f
C51 VDD1.n35 B 0.008325f
C52 VDD1.n36 B 0.007863f
C53 VDD1.n37 B 0.034222f
C54 VDD1.n38 B 0.034073f
C55 VDD1.n39 B 0.021554f
C56 VDD1.n40 B 0.014632f
C57 VDD1.n41 B 0.007863f
C58 VDD1.n42 B 0.018585f
C59 VDD1.n43 B 0.008325f
C60 VDD1.n44 B 0.014632f
C61 VDD1.n45 B 0.007863f
C62 VDD1.n46 B 0.018585f
C63 VDD1.n47 B 0.008325f
C64 VDD1.n48 B 0.014632f
C65 VDD1.n49 B 0.007863f
C66 VDD1.n50 B 0.013939f
C67 VDD1.n51 B 0.010979f
C68 VDD1.t1 B 0.030294f
C69 VDD1.n52 B 0.067834f
C70 VDD1.n53 B 0.446281f
C71 VDD1.n54 B 0.007863f
C72 VDD1.n55 B 0.008325f
C73 VDD1.n56 B 0.018585f
C74 VDD1.n57 B 0.018585f
C75 VDD1.n58 B 0.008325f
C76 VDD1.n59 B 0.007863f
C77 VDD1.n60 B 0.014632f
C78 VDD1.n61 B 0.014632f
C79 VDD1.n62 B 0.007863f
C80 VDD1.n63 B 0.008325f
C81 VDD1.n64 B 0.018585f
C82 VDD1.n65 B 0.018585f
C83 VDD1.n66 B 0.008325f
C84 VDD1.n67 B 0.007863f
C85 VDD1.n68 B 0.014632f
C86 VDD1.n69 B 0.014632f
C87 VDD1.n70 B 0.007863f
C88 VDD1.n71 B 0.008325f
C89 VDD1.n72 B 0.018585f
C90 VDD1.n73 B 0.041979f
C91 VDD1.n74 B 0.008325f
C92 VDD1.n75 B 0.007863f
C93 VDD1.n76 B 0.034222f
C94 VDD1.n77 B 0.301981f
C95 VP.t1 B 0.817433f
C96 VP.t0 B 0.718448f
C97 VP.n0 B 2.2491f
C98 VDD2.n0 B 0.022441f
C99 VDD2.n1 B 0.015234f
C100 VDD2.n2 B 0.008186f
C101 VDD2.n3 B 0.019349f
C102 VDD2.n4 B 0.008668f
C103 VDD2.n5 B 0.015234f
C104 VDD2.n6 B 0.008186f
C105 VDD2.n7 B 0.019349f
C106 VDD2.n8 B 0.008668f
C107 VDD2.n9 B 0.015234f
C108 VDD2.n10 B 0.008186f
C109 VDD2.n11 B 0.014512f
C110 VDD2.n12 B 0.01143f
C111 VDD2.t0 B 0.03154f
C112 VDD2.n13 B 0.070623f
C113 VDD2.n14 B 0.464633f
C114 VDD2.n15 B 0.008186f
C115 VDD2.n16 B 0.008668f
C116 VDD2.n17 B 0.019349f
C117 VDD2.n18 B 0.019349f
C118 VDD2.n19 B 0.008668f
C119 VDD2.n20 B 0.008186f
C120 VDD2.n21 B 0.015234f
C121 VDD2.n22 B 0.015234f
C122 VDD2.n23 B 0.008186f
C123 VDD2.n24 B 0.008668f
C124 VDD2.n25 B 0.019349f
C125 VDD2.n26 B 0.019349f
C126 VDD2.n27 B 0.008668f
C127 VDD2.n28 B 0.008186f
C128 VDD2.n29 B 0.015234f
C129 VDD2.n30 B 0.015234f
C130 VDD2.n31 B 0.008186f
C131 VDD2.n32 B 0.008668f
C132 VDD2.n33 B 0.019349f
C133 VDD2.n34 B 0.043705f
C134 VDD2.n35 B 0.008668f
C135 VDD2.n36 B 0.008186f
C136 VDD2.n37 B 0.035629f
C137 VDD2.n38 B 0.294875f
C138 VDD2.n39 B 0.022441f
C139 VDD2.n40 B 0.015234f
C140 VDD2.n41 B 0.008186f
C141 VDD2.n42 B 0.019349f
C142 VDD2.n43 B 0.008668f
C143 VDD2.n44 B 0.015234f
C144 VDD2.n45 B 0.008186f
C145 VDD2.n46 B 0.019349f
C146 VDD2.n47 B 0.008668f
C147 VDD2.n48 B 0.015234f
C148 VDD2.n49 B 0.008186f
C149 VDD2.n50 B 0.014512f
C150 VDD2.n51 B 0.01143f
C151 VDD2.t1 B 0.03154f
C152 VDD2.n52 B 0.070623f
C153 VDD2.n53 B 0.464633f
C154 VDD2.n54 B 0.008186f
C155 VDD2.n55 B 0.008668f
C156 VDD2.n56 B 0.019349f
C157 VDD2.n57 B 0.019349f
C158 VDD2.n58 B 0.008668f
C159 VDD2.n59 B 0.008186f
C160 VDD2.n60 B 0.015234f
C161 VDD2.n61 B 0.015234f
C162 VDD2.n62 B 0.008186f
C163 VDD2.n63 B 0.008668f
C164 VDD2.n64 B 0.019349f
C165 VDD2.n65 B 0.019349f
C166 VDD2.n66 B 0.008668f
C167 VDD2.n67 B 0.008186f
C168 VDD2.n68 B 0.015234f
C169 VDD2.n69 B 0.015234f
C170 VDD2.n70 B 0.008186f
C171 VDD2.n71 B 0.008668f
C172 VDD2.n72 B 0.019349f
C173 VDD2.n73 B 0.043705f
C174 VDD2.n74 B 0.008668f
C175 VDD2.n75 B 0.008186f
C176 VDD2.n76 B 0.035629f
C177 VDD2.n77 B 0.03517f
C178 VDD2.n78 B 1.36746f
C179 VTAIL.n0 B 0.024396f
C180 VTAIL.n1 B 0.016562f
C181 VTAIL.n2 B 0.0089f
C182 VTAIL.n3 B 0.021035f
C183 VTAIL.n4 B 0.009423f
C184 VTAIL.n5 B 0.016562f
C185 VTAIL.n6 B 0.0089f
C186 VTAIL.n7 B 0.021035f
C187 VTAIL.n8 B 0.009423f
C188 VTAIL.n9 B 0.016562f
C189 VTAIL.n10 B 0.0089f
C190 VTAIL.n11 B 0.015777f
C191 VTAIL.n12 B 0.012426f
C192 VTAIL.t1 B 0.034289f
C193 VTAIL.n13 B 0.076778f
C194 VTAIL.n14 B 0.505126f
C195 VTAIL.n15 B 0.0089f
C196 VTAIL.n16 B 0.009423f
C197 VTAIL.n17 B 0.021035f
C198 VTAIL.n18 B 0.021035f
C199 VTAIL.n19 B 0.009423f
C200 VTAIL.n20 B 0.0089f
C201 VTAIL.n21 B 0.016562f
C202 VTAIL.n22 B 0.016562f
C203 VTAIL.n23 B 0.0089f
C204 VTAIL.n24 B 0.009423f
C205 VTAIL.n25 B 0.021035f
C206 VTAIL.n26 B 0.021035f
C207 VTAIL.n27 B 0.009423f
C208 VTAIL.n28 B 0.0089f
C209 VTAIL.n29 B 0.016562f
C210 VTAIL.n30 B 0.016562f
C211 VTAIL.n31 B 0.0089f
C212 VTAIL.n32 B 0.009423f
C213 VTAIL.n33 B 0.021035f
C214 VTAIL.n34 B 0.047514f
C215 VTAIL.n35 B 0.009423f
C216 VTAIL.n36 B 0.0089f
C217 VTAIL.n37 B 0.038734f
C218 VTAIL.n38 B 0.026803f
C219 VTAIL.n39 B 0.742092f
C220 VTAIL.n40 B 0.024396f
C221 VTAIL.n41 B 0.016562f
C222 VTAIL.n42 B 0.0089f
C223 VTAIL.n43 B 0.021035f
C224 VTAIL.n44 B 0.009423f
C225 VTAIL.n45 B 0.016562f
C226 VTAIL.n46 B 0.0089f
C227 VTAIL.n47 B 0.021035f
C228 VTAIL.n48 B 0.009423f
C229 VTAIL.n49 B 0.016562f
C230 VTAIL.n50 B 0.0089f
C231 VTAIL.n51 B 0.015777f
C232 VTAIL.n52 B 0.012426f
C233 VTAIL.t3 B 0.034289f
C234 VTAIL.n53 B 0.076778f
C235 VTAIL.n54 B 0.505126f
C236 VTAIL.n55 B 0.0089f
C237 VTAIL.n56 B 0.009423f
C238 VTAIL.n57 B 0.021035f
C239 VTAIL.n58 B 0.021035f
C240 VTAIL.n59 B 0.009423f
C241 VTAIL.n60 B 0.0089f
C242 VTAIL.n61 B 0.016562f
C243 VTAIL.n62 B 0.016562f
C244 VTAIL.n63 B 0.0089f
C245 VTAIL.n64 B 0.009423f
C246 VTAIL.n65 B 0.021035f
C247 VTAIL.n66 B 0.021035f
C248 VTAIL.n67 B 0.009423f
C249 VTAIL.n68 B 0.0089f
C250 VTAIL.n69 B 0.016562f
C251 VTAIL.n70 B 0.016562f
C252 VTAIL.n71 B 0.0089f
C253 VTAIL.n72 B 0.009423f
C254 VTAIL.n73 B 0.021035f
C255 VTAIL.n74 B 0.047514f
C256 VTAIL.n75 B 0.009423f
C257 VTAIL.n76 B 0.0089f
C258 VTAIL.n77 B 0.038734f
C259 VTAIL.n78 B 0.026803f
C260 VTAIL.n79 B 0.753479f
C261 VTAIL.n80 B 0.024396f
C262 VTAIL.n81 B 0.016562f
C263 VTAIL.n82 B 0.0089f
C264 VTAIL.n83 B 0.021035f
C265 VTAIL.n84 B 0.009423f
C266 VTAIL.n85 B 0.016562f
C267 VTAIL.n86 B 0.0089f
C268 VTAIL.n87 B 0.021035f
C269 VTAIL.n88 B 0.009423f
C270 VTAIL.n89 B 0.016562f
C271 VTAIL.n90 B 0.0089f
C272 VTAIL.n91 B 0.015777f
C273 VTAIL.n92 B 0.012426f
C274 VTAIL.t0 B 0.034289f
C275 VTAIL.n93 B 0.076778f
C276 VTAIL.n94 B 0.505126f
C277 VTAIL.n95 B 0.0089f
C278 VTAIL.n96 B 0.009423f
C279 VTAIL.n97 B 0.021035f
C280 VTAIL.n98 B 0.021035f
C281 VTAIL.n99 B 0.009423f
C282 VTAIL.n100 B 0.0089f
C283 VTAIL.n101 B 0.016562f
C284 VTAIL.n102 B 0.016562f
C285 VTAIL.n103 B 0.0089f
C286 VTAIL.n104 B 0.009423f
C287 VTAIL.n105 B 0.021035f
C288 VTAIL.n106 B 0.021035f
C289 VTAIL.n107 B 0.009423f
C290 VTAIL.n108 B 0.0089f
C291 VTAIL.n109 B 0.016562f
C292 VTAIL.n110 B 0.016562f
C293 VTAIL.n111 B 0.0089f
C294 VTAIL.n112 B 0.009423f
C295 VTAIL.n113 B 0.021035f
C296 VTAIL.n114 B 0.047514f
C297 VTAIL.n115 B 0.009423f
C298 VTAIL.n116 B 0.0089f
C299 VTAIL.n117 B 0.038734f
C300 VTAIL.n118 B 0.026803f
C301 VTAIL.n119 B 0.695512f
C302 VTAIL.n120 B 0.024396f
C303 VTAIL.n121 B 0.016562f
C304 VTAIL.n122 B 0.0089f
C305 VTAIL.n123 B 0.021035f
C306 VTAIL.n124 B 0.009423f
C307 VTAIL.n125 B 0.016562f
C308 VTAIL.n126 B 0.0089f
C309 VTAIL.n127 B 0.021035f
C310 VTAIL.n128 B 0.009423f
C311 VTAIL.n129 B 0.016562f
C312 VTAIL.n130 B 0.0089f
C313 VTAIL.n131 B 0.015777f
C314 VTAIL.n132 B 0.012426f
C315 VTAIL.t2 B 0.034289f
C316 VTAIL.n133 B 0.076778f
C317 VTAIL.n134 B 0.505126f
C318 VTAIL.n135 B 0.0089f
C319 VTAIL.n136 B 0.009423f
C320 VTAIL.n137 B 0.021035f
C321 VTAIL.n138 B 0.021035f
C322 VTAIL.n139 B 0.009423f
C323 VTAIL.n140 B 0.0089f
C324 VTAIL.n141 B 0.016562f
C325 VTAIL.n142 B 0.016562f
C326 VTAIL.n143 B 0.0089f
C327 VTAIL.n144 B 0.009423f
C328 VTAIL.n145 B 0.021035f
C329 VTAIL.n146 B 0.021035f
C330 VTAIL.n147 B 0.009423f
C331 VTAIL.n148 B 0.0089f
C332 VTAIL.n149 B 0.016562f
C333 VTAIL.n150 B 0.016562f
C334 VTAIL.n151 B 0.0089f
C335 VTAIL.n152 B 0.009423f
C336 VTAIL.n153 B 0.021035f
C337 VTAIL.n154 B 0.047514f
C338 VTAIL.n155 B 0.009423f
C339 VTAIL.n156 B 0.0089f
C340 VTAIL.n157 B 0.038734f
C341 VTAIL.n158 B 0.026803f
C342 VTAIL.n159 B 0.652843f
C343 VN.t1 B 0.710418f
C344 VN.t0 B 0.810914f
.ends

