* NGSPICE file created from diff_pair_sample_1019.ext - technology: sky130A

.subckt diff_pair_sample_1019 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=1.67
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=1.67
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=7.3398 ps=38.42 w=18.82 l=1.67
X3 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=7.3398 ps=38.42 w=18.82 l=1.67
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=7.3398 ps=38.42 w=18.82 l=1.67
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=7.3398 ps=38.42 w=18.82 l=1.67
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=1.67
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=1.67
R0 B.n838 B.n837 585
R1 B.n839 B.n838 585
R2 B.n374 B.n107 585
R3 B.n373 B.n372 585
R4 B.n371 B.n370 585
R5 B.n369 B.n368 585
R6 B.n367 B.n366 585
R7 B.n365 B.n364 585
R8 B.n363 B.n362 585
R9 B.n361 B.n360 585
R10 B.n359 B.n358 585
R11 B.n357 B.n356 585
R12 B.n355 B.n354 585
R13 B.n353 B.n352 585
R14 B.n351 B.n350 585
R15 B.n349 B.n348 585
R16 B.n347 B.n346 585
R17 B.n345 B.n344 585
R18 B.n343 B.n342 585
R19 B.n341 B.n340 585
R20 B.n339 B.n338 585
R21 B.n337 B.n336 585
R22 B.n335 B.n334 585
R23 B.n333 B.n332 585
R24 B.n331 B.n330 585
R25 B.n329 B.n328 585
R26 B.n327 B.n326 585
R27 B.n325 B.n324 585
R28 B.n323 B.n322 585
R29 B.n321 B.n320 585
R30 B.n319 B.n318 585
R31 B.n317 B.n316 585
R32 B.n315 B.n314 585
R33 B.n313 B.n312 585
R34 B.n311 B.n310 585
R35 B.n309 B.n308 585
R36 B.n307 B.n306 585
R37 B.n305 B.n304 585
R38 B.n303 B.n302 585
R39 B.n301 B.n300 585
R40 B.n299 B.n298 585
R41 B.n297 B.n296 585
R42 B.n295 B.n294 585
R43 B.n293 B.n292 585
R44 B.n291 B.n290 585
R45 B.n289 B.n288 585
R46 B.n287 B.n286 585
R47 B.n285 B.n284 585
R48 B.n283 B.n282 585
R49 B.n281 B.n280 585
R50 B.n279 B.n278 585
R51 B.n277 B.n276 585
R52 B.n275 B.n274 585
R53 B.n273 B.n272 585
R54 B.n271 B.n270 585
R55 B.n269 B.n268 585
R56 B.n267 B.n266 585
R57 B.n265 B.n264 585
R58 B.n263 B.n262 585
R59 B.n261 B.n260 585
R60 B.n259 B.n258 585
R61 B.n257 B.n256 585
R62 B.n255 B.n254 585
R63 B.n252 B.n251 585
R64 B.n250 B.n249 585
R65 B.n248 B.n247 585
R66 B.n246 B.n245 585
R67 B.n244 B.n243 585
R68 B.n242 B.n241 585
R69 B.n240 B.n239 585
R70 B.n238 B.n237 585
R71 B.n236 B.n235 585
R72 B.n234 B.n233 585
R73 B.n232 B.n231 585
R74 B.n230 B.n229 585
R75 B.n228 B.n227 585
R76 B.n226 B.n225 585
R77 B.n224 B.n223 585
R78 B.n222 B.n221 585
R79 B.n220 B.n219 585
R80 B.n218 B.n217 585
R81 B.n216 B.n215 585
R82 B.n214 B.n213 585
R83 B.n212 B.n211 585
R84 B.n210 B.n209 585
R85 B.n208 B.n207 585
R86 B.n206 B.n205 585
R87 B.n204 B.n203 585
R88 B.n202 B.n201 585
R89 B.n200 B.n199 585
R90 B.n198 B.n197 585
R91 B.n196 B.n195 585
R92 B.n194 B.n193 585
R93 B.n192 B.n191 585
R94 B.n190 B.n189 585
R95 B.n188 B.n187 585
R96 B.n186 B.n185 585
R97 B.n184 B.n183 585
R98 B.n182 B.n181 585
R99 B.n180 B.n179 585
R100 B.n178 B.n177 585
R101 B.n176 B.n175 585
R102 B.n174 B.n173 585
R103 B.n172 B.n171 585
R104 B.n170 B.n169 585
R105 B.n168 B.n167 585
R106 B.n166 B.n165 585
R107 B.n164 B.n163 585
R108 B.n162 B.n161 585
R109 B.n160 B.n159 585
R110 B.n158 B.n157 585
R111 B.n156 B.n155 585
R112 B.n154 B.n153 585
R113 B.n152 B.n151 585
R114 B.n150 B.n149 585
R115 B.n148 B.n147 585
R116 B.n146 B.n145 585
R117 B.n144 B.n143 585
R118 B.n142 B.n141 585
R119 B.n140 B.n139 585
R120 B.n138 B.n137 585
R121 B.n136 B.n135 585
R122 B.n134 B.n133 585
R123 B.n132 B.n131 585
R124 B.n130 B.n129 585
R125 B.n128 B.n127 585
R126 B.n126 B.n125 585
R127 B.n124 B.n123 585
R128 B.n122 B.n121 585
R129 B.n120 B.n119 585
R130 B.n118 B.n117 585
R131 B.n116 B.n115 585
R132 B.n114 B.n113 585
R133 B.n39 B.n38 585
R134 B.n836 B.n40 585
R135 B.n840 B.n40 585
R136 B.n835 B.n834 585
R137 B.n834 B.n36 585
R138 B.n833 B.n35 585
R139 B.n846 B.n35 585
R140 B.n832 B.n34 585
R141 B.n847 B.n34 585
R142 B.n831 B.n33 585
R143 B.n848 B.n33 585
R144 B.n830 B.n829 585
R145 B.n829 B.n29 585
R146 B.n828 B.n28 585
R147 B.n854 B.n28 585
R148 B.n827 B.n27 585
R149 B.n855 B.n27 585
R150 B.n826 B.n26 585
R151 B.n856 B.n26 585
R152 B.n825 B.n824 585
R153 B.n824 B.n22 585
R154 B.n823 B.n21 585
R155 B.n862 B.n21 585
R156 B.n822 B.n20 585
R157 B.n863 B.n20 585
R158 B.n821 B.n19 585
R159 B.n864 B.n19 585
R160 B.n820 B.n819 585
R161 B.n819 B.n15 585
R162 B.n818 B.n14 585
R163 B.n870 B.n14 585
R164 B.n817 B.n13 585
R165 B.n871 B.n13 585
R166 B.n816 B.n12 585
R167 B.n872 B.n12 585
R168 B.n815 B.n814 585
R169 B.n814 B.n8 585
R170 B.n813 B.n7 585
R171 B.n878 B.n7 585
R172 B.n812 B.n6 585
R173 B.n879 B.n6 585
R174 B.n811 B.n5 585
R175 B.n880 B.n5 585
R176 B.n810 B.n809 585
R177 B.n809 B.n4 585
R178 B.n808 B.n375 585
R179 B.n808 B.n807 585
R180 B.n798 B.n376 585
R181 B.n377 B.n376 585
R182 B.n800 B.n799 585
R183 B.n801 B.n800 585
R184 B.n797 B.n381 585
R185 B.n385 B.n381 585
R186 B.n796 B.n795 585
R187 B.n795 B.n794 585
R188 B.n383 B.n382 585
R189 B.n384 B.n383 585
R190 B.n787 B.n786 585
R191 B.n788 B.n787 585
R192 B.n785 B.n390 585
R193 B.n390 B.n389 585
R194 B.n784 B.n783 585
R195 B.n783 B.n782 585
R196 B.n392 B.n391 585
R197 B.n393 B.n392 585
R198 B.n775 B.n774 585
R199 B.n776 B.n775 585
R200 B.n773 B.n398 585
R201 B.n398 B.n397 585
R202 B.n772 B.n771 585
R203 B.n771 B.n770 585
R204 B.n400 B.n399 585
R205 B.n401 B.n400 585
R206 B.n763 B.n762 585
R207 B.n764 B.n763 585
R208 B.n761 B.n406 585
R209 B.n406 B.n405 585
R210 B.n760 B.n759 585
R211 B.n759 B.n758 585
R212 B.n408 B.n407 585
R213 B.n409 B.n408 585
R214 B.n751 B.n750 585
R215 B.n752 B.n751 585
R216 B.n412 B.n411 585
R217 B.n485 B.n483 585
R218 B.n486 B.n482 585
R219 B.n486 B.n413 585
R220 B.n489 B.n488 585
R221 B.n490 B.n481 585
R222 B.n492 B.n491 585
R223 B.n494 B.n480 585
R224 B.n497 B.n496 585
R225 B.n498 B.n479 585
R226 B.n500 B.n499 585
R227 B.n502 B.n478 585
R228 B.n505 B.n504 585
R229 B.n506 B.n477 585
R230 B.n508 B.n507 585
R231 B.n510 B.n476 585
R232 B.n513 B.n512 585
R233 B.n514 B.n475 585
R234 B.n516 B.n515 585
R235 B.n518 B.n474 585
R236 B.n521 B.n520 585
R237 B.n522 B.n473 585
R238 B.n524 B.n523 585
R239 B.n526 B.n472 585
R240 B.n529 B.n528 585
R241 B.n530 B.n471 585
R242 B.n532 B.n531 585
R243 B.n534 B.n470 585
R244 B.n537 B.n536 585
R245 B.n538 B.n469 585
R246 B.n540 B.n539 585
R247 B.n542 B.n468 585
R248 B.n545 B.n544 585
R249 B.n546 B.n467 585
R250 B.n548 B.n547 585
R251 B.n550 B.n466 585
R252 B.n553 B.n552 585
R253 B.n554 B.n465 585
R254 B.n556 B.n555 585
R255 B.n558 B.n464 585
R256 B.n561 B.n560 585
R257 B.n562 B.n463 585
R258 B.n564 B.n563 585
R259 B.n566 B.n462 585
R260 B.n569 B.n568 585
R261 B.n570 B.n461 585
R262 B.n572 B.n571 585
R263 B.n574 B.n460 585
R264 B.n577 B.n576 585
R265 B.n578 B.n459 585
R266 B.n580 B.n579 585
R267 B.n582 B.n458 585
R268 B.n585 B.n584 585
R269 B.n586 B.n457 585
R270 B.n588 B.n587 585
R271 B.n590 B.n456 585
R272 B.n593 B.n592 585
R273 B.n594 B.n455 585
R274 B.n596 B.n595 585
R275 B.n598 B.n454 585
R276 B.n601 B.n600 585
R277 B.n602 B.n453 585
R278 B.n607 B.n606 585
R279 B.n609 B.n452 585
R280 B.n612 B.n611 585
R281 B.n613 B.n451 585
R282 B.n615 B.n614 585
R283 B.n617 B.n450 585
R284 B.n620 B.n619 585
R285 B.n621 B.n449 585
R286 B.n623 B.n622 585
R287 B.n625 B.n448 585
R288 B.n628 B.n627 585
R289 B.n629 B.n444 585
R290 B.n631 B.n630 585
R291 B.n633 B.n443 585
R292 B.n636 B.n635 585
R293 B.n637 B.n442 585
R294 B.n639 B.n638 585
R295 B.n641 B.n441 585
R296 B.n644 B.n643 585
R297 B.n645 B.n440 585
R298 B.n647 B.n646 585
R299 B.n649 B.n439 585
R300 B.n652 B.n651 585
R301 B.n653 B.n438 585
R302 B.n655 B.n654 585
R303 B.n657 B.n437 585
R304 B.n660 B.n659 585
R305 B.n661 B.n436 585
R306 B.n663 B.n662 585
R307 B.n665 B.n435 585
R308 B.n668 B.n667 585
R309 B.n669 B.n434 585
R310 B.n671 B.n670 585
R311 B.n673 B.n433 585
R312 B.n676 B.n675 585
R313 B.n677 B.n432 585
R314 B.n679 B.n678 585
R315 B.n681 B.n431 585
R316 B.n684 B.n683 585
R317 B.n685 B.n430 585
R318 B.n687 B.n686 585
R319 B.n689 B.n429 585
R320 B.n692 B.n691 585
R321 B.n693 B.n428 585
R322 B.n695 B.n694 585
R323 B.n697 B.n427 585
R324 B.n700 B.n699 585
R325 B.n701 B.n426 585
R326 B.n703 B.n702 585
R327 B.n705 B.n425 585
R328 B.n708 B.n707 585
R329 B.n709 B.n424 585
R330 B.n711 B.n710 585
R331 B.n713 B.n423 585
R332 B.n716 B.n715 585
R333 B.n717 B.n422 585
R334 B.n719 B.n718 585
R335 B.n721 B.n421 585
R336 B.n724 B.n723 585
R337 B.n725 B.n420 585
R338 B.n727 B.n726 585
R339 B.n729 B.n419 585
R340 B.n732 B.n731 585
R341 B.n733 B.n418 585
R342 B.n735 B.n734 585
R343 B.n737 B.n417 585
R344 B.n740 B.n739 585
R345 B.n741 B.n416 585
R346 B.n743 B.n742 585
R347 B.n745 B.n415 585
R348 B.n748 B.n747 585
R349 B.n749 B.n414 585
R350 B.n754 B.n753 585
R351 B.n753 B.n752 585
R352 B.n755 B.n410 585
R353 B.n410 B.n409 585
R354 B.n757 B.n756 585
R355 B.n758 B.n757 585
R356 B.n404 B.n403 585
R357 B.n405 B.n404 585
R358 B.n766 B.n765 585
R359 B.n765 B.n764 585
R360 B.n767 B.n402 585
R361 B.n402 B.n401 585
R362 B.n769 B.n768 585
R363 B.n770 B.n769 585
R364 B.n396 B.n395 585
R365 B.n397 B.n396 585
R366 B.n778 B.n777 585
R367 B.n777 B.n776 585
R368 B.n779 B.n394 585
R369 B.n394 B.n393 585
R370 B.n781 B.n780 585
R371 B.n782 B.n781 585
R372 B.n388 B.n387 585
R373 B.n389 B.n388 585
R374 B.n790 B.n789 585
R375 B.n789 B.n788 585
R376 B.n791 B.n386 585
R377 B.n386 B.n384 585
R378 B.n793 B.n792 585
R379 B.n794 B.n793 585
R380 B.n380 B.n379 585
R381 B.n385 B.n380 585
R382 B.n803 B.n802 585
R383 B.n802 B.n801 585
R384 B.n804 B.n378 585
R385 B.n378 B.n377 585
R386 B.n806 B.n805 585
R387 B.n807 B.n806 585
R388 B.n2 B.n0 585
R389 B.n4 B.n2 585
R390 B.n3 B.n1 585
R391 B.n879 B.n3 585
R392 B.n877 B.n876 585
R393 B.n878 B.n877 585
R394 B.n875 B.n9 585
R395 B.n9 B.n8 585
R396 B.n874 B.n873 585
R397 B.n873 B.n872 585
R398 B.n11 B.n10 585
R399 B.n871 B.n11 585
R400 B.n869 B.n868 585
R401 B.n870 B.n869 585
R402 B.n867 B.n16 585
R403 B.n16 B.n15 585
R404 B.n866 B.n865 585
R405 B.n865 B.n864 585
R406 B.n18 B.n17 585
R407 B.n863 B.n18 585
R408 B.n861 B.n860 585
R409 B.n862 B.n861 585
R410 B.n859 B.n23 585
R411 B.n23 B.n22 585
R412 B.n858 B.n857 585
R413 B.n857 B.n856 585
R414 B.n25 B.n24 585
R415 B.n855 B.n25 585
R416 B.n853 B.n852 585
R417 B.n854 B.n853 585
R418 B.n851 B.n30 585
R419 B.n30 B.n29 585
R420 B.n850 B.n849 585
R421 B.n849 B.n848 585
R422 B.n32 B.n31 585
R423 B.n847 B.n32 585
R424 B.n845 B.n844 585
R425 B.n846 B.n845 585
R426 B.n843 B.n37 585
R427 B.n37 B.n36 585
R428 B.n842 B.n841 585
R429 B.n841 B.n840 585
R430 B.n882 B.n881 585
R431 B.n881 B.n880 585
R432 B.n445 B.t13 477.615
R433 B.n603 B.t2 477.615
R434 B.n110 B.t6 477.615
R435 B.n108 B.t10 477.615
R436 B.n753 B.n412 473.281
R437 B.n841 B.n39 473.281
R438 B.n751 B.n414 473.281
R439 B.n838 B.n40 473.281
R440 B.n445 B.t15 438.308
R441 B.n108 B.t11 438.308
R442 B.n603 B.t5 438.308
R443 B.n110 B.t8 438.308
R444 B.n446 B.t14 399.521
R445 B.n109 B.t12 399.521
R446 B.n604 B.t4 399.521
R447 B.n111 B.t9 399.521
R448 B.n839 B.n106 256.663
R449 B.n839 B.n105 256.663
R450 B.n839 B.n104 256.663
R451 B.n839 B.n103 256.663
R452 B.n839 B.n102 256.663
R453 B.n839 B.n101 256.663
R454 B.n839 B.n100 256.663
R455 B.n839 B.n99 256.663
R456 B.n839 B.n98 256.663
R457 B.n839 B.n97 256.663
R458 B.n839 B.n96 256.663
R459 B.n839 B.n95 256.663
R460 B.n839 B.n94 256.663
R461 B.n839 B.n93 256.663
R462 B.n839 B.n92 256.663
R463 B.n839 B.n91 256.663
R464 B.n839 B.n90 256.663
R465 B.n839 B.n89 256.663
R466 B.n839 B.n88 256.663
R467 B.n839 B.n87 256.663
R468 B.n839 B.n86 256.663
R469 B.n839 B.n85 256.663
R470 B.n839 B.n84 256.663
R471 B.n839 B.n83 256.663
R472 B.n839 B.n82 256.663
R473 B.n839 B.n81 256.663
R474 B.n839 B.n80 256.663
R475 B.n839 B.n79 256.663
R476 B.n839 B.n78 256.663
R477 B.n839 B.n77 256.663
R478 B.n839 B.n76 256.663
R479 B.n839 B.n75 256.663
R480 B.n839 B.n74 256.663
R481 B.n839 B.n73 256.663
R482 B.n839 B.n72 256.663
R483 B.n839 B.n71 256.663
R484 B.n839 B.n70 256.663
R485 B.n839 B.n69 256.663
R486 B.n839 B.n68 256.663
R487 B.n839 B.n67 256.663
R488 B.n839 B.n66 256.663
R489 B.n839 B.n65 256.663
R490 B.n839 B.n64 256.663
R491 B.n839 B.n63 256.663
R492 B.n839 B.n62 256.663
R493 B.n839 B.n61 256.663
R494 B.n839 B.n60 256.663
R495 B.n839 B.n59 256.663
R496 B.n839 B.n58 256.663
R497 B.n839 B.n57 256.663
R498 B.n839 B.n56 256.663
R499 B.n839 B.n55 256.663
R500 B.n839 B.n54 256.663
R501 B.n839 B.n53 256.663
R502 B.n839 B.n52 256.663
R503 B.n839 B.n51 256.663
R504 B.n839 B.n50 256.663
R505 B.n839 B.n49 256.663
R506 B.n839 B.n48 256.663
R507 B.n839 B.n47 256.663
R508 B.n839 B.n46 256.663
R509 B.n839 B.n45 256.663
R510 B.n839 B.n44 256.663
R511 B.n839 B.n43 256.663
R512 B.n839 B.n42 256.663
R513 B.n839 B.n41 256.663
R514 B.n484 B.n413 256.663
R515 B.n487 B.n413 256.663
R516 B.n493 B.n413 256.663
R517 B.n495 B.n413 256.663
R518 B.n501 B.n413 256.663
R519 B.n503 B.n413 256.663
R520 B.n509 B.n413 256.663
R521 B.n511 B.n413 256.663
R522 B.n517 B.n413 256.663
R523 B.n519 B.n413 256.663
R524 B.n525 B.n413 256.663
R525 B.n527 B.n413 256.663
R526 B.n533 B.n413 256.663
R527 B.n535 B.n413 256.663
R528 B.n541 B.n413 256.663
R529 B.n543 B.n413 256.663
R530 B.n549 B.n413 256.663
R531 B.n551 B.n413 256.663
R532 B.n557 B.n413 256.663
R533 B.n559 B.n413 256.663
R534 B.n565 B.n413 256.663
R535 B.n567 B.n413 256.663
R536 B.n573 B.n413 256.663
R537 B.n575 B.n413 256.663
R538 B.n581 B.n413 256.663
R539 B.n583 B.n413 256.663
R540 B.n589 B.n413 256.663
R541 B.n591 B.n413 256.663
R542 B.n597 B.n413 256.663
R543 B.n599 B.n413 256.663
R544 B.n608 B.n413 256.663
R545 B.n610 B.n413 256.663
R546 B.n616 B.n413 256.663
R547 B.n618 B.n413 256.663
R548 B.n624 B.n413 256.663
R549 B.n626 B.n413 256.663
R550 B.n632 B.n413 256.663
R551 B.n634 B.n413 256.663
R552 B.n640 B.n413 256.663
R553 B.n642 B.n413 256.663
R554 B.n648 B.n413 256.663
R555 B.n650 B.n413 256.663
R556 B.n656 B.n413 256.663
R557 B.n658 B.n413 256.663
R558 B.n664 B.n413 256.663
R559 B.n666 B.n413 256.663
R560 B.n672 B.n413 256.663
R561 B.n674 B.n413 256.663
R562 B.n680 B.n413 256.663
R563 B.n682 B.n413 256.663
R564 B.n688 B.n413 256.663
R565 B.n690 B.n413 256.663
R566 B.n696 B.n413 256.663
R567 B.n698 B.n413 256.663
R568 B.n704 B.n413 256.663
R569 B.n706 B.n413 256.663
R570 B.n712 B.n413 256.663
R571 B.n714 B.n413 256.663
R572 B.n720 B.n413 256.663
R573 B.n722 B.n413 256.663
R574 B.n728 B.n413 256.663
R575 B.n730 B.n413 256.663
R576 B.n736 B.n413 256.663
R577 B.n738 B.n413 256.663
R578 B.n744 B.n413 256.663
R579 B.n746 B.n413 256.663
R580 B.n753 B.n410 163.367
R581 B.n757 B.n410 163.367
R582 B.n757 B.n404 163.367
R583 B.n765 B.n404 163.367
R584 B.n765 B.n402 163.367
R585 B.n769 B.n402 163.367
R586 B.n769 B.n396 163.367
R587 B.n777 B.n396 163.367
R588 B.n777 B.n394 163.367
R589 B.n781 B.n394 163.367
R590 B.n781 B.n388 163.367
R591 B.n789 B.n388 163.367
R592 B.n789 B.n386 163.367
R593 B.n793 B.n386 163.367
R594 B.n793 B.n380 163.367
R595 B.n802 B.n380 163.367
R596 B.n802 B.n378 163.367
R597 B.n806 B.n378 163.367
R598 B.n806 B.n2 163.367
R599 B.n881 B.n2 163.367
R600 B.n881 B.n3 163.367
R601 B.n877 B.n3 163.367
R602 B.n877 B.n9 163.367
R603 B.n873 B.n9 163.367
R604 B.n873 B.n11 163.367
R605 B.n869 B.n11 163.367
R606 B.n869 B.n16 163.367
R607 B.n865 B.n16 163.367
R608 B.n865 B.n18 163.367
R609 B.n861 B.n18 163.367
R610 B.n861 B.n23 163.367
R611 B.n857 B.n23 163.367
R612 B.n857 B.n25 163.367
R613 B.n853 B.n25 163.367
R614 B.n853 B.n30 163.367
R615 B.n849 B.n30 163.367
R616 B.n849 B.n32 163.367
R617 B.n845 B.n32 163.367
R618 B.n845 B.n37 163.367
R619 B.n841 B.n37 163.367
R620 B.n486 B.n485 163.367
R621 B.n488 B.n486 163.367
R622 B.n492 B.n481 163.367
R623 B.n496 B.n494 163.367
R624 B.n500 B.n479 163.367
R625 B.n504 B.n502 163.367
R626 B.n508 B.n477 163.367
R627 B.n512 B.n510 163.367
R628 B.n516 B.n475 163.367
R629 B.n520 B.n518 163.367
R630 B.n524 B.n473 163.367
R631 B.n528 B.n526 163.367
R632 B.n532 B.n471 163.367
R633 B.n536 B.n534 163.367
R634 B.n540 B.n469 163.367
R635 B.n544 B.n542 163.367
R636 B.n548 B.n467 163.367
R637 B.n552 B.n550 163.367
R638 B.n556 B.n465 163.367
R639 B.n560 B.n558 163.367
R640 B.n564 B.n463 163.367
R641 B.n568 B.n566 163.367
R642 B.n572 B.n461 163.367
R643 B.n576 B.n574 163.367
R644 B.n580 B.n459 163.367
R645 B.n584 B.n582 163.367
R646 B.n588 B.n457 163.367
R647 B.n592 B.n590 163.367
R648 B.n596 B.n455 163.367
R649 B.n600 B.n598 163.367
R650 B.n607 B.n453 163.367
R651 B.n611 B.n609 163.367
R652 B.n615 B.n451 163.367
R653 B.n619 B.n617 163.367
R654 B.n623 B.n449 163.367
R655 B.n627 B.n625 163.367
R656 B.n631 B.n444 163.367
R657 B.n635 B.n633 163.367
R658 B.n639 B.n442 163.367
R659 B.n643 B.n641 163.367
R660 B.n647 B.n440 163.367
R661 B.n651 B.n649 163.367
R662 B.n655 B.n438 163.367
R663 B.n659 B.n657 163.367
R664 B.n663 B.n436 163.367
R665 B.n667 B.n665 163.367
R666 B.n671 B.n434 163.367
R667 B.n675 B.n673 163.367
R668 B.n679 B.n432 163.367
R669 B.n683 B.n681 163.367
R670 B.n687 B.n430 163.367
R671 B.n691 B.n689 163.367
R672 B.n695 B.n428 163.367
R673 B.n699 B.n697 163.367
R674 B.n703 B.n426 163.367
R675 B.n707 B.n705 163.367
R676 B.n711 B.n424 163.367
R677 B.n715 B.n713 163.367
R678 B.n719 B.n422 163.367
R679 B.n723 B.n721 163.367
R680 B.n727 B.n420 163.367
R681 B.n731 B.n729 163.367
R682 B.n735 B.n418 163.367
R683 B.n739 B.n737 163.367
R684 B.n743 B.n416 163.367
R685 B.n747 B.n745 163.367
R686 B.n751 B.n408 163.367
R687 B.n759 B.n408 163.367
R688 B.n759 B.n406 163.367
R689 B.n763 B.n406 163.367
R690 B.n763 B.n400 163.367
R691 B.n771 B.n400 163.367
R692 B.n771 B.n398 163.367
R693 B.n775 B.n398 163.367
R694 B.n775 B.n392 163.367
R695 B.n783 B.n392 163.367
R696 B.n783 B.n390 163.367
R697 B.n787 B.n390 163.367
R698 B.n787 B.n383 163.367
R699 B.n795 B.n383 163.367
R700 B.n795 B.n381 163.367
R701 B.n800 B.n381 163.367
R702 B.n800 B.n376 163.367
R703 B.n808 B.n376 163.367
R704 B.n809 B.n808 163.367
R705 B.n809 B.n5 163.367
R706 B.n6 B.n5 163.367
R707 B.n7 B.n6 163.367
R708 B.n814 B.n7 163.367
R709 B.n814 B.n12 163.367
R710 B.n13 B.n12 163.367
R711 B.n14 B.n13 163.367
R712 B.n819 B.n14 163.367
R713 B.n819 B.n19 163.367
R714 B.n20 B.n19 163.367
R715 B.n21 B.n20 163.367
R716 B.n824 B.n21 163.367
R717 B.n824 B.n26 163.367
R718 B.n27 B.n26 163.367
R719 B.n28 B.n27 163.367
R720 B.n829 B.n28 163.367
R721 B.n829 B.n33 163.367
R722 B.n34 B.n33 163.367
R723 B.n35 B.n34 163.367
R724 B.n834 B.n35 163.367
R725 B.n834 B.n40 163.367
R726 B.n115 B.n114 163.367
R727 B.n119 B.n118 163.367
R728 B.n123 B.n122 163.367
R729 B.n127 B.n126 163.367
R730 B.n131 B.n130 163.367
R731 B.n135 B.n134 163.367
R732 B.n139 B.n138 163.367
R733 B.n143 B.n142 163.367
R734 B.n147 B.n146 163.367
R735 B.n151 B.n150 163.367
R736 B.n155 B.n154 163.367
R737 B.n159 B.n158 163.367
R738 B.n163 B.n162 163.367
R739 B.n167 B.n166 163.367
R740 B.n171 B.n170 163.367
R741 B.n175 B.n174 163.367
R742 B.n179 B.n178 163.367
R743 B.n183 B.n182 163.367
R744 B.n187 B.n186 163.367
R745 B.n191 B.n190 163.367
R746 B.n195 B.n194 163.367
R747 B.n199 B.n198 163.367
R748 B.n203 B.n202 163.367
R749 B.n207 B.n206 163.367
R750 B.n211 B.n210 163.367
R751 B.n215 B.n214 163.367
R752 B.n219 B.n218 163.367
R753 B.n223 B.n222 163.367
R754 B.n227 B.n226 163.367
R755 B.n231 B.n230 163.367
R756 B.n235 B.n234 163.367
R757 B.n239 B.n238 163.367
R758 B.n243 B.n242 163.367
R759 B.n247 B.n246 163.367
R760 B.n251 B.n250 163.367
R761 B.n256 B.n255 163.367
R762 B.n260 B.n259 163.367
R763 B.n264 B.n263 163.367
R764 B.n268 B.n267 163.367
R765 B.n272 B.n271 163.367
R766 B.n276 B.n275 163.367
R767 B.n280 B.n279 163.367
R768 B.n284 B.n283 163.367
R769 B.n288 B.n287 163.367
R770 B.n292 B.n291 163.367
R771 B.n296 B.n295 163.367
R772 B.n300 B.n299 163.367
R773 B.n304 B.n303 163.367
R774 B.n308 B.n307 163.367
R775 B.n312 B.n311 163.367
R776 B.n316 B.n315 163.367
R777 B.n320 B.n319 163.367
R778 B.n324 B.n323 163.367
R779 B.n328 B.n327 163.367
R780 B.n332 B.n331 163.367
R781 B.n336 B.n335 163.367
R782 B.n340 B.n339 163.367
R783 B.n344 B.n343 163.367
R784 B.n348 B.n347 163.367
R785 B.n352 B.n351 163.367
R786 B.n356 B.n355 163.367
R787 B.n360 B.n359 163.367
R788 B.n364 B.n363 163.367
R789 B.n368 B.n367 163.367
R790 B.n372 B.n371 163.367
R791 B.n838 B.n107 163.367
R792 B.n484 B.n412 71.676
R793 B.n488 B.n487 71.676
R794 B.n493 B.n492 71.676
R795 B.n496 B.n495 71.676
R796 B.n501 B.n500 71.676
R797 B.n504 B.n503 71.676
R798 B.n509 B.n508 71.676
R799 B.n512 B.n511 71.676
R800 B.n517 B.n516 71.676
R801 B.n520 B.n519 71.676
R802 B.n525 B.n524 71.676
R803 B.n528 B.n527 71.676
R804 B.n533 B.n532 71.676
R805 B.n536 B.n535 71.676
R806 B.n541 B.n540 71.676
R807 B.n544 B.n543 71.676
R808 B.n549 B.n548 71.676
R809 B.n552 B.n551 71.676
R810 B.n557 B.n556 71.676
R811 B.n560 B.n559 71.676
R812 B.n565 B.n564 71.676
R813 B.n568 B.n567 71.676
R814 B.n573 B.n572 71.676
R815 B.n576 B.n575 71.676
R816 B.n581 B.n580 71.676
R817 B.n584 B.n583 71.676
R818 B.n589 B.n588 71.676
R819 B.n592 B.n591 71.676
R820 B.n597 B.n596 71.676
R821 B.n600 B.n599 71.676
R822 B.n608 B.n607 71.676
R823 B.n611 B.n610 71.676
R824 B.n616 B.n615 71.676
R825 B.n619 B.n618 71.676
R826 B.n624 B.n623 71.676
R827 B.n627 B.n626 71.676
R828 B.n632 B.n631 71.676
R829 B.n635 B.n634 71.676
R830 B.n640 B.n639 71.676
R831 B.n643 B.n642 71.676
R832 B.n648 B.n647 71.676
R833 B.n651 B.n650 71.676
R834 B.n656 B.n655 71.676
R835 B.n659 B.n658 71.676
R836 B.n664 B.n663 71.676
R837 B.n667 B.n666 71.676
R838 B.n672 B.n671 71.676
R839 B.n675 B.n674 71.676
R840 B.n680 B.n679 71.676
R841 B.n683 B.n682 71.676
R842 B.n688 B.n687 71.676
R843 B.n691 B.n690 71.676
R844 B.n696 B.n695 71.676
R845 B.n699 B.n698 71.676
R846 B.n704 B.n703 71.676
R847 B.n707 B.n706 71.676
R848 B.n712 B.n711 71.676
R849 B.n715 B.n714 71.676
R850 B.n720 B.n719 71.676
R851 B.n723 B.n722 71.676
R852 B.n728 B.n727 71.676
R853 B.n731 B.n730 71.676
R854 B.n736 B.n735 71.676
R855 B.n739 B.n738 71.676
R856 B.n744 B.n743 71.676
R857 B.n747 B.n746 71.676
R858 B.n41 B.n39 71.676
R859 B.n115 B.n42 71.676
R860 B.n119 B.n43 71.676
R861 B.n123 B.n44 71.676
R862 B.n127 B.n45 71.676
R863 B.n131 B.n46 71.676
R864 B.n135 B.n47 71.676
R865 B.n139 B.n48 71.676
R866 B.n143 B.n49 71.676
R867 B.n147 B.n50 71.676
R868 B.n151 B.n51 71.676
R869 B.n155 B.n52 71.676
R870 B.n159 B.n53 71.676
R871 B.n163 B.n54 71.676
R872 B.n167 B.n55 71.676
R873 B.n171 B.n56 71.676
R874 B.n175 B.n57 71.676
R875 B.n179 B.n58 71.676
R876 B.n183 B.n59 71.676
R877 B.n187 B.n60 71.676
R878 B.n191 B.n61 71.676
R879 B.n195 B.n62 71.676
R880 B.n199 B.n63 71.676
R881 B.n203 B.n64 71.676
R882 B.n207 B.n65 71.676
R883 B.n211 B.n66 71.676
R884 B.n215 B.n67 71.676
R885 B.n219 B.n68 71.676
R886 B.n223 B.n69 71.676
R887 B.n227 B.n70 71.676
R888 B.n231 B.n71 71.676
R889 B.n235 B.n72 71.676
R890 B.n239 B.n73 71.676
R891 B.n243 B.n74 71.676
R892 B.n247 B.n75 71.676
R893 B.n251 B.n76 71.676
R894 B.n256 B.n77 71.676
R895 B.n260 B.n78 71.676
R896 B.n264 B.n79 71.676
R897 B.n268 B.n80 71.676
R898 B.n272 B.n81 71.676
R899 B.n276 B.n82 71.676
R900 B.n280 B.n83 71.676
R901 B.n284 B.n84 71.676
R902 B.n288 B.n85 71.676
R903 B.n292 B.n86 71.676
R904 B.n296 B.n87 71.676
R905 B.n300 B.n88 71.676
R906 B.n304 B.n89 71.676
R907 B.n308 B.n90 71.676
R908 B.n312 B.n91 71.676
R909 B.n316 B.n92 71.676
R910 B.n320 B.n93 71.676
R911 B.n324 B.n94 71.676
R912 B.n328 B.n95 71.676
R913 B.n332 B.n96 71.676
R914 B.n336 B.n97 71.676
R915 B.n340 B.n98 71.676
R916 B.n344 B.n99 71.676
R917 B.n348 B.n100 71.676
R918 B.n352 B.n101 71.676
R919 B.n356 B.n102 71.676
R920 B.n360 B.n103 71.676
R921 B.n364 B.n104 71.676
R922 B.n368 B.n105 71.676
R923 B.n372 B.n106 71.676
R924 B.n107 B.n106 71.676
R925 B.n371 B.n105 71.676
R926 B.n367 B.n104 71.676
R927 B.n363 B.n103 71.676
R928 B.n359 B.n102 71.676
R929 B.n355 B.n101 71.676
R930 B.n351 B.n100 71.676
R931 B.n347 B.n99 71.676
R932 B.n343 B.n98 71.676
R933 B.n339 B.n97 71.676
R934 B.n335 B.n96 71.676
R935 B.n331 B.n95 71.676
R936 B.n327 B.n94 71.676
R937 B.n323 B.n93 71.676
R938 B.n319 B.n92 71.676
R939 B.n315 B.n91 71.676
R940 B.n311 B.n90 71.676
R941 B.n307 B.n89 71.676
R942 B.n303 B.n88 71.676
R943 B.n299 B.n87 71.676
R944 B.n295 B.n86 71.676
R945 B.n291 B.n85 71.676
R946 B.n287 B.n84 71.676
R947 B.n283 B.n83 71.676
R948 B.n279 B.n82 71.676
R949 B.n275 B.n81 71.676
R950 B.n271 B.n80 71.676
R951 B.n267 B.n79 71.676
R952 B.n263 B.n78 71.676
R953 B.n259 B.n77 71.676
R954 B.n255 B.n76 71.676
R955 B.n250 B.n75 71.676
R956 B.n246 B.n74 71.676
R957 B.n242 B.n73 71.676
R958 B.n238 B.n72 71.676
R959 B.n234 B.n71 71.676
R960 B.n230 B.n70 71.676
R961 B.n226 B.n69 71.676
R962 B.n222 B.n68 71.676
R963 B.n218 B.n67 71.676
R964 B.n214 B.n66 71.676
R965 B.n210 B.n65 71.676
R966 B.n206 B.n64 71.676
R967 B.n202 B.n63 71.676
R968 B.n198 B.n62 71.676
R969 B.n194 B.n61 71.676
R970 B.n190 B.n60 71.676
R971 B.n186 B.n59 71.676
R972 B.n182 B.n58 71.676
R973 B.n178 B.n57 71.676
R974 B.n174 B.n56 71.676
R975 B.n170 B.n55 71.676
R976 B.n166 B.n54 71.676
R977 B.n162 B.n53 71.676
R978 B.n158 B.n52 71.676
R979 B.n154 B.n51 71.676
R980 B.n150 B.n50 71.676
R981 B.n146 B.n49 71.676
R982 B.n142 B.n48 71.676
R983 B.n138 B.n47 71.676
R984 B.n134 B.n46 71.676
R985 B.n130 B.n45 71.676
R986 B.n126 B.n44 71.676
R987 B.n122 B.n43 71.676
R988 B.n118 B.n42 71.676
R989 B.n114 B.n41 71.676
R990 B.n485 B.n484 71.676
R991 B.n487 B.n481 71.676
R992 B.n494 B.n493 71.676
R993 B.n495 B.n479 71.676
R994 B.n502 B.n501 71.676
R995 B.n503 B.n477 71.676
R996 B.n510 B.n509 71.676
R997 B.n511 B.n475 71.676
R998 B.n518 B.n517 71.676
R999 B.n519 B.n473 71.676
R1000 B.n526 B.n525 71.676
R1001 B.n527 B.n471 71.676
R1002 B.n534 B.n533 71.676
R1003 B.n535 B.n469 71.676
R1004 B.n542 B.n541 71.676
R1005 B.n543 B.n467 71.676
R1006 B.n550 B.n549 71.676
R1007 B.n551 B.n465 71.676
R1008 B.n558 B.n557 71.676
R1009 B.n559 B.n463 71.676
R1010 B.n566 B.n565 71.676
R1011 B.n567 B.n461 71.676
R1012 B.n574 B.n573 71.676
R1013 B.n575 B.n459 71.676
R1014 B.n582 B.n581 71.676
R1015 B.n583 B.n457 71.676
R1016 B.n590 B.n589 71.676
R1017 B.n591 B.n455 71.676
R1018 B.n598 B.n597 71.676
R1019 B.n599 B.n453 71.676
R1020 B.n609 B.n608 71.676
R1021 B.n610 B.n451 71.676
R1022 B.n617 B.n616 71.676
R1023 B.n618 B.n449 71.676
R1024 B.n625 B.n624 71.676
R1025 B.n626 B.n444 71.676
R1026 B.n633 B.n632 71.676
R1027 B.n634 B.n442 71.676
R1028 B.n641 B.n640 71.676
R1029 B.n642 B.n440 71.676
R1030 B.n649 B.n648 71.676
R1031 B.n650 B.n438 71.676
R1032 B.n657 B.n656 71.676
R1033 B.n658 B.n436 71.676
R1034 B.n665 B.n664 71.676
R1035 B.n666 B.n434 71.676
R1036 B.n673 B.n672 71.676
R1037 B.n674 B.n432 71.676
R1038 B.n681 B.n680 71.676
R1039 B.n682 B.n430 71.676
R1040 B.n689 B.n688 71.676
R1041 B.n690 B.n428 71.676
R1042 B.n697 B.n696 71.676
R1043 B.n698 B.n426 71.676
R1044 B.n705 B.n704 71.676
R1045 B.n706 B.n424 71.676
R1046 B.n713 B.n712 71.676
R1047 B.n714 B.n422 71.676
R1048 B.n721 B.n720 71.676
R1049 B.n722 B.n420 71.676
R1050 B.n729 B.n728 71.676
R1051 B.n730 B.n418 71.676
R1052 B.n737 B.n736 71.676
R1053 B.n738 B.n416 71.676
R1054 B.n745 B.n744 71.676
R1055 B.n746 B.n414 71.676
R1056 B.n447 B.n446 59.5399
R1057 B.n605 B.n604 59.5399
R1058 B.n112 B.n111 59.5399
R1059 B.n253 B.n109 59.5399
R1060 B.n752 B.n413 52.501
R1061 B.n840 B.n839 52.501
R1062 B.n446 B.n445 38.7884
R1063 B.n604 B.n603 38.7884
R1064 B.n111 B.n110 38.7884
R1065 B.n109 B.n108 38.7884
R1066 B.n752 B.n409 31.0443
R1067 B.n758 B.n409 31.0443
R1068 B.n758 B.n405 31.0443
R1069 B.n764 B.n405 31.0443
R1070 B.n764 B.n401 31.0443
R1071 B.n770 B.n401 31.0443
R1072 B.n776 B.n397 31.0443
R1073 B.n776 B.n393 31.0443
R1074 B.n782 B.n393 31.0443
R1075 B.n782 B.n389 31.0443
R1076 B.n788 B.n389 31.0443
R1077 B.n788 B.n384 31.0443
R1078 B.n794 B.n384 31.0443
R1079 B.n794 B.n385 31.0443
R1080 B.n801 B.n377 31.0443
R1081 B.n807 B.n377 31.0443
R1082 B.n807 B.n4 31.0443
R1083 B.n880 B.n4 31.0443
R1084 B.n880 B.n879 31.0443
R1085 B.n879 B.n878 31.0443
R1086 B.n878 B.n8 31.0443
R1087 B.n872 B.n8 31.0443
R1088 B.n871 B.n870 31.0443
R1089 B.n870 B.n15 31.0443
R1090 B.n864 B.n15 31.0443
R1091 B.n864 B.n863 31.0443
R1092 B.n863 B.n862 31.0443
R1093 B.n862 B.n22 31.0443
R1094 B.n856 B.n22 31.0443
R1095 B.n856 B.n855 31.0443
R1096 B.n854 B.n29 31.0443
R1097 B.n848 B.n29 31.0443
R1098 B.n848 B.n847 31.0443
R1099 B.n847 B.n846 31.0443
R1100 B.n846 B.n36 31.0443
R1101 B.n840 B.n36 31.0443
R1102 B.n842 B.n38 30.7517
R1103 B.n837 B.n836 30.7517
R1104 B.n750 B.n749 30.7517
R1105 B.n754 B.n411 30.7517
R1106 B.t3 B.n397 19.6311
R1107 B.n855 B.t7 19.6311
R1108 B B.n882 18.0485
R1109 B.n801 B.t1 16.892
R1110 B.n872 B.t0 16.892
R1111 B.n385 B.t1 14.1528
R1112 B.t0 B.n871 14.1528
R1113 B.n770 B.t3 11.4137
R1114 B.t7 B.n854 11.4137
R1115 B.n113 B.n38 10.6151
R1116 B.n116 B.n113 10.6151
R1117 B.n117 B.n116 10.6151
R1118 B.n120 B.n117 10.6151
R1119 B.n121 B.n120 10.6151
R1120 B.n124 B.n121 10.6151
R1121 B.n125 B.n124 10.6151
R1122 B.n128 B.n125 10.6151
R1123 B.n129 B.n128 10.6151
R1124 B.n132 B.n129 10.6151
R1125 B.n133 B.n132 10.6151
R1126 B.n136 B.n133 10.6151
R1127 B.n137 B.n136 10.6151
R1128 B.n140 B.n137 10.6151
R1129 B.n141 B.n140 10.6151
R1130 B.n144 B.n141 10.6151
R1131 B.n145 B.n144 10.6151
R1132 B.n148 B.n145 10.6151
R1133 B.n149 B.n148 10.6151
R1134 B.n152 B.n149 10.6151
R1135 B.n153 B.n152 10.6151
R1136 B.n156 B.n153 10.6151
R1137 B.n157 B.n156 10.6151
R1138 B.n160 B.n157 10.6151
R1139 B.n161 B.n160 10.6151
R1140 B.n164 B.n161 10.6151
R1141 B.n165 B.n164 10.6151
R1142 B.n168 B.n165 10.6151
R1143 B.n169 B.n168 10.6151
R1144 B.n172 B.n169 10.6151
R1145 B.n173 B.n172 10.6151
R1146 B.n176 B.n173 10.6151
R1147 B.n177 B.n176 10.6151
R1148 B.n180 B.n177 10.6151
R1149 B.n181 B.n180 10.6151
R1150 B.n184 B.n181 10.6151
R1151 B.n185 B.n184 10.6151
R1152 B.n188 B.n185 10.6151
R1153 B.n189 B.n188 10.6151
R1154 B.n192 B.n189 10.6151
R1155 B.n193 B.n192 10.6151
R1156 B.n196 B.n193 10.6151
R1157 B.n197 B.n196 10.6151
R1158 B.n200 B.n197 10.6151
R1159 B.n201 B.n200 10.6151
R1160 B.n204 B.n201 10.6151
R1161 B.n205 B.n204 10.6151
R1162 B.n208 B.n205 10.6151
R1163 B.n209 B.n208 10.6151
R1164 B.n212 B.n209 10.6151
R1165 B.n213 B.n212 10.6151
R1166 B.n216 B.n213 10.6151
R1167 B.n217 B.n216 10.6151
R1168 B.n220 B.n217 10.6151
R1169 B.n221 B.n220 10.6151
R1170 B.n224 B.n221 10.6151
R1171 B.n225 B.n224 10.6151
R1172 B.n228 B.n225 10.6151
R1173 B.n229 B.n228 10.6151
R1174 B.n232 B.n229 10.6151
R1175 B.n233 B.n232 10.6151
R1176 B.n237 B.n236 10.6151
R1177 B.n240 B.n237 10.6151
R1178 B.n241 B.n240 10.6151
R1179 B.n244 B.n241 10.6151
R1180 B.n245 B.n244 10.6151
R1181 B.n248 B.n245 10.6151
R1182 B.n249 B.n248 10.6151
R1183 B.n252 B.n249 10.6151
R1184 B.n257 B.n254 10.6151
R1185 B.n258 B.n257 10.6151
R1186 B.n261 B.n258 10.6151
R1187 B.n262 B.n261 10.6151
R1188 B.n265 B.n262 10.6151
R1189 B.n266 B.n265 10.6151
R1190 B.n269 B.n266 10.6151
R1191 B.n270 B.n269 10.6151
R1192 B.n273 B.n270 10.6151
R1193 B.n274 B.n273 10.6151
R1194 B.n277 B.n274 10.6151
R1195 B.n278 B.n277 10.6151
R1196 B.n281 B.n278 10.6151
R1197 B.n282 B.n281 10.6151
R1198 B.n285 B.n282 10.6151
R1199 B.n286 B.n285 10.6151
R1200 B.n289 B.n286 10.6151
R1201 B.n290 B.n289 10.6151
R1202 B.n293 B.n290 10.6151
R1203 B.n294 B.n293 10.6151
R1204 B.n297 B.n294 10.6151
R1205 B.n298 B.n297 10.6151
R1206 B.n301 B.n298 10.6151
R1207 B.n302 B.n301 10.6151
R1208 B.n305 B.n302 10.6151
R1209 B.n306 B.n305 10.6151
R1210 B.n309 B.n306 10.6151
R1211 B.n310 B.n309 10.6151
R1212 B.n313 B.n310 10.6151
R1213 B.n314 B.n313 10.6151
R1214 B.n317 B.n314 10.6151
R1215 B.n318 B.n317 10.6151
R1216 B.n321 B.n318 10.6151
R1217 B.n322 B.n321 10.6151
R1218 B.n325 B.n322 10.6151
R1219 B.n326 B.n325 10.6151
R1220 B.n329 B.n326 10.6151
R1221 B.n330 B.n329 10.6151
R1222 B.n333 B.n330 10.6151
R1223 B.n334 B.n333 10.6151
R1224 B.n337 B.n334 10.6151
R1225 B.n338 B.n337 10.6151
R1226 B.n341 B.n338 10.6151
R1227 B.n342 B.n341 10.6151
R1228 B.n345 B.n342 10.6151
R1229 B.n346 B.n345 10.6151
R1230 B.n349 B.n346 10.6151
R1231 B.n350 B.n349 10.6151
R1232 B.n353 B.n350 10.6151
R1233 B.n354 B.n353 10.6151
R1234 B.n357 B.n354 10.6151
R1235 B.n358 B.n357 10.6151
R1236 B.n361 B.n358 10.6151
R1237 B.n362 B.n361 10.6151
R1238 B.n365 B.n362 10.6151
R1239 B.n366 B.n365 10.6151
R1240 B.n369 B.n366 10.6151
R1241 B.n370 B.n369 10.6151
R1242 B.n373 B.n370 10.6151
R1243 B.n374 B.n373 10.6151
R1244 B.n837 B.n374 10.6151
R1245 B.n750 B.n407 10.6151
R1246 B.n760 B.n407 10.6151
R1247 B.n761 B.n760 10.6151
R1248 B.n762 B.n761 10.6151
R1249 B.n762 B.n399 10.6151
R1250 B.n772 B.n399 10.6151
R1251 B.n773 B.n772 10.6151
R1252 B.n774 B.n773 10.6151
R1253 B.n774 B.n391 10.6151
R1254 B.n784 B.n391 10.6151
R1255 B.n785 B.n784 10.6151
R1256 B.n786 B.n785 10.6151
R1257 B.n786 B.n382 10.6151
R1258 B.n796 B.n382 10.6151
R1259 B.n797 B.n796 10.6151
R1260 B.n799 B.n797 10.6151
R1261 B.n799 B.n798 10.6151
R1262 B.n798 B.n375 10.6151
R1263 B.n810 B.n375 10.6151
R1264 B.n811 B.n810 10.6151
R1265 B.n812 B.n811 10.6151
R1266 B.n813 B.n812 10.6151
R1267 B.n815 B.n813 10.6151
R1268 B.n816 B.n815 10.6151
R1269 B.n817 B.n816 10.6151
R1270 B.n818 B.n817 10.6151
R1271 B.n820 B.n818 10.6151
R1272 B.n821 B.n820 10.6151
R1273 B.n822 B.n821 10.6151
R1274 B.n823 B.n822 10.6151
R1275 B.n825 B.n823 10.6151
R1276 B.n826 B.n825 10.6151
R1277 B.n827 B.n826 10.6151
R1278 B.n828 B.n827 10.6151
R1279 B.n830 B.n828 10.6151
R1280 B.n831 B.n830 10.6151
R1281 B.n832 B.n831 10.6151
R1282 B.n833 B.n832 10.6151
R1283 B.n835 B.n833 10.6151
R1284 B.n836 B.n835 10.6151
R1285 B.n483 B.n411 10.6151
R1286 B.n483 B.n482 10.6151
R1287 B.n489 B.n482 10.6151
R1288 B.n490 B.n489 10.6151
R1289 B.n491 B.n490 10.6151
R1290 B.n491 B.n480 10.6151
R1291 B.n497 B.n480 10.6151
R1292 B.n498 B.n497 10.6151
R1293 B.n499 B.n498 10.6151
R1294 B.n499 B.n478 10.6151
R1295 B.n505 B.n478 10.6151
R1296 B.n506 B.n505 10.6151
R1297 B.n507 B.n506 10.6151
R1298 B.n507 B.n476 10.6151
R1299 B.n513 B.n476 10.6151
R1300 B.n514 B.n513 10.6151
R1301 B.n515 B.n514 10.6151
R1302 B.n515 B.n474 10.6151
R1303 B.n521 B.n474 10.6151
R1304 B.n522 B.n521 10.6151
R1305 B.n523 B.n522 10.6151
R1306 B.n523 B.n472 10.6151
R1307 B.n529 B.n472 10.6151
R1308 B.n530 B.n529 10.6151
R1309 B.n531 B.n530 10.6151
R1310 B.n531 B.n470 10.6151
R1311 B.n537 B.n470 10.6151
R1312 B.n538 B.n537 10.6151
R1313 B.n539 B.n538 10.6151
R1314 B.n539 B.n468 10.6151
R1315 B.n545 B.n468 10.6151
R1316 B.n546 B.n545 10.6151
R1317 B.n547 B.n546 10.6151
R1318 B.n547 B.n466 10.6151
R1319 B.n553 B.n466 10.6151
R1320 B.n554 B.n553 10.6151
R1321 B.n555 B.n554 10.6151
R1322 B.n555 B.n464 10.6151
R1323 B.n561 B.n464 10.6151
R1324 B.n562 B.n561 10.6151
R1325 B.n563 B.n562 10.6151
R1326 B.n563 B.n462 10.6151
R1327 B.n569 B.n462 10.6151
R1328 B.n570 B.n569 10.6151
R1329 B.n571 B.n570 10.6151
R1330 B.n571 B.n460 10.6151
R1331 B.n577 B.n460 10.6151
R1332 B.n578 B.n577 10.6151
R1333 B.n579 B.n578 10.6151
R1334 B.n579 B.n458 10.6151
R1335 B.n585 B.n458 10.6151
R1336 B.n586 B.n585 10.6151
R1337 B.n587 B.n586 10.6151
R1338 B.n587 B.n456 10.6151
R1339 B.n593 B.n456 10.6151
R1340 B.n594 B.n593 10.6151
R1341 B.n595 B.n594 10.6151
R1342 B.n595 B.n454 10.6151
R1343 B.n601 B.n454 10.6151
R1344 B.n602 B.n601 10.6151
R1345 B.n606 B.n602 10.6151
R1346 B.n612 B.n452 10.6151
R1347 B.n613 B.n612 10.6151
R1348 B.n614 B.n613 10.6151
R1349 B.n614 B.n450 10.6151
R1350 B.n620 B.n450 10.6151
R1351 B.n621 B.n620 10.6151
R1352 B.n622 B.n621 10.6151
R1353 B.n622 B.n448 10.6151
R1354 B.n629 B.n628 10.6151
R1355 B.n630 B.n629 10.6151
R1356 B.n630 B.n443 10.6151
R1357 B.n636 B.n443 10.6151
R1358 B.n637 B.n636 10.6151
R1359 B.n638 B.n637 10.6151
R1360 B.n638 B.n441 10.6151
R1361 B.n644 B.n441 10.6151
R1362 B.n645 B.n644 10.6151
R1363 B.n646 B.n645 10.6151
R1364 B.n646 B.n439 10.6151
R1365 B.n652 B.n439 10.6151
R1366 B.n653 B.n652 10.6151
R1367 B.n654 B.n653 10.6151
R1368 B.n654 B.n437 10.6151
R1369 B.n660 B.n437 10.6151
R1370 B.n661 B.n660 10.6151
R1371 B.n662 B.n661 10.6151
R1372 B.n662 B.n435 10.6151
R1373 B.n668 B.n435 10.6151
R1374 B.n669 B.n668 10.6151
R1375 B.n670 B.n669 10.6151
R1376 B.n670 B.n433 10.6151
R1377 B.n676 B.n433 10.6151
R1378 B.n677 B.n676 10.6151
R1379 B.n678 B.n677 10.6151
R1380 B.n678 B.n431 10.6151
R1381 B.n684 B.n431 10.6151
R1382 B.n685 B.n684 10.6151
R1383 B.n686 B.n685 10.6151
R1384 B.n686 B.n429 10.6151
R1385 B.n692 B.n429 10.6151
R1386 B.n693 B.n692 10.6151
R1387 B.n694 B.n693 10.6151
R1388 B.n694 B.n427 10.6151
R1389 B.n700 B.n427 10.6151
R1390 B.n701 B.n700 10.6151
R1391 B.n702 B.n701 10.6151
R1392 B.n702 B.n425 10.6151
R1393 B.n708 B.n425 10.6151
R1394 B.n709 B.n708 10.6151
R1395 B.n710 B.n709 10.6151
R1396 B.n710 B.n423 10.6151
R1397 B.n716 B.n423 10.6151
R1398 B.n717 B.n716 10.6151
R1399 B.n718 B.n717 10.6151
R1400 B.n718 B.n421 10.6151
R1401 B.n724 B.n421 10.6151
R1402 B.n725 B.n724 10.6151
R1403 B.n726 B.n725 10.6151
R1404 B.n726 B.n419 10.6151
R1405 B.n732 B.n419 10.6151
R1406 B.n733 B.n732 10.6151
R1407 B.n734 B.n733 10.6151
R1408 B.n734 B.n417 10.6151
R1409 B.n740 B.n417 10.6151
R1410 B.n741 B.n740 10.6151
R1411 B.n742 B.n741 10.6151
R1412 B.n742 B.n415 10.6151
R1413 B.n748 B.n415 10.6151
R1414 B.n749 B.n748 10.6151
R1415 B.n755 B.n754 10.6151
R1416 B.n756 B.n755 10.6151
R1417 B.n756 B.n403 10.6151
R1418 B.n766 B.n403 10.6151
R1419 B.n767 B.n766 10.6151
R1420 B.n768 B.n767 10.6151
R1421 B.n768 B.n395 10.6151
R1422 B.n778 B.n395 10.6151
R1423 B.n779 B.n778 10.6151
R1424 B.n780 B.n779 10.6151
R1425 B.n780 B.n387 10.6151
R1426 B.n790 B.n387 10.6151
R1427 B.n791 B.n790 10.6151
R1428 B.n792 B.n791 10.6151
R1429 B.n792 B.n379 10.6151
R1430 B.n803 B.n379 10.6151
R1431 B.n804 B.n803 10.6151
R1432 B.n805 B.n804 10.6151
R1433 B.n805 B.n0 10.6151
R1434 B.n876 B.n1 10.6151
R1435 B.n876 B.n875 10.6151
R1436 B.n875 B.n874 10.6151
R1437 B.n874 B.n10 10.6151
R1438 B.n868 B.n10 10.6151
R1439 B.n868 B.n867 10.6151
R1440 B.n867 B.n866 10.6151
R1441 B.n866 B.n17 10.6151
R1442 B.n860 B.n17 10.6151
R1443 B.n860 B.n859 10.6151
R1444 B.n859 B.n858 10.6151
R1445 B.n858 B.n24 10.6151
R1446 B.n852 B.n24 10.6151
R1447 B.n852 B.n851 10.6151
R1448 B.n851 B.n850 10.6151
R1449 B.n850 B.n31 10.6151
R1450 B.n844 B.n31 10.6151
R1451 B.n844 B.n843 10.6151
R1452 B.n843 B.n842 10.6151
R1453 B.n236 B.n112 6.5566
R1454 B.n253 B.n252 6.5566
R1455 B.n605 B.n452 6.5566
R1456 B.n448 B.n447 6.5566
R1457 B.n233 B.n112 4.05904
R1458 B.n254 B.n253 4.05904
R1459 B.n606 B.n605 4.05904
R1460 B.n628 B.n447 4.05904
R1461 B.n882 B.n0 2.81026
R1462 B.n882 B.n1 2.81026
R1463 VP.n0 VP.t1 377.837
R1464 VP.n0 VP.t0 330.481
R1465 VP VP.n0 0.241678
R1466 VTAIL.n414 VTAIL.n413 289.615
R1467 VTAIL.n102 VTAIL.n101 289.615
R1468 VTAIL.n310 VTAIL.n309 289.615
R1469 VTAIL.n206 VTAIL.n205 289.615
R1470 VTAIL.n347 VTAIL.n346 185
R1471 VTAIL.n349 VTAIL.n348 185
R1472 VTAIL.n342 VTAIL.n341 185
R1473 VTAIL.n355 VTAIL.n354 185
R1474 VTAIL.n357 VTAIL.n356 185
R1475 VTAIL.n338 VTAIL.n337 185
R1476 VTAIL.n364 VTAIL.n363 185
R1477 VTAIL.n365 VTAIL.n336 185
R1478 VTAIL.n367 VTAIL.n366 185
R1479 VTAIL.n334 VTAIL.n333 185
R1480 VTAIL.n373 VTAIL.n372 185
R1481 VTAIL.n375 VTAIL.n374 185
R1482 VTAIL.n330 VTAIL.n329 185
R1483 VTAIL.n381 VTAIL.n380 185
R1484 VTAIL.n383 VTAIL.n382 185
R1485 VTAIL.n326 VTAIL.n325 185
R1486 VTAIL.n389 VTAIL.n388 185
R1487 VTAIL.n391 VTAIL.n390 185
R1488 VTAIL.n322 VTAIL.n321 185
R1489 VTAIL.n397 VTAIL.n396 185
R1490 VTAIL.n399 VTAIL.n398 185
R1491 VTAIL.n318 VTAIL.n317 185
R1492 VTAIL.n405 VTAIL.n404 185
R1493 VTAIL.n407 VTAIL.n406 185
R1494 VTAIL.n314 VTAIL.n313 185
R1495 VTAIL.n413 VTAIL.n412 185
R1496 VTAIL.n35 VTAIL.n34 185
R1497 VTAIL.n37 VTAIL.n36 185
R1498 VTAIL.n30 VTAIL.n29 185
R1499 VTAIL.n43 VTAIL.n42 185
R1500 VTAIL.n45 VTAIL.n44 185
R1501 VTAIL.n26 VTAIL.n25 185
R1502 VTAIL.n52 VTAIL.n51 185
R1503 VTAIL.n53 VTAIL.n24 185
R1504 VTAIL.n55 VTAIL.n54 185
R1505 VTAIL.n22 VTAIL.n21 185
R1506 VTAIL.n61 VTAIL.n60 185
R1507 VTAIL.n63 VTAIL.n62 185
R1508 VTAIL.n18 VTAIL.n17 185
R1509 VTAIL.n69 VTAIL.n68 185
R1510 VTAIL.n71 VTAIL.n70 185
R1511 VTAIL.n14 VTAIL.n13 185
R1512 VTAIL.n77 VTAIL.n76 185
R1513 VTAIL.n79 VTAIL.n78 185
R1514 VTAIL.n10 VTAIL.n9 185
R1515 VTAIL.n85 VTAIL.n84 185
R1516 VTAIL.n87 VTAIL.n86 185
R1517 VTAIL.n6 VTAIL.n5 185
R1518 VTAIL.n93 VTAIL.n92 185
R1519 VTAIL.n95 VTAIL.n94 185
R1520 VTAIL.n2 VTAIL.n1 185
R1521 VTAIL.n101 VTAIL.n100 185
R1522 VTAIL.n309 VTAIL.n308 185
R1523 VTAIL.n210 VTAIL.n209 185
R1524 VTAIL.n303 VTAIL.n302 185
R1525 VTAIL.n301 VTAIL.n300 185
R1526 VTAIL.n214 VTAIL.n213 185
R1527 VTAIL.n295 VTAIL.n294 185
R1528 VTAIL.n293 VTAIL.n292 185
R1529 VTAIL.n218 VTAIL.n217 185
R1530 VTAIL.n287 VTAIL.n286 185
R1531 VTAIL.n285 VTAIL.n284 185
R1532 VTAIL.n222 VTAIL.n221 185
R1533 VTAIL.n279 VTAIL.n278 185
R1534 VTAIL.n277 VTAIL.n276 185
R1535 VTAIL.n226 VTAIL.n225 185
R1536 VTAIL.n271 VTAIL.n270 185
R1537 VTAIL.n269 VTAIL.n268 185
R1538 VTAIL.n230 VTAIL.n229 185
R1539 VTAIL.n234 VTAIL.n232 185
R1540 VTAIL.n263 VTAIL.n262 185
R1541 VTAIL.n261 VTAIL.n260 185
R1542 VTAIL.n236 VTAIL.n235 185
R1543 VTAIL.n255 VTAIL.n254 185
R1544 VTAIL.n253 VTAIL.n252 185
R1545 VTAIL.n240 VTAIL.n239 185
R1546 VTAIL.n247 VTAIL.n246 185
R1547 VTAIL.n245 VTAIL.n244 185
R1548 VTAIL.n205 VTAIL.n204 185
R1549 VTAIL.n106 VTAIL.n105 185
R1550 VTAIL.n199 VTAIL.n198 185
R1551 VTAIL.n197 VTAIL.n196 185
R1552 VTAIL.n110 VTAIL.n109 185
R1553 VTAIL.n191 VTAIL.n190 185
R1554 VTAIL.n189 VTAIL.n188 185
R1555 VTAIL.n114 VTAIL.n113 185
R1556 VTAIL.n183 VTAIL.n182 185
R1557 VTAIL.n181 VTAIL.n180 185
R1558 VTAIL.n118 VTAIL.n117 185
R1559 VTAIL.n175 VTAIL.n174 185
R1560 VTAIL.n173 VTAIL.n172 185
R1561 VTAIL.n122 VTAIL.n121 185
R1562 VTAIL.n167 VTAIL.n166 185
R1563 VTAIL.n165 VTAIL.n164 185
R1564 VTAIL.n126 VTAIL.n125 185
R1565 VTAIL.n130 VTAIL.n128 185
R1566 VTAIL.n159 VTAIL.n158 185
R1567 VTAIL.n157 VTAIL.n156 185
R1568 VTAIL.n132 VTAIL.n131 185
R1569 VTAIL.n151 VTAIL.n150 185
R1570 VTAIL.n149 VTAIL.n148 185
R1571 VTAIL.n136 VTAIL.n135 185
R1572 VTAIL.n143 VTAIL.n142 185
R1573 VTAIL.n141 VTAIL.n140 185
R1574 VTAIL.n345 VTAIL.t1 149.524
R1575 VTAIL.n33 VTAIL.t3 149.524
R1576 VTAIL.n243 VTAIL.t2 149.524
R1577 VTAIL.n139 VTAIL.t0 149.524
R1578 VTAIL.n348 VTAIL.n347 104.615
R1579 VTAIL.n348 VTAIL.n341 104.615
R1580 VTAIL.n355 VTAIL.n341 104.615
R1581 VTAIL.n356 VTAIL.n355 104.615
R1582 VTAIL.n356 VTAIL.n337 104.615
R1583 VTAIL.n364 VTAIL.n337 104.615
R1584 VTAIL.n365 VTAIL.n364 104.615
R1585 VTAIL.n366 VTAIL.n365 104.615
R1586 VTAIL.n366 VTAIL.n333 104.615
R1587 VTAIL.n373 VTAIL.n333 104.615
R1588 VTAIL.n374 VTAIL.n373 104.615
R1589 VTAIL.n374 VTAIL.n329 104.615
R1590 VTAIL.n381 VTAIL.n329 104.615
R1591 VTAIL.n382 VTAIL.n381 104.615
R1592 VTAIL.n382 VTAIL.n325 104.615
R1593 VTAIL.n389 VTAIL.n325 104.615
R1594 VTAIL.n390 VTAIL.n389 104.615
R1595 VTAIL.n390 VTAIL.n321 104.615
R1596 VTAIL.n397 VTAIL.n321 104.615
R1597 VTAIL.n398 VTAIL.n397 104.615
R1598 VTAIL.n398 VTAIL.n317 104.615
R1599 VTAIL.n405 VTAIL.n317 104.615
R1600 VTAIL.n406 VTAIL.n405 104.615
R1601 VTAIL.n406 VTAIL.n313 104.615
R1602 VTAIL.n413 VTAIL.n313 104.615
R1603 VTAIL.n36 VTAIL.n35 104.615
R1604 VTAIL.n36 VTAIL.n29 104.615
R1605 VTAIL.n43 VTAIL.n29 104.615
R1606 VTAIL.n44 VTAIL.n43 104.615
R1607 VTAIL.n44 VTAIL.n25 104.615
R1608 VTAIL.n52 VTAIL.n25 104.615
R1609 VTAIL.n53 VTAIL.n52 104.615
R1610 VTAIL.n54 VTAIL.n53 104.615
R1611 VTAIL.n54 VTAIL.n21 104.615
R1612 VTAIL.n61 VTAIL.n21 104.615
R1613 VTAIL.n62 VTAIL.n61 104.615
R1614 VTAIL.n62 VTAIL.n17 104.615
R1615 VTAIL.n69 VTAIL.n17 104.615
R1616 VTAIL.n70 VTAIL.n69 104.615
R1617 VTAIL.n70 VTAIL.n13 104.615
R1618 VTAIL.n77 VTAIL.n13 104.615
R1619 VTAIL.n78 VTAIL.n77 104.615
R1620 VTAIL.n78 VTAIL.n9 104.615
R1621 VTAIL.n85 VTAIL.n9 104.615
R1622 VTAIL.n86 VTAIL.n85 104.615
R1623 VTAIL.n86 VTAIL.n5 104.615
R1624 VTAIL.n93 VTAIL.n5 104.615
R1625 VTAIL.n94 VTAIL.n93 104.615
R1626 VTAIL.n94 VTAIL.n1 104.615
R1627 VTAIL.n101 VTAIL.n1 104.615
R1628 VTAIL.n309 VTAIL.n209 104.615
R1629 VTAIL.n302 VTAIL.n209 104.615
R1630 VTAIL.n302 VTAIL.n301 104.615
R1631 VTAIL.n301 VTAIL.n213 104.615
R1632 VTAIL.n294 VTAIL.n213 104.615
R1633 VTAIL.n294 VTAIL.n293 104.615
R1634 VTAIL.n293 VTAIL.n217 104.615
R1635 VTAIL.n286 VTAIL.n217 104.615
R1636 VTAIL.n286 VTAIL.n285 104.615
R1637 VTAIL.n285 VTAIL.n221 104.615
R1638 VTAIL.n278 VTAIL.n221 104.615
R1639 VTAIL.n278 VTAIL.n277 104.615
R1640 VTAIL.n277 VTAIL.n225 104.615
R1641 VTAIL.n270 VTAIL.n225 104.615
R1642 VTAIL.n270 VTAIL.n269 104.615
R1643 VTAIL.n269 VTAIL.n229 104.615
R1644 VTAIL.n234 VTAIL.n229 104.615
R1645 VTAIL.n262 VTAIL.n234 104.615
R1646 VTAIL.n262 VTAIL.n261 104.615
R1647 VTAIL.n261 VTAIL.n235 104.615
R1648 VTAIL.n254 VTAIL.n235 104.615
R1649 VTAIL.n254 VTAIL.n253 104.615
R1650 VTAIL.n253 VTAIL.n239 104.615
R1651 VTAIL.n246 VTAIL.n239 104.615
R1652 VTAIL.n246 VTAIL.n245 104.615
R1653 VTAIL.n205 VTAIL.n105 104.615
R1654 VTAIL.n198 VTAIL.n105 104.615
R1655 VTAIL.n198 VTAIL.n197 104.615
R1656 VTAIL.n197 VTAIL.n109 104.615
R1657 VTAIL.n190 VTAIL.n109 104.615
R1658 VTAIL.n190 VTAIL.n189 104.615
R1659 VTAIL.n189 VTAIL.n113 104.615
R1660 VTAIL.n182 VTAIL.n113 104.615
R1661 VTAIL.n182 VTAIL.n181 104.615
R1662 VTAIL.n181 VTAIL.n117 104.615
R1663 VTAIL.n174 VTAIL.n117 104.615
R1664 VTAIL.n174 VTAIL.n173 104.615
R1665 VTAIL.n173 VTAIL.n121 104.615
R1666 VTAIL.n166 VTAIL.n121 104.615
R1667 VTAIL.n166 VTAIL.n165 104.615
R1668 VTAIL.n165 VTAIL.n125 104.615
R1669 VTAIL.n130 VTAIL.n125 104.615
R1670 VTAIL.n158 VTAIL.n130 104.615
R1671 VTAIL.n158 VTAIL.n157 104.615
R1672 VTAIL.n157 VTAIL.n131 104.615
R1673 VTAIL.n150 VTAIL.n131 104.615
R1674 VTAIL.n150 VTAIL.n149 104.615
R1675 VTAIL.n149 VTAIL.n135 104.615
R1676 VTAIL.n142 VTAIL.n135 104.615
R1677 VTAIL.n142 VTAIL.n141 104.615
R1678 VTAIL.n347 VTAIL.t1 52.3082
R1679 VTAIL.n35 VTAIL.t3 52.3082
R1680 VTAIL.n245 VTAIL.t2 52.3082
R1681 VTAIL.n141 VTAIL.t0 52.3082
R1682 VTAIL.n415 VTAIL.n414 36.0641
R1683 VTAIL.n103 VTAIL.n102 36.0641
R1684 VTAIL.n311 VTAIL.n310 36.0641
R1685 VTAIL.n207 VTAIL.n206 36.0641
R1686 VTAIL.n207 VTAIL.n103 32.0393
R1687 VTAIL.n415 VTAIL.n311 30.3152
R1688 VTAIL.n367 VTAIL.n334 13.1884
R1689 VTAIL.n55 VTAIL.n22 13.1884
R1690 VTAIL.n232 VTAIL.n230 13.1884
R1691 VTAIL.n128 VTAIL.n126 13.1884
R1692 VTAIL.n368 VTAIL.n336 12.8005
R1693 VTAIL.n372 VTAIL.n371 12.8005
R1694 VTAIL.n412 VTAIL.n312 12.8005
R1695 VTAIL.n56 VTAIL.n24 12.8005
R1696 VTAIL.n60 VTAIL.n59 12.8005
R1697 VTAIL.n100 VTAIL.n0 12.8005
R1698 VTAIL.n308 VTAIL.n208 12.8005
R1699 VTAIL.n268 VTAIL.n267 12.8005
R1700 VTAIL.n264 VTAIL.n263 12.8005
R1701 VTAIL.n204 VTAIL.n104 12.8005
R1702 VTAIL.n164 VTAIL.n163 12.8005
R1703 VTAIL.n160 VTAIL.n159 12.8005
R1704 VTAIL.n363 VTAIL.n362 12.0247
R1705 VTAIL.n375 VTAIL.n332 12.0247
R1706 VTAIL.n411 VTAIL.n314 12.0247
R1707 VTAIL.n51 VTAIL.n50 12.0247
R1708 VTAIL.n63 VTAIL.n20 12.0247
R1709 VTAIL.n99 VTAIL.n2 12.0247
R1710 VTAIL.n307 VTAIL.n210 12.0247
R1711 VTAIL.n271 VTAIL.n228 12.0247
R1712 VTAIL.n260 VTAIL.n233 12.0247
R1713 VTAIL.n203 VTAIL.n106 12.0247
R1714 VTAIL.n167 VTAIL.n124 12.0247
R1715 VTAIL.n156 VTAIL.n129 12.0247
R1716 VTAIL.n361 VTAIL.n338 11.249
R1717 VTAIL.n376 VTAIL.n330 11.249
R1718 VTAIL.n408 VTAIL.n407 11.249
R1719 VTAIL.n49 VTAIL.n26 11.249
R1720 VTAIL.n64 VTAIL.n18 11.249
R1721 VTAIL.n96 VTAIL.n95 11.249
R1722 VTAIL.n304 VTAIL.n303 11.249
R1723 VTAIL.n272 VTAIL.n226 11.249
R1724 VTAIL.n259 VTAIL.n236 11.249
R1725 VTAIL.n200 VTAIL.n199 11.249
R1726 VTAIL.n168 VTAIL.n122 11.249
R1727 VTAIL.n155 VTAIL.n132 11.249
R1728 VTAIL.n358 VTAIL.n357 10.4732
R1729 VTAIL.n380 VTAIL.n379 10.4732
R1730 VTAIL.n404 VTAIL.n316 10.4732
R1731 VTAIL.n46 VTAIL.n45 10.4732
R1732 VTAIL.n68 VTAIL.n67 10.4732
R1733 VTAIL.n92 VTAIL.n4 10.4732
R1734 VTAIL.n300 VTAIL.n212 10.4732
R1735 VTAIL.n276 VTAIL.n275 10.4732
R1736 VTAIL.n256 VTAIL.n255 10.4732
R1737 VTAIL.n196 VTAIL.n108 10.4732
R1738 VTAIL.n172 VTAIL.n171 10.4732
R1739 VTAIL.n152 VTAIL.n151 10.4732
R1740 VTAIL.n346 VTAIL.n345 10.2747
R1741 VTAIL.n34 VTAIL.n33 10.2747
R1742 VTAIL.n244 VTAIL.n243 10.2747
R1743 VTAIL.n140 VTAIL.n139 10.2747
R1744 VTAIL.n354 VTAIL.n340 9.69747
R1745 VTAIL.n383 VTAIL.n328 9.69747
R1746 VTAIL.n403 VTAIL.n318 9.69747
R1747 VTAIL.n42 VTAIL.n28 9.69747
R1748 VTAIL.n71 VTAIL.n16 9.69747
R1749 VTAIL.n91 VTAIL.n6 9.69747
R1750 VTAIL.n299 VTAIL.n214 9.69747
R1751 VTAIL.n279 VTAIL.n224 9.69747
R1752 VTAIL.n252 VTAIL.n238 9.69747
R1753 VTAIL.n195 VTAIL.n110 9.69747
R1754 VTAIL.n175 VTAIL.n120 9.69747
R1755 VTAIL.n148 VTAIL.n134 9.69747
R1756 VTAIL.n410 VTAIL.n312 9.45567
R1757 VTAIL.n98 VTAIL.n0 9.45567
R1758 VTAIL.n306 VTAIL.n208 9.45567
R1759 VTAIL.n202 VTAIL.n104 9.45567
R1760 VTAIL.n393 VTAIL.n392 9.3005
R1761 VTAIL.n395 VTAIL.n394 9.3005
R1762 VTAIL.n320 VTAIL.n319 9.3005
R1763 VTAIL.n401 VTAIL.n400 9.3005
R1764 VTAIL.n403 VTAIL.n402 9.3005
R1765 VTAIL.n316 VTAIL.n315 9.3005
R1766 VTAIL.n409 VTAIL.n408 9.3005
R1767 VTAIL.n411 VTAIL.n410 9.3005
R1768 VTAIL.n387 VTAIL.n386 9.3005
R1769 VTAIL.n385 VTAIL.n384 9.3005
R1770 VTAIL.n328 VTAIL.n327 9.3005
R1771 VTAIL.n379 VTAIL.n378 9.3005
R1772 VTAIL.n377 VTAIL.n376 9.3005
R1773 VTAIL.n332 VTAIL.n331 9.3005
R1774 VTAIL.n371 VTAIL.n370 9.3005
R1775 VTAIL.n344 VTAIL.n343 9.3005
R1776 VTAIL.n351 VTAIL.n350 9.3005
R1777 VTAIL.n353 VTAIL.n352 9.3005
R1778 VTAIL.n340 VTAIL.n339 9.3005
R1779 VTAIL.n359 VTAIL.n358 9.3005
R1780 VTAIL.n361 VTAIL.n360 9.3005
R1781 VTAIL.n362 VTAIL.n335 9.3005
R1782 VTAIL.n369 VTAIL.n368 9.3005
R1783 VTAIL.n324 VTAIL.n323 9.3005
R1784 VTAIL.n81 VTAIL.n80 9.3005
R1785 VTAIL.n83 VTAIL.n82 9.3005
R1786 VTAIL.n8 VTAIL.n7 9.3005
R1787 VTAIL.n89 VTAIL.n88 9.3005
R1788 VTAIL.n91 VTAIL.n90 9.3005
R1789 VTAIL.n4 VTAIL.n3 9.3005
R1790 VTAIL.n97 VTAIL.n96 9.3005
R1791 VTAIL.n99 VTAIL.n98 9.3005
R1792 VTAIL.n75 VTAIL.n74 9.3005
R1793 VTAIL.n73 VTAIL.n72 9.3005
R1794 VTAIL.n16 VTAIL.n15 9.3005
R1795 VTAIL.n67 VTAIL.n66 9.3005
R1796 VTAIL.n65 VTAIL.n64 9.3005
R1797 VTAIL.n20 VTAIL.n19 9.3005
R1798 VTAIL.n59 VTAIL.n58 9.3005
R1799 VTAIL.n32 VTAIL.n31 9.3005
R1800 VTAIL.n39 VTAIL.n38 9.3005
R1801 VTAIL.n41 VTAIL.n40 9.3005
R1802 VTAIL.n28 VTAIL.n27 9.3005
R1803 VTAIL.n47 VTAIL.n46 9.3005
R1804 VTAIL.n49 VTAIL.n48 9.3005
R1805 VTAIL.n50 VTAIL.n23 9.3005
R1806 VTAIL.n57 VTAIL.n56 9.3005
R1807 VTAIL.n12 VTAIL.n11 9.3005
R1808 VTAIL.n307 VTAIL.n306 9.3005
R1809 VTAIL.n305 VTAIL.n304 9.3005
R1810 VTAIL.n212 VTAIL.n211 9.3005
R1811 VTAIL.n299 VTAIL.n298 9.3005
R1812 VTAIL.n297 VTAIL.n296 9.3005
R1813 VTAIL.n216 VTAIL.n215 9.3005
R1814 VTAIL.n291 VTAIL.n290 9.3005
R1815 VTAIL.n289 VTAIL.n288 9.3005
R1816 VTAIL.n220 VTAIL.n219 9.3005
R1817 VTAIL.n283 VTAIL.n282 9.3005
R1818 VTAIL.n281 VTAIL.n280 9.3005
R1819 VTAIL.n224 VTAIL.n223 9.3005
R1820 VTAIL.n275 VTAIL.n274 9.3005
R1821 VTAIL.n273 VTAIL.n272 9.3005
R1822 VTAIL.n228 VTAIL.n227 9.3005
R1823 VTAIL.n267 VTAIL.n266 9.3005
R1824 VTAIL.n265 VTAIL.n264 9.3005
R1825 VTAIL.n233 VTAIL.n231 9.3005
R1826 VTAIL.n259 VTAIL.n258 9.3005
R1827 VTAIL.n257 VTAIL.n256 9.3005
R1828 VTAIL.n238 VTAIL.n237 9.3005
R1829 VTAIL.n251 VTAIL.n250 9.3005
R1830 VTAIL.n249 VTAIL.n248 9.3005
R1831 VTAIL.n242 VTAIL.n241 9.3005
R1832 VTAIL.n138 VTAIL.n137 9.3005
R1833 VTAIL.n145 VTAIL.n144 9.3005
R1834 VTAIL.n147 VTAIL.n146 9.3005
R1835 VTAIL.n134 VTAIL.n133 9.3005
R1836 VTAIL.n153 VTAIL.n152 9.3005
R1837 VTAIL.n155 VTAIL.n154 9.3005
R1838 VTAIL.n129 VTAIL.n127 9.3005
R1839 VTAIL.n161 VTAIL.n160 9.3005
R1840 VTAIL.n187 VTAIL.n186 9.3005
R1841 VTAIL.n112 VTAIL.n111 9.3005
R1842 VTAIL.n193 VTAIL.n192 9.3005
R1843 VTAIL.n195 VTAIL.n194 9.3005
R1844 VTAIL.n108 VTAIL.n107 9.3005
R1845 VTAIL.n201 VTAIL.n200 9.3005
R1846 VTAIL.n203 VTAIL.n202 9.3005
R1847 VTAIL.n185 VTAIL.n184 9.3005
R1848 VTAIL.n116 VTAIL.n115 9.3005
R1849 VTAIL.n179 VTAIL.n178 9.3005
R1850 VTAIL.n177 VTAIL.n176 9.3005
R1851 VTAIL.n120 VTAIL.n119 9.3005
R1852 VTAIL.n171 VTAIL.n170 9.3005
R1853 VTAIL.n169 VTAIL.n168 9.3005
R1854 VTAIL.n124 VTAIL.n123 9.3005
R1855 VTAIL.n163 VTAIL.n162 9.3005
R1856 VTAIL.n353 VTAIL.n342 8.92171
R1857 VTAIL.n384 VTAIL.n326 8.92171
R1858 VTAIL.n400 VTAIL.n399 8.92171
R1859 VTAIL.n41 VTAIL.n30 8.92171
R1860 VTAIL.n72 VTAIL.n14 8.92171
R1861 VTAIL.n88 VTAIL.n87 8.92171
R1862 VTAIL.n296 VTAIL.n295 8.92171
R1863 VTAIL.n280 VTAIL.n222 8.92171
R1864 VTAIL.n251 VTAIL.n240 8.92171
R1865 VTAIL.n192 VTAIL.n191 8.92171
R1866 VTAIL.n176 VTAIL.n118 8.92171
R1867 VTAIL.n147 VTAIL.n136 8.92171
R1868 VTAIL.n350 VTAIL.n349 8.14595
R1869 VTAIL.n388 VTAIL.n387 8.14595
R1870 VTAIL.n396 VTAIL.n320 8.14595
R1871 VTAIL.n38 VTAIL.n37 8.14595
R1872 VTAIL.n76 VTAIL.n75 8.14595
R1873 VTAIL.n84 VTAIL.n8 8.14595
R1874 VTAIL.n292 VTAIL.n216 8.14595
R1875 VTAIL.n284 VTAIL.n283 8.14595
R1876 VTAIL.n248 VTAIL.n247 8.14595
R1877 VTAIL.n188 VTAIL.n112 8.14595
R1878 VTAIL.n180 VTAIL.n179 8.14595
R1879 VTAIL.n144 VTAIL.n143 8.14595
R1880 VTAIL.n346 VTAIL.n344 7.3702
R1881 VTAIL.n391 VTAIL.n324 7.3702
R1882 VTAIL.n395 VTAIL.n322 7.3702
R1883 VTAIL.n34 VTAIL.n32 7.3702
R1884 VTAIL.n79 VTAIL.n12 7.3702
R1885 VTAIL.n83 VTAIL.n10 7.3702
R1886 VTAIL.n291 VTAIL.n218 7.3702
R1887 VTAIL.n287 VTAIL.n220 7.3702
R1888 VTAIL.n244 VTAIL.n242 7.3702
R1889 VTAIL.n187 VTAIL.n114 7.3702
R1890 VTAIL.n183 VTAIL.n116 7.3702
R1891 VTAIL.n140 VTAIL.n138 7.3702
R1892 VTAIL.n392 VTAIL.n391 6.59444
R1893 VTAIL.n392 VTAIL.n322 6.59444
R1894 VTAIL.n80 VTAIL.n79 6.59444
R1895 VTAIL.n80 VTAIL.n10 6.59444
R1896 VTAIL.n288 VTAIL.n218 6.59444
R1897 VTAIL.n288 VTAIL.n287 6.59444
R1898 VTAIL.n184 VTAIL.n114 6.59444
R1899 VTAIL.n184 VTAIL.n183 6.59444
R1900 VTAIL.n349 VTAIL.n344 5.81868
R1901 VTAIL.n388 VTAIL.n324 5.81868
R1902 VTAIL.n396 VTAIL.n395 5.81868
R1903 VTAIL.n37 VTAIL.n32 5.81868
R1904 VTAIL.n76 VTAIL.n12 5.81868
R1905 VTAIL.n84 VTAIL.n83 5.81868
R1906 VTAIL.n292 VTAIL.n291 5.81868
R1907 VTAIL.n284 VTAIL.n220 5.81868
R1908 VTAIL.n247 VTAIL.n242 5.81868
R1909 VTAIL.n188 VTAIL.n187 5.81868
R1910 VTAIL.n180 VTAIL.n116 5.81868
R1911 VTAIL.n143 VTAIL.n138 5.81868
R1912 VTAIL.n350 VTAIL.n342 5.04292
R1913 VTAIL.n387 VTAIL.n326 5.04292
R1914 VTAIL.n399 VTAIL.n320 5.04292
R1915 VTAIL.n38 VTAIL.n30 5.04292
R1916 VTAIL.n75 VTAIL.n14 5.04292
R1917 VTAIL.n87 VTAIL.n8 5.04292
R1918 VTAIL.n295 VTAIL.n216 5.04292
R1919 VTAIL.n283 VTAIL.n222 5.04292
R1920 VTAIL.n248 VTAIL.n240 5.04292
R1921 VTAIL.n191 VTAIL.n112 5.04292
R1922 VTAIL.n179 VTAIL.n118 5.04292
R1923 VTAIL.n144 VTAIL.n136 5.04292
R1924 VTAIL.n354 VTAIL.n353 4.26717
R1925 VTAIL.n384 VTAIL.n383 4.26717
R1926 VTAIL.n400 VTAIL.n318 4.26717
R1927 VTAIL.n42 VTAIL.n41 4.26717
R1928 VTAIL.n72 VTAIL.n71 4.26717
R1929 VTAIL.n88 VTAIL.n6 4.26717
R1930 VTAIL.n296 VTAIL.n214 4.26717
R1931 VTAIL.n280 VTAIL.n279 4.26717
R1932 VTAIL.n252 VTAIL.n251 4.26717
R1933 VTAIL.n192 VTAIL.n110 4.26717
R1934 VTAIL.n176 VTAIL.n175 4.26717
R1935 VTAIL.n148 VTAIL.n147 4.26717
R1936 VTAIL.n357 VTAIL.n340 3.49141
R1937 VTAIL.n380 VTAIL.n328 3.49141
R1938 VTAIL.n404 VTAIL.n403 3.49141
R1939 VTAIL.n45 VTAIL.n28 3.49141
R1940 VTAIL.n68 VTAIL.n16 3.49141
R1941 VTAIL.n92 VTAIL.n91 3.49141
R1942 VTAIL.n300 VTAIL.n299 3.49141
R1943 VTAIL.n276 VTAIL.n224 3.49141
R1944 VTAIL.n255 VTAIL.n238 3.49141
R1945 VTAIL.n196 VTAIL.n195 3.49141
R1946 VTAIL.n172 VTAIL.n120 3.49141
R1947 VTAIL.n151 VTAIL.n134 3.49141
R1948 VTAIL.n345 VTAIL.n343 2.84303
R1949 VTAIL.n33 VTAIL.n31 2.84303
R1950 VTAIL.n243 VTAIL.n241 2.84303
R1951 VTAIL.n139 VTAIL.n137 2.84303
R1952 VTAIL.n358 VTAIL.n338 2.71565
R1953 VTAIL.n379 VTAIL.n330 2.71565
R1954 VTAIL.n407 VTAIL.n316 2.71565
R1955 VTAIL.n46 VTAIL.n26 2.71565
R1956 VTAIL.n67 VTAIL.n18 2.71565
R1957 VTAIL.n95 VTAIL.n4 2.71565
R1958 VTAIL.n303 VTAIL.n212 2.71565
R1959 VTAIL.n275 VTAIL.n226 2.71565
R1960 VTAIL.n256 VTAIL.n236 2.71565
R1961 VTAIL.n199 VTAIL.n108 2.71565
R1962 VTAIL.n171 VTAIL.n122 2.71565
R1963 VTAIL.n152 VTAIL.n132 2.71565
R1964 VTAIL.n363 VTAIL.n361 1.93989
R1965 VTAIL.n376 VTAIL.n375 1.93989
R1966 VTAIL.n408 VTAIL.n314 1.93989
R1967 VTAIL.n51 VTAIL.n49 1.93989
R1968 VTAIL.n64 VTAIL.n63 1.93989
R1969 VTAIL.n96 VTAIL.n2 1.93989
R1970 VTAIL.n304 VTAIL.n210 1.93989
R1971 VTAIL.n272 VTAIL.n271 1.93989
R1972 VTAIL.n260 VTAIL.n259 1.93989
R1973 VTAIL.n200 VTAIL.n106 1.93989
R1974 VTAIL.n168 VTAIL.n167 1.93989
R1975 VTAIL.n156 VTAIL.n155 1.93989
R1976 VTAIL.n311 VTAIL.n207 1.3324
R1977 VTAIL.n362 VTAIL.n336 1.16414
R1978 VTAIL.n372 VTAIL.n332 1.16414
R1979 VTAIL.n412 VTAIL.n411 1.16414
R1980 VTAIL.n50 VTAIL.n24 1.16414
R1981 VTAIL.n60 VTAIL.n20 1.16414
R1982 VTAIL.n100 VTAIL.n99 1.16414
R1983 VTAIL.n308 VTAIL.n307 1.16414
R1984 VTAIL.n268 VTAIL.n228 1.16414
R1985 VTAIL.n263 VTAIL.n233 1.16414
R1986 VTAIL.n204 VTAIL.n203 1.16414
R1987 VTAIL.n164 VTAIL.n124 1.16414
R1988 VTAIL.n159 VTAIL.n129 1.16414
R1989 VTAIL VTAIL.n103 0.959552
R1990 VTAIL.n368 VTAIL.n367 0.388379
R1991 VTAIL.n371 VTAIL.n334 0.388379
R1992 VTAIL.n414 VTAIL.n312 0.388379
R1993 VTAIL.n56 VTAIL.n55 0.388379
R1994 VTAIL.n59 VTAIL.n22 0.388379
R1995 VTAIL.n102 VTAIL.n0 0.388379
R1996 VTAIL.n310 VTAIL.n208 0.388379
R1997 VTAIL.n267 VTAIL.n230 0.388379
R1998 VTAIL.n264 VTAIL.n232 0.388379
R1999 VTAIL.n206 VTAIL.n104 0.388379
R2000 VTAIL.n163 VTAIL.n126 0.388379
R2001 VTAIL.n160 VTAIL.n128 0.388379
R2002 VTAIL VTAIL.n415 0.373345
R2003 VTAIL.n351 VTAIL.n343 0.155672
R2004 VTAIL.n352 VTAIL.n351 0.155672
R2005 VTAIL.n352 VTAIL.n339 0.155672
R2006 VTAIL.n359 VTAIL.n339 0.155672
R2007 VTAIL.n360 VTAIL.n359 0.155672
R2008 VTAIL.n360 VTAIL.n335 0.155672
R2009 VTAIL.n369 VTAIL.n335 0.155672
R2010 VTAIL.n370 VTAIL.n369 0.155672
R2011 VTAIL.n370 VTAIL.n331 0.155672
R2012 VTAIL.n377 VTAIL.n331 0.155672
R2013 VTAIL.n378 VTAIL.n377 0.155672
R2014 VTAIL.n378 VTAIL.n327 0.155672
R2015 VTAIL.n385 VTAIL.n327 0.155672
R2016 VTAIL.n386 VTAIL.n385 0.155672
R2017 VTAIL.n386 VTAIL.n323 0.155672
R2018 VTAIL.n393 VTAIL.n323 0.155672
R2019 VTAIL.n394 VTAIL.n393 0.155672
R2020 VTAIL.n394 VTAIL.n319 0.155672
R2021 VTAIL.n401 VTAIL.n319 0.155672
R2022 VTAIL.n402 VTAIL.n401 0.155672
R2023 VTAIL.n402 VTAIL.n315 0.155672
R2024 VTAIL.n409 VTAIL.n315 0.155672
R2025 VTAIL.n410 VTAIL.n409 0.155672
R2026 VTAIL.n39 VTAIL.n31 0.155672
R2027 VTAIL.n40 VTAIL.n39 0.155672
R2028 VTAIL.n40 VTAIL.n27 0.155672
R2029 VTAIL.n47 VTAIL.n27 0.155672
R2030 VTAIL.n48 VTAIL.n47 0.155672
R2031 VTAIL.n48 VTAIL.n23 0.155672
R2032 VTAIL.n57 VTAIL.n23 0.155672
R2033 VTAIL.n58 VTAIL.n57 0.155672
R2034 VTAIL.n58 VTAIL.n19 0.155672
R2035 VTAIL.n65 VTAIL.n19 0.155672
R2036 VTAIL.n66 VTAIL.n65 0.155672
R2037 VTAIL.n66 VTAIL.n15 0.155672
R2038 VTAIL.n73 VTAIL.n15 0.155672
R2039 VTAIL.n74 VTAIL.n73 0.155672
R2040 VTAIL.n74 VTAIL.n11 0.155672
R2041 VTAIL.n81 VTAIL.n11 0.155672
R2042 VTAIL.n82 VTAIL.n81 0.155672
R2043 VTAIL.n82 VTAIL.n7 0.155672
R2044 VTAIL.n89 VTAIL.n7 0.155672
R2045 VTAIL.n90 VTAIL.n89 0.155672
R2046 VTAIL.n90 VTAIL.n3 0.155672
R2047 VTAIL.n97 VTAIL.n3 0.155672
R2048 VTAIL.n98 VTAIL.n97 0.155672
R2049 VTAIL.n306 VTAIL.n305 0.155672
R2050 VTAIL.n305 VTAIL.n211 0.155672
R2051 VTAIL.n298 VTAIL.n211 0.155672
R2052 VTAIL.n298 VTAIL.n297 0.155672
R2053 VTAIL.n297 VTAIL.n215 0.155672
R2054 VTAIL.n290 VTAIL.n215 0.155672
R2055 VTAIL.n290 VTAIL.n289 0.155672
R2056 VTAIL.n289 VTAIL.n219 0.155672
R2057 VTAIL.n282 VTAIL.n219 0.155672
R2058 VTAIL.n282 VTAIL.n281 0.155672
R2059 VTAIL.n281 VTAIL.n223 0.155672
R2060 VTAIL.n274 VTAIL.n223 0.155672
R2061 VTAIL.n274 VTAIL.n273 0.155672
R2062 VTAIL.n273 VTAIL.n227 0.155672
R2063 VTAIL.n266 VTAIL.n227 0.155672
R2064 VTAIL.n266 VTAIL.n265 0.155672
R2065 VTAIL.n265 VTAIL.n231 0.155672
R2066 VTAIL.n258 VTAIL.n231 0.155672
R2067 VTAIL.n258 VTAIL.n257 0.155672
R2068 VTAIL.n257 VTAIL.n237 0.155672
R2069 VTAIL.n250 VTAIL.n237 0.155672
R2070 VTAIL.n250 VTAIL.n249 0.155672
R2071 VTAIL.n249 VTAIL.n241 0.155672
R2072 VTAIL.n202 VTAIL.n201 0.155672
R2073 VTAIL.n201 VTAIL.n107 0.155672
R2074 VTAIL.n194 VTAIL.n107 0.155672
R2075 VTAIL.n194 VTAIL.n193 0.155672
R2076 VTAIL.n193 VTAIL.n111 0.155672
R2077 VTAIL.n186 VTAIL.n111 0.155672
R2078 VTAIL.n186 VTAIL.n185 0.155672
R2079 VTAIL.n185 VTAIL.n115 0.155672
R2080 VTAIL.n178 VTAIL.n115 0.155672
R2081 VTAIL.n178 VTAIL.n177 0.155672
R2082 VTAIL.n177 VTAIL.n119 0.155672
R2083 VTAIL.n170 VTAIL.n119 0.155672
R2084 VTAIL.n170 VTAIL.n169 0.155672
R2085 VTAIL.n169 VTAIL.n123 0.155672
R2086 VTAIL.n162 VTAIL.n123 0.155672
R2087 VTAIL.n162 VTAIL.n161 0.155672
R2088 VTAIL.n161 VTAIL.n127 0.155672
R2089 VTAIL.n154 VTAIL.n127 0.155672
R2090 VTAIL.n154 VTAIL.n153 0.155672
R2091 VTAIL.n153 VTAIL.n133 0.155672
R2092 VTAIL.n146 VTAIL.n133 0.155672
R2093 VTAIL.n146 VTAIL.n145 0.155672
R2094 VTAIL.n145 VTAIL.n137 0.155672
R2095 VDD1.n102 VDD1.n101 289.615
R2096 VDD1.n205 VDD1.n204 289.615
R2097 VDD1.n101 VDD1.n100 185
R2098 VDD1.n2 VDD1.n1 185
R2099 VDD1.n95 VDD1.n94 185
R2100 VDD1.n93 VDD1.n92 185
R2101 VDD1.n6 VDD1.n5 185
R2102 VDD1.n87 VDD1.n86 185
R2103 VDD1.n85 VDD1.n84 185
R2104 VDD1.n10 VDD1.n9 185
R2105 VDD1.n79 VDD1.n78 185
R2106 VDD1.n77 VDD1.n76 185
R2107 VDD1.n14 VDD1.n13 185
R2108 VDD1.n71 VDD1.n70 185
R2109 VDD1.n69 VDD1.n68 185
R2110 VDD1.n18 VDD1.n17 185
R2111 VDD1.n63 VDD1.n62 185
R2112 VDD1.n61 VDD1.n60 185
R2113 VDD1.n22 VDD1.n21 185
R2114 VDD1.n26 VDD1.n24 185
R2115 VDD1.n55 VDD1.n54 185
R2116 VDD1.n53 VDD1.n52 185
R2117 VDD1.n28 VDD1.n27 185
R2118 VDD1.n47 VDD1.n46 185
R2119 VDD1.n45 VDD1.n44 185
R2120 VDD1.n32 VDD1.n31 185
R2121 VDD1.n39 VDD1.n38 185
R2122 VDD1.n37 VDD1.n36 185
R2123 VDD1.n138 VDD1.n137 185
R2124 VDD1.n140 VDD1.n139 185
R2125 VDD1.n133 VDD1.n132 185
R2126 VDD1.n146 VDD1.n145 185
R2127 VDD1.n148 VDD1.n147 185
R2128 VDD1.n129 VDD1.n128 185
R2129 VDD1.n155 VDD1.n154 185
R2130 VDD1.n156 VDD1.n127 185
R2131 VDD1.n158 VDD1.n157 185
R2132 VDD1.n125 VDD1.n124 185
R2133 VDD1.n164 VDD1.n163 185
R2134 VDD1.n166 VDD1.n165 185
R2135 VDD1.n121 VDD1.n120 185
R2136 VDD1.n172 VDD1.n171 185
R2137 VDD1.n174 VDD1.n173 185
R2138 VDD1.n117 VDD1.n116 185
R2139 VDD1.n180 VDD1.n179 185
R2140 VDD1.n182 VDD1.n181 185
R2141 VDD1.n113 VDD1.n112 185
R2142 VDD1.n188 VDD1.n187 185
R2143 VDD1.n190 VDD1.n189 185
R2144 VDD1.n109 VDD1.n108 185
R2145 VDD1.n196 VDD1.n195 185
R2146 VDD1.n198 VDD1.n197 185
R2147 VDD1.n105 VDD1.n104 185
R2148 VDD1.n204 VDD1.n203 185
R2149 VDD1.n35 VDD1.t0 149.524
R2150 VDD1.n136 VDD1.t1 149.524
R2151 VDD1.n101 VDD1.n1 104.615
R2152 VDD1.n94 VDD1.n1 104.615
R2153 VDD1.n94 VDD1.n93 104.615
R2154 VDD1.n93 VDD1.n5 104.615
R2155 VDD1.n86 VDD1.n5 104.615
R2156 VDD1.n86 VDD1.n85 104.615
R2157 VDD1.n85 VDD1.n9 104.615
R2158 VDD1.n78 VDD1.n9 104.615
R2159 VDD1.n78 VDD1.n77 104.615
R2160 VDD1.n77 VDD1.n13 104.615
R2161 VDD1.n70 VDD1.n13 104.615
R2162 VDD1.n70 VDD1.n69 104.615
R2163 VDD1.n69 VDD1.n17 104.615
R2164 VDD1.n62 VDD1.n17 104.615
R2165 VDD1.n62 VDD1.n61 104.615
R2166 VDD1.n61 VDD1.n21 104.615
R2167 VDD1.n26 VDD1.n21 104.615
R2168 VDD1.n54 VDD1.n26 104.615
R2169 VDD1.n54 VDD1.n53 104.615
R2170 VDD1.n53 VDD1.n27 104.615
R2171 VDD1.n46 VDD1.n27 104.615
R2172 VDD1.n46 VDD1.n45 104.615
R2173 VDD1.n45 VDD1.n31 104.615
R2174 VDD1.n38 VDD1.n31 104.615
R2175 VDD1.n38 VDD1.n37 104.615
R2176 VDD1.n139 VDD1.n138 104.615
R2177 VDD1.n139 VDD1.n132 104.615
R2178 VDD1.n146 VDD1.n132 104.615
R2179 VDD1.n147 VDD1.n146 104.615
R2180 VDD1.n147 VDD1.n128 104.615
R2181 VDD1.n155 VDD1.n128 104.615
R2182 VDD1.n156 VDD1.n155 104.615
R2183 VDD1.n157 VDD1.n156 104.615
R2184 VDD1.n157 VDD1.n124 104.615
R2185 VDD1.n164 VDD1.n124 104.615
R2186 VDD1.n165 VDD1.n164 104.615
R2187 VDD1.n165 VDD1.n120 104.615
R2188 VDD1.n172 VDD1.n120 104.615
R2189 VDD1.n173 VDD1.n172 104.615
R2190 VDD1.n173 VDD1.n116 104.615
R2191 VDD1.n180 VDD1.n116 104.615
R2192 VDD1.n181 VDD1.n180 104.615
R2193 VDD1.n181 VDD1.n112 104.615
R2194 VDD1.n188 VDD1.n112 104.615
R2195 VDD1.n189 VDD1.n188 104.615
R2196 VDD1.n189 VDD1.n108 104.615
R2197 VDD1.n196 VDD1.n108 104.615
R2198 VDD1.n197 VDD1.n196 104.615
R2199 VDD1.n197 VDD1.n104 104.615
R2200 VDD1.n204 VDD1.n104 104.615
R2201 VDD1 VDD1.n205 97.0307
R2202 VDD1 VDD1.n102 53.2321
R2203 VDD1.n37 VDD1.t0 52.3082
R2204 VDD1.n138 VDD1.t1 52.3082
R2205 VDD1.n24 VDD1.n22 13.1884
R2206 VDD1.n158 VDD1.n125 13.1884
R2207 VDD1.n100 VDD1.n0 12.8005
R2208 VDD1.n60 VDD1.n59 12.8005
R2209 VDD1.n56 VDD1.n55 12.8005
R2210 VDD1.n159 VDD1.n127 12.8005
R2211 VDD1.n163 VDD1.n162 12.8005
R2212 VDD1.n203 VDD1.n103 12.8005
R2213 VDD1.n99 VDD1.n2 12.0247
R2214 VDD1.n63 VDD1.n20 12.0247
R2215 VDD1.n52 VDD1.n25 12.0247
R2216 VDD1.n154 VDD1.n153 12.0247
R2217 VDD1.n166 VDD1.n123 12.0247
R2218 VDD1.n202 VDD1.n105 12.0247
R2219 VDD1.n96 VDD1.n95 11.249
R2220 VDD1.n64 VDD1.n18 11.249
R2221 VDD1.n51 VDD1.n28 11.249
R2222 VDD1.n152 VDD1.n129 11.249
R2223 VDD1.n167 VDD1.n121 11.249
R2224 VDD1.n199 VDD1.n198 11.249
R2225 VDD1.n92 VDD1.n4 10.4732
R2226 VDD1.n68 VDD1.n67 10.4732
R2227 VDD1.n48 VDD1.n47 10.4732
R2228 VDD1.n149 VDD1.n148 10.4732
R2229 VDD1.n171 VDD1.n170 10.4732
R2230 VDD1.n195 VDD1.n107 10.4732
R2231 VDD1.n36 VDD1.n35 10.2747
R2232 VDD1.n137 VDD1.n136 10.2747
R2233 VDD1.n91 VDD1.n6 9.69747
R2234 VDD1.n71 VDD1.n16 9.69747
R2235 VDD1.n44 VDD1.n30 9.69747
R2236 VDD1.n145 VDD1.n131 9.69747
R2237 VDD1.n174 VDD1.n119 9.69747
R2238 VDD1.n194 VDD1.n109 9.69747
R2239 VDD1.n98 VDD1.n0 9.45567
R2240 VDD1.n201 VDD1.n103 9.45567
R2241 VDD1.n99 VDD1.n98 9.3005
R2242 VDD1.n97 VDD1.n96 9.3005
R2243 VDD1.n4 VDD1.n3 9.3005
R2244 VDD1.n91 VDD1.n90 9.3005
R2245 VDD1.n89 VDD1.n88 9.3005
R2246 VDD1.n8 VDD1.n7 9.3005
R2247 VDD1.n83 VDD1.n82 9.3005
R2248 VDD1.n81 VDD1.n80 9.3005
R2249 VDD1.n12 VDD1.n11 9.3005
R2250 VDD1.n75 VDD1.n74 9.3005
R2251 VDD1.n73 VDD1.n72 9.3005
R2252 VDD1.n16 VDD1.n15 9.3005
R2253 VDD1.n67 VDD1.n66 9.3005
R2254 VDD1.n65 VDD1.n64 9.3005
R2255 VDD1.n20 VDD1.n19 9.3005
R2256 VDD1.n59 VDD1.n58 9.3005
R2257 VDD1.n57 VDD1.n56 9.3005
R2258 VDD1.n25 VDD1.n23 9.3005
R2259 VDD1.n51 VDD1.n50 9.3005
R2260 VDD1.n49 VDD1.n48 9.3005
R2261 VDD1.n30 VDD1.n29 9.3005
R2262 VDD1.n43 VDD1.n42 9.3005
R2263 VDD1.n41 VDD1.n40 9.3005
R2264 VDD1.n34 VDD1.n33 9.3005
R2265 VDD1.n184 VDD1.n183 9.3005
R2266 VDD1.n186 VDD1.n185 9.3005
R2267 VDD1.n111 VDD1.n110 9.3005
R2268 VDD1.n192 VDD1.n191 9.3005
R2269 VDD1.n194 VDD1.n193 9.3005
R2270 VDD1.n107 VDD1.n106 9.3005
R2271 VDD1.n200 VDD1.n199 9.3005
R2272 VDD1.n202 VDD1.n201 9.3005
R2273 VDD1.n178 VDD1.n177 9.3005
R2274 VDD1.n176 VDD1.n175 9.3005
R2275 VDD1.n119 VDD1.n118 9.3005
R2276 VDD1.n170 VDD1.n169 9.3005
R2277 VDD1.n168 VDD1.n167 9.3005
R2278 VDD1.n123 VDD1.n122 9.3005
R2279 VDD1.n162 VDD1.n161 9.3005
R2280 VDD1.n135 VDD1.n134 9.3005
R2281 VDD1.n142 VDD1.n141 9.3005
R2282 VDD1.n144 VDD1.n143 9.3005
R2283 VDD1.n131 VDD1.n130 9.3005
R2284 VDD1.n150 VDD1.n149 9.3005
R2285 VDD1.n152 VDD1.n151 9.3005
R2286 VDD1.n153 VDD1.n126 9.3005
R2287 VDD1.n160 VDD1.n159 9.3005
R2288 VDD1.n115 VDD1.n114 9.3005
R2289 VDD1.n88 VDD1.n87 8.92171
R2290 VDD1.n72 VDD1.n14 8.92171
R2291 VDD1.n43 VDD1.n32 8.92171
R2292 VDD1.n144 VDD1.n133 8.92171
R2293 VDD1.n175 VDD1.n117 8.92171
R2294 VDD1.n191 VDD1.n190 8.92171
R2295 VDD1.n84 VDD1.n8 8.14595
R2296 VDD1.n76 VDD1.n75 8.14595
R2297 VDD1.n40 VDD1.n39 8.14595
R2298 VDD1.n141 VDD1.n140 8.14595
R2299 VDD1.n179 VDD1.n178 8.14595
R2300 VDD1.n187 VDD1.n111 8.14595
R2301 VDD1.n83 VDD1.n10 7.3702
R2302 VDD1.n79 VDD1.n12 7.3702
R2303 VDD1.n36 VDD1.n34 7.3702
R2304 VDD1.n137 VDD1.n135 7.3702
R2305 VDD1.n182 VDD1.n115 7.3702
R2306 VDD1.n186 VDD1.n113 7.3702
R2307 VDD1.n80 VDD1.n10 6.59444
R2308 VDD1.n80 VDD1.n79 6.59444
R2309 VDD1.n183 VDD1.n182 6.59444
R2310 VDD1.n183 VDD1.n113 6.59444
R2311 VDD1.n84 VDD1.n83 5.81868
R2312 VDD1.n76 VDD1.n12 5.81868
R2313 VDD1.n39 VDD1.n34 5.81868
R2314 VDD1.n140 VDD1.n135 5.81868
R2315 VDD1.n179 VDD1.n115 5.81868
R2316 VDD1.n187 VDD1.n186 5.81868
R2317 VDD1.n87 VDD1.n8 5.04292
R2318 VDD1.n75 VDD1.n14 5.04292
R2319 VDD1.n40 VDD1.n32 5.04292
R2320 VDD1.n141 VDD1.n133 5.04292
R2321 VDD1.n178 VDD1.n117 5.04292
R2322 VDD1.n190 VDD1.n111 5.04292
R2323 VDD1.n88 VDD1.n6 4.26717
R2324 VDD1.n72 VDD1.n71 4.26717
R2325 VDD1.n44 VDD1.n43 4.26717
R2326 VDD1.n145 VDD1.n144 4.26717
R2327 VDD1.n175 VDD1.n174 4.26717
R2328 VDD1.n191 VDD1.n109 4.26717
R2329 VDD1.n92 VDD1.n91 3.49141
R2330 VDD1.n68 VDD1.n16 3.49141
R2331 VDD1.n47 VDD1.n30 3.49141
R2332 VDD1.n148 VDD1.n131 3.49141
R2333 VDD1.n171 VDD1.n119 3.49141
R2334 VDD1.n195 VDD1.n194 3.49141
R2335 VDD1.n136 VDD1.n134 2.84303
R2336 VDD1.n35 VDD1.n33 2.84303
R2337 VDD1.n95 VDD1.n4 2.71565
R2338 VDD1.n67 VDD1.n18 2.71565
R2339 VDD1.n48 VDD1.n28 2.71565
R2340 VDD1.n149 VDD1.n129 2.71565
R2341 VDD1.n170 VDD1.n121 2.71565
R2342 VDD1.n198 VDD1.n107 2.71565
R2343 VDD1.n96 VDD1.n2 1.93989
R2344 VDD1.n64 VDD1.n63 1.93989
R2345 VDD1.n52 VDD1.n51 1.93989
R2346 VDD1.n154 VDD1.n152 1.93989
R2347 VDD1.n167 VDD1.n166 1.93989
R2348 VDD1.n199 VDD1.n105 1.93989
R2349 VDD1.n100 VDD1.n99 1.16414
R2350 VDD1.n60 VDD1.n20 1.16414
R2351 VDD1.n55 VDD1.n25 1.16414
R2352 VDD1.n153 VDD1.n127 1.16414
R2353 VDD1.n163 VDD1.n123 1.16414
R2354 VDD1.n203 VDD1.n202 1.16414
R2355 VDD1.n102 VDD1.n0 0.388379
R2356 VDD1.n59 VDD1.n22 0.388379
R2357 VDD1.n56 VDD1.n24 0.388379
R2358 VDD1.n159 VDD1.n158 0.388379
R2359 VDD1.n162 VDD1.n125 0.388379
R2360 VDD1.n205 VDD1.n103 0.388379
R2361 VDD1.n98 VDD1.n97 0.155672
R2362 VDD1.n97 VDD1.n3 0.155672
R2363 VDD1.n90 VDD1.n3 0.155672
R2364 VDD1.n90 VDD1.n89 0.155672
R2365 VDD1.n89 VDD1.n7 0.155672
R2366 VDD1.n82 VDD1.n7 0.155672
R2367 VDD1.n82 VDD1.n81 0.155672
R2368 VDD1.n81 VDD1.n11 0.155672
R2369 VDD1.n74 VDD1.n11 0.155672
R2370 VDD1.n74 VDD1.n73 0.155672
R2371 VDD1.n73 VDD1.n15 0.155672
R2372 VDD1.n66 VDD1.n15 0.155672
R2373 VDD1.n66 VDD1.n65 0.155672
R2374 VDD1.n65 VDD1.n19 0.155672
R2375 VDD1.n58 VDD1.n19 0.155672
R2376 VDD1.n58 VDD1.n57 0.155672
R2377 VDD1.n57 VDD1.n23 0.155672
R2378 VDD1.n50 VDD1.n23 0.155672
R2379 VDD1.n50 VDD1.n49 0.155672
R2380 VDD1.n49 VDD1.n29 0.155672
R2381 VDD1.n42 VDD1.n29 0.155672
R2382 VDD1.n42 VDD1.n41 0.155672
R2383 VDD1.n41 VDD1.n33 0.155672
R2384 VDD1.n142 VDD1.n134 0.155672
R2385 VDD1.n143 VDD1.n142 0.155672
R2386 VDD1.n143 VDD1.n130 0.155672
R2387 VDD1.n150 VDD1.n130 0.155672
R2388 VDD1.n151 VDD1.n150 0.155672
R2389 VDD1.n151 VDD1.n126 0.155672
R2390 VDD1.n160 VDD1.n126 0.155672
R2391 VDD1.n161 VDD1.n160 0.155672
R2392 VDD1.n161 VDD1.n122 0.155672
R2393 VDD1.n168 VDD1.n122 0.155672
R2394 VDD1.n169 VDD1.n168 0.155672
R2395 VDD1.n169 VDD1.n118 0.155672
R2396 VDD1.n176 VDD1.n118 0.155672
R2397 VDD1.n177 VDD1.n176 0.155672
R2398 VDD1.n177 VDD1.n114 0.155672
R2399 VDD1.n184 VDD1.n114 0.155672
R2400 VDD1.n185 VDD1.n184 0.155672
R2401 VDD1.n185 VDD1.n110 0.155672
R2402 VDD1.n192 VDD1.n110 0.155672
R2403 VDD1.n193 VDD1.n192 0.155672
R2404 VDD1.n193 VDD1.n106 0.155672
R2405 VDD1.n200 VDD1.n106 0.155672
R2406 VDD1.n201 VDD1.n200 0.155672
R2407 VN VN.t1 378.029
R2408 VN VN.t0 330.721
R2409 VDD2.n205 VDD2.n204 289.615
R2410 VDD2.n102 VDD2.n101 289.615
R2411 VDD2.n204 VDD2.n203 185
R2412 VDD2.n105 VDD2.n104 185
R2413 VDD2.n198 VDD2.n197 185
R2414 VDD2.n196 VDD2.n195 185
R2415 VDD2.n109 VDD2.n108 185
R2416 VDD2.n190 VDD2.n189 185
R2417 VDD2.n188 VDD2.n187 185
R2418 VDD2.n113 VDD2.n112 185
R2419 VDD2.n182 VDD2.n181 185
R2420 VDD2.n180 VDD2.n179 185
R2421 VDD2.n117 VDD2.n116 185
R2422 VDD2.n174 VDD2.n173 185
R2423 VDD2.n172 VDD2.n171 185
R2424 VDD2.n121 VDD2.n120 185
R2425 VDD2.n166 VDD2.n165 185
R2426 VDD2.n164 VDD2.n163 185
R2427 VDD2.n125 VDD2.n124 185
R2428 VDD2.n129 VDD2.n127 185
R2429 VDD2.n158 VDD2.n157 185
R2430 VDD2.n156 VDD2.n155 185
R2431 VDD2.n131 VDD2.n130 185
R2432 VDD2.n150 VDD2.n149 185
R2433 VDD2.n148 VDD2.n147 185
R2434 VDD2.n135 VDD2.n134 185
R2435 VDD2.n142 VDD2.n141 185
R2436 VDD2.n140 VDD2.n139 185
R2437 VDD2.n35 VDD2.n34 185
R2438 VDD2.n37 VDD2.n36 185
R2439 VDD2.n30 VDD2.n29 185
R2440 VDD2.n43 VDD2.n42 185
R2441 VDD2.n45 VDD2.n44 185
R2442 VDD2.n26 VDD2.n25 185
R2443 VDD2.n52 VDD2.n51 185
R2444 VDD2.n53 VDD2.n24 185
R2445 VDD2.n55 VDD2.n54 185
R2446 VDD2.n22 VDD2.n21 185
R2447 VDD2.n61 VDD2.n60 185
R2448 VDD2.n63 VDD2.n62 185
R2449 VDD2.n18 VDD2.n17 185
R2450 VDD2.n69 VDD2.n68 185
R2451 VDD2.n71 VDD2.n70 185
R2452 VDD2.n14 VDD2.n13 185
R2453 VDD2.n77 VDD2.n76 185
R2454 VDD2.n79 VDD2.n78 185
R2455 VDD2.n10 VDD2.n9 185
R2456 VDD2.n85 VDD2.n84 185
R2457 VDD2.n87 VDD2.n86 185
R2458 VDD2.n6 VDD2.n5 185
R2459 VDD2.n93 VDD2.n92 185
R2460 VDD2.n95 VDD2.n94 185
R2461 VDD2.n2 VDD2.n1 185
R2462 VDD2.n101 VDD2.n100 185
R2463 VDD2.n138 VDD2.t0 149.524
R2464 VDD2.n33 VDD2.t1 149.524
R2465 VDD2.n204 VDD2.n104 104.615
R2466 VDD2.n197 VDD2.n104 104.615
R2467 VDD2.n197 VDD2.n196 104.615
R2468 VDD2.n196 VDD2.n108 104.615
R2469 VDD2.n189 VDD2.n108 104.615
R2470 VDD2.n189 VDD2.n188 104.615
R2471 VDD2.n188 VDD2.n112 104.615
R2472 VDD2.n181 VDD2.n112 104.615
R2473 VDD2.n181 VDD2.n180 104.615
R2474 VDD2.n180 VDD2.n116 104.615
R2475 VDD2.n173 VDD2.n116 104.615
R2476 VDD2.n173 VDD2.n172 104.615
R2477 VDD2.n172 VDD2.n120 104.615
R2478 VDD2.n165 VDD2.n120 104.615
R2479 VDD2.n165 VDD2.n164 104.615
R2480 VDD2.n164 VDD2.n124 104.615
R2481 VDD2.n129 VDD2.n124 104.615
R2482 VDD2.n157 VDD2.n129 104.615
R2483 VDD2.n157 VDD2.n156 104.615
R2484 VDD2.n156 VDD2.n130 104.615
R2485 VDD2.n149 VDD2.n130 104.615
R2486 VDD2.n149 VDD2.n148 104.615
R2487 VDD2.n148 VDD2.n134 104.615
R2488 VDD2.n141 VDD2.n134 104.615
R2489 VDD2.n141 VDD2.n140 104.615
R2490 VDD2.n36 VDD2.n35 104.615
R2491 VDD2.n36 VDD2.n29 104.615
R2492 VDD2.n43 VDD2.n29 104.615
R2493 VDD2.n44 VDD2.n43 104.615
R2494 VDD2.n44 VDD2.n25 104.615
R2495 VDD2.n52 VDD2.n25 104.615
R2496 VDD2.n53 VDD2.n52 104.615
R2497 VDD2.n54 VDD2.n53 104.615
R2498 VDD2.n54 VDD2.n21 104.615
R2499 VDD2.n61 VDD2.n21 104.615
R2500 VDD2.n62 VDD2.n61 104.615
R2501 VDD2.n62 VDD2.n17 104.615
R2502 VDD2.n69 VDD2.n17 104.615
R2503 VDD2.n70 VDD2.n69 104.615
R2504 VDD2.n70 VDD2.n13 104.615
R2505 VDD2.n77 VDD2.n13 104.615
R2506 VDD2.n78 VDD2.n77 104.615
R2507 VDD2.n78 VDD2.n9 104.615
R2508 VDD2.n85 VDD2.n9 104.615
R2509 VDD2.n86 VDD2.n85 104.615
R2510 VDD2.n86 VDD2.n5 104.615
R2511 VDD2.n93 VDD2.n5 104.615
R2512 VDD2.n94 VDD2.n93 104.615
R2513 VDD2.n94 VDD2.n1 104.615
R2514 VDD2.n101 VDD2.n1 104.615
R2515 VDD2.n206 VDD2.n102 96.0748
R2516 VDD2.n206 VDD2.n205 52.7429
R2517 VDD2.n140 VDD2.t0 52.3082
R2518 VDD2.n35 VDD2.t1 52.3082
R2519 VDD2.n127 VDD2.n125 13.1884
R2520 VDD2.n55 VDD2.n22 13.1884
R2521 VDD2.n203 VDD2.n103 12.8005
R2522 VDD2.n163 VDD2.n162 12.8005
R2523 VDD2.n159 VDD2.n158 12.8005
R2524 VDD2.n56 VDD2.n24 12.8005
R2525 VDD2.n60 VDD2.n59 12.8005
R2526 VDD2.n100 VDD2.n0 12.8005
R2527 VDD2.n202 VDD2.n105 12.0247
R2528 VDD2.n166 VDD2.n123 12.0247
R2529 VDD2.n155 VDD2.n128 12.0247
R2530 VDD2.n51 VDD2.n50 12.0247
R2531 VDD2.n63 VDD2.n20 12.0247
R2532 VDD2.n99 VDD2.n2 12.0247
R2533 VDD2.n199 VDD2.n198 11.249
R2534 VDD2.n167 VDD2.n121 11.249
R2535 VDD2.n154 VDD2.n131 11.249
R2536 VDD2.n49 VDD2.n26 11.249
R2537 VDD2.n64 VDD2.n18 11.249
R2538 VDD2.n96 VDD2.n95 11.249
R2539 VDD2.n195 VDD2.n107 10.4732
R2540 VDD2.n171 VDD2.n170 10.4732
R2541 VDD2.n151 VDD2.n150 10.4732
R2542 VDD2.n46 VDD2.n45 10.4732
R2543 VDD2.n68 VDD2.n67 10.4732
R2544 VDD2.n92 VDD2.n4 10.4732
R2545 VDD2.n139 VDD2.n138 10.2747
R2546 VDD2.n34 VDD2.n33 10.2747
R2547 VDD2.n194 VDD2.n109 9.69747
R2548 VDD2.n174 VDD2.n119 9.69747
R2549 VDD2.n147 VDD2.n133 9.69747
R2550 VDD2.n42 VDD2.n28 9.69747
R2551 VDD2.n71 VDD2.n16 9.69747
R2552 VDD2.n91 VDD2.n6 9.69747
R2553 VDD2.n201 VDD2.n103 9.45567
R2554 VDD2.n98 VDD2.n0 9.45567
R2555 VDD2.n202 VDD2.n201 9.3005
R2556 VDD2.n200 VDD2.n199 9.3005
R2557 VDD2.n107 VDD2.n106 9.3005
R2558 VDD2.n194 VDD2.n193 9.3005
R2559 VDD2.n192 VDD2.n191 9.3005
R2560 VDD2.n111 VDD2.n110 9.3005
R2561 VDD2.n186 VDD2.n185 9.3005
R2562 VDD2.n184 VDD2.n183 9.3005
R2563 VDD2.n115 VDD2.n114 9.3005
R2564 VDD2.n178 VDD2.n177 9.3005
R2565 VDD2.n176 VDD2.n175 9.3005
R2566 VDD2.n119 VDD2.n118 9.3005
R2567 VDD2.n170 VDD2.n169 9.3005
R2568 VDD2.n168 VDD2.n167 9.3005
R2569 VDD2.n123 VDD2.n122 9.3005
R2570 VDD2.n162 VDD2.n161 9.3005
R2571 VDD2.n160 VDD2.n159 9.3005
R2572 VDD2.n128 VDD2.n126 9.3005
R2573 VDD2.n154 VDD2.n153 9.3005
R2574 VDD2.n152 VDD2.n151 9.3005
R2575 VDD2.n133 VDD2.n132 9.3005
R2576 VDD2.n146 VDD2.n145 9.3005
R2577 VDD2.n144 VDD2.n143 9.3005
R2578 VDD2.n137 VDD2.n136 9.3005
R2579 VDD2.n81 VDD2.n80 9.3005
R2580 VDD2.n83 VDD2.n82 9.3005
R2581 VDD2.n8 VDD2.n7 9.3005
R2582 VDD2.n89 VDD2.n88 9.3005
R2583 VDD2.n91 VDD2.n90 9.3005
R2584 VDD2.n4 VDD2.n3 9.3005
R2585 VDD2.n97 VDD2.n96 9.3005
R2586 VDD2.n99 VDD2.n98 9.3005
R2587 VDD2.n75 VDD2.n74 9.3005
R2588 VDD2.n73 VDD2.n72 9.3005
R2589 VDD2.n16 VDD2.n15 9.3005
R2590 VDD2.n67 VDD2.n66 9.3005
R2591 VDD2.n65 VDD2.n64 9.3005
R2592 VDD2.n20 VDD2.n19 9.3005
R2593 VDD2.n59 VDD2.n58 9.3005
R2594 VDD2.n32 VDD2.n31 9.3005
R2595 VDD2.n39 VDD2.n38 9.3005
R2596 VDD2.n41 VDD2.n40 9.3005
R2597 VDD2.n28 VDD2.n27 9.3005
R2598 VDD2.n47 VDD2.n46 9.3005
R2599 VDD2.n49 VDD2.n48 9.3005
R2600 VDD2.n50 VDD2.n23 9.3005
R2601 VDD2.n57 VDD2.n56 9.3005
R2602 VDD2.n12 VDD2.n11 9.3005
R2603 VDD2.n191 VDD2.n190 8.92171
R2604 VDD2.n175 VDD2.n117 8.92171
R2605 VDD2.n146 VDD2.n135 8.92171
R2606 VDD2.n41 VDD2.n30 8.92171
R2607 VDD2.n72 VDD2.n14 8.92171
R2608 VDD2.n88 VDD2.n87 8.92171
R2609 VDD2.n187 VDD2.n111 8.14595
R2610 VDD2.n179 VDD2.n178 8.14595
R2611 VDD2.n143 VDD2.n142 8.14595
R2612 VDD2.n38 VDD2.n37 8.14595
R2613 VDD2.n76 VDD2.n75 8.14595
R2614 VDD2.n84 VDD2.n8 8.14595
R2615 VDD2.n186 VDD2.n113 7.3702
R2616 VDD2.n182 VDD2.n115 7.3702
R2617 VDD2.n139 VDD2.n137 7.3702
R2618 VDD2.n34 VDD2.n32 7.3702
R2619 VDD2.n79 VDD2.n12 7.3702
R2620 VDD2.n83 VDD2.n10 7.3702
R2621 VDD2.n183 VDD2.n113 6.59444
R2622 VDD2.n183 VDD2.n182 6.59444
R2623 VDD2.n80 VDD2.n79 6.59444
R2624 VDD2.n80 VDD2.n10 6.59444
R2625 VDD2.n187 VDD2.n186 5.81868
R2626 VDD2.n179 VDD2.n115 5.81868
R2627 VDD2.n142 VDD2.n137 5.81868
R2628 VDD2.n37 VDD2.n32 5.81868
R2629 VDD2.n76 VDD2.n12 5.81868
R2630 VDD2.n84 VDD2.n83 5.81868
R2631 VDD2.n190 VDD2.n111 5.04292
R2632 VDD2.n178 VDD2.n117 5.04292
R2633 VDD2.n143 VDD2.n135 5.04292
R2634 VDD2.n38 VDD2.n30 5.04292
R2635 VDD2.n75 VDD2.n14 5.04292
R2636 VDD2.n87 VDD2.n8 5.04292
R2637 VDD2.n191 VDD2.n109 4.26717
R2638 VDD2.n175 VDD2.n174 4.26717
R2639 VDD2.n147 VDD2.n146 4.26717
R2640 VDD2.n42 VDD2.n41 4.26717
R2641 VDD2.n72 VDD2.n71 4.26717
R2642 VDD2.n88 VDD2.n6 4.26717
R2643 VDD2.n195 VDD2.n194 3.49141
R2644 VDD2.n171 VDD2.n119 3.49141
R2645 VDD2.n150 VDD2.n133 3.49141
R2646 VDD2.n45 VDD2.n28 3.49141
R2647 VDD2.n68 VDD2.n16 3.49141
R2648 VDD2.n92 VDD2.n91 3.49141
R2649 VDD2.n33 VDD2.n31 2.84303
R2650 VDD2.n138 VDD2.n136 2.84303
R2651 VDD2.n198 VDD2.n107 2.71565
R2652 VDD2.n170 VDD2.n121 2.71565
R2653 VDD2.n151 VDD2.n131 2.71565
R2654 VDD2.n46 VDD2.n26 2.71565
R2655 VDD2.n67 VDD2.n18 2.71565
R2656 VDD2.n95 VDD2.n4 2.71565
R2657 VDD2.n199 VDD2.n105 1.93989
R2658 VDD2.n167 VDD2.n166 1.93989
R2659 VDD2.n155 VDD2.n154 1.93989
R2660 VDD2.n51 VDD2.n49 1.93989
R2661 VDD2.n64 VDD2.n63 1.93989
R2662 VDD2.n96 VDD2.n2 1.93989
R2663 VDD2.n203 VDD2.n202 1.16414
R2664 VDD2.n163 VDD2.n123 1.16414
R2665 VDD2.n158 VDD2.n128 1.16414
R2666 VDD2.n50 VDD2.n24 1.16414
R2667 VDD2.n60 VDD2.n20 1.16414
R2668 VDD2.n100 VDD2.n99 1.16414
R2669 VDD2 VDD2.n206 0.489724
R2670 VDD2.n205 VDD2.n103 0.388379
R2671 VDD2.n162 VDD2.n125 0.388379
R2672 VDD2.n159 VDD2.n127 0.388379
R2673 VDD2.n56 VDD2.n55 0.388379
R2674 VDD2.n59 VDD2.n22 0.388379
R2675 VDD2.n102 VDD2.n0 0.388379
R2676 VDD2.n201 VDD2.n200 0.155672
R2677 VDD2.n200 VDD2.n106 0.155672
R2678 VDD2.n193 VDD2.n106 0.155672
R2679 VDD2.n193 VDD2.n192 0.155672
R2680 VDD2.n192 VDD2.n110 0.155672
R2681 VDD2.n185 VDD2.n110 0.155672
R2682 VDD2.n185 VDD2.n184 0.155672
R2683 VDD2.n184 VDD2.n114 0.155672
R2684 VDD2.n177 VDD2.n114 0.155672
R2685 VDD2.n177 VDD2.n176 0.155672
R2686 VDD2.n176 VDD2.n118 0.155672
R2687 VDD2.n169 VDD2.n118 0.155672
R2688 VDD2.n169 VDD2.n168 0.155672
R2689 VDD2.n168 VDD2.n122 0.155672
R2690 VDD2.n161 VDD2.n122 0.155672
R2691 VDD2.n161 VDD2.n160 0.155672
R2692 VDD2.n160 VDD2.n126 0.155672
R2693 VDD2.n153 VDD2.n126 0.155672
R2694 VDD2.n153 VDD2.n152 0.155672
R2695 VDD2.n152 VDD2.n132 0.155672
R2696 VDD2.n145 VDD2.n132 0.155672
R2697 VDD2.n145 VDD2.n144 0.155672
R2698 VDD2.n144 VDD2.n136 0.155672
R2699 VDD2.n39 VDD2.n31 0.155672
R2700 VDD2.n40 VDD2.n39 0.155672
R2701 VDD2.n40 VDD2.n27 0.155672
R2702 VDD2.n47 VDD2.n27 0.155672
R2703 VDD2.n48 VDD2.n47 0.155672
R2704 VDD2.n48 VDD2.n23 0.155672
R2705 VDD2.n57 VDD2.n23 0.155672
R2706 VDD2.n58 VDD2.n57 0.155672
R2707 VDD2.n58 VDD2.n19 0.155672
R2708 VDD2.n65 VDD2.n19 0.155672
R2709 VDD2.n66 VDD2.n65 0.155672
R2710 VDD2.n66 VDD2.n15 0.155672
R2711 VDD2.n73 VDD2.n15 0.155672
R2712 VDD2.n74 VDD2.n73 0.155672
R2713 VDD2.n74 VDD2.n11 0.155672
R2714 VDD2.n81 VDD2.n11 0.155672
R2715 VDD2.n82 VDD2.n81 0.155672
R2716 VDD2.n82 VDD2.n7 0.155672
R2717 VDD2.n89 VDD2.n7 0.155672
R2718 VDD2.n90 VDD2.n89 0.155672
R2719 VDD2.n90 VDD2.n3 0.155672
R2720 VDD2.n97 VDD2.n3 0.155672
R2721 VDD2.n98 VDD2.n97 0.155672
C0 VP VDD1 4.02068f
C1 VP VDD2 0.295158f
C2 VN VDD1 0.148029f
C3 VTAIL VDD1 7.00856f
C4 VN VDD2 3.87833f
C5 VTAIL VDD2 7.04928f
C6 VP VN 6.28262f
C7 VP VTAIL 3.20084f
C8 VDD1 VDD2 0.56651f
C9 VN VTAIL 3.18629f
C10 VDD2 B 5.33035f
C11 VDD1 B 8.4233f
C12 VTAIL B 9.575613f
C13 VN B 11.661099f
C14 VP B 5.71516f
C15 VDD2.n0 B 0.011222f
C16 VDD2.n1 B 0.025261f
C17 VDD2.n2 B 0.011316f
C18 VDD2.n3 B 0.019889f
C19 VDD2.n4 B 0.010687f
C20 VDD2.n5 B 0.025261f
C21 VDD2.n6 B 0.011316f
C22 VDD2.n7 B 0.019889f
C23 VDD2.n8 B 0.010687f
C24 VDD2.n9 B 0.025261f
C25 VDD2.n10 B 0.011316f
C26 VDD2.n11 B 0.019889f
C27 VDD2.n12 B 0.010687f
C28 VDD2.n13 B 0.025261f
C29 VDD2.n14 B 0.011316f
C30 VDD2.n15 B 0.019889f
C31 VDD2.n16 B 0.010687f
C32 VDD2.n17 B 0.025261f
C33 VDD2.n18 B 0.011316f
C34 VDD2.n19 B 0.019889f
C35 VDD2.n20 B 0.010687f
C36 VDD2.n21 B 0.025261f
C37 VDD2.n22 B 0.011002f
C38 VDD2.n23 B 0.019889f
C39 VDD2.n24 B 0.011316f
C40 VDD2.n25 B 0.025261f
C41 VDD2.n26 B 0.011316f
C42 VDD2.n27 B 0.019889f
C43 VDD2.n28 B 0.010687f
C44 VDD2.n29 B 0.025261f
C45 VDD2.n30 B 0.011316f
C46 VDD2.n31 B 1.60665f
C47 VDD2.n32 B 0.010687f
C48 VDD2.t1 B 0.043394f
C49 VDD2.n33 B 0.195468f
C50 VDD2.n34 B 0.017857f
C51 VDD2.n35 B 0.018946f
C52 VDD2.n36 B 0.025261f
C53 VDD2.n37 B 0.011316f
C54 VDD2.n38 B 0.010687f
C55 VDD2.n39 B 0.019889f
C56 VDD2.n40 B 0.019889f
C57 VDD2.n41 B 0.010687f
C58 VDD2.n42 B 0.011316f
C59 VDD2.n43 B 0.025261f
C60 VDD2.n44 B 0.025261f
C61 VDD2.n45 B 0.011316f
C62 VDD2.n46 B 0.010687f
C63 VDD2.n47 B 0.019889f
C64 VDD2.n48 B 0.019889f
C65 VDD2.n49 B 0.010687f
C66 VDD2.n50 B 0.010687f
C67 VDD2.n51 B 0.011316f
C68 VDD2.n52 B 0.025261f
C69 VDD2.n53 B 0.025261f
C70 VDD2.n54 B 0.025261f
C71 VDD2.n55 B 0.011002f
C72 VDD2.n56 B 0.010687f
C73 VDD2.n57 B 0.019889f
C74 VDD2.n58 B 0.019889f
C75 VDD2.n59 B 0.010687f
C76 VDD2.n60 B 0.011316f
C77 VDD2.n61 B 0.025261f
C78 VDD2.n62 B 0.025261f
C79 VDD2.n63 B 0.011316f
C80 VDD2.n64 B 0.010687f
C81 VDD2.n65 B 0.019889f
C82 VDD2.n66 B 0.019889f
C83 VDD2.n67 B 0.010687f
C84 VDD2.n68 B 0.011316f
C85 VDD2.n69 B 0.025261f
C86 VDD2.n70 B 0.025261f
C87 VDD2.n71 B 0.011316f
C88 VDD2.n72 B 0.010687f
C89 VDD2.n73 B 0.019889f
C90 VDD2.n74 B 0.019889f
C91 VDD2.n75 B 0.010687f
C92 VDD2.n76 B 0.011316f
C93 VDD2.n77 B 0.025261f
C94 VDD2.n78 B 0.025261f
C95 VDD2.n79 B 0.011316f
C96 VDD2.n80 B 0.010687f
C97 VDD2.n81 B 0.019889f
C98 VDD2.n82 B 0.019889f
C99 VDD2.n83 B 0.010687f
C100 VDD2.n84 B 0.011316f
C101 VDD2.n85 B 0.025261f
C102 VDD2.n86 B 0.025261f
C103 VDD2.n87 B 0.011316f
C104 VDD2.n88 B 0.010687f
C105 VDD2.n89 B 0.019889f
C106 VDD2.n90 B 0.019889f
C107 VDD2.n91 B 0.010687f
C108 VDD2.n92 B 0.011316f
C109 VDD2.n93 B 0.025261f
C110 VDD2.n94 B 0.025261f
C111 VDD2.n95 B 0.011316f
C112 VDD2.n96 B 0.010687f
C113 VDD2.n97 B 0.019889f
C114 VDD2.n98 B 0.051949f
C115 VDD2.n99 B 0.010687f
C116 VDD2.n100 B 0.011316f
C117 VDD2.n101 B 0.052312f
C118 VDD2.n102 B 0.723019f
C119 VDD2.n103 B 0.011222f
C120 VDD2.n104 B 0.025261f
C121 VDD2.n105 B 0.011316f
C122 VDD2.n106 B 0.019889f
C123 VDD2.n107 B 0.010687f
C124 VDD2.n108 B 0.025261f
C125 VDD2.n109 B 0.011316f
C126 VDD2.n110 B 0.019889f
C127 VDD2.n111 B 0.010687f
C128 VDD2.n112 B 0.025261f
C129 VDD2.n113 B 0.011316f
C130 VDD2.n114 B 0.019889f
C131 VDD2.n115 B 0.010687f
C132 VDD2.n116 B 0.025261f
C133 VDD2.n117 B 0.011316f
C134 VDD2.n118 B 0.019889f
C135 VDD2.n119 B 0.010687f
C136 VDD2.n120 B 0.025261f
C137 VDD2.n121 B 0.011316f
C138 VDD2.n122 B 0.019889f
C139 VDD2.n123 B 0.010687f
C140 VDD2.n124 B 0.025261f
C141 VDD2.n125 B 0.011002f
C142 VDD2.n126 B 0.019889f
C143 VDD2.n127 B 0.011002f
C144 VDD2.n128 B 0.010687f
C145 VDD2.n129 B 0.025261f
C146 VDD2.n130 B 0.025261f
C147 VDD2.n131 B 0.011316f
C148 VDD2.n132 B 0.019889f
C149 VDD2.n133 B 0.010687f
C150 VDD2.n134 B 0.025261f
C151 VDD2.n135 B 0.011316f
C152 VDD2.n136 B 1.60665f
C153 VDD2.n137 B 0.010687f
C154 VDD2.t0 B 0.043394f
C155 VDD2.n138 B 0.195468f
C156 VDD2.n139 B 0.017857f
C157 VDD2.n140 B 0.018946f
C158 VDD2.n141 B 0.025261f
C159 VDD2.n142 B 0.011316f
C160 VDD2.n143 B 0.010687f
C161 VDD2.n144 B 0.019889f
C162 VDD2.n145 B 0.019889f
C163 VDD2.n146 B 0.010687f
C164 VDD2.n147 B 0.011316f
C165 VDD2.n148 B 0.025261f
C166 VDD2.n149 B 0.025261f
C167 VDD2.n150 B 0.011316f
C168 VDD2.n151 B 0.010687f
C169 VDD2.n152 B 0.019889f
C170 VDD2.n153 B 0.019889f
C171 VDD2.n154 B 0.010687f
C172 VDD2.n155 B 0.011316f
C173 VDD2.n156 B 0.025261f
C174 VDD2.n157 B 0.025261f
C175 VDD2.n158 B 0.011316f
C176 VDD2.n159 B 0.010687f
C177 VDD2.n160 B 0.019889f
C178 VDD2.n161 B 0.019889f
C179 VDD2.n162 B 0.010687f
C180 VDD2.n163 B 0.011316f
C181 VDD2.n164 B 0.025261f
C182 VDD2.n165 B 0.025261f
C183 VDD2.n166 B 0.011316f
C184 VDD2.n167 B 0.010687f
C185 VDD2.n168 B 0.019889f
C186 VDD2.n169 B 0.019889f
C187 VDD2.n170 B 0.010687f
C188 VDD2.n171 B 0.011316f
C189 VDD2.n172 B 0.025261f
C190 VDD2.n173 B 0.025261f
C191 VDD2.n174 B 0.011316f
C192 VDD2.n175 B 0.010687f
C193 VDD2.n176 B 0.019889f
C194 VDD2.n177 B 0.019889f
C195 VDD2.n178 B 0.010687f
C196 VDD2.n179 B 0.011316f
C197 VDD2.n180 B 0.025261f
C198 VDD2.n181 B 0.025261f
C199 VDD2.n182 B 0.011316f
C200 VDD2.n183 B 0.010687f
C201 VDD2.n184 B 0.019889f
C202 VDD2.n185 B 0.019889f
C203 VDD2.n186 B 0.010687f
C204 VDD2.n187 B 0.011316f
C205 VDD2.n188 B 0.025261f
C206 VDD2.n189 B 0.025261f
C207 VDD2.n190 B 0.011316f
C208 VDD2.n191 B 0.010687f
C209 VDD2.n192 B 0.019889f
C210 VDD2.n193 B 0.019889f
C211 VDD2.n194 B 0.010687f
C212 VDD2.n195 B 0.011316f
C213 VDD2.n196 B 0.025261f
C214 VDD2.n197 B 0.025261f
C215 VDD2.n198 B 0.011316f
C216 VDD2.n199 B 0.010687f
C217 VDD2.n200 B 0.019889f
C218 VDD2.n201 B 0.051949f
C219 VDD2.n202 B 0.010687f
C220 VDD2.n203 B 0.011316f
C221 VDD2.n204 B 0.052312f
C222 VDD2.n205 B 0.057967f
C223 VDD2.n206 B 2.87114f
C224 VN.t0 B 3.55842f
C225 VN.t1 B 3.94973f
C226 VDD1.n0 B 0.011249f
C227 VDD1.n1 B 0.025322f
C228 VDD1.n2 B 0.011343f
C229 VDD1.n3 B 0.019937f
C230 VDD1.n4 B 0.010713f
C231 VDD1.n5 B 0.025322f
C232 VDD1.n6 B 0.011343f
C233 VDD1.n7 B 0.019937f
C234 VDD1.n8 B 0.010713f
C235 VDD1.n9 B 0.025322f
C236 VDD1.n10 B 0.011343f
C237 VDD1.n11 B 0.019937f
C238 VDD1.n12 B 0.010713f
C239 VDD1.n13 B 0.025322f
C240 VDD1.n14 B 0.011343f
C241 VDD1.n15 B 0.019937f
C242 VDD1.n16 B 0.010713f
C243 VDD1.n17 B 0.025322f
C244 VDD1.n18 B 0.011343f
C245 VDD1.n19 B 0.019937f
C246 VDD1.n20 B 0.010713f
C247 VDD1.n21 B 0.025322f
C248 VDD1.n22 B 0.011028f
C249 VDD1.n23 B 0.019937f
C250 VDD1.n24 B 0.011028f
C251 VDD1.n25 B 0.010713f
C252 VDD1.n26 B 0.025322f
C253 VDD1.n27 B 0.025322f
C254 VDD1.n28 B 0.011343f
C255 VDD1.n29 B 0.019937f
C256 VDD1.n30 B 0.010713f
C257 VDD1.n31 B 0.025322f
C258 VDD1.n32 B 0.011343f
C259 VDD1.n33 B 1.61053f
C260 VDD1.n34 B 0.010713f
C261 VDD1.t0 B 0.043499f
C262 VDD1.n35 B 0.195941f
C263 VDD1.n36 B 0.017901f
C264 VDD1.n37 B 0.018991f
C265 VDD1.n38 B 0.025322f
C266 VDD1.n39 B 0.011343f
C267 VDD1.n40 B 0.010713f
C268 VDD1.n41 B 0.019937f
C269 VDD1.n42 B 0.019937f
C270 VDD1.n43 B 0.010713f
C271 VDD1.n44 B 0.011343f
C272 VDD1.n45 B 0.025322f
C273 VDD1.n46 B 0.025322f
C274 VDD1.n47 B 0.011343f
C275 VDD1.n48 B 0.010713f
C276 VDD1.n49 B 0.019937f
C277 VDD1.n50 B 0.019937f
C278 VDD1.n51 B 0.010713f
C279 VDD1.n52 B 0.011343f
C280 VDD1.n53 B 0.025322f
C281 VDD1.n54 B 0.025322f
C282 VDD1.n55 B 0.011343f
C283 VDD1.n56 B 0.010713f
C284 VDD1.n57 B 0.019937f
C285 VDD1.n58 B 0.019937f
C286 VDD1.n59 B 0.010713f
C287 VDD1.n60 B 0.011343f
C288 VDD1.n61 B 0.025322f
C289 VDD1.n62 B 0.025322f
C290 VDD1.n63 B 0.011343f
C291 VDD1.n64 B 0.010713f
C292 VDD1.n65 B 0.019937f
C293 VDD1.n66 B 0.019937f
C294 VDD1.n67 B 0.010713f
C295 VDD1.n68 B 0.011343f
C296 VDD1.n69 B 0.025322f
C297 VDD1.n70 B 0.025322f
C298 VDD1.n71 B 0.011343f
C299 VDD1.n72 B 0.010713f
C300 VDD1.n73 B 0.019937f
C301 VDD1.n74 B 0.019937f
C302 VDD1.n75 B 0.010713f
C303 VDD1.n76 B 0.011343f
C304 VDD1.n77 B 0.025322f
C305 VDD1.n78 B 0.025322f
C306 VDD1.n79 B 0.011343f
C307 VDD1.n80 B 0.010713f
C308 VDD1.n81 B 0.019937f
C309 VDD1.n82 B 0.019937f
C310 VDD1.n83 B 0.010713f
C311 VDD1.n84 B 0.011343f
C312 VDD1.n85 B 0.025322f
C313 VDD1.n86 B 0.025322f
C314 VDD1.n87 B 0.011343f
C315 VDD1.n88 B 0.010713f
C316 VDD1.n89 B 0.019937f
C317 VDD1.n90 B 0.019937f
C318 VDD1.n91 B 0.010713f
C319 VDD1.n92 B 0.011343f
C320 VDD1.n93 B 0.025322f
C321 VDD1.n94 B 0.025322f
C322 VDD1.n95 B 0.011343f
C323 VDD1.n96 B 0.010713f
C324 VDD1.n97 B 0.019937f
C325 VDD1.n98 B 0.052074f
C326 VDD1.n99 B 0.010713f
C327 VDD1.n100 B 0.011343f
C328 VDD1.n101 B 0.052439f
C329 VDD1.n102 B 0.058777f
C330 VDD1.n103 B 0.011249f
C331 VDD1.n104 B 0.025322f
C332 VDD1.n105 B 0.011343f
C333 VDD1.n106 B 0.019937f
C334 VDD1.n107 B 0.010713f
C335 VDD1.n108 B 0.025322f
C336 VDD1.n109 B 0.011343f
C337 VDD1.n110 B 0.019937f
C338 VDD1.n111 B 0.010713f
C339 VDD1.n112 B 0.025322f
C340 VDD1.n113 B 0.011343f
C341 VDD1.n114 B 0.019937f
C342 VDD1.n115 B 0.010713f
C343 VDD1.n116 B 0.025322f
C344 VDD1.n117 B 0.011343f
C345 VDD1.n118 B 0.019937f
C346 VDD1.n119 B 0.010713f
C347 VDD1.n120 B 0.025322f
C348 VDD1.n121 B 0.011343f
C349 VDD1.n122 B 0.019937f
C350 VDD1.n123 B 0.010713f
C351 VDD1.n124 B 0.025322f
C352 VDD1.n125 B 0.011028f
C353 VDD1.n126 B 0.019937f
C354 VDD1.n127 B 0.011343f
C355 VDD1.n128 B 0.025322f
C356 VDD1.n129 B 0.011343f
C357 VDD1.n130 B 0.019937f
C358 VDD1.n131 B 0.010713f
C359 VDD1.n132 B 0.025322f
C360 VDD1.n133 B 0.011343f
C361 VDD1.n134 B 1.61053f
C362 VDD1.n135 B 0.010713f
C363 VDD1.t1 B 0.043499f
C364 VDD1.n136 B 0.195941f
C365 VDD1.n137 B 0.017901f
C366 VDD1.n138 B 0.018991f
C367 VDD1.n139 B 0.025322f
C368 VDD1.n140 B 0.011343f
C369 VDD1.n141 B 0.010713f
C370 VDD1.n142 B 0.019937f
C371 VDD1.n143 B 0.019937f
C372 VDD1.n144 B 0.010713f
C373 VDD1.n145 B 0.011343f
C374 VDD1.n146 B 0.025322f
C375 VDD1.n147 B 0.025322f
C376 VDD1.n148 B 0.011343f
C377 VDD1.n149 B 0.010713f
C378 VDD1.n150 B 0.019937f
C379 VDD1.n151 B 0.019937f
C380 VDD1.n152 B 0.010713f
C381 VDD1.n153 B 0.010713f
C382 VDD1.n154 B 0.011343f
C383 VDD1.n155 B 0.025322f
C384 VDD1.n156 B 0.025322f
C385 VDD1.n157 B 0.025322f
C386 VDD1.n158 B 0.011028f
C387 VDD1.n159 B 0.010713f
C388 VDD1.n160 B 0.019937f
C389 VDD1.n161 B 0.019937f
C390 VDD1.n162 B 0.010713f
C391 VDD1.n163 B 0.011343f
C392 VDD1.n164 B 0.025322f
C393 VDD1.n165 B 0.025322f
C394 VDD1.n166 B 0.011343f
C395 VDD1.n167 B 0.010713f
C396 VDD1.n168 B 0.019937f
C397 VDD1.n169 B 0.019937f
C398 VDD1.n170 B 0.010713f
C399 VDD1.n171 B 0.011343f
C400 VDD1.n172 B 0.025322f
C401 VDD1.n173 B 0.025322f
C402 VDD1.n174 B 0.011343f
C403 VDD1.n175 B 0.010713f
C404 VDD1.n176 B 0.019937f
C405 VDD1.n177 B 0.019937f
C406 VDD1.n178 B 0.010713f
C407 VDD1.n179 B 0.011343f
C408 VDD1.n180 B 0.025322f
C409 VDD1.n181 B 0.025322f
C410 VDD1.n182 B 0.011343f
C411 VDD1.n183 B 0.010713f
C412 VDD1.n184 B 0.019937f
C413 VDD1.n185 B 0.019937f
C414 VDD1.n186 B 0.010713f
C415 VDD1.n187 B 0.011343f
C416 VDD1.n188 B 0.025322f
C417 VDD1.n189 B 0.025322f
C418 VDD1.n190 B 0.011343f
C419 VDD1.n191 B 0.010713f
C420 VDD1.n192 B 0.019937f
C421 VDD1.n193 B 0.019937f
C422 VDD1.n194 B 0.010713f
C423 VDD1.n195 B 0.011343f
C424 VDD1.n196 B 0.025322f
C425 VDD1.n197 B 0.025322f
C426 VDD1.n198 B 0.011343f
C427 VDD1.n199 B 0.010713f
C428 VDD1.n200 B 0.019937f
C429 VDD1.n201 B 0.052074f
C430 VDD1.n202 B 0.010713f
C431 VDD1.n203 B 0.011343f
C432 VDD1.n204 B 0.052439f
C433 VDD1.n205 B 0.759939f
C434 VTAIL.n0 B 0.010994f
C435 VTAIL.n1 B 0.024748f
C436 VTAIL.n2 B 0.011086f
C437 VTAIL.n3 B 0.019485f
C438 VTAIL.n4 B 0.01047f
C439 VTAIL.n5 B 0.024748f
C440 VTAIL.n6 B 0.011086f
C441 VTAIL.n7 B 0.019485f
C442 VTAIL.n8 B 0.01047f
C443 VTAIL.n9 B 0.024748f
C444 VTAIL.n10 B 0.011086f
C445 VTAIL.n11 B 0.019485f
C446 VTAIL.n12 B 0.01047f
C447 VTAIL.n13 B 0.024748f
C448 VTAIL.n14 B 0.011086f
C449 VTAIL.n15 B 0.019485f
C450 VTAIL.n16 B 0.01047f
C451 VTAIL.n17 B 0.024748f
C452 VTAIL.n18 B 0.011086f
C453 VTAIL.n19 B 0.019485f
C454 VTAIL.n20 B 0.01047f
C455 VTAIL.n21 B 0.024748f
C456 VTAIL.n22 B 0.010778f
C457 VTAIL.n23 B 0.019485f
C458 VTAIL.n24 B 0.011086f
C459 VTAIL.n25 B 0.024748f
C460 VTAIL.n26 B 0.011086f
C461 VTAIL.n27 B 0.019485f
C462 VTAIL.n28 B 0.01047f
C463 VTAIL.n29 B 0.024748f
C464 VTAIL.n30 B 0.011086f
C465 VTAIL.n31 B 1.57403f
C466 VTAIL.n32 B 0.01047f
C467 VTAIL.t3 B 0.042513f
C468 VTAIL.n33 B 0.1915f
C469 VTAIL.n34 B 0.017495f
C470 VTAIL.n35 B 0.018561f
C471 VTAIL.n36 B 0.024748f
C472 VTAIL.n37 B 0.011086f
C473 VTAIL.n38 B 0.01047f
C474 VTAIL.n39 B 0.019485f
C475 VTAIL.n40 B 0.019485f
C476 VTAIL.n41 B 0.01047f
C477 VTAIL.n42 B 0.011086f
C478 VTAIL.n43 B 0.024748f
C479 VTAIL.n44 B 0.024748f
C480 VTAIL.n45 B 0.011086f
C481 VTAIL.n46 B 0.01047f
C482 VTAIL.n47 B 0.019485f
C483 VTAIL.n48 B 0.019485f
C484 VTAIL.n49 B 0.01047f
C485 VTAIL.n50 B 0.01047f
C486 VTAIL.n51 B 0.011086f
C487 VTAIL.n52 B 0.024748f
C488 VTAIL.n53 B 0.024748f
C489 VTAIL.n54 B 0.024748f
C490 VTAIL.n55 B 0.010778f
C491 VTAIL.n56 B 0.01047f
C492 VTAIL.n57 B 0.019485f
C493 VTAIL.n58 B 0.019485f
C494 VTAIL.n59 B 0.01047f
C495 VTAIL.n60 B 0.011086f
C496 VTAIL.n61 B 0.024748f
C497 VTAIL.n62 B 0.024748f
C498 VTAIL.n63 B 0.011086f
C499 VTAIL.n64 B 0.01047f
C500 VTAIL.n65 B 0.019485f
C501 VTAIL.n66 B 0.019485f
C502 VTAIL.n67 B 0.01047f
C503 VTAIL.n68 B 0.011086f
C504 VTAIL.n69 B 0.024748f
C505 VTAIL.n70 B 0.024748f
C506 VTAIL.n71 B 0.011086f
C507 VTAIL.n72 B 0.01047f
C508 VTAIL.n73 B 0.019485f
C509 VTAIL.n74 B 0.019485f
C510 VTAIL.n75 B 0.01047f
C511 VTAIL.n76 B 0.011086f
C512 VTAIL.n77 B 0.024748f
C513 VTAIL.n78 B 0.024748f
C514 VTAIL.n79 B 0.011086f
C515 VTAIL.n80 B 0.01047f
C516 VTAIL.n81 B 0.019485f
C517 VTAIL.n82 B 0.019485f
C518 VTAIL.n83 B 0.01047f
C519 VTAIL.n84 B 0.011086f
C520 VTAIL.n85 B 0.024748f
C521 VTAIL.n86 B 0.024748f
C522 VTAIL.n87 B 0.011086f
C523 VTAIL.n88 B 0.01047f
C524 VTAIL.n89 B 0.019485f
C525 VTAIL.n90 B 0.019485f
C526 VTAIL.n91 B 0.01047f
C527 VTAIL.n92 B 0.011086f
C528 VTAIL.n93 B 0.024748f
C529 VTAIL.n94 B 0.024748f
C530 VTAIL.n95 B 0.011086f
C531 VTAIL.n96 B 0.01047f
C532 VTAIL.n97 B 0.019485f
C533 VTAIL.n98 B 0.050894f
C534 VTAIL.n99 B 0.01047f
C535 VTAIL.n100 B 0.011086f
C536 VTAIL.n101 B 0.05125f
C537 VTAIL.n102 B 0.043373f
C538 VTAIL.n103 B 1.57966f
C539 VTAIL.n104 B 0.010994f
C540 VTAIL.n105 B 0.024748f
C541 VTAIL.n106 B 0.011086f
C542 VTAIL.n107 B 0.019485f
C543 VTAIL.n108 B 0.01047f
C544 VTAIL.n109 B 0.024748f
C545 VTAIL.n110 B 0.011086f
C546 VTAIL.n111 B 0.019485f
C547 VTAIL.n112 B 0.01047f
C548 VTAIL.n113 B 0.024748f
C549 VTAIL.n114 B 0.011086f
C550 VTAIL.n115 B 0.019485f
C551 VTAIL.n116 B 0.01047f
C552 VTAIL.n117 B 0.024748f
C553 VTAIL.n118 B 0.011086f
C554 VTAIL.n119 B 0.019485f
C555 VTAIL.n120 B 0.01047f
C556 VTAIL.n121 B 0.024748f
C557 VTAIL.n122 B 0.011086f
C558 VTAIL.n123 B 0.019485f
C559 VTAIL.n124 B 0.01047f
C560 VTAIL.n125 B 0.024748f
C561 VTAIL.n126 B 0.010778f
C562 VTAIL.n127 B 0.019485f
C563 VTAIL.n128 B 0.010778f
C564 VTAIL.n129 B 0.01047f
C565 VTAIL.n130 B 0.024748f
C566 VTAIL.n131 B 0.024748f
C567 VTAIL.n132 B 0.011086f
C568 VTAIL.n133 B 0.019485f
C569 VTAIL.n134 B 0.01047f
C570 VTAIL.n135 B 0.024748f
C571 VTAIL.n136 B 0.011086f
C572 VTAIL.n137 B 1.57403f
C573 VTAIL.n138 B 0.01047f
C574 VTAIL.t0 B 0.042513f
C575 VTAIL.n139 B 0.1915f
C576 VTAIL.n140 B 0.017495f
C577 VTAIL.n141 B 0.018561f
C578 VTAIL.n142 B 0.024748f
C579 VTAIL.n143 B 0.011086f
C580 VTAIL.n144 B 0.01047f
C581 VTAIL.n145 B 0.019485f
C582 VTAIL.n146 B 0.019485f
C583 VTAIL.n147 B 0.01047f
C584 VTAIL.n148 B 0.011086f
C585 VTAIL.n149 B 0.024748f
C586 VTAIL.n150 B 0.024748f
C587 VTAIL.n151 B 0.011086f
C588 VTAIL.n152 B 0.01047f
C589 VTAIL.n153 B 0.019485f
C590 VTAIL.n154 B 0.019485f
C591 VTAIL.n155 B 0.01047f
C592 VTAIL.n156 B 0.011086f
C593 VTAIL.n157 B 0.024748f
C594 VTAIL.n158 B 0.024748f
C595 VTAIL.n159 B 0.011086f
C596 VTAIL.n160 B 0.01047f
C597 VTAIL.n161 B 0.019485f
C598 VTAIL.n162 B 0.019485f
C599 VTAIL.n163 B 0.01047f
C600 VTAIL.n164 B 0.011086f
C601 VTAIL.n165 B 0.024748f
C602 VTAIL.n166 B 0.024748f
C603 VTAIL.n167 B 0.011086f
C604 VTAIL.n168 B 0.01047f
C605 VTAIL.n169 B 0.019485f
C606 VTAIL.n170 B 0.019485f
C607 VTAIL.n171 B 0.01047f
C608 VTAIL.n172 B 0.011086f
C609 VTAIL.n173 B 0.024748f
C610 VTAIL.n174 B 0.024748f
C611 VTAIL.n175 B 0.011086f
C612 VTAIL.n176 B 0.01047f
C613 VTAIL.n177 B 0.019485f
C614 VTAIL.n178 B 0.019485f
C615 VTAIL.n179 B 0.01047f
C616 VTAIL.n180 B 0.011086f
C617 VTAIL.n181 B 0.024748f
C618 VTAIL.n182 B 0.024748f
C619 VTAIL.n183 B 0.011086f
C620 VTAIL.n184 B 0.01047f
C621 VTAIL.n185 B 0.019485f
C622 VTAIL.n186 B 0.019485f
C623 VTAIL.n187 B 0.01047f
C624 VTAIL.n188 B 0.011086f
C625 VTAIL.n189 B 0.024748f
C626 VTAIL.n190 B 0.024748f
C627 VTAIL.n191 B 0.011086f
C628 VTAIL.n192 B 0.01047f
C629 VTAIL.n193 B 0.019485f
C630 VTAIL.n194 B 0.019485f
C631 VTAIL.n195 B 0.01047f
C632 VTAIL.n196 B 0.011086f
C633 VTAIL.n197 B 0.024748f
C634 VTAIL.n198 B 0.024748f
C635 VTAIL.n199 B 0.011086f
C636 VTAIL.n200 B 0.01047f
C637 VTAIL.n201 B 0.019485f
C638 VTAIL.n202 B 0.050894f
C639 VTAIL.n203 B 0.01047f
C640 VTAIL.n204 B 0.011086f
C641 VTAIL.n205 B 0.05125f
C642 VTAIL.n206 B 0.043373f
C643 VTAIL.n207 B 1.60307f
C644 VTAIL.n208 B 0.010994f
C645 VTAIL.n209 B 0.024748f
C646 VTAIL.n210 B 0.011086f
C647 VTAIL.n211 B 0.019485f
C648 VTAIL.n212 B 0.01047f
C649 VTAIL.n213 B 0.024748f
C650 VTAIL.n214 B 0.011086f
C651 VTAIL.n215 B 0.019485f
C652 VTAIL.n216 B 0.01047f
C653 VTAIL.n217 B 0.024748f
C654 VTAIL.n218 B 0.011086f
C655 VTAIL.n219 B 0.019485f
C656 VTAIL.n220 B 0.01047f
C657 VTAIL.n221 B 0.024748f
C658 VTAIL.n222 B 0.011086f
C659 VTAIL.n223 B 0.019485f
C660 VTAIL.n224 B 0.01047f
C661 VTAIL.n225 B 0.024748f
C662 VTAIL.n226 B 0.011086f
C663 VTAIL.n227 B 0.019485f
C664 VTAIL.n228 B 0.01047f
C665 VTAIL.n229 B 0.024748f
C666 VTAIL.n230 B 0.010778f
C667 VTAIL.n231 B 0.019485f
C668 VTAIL.n232 B 0.010778f
C669 VTAIL.n233 B 0.01047f
C670 VTAIL.n234 B 0.024748f
C671 VTAIL.n235 B 0.024748f
C672 VTAIL.n236 B 0.011086f
C673 VTAIL.n237 B 0.019485f
C674 VTAIL.n238 B 0.01047f
C675 VTAIL.n239 B 0.024748f
C676 VTAIL.n240 B 0.011086f
C677 VTAIL.n241 B 1.57403f
C678 VTAIL.n242 B 0.01047f
C679 VTAIL.t2 B 0.042513f
C680 VTAIL.n243 B 0.1915f
C681 VTAIL.n244 B 0.017495f
C682 VTAIL.n245 B 0.018561f
C683 VTAIL.n246 B 0.024748f
C684 VTAIL.n247 B 0.011086f
C685 VTAIL.n248 B 0.01047f
C686 VTAIL.n249 B 0.019485f
C687 VTAIL.n250 B 0.019485f
C688 VTAIL.n251 B 0.01047f
C689 VTAIL.n252 B 0.011086f
C690 VTAIL.n253 B 0.024748f
C691 VTAIL.n254 B 0.024748f
C692 VTAIL.n255 B 0.011086f
C693 VTAIL.n256 B 0.01047f
C694 VTAIL.n257 B 0.019485f
C695 VTAIL.n258 B 0.019485f
C696 VTAIL.n259 B 0.01047f
C697 VTAIL.n260 B 0.011086f
C698 VTAIL.n261 B 0.024748f
C699 VTAIL.n262 B 0.024748f
C700 VTAIL.n263 B 0.011086f
C701 VTAIL.n264 B 0.01047f
C702 VTAIL.n265 B 0.019485f
C703 VTAIL.n266 B 0.019485f
C704 VTAIL.n267 B 0.01047f
C705 VTAIL.n268 B 0.011086f
C706 VTAIL.n269 B 0.024748f
C707 VTAIL.n270 B 0.024748f
C708 VTAIL.n271 B 0.011086f
C709 VTAIL.n272 B 0.01047f
C710 VTAIL.n273 B 0.019485f
C711 VTAIL.n274 B 0.019485f
C712 VTAIL.n275 B 0.01047f
C713 VTAIL.n276 B 0.011086f
C714 VTAIL.n277 B 0.024748f
C715 VTAIL.n278 B 0.024748f
C716 VTAIL.n279 B 0.011086f
C717 VTAIL.n280 B 0.01047f
C718 VTAIL.n281 B 0.019485f
C719 VTAIL.n282 B 0.019485f
C720 VTAIL.n283 B 0.01047f
C721 VTAIL.n284 B 0.011086f
C722 VTAIL.n285 B 0.024748f
C723 VTAIL.n286 B 0.024748f
C724 VTAIL.n287 B 0.011086f
C725 VTAIL.n288 B 0.01047f
C726 VTAIL.n289 B 0.019485f
C727 VTAIL.n290 B 0.019485f
C728 VTAIL.n291 B 0.01047f
C729 VTAIL.n292 B 0.011086f
C730 VTAIL.n293 B 0.024748f
C731 VTAIL.n294 B 0.024748f
C732 VTAIL.n295 B 0.011086f
C733 VTAIL.n296 B 0.01047f
C734 VTAIL.n297 B 0.019485f
C735 VTAIL.n298 B 0.019485f
C736 VTAIL.n299 B 0.01047f
C737 VTAIL.n300 B 0.011086f
C738 VTAIL.n301 B 0.024748f
C739 VTAIL.n302 B 0.024748f
C740 VTAIL.n303 B 0.011086f
C741 VTAIL.n304 B 0.01047f
C742 VTAIL.n305 B 0.019485f
C743 VTAIL.n306 B 0.050894f
C744 VTAIL.n307 B 0.01047f
C745 VTAIL.n308 B 0.011086f
C746 VTAIL.n309 B 0.05125f
C747 VTAIL.n310 B 0.043373f
C748 VTAIL.n311 B 1.49482f
C749 VTAIL.n312 B 0.010994f
C750 VTAIL.n313 B 0.024748f
C751 VTAIL.n314 B 0.011086f
C752 VTAIL.n315 B 0.019485f
C753 VTAIL.n316 B 0.01047f
C754 VTAIL.n317 B 0.024748f
C755 VTAIL.n318 B 0.011086f
C756 VTAIL.n319 B 0.019485f
C757 VTAIL.n320 B 0.01047f
C758 VTAIL.n321 B 0.024748f
C759 VTAIL.n322 B 0.011086f
C760 VTAIL.n323 B 0.019485f
C761 VTAIL.n324 B 0.01047f
C762 VTAIL.n325 B 0.024748f
C763 VTAIL.n326 B 0.011086f
C764 VTAIL.n327 B 0.019485f
C765 VTAIL.n328 B 0.01047f
C766 VTAIL.n329 B 0.024748f
C767 VTAIL.n330 B 0.011086f
C768 VTAIL.n331 B 0.019485f
C769 VTAIL.n332 B 0.01047f
C770 VTAIL.n333 B 0.024748f
C771 VTAIL.n334 B 0.010778f
C772 VTAIL.n335 B 0.019485f
C773 VTAIL.n336 B 0.011086f
C774 VTAIL.n337 B 0.024748f
C775 VTAIL.n338 B 0.011086f
C776 VTAIL.n339 B 0.019485f
C777 VTAIL.n340 B 0.01047f
C778 VTAIL.n341 B 0.024748f
C779 VTAIL.n342 B 0.011086f
C780 VTAIL.n343 B 1.57403f
C781 VTAIL.n344 B 0.01047f
C782 VTAIL.t1 B 0.042513f
C783 VTAIL.n345 B 0.1915f
C784 VTAIL.n346 B 0.017495f
C785 VTAIL.n347 B 0.018561f
C786 VTAIL.n348 B 0.024748f
C787 VTAIL.n349 B 0.011086f
C788 VTAIL.n350 B 0.01047f
C789 VTAIL.n351 B 0.019485f
C790 VTAIL.n352 B 0.019485f
C791 VTAIL.n353 B 0.01047f
C792 VTAIL.n354 B 0.011086f
C793 VTAIL.n355 B 0.024748f
C794 VTAIL.n356 B 0.024748f
C795 VTAIL.n357 B 0.011086f
C796 VTAIL.n358 B 0.01047f
C797 VTAIL.n359 B 0.019485f
C798 VTAIL.n360 B 0.019485f
C799 VTAIL.n361 B 0.01047f
C800 VTAIL.n362 B 0.01047f
C801 VTAIL.n363 B 0.011086f
C802 VTAIL.n364 B 0.024748f
C803 VTAIL.n365 B 0.024748f
C804 VTAIL.n366 B 0.024748f
C805 VTAIL.n367 B 0.010778f
C806 VTAIL.n368 B 0.01047f
C807 VTAIL.n369 B 0.019485f
C808 VTAIL.n370 B 0.019485f
C809 VTAIL.n371 B 0.01047f
C810 VTAIL.n372 B 0.011086f
C811 VTAIL.n373 B 0.024748f
C812 VTAIL.n374 B 0.024748f
C813 VTAIL.n375 B 0.011086f
C814 VTAIL.n376 B 0.01047f
C815 VTAIL.n377 B 0.019485f
C816 VTAIL.n378 B 0.019485f
C817 VTAIL.n379 B 0.01047f
C818 VTAIL.n380 B 0.011086f
C819 VTAIL.n381 B 0.024748f
C820 VTAIL.n382 B 0.024748f
C821 VTAIL.n383 B 0.011086f
C822 VTAIL.n384 B 0.01047f
C823 VTAIL.n385 B 0.019485f
C824 VTAIL.n386 B 0.019485f
C825 VTAIL.n387 B 0.01047f
C826 VTAIL.n388 B 0.011086f
C827 VTAIL.n389 B 0.024748f
C828 VTAIL.n390 B 0.024748f
C829 VTAIL.n391 B 0.011086f
C830 VTAIL.n392 B 0.01047f
C831 VTAIL.n393 B 0.019485f
C832 VTAIL.n394 B 0.019485f
C833 VTAIL.n395 B 0.01047f
C834 VTAIL.n396 B 0.011086f
C835 VTAIL.n397 B 0.024748f
C836 VTAIL.n398 B 0.024748f
C837 VTAIL.n399 B 0.011086f
C838 VTAIL.n400 B 0.01047f
C839 VTAIL.n401 B 0.019485f
C840 VTAIL.n402 B 0.019485f
C841 VTAIL.n403 B 0.01047f
C842 VTAIL.n404 B 0.011086f
C843 VTAIL.n405 B 0.024748f
C844 VTAIL.n406 B 0.024748f
C845 VTAIL.n407 B 0.011086f
C846 VTAIL.n408 B 0.01047f
C847 VTAIL.n409 B 0.019485f
C848 VTAIL.n410 B 0.050894f
C849 VTAIL.n411 B 0.01047f
C850 VTAIL.n412 B 0.011086f
C851 VTAIL.n413 B 0.05125f
C852 VTAIL.n414 B 0.043373f
C853 VTAIL.n415 B 1.43461f
C854 VP.t1 B 3.99173f
C855 VP.t0 B 3.59858f
C856 VP.n0 B 5.85471f
.ends

