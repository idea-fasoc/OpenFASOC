* NGSPICE file created from diff_pair_sample_0320.ext - technology: sky130A

.subckt diff_pair_sample_0320 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0 ps=0 w=5.33 l=1.23
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0 ps=0 w=5.33 l=1.23
X2 VDD1.t3 VP.t0 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.87945 pd=5.66 as=2.0787 ps=11.44 w=5.33 l=1.23
X3 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0.87945 ps=5.66 w=5.33 l=1.23
X4 VDD1.t1 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.87945 pd=5.66 as=2.0787 ps=11.44 w=5.33 l=1.23
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0 ps=0 w=5.33 l=1.23
X6 VDD2.t3 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.87945 pd=5.66 as=2.0787 ps=11.44 w=5.33 l=1.23
X7 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.87945 pd=5.66 as=2.0787 ps=11.44 w=5.33 l=1.23
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0 ps=0 w=5.33 l=1.23
X9 VTAIL.t1 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0.87945 ps=5.66 w=5.33 l=1.23
X10 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0.87945 ps=5.66 w=5.33 l=1.23
X11 VTAIL.t7 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0787 pd=11.44 as=0.87945 ps=5.66 w=5.33 l=1.23
R0 B.n355 B.n354 585
R1 B.n356 B.n76 585
R2 B.n358 B.n357 585
R3 B.n360 B.n75 585
R4 B.n363 B.n362 585
R5 B.n364 B.n74 585
R6 B.n366 B.n365 585
R7 B.n368 B.n73 585
R8 B.n371 B.n370 585
R9 B.n372 B.n72 585
R10 B.n374 B.n373 585
R11 B.n376 B.n71 585
R12 B.n379 B.n378 585
R13 B.n380 B.n70 585
R14 B.n382 B.n381 585
R15 B.n384 B.n69 585
R16 B.n387 B.n386 585
R17 B.n388 B.n68 585
R18 B.n390 B.n389 585
R19 B.n392 B.n67 585
R20 B.n394 B.n393 585
R21 B.n396 B.n395 585
R22 B.n399 B.n398 585
R23 B.n400 B.n62 585
R24 B.n402 B.n401 585
R25 B.n404 B.n61 585
R26 B.n407 B.n406 585
R27 B.n408 B.n60 585
R28 B.n410 B.n409 585
R29 B.n412 B.n59 585
R30 B.n414 B.n413 585
R31 B.n416 B.n415 585
R32 B.n419 B.n418 585
R33 B.n420 B.n54 585
R34 B.n422 B.n421 585
R35 B.n424 B.n53 585
R36 B.n427 B.n426 585
R37 B.n428 B.n52 585
R38 B.n430 B.n429 585
R39 B.n432 B.n51 585
R40 B.n435 B.n434 585
R41 B.n436 B.n50 585
R42 B.n438 B.n437 585
R43 B.n440 B.n49 585
R44 B.n443 B.n442 585
R45 B.n444 B.n48 585
R46 B.n446 B.n445 585
R47 B.n448 B.n47 585
R48 B.n451 B.n450 585
R49 B.n452 B.n46 585
R50 B.n454 B.n453 585
R51 B.n456 B.n45 585
R52 B.n459 B.n458 585
R53 B.n460 B.n44 585
R54 B.n352 B.n42 585
R55 B.n463 B.n42 585
R56 B.n351 B.n41 585
R57 B.n464 B.n41 585
R58 B.n350 B.n40 585
R59 B.n465 B.n40 585
R60 B.n349 B.n348 585
R61 B.n348 B.n36 585
R62 B.n347 B.n35 585
R63 B.n471 B.n35 585
R64 B.n346 B.n34 585
R65 B.n472 B.n34 585
R66 B.n345 B.n33 585
R67 B.n473 B.n33 585
R68 B.n344 B.n343 585
R69 B.n343 B.n29 585
R70 B.n342 B.n28 585
R71 B.n479 B.n28 585
R72 B.n341 B.n27 585
R73 B.n480 B.n27 585
R74 B.n340 B.n26 585
R75 B.n481 B.n26 585
R76 B.n339 B.n338 585
R77 B.n338 B.n22 585
R78 B.n337 B.n21 585
R79 B.n487 B.n21 585
R80 B.n336 B.n20 585
R81 B.n488 B.n20 585
R82 B.n335 B.n19 585
R83 B.n489 B.n19 585
R84 B.n334 B.n333 585
R85 B.n333 B.n15 585
R86 B.n332 B.n14 585
R87 B.n495 B.n14 585
R88 B.n331 B.n13 585
R89 B.n496 B.n13 585
R90 B.n330 B.n12 585
R91 B.n497 B.n12 585
R92 B.n329 B.n328 585
R93 B.n328 B.n8 585
R94 B.n327 B.n7 585
R95 B.n503 B.n7 585
R96 B.n326 B.n6 585
R97 B.n504 B.n6 585
R98 B.n325 B.n5 585
R99 B.n505 B.n5 585
R100 B.n324 B.n323 585
R101 B.n323 B.n4 585
R102 B.n322 B.n77 585
R103 B.n322 B.n321 585
R104 B.n312 B.n78 585
R105 B.n79 B.n78 585
R106 B.n314 B.n313 585
R107 B.n315 B.n314 585
R108 B.n311 B.n84 585
R109 B.n84 B.n83 585
R110 B.n310 B.n309 585
R111 B.n309 B.n308 585
R112 B.n86 B.n85 585
R113 B.n87 B.n86 585
R114 B.n301 B.n300 585
R115 B.n302 B.n301 585
R116 B.n299 B.n91 585
R117 B.n95 B.n91 585
R118 B.n298 B.n297 585
R119 B.n297 B.n296 585
R120 B.n93 B.n92 585
R121 B.n94 B.n93 585
R122 B.n289 B.n288 585
R123 B.n290 B.n289 585
R124 B.n287 B.n100 585
R125 B.n100 B.n99 585
R126 B.n286 B.n285 585
R127 B.n285 B.n284 585
R128 B.n102 B.n101 585
R129 B.n103 B.n102 585
R130 B.n277 B.n276 585
R131 B.n278 B.n277 585
R132 B.n275 B.n107 585
R133 B.n111 B.n107 585
R134 B.n274 B.n273 585
R135 B.n273 B.n272 585
R136 B.n109 B.n108 585
R137 B.n110 B.n109 585
R138 B.n265 B.n264 585
R139 B.n266 B.n265 585
R140 B.n263 B.n116 585
R141 B.n116 B.n115 585
R142 B.n262 B.n261 585
R143 B.n261 B.n260 585
R144 B.n257 B.n120 585
R145 B.n256 B.n255 585
R146 B.n253 B.n121 585
R147 B.n253 B.n119 585
R148 B.n252 B.n251 585
R149 B.n250 B.n249 585
R150 B.n248 B.n123 585
R151 B.n246 B.n245 585
R152 B.n244 B.n124 585
R153 B.n243 B.n242 585
R154 B.n240 B.n125 585
R155 B.n238 B.n237 585
R156 B.n236 B.n126 585
R157 B.n235 B.n234 585
R158 B.n232 B.n127 585
R159 B.n230 B.n229 585
R160 B.n228 B.n128 585
R161 B.n227 B.n226 585
R162 B.n224 B.n129 585
R163 B.n222 B.n221 585
R164 B.n220 B.n130 585
R165 B.n219 B.n218 585
R166 B.n216 B.n131 585
R167 B.n214 B.n213 585
R168 B.n212 B.n132 585
R169 B.n211 B.n210 585
R170 B.n208 B.n136 585
R171 B.n206 B.n205 585
R172 B.n204 B.n137 585
R173 B.n203 B.n202 585
R174 B.n200 B.n138 585
R175 B.n198 B.n197 585
R176 B.n196 B.n139 585
R177 B.n194 B.n193 585
R178 B.n191 B.n142 585
R179 B.n189 B.n188 585
R180 B.n187 B.n143 585
R181 B.n186 B.n185 585
R182 B.n183 B.n144 585
R183 B.n181 B.n180 585
R184 B.n179 B.n145 585
R185 B.n178 B.n177 585
R186 B.n175 B.n146 585
R187 B.n173 B.n172 585
R188 B.n171 B.n147 585
R189 B.n170 B.n169 585
R190 B.n167 B.n148 585
R191 B.n165 B.n164 585
R192 B.n163 B.n149 585
R193 B.n162 B.n161 585
R194 B.n159 B.n150 585
R195 B.n157 B.n156 585
R196 B.n155 B.n151 585
R197 B.n154 B.n153 585
R198 B.n118 B.n117 585
R199 B.n119 B.n118 585
R200 B.n259 B.n258 585
R201 B.n260 B.n259 585
R202 B.n114 B.n113 585
R203 B.n115 B.n114 585
R204 B.n268 B.n267 585
R205 B.n267 B.n266 585
R206 B.n269 B.n112 585
R207 B.n112 B.n110 585
R208 B.n271 B.n270 585
R209 B.n272 B.n271 585
R210 B.n106 B.n105 585
R211 B.n111 B.n106 585
R212 B.n280 B.n279 585
R213 B.n279 B.n278 585
R214 B.n281 B.n104 585
R215 B.n104 B.n103 585
R216 B.n283 B.n282 585
R217 B.n284 B.n283 585
R218 B.n98 B.n97 585
R219 B.n99 B.n98 585
R220 B.n292 B.n291 585
R221 B.n291 B.n290 585
R222 B.n293 B.n96 585
R223 B.n96 B.n94 585
R224 B.n295 B.n294 585
R225 B.n296 B.n295 585
R226 B.n90 B.n89 585
R227 B.n95 B.n90 585
R228 B.n304 B.n303 585
R229 B.n303 B.n302 585
R230 B.n305 B.n88 585
R231 B.n88 B.n87 585
R232 B.n307 B.n306 585
R233 B.n308 B.n307 585
R234 B.n82 B.n81 585
R235 B.n83 B.n82 585
R236 B.n317 B.n316 585
R237 B.n316 B.n315 585
R238 B.n318 B.n80 585
R239 B.n80 B.n79 585
R240 B.n320 B.n319 585
R241 B.n321 B.n320 585
R242 B.n2 B.n0 585
R243 B.n4 B.n2 585
R244 B.n3 B.n1 585
R245 B.n504 B.n3 585
R246 B.n502 B.n501 585
R247 B.n503 B.n502 585
R248 B.n500 B.n9 585
R249 B.n9 B.n8 585
R250 B.n499 B.n498 585
R251 B.n498 B.n497 585
R252 B.n11 B.n10 585
R253 B.n496 B.n11 585
R254 B.n494 B.n493 585
R255 B.n495 B.n494 585
R256 B.n492 B.n16 585
R257 B.n16 B.n15 585
R258 B.n491 B.n490 585
R259 B.n490 B.n489 585
R260 B.n18 B.n17 585
R261 B.n488 B.n18 585
R262 B.n486 B.n485 585
R263 B.n487 B.n486 585
R264 B.n484 B.n23 585
R265 B.n23 B.n22 585
R266 B.n483 B.n482 585
R267 B.n482 B.n481 585
R268 B.n25 B.n24 585
R269 B.n480 B.n25 585
R270 B.n478 B.n477 585
R271 B.n479 B.n478 585
R272 B.n476 B.n30 585
R273 B.n30 B.n29 585
R274 B.n475 B.n474 585
R275 B.n474 B.n473 585
R276 B.n32 B.n31 585
R277 B.n472 B.n32 585
R278 B.n470 B.n469 585
R279 B.n471 B.n470 585
R280 B.n468 B.n37 585
R281 B.n37 B.n36 585
R282 B.n467 B.n466 585
R283 B.n466 B.n465 585
R284 B.n39 B.n38 585
R285 B.n464 B.n39 585
R286 B.n462 B.n461 585
R287 B.n463 B.n462 585
R288 B.n507 B.n506 585
R289 B.n506 B.n505 585
R290 B.n259 B.n120 444.452
R291 B.n462 B.n44 444.452
R292 B.n261 B.n118 444.452
R293 B.n354 B.n42 444.452
R294 B.n140 B.t12 308.704
R295 B.n133 B.t8 308.704
R296 B.n55 B.t15 308.704
R297 B.n63 B.t4 308.704
R298 B.n353 B.n43 256.663
R299 B.n359 B.n43 256.663
R300 B.n361 B.n43 256.663
R301 B.n367 B.n43 256.663
R302 B.n369 B.n43 256.663
R303 B.n375 B.n43 256.663
R304 B.n377 B.n43 256.663
R305 B.n383 B.n43 256.663
R306 B.n385 B.n43 256.663
R307 B.n391 B.n43 256.663
R308 B.n66 B.n43 256.663
R309 B.n397 B.n43 256.663
R310 B.n403 B.n43 256.663
R311 B.n405 B.n43 256.663
R312 B.n411 B.n43 256.663
R313 B.n58 B.n43 256.663
R314 B.n417 B.n43 256.663
R315 B.n423 B.n43 256.663
R316 B.n425 B.n43 256.663
R317 B.n431 B.n43 256.663
R318 B.n433 B.n43 256.663
R319 B.n439 B.n43 256.663
R320 B.n441 B.n43 256.663
R321 B.n447 B.n43 256.663
R322 B.n449 B.n43 256.663
R323 B.n455 B.n43 256.663
R324 B.n457 B.n43 256.663
R325 B.n254 B.n119 256.663
R326 B.n122 B.n119 256.663
R327 B.n247 B.n119 256.663
R328 B.n241 B.n119 256.663
R329 B.n239 B.n119 256.663
R330 B.n233 B.n119 256.663
R331 B.n231 B.n119 256.663
R332 B.n225 B.n119 256.663
R333 B.n223 B.n119 256.663
R334 B.n217 B.n119 256.663
R335 B.n215 B.n119 256.663
R336 B.n209 B.n119 256.663
R337 B.n207 B.n119 256.663
R338 B.n201 B.n119 256.663
R339 B.n199 B.n119 256.663
R340 B.n192 B.n119 256.663
R341 B.n190 B.n119 256.663
R342 B.n184 B.n119 256.663
R343 B.n182 B.n119 256.663
R344 B.n176 B.n119 256.663
R345 B.n174 B.n119 256.663
R346 B.n168 B.n119 256.663
R347 B.n166 B.n119 256.663
R348 B.n160 B.n119 256.663
R349 B.n158 B.n119 256.663
R350 B.n152 B.n119 256.663
R351 B.n140 B.t14 197.798
R352 B.n63 B.t6 197.798
R353 B.n133 B.t11 197.798
R354 B.n55 B.t16 197.798
R355 B.n141 B.t13 167.543
R356 B.n64 B.t7 167.543
R357 B.n134 B.t10 167.543
R358 B.n56 B.t17 167.543
R359 B.n259 B.n114 163.367
R360 B.n267 B.n114 163.367
R361 B.n267 B.n112 163.367
R362 B.n271 B.n112 163.367
R363 B.n271 B.n106 163.367
R364 B.n279 B.n106 163.367
R365 B.n279 B.n104 163.367
R366 B.n283 B.n104 163.367
R367 B.n283 B.n98 163.367
R368 B.n291 B.n98 163.367
R369 B.n291 B.n96 163.367
R370 B.n295 B.n96 163.367
R371 B.n295 B.n90 163.367
R372 B.n303 B.n90 163.367
R373 B.n303 B.n88 163.367
R374 B.n307 B.n88 163.367
R375 B.n307 B.n82 163.367
R376 B.n316 B.n82 163.367
R377 B.n316 B.n80 163.367
R378 B.n320 B.n80 163.367
R379 B.n320 B.n2 163.367
R380 B.n506 B.n2 163.367
R381 B.n506 B.n3 163.367
R382 B.n502 B.n3 163.367
R383 B.n502 B.n9 163.367
R384 B.n498 B.n9 163.367
R385 B.n498 B.n11 163.367
R386 B.n494 B.n11 163.367
R387 B.n494 B.n16 163.367
R388 B.n490 B.n16 163.367
R389 B.n490 B.n18 163.367
R390 B.n486 B.n18 163.367
R391 B.n486 B.n23 163.367
R392 B.n482 B.n23 163.367
R393 B.n482 B.n25 163.367
R394 B.n478 B.n25 163.367
R395 B.n478 B.n30 163.367
R396 B.n474 B.n30 163.367
R397 B.n474 B.n32 163.367
R398 B.n470 B.n32 163.367
R399 B.n470 B.n37 163.367
R400 B.n466 B.n37 163.367
R401 B.n466 B.n39 163.367
R402 B.n462 B.n39 163.367
R403 B.n255 B.n253 163.367
R404 B.n253 B.n252 163.367
R405 B.n249 B.n248 163.367
R406 B.n246 B.n124 163.367
R407 B.n242 B.n240 163.367
R408 B.n238 B.n126 163.367
R409 B.n234 B.n232 163.367
R410 B.n230 B.n128 163.367
R411 B.n226 B.n224 163.367
R412 B.n222 B.n130 163.367
R413 B.n218 B.n216 163.367
R414 B.n214 B.n132 163.367
R415 B.n210 B.n208 163.367
R416 B.n206 B.n137 163.367
R417 B.n202 B.n200 163.367
R418 B.n198 B.n139 163.367
R419 B.n193 B.n191 163.367
R420 B.n189 B.n143 163.367
R421 B.n185 B.n183 163.367
R422 B.n181 B.n145 163.367
R423 B.n177 B.n175 163.367
R424 B.n173 B.n147 163.367
R425 B.n169 B.n167 163.367
R426 B.n165 B.n149 163.367
R427 B.n161 B.n159 163.367
R428 B.n157 B.n151 163.367
R429 B.n153 B.n118 163.367
R430 B.n261 B.n116 163.367
R431 B.n265 B.n116 163.367
R432 B.n265 B.n109 163.367
R433 B.n273 B.n109 163.367
R434 B.n273 B.n107 163.367
R435 B.n277 B.n107 163.367
R436 B.n277 B.n102 163.367
R437 B.n285 B.n102 163.367
R438 B.n285 B.n100 163.367
R439 B.n289 B.n100 163.367
R440 B.n289 B.n93 163.367
R441 B.n297 B.n93 163.367
R442 B.n297 B.n91 163.367
R443 B.n301 B.n91 163.367
R444 B.n301 B.n86 163.367
R445 B.n309 B.n86 163.367
R446 B.n309 B.n84 163.367
R447 B.n314 B.n84 163.367
R448 B.n314 B.n78 163.367
R449 B.n322 B.n78 163.367
R450 B.n323 B.n322 163.367
R451 B.n323 B.n5 163.367
R452 B.n6 B.n5 163.367
R453 B.n7 B.n6 163.367
R454 B.n328 B.n7 163.367
R455 B.n328 B.n12 163.367
R456 B.n13 B.n12 163.367
R457 B.n14 B.n13 163.367
R458 B.n333 B.n14 163.367
R459 B.n333 B.n19 163.367
R460 B.n20 B.n19 163.367
R461 B.n21 B.n20 163.367
R462 B.n338 B.n21 163.367
R463 B.n338 B.n26 163.367
R464 B.n27 B.n26 163.367
R465 B.n28 B.n27 163.367
R466 B.n343 B.n28 163.367
R467 B.n343 B.n33 163.367
R468 B.n34 B.n33 163.367
R469 B.n35 B.n34 163.367
R470 B.n348 B.n35 163.367
R471 B.n348 B.n40 163.367
R472 B.n41 B.n40 163.367
R473 B.n42 B.n41 163.367
R474 B.n458 B.n456 163.367
R475 B.n454 B.n46 163.367
R476 B.n450 B.n448 163.367
R477 B.n446 B.n48 163.367
R478 B.n442 B.n440 163.367
R479 B.n438 B.n50 163.367
R480 B.n434 B.n432 163.367
R481 B.n430 B.n52 163.367
R482 B.n426 B.n424 163.367
R483 B.n422 B.n54 163.367
R484 B.n418 B.n416 163.367
R485 B.n413 B.n412 163.367
R486 B.n410 B.n60 163.367
R487 B.n406 B.n404 163.367
R488 B.n402 B.n62 163.367
R489 B.n398 B.n396 163.367
R490 B.n393 B.n392 163.367
R491 B.n390 B.n68 163.367
R492 B.n386 B.n384 163.367
R493 B.n382 B.n70 163.367
R494 B.n378 B.n376 163.367
R495 B.n374 B.n72 163.367
R496 B.n370 B.n368 163.367
R497 B.n366 B.n74 163.367
R498 B.n362 B.n360 163.367
R499 B.n358 B.n76 163.367
R500 B.n260 B.n119 119.284
R501 B.n463 B.n43 119.284
R502 B.n254 B.n120 71.676
R503 B.n252 B.n122 71.676
R504 B.n248 B.n247 71.676
R505 B.n241 B.n124 71.676
R506 B.n240 B.n239 71.676
R507 B.n233 B.n126 71.676
R508 B.n232 B.n231 71.676
R509 B.n225 B.n128 71.676
R510 B.n224 B.n223 71.676
R511 B.n217 B.n130 71.676
R512 B.n216 B.n215 71.676
R513 B.n209 B.n132 71.676
R514 B.n208 B.n207 71.676
R515 B.n201 B.n137 71.676
R516 B.n200 B.n199 71.676
R517 B.n192 B.n139 71.676
R518 B.n191 B.n190 71.676
R519 B.n184 B.n143 71.676
R520 B.n183 B.n182 71.676
R521 B.n176 B.n145 71.676
R522 B.n175 B.n174 71.676
R523 B.n168 B.n147 71.676
R524 B.n167 B.n166 71.676
R525 B.n160 B.n149 71.676
R526 B.n159 B.n158 71.676
R527 B.n152 B.n151 71.676
R528 B.n457 B.n44 71.676
R529 B.n456 B.n455 71.676
R530 B.n449 B.n46 71.676
R531 B.n448 B.n447 71.676
R532 B.n441 B.n48 71.676
R533 B.n440 B.n439 71.676
R534 B.n433 B.n50 71.676
R535 B.n432 B.n431 71.676
R536 B.n425 B.n52 71.676
R537 B.n424 B.n423 71.676
R538 B.n417 B.n54 71.676
R539 B.n416 B.n58 71.676
R540 B.n412 B.n411 71.676
R541 B.n405 B.n60 71.676
R542 B.n404 B.n403 71.676
R543 B.n397 B.n62 71.676
R544 B.n396 B.n66 71.676
R545 B.n392 B.n391 71.676
R546 B.n385 B.n68 71.676
R547 B.n384 B.n383 71.676
R548 B.n377 B.n70 71.676
R549 B.n376 B.n375 71.676
R550 B.n369 B.n72 71.676
R551 B.n368 B.n367 71.676
R552 B.n361 B.n74 71.676
R553 B.n360 B.n359 71.676
R554 B.n353 B.n76 71.676
R555 B.n354 B.n353 71.676
R556 B.n359 B.n358 71.676
R557 B.n362 B.n361 71.676
R558 B.n367 B.n366 71.676
R559 B.n370 B.n369 71.676
R560 B.n375 B.n374 71.676
R561 B.n378 B.n377 71.676
R562 B.n383 B.n382 71.676
R563 B.n386 B.n385 71.676
R564 B.n391 B.n390 71.676
R565 B.n393 B.n66 71.676
R566 B.n398 B.n397 71.676
R567 B.n403 B.n402 71.676
R568 B.n406 B.n405 71.676
R569 B.n411 B.n410 71.676
R570 B.n413 B.n58 71.676
R571 B.n418 B.n417 71.676
R572 B.n423 B.n422 71.676
R573 B.n426 B.n425 71.676
R574 B.n431 B.n430 71.676
R575 B.n434 B.n433 71.676
R576 B.n439 B.n438 71.676
R577 B.n442 B.n441 71.676
R578 B.n447 B.n446 71.676
R579 B.n450 B.n449 71.676
R580 B.n455 B.n454 71.676
R581 B.n458 B.n457 71.676
R582 B.n255 B.n254 71.676
R583 B.n249 B.n122 71.676
R584 B.n247 B.n246 71.676
R585 B.n242 B.n241 71.676
R586 B.n239 B.n238 71.676
R587 B.n234 B.n233 71.676
R588 B.n231 B.n230 71.676
R589 B.n226 B.n225 71.676
R590 B.n223 B.n222 71.676
R591 B.n218 B.n217 71.676
R592 B.n215 B.n214 71.676
R593 B.n210 B.n209 71.676
R594 B.n207 B.n206 71.676
R595 B.n202 B.n201 71.676
R596 B.n199 B.n198 71.676
R597 B.n193 B.n192 71.676
R598 B.n190 B.n189 71.676
R599 B.n185 B.n184 71.676
R600 B.n182 B.n181 71.676
R601 B.n177 B.n176 71.676
R602 B.n174 B.n173 71.676
R603 B.n169 B.n168 71.676
R604 B.n166 B.n165 71.676
R605 B.n161 B.n160 71.676
R606 B.n158 B.n157 71.676
R607 B.n153 B.n152 71.676
R608 B.n260 B.n115 70.5333
R609 B.n266 B.n115 70.5333
R610 B.n266 B.n110 70.5333
R611 B.n272 B.n110 70.5333
R612 B.n272 B.n111 70.5333
R613 B.n278 B.n103 70.5333
R614 B.n284 B.n103 70.5333
R615 B.n284 B.n99 70.5333
R616 B.n290 B.n99 70.5333
R617 B.n290 B.n94 70.5333
R618 B.n296 B.n94 70.5333
R619 B.n296 B.n95 70.5333
R620 B.n302 B.n87 70.5333
R621 B.n308 B.n87 70.5333
R622 B.n308 B.n83 70.5333
R623 B.n315 B.n83 70.5333
R624 B.n321 B.n79 70.5333
R625 B.n321 B.n4 70.5333
R626 B.n505 B.n4 70.5333
R627 B.n505 B.n504 70.5333
R628 B.n504 B.n503 70.5333
R629 B.n503 B.n8 70.5333
R630 B.n497 B.n496 70.5333
R631 B.n496 B.n495 70.5333
R632 B.n495 B.n15 70.5333
R633 B.n489 B.n15 70.5333
R634 B.n488 B.n487 70.5333
R635 B.n487 B.n22 70.5333
R636 B.n481 B.n22 70.5333
R637 B.n481 B.n480 70.5333
R638 B.n480 B.n479 70.5333
R639 B.n479 B.n29 70.5333
R640 B.n473 B.n29 70.5333
R641 B.n472 B.n471 70.5333
R642 B.n471 B.n36 70.5333
R643 B.n465 B.n36 70.5333
R644 B.n465 B.n464 70.5333
R645 B.n464 B.n463 70.5333
R646 B.t3 B.n79 63.2725
R647 B.t0 B.n8 63.2725
R648 B.n195 B.n141 59.5399
R649 B.n135 B.n134 59.5399
R650 B.n57 B.n56 59.5399
R651 B.n65 B.n64 59.5399
R652 B.n111 B.t9 50.8256
R653 B.t5 B.n472 50.8256
R654 B.n95 B.t2 36.3041
R655 B.t1 B.n488 36.3041
R656 B.n302 B.t2 34.2296
R657 B.n489 B.t1 34.2296
R658 B.n141 B.n140 30.255
R659 B.n134 B.n133 30.255
R660 B.n56 B.n55 30.255
R661 B.n64 B.n63 30.255
R662 B.n355 B.n352 28.8785
R663 B.n461 B.n460 28.8785
R664 B.n262 B.n117 28.8785
R665 B.n258 B.n257 28.8785
R666 B.n278 B.t9 19.7082
R667 B.n473 B.t5 19.7082
R668 B B.n507 18.0485
R669 B.n460 B.n459 10.6151
R670 B.n459 B.n45 10.6151
R671 B.n453 B.n45 10.6151
R672 B.n453 B.n452 10.6151
R673 B.n452 B.n451 10.6151
R674 B.n451 B.n47 10.6151
R675 B.n445 B.n47 10.6151
R676 B.n445 B.n444 10.6151
R677 B.n444 B.n443 10.6151
R678 B.n443 B.n49 10.6151
R679 B.n437 B.n49 10.6151
R680 B.n437 B.n436 10.6151
R681 B.n436 B.n435 10.6151
R682 B.n435 B.n51 10.6151
R683 B.n429 B.n51 10.6151
R684 B.n429 B.n428 10.6151
R685 B.n428 B.n427 10.6151
R686 B.n427 B.n53 10.6151
R687 B.n421 B.n53 10.6151
R688 B.n421 B.n420 10.6151
R689 B.n420 B.n419 10.6151
R690 B.n415 B.n414 10.6151
R691 B.n414 B.n59 10.6151
R692 B.n409 B.n59 10.6151
R693 B.n409 B.n408 10.6151
R694 B.n408 B.n407 10.6151
R695 B.n407 B.n61 10.6151
R696 B.n401 B.n61 10.6151
R697 B.n401 B.n400 10.6151
R698 B.n400 B.n399 10.6151
R699 B.n395 B.n394 10.6151
R700 B.n394 B.n67 10.6151
R701 B.n389 B.n67 10.6151
R702 B.n389 B.n388 10.6151
R703 B.n388 B.n387 10.6151
R704 B.n387 B.n69 10.6151
R705 B.n381 B.n69 10.6151
R706 B.n381 B.n380 10.6151
R707 B.n380 B.n379 10.6151
R708 B.n379 B.n71 10.6151
R709 B.n373 B.n71 10.6151
R710 B.n373 B.n372 10.6151
R711 B.n372 B.n371 10.6151
R712 B.n371 B.n73 10.6151
R713 B.n365 B.n73 10.6151
R714 B.n365 B.n364 10.6151
R715 B.n364 B.n363 10.6151
R716 B.n363 B.n75 10.6151
R717 B.n357 B.n75 10.6151
R718 B.n357 B.n356 10.6151
R719 B.n356 B.n355 10.6151
R720 B.n263 B.n262 10.6151
R721 B.n264 B.n263 10.6151
R722 B.n264 B.n108 10.6151
R723 B.n274 B.n108 10.6151
R724 B.n275 B.n274 10.6151
R725 B.n276 B.n275 10.6151
R726 B.n276 B.n101 10.6151
R727 B.n286 B.n101 10.6151
R728 B.n287 B.n286 10.6151
R729 B.n288 B.n287 10.6151
R730 B.n288 B.n92 10.6151
R731 B.n298 B.n92 10.6151
R732 B.n299 B.n298 10.6151
R733 B.n300 B.n299 10.6151
R734 B.n300 B.n85 10.6151
R735 B.n310 B.n85 10.6151
R736 B.n311 B.n310 10.6151
R737 B.n313 B.n311 10.6151
R738 B.n313 B.n312 10.6151
R739 B.n312 B.n77 10.6151
R740 B.n324 B.n77 10.6151
R741 B.n325 B.n324 10.6151
R742 B.n326 B.n325 10.6151
R743 B.n327 B.n326 10.6151
R744 B.n329 B.n327 10.6151
R745 B.n330 B.n329 10.6151
R746 B.n331 B.n330 10.6151
R747 B.n332 B.n331 10.6151
R748 B.n334 B.n332 10.6151
R749 B.n335 B.n334 10.6151
R750 B.n336 B.n335 10.6151
R751 B.n337 B.n336 10.6151
R752 B.n339 B.n337 10.6151
R753 B.n340 B.n339 10.6151
R754 B.n341 B.n340 10.6151
R755 B.n342 B.n341 10.6151
R756 B.n344 B.n342 10.6151
R757 B.n345 B.n344 10.6151
R758 B.n346 B.n345 10.6151
R759 B.n347 B.n346 10.6151
R760 B.n349 B.n347 10.6151
R761 B.n350 B.n349 10.6151
R762 B.n351 B.n350 10.6151
R763 B.n352 B.n351 10.6151
R764 B.n257 B.n256 10.6151
R765 B.n256 B.n121 10.6151
R766 B.n251 B.n121 10.6151
R767 B.n251 B.n250 10.6151
R768 B.n250 B.n123 10.6151
R769 B.n245 B.n123 10.6151
R770 B.n245 B.n244 10.6151
R771 B.n244 B.n243 10.6151
R772 B.n243 B.n125 10.6151
R773 B.n237 B.n125 10.6151
R774 B.n237 B.n236 10.6151
R775 B.n236 B.n235 10.6151
R776 B.n235 B.n127 10.6151
R777 B.n229 B.n127 10.6151
R778 B.n229 B.n228 10.6151
R779 B.n228 B.n227 10.6151
R780 B.n227 B.n129 10.6151
R781 B.n221 B.n129 10.6151
R782 B.n221 B.n220 10.6151
R783 B.n220 B.n219 10.6151
R784 B.n219 B.n131 10.6151
R785 B.n213 B.n212 10.6151
R786 B.n212 B.n211 10.6151
R787 B.n211 B.n136 10.6151
R788 B.n205 B.n136 10.6151
R789 B.n205 B.n204 10.6151
R790 B.n204 B.n203 10.6151
R791 B.n203 B.n138 10.6151
R792 B.n197 B.n138 10.6151
R793 B.n197 B.n196 10.6151
R794 B.n194 B.n142 10.6151
R795 B.n188 B.n142 10.6151
R796 B.n188 B.n187 10.6151
R797 B.n187 B.n186 10.6151
R798 B.n186 B.n144 10.6151
R799 B.n180 B.n144 10.6151
R800 B.n180 B.n179 10.6151
R801 B.n179 B.n178 10.6151
R802 B.n178 B.n146 10.6151
R803 B.n172 B.n146 10.6151
R804 B.n172 B.n171 10.6151
R805 B.n171 B.n170 10.6151
R806 B.n170 B.n148 10.6151
R807 B.n164 B.n148 10.6151
R808 B.n164 B.n163 10.6151
R809 B.n163 B.n162 10.6151
R810 B.n162 B.n150 10.6151
R811 B.n156 B.n150 10.6151
R812 B.n156 B.n155 10.6151
R813 B.n155 B.n154 10.6151
R814 B.n154 B.n117 10.6151
R815 B.n258 B.n113 10.6151
R816 B.n268 B.n113 10.6151
R817 B.n269 B.n268 10.6151
R818 B.n270 B.n269 10.6151
R819 B.n270 B.n105 10.6151
R820 B.n280 B.n105 10.6151
R821 B.n281 B.n280 10.6151
R822 B.n282 B.n281 10.6151
R823 B.n282 B.n97 10.6151
R824 B.n292 B.n97 10.6151
R825 B.n293 B.n292 10.6151
R826 B.n294 B.n293 10.6151
R827 B.n294 B.n89 10.6151
R828 B.n304 B.n89 10.6151
R829 B.n305 B.n304 10.6151
R830 B.n306 B.n305 10.6151
R831 B.n306 B.n81 10.6151
R832 B.n317 B.n81 10.6151
R833 B.n318 B.n317 10.6151
R834 B.n319 B.n318 10.6151
R835 B.n319 B.n0 10.6151
R836 B.n501 B.n1 10.6151
R837 B.n501 B.n500 10.6151
R838 B.n500 B.n499 10.6151
R839 B.n499 B.n10 10.6151
R840 B.n493 B.n10 10.6151
R841 B.n493 B.n492 10.6151
R842 B.n492 B.n491 10.6151
R843 B.n491 B.n17 10.6151
R844 B.n485 B.n17 10.6151
R845 B.n485 B.n484 10.6151
R846 B.n484 B.n483 10.6151
R847 B.n483 B.n24 10.6151
R848 B.n477 B.n24 10.6151
R849 B.n477 B.n476 10.6151
R850 B.n476 B.n475 10.6151
R851 B.n475 B.n31 10.6151
R852 B.n469 B.n31 10.6151
R853 B.n469 B.n468 10.6151
R854 B.n468 B.n467 10.6151
R855 B.n467 B.n38 10.6151
R856 B.n461 B.n38 10.6151
R857 B.n419 B.n57 9.36635
R858 B.n395 B.n65 9.36635
R859 B.n135 B.n131 9.36635
R860 B.n195 B.n194 9.36635
R861 B.n315 B.t3 7.26123
R862 B.n497 B.t0 7.26123
R863 B.n507 B.n0 2.81026
R864 B.n507 B.n1 2.81026
R865 B.n415 B.n57 1.24928
R866 B.n399 B.n65 1.24928
R867 B.n213 B.n135 1.24928
R868 B.n196 B.n195 1.24928
R869 VP.n4 VP.n3 172.065
R870 VP.n10 VP.n9 172.065
R871 VP.n8 VP.n0 161.3
R872 VP.n7 VP.n6 161.3
R873 VP.n5 VP.n1 161.3
R874 VP.n2 VP.t3 140.919
R875 VP.n2 VP.t0 140.698
R876 VP.n3 VP.t1 104.433
R877 VP.n9 VP.t2 104.433
R878 VP.n4 VP.n2 55.289
R879 VP.n7 VP.n1 40.4934
R880 VP.n8 VP.n7 40.4934
R881 VP.n3 VP.n1 13.702
R882 VP.n9 VP.n8 13.702
R883 VP.n5 VP.n4 0.189894
R884 VP.n6 VP.n5 0.189894
R885 VP.n6 VP.n0 0.189894
R886 VP.n10 VP.n0 0.189894
R887 VP VP.n10 0.0516364
R888 VTAIL.n218 VTAIL.n196 289.615
R889 VTAIL.n22 VTAIL.n0 289.615
R890 VTAIL.n50 VTAIL.n28 289.615
R891 VTAIL.n78 VTAIL.n56 289.615
R892 VTAIL.n190 VTAIL.n168 289.615
R893 VTAIL.n162 VTAIL.n140 289.615
R894 VTAIL.n134 VTAIL.n112 289.615
R895 VTAIL.n106 VTAIL.n84 289.615
R896 VTAIL.n204 VTAIL.n203 185
R897 VTAIL.n209 VTAIL.n208 185
R898 VTAIL.n211 VTAIL.n210 185
R899 VTAIL.n200 VTAIL.n199 185
R900 VTAIL.n217 VTAIL.n216 185
R901 VTAIL.n219 VTAIL.n218 185
R902 VTAIL.n8 VTAIL.n7 185
R903 VTAIL.n13 VTAIL.n12 185
R904 VTAIL.n15 VTAIL.n14 185
R905 VTAIL.n4 VTAIL.n3 185
R906 VTAIL.n21 VTAIL.n20 185
R907 VTAIL.n23 VTAIL.n22 185
R908 VTAIL.n36 VTAIL.n35 185
R909 VTAIL.n41 VTAIL.n40 185
R910 VTAIL.n43 VTAIL.n42 185
R911 VTAIL.n32 VTAIL.n31 185
R912 VTAIL.n49 VTAIL.n48 185
R913 VTAIL.n51 VTAIL.n50 185
R914 VTAIL.n64 VTAIL.n63 185
R915 VTAIL.n69 VTAIL.n68 185
R916 VTAIL.n71 VTAIL.n70 185
R917 VTAIL.n60 VTAIL.n59 185
R918 VTAIL.n77 VTAIL.n76 185
R919 VTAIL.n79 VTAIL.n78 185
R920 VTAIL.n191 VTAIL.n190 185
R921 VTAIL.n189 VTAIL.n188 185
R922 VTAIL.n172 VTAIL.n171 185
R923 VTAIL.n183 VTAIL.n182 185
R924 VTAIL.n181 VTAIL.n180 185
R925 VTAIL.n176 VTAIL.n175 185
R926 VTAIL.n163 VTAIL.n162 185
R927 VTAIL.n161 VTAIL.n160 185
R928 VTAIL.n144 VTAIL.n143 185
R929 VTAIL.n155 VTAIL.n154 185
R930 VTAIL.n153 VTAIL.n152 185
R931 VTAIL.n148 VTAIL.n147 185
R932 VTAIL.n135 VTAIL.n134 185
R933 VTAIL.n133 VTAIL.n132 185
R934 VTAIL.n116 VTAIL.n115 185
R935 VTAIL.n127 VTAIL.n126 185
R936 VTAIL.n125 VTAIL.n124 185
R937 VTAIL.n120 VTAIL.n119 185
R938 VTAIL.n107 VTAIL.n106 185
R939 VTAIL.n105 VTAIL.n104 185
R940 VTAIL.n88 VTAIL.n87 185
R941 VTAIL.n99 VTAIL.n98 185
R942 VTAIL.n97 VTAIL.n96 185
R943 VTAIL.n92 VTAIL.n91 185
R944 VTAIL.n205 VTAIL.t0 147.672
R945 VTAIL.n9 VTAIL.t1 147.672
R946 VTAIL.n37 VTAIL.t5 147.672
R947 VTAIL.n65 VTAIL.t6 147.672
R948 VTAIL.n177 VTAIL.t4 147.672
R949 VTAIL.n149 VTAIL.t7 147.672
R950 VTAIL.n121 VTAIL.t3 147.672
R951 VTAIL.n93 VTAIL.t2 147.672
R952 VTAIL.n209 VTAIL.n203 104.615
R953 VTAIL.n210 VTAIL.n209 104.615
R954 VTAIL.n210 VTAIL.n199 104.615
R955 VTAIL.n217 VTAIL.n199 104.615
R956 VTAIL.n218 VTAIL.n217 104.615
R957 VTAIL.n13 VTAIL.n7 104.615
R958 VTAIL.n14 VTAIL.n13 104.615
R959 VTAIL.n14 VTAIL.n3 104.615
R960 VTAIL.n21 VTAIL.n3 104.615
R961 VTAIL.n22 VTAIL.n21 104.615
R962 VTAIL.n41 VTAIL.n35 104.615
R963 VTAIL.n42 VTAIL.n41 104.615
R964 VTAIL.n42 VTAIL.n31 104.615
R965 VTAIL.n49 VTAIL.n31 104.615
R966 VTAIL.n50 VTAIL.n49 104.615
R967 VTAIL.n69 VTAIL.n63 104.615
R968 VTAIL.n70 VTAIL.n69 104.615
R969 VTAIL.n70 VTAIL.n59 104.615
R970 VTAIL.n77 VTAIL.n59 104.615
R971 VTAIL.n78 VTAIL.n77 104.615
R972 VTAIL.n190 VTAIL.n189 104.615
R973 VTAIL.n189 VTAIL.n171 104.615
R974 VTAIL.n182 VTAIL.n171 104.615
R975 VTAIL.n182 VTAIL.n181 104.615
R976 VTAIL.n181 VTAIL.n175 104.615
R977 VTAIL.n162 VTAIL.n161 104.615
R978 VTAIL.n161 VTAIL.n143 104.615
R979 VTAIL.n154 VTAIL.n143 104.615
R980 VTAIL.n154 VTAIL.n153 104.615
R981 VTAIL.n153 VTAIL.n147 104.615
R982 VTAIL.n134 VTAIL.n133 104.615
R983 VTAIL.n133 VTAIL.n115 104.615
R984 VTAIL.n126 VTAIL.n115 104.615
R985 VTAIL.n126 VTAIL.n125 104.615
R986 VTAIL.n125 VTAIL.n119 104.615
R987 VTAIL.n106 VTAIL.n105 104.615
R988 VTAIL.n105 VTAIL.n87 104.615
R989 VTAIL.n98 VTAIL.n87 104.615
R990 VTAIL.n98 VTAIL.n97 104.615
R991 VTAIL.n97 VTAIL.n91 104.615
R992 VTAIL.t0 VTAIL.n203 52.3082
R993 VTAIL.t1 VTAIL.n7 52.3082
R994 VTAIL.t5 VTAIL.n35 52.3082
R995 VTAIL.t6 VTAIL.n63 52.3082
R996 VTAIL.t4 VTAIL.n175 52.3082
R997 VTAIL.t7 VTAIL.n147 52.3082
R998 VTAIL.t3 VTAIL.n119 52.3082
R999 VTAIL.t2 VTAIL.n91 52.3082
R1000 VTAIL.n223 VTAIL.n222 33.155
R1001 VTAIL.n27 VTAIL.n26 33.155
R1002 VTAIL.n55 VTAIL.n54 33.155
R1003 VTAIL.n83 VTAIL.n82 33.155
R1004 VTAIL.n195 VTAIL.n194 33.155
R1005 VTAIL.n167 VTAIL.n166 33.155
R1006 VTAIL.n139 VTAIL.n138 33.155
R1007 VTAIL.n111 VTAIL.n110 33.155
R1008 VTAIL.n223 VTAIL.n195 18.3065
R1009 VTAIL.n111 VTAIL.n83 18.3065
R1010 VTAIL.n205 VTAIL.n204 15.6666
R1011 VTAIL.n9 VTAIL.n8 15.6666
R1012 VTAIL.n37 VTAIL.n36 15.6666
R1013 VTAIL.n65 VTAIL.n64 15.6666
R1014 VTAIL.n177 VTAIL.n176 15.6666
R1015 VTAIL.n149 VTAIL.n148 15.6666
R1016 VTAIL.n121 VTAIL.n120 15.6666
R1017 VTAIL.n93 VTAIL.n92 15.6666
R1018 VTAIL.n208 VTAIL.n207 12.8005
R1019 VTAIL.n12 VTAIL.n11 12.8005
R1020 VTAIL.n40 VTAIL.n39 12.8005
R1021 VTAIL.n68 VTAIL.n67 12.8005
R1022 VTAIL.n180 VTAIL.n179 12.8005
R1023 VTAIL.n152 VTAIL.n151 12.8005
R1024 VTAIL.n124 VTAIL.n123 12.8005
R1025 VTAIL.n96 VTAIL.n95 12.8005
R1026 VTAIL.n211 VTAIL.n202 12.0247
R1027 VTAIL.n15 VTAIL.n6 12.0247
R1028 VTAIL.n43 VTAIL.n34 12.0247
R1029 VTAIL.n71 VTAIL.n62 12.0247
R1030 VTAIL.n183 VTAIL.n174 12.0247
R1031 VTAIL.n155 VTAIL.n146 12.0247
R1032 VTAIL.n127 VTAIL.n118 12.0247
R1033 VTAIL.n99 VTAIL.n90 12.0247
R1034 VTAIL.n212 VTAIL.n200 11.249
R1035 VTAIL.n16 VTAIL.n4 11.249
R1036 VTAIL.n44 VTAIL.n32 11.249
R1037 VTAIL.n72 VTAIL.n60 11.249
R1038 VTAIL.n184 VTAIL.n172 11.249
R1039 VTAIL.n156 VTAIL.n144 11.249
R1040 VTAIL.n128 VTAIL.n116 11.249
R1041 VTAIL.n100 VTAIL.n88 11.249
R1042 VTAIL.n216 VTAIL.n215 10.4732
R1043 VTAIL.n20 VTAIL.n19 10.4732
R1044 VTAIL.n48 VTAIL.n47 10.4732
R1045 VTAIL.n76 VTAIL.n75 10.4732
R1046 VTAIL.n188 VTAIL.n187 10.4732
R1047 VTAIL.n160 VTAIL.n159 10.4732
R1048 VTAIL.n132 VTAIL.n131 10.4732
R1049 VTAIL.n104 VTAIL.n103 10.4732
R1050 VTAIL.n219 VTAIL.n198 9.69747
R1051 VTAIL.n23 VTAIL.n2 9.69747
R1052 VTAIL.n51 VTAIL.n30 9.69747
R1053 VTAIL.n79 VTAIL.n58 9.69747
R1054 VTAIL.n191 VTAIL.n170 9.69747
R1055 VTAIL.n163 VTAIL.n142 9.69747
R1056 VTAIL.n135 VTAIL.n114 9.69747
R1057 VTAIL.n107 VTAIL.n86 9.69747
R1058 VTAIL.n222 VTAIL.n221 9.45567
R1059 VTAIL.n26 VTAIL.n25 9.45567
R1060 VTAIL.n54 VTAIL.n53 9.45567
R1061 VTAIL.n82 VTAIL.n81 9.45567
R1062 VTAIL.n194 VTAIL.n193 9.45567
R1063 VTAIL.n166 VTAIL.n165 9.45567
R1064 VTAIL.n138 VTAIL.n137 9.45567
R1065 VTAIL.n110 VTAIL.n109 9.45567
R1066 VTAIL.n221 VTAIL.n220 9.3005
R1067 VTAIL.n198 VTAIL.n197 9.3005
R1068 VTAIL.n215 VTAIL.n214 9.3005
R1069 VTAIL.n213 VTAIL.n212 9.3005
R1070 VTAIL.n202 VTAIL.n201 9.3005
R1071 VTAIL.n207 VTAIL.n206 9.3005
R1072 VTAIL.n25 VTAIL.n24 9.3005
R1073 VTAIL.n2 VTAIL.n1 9.3005
R1074 VTAIL.n19 VTAIL.n18 9.3005
R1075 VTAIL.n17 VTAIL.n16 9.3005
R1076 VTAIL.n6 VTAIL.n5 9.3005
R1077 VTAIL.n11 VTAIL.n10 9.3005
R1078 VTAIL.n53 VTAIL.n52 9.3005
R1079 VTAIL.n30 VTAIL.n29 9.3005
R1080 VTAIL.n47 VTAIL.n46 9.3005
R1081 VTAIL.n45 VTAIL.n44 9.3005
R1082 VTAIL.n34 VTAIL.n33 9.3005
R1083 VTAIL.n39 VTAIL.n38 9.3005
R1084 VTAIL.n81 VTAIL.n80 9.3005
R1085 VTAIL.n58 VTAIL.n57 9.3005
R1086 VTAIL.n75 VTAIL.n74 9.3005
R1087 VTAIL.n73 VTAIL.n72 9.3005
R1088 VTAIL.n62 VTAIL.n61 9.3005
R1089 VTAIL.n67 VTAIL.n66 9.3005
R1090 VTAIL.n193 VTAIL.n192 9.3005
R1091 VTAIL.n170 VTAIL.n169 9.3005
R1092 VTAIL.n187 VTAIL.n186 9.3005
R1093 VTAIL.n185 VTAIL.n184 9.3005
R1094 VTAIL.n174 VTAIL.n173 9.3005
R1095 VTAIL.n179 VTAIL.n178 9.3005
R1096 VTAIL.n165 VTAIL.n164 9.3005
R1097 VTAIL.n142 VTAIL.n141 9.3005
R1098 VTAIL.n159 VTAIL.n158 9.3005
R1099 VTAIL.n157 VTAIL.n156 9.3005
R1100 VTAIL.n146 VTAIL.n145 9.3005
R1101 VTAIL.n151 VTAIL.n150 9.3005
R1102 VTAIL.n137 VTAIL.n136 9.3005
R1103 VTAIL.n114 VTAIL.n113 9.3005
R1104 VTAIL.n131 VTAIL.n130 9.3005
R1105 VTAIL.n129 VTAIL.n128 9.3005
R1106 VTAIL.n118 VTAIL.n117 9.3005
R1107 VTAIL.n123 VTAIL.n122 9.3005
R1108 VTAIL.n109 VTAIL.n108 9.3005
R1109 VTAIL.n86 VTAIL.n85 9.3005
R1110 VTAIL.n103 VTAIL.n102 9.3005
R1111 VTAIL.n101 VTAIL.n100 9.3005
R1112 VTAIL.n90 VTAIL.n89 9.3005
R1113 VTAIL.n95 VTAIL.n94 9.3005
R1114 VTAIL.n220 VTAIL.n196 8.92171
R1115 VTAIL.n24 VTAIL.n0 8.92171
R1116 VTAIL.n52 VTAIL.n28 8.92171
R1117 VTAIL.n80 VTAIL.n56 8.92171
R1118 VTAIL.n192 VTAIL.n168 8.92171
R1119 VTAIL.n164 VTAIL.n140 8.92171
R1120 VTAIL.n136 VTAIL.n112 8.92171
R1121 VTAIL.n108 VTAIL.n84 8.92171
R1122 VTAIL.n222 VTAIL.n196 5.04292
R1123 VTAIL.n26 VTAIL.n0 5.04292
R1124 VTAIL.n54 VTAIL.n28 5.04292
R1125 VTAIL.n82 VTAIL.n56 5.04292
R1126 VTAIL.n194 VTAIL.n168 5.04292
R1127 VTAIL.n166 VTAIL.n140 5.04292
R1128 VTAIL.n138 VTAIL.n112 5.04292
R1129 VTAIL.n110 VTAIL.n84 5.04292
R1130 VTAIL.n206 VTAIL.n205 4.38687
R1131 VTAIL.n10 VTAIL.n9 4.38687
R1132 VTAIL.n38 VTAIL.n37 4.38687
R1133 VTAIL.n66 VTAIL.n65 4.38687
R1134 VTAIL.n178 VTAIL.n177 4.38687
R1135 VTAIL.n150 VTAIL.n149 4.38687
R1136 VTAIL.n122 VTAIL.n121 4.38687
R1137 VTAIL.n94 VTAIL.n93 4.38687
R1138 VTAIL.n220 VTAIL.n219 4.26717
R1139 VTAIL.n24 VTAIL.n23 4.26717
R1140 VTAIL.n52 VTAIL.n51 4.26717
R1141 VTAIL.n80 VTAIL.n79 4.26717
R1142 VTAIL.n192 VTAIL.n191 4.26717
R1143 VTAIL.n164 VTAIL.n163 4.26717
R1144 VTAIL.n136 VTAIL.n135 4.26717
R1145 VTAIL.n108 VTAIL.n107 4.26717
R1146 VTAIL.n216 VTAIL.n198 3.49141
R1147 VTAIL.n20 VTAIL.n2 3.49141
R1148 VTAIL.n48 VTAIL.n30 3.49141
R1149 VTAIL.n76 VTAIL.n58 3.49141
R1150 VTAIL.n188 VTAIL.n170 3.49141
R1151 VTAIL.n160 VTAIL.n142 3.49141
R1152 VTAIL.n132 VTAIL.n114 3.49141
R1153 VTAIL.n104 VTAIL.n86 3.49141
R1154 VTAIL.n215 VTAIL.n200 2.71565
R1155 VTAIL.n19 VTAIL.n4 2.71565
R1156 VTAIL.n47 VTAIL.n32 2.71565
R1157 VTAIL.n75 VTAIL.n60 2.71565
R1158 VTAIL.n187 VTAIL.n172 2.71565
R1159 VTAIL.n159 VTAIL.n144 2.71565
R1160 VTAIL.n131 VTAIL.n116 2.71565
R1161 VTAIL.n103 VTAIL.n88 2.71565
R1162 VTAIL.n212 VTAIL.n211 1.93989
R1163 VTAIL.n16 VTAIL.n15 1.93989
R1164 VTAIL.n44 VTAIL.n43 1.93989
R1165 VTAIL.n72 VTAIL.n71 1.93989
R1166 VTAIL.n184 VTAIL.n183 1.93989
R1167 VTAIL.n156 VTAIL.n155 1.93989
R1168 VTAIL.n128 VTAIL.n127 1.93989
R1169 VTAIL.n100 VTAIL.n99 1.93989
R1170 VTAIL.n139 VTAIL.n111 1.34533
R1171 VTAIL.n195 VTAIL.n167 1.34533
R1172 VTAIL.n83 VTAIL.n55 1.34533
R1173 VTAIL.n208 VTAIL.n202 1.16414
R1174 VTAIL.n12 VTAIL.n6 1.16414
R1175 VTAIL.n40 VTAIL.n34 1.16414
R1176 VTAIL.n68 VTAIL.n62 1.16414
R1177 VTAIL.n180 VTAIL.n174 1.16414
R1178 VTAIL.n152 VTAIL.n146 1.16414
R1179 VTAIL.n124 VTAIL.n118 1.16414
R1180 VTAIL.n96 VTAIL.n90 1.16414
R1181 VTAIL VTAIL.n27 0.731103
R1182 VTAIL VTAIL.n223 0.614724
R1183 VTAIL.n167 VTAIL.n139 0.470328
R1184 VTAIL.n55 VTAIL.n27 0.470328
R1185 VTAIL.n207 VTAIL.n204 0.388379
R1186 VTAIL.n11 VTAIL.n8 0.388379
R1187 VTAIL.n39 VTAIL.n36 0.388379
R1188 VTAIL.n67 VTAIL.n64 0.388379
R1189 VTAIL.n179 VTAIL.n176 0.388379
R1190 VTAIL.n151 VTAIL.n148 0.388379
R1191 VTAIL.n123 VTAIL.n120 0.388379
R1192 VTAIL.n95 VTAIL.n92 0.388379
R1193 VTAIL.n206 VTAIL.n201 0.155672
R1194 VTAIL.n213 VTAIL.n201 0.155672
R1195 VTAIL.n214 VTAIL.n213 0.155672
R1196 VTAIL.n214 VTAIL.n197 0.155672
R1197 VTAIL.n221 VTAIL.n197 0.155672
R1198 VTAIL.n10 VTAIL.n5 0.155672
R1199 VTAIL.n17 VTAIL.n5 0.155672
R1200 VTAIL.n18 VTAIL.n17 0.155672
R1201 VTAIL.n18 VTAIL.n1 0.155672
R1202 VTAIL.n25 VTAIL.n1 0.155672
R1203 VTAIL.n38 VTAIL.n33 0.155672
R1204 VTAIL.n45 VTAIL.n33 0.155672
R1205 VTAIL.n46 VTAIL.n45 0.155672
R1206 VTAIL.n46 VTAIL.n29 0.155672
R1207 VTAIL.n53 VTAIL.n29 0.155672
R1208 VTAIL.n66 VTAIL.n61 0.155672
R1209 VTAIL.n73 VTAIL.n61 0.155672
R1210 VTAIL.n74 VTAIL.n73 0.155672
R1211 VTAIL.n74 VTAIL.n57 0.155672
R1212 VTAIL.n81 VTAIL.n57 0.155672
R1213 VTAIL.n193 VTAIL.n169 0.155672
R1214 VTAIL.n186 VTAIL.n169 0.155672
R1215 VTAIL.n186 VTAIL.n185 0.155672
R1216 VTAIL.n185 VTAIL.n173 0.155672
R1217 VTAIL.n178 VTAIL.n173 0.155672
R1218 VTAIL.n165 VTAIL.n141 0.155672
R1219 VTAIL.n158 VTAIL.n141 0.155672
R1220 VTAIL.n158 VTAIL.n157 0.155672
R1221 VTAIL.n157 VTAIL.n145 0.155672
R1222 VTAIL.n150 VTAIL.n145 0.155672
R1223 VTAIL.n137 VTAIL.n113 0.155672
R1224 VTAIL.n130 VTAIL.n113 0.155672
R1225 VTAIL.n130 VTAIL.n129 0.155672
R1226 VTAIL.n129 VTAIL.n117 0.155672
R1227 VTAIL.n122 VTAIL.n117 0.155672
R1228 VTAIL.n109 VTAIL.n85 0.155672
R1229 VTAIL.n102 VTAIL.n85 0.155672
R1230 VTAIL.n102 VTAIL.n101 0.155672
R1231 VTAIL.n101 VTAIL.n89 0.155672
R1232 VTAIL.n94 VTAIL.n89 0.155672
R1233 VDD1 VDD1.n1 102.493
R1234 VDD1 VDD1.n0 69.683
R1235 VDD1.n0 VDD1.t0 3.71532
R1236 VDD1.n0 VDD1.t3 3.71532
R1237 VDD1.n1 VDD1.t2 3.71532
R1238 VDD1.n1 VDD1.t1 3.71532
R1239 VN.n0 VN.t2 140.919
R1240 VN.n1 VN.t1 140.919
R1241 VN.n0 VN.t0 140.698
R1242 VN.n1 VN.t3 140.698
R1243 VN VN.n1 55.6697
R1244 VN VN.n0 18.3553
R1245 VDD2.n2 VDD2.n0 101.969
R1246 VDD2.n2 VDD2.n1 69.6248
R1247 VDD2.n1 VDD2.t0 3.71532
R1248 VDD2.n1 VDD2.t2 3.71532
R1249 VDD2.n0 VDD2.t1 3.71532
R1250 VDD2.n0 VDD2.t3 3.71532
R1251 VDD2 VDD2.n2 0.0586897
C0 VDD2 VDD1 0.691651f
C1 VN VTAIL 1.96017f
C2 VP VTAIL 1.97428f
C3 VDD2 VN 1.92083f
C4 VDD2 VP 0.310844f
C5 VDD2 VTAIL 3.57616f
C6 VN VDD1 0.147575f
C7 VP VDD1 2.07979f
C8 VN VP 3.97004f
C9 VDD1 VTAIL 3.53114f
C10 VDD2 B 2.425495f
C11 VDD1 B 5.43062f
C12 VTAIL B 5.14135f
C13 VN B 6.67091f
C14 VP B 5.475414f
C15 VDD2.t1 B 0.074685f
C16 VDD2.t3 B 0.074685f
C17 VDD2.n0 B 0.853927f
C18 VDD2.t0 B 0.074685f
C19 VDD2.t2 B 0.074685f
C20 VDD2.n1 B 0.613643f
C21 VDD2.n2 B 1.75304f
C22 VN.t2 B 0.420088f
C23 VN.t0 B 0.419727f
C24 VN.n0 B 0.345079f
C25 VN.t1 B 0.420088f
C26 VN.t3 B 0.419727f
C27 VN.n1 B 0.884616f
C28 VDD1.t0 B 0.114101f
C29 VDD1.t3 B 0.114101f
C30 VDD1.n0 B 0.937794f
C31 VDD1.t2 B 0.114101f
C32 VDD1.t1 B 0.114101f
C33 VDD1.n1 B 1.32641f
C34 VTAIL.n0 B 0.016893f
C35 VTAIL.n1 B 0.011961f
C36 VTAIL.n2 B 0.006427f
C37 VTAIL.n3 B 0.015191f
C38 VTAIL.n4 B 0.006805f
C39 VTAIL.n5 B 0.011961f
C40 VTAIL.n6 B 0.006427f
C41 VTAIL.n7 B 0.011394f
C42 VTAIL.n8 B 0.008972f
C43 VTAIL.t1 B 0.024818f
C44 VTAIL.n9 B 0.049338f
C45 VTAIL.n10 B 0.24762f
C46 VTAIL.n11 B 0.006427f
C47 VTAIL.n12 B 0.006805f
C48 VTAIL.n13 B 0.015191f
C49 VTAIL.n14 B 0.015191f
C50 VTAIL.n15 B 0.006805f
C51 VTAIL.n16 B 0.006427f
C52 VTAIL.n17 B 0.011961f
C53 VTAIL.n18 B 0.011961f
C54 VTAIL.n19 B 0.006427f
C55 VTAIL.n20 B 0.006805f
C56 VTAIL.n21 B 0.015191f
C57 VTAIL.n22 B 0.03303f
C58 VTAIL.n23 B 0.006805f
C59 VTAIL.n24 B 0.006427f
C60 VTAIL.n25 B 0.028464f
C61 VTAIL.n26 B 0.018521f
C62 VTAIL.n27 B 0.056941f
C63 VTAIL.n28 B 0.016893f
C64 VTAIL.n29 B 0.011961f
C65 VTAIL.n30 B 0.006427f
C66 VTAIL.n31 B 0.015191f
C67 VTAIL.n32 B 0.006805f
C68 VTAIL.n33 B 0.011961f
C69 VTAIL.n34 B 0.006427f
C70 VTAIL.n35 B 0.011394f
C71 VTAIL.n36 B 0.008972f
C72 VTAIL.t5 B 0.024818f
C73 VTAIL.n37 B 0.049338f
C74 VTAIL.n38 B 0.24762f
C75 VTAIL.n39 B 0.006427f
C76 VTAIL.n40 B 0.006805f
C77 VTAIL.n41 B 0.015191f
C78 VTAIL.n42 B 0.015191f
C79 VTAIL.n43 B 0.006805f
C80 VTAIL.n44 B 0.006427f
C81 VTAIL.n45 B 0.011961f
C82 VTAIL.n46 B 0.011961f
C83 VTAIL.n47 B 0.006427f
C84 VTAIL.n48 B 0.006805f
C85 VTAIL.n49 B 0.015191f
C86 VTAIL.n50 B 0.03303f
C87 VTAIL.n51 B 0.006805f
C88 VTAIL.n52 B 0.006427f
C89 VTAIL.n53 B 0.028464f
C90 VTAIL.n54 B 0.018521f
C91 VTAIL.n55 B 0.080614f
C92 VTAIL.n56 B 0.016893f
C93 VTAIL.n57 B 0.011961f
C94 VTAIL.n58 B 0.006427f
C95 VTAIL.n59 B 0.015191f
C96 VTAIL.n60 B 0.006805f
C97 VTAIL.n61 B 0.011961f
C98 VTAIL.n62 B 0.006427f
C99 VTAIL.n63 B 0.011394f
C100 VTAIL.n64 B 0.008972f
C101 VTAIL.t6 B 0.024818f
C102 VTAIL.n65 B 0.049338f
C103 VTAIL.n66 B 0.24762f
C104 VTAIL.n67 B 0.006427f
C105 VTAIL.n68 B 0.006805f
C106 VTAIL.n69 B 0.015191f
C107 VTAIL.n70 B 0.015191f
C108 VTAIL.n71 B 0.006805f
C109 VTAIL.n72 B 0.006427f
C110 VTAIL.n73 B 0.011961f
C111 VTAIL.n74 B 0.011961f
C112 VTAIL.n75 B 0.006427f
C113 VTAIL.n76 B 0.006805f
C114 VTAIL.n77 B 0.015191f
C115 VTAIL.n78 B 0.03303f
C116 VTAIL.n79 B 0.006805f
C117 VTAIL.n80 B 0.006427f
C118 VTAIL.n81 B 0.028464f
C119 VTAIL.n82 B 0.018521f
C120 VTAIL.n83 B 0.453894f
C121 VTAIL.n84 B 0.016893f
C122 VTAIL.n85 B 0.011961f
C123 VTAIL.n86 B 0.006427f
C124 VTAIL.n87 B 0.015191f
C125 VTAIL.n88 B 0.006805f
C126 VTAIL.n89 B 0.011961f
C127 VTAIL.n90 B 0.006427f
C128 VTAIL.n91 B 0.011394f
C129 VTAIL.n92 B 0.008972f
C130 VTAIL.t2 B 0.024818f
C131 VTAIL.n93 B 0.049338f
C132 VTAIL.n94 B 0.24762f
C133 VTAIL.n95 B 0.006427f
C134 VTAIL.n96 B 0.006805f
C135 VTAIL.n97 B 0.015191f
C136 VTAIL.n98 B 0.015191f
C137 VTAIL.n99 B 0.006805f
C138 VTAIL.n100 B 0.006427f
C139 VTAIL.n101 B 0.011961f
C140 VTAIL.n102 B 0.011961f
C141 VTAIL.n103 B 0.006427f
C142 VTAIL.n104 B 0.006805f
C143 VTAIL.n105 B 0.015191f
C144 VTAIL.n106 B 0.03303f
C145 VTAIL.n107 B 0.006805f
C146 VTAIL.n108 B 0.006427f
C147 VTAIL.n109 B 0.028464f
C148 VTAIL.n110 B 0.018521f
C149 VTAIL.n111 B 0.453894f
C150 VTAIL.n112 B 0.016893f
C151 VTAIL.n113 B 0.011961f
C152 VTAIL.n114 B 0.006427f
C153 VTAIL.n115 B 0.015191f
C154 VTAIL.n116 B 0.006805f
C155 VTAIL.n117 B 0.011961f
C156 VTAIL.n118 B 0.006427f
C157 VTAIL.n119 B 0.011394f
C158 VTAIL.n120 B 0.008972f
C159 VTAIL.t3 B 0.024818f
C160 VTAIL.n121 B 0.049338f
C161 VTAIL.n122 B 0.24762f
C162 VTAIL.n123 B 0.006427f
C163 VTAIL.n124 B 0.006805f
C164 VTAIL.n125 B 0.015191f
C165 VTAIL.n126 B 0.015191f
C166 VTAIL.n127 B 0.006805f
C167 VTAIL.n128 B 0.006427f
C168 VTAIL.n129 B 0.011961f
C169 VTAIL.n130 B 0.011961f
C170 VTAIL.n131 B 0.006427f
C171 VTAIL.n132 B 0.006805f
C172 VTAIL.n133 B 0.015191f
C173 VTAIL.n134 B 0.03303f
C174 VTAIL.n135 B 0.006805f
C175 VTAIL.n136 B 0.006427f
C176 VTAIL.n137 B 0.028464f
C177 VTAIL.n138 B 0.018521f
C178 VTAIL.n139 B 0.080614f
C179 VTAIL.n140 B 0.016893f
C180 VTAIL.n141 B 0.011961f
C181 VTAIL.n142 B 0.006427f
C182 VTAIL.n143 B 0.015191f
C183 VTAIL.n144 B 0.006805f
C184 VTAIL.n145 B 0.011961f
C185 VTAIL.n146 B 0.006427f
C186 VTAIL.n147 B 0.011394f
C187 VTAIL.n148 B 0.008972f
C188 VTAIL.t7 B 0.024818f
C189 VTAIL.n149 B 0.049338f
C190 VTAIL.n150 B 0.24762f
C191 VTAIL.n151 B 0.006427f
C192 VTAIL.n152 B 0.006805f
C193 VTAIL.n153 B 0.015191f
C194 VTAIL.n154 B 0.015191f
C195 VTAIL.n155 B 0.006805f
C196 VTAIL.n156 B 0.006427f
C197 VTAIL.n157 B 0.011961f
C198 VTAIL.n158 B 0.011961f
C199 VTAIL.n159 B 0.006427f
C200 VTAIL.n160 B 0.006805f
C201 VTAIL.n161 B 0.015191f
C202 VTAIL.n162 B 0.03303f
C203 VTAIL.n163 B 0.006805f
C204 VTAIL.n164 B 0.006427f
C205 VTAIL.n165 B 0.028464f
C206 VTAIL.n166 B 0.018521f
C207 VTAIL.n167 B 0.080614f
C208 VTAIL.n168 B 0.016893f
C209 VTAIL.n169 B 0.011961f
C210 VTAIL.n170 B 0.006427f
C211 VTAIL.n171 B 0.015191f
C212 VTAIL.n172 B 0.006805f
C213 VTAIL.n173 B 0.011961f
C214 VTAIL.n174 B 0.006427f
C215 VTAIL.n175 B 0.011394f
C216 VTAIL.n176 B 0.008972f
C217 VTAIL.t4 B 0.024818f
C218 VTAIL.n177 B 0.049338f
C219 VTAIL.n178 B 0.24762f
C220 VTAIL.n179 B 0.006427f
C221 VTAIL.n180 B 0.006805f
C222 VTAIL.n181 B 0.015191f
C223 VTAIL.n182 B 0.015191f
C224 VTAIL.n183 B 0.006805f
C225 VTAIL.n184 B 0.006427f
C226 VTAIL.n185 B 0.011961f
C227 VTAIL.n186 B 0.011961f
C228 VTAIL.n187 B 0.006427f
C229 VTAIL.n188 B 0.006805f
C230 VTAIL.n189 B 0.015191f
C231 VTAIL.n190 B 0.03303f
C232 VTAIL.n191 B 0.006805f
C233 VTAIL.n192 B 0.006427f
C234 VTAIL.n193 B 0.028464f
C235 VTAIL.n194 B 0.018521f
C236 VTAIL.n195 B 0.453894f
C237 VTAIL.n196 B 0.016893f
C238 VTAIL.n197 B 0.011961f
C239 VTAIL.n198 B 0.006427f
C240 VTAIL.n199 B 0.015191f
C241 VTAIL.n200 B 0.006805f
C242 VTAIL.n201 B 0.011961f
C243 VTAIL.n202 B 0.006427f
C244 VTAIL.n203 B 0.011394f
C245 VTAIL.n204 B 0.008972f
C246 VTAIL.t0 B 0.024818f
C247 VTAIL.n205 B 0.049338f
C248 VTAIL.n206 B 0.24762f
C249 VTAIL.n207 B 0.006427f
C250 VTAIL.n208 B 0.006805f
C251 VTAIL.n209 B 0.015191f
C252 VTAIL.n210 B 0.015191f
C253 VTAIL.n211 B 0.006805f
C254 VTAIL.n212 B 0.006427f
C255 VTAIL.n213 B 0.011961f
C256 VTAIL.n214 B 0.011961f
C257 VTAIL.n215 B 0.006427f
C258 VTAIL.n216 B 0.006805f
C259 VTAIL.n217 B 0.015191f
C260 VTAIL.n218 B 0.03303f
C261 VTAIL.n219 B 0.006805f
C262 VTAIL.n220 B 0.006427f
C263 VTAIL.n221 B 0.028464f
C264 VTAIL.n222 B 0.018521f
C265 VTAIL.n223 B 0.425736f
C266 VP.n0 B 0.032448f
C267 VP.t2 B 0.55888f
C268 VP.n1 B 0.051354f
C269 VP.t3 B 0.645425f
C270 VP.t0 B 0.644869f
C271 VP.n2 B 1.34196f
C272 VP.t1 B 0.55888f
C273 VP.n3 B 0.28583f
C274 VP.n4 B 1.50997f
C275 VP.n5 B 0.032448f
C276 VP.n6 B 0.032448f
C277 VP.n7 B 0.026231f
C278 VP.n8 B 0.051354f
C279 VP.n9 B 0.28583f
C280 VP.n10 B 0.028967f
.ends

