* NGSPICE file created from diff_pair_sample_0769.ext - technology: sky130A

.subckt diff_pair_sample_0769 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=0 ps=0 w=7.12 l=3.76
X1 VDD2.t9 VN.t0 VTAIL.t18 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X2 VTAIL.t17 VN.t1 VDD2.t8 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X3 VDD2.t7 VN.t2 VTAIL.t10 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=2.7768 ps=15.02 w=7.12 l=3.76
X4 VTAIL.t11 VN.t3 VDD2.t6 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X5 VTAIL.t19 VP.t0 VDD1.t9 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X6 VTAIL.t2 VP.t1 VDD1.t8 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X7 VDD1.t7 VP.t2 VTAIL.t0 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=1.1748 ps=7.45 w=7.12 l=3.76
X8 VDD2.t5 VN.t4 VTAIL.t9 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=1.1748 ps=7.45 w=7.12 l=3.76
X9 VDD1.t6 VP.t3 VTAIL.t1 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=1.1748 ps=7.45 w=7.12 l=3.76
X10 B.t8 B.t6 B.t7 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=0 ps=0 w=7.12 l=3.76
X11 VDD1.t5 VP.t4 VTAIL.t3 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X12 VDD2.t4 VN.t5 VTAIL.t12 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=1.1748 ps=7.45 w=7.12 l=3.76
X13 VDD2.t3 VN.t6 VTAIL.t16 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=2.7768 ps=15.02 w=7.12 l=3.76
X14 B.t5 B.t3 B.t4 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=0 ps=0 w=7.12 l=3.76
X15 VTAIL.t13 VN.t7 VDD2.t2 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X16 VDD1.t4 VP.t5 VTAIL.t6 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=2.7768 ps=15.02 w=7.12 l=3.76
X17 VDD2.t1 VN.t8 VTAIL.t14 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X18 VTAIL.t5 VP.t6 VDD1.t3 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X19 B.t2 B.t0 B.t1 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=2.7768 pd=15.02 as=0 ps=0 w=7.12 l=3.76
X20 VDD1.t2 VP.t7 VTAIL.t4 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=2.7768 ps=15.02 w=7.12 l=3.76
X21 VDD1.t1 VP.t8 VTAIL.t7 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X22 VTAIL.t15 VN.t9 VDD2.t0 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
X23 VTAIL.t8 VP.t9 VDD1.t0 w_n5878_n2392# sky130_fd_pr__pfet_01v8 ad=1.1748 pd=7.45 as=1.1748 ps=7.45 w=7.12 l=3.76
R0 B.n451 B.n160 585
R1 B.n450 B.n449 585
R2 B.n448 B.n161 585
R3 B.n447 B.n446 585
R4 B.n445 B.n162 585
R5 B.n444 B.n443 585
R6 B.n442 B.n163 585
R7 B.n441 B.n440 585
R8 B.n439 B.n164 585
R9 B.n438 B.n437 585
R10 B.n436 B.n165 585
R11 B.n435 B.n434 585
R12 B.n433 B.n166 585
R13 B.n432 B.n431 585
R14 B.n430 B.n167 585
R15 B.n429 B.n428 585
R16 B.n427 B.n168 585
R17 B.n426 B.n425 585
R18 B.n424 B.n169 585
R19 B.n423 B.n422 585
R20 B.n421 B.n170 585
R21 B.n420 B.n419 585
R22 B.n418 B.n171 585
R23 B.n417 B.n416 585
R24 B.n415 B.n172 585
R25 B.n414 B.n413 585
R26 B.n412 B.n173 585
R27 B.n411 B.n410 585
R28 B.n406 B.n174 585
R29 B.n405 B.n404 585
R30 B.n403 B.n175 585
R31 B.n402 B.n401 585
R32 B.n400 B.n176 585
R33 B.n399 B.n398 585
R34 B.n397 B.n177 585
R35 B.n396 B.n395 585
R36 B.n394 B.n178 585
R37 B.n392 B.n391 585
R38 B.n390 B.n181 585
R39 B.n389 B.n388 585
R40 B.n387 B.n182 585
R41 B.n386 B.n385 585
R42 B.n384 B.n183 585
R43 B.n383 B.n382 585
R44 B.n381 B.n184 585
R45 B.n380 B.n379 585
R46 B.n378 B.n185 585
R47 B.n377 B.n376 585
R48 B.n375 B.n186 585
R49 B.n374 B.n373 585
R50 B.n372 B.n187 585
R51 B.n371 B.n370 585
R52 B.n369 B.n188 585
R53 B.n368 B.n367 585
R54 B.n366 B.n189 585
R55 B.n365 B.n364 585
R56 B.n363 B.n190 585
R57 B.n362 B.n361 585
R58 B.n360 B.n191 585
R59 B.n359 B.n358 585
R60 B.n357 B.n192 585
R61 B.n356 B.n355 585
R62 B.n354 B.n193 585
R63 B.n353 B.n352 585
R64 B.n453 B.n452 585
R65 B.n454 B.n159 585
R66 B.n456 B.n455 585
R67 B.n457 B.n158 585
R68 B.n459 B.n458 585
R69 B.n460 B.n157 585
R70 B.n462 B.n461 585
R71 B.n463 B.n156 585
R72 B.n465 B.n464 585
R73 B.n466 B.n155 585
R74 B.n468 B.n467 585
R75 B.n469 B.n154 585
R76 B.n471 B.n470 585
R77 B.n472 B.n153 585
R78 B.n474 B.n473 585
R79 B.n475 B.n152 585
R80 B.n477 B.n476 585
R81 B.n478 B.n151 585
R82 B.n480 B.n479 585
R83 B.n481 B.n150 585
R84 B.n483 B.n482 585
R85 B.n484 B.n149 585
R86 B.n486 B.n485 585
R87 B.n487 B.n148 585
R88 B.n489 B.n488 585
R89 B.n490 B.n147 585
R90 B.n492 B.n491 585
R91 B.n493 B.n146 585
R92 B.n495 B.n494 585
R93 B.n496 B.n145 585
R94 B.n498 B.n497 585
R95 B.n499 B.n144 585
R96 B.n501 B.n500 585
R97 B.n502 B.n143 585
R98 B.n504 B.n503 585
R99 B.n505 B.n142 585
R100 B.n507 B.n506 585
R101 B.n508 B.n141 585
R102 B.n510 B.n509 585
R103 B.n511 B.n140 585
R104 B.n513 B.n512 585
R105 B.n514 B.n139 585
R106 B.n516 B.n515 585
R107 B.n517 B.n138 585
R108 B.n519 B.n518 585
R109 B.n520 B.n137 585
R110 B.n522 B.n521 585
R111 B.n523 B.n136 585
R112 B.n525 B.n524 585
R113 B.n526 B.n135 585
R114 B.n528 B.n527 585
R115 B.n529 B.n134 585
R116 B.n531 B.n530 585
R117 B.n532 B.n133 585
R118 B.n534 B.n533 585
R119 B.n535 B.n132 585
R120 B.n537 B.n536 585
R121 B.n538 B.n131 585
R122 B.n540 B.n539 585
R123 B.n541 B.n130 585
R124 B.n543 B.n542 585
R125 B.n544 B.n129 585
R126 B.n546 B.n545 585
R127 B.n547 B.n128 585
R128 B.n549 B.n548 585
R129 B.n550 B.n127 585
R130 B.n552 B.n551 585
R131 B.n553 B.n126 585
R132 B.n555 B.n554 585
R133 B.n556 B.n125 585
R134 B.n558 B.n557 585
R135 B.n559 B.n124 585
R136 B.n561 B.n560 585
R137 B.n562 B.n123 585
R138 B.n564 B.n563 585
R139 B.n565 B.n122 585
R140 B.n567 B.n566 585
R141 B.n568 B.n121 585
R142 B.n570 B.n569 585
R143 B.n571 B.n120 585
R144 B.n573 B.n572 585
R145 B.n574 B.n119 585
R146 B.n576 B.n575 585
R147 B.n577 B.n118 585
R148 B.n579 B.n578 585
R149 B.n580 B.n117 585
R150 B.n582 B.n581 585
R151 B.n583 B.n116 585
R152 B.n585 B.n584 585
R153 B.n586 B.n115 585
R154 B.n588 B.n587 585
R155 B.n589 B.n114 585
R156 B.n591 B.n590 585
R157 B.n592 B.n113 585
R158 B.n594 B.n593 585
R159 B.n595 B.n112 585
R160 B.n597 B.n596 585
R161 B.n598 B.n111 585
R162 B.n600 B.n599 585
R163 B.n601 B.n110 585
R164 B.n603 B.n602 585
R165 B.n604 B.n109 585
R166 B.n606 B.n605 585
R167 B.n607 B.n108 585
R168 B.n609 B.n608 585
R169 B.n610 B.n107 585
R170 B.n612 B.n611 585
R171 B.n613 B.n106 585
R172 B.n615 B.n614 585
R173 B.n616 B.n105 585
R174 B.n618 B.n617 585
R175 B.n619 B.n104 585
R176 B.n621 B.n620 585
R177 B.n622 B.n103 585
R178 B.n624 B.n623 585
R179 B.n625 B.n102 585
R180 B.n627 B.n626 585
R181 B.n628 B.n101 585
R182 B.n630 B.n629 585
R183 B.n631 B.n100 585
R184 B.n633 B.n632 585
R185 B.n634 B.n99 585
R186 B.n636 B.n635 585
R187 B.n637 B.n98 585
R188 B.n639 B.n638 585
R189 B.n640 B.n97 585
R190 B.n642 B.n641 585
R191 B.n643 B.n96 585
R192 B.n645 B.n644 585
R193 B.n646 B.n95 585
R194 B.n648 B.n647 585
R195 B.n649 B.n94 585
R196 B.n651 B.n650 585
R197 B.n652 B.n93 585
R198 B.n654 B.n653 585
R199 B.n655 B.n92 585
R200 B.n657 B.n656 585
R201 B.n658 B.n91 585
R202 B.n660 B.n659 585
R203 B.n661 B.n90 585
R204 B.n663 B.n662 585
R205 B.n664 B.n89 585
R206 B.n666 B.n665 585
R207 B.n667 B.n88 585
R208 B.n669 B.n668 585
R209 B.n670 B.n87 585
R210 B.n672 B.n671 585
R211 B.n673 B.n86 585
R212 B.n675 B.n674 585
R213 B.n676 B.n85 585
R214 B.n678 B.n677 585
R215 B.n679 B.n84 585
R216 B.n681 B.n680 585
R217 B.n682 B.n83 585
R218 B.n684 B.n683 585
R219 B.n685 B.n82 585
R220 B.n687 B.n686 585
R221 B.n688 B.n81 585
R222 B.n690 B.n689 585
R223 B.n691 B.n80 585
R224 B.n693 B.n692 585
R225 B.n694 B.n79 585
R226 B.n791 B.n42 585
R227 B.n790 B.n789 585
R228 B.n788 B.n43 585
R229 B.n787 B.n786 585
R230 B.n785 B.n44 585
R231 B.n784 B.n783 585
R232 B.n782 B.n45 585
R233 B.n781 B.n780 585
R234 B.n779 B.n46 585
R235 B.n778 B.n777 585
R236 B.n776 B.n47 585
R237 B.n775 B.n774 585
R238 B.n773 B.n48 585
R239 B.n772 B.n771 585
R240 B.n770 B.n49 585
R241 B.n769 B.n768 585
R242 B.n767 B.n50 585
R243 B.n766 B.n765 585
R244 B.n764 B.n51 585
R245 B.n763 B.n762 585
R246 B.n761 B.n52 585
R247 B.n760 B.n759 585
R248 B.n758 B.n53 585
R249 B.n757 B.n756 585
R250 B.n755 B.n54 585
R251 B.n754 B.n753 585
R252 B.n752 B.n55 585
R253 B.n750 B.n749 585
R254 B.n748 B.n58 585
R255 B.n747 B.n746 585
R256 B.n745 B.n59 585
R257 B.n744 B.n743 585
R258 B.n742 B.n60 585
R259 B.n741 B.n740 585
R260 B.n739 B.n61 585
R261 B.n738 B.n737 585
R262 B.n736 B.n62 585
R263 B.n735 B.n734 585
R264 B.n733 B.n63 585
R265 B.n732 B.n731 585
R266 B.n730 B.n67 585
R267 B.n729 B.n728 585
R268 B.n727 B.n68 585
R269 B.n726 B.n725 585
R270 B.n724 B.n69 585
R271 B.n723 B.n722 585
R272 B.n721 B.n70 585
R273 B.n720 B.n719 585
R274 B.n718 B.n71 585
R275 B.n717 B.n716 585
R276 B.n715 B.n72 585
R277 B.n714 B.n713 585
R278 B.n712 B.n73 585
R279 B.n711 B.n710 585
R280 B.n709 B.n74 585
R281 B.n708 B.n707 585
R282 B.n706 B.n75 585
R283 B.n705 B.n704 585
R284 B.n703 B.n76 585
R285 B.n702 B.n701 585
R286 B.n700 B.n77 585
R287 B.n699 B.n698 585
R288 B.n697 B.n78 585
R289 B.n696 B.n695 585
R290 B.n793 B.n792 585
R291 B.n794 B.n41 585
R292 B.n796 B.n795 585
R293 B.n797 B.n40 585
R294 B.n799 B.n798 585
R295 B.n800 B.n39 585
R296 B.n802 B.n801 585
R297 B.n803 B.n38 585
R298 B.n805 B.n804 585
R299 B.n806 B.n37 585
R300 B.n808 B.n807 585
R301 B.n809 B.n36 585
R302 B.n811 B.n810 585
R303 B.n812 B.n35 585
R304 B.n814 B.n813 585
R305 B.n815 B.n34 585
R306 B.n817 B.n816 585
R307 B.n818 B.n33 585
R308 B.n820 B.n819 585
R309 B.n821 B.n32 585
R310 B.n823 B.n822 585
R311 B.n824 B.n31 585
R312 B.n826 B.n825 585
R313 B.n827 B.n30 585
R314 B.n829 B.n828 585
R315 B.n830 B.n29 585
R316 B.n832 B.n831 585
R317 B.n833 B.n28 585
R318 B.n835 B.n834 585
R319 B.n836 B.n27 585
R320 B.n838 B.n837 585
R321 B.n839 B.n26 585
R322 B.n841 B.n840 585
R323 B.n842 B.n25 585
R324 B.n844 B.n843 585
R325 B.n845 B.n24 585
R326 B.n847 B.n846 585
R327 B.n848 B.n23 585
R328 B.n850 B.n849 585
R329 B.n851 B.n22 585
R330 B.n853 B.n852 585
R331 B.n854 B.n21 585
R332 B.n856 B.n855 585
R333 B.n857 B.n20 585
R334 B.n859 B.n858 585
R335 B.n860 B.n19 585
R336 B.n862 B.n861 585
R337 B.n863 B.n18 585
R338 B.n865 B.n864 585
R339 B.n866 B.n17 585
R340 B.n868 B.n867 585
R341 B.n869 B.n16 585
R342 B.n871 B.n870 585
R343 B.n872 B.n15 585
R344 B.n874 B.n873 585
R345 B.n875 B.n14 585
R346 B.n877 B.n876 585
R347 B.n878 B.n13 585
R348 B.n880 B.n879 585
R349 B.n881 B.n12 585
R350 B.n883 B.n882 585
R351 B.n884 B.n11 585
R352 B.n886 B.n885 585
R353 B.n887 B.n10 585
R354 B.n889 B.n888 585
R355 B.n890 B.n9 585
R356 B.n892 B.n891 585
R357 B.n893 B.n8 585
R358 B.n895 B.n894 585
R359 B.n896 B.n7 585
R360 B.n898 B.n897 585
R361 B.n899 B.n6 585
R362 B.n901 B.n900 585
R363 B.n902 B.n5 585
R364 B.n904 B.n903 585
R365 B.n905 B.n4 585
R366 B.n907 B.n906 585
R367 B.n908 B.n3 585
R368 B.n910 B.n909 585
R369 B.n911 B.n0 585
R370 B.n2 B.n1 585
R371 B.n234 B.n233 585
R372 B.n236 B.n235 585
R373 B.n237 B.n232 585
R374 B.n239 B.n238 585
R375 B.n240 B.n231 585
R376 B.n242 B.n241 585
R377 B.n243 B.n230 585
R378 B.n245 B.n244 585
R379 B.n246 B.n229 585
R380 B.n248 B.n247 585
R381 B.n249 B.n228 585
R382 B.n251 B.n250 585
R383 B.n252 B.n227 585
R384 B.n254 B.n253 585
R385 B.n255 B.n226 585
R386 B.n257 B.n256 585
R387 B.n258 B.n225 585
R388 B.n260 B.n259 585
R389 B.n261 B.n224 585
R390 B.n263 B.n262 585
R391 B.n264 B.n223 585
R392 B.n266 B.n265 585
R393 B.n267 B.n222 585
R394 B.n269 B.n268 585
R395 B.n270 B.n221 585
R396 B.n272 B.n271 585
R397 B.n273 B.n220 585
R398 B.n275 B.n274 585
R399 B.n276 B.n219 585
R400 B.n278 B.n277 585
R401 B.n279 B.n218 585
R402 B.n281 B.n280 585
R403 B.n282 B.n217 585
R404 B.n284 B.n283 585
R405 B.n285 B.n216 585
R406 B.n287 B.n286 585
R407 B.n288 B.n215 585
R408 B.n290 B.n289 585
R409 B.n291 B.n214 585
R410 B.n293 B.n292 585
R411 B.n294 B.n213 585
R412 B.n296 B.n295 585
R413 B.n297 B.n212 585
R414 B.n299 B.n298 585
R415 B.n300 B.n211 585
R416 B.n302 B.n301 585
R417 B.n303 B.n210 585
R418 B.n305 B.n304 585
R419 B.n306 B.n209 585
R420 B.n308 B.n307 585
R421 B.n309 B.n208 585
R422 B.n311 B.n310 585
R423 B.n312 B.n207 585
R424 B.n314 B.n313 585
R425 B.n315 B.n206 585
R426 B.n317 B.n316 585
R427 B.n318 B.n205 585
R428 B.n320 B.n319 585
R429 B.n321 B.n204 585
R430 B.n323 B.n322 585
R431 B.n324 B.n203 585
R432 B.n326 B.n325 585
R433 B.n327 B.n202 585
R434 B.n329 B.n328 585
R435 B.n330 B.n201 585
R436 B.n332 B.n331 585
R437 B.n333 B.n200 585
R438 B.n335 B.n334 585
R439 B.n336 B.n199 585
R440 B.n338 B.n337 585
R441 B.n339 B.n198 585
R442 B.n341 B.n340 585
R443 B.n342 B.n197 585
R444 B.n344 B.n343 585
R445 B.n345 B.n196 585
R446 B.n347 B.n346 585
R447 B.n348 B.n195 585
R448 B.n350 B.n349 585
R449 B.n351 B.n194 585
R450 B.n353 B.n194 473.281
R451 B.n453 B.n160 473.281
R452 B.n695 B.n694 473.281
R453 B.n792 B.n791 473.281
R454 B.n913 B.n912 256.663
R455 B.n179 B.t9 254.948
R456 B.n407 B.t0 254.948
R457 B.n64 B.t3 254.948
R458 B.n56 B.t6 254.948
R459 B.n912 B.n911 235.042
R460 B.n912 B.n2 235.042
R461 B.n407 B.t1 195.066
R462 B.n64 B.t5 195.066
R463 B.n179 B.t10 195.059
R464 B.n56 B.t8 195.059
R465 B.n354 B.n353 163.367
R466 B.n355 B.n354 163.367
R467 B.n355 B.n192 163.367
R468 B.n359 B.n192 163.367
R469 B.n360 B.n359 163.367
R470 B.n361 B.n360 163.367
R471 B.n361 B.n190 163.367
R472 B.n365 B.n190 163.367
R473 B.n366 B.n365 163.367
R474 B.n367 B.n366 163.367
R475 B.n367 B.n188 163.367
R476 B.n371 B.n188 163.367
R477 B.n372 B.n371 163.367
R478 B.n373 B.n372 163.367
R479 B.n373 B.n186 163.367
R480 B.n377 B.n186 163.367
R481 B.n378 B.n377 163.367
R482 B.n379 B.n378 163.367
R483 B.n379 B.n184 163.367
R484 B.n383 B.n184 163.367
R485 B.n384 B.n383 163.367
R486 B.n385 B.n384 163.367
R487 B.n385 B.n182 163.367
R488 B.n389 B.n182 163.367
R489 B.n390 B.n389 163.367
R490 B.n391 B.n390 163.367
R491 B.n391 B.n178 163.367
R492 B.n396 B.n178 163.367
R493 B.n397 B.n396 163.367
R494 B.n398 B.n397 163.367
R495 B.n398 B.n176 163.367
R496 B.n402 B.n176 163.367
R497 B.n403 B.n402 163.367
R498 B.n404 B.n403 163.367
R499 B.n404 B.n174 163.367
R500 B.n411 B.n174 163.367
R501 B.n412 B.n411 163.367
R502 B.n413 B.n412 163.367
R503 B.n413 B.n172 163.367
R504 B.n417 B.n172 163.367
R505 B.n418 B.n417 163.367
R506 B.n419 B.n418 163.367
R507 B.n419 B.n170 163.367
R508 B.n423 B.n170 163.367
R509 B.n424 B.n423 163.367
R510 B.n425 B.n424 163.367
R511 B.n425 B.n168 163.367
R512 B.n429 B.n168 163.367
R513 B.n430 B.n429 163.367
R514 B.n431 B.n430 163.367
R515 B.n431 B.n166 163.367
R516 B.n435 B.n166 163.367
R517 B.n436 B.n435 163.367
R518 B.n437 B.n436 163.367
R519 B.n437 B.n164 163.367
R520 B.n441 B.n164 163.367
R521 B.n442 B.n441 163.367
R522 B.n443 B.n442 163.367
R523 B.n443 B.n162 163.367
R524 B.n447 B.n162 163.367
R525 B.n448 B.n447 163.367
R526 B.n449 B.n448 163.367
R527 B.n449 B.n160 163.367
R528 B.n694 B.n693 163.367
R529 B.n693 B.n80 163.367
R530 B.n689 B.n80 163.367
R531 B.n689 B.n688 163.367
R532 B.n688 B.n687 163.367
R533 B.n687 B.n82 163.367
R534 B.n683 B.n82 163.367
R535 B.n683 B.n682 163.367
R536 B.n682 B.n681 163.367
R537 B.n681 B.n84 163.367
R538 B.n677 B.n84 163.367
R539 B.n677 B.n676 163.367
R540 B.n676 B.n675 163.367
R541 B.n675 B.n86 163.367
R542 B.n671 B.n86 163.367
R543 B.n671 B.n670 163.367
R544 B.n670 B.n669 163.367
R545 B.n669 B.n88 163.367
R546 B.n665 B.n88 163.367
R547 B.n665 B.n664 163.367
R548 B.n664 B.n663 163.367
R549 B.n663 B.n90 163.367
R550 B.n659 B.n90 163.367
R551 B.n659 B.n658 163.367
R552 B.n658 B.n657 163.367
R553 B.n657 B.n92 163.367
R554 B.n653 B.n92 163.367
R555 B.n653 B.n652 163.367
R556 B.n652 B.n651 163.367
R557 B.n651 B.n94 163.367
R558 B.n647 B.n94 163.367
R559 B.n647 B.n646 163.367
R560 B.n646 B.n645 163.367
R561 B.n645 B.n96 163.367
R562 B.n641 B.n96 163.367
R563 B.n641 B.n640 163.367
R564 B.n640 B.n639 163.367
R565 B.n639 B.n98 163.367
R566 B.n635 B.n98 163.367
R567 B.n635 B.n634 163.367
R568 B.n634 B.n633 163.367
R569 B.n633 B.n100 163.367
R570 B.n629 B.n100 163.367
R571 B.n629 B.n628 163.367
R572 B.n628 B.n627 163.367
R573 B.n627 B.n102 163.367
R574 B.n623 B.n102 163.367
R575 B.n623 B.n622 163.367
R576 B.n622 B.n621 163.367
R577 B.n621 B.n104 163.367
R578 B.n617 B.n104 163.367
R579 B.n617 B.n616 163.367
R580 B.n616 B.n615 163.367
R581 B.n615 B.n106 163.367
R582 B.n611 B.n106 163.367
R583 B.n611 B.n610 163.367
R584 B.n610 B.n609 163.367
R585 B.n609 B.n108 163.367
R586 B.n605 B.n108 163.367
R587 B.n605 B.n604 163.367
R588 B.n604 B.n603 163.367
R589 B.n603 B.n110 163.367
R590 B.n599 B.n110 163.367
R591 B.n599 B.n598 163.367
R592 B.n598 B.n597 163.367
R593 B.n597 B.n112 163.367
R594 B.n593 B.n112 163.367
R595 B.n593 B.n592 163.367
R596 B.n592 B.n591 163.367
R597 B.n591 B.n114 163.367
R598 B.n587 B.n114 163.367
R599 B.n587 B.n586 163.367
R600 B.n586 B.n585 163.367
R601 B.n585 B.n116 163.367
R602 B.n581 B.n116 163.367
R603 B.n581 B.n580 163.367
R604 B.n580 B.n579 163.367
R605 B.n579 B.n118 163.367
R606 B.n575 B.n118 163.367
R607 B.n575 B.n574 163.367
R608 B.n574 B.n573 163.367
R609 B.n573 B.n120 163.367
R610 B.n569 B.n120 163.367
R611 B.n569 B.n568 163.367
R612 B.n568 B.n567 163.367
R613 B.n567 B.n122 163.367
R614 B.n563 B.n122 163.367
R615 B.n563 B.n562 163.367
R616 B.n562 B.n561 163.367
R617 B.n561 B.n124 163.367
R618 B.n557 B.n124 163.367
R619 B.n557 B.n556 163.367
R620 B.n556 B.n555 163.367
R621 B.n555 B.n126 163.367
R622 B.n551 B.n126 163.367
R623 B.n551 B.n550 163.367
R624 B.n550 B.n549 163.367
R625 B.n549 B.n128 163.367
R626 B.n545 B.n128 163.367
R627 B.n545 B.n544 163.367
R628 B.n544 B.n543 163.367
R629 B.n543 B.n130 163.367
R630 B.n539 B.n130 163.367
R631 B.n539 B.n538 163.367
R632 B.n538 B.n537 163.367
R633 B.n537 B.n132 163.367
R634 B.n533 B.n132 163.367
R635 B.n533 B.n532 163.367
R636 B.n532 B.n531 163.367
R637 B.n531 B.n134 163.367
R638 B.n527 B.n134 163.367
R639 B.n527 B.n526 163.367
R640 B.n526 B.n525 163.367
R641 B.n525 B.n136 163.367
R642 B.n521 B.n136 163.367
R643 B.n521 B.n520 163.367
R644 B.n520 B.n519 163.367
R645 B.n519 B.n138 163.367
R646 B.n515 B.n138 163.367
R647 B.n515 B.n514 163.367
R648 B.n514 B.n513 163.367
R649 B.n513 B.n140 163.367
R650 B.n509 B.n140 163.367
R651 B.n509 B.n508 163.367
R652 B.n508 B.n507 163.367
R653 B.n507 B.n142 163.367
R654 B.n503 B.n142 163.367
R655 B.n503 B.n502 163.367
R656 B.n502 B.n501 163.367
R657 B.n501 B.n144 163.367
R658 B.n497 B.n144 163.367
R659 B.n497 B.n496 163.367
R660 B.n496 B.n495 163.367
R661 B.n495 B.n146 163.367
R662 B.n491 B.n146 163.367
R663 B.n491 B.n490 163.367
R664 B.n490 B.n489 163.367
R665 B.n489 B.n148 163.367
R666 B.n485 B.n148 163.367
R667 B.n485 B.n484 163.367
R668 B.n484 B.n483 163.367
R669 B.n483 B.n150 163.367
R670 B.n479 B.n150 163.367
R671 B.n479 B.n478 163.367
R672 B.n478 B.n477 163.367
R673 B.n477 B.n152 163.367
R674 B.n473 B.n152 163.367
R675 B.n473 B.n472 163.367
R676 B.n472 B.n471 163.367
R677 B.n471 B.n154 163.367
R678 B.n467 B.n154 163.367
R679 B.n467 B.n466 163.367
R680 B.n466 B.n465 163.367
R681 B.n465 B.n156 163.367
R682 B.n461 B.n156 163.367
R683 B.n461 B.n460 163.367
R684 B.n460 B.n459 163.367
R685 B.n459 B.n158 163.367
R686 B.n455 B.n158 163.367
R687 B.n455 B.n454 163.367
R688 B.n454 B.n453 163.367
R689 B.n791 B.n790 163.367
R690 B.n790 B.n43 163.367
R691 B.n786 B.n43 163.367
R692 B.n786 B.n785 163.367
R693 B.n785 B.n784 163.367
R694 B.n784 B.n45 163.367
R695 B.n780 B.n45 163.367
R696 B.n780 B.n779 163.367
R697 B.n779 B.n778 163.367
R698 B.n778 B.n47 163.367
R699 B.n774 B.n47 163.367
R700 B.n774 B.n773 163.367
R701 B.n773 B.n772 163.367
R702 B.n772 B.n49 163.367
R703 B.n768 B.n49 163.367
R704 B.n768 B.n767 163.367
R705 B.n767 B.n766 163.367
R706 B.n766 B.n51 163.367
R707 B.n762 B.n51 163.367
R708 B.n762 B.n761 163.367
R709 B.n761 B.n760 163.367
R710 B.n760 B.n53 163.367
R711 B.n756 B.n53 163.367
R712 B.n756 B.n755 163.367
R713 B.n755 B.n754 163.367
R714 B.n754 B.n55 163.367
R715 B.n749 B.n55 163.367
R716 B.n749 B.n748 163.367
R717 B.n748 B.n747 163.367
R718 B.n747 B.n59 163.367
R719 B.n743 B.n59 163.367
R720 B.n743 B.n742 163.367
R721 B.n742 B.n741 163.367
R722 B.n741 B.n61 163.367
R723 B.n737 B.n61 163.367
R724 B.n737 B.n736 163.367
R725 B.n736 B.n735 163.367
R726 B.n735 B.n63 163.367
R727 B.n731 B.n63 163.367
R728 B.n731 B.n730 163.367
R729 B.n730 B.n729 163.367
R730 B.n729 B.n68 163.367
R731 B.n725 B.n68 163.367
R732 B.n725 B.n724 163.367
R733 B.n724 B.n723 163.367
R734 B.n723 B.n70 163.367
R735 B.n719 B.n70 163.367
R736 B.n719 B.n718 163.367
R737 B.n718 B.n717 163.367
R738 B.n717 B.n72 163.367
R739 B.n713 B.n72 163.367
R740 B.n713 B.n712 163.367
R741 B.n712 B.n711 163.367
R742 B.n711 B.n74 163.367
R743 B.n707 B.n74 163.367
R744 B.n707 B.n706 163.367
R745 B.n706 B.n705 163.367
R746 B.n705 B.n76 163.367
R747 B.n701 B.n76 163.367
R748 B.n701 B.n700 163.367
R749 B.n700 B.n699 163.367
R750 B.n699 B.n78 163.367
R751 B.n695 B.n78 163.367
R752 B.n792 B.n41 163.367
R753 B.n796 B.n41 163.367
R754 B.n797 B.n796 163.367
R755 B.n798 B.n797 163.367
R756 B.n798 B.n39 163.367
R757 B.n802 B.n39 163.367
R758 B.n803 B.n802 163.367
R759 B.n804 B.n803 163.367
R760 B.n804 B.n37 163.367
R761 B.n808 B.n37 163.367
R762 B.n809 B.n808 163.367
R763 B.n810 B.n809 163.367
R764 B.n810 B.n35 163.367
R765 B.n814 B.n35 163.367
R766 B.n815 B.n814 163.367
R767 B.n816 B.n815 163.367
R768 B.n816 B.n33 163.367
R769 B.n820 B.n33 163.367
R770 B.n821 B.n820 163.367
R771 B.n822 B.n821 163.367
R772 B.n822 B.n31 163.367
R773 B.n826 B.n31 163.367
R774 B.n827 B.n826 163.367
R775 B.n828 B.n827 163.367
R776 B.n828 B.n29 163.367
R777 B.n832 B.n29 163.367
R778 B.n833 B.n832 163.367
R779 B.n834 B.n833 163.367
R780 B.n834 B.n27 163.367
R781 B.n838 B.n27 163.367
R782 B.n839 B.n838 163.367
R783 B.n840 B.n839 163.367
R784 B.n840 B.n25 163.367
R785 B.n844 B.n25 163.367
R786 B.n845 B.n844 163.367
R787 B.n846 B.n845 163.367
R788 B.n846 B.n23 163.367
R789 B.n850 B.n23 163.367
R790 B.n851 B.n850 163.367
R791 B.n852 B.n851 163.367
R792 B.n852 B.n21 163.367
R793 B.n856 B.n21 163.367
R794 B.n857 B.n856 163.367
R795 B.n858 B.n857 163.367
R796 B.n858 B.n19 163.367
R797 B.n862 B.n19 163.367
R798 B.n863 B.n862 163.367
R799 B.n864 B.n863 163.367
R800 B.n864 B.n17 163.367
R801 B.n868 B.n17 163.367
R802 B.n869 B.n868 163.367
R803 B.n870 B.n869 163.367
R804 B.n870 B.n15 163.367
R805 B.n874 B.n15 163.367
R806 B.n875 B.n874 163.367
R807 B.n876 B.n875 163.367
R808 B.n876 B.n13 163.367
R809 B.n880 B.n13 163.367
R810 B.n881 B.n880 163.367
R811 B.n882 B.n881 163.367
R812 B.n882 B.n11 163.367
R813 B.n886 B.n11 163.367
R814 B.n887 B.n886 163.367
R815 B.n888 B.n887 163.367
R816 B.n888 B.n9 163.367
R817 B.n892 B.n9 163.367
R818 B.n893 B.n892 163.367
R819 B.n894 B.n893 163.367
R820 B.n894 B.n7 163.367
R821 B.n898 B.n7 163.367
R822 B.n899 B.n898 163.367
R823 B.n900 B.n899 163.367
R824 B.n900 B.n5 163.367
R825 B.n904 B.n5 163.367
R826 B.n905 B.n904 163.367
R827 B.n906 B.n905 163.367
R828 B.n906 B.n3 163.367
R829 B.n910 B.n3 163.367
R830 B.n911 B.n910 163.367
R831 B.n234 B.n2 163.367
R832 B.n235 B.n234 163.367
R833 B.n235 B.n232 163.367
R834 B.n239 B.n232 163.367
R835 B.n240 B.n239 163.367
R836 B.n241 B.n240 163.367
R837 B.n241 B.n230 163.367
R838 B.n245 B.n230 163.367
R839 B.n246 B.n245 163.367
R840 B.n247 B.n246 163.367
R841 B.n247 B.n228 163.367
R842 B.n251 B.n228 163.367
R843 B.n252 B.n251 163.367
R844 B.n253 B.n252 163.367
R845 B.n253 B.n226 163.367
R846 B.n257 B.n226 163.367
R847 B.n258 B.n257 163.367
R848 B.n259 B.n258 163.367
R849 B.n259 B.n224 163.367
R850 B.n263 B.n224 163.367
R851 B.n264 B.n263 163.367
R852 B.n265 B.n264 163.367
R853 B.n265 B.n222 163.367
R854 B.n269 B.n222 163.367
R855 B.n270 B.n269 163.367
R856 B.n271 B.n270 163.367
R857 B.n271 B.n220 163.367
R858 B.n275 B.n220 163.367
R859 B.n276 B.n275 163.367
R860 B.n277 B.n276 163.367
R861 B.n277 B.n218 163.367
R862 B.n281 B.n218 163.367
R863 B.n282 B.n281 163.367
R864 B.n283 B.n282 163.367
R865 B.n283 B.n216 163.367
R866 B.n287 B.n216 163.367
R867 B.n288 B.n287 163.367
R868 B.n289 B.n288 163.367
R869 B.n289 B.n214 163.367
R870 B.n293 B.n214 163.367
R871 B.n294 B.n293 163.367
R872 B.n295 B.n294 163.367
R873 B.n295 B.n212 163.367
R874 B.n299 B.n212 163.367
R875 B.n300 B.n299 163.367
R876 B.n301 B.n300 163.367
R877 B.n301 B.n210 163.367
R878 B.n305 B.n210 163.367
R879 B.n306 B.n305 163.367
R880 B.n307 B.n306 163.367
R881 B.n307 B.n208 163.367
R882 B.n311 B.n208 163.367
R883 B.n312 B.n311 163.367
R884 B.n313 B.n312 163.367
R885 B.n313 B.n206 163.367
R886 B.n317 B.n206 163.367
R887 B.n318 B.n317 163.367
R888 B.n319 B.n318 163.367
R889 B.n319 B.n204 163.367
R890 B.n323 B.n204 163.367
R891 B.n324 B.n323 163.367
R892 B.n325 B.n324 163.367
R893 B.n325 B.n202 163.367
R894 B.n329 B.n202 163.367
R895 B.n330 B.n329 163.367
R896 B.n331 B.n330 163.367
R897 B.n331 B.n200 163.367
R898 B.n335 B.n200 163.367
R899 B.n336 B.n335 163.367
R900 B.n337 B.n336 163.367
R901 B.n337 B.n198 163.367
R902 B.n341 B.n198 163.367
R903 B.n342 B.n341 163.367
R904 B.n343 B.n342 163.367
R905 B.n343 B.n196 163.367
R906 B.n347 B.n196 163.367
R907 B.n348 B.n347 163.367
R908 B.n349 B.n348 163.367
R909 B.n349 B.n194 163.367
R910 B.n408 B.t2 115.745
R911 B.n65 B.t4 115.745
R912 B.n180 B.t11 115.737
R913 B.n57 B.t7 115.737
R914 B.n180 B.n179 79.3217
R915 B.n408 B.n407 79.3217
R916 B.n65 B.n64 79.3217
R917 B.n57 B.n56 79.3217
R918 B.n393 B.n180 59.5399
R919 B.n409 B.n408 59.5399
R920 B.n66 B.n65 59.5399
R921 B.n751 B.n57 59.5399
R922 B.n793 B.n42 30.7517
R923 B.n696 B.n79 30.7517
R924 B.n452 B.n451 30.7517
R925 B.n352 B.n351 30.7517
R926 B B.n913 18.0485
R927 B.n794 B.n793 10.6151
R928 B.n795 B.n794 10.6151
R929 B.n795 B.n40 10.6151
R930 B.n799 B.n40 10.6151
R931 B.n800 B.n799 10.6151
R932 B.n801 B.n800 10.6151
R933 B.n801 B.n38 10.6151
R934 B.n805 B.n38 10.6151
R935 B.n806 B.n805 10.6151
R936 B.n807 B.n806 10.6151
R937 B.n807 B.n36 10.6151
R938 B.n811 B.n36 10.6151
R939 B.n812 B.n811 10.6151
R940 B.n813 B.n812 10.6151
R941 B.n813 B.n34 10.6151
R942 B.n817 B.n34 10.6151
R943 B.n818 B.n817 10.6151
R944 B.n819 B.n818 10.6151
R945 B.n819 B.n32 10.6151
R946 B.n823 B.n32 10.6151
R947 B.n824 B.n823 10.6151
R948 B.n825 B.n824 10.6151
R949 B.n825 B.n30 10.6151
R950 B.n829 B.n30 10.6151
R951 B.n830 B.n829 10.6151
R952 B.n831 B.n830 10.6151
R953 B.n831 B.n28 10.6151
R954 B.n835 B.n28 10.6151
R955 B.n836 B.n835 10.6151
R956 B.n837 B.n836 10.6151
R957 B.n837 B.n26 10.6151
R958 B.n841 B.n26 10.6151
R959 B.n842 B.n841 10.6151
R960 B.n843 B.n842 10.6151
R961 B.n843 B.n24 10.6151
R962 B.n847 B.n24 10.6151
R963 B.n848 B.n847 10.6151
R964 B.n849 B.n848 10.6151
R965 B.n849 B.n22 10.6151
R966 B.n853 B.n22 10.6151
R967 B.n854 B.n853 10.6151
R968 B.n855 B.n854 10.6151
R969 B.n855 B.n20 10.6151
R970 B.n859 B.n20 10.6151
R971 B.n860 B.n859 10.6151
R972 B.n861 B.n860 10.6151
R973 B.n861 B.n18 10.6151
R974 B.n865 B.n18 10.6151
R975 B.n866 B.n865 10.6151
R976 B.n867 B.n866 10.6151
R977 B.n867 B.n16 10.6151
R978 B.n871 B.n16 10.6151
R979 B.n872 B.n871 10.6151
R980 B.n873 B.n872 10.6151
R981 B.n873 B.n14 10.6151
R982 B.n877 B.n14 10.6151
R983 B.n878 B.n877 10.6151
R984 B.n879 B.n878 10.6151
R985 B.n879 B.n12 10.6151
R986 B.n883 B.n12 10.6151
R987 B.n884 B.n883 10.6151
R988 B.n885 B.n884 10.6151
R989 B.n885 B.n10 10.6151
R990 B.n889 B.n10 10.6151
R991 B.n890 B.n889 10.6151
R992 B.n891 B.n890 10.6151
R993 B.n891 B.n8 10.6151
R994 B.n895 B.n8 10.6151
R995 B.n896 B.n895 10.6151
R996 B.n897 B.n896 10.6151
R997 B.n897 B.n6 10.6151
R998 B.n901 B.n6 10.6151
R999 B.n902 B.n901 10.6151
R1000 B.n903 B.n902 10.6151
R1001 B.n903 B.n4 10.6151
R1002 B.n907 B.n4 10.6151
R1003 B.n908 B.n907 10.6151
R1004 B.n909 B.n908 10.6151
R1005 B.n909 B.n0 10.6151
R1006 B.n789 B.n42 10.6151
R1007 B.n789 B.n788 10.6151
R1008 B.n788 B.n787 10.6151
R1009 B.n787 B.n44 10.6151
R1010 B.n783 B.n44 10.6151
R1011 B.n783 B.n782 10.6151
R1012 B.n782 B.n781 10.6151
R1013 B.n781 B.n46 10.6151
R1014 B.n777 B.n46 10.6151
R1015 B.n777 B.n776 10.6151
R1016 B.n776 B.n775 10.6151
R1017 B.n775 B.n48 10.6151
R1018 B.n771 B.n48 10.6151
R1019 B.n771 B.n770 10.6151
R1020 B.n770 B.n769 10.6151
R1021 B.n769 B.n50 10.6151
R1022 B.n765 B.n50 10.6151
R1023 B.n765 B.n764 10.6151
R1024 B.n764 B.n763 10.6151
R1025 B.n763 B.n52 10.6151
R1026 B.n759 B.n52 10.6151
R1027 B.n759 B.n758 10.6151
R1028 B.n758 B.n757 10.6151
R1029 B.n757 B.n54 10.6151
R1030 B.n753 B.n54 10.6151
R1031 B.n753 B.n752 10.6151
R1032 B.n750 B.n58 10.6151
R1033 B.n746 B.n58 10.6151
R1034 B.n746 B.n745 10.6151
R1035 B.n745 B.n744 10.6151
R1036 B.n744 B.n60 10.6151
R1037 B.n740 B.n60 10.6151
R1038 B.n740 B.n739 10.6151
R1039 B.n739 B.n738 10.6151
R1040 B.n738 B.n62 10.6151
R1041 B.n734 B.n733 10.6151
R1042 B.n733 B.n732 10.6151
R1043 B.n732 B.n67 10.6151
R1044 B.n728 B.n67 10.6151
R1045 B.n728 B.n727 10.6151
R1046 B.n727 B.n726 10.6151
R1047 B.n726 B.n69 10.6151
R1048 B.n722 B.n69 10.6151
R1049 B.n722 B.n721 10.6151
R1050 B.n721 B.n720 10.6151
R1051 B.n720 B.n71 10.6151
R1052 B.n716 B.n71 10.6151
R1053 B.n716 B.n715 10.6151
R1054 B.n715 B.n714 10.6151
R1055 B.n714 B.n73 10.6151
R1056 B.n710 B.n73 10.6151
R1057 B.n710 B.n709 10.6151
R1058 B.n709 B.n708 10.6151
R1059 B.n708 B.n75 10.6151
R1060 B.n704 B.n75 10.6151
R1061 B.n704 B.n703 10.6151
R1062 B.n703 B.n702 10.6151
R1063 B.n702 B.n77 10.6151
R1064 B.n698 B.n77 10.6151
R1065 B.n698 B.n697 10.6151
R1066 B.n697 B.n696 10.6151
R1067 B.n692 B.n79 10.6151
R1068 B.n692 B.n691 10.6151
R1069 B.n691 B.n690 10.6151
R1070 B.n690 B.n81 10.6151
R1071 B.n686 B.n81 10.6151
R1072 B.n686 B.n685 10.6151
R1073 B.n685 B.n684 10.6151
R1074 B.n684 B.n83 10.6151
R1075 B.n680 B.n83 10.6151
R1076 B.n680 B.n679 10.6151
R1077 B.n679 B.n678 10.6151
R1078 B.n678 B.n85 10.6151
R1079 B.n674 B.n85 10.6151
R1080 B.n674 B.n673 10.6151
R1081 B.n673 B.n672 10.6151
R1082 B.n672 B.n87 10.6151
R1083 B.n668 B.n87 10.6151
R1084 B.n668 B.n667 10.6151
R1085 B.n667 B.n666 10.6151
R1086 B.n666 B.n89 10.6151
R1087 B.n662 B.n89 10.6151
R1088 B.n662 B.n661 10.6151
R1089 B.n661 B.n660 10.6151
R1090 B.n660 B.n91 10.6151
R1091 B.n656 B.n91 10.6151
R1092 B.n656 B.n655 10.6151
R1093 B.n655 B.n654 10.6151
R1094 B.n654 B.n93 10.6151
R1095 B.n650 B.n93 10.6151
R1096 B.n650 B.n649 10.6151
R1097 B.n649 B.n648 10.6151
R1098 B.n648 B.n95 10.6151
R1099 B.n644 B.n95 10.6151
R1100 B.n644 B.n643 10.6151
R1101 B.n643 B.n642 10.6151
R1102 B.n642 B.n97 10.6151
R1103 B.n638 B.n97 10.6151
R1104 B.n638 B.n637 10.6151
R1105 B.n637 B.n636 10.6151
R1106 B.n636 B.n99 10.6151
R1107 B.n632 B.n99 10.6151
R1108 B.n632 B.n631 10.6151
R1109 B.n631 B.n630 10.6151
R1110 B.n630 B.n101 10.6151
R1111 B.n626 B.n101 10.6151
R1112 B.n626 B.n625 10.6151
R1113 B.n625 B.n624 10.6151
R1114 B.n624 B.n103 10.6151
R1115 B.n620 B.n103 10.6151
R1116 B.n620 B.n619 10.6151
R1117 B.n619 B.n618 10.6151
R1118 B.n618 B.n105 10.6151
R1119 B.n614 B.n105 10.6151
R1120 B.n614 B.n613 10.6151
R1121 B.n613 B.n612 10.6151
R1122 B.n612 B.n107 10.6151
R1123 B.n608 B.n107 10.6151
R1124 B.n608 B.n607 10.6151
R1125 B.n607 B.n606 10.6151
R1126 B.n606 B.n109 10.6151
R1127 B.n602 B.n109 10.6151
R1128 B.n602 B.n601 10.6151
R1129 B.n601 B.n600 10.6151
R1130 B.n600 B.n111 10.6151
R1131 B.n596 B.n111 10.6151
R1132 B.n596 B.n595 10.6151
R1133 B.n595 B.n594 10.6151
R1134 B.n594 B.n113 10.6151
R1135 B.n590 B.n113 10.6151
R1136 B.n590 B.n589 10.6151
R1137 B.n589 B.n588 10.6151
R1138 B.n588 B.n115 10.6151
R1139 B.n584 B.n115 10.6151
R1140 B.n584 B.n583 10.6151
R1141 B.n583 B.n582 10.6151
R1142 B.n582 B.n117 10.6151
R1143 B.n578 B.n117 10.6151
R1144 B.n578 B.n577 10.6151
R1145 B.n577 B.n576 10.6151
R1146 B.n576 B.n119 10.6151
R1147 B.n572 B.n119 10.6151
R1148 B.n572 B.n571 10.6151
R1149 B.n571 B.n570 10.6151
R1150 B.n570 B.n121 10.6151
R1151 B.n566 B.n121 10.6151
R1152 B.n566 B.n565 10.6151
R1153 B.n565 B.n564 10.6151
R1154 B.n564 B.n123 10.6151
R1155 B.n560 B.n123 10.6151
R1156 B.n560 B.n559 10.6151
R1157 B.n559 B.n558 10.6151
R1158 B.n558 B.n125 10.6151
R1159 B.n554 B.n125 10.6151
R1160 B.n554 B.n553 10.6151
R1161 B.n553 B.n552 10.6151
R1162 B.n552 B.n127 10.6151
R1163 B.n548 B.n127 10.6151
R1164 B.n548 B.n547 10.6151
R1165 B.n547 B.n546 10.6151
R1166 B.n546 B.n129 10.6151
R1167 B.n542 B.n129 10.6151
R1168 B.n542 B.n541 10.6151
R1169 B.n541 B.n540 10.6151
R1170 B.n540 B.n131 10.6151
R1171 B.n536 B.n131 10.6151
R1172 B.n536 B.n535 10.6151
R1173 B.n535 B.n534 10.6151
R1174 B.n534 B.n133 10.6151
R1175 B.n530 B.n133 10.6151
R1176 B.n530 B.n529 10.6151
R1177 B.n529 B.n528 10.6151
R1178 B.n528 B.n135 10.6151
R1179 B.n524 B.n135 10.6151
R1180 B.n524 B.n523 10.6151
R1181 B.n523 B.n522 10.6151
R1182 B.n522 B.n137 10.6151
R1183 B.n518 B.n137 10.6151
R1184 B.n518 B.n517 10.6151
R1185 B.n517 B.n516 10.6151
R1186 B.n516 B.n139 10.6151
R1187 B.n512 B.n139 10.6151
R1188 B.n512 B.n511 10.6151
R1189 B.n511 B.n510 10.6151
R1190 B.n510 B.n141 10.6151
R1191 B.n506 B.n141 10.6151
R1192 B.n506 B.n505 10.6151
R1193 B.n505 B.n504 10.6151
R1194 B.n504 B.n143 10.6151
R1195 B.n500 B.n143 10.6151
R1196 B.n500 B.n499 10.6151
R1197 B.n499 B.n498 10.6151
R1198 B.n498 B.n145 10.6151
R1199 B.n494 B.n145 10.6151
R1200 B.n494 B.n493 10.6151
R1201 B.n493 B.n492 10.6151
R1202 B.n492 B.n147 10.6151
R1203 B.n488 B.n147 10.6151
R1204 B.n488 B.n487 10.6151
R1205 B.n487 B.n486 10.6151
R1206 B.n486 B.n149 10.6151
R1207 B.n482 B.n149 10.6151
R1208 B.n482 B.n481 10.6151
R1209 B.n481 B.n480 10.6151
R1210 B.n480 B.n151 10.6151
R1211 B.n476 B.n151 10.6151
R1212 B.n476 B.n475 10.6151
R1213 B.n475 B.n474 10.6151
R1214 B.n474 B.n153 10.6151
R1215 B.n470 B.n153 10.6151
R1216 B.n470 B.n469 10.6151
R1217 B.n469 B.n468 10.6151
R1218 B.n468 B.n155 10.6151
R1219 B.n464 B.n155 10.6151
R1220 B.n464 B.n463 10.6151
R1221 B.n463 B.n462 10.6151
R1222 B.n462 B.n157 10.6151
R1223 B.n458 B.n157 10.6151
R1224 B.n458 B.n457 10.6151
R1225 B.n457 B.n456 10.6151
R1226 B.n456 B.n159 10.6151
R1227 B.n452 B.n159 10.6151
R1228 B.n233 B.n1 10.6151
R1229 B.n236 B.n233 10.6151
R1230 B.n237 B.n236 10.6151
R1231 B.n238 B.n237 10.6151
R1232 B.n238 B.n231 10.6151
R1233 B.n242 B.n231 10.6151
R1234 B.n243 B.n242 10.6151
R1235 B.n244 B.n243 10.6151
R1236 B.n244 B.n229 10.6151
R1237 B.n248 B.n229 10.6151
R1238 B.n249 B.n248 10.6151
R1239 B.n250 B.n249 10.6151
R1240 B.n250 B.n227 10.6151
R1241 B.n254 B.n227 10.6151
R1242 B.n255 B.n254 10.6151
R1243 B.n256 B.n255 10.6151
R1244 B.n256 B.n225 10.6151
R1245 B.n260 B.n225 10.6151
R1246 B.n261 B.n260 10.6151
R1247 B.n262 B.n261 10.6151
R1248 B.n262 B.n223 10.6151
R1249 B.n266 B.n223 10.6151
R1250 B.n267 B.n266 10.6151
R1251 B.n268 B.n267 10.6151
R1252 B.n268 B.n221 10.6151
R1253 B.n272 B.n221 10.6151
R1254 B.n273 B.n272 10.6151
R1255 B.n274 B.n273 10.6151
R1256 B.n274 B.n219 10.6151
R1257 B.n278 B.n219 10.6151
R1258 B.n279 B.n278 10.6151
R1259 B.n280 B.n279 10.6151
R1260 B.n280 B.n217 10.6151
R1261 B.n284 B.n217 10.6151
R1262 B.n285 B.n284 10.6151
R1263 B.n286 B.n285 10.6151
R1264 B.n286 B.n215 10.6151
R1265 B.n290 B.n215 10.6151
R1266 B.n291 B.n290 10.6151
R1267 B.n292 B.n291 10.6151
R1268 B.n292 B.n213 10.6151
R1269 B.n296 B.n213 10.6151
R1270 B.n297 B.n296 10.6151
R1271 B.n298 B.n297 10.6151
R1272 B.n298 B.n211 10.6151
R1273 B.n302 B.n211 10.6151
R1274 B.n303 B.n302 10.6151
R1275 B.n304 B.n303 10.6151
R1276 B.n304 B.n209 10.6151
R1277 B.n308 B.n209 10.6151
R1278 B.n309 B.n308 10.6151
R1279 B.n310 B.n309 10.6151
R1280 B.n310 B.n207 10.6151
R1281 B.n314 B.n207 10.6151
R1282 B.n315 B.n314 10.6151
R1283 B.n316 B.n315 10.6151
R1284 B.n316 B.n205 10.6151
R1285 B.n320 B.n205 10.6151
R1286 B.n321 B.n320 10.6151
R1287 B.n322 B.n321 10.6151
R1288 B.n322 B.n203 10.6151
R1289 B.n326 B.n203 10.6151
R1290 B.n327 B.n326 10.6151
R1291 B.n328 B.n327 10.6151
R1292 B.n328 B.n201 10.6151
R1293 B.n332 B.n201 10.6151
R1294 B.n333 B.n332 10.6151
R1295 B.n334 B.n333 10.6151
R1296 B.n334 B.n199 10.6151
R1297 B.n338 B.n199 10.6151
R1298 B.n339 B.n338 10.6151
R1299 B.n340 B.n339 10.6151
R1300 B.n340 B.n197 10.6151
R1301 B.n344 B.n197 10.6151
R1302 B.n345 B.n344 10.6151
R1303 B.n346 B.n345 10.6151
R1304 B.n346 B.n195 10.6151
R1305 B.n350 B.n195 10.6151
R1306 B.n351 B.n350 10.6151
R1307 B.n352 B.n193 10.6151
R1308 B.n356 B.n193 10.6151
R1309 B.n357 B.n356 10.6151
R1310 B.n358 B.n357 10.6151
R1311 B.n358 B.n191 10.6151
R1312 B.n362 B.n191 10.6151
R1313 B.n363 B.n362 10.6151
R1314 B.n364 B.n363 10.6151
R1315 B.n364 B.n189 10.6151
R1316 B.n368 B.n189 10.6151
R1317 B.n369 B.n368 10.6151
R1318 B.n370 B.n369 10.6151
R1319 B.n370 B.n187 10.6151
R1320 B.n374 B.n187 10.6151
R1321 B.n375 B.n374 10.6151
R1322 B.n376 B.n375 10.6151
R1323 B.n376 B.n185 10.6151
R1324 B.n380 B.n185 10.6151
R1325 B.n381 B.n380 10.6151
R1326 B.n382 B.n381 10.6151
R1327 B.n382 B.n183 10.6151
R1328 B.n386 B.n183 10.6151
R1329 B.n387 B.n386 10.6151
R1330 B.n388 B.n387 10.6151
R1331 B.n388 B.n181 10.6151
R1332 B.n392 B.n181 10.6151
R1333 B.n395 B.n394 10.6151
R1334 B.n395 B.n177 10.6151
R1335 B.n399 B.n177 10.6151
R1336 B.n400 B.n399 10.6151
R1337 B.n401 B.n400 10.6151
R1338 B.n401 B.n175 10.6151
R1339 B.n405 B.n175 10.6151
R1340 B.n406 B.n405 10.6151
R1341 B.n410 B.n406 10.6151
R1342 B.n414 B.n173 10.6151
R1343 B.n415 B.n414 10.6151
R1344 B.n416 B.n415 10.6151
R1345 B.n416 B.n171 10.6151
R1346 B.n420 B.n171 10.6151
R1347 B.n421 B.n420 10.6151
R1348 B.n422 B.n421 10.6151
R1349 B.n422 B.n169 10.6151
R1350 B.n426 B.n169 10.6151
R1351 B.n427 B.n426 10.6151
R1352 B.n428 B.n427 10.6151
R1353 B.n428 B.n167 10.6151
R1354 B.n432 B.n167 10.6151
R1355 B.n433 B.n432 10.6151
R1356 B.n434 B.n433 10.6151
R1357 B.n434 B.n165 10.6151
R1358 B.n438 B.n165 10.6151
R1359 B.n439 B.n438 10.6151
R1360 B.n440 B.n439 10.6151
R1361 B.n440 B.n163 10.6151
R1362 B.n444 B.n163 10.6151
R1363 B.n445 B.n444 10.6151
R1364 B.n446 B.n445 10.6151
R1365 B.n446 B.n161 10.6151
R1366 B.n450 B.n161 10.6151
R1367 B.n451 B.n450 10.6151
R1368 B.n752 B.n751 9.36635
R1369 B.n734 B.n66 9.36635
R1370 B.n393 B.n392 9.36635
R1371 B.n409 B.n173 9.36635
R1372 B.n913 B.n0 8.11757
R1373 B.n913 B.n1 8.11757
R1374 B.n751 B.n750 1.24928
R1375 B.n66 B.n62 1.24928
R1376 B.n394 B.n393 1.24928
R1377 B.n410 B.n409 1.24928
R1378 VN.n105 VN.n54 161.3
R1379 VN.n104 VN.n103 161.3
R1380 VN.n102 VN.n55 161.3
R1381 VN.n101 VN.n100 161.3
R1382 VN.n99 VN.n56 161.3
R1383 VN.n98 VN.n97 161.3
R1384 VN.n96 VN.n57 161.3
R1385 VN.n95 VN.n94 161.3
R1386 VN.n92 VN.n58 161.3
R1387 VN.n91 VN.n90 161.3
R1388 VN.n89 VN.n59 161.3
R1389 VN.n88 VN.n87 161.3
R1390 VN.n86 VN.n60 161.3
R1391 VN.n85 VN.n84 161.3
R1392 VN.n83 VN.n61 161.3
R1393 VN.n82 VN.n81 161.3
R1394 VN.n79 VN.n62 161.3
R1395 VN.n78 VN.n77 161.3
R1396 VN.n76 VN.n63 161.3
R1397 VN.n75 VN.n74 161.3
R1398 VN.n73 VN.n64 161.3
R1399 VN.n72 VN.n71 161.3
R1400 VN.n70 VN.n65 161.3
R1401 VN.n69 VN.n68 161.3
R1402 VN.n51 VN.n0 161.3
R1403 VN.n50 VN.n49 161.3
R1404 VN.n48 VN.n1 161.3
R1405 VN.n47 VN.n46 161.3
R1406 VN.n45 VN.n2 161.3
R1407 VN.n44 VN.n43 161.3
R1408 VN.n42 VN.n3 161.3
R1409 VN.n41 VN.n40 161.3
R1410 VN.n38 VN.n4 161.3
R1411 VN.n37 VN.n36 161.3
R1412 VN.n35 VN.n5 161.3
R1413 VN.n34 VN.n33 161.3
R1414 VN.n32 VN.n6 161.3
R1415 VN.n31 VN.n30 161.3
R1416 VN.n29 VN.n7 161.3
R1417 VN.n28 VN.n27 161.3
R1418 VN.n25 VN.n8 161.3
R1419 VN.n24 VN.n23 161.3
R1420 VN.n22 VN.n9 161.3
R1421 VN.n21 VN.n20 161.3
R1422 VN.n19 VN.n10 161.3
R1423 VN.n18 VN.n17 161.3
R1424 VN.n16 VN.n11 161.3
R1425 VN.n15 VN.n14 161.3
R1426 VN.n12 VN.t5 78.0002
R1427 VN.n66 VN.t6 78.0002
R1428 VN.n53 VN.n52 61.2309
R1429 VN.n107 VN.n106 61.2309
R1430 VN.n13 VN.n12 58.5323
R1431 VN.n67 VN.n66 58.5323
R1432 VN.n20 VN.n19 56.5617
R1433 VN.n33 VN.n32 56.5617
R1434 VN.n74 VN.n73 56.5617
R1435 VN.n87 VN.n86 56.5617
R1436 VN VN.n107 55.9627
R1437 VN.n46 VN.n45 51.7179
R1438 VN.n100 VN.n99 51.7179
R1439 VN.n13 VN.t1 45.6367
R1440 VN.n26 VN.t8 45.6367
R1441 VN.n39 VN.t9 45.6367
R1442 VN.n52 VN.t2 45.6367
R1443 VN.n67 VN.t3 45.6367
R1444 VN.n80 VN.t0 45.6367
R1445 VN.n93 VN.t7 45.6367
R1446 VN.n106 VN.t4 45.6367
R1447 VN.n46 VN.n1 29.4362
R1448 VN.n100 VN.n55 29.4362
R1449 VN.n14 VN.n11 24.5923
R1450 VN.n18 VN.n11 24.5923
R1451 VN.n19 VN.n18 24.5923
R1452 VN.n20 VN.n9 24.5923
R1453 VN.n24 VN.n9 24.5923
R1454 VN.n25 VN.n24 24.5923
R1455 VN.n27 VN.n7 24.5923
R1456 VN.n31 VN.n7 24.5923
R1457 VN.n32 VN.n31 24.5923
R1458 VN.n33 VN.n5 24.5923
R1459 VN.n37 VN.n5 24.5923
R1460 VN.n38 VN.n37 24.5923
R1461 VN.n40 VN.n3 24.5923
R1462 VN.n44 VN.n3 24.5923
R1463 VN.n45 VN.n44 24.5923
R1464 VN.n50 VN.n1 24.5923
R1465 VN.n51 VN.n50 24.5923
R1466 VN.n73 VN.n72 24.5923
R1467 VN.n72 VN.n65 24.5923
R1468 VN.n68 VN.n65 24.5923
R1469 VN.n86 VN.n85 24.5923
R1470 VN.n85 VN.n61 24.5923
R1471 VN.n81 VN.n61 24.5923
R1472 VN.n79 VN.n78 24.5923
R1473 VN.n78 VN.n63 24.5923
R1474 VN.n74 VN.n63 24.5923
R1475 VN.n99 VN.n98 24.5923
R1476 VN.n98 VN.n57 24.5923
R1477 VN.n94 VN.n57 24.5923
R1478 VN.n92 VN.n91 24.5923
R1479 VN.n91 VN.n59 24.5923
R1480 VN.n87 VN.n59 24.5923
R1481 VN.n105 VN.n104 24.5923
R1482 VN.n104 VN.n55 24.5923
R1483 VN.n52 VN.n51 21.1495
R1484 VN.n106 VN.n105 21.1495
R1485 VN.n14 VN.n13 16.7229
R1486 VN.n39 VN.n38 16.7229
R1487 VN.n68 VN.n67 16.7229
R1488 VN.n93 VN.n92 16.7229
R1489 VN.n26 VN.n25 12.2964
R1490 VN.n27 VN.n26 12.2964
R1491 VN.n81 VN.n80 12.2964
R1492 VN.n80 VN.n79 12.2964
R1493 VN.n40 VN.n39 7.86989
R1494 VN.n94 VN.n93 7.86989
R1495 VN.n69 VN.n66 2.63944
R1496 VN.n15 VN.n12 2.63944
R1497 VN.n107 VN.n54 0.417304
R1498 VN.n53 VN.n0 0.417304
R1499 VN VN.n53 0.394524
R1500 VN.n103 VN.n54 0.189894
R1501 VN.n103 VN.n102 0.189894
R1502 VN.n102 VN.n101 0.189894
R1503 VN.n101 VN.n56 0.189894
R1504 VN.n97 VN.n56 0.189894
R1505 VN.n97 VN.n96 0.189894
R1506 VN.n96 VN.n95 0.189894
R1507 VN.n95 VN.n58 0.189894
R1508 VN.n90 VN.n58 0.189894
R1509 VN.n90 VN.n89 0.189894
R1510 VN.n89 VN.n88 0.189894
R1511 VN.n88 VN.n60 0.189894
R1512 VN.n84 VN.n60 0.189894
R1513 VN.n84 VN.n83 0.189894
R1514 VN.n83 VN.n82 0.189894
R1515 VN.n82 VN.n62 0.189894
R1516 VN.n77 VN.n62 0.189894
R1517 VN.n77 VN.n76 0.189894
R1518 VN.n76 VN.n75 0.189894
R1519 VN.n75 VN.n64 0.189894
R1520 VN.n71 VN.n64 0.189894
R1521 VN.n71 VN.n70 0.189894
R1522 VN.n70 VN.n69 0.189894
R1523 VN.n16 VN.n15 0.189894
R1524 VN.n17 VN.n16 0.189894
R1525 VN.n17 VN.n10 0.189894
R1526 VN.n21 VN.n10 0.189894
R1527 VN.n22 VN.n21 0.189894
R1528 VN.n23 VN.n22 0.189894
R1529 VN.n23 VN.n8 0.189894
R1530 VN.n28 VN.n8 0.189894
R1531 VN.n29 VN.n28 0.189894
R1532 VN.n30 VN.n29 0.189894
R1533 VN.n30 VN.n6 0.189894
R1534 VN.n34 VN.n6 0.189894
R1535 VN.n35 VN.n34 0.189894
R1536 VN.n36 VN.n35 0.189894
R1537 VN.n36 VN.n4 0.189894
R1538 VN.n41 VN.n4 0.189894
R1539 VN.n42 VN.n41 0.189894
R1540 VN.n43 VN.n42 0.189894
R1541 VN.n43 VN.n2 0.189894
R1542 VN.n47 VN.n2 0.189894
R1543 VN.n48 VN.n47 0.189894
R1544 VN.n49 VN.n48 0.189894
R1545 VN.n49 VN.n0 0.189894
R1546 VTAIL.n11 VTAIL.t16 75.4284
R1547 VTAIL.n17 VTAIL.t10 75.4282
R1548 VTAIL.n2 VTAIL.t6 75.4282
R1549 VTAIL.n16 VTAIL.t4 75.4282
R1550 VTAIL.n15 VTAIL.n14 70.8631
R1551 VTAIL.n13 VTAIL.n12 70.8631
R1552 VTAIL.n10 VTAIL.n9 70.8631
R1553 VTAIL.n8 VTAIL.n7 70.8631
R1554 VTAIL.n19 VTAIL.n18 70.863
R1555 VTAIL.n1 VTAIL.n0 70.863
R1556 VTAIL.n4 VTAIL.n3 70.863
R1557 VTAIL.n6 VTAIL.n5 70.863
R1558 VTAIL.n8 VTAIL.n6 25.5565
R1559 VTAIL.n17 VTAIL.n16 22.0307
R1560 VTAIL.n18 VTAIL.t14 4.56581
R1561 VTAIL.n18 VTAIL.t15 4.56581
R1562 VTAIL.n0 VTAIL.t12 4.56581
R1563 VTAIL.n0 VTAIL.t17 4.56581
R1564 VTAIL.n3 VTAIL.t3 4.56581
R1565 VTAIL.n3 VTAIL.t8 4.56581
R1566 VTAIL.n5 VTAIL.t0 4.56581
R1567 VTAIL.n5 VTAIL.t5 4.56581
R1568 VTAIL.n14 VTAIL.t7 4.56581
R1569 VTAIL.n14 VTAIL.t19 4.56581
R1570 VTAIL.n12 VTAIL.t1 4.56581
R1571 VTAIL.n12 VTAIL.t2 4.56581
R1572 VTAIL.n9 VTAIL.t18 4.56581
R1573 VTAIL.n9 VTAIL.t11 4.56581
R1574 VTAIL.n7 VTAIL.t9 4.56581
R1575 VTAIL.n7 VTAIL.t13 4.56581
R1576 VTAIL.n10 VTAIL.n8 3.52636
R1577 VTAIL.n11 VTAIL.n10 3.52636
R1578 VTAIL.n15 VTAIL.n13 3.52636
R1579 VTAIL.n16 VTAIL.n15 3.52636
R1580 VTAIL.n6 VTAIL.n4 3.52636
R1581 VTAIL.n4 VTAIL.n2 3.52636
R1582 VTAIL.n19 VTAIL.n17 3.52636
R1583 VTAIL VTAIL.n1 2.70309
R1584 VTAIL.n13 VTAIL.n11 2.23326
R1585 VTAIL.n2 VTAIL.n1 2.23326
R1586 VTAIL VTAIL.n19 0.823776
R1587 VDD2.n1 VDD2.t4 95.6328
R1588 VDD2.n4 VDD2.t5 92.1072
R1589 VDD2.n3 VDD2.n2 90.1309
R1590 VDD2 VDD2.n7 90.1279
R1591 VDD2.n6 VDD2.n5 87.5419
R1592 VDD2.n1 VDD2.n0 87.5418
R1593 VDD2.n4 VDD2.n3 46.6011
R1594 VDD2.n7 VDD2.t6 4.56581
R1595 VDD2.n7 VDD2.t3 4.56581
R1596 VDD2.n5 VDD2.t2 4.56581
R1597 VDD2.n5 VDD2.t9 4.56581
R1598 VDD2.n2 VDD2.t0 4.56581
R1599 VDD2.n2 VDD2.t7 4.56581
R1600 VDD2.n0 VDD2.t8 4.56581
R1601 VDD2.n0 VDD2.t1 4.56581
R1602 VDD2.n6 VDD2.n4 3.52636
R1603 VDD2 VDD2.n6 0.940155
R1604 VDD2.n3 VDD2.n1 0.826619
R1605 VP.n31 VP.n30 161.3
R1606 VP.n32 VP.n27 161.3
R1607 VP.n34 VP.n33 161.3
R1608 VP.n35 VP.n26 161.3
R1609 VP.n37 VP.n36 161.3
R1610 VP.n38 VP.n25 161.3
R1611 VP.n40 VP.n39 161.3
R1612 VP.n41 VP.n24 161.3
R1613 VP.n44 VP.n43 161.3
R1614 VP.n45 VP.n23 161.3
R1615 VP.n47 VP.n46 161.3
R1616 VP.n48 VP.n22 161.3
R1617 VP.n50 VP.n49 161.3
R1618 VP.n51 VP.n21 161.3
R1619 VP.n53 VP.n52 161.3
R1620 VP.n54 VP.n20 161.3
R1621 VP.n57 VP.n56 161.3
R1622 VP.n58 VP.n19 161.3
R1623 VP.n60 VP.n59 161.3
R1624 VP.n61 VP.n18 161.3
R1625 VP.n63 VP.n62 161.3
R1626 VP.n64 VP.n17 161.3
R1627 VP.n66 VP.n65 161.3
R1628 VP.n67 VP.n16 161.3
R1629 VP.n122 VP.n0 161.3
R1630 VP.n121 VP.n120 161.3
R1631 VP.n119 VP.n1 161.3
R1632 VP.n118 VP.n117 161.3
R1633 VP.n116 VP.n2 161.3
R1634 VP.n115 VP.n114 161.3
R1635 VP.n113 VP.n3 161.3
R1636 VP.n112 VP.n111 161.3
R1637 VP.n109 VP.n4 161.3
R1638 VP.n108 VP.n107 161.3
R1639 VP.n106 VP.n5 161.3
R1640 VP.n105 VP.n104 161.3
R1641 VP.n103 VP.n6 161.3
R1642 VP.n102 VP.n101 161.3
R1643 VP.n100 VP.n7 161.3
R1644 VP.n99 VP.n98 161.3
R1645 VP.n96 VP.n8 161.3
R1646 VP.n95 VP.n94 161.3
R1647 VP.n93 VP.n9 161.3
R1648 VP.n92 VP.n91 161.3
R1649 VP.n90 VP.n10 161.3
R1650 VP.n89 VP.n88 161.3
R1651 VP.n87 VP.n11 161.3
R1652 VP.n86 VP.n85 161.3
R1653 VP.n83 VP.n12 161.3
R1654 VP.n82 VP.n81 161.3
R1655 VP.n80 VP.n13 161.3
R1656 VP.n79 VP.n78 161.3
R1657 VP.n77 VP.n14 161.3
R1658 VP.n76 VP.n75 161.3
R1659 VP.n74 VP.n15 161.3
R1660 VP.n73 VP.n72 161.3
R1661 VP.n28 VP.t3 77.9999
R1662 VP.n71 VP.n70 61.2309
R1663 VP.n124 VP.n123 61.2309
R1664 VP.n69 VP.n68 61.2309
R1665 VP.n29 VP.n28 58.5323
R1666 VP.n91 VP.n90 56.5617
R1667 VP.n104 VP.n103 56.5617
R1668 VP.n49 VP.n48 56.5617
R1669 VP.n36 VP.n35 56.5617
R1670 VP.n70 VP.n69 55.9249
R1671 VP.n78 VP.n77 51.7179
R1672 VP.n117 VP.n116 51.7179
R1673 VP.n62 VP.n61 51.7179
R1674 VP.n71 VP.t2 45.6367
R1675 VP.n84 VP.t6 45.6367
R1676 VP.n97 VP.t4 45.6367
R1677 VP.n110 VP.t9 45.6367
R1678 VP.n123 VP.t5 45.6367
R1679 VP.n68 VP.t7 45.6367
R1680 VP.n55 VP.t0 45.6367
R1681 VP.n42 VP.t8 45.6367
R1682 VP.n29 VP.t1 45.6367
R1683 VP.n77 VP.n76 29.4362
R1684 VP.n117 VP.n1 29.4362
R1685 VP.n62 VP.n17 29.4362
R1686 VP.n72 VP.n15 24.5923
R1687 VP.n76 VP.n15 24.5923
R1688 VP.n78 VP.n13 24.5923
R1689 VP.n82 VP.n13 24.5923
R1690 VP.n83 VP.n82 24.5923
R1691 VP.n85 VP.n11 24.5923
R1692 VP.n89 VP.n11 24.5923
R1693 VP.n90 VP.n89 24.5923
R1694 VP.n91 VP.n9 24.5923
R1695 VP.n95 VP.n9 24.5923
R1696 VP.n96 VP.n95 24.5923
R1697 VP.n98 VP.n7 24.5923
R1698 VP.n102 VP.n7 24.5923
R1699 VP.n103 VP.n102 24.5923
R1700 VP.n104 VP.n5 24.5923
R1701 VP.n108 VP.n5 24.5923
R1702 VP.n109 VP.n108 24.5923
R1703 VP.n111 VP.n3 24.5923
R1704 VP.n115 VP.n3 24.5923
R1705 VP.n116 VP.n115 24.5923
R1706 VP.n121 VP.n1 24.5923
R1707 VP.n122 VP.n121 24.5923
R1708 VP.n66 VP.n17 24.5923
R1709 VP.n67 VP.n66 24.5923
R1710 VP.n49 VP.n21 24.5923
R1711 VP.n53 VP.n21 24.5923
R1712 VP.n54 VP.n53 24.5923
R1713 VP.n56 VP.n19 24.5923
R1714 VP.n60 VP.n19 24.5923
R1715 VP.n61 VP.n60 24.5923
R1716 VP.n36 VP.n25 24.5923
R1717 VP.n40 VP.n25 24.5923
R1718 VP.n41 VP.n40 24.5923
R1719 VP.n43 VP.n23 24.5923
R1720 VP.n47 VP.n23 24.5923
R1721 VP.n48 VP.n47 24.5923
R1722 VP.n30 VP.n27 24.5923
R1723 VP.n34 VP.n27 24.5923
R1724 VP.n35 VP.n34 24.5923
R1725 VP.n72 VP.n71 21.1495
R1726 VP.n123 VP.n122 21.1495
R1727 VP.n68 VP.n67 21.1495
R1728 VP.n85 VP.n84 16.7229
R1729 VP.n110 VP.n109 16.7229
R1730 VP.n55 VP.n54 16.7229
R1731 VP.n30 VP.n29 16.7229
R1732 VP.n97 VP.n96 12.2964
R1733 VP.n98 VP.n97 12.2964
R1734 VP.n42 VP.n41 12.2964
R1735 VP.n43 VP.n42 12.2964
R1736 VP.n84 VP.n83 7.86989
R1737 VP.n111 VP.n110 7.86989
R1738 VP.n56 VP.n55 7.86989
R1739 VP.n31 VP.n28 2.63942
R1740 VP.n69 VP.n16 0.417304
R1741 VP.n73 VP.n70 0.417304
R1742 VP.n124 VP.n0 0.417304
R1743 VP VP.n124 0.394524
R1744 VP.n32 VP.n31 0.189894
R1745 VP.n33 VP.n32 0.189894
R1746 VP.n33 VP.n26 0.189894
R1747 VP.n37 VP.n26 0.189894
R1748 VP.n38 VP.n37 0.189894
R1749 VP.n39 VP.n38 0.189894
R1750 VP.n39 VP.n24 0.189894
R1751 VP.n44 VP.n24 0.189894
R1752 VP.n45 VP.n44 0.189894
R1753 VP.n46 VP.n45 0.189894
R1754 VP.n46 VP.n22 0.189894
R1755 VP.n50 VP.n22 0.189894
R1756 VP.n51 VP.n50 0.189894
R1757 VP.n52 VP.n51 0.189894
R1758 VP.n52 VP.n20 0.189894
R1759 VP.n57 VP.n20 0.189894
R1760 VP.n58 VP.n57 0.189894
R1761 VP.n59 VP.n58 0.189894
R1762 VP.n59 VP.n18 0.189894
R1763 VP.n63 VP.n18 0.189894
R1764 VP.n64 VP.n63 0.189894
R1765 VP.n65 VP.n64 0.189894
R1766 VP.n65 VP.n16 0.189894
R1767 VP.n74 VP.n73 0.189894
R1768 VP.n75 VP.n74 0.189894
R1769 VP.n75 VP.n14 0.189894
R1770 VP.n79 VP.n14 0.189894
R1771 VP.n80 VP.n79 0.189894
R1772 VP.n81 VP.n80 0.189894
R1773 VP.n81 VP.n12 0.189894
R1774 VP.n86 VP.n12 0.189894
R1775 VP.n87 VP.n86 0.189894
R1776 VP.n88 VP.n87 0.189894
R1777 VP.n88 VP.n10 0.189894
R1778 VP.n92 VP.n10 0.189894
R1779 VP.n93 VP.n92 0.189894
R1780 VP.n94 VP.n93 0.189894
R1781 VP.n94 VP.n8 0.189894
R1782 VP.n99 VP.n8 0.189894
R1783 VP.n100 VP.n99 0.189894
R1784 VP.n101 VP.n100 0.189894
R1785 VP.n101 VP.n6 0.189894
R1786 VP.n105 VP.n6 0.189894
R1787 VP.n106 VP.n105 0.189894
R1788 VP.n107 VP.n106 0.189894
R1789 VP.n107 VP.n4 0.189894
R1790 VP.n112 VP.n4 0.189894
R1791 VP.n113 VP.n112 0.189894
R1792 VP.n114 VP.n113 0.189894
R1793 VP.n114 VP.n2 0.189894
R1794 VP.n118 VP.n2 0.189894
R1795 VP.n119 VP.n118 0.189894
R1796 VP.n120 VP.n119 0.189894
R1797 VP.n120 VP.n0 0.189894
R1798 VDD1.n1 VDD1.t6 95.6331
R1799 VDD1.n3 VDD1.t7 95.6328
R1800 VDD1.n5 VDD1.n4 90.1309
R1801 VDD1.n1 VDD1.n0 87.5419
R1802 VDD1.n3 VDD1.n2 87.5418
R1803 VDD1.n7 VDD1.n6 87.5417
R1804 VDD1.n7 VDD1.n5 48.947
R1805 VDD1.n6 VDD1.t9 4.56581
R1806 VDD1.n6 VDD1.t2 4.56581
R1807 VDD1.n0 VDD1.t8 4.56581
R1808 VDD1.n0 VDD1.t1 4.56581
R1809 VDD1.n4 VDD1.t0 4.56581
R1810 VDD1.n4 VDD1.t4 4.56581
R1811 VDD1.n2 VDD1.t3 4.56581
R1812 VDD1.n2 VDD1.t5 4.56581
R1813 VDD1 VDD1.n7 2.58671
R1814 VDD1 VDD1.n1 0.940155
R1815 VDD1.n5 VDD1.n3 0.826619
C0 w_n5878_n2392# VDD2 3.09974f
C1 VDD1 B 2.53665f
C2 VN VDD2 6.95802f
C3 VN w_n5878_n2392# 12.8277f
C4 VTAIL B 3.0022f
C5 VP VDD1 7.52994f
C6 VP VTAIL 8.61365f
C7 VDD1 VDD2 2.93036f
C8 VP B 2.82474f
C9 w_n5878_n2392# VDD1 2.8959f
C10 VN VDD1 0.156427f
C11 VTAIL VDD2 9.1442f
C12 VTAIL w_n5878_n2392# 2.72357f
C13 VN VTAIL 8.59923f
C14 B VDD2 2.69974f
C15 w_n5878_n2392# B 11.132f
C16 VN B 1.52545f
C17 VP VDD2 0.731483f
C18 VP w_n5878_n2392# 13.5966f
C19 VP VN 9.20185f
C20 VTAIL VDD1 9.08377f
C21 VDD2 VSUBS 2.569056f
C22 VDD1 VSUBS 2.339155f
C23 VTAIL VSUBS 0.82964f
C24 VN VSUBS 9.38395f
C25 VP VSUBS 5.262846f
C26 B VSUBS 6.393545f
C27 w_n5878_n2392# VSUBS 0.174859p
C28 VDD1.t6 VSUBS 1.82279f
C29 VDD1.t8 VSUBS 0.193011f
C30 VDD1.t1 VSUBS 0.193011f
C31 VDD1.n0 VSUBS 1.33986f
C32 VDD1.n1 VSUBS 2.10853f
C33 VDD1.t7 VSUBS 1.82278f
C34 VDD1.t3 VSUBS 0.193011f
C35 VDD1.t5 VSUBS 0.193011f
C36 VDD1.n2 VSUBS 1.33986f
C37 VDD1.n3 VSUBS 2.09695f
C38 VDD1.t0 VSUBS 0.193011f
C39 VDD1.t4 VSUBS 0.193011f
C40 VDD1.n4 VSUBS 1.37646f
C41 VDD1.n5 VSUBS 4.91386f
C42 VDD1.t9 VSUBS 0.193011f
C43 VDD1.t2 VSUBS 0.193011f
C44 VDD1.n6 VSUBS 1.33986f
C45 VDD1.n7 VSUBS 4.80524f
C46 VP.n0 VSUBS 0.059736f
C47 VP.t5 VSUBS 2.27174f
C48 VP.n1 VSUBS 0.062737f
C49 VP.n2 VSUBS 0.031767f
C50 VP.n3 VSUBS 0.058909f
C51 VP.n4 VSUBS 0.031767f
C52 VP.t9 VSUBS 2.27174f
C53 VP.n5 VSUBS 0.058909f
C54 VP.n6 VSUBS 0.031767f
C55 VP.n7 VSUBS 0.058909f
C56 VP.n8 VSUBS 0.031767f
C57 VP.t4 VSUBS 2.27174f
C58 VP.n9 VSUBS 0.058909f
C59 VP.n10 VSUBS 0.031767f
C60 VP.n11 VSUBS 0.058909f
C61 VP.n12 VSUBS 0.031767f
C62 VP.t6 VSUBS 2.27174f
C63 VP.n13 VSUBS 0.058909f
C64 VP.n14 VSUBS 0.031767f
C65 VP.n15 VSUBS 0.058909f
C66 VP.n16 VSUBS 0.059736f
C67 VP.t7 VSUBS 2.27174f
C68 VP.n17 VSUBS 0.062737f
C69 VP.n18 VSUBS 0.031767f
C70 VP.n19 VSUBS 0.058909f
C71 VP.n20 VSUBS 0.031767f
C72 VP.t0 VSUBS 2.27174f
C73 VP.n21 VSUBS 0.058909f
C74 VP.n22 VSUBS 0.031767f
C75 VP.n23 VSUBS 0.058909f
C76 VP.n24 VSUBS 0.031767f
C77 VP.t8 VSUBS 2.27174f
C78 VP.n25 VSUBS 0.058909f
C79 VP.n26 VSUBS 0.031767f
C80 VP.n27 VSUBS 0.058909f
C81 VP.t3 VSUBS 2.7145f
C82 VP.n28 VSUBS 0.90412f
C83 VP.t1 VSUBS 2.27174f
C84 VP.n29 VSUBS 0.9417f
C85 VP.n30 VSUBS 0.049603f
C86 VP.n31 VSUBS 0.413344f
C87 VP.n32 VSUBS 0.031767f
C88 VP.n33 VSUBS 0.031767f
C89 VP.n34 VSUBS 0.058909f
C90 VP.n35 VSUBS 0.042223f
C91 VP.n36 VSUBS 0.050133f
C92 VP.n37 VSUBS 0.031767f
C93 VP.n38 VSUBS 0.031767f
C94 VP.n39 VSUBS 0.031767f
C95 VP.n40 VSUBS 0.058909f
C96 VP.n41 VSUBS 0.044368f
C97 VP.n42 VSUBS 0.823522f
C98 VP.n43 VSUBS 0.044368f
C99 VP.n44 VSUBS 0.031767f
C100 VP.n45 VSUBS 0.031767f
C101 VP.n46 VSUBS 0.031767f
C102 VP.n47 VSUBS 0.058909f
C103 VP.n48 VSUBS 0.050133f
C104 VP.n49 VSUBS 0.042223f
C105 VP.n50 VSUBS 0.031767f
C106 VP.n51 VSUBS 0.031767f
C107 VP.n52 VSUBS 0.031767f
C108 VP.n53 VSUBS 0.058909f
C109 VP.n54 VSUBS 0.049603f
C110 VP.n55 VSUBS 0.823522f
C111 VP.n56 VSUBS 0.039133f
C112 VP.n57 VSUBS 0.031767f
C113 VP.n58 VSUBS 0.031767f
C114 VP.n59 VSUBS 0.031767f
C115 VP.n60 VSUBS 0.058909f
C116 VP.n61 VSUBS 0.057078f
C117 VP.n62 VSUBS 0.031449f
C118 VP.n63 VSUBS 0.031767f
C119 VP.n64 VSUBS 0.031767f
C120 VP.n65 VSUBS 0.031767f
C121 VP.n66 VSUBS 0.058909f
C122 VP.n67 VSUBS 0.054837f
C123 VP.n68 VSUBS 0.957988f
C124 VP.n69 VSUBS 2.1496f
C125 VP.n70 VSUBS 2.17008f
C126 VP.t2 VSUBS 2.27174f
C127 VP.n71 VSUBS 0.957988f
C128 VP.n72 VSUBS 0.054837f
C129 VP.n73 VSUBS 0.059736f
C130 VP.n74 VSUBS 0.031767f
C131 VP.n75 VSUBS 0.031767f
C132 VP.n76 VSUBS 0.062737f
C133 VP.n77 VSUBS 0.031449f
C134 VP.n78 VSUBS 0.057078f
C135 VP.n79 VSUBS 0.031767f
C136 VP.n80 VSUBS 0.031767f
C137 VP.n81 VSUBS 0.031767f
C138 VP.n82 VSUBS 0.058909f
C139 VP.n83 VSUBS 0.039133f
C140 VP.n84 VSUBS 0.823522f
C141 VP.n85 VSUBS 0.049603f
C142 VP.n86 VSUBS 0.031767f
C143 VP.n87 VSUBS 0.031767f
C144 VP.n88 VSUBS 0.031767f
C145 VP.n89 VSUBS 0.058909f
C146 VP.n90 VSUBS 0.042223f
C147 VP.n91 VSUBS 0.050133f
C148 VP.n92 VSUBS 0.031767f
C149 VP.n93 VSUBS 0.031767f
C150 VP.n94 VSUBS 0.031767f
C151 VP.n95 VSUBS 0.058909f
C152 VP.n96 VSUBS 0.044368f
C153 VP.n97 VSUBS 0.823522f
C154 VP.n98 VSUBS 0.044368f
C155 VP.n99 VSUBS 0.031767f
C156 VP.n100 VSUBS 0.031767f
C157 VP.n101 VSUBS 0.031767f
C158 VP.n102 VSUBS 0.058909f
C159 VP.n103 VSUBS 0.050133f
C160 VP.n104 VSUBS 0.042223f
C161 VP.n105 VSUBS 0.031767f
C162 VP.n106 VSUBS 0.031767f
C163 VP.n107 VSUBS 0.031767f
C164 VP.n108 VSUBS 0.058909f
C165 VP.n109 VSUBS 0.049603f
C166 VP.n110 VSUBS 0.823522f
C167 VP.n111 VSUBS 0.039133f
C168 VP.n112 VSUBS 0.031767f
C169 VP.n113 VSUBS 0.031767f
C170 VP.n114 VSUBS 0.031767f
C171 VP.n115 VSUBS 0.058909f
C172 VP.n116 VSUBS 0.057078f
C173 VP.n117 VSUBS 0.031449f
C174 VP.n118 VSUBS 0.031767f
C175 VP.n119 VSUBS 0.031767f
C176 VP.n120 VSUBS 0.031767f
C177 VP.n121 VSUBS 0.058909f
C178 VP.n122 VSUBS 0.054837f
C179 VP.n123 VSUBS 0.957988f
C180 VP.n124 VSUBS 0.09669f
C181 VDD2.t4 VSUBS 1.82475f
C182 VDD2.t8 VSUBS 0.193219f
C183 VDD2.t1 VSUBS 0.193219f
C184 VDD2.n0 VSUBS 1.3413f
C185 VDD2.n1 VSUBS 2.09921f
C186 VDD2.t0 VSUBS 0.193219f
C187 VDD2.t7 VSUBS 0.193219f
C188 VDD2.n2 VSUBS 1.37794f
C189 VDD2.n3 VSUBS 4.70944f
C190 VDD2.t5 VSUBS 1.78524f
C191 VDD2.n4 VSUBS 4.69013f
C192 VDD2.t2 VSUBS 0.193219f
C193 VDD2.t9 VSUBS 0.193219f
C194 VDD2.n5 VSUBS 1.34131f
C195 VDD2.n6 VSUBS 1.07872f
C196 VDD2.t6 VSUBS 0.193219f
C197 VDD2.t3 VSUBS 0.193219f
C198 VDD2.n7 VSUBS 1.37788f
C199 VTAIL.t12 VSUBS 0.18951f
C200 VTAIL.t17 VSUBS 0.18951f
C201 VTAIL.n0 VSUBS 1.18212f
C202 VTAIL.n1 VSUBS 1.19667f
C203 VTAIL.t6 VSUBS 1.6076f
C204 VTAIL.n2 VSUBS 1.37738f
C205 VTAIL.t3 VSUBS 0.18951f
C206 VTAIL.t8 VSUBS 0.18951f
C207 VTAIL.n3 VSUBS 1.18212f
C208 VTAIL.n4 VSUBS 1.42636f
C209 VTAIL.t0 VSUBS 0.18951f
C210 VTAIL.t5 VSUBS 0.18951f
C211 VTAIL.n5 VSUBS 1.18212f
C212 VTAIL.n6 VSUBS 2.93272f
C213 VTAIL.t9 VSUBS 0.18951f
C214 VTAIL.t13 VSUBS 0.18951f
C215 VTAIL.n7 VSUBS 1.18212f
C216 VTAIL.n8 VSUBS 2.93271f
C217 VTAIL.t18 VSUBS 0.18951f
C218 VTAIL.t11 VSUBS 0.18951f
C219 VTAIL.n9 VSUBS 1.18212f
C220 VTAIL.n10 VSUBS 1.42636f
C221 VTAIL.t16 VSUBS 1.60761f
C222 VTAIL.n11 VSUBS 1.37737f
C223 VTAIL.t1 VSUBS 0.18951f
C224 VTAIL.t2 VSUBS 0.18951f
C225 VTAIL.n12 VSUBS 1.18212f
C226 VTAIL.n13 VSUBS 1.28601f
C227 VTAIL.t7 VSUBS 0.18951f
C228 VTAIL.t19 VSUBS 0.18951f
C229 VTAIL.n14 VSUBS 1.18212f
C230 VTAIL.n15 VSUBS 1.42636f
C231 VTAIL.t4 VSUBS 1.6076f
C232 VTAIL.n16 VSUBS 2.64141f
C233 VTAIL.t10 VSUBS 1.6076f
C234 VTAIL.n17 VSUBS 2.64141f
C235 VTAIL.t14 VSUBS 0.18951f
C236 VTAIL.t15 VSUBS 0.18951f
C237 VTAIL.n18 VSUBS 1.18212f
C238 VTAIL.n19 VSUBS 1.13305f
C239 VN.n0 VSUBS 0.053805f
C240 VN.t2 VSUBS 2.04619f
C241 VN.n1 VSUBS 0.056508f
C242 VN.n2 VSUBS 0.028613f
C243 VN.n3 VSUBS 0.05306f
C244 VN.n4 VSUBS 0.028613f
C245 VN.t9 VSUBS 2.04619f
C246 VN.n5 VSUBS 0.05306f
C247 VN.n6 VSUBS 0.028613f
C248 VN.n7 VSUBS 0.05306f
C249 VN.n8 VSUBS 0.028613f
C250 VN.t8 VSUBS 2.04619f
C251 VN.n9 VSUBS 0.05306f
C252 VN.n10 VSUBS 0.028613f
C253 VN.n11 VSUBS 0.05306f
C254 VN.t5 VSUBS 2.445f
C255 VN.n12 VSUBS 0.814351f
C256 VN.t1 VSUBS 2.04619f
C257 VN.n13 VSUBS 0.848203f
C258 VN.n14 VSUBS 0.044678f
C259 VN.n15 VSUBS 0.372304f
C260 VN.n16 VSUBS 0.028613f
C261 VN.n17 VSUBS 0.028613f
C262 VN.n18 VSUBS 0.05306f
C263 VN.n19 VSUBS 0.038031f
C264 VN.n20 VSUBS 0.045155f
C265 VN.n21 VSUBS 0.028613f
C266 VN.n22 VSUBS 0.028613f
C267 VN.n23 VSUBS 0.028613f
C268 VN.n24 VSUBS 0.05306f
C269 VN.n25 VSUBS 0.039963f
C270 VN.n26 VSUBS 0.741758f
C271 VN.n27 VSUBS 0.039963f
C272 VN.n28 VSUBS 0.028613f
C273 VN.n29 VSUBS 0.028613f
C274 VN.n30 VSUBS 0.028613f
C275 VN.n31 VSUBS 0.05306f
C276 VN.n32 VSUBS 0.045155f
C277 VN.n33 VSUBS 0.038031f
C278 VN.n34 VSUBS 0.028613f
C279 VN.n35 VSUBS 0.028613f
C280 VN.n36 VSUBS 0.028613f
C281 VN.n37 VSUBS 0.05306f
C282 VN.n38 VSUBS 0.044678f
C283 VN.n39 VSUBS 0.741758f
C284 VN.n40 VSUBS 0.035248f
C285 VN.n41 VSUBS 0.028613f
C286 VN.n42 VSUBS 0.028613f
C287 VN.n43 VSUBS 0.028613f
C288 VN.n44 VSUBS 0.05306f
C289 VN.n45 VSUBS 0.051411f
C290 VN.n46 VSUBS 0.028327f
C291 VN.n47 VSUBS 0.028613f
C292 VN.n48 VSUBS 0.028613f
C293 VN.n49 VSUBS 0.028613f
C294 VN.n50 VSUBS 0.05306f
C295 VN.n51 VSUBS 0.049393f
C296 VN.n52 VSUBS 0.862874f
C297 VN.n53 VSUBS 0.08709f
C298 VN.n54 VSUBS 0.053805f
C299 VN.t4 VSUBS 2.04619f
C300 VN.n55 VSUBS 0.056508f
C301 VN.n56 VSUBS 0.028613f
C302 VN.n57 VSUBS 0.05306f
C303 VN.n58 VSUBS 0.028613f
C304 VN.t7 VSUBS 2.04619f
C305 VN.n59 VSUBS 0.05306f
C306 VN.n60 VSUBS 0.028613f
C307 VN.n61 VSUBS 0.05306f
C308 VN.n62 VSUBS 0.028613f
C309 VN.t0 VSUBS 2.04619f
C310 VN.n63 VSUBS 0.05306f
C311 VN.n64 VSUBS 0.028613f
C312 VN.n65 VSUBS 0.05306f
C313 VN.t6 VSUBS 2.445f
C314 VN.n66 VSUBS 0.814351f
C315 VN.t3 VSUBS 2.04619f
C316 VN.n67 VSUBS 0.848203f
C317 VN.n68 VSUBS 0.044678f
C318 VN.n69 VSUBS 0.372304f
C319 VN.n70 VSUBS 0.028613f
C320 VN.n71 VSUBS 0.028613f
C321 VN.n72 VSUBS 0.05306f
C322 VN.n73 VSUBS 0.038031f
C323 VN.n74 VSUBS 0.045155f
C324 VN.n75 VSUBS 0.028613f
C325 VN.n76 VSUBS 0.028613f
C326 VN.n77 VSUBS 0.028613f
C327 VN.n78 VSUBS 0.05306f
C328 VN.n79 VSUBS 0.039963f
C329 VN.n80 VSUBS 0.741758f
C330 VN.n81 VSUBS 0.039963f
C331 VN.n82 VSUBS 0.028613f
C332 VN.n83 VSUBS 0.028613f
C333 VN.n84 VSUBS 0.028613f
C334 VN.n85 VSUBS 0.05306f
C335 VN.n86 VSUBS 0.045155f
C336 VN.n87 VSUBS 0.038031f
C337 VN.n88 VSUBS 0.028613f
C338 VN.n89 VSUBS 0.028613f
C339 VN.n90 VSUBS 0.028613f
C340 VN.n91 VSUBS 0.05306f
C341 VN.n92 VSUBS 0.044678f
C342 VN.n93 VSUBS 0.741758f
C343 VN.n94 VSUBS 0.035248f
C344 VN.n95 VSUBS 0.028613f
C345 VN.n96 VSUBS 0.028613f
C346 VN.n97 VSUBS 0.028613f
C347 VN.n98 VSUBS 0.05306f
C348 VN.n99 VSUBS 0.051411f
C349 VN.n100 VSUBS 0.028327f
C350 VN.n101 VSUBS 0.028613f
C351 VN.n102 VSUBS 0.028613f
C352 VN.n103 VSUBS 0.028613f
C353 VN.n104 VSUBS 0.05306f
C354 VN.n105 VSUBS 0.049393f
C355 VN.n106 VSUBS 0.862874f
C356 VN.n107 VSUBS 1.94307f
C357 B.n0 VSUBS 0.009508f
C358 B.n1 VSUBS 0.009508f
C359 B.n2 VSUBS 0.014062f
C360 B.n3 VSUBS 0.010776f
C361 B.n4 VSUBS 0.010776f
C362 B.n5 VSUBS 0.010776f
C363 B.n6 VSUBS 0.010776f
C364 B.n7 VSUBS 0.010776f
C365 B.n8 VSUBS 0.010776f
C366 B.n9 VSUBS 0.010776f
C367 B.n10 VSUBS 0.010776f
C368 B.n11 VSUBS 0.010776f
C369 B.n12 VSUBS 0.010776f
C370 B.n13 VSUBS 0.010776f
C371 B.n14 VSUBS 0.010776f
C372 B.n15 VSUBS 0.010776f
C373 B.n16 VSUBS 0.010776f
C374 B.n17 VSUBS 0.010776f
C375 B.n18 VSUBS 0.010776f
C376 B.n19 VSUBS 0.010776f
C377 B.n20 VSUBS 0.010776f
C378 B.n21 VSUBS 0.010776f
C379 B.n22 VSUBS 0.010776f
C380 B.n23 VSUBS 0.010776f
C381 B.n24 VSUBS 0.010776f
C382 B.n25 VSUBS 0.010776f
C383 B.n26 VSUBS 0.010776f
C384 B.n27 VSUBS 0.010776f
C385 B.n28 VSUBS 0.010776f
C386 B.n29 VSUBS 0.010776f
C387 B.n30 VSUBS 0.010776f
C388 B.n31 VSUBS 0.010776f
C389 B.n32 VSUBS 0.010776f
C390 B.n33 VSUBS 0.010776f
C391 B.n34 VSUBS 0.010776f
C392 B.n35 VSUBS 0.010776f
C393 B.n36 VSUBS 0.010776f
C394 B.n37 VSUBS 0.010776f
C395 B.n38 VSUBS 0.010776f
C396 B.n39 VSUBS 0.010776f
C397 B.n40 VSUBS 0.010776f
C398 B.n41 VSUBS 0.010776f
C399 B.n42 VSUBS 0.024592f
C400 B.n43 VSUBS 0.010776f
C401 B.n44 VSUBS 0.010776f
C402 B.n45 VSUBS 0.010776f
C403 B.n46 VSUBS 0.010776f
C404 B.n47 VSUBS 0.010776f
C405 B.n48 VSUBS 0.010776f
C406 B.n49 VSUBS 0.010776f
C407 B.n50 VSUBS 0.010776f
C408 B.n51 VSUBS 0.010776f
C409 B.n52 VSUBS 0.010776f
C410 B.n53 VSUBS 0.010776f
C411 B.n54 VSUBS 0.010776f
C412 B.n55 VSUBS 0.010776f
C413 B.t7 VSUBS 0.331088f
C414 B.t8 VSUBS 0.372512f
C415 B.t6 VSUBS 1.96771f
C416 B.n56 VSUBS 0.222794f
C417 B.n57 VSUBS 0.117236f
C418 B.n58 VSUBS 0.010776f
C419 B.n59 VSUBS 0.010776f
C420 B.n60 VSUBS 0.010776f
C421 B.n61 VSUBS 0.010776f
C422 B.n62 VSUBS 0.006022f
C423 B.n63 VSUBS 0.010776f
C424 B.t4 VSUBS 0.331086f
C425 B.t5 VSUBS 0.372509f
C426 B.t3 VSUBS 1.96771f
C427 B.n64 VSUBS 0.222796f
C428 B.n65 VSUBS 0.117238f
C429 B.n66 VSUBS 0.024967f
C430 B.n67 VSUBS 0.010776f
C431 B.n68 VSUBS 0.010776f
C432 B.n69 VSUBS 0.010776f
C433 B.n70 VSUBS 0.010776f
C434 B.n71 VSUBS 0.010776f
C435 B.n72 VSUBS 0.010776f
C436 B.n73 VSUBS 0.010776f
C437 B.n74 VSUBS 0.010776f
C438 B.n75 VSUBS 0.010776f
C439 B.n76 VSUBS 0.010776f
C440 B.n77 VSUBS 0.010776f
C441 B.n78 VSUBS 0.010776f
C442 B.n79 VSUBS 0.0239f
C443 B.n80 VSUBS 0.010776f
C444 B.n81 VSUBS 0.010776f
C445 B.n82 VSUBS 0.010776f
C446 B.n83 VSUBS 0.010776f
C447 B.n84 VSUBS 0.010776f
C448 B.n85 VSUBS 0.010776f
C449 B.n86 VSUBS 0.010776f
C450 B.n87 VSUBS 0.010776f
C451 B.n88 VSUBS 0.010776f
C452 B.n89 VSUBS 0.010776f
C453 B.n90 VSUBS 0.010776f
C454 B.n91 VSUBS 0.010776f
C455 B.n92 VSUBS 0.010776f
C456 B.n93 VSUBS 0.010776f
C457 B.n94 VSUBS 0.010776f
C458 B.n95 VSUBS 0.010776f
C459 B.n96 VSUBS 0.010776f
C460 B.n97 VSUBS 0.010776f
C461 B.n98 VSUBS 0.010776f
C462 B.n99 VSUBS 0.010776f
C463 B.n100 VSUBS 0.010776f
C464 B.n101 VSUBS 0.010776f
C465 B.n102 VSUBS 0.010776f
C466 B.n103 VSUBS 0.010776f
C467 B.n104 VSUBS 0.010776f
C468 B.n105 VSUBS 0.010776f
C469 B.n106 VSUBS 0.010776f
C470 B.n107 VSUBS 0.010776f
C471 B.n108 VSUBS 0.010776f
C472 B.n109 VSUBS 0.010776f
C473 B.n110 VSUBS 0.010776f
C474 B.n111 VSUBS 0.010776f
C475 B.n112 VSUBS 0.010776f
C476 B.n113 VSUBS 0.010776f
C477 B.n114 VSUBS 0.010776f
C478 B.n115 VSUBS 0.010776f
C479 B.n116 VSUBS 0.010776f
C480 B.n117 VSUBS 0.010776f
C481 B.n118 VSUBS 0.010776f
C482 B.n119 VSUBS 0.010776f
C483 B.n120 VSUBS 0.010776f
C484 B.n121 VSUBS 0.010776f
C485 B.n122 VSUBS 0.010776f
C486 B.n123 VSUBS 0.010776f
C487 B.n124 VSUBS 0.010776f
C488 B.n125 VSUBS 0.010776f
C489 B.n126 VSUBS 0.010776f
C490 B.n127 VSUBS 0.010776f
C491 B.n128 VSUBS 0.010776f
C492 B.n129 VSUBS 0.010776f
C493 B.n130 VSUBS 0.010776f
C494 B.n131 VSUBS 0.010776f
C495 B.n132 VSUBS 0.010776f
C496 B.n133 VSUBS 0.010776f
C497 B.n134 VSUBS 0.010776f
C498 B.n135 VSUBS 0.010776f
C499 B.n136 VSUBS 0.010776f
C500 B.n137 VSUBS 0.010776f
C501 B.n138 VSUBS 0.010776f
C502 B.n139 VSUBS 0.010776f
C503 B.n140 VSUBS 0.010776f
C504 B.n141 VSUBS 0.010776f
C505 B.n142 VSUBS 0.010776f
C506 B.n143 VSUBS 0.010776f
C507 B.n144 VSUBS 0.010776f
C508 B.n145 VSUBS 0.010776f
C509 B.n146 VSUBS 0.010776f
C510 B.n147 VSUBS 0.010776f
C511 B.n148 VSUBS 0.010776f
C512 B.n149 VSUBS 0.010776f
C513 B.n150 VSUBS 0.010776f
C514 B.n151 VSUBS 0.010776f
C515 B.n152 VSUBS 0.010776f
C516 B.n153 VSUBS 0.010776f
C517 B.n154 VSUBS 0.010776f
C518 B.n155 VSUBS 0.010776f
C519 B.n156 VSUBS 0.010776f
C520 B.n157 VSUBS 0.010776f
C521 B.n158 VSUBS 0.010776f
C522 B.n159 VSUBS 0.010776f
C523 B.n160 VSUBS 0.024592f
C524 B.n161 VSUBS 0.010776f
C525 B.n162 VSUBS 0.010776f
C526 B.n163 VSUBS 0.010776f
C527 B.n164 VSUBS 0.010776f
C528 B.n165 VSUBS 0.010776f
C529 B.n166 VSUBS 0.010776f
C530 B.n167 VSUBS 0.010776f
C531 B.n168 VSUBS 0.010776f
C532 B.n169 VSUBS 0.010776f
C533 B.n170 VSUBS 0.010776f
C534 B.n171 VSUBS 0.010776f
C535 B.n172 VSUBS 0.010776f
C536 B.n173 VSUBS 0.010142f
C537 B.n174 VSUBS 0.010776f
C538 B.n175 VSUBS 0.010776f
C539 B.n176 VSUBS 0.010776f
C540 B.n177 VSUBS 0.010776f
C541 B.n178 VSUBS 0.010776f
C542 B.t11 VSUBS 0.331088f
C543 B.t10 VSUBS 0.372512f
C544 B.t9 VSUBS 1.96771f
C545 B.n179 VSUBS 0.222794f
C546 B.n180 VSUBS 0.117236f
C547 B.n181 VSUBS 0.010776f
C548 B.n182 VSUBS 0.010776f
C549 B.n183 VSUBS 0.010776f
C550 B.n184 VSUBS 0.010776f
C551 B.n185 VSUBS 0.010776f
C552 B.n186 VSUBS 0.010776f
C553 B.n187 VSUBS 0.010776f
C554 B.n188 VSUBS 0.010776f
C555 B.n189 VSUBS 0.010776f
C556 B.n190 VSUBS 0.010776f
C557 B.n191 VSUBS 0.010776f
C558 B.n192 VSUBS 0.010776f
C559 B.n193 VSUBS 0.010776f
C560 B.n194 VSUBS 0.0239f
C561 B.n195 VSUBS 0.010776f
C562 B.n196 VSUBS 0.010776f
C563 B.n197 VSUBS 0.010776f
C564 B.n198 VSUBS 0.010776f
C565 B.n199 VSUBS 0.010776f
C566 B.n200 VSUBS 0.010776f
C567 B.n201 VSUBS 0.010776f
C568 B.n202 VSUBS 0.010776f
C569 B.n203 VSUBS 0.010776f
C570 B.n204 VSUBS 0.010776f
C571 B.n205 VSUBS 0.010776f
C572 B.n206 VSUBS 0.010776f
C573 B.n207 VSUBS 0.010776f
C574 B.n208 VSUBS 0.010776f
C575 B.n209 VSUBS 0.010776f
C576 B.n210 VSUBS 0.010776f
C577 B.n211 VSUBS 0.010776f
C578 B.n212 VSUBS 0.010776f
C579 B.n213 VSUBS 0.010776f
C580 B.n214 VSUBS 0.010776f
C581 B.n215 VSUBS 0.010776f
C582 B.n216 VSUBS 0.010776f
C583 B.n217 VSUBS 0.010776f
C584 B.n218 VSUBS 0.010776f
C585 B.n219 VSUBS 0.010776f
C586 B.n220 VSUBS 0.010776f
C587 B.n221 VSUBS 0.010776f
C588 B.n222 VSUBS 0.010776f
C589 B.n223 VSUBS 0.010776f
C590 B.n224 VSUBS 0.010776f
C591 B.n225 VSUBS 0.010776f
C592 B.n226 VSUBS 0.010776f
C593 B.n227 VSUBS 0.010776f
C594 B.n228 VSUBS 0.010776f
C595 B.n229 VSUBS 0.010776f
C596 B.n230 VSUBS 0.010776f
C597 B.n231 VSUBS 0.010776f
C598 B.n232 VSUBS 0.010776f
C599 B.n233 VSUBS 0.010776f
C600 B.n234 VSUBS 0.010776f
C601 B.n235 VSUBS 0.010776f
C602 B.n236 VSUBS 0.010776f
C603 B.n237 VSUBS 0.010776f
C604 B.n238 VSUBS 0.010776f
C605 B.n239 VSUBS 0.010776f
C606 B.n240 VSUBS 0.010776f
C607 B.n241 VSUBS 0.010776f
C608 B.n242 VSUBS 0.010776f
C609 B.n243 VSUBS 0.010776f
C610 B.n244 VSUBS 0.010776f
C611 B.n245 VSUBS 0.010776f
C612 B.n246 VSUBS 0.010776f
C613 B.n247 VSUBS 0.010776f
C614 B.n248 VSUBS 0.010776f
C615 B.n249 VSUBS 0.010776f
C616 B.n250 VSUBS 0.010776f
C617 B.n251 VSUBS 0.010776f
C618 B.n252 VSUBS 0.010776f
C619 B.n253 VSUBS 0.010776f
C620 B.n254 VSUBS 0.010776f
C621 B.n255 VSUBS 0.010776f
C622 B.n256 VSUBS 0.010776f
C623 B.n257 VSUBS 0.010776f
C624 B.n258 VSUBS 0.010776f
C625 B.n259 VSUBS 0.010776f
C626 B.n260 VSUBS 0.010776f
C627 B.n261 VSUBS 0.010776f
C628 B.n262 VSUBS 0.010776f
C629 B.n263 VSUBS 0.010776f
C630 B.n264 VSUBS 0.010776f
C631 B.n265 VSUBS 0.010776f
C632 B.n266 VSUBS 0.010776f
C633 B.n267 VSUBS 0.010776f
C634 B.n268 VSUBS 0.010776f
C635 B.n269 VSUBS 0.010776f
C636 B.n270 VSUBS 0.010776f
C637 B.n271 VSUBS 0.010776f
C638 B.n272 VSUBS 0.010776f
C639 B.n273 VSUBS 0.010776f
C640 B.n274 VSUBS 0.010776f
C641 B.n275 VSUBS 0.010776f
C642 B.n276 VSUBS 0.010776f
C643 B.n277 VSUBS 0.010776f
C644 B.n278 VSUBS 0.010776f
C645 B.n279 VSUBS 0.010776f
C646 B.n280 VSUBS 0.010776f
C647 B.n281 VSUBS 0.010776f
C648 B.n282 VSUBS 0.010776f
C649 B.n283 VSUBS 0.010776f
C650 B.n284 VSUBS 0.010776f
C651 B.n285 VSUBS 0.010776f
C652 B.n286 VSUBS 0.010776f
C653 B.n287 VSUBS 0.010776f
C654 B.n288 VSUBS 0.010776f
C655 B.n289 VSUBS 0.010776f
C656 B.n290 VSUBS 0.010776f
C657 B.n291 VSUBS 0.010776f
C658 B.n292 VSUBS 0.010776f
C659 B.n293 VSUBS 0.010776f
C660 B.n294 VSUBS 0.010776f
C661 B.n295 VSUBS 0.010776f
C662 B.n296 VSUBS 0.010776f
C663 B.n297 VSUBS 0.010776f
C664 B.n298 VSUBS 0.010776f
C665 B.n299 VSUBS 0.010776f
C666 B.n300 VSUBS 0.010776f
C667 B.n301 VSUBS 0.010776f
C668 B.n302 VSUBS 0.010776f
C669 B.n303 VSUBS 0.010776f
C670 B.n304 VSUBS 0.010776f
C671 B.n305 VSUBS 0.010776f
C672 B.n306 VSUBS 0.010776f
C673 B.n307 VSUBS 0.010776f
C674 B.n308 VSUBS 0.010776f
C675 B.n309 VSUBS 0.010776f
C676 B.n310 VSUBS 0.010776f
C677 B.n311 VSUBS 0.010776f
C678 B.n312 VSUBS 0.010776f
C679 B.n313 VSUBS 0.010776f
C680 B.n314 VSUBS 0.010776f
C681 B.n315 VSUBS 0.010776f
C682 B.n316 VSUBS 0.010776f
C683 B.n317 VSUBS 0.010776f
C684 B.n318 VSUBS 0.010776f
C685 B.n319 VSUBS 0.010776f
C686 B.n320 VSUBS 0.010776f
C687 B.n321 VSUBS 0.010776f
C688 B.n322 VSUBS 0.010776f
C689 B.n323 VSUBS 0.010776f
C690 B.n324 VSUBS 0.010776f
C691 B.n325 VSUBS 0.010776f
C692 B.n326 VSUBS 0.010776f
C693 B.n327 VSUBS 0.010776f
C694 B.n328 VSUBS 0.010776f
C695 B.n329 VSUBS 0.010776f
C696 B.n330 VSUBS 0.010776f
C697 B.n331 VSUBS 0.010776f
C698 B.n332 VSUBS 0.010776f
C699 B.n333 VSUBS 0.010776f
C700 B.n334 VSUBS 0.010776f
C701 B.n335 VSUBS 0.010776f
C702 B.n336 VSUBS 0.010776f
C703 B.n337 VSUBS 0.010776f
C704 B.n338 VSUBS 0.010776f
C705 B.n339 VSUBS 0.010776f
C706 B.n340 VSUBS 0.010776f
C707 B.n341 VSUBS 0.010776f
C708 B.n342 VSUBS 0.010776f
C709 B.n343 VSUBS 0.010776f
C710 B.n344 VSUBS 0.010776f
C711 B.n345 VSUBS 0.010776f
C712 B.n346 VSUBS 0.010776f
C713 B.n347 VSUBS 0.010776f
C714 B.n348 VSUBS 0.010776f
C715 B.n349 VSUBS 0.010776f
C716 B.n350 VSUBS 0.010776f
C717 B.n351 VSUBS 0.0239f
C718 B.n352 VSUBS 0.024592f
C719 B.n353 VSUBS 0.024592f
C720 B.n354 VSUBS 0.010776f
C721 B.n355 VSUBS 0.010776f
C722 B.n356 VSUBS 0.010776f
C723 B.n357 VSUBS 0.010776f
C724 B.n358 VSUBS 0.010776f
C725 B.n359 VSUBS 0.010776f
C726 B.n360 VSUBS 0.010776f
C727 B.n361 VSUBS 0.010776f
C728 B.n362 VSUBS 0.010776f
C729 B.n363 VSUBS 0.010776f
C730 B.n364 VSUBS 0.010776f
C731 B.n365 VSUBS 0.010776f
C732 B.n366 VSUBS 0.010776f
C733 B.n367 VSUBS 0.010776f
C734 B.n368 VSUBS 0.010776f
C735 B.n369 VSUBS 0.010776f
C736 B.n370 VSUBS 0.010776f
C737 B.n371 VSUBS 0.010776f
C738 B.n372 VSUBS 0.010776f
C739 B.n373 VSUBS 0.010776f
C740 B.n374 VSUBS 0.010776f
C741 B.n375 VSUBS 0.010776f
C742 B.n376 VSUBS 0.010776f
C743 B.n377 VSUBS 0.010776f
C744 B.n378 VSUBS 0.010776f
C745 B.n379 VSUBS 0.010776f
C746 B.n380 VSUBS 0.010776f
C747 B.n381 VSUBS 0.010776f
C748 B.n382 VSUBS 0.010776f
C749 B.n383 VSUBS 0.010776f
C750 B.n384 VSUBS 0.010776f
C751 B.n385 VSUBS 0.010776f
C752 B.n386 VSUBS 0.010776f
C753 B.n387 VSUBS 0.010776f
C754 B.n388 VSUBS 0.010776f
C755 B.n389 VSUBS 0.010776f
C756 B.n390 VSUBS 0.010776f
C757 B.n391 VSUBS 0.010776f
C758 B.n392 VSUBS 0.010142f
C759 B.n393 VSUBS 0.024967f
C760 B.n394 VSUBS 0.006022f
C761 B.n395 VSUBS 0.010776f
C762 B.n396 VSUBS 0.010776f
C763 B.n397 VSUBS 0.010776f
C764 B.n398 VSUBS 0.010776f
C765 B.n399 VSUBS 0.010776f
C766 B.n400 VSUBS 0.010776f
C767 B.n401 VSUBS 0.010776f
C768 B.n402 VSUBS 0.010776f
C769 B.n403 VSUBS 0.010776f
C770 B.n404 VSUBS 0.010776f
C771 B.n405 VSUBS 0.010776f
C772 B.n406 VSUBS 0.010776f
C773 B.t2 VSUBS 0.331086f
C774 B.t1 VSUBS 0.372509f
C775 B.t0 VSUBS 1.96771f
C776 B.n407 VSUBS 0.222796f
C777 B.n408 VSUBS 0.117238f
C778 B.n409 VSUBS 0.024967f
C779 B.n410 VSUBS 0.006022f
C780 B.n411 VSUBS 0.010776f
C781 B.n412 VSUBS 0.010776f
C782 B.n413 VSUBS 0.010776f
C783 B.n414 VSUBS 0.010776f
C784 B.n415 VSUBS 0.010776f
C785 B.n416 VSUBS 0.010776f
C786 B.n417 VSUBS 0.010776f
C787 B.n418 VSUBS 0.010776f
C788 B.n419 VSUBS 0.010776f
C789 B.n420 VSUBS 0.010776f
C790 B.n421 VSUBS 0.010776f
C791 B.n422 VSUBS 0.010776f
C792 B.n423 VSUBS 0.010776f
C793 B.n424 VSUBS 0.010776f
C794 B.n425 VSUBS 0.010776f
C795 B.n426 VSUBS 0.010776f
C796 B.n427 VSUBS 0.010776f
C797 B.n428 VSUBS 0.010776f
C798 B.n429 VSUBS 0.010776f
C799 B.n430 VSUBS 0.010776f
C800 B.n431 VSUBS 0.010776f
C801 B.n432 VSUBS 0.010776f
C802 B.n433 VSUBS 0.010776f
C803 B.n434 VSUBS 0.010776f
C804 B.n435 VSUBS 0.010776f
C805 B.n436 VSUBS 0.010776f
C806 B.n437 VSUBS 0.010776f
C807 B.n438 VSUBS 0.010776f
C808 B.n439 VSUBS 0.010776f
C809 B.n440 VSUBS 0.010776f
C810 B.n441 VSUBS 0.010776f
C811 B.n442 VSUBS 0.010776f
C812 B.n443 VSUBS 0.010776f
C813 B.n444 VSUBS 0.010776f
C814 B.n445 VSUBS 0.010776f
C815 B.n446 VSUBS 0.010776f
C816 B.n447 VSUBS 0.010776f
C817 B.n448 VSUBS 0.010776f
C818 B.n449 VSUBS 0.010776f
C819 B.n450 VSUBS 0.010776f
C820 B.n451 VSUBS 0.02324f
C821 B.n452 VSUBS 0.025252f
C822 B.n453 VSUBS 0.0239f
C823 B.n454 VSUBS 0.010776f
C824 B.n455 VSUBS 0.010776f
C825 B.n456 VSUBS 0.010776f
C826 B.n457 VSUBS 0.010776f
C827 B.n458 VSUBS 0.010776f
C828 B.n459 VSUBS 0.010776f
C829 B.n460 VSUBS 0.010776f
C830 B.n461 VSUBS 0.010776f
C831 B.n462 VSUBS 0.010776f
C832 B.n463 VSUBS 0.010776f
C833 B.n464 VSUBS 0.010776f
C834 B.n465 VSUBS 0.010776f
C835 B.n466 VSUBS 0.010776f
C836 B.n467 VSUBS 0.010776f
C837 B.n468 VSUBS 0.010776f
C838 B.n469 VSUBS 0.010776f
C839 B.n470 VSUBS 0.010776f
C840 B.n471 VSUBS 0.010776f
C841 B.n472 VSUBS 0.010776f
C842 B.n473 VSUBS 0.010776f
C843 B.n474 VSUBS 0.010776f
C844 B.n475 VSUBS 0.010776f
C845 B.n476 VSUBS 0.010776f
C846 B.n477 VSUBS 0.010776f
C847 B.n478 VSUBS 0.010776f
C848 B.n479 VSUBS 0.010776f
C849 B.n480 VSUBS 0.010776f
C850 B.n481 VSUBS 0.010776f
C851 B.n482 VSUBS 0.010776f
C852 B.n483 VSUBS 0.010776f
C853 B.n484 VSUBS 0.010776f
C854 B.n485 VSUBS 0.010776f
C855 B.n486 VSUBS 0.010776f
C856 B.n487 VSUBS 0.010776f
C857 B.n488 VSUBS 0.010776f
C858 B.n489 VSUBS 0.010776f
C859 B.n490 VSUBS 0.010776f
C860 B.n491 VSUBS 0.010776f
C861 B.n492 VSUBS 0.010776f
C862 B.n493 VSUBS 0.010776f
C863 B.n494 VSUBS 0.010776f
C864 B.n495 VSUBS 0.010776f
C865 B.n496 VSUBS 0.010776f
C866 B.n497 VSUBS 0.010776f
C867 B.n498 VSUBS 0.010776f
C868 B.n499 VSUBS 0.010776f
C869 B.n500 VSUBS 0.010776f
C870 B.n501 VSUBS 0.010776f
C871 B.n502 VSUBS 0.010776f
C872 B.n503 VSUBS 0.010776f
C873 B.n504 VSUBS 0.010776f
C874 B.n505 VSUBS 0.010776f
C875 B.n506 VSUBS 0.010776f
C876 B.n507 VSUBS 0.010776f
C877 B.n508 VSUBS 0.010776f
C878 B.n509 VSUBS 0.010776f
C879 B.n510 VSUBS 0.010776f
C880 B.n511 VSUBS 0.010776f
C881 B.n512 VSUBS 0.010776f
C882 B.n513 VSUBS 0.010776f
C883 B.n514 VSUBS 0.010776f
C884 B.n515 VSUBS 0.010776f
C885 B.n516 VSUBS 0.010776f
C886 B.n517 VSUBS 0.010776f
C887 B.n518 VSUBS 0.010776f
C888 B.n519 VSUBS 0.010776f
C889 B.n520 VSUBS 0.010776f
C890 B.n521 VSUBS 0.010776f
C891 B.n522 VSUBS 0.010776f
C892 B.n523 VSUBS 0.010776f
C893 B.n524 VSUBS 0.010776f
C894 B.n525 VSUBS 0.010776f
C895 B.n526 VSUBS 0.010776f
C896 B.n527 VSUBS 0.010776f
C897 B.n528 VSUBS 0.010776f
C898 B.n529 VSUBS 0.010776f
C899 B.n530 VSUBS 0.010776f
C900 B.n531 VSUBS 0.010776f
C901 B.n532 VSUBS 0.010776f
C902 B.n533 VSUBS 0.010776f
C903 B.n534 VSUBS 0.010776f
C904 B.n535 VSUBS 0.010776f
C905 B.n536 VSUBS 0.010776f
C906 B.n537 VSUBS 0.010776f
C907 B.n538 VSUBS 0.010776f
C908 B.n539 VSUBS 0.010776f
C909 B.n540 VSUBS 0.010776f
C910 B.n541 VSUBS 0.010776f
C911 B.n542 VSUBS 0.010776f
C912 B.n543 VSUBS 0.010776f
C913 B.n544 VSUBS 0.010776f
C914 B.n545 VSUBS 0.010776f
C915 B.n546 VSUBS 0.010776f
C916 B.n547 VSUBS 0.010776f
C917 B.n548 VSUBS 0.010776f
C918 B.n549 VSUBS 0.010776f
C919 B.n550 VSUBS 0.010776f
C920 B.n551 VSUBS 0.010776f
C921 B.n552 VSUBS 0.010776f
C922 B.n553 VSUBS 0.010776f
C923 B.n554 VSUBS 0.010776f
C924 B.n555 VSUBS 0.010776f
C925 B.n556 VSUBS 0.010776f
C926 B.n557 VSUBS 0.010776f
C927 B.n558 VSUBS 0.010776f
C928 B.n559 VSUBS 0.010776f
C929 B.n560 VSUBS 0.010776f
C930 B.n561 VSUBS 0.010776f
C931 B.n562 VSUBS 0.010776f
C932 B.n563 VSUBS 0.010776f
C933 B.n564 VSUBS 0.010776f
C934 B.n565 VSUBS 0.010776f
C935 B.n566 VSUBS 0.010776f
C936 B.n567 VSUBS 0.010776f
C937 B.n568 VSUBS 0.010776f
C938 B.n569 VSUBS 0.010776f
C939 B.n570 VSUBS 0.010776f
C940 B.n571 VSUBS 0.010776f
C941 B.n572 VSUBS 0.010776f
C942 B.n573 VSUBS 0.010776f
C943 B.n574 VSUBS 0.010776f
C944 B.n575 VSUBS 0.010776f
C945 B.n576 VSUBS 0.010776f
C946 B.n577 VSUBS 0.010776f
C947 B.n578 VSUBS 0.010776f
C948 B.n579 VSUBS 0.010776f
C949 B.n580 VSUBS 0.010776f
C950 B.n581 VSUBS 0.010776f
C951 B.n582 VSUBS 0.010776f
C952 B.n583 VSUBS 0.010776f
C953 B.n584 VSUBS 0.010776f
C954 B.n585 VSUBS 0.010776f
C955 B.n586 VSUBS 0.010776f
C956 B.n587 VSUBS 0.010776f
C957 B.n588 VSUBS 0.010776f
C958 B.n589 VSUBS 0.010776f
C959 B.n590 VSUBS 0.010776f
C960 B.n591 VSUBS 0.010776f
C961 B.n592 VSUBS 0.010776f
C962 B.n593 VSUBS 0.010776f
C963 B.n594 VSUBS 0.010776f
C964 B.n595 VSUBS 0.010776f
C965 B.n596 VSUBS 0.010776f
C966 B.n597 VSUBS 0.010776f
C967 B.n598 VSUBS 0.010776f
C968 B.n599 VSUBS 0.010776f
C969 B.n600 VSUBS 0.010776f
C970 B.n601 VSUBS 0.010776f
C971 B.n602 VSUBS 0.010776f
C972 B.n603 VSUBS 0.010776f
C973 B.n604 VSUBS 0.010776f
C974 B.n605 VSUBS 0.010776f
C975 B.n606 VSUBS 0.010776f
C976 B.n607 VSUBS 0.010776f
C977 B.n608 VSUBS 0.010776f
C978 B.n609 VSUBS 0.010776f
C979 B.n610 VSUBS 0.010776f
C980 B.n611 VSUBS 0.010776f
C981 B.n612 VSUBS 0.010776f
C982 B.n613 VSUBS 0.010776f
C983 B.n614 VSUBS 0.010776f
C984 B.n615 VSUBS 0.010776f
C985 B.n616 VSUBS 0.010776f
C986 B.n617 VSUBS 0.010776f
C987 B.n618 VSUBS 0.010776f
C988 B.n619 VSUBS 0.010776f
C989 B.n620 VSUBS 0.010776f
C990 B.n621 VSUBS 0.010776f
C991 B.n622 VSUBS 0.010776f
C992 B.n623 VSUBS 0.010776f
C993 B.n624 VSUBS 0.010776f
C994 B.n625 VSUBS 0.010776f
C995 B.n626 VSUBS 0.010776f
C996 B.n627 VSUBS 0.010776f
C997 B.n628 VSUBS 0.010776f
C998 B.n629 VSUBS 0.010776f
C999 B.n630 VSUBS 0.010776f
C1000 B.n631 VSUBS 0.010776f
C1001 B.n632 VSUBS 0.010776f
C1002 B.n633 VSUBS 0.010776f
C1003 B.n634 VSUBS 0.010776f
C1004 B.n635 VSUBS 0.010776f
C1005 B.n636 VSUBS 0.010776f
C1006 B.n637 VSUBS 0.010776f
C1007 B.n638 VSUBS 0.010776f
C1008 B.n639 VSUBS 0.010776f
C1009 B.n640 VSUBS 0.010776f
C1010 B.n641 VSUBS 0.010776f
C1011 B.n642 VSUBS 0.010776f
C1012 B.n643 VSUBS 0.010776f
C1013 B.n644 VSUBS 0.010776f
C1014 B.n645 VSUBS 0.010776f
C1015 B.n646 VSUBS 0.010776f
C1016 B.n647 VSUBS 0.010776f
C1017 B.n648 VSUBS 0.010776f
C1018 B.n649 VSUBS 0.010776f
C1019 B.n650 VSUBS 0.010776f
C1020 B.n651 VSUBS 0.010776f
C1021 B.n652 VSUBS 0.010776f
C1022 B.n653 VSUBS 0.010776f
C1023 B.n654 VSUBS 0.010776f
C1024 B.n655 VSUBS 0.010776f
C1025 B.n656 VSUBS 0.010776f
C1026 B.n657 VSUBS 0.010776f
C1027 B.n658 VSUBS 0.010776f
C1028 B.n659 VSUBS 0.010776f
C1029 B.n660 VSUBS 0.010776f
C1030 B.n661 VSUBS 0.010776f
C1031 B.n662 VSUBS 0.010776f
C1032 B.n663 VSUBS 0.010776f
C1033 B.n664 VSUBS 0.010776f
C1034 B.n665 VSUBS 0.010776f
C1035 B.n666 VSUBS 0.010776f
C1036 B.n667 VSUBS 0.010776f
C1037 B.n668 VSUBS 0.010776f
C1038 B.n669 VSUBS 0.010776f
C1039 B.n670 VSUBS 0.010776f
C1040 B.n671 VSUBS 0.010776f
C1041 B.n672 VSUBS 0.010776f
C1042 B.n673 VSUBS 0.010776f
C1043 B.n674 VSUBS 0.010776f
C1044 B.n675 VSUBS 0.010776f
C1045 B.n676 VSUBS 0.010776f
C1046 B.n677 VSUBS 0.010776f
C1047 B.n678 VSUBS 0.010776f
C1048 B.n679 VSUBS 0.010776f
C1049 B.n680 VSUBS 0.010776f
C1050 B.n681 VSUBS 0.010776f
C1051 B.n682 VSUBS 0.010776f
C1052 B.n683 VSUBS 0.010776f
C1053 B.n684 VSUBS 0.010776f
C1054 B.n685 VSUBS 0.010776f
C1055 B.n686 VSUBS 0.010776f
C1056 B.n687 VSUBS 0.010776f
C1057 B.n688 VSUBS 0.010776f
C1058 B.n689 VSUBS 0.010776f
C1059 B.n690 VSUBS 0.010776f
C1060 B.n691 VSUBS 0.010776f
C1061 B.n692 VSUBS 0.010776f
C1062 B.n693 VSUBS 0.010776f
C1063 B.n694 VSUBS 0.0239f
C1064 B.n695 VSUBS 0.024592f
C1065 B.n696 VSUBS 0.024592f
C1066 B.n697 VSUBS 0.010776f
C1067 B.n698 VSUBS 0.010776f
C1068 B.n699 VSUBS 0.010776f
C1069 B.n700 VSUBS 0.010776f
C1070 B.n701 VSUBS 0.010776f
C1071 B.n702 VSUBS 0.010776f
C1072 B.n703 VSUBS 0.010776f
C1073 B.n704 VSUBS 0.010776f
C1074 B.n705 VSUBS 0.010776f
C1075 B.n706 VSUBS 0.010776f
C1076 B.n707 VSUBS 0.010776f
C1077 B.n708 VSUBS 0.010776f
C1078 B.n709 VSUBS 0.010776f
C1079 B.n710 VSUBS 0.010776f
C1080 B.n711 VSUBS 0.010776f
C1081 B.n712 VSUBS 0.010776f
C1082 B.n713 VSUBS 0.010776f
C1083 B.n714 VSUBS 0.010776f
C1084 B.n715 VSUBS 0.010776f
C1085 B.n716 VSUBS 0.010776f
C1086 B.n717 VSUBS 0.010776f
C1087 B.n718 VSUBS 0.010776f
C1088 B.n719 VSUBS 0.010776f
C1089 B.n720 VSUBS 0.010776f
C1090 B.n721 VSUBS 0.010776f
C1091 B.n722 VSUBS 0.010776f
C1092 B.n723 VSUBS 0.010776f
C1093 B.n724 VSUBS 0.010776f
C1094 B.n725 VSUBS 0.010776f
C1095 B.n726 VSUBS 0.010776f
C1096 B.n727 VSUBS 0.010776f
C1097 B.n728 VSUBS 0.010776f
C1098 B.n729 VSUBS 0.010776f
C1099 B.n730 VSUBS 0.010776f
C1100 B.n731 VSUBS 0.010776f
C1101 B.n732 VSUBS 0.010776f
C1102 B.n733 VSUBS 0.010776f
C1103 B.n734 VSUBS 0.010142f
C1104 B.n735 VSUBS 0.010776f
C1105 B.n736 VSUBS 0.010776f
C1106 B.n737 VSUBS 0.010776f
C1107 B.n738 VSUBS 0.010776f
C1108 B.n739 VSUBS 0.010776f
C1109 B.n740 VSUBS 0.010776f
C1110 B.n741 VSUBS 0.010776f
C1111 B.n742 VSUBS 0.010776f
C1112 B.n743 VSUBS 0.010776f
C1113 B.n744 VSUBS 0.010776f
C1114 B.n745 VSUBS 0.010776f
C1115 B.n746 VSUBS 0.010776f
C1116 B.n747 VSUBS 0.010776f
C1117 B.n748 VSUBS 0.010776f
C1118 B.n749 VSUBS 0.010776f
C1119 B.n750 VSUBS 0.006022f
C1120 B.n751 VSUBS 0.024967f
C1121 B.n752 VSUBS 0.010142f
C1122 B.n753 VSUBS 0.010776f
C1123 B.n754 VSUBS 0.010776f
C1124 B.n755 VSUBS 0.010776f
C1125 B.n756 VSUBS 0.010776f
C1126 B.n757 VSUBS 0.010776f
C1127 B.n758 VSUBS 0.010776f
C1128 B.n759 VSUBS 0.010776f
C1129 B.n760 VSUBS 0.010776f
C1130 B.n761 VSUBS 0.010776f
C1131 B.n762 VSUBS 0.010776f
C1132 B.n763 VSUBS 0.010776f
C1133 B.n764 VSUBS 0.010776f
C1134 B.n765 VSUBS 0.010776f
C1135 B.n766 VSUBS 0.010776f
C1136 B.n767 VSUBS 0.010776f
C1137 B.n768 VSUBS 0.010776f
C1138 B.n769 VSUBS 0.010776f
C1139 B.n770 VSUBS 0.010776f
C1140 B.n771 VSUBS 0.010776f
C1141 B.n772 VSUBS 0.010776f
C1142 B.n773 VSUBS 0.010776f
C1143 B.n774 VSUBS 0.010776f
C1144 B.n775 VSUBS 0.010776f
C1145 B.n776 VSUBS 0.010776f
C1146 B.n777 VSUBS 0.010776f
C1147 B.n778 VSUBS 0.010776f
C1148 B.n779 VSUBS 0.010776f
C1149 B.n780 VSUBS 0.010776f
C1150 B.n781 VSUBS 0.010776f
C1151 B.n782 VSUBS 0.010776f
C1152 B.n783 VSUBS 0.010776f
C1153 B.n784 VSUBS 0.010776f
C1154 B.n785 VSUBS 0.010776f
C1155 B.n786 VSUBS 0.010776f
C1156 B.n787 VSUBS 0.010776f
C1157 B.n788 VSUBS 0.010776f
C1158 B.n789 VSUBS 0.010776f
C1159 B.n790 VSUBS 0.010776f
C1160 B.n791 VSUBS 0.024592f
C1161 B.n792 VSUBS 0.0239f
C1162 B.n793 VSUBS 0.0239f
C1163 B.n794 VSUBS 0.010776f
C1164 B.n795 VSUBS 0.010776f
C1165 B.n796 VSUBS 0.010776f
C1166 B.n797 VSUBS 0.010776f
C1167 B.n798 VSUBS 0.010776f
C1168 B.n799 VSUBS 0.010776f
C1169 B.n800 VSUBS 0.010776f
C1170 B.n801 VSUBS 0.010776f
C1171 B.n802 VSUBS 0.010776f
C1172 B.n803 VSUBS 0.010776f
C1173 B.n804 VSUBS 0.010776f
C1174 B.n805 VSUBS 0.010776f
C1175 B.n806 VSUBS 0.010776f
C1176 B.n807 VSUBS 0.010776f
C1177 B.n808 VSUBS 0.010776f
C1178 B.n809 VSUBS 0.010776f
C1179 B.n810 VSUBS 0.010776f
C1180 B.n811 VSUBS 0.010776f
C1181 B.n812 VSUBS 0.010776f
C1182 B.n813 VSUBS 0.010776f
C1183 B.n814 VSUBS 0.010776f
C1184 B.n815 VSUBS 0.010776f
C1185 B.n816 VSUBS 0.010776f
C1186 B.n817 VSUBS 0.010776f
C1187 B.n818 VSUBS 0.010776f
C1188 B.n819 VSUBS 0.010776f
C1189 B.n820 VSUBS 0.010776f
C1190 B.n821 VSUBS 0.010776f
C1191 B.n822 VSUBS 0.010776f
C1192 B.n823 VSUBS 0.010776f
C1193 B.n824 VSUBS 0.010776f
C1194 B.n825 VSUBS 0.010776f
C1195 B.n826 VSUBS 0.010776f
C1196 B.n827 VSUBS 0.010776f
C1197 B.n828 VSUBS 0.010776f
C1198 B.n829 VSUBS 0.010776f
C1199 B.n830 VSUBS 0.010776f
C1200 B.n831 VSUBS 0.010776f
C1201 B.n832 VSUBS 0.010776f
C1202 B.n833 VSUBS 0.010776f
C1203 B.n834 VSUBS 0.010776f
C1204 B.n835 VSUBS 0.010776f
C1205 B.n836 VSUBS 0.010776f
C1206 B.n837 VSUBS 0.010776f
C1207 B.n838 VSUBS 0.010776f
C1208 B.n839 VSUBS 0.010776f
C1209 B.n840 VSUBS 0.010776f
C1210 B.n841 VSUBS 0.010776f
C1211 B.n842 VSUBS 0.010776f
C1212 B.n843 VSUBS 0.010776f
C1213 B.n844 VSUBS 0.010776f
C1214 B.n845 VSUBS 0.010776f
C1215 B.n846 VSUBS 0.010776f
C1216 B.n847 VSUBS 0.010776f
C1217 B.n848 VSUBS 0.010776f
C1218 B.n849 VSUBS 0.010776f
C1219 B.n850 VSUBS 0.010776f
C1220 B.n851 VSUBS 0.010776f
C1221 B.n852 VSUBS 0.010776f
C1222 B.n853 VSUBS 0.010776f
C1223 B.n854 VSUBS 0.010776f
C1224 B.n855 VSUBS 0.010776f
C1225 B.n856 VSUBS 0.010776f
C1226 B.n857 VSUBS 0.010776f
C1227 B.n858 VSUBS 0.010776f
C1228 B.n859 VSUBS 0.010776f
C1229 B.n860 VSUBS 0.010776f
C1230 B.n861 VSUBS 0.010776f
C1231 B.n862 VSUBS 0.010776f
C1232 B.n863 VSUBS 0.010776f
C1233 B.n864 VSUBS 0.010776f
C1234 B.n865 VSUBS 0.010776f
C1235 B.n866 VSUBS 0.010776f
C1236 B.n867 VSUBS 0.010776f
C1237 B.n868 VSUBS 0.010776f
C1238 B.n869 VSUBS 0.010776f
C1239 B.n870 VSUBS 0.010776f
C1240 B.n871 VSUBS 0.010776f
C1241 B.n872 VSUBS 0.010776f
C1242 B.n873 VSUBS 0.010776f
C1243 B.n874 VSUBS 0.010776f
C1244 B.n875 VSUBS 0.010776f
C1245 B.n876 VSUBS 0.010776f
C1246 B.n877 VSUBS 0.010776f
C1247 B.n878 VSUBS 0.010776f
C1248 B.n879 VSUBS 0.010776f
C1249 B.n880 VSUBS 0.010776f
C1250 B.n881 VSUBS 0.010776f
C1251 B.n882 VSUBS 0.010776f
C1252 B.n883 VSUBS 0.010776f
C1253 B.n884 VSUBS 0.010776f
C1254 B.n885 VSUBS 0.010776f
C1255 B.n886 VSUBS 0.010776f
C1256 B.n887 VSUBS 0.010776f
C1257 B.n888 VSUBS 0.010776f
C1258 B.n889 VSUBS 0.010776f
C1259 B.n890 VSUBS 0.010776f
C1260 B.n891 VSUBS 0.010776f
C1261 B.n892 VSUBS 0.010776f
C1262 B.n893 VSUBS 0.010776f
C1263 B.n894 VSUBS 0.010776f
C1264 B.n895 VSUBS 0.010776f
C1265 B.n896 VSUBS 0.010776f
C1266 B.n897 VSUBS 0.010776f
C1267 B.n898 VSUBS 0.010776f
C1268 B.n899 VSUBS 0.010776f
C1269 B.n900 VSUBS 0.010776f
C1270 B.n901 VSUBS 0.010776f
C1271 B.n902 VSUBS 0.010776f
C1272 B.n903 VSUBS 0.010776f
C1273 B.n904 VSUBS 0.010776f
C1274 B.n905 VSUBS 0.010776f
C1275 B.n906 VSUBS 0.010776f
C1276 B.n907 VSUBS 0.010776f
C1277 B.n908 VSUBS 0.010776f
C1278 B.n909 VSUBS 0.010776f
C1279 B.n910 VSUBS 0.010776f
C1280 B.n911 VSUBS 0.014062f
C1281 B.n912 VSUBS 0.01498f
C1282 B.n913 VSUBS 0.029789f
.ends

