* NGSPICE file created from diff_pair_sample_1280.ext - technology: sky130A

.subckt diff_pair_sample_1280 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=2.19285 ps=13.62 w=13.29 l=2.73
X1 VTAIL.t13 VP.t1 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X2 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X3 VTAIL.t12 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=2.19285 ps=13.62 w=13.29 l=2.73
X4 VDD1.t1 VP.t3 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X5 VDD2.t6 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X6 VDD2.t5 VN.t2 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=5.1831 ps=27.36 w=13.29 l=2.73
X7 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=2.73
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=2.73
X9 VDD1.t0 VP.t4 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=5.1831 ps=27.36 w=13.29 l=2.73
X10 VDD1.t4 VP.t5 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X11 VTAIL.t2 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=2.19285 ps=13.62 w=13.29 l=2.73
X12 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=5.1831 ps=27.36 w=13.29 l=2.73
X13 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=2.19285 ps=13.62 w=13.29 l=2.73
X14 VTAIL.t8 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=2.73
X16 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=5.1831 ps=27.36 w=13.29 l=2.73
X17 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X18 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.19285 pd=13.62 as=2.19285 ps=13.62 w=13.29 l=2.73
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1831 pd=27.36 as=0 ps=0 w=13.29 l=2.73
R0 VP.n21 VP.n20 161.3
R1 VP.n22 VP.n17 161.3
R2 VP.n24 VP.n23 161.3
R3 VP.n25 VP.n16 161.3
R4 VP.n27 VP.n26 161.3
R5 VP.n28 VP.n15 161.3
R6 VP.n30 VP.n29 161.3
R7 VP.n32 VP.n31 161.3
R8 VP.n33 VP.n13 161.3
R9 VP.n35 VP.n34 161.3
R10 VP.n36 VP.n12 161.3
R11 VP.n38 VP.n37 161.3
R12 VP.n39 VP.n11 161.3
R13 VP.n72 VP.n0 161.3
R14 VP.n71 VP.n70 161.3
R15 VP.n69 VP.n1 161.3
R16 VP.n68 VP.n67 161.3
R17 VP.n66 VP.n2 161.3
R18 VP.n65 VP.n64 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n61 VP.n4 161.3
R21 VP.n60 VP.n59 161.3
R22 VP.n58 VP.n5 161.3
R23 VP.n57 VP.n56 161.3
R24 VP.n55 VP.n6 161.3
R25 VP.n54 VP.n53 161.3
R26 VP.n52 VP.n51 161.3
R27 VP.n50 VP.n8 161.3
R28 VP.n49 VP.n48 161.3
R29 VP.n47 VP.n9 161.3
R30 VP.n46 VP.n45 161.3
R31 VP.n44 VP.n10 161.3
R32 VP.n19 VP.t0 148.993
R33 VP.n43 VP.t2 117.323
R34 VP.n7 VP.t5 117.323
R35 VP.n3 VP.t1 117.323
R36 VP.n73 VP.t4 117.323
R37 VP.n40 VP.t7 117.323
R38 VP.n14 VP.t6 117.323
R39 VP.n18 VP.t3 117.323
R40 VP.n43 VP.n42 106.353
R41 VP.n74 VP.n73 106.353
R42 VP.n41 VP.n40 106.353
R43 VP.n19 VP.n18 71.7459
R44 VP.n42 VP.n41 52.4466
R45 VP.n49 VP.n9 46.321
R46 VP.n67 VP.n1 46.321
R47 VP.n34 VP.n12 46.321
R48 VP.n56 VP.n5 40.4934
R49 VP.n60 VP.n5 40.4934
R50 VP.n27 VP.n16 40.4934
R51 VP.n23 VP.n16 40.4934
R52 VP.n50 VP.n49 34.6658
R53 VP.n67 VP.n66 34.6658
R54 VP.n34 VP.n33 34.6658
R55 VP.n45 VP.n44 24.4675
R56 VP.n45 VP.n9 24.4675
R57 VP.n51 VP.n50 24.4675
R58 VP.n55 VP.n54 24.4675
R59 VP.n56 VP.n55 24.4675
R60 VP.n61 VP.n60 24.4675
R61 VP.n62 VP.n61 24.4675
R62 VP.n66 VP.n65 24.4675
R63 VP.n71 VP.n1 24.4675
R64 VP.n72 VP.n71 24.4675
R65 VP.n38 VP.n12 24.4675
R66 VP.n39 VP.n38 24.4675
R67 VP.n28 VP.n27 24.4675
R68 VP.n29 VP.n28 24.4675
R69 VP.n33 VP.n32 24.4675
R70 VP.n22 VP.n21 24.4675
R71 VP.n23 VP.n22 24.4675
R72 VP.n51 VP.n7 22.9995
R73 VP.n65 VP.n3 22.9995
R74 VP.n32 VP.n14 22.9995
R75 VP.n20 VP.n19 7.21203
R76 VP.n44 VP.n43 4.40456
R77 VP.n73 VP.n72 4.40456
R78 VP.n40 VP.n39 4.40456
R79 VP.n54 VP.n7 1.46852
R80 VP.n62 VP.n3 1.46852
R81 VP.n29 VP.n14 1.46852
R82 VP.n21 VP.n18 1.46852
R83 VP.n41 VP.n11 0.278367
R84 VP.n42 VP.n10 0.278367
R85 VP.n74 VP.n0 0.278367
R86 VP.n20 VP.n17 0.189894
R87 VP.n24 VP.n17 0.189894
R88 VP.n25 VP.n24 0.189894
R89 VP.n26 VP.n25 0.189894
R90 VP.n26 VP.n15 0.189894
R91 VP.n30 VP.n15 0.189894
R92 VP.n31 VP.n30 0.189894
R93 VP.n31 VP.n13 0.189894
R94 VP.n35 VP.n13 0.189894
R95 VP.n36 VP.n35 0.189894
R96 VP.n37 VP.n36 0.189894
R97 VP.n37 VP.n11 0.189894
R98 VP.n46 VP.n10 0.189894
R99 VP.n47 VP.n46 0.189894
R100 VP.n48 VP.n47 0.189894
R101 VP.n48 VP.n8 0.189894
R102 VP.n52 VP.n8 0.189894
R103 VP.n53 VP.n52 0.189894
R104 VP.n53 VP.n6 0.189894
R105 VP.n57 VP.n6 0.189894
R106 VP.n58 VP.n57 0.189894
R107 VP.n59 VP.n58 0.189894
R108 VP.n59 VP.n4 0.189894
R109 VP.n63 VP.n4 0.189894
R110 VP.n64 VP.n63 0.189894
R111 VP.n64 VP.n2 0.189894
R112 VP.n68 VP.n2 0.189894
R113 VP.n69 VP.n68 0.189894
R114 VP.n70 VP.n69 0.189894
R115 VP.n70 VP.n0 0.189894
R116 VP VP.n74 0.153454
R117 VDD1 VDD1.n0 64.2422
R118 VDD1.n3 VDD1.n2 64.1285
R119 VDD1.n3 VDD1.n1 64.1285
R120 VDD1.n5 VDD1.n4 62.8649
R121 VDD1.n5 VDD1.n3 47.6259
R122 VDD1.n4 VDD1.t3 1.49034
R123 VDD1.n4 VDD1.t2 1.49034
R124 VDD1.n0 VDD1.t7 1.49034
R125 VDD1.n0 VDD1.t1 1.49034
R126 VDD1.n2 VDD1.t6 1.49034
R127 VDD1.n2 VDD1.t0 1.49034
R128 VDD1.n1 VDD1.t5 1.49034
R129 VDD1.n1 VDD1.t4 1.49034
R130 VDD1 VDD1.n5 1.26128
R131 VTAIL.n578 VTAIL.n512 214.453
R132 VTAIL.n68 VTAIL.n2 214.453
R133 VTAIL.n140 VTAIL.n74 214.453
R134 VTAIL.n214 VTAIL.n148 214.453
R135 VTAIL.n506 VTAIL.n440 214.453
R136 VTAIL.n432 VTAIL.n366 214.453
R137 VTAIL.n360 VTAIL.n294 214.453
R138 VTAIL.n286 VTAIL.n220 214.453
R139 VTAIL.n537 VTAIL.n536 185
R140 VTAIL.n539 VTAIL.n538 185
R141 VTAIL.n532 VTAIL.n531 185
R142 VTAIL.n545 VTAIL.n544 185
R143 VTAIL.n547 VTAIL.n546 185
R144 VTAIL.n528 VTAIL.n527 185
R145 VTAIL.n553 VTAIL.n552 185
R146 VTAIL.n555 VTAIL.n554 185
R147 VTAIL.n524 VTAIL.n523 185
R148 VTAIL.n561 VTAIL.n560 185
R149 VTAIL.n563 VTAIL.n562 185
R150 VTAIL.n520 VTAIL.n519 185
R151 VTAIL.n569 VTAIL.n568 185
R152 VTAIL.n571 VTAIL.n570 185
R153 VTAIL.n516 VTAIL.n515 185
R154 VTAIL.n577 VTAIL.n576 185
R155 VTAIL.n579 VTAIL.n578 185
R156 VTAIL.n27 VTAIL.n26 185
R157 VTAIL.n29 VTAIL.n28 185
R158 VTAIL.n22 VTAIL.n21 185
R159 VTAIL.n35 VTAIL.n34 185
R160 VTAIL.n37 VTAIL.n36 185
R161 VTAIL.n18 VTAIL.n17 185
R162 VTAIL.n43 VTAIL.n42 185
R163 VTAIL.n45 VTAIL.n44 185
R164 VTAIL.n14 VTAIL.n13 185
R165 VTAIL.n51 VTAIL.n50 185
R166 VTAIL.n53 VTAIL.n52 185
R167 VTAIL.n10 VTAIL.n9 185
R168 VTAIL.n59 VTAIL.n58 185
R169 VTAIL.n61 VTAIL.n60 185
R170 VTAIL.n6 VTAIL.n5 185
R171 VTAIL.n67 VTAIL.n66 185
R172 VTAIL.n69 VTAIL.n68 185
R173 VTAIL.n99 VTAIL.n98 185
R174 VTAIL.n101 VTAIL.n100 185
R175 VTAIL.n94 VTAIL.n93 185
R176 VTAIL.n107 VTAIL.n106 185
R177 VTAIL.n109 VTAIL.n108 185
R178 VTAIL.n90 VTAIL.n89 185
R179 VTAIL.n115 VTAIL.n114 185
R180 VTAIL.n117 VTAIL.n116 185
R181 VTAIL.n86 VTAIL.n85 185
R182 VTAIL.n123 VTAIL.n122 185
R183 VTAIL.n125 VTAIL.n124 185
R184 VTAIL.n82 VTAIL.n81 185
R185 VTAIL.n131 VTAIL.n130 185
R186 VTAIL.n133 VTAIL.n132 185
R187 VTAIL.n78 VTAIL.n77 185
R188 VTAIL.n139 VTAIL.n138 185
R189 VTAIL.n141 VTAIL.n140 185
R190 VTAIL.n173 VTAIL.n172 185
R191 VTAIL.n175 VTAIL.n174 185
R192 VTAIL.n168 VTAIL.n167 185
R193 VTAIL.n181 VTAIL.n180 185
R194 VTAIL.n183 VTAIL.n182 185
R195 VTAIL.n164 VTAIL.n163 185
R196 VTAIL.n189 VTAIL.n188 185
R197 VTAIL.n191 VTAIL.n190 185
R198 VTAIL.n160 VTAIL.n159 185
R199 VTAIL.n197 VTAIL.n196 185
R200 VTAIL.n199 VTAIL.n198 185
R201 VTAIL.n156 VTAIL.n155 185
R202 VTAIL.n205 VTAIL.n204 185
R203 VTAIL.n207 VTAIL.n206 185
R204 VTAIL.n152 VTAIL.n151 185
R205 VTAIL.n213 VTAIL.n212 185
R206 VTAIL.n215 VTAIL.n214 185
R207 VTAIL.n507 VTAIL.n506 185
R208 VTAIL.n505 VTAIL.n504 185
R209 VTAIL.n444 VTAIL.n443 185
R210 VTAIL.n499 VTAIL.n498 185
R211 VTAIL.n497 VTAIL.n496 185
R212 VTAIL.n448 VTAIL.n447 185
R213 VTAIL.n491 VTAIL.n490 185
R214 VTAIL.n489 VTAIL.n488 185
R215 VTAIL.n452 VTAIL.n451 185
R216 VTAIL.n483 VTAIL.n482 185
R217 VTAIL.n481 VTAIL.n480 185
R218 VTAIL.n456 VTAIL.n455 185
R219 VTAIL.n475 VTAIL.n474 185
R220 VTAIL.n473 VTAIL.n472 185
R221 VTAIL.n460 VTAIL.n459 185
R222 VTAIL.n467 VTAIL.n466 185
R223 VTAIL.n465 VTAIL.n464 185
R224 VTAIL.n433 VTAIL.n432 185
R225 VTAIL.n431 VTAIL.n430 185
R226 VTAIL.n370 VTAIL.n369 185
R227 VTAIL.n425 VTAIL.n424 185
R228 VTAIL.n423 VTAIL.n422 185
R229 VTAIL.n374 VTAIL.n373 185
R230 VTAIL.n417 VTAIL.n416 185
R231 VTAIL.n415 VTAIL.n414 185
R232 VTAIL.n378 VTAIL.n377 185
R233 VTAIL.n409 VTAIL.n408 185
R234 VTAIL.n407 VTAIL.n406 185
R235 VTAIL.n382 VTAIL.n381 185
R236 VTAIL.n401 VTAIL.n400 185
R237 VTAIL.n399 VTAIL.n398 185
R238 VTAIL.n386 VTAIL.n385 185
R239 VTAIL.n393 VTAIL.n392 185
R240 VTAIL.n391 VTAIL.n390 185
R241 VTAIL.n361 VTAIL.n360 185
R242 VTAIL.n359 VTAIL.n358 185
R243 VTAIL.n298 VTAIL.n297 185
R244 VTAIL.n353 VTAIL.n352 185
R245 VTAIL.n351 VTAIL.n350 185
R246 VTAIL.n302 VTAIL.n301 185
R247 VTAIL.n345 VTAIL.n344 185
R248 VTAIL.n343 VTAIL.n342 185
R249 VTAIL.n306 VTAIL.n305 185
R250 VTAIL.n337 VTAIL.n336 185
R251 VTAIL.n335 VTAIL.n334 185
R252 VTAIL.n310 VTAIL.n309 185
R253 VTAIL.n329 VTAIL.n328 185
R254 VTAIL.n327 VTAIL.n326 185
R255 VTAIL.n314 VTAIL.n313 185
R256 VTAIL.n321 VTAIL.n320 185
R257 VTAIL.n319 VTAIL.n318 185
R258 VTAIL.n287 VTAIL.n286 185
R259 VTAIL.n285 VTAIL.n284 185
R260 VTAIL.n224 VTAIL.n223 185
R261 VTAIL.n279 VTAIL.n278 185
R262 VTAIL.n277 VTAIL.n276 185
R263 VTAIL.n228 VTAIL.n227 185
R264 VTAIL.n271 VTAIL.n270 185
R265 VTAIL.n269 VTAIL.n268 185
R266 VTAIL.n232 VTAIL.n231 185
R267 VTAIL.n263 VTAIL.n262 185
R268 VTAIL.n261 VTAIL.n260 185
R269 VTAIL.n236 VTAIL.n235 185
R270 VTAIL.n255 VTAIL.n254 185
R271 VTAIL.n253 VTAIL.n252 185
R272 VTAIL.n240 VTAIL.n239 185
R273 VTAIL.n247 VTAIL.n246 185
R274 VTAIL.n245 VTAIL.n244 185
R275 VTAIL.n535 VTAIL.t15 147.659
R276 VTAIL.n25 VTAIL.t2 147.659
R277 VTAIL.n97 VTAIL.t10 147.659
R278 VTAIL.n171 VTAIL.t12 147.659
R279 VTAIL.n463 VTAIL.t7 147.659
R280 VTAIL.n389 VTAIL.t14 147.659
R281 VTAIL.n317 VTAIL.t0 147.659
R282 VTAIL.n243 VTAIL.t1 147.659
R283 VTAIL.n538 VTAIL.n537 104.615
R284 VTAIL.n538 VTAIL.n531 104.615
R285 VTAIL.n545 VTAIL.n531 104.615
R286 VTAIL.n546 VTAIL.n545 104.615
R287 VTAIL.n546 VTAIL.n527 104.615
R288 VTAIL.n553 VTAIL.n527 104.615
R289 VTAIL.n554 VTAIL.n553 104.615
R290 VTAIL.n554 VTAIL.n523 104.615
R291 VTAIL.n561 VTAIL.n523 104.615
R292 VTAIL.n562 VTAIL.n561 104.615
R293 VTAIL.n562 VTAIL.n519 104.615
R294 VTAIL.n569 VTAIL.n519 104.615
R295 VTAIL.n570 VTAIL.n569 104.615
R296 VTAIL.n570 VTAIL.n515 104.615
R297 VTAIL.n577 VTAIL.n515 104.615
R298 VTAIL.n578 VTAIL.n577 104.615
R299 VTAIL.n28 VTAIL.n27 104.615
R300 VTAIL.n28 VTAIL.n21 104.615
R301 VTAIL.n35 VTAIL.n21 104.615
R302 VTAIL.n36 VTAIL.n35 104.615
R303 VTAIL.n36 VTAIL.n17 104.615
R304 VTAIL.n43 VTAIL.n17 104.615
R305 VTAIL.n44 VTAIL.n43 104.615
R306 VTAIL.n44 VTAIL.n13 104.615
R307 VTAIL.n51 VTAIL.n13 104.615
R308 VTAIL.n52 VTAIL.n51 104.615
R309 VTAIL.n52 VTAIL.n9 104.615
R310 VTAIL.n59 VTAIL.n9 104.615
R311 VTAIL.n60 VTAIL.n59 104.615
R312 VTAIL.n60 VTAIL.n5 104.615
R313 VTAIL.n67 VTAIL.n5 104.615
R314 VTAIL.n68 VTAIL.n67 104.615
R315 VTAIL.n100 VTAIL.n99 104.615
R316 VTAIL.n100 VTAIL.n93 104.615
R317 VTAIL.n107 VTAIL.n93 104.615
R318 VTAIL.n108 VTAIL.n107 104.615
R319 VTAIL.n108 VTAIL.n89 104.615
R320 VTAIL.n115 VTAIL.n89 104.615
R321 VTAIL.n116 VTAIL.n115 104.615
R322 VTAIL.n116 VTAIL.n85 104.615
R323 VTAIL.n123 VTAIL.n85 104.615
R324 VTAIL.n124 VTAIL.n123 104.615
R325 VTAIL.n124 VTAIL.n81 104.615
R326 VTAIL.n131 VTAIL.n81 104.615
R327 VTAIL.n132 VTAIL.n131 104.615
R328 VTAIL.n132 VTAIL.n77 104.615
R329 VTAIL.n139 VTAIL.n77 104.615
R330 VTAIL.n140 VTAIL.n139 104.615
R331 VTAIL.n174 VTAIL.n173 104.615
R332 VTAIL.n174 VTAIL.n167 104.615
R333 VTAIL.n181 VTAIL.n167 104.615
R334 VTAIL.n182 VTAIL.n181 104.615
R335 VTAIL.n182 VTAIL.n163 104.615
R336 VTAIL.n189 VTAIL.n163 104.615
R337 VTAIL.n190 VTAIL.n189 104.615
R338 VTAIL.n190 VTAIL.n159 104.615
R339 VTAIL.n197 VTAIL.n159 104.615
R340 VTAIL.n198 VTAIL.n197 104.615
R341 VTAIL.n198 VTAIL.n155 104.615
R342 VTAIL.n205 VTAIL.n155 104.615
R343 VTAIL.n206 VTAIL.n205 104.615
R344 VTAIL.n206 VTAIL.n151 104.615
R345 VTAIL.n213 VTAIL.n151 104.615
R346 VTAIL.n214 VTAIL.n213 104.615
R347 VTAIL.n506 VTAIL.n505 104.615
R348 VTAIL.n505 VTAIL.n443 104.615
R349 VTAIL.n498 VTAIL.n443 104.615
R350 VTAIL.n498 VTAIL.n497 104.615
R351 VTAIL.n497 VTAIL.n447 104.615
R352 VTAIL.n490 VTAIL.n447 104.615
R353 VTAIL.n490 VTAIL.n489 104.615
R354 VTAIL.n489 VTAIL.n451 104.615
R355 VTAIL.n482 VTAIL.n451 104.615
R356 VTAIL.n482 VTAIL.n481 104.615
R357 VTAIL.n481 VTAIL.n455 104.615
R358 VTAIL.n474 VTAIL.n455 104.615
R359 VTAIL.n474 VTAIL.n473 104.615
R360 VTAIL.n473 VTAIL.n459 104.615
R361 VTAIL.n466 VTAIL.n459 104.615
R362 VTAIL.n466 VTAIL.n465 104.615
R363 VTAIL.n432 VTAIL.n431 104.615
R364 VTAIL.n431 VTAIL.n369 104.615
R365 VTAIL.n424 VTAIL.n369 104.615
R366 VTAIL.n424 VTAIL.n423 104.615
R367 VTAIL.n423 VTAIL.n373 104.615
R368 VTAIL.n416 VTAIL.n373 104.615
R369 VTAIL.n416 VTAIL.n415 104.615
R370 VTAIL.n415 VTAIL.n377 104.615
R371 VTAIL.n408 VTAIL.n377 104.615
R372 VTAIL.n408 VTAIL.n407 104.615
R373 VTAIL.n407 VTAIL.n381 104.615
R374 VTAIL.n400 VTAIL.n381 104.615
R375 VTAIL.n400 VTAIL.n399 104.615
R376 VTAIL.n399 VTAIL.n385 104.615
R377 VTAIL.n392 VTAIL.n385 104.615
R378 VTAIL.n392 VTAIL.n391 104.615
R379 VTAIL.n360 VTAIL.n359 104.615
R380 VTAIL.n359 VTAIL.n297 104.615
R381 VTAIL.n352 VTAIL.n297 104.615
R382 VTAIL.n352 VTAIL.n351 104.615
R383 VTAIL.n351 VTAIL.n301 104.615
R384 VTAIL.n344 VTAIL.n301 104.615
R385 VTAIL.n344 VTAIL.n343 104.615
R386 VTAIL.n343 VTAIL.n305 104.615
R387 VTAIL.n336 VTAIL.n305 104.615
R388 VTAIL.n336 VTAIL.n335 104.615
R389 VTAIL.n335 VTAIL.n309 104.615
R390 VTAIL.n328 VTAIL.n309 104.615
R391 VTAIL.n328 VTAIL.n327 104.615
R392 VTAIL.n327 VTAIL.n313 104.615
R393 VTAIL.n320 VTAIL.n313 104.615
R394 VTAIL.n320 VTAIL.n319 104.615
R395 VTAIL.n286 VTAIL.n285 104.615
R396 VTAIL.n285 VTAIL.n223 104.615
R397 VTAIL.n278 VTAIL.n223 104.615
R398 VTAIL.n278 VTAIL.n277 104.615
R399 VTAIL.n277 VTAIL.n227 104.615
R400 VTAIL.n270 VTAIL.n227 104.615
R401 VTAIL.n270 VTAIL.n269 104.615
R402 VTAIL.n269 VTAIL.n231 104.615
R403 VTAIL.n262 VTAIL.n231 104.615
R404 VTAIL.n262 VTAIL.n261 104.615
R405 VTAIL.n261 VTAIL.n235 104.615
R406 VTAIL.n254 VTAIL.n235 104.615
R407 VTAIL.n254 VTAIL.n253 104.615
R408 VTAIL.n253 VTAIL.n239 104.615
R409 VTAIL.n246 VTAIL.n239 104.615
R410 VTAIL.n246 VTAIL.n245 104.615
R411 VTAIL.n537 VTAIL.t15 52.3082
R412 VTAIL.n27 VTAIL.t2 52.3082
R413 VTAIL.n99 VTAIL.t10 52.3082
R414 VTAIL.n173 VTAIL.t12 52.3082
R415 VTAIL.n465 VTAIL.t7 52.3082
R416 VTAIL.n391 VTAIL.t14 52.3082
R417 VTAIL.n319 VTAIL.t0 52.3082
R418 VTAIL.n245 VTAIL.t1 52.3082
R419 VTAIL.n439 VTAIL.n438 46.1863
R420 VTAIL.n293 VTAIL.n292 46.1863
R421 VTAIL.n1 VTAIL.n0 46.1861
R422 VTAIL.n147 VTAIL.n146 46.1861
R423 VTAIL.n583 VTAIL.n582 33.9308
R424 VTAIL.n73 VTAIL.n72 33.9308
R425 VTAIL.n145 VTAIL.n144 33.9308
R426 VTAIL.n219 VTAIL.n218 33.9308
R427 VTAIL.n511 VTAIL.n510 33.9308
R428 VTAIL.n437 VTAIL.n436 33.9308
R429 VTAIL.n365 VTAIL.n364 33.9308
R430 VTAIL.n291 VTAIL.n290 33.9308
R431 VTAIL.n583 VTAIL.n511 26.4617
R432 VTAIL.n291 VTAIL.n219 26.4617
R433 VTAIL.n536 VTAIL.n535 15.6677
R434 VTAIL.n26 VTAIL.n25 15.6677
R435 VTAIL.n98 VTAIL.n97 15.6677
R436 VTAIL.n172 VTAIL.n171 15.6677
R437 VTAIL.n464 VTAIL.n463 15.6677
R438 VTAIL.n390 VTAIL.n389 15.6677
R439 VTAIL.n318 VTAIL.n317 15.6677
R440 VTAIL.n244 VTAIL.n243 15.6677
R441 VTAIL.n539 VTAIL.n534 12.8005
R442 VTAIL.n580 VTAIL.n579 12.8005
R443 VTAIL.n29 VTAIL.n24 12.8005
R444 VTAIL.n70 VTAIL.n69 12.8005
R445 VTAIL.n101 VTAIL.n96 12.8005
R446 VTAIL.n142 VTAIL.n141 12.8005
R447 VTAIL.n175 VTAIL.n170 12.8005
R448 VTAIL.n216 VTAIL.n215 12.8005
R449 VTAIL.n508 VTAIL.n507 12.8005
R450 VTAIL.n467 VTAIL.n462 12.8005
R451 VTAIL.n434 VTAIL.n433 12.8005
R452 VTAIL.n393 VTAIL.n388 12.8005
R453 VTAIL.n362 VTAIL.n361 12.8005
R454 VTAIL.n321 VTAIL.n316 12.8005
R455 VTAIL.n288 VTAIL.n287 12.8005
R456 VTAIL.n247 VTAIL.n242 12.8005
R457 VTAIL.n540 VTAIL.n532 12.0247
R458 VTAIL.n576 VTAIL.n514 12.0247
R459 VTAIL.n30 VTAIL.n22 12.0247
R460 VTAIL.n66 VTAIL.n4 12.0247
R461 VTAIL.n102 VTAIL.n94 12.0247
R462 VTAIL.n138 VTAIL.n76 12.0247
R463 VTAIL.n176 VTAIL.n168 12.0247
R464 VTAIL.n212 VTAIL.n150 12.0247
R465 VTAIL.n504 VTAIL.n442 12.0247
R466 VTAIL.n468 VTAIL.n460 12.0247
R467 VTAIL.n430 VTAIL.n368 12.0247
R468 VTAIL.n394 VTAIL.n386 12.0247
R469 VTAIL.n358 VTAIL.n296 12.0247
R470 VTAIL.n322 VTAIL.n314 12.0247
R471 VTAIL.n284 VTAIL.n222 12.0247
R472 VTAIL.n248 VTAIL.n240 12.0247
R473 VTAIL.n544 VTAIL.n543 11.249
R474 VTAIL.n575 VTAIL.n516 11.249
R475 VTAIL.n34 VTAIL.n33 11.249
R476 VTAIL.n65 VTAIL.n6 11.249
R477 VTAIL.n106 VTAIL.n105 11.249
R478 VTAIL.n137 VTAIL.n78 11.249
R479 VTAIL.n180 VTAIL.n179 11.249
R480 VTAIL.n211 VTAIL.n152 11.249
R481 VTAIL.n503 VTAIL.n444 11.249
R482 VTAIL.n472 VTAIL.n471 11.249
R483 VTAIL.n429 VTAIL.n370 11.249
R484 VTAIL.n398 VTAIL.n397 11.249
R485 VTAIL.n357 VTAIL.n298 11.249
R486 VTAIL.n326 VTAIL.n325 11.249
R487 VTAIL.n283 VTAIL.n224 11.249
R488 VTAIL.n252 VTAIL.n251 11.249
R489 VTAIL.n547 VTAIL.n530 10.4732
R490 VTAIL.n572 VTAIL.n571 10.4732
R491 VTAIL.n37 VTAIL.n20 10.4732
R492 VTAIL.n62 VTAIL.n61 10.4732
R493 VTAIL.n109 VTAIL.n92 10.4732
R494 VTAIL.n134 VTAIL.n133 10.4732
R495 VTAIL.n183 VTAIL.n166 10.4732
R496 VTAIL.n208 VTAIL.n207 10.4732
R497 VTAIL.n500 VTAIL.n499 10.4732
R498 VTAIL.n475 VTAIL.n458 10.4732
R499 VTAIL.n426 VTAIL.n425 10.4732
R500 VTAIL.n401 VTAIL.n384 10.4732
R501 VTAIL.n354 VTAIL.n353 10.4732
R502 VTAIL.n329 VTAIL.n312 10.4732
R503 VTAIL.n280 VTAIL.n279 10.4732
R504 VTAIL.n255 VTAIL.n238 10.4732
R505 VTAIL.n548 VTAIL.n528 9.69747
R506 VTAIL.n568 VTAIL.n518 9.69747
R507 VTAIL.n38 VTAIL.n18 9.69747
R508 VTAIL.n58 VTAIL.n8 9.69747
R509 VTAIL.n110 VTAIL.n90 9.69747
R510 VTAIL.n130 VTAIL.n80 9.69747
R511 VTAIL.n184 VTAIL.n164 9.69747
R512 VTAIL.n204 VTAIL.n154 9.69747
R513 VTAIL.n496 VTAIL.n446 9.69747
R514 VTAIL.n476 VTAIL.n456 9.69747
R515 VTAIL.n422 VTAIL.n372 9.69747
R516 VTAIL.n402 VTAIL.n382 9.69747
R517 VTAIL.n350 VTAIL.n300 9.69747
R518 VTAIL.n330 VTAIL.n310 9.69747
R519 VTAIL.n276 VTAIL.n226 9.69747
R520 VTAIL.n256 VTAIL.n236 9.69747
R521 VTAIL.n582 VTAIL.n581 9.45567
R522 VTAIL.n72 VTAIL.n71 9.45567
R523 VTAIL.n144 VTAIL.n143 9.45567
R524 VTAIL.n218 VTAIL.n217 9.45567
R525 VTAIL.n510 VTAIL.n509 9.45567
R526 VTAIL.n436 VTAIL.n435 9.45567
R527 VTAIL.n364 VTAIL.n363 9.45567
R528 VTAIL.n290 VTAIL.n289 9.45567
R529 VTAIL.n557 VTAIL.n556 9.3005
R530 VTAIL.n526 VTAIL.n525 9.3005
R531 VTAIL.n551 VTAIL.n550 9.3005
R532 VTAIL.n549 VTAIL.n548 9.3005
R533 VTAIL.n530 VTAIL.n529 9.3005
R534 VTAIL.n543 VTAIL.n542 9.3005
R535 VTAIL.n541 VTAIL.n540 9.3005
R536 VTAIL.n534 VTAIL.n533 9.3005
R537 VTAIL.n559 VTAIL.n558 9.3005
R538 VTAIL.n522 VTAIL.n521 9.3005
R539 VTAIL.n565 VTAIL.n564 9.3005
R540 VTAIL.n567 VTAIL.n566 9.3005
R541 VTAIL.n518 VTAIL.n517 9.3005
R542 VTAIL.n573 VTAIL.n572 9.3005
R543 VTAIL.n575 VTAIL.n574 9.3005
R544 VTAIL.n514 VTAIL.n513 9.3005
R545 VTAIL.n581 VTAIL.n580 9.3005
R546 VTAIL.n47 VTAIL.n46 9.3005
R547 VTAIL.n16 VTAIL.n15 9.3005
R548 VTAIL.n41 VTAIL.n40 9.3005
R549 VTAIL.n39 VTAIL.n38 9.3005
R550 VTAIL.n20 VTAIL.n19 9.3005
R551 VTAIL.n33 VTAIL.n32 9.3005
R552 VTAIL.n31 VTAIL.n30 9.3005
R553 VTAIL.n24 VTAIL.n23 9.3005
R554 VTAIL.n49 VTAIL.n48 9.3005
R555 VTAIL.n12 VTAIL.n11 9.3005
R556 VTAIL.n55 VTAIL.n54 9.3005
R557 VTAIL.n57 VTAIL.n56 9.3005
R558 VTAIL.n8 VTAIL.n7 9.3005
R559 VTAIL.n63 VTAIL.n62 9.3005
R560 VTAIL.n65 VTAIL.n64 9.3005
R561 VTAIL.n4 VTAIL.n3 9.3005
R562 VTAIL.n71 VTAIL.n70 9.3005
R563 VTAIL.n119 VTAIL.n118 9.3005
R564 VTAIL.n88 VTAIL.n87 9.3005
R565 VTAIL.n113 VTAIL.n112 9.3005
R566 VTAIL.n111 VTAIL.n110 9.3005
R567 VTAIL.n92 VTAIL.n91 9.3005
R568 VTAIL.n105 VTAIL.n104 9.3005
R569 VTAIL.n103 VTAIL.n102 9.3005
R570 VTAIL.n96 VTAIL.n95 9.3005
R571 VTAIL.n121 VTAIL.n120 9.3005
R572 VTAIL.n84 VTAIL.n83 9.3005
R573 VTAIL.n127 VTAIL.n126 9.3005
R574 VTAIL.n129 VTAIL.n128 9.3005
R575 VTAIL.n80 VTAIL.n79 9.3005
R576 VTAIL.n135 VTAIL.n134 9.3005
R577 VTAIL.n137 VTAIL.n136 9.3005
R578 VTAIL.n76 VTAIL.n75 9.3005
R579 VTAIL.n143 VTAIL.n142 9.3005
R580 VTAIL.n193 VTAIL.n192 9.3005
R581 VTAIL.n162 VTAIL.n161 9.3005
R582 VTAIL.n187 VTAIL.n186 9.3005
R583 VTAIL.n185 VTAIL.n184 9.3005
R584 VTAIL.n166 VTAIL.n165 9.3005
R585 VTAIL.n179 VTAIL.n178 9.3005
R586 VTAIL.n177 VTAIL.n176 9.3005
R587 VTAIL.n170 VTAIL.n169 9.3005
R588 VTAIL.n195 VTAIL.n194 9.3005
R589 VTAIL.n158 VTAIL.n157 9.3005
R590 VTAIL.n201 VTAIL.n200 9.3005
R591 VTAIL.n203 VTAIL.n202 9.3005
R592 VTAIL.n154 VTAIL.n153 9.3005
R593 VTAIL.n209 VTAIL.n208 9.3005
R594 VTAIL.n211 VTAIL.n210 9.3005
R595 VTAIL.n150 VTAIL.n149 9.3005
R596 VTAIL.n217 VTAIL.n216 9.3005
R597 VTAIL.n450 VTAIL.n449 9.3005
R598 VTAIL.n493 VTAIL.n492 9.3005
R599 VTAIL.n495 VTAIL.n494 9.3005
R600 VTAIL.n446 VTAIL.n445 9.3005
R601 VTAIL.n501 VTAIL.n500 9.3005
R602 VTAIL.n503 VTAIL.n502 9.3005
R603 VTAIL.n442 VTAIL.n441 9.3005
R604 VTAIL.n509 VTAIL.n508 9.3005
R605 VTAIL.n487 VTAIL.n486 9.3005
R606 VTAIL.n485 VTAIL.n484 9.3005
R607 VTAIL.n454 VTAIL.n453 9.3005
R608 VTAIL.n479 VTAIL.n478 9.3005
R609 VTAIL.n477 VTAIL.n476 9.3005
R610 VTAIL.n458 VTAIL.n457 9.3005
R611 VTAIL.n471 VTAIL.n470 9.3005
R612 VTAIL.n469 VTAIL.n468 9.3005
R613 VTAIL.n462 VTAIL.n461 9.3005
R614 VTAIL.n376 VTAIL.n375 9.3005
R615 VTAIL.n419 VTAIL.n418 9.3005
R616 VTAIL.n421 VTAIL.n420 9.3005
R617 VTAIL.n372 VTAIL.n371 9.3005
R618 VTAIL.n427 VTAIL.n426 9.3005
R619 VTAIL.n429 VTAIL.n428 9.3005
R620 VTAIL.n368 VTAIL.n367 9.3005
R621 VTAIL.n435 VTAIL.n434 9.3005
R622 VTAIL.n413 VTAIL.n412 9.3005
R623 VTAIL.n411 VTAIL.n410 9.3005
R624 VTAIL.n380 VTAIL.n379 9.3005
R625 VTAIL.n405 VTAIL.n404 9.3005
R626 VTAIL.n403 VTAIL.n402 9.3005
R627 VTAIL.n384 VTAIL.n383 9.3005
R628 VTAIL.n397 VTAIL.n396 9.3005
R629 VTAIL.n395 VTAIL.n394 9.3005
R630 VTAIL.n388 VTAIL.n387 9.3005
R631 VTAIL.n304 VTAIL.n303 9.3005
R632 VTAIL.n347 VTAIL.n346 9.3005
R633 VTAIL.n349 VTAIL.n348 9.3005
R634 VTAIL.n300 VTAIL.n299 9.3005
R635 VTAIL.n355 VTAIL.n354 9.3005
R636 VTAIL.n357 VTAIL.n356 9.3005
R637 VTAIL.n296 VTAIL.n295 9.3005
R638 VTAIL.n363 VTAIL.n362 9.3005
R639 VTAIL.n341 VTAIL.n340 9.3005
R640 VTAIL.n339 VTAIL.n338 9.3005
R641 VTAIL.n308 VTAIL.n307 9.3005
R642 VTAIL.n333 VTAIL.n332 9.3005
R643 VTAIL.n331 VTAIL.n330 9.3005
R644 VTAIL.n312 VTAIL.n311 9.3005
R645 VTAIL.n325 VTAIL.n324 9.3005
R646 VTAIL.n323 VTAIL.n322 9.3005
R647 VTAIL.n316 VTAIL.n315 9.3005
R648 VTAIL.n230 VTAIL.n229 9.3005
R649 VTAIL.n273 VTAIL.n272 9.3005
R650 VTAIL.n275 VTAIL.n274 9.3005
R651 VTAIL.n226 VTAIL.n225 9.3005
R652 VTAIL.n281 VTAIL.n280 9.3005
R653 VTAIL.n283 VTAIL.n282 9.3005
R654 VTAIL.n222 VTAIL.n221 9.3005
R655 VTAIL.n289 VTAIL.n288 9.3005
R656 VTAIL.n267 VTAIL.n266 9.3005
R657 VTAIL.n265 VTAIL.n264 9.3005
R658 VTAIL.n234 VTAIL.n233 9.3005
R659 VTAIL.n259 VTAIL.n258 9.3005
R660 VTAIL.n257 VTAIL.n256 9.3005
R661 VTAIL.n238 VTAIL.n237 9.3005
R662 VTAIL.n251 VTAIL.n250 9.3005
R663 VTAIL.n249 VTAIL.n248 9.3005
R664 VTAIL.n242 VTAIL.n241 9.3005
R665 VTAIL.n552 VTAIL.n551 8.92171
R666 VTAIL.n567 VTAIL.n520 8.92171
R667 VTAIL.n42 VTAIL.n41 8.92171
R668 VTAIL.n57 VTAIL.n10 8.92171
R669 VTAIL.n114 VTAIL.n113 8.92171
R670 VTAIL.n129 VTAIL.n82 8.92171
R671 VTAIL.n188 VTAIL.n187 8.92171
R672 VTAIL.n203 VTAIL.n156 8.92171
R673 VTAIL.n495 VTAIL.n448 8.92171
R674 VTAIL.n480 VTAIL.n479 8.92171
R675 VTAIL.n421 VTAIL.n374 8.92171
R676 VTAIL.n406 VTAIL.n405 8.92171
R677 VTAIL.n349 VTAIL.n302 8.92171
R678 VTAIL.n334 VTAIL.n333 8.92171
R679 VTAIL.n275 VTAIL.n228 8.92171
R680 VTAIL.n260 VTAIL.n259 8.92171
R681 VTAIL.n582 VTAIL.n512 8.2187
R682 VTAIL.n72 VTAIL.n2 8.2187
R683 VTAIL.n144 VTAIL.n74 8.2187
R684 VTAIL.n218 VTAIL.n148 8.2187
R685 VTAIL.n510 VTAIL.n440 8.2187
R686 VTAIL.n436 VTAIL.n366 8.2187
R687 VTAIL.n364 VTAIL.n294 8.2187
R688 VTAIL.n290 VTAIL.n220 8.2187
R689 VTAIL.n555 VTAIL.n526 8.14595
R690 VTAIL.n564 VTAIL.n563 8.14595
R691 VTAIL.n45 VTAIL.n16 8.14595
R692 VTAIL.n54 VTAIL.n53 8.14595
R693 VTAIL.n117 VTAIL.n88 8.14595
R694 VTAIL.n126 VTAIL.n125 8.14595
R695 VTAIL.n191 VTAIL.n162 8.14595
R696 VTAIL.n200 VTAIL.n199 8.14595
R697 VTAIL.n492 VTAIL.n491 8.14595
R698 VTAIL.n483 VTAIL.n454 8.14595
R699 VTAIL.n418 VTAIL.n417 8.14595
R700 VTAIL.n409 VTAIL.n380 8.14595
R701 VTAIL.n346 VTAIL.n345 8.14595
R702 VTAIL.n337 VTAIL.n308 8.14595
R703 VTAIL.n272 VTAIL.n271 8.14595
R704 VTAIL.n263 VTAIL.n234 8.14595
R705 VTAIL.n556 VTAIL.n524 7.3702
R706 VTAIL.n560 VTAIL.n522 7.3702
R707 VTAIL.n46 VTAIL.n14 7.3702
R708 VTAIL.n50 VTAIL.n12 7.3702
R709 VTAIL.n118 VTAIL.n86 7.3702
R710 VTAIL.n122 VTAIL.n84 7.3702
R711 VTAIL.n192 VTAIL.n160 7.3702
R712 VTAIL.n196 VTAIL.n158 7.3702
R713 VTAIL.n488 VTAIL.n450 7.3702
R714 VTAIL.n484 VTAIL.n452 7.3702
R715 VTAIL.n414 VTAIL.n376 7.3702
R716 VTAIL.n410 VTAIL.n378 7.3702
R717 VTAIL.n342 VTAIL.n304 7.3702
R718 VTAIL.n338 VTAIL.n306 7.3702
R719 VTAIL.n268 VTAIL.n230 7.3702
R720 VTAIL.n264 VTAIL.n232 7.3702
R721 VTAIL.n559 VTAIL.n524 6.59444
R722 VTAIL.n560 VTAIL.n559 6.59444
R723 VTAIL.n49 VTAIL.n14 6.59444
R724 VTAIL.n50 VTAIL.n49 6.59444
R725 VTAIL.n121 VTAIL.n86 6.59444
R726 VTAIL.n122 VTAIL.n121 6.59444
R727 VTAIL.n195 VTAIL.n160 6.59444
R728 VTAIL.n196 VTAIL.n195 6.59444
R729 VTAIL.n488 VTAIL.n487 6.59444
R730 VTAIL.n487 VTAIL.n452 6.59444
R731 VTAIL.n414 VTAIL.n413 6.59444
R732 VTAIL.n413 VTAIL.n378 6.59444
R733 VTAIL.n342 VTAIL.n341 6.59444
R734 VTAIL.n341 VTAIL.n306 6.59444
R735 VTAIL.n268 VTAIL.n267 6.59444
R736 VTAIL.n267 VTAIL.n232 6.59444
R737 VTAIL.n556 VTAIL.n555 5.81868
R738 VTAIL.n563 VTAIL.n522 5.81868
R739 VTAIL.n46 VTAIL.n45 5.81868
R740 VTAIL.n53 VTAIL.n12 5.81868
R741 VTAIL.n118 VTAIL.n117 5.81868
R742 VTAIL.n125 VTAIL.n84 5.81868
R743 VTAIL.n192 VTAIL.n191 5.81868
R744 VTAIL.n199 VTAIL.n158 5.81868
R745 VTAIL.n491 VTAIL.n450 5.81868
R746 VTAIL.n484 VTAIL.n483 5.81868
R747 VTAIL.n417 VTAIL.n376 5.81868
R748 VTAIL.n410 VTAIL.n409 5.81868
R749 VTAIL.n345 VTAIL.n304 5.81868
R750 VTAIL.n338 VTAIL.n337 5.81868
R751 VTAIL.n271 VTAIL.n230 5.81868
R752 VTAIL.n264 VTAIL.n263 5.81868
R753 VTAIL.n580 VTAIL.n512 5.3904
R754 VTAIL.n70 VTAIL.n2 5.3904
R755 VTAIL.n142 VTAIL.n74 5.3904
R756 VTAIL.n216 VTAIL.n148 5.3904
R757 VTAIL.n508 VTAIL.n440 5.3904
R758 VTAIL.n434 VTAIL.n366 5.3904
R759 VTAIL.n362 VTAIL.n294 5.3904
R760 VTAIL.n288 VTAIL.n220 5.3904
R761 VTAIL.n552 VTAIL.n526 5.04292
R762 VTAIL.n564 VTAIL.n520 5.04292
R763 VTAIL.n42 VTAIL.n16 5.04292
R764 VTAIL.n54 VTAIL.n10 5.04292
R765 VTAIL.n114 VTAIL.n88 5.04292
R766 VTAIL.n126 VTAIL.n82 5.04292
R767 VTAIL.n188 VTAIL.n162 5.04292
R768 VTAIL.n200 VTAIL.n156 5.04292
R769 VTAIL.n492 VTAIL.n448 5.04292
R770 VTAIL.n480 VTAIL.n454 5.04292
R771 VTAIL.n418 VTAIL.n374 5.04292
R772 VTAIL.n406 VTAIL.n380 5.04292
R773 VTAIL.n346 VTAIL.n302 5.04292
R774 VTAIL.n334 VTAIL.n308 5.04292
R775 VTAIL.n272 VTAIL.n228 5.04292
R776 VTAIL.n260 VTAIL.n234 5.04292
R777 VTAIL.n535 VTAIL.n533 4.38563
R778 VTAIL.n25 VTAIL.n23 4.38563
R779 VTAIL.n97 VTAIL.n95 4.38563
R780 VTAIL.n171 VTAIL.n169 4.38563
R781 VTAIL.n463 VTAIL.n461 4.38563
R782 VTAIL.n389 VTAIL.n387 4.38563
R783 VTAIL.n317 VTAIL.n315 4.38563
R784 VTAIL.n243 VTAIL.n241 4.38563
R785 VTAIL.n551 VTAIL.n528 4.26717
R786 VTAIL.n568 VTAIL.n567 4.26717
R787 VTAIL.n41 VTAIL.n18 4.26717
R788 VTAIL.n58 VTAIL.n57 4.26717
R789 VTAIL.n113 VTAIL.n90 4.26717
R790 VTAIL.n130 VTAIL.n129 4.26717
R791 VTAIL.n187 VTAIL.n164 4.26717
R792 VTAIL.n204 VTAIL.n203 4.26717
R793 VTAIL.n496 VTAIL.n495 4.26717
R794 VTAIL.n479 VTAIL.n456 4.26717
R795 VTAIL.n422 VTAIL.n421 4.26717
R796 VTAIL.n405 VTAIL.n382 4.26717
R797 VTAIL.n350 VTAIL.n349 4.26717
R798 VTAIL.n333 VTAIL.n310 4.26717
R799 VTAIL.n276 VTAIL.n275 4.26717
R800 VTAIL.n259 VTAIL.n236 4.26717
R801 VTAIL.n548 VTAIL.n547 3.49141
R802 VTAIL.n571 VTAIL.n518 3.49141
R803 VTAIL.n38 VTAIL.n37 3.49141
R804 VTAIL.n61 VTAIL.n8 3.49141
R805 VTAIL.n110 VTAIL.n109 3.49141
R806 VTAIL.n133 VTAIL.n80 3.49141
R807 VTAIL.n184 VTAIL.n183 3.49141
R808 VTAIL.n207 VTAIL.n154 3.49141
R809 VTAIL.n499 VTAIL.n446 3.49141
R810 VTAIL.n476 VTAIL.n475 3.49141
R811 VTAIL.n425 VTAIL.n372 3.49141
R812 VTAIL.n402 VTAIL.n401 3.49141
R813 VTAIL.n353 VTAIL.n300 3.49141
R814 VTAIL.n330 VTAIL.n329 3.49141
R815 VTAIL.n279 VTAIL.n226 3.49141
R816 VTAIL.n256 VTAIL.n255 3.49141
R817 VTAIL.n544 VTAIL.n530 2.71565
R818 VTAIL.n572 VTAIL.n516 2.71565
R819 VTAIL.n34 VTAIL.n20 2.71565
R820 VTAIL.n62 VTAIL.n6 2.71565
R821 VTAIL.n106 VTAIL.n92 2.71565
R822 VTAIL.n134 VTAIL.n78 2.71565
R823 VTAIL.n180 VTAIL.n166 2.71565
R824 VTAIL.n208 VTAIL.n152 2.71565
R825 VTAIL.n500 VTAIL.n444 2.71565
R826 VTAIL.n472 VTAIL.n458 2.71565
R827 VTAIL.n426 VTAIL.n370 2.71565
R828 VTAIL.n398 VTAIL.n384 2.71565
R829 VTAIL.n354 VTAIL.n298 2.71565
R830 VTAIL.n326 VTAIL.n312 2.71565
R831 VTAIL.n280 VTAIL.n224 2.71565
R832 VTAIL.n252 VTAIL.n238 2.71565
R833 VTAIL.n293 VTAIL.n291 2.63843
R834 VTAIL.n365 VTAIL.n293 2.63843
R835 VTAIL.n439 VTAIL.n437 2.63843
R836 VTAIL.n511 VTAIL.n439 2.63843
R837 VTAIL.n219 VTAIL.n147 2.63843
R838 VTAIL.n147 VTAIL.n145 2.63843
R839 VTAIL.n73 VTAIL.n1 2.63843
R840 VTAIL VTAIL.n583 2.58024
R841 VTAIL.n543 VTAIL.n532 1.93989
R842 VTAIL.n576 VTAIL.n575 1.93989
R843 VTAIL.n33 VTAIL.n22 1.93989
R844 VTAIL.n66 VTAIL.n65 1.93989
R845 VTAIL.n105 VTAIL.n94 1.93989
R846 VTAIL.n138 VTAIL.n137 1.93989
R847 VTAIL.n179 VTAIL.n168 1.93989
R848 VTAIL.n212 VTAIL.n211 1.93989
R849 VTAIL.n504 VTAIL.n503 1.93989
R850 VTAIL.n471 VTAIL.n460 1.93989
R851 VTAIL.n430 VTAIL.n429 1.93989
R852 VTAIL.n397 VTAIL.n386 1.93989
R853 VTAIL.n358 VTAIL.n357 1.93989
R854 VTAIL.n325 VTAIL.n314 1.93989
R855 VTAIL.n284 VTAIL.n283 1.93989
R856 VTAIL.n251 VTAIL.n240 1.93989
R857 VTAIL.n0 VTAIL.t6 1.49034
R858 VTAIL.n0 VTAIL.t4 1.49034
R859 VTAIL.n146 VTAIL.t9 1.49034
R860 VTAIL.n146 VTAIL.t13 1.49034
R861 VTAIL.n438 VTAIL.t11 1.49034
R862 VTAIL.n438 VTAIL.t8 1.49034
R863 VTAIL.n292 VTAIL.t3 1.49034
R864 VTAIL.n292 VTAIL.t5 1.49034
R865 VTAIL.n540 VTAIL.n539 1.16414
R866 VTAIL.n579 VTAIL.n514 1.16414
R867 VTAIL.n30 VTAIL.n29 1.16414
R868 VTAIL.n69 VTAIL.n4 1.16414
R869 VTAIL.n102 VTAIL.n101 1.16414
R870 VTAIL.n141 VTAIL.n76 1.16414
R871 VTAIL.n176 VTAIL.n175 1.16414
R872 VTAIL.n215 VTAIL.n150 1.16414
R873 VTAIL.n507 VTAIL.n442 1.16414
R874 VTAIL.n468 VTAIL.n467 1.16414
R875 VTAIL.n433 VTAIL.n368 1.16414
R876 VTAIL.n394 VTAIL.n393 1.16414
R877 VTAIL.n361 VTAIL.n296 1.16414
R878 VTAIL.n322 VTAIL.n321 1.16414
R879 VTAIL.n287 VTAIL.n222 1.16414
R880 VTAIL.n248 VTAIL.n247 1.16414
R881 VTAIL.n437 VTAIL.n365 0.470328
R882 VTAIL.n145 VTAIL.n73 0.470328
R883 VTAIL.n536 VTAIL.n534 0.388379
R884 VTAIL.n26 VTAIL.n24 0.388379
R885 VTAIL.n98 VTAIL.n96 0.388379
R886 VTAIL.n172 VTAIL.n170 0.388379
R887 VTAIL.n464 VTAIL.n462 0.388379
R888 VTAIL.n390 VTAIL.n388 0.388379
R889 VTAIL.n318 VTAIL.n316 0.388379
R890 VTAIL.n244 VTAIL.n242 0.388379
R891 VTAIL.n541 VTAIL.n533 0.155672
R892 VTAIL.n542 VTAIL.n541 0.155672
R893 VTAIL.n542 VTAIL.n529 0.155672
R894 VTAIL.n549 VTAIL.n529 0.155672
R895 VTAIL.n550 VTAIL.n549 0.155672
R896 VTAIL.n550 VTAIL.n525 0.155672
R897 VTAIL.n557 VTAIL.n525 0.155672
R898 VTAIL.n558 VTAIL.n557 0.155672
R899 VTAIL.n558 VTAIL.n521 0.155672
R900 VTAIL.n565 VTAIL.n521 0.155672
R901 VTAIL.n566 VTAIL.n565 0.155672
R902 VTAIL.n566 VTAIL.n517 0.155672
R903 VTAIL.n573 VTAIL.n517 0.155672
R904 VTAIL.n574 VTAIL.n573 0.155672
R905 VTAIL.n574 VTAIL.n513 0.155672
R906 VTAIL.n581 VTAIL.n513 0.155672
R907 VTAIL.n31 VTAIL.n23 0.155672
R908 VTAIL.n32 VTAIL.n31 0.155672
R909 VTAIL.n32 VTAIL.n19 0.155672
R910 VTAIL.n39 VTAIL.n19 0.155672
R911 VTAIL.n40 VTAIL.n39 0.155672
R912 VTAIL.n40 VTAIL.n15 0.155672
R913 VTAIL.n47 VTAIL.n15 0.155672
R914 VTAIL.n48 VTAIL.n47 0.155672
R915 VTAIL.n48 VTAIL.n11 0.155672
R916 VTAIL.n55 VTAIL.n11 0.155672
R917 VTAIL.n56 VTAIL.n55 0.155672
R918 VTAIL.n56 VTAIL.n7 0.155672
R919 VTAIL.n63 VTAIL.n7 0.155672
R920 VTAIL.n64 VTAIL.n63 0.155672
R921 VTAIL.n64 VTAIL.n3 0.155672
R922 VTAIL.n71 VTAIL.n3 0.155672
R923 VTAIL.n103 VTAIL.n95 0.155672
R924 VTAIL.n104 VTAIL.n103 0.155672
R925 VTAIL.n104 VTAIL.n91 0.155672
R926 VTAIL.n111 VTAIL.n91 0.155672
R927 VTAIL.n112 VTAIL.n111 0.155672
R928 VTAIL.n112 VTAIL.n87 0.155672
R929 VTAIL.n119 VTAIL.n87 0.155672
R930 VTAIL.n120 VTAIL.n119 0.155672
R931 VTAIL.n120 VTAIL.n83 0.155672
R932 VTAIL.n127 VTAIL.n83 0.155672
R933 VTAIL.n128 VTAIL.n127 0.155672
R934 VTAIL.n128 VTAIL.n79 0.155672
R935 VTAIL.n135 VTAIL.n79 0.155672
R936 VTAIL.n136 VTAIL.n135 0.155672
R937 VTAIL.n136 VTAIL.n75 0.155672
R938 VTAIL.n143 VTAIL.n75 0.155672
R939 VTAIL.n177 VTAIL.n169 0.155672
R940 VTAIL.n178 VTAIL.n177 0.155672
R941 VTAIL.n178 VTAIL.n165 0.155672
R942 VTAIL.n185 VTAIL.n165 0.155672
R943 VTAIL.n186 VTAIL.n185 0.155672
R944 VTAIL.n186 VTAIL.n161 0.155672
R945 VTAIL.n193 VTAIL.n161 0.155672
R946 VTAIL.n194 VTAIL.n193 0.155672
R947 VTAIL.n194 VTAIL.n157 0.155672
R948 VTAIL.n201 VTAIL.n157 0.155672
R949 VTAIL.n202 VTAIL.n201 0.155672
R950 VTAIL.n202 VTAIL.n153 0.155672
R951 VTAIL.n209 VTAIL.n153 0.155672
R952 VTAIL.n210 VTAIL.n209 0.155672
R953 VTAIL.n210 VTAIL.n149 0.155672
R954 VTAIL.n217 VTAIL.n149 0.155672
R955 VTAIL.n509 VTAIL.n441 0.155672
R956 VTAIL.n502 VTAIL.n441 0.155672
R957 VTAIL.n502 VTAIL.n501 0.155672
R958 VTAIL.n501 VTAIL.n445 0.155672
R959 VTAIL.n494 VTAIL.n445 0.155672
R960 VTAIL.n494 VTAIL.n493 0.155672
R961 VTAIL.n493 VTAIL.n449 0.155672
R962 VTAIL.n486 VTAIL.n449 0.155672
R963 VTAIL.n486 VTAIL.n485 0.155672
R964 VTAIL.n485 VTAIL.n453 0.155672
R965 VTAIL.n478 VTAIL.n453 0.155672
R966 VTAIL.n478 VTAIL.n477 0.155672
R967 VTAIL.n477 VTAIL.n457 0.155672
R968 VTAIL.n470 VTAIL.n457 0.155672
R969 VTAIL.n470 VTAIL.n469 0.155672
R970 VTAIL.n469 VTAIL.n461 0.155672
R971 VTAIL.n435 VTAIL.n367 0.155672
R972 VTAIL.n428 VTAIL.n367 0.155672
R973 VTAIL.n428 VTAIL.n427 0.155672
R974 VTAIL.n427 VTAIL.n371 0.155672
R975 VTAIL.n420 VTAIL.n371 0.155672
R976 VTAIL.n420 VTAIL.n419 0.155672
R977 VTAIL.n419 VTAIL.n375 0.155672
R978 VTAIL.n412 VTAIL.n375 0.155672
R979 VTAIL.n412 VTAIL.n411 0.155672
R980 VTAIL.n411 VTAIL.n379 0.155672
R981 VTAIL.n404 VTAIL.n379 0.155672
R982 VTAIL.n404 VTAIL.n403 0.155672
R983 VTAIL.n403 VTAIL.n383 0.155672
R984 VTAIL.n396 VTAIL.n383 0.155672
R985 VTAIL.n396 VTAIL.n395 0.155672
R986 VTAIL.n395 VTAIL.n387 0.155672
R987 VTAIL.n363 VTAIL.n295 0.155672
R988 VTAIL.n356 VTAIL.n295 0.155672
R989 VTAIL.n356 VTAIL.n355 0.155672
R990 VTAIL.n355 VTAIL.n299 0.155672
R991 VTAIL.n348 VTAIL.n299 0.155672
R992 VTAIL.n348 VTAIL.n347 0.155672
R993 VTAIL.n347 VTAIL.n303 0.155672
R994 VTAIL.n340 VTAIL.n303 0.155672
R995 VTAIL.n340 VTAIL.n339 0.155672
R996 VTAIL.n339 VTAIL.n307 0.155672
R997 VTAIL.n332 VTAIL.n307 0.155672
R998 VTAIL.n332 VTAIL.n331 0.155672
R999 VTAIL.n331 VTAIL.n311 0.155672
R1000 VTAIL.n324 VTAIL.n311 0.155672
R1001 VTAIL.n324 VTAIL.n323 0.155672
R1002 VTAIL.n323 VTAIL.n315 0.155672
R1003 VTAIL.n289 VTAIL.n221 0.155672
R1004 VTAIL.n282 VTAIL.n221 0.155672
R1005 VTAIL.n282 VTAIL.n281 0.155672
R1006 VTAIL.n281 VTAIL.n225 0.155672
R1007 VTAIL.n274 VTAIL.n225 0.155672
R1008 VTAIL.n274 VTAIL.n273 0.155672
R1009 VTAIL.n273 VTAIL.n229 0.155672
R1010 VTAIL.n266 VTAIL.n229 0.155672
R1011 VTAIL.n266 VTAIL.n265 0.155672
R1012 VTAIL.n265 VTAIL.n233 0.155672
R1013 VTAIL.n258 VTAIL.n233 0.155672
R1014 VTAIL.n258 VTAIL.n257 0.155672
R1015 VTAIL.n257 VTAIL.n237 0.155672
R1016 VTAIL.n250 VTAIL.n237 0.155672
R1017 VTAIL.n250 VTAIL.n249 0.155672
R1018 VTAIL.n249 VTAIL.n241 0.155672
R1019 VTAIL VTAIL.n1 0.0586897
R1020 B.n937 B.n936 585
R1021 B.n350 B.n147 585
R1022 B.n349 B.n348 585
R1023 B.n347 B.n346 585
R1024 B.n345 B.n344 585
R1025 B.n343 B.n342 585
R1026 B.n341 B.n340 585
R1027 B.n339 B.n338 585
R1028 B.n337 B.n336 585
R1029 B.n335 B.n334 585
R1030 B.n333 B.n332 585
R1031 B.n331 B.n330 585
R1032 B.n329 B.n328 585
R1033 B.n327 B.n326 585
R1034 B.n325 B.n324 585
R1035 B.n323 B.n322 585
R1036 B.n321 B.n320 585
R1037 B.n319 B.n318 585
R1038 B.n317 B.n316 585
R1039 B.n315 B.n314 585
R1040 B.n313 B.n312 585
R1041 B.n311 B.n310 585
R1042 B.n309 B.n308 585
R1043 B.n307 B.n306 585
R1044 B.n305 B.n304 585
R1045 B.n303 B.n302 585
R1046 B.n301 B.n300 585
R1047 B.n299 B.n298 585
R1048 B.n297 B.n296 585
R1049 B.n295 B.n294 585
R1050 B.n293 B.n292 585
R1051 B.n291 B.n290 585
R1052 B.n289 B.n288 585
R1053 B.n287 B.n286 585
R1054 B.n285 B.n284 585
R1055 B.n283 B.n282 585
R1056 B.n281 B.n280 585
R1057 B.n279 B.n278 585
R1058 B.n277 B.n276 585
R1059 B.n275 B.n274 585
R1060 B.n273 B.n272 585
R1061 B.n271 B.n270 585
R1062 B.n269 B.n268 585
R1063 B.n267 B.n266 585
R1064 B.n265 B.n264 585
R1065 B.n262 B.n261 585
R1066 B.n260 B.n259 585
R1067 B.n258 B.n257 585
R1068 B.n256 B.n255 585
R1069 B.n254 B.n253 585
R1070 B.n252 B.n251 585
R1071 B.n250 B.n249 585
R1072 B.n248 B.n247 585
R1073 B.n246 B.n245 585
R1074 B.n244 B.n243 585
R1075 B.n241 B.n240 585
R1076 B.n239 B.n238 585
R1077 B.n237 B.n236 585
R1078 B.n235 B.n234 585
R1079 B.n233 B.n232 585
R1080 B.n231 B.n230 585
R1081 B.n229 B.n228 585
R1082 B.n227 B.n226 585
R1083 B.n225 B.n224 585
R1084 B.n223 B.n222 585
R1085 B.n221 B.n220 585
R1086 B.n219 B.n218 585
R1087 B.n217 B.n216 585
R1088 B.n215 B.n214 585
R1089 B.n213 B.n212 585
R1090 B.n211 B.n210 585
R1091 B.n209 B.n208 585
R1092 B.n207 B.n206 585
R1093 B.n205 B.n204 585
R1094 B.n203 B.n202 585
R1095 B.n201 B.n200 585
R1096 B.n199 B.n198 585
R1097 B.n197 B.n196 585
R1098 B.n195 B.n194 585
R1099 B.n193 B.n192 585
R1100 B.n191 B.n190 585
R1101 B.n189 B.n188 585
R1102 B.n187 B.n186 585
R1103 B.n185 B.n184 585
R1104 B.n183 B.n182 585
R1105 B.n181 B.n180 585
R1106 B.n179 B.n178 585
R1107 B.n177 B.n176 585
R1108 B.n175 B.n174 585
R1109 B.n173 B.n172 585
R1110 B.n171 B.n170 585
R1111 B.n169 B.n168 585
R1112 B.n167 B.n166 585
R1113 B.n165 B.n164 585
R1114 B.n163 B.n162 585
R1115 B.n161 B.n160 585
R1116 B.n159 B.n158 585
R1117 B.n157 B.n156 585
R1118 B.n155 B.n154 585
R1119 B.n153 B.n152 585
R1120 B.n935 B.n97 585
R1121 B.n940 B.n97 585
R1122 B.n934 B.n96 585
R1123 B.n941 B.n96 585
R1124 B.n933 B.n932 585
R1125 B.n932 B.n92 585
R1126 B.n931 B.n91 585
R1127 B.n947 B.n91 585
R1128 B.n930 B.n90 585
R1129 B.n948 B.n90 585
R1130 B.n929 B.n89 585
R1131 B.n949 B.n89 585
R1132 B.n928 B.n927 585
R1133 B.n927 B.n85 585
R1134 B.n926 B.n84 585
R1135 B.n955 B.n84 585
R1136 B.n925 B.n83 585
R1137 B.n956 B.n83 585
R1138 B.n924 B.n82 585
R1139 B.n957 B.n82 585
R1140 B.n923 B.n922 585
R1141 B.n922 B.n78 585
R1142 B.n921 B.n77 585
R1143 B.n963 B.n77 585
R1144 B.n920 B.n76 585
R1145 B.n964 B.n76 585
R1146 B.n919 B.n75 585
R1147 B.n965 B.n75 585
R1148 B.n918 B.n917 585
R1149 B.n917 B.n71 585
R1150 B.n916 B.n70 585
R1151 B.n971 B.n70 585
R1152 B.n915 B.n69 585
R1153 B.n972 B.n69 585
R1154 B.n914 B.n68 585
R1155 B.n973 B.n68 585
R1156 B.n913 B.n912 585
R1157 B.n912 B.n64 585
R1158 B.n911 B.n63 585
R1159 B.n979 B.n63 585
R1160 B.n910 B.n62 585
R1161 B.n980 B.n62 585
R1162 B.n909 B.n61 585
R1163 B.n981 B.n61 585
R1164 B.n908 B.n907 585
R1165 B.n907 B.n57 585
R1166 B.n906 B.n56 585
R1167 B.n987 B.n56 585
R1168 B.n905 B.n55 585
R1169 B.n988 B.n55 585
R1170 B.n904 B.n54 585
R1171 B.n989 B.n54 585
R1172 B.n903 B.n902 585
R1173 B.n902 B.n50 585
R1174 B.n901 B.n49 585
R1175 B.n995 B.n49 585
R1176 B.n900 B.n48 585
R1177 B.n996 B.n48 585
R1178 B.n899 B.n47 585
R1179 B.n997 B.n47 585
R1180 B.n898 B.n897 585
R1181 B.n897 B.n43 585
R1182 B.n896 B.n42 585
R1183 B.n1003 B.n42 585
R1184 B.n895 B.n41 585
R1185 B.n1004 B.n41 585
R1186 B.n894 B.n40 585
R1187 B.n1005 B.n40 585
R1188 B.n893 B.n892 585
R1189 B.n892 B.n36 585
R1190 B.n891 B.n35 585
R1191 B.n1011 B.n35 585
R1192 B.n890 B.n34 585
R1193 B.n1012 B.n34 585
R1194 B.n889 B.n33 585
R1195 B.n1013 B.n33 585
R1196 B.n888 B.n887 585
R1197 B.n887 B.n29 585
R1198 B.n886 B.n28 585
R1199 B.n1019 B.n28 585
R1200 B.n885 B.n27 585
R1201 B.n1020 B.n27 585
R1202 B.n884 B.n26 585
R1203 B.n1021 B.n26 585
R1204 B.n883 B.n882 585
R1205 B.n882 B.n22 585
R1206 B.n881 B.n21 585
R1207 B.n1027 B.n21 585
R1208 B.n880 B.n20 585
R1209 B.n1028 B.n20 585
R1210 B.n879 B.n19 585
R1211 B.n1029 B.n19 585
R1212 B.n878 B.n877 585
R1213 B.n877 B.n18 585
R1214 B.n876 B.n14 585
R1215 B.n1035 B.n14 585
R1216 B.n875 B.n13 585
R1217 B.n1036 B.n13 585
R1218 B.n874 B.n12 585
R1219 B.n1037 B.n12 585
R1220 B.n873 B.n872 585
R1221 B.n872 B.n8 585
R1222 B.n871 B.n7 585
R1223 B.n1043 B.n7 585
R1224 B.n870 B.n6 585
R1225 B.n1044 B.n6 585
R1226 B.n869 B.n5 585
R1227 B.n1045 B.n5 585
R1228 B.n868 B.n867 585
R1229 B.n867 B.n4 585
R1230 B.n866 B.n351 585
R1231 B.n866 B.n865 585
R1232 B.n856 B.n352 585
R1233 B.n353 B.n352 585
R1234 B.n858 B.n857 585
R1235 B.n859 B.n858 585
R1236 B.n855 B.n358 585
R1237 B.n358 B.n357 585
R1238 B.n854 B.n853 585
R1239 B.n853 B.n852 585
R1240 B.n360 B.n359 585
R1241 B.n845 B.n360 585
R1242 B.n844 B.n843 585
R1243 B.n846 B.n844 585
R1244 B.n842 B.n365 585
R1245 B.n365 B.n364 585
R1246 B.n841 B.n840 585
R1247 B.n840 B.n839 585
R1248 B.n367 B.n366 585
R1249 B.n368 B.n367 585
R1250 B.n832 B.n831 585
R1251 B.n833 B.n832 585
R1252 B.n830 B.n373 585
R1253 B.n373 B.n372 585
R1254 B.n829 B.n828 585
R1255 B.n828 B.n827 585
R1256 B.n375 B.n374 585
R1257 B.n376 B.n375 585
R1258 B.n820 B.n819 585
R1259 B.n821 B.n820 585
R1260 B.n818 B.n381 585
R1261 B.n381 B.n380 585
R1262 B.n817 B.n816 585
R1263 B.n816 B.n815 585
R1264 B.n383 B.n382 585
R1265 B.n384 B.n383 585
R1266 B.n808 B.n807 585
R1267 B.n809 B.n808 585
R1268 B.n806 B.n389 585
R1269 B.n389 B.n388 585
R1270 B.n805 B.n804 585
R1271 B.n804 B.n803 585
R1272 B.n391 B.n390 585
R1273 B.n392 B.n391 585
R1274 B.n796 B.n795 585
R1275 B.n797 B.n796 585
R1276 B.n794 B.n396 585
R1277 B.n400 B.n396 585
R1278 B.n793 B.n792 585
R1279 B.n792 B.n791 585
R1280 B.n398 B.n397 585
R1281 B.n399 B.n398 585
R1282 B.n784 B.n783 585
R1283 B.n785 B.n784 585
R1284 B.n782 B.n405 585
R1285 B.n405 B.n404 585
R1286 B.n781 B.n780 585
R1287 B.n780 B.n779 585
R1288 B.n407 B.n406 585
R1289 B.n408 B.n407 585
R1290 B.n772 B.n771 585
R1291 B.n773 B.n772 585
R1292 B.n770 B.n413 585
R1293 B.n413 B.n412 585
R1294 B.n769 B.n768 585
R1295 B.n768 B.n767 585
R1296 B.n415 B.n414 585
R1297 B.n416 B.n415 585
R1298 B.n760 B.n759 585
R1299 B.n761 B.n760 585
R1300 B.n758 B.n421 585
R1301 B.n421 B.n420 585
R1302 B.n757 B.n756 585
R1303 B.n756 B.n755 585
R1304 B.n423 B.n422 585
R1305 B.n424 B.n423 585
R1306 B.n748 B.n747 585
R1307 B.n749 B.n748 585
R1308 B.n746 B.n429 585
R1309 B.n429 B.n428 585
R1310 B.n745 B.n744 585
R1311 B.n744 B.n743 585
R1312 B.n431 B.n430 585
R1313 B.n432 B.n431 585
R1314 B.n736 B.n735 585
R1315 B.n737 B.n736 585
R1316 B.n734 B.n437 585
R1317 B.n437 B.n436 585
R1318 B.n733 B.n732 585
R1319 B.n732 B.n731 585
R1320 B.n439 B.n438 585
R1321 B.n440 B.n439 585
R1322 B.n724 B.n723 585
R1323 B.n725 B.n724 585
R1324 B.n722 B.n445 585
R1325 B.n445 B.n444 585
R1326 B.n721 B.n720 585
R1327 B.n720 B.n719 585
R1328 B.n447 B.n446 585
R1329 B.n448 B.n447 585
R1330 B.n712 B.n711 585
R1331 B.n713 B.n712 585
R1332 B.n710 B.n453 585
R1333 B.n453 B.n452 585
R1334 B.n705 B.n704 585
R1335 B.n703 B.n505 585
R1336 B.n702 B.n504 585
R1337 B.n707 B.n504 585
R1338 B.n701 B.n700 585
R1339 B.n699 B.n698 585
R1340 B.n697 B.n696 585
R1341 B.n695 B.n694 585
R1342 B.n693 B.n692 585
R1343 B.n691 B.n690 585
R1344 B.n689 B.n688 585
R1345 B.n687 B.n686 585
R1346 B.n685 B.n684 585
R1347 B.n683 B.n682 585
R1348 B.n681 B.n680 585
R1349 B.n679 B.n678 585
R1350 B.n677 B.n676 585
R1351 B.n675 B.n674 585
R1352 B.n673 B.n672 585
R1353 B.n671 B.n670 585
R1354 B.n669 B.n668 585
R1355 B.n667 B.n666 585
R1356 B.n665 B.n664 585
R1357 B.n663 B.n662 585
R1358 B.n661 B.n660 585
R1359 B.n659 B.n658 585
R1360 B.n657 B.n656 585
R1361 B.n655 B.n654 585
R1362 B.n653 B.n652 585
R1363 B.n651 B.n650 585
R1364 B.n649 B.n648 585
R1365 B.n647 B.n646 585
R1366 B.n645 B.n644 585
R1367 B.n643 B.n642 585
R1368 B.n641 B.n640 585
R1369 B.n639 B.n638 585
R1370 B.n637 B.n636 585
R1371 B.n635 B.n634 585
R1372 B.n633 B.n632 585
R1373 B.n631 B.n630 585
R1374 B.n629 B.n628 585
R1375 B.n627 B.n626 585
R1376 B.n625 B.n624 585
R1377 B.n623 B.n622 585
R1378 B.n621 B.n620 585
R1379 B.n619 B.n618 585
R1380 B.n617 B.n616 585
R1381 B.n615 B.n614 585
R1382 B.n613 B.n612 585
R1383 B.n611 B.n610 585
R1384 B.n609 B.n608 585
R1385 B.n607 B.n606 585
R1386 B.n605 B.n604 585
R1387 B.n603 B.n602 585
R1388 B.n601 B.n600 585
R1389 B.n599 B.n598 585
R1390 B.n597 B.n596 585
R1391 B.n595 B.n594 585
R1392 B.n593 B.n592 585
R1393 B.n591 B.n590 585
R1394 B.n589 B.n588 585
R1395 B.n587 B.n586 585
R1396 B.n585 B.n584 585
R1397 B.n583 B.n582 585
R1398 B.n581 B.n580 585
R1399 B.n579 B.n578 585
R1400 B.n577 B.n576 585
R1401 B.n575 B.n574 585
R1402 B.n573 B.n572 585
R1403 B.n571 B.n570 585
R1404 B.n569 B.n568 585
R1405 B.n567 B.n566 585
R1406 B.n565 B.n564 585
R1407 B.n563 B.n562 585
R1408 B.n561 B.n560 585
R1409 B.n559 B.n558 585
R1410 B.n557 B.n556 585
R1411 B.n555 B.n554 585
R1412 B.n553 B.n552 585
R1413 B.n551 B.n550 585
R1414 B.n549 B.n548 585
R1415 B.n547 B.n546 585
R1416 B.n545 B.n544 585
R1417 B.n543 B.n542 585
R1418 B.n541 B.n540 585
R1419 B.n539 B.n538 585
R1420 B.n537 B.n536 585
R1421 B.n535 B.n534 585
R1422 B.n533 B.n532 585
R1423 B.n531 B.n530 585
R1424 B.n529 B.n528 585
R1425 B.n527 B.n526 585
R1426 B.n525 B.n524 585
R1427 B.n523 B.n522 585
R1428 B.n521 B.n520 585
R1429 B.n519 B.n518 585
R1430 B.n517 B.n516 585
R1431 B.n515 B.n514 585
R1432 B.n513 B.n512 585
R1433 B.n455 B.n454 585
R1434 B.n709 B.n708 585
R1435 B.n708 B.n707 585
R1436 B.n451 B.n450 585
R1437 B.n452 B.n451 585
R1438 B.n715 B.n714 585
R1439 B.n714 B.n713 585
R1440 B.n716 B.n449 585
R1441 B.n449 B.n448 585
R1442 B.n718 B.n717 585
R1443 B.n719 B.n718 585
R1444 B.n443 B.n442 585
R1445 B.n444 B.n443 585
R1446 B.n727 B.n726 585
R1447 B.n726 B.n725 585
R1448 B.n728 B.n441 585
R1449 B.n441 B.n440 585
R1450 B.n730 B.n729 585
R1451 B.n731 B.n730 585
R1452 B.n435 B.n434 585
R1453 B.n436 B.n435 585
R1454 B.n739 B.n738 585
R1455 B.n738 B.n737 585
R1456 B.n740 B.n433 585
R1457 B.n433 B.n432 585
R1458 B.n742 B.n741 585
R1459 B.n743 B.n742 585
R1460 B.n427 B.n426 585
R1461 B.n428 B.n427 585
R1462 B.n751 B.n750 585
R1463 B.n750 B.n749 585
R1464 B.n752 B.n425 585
R1465 B.n425 B.n424 585
R1466 B.n754 B.n753 585
R1467 B.n755 B.n754 585
R1468 B.n419 B.n418 585
R1469 B.n420 B.n419 585
R1470 B.n763 B.n762 585
R1471 B.n762 B.n761 585
R1472 B.n764 B.n417 585
R1473 B.n417 B.n416 585
R1474 B.n766 B.n765 585
R1475 B.n767 B.n766 585
R1476 B.n411 B.n410 585
R1477 B.n412 B.n411 585
R1478 B.n775 B.n774 585
R1479 B.n774 B.n773 585
R1480 B.n776 B.n409 585
R1481 B.n409 B.n408 585
R1482 B.n778 B.n777 585
R1483 B.n779 B.n778 585
R1484 B.n403 B.n402 585
R1485 B.n404 B.n403 585
R1486 B.n787 B.n786 585
R1487 B.n786 B.n785 585
R1488 B.n788 B.n401 585
R1489 B.n401 B.n399 585
R1490 B.n790 B.n789 585
R1491 B.n791 B.n790 585
R1492 B.n395 B.n394 585
R1493 B.n400 B.n395 585
R1494 B.n799 B.n798 585
R1495 B.n798 B.n797 585
R1496 B.n800 B.n393 585
R1497 B.n393 B.n392 585
R1498 B.n802 B.n801 585
R1499 B.n803 B.n802 585
R1500 B.n387 B.n386 585
R1501 B.n388 B.n387 585
R1502 B.n811 B.n810 585
R1503 B.n810 B.n809 585
R1504 B.n812 B.n385 585
R1505 B.n385 B.n384 585
R1506 B.n814 B.n813 585
R1507 B.n815 B.n814 585
R1508 B.n379 B.n378 585
R1509 B.n380 B.n379 585
R1510 B.n823 B.n822 585
R1511 B.n822 B.n821 585
R1512 B.n824 B.n377 585
R1513 B.n377 B.n376 585
R1514 B.n826 B.n825 585
R1515 B.n827 B.n826 585
R1516 B.n371 B.n370 585
R1517 B.n372 B.n371 585
R1518 B.n835 B.n834 585
R1519 B.n834 B.n833 585
R1520 B.n836 B.n369 585
R1521 B.n369 B.n368 585
R1522 B.n838 B.n837 585
R1523 B.n839 B.n838 585
R1524 B.n363 B.n362 585
R1525 B.n364 B.n363 585
R1526 B.n848 B.n847 585
R1527 B.n847 B.n846 585
R1528 B.n849 B.n361 585
R1529 B.n845 B.n361 585
R1530 B.n851 B.n850 585
R1531 B.n852 B.n851 585
R1532 B.n356 B.n355 585
R1533 B.n357 B.n356 585
R1534 B.n861 B.n860 585
R1535 B.n860 B.n859 585
R1536 B.n862 B.n354 585
R1537 B.n354 B.n353 585
R1538 B.n864 B.n863 585
R1539 B.n865 B.n864 585
R1540 B.n2 B.n0 585
R1541 B.n4 B.n2 585
R1542 B.n3 B.n1 585
R1543 B.n1044 B.n3 585
R1544 B.n1042 B.n1041 585
R1545 B.n1043 B.n1042 585
R1546 B.n1040 B.n9 585
R1547 B.n9 B.n8 585
R1548 B.n1039 B.n1038 585
R1549 B.n1038 B.n1037 585
R1550 B.n11 B.n10 585
R1551 B.n1036 B.n11 585
R1552 B.n1034 B.n1033 585
R1553 B.n1035 B.n1034 585
R1554 B.n1032 B.n15 585
R1555 B.n18 B.n15 585
R1556 B.n1031 B.n1030 585
R1557 B.n1030 B.n1029 585
R1558 B.n17 B.n16 585
R1559 B.n1028 B.n17 585
R1560 B.n1026 B.n1025 585
R1561 B.n1027 B.n1026 585
R1562 B.n1024 B.n23 585
R1563 B.n23 B.n22 585
R1564 B.n1023 B.n1022 585
R1565 B.n1022 B.n1021 585
R1566 B.n25 B.n24 585
R1567 B.n1020 B.n25 585
R1568 B.n1018 B.n1017 585
R1569 B.n1019 B.n1018 585
R1570 B.n1016 B.n30 585
R1571 B.n30 B.n29 585
R1572 B.n1015 B.n1014 585
R1573 B.n1014 B.n1013 585
R1574 B.n32 B.n31 585
R1575 B.n1012 B.n32 585
R1576 B.n1010 B.n1009 585
R1577 B.n1011 B.n1010 585
R1578 B.n1008 B.n37 585
R1579 B.n37 B.n36 585
R1580 B.n1007 B.n1006 585
R1581 B.n1006 B.n1005 585
R1582 B.n39 B.n38 585
R1583 B.n1004 B.n39 585
R1584 B.n1002 B.n1001 585
R1585 B.n1003 B.n1002 585
R1586 B.n1000 B.n44 585
R1587 B.n44 B.n43 585
R1588 B.n999 B.n998 585
R1589 B.n998 B.n997 585
R1590 B.n46 B.n45 585
R1591 B.n996 B.n46 585
R1592 B.n994 B.n993 585
R1593 B.n995 B.n994 585
R1594 B.n992 B.n51 585
R1595 B.n51 B.n50 585
R1596 B.n991 B.n990 585
R1597 B.n990 B.n989 585
R1598 B.n53 B.n52 585
R1599 B.n988 B.n53 585
R1600 B.n986 B.n985 585
R1601 B.n987 B.n986 585
R1602 B.n984 B.n58 585
R1603 B.n58 B.n57 585
R1604 B.n983 B.n982 585
R1605 B.n982 B.n981 585
R1606 B.n60 B.n59 585
R1607 B.n980 B.n60 585
R1608 B.n978 B.n977 585
R1609 B.n979 B.n978 585
R1610 B.n976 B.n65 585
R1611 B.n65 B.n64 585
R1612 B.n975 B.n974 585
R1613 B.n974 B.n973 585
R1614 B.n67 B.n66 585
R1615 B.n972 B.n67 585
R1616 B.n970 B.n969 585
R1617 B.n971 B.n970 585
R1618 B.n968 B.n72 585
R1619 B.n72 B.n71 585
R1620 B.n967 B.n966 585
R1621 B.n966 B.n965 585
R1622 B.n74 B.n73 585
R1623 B.n964 B.n74 585
R1624 B.n962 B.n961 585
R1625 B.n963 B.n962 585
R1626 B.n960 B.n79 585
R1627 B.n79 B.n78 585
R1628 B.n959 B.n958 585
R1629 B.n958 B.n957 585
R1630 B.n81 B.n80 585
R1631 B.n956 B.n81 585
R1632 B.n954 B.n953 585
R1633 B.n955 B.n954 585
R1634 B.n952 B.n86 585
R1635 B.n86 B.n85 585
R1636 B.n951 B.n950 585
R1637 B.n950 B.n949 585
R1638 B.n88 B.n87 585
R1639 B.n948 B.n88 585
R1640 B.n946 B.n945 585
R1641 B.n947 B.n946 585
R1642 B.n944 B.n93 585
R1643 B.n93 B.n92 585
R1644 B.n943 B.n942 585
R1645 B.n942 B.n941 585
R1646 B.n95 B.n94 585
R1647 B.n940 B.n95 585
R1648 B.n1047 B.n1046 585
R1649 B.n1046 B.n1045 585
R1650 B.n705 B.n451 550.159
R1651 B.n152 B.n95 550.159
R1652 B.n708 B.n453 550.159
R1653 B.n937 B.n97 550.159
R1654 B.n509 B.t11 363.421
R1655 B.n148 B.t14 363.421
R1656 B.n506 B.t18 363.421
R1657 B.n150 B.t20 363.421
R1658 B.n509 B.t8 325.558
R1659 B.n506 B.t16 325.558
R1660 B.n150 B.t19 325.558
R1661 B.n148 B.t12 325.558
R1662 B.n510 B.t10 304.075
R1663 B.n149 B.t15 304.075
R1664 B.n507 B.t17 304.075
R1665 B.n151 B.t21 304.075
R1666 B.n939 B.n938 256.663
R1667 B.n939 B.n146 256.663
R1668 B.n939 B.n145 256.663
R1669 B.n939 B.n144 256.663
R1670 B.n939 B.n143 256.663
R1671 B.n939 B.n142 256.663
R1672 B.n939 B.n141 256.663
R1673 B.n939 B.n140 256.663
R1674 B.n939 B.n139 256.663
R1675 B.n939 B.n138 256.663
R1676 B.n939 B.n137 256.663
R1677 B.n939 B.n136 256.663
R1678 B.n939 B.n135 256.663
R1679 B.n939 B.n134 256.663
R1680 B.n939 B.n133 256.663
R1681 B.n939 B.n132 256.663
R1682 B.n939 B.n131 256.663
R1683 B.n939 B.n130 256.663
R1684 B.n939 B.n129 256.663
R1685 B.n939 B.n128 256.663
R1686 B.n939 B.n127 256.663
R1687 B.n939 B.n126 256.663
R1688 B.n939 B.n125 256.663
R1689 B.n939 B.n124 256.663
R1690 B.n939 B.n123 256.663
R1691 B.n939 B.n122 256.663
R1692 B.n939 B.n121 256.663
R1693 B.n939 B.n120 256.663
R1694 B.n939 B.n119 256.663
R1695 B.n939 B.n118 256.663
R1696 B.n939 B.n117 256.663
R1697 B.n939 B.n116 256.663
R1698 B.n939 B.n115 256.663
R1699 B.n939 B.n114 256.663
R1700 B.n939 B.n113 256.663
R1701 B.n939 B.n112 256.663
R1702 B.n939 B.n111 256.663
R1703 B.n939 B.n110 256.663
R1704 B.n939 B.n109 256.663
R1705 B.n939 B.n108 256.663
R1706 B.n939 B.n107 256.663
R1707 B.n939 B.n106 256.663
R1708 B.n939 B.n105 256.663
R1709 B.n939 B.n104 256.663
R1710 B.n939 B.n103 256.663
R1711 B.n939 B.n102 256.663
R1712 B.n939 B.n101 256.663
R1713 B.n939 B.n100 256.663
R1714 B.n939 B.n99 256.663
R1715 B.n939 B.n98 256.663
R1716 B.n707 B.n706 256.663
R1717 B.n707 B.n456 256.663
R1718 B.n707 B.n457 256.663
R1719 B.n707 B.n458 256.663
R1720 B.n707 B.n459 256.663
R1721 B.n707 B.n460 256.663
R1722 B.n707 B.n461 256.663
R1723 B.n707 B.n462 256.663
R1724 B.n707 B.n463 256.663
R1725 B.n707 B.n464 256.663
R1726 B.n707 B.n465 256.663
R1727 B.n707 B.n466 256.663
R1728 B.n707 B.n467 256.663
R1729 B.n707 B.n468 256.663
R1730 B.n707 B.n469 256.663
R1731 B.n707 B.n470 256.663
R1732 B.n707 B.n471 256.663
R1733 B.n707 B.n472 256.663
R1734 B.n707 B.n473 256.663
R1735 B.n707 B.n474 256.663
R1736 B.n707 B.n475 256.663
R1737 B.n707 B.n476 256.663
R1738 B.n707 B.n477 256.663
R1739 B.n707 B.n478 256.663
R1740 B.n707 B.n479 256.663
R1741 B.n707 B.n480 256.663
R1742 B.n707 B.n481 256.663
R1743 B.n707 B.n482 256.663
R1744 B.n707 B.n483 256.663
R1745 B.n707 B.n484 256.663
R1746 B.n707 B.n485 256.663
R1747 B.n707 B.n486 256.663
R1748 B.n707 B.n487 256.663
R1749 B.n707 B.n488 256.663
R1750 B.n707 B.n489 256.663
R1751 B.n707 B.n490 256.663
R1752 B.n707 B.n491 256.663
R1753 B.n707 B.n492 256.663
R1754 B.n707 B.n493 256.663
R1755 B.n707 B.n494 256.663
R1756 B.n707 B.n495 256.663
R1757 B.n707 B.n496 256.663
R1758 B.n707 B.n497 256.663
R1759 B.n707 B.n498 256.663
R1760 B.n707 B.n499 256.663
R1761 B.n707 B.n500 256.663
R1762 B.n707 B.n501 256.663
R1763 B.n707 B.n502 256.663
R1764 B.n707 B.n503 256.663
R1765 B.n714 B.n451 163.367
R1766 B.n714 B.n449 163.367
R1767 B.n718 B.n449 163.367
R1768 B.n718 B.n443 163.367
R1769 B.n726 B.n443 163.367
R1770 B.n726 B.n441 163.367
R1771 B.n730 B.n441 163.367
R1772 B.n730 B.n435 163.367
R1773 B.n738 B.n435 163.367
R1774 B.n738 B.n433 163.367
R1775 B.n742 B.n433 163.367
R1776 B.n742 B.n427 163.367
R1777 B.n750 B.n427 163.367
R1778 B.n750 B.n425 163.367
R1779 B.n754 B.n425 163.367
R1780 B.n754 B.n419 163.367
R1781 B.n762 B.n419 163.367
R1782 B.n762 B.n417 163.367
R1783 B.n766 B.n417 163.367
R1784 B.n766 B.n411 163.367
R1785 B.n774 B.n411 163.367
R1786 B.n774 B.n409 163.367
R1787 B.n778 B.n409 163.367
R1788 B.n778 B.n403 163.367
R1789 B.n786 B.n403 163.367
R1790 B.n786 B.n401 163.367
R1791 B.n790 B.n401 163.367
R1792 B.n790 B.n395 163.367
R1793 B.n798 B.n395 163.367
R1794 B.n798 B.n393 163.367
R1795 B.n802 B.n393 163.367
R1796 B.n802 B.n387 163.367
R1797 B.n810 B.n387 163.367
R1798 B.n810 B.n385 163.367
R1799 B.n814 B.n385 163.367
R1800 B.n814 B.n379 163.367
R1801 B.n822 B.n379 163.367
R1802 B.n822 B.n377 163.367
R1803 B.n826 B.n377 163.367
R1804 B.n826 B.n371 163.367
R1805 B.n834 B.n371 163.367
R1806 B.n834 B.n369 163.367
R1807 B.n838 B.n369 163.367
R1808 B.n838 B.n363 163.367
R1809 B.n847 B.n363 163.367
R1810 B.n847 B.n361 163.367
R1811 B.n851 B.n361 163.367
R1812 B.n851 B.n356 163.367
R1813 B.n860 B.n356 163.367
R1814 B.n860 B.n354 163.367
R1815 B.n864 B.n354 163.367
R1816 B.n864 B.n2 163.367
R1817 B.n1046 B.n2 163.367
R1818 B.n1046 B.n3 163.367
R1819 B.n1042 B.n3 163.367
R1820 B.n1042 B.n9 163.367
R1821 B.n1038 B.n9 163.367
R1822 B.n1038 B.n11 163.367
R1823 B.n1034 B.n11 163.367
R1824 B.n1034 B.n15 163.367
R1825 B.n1030 B.n15 163.367
R1826 B.n1030 B.n17 163.367
R1827 B.n1026 B.n17 163.367
R1828 B.n1026 B.n23 163.367
R1829 B.n1022 B.n23 163.367
R1830 B.n1022 B.n25 163.367
R1831 B.n1018 B.n25 163.367
R1832 B.n1018 B.n30 163.367
R1833 B.n1014 B.n30 163.367
R1834 B.n1014 B.n32 163.367
R1835 B.n1010 B.n32 163.367
R1836 B.n1010 B.n37 163.367
R1837 B.n1006 B.n37 163.367
R1838 B.n1006 B.n39 163.367
R1839 B.n1002 B.n39 163.367
R1840 B.n1002 B.n44 163.367
R1841 B.n998 B.n44 163.367
R1842 B.n998 B.n46 163.367
R1843 B.n994 B.n46 163.367
R1844 B.n994 B.n51 163.367
R1845 B.n990 B.n51 163.367
R1846 B.n990 B.n53 163.367
R1847 B.n986 B.n53 163.367
R1848 B.n986 B.n58 163.367
R1849 B.n982 B.n58 163.367
R1850 B.n982 B.n60 163.367
R1851 B.n978 B.n60 163.367
R1852 B.n978 B.n65 163.367
R1853 B.n974 B.n65 163.367
R1854 B.n974 B.n67 163.367
R1855 B.n970 B.n67 163.367
R1856 B.n970 B.n72 163.367
R1857 B.n966 B.n72 163.367
R1858 B.n966 B.n74 163.367
R1859 B.n962 B.n74 163.367
R1860 B.n962 B.n79 163.367
R1861 B.n958 B.n79 163.367
R1862 B.n958 B.n81 163.367
R1863 B.n954 B.n81 163.367
R1864 B.n954 B.n86 163.367
R1865 B.n950 B.n86 163.367
R1866 B.n950 B.n88 163.367
R1867 B.n946 B.n88 163.367
R1868 B.n946 B.n93 163.367
R1869 B.n942 B.n93 163.367
R1870 B.n942 B.n95 163.367
R1871 B.n505 B.n504 163.367
R1872 B.n700 B.n504 163.367
R1873 B.n698 B.n697 163.367
R1874 B.n694 B.n693 163.367
R1875 B.n690 B.n689 163.367
R1876 B.n686 B.n685 163.367
R1877 B.n682 B.n681 163.367
R1878 B.n678 B.n677 163.367
R1879 B.n674 B.n673 163.367
R1880 B.n670 B.n669 163.367
R1881 B.n666 B.n665 163.367
R1882 B.n662 B.n661 163.367
R1883 B.n658 B.n657 163.367
R1884 B.n654 B.n653 163.367
R1885 B.n650 B.n649 163.367
R1886 B.n646 B.n645 163.367
R1887 B.n642 B.n641 163.367
R1888 B.n638 B.n637 163.367
R1889 B.n634 B.n633 163.367
R1890 B.n630 B.n629 163.367
R1891 B.n626 B.n625 163.367
R1892 B.n622 B.n621 163.367
R1893 B.n618 B.n617 163.367
R1894 B.n614 B.n613 163.367
R1895 B.n610 B.n609 163.367
R1896 B.n606 B.n605 163.367
R1897 B.n602 B.n601 163.367
R1898 B.n598 B.n597 163.367
R1899 B.n594 B.n593 163.367
R1900 B.n590 B.n589 163.367
R1901 B.n586 B.n585 163.367
R1902 B.n582 B.n581 163.367
R1903 B.n578 B.n577 163.367
R1904 B.n574 B.n573 163.367
R1905 B.n570 B.n569 163.367
R1906 B.n566 B.n565 163.367
R1907 B.n562 B.n561 163.367
R1908 B.n558 B.n557 163.367
R1909 B.n554 B.n553 163.367
R1910 B.n550 B.n549 163.367
R1911 B.n546 B.n545 163.367
R1912 B.n542 B.n541 163.367
R1913 B.n538 B.n537 163.367
R1914 B.n534 B.n533 163.367
R1915 B.n530 B.n529 163.367
R1916 B.n526 B.n525 163.367
R1917 B.n522 B.n521 163.367
R1918 B.n518 B.n517 163.367
R1919 B.n514 B.n513 163.367
R1920 B.n708 B.n455 163.367
R1921 B.n712 B.n453 163.367
R1922 B.n712 B.n447 163.367
R1923 B.n720 B.n447 163.367
R1924 B.n720 B.n445 163.367
R1925 B.n724 B.n445 163.367
R1926 B.n724 B.n439 163.367
R1927 B.n732 B.n439 163.367
R1928 B.n732 B.n437 163.367
R1929 B.n736 B.n437 163.367
R1930 B.n736 B.n431 163.367
R1931 B.n744 B.n431 163.367
R1932 B.n744 B.n429 163.367
R1933 B.n748 B.n429 163.367
R1934 B.n748 B.n423 163.367
R1935 B.n756 B.n423 163.367
R1936 B.n756 B.n421 163.367
R1937 B.n760 B.n421 163.367
R1938 B.n760 B.n415 163.367
R1939 B.n768 B.n415 163.367
R1940 B.n768 B.n413 163.367
R1941 B.n772 B.n413 163.367
R1942 B.n772 B.n407 163.367
R1943 B.n780 B.n407 163.367
R1944 B.n780 B.n405 163.367
R1945 B.n784 B.n405 163.367
R1946 B.n784 B.n398 163.367
R1947 B.n792 B.n398 163.367
R1948 B.n792 B.n396 163.367
R1949 B.n796 B.n396 163.367
R1950 B.n796 B.n391 163.367
R1951 B.n804 B.n391 163.367
R1952 B.n804 B.n389 163.367
R1953 B.n808 B.n389 163.367
R1954 B.n808 B.n383 163.367
R1955 B.n816 B.n383 163.367
R1956 B.n816 B.n381 163.367
R1957 B.n820 B.n381 163.367
R1958 B.n820 B.n375 163.367
R1959 B.n828 B.n375 163.367
R1960 B.n828 B.n373 163.367
R1961 B.n832 B.n373 163.367
R1962 B.n832 B.n367 163.367
R1963 B.n840 B.n367 163.367
R1964 B.n840 B.n365 163.367
R1965 B.n844 B.n365 163.367
R1966 B.n844 B.n360 163.367
R1967 B.n853 B.n360 163.367
R1968 B.n853 B.n358 163.367
R1969 B.n858 B.n358 163.367
R1970 B.n858 B.n352 163.367
R1971 B.n866 B.n352 163.367
R1972 B.n867 B.n866 163.367
R1973 B.n867 B.n5 163.367
R1974 B.n6 B.n5 163.367
R1975 B.n7 B.n6 163.367
R1976 B.n872 B.n7 163.367
R1977 B.n872 B.n12 163.367
R1978 B.n13 B.n12 163.367
R1979 B.n14 B.n13 163.367
R1980 B.n877 B.n14 163.367
R1981 B.n877 B.n19 163.367
R1982 B.n20 B.n19 163.367
R1983 B.n21 B.n20 163.367
R1984 B.n882 B.n21 163.367
R1985 B.n882 B.n26 163.367
R1986 B.n27 B.n26 163.367
R1987 B.n28 B.n27 163.367
R1988 B.n887 B.n28 163.367
R1989 B.n887 B.n33 163.367
R1990 B.n34 B.n33 163.367
R1991 B.n35 B.n34 163.367
R1992 B.n892 B.n35 163.367
R1993 B.n892 B.n40 163.367
R1994 B.n41 B.n40 163.367
R1995 B.n42 B.n41 163.367
R1996 B.n897 B.n42 163.367
R1997 B.n897 B.n47 163.367
R1998 B.n48 B.n47 163.367
R1999 B.n49 B.n48 163.367
R2000 B.n902 B.n49 163.367
R2001 B.n902 B.n54 163.367
R2002 B.n55 B.n54 163.367
R2003 B.n56 B.n55 163.367
R2004 B.n907 B.n56 163.367
R2005 B.n907 B.n61 163.367
R2006 B.n62 B.n61 163.367
R2007 B.n63 B.n62 163.367
R2008 B.n912 B.n63 163.367
R2009 B.n912 B.n68 163.367
R2010 B.n69 B.n68 163.367
R2011 B.n70 B.n69 163.367
R2012 B.n917 B.n70 163.367
R2013 B.n917 B.n75 163.367
R2014 B.n76 B.n75 163.367
R2015 B.n77 B.n76 163.367
R2016 B.n922 B.n77 163.367
R2017 B.n922 B.n82 163.367
R2018 B.n83 B.n82 163.367
R2019 B.n84 B.n83 163.367
R2020 B.n927 B.n84 163.367
R2021 B.n927 B.n89 163.367
R2022 B.n90 B.n89 163.367
R2023 B.n91 B.n90 163.367
R2024 B.n932 B.n91 163.367
R2025 B.n932 B.n96 163.367
R2026 B.n97 B.n96 163.367
R2027 B.n156 B.n155 163.367
R2028 B.n160 B.n159 163.367
R2029 B.n164 B.n163 163.367
R2030 B.n168 B.n167 163.367
R2031 B.n172 B.n171 163.367
R2032 B.n176 B.n175 163.367
R2033 B.n180 B.n179 163.367
R2034 B.n184 B.n183 163.367
R2035 B.n188 B.n187 163.367
R2036 B.n192 B.n191 163.367
R2037 B.n196 B.n195 163.367
R2038 B.n200 B.n199 163.367
R2039 B.n204 B.n203 163.367
R2040 B.n208 B.n207 163.367
R2041 B.n212 B.n211 163.367
R2042 B.n216 B.n215 163.367
R2043 B.n220 B.n219 163.367
R2044 B.n224 B.n223 163.367
R2045 B.n228 B.n227 163.367
R2046 B.n232 B.n231 163.367
R2047 B.n236 B.n235 163.367
R2048 B.n240 B.n239 163.367
R2049 B.n245 B.n244 163.367
R2050 B.n249 B.n248 163.367
R2051 B.n253 B.n252 163.367
R2052 B.n257 B.n256 163.367
R2053 B.n261 B.n260 163.367
R2054 B.n266 B.n265 163.367
R2055 B.n270 B.n269 163.367
R2056 B.n274 B.n273 163.367
R2057 B.n278 B.n277 163.367
R2058 B.n282 B.n281 163.367
R2059 B.n286 B.n285 163.367
R2060 B.n290 B.n289 163.367
R2061 B.n294 B.n293 163.367
R2062 B.n298 B.n297 163.367
R2063 B.n302 B.n301 163.367
R2064 B.n306 B.n305 163.367
R2065 B.n310 B.n309 163.367
R2066 B.n314 B.n313 163.367
R2067 B.n318 B.n317 163.367
R2068 B.n322 B.n321 163.367
R2069 B.n326 B.n325 163.367
R2070 B.n330 B.n329 163.367
R2071 B.n334 B.n333 163.367
R2072 B.n338 B.n337 163.367
R2073 B.n342 B.n341 163.367
R2074 B.n346 B.n345 163.367
R2075 B.n348 B.n147 163.367
R2076 B.n707 B.n452 77.6197
R2077 B.n940 B.n939 77.6197
R2078 B.n706 B.n705 71.676
R2079 B.n700 B.n456 71.676
R2080 B.n697 B.n457 71.676
R2081 B.n693 B.n458 71.676
R2082 B.n689 B.n459 71.676
R2083 B.n685 B.n460 71.676
R2084 B.n681 B.n461 71.676
R2085 B.n677 B.n462 71.676
R2086 B.n673 B.n463 71.676
R2087 B.n669 B.n464 71.676
R2088 B.n665 B.n465 71.676
R2089 B.n661 B.n466 71.676
R2090 B.n657 B.n467 71.676
R2091 B.n653 B.n468 71.676
R2092 B.n649 B.n469 71.676
R2093 B.n645 B.n470 71.676
R2094 B.n641 B.n471 71.676
R2095 B.n637 B.n472 71.676
R2096 B.n633 B.n473 71.676
R2097 B.n629 B.n474 71.676
R2098 B.n625 B.n475 71.676
R2099 B.n621 B.n476 71.676
R2100 B.n617 B.n477 71.676
R2101 B.n613 B.n478 71.676
R2102 B.n609 B.n479 71.676
R2103 B.n605 B.n480 71.676
R2104 B.n601 B.n481 71.676
R2105 B.n597 B.n482 71.676
R2106 B.n593 B.n483 71.676
R2107 B.n589 B.n484 71.676
R2108 B.n585 B.n485 71.676
R2109 B.n581 B.n486 71.676
R2110 B.n577 B.n487 71.676
R2111 B.n573 B.n488 71.676
R2112 B.n569 B.n489 71.676
R2113 B.n565 B.n490 71.676
R2114 B.n561 B.n491 71.676
R2115 B.n557 B.n492 71.676
R2116 B.n553 B.n493 71.676
R2117 B.n549 B.n494 71.676
R2118 B.n545 B.n495 71.676
R2119 B.n541 B.n496 71.676
R2120 B.n537 B.n497 71.676
R2121 B.n533 B.n498 71.676
R2122 B.n529 B.n499 71.676
R2123 B.n525 B.n500 71.676
R2124 B.n521 B.n501 71.676
R2125 B.n517 B.n502 71.676
R2126 B.n513 B.n503 71.676
R2127 B.n152 B.n98 71.676
R2128 B.n156 B.n99 71.676
R2129 B.n160 B.n100 71.676
R2130 B.n164 B.n101 71.676
R2131 B.n168 B.n102 71.676
R2132 B.n172 B.n103 71.676
R2133 B.n176 B.n104 71.676
R2134 B.n180 B.n105 71.676
R2135 B.n184 B.n106 71.676
R2136 B.n188 B.n107 71.676
R2137 B.n192 B.n108 71.676
R2138 B.n196 B.n109 71.676
R2139 B.n200 B.n110 71.676
R2140 B.n204 B.n111 71.676
R2141 B.n208 B.n112 71.676
R2142 B.n212 B.n113 71.676
R2143 B.n216 B.n114 71.676
R2144 B.n220 B.n115 71.676
R2145 B.n224 B.n116 71.676
R2146 B.n228 B.n117 71.676
R2147 B.n232 B.n118 71.676
R2148 B.n236 B.n119 71.676
R2149 B.n240 B.n120 71.676
R2150 B.n245 B.n121 71.676
R2151 B.n249 B.n122 71.676
R2152 B.n253 B.n123 71.676
R2153 B.n257 B.n124 71.676
R2154 B.n261 B.n125 71.676
R2155 B.n266 B.n126 71.676
R2156 B.n270 B.n127 71.676
R2157 B.n274 B.n128 71.676
R2158 B.n278 B.n129 71.676
R2159 B.n282 B.n130 71.676
R2160 B.n286 B.n131 71.676
R2161 B.n290 B.n132 71.676
R2162 B.n294 B.n133 71.676
R2163 B.n298 B.n134 71.676
R2164 B.n302 B.n135 71.676
R2165 B.n306 B.n136 71.676
R2166 B.n310 B.n137 71.676
R2167 B.n314 B.n138 71.676
R2168 B.n318 B.n139 71.676
R2169 B.n322 B.n140 71.676
R2170 B.n326 B.n141 71.676
R2171 B.n330 B.n142 71.676
R2172 B.n334 B.n143 71.676
R2173 B.n338 B.n144 71.676
R2174 B.n342 B.n145 71.676
R2175 B.n346 B.n146 71.676
R2176 B.n938 B.n147 71.676
R2177 B.n938 B.n937 71.676
R2178 B.n348 B.n146 71.676
R2179 B.n345 B.n145 71.676
R2180 B.n341 B.n144 71.676
R2181 B.n337 B.n143 71.676
R2182 B.n333 B.n142 71.676
R2183 B.n329 B.n141 71.676
R2184 B.n325 B.n140 71.676
R2185 B.n321 B.n139 71.676
R2186 B.n317 B.n138 71.676
R2187 B.n313 B.n137 71.676
R2188 B.n309 B.n136 71.676
R2189 B.n305 B.n135 71.676
R2190 B.n301 B.n134 71.676
R2191 B.n297 B.n133 71.676
R2192 B.n293 B.n132 71.676
R2193 B.n289 B.n131 71.676
R2194 B.n285 B.n130 71.676
R2195 B.n281 B.n129 71.676
R2196 B.n277 B.n128 71.676
R2197 B.n273 B.n127 71.676
R2198 B.n269 B.n126 71.676
R2199 B.n265 B.n125 71.676
R2200 B.n260 B.n124 71.676
R2201 B.n256 B.n123 71.676
R2202 B.n252 B.n122 71.676
R2203 B.n248 B.n121 71.676
R2204 B.n244 B.n120 71.676
R2205 B.n239 B.n119 71.676
R2206 B.n235 B.n118 71.676
R2207 B.n231 B.n117 71.676
R2208 B.n227 B.n116 71.676
R2209 B.n223 B.n115 71.676
R2210 B.n219 B.n114 71.676
R2211 B.n215 B.n113 71.676
R2212 B.n211 B.n112 71.676
R2213 B.n207 B.n111 71.676
R2214 B.n203 B.n110 71.676
R2215 B.n199 B.n109 71.676
R2216 B.n195 B.n108 71.676
R2217 B.n191 B.n107 71.676
R2218 B.n187 B.n106 71.676
R2219 B.n183 B.n105 71.676
R2220 B.n179 B.n104 71.676
R2221 B.n175 B.n103 71.676
R2222 B.n171 B.n102 71.676
R2223 B.n167 B.n101 71.676
R2224 B.n163 B.n100 71.676
R2225 B.n159 B.n99 71.676
R2226 B.n155 B.n98 71.676
R2227 B.n706 B.n505 71.676
R2228 B.n698 B.n456 71.676
R2229 B.n694 B.n457 71.676
R2230 B.n690 B.n458 71.676
R2231 B.n686 B.n459 71.676
R2232 B.n682 B.n460 71.676
R2233 B.n678 B.n461 71.676
R2234 B.n674 B.n462 71.676
R2235 B.n670 B.n463 71.676
R2236 B.n666 B.n464 71.676
R2237 B.n662 B.n465 71.676
R2238 B.n658 B.n466 71.676
R2239 B.n654 B.n467 71.676
R2240 B.n650 B.n468 71.676
R2241 B.n646 B.n469 71.676
R2242 B.n642 B.n470 71.676
R2243 B.n638 B.n471 71.676
R2244 B.n634 B.n472 71.676
R2245 B.n630 B.n473 71.676
R2246 B.n626 B.n474 71.676
R2247 B.n622 B.n475 71.676
R2248 B.n618 B.n476 71.676
R2249 B.n614 B.n477 71.676
R2250 B.n610 B.n478 71.676
R2251 B.n606 B.n479 71.676
R2252 B.n602 B.n480 71.676
R2253 B.n598 B.n481 71.676
R2254 B.n594 B.n482 71.676
R2255 B.n590 B.n483 71.676
R2256 B.n586 B.n484 71.676
R2257 B.n582 B.n485 71.676
R2258 B.n578 B.n486 71.676
R2259 B.n574 B.n487 71.676
R2260 B.n570 B.n488 71.676
R2261 B.n566 B.n489 71.676
R2262 B.n562 B.n490 71.676
R2263 B.n558 B.n491 71.676
R2264 B.n554 B.n492 71.676
R2265 B.n550 B.n493 71.676
R2266 B.n546 B.n494 71.676
R2267 B.n542 B.n495 71.676
R2268 B.n538 B.n496 71.676
R2269 B.n534 B.n497 71.676
R2270 B.n530 B.n498 71.676
R2271 B.n526 B.n499 71.676
R2272 B.n522 B.n500 71.676
R2273 B.n518 B.n501 71.676
R2274 B.n514 B.n502 71.676
R2275 B.n503 B.n455 71.676
R2276 B.n511 B.n510 59.5399
R2277 B.n508 B.n507 59.5399
R2278 B.n242 B.n151 59.5399
R2279 B.n263 B.n149 59.5399
R2280 B.n510 B.n509 59.346
R2281 B.n507 B.n506 59.346
R2282 B.n151 B.n150 59.346
R2283 B.n149 B.n148 59.346
R2284 B.n713 B.n452 40.2914
R2285 B.n713 B.n448 40.2914
R2286 B.n719 B.n448 40.2914
R2287 B.n719 B.n444 40.2914
R2288 B.n725 B.n444 40.2914
R2289 B.n725 B.n440 40.2914
R2290 B.n731 B.n440 40.2914
R2291 B.n737 B.n436 40.2914
R2292 B.n737 B.n432 40.2914
R2293 B.n743 B.n432 40.2914
R2294 B.n743 B.n428 40.2914
R2295 B.n749 B.n428 40.2914
R2296 B.n749 B.n424 40.2914
R2297 B.n755 B.n424 40.2914
R2298 B.n755 B.n420 40.2914
R2299 B.n761 B.n420 40.2914
R2300 B.n761 B.n416 40.2914
R2301 B.n767 B.n416 40.2914
R2302 B.n773 B.n412 40.2914
R2303 B.n773 B.n408 40.2914
R2304 B.n779 B.n408 40.2914
R2305 B.n779 B.n404 40.2914
R2306 B.n785 B.n404 40.2914
R2307 B.n785 B.n399 40.2914
R2308 B.n791 B.n399 40.2914
R2309 B.n791 B.n400 40.2914
R2310 B.n797 B.n392 40.2914
R2311 B.n803 B.n392 40.2914
R2312 B.n803 B.n388 40.2914
R2313 B.n809 B.n388 40.2914
R2314 B.n809 B.n384 40.2914
R2315 B.n815 B.n384 40.2914
R2316 B.n815 B.n380 40.2914
R2317 B.n821 B.n380 40.2914
R2318 B.n827 B.n376 40.2914
R2319 B.n827 B.n372 40.2914
R2320 B.n833 B.n372 40.2914
R2321 B.n833 B.n368 40.2914
R2322 B.n839 B.n368 40.2914
R2323 B.n839 B.n364 40.2914
R2324 B.n846 B.n364 40.2914
R2325 B.n846 B.n845 40.2914
R2326 B.n852 B.n357 40.2914
R2327 B.n859 B.n357 40.2914
R2328 B.n859 B.n353 40.2914
R2329 B.n865 B.n353 40.2914
R2330 B.n865 B.n4 40.2914
R2331 B.n1045 B.n4 40.2914
R2332 B.n1045 B.n1044 40.2914
R2333 B.n1044 B.n1043 40.2914
R2334 B.n1043 B.n8 40.2914
R2335 B.n1037 B.n8 40.2914
R2336 B.n1037 B.n1036 40.2914
R2337 B.n1036 B.n1035 40.2914
R2338 B.n1029 B.n18 40.2914
R2339 B.n1029 B.n1028 40.2914
R2340 B.n1028 B.n1027 40.2914
R2341 B.n1027 B.n22 40.2914
R2342 B.n1021 B.n22 40.2914
R2343 B.n1021 B.n1020 40.2914
R2344 B.n1020 B.n1019 40.2914
R2345 B.n1019 B.n29 40.2914
R2346 B.n1013 B.n1012 40.2914
R2347 B.n1012 B.n1011 40.2914
R2348 B.n1011 B.n36 40.2914
R2349 B.n1005 B.n36 40.2914
R2350 B.n1005 B.n1004 40.2914
R2351 B.n1004 B.n1003 40.2914
R2352 B.n1003 B.n43 40.2914
R2353 B.n997 B.n43 40.2914
R2354 B.n996 B.n995 40.2914
R2355 B.n995 B.n50 40.2914
R2356 B.n989 B.n50 40.2914
R2357 B.n989 B.n988 40.2914
R2358 B.n988 B.n987 40.2914
R2359 B.n987 B.n57 40.2914
R2360 B.n981 B.n57 40.2914
R2361 B.n981 B.n980 40.2914
R2362 B.n979 B.n64 40.2914
R2363 B.n973 B.n64 40.2914
R2364 B.n973 B.n972 40.2914
R2365 B.n972 B.n971 40.2914
R2366 B.n971 B.n71 40.2914
R2367 B.n965 B.n71 40.2914
R2368 B.n965 B.n964 40.2914
R2369 B.n964 B.n963 40.2914
R2370 B.n963 B.n78 40.2914
R2371 B.n957 B.n78 40.2914
R2372 B.n957 B.n956 40.2914
R2373 B.n955 B.n85 40.2914
R2374 B.n949 B.n85 40.2914
R2375 B.n949 B.n948 40.2914
R2376 B.n948 B.n947 40.2914
R2377 B.n947 B.n92 40.2914
R2378 B.n941 B.n92 40.2914
R2379 B.n941 B.n940 40.2914
R2380 B.n767 B.t1 36.1438
R2381 B.n400 B.t3 36.1438
R2382 B.n821 B.t5 36.1438
R2383 B.n845 B.t0 36.1438
R2384 B.n18 B.t2 36.1438
R2385 B.n1013 B.t6 36.1438
R2386 B.t4 B.n996 36.1438
R2387 B.t7 B.n979 36.1438
R2388 B.n153 B.n94 35.7468
R2389 B.n710 B.n709 35.7468
R2390 B.n704 B.n450 35.7468
R2391 B.n936 B.n935 35.7468
R2392 B.n731 B.t9 27.8486
R2393 B.t13 B.n955 27.8486
R2394 B B.n1047 18.0485
R2395 B.t9 B.n436 12.4433
R2396 B.n956 B.t13 12.4433
R2397 B.n154 B.n153 10.6151
R2398 B.n157 B.n154 10.6151
R2399 B.n158 B.n157 10.6151
R2400 B.n161 B.n158 10.6151
R2401 B.n162 B.n161 10.6151
R2402 B.n165 B.n162 10.6151
R2403 B.n166 B.n165 10.6151
R2404 B.n169 B.n166 10.6151
R2405 B.n170 B.n169 10.6151
R2406 B.n173 B.n170 10.6151
R2407 B.n174 B.n173 10.6151
R2408 B.n177 B.n174 10.6151
R2409 B.n178 B.n177 10.6151
R2410 B.n181 B.n178 10.6151
R2411 B.n182 B.n181 10.6151
R2412 B.n185 B.n182 10.6151
R2413 B.n186 B.n185 10.6151
R2414 B.n189 B.n186 10.6151
R2415 B.n190 B.n189 10.6151
R2416 B.n193 B.n190 10.6151
R2417 B.n194 B.n193 10.6151
R2418 B.n197 B.n194 10.6151
R2419 B.n198 B.n197 10.6151
R2420 B.n201 B.n198 10.6151
R2421 B.n202 B.n201 10.6151
R2422 B.n205 B.n202 10.6151
R2423 B.n206 B.n205 10.6151
R2424 B.n209 B.n206 10.6151
R2425 B.n210 B.n209 10.6151
R2426 B.n213 B.n210 10.6151
R2427 B.n214 B.n213 10.6151
R2428 B.n217 B.n214 10.6151
R2429 B.n218 B.n217 10.6151
R2430 B.n221 B.n218 10.6151
R2431 B.n222 B.n221 10.6151
R2432 B.n225 B.n222 10.6151
R2433 B.n226 B.n225 10.6151
R2434 B.n229 B.n226 10.6151
R2435 B.n230 B.n229 10.6151
R2436 B.n233 B.n230 10.6151
R2437 B.n234 B.n233 10.6151
R2438 B.n237 B.n234 10.6151
R2439 B.n238 B.n237 10.6151
R2440 B.n241 B.n238 10.6151
R2441 B.n246 B.n243 10.6151
R2442 B.n247 B.n246 10.6151
R2443 B.n250 B.n247 10.6151
R2444 B.n251 B.n250 10.6151
R2445 B.n254 B.n251 10.6151
R2446 B.n255 B.n254 10.6151
R2447 B.n258 B.n255 10.6151
R2448 B.n259 B.n258 10.6151
R2449 B.n262 B.n259 10.6151
R2450 B.n267 B.n264 10.6151
R2451 B.n268 B.n267 10.6151
R2452 B.n271 B.n268 10.6151
R2453 B.n272 B.n271 10.6151
R2454 B.n275 B.n272 10.6151
R2455 B.n276 B.n275 10.6151
R2456 B.n279 B.n276 10.6151
R2457 B.n280 B.n279 10.6151
R2458 B.n283 B.n280 10.6151
R2459 B.n284 B.n283 10.6151
R2460 B.n287 B.n284 10.6151
R2461 B.n288 B.n287 10.6151
R2462 B.n291 B.n288 10.6151
R2463 B.n292 B.n291 10.6151
R2464 B.n295 B.n292 10.6151
R2465 B.n296 B.n295 10.6151
R2466 B.n299 B.n296 10.6151
R2467 B.n300 B.n299 10.6151
R2468 B.n303 B.n300 10.6151
R2469 B.n304 B.n303 10.6151
R2470 B.n307 B.n304 10.6151
R2471 B.n308 B.n307 10.6151
R2472 B.n311 B.n308 10.6151
R2473 B.n312 B.n311 10.6151
R2474 B.n315 B.n312 10.6151
R2475 B.n316 B.n315 10.6151
R2476 B.n319 B.n316 10.6151
R2477 B.n320 B.n319 10.6151
R2478 B.n323 B.n320 10.6151
R2479 B.n324 B.n323 10.6151
R2480 B.n327 B.n324 10.6151
R2481 B.n328 B.n327 10.6151
R2482 B.n331 B.n328 10.6151
R2483 B.n332 B.n331 10.6151
R2484 B.n335 B.n332 10.6151
R2485 B.n336 B.n335 10.6151
R2486 B.n339 B.n336 10.6151
R2487 B.n340 B.n339 10.6151
R2488 B.n343 B.n340 10.6151
R2489 B.n344 B.n343 10.6151
R2490 B.n347 B.n344 10.6151
R2491 B.n349 B.n347 10.6151
R2492 B.n350 B.n349 10.6151
R2493 B.n936 B.n350 10.6151
R2494 B.n711 B.n710 10.6151
R2495 B.n711 B.n446 10.6151
R2496 B.n721 B.n446 10.6151
R2497 B.n722 B.n721 10.6151
R2498 B.n723 B.n722 10.6151
R2499 B.n723 B.n438 10.6151
R2500 B.n733 B.n438 10.6151
R2501 B.n734 B.n733 10.6151
R2502 B.n735 B.n734 10.6151
R2503 B.n735 B.n430 10.6151
R2504 B.n745 B.n430 10.6151
R2505 B.n746 B.n745 10.6151
R2506 B.n747 B.n746 10.6151
R2507 B.n747 B.n422 10.6151
R2508 B.n757 B.n422 10.6151
R2509 B.n758 B.n757 10.6151
R2510 B.n759 B.n758 10.6151
R2511 B.n759 B.n414 10.6151
R2512 B.n769 B.n414 10.6151
R2513 B.n770 B.n769 10.6151
R2514 B.n771 B.n770 10.6151
R2515 B.n771 B.n406 10.6151
R2516 B.n781 B.n406 10.6151
R2517 B.n782 B.n781 10.6151
R2518 B.n783 B.n782 10.6151
R2519 B.n783 B.n397 10.6151
R2520 B.n793 B.n397 10.6151
R2521 B.n794 B.n793 10.6151
R2522 B.n795 B.n794 10.6151
R2523 B.n795 B.n390 10.6151
R2524 B.n805 B.n390 10.6151
R2525 B.n806 B.n805 10.6151
R2526 B.n807 B.n806 10.6151
R2527 B.n807 B.n382 10.6151
R2528 B.n817 B.n382 10.6151
R2529 B.n818 B.n817 10.6151
R2530 B.n819 B.n818 10.6151
R2531 B.n819 B.n374 10.6151
R2532 B.n829 B.n374 10.6151
R2533 B.n830 B.n829 10.6151
R2534 B.n831 B.n830 10.6151
R2535 B.n831 B.n366 10.6151
R2536 B.n841 B.n366 10.6151
R2537 B.n842 B.n841 10.6151
R2538 B.n843 B.n842 10.6151
R2539 B.n843 B.n359 10.6151
R2540 B.n854 B.n359 10.6151
R2541 B.n855 B.n854 10.6151
R2542 B.n857 B.n855 10.6151
R2543 B.n857 B.n856 10.6151
R2544 B.n856 B.n351 10.6151
R2545 B.n868 B.n351 10.6151
R2546 B.n869 B.n868 10.6151
R2547 B.n870 B.n869 10.6151
R2548 B.n871 B.n870 10.6151
R2549 B.n873 B.n871 10.6151
R2550 B.n874 B.n873 10.6151
R2551 B.n875 B.n874 10.6151
R2552 B.n876 B.n875 10.6151
R2553 B.n878 B.n876 10.6151
R2554 B.n879 B.n878 10.6151
R2555 B.n880 B.n879 10.6151
R2556 B.n881 B.n880 10.6151
R2557 B.n883 B.n881 10.6151
R2558 B.n884 B.n883 10.6151
R2559 B.n885 B.n884 10.6151
R2560 B.n886 B.n885 10.6151
R2561 B.n888 B.n886 10.6151
R2562 B.n889 B.n888 10.6151
R2563 B.n890 B.n889 10.6151
R2564 B.n891 B.n890 10.6151
R2565 B.n893 B.n891 10.6151
R2566 B.n894 B.n893 10.6151
R2567 B.n895 B.n894 10.6151
R2568 B.n896 B.n895 10.6151
R2569 B.n898 B.n896 10.6151
R2570 B.n899 B.n898 10.6151
R2571 B.n900 B.n899 10.6151
R2572 B.n901 B.n900 10.6151
R2573 B.n903 B.n901 10.6151
R2574 B.n904 B.n903 10.6151
R2575 B.n905 B.n904 10.6151
R2576 B.n906 B.n905 10.6151
R2577 B.n908 B.n906 10.6151
R2578 B.n909 B.n908 10.6151
R2579 B.n910 B.n909 10.6151
R2580 B.n911 B.n910 10.6151
R2581 B.n913 B.n911 10.6151
R2582 B.n914 B.n913 10.6151
R2583 B.n915 B.n914 10.6151
R2584 B.n916 B.n915 10.6151
R2585 B.n918 B.n916 10.6151
R2586 B.n919 B.n918 10.6151
R2587 B.n920 B.n919 10.6151
R2588 B.n921 B.n920 10.6151
R2589 B.n923 B.n921 10.6151
R2590 B.n924 B.n923 10.6151
R2591 B.n925 B.n924 10.6151
R2592 B.n926 B.n925 10.6151
R2593 B.n928 B.n926 10.6151
R2594 B.n929 B.n928 10.6151
R2595 B.n930 B.n929 10.6151
R2596 B.n931 B.n930 10.6151
R2597 B.n933 B.n931 10.6151
R2598 B.n934 B.n933 10.6151
R2599 B.n935 B.n934 10.6151
R2600 B.n704 B.n703 10.6151
R2601 B.n703 B.n702 10.6151
R2602 B.n702 B.n701 10.6151
R2603 B.n701 B.n699 10.6151
R2604 B.n699 B.n696 10.6151
R2605 B.n696 B.n695 10.6151
R2606 B.n695 B.n692 10.6151
R2607 B.n692 B.n691 10.6151
R2608 B.n691 B.n688 10.6151
R2609 B.n688 B.n687 10.6151
R2610 B.n687 B.n684 10.6151
R2611 B.n684 B.n683 10.6151
R2612 B.n683 B.n680 10.6151
R2613 B.n680 B.n679 10.6151
R2614 B.n679 B.n676 10.6151
R2615 B.n676 B.n675 10.6151
R2616 B.n675 B.n672 10.6151
R2617 B.n672 B.n671 10.6151
R2618 B.n671 B.n668 10.6151
R2619 B.n668 B.n667 10.6151
R2620 B.n667 B.n664 10.6151
R2621 B.n664 B.n663 10.6151
R2622 B.n663 B.n660 10.6151
R2623 B.n660 B.n659 10.6151
R2624 B.n659 B.n656 10.6151
R2625 B.n656 B.n655 10.6151
R2626 B.n655 B.n652 10.6151
R2627 B.n652 B.n651 10.6151
R2628 B.n651 B.n648 10.6151
R2629 B.n648 B.n647 10.6151
R2630 B.n647 B.n644 10.6151
R2631 B.n644 B.n643 10.6151
R2632 B.n643 B.n640 10.6151
R2633 B.n640 B.n639 10.6151
R2634 B.n639 B.n636 10.6151
R2635 B.n636 B.n635 10.6151
R2636 B.n635 B.n632 10.6151
R2637 B.n632 B.n631 10.6151
R2638 B.n631 B.n628 10.6151
R2639 B.n628 B.n627 10.6151
R2640 B.n627 B.n624 10.6151
R2641 B.n624 B.n623 10.6151
R2642 B.n623 B.n620 10.6151
R2643 B.n620 B.n619 10.6151
R2644 B.n616 B.n615 10.6151
R2645 B.n615 B.n612 10.6151
R2646 B.n612 B.n611 10.6151
R2647 B.n611 B.n608 10.6151
R2648 B.n608 B.n607 10.6151
R2649 B.n607 B.n604 10.6151
R2650 B.n604 B.n603 10.6151
R2651 B.n603 B.n600 10.6151
R2652 B.n600 B.n599 10.6151
R2653 B.n596 B.n595 10.6151
R2654 B.n595 B.n592 10.6151
R2655 B.n592 B.n591 10.6151
R2656 B.n591 B.n588 10.6151
R2657 B.n588 B.n587 10.6151
R2658 B.n587 B.n584 10.6151
R2659 B.n584 B.n583 10.6151
R2660 B.n583 B.n580 10.6151
R2661 B.n580 B.n579 10.6151
R2662 B.n579 B.n576 10.6151
R2663 B.n576 B.n575 10.6151
R2664 B.n575 B.n572 10.6151
R2665 B.n572 B.n571 10.6151
R2666 B.n571 B.n568 10.6151
R2667 B.n568 B.n567 10.6151
R2668 B.n567 B.n564 10.6151
R2669 B.n564 B.n563 10.6151
R2670 B.n563 B.n560 10.6151
R2671 B.n560 B.n559 10.6151
R2672 B.n559 B.n556 10.6151
R2673 B.n556 B.n555 10.6151
R2674 B.n555 B.n552 10.6151
R2675 B.n552 B.n551 10.6151
R2676 B.n551 B.n548 10.6151
R2677 B.n548 B.n547 10.6151
R2678 B.n547 B.n544 10.6151
R2679 B.n544 B.n543 10.6151
R2680 B.n543 B.n540 10.6151
R2681 B.n540 B.n539 10.6151
R2682 B.n539 B.n536 10.6151
R2683 B.n536 B.n535 10.6151
R2684 B.n535 B.n532 10.6151
R2685 B.n532 B.n531 10.6151
R2686 B.n531 B.n528 10.6151
R2687 B.n528 B.n527 10.6151
R2688 B.n527 B.n524 10.6151
R2689 B.n524 B.n523 10.6151
R2690 B.n523 B.n520 10.6151
R2691 B.n520 B.n519 10.6151
R2692 B.n519 B.n516 10.6151
R2693 B.n516 B.n515 10.6151
R2694 B.n515 B.n512 10.6151
R2695 B.n512 B.n454 10.6151
R2696 B.n709 B.n454 10.6151
R2697 B.n715 B.n450 10.6151
R2698 B.n716 B.n715 10.6151
R2699 B.n717 B.n716 10.6151
R2700 B.n717 B.n442 10.6151
R2701 B.n727 B.n442 10.6151
R2702 B.n728 B.n727 10.6151
R2703 B.n729 B.n728 10.6151
R2704 B.n729 B.n434 10.6151
R2705 B.n739 B.n434 10.6151
R2706 B.n740 B.n739 10.6151
R2707 B.n741 B.n740 10.6151
R2708 B.n741 B.n426 10.6151
R2709 B.n751 B.n426 10.6151
R2710 B.n752 B.n751 10.6151
R2711 B.n753 B.n752 10.6151
R2712 B.n753 B.n418 10.6151
R2713 B.n763 B.n418 10.6151
R2714 B.n764 B.n763 10.6151
R2715 B.n765 B.n764 10.6151
R2716 B.n765 B.n410 10.6151
R2717 B.n775 B.n410 10.6151
R2718 B.n776 B.n775 10.6151
R2719 B.n777 B.n776 10.6151
R2720 B.n777 B.n402 10.6151
R2721 B.n787 B.n402 10.6151
R2722 B.n788 B.n787 10.6151
R2723 B.n789 B.n788 10.6151
R2724 B.n789 B.n394 10.6151
R2725 B.n799 B.n394 10.6151
R2726 B.n800 B.n799 10.6151
R2727 B.n801 B.n800 10.6151
R2728 B.n801 B.n386 10.6151
R2729 B.n811 B.n386 10.6151
R2730 B.n812 B.n811 10.6151
R2731 B.n813 B.n812 10.6151
R2732 B.n813 B.n378 10.6151
R2733 B.n823 B.n378 10.6151
R2734 B.n824 B.n823 10.6151
R2735 B.n825 B.n824 10.6151
R2736 B.n825 B.n370 10.6151
R2737 B.n835 B.n370 10.6151
R2738 B.n836 B.n835 10.6151
R2739 B.n837 B.n836 10.6151
R2740 B.n837 B.n362 10.6151
R2741 B.n848 B.n362 10.6151
R2742 B.n849 B.n848 10.6151
R2743 B.n850 B.n849 10.6151
R2744 B.n850 B.n355 10.6151
R2745 B.n861 B.n355 10.6151
R2746 B.n862 B.n861 10.6151
R2747 B.n863 B.n862 10.6151
R2748 B.n863 B.n0 10.6151
R2749 B.n1041 B.n1 10.6151
R2750 B.n1041 B.n1040 10.6151
R2751 B.n1040 B.n1039 10.6151
R2752 B.n1039 B.n10 10.6151
R2753 B.n1033 B.n10 10.6151
R2754 B.n1033 B.n1032 10.6151
R2755 B.n1032 B.n1031 10.6151
R2756 B.n1031 B.n16 10.6151
R2757 B.n1025 B.n16 10.6151
R2758 B.n1025 B.n1024 10.6151
R2759 B.n1024 B.n1023 10.6151
R2760 B.n1023 B.n24 10.6151
R2761 B.n1017 B.n24 10.6151
R2762 B.n1017 B.n1016 10.6151
R2763 B.n1016 B.n1015 10.6151
R2764 B.n1015 B.n31 10.6151
R2765 B.n1009 B.n31 10.6151
R2766 B.n1009 B.n1008 10.6151
R2767 B.n1008 B.n1007 10.6151
R2768 B.n1007 B.n38 10.6151
R2769 B.n1001 B.n38 10.6151
R2770 B.n1001 B.n1000 10.6151
R2771 B.n1000 B.n999 10.6151
R2772 B.n999 B.n45 10.6151
R2773 B.n993 B.n45 10.6151
R2774 B.n993 B.n992 10.6151
R2775 B.n992 B.n991 10.6151
R2776 B.n991 B.n52 10.6151
R2777 B.n985 B.n52 10.6151
R2778 B.n985 B.n984 10.6151
R2779 B.n984 B.n983 10.6151
R2780 B.n983 B.n59 10.6151
R2781 B.n977 B.n59 10.6151
R2782 B.n977 B.n976 10.6151
R2783 B.n976 B.n975 10.6151
R2784 B.n975 B.n66 10.6151
R2785 B.n969 B.n66 10.6151
R2786 B.n969 B.n968 10.6151
R2787 B.n968 B.n967 10.6151
R2788 B.n967 B.n73 10.6151
R2789 B.n961 B.n73 10.6151
R2790 B.n961 B.n960 10.6151
R2791 B.n960 B.n959 10.6151
R2792 B.n959 B.n80 10.6151
R2793 B.n953 B.n80 10.6151
R2794 B.n953 B.n952 10.6151
R2795 B.n952 B.n951 10.6151
R2796 B.n951 B.n87 10.6151
R2797 B.n945 B.n87 10.6151
R2798 B.n945 B.n944 10.6151
R2799 B.n944 B.n943 10.6151
R2800 B.n943 B.n94 10.6151
R2801 B.n242 B.n241 9.36635
R2802 B.n264 B.n263 9.36635
R2803 B.n619 B.n508 9.36635
R2804 B.n596 B.n511 9.36635
R2805 B.t1 B.n412 4.14809
R2806 B.n797 B.t3 4.14809
R2807 B.t5 B.n376 4.14809
R2808 B.n852 B.t0 4.14809
R2809 B.n1035 B.t2 4.14809
R2810 B.t6 B.n29 4.14809
R2811 B.n997 B.t4 4.14809
R2812 B.n980 B.t7 4.14809
R2813 B.n1047 B.n0 2.81026
R2814 B.n1047 B.n1 2.81026
R2815 B.n243 B.n242 1.24928
R2816 B.n263 B.n262 1.24928
R2817 B.n616 B.n508 1.24928
R2818 B.n599 B.n511 1.24928
R2819 VN.n59 VN.n31 161.3
R2820 VN.n58 VN.n57 161.3
R2821 VN.n56 VN.n32 161.3
R2822 VN.n55 VN.n54 161.3
R2823 VN.n53 VN.n33 161.3
R2824 VN.n52 VN.n51 161.3
R2825 VN.n50 VN.n49 161.3
R2826 VN.n48 VN.n35 161.3
R2827 VN.n47 VN.n46 161.3
R2828 VN.n45 VN.n36 161.3
R2829 VN.n44 VN.n43 161.3
R2830 VN.n42 VN.n37 161.3
R2831 VN.n41 VN.n40 161.3
R2832 VN.n28 VN.n0 161.3
R2833 VN.n27 VN.n26 161.3
R2834 VN.n25 VN.n1 161.3
R2835 VN.n24 VN.n23 161.3
R2836 VN.n22 VN.n2 161.3
R2837 VN.n21 VN.n20 161.3
R2838 VN.n19 VN.n18 161.3
R2839 VN.n17 VN.n4 161.3
R2840 VN.n16 VN.n15 161.3
R2841 VN.n14 VN.n5 161.3
R2842 VN.n13 VN.n12 161.3
R2843 VN.n11 VN.n6 161.3
R2844 VN.n10 VN.n9 161.3
R2845 VN.n8 VN.t3 148.993
R2846 VN.n39 VN.t4 148.993
R2847 VN.n7 VN.t0 117.323
R2848 VN.n3 VN.t6 117.323
R2849 VN.n29 VN.t2 117.323
R2850 VN.n38 VN.t7 117.323
R2851 VN.n34 VN.t1 117.323
R2852 VN.n60 VN.t5 117.323
R2853 VN.n30 VN.n29 106.353
R2854 VN.n61 VN.n60 106.353
R2855 VN.n8 VN.n7 71.7459
R2856 VN.n39 VN.n38 71.7459
R2857 VN VN.n61 52.7254
R2858 VN.n23 VN.n1 46.321
R2859 VN.n54 VN.n32 46.321
R2860 VN.n12 VN.n5 40.4934
R2861 VN.n16 VN.n5 40.4934
R2862 VN.n43 VN.n36 40.4934
R2863 VN.n47 VN.n36 40.4934
R2864 VN.n23 VN.n22 34.6658
R2865 VN.n54 VN.n53 34.6658
R2866 VN.n11 VN.n10 24.4675
R2867 VN.n12 VN.n11 24.4675
R2868 VN.n17 VN.n16 24.4675
R2869 VN.n18 VN.n17 24.4675
R2870 VN.n22 VN.n21 24.4675
R2871 VN.n27 VN.n1 24.4675
R2872 VN.n28 VN.n27 24.4675
R2873 VN.n43 VN.n42 24.4675
R2874 VN.n42 VN.n41 24.4675
R2875 VN.n53 VN.n52 24.4675
R2876 VN.n49 VN.n48 24.4675
R2877 VN.n48 VN.n47 24.4675
R2878 VN.n59 VN.n58 24.4675
R2879 VN.n58 VN.n32 24.4675
R2880 VN.n21 VN.n3 22.9995
R2881 VN.n52 VN.n34 22.9995
R2882 VN.n40 VN.n39 7.21203
R2883 VN.n9 VN.n8 7.21203
R2884 VN.n29 VN.n28 4.40456
R2885 VN.n60 VN.n59 4.40456
R2886 VN.n10 VN.n7 1.46852
R2887 VN.n18 VN.n3 1.46852
R2888 VN.n41 VN.n38 1.46852
R2889 VN.n49 VN.n34 1.46852
R2890 VN.n61 VN.n31 0.278367
R2891 VN.n30 VN.n0 0.278367
R2892 VN.n57 VN.n31 0.189894
R2893 VN.n57 VN.n56 0.189894
R2894 VN.n56 VN.n55 0.189894
R2895 VN.n55 VN.n33 0.189894
R2896 VN.n51 VN.n33 0.189894
R2897 VN.n51 VN.n50 0.189894
R2898 VN.n50 VN.n35 0.189894
R2899 VN.n46 VN.n35 0.189894
R2900 VN.n46 VN.n45 0.189894
R2901 VN.n45 VN.n44 0.189894
R2902 VN.n44 VN.n37 0.189894
R2903 VN.n40 VN.n37 0.189894
R2904 VN.n9 VN.n6 0.189894
R2905 VN.n13 VN.n6 0.189894
R2906 VN.n14 VN.n13 0.189894
R2907 VN.n15 VN.n14 0.189894
R2908 VN.n15 VN.n4 0.189894
R2909 VN.n19 VN.n4 0.189894
R2910 VN.n20 VN.n19 0.189894
R2911 VN.n20 VN.n2 0.189894
R2912 VN.n24 VN.n2 0.189894
R2913 VN.n25 VN.n24 0.189894
R2914 VN.n26 VN.n25 0.189894
R2915 VN.n26 VN.n0 0.189894
R2916 VN VN.n30 0.153454
R2917 VDD2.n2 VDD2.n1 64.1285
R2918 VDD2.n2 VDD2.n0 64.1285
R2919 VDD2 VDD2.n5 64.1257
R2920 VDD2.n4 VDD2.n3 62.8651
R2921 VDD2.n4 VDD2.n2 47.0429
R2922 VDD2.n5 VDD2.t0 1.49034
R2923 VDD2.n5 VDD2.t3 1.49034
R2924 VDD2.n3 VDD2.t2 1.49034
R2925 VDD2.n3 VDD2.t6 1.49034
R2926 VDD2.n1 VDD2.t1 1.49034
R2927 VDD2.n1 VDD2.t5 1.49034
R2928 VDD2.n0 VDD2.t4 1.49034
R2929 VDD2.n0 VDD2.t7 1.49034
R2930 VDD2 VDD2.n4 1.37766
C0 VDD1 VP 10.055201f
C1 VN VTAIL 10.0537f
C2 VDD2 VN 9.675079f
C3 VDD2 VTAIL 8.58524f
C4 VDD1 VN 0.151684f
C5 VDD1 VTAIL 8.52995f
C6 VP VN 8.06101f
C7 VDD1 VDD2 1.84312f
C8 VP VTAIL 10.0678f
C9 VDD2 VP 0.533225f
C10 VDD2 B 5.561494f
C11 VDD1 B 6.011205f
C12 VTAIL B 11.344266f
C13 VN B 16.110828f
C14 VP B 14.688339f
C15 VDD2.t4 B 0.255358f
C16 VDD2.t7 B 0.255358f
C17 VDD2.n0 B 2.3065f
C18 VDD2.t1 B 0.255358f
C19 VDD2.t5 B 0.255358f
C20 VDD2.n1 B 2.3065f
C21 VDD2.n2 B 3.33046f
C22 VDD2.t2 B 0.255358f
C23 VDD2.t6 B 0.255358f
C24 VDD2.n3 B 2.29644f
C25 VDD2.n4 B 3.00367f
C26 VDD2.t0 B 0.255358f
C27 VDD2.t3 B 0.255358f
C28 VDD2.n5 B 2.30646f
C29 VN.n0 B 0.028063f
C30 VN.t2 B 2.11002f
C31 VN.n1 B 0.040594f
C32 VN.n2 B 0.021286f
C33 VN.t6 B 2.11002f
C34 VN.n3 B 0.741019f
C35 VN.n4 B 0.021286f
C36 VN.n5 B 0.017208f
C37 VN.n6 B 0.021286f
C38 VN.t0 B 2.11002f
C39 VN.n7 B 0.797131f
C40 VN.t3 B 2.29603f
C41 VN.n8 B 0.782838f
C42 VN.n9 B 0.208482f
C43 VN.n10 B 0.02126f
C44 VN.n11 B 0.039671f
C45 VN.n12 B 0.042305f
C46 VN.n13 B 0.021286f
C47 VN.n14 B 0.021286f
C48 VN.n15 B 0.021286f
C49 VN.n16 B 0.042305f
C50 VN.n17 B 0.039671f
C51 VN.n18 B 0.02126f
C52 VN.n19 B 0.021286f
C53 VN.n20 B 0.021286f
C54 VN.n21 B 0.038496f
C55 VN.n22 B 0.043012f
C56 VN.n23 B 0.018213f
C57 VN.n24 B 0.021286f
C58 VN.n25 B 0.021286f
C59 VN.n26 B 0.021286f
C60 VN.n27 B 0.039671f
C61 VN.n28 B 0.023611f
C62 VN.n29 B 0.809609f
C63 VN.n30 B 0.038425f
C64 VN.n31 B 0.028063f
C65 VN.t5 B 2.11002f
C66 VN.n32 B 0.040594f
C67 VN.n33 B 0.021286f
C68 VN.t1 B 2.11002f
C69 VN.n34 B 0.741019f
C70 VN.n35 B 0.021286f
C71 VN.n36 B 0.017208f
C72 VN.n37 B 0.021286f
C73 VN.t7 B 2.11002f
C74 VN.n38 B 0.797131f
C75 VN.t4 B 2.29603f
C76 VN.n39 B 0.782838f
C77 VN.n40 B 0.208482f
C78 VN.n41 B 0.02126f
C79 VN.n42 B 0.039671f
C80 VN.n43 B 0.042305f
C81 VN.n44 B 0.021286f
C82 VN.n45 B 0.021286f
C83 VN.n46 B 0.021286f
C84 VN.n47 B 0.042305f
C85 VN.n48 B 0.039671f
C86 VN.n49 B 0.02126f
C87 VN.n50 B 0.021286f
C88 VN.n51 B 0.021286f
C89 VN.n52 B 0.038496f
C90 VN.n53 B 0.043012f
C91 VN.n54 B 0.018213f
C92 VN.n55 B 0.021286f
C93 VN.n56 B 0.021286f
C94 VN.n57 B 0.021286f
C95 VN.n58 B 0.039671f
C96 VN.n59 B 0.023611f
C97 VN.n60 B 0.809609f
C98 VN.n61 B 1.28445f
C99 VTAIL.t6 B 0.205677f
C100 VTAIL.t4 B 0.205677f
C101 VTAIL.n0 B 1.79421f
C102 VTAIL.n1 B 0.356189f
C103 VTAIL.n2 B 0.026049f
C104 VTAIL.n3 B 0.019584f
C105 VTAIL.n4 B 0.010524f
C106 VTAIL.n5 B 0.024874f
C107 VTAIL.n6 B 0.011143f
C108 VTAIL.n7 B 0.019584f
C109 VTAIL.n8 B 0.010524f
C110 VTAIL.n9 B 0.024874f
C111 VTAIL.n10 B 0.011143f
C112 VTAIL.n11 B 0.019584f
C113 VTAIL.n12 B 0.010524f
C114 VTAIL.n13 B 0.024874f
C115 VTAIL.n14 B 0.011143f
C116 VTAIL.n15 B 0.019584f
C117 VTAIL.n16 B 0.010524f
C118 VTAIL.n17 B 0.024874f
C119 VTAIL.n18 B 0.011143f
C120 VTAIL.n19 B 0.019584f
C121 VTAIL.n20 B 0.010524f
C122 VTAIL.n21 B 0.024874f
C123 VTAIL.n22 B 0.011143f
C124 VTAIL.n23 B 1.1207f
C125 VTAIL.n24 B 0.010524f
C126 VTAIL.t2 B 0.0409f
C127 VTAIL.n25 B 0.119336f
C128 VTAIL.n26 B 0.014694f
C129 VTAIL.n27 B 0.018656f
C130 VTAIL.n28 B 0.024874f
C131 VTAIL.n29 B 0.011143f
C132 VTAIL.n30 B 0.010524f
C133 VTAIL.n31 B 0.019584f
C134 VTAIL.n32 B 0.019584f
C135 VTAIL.n33 B 0.010524f
C136 VTAIL.n34 B 0.011143f
C137 VTAIL.n35 B 0.024874f
C138 VTAIL.n36 B 0.024874f
C139 VTAIL.n37 B 0.011143f
C140 VTAIL.n38 B 0.010524f
C141 VTAIL.n39 B 0.019584f
C142 VTAIL.n40 B 0.019584f
C143 VTAIL.n41 B 0.010524f
C144 VTAIL.n42 B 0.011143f
C145 VTAIL.n43 B 0.024874f
C146 VTAIL.n44 B 0.024874f
C147 VTAIL.n45 B 0.011143f
C148 VTAIL.n46 B 0.010524f
C149 VTAIL.n47 B 0.019584f
C150 VTAIL.n48 B 0.019584f
C151 VTAIL.n49 B 0.010524f
C152 VTAIL.n50 B 0.011143f
C153 VTAIL.n51 B 0.024874f
C154 VTAIL.n52 B 0.024874f
C155 VTAIL.n53 B 0.011143f
C156 VTAIL.n54 B 0.010524f
C157 VTAIL.n55 B 0.019584f
C158 VTAIL.n56 B 0.019584f
C159 VTAIL.n57 B 0.010524f
C160 VTAIL.n58 B 0.011143f
C161 VTAIL.n59 B 0.024874f
C162 VTAIL.n60 B 0.024874f
C163 VTAIL.n61 B 0.011143f
C164 VTAIL.n62 B 0.010524f
C165 VTAIL.n63 B 0.019584f
C166 VTAIL.n64 B 0.019584f
C167 VTAIL.n65 B 0.010524f
C168 VTAIL.n66 B 0.011143f
C169 VTAIL.n67 B 0.024874f
C170 VTAIL.n68 B 0.05018f
C171 VTAIL.n69 B 0.011143f
C172 VTAIL.n70 B 0.020577f
C173 VTAIL.n71 B 0.047676f
C174 VTAIL.n72 B 0.050803f
C175 VTAIL.n73 B 0.214202f
C176 VTAIL.n74 B 0.026049f
C177 VTAIL.n75 B 0.019584f
C178 VTAIL.n76 B 0.010524f
C179 VTAIL.n77 B 0.024874f
C180 VTAIL.n78 B 0.011143f
C181 VTAIL.n79 B 0.019584f
C182 VTAIL.n80 B 0.010524f
C183 VTAIL.n81 B 0.024874f
C184 VTAIL.n82 B 0.011143f
C185 VTAIL.n83 B 0.019584f
C186 VTAIL.n84 B 0.010524f
C187 VTAIL.n85 B 0.024874f
C188 VTAIL.n86 B 0.011143f
C189 VTAIL.n87 B 0.019584f
C190 VTAIL.n88 B 0.010524f
C191 VTAIL.n89 B 0.024874f
C192 VTAIL.n90 B 0.011143f
C193 VTAIL.n91 B 0.019584f
C194 VTAIL.n92 B 0.010524f
C195 VTAIL.n93 B 0.024874f
C196 VTAIL.n94 B 0.011143f
C197 VTAIL.n95 B 1.1207f
C198 VTAIL.n96 B 0.010524f
C199 VTAIL.t10 B 0.0409f
C200 VTAIL.n97 B 0.119336f
C201 VTAIL.n98 B 0.014694f
C202 VTAIL.n99 B 0.018656f
C203 VTAIL.n100 B 0.024874f
C204 VTAIL.n101 B 0.011143f
C205 VTAIL.n102 B 0.010524f
C206 VTAIL.n103 B 0.019584f
C207 VTAIL.n104 B 0.019584f
C208 VTAIL.n105 B 0.010524f
C209 VTAIL.n106 B 0.011143f
C210 VTAIL.n107 B 0.024874f
C211 VTAIL.n108 B 0.024874f
C212 VTAIL.n109 B 0.011143f
C213 VTAIL.n110 B 0.010524f
C214 VTAIL.n111 B 0.019584f
C215 VTAIL.n112 B 0.019584f
C216 VTAIL.n113 B 0.010524f
C217 VTAIL.n114 B 0.011143f
C218 VTAIL.n115 B 0.024874f
C219 VTAIL.n116 B 0.024874f
C220 VTAIL.n117 B 0.011143f
C221 VTAIL.n118 B 0.010524f
C222 VTAIL.n119 B 0.019584f
C223 VTAIL.n120 B 0.019584f
C224 VTAIL.n121 B 0.010524f
C225 VTAIL.n122 B 0.011143f
C226 VTAIL.n123 B 0.024874f
C227 VTAIL.n124 B 0.024874f
C228 VTAIL.n125 B 0.011143f
C229 VTAIL.n126 B 0.010524f
C230 VTAIL.n127 B 0.019584f
C231 VTAIL.n128 B 0.019584f
C232 VTAIL.n129 B 0.010524f
C233 VTAIL.n130 B 0.011143f
C234 VTAIL.n131 B 0.024874f
C235 VTAIL.n132 B 0.024874f
C236 VTAIL.n133 B 0.011143f
C237 VTAIL.n134 B 0.010524f
C238 VTAIL.n135 B 0.019584f
C239 VTAIL.n136 B 0.019584f
C240 VTAIL.n137 B 0.010524f
C241 VTAIL.n138 B 0.011143f
C242 VTAIL.n139 B 0.024874f
C243 VTAIL.n140 B 0.05018f
C244 VTAIL.n141 B 0.011143f
C245 VTAIL.n142 B 0.020577f
C246 VTAIL.n143 B 0.047676f
C247 VTAIL.n144 B 0.050803f
C248 VTAIL.n145 B 0.214202f
C249 VTAIL.t9 B 0.205677f
C250 VTAIL.t13 B 0.205677f
C251 VTAIL.n146 B 1.79421f
C252 VTAIL.n147 B 0.518983f
C253 VTAIL.n148 B 0.026049f
C254 VTAIL.n149 B 0.019584f
C255 VTAIL.n150 B 0.010524f
C256 VTAIL.n151 B 0.024874f
C257 VTAIL.n152 B 0.011143f
C258 VTAIL.n153 B 0.019584f
C259 VTAIL.n154 B 0.010524f
C260 VTAIL.n155 B 0.024874f
C261 VTAIL.n156 B 0.011143f
C262 VTAIL.n157 B 0.019584f
C263 VTAIL.n158 B 0.010524f
C264 VTAIL.n159 B 0.024874f
C265 VTAIL.n160 B 0.011143f
C266 VTAIL.n161 B 0.019584f
C267 VTAIL.n162 B 0.010524f
C268 VTAIL.n163 B 0.024874f
C269 VTAIL.n164 B 0.011143f
C270 VTAIL.n165 B 0.019584f
C271 VTAIL.n166 B 0.010524f
C272 VTAIL.n167 B 0.024874f
C273 VTAIL.n168 B 0.011143f
C274 VTAIL.n169 B 1.1207f
C275 VTAIL.n170 B 0.010524f
C276 VTAIL.t12 B 0.0409f
C277 VTAIL.n171 B 0.119336f
C278 VTAIL.n172 B 0.014694f
C279 VTAIL.n173 B 0.018656f
C280 VTAIL.n174 B 0.024874f
C281 VTAIL.n175 B 0.011143f
C282 VTAIL.n176 B 0.010524f
C283 VTAIL.n177 B 0.019584f
C284 VTAIL.n178 B 0.019584f
C285 VTAIL.n179 B 0.010524f
C286 VTAIL.n180 B 0.011143f
C287 VTAIL.n181 B 0.024874f
C288 VTAIL.n182 B 0.024874f
C289 VTAIL.n183 B 0.011143f
C290 VTAIL.n184 B 0.010524f
C291 VTAIL.n185 B 0.019584f
C292 VTAIL.n186 B 0.019584f
C293 VTAIL.n187 B 0.010524f
C294 VTAIL.n188 B 0.011143f
C295 VTAIL.n189 B 0.024874f
C296 VTAIL.n190 B 0.024874f
C297 VTAIL.n191 B 0.011143f
C298 VTAIL.n192 B 0.010524f
C299 VTAIL.n193 B 0.019584f
C300 VTAIL.n194 B 0.019584f
C301 VTAIL.n195 B 0.010524f
C302 VTAIL.n196 B 0.011143f
C303 VTAIL.n197 B 0.024874f
C304 VTAIL.n198 B 0.024874f
C305 VTAIL.n199 B 0.011143f
C306 VTAIL.n200 B 0.010524f
C307 VTAIL.n201 B 0.019584f
C308 VTAIL.n202 B 0.019584f
C309 VTAIL.n203 B 0.010524f
C310 VTAIL.n204 B 0.011143f
C311 VTAIL.n205 B 0.024874f
C312 VTAIL.n206 B 0.024874f
C313 VTAIL.n207 B 0.011143f
C314 VTAIL.n208 B 0.010524f
C315 VTAIL.n209 B 0.019584f
C316 VTAIL.n210 B 0.019584f
C317 VTAIL.n211 B 0.010524f
C318 VTAIL.n212 B 0.011143f
C319 VTAIL.n213 B 0.024874f
C320 VTAIL.n214 B 0.05018f
C321 VTAIL.n215 B 0.011143f
C322 VTAIL.n216 B 0.020577f
C323 VTAIL.n217 B 0.047676f
C324 VTAIL.n218 B 0.050803f
C325 VTAIL.n219 B 1.34003f
C326 VTAIL.n220 B 0.026049f
C327 VTAIL.n221 B 0.019584f
C328 VTAIL.n222 B 0.010524f
C329 VTAIL.n223 B 0.024874f
C330 VTAIL.n224 B 0.011143f
C331 VTAIL.n225 B 0.019584f
C332 VTAIL.n226 B 0.010524f
C333 VTAIL.n227 B 0.024874f
C334 VTAIL.n228 B 0.011143f
C335 VTAIL.n229 B 0.019584f
C336 VTAIL.n230 B 0.010524f
C337 VTAIL.n231 B 0.024874f
C338 VTAIL.n232 B 0.011143f
C339 VTAIL.n233 B 0.019584f
C340 VTAIL.n234 B 0.010524f
C341 VTAIL.n235 B 0.024874f
C342 VTAIL.n236 B 0.011143f
C343 VTAIL.n237 B 0.019584f
C344 VTAIL.n238 B 0.010524f
C345 VTAIL.n239 B 0.024874f
C346 VTAIL.n240 B 0.011143f
C347 VTAIL.n241 B 1.1207f
C348 VTAIL.n242 B 0.010524f
C349 VTAIL.t1 B 0.0409f
C350 VTAIL.n243 B 0.119336f
C351 VTAIL.n244 B 0.014694f
C352 VTAIL.n245 B 0.018656f
C353 VTAIL.n246 B 0.024874f
C354 VTAIL.n247 B 0.011143f
C355 VTAIL.n248 B 0.010524f
C356 VTAIL.n249 B 0.019584f
C357 VTAIL.n250 B 0.019584f
C358 VTAIL.n251 B 0.010524f
C359 VTAIL.n252 B 0.011143f
C360 VTAIL.n253 B 0.024874f
C361 VTAIL.n254 B 0.024874f
C362 VTAIL.n255 B 0.011143f
C363 VTAIL.n256 B 0.010524f
C364 VTAIL.n257 B 0.019584f
C365 VTAIL.n258 B 0.019584f
C366 VTAIL.n259 B 0.010524f
C367 VTAIL.n260 B 0.011143f
C368 VTAIL.n261 B 0.024874f
C369 VTAIL.n262 B 0.024874f
C370 VTAIL.n263 B 0.011143f
C371 VTAIL.n264 B 0.010524f
C372 VTAIL.n265 B 0.019584f
C373 VTAIL.n266 B 0.019584f
C374 VTAIL.n267 B 0.010524f
C375 VTAIL.n268 B 0.011143f
C376 VTAIL.n269 B 0.024874f
C377 VTAIL.n270 B 0.024874f
C378 VTAIL.n271 B 0.011143f
C379 VTAIL.n272 B 0.010524f
C380 VTAIL.n273 B 0.019584f
C381 VTAIL.n274 B 0.019584f
C382 VTAIL.n275 B 0.010524f
C383 VTAIL.n276 B 0.011143f
C384 VTAIL.n277 B 0.024874f
C385 VTAIL.n278 B 0.024874f
C386 VTAIL.n279 B 0.011143f
C387 VTAIL.n280 B 0.010524f
C388 VTAIL.n281 B 0.019584f
C389 VTAIL.n282 B 0.019584f
C390 VTAIL.n283 B 0.010524f
C391 VTAIL.n284 B 0.011143f
C392 VTAIL.n285 B 0.024874f
C393 VTAIL.n286 B 0.05018f
C394 VTAIL.n287 B 0.011143f
C395 VTAIL.n288 B 0.020577f
C396 VTAIL.n289 B 0.047676f
C397 VTAIL.n290 B 0.050803f
C398 VTAIL.n291 B 1.34003f
C399 VTAIL.t3 B 0.205677f
C400 VTAIL.t5 B 0.205677f
C401 VTAIL.n292 B 1.79422f
C402 VTAIL.n293 B 0.518973f
C403 VTAIL.n294 B 0.026049f
C404 VTAIL.n295 B 0.019584f
C405 VTAIL.n296 B 0.010524f
C406 VTAIL.n297 B 0.024874f
C407 VTAIL.n298 B 0.011143f
C408 VTAIL.n299 B 0.019584f
C409 VTAIL.n300 B 0.010524f
C410 VTAIL.n301 B 0.024874f
C411 VTAIL.n302 B 0.011143f
C412 VTAIL.n303 B 0.019584f
C413 VTAIL.n304 B 0.010524f
C414 VTAIL.n305 B 0.024874f
C415 VTAIL.n306 B 0.011143f
C416 VTAIL.n307 B 0.019584f
C417 VTAIL.n308 B 0.010524f
C418 VTAIL.n309 B 0.024874f
C419 VTAIL.n310 B 0.011143f
C420 VTAIL.n311 B 0.019584f
C421 VTAIL.n312 B 0.010524f
C422 VTAIL.n313 B 0.024874f
C423 VTAIL.n314 B 0.011143f
C424 VTAIL.n315 B 1.1207f
C425 VTAIL.n316 B 0.010524f
C426 VTAIL.t0 B 0.0409f
C427 VTAIL.n317 B 0.119336f
C428 VTAIL.n318 B 0.014694f
C429 VTAIL.n319 B 0.018656f
C430 VTAIL.n320 B 0.024874f
C431 VTAIL.n321 B 0.011143f
C432 VTAIL.n322 B 0.010524f
C433 VTAIL.n323 B 0.019584f
C434 VTAIL.n324 B 0.019584f
C435 VTAIL.n325 B 0.010524f
C436 VTAIL.n326 B 0.011143f
C437 VTAIL.n327 B 0.024874f
C438 VTAIL.n328 B 0.024874f
C439 VTAIL.n329 B 0.011143f
C440 VTAIL.n330 B 0.010524f
C441 VTAIL.n331 B 0.019584f
C442 VTAIL.n332 B 0.019584f
C443 VTAIL.n333 B 0.010524f
C444 VTAIL.n334 B 0.011143f
C445 VTAIL.n335 B 0.024874f
C446 VTAIL.n336 B 0.024874f
C447 VTAIL.n337 B 0.011143f
C448 VTAIL.n338 B 0.010524f
C449 VTAIL.n339 B 0.019584f
C450 VTAIL.n340 B 0.019584f
C451 VTAIL.n341 B 0.010524f
C452 VTAIL.n342 B 0.011143f
C453 VTAIL.n343 B 0.024874f
C454 VTAIL.n344 B 0.024874f
C455 VTAIL.n345 B 0.011143f
C456 VTAIL.n346 B 0.010524f
C457 VTAIL.n347 B 0.019584f
C458 VTAIL.n348 B 0.019584f
C459 VTAIL.n349 B 0.010524f
C460 VTAIL.n350 B 0.011143f
C461 VTAIL.n351 B 0.024874f
C462 VTAIL.n352 B 0.024874f
C463 VTAIL.n353 B 0.011143f
C464 VTAIL.n354 B 0.010524f
C465 VTAIL.n355 B 0.019584f
C466 VTAIL.n356 B 0.019584f
C467 VTAIL.n357 B 0.010524f
C468 VTAIL.n358 B 0.011143f
C469 VTAIL.n359 B 0.024874f
C470 VTAIL.n360 B 0.05018f
C471 VTAIL.n361 B 0.011143f
C472 VTAIL.n362 B 0.020577f
C473 VTAIL.n363 B 0.047676f
C474 VTAIL.n364 B 0.050803f
C475 VTAIL.n365 B 0.214202f
C476 VTAIL.n366 B 0.026049f
C477 VTAIL.n367 B 0.019584f
C478 VTAIL.n368 B 0.010524f
C479 VTAIL.n369 B 0.024874f
C480 VTAIL.n370 B 0.011143f
C481 VTAIL.n371 B 0.019584f
C482 VTAIL.n372 B 0.010524f
C483 VTAIL.n373 B 0.024874f
C484 VTAIL.n374 B 0.011143f
C485 VTAIL.n375 B 0.019584f
C486 VTAIL.n376 B 0.010524f
C487 VTAIL.n377 B 0.024874f
C488 VTAIL.n378 B 0.011143f
C489 VTAIL.n379 B 0.019584f
C490 VTAIL.n380 B 0.010524f
C491 VTAIL.n381 B 0.024874f
C492 VTAIL.n382 B 0.011143f
C493 VTAIL.n383 B 0.019584f
C494 VTAIL.n384 B 0.010524f
C495 VTAIL.n385 B 0.024874f
C496 VTAIL.n386 B 0.011143f
C497 VTAIL.n387 B 1.1207f
C498 VTAIL.n388 B 0.010524f
C499 VTAIL.t14 B 0.0409f
C500 VTAIL.n389 B 0.119336f
C501 VTAIL.n390 B 0.014694f
C502 VTAIL.n391 B 0.018656f
C503 VTAIL.n392 B 0.024874f
C504 VTAIL.n393 B 0.011143f
C505 VTAIL.n394 B 0.010524f
C506 VTAIL.n395 B 0.019584f
C507 VTAIL.n396 B 0.019584f
C508 VTAIL.n397 B 0.010524f
C509 VTAIL.n398 B 0.011143f
C510 VTAIL.n399 B 0.024874f
C511 VTAIL.n400 B 0.024874f
C512 VTAIL.n401 B 0.011143f
C513 VTAIL.n402 B 0.010524f
C514 VTAIL.n403 B 0.019584f
C515 VTAIL.n404 B 0.019584f
C516 VTAIL.n405 B 0.010524f
C517 VTAIL.n406 B 0.011143f
C518 VTAIL.n407 B 0.024874f
C519 VTAIL.n408 B 0.024874f
C520 VTAIL.n409 B 0.011143f
C521 VTAIL.n410 B 0.010524f
C522 VTAIL.n411 B 0.019584f
C523 VTAIL.n412 B 0.019584f
C524 VTAIL.n413 B 0.010524f
C525 VTAIL.n414 B 0.011143f
C526 VTAIL.n415 B 0.024874f
C527 VTAIL.n416 B 0.024874f
C528 VTAIL.n417 B 0.011143f
C529 VTAIL.n418 B 0.010524f
C530 VTAIL.n419 B 0.019584f
C531 VTAIL.n420 B 0.019584f
C532 VTAIL.n421 B 0.010524f
C533 VTAIL.n422 B 0.011143f
C534 VTAIL.n423 B 0.024874f
C535 VTAIL.n424 B 0.024874f
C536 VTAIL.n425 B 0.011143f
C537 VTAIL.n426 B 0.010524f
C538 VTAIL.n427 B 0.019584f
C539 VTAIL.n428 B 0.019584f
C540 VTAIL.n429 B 0.010524f
C541 VTAIL.n430 B 0.011143f
C542 VTAIL.n431 B 0.024874f
C543 VTAIL.n432 B 0.05018f
C544 VTAIL.n433 B 0.011143f
C545 VTAIL.n434 B 0.020577f
C546 VTAIL.n435 B 0.047676f
C547 VTAIL.n436 B 0.050803f
C548 VTAIL.n437 B 0.214202f
C549 VTAIL.t11 B 0.205677f
C550 VTAIL.t8 B 0.205677f
C551 VTAIL.n438 B 1.79422f
C552 VTAIL.n439 B 0.518973f
C553 VTAIL.n440 B 0.026049f
C554 VTAIL.n441 B 0.019584f
C555 VTAIL.n442 B 0.010524f
C556 VTAIL.n443 B 0.024874f
C557 VTAIL.n444 B 0.011143f
C558 VTAIL.n445 B 0.019584f
C559 VTAIL.n446 B 0.010524f
C560 VTAIL.n447 B 0.024874f
C561 VTAIL.n448 B 0.011143f
C562 VTAIL.n449 B 0.019584f
C563 VTAIL.n450 B 0.010524f
C564 VTAIL.n451 B 0.024874f
C565 VTAIL.n452 B 0.011143f
C566 VTAIL.n453 B 0.019584f
C567 VTAIL.n454 B 0.010524f
C568 VTAIL.n455 B 0.024874f
C569 VTAIL.n456 B 0.011143f
C570 VTAIL.n457 B 0.019584f
C571 VTAIL.n458 B 0.010524f
C572 VTAIL.n459 B 0.024874f
C573 VTAIL.n460 B 0.011143f
C574 VTAIL.n461 B 1.1207f
C575 VTAIL.n462 B 0.010524f
C576 VTAIL.t7 B 0.0409f
C577 VTAIL.n463 B 0.119336f
C578 VTAIL.n464 B 0.014694f
C579 VTAIL.n465 B 0.018656f
C580 VTAIL.n466 B 0.024874f
C581 VTAIL.n467 B 0.011143f
C582 VTAIL.n468 B 0.010524f
C583 VTAIL.n469 B 0.019584f
C584 VTAIL.n470 B 0.019584f
C585 VTAIL.n471 B 0.010524f
C586 VTAIL.n472 B 0.011143f
C587 VTAIL.n473 B 0.024874f
C588 VTAIL.n474 B 0.024874f
C589 VTAIL.n475 B 0.011143f
C590 VTAIL.n476 B 0.010524f
C591 VTAIL.n477 B 0.019584f
C592 VTAIL.n478 B 0.019584f
C593 VTAIL.n479 B 0.010524f
C594 VTAIL.n480 B 0.011143f
C595 VTAIL.n481 B 0.024874f
C596 VTAIL.n482 B 0.024874f
C597 VTAIL.n483 B 0.011143f
C598 VTAIL.n484 B 0.010524f
C599 VTAIL.n485 B 0.019584f
C600 VTAIL.n486 B 0.019584f
C601 VTAIL.n487 B 0.010524f
C602 VTAIL.n488 B 0.011143f
C603 VTAIL.n489 B 0.024874f
C604 VTAIL.n490 B 0.024874f
C605 VTAIL.n491 B 0.011143f
C606 VTAIL.n492 B 0.010524f
C607 VTAIL.n493 B 0.019584f
C608 VTAIL.n494 B 0.019584f
C609 VTAIL.n495 B 0.010524f
C610 VTAIL.n496 B 0.011143f
C611 VTAIL.n497 B 0.024874f
C612 VTAIL.n498 B 0.024874f
C613 VTAIL.n499 B 0.011143f
C614 VTAIL.n500 B 0.010524f
C615 VTAIL.n501 B 0.019584f
C616 VTAIL.n502 B 0.019584f
C617 VTAIL.n503 B 0.010524f
C618 VTAIL.n504 B 0.011143f
C619 VTAIL.n505 B 0.024874f
C620 VTAIL.n506 B 0.05018f
C621 VTAIL.n507 B 0.011143f
C622 VTAIL.n508 B 0.020577f
C623 VTAIL.n509 B 0.047676f
C624 VTAIL.n510 B 0.050803f
C625 VTAIL.n511 B 1.34003f
C626 VTAIL.n512 B 0.026049f
C627 VTAIL.n513 B 0.019584f
C628 VTAIL.n514 B 0.010524f
C629 VTAIL.n515 B 0.024874f
C630 VTAIL.n516 B 0.011143f
C631 VTAIL.n517 B 0.019584f
C632 VTAIL.n518 B 0.010524f
C633 VTAIL.n519 B 0.024874f
C634 VTAIL.n520 B 0.011143f
C635 VTAIL.n521 B 0.019584f
C636 VTAIL.n522 B 0.010524f
C637 VTAIL.n523 B 0.024874f
C638 VTAIL.n524 B 0.011143f
C639 VTAIL.n525 B 0.019584f
C640 VTAIL.n526 B 0.010524f
C641 VTAIL.n527 B 0.024874f
C642 VTAIL.n528 B 0.011143f
C643 VTAIL.n529 B 0.019584f
C644 VTAIL.n530 B 0.010524f
C645 VTAIL.n531 B 0.024874f
C646 VTAIL.n532 B 0.011143f
C647 VTAIL.n533 B 1.1207f
C648 VTAIL.n534 B 0.010524f
C649 VTAIL.t15 B 0.0409f
C650 VTAIL.n535 B 0.119336f
C651 VTAIL.n536 B 0.014694f
C652 VTAIL.n537 B 0.018656f
C653 VTAIL.n538 B 0.024874f
C654 VTAIL.n539 B 0.011143f
C655 VTAIL.n540 B 0.010524f
C656 VTAIL.n541 B 0.019584f
C657 VTAIL.n542 B 0.019584f
C658 VTAIL.n543 B 0.010524f
C659 VTAIL.n544 B 0.011143f
C660 VTAIL.n545 B 0.024874f
C661 VTAIL.n546 B 0.024874f
C662 VTAIL.n547 B 0.011143f
C663 VTAIL.n548 B 0.010524f
C664 VTAIL.n549 B 0.019584f
C665 VTAIL.n550 B 0.019584f
C666 VTAIL.n551 B 0.010524f
C667 VTAIL.n552 B 0.011143f
C668 VTAIL.n553 B 0.024874f
C669 VTAIL.n554 B 0.024874f
C670 VTAIL.n555 B 0.011143f
C671 VTAIL.n556 B 0.010524f
C672 VTAIL.n557 B 0.019584f
C673 VTAIL.n558 B 0.019584f
C674 VTAIL.n559 B 0.010524f
C675 VTAIL.n560 B 0.011143f
C676 VTAIL.n561 B 0.024874f
C677 VTAIL.n562 B 0.024874f
C678 VTAIL.n563 B 0.011143f
C679 VTAIL.n564 B 0.010524f
C680 VTAIL.n565 B 0.019584f
C681 VTAIL.n566 B 0.019584f
C682 VTAIL.n567 B 0.010524f
C683 VTAIL.n568 B 0.011143f
C684 VTAIL.n569 B 0.024874f
C685 VTAIL.n570 B 0.024874f
C686 VTAIL.n571 B 0.011143f
C687 VTAIL.n572 B 0.010524f
C688 VTAIL.n573 B 0.019584f
C689 VTAIL.n574 B 0.019584f
C690 VTAIL.n575 B 0.010524f
C691 VTAIL.n576 B 0.011143f
C692 VTAIL.n577 B 0.024874f
C693 VTAIL.n578 B 0.05018f
C694 VTAIL.n579 B 0.011143f
C695 VTAIL.n580 B 0.020577f
C696 VTAIL.n581 B 0.047676f
C697 VTAIL.n582 B 0.050803f
C698 VTAIL.n583 B 1.33636f
C699 VDD1.t7 B 0.258277f
C700 VDD1.t1 B 0.258277f
C701 VDD1.n0 B 2.33395f
C702 VDD1.t5 B 0.258277f
C703 VDD1.t4 B 0.258277f
C704 VDD1.n1 B 2.33286f
C705 VDD1.t6 B 0.258277f
C706 VDD1.t0 B 0.258277f
C707 VDD1.n2 B 2.33286f
C708 VDD1.n3 B 3.41963f
C709 VDD1.t3 B 0.258277f
C710 VDD1.t2 B 0.258277f
C711 VDD1.n4 B 2.32268f
C712 VDD1.n5 B 3.06851f
C713 VP.n0 B 0.028496f
C714 VP.t4 B 2.14257f
C715 VP.n1 B 0.04122f
C716 VP.n2 B 0.021614f
C717 VP.t1 B 2.14257f
C718 VP.n3 B 0.75245f
C719 VP.n4 B 0.021614f
C720 VP.n5 B 0.017473f
C721 VP.n6 B 0.021614f
C722 VP.t5 B 2.14257f
C723 VP.n7 B 0.75245f
C724 VP.n8 B 0.021614f
C725 VP.n9 B 0.04122f
C726 VP.n10 B 0.028496f
C727 VP.t2 B 2.14257f
C728 VP.n11 B 0.028496f
C729 VP.t7 B 2.14257f
C730 VP.n12 B 0.04122f
C731 VP.n13 B 0.021614f
C732 VP.t6 B 2.14257f
C733 VP.n14 B 0.75245f
C734 VP.n15 B 0.021614f
C735 VP.n16 B 0.017473f
C736 VP.n17 B 0.021614f
C737 VP.t3 B 2.14257f
C738 VP.n18 B 0.809428f
C739 VP.t0 B 2.33145f
C740 VP.n19 B 0.794914f
C741 VP.n20 B 0.211698f
C742 VP.n21 B 0.021588f
C743 VP.n22 B 0.040283f
C744 VP.n23 B 0.042958f
C745 VP.n24 B 0.021614f
C746 VP.n25 B 0.021614f
C747 VP.n26 B 0.021614f
C748 VP.n27 B 0.042958f
C749 VP.n28 B 0.040283f
C750 VP.n29 B 0.021588f
C751 VP.n30 B 0.021614f
C752 VP.n31 B 0.021614f
C753 VP.n32 B 0.03909f
C754 VP.n33 B 0.043675f
C755 VP.n34 B 0.018493f
C756 VP.n35 B 0.021614f
C757 VP.n36 B 0.021614f
C758 VP.n37 B 0.021614f
C759 VP.n38 B 0.040283f
C760 VP.n39 B 0.023975f
C761 VP.n40 B 0.822098f
C762 VP.n41 B 1.29274f
C763 VP.n42 B 1.30755f
C764 VP.n43 B 0.822098f
C765 VP.n44 B 0.023975f
C766 VP.n45 B 0.040283f
C767 VP.n46 B 0.021614f
C768 VP.n47 B 0.021614f
C769 VP.n48 B 0.021614f
C770 VP.n49 B 0.018493f
C771 VP.n50 B 0.043675f
C772 VP.n51 B 0.03909f
C773 VP.n52 B 0.021614f
C774 VP.n53 B 0.021614f
C775 VP.n54 B 0.021588f
C776 VP.n55 B 0.040283f
C777 VP.n56 B 0.042958f
C778 VP.n57 B 0.021614f
C779 VP.n58 B 0.021614f
C780 VP.n59 B 0.021614f
C781 VP.n60 B 0.042958f
C782 VP.n61 B 0.040283f
C783 VP.n62 B 0.021588f
C784 VP.n63 B 0.021614f
C785 VP.n64 B 0.021614f
C786 VP.n65 B 0.03909f
C787 VP.n66 B 0.043675f
C788 VP.n67 B 0.018493f
C789 VP.n68 B 0.021614f
C790 VP.n69 B 0.021614f
C791 VP.n70 B 0.021614f
C792 VP.n71 B 0.040283f
C793 VP.n72 B 0.023975f
C794 VP.n73 B 0.822098f
C795 VP.n74 B 0.039018f
.ends

