* NGSPICE file created from diff_pair_sample_1627.ext - technology: sky130A

.subckt diff_pair_sample_1627 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X1 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X2 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=1.11
X3 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=1.11
X4 VTAIL.t11 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X5 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=1.11
X6 VDD2.t6 VN.t1 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X7 VTAIL.t14 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=1.11
X8 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=1.11
X9 VTAIL.t3 VN.t3 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X10 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X11 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=1.11
X12 VDD1.t4 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=1.11
X13 VDD1.t3 VP.t4 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=2.9523 ps=15.92 w=7.57 l=1.11
X14 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=1.11
X15 VDD1.t2 VP.t5 VTAIL.t13 B.t21 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X16 VTAIL.t7 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=1.11
X17 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=1.24905 ps=7.9 w=7.57 l=1.11
X18 VTAIL.t8 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.24905 pd=7.9 as=1.24905 ps=7.9 w=7.57 l=1.11
X19 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9523 pd=15.92 as=0 ps=0 w=7.57 l=1.11
R0 VP.n7 VP.t6 222.696
R1 VP.n17 VP.t2 199.965
R2 VP.n29 VP.t3 199.965
R3 VP.n15 VP.t4 199.965
R4 VP.n22 VP.t0 164.358
R5 VP.n1 VP.t1 164.358
R6 VP.n5 VP.t7 164.358
R7 VP.n8 VP.t5 164.358
R8 VP.n9 VP.n6 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n4 161.3
R12 VP.n28 VP.n0 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n25 VP.n24 161.3
R15 VP.n23 VP.n2 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n19 VP.n3 161.3
R18 VP.n16 VP.n15 80.6037
R19 VP.n30 VP.n29 80.6037
R20 VP.n18 VP.n17 80.6037
R21 VP.n24 VP.n23 56.5193
R22 VP.n10 VP.n9 56.5193
R23 VP.n17 VP.n3 49.4239
R24 VP.n29 VP.n28 49.4239
R25 VP.n15 VP.n14 49.4239
R26 VP.n18 VP.n16 40.7438
R27 VP.n8 VP.n7 33.8527
R28 VP.n7 VP.n6 28.2774
R29 VP.n21 VP.n3 24.4675
R30 VP.n28 VP.n27 24.4675
R31 VP.n14 VP.n13 24.4675
R32 VP.n23 VP.n22 22.9995
R33 VP.n24 VP.n1 22.9995
R34 VP.n10 VP.n5 22.9995
R35 VP.n9 VP.n8 22.9995
R36 VP.n22 VP.n21 1.46852
R37 VP.n27 VP.n1 1.46852
R38 VP.n13 VP.n5 1.46852
R39 VP.n16 VP.n4 0.285035
R40 VP.n19 VP.n18 0.285035
R41 VP.n30 VP.n0 0.285035
R42 VP.n11 VP.n6 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n20 VP.n2 0.189894
R47 VP.n25 VP.n2 0.189894
R48 VP.n26 VP.n25 0.189894
R49 VP.n26 VP.n0 0.189894
R50 VP VP.n30 0.146778
R51 VTAIL.n11 VTAIL.t7 52.7493
R52 VTAIL.n10 VTAIL.t2 52.7493
R53 VTAIL.n7 VTAIL.t5 52.7493
R54 VTAIL.n15 VTAIL.t1 52.7491
R55 VTAIL.n2 VTAIL.t4 52.7491
R56 VTAIL.n3 VTAIL.t12 52.7491
R57 VTAIL.n6 VTAIL.t14 52.7491
R58 VTAIL.n14 VTAIL.t9 52.7491
R59 VTAIL.n13 VTAIL.n12 50.1337
R60 VTAIL.n9 VTAIL.n8 50.1337
R61 VTAIL.n1 VTAIL.n0 50.1335
R62 VTAIL.n5 VTAIL.n4 50.1335
R63 VTAIL.n15 VTAIL.n14 20.1341
R64 VTAIL.n7 VTAIL.n6 20.1341
R65 VTAIL.n0 VTAIL.t15 2.61609
R66 VTAIL.n0 VTAIL.t6 2.61609
R67 VTAIL.n4 VTAIL.t10 2.61609
R68 VTAIL.n4 VTAIL.t11 2.61609
R69 VTAIL.n12 VTAIL.t13 2.61609
R70 VTAIL.n12 VTAIL.t8 2.61609
R71 VTAIL.n8 VTAIL.t0 2.61609
R72 VTAIL.n8 VTAIL.t3 2.61609
R73 VTAIL.n9 VTAIL.n7 1.24188
R74 VTAIL.n10 VTAIL.n9 1.24188
R75 VTAIL.n13 VTAIL.n11 1.24188
R76 VTAIL.n14 VTAIL.n13 1.24188
R77 VTAIL.n6 VTAIL.n5 1.24188
R78 VTAIL.n5 VTAIL.n3 1.24188
R79 VTAIL.n2 VTAIL.n1 1.24188
R80 VTAIL VTAIL.n15 1.18369
R81 VTAIL.n11 VTAIL.n10 0.470328
R82 VTAIL.n3 VTAIL.n2 0.470328
R83 VTAIL VTAIL.n1 0.0586897
R84 VDD1 VDD1.n0 67.4914
R85 VDD1.n3 VDD1.n2 67.3776
R86 VDD1.n3 VDD1.n1 67.3776
R87 VDD1.n5 VDD1.n4 66.8123
R88 VDD1.n5 VDD1.n3 36.4104
R89 VDD1.n4 VDD1.t0 2.61609
R90 VDD1.n4 VDD1.t3 2.61609
R91 VDD1.n0 VDD1.t1 2.61609
R92 VDD1.n0 VDD1.t2 2.61609
R93 VDD1.n2 VDD1.t6 2.61609
R94 VDD1.n2 VDD1.t4 2.61609
R95 VDD1.n1 VDD1.t5 2.61609
R96 VDD1.n1 VDD1.t7 2.61609
R97 VDD1 VDD1.n5 0.563
R98 B.n581 B.n580 585
R99 B.n582 B.n581 585
R100 B.n226 B.n89 585
R101 B.n225 B.n224 585
R102 B.n223 B.n222 585
R103 B.n221 B.n220 585
R104 B.n219 B.n218 585
R105 B.n217 B.n216 585
R106 B.n215 B.n214 585
R107 B.n213 B.n212 585
R108 B.n211 B.n210 585
R109 B.n209 B.n208 585
R110 B.n207 B.n206 585
R111 B.n205 B.n204 585
R112 B.n203 B.n202 585
R113 B.n201 B.n200 585
R114 B.n199 B.n198 585
R115 B.n197 B.n196 585
R116 B.n195 B.n194 585
R117 B.n193 B.n192 585
R118 B.n191 B.n190 585
R119 B.n189 B.n188 585
R120 B.n187 B.n186 585
R121 B.n185 B.n184 585
R122 B.n183 B.n182 585
R123 B.n181 B.n180 585
R124 B.n179 B.n178 585
R125 B.n177 B.n176 585
R126 B.n175 B.n174 585
R127 B.n173 B.n172 585
R128 B.n171 B.n170 585
R129 B.n169 B.n168 585
R130 B.n167 B.n166 585
R131 B.n165 B.n164 585
R132 B.n163 B.n162 585
R133 B.n161 B.n160 585
R134 B.n159 B.n158 585
R135 B.n157 B.n156 585
R136 B.n155 B.n154 585
R137 B.n152 B.n151 585
R138 B.n150 B.n149 585
R139 B.n148 B.n147 585
R140 B.n146 B.n145 585
R141 B.n144 B.n143 585
R142 B.n142 B.n141 585
R143 B.n140 B.n139 585
R144 B.n138 B.n137 585
R145 B.n136 B.n135 585
R146 B.n134 B.n133 585
R147 B.n132 B.n131 585
R148 B.n130 B.n129 585
R149 B.n128 B.n127 585
R150 B.n126 B.n125 585
R151 B.n124 B.n123 585
R152 B.n122 B.n121 585
R153 B.n120 B.n119 585
R154 B.n118 B.n117 585
R155 B.n116 B.n115 585
R156 B.n114 B.n113 585
R157 B.n112 B.n111 585
R158 B.n110 B.n109 585
R159 B.n108 B.n107 585
R160 B.n106 B.n105 585
R161 B.n104 B.n103 585
R162 B.n102 B.n101 585
R163 B.n100 B.n99 585
R164 B.n98 B.n97 585
R165 B.n96 B.n95 585
R166 B.n579 B.n55 585
R167 B.n583 B.n55 585
R168 B.n578 B.n54 585
R169 B.n584 B.n54 585
R170 B.n577 B.n576 585
R171 B.n576 B.n50 585
R172 B.n575 B.n49 585
R173 B.n590 B.n49 585
R174 B.n574 B.n48 585
R175 B.n591 B.n48 585
R176 B.n573 B.n47 585
R177 B.n592 B.n47 585
R178 B.n572 B.n571 585
R179 B.n571 B.n43 585
R180 B.n570 B.n42 585
R181 B.n598 B.n42 585
R182 B.n569 B.n41 585
R183 B.n599 B.n41 585
R184 B.n568 B.n40 585
R185 B.n600 B.n40 585
R186 B.n567 B.n566 585
R187 B.n566 B.n36 585
R188 B.n565 B.n35 585
R189 B.n606 B.n35 585
R190 B.n564 B.n34 585
R191 B.n607 B.n34 585
R192 B.n563 B.n33 585
R193 B.n608 B.n33 585
R194 B.n562 B.n561 585
R195 B.n561 B.n29 585
R196 B.n560 B.n28 585
R197 B.n614 B.n28 585
R198 B.n559 B.n27 585
R199 B.n615 B.n27 585
R200 B.n558 B.n26 585
R201 B.n616 B.n26 585
R202 B.n557 B.n556 585
R203 B.n556 B.n22 585
R204 B.n555 B.n21 585
R205 B.n622 B.n21 585
R206 B.n554 B.n20 585
R207 B.n623 B.n20 585
R208 B.n553 B.n19 585
R209 B.n624 B.n19 585
R210 B.n552 B.n551 585
R211 B.n551 B.n15 585
R212 B.n550 B.n14 585
R213 B.n630 B.n14 585
R214 B.n549 B.n13 585
R215 B.n631 B.n13 585
R216 B.n548 B.n12 585
R217 B.n632 B.n12 585
R218 B.n547 B.n546 585
R219 B.n546 B.n8 585
R220 B.n545 B.n7 585
R221 B.n638 B.n7 585
R222 B.n544 B.n6 585
R223 B.n639 B.n6 585
R224 B.n543 B.n5 585
R225 B.n640 B.n5 585
R226 B.n542 B.n541 585
R227 B.n541 B.n4 585
R228 B.n540 B.n227 585
R229 B.n540 B.n539 585
R230 B.n530 B.n228 585
R231 B.n229 B.n228 585
R232 B.n532 B.n531 585
R233 B.n533 B.n532 585
R234 B.n529 B.n234 585
R235 B.n234 B.n233 585
R236 B.n528 B.n527 585
R237 B.n527 B.n526 585
R238 B.n236 B.n235 585
R239 B.n237 B.n236 585
R240 B.n519 B.n518 585
R241 B.n520 B.n519 585
R242 B.n517 B.n242 585
R243 B.n242 B.n241 585
R244 B.n516 B.n515 585
R245 B.n515 B.n514 585
R246 B.n244 B.n243 585
R247 B.n245 B.n244 585
R248 B.n507 B.n506 585
R249 B.n508 B.n507 585
R250 B.n505 B.n249 585
R251 B.n253 B.n249 585
R252 B.n504 B.n503 585
R253 B.n503 B.n502 585
R254 B.n251 B.n250 585
R255 B.n252 B.n251 585
R256 B.n495 B.n494 585
R257 B.n496 B.n495 585
R258 B.n493 B.n257 585
R259 B.n261 B.n257 585
R260 B.n492 B.n491 585
R261 B.n491 B.n490 585
R262 B.n259 B.n258 585
R263 B.n260 B.n259 585
R264 B.n483 B.n482 585
R265 B.n484 B.n483 585
R266 B.n481 B.n266 585
R267 B.n266 B.n265 585
R268 B.n480 B.n479 585
R269 B.n479 B.n478 585
R270 B.n268 B.n267 585
R271 B.n269 B.n268 585
R272 B.n471 B.n470 585
R273 B.n472 B.n471 585
R274 B.n469 B.n274 585
R275 B.n274 B.n273 585
R276 B.n468 B.n467 585
R277 B.n467 B.n466 585
R278 B.n276 B.n275 585
R279 B.n277 B.n276 585
R280 B.n459 B.n458 585
R281 B.n460 B.n459 585
R282 B.n457 B.n282 585
R283 B.n282 B.n281 585
R284 B.n451 B.n450 585
R285 B.n449 B.n317 585
R286 B.n448 B.n316 585
R287 B.n453 B.n316 585
R288 B.n447 B.n446 585
R289 B.n445 B.n444 585
R290 B.n443 B.n442 585
R291 B.n441 B.n440 585
R292 B.n439 B.n438 585
R293 B.n437 B.n436 585
R294 B.n435 B.n434 585
R295 B.n433 B.n432 585
R296 B.n431 B.n430 585
R297 B.n429 B.n428 585
R298 B.n427 B.n426 585
R299 B.n425 B.n424 585
R300 B.n423 B.n422 585
R301 B.n421 B.n420 585
R302 B.n419 B.n418 585
R303 B.n417 B.n416 585
R304 B.n415 B.n414 585
R305 B.n413 B.n412 585
R306 B.n411 B.n410 585
R307 B.n409 B.n408 585
R308 B.n407 B.n406 585
R309 B.n405 B.n404 585
R310 B.n403 B.n402 585
R311 B.n401 B.n400 585
R312 B.n399 B.n398 585
R313 B.n397 B.n396 585
R314 B.n395 B.n394 585
R315 B.n393 B.n392 585
R316 B.n391 B.n390 585
R317 B.n389 B.n388 585
R318 B.n387 B.n386 585
R319 B.n385 B.n384 585
R320 B.n383 B.n382 585
R321 B.n381 B.n380 585
R322 B.n379 B.n378 585
R323 B.n376 B.n375 585
R324 B.n374 B.n373 585
R325 B.n372 B.n371 585
R326 B.n370 B.n369 585
R327 B.n368 B.n367 585
R328 B.n366 B.n365 585
R329 B.n364 B.n363 585
R330 B.n362 B.n361 585
R331 B.n360 B.n359 585
R332 B.n358 B.n357 585
R333 B.n356 B.n355 585
R334 B.n354 B.n353 585
R335 B.n352 B.n351 585
R336 B.n350 B.n349 585
R337 B.n348 B.n347 585
R338 B.n346 B.n345 585
R339 B.n344 B.n343 585
R340 B.n342 B.n341 585
R341 B.n340 B.n339 585
R342 B.n338 B.n337 585
R343 B.n336 B.n335 585
R344 B.n334 B.n333 585
R345 B.n332 B.n331 585
R346 B.n330 B.n329 585
R347 B.n328 B.n327 585
R348 B.n326 B.n325 585
R349 B.n324 B.n323 585
R350 B.n284 B.n283 585
R351 B.n456 B.n455 585
R352 B.n280 B.n279 585
R353 B.n281 B.n280 585
R354 B.n462 B.n461 585
R355 B.n461 B.n460 585
R356 B.n463 B.n278 585
R357 B.n278 B.n277 585
R358 B.n465 B.n464 585
R359 B.n466 B.n465 585
R360 B.n272 B.n271 585
R361 B.n273 B.n272 585
R362 B.n474 B.n473 585
R363 B.n473 B.n472 585
R364 B.n475 B.n270 585
R365 B.n270 B.n269 585
R366 B.n477 B.n476 585
R367 B.n478 B.n477 585
R368 B.n264 B.n263 585
R369 B.n265 B.n264 585
R370 B.n486 B.n485 585
R371 B.n485 B.n484 585
R372 B.n487 B.n262 585
R373 B.n262 B.n260 585
R374 B.n489 B.n488 585
R375 B.n490 B.n489 585
R376 B.n256 B.n255 585
R377 B.n261 B.n256 585
R378 B.n498 B.n497 585
R379 B.n497 B.n496 585
R380 B.n499 B.n254 585
R381 B.n254 B.n252 585
R382 B.n501 B.n500 585
R383 B.n502 B.n501 585
R384 B.n248 B.n247 585
R385 B.n253 B.n248 585
R386 B.n510 B.n509 585
R387 B.n509 B.n508 585
R388 B.n511 B.n246 585
R389 B.n246 B.n245 585
R390 B.n513 B.n512 585
R391 B.n514 B.n513 585
R392 B.n240 B.n239 585
R393 B.n241 B.n240 585
R394 B.n522 B.n521 585
R395 B.n521 B.n520 585
R396 B.n523 B.n238 585
R397 B.n238 B.n237 585
R398 B.n525 B.n524 585
R399 B.n526 B.n525 585
R400 B.n232 B.n231 585
R401 B.n233 B.n232 585
R402 B.n535 B.n534 585
R403 B.n534 B.n533 585
R404 B.n536 B.n230 585
R405 B.n230 B.n229 585
R406 B.n538 B.n537 585
R407 B.n539 B.n538 585
R408 B.n2 B.n0 585
R409 B.n4 B.n2 585
R410 B.n3 B.n1 585
R411 B.n639 B.n3 585
R412 B.n637 B.n636 585
R413 B.n638 B.n637 585
R414 B.n635 B.n9 585
R415 B.n9 B.n8 585
R416 B.n634 B.n633 585
R417 B.n633 B.n632 585
R418 B.n11 B.n10 585
R419 B.n631 B.n11 585
R420 B.n629 B.n628 585
R421 B.n630 B.n629 585
R422 B.n627 B.n16 585
R423 B.n16 B.n15 585
R424 B.n626 B.n625 585
R425 B.n625 B.n624 585
R426 B.n18 B.n17 585
R427 B.n623 B.n18 585
R428 B.n621 B.n620 585
R429 B.n622 B.n621 585
R430 B.n619 B.n23 585
R431 B.n23 B.n22 585
R432 B.n618 B.n617 585
R433 B.n617 B.n616 585
R434 B.n25 B.n24 585
R435 B.n615 B.n25 585
R436 B.n613 B.n612 585
R437 B.n614 B.n613 585
R438 B.n611 B.n30 585
R439 B.n30 B.n29 585
R440 B.n610 B.n609 585
R441 B.n609 B.n608 585
R442 B.n32 B.n31 585
R443 B.n607 B.n32 585
R444 B.n605 B.n604 585
R445 B.n606 B.n605 585
R446 B.n603 B.n37 585
R447 B.n37 B.n36 585
R448 B.n602 B.n601 585
R449 B.n601 B.n600 585
R450 B.n39 B.n38 585
R451 B.n599 B.n39 585
R452 B.n597 B.n596 585
R453 B.n598 B.n597 585
R454 B.n595 B.n44 585
R455 B.n44 B.n43 585
R456 B.n594 B.n593 585
R457 B.n593 B.n592 585
R458 B.n46 B.n45 585
R459 B.n591 B.n46 585
R460 B.n589 B.n588 585
R461 B.n590 B.n589 585
R462 B.n587 B.n51 585
R463 B.n51 B.n50 585
R464 B.n586 B.n585 585
R465 B.n585 B.n584 585
R466 B.n53 B.n52 585
R467 B.n583 B.n53 585
R468 B.n642 B.n641 585
R469 B.n641 B.n640 585
R470 B.n451 B.n280 526.135
R471 B.n95 B.n53 526.135
R472 B.n455 B.n282 526.135
R473 B.n581 B.n55 526.135
R474 B.n321 B.t7 367.978
R475 B.n318 B.t11 367.978
R476 B.n93 B.t14 367.978
R477 B.n90 B.t18 367.978
R478 B.n582 B.n88 256.663
R479 B.n582 B.n87 256.663
R480 B.n582 B.n86 256.663
R481 B.n582 B.n85 256.663
R482 B.n582 B.n84 256.663
R483 B.n582 B.n83 256.663
R484 B.n582 B.n82 256.663
R485 B.n582 B.n81 256.663
R486 B.n582 B.n80 256.663
R487 B.n582 B.n79 256.663
R488 B.n582 B.n78 256.663
R489 B.n582 B.n77 256.663
R490 B.n582 B.n76 256.663
R491 B.n582 B.n75 256.663
R492 B.n582 B.n74 256.663
R493 B.n582 B.n73 256.663
R494 B.n582 B.n72 256.663
R495 B.n582 B.n71 256.663
R496 B.n582 B.n70 256.663
R497 B.n582 B.n69 256.663
R498 B.n582 B.n68 256.663
R499 B.n582 B.n67 256.663
R500 B.n582 B.n66 256.663
R501 B.n582 B.n65 256.663
R502 B.n582 B.n64 256.663
R503 B.n582 B.n63 256.663
R504 B.n582 B.n62 256.663
R505 B.n582 B.n61 256.663
R506 B.n582 B.n60 256.663
R507 B.n582 B.n59 256.663
R508 B.n582 B.n58 256.663
R509 B.n582 B.n57 256.663
R510 B.n582 B.n56 256.663
R511 B.n453 B.n452 256.663
R512 B.n453 B.n285 256.663
R513 B.n453 B.n286 256.663
R514 B.n453 B.n287 256.663
R515 B.n453 B.n288 256.663
R516 B.n453 B.n289 256.663
R517 B.n453 B.n290 256.663
R518 B.n453 B.n291 256.663
R519 B.n453 B.n292 256.663
R520 B.n453 B.n293 256.663
R521 B.n453 B.n294 256.663
R522 B.n453 B.n295 256.663
R523 B.n453 B.n296 256.663
R524 B.n453 B.n297 256.663
R525 B.n453 B.n298 256.663
R526 B.n453 B.n299 256.663
R527 B.n453 B.n300 256.663
R528 B.n453 B.n301 256.663
R529 B.n453 B.n302 256.663
R530 B.n453 B.n303 256.663
R531 B.n453 B.n304 256.663
R532 B.n453 B.n305 256.663
R533 B.n453 B.n306 256.663
R534 B.n453 B.n307 256.663
R535 B.n453 B.n308 256.663
R536 B.n453 B.n309 256.663
R537 B.n453 B.n310 256.663
R538 B.n453 B.n311 256.663
R539 B.n453 B.n312 256.663
R540 B.n453 B.n313 256.663
R541 B.n453 B.n314 256.663
R542 B.n453 B.n315 256.663
R543 B.n454 B.n453 256.663
R544 B.n461 B.n280 163.367
R545 B.n461 B.n278 163.367
R546 B.n465 B.n278 163.367
R547 B.n465 B.n272 163.367
R548 B.n473 B.n272 163.367
R549 B.n473 B.n270 163.367
R550 B.n477 B.n270 163.367
R551 B.n477 B.n264 163.367
R552 B.n485 B.n264 163.367
R553 B.n485 B.n262 163.367
R554 B.n489 B.n262 163.367
R555 B.n489 B.n256 163.367
R556 B.n497 B.n256 163.367
R557 B.n497 B.n254 163.367
R558 B.n501 B.n254 163.367
R559 B.n501 B.n248 163.367
R560 B.n509 B.n248 163.367
R561 B.n509 B.n246 163.367
R562 B.n513 B.n246 163.367
R563 B.n513 B.n240 163.367
R564 B.n521 B.n240 163.367
R565 B.n521 B.n238 163.367
R566 B.n525 B.n238 163.367
R567 B.n525 B.n232 163.367
R568 B.n534 B.n232 163.367
R569 B.n534 B.n230 163.367
R570 B.n538 B.n230 163.367
R571 B.n538 B.n2 163.367
R572 B.n641 B.n2 163.367
R573 B.n641 B.n3 163.367
R574 B.n637 B.n3 163.367
R575 B.n637 B.n9 163.367
R576 B.n633 B.n9 163.367
R577 B.n633 B.n11 163.367
R578 B.n629 B.n11 163.367
R579 B.n629 B.n16 163.367
R580 B.n625 B.n16 163.367
R581 B.n625 B.n18 163.367
R582 B.n621 B.n18 163.367
R583 B.n621 B.n23 163.367
R584 B.n617 B.n23 163.367
R585 B.n617 B.n25 163.367
R586 B.n613 B.n25 163.367
R587 B.n613 B.n30 163.367
R588 B.n609 B.n30 163.367
R589 B.n609 B.n32 163.367
R590 B.n605 B.n32 163.367
R591 B.n605 B.n37 163.367
R592 B.n601 B.n37 163.367
R593 B.n601 B.n39 163.367
R594 B.n597 B.n39 163.367
R595 B.n597 B.n44 163.367
R596 B.n593 B.n44 163.367
R597 B.n593 B.n46 163.367
R598 B.n589 B.n46 163.367
R599 B.n589 B.n51 163.367
R600 B.n585 B.n51 163.367
R601 B.n585 B.n53 163.367
R602 B.n317 B.n316 163.367
R603 B.n446 B.n316 163.367
R604 B.n444 B.n443 163.367
R605 B.n440 B.n439 163.367
R606 B.n436 B.n435 163.367
R607 B.n432 B.n431 163.367
R608 B.n428 B.n427 163.367
R609 B.n424 B.n423 163.367
R610 B.n420 B.n419 163.367
R611 B.n416 B.n415 163.367
R612 B.n412 B.n411 163.367
R613 B.n408 B.n407 163.367
R614 B.n404 B.n403 163.367
R615 B.n400 B.n399 163.367
R616 B.n396 B.n395 163.367
R617 B.n392 B.n391 163.367
R618 B.n388 B.n387 163.367
R619 B.n384 B.n383 163.367
R620 B.n380 B.n379 163.367
R621 B.n375 B.n374 163.367
R622 B.n371 B.n370 163.367
R623 B.n367 B.n366 163.367
R624 B.n363 B.n362 163.367
R625 B.n359 B.n358 163.367
R626 B.n355 B.n354 163.367
R627 B.n351 B.n350 163.367
R628 B.n347 B.n346 163.367
R629 B.n343 B.n342 163.367
R630 B.n339 B.n338 163.367
R631 B.n335 B.n334 163.367
R632 B.n331 B.n330 163.367
R633 B.n327 B.n326 163.367
R634 B.n323 B.n284 163.367
R635 B.n459 B.n282 163.367
R636 B.n459 B.n276 163.367
R637 B.n467 B.n276 163.367
R638 B.n467 B.n274 163.367
R639 B.n471 B.n274 163.367
R640 B.n471 B.n268 163.367
R641 B.n479 B.n268 163.367
R642 B.n479 B.n266 163.367
R643 B.n483 B.n266 163.367
R644 B.n483 B.n259 163.367
R645 B.n491 B.n259 163.367
R646 B.n491 B.n257 163.367
R647 B.n495 B.n257 163.367
R648 B.n495 B.n251 163.367
R649 B.n503 B.n251 163.367
R650 B.n503 B.n249 163.367
R651 B.n507 B.n249 163.367
R652 B.n507 B.n244 163.367
R653 B.n515 B.n244 163.367
R654 B.n515 B.n242 163.367
R655 B.n519 B.n242 163.367
R656 B.n519 B.n236 163.367
R657 B.n527 B.n236 163.367
R658 B.n527 B.n234 163.367
R659 B.n532 B.n234 163.367
R660 B.n532 B.n228 163.367
R661 B.n540 B.n228 163.367
R662 B.n541 B.n540 163.367
R663 B.n541 B.n5 163.367
R664 B.n6 B.n5 163.367
R665 B.n7 B.n6 163.367
R666 B.n546 B.n7 163.367
R667 B.n546 B.n12 163.367
R668 B.n13 B.n12 163.367
R669 B.n14 B.n13 163.367
R670 B.n551 B.n14 163.367
R671 B.n551 B.n19 163.367
R672 B.n20 B.n19 163.367
R673 B.n21 B.n20 163.367
R674 B.n556 B.n21 163.367
R675 B.n556 B.n26 163.367
R676 B.n27 B.n26 163.367
R677 B.n28 B.n27 163.367
R678 B.n561 B.n28 163.367
R679 B.n561 B.n33 163.367
R680 B.n34 B.n33 163.367
R681 B.n35 B.n34 163.367
R682 B.n566 B.n35 163.367
R683 B.n566 B.n40 163.367
R684 B.n41 B.n40 163.367
R685 B.n42 B.n41 163.367
R686 B.n571 B.n42 163.367
R687 B.n571 B.n47 163.367
R688 B.n48 B.n47 163.367
R689 B.n49 B.n48 163.367
R690 B.n576 B.n49 163.367
R691 B.n576 B.n54 163.367
R692 B.n55 B.n54 163.367
R693 B.n99 B.n98 163.367
R694 B.n103 B.n102 163.367
R695 B.n107 B.n106 163.367
R696 B.n111 B.n110 163.367
R697 B.n115 B.n114 163.367
R698 B.n119 B.n118 163.367
R699 B.n123 B.n122 163.367
R700 B.n127 B.n126 163.367
R701 B.n131 B.n130 163.367
R702 B.n135 B.n134 163.367
R703 B.n139 B.n138 163.367
R704 B.n143 B.n142 163.367
R705 B.n147 B.n146 163.367
R706 B.n151 B.n150 163.367
R707 B.n156 B.n155 163.367
R708 B.n160 B.n159 163.367
R709 B.n164 B.n163 163.367
R710 B.n168 B.n167 163.367
R711 B.n172 B.n171 163.367
R712 B.n176 B.n175 163.367
R713 B.n180 B.n179 163.367
R714 B.n184 B.n183 163.367
R715 B.n188 B.n187 163.367
R716 B.n192 B.n191 163.367
R717 B.n196 B.n195 163.367
R718 B.n200 B.n199 163.367
R719 B.n204 B.n203 163.367
R720 B.n208 B.n207 163.367
R721 B.n212 B.n211 163.367
R722 B.n216 B.n215 163.367
R723 B.n220 B.n219 163.367
R724 B.n224 B.n223 163.367
R725 B.n581 B.n89 163.367
R726 B.n453 B.n281 122.46
R727 B.n583 B.n582 122.46
R728 B.n321 B.t10 98.4231
R729 B.n90 B.t19 98.4231
R730 B.n318 B.t13 98.4144
R731 B.n93 B.t16 98.4144
R732 B.n452 B.n451 71.676
R733 B.n446 B.n285 71.676
R734 B.n443 B.n286 71.676
R735 B.n439 B.n287 71.676
R736 B.n435 B.n288 71.676
R737 B.n431 B.n289 71.676
R738 B.n427 B.n290 71.676
R739 B.n423 B.n291 71.676
R740 B.n419 B.n292 71.676
R741 B.n415 B.n293 71.676
R742 B.n411 B.n294 71.676
R743 B.n407 B.n295 71.676
R744 B.n403 B.n296 71.676
R745 B.n399 B.n297 71.676
R746 B.n395 B.n298 71.676
R747 B.n391 B.n299 71.676
R748 B.n387 B.n300 71.676
R749 B.n383 B.n301 71.676
R750 B.n379 B.n302 71.676
R751 B.n374 B.n303 71.676
R752 B.n370 B.n304 71.676
R753 B.n366 B.n305 71.676
R754 B.n362 B.n306 71.676
R755 B.n358 B.n307 71.676
R756 B.n354 B.n308 71.676
R757 B.n350 B.n309 71.676
R758 B.n346 B.n310 71.676
R759 B.n342 B.n311 71.676
R760 B.n338 B.n312 71.676
R761 B.n334 B.n313 71.676
R762 B.n330 B.n314 71.676
R763 B.n326 B.n315 71.676
R764 B.n454 B.n284 71.676
R765 B.n95 B.n56 71.676
R766 B.n99 B.n57 71.676
R767 B.n103 B.n58 71.676
R768 B.n107 B.n59 71.676
R769 B.n111 B.n60 71.676
R770 B.n115 B.n61 71.676
R771 B.n119 B.n62 71.676
R772 B.n123 B.n63 71.676
R773 B.n127 B.n64 71.676
R774 B.n131 B.n65 71.676
R775 B.n135 B.n66 71.676
R776 B.n139 B.n67 71.676
R777 B.n143 B.n68 71.676
R778 B.n147 B.n69 71.676
R779 B.n151 B.n70 71.676
R780 B.n156 B.n71 71.676
R781 B.n160 B.n72 71.676
R782 B.n164 B.n73 71.676
R783 B.n168 B.n74 71.676
R784 B.n172 B.n75 71.676
R785 B.n176 B.n76 71.676
R786 B.n180 B.n77 71.676
R787 B.n184 B.n78 71.676
R788 B.n188 B.n79 71.676
R789 B.n192 B.n80 71.676
R790 B.n196 B.n81 71.676
R791 B.n200 B.n82 71.676
R792 B.n204 B.n83 71.676
R793 B.n208 B.n84 71.676
R794 B.n212 B.n85 71.676
R795 B.n216 B.n86 71.676
R796 B.n220 B.n87 71.676
R797 B.n224 B.n88 71.676
R798 B.n89 B.n88 71.676
R799 B.n223 B.n87 71.676
R800 B.n219 B.n86 71.676
R801 B.n215 B.n85 71.676
R802 B.n211 B.n84 71.676
R803 B.n207 B.n83 71.676
R804 B.n203 B.n82 71.676
R805 B.n199 B.n81 71.676
R806 B.n195 B.n80 71.676
R807 B.n191 B.n79 71.676
R808 B.n187 B.n78 71.676
R809 B.n183 B.n77 71.676
R810 B.n179 B.n76 71.676
R811 B.n175 B.n75 71.676
R812 B.n171 B.n74 71.676
R813 B.n167 B.n73 71.676
R814 B.n163 B.n72 71.676
R815 B.n159 B.n71 71.676
R816 B.n155 B.n70 71.676
R817 B.n150 B.n69 71.676
R818 B.n146 B.n68 71.676
R819 B.n142 B.n67 71.676
R820 B.n138 B.n66 71.676
R821 B.n134 B.n65 71.676
R822 B.n130 B.n64 71.676
R823 B.n126 B.n63 71.676
R824 B.n122 B.n62 71.676
R825 B.n118 B.n61 71.676
R826 B.n114 B.n60 71.676
R827 B.n110 B.n59 71.676
R828 B.n106 B.n58 71.676
R829 B.n102 B.n57 71.676
R830 B.n98 B.n56 71.676
R831 B.n452 B.n317 71.676
R832 B.n444 B.n285 71.676
R833 B.n440 B.n286 71.676
R834 B.n436 B.n287 71.676
R835 B.n432 B.n288 71.676
R836 B.n428 B.n289 71.676
R837 B.n424 B.n290 71.676
R838 B.n420 B.n291 71.676
R839 B.n416 B.n292 71.676
R840 B.n412 B.n293 71.676
R841 B.n408 B.n294 71.676
R842 B.n404 B.n295 71.676
R843 B.n400 B.n296 71.676
R844 B.n396 B.n297 71.676
R845 B.n392 B.n298 71.676
R846 B.n388 B.n299 71.676
R847 B.n384 B.n300 71.676
R848 B.n380 B.n301 71.676
R849 B.n375 B.n302 71.676
R850 B.n371 B.n303 71.676
R851 B.n367 B.n304 71.676
R852 B.n363 B.n305 71.676
R853 B.n359 B.n306 71.676
R854 B.n355 B.n307 71.676
R855 B.n351 B.n308 71.676
R856 B.n347 B.n309 71.676
R857 B.n343 B.n310 71.676
R858 B.n339 B.n311 71.676
R859 B.n335 B.n312 71.676
R860 B.n331 B.n313 71.676
R861 B.n327 B.n314 71.676
R862 B.n323 B.n315 71.676
R863 B.n455 B.n454 71.676
R864 B.n322 B.t9 70.4958
R865 B.n91 B.t20 70.4958
R866 B.n319 B.t12 70.4871
R867 B.n94 B.t17 70.4871
R868 B.n377 B.n322 59.5399
R869 B.n320 B.n319 59.5399
R870 B.n153 B.n94 59.5399
R871 B.n92 B.n91 59.5399
R872 B.n460 B.n281 58.2333
R873 B.n460 B.n277 58.2333
R874 B.n466 B.n277 58.2333
R875 B.n466 B.n273 58.2333
R876 B.n472 B.n273 58.2333
R877 B.n478 B.n269 58.2333
R878 B.n478 B.n265 58.2333
R879 B.n484 B.n265 58.2333
R880 B.n484 B.n260 58.2333
R881 B.n490 B.n260 58.2333
R882 B.n490 B.n261 58.2333
R883 B.n496 B.n252 58.2333
R884 B.n502 B.n252 58.2333
R885 B.n502 B.n253 58.2333
R886 B.n508 B.n245 58.2333
R887 B.n514 B.n245 58.2333
R888 B.n514 B.n241 58.2333
R889 B.n520 B.n241 58.2333
R890 B.n526 B.n237 58.2333
R891 B.n526 B.n233 58.2333
R892 B.n533 B.n233 58.2333
R893 B.n539 B.n229 58.2333
R894 B.n539 B.n4 58.2333
R895 B.n640 B.n4 58.2333
R896 B.n640 B.n639 58.2333
R897 B.n639 B.n638 58.2333
R898 B.n638 B.n8 58.2333
R899 B.n632 B.n631 58.2333
R900 B.n631 B.n630 58.2333
R901 B.n630 B.n15 58.2333
R902 B.n624 B.n623 58.2333
R903 B.n623 B.n622 58.2333
R904 B.n622 B.n22 58.2333
R905 B.n616 B.n22 58.2333
R906 B.n615 B.n614 58.2333
R907 B.n614 B.n29 58.2333
R908 B.n608 B.n29 58.2333
R909 B.n607 B.n606 58.2333
R910 B.n606 B.n36 58.2333
R911 B.n600 B.n36 58.2333
R912 B.n600 B.n599 58.2333
R913 B.n599 B.n598 58.2333
R914 B.n598 B.n43 58.2333
R915 B.n592 B.n591 58.2333
R916 B.n591 B.n590 58.2333
R917 B.n590 B.n50 58.2333
R918 B.n584 B.n50 58.2333
R919 B.n584 B.n583 58.2333
R920 B.t3 B.n237 55.6642
R921 B.t21 B.n15 55.6642
R922 B.t8 B.n269 50.526
R923 B.t15 B.n43 50.526
R924 B.n253 B.t0 47.1005
R925 B.t6 B.n615 47.1005
R926 B.t2 B.n229 41.9624
R927 B.t4 B.n8 41.9624
R928 B.n96 B.n52 34.1859
R929 B.n580 B.n579 34.1859
R930 B.n457 B.n456 34.1859
R931 B.n450 B.n279 34.1859
R932 B.n261 B.t5 33.3987
R933 B.t1 B.n607 33.3987
R934 B.n322 B.n321 27.9278
R935 B.n319 B.n318 27.9278
R936 B.n94 B.n93 27.9278
R937 B.n91 B.n90 27.9278
R938 B.n496 B.t5 24.8351
R939 B.n608 B.t1 24.8351
R940 B B.n642 18.0485
R941 B.n533 B.t2 16.2714
R942 B.n632 B.t4 16.2714
R943 B.n508 B.t0 11.1332
R944 B.n616 B.t6 11.1332
R945 B.n97 B.n96 10.6151
R946 B.n100 B.n97 10.6151
R947 B.n101 B.n100 10.6151
R948 B.n104 B.n101 10.6151
R949 B.n105 B.n104 10.6151
R950 B.n108 B.n105 10.6151
R951 B.n109 B.n108 10.6151
R952 B.n112 B.n109 10.6151
R953 B.n113 B.n112 10.6151
R954 B.n116 B.n113 10.6151
R955 B.n117 B.n116 10.6151
R956 B.n120 B.n117 10.6151
R957 B.n121 B.n120 10.6151
R958 B.n124 B.n121 10.6151
R959 B.n125 B.n124 10.6151
R960 B.n128 B.n125 10.6151
R961 B.n129 B.n128 10.6151
R962 B.n132 B.n129 10.6151
R963 B.n133 B.n132 10.6151
R964 B.n136 B.n133 10.6151
R965 B.n137 B.n136 10.6151
R966 B.n140 B.n137 10.6151
R967 B.n141 B.n140 10.6151
R968 B.n144 B.n141 10.6151
R969 B.n145 B.n144 10.6151
R970 B.n148 B.n145 10.6151
R971 B.n149 B.n148 10.6151
R972 B.n152 B.n149 10.6151
R973 B.n157 B.n154 10.6151
R974 B.n158 B.n157 10.6151
R975 B.n161 B.n158 10.6151
R976 B.n162 B.n161 10.6151
R977 B.n165 B.n162 10.6151
R978 B.n166 B.n165 10.6151
R979 B.n169 B.n166 10.6151
R980 B.n170 B.n169 10.6151
R981 B.n174 B.n173 10.6151
R982 B.n177 B.n174 10.6151
R983 B.n178 B.n177 10.6151
R984 B.n181 B.n178 10.6151
R985 B.n182 B.n181 10.6151
R986 B.n185 B.n182 10.6151
R987 B.n186 B.n185 10.6151
R988 B.n189 B.n186 10.6151
R989 B.n190 B.n189 10.6151
R990 B.n193 B.n190 10.6151
R991 B.n194 B.n193 10.6151
R992 B.n197 B.n194 10.6151
R993 B.n198 B.n197 10.6151
R994 B.n201 B.n198 10.6151
R995 B.n202 B.n201 10.6151
R996 B.n205 B.n202 10.6151
R997 B.n206 B.n205 10.6151
R998 B.n209 B.n206 10.6151
R999 B.n210 B.n209 10.6151
R1000 B.n213 B.n210 10.6151
R1001 B.n214 B.n213 10.6151
R1002 B.n217 B.n214 10.6151
R1003 B.n218 B.n217 10.6151
R1004 B.n221 B.n218 10.6151
R1005 B.n222 B.n221 10.6151
R1006 B.n225 B.n222 10.6151
R1007 B.n226 B.n225 10.6151
R1008 B.n580 B.n226 10.6151
R1009 B.n458 B.n457 10.6151
R1010 B.n458 B.n275 10.6151
R1011 B.n468 B.n275 10.6151
R1012 B.n469 B.n468 10.6151
R1013 B.n470 B.n469 10.6151
R1014 B.n470 B.n267 10.6151
R1015 B.n480 B.n267 10.6151
R1016 B.n481 B.n480 10.6151
R1017 B.n482 B.n481 10.6151
R1018 B.n482 B.n258 10.6151
R1019 B.n492 B.n258 10.6151
R1020 B.n493 B.n492 10.6151
R1021 B.n494 B.n493 10.6151
R1022 B.n494 B.n250 10.6151
R1023 B.n504 B.n250 10.6151
R1024 B.n505 B.n504 10.6151
R1025 B.n506 B.n505 10.6151
R1026 B.n506 B.n243 10.6151
R1027 B.n516 B.n243 10.6151
R1028 B.n517 B.n516 10.6151
R1029 B.n518 B.n517 10.6151
R1030 B.n518 B.n235 10.6151
R1031 B.n528 B.n235 10.6151
R1032 B.n529 B.n528 10.6151
R1033 B.n531 B.n529 10.6151
R1034 B.n531 B.n530 10.6151
R1035 B.n530 B.n227 10.6151
R1036 B.n542 B.n227 10.6151
R1037 B.n543 B.n542 10.6151
R1038 B.n544 B.n543 10.6151
R1039 B.n545 B.n544 10.6151
R1040 B.n547 B.n545 10.6151
R1041 B.n548 B.n547 10.6151
R1042 B.n549 B.n548 10.6151
R1043 B.n550 B.n549 10.6151
R1044 B.n552 B.n550 10.6151
R1045 B.n553 B.n552 10.6151
R1046 B.n554 B.n553 10.6151
R1047 B.n555 B.n554 10.6151
R1048 B.n557 B.n555 10.6151
R1049 B.n558 B.n557 10.6151
R1050 B.n559 B.n558 10.6151
R1051 B.n560 B.n559 10.6151
R1052 B.n562 B.n560 10.6151
R1053 B.n563 B.n562 10.6151
R1054 B.n564 B.n563 10.6151
R1055 B.n565 B.n564 10.6151
R1056 B.n567 B.n565 10.6151
R1057 B.n568 B.n567 10.6151
R1058 B.n569 B.n568 10.6151
R1059 B.n570 B.n569 10.6151
R1060 B.n572 B.n570 10.6151
R1061 B.n573 B.n572 10.6151
R1062 B.n574 B.n573 10.6151
R1063 B.n575 B.n574 10.6151
R1064 B.n577 B.n575 10.6151
R1065 B.n578 B.n577 10.6151
R1066 B.n579 B.n578 10.6151
R1067 B.n450 B.n449 10.6151
R1068 B.n449 B.n448 10.6151
R1069 B.n448 B.n447 10.6151
R1070 B.n447 B.n445 10.6151
R1071 B.n445 B.n442 10.6151
R1072 B.n442 B.n441 10.6151
R1073 B.n441 B.n438 10.6151
R1074 B.n438 B.n437 10.6151
R1075 B.n437 B.n434 10.6151
R1076 B.n434 B.n433 10.6151
R1077 B.n433 B.n430 10.6151
R1078 B.n430 B.n429 10.6151
R1079 B.n429 B.n426 10.6151
R1080 B.n426 B.n425 10.6151
R1081 B.n425 B.n422 10.6151
R1082 B.n422 B.n421 10.6151
R1083 B.n421 B.n418 10.6151
R1084 B.n418 B.n417 10.6151
R1085 B.n417 B.n414 10.6151
R1086 B.n414 B.n413 10.6151
R1087 B.n413 B.n410 10.6151
R1088 B.n410 B.n409 10.6151
R1089 B.n409 B.n406 10.6151
R1090 B.n406 B.n405 10.6151
R1091 B.n405 B.n402 10.6151
R1092 B.n402 B.n401 10.6151
R1093 B.n401 B.n398 10.6151
R1094 B.n398 B.n397 10.6151
R1095 B.n394 B.n393 10.6151
R1096 B.n393 B.n390 10.6151
R1097 B.n390 B.n389 10.6151
R1098 B.n389 B.n386 10.6151
R1099 B.n386 B.n385 10.6151
R1100 B.n385 B.n382 10.6151
R1101 B.n382 B.n381 10.6151
R1102 B.n381 B.n378 10.6151
R1103 B.n376 B.n373 10.6151
R1104 B.n373 B.n372 10.6151
R1105 B.n372 B.n369 10.6151
R1106 B.n369 B.n368 10.6151
R1107 B.n368 B.n365 10.6151
R1108 B.n365 B.n364 10.6151
R1109 B.n364 B.n361 10.6151
R1110 B.n361 B.n360 10.6151
R1111 B.n360 B.n357 10.6151
R1112 B.n357 B.n356 10.6151
R1113 B.n356 B.n353 10.6151
R1114 B.n353 B.n352 10.6151
R1115 B.n352 B.n349 10.6151
R1116 B.n349 B.n348 10.6151
R1117 B.n348 B.n345 10.6151
R1118 B.n345 B.n344 10.6151
R1119 B.n344 B.n341 10.6151
R1120 B.n341 B.n340 10.6151
R1121 B.n340 B.n337 10.6151
R1122 B.n337 B.n336 10.6151
R1123 B.n336 B.n333 10.6151
R1124 B.n333 B.n332 10.6151
R1125 B.n332 B.n329 10.6151
R1126 B.n329 B.n328 10.6151
R1127 B.n328 B.n325 10.6151
R1128 B.n325 B.n324 10.6151
R1129 B.n324 B.n283 10.6151
R1130 B.n456 B.n283 10.6151
R1131 B.n462 B.n279 10.6151
R1132 B.n463 B.n462 10.6151
R1133 B.n464 B.n463 10.6151
R1134 B.n464 B.n271 10.6151
R1135 B.n474 B.n271 10.6151
R1136 B.n475 B.n474 10.6151
R1137 B.n476 B.n475 10.6151
R1138 B.n476 B.n263 10.6151
R1139 B.n486 B.n263 10.6151
R1140 B.n487 B.n486 10.6151
R1141 B.n488 B.n487 10.6151
R1142 B.n488 B.n255 10.6151
R1143 B.n498 B.n255 10.6151
R1144 B.n499 B.n498 10.6151
R1145 B.n500 B.n499 10.6151
R1146 B.n500 B.n247 10.6151
R1147 B.n510 B.n247 10.6151
R1148 B.n511 B.n510 10.6151
R1149 B.n512 B.n511 10.6151
R1150 B.n512 B.n239 10.6151
R1151 B.n522 B.n239 10.6151
R1152 B.n523 B.n522 10.6151
R1153 B.n524 B.n523 10.6151
R1154 B.n524 B.n231 10.6151
R1155 B.n535 B.n231 10.6151
R1156 B.n536 B.n535 10.6151
R1157 B.n537 B.n536 10.6151
R1158 B.n537 B.n0 10.6151
R1159 B.n636 B.n1 10.6151
R1160 B.n636 B.n635 10.6151
R1161 B.n635 B.n634 10.6151
R1162 B.n634 B.n10 10.6151
R1163 B.n628 B.n10 10.6151
R1164 B.n628 B.n627 10.6151
R1165 B.n627 B.n626 10.6151
R1166 B.n626 B.n17 10.6151
R1167 B.n620 B.n17 10.6151
R1168 B.n620 B.n619 10.6151
R1169 B.n619 B.n618 10.6151
R1170 B.n618 B.n24 10.6151
R1171 B.n612 B.n24 10.6151
R1172 B.n612 B.n611 10.6151
R1173 B.n611 B.n610 10.6151
R1174 B.n610 B.n31 10.6151
R1175 B.n604 B.n31 10.6151
R1176 B.n604 B.n603 10.6151
R1177 B.n603 B.n602 10.6151
R1178 B.n602 B.n38 10.6151
R1179 B.n596 B.n38 10.6151
R1180 B.n596 B.n595 10.6151
R1181 B.n595 B.n594 10.6151
R1182 B.n594 B.n45 10.6151
R1183 B.n588 B.n45 10.6151
R1184 B.n588 B.n587 10.6151
R1185 B.n587 B.n586 10.6151
R1186 B.n586 B.n52 10.6151
R1187 B.n472 B.t8 7.70778
R1188 B.n592 B.t15 7.70778
R1189 B.n154 B.n153 6.5566
R1190 B.n170 B.n92 6.5566
R1191 B.n394 B.n320 6.5566
R1192 B.n378 B.n377 6.5566
R1193 B.n153 B.n152 4.05904
R1194 B.n173 B.n92 4.05904
R1195 B.n397 B.n320 4.05904
R1196 B.n377 B.n376 4.05904
R1197 B.n642 B.n0 2.81026
R1198 B.n642 B.n1 2.81026
R1199 B.n520 B.t3 2.56959
R1200 B.n624 B.t21 2.56959
R1201 VN.n3 VN.t6 222.696
R1202 VN.n16 VN.t2 222.696
R1203 VN.n11 VN.t5 199.965
R1204 VN.n24 VN.t7 199.965
R1205 VN.n4 VN.t1 164.358
R1206 VN.n1 VN.t0 164.358
R1207 VN.n17 VN.t3 164.358
R1208 VN.n14 VN.t4 164.358
R1209 VN.n23 VN.n13 161.3
R1210 VN.n22 VN.n21 161.3
R1211 VN.n20 VN.n19 161.3
R1212 VN.n18 VN.n15 161.3
R1213 VN.n10 VN.n0 161.3
R1214 VN.n9 VN.n8 161.3
R1215 VN.n7 VN.n6 161.3
R1216 VN.n5 VN.n2 161.3
R1217 VN.n25 VN.n24 80.6037
R1218 VN.n12 VN.n11 80.6037
R1219 VN.n6 VN.n5 56.5193
R1220 VN.n19 VN.n18 56.5193
R1221 VN.n11 VN.n10 49.4239
R1222 VN.n24 VN.n23 49.4239
R1223 VN VN.n25 41.0294
R1224 VN.n4 VN.n3 33.8527
R1225 VN.n17 VN.n16 33.8527
R1226 VN.n16 VN.n15 28.2774
R1227 VN.n3 VN.n2 28.2774
R1228 VN.n10 VN.n9 24.4675
R1229 VN.n23 VN.n22 24.4675
R1230 VN.n5 VN.n4 22.9995
R1231 VN.n6 VN.n1 22.9995
R1232 VN.n18 VN.n17 22.9995
R1233 VN.n19 VN.n14 22.9995
R1234 VN.n9 VN.n1 1.46852
R1235 VN.n22 VN.n14 1.46852
R1236 VN.n25 VN.n13 0.285035
R1237 VN.n12 VN.n0 0.285035
R1238 VN.n21 VN.n13 0.189894
R1239 VN.n21 VN.n20 0.189894
R1240 VN.n20 VN.n15 0.189894
R1241 VN.n7 VN.n2 0.189894
R1242 VN.n8 VN.n7 0.189894
R1243 VN.n8 VN.n0 0.189894
R1244 VN VN.n12 0.146778
R1245 VDD2.n2 VDD2.n1 67.3776
R1246 VDD2.n2 VDD2.n0 67.3776
R1247 VDD2 VDD2.n5 67.3748
R1248 VDD2.n4 VDD2.n3 66.8125
R1249 VDD2.n4 VDD2.n2 35.8274
R1250 VDD2.n5 VDD2.t4 2.61609
R1251 VDD2.n5 VDD2.t5 2.61609
R1252 VDD2.n3 VDD2.t0 2.61609
R1253 VDD2.n3 VDD2.t3 2.61609
R1254 VDD2.n1 VDD2.t7 2.61609
R1255 VDD2.n1 VDD2.t2 2.61609
R1256 VDD2.n0 VDD2.t1 2.61609
R1257 VDD2.n0 VDD2.t6 2.61609
R1258 VDD2 VDD2.n4 0.679379
C0 VDD1 VN 0.14909f
C1 VDD1 VP 4.64181f
C2 VN VTAIL 4.51757f
C3 VN VDD2 4.43037f
C4 VTAIL VP 4.53167f
C5 VDD2 VP 0.361175f
C6 VDD1 VTAIL 6.75084f
C7 VDD1 VDD2 1.03155f
C8 VDD2 VTAIL 6.79527f
C9 VN VP 5.01906f
C10 VDD2 B 3.533987f
C11 VDD1 B 3.813775f
C12 VTAIL B 6.782642f
C13 VN B 9.5317f
C14 VP B 7.951651f
C15 VDD2.t1 B 0.152046f
C16 VDD2.t6 B 0.152046f
C17 VDD2.n0 B 1.31396f
C18 VDD2.t7 B 0.152046f
C19 VDD2.t2 B 0.152046f
C20 VDD2.n1 B 1.31396f
C21 VDD2.n2 B 2.16155f
C22 VDD2.t0 B 0.152046f
C23 VDD2.t3 B 0.152046f
C24 VDD2.n3 B 1.31095f
C25 VDD2.n4 B 2.11216f
C26 VDD2.t4 B 0.152046f
C27 VDD2.t5 B 0.152046f
C28 VDD2.n5 B 1.31394f
C29 VN.n0 B 0.049183f
C30 VN.t0 B 0.829738f
C31 VN.n1 B 0.323234f
C32 VN.n2 B 0.19226f
C33 VN.t1 B 0.829738f
C34 VN.t6 B 0.932802f
C35 VN.n3 B 0.372196f
C36 VN.n4 B 0.381392f
C37 VN.n5 B 0.051772f
C38 VN.n6 B 0.051772f
C39 VN.n7 B 0.036859f
C40 VN.n8 B 0.036859f
C41 VN.n9 B 0.036815f
C42 VN.n10 B 0.04544f
C43 VN.t5 B 0.892417f
C44 VN.n11 B 0.386679f
C45 VN.n12 B 0.03452f
C46 VN.n13 B 0.049183f
C47 VN.t4 B 0.829738f
C48 VN.n14 B 0.323234f
C49 VN.n15 B 0.19226f
C50 VN.t3 B 0.829738f
C51 VN.t2 B 0.932802f
C52 VN.n16 B 0.372196f
C53 VN.n17 B 0.381392f
C54 VN.n18 B 0.051772f
C55 VN.n19 B 0.051772f
C56 VN.n20 B 0.036859f
C57 VN.n21 B 0.036859f
C58 VN.n22 B 0.036815f
C59 VN.n23 B 0.04544f
C60 VN.t7 B 0.892417f
C61 VN.n24 B 0.386679f
C62 VN.n25 B 1.47947f
C63 VDD1.t1 B 0.153474f
C64 VDD1.t2 B 0.153474f
C65 VDD1.n0 B 1.327f
C66 VDD1.t5 B 0.153474f
C67 VDD1.t7 B 0.153474f
C68 VDD1.n1 B 1.32631f
C69 VDD1.t6 B 0.153474f
C70 VDD1.t4 B 0.153474f
C71 VDD1.n2 B 1.32631f
C72 VDD1.n3 B 2.23647f
C73 VDD1.t0 B 0.153474f
C74 VDD1.t3 B 0.153474f
C75 VDD1.n4 B 1.32326f
C76 VDD1.n5 B 2.16254f
C77 VTAIL.t15 B 0.122888f
C78 VTAIL.t6 B 0.122888f
C79 VTAIL.n0 B 1.00694f
C80 VTAIL.n1 B 0.272728f
C81 VTAIL.t4 B 1.28164f
C82 VTAIL.n2 B 0.360432f
C83 VTAIL.t12 B 1.28164f
C84 VTAIL.n3 B 0.360432f
C85 VTAIL.t10 B 0.122888f
C86 VTAIL.t11 B 0.122888f
C87 VTAIL.n4 B 1.00694f
C88 VTAIL.n5 B 0.351048f
C89 VTAIL.t14 B 1.28164f
C90 VTAIL.n6 B 1.12252f
C91 VTAIL.t5 B 1.28164f
C92 VTAIL.n7 B 1.12252f
C93 VTAIL.t0 B 0.122888f
C94 VTAIL.t3 B 0.122888f
C95 VTAIL.n8 B 1.00695f
C96 VTAIL.n9 B 0.351045f
C97 VTAIL.t2 B 1.28164f
C98 VTAIL.n10 B 0.360429f
C99 VTAIL.t7 B 1.28164f
C100 VTAIL.n11 B 0.360429f
C101 VTAIL.t13 B 0.122888f
C102 VTAIL.t8 B 0.122888f
C103 VTAIL.n12 B 1.00695f
C104 VTAIL.n13 B 0.351045f
C105 VTAIL.t9 B 1.28164f
C106 VTAIL.n14 B 1.12252f
C107 VTAIL.t1 B 1.28164f
C108 VTAIL.n15 B 1.11867f
C109 VP.n0 B 0.050077f
C110 VP.t1 B 0.844826f
C111 VP.n1 B 0.329112f
C112 VP.n2 B 0.037529f
C113 VP.t0 B 0.844826f
C114 VP.n3 B 0.046266f
C115 VP.n4 B 0.050077f
C116 VP.t4 B 0.908645f
C117 VP.t7 B 0.844826f
C118 VP.n5 B 0.329112f
C119 VP.n6 B 0.195756f
C120 VP.t5 B 0.844826f
C121 VP.t6 B 0.949764f
C122 VP.n7 B 0.378964f
C123 VP.n8 B 0.388327f
C124 VP.n9 B 0.052713f
C125 VP.n10 B 0.052713f
C126 VP.n11 B 0.037529f
C127 VP.n12 B 0.037529f
C128 VP.n13 B 0.037484f
C129 VP.n14 B 0.046266f
C130 VP.n15 B 0.393711f
C131 VP.n16 B 1.4852f
C132 VP.t2 B 0.908645f
C133 VP.n17 B 0.393711f
C134 VP.n18 B 1.51831f
C135 VP.n19 B 0.050077f
C136 VP.n20 B 0.037529f
C137 VP.n21 B 0.037484f
C138 VP.n22 B 0.329112f
C139 VP.n23 B 0.052713f
C140 VP.n24 B 0.052713f
C141 VP.n25 B 0.037529f
C142 VP.n26 B 0.037529f
C143 VP.n27 B 0.037484f
C144 VP.n28 B 0.046266f
C145 VP.t3 B 0.908645f
C146 VP.n29 B 0.393711f
C147 VP.n30 B 0.035147f
.ends

