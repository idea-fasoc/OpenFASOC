* NGSPICE file created from diff_pair_sample_1477.ext - technology: sky130A

.subckt diff_pair_sample_1477 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.3627 ps=2.64 w=0.93 l=1.32
X1 VDD2.t7 VN.t0 VTAIL.t7 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.3627 ps=2.64 w=0.93 l=1.32
X2 VTAIL.t11 VP.t1 VDD1.t6 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0.15345 ps=1.26 w=0.93 l=1.32
X3 VTAIL.t15 VP.t2 VDD1.t5 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0.15345 ps=1.26 w=0.93 l=1.32
X4 B.t11 B.t9 B.t10 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0 ps=0 w=0.93 l=1.32
X5 VDD2.t6 VN.t1 VTAIL.t1 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X6 VDD1.t4 VP.t3 VTAIL.t8 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.3627 ps=2.64 w=0.93 l=1.32
X7 VDD2.t5 VN.t2 VTAIL.t4 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X8 VDD2.t4 VN.t3 VTAIL.t2 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.3627 ps=2.64 w=0.93 l=1.32
X9 VDD1.t3 VP.t4 VTAIL.t12 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X10 B.t8 B.t6 B.t7 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0 ps=0 w=0.93 l=1.32
X11 B.t5 B.t3 B.t4 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0 ps=0 w=0.93 l=1.32
X12 VTAIL.t9 VP.t5 VDD1.t2 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X13 VTAIL.t3 VN.t4 VDD2.t3 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X14 VTAIL.t10 VP.t6 VDD1.t1 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X15 VTAIL.t5 VN.t5 VDD2.t2 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X16 VTAIL.t0 VN.t6 VDD2.t1 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0.15345 ps=1.26 w=0.93 l=1.32
X17 VDD1.t0 VP.t7 VTAIL.t14 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.15345 pd=1.26 as=0.15345 ps=1.26 w=0.93 l=1.32
X18 VTAIL.t6 VN.t7 VDD2.t0 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0.15345 ps=1.26 w=0.93 l=1.32
X19 B.t2 B.t0 B.t1 w_n2620_n1154# sky130_fd_pr__pfet_01v8 ad=0.3627 pd=2.64 as=0 ps=0 w=0.93 l=1.32
R0 VP.n25 VP.n5 174.757
R1 VP.n44 VP.n43 174.757
R2 VP.n24 VP.n23 174.757
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n42 VP.n0 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n39 VP.n1 161.3
R13 VP.n38 VP.n37 161.3
R14 VP.n35 VP.n2 161.3
R15 VP.n34 VP.n33 161.3
R16 VP.n32 VP.n3 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n28 VP.n4 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n11 VP.n10 61.745
R21 VP.n35 VP.n34 56.5193
R22 VP.n15 VP.n14 56.5193
R23 VP.n30 VP.n28 50.2061
R24 VP.n41 VP.n1 50.2061
R25 VP.n21 VP.n7 50.2061
R26 VP.n11 VP.t2 45.0385
R27 VP.n25 VP.n24 36.4172
R28 VP.n28 VP.n27 30.7807
R29 VP.n42 VP.n41 30.7807
R30 VP.n22 VP.n21 30.7807
R31 VP.n12 VP.n11 27.4982
R32 VP.n34 VP.n3 24.4675
R33 VP.n37 VP.n35 24.4675
R34 VP.n17 VP.n15 24.4675
R35 VP.n14 VP.n9 24.4675
R36 VP.n30 VP.n29 20.7975
R37 VP.n36 VP.n1 20.7975
R38 VP.n16 VP.n7 20.7975
R39 VP.n5 VP.t1 16.98
R40 VP.n29 VP.t7 16.98
R41 VP.n36 VP.t5 16.98
R42 VP.n43 VP.t3 16.98
R43 VP.n23 VP.t0 16.98
R44 VP.n16 VP.t6 16.98
R45 VP.n10 VP.t4 16.98
R46 VP.n27 VP.n5 11.0107
R47 VP.n43 VP.n42 11.0107
R48 VP.n23 VP.n22 11.0107
R49 VP.n29 VP.n3 3.67055
R50 VP.n37 VP.n36 3.67055
R51 VP.n17 VP.n16 3.67055
R52 VP.n10 VP.n9 3.67055
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VTAIL.n14 VTAIL.t13 657.048
R73 VTAIL.n11 VTAIL.t15 657.048
R74 VTAIL.n10 VTAIL.t2 657.048
R75 VTAIL.n7 VTAIL.t0 657.048
R76 VTAIL.n15 VTAIL.t7 657.048
R77 VTAIL.n2 VTAIL.t6 657.048
R78 VTAIL.n3 VTAIL.t8 657.048
R79 VTAIL.n6 VTAIL.t11 657.048
R80 VTAIL.n13 VTAIL.n12 622.096
R81 VTAIL.n9 VTAIL.n8 622.096
R82 VTAIL.n1 VTAIL.n0 622.096
R83 VTAIL.n5 VTAIL.n4 622.096
R84 VTAIL.n0 VTAIL.t1 34.9521
R85 VTAIL.n0 VTAIL.t3 34.9521
R86 VTAIL.n4 VTAIL.t14 34.9521
R87 VTAIL.n4 VTAIL.t9 34.9521
R88 VTAIL.n12 VTAIL.t12 34.9521
R89 VTAIL.n12 VTAIL.t10 34.9521
R90 VTAIL.n8 VTAIL.t4 34.9521
R91 VTAIL.n8 VTAIL.t5 34.9521
R92 VTAIL.n15 VTAIL.n14 14.591
R93 VTAIL.n7 VTAIL.n6 14.591
R94 VTAIL.n9 VTAIL.n7 1.42291
R95 VTAIL.n10 VTAIL.n9 1.42291
R96 VTAIL.n13 VTAIL.n11 1.42291
R97 VTAIL.n14 VTAIL.n13 1.42291
R98 VTAIL.n6 VTAIL.n5 1.42291
R99 VTAIL.n5 VTAIL.n3 1.42291
R100 VTAIL.n2 VTAIL.n1 1.42291
R101 VTAIL VTAIL.n15 1.36472
R102 VTAIL.n11 VTAIL.n10 0.470328
R103 VTAIL.n3 VTAIL.n2 0.470328
R104 VTAIL VTAIL.n1 0.0586897
R105 VDD1 VDD1.n0 639.544
R106 VDD1.n3 VDD1.n2 639.431
R107 VDD1.n3 VDD1.n1 639.431
R108 VDD1.n5 VDD1.n4 638.775
R109 VDD1.n4 VDD1.t1 34.9521
R110 VDD1.n4 VDD1.t7 34.9521
R111 VDD1.n0 VDD1.t5 34.9521
R112 VDD1.n0 VDD1.t3 34.9521
R113 VDD1.n2 VDD1.t2 34.9521
R114 VDD1.n2 VDD1.t4 34.9521
R115 VDD1.n1 VDD1.t6 34.9521
R116 VDD1.n1 VDD1.t0 34.9521
R117 VDD1.n5 VDD1.n3 31.5009
R118 VDD1 VDD1.n5 0.653517
R119 VN.n18 VN.n17 174.757
R120 VN.n37 VN.n36 174.757
R121 VN.n35 VN.n19 161.3
R122 VN.n34 VN.n33 161.3
R123 VN.n32 VN.n20 161.3
R124 VN.n31 VN.n30 161.3
R125 VN.n29 VN.n21 161.3
R126 VN.n28 VN.n27 161.3
R127 VN.n26 VN.n23 161.3
R128 VN.n16 VN.n0 161.3
R129 VN.n15 VN.n14 161.3
R130 VN.n13 VN.n1 161.3
R131 VN.n12 VN.n11 161.3
R132 VN.n9 VN.n2 161.3
R133 VN.n8 VN.n7 161.3
R134 VN.n6 VN.n3 161.3
R135 VN.n5 VN.n4 61.745
R136 VN.n25 VN.n24 61.745
R137 VN.n9 VN.n8 56.5193
R138 VN.n29 VN.n28 56.5193
R139 VN.n15 VN.n1 50.2061
R140 VN.n34 VN.n20 50.2061
R141 VN.n5 VN.t7 45.0385
R142 VN.n25 VN.t3 45.0385
R143 VN VN.n37 36.7978
R144 VN.n16 VN.n15 30.7807
R145 VN.n35 VN.n34 30.7807
R146 VN.n26 VN.n25 27.4982
R147 VN.n6 VN.n5 27.4982
R148 VN.n8 VN.n3 24.4675
R149 VN.n11 VN.n9 24.4675
R150 VN.n28 VN.n23 24.4675
R151 VN.n30 VN.n29 24.4675
R152 VN.n10 VN.n1 20.7975
R153 VN.n22 VN.n20 20.7975
R154 VN.n4 VN.t1 16.98
R155 VN.n10 VN.t4 16.98
R156 VN.n17 VN.t0 16.98
R157 VN.n24 VN.t5 16.98
R158 VN.n22 VN.t2 16.98
R159 VN.n36 VN.t6 16.98
R160 VN.n17 VN.n16 11.0107
R161 VN.n36 VN.n35 11.0107
R162 VN.n4 VN.n3 3.67055
R163 VN.n11 VN.n10 3.67055
R164 VN.n24 VN.n23 3.67055
R165 VN.n30 VN.n22 3.67055
R166 VN.n37 VN.n19 0.189894
R167 VN.n33 VN.n19 0.189894
R168 VN.n33 VN.n32 0.189894
R169 VN.n32 VN.n31 0.189894
R170 VN.n31 VN.n21 0.189894
R171 VN.n27 VN.n21 0.189894
R172 VN.n27 VN.n26 0.189894
R173 VN.n7 VN.n6 0.189894
R174 VN.n7 VN.n2 0.189894
R175 VN.n12 VN.n2 0.189894
R176 VN.n13 VN.n12 0.189894
R177 VN.n14 VN.n13 0.189894
R178 VN.n14 VN.n0 0.189894
R179 VN.n18 VN.n0 0.189894
R180 VN VN.n18 0.0516364
R181 VDD2.n2 VDD2.n1 639.431
R182 VDD2.n2 VDD2.n0 639.431
R183 VDD2 VDD2.n5 639.428
R184 VDD2.n4 VDD2.n3 638.775
R185 VDD2.n5 VDD2.t2 34.9521
R186 VDD2.n5 VDD2.t4 34.9521
R187 VDD2.n3 VDD2.t1 34.9521
R188 VDD2.n3 VDD2.t5 34.9521
R189 VDD2.n1 VDD2.t3 34.9521
R190 VDD2.n1 VDD2.t7 34.9521
R191 VDD2.n0 VDD2.t0 34.9521
R192 VDD2.n0 VDD2.t6 34.9521
R193 VDD2.n4 VDD2.n2 30.9179
R194 VDD2 VDD2.n4 0.769897
R195 B.n160 B.t10 679.88
R196 B.n75 B.t4 679.88
R197 B.n31 B.t2 679.88
R198 B.n24 B.t8 679.88
R199 B.n161 B.t11 647.88
R200 B.n76 B.t5 647.88
R201 B.n32 B.t1 647.88
R202 B.n25 B.t7 647.88
R203 B.n193 B.n70 585
R204 B.n192 B.n191 585
R205 B.n190 B.n71 585
R206 B.n189 B.n188 585
R207 B.n187 B.n72 585
R208 B.n186 B.n185 585
R209 B.n184 B.n73 585
R210 B.n183 B.n182 585
R211 B.n181 B.n74 585
R212 B.n179 B.n178 585
R213 B.n177 B.n77 585
R214 B.n176 B.n175 585
R215 B.n174 B.n78 585
R216 B.n173 B.n172 585
R217 B.n171 B.n79 585
R218 B.n170 B.n169 585
R219 B.n168 B.n80 585
R220 B.n167 B.n166 585
R221 B.n165 B.n81 585
R222 B.n164 B.n163 585
R223 B.n159 B.n82 585
R224 B.n158 B.n157 585
R225 B.n156 B.n83 585
R226 B.n155 B.n154 585
R227 B.n153 B.n84 585
R228 B.n152 B.n151 585
R229 B.n150 B.n85 585
R230 B.n149 B.n148 585
R231 B.n195 B.n194 585
R232 B.n196 B.n69 585
R233 B.n198 B.n197 585
R234 B.n199 B.n68 585
R235 B.n201 B.n200 585
R236 B.n202 B.n67 585
R237 B.n204 B.n203 585
R238 B.n205 B.n66 585
R239 B.n207 B.n206 585
R240 B.n208 B.n65 585
R241 B.n210 B.n209 585
R242 B.n211 B.n64 585
R243 B.n213 B.n212 585
R244 B.n214 B.n63 585
R245 B.n216 B.n215 585
R246 B.n217 B.n62 585
R247 B.n219 B.n218 585
R248 B.n220 B.n61 585
R249 B.n222 B.n221 585
R250 B.n223 B.n60 585
R251 B.n225 B.n224 585
R252 B.n226 B.n59 585
R253 B.n228 B.n227 585
R254 B.n229 B.n58 585
R255 B.n231 B.n230 585
R256 B.n232 B.n57 585
R257 B.n234 B.n233 585
R258 B.n235 B.n56 585
R259 B.n237 B.n236 585
R260 B.n238 B.n55 585
R261 B.n240 B.n239 585
R262 B.n241 B.n54 585
R263 B.n243 B.n242 585
R264 B.n244 B.n53 585
R265 B.n246 B.n245 585
R266 B.n247 B.n52 585
R267 B.n249 B.n248 585
R268 B.n250 B.n51 585
R269 B.n252 B.n251 585
R270 B.n253 B.n50 585
R271 B.n255 B.n254 585
R272 B.n256 B.n49 585
R273 B.n258 B.n257 585
R274 B.n259 B.n48 585
R275 B.n261 B.n260 585
R276 B.n262 B.n47 585
R277 B.n264 B.n263 585
R278 B.n265 B.n46 585
R279 B.n267 B.n266 585
R280 B.n268 B.n45 585
R281 B.n270 B.n269 585
R282 B.n271 B.n44 585
R283 B.n273 B.n272 585
R284 B.n274 B.n43 585
R285 B.n276 B.n275 585
R286 B.n277 B.n42 585
R287 B.n279 B.n278 585
R288 B.n280 B.n41 585
R289 B.n282 B.n281 585
R290 B.n283 B.n40 585
R291 B.n285 B.n284 585
R292 B.n286 B.n39 585
R293 B.n288 B.n287 585
R294 B.n289 B.n38 585
R295 B.n291 B.n290 585
R296 B.n292 B.n37 585
R297 B.n335 B.n18 585
R298 B.n334 B.n333 585
R299 B.n332 B.n19 585
R300 B.n331 B.n330 585
R301 B.n329 B.n20 585
R302 B.n328 B.n327 585
R303 B.n326 B.n21 585
R304 B.n325 B.n324 585
R305 B.n323 B.n22 585
R306 B.n322 B.n321 585
R307 B.n320 B.n23 585
R308 B.n319 B.n318 585
R309 B.n317 B.n27 585
R310 B.n316 B.n315 585
R311 B.n314 B.n28 585
R312 B.n313 B.n312 585
R313 B.n311 B.n29 585
R314 B.n310 B.n309 585
R315 B.n308 B.n30 585
R316 B.n306 B.n305 585
R317 B.n304 B.n33 585
R318 B.n303 B.n302 585
R319 B.n301 B.n34 585
R320 B.n300 B.n299 585
R321 B.n298 B.n35 585
R322 B.n297 B.n296 585
R323 B.n295 B.n36 585
R324 B.n294 B.n293 585
R325 B.n337 B.n336 585
R326 B.n338 B.n17 585
R327 B.n340 B.n339 585
R328 B.n341 B.n16 585
R329 B.n343 B.n342 585
R330 B.n344 B.n15 585
R331 B.n346 B.n345 585
R332 B.n347 B.n14 585
R333 B.n349 B.n348 585
R334 B.n350 B.n13 585
R335 B.n352 B.n351 585
R336 B.n353 B.n12 585
R337 B.n355 B.n354 585
R338 B.n356 B.n11 585
R339 B.n358 B.n357 585
R340 B.n359 B.n10 585
R341 B.n361 B.n360 585
R342 B.n362 B.n9 585
R343 B.n364 B.n363 585
R344 B.n365 B.n8 585
R345 B.n367 B.n366 585
R346 B.n368 B.n7 585
R347 B.n370 B.n369 585
R348 B.n371 B.n6 585
R349 B.n373 B.n372 585
R350 B.n374 B.n5 585
R351 B.n376 B.n375 585
R352 B.n377 B.n4 585
R353 B.n379 B.n378 585
R354 B.n380 B.n3 585
R355 B.n382 B.n381 585
R356 B.n383 B.n0 585
R357 B.n2 B.n1 585
R358 B.n102 B.n101 585
R359 B.n104 B.n103 585
R360 B.n105 B.n100 585
R361 B.n107 B.n106 585
R362 B.n108 B.n99 585
R363 B.n110 B.n109 585
R364 B.n111 B.n98 585
R365 B.n113 B.n112 585
R366 B.n114 B.n97 585
R367 B.n116 B.n115 585
R368 B.n117 B.n96 585
R369 B.n119 B.n118 585
R370 B.n120 B.n95 585
R371 B.n122 B.n121 585
R372 B.n123 B.n94 585
R373 B.n125 B.n124 585
R374 B.n126 B.n93 585
R375 B.n128 B.n127 585
R376 B.n129 B.n92 585
R377 B.n131 B.n130 585
R378 B.n132 B.n91 585
R379 B.n134 B.n133 585
R380 B.n135 B.n90 585
R381 B.n137 B.n136 585
R382 B.n138 B.n89 585
R383 B.n140 B.n139 585
R384 B.n141 B.n88 585
R385 B.n143 B.n142 585
R386 B.n144 B.n87 585
R387 B.n146 B.n145 585
R388 B.n147 B.n86 585
R389 B.n149 B.n86 454.062
R390 B.n195 B.n70 454.062
R391 B.n293 B.n292 454.062
R392 B.n336 B.n335 454.062
R393 B.n385 B.n384 256.663
R394 B.n384 B.n383 235.042
R395 B.n384 B.n2 235.042
R396 B.n75 B.t3 222.321
R397 B.n31 B.t0 222.321
R398 B.n160 B.t9 221.817
R399 B.n24 B.t6 221.817
R400 B.n150 B.n149 163.367
R401 B.n151 B.n150 163.367
R402 B.n151 B.n84 163.367
R403 B.n155 B.n84 163.367
R404 B.n156 B.n155 163.367
R405 B.n157 B.n156 163.367
R406 B.n157 B.n82 163.367
R407 B.n164 B.n82 163.367
R408 B.n165 B.n164 163.367
R409 B.n166 B.n165 163.367
R410 B.n166 B.n80 163.367
R411 B.n170 B.n80 163.367
R412 B.n171 B.n170 163.367
R413 B.n172 B.n171 163.367
R414 B.n172 B.n78 163.367
R415 B.n176 B.n78 163.367
R416 B.n177 B.n176 163.367
R417 B.n178 B.n177 163.367
R418 B.n178 B.n74 163.367
R419 B.n183 B.n74 163.367
R420 B.n184 B.n183 163.367
R421 B.n185 B.n184 163.367
R422 B.n185 B.n72 163.367
R423 B.n189 B.n72 163.367
R424 B.n190 B.n189 163.367
R425 B.n191 B.n190 163.367
R426 B.n191 B.n70 163.367
R427 B.n292 B.n291 163.367
R428 B.n291 B.n38 163.367
R429 B.n287 B.n38 163.367
R430 B.n287 B.n286 163.367
R431 B.n286 B.n285 163.367
R432 B.n285 B.n40 163.367
R433 B.n281 B.n40 163.367
R434 B.n281 B.n280 163.367
R435 B.n280 B.n279 163.367
R436 B.n279 B.n42 163.367
R437 B.n275 B.n42 163.367
R438 B.n275 B.n274 163.367
R439 B.n274 B.n273 163.367
R440 B.n273 B.n44 163.367
R441 B.n269 B.n44 163.367
R442 B.n269 B.n268 163.367
R443 B.n268 B.n267 163.367
R444 B.n267 B.n46 163.367
R445 B.n263 B.n46 163.367
R446 B.n263 B.n262 163.367
R447 B.n262 B.n261 163.367
R448 B.n261 B.n48 163.367
R449 B.n257 B.n48 163.367
R450 B.n257 B.n256 163.367
R451 B.n256 B.n255 163.367
R452 B.n255 B.n50 163.367
R453 B.n251 B.n50 163.367
R454 B.n251 B.n250 163.367
R455 B.n250 B.n249 163.367
R456 B.n249 B.n52 163.367
R457 B.n245 B.n52 163.367
R458 B.n245 B.n244 163.367
R459 B.n244 B.n243 163.367
R460 B.n243 B.n54 163.367
R461 B.n239 B.n54 163.367
R462 B.n239 B.n238 163.367
R463 B.n238 B.n237 163.367
R464 B.n237 B.n56 163.367
R465 B.n233 B.n56 163.367
R466 B.n233 B.n232 163.367
R467 B.n232 B.n231 163.367
R468 B.n231 B.n58 163.367
R469 B.n227 B.n58 163.367
R470 B.n227 B.n226 163.367
R471 B.n226 B.n225 163.367
R472 B.n225 B.n60 163.367
R473 B.n221 B.n60 163.367
R474 B.n221 B.n220 163.367
R475 B.n220 B.n219 163.367
R476 B.n219 B.n62 163.367
R477 B.n215 B.n62 163.367
R478 B.n215 B.n214 163.367
R479 B.n214 B.n213 163.367
R480 B.n213 B.n64 163.367
R481 B.n209 B.n64 163.367
R482 B.n209 B.n208 163.367
R483 B.n208 B.n207 163.367
R484 B.n207 B.n66 163.367
R485 B.n203 B.n66 163.367
R486 B.n203 B.n202 163.367
R487 B.n202 B.n201 163.367
R488 B.n201 B.n68 163.367
R489 B.n197 B.n68 163.367
R490 B.n197 B.n196 163.367
R491 B.n196 B.n195 163.367
R492 B.n335 B.n334 163.367
R493 B.n334 B.n19 163.367
R494 B.n330 B.n19 163.367
R495 B.n330 B.n329 163.367
R496 B.n329 B.n328 163.367
R497 B.n328 B.n21 163.367
R498 B.n324 B.n21 163.367
R499 B.n324 B.n323 163.367
R500 B.n323 B.n322 163.367
R501 B.n322 B.n23 163.367
R502 B.n318 B.n23 163.367
R503 B.n318 B.n317 163.367
R504 B.n317 B.n316 163.367
R505 B.n316 B.n28 163.367
R506 B.n312 B.n28 163.367
R507 B.n312 B.n311 163.367
R508 B.n311 B.n310 163.367
R509 B.n310 B.n30 163.367
R510 B.n305 B.n30 163.367
R511 B.n305 B.n304 163.367
R512 B.n304 B.n303 163.367
R513 B.n303 B.n34 163.367
R514 B.n299 B.n34 163.367
R515 B.n299 B.n298 163.367
R516 B.n298 B.n297 163.367
R517 B.n297 B.n36 163.367
R518 B.n293 B.n36 163.367
R519 B.n336 B.n17 163.367
R520 B.n340 B.n17 163.367
R521 B.n341 B.n340 163.367
R522 B.n342 B.n341 163.367
R523 B.n342 B.n15 163.367
R524 B.n346 B.n15 163.367
R525 B.n347 B.n346 163.367
R526 B.n348 B.n347 163.367
R527 B.n348 B.n13 163.367
R528 B.n352 B.n13 163.367
R529 B.n353 B.n352 163.367
R530 B.n354 B.n353 163.367
R531 B.n354 B.n11 163.367
R532 B.n358 B.n11 163.367
R533 B.n359 B.n358 163.367
R534 B.n360 B.n359 163.367
R535 B.n360 B.n9 163.367
R536 B.n364 B.n9 163.367
R537 B.n365 B.n364 163.367
R538 B.n366 B.n365 163.367
R539 B.n366 B.n7 163.367
R540 B.n370 B.n7 163.367
R541 B.n371 B.n370 163.367
R542 B.n372 B.n371 163.367
R543 B.n372 B.n5 163.367
R544 B.n376 B.n5 163.367
R545 B.n377 B.n376 163.367
R546 B.n378 B.n377 163.367
R547 B.n378 B.n3 163.367
R548 B.n382 B.n3 163.367
R549 B.n383 B.n382 163.367
R550 B.n102 B.n2 163.367
R551 B.n103 B.n102 163.367
R552 B.n103 B.n100 163.367
R553 B.n107 B.n100 163.367
R554 B.n108 B.n107 163.367
R555 B.n109 B.n108 163.367
R556 B.n109 B.n98 163.367
R557 B.n113 B.n98 163.367
R558 B.n114 B.n113 163.367
R559 B.n115 B.n114 163.367
R560 B.n115 B.n96 163.367
R561 B.n119 B.n96 163.367
R562 B.n120 B.n119 163.367
R563 B.n121 B.n120 163.367
R564 B.n121 B.n94 163.367
R565 B.n125 B.n94 163.367
R566 B.n126 B.n125 163.367
R567 B.n127 B.n126 163.367
R568 B.n127 B.n92 163.367
R569 B.n131 B.n92 163.367
R570 B.n132 B.n131 163.367
R571 B.n133 B.n132 163.367
R572 B.n133 B.n90 163.367
R573 B.n137 B.n90 163.367
R574 B.n138 B.n137 163.367
R575 B.n139 B.n138 163.367
R576 B.n139 B.n88 163.367
R577 B.n143 B.n88 163.367
R578 B.n144 B.n143 163.367
R579 B.n145 B.n144 163.367
R580 B.n145 B.n86 163.367
R581 B.n162 B.n161 59.5399
R582 B.n180 B.n76 59.5399
R583 B.n307 B.n32 59.5399
R584 B.n26 B.n25 59.5399
R585 B.n161 B.n160 32.0005
R586 B.n76 B.n75 32.0005
R587 B.n32 B.n31 32.0005
R588 B.n25 B.n24 32.0005
R589 B.n337 B.n18 29.5029
R590 B.n294 B.n37 29.5029
R591 B.n194 B.n193 29.5029
R592 B.n148 B.n147 29.5029
R593 B B.n385 18.0485
R594 B.n338 B.n337 10.6151
R595 B.n339 B.n338 10.6151
R596 B.n339 B.n16 10.6151
R597 B.n343 B.n16 10.6151
R598 B.n344 B.n343 10.6151
R599 B.n345 B.n344 10.6151
R600 B.n345 B.n14 10.6151
R601 B.n349 B.n14 10.6151
R602 B.n350 B.n349 10.6151
R603 B.n351 B.n350 10.6151
R604 B.n351 B.n12 10.6151
R605 B.n355 B.n12 10.6151
R606 B.n356 B.n355 10.6151
R607 B.n357 B.n356 10.6151
R608 B.n357 B.n10 10.6151
R609 B.n361 B.n10 10.6151
R610 B.n362 B.n361 10.6151
R611 B.n363 B.n362 10.6151
R612 B.n363 B.n8 10.6151
R613 B.n367 B.n8 10.6151
R614 B.n368 B.n367 10.6151
R615 B.n369 B.n368 10.6151
R616 B.n369 B.n6 10.6151
R617 B.n373 B.n6 10.6151
R618 B.n374 B.n373 10.6151
R619 B.n375 B.n374 10.6151
R620 B.n375 B.n4 10.6151
R621 B.n379 B.n4 10.6151
R622 B.n380 B.n379 10.6151
R623 B.n381 B.n380 10.6151
R624 B.n381 B.n0 10.6151
R625 B.n333 B.n18 10.6151
R626 B.n333 B.n332 10.6151
R627 B.n332 B.n331 10.6151
R628 B.n331 B.n20 10.6151
R629 B.n327 B.n20 10.6151
R630 B.n327 B.n326 10.6151
R631 B.n326 B.n325 10.6151
R632 B.n325 B.n22 10.6151
R633 B.n321 B.n320 10.6151
R634 B.n320 B.n319 10.6151
R635 B.n319 B.n27 10.6151
R636 B.n315 B.n27 10.6151
R637 B.n315 B.n314 10.6151
R638 B.n314 B.n313 10.6151
R639 B.n313 B.n29 10.6151
R640 B.n309 B.n29 10.6151
R641 B.n309 B.n308 10.6151
R642 B.n306 B.n33 10.6151
R643 B.n302 B.n33 10.6151
R644 B.n302 B.n301 10.6151
R645 B.n301 B.n300 10.6151
R646 B.n300 B.n35 10.6151
R647 B.n296 B.n35 10.6151
R648 B.n296 B.n295 10.6151
R649 B.n295 B.n294 10.6151
R650 B.n290 B.n37 10.6151
R651 B.n290 B.n289 10.6151
R652 B.n289 B.n288 10.6151
R653 B.n288 B.n39 10.6151
R654 B.n284 B.n39 10.6151
R655 B.n284 B.n283 10.6151
R656 B.n283 B.n282 10.6151
R657 B.n282 B.n41 10.6151
R658 B.n278 B.n41 10.6151
R659 B.n278 B.n277 10.6151
R660 B.n277 B.n276 10.6151
R661 B.n276 B.n43 10.6151
R662 B.n272 B.n43 10.6151
R663 B.n272 B.n271 10.6151
R664 B.n271 B.n270 10.6151
R665 B.n270 B.n45 10.6151
R666 B.n266 B.n45 10.6151
R667 B.n266 B.n265 10.6151
R668 B.n265 B.n264 10.6151
R669 B.n264 B.n47 10.6151
R670 B.n260 B.n47 10.6151
R671 B.n260 B.n259 10.6151
R672 B.n259 B.n258 10.6151
R673 B.n258 B.n49 10.6151
R674 B.n254 B.n49 10.6151
R675 B.n254 B.n253 10.6151
R676 B.n253 B.n252 10.6151
R677 B.n252 B.n51 10.6151
R678 B.n248 B.n51 10.6151
R679 B.n248 B.n247 10.6151
R680 B.n247 B.n246 10.6151
R681 B.n246 B.n53 10.6151
R682 B.n242 B.n53 10.6151
R683 B.n242 B.n241 10.6151
R684 B.n241 B.n240 10.6151
R685 B.n240 B.n55 10.6151
R686 B.n236 B.n55 10.6151
R687 B.n236 B.n235 10.6151
R688 B.n235 B.n234 10.6151
R689 B.n234 B.n57 10.6151
R690 B.n230 B.n57 10.6151
R691 B.n230 B.n229 10.6151
R692 B.n229 B.n228 10.6151
R693 B.n228 B.n59 10.6151
R694 B.n224 B.n59 10.6151
R695 B.n224 B.n223 10.6151
R696 B.n223 B.n222 10.6151
R697 B.n222 B.n61 10.6151
R698 B.n218 B.n61 10.6151
R699 B.n218 B.n217 10.6151
R700 B.n217 B.n216 10.6151
R701 B.n216 B.n63 10.6151
R702 B.n212 B.n63 10.6151
R703 B.n212 B.n211 10.6151
R704 B.n211 B.n210 10.6151
R705 B.n210 B.n65 10.6151
R706 B.n206 B.n65 10.6151
R707 B.n206 B.n205 10.6151
R708 B.n205 B.n204 10.6151
R709 B.n204 B.n67 10.6151
R710 B.n200 B.n67 10.6151
R711 B.n200 B.n199 10.6151
R712 B.n199 B.n198 10.6151
R713 B.n198 B.n69 10.6151
R714 B.n194 B.n69 10.6151
R715 B.n101 B.n1 10.6151
R716 B.n104 B.n101 10.6151
R717 B.n105 B.n104 10.6151
R718 B.n106 B.n105 10.6151
R719 B.n106 B.n99 10.6151
R720 B.n110 B.n99 10.6151
R721 B.n111 B.n110 10.6151
R722 B.n112 B.n111 10.6151
R723 B.n112 B.n97 10.6151
R724 B.n116 B.n97 10.6151
R725 B.n117 B.n116 10.6151
R726 B.n118 B.n117 10.6151
R727 B.n118 B.n95 10.6151
R728 B.n122 B.n95 10.6151
R729 B.n123 B.n122 10.6151
R730 B.n124 B.n123 10.6151
R731 B.n124 B.n93 10.6151
R732 B.n128 B.n93 10.6151
R733 B.n129 B.n128 10.6151
R734 B.n130 B.n129 10.6151
R735 B.n130 B.n91 10.6151
R736 B.n134 B.n91 10.6151
R737 B.n135 B.n134 10.6151
R738 B.n136 B.n135 10.6151
R739 B.n136 B.n89 10.6151
R740 B.n140 B.n89 10.6151
R741 B.n141 B.n140 10.6151
R742 B.n142 B.n141 10.6151
R743 B.n142 B.n87 10.6151
R744 B.n146 B.n87 10.6151
R745 B.n147 B.n146 10.6151
R746 B.n148 B.n85 10.6151
R747 B.n152 B.n85 10.6151
R748 B.n153 B.n152 10.6151
R749 B.n154 B.n153 10.6151
R750 B.n154 B.n83 10.6151
R751 B.n158 B.n83 10.6151
R752 B.n159 B.n158 10.6151
R753 B.n163 B.n159 10.6151
R754 B.n167 B.n81 10.6151
R755 B.n168 B.n167 10.6151
R756 B.n169 B.n168 10.6151
R757 B.n169 B.n79 10.6151
R758 B.n173 B.n79 10.6151
R759 B.n174 B.n173 10.6151
R760 B.n175 B.n174 10.6151
R761 B.n175 B.n77 10.6151
R762 B.n179 B.n77 10.6151
R763 B.n182 B.n181 10.6151
R764 B.n182 B.n73 10.6151
R765 B.n186 B.n73 10.6151
R766 B.n187 B.n186 10.6151
R767 B.n188 B.n187 10.6151
R768 B.n188 B.n71 10.6151
R769 B.n192 B.n71 10.6151
R770 B.n193 B.n192 10.6151
R771 B.n26 B.n22 9.52245
R772 B.n307 B.n306 9.52245
R773 B.n163 B.n162 9.52245
R774 B.n181 B.n180 9.52245
R775 B.n385 B.n0 8.11757
R776 B.n385 B.n1 8.11757
R777 B.n321 B.n26 1.09318
R778 B.n308 B.n307 1.09318
R779 B.n162 B.n81 1.09318
R780 B.n180 B.n179 1.09318
C0 B VP 1.32978f
C1 VN VDD2 0.953778f
C2 w_n2620_n1154# B 5.07606f
C3 VTAIL VP 1.63402f
C4 w_n2620_n1154# VTAIL 1.43263f
C5 VDD1 B 0.959854f
C6 VDD2 B 1.01615f
C7 VDD1 VTAIL 3.19668f
C8 VN B 0.77404f
C9 VDD2 VTAIL 3.24252f
C10 w_n2620_n1154# VP 5.08602f
C11 VN VTAIL 1.61991f
C12 VDD1 VP 1.18683f
C13 VDD1 w_n2620_n1154# 1.2197f
C14 VDD2 VP 0.392016f
C15 VTAIL B 0.925897f
C16 VDD2 w_n2620_n1154# 1.27952f
C17 VN VP 4.05848f
C18 VN w_n2620_n1154# 4.75764f
C19 VDD1 VDD2 1.1362f
C20 VDD1 VN 0.156468f
C21 VDD2 VSUBS 0.77794f
C22 VDD1 VSUBS 1.182192f
C23 VTAIL VSUBS 0.325725f
C24 VN VSUBS 4.58362f
C25 VP VSUBS 1.695558f
C26 B VSUBS 2.490729f
C27 w_n2620_n1154# VSUBS 39.017002f
C28 B.n0 VSUBS 0.00882f
C29 B.n1 VSUBS 0.00882f
C30 B.n2 VSUBS 0.013045f
C31 B.n3 VSUBS 0.009996f
C32 B.n4 VSUBS 0.009996f
C33 B.n5 VSUBS 0.009996f
C34 B.n6 VSUBS 0.009996f
C35 B.n7 VSUBS 0.009996f
C36 B.n8 VSUBS 0.009996f
C37 B.n9 VSUBS 0.009996f
C38 B.n10 VSUBS 0.009996f
C39 B.n11 VSUBS 0.009996f
C40 B.n12 VSUBS 0.009996f
C41 B.n13 VSUBS 0.009996f
C42 B.n14 VSUBS 0.009996f
C43 B.n15 VSUBS 0.009996f
C44 B.n16 VSUBS 0.009996f
C45 B.n17 VSUBS 0.009996f
C46 B.n18 VSUBS 0.022558f
C47 B.n19 VSUBS 0.009996f
C48 B.n20 VSUBS 0.009996f
C49 B.n21 VSUBS 0.009996f
C50 B.n22 VSUBS 0.009482f
C51 B.n23 VSUBS 0.009996f
C52 B.t7 VSUBS 0.025745f
C53 B.t8 VSUBS 0.02772f
C54 B.t6 VSUBS 0.089513f
C55 B.n24 VSUBS 0.065847f
C56 B.n25 VSUBS 0.056231f
C57 B.n26 VSUBS 0.023161f
C58 B.n27 VSUBS 0.009996f
C59 B.n28 VSUBS 0.009996f
C60 B.n29 VSUBS 0.009996f
C61 B.n30 VSUBS 0.009996f
C62 B.t1 VSUBS 0.025745f
C63 B.t2 VSUBS 0.02772f
C64 B.t0 VSUBS 0.089507f
C65 B.n31 VSUBS 0.065854f
C66 B.n32 VSUBS 0.056231f
C67 B.n33 VSUBS 0.009996f
C68 B.n34 VSUBS 0.009996f
C69 B.n35 VSUBS 0.009996f
C70 B.n36 VSUBS 0.009996f
C71 B.n37 VSUBS 0.02125f
C72 B.n38 VSUBS 0.009996f
C73 B.n39 VSUBS 0.009996f
C74 B.n40 VSUBS 0.009996f
C75 B.n41 VSUBS 0.009996f
C76 B.n42 VSUBS 0.009996f
C77 B.n43 VSUBS 0.009996f
C78 B.n44 VSUBS 0.009996f
C79 B.n45 VSUBS 0.009996f
C80 B.n46 VSUBS 0.009996f
C81 B.n47 VSUBS 0.009996f
C82 B.n48 VSUBS 0.009996f
C83 B.n49 VSUBS 0.009996f
C84 B.n50 VSUBS 0.009996f
C85 B.n51 VSUBS 0.009996f
C86 B.n52 VSUBS 0.009996f
C87 B.n53 VSUBS 0.009996f
C88 B.n54 VSUBS 0.009996f
C89 B.n55 VSUBS 0.009996f
C90 B.n56 VSUBS 0.009996f
C91 B.n57 VSUBS 0.009996f
C92 B.n58 VSUBS 0.009996f
C93 B.n59 VSUBS 0.009996f
C94 B.n60 VSUBS 0.009996f
C95 B.n61 VSUBS 0.009996f
C96 B.n62 VSUBS 0.009996f
C97 B.n63 VSUBS 0.009996f
C98 B.n64 VSUBS 0.009996f
C99 B.n65 VSUBS 0.009996f
C100 B.n66 VSUBS 0.009996f
C101 B.n67 VSUBS 0.009996f
C102 B.n68 VSUBS 0.009996f
C103 B.n69 VSUBS 0.009996f
C104 B.n70 VSUBS 0.022558f
C105 B.n71 VSUBS 0.009996f
C106 B.n72 VSUBS 0.009996f
C107 B.n73 VSUBS 0.009996f
C108 B.n74 VSUBS 0.009996f
C109 B.t5 VSUBS 0.025745f
C110 B.t4 VSUBS 0.02772f
C111 B.t3 VSUBS 0.089507f
C112 B.n75 VSUBS 0.065854f
C113 B.n76 VSUBS 0.056231f
C114 B.n77 VSUBS 0.009996f
C115 B.n78 VSUBS 0.009996f
C116 B.n79 VSUBS 0.009996f
C117 B.n80 VSUBS 0.009996f
C118 B.n81 VSUBS 0.005513f
C119 B.n82 VSUBS 0.009996f
C120 B.n83 VSUBS 0.009996f
C121 B.n84 VSUBS 0.009996f
C122 B.n85 VSUBS 0.009996f
C123 B.n86 VSUBS 0.02125f
C124 B.n87 VSUBS 0.009996f
C125 B.n88 VSUBS 0.009996f
C126 B.n89 VSUBS 0.009996f
C127 B.n90 VSUBS 0.009996f
C128 B.n91 VSUBS 0.009996f
C129 B.n92 VSUBS 0.009996f
C130 B.n93 VSUBS 0.009996f
C131 B.n94 VSUBS 0.009996f
C132 B.n95 VSUBS 0.009996f
C133 B.n96 VSUBS 0.009996f
C134 B.n97 VSUBS 0.009996f
C135 B.n98 VSUBS 0.009996f
C136 B.n99 VSUBS 0.009996f
C137 B.n100 VSUBS 0.009996f
C138 B.n101 VSUBS 0.009996f
C139 B.n102 VSUBS 0.009996f
C140 B.n103 VSUBS 0.009996f
C141 B.n104 VSUBS 0.009996f
C142 B.n105 VSUBS 0.009996f
C143 B.n106 VSUBS 0.009996f
C144 B.n107 VSUBS 0.009996f
C145 B.n108 VSUBS 0.009996f
C146 B.n109 VSUBS 0.009996f
C147 B.n110 VSUBS 0.009996f
C148 B.n111 VSUBS 0.009996f
C149 B.n112 VSUBS 0.009996f
C150 B.n113 VSUBS 0.009996f
C151 B.n114 VSUBS 0.009996f
C152 B.n115 VSUBS 0.009996f
C153 B.n116 VSUBS 0.009996f
C154 B.n117 VSUBS 0.009996f
C155 B.n118 VSUBS 0.009996f
C156 B.n119 VSUBS 0.009996f
C157 B.n120 VSUBS 0.009996f
C158 B.n121 VSUBS 0.009996f
C159 B.n122 VSUBS 0.009996f
C160 B.n123 VSUBS 0.009996f
C161 B.n124 VSUBS 0.009996f
C162 B.n125 VSUBS 0.009996f
C163 B.n126 VSUBS 0.009996f
C164 B.n127 VSUBS 0.009996f
C165 B.n128 VSUBS 0.009996f
C166 B.n129 VSUBS 0.009996f
C167 B.n130 VSUBS 0.009996f
C168 B.n131 VSUBS 0.009996f
C169 B.n132 VSUBS 0.009996f
C170 B.n133 VSUBS 0.009996f
C171 B.n134 VSUBS 0.009996f
C172 B.n135 VSUBS 0.009996f
C173 B.n136 VSUBS 0.009996f
C174 B.n137 VSUBS 0.009996f
C175 B.n138 VSUBS 0.009996f
C176 B.n139 VSUBS 0.009996f
C177 B.n140 VSUBS 0.009996f
C178 B.n141 VSUBS 0.009996f
C179 B.n142 VSUBS 0.009996f
C180 B.n143 VSUBS 0.009996f
C181 B.n144 VSUBS 0.009996f
C182 B.n145 VSUBS 0.009996f
C183 B.n146 VSUBS 0.009996f
C184 B.n147 VSUBS 0.02125f
C185 B.n148 VSUBS 0.022558f
C186 B.n149 VSUBS 0.022558f
C187 B.n150 VSUBS 0.009996f
C188 B.n151 VSUBS 0.009996f
C189 B.n152 VSUBS 0.009996f
C190 B.n153 VSUBS 0.009996f
C191 B.n154 VSUBS 0.009996f
C192 B.n155 VSUBS 0.009996f
C193 B.n156 VSUBS 0.009996f
C194 B.n157 VSUBS 0.009996f
C195 B.n158 VSUBS 0.009996f
C196 B.n159 VSUBS 0.009996f
C197 B.t11 VSUBS 0.025745f
C198 B.t10 VSUBS 0.02772f
C199 B.t9 VSUBS 0.089513f
C200 B.n160 VSUBS 0.065847f
C201 B.n161 VSUBS 0.056231f
C202 B.n162 VSUBS 0.023161f
C203 B.n163 VSUBS 0.009482f
C204 B.n164 VSUBS 0.009996f
C205 B.n165 VSUBS 0.009996f
C206 B.n166 VSUBS 0.009996f
C207 B.n167 VSUBS 0.009996f
C208 B.n168 VSUBS 0.009996f
C209 B.n169 VSUBS 0.009996f
C210 B.n170 VSUBS 0.009996f
C211 B.n171 VSUBS 0.009996f
C212 B.n172 VSUBS 0.009996f
C213 B.n173 VSUBS 0.009996f
C214 B.n174 VSUBS 0.009996f
C215 B.n175 VSUBS 0.009996f
C216 B.n176 VSUBS 0.009996f
C217 B.n177 VSUBS 0.009996f
C218 B.n178 VSUBS 0.009996f
C219 B.n179 VSUBS 0.005513f
C220 B.n180 VSUBS 0.023161f
C221 B.n181 VSUBS 0.009482f
C222 B.n182 VSUBS 0.009996f
C223 B.n183 VSUBS 0.009996f
C224 B.n184 VSUBS 0.009996f
C225 B.n185 VSUBS 0.009996f
C226 B.n186 VSUBS 0.009996f
C227 B.n187 VSUBS 0.009996f
C228 B.n188 VSUBS 0.009996f
C229 B.n189 VSUBS 0.009996f
C230 B.n190 VSUBS 0.009996f
C231 B.n191 VSUBS 0.009996f
C232 B.n192 VSUBS 0.009996f
C233 B.n193 VSUBS 0.02125f
C234 B.n194 VSUBS 0.022558f
C235 B.n195 VSUBS 0.02125f
C236 B.n196 VSUBS 0.009996f
C237 B.n197 VSUBS 0.009996f
C238 B.n198 VSUBS 0.009996f
C239 B.n199 VSUBS 0.009996f
C240 B.n200 VSUBS 0.009996f
C241 B.n201 VSUBS 0.009996f
C242 B.n202 VSUBS 0.009996f
C243 B.n203 VSUBS 0.009996f
C244 B.n204 VSUBS 0.009996f
C245 B.n205 VSUBS 0.009996f
C246 B.n206 VSUBS 0.009996f
C247 B.n207 VSUBS 0.009996f
C248 B.n208 VSUBS 0.009996f
C249 B.n209 VSUBS 0.009996f
C250 B.n210 VSUBS 0.009996f
C251 B.n211 VSUBS 0.009996f
C252 B.n212 VSUBS 0.009996f
C253 B.n213 VSUBS 0.009996f
C254 B.n214 VSUBS 0.009996f
C255 B.n215 VSUBS 0.009996f
C256 B.n216 VSUBS 0.009996f
C257 B.n217 VSUBS 0.009996f
C258 B.n218 VSUBS 0.009996f
C259 B.n219 VSUBS 0.009996f
C260 B.n220 VSUBS 0.009996f
C261 B.n221 VSUBS 0.009996f
C262 B.n222 VSUBS 0.009996f
C263 B.n223 VSUBS 0.009996f
C264 B.n224 VSUBS 0.009996f
C265 B.n225 VSUBS 0.009996f
C266 B.n226 VSUBS 0.009996f
C267 B.n227 VSUBS 0.009996f
C268 B.n228 VSUBS 0.009996f
C269 B.n229 VSUBS 0.009996f
C270 B.n230 VSUBS 0.009996f
C271 B.n231 VSUBS 0.009996f
C272 B.n232 VSUBS 0.009996f
C273 B.n233 VSUBS 0.009996f
C274 B.n234 VSUBS 0.009996f
C275 B.n235 VSUBS 0.009996f
C276 B.n236 VSUBS 0.009996f
C277 B.n237 VSUBS 0.009996f
C278 B.n238 VSUBS 0.009996f
C279 B.n239 VSUBS 0.009996f
C280 B.n240 VSUBS 0.009996f
C281 B.n241 VSUBS 0.009996f
C282 B.n242 VSUBS 0.009996f
C283 B.n243 VSUBS 0.009996f
C284 B.n244 VSUBS 0.009996f
C285 B.n245 VSUBS 0.009996f
C286 B.n246 VSUBS 0.009996f
C287 B.n247 VSUBS 0.009996f
C288 B.n248 VSUBS 0.009996f
C289 B.n249 VSUBS 0.009996f
C290 B.n250 VSUBS 0.009996f
C291 B.n251 VSUBS 0.009996f
C292 B.n252 VSUBS 0.009996f
C293 B.n253 VSUBS 0.009996f
C294 B.n254 VSUBS 0.009996f
C295 B.n255 VSUBS 0.009996f
C296 B.n256 VSUBS 0.009996f
C297 B.n257 VSUBS 0.009996f
C298 B.n258 VSUBS 0.009996f
C299 B.n259 VSUBS 0.009996f
C300 B.n260 VSUBS 0.009996f
C301 B.n261 VSUBS 0.009996f
C302 B.n262 VSUBS 0.009996f
C303 B.n263 VSUBS 0.009996f
C304 B.n264 VSUBS 0.009996f
C305 B.n265 VSUBS 0.009996f
C306 B.n266 VSUBS 0.009996f
C307 B.n267 VSUBS 0.009996f
C308 B.n268 VSUBS 0.009996f
C309 B.n269 VSUBS 0.009996f
C310 B.n270 VSUBS 0.009996f
C311 B.n271 VSUBS 0.009996f
C312 B.n272 VSUBS 0.009996f
C313 B.n273 VSUBS 0.009996f
C314 B.n274 VSUBS 0.009996f
C315 B.n275 VSUBS 0.009996f
C316 B.n276 VSUBS 0.009996f
C317 B.n277 VSUBS 0.009996f
C318 B.n278 VSUBS 0.009996f
C319 B.n279 VSUBS 0.009996f
C320 B.n280 VSUBS 0.009996f
C321 B.n281 VSUBS 0.009996f
C322 B.n282 VSUBS 0.009996f
C323 B.n283 VSUBS 0.009996f
C324 B.n284 VSUBS 0.009996f
C325 B.n285 VSUBS 0.009996f
C326 B.n286 VSUBS 0.009996f
C327 B.n287 VSUBS 0.009996f
C328 B.n288 VSUBS 0.009996f
C329 B.n289 VSUBS 0.009996f
C330 B.n290 VSUBS 0.009996f
C331 B.n291 VSUBS 0.009996f
C332 B.n292 VSUBS 0.02125f
C333 B.n293 VSUBS 0.022558f
C334 B.n294 VSUBS 0.022558f
C335 B.n295 VSUBS 0.009996f
C336 B.n296 VSUBS 0.009996f
C337 B.n297 VSUBS 0.009996f
C338 B.n298 VSUBS 0.009996f
C339 B.n299 VSUBS 0.009996f
C340 B.n300 VSUBS 0.009996f
C341 B.n301 VSUBS 0.009996f
C342 B.n302 VSUBS 0.009996f
C343 B.n303 VSUBS 0.009996f
C344 B.n304 VSUBS 0.009996f
C345 B.n305 VSUBS 0.009996f
C346 B.n306 VSUBS 0.009482f
C347 B.n307 VSUBS 0.023161f
C348 B.n308 VSUBS 0.005513f
C349 B.n309 VSUBS 0.009996f
C350 B.n310 VSUBS 0.009996f
C351 B.n311 VSUBS 0.009996f
C352 B.n312 VSUBS 0.009996f
C353 B.n313 VSUBS 0.009996f
C354 B.n314 VSUBS 0.009996f
C355 B.n315 VSUBS 0.009996f
C356 B.n316 VSUBS 0.009996f
C357 B.n317 VSUBS 0.009996f
C358 B.n318 VSUBS 0.009996f
C359 B.n319 VSUBS 0.009996f
C360 B.n320 VSUBS 0.009996f
C361 B.n321 VSUBS 0.005513f
C362 B.n322 VSUBS 0.009996f
C363 B.n323 VSUBS 0.009996f
C364 B.n324 VSUBS 0.009996f
C365 B.n325 VSUBS 0.009996f
C366 B.n326 VSUBS 0.009996f
C367 B.n327 VSUBS 0.009996f
C368 B.n328 VSUBS 0.009996f
C369 B.n329 VSUBS 0.009996f
C370 B.n330 VSUBS 0.009996f
C371 B.n331 VSUBS 0.009996f
C372 B.n332 VSUBS 0.009996f
C373 B.n333 VSUBS 0.009996f
C374 B.n334 VSUBS 0.009996f
C375 B.n335 VSUBS 0.022558f
C376 B.n336 VSUBS 0.02125f
C377 B.n337 VSUBS 0.02125f
C378 B.n338 VSUBS 0.009996f
C379 B.n339 VSUBS 0.009996f
C380 B.n340 VSUBS 0.009996f
C381 B.n341 VSUBS 0.009996f
C382 B.n342 VSUBS 0.009996f
C383 B.n343 VSUBS 0.009996f
C384 B.n344 VSUBS 0.009996f
C385 B.n345 VSUBS 0.009996f
C386 B.n346 VSUBS 0.009996f
C387 B.n347 VSUBS 0.009996f
C388 B.n348 VSUBS 0.009996f
C389 B.n349 VSUBS 0.009996f
C390 B.n350 VSUBS 0.009996f
C391 B.n351 VSUBS 0.009996f
C392 B.n352 VSUBS 0.009996f
C393 B.n353 VSUBS 0.009996f
C394 B.n354 VSUBS 0.009996f
C395 B.n355 VSUBS 0.009996f
C396 B.n356 VSUBS 0.009996f
C397 B.n357 VSUBS 0.009996f
C398 B.n358 VSUBS 0.009996f
C399 B.n359 VSUBS 0.009996f
C400 B.n360 VSUBS 0.009996f
C401 B.n361 VSUBS 0.009996f
C402 B.n362 VSUBS 0.009996f
C403 B.n363 VSUBS 0.009996f
C404 B.n364 VSUBS 0.009996f
C405 B.n365 VSUBS 0.009996f
C406 B.n366 VSUBS 0.009996f
C407 B.n367 VSUBS 0.009996f
C408 B.n368 VSUBS 0.009996f
C409 B.n369 VSUBS 0.009996f
C410 B.n370 VSUBS 0.009996f
C411 B.n371 VSUBS 0.009996f
C412 B.n372 VSUBS 0.009996f
C413 B.n373 VSUBS 0.009996f
C414 B.n374 VSUBS 0.009996f
C415 B.n375 VSUBS 0.009996f
C416 B.n376 VSUBS 0.009996f
C417 B.n377 VSUBS 0.009996f
C418 B.n378 VSUBS 0.009996f
C419 B.n379 VSUBS 0.009996f
C420 B.n380 VSUBS 0.009996f
C421 B.n381 VSUBS 0.009996f
C422 B.n382 VSUBS 0.009996f
C423 B.n383 VSUBS 0.013045f
C424 B.n384 VSUBS 0.013896f
C425 B.n385 VSUBS 0.027634f
C426 VDD2.t0 VSUBS 0.01372f
C427 VDD2.t6 VSUBS 0.01372f
C428 VDD2.n0 VSUBS 0.037371f
C429 VDD2.t3 VSUBS 0.01372f
C430 VDD2.t7 VSUBS 0.01372f
C431 VDD2.n1 VSUBS 0.037371f
C432 VDD2.n2 VSUBS 1.38227f
C433 VDD2.t1 VSUBS 0.01372f
C434 VDD2.t5 VSUBS 0.01372f
C435 VDD2.n3 VSUBS 0.03709f
C436 VDD2.n4 VSUBS 1.20016f
C437 VDD2.t2 VSUBS 0.01372f
C438 VDD2.t4 VSUBS 0.01372f
C439 VDD2.n5 VSUBS 0.037369f
C440 VN.n0 VSUBS 0.056516f
C441 VN.t0 VSUBS 0.123349f
C442 VN.n1 VSUBS 0.095924f
C443 VN.n2 VSUBS 0.056516f
C444 VN.n3 VSUBS 0.061126f
C445 VN.t7 VSUBS 0.308399f
C446 VN.t1 VSUBS 0.123349f
C447 VN.n4 VSUBS 0.193128f
C448 VN.n5 VSUBS 0.193713f
C449 VN.n6 VSUBS 0.297653f
C450 VN.n7 VSUBS 0.056516f
C451 VN.n8 VSUBS 0.082503f
C452 VN.n9 VSUBS 0.082503f
C453 VN.t4 VSUBS 0.123349f
C454 VN.n10 VSUBS 0.116808f
C455 VN.n11 VSUBS 0.061126f
C456 VN.n12 VSUBS 0.056516f
C457 VN.n13 VSUBS 0.056516f
C458 VN.n14 VSUBS 0.056516f
C459 VN.n15 VSUBS 0.053389f
C460 VN.n16 VSUBS 0.084617f
C461 VN.n17 VSUBS 0.218346f
C462 VN.n18 VSUBS 0.052269f
C463 VN.n19 VSUBS 0.056516f
C464 VN.t6 VSUBS 0.123349f
C465 VN.n20 VSUBS 0.095924f
C466 VN.n21 VSUBS 0.056516f
C467 VN.t2 VSUBS 0.123349f
C468 VN.n22 VSUBS 0.116808f
C469 VN.n23 VSUBS 0.061126f
C470 VN.t3 VSUBS 0.308399f
C471 VN.t5 VSUBS 0.123349f
C472 VN.n24 VSUBS 0.193128f
C473 VN.n25 VSUBS 0.193713f
C474 VN.n26 VSUBS 0.297653f
C475 VN.n27 VSUBS 0.056516f
C476 VN.n28 VSUBS 0.082503f
C477 VN.n29 VSUBS 0.082503f
C478 VN.n30 VSUBS 0.061126f
C479 VN.n31 VSUBS 0.056516f
C480 VN.n32 VSUBS 0.056516f
C481 VN.n33 VSUBS 0.056516f
C482 VN.n34 VSUBS 0.053389f
C483 VN.n35 VSUBS 0.084617f
C484 VN.n36 VSUBS 0.218346f
C485 VN.n37 VSUBS 1.86146f
C486 VDD1.t5 VSUBS 0.013431f
C487 VDD1.t3 VSUBS 0.013431f
C488 VDD1.n0 VSUBS 0.036637f
C489 VDD1.t6 VSUBS 0.013431f
C490 VDD1.t0 VSUBS 0.013431f
C491 VDD1.n1 VSUBS 0.036582f
C492 VDD1.t2 VSUBS 0.013431f
C493 VDD1.t4 VSUBS 0.013431f
C494 VDD1.n2 VSUBS 0.036582f
C495 VDD1.n3 VSUBS 1.3919f
C496 VDD1.t1 VSUBS 0.013431f
C497 VDD1.t7 VSUBS 0.013431f
C498 VDD1.n4 VSUBS 0.036307f
C499 VDD1.n5 VSUBS 1.19669f
C500 VTAIL.t1 VSUBS 0.016653f
C501 VTAIL.t3 VSUBS 0.016653f
C502 VTAIL.n0 VSUBS 0.040546f
C503 VTAIL.n1 VSUBS 0.252871f
C504 VTAIL.t6 VSUBS 0.082276f
C505 VTAIL.n2 VSUBS 0.286614f
C506 VTAIL.t8 VSUBS 0.082276f
C507 VTAIL.n3 VSUBS 0.286614f
C508 VTAIL.t14 VSUBS 0.016653f
C509 VTAIL.t9 VSUBS 0.016653f
C510 VTAIL.n4 VSUBS 0.040546f
C511 VTAIL.n5 VSUBS 0.352479f
C512 VTAIL.t11 VSUBS 0.082276f
C513 VTAIL.n6 VSUBS 0.722505f
C514 VTAIL.t0 VSUBS 0.082276f
C515 VTAIL.n7 VSUBS 0.722505f
C516 VTAIL.t4 VSUBS 0.016653f
C517 VTAIL.t5 VSUBS 0.016653f
C518 VTAIL.n8 VSUBS 0.040546f
C519 VTAIL.n9 VSUBS 0.352479f
C520 VTAIL.t2 VSUBS 0.082276f
C521 VTAIL.n10 VSUBS 0.286614f
C522 VTAIL.t15 VSUBS 0.082276f
C523 VTAIL.n11 VSUBS 0.286614f
C524 VTAIL.t12 VSUBS 0.016653f
C525 VTAIL.t10 VSUBS 0.016653f
C526 VTAIL.n12 VSUBS 0.040546f
C527 VTAIL.n13 VSUBS 0.352479f
C528 VTAIL.t13 VSUBS 0.082276f
C529 VTAIL.n14 VSUBS 0.722505f
C530 VTAIL.t7 VSUBS 0.082276f
C531 VTAIL.n15 VSUBS 0.718256f
C532 VP.n0 VSUBS 0.058947f
C533 VP.t3 VSUBS 0.128656f
C534 VP.n1 VSUBS 0.100051f
C535 VP.n2 VSUBS 0.058947f
C536 VP.n3 VSUBS 0.063756f
C537 VP.n4 VSUBS 0.058947f
C538 VP.t1 VSUBS 0.128656f
C539 VP.n5 VSUBS 0.227739f
C540 VP.n6 VSUBS 0.058947f
C541 VP.t0 VSUBS 0.128656f
C542 VP.n7 VSUBS 0.100051f
C543 VP.n8 VSUBS 0.058947f
C544 VP.n9 VSUBS 0.063756f
C545 VP.t2 VSUBS 0.321666f
C546 VP.t4 VSUBS 0.128656f
C547 VP.n10 VSUBS 0.201436f
C548 VP.n11 VSUBS 0.202046f
C549 VP.n12 VSUBS 0.310458f
C550 VP.n13 VSUBS 0.058947f
C551 VP.n14 VSUBS 0.086052f
C552 VP.n15 VSUBS 0.086052f
C553 VP.t6 VSUBS 0.128656f
C554 VP.n16 VSUBS 0.121833f
C555 VP.n17 VSUBS 0.063756f
C556 VP.n18 VSUBS 0.058947f
C557 VP.n19 VSUBS 0.058947f
C558 VP.n20 VSUBS 0.058947f
C559 VP.n21 VSUBS 0.055686f
C560 VP.n22 VSUBS 0.088257f
C561 VP.n23 VSUBS 0.227739f
C562 VP.n24 VSUBS 1.90247f
C563 VP.n25 VSUBS 1.96066f
C564 VP.n26 VSUBS 0.058947f
C565 VP.n27 VSUBS 0.088257f
C566 VP.n28 VSUBS 0.055686f
C567 VP.t7 VSUBS 0.128656f
C568 VP.n29 VSUBS 0.121833f
C569 VP.n30 VSUBS 0.100051f
C570 VP.n31 VSUBS 0.058947f
C571 VP.n32 VSUBS 0.058947f
C572 VP.n33 VSUBS 0.058947f
C573 VP.n34 VSUBS 0.086052f
C574 VP.n35 VSUBS 0.086052f
C575 VP.t5 VSUBS 0.128656f
C576 VP.n36 VSUBS 0.121833f
C577 VP.n37 VSUBS 0.063756f
C578 VP.n38 VSUBS 0.058947f
C579 VP.n39 VSUBS 0.058947f
C580 VP.n40 VSUBS 0.058947f
C581 VP.n41 VSUBS 0.055686f
C582 VP.n42 VSUBS 0.088257f
C583 VP.n43 VSUBS 0.227739f
C584 VP.n44 VSUBS 0.054517f
.ends

