* NGSPICE file created from diff_pair_sample_0358.ext - technology: sky130A

.subckt diff_pair_sample_0358 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.46
X1 VTAIL.t14 VN.t0 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.46
X2 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.46
X3 VDD2.t4 VN.t1 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X4 VDD2.t3 VN.t2 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.46
X5 VDD1.t7 VP.t0 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.46
X6 VTAIL.t2 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.46
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.46
X8 VDD2.t2 VN.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X9 VTAIL.t10 VN.t4 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.46
X10 VTAIL.t3 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X11 VDD1.t4 VP.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X12 VDD2.t0 VN.t5 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.46
X13 VTAIL.t8 VN.t6 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X14 VTAIL.t1 VP.t4 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X15 VTAIL.t7 VN.t7 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X16 VDD1.t2 VP.t5 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.46
X17 VTAIL.t6 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.46
X18 VDD1.t0 VP.t7 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.46
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.46
R0 B.n97 B.t19 953.509
R1 B.n94 B.t15 953.509
R2 B.n395 B.t12 953.509
R3 B.n393 B.t8 953.509
R4 B.n695 B.n694 585
R5 B.n304 B.n92 585
R6 B.n303 B.n302 585
R7 B.n301 B.n300 585
R8 B.n299 B.n298 585
R9 B.n297 B.n296 585
R10 B.n295 B.n294 585
R11 B.n293 B.n292 585
R12 B.n291 B.n290 585
R13 B.n289 B.n288 585
R14 B.n287 B.n286 585
R15 B.n285 B.n284 585
R16 B.n283 B.n282 585
R17 B.n281 B.n280 585
R18 B.n279 B.n278 585
R19 B.n277 B.n276 585
R20 B.n275 B.n274 585
R21 B.n273 B.n272 585
R22 B.n271 B.n270 585
R23 B.n269 B.n268 585
R24 B.n267 B.n266 585
R25 B.n265 B.n264 585
R26 B.n263 B.n262 585
R27 B.n261 B.n260 585
R28 B.n259 B.n258 585
R29 B.n257 B.n256 585
R30 B.n255 B.n254 585
R31 B.n253 B.n252 585
R32 B.n251 B.n250 585
R33 B.n249 B.n248 585
R34 B.n247 B.n246 585
R35 B.n245 B.n244 585
R36 B.n243 B.n242 585
R37 B.n241 B.n240 585
R38 B.n239 B.n238 585
R39 B.n237 B.n236 585
R40 B.n235 B.n234 585
R41 B.n233 B.n232 585
R42 B.n231 B.n230 585
R43 B.n229 B.n228 585
R44 B.n227 B.n226 585
R45 B.n225 B.n224 585
R46 B.n223 B.n222 585
R47 B.n221 B.n220 585
R48 B.n219 B.n218 585
R49 B.n217 B.n216 585
R50 B.n215 B.n214 585
R51 B.n213 B.n212 585
R52 B.n211 B.n210 585
R53 B.n209 B.n208 585
R54 B.n207 B.n206 585
R55 B.n205 B.n204 585
R56 B.n203 B.n202 585
R57 B.n201 B.n200 585
R58 B.n199 B.n198 585
R59 B.n197 B.n196 585
R60 B.n195 B.n194 585
R61 B.n193 B.n192 585
R62 B.n191 B.n190 585
R63 B.n189 B.n188 585
R64 B.n187 B.n186 585
R65 B.n185 B.n184 585
R66 B.n183 B.n182 585
R67 B.n181 B.n180 585
R68 B.n179 B.n178 585
R69 B.n177 B.n176 585
R70 B.n175 B.n174 585
R71 B.n173 B.n172 585
R72 B.n171 B.n170 585
R73 B.n169 B.n168 585
R74 B.n167 B.n166 585
R75 B.n165 B.n164 585
R76 B.n163 B.n162 585
R77 B.n161 B.n160 585
R78 B.n159 B.n158 585
R79 B.n157 B.n156 585
R80 B.n155 B.n154 585
R81 B.n153 B.n152 585
R82 B.n151 B.n150 585
R83 B.n149 B.n148 585
R84 B.n147 B.n146 585
R85 B.n145 B.n144 585
R86 B.n143 B.n142 585
R87 B.n141 B.n140 585
R88 B.n139 B.n138 585
R89 B.n137 B.n136 585
R90 B.n135 B.n134 585
R91 B.n133 B.n132 585
R92 B.n131 B.n130 585
R93 B.n129 B.n128 585
R94 B.n127 B.n126 585
R95 B.n125 B.n124 585
R96 B.n123 B.n122 585
R97 B.n121 B.n120 585
R98 B.n119 B.n118 585
R99 B.n117 B.n116 585
R100 B.n115 B.n114 585
R101 B.n113 B.n112 585
R102 B.n111 B.n110 585
R103 B.n109 B.n108 585
R104 B.n107 B.n106 585
R105 B.n105 B.n104 585
R106 B.n103 B.n102 585
R107 B.n101 B.n100 585
R108 B.n40 B.n39 585
R109 B.n700 B.n699 585
R110 B.n693 B.n93 585
R111 B.n93 B.n37 585
R112 B.n692 B.n36 585
R113 B.n704 B.n36 585
R114 B.n691 B.n35 585
R115 B.n705 B.n35 585
R116 B.n690 B.n34 585
R117 B.n706 B.n34 585
R118 B.n689 B.n688 585
R119 B.n688 B.n33 585
R120 B.n687 B.n29 585
R121 B.n712 B.n29 585
R122 B.n686 B.n28 585
R123 B.n713 B.n28 585
R124 B.n685 B.n27 585
R125 B.n714 B.n27 585
R126 B.n684 B.n683 585
R127 B.n683 B.n23 585
R128 B.n682 B.n22 585
R129 B.n720 B.n22 585
R130 B.n681 B.n21 585
R131 B.n721 B.n21 585
R132 B.n680 B.n20 585
R133 B.n722 B.n20 585
R134 B.n679 B.n678 585
R135 B.n678 B.n19 585
R136 B.n677 B.n15 585
R137 B.n728 B.n15 585
R138 B.n676 B.n14 585
R139 B.n729 B.n14 585
R140 B.n675 B.n13 585
R141 B.n730 B.n13 585
R142 B.n674 B.n673 585
R143 B.n673 B.n12 585
R144 B.n672 B.n671 585
R145 B.n672 B.n8 585
R146 B.n670 B.n7 585
R147 B.n737 B.n7 585
R148 B.n669 B.n6 585
R149 B.n738 B.n6 585
R150 B.n668 B.n5 585
R151 B.n739 B.n5 585
R152 B.n667 B.n666 585
R153 B.n666 B.n4 585
R154 B.n665 B.n305 585
R155 B.n665 B.n664 585
R156 B.n654 B.n306 585
R157 B.n657 B.n306 585
R158 B.n656 B.n655 585
R159 B.n658 B.n656 585
R160 B.n653 B.n310 585
R161 B.n313 B.n310 585
R162 B.n652 B.n651 585
R163 B.n651 B.n650 585
R164 B.n312 B.n311 585
R165 B.n643 B.n312 585
R166 B.n642 B.n641 585
R167 B.n644 B.n642 585
R168 B.n640 B.n318 585
R169 B.n318 B.n317 585
R170 B.n639 B.n638 585
R171 B.n638 B.n637 585
R172 B.n320 B.n319 585
R173 B.n321 B.n320 585
R174 B.n630 B.n629 585
R175 B.n631 B.n630 585
R176 B.n628 B.n326 585
R177 B.n326 B.n325 585
R178 B.n627 B.n626 585
R179 B.n626 B.n625 585
R180 B.n328 B.n327 585
R181 B.n618 B.n328 585
R182 B.n617 B.n616 585
R183 B.n619 B.n617 585
R184 B.n615 B.n333 585
R185 B.n333 B.n332 585
R186 B.n614 B.n613 585
R187 B.n613 B.n612 585
R188 B.n335 B.n334 585
R189 B.n336 B.n335 585
R190 B.n608 B.n607 585
R191 B.n339 B.n338 585
R192 B.n604 B.n603 585
R193 B.n605 B.n604 585
R194 B.n602 B.n392 585
R195 B.n601 B.n600 585
R196 B.n599 B.n598 585
R197 B.n597 B.n596 585
R198 B.n595 B.n594 585
R199 B.n593 B.n592 585
R200 B.n591 B.n590 585
R201 B.n589 B.n588 585
R202 B.n587 B.n586 585
R203 B.n585 B.n584 585
R204 B.n583 B.n582 585
R205 B.n581 B.n580 585
R206 B.n579 B.n578 585
R207 B.n577 B.n576 585
R208 B.n575 B.n574 585
R209 B.n573 B.n572 585
R210 B.n571 B.n570 585
R211 B.n569 B.n568 585
R212 B.n567 B.n566 585
R213 B.n565 B.n564 585
R214 B.n563 B.n562 585
R215 B.n561 B.n560 585
R216 B.n559 B.n558 585
R217 B.n557 B.n556 585
R218 B.n555 B.n554 585
R219 B.n553 B.n552 585
R220 B.n551 B.n550 585
R221 B.n549 B.n548 585
R222 B.n547 B.n546 585
R223 B.n545 B.n544 585
R224 B.n543 B.n542 585
R225 B.n541 B.n540 585
R226 B.n539 B.n538 585
R227 B.n537 B.n536 585
R228 B.n535 B.n534 585
R229 B.n533 B.n532 585
R230 B.n531 B.n530 585
R231 B.n529 B.n528 585
R232 B.n527 B.n526 585
R233 B.n525 B.n524 585
R234 B.n523 B.n522 585
R235 B.n521 B.n520 585
R236 B.n519 B.n518 585
R237 B.n517 B.n516 585
R238 B.n515 B.n514 585
R239 B.n512 B.n511 585
R240 B.n510 B.n509 585
R241 B.n508 B.n507 585
R242 B.n506 B.n505 585
R243 B.n504 B.n503 585
R244 B.n502 B.n501 585
R245 B.n500 B.n499 585
R246 B.n498 B.n497 585
R247 B.n496 B.n495 585
R248 B.n494 B.n493 585
R249 B.n491 B.n490 585
R250 B.n489 B.n488 585
R251 B.n487 B.n486 585
R252 B.n485 B.n484 585
R253 B.n483 B.n482 585
R254 B.n481 B.n480 585
R255 B.n479 B.n478 585
R256 B.n477 B.n476 585
R257 B.n475 B.n474 585
R258 B.n473 B.n472 585
R259 B.n471 B.n470 585
R260 B.n469 B.n468 585
R261 B.n467 B.n466 585
R262 B.n465 B.n464 585
R263 B.n463 B.n462 585
R264 B.n461 B.n460 585
R265 B.n459 B.n458 585
R266 B.n457 B.n456 585
R267 B.n455 B.n454 585
R268 B.n453 B.n452 585
R269 B.n451 B.n450 585
R270 B.n449 B.n448 585
R271 B.n447 B.n446 585
R272 B.n445 B.n444 585
R273 B.n443 B.n442 585
R274 B.n441 B.n440 585
R275 B.n439 B.n438 585
R276 B.n437 B.n436 585
R277 B.n435 B.n434 585
R278 B.n433 B.n432 585
R279 B.n431 B.n430 585
R280 B.n429 B.n428 585
R281 B.n427 B.n426 585
R282 B.n425 B.n424 585
R283 B.n423 B.n422 585
R284 B.n421 B.n420 585
R285 B.n419 B.n418 585
R286 B.n417 B.n416 585
R287 B.n415 B.n414 585
R288 B.n413 B.n412 585
R289 B.n411 B.n410 585
R290 B.n409 B.n408 585
R291 B.n407 B.n406 585
R292 B.n405 B.n404 585
R293 B.n403 B.n402 585
R294 B.n401 B.n400 585
R295 B.n399 B.n398 585
R296 B.n397 B.n391 585
R297 B.n605 B.n391 585
R298 B.n609 B.n337 585
R299 B.n337 B.n336 585
R300 B.n611 B.n610 585
R301 B.n612 B.n611 585
R302 B.n331 B.n330 585
R303 B.n332 B.n331 585
R304 B.n621 B.n620 585
R305 B.n620 B.n619 585
R306 B.n622 B.n329 585
R307 B.n618 B.n329 585
R308 B.n624 B.n623 585
R309 B.n625 B.n624 585
R310 B.n324 B.n323 585
R311 B.n325 B.n324 585
R312 B.n633 B.n632 585
R313 B.n632 B.n631 585
R314 B.n634 B.n322 585
R315 B.n322 B.n321 585
R316 B.n636 B.n635 585
R317 B.n637 B.n636 585
R318 B.n316 B.n315 585
R319 B.n317 B.n316 585
R320 B.n646 B.n645 585
R321 B.n645 B.n644 585
R322 B.n647 B.n314 585
R323 B.n643 B.n314 585
R324 B.n649 B.n648 585
R325 B.n650 B.n649 585
R326 B.n309 B.n308 585
R327 B.n313 B.n309 585
R328 B.n660 B.n659 585
R329 B.n659 B.n658 585
R330 B.n661 B.n307 585
R331 B.n657 B.n307 585
R332 B.n663 B.n662 585
R333 B.n664 B.n663 585
R334 B.n3 B.n0 585
R335 B.n4 B.n3 585
R336 B.n736 B.n1 585
R337 B.n737 B.n736 585
R338 B.n735 B.n734 585
R339 B.n735 B.n8 585
R340 B.n733 B.n9 585
R341 B.n12 B.n9 585
R342 B.n732 B.n731 585
R343 B.n731 B.n730 585
R344 B.n11 B.n10 585
R345 B.n729 B.n11 585
R346 B.n727 B.n726 585
R347 B.n728 B.n727 585
R348 B.n725 B.n16 585
R349 B.n19 B.n16 585
R350 B.n724 B.n723 585
R351 B.n723 B.n722 585
R352 B.n18 B.n17 585
R353 B.n721 B.n18 585
R354 B.n719 B.n718 585
R355 B.n720 B.n719 585
R356 B.n717 B.n24 585
R357 B.n24 B.n23 585
R358 B.n716 B.n715 585
R359 B.n715 B.n714 585
R360 B.n26 B.n25 585
R361 B.n713 B.n26 585
R362 B.n711 B.n710 585
R363 B.n712 B.n711 585
R364 B.n709 B.n30 585
R365 B.n33 B.n30 585
R366 B.n708 B.n707 585
R367 B.n707 B.n706 585
R368 B.n32 B.n31 585
R369 B.n705 B.n32 585
R370 B.n703 B.n702 585
R371 B.n704 B.n703 585
R372 B.n701 B.n38 585
R373 B.n38 B.n37 585
R374 B.n740 B.n739 585
R375 B.n738 B.n2 585
R376 B.n699 B.n38 535.745
R377 B.n695 B.n93 535.745
R378 B.n391 B.n335 535.745
R379 B.n607 B.n337 535.745
R380 B.n94 B.t17 336.346
R381 B.n395 B.t14 336.346
R382 B.n97 B.t20 336.346
R383 B.n393 B.t11 336.346
R384 B.n95 B.t18 321.024
R385 B.n396 B.t13 321.024
R386 B.n98 B.t21 321.024
R387 B.n394 B.t10 321.024
R388 B.n697 B.n696 256.663
R389 B.n697 B.n91 256.663
R390 B.n697 B.n90 256.663
R391 B.n697 B.n89 256.663
R392 B.n697 B.n88 256.663
R393 B.n697 B.n87 256.663
R394 B.n697 B.n86 256.663
R395 B.n697 B.n85 256.663
R396 B.n697 B.n84 256.663
R397 B.n697 B.n83 256.663
R398 B.n697 B.n82 256.663
R399 B.n697 B.n81 256.663
R400 B.n697 B.n80 256.663
R401 B.n697 B.n79 256.663
R402 B.n697 B.n78 256.663
R403 B.n697 B.n77 256.663
R404 B.n697 B.n76 256.663
R405 B.n697 B.n75 256.663
R406 B.n697 B.n74 256.663
R407 B.n697 B.n73 256.663
R408 B.n697 B.n72 256.663
R409 B.n697 B.n71 256.663
R410 B.n697 B.n70 256.663
R411 B.n697 B.n69 256.663
R412 B.n697 B.n68 256.663
R413 B.n697 B.n67 256.663
R414 B.n697 B.n66 256.663
R415 B.n697 B.n65 256.663
R416 B.n697 B.n64 256.663
R417 B.n697 B.n63 256.663
R418 B.n697 B.n62 256.663
R419 B.n697 B.n61 256.663
R420 B.n697 B.n60 256.663
R421 B.n697 B.n59 256.663
R422 B.n697 B.n58 256.663
R423 B.n697 B.n57 256.663
R424 B.n697 B.n56 256.663
R425 B.n697 B.n55 256.663
R426 B.n697 B.n54 256.663
R427 B.n697 B.n53 256.663
R428 B.n697 B.n52 256.663
R429 B.n697 B.n51 256.663
R430 B.n697 B.n50 256.663
R431 B.n697 B.n49 256.663
R432 B.n697 B.n48 256.663
R433 B.n697 B.n47 256.663
R434 B.n697 B.n46 256.663
R435 B.n697 B.n45 256.663
R436 B.n697 B.n44 256.663
R437 B.n697 B.n43 256.663
R438 B.n697 B.n42 256.663
R439 B.n697 B.n41 256.663
R440 B.n698 B.n697 256.663
R441 B.n606 B.n605 256.663
R442 B.n605 B.n340 256.663
R443 B.n605 B.n341 256.663
R444 B.n605 B.n342 256.663
R445 B.n605 B.n343 256.663
R446 B.n605 B.n344 256.663
R447 B.n605 B.n345 256.663
R448 B.n605 B.n346 256.663
R449 B.n605 B.n347 256.663
R450 B.n605 B.n348 256.663
R451 B.n605 B.n349 256.663
R452 B.n605 B.n350 256.663
R453 B.n605 B.n351 256.663
R454 B.n605 B.n352 256.663
R455 B.n605 B.n353 256.663
R456 B.n605 B.n354 256.663
R457 B.n605 B.n355 256.663
R458 B.n605 B.n356 256.663
R459 B.n605 B.n357 256.663
R460 B.n605 B.n358 256.663
R461 B.n605 B.n359 256.663
R462 B.n605 B.n360 256.663
R463 B.n605 B.n361 256.663
R464 B.n605 B.n362 256.663
R465 B.n605 B.n363 256.663
R466 B.n605 B.n364 256.663
R467 B.n605 B.n365 256.663
R468 B.n605 B.n366 256.663
R469 B.n605 B.n367 256.663
R470 B.n605 B.n368 256.663
R471 B.n605 B.n369 256.663
R472 B.n605 B.n370 256.663
R473 B.n605 B.n371 256.663
R474 B.n605 B.n372 256.663
R475 B.n605 B.n373 256.663
R476 B.n605 B.n374 256.663
R477 B.n605 B.n375 256.663
R478 B.n605 B.n376 256.663
R479 B.n605 B.n377 256.663
R480 B.n605 B.n378 256.663
R481 B.n605 B.n379 256.663
R482 B.n605 B.n380 256.663
R483 B.n605 B.n381 256.663
R484 B.n605 B.n382 256.663
R485 B.n605 B.n383 256.663
R486 B.n605 B.n384 256.663
R487 B.n605 B.n385 256.663
R488 B.n605 B.n386 256.663
R489 B.n605 B.n387 256.663
R490 B.n605 B.n388 256.663
R491 B.n605 B.n389 256.663
R492 B.n605 B.n390 256.663
R493 B.n742 B.n741 256.663
R494 B.n100 B.n40 163.367
R495 B.n104 B.n103 163.367
R496 B.n108 B.n107 163.367
R497 B.n112 B.n111 163.367
R498 B.n116 B.n115 163.367
R499 B.n120 B.n119 163.367
R500 B.n124 B.n123 163.367
R501 B.n128 B.n127 163.367
R502 B.n132 B.n131 163.367
R503 B.n136 B.n135 163.367
R504 B.n140 B.n139 163.367
R505 B.n144 B.n143 163.367
R506 B.n148 B.n147 163.367
R507 B.n152 B.n151 163.367
R508 B.n156 B.n155 163.367
R509 B.n160 B.n159 163.367
R510 B.n164 B.n163 163.367
R511 B.n168 B.n167 163.367
R512 B.n172 B.n171 163.367
R513 B.n176 B.n175 163.367
R514 B.n180 B.n179 163.367
R515 B.n184 B.n183 163.367
R516 B.n188 B.n187 163.367
R517 B.n192 B.n191 163.367
R518 B.n196 B.n195 163.367
R519 B.n200 B.n199 163.367
R520 B.n204 B.n203 163.367
R521 B.n208 B.n207 163.367
R522 B.n212 B.n211 163.367
R523 B.n216 B.n215 163.367
R524 B.n220 B.n219 163.367
R525 B.n224 B.n223 163.367
R526 B.n228 B.n227 163.367
R527 B.n232 B.n231 163.367
R528 B.n236 B.n235 163.367
R529 B.n240 B.n239 163.367
R530 B.n244 B.n243 163.367
R531 B.n248 B.n247 163.367
R532 B.n252 B.n251 163.367
R533 B.n256 B.n255 163.367
R534 B.n260 B.n259 163.367
R535 B.n264 B.n263 163.367
R536 B.n268 B.n267 163.367
R537 B.n272 B.n271 163.367
R538 B.n276 B.n275 163.367
R539 B.n280 B.n279 163.367
R540 B.n284 B.n283 163.367
R541 B.n288 B.n287 163.367
R542 B.n292 B.n291 163.367
R543 B.n296 B.n295 163.367
R544 B.n300 B.n299 163.367
R545 B.n302 B.n92 163.367
R546 B.n613 B.n335 163.367
R547 B.n613 B.n333 163.367
R548 B.n617 B.n333 163.367
R549 B.n617 B.n328 163.367
R550 B.n626 B.n328 163.367
R551 B.n626 B.n326 163.367
R552 B.n630 B.n326 163.367
R553 B.n630 B.n320 163.367
R554 B.n638 B.n320 163.367
R555 B.n638 B.n318 163.367
R556 B.n642 B.n318 163.367
R557 B.n642 B.n312 163.367
R558 B.n651 B.n312 163.367
R559 B.n651 B.n310 163.367
R560 B.n656 B.n310 163.367
R561 B.n656 B.n306 163.367
R562 B.n665 B.n306 163.367
R563 B.n666 B.n665 163.367
R564 B.n666 B.n5 163.367
R565 B.n6 B.n5 163.367
R566 B.n7 B.n6 163.367
R567 B.n672 B.n7 163.367
R568 B.n673 B.n672 163.367
R569 B.n673 B.n13 163.367
R570 B.n14 B.n13 163.367
R571 B.n15 B.n14 163.367
R572 B.n678 B.n15 163.367
R573 B.n678 B.n20 163.367
R574 B.n21 B.n20 163.367
R575 B.n22 B.n21 163.367
R576 B.n683 B.n22 163.367
R577 B.n683 B.n27 163.367
R578 B.n28 B.n27 163.367
R579 B.n29 B.n28 163.367
R580 B.n688 B.n29 163.367
R581 B.n688 B.n34 163.367
R582 B.n35 B.n34 163.367
R583 B.n36 B.n35 163.367
R584 B.n93 B.n36 163.367
R585 B.n604 B.n339 163.367
R586 B.n604 B.n392 163.367
R587 B.n600 B.n599 163.367
R588 B.n596 B.n595 163.367
R589 B.n592 B.n591 163.367
R590 B.n588 B.n587 163.367
R591 B.n584 B.n583 163.367
R592 B.n580 B.n579 163.367
R593 B.n576 B.n575 163.367
R594 B.n572 B.n571 163.367
R595 B.n568 B.n567 163.367
R596 B.n564 B.n563 163.367
R597 B.n560 B.n559 163.367
R598 B.n556 B.n555 163.367
R599 B.n552 B.n551 163.367
R600 B.n548 B.n547 163.367
R601 B.n544 B.n543 163.367
R602 B.n540 B.n539 163.367
R603 B.n536 B.n535 163.367
R604 B.n532 B.n531 163.367
R605 B.n528 B.n527 163.367
R606 B.n524 B.n523 163.367
R607 B.n520 B.n519 163.367
R608 B.n516 B.n515 163.367
R609 B.n511 B.n510 163.367
R610 B.n507 B.n506 163.367
R611 B.n503 B.n502 163.367
R612 B.n499 B.n498 163.367
R613 B.n495 B.n494 163.367
R614 B.n490 B.n489 163.367
R615 B.n486 B.n485 163.367
R616 B.n482 B.n481 163.367
R617 B.n478 B.n477 163.367
R618 B.n474 B.n473 163.367
R619 B.n470 B.n469 163.367
R620 B.n466 B.n465 163.367
R621 B.n462 B.n461 163.367
R622 B.n458 B.n457 163.367
R623 B.n454 B.n453 163.367
R624 B.n450 B.n449 163.367
R625 B.n446 B.n445 163.367
R626 B.n442 B.n441 163.367
R627 B.n438 B.n437 163.367
R628 B.n434 B.n433 163.367
R629 B.n430 B.n429 163.367
R630 B.n426 B.n425 163.367
R631 B.n422 B.n421 163.367
R632 B.n418 B.n417 163.367
R633 B.n414 B.n413 163.367
R634 B.n410 B.n409 163.367
R635 B.n406 B.n405 163.367
R636 B.n402 B.n401 163.367
R637 B.n398 B.n391 163.367
R638 B.n611 B.n337 163.367
R639 B.n611 B.n331 163.367
R640 B.n620 B.n331 163.367
R641 B.n620 B.n329 163.367
R642 B.n624 B.n329 163.367
R643 B.n624 B.n324 163.367
R644 B.n632 B.n324 163.367
R645 B.n632 B.n322 163.367
R646 B.n636 B.n322 163.367
R647 B.n636 B.n316 163.367
R648 B.n645 B.n316 163.367
R649 B.n645 B.n314 163.367
R650 B.n649 B.n314 163.367
R651 B.n649 B.n309 163.367
R652 B.n659 B.n309 163.367
R653 B.n659 B.n307 163.367
R654 B.n663 B.n307 163.367
R655 B.n663 B.n3 163.367
R656 B.n740 B.n3 163.367
R657 B.n736 B.n2 163.367
R658 B.n736 B.n735 163.367
R659 B.n735 B.n9 163.367
R660 B.n731 B.n9 163.367
R661 B.n731 B.n11 163.367
R662 B.n727 B.n11 163.367
R663 B.n727 B.n16 163.367
R664 B.n723 B.n16 163.367
R665 B.n723 B.n18 163.367
R666 B.n719 B.n18 163.367
R667 B.n719 B.n24 163.367
R668 B.n715 B.n24 163.367
R669 B.n715 B.n26 163.367
R670 B.n711 B.n26 163.367
R671 B.n711 B.n30 163.367
R672 B.n707 B.n30 163.367
R673 B.n707 B.n32 163.367
R674 B.n703 B.n32 163.367
R675 B.n703 B.n38 163.367
R676 B.n605 B.n336 78.3505
R677 B.n697 B.n37 78.3505
R678 B.n699 B.n698 71.676
R679 B.n100 B.n41 71.676
R680 B.n104 B.n42 71.676
R681 B.n108 B.n43 71.676
R682 B.n112 B.n44 71.676
R683 B.n116 B.n45 71.676
R684 B.n120 B.n46 71.676
R685 B.n124 B.n47 71.676
R686 B.n128 B.n48 71.676
R687 B.n132 B.n49 71.676
R688 B.n136 B.n50 71.676
R689 B.n140 B.n51 71.676
R690 B.n144 B.n52 71.676
R691 B.n148 B.n53 71.676
R692 B.n152 B.n54 71.676
R693 B.n156 B.n55 71.676
R694 B.n160 B.n56 71.676
R695 B.n164 B.n57 71.676
R696 B.n168 B.n58 71.676
R697 B.n172 B.n59 71.676
R698 B.n176 B.n60 71.676
R699 B.n180 B.n61 71.676
R700 B.n184 B.n62 71.676
R701 B.n188 B.n63 71.676
R702 B.n192 B.n64 71.676
R703 B.n196 B.n65 71.676
R704 B.n200 B.n66 71.676
R705 B.n204 B.n67 71.676
R706 B.n208 B.n68 71.676
R707 B.n212 B.n69 71.676
R708 B.n216 B.n70 71.676
R709 B.n220 B.n71 71.676
R710 B.n224 B.n72 71.676
R711 B.n228 B.n73 71.676
R712 B.n232 B.n74 71.676
R713 B.n236 B.n75 71.676
R714 B.n240 B.n76 71.676
R715 B.n244 B.n77 71.676
R716 B.n248 B.n78 71.676
R717 B.n252 B.n79 71.676
R718 B.n256 B.n80 71.676
R719 B.n260 B.n81 71.676
R720 B.n264 B.n82 71.676
R721 B.n268 B.n83 71.676
R722 B.n272 B.n84 71.676
R723 B.n276 B.n85 71.676
R724 B.n280 B.n86 71.676
R725 B.n284 B.n87 71.676
R726 B.n288 B.n88 71.676
R727 B.n292 B.n89 71.676
R728 B.n296 B.n90 71.676
R729 B.n300 B.n91 71.676
R730 B.n696 B.n92 71.676
R731 B.n696 B.n695 71.676
R732 B.n302 B.n91 71.676
R733 B.n299 B.n90 71.676
R734 B.n295 B.n89 71.676
R735 B.n291 B.n88 71.676
R736 B.n287 B.n87 71.676
R737 B.n283 B.n86 71.676
R738 B.n279 B.n85 71.676
R739 B.n275 B.n84 71.676
R740 B.n271 B.n83 71.676
R741 B.n267 B.n82 71.676
R742 B.n263 B.n81 71.676
R743 B.n259 B.n80 71.676
R744 B.n255 B.n79 71.676
R745 B.n251 B.n78 71.676
R746 B.n247 B.n77 71.676
R747 B.n243 B.n76 71.676
R748 B.n239 B.n75 71.676
R749 B.n235 B.n74 71.676
R750 B.n231 B.n73 71.676
R751 B.n227 B.n72 71.676
R752 B.n223 B.n71 71.676
R753 B.n219 B.n70 71.676
R754 B.n215 B.n69 71.676
R755 B.n211 B.n68 71.676
R756 B.n207 B.n67 71.676
R757 B.n203 B.n66 71.676
R758 B.n199 B.n65 71.676
R759 B.n195 B.n64 71.676
R760 B.n191 B.n63 71.676
R761 B.n187 B.n62 71.676
R762 B.n183 B.n61 71.676
R763 B.n179 B.n60 71.676
R764 B.n175 B.n59 71.676
R765 B.n171 B.n58 71.676
R766 B.n167 B.n57 71.676
R767 B.n163 B.n56 71.676
R768 B.n159 B.n55 71.676
R769 B.n155 B.n54 71.676
R770 B.n151 B.n53 71.676
R771 B.n147 B.n52 71.676
R772 B.n143 B.n51 71.676
R773 B.n139 B.n50 71.676
R774 B.n135 B.n49 71.676
R775 B.n131 B.n48 71.676
R776 B.n127 B.n47 71.676
R777 B.n123 B.n46 71.676
R778 B.n119 B.n45 71.676
R779 B.n115 B.n44 71.676
R780 B.n111 B.n43 71.676
R781 B.n107 B.n42 71.676
R782 B.n103 B.n41 71.676
R783 B.n698 B.n40 71.676
R784 B.n607 B.n606 71.676
R785 B.n392 B.n340 71.676
R786 B.n599 B.n341 71.676
R787 B.n595 B.n342 71.676
R788 B.n591 B.n343 71.676
R789 B.n587 B.n344 71.676
R790 B.n583 B.n345 71.676
R791 B.n579 B.n346 71.676
R792 B.n575 B.n347 71.676
R793 B.n571 B.n348 71.676
R794 B.n567 B.n349 71.676
R795 B.n563 B.n350 71.676
R796 B.n559 B.n351 71.676
R797 B.n555 B.n352 71.676
R798 B.n551 B.n353 71.676
R799 B.n547 B.n354 71.676
R800 B.n543 B.n355 71.676
R801 B.n539 B.n356 71.676
R802 B.n535 B.n357 71.676
R803 B.n531 B.n358 71.676
R804 B.n527 B.n359 71.676
R805 B.n523 B.n360 71.676
R806 B.n519 B.n361 71.676
R807 B.n515 B.n362 71.676
R808 B.n510 B.n363 71.676
R809 B.n506 B.n364 71.676
R810 B.n502 B.n365 71.676
R811 B.n498 B.n366 71.676
R812 B.n494 B.n367 71.676
R813 B.n489 B.n368 71.676
R814 B.n485 B.n369 71.676
R815 B.n481 B.n370 71.676
R816 B.n477 B.n371 71.676
R817 B.n473 B.n372 71.676
R818 B.n469 B.n373 71.676
R819 B.n465 B.n374 71.676
R820 B.n461 B.n375 71.676
R821 B.n457 B.n376 71.676
R822 B.n453 B.n377 71.676
R823 B.n449 B.n378 71.676
R824 B.n445 B.n379 71.676
R825 B.n441 B.n380 71.676
R826 B.n437 B.n381 71.676
R827 B.n433 B.n382 71.676
R828 B.n429 B.n383 71.676
R829 B.n425 B.n384 71.676
R830 B.n421 B.n385 71.676
R831 B.n417 B.n386 71.676
R832 B.n413 B.n387 71.676
R833 B.n409 B.n388 71.676
R834 B.n405 B.n389 71.676
R835 B.n401 B.n390 71.676
R836 B.n606 B.n339 71.676
R837 B.n600 B.n340 71.676
R838 B.n596 B.n341 71.676
R839 B.n592 B.n342 71.676
R840 B.n588 B.n343 71.676
R841 B.n584 B.n344 71.676
R842 B.n580 B.n345 71.676
R843 B.n576 B.n346 71.676
R844 B.n572 B.n347 71.676
R845 B.n568 B.n348 71.676
R846 B.n564 B.n349 71.676
R847 B.n560 B.n350 71.676
R848 B.n556 B.n351 71.676
R849 B.n552 B.n352 71.676
R850 B.n548 B.n353 71.676
R851 B.n544 B.n354 71.676
R852 B.n540 B.n355 71.676
R853 B.n536 B.n356 71.676
R854 B.n532 B.n357 71.676
R855 B.n528 B.n358 71.676
R856 B.n524 B.n359 71.676
R857 B.n520 B.n360 71.676
R858 B.n516 B.n361 71.676
R859 B.n511 B.n362 71.676
R860 B.n507 B.n363 71.676
R861 B.n503 B.n364 71.676
R862 B.n499 B.n365 71.676
R863 B.n495 B.n366 71.676
R864 B.n490 B.n367 71.676
R865 B.n486 B.n368 71.676
R866 B.n482 B.n369 71.676
R867 B.n478 B.n370 71.676
R868 B.n474 B.n371 71.676
R869 B.n470 B.n372 71.676
R870 B.n466 B.n373 71.676
R871 B.n462 B.n374 71.676
R872 B.n458 B.n375 71.676
R873 B.n454 B.n376 71.676
R874 B.n450 B.n377 71.676
R875 B.n446 B.n378 71.676
R876 B.n442 B.n379 71.676
R877 B.n438 B.n380 71.676
R878 B.n434 B.n381 71.676
R879 B.n430 B.n382 71.676
R880 B.n426 B.n383 71.676
R881 B.n422 B.n384 71.676
R882 B.n418 B.n385 71.676
R883 B.n414 B.n386 71.676
R884 B.n410 B.n387 71.676
R885 B.n406 B.n388 71.676
R886 B.n402 B.n389 71.676
R887 B.n398 B.n390 71.676
R888 B.n741 B.n740 71.676
R889 B.n741 B.n2 71.676
R890 B.n99 B.n98 59.5399
R891 B.n96 B.n95 59.5399
R892 B.n492 B.n396 59.5399
R893 B.n513 B.n394 59.5399
R894 B.n612 B.n336 38.33
R895 B.n612 B.n332 38.33
R896 B.n619 B.n332 38.33
R897 B.n619 B.n618 38.33
R898 B.n625 B.n325 38.33
R899 B.n631 B.n325 38.33
R900 B.n631 B.n321 38.33
R901 B.n637 B.n321 38.33
R902 B.n644 B.n317 38.33
R903 B.n644 B.n643 38.33
R904 B.n650 B.n313 38.33
R905 B.n658 B.n657 38.33
R906 B.n664 B.n4 38.33
R907 B.n739 B.n4 38.33
R908 B.n739 B.n738 38.33
R909 B.n738 B.n737 38.33
R910 B.n737 B.n8 38.33
R911 B.n730 B.n12 38.33
R912 B.n729 B.n728 38.33
R913 B.n722 B.n19 38.33
R914 B.n722 B.n721 38.33
R915 B.n720 B.n23 38.33
R916 B.n714 B.n23 38.33
R917 B.n714 B.n713 38.33
R918 B.n713 B.n712 38.33
R919 B.n706 B.n33 38.33
R920 B.n706 B.n705 38.33
R921 B.n705 B.n704 38.33
R922 B.n704 B.n37 38.33
R923 B.n650 B.t4 34.948
R924 B.n728 B.t0 34.948
R925 B.n609 B.n608 34.8103
R926 B.n397 B.n334 34.8103
R927 B.n694 B.n693 34.8103
R928 B.n701 B.n700 34.8103
R929 B.n625 B.t9 29.3113
R930 B.n637 B.t1 29.3113
R931 B.t7 B.n720 29.3113
R932 B.n712 B.t16 29.3113
R933 B.n657 B.t6 28.1839
R934 B.n12 B.t3 28.1839
R935 B.n658 B.t5 22.5473
R936 B.n730 B.t2 22.5473
R937 B B.n742 18.0485
R938 B.n313 B.t5 15.7832
R939 B.t2 B.n729 15.7832
R940 B.n98 B.n97 15.3217
R941 B.n95 B.n94 15.3217
R942 B.n396 B.n395 15.3217
R943 B.n394 B.n393 15.3217
R944 B.n610 B.n609 10.6151
R945 B.n610 B.n330 10.6151
R946 B.n621 B.n330 10.6151
R947 B.n622 B.n621 10.6151
R948 B.n623 B.n622 10.6151
R949 B.n623 B.n323 10.6151
R950 B.n633 B.n323 10.6151
R951 B.n634 B.n633 10.6151
R952 B.n635 B.n634 10.6151
R953 B.n635 B.n315 10.6151
R954 B.n646 B.n315 10.6151
R955 B.n647 B.n646 10.6151
R956 B.n648 B.n647 10.6151
R957 B.n648 B.n308 10.6151
R958 B.n660 B.n308 10.6151
R959 B.n661 B.n660 10.6151
R960 B.n662 B.n661 10.6151
R961 B.n662 B.n0 10.6151
R962 B.n608 B.n338 10.6151
R963 B.n603 B.n338 10.6151
R964 B.n603 B.n602 10.6151
R965 B.n602 B.n601 10.6151
R966 B.n601 B.n598 10.6151
R967 B.n598 B.n597 10.6151
R968 B.n597 B.n594 10.6151
R969 B.n594 B.n593 10.6151
R970 B.n593 B.n590 10.6151
R971 B.n590 B.n589 10.6151
R972 B.n589 B.n586 10.6151
R973 B.n586 B.n585 10.6151
R974 B.n585 B.n582 10.6151
R975 B.n582 B.n581 10.6151
R976 B.n581 B.n578 10.6151
R977 B.n578 B.n577 10.6151
R978 B.n577 B.n574 10.6151
R979 B.n574 B.n573 10.6151
R980 B.n573 B.n570 10.6151
R981 B.n570 B.n569 10.6151
R982 B.n569 B.n566 10.6151
R983 B.n566 B.n565 10.6151
R984 B.n565 B.n562 10.6151
R985 B.n562 B.n561 10.6151
R986 B.n561 B.n558 10.6151
R987 B.n558 B.n557 10.6151
R988 B.n557 B.n554 10.6151
R989 B.n554 B.n553 10.6151
R990 B.n553 B.n550 10.6151
R991 B.n550 B.n549 10.6151
R992 B.n549 B.n546 10.6151
R993 B.n546 B.n545 10.6151
R994 B.n545 B.n542 10.6151
R995 B.n542 B.n541 10.6151
R996 B.n541 B.n538 10.6151
R997 B.n538 B.n537 10.6151
R998 B.n537 B.n534 10.6151
R999 B.n534 B.n533 10.6151
R1000 B.n533 B.n530 10.6151
R1001 B.n530 B.n529 10.6151
R1002 B.n529 B.n526 10.6151
R1003 B.n526 B.n525 10.6151
R1004 B.n525 B.n522 10.6151
R1005 B.n522 B.n521 10.6151
R1006 B.n521 B.n518 10.6151
R1007 B.n518 B.n517 10.6151
R1008 B.n517 B.n514 10.6151
R1009 B.n512 B.n509 10.6151
R1010 B.n509 B.n508 10.6151
R1011 B.n508 B.n505 10.6151
R1012 B.n505 B.n504 10.6151
R1013 B.n504 B.n501 10.6151
R1014 B.n501 B.n500 10.6151
R1015 B.n500 B.n497 10.6151
R1016 B.n497 B.n496 10.6151
R1017 B.n496 B.n493 10.6151
R1018 B.n491 B.n488 10.6151
R1019 B.n488 B.n487 10.6151
R1020 B.n487 B.n484 10.6151
R1021 B.n484 B.n483 10.6151
R1022 B.n483 B.n480 10.6151
R1023 B.n480 B.n479 10.6151
R1024 B.n479 B.n476 10.6151
R1025 B.n476 B.n475 10.6151
R1026 B.n475 B.n472 10.6151
R1027 B.n472 B.n471 10.6151
R1028 B.n471 B.n468 10.6151
R1029 B.n468 B.n467 10.6151
R1030 B.n467 B.n464 10.6151
R1031 B.n464 B.n463 10.6151
R1032 B.n463 B.n460 10.6151
R1033 B.n460 B.n459 10.6151
R1034 B.n459 B.n456 10.6151
R1035 B.n456 B.n455 10.6151
R1036 B.n455 B.n452 10.6151
R1037 B.n452 B.n451 10.6151
R1038 B.n451 B.n448 10.6151
R1039 B.n448 B.n447 10.6151
R1040 B.n447 B.n444 10.6151
R1041 B.n444 B.n443 10.6151
R1042 B.n443 B.n440 10.6151
R1043 B.n440 B.n439 10.6151
R1044 B.n439 B.n436 10.6151
R1045 B.n436 B.n435 10.6151
R1046 B.n435 B.n432 10.6151
R1047 B.n432 B.n431 10.6151
R1048 B.n431 B.n428 10.6151
R1049 B.n428 B.n427 10.6151
R1050 B.n427 B.n424 10.6151
R1051 B.n424 B.n423 10.6151
R1052 B.n423 B.n420 10.6151
R1053 B.n420 B.n419 10.6151
R1054 B.n419 B.n416 10.6151
R1055 B.n416 B.n415 10.6151
R1056 B.n415 B.n412 10.6151
R1057 B.n412 B.n411 10.6151
R1058 B.n411 B.n408 10.6151
R1059 B.n408 B.n407 10.6151
R1060 B.n407 B.n404 10.6151
R1061 B.n404 B.n403 10.6151
R1062 B.n403 B.n400 10.6151
R1063 B.n400 B.n399 10.6151
R1064 B.n399 B.n397 10.6151
R1065 B.n614 B.n334 10.6151
R1066 B.n615 B.n614 10.6151
R1067 B.n616 B.n615 10.6151
R1068 B.n616 B.n327 10.6151
R1069 B.n627 B.n327 10.6151
R1070 B.n628 B.n627 10.6151
R1071 B.n629 B.n628 10.6151
R1072 B.n629 B.n319 10.6151
R1073 B.n639 B.n319 10.6151
R1074 B.n640 B.n639 10.6151
R1075 B.n641 B.n640 10.6151
R1076 B.n641 B.n311 10.6151
R1077 B.n652 B.n311 10.6151
R1078 B.n653 B.n652 10.6151
R1079 B.n655 B.n653 10.6151
R1080 B.n655 B.n654 10.6151
R1081 B.n654 B.n305 10.6151
R1082 B.n667 B.n305 10.6151
R1083 B.n668 B.n667 10.6151
R1084 B.n669 B.n668 10.6151
R1085 B.n670 B.n669 10.6151
R1086 B.n671 B.n670 10.6151
R1087 B.n674 B.n671 10.6151
R1088 B.n675 B.n674 10.6151
R1089 B.n676 B.n675 10.6151
R1090 B.n677 B.n676 10.6151
R1091 B.n679 B.n677 10.6151
R1092 B.n680 B.n679 10.6151
R1093 B.n681 B.n680 10.6151
R1094 B.n682 B.n681 10.6151
R1095 B.n684 B.n682 10.6151
R1096 B.n685 B.n684 10.6151
R1097 B.n686 B.n685 10.6151
R1098 B.n687 B.n686 10.6151
R1099 B.n689 B.n687 10.6151
R1100 B.n690 B.n689 10.6151
R1101 B.n691 B.n690 10.6151
R1102 B.n692 B.n691 10.6151
R1103 B.n693 B.n692 10.6151
R1104 B.n734 B.n1 10.6151
R1105 B.n734 B.n733 10.6151
R1106 B.n733 B.n732 10.6151
R1107 B.n732 B.n10 10.6151
R1108 B.n726 B.n10 10.6151
R1109 B.n726 B.n725 10.6151
R1110 B.n725 B.n724 10.6151
R1111 B.n724 B.n17 10.6151
R1112 B.n718 B.n17 10.6151
R1113 B.n718 B.n717 10.6151
R1114 B.n717 B.n716 10.6151
R1115 B.n716 B.n25 10.6151
R1116 B.n710 B.n25 10.6151
R1117 B.n710 B.n709 10.6151
R1118 B.n709 B.n708 10.6151
R1119 B.n708 B.n31 10.6151
R1120 B.n702 B.n31 10.6151
R1121 B.n702 B.n701 10.6151
R1122 B.n700 B.n39 10.6151
R1123 B.n101 B.n39 10.6151
R1124 B.n102 B.n101 10.6151
R1125 B.n105 B.n102 10.6151
R1126 B.n106 B.n105 10.6151
R1127 B.n109 B.n106 10.6151
R1128 B.n110 B.n109 10.6151
R1129 B.n113 B.n110 10.6151
R1130 B.n114 B.n113 10.6151
R1131 B.n117 B.n114 10.6151
R1132 B.n118 B.n117 10.6151
R1133 B.n121 B.n118 10.6151
R1134 B.n122 B.n121 10.6151
R1135 B.n125 B.n122 10.6151
R1136 B.n126 B.n125 10.6151
R1137 B.n129 B.n126 10.6151
R1138 B.n130 B.n129 10.6151
R1139 B.n133 B.n130 10.6151
R1140 B.n134 B.n133 10.6151
R1141 B.n137 B.n134 10.6151
R1142 B.n138 B.n137 10.6151
R1143 B.n141 B.n138 10.6151
R1144 B.n142 B.n141 10.6151
R1145 B.n145 B.n142 10.6151
R1146 B.n146 B.n145 10.6151
R1147 B.n149 B.n146 10.6151
R1148 B.n150 B.n149 10.6151
R1149 B.n153 B.n150 10.6151
R1150 B.n154 B.n153 10.6151
R1151 B.n157 B.n154 10.6151
R1152 B.n158 B.n157 10.6151
R1153 B.n161 B.n158 10.6151
R1154 B.n162 B.n161 10.6151
R1155 B.n165 B.n162 10.6151
R1156 B.n166 B.n165 10.6151
R1157 B.n169 B.n166 10.6151
R1158 B.n170 B.n169 10.6151
R1159 B.n173 B.n170 10.6151
R1160 B.n174 B.n173 10.6151
R1161 B.n177 B.n174 10.6151
R1162 B.n178 B.n177 10.6151
R1163 B.n181 B.n178 10.6151
R1164 B.n182 B.n181 10.6151
R1165 B.n185 B.n182 10.6151
R1166 B.n186 B.n185 10.6151
R1167 B.n189 B.n186 10.6151
R1168 B.n190 B.n189 10.6151
R1169 B.n194 B.n193 10.6151
R1170 B.n197 B.n194 10.6151
R1171 B.n198 B.n197 10.6151
R1172 B.n201 B.n198 10.6151
R1173 B.n202 B.n201 10.6151
R1174 B.n205 B.n202 10.6151
R1175 B.n206 B.n205 10.6151
R1176 B.n209 B.n206 10.6151
R1177 B.n210 B.n209 10.6151
R1178 B.n214 B.n213 10.6151
R1179 B.n217 B.n214 10.6151
R1180 B.n218 B.n217 10.6151
R1181 B.n221 B.n218 10.6151
R1182 B.n222 B.n221 10.6151
R1183 B.n225 B.n222 10.6151
R1184 B.n226 B.n225 10.6151
R1185 B.n229 B.n226 10.6151
R1186 B.n230 B.n229 10.6151
R1187 B.n233 B.n230 10.6151
R1188 B.n234 B.n233 10.6151
R1189 B.n237 B.n234 10.6151
R1190 B.n238 B.n237 10.6151
R1191 B.n241 B.n238 10.6151
R1192 B.n242 B.n241 10.6151
R1193 B.n245 B.n242 10.6151
R1194 B.n246 B.n245 10.6151
R1195 B.n249 B.n246 10.6151
R1196 B.n250 B.n249 10.6151
R1197 B.n253 B.n250 10.6151
R1198 B.n254 B.n253 10.6151
R1199 B.n257 B.n254 10.6151
R1200 B.n258 B.n257 10.6151
R1201 B.n261 B.n258 10.6151
R1202 B.n262 B.n261 10.6151
R1203 B.n265 B.n262 10.6151
R1204 B.n266 B.n265 10.6151
R1205 B.n269 B.n266 10.6151
R1206 B.n270 B.n269 10.6151
R1207 B.n273 B.n270 10.6151
R1208 B.n274 B.n273 10.6151
R1209 B.n277 B.n274 10.6151
R1210 B.n278 B.n277 10.6151
R1211 B.n281 B.n278 10.6151
R1212 B.n282 B.n281 10.6151
R1213 B.n285 B.n282 10.6151
R1214 B.n286 B.n285 10.6151
R1215 B.n289 B.n286 10.6151
R1216 B.n290 B.n289 10.6151
R1217 B.n293 B.n290 10.6151
R1218 B.n294 B.n293 10.6151
R1219 B.n297 B.n294 10.6151
R1220 B.n298 B.n297 10.6151
R1221 B.n301 B.n298 10.6151
R1222 B.n303 B.n301 10.6151
R1223 B.n304 B.n303 10.6151
R1224 B.n694 B.n304 10.6151
R1225 B.n664 B.t6 10.1465
R1226 B.t3 B.n8 10.1465
R1227 B.n514 B.n513 9.36635
R1228 B.n492 B.n491 9.36635
R1229 B.n190 B.n99 9.36635
R1230 B.n213 B.n96 9.36635
R1231 B.n618 B.t9 9.0192
R1232 B.t1 B.n317 9.0192
R1233 B.n721 B.t7 9.0192
R1234 B.n33 B.t16 9.0192
R1235 B.n742 B.n0 8.11757
R1236 B.n742 B.n1 8.11757
R1237 B.n643 B.t4 3.38251
R1238 B.n19 B.t0 3.38251
R1239 B.n513 B.n512 1.24928
R1240 B.n493 B.n492 1.24928
R1241 B.n193 B.n99 1.24928
R1242 B.n210 B.n96 1.24928
R1243 VN.n2 VN.t0 853.48
R1244 VN.n10 VN.t5 853.48
R1245 VN.n1 VN.t1 832.499
R1246 VN.n5 VN.t7 832.499
R1247 VN.n6 VN.t2 832.499
R1248 VN.n9 VN.t6 832.499
R1249 VN.n13 VN.t3 832.499
R1250 VN.n14 VN.t4 832.499
R1251 VN.n7 VN.n6 161.3
R1252 VN.n15 VN.n14 161.3
R1253 VN.n13 VN.n8 161.3
R1254 VN.n12 VN.n11 161.3
R1255 VN.n5 VN.n0 161.3
R1256 VN.n4 VN.n3 161.3
R1257 VN.n11 VN.n10 70.4033
R1258 VN.n3 VN.n2 70.4033
R1259 VN.n6 VN.n5 48.2005
R1260 VN.n14 VN.n13 48.2005
R1261 VN VN.n15 42.9948
R1262 VN.n4 VN.n1 24.1005
R1263 VN.n5 VN.n4 24.1005
R1264 VN.n13 VN.n12 24.1005
R1265 VN.n12 VN.n9 24.1005
R1266 VN.n10 VN.n9 20.9576
R1267 VN.n2 VN.n1 20.9576
R1268 VN.n15 VN.n8 0.189894
R1269 VN.n11 VN.n8 0.189894
R1270 VN.n3 VN.n0 0.189894
R1271 VN.n7 VN.n0 0.189894
R1272 VN VN.n7 0.0516364
R1273 VDD2.n2 VDD2.n1 60.9376
R1274 VDD2.n2 VDD2.n0 60.9376
R1275 VDD2 VDD2.n5 60.9348
R1276 VDD2.n4 VDD2.n3 60.6524
R1277 VDD2.n4 VDD2.n2 39.0558
R1278 VDD2.n5 VDD2.t7 1.39095
R1279 VDD2.n5 VDD2.t0 1.39095
R1280 VDD2.n3 VDD2.t6 1.39095
R1281 VDD2.n3 VDD2.t2 1.39095
R1282 VDD2.n1 VDD2.t1 1.39095
R1283 VDD2.n1 VDD2.t3 1.39095
R1284 VDD2.n0 VDD2.t5 1.39095
R1285 VDD2.n0 VDD2.t4 1.39095
R1286 VDD2 VDD2.n4 0.399207
R1287 VTAIL.n626 VTAIL.n554 289.615
R1288 VTAIL.n74 VTAIL.n2 289.615
R1289 VTAIL.n152 VTAIL.n80 289.615
R1290 VTAIL.n232 VTAIL.n160 289.615
R1291 VTAIL.n548 VTAIL.n476 289.615
R1292 VTAIL.n468 VTAIL.n396 289.615
R1293 VTAIL.n390 VTAIL.n318 289.615
R1294 VTAIL.n310 VTAIL.n238 289.615
R1295 VTAIL.n578 VTAIL.n577 185
R1296 VTAIL.n583 VTAIL.n582 185
R1297 VTAIL.n585 VTAIL.n584 185
R1298 VTAIL.n574 VTAIL.n573 185
R1299 VTAIL.n591 VTAIL.n590 185
R1300 VTAIL.n593 VTAIL.n592 185
R1301 VTAIL.n570 VTAIL.n569 185
R1302 VTAIL.n600 VTAIL.n599 185
R1303 VTAIL.n601 VTAIL.n568 185
R1304 VTAIL.n603 VTAIL.n602 185
R1305 VTAIL.n566 VTAIL.n565 185
R1306 VTAIL.n609 VTAIL.n608 185
R1307 VTAIL.n611 VTAIL.n610 185
R1308 VTAIL.n562 VTAIL.n561 185
R1309 VTAIL.n617 VTAIL.n616 185
R1310 VTAIL.n619 VTAIL.n618 185
R1311 VTAIL.n558 VTAIL.n557 185
R1312 VTAIL.n625 VTAIL.n624 185
R1313 VTAIL.n627 VTAIL.n626 185
R1314 VTAIL.n26 VTAIL.n25 185
R1315 VTAIL.n31 VTAIL.n30 185
R1316 VTAIL.n33 VTAIL.n32 185
R1317 VTAIL.n22 VTAIL.n21 185
R1318 VTAIL.n39 VTAIL.n38 185
R1319 VTAIL.n41 VTAIL.n40 185
R1320 VTAIL.n18 VTAIL.n17 185
R1321 VTAIL.n48 VTAIL.n47 185
R1322 VTAIL.n49 VTAIL.n16 185
R1323 VTAIL.n51 VTAIL.n50 185
R1324 VTAIL.n14 VTAIL.n13 185
R1325 VTAIL.n57 VTAIL.n56 185
R1326 VTAIL.n59 VTAIL.n58 185
R1327 VTAIL.n10 VTAIL.n9 185
R1328 VTAIL.n65 VTAIL.n64 185
R1329 VTAIL.n67 VTAIL.n66 185
R1330 VTAIL.n6 VTAIL.n5 185
R1331 VTAIL.n73 VTAIL.n72 185
R1332 VTAIL.n75 VTAIL.n74 185
R1333 VTAIL.n104 VTAIL.n103 185
R1334 VTAIL.n109 VTAIL.n108 185
R1335 VTAIL.n111 VTAIL.n110 185
R1336 VTAIL.n100 VTAIL.n99 185
R1337 VTAIL.n117 VTAIL.n116 185
R1338 VTAIL.n119 VTAIL.n118 185
R1339 VTAIL.n96 VTAIL.n95 185
R1340 VTAIL.n126 VTAIL.n125 185
R1341 VTAIL.n127 VTAIL.n94 185
R1342 VTAIL.n129 VTAIL.n128 185
R1343 VTAIL.n92 VTAIL.n91 185
R1344 VTAIL.n135 VTAIL.n134 185
R1345 VTAIL.n137 VTAIL.n136 185
R1346 VTAIL.n88 VTAIL.n87 185
R1347 VTAIL.n143 VTAIL.n142 185
R1348 VTAIL.n145 VTAIL.n144 185
R1349 VTAIL.n84 VTAIL.n83 185
R1350 VTAIL.n151 VTAIL.n150 185
R1351 VTAIL.n153 VTAIL.n152 185
R1352 VTAIL.n184 VTAIL.n183 185
R1353 VTAIL.n189 VTAIL.n188 185
R1354 VTAIL.n191 VTAIL.n190 185
R1355 VTAIL.n180 VTAIL.n179 185
R1356 VTAIL.n197 VTAIL.n196 185
R1357 VTAIL.n199 VTAIL.n198 185
R1358 VTAIL.n176 VTAIL.n175 185
R1359 VTAIL.n206 VTAIL.n205 185
R1360 VTAIL.n207 VTAIL.n174 185
R1361 VTAIL.n209 VTAIL.n208 185
R1362 VTAIL.n172 VTAIL.n171 185
R1363 VTAIL.n215 VTAIL.n214 185
R1364 VTAIL.n217 VTAIL.n216 185
R1365 VTAIL.n168 VTAIL.n167 185
R1366 VTAIL.n223 VTAIL.n222 185
R1367 VTAIL.n225 VTAIL.n224 185
R1368 VTAIL.n164 VTAIL.n163 185
R1369 VTAIL.n231 VTAIL.n230 185
R1370 VTAIL.n233 VTAIL.n232 185
R1371 VTAIL.n549 VTAIL.n548 185
R1372 VTAIL.n547 VTAIL.n546 185
R1373 VTAIL.n480 VTAIL.n479 185
R1374 VTAIL.n541 VTAIL.n540 185
R1375 VTAIL.n539 VTAIL.n538 185
R1376 VTAIL.n484 VTAIL.n483 185
R1377 VTAIL.n533 VTAIL.n532 185
R1378 VTAIL.n531 VTAIL.n530 185
R1379 VTAIL.n488 VTAIL.n487 185
R1380 VTAIL.n525 VTAIL.n524 185
R1381 VTAIL.n523 VTAIL.n490 185
R1382 VTAIL.n522 VTAIL.n521 185
R1383 VTAIL.n493 VTAIL.n491 185
R1384 VTAIL.n516 VTAIL.n515 185
R1385 VTAIL.n514 VTAIL.n513 185
R1386 VTAIL.n497 VTAIL.n496 185
R1387 VTAIL.n508 VTAIL.n507 185
R1388 VTAIL.n506 VTAIL.n505 185
R1389 VTAIL.n501 VTAIL.n500 185
R1390 VTAIL.n469 VTAIL.n468 185
R1391 VTAIL.n467 VTAIL.n466 185
R1392 VTAIL.n400 VTAIL.n399 185
R1393 VTAIL.n461 VTAIL.n460 185
R1394 VTAIL.n459 VTAIL.n458 185
R1395 VTAIL.n404 VTAIL.n403 185
R1396 VTAIL.n453 VTAIL.n452 185
R1397 VTAIL.n451 VTAIL.n450 185
R1398 VTAIL.n408 VTAIL.n407 185
R1399 VTAIL.n445 VTAIL.n444 185
R1400 VTAIL.n443 VTAIL.n410 185
R1401 VTAIL.n442 VTAIL.n441 185
R1402 VTAIL.n413 VTAIL.n411 185
R1403 VTAIL.n436 VTAIL.n435 185
R1404 VTAIL.n434 VTAIL.n433 185
R1405 VTAIL.n417 VTAIL.n416 185
R1406 VTAIL.n428 VTAIL.n427 185
R1407 VTAIL.n426 VTAIL.n425 185
R1408 VTAIL.n421 VTAIL.n420 185
R1409 VTAIL.n391 VTAIL.n390 185
R1410 VTAIL.n389 VTAIL.n388 185
R1411 VTAIL.n322 VTAIL.n321 185
R1412 VTAIL.n383 VTAIL.n382 185
R1413 VTAIL.n381 VTAIL.n380 185
R1414 VTAIL.n326 VTAIL.n325 185
R1415 VTAIL.n375 VTAIL.n374 185
R1416 VTAIL.n373 VTAIL.n372 185
R1417 VTAIL.n330 VTAIL.n329 185
R1418 VTAIL.n367 VTAIL.n366 185
R1419 VTAIL.n365 VTAIL.n332 185
R1420 VTAIL.n364 VTAIL.n363 185
R1421 VTAIL.n335 VTAIL.n333 185
R1422 VTAIL.n358 VTAIL.n357 185
R1423 VTAIL.n356 VTAIL.n355 185
R1424 VTAIL.n339 VTAIL.n338 185
R1425 VTAIL.n350 VTAIL.n349 185
R1426 VTAIL.n348 VTAIL.n347 185
R1427 VTAIL.n343 VTAIL.n342 185
R1428 VTAIL.n311 VTAIL.n310 185
R1429 VTAIL.n309 VTAIL.n308 185
R1430 VTAIL.n242 VTAIL.n241 185
R1431 VTAIL.n303 VTAIL.n302 185
R1432 VTAIL.n301 VTAIL.n300 185
R1433 VTAIL.n246 VTAIL.n245 185
R1434 VTAIL.n295 VTAIL.n294 185
R1435 VTAIL.n293 VTAIL.n292 185
R1436 VTAIL.n250 VTAIL.n249 185
R1437 VTAIL.n287 VTAIL.n286 185
R1438 VTAIL.n285 VTAIL.n252 185
R1439 VTAIL.n284 VTAIL.n283 185
R1440 VTAIL.n255 VTAIL.n253 185
R1441 VTAIL.n278 VTAIL.n277 185
R1442 VTAIL.n276 VTAIL.n275 185
R1443 VTAIL.n259 VTAIL.n258 185
R1444 VTAIL.n270 VTAIL.n269 185
R1445 VTAIL.n268 VTAIL.n267 185
R1446 VTAIL.n263 VTAIL.n262 185
R1447 VTAIL.n579 VTAIL.t12 149.524
R1448 VTAIL.n27 VTAIL.t14 149.524
R1449 VTAIL.n105 VTAIL.t5 149.524
R1450 VTAIL.n185 VTAIL.t2 149.524
R1451 VTAIL.n502 VTAIL.t15 149.524
R1452 VTAIL.n422 VTAIL.t6 149.524
R1453 VTAIL.n344 VTAIL.t9 149.524
R1454 VTAIL.n264 VTAIL.t10 149.524
R1455 VTAIL.n583 VTAIL.n577 104.615
R1456 VTAIL.n584 VTAIL.n583 104.615
R1457 VTAIL.n584 VTAIL.n573 104.615
R1458 VTAIL.n591 VTAIL.n573 104.615
R1459 VTAIL.n592 VTAIL.n591 104.615
R1460 VTAIL.n592 VTAIL.n569 104.615
R1461 VTAIL.n600 VTAIL.n569 104.615
R1462 VTAIL.n601 VTAIL.n600 104.615
R1463 VTAIL.n602 VTAIL.n601 104.615
R1464 VTAIL.n602 VTAIL.n565 104.615
R1465 VTAIL.n609 VTAIL.n565 104.615
R1466 VTAIL.n610 VTAIL.n609 104.615
R1467 VTAIL.n610 VTAIL.n561 104.615
R1468 VTAIL.n617 VTAIL.n561 104.615
R1469 VTAIL.n618 VTAIL.n617 104.615
R1470 VTAIL.n618 VTAIL.n557 104.615
R1471 VTAIL.n625 VTAIL.n557 104.615
R1472 VTAIL.n626 VTAIL.n625 104.615
R1473 VTAIL.n31 VTAIL.n25 104.615
R1474 VTAIL.n32 VTAIL.n31 104.615
R1475 VTAIL.n32 VTAIL.n21 104.615
R1476 VTAIL.n39 VTAIL.n21 104.615
R1477 VTAIL.n40 VTAIL.n39 104.615
R1478 VTAIL.n40 VTAIL.n17 104.615
R1479 VTAIL.n48 VTAIL.n17 104.615
R1480 VTAIL.n49 VTAIL.n48 104.615
R1481 VTAIL.n50 VTAIL.n49 104.615
R1482 VTAIL.n50 VTAIL.n13 104.615
R1483 VTAIL.n57 VTAIL.n13 104.615
R1484 VTAIL.n58 VTAIL.n57 104.615
R1485 VTAIL.n58 VTAIL.n9 104.615
R1486 VTAIL.n65 VTAIL.n9 104.615
R1487 VTAIL.n66 VTAIL.n65 104.615
R1488 VTAIL.n66 VTAIL.n5 104.615
R1489 VTAIL.n73 VTAIL.n5 104.615
R1490 VTAIL.n74 VTAIL.n73 104.615
R1491 VTAIL.n109 VTAIL.n103 104.615
R1492 VTAIL.n110 VTAIL.n109 104.615
R1493 VTAIL.n110 VTAIL.n99 104.615
R1494 VTAIL.n117 VTAIL.n99 104.615
R1495 VTAIL.n118 VTAIL.n117 104.615
R1496 VTAIL.n118 VTAIL.n95 104.615
R1497 VTAIL.n126 VTAIL.n95 104.615
R1498 VTAIL.n127 VTAIL.n126 104.615
R1499 VTAIL.n128 VTAIL.n127 104.615
R1500 VTAIL.n128 VTAIL.n91 104.615
R1501 VTAIL.n135 VTAIL.n91 104.615
R1502 VTAIL.n136 VTAIL.n135 104.615
R1503 VTAIL.n136 VTAIL.n87 104.615
R1504 VTAIL.n143 VTAIL.n87 104.615
R1505 VTAIL.n144 VTAIL.n143 104.615
R1506 VTAIL.n144 VTAIL.n83 104.615
R1507 VTAIL.n151 VTAIL.n83 104.615
R1508 VTAIL.n152 VTAIL.n151 104.615
R1509 VTAIL.n189 VTAIL.n183 104.615
R1510 VTAIL.n190 VTAIL.n189 104.615
R1511 VTAIL.n190 VTAIL.n179 104.615
R1512 VTAIL.n197 VTAIL.n179 104.615
R1513 VTAIL.n198 VTAIL.n197 104.615
R1514 VTAIL.n198 VTAIL.n175 104.615
R1515 VTAIL.n206 VTAIL.n175 104.615
R1516 VTAIL.n207 VTAIL.n206 104.615
R1517 VTAIL.n208 VTAIL.n207 104.615
R1518 VTAIL.n208 VTAIL.n171 104.615
R1519 VTAIL.n215 VTAIL.n171 104.615
R1520 VTAIL.n216 VTAIL.n215 104.615
R1521 VTAIL.n216 VTAIL.n167 104.615
R1522 VTAIL.n223 VTAIL.n167 104.615
R1523 VTAIL.n224 VTAIL.n223 104.615
R1524 VTAIL.n224 VTAIL.n163 104.615
R1525 VTAIL.n231 VTAIL.n163 104.615
R1526 VTAIL.n232 VTAIL.n231 104.615
R1527 VTAIL.n548 VTAIL.n547 104.615
R1528 VTAIL.n547 VTAIL.n479 104.615
R1529 VTAIL.n540 VTAIL.n479 104.615
R1530 VTAIL.n540 VTAIL.n539 104.615
R1531 VTAIL.n539 VTAIL.n483 104.615
R1532 VTAIL.n532 VTAIL.n483 104.615
R1533 VTAIL.n532 VTAIL.n531 104.615
R1534 VTAIL.n531 VTAIL.n487 104.615
R1535 VTAIL.n524 VTAIL.n487 104.615
R1536 VTAIL.n524 VTAIL.n523 104.615
R1537 VTAIL.n523 VTAIL.n522 104.615
R1538 VTAIL.n522 VTAIL.n491 104.615
R1539 VTAIL.n515 VTAIL.n491 104.615
R1540 VTAIL.n515 VTAIL.n514 104.615
R1541 VTAIL.n514 VTAIL.n496 104.615
R1542 VTAIL.n507 VTAIL.n496 104.615
R1543 VTAIL.n507 VTAIL.n506 104.615
R1544 VTAIL.n506 VTAIL.n500 104.615
R1545 VTAIL.n468 VTAIL.n467 104.615
R1546 VTAIL.n467 VTAIL.n399 104.615
R1547 VTAIL.n460 VTAIL.n399 104.615
R1548 VTAIL.n460 VTAIL.n459 104.615
R1549 VTAIL.n459 VTAIL.n403 104.615
R1550 VTAIL.n452 VTAIL.n403 104.615
R1551 VTAIL.n452 VTAIL.n451 104.615
R1552 VTAIL.n451 VTAIL.n407 104.615
R1553 VTAIL.n444 VTAIL.n407 104.615
R1554 VTAIL.n444 VTAIL.n443 104.615
R1555 VTAIL.n443 VTAIL.n442 104.615
R1556 VTAIL.n442 VTAIL.n411 104.615
R1557 VTAIL.n435 VTAIL.n411 104.615
R1558 VTAIL.n435 VTAIL.n434 104.615
R1559 VTAIL.n434 VTAIL.n416 104.615
R1560 VTAIL.n427 VTAIL.n416 104.615
R1561 VTAIL.n427 VTAIL.n426 104.615
R1562 VTAIL.n426 VTAIL.n420 104.615
R1563 VTAIL.n390 VTAIL.n389 104.615
R1564 VTAIL.n389 VTAIL.n321 104.615
R1565 VTAIL.n382 VTAIL.n321 104.615
R1566 VTAIL.n382 VTAIL.n381 104.615
R1567 VTAIL.n381 VTAIL.n325 104.615
R1568 VTAIL.n374 VTAIL.n325 104.615
R1569 VTAIL.n374 VTAIL.n373 104.615
R1570 VTAIL.n373 VTAIL.n329 104.615
R1571 VTAIL.n366 VTAIL.n329 104.615
R1572 VTAIL.n366 VTAIL.n365 104.615
R1573 VTAIL.n365 VTAIL.n364 104.615
R1574 VTAIL.n364 VTAIL.n333 104.615
R1575 VTAIL.n357 VTAIL.n333 104.615
R1576 VTAIL.n357 VTAIL.n356 104.615
R1577 VTAIL.n356 VTAIL.n338 104.615
R1578 VTAIL.n349 VTAIL.n338 104.615
R1579 VTAIL.n349 VTAIL.n348 104.615
R1580 VTAIL.n348 VTAIL.n342 104.615
R1581 VTAIL.n310 VTAIL.n309 104.615
R1582 VTAIL.n309 VTAIL.n241 104.615
R1583 VTAIL.n302 VTAIL.n241 104.615
R1584 VTAIL.n302 VTAIL.n301 104.615
R1585 VTAIL.n301 VTAIL.n245 104.615
R1586 VTAIL.n294 VTAIL.n245 104.615
R1587 VTAIL.n294 VTAIL.n293 104.615
R1588 VTAIL.n293 VTAIL.n249 104.615
R1589 VTAIL.n286 VTAIL.n249 104.615
R1590 VTAIL.n286 VTAIL.n285 104.615
R1591 VTAIL.n285 VTAIL.n284 104.615
R1592 VTAIL.n284 VTAIL.n253 104.615
R1593 VTAIL.n277 VTAIL.n253 104.615
R1594 VTAIL.n277 VTAIL.n276 104.615
R1595 VTAIL.n276 VTAIL.n258 104.615
R1596 VTAIL.n269 VTAIL.n258 104.615
R1597 VTAIL.n269 VTAIL.n268 104.615
R1598 VTAIL.n268 VTAIL.n262 104.615
R1599 VTAIL.t12 VTAIL.n577 52.3082
R1600 VTAIL.t14 VTAIL.n25 52.3082
R1601 VTAIL.t5 VTAIL.n103 52.3082
R1602 VTAIL.t2 VTAIL.n183 52.3082
R1603 VTAIL.t15 VTAIL.n500 52.3082
R1604 VTAIL.t6 VTAIL.n420 52.3082
R1605 VTAIL.t9 VTAIL.n342 52.3082
R1606 VTAIL.t10 VTAIL.n262 52.3082
R1607 VTAIL.n475 VTAIL.n474 43.9736
R1608 VTAIL.n317 VTAIL.n316 43.9736
R1609 VTAIL.n1 VTAIL.n0 43.9736
R1610 VTAIL.n159 VTAIL.n158 43.9736
R1611 VTAIL.n631 VTAIL.n630 31.4096
R1612 VTAIL.n79 VTAIL.n78 31.4096
R1613 VTAIL.n157 VTAIL.n156 31.4096
R1614 VTAIL.n237 VTAIL.n236 31.4096
R1615 VTAIL.n553 VTAIL.n552 31.4096
R1616 VTAIL.n473 VTAIL.n472 31.4096
R1617 VTAIL.n395 VTAIL.n394 31.4096
R1618 VTAIL.n315 VTAIL.n314 31.4096
R1619 VTAIL.n631 VTAIL.n553 25.3238
R1620 VTAIL.n315 VTAIL.n237 25.3238
R1621 VTAIL.n603 VTAIL.n568 13.1884
R1622 VTAIL.n51 VTAIL.n16 13.1884
R1623 VTAIL.n129 VTAIL.n94 13.1884
R1624 VTAIL.n209 VTAIL.n174 13.1884
R1625 VTAIL.n525 VTAIL.n490 13.1884
R1626 VTAIL.n445 VTAIL.n410 13.1884
R1627 VTAIL.n367 VTAIL.n332 13.1884
R1628 VTAIL.n287 VTAIL.n252 13.1884
R1629 VTAIL.n599 VTAIL.n598 12.8005
R1630 VTAIL.n604 VTAIL.n566 12.8005
R1631 VTAIL.n47 VTAIL.n46 12.8005
R1632 VTAIL.n52 VTAIL.n14 12.8005
R1633 VTAIL.n125 VTAIL.n124 12.8005
R1634 VTAIL.n130 VTAIL.n92 12.8005
R1635 VTAIL.n205 VTAIL.n204 12.8005
R1636 VTAIL.n210 VTAIL.n172 12.8005
R1637 VTAIL.n526 VTAIL.n488 12.8005
R1638 VTAIL.n521 VTAIL.n492 12.8005
R1639 VTAIL.n446 VTAIL.n408 12.8005
R1640 VTAIL.n441 VTAIL.n412 12.8005
R1641 VTAIL.n368 VTAIL.n330 12.8005
R1642 VTAIL.n363 VTAIL.n334 12.8005
R1643 VTAIL.n288 VTAIL.n250 12.8005
R1644 VTAIL.n283 VTAIL.n254 12.8005
R1645 VTAIL.n597 VTAIL.n570 12.0247
R1646 VTAIL.n608 VTAIL.n607 12.0247
R1647 VTAIL.n45 VTAIL.n18 12.0247
R1648 VTAIL.n56 VTAIL.n55 12.0247
R1649 VTAIL.n123 VTAIL.n96 12.0247
R1650 VTAIL.n134 VTAIL.n133 12.0247
R1651 VTAIL.n203 VTAIL.n176 12.0247
R1652 VTAIL.n214 VTAIL.n213 12.0247
R1653 VTAIL.n530 VTAIL.n529 12.0247
R1654 VTAIL.n520 VTAIL.n493 12.0247
R1655 VTAIL.n450 VTAIL.n449 12.0247
R1656 VTAIL.n440 VTAIL.n413 12.0247
R1657 VTAIL.n372 VTAIL.n371 12.0247
R1658 VTAIL.n362 VTAIL.n335 12.0247
R1659 VTAIL.n292 VTAIL.n291 12.0247
R1660 VTAIL.n282 VTAIL.n255 12.0247
R1661 VTAIL.n594 VTAIL.n593 11.249
R1662 VTAIL.n611 VTAIL.n564 11.249
R1663 VTAIL.n42 VTAIL.n41 11.249
R1664 VTAIL.n59 VTAIL.n12 11.249
R1665 VTAIL.n120 VTAIL.n119 11.249
R1666 VTAIL.n137 VTAIL.n90 11.249
R1667 VTAIL.n200 VTAIL.n199 11.249
R1668 VTAIL.n217 VTAIL.n170 11.249
R1669 VTAIL.n533 VTAIL.n486 11.249
R1670 VTAIL.n517 VTAIL.n516 11.249
R1671 VTAIL.n453 VTAIL.n406 11.249
R1672 VTAIL.n437 VTAIL.n436 11.249
R1673 VTAIL.n375 VTAIL.n328 11.249
R1674 VTAIL.n359 VTAIL.n358 11.249
R1675 VTAIL.n295 VTAIL.n248 11.249
R1676 VTAIL.n279 VTAIL.n278 11.249
R1677 VTAIL.n590 VTAIL.n572 10.4732
R1678 VTAIL.n612 VTAIL.n562 10.4732
R1679 VTAIL.n38 VTAIL.n20 10.4732
R1680 VTAIL.n60 VTAIL.n10 10.4732
R1681 VTAIL.n116 VTAIL.n98 10.4732
R1682 VTAIL.n138 VTAIL.n88 10.4732
R1683 VTAIL.n196 VTAIL.n178 10.4732
R1684 VTAIL.n218 VTAIL.n168 10.4732
R1685 VTAIL.n534 VTAIL.n484 10.4732
R1686 VTAIL.n513 VTAIL.n495 10.4732
R1687 VTAIL.n454 VTAIL.n404 10.4732
R1688 VTAIL.n433 VTAIL.n415 10.4732
R1689 VTAIL.n376 VTAIL.n326 10.4732
R1690 VTAIL.n355 VTAIL.n337 10.4732
R1691 VTAIL.n296 VTAIL.n246 10.4732
R1692 VTAIL.n275 VTAIL.n257 10.4732
R1693 VTAIL.n579 VTAIL.n578 10.2747
R1694 VTAIL.n27 VTAIL.n26 10.2747
R1695 VTAIL.n105 VTAIL.n104 10.2747
R1696 VTAIL.n185 VTAIL.n184 10.2747
R1697 VTAIL.n502 VTAIL.n501 10.2747
R1698 VTAIL.n422 VTAIL.n421 10.2747
R1699 VTAIL.n344 VTAIL.n343 10.2747
R1700 VTAIL.n264 VTAIL.n263 10.2747
R1701 VTAIL.n589 VTAIL.n574 9.69747
R1702 VTAIL.n616 VTAIL.n615 9.69747
R1703 VTAIL.n37 VTAIL.n22 9.69747
R1704 VTAIL.n64 VTAIL.n63 9.69747
R1705 VTAIL.n115 VTAIL.n100 9.69747
R1706 VTAIL.n142 VTAIL.n141 9.69747
R1707 VTAIL.n195 VTAIL.n180 9.69747
R1708 VTAIL.n222 VTAIL.n221 9.69747
R1709 VTAIL.n538 VTAIL.n537 9.69747
R1710 VTAIL.n512 VTAIL.n497 9.69747
R1711 VTAIL.n458 VTAIL.n457 9.69747
R1712 VTAIL.n432 VTAIL.n417 9.69747
R1713 VTAIL.n380 VTAIL.n379 9.69747
R1714 VTAIL.n354 VTAIL.n339 9.69747
R1715 VTAIL.n300 VTAIL.n299 9.69747
R1716 VTAIL.n274 VTAIL.n259 9.69747
R1717 VTAIL.n630 VTAIL.n629 9.45567
R1718 VTAIL.n78 VTAIL.n77 9.45567
R1719 VTAIL.n156 VTAIL.n155 9.45567
R1720 VTAIL.n236 VTAIL.n235 9.45567
R1721 VTAIL.n552 VTAIL.n551 9.45567
R1722 VTAIL.n472 VTAIL.n471 9.45567
R1723 VTAIL.n394 VTAIL.n393 9.45567
R1724 VTAIL.n314 VTAIL.n313 9.45567
R1725 VTAIL.n556 VTAIL.n555 9.3005
R1726 VTAIL.n629 VTAIL.n628 9.3005
R1727 VTAIL.n621 VTAIL.n620 9.3005
R1728 VTAIL.n560 VTAIL.n559 9.3005
R1729 VTAIL.n615 VTAIL.n614 9.3005
R1730 VTAIL.n613 VTAIL.n612 9.3005
R1731 VTAIL.n564 VTAIL.n563 9.3005
R1732 VTAIL.n607 VTAIL.n606 9.3005
R1733 VTAIL.n605 VTAIL.n604 9.3005
R1734 VTAIL.n581 VTAIL.n580 9.3005
R1735 VTAIL.n576 VTAIL.n575 9.3005
R1736 VTAIL.n587 VTAIL.n586 9.3005
R1737 VTAIL.n589 VTAIL.n588 9.3005
R1738 VTAIL.n572 VTAIL.n571 9.3005
R1739 VTAIL.n595 VTAIL.n594 9.3005
R1740 VTAIL.n597 VTAIL.n596 9.3005
R1741 VTAIL.n598 VTAIL.n567 9.3005
R1742 VTAIL.n623 VTAIL.n622 9.3005
R1743 VTAIL.n4 VTAIL.n3 9.3005
R1744 VTAIL.n77 VTAIL.n76 9.3005
R1745 VTAIL.n69 VTAIL.n68 9.3005
R1746 VTAIL.n8 VTAIL.n7 9.3005
R1747 VTAIL.n63 VTAIL.n62 9.3005
R1748 VTAIL.n61 VTAIL.n60 9.3005
R1749 VTAIL.n12 VTAIL.n11 9.3005
R1750 VTAIL.n55 VTAIL.n54 9.3005
R1751 VTAIL.n53 VTAIL.n52 9.3005
R1752 VTAIL.n29 VTAIL.n28 9.3005
R1753 VTAIL.n24 VTAIL.n23 9.3005
R1754 VTAIL.n35 VTAIL.n34 9.3005
R1755 VTAIL.n37 VTAIL.n36 9.3005
R1756 VTAIL.n20 VTAIL.n19 9.3005
R1757 VTAIL.n43 VTAIL.n42 9.3005
R1758 VTAIL.n45 VTAIL.n44 9.3005
R1759 VTAIL.n46 VTAIL.n15 9.3005
R1760 VTAIL.n71 VTAIL.n70 9.3005
R1761 VTAIL.n82 VTAIL.n81 9.3005
R1762 VTAIL.n155 VTAIL.n154 9.3005
R1763 VTAIL.n147 VTAIL.n146 9.3005
R1764 VTAIL.n86 VTAIL.n85 9.3005
R1765 VTAIL.n141 VTAIL.n140 9.3005
R1766 VTAIL.n139 VTAIL.n138 9.3005
R1767 VTAIL.n90 VTAIL.n89 9.3005
R1768 VTAIL.n133 VTAIL.n132 9.3005
R1769 VTAIL.n131 VTAIL.n130 9.3005
R1770 VTAIL.n107 VTAIL.n106 9.3005
R1771 VTAIL.n102 VTAIL.n101 9.3005
R1772 VTAIL.n113 VTAIL.n112 9.3005
R1773 VTAIL.n115 VTAIL.n114 9.3005
R1774 VTAIL.n98 VTAIL.n97 9.3005
R1775 VTAIL.n121 VTAIL.n120 9.3005
R1776 VTAIL.n123 VTAIL.n122 9.3005
R1777 VTAIL.n124 VTAIL.n93 9.3005
R1778 VTAIL.n149 VTAIL.n148 9.3005
R1779 VTAIL.n162 VTAIL.n161 9.3005
R1780 VTAIL.n235 VTAIL.n234 9.3005
R1781 VTAIL.n227 VTAIL.n226 9.3005
R1782 VTAIL.n166 VTAIL.n165 9.3005
R1783 VTAIL.n221 VTAIL.n220 9.3005
R1784 VTAIL.n219 VTAIL.n218 9.3005
R1785 VTAIL.n170 VTAIL.n169 9.3005
R1786 VTAIL.n213 VTAIL.n212 9.3005
R1787 VTAIL.n211 VTAIL.n210 9.3005
R1788 VTAIL.n187 VTAIL.n186 9.3005
R1789 VTAIL.n182 VTAIL.n181 9.3005
R1790 VTAIL.n193 VTAIL.n192 9.3005
R1791 VTAIL.n195 VTAIL.n194 9.3005
R1792 VTAIL.n178 VTAIL.n177 9.3005
R1793 VTAIL.n201 VTAIL.n200 9.3005
R1794 VTAIL.n203 VTAIL.n202 9.3005
R1795 VTAIL.n204 VTAIL.n173 9.3005
R1796 VTAIL.n229 VTAIL.n228 9.3005
R1797 VTAIL.n478 VTAIL.n477 9.3005
R1798 VTAIL.n545 VTAIL.n544 9.3005
R1799 VTAIL.n543 VTAIL.n542 9.3005
R1800 VTAIL.n482 VTAIL.n481 9.3005
R1801 VTAIL.n537 VTAIL.n536 9.3005
R1802 VTAIL.n535 VTAIL.n534 9.3005
R1803 VTAIL.n486 VTAIL.n485 9.3005
R1804 VTAIL.n529 VTAIL.n528 9.3005
R1805 VTAIL.n527 VTAIL.n526 9.3005
R1806 VTAIL.n492 VTAIL.n489 9.3005
R1807 VTAIL.n520 VTAIL.n519 9.3005
R1808 VTAIL.n518 VTAIL.n517 9.3005
R1809 VTAIL.n495 VTAIL.n494 9.3005
R1810 VTAIL.n512 VTAIL.n511 9.3005
R1811 VTAIL.n510 VTAIL.n509 9.3005
R1812 VTAIL.n499 VTAIL.n498 9.3005
R1813 VTAIL.n504 VTAIL.n503 9.3005
R1814 VTAIL.n551 VTAIL.n550 9.3005
R1815 VTAIL.n424 VTAIL.n423 9.3005
R1816 VTAIL.n419 VTAIL.n418 9.3005
R1817 VTAIL.n430 VTAIL.n429 9.3005
R1818 VTAIL.n432 VTAIL.n431 9.3005
R1819 VTAIL.n415 VTAIL.n414 9.3005
R1820 VTAIL.n438 VTAIL.n437 9.3005
R1821 VTAIL.n440 VTAIL.n439 9.3005
R1822 VTAIL.n412 VTAIL.n409 9.3005
R1823 VTAIL.n471 VTAIL.n470 9.3005
R1824 VTAIL.n398 VTAIL.n397 9.3005
R1825 VTAIL.n465 VTAIL.n464 9.3005
R1826 VTAIL.n463 VTAIL.n462 9.3005
R1827 VTAIL.n402 VTAIL.n401 9.3005
R1828 VTAIL.n457 VTAIL.n456 9.3005
R1829 VTAIL.n455 VTAIL.n454 9.3005
R1830 VTAIL.n406 VTAIL.n405 9.3005
R1831 VTAIL.n449 VTAIL.n448 9.3005
R1832 VTAIL.n447 VTAIL.n446 9.3005
R1833 VTAIL.n346 VTAIL.n345 9.3005
R1834 VTAIL.n341 VTAIL.n340 9.3005
R1835 VTAIL.n352 VTAIL.n351 9.3005
R1836 VTAIL.n354 VTAIL.n353 9.3005
R1837 VTAIL.n337 VTAIL.n336 9.3005
R1838 VTAIL.n360 VTAIL.n359 9.3005
R1839 VTAIL.n362 VTAIL.n361 9.3005
R1840 VTAIL.n334 VTAIL.n331 9.3005
R1841 VTAIL.n393 VTAIL.n392 9.3005
R1842 VTAIL.n320 VTAIL.n319 9.3005
R1843 VTAIL.n387 VTAIL.n386 9.3005
R1844 VTAIL.n385 VTAIL.n384 9.3005
R1845 VTAIL.n324 VTAIL.n323 9.3005
R1846 VTAIL.n379 VTAIL.n378 9.3005
R1847 VTAIL.n377 VTAIL.n376 9.3005
R1848 VTAIL.n328 VTAIL.n327 9.3005
R1849 VTAIL.n371 VTAIL.n370 9.3005
R1850 VTAIL.n369 VTAIL.n368 9.3005
R1851 VTAIL.n266 VTAIL.n265 9.3005
R1852 VTAIL.n261 VTAIL.n260 9.3005
R1853 VTAIL.n272 VTAIL.n271 9.3005
R1854 VTAIL.n274 VTAIL.n273 9.3005
R1855 VTAIL.n257 VTAIL.n256 9.3005
R1856 VTAIL.n280 VTAIL.n279 9.3005
R1857 VTAIL.n282 VTAIL.n281 9.3005
R1858 VTAIL.n254 VTAIL.n251 9.3005
R1859 VTAIL.n313 VTAIL.n312 9.3005
R1860 VTAIL.n240 VTAIL.n239 9.3005
R1861 VTAIL.n307 VTAIL.n306 9.3005
R1862 VTAIL.n305 VTAIL.n304 9.3005
R1863 VTAIL.n244 VTAIL.n243 9.3005
R1864 VTAIL.n299 VTAIL.n298 9.3005
R1865 VTAIL.n297 VTAIL.n296 9.3005
R1866 VTAIL.n248 VTAIL.n247 9.3005
R1867 VTAIL.n291 VTAIL.n290 9.3005
R1868 VTAIL.n289 VTAIL.n288 9.3005
R1869 VTAIL.n586 VTAIL.n585 8.92171
R1870 VTAIL.n619 VTAIL.n560 8.92171
R1871 VTAIL.n34 VTAIL.n33 8.92171
R1872 VTAIL.n67 VTAIL.n8 8.92171
R1873 VTAIL.n112 VTAIL.n111 8.92171
R1874 VTAIL.n145 VTAIL.n86 8.92171
R1875 VTAIL.n192 VTAIL.n191 8.92171
R1876 VTAIL.n225 VTAIL.n166 8.92171
R1877 VTAIL.n541 VTAIL.n482 8.92171
R1878 VTAIL.n509 VTAIL.n508 8.92171
R1879 VTAIL.n461 VTAIL.n402 8.92171
R1880 VTAIL.n429 VTAIL.n428 8.92171
R1881 VTAIL.n383 VTAIL.n324 8.92171
R1882 VTAIL.n351 VTAIL.n350 8.92171
R1883 VTAIL.n303 VTAIL.n244 8.92171
R1884 VTAIL.n271 VTAIL.n270 8.92171
R1885 VTAIL.n582 VTAIL.n576 8.14595
R1886 VTAIL.n620 VTAIL.n558 8.14595
R1887 VTAIL.n630 VTAIL.n554 8.14595
R1888 VTAIL.n30 VTAIL.n24 8.14595
R1889 VTAIL.n68 VTAIL.n6 8.14595
R1890 VTAIL.n78 VTAIL.n2 8.14595
R1891 VTAIL.n108 VTAIL.n102 8.14595
R1892 VTAIL.n146 VTAIL.n84 8.14595
R1893 VTAIL.n156 VTAIL.n80 8.14595
R1894 VTAIL.n188 VTAIL.n182 8.14595
R1895 VTAIL.n226 VTAIL.n164 8.14595
R1896 VTAIL.n236 VTAIL.n160 8.14595
R1897 VTAIL.n552 VTAIL.n476 8.14595
R1898 VTAIL.n542 VTAIL.n480 8.14595
R1899 VTAIL.n505 VTAIL.n499 8.14595
R1900 VTAIL.n472 VTAIL.n396 8.14595
R1901 VTAIL.n462 VTAIL.n400 8.14595
R1902 VTAIL.n425 VTAIL.n419 8.14595
R1903 VTAIL.n394 VTAIL.n318 8.14595
R1904 VTAIL.n384 VTAIL.n322 8.14595
R1905 VTAIL.n347 VTAIL.n341 8.14595
R1906 VTAIL.n314 VTAIL.n238 8.14595
R1907 VTAIL.n304 VTAIL.n242 8.14595
R1908 VTAIL.n267 VTAIL.n261 8.14595
R1909 VTAIL.n581 VTAIL.n578 7.3702
R1910 VTAIL.n624 VTAIL.n623 7.3702
R1911 VTAIL.n628 VTAIL.n627 7.3702
R1912 VTAIL.n29 VTAIL.n26 7.3702
R1913 VTAIL.n72 VTAIL.n71 7.3702
R1914 VTAIL.n76 VTAIL.n75 7.3702
R1915 VTAIL.n107 VTAIL.n104 7.3702
R1916 VTAIL.n150 VTAIL.n149 7.3702
R1917 VTAIL.n154 VTAIL.n153 7.3702
R1918 VTAIL.n187 VTAIL.n184 7.3702
R1919 VTAIL.n230 VTAIL.n229 7.3702
R1920 VTAIL.n234 VTAIL.n233 7.3702
R1921 VTAIL.n550 VTAIL.n549 7.3702
R1922 VTAIL.n546 VTAIL.n545 7.3702
R1923 VTAIL.n504 VTAIL.n501 7.3702
R1924 VTAIL.n470 VTAIL.n469 7.3702
R1925 VTAIL.n466 VTAIL.n465 7.3702
R1926 VTAIL.n424 VTAIL.n421 7.3702
R1927 VTAIL.n392 VTAIL.n391 7.3702
R1928 VTAIL.n388 VTAIL.n387 7.3702
R1929 VTAIL.n346 VTAIL.n343 7.3702
R1930 VTAIL.n312 VTAIL.n311 7.3702
R1931 VTAIL.n308 VTAIL.n307 7.3702
R1932 VTAIL.n266 VTAIL.n263 7.3702
R1933 VTAIL.n624 VTAIL.n556 6.59444
R1934 VTAIL.n627 VTAIL.n556 6.59444
R1935 VTAIL.n72 VTAIL.n4 6.59444
R1936 VTAIL.n75 VTAIL.n4 6.59444
R1937 VTAIL.n150 VTAIL.n82 6.59444
R1938 VTAIL.n153 VTAIL.n82 6.59444
R1939 VTAIL.n230 VTAIL.n162 6.59444
R1940 VTAIL.n233 VTAIL.n162 6.59444
R1941 VTAIL.n549 VTAIL.n478 6.59444
R1942 VTAIL.n546 VTAIL.n478 6.59444
R1943 VTAIL.n469 VTAIL.n398 6.59444
R1944 VTAIL.n466 VTAIL.n398 6.59444
R1945 VTAIL.n391 VTAIL.n320 6.59444
R1946 VTAIL.n388 VTAIL.n320 6.59444
R1947 VTAIL.n311 VTAIL.n240 6.59444
R1948 VTAIL.n308 VTAIL.n240 6.59444
R1949 VTAIL.n582 VTAIL.n581 5.81868
R1950 VTAIL.n623 VTAIL.n558 5.81868
R1951 VTAIL.n628 VTAIL.n554 5.81868
R1952 VTAIL.n30 VTAIL.n29 5.81868
R1953 VTAIL.n71 VTAIL.n6 5.81868
R1954 VTAIL.n76 VTAIL.n2 5.81868
R1955 VTAIL.n108 VTAIL.n107 5.81868
R1956 VTAIL.n149 VTAIL.n84 5.81868
R1957 VTAIL.n154 VTAIL.n80 5.81868
R1958 VTAIL.n188 VTAIL.n187 5.81868
R1959 VTAIL.n229 VTAIL.n164 5.81868
R1960 VTAIL.n234 VTAIL.n160 5.81868
R1961 VTAIL.n550 VTAIL.n476 5.81868
R1962 VTAIL.n545 VTAIL.n480 5.81868
R1963 VTAIL.n505 VTAIL.n504 5.81868
R1964 VTAIL.n470 VTAIL.n396 5.81868
R1965 VTAIL.n465 VTAIL.n400 5.81868
R1966 VTAIL.n425 VTAIL.n424 5.81868
R1967 VTAIL.n392 VTAIL.n318 5.81868
R1968 VTAIL.n387 VTAIL.n322 5.81868
R1969 VTAIL.n347 VTAIL.n346 5.81868
R1970 VTAIL.n312 VTAIL.n238 5.81868
R1971 VTAIL.n307 VTAIL.n242 5.81868
R1972 VTAIL.n267 VTAIL.n266 5.81868
R1973 VTAIL.n585 VTAIL.n576 5.04292
R1974 VTAIL.n620 VTAIL.n619 5.04292
R1975 VTAIL.n33 VTAIL.n24 5.04292
R1976 VTAIL.n68 VTAIL.n67 5.04292
R1977 VTAIL.n111 VTAIL.n102 5.04292
R1978 VTAIL.n146 VTAIL.n145 5.04292
R1979 VTAIL.n191 VTAIL.n182 5.04292
R1980 VTAIL.n226 VTAIL.n225 5.04292
R1981 VTAIL.n542 VTAIL.n541 5.04292
R1982 VTAIL.n508 VTAIL.n499 5.04292
R1983 VTAIL.n462 VTAIL.n461 5.04292
R1984 VTAIL.n428 VTAIL.n419 5.04292
R1985 VTAIL.n384 VTAIL.n383 5.04292
R1986 VTAIL.n350 VTAIL.n341 5.04292
R1987 VTAIL.n304 VTAIL.n303 5.04292
R1988 VTAIL.n270 VTAIL.n261 5.04292
R1989 VTAIL.n586 VTAIL.n574 4.26717
R1990 VTAIL.n616 VTAIL.n560 4.26717
R1991 VTAIL.n34 VTAIL.n22 4.26717
R1992 VTAIL.n64 VTAIL.n8 4.26717
R1993 VTAIL.n112 VTAIL.n100 4.26717
R1994 VTAIL.n142 VTAIL.n86 4.26717
R1995 VTAIL.n192 VTAIL.n180 4.26717
R1996 VTAIL.n222 VTAIL.n166 4.26717
R1997 VTAIL.n538 VTAIL.n482 4.26717
R1998 VTAIL.n509 VTAIL.n497 4.26717
R1999 VTAIL.n458 VTAIL.n402 4.26717
R2000 VTAIL.n429 VTAIL.n417 4.26717
R2001 VTAIL.n380 VTAIL.n324 4.26717
R2002 VTAIL.n351 VTAIL.n339 4.26717
R2003 VTAIL.n300 VTAIL.n244 4.26717
R2004 VTAIL.n271 VTAIL.n259 4.26717
R2005 VTAIL.n590 VTAIL.n589 3.49141
R2006 VTAIL.n615 VTAIL.n562 3.49141
R2007 VTAIL.n38 VTAIL.n37 3.49141
R2008 VTAIL.n63 VTAIL.n10 3.49141
R2009 VTAIL.n116 VTAIL.n115 3.49141
R2010 VTAIL.n141 VTAIL.n88 3.49141
R2011 VTAIL.n196 VTAIL.n195 3.49141
R2012 VTAIL.n221 VTAIL.n168 3.49141
R2013 VTAIL.n537 VTAIL.n484 3.49141
R2014 VTAIL.n513 VTAIL.n512 3.49141
R2015 VTAIL.n457 VTAIL.n404 3.49141
R2016 VTAIL.n433 VTAIL.n432 3.49141
R2017 VTAIL.n379 VTAIL.n326 3.49141
R2018 VTAIL.n355 VTAIL.n354 3.49141
R2019 VTAIL.n299 VTAIL.n246 3.49141
R2020 VTAIL.n275 VTAIL.n274 3.49141
R2021 VTAIL.n580 VTAIL.n579 2.84303
R2022 VTAIL.n28 VTAIL.n27 2.84303
R2023 VTAIL.n106 VTAIL.n105 2.84303
R2024 VTAIL.n186 VTAIL.n185 2.84303
R2025 VTAIL.n423 VTAIL.n422 2.84303
R2026 VTAIL.n345 VTAIL.n344 2.84303
R2027 VTAIL.n265 VTAIL.n264 2.84303
R2028 VTAIL.n503 VTAIL.n502 2.84303
R2029 VTAIL.n593 VTAIL.n572 2.71565
R2030 VTAIL.n612 VTAIL.n611 2.71565
R2031 VTAIL.n41 VTAIL.n20 2.71565
R2032 VTAIL.n60 VTAIL.n59 2.71565
R2033 VTAIL.n119 VTAIL.n98 2.71565
R2034 VTAIL.n138 VTAIL.n137 2.71565
R2035 VTAIL.n199 VTAIL.n178 2.71565
R2036 VTAIL.n218 VTAIL.n217 2.71565
R2037 VTAIL.n534 VTAIL.n533 2.71565
R2038 VTAIL.n516 VTAIL.n495 2.71565
R2039 VTAIL.n454 VTAIL.n453 2.71565
R2040 VTAIL.n436 VTAIL.n415 2.71565
R2041 VTAIL.n376 VTAIL.n375 2.71565
R2042 VTAIL.n358 VTAIL.n337 2.71565
R2043 VTAIL.n296 VTAIL.n295 2.71565
R2044 VTAIL.n278 VTAIL.n257 2.71565
R2045 VTAIL.n594 VTAIL.n570 1.93989
R2046 VTAIL.n608 VTAIL.n564 1.93989
R2047 VTAIL.n42 VTAIL.n18 1.93989
R2048 VTAIL.n56 VTAIL.n12 1.93989
R2049 VTAIL.n120 VTAIL.n96 1.93989
R2050 VTAIL.n134 VTAIL.n90 1.93989
R2051 VTAIL.n200 VTAIL.n176 1.93989
R2052 VTAIL.n214 VTAIL.n170 1.93989
R2053 VTAIL.n530 VTAIL.n486 1.93989
R2054 VTAIL.n517 VTAIL.n493 1.93989
R2055 VTAIL.n450 VTAIL.n406 1.93989
R2056 VTAIL.n437 VTAIL.n413 1.93989
R2057 VTAIL.n372 VTAIL.n328 1.93989
R2058 VTAIL.n359 VTAIL.n335 1.93989
R2059 VTAIL.n292 VTAIL.n248 1.93989
R2060 VTAIL.n279 VTAIL.n255 1.93989
R2061 VTAIL.n0 VTAIL.t13 1.39095
R2062 VTAIL.n0 VTAIL.t7 1.39095
R2063 VTAIL.n158 VTAIL.t0 1.39095
R2064 VTAIL.n158 VTAIL.t3 1.39095
R2065 VTAIL.n474 VTAIL.t4 1.39095
R2066 VTAIL.n474 VTAIL.t1 1.39095
R2067 VTAIL.n316 VTAIL.t11 1.39095
R2068 VTAIL.n316 VTAIL.t8 1.39095
R2069 VTAIL.n599 VTAIL.n597 1.16414
R2070 VTAIL.n607 VTAIL.n566 1.16414
R2071 VTAIL.n47 VTAIL.n45 1.16414
R2072 VTAIL.n55 VTAIL.n14 1.16414
R2073 VTAIL.n125 VTAIL.n123 1.16414
R2074 VTAIL.n133 VTAIL.n92 1.16414
R2075 VTAIL.n205 VTAIL.n203 1.16414
R2076 VTAIL.n213 VTAIL.n172 1.16414
R2077 VTAIL.n529 VTAIL.n488 1.16414
R2078 VTAIL.n521 VTAIL.n520 1.16414
R2079 VTAIL.n449 VTAIL.n408 1.16414
R2080 VTAIL.n441 VTAIL.n440 1.16414
R2081 VTAIL.n371 VTAIL.n330 1.16414
R2082 VTAIL.n363 VTAIL.n362 1.16414
R2083 VTAIL.n291 VTAIL.n250 1.16414
R2084 VTAIL.n283 VTAIL.n282 1.16414
R2085 VTAIL.n317 VTAIL.n315 0.681535
R2086 VTAIL.n395 VTAIL.n317 0.681535
R2087 VTAIL.n475 VTAIL.n473 0.681535
R2088 VTAIL.n553 VTAIL.n475 0.681535
R2089 VTAIL.n237 VTAIL.n159 0.681535
R2090 VTAIL.n159 VTAIL.n157 0.681535
R2091 VTAIL.n79 VTAIL.n1 0.681535
R2092 VTAIL VTAIL.n631 0.623345
R2093 VTAIL.n473 VTAIL.n395 0.470328
R2094 VTAIL.n157 VTAIL.n79 0.470328
R2095 VTAIL.n598 VTAIL.n568 0.388379
R2096 VTAIL.n604 VTAIL.n603 0.388379
R2097 VTAIL.n46 VTAIL.n16 0.388379
R2098 VTAIL.n52 VTAIL.n51 0.388379
R2099 VTAIL.n124 VTAIL.n94 0.388379
R2100 VTAIL.n130 VTAIL.n129 0.388379
R2101 VTAIL.n204 VTAIL.n174 0.388379
R2102 VTAIL.n210 VTAIL.n209 0.388379
R2103 VTAIL.n526 VTAIL.n525 0.388379
R2104 VTAIL.n492 VTAIL.n490 0.388379
R2105 VTAIL.n446 VTAIL.n445 0.388379
R2106 VTAIL.n412 VTAIL.n410 0.388379
R2107 VTAIL.n368 VTAIL.n367 0.388379
R2108 VTAIL.n334 VTAIL.n332 0.388379
R2109 VTAIL.n288 VTAIL.n287 0.388379
R2110 VTAIL.n254 VTAIL.n252 0.388379
R2111 VTAIL.n580 VTAIL.n575 0.155672
R2112 VTAIL.n587 VTAIL.n575 0.155672
R2113 VTAIL.n588 VTAIL.n587 0.155672
R2114 VTAIL.n588 VTAIL.n571 0.155672
R2115 VTAIL.n595 VTAIL.n571 0.155672
R2116 VTAIL.n596 VTAIL.n595 0.155672
R2117 VTAIL.n596 VTAIL.n567 0.155672
R2118 VTAIL.n605 VTAIL.n567 0.155672
R2119 VTAIL.n606 VTAIL.n605 0.155672
R2120 VTAIL.n606 VTAIL.n563 0.155672
R2121 VTAIL.n613 VTAIL.n563 0.155672
R2122 VTAIL.n614 VTAIL.n613 0.155672
R2123 VTAIL.n614 VTAIL.n559 0.155672
R2124 VTAIL.n621 VTAIL.n559 0.155672
R2125 VTAIL.n622 VTAIL.n621 0.155672
R2126 VTAIL.n622 VTAIL.n555 0.155672
R2127 VTAIL.n629 VTAIL.n555 0.155672
R2128 VTAIL.n28 VTAIL.n23 0.155672
R2129 VTAIL.n35 VTAIL.n23 0.155672
R2130 VTAIL.n36 VTAIL.n35 0.155672
R2131 VTAIL.n36 VTAIL.n19 0.155672
R2132 VTAIL.n43 VTAIL.n19 0.155672
R2133 VTAIL.n44 VTAIL.n43 0.155672
R2134 VTAIL.n44 VTAIL.n15 0.155672
R2135 VTAIL.n53 VTAIL.n15 0.155672
R2136 VTAIL.n54 VTAIL.n53 0.155672
R2137 VTAIL.n54 VTAIL.n11 0.155672
R2138 VTAIL.n61 VTAIL.n11 0.155672
R2139 VTAIL.n62 VTAIL.n61 0.155672
R2140 VTAIL.n62 VTAIL.n7 0.155672
R2141 VTAIL.n69 VTAIL.n7 0.155672
R2142 VTAIL.n70 VTAIL.n69 0.155672
R2143 VTAIL.n70 VTAIL.n3 0.155672
R2144 VTAIL.n77 VTAIL.n3 0.155672
R2145 VTAIL.n106 VTAIL.n101 0.155672
R2146 VTAIL.n113 VTAIL.n101 0.155672
R2147 VTAIL.n114 VTAIL.n113 0.155672
R2148 VTAIL.n114 VTAIL.n97 0.155672
R2149 VTAIL.n121 VTAIL.n97 0.155672
R2150 VTAIL.n122 VTAIL.n121 0.155672
R2151 VTAIL.n122 VTAIL.n93 0.155672
R2152 VTAIL.n131 VTAIL.n93 0.155672
R2153 VTAIL.n132 VTAIL.n131 0.155672
R2154 VTAIL.n132 VTAIL.n89 0.155672
R2155 VTAIL.n139 VTAIL.n89 0.155672
R2156 VTAIL.n140 VTAIL.n139 0.155672
R2157 VTAIL.n140 VTAIL.n85 0.155672
R2158 VTAIL.n147 VTAIL.n85 0.155672
R2159 VTAIL.n148 VTAIL.n147 0.155672
R2160 VTAIL.n148 VTAIL.n81 0.155672
R2161 VTAIL.n155 VTAIL.n81 0.155672
R2162 VTAIL.n186 VTAIL.n181 0.155672
R2163 VTAIL.n193 VTAIL.n181 0.155672
R2164 VTAIL.n194 VTAIL.n193 0.155672
R2165 VTAIL.n194 VTAIL.n177 0.155672
R2166 VTAIL.n201 VTAIL.n177 0.155672
R2167 VTAIL.n202 VTAIL.n201 0.155672
R2168 VTAIL.n202 VTAIL.n173 0.155672
R2169 VTAIL.n211 VTAIL.n173 0.155672
R2170 VTAIL.n212 VTAIL.n211 0.155672
R2171 VTAIL.n212 VTAIL.n169 0.155672
R2172 VTAIL.n219 VTAIL.n169 0.155672
R2173 VTAIL.n220 VTAIL.n219 0.155672
R2174 VTAIL.n220 VTAIL.n165 0.155672
R2175 VTAIL.n227 VTAIL.n165 0.155672
R2176 VTAIL.n228 VTAIL.n227 0.155672
R2177 VTAIL.n228 VTAIL.n161 0.155672
R2178 VTAIL.n235 VTAIL.n161 0.155672
R2179 VTAIL.n551 VTAIL.n477 0.155672
R2180 VTAIL.n544 VTAIL.n477 0.155672
R2181 VTAIL.n544 VTAIL.n543 0.155672
R2182 VTAIL.n543 VTAIL.n481 0.155672
R2183 VTAIL.n536 VTAIL.n481 0.155672
R2184 VTAIL.n536 VTAIL.n535 0.155672
R2185 VTAIL.n535 VTAIL.n485 0.155672
R2186 VTAIL.n528 VTAIL.n485 0.155672
R2187 VTAIL.n528 VTAIL.n527 0.155672
R2188 VTAIL.n527 VTAIL.n489 0.155672
R2189 VTAIL.n519 VTAIL.n489 0.155672
R2190 VTAIL.n519 VTAIL.n518 0.155672
R2191 VTAIL.n518 VTAIL.n494 0.155672
R2192 VTAIL.n511 VTAIL.n494 0.155672
R2193 VTAIL.n511 VTAIL.n510 0.155672
R2194 VTAIL.n510 VTAIL.n498 0.155672
R2195 VTAIL.n503 VTAIL.n498 0.155672
R2196 VTAIL.n471 VTAIL.n397 0.155672
R2197 VTAIL.n464 VTAIL.n397 0.155672
R2198 VTAIL.n464 VTAIL.n463 0.155672
R2199 VTAIL.n463 VTAIL.n401 0.155672
R2200 VTAIL.n456 VTAIL.n401 0.155672
R2201 VTAIL.n456 VTAIL.n455 0.155672
R2202 VTAIL.n455 VTAIL.n405 0.155672
R2203 VTAIL.n448 VTAIL.n405 0.155672
R2204 VTAIL.n448 VTAIL.n447 0.155672
R2205 VTAIL.n447 VTAIL.n409 0.155672
R2206 VTAIL.n439 VTAIL.n409 0.155672
R2207 VTAIL.n439 VTAIL.n438 0.155672
R2208 VTAIL.n438 VTAIL.n414 0.155672
R2209 VTAIL.n431 VTAIL.n414 0.155672
R2210 VTAIL.n431 VTAIL.n430 0.155672
R2211 VTAIL.n430 VTAIL.n418 0.155672
R2212 VTAIL.n423 VTAIL.n418 0.155672
R2213 VTAIL.n393 VTAIL.n319 0.155672
R2214 VTAIL.n386 VTAIL.n319 0.155672
R2215 VTAIL.n386 VTAIL.n385 0.155672
R2216 VTAIL.n385 VTAIL.n323 0.155672
R2217 VTAIL.n378 VTAIL.n323 0.155672
R2218 VTAIL.n378 VTAIL.n377 0.155672
R2219 VTAIL.n377 VTAIL.n327 0.155672
R2220 VTAIL.n370 VTAIL.n327 0.155672
R2221 VTAIL.n370 VTAIL.n369 0.155672
R2222 VTAIL.n369 VTAIL.n331 0.155672
R2223 VTAIL.n361 VTAIL.n331 0.155672
R2224 VTAIL.n361 VTAIL.n360 0.155672
R2225 VTAIL.n360 VTAIL.n336 0.155672
R2226 VTAIL.n353 VTAIL.n336 0.155672
R2227 VTAIL.n353 VTAIL.n352 0.155672
R2228 VTAIL.n352 VTAIL.n340 0.155672
R2229 VTAIL.n345 VTAIL.n340 0.155672
R2230 VTAIL.n313 VTAIL.n239 0.155672
R2231 VTAIL.n306 VTAIL.n239 0.155672
R2232 VTAIL.n306 VTAIL.n305 0.155672
R2233 VTAIL.n305 VTAIL.n243 0.155672
R2234 VTAIL.n298 VTAIL.n243 0.155672
R2235 VTAIL.n298 VTAIL.n297 0.155672
R2236 VTAIL.n297 VTAIL.n247 0.155672
R2237 VTAIL.n290 VTAIL.n247 0.155672
R2238 VTAIL.n290 VTAIL.n289 0.155672
R2239 VTAIL.n289 VTAIL.n251 0.155672
R2240 VTAIL.n281 VTAIL.n251 0.155672
R2241 VTAIL.n281 VTAIL.n280 0.155672
R2242 VTAIL.n280 VTAIL.n256 0.155672
R2243 VTAIL.n273 VTAIL.n256 0.155672
R2244 VTAIL.n273 VTAIL.n272 0.155672
R2245 VTAIL.n272 VTAIL.n260 0.155672
R2246 VTAIL.n265 VTAIL.n260 0.155672
R2247 VTAIL VTAIL.n1 0.0586897
R2248 VP.n4 VP.t6 853.48
R2249 VP.n10 VP.t1 832.499
R2250 VP.n1 VP.t7 832.499
R2251 VP.n15 VP.t2 832.499
R2252 VP.n16 VP.t0 832.499
R2253 VP.n8 VP.t5 832.499
R2254 VP.n7 VP.t4 832.499
R2255 VP.n3 VP.t3 832.499
R2256 VP.n17 VP.n16 161.3
R2257 VP.n6 VP.n5 161.3
R2258 VP.n7 VP.n2 161.3
R2259 VP.n9 VP.n8 161.3
R2260 VP.n15 VP.n0 161.3
R2261 VP.n14 VP.n13 161.3
R2262 VP.n12 VP.n1 161.3
R2263 VP.n11 VP.n10 161.3
R2264 VP.n5 VP.n4 70.4033
R2265 VP.n10 VP.n1 48.2005
R2266 VP.n16 VP.n15 48.2005
R2267 VP.n8 VP.n7 48.2005
R2268 VP.n11 VP.n9 42.6141
R2269 VP.n14 VP.n1 24.1005
R2270 VP.n15 VP.n14 24.1005
R2271 VP.n6 VP.n3 24.1005
R2272 VP.n7 VP.n6 24.1005
R2273 VP.n4 VP.n3 20.9576
R2274 VP.n5 VP.n2 0.189894
R2275 VP.n9 VP.n2 0.189894
R2276 VP.n12 VP.n11 0.189894
R2277 VP.n13 VP.n12 0.189894
R2278 VP.n13 VP.n0 0.189894
R2279 VP.n17 VP.n0 0.189894
R2280 VP VP.n17 0.0516364
R2281 VDD1 VDD1.n0 61.0511
R2282 VDD1.n3 VDD1.n2 60.9376
R2283 VDD1.n3 VDD1.n1 60.9376
R2284 VDD1.n5 VDD1.n4 60.6524
R2285 VDD1.n5 VDD1.n3 39.6388
R2286 VDD1.n4 VDD1.t3 1.39095
R2287 VDD1.n4 VDD1.t2 1.39095
R2288 VDD1.n0 VDD1.t1 1.39095
R2289 VDD1.n0 VDD1.t4 1.39095
R2290 VDD1.n2 VDD1.t5 1.39095
R2291 VDD1.n2 VDD1.t7 1.39095
R2292 VDD1.n1 VDD1.t6 1.39095
R2293 VDD1.n1 VDD1.t0 1.39095
R2294 VDD1 VDD1.n5 0.282828
C0 VDD2 VP 0.291656f
C1 VDD1 VP 5.23952f
C2 VP VN 5.46331f
C3 VDD1 VDD2 0.709053f
C4 VP VTAIL 4.68494f
C5 VDD2 VN 5.09574f
C6 VDD2 VTAIL 15.6547f
C7 VDD1 VN 0.147563f
C8 VDD1 VTAIL 15.6146f
C9 VN VTAIL 4.67083f
C10 VDD2 B 3.458879f
C11 VDD1 B 3.666906f
C12 VTAIL B 9.913359f
C13 VN B 8.101939f
C14 VP B 5.844716f
C15 VDD1.t1 B 0.336637f
C16 VDD1.t4 B 0.336637f
C17 VDD1.n0 B 3.02932f
C18 VDD1.t6 B 0.336637f
C19 VDD1.t0 B 0.336637f
C20 VDD1.n1 B 3.0286f
C21 VDD1.t5 B 0.336637f
C22 VDD1.t7 B 0.336637f
C23 VDD1.n2 B 3.0286f
C24 VDD1.n3 B 2.67164f
C25 VDD1.t3 B 0.336637f
C26 VDD1.t2 B 0.336637f
C27 VDD1.n4 B 3.02691f
C28 VDD1.n5 B 2.8901f
C29 VP.n0 B 0.050913f
C30 VP.t7 B 0.948839f
C31 VP.n1 B 0.37881f
C32 VP.n2 B 0.050913f
C33 VP.t5 B 0.948839f
C34 VP.t4 B 0.948839f
C35 VP.t3 B 0.948839f
C36 VP.n3 B 0.37881f
C37 VP.t6 B 0.958026f
C38 VP.n4 B 0.364817f
C39 VP.n5 B 0.162723f
C40 VP.n6 B 0.011553f
C41 VP.n7 B 0.37881f
C42 VP.n8 B 0.37363f
C43 VP.n9 B 2.15279f
C44 VP.t1 B 0.948839f
C45 VP.n10 B 0.37363f
C46 VP.n11 B 2.19561f
C47 VP.n12 B 0.050913f
C48 VP.n13 B 0.050913f
C49 VP.n14 B 0.011553f
C50 VP.t2 B 0.948839f
C51 VP.n15 B 0.37881f
C52 VP.t0 B 0.948839f
C53 VP.n16 B 0.37363f
C54 VP.n17 B 0.039455f
C55 VTAIL.t13 B 0.241412f
C56 VTAIL.t7 B 0.241412f
C57 VTAIL.n0 B 2.10358f
C58 VTAIL.n1 B 0.270016f
C59 VTAIL.n2 B 0.031312f
C60 VTAIL.n3 B 0.021453f
C61 VTAIL.n4 B 0.011528f
C62 VTAIL.n5 B 0.027248f
C63 VTAIL.n6 B 0.012206f
C64 VTAIL.n7 B 0.021453f
C65 VTAIL.n8 B 0.011528f
C66 VTAIL.n9 B 0.027248f
C67 VTAIL.n10 B 0.012206f
C68 VTAIL.n11 B 0.021453f
C69 VTAIL.n12 B 0.011528f
C70 VTAIL.n13 B 0.027248f
C71 VTAIL.n14 B 0.012206f
C72 VTAIL.n15 B 0.021453f
C73 VTAIL.n16 B 0.011867f
C74 VTAIL.n17 B 0.027248f
C75 VTAIL.n18 B 0.012206f
C76 VTAIL.n19 B 0.021453f
C77 VTAIL.n20 B 0.011528f
C78 VTAIL.n21 B 0.027248f
C79 VTAIL.n22 B 0.012206f
C80 VTAIL.n23 B 0.021453f
C81 VTAIL.n24 B 0.011528f
C82 VTAIL.n25 B 0.020436f
C83 VTAIL.n26 B 0.019262f
C84 VTAIL.t14 B 0.046279f
C85 VTAIL.n27 B 0.173125f
C86 VTAIL.n28 B 1.29603f
C87 VTAIL.n29 B 0.011528f
C88 VTAIL.n30 B 0.012206f
C89 VTAIL.n31 B 0.027248f
C90 VTAIL.n32 B 0.027248f
C91 VTAIL.n33 B 0.012206f
C92 VTAIL.n34 B 0.011528f
C93 VTAIL.n35 B 0.021453f
C94 VTAIL.n36 B 0.021453f
C95 VTAIL.n37 B 0.011528f
C96 VTAIL.n38 B 0.012206f
C97 VTAIL.n39 B 0.027248f
C98 VTAIL.n40 B 0.027248f
C99 VTAIL.n41 B 0.012206f
C100 VTAIL.n42 B 0.011528f
C101 VTAIL.n43 B 0.021453f
C102 VTAIL.n44 B 0.021453f
C103 VTAIL.n45 B 0.011528f
C104 VTAIL.n46 B 0.011528f
C105 VTAIL.n47 B 0.012206f
C106 VTAIL.n48 B 0.027248f
C107 VTAIL.n49 B 0.027248f
C108 VTAIL.n50 B 0.027248f
C109 VTAIL.n51 B 0.011867f
C110 VTAIL.n52 B 0.011528f
C111 VTAIL.n53 B 0.021453f
C112 VTAIL.n54 B 0.021453f
C113 VTAIL.n55 B 0.011528f
C114 VTAIL.n56 B 0.012206f
C115 VTAIL.n57 B 0.027248f
C116 VTAIL.n58 B 0.027248f
C117 VTAIL.n59 B 0.012206f
C118 VTAIL.n60 B 0.011528f
C119 VTAIL.n61 B 0.021453f
C120 VTAIL.n62 B 0.021453f
C121 VTAIL.n63 B 0.011528f
C122 VTAIL.n64 B 0.012206f
C123 VTAIL.n65 B 0.027248f
C124 VTAIL.n66 B 0.027248f
C125 VTAIL.n67 B 0.012206f
C126 VTAIL.n68 B 0.011528f
C127 VTAIL.n69 B 0.021453f
C128 VTAIL.n70 B 0.021453f
C129 VTAIL.n71 B 0.011528f
C130 VTAIL.n72 B 0.012206f
C131 VTAIL.n73 B 0.027248f
C132 VTAIL.n74 B 0.061035f
C133 VTAIL.n75 B 0.012206f
C134 VTAIL.n76 B 0.011528f
C135 VTAIL.n77 B 0.048416f
C136 VTAIL.n78 B 0.034326f
C137 VTAIL.n79 B 0.097218f
C138 VTAIL.n80 B 0.031312f
C139 VTAIL.n81 B 0.021453f
C140 VTAIL.n82 B 0.011528f
C141 VTAIL.n83 B 0.027248f
C142 VTAIL.n84 B 0.012206f
C143 VTAIL.n85 B 0.021453f
C144 VTAIL.n86 B 0.011528f
C145 VTAIL.n87 B 0.027248f
C146 VTAIL.n88 B 0.012206f
C147 VTAIL.n89 B 0.021453f
C148 VTAIL.n90 B 0.011528f
C149 VTAIL.n91 B 0.027248f
C150 VTAIL.n92 B 0.012206f
C151 VTAIL.n93 B 0.021453f
C152 VTAIL.n94 B 0.011867f
C153 VTAIL.n95 B 0.027248f
C154 VTAIL.n96 B 0.012206f
C155 VTAIL.n97 B 0.021453f
C156 VTAIL.n98 B 0.011528f
C157 VTAIL.n99 B 0.027248f
C158 VTAIL.n100 B 0.012206f
C159 VTAIL.n101 B 0.021453f
C160 VTAIL.n102 B 0.011528f
C161 VTAIL.n103 B 0.020436f
C162 VTAIL.n104 B 0.019262f
C163 VTAIL.t5 B 0.046279f
C164 VTAIL.n105 B 0.173125f
C165 VTAIL.n106 B 1.29603f
C166 VTAIL.n107 B 0.011528f
C167 VTAIL.n108 B 0.012206f
C168 VTAIL.n109 B 0.027248f
C169 VTAIL.n110 B 0.027248f
C170 VTAIL.n111 B 0.012206f
C171 VTAIL.n112 B 0.011528f
C172 VTAIL.n113 B 0.021453f
C173 VTAIL.n114 B 0.021453f
C174 VTAIL.n115 B 0.011528f
C175 VTAIL.n116 B 0.012206f
C176 VTAIL.n117 B 0.027248f
C177 VTAIL.n118 B 0.027248f
C178 VTAIL.n119 B 0.012206f
C179 VTAIL.n120 B 0.011528f
C180 VTAIL.n121 B 0.021453f
C181 VTAIL.n122 B 0.021453f
C182 VTAIL.n123 B 0.011528f
C183 VTAIL.n124 B 0.011528f
C184 VTAIL.n125 B 0.012206f
C185 VTAIL.n126 B 0.027248f
C186 VTAIL.n127 B 0.027248f
C187 VTAIL.n128 B 0.027248f
C188 VTAIL.n129 B 0.011867f
C189 VTAIL.n130 B 0.011528f
C190 VTAIL.n131 B 0.021453f
C191 VTAIL.n132 B 0.021453f
C192 VTAIL.n133 B 0.011528f
C193 VTAIL.n134 B 0.012206f
C194 VTAIL.n135 B 0.027248f
C195 VTAIL.n136 B 0.027248f
C196 VTAIL.n137 B 0.012206f
C197 VTAIL.n138 B 0.011528f
C198 VTAIL.n139 B 0.021453f
C199 VTAIL.n140 B 0.021453f
C200 VTAIL.n141 B 0.011528f
C201 VTAIL.n142 B 0.012206f
C202 VTAIL.n143 B 0.027248f
C203 VTAIL.n144 B 0.027248f
C204 VTAIL.n145 B 0.012206f
C205 VTAIL.n146 B 0.011528f
C206 VTAIL.n147 B 0.021453f
C207 VTAIL.n148 B 0.021453f
C208 VTAIL.n149 B 0.011528f
C209 VTAIL.n150 B 0.012206f
C210 VTAIL.n151 B 0.027248f
C211 VTAIL.n152 B 0.061035f
C212 VTAIL.n153 B 0.012206f
C213 VTAIL.n154 B 0.011528f
C214 VTAIL.n155 B 0.048416f
C215 VTAIL.n156 B 0.034326f
C216 VTAIL.n157 B 0.097218f
C217 VTAIL.t0 B 0.241412f
C218 VTAIL.t3 B 0.241412f
C219 VTAIL.n158 B 2.10358f
C220 VTAIL.n159 B 0.313071f
C221 VTAIL.n160 B 0.031312f
C222 VTAIL.n161 B 0.021453f
C223 VTAIL.n162 B 0.011528f
C224 VTAIL.n163 B 0.027248f
C225 VTAIL.n164 B 0.012206f
C226 VTAIL.n165 B 0.021453f
C227 VTAIL.n166 B 0.011528f
C228 VTAIL.n167 B 0.027248f
C229 VTAIL.n168 B 0.012206f
C230 VTAIL.n169 B 0.021453f
C231 VTAIL.n170 B 0.011528f
C232 VTAIL.n171 B 0.027248f
C233 VTAIL.n172 B 0.012206f
C234 VTAIL.n173 B 0.021453f
C235 VTAIL.n174 B 0.011867f
C236 VTAIL.n175 B 0.027248f
C237 VTAIL.n176 B 0.012206f
C238 VTAIL.n177 B 0.021453f
C239 VTAIL.n178 B 0.011528f
C240 VTAIL.n179 B 0.027248f
C241 VTAIL.n180 B 0.012206f
C242 VTAIL.n181 B 0.021453f
C243 VTAIL.n182 B 0.011528f
C244 VTAIL.n183 B 0.020436f
C245 VTAIL.n184 B 0.019262f
C246 VTAIL.t2 B 0.046279f
C247 VTAIL.n185 B 0.173125f
C248 VTAIL.n186 B 1.29603f
C249 VTAIL.n187 B 0.011528f
C250 VTAIL.n188 B 0.012206f
C251 VTAIL.n189 B 0.027248f
C252 VTAIL.n190 B 0.027248f
C253 VTAIL.n191 B 0.012206f
C254 VTAIL.n192 B 0.011528f
C255 VTAIL.n193 B 0.021453f
C256 VTAIL.n194 B 0.021453f
C257 VTAIL.n195 B 0.011528f
C258 VTAIL.n196 B 0.012206f
C259 VTAIL.n197 B 0.027248f
C260 VTAIL.n198 B 0.027248f
C261 VTAIL.n199 B 0.012206f
C262 VTAIL.n200 B 0.011528f
C263 VTAIL.n201 B 0.021453f
C264 VTAIL.n202 B 0.021453f
C265 VTAIL.n203 B 0.011528f
C266 VTAIL.n204 B 0.011528f
C267 VTAIL.n205 B 0.012206f
C268 VTAIL.n206 B 0.027248f
C269 VTAIL.n207 B 0.027248f
C270 VTAIL.n208 B 0.027248f
C271 VTAIL.n209 B 0.011867f
C272 VTAIL.n210 B 0.011528f
C273 VTAIL.n211 B 0.021453f
C274 VTAIL.n212 B 0.021453f
C275 VTAIL.n213 B 0.011528f
C276 VTAIL.n214 B 0.012206f
C277 VTAIL.n215 B 0.027248f
C278 VTAIL.n216 B 0.027248f
C279 VTAIL.n217 B 0.012206f
C280 VTAIL.n218 B 0.011528f
C281 VTAIL.n219 B 0.021453f
C282 VTAIL.n220 B 0.021453f
C283 VTAIL.n221 B 0.011528f
C284 VTAIL.n222 B 0.012206f
C285 VTAIL.n223 B 0.027248f
C286 VTAIL.n224 B 0.027248f
C287 VTAIL.n225 B 0.012206f
C288 VTAIL.n226 B 0.011528f
C289 VTAIL.n227 B 0.021453f
C290 VTAIL.n228 B 0.021453f
C291 VTAIL.n229 B 0.011528f
C292 VTAIL.n230 B 0.012206f
C293 VTAIL.n231 B 0.027248f
C294 VTAIL.n232 B 0.061035f
C295 VTAIL.n233 B 0.012206f
C296 VTAIL.n234 B 0.011528f
C297 VTAIL.n235 B 0.048416f
C298 VTAIL.n236 B 0.034326f
C299 VTAIL.n237 B 1.25183f
C300 VTAIL.n238 B 0.031312f
C301 VTAIL.n239 B 0.021453f
C302 VTAIL.n240 B 0.011528f
C303 VTAIL.n241 B 0.027248f
C304 VTAIL.n242 B 0.012206f
C305 VTAIL.n243 B 0.021453f
C306 VTAIL.n244 B 0.011528f
C307 VTAIL.n245 B 0.027248f
C308 VTAIL.n246 B 0.012206f
C309 VTAIL.n247 B 0.021453f
C310 VTAIL.n248 B 0.011528f
C311 VTAIL.n249 B 0.027248f
C312 VTAIL.n250 B 0.012206f
C313 VTAIL.n251 B 0.021453f
C314 VTAIL.n252 B 0.011867f
C315 VTAIL.n253 B 0.027248f
C316 VTAIL.n254 B 0.011528f
C317 VTAIL.n255 B 0.012206f
C318 VTAIL.n256 B 0.021453f
C319 VTAIL.n257 B 0.011528f
C320 VTAIL.n258 B 0.027248f
C321 VTAIL.n259 B 0.012206f
C322 VTAIL.n260 B 0.021453f
C323 VTAIL.n261 B 0.011528f
C324 VTAIL.n262 B 0.020436f
C325 VTAIL.n263 B 0.019262f
C326 VTAIL.t10 B 0.046279f
C327 VTAIL.n264 B 0.173125f
C328 VTAIL.n265 B 1.29603f
C329 VTAIL.n266 B 0.011528f
C330 VTAIL.n267 B 0.012206f
C331 VTAIL.n268 B 0.027248f
C332 VTAIL.n269 B 0.027248f
C333 VTAIL.n270 B 0.012206f
C334 VTAIL.n271 B 0.011528f
C335 VTAIL.n272 B 0.021453f
C336 VTAIL.n273 B 0.021453f
C337 VTAIL.n274 B 0.011528f
C338 VTAIL.n275 B 0.012206f
C339 VTAIL.n276 B 0.027248f
C340 VTAIL.n277 B 0.027248f
C341 VTAIL.n278 B 0.012206f
C342 VTAIL.n279 B 0.011528f
C343 VTAIL.n280 B 0.021453f
C344 VTAIL.n281 B 0.021453f
C345 VTAIL.n282 B 0.011528f
C346 VTAIL.n283 B 0.012206f
C347 VTAIL.n284 B 0.027248f
C348 VTAIL.n285 B 0.027248f
C349 VTAIL.n286 B 0.027248f
C350 VTAIL.n287 B 0.011867f
C351 VTAIL.n288 B 0.011528f
C352 VTAIL.n289 B 0.021453f
C353 VTAIL.n290 B 0.021453f
C354 VTAIL.n291 B 0.011528f
C355 VTAIL.n292 B 0.012206f
C356 VTAIL.n293 B 0.027248f
C357 VTAIL.n294 B 0.027248f
C358 VTAIL.n295 B 0.012206f
C359 VTAIL.n296 B 0.011528f
C360 VTAIL.n297 B 0.021453f
C361 VTAIL.n298 B 0.021453f
C362 VTAIL.n299 B 0.011528f
C363 VTAIL.n300 B 0.012206f
C364 VTAIL.n301 B 0.027248f
C365 VTAIL.n302 B 0.027248f
C366 VTAIL.n303 B 0.012206f
C367 VTAIL.n304 B 0.011528f
C368 VTAIL.n305 B 0.021453f
C369 VTAIL.n306 B 0.021453f
C370 VTAIL.n307 B 0.011528f
C371 VTAIL.n308 B 0.012206f
C372 VTAIL.n309 B 0.027248f
C373 VTAIL.n310 B 0.061035f
C374 VTAIL.n311 B 0.012206f
C375 VTAIL.n312 B 0.011528f
C376 VTAIL.n313 B 0.048416f
C377 VTAIL.n314 B 0.034326f
C378 VTAIL.n315 B 1.25183f
C379 VTAIL.t11 B 0.241412f
C380 VTAIL.t8 B 0.241412f
C381 VTAIL.n316 B 2.10359f
C382 VTAIL.n317 B 0.313068f
C383 VTAIL.n318 B 0.031312f
C384 VTAIL.n319 B 0.021453f
C385 VTAIL.n320 B 0.011528f
C386 VTAIL.n321 B 0.027248f
C387 VTAIL.n322 B 0.012206f
C388 VTAIL.n323 B 0.021453f
C389 VTAIL.n324 B 0.011528f
C390 VTAIL.n325 B 0.027248f
C391 VTAIL.n326 B 0.012206f
C392 VTAIL.n327 B 0.021453f
C393 VTAIL.n328 B 0.011528f
C394 VTAIL.n329 B 0.027248f
C395 VTAIL.n330 B 0.012206f
C396 VTAIL.n331 B 0.021453f
C397 VTAIL.n332 B 0.011867f
C398 VTAIL.n333 B 0.027248f
C399 VTAIL.n334 B 0.011528f
C400 VTAIL.n335 B 0.012206f
C401 VTAIL.n336 B 0.021453f
C402 VTAIL.n337 B 0.011528f
C403 VTAIL.n338 B 0.027248f
C404 VTAIL.n339 B 0.012206f
C405 VTAIL.n340 B 0.021453f
C406 VTAIL.n341 B 0.011528f
C407 VTAIL.n342 B 0.020436f
C408 VTAIL.n343 B 0.019262f
C409 VTAIL.t9 B 0.046279f
C410 VTAIL.n344 B 0.173125f
C411 VTAIL.n345 B 1.29603f
C412 VTAIL.n346 B 0.011528f
C413 VTAIL.n347 B 0.012206f
C414 VTAIL.n348 B 0.027248f
C415 VTAIL.n349 B 0.027248f
C416 VTAIL.n350 B 0.012206f
C417 VTAIL.n351 B 0.011528f
C418 VTAIL.n352 B 0.021453f
C419 VTAIL.n353 B 0.021453f
C420 VTAIL.n354 B 0.011528f
C421 VTAIL.n355 B 0.012206f
C422 VTAIL.n356 B 0.027248f
C423 VTAIL.n357 B 0.027248f
C424 VTAIL.n358 B 0.012206f
C425 VTAIL.n359 B 0.011528f
C426 VTAIL.n360 B 0.021453f
C427 VTAIL.n361 B 0.021453f
C428 VTAIL.n362 B 0.011528f
C429 VTAIL.n363 B 0.012206f
C430 VTAIL.n364 B 0.027248f
C431 VTAIL.n365 B 0.027248f
C432 VTAIL.n366 B 0.027248f
C433 VTAIL.n367 B 0.011867f
C434 VTAIL.n368 B 0.011528f
C435 VTAIL.n369 B 0.021453f
C436 VTAIL.n370 B 0.021453f
C437 VTAIL.n371 B 0.011528f
C438 VTAIL.n372 B 0.012206f
C439 VTAIL.n373 B 0.027248f
C440 VTAIL.n374 B 0.027248f
C441 VTAIL.n375 B 0.012206f
C442 VTAIL.n376 B 0.011528f
C443 VTAIL.n377 B 0.021453f
C444 VTAIL.n378 B 0.021453f
C445 VTAIL.n379 B 0.011528f
C446 VTAIL.n380 B 0.012206f
C447 VTAIL.n381 B 0.027248f
C448 VTAIL.n382 B 0.027248f
C449 VTAIL.n383 B 0.012206f
C450 VTAIL.n384 B 0.011528f
C451 VTAIL.n385 B 0.021453f
C452 VTAIL.n386 B 0.021453f
C453 VTAIL.n387 B 0.011528f
C454 VTAIL.n388 B 0.012206f
C455 VTAIL.n389 B 0.027248f
C456 VTAIL.n390 B 0.061035f
C457 VTAIL.n391 B 0.012206f
C458 VTAIL.n392 B 0.011528f
C459 VTAIL.n393 B 0.048416f
C460 VTAIL.n394 B 0.034326f
C461 VTAIL.n395 B 0.097218f
C462 VTAIL.n396 B 0.031312f
C463 VTAIL.n397 B 0.021453f
C464 VTAIL.n398 B 0.011528f
C465 VTAIL.n399 B 0.027248f
C466 VTAIL.n400 B 0.012206f
C467 VTAIL.n401 B 0.021453f
C468 VTAIL.n402 B 0.011528f
C469 VTAIL.n403 B 0.027248f
C470 VTAIL.n404 B 0.012206f
C471 VTAIL.n405 B 0.021453f
C472 VTAIL.n406 B 0.011528f
C473 VTAIL.n407 B 0.027248f
C474 VTAIL.n408 B 0.012206f
C475 VTAIL.n409 B 0.021453f
C476 VTAIL.n410 B 0.011867f
C477 VTAIL.n411 B 0.027248f
C478 VTAIL.n412 B 0.011528f
C479 VTAIL.n413 B 0.012206f
C480 VTAIL.n414 B 0.021453f
C481 VTAIL.n415 B 0.011528f
C482 VTAIL.n416 B 0.027248f
C483 VTAIL.n417 B 0.012206f
C484 VTAIL.n418 B 0.021453f
C485 VTAIL.n419 B 0.011528f
C486 VTAIL.n420 B 0.020436f
C487 VTAIL.n421 B 0.019262f
C488 VTAIL.t6 B 0.046279f
C489 VTAIL.n422 B 0.173125f
C490 VTAIL.n423 B 1.29603f
C491 VTAIL.n424 B 0.011528f
C492 VTAIL.n425 B 0.012206f
C493 VTAIL.n426 B 0.027248f
C494 VTAIL.n427 B 0.027248f
C495 VTAIL.n428 B 0.012206f
C496 VTAIL.n429 B 0.011528f
C497 VTAIL.n430 B 0.021453f
C498 VTAIL.n431 B 0.021453f
C499 VTAIL.n432 B 0.011528f
C500 VTAIL.n433 B 0.012206f
C501 VTAIL.n434 B 0.027248f
C502 VTAIL.n435 B 0.027248f
C503 VTAIL.n436 B 0.012206f
C504 VTAIL.n437 B 0.011528f
C505 VTAIL.n438 B 0.021453f
C506 VTAIL.n439 B 0.021453f
C507 VTAIL.n440 B 0.011528f
C508 VTAIL.n441 B 0.012206f
C509 VTAIL.n442 B 0.027248f
C510 VTAIL.n443 B 0.027248f
C511 VTAIL.n444 B 0.027248f
C512 VTAIL.n445 B 0.011867f
C513 VTAIL.n446 B 0.011528f
C514 VTAIL.n447 B 0.021453f
C515 VTAIL.n448 B 0.021453f
C516 VTAIL.n449 B 0.011528f
C517 VTAIL.n450 B 0.012206f
C518 VTAIL.n451 B 0.027248f
C519 VTAIL.n452 B 0.027248f
C520 VTAIL.n453 B 0.012206f
C521 VTAIL.n454 B 0.011528f
C522 VTAIL.n455 B 0.021453f
C523 VTAIL.n456 B 0.021453f
C524 VTAIL.n457 B 0.011528f
C525 VTAIL.n458 B 0.012206f
C526 VTAIL.n459 B 0.027248f
C527 VTAIL.n460 B 0.027248f
C528 VTAIL.n461 B 0.012206f
C529 VTAIL.n462 B 0.011528f
C530 VTAIL.n463 B 0.021453f
C531 VTAIL.n464 B 0.021453f
C532 VTAIL.n465 B 0.011528f
C533 VTAIL.n466 B 0.012206f
C534 VTAIL.n467 B 0.027248f
C535 VTAIL.n468 B 0.061035f
C536 VTAIL.n469 B 0.012206f
C537 VTAIL.n470 B 0.011528f
C538 VTAIL.n471 B 0.048416f
C539 VTAIL.n472 B 0.034326f
C540 VTAIL.n473 B 0.097218f
C541 VTAIL.t4 B 0.241412f
C542 VTAIL.t1 B 0.241412f
C543 VTAIL.n474 B 2.10359f
C544 VTAIL.n475 B 0.313068f
C545 VTAIL.n476 B 0.031312f
C546 VTAIL.n477 B 0.021453f
C547 VTAIL.n478 B 0.011528f
C548 VTAIL.n479 B 0.027248f
C549 VTAIL.n480 B 0.012206f
C550 VTAIL.n481 B 0.021453f
C551 VTAIL.n482 B 0.011528f
C552 VTAIL.n483 B 0.027248f
C553 VTAIL.n484 B 0.012206f
C554 VTAIL.n485 B 0.021453f
C555 VTAIL.n486 B 0.011528f
C556 VTAIL.n487 B 0.027248f
C557 VTAIL.n488 B 0.012206f
C558 VTAIL.n489 B 0.021453f
C559 VTAIL.n490 B 0.011867f
C560 VTAIL.n491 B 0.027248f
C561 VTAIL.n492 B 0.011528f
C562 VTAIL.n493 B 0.012206f
C563 VTAIL.n494 B 0.021453f
C564 VTAIL.n495 B 0.011528f
C565 VTAIL.n496 B 0.027248f
C566 VTAIL.n497 B 0.012206f
C567 VTAIL.n498 B 0.021453f
C568 VTAIL.n499 B 0.011528f
C569 VTAIL.n500 B 0.020436f
C570 VTAIL.n501 B 0.019262f
C571 VTAIL.t15 B 0.046279f
C572 VTAIL.n502 B 0.173125f
C573 VTAIL.n503 B 1.29603f
C574 VTAIL.n504 B 0.011528f
C575 VTAIL.n505 B 0.012206f
C576 VTAIL.n506 B 0.027248f
C577 VTAIL.n507 B 0.027248f
C578 VTAIL.n508 B 0.012206f
C579 VTAIL.n509 B 0.011528f
C580 VTAIL.n510 B 0.021453f
C581 VTAIL.n511 B 0.021453f
C582 VTAIL.n512 B 0.011528f
C583 VTAIL.n513 B 0.012206f
C584 VTAIL.n514 B 0.027248f
C585 VTAIL.n515 B 0.027248f
C586 VTAIL.n516 B 0.012206f
C587 VTAIL.n517 B 0.011528f
C588 VTAIL.n518 B 0.021453f
C589 VTAIL.n519 B 0.021453f
C590 VTAIL.n520 B 0.011528f
C591 VTAIL.n521 B 0.012206f
C592 VTAIL.n522 B 0.027248f
C593 VTAIL.n523 B 0.027248f
C594 VTAIL.n524 B 0.027248f
C595 VTAIL.n525 B 0.011867f
C596 VTAIL.n526 B 0.011528f
C597 VTAIL.n527 B 0.021453f
C598 VTAIL.n528 B 0.021453f
C599 VTAIL.n529 B 0.011528f
C600 VTAIL.n530 B 0.012206f
C601 VTAIL.n531 B 0.027248f
C602 VTAIL.n532 B 0.027248f
C603 VTAIL.n533 B 0.012206f
C604 VTAIL.n534 B 0.011528f
C605 VTAIL.n535 B 0.021453f
C606 VTAIL.n536 B 0.021453f
C607 VTAIL.n537 B 0.011528f
C608 VTAIL.n538 B 0.012206f
C609 VTAIL.n539 B 0.027248f
C610 VTAIL.n540 B 0.027248f
C611 VTAIL.n541 B 0.012206f
C612 VTAIL.n542 B 0.011528f
C613 VTAIL.n543 B 0.021453f
C614 VTAIL.n544 B 0.021453f
C615 VTAIL.n545 B 0.011528f
C616 VTAIL.n546 B 0.012206f
C617 VTAIL.n547 B 0.027248f
C618 VTAIL.n548 B 0.061035f
C619 VTAIL.n549 B 0.012206f
C620 VTAIL.n550 B 0.011528f
C621 VTAIL.n551 B 0.048416f
C622 VTAIL.n552 B 0.034326f
C623 VTAIL.n553 B 1.25183f
C624 VTAIL.n554 B 0.031312f
C625 VTAIL.n555 B 0.021453f
C626 VTAIL.n556 B 0.011528f
C627 VTAIL.n557 B 0.027248f
C628 VTAIL.n558 B 0.012206f
C629 VTAIL.n559 B 0.021453f
C630 VTAIL.n560 B 0.011528f
C631 VTAIL.n561 B 0.027248f
C632 VTAIL.n562 B 0.012206f
C633 VTAIL.n563 B 0.021453f
C634 VTAIL.n564 B 0.011528f
C635 VTAIL.n565 B 0.027248f
C636 VTAIL.n566 B 0.012206f
C637 VTAIL.n567 B 0.021453f
C638 VTAIL.n568 B 0.011867f
C639 VTAIL.n569 B 0.027248f
C640 VTAIL.n570 B 0.012206f
C641 VTAIL.n571 B 0.021453f
C642 VTAIL.n572 B 0.011528f
C643 VTAIL.n573 B 0.027248f
C644 VTAIL.n574 B 0.012206f
C645 VTAIL.n575 B 0.021453f
C646 VTAIL.n576 B 0.011528f
C647 VTAIL.n577 B 0.020436f
C648 VTAIL.n578 B 0.019262f
C649 VTAIL.t12 B 0.046279f
C650 VTAIL.n579 B 0.173125f
C651 VTAIL.n580 B 1.29603f
C652 VTAIL.n581 B 0.011528f
C653 VTAIL.n582 B 0.012206f
C654 VTAIL.n583 B 0.027248f
C655 VTAIL.n584 B 0.027248f
C656 VTAIL.n585 B 0.012206f
C657 VTAIL.n586 B 0.011528f
C658 VTAIL.n587 B 0.021453f
C659 VTAIL.n588 B 0.021453f
C660 VTAIL.n589 B 0.011528f
C661 VTAIL.n590 B 0.012206f
C662 VTAIL.n591 B 0.027248f
C663 VTAIL.n592 B 0.027248f
C664 VTAIL.n593 B 0.012206f
C665 VTAIL.n594 B 0.011528f
C666 VTAIL.n595 B 0.021453f
C667 VTAIL.n596 B 0.021453f
C668 VTAIL.n597 B 0.011528f
C669 VTAIL.n598 B 0.011528f
C670 VTAIL.n599 B 0.012206f
C671 VTAIL.n600 B 0.027248f
C672 VTAIL.n601 B 0.027248f
C673 VTAIL.n602 B 0.027248f
C674 VTAIL.n603 B 0.011867f
C675 VTAIL.n604 B 0.011528f
C676 VTAIL.n605 B 0.021453f
C677 VTAIL.n606 B 0.021453f
C678 VTAIL.n607 B 0.011528f
C679 VTAIL.n608 B 0.012206f
C680 VTAIL.n609 B 0.027248f
C681 VTAIL.n610 B 0.027248f
C682 VTAIL.n611 B 0.012206f
C683 VTAIL.n612 B 0.011528f
C684 VTAIL.n613 B 0.021453f
C685 VTAIL.n614 B 0.021453f
C686 VTAIL.n615 B 0.011528f
C687 VTAIL.n616 B 0.012206f
C688 VTAIL.n617 B 0.027248f
C689 VTAIL.n618 B 0.027248f
C690 VTAIL.n619 B 0.012206f
C691 VTAIL.n620 B 0.011528f
C692 VTAIL.n621 B 0.021453f
C693 VTAIL.n622 B 0.021453f
C694 VTAIL.n623 B 0.011528f
C695 VTAIL.n624 B 0.012206f
C696 VTAIL.n625 B 0.027248f
C697 VTAIL.n626 B 0.061035f
C698 VTAIL.n627 B 0.012206f
C699 VTAIL.n628 B 0.011528f
C700 VTAIL.n629 B 0.048416f
C701 VTAIL.n630 B 0.034326f
C702 VTAIL.n631 B 1.24781f
C703 VDD2.t5 B 0.338435f
C704 VDD2.t4 B 0.338435f
C705 VDD2.n0 B 3.04477f
C706 VDD2.t1 B 0.338435f
C707 VDD2.t3 B 0.338435f
C708 VDD2.n1 B 3.04477f
C709 VDD2.n2 B 2.62165f
C710 VDD2.t6 B 0.338435f
C711 VDD2.t2 B 0.338435f
C712 VDD2.n3 B 3.04308f
C713 VDD2.n4 B 2.86999f
C714 VDD2.t7 B 0.338435f
C715 VDD2.t0 B 0.338435f
C716 VDD2.n5 B 3.04474f
C717 VN.n0 B 0.050348f
C718 VN.t1 B 0.938317f
C719 VN.n1 B 0.374609f
C720 VN.t0 B 0.947402f
C721 VN.n2 B 0.360771f
C722 VN.n3 B 0.160919f
C723 VN.n4 B 0.011425f
C724 VN.t7 B 0.938317f
C725 VN.n5 B 0.374609f
C726 VN.t2 B 0.938317f
C727 VN.n6 B 0.369487f
C728 VN.n7 B 0.039018f
C729 VN.n8 B 0.050348f
C730 VN.t6 B 0.938317f
C731 VN.n9 B 0.374609f
C732 VN.t5 B 0.947402f
C733 VN.n10 B 0.360771f
C734 VN.n11 B 0.160919f
C735 VN.n12 B 0.011425f
C736 VN.t3 B 0.938317f
C737 VN.n13 B 0.374609f
C738 VN.t4 B 0.938317f
C739 VN.n14 B 0.369487f
C740 VN.n15 B 2.16194f
.ends

