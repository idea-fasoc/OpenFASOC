* NGSPICE file created from diff_pair_sample_0113.ext - technology: sky130A

.subckt diff_pair_sample_0113 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=0 ps=0 w=12.13 l=3.17
X1 B.t8 B.t6 B.t7 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=0 ps=0 w=12.13 l=3.17
X2 B.t5 B.t3 B.t4 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=0 ps=0 w=12.13 l=3.17
X3 VDD1.t7 VP.t0 VTAIL.t9 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=4.7307 ps=25.04 w=12.13 l=3.17
X4 B.t2 B.t0 B.t1 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=0 ps=0 w=12.13 l=3.17
X5 VDD1.t6 VP.t1 VTAIL.t15 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X6 VTAIL.t4 VN.t0 VDD2.t7 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X7 VDD2.t6 VN.t1 VTAIL.t0 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X8 VDD2.t5 VN.t2 VTAIL.t6 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X9 VDD2.t4 VN.t3 VTAIL.t3 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=4.7307 ps=25.04 w=12.13 l=3.17
X10 VTAIL.t11 VP.t2 VDD1.t5 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=2.00145 ps=12.46 w=12.13 l=3.17
X11 VTAIL.t12 VP.t3 VDD1.t4 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X12 VTAIL.t5 VN.t4 VDD2.t3 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X13 VDD1.t3 VP.t4 VTAIL.t13 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X14 VDD1.t2 VP.t5 VTAIL.t14 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=4.7307 ps=25.04 w=12.13 l=3.17
X15 VDD2.t2 VN.t5 VTAIL.t2 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=4.7307 ps=25.04 w=12.13 l=3.17
X16 VTAIL.t8 VP.t6 VDD1.t1 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=2.00145 pd=12.46 as=2.00145 ps=12.46 w=12.13 l=3.17
X17 VTAIL.t10 VP.t7 VDD1.t0 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=2.00145 ps=12.46 w=12.13 l=3.17
X18 VTAIL.t7 VN.t6 VDD2.t1 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=2.00145 ps=12.46 w=12.13 l=3.17
X19 VTAIL.t1 VN.t7 VDD2.t0 w_n4470_n3394# sky130_fd_pr__pfet_01v8 ad=4.7307 pd=25.04 as=2.00145 ps=12.46 w=12.13 l=3.17
R0 B.n453 B.n452 585
R1 B.n451 B.n144 585
R2 B.n450 B.n449 585
R3 B.n448 B.n145 585
R4 B.n447 B.n446 585
R5 B.n445 B.n146 585
R6 B.n444 B.n443 585
R7 B.n442 B.n147 585
R8 B.n441 B.n440 585
R9 B.n439 B.n148 585
R10 B.n438 B.n437 585
R11 B.n436 B.n149 585
R12 B.n435 B.n434 585
R13 B.n433 B.n150 585
R14 B.n432 B.n431 585
R15 B.n430 B.n151 585
R16 B.n429 B.n428 585
R17 B.n427 B.n152 585
R18 B.n426 B.n425 585
R19 B.n424 B.n153 585
R20 B.n423 B.n422 585
R21 B.n421 B.n154 585
R22 B.n420 B.n419 585
R23 B.n418 B.n155 585
R24 B.n417 B.n416 585
R25 B.n415 B.n156 585
R26 B.n414 B.n413 585
R27 B.n412 B.n157 585
R28 B.n411 B.n410 585
R29 B.n409 B.n158 585
R30 B.n408 B.n407 585
R31 B.n406 B.n159 585
R32 B.n405 B.n404 585
R33 B.n403 B.n160 585
R34 B.n402 B.n401 585
R35 B.n400 B.n161 585
R36 B.n399 B.n398 585
R37 B.n397 B.n162 585
R38 B.n396 B.n395 585
R39 B.n394 B.n163 585
R40 B.n393 B.n392 585
R41 B.n391 B.n164 585
R42 B.n389 B.n388 585
R43 B.n387 B.n167 585
R44 B.n386 B.n385 585
R45 B.n384 B.n168 585
R46 B.n383 B.n382 585
R47 B.n381 B.n169 585
R48 B.n380 B.n379 585
R49 B.n378 B.n170 585
R50 B.n377 B.n376 585
R51 B.n375 B.n171 585
R52 B.n374 B.n373 585
R53 B.n369 B.n172 585
R54 B.n368 B.n367 585
R55 B.n366 B.n173 585
R56 B.n365 B.n364 585
R57 B.n363 B.n174 585
R58 B.n362 B.n361 585
R59 B.n360 B.n175 585
R60 B.n359 B.n358 585
R61 B.n357 B.n176 585
R62 B.n356 B.n355 585
R63 B.n354 B.n177 585
R64 B.n353 B.n352 585
R65 B.n351 B.n178 585
R66 B.n350 B.n349 585
R67 B.n348 B.n179 585
R68 B.n347 B.n346 585
R69 B.n345 B.n180 585
R70 B.n344 B.n343 585
R71 B.n342 B.n181 585
R72 B.n341 B.n340 585
R73 B.n339 B.n182 585
R74 B.n338 B.n337 585
R75 B.n336 B.n183 585
R76 B.n335 B.n334 585
R77 B.n333 B.n184 585
R78 B.n332 B.n331 585
R79 B.n330 B.n185 585
R80 B.n329 B.n328 585
R81 B.n327 B.n186 585
R82 B.n326 B.n325 585
R83 B.n324 B.n187 585
R84 B.n323 B.n322 585
R85 B.n321 B.n188 585
R86 B.n320 B.n319 585
R87 B.n318 B.n189 585
R88 B.n317 B.n316 585
R89 B.n315 B.n190 585
R90 B.n314 B.n313 585
R91 B.n312 B.n191 585
R92 B.n311 B.n310 585
R93 B.n309 B.n192 585
R94 B.n454 B.n143 585
R95 B.n456 B.n455 585
R96 B.n457 B.n142 585
R97 B.n459 B.n458 585
R98 B.n460 B.n141 585
R99 B.n462 B.n461 585
R100 B.n463 B.n140 585
R101 B.n465 B.n464 585
R102 B.n466 B.n139 585
R103 B.n468 B.n467 585
R104 B.n469 B.n138 585
R105 B.n471 B.n470 585
R106 B.n472 B.n137 585
R107 B.n474 B.n473 585
R108 B.n475 B.n136 585
R109 B.n477 B.n476 585
R110 B.n478 B.n135 585
R111 B.n480 B.n479 585
R112 B.n481 B.n134 585
R113 B.n483 B.n482 585
R114 B.n484 B.n133 585
R115 B.n486 B.n485 585
R116 B.n487 B.n132 585
R117 B.n489 B.n488 585
R118 B.n490 B.n131 585
R119 B.n492 B.n491 585
R120 B.n493 B.n130 585
R121 B.n495 B.n494 585
R122 B.n496 B.n129 585
R123 B.n498 B.n497 585
R124 B.n499 B.n128 585
R125 B.n501 B.n500 585
R126 B.n502 B.n127 585
R127 B.n504 B.n503 585
R128 B.n505 B.n126 585
R129 B.n507 B.n506 585
R130 B.n508 B.n125 585
R131 B.n510 B.n509 585
R132 B.n511 B.n124 585
R133 B.n513 B.n512 585
R134 B.n514 B.n123 585
R135 B.n516 B.n515 585
R136 B.n517 B.n122 585
R137 B.n519 B.n518 585
R138 B.n520 B.n121 585
R139 B.n522 B.n521 585
R140 B.n523 B.n120 585
R141 B.n525 B.n524 585
R142 B.n526 B.n119 585
R143 B.n528 B.n527 585
R144 B.n529 B.n118 585
R145 B.n531 B.n530 585
R146 B.n532 B.n117 585
R147 B.n534 B.n533 585
R148 B.n535 B.n116 585
R149 B.n537 B.n536 585
R150 B.n538 B.n115 585
R151 B.n540 B.n539 585
R152 B.n541 B.n114 585
R153 B.n543 B.n542 585
R154 B.n544 B.n113 585
R155 B.n546 B.n545 585
R156 B.n547 B.n112 585
R157 B.n549 B.n548 585
R158 B.n550 B.n111 585
R159 B.n552 B.n551 585
R160 B.n553 B.n110 585
R161 B.n555 B.n554 585
R162 B.n556 B.n109 585
R163 B.n558 B.n557 585
R164 B.n559 B.n108 585
R165 B.n561 B.n560 585
R166 B.n562 B.n107 585
R167 B.n564 B.n563 585
R168 B.n565 B.n106 585
R169 B.n567 B.n566 585
R170 B.n568 B.n105 585
R171 B.n570 B.n569 585
R172 B.n571 B.n104 585
R173 B.n573 B.n572 585
R174 B.n574 B.n103 585
R175 B.n576 B.n575 585
R176 B.n577 B.n102 585
R177 B.n579 B.n578 585
R178 B.n580 B.n101 585
R179 B.n582 B.n581 585
R180 B.n583 B.n100 585
R181 B.n585 B.n584 585
R182 B.n586 B.n99 585
R183 B.n588 B.n587 585
R184 B.n589 B.n98 585
R185 B.n591 B.n590 585
R186 B.n592 B.n97 585
R187 B.n594 B.n593 585
R188 B.n595 B.n96 585
R189 B.n597 B.n596 585
R190 B.n598 B.n95 585
R191 B.n600 B.n599 585
R192 B.n601 B.n94 585
R193 B.n603 B.n602 585
R194 B.n604 B.n93 585
R195 B.n606 B.n605 585
R196 B.n607 B.n92 585
R197 B.n609 B.n608 585
R198 B.n610 B.n91 585
R199 B.n612 B.n611 585
R200 B.n613 B.n90 585
R201 B.n615 B.n614 585
R202 B.n616 B.n89 585
R203 B.n618 B.n617 585
R204 B.n619 B.n88 585
R205 B.n621 B.n620 585
R206 B.n622 B.n87 585
R207 B.n624 B.n623 585
R208 B.n625 B.n86 585
R209 B.n627 B.n626 585
R210 B.n628 B.n85 585
R211 B.n630 B.n629 585
R212 B.n631 B.n84 585
R213 B.n633 B.n632 585
R214 B.n775 B.n774 585
R215 B.n773 B.n32 585
R216 B.n772 B.n771 585
R217 B.n770 B.n33 585
R218 B.n769 B.n768 585
R219 B.n767 B.n34 585
R220 B.n766 B.n765 585
R221 B.n764 B.n35 585
R222 B.n763 B.n762 585
R223 B.n761 B.n36 585
R224 B.n760 B.n759 585
R225 B.n758 B.n37 585
R226 B.n757 B.n756 585
R227 B.n755 B.n38 585
R228 B.n754 B.n753 585
R229 B.n752 B.n39 585
R230 B.n751 B.n750 585
R231 B.n749 B.n40 585
R232 B.n748 B.n747 585
R233 B.n746 B.n41 585
R234 B.n745 B.n744 585
R235 B.n743 B.n42 585
R236 B.n742 B.n741 585
R237 B.n740 B.n43 585
R238 B.n739 B.n738 585
R239 B.n737 B.n44 585
R240 B.n736 B.n735 585
R241 B.n734 B.n45 585
R242 B.n733 B.n732 585
R243 B.n731 B.n46 585
R244 B.n730 B.n729 585
R245 B.n728 B.n47 585
R246 B.n727 B.n726 585
R247 B.n725 B.n48 585
R248 B.n724 B.n723 585
R249 B.n722 B.n49 585
R250 B.n721 B.n720 585
R251 B.n719 B.n50 585
R252 B.n718 B.n717 585
R253 B.n716 B.n51 585
R254 B.n715 B.n714 585
R255 B.n713 B.n52 585
R256 B.n712 B.n711 585
R257 B.n710 B.n53 585
R258 B.n709 B.n708 585
R259 B.n707 B.n57 585
R260 B.n706 B.n705 585
R261 B.n704 B.n58 585
R262 B.n703 B.n702 585
R263 B.n701 B.n59 585
R264 B.n700 B.n699 585
R265 B.n698 B.n60 585
R266 B.n696 B.n695 585
R267 B.n694 B.n63 585
R268 B.n693 B.n692 585
R269 B.n691 B.n64 585
R270 B.n690 B.n689 585
R271 B.n688 B.n65 585
R272 B.n687 B.n686 585
R273 B.n685 B.n66 585
R274 B.n684 B.n683 585
R275 B.n682 B.n67 585
R276 B.n681 B.n680 585
R277 B.n679 B.n68 585
R278 B.n678 B.n677 585
R279 B.n676 B.n69 585
R280 B.n675 B.n674 585
R281 B.n673 B.n70 585
R282 B.n672 B.n671 585
R283 B.n670 B.n71 585
R284 B.n669 B.n668 585
R285 B.n667 B.n72 585
R286 B.n666 B.n665 585
R287 B.n664 B.n73 585
R288 B.n663 B.n662 585
R289 B.n661 B.n74 585
R290 B.n660 B.n659 585
R291 B.n658 B.n75 585
R292 B.n657 B.n656 585
R293 B.n655 B.n76 585
R294 B.n654 B.n653 585
R295 B.n652 B.n77 585
R296 B.n651 B.n650 585
R297 B.n649 B.n78 585
R298 B.n648 B.n647 585
R299 B.n646 B.n79 585
R300 B.n645 B.n644 585
R301 B.n643 B.n80 585
R302 B.n642 B.n641 585
R303 B.n640 B.n81 585
R304 B.n639 B.n638 585
R305 B.n637 B.n82 585
R306 B.n636 B.n635 585
R307 B.n634 B.n83 585
R308 B.n776 B.n31 585
R309 B.n778 B.n777 585
R310 B.n779 B.n30 585
R311 B.n781 B.n780 585
R312 B.n782 B.n29 585
R313 B.n784 B.n783 585
R314 B.n785 B.n28 585
R315 B.n787 B.n786 585
R316 B.n788 B.n27 585
R317 B.n790 B.n789 585
R318 B.n791 B.n26 585
R319 B.n793 B.n792 585
R320 B.n794 B.n25 585
R321 B.n796 B.n795 585
R322 B.n797 B.n24 585
R323 B.n799 B.n798 585
R324 B.n800 B.n23 585
R325 B.n802 B.n801 585
R326 B.n803 B.n22 585
R327 B.n805 B.n804 585
R328 B.n806 B.n21 585
R329 B.n808 B.n807 585
R330 B.n809 B.n20 585
R331 B.n811 B.n810 585
R332 B.n812 B.n19 585
R333 B.n814 B.n813 585
R334 B.n815 B.n18 585
R335 B.n817 B.n816 585
R336 B.n818 B.n17 585
R337 B.n820 B.n819 585
R338 B.n821 B.n16 585
R339 B.n823 B.n822 585
R340 B.n824 B.n15 585
R341 B.n826 B.n825 585
R342 B.n827 B.n14 585
R343 B.n829 B.n828 585
R344 B.n830 B.n13 585
R345 B.n832 B.n831 585
R346 B.n833 B.n12 585
R347 B.n835 B.n834 585
R348 B.n836 B.n11 585
R349 B.n838 B.n837 585
R350 B.n839 B.n10 585
R351 B.n841 B.n840 585
R352 B.n842 B.n9 585
R353 B.n844 B.n843 585
R354 B.n845 B.n8 585
R355 B.n847 B.n846 585
R356 B.n848 B.n7 585
R357 B.n850 B.n849 585
R358 B.n851 B.n6 585
R359 B.n853 B.n852 585
R360 B.n854 B.n5 585
R361 B.n856 B.n855 585
R362 B.n857 B.n4 585
R363 B.n859 B.n858 585
R364 B.n860 B.n3 585
R365 B.n862 B.n861 585
R366 B.n863 B.n0 585
R367 B.n2 B.n1 585
R368 B.n222 B.n221 585
R369 B.n224 B.n223 585
R370 B.n225 B.n220 585
R371 B.n227 B.n226 585
R372 B.n228 B.n219 585
R373 B.n230 B.n229 585
R374 B.n231 B.n218 585
R375 B.n233 B.n232 585
R376 B.n234 B.n217 585
R377 B.n236 B.n235 585
R378 B.n237 B.n216 585
R379 B.n239 B.n238 585
R380 B.n240 B.n215 585
R381 B.n242 B.n241 585
R382 B.n243 B.n214 585
R383 B.n245 B.n244 585
R384 B.n246 B.n213 585
R385 B.n248 B.n247 585
R386 B.n249 B.n212 585
R387 B.n251 B.n250 585
R388 B.n252 B.n211 585
R389 B.n254 B.n253 585
R390 B.n255 B.n210 585
R391 B.n257 B.n256 585
R392 B.n258 B.n209 585
R393 B.n260 B.n259 585
R394 B.n261 B.n208 585
R395 B.n263 B.n262 585
R396 B.n264 B.n207 585
R397 B.n266 B.n265 585
R398 B.n267 B.n206 585
R399 B.n269 B.n268 585
R400 B.n270 B.n205 585
R401 B.n272 B.n271 585
R402 B.n273 B.n204 585
R403 B.n275 B.n274 585
R404 B.n276 B.n203 585
R405 B.n278 B.n277 585
R406 B.n279 B.n202 585
R407 B.n281 B.n280 585
R408 B.n282 B.n201 585
R409 B.n284 B.n283 585
R410 B.n285 B.n200 585
R411 B.n287 B.n286 585
R412 B.n288 B.n199 585
R413 B.n290 B.n289 585
R414 B.n291 B.n198 585
R415 B.n293 B.n292 585
R416 B.n294 B.n197 585
R417 B.n296 B.n295 585
R418 B.n297 B.n196 585
R419 B.n299 B.n298 585
R420 B.n300 B.n195 585
R421 B.n302 B.n301 585
R422 B.n303 B.n194 585
R423 B.n305 B.n304 585
R424 B.n306 B.n193 585
R425 B.n308 B.n307 585
R426 B.n307 B.n192 478.086
R427 B.n454 B.n453 478.086
R428 B.n634 B.n633 478.086
R429 B.n774 B.n31 478.086
R430 B.n165 B.t7 445.93
R431 B.n61 B.t5 445.93
R432 B.n370 B.t10 445.93
R433 B.n54 B.t2 445.93
R434 B.n166 B.t8 378.051
R435 B.n62 B.t4 378.051
R436 B.n371 B.t11 378.051
R437 B.n55 B.t1 378.051
R438 B.n370 B.t9 300.99
R439 B.n165 B.t6 300.99
R440 B.n61 B.t3 300.99
R441 B.n54 B.t0 300.99
R442 B.n865 B.n864 256.663
R443 B.n864 B.n863 235.042
R444 B.n864 B.n2 235.042
R445 B.n311 B.n192 163.367
R446 B.n312 B.n311 163.367
R447 B.n313 B.n312 163.367
R448 B.n313 B.n190 163.367
R449 B.n317 B.n190 163.367
R450 B.n318 B.n317 163.367
R451 B.n319 B.n318 163.367
R452 B.n319 B.n188 163.367
R453 B.n323 B.n188 163.367
R454 B.n324 B.n323 163.367
R455 B.n325 B.n324 163.367
R456 B.n325 B.n186 163.367
R457 B.n329 B.n186 163.367
R458 B.n330 B.n329 163.367
R459 B.n331 B.n330 163.367
R460 B.n331 B.n184 163.367
R461 B.n335 B.n184 163.367
R462 B.n336 B.n335 163.367
R463 B.n337 B.n336 163.367
R464 B.n337 B.n182 163.367
R465 B.n341 B.n182 163.367
R466 B.n342 B.n341 163.367
R467 B.n343 B.n342 163.367
R468 B.n343 B.n180 163.367
R469 B.n347 B.n180 163.367
R470 B.n348 B.n347 163.367
R471 B.n349 B.n348 163.367
R472 B.n349 B.n178 163.367
R473 B.n353 B.n178 163.367
R474 B.n354 B.n353 163.367
R475 B.n355 B.n354 163.367
R476 B.n355 B.n176 163.367
R477 B.n359 B.n176 163.367
R478 B.n360 B.n359 163.367
R479 B.n361 B.n360 163.367
R480 B.n361 B.n174 163.367
R481 B.n365 B.n174 163.367
R482 B.n366 B.n365 163.367
R483 B.n367 B.n366 163.367
R484 B.n367 B.n172 163.367
R485 B.n374 B.n172 163.367
R486 B.n375 B.n374 163.367
R487 B.n376 B.n375 163.367
R488 B.n376 B.n170 163.367
R489 B.n380 B.n170 163.367
R490 B.n381 B.n380 163.367
R491 B.n382 B.n381 163.367
R492 B.n382 B.n168 163.367
R493 B.n386 B.n168 163.367
R494 B.n387 B.n386 163.367
R495 B.n388 B.n387 163.367
R496 B.n388 B.n164 163.367
R497 B.n393 B.n164 163.367
R498 B.n394 B.n393 163.367
R499 B.n395 B.n394 163.367
R500 B.n395 B.n162 163.367
R501 B.n399 B.n162 163.367
R502 B.n400 B.n399 163.367
R503 B.n401 B.n400 163.367
R504 B.n401 B.n160 163.367
R505 B.n405 B.n160 163.367
R506 B.n406 B.n405 163.367
R507 B.n407 B.n406 163.367
R508 B.n407 B.n158 163.367
R509 B.n411 B.n158 163.367
R510 B.n412 B.n411 163.367
R511 B.n413 B.n412 163.367
R512 B.n413 B.n156 163.367
R513 B.n417 B.n156 163.367
R514 B.n418 B.n417 163.367
R515 B.n419 B.n418 163.367
R516 B.n419 B.n154 163.367
R517 B.n423 B.n154 163.367
R518 B.n424 B.n423 163.367
R519 B.n425 B.n424 163.367
R520 B.n425 B.n152 163.367
R521 B.n429 B.n152 163.367
R522 B.n430 B.n429 163.367
R523 B.n431 B.n430 163.367
R524 B.n431 B.n150 163.367
R525 B.n435 B.n150 163.367
R526 B.n436 B.n435 163.367
R527 B.n437 B.n436 163.367
R528 B.n437 B.n148 163.367
R529 B.n441 B.n148 163.367
R530 B.n442 B.n441 163.367
R531 B.n443 B.n442 163.367
R532 B.n443 B.n146 163.367
R533 B.n447 B.n146 163.367
R534 B.n448 B.n447 163.367
R535 B.n449 B.n448 163.367
R536 B.n449 B.n144 163.367
R537 B.n453 B.n144 163.367
R538 B.n633 B.n84 163.367
R539 B.n629 B.n84 163.367
R540 B.n629 B.n628 163.367
R541 B.n628 B.n627 163.367
R542 B.n627 B.n86 163.367
R543 B.n623 B.n86 163.367
R544 B.n623 B.n622 163.367
R545 B.n622 B.n621 163.367
R546 B.n621 B.n88 163.367
R547 B.n617 B.n88 163.367
R548 B.n617 B.n616 163.367
R549 B.n616 B.n615 163.367
R550 B.n615 B.n90 163.367
R551 B.n611 B.n90 163.367
R552 B.n611 B.n610 163.367
R553 B.n610 B.n609 163.367
R554 B.n609 B.n92 163.367
R555 B.n605 B.n92 163.367
R556 B.n605 B.n604 163.367
R557 B.n604 B.n603 163.367
R558 B.n603 B.n94 163.367
R559 B.n599 B.n94 163.367
R560 B.n599 B.n598 163.367
R561 B.n598 B.n597 163.367
R562 B.n597 B.n96 163.367
R563 B.n593 B.n96 163.367
R564 B.n593 B.n592 163.367
R565 B.n592 B.n591 163.367
R566 B.n591 B.n98 163.367
R567 B.n587 B.n98 163.367
R568 B.n587 B.n586 163.367
R569 B.n586 B.n585 163.367
R570 B.n585 B.n100 163.367
R571 B.n581 B.n100 163.367
R572 B.n581 B.n580 163.367
R573 B.n580 B.n579 163.367
R574 B.n579 B.n102 163.367
R575 B.n575 B.n102 163.367
R576 B.n575 B.n574 163.367
R577 B.n574 B.n573 163.367
R578 B.n573 B.n104 163.367
R579 B.n569 B.n104 163.367
R580 B.n569 B.n568 163.367
R581 B.n568 B.n567 163.367
R582 B.n567 B.n106 163.367
R583 B.n563 B.n106 163.367
R584 B.n563 B.n562 163.367
R585 B.n562 B.n561 163.367
R586 B.n561 B.n108 163.367
R587 B.n557 B.n108 163.367
R588 B.n557 B.n556 163.367
R589 B.n556 B.n555 163.367
R590 B.n555 B.n110 163.367
R591 B.n551 B.n110 163.367
R592 B.n551 B.n550 163.367
R593 B.n550 B.n549 163.367
R594 B.n549 B.n112 163.367
R595 B.n545 B.n112 163.367
R596 B.n545 B.n544 163.367
R597 B.n544 B.n543 163.367
R598 B.n543 B.n114 163.367
R599 B.n539 B.n114 163.367
R600 B.n539 B.n538 163.367
R601 B.n538 B.n537 163.367
R602 B.n537 B.n116 163.367
R603 B.n533 B.n116 163.367
R604 B.n533 B.n532 163.367
R605 B.n532 B.n531 163.367
R606 B.n531 B.n118 163.367
R607 B.n527 B.n118 163.367
R608 B.n527 B.n526 163.367
R609 B.n526 B.n525 163.367
R610 B.n525 B.n120 163.367
R611 B.n521 B.n120 163.367
R612 B.n521 B.n520 163.367
R613 B.n520 B.n519 163.367
R614 B.n519 B.n122 163.367
R615 B.n515 B.n122 163.367
R616 B.n515 B.n514 163.367
R617 B.n514 B.n513 163.367
R618 B.n513 B.n124 163.367
R619 B.n509 B.n124 163.367
R620 B.n509 B.n508 163.367
R621 B.n508 B.n507 163.367
R622 B.n507 B.n126 163.367
R623 B.n503 B.n126 163.367
R624 B.n503 B.n502 163.367
R625 B.n502 B.n501 163.367
R626 B.n501 B.n128 163.367
R627 B.n497 B.n128 163.367
R628 B.n497 B.n496 163.367
R629 B.n496 B.n495 163.367
R630 B.n495 B.n130 163.367
R631 B.n491 B.n130 163.367
R632 B.n491 B.n490 163.367
R633 B.n490 B.n489 163.367
R634 B.n489 B.n132 163.367
R635 B.n485 B.n132 163.367
R636 B.n485 B.n484 163.367
R637 B.n484 B.n483 163.367
R638 B.n483 B.n134 163.367
R639 B.n479 B.n134 163.367
R640 B.n479 B.n478 163.367
R641 B.n478 B.n477 163.367
R642 B.n477 B.n136 163.367
R643 B.n473 B.n136 163.367
R644 B.n473 B.n472 163.367
R645 B.n472 B.n471 163.367
R646 B.n471 B.n138 163.367
R647 B.n467 B.n138 163.367
R648 B.n467 B.n466 163.367
R649 B.n466 B.n465 163.367
R650 B.n465 B.n140 163.367
R651 B.n461 B.n140 163.367
R652 B.n461 B.n460 163.367
R653 B.n460 B.n459 163.367
R654 B.n459 B.n142 163.367
R655 B.n455 B.n142 163.367
R656 B.n455 B.n454 163.367
R657 B.n774 B.n773 163.367
R658 B.n773 B.n772 163.367
R659 B.n772 B.n33 163.367
R660 B.n768 B.n33 163.367
R661 B.n768 B.n767 163.367
R662 B.n767 B.n766 163.367
R663 B.n766 B.n35 163.367
R664 B.n762 B.n35 163.367
R665 B.n762 B.n761 163.367
R666 B.n761 B.n760 163.367
R667 B.n760 B.n37 163.367
R668 B.n756 B.n37 163.367
R669 B.n756 B.n755 163.367
R670 B.n755 B.n754 163.367
R671 B.n754 B.n39 163.367
R672 B.n750 B.n39 163.367
R673 B.n750 B.n749 163.367
R674 B.n749 B.n748 163.367
R675 B.n748 B.n41 163.367
R676 B.n744 B.n41 163.367
R677 B.n744 B.n743 163.367
R678 B.n743 B.n742 163.367
R679 B.n742 B.n43 163.367
R680 B.n738 B.n43 163.367
R681 B.n738 B.n737 163.367
R682 B.n737 B.n736 163.367
R683 B.n736 B.n45 163.367
R684 B.n732 B.n45 163.367
R685 B.n732 B.n731 163.367
R686 B.n731 B.n730 163.367
R687 B.n730 B.n47 163.367
R688 B.n726 B.n47 163.367
R689 B.n726 B.n725 163.367
R690 B.n725 B.n724 163.367
R691 B.n724 B.n49 163.367
R692 B.n720 B.n49 163.367
R693 B.n720 B.n719 163.367
R694 B.n719 B.n718 163.367
R695 B.n718 B.n51 163.367
R696 B.n714 B.n51 163.367
R697 B.n714 B.n713 163.367
R698 B.n713 B.n712 163.367
R699 B.n712 B.n53 163.367
R700 B.n708 B.n53 163.367
R701 B.n708 B.n707 163.367
R702 B.n707 B.n706 163.367
R703 B.n706 B.n58 163.367
R704 B.n702 B.n58 163.367
R705 B.n702 B.n701 163.367
R706 B.n701 B.n700 163.367
R707 B.n700 B.n60 163.367
R708 B.n695 B.n60 163.367
R709 B.n695 B.n694 163.367
R710 B.n694 B.n693 163.367
R711 B.n693 B.n64 163.367
R712 B.n689 B.n64 163.367
R713 B.n689 B.n688 163.367
R714 B.n688 B.n687 163.367
R715 B.n687 B.n66 163.367
R716 B.n683 B.n66 163.367
R717 B.n683 B.n682 163.367
R718 B.n682 B.n681 163.367
R719 B.n681 B.n68 163.367
R720 B.n677 B.n68 163.367
R721 B.n677 B.n676 163.367
R722 B.n676 B.n675 163.367
R723 B.n675 B.n70 163.367
R724 B.n671 B.n70 163.367
R725 B.n671 B.n670 163.367
R726 B.n670 B.n669 163.367
R727 B.n669 B.n72 163.367
R728 B.n665 B.n72 163.367
R729 B.n665 B.n664 163.367
R730 B.n664 B.n663 163.367
R731 B.n663 B.n74 163.367
R732 B.n659 B.n74 163.367
R733 B.n659 B.n658 163.367
R734 B.n658 B.n657 163.367
R735 B.n657 B.n76 163.367
R736 B.n653 B.n76 163.367
R737 B.n653 B.n652 163.367
R738 B.n652 B.n651 163.367
R739 B.n651 B.n78 163.367
R740 B.n647 B.n78 163.367
R741 B.n647 B.n646 163.367
R742 B.n646 B.n645 163.367
R743 B.n645 B.n80 163.367
R744 B.n641 B.n80 163.367
R745 B.n641 B.n640 163.367
R746 B.n640 B.n639 163.367
R747 B.n639 B.n82 163.367
R748 B.n635 B.n82 163.367
R749 B.n635 B.n634 163.367
R750 B.n778 B.n31 163.367
R751 B.n779 B.n778 163.367
R752 B.n780 B.n779 163.367
R753 B.n780 B.n29 163.367
R754 B.n784 B.n29 163.367
R755 B.n785 B.n784 163.367
R756 B.n786 B.n785 163.367
R757 B.n786 B.n27 163.367
R758 B.n790 B.n27 163.367
R759 B.n791 B.n790 163.367
R760 B.n792 B.n791 163.367
R761 B.n792 B.n25 163.367
R762 B.n796 B.n25 163.367
R763 B.n797 B.n796 163.367
R764 B.n798 B.n797 163.367
R765 B.n798 B.n23 163.367
R766 B.n802 B.n23 163.367
R767 B.n803 B.n802 163.367
R768 B.n804 B.n803 163.367
R769 B.n804 B.n21 163.367
R770 B.n808 B.n21 163.367
R771 B.n809 B.n808 163.367
R772 B.n810 B.n809 163.367
R773 B.n810 B.n19 163.367
R774 B.n814 B.n19 163.367
R775 B.n815 B.n814 163.367
R776 B.n816 B.n815 163.367
R777 B.n816 B.n17 163.367
R778 B.n820 B.n17 163.367
R779 B.n821 B.n820 163.367
R780 B.n822 B.n821 163.367
R781 B.n822 B.n15 163.367
R782 B.n826 B.n15 163.367
R783 B.n827 B.n826 163.367
R784 B.n828 B.n827 163.367
R785 B.n828 B.n13 163.367
R786 B.n832 B.n13 163.367
R787 B.n833 B.n832 163.367
R788 B.n834 B.n833 163.367
R789 B.n834 B.n11 163.367
R790 B.n838 B.n11 163.367
R791 B.n839 B.n838 163.367
R792 B.n840 B.n839 163.367
R793 B.n840 B.n9 163.367
R794 B.n844 B.n9 163.367
R795 B.n845 B.n844 163.367
R796 B.n846 B.n845 163.367
R797 B.n846 B.n7 163.367
R798 B.n850 B.n7 163.367
R799 B.n851 B.n850 163.367
R800 B.n852 B.n851 163.367
R801 B.n852 B.n5 163.367
R802 B.n856 B.n5 163.367
R803 B.n857 B.n856 163.367
R804 B.n858 B.n857 163.367
R805 B.n858 B.n3 163.367
R806 B.n862 B.n3 163.367
R807 B.n863 B.n862 163.367
R808 B.n222 B.n2 163.367
R809 B.n223 B.n222 163.367
R810 B.n223 B.n220 163.367
R811 B.n227 B.n220 163.367
R812 B.n228 B.n227 163.367
R813 B.n229 B.n228 163.367
R814 B.n229 B.n218 163.367
R815 B.n233 B.n218 163.367
R816 B.n234 B.n233 163.367
R817 B.n235 B.n234 163.367
R818 B.n235 B.n216 163.367
R819 B.n239 B.n216 163.367
R820 B.n240 B.n239 163.367
R821 B.n241 B.n240 163.367
R822 B.n241 B.n214 163.367
R823 B.n245 B.n214 163.367
R824 B.n246 B.n245 163.367
R825 B.n247 B.n246 163.367
R826 B.n247 B.n212 163.367
R827 B.n251 B.n212 163.367
R828 B.n252 B.n251 163.367
R829 B.n253 B.n252 163.367
R830 B.n253 B.n210 163.367
R831 B.n257 B.n210 163.367
R832 B.n258 B.n257 163.367
R833 B.n259 B.n258 163.367
R834 B.n259 B.n208 163.367
R835 B.n263 B.n208 163.367
R836 B.n264 B.n263 163.367
R837 B.n265 B.n264 163.367
R838 B.n265 B.n206 163.367
R839 B.n269 B.n206 163.367
R840 B.n270 B.n269 163.367
R841 B.n271 B.n270 163.367
R842 B.n271 B.n204 163.367
R843 B.n275 B.n204 163.367
R844 B.n276 B.n275 163.367
R845 B.n277 B.n276 163.367
R846 B.n277 B.n202 163.367
R847 B.n281 B.n202 163.367
R848 B.n282 B.n281 163.367
R849 B.n283 B.n282 163.367
R850 B.n283 B.n200 163.367
R851 B.n287 B.n200 163.367
R852 B.n288 B.n287 163.367
R853 B.n289 B.n288 163.367
R854 B.n289 B.n198 163.367
R855 B.n293 B.n198 163.367
R856 B.n294 B.n293 163.367
R857 B.n295 B.n294 163.367
R858 B.n295 B.n196 163.367
R859 B.n299 B.n196 163.367
R860 B.n300 B.n299 163.367
R861 B.n301 B.n300 163.367
R862 B.n301 B.n194 163.367
R863 B.n305 B.n194 163.367
R864 B.n306 B.n305 163.367
R865 B.n307 B.n306 163.367
R866 B.n371 B.n370 67.8793
R867 B.n166 B.n165 67.8793
R868 B.n62 B.n61 67.8793
R869 B.n55 B.n54 67.8793
R870 B.n372 B.n371 59.5399
R871 B.n390 B.n166 59.5399
R872 B.n697 B.n62 59.5399
R873 B.n56 B.n55 59.5399
R874 B.n776 B.n775 31.0639
R875 B.n632 B.n83 31.0639
R876 B.n452 B.n143 31.0639
R877 B.n309 B.n308 31.0639
R878 B B.n865 18.0485
R879 B.n777 B.n776 10.6151
R880 B.n777 B.n30 10.6151
R881 B.n781 B.n30 10.6151
R882 B.n782 B.n781 10.6151
R883 B.n783 B.n782 10.6151
R884 B.n783 B.n28 10.6151
R885 B.n787 B.n28 10.6151
R886 B.n788 B.n787 10.6151
R887 B.n789 B.n788 10.6151
R888 B.n789 B.n26 10.6151
R889 B.n793 B.n26 10.6151
R890 B.n794 B.n793 10.6151
R891 B.n795 B.n794 10.6151
R892 B.n795 B.n24 10.6151
R893 B.n799 B.n24 10.6151
R894 B.n800 B.n799 10.6151
R895 B.n801 B.n800 10.6151
R896 B.n801 B.n22 10.6151
R897 B.n805 B.n22 10.6151
R898 B.n806 B.n805 10.6151
R899 B.n807 B.n806 10.6151
R900 B.n807 B.n20 10.6151
R901 B.n811 B.n20 10.6151
R902 B.n812 B.n811 10.6151
R903 B.n813 B.n812 10.6151
R904 B.n813 B.n18 10.6151
R905 B.n817 B.n18 10.6151
R906 B.n818 B.n817 10.6151
R907 B.n819 B.n818 10.6151
R908 B.n819 B.n16 10.6151
R909 B.n823 B.n16 10.6151
R910 B.n824 B.n823 10.6151
R911 B.n825 B.n824 10.6151
R912 B.n825 B.n14 10.6151
R913 B.n829 B.n14 10.6151
R914 B.n830 B.n829 10.6151
R915 B.n831 B.n830 10.6151
R916 B.n831 B.n12 10.6151
R917 B.n835 B.n12 10.6151
R918 B.n836 B.n835 10.6151
R919 B.n837 B.n836 10.6151
R920 B.n837 B.n10 10.6151
R921 B.n841 B.n10 10.6151
R922 B.n842 B.n841 10.6151
R923 B.n843 B.n842 10.6151
R924 B.n843 B.n8 10.6151
R925 B.n847 B.n8 10.6151
R926 B.n848 B.n847 10.6151
R927 B.n849 B.n848 10.6151
R928 B.n849 B.n6 10.6151
R929 B.n853 B.n6 10.6151
R930 B.n854 B.n853 10.6151
R931 B.n855 B.n854 10.6151
R932 B.n855 B.n4 10.6151
R933 B.n859 B.n4 10.6151
R934 B.n860 B.n859 10.6151
R935 B.n861 B.n860 10.6151
R936 B.n861 B.n0 10.6151
R937 B.n775 B.n32 10.6151
R938 B.n771 B.n32 10.6151
R939 B.n771 B.n770 10.6151
R940 B.n770 B.n769 10.6151
R941 B.n769 B.n34 10.6151
R942 B.n765 B.n34 10.6151
R943 B.n765 B.n764 10.6151
R944 B.n764 B.n763 10.6151
R945 B.n763 B.n36 10.6151
R946 B.n759 B.n36 10.6151
R947 B.n759 B.n758 10.6151
R948 B.n758 B.n757 10.6151
R949 B.n757 B.n38 10.6151
R950 B.n753 B.n38 10.6151
R951 B.n753 B.n752 10.6151
R952 B.n752 B.n751 10.6151
R953 B.n751 B.n40 10.6151
R954 B.n747 B.n40 10.6151
R955 B.n747 B.n746 10.6151
R956 B.n746 B.n745 10.6151
R957 B.n745 B.n42 10.6151
R958 B.n741 B.n42 10.6151
R959 B.n741 B.n740 10.6151
R960 B.n740 B.n739 10.6151
R961 B.n739 B.n44 10.6151
R962 B.n735 B.n44 10.6151
R963 B.n735 B.n734 10.6151
R964 B.n734 B.n733 10.6151
R965 B.n733 B.n46 10.6151
R966 B.n729 B.n46 10.6151
R967 B.n729 B.n728 10.6151
R968 B.n728 B.n727 10.6151
R969 B.n727 B.n48 10.6151
R970 B.n723 B.n48 10.6151
R971 B.n723 B.n722 10.6151
R972 B.n722 B.n721 10.6151
R973 B.n721 B.n50 10.6151
R974 B.n717 B.n50 10.6151
R975 B.n717 B.n716 10.6151
R976 B.n716 B.n715 10.6151
R977 B.n715 B.n52 10.6151
R978 B.n711 B.n710 10.6151
R979 B.n710 B.n709 10.6151
R980 B.n709 B.n57 10.6151
R981 B.n705 B.n57 10.6151
R982 B.n705 B.n704 10.6151
R983 B.n704 B.n703 10.6151
R984 B.n703 B.n59 10.6151
R985 B.n699 B.n59 10.6151
R986 B.n699 B.n698 10.6151
R987 B.n696 B.n63 10.6151
R988 B.n692 B.n63 10.6151
R989 B.n692 B.n691 10.6151
R990 B.n691 B.n690 10.6151
R991 B.n690 B.n65 10.6151
R992 B.n686 B.n65 10.6151
R993 B.n686 B.n685 10.6151
R994 B.n685 B.n684 10.6151
R995 B.n684 B.n67 10.6151
R996 B.n680 B.n67 10.6151
R997 B.n680 B.n679 10.6151
R998 B.n679 B.n678 10.6151
R999 B.n678 B.n69 10.6151
R1000 B.n674 B.n69 10.6151
R1001 B.n674 B.n673 10.6151
R1002 B.n673 B.n672 10.6151
R1003 B.n672 B.n71 10.6151
R1004 B.n668 B.n71 10.6151
R1005 B.n668 B.n667 10.6151
R1006 B.n667 B.n666 10.6151
R1007 B.n666 B.n73 10.6151
R1008 B.n662 B.n73 10.6151
R1009 B.n662 B.n661 10.6151
R1010 B.n661 B.n660 10.6151
R1011 B.n660 B.n75 10.6151
R1012 B.n656 B.n75 10.6151
R1013 B.n656 B.n655 10.6151
R1014 B.n655 B.n654 10.6151
R1015 B.n654 B.n77 10.6151
R1016 B.n650 B.n77 10.6151
R1017 B.n650 B.n649 10.6151
R1018 B.n649 B.n648 10.6151
R1019 B.n648 B.n79 10.6151
R1020 B.n644 B.n79 10.6151
R1021 B.n644 B.n643 10.6151
R1022 B.n643 B.n642 10.6151
R1023 B.n642 B.n81 10.6151
R1024 B.n638 B.n81 10.6151
R1025 B.n638 B.n637 10.6151
R1026 B.n637 B.n636 10.6151
R1027 B.n636 B.n83 10.6151
R1028 B.n632 B.n631 10.6151
R1029 B.n631 B.n630 10.6151
R1030 B.n630 B.n85 10.6151
R1031 B.n626 B.n85 10.6151
R1032 B.n626 B.n625 10.6151
R1033 B.n625 B.n624 10.6151
R1034 B.n624 B.n87 10.6151
R1035 B.n620 B.n87 10.6151
R1036 B.n620 B.n619 10.6151
R1037 B.n619 B.n618 10.6151
R1038 B.n618 B.n89 10.6151
R1039 B.n614 B.n89 10.6151
R1040 B.n614 B.n613 10.6151
R1041 B.n613 B.n612 10.6151
R1042 B.n612 B.n91 10.6151
R1043 B.n608 B.n91 10.6151
R1044 B.n608 B.n607 10.6151
R1045 B.n607 B.n606 10.6151
R1046 B.n606 B.n93 10.6151
R1047 B.n602 B.n93 10.6151
R1048 B.n602 B.n601 10.6151
R1049 B.n601 B.n600 10.6151
R1050 B.n600 B.n95 10.6151
R1051 B.n596 B.n95 10.6151
R1052 B.n596 B.n595 10.6151
R1053 B.n595 B.n594 10.6151
R1054 B.n594 B.n97 10.6151
R1055 B.n590 B.n97 10.6151
R1056 B.n590 B.n589 10.6151
R1057 B.n589 B.n588 10.6151
R1058 B.n588 B.n99 10.6151
R1059 B.n584 B.n99 10.6151
R1060 B.n584 B.n583 10.6151
R1061 B.n583 B.n582 10.6151
R1062 B.n582 B.n101 10.6151
R1063 B.n578 B.n101 10.6151
R1064 B.n578 B.n577 10.6151
R1065 B.n577 B.n576 10.6151
R1066 B.n576 B.n103 10.6151
R1067 B.n572 B.n103 10.6151
R1068 B.n572 B.n571 10.6151
R1069 B.n571 B.n570 10.6151
R1070 B.n570 B.n105 10.6151
R1071 B.n566 B.n105 10.6151
R1072 B.n566 B.n565 10.6151
R1073 B.n565 B.n564 10.6151
R1074 B.n564 B.n107 10.6151
R1075 B.n560 B.n107 10.6151
R1076 B.n560 B.n559 10.6151
R1077 B.n559 B.n558 10.6151
R1078 B.n558 B.n109 10.6151
R1079 B.n554 B.n109 10.6151
R1080 B.n554 B.n553 10.6151
R1081 B.n553 B.n552 10.6151
R1082 B.n552 B.n111 10.6151
R1083 B.n548 B.n111 10.6151
R1084 B.n548 B.n547 10.6151
R1085 B.n547 B.n546 10.6151
R1086 B.n546 B.n113 10.6151
R1087 B.n542 B.n113 10.6151
R1088 B.n542 B.n541 10.6151
R1089 B.n541 B.n540 10.6151
R1090 B.n540 B.n115 10.6151
R1091 B.n536 B.n115 10.6151
R1092 B.n536 B.n535 10.6151
R1093 B.n535 B.n534 10.6151
R1094 B.n534 B.n117 10.6151
R1095 B.n530 B.n117 10.6151
R1096 B.n530 B.n529 10.6151
R1097 B.n529 B.n528 10.6151
R1098 B.n528 B.n119 10.6151
R1099 B.n524 B.n119 10.6151
R1100 B.n524 B.n523 10.6151
R1101 B.n523 B.n522 10.6151
R1102 B.n522 B.n121 10.6151
R1103 B.n518 B.n121 10.6151
R1104 B.n518 B.n517 10.6151
R1105 B.n517 B.n516 10.6151
R1106 B.n516 B.n123 10.6151
R1107 B.n512 B.n123 10.6151
R1108 B.n512 B.n511 10.6151
R1109 B.n511 B.n510 10.6151
R1110 B.n510 B.n125 10.6151
R1111 B.n506 B.n125 10.6151
R1112 B.n506 B.n505 10.6151
R1113 B.n505 B.n504 10.6151
R1114 B.n504 B.n127 10.6151
R1115 B.n500 B.n127 10.6151
R1116 B.n500 B.n499 10.6151
R1117 B.n499 B.n498 10.6151
R1118 B.n498 B.n129 10.6151
R1119 B.n494 B.n129 10.6151
R1120 B.n494 B.n493 10.6151
R1121 B.n493 B.n492 10.6151
R1122 B.n492 B.n131 10.6151
R1123 B.n488 B.n131 10.6151
R1124 B.n488 B.n487 10.6151
R1125 B.n487 B.n486 10.6151
R1126 B.n486 B.n133 10.6151
R1127 B.n482 B.n133 10.6151
R1128 B.n482 B.n481 10.6151
R1129 B.n481 B.n480 10.6151
R1130 B.n480 B.n135 10.6151
R1131 B.n476 B.n135 10.6151
R1132 B.n476 B.n475 10.6151
R1133 B.n475 B.n474 10.6151
R1134 B.n474 B.n137 10.6151
R1135 B.n470 B.n137 10.6151
R1136 B.n470 B.n469 10.6151
R1137 B.n469 B.n468 10.6151
R1138 B.n468 B.n139 10.6151
R1139 B.n464 B.n139 10.6151
R1140 B.n464 B.n463 10.6151
R1141 B.n463 B.n462 10.6151
R1142 B.n462 B.n141 10.6151
R1143 B.n458 B.n141 10.6151
R1144 B.n458 B.n457 10.6151
R1145 B.n457 B.n456 10.6151
R1146 B.n456 B.n143 10.6151
R1147 B.n221 B.n1 10.6151
R1148 B.n224 B.n221 10.6151
R1149 B.n225 B.n224 10.6151
R1150 B.n226 B.n225 10.6151
R1151 B.n226 B.n219 10.6151
R1152 B.n230 B.n219 10.6151
R1153 B.n231 B.n230 10.6151
R1154 B.n232 B.n231 10.6151
R1155 B.n232 B.n217 10.6151
R1156 B.n236 B.n217 10.6151
R1157 B.n237 B.n236 10.6151
R1158 B.n238 B.n237 10.6151
R1159 B.n238 B.n215 10.6151
R1160 B.n242 B.n215 10.6151
R1161 B.n243 B.n242 10.6151
R1162 B.n244 B.n243 10.6151
R1163 B.n244 B.n213 10.6151
R1164 B.n248 B.n213 10.6151
R1165 B.n249 B.n248 10.6151
R1166 B.n250 B.n249 10.6151
R1167 B.n250 B.n211 10.6151
R1168 B.n254 B.n211 10.6151
R1169 B.n255 B.n254 10.6151
R1170 B.n256 B.n255 10.6151
R1171 B.n256 B.n209 10.6151
R1172 B.n260 B.n209 10.6151
R1173 B.n261 B.n260 10.6151
R1174 B.n262 B.n261 10.6151
R1175 B.n262 B.n207 10.6151
R1176 B.n266 B.n207 10.6151
R1177 B.n267 B.n266 10.6151
R1178 B.n268 B.n267 10.6151
R1179 B.n268 B.n205 10.6151
R1180 B.n272 B.n205 10.6151
R1181 B.n273 B.n272 10.6151
R1182 B.n274 B.n273 10.6151
R1183 B.n274 B.n203 10.6151
R1184 B.n278 B.n203 10.6151
R1185 B.n279 B.n278 10.6151
R1186 B.n280 B.n279 10.6151
R1187 B.n280 B.n201 10.6151
R1188 B.n284 B.n201 10.6151
R1189 B.n285 B.n284 10.6151
R1190 B.n286 B.n285 10.6151
R1191 B.n286 B.n199 10.6151
R1192 B.n290 B.n199 10.6151
R1193 B.n291 B.n290 10.6151
R1194 B.n292 B.n291 10.6151
R1195 B.n292 B.n197 10.6151
R1196 B.n296 B.n197 10.6151
R1197 B.n297 B.n296 10.6151
R1198 B.n298 B.n297 10.6151
R1199 B.n298 B.n195 10.6151
R1200 B.n302 B.n195 10.6151
R1201 B.n303 B.n302 10.6151
R1202 B.n304 B.n303 10.6151
R1203 B.n304 B.n193 10.6151
R1204 B.n308 B.n193 10.6151
R1205 B.n310 B.n309 10.6151
R1206 B.n310 B.n191 10.6151
R1207 B.n314 B.n191 10.6151
R1208 B.n315 B.n314 10.6151
R1209 B.n316 B.n315 10.6151
R1210 B.n316 B.n189 10.6151
R1211 B.n320 B.n189 10.6151
R1212 B.n321 B.n320 10.6151
R1213 B.n322 B.n321 10.6151
R1214 B.n322 B.n187 10.6151
R1215 B.n326 B.n187 10.6151
R1216 B.n327 B.n326 10.6151
R1217 B.n328 B.n327 10.6151
R1218 B.n328 B.n185 10.6151
R1219 B.n332 B.n185 10.6151
R1220 B.n333 B.n332 10.6151
R1221 B.n334 B.n333 10.6151
R1222 B.n334 B.n183 10.6151
R1223 B.n338 B.n183 10.6151
R1224 B.n339 B.n338 10.6151
R1225 B.n340 B.n339 10.6151
R1226 B.n340 B.n181 10.6151
R1227 B.n344 B.n181 10.6151
R1228 B.n345 B.n344 10.6151
R1229 B.n346 B.n345 10.6151
R1230 B.n346 B.n179 10.6151
R1231 B.n350 B.n179 10.6151
R1232 B.n351 B.n350 10.6151
R1233 B.n352 B.n351 10.6151
R1234 B.n352 B.n177 10.6151
R1235 B.n356 B.n177 10.6151
R1236 B.n357 B.n356 10.6151
R1237 B.n358 B.n357 10.6151
R1238 B.n358 B.n175 10.6151
R1239 B.n362 B.n175 10.6151
R1240 B.n363 B.n362 10.6151
R1241 B.n364 B.n363 10.6151
R1242 B.n364 B.n173 10.6151
R1243 B.n368 B.n173 10.6151
R1244 B.n369 B.n368 10.6151
R1245 B.n373 B.n369 10.6151
R1246 B.n377 B.n171 10.6151
R1247 B.n378 B.n377 10.6151
R1248 B.n379 B.n378 10.6151
R1249 B.n379 B.n169 10.6151
R1250 B.n383 B.n169 10.6151
R1251 B.n384 B.n383 10.6151
R1252 B.n385 B.n384 10.6151
R1253 B.n385 B.n167 10.6151
R1254 B.n389 B.n167 10.6151
R1255 B.n392 B.n391 10.6151
R1256 B.n392 B.n163 10.6151
R1257 B.n396 B.n163 10.6151
R1258 B.n397 B.n396 10.6151
R1259 B.n398 B.n397 10.6151
R1260 B.n398 B.n161 10.6151
R1261 B.n402 B.n161 10.6151
R1262 B.n403 B.n402 10.6151
R1263 B.n404 B.n403 10.6151
R1264 B.n404 B.n159 10.6151
R1265 B.n408 B.n159 10.6151
R1266 B.n409 B.n408 10.6151
R1267 B.n410 B.n409 10.6151
R1268 B.n410 B.n157 10.6151
R1269 B.n414 B.n157 10.6151
R1270 B.n415 B.n414 10.6151
R1271 B.n416 B.n415 10.6151
R1272 B.n416 B.n155 10.6151
R1273 B.n420 B.n155 10.6151
R1274 B.n421 B.n420 10.6151
R1275 B.n422 B.n421 10.6151
R1276 B.n422 B.n153 10.6151
R1277 B.n426 B.n153 10.6151
R1278 B.n427 B.n426 10.6151
R1279 B.n428 B.n427 10.6151
R1280 B.n428 B.n151 10.6151
R1281 B.n432 B.n151 10.6151
R1282 B.n433 B.n432 10.6151
R1283 B.n434 B.n433 10.6151
R1284 B.n434 B.n149 10.6151
R1285 B.n438 B.n149 10.6151
R1286 B.n439 B.n438 10.6151
R1287 B.n440 B.n439 10.6151
R1288 B.n440 B.n147 10.6151
R1289 B.n444 B.n147 10.6151
R1290 B.n445 B.n444 10.6151
R1291 B.n446 B.n445 10.6151
R1292 B.n446 B.n145 10.6151
R1293 B.n450 B.n145 10.6151
R1294 B.n451 B.n450 10.6151
R1295 B.n452 B.n451 10.6151
R1296 B.n56 B.n52 9.36635
R1297 B.n697 B.n696 9.36635
R1298 B.n373 B.n372 9.36635
R1299 B.n391 B.n390 9.36635
R1300 B.n865 B.n0 8.11757
R1301 B.n865 B.n1 8.11757
R1302 B.n711 B.n56 1.24928
R1303 B.n698 B.n697 1.24928
R1304 B.n372 B.n171 1.24928
R1305 B.n390 B.n389 1.24928
R1306 VP.n24 VP.n23 161.3
R1307 VP.n25 VP.n20 161.3
R1308 VP.n27 VP.n26 161.3
R1309 VP.n28 VP.n19 161.3
R1310 VP.n30 VP.n29 161.3
R1311 VP.n31 VP.n18 161.3
R1312 VP.n33 VP.n32 161.3
R1313 VP.n35 VP.n34 161.3
R1314 VP.n36 VP.n16 161.3
R1315 VP.n38 VP.n37 161.3
R1316 VP.n39 VP.n15 161.3
R1317 VP.n41 VP.n40 161.3
R1318 VP.n42 VP.n14 161.3
R1319 VP.n44 VP.n43 161.3
R1320 VP.n79 VP.n78 161.3
R1321 VP.n77 VP.n1 161.3
R1322 VP.n76 VP.n75 161.3
R1323 VP.n74 VP.n2 161.3
R1324 VP.n73 VP.n72 161.3
R1325 VP.n71 VP.n3 161.3
R1326 VP.n70 VP.n69 161.3
R1327 VP.n68 VP.n67 161.3
R1328 VP.n66 VP.n5 161.3
R1329 VP.n65 VP.n64 161.3
R1330 VP.n63 VP.n6 161.3
R1331 VP.n62 VP.n61 161.3
R1332 VP.n60 VP.n7 161.3
R1333 VP.n59 VP.n58 161.3
R1334 VP.n57 VP.n56 161.3
R1335 VP.n55 VP.n9 161.3
R1336 VP.n54 VP.n53 161.3
R1337 VP.n52 VP.n10 161.3
R1338 VP.n51 VP.n50 161.3
R1339 VP.n49 VP.n11 161.3
R1340 VP.n48 VP.n47 161.3
R1341 VP.n22 VP.t2 124.856
R1342 VP.n12 VP.t7 92.2191
R1343 VP.n8 VP.t4 92.2191
R1344 VP.n4 VP.t3 92.2191
R1345 VP.n0 VP.t0 92.2191
R1346 VP.n13 VP.t5 92.2191
R1347 VP.n17 VP.t6 92.2191
R1348 VP.n21 VP.t1 92.2191
R1349 VP.n46 VP.n12 77.8339
R1350 VP.n80 VP.n0 77.8339
R1351 VP.n45 VP.n13 77.8339
R1352 VP.n22 VP.n21 62.0322
R1353 VP.n46 VP.n45 53.7039
R1354 VP.n50 VP.n10 40.4934
R1355 VP.n54 VP.n10 40.4934
R1356 VP.n61 VP.n6 40.4934
R1357 VP.n65 VP.n6 40.4934
R1358 VP.n72 VP.n2 40.4934
R1359 VP.n76 VP.n2 40.4934
R1360 VP.n41 VP.n15 40.4934
R1361 VP.n37 VP.n15 40.4934
R1362 VP.n30 VP.n19 40.4934
R1363 VP.n26 VP.n19 40.4934
R1364 VP.n49 VP.n48 24.4675
R1365 VP.n50 VP.n49 24.4675
R1366 VP.n55 VP.n54 24.4675
R1367 VP.n56 VP.n55 24.4675
R1368 VP.n60 VP.n59 24.4675
R1369 VP.n61 VP.n60 24.4675
R1370 VP.n66 VP.n65 24.4675
R1371 VP.n67 VP.n66 24.4675
R1372 VP.n71 VP.n70 24.4675
R1373 VP.n72 VP.n71 24.4675
R1374 VP.n77 VP.n76 24.4675
R1375 VP.n78 VP.n77 24.4675
R1376 VP.n42 VP.n41 24.4675
R1377 VP.n43 VP.n42 24.4675
R1378 VP.n31 VP.n30 24.4675
R1379 VP.n32 VP.n31 24.4675
R1380 VP.n36 VP.n35 24.4675
R1381 VP.n37 VP.n36 24.4675
R1382 VP.n25 VP.n24 24.4675
R1383 VP.n26 VP.n25 24.4675
R1384 VP.n48 VP.n12 12.234
R1385 VP.n56 VP.n8 12.234
R1386 VP.n59 VP.n8 12.234
R1387 VP.n67 VP.n4 12.234
R1388 VP.n70 VP.n4 12.234
R1389 VP.n78 VP.n0 12.234
R1390 VP.n43 VP.n13 12.234
R1391 VP.n32 VP.n17 12.234
R1392 VP.n35 VP.n17 12.234
R1393 VP.n24 VP.n21 12.234
R1394 VP.n23 VP.n22 4.27755
R1395 VP.n45 VP.n44 0.354971
R1396 VP.n47 VP.n46 0.354971
R1397 VP.n80 VP.n79 0.354971
R1398 VP VP.n80 0.26696
R1399 VP.n23 VP.n20 0.189894
R1400 VP.n27 VP.n20 0.189894
R1401 VP.n28 VP.n27 0.189894
R1402 VP.n29 VP.n28 0.189894
R1403 VP.n29 VP.n18 0.189894
R1404 VP.n33 VP.n18 0.189894
R1405 VP.n34 VP.n33 0.189894
R1406 VP.n34 VP.n16 0.189894
R1407 VP.n38 VP.n16 0.189894
R1408 VP.n39 VP.n38 0.189894
R1409 VP.n40 VP.n39 0.189894
R1410 VP.n40 VP.n14 0.189894
R1411 VP.n44 VP.n14 0.189894
R1412 VP.n47 VP.n11 0.189894
R1413 VP.n51 VP.n11 0.189894
R1414 VP.n52 VP.n51 0.189894
R1415 VP.n53 VP.n52 0.189894
R1416 VP.n53 VP.n9 0.189894
R1417 VP.n57 VP.n9 0.189894
R1418 VP.n58 VP.n57 0.189894
R1419 VP.n58 VP.n7 0.189894
R1420 VP.n62 VP.n7 0.189894
R1421 VP.n63 VP.n62 0.189894
R1422 VP.n64 VP.n63 0.189894
R1423 VP.n64 VP.n5 0.189894
R1424 VP.n68 VP.n5 0.189894
R1425 VP.n69 VP.n68 0.189894
R1426 VP.n69 VP.n3 0.189894
R1427 VP.n73 VP.n3 0.189894
R1428 VP.n74 VP.n73 0.189894
R1429 VP.n75 VP.n74 0.189894
R1430 VP.n75 VP.n1 0.189894
R1431 VP.n79 VP.n1 0.189894
R1432 VTAIL.n530 VTAIL.n470 756.745
R1433 VTAIL.n62 VTAIL.n2 756.745
R1434 VTAIL.n128 VTAIL.n68 756.745
R1435 VTAIL.n196 VTAIL.n136 756.745
R1436 VTAIL.n464 VTAIL.n404 756.745
R1437 VTAIL.n396 VTAIL.n336 756.745
R1438 VTAIL.n330 VTAIL.n270 756.745
R1439 VTAIL.n262 VTAIL.n202 756.745
R1440 VTAIL.n490 VTAIL.n489 585
R1441 VTAIL.n495 VTAIL.n494 585
R1442 VTAIL.n497 VTAIL.n496 585
R1443 VTAIL.n486 VTAIL.n485 585
R1444 VTAIL.n503 VTAIL.n502 585
R1445 VTAIL.n505 VTAIL.n504 585
R1446 VTAIL.n482 VTAIL.n481 585
R1447 VTAIL.n512 VTAIL.n511 585
R1448 VTAIL.n513 VTAIL.n480 585
R1449 VTAIL.n515 VTAIL.n514 585
R1450 VTAIL.n478 VTAIL.n477 585
R1451 VTAIL.n521 VTAIL.n520 585
R1452 VTAIL.n523 VTAIL.n522 585
R1453 VTAIL.n474 VTAIL.n473 585
R1454 VTAIL.n529 VTAIL.n528 585
R1455 VTAIL.n531 VTAIL.n530 585
R1456 VTAIL.n22 VTAIL.n21 585
R1457 VTAIL.n27 VTAIL.n26 585
R1458 VTAIL.n29 VTAIL.n28 585
R1459 VTAIL.n18 VTAIL.n17 585
R1460 VTAIL.n35 VTAIL.n34 585
R1461 VTAIL.n37 VTAIL.n36 585
R1462 VTAIL.n14 VTAIL.n13 585
R1463 VTAIL.n44 VTAIL.n43 585
R1464 VTAIL.n45 VTAIL.n12 585
R1465 VTAIL.n47 VTAIL.n46 585
R1466 VTAIL.n10 VTAIL.n9 585
R1467 VTAIL.n53 VTAIL.n52 585
R1468 VTAIL.n55 VTAIL.n54 585
R1469 VTAIL.n6 VTAIL.n5 585
R1470 VTAIL.n61 VTAIL.n60 585
R1471 VTAIL.n63 VTAIL.n62 585
R1472 VTAIL.n88 VTAIL.n87 585
R1473 VTAIL.n93 VTAIL.n92 585
R1474 VTAIL.n95 VTAIL.n94 585
R1475 VTAIL.n84 VTAIL.n83 585
R1476 VTAIL.n101 VTAIL.n100 585
R1477 VTAIL.n103 VTAIL.n102 585
R1478 VTAIL.n80 VTAIL.n79 585
R1479 VTAIL.n110 VTAIL.n109 585
R1480 VTAIL.n111 VTAIL.n78 585
R1481 VTAIL.n113 VTAIL.n112 585
R1482 VTAIL.n76 VTAIL.n75 585
R1483 VTAIL.n119 VTAIL.n118 585
R1484 VTAIL.n121 VTAIL.n120 585
R1485 VTAIL.n72 VTAIL.n71 585
R1486 VTAIL.n127 VTAIL.n126 585
R1487 VTAIL.n129 VTAIL.n128 585
R1488 VTAIL.n156 VTAIL.n155 585
R1489 VTAIL.n161 VTAIL.n160 585
R1490 VTAIL.n163 VTAIL.n162 585
R1491 VTAIL.n152 VTAIL.n151 585
R1492 VTAIL.n169 VTAIL.n168 585
R1493 VTAIL.n171 VTAIL.n170 585
R1494 VTAIL.n148 VTAIL.n147 585
R1495 VTAIL.n178 VTAIL.n177 585
R1496 VTAIL.n179 VTAIL.n146 585
R1497 VTAIL.n181 VTAIL.n180 585
R1498 VTAIL.n144 VTAIL.n143 585
R1499 VTAIL.n187 VTAIL.n186 585
R1500 VTAIL.n189 VTAIL.n188 585
R1501 VTAIL.n140 VTAIL.n139 585
R1502 VTAIL.n195 VTAIL.n194 585
R1503 VTAIL.n197 VTAIL.n196 585
R1504 VTAIL.n465 VTAIL.n464 585
R1505 VTAIL.n463 VTAIL.n462 585
R1506 VTAIL.n408 VTAIL.n407 585
R1507 VTAIL.n457 VTAIL.n456 585
R1508 VTAIL.n455 VTAIL.n454 585
R1509 VTAIL.n412 VTAIL.n411 585
R1510 VTAIL.n449 VTAIL.n448 585
R1511 VTAIL.n447 VTAIL.n414 585
R1512 VTAIL.n446 VTAIL.n445 585
R1513 VTAIL.n417 VTAIL.n415 585
R1514 VTAIL.n440 VTAIL.n439 585
R1515 VTAIL.n438 VTAIL.n437 585
R1516 VTAIL.n421 VTAIL.n420 585
R1517 VTAIL.n432 VTAIL.n431 585
R1518 VTAIL.n430 VTAIL.n429 585
R1519 VTAIL.n425 VTAIL.n424 585
R1520 VTAIL.n397 VTAIL.n396 585
R1521 VTAIL.n395 VTAIL.n394 585
R1522 VTAIL.n340 VTAIL.n339 585
R1523 VTAIL.n389 VTAIL.n388 585
R1524 VTAIL.n387 VTAIL.n386 585
R1525 VTAIL.n344 VTAIL.n343 585
R1526 VTAIL.n381 VTAIL.n380 585
R1527 VTAIL.n379 VTAIL.n346 585
R1528 VTAIL.n378 VTAIL.n377 585
R1529 VTAIL.n349 VTAIL.n347 585
R1530 VTAIL.n372 VTAIL.n371 585
R1531 VTAIL.n370 VTAIL.n369 585
R1532 VTAIL.n353 VTAIL.n352 585
R1533 VTAIL.n364 VTAIL.n363 585
R1534 VTAIL.n362 VTAIL.n361 585
R1535 VTAIL.n357 VTAIL.n356 585
R1536 VTAIL.n331 VTAIL.n330 585
R1537 VTAIL.n329 VTAIL.n328 585
R1538 VTAIL.n274 VTAIL.n273 585
R1539 VTAIL.n323 VTAIL.n322 585
R1540 VTAIL.n321 VTAIL.n320 585
R1541 VTAIL.n278 VTAIL.n277 585
R1542 VTAIL.n315 VTAIL.n314 585
R1543 VTAIL.n313 VTAIL.n280 585
R1544 VTAIL.n312 VTAIL.n311 585
R1545 VTAIL.n283 VTAIL.n281 585
R1546 VTAIL.n306 VTAIL.n305 585
R1547 VTAIL.n304 VTAIL.n303 585
R1548 VTAIL.n287 VTAIL.n286 585
R1549 VTAIL.n298 VTAIL.n297 585
R1550 VTAIL.n296 VTAIL.n295 585
R1551 VTAIL.n291 VTAIL.n290 585
R1552 VTAIL.n263 VTAIL.n262 585
R1553 VTAIL.n261 VTAIL.n260 585
R1554 VTAIL.n206 VTAIL.n205 585
R1555 VTAIL.n255 VTAIL.n254 585
R1556 VTAIL.n253 VTAIL.n252 585
R1557 VTAIL.n210 VTAIL.n209 585
R1558 VTAIL.n247 VTAIL.n246 585
R1559 VTAIL.n245 VTAIL.n212 585
R1560 VTAIL.n244 VTAIL.n243 585
R1561 VTAIL.n215 VTAIL.n213 585
R1562 VTAIL.n238 VTAIL.n237 585
R1563 VTAIL.n236 VTAIL.n235 585
R1564 VTAIL.n219 VTAIL.n218 585
R1565 VTAIL.n230 VTAIL.n229 585
R1566 VTAIL.n228 VTAIL.n227 585
R1567 VTAIL.n223 VTAIL.n222 585
R1568 VTAIL.n491 VTAIL.t2 329.036
R1569 VTAIL.n23 VTAIL.t1 329.036
R1570 VTAIL.n89 VTAIL.t9 329.036
R1571 VTAIL.n157 VTAIL.t10 329.036
R1572 VTAIL.n426 VTAIL.t14 329.036
R1573 VTAIL.n358 VTAIL.t11 329.036
R1574 VTAIL.n292 VTAIL.t3 329.036
R1575 VTAIL.n224 VTAIL.t7 329.036
R1576 VTAIL.n495 VTAIL.n489 171.744
R1577 VTAIL.n496 VTAIL.n495 171.744
R1578 VTAIL.n496 VTAIL.n485 171.744
R1579 VTAIL.n503 VTAIL.n485 171.744
R1580 VTAIL.n504 VTAIL.n503 171.744
R1581 VTAIL.n504 VTAIL.n481 171.744
R1582 VTAIL.n512 VTAIL.n481 171.744
R1583 VTAIL.n513 VTAIL.n512 171.744
R1584 VTAIL.n514 VTAIL.n513 171.744
R1585 VTAIL.n514 VTAIL.n477 171.744
R1586 VTAIL.n521 VTAIL.n477 171.744
R1587 VTAIL.n522 VTAIL.n521 171.744
R1588 VTAIL.n522 VTAIL.n473 171.744
R1589 VTAIL.n529 VTAIL.n473 171.744
R1590 VTAIL.n530 VTAIL.n529 171.744
R1591 VTAIL.n27 VTAIL.n21 171.744
R1592 VTAIL.n28 VTAIL.n27 171.744
R1593 VTAIL.n28 VTAIL.n17 171.744
R1594 VTAIL.n35 VTAIL.n17 171.744
R1595 VTAIL.n36 VTAIL.n35 171.744
R1596 VTAIL.n36 VTAIL.n13 171.744
R1597 VTAIL.n44 VTAIL.n13 171.744
R1598 VTAIL.n45 VTAIL.n44 171.744
R1599 VTAIL.n46 VTAIL.n45 171.744
R1600 VTAIL.n46 VTAIL.n9 171.744
R1601 VTAIL.n53 VTAIL.n9 171.744
R1602 VTAIL.n54 VTAIL.n53 171.744
R1603 VTAIL.n54 VTAIL.n5 171.744
R1604 VTAIL.n61 VTAIL.n5 171.744
R1605 VTAIL.n62 VTAIL.n61 171.744
R1606 VTAIL.n93 VTAIL.n87 171.744
R1607 VTAIL.n94 VTAIL.n93 171.744
R1608 VTAIL.n94 VTAIL.n83 171.744
R1609 VTAIL.n101 VTAIL.n83 171.744
R1610 VTAIL.n102 VTAIL.n101 171.744
R1611 VTAIL.n102 VTAIL.n79 171.744
R1612 VTAIL.n110 VTAIL.n79 171.744
R1613 VTAIL.n111 VTAIL.n110 171.744
R1614 VTAIL.n112 VTAIL.n111 171.744
R1615 VTAIL.n112 VTAIL.n75 171.744
R1616 VTAIL.n119 VTAIL.n75 171.744
R1617 VTAIL.n120 VTAIL.n119 171.744
R1618 VTAIL.n120 VTAIL.n71 171.744
R1619 VTAIL.n127 VTAIL.n71 171.744
R1620 VTAIL.n128 VTAIL.n127 171.744
R1621 VTAIL.n161 VTAIL.n155 171.744
R1622 VTAIL.n162 VTAIL.n161 171.744
R1623 VTAIL.n162 VTAIL.n151 171.744
R1624 VTAIL.n169 VTAIL.n151 171.744
R1625 VTAIL.n170 VTAIL.n169 171.744
R1626 VTAIL.n170 VTAIL.n147 171.744
R1627 VTAIL.n178 VTAIL.n147 171.744
R1628 VTAIL.n179 VTAIL.n178 171.744
R1629 VTAIL.n180 VTAIL.n179 171.744
R1630 VTAIL.n180 VTAIL.n143 171.744
R1631 VTAIL.n187 VTAIL.n143 171.744
R1632 VTAIL.n188 VTAIL.n187 171.744
R1633 VTAIL.n188 VTAIL.n139 171.744
R1634 VTAIL.n195 VTAIL.n139 171.744
R1635 VTAIL.n196 VTAIL.n195 171.744
R1636 VTAIL.n464 VTAIL.n463 171.744
R1637 VTAIL.n463 VTAIL.n407 171.744
R1638 VTAIL.n456 VTAIL.n407 171.744
R1639 VTAIL.n456 VTAIL.n455 171.744
R1640 VTAIL.n455 VTAIL.n411 171.744
R1641 VTAIL.n448 VTAIL.n411 171.744
R1642 VTAIL.n448 VTAIL.n447 171.744
R1643 VTAIL.n447 VTAIL.n446 171.744
R1644 VTAIL.n446 VTAIL.n415 171.744
R1645 VTAIL.n439 VTAIL.n415 171.744
R1646 VTAIL.n439 VTAIL.n438 171.744
R1647 VTAIL.n438 VTAIL.n420 171.744
R1648 VTAIL.n431 VTAIL.n420 171.744
R1649 VTAIL.n431 VTAIL.n430 171.744
R1650 VTAIL.n430 VTAIL.n424 171.744
R1651 VTAIL.n396 VTAIL.n395 171.744
R1652 VTAIL.n395 VTAIL.n339 171.744
R1653 VTAIL.n388 VTAIL.n339 171.744
R1654 VTAIL.n388 VTAIL.n387 171.744
R1655 VTAIL.n387 VTAIL.n343 171.744
R1656 VTAIL.n380 VTAIL.n343 171.744
R1657 VTAIL.n380 VTAIL.n379 171.744
R1658 VTAIL.n379 VTAIL.n378 171.744
R1659 VTAIL.n378 VTAIL.n347 171.744
R1660 VTAIL.n371 VTAIL.n347 171.744
R1661 VTAIL.n371 VTAIL.n370 171.744
R1662 VTAIL.n370 VTAIL.n352 171.744
R1663 VTAIL.n363 VTAIL.n352 171.744
R1664 VTAIL.n363 VTAIL.n362 171.744
R1665 VTAIL.n362 VTAIL.n356 171.744
R1666 VTAIL.n330 VTAIL.n329 171.744
R1667 VTAIL.n329 VTAIL.n273 171.744
R1668 VTAIL.n322 VTAIL.n273 171.744
R1669 VTAIL.n322 VTAIL.n321 171.744
R1670 VTAIL.n321 VTAIL.n277 171.744
R1671 VTAIL.n314 VTAIL.n277 171.744
R1672 VTAIL.n314 VTAIL.n313 171.744
R1673 VTAIL.n313 VTAIL.n312 171.744
R1674 VTAIL.n312 VTAIL.n281 171.744
R1675 VTAIL.n305 VTAIL.n281 171.744
R1676 VTAIL.n305 VTAIL.n304 171.744
R1677 VTAIL.n304 VTAIL.n286 171.744
R1678 VTAIL.n297 VTAIL.n286 171.744
R1679 VTAIL.n297 VTAIL.n296 171.744
R1680 VTAIL.n296 VTAIL.n290 171.744
R1681 VTAIL.n262 VTAIL.n261 171.744
R1682 VTAIL.n261 VTAIL.n205 171.744
R1683 VTAIL.n254 VTAIL.n205 171.744
R1684 VTAIL.n254 VTAIL.n253 171.744
R1685 VTAIL.n253 VTAIL.n209 171.744
R1686 VTAIL.n246 VTAIL.n209 171.744
R1687 VTAIL.n246 VTAIL.n245 171.744
R1688 VTAIL.n245 VTAIL.n244 171.744
R1689 VTAIL.n244 VTAIL.n213 171.744
R1690 VTAIL.n237 VTAIL.n213 171.744
R1691 VTAIL.n237 VTAIL.n236 171.744
R1692 VTAIL.n236 VTAIL.n218 171.744
R1693 VTAIL.n229 VTAIL.n218 171.744
R1694 VTAIL.n229 VTAIL.n228 171.744
R1695 VTAIL.n228 VTAIL.n222 171.744
R1696 VTAIL.t2 VTAIL.n489 85.8723
R1697 VTAIL.t1 VTAIL.n21 85.8723
R1698 VTAIL.t9 VTAIL.n87 85.8723
R1699 VTAIL.t10 VTAIL.n155 85.8723
R1700 VTAIL.t14 VTAIL.n424 85.8723
R1701 VTAIL.t11 VTAIL.n356 85.8723
R1702 VTAIL.t3 VTAIL.n290 85.8723
R1703 VTAIL.t7 VTAIL.n222 85.8723
R1704 VTAIL.n403 VTAIL.n402 57.3544
R1705 VTAIL.n269 VTAIL.n268 57.3544
R1706 VTAIL.n1 VTAIL.n0 57.3542
R1707 VTAIL.n135 VTAIL.n134 57.3542
R1708 VTAIL.n535 VTAIL.n534 32.3793
R1709 VTAIL.n67 VTAIL.n66 32.3793
R1710 VTAIL.n133 VTAIL.n132 32.3793
R1711 VTAIL.n201 VTAIL.n200 32.3793
R1712 VTAIL.n469 VTAIL.n468 32.3793
R1713 VTAIL.n401 VTAIL.n400 32.3793
R1714 VTAIL.n335 VTAIL.n334 32.3793
R1715 VTAIL.n267 VTAIL.n266 32.3793
R1716 VTAIL.n535 VTAIL.n469 25.841
R1717 VTAIL.n267 VTAIL.n201 25.841
R1718 VTAIL.n515 VTAIL.n480 13.1884
R1719 VTAIL.n47 VTAIL.n12 13.1884
R1720 VTAIL.n113 VTAIL.n78 13.1884
R1721 VTAIL.n181 VTAIL.n146 13.1884
R1722 VTAIL.n449 VTAIL.n414 13.1884
R1723 VTAIL.n381 VTAIL.n346 13.1884
R1724 VTAIL.n315 VTAIL.n280 13.1884
R1725 VTAIL.n247 VTAIL.n212 13.1884
R1726 VTAIL.n511 VTAIL.n510 12.8005
R1727 VTAIL.n516 VTAIL.n478 12.8005
R1728 VTAIL.n43 VTAIL.n42 12.8005
R1729 VTAIL.n48 VTAIL.n10 12.8005
R1730 VTAIL.n109 VTAIL.n108 12.8005
R1731 VTAIL.n114 VTAIL.n76 12.8005
R1732 VTAIL.n177 VTAIL.n176 12.8005
R1733 VTAIL.n182 VTAIL.n144 12.8005
R1734 VTAIL.n450 VTAIL.n412 12.8005
R1735 VTAIL.n445 VTAIL.n416 12.8005
R1736 VTAIL.n382 VTAIL.n344 12.8005
R1737 VTAIL.n377 VTAIL.n348 12.8005
R1738 VTAIL.n316 VTAIL.n278 12.8005
R1739 VTAIL.n311 VTAIL.n282 12.8005
R1740 VTAIL.n248 VTAIL.n210 12.8005
R1741 VTAIL.n243 VTAIL.n214 12.8005
R1742 VTAIL.n509 VTAIL.n482 12.0247
R1743 VTAIL.n520 VTAIL.n519 12.0247
R1744 VTAIL.n41 VTAIL.n14 12.0247
R1745 VTAIL.n52 VTAIL.n51 12.0247
R1746 VTAIL.n107 VTAIL.n80 12.0247
R1747 VTAIL.n118 VTAIL.n117 12.0247
R1748 VTAIL.n175 VTAIL.n148 12.0247
R1749 VTAIL.n186 VTAIL.n185 12.0247
R1750 VTAIL.n454 VTAIL.n453 12.0247
R1751 VTAIL.n444 VTAIL.n417 12.0247
R1752 VTAIL.n386 VTAIL.n385 12.0247
R1753 VTAIL.n376 VTAIL.n349 12.0247
R1754 VTAIL.n320 VTAIL.n319 12.0247
R1755 VTAIL.n310 VTAIL.n283 12.0247
R1756 VTAIL.n252 VTAIL.n251 12.0247
R1757 VTAIL.n242 VTAIL.n215 12.0247
R1758 VTAIL.n506 VTAIL.n505 11.249
R1759 VTAIL.n523 VTAIL.n476 11.249
R1760 VTAIL.n38 VTAIL.n37 11.249
R1761 VTAIL.n55 VTAIL.n8 11.249
R1762 VTAIL.n104 VTAIL.n103 11.249
R1763 VTAIL.n121 VTAIL.n74 11.249
R1764 VTAIL.n172 VTAIL.n171 11.249
R1765 VTAIL.n189 VTAIL.n142 11.249
R1766 VTAIL.n457 VTAIL.n410 11.249
R1767 VTAIL.n441 VTAIL.n440 11.249
R1768 VTAIL.n389 VTAIL.n342 11.249
R1769 VTAIL.n373 VTAIL.n372 11.249
R1770 VTAIL.n323 VTAIL.n276 11.249
R1771 VTAIL.n307 VTAIL.n306 11.249
R1772 VTAIL.n255 VTAIL.n208 11.249
R1773 VTAIL.n239 VTAIL.n238 11.249
R1774 VTAIL.n491 VTAIL.n490 10.7239
R1775 VTAIL.n23 VTAIL.n22 10.7239
R1776 VTAIL.n89 VTAIL.n88 10.7239
R1777 VTAIL.n157 VTAIL.n156 10.7239
R1778 VTAIL.n426 VTAIL.n425 10.7239
R1779 VTAIL.n358 VTAIL.n357 10.7239
R1780 VTAIL.n292 VTAIL.n291 10.7239
R1781 VTAIL.n224 VTAIL.n223 10.7239
R1782 VTAIL.n502 VTAIL.n484 10.4732
R1783 VTAIL.n524 VTAIL.n474 10.4732
R1784 VTAIL.n34 VTAIL.n16 10.4732
R1785 VTAIL.n56 VTAIL.n6 10.4732
R1786 VTAIL.n100 VTAIL.n82 10.4732
R1787 VTAIL.n122 VTAIL.n72 10.4732
R1788 VTAIL.n168 VTAIL.n150 10.4732
R1789 VTAIL.n190 VTAIL.n140 10.4732
R1790 VTAIL.n458 VTAIL.n408 10.4732
R1791 VTAIL.n437 VTAIL.n419 10.4732
R1792 VTAIL.n390 VTAIL.n340 10.4732
R1793 VTAIL.n369 VTAIL.n351 10.4732
R1794 VTAIL.n324 VTAIL.n274 10.4732
R1795 VTAIL.n303 VTAIL.n285 10.4732
R1796 VTAIL.n256 VTAIL.n206 10.4732
R1797 VTAIL.n235 VTAIL.n217 10.4732
R1798 VTAIL.n501 VTAIL.n486 9.69747
R1799 VTAIL.n528 VTAIL.n527 9.69747
R1800 VTAIL.n33 VTAIL.n18 9.69747
R1801 VTAIL.n60 VTAIL.n59 9.69747
R1802 VTAIL.n99 VTAIL.n84 9.69747
R1803 VTAIL.n126 VTAIL.n125 9.69747
R1804 VTAIL.n167 VTAIL.n152 9.69747
R1805 VTAIL.n194 VTAIL.n193 9.69747
R1806 VTAIL.n462 VTAIL.n461 9.69747
R1807 VTAIL.n436 VTAIL.n421 9.69747
R1808 VTAIL.n394 VTAIL.n393 9.69747
R1809 VTAIL.n368 VTAIL.n353 9.69747
R1810 VTAIL.n328 VTAIL.n327 9.69747
R1811 VTAIL.n302 VTAIL.n287 9.69747
R1812 VTAIL.n260 VTAIL.n259 9.69747
R1813 VTAIL.n234 VTAIL.n219 9.69747
R1814 VTAIL.n534 VTAIL.n533 9.45567
R1815 VTAIL.n66 VTAIL.n65 9.45567
R1816 VTAIL.n132 VTAIL.n131 9.45567
R1817 VTAIL.n200 VTAIL.n199 9.45567
R1818 VTAIL.n468 VTAIL.n467 9.45567
R1819 VTAIL.n400 VTAIL.n399 9.45567
R1820 VTAIL.n334 VTAIL.n333 9.45567
R1821 VTAIL.n266 VTAIL.n265 9.45567
R1822 VTAIL.n533 VTAIL.n532 9.3005
R1823 VTAIL.n472 VTAIL.n471 9.3005
R1824 VTAIL.n527 VTAIL.n526 9.3005
R1825 VTAIL.n525 VTAIL.n524 9.3005
R1826 VTAIL.n476 VTAIL.n475 9.3005
R1827 VTAIL.n519 VTAIL.n518 9.3005
R1828 VTAIL.n517 VTAIL.n516 9.3005
R1829 VTAIL.n493 VTAIL.n492 9.3005
R1830 VTAIL.n488 VTAIL.n487 9.3005
R1831 VTAIL.n499 VTAIL.n498 9.3005
R1832 VTAIL.n501 VTAIL.n500 9.3005
R1833 VTAIL.n484 VTAIL.n483 9.3005
R1834 VTAIL.n507 VTAIL.n506 9.3005
R1835 VTAIL.n509 VTAIL.n508 9.3005
R1836 VTAIL.n510 VTAIL.n479 9.3005
R1837 VTAIL.n65 VTAIL.n64 9.3005
R1838 VTAIL.n4 VTAIL.n3 9.3005
R1839 VTAIL.n59 VTAIL.n58 9.3005
R1840 VTAIL.n57 VTAIL.n56 9.3005
R1841 VTAIL.n8 VTAIL.n7 9.3005
R1842 VTAIL.n51 VTAIL.n50 9.3005
R1843 VTAIL.n49 VTAIL.n48 9.3005
R1844 VTAIL.n25 VTAIL.n24 9.3005
R1845 VTAIL.n20 VTAIL.n19 9.3005
R1846 VTAIL.n31 VTAIL.n30 9.3005
R1847 VTAIL.n33 VTAIL.n32 9.3005
R1848 VTAIL.n16 VTAIL.n15 9.3005
R1849 VTAIL.n39 VTAIL.n38 9.3005
R1850 VTAIL.n41 VTAIL.n40 9.3005
R1851 VTAIL.n42 VTAIL.n11 9.3005
R1852 VTAIL.n131 VTAIL.n130 9.3005
R1853 VTAIL.n70 VTAIL.n69 9.3005
R1854 VTAIL.n125 VTAIL.n124 9.3005
R1855 VTAIL.n123 VTAIL.n122 9.3005
R1856 VTAIL.n74 VTAIL.n73 9.3005
R1857 VTAIL.n117 VTAIL.n116 9.3005
R1858 VTAIL.n115 VTAIL.n114 9.3005
R1859 VTAIL.n91 VTAIL.n90 9.3005
R1860 VTAIL.n86 VTAIL.n85 9.3005
R1861 VTAIL.n97 VTAIL.n96 9.3005
R1862 VTAIL.n99 VTAIL.n98 9.3005
R1863 VTAIL.n82 VTAIL.n81 9.3005
R1864 VTAIL.n105 VTAIL.n104 9.3005
R1865 VTAIL.n107 VTAIL.n106 9.3005
R1866 VTAIL.n108 VTAIL.n77 9.3005
R1867 VTAIL.n199 VTAIL.n198 9.3005
R1868 VTAIL.n138 VTAIL.n137 9.3005
R1869 VTAIL.n193 VTAIL.n192 9.3005
R1870 VTAIL.n191 VTAIL.n190 9.3005
R1871 VTAIL.n142 VTAIL.n141 9.3005
R1872 VTAIL.n185 VTAIL.n184 9.3005
R1873 VTAIL.n183 VTAIL.n182 9.3005
R1874 VTAIL.n159 VTAIL.n158 9.3005
R1875 VTAIL.n154 VTAIL.n153 9.3005
R1876 VTAIL.n165 VTAIL.n164 9.3005
R1877 VTAIL.n167 VTAIL.n166 9.3005
R1878 VTAIL.n150 VTAIL.n149 9.3005
R1879 VTAIL.n173 VTAIL.n172 9.3005
R1880 VTAIL.n175 VTAIL.n174 9.3005
R1881 VTAIL.n176 VTAIL.n145 9.3005
R1882 VTAIL.n428 VTAIL.n427 9.3005
R1883 VTAIL.n423 VTAIL.n422 9.3005
R1884 VTAIL.n434 VTAIL.n433 9.3005
R1885 VTAIL.n436 VTAIL.n435 9.3005
R1886 VTAIL.n419 VTAIL.n418 9.3005
R1887 VTAIL.n442 VTAIL.n441 9.3005
R1888 VTAIL.n444 VTAIL.n443 9.3005
R1889 VTAIL.n416 VTAIL.n413 9.3005
R1890 VTAIL.n467 VTAIL.n466 9.3005
R1891 VTAIL.n406 VTAIL.n405 9.3005
R1892 VTAIL.n461 VTAIL.n460 9.3005
R1893 VTAIL.n459 VTAIL.n458 9.3005
R1894 VTAIL.n410 VTAIL.n409 9.3005
R1895 VTAIL.n453 VTAIL.n452 9.3005
R1896 VTAIL.n451 VTAIL.n450 9.3005
R1897 VTAIL.n360 VTAIL.n359 9.3005
R1898 VTAIL.n355 VTAIL.n354 9.3005
R1899 VTAIL.n366 VTAIL.n365 9.3005
R1900 VTAIL.n368 VTAIL.n367 9.3005
R1901 VTAIL.n351 VTAIL.n350 9.3005
R1902 VTAIL.n374 VTAIL.n373 9.3005
R1903 VTAIL.n376 VTAIL.n375 9.3005
R1904 VTAIL.n348 VTAIL.n345 9.3005
R1905 VTAIL.n399 VTAIL.n398 9.3005
R1906 VTAIL.n338 VTAIL.n337 9.3005
R1907 VTAIL.n393 VTAIL.n392 9.3005
R1908 VTAIL.n391 VTAIL.n390 9.3005
R1909 VTAIL.n342 VTAIL.n341 9.3005
R1910 VTAIL.n385 VTAIL.n384 9.3005
R1911 VTAIL.n383 VTAIL.n382 9.3005
R1912 VTAIL.n294 VTAIL.n293 9.3005
R1913 VTAIL.n289 VTAIL.n288 9.3005
R1914 VTAIL.n300 VTAIL.n299 9.3005
R1915 VTAIL.n302 VTAIL.n301 9.3005
R1916 VTAIL.n285 VTAIL.n284 9.3005
R1917 VTAIL.n308 VTAIL.n307 9.3005
R1918 VTAIL.n310 VTAIL.n309 9.3005
R1919 VTAIL.n282 VTAIL.n279 9.3005
R1920 VTAIL.n333 VTAIL.n332 9.3005
R1921 VTAIL.n272 VTAIL.n271 9.3005
R1922 VTAIL.n327 VTAIL.n326 9.3005
R1923 VTAIL.n325 VTAIL.n324 9.3005
R1924 VTAIL.n276 VTAIL.n275 9.3005
R1925 VTAIL.n319 VTAIL.n318 9.3005
R1926 VTAIL.n317 VTAIL.n316 9.3005
R1927 VTAIL.n226 VTAIL.n225 9.3005
R1928 VTAIL.n221 VTAIL.n220 9.3005
R1929 VTAIL.n232 VTAIL.n231 9.3005
R1930 VTAIL.n234 VTAIL.n233 9.3005
R1931 VTAIL.n217 VTAIL.n216 9.3005
R1932 VTAIL.n240 VTAIL.n239 9.3005
R1933 VTAIL.n242 VTAIL.n241 9.3005
R1934 VTAIL.n214 VTAIL.n211 9.3005
R1935 VTAIL.n265 VTAIL.n264 9.3005
R1936 VTAIL.n204 VTAIL.n203 9.3005
R1937 VTAIL.n259 VTAIL.n258 9.3005
R1938 VTAIL.n257 VTAIL.n256 9.3005
R1939 VTAIL.n208 VTAIL.n207 9.3005
R1940 VTAIL.n251 VTAIL.n250 9.3005
R1941 VTAIL.n249 VTAIL.n248 9.3005
R1942 VTAIL.n498 VTAIL.n497 8.92171
R1943 VTAIL.n531 VTAIL.n472 8.92171
R1944 VTAIL.n30 VTAIL.n29 8.92171
R1945 VTAIL.n63 VTAIL.n4 8.92171
R1946 VTAIL.n96 VTAIL.n95 8.92171
R1947 VTAIL.n129 VTAIL.n70 8.92171
R1948 VTAIL.n164 VTAIL.n163 8.92171
R1949 VTAIL.n197 VTAIL.n138 8.92171
R1950 VTAIL.n465 VTAIL.n406 8.92171
R1951 VTAIL.n433 VTAIL.n432 8.92171
R1952 VTAIL.n397 VTAIL.n338 8.92171
R1953 VTAIL.n365 VTAIL.n364 8.92171
R1954 VTAIL.n331 VTAIL.n272 8.92171
R1955 VTAIL.n299 VTAIL.n298 8.92171
R1956 VTAIL.n263 VTAIL.n204 8.92171
R1957 VTAIL.n231 VTAIL.n230 8.92171
R1958 VTAIL.n494 VTAIL.n488 8.14595
R1959 VTAIL.n532 VTAIL.n470 8.14595
R1960 VTAIL.n26 VTAIL.n20 8.14595
R1961 VTAIL.n64 VTAIL.n2 8.14595
R1962 VTAIL.n92 VTAIL.n86 8.14595
R1963 VTAIL.n130 VTAIL.n68 8.14595
R1964 VTAIL.n160 VTAIL.n154 8.14595
R1965 VTAIL.n198 VTAIL.n136 8.14595
R1966 VTAIL.n466 VTAIL.n404 8.14595
R1967 VTAIL.n429 VTAIL.n423 8.14595
R1968 VTAIL.n398 VTAIL.n336 8.14595
R1969 VTAIL.n361 VTAIL.n355 8.14595
R1970 VTAIL.n332 VTAIL.n270 8.14595
R1971 VTAIL.n295 VTAIL.n289 8.14595
R1972 VTAIL.n264 VTAIL.n202 8.14595
R1973 VTAIL.n227 VTAIL.n221 8.14595
R1974 VTAIL.n493 VTAIL.n490 7.3702
R1975 VTAIL.n25 VTAIL.n22 7.3702
R1976 VTAIL.n91 VTAIL.n88 7.3702
R1977 VTAIL.n159 VTAIL.n156 7.3702
R1978 VTAIL.n428 VTAIL.n425 7.3702
R1979 VTAIL.n360 VTAIL.n357 7.3702
R1980 VTAIL.n294 VTAIL.n291 7.3702
R1981 VTAIL.n226 VTAIL.n223 7.3702
R1982 VTAIL.n494 VTAIL.n493 5.81868
R1983 VTAIL.n534 VTAIL.n470 5.81868
R1984 VTAIL.n26 VTAIL.n25 5.81868
R1985 VTAIL.n66 VTAIL.n2 5.81868
R1986 VTAIL.n92 VTAIL.n91 5.81868
R1987 VTAIL.n132 VTAIL.n68 5.81868
R1988 VTAIL.n160 VTAIL.n159 5.81868
R1989 VTAIL.n200 VTAIL.n136 5.81868
R1990 VTAIL.n468 VTAIL.n404 5.81868
R1991 VTAIL.n429 VTAIL.n428 5.81868
R1992 VTAIL.n400 VTAIL.n336 5.81868
R1993 VTAIL.n361 VTAIL.n360 5.81868
R1994 VTAIL.n334 VTAIL.n270 5.81868
R1995 VTAIL.n295 VTAIL.n294 5.81868
R1996 VTAIL.n266 VTAIL.n202 5.81868
R1997 VTAIL.n227 VTAIL.n226 5.81868
R1998 VTAIL.n497 VTAIL.n488 5.04292
R1999 VTAIL.n532 VTAIL.n531 5.04292
R2000 VTAIL.n29 VTAIL.n20 5.04292
R2001 VTAIL.n64 VTAIL.n63 5.04292
R2002 VTAIL.n95 VTAIL.n86 5.04292
R2003 VTAIL.n130 VTAIL.n129 5.04292
R2004 VTAIL.n163 VTAIL.n154 5.04292
R2005 VTAIL.n198 VTAIL.n197 5.04292
R2006 VTAIL.n466 VTAIL.n465 5.04292
R2007 VTAIL.n432 VTAIL.n423 5.04292
R2008 VTAIL.n398 VTAIL.n397 5.04292
R2009 VTAIL.n364 VTAIL.n355 5.04292
R2010 VTAIL.n332 VTAIL.n331 5.04292
R2011 VTAIL.n298 VTAIL.n289 5.04292
R2012 VTAIL.n264 VTAIL.n263 5.04292
R2013 VTAIL.n230 VTAIL.n221 5.04292
R2014 VTAIL.n498 VTAIL.n486 4.26717
R2015 VTAIL.n528 VTAIL.n472 4.26717
R2016 VTAIL.n30 VTAIL.n18 4.26717
R2017 VTAIL.n60 VTAIL.n4 4.26717
R2018 VTAIL.n96 VTAIL.n84 4.26717
R2019 VTAIL.n126 VTAIL.n70 4.26717
R2020 VTAIL.n164 VTAIL.n152 4.26717
R2021 VTAIL.n194 VTAIL.n138 4.26717
R2022 VTAIL.n462 VTAIL.n406 4.26717
R2023 VTAIL.n433 VTAIL.n421 4.26717
R2024 VTAIL.n394 VTAIL.n338 4.26717
R2025 VTAIL.n365 VTAIL.n353 4.26717
R2026 VTAIL.n328 VTAIL.n272 4.26717
R2027 VTAIL.n299 VTAIL.n287 4.26717
R2028 VTAIL.n260 VTAIL.n204 4.26717
R2029 VTAIL.n231 VTAIL.n219 4.26717
R2030 VTAIL.n502 VTAIL.n501 3.49141
R2031 VTAIL.n527 VTAIL.n474 3.49141
R2032 VTAIL.n34 VTAIL.n33 3.49141
R2033 VTAIL.n59 VTAIL.n6 3.49141
R2034 VTAIL.n100 VTAIL.n99 3.49141
R2035 VTAIL.n125 VTAIL.n72 3.49141
R2036 VTAIL.n168 VTAIL.n167 3.49141
R2037 VTAIL.n193 VTAIL.n140 3.49141
R2038 VTAIL.n461 VTAIL.n408 3.49141
R2039 VTAIL.n437 VTAIL.n436 3.49141
R2040 VTAIL.n393 VTAIL.n340 3.49141
R2041 VTAIL.n369 VTAIL.n368 3.49141
R2042 VTAIL.n327 VTAIL.n274 3.49141
R2043 VTAIL.n303 VTAIL.n302 3.49141
R2044 VTAIL.n259 VTAIL.n206 3.49141
R2045 VTAIL.n235 VTAIL.n234 3.49141
R2046 VTAIL.n269 VTAIL.n267 3.01774
R2047 VTAIL.n335 VTAIL.n269 3.01774
R2048 VTAIL.n403 VTAIL.n401 3.01774
R2049 VTAIL.n469 VTAIL.n403 3.01774
R2050 VTAIL.n201 VTAIL.n135 3.01774
R2051 VTAIL.n135 VTAIL.n133 3.01774
R2052 VTAIL.n67 VTAIL.n1 3.01774
R2053 VTAIL VTAIL.n535 2.95955
R2054 VTAIL.n505 VTAIL.n484 2.71565
R2055 VTAIL.n524 VTAIL.n523 2.71565
R2056 VTAIL.n37 VTAIL.n16 2.71565
R2057 VTAIL.n56 VTAIL.n55 2.71565
R2058 VTAIL.n103 VTAIL.n82 2.71565
R2059 VTAIL.n122 VTAIL.n121 2.71565
R2060 VTAIL.n171 VTAIL.n150 2.71565
R2061 VTAIL.n190 VTAIL.n189 2.71565
R2062 VTAIL.n458 VTAIL.n457 2.71565
R2063 VTAIL.n440 VTAIL.n419 2.71565
R2064 VTAIL.n390 VTAIL.n389 2.71565
R2065 VTAIL.n372 VTAIL.n351 2.71565
R2066 VTAIL.n324 VTAIL.n323 2.71565
R2067 VTAIL.n306 VTAIL.n285 2.71565
R2068 VTAIL.n256 VTAIL.n255 2.71565
R2069 VTAIL.n238 VTAIL.n217 2.71565
R2070 VTAIL.n0 VTAIL.t6 2.68022
R2071 VTAIL.n0 VTAIL.t5 2.68022
R2072 VTAIL.n134 VTAIL.t13 2.68022
R2073 VTAIL.n134 VTAIL.t12 2.68022
R2074 VTAIL.n402 VTAIL.t15 2.68022
R2075 VTAIL.n402 VTAIL.t8 2.68022
R2076 VTAIL.n268 VTAIL.t0 2.68022
R2077 VTAIL.n268 VTAIL.t4 2.68022
R2078 VTAIL.n427 VTAIL.n426 2.41282
R2079 VTAIL.n359 VTAIL.n358 2.41282
R2080 VTAIL.n293 VTAIL.n292 2.41282
R2081 VTAIL.n225 VTAIL.n224 2.41282
R2082 VTAIL.n492 VTAIL.n491 2.41282
R2083 VTAIL.n24 VTAIL.n23 2.41282
R2084 VTAIL.n90 VTAIL.n89 2.41282
R2085 VTAIL.n158 VTAIL.n157 2.41282
R2086 VTAIL.n506 VTAIL.n482 1.93989
R2087 VTAIL.n520 VTAIL.n476 1.93989
R2088 VTAIL.n38 VTAIL.n14 1.93989
R2089 VTAIL.n52 VTAIL.n8 1.93989
R2090 VTAIL.n104 VTAIL.n80 1.93989
R2091 VTAIL.n118 VTAIL.n74 1.93989
R2092 VTAIL.n172 VTAIL.n148 1.93989
R2093 VTAIL.n186 VTAIL.n142 1.93989
R2094 VTAIL.n454 VTAIL.n410 1.93989
R2095 VTAIL.n441 VTAIL.n417 1.93989
R2096 VTAIL.n386 VTAIL.n342 1.93989
R2097 VTAIL.n373 VTAIL.n349 1.93989
R2098 VTAIL.n320 VTAIL.n276 1.93989
R2099 VTAIL.n307 VTAIL.n283 1.93989
R2100 VTAIL.n252 VTAIL.n208 1.93989
R2101 VTAIL.n239 VTAIL.n215 1.93989
R2102 VTAIL.n511 VTAIL.n509 1.16414
R2103 VTAIL.n519 VTAIL.n478 1.16414
R2104 VTAIL.n43 VTAIL.n41 1.16414
R2105 VTAIL.n51 VTAIL.n10 1.16414
R2106 VTAIL.n109 VTAIL.n107 1.16414
R2107 VTAIL.n117 VTAIL.n76 1.16414
R2108 VTAIL.n177 VTAIL.n175 1.16414
R2109 VTAIL.n185 VTAIL.n144 1.16414
R2110 VTAIL.n453 VTAIL.n412 1.16414
R2111 VTAIL.n445 VTAIL.n444 1.16414
R2112 VTAIL.n385 VTAIL.n344 1.16414
R2113 VTAIL.n377 VTAIL.n376 1.16414
R2114 VTAIL.n319 VTAIL.n278 1.16414
R2115 VTAIL.n311 VTAIL.n310 1.16414
R2116 VTAIL.n251 VTAIL.n210 1.16414
R2117 VTAIL.n243 VTAIL.n242 1.16414
R2118 VTAIL.n401 VTAIL.n335 0.470328
R2119 VTAIL.n133 VTAIL.n67 0.470328
R2120 VTAIL.n510 VTAIL.n480 0.388379
R2121 VTAIL.n516 VTAIL.n515 0.388379
R2122 VTAIL.n42 VTAIL.n12 0.388379
R2123 VTAIL.n48 VTAIL.n47 0.388379
R2124 VTAIL.n108 VTAIL.n78 0.388379
R2125 VTAIL.n114 VTAIL.n113 0.388379
R2126 VTAIL.n176 VTAIL.n146 0.388379
R2127 VTAIL.n182 VTAIL.n181 0.388379
R2128 VTAIL.n450 VTAIL.n449 0.388379
R2129 VTAIL.n416 VTAIL.n414 0.388379
R2130 VTAIL.n382 VTAIL.n381 0.388379
R2131 VTAIL.n348 VTAIL.n346 0.388379
R2132 VTAIL.n316 VTAIL.n315 0.388379
R2133 VTAIL.n282 VTAIL.n280 0.388379
R2134 VTAIL.n248 VTAIL.n247 0.388379
R2135 VTAIL.n214 VTAIL.n212 0.388379
R2136 VTAIL.n492 VTAIL.n487 0.155672
R2137 VTAIL.n499 VTAIL.n487 0.155672
R2138 VTAIL.n500 VTAIL.n499 0.155672
R2139 VTAIL.n500 VTAIL.n483 0.155672
R2140 VTAIL.n507 VTAIL.n483 0.155672
R2141 VTAIL.n508 VTAIL.n507 0.155672
R2142 VTAIL.n508 VTAIL.n479 0.155672
R2143 VTAIL.n517 VTAIL.n479 0.155672
R2144 VTAIL.n518 VTAIL.n517 0.155672
R2145 VTAIL.n518 VTAIL.n475 0.155672
R2146 VTAIL.n525 VTAIL.n475 0.155672
R2147 VTAIL.n526 VTAIL.n525 0.155672
R2148 VTAIL.n526 VTAIL.n471 0.155672
R2149 VTAIL.n533 VTAIL.n471 0.155672
R2150 VTAIL.n24 VTAIL.n19 0.155672
R2151 VTAIL.n31 VTAIL.n19 0.155672
R2152 VTAIL.n32 VTAIL.n31 0.155672
R2153 VTAIL.n32 VTAIL.n15 0.155672
R2154 VTAIL.n39 VTAIL.n15 0.155672
R2155 VTAIL.n40 VTAIL.n39 0.155672
R2156 VTAIL.n40 VTAIL.n11 0.155672
R2157 VTAIL.n49 VTAIL.n11 0.155672
R2158 VTAIL.n50 VTAIL.n49 0.155672
R2159 VTAIL.n50 VTAIL.n7 0.155672
R2160 VTAIL.n57 VTAIL.n7 0.155672
R2161 VTAIL.n58 VTAIL.n57 0.155672
R2162 VTAIL.n58 VTAIL.n3 0.155672
R2163 VTAIL.n65 VTAIL.n3 0.155672
R2164 VTAIL.n90 VTAIL.n85 0.155672
R2165 VTAIL.n97 VTAIL.n85 0.155672
R2166 VTAIL.n98 VTAIL.n97 0.155672
R2167 VTAIL.n98 VTAIL.n81 0.155672
R2168 VTAIL.n105 VTAIL.n81 0.155672
R2169 VTAIL.n106 VTAIL.n105 0.155672
R2170 VTAIL.n106 VTAIL.n77 0.155672
R2171 VTAIL.n115 VTAIL.n77 0.155672
R2172 VTAIL.n116 VTAIL.n115 0.155672
R2173 VTAIL.n116 VTAIL.n73 0.155672
R2174 VTAIL.n123 VTAIL.n73 0.155672
R2175 VTAIL.n124 VTAIL.n123 0.155672
R2176 VTAIL.n124 VTAIL.n69 0.155672
R2177 VTAIL.n131 VTAIL.n69 0.155672
R2178 VTAIL.n158 VTAIL.n153 0.155672
R2179 VTAIL.n165 VTAIL.n153 0.155672
R2180 VTAIL.n166 VTAIL.n165 0.155672
R2181 VTAIL.n166 VTAIL.n149 0.155672
R2182 VTAIL.n173 VTAIL.n149 0.155672
R2183 VTAIL.n174 VTAIL.n173 0.155672
R2184 VTAIL.n174 VTAIL.n145 0.155672
R2185 VTAIL.n183 VTAIL.n145 0.155672
R2186 VTAIL.n184 VTAIL.n183 0.155672
R2187 VTAIL.n184 VTAIL.n141 0.155672
R2188 VTAIL.n191 VTAIL.n141 0.155672
R2189 VTAIL.n192 VTAIL.n191 0.155672
R2190 VTAIL.n192 VTAIL.n137 0.155672
R2191 VTAIL.n199 VTAIL.n137 0.155672
R2192 VTAIL.n467 VTAIL.n405 0.155672
R2193 VTAIL.n460 VTAIL.n405 0.155672
R2194 VTAIL.n460 VTAIL.n459 0.155672
R2195 VTAIL.n459 VTAIL.n409 0.155672
R2196 VTAIL.n452 VTAIL.n409 0.155672
R2197 VTAIL.n452 VTAIL.n451 0.155672
R2198 VTAIL.n451 VTAIL.n413 0.155672
R2199 VTAIL.n443 VTAIL.n413 0.155672
R2200 VTAIL.n443 VTAIL.n442 0.155672
R2201 VTAIL.n442 VTAIL.n418 0.155672
R2202 VTAIL.n435 VTAIL.n418 0.155672
R2203 VTAIL.n435 VTAIL.n434 0.155672
R2204 VTAIL.n434 VTAIL.n422 0.155672
R2205 VTAIL.n427 VTAIL.n422 0.155672
R2206 VTAIL.n399 VTAIL.n337 0.155672
R2207 VTAIL.n392 VTAIL.n337 0.155672
R2208 VTAIL.n392 VTAIL.n391 0.155672
R2209 VTAIL.n391 VTAIL.n341 0.155672
R2210 VTAIL.n384 VTAIL.n341 0.155672
R2211 VTAIL.n384 VTAIL.n383 0.155672
R2212 VTAIL.n383 VTAIL.n345 0.155672
R2213 VTAIL.n375 VTAIL.n345 0.155672
R2214 VTAIL.n375 VTAIL.n374 0.155672
R2215 VTAIL.n374 VTAIL.n350 0.155672
R2216 VTAIL.n367 VTAIL.n350 0.155672
R2217 VTAIL.n367 VTAIL.n366 0.155672
R2218 VTAIL.n366 VTAIL.n354 0.155672
R2219 VTAIL.n359 VTAIL.n354 0.155672
R2220 VTAIL.n333 VTAIL.n271 0.155672
R2221 VTAIL.n326 VTAIL.n271 0.155672
R2222 VTAIL.n326 VTAIL.n325 0.155672
R2223 VTAIL.n325 VTAIL.n275 0.155672
R2224 VTAIL.n318 VTAIL.n275 0.155672
R2225 VTAIL.n318 VTAIL.n317 0.155672
R2226 VTAIL.n317 VTAIL.n279 0.155672
R2227 VTAIL.n309 VTAIL.n279 0.155672
R2228 VTAIL.n309 VTAIL.n308 0.155672
R2229 VTAIL.n308 VTAIL.n284 0.155672
R2230 VTAIL.n301 VTAIL.n284 0.155672
R2231 VTAIL.n301 VTAIL.n300 0.155672
R2232 VTAIL.n300 VTAIL.n288 0.155672
R2233 VTAIL.n293 VTAIL.n288 0.155672
R2234 VTAIL.n265 VTAIL.n203 0.155672
R2235 VTAIL.n258 VTAIL.n203 0.155672
R2236 VTAIL.n258 VTAIL.n257 0.155672
R2237 VTAIL.n257 VTAIL.n207 0.155672
R2238 VTAIL.n250 VTAIL.n207 0.155672
R2239 VTAIL.n250 VTAIL.n249 0.155672
R2240 VTAIL.n249 VTAIL.n211 0.155672
R2241 VTAIL.n241 VTAIL.n211 0.155672
R2242 VTAIL.n241 VTAIL.n240 0.155672
R2243 VTAIL.n240 VTAIL.n216 0.155672
R2244 VTAIL.n233 VTAIL.n216 0.155672
R2245 VTAIL.n233 VTAIL.n232 0.155672
R2246 VTAIL.n232 VTAIL.n220 0.155672
R2247 VTAIL.n225 VTAIL.n220 0.155672
R2248 VTAIL VTAIL.n1 0.0586897
R2249 VDD1 VDD1.n0 75.6
R2250 VDD1.n3 VDD1.n2 75.4862
R2251 VDD1.n3 VDD1.n1 75.4862
R2252 VDD1.n5 VDD1.n4 74.033
R2253 VDD1.n5 VDD1.n3 48.3328
R2254 VDD1.n4 VDD1.t1 2.68022
R2255 VDD1.n4 VDD1.t2 2.68022
R2256 VDD1.n0 VDD1.t5 2.68022
R2257 VDD1.n0 VDD1.t6 2.68022
R2258 VDD1.n2 VDD1.t4 2.68022
R2259 VDD1.n2 VDD1.t7 2.68022
R2260 VDD1.n1 VDD1.t0 2.68022
R2261 VDD1.n1 VDD1.t3 2.68022
R2262 VDD1 VDD1.n5 1.45093
R2263 VN.n64 VN.n63 161.3
R2264 VN.n62 VN.n34 161.3
R2265 VN.n61 VN.n60 161.3
R2266 VN.n59 VN.n35 161.3
R2267 VN.n58 VN.n57 161.3
R2268 VN.n56 VN.n36 161.3
R2269 VN.n55 VN.n54 161.3
R2270 VN.n53 VN.n52 161.3
R2271 VN.n51 VN.n38 161.3
R2272 VN.n50 VN.n49 161.3
R2273 VN.n48 VN.n39 161.3
R2274 VN.n47 VN.n46 161.3
R2275 VN.n45 VN.n40 161.3
R2276 VN.n44 VN.n43 161.3
R2277 VN.n31 VN.n30 161.3
R2278 VN.n29 VN.n1 161.3
R2279 VN.n28 VN.n27 161.3
R2280 VN.n26 VN.n2 161.3
R2281 VN.n25 VN.n24 161.3
R2282 VN.n23 VN.n3 161.3
R2283 VN.n22 VN.n21 161.3
R2284 VN.n20 VN.n19 161.3
R2285 VN.n18 VN.n5 161.3
R2286 VN.n17 VN.n16 161.3
R2287 VN.n15 VN.n6 161.3
R2288 VN.n14 VN.n13 161.3
R2289 VN.n12 VN.n7 161.3
R2290 VN.n11 VN.n10 161.3
R2291 VN.n42 VN.t3 124.856
R2292 VN.n9 VN.t7 124.856
R2293 VN.n8 VN.t2 92.2191
R2294 VN.n4 VN.t4 92.2191
R2295 VN.n0 VN.t5 92.2191
R2296 VN.n41 VN.t0 92.2191
R2297 VN.n37 VN.t1 92.2191
R2298 VN.n33 VN.t6 92.2191
R2299 VN.n32 VN.n0 77.8339
R2300 VN.n65 VN.n33 77.8339
R2301 VN.n9 VN.n8 62.0322
R2302 VN.n42 VN.n41 62.0322
R2303 VN VN.n65 53.8692
R2304 VN.n13 VN.n6 40.4934
R2305 VN.n17 VN.n6 40.4934
R2306 VN.n24 VN.n2 40.4934
R2307 VN.n28 VN.n2 40.4934
R2308 VN.n46 VN.n39 40.4934
R2309 VN.n50 VN.n39 40.4934
R2310 VN.n57 VN.n35 40.4934
R2311 VN.n61 VN.n35 40.4934
R2312 VN.n12 VN.n11 24.4675
R2313 VN.n13 VN.n12 24.4675
R2314 VN.n18 VN.n17 24.4675
R2315 VN.n19 VN.n18 24.4675
R2316 VN.n23 VN.n22 24.4675
R2317 VN.n24 VN.n23 24.4675
R2318 VN.n29 VN.n28 24.4675
R2319 VN.n30 VN.n29 24.4675
R2320 VN.n46 VN.n45 24.4675
R2321 VN.n45 VN.n44 24.4675
R2322 VN.n57 VN.n56 24.4675
R2323 VN.n56 VN.n55 24.4675
R2324 VN.n52 VN.n51 24.4675
R2325 VN.n51 VN.n50 24.4675
R2326 VN.n63 VN.n62 24.4675
R2327 VN.n62 VN.n61 24.4675
R2328 VN.n11 VN.n8 12.234
R2329 VN.n19 VN.n4 12.234
R2330 VN.n22 VN.n4 12.234
R2331 VN.n30 VN.n0 12.234
R2332 VN.n44 VN.n41 12.234
R2333 VN.n55 VN.n37 12.234
R2334 VN.n52 VN.n37 12.234
R2335 VN.n63 VN.n33 12.234
R2336 VN.n10 VN.n9 4.27758
R2337 VN.n43 VN.n42 4.27758
R2338 VN.n65 VN.n64 0.354971
R2339 VN.n32 VN.n31 0.354971
R2340 VN VN.n32 0.26696
R2341 VN.n64 VN.n34 0.189894
R2342 VN.n60 VN.n34 0.189894
R2343 VN.n60 VN.n59 0.189894
R2344 VN.n59 VN.n58 0.189894
R2345 VN.n58 VN.n36 0.189894
R2346 VN.n54 VN.n36 0.189894
R2347 VN.n54 VN.n53 0.189894
R2348 VN.n53 VN.n38 0.189894
R2349 VN.n49 VN.n38 0.189894
R2350 VN.n49 VN.n48 0.189894
R2351 VN.n48 VN.n47 0.189894
R2352 VN.n47 VN.n40 0.189894
R2353 VN.n43 VN.n40 0.189894
R2354 VN.n10 VN.n7 0.189894
R2355 VN.n14 VN.n7 0.189894
R2356 VN.n15 VN.n14 0.189894
R2357 VN.n16 VN.n15 0.189894
R2358 VN.n16 VN.n5 0.189894
R2359 VN.n20 VN.n5 0.189894
R2360 VN.n21 VN.n20 0.189894
R2361 VN.n21 VN.n3 0.189894
R2362 VN.n25 VN.n3 0.189894
R2363 VN.n26 VN.n25 0.189894
R2364 VN.n27 VN.n26 0.189894
R2365 VN.n27 VN.n1 0.189894
R2366 VN.n31 VN.n1 0.189894
R2367 VDD2.n2 VDD2.n1 75.4862
R2368 VDD2.n2 VDD2.n0 75.4862
R2369 VDD2 VDD2.n5 75.4834
R2370 VDD2.n4 VDD2.n3 74.0332
R2371 VDD2.n4 VDD2.n2 47.7498
R2372 VDD2.n5 VDD2.t7 2.68022
R2373 VDD2.n5 VDD2.t4 2.68022
R2374 VDD2.n3 VDD2.t1 2.68022
R2375 VDD2.n3 VDD2.t6 2.68022
R2376 VDD2.n1 VDD2.t3 2.68022
R2377 VDD2.n1 VDD2.t2 2.68022
R2378 VDD2.n0 VDD2.t0 2.68022
R2379 VDD2.n0 VDD2.t5 2.68022
R2380 VDD2 VDD2.n4 1.56731
C0 w_n4470_n3394# VP 9.859179f
C1 B VTAIL 5.27303f
C2 w_n4470_n3394# VN 9.277201f
C3 B VP 2.33803f
C4 VP VTAIL 9.70109f
C5 B VN 1.35939f
C6 VDD1 w_n4470_n3394# 2.13462f
C7 VN VTAIL 9.686991f
C8 VDD1 B 1.82642f
C9 VP VN 8.38855f
C10 VDD2 w_n4470_n3394# 2.27324f
C11 VDD1 VTAIL 8.30332f
C12 VDD2 B 1.94038f
C13 VDD1 VP 9.53685f
C14 VDD2 VTAIL 8.36156f
C15 VDD1 VN 0.152283f
C16 VDD2 VP 0.579849f
C17 VDD2 VN 9.11096f
C18 VDD1 VDD2 2.07101f
C19 w_n4470_n3394# B 11.0247f
C20 w_n4470_n3394# VTAIL 4.2815f
C21 VDD2 VSUBS 2.190166f
C22 VDD1 VSUBS 2.93048f
C23 VTAIL VSUBS 1.44465f
C24 VN VSUBS 7.50389f
C25 VP VSUBS 4.176874f
C26 B VSUBS 5.650599f
C27 w_n4470_n3394# VSUBS 0.186721p
C28 VDD2.t0 VSUBS 0.290142f
C29 VDD2.t5 VSUBS 0.290142f
C30 VDD2.n0 VSUBS 2.28807f
C31 VDD2.t3 VSUBS 0.290142f
C32 VDD2.t2 VSUBS 0.290142f
C33 VDD2.n1 VSUBS 2.28807f
C34 VDD2.n2 VSUBS 5.01075f
C35 VDD2.t1 VSUBS 0.290142f
C36 VDD2.t6 VSUBS 0.290142f
C37 VDD2.n3 VSUBS 2.26848f
C38 VDD2.n4 VSUBS 4.1435f
C39 VDD2.t7 VSUBS 0.290142f
C40 VDD2.t4 VSUBS 0.290142f
C41 VDD2.n5 VSUBS 2.28802f
C42 VN.t5 VSUBS 2.73907f
C43 VN.n0 VSUBS 1.05821f
C44 VN.n1 VSUBS 0.026136f
C45 VN.n2 VSUBS 0.021129f
C46 VN.n3 VSUBS 0.026136f
C47 VN.t4 VSUBS 2.73907f
C48 VN.n4 VSUBS 0.96287f
C49 VN.n5 VSUBS 0.026136f
C50 VN.n6 VSUBS 0.021129f
C51 VN.n7 VSUBS 0.026136f
C52 VN.t2 VSUBS 2.73907f
C53 VN.n8 VSUBS 1.04852f
C54 VN.t7 VSUBS 3.03791f
C55 VN.n9 VSUBS 1.00285f
C56 VN.n10 VSUBS 0.303865f
C57 VN.n11 VSUBS 0.036687f
C58 VN.n12 VSUBS 0.048711f
C59 VN.n13 VSUBS 0.051946f
C60 VN.n14 VSUBS 0.026136f
C61 VN.n15 VSUBS 0.026136f
C62 VN.n16 VSUBS 0.026136f
C63 VN.n17 VSUBS 0.051946f
C64 VN.n18 VSUBS 0.048711f
C65 VN.n19 VSUBS 0.036687f
C66 VN.n20 VSUBS 0.026136f
C67 VN.n21 VSUBS 0.026136f
C68 VN.n22 VSUBS 0.036687f
C69 VN.n23 VSUBS 0.048711f
C70 VN.n24 VSUBS 0.051946f
C71 VN.n25 VSUBS 0.026136f
C72 VN.n26 VSUBS 0.026136f
C73 VN.n27 VSUBS 0.026136f
C74 VN.n28 VSUBS 0.051946f
C75 VN.n29 VSUBS 0.048711f
C76 VN.n30 VSUBS 0.036687f
C77 VN.n31 VSUBS 0.042183f
C78 VN.n32 VSUBS 0.064182f
C79 VN.t6 VSUBS 2.73907f
C80 VN.n33 VSUBS 1.05821f
C81 VN.n34 VSUBS 0.026136f
C82 VN.n35 VSUBS 0.021129f
C83 VN.n36 VSUBS 0.026136f
C84 VN.t1 VSUBS 2.73907f
C85 VN.n37 VSUBS 0.96287f
C86 VN.n38 VSUBS 0.026136f
C87 VN.n39 VSUBS 0.021129f
C88 VN.n40 VSUBS 0.026136f
C89 VN.t0 VSUBS 2.73907f
C90 VN.n41 VSUBS 1.04852f
C91 VN.t3 VSUBS 3.03791f
C92 VN.n42 VSUBS 1.00285f
C93 VN.n43 VSUBS 0.303865f
C94 VN.n44 VSUBS 0.036687f
C95 VN.n45 VSUBS 0.048711f
C96 VN.n46 VSUBS 0.051946f
C97 VN.n47 VSUBS 0.026136f
C98 VN.n48 VSUBS 0.026136f
C99 VN.n49 VSUBS 0.026136f
C100 VN.n50 VSUBS 0.051946f
C101 VN.n51 VSUBS 0.048711f
C102 VN.n52 VSUBS 0.036687f
C103 VN.n53 VSUBS 0.026136f
C104 VN.n54 VSUBS 0.026136f
C105 VN.n55 VSUBS 0.036687f
C106 VN.n56 VSUBS 0.048711f
C107 VN.n57 VSUBS 0.051946f
C108 VN.n58 VSUBS 0.026136f
C109 VN.n59 VSUBS 0.026136f
C110 VN.n60 VSUBS 0.026136f
C111 VN.n61 VSUBS 0.051946f
C112 VN.n62 VSUBS 0.048711f
C113 VN.n63 VSUBS 0.036687f
C114 VN.n64 VSUBS 0.042183f
C115 VN.n65 VSUBS 1.65446f
C116 VDD1.t5 VSUBS 0.289986f
C117 VDD1.t6 VSUBS 0.289986f
C118 VDD1.n0 VSUBS 2.28857f
C119 VDD1.t0 VSUBS 0.289986f
C120 VDD1.t3 VSUBS 0.289986f
C121 VDD1.n1 VSUBS 2.28685f
C122 VDD1.t4 VSUBS 0.289986f
C123 VDD1.t7 VSUBS 0.289986f
C124 VDD1.n2 VSUBS 2.28685f
C125 VDD1.n3 VSUBS 5.0707f
C126 VDD1.t1 VSUBS 0.289986f
C127 VDD1.t2 VSUBS 0.289986f
C128 VDD1.n4 VSUBS 2.26726f
C129 VDD1.n5 VSUBS 4.17904f
C130 VTAIL.t6 VSUBS 0.245527f
C131 VTAIL.t5 VSUBS 0.245527f
C132 VTAIL.n0 VSUBS 1.78098f
C133 VTAIL.n1 VSUBS 0.839448f
C134 VTAIL.n2 VSUBS 0.028146f
C135 VTAIL.n3 VSUBS 0.025615f
C136 VTAIL.n4 VSUBS 0.013764f
C137 VTAIL.n5 VSUBS 0.032533f
C138 VTAIL.n6 VSUBS 0.014574f
C139 VTAIL.n7 VSUBS 0.025615f
C140 VTAIL.n8 VSUBS 0.013764f
C141 VTAIL.n9 VSUBS 0.032533f
C142 VTAIL.n10 VSUBS 0.014574f
C143 VTAIL.n11 VSUBS 0.025615f
C144 VTAIL.n12 VSUBS 0.014169f
C145 VTAIL.n13 VSUBS 0.032533f
C146 VTAIL.n14 VSUBS 0.014574f
C147 VTAIL.n15 VSUBS 0.025615f
C148 VTAIL.n16 VSUBS 0.013764f
C149 VTAIL.n17 VSUBS 0.032533f
C150 VTAIL.n18 VSUBS 0.014574f
C151 VTAIL.n19 VSUBS 0.025615f
C152 VTAIL.n20 VSUBS 0.013764f
C153 VTAIL.n21 VSUBS 0.0244f
C154 VTAIL.n22 VSUBS 0.024473f
C155 VTAIL.t1 VSUBS 0.070117f
C156 VTAIL.n23 VSUBS 0.203235f
C157 VTAIL.n24 VSUBS 1.27311f
C158 VTAIL.n25 VSUBS 0.013764f
C159 VTAIL.n26 VSUBS 0.014574f
C160 VTAIL.n27 VSUBS 0.032533f
C161 VTAIL.n28 VSUBS 0.032533f
C162 VTAIL.n29 VSUBS 0.014574f
C163 VTAIL.n30 VSUBS 0.013764f
C164 VTAIL.n31 VSUBS 0.025615f
C165 VTAIL.n32 VSUBS 0.025615f
C166 VTAIL.n33 VSUBS 0.013764f
C167 VTAIL.n34 VSUBS 0.014574f
C168 VTAIL.n35 VSUBS 0.032533f
C169 VTAIL.n36 VSUBS 0.032533f
C170 VTAIL.n37 VSUBS 0.014574f
C171 VTAIL.n38 VSUBS 0.013764f
C172 VTAIL.n39 VSUBS 0.025615f
C173 VTAIL.n40 VSUBS 0.025615f
C174 VTAIL.n41 VSUBS 0.013764f
C175 VTAIL.n42 VSUBS 0.013764f
C176 VTAIL.n43 VSUBS 0.014574f
C177 VTAIL.n44 VSUBS 0.032533f
C178 VTAIL.n45 VSUBS 0.032533f
C179 VTAIL.n46 VSUBS 0.032533f
C180 VTAIL.n47 VSUBS 0.014169f
C181 VTAIL.n48 VSUBS 0.013764f
C182 VTAIL.n49 VSUBS 0.025615f
C183 VTAIL.n50 VSUBS 0.025615f
C184 VTAIL.n51 VSUBS 0.013764f
C185 VTAIL.n52 VSUBS 0.014574f
C186 VTAIL.n53 VSUBS 0.032533f
C187 VTAIL.n54 VSUBS 0.032533f
C188 VTAIL.n55 VSUBS 0.014574f
C189 VTAIL.n56 VSUBS 0.013764f
C190 VTAIL.n57 VSUBS 0.025615f
C191 VTAIL.n58 VSUBS 0.025615f
C192 VTAIL.n59 VSUBS 0.013764f
C193 VTAIL.n60 VSUBS 0.014574f
C194 VTAIL.n61 VSUBS 0.032533f
C195 VTAIL.n62 VSUBS 0.078765f
C196 VTAIL.n63 VSUBS 0.014574f
C197 VTAIL.n64 VSUBS 0.013764f
C198 VTAIL.n65 VSUBS 0.059557f
C199 VTAIL.n66 VSUBS 0.039621f
C200 VTAIL.n67 VSUBS 0.309881f
C201 VTAIL.n68 VSUBS 0.028146f
C202 VTAIL.n69 VSUBS 0.025615f
C203 VTAIL.n70 VSUBS 0.013764f
C204 VTAIL.n71 VSUBS 0.032533f
C205 VTAIL.n72 VSUBS 0.014574f
C206 VTAIL.n73 VSUBS 0.025615f
C207 VTAIL.n74 VSUBS 0.013764f
C208 VTAIL.n75 VSUBS 0.032533f
C209 VTAIL.n76 VSUBS 0.014574f
C210 VTAIL.n77 VSUBS 0.025615f
C211 VTAIL.n78 VSUBS 0.014169f
C212 VTAIL.n79 VSUBS 0.032533f
C213 VTAIL.n80 VSUBS 0.014574f
C214 VTAIL.n81 VSUBS 0.025615f
C215 VTAIL.n82 VSUBS 0.013764f
C216 VTAIL.n83 VSUBS 0.032533f
C217 VTAIL.n84 VSUBS 0.014574f
C218 VTAIL.n85 VSUBS 0.025615f
C219 VTAIL.n86 VSUBS 0.013764f
C220 VTAIL.n87 VSUBS 0.0244f
C221 VTAIL.n88 VSUBS 0.024473f
C222 VTAIL.t9 VSUBS 0.070117f
C223 VTAIL.n89 VSUBS 0.203235f
C224 VTAIL.n90 VSUBS 1.27311f
C225 VTAIL.n91 VSUBS 0.013764f
C226 VTAIL.n92 VSUBS 0.014574f
C227 VTAIL.n93 VSUBS 0.032533f
C228 VTAIL.n94 VSUBS 0.032533f
C229 VTAIL.n95 VSUBS 0.014574f
C230 VTAIL.n96 VSUBS 0.013764f
C231 VTAIL.n97 VSUBS 0.025615f
C232 VTAIL.n98 VSUBS 0.025615f
C233 VTAIL.n99 VSUBS 0.013764f
C234 VTAIL.n100 VSUBS 0.014574f
C235 VTAIL.n101 VSUBS 0.032533f
C236 VTAIL.n102 VSUBS 0.032533f
C237 VTAIL.n103 VSUBS 0.014574f
C238 VTAIL.n104 VSUBS 0.013764f
C239 VTAIL.n105 VSUBS 0.025615f
C240 VTAIL.n106 VSUBS 0.025615f
C241 VTAIL.n107 VSUBS 0.013764f
C242 VTAIL.n108 VSUBS 0.013764f
C243 VTAIL.n109 VSUBS 0.014574f
C244 VTAIL.n110 VSUBS 0.032533f
C245 VTAIL.n111 VSUBS 0.032533f
C246 VTAIL.n112 VSUBS 0.032533f
C247 VTAIL.n113 VSUBS 0.014169f
C248 VTAIL.n114 VSUBS 0.013764f
C249 VTAIL.n115 VSUBS 0.025615f
C250 VTAIL.n116 VSUBS 0.025615f
C251 VTAIL.n117 VSUBS 0.013764f
C252 VTAIL.n118 VSUBS 0.014574f
C253 VTAIL.n119 VSUBS 0.032533f
C254 VTAIL.n120 VSUBS 0.032533f
C255 VTAIL.n121 VSUBS 0.014574f
C256 VTAIL.n122 VSUBS 0.013764f
C257 VTAIL.n123 VSUBS 0.025615f
C258 VTAIL.n124 VSUBS 0.025615f
C259 VTAIL.n125 VSUBS 0.013764f
C260 VTAIL.n126 VSUBS 0.014574f
C261 VTAIL.n127 VSUBS 0.032533f
C262 VTAIL.n128 VSUBS 0.078765f
C263 VTAIL.n129 VSUBS 0.014574f
C264 VTAIL.n130 VSUBS 0.013764f
C265 VTAIL.n131 VSUBS 0.059557f
C266 VTAIL.n132 VSUBS 0.039621f
C267 VTAIL.n133 VSUBS 0.309881f
C268 VTAIL.t13 VSUBS 0.245527f
C269 VTAIL.t12 VSUBS 0.245527f
C270 VTAIL.n134 VSUBS 1.78098f
C271 VTAIL.n135 VSUBS 1.08367f
C272 VTAIL.n136 VSUBS 0.028146f
C273 VTAIL.n137 VSUBS 0.025615f
C274 VTAIL.n138 VSUBS 0.013764f
C275 VTAIL.n139 VSUBS 0.032533f
C276 VTAIL.n140 VSUBS 0.014574f
C277 VTAIL.n141 VSUBS 0.025615f
C278 VTAIL.n142 VSUBS 0.013764f
C279 VTAIL.n143 VSUBS 0.032533f
C280 VTAIL.n144 VSUBS 0.014574f
C281 VTAIL.n145 VSUBS 0.025615f
C282 VTAIL.n146 VSUBS 0.014169f
C283 VTAIL.n147 VSUBS 0.032533f
C284 VTAIL.n148 VSUBS 0.014574f
C285 VTAIL.n149 VSUBS 0.025615f
C286 VTAIL.n150 VSUBS 0.013764f
C287 VTAIL.n151 VSUBS 0.032533f
C288 VTAIL.n152 VSUBS 0.014574f
C289 VTAIL.n153 VSUBS 0.025615f
C290 VTAIL.n154 VSUBS 0.013764f
C291 VTAIL.n155 VSUBS 0.0244f
C292 VTAIL.n156 VSUBS 0.024473f
C293 VTAIL.t10 VSUBS 0.070117f
C294 VTAIL.n157 VSUBS 0.203235f
C295 VTAIL.n158 VSUBS 1.27311f
C296 VTAIL.n159 VSUBS 0.013764f
C297 VTAIL.n160 VSUBS 0.014574f
C298 VTAIL.n161 VSUBS 0.032533f
C299 VTAIL.n162 VSUBS 0.032533f
C300 VTAIL.n163 VSUBS 0.014574f
C301 VTAIL.n164 VSUBS 0.013764f
C302 VTAIL.n165 VSUBS 0.025615f
C303 VTAIL.n166 VSUBS 0.025615f
C304 VTAIL.n167 VSUBS 0.013764f
C305 VTAIL.n168 VSUBS 0.014574f
C306 VTAIL.n169 VSUBS 0.032533f
C307 VTAIL.n170 VSUBS 0.032533f
C308 VTAIL.n171 VSUBS 0.014574f
C309 VTAIL.n172 VSUBS 0.013764f
C310 VTAIL.n173 VSUBS 0.025615f
C311 VTAIL.n174 VSUBS 0.025615f
C312 VTAIL.n175 VSUBS 0.013764f
C313 VTAIL.n176 VSUBS 0.013764f
C314 VTAIL.n177 VSUBS 0.014574f
C315 VTAIL.n178 VSUBS 0.032533f
C316 VTAIL.n179 VSUBS 0.032533f
C317 VTAIL.n180 VSUBS 0.032533f
C318 VTAIL.n181 VSUBS 0.014169f
C319 VTAIL.n182 VSUBS 0.013764f
C320 VTAIL.n183 VSUBS 0.025615f
C321 VTAIL.n184 VSUBS 0.025615f
C322 VTAIL.n185 VSUBS 0.013764f
C323 VTAIL.n186 VSUBS 0.014574f
C324 VTAIL.n187 VSUBS 0.032533f
C325 VTAIL.n188 VSUBS 0.032533f
C326 VTAIL.n189 VSUBS 0.014574f
C327 VTAIL.n190 VSUBS 0.013764f
C328 VTAIL.n191 VSUBS 0.025615f
C329 VTAIL.n192 VSUBS 0.025615f
C330 VTAIL.n193 VSUBS 0.013764f
C331 VTAIL.n194 VSUBS 0.014574f
C332 VTAIL.n195 VSUBS 0.032533f
C333 VTAIL.n196 VSUBS 0.078765f
C334 VTAIL.n197 VSUBS 0.014574f
C335 VTAIL.n198 VSUBS 0.013764f
C336 VTAIL.n199 VSUBS 0.059557f
C337 VTAIL.n200 VSUBS 0.039621f
C338 VTAIL.n201 VSUBS 1.73114f
C339 VTAIL.n202 VSUBS 0.028146f
C340 VTAIL.n203 VSUBS 0.025615f
C341 VTAIL.n204 VSUBS 0.013764f
C342 VTAIL.n205 VSUBS 0.032533f
C343 VTAIL.n206 VSUBS 0.014574f
C344 VTAIL.n207 VSUBS 0.025615f
C345 VTAIL.n208 VSUBS 0.013764f
C346 VTAIL.n209 VSUBS 0.032533f
C347 VTAIL.n210 VSUBS 0.014574f
C348 VTAIL.n211 VSUBS 0.025615f
C349 VTAIL.n212 VSUBS 0.014169f
C350 VTAIL.n213 VSUBS 0.032533f
C351 VTAIL.n214 VSUBS 0.013764f
C352 VTAIL.n215 VSUBS 0.014574f
C353 VTAIL.n216 VSUBS 0.025615f
C354 VTAIL.n217 VSUBS 0.013764f
C355 VTAIL.n218 VSUBS 0.032533f
C356 VTAIL.n219 VSUBS 0.014574f
C357 VTAIL.n220 VSUBS 0.025615f
C358 VTAIL.n221 VSUBS 0.013764f
C359 VTAIL.n222 VSUBS 0.0244f
C360 VTAIL.n223 VSUBS 0.024473f
C361 VTAIL.t7 VSUBS 0.070117f
C362 VTAIL.n224 VSUBS 0.203235f
C363 VTAIL.n225 VSUBS 1.27311f
C364 VTAIL.n226 VSUBS 0.013764f
C365 VTAIL.n227 VSUBS 0.014574f
C366 VTAIL.n228 VSUBS 0.032533f
C367 VTAIL.n229 VSUBS 0.032533f
C368 VTAIL.n230 VSUBS 0.014574f
C369 VTAIL.n231 VSUBS 0.013764f
C370 VTAIL.n232 VSUBS 0.025615f
C371 VTAIL.n233 VSUBS 0.025615f
C372 VTAIL.n234 VSUBS 0.013764f
C373 VTAIL.n235 VSUBS 0.014574f
C374 VTAIL.n236 VSUBS 0.032533f
C375 VTAIL.n237 VSUBS 0.032533f
C376 VTAIL.n238 VSUBS 0.014574f
C377 VTAIL.n239 VSUBS 0.013764f
C378 VTAIL.n240 VSUBS 0.025615f
C379 VTAIL.n241 VSUBS 0.025615f
C380 VTAIL.n242 VSUBS 0.013764f
C381 VTAIL.n243 VSUBS 0.014574f
C382 VTAIL.n244 VSUBS 0.032533f
C383 VTAIL.n245 VSUBS 0.032533f
C384 VTAIL.n246 VSUBS 0.032533f
C385 VTAIL.n247 VSUBS 0.014169f
C386 VTAIL.n248 VSUBS 0.013764f
C387 VTAIL.n249 VSUBS 0.025615f
C388 VTAIL.n250 VSUBS 0.025615f
C389 VTAIL.n251 VSUBS 0.013764f
C390 VTAIL.n252 VSUBS 0.014574f
C391 VTAIL.n253 VSUBS 0.032533f
C392 VTAIL.n254 VSUBS 0.032533f
C393 VTAIL.n255 VSUBS 0.014574f
C394 VTAIL.n256 VSUBS 0.013764f
C395 VTAIL.n257 VSUBS 0.025615f
C396 VTAIL.n258 VSUBS 0.025615f
C397 VTAIL.n259 VSUBS 0.013764f
C398 VTAIL.n260 VSUBS 0.014574f
C399 VTAIL.n261 VSUBS 0.032533f
C400 VTAIL.n262 VSUBS 0.078765f
C401 VTAIL.n263 VSUBS 0.014574f
C402 VTAIL.n264 VSUBS 0.013764f
C403 VTAIL.n265 VSUBS 0.059557f
C404 VTAIL.n266 VSUBS 0.039621f
C405 VTAIL.n267 VSUBS 1.73114f
C406 VTAIL.t0 VSUBS 0.245527f
C407 VTAIL.t4 VSUBS 0.245527f
C408 VTAIL.n268 VSUBS 1.78099f
C409 VTAIL.n269 VSUBS 1.08366f
C410 VTAIL.n270 VSUBS 0.028146f
C411 VTAIL.n271 VSUBS 0.025615f
C412 VTAIL.n272 VSUBS 0.013764f
C413 VTAIL.n273 VSUBS 0.032533f
C414 VTAIL.n274 VSUBS 0.014574f
C415 VTAIL.n275 VSUBS 0.025615f
C416 VTAIL.n276 VSUBS 0.013764f
C417 VTAIL.n277 VSUBS 0.032533f
C418 VTAIL.n278 VSUBS 0.014574f
C419 VTAIL.n279 VSUBS 0.025615f
C420 VTAIL.n280 VSUBS 0.014169f
C421 VTAIL.n281 VSUBS 0.032533f
C422 VTAIL.n282 VSUBS 0.013764f
C423 VTAIL.n283 VSUBS 0.014574f
C424 VTAIL.n284 VSUBS 0.025615f
C425 VTAIL.n285 VSUBS 0.013764f
C426 VTAIL.n286 VSUBS 0.032533f
C427 VTAIL.n287 VSUBS 0.014574f
C428 VTAIL.n288 VSUBS 0.025615f
C429 VTAIL.n289 VSUBS 0.013764f
C430 VTAIL.n290 VSUBS 0.0244f
C431 VTAIL.n291 VSUBS 0.024473f
C432 VTAIL.t3 VSUBS 0.070117f
C433 VTAIL.n292 VSUBS 0.203235f
C434 VTAIL.n293 VSUBS 1.27311f
C435 VTAIL.n294 VSUBS 0.013764f
C436 VTAIL.n295 VSUBS 0.014574f
C437 VTAIL.n296 VSUBS 0.032533f
C438 VTAIL.n297 VSUBS 0.032533f
C439 VTAIL.n298 VSUBS 0.014574f
C440 VTAIL.n299 VSUBS 0.013764f
C441 VTAIL.n300 VSUBS 0.025615f
C442 VTAIL.n301 VSUBS 0.025615f
C443 VTAIL.n302 VSUBS 0.013764f
C444 VTAIL.n303 VSUBS 0.014574f
C445 VTAIL.n304 VSUBS 0.032533f
C446 VTAIL.n305 VSUBS 0.032533f
C447 VTAIL.n306 VSUBS 0.014574f
C448 VTAIL.n307 VSUBS 0.013764f
C449 VTAIL.n308 VSUBS 0.025615f
C450 VTAIL.n309 VSUBS 0.025615f
C451 VTAIL.n310 VSUBS 0.013764f
C452 VTAIL.n311 VSUBS 0.014574f
C453 VTAIL.n312 VSUBS 0.032533f
C454 VTAIL.n313 VSUBS 0.032533f
C455 VTAIL.n314 VSUBS 0.032533f
C456 VTAIL.n315 VSUBS 0.014169f
C457 VTAIL.n316 VSUBS 0.013764f
C458 VTAIL.n317 VSUBS 0.025615f
C459 VTAIL.n318 VSUBS 0.025615f
C460 VTAIL.n319 VSUBS 0.013764f
C461 VTAIL.n320 VSUBS 0.014574f
C462 VTAIL.n321 VSUBS 0.032533f
C463 VTAIL.n322 VSUBS 0.032533f
C464 VTAIL.n323 VSUBS 0.014574f
C465 VTAIL.n324 VSUBS 0.013764f
C466 VTAIL.n325 VSUBS 0.025615f
C467 VTAIL.n326 VSUBS 0.025615f
C468 VTAIL.n327 VSUBS 0.013764f
C469 VTAIL.n328 VSUBS 0.014574f
C470 VTAIL.n329 VSUBS 0.032533f
C471 VTAIL.n330 VSUBS 0.078765f
C472 VTAIL.n331 VSUBS 0.014574f
C473 VTAIL.n332 VSUBS 0.013764f
C474 VTAIL.n333 VSUBS 0.059557f
C475 VTAIL.n334 VSUBS 0.039621f
C476 VTAIL.n335 VSUBS 0.309881f
C477 VTAIL.n336 VSUBS 0.028146f
C478 VTAIL.n337 VSUBS 0.025615f
C479 VTAIL.n338 VSUBS 0.013764f
C480 VTAIL.n339 VSUBS 0.032533f
C481 VTAIL.n340 VSUBS 0.014574f
C482 VTAIL.n341 VSUBS 0.025615f
C483 VTAIL.n342 VSUBS 0.013764f
C484 VTAIL.n343 VSUBS 0.032533f
C485 VTAIL.n344 VSUBS 0.014574f
C486 VTAIL.n345 VSUBS 0.025615f
C487 VTAIL.n346 VSUBS 0.014169f
C488 VTAIL.n347 VSUBS 0.032533f
C489 VTAIL.n348 VSUBS 0.013764f
C490 VTAIL.n349 VSUBS 0.014574f
C491 VTAIL.n350 VSUBS 0.025615f
C492 VTAIL.n351 VSUBS 0.013764f
C493 VTAIL.n352 VSUBS 0.032533f
C494 VTAIL.n353 VSUBS 0.014574f
C495 VTAIL.n354 VSUBS 0.025615f
C496 VTAIL.n355 VSUBS 0.013764f
C497 VTAIL.n356 VSUBS 0.0244f
C498 VTAIL.n357 VSUBS 0.024473f
C499 VTAIL.t11 VSUBS 0.070117f
C500 VTAIL.n358 VSUBS 0.203235f
C501 VTAIL.n359 VSUBS 1.27311f
C502 VTAIL.n360 VSUBS 0.013764f
C503 VTAIL.n361 VSUBS 0.014574f
C504 VTAIL.n362 VSUBS 0.032533f
C505 VTAIL.n363 VSUBS 0.032533f
C506 VTAIL.n364 VSUBS 0.014574f
C507 VTAIL.n365 VSUBS 0.013764f
C508 VTAIL.n366 VSUBS 0.025615f
C509 VTAIL.n367 VSUBS 0.025615f
C510 VTAIL.n368 VSUBS 0.013764f
C511 VTAIL.n369 VSUBS 0.014574f
C512 VTAIL.n370 VSUBS 0.032533f
C513 VTAIL.n371 VSUBS 0.032533f
C514 VTAIL.n372 VSUBS 0.014574f
C515 VTAIL.n373 VSUBS 0.013764f
C516 VTAIL.n374 VSUBS 0.025615f
C517 VTAIL.n375 VSUBS 0.025615f
C518 VTAIL.n376 VSUBS 0.013764f
C519 VTAIL.n377 VSUBS 0.014574f
C520 VTAIL.n378 VSUBS 0.032533f
C521 VTAIL.n379 VSUBS 0.032533f
C522 VTAIL.n380 VSUBS 0.032533f
C523 VTAIL.n381 VSUBS 0.014169f
C524 VTAIL.n382 VSUBS 0.013764f
C525 VTAIL.n383 VSUBS 0.025615f
C526 VTAIL.n384 VSUBS 0.025615f
C527 VTAIL.n385 VSUBS 0.013764f
C528 VTAIL.n386 VSUBS 0.014574f
C529 VTAIL.n387 VSUBS 0.032533f
C530 VTAIL.n388 VSUBS 0.032533f
C531 VTAIL.n389 VSUBS 0.014574f
C532 VTAIL.n390 VSUBS 0.013764f
C533 VTAIL.n391 VSUBS 0.025615f
C534 VTAIL.n392 VSUBS 0.025615f
C535 VTAIL.n393 VSUBS 0.013764f
C536 VTAIL.n394 VSUBS 0.014574f
C537 VTAIL.n395 VSUBS 0.032533f
C538 VTAIL.n396 VSUBS 0.078765f
C539 VTAIL.n397 VSUBS 0.014574f
C540 VTAIL.n398 VSUBS 0.013764f
C541 VTAIL.n399 VSUBS 0.059557f
C542 VTAIL.n400 VSUBS 0.039621f
C543 VTAIL.n401 VSUBS 0.309881f
C544 VTAIL.t15 VSUBS 0.245527f
C545 VTAIL.t8 VSUBS 0.245527f
C546 VTAIL.n402 VSUBS 1.78099f
C547 VTAIL.n403 VSUBS 1.08366f
C548 VTAIL.n404 VSUBS 0.028146f
C549 VTAIL.n405 VSUBS 0.025615f
C550 VTAIL.n406 VSUBS 0.013764f
C551 VTAIL.n407 VSUBS 0.032533f
C552 VTAIL.n408 VSUBS 0.014574f
C553 VTAIL.n409 VSUBS 0.025615f
C554 VTAIL.n410 VSUBS 0.013764f
C555 VTAIL.n411 VSUBS 0.032533f
C556 VTAIL.n412 VSUBS 0.014574f
C557 VTAIL.n413 VSUBS 0.025615f
C558 VTAIL.n414 VSUBS 0.014169f
C559 VTAIL.n415 VSUBS 0.032533f
C560 VTAIL.n416 VSUBS 0.013764f
C561 VTAIL.n417 VSUBS 0.014574f
C562 VTAIL.n418 VSUBS 0.025615f
C563 VTAIL.n419 VSUBS 0.013764f
C564 VTAIL.n420 VSUBS 0.032533f
C565 VTAIL.n421 VSUBS 0.014574f
C566 VTAIL.n422 VSUBS 0.025615f
C567 VTAIL.n423 VSUBS 0.013764f
C568 VTAIL.n424 VSUBS 0.0244f
C569 VTAIL.n425 VSUBS 0.024473f
C570 VTAIL.t14 VSUBS 0.070117f
C571 VTAIL.n426 VSUBS 0.203235f
C572 VTAIL.n427 VSUBS 1.27311f
C573 VTAIL.n428 VSUBS 0.013764f
C574 VTAIL.n429 VSUBS 0.014574f
C575 VTAIL.n430 VSUBS 0.032533f
C576 VTAIL.n431 VSUBS 0.032533f
C577 VTAIL.n432 VSUBS 0.014574f
C578 VTAIL.n433 VSUBS 0.013764f
C579 VTAIL.n434 VSUBS 0.025615f
C580 VTAIL.n435 VSUBS 0.025615f
C581 VTAIL.n436 VSUBS 0.013764f
C582 VTAIL.n437 VSUBS 0.014574f
C583 VTAIL.n438 VSUBS 0.032533f
C584 VTAIL.n439 VSUBS 0.032533f
C585 VTAIL.n440 VSUBS 0.014574f
C586 VTAIL.n441 VSUBS 0.013764f
C587 VTAIL.n442 VSUBS 0.025615f
C588 VTAIL.n443 VSUBS 0.025615f
C589 VTAIL.n444 VSUBS 0.013764f
C590 VTAIL.n445 VSUBS 0.014574f
C591 VTAIL.n446 VSUBS 0.032533f
C592 VTAIL.n447 VSUBS 0.032533f
C593 VTAIL.n448 VSUBS 0.032533f
C594 VTAIL.n449 VSUBS 0.014169f
C595 VTAIL.n450 VSUBS 0.013764f
C596 VTAIL.n451 VSUBS 0.025615f
C597 VTAIL.n452 VSUBS 0.025615f
C598 VTAIL.n453 VSUBS 0.013764f
C599 VTAIL.n454 VSUBS 0.014574f
C600 VTAIL.n455 VSUBS 0.032533f
C601 VTAIL.n456 VSUBS 0.032533f
C602 VTAIL.n457 VSUBS 0.014574f
C603 VTAIL.n458 VSUBS 0.013764f
C604 VTAIL.n459 VSUBS 0.025615f
C605 VTAIL.n460 VSUBS 0.025615f
C606 VTAIL.n461 VSUBS 0.013764f
C607 VTAIL.n462 VSUBS 0.014574f
C608 VTAIL.n463 VSUBS 0.032533f
C609 VTAIL.n464 VSUBS 0.078765f
C610 VTAIL.n465 VSUBS 0.014574f
C611 VTAIL.n466 VSUBS 0.013764f
C612 VTAIL.n467 VSUBS 0.059557f
C613 VTAIL.n468 VSUBS 0.039621f
C614 VTAIL.n469 VSUBS 1.73114f
C615 VTAIL.n470 VSUBS 0.028146f
C616 VTAIL.n471 VSUBS 0.025615f
C617 VTAIL.n472 VSUBS 0.013764f
C618 VTAIL.n473 VSUBS 0.032533f
C619 VTAIL.n474 VSUBS 0.014574f
C620 VTAIL.n475 VSUBS 0.025615f
C621 VTAIL.n476 VSUBS 0.013764f
C622 VTAIL.n477 VSUBS 0.032533f
C623 VTAIL.n478 VSUBS 0.014574f
C624 VTAIL.n479 VSUBS 0.025615f
C625 VTAIL.n480 VSUBS 0.014169f
C626 VTAIL.n481 VSUBS 0.032533f
C627 VTAIL.n482 VSUBS 0.014574f
C628 VTAIL.n483 VSUBS 0.025615f
C629 VTAIL.n484 VSUBS 0.013764f
C630 VTAIL.n485 VSUBS 0.032533f
C631 VTAIL.n486 VSUBS 0.014574f
C632 VTAIL.n487 VSUBS 0.025615f
C633 VTAIL.n488 VSUBS 0.013764f
C634 VTAIL.n489 VSUBS 0.0244f
C635 VTAIL.n490 VSUBS 0.024473f
C636 VTAIL.t2 VSUBS 0.070117f
C637 VTAIL.n491 VSUBS 0.203235f
C638 VTAIL.n492 VSUBS 1.27311f
C639 VTAIL.n493 VSUBS 0.013764f
C640 VTAIL.n494 VSUBS 0.014574f
C641 VTAIL.n495 VSUBS 0.032533f
C642 VTAIL.n496 VSUBS 0.032533f
C643 VTAIL.n497 VSUBS 0.014574f
C644 VTAIL.n498 VSUBS 0.013764f
C645 VTAIL.n499 VSUBS 0.025615f
C646 VTAIL.n500 VSUBS 0.025615f
C647 VTAIL.n501 VSUBS 0.013764f
C648 VTAIL.n502 VSUBS 0.014574f
C649 VTAIL.n503 VSUBS 0.032533f
C650 VTAIL.n504 VSUBS 0.032533f
C651 VTAIL.n505 VSUBS 0.014574f
C652 VTAIL.n506 VSUBS 0.013764f
C653 VTAIL.n507 VSUBS 0.025615f
C654 VTAIL.n508 VSUBS 0.025615f
C655 VTAIL.n509 VSUBS 0.013764f
C656 VTAIL.n510 VSUBS 0.013764f
C657 VTAIL.n511 VSUBS 0.014574f
C658 VTAIL.n512 VSUBS 0.032533f
C659 VTAIL.n513 VSUBS 0.032533f
C660 VTAIL.n514 VSUBS 0.032533f
C661 VTAIL.n515 VSUBS 0.014169f
C662 VTAIL.n516 VSUBS 0.013764f
C663 VTAIL.n517 VSUBS 0.025615f
C664 VTAIL.n518 VSUBS 0.025615f
C665 VTAIL.n519 VSUBS 0.013764f
C666 VTAIL.n520 VSUBS 0.014574f
C667 VTAIL.n521 VSUBS 0.032533f
C668 VTAIL.n522 VSUBS 0.032533f
C669 VTAIL.n523 VSUBS 0.014574f
C670 VTAIL.n524 VSUBS 0.013764f
C671 VTAIL.n525 VSUBS 0.025615f
C672 VTAIL.n526 VSUBS 0.025615f
C673 VTAIL.n527 VSUBS 0.013764f
C674 VTAIL.n528 VSUBS 0.014574f
C675 VTAIL.n529 VSUBS 0.032533f
C676 VTAIL.n530 VSUBS 0.078765f
C677 VTAIL.n531 VSUBS 0.014574f
C678 VTAIL.n532 VSUBS 0.013764f
C679 VTAIL.n533 VSUBS 0.059557f
C680 VTAIL.n534 VSUBS 0.039621f
C681 VTAIL.n535 VSUBS 1.72634f
C682 VP.t0 VSUBS 2.98972f
C683 VP.n0 VSUBS 1.15505f
C684 VP.n1 VSUBS 0.028528f
C685 VP.n2 VSUBS 0.023062f
C686 VP.n3 VSUBS 0.028528f
C687 VP.t3 VSUBS 2.98972f
C688 VP.n4 VSUBS 1.05098f
C689 VP.n5 VSUBS 0.028528f
C690 VP.n6 VSUBS 0.023062f
C691 VP.n7 VSUBS 0.028528f
C692 VP.t4 VSUBS 2.98972f
C693 VP.n8 VSUBS 1.05098f
C694 VP.n9 VSUBS 0.028528f
C695 VP.n10 VSUBS 0.023062f
C696 VP.n11 VSUBS 0.028528f
C697 VP.t7 VSUBS 2.98972f
C698 VP.n12 VSUBS 1.15505f
C699 VP.t5 VSUBS 2.98972f
C700 VP.n13 VSUBS 1.15505f
C701 VP.n14 VSUBS 0.028528f
C702 VP.n15 VSUBS 0.023062f
C703 VP.n16 VSUBS 0.028528f
C704 VP.t6 VSUBS 2.98972f
C705 VP.n17 VSUBS 1.05098f
C706 VP.n18 VSUBS 0.028528f
C707 VP.n19 VSUBS 0.023062f
C708 VP.n20 VSUBS 0.028528f
C709 VP.t1 VSUBS 2.98972f
C710 VP.n21 VSUBS 1.14446f
C711 VP.t2 VSUBS 3.31591f
C712 VP.n22 VSUBS 1.09462f
C713 VP.n23 VSUBS 0.331672f
C714 VP.n24 VSUBS 0.040044f
C715 VP.n25 VSUBS 0.053169f
C716 VP.n26 VSUBS 0.056699f
C717 VP.n27 VSUBS 0.028528f
C718 VP.n28 VSUBS 0.028528f
C719 VP.n29 VSUBS 0.028528f
C720 VP.n30 VSUBS 0.056699f
C721 VP.n31 VSUBS 0.053169f
C722 VP.n32 VSUBS 0.040044f
C723 VP.n33 VSUBS 0.028528f
C724 VP.n34 VSUBS 0.028528f
C725 VP.n35 VSUBS 0.040044f
C726 VP.n36 VSUBS 0.053169f
C727 VP.n37 VSUBS 0.056699f
C728 VP.n38 VSUBS 0.028528f
C729 VP.n39 VSUBS 0.028528f
C730 VP.n40 VSUBS 0.028528f
C731 VP.n41 VSUBS 0.056699f
C732 VP.n42 VSUBS 0.053169f
C733 VP.n43 VSUBS 0.040044f
C734 VP.n44 VSUBS 0.046044f
C735 VP.n45 VSUBS 1.79445f
C736 VP.n46 VSUBS 1.81355f
C737 VP.n47 VSUBS 0.046044f
C738 VP.n48 VSUBS 0.040044f
C739 VP.n49 VSUBS 0.053169f
C740 VP.n50 VSUBS 0.056699f
C741 VP.n51 VSUBS 0.028528f
C742 VP.n52 VSUBS 0.028528f
C743 VP.n53 VSUBS 0.028528f
C744 VP.n54 VSUBS 0.056699f
C745 VP.n55 VSUBS 0.053169f
C746 VP.n56 VSUBS 0.040044f
C747 VP.n57 VSUBS 0.028528f
C748 VP.n58 VSUBS 0.028528f
C749 VP.n59 VSUBS 0.040044f
C750 VP.n60 VSUBS 0.053169f
C751 VP.n61 VSUBS 0.056699f
C752 VP.n62 VSUBS 0.028528f
C753 VP.n63 VSUBS 0.028528f
C754 VP.n64 VSUBS 0.028528f
C755 VP.n65 VSUBS 0.056699f
C756 VP.n66 VSUBS 0.053169f
C757 VP.n67 VSUBS 0.040044f
C758 VP.n68 VSUBS 0.028528f
C759 VP.n69 VSUBS 0.028528f
C760 VP.n70 VSUBS 0.040044f
C761 VP.n71 VSUBS 0.053169f
C762 VP.n72 VSUBS 0.056699f
C763 VP.n73 VSUBS 0.028528f
C764 VP.n74 VSUBS 0.028528f
C765 VP.n75 VSUBS 0.028528f
C766 VP.n76 VSUBS 0.056699f
C767 VP.n77 VSUBS 0.053169f
C768 VP.n78 VSUBS 0.040044f
C769 VP.n79 VSUBS 0.046044f
C770 VP.n80 VSUBS 0.070055f
C771 B.n0 VSUBS 0.006462f
C772 B.n1 VSUBS 0.006462f
C773 B.n2 VSUBS 0.009557f
C774 B.n3 VSUBS 0.007324f
C775 B.n4 VSUBS 0.007324f
C776 B.n5 VSUBS 0.007324f
C777 B.n6 VSUBS 0.007324f
C778 B.n7 VSUBS 0.007324f
C779 B.n8 VSUBS 0.007324f
C780 B.n9 VSUBS 0.007324f
C781 B.n10 VSUBS 0.007324f
C782 B.n11 VSUBS 0.007324f
C783 B.n12 VSUBS 0.007324f
C784 B.n13 VSUBS 0.007324f
C785 B.n14 VSUBS 0.007324f
C786 B.n15 VSUBS 0.007324f
C787 B.n16 VSUBS 0.007324f
C788 B.n17 VSUBS 0.007324f
C789 B.n18 VSUBS 0.007324f
C790 B.n19 VSUBS 0.007324f
C791 B.n20 VSUBS 0.007324f
C792 B.n21 VSUBS 0.007324f
C793 B.n22 VSUBS 0.007324f
C794 B.n23 VSUBS 0.007324f
C795 B.n24 VSUBS 0.007324f
C796 B.n25 VSUBS 0.007324f
C797 B.n26 VSUBS 0.007324f
C798 B.n27 VSUBS 0.007324f
C799 B.n28 VSUBS 0.007324f
C800 B.n29 VSUBS 0.007324f
C801 B.n30 VSUBS 0.007324f
C802 B.n31 VSUBS 0.015931f
C803 B.n32 VSUBS 0.007324f
C804 B.n33 VSUBS 0.007324f
C805 B.n34 VSUBS 0.007324f
C806 B.n35 VSUBS 0.007324f
C807 B.n36 VSUBS 0.007324f
C808 B.n37 VSUBS 0.007324f
C809 B.n38 VSUBS 0.007324f
C810 B.n39 VSUBS 0.007324f
C811 B.n40 VSUBS 0.007324f
C812 B.n41 VSUBS 0.007324f
C813 B.n42 VSUBS 0.007324f
C814 B.n43 VSUBS 0.007324f
C815 B.n44 VSUBS 0.007324f
C816 B.n45 VSUBS 0.007324f
C817 B.n46 VSUBS 0.007324f
C818 B.n47 VSUBS 0.007324f
C819 B.n48 VSUBS 0.007324f
C820 B.n49 VSUBS 0.007324f
C821 B.n50 VSUBS 0.007324f
C822 B.n51 VSUBS 0.007324f
C823 B.n52 VSUBS 0.006893f
C824 B.n53 VSUBS 0.007324f
C825 B.t1 VSUBS 0.223906f
C826 B.t2 VSUBS 0.263071f
C827 B.t0 VSUBS 1.85501f
C828 B.n54 VSUBS 0.419354f
C829 B.n55 VSUBS 0.267745f
C830 B.n56 VSUBS 0.016968f
C831 B.n57 VSUBS 0.007324f
C832 B.n58 VSUBS 0.007324f
C833 B.n59 VSUBS 0.007324f
C834 B.n60 VSUBS 0.007324f
C835 B.t4 VSUBS 0.223909f
C836 B.t5 VSUBS 0.263074f
C837 B.t3 VSUBS 1.85501f
C838 B.n61 VSUBS 0.419351f
C839 B.n62 VSUBS 0.267742f
C840 B.n63 VSUBS 0.007324f
C841 B.n64 VSUBS 0.007324f
C842 B.n65 VSUBS 0.007324f
C843 B.n66 VSUBS 0.007324f
C844 B.n67 VSUBS 0.007324f
C845 B.n68 VSUBS 0.007324f
C846 B.n69 VSUBS 0.007324f
C847 B.n70 VSUBS 0.007324f
C848 B.n71 VSUBS 0.007324f
C849 B.n72 VSUBS 0.007324f
C850 B.n73 VSUBS 0.007324f
C851 B.n74 VSUBS 0.007324f
C852 B.n75 VSUBS 0.007324f
C853 B.n76 VSUBS 0.007324f
C854 B.n77 VSUBS 0.007324f
C855 B.n78 VSUBS 0.007324f
C856 B.n79 VSUBS 0.007324f
C857 B.n80 VSUBS 0.007324f
C858 B.n81 VSUBS 0.007324f
C859 B.n82 VSUBS 0.007324f
C860 B.n83 VSUBS 0.017241f
C861 B.n84 VSUBS 0.007324f
C862 B.n85 VSUBS 0.007324f
C863 B.n86 VSUBS 0.007324f
C864 B.n87 VSUBS 0.007324f
C865 B.n88 VSUBS 0.007324f
C866 B.n89 VSUBS 0.007324f
C867 B.n90 VSUBS 0.007324f
C868 B.n91 VSUBS 0.007324f
C869 B.n92 VSUBS 0.007324f
C870 B.n93 VSUBS 0.007324f
C871 B.n94 VSUBS 0.007324f
C872 B.n95 VSUBS 0.007324f
C873 B.n96 VSUBS 0.007324f
C874 B.n97 VSUBS 0.007324f
C875 B.n98 VSUBS 0.007324f
C876 B.n99 VSUBS 0.007324f
C877 B.n100 VSUBS 0.007324f
C878 B.n101 VSUBS 0.007324f
C879 B.n102 VSUBS 0.007324f
C880 B.n103 VSUBS 0.007324f
C881 B.n104 VSUBS 0.007324f
C882 B.n105 VSUBS 0.007324f
C883 B.n106 VSUBS 0.007324f
C884 B.n107 VSUBS 0.007324f
C885 B.n108 VSUBS 0.007324f
C886 B.n109 VSUBS 0.007324f
C887 B.n110 VSUBS 0.007324f
C888 B.n111 VSUBS 0.007324f
C889 B.n112 VSUBS 0.007324f
C890 B.n113 VSUBS 0.007324f
C891 B.n114 VSUBS 0.007324f
C892 B.n115 VSUBS 0.007324f
C893 B.n116 VSUBS 0.007324f
C894 B.n117 VSUBS 0.007324f
C895 B.n118 VSUBS 0.007324f
C896 B.n119 VSUBS 0.007324f
C897 B.n120 VSUBS 0.007324f
C898 B.n121 VSUBS 0.007324f
C899 B.n122 VSUBS 0.007324f
C900 B.n123 VSUBS 0.007324f
C901 B.n124 VSUBS 0.007324f
C902 B.n125 VSUBS 0.007324f
C903 B.n126 VSUBS 0.007324f
C904 B.n127 VSUBS 0.007324f
C905 B.n128 VSUBS 0.007324f
C906 B.n129 VSUBS 0.007324f
C907 B.n130 VSUBS 0.007324f
C908 B.n131 VSUBS 0.007324f
C909 B.n132 VSUBS 0.007324f
C910 B.n133 VSUBS 0.007324f
C911 B.n134 VSUBS 0.007324f
C912 B.n135 VSUBS 0.007324f
C913 B.n136 VSUBS 0.007324f
C914 B.n137 VSUBS 0.007324f
C915 B.n138 VSUBS 0.007324f
C916 B.n139 VSUBS 0.007324f
C917 B.n140 VSUBS 0.007324f
C918 B.n141 VSUBS 0.007324f
C919 B.n142 VSUBS 0.007324f
C920 B.n143 VSUBS 0.016841f
C921 B.n144 VSUBS 0.007324f
C922 B.n145 VSUBS 0.007324f
C923 B.n146 VSUBS 0.007324f
C924 B.n147 VSUBS 0.007324f
C925 B.n148 VSUBS 0.007324f
C926 B.n149 VSUBS 0.007324f
C927 B.n150 VSUBS 0.007324f
C928 B.n151 VSUBS 0.007324f
C929 B.n152 VSUBS 0.007324f
C930 B.n153 VSUBS 0.007324f
C931 B.n154 VSUBS 0.007324f
C932 B.n155 VSUBS 0.007324f
C933 B.n156 VSUBS 0.007324f
C934 B.n157 VSUBS 0.007324f
C935 B.n158 VSUBS 0.007324f
C936 B.n159 VSUBS 0.007324f
C937 B.n160 VSUBS 0.007324f
C938 B.n161 VSUBS 0.007324f
C939 B.n162 VSUBS 0.007324f
C940 B.n163 VSUBS 0.007324f
C941 B.n164 VSUBS 0.007324f
C942 B.t8 VSUBS 0.223909f
C943 B.t7 VSUBS 0.263074f
C944 B.t6 VSUBS 1.85501f
C945 B.n165 VSUBS 0.419351f
C946 B.n166 VSUBS 0.267742f
C947 B.n167 VSUBS 0.007324f
C948 B.n168 VSUBS 0.007324f
C949 B.n169 VSUBS 0.007324f
C950 B.n170 VSUBS 0.007324f
C951 B.n171 VSUBS 0.004093f
C952 B.n172 VSUBS 0.007324f
C953 B.n173 VSUBS 0.007324f
C954 B.n174 VSUBS 0.007324f
C955 B.n175 VSUBS 0.007324f
C956 B.n176 VSUBS 0.007324f
C957 B.n177 VSUBS 0.007324f
C958 B.n178 VSUBS 0.007324f
C959 B.n179 VSUBS 0.007324f
C960 B.n180 VSUBS 0.007324f
C961 B.n181 VSUBS 0.007324f
C962 B.n182 VSUBS 0.007324f
C963 B.n183 VSUBS 0.007324f
C964 B.n184 VSUBS 0.007324f
C965 B.n185 VSUBS 0.007324f
C966 B.n186 VSUBS 0.007324f
C967 B.n187 VSUBS 0.007324f
C968 B.n188 VSUBS 0.007324f
C969 B.n189 VSUBS 0.007324f
C970 B.n190 VSUBS 0.007324f
C971 B.n191 VSUBS 0.007324f
C972 B.n192 VSUBS 0.017241f
C973 B.n193 VSUBS 0.007324f
C974 B.n194 VSUBS 0.007324f
C975 B.n195 VSUBS 0.007324f
C976 B.n196 VSUBS 0.007324f
C977 B.n197 VSUBS 0.007324f
C978 B.n198 VSUBS 0.007324f
C979 B.n199 VSUBS 0.007324f
C980 B.n200 VSUBS 0.007324f
C981 B.n201 VSUBS 0.007324f
C982 B.n202 VSUBS 0.007324f
C983 B.n203 VSUBS 0.007324f
C984 B.n204 VSUBS 0.007324f
C985 B.n205 VSUBS 0.007324f
C986 B.n206 VSUBS 0.007324f
C987 B.n207 VSUBS 0.007324f
C988 B.n208 VSUBS 0.007324f
C989 B.n209 VSUBS 0.007324f
C990 B.n210 VSUBS 0.007324f
C991 B.n211 VSUBS 0.007324f
C992 B.n212 VSUBS 0.007324f
C993 B.n213 VSUBS 0.007324f
C994 B.n214 VSUBS 0.007324f
C995 B.n215 VSUBS 0.007324f
C996 B.n216 VSUBS 0.007324f
C997 B.n217 VSUBS 0.007324f
C998 B.n218 VSUBS 0.007324f
C999 B.n219 VSUBS 0.007324f
C1000 B.n220 VSUBS 0.007324f
C1001 B.n221 VSUBS 0.007324f
C1002 B.n222 VSUBS 0.007324f
C1003 B.n223 VSUBS 0.007324f
C1004 B.n224 VSUBS 0.007324f
C1005 B.n225 VSUBS 0.007324f
C1006 B.n226 VSUBS 0.007324f
C1007 B.n227 VSUBS 0.007324f
C1008 B.n228 VSUBS 0.007324f
C1009 B.n229 VSUBS 0.007324f
C1010 B.n230 VSUBS 0.007324f
C1011 B.n231 VSUBS 0.007324f
C1012 B.n232 VSUBS 0.007324f
C1013 B.n233 VSUBS 0.007324f
C1014 B.n234 VSUBS 0.007324f
C1015 B.n235 VSUBS 0.007324f
C1016 B.n236 VSUBS 0.007324f
C1017 B.n237 VSUBS 0.007324f
C1018 B.n238 VSUBS 0.007324f
C1019 B.n239 VSUBS 0.007324f
C1020 B.n240 VSUBS 0.007324f
C1021 B.n241 VSUBS 0.007324f
C1022 B.n242 VSUBS 0.007324f
C1023 B.n243 VSUBS 0.007324f
C1024 B.n244 VSUBS 0.007324f
C1025 B.n245 VSUBS 0.007324f
C1026 B.n246 VSUBS 0.007324f
C1027 B.n247 VSUBS 0.007324f
C1028 B.n248 VSUBS 0.007324f
C1029 B.n249 VSUBS 0.007324f
C1030 B.n250 VSUBS 0.007324f
C1031 B.n251 VSUBS 0.007324f
C1032 B.n252 VSUBS 0.007324f
C1033 B.n253 VSUBS 0.007324f
C1034 B.n254 VSUBS 0.007324f
C1035 B.n255 VSUBS 0.007324f
C1036 B.n256 VSUBS 0.007324f
C1037 B.n257 VSUBS 0.007324f
C1038 B.n258 VSUBS 0.007324f
C1039 B.n259 VSUBS 0.007324f
C1040 B.n260 VSUBS 0.007324f
C1041 B.n261 VSUBS 0.007324f
C1042 B.n262 VSUBS 0.007324f
C1043 B.n263 VSUBS 0.007324f
C1044 B.n264 VSUBS 0.007324f
C1045 B.n265 VSUBS 0.007324f
C1046 B.n266 VSUBS 0.007324f
C1047 B.n267 VSUBS 0.007324f
C1048 B.n268 VSUBS 0.007324f
C1049 B.n269 VSUBS 0.007324f
C1050 B.n270 VSUBS 0.007324f
C1051 B.n271 VSUBS 0.007324f
C1052 B.n272 VSUBS 0.007324f
C1053 B.n273 VSUBS 0.007324f
C1054 B.n274 VSUBS 0.007324f
C1055 B.n275 VSUBS 0.007324f
C1056 B.n276 VSUBS 0.007324f
C1057 B.n277 VSUBS 0.007324f
C1058 B.n278 VSUBS 0.007324f
C1059 B.n279 VSUBS 0.007324f
C1060 B.n280 VSUBS 0.007324f
C1061 B.n281 VSUBS 0.007324f
C1062 B.n282 VSUBS 0.007324f
C1063 B.n283 VSUBS 0.007324f
C1064 B.n284 VSUBS 0.007324f
C1065 B.n285 VSUBS 0.007324f
C1066 B.n286 VSUBS 0.007324f
C1067 B.n287 VSUBS 0.007324f
C1068 B.n288 VSUBS 0.007324f
C1069 B.n289 VSUBS 0.007324f
C1070 B.n290 VSUBS 0.007324f
C1071 B.n291 VSUBS 0.007324f
C1072 B.n292 VSUBS 0.007324f
C1073 B.n293 VSUBS 0.007324f
C1074 B.n294 VSUBS 0.007324f
C1075 B.n295 VSUBS 0.007324f
C1076 B.n296 VSUBS 0.007324f
C1077 B.n297 VSUBS 0.007324f
C1078 B.n298 VSUBS 0.007324f
C1079 B.n299 VSUBS 0.007324f
C1080 B.n300 VSUBS 0.007324f
C1081 B.n301 VSUBS 0.007324f
C1082 B.n302 VSUBS 0.007324f
C1083 B.n303 VSUBS 0.007324f
C1084 B.n304 VSUBS 0.007324f
C1085 B.n305 VSUBS 0.007324f
C1086 B.n306 VSUBS 0.007324f
C1087 B.n307 VSUBS 0.015931f
C1088 B.n308 VSUBS 0.015931f
C1089 B.n309 VSUBS 0.017241f
C1090 B.n310 VSUBS 0.007324f
C1091 B.n311 VSUBS 0.007324f
C1092 B.n312 VSUBS 0.007324f
C1093 B.n313 VSUBS 0.007324f
C1094 B.n314 VSUBS 0.007324f
C1095 B.n315 VSUBS 0.007324f
C1096 B.n316 VSUBS 0.007324f
C1097 B.n317 VSUBS 0.007324f
C1098 B.n318 VSUBS 0.007324f
C1099 B.n319 VSUBS 0.007324f
C1100 B.n320 VSUBS 0.007324f
C1101 B.n321 VSUBS 0.007324f
C1102 B.n322 VSUBS 0.007324f
C1103 B.n323 VSUBS 0.007324f
C1104 B.n324 VSUBS 0.007324f
C1105 B.n325 VSUBS 0.007324f
C1106 B.n326 VSUBS 0.007324f
C1107 B.n327 VSUBS 0.007324f
C1108 B.n328 VSUBS 0.007324f
C1109 B.n329 VSUBS 0.007324f
C1110 B.n330 VSUBS 0.007324f
C1111 B.n331 VSUBS 0.007324f
C1112 B.n332 VSUBS 0.007324f
C1113 B.n333 VSUBS 0.007324f
C1114 B.n334 VSUBS 0.007324f
C1115 B.n335 VSUBS 0.007324f
C1116 B.n336 VSUBS 0.007324f
C1117 B.n337 VSUBS 0.007324f
C1118 B.n338 VSUBS 0.007324f
C1119 B.n339 VSUBS 0.007324f
C1120 B.n340 VSUBS 0.007324f
C1121 B.n341 VSUBS 0.007324f
C1122 B.n342 VSUBS 0.007324f
C1123 B.n343 VSUBS 0.007324f
C1124 B.n344 VSUBS 0.007324f
C1125 B.n345 VSUBS 0.007324f
C1126 B.n346 VSUBS 0.007324f
C1127 B.n347 VSUBS 0.007324f
C1128 B.n348 VSUBS 0.007324f
C1129 B.n349 VSUBS 0.007324f
C1130 B.n350 VSUBS 0.007324f
C1131 B.n351 VSUBS 0.007324f
C1132 B.n352 VSUBS 0.007324f
C1133 B.n353 VSUBS 0.007324f
C1134 B.n354 VSUBS 0.007324f
C1135 B.n355 VSUBS 0.007324f
C1136 B.n356 VSUBS 0.007324f
C1137 B.n357 VSUBS 0.007324f
C1138 B.n358 VSUBS 0.007324f
C1139 B.n359 VSUBS 0.007324f
C1140 B.n360 VSUBS 0.007324f
C1141 B.n361 VSUBS 0.007324f
C1142 B.n362 VSUBS 0.007324f
C1143 B.n363 VSUBS 0.007324f
C1144 B.n364 VSUBS 0.007324f
C1145 B.n365 VSUBS 0.007324f
C1146 B.n366 VSUBS 0.007324f
C1147 B.n367 VSUBS 0.007324f
C1148 B.n368 VSUBS 0.007324f
C1149 B.n369 VSUBS 0.007324f
C1150 B.t11 VSUBS 0.223906f
C1151 B.t10 VSUBS 0.263071f
C1152 B.t9 VSUBS 1.85501f
C1153 B.n370 VSUBS 0.419354f
C1154 B.n371 VSUBS 0.267745f
C1155 B.n372 VSUBS 0.016968f
C1156 B.n373 VSUBS 0.006893f
C1157 B.n374 VSUBS 0.007324f
C1158 B.n375 VSUBS 0.007324f
C1159 B.n376 VSUBS 0.007324f
C1160 B.n377 VSUBS 0.007324f
C1161 B.n378 VSUBS 0.007324f
C1162 B.n379 VSUBS 0.007324f
C1163 B.n380 VSUBS 0.007324f
C1164 B.n381 VSUBS 0.007324f
C1165 B.n382 VSUBS 0.007324f
C1166 B.n383 VSUBS 0.007324f
C1167 B.n384 VSUBS 0.007324f
C1168 B.n385 VSUBS 0.007324f
C1169 B.n386 VSUBS 0.007324f
C1170 B.n387 VSUBS 0.007324f
C1171 B.n388 VSUBS 0.007324f
C1172 B.n389 VSUBS 0.004093f
C1173 B.n390 VSUBS 0.016968f
C1174 B.n391 VSUBS 0.006893f
C1175 B.n392 VSUBS 0.007324f
C1176 B.n393 VSUBS 0.007324f
C1177 B.n394 VSUBS 0.007324f
C1178 B.n395 VSUBS 0.007324f
C1179 B.n396 VSUBS 0.007324f
C1180 B.n397 VSUBS 0.007324f
C1181 B.n398 VSUBS 0.007324f
C1182 B.n399 VSUBS 0.007324f
C1183 B.n400 VSUBS 0.007324f
C1184 B.n401 VSUBS 0.007324f
C1185 B.n402 VSUBS 0.007324f
C1186 B.n403 VSUBS 0.007324f
C1187 B.n404 VSUBS 0.007324f
C1188 B.n405 VSUBS 0.007324f
C1189 B.n406 VSUBS 0.007324f
C1190 B.n407 VSUBS 0.007324f
C1191 B.n408 VSUBS 0.007324f
C1192 B.n409 VSUBS 0.007324f
C1193 B.n410 VSUBS 0.007324f
C1194 B.n411 VSUBS 0.007324f
C1195 B.n412 VSUBS 0.007324f
C1196 B.n413 VSUBS 0.007324f
C1197 B.n414 VSUBS 0.007324f
C1198 B.n415 VSUBS 0.007324f
C1199 B.n416 VSUBS 0.007324f
C1200 B.n417 VSUBS 0.007324f
C1201 B.n418 VSUBS 0.007324f
C1202 B.n419 VSUBS 0.007324f
C1203 B.n420 VSUBS 0.007324f
C1204 B.n421 VSUBS 0.007324f
C1205 B.n422 VSUBS 0.007324f
C1206 B.n423 VSUBS 0.007324f
C1207 B.n424 VSUBS 0.007324f
C1208 B.n425 VSUBS 0.007324f
C1209 B.n426 VSUBS 0.007324f
C1210 B.n427 VSUBS 0.007324f
C1211 B.n428 VSUBS 0.007324f
C1212 B.n429 VSUBS 0.007324f
C1213 B.n430 VSUBS 0.007324f
C1214 B.n431 VSUBS 0.007324f
C1215 B.n432 VSUBS 0.007324f
C1216 B.n433 VSUBS 0.007324f
C1217 B.n434 VSUBS 0.007324f
C1218 B.n435 VSUBS 0.007324f
C1219 B.n436 VSUBS 0.007324f
C1220 B.n437 VSUBS 0.007324f
C1221 B.n438 VSUBS 0.007324f
C1222 B.n439 VSUBS 0.007324f
C1223 B.n440 VSUBS 0.007324f
C1224 B.n441 VSUBS 0.007324f
C1225 B.n442 VSUBS 0.007324f
C1226 B.n443 VSUBS 0.007324f
C1227 B.n444 VSUBS 0.007324f
C1228 B.n445 VSUBS 0.007324f
C1229 B.n446 VSUBS 0.007324f
C1230 B.n447 VSUBS 0.007324f
C1231 B.n448 VSUBS 0.007324f
C1232 B.n449 VSUBS 0.007324f
C1233 B.n450 VSUBS 0.007324f
C1234 B.n451 VSUBS 0.007324f
C1235 B.n452 VSUBS 0.016331f
C1236 B.n453 VSUBS 0.017241f
C1237 B.n454 VSUBS 0.015931f
C1238 B.n455 VSUBS 0.007324f
C1239 B.n456 VSUBS 0.007324f
C1240 B.n457 VSUBS 0.007324f
C1241 B.n458 VSUBS 0.007324f
C1242 B.n459 VSUBS 0.007324f
C1243 B.n460 VSUBS 0.007324f
C1244 B.n461 VSUBS 0.007324f
C1245 B.n462 VSUBS 0.007324f
C1246 B.n463 VSUBS 0.007324f
C1247 B.n464 VSUBS 0.007324f
C1248 B.n465 VSUBS 0.007324f
C1249 B.n466 VSUBS 0.007324f
C1250 B.n467 VSUBS 0.007324f
C1251 B.n468 VSUBS 0.007324f
C1252 B.n469 VSUBS 0.007324f
C1253 B.n470 VSUBS 0.007324f
C1254 B.n471 VSUBS 0.007324f
C1255 B.n472 VSUBS 0.007324f
C1256 B.n473 VSUBS 0.007324f
C1257 B.n474 VSUBS 0.007324f
C1258 B.n475 VSUBS 0.007324f
C1259 B.n476 VSUBS 0.007324f
C1260 B.n477 VSUBS 0.007324f
C1261 B.n478 VSUBS 0.007324f
C1262 B.n479 VSUBS 0.007324f
C1263 B.n480 VSUBS 0.007324f
C1264 B.n481 VSUBS 0.007324f
C1265 B.n482 VSUBS 0.007324f
C1266 B.n483 VSUBS 0.007324f
C1267 B.n484 VSUBS 0.007324f
C1268 B.n485 VSUBS 0.007324f
C1269 B.n486 VSUBS 0.007324f
C1270 B.n487 VSUBS 0.007324f
C1271 B.n488 VSUBS 0.007324f
C1272 B.n489 VSUBS 0.007324f
C1273 B.n490 VSUBS 0.007324f
C1274 B.n491 VSUBS 0.007324f
C1275 B.n492 VSUBS 0.007324f
C1276 B.n493 VSUBS 0.007324f
C1277 B.n494 VSUBS 0.007324f
C1278 B.n495 VSUBS 0.007324f
C1279 B.n496 VSUBS 0.007324f
C1280 B.n497 VSUBS 0.007324f
C1281 B.n498 VSUBS 0.007324f
C1282 B.n499 VSUBS 0.007324f
C1283 B.n500 VSUBS 0.007324f
C1284 B.n501 VSUBS 0.007324f
C1285 B.n502 VSUBS 0.007324f
C1286 B.n503 VSUBS 0.007324f
C1287 B.n504 VSUBS 0.007324f
C1288 B.n505 VSUBS 0.007324f
C1289 B.n506 VSUBS 0.007324f
C1290 B.n507 VSUBS 0.007324f
C1291 B.n508 VSUBS 0.007324f
C1292 B.n509 VSUBS 0.007324f
C1293 B.n510 VSUBS 0.007324f
C1294 B.n511 VSUBS 0.007324f
C1295 B.n512 VSUBS 0.007324f
C1296 B.n513 VSUBS 0.007324f
C1297 B.n514 VSUBS 0.007324f
C1298 B.n515 VSUBS 0.007324f
C1299 B.n516 VSUBS 0.007324f
C1300 B.n517 VSUBS 0.007324f
C1301 B.n518 VSUBS 0.007324f
C1302 B.n519 VSUBS 0.007324f
C1303 B.n520 VSUBS 0.007324f
C1304 B.n521 VSUBS 0.007324f
C1305 B.n522 VSUBS 0.007324f
C1306 B.n523 VSUBS 0.007324f
C1307 B.n524 VSUBS 0.007324f
C1308 B.n525 VSUBS 0.007324f
C1309 B.n526 VSUBS 0.007324f
C1310 B.n527 VSUBS 0.007324f
C1311 B.n528 VSUBS 0.007324f
C1312 B.n529 VSUBS 0.007324f
C1313 B.n530 VSUBS 0.007324f
C1314 B.n531 VSUBS 0.007324f
C1315 B.n532 VSUBS 0.007324f
C1316 B.n533 VSUBS 0.007324f
C1317 B.n534 VSUBS 0.007324f
C1318 B.n535 VSUBS 0.007324f
C1319 B.n536 VSUBS 0.007324f
C1320 B.n537 VSUBS 0.007324f
C1321 B.n538 VSUBS 0.007324f
C1322 B.n539 VSUBS 0.007324f
C1323 B.n540 VSUBS 0.007324f
C1324 B.n541 VSUBS 0.007324f
C1325 B.n542 VSUBS 0.007324f
C1326 B.n543 VSUBS 0.007324f
C1327 B.n544 VSUBS 0.007324f
C1328 B.n545 VSUBS 0.007324f
C1329 B.n546 VSUBS 0.007324f
C1330 B.n547 VSUBS 0.007324f
C1331 B.n548 VSUBS 0.007324f
C1332 B.n549 VSUBS 0.007324f
C1333 B.n550 VSUBS 0.007324f
C1334 B.n551 VSUBS 0.007324f
C1335 B.n552 VSUBS 0.007324f
C1336 B.n553 VSUBS 0.007324f
C1337 B.n554 VSUBS 0.007324f
C1338 B.n555 VSUBS 0.007324f
C1339 B.n556 VSUBS 0.007324f
C1340 B.n557 VSUBS 0.007324f
C1341 B.n558 VSUBS 0.007324f
C1342 B.n559 VSUBS 0.007324f
C1343 B.n560 VSUBS 0.007324f
C1344 B.n561 VSUBS 0.007324f
C1345 B.n562 VSUBS 0.007324f
C1346 B.n563 VSUBS 0.007324f
C1347 B.n564 VSUBS 0.007324f
C1348 B.n565 VSUBS 0.007324f
C1349 B.n566 VSUBS 0.007324f
C1350 B.n567 VSUBS 0.007324f
C1351 B.n568 VSUBS 0.007324f
C1352 B.n569 VSUBS 0.007324f
C1353 B.n570 VSUBS 0.007324f
C1354 B.n571 VSUBS 0.007324f
C1355 B.n572 VSUBS 0.007324f
C1356 B.n573 VSUBS 0.007324f
C1357 B.n574 VSUBS 0.007324f
C1358 B.n575 VSUBS 0.007324f
C1359 B.n576 VSUBS 0.007324f
C1360 B.n577 VSUBS 0.007324f
C1361 B.n578 VSUBS 0.007324f
C1362 B.n579 VSUBS 0.007324f
C1363 B.n580 VSUBS 0.007324f
C1364 B.n581 VSUBS 0.007324f
C1365 B.n582 VSUBS 0.007324f
C1366 B.n583 VSUBS 0.007324f
C1367 B.n584 VSUBS 0.007324f
C1368 B.n585 VSUBS 0.007324f
C1369 B.n586 VSUBS 0.007324f
C1370 B.n587 VSUBS 0.007324f
C1371 B.n588 VSUBS 0.007324f
C1372 B.n589 VSUBS 0.007324f
C1373 B.n590 VSUBS 0.007324f
C1374 B.n591 VSUBS 0.007324f
C1375 B.n592 VSUBS 0.007324f
C1376 B.n593 VSUBS 0.007324f
C1377 B.n594 VSUBS 0.007324f
C1378 B.n595 VSUBS 0.007324f
C1379 B.n596 VSUBS 0.007324f
C1380 B.n597 VSUBS 0.007324f
C1381 B.n598 VSUBS 0.007324f
C1382 B.n599 VSUBS 0.007324f
C1383 B.n600 VSUBS 0.007324f
C1384 B.n601 VSUBS 0.007324f
C1385 B.n602 VSUBS 0.007324f
C1386 B.n603 VSUBS 0.007324f
C1387 B.n604 VSUBS 0.007324f
C1388 B.n605 VSUBS 0.007324f
C1389 B.n606 VSUBS 0.007324f
C1390 B.n607 VSUBS 0.007324f
C1391 B.n608 VSUBS 0.007324f
C1392 B.n609 VSUBS 0.007324f
C1393 B.n610 VSUBS 0.007324f
C1394 B.n611 VSUBS 0.007324f
C1395 B.n612 VSUBS 0.007324f
C1396 B.n613 VSUBS 0.007324f
C1397 B.n614 VSUBS 0.007324f
C1398 B.n615 VSUBS 0.007324f
C1399 B.n616 VSUBS 0.007324f
C1400 B.n617 VSUBS 0.007324f
C1401 B.n618 VSUBS 0.007324f
C1402 B.n619 VSUBS 0.007324f
C1403 B.n620 VSUBS 0.007324f
C1404 B.n621 VSUBS 0.007324f
C1405 B.n622 VSUBS 0.007324f
C1406 B.n623 VSUBS 0.007324f
C1407 B.n624 VSUBS 0.007324f
C1408 B.n625 VSUBS 0.007324f
C1409 B.n626 VSUBS 0.007324f
C1410 B.n627 VSUBS 0.007324f
C1411 B.n628 VSUBS 0.007324f
C1412 B.n629 VSUBS 0.007324f
C1413 B.n630 VSUBS 0.007324f
C1414 B.n631 VSUBS 0.007324f
C1415 B.n632 VSUBS 0.015931f
C1416 B.n633 VSUBS 0.015931f
C1417 B.n634 VSUBS 0.017241f
C1418 B.n635 VSUBS 0.007324f
C1419 B.n636 VSUBS 0.007324f
C1420 B.n637 VSUBS 0.007324f
C1421 B.n638 VSUBS 0.007324f
C1422 B.n639 VSUBS 0.007324f
C1423 B.n640 VSUBS 0.007324f
C1424 B.n641 VSUBS 0.007324f
C1425 B.n642 VSUBS 0.007324f
C1426 B.n643 VSUBS 0.007324f
C1427 B.n644 VSUBS 0.007324f
C1428 B.n645 VSUBS 0.007324f
C1429 B.n646 VSUBS 0.007324f
C1430 B.n647 VSUBS 0.007324f
C1431 B.n648 VSUBS 0.007324f
C1432 B.n649 VSUBS 0.007324f
C1433 B.n650 VSUBS 0.007324f
C1434 B.n651 VSUBS 0.007324f
C1435 B.n652 VSUBS 0.007324f
C1436 B.n653 VSUBS 0.007324f
C1437 B.n654 VSUBS 0.007324f
C1438 B.n655 VSUBS 0.007324f
C1439 B.n656 VSUBS 0.007324f
C1440 B.n657 VSUBS 0.007324f
C1441 B.n658 VSUBS 0.007324f
C1442 B.n659 VSUBS 0.007324f
C1443 B.n660 VSUBS 0.007324f
C1444 B.n661 VSUBS 0.007324f
C1445 B.n662 VSUBS 0.007324f
C1446 B.n663 VSUBS 0.007324f
C1447 B.n664 VSUBS 0.007324f
C1448 B.n665 VSUBS 0.007324f
C1449 B.n666 VSUBS 0.007324f
C1450 B.n667 VSUBS 0.007324f
C1451 B.n668 VSUBS 0.007324f
C1452 B.n669 VSUBS 0.007324f
C1453 B.n670 VSUBS 0.007324f
C1454 B.n671 VSUBS 0.007324f
C1455 B.n672 VSUBS 0.007324f
C1456 B.n673 VSUBS 0.007324f
C1457 B.n674 VSUBS 0.007324f
C1458 B.n675 VSUBS 0.007324f
C1459 B.n676 VSUBS 0.007324f
C1460 B.n677 VSUBS 0.007324f
C1461 B.n678 VSUBS 0.007324f
C1462 B.n679 VSUBS 0.007324f
C1463 B.n680 VSUBS 0.007324f
C1464 B.n681 VSUBS 0.007324f
C1465 B.n682 VSUBS 0.007324f
C1466 B.n683 VSUBS 0.007324f
C1467 B.n684 VSUBS 0.007324f
C1468 B.n685 VSUBS 0.007324f
C1469 B.n686 VSUBS 0.007324f
C1470 B.n687 VSUBS 0.007324f
C1471 B.n688 VSUBS 0.007324f
C1472 B.n689 VSUBS 0.007324f
C1473 B.n690 VSUBS 0.007324f
C1474 B.n691 VSUBS 0.007324f
C1475 B.n692 VSUBS 0.007324f
C1476 B.n693 VSUBS 0.007324f
C1477 B.n694 VSUBS 0.007324f
C1478 B.n695 VSUBS 0.007324f
C1479 B.n696 VSUBS 0.006893f
C1480 B.n697 VSUBS 0.016968f
C1481 B.n698 VSUBS 0.004093f
C1482 B.n699 VSUBS 0.007324f
C1483 B.n700 VSUBS 0.007324f
C1484 B.n701 VSUBS 0.007324f
C1485 B.n702 VSUBS 0.007324f
C1486 B.n703 VSUBS 0.007324f
C1487 B.n704 VSUBS 0.007324f
C1488 B.n705 VSUBS 0.007324f
C1489 B.n706 VSUBS 0.007324f
C1490 B.n707 VSUBS 0.007324f
C1491 B.n708 VSUBS 0.007324f
C1492 B.n709 VSUBS 0.007324f
C1493 B.n710 VSUBS 0.007324f
C1494 B.n711 VSUBS 0.004093f
C1495 B.n712 VSUBS 0.007324f
C1496 B.n713 VSUBS 0.007324f
C1497 B.n714 VSUBS 0.007324f
C1498 B.n715 VSUBS 0.007324f
C1499 B.n716 VSUBS 0.007324f
C1500 B.n717 VSUBS 0.007324f
C1501 B.n718 VSUBS 0.007324f
C1502 B.n719 VSUBS 0.007324f
C1503 B.n720 VSUBS 0.007324f
C1504 B.n721 VSUBS 0.007324f
C1505 B.n722 VSUBS 0.007324f
C1506 B.n723 VSUBS 0.007324f
C1507 B.n724 VSUBS 0.007324f
C1508 B.n725 VSUBS 0.007324f
C1509 B.n726 VSUBS 0.007324f
C1510 B.n727 VSUBS 0.007324f
C1511 B.n728 VSUBS 0.007324f
C1512 B.n729 VSUBS 0.007324f
C1513 B.n730 VSUBS 0.007324f
C1514 B.n731 VSUBS 0.007324f
C1515 B.n732 VSUBS 0.007324f
C1516 B.n733 VSUBS 0.007324f
C1517 B.n734 VSUBS 0.007324f
C1518 B.n735 VSUBS 0.007324f
C1519 B.n736 VSUBS 0.007324f
C1520 B.n737 VSUBS 0.007324f
C1521 B.n738 VSUBS 0.007324f
C1522 B.n739 VSUBS 0.007324f
C1523 B.n740 VSUBS 0.007324f
C1524 B.n741 VSUBS 0.007324f
C1525 B.n742 VSUBS 0.007324f
C1526 B.n743 VSUBS 0.007324f
C1527 B.n744 VSUBS 0.007324f
C1528 B.n745 VSUBS 0.007324f
C1529 B.n746 VSUBS 0.007324f
C1530 B.n747 VSUBS 0.007324f
C1531 B.n748 VSUBS 0.007324f
C1532 B.n749 VSUBS 0.007324f
C1533 B.n750 VSUBS 0.007324f
C1534 B.n751 VSUBS 0.007324f
C1535 B.n752 VSUBS 0.007324f
C1536 B.n753 VSUBS 0.007324f
C1537 B.n754 VSUBS 0.007324f
C1538 B.n755 VSUBS 0.007324f
C1539 B.n756 VSUBS 0.007324f
C1540 B.n757 VSUBS 0.007324f
C1541 B.n758 VSUBS 0.007324f
C1542 B.n759 VSUBS 0.007324f
C1543 B.n760 VSUBS 0.007324f
C1544 B.n761 VSUBS 0.007324f
C1545 B.n762 VSUBS 0.007324f
C1546 B.n763 VSUBS 0.007324f
C1547 B.n764 VSUBS 0.007324f
C1548 B.n765 VSUBS 0.007324f
C1549 B.n766 VSUBS 0.007324f
C1550 B.n767 VSUBS 0.007324f
C1551 B.n768 VSUBS 0.007324f
C1552 B.n769 VSUBS 0.007324f
C1553 B.n770 VSUBS 0.007324f
C1554 B.n771 VSUBS 0.007324f
C1555 B.n772 VSUBS 0.007324f
C1556 B.n773 VSUBS 0.007324f
C1557 B.n774 VSUBS 0.017241f
C1558 B.n775 VSUBS 0.017241f
C1559 B.n776 VSUBS 0.015931f
C1560 B.n777 VSUBS 0.007324f
C1561 B.n778 VSUBS 0.007324f
C1562 B.n779 VSUBS 0.007324f
C1563 B.n780 VSUBS 0.007324f
C1564 B.n781 VSUBS 0.007324f
C1565 B.n782 VSUBS 0.007324f
C1566 B.n783 VSUBS 0.007324f
C1567 B.n784 VSUBS 0.007324f
C1568 B.n785 VSUBS 0.007324f
C1569 B.n786 VSUBS 0.007324f
C1570 B.n787 VSUBS 0.007324f
C1571 B.n788 VSUBS 0.007324f
C1572 B.n789 VSUBS 0.007324f
C1573 B.n790 VSUBS 0.007324f
C1574 B.n791 VSUBS 0.007324f
C1575 B.n792 VSUBS 0.007324f
C1576 B.n793 VSUBS 0.007324f
C1577 B.n794 VSUBS 0.007324f
C1578 B.n795 VSUBS 0.007324f
C1579 B.n796 VSUBS 0.007324f
C1580 B.n797 VSUBS 0.007324f
C1581 B.n798 VSUBS 0.007324f
C1582 B.n799 VSUBS 0.007324f
C1583 B.n800 VSUBS 0.007324f
C1584 B.n801 VSUBS 0.007324f
C1585 B.n802 VSUBS 0.007324f
C1586 B.n803 VSUBS 0.007324f
C1587 B.n804 VSUBS 0.007324f
C1588 B.n805 VSUBS 0.007324f
C1589 B.n806 VSUBS 0.007324f
C1590 B.n807 VSUBS 0.007324f
C1591 B.n808 VSUBS 0.007324f
C1592 B.n809 VSUBS 0.007324f
C1593 B.n810 VSUBS 0.007324f
C1594 B.n811 VSUBS 0.007324f
C1595 B.n812 VSUBS 0.007324f
C1596 B.n813 VSUBS 0.007324f
C1597 B.n814 VSUBS 0.007324f
C1598 B.n815 VSUBS 0.007324f
C1599 B.n816 VSUBS 0.007324f
C1600 B.n817 VSUBS 0.007324f
C1601 B.n818 VSUBS 0.007324f
C1602 B.n819 VSUBS 0.007324f
C1603 B.n820 VSUBS 0.007324f
C1604 B.n821 VSUBS 0.007324f
C1605 B.n822 VSUBS 0.007324f
C1606 B.n823 VSUBS 0.007324f
C1607 B.n824 VSUBS 0.007324f
C1608 B.n825 VSUBS 0.007324f
C1609 B.n826 VSUBS 0.007324f
C1610 B.n827 VSUBS 0.007324f
C1611 B.n828 VSUBS 0.007324f
C1612 B.n829 VSUBS 0.007324f
C1613 B.n830 VSUBS 0.007324f
C1614 B.n831 VSUBS 0.007324f
C1615 B.n832 VSUBS 0.007324f
C1616 B.n833 VSUBS 0.007324f
C1617 B.n834 VSUBS 0.007324f
C1618 B.n835 VSUBS 0.007324f
C1619 B.n836 VSUBS 0.007324f
C1620 B.n837 VSUBS 0.007324f
C1621 B.n838 VSUBS 0.007324f
C1622 B.n839 VSUBS 0.007324f
C1623 B.n840 VSUBS 0.007324f
C1624 B.n841 VSUBS 0.007324f
C1625 B.n842 VSUBS 0.007324f
C1626 B.n843 VSUBS 0.007324f
C1627 B.n844 VSUBS 0.007324f
C1628 B.n845 VSUBS 0.007324f
C1629 B.n846 VSUBS 0.007324f
C1630 B.n847 VSUBS 0.007324f
C1631 B.n848 VSUBS 0.007324f
C1632 B.n849 VSUBS 0.007324f
C1633 B.n850 VSUBS 0.007324f
C1634 B.n851 VSUBS 0.007324f
C1635 B.n852 VSUBS 0.007324f
C1636 B.n853 VSUBS 0.007324f
C1637 B.n854 VSUBS 0.007324f
C1638 B.n855 VSUBS 0.007324f
C1639 B.n856 VSUBS 0.007324f
C1640 B.n857 VSUBS 0.007324f
C1641 B.n858 VSUBS 0.007324f
C1642 B.n859 VSUBS 0.007324f
C1643 B.n860 VSUBS 0.007324f
C1644 B.n861 VSUBS 0.007324f
C1645 B.n862 VSUBS 0.007324f
C1646 B.n863 VSUBS 0.009557f
C1647 B.n864 VSUBS 0.010181f
C1648 B.n865 VSUBS 0.020245f
.ends

