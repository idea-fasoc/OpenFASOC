* NGSPICE file created from diff_pair_sample_0670.ext - technology: sky130A

.subckt diff_pair_sample_0670 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=1.96
X1 VDD1.t5 VP.t0 VTAIL.t8 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=1.96
X2 VDD2.t5 VN.t0 VTAIL.t5 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=1.96
X3 VDD1.t4 VP.t1 VTAIL.t9 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=1.96
X4 VDD2.t4 VN.t1 VTAIL.t2 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=1.96
X5 B.t8 B.t6 B.t7 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=1.96
X6 B.t5 B.t3 B.t4 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=1.96
X7 VDD2.t3 VN.t2 VTAIL.t3 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=1.96
X8 B.t2 B.t0 B.t1 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0 ps=0 w=1.6 l=1.96
X9 VTAIL.t4 VN.t3 VDD2.t2 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=1.96
X10 VTAIL.t6 VP.t2 VDD1.t3 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=1.96
X11 VDD2.t1 VN.t4 VTAIL.t1 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=1.96
X12 VTAIL.t11 VP.t3 VDD1.t2 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=1.96
X13 VDD1.t1 VP.t4 VTAIL.t10 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.624 pd=3.98 as=0.264 ps=1.93 w=1.6 l=1.96
X14 VDD1.t0 VP.t5 VTAIL.t7 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.624 ps=3.98 w=1.6 l=1.96
X15 VTAIL.t0 VN.t5 VDD2.t0 w_n2802_n1288# sky130_fd_pr__pfet_01v8 ad=0.264 pd=1.93 as=0.264 ps=1.93 w=1.6 l=1.96
R0 B.n321 B.n320 585
R1 B.n322 B.n39 585
R2 B.n324 B.n323 585
R3 B.n325 B.n38 585
R4 B.n327 B.n326 585
R5 B.n328 B.n37 585
R6 B.n330 B.n329 585
R7 B.n331 B.n36 585
R8 B.n333 B.n332 585
R9 B.n334 B.n35 585
R10 B.n336 B.n335 585
R11 B.n338 B.n337 585
R12 B.n339 B.n31 585
R13 B.n341 B.n340 585
R14 B.n342 B.n30 585
R15 B.n344 B.n343 585
R16 B.n345 B.n29 585
R17 B.n347 B.n346 585
R18 B.n348 B.n28 585
R19 B.n350 B.n349 585
R20 B.n351 B.n25 585
R21 B.n354 B.n353 585
R22 B.n355 B.n24 585
R23 B.n357 B.n356 585
R24 B.n358 B.n23 585
R25 B.n360 B.n359 585
R26 B.n361 B.n22 585
R27 B.n363 B.n362 585
R28 B.n364 B.n21 585
R29 B.n366 B.n365 585
R30 B.n367 B.n20 585
R31 B.n369 B.n368 585
R32 B.n319 B.n40 585
R33 B.n318 B.n317 585
R34 B.n316 B.n41 585
R35 B.n315 B.n314 585
R36 B.n313 B.n42 585
R37 B.n312 B.n311 585
R38 B.n310 B.n43 585
R39 B.n309 B.n308 585
R40 B.n307 B.n44 585
R41 B.n306 B.n305 585
R42 B.n304 B.n45 585
R43 B.n303 B.n302 585
R44 B.n301 B.n46 585
R45 B.n300 B.n299 585
R46 B.n298 B.n47 585
R47 B.n297 B.n296 585
R48 B.n295 B.n48 585
R49 B.n294 B.n293 585
R50 B.n292 B.n49 585
R51 B.n291 B.n290 585
R52 B.n289 B.n50 585
R53 B.n288 B.n287 585
R54 B.n286 B.n51 585
R55 B.n285 B.n284 585
R56 B.n283 B.n52 585
R57 B.n282 B.n281 585
R58 B.n280 B.n53 585
R59 B.n279 B.n278 585
R60 B.n277 B.n54 585
R61 B.n276 B.n275 585
R62 B.n274 B.n55 585
R63 B.n273 B.n272 585
R64 B.n271 B.n56 585
R65 B.n270 B.n269 585
R66 B.n268 B.n57 585
R67 B.n267 B.n266 585
R68 B.n265 B.n58 585
R69 B.n264 B.n263 585
R70 B.n262 B.n59 585
R71 B.n261 B.n260 585
R72 B.n259 B.n60 585
R73 B.n258 B.n257 585
R74 B.n256 B.n61 585
R75 B.n255 B.n254 585
R76 B.n253 B.n62 585
R77 B.n252 B.n251 585
R78 B.n250 B.n63 585
R79 B.n249 B.n248 585
R80 B.n247 B.n64 585
R81 B.n246 B.n245 585
R82 B.n244 B.n65 585
R83 B.n243 B.n242 585
R84 B.n241 B.n66 585
R85 B.n240 B.n239 585
R86 B.n238 B.n67 585
R87 B.n237 B.n236 585
R88 B.n235 B.n68 585
R89 B.n234 B.n233 585
R90 B.n232 B.n69 585
R91 B.n231 B.n230 585
R92 B.n229 B.n70 585
R93 B.n228 B.n227 585
R94 B.n226 B.n71 585
R95 B.n225 B.n224 585
R96 B.n223 B.n72 585
R97 B.n222 B.n221 585
R98 B.n220 B.n73 585
R99 B.n219 B.n218 585
R100 B.n217 B.n74 585
R101 B.n216 B.n215 585
R102 B.n214 B.n75 585
R103 B.n165 B.n164 585
R104 B.n166 B.n95 585
R105 B.n168 B.n167 585
R106 B.n169 B.n94 585
R107 B.n171 B.n170 585
R108 B.n172 B.n93 585
R109 B.n174 B.n173 585
R110 B.n175 B.n92 585
R111 B.n177 B.n176 585
R112 B.n178 B.n91 585
R113 B.n180 B.n179 585
R114 B.n182 B.n181 585
R115 B.n183 B.n87 585
R116 B.n185 B.n184 585
R117 B.n186 B.n86 585
R118 B.n188 B.n187 585
R119 B.n189 B.n85 585
R120 B.n191 B.n190 585
R121 B.n192 B.n84 585
R122 B.n194 B.n193 585
R123 B.n195 B.n81 585
R124 B.n198 B.n197 585
R125 B.n199 B.n80 585
R126 B.n201 B.n200 585
R127 B.n202 B.n79 585
R128 B.n204 B.n203 585
R129 B.n205 B.n78 585
R130 B.n207 B.n206 585
R131 B.n208 B.n77 585
R132 B.n210 B.n209 585
R133 B.n211 B.n76 585
R134 B.n213 B.n212 585
R135 B.n163 B.n96 585
R136 B.n162 B.n161 585
R137 B.n160 B.n97 585
R138 B.n159 B.n158 585
R139 B.n157 B.n98 585
R140 B.n156 B.n155 585
R141 B.n154 B.n99 585
R142 B.n153 B.n152 585
R143 B.n151 B.n100 585
R144 B.n150 B.n149 585
R145 B.n148 B.n101 585
R146 B.n147 B.n146 585
R147 B.n145 B.n102 585
R148 B.n144 B.n143 585
R149 B.n142 B.n103 585
R150 B.n141 B.n140 585
R151 B.n139 B.n104 585
R152 B.n138 B.n137 585
R153 B.n136 B.n105 585
R154 B.n135 B.n134 585
R155 B.n133 B.n106 585
R156 B.n132 B.n131 585
R157 B.n130 B.n107 585
R158 B.n129 B.n128 585
R159 B.n127 B.n108 585
R160 B.n126 B.n125 585
R161 B.n124 B.n109 585
R162 B.n123 B.n122 585
R163 B.n121 B.n110 585
R164 B.n120 B.n119 585
R165 B.n118 B.n111 585
R166 B.n117 B.n116 585
R167 B.n115 B.n112 585
R168 B.n114 B.n113 585
R169 B.n2 B.n0 585
R170 B.n421 B.n1 585
R171 B.n420 B.n419 585
R172 B.n418 B.n3 585
R173 B.n417 B.n416 585
R174 B.n415 B.n4 585
R175 B.n414 B.n413 585
R176 B.n412 B.n5 585
R177 B.n411 B.n410 585
R178 B.n409 B.n6 585
R179 B.n408 B.n407 585
R180 B.n406 B.n7 585
R181 B.n405 B.n404 585
R182 B.n403 B.n8 585
R183 B.n402 B.n401 585
R184 B.n400 B.n9 585
R185 B.n399 B.n398 585
R186 B.n397 B.n10 585
R187 B.n396 B.n395 585
R188 B.n394 B.n11 585
R189 B.n393 B.n392 585
R190 B.n391 B.n12 585
R191 B.n390 B.n389 585
R192 B.n388 B.n13 585
R193 B.n387 B.n386 585
R194 B.n385 B.n14 585
R195 B.n384 B.n383 585
R196 B.n382 B.n15 585
R197 B.n381 B.n380 585
R198 B.n379 B.n16 585
R199 B.n378 B.n377 585
R200 B.n376 B.n17 585
R201 B.n375 B.n374 585
R202 B.n373 B.n18 585
R203 B.n372 B.n371 585
R204 B.n370 B.n19 585
R205 B.n423 B.n422 585
R206 B.n164 B.n163 478.086
R207 B.n368 B.n19 478.086
R208 B.n212 B.n75 478.086
R209 B.n320 B.n319 478.086
R210 B.n82 B.t11 294.445
R211 B.n32 B.t1 294.445
R212 B.n88 B.t5 294.445
R213 B.n26 B.t7 294.445
R214 B.n83 B.t10 250.032
R215 B.n33 B.t2 250.032
R216 B.n89 B.t4 250.032
R217 B.n27 B.t8 250.032
R218 B.n82 B.t9 226.495
R219 B.n88 B.t3 226.495
R220 B.n26 B.t6 226.495
R221 B.n32 B.t0 226.495
R222 B.n163 B.n162 163.367
R223 B.n162 B.n97 163.367
R224 B.n158 B.n97 163.367
R225 B.n158 B.n157 163.367
R226 B.n157 B.n156 163.367
R227 B.n156 B.n99 163.367
R228 B.n152 B.n99 163.367
R229 B.n152 B.n151 163.367
R230 B.n151 B.n150 163.367
R231 B.n150 B.n101 163.367
R232 B.n146 B.n101 163.367
R233 B.n146 B.n145 163.367
R234 B.n145 B.n144 163.367
R235 B.n144 B.n103 163.367
R236 B.n140 B.n103 163.367
R237 B.n140 B.n139 163.367
R238 B.n139 B.n138 163.367
R239 B.n138 B.n105 163.367
R240 B.n134 B.n105 163.367
R241 B.n134 B.n133 163.367
R242 B.n133 B.n132 163.367
R243 B.n132 B.n107 163.367
R244 B.n128 B.n107 163.367
R245 B.n128 B.n127 163.367
R246 B.n127 B.n126 163.367
R247 B.n126 B.n109 163.367
R248 B.n122 B.n109 163.367
R249 B.n122 B.n121 163.367
R250 B.n121 B.n120 163.367
R251 B.n120 B.n111 163.367
R252 B.n116 B.n111 163.367
R253 B.n116 B.n115 163.367
R254 B.n115 B.n114 163.367
R255 B.n114 B.n2 163.367
R256 B.n422 B.n2 163.367
R257 B.n422 B.n421 163.367
R258 B.n421 B.n420 163.367
R259 B.n420 B.n3 163.367
R260 B.n416 B.n3 163.367
R261 B.n416 B.n415 163.367
R262 B.n415 B.n414 163.367
R263 B.n414 B.n5 163.367
R264 B.n410 B.n5 163.367
R265 B.n410 B.n409 163.367
R266 B.n409 B.n408 163.367
R267 B.n408 B.n7 163.367
R268 B.n404 B.n7 163.367
R269 B.n404 B.n403 163.367
R270 B.n403 B.n402 163.367
R271 B.n402 B.n9 163.367
R272 B.n398 B.n9 163.367
R273 B.n398 B.n397 163.367
R274 B.n397 B.n396 163.367
R275 B.n396 B.n11 163.367
R276 B.n392 B.n11 163.367
R277 B.n392 B.n391 163.367
R278 B.n391 B.n390 163.367
R279 B.n390 B.n13 163.367
R280 B.n386 B.n13 163.367
R281 B.n386 B.n385 163.367
R282 B.n385 B.n384 163.367
R283 B.n384 B.n15 163.367
R284 B.n380 B.n15 163.367
R285 B.n380 B.n379 163.367
R286 B.n379 B.n378 163.367
R287 B.n378 B.n17 163.367
R288 B.n374 B.n17 163.367
R289 B.n374 B.n373 163.367
R290 B.n373 B.n372 163.367
R291 B.n372 B.n19 163.367
R292 B.n164 B.n95 163.367
R293 B.n168 B.n95 163.367
R294 B.n169 B.n168 163.367
R295 B.n170 B.n169 163.367
R296 B.n170 B.n93 163.367
R297 B.n174 B.n93 163.367
R298 B.n175 B.n174 163.367
R299 B.n176 B.n175 163.367
R300 B.n176 B.n91 163.367
R301 B.n180 B.n91 163.367
R302 B.n181 B.n180 163.367
R303 B.n181 B.n87 163.367
R304 B.n185 B.n87 163.367
R305 B.n186 B.n185 163.367
R306 B.n187 B.n186 163.367
R307 B.n187 B.n85 163.367
R308 B.n191 B.n85 163.367
R309 B.n192 B.n191 163.367
R310 B.n193 B.n192 163.367
R311 B.n193 B.n81 163.367
R312 B.n198 B.n81 163.367
R313 B.n199 B.n198 163.367
R314 B.n200 B.n199 163.367
R315 B.n200 B.n79 163.367
R316 B.n204 B.n79 163.367
R317 B.n205 B.n204 163.367
R318 B.n206 B.n205 163.367
R319 B.n206 B.n77 163.367
R320 B.n210 B.n77 163.367
R321 B.n211 B.n210 163.367
R322 B.n212 B.n211 163.367
R323 B.n216 B.n75 163.367
R324 B.n217 B.n216 163.367
R325 B.n218 B.n217 163.367
R326 B.n218 B.n73 163.367
R327 B.n222 B.n73 163.367
R328 B.n223 B.n222 163.367
R329 B.n224 B.n223 163.367
R330 B.n224 B.n71 163.367
R331 B.n228 B.n71 163.367
R332 B.n229 B.n228 163.367
R333 B.n230 B.n229 163.367
R334 B.n230 B.n69 163.367
R335 B.n234 B.n69 163.367
R336 B.n235 B.n234 163.367
R337 B.n236 B.n235 163.367
R338 B.n236 B.n67 163.367
R339 B.n240 B.n67 163.367
R340 B.n241 B.n240 163.367
R341 B.n242 B.n241 163.367
R342 B.n242 B.n65 163.367
R343 B.n246 B.n65 163.367
R344 B.n247 B.n246 163.367
R345 B.n248 B.n247 163.367
R346 B.n248 B.n63 163.367
R347 B.n252 B.n63 163.367
R348 B.n253 B.n252 163.367
R349 B.n254 B.n253 163.367
R350 B.n254 B.n61 163.367
R351 B.n258 B.n61 163.367
R352 B.n259 B.n258 163.367
R353 B.n260 B.n259 163.367
R354 B.n260 B.n59 163.367
R355 B.n264 B.n59 163.367
R356 B.n265 B.n264 163.367
R357 B.n266 B.n265 163.367
R358 B.n266 B.n57 163.367
R359 B.n270 B.n57 163.367
R360 B.n271 B.n270 163.367
R361 B.n272 B.n271 163.367
R362 B.n272 B.n55 163.367
R363 B.n276 B.n55 163.367
R364 B.n277 B.n276 163.367
R365 B.n278 B.n277 163.367
R366 B.n278 B.n53 163.367
R367 B.n282 B.n53 163.367
R368 B.n283 B.n282 163.367
R369 B.n284 B.n283 163.367
R370 B.n284 B.n51 163.367
R371 B.n288 B.n51 163.367
R372 B.n289 B.n288 163.367
R373 B.n290 B.n289 163.367
R374 B.n290 B.n49 163.367
R375 B.n294 B.n49 163.367
R376 B.n295 B.n294 163.367
R377 B.n296 B.n295 163.367
R378 B.n296 B.n47 163.367
R379 B.n300 B.n47 163.367
R380 B.n301 B.n300 163.367
R381 B.n302 B.n301 163.367
R382 B.n302 B.n45 163.367
R383 B.n306 B.n45 163.367
R384 B.n307 B.n306 163.367
R385 B.n308 B.n307 163.367
R386 B.n308 B.n43 163.367
R387 B.n312 B.n43 163.367
R388 B.n313 B.n312 163.367
R389 B.n314 B.n313 163.367
R390 B.n314 B.n41 163.367
R391 B.n318 B.n41 163.367
R392 B.n319 B.n318 163.367
R393 B.n368 B.n367 163.367
R394 B.n367 B.n366 163.367
R395 B.n366 B.n21 163.367
R396 B.n362 B.n21 163.367
R397 B.n362 B.n361 163.367
R398 B.n361 B.n360 163.367
R399 B.n360 B.n23 163.367
R400 B.n356 B.n23 163.367
R401 B.n356 B.n355 163.367
R402 B.n355 B.n354 163.367
R403 B.n354 B.n25 163.367
R404 B.n349 B.n25 163.367
R405 B.n349 B.n348 163.367
R406 B.n348 B.n347 163.367
R407 B.n347 B.n29 163.367
R408 B.n343 B.n29 163.367
R409 B.n343 B.n342 163.367
R410 B.n342 B.n341 163.367
R411 B.n341 B.n31 163.367
R412 B.n337 B.n31 163.367
R413 B.n337 B.n336 163.367
R414 B.n336 B.n35 163.367
R415 B.n332 B.n35 163.367
R416 B.n332 B.n331 163.367
R417 B.n331 B.n330 163.367
R418 B.n330 B.n37 163.367
R419 B.n326 B.n37 163.367
R420 B.n326 B.n325 163.367
R421 B.n325 B.n324 163.367
R422 B.n324 B.n39 163.367
R423 B.n320 B.n39 163.367
R424 B.n196 B.n83 59.5399
R425 B.n90 B.n89 59.5399
R426 B.n352 B.n27 59.5399
R427 B.n34 B.n33 59.5399
R428 B.n83 B.n82 44.4126
R429 B.n89 B.n88 44.4126
R430 B.n27 B.n26 44.4126
R431 B.n33 B.n32 44.4126
R432 B.n370 B.n369 31.0639
R433 B.n321 B.n40 31.0639
R434 B.n214 B.n213 31.0639
R435 B.n165 B.n96 31.0639
R436 B B.n423 18.0485
R437 B.n369 B.n20 10.6151
R438 B.n365 B.n20 10.6151
R439 B.n365 B.n364 10.6151
R440 B.n364 B.n363 10.6151
R441 B.n363 B.n22 10.6151
R442 B.n359 B.n22 10.6151
R443 B.n359 B.n358 10.6151
R444 B.n358 B.n357 10.6151
R445 B.n357 B.n24 10.6151
R446 B.n353 B.n24 10.6151
R447 B.n351 B.n350 10.6151
R448 B.n350 B.n28 10.6151
R449 B.n346 B.n28 10.6151
R450 B.n346 B.n345 10.6151
R451 B.n345 B.n344 10.6151
R452 B.n344 B.n30 10.6151
R453 B.n340 B.n30 10.6151
R454 B.n340 B.n339 10.6151
R455 B.n339 B.n338 10.6151
R456 B.n335 B.n334 10.6151
R457 B.n334 B.n333 10.6151
R458 B.n333 B.n36 10.6151
R459 B.n329 B.n36 10.6151
R460 B.n329 B.n328 10.6151
R461 B.n328 B.n327 10.6151
R462 B.n327 B.n38 10.6151
R463 B.n323 B.n38 10.6151
R464 B.n323 B.n322 10.6151
R465 B.n322 B.n321 10.6151
R466 B.n215 B.n214 10.6151
R467 B.n215 B.n74 10.6151
R468 B.n219 B.n74 10.6151
R469 B.n220 B.n219 10.6151
R470 B.n221 B.n220 10.6151
R471 B.n221 B.n72 10.6151
R472 B.n225 B.n72 10.6151
R473 B.n226 B.n225 10.6151
R474 B.n227 B.n226 10.6151
R475 B.n227 B.n70 10.6151
R476 B.n231 B.n70 10.6151
R477 B.n232 B.n231 10.6151
R478 B.n233 B.n232 10.6151
R479 B.n233 B.n68 10.6151
R480 B.n237 B.n68 10.6151
R481 B.n238 B.n237 10.6151
R482 B.n239 B.n238 10.6151
R483 B.n239 B.n66 10.6151
R484 B.n243 B.n66 10.6151
R485 B.n244 B.n243 10.6151
R486 B.n245 B.n244 10.6151
R487 B.n245 B.n64 10.6151
R488 B.n249 B.n64 10.6151
R489 B.n250 B.n249 10.6151
R490 B.n251 B.n250 10.6151
R491 B.n251 B.n62 10.6151
R492 B.n255 B.n62 10.6151
R493 B.n256 B.n255 10.6151
R494 B.n257 B.n256 10.6151
R495 B.n257 B.n60 10.6151
R496 B.n261 B.n60 10.6151
R497 B.n262 B.n261 10.6151
R498 B.n263 B.n262 10.6151
R499 B.n263 B.n58 10.6151
R500 B.n267 B.n58 10.6151
R501 B.n268 B.n267 10.6151
R502 B.n269 B.n268 10.6151
R503 B.n269 B.n56 10.6151
R504 B.n273 B.n56 10.6151
R505 B.n274 B.n273 10.6151
R506 B.n275 B.n274 10.6151
R507 B.n275 B.n54 10.6151
R508 B.n279 B.n54 10.6151
R509 B.n280 B.n279 10.6151
R510 B.n281 B.n280 10.6151
R511 B.n281 B.n52 10.6151
R512 B.n285 B.n52 10.6151
R513 B.n286 B.n285 10.6151
R514 B.n287 B.n286 10.6151
R515 B.n287 B.n50 10.6151
R516 B.n291 B.n50 10.6151
R517 B.n292 B.n291 10.6151
R518 B.n293 B.n292 10.6151
R519 B.n293 B.n48 10.6151
R520 B.n297 B.n48 10.6151
R521 B.n298 B.n297 10.6151
R522 B.n299 B.n298 10.6151
R523 B.n299 B.n46 10.6151
R524 B.n303 B.n46 10.6151
R525 B.n304 B.n303 10.6151
R526 B.n305 B.n304 10.6151
R527 B.n305 B.n44 10.6151
R528 B.n309 B.n44 10.6151
R529 B.n310 B.n309 10.6151
R530 B.n311 B.n310 10.6151
R531 B.n311 B.n42 10.6151
R532 B.n315 B.n42 10.6151
R533 B.n316 B.n315 10.6151
R534 B.n317 B.n316 10.6151
R535 B.n317 B.n40 10.6151
R536 B.n166 B.n165 10.6151
R537 B.n167 B.n166 10.6151
R538 B.n167 B.n94 10.6151
R539 B.n171 B.n94 10.6151
R540 B.n172 B.n171 10.6151
R541 B.n173 B.n172 10.6151
R542 B.n173 B.n92 10.6151
R543 B.n177 B.n92 10.6151
R544 B.n178 B.n177 10.6151
R545 B.n179 B.n178 10.6151
R546 B.n183 B.n182 10.6151
R547 B.n184 B.n183 10.6151
R548 B.n184 B.n86 10.6151
R549 B.n188 B.n86 10.6151
R550 B.n189 B.n188 10.6151
R551 B.n190 B.n189 10.6151
R552 B.n190 B.n84 10.6151
R553 B.n194 B.n84 10.6151
R554 B.n195 B.n194 10.6151
R555 B.n197 B.n80 10.6151
R556 B.n201 B.n80 10.6151
R557 B.n202 B.n201 10.6151
R558 B.n203 B.n202 10.6151
R559 B.n203 B.n78 10.6151
R560 B.n207 B.n78 10.6151
R561 B.n208 B.n207 10.6151
R562 B.n209 B.n208 10.6151
R563 B.n209 B.n76 10.6151
R564 B.n213 B.n76 10.6151
R565 B.n161 B.n96 10.6151
R566 B.n161 B.n160 10.6151
R567 B.n160 B.n159 10.6151
R568 B.n159 B.n98 10.6151
R569 B.n155 B.n98 10.6151
R570 B.n155 B.n154 10.6151
R571 B.n154 B.n153 10.6151
R572 B.n153 B.n100 10.6151
R573 B.n149 B.n100 10.6151
R574 B.n149 B.n148 10.6151
R575 B.n148 B.n147 10.6151
R576 B.n147 B.n102 10.6151
R577 B.n143 B.n102 10.6151
R578 B.n143 B.n142 10.6151
R579 B.n142 B.n141 10.6151
R580 B.n141 B.n104 10.6151
R581 B.n137 B.n104 10.6151
R582 B.n137 B.n136 10.6151
R583 B.n136 B.n135 10.6151
R584 B.n135 B.n106 10.6151
R585 B.n131 B.n106 10.6151
R586 B.n131 B.n130 10.6151
R587 B.n130 B.n129 10.6151
R588 B.n129 B.n108 10.6151
R589 B.n125 B.n108 10.6151
R590 B.n125 B.n124 10.6151
R591 B.n124 B.n123 10.6151
R592 B.n123 B.n110 10.6151
R593 B.n119 B.n110 10.6151
R594 B.n119 B.n118 10.6151
R595 B.n118 B.n117 10.6151
R596 B.n117 B.n112 10.6151
R597 B.n113 B.n112 10.6151
R598 B.n113 B.n0 10.6151
R599 B.n419 B.n1 10.6151
R600 B.n419 B.n418 10.6151
R601 B.n418 B.n417 10.6151
R602 B.n417 B.n4 10.6151
R603 B.n413 B.n4 10.6151
R604 B.n413 B.n412 10.6151
R605 B.n412 B.n411 10.6151
R606 B.n411 B.n6 10.6151
R607 B.n407 B.n6 10.6151
R608 B.n407 B.n406 10.6151
R609 B.n406 B.n405 10.6151
R610 B.n405 B.n8 10.6151
R611 B.n401 B.n8 10.6151
R612 B.n401 B.n400 10.6151
R613 B.n400 B.n399 10.6151
R614 B.n399 B.n10 10.6151
R615 B.n395 B.n10 10.6151
R616 B.n395 B.n394 10.6151
R617 B.n394 B.n393 10.6151
R618 B.n393 B.n12 10.6151
R619 B.n389 B.n12 10.6151
R620 B.n389 B.n388 10.6151
R621 B.n388 B.n387 10.6151
R622 B.n387 B.n14 10.6151
R623 B.n383 B.n14 10.6151
R624 B.n383 B.n382 10.6151
R625 B.n382 B.n381 10.6151
R626 B.n381 B.n16 10.6151
R627 B.n377 B.n16 10.6151
R628 B.n377 B.n376 10.6151
R629 B.n376 B.n375 10.6151
R630 B.n375 B.n18 10.6151
R631 B.n371 B.n18 10.6151
R632 B.n371 B.n370 10.6151
R633 B.n353 B.n352 9.36635
R634 B.n335 B.n34 9.36635
R635 B.n179 B.n90 9.36635
R636 B.n197 B.n196 9.36635
R637 B.n423 B.n0 2.81026
R638 B.n423 B.n1 2.81026
R639 B.n352 B.n351 1.24928
R640 B.n338 B.n34 1.24928
R641 B.n182 B.n90 1.24928
R642 B.n196 B.n195 1.24928
R643 VP.n20 VP.n5 183.696
R644 VP.n38 VP.n37 183.696
R645 VP.n19 VP.n18 183.696
R646 VP.n11 VP.n8 161.3
R647 VP.n13 VP.n12 161.3
R648 VP.n14 VP.n7 161.3
R649 VP.n16 VP.n15 161.3
R650 VP.n17 VP.n6 161.3
R651 VP.n36 VP.n0 161.3
R652 VP.n35 VP.n34 161.3
R653 VP.n33 VP.n1 161.3
R654 VP.n32 VP.n31 161.3
R655 VP.n30 VP.n2 161.3
R656 VP.n28 VP.n27 161.3
R657 VP.n26 VP.n3 161.3
R658 VP.n25 VP.n24 161.3
R659 VP.n23 VP.n4 161.3
R660 VP.n22 VP.n21 161.3
R661 VP.n10 VP.n9 57.7491
R662 VP.n9 VP.t4 52.3214
R663 VP.n24 VP.n3 50.6348
R664 VP.n31 VP.n1 50.6348
R665 VP.n12 VP.n7 50.6348
R666 VP.n20 VP.n19 38.2013
R667 VP.n24 VP.n23 30.1864
R668 VP.n35 VP.n1 30.1864
R669 VP.n16 VP.n7 30.1864
R670 VP.n23 VP.n22 24.3439
R671 VP.n28 VP.n3 24.3439
R672 VP.n31 VP.n30 24.3439
R673 VP.n36 VP.n35 24.3439
R674 VP.n17 VP.n16 24.3439
R675 VP.n12 VP.n11 24.3439
R676 VP.n5 VP.t0 19.674
R677 VP.n29 VP.t3 19.674
R678 VP.n37 VP.t1 19.674
R679 VP.n18 VP.t5 19.674
R680 VP.n10 VP.t2 19.674
R681 VP.n9 VP.n8 12.5052
R682 VP.n29 VP.n28 12.1722
R683 VP.n30 VP.n29 12.1722
R684 VP.n11 VP.n10 12.1722
R685 VP.n22 VP.n5 1.94797
R686 VP.n37 VP.n36 1.94797
R687 VP.n18 VP.n17 1.94797
R688 VP.n13 VP.n8 0.189894
R689 VP.n14 VP.n13 0.189894
R690 VP.n15 VP.n14 0.189894
R691 VP.n15 VP.n6 0.189894
R692 VP.n19 VP.n6 0.189894
R693 VP.n21 VP.n20 0.189894
R694 VP.n21 VP.n4 0.189894
R695 VP.n25 VP.n4 0.189894
R696 VP.n26 VP.n25 0.189894
R697 VP.n27 VP.n26 0.189894
R698 VP.n27 VP.n2 0.189894
R699 VP.n32 VP.n2 0.189894
R700 VP.n33 VP.n32 0.189894
R701 VP.n34 VP.n33 0.189894
R702 VP.n34 VP.n0 0.189894
R703 VP.n38 VP.n0 0.189894
R704 VP VP.n38 0.0516364
R705 VTAIL.n11 VTAIL.t2 252.196
R706 VTAIL.n2 VTAIL.t9 252.196
R707 VTAIL.n10 VTAIL.t7 252.196
R708 VTAIL.n7 VTAIL.t3 252.196
R709 VTAIL.n1 VTAIL.n0 231.881
R710 VTAIL.n4 VTAIL.n3 231.881
R711 VTAIL.n9 VTAIL.n8 231.881
R712 VTAIL.n6 VTAIL.n5 231.881
R713 VTAIL.n0 VTAIL.t5 20.3161
R714 VTAIL.n0 VTAIL.t0 20.3161
R715 VTAIL.n3 VTAIL.t8 20.3161
R716 VTAIL.n3 VTAIL.t11 20.3161
R717 VTAIL.n8 VTAIL.t10 20.3161
R718 VTAIL.n8 VTAIL.t6 20.3161
R719 VTAIL.n5 VTAIL.t1 20.3161
R720 VTAIL.n5 VTAIL.t4 20.3161
R721 VTAIL.n6 VTAIL.n4 17.6945
R722 VTAIL.n11 VTAIL.n10 15.7203
R723 VTAIL.n7 VTAIL.n6 1.97464
R724 VTAIL.n10 VTAIL.n9 1.97464
R725 VTAIL.n4 VTAIL.n2 1.97464
R726 VTAIL.n9 VTAIL.n7 1.4574
R727 VTAIL.n2 VTAIL.n1 1.4574
R728 VTAIL VTAIL.n11 1.42291
R729 VTAIL VTAIL.n1 0.552224
R730 VDD1 VDD1.t1 270.414
R731 VDD1.n1 VDD1.t5 270.3
R732 VDD1.n1 VDD1.n0 248.999
R733 VDD1.n3 VDD1.n2 248.56
R734 VDD1.n3 VDD1.n1 33.0806
R735 VDD1.n2 VDD1.t3 20.3161
R736 VDD1.n2 VDD1.t0 20.3161
R737 VDD1.n0 VDD1.t2 20.3161
R738 VDD1.n0 VDD1.t4 20.3161
R739 VDD1 VDD1.n3 0.435845
R740 VN.n13 VN.n12 183.696
R741 VN.n27 VN.n26 183.696
R742 VN.n25 VN.n14 161.3
R743 VN.n24 VN.n23 161.3
R744 VN.n22 VN.n15 161.3
R745 VN.n21 VN.n20 161.3
R746 VN.n19 VN.n16 161.3
R747 VN.n11 VN.n0 161.3
R748 VN.n10 VN.n9 161.3
R749 VN.n8 VN.n1 161.3
R750 VN.n7 VN.n6 161.3
R751 VN.n5 VN.n2 161.3
R752 VN.n4 VN.n3 57.7491
R753 VN.n18 VN.n17 57.7491
R754 VN.n3 VN.t0 52.3214
R755 VN.n17 VN.t2 52.3214
R756 VN.n6 VN.n1 50.6348
R757 VN.n20 VN.n15 50.6348
R758 VN VN.n27 38.5819
R759 VN.n10 VN.n1 30.1864
R760 VN.n24 VN.n15 30.1864
R761 VN.n6 VN.n5 24.3439
R762 VN.n11 VN.n10 24.3439
R763 VN.n20 VN.n19 24.3439
R764 VN.n25 VN.n24 24.3439
R765 VN.n4 VN.t5 19.674
R766 VN.n12 VN.t1 19.674
R767 VN.n18 VN.t3 19.674
R768 VN.n26 VN.t4 19.674
R769 VN.n17 VN.n16 12.5052
R770 VN.n3 VN.n2 12.5052
R771 VN.n5 VN.n4 12.1722
R772 VN.n19 VN.n18 12.1722
R773 VN.n12 VN.n11 1.94797
R774 VN.n26 VN.n25 1.94797
R775 VN.n27 VN.n14 0.189894
R776 VN.n23 VN.n14 0.189894
R777 VN.n23 VN.n22 0.189894
R778 VN.n22 VN.n21 0.189894
R779 VN.n21 VN.n16 0.189894
R780 VN.n7 VN.n2 0.189894
R781 VN.n8 VN.n7 0.189894
R782 VN.n9 VN.n8 0.189894
R783 VN.n9 VN.n0 0.189894
R784 VN.n13 VN.n0 0.189894
R785 VN VN.n13 0.0516364
R786 VDD2.n1 VDD2.t5 270.3
R787 VDD2.n2 VDD2.t1 268.875
R788 VDD2.n1 VDD2.n0 248.999
R789 VDD2 VDD2.n3 248.995
R790 VDD2.n2 VDD2.n1 31.5106
R791 VDD2.n3 VDD2.t2 20.3161
R792 VDD2.n3 VDD2.t3 20.3161
R793 VDD2.n0 VDD2.t0 20.3161
R794 VDD2.n0 VDD2.t4 20.3161
R795 VDD2 VDD2.n2 1.53929
C0 VP w_n2802_n1288# 5.29987f
C1 B VN 0.884856f
C2 VP VN 4.389f
C3 w_n2802_n1288# VTAIL 1.38094f
C4 VDD1 VDD2 1.17967f
C5 VN VTAIL 1.8436f
C6 B VDD1 1.11367f
C7 VDD1 VP 1.42136f
C8 B VDD2 1.17277f
C9 VP VDD2 0.410802f
C10 VDD1 VTAIL 3.51195f
C11 VN w_n2802_n1288# 4.94526f
C12 B VP 1.48257f
C13 VDD2 VTAIL 3.56078f
C14 B VTAIL 1.10666f
C15 VDD1 w_n2802_n1288# 1.39529f
C16 VP VTAIL 1.85774f
C17 VDD1 VN 0.156475f
C18 VDD2 w_n2802_n1288# 1.45914f
C19 B w_n2802_n1288# 5.90458f
C20 VDD2 VN 1.16951f
C21 VDD2 VSUBS 0.893657f
C22 VDD1 VSUBS 1.257078f
C23 VTAIL VSUBS 0.373959f
C24 VN VSUBS 4.61466f
C25 VP VSUBS 1.857755f
C26 B VSUBS 2.949443f
C27 w_n2802_n1288# VSUBS 46.232998f
C28 VDD2.t5 VSUBS 0.134073f
C29 VDD2.t0 VSUBS 0.021932f
C30 VDD2.t4 VSUBS 0.021932f
C31 VDD2.n0 VSUBS 0.082453f
C32 VDD2.n1 VSUBS 1.42456f
C33 VDD2.t1 VSUBS 0.132666f
C34 VDD2.n2 VSUBS 1.23369f
C35 VDD2.t2 VSUBS 0.021932f
C36 VDD2.t3 VSUBS 0.021932f
C37 VDD2.n3 VSUBS 0.082448f
C38 VN.n0 VSUBS 0.046469f
C39 VN.t1 VSUBS 0.323315f
C40 VN.n1 VSUBS 0.044686f
C41 VN.n2 VSUBS 0.347144f
C42 VN.t5 VSUBS 0.323315f
C43 VN.t0 VSUBS 0.581638f
C44 VN.n3 VSUBS 0.27062f
C45 VN.n4 VSUBS 0.289267f
C46 VN.n5 VSUBS 0.065554f
C47 VN.n6 VSUBS 0.085256f
C48 VN.n7 VSUBS 0.046469f
C49 VN.n8 VSUBS 0.046469f
C50 VN.n9 VSUBS 0.046469f
C51 VN.n10 VSUBS 0.093363f
C52 VN.n11 VSUBS 0.047504f
C53 VN.n12 VSUBS 0.293274f
C54 VN.n13 VSUBS 0.051863f
C55 VN.n14 VSUBS 0.046469f
C56 VN.t4 VSUBS 0.323315f
C57 VN.n15 VSUBS 0.044686f
C58 VN.n16 VSUBS 0.347144f
C59 VN.t3 VSUBS 0.323315f
C60 VN.t2 VSUBS 0.581638f
C61 VN.n17 VSUBS 0.27062f
C62 VN.n18 VSUBS 0.289267f
C63 VN.n19 VSUBS 0.065554f
C64 VN.n20 VSUBS 0.085256f
C65 VN.n21 VSUBS 0.046469f
C66 VN.n22 VSUBS 0.046469f
C67 VN.n23 VSUBS 0.046469f
C68 VN.n24 VSUBS 0.093363f
C69 VN.n25 VSUBS 0.047504f
C70 VN.n26 VSUBS 0.293274f
C71 VN.n27 VSUBS 1.67542f
C72 VDD1.t1 VSUBS 0.128209f
C73 VDD1.t5 VSUBS 0.128069f
C74 VDD1.t2 VSUBS 0.02095f
C75 VDD1.t4 VSUBS 0.02095f
C76 VDD1.n0 VSUBS 0.078761f
C77 VDD1.n1 VSUBS 1.42568f
C78 VDD1.t3 VSUBS 0.02095f
C79 VDD1.t0 VSUBS 0.02095f
C80 VDD1.n2 VSUBS 0.078234f
C81 VDD1.n3 VSUBS 1.21258f
C82 VTAIL.t5 VSUBS 0.028997f
C83 VTAIL.t0 VSUBS 0.028997f
C84 VTAIL.n0 VSUBS 0.092344f
C85 VTAIL.n1 VSUBS 0.359188f
C86 VTAIL.t9 VSUBS 0.159953f
C87 VTAIL.n2 VSUBS 0.475776f
C88 VTAIL.t8 VSUBS 0.028997f
C89 VTAIL.t11 VSUBS 0.028997f
C90 VTAIL.n3 VSUBS 0.092344f
C91 VTAIL.n4 VSUBS 1.06188f
C92 VTAIL.t1 VSUBS 0.028997f
C93 VTAIL.t4 VSUBS 0.028997f
C94 VTAIL.n5 VSUBS 0.092344f
C95 VTAIL.n6 VSUBS 1.06188f
C96 VTAIL.t3 VSUBS 0.159954f
C97 VTAIL.n7 VSUBS 0.475776f
C98 VTAIL.t10 VSUBS 0.028997f
C99 VTAIL.t6 VSUBS 0.028997f
C100 VTAIL.n8 VSUBS 0.092344f
C101 VTAIL.n9 VSUBS 0.464303f
C102 VTAIL.t7 VSUBS 0.159954f
C103 VTAIL.n10 VSUBS 0.927462f
C104 VTAIL.t2 VSUBS 0.159953f
C105 VTAIL.n11 VSUBS 0.88669f
C106 VP.n0 VSUBS 0.048811f
C107 VP.t1 VSUBS 0.339607f
C108 VP.n1 VSUBS 0.046938f
C109 VP.n2 VSUBS 0.048811f
C110 VP.t3 VSUBS 0.339607f
C111 VP.n3 VSUBS 0.089552f
C112 VP.n4 VSUBS 0.048811f
C113 VP.t0 VSUBS 0.339607f
C114 VP.n5 VSUBS 0.308051f
C115 VP.n6 VSUBS 0.048811f
C116 VP.t5 VSUBS 0.339607f
C117 VP.n7 VSUBS 0.046938f
C118 VP.n8 VSUBS 0.364636f
C119 VP.t2 VSUBS 0.339607f
C120 VP.t4 VSUBS 0.610946f
C121 VP.n9 VSUBS 0.284257f
C122 VP.n10 VSUBS 0.303842f
C123 VP.n11 VSUBS 0.068857f
C124 VP.n12 VSUBS 0.089552f
C125 VP.n13 VSUBS 0.048811f
C126 VP.n14 VSUBS 0.048811f
C127 VP.n15 VSUBS 0.048811f
C128 VP.n16 VSUBS 0.098067f
C129 VP.n17 VSUBS 0.049897f
C130 VP.n18 VSUBS 0.308051f
C131 VP.n19 VSUBS 1.7276f
C132 VP.n20 VSUBS 1.7734f
C133 VP.n21 VSUBS 0.048811f
C134 VP.n22 VSUBS 0.049897f
C135 VP.n23 VSUBS 0.098067f
C136 VP.n24 VSUBS 0.046938f
C137 VP.n25 VSUBS 0.048811f
C138 VP.n26 VSUBS 0.048811f
C139 VP.n27 VSUBS 0.048811f
C140 VP.n28 VSUBS 0.068857f
C141 VP.n29 VSUBS 0.188133f
C142 VP.n30 VSUBS 0.068857f
C143 VP.n31 VSUBS 0.089552f
C144 VP.n32 VSUBS 0.048811f
C145 VP.n33 VSUBS 0.048811f
C146 VP.n34 VSUBS 0.048811f
C147 VP.n35 VSUBS 0.098067f
C148 VP.n36 VSUBS 0.049897f
C149 VP.n37 VSUBS 0.308051f
C150 VP.n38 VSUBS 0.054477f
C151 B.n0 VSUBS 0.005868f
C152 B.n1 VSUBS 0.005868f
C153 B.n2 VSUBS 0.00928f
C154 B.n3 VSUBS 0.00928f
C155 B.n4 VSUBS 0.00928f
C156 B.n5 VSUBS 0.00928f
C157 B.n6 VSUBS 0.00928f
C158 B.n7 VSUBS 0.00928f
C159 B.n8 VSUBS 0.00928f
C160 B.n9 VSUBS 0.00928f
C161 B.n10 VSUBS 0.00928f
C162 B.n11 VSUBS 0.00928f
C163 B.n12 VSUBS 0.00928f
C164 B.n13 VSUBS 0.00928f
C165 B.n14 VSUBS 0.00928f
C166 B.n15 VSUBS 0.00928f
C167 B.n16 VSUBS 0.00928f
C168 B.n17 VSUBS 0.00928f
C169 B.n18 VSUBS 0.00928f
C170 B.n19 VSUBS 0.020243f
C171 B.n20 VSUBS 0.00928f
C172 B.n21 VSUBS 0.00928f
C173 B.n22 VSUBS 0.00928f
C174 B.n23 VSUBS 0.00928f
C175 B.n24 VSUBS 0.00928f
C176 B.n25 VSUBS 0.00928f
C177 B.t8 VSUBS 0.043469f
C178 B.t7 VSUBS 0.051752f
C179 B.t6 VSUBS 0.20575f
C180 B.n26 VSUBS 0.082056f
C181 B.n27 VSUBS 0.068152f
C182 B.n28 VSUBS 0.00928f
C183 B.n29 VSUBS 0.00928f
C184 B.n30 VSUBS 0.00928f
C185 B.n31 VSUBS 0.00928f
C186 B.t2 VSUBS 0.043469f
C187 B.t1 VSUBS 0.051752f
C188 B.t0 VSUBS 0.20575f
C189 B.n32 VSUBS 0.082056f
C190 B.n33 VSUBS 0.068152f
C191 B.n34 VSUBS 0.021501f
C192 B.n35 VSUBS 0.00928f
C193 B.n36 VSUBS 0.00928f
C194 B.n37 VSUBS 0.00928f
C195 B.n38 VSUBS 0.00928f
C196 B.n39 VSUBS 0.00928f
C197 B.n40 VSUBS 0.021396f
C198 B.n41 VSUBS 0.00928f
C199 B.n42 VSUBS 0.00928f
C200 B.n43 VSUBS 0.00928f
C201 B.n44 VSUBS 0.00928f
C202 B.n45 VSUBS 0.00928f
C203 B.n46 VSUBS 0.00928f
C204 B.n47 VSUBS 0.00928f
C205 B.n48 VSUBS 0.00928f
C206 B.n49 VSUBS 0.00928f
C207 B.n50 VSUBS 0.00928f
C208 B.n51 VSUBS 0.00928f
C209 B.n52 VSUBS 0.00928f
C210 B.n53 VSUBS 0.00928f
C211 B.n54 VSUBS 0.00928f
C212 B.n55 VSUBS 0.00928f
C213 B.n56 VSUBS 0.00928f
C214 B.n57 VSUBS 0.00928f
C215 B.n58 VSUBS 0.00928f
C216 B.n59 VSUBS 0.00928f
C217 B.n60 VSUBS 0.00928f
C218 B.n61 VSUBS 0.00928f
C219 B.n62 VSUBS 0.00928f
C220 B.n63 VSUBS 0.00928f
C221 B.n64 VSUBS 0.00928f
C222 B.n65 VSUBS 0.00928f
C223 B.n66 VSUBS 0.00928f
C224 B.n67 VSUBS 0.00928f
C225 B.n68 VSUBS 0.00928f
C226 B.n69 VSUBS 0.00928f
C227 B.n70 VSUBS 0.00928f
C228 B.n71 VSUBS 0.00928f
C229 B.n72 VSUBS 0.00928f
C230 B.n73 VSUBS 0.00928f
C231 B.n74 VSUBS 0.00928f
C232 B.n75 VSUBS 0.020243f
C233 B.n76 VSUBS 0.00928f
C234 B.n77 VSUBS 0.00928f
C235 B.n78 VSUBS 0.00928f
C236 B.n79 VSUBS 0.00928f
C237 B.n80 VSUBS 0.00928f
C238 B.n81 VSUBS 0.00928f
C239 B.t10 VSUBS 0.043469f
C240 B.t11 VSUBS 0.051752f
C241 B.t9 VSUBS 0.20575f
C242 B.n82 VSUBS 0.082056f
C243 B.n83 VSUBS 0.068152f
C244 B.n84 VSUBS 0.00928f
C245 B.n85 VSUBS 0.00928f
C246 B.n86 VSUBS 0.00928f
C247 B.n87 VSUBS 0.00928f
C248 B.t4 VSUBS 0.043469f
C249 B.t5 VSUBS 0.051752f
C250 B.t3 VSUBS 0.20575f
C251 B.n88 VSUBS 0.082056f
C252 B.n89 VSUBS 0.068152f
C253 B.n90 VSUBS 0.021501f
C254 B.n91 VSUBS 0.00928f
C255 B.n92 VSUBS 0.00928f
C256 B.n93 VSUBS 0.00928f
C257 B.n94 VSUBS 0.00928f
C258 B.n95 VSUBS 0.00928f
C259 B.n96 VSUBS 0.020243f
C260 B.n97 VSUBS 0.00928f
C261 B.n98 VSUBS 0.00928f
C262 B.n99 VSUBS 0.00928f
C263 B.n100 VSUBS 0.00928f
C264 B.n101 VSUBS 0.00928f
C265 B.n102 VSUBS 0.00928f
C266 B.n103 VSUBS 0.00928f
C267 B.n104 VSUBS 0.00928f
C268 B.n105 VSUBS 0.00928f
C269 B.n106 VSUBS 0.00928f
C270 B.n107 VSUBS 0.00928f
C271 B.n108 VSUBS 0.00928f
C272 B.n109 VSUBS 0.00928f
C273 B.n110 VSUBS 0.00928f
C274 B.n111 VSUBS 0.00928f
C275 B.n112 VSUBS 0.00928f
C276 B.n113 VSUBS 0.00928f
C277 B.n114 VSUBS 0.00928f
C278 B.n115 VSUBS 0.00928f
C279 B.n116 VSUBS 0.00928f
C280 B.n117 VSUBS 0.00928f
C281 B.n118 VSUBS 0.00928f
C282 B.n119 VSUBS 0.00928f
C283 B.n120 VSUBS 0.00928f
C284 B.n121 VSUBS 0.00928f
C285 B.n122 VSUBS 0.00928f
C286 B.n123 VSUBS 0.00928f
C287 B.n124 VSUBS 0.00928f
C288 B.n125 VSUBS 0.00928f
C289 B.n126 VSUBS 0.00928f
C290 B.n127 VSUBS 0.00928f
C291 B.n128 VSUBS 0.00928f
C292 B.n129 VSUBS 0.00928f
C293 B.n130 VSUBS 0.00928f
C294 B.n131 VSUBS 0.00928f
C295 B.n132 VSUBS 0.00928f
C296 B.n133 VSUBS 0.00928f
C297 B.n134 VSUBS 0.00928f
C298 B.n135 VSUBS 0.00928f
C299 B.n136 VSUBS 0.00928f
C300 B.n137 VSUBS 0.00928f
C301 B.n138 VSUBS 0.00928f
C302 B.n139 VSUBS 0.00928f
C303 B.n140 VSUBS 0.00928f
C304 B.n141 VSUBS 0.00928f
C305 B.n142 VSUBS 0.00928f
C306 B.n143 VSUBS 0.00928f
C307 B.n144 VSUBS 0.00928f
C308 B.n145 VSUBS 0.00928f
C309 B.n146 VSUBS 0.00928f
C310 B.n147 VSUBS 0.00928f
C311 B.n148 VSUBS 0.00928f
C312 B.n149 VSUBS 0.00928f
C313 B.n150 VSUBS 0.00928f
C314 B.n151 VSUBS 0.00928f
C315 B.n152 VSUBS 0.00928f
C316 B.n153 VSUBS 0.00928f
C317 B.n154 VSUBS 0.00928f
C318 B.n155 VSUBS 0.00928f
C319 B.n156 VSUBS 0.00928f
C320 B.n157 VSUBS 0.00928f
C321 B.n158 VSUBS 0.00928f
C322 B.n159 VSUBS 0.00928f
C323 B.n160 VSUBS 0.00928f
C324 B.n161 VSUBS 0.00928f
C325 B.n162 VSUBS 0.00928f
C326 B.n163 VSUBS 0.020243f
C327 B.n164 VSUBS 0.02179f
C328 B.n165 VSUBS 0.02179f
C329 B.n166 VSUBS 0.00928f
C330 B.n167 VSUBS 0.00928f
C331 B.n168 VSUBS 0.00928f
C332 B.n169 VSUBS 0.00928f
C333 B.n170 VSUBS 0.00928f
C334 B.n171 VSUBS 0.00928f
C335 B.n172 VSUBS 0.00928f
C336 B.n173 VSUBS 0.00928f
C337 B.n174 VSUBS 0.00928f
C338 B.n175 VSUBS 0.00928f
C339 B.n176 VSUBS 0.00928f
C340 B.n177 VSUBS 0.00928f
C341 B.n178 VSUBS 0.00928f
C342 B.n179 VSUBS 0.008734f
C343 B.n180 VSUBS 0.00928f
C344 B.n181 VSUBS 0.00928f
C345 B.n182 VSUBS 0.005186f
C346 B.n183 VSUBS 0.00928f
C347 B.n184 VSUBS 0.00928f
C348 B.n185 VSUBS 0.00928f
C349 B.n186 VSUBS 0.00928f
C350 B.n187 VSUBS 0.00928f
C351 B.n188 VSUBS 0.00928f
C352 B.n189 VSUBS 0.00928f
C353 B.n190 VSUBS 0.00928f
C354 B.n191 VSUBS 0.00928f
C355 B.n192 VSUBS 0.00928f
C356 B.n193 VSUBS 0.00928f
C357 B.n194 VSUBS 0.00928f
C358 B.n195 VSUBS 0.005186f
C359 B.n196 VSUBS 0.021501f
C360 B.n197 VSUBS 0.008734f
C361 B.n198 VSUBS 0.00928f
C362 B.n199 VSUBS 0.00928f
C363 B.n200 VSUBS 0.00928f
C364 B.n201 VSUBS 0.00928f
C365 B.n202 VSUBS 0.00928f
C366 B.n203 VSUBS 0.00928f
C367 B.n204 VSUBS 0.00928f
C368 B.n205 VSUBS 0.00928f
C369 B.n206 VSUBS 0.00928f
C370 B.n207 VSUBS 0.00928f
C371 B.n208 VSUBS 0.00928f
C372 B.n209 VSUBS 0.00928f
C373 B.n210 VSUBS 0.00928f
C374 B.n211 VSUBS 0.00928f
C375 B.n212 VSUBS 0.02179f
C376 B.n213 VSUBS 0.02179f
C377 B.n214 VSUBS 0.020243f
C378 B.n215 VSUBS 0.00928f
C379 B.n216 VSUBS 0.00928f
C380 B.n217 VSUBS 0.00928f
C381 B.n218 VSUBS 0.00928f
C382 B.n219 VSUBS 0.00928f
C383 B.n220 VSUBS 0.00928f
C384 B.n221 VSUBS 0.00928f
C385 B.n222 VSUBS 0.00928f
C386 B.n223 VSUBS 0.00928f
C387 B.n224 VSUBS 0.00928f
C388 B.n225 VSUBS 0.00928f
C389 B.n226 VSUBS 0.00928f
C390 B.n227 VSUBS 0.00928f
C391 B.n228 VSUBS 0.00928f
C392 B.n229 VSUBS 0.00928f
C393 B.n230 VSUBS 0.00928f
C394 B.n231 VSUBS 0.00928f
C395 B.n232 VSUBS 0.00928f
C396 B.n233 VSUBS 0.00928f
C397 B.n234 VSUBS 0.00928f
C398 B.n235 VSUBS 0.00928f
C399 B.n236 VSUBS 0.00928f
C400 B.n237 VSUBS 0.00928f
C401 B.n238 VSUBS 0.00928f
C402 B.n239 VSUBS 0.00928f
C403 B.n240 VSUBS 0.00928f
C404 B.n241 VSUBS 0.00928f
C405 B.n242 VSUBS 0.00928f
C406 B.n243 VSUBS 0.00928f
C407 B.n244 VSUBS 0.00928f
C408 B.n245 VSUBS 0.00928f
C409 B.n246 VSUBS 0.00928f
C410 B.n247 VSUBS 0.00928f
C411 B.n248 VSUBS 0.00928f
C412 B.n249 VSUBS 0.00928f
C413 B.n250 VSUBS 0.00928f
C414 B.n251 VSUBS 0.00928f
C415 B.n252 VSUBS 0.00928f
C416 B.n253 VSUBS 0.00928f
C417 B.n254 VSUBS 0.00928f
C418 B.n255 VSUBS 0.00928f
C419 B.n256 VSUBS 0.00928f
C420 B.n257 VSUBS 0.00928f
C421 B.n258 VSUBS 0.00928f
C422 B.n259 VSUBS 0.00928f
C423 B.n260 VSUBS 0.00928f
C424 B.n261 VSUBS 0.00928f
C425 B.n262 VSUBS 0.00928f
C426 B.n263 VSUBS 0.00928f
C427 B.n264 VSUBS 0.00928f
C428 B.n265 VSUBS 0.00928f
C429 B.n266 VSUBS 0.00928f
C430 B.n267 VSUBS 0.00928f
C431 B.n268 VSUBS 0.00928f
C432 B.n269 VSUBS 0.00928f
C433 B.n270 VSUBS 0.00928f
C434 B.n271 VSUBS 0.00928f
C435 B.n272 VSUBS 0.00928f
C436 B.n273 VSUBS 0.00928f
C437 B.n274 VSUBS 0.00928f
C438 B.n275 VSUBS 0.00928f
C439 B.n276 VSUBS 0.00928f
C440 B.n277 VSUBS 0.00928f
C441 B.n278 VSUBS 0.00928f
C442 B.n279 VSUBS 0.00928f
C443 B.n280 VSUBS 0.00928f
C444 B.n281 VSUBS 0.00928f
C445 B.n282 VSUBS 0.00928f
C446 B.n283 VSUBS 0.00928f
C447 B.n284 VSUBS 0.00928f
C448 B.n285 VSUBS 0.00928f
C449 B.n286 VSUBS 0.00928f
C450 B.n287 VSUBS 0.00928f
C451 B.n288 VSUBS 0.00928f
C452 B.n289 VSUBS 0.00928f
C453 B.n290 VSUBS 0.00928f
C454 B.n291 VSUBS 0.00928f
C455 B.n292 VSUBS 0.00928f
C456 B.n293 VSUBS 0.00928f
C457 B.n294 VSUBS 0.00928f
C458 B.n295 VSUBS 0.00928f
C459 B.n296 VSUBS 0.00928f
C460 B.n297 VSUBS 0.00928f
C461 B.n298 VSUBS 0.00928f
C462 B.n299 VSUBS 0.00928f
C463 B.n300 VSUBS 0.00928f
C464 B.n301 VSUBS 0.00928f
C465 B.n302 VSUBS 0.00928f
C466 B.n303 VSUBS 0.00928f
C467 B.n304 VSUBS 0.00928f
C468 B.n305 VSUBS 0.00928f
C469 B.n306 VSUBS 0.00928f
C470 B.n307 VSUBS 0.00928f
C471 B.n308 VSUBS 0.00928f
C472 B.n309 VSUBS 0.00928f
C473 B.n310 VSUBS 0.00928f
C474 B.n311 VSUBS 0.00928f
C475 B.n312 VSUBS 0.00928f
C476 B.n313 VSUBS 0.00928f
C477 B.n314 VSUBS 0.00928f
C478 B.n315 VSUBS 0.00928f
C479 B.n316 VSUBS 0.00928f
C480 B.n317 VSUBS 0.00928f
C481 B.n318 VSUBS 0.00928f
C482 B.n319 VSUBS 0.020243f
C483 B.n320 VSUBS 0.02179f
C484 B.n321 VSUBS 0.020637f
C485 B.n322 VSUBS 0.00928f
C486 B.n323 VSUBS 0.00928f
C487 B.n324 VSUBS 0.00928f
C488 B.n325 VSUBS 0.00928f
C489 B.n326 VSUBS 0.00928f
C490 B.n327 VSUBS 0.00928f
C491 B.n328 VSUBS 0.00928f
C492 B.n329 VSUBS 0.00928f
C493 B.n330 VSUBS 0.00928f
C494 B.n331 VSUBS 0.00928f
C495 B.n332 VSUBS 0.00928f
C496 B.n333 VSUBS 0.00928f
C497 B.n334 VSUBS 0.00928f
C498 B.n335 VSUBS 0.008734f
C499 B.n336 VSUBS 0.00928f
C500 B.n337 VSUBS 0.00928f
C501 B.n338 VSUBS 0.005186f
C502 B.n339 VSUBS 0.00928f
C503 B.n340 VSUBS 0.00928f
C504 B.n341 VSUBS 0.00928f
C505 B.n342 VSUBS 0.00928f
C506 B.n343 VSUBS 0.00928f
C507 B.n344 VSUBS 0.00928f
C508 B.n345 VSUBS 0.00928f
C509 B.n346 VSUBS 0.00928f
C510 B.n347 VSUBS 0.00928f
C511 B.n348 VSUBS 0.00928f
C512 B.n349 VSUBS 0.00928f
C513 B.n350 VSUBS 0.00928f
C514 B.n351 VSUBS 0.005186f
C515 B.n352 VSUBS 0.021501f
C516 B.n353 VSUBS 0.008734f
C517 B.n354 VSUBS 0.00928f
C518 B.n355 VSUBS 0.00928f
C519 B.n356 VSUBS 0.00928f
C520 B.n357 VSUBS 0.00928f
C521 B.n358 VSUBS 0.00928f
C522 B.n359 VSUBS 0.00928f
C523 B.n360 VSUBS 0.00928f
C524 B.n361 VSUBS 0.00928f
C525 B.n362 VSUBS 0.00928f
C526 B.n363 VSUBS 0.00928f
C527 B.n364 VSUBS 0.00928f
C528 B.n365 VSUBS 0.00928f
C529 B.n366 VSUBS 0.00928f
C530 B.n367 VSUBS 0.00928f
C531 B.n368 VSUBS 0.02179f
C532 B.n369 VSUBS 0.02179f
C533 B.n370 VSUBS 0.020243f
C534 B.n371 VSUBS 0.00928f
C535 B.n372 VSUBS 0.00928f
C536 B.n373 VSUBS 0.00928f
C537 B.n374 VSUBS 0.00928f
C538 B.n375 VSUBS 0.00928f
C539 B.n376 VSUBS 0.00928f
C540 B.n377 VSUBS 0.00928f
C541 B.n378 VSUBS 0.00928f
C542 B.n379 VSUBS 0.00928f
C543 B.n380 VSUBS 0.00928f
C544 B.n381 VSUBS 0.00928f
C545 B.n382 VSUBS 0.00928f
C546 B.n383 VSUBS 0.00928f
C547 B.n384 VSUBS 0.00928f
C548 B.n385 VSUBS 0.00928f
C549 B.n386 VSUBS 0.00928f
C550 B.n387 VSUBS 0.00928f
C551 B.n388 VSUBS 0.00928f
C552 B.n389 VSUBS 0.00928f
C553 B.n390 VSUBS 0.00928f
C554 B.n391 VSUBS 0.00928f
C555 B.n392 VSUBS 0.00928f
C556 B.n393 VSUBS 0.00928f
C557 B.n394 VSUBS 0.00928f
C558 B.n395 VSUBS 0.00928f
C559 B.n396 VSUBS 0.00928f
C560 B.n397 VSUBS 0.00928f
C561 B.n398 VSUBS 0.00928f
C562 B.n399 VSUBS 0.00928f
C563 B.n400 VSUBS 0.00928f
C564 B.n401 VSUBS 0.00928f
C565 B.n402 VSUBS 0.00928f
C566 B.n403 VSUBS 0.00928f
C567 B.n404 VSUBS 0.00928f
C568 B.n405 VSUBS 0.00928f
C569 B.n406 VSUBS 0.00928f
C570 B.n407 VSUBS 0.00928f
C571 B.n408 VSUBS 0.00928f
C572 B.n409 VSUBS 0.00928f
C573 B.n410 VSUBS 0.00928f
C574 B.n411 VSUBS 0.00928f
C575 B.n412 VSUBS 0.00928f
C576 B.n413 VSUBS 0.00928f
C577 B.n414 VSUBS 0.00928f
C578 B.n415 VSUBS 0.00928f
C579 B.n416 VSUBS 0.00928f
C580 B.n417 VSUBS 0.00928f
C581 B.n418 VSUBS 0.00928f
C582 B.n419 VSUBS 0.00928f
C583 B.n420 VSUBS 0.00928f
C584 B.n421 VSUBS 0.00928f
C585 B.n422 VSUBS 0.00928f
C586 B.n423 VSUBS 0.021013f
.ends

