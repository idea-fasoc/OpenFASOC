* NGSPICE file created from diff_pair_sample_0631.ext - technology: sky130A

.subckt diff_pair_sample_0631 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VN.t0 VDD2.t2 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=1.63845 ps=10.26 w=9.93 l=3.6
X1 B.t11 B.t9 B.t10 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=3.6
X2 B.t8 B.t6 B.t7 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=3.6
X3 B.t5 B.t3 B.t4 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=3.6
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=1.63845 pd=10.26 as=3.8727 ps=20.64 w=9.93 l=3.6
X5 B.t2 B.t0 B.t1 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=0 ps=0 w=9.93 l=3.6
X6 VTAIL.t2 VN.t2 VDD2.t3 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=1.63845 ps=10.26 w=9.93 l=3.6
X7 VTAIL.t7 VP.t0 VDD1.t3 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=1.63845 ps=10.26 w=9.93 l=3.6
X8 VDD1.t2 VP.t1 VTAIL.t0 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=1.63845 pd=10.26 as=3.8727 ps=20.64 w=9.93 l=3.6
X9 VTAIL.t5 VP.t2 VDD1.t1 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=3.8727 pd=20.64 as=1.63845 ps=10.26 w=9.93 l=3.6
X10 VDD1.t0 VP.t3 VTAIL.t6 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=1.63845 pd=10.26 as=3.8727 ps=20.64 w=9.93 l=3.6
X11 VDD2.t1 VN.t3 VTAIL.t1 w_n3328_n2954# sky130_fd_pr__pfet_01v8 ad=1.63845 pd=10.26 as=3.8727 ps=20.64 w=9.93 l=3.6
R0 VN.n1 VN.t1 101.349
R1 VN.n0 VN.t0 101.349
R2 VN.n0 VN.t3 100.105
R3 VN.n1 VN.t2 100.105
R4 VN VN.n1 50.1709
R5 VN VN.n0 2.09897
R6 VDD2.n2 VDD2.n0 118.975
R7 VDD2.n2 VDD2.n1 76.537
R8 VDD2.n1 VDD2.t3 3.27391
R9 VDD2.n1 VDD2.t0 3.27391
R10 VDD2.n0 VDD2.t2 3.27391
R11 VDD2.n0 VDD2.t1 3.27391
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n426 VTAIL.n378 756.745
R14 VTAIL.n48 VTAIL.n0 756.745
R15 VTAIL.n102 VTAIL.n54 756.745
R16 VTAIL.n156 VTAIL.n108 756.745
R17 VTAIL.n372 VTAIL.n324 756.745
R18 VTAIL.n318 VTAIL.n270 756.745
R19 VTAIL.n264 VTAIL.n216 756.745
R20 VTAIL.n210 VTAIL.n162 756.745
R21 VTAIL.n394 VTAIL.n393 585
R22 VTAIL.n399 VTAIL.n398 585
R23 VTAIL.n401 VTAIL.n400 585
R24 VTAIL.n390 VTAIL.n389 585
R25 VTAIL.n407 VTAIL.n406 585
R26 VTAIL.n409 VTAIL.n408 585
R27 VTAIL.n386 VTAIL.n385 585
R28 VTAIL.n416 VTAIL.n415 585
R29 VTAIL.n417 VTAIL.n384 585
R30 VTAIL.n419 VTAIL.n418 585
R31 VTAIL.n382 VTAIL.n381 585
R32 VTAIL.n425 VTAIL.n424 585
R33 VTAIL.n427 VTAIL.n426 585
R34 VTAIL.n16 VTAIL.n15 585
R35 VTAIL.n21 VTAIL.n20 585
R36 VTAIL.n23 VTAIL.n22 585
R37 VTAIL.n12 VTAIL.n11 585
R38 VTAIL.n29 VTAIL.n28 585
R39 VTAIL.n31 VTAIL.n30 585
R40 VTAIL.n8 VTAIL.n7 585
R41 VTAIL.n38 VTAIL.n37 585
R42 VTAIL.n39 VTAIL.n6 585
R43 VTAIL.n41 VTAIL.n40 585
R44 VTAIL.n4 VTAIL.n3 585
R45 VTAIL.n47 VTAIL.n46 585
R46 VTAIL.n49 VTAIL.n48 585
R47 VTAIL.n70 VTAIL.n69 585
R48 VTAIL.n75 VTAIL.n74 585
R49 VTAIL.n77 VTAIL.n76 585
R50 VTAIL.n66 VTAIL.n65 585
R51 VTAIL.n83 VTAIL.n82 585
R52 VTAIL.n85 VTAIL.n84 585
R53 VTAIL.n62 VTAIL.n61 585
R54 VTAIL.n92 VTAIL.n91 585
R55 VTAIL.n93 VTAIL.n60 585
R56 VTAIL.n95 VTAIL.n94 585
R57 VTAIL.n58 VTAIL.n57 585
R58 VTAIL.n101 VTAIL.n100 585
R59 VTAIL.n103 VTAIL.n102 585
R60 VTAIL.n124 VTAIL.n123 585
R61 VTAIL.n129 VTAIL.n128 585
R62 VTAIL.n131 VTAIL.n130 585
R63 VTAIL.n120 VTAIL.n119 585
R64 VTAIL.n137 VTAIL.n136 585
R65 VTAIL.n139 VTAIL.n138 585
R66 VTAIL.n116 VTAIL.n115 585
R67 VTAIL.n146 VTAIL.n145 585
R68 VTAIL.n147 VTAIL.n114 585
R69 VTAIL.n149 VTAIL.n148 585
R70 VTAIL.n112 VTAIL.n111 585
R71 VTAIL.n155 VTAIL.n154 585
R72 VTAIL.n157 VTAIL.n156 585
R73 VTAIL.n373 VTAIL.n372 585
R74 VTAIL.n371 VTAIL.n370 585
R75 VTAIL.n328 VTAIL.n327 585
R76 VTAIL.n365 VTAIL.n364 585
R77 VTAIL.n363 VTAIL.n330 585
R78 VTAIL.n362 VTAIL.n361 585
R79 VTAIL.n333 VTAIL.n331 585
R80 VTAIL.n356 VTAIL.n355 585
R81 VTAIL.n354 VTAIL.n353 585
R82 VTAIL.n337 VTAIL.n336 585
R83 VTAIL.n348 VTAIL.n347 585
R84 VTAIL.n346 VTAIL.n345 585
R85 VTAIL.n341 VTAIL.n340 585
R86 VTAIL.n319 VTAIL.n318 585
R87 VTAIL.n317 VTAIL.n316 585
R88 VTAIL.n274 VTAIL.n273 585
R89 VTAIL.n311 VTAIL.n310 585
R90 VTAIL.n309 VTAIL.n276 585
R91 VTAIL.n308 VTAIL.n307 585
R92 VTAIL.n279 VTAIL.n277 585
R93 VTAIL.n302 VTAIL.n301 585
R94 VTAIL.n300 VTAIL.n299 585
R95 VTAIL.n283 VTAIL.n282 585
R96 VTAIL.n294 VTAIL.n293 585
R97 VTAIL.n292 VTAIL.n291 585
R98 VTAIL.n287 VTAIL.n286 585
R99 VTAIL.n265 VTAIL.n264 585
R100 VTAIL.n263 VTAIL.n262 585
R101 VTAIL.n220 VTAIL.n219 585
R102 VTAIL.n257 VTAIL.n256 585
R103 VTAIL.n255 VTAIL.n222 585
R104 VTAIL.n254 VTAIL.n253 585
R105 VTAIL.n225 VTAIL.n223 585
R106 VTAIL.n248 VTAIL.n247 585
R107 VTAIL.n246 VTAIL.n245 585
R108 VTAIL.n229 VTAIL.n228 585
R109 VTAIL.n240 VTAIL.n239 585
R110 VTAIL.n238 VTAIL.n237 585
R111 VTAIL.n233 VTAIL.n232 585
R112 VTAIL.n211 VTAIL.n210 585
R113 VTAIL.n209 VTAIL.n208 585
R114 VTAIL.n166 VTAIL.n165 585
R115 VTAIL.n203 VTAIL.n202 585
R116 VTAIL.n201 VTAIL.n168 585
R117 VTAIL.n200 VTAIL.n199 585
R118 VTAIL.n171 VTAIL.n169 585
R119 VTAIL.n194 VTAIL.n193 585
R120 VTAIL.n192 VTAIL.n191 585
R121 VTAIL.n175 VTAIL.n174 585
R122 VTAIL.n186 VTAIL.n185 585
R123 VTAIL.n184 VTAIL.n183 585
R124 VTAIL.n179 VTAIL.n178 585
R125 VTAIL.n395 VTAIL.t1 329.038
R126 VTAIL.n17 VTAIL.t4 329.038
R127 VTAIL.n71 VTAIL.t6 329.038
R128 VTAIL.n125 VTAIL.t5 329.038
R129 VTAIL.n342 VTAIL.t0 329.038
R130 VTAIL.n288 VTAIL.t7 329.038
R131 VTAIL.n234 VTAIL.t3 329.038
R132 VTAIL.n180 VTAIL.t2 329.038
R133 VTAIL.n399 VTAIL.n393 171.744
R134 VTAIL.n400 VTAIL.n399 171.744
R135 VTAIL.n400 VTAIL.n389 171.744
R136 VTAIL.n407 VTAIL.n389 171.744
R137 VTAIL.n408 VTAIL.n407 171.744
R138 VTAIL.n408 VTAIL.n385 171.744
R139 VTAIL.n416 VTAIL.n385 171.744
R140 VTAIL.n417 VTAIL.n416 171.744
R141 VTAIL.n418 VTAIL.n417 171.744
R142 VTAIL.n418 VTAIL.n381 171.744
R143 VTAIL.n425 VTAIL.n381 171.744
R144 VTAIL.n426 VTAIL.n425 171.744
R145 VTAIL.n21 VTAIL.n15 171.744
R146 VTAIL.n22 VTAIL.n21 171.744
R147 VTAIL.n22 VTAIL.n11 171.744
R148 VTAIL.n29 VTAIL.n11 171.744
R149 VTAIL.n30 VTAIL.n29 171.744
R150 VTAIL.n30 VTAIL.n7 171.744
R151 VTAIL.n38 VTAIL.n7 171.744
R152 VTAIL.n39 VTAIL.n38 171.744
R153 VTAIL.n40 VTAIL.n39 171.744
R154 VTAIL.n40 VTAIL.n3 171.744
R155 VTAIL.n47 VTAIL.n3 171.744
R156 VTAIL.n48 VTAIL.n47 171.744
R157 VTAIL.n75 VTAIL.n69 171.744
R158 VTAIL.n76 VTAIL.n75 171.744
R159 VTAIL.n76 VTAIL.n65 171.744
R160 VTAIL.n83 VTAIL.n65 171.744
R161 VTAIL.n84 VTAIL.n83 171.744
R162 VTAIL.n84 VTAIL.n61 171.744
R163 VTAIL.n92 VTAIL.n61 171.744
R164 VTAIL.n93 VTAIL.n92 171.744
R165 VTAIL.n94 VTAIL.n93 171.744
R166 VTAIL.n94 VTAIL.n57 171.744
R167 VTAIL.n101 VTAIL.n57 171.744
R168 VTAIL.n102 VTAIL.n101 171.744
R169 VTAIL.n129 VTAIL.n123 171.744
R170 VTAIL.n130 VTAIL.n129 171.744
R171 VTAIL.n130 VTAIL.n119 171.744
R172 VTAIL.n137 VTAIL.n119 171.744
R173 VTAIL.n138 VTAIL.n137 171.744
R174 VTAIL.n138 VTAIL.n115 171.744
R175 VTAIL.n146 VTAIL.n115 171.744
R176 VTAIL.n147 VTAIL.n146 171.744
R177 VTAIL.n148 VTAIL.n147 171.744
R178 VTAIL.n148 VTAIL.n111 171.744
R179 VTAIL.n155 VTAIL.n111 171.744
R180 VTAIL.n156 VTAIL.n155 171.744
R181 VTAIL.n372 VTAIL.n371 171.744
R182 VTAIL.n371 VTAIL.n327 171.744
R183 VTAIL.n364 VTAIL.n327 171.744
R184 VTAIL.n364 VTAIL.n363 171.744
R185 VTAIL.n363 VTAIL.n362 171.744
R186 VTAIL.n362 VTAIL.n331 171.744
R187 VTAIL.n355 VTAIL.n331 171.744
R188 VTAIL.n355 VTAIL.n354 171.744
R189 VTAIL.n354 VTAIL.n336 171.744
R190 VTAIL.n347 VTAIL.n336 171.744
R191 VTAIL.n347 VTAIL.n346 171.744
R192 VTAIL.n346 VTAIL.n340 171.744
R193 VTAIL.n318 VTAIL.n317 171.744
R194 VTAIL.n317 VTAIL.n273 171.744
R195 VTAIL.n310 VTAIL.n273 171.744
R196 VTAIL.n310 VTAIL.n309 171.744
R197 VTAIL.n309 VTAIL.n308 171.744
R198 VTAIL.n308 VTAIL.n277 171.744
R199 VTAIL.n301 VTAIL.n277 171.744
R200 VTAIL.n301 VTAIL.n300 171.744
R201 VTAIL.n300 VTAIL.n282 171.744
R202 VTAIL.n293 VTAIL.n282 171.744
R203 VTAIL.n293 VTAIL.n292 171.744
R204 VTAIL.n292 VTAIL.n286 171.744
R205 VTAIL.n264 VTAIL.n263 171.744
R206 VTAIL.n263 VTAIL.n219 171.744
R207 VTAIL.n256 VTAIL.n219 171.744
R208 VTAIL.n256 VTAIL.n255 171.744
R209 VTAIL.n255 VTAIL.n254 171.744
R210 VTAIL.n254 VTAIL.n223 171.744
R211 VTAIL.n247 VTAIL.n223 171.744
R212 VTAIL.n247 VTAIL.n246 171.744
R213 VTAIL.n246 VTAIL.n228 171.744
R214 VTAIL.n239 VTAIL.n228 171.744
R215 VTAIL.n239 VTAIL.n238 171.744
R216 VTAIL.n238 VTAIL.n232 171.744
R217 VTAIL.n210 VTAIL.n209 171.744
R218 VTAIL.n209 VTAIL.n165 171.744
R219 VTAIL.n202 VTAIL.n165 171.744
R220 VTAIL.n202 VTAIL.n201 171.744
R221 VTAIL.n201 VTAIL.n200 171.744
R222 VTAIL.n200 VTAIL.n169 171.744
R223 VTAIL.n193 VTAIL.n169 171.744
R224 VTAIL.n193 VTAIL.n192 171.744
R225 VTAIL.n192 VTAIL.n174 171.744
R226 VTAIL.n185 VTAIL.n174 171.744
R227 VTAIL.n185 VTAIL.n184 171.744
R228 VTAIL.n184 VTAIL.n178 171.744
R229 VTAIL.t1 VTAIL.n393 85.8723
R230 VTAIL.t4 VTAIL.n15 85.8723
R231 VTAIL.t6 VTAIL.n69 85.8723
R232 VTAIL.t5 VTAIL.n123 85.8723
R233 VTAIL.t0 VTAIL.n340 85.8723
R234 VTAIL.t7 VTAIL.n286 85.8723
R235 VTAIL.t3 VTAIL.n232 85.8723
R236 VTAIL.t2 VTAIL.n178 85.8723
R237 VTAIL.n431 VTAIL.n430 31.6035
R238 VTAIL.n53 VTAIL.n52 31.6035
R239 VTAIL.n107 VTAIL.n106 31.6035
R240 VTAIL.n161 VTAIL.n160 31.6035
R241 VTAIL.n377 VTAIL.n376 31.6035
R242 VTAIL.n323 VTAIL.n322 31.6035
R243 VTAIL.n269 VTAIL.n268 31.6035
R244 VTAIL.n215 VTAIL.n214 31.6035
R245 VTAIL.n431 VTAIL.n377 24.3152
R246 VTAIL.n215 VTAIL.n161 24.3152
R247 VTAIL.n419 VTAIL.n384 13.1884
R248 VTAIL.n41 VTAIL.n6 13.1884
R249 VTAIL.n95 VTAIL.n60 13.1884
R250 VTAIL.n149 VTAIL.n114 13.1884
R251 VTAIL.n365 VTAIL.n330 13.1884
R252 VTAIL.n311 VTAIL.n276 13.1884
R253 VTAIL.n257 VTAIL.n222 13.1884
R254 VTAIL.n203 VTAIL.n168 13.1884
R255 VTAIL.n415 VTAIL.n414 12.8005
R256 VTAIL.n420 VTAIL.n382 12.8005
R257 VTAIL.n37 VTAIL.n36 12.8005
R258 VTAIL.n42 VTAIL.n4 12.8005
R259 VTAIL.n91 VTAIL.n90 12.8005
R260 VTAIL.n96 VTAIL.n58 12.8005
R261 VTAIL.n145 VTAIL.n144 12.8005
R262 VTAIL.n150 VTAIL.n112 12.8005
R263 VTAIL.n366 VTAIL.n328 12.8005
R264 VTAIL.n361 VTAIL.n332 12.8005
R265 VTAIL.n312 VTAIL.n274 12.8005
R266 VTAIL.n307 VTAIL.n278 12.8005
R267 VTAIL.n258 VTAIL.n220 12.8005
R268 VTAIL.n253 VTAIL.n224 12.8005
R269 VTAIL.n204 VTAIL.n166 12.8005
R270 VTAIL.n199 VTAIL.n170 12.8005
R271 VTAIL.n413 VTAIL.n386 12.0247
R272 VTAIL.n424 VTAIL.n423 12.0247
R273 VTAIL.n35 VTAIL.n8 12.0247
R274 VTAIL.n46 VTAIL.n45 12.0247
R275 VTAIL.n89 VTAIL.n62 12.0247
R276 VTAIL.n100 VTAIL.n99 12.0247
R277 VTAIL.n143 VTAIL.n116 12.0247
R278 VTAIL.n154 VTAIL.n153 12.0247
R279 VTAIL.n370 VTAIL.n369 12.0247
R280 VTAIL.n360 VTAIL.n333 12.0247
R281 VTAIL.n316 VTAIL.n315 12.0247
R282 VTAIL.n306 VTAIL.n279 12.0247
R283 VTAIL.n262 VTAIL.n261 12.0247
R284 VTAIL.n252 VTAIL.n225 12.0247
R285 VTAIL.n208 VTAIL.n207 12.0247
R286 VTAIL.n198 VTAIL.n171 12.0247
R287 VTAIL.n410 VTAIL.n409 11.249
R288 VTAIL.n427 VTAIL.n380 11.249
R289 VTAIL.n32 VTAIL.n31 11.249
R290 VTAIL.n49 VTAIL.n2 11.249
R291 VTAIL.n86 VTAIL.n85 11.249
R292 VTAIL.n103 VTAIL.n56 11.249
R293 VTAIL.n140 VTAIL.n139 11.249
R294 VTAIL.n157 VTAIL.n110 11.249
R295 VTAIL.n373 VTAIL.n326 11.249
R296 VTAIL.n357 VTAIL.n356 11.249
R297 VTAIL.n319 VTAIL.n272 11.249
R298 VTAIL.n303 VTAIL.n302 11.249
R299 VTAIL.n265 VTAIL.n218 11.249
R300 VTAIL.n249 VTAIL.n248 11.249
R301 VTAIL.n211 VTAIL.n164 11.249
R302 VTAIL.n195 VTAIL.n194 11.249
R303 VTAIL.n395 VTAIL.n394 10.7239
R304 VTAIL.n17 VTAIL.n16 10.7239
R305 VTAIL.n71 VTAIL.n70 10.7239
R306 VTAIL.n125 VTAIL.n124 10.7239
R307 VTAIL.n342 VTAIL.n341 10.7239
R308 VTAIL.n288 VTAIL.n287 10.7239
R309 VTAIL.n234 VTAIL.n233 10.7239
R310 VTAIL.n180 VTAIL.n179 10.7239
R311 VTAIL.n406 VTAIL.n388 10.4732
R312 VTAIL.n428 VTAIL.n378 10.4732
R313 VTAIL.n28 VTAIL.n10 10.4732
R314 VTAIL.n50 VTAIL.n0 10.4732
R315 VTAIL.n82 VTAIL.n64 10.4732
R316 VTAIL.n104 VTAIL.n54 10.4732
R317 VTAIL.n136 VTAIL.n118 10.4732
R318 VTAIL.n158 VTAIL.n108 10.4732
R319 VTAIL.n374 VTAIL.n324 10.4732
R320 VTAIL.n353 VTAIL.n335 10.4732
R321 VTAIL.n320 VTAIL.n270 10.4732
R322 VTAIL.n299 VTAIL.n281 10.4732
R323 VTAIL.n266 VTAIL.n216 10.4732
R324 VTAIL.n245 VTAIL.n227 10.4732
R325 VTAIL.n212 VTAIL.n162 10.4732
R326 VTAIL.n191 VTAIL.n173 10.4732
R327 VTAIL.n405 VTAIL.n390 9.69747
R328 VTAIL.n27 VTAIL.n12 9.69747
R329 VTAIL.n81 VTAIL.n66 9.69747
R330 VTAIL.n135 VTAIL.n120 9.69747
R331 VTAIL.n352 VTAIL.n337 9.69747
R332 VTAIL.n298 VTAIL.n283 9.69747
R333 VTAIL.n244 VTAIL.n229 9.69747
R334 VTAIL.n190 VTAIL.n175 9.69747
R335 VTAIL.n430 VTAIL.n429 9.45567
R336 VTAIL.n52 VTAIL.n51 9.45567
R337 VTAIL.n106 VTAIL.n105 9.45567
R338 VTAIL.n160 VTAIL.n159 9.45567
R339 VTAIL.n376 VTAIL.n375 9.45567
R340 VTAIL.n322 VTAIL.n321 9.45567
R341 VTAIL.n268 VTAIL.n267 9.45567
R342 VTAIL.n214 VTAIL.n213 9.45567
R343 VTAIL.n429 VTAIL.n428 9.3005
R344 VTAIL.n380 VTAIL.n379 9.3005
R345 VTAIL.n423 VTAIL.n422 9.3005
R346 VTAIL.n421 VTAIL.n420 9.3005
R347 VTAIL.n397 VTAIL.n396 9.3005
R348 VTAIL.n392 VTAIL.n391 9.3005
R349 VTAIL.n403 VTAIL.n402 9.3005
R350 VTAIL.n405 VTAIL.n404 9.3005
R351 VTAIL.n388 VTAIL.n387 9.3005
R352 VTAIL.n411 VTAIL.n410 9.3005
R353 VTAIL.n413 VTAIL.n412 9.3005
R354 VTAIL.n414 VTAIL.n383 9.3005
R355 VTAIL.n51 VTAIL.n50 9.3005
R356 VTAIL.n2 VTAIL.n1 9.3005
R357 VTAIL.n45 VTAIL.n44 9.3005
R358 VTAIL.n43 VTAIL.n42 9.3005
R359 VTAIL.n19 VTAIL.n18 9.3005
R360 VTAIL.n14 VTAIL.n13 9.3005
R361 VTAIL.n25 VTAIL.n24 9.3005
R362 VTAIL.n27 VTAIL.n26 9.3005
R363 VTAIL.n10 VTAIL.n9 9.3005
R364 VTAIL.n33 VTAIL.n32 9.3005
R365 VTAIL.n35 VTAIL.n34 9.3005
R366 VTAIL.n36 VTAIL.n5 9.3005
R367 VTAIL.n105 VTAIL.n104 9.3005
R368 VTAIL.n56 VTAIL.n55 9.3005
R369 VTAIL.n99 VTAIL.n98 9.3005
R370 VTAIL.n97 VTAIL.n96 9.3005
R371 VTAIL.n73 VTAIL.n72 9.3005
R372 VTAIL.n68 VTAIL.n67 9.3005
R373 VTAIL.n79 VTAIL.n78 9.3005
R374 VTAIL.n81 VTAIL.n80 9.3005
R375 VTAIL.n64 VTAIL.n63 9.3005
R376 VTAIL.n87 VTAIL.n86 9.3005
R377 VTAIL.n89 VTAIL.n88 9.3005
R378 VTAIL.n90 VTAIL.n59 9.3005
R379 VTAIL.n159 VTAIL.n158 9.3005
R380 VTAIL.n110 VTAIL.n109 9.3005
R381 VTAIL.n153 VTAIL.n152 9.3005
R382 VTAIL.n151 VTAIL.n150 9.3005
R383 VTAIL.n127 VTAIL.n126 9.3005
R384 VTAIL.n122 VTAIL.n121 9.3005
R385 VTAIL.n133 VTAIL.n132 9.3005
R386 VTAIL.n135 VTAIL.n134 9.3005
R387 VTAIL.n118 VTAIL.n117 9.3005
R388 VTAIL.n141 VTAIL.n140 9.3005
R389 VTAIL.n143 VTAIL.n142 9.3005
R390 VTAIL.n144 VTAIL.n113 9.3005
R391 VTAIL.n344 VTAIL.n343 9.3005
R392 VTAIL.n339 VTAIL.n338 9.3005
R393 VTAIL.n350 VTAIL.n349 9.3005
R394 VTAIL.n352 VTAIL.n351 9.3005
R395 VTAIL.n335 VTAIL.n334 9.3005
R396 VTAIL.n358 VTAIL.n357 9.3005
R397 VTAIL.n360 VTAIL.n359 9.3005
R398 VTAIL.n332 VTAIL.n329 9.3005
R399 VTAIL.n375 VTAIL.n374 9.3005
R400 VTAIL.n326 VTAIL.n325 9.3005
R401 VTAIL.n369 VTAIL.n368 9.3005
R402 VTAIL.n367 VTAIL.n366 9.3005
R403 VTAIL.n290 VTAIL.n289 9.3005
R404 VTAIL.n285 VTAIL.n284 9.3005
R405 VTAIL.n296 VTAIL.n295 9.3005
R406 VTAIL.n298 VTAIL.n297 9.3005
R407 VTAIL.n281 VTAIL.n280 9.3005
R408 VTAIL.n304 VTAIL.n303 9.3005
R409 VTAIL.n306 VTAIL.n305 9.3005
R410 VTAIL.n278 VTAIL.n275 9.3005
R411 VTAIL.n321 VTAIL.n320 9.3005
R412 VTAIL.n272 VTAIL.n271 9.3005
R413 VTAIL.n315 VTAIL.n314 9.3005
R414 VTAIL.n313 VTAIL.n312 9.3005
R415 VTAIL.n236 VTAIL.n235 9.3005
R416 VTAIL.n231 VTAIL.n230 9.3005
R417 VTAIL.n242 VTAIL.n241 9.3005
R418 VTAIL.n244 VTAIL.n243 9.3005
R419 VTAIL.n227 VTAIL.n226 9.3005
R420 VTAIL.n250 VTAIL.n249 9.3005
R421 VTAIL.n252 VTAIL.n251 9.3005
R422 VTAIL.n224 VTAIL.n221 9.3005
R423 VTAIL.n267 VTAIL.n266 9.3005
R424 VTAIL.n218 VTAIL.n217 9.3005
R425 VTAIL.n261 VTAIL.n260 9.3005
R426 VTAIL.n259 VTAIL.n258 9.3005
R427 VTAIL.n182 VTAIL.n181 9.3005
R428 VTAIL.n177 VTAIL.n176 9.3005
R429 VTAIL.n188 VTAIL.n187 9.3005
R430 VTAIL.n190 VTAIL.n189 9.3005
R431 VTAIL.n173 VTAIL.n172 9.3005
R432 VTAIL.n196 VTAIL.n195 9.3005
R433 VTAIL.n198 VTAIL.n197 9.3005
R434 VTAIL.n170 VTAIL.n167 9.3005
R435 VTAIL.n213 VTAIL.n212 9.3005
R436 VTAIL.n164 VTAIL.n163 9.3005
R437 VTAIL.n207 VTAIL.n206 9.3005
R438 VTAIL.n205 VTAIL.n204 9.3005
R439 VTAIL.n402 VTAIL.n401 8.92171
R440 VTAIL.n24 VTAIL.n23 8.92171
R441 VTAIL.n78 VTAIL.n77 8.92171
R442 VTAIL.n132 VTAIL.n131 8.92171
R443 VTAIL.n349 VTAIL.n348 8.92171
R444 VTAIL.n295 VTAIL.n294 8.92171
R445 VTAIL.n241 VTAIL.n240 8.92171
R446 VTAIL.n187 VTAIL.n186 8.92171
R447 VTAIL.n398 VTAIL.n392 8.14595
R448 VTAIL.n20 VTAIL.n14 8.14595
R449 VTAIL.n74 VTAIL.n68 8.14595
R450 VTAIL.n128 VTAIL.n122 8.14595
R451 VTAIL.n345 VTAIL.n339 8.14595
R452 VTAIL.n291 VTAIL.n285 8.14595
R453 VTAIL.n237 VTAIL.n231 8.14595
R454 VTAIL.n183 VTAIL.n177 8.14595
R455 VTAIL.n397 VTAIL.n394 7.3702
R456 VTAIL.n19 VTAIL.n16 7.3702
R457 VTAIL.n73 VTAIL.n70 7.3702
R458 VTAIL.n127 VTAIL.n124 7.3702
R459 VTAIL.n344 VTAIL.n341 7.3702
R460 VTAIL.n290 VTAIL.n287 7.3702
R461 VTAIL.n236 VTAIL.n233 7.3702
R462 VTAIL.n182 VTAIL.n179 7.3702
R463 VTAIL.n398 VTAIL.n397 5.81868
R464 VTAIL.n20 VTAIL.n19 5.81868
R465 VTAIL.n74 VTAIL.n73 5.81868
R466 VTAIL.n128 VTAIL.n127 5.81868
R467 VTAIL.n345 VTAIL.n344 5.81868
R468 VTAIL.n291 VTAIL.n290 5.81868
R469 VTAIL.n237 VTAIL.n236 5.81868
R470 VTAIL.n183 VTAIL.n182 5.81868
R471 VTAIL.n401 VTAIL.n392 5.04292
R472 VTAIL.n23 VTAIL.n14 5.04292
R473 VTAIL.n77 VTAIL.n68 5.04292
R474 VTAIL.n131 VTAIL.n122 5.04292
R475 VTAIL.n348 VTAIL.n339 5.04292
R476 VTAIL.n294 VTAIL.n285 5.04292
R477 VTAIL.n240 VTAIL.n231 5.04292
R478 VTAIL.n186 VTAIL.n177 5.04292
R479 VTAIL.n402 VTAIL.n390 4.26717
R480 VTAIL.n24 VTAIL.n12 4.26717
R481 VTAIL.n78 VTAIL.n66 4.26717
R482 VTAIL.n132 VTAIL.n120 4.26717
R483 VTAIL.n349 VTAIL.n337 4.26717
R484 VTAIL.n295 VTAIL.n283 4.26717
R485 VTAIL.n241 VTAIL.n229 4.26717
R486 VTAIL.n187 VTAIL.n175 4.26717
R487 VTAIL.n406 VTAIL.n405 3.49141
R488 VTAIL.n430 VTAIL.n378 3.49141
R489 VTAIL.n28 VTAIL.n27 3.49141
R490 VTAIL.n52 VTAIL.n0 3.49141
R491 VTAIL.n82 VTAIL.n81 3.49141
R492 VTAIL.n106 VTAIL.n54 3.49141
R493 VTAIL.n136 VTAIL.n135 3.49141
R494 VTAIL.n160 VTAIL.n108 3.49141
R495 VTAIL.n376 VTAIL.n324 3.49141
R496 VTAIL.n353 VTAIL.n352 3.49141
R497 VTAIL.n322 VTAIL.n270 3.49141
R498 VTAIL.n299 VTAIL.n298 3.49141
R499 VTAIL.n268 VTAIL.n216 3.49141
R500 VTAIL.n245 VTAIL.n244 3.49141
R501 VTAIL.n214 VTAIL.n162 3.49141
R502 VTAIL.n191 VTAIL.n190 3.49141
R503 VTAIL.n269 VTAIL.n215 3.38843
R504 VTAIL.n377 VTAIL.n323 3.38843
R505 VTAIL.n161 VTAIL.n107 3.38843
R506 VTAIL.n409 VTAIL.n388 2.71565
R507 VTAIL.n428 VTAIL.n427 2.71565
R508 VTAIL.n31 VTAIL.n10 2.71565
R509 VTAIL.n50 VTAIL.n49 2.71565
R510 VTAIL.n85 VTAIL.n64 2.71565
R511 VTAIL.n104 VTAIL.n103 2.71565
R512 VTAIL.n139 VTAIL.n118 2.71565
R513 VTAIL.n158 VTAIL.n157 2.71565
R514 VTAIL.n374 VTAIL.n373 2.71565
R515 VTAIL.n356 VTAIL.n335 2.71565
R516 VTAIL.n320 VTAIL.n319 2.71565
R517 VTAIL.n302 VTAIL.n281 2.71565
R518 VTAIL.n266 VTAIL.n265 2.71565
R519 VTAIL.n248 VTAIL.n227 2.71565
R520 VTAIL.n212 VTAIL.n211 2.71565
R521 VTAIL.n194 VTAIL.n173 2.71565
R522 VTAIL.n396 VTAIL.n395 2.41283
R523 VTAIL.n18 VTAIL.n17 2.41283
R524 VTAIL.n72 VTAIL.n71 2.41283
R525 VTAIL.n126 VTAIL.n125 2.41283
R526 VTAIL.n343 VTAIL.n342 2.41283
R527 VTAIL.n289 VTAIL.n288 2.41283
R528 VTAIL.n235 VTAIL.n234 2.41283
R529 VTAIL.n181 VTAIL.n180 2.41283
R530 VTAIL.n410 VTAIL.n386 1.93989
R531 VTAIL.n424 VTAIL.n380 1.93989
R532 VTAIL.n32 VTAIL.n8 1.93989
R533 VTAIL.n46 VTAIL.n2 1.93989
R534 VTAIL.n86 VTAIL.n62 1.93989
R535 VTAIL.n100 VTAIL.n56 1.93989
R536 VTAIL.n140 VTAIL.n116 1.93989
R537 VTAIL.n154 VTAIL.n110 1.93989
R538 VTAIL.n370 VTAIL.n326 1.93989
R539 VTAIL.n357 VTAIL.n333 1.93989
R540 VTAIL.n316 VTAIL.n272 1.93989
R541 VTAIL.n303 VTAIL.n279 1.93989
R542 VTAIL.n262 VTAIL.n218 1.93989
R543 VTAIL.n249 VTAIL.n225 1.93989
R544 VTAIL.n208 VTAIL.n164 1.93989
R545 VTAIL.n195 VTAIL.n171 1.93989
R546 VTAIL VTAIL.n53 1.75266
R547 VTAIL VTAIL.n431 1.63628
R548 VTAIL.n415 VTAIL.n413 1.16414
R549 VTAIL.n423 VTAIL.n382 1.16414
R550 VTAIL.n37 VTAIL.n35 1.16414
R551 VTAIL.n45 VTAIL.n4 1.16414
R552 VTAIL.n91 VTAIL.n89 1.16414
R553 VTAIL.n99 VTAIL.n58 1.16414
R554 VTAIL.n145 VTAIL.n143 1.16414
R555 VTAIL.n153 VTAIL.n112 1.16414
R556 VTAIL.n369 VTAIL.n328 1.16414
R557 VTAIL.n361 VTAIL.n360 1.16414
R558 VTAIL.n315 VTAIL.n274 1.16414
R559 VTAIL.n307 VTAIL.n306 1.16414
R560 VTAIL.n261 VTAIL.n220 1.16414
R561 VTAIL.n253 VTAIL.n252 1.16414
R562 VTAIL.n207 VTAIL.n166 1.16414
R563 VTAIL.n199 VTAIL.n198 1.16414
R564 VTAIL.n323 VTAIL.n269 0.470328
R565 VTAIL.n107 VTAIL.n53 0.470328
R566 VTAIL.n414 VTAIL.n384 0.388379
R567 VTAIL.n420 VTAIL.n419 0.388379
R568 VTAIL.n36 VTAIL.n6 0.388379
R569 VTAIL.n42 VTAIL.n41 0.388379
R570 VTAIL.n90 VTAIL.n60 0.388379
R571 VTAIL.n96 VTAIL.n95 0.388379
R572 VTAIL.n144 VTAIL.n114 0.388379
R573 VTAIL.n150 VTAIL.n149 0.388379
R574 VTAIL.n366 VTAIL.n365 0.388379
R575 VTAIL.n332 VTAIL.n330 0.388379
R576 VTAIL.n312 VTAIL.n311 0.388379
R577 VTAIL.n278 VTAIL.n276 0.388379
R578 VTAIL.n258 VTAIL.n257 0.388379
R579 VTAIL.n224 VTAIL.n222 0.388379
R580 VTAIL.n204 VTAIL.n203 0.388379
R581 VTAIL.n170 VTAIL.n168 0.388379
R582 VTAIL.n396 VTAIL.n391 0.155672
R583 VTAIL.n403 VTAIL.n391 0.155672
R584 VTAIL.n404 VTAIL.n403 0.155672
R585 VTAIL.n404 VTAIL.n387 0.155672
R586 VTAIL.n411 VTAIL.n387 0.155672
R587 VTAIL.n412 VTAIL.n411 0.155672
R588 VTAIL.n412 VTAIL.n383 0.155672
R589 VTAIL.n421 VTAIL.n383 0.155672
R590 VTAIL.n422 VTAIL.n421 0.155672
R591 VTAIL.n422 VTAIL.n379 0.155672
R592 VTAIL.n429 VTAIL.n379 0.155672
R593 VTAIL.n18 VTAIL.n13 0.155672
R594 VTAIL.n25 VTAIL.n13 0.155672
R595 VTAIL.n26 VTAIL.n25 0.155672
R596 VTAIL.n26 VTAIL.n9 0.155672
R597 VTAIL.n33 VTAIL.n9 0.155672
R598 VTAIL.n34 VTAIL.n33 0.155672
R599 VTAIL.n34 VTAIL.n5 0.155672
R600 VTAIL.n43 VTAIL.n5 0.155672
R601 VTAIL.n44 VTAIL.n43 0.155672
R602 VTAIL.n44 VTAIL.n1 0.155672
R603 VTAIL.n51 VTAIL.n1 0.155672
R604 VTAIL.n72 VTAIL.n67 0.155672
R605 VTAIL.n79 VTAIL.n67 0.155672
R606 VTAIL.n80 VTAIL.n79 0.155672
R607 VTAIL.n80 VTAIL.n63 0.155672
R608 VTAIL.n87 VTAIL.n63 0.155672
R609 VTAIL.n88 VTAIL.n87 0.155672
R610 VTAIL.n88 VTAIL.n59 0.155672
R611 VTAIL.n97 VTAIL.n59 0.155672
R612 VTAIL.n98 VTAIL.n97 0.155672
R613 VTAIL.n98 VTAIL.n55 0.155672
R614 VTAIL.n105 VTAIL.n55 0.155672
R615 VTAIL.n126 VTAIL.n121 0.155672
R616 VTAIL.n133 VTAIL.n121 0.155672
R617 VTAIL.n134 VTAIL.n133 0.155672
R618 VTAIL.n134 VTAIL.n117 0.155672
R619 VTAIL.n141 VTAIL.n117 0.155672
R620 VTAIL.n142 VTAIL.n141 0.155672
R621 VTAIL.n142 VTAIL.n113 0.155672
R622 VTAIL.n151 VTAIL.n113 0.155672
R623 VTAIL.n152 VTAIL.n151 0.155672
R624 VTAIL.n152 VTAIL.n109 0.155672
R625 VTAIL.n159 VTAIL.n109 0.155672
R626 VTAIL.n375 VTAIL.n325 0.155672
R627 VTAIL.n368 VTAIL.n325 0.155672
R628 VTAIL.n368 VTAIL.n367 0.155672
R629 VTAIL.n367 VTAIL.n329 0.155672
R630 VTAIL.n359 VTAIL.n329 0.155672
R631 VTAIL.n359 VTAIL.n358 0.155672
R632 VTAIL.n358 VTAIL.n334 0.155672
R633 VTAIL.n351 VTAIL.n334 0.155672
R634 VTAIL.n351 VTAIL.n350 0.155672
R635 VTAIL.n350 VTAIL.n338 0.155672
R636 VTAIL.n343 VTAIL.n338 0.155672
R637 VTAIL.n321 VTAIL.n271 0.155672
R638 VTAIL.n314 VTAIL.n271 0.155672
R639 VTAIL.n314 VTAIL.n313 0.155672
R640 VTAIL.n313 VTAIL.n275 0.155672
R641 VTAIL.n305 VTAIL.n275 0.155672
R642 VTAIL.n305 VTAIL.n304 0.155672
R643 VTAIL.n304 VTAIL.n280 0.155672
R644 VTAIL.n297 VTAIL.n280 0.155672
R645 VTAIL.n297 VTAIL.n296 0.155672
R646 VTAIL.n296 VTAIL.n284 0.155672
R647 VTAIL.n289 VTAIL.n284 0.155672
R648 VTAIL.n267 VTAIL.n217 0.155672
R649 VTAIL.n260 VTAIL.n217 0.155672
R650 VTAIL.n260 VTAIL.n259 0.155672
R651 VTAIL.n259 VTAIL.n221 0.155672
R652 VTAIL.n251 VTAIL.n221 0.155672
R653 VTAIL.n251 VTAIL.n250 0.155672
R654 VTAIL.n250 VTAIL.n226 0.155672
R655 VTAIL.n243 VTAIL.n226 0.155672
R656 VTAIL.n243 VTAIL.n242 0.155672
R657 VTAIL.n242 VTAIL.n230 0.155672
R658 VTAIL.n235 VTAIL.n230 0.155672
R659 VTAIL.n213 VTAIL.n163 0.155672
R660 VTAIL.n206 VTAIL.n163 0.155672
R661 VTAIL.n206 VTAIL.n205 0.155672
R662 VTAIL.n205 VTAIL.n167 0.155672
R663 VTAIL.n197 VTAIL.n167 0.155672
R664 VTAIL.n197 VTAIL.n196 0.155672
R665 VTAIL.n196 VTAIL.n172 0.155672
R666 VTAIL.n189 VTAIL.n172 0.155672
R667 VTAIL.n189 VTAIL.n188 0.155672
R668 VTAIL.n188 VTAIL.n176 0.155672
R669 VTAIL.n181 VTAIL.n176 0.155672
R670 B.n495 B.n68 585
R671 B.n497 B.n496 585
R672 B.n498 B.n67 585
R673 B.n500 B.n499 585
R674 B.n501 B.n66 585
R675 B.n503 B.n502 585
R676 B.n504 B.n65 585
R677 B.n506 B.n505 585
R678 B.n507 B.n64 585
R679 B.n509 B.n508 585
R680 B.n510 B.n63 585
R681 B.n512 B.n511 585
R682 B.n513 B.n62 585
R683 B.n515 B.n514 585
R684 B.n516 B.n61 585
R685 B.n518 B.n517 585
R686 B.n519 B.n60 585
R687 B.n521 B.n520 585
R688 B.n522 B.n59 585
R689 B.n524 B.n523 585
R690 B.n525 B.n58 585
R691 B.n527 B.n526 585
R692 B.n528 B.n57 585
R693 B.n530 B.n529 585
R694 B.n531 B.n56 585
R695 B.n533 B.n532 585
R696 B.n534 B.n55 585
R697 B.n536 B.n535 585
R698 B.n537 B.n54 585
R699 B.n539 B.n538 585
R700 B.n540 B.n53 585
R701 B.n542 B.n541 585
R702 B.n543 B.n52 585
R703 B.n545 B.n544 585
R704 B.n546 B.n51 585
R705 B.n548 B.n547 585
R706 B.n550 B.n549 585
R707 B.n551 B.n47 585
R708 B.n553 B.n552 585
R709 B.n554 B.n46 585
R710 B.n556 B.n555 585
R711 B.n557 B.n45 585
R712 B.n559 B.n558 585
R713 B.n560 B.n44 585
R714 B.n562 B.n561 585
R715 B.n564 B.n41 585
R716 B.n566 B.n565 585
R717 B.n567 B.n40 585
R718 B.n569 B.n568 585
R719 B.n570 B.n39 585
R720 B.n572 B.n571 585
R721 B.n573 B.n38 585
R722 B.n575 B.n574 585
R723 B.n576 B.n37 585
R724 B.n578 B.n577 585
R725 B.n579 B.n36 585
R726 B.n581 B.n580 585
R727 B.n582 B.n35 585
R728 B.n584 B.n583 585
R729 B.n585 B.n34 585
R730 B.n587 B.n586 585
R731 B.n588 B.n33 585
R732 B.n590 B.n589 585
R733 B.n591 B.n32 585
R734 B.n593 B.n592 585
R735 B.n594 B.n31 585
R736 B.n596 B.n595 585
R737 B.n597 B.n30 585
R738 B.n599 B.n598 585
R739 B.n600 B.n29 585
R740 B.n602 B.n601 585
R741 B.n603 B.n28 585
R742 B.n605 B.n604 585
R743 B.n606 B.n27 585
R744 B.n608 B.n607 585
R745 B.n609 B.n26 585
R746 B.n611 B.n610 585
R747 B.n612 B.n25 585
R748 B.n614 B.n613 585
R749 B.n615 B.n24 585
R750 B.n617 B.n616 585
R751 B.n494 B.n493 585
R752 B.n492 B.n69 585
R753 B.n491 B.n490 585
R754 B.n489 B.n70 585
R755 B.n488 B.n487 585
R756 B.n486 B.n71 585
R757 B.n485 B.n484 585
R758 B.n483 B.n72 585
R759 B.n482 B.n481 585
R760 B.n480 B.n73 585
R761 B.n479 B.n478 585
R762 B.n477 B.n74 585
R763 B.n476 B.n475 585
R764 B.n474 B.n75 585
R765 B.n473 B.n472 585
R766 B.n471 B.n76 585
R767 B.n470 B.n469 585
R768 B.n468 B.n77 585
R769 B.n467 B.n466 585
R770 B.n465 B.n78 585
R771 B.n464 B.n463 585
R772 B.n462 B.n79 585
R773 B.n461 B.n460 585
R774 B.n459 B.n80 585
R775 B.n458 B.n457 585
R776 B.n456 B.n81 585
R777 B.n455 B.n454 585
R778 B.n453 B.n82 585
R779 B.n452 B.n451 585
R780 B.n450 B.n83 585
R781 B.n449 B.n448 585
R782 B.n447 B.n84 585
R783 B.n446 B.n445 585
R784 B.n444 B.n85 585
R785 B.n443 B.n442 585
R786 B.n441 B.n86 585
R787 B.n440 B.n439 585
R788 B.n438 B.n87 585
R789 B.n437 B.n436 585
R790 B.n435 B.n88 585
R791 B.n434 B.n433 585
R792 B.n432 B.n89 585
R793 B.n431 B.n430 585
R794 B.n429 B.n90 585
R795 B.n428 B.n427 585
R796 B.n426 B.n91 585
R797 B.n425 B.n424 585
R798 B.n423 B.n92 585
R799 B.n422 B.n421 585
R800 B.n420 B.n93 585
R801 B.n419 B.n418 585
R802 B.n417 B.n94 585
R803 B.n416 B.n415 585
R804 B.n414 B.n95 585
R805 B.n413 B.n412 585
R806 B.n411 B.n96 585
R807 B.n410 B.n409 585
R808 B.n408 B.n97 585
R809 B.n407 B.n406 585
R810 B.n405 B.n98 585
R811 B.n404 B.n403 585
R812 B.n402 B.n99 585
R813 B.n401 B.n400 585
R814 B.n399 B.n100 585
R815 B.n398 B.n397 585
R816 B.n396 B.n101 585
R817 B.n395 B.n394 585
R818 B.n393 B.n102 585
R819 B.n392 B.n391 585
R820 B.n390 B.n103 585
R821 B.n389 B.n388 585
R822 B.n387 B.n104 585
R823 B.n386 B.n385 585
R824 B.n384 B.n105 585
R825 B.n383 B.n382 585
R826 B.n381 B.n106 585
R827 B.n380 B.n379 585
R828 B.n378 B.n107 585
R829 B.n377 B.n376 585
R830 B.n375 B.n108 585
R831 B.n374 B.n373 585
R832 B.n372 B.n109 585
R833 B.n371 B.n370 585
R834 B.n369 B.n110 585
R835 B.n368 B.n367 585
R836 B.n366 B.n111 585
R837 B.n365 B.n364 585
R838 B.n242 B.n241 585
R839 B.n243 B.n156 585
R840 B.n245 B.n244 585
R841 B.n246 B.n155 585
R842 B.n248 B.n247 585
R843 B.n249 B.n154 585
R844 B.n251 B.n250 585
R845 B.n252 B.n153 585
R846 B.n254 B.n253 585
R847 B.n255 B.n152 585
R848 B.n257 B.n256 585
R849 B.n258 B.n151 585
R850 B.n260 B.n259 585
R851 B.n261 B.n150 585
R852 B.n263 B.n262 585
R853 B.n264 B.n149 585
R854 B.n266 B.n265 585
R855 B.n267 B.n148 585
R856 B.n269 B.n268 585
R857 B.n270 B.n147 585
R858 B.n272 B.n271 585
R859 B.n273 B.n146 585
R860 B.n275 B.n274 585
R861 B.n276 B.n145 585
R862 B.n278 B.n277 585
R863 B.n279 B.n144 585
R864 B.n281 B.n280 585
R865 B.n282 B.n143 585
R866 B.n284 B.n283 585
R867 B.n285 B.n142 585
R868 B.n287 B.n286 585
R869 B.n288 B.n141 585
R870 B.n290 B.n289 585
R871 B.n291 B.n140 585
R872 B.n293 B.n292 585
R873 B.n294 B.n137 585
R874 B.n297 B.n296 585
R875 B.n298 B.n136 585
R876 B.n300 B.n299 585
R877 B.n301 B.n135 585
R878 B.n303 B.n302 585
R879 B.n304 B.n134 585
R880 B.n306 B.n305 585
R881 B.n307 B.n133 585
R882 B.n309 B.n308 585
R883 B.n311 B.n310 585
R884 B.n312 B.n129 585
R885 B.n314 B.n313 585
R886 B.n315 B.n128 585
R887 B.n317 B.n316 585
R888 B.n318 B.n127 585
R889 B.n320 B.n319 585
R890 B.n321 B.n126 585
R891 B.n323 B.n322 585
R892 B.n324 B.n125 585
R893 B.n326 B.n325 585
R894 B.n327 B.n124 585
R895 B.n329 B.n328 585
R896 B.n330 B.n123 585
R897 B.n332 B.n331 585
R898 B.n333 B.n122 585
R899 B.n335 B.n334 585
R900 B.n336 B.n121 585
R901 B.n338 B.n337 585
R902 B.n339 B.n120 585
R903 B.n341 B.n340 585
R904 B.n342 B.n119 585
R905 B.n344 B.n343 585
R906 B.n345 B.n118 585
R907 B.n347 B.n346 585
R908 B.n348 B.n117 585
R909 B.n350 B.n349 585
R910 B.n351 B.n116 585
R911 B.n353 B.n352 585
R912 B.n354 B.n115 585
R913 B.n356 B.n355 585
R914 B.n357 B.n114 585
R915 B.n359 B.n358 585
R916 B.n360 B.n113 585
R917 B.n362 B.n361 585
R918 B.n363 B.n112 585
R919 B.n240 B.n157 585
R920 B.n239 B.n238 585
R921 B.n237 B.n158 585
R922 B.n236 B.n235 585
R923 B.n234 B.n159 585
R924 B.n233 B.n232 585
R925 B.n231 B.n160 585
R926 B.n230 B.n229 585
R927 B.n228 B.n161 585
R928 B.n227 B.n226 585
R929 B.n225 B.n162 585
R930 B.n224 B.n223 585
R931 B.n222 B.n163 585
R932 B.n221 B.n220 585
R933 B.n219 B.n164 585
R934 B.n218 B.n217 585
R935 B.n216 B.n165 585
R936 B.n215 B.n214 585
R937 B.n213 B.n166 585
R938 B.n212 B.n211 585
R939 B.n210 B.n167 585
R940 B.n209 B.n208 585
R941 B.n207 B.n168 585
R942 B.n206 B.n205 585
R943 B.n204 B.n169 585
R944 B.n203 B.n202 585
R945 B.n201 B.n170 585
R946 B.n200 B.n199 585
R947 B.n198 B.n171 585
R948 B.n197 B.n196 585
R949 B.n195 B.n172 585
R950 B.n194 B.n193 585
R951 B.n192 B.n173 585
R952 B.n191 B.n190 585
R953 B.n189 B.n174 585
R954 B.n188 B.n187 585
R955 B.n186 B.n175 585
R956 B.n185 B.n184 585
R957 B.n183 B.n176 585
R958 B.n182 B.n181 585
R959 B.n180 B.n177 585
R960 B.n179 B.n178 585
R961 B.n2 B.n0 585
R962 B.n681 B.n1 585
R963 B.n680 B.n679 585
R964 B.n678 B.n3 585
R965 B.n677 B.n676 585
R966 B.n675 B.n4 585
R967 B.n674 B.n673 585
R968 B.n672 B.n5 585
R969 B.n671 B.n670 585
R970 B.n669 B.n6 585
R971 B.n668 B.n667 585
R972 B.n666 B.n7 585
R973 B.n665 B.n664 585
R974 B.n663 B.n8 585
R975 B.n662 B.n661 585
R976 B.n660 B.n9 585
R977 B.n659 B.n658 585
R978 B.n657 B.n10 585
R979 B.n656 B.n655 585
R980 B.n654 B.n11 585
R981 B.n653 B.n652 585
R982 B.n651 B.n12 585
R983 B.n650 B.n649 585
R984 B.n648 B.n13 585
R985 B.n647 B.n646 585
R986 B.n645 B.n14 585
R987 B.n644 B.n643 585
R988 B.n642 B.n15 585
R989 B.n641 B.n640 585
R990 B.n639 B.n16 585
R991 B.n638 B.n637 585
R992 B.n636 B.n17 585
R993 B.n635 B.n634 585
R994 B.n633 B.n18 585
R995 B.n632 B.n631 585
R996 B.n630 B.n19 585
R997 B.n629 B.n628 585
R998 B.n627 B.n20 585
R999 B.n626 B.n625 585
R1000 B.n624 B.n21 585
R1001 B.n623 B.n622 585
R1002 B.n621 B.n22 585
R1003 B.n620 B.n619 585
R1004 B.n618 B.n23 585
R1005 B.n683 B.n682 585
R1006 B.n242 B.n157 434.841
R1007 B.n616 B.n23 434.841
R1008 B.n364 B.n363 434.841
R1009 B.n495 B.n494 434.841
R1010 B.n130 B.t8 414.437
R1011 B.n48 B.t1 414.437
R1012 B.n138 B.t5 414.437
R1013 B.n42 B.t10 414.437
R1014 B.n131 B.t7 338.219
R1015 B.n49 B.t2 338.219
R1016 B.n139 B.t4 338.219
R1017 B.n43 B.t11 338.219
R1018 B.n130 B.t6 275.658
R1019 B.n138 B.t3 275.658
R1020 B.n42 B.t9 275.658
R1021 B.n48 B.t0 275.658
R1022 B.n238 B.n157 163.367
R1023 B.n238 B.n237 163.367
R1024 B.n237 B.n236 163.367
R1025 B.n236 B.n159 163.367
R1026 B.n232 B.n159 163.367
R1027 B.n232 B.n231 163.367
R1028 B.n231 B.n230 163.367
R1029 B.n230 B.n161 163.367
R1030 B.n226 B.n161 163.367
R1031 B.n226 B.n225 163.367
R1032 B.n225 B.n224 163.367
R1033 B.n224 B.n163 163.367
R1034 B.n220 B.n163 163.367
R1035 B.n220 B.n219 163.367
R1036 B.n219 B.n218 163.367
R1037 B.n218 B.n165 163.367
R1038 B.n214 B.n165 163.367
R1039 B.n214 B.n213 163.367
R1040 B.n213 B.n212 163.367
R1041 B.n212 B.n167 163.367
R1042 B.n208 B.n167 163.367
R1043 B.n208 B.n207 163.367
R1044 B.n207 B.n206 163.367
R1045 B.n206 B.n169 163.367
R1046 B.n202 B.n169 163.367
R1047 B.n202 B.n201 163.367
R1048 B.n201 B.n200 163.367
R1049 B.n200 B.n171 163.367
R1050 B.n196 B.n171 163.367
R1051 B.n196 B.n195 163.367
R1052 B.n195 B.n194 163.367
R1053 B.n194 B.n173 163.367
R1054 B.n190 B.n173 163.367
R1055 B.n190 B.n189 163.367
R1056 B.n189 B.n188 163.367
R1057 B.n188 B.n175 163.367
R1058 B.n184 B.n175 163.367
R1059 B.n184 B.n183 163.367
R1060 B.n183 B.n182 163.367
R1061 B.n182 B.n177 163.367
R1062 B.n178 B.n177 163.367
R1063 B.n178 B.n2 163.367
R1064 B.n682 B.n2 163.367
R1065 B.n682 B.n681 163.367
R1066 B.n681 B.n680 163.367
R1067 B.n680 B.n3 163.367
R1068 B.n676 B.n3 163.367
R1069 B.n676 B.n675 163.367
R1070 B.n675 B.n674 163.367
R1071 B.n674 B.n5 163.367
R1072 B.n670 B.n5 163.367
R1073 B.n670 B.n669 163.367
R1074 B.n669 B.n668 163.367
R1075 B.n668 B.n7 163.367
R1076 B.n664 B.n7 163.367
R1077 B.n664 B.n663 163.367
R1078 B.n663 B.n662 163.367
R1079 B.n662 B.n9 163.367
R1080 B.n658 B.n9 163.367
R1081 B.n658 B.n657 163.367
R1082 B.n657 B.n656 163.367
R1083 B.n656 B.n11 163.367
R1084 B.n652 B.n11 163.367
R1085 B.n652 B.n651 163.367
R1086 B.n651 B.n650 163.367
R1087 B.n650 B.n13 163.367
R1088 B.n646 B.n13 163.367
R1089 B.n646 B.n645 163.367
R1090 B.n645 B.n644 163.367
R1091 B.n644 B.n15 163.367
R1092 B.n640 B.n15 163.367
R1093 B.n640 B.n639 163.367
R1094 B.n639 B.n638 163.367
R1095 B.n638 B.n17 163.367
R1096 B.n634 B.n17 163.367
R1097 B.n634 B.n633 163.367
R1098 B.n633 B.n632 163.367
R1099 B.n632 B.n19 163.367
R1100 B.n628 B.n19 163.367
R1101 B.n628 B.n627 163.367
R1102 B.n627 B.n626 163.367
R1103 B.n626 B.n21 163.367
R1104 B.n622 B.n21 163.367
R1105 B.n622 B.n621 163.367
R1106 B.n621 B.n620 163.367
R1107 B.n620 B.n23 163.367
R1108 B.n243 B.n242 163.367
R1109 B.n244 B.n243 163.367
R1110 B.n244 B.n155 163.367
R1111 B.n248 B.n155 163.367
R1112 B.n249 B.n248 163.367
R1113 B.n250 B.n249 163.367
R1114 B.n250 B.n153 163.367
R1115 B.n254 B.n153 163.367
R1116 B.n255 B.n254 163.367
R1117 B.n256 B.n255 163.367
R1118 B.n256 B.n151 163.367
R1119 B.n260 B.n151 163.367
R1120 B.n261 B.n260 163.367
R1121 B.n262 B.n261 163.367
R1122 B.n262 B.n149 163.367
R1123 B.n266 B.n149 163.367
R1124 B.n267 B.n266 163.367
R1125 B.n268 B.n267 163.367
R1126 B.n268 B.n147 163.367
R1127 B.n272 B.n147 163.367
R1128 B.n273 B.n272 163.367
R1129 B.n274 B.n273 163.367
R1130 B.n274 B.n145 163.367
R1131 B.n278 B.n145 163.367
R1132 B.n279 B.n278 163.367
R1133 B.n280 B.n279 163.367
R1134 B.n280 B.n143 163.367
R1135 B.n284 B.n143 163.367
R1136 B.n285 B.n284 163.367
R1137 B.n286 B.n285 163.367
R1138 B.n286 B.n141 163.367
R1139 B.n290 B.n141 163.367
R1140 B.n291 B.n290 163.367
R1141 B.n292 B.n291 163.367
R1142 B.n292 B.n137 163.367
R1143 B.n297 B.n137 163.367
R1144 B.n298 B.n297 163.367
R1145 B.n299 B.n298 163.367
R1146 B.n299 B.n135 163.367
R1147 B.n303 B.n135 163.367
R1148 B.n304 B.n303 163.367
R1149 B.n305 B.n304 163.367
R1150 B.n305 B.n133 163.367
R1151 B.n309 B.n133 163.367
R1152 B.n310 B.n309 163.367
R1153 B.n310 B.n129 163.367
R1154 B.n314 B.n129 163.367
R1155 B.n315 B.n314 163.367
R1156 B.n316 B.n315 163.367
R1157 B.n316 B.n127 163.367
R1158 B.n320 B.n127 163.367
R1159 B.n321 B.n320 163.367
R1160 B.n322 B.n321 163.367
R1161 B.n322 B.n125 163.367
R1162 B.n326 B.n125 163.367
R1163 B.n327 B.n326 163.367
R1164 B.n328 B.n327 163.367
R1165 B.n328 B.n123 163.367
R1166 B.n332 B.n123 163.367
R1167 B.n333 B.n332 163.367
R1168 B.n334 B.n333 163.367
R1169 B.n334 B.n121 163.367
R1170 B.n338 B.n121 163.367
R1171 B.n339 B.n338 163.367
R1172 B.n340 B.n339 163.367
R1173 B.n340 B.n119 163.367
R1174 B.n344 B.n119 163.367
R1175 B.n345 B.n344 163.367
R1176 B.n346 B.n345 163.367
R1177 B.n346 B.n117 163.367
R1178 B.n350 B.n117 163.367
R1179 B.n351 B.n350 163.367
R1180 B.n352 B.n351 163.367
R1181 B.n352 B.n115 163.367
R1182 B.n356 B.n115 163.367
R1183 B.n357 B.n356 163.367
R1184 B.n358 B.n357 163.367
R1185 B.n358 B.n113 163.367
R1186 B.n362 B.n113 163.367
R1187 B.n363 B.n362 163.367
R1188 B.n364 B.n111 163.367
R1189 B.n368 B.n111 163.367
R1190 B.n369 B.n368 163.367
R1191 B.n370 B.n369 163.367
R1192 B.n370 B.n109 163.367
R1193 B.n374 B.n109 163.367
R1194 B.n375 B.n374 163.367
R1195 B.n376 B.n375 163.367
R1196 B.n376 B.n107 163.367
R1197 B.n380 B.n107 163.367
R1198 B.n381 B.n380 163.367
R1199 B.n382 B.n381 163.367
R1200 B.n382 B.n105 163.367
R1201 B.n386 B.n105 163.367
R1202 B.n387 B.n386 163.367
R1203 B.n388 B.n387 163.367
R1204 B.n388 B.n103 163.367
R1205 B.n392 B.n103 163.367
R1206 B.n393 B.n392 163.367
R1207 B.n394 B.n393 163.367
R1208 B.n394 B.n101 163.367
R1209 B.n398 B.n101 163.367
R1210 B.n399 B.n398 163.367
R1211 B.n400 B.n399 163.367
R1212 B.n400 B.n99 163.367
R1213 B.n404 B.n99 163.367
R1214 B.n405 B.n404 163.367
R1215 B.n406 B.n405 163.367
R1216 B.n406 B.n97 163.367
R1217 B.n410 B.n97 163.367
R1218 B.n411 B.n410 163.367
R1219 B.n412 B.n411 163.367
R1220 B.n412 B.n95 163.367
R1221 B.n416 B.n95 163.367
R1222 B.n417 B.n416 163.367
R1223 B.n418 B.n417 163.367
R1224 B.n418 B.n93 163.367
R1225 B.n422 B.n93 163.367
R1226 B.n423 B.n422 163.367
R1227 B.n424 B.n423 163.367
R1228 B.n424 B.n91 163.367
R1229 B.n428 B.n91 163.367
R1230 B.n429 B.n428 163.367
R1231 B.n430 B.n429 163.367
R1232 B.n430 B.n89 163.367
R1233 B.n434 B.n89 163.367
R1234 B.n435 B.n434 163.367
R1235 B.n436 B.n435 163.367
R1236 B.n436 B.n87 163.367
R1237 B.n440 B.n87 163.367
R1238 B.n441 B.n440 163.367
R1239 B.n442 B.n441 163.367
R1240 B.n442 B.n85 163.367
R1241 B.n446 B.n85 163.367
R1242 B.n447 B.n446 163.367
R1243 B.n448 B.n447 163.367
R1244 B.n448 B.n83 163.367
R1245 B.n452 B.n83 163.367
R1246 B.n453 B.n452 163.367
R1247 B.n454 B.n453 163.367
R1248 B.n454 B.n81 163.367
R1249 B.n458 B.n81 163.367
R1250 B.n459 B.n458 163.367
R1251 B.n460 B.n459 163.367
R1252 B.n460 B.n79 163.367
R1253 B.n464 B.n79 163.367
R1254 B.n465 B.n464 163.367
R1255 B.n466 B.n465 163.367
R1256 B.n466 B.n77 163.367
R1257 B.n470 B.n77 163.367
R1258 B.n471 B.n470 163.367
R1259 B.n472 B.n471 163.367
R1260 B.n472 B.n75 163.367
R1261 B.n476 B.n75 163.367
R1262 B.n477 B.n476 163.367
R1263 B.n478 B.n477 163.367
R1264 B.n478 B.n73 163.367
R1265 B.n482 B.n73 163.367
R1266 B.n483 B.n482 163.367
R1267 B.n484 B.n483 163.367
R1268 B.n484 B.n71 163.367
R1269 B.n488 B.n71 163.367
R1270 B.n489 B.n488 163.367
R1271 B.n490 B.n489 163.367
R1272 B.n490 B.n69 163.367
R1273 B.n494 B.n69 163.367
R1274 B.n616 B.n615 163.367
R1275 B.n615 B.n614 163.367
R1276 B.n614 B.n25 163.367
R1277 B.n610 B.n25 163.367
R1278 B.n610 B.n609 163.367
R1279 B.n609 B.n608 163.367
R1280 B.n608 B.n27 163.367
R1281 B.n604 B.n27 163.367
R1282 B.n604 B.n603 163.367
R1283 B.n603 B.n602 163.367
R1284 B.n602 B.n29 163.367
R1285 B.n598 B.n29 163.367
R1286 B.n598 B.n597 163.367
R1287 B.n597 B.n596 163.367
R1288 B.n596 B.n31 163.367
R1289 B.n592 B.n31 163.367
R1290 B.n592 B.n591 163.367
R1291 B.n591 B.n590 163.367
R1292 B.n590 B.n33 163.367
R1293 B.n586 B.n33 163.367
R1294 B.n586 B.n585 163.367
R1295 B.n585 B.n584 163.367
R1296 B.n584 B.n35 163.367
R1297 B.n580 B.n35 163.367
R1298 B.n580 B.n579 163.367
R1299 B.n579 B.n578 163.367
R1300 B.n578 B.n37 163.367
R1301 B.n574 B.n37 163.367
R1302 B.n574 B.n573 163.367
R1303 B.n573 B.n572 163.367
R1304 B.n572 B.n39 163.367
R1305 B.n568 B.n39 163.367
R1306 B.n568 B.n567 163.367
R1307 B.n567 B.n566 163.367
R1308 B.n566 B.n41 163.367
R1309 B.n561 B.n41 163.367
R1310 B.n561 B.n560 163.367
R1311 B.n560 B.n559 163.367
R1312 B.n559 B.n45 163.367
R1313 B.n555 B.n45 163.367
R1314 B.n555 B.n554 163.367
R1315 B.n554 B.n553 163.367
R1316 B.n553 B.n47 163.367
R1317 B.n549 B.n47 163.367
R1318 B.n549 B.n548 163.367
R1319 B.n548 B.n51 163.367
R1320 B.n544 B.n51 163.367
R1321 B.n544 B.n543 163.367
R1322 B.n543 B.n542 163.367
R1323 B.n542 B.n53 163.367
R1324 B.n538 B.n53 163.367
R1325 B.n538 B.n537 163.367
R1326 B.n537 B.n536 163.367
R1327 B.n536 B.n55 163.367
R1328 B.n532 B.n55 163.367
R1329 B.n532 B.n531 163.367
R1330 B.n531 B.n530 163.367
R1331 B.n530 B.n57 163.367
R1332 B.n526 B.n57 163.367
R1333 B.n526 B.n525 163.367
R1334 B.n525 B.n524 163.367
R1335 B.n524 B.n59 163.367
R1336 B.n520 B.n59 163.367
R1337 B.n520 B.n519 163.367
R1338 B.n519 B.n518 163.367
R1339 B.n518 B.n61 163.367
R1340 B.n514 B.n61 163.367
R1341 B.n514 B.n513 163.367
R1342 B.n513 B.n512 163.367
R1343 B.n512 B.n63 163.367
R1344 B.n508 B.n63 163.367
R1345 B.n508 B.n507 163.367
R1346 B.n507 B.n506 163.367
R1347 B.n506 B.n65 163.367
R1348 B.n502 B.n65 163.367
R1349 B.n502 B.n501 163.367
R1350 B.n501 B.n500 163.367
R1351 B.n500 B.n67 163.367
R1352 B.n496 B.n67 163.367
R1353 B.n496 B.n495 163.367
R1354 B.n131 B.n130 76.2187
R1355 B.n139 B.n138 76.2187
R1356 B.n43 B.n42 76.2187
R1357 B.n49 B.n48 76.2187
R1358 B.n132 B.n131 59.5399
R1359 B.n295 B.n139 59.5399
R1360 B.n563 B.n43 59.5399
R1361 B.n50 B.n49 59.5399
R1362 B.n618 B.n617 28.2542
R1363 B.n365 B.n112 28.2542
R1364 B.n241 B.n240 28.2542
R1365 B.n493 B.n68 28.2542
R1366 B B.n683 18.0485
R1367 B.n617 B.n24 10.6151
R1368 B.n613 B.n24 10.6151
R1369 B.n613 B.n612 10.6151
R1370 B.n612 B.n611 10.6151
R1371 B.n611 B.n26 10.6151
R1372 B.n607 B.n26 10.6151
R1373 B.n607 B.n606 10.6151
R1374 B.n606 B.n605 10.6151
R1375 B.n605 B.n28 10.6151
R1376 B.n601 B.n28 10.6151
R1377 B.n601 B.n600 10.6151
R1378 B.n600 B.n599 10.6151
R1379 B.n599 B.n30 10.6151
R1380 B.n595 B.n30 10.6151
R1381 B.n595 B.n594 10.6151
R1382 B.n594 B.n593 10.6151
R1383 B.n593 B.n32 10.6151
R1384 B.n589 B.n32 10.6151
R1385 B.n589 B.n588 10.6151
R1386 B.n588 B.n587 10.6151
R1387 B.n587 B.n34 10.6151
R1388 B.n583 B.n34 10.6151
R1389 B.n583 B.n582 10.6151
R1390 B.n582 B.n581 10.6151
R1391 B.n581 B.n36 10.6151
R1392 B.n577 B.n36 10.6151
R1393 B.n577 B.n576 10.6151
R1394 B.n576 B.n575 10.6151
R1395 B.n575 B.n38 10.6151
R1396 B.n571 B.n38 10.6151
R1397 B.n571 B.n570 10.6151
R1398 B.n570 B.n569 10.6151
R1399 B.n569 B.n40 10.6151
R1400 B.n565 B.n40 10.6151
R1401 B.n565 B.n564 10.6151
R1402 B.n562 B.n44 10.6151
R1403 B.n558 B.n44 10.6151
R1404 B.n558 B.n557 10.6151
R1405 B.n557 B.n556 10.6151
R1406 B.n556 B.n46 10.6151
R1407 B.n552 B.n46 10.6151
R1408 B.n552 B.n551 10.6151
R1409 B.n551 B.n550 10.6151
R1410 B.n547 B.n546 10.6151
R1411 B.n546 B.n545 10.6151
R1412 B.n545 B.n52 10.6151
R1413 B.n541 B.n52 10.6151
R1414 B.n541 B.n540 10.6151
R1415 B.n540 B.n539 10.6151
R1416 B.n539 B.n54 10.6151
R1417 B.n535 B.n54 10.6151
R1418 B.n535 B.n534 10.6151
R1419 B.n534 B.n533 10.6151
R1420 B.n533 B.n56 10.6151
R1421 B.n529 B.n56 10.6151
R1422 B.n529 B.n528 10.6151
R1423 B.n528 B.n527 10.6151
R1424 B.n527 B.n58 10.6151
R1425 B.n523 B.n58 10.6151
R1426 B.n523 B.n522 10.6151
R1427 B.n522 B.n521 10.6151
R1428 B.n521 B.n60 10.6151
R1429 B.n517 B.n60 10.6151
R1430 B.n517 B.n516 10.6151
R1431 B.n516 B.n515 10.6151
R1432 B.n515 B.n62 10.6151
R1433 B.n511 B.n62 10.6151
R1434 B.n511 B.n510 10.6151
R1435 B.n510 B.n509 10.6151
R1436 B.n509 B.n64 10.6151
R1437 B.n505 B.n64 10.6151
R1438 B.n505 B.n504 10.6151
R1439 B.n504 B.n503 10.6151
R1440 B.n503 B.n66 10.6151
R1441 B.n499 B.n66 10.6151
R1442 B.n499 B.n498 10.6151
R1443 B.n498 B.n497 10.6151
R1444 B.n497 B.n68 10.6151
R1445 B.n366 B.n365 10.6151
R1446 B.n367 B.n366 10.6151
R1447 B.n367 B.n110 10.6151
R1448 B.n371 B.n110 10.6151
R1449 B.n372 B.n371 10.6151
R1450 B.n373 B.n372 10.6151
R1451 B.n373 B.n108 10.6151
R1452 B.n377 B.n108 10.6151
R1453 B.n378 B.n377 10.6151
R1454 B.n379 B.n378 10.6151
R1455 B.n379 B.n106 10.6151
R1456 B.n383 B.n106 10.6151
R1457 B.n384 B.n383 10.6151
R1458 B.n385 B.n384 10.6151
R1459 B.n385 B.n104 10.6151
R1460 B.n389 B.n104 10.6151
R1461 B.n390 B.n389 10.6151
R1462 B.n391 B.n390 10.6151
R1463 B.n391 B.n102 10.6151
R1464 B.n395 B.n102 10.6151
R1465 B.n396 B.n395 10.6151
R1466 B.n397 B.n396 10.6151
R1467 B.n397 B.n100 10.6151
R1468 B.n401 B.n100 10.6151
R1469 B.n402 B.n401 10.6151
R1470 B.n403 B.n402 10.6151
R1471 B.n403 B.n98 10.6151
R1472 B.n407 B.n98 10.6151
R1473 B.n408 B.n407 10.6151
R1474 B.n409 B.n408 10.6151
R1475 B.n409 B.n96 10.6151
R1476 B.n413 B.n96 10.6151
R1477 B.n414 B.n413 10.6151
R1478 B.n415 B.n414 10.6151
R1479 B.n415 B.n94 10.6151
R1480 B.n419 B.n94 10.6151
R1481 B.n420 B.n419 10.6151
R1482 B.n421 B.n420 10.6151
R1483 B.n421 B.n92 10.6151
R1484 B.n425 B.n92 10.6151
R1485 B.n426 B.n425 10.6151
R1486 B.n427 B.n426 10.6151
R1487 B.n427 B.n90 10.6151
R1488 B.n431 B.n90 10.6151
R1489 B.n432 B.n431 10.6151
R1490 B.n433 B.n432 10.6151
R1491 B.n433 B.n88 10.6151
R1492 B.n437 B.n88 10.6151
R1493 B.n438 B.n437 10.6151
R1494 B.n439 B.n438 10.6151
R1495 B.n439 B.n86 10.6151
R1496 B.n443 B.n86 10.6151
R1497 B.n444 B.n443 10.6151
R1498 B.n445 B.n444 10.6151
R1499 B.n445 B.n84 10.6151
R1500 B.n449 B.n84 10.6151
R1501 B.n450 B.n449 10.6151
R1502 B.n451 B.n450 10.6151
R1503 B.n451 B.n82 10.6151
R1504 B.n455 B.n82 10.6151
R1505 B.n456 B.n455 10.6151
R1506 B.n457 B.n456 10.6151
R1507 B.n457 B.n80 10.6151
R1508 B.n461 B.n80 10.6151
R1509 B.n462 B.n461 10.6151
R1510 B.n463 B.n462 10.6151
R1511 B.n463 B.n78 10.6151
R1512 B.n467 B.n78 10.6151
R1513 B.n468 B.n467 10.6151
R1514 B.n469 B.n468 10.6151
R1515 B.n469 B.n76 10.6151
R1516 B.n473 B.n76 10.6151
R1517 B.n474 B.n473 10.6151
R1518 B.n475 B.n474 10.6151
R1519 B.n475 B.n74 10.6151
R1520 B.n479 B.n74 10.6151
R1521 B.n480 B.n479 10.6151
R1522 B.n481 B.n480 10.6151
R1523 B.n481 B.n72 10.6151
R1524 B.n485 B.n72 10.6151
R1525 B.n486 B.n485 10.6151
R1526 B.n487 B.n486 10.6151
R1527 B.n487 B.n70 10.6151
R1528 B.n491 B.n70 10.6151
R1529 B.n492 B.n491 10.6151
R1530 B.n493 B.n492 10.6151
R1531 B.n241 B.n156 10.6151
R1532 B.n245 B.n156 10.6151
R1533 B.n246 B.n245 10.6151
R1534 B.n247 B.n246 10.6151
R1535 B.n247 B.n154 10.6151
R1536 B.n251 B.n154 10.6151
R1537 B.n252 B.n251 10.6151
R1538 B.n253 B.n252 10.6151
R1539 B.n253 B.n152 10.6151
R1540 B.n257 B.n152 10.6151
R1541 B.n258 B.n257 10.6151
R1542 B.n259 B.n258 10.6151
R1543 B.n259 B.n150 10.6151
R1544 B.n263 B.n150 10.6151
R1545 B.n264 B.n263 10.6151
R1546 B.n265 B.n264 10.6151
R1547 B.n265 B.n148 10.6151
R1548 B.n269 B.n148 10.6151
R1549 B.n270 B.n269 10.6151
R1550 B.n271 B.n270 10.6151
R1551 B.n271 B.n146 10.6151
R1552 B.n275 B.n146 10.6151
R1553 B.n276 B.n275 10.6151
R1554 B.n277 B.n276 10.6151
R1555 B.n277 B.n144 10.6151
R1556 B.n281 B.n144 10.6151
R1557 B.n282 B.n281 10.6151
R1558 B.n283 B.n282 10.6151
R1559 B.n283 B.n142 10.6151
R1560 B.n287 B.n142 10.6151
R1561 B.n288 B.n287 10.6151
R1562 B.n289 B.n288 10.6151
R1563 B.n289 B.n140 10.6151
R1564 B.n293 B.n140 10.6151
R1565 B.n294 B.n293 10.6151
R1566 B.n296 B.n136 10.6151
R1567 B.n300 B.n136 10.6151
R1568 B.n301 B.n300 10.6151
R1569 B.n302 B.n301 10.6151
R1570 B.n302 B.n134 10.6151
R1571 B.n306 B.n134 10.6151
R1572 B.n307 B.n306 10.6151
R1573 B.n308 B.n307 10.6151
R1574 B.n312 B.n311 10.6151
R1575 B.n313 B.n312 10.6151
R1576 B.n313 B.n128 10.6151
R1577 B.n317 B.n128 10.6151
R1578 B.n318 B.n317 10.6151
R1579 B.n319 B.n318 10.6151
R1580 B.n319 B.n126 10.6151
R1581 B.n323 B.n126 10.6151
R1582 B.n324 B.n323 10.6151
R1583 B.n325 B.n324 10.6151
R1584 B.n325 B.n124 10.6151
R1585 B.n329 B.n124 10.6151
R1586 B.n330 B.n329 10.6151
R1587 B.n331 B.n330 10.6151
R1588 B.n331 B.n122 10.6151
R1589 B.n335 B.n122 10.6151
R1590 B.n336 B.n335 10.6151
R1591 B.n337 B.n336 10.6151
R1592 B.n337 B.n120 10.6151
R1593 B.n341 B.n120 10.6151
R1594 B.n342 B.n341 10.6151
R1595 B.n343 B.n342 10.6151
R1596 B.n343 B.n118 10.6151
R1597 B.n347 B.n118 10.6151
R1598 B.n348 B.n347 10.6151
R1599 B.n349 B.n348 10.6151
R1600 B.n349 B.n116 10.6151
R1601 B.n353 B.n116 10.6151
R1602 B.n354 B.n353 10.6151
R1603 B.n355 B.n354 10.6151
R1604 B.n355 B.n114 10.6151
R1605 B.n359 B.n114 10.6151
R1606 B.n360 B.n359 10.6151
R1607 B.n361 B.n360 10.6151
R1608 B.n361 B.n112 10.6151
R1609 B.n240 B.n239 10.6151
R1610 B.n239 B.n158 10.6151
R1611 B.n235 B.n158 10.6151
R1612 B.n235 B.n234 10.6151
R1613 B.n234 B.n233 10.6151
R1614 B.n233 B.n160 10.6151
R1615 B.n229 B.n160 10.6151
R1616 B.n229 B.n228 10.6151
R1617 B.n228 B.n227 10.6151
R1618 B.n227 B.n162 10.6151
R1619 B.n223 B.n162 10.6151
R1620 B.n223 B.n222 10.6151
R1621 B.n222 B.n221 10.6151
R1622 B.n221 B.n164 10.6151
R1623 B.n217 B.n164 10.6151
R1624 B.n217 B.n216 10.6151
R1625 B.n216 B.n215 10.6151
R1626 B.n215 B.n166 10.6151
R1627 B.n211 B.n166 10.6151
R1628 B.n211 B.n210 10.6151
R1629 B.n210 B.n209 10.6151
R1630 B.n209 B.n168 10.6151
R1631 B.n205 B.n168 10.6151
R1632 B.n205 B.n204 10.6151
R1633 B.n204 B.n203 10.6151
R1634 B.n203 B.n170 10.6151
R1635 B.n199 B.n170 10.6151
R1636 B.n199 B.n198 10.6151
R1637 B.n198 B.n197 10.6151
R1638 B.n197 B.n172 10.6151
R1639 B.n193 B.n172 10.6151
R1640 B.n193 B.n192 10.6151
R1641 B.n192 B.n191 10.6151
R1642 B.n191 B.n174 10.6151
R1643 B.n187 B.n174 10.6151
R1644 B.n187 B.n186 10.6151
R1645 B.n186 B.n185 10.6151
R1646 B.n185 B.n176 10.6151
R1647 B.n181 B.n176 10.6151
R1648 B.n181 B.n180 10.6151
R1649 B.n180 B.n179 10.6151
R1650 B.n179 B.n0 10.6151
R1651 B.n679 B.n1 10.6151
R1652 B.n679 B.n678 10.6151
R1653 B.n678 B.n677 10.6151
R1654 B.n677 B.n4 10.6151
R1655 B.n673 B.n4 10.6151
R1656 B.n673 B.n672 10.6151
R1657 B.n672 B.n671 10.6151
R1658 B.n671 B.n6 10.6151
R1659 B.n667 B.n6 10.6151
R1660 B.n667 B.n666 10.6151
R1661 B.n666 B.n665 10.6151
R1662 B.n665 B.n8 10.6151
R1663 B.n661 B.n8 10.6151
R1664 B.n661 B.n660 10.6151
R1665 B.n660 B.n659 10.6151
R1666 B.n659 B.n10 10.6151
R1667 B.n655 B.n10 10.6151
R1668 B.n655 B.n654 10.6151
R1669 B.n654 B.n653 10.6151
R1670 B.n653 B.n12 10.6151
R1671 B.n649 B.n12 10.6151
R1672 B.n649 B.n648 10.6151
R1673 B.n648 B.n647 10.6151
R1674 B.n647 B.n14 10.6151
R1675 B.n643 B.n14 10.6151
R1676 B.n643 B.n642 10.6151
R1677 B.n642 B.n641 10.6151
R1678 B.n641 B.n16 10.6151
R1679 B.n637 B.n16 10.6151
R1680 B.n637 B.n636 10.6151
R1681 B.n636 B.n635 10.6151
R1682 B.n635 B.n18 10.6151
R1683 B.n631 B.n18 10.6151
R1684 B.n631 B.n630 10.6151
R1685 B.n630 B.n629 10.6151
R1686 B.n629 B.n20 10.6151
R1687 B.n625 B.n20 10.6151
R1688 B.n625 B.n624 10.6151
R1689 B.n624 B.n623 10.6151
R1690 B.n623 B.n22 10.6151
R1691 B.n619 B.n22 10.6151
R1692 B.n619 B.n618 10.6151
R1693 B.n563 B.n562 6.5566
R1694 B.n550 B.n50 6.5566
R1695 B.n296 B.n295 6.5566
R1696 B.n308 B.n132 6.5566
R1697 B.n564 B.n563 4.05904
R1698 B.n547 B.n50 4.05904
R1699 B.n295 B.n294 4.05904
R1700 B.n311 B.n132 4.05904
R1701 B.n683 B.n0 2.81026
R1702 B.n683 B.n1 2.81026
R1703 VP.n19 VP.n18 161.3
R1704 VP.n17 VP.n1 161.3
R1705 VP.n16 VP.n15 161.3
R1706 VP.n14 VP.n2 161.3
R1707 VP.n13 VP.n12 161.3
R1708 VP.n11 VP.n3 161.3
R1709 VP.n10 VP.n9 161.3
R1710 VP.n8 VP.n4 161.3
R1711 VP.n5 VP.t0 101.349
R1712 VP.n5 VP.t1 100.105
R1713 VP.n7 VP.n6 79.5466
R1714 VP.n20 VP.n0 79.5466
R1715 VP.n6 VP.t2 66.4763
R1716 VP.n0 VP.t3 66.4763
R1717 VP.n12 VP.n2 56.5193
R1718 VP.n7 VP.n5 50.0056
R1719 VP.n10 VP.n4 24.4675
R1720 VP.n11 VP.n10 24.4675
R1721 VP.n12 VP.n11 24.4675
R1722 VP.n16 VP.n2 24.4675
R1723 VP.n17 VP.n16 24.4675
R1724 VP.n18 VP.n17 24.4675
R1725 VP.n6 VP.n4 10.5213
R1726 VP.n18 VP.n0 10.5213
R1727 VP.n8 VP.n7 0.354971
R1728 VP.n20 VP.n19 0.354971
R1729 VP VP.n20 0.26696
R1730 VP.n9 VP.n8 0.189894
R1731 VP.n9 VP.n3 0.189894
R1732 VP.n13 VP.n3 0.189894
R1733 VP.n14 VP.n13 0.189894
R1734 VP.n15 VP.n14 0.189894
R1735 VP.n15 VP.n1 0.189894
R1736 VP.n19 VP.n1 0.189894
R1737 VDD1 VDD1.n1 119.501
R1738 VDD1 VDD1.n0 76.5952
R1739 VDD1.n0 VDD1.t3 3.27391
R1740 VDD1.n0 VDD1.t2 3.27391
R1741 VDD1.n1 VDD1.t1 3.27391
R1742 VDD1.n1 VDD1.t0 3.27391
C0 B VTAIL 4.64189f
C1 B w_n3328_n2954# 9.89496f
C2 B VDD1 1.38308f
C3 B VDD2 1.45178f
C4 VN B 1.27414f
C5 VTAIL VP 4.36177f
C6 w_n3328_n2954# VP 6.20668f
C7 VDD1 VP 4.49488f
C8 w_n3328_n2954# VTAIL 3.55641f
C9 VDD1 VTAIL 5.23703f
C10 VDD2 VP 0.458089f
C11 VN VP 6.52705f
C12 w_n3328_n2954# VDD1 1.58739f
C13 VDD2 VTAIL 5.29794f
C14 VN VTAIL 4.34766f
C15 w_n3328_n2954# VDD2 1.66556f
C16 VN w_n3328_n2954# 5.77632f
C17 VDD2 VDD1 1.26764f
C18 VN VDD1 0.150056f
C19 VN VDD2 4.18784f
C20 B VP 1.99295f
C21 VDD2 VSUBS 1.064234f
C22 VDD1 VSUBS 6.05901f
C23 VTAIL VSUBS 1.253445f
C24 VN VSUBS 5.98822f
C25 VP VSUBS 2.741485f
C26 B VSUBS 4.961504f
C27 w_n3328_n2954# VSUBS 0.121445p
C28 VDD1.t3 VSUBS 0.218154f
C29 VDD1.t2 VSUBS 0.218154f
C30 VDD1.n0 VSUBS 1.64342f
C31 VDD1.t1 VSUBS 0.218154f
C32 VDD1.t0 VSUBS 0.218154f
C33 VDD1.n1 VSUBS 2.3576f
C34 VP.t3 VSUBS 2.97025f
C35 VP.n0 VSUBS 1.17517f
C36 VP.n1 VSUBS 0.030678f
C37 VP.n2 VSUBS 0.044785f
C38 VP.n3 VSUBS 0.030678f
C39 VP.n4 VSUBS 0.041085f
C40 VP.t0 VSUBS 3.41668f
C41 VP.t1 VSUBS 3.40154f
C42 VP.n5 VSUBS 3.89651f
C43 VP.t2 VSUBS 2.97025f
C44 VP.n6 VSUBS 1.17517f
C45 VP.n7 VSUBS 1.76083f
C46 VP.n8 VSUBS 0.049514f
C47 VP.n9 VSUBS 0.030678f
C48 VP.n10 VSUBS 0.057176f
C49 VP.n11 VSUBS 0.057176f
C50 VP.n12 VSUBS 0.044785f
C51 VP.n13 VSUBS 0.030678f
C52 VP.n14 VSUBS 0.030678f
C53 VP.n15 VSUBS 0.030678f
C54 VP.n16 VSUBS 0.057176f
C55 VP.n17 VSUBS 0.057176f
C56 VP.n18 VSUBS 0.041085f
C57 VP.n19 VSUBS 0.049514f
C58 VP.n20 VSUBS 0.083253f
C59 B.n0 VSUBS 0.004188f
C60 B.n1 VSUBS 0.004188f
C61 B.n2 VSUBS 0.006624f
C62 B.n3 VSUBS 0.006624f
C63 B.n4 VSUBS 0.006624f
C64 B.n5 VSUBS 0.006624f
C65 B.n6 VSUBS 0.006624f
C66 B.n7 VSUBS 0.006624f
C67 B.n8 VSUBS 0.006624f
C68 B.n9 VSUBS 0.006624f
C69 B.n10 VSUBS 0.006624f
C70 B.n11 VSUBS 0.006624f
C71 B.n12 VSUBS 0.006624f
C72 B.n13 VSUBS 0.006624f
C73 B.n14 VSUBS 0.006624f
C74 B.n15 VSUBS 0.006624f
C75 B.n16 VSUBS 0.006624f
C76 B.n17 VSUBS 0.006624f
C77 B.n18 VSUBS 0.006624f
C78 B.n19 VSUBS 0.006624f
C79 B.n20 VSUBS 0.006624f
C80 B.n21 VSUBS 0.006624f
C81 B.n22 VSUBS 0.006624f
C82 B.n23 VSUBS 0.013716f
C83 B.n24 VSUBS 0.006624f
C84 B.n25 VSUBS 0.006624f
C85 B.n26 VSUBS 0.006624f
C86 B.n27 VSUBS 0.006624f
C87 B.n28 VSUBS 0.006624f
C88 B.n29 VSUBS 0.006624f
C89 B.n30 VSUBS 0.006624f
C90 B.n31 VSUBS 0.006624f
C91 B.n32 VSUBS 0.006624f
C92 B.n33 VSUBS 0.006624f
C93 B.n34 VSUBS 0.006624f
C94 B.n35 VSUBS 0.006624f
C95 B.n36 VSUBS 0.006624f
C96 B.n37 VSUBS 0.006624f
C97 B.n38 VSUBS 0.006624f
C98 B.n39 VSUBS 0.006624f
C99 B.n40 VSUBS 0.006624f
C100 B.n41 VSUBS 0.006624f
C101 B.t11 VSUBS 0.156972f
C102 B.t10 VSUBS 0.194609f
C103 B.t9 VSUBS 1.58806f
C104 B.n42 VSUBS 0.313496f
C105 B.n43 VSUBS 0.2141f
C106 B.n44 VSUBS 0.006624f
C107 B.n45 VSUBS 0.006624f
C108 B.n46 VSUBS 0.006624f
C109 B.n47 VSUBS 0.006624f
C110 B.t2 VSUBS 0.156974f
C111 B.t1 VSUBS 0.194611f
C112 B.t0 VSUBS 1.58806f
C113 B.n48 VSUBS 0.313493f
C114 B.n49 VSUBS 0.214097f
C115 B.n50 VSUBS 0.015346f
C116 B.n51 VSUBS 0.006624f
C117 B.n52 VSUBS 0.006624f
C118 B.n53 VSUBS 0.006624f
C119 B.n54 VSUBS 0.006624f
C120 B.n55 VSUBS 0.006624f
C121 B.n56 VSUBS 0.006624f
C122 B.n57 VSUBS 0.006624f
C123 B.n58 VSUBS 0.006624f
C124 B.n59 VSUBS 0.006624f
C125 B.n60 VSUBS 0.006624f
C126 B.n61 VSUBS 0.006624f
C127 B.n62 VSUBS 0.006624f
C128 B.n63 VSUBS 0.006624f
C129 B.n64 VSUBS 0.006624f
C130 B.n65 VSUBS 0.006624f
C131 B.n66 VSUBS 0.006624f
C132 B.n67 VSUBS 0.006624f
C133 B.n68 VSUBS 0.013627f
C134 B.n69 VSUBS 0.006624f
C135 B.n70 VSUBS 0.006624f
C136 B.n71 VSUBS 0.006624f
C137 B.n72 VSUBS 0.006624f
C138 B.n73 VSUBS 0.006624f
C139 B.n74 VSUBS 0.006624f
C140 B.n75 VSUBS 0.006624f
C141 B.n76 VSUBS 0.006624f
C142 B.n77 VSUBS 0.006624f
C143 B.n78 VSUBS 0.006624f
C144 B.n79 VSUBS 0.006624f
C145 B.n80 VSUBS 0.006624f
C146 B.n81 VSUBS 0.006624f
C147 B.n82 VSUBS 0.006624f
C148 B.n83 VSUBS 0.006624f
C149 B.n84 VSUBS 0.006624f
C150 B.n85 VSUBS 0.006624f
C151 B.n86 VSUBS 0.006624f
C152 B.n87 VSUBS 0.006624f
C153 B.n88 VSUBS 0.006624f
C154 B.n89 VSUBS 0.006624f
C155 B.n90 VSUBS 0.006624f
C156 B.n91 VSUBS 0.006624f
C157 B.n92 VSUBS 0.006624f
C158 B.n93 VSUBS 0.006624f
C159 B.n94 VSUBS 0.006624f
C160 B.n95 VSUBS 0.006624f
C161 B.n96 VSUBS 0.006624f
C162 B.n97 VSUBS 0.006624f
C163 B.n98 VSUBS 0.006624f
C164 B.n99 VSUBS 0.006624f
C165 B.n100 VSUBS 0.006624f
C166 B.n101 VSUBS 0.006624f
C167 B.n102 VSUBS 0.006624f
C168 B.n103 VSUBS 0.006624f
C169 B.n104 VSUBS 0.006624f
C170 B.n105 VSUBS 0.006624f
C171 B.n106 VSUBS 0.006624f
C172 B.n107 VSUBS 0.006624f
C173 B.n108 VSUBS 0.006624f
C174 B.n109 VSUBS 0.006624f
C175 B.n110 VSUBS 0.006624f
C176 B.n111 VSUBS 0.006624f
C177 B.n112 VSUBS 0.014532f
C178 B.n113 VSUBS 0.006624f
C179 B.n114 VSUBS 0.006624f
C180 B.n115 VSUBS 0.006624f
C181 B.n116 VSUBS 0.006624f
C182 B.n117 VSUBS 0.006624f
C183 B.n118 VSUBS 0.006624f
C184 B.n119 VSUBS 0.006624f
C185 B.n120 VSUBS 0.006624f
C186 B.n121 VSUBS 0.006624f
C187 B.n122 VSUBS 0.006624f
C188 B.n123 VSUBS 0.006624f
C189 B.n124 VSUBS 0.006624f
C190 B.n125 VSUBS 0.006624f
C191 B.n126 VSUBS 0.006624f
C192 B.n127 VSUBS 0.006624f
C193 B.n128 VSUBS 0.006624f
C194 B.n129 VSUBS 0.006624f
C195 B.t7 VSUBS 0.156974f
C196 B.t8 VSUBS 0.194611f
C197 B.t6 VSUBS 1.58806f
C198 B.n130 VSUBS 0.313493f
C199 B.n131 VSUBS 0.214097f
C200 B.n132 VSUBS 0.015346f
C201 B.n133 VSUBS 0.006624f
C202 B.n134 VSUBS 0.006624f
C203 B.n135 VSUBS 0.006624f
C204 B.n136 VSUBS 0.006624f
C205 B.n137 VSUBS 0.006624f
C206 B.t4 VSUBS 0.156972f
C207 B.t5 VSUBS 0.194609f
C208 B.t3 VSUBS 1.58806f
C209 B.n138 VSUBS 0.313496f
C210 B.n139 VSUBS 0.2141f
C211 B.n140 VSUBS 0.006624f
C212 B.n141 VSUBS 0.006624f
C213 B.n142 VSUBS 0.006624f
C214 B.n143 VSUBS 0.006624f
C215 B.n144 VSUBS 0.006624f
C216 B.n145 VSUBS 0.006624f
C217 B.n146 VSUBS 0.006624f
C218 B.n147 VSUBS 0.006624f
C219 B.n148 VSUBS 0.006624f
C220 B.n149 VSUBS 0.006624f
C221 B.n150 VSUBS 0.006624f
C222 B.n151 VSUBS 0.006624f
C223 B.n152 VSUBS 0.006624f
C224 B.n153 VSUBS 0.006624f
C225 B.n154 VSUBS 0.006624f
C226 B.n155 VSUBS 0.006624f
C227 B.n156 VSUBS 0.006624f
C228 B.n157 VSUBS 0.013716f
C229 B.n158 VSUBS 0.006624f
C230 B.n159 VSUBS 0.006624f
C231 B.n160 VSUBS 0.006624f
C232 B.n161 VSUBS 0.006624f
C233 B.n162 VSUBS 0.006624f
C234 B.n163 VSUBS 0.006624f
C235 B.n164 VSUBS 0.006624f
C236 B.n165 VSUBS 0.006624f
C237 B.n166 VSUBS 0.006624f
C238 B.n167 VSUBS 0.006624f
C239 B.n168 VSUBS 0.006624f
C240 B.n169 VSUBS 0.006624f
C241 B.n170 VSUBS 0.006624f
C242 B.n171 VSUBS 0.006624f
C243 B.n172 VSUBS 0.006624f
C244 B.n173 VSUBS 0.006624f
C245 B.n174 VSUBS 0.006624f
C246 B.n175 VSUBS 0.006624f
C247 B.n176 VSUBS 0.006624f
C248 B.n177 VSUBS 0.006624f
C249 B.n178 VSUBS 0.006624f
C250 B.n179 VSUBS 0.006624f
C251 B.n180 VSUBS 0.006624f
C252 B.n181 VSUBS 0.006624f
C253 B.n182 VSUBS 0.006624f
C254 B.n183 VSUBS 0.006624f
C255 B.n184 VSUBS 0.006624f
C256 B.n185 VSUBS 0.006624f
C257 B.n186 VSUBS 0.006624f
C258 B.n187 VSUBS 0.006624f
C259 B.n188 VSUBS 0.006624f
C260 B.n189 VSUBS 0.006624f
C261 B.n190 VSUBS 0.006624f
C262 B.n191 VSUBS 0.006624f
C263 B.n192 VSUBS 0.006624f
C264 B.n193 VSUBS 0.006624f
C265 B.n194 VSUBS 0.006624f
C266 B.n195 VSUBS 0.006624f
C267 B.n196 VSUBS 0.006624f
C268 B.n197 VSUBS 0.006624f
C269 B.n198 VSUBS 0.006624f
C270 B.n199 VSUBS 0.006624f
C271 B.n200 VSUBS 0.006624f
C272 B.n201 VSUBS 0.006624f
C273 B.n202 VSUBS 0.006624f
C274 B.n203 VSUBS 0.006624f
C275 B.n204 VSUBS 0.006624f
C276 B.n205 VSUBS 0.006624f
C277 B.n206 VSUBS 0.006624f
C278 B.n207 VSUBS 0.006624f
C279 B.n208 VSUBS 0.006624f
C280 B.n209 VSUBS 0.006624f
C281 B.n210 VSUBS 0.006624f
C282 B.n211 VSUBS 0.006624f
C283 B.n212 VSUBS 0.006624f
C284 B.n213 VSUBS 0.006624f
C285 B.n214 VSUBS 0.006624f
C286 B.n215 VSUBS 0.006624f
C287 B.n216 VSUBS 0.006624f
C288 B.n217 VSUBS 0.006624f
C289 B.n218 VSUBS 0.006624f
C290 B.n219 VSUBS 0.006624f
C291 B.n220 VSUBS 0.006624f
C292 B.n221 VSUBS 0.006624f
C293 B.n222 VSUBS 0.006624f
C294 B.n223 VSUBS 0.006624f
C295 B.n224 VSUBS 0.006624f
C296 B.n225 VSUBS 0.006624f
C297 B.n226 VSUBS 0.006624f
C298 B.n227 VSUBS 0.006624f
C299 B.n228 VSUBS 0.006624f
C300 B.n229 VSUBS 0.006624f
C301 B.n230 VSUBS 0.006624f
C302 B.n231 VSUBS 0.006624f
C303 B.n232 VSUBS 0.006624f
C304 B.n233 VSUBS 0.006624f
C305 B.n234 VSUBS 0.006624f
C306 B.n235 VSUBS 0.006624f
C307 B.n236 VSUBS 0.006624f
C308 B.n237 VSUBS 0.006624f
C309 B.n238 VSUBS 0.006624f
C310 B.n239 VSUBS 0.006624f
C311 B.n240 VSUBS 0.013716f
C312 B.n241 VSUBS 0.014532f
C313 B.n242 VSUBS 0.014532f
C314 B.n243 VSUBS 0.006624f
C315 B.n244 VSUBS 0.006624f
C316 B.n245 VSUBS 0.006624f
C317 B.n246 VSUBS 0.006624f
C318 B.n247 VSUBS 0.006624f
C319 B.n248 VSUBS 0.006624f
C320 B.n249 VSUBS 0.006624f
C321 B.n250 VSUBS 0.006624f
C322 B.n251 VSUBS 0.006624f
C323 B.n252 VSUBS 0.006624f
C324 B.n253 VSUBS 0.006624f
C325 B.n254 VSUBS 0.006624f
C326 B.n255 VSUBS 0.006624f
C327 B.n256 VSUBS 0.006624f
C328 B.n257 VSUBS 0.006624f
C329 B.n258 VSUBS 0.006624f
C330 B.n259 VSUBS 0.006624f
C331 B.n260 VSUBS 0.006624f
C332 B.n261 VSUBS 0.006624f
C333 B.n262 VSUBS 0.006624f
C334 B.n263 VSUBS 0.006624f
C335 B.n264 VSUBS 0.006624f
C336 B.n265 VSUBS 0.006624f
C337 B.n266 VSUBS 0.006624f
C338 B.n267 VSUBS 0.006624f
C339 B.n268 VSUBS 0.006624f
C340 B.n269 VSUBS 0.006624f
C341 B.n270 VSUBS 0.006624f
C342 B.n271 VSUBS 0.006624f
C343 B.n272 VSUBS 0.006624f
C344 B.n273 VSUBS 0.006624f
C345 B.n274 VSUBS 0.006624f
C346 B.n275 VSUBS 0.006624f
C347 B.n276 VSUBS 0.006624f
C348 B.n277 VSUBS 0.006624f
C349 B.n278 VSUBS 0.006624f
C350 B.n279 VSUBS 0.006624f
C351 B.n280 VSUBS 0.006624f
C352 B.n281 VSUBS 0.006624f
C353 B.n282 VSUBS 0.006624f
C354 B.n283 VSUBS 0.006624f
C355 B.n284 VSUBS 0.006624f
C356 B.n285 VSUBS 0.006624f
C357 B.n286 VSUBS 0.006624f
C358 B.n287 VSUBS 0.006624f
C359 B.n288 VSUBS 0.006624f
C360 B.n289 VSUBS 0.006624f
C361 B.n290 VSUBS 0.006624f
C362 B.n291 VSUBS 0.006624f
C363 B.n292 VSUBS 0.006624f
C364 B.n293 VSUBS 0.006624f
C365 B.n294 VSUBS 0.004578f
C366 B.n295 VSUBS 0.015346f
C367 B.n296 VSUBS 0.005357f
C368 B.n297 VSUBS 0.006624f
C369 B.n298 VSUBS 0.006624f
C370 B.n299 VSUBS 0.006624f
C371 B.n300 VSUBS 0.006624f
C372 B.n301 VSUBS 0.006624f
C373 B.n302 VSUBS 0.006624f
C374 B.n303 VSUBS 0.006624f
C375 B.n304 VSUBS 0.006624f
C376 B.n305 VSUBS 0.006624f
C377 B.n306 VSUBS 0.006624f
C378 B.n307 VSUBS 0.006624f
C379 B.n308 VSUBS 0.005357f
C380 B.n309 VSUBS 0.006624f
C381 B.n310 VSUBS 0.006624f
C382 B.n311 VSUBS 0.004578f
C383 B.n312 VSUBS 0.006624f
C384 B.n313 VSUBS 0.006624f
C385 B.n314 VSUBS 0.006624f
C386 B.n315 VSUBS 0.006624f
C387 B.n316 VSUBS 0.006624f
C388 B.n317 VSUBS 0.006624f
C389 B.n318 VSUBS 0.006624f
C390 B.n319 VSUBS 0.006624f
C391 B.n320 VSUBS 0.006624f
C392 B.n321 VSUBS 0.006624f
C393 B.n322 VSUBS 0.006624f
C394 B.n323 VSUBS 0.006624f
C395 B.n324 VSUBS 0.006624f
C396 B.n325 VSUBS 0.006624f
C397 B.n326 VSUBS 0.006624f
C398 B.n327 VSUBS 0.006624f
C399 B.n328 VSUBS 0.006624f
C400 B.n329 VSUBS 0.006624f
C401 B.n330 VSUBS 0.006624f
C402 B.n331 VSUBS 0.006624f
C403 B.n332 VSUBS 0.006624f
C404 B.n333 VSUBS 0.006624f
C405 B.n334 VSUBS 0.006624f
C406 B.n335 VSUBS 0.006624f
C407 B.n336 VSUBS 0.006624f
C408 B.n337 VSUBS 0.006624f
C409 B.n338 VSUBS 0.006624f
C410 B.n339 VSUBS 0.006624f
C411 B.n340 VSUBS 0.006624f
C412 B.n341 VSUBS 0.006624f
C413 B.n342 VSUBS 0.006624f
C414 B.n343 VSUBS 0.006624f
C415 B.n344 VSUBS 0.006624f
C416 B.n345 VSUBS 0.006624f
C417 B.n346 VSUBS 0.006624f
C418 B.n347 VSUBS 0.006624f
C419 B.n348 VSUBS 0.006624f
C420 B.n349 VSUBS 0.006624f
C421 B.n350 VSUBS 0.006624f
C422 B.n351 VSUBS 0.006624f
C423 B.n352 VSUBS 0.006624f
C424 B.n353 VSUBS 0.006624f
C425 B.n354 VSUBS 0.006624f
C426 B.n355 VSUBS 0.006624f
C427 B.n356 VSUBS 0.006624f
C428 B.n357 VSUBS 0.006624f
C429 B.n358 VSUBS 0.006624f
C430 B.n359 VSUBS 0.006624f
C431 B.n360 VSUBS 0.006624f
C432 B.n361 VSUBS 0.006624f
C433 B.n362 VSUBS 0.006624f
C434 B.n363 VSUBS 0.014532f
C435 B.n364 VSUBS 0.013716f
C436 B.n365 VSUBS 0.013716f
C437 B.n366 VSUBS 0.006624f
C438 B.n367 VSUBS 0.006624f
C439 B.n368 VSUBS 0.006624f
C440 B.n369 VSUBS 0.006624f
C441 B.n370 VSUBS 0.006624f
C442 B.n371 VSUBS 0.006624f
C443 B.n372 VSUBS 0.006624f
C444 B.n373 VSUBS 0.006624f
C445 B.n374 VSUBS 0.006624f
C446 B.n375 VSUBS 0.006624f
C447 B.n376 VSUBS 0.006624f
C448 B.n377 VSUBS 0.006624f
C449 B.n378 VSUBS 0.006624f
C450 B.n379 VSUBS 0.006624f
C451 B.n380 VSUBS 0.006624f
C452 B.n381 VSUBS 0.006624f
C453 B.n382 VSUBS 0.006624f
C454 B.n383 VSUBS 0.006624f
C455 B.n384 VSUBS 0.006624f
C456 B.n385 VSUBS 0.006624f
C457 B.n386 VSUBS 0.006624f
C458 B.n387 VSUBS 0.006624f
C459 B.n388 VSUBS 0.006624f
C460 B.n389 VSUBS 0.006624f
C461 B.n390 VSUBS 0.006624f
C462 B.n391 VSUBS 0.006624f
C463 B.n392 VSUBS 0.006624f
C464 B.n393 VSUBS 0.006624f
C465 B.n394 VSUBS 0.006624f
C466 B.n395 VSUBS 0.006624f
C467 B.n396 VSUBS 0.006624f
C468 B.n397 VSUBS 0.006624f
C469 B.n398 VSUBS 0.006624f
C470 B.n399 VSUBS 0.006624f
C471 B.n400 VSUBS 0.006624f
C472 B.n401 VSUBS 0.006624f
C473 B.n402 VSUBS 0.006624f
C474 B.n403 VSUBS 0.006624f
C475 B.n404 VSUBS 0.006624f
C476 B.n405 VSUBS 0.006624f
C477 B.n406 VSUBS 0.006624f
C478 B.n407 VSUBS 0.006624f
C479 B.n408 VSUBS 0.006624f
C480 B.n409 VSUBS 0.006624f
C481 B.n410 VSUBS 0.006624f
C482 B.n411 VSUBS 0.006624f
C483 B.n412 VSUBS 0.006624f
C484 B.n413 VSUBS 0.006624f
C485 B.n414 VSUBS 0.006624f
C486 B.n415 VSUBS 0.006624f
C487 B.n416 VSUBS 0.006624f
C488 B.n417 VSUBS 0.006624f
C489 B.n418 VSUBS 0.006624f
C490 B.n419 VSUBS 0.006624f
C491 B.n420 VSUBS 0.006624f
C492 B.n421 VSUBS 0.006624f
C493 B.n422 VSUBS 0.006624f
C494 B.n423 VSUBS 0.006624f
C495 B.n424 VSUBS 0.006624f
C496 B.n425 VSUBS 0.006624f
C497 B.n426 VSUBS 0.006624f
C498 B.n427 VSUBS 0.006624f
C499 B.n428 VSUBS 0.006624f
C500 B.n429 VSUBS 0.006624f
C501 B.n430 VSUBS 0.006624f
C502 B.n431 VSUBS 0.006624f
C503 B.n432 VSUBS 0.006624f
C504 B.n433 VSUBS 0.006624f
C505 B.n434 VSUBS 0.006624f
C506 B.n435 VSUBS 0.006624f
C507 B.n436 VSUBS 0.006624f
C508 B.n437 VSUBS 0.006624f
C509 B.n438 VSUBS 0.006624f
C510 B.n439 VSUBS 0.006624f
C511 B.n440 VSUBS 0.006624f
C512 B.n441 VSUBS 0.006624f
C513 B.n442 VSUBS 0.006624f
C514 B.n443 VSUBS 0.006624f
C515 B.n444 VSUBS 0.006624f
C516 B.n445 VSUBS 0.006624f
C517 B.n446 VSUBS 0.006624f
C518 B.n447 VSUBS 0.006624f
C519 B.n448 VSUBS 0.006624f
C520 B.n449 VSUBS 0.006624f
C521 B.n450 VSUBS 0.006624f
C522 B.n451 VSUBS 0.006624f
C523 B.n452 VSUBS 0.006624f
C524 B.n453 VSUBS 0.006624f
C525 B.n454 VSUBS 0.006624f
C526 B.n455 VSUBS 0.006624f
C527 B.n456 VSUBS 0.006624f
C528 B.n457 VSUBS 0.006624f
C529 B.n458 VSUBS 0.006624f
C530 B.n459 VSUBS 0.006624f
C531 B.n460 VSUBS 0.006624f
C532 B.n461 VSUBS 0.006624f
C533 B.n462 VSUBS 0.006624f
C534 B.n463 VSUBS 0.006624f
C535 B.n464 VSUBS 0.006624f
C536 B.n465 VSUBS 0.006624f
C537 B.n466 VSUBS 0.006624f
C538 B.n467 VSUBS 0.006624f
C539 B.n468 VSUBS 0.006624f
C540 B.n469 VSUBS 0.006624f
C541 B.n470 VSUBS 0.006624f
C542 B.n471 VSUBS 0.006624f
C543 B.n472 VSUBS 0.006624f
C544 B.n473 VSUBS 0.006624f
C545 B.n474 VSUBS 0.006624f
C546 B.n475 VSUBS 0.006624f
C547 B.n476 VSUBS 0.006624f
C548 B.n477 VSUBS 0.006624f
C549 B.n478 VSUBS 0.006624f
C550 B.n479 VSUBS 0.006624f
C551 B.n480 VSUBS 0.006624f
C552 B.n481 VSUBS 0.006624f
C553 B.n482 VSUBS 0.006624f
C554 B.n483 VSUBS 0.006624f
C555 B.n484 VSUBS 0.006624f
C556 B.n485 VSUBS 0.006624f
C557 B.n486 VSUBS 0.006624f
C558 B.n487 VSUBS 0.006624f
C559 B.n488 VSUBS 0.006624f
C560 B.n489 VSUBS 0.006624f
C561 B.n490 VSUBS 0.006624f
C562 B.n491 VSUBS 0.006624f
C563 B.n492 VSUBS 0.006624f
C564 B.n493 VSUBS 0.01462f
C565 B.n494 VSUBS 0.013716f
C566 B.n495 VSUBS 0.014532f
C567 B.n496 VSUBS 0.006624f
C568 B.n497 VSUBS 0.006624f
C569 B.n498 VSUBS 0.006624f
C570 B.n499 VSUBS 0.006624f
C571 B.n500 VSUBS 0.006624f
C572 B.n501 VSUBS 0.006624f
C573 B.n502 VSUBS 0.006624f
C574 B.n503 VSUBS 0.006624f
C575 B.n504 VSUBS 0.006624f
C576 B.n505 VSUBS 0.006624f
C577 B.n506 VSUBS 0.006624f
C578 B.n507 VSUBS 0.006624f
C579 B.n508 VSUBS 0.006624f
C580 B.n509 VSUBS 0.006624f
C581 B.n510 VSUBS 0.006624f
C582 B.n511 VSUBS 0.006624f
C583 B.n512 VSUBS 0.006624f
C584 B.n513 VSUBS 0.006624f
C585 B.n514 VSUBS 0.006624f
C586 B.n515 VSUBS 0.006624f
C587 B.n516 VSUBS 0.006624f
C588 B.n517 VSUBS 0.006624f
C589 B.n518 VSUBS 0.006624f
C590 B.n519 VSUBS 0.006624f
C591 B.n520 VSUBS 0.006624f
C592 B.n521 VSUBS 0.006624f
C593 B.n522 VSUBS 0.006624f
C594 B.n523 VSUBS 0.006624f
C595 B.n524 VSUBS 0.006624f
C596 B.n525 VSUBS 0.006624f
C597 B.n526 VSUBS 0.006624f
C598 B.n527 VSUBS 0.006624f
C599 B.n528 VSUBS 0.006624f
C600 B.n529 VSUBS 0.006624f
C601 B.n530 VSUBS 0.006624f
C602 B.n531 VSUBS 0.006624f
C603 B.n532 VSUBS 0.006624f
C604 B.n533 VSUBS 0.006624f
C605 B.n534 VSUBS 0.006624f
C606 B.n535 VSUBS 0.006624f
C607 B.n536 VSUBS 0.006624f
C608 B.n537 VSUBS 0.006624f
C609 B.n538 VSUBS 0.006624f
C610 B.n539 VSUBS 0.006624f
C611 B.n540 VSUBS 0.006624f
C612 B.n541 VSUBS 0.006624f
C613 B.n542 VSUBS 0.006624f
C614 B.n543 VSUBS 0.006624f
C615 B.n544 VSUBS 0.006624f
C616 B.n545 VSUBS 0.006624f
C617 B.n546 VSUBS 0.006624f
C618 B.n547 VSUBS 0.004578f
C619 B.n548 VSUBS 0.006624f
C620 B.n549 VSUBS 0.006624f
C621 B.n550 VSUBS 0.005357f
C622 B.n551 VSUBS 0.006624f
C623 B.n552 VSUBS 0.006624f
C624 B.n553 VSUBS 0.006624f
C625 B.n554 VSUBS 0.006624f
C626 B.n555 VSUBS 0.006624f
C627 B.n556 VSUBS 0.006624f
C628 B.n557 VSUBS 0.006624f
C629 B.n558 VSUBS 0.006624f
C630 B.n559 VSUBS 0.006624f
C631 B.n560 VSUBS 0.006624f
C632 B.n561 VSUBS 0.006624f
C633 B.n562 VSUBS 0.005357f
C634 B.n563 VSUBS 0.015346f
C635 B.n564 VSUBS 0.004578f
C636 B.n565 VSUBS 0.006624f
C637 B.n566 VSUBS 0.006624f
C638 B.n567 VSUBS 0.006624f
C639 B.n568 VSUBS 0.006624f
C640 B.n569 VSUBS 0.006624f
C641 B.n570 VSUBS 0.006624f
C642 B.n571 VSUBS 0.006624f
C643 B.n572 VSUBS 0.006624f
C644 B.n573 VSUBS 0.006624f
C645 B.n574 VSUBS 0.006624f
C646 B.n575 VSUBS 0.006624f
C647 B.n576 VSUBS 0.006624f
C648 B.n577 VSUBS 0.006624f
C649 B.n578 VSUBS 0.006624f
C650 B.n579 VSUBS 0.006624f
C651 B.n580 VSUBS 0.006624f
C652 B.n581 VSUBS 0.006624f
C653 B.n582 VSUBS 0.006624f
C654 B.n583 VSUBS 0.006624f
C655 B.n584 VSUBS 0.006624f
C656 B.n585 VSUBS 0.006624f
C657 B.n586 VSUBS 0.006624f
C658 B.n587 VSUBS 0.006624f
C659 B.n588 VSUBS 0.006624f
C660 B.n589 VSUBS 0.006624f
C661 B.n590 VSUBS 0.006624f
C662 B.n591 VSUBS 0.006624f
C663 B.n592 VSUBS 0.006624f
C664 B.n593 VSUBS 0.006624f
C665 B.n594 VSUBS 0.006624f
C666 B.n595 VSUBS 0.006624f
C667 B.n596 VSUBS 0.006624f
C668 B.n597 VSUBS 0.006624f
C669 B.n598 VSUBS 0.006624f
C670 B.n599 VSUBS 0.006624f
C671 B.n600 VSUBS 0.006624f
C672 B.n601 VSUBS 0.006624f
C673 B.n602 VSUBS 0.006624f
C674 B.n603 VSUBS 0.006624f
C675 B.n604 VSUBS 0.006624f
C676 B.n605 VSUBS 0.006624f
C677 B.n606 VSUBS 0.006624f
C678 B.n607 VSUBS 0.006624f
C679 B.n608 VSUBS 0.006624f
C680 B.n609 VSUBS 0.006624f
C681 B.n610 VSUBS 0.006624f
C682 B.n611 VSUBS 0.006624f
C683 B.n612 VSUBS 0.006624f
C684 B.n613 VSUBS 0.006624f
C685 B.n614 VSUBS 0.006624f
C686 B.n615 VSUBS 0.006624f
C687 B.n616 VSUBS 0.014532f
C688 B.n617 VSUBS 0.014532f
C689 B.n618 VSUBS 0.013716f
C690 B.n619 VSUBS 0.006624f
C691 B.n620 VSUBS 0.006624f
C692 B.n621 VSUBS 0.006624f
C693 B.n622 VSUBS 0.006624f
C694 B.n623 VSUBS 0.006624f
C695 B.n624 VSUBS 0.006624f
C696 B.n625 VSUBS 0.006624f
C697 B.n626 VSUBS 0.006624f
C698 B.n627 VSUBS 0.006624f
C699 B.n628 VSUBS 0.006624f
C700 B.n629 VSUBS 0.006624f
C701 B.n630 VSUBS 0.006624f
C702 B.n631 VSUBS 0.006624f
C703 B.n632 VSUBS 0.006624f
C704 B.n633 VSUBS 0.006624f
C705 B.n634 VSUBS 0.006624f
C706 B.n635 VSUBS 0.006624f
C707 B.n636 VSUBS 0.006624f
C708 B.n637 VSUBS 0.006624f
C709 B.n638 VSUBS 0.006624f
C710 B.n639 VSUBS 0.006624f
C711 B.n640 VSUBS 0.006624f
C712 B.n641 VSUBS 0.006624f
C713 B.n642 VSUBS 0.006624f
C714 B.n643 VSUBS 0.006624f
C715 B.n644 VSUBS 0.006624f
C716 B.n645 VSUBS 0.006624f
C717 B.n646 VSUBS 0.006624f
C718 B.n647 VSUBS 0.006624f
C719 B.n648 VSUBS 0.006624f
C720 B.n649 VSUBS 0.006624f
C721 B.n650 VSUBS 0.006624f
C722 B.n651 VSUBS 0.006624f
C723 B.n652 VSUBS 0.006624f
C724 B.n653 VSUBS 0.006624f
C725 B.n654 VSUBS 0.006624f
C726 B.n655 VSUBS 0.006624f
C727 B.n656 VSUBS 0.006624f
C728 B.n657 VSUBS 0.006624f
C729 B.n658 VSUBS 0.006624f
C730 B.n659 VSUBS 0.006624f
C731 B.n660 VSUBS 0.006624f
C732 B.n661 VSUBS 0.006624f
C733 B.n662 VSUBS 0.006624f
C734 B.n663 VSUBS 0.006624f
C735 B.n664 VSUBS 0.006624f
C736 B.n665 VSUBS 0.006624f
C737 B.n666 VSUBS 0.006624f
C738 B.n667 VSUBS 0.006624f
C739 B.n668 VSUBS 0.006624f
C740 B.n669 VSUBS 0.006624f
C741 B.n670 VSUBS 0.006624f
C742 B.n671 VSUBS 0.006624f
C743 B.n672 VSUBS 0.006624f
C744 B.n673 VSUBS 0.006624f
C745 B.n674 VSUBS 0.006624f
C746 B.n675 VSUBS 0.006624f
C747 B.n676 VSUBS 0.006624f
C748 B.n677 VSUBS 0.006624f
C749 B.n678 VSUBS 0.006624f
C750 B.n679 VSUBS 0.006624f
C751 B.n680 VSUBS 0.006624f
C752 B.n681 VSUBS 0.006624f
C753 B.n682 VSUBS 0.006624f
C754 B.n683 VSUBS 0.014998f
C755 VTAIL.n0 VSUBS 0.026164f
C756 VTAIL.n1 VSUBS 0.025377f
C757 VTAIL.n2 VSUBS 0.013636f
C758 VTAIL.n3 VSUBS 0.032231f
C759 VTAIL.n4 VSUBS 0.014438f
C760 VTAIL.n5 VSUBS 0.025377f
C761 VTAIL.n6 VSUBS 0.014037f
C762 VTAIL.n7 VSUBS 0.032231f
C763 VTAIL.n8 VSUBS 0.014438f
C764 VTAIL.n9 VSUBS 0.025377f
C765 VTAIL.n10 VSUBS 0.013636f
C766 VTAIL.n11 VSUBS 0.032231f
C767 VTAIL.n12 VSUBS 0.014438f
C768 VTAIL.n13 VSUBS 0.025377f
C769 VTAIL.n14 VSUBS 0.013636f
C770 VTAIL.n15 VSUBS 0.024173f
C771 VTAIL.n16 VSUBS 0.024246f
C772 VTAIL.t4 VSUBS 0.069292f
C773 VTAIL.n17 VSUBS 0.176117f
C774 VTAIL.n18 VSUBS 1.01664f
C775 VTAIL.n19 VSUBS 0.013636f
C776 VTAIL.n20 VSUBS 0.014438f
C777 VTAIL.n21 VSUBS 0.032231f
C778 VTAIL.n22 VSUBS 0.032231f
C779 VTAIL.n23 VSUBS 0.014438f
C780 VTAIL.n24 VSUBS 0.013636f
C781 VTAIL.n25 VSUBS 0.025377f
C782 VTAIL.n26 VSUBS 0.025377f
C783 VTAIL.n27 VSUBS 0.013636f
C784 VTAIL.n28 VSUBS 0.014438f
C785 VTAIL.n29 VSUBS 0.032231f
C786 VTAIL.n30 VSUBS 0.032231f
C787 VTAIL.n31 VSUBS 0.014438f
C788 VTAIL.n32 VSUBS 0.013636f
C789 VTAIL.n33 VSUBS 0.025377f
C790 VTAIL.n34 VSUBS 0.025377f
C791 VTAIL.n35 VSUBS 0.013636f
C792 VTAIL.n36 VSUBS 0.013636f
C793 VTAIL.n37 VSUBS 0.014438f
C794 VTAIL.n38 VSUBS 0.032231f
C795 VTAIL.n39 VSUBS 0.032231f
C796 VTAIL.n40 VSUBS 0.032231f
C797 VTAIL.n41 VSUBS 0.014037f
C798 VTAIL.n42 VSUBS 0.013636f
C799 VTAIL.n43 VSUBS 0.025377f
C800 VTAIL.n44 VSUBS 0.025377f
C801 VTAIL.n45 VSUBS 0.013636f
C802 VTAIL.n46 VSUBS 0.014438f
C803 VTAIL.n47 VSUBS 0.032231f
C804 VTAIL.n48 VSUBS 0.072171f
C805 VTAIL.n49 VSUBS 0.014438f
C806 VTAIL.n50 VSUBS 0.013636f
C807 VTAIL.n51 VSUBS 0.057617f
C808 VTAIL.n52 VSUBS 0.036002f
C809 VTAIL.n53 VSUBS 0.202776f
C810 VTAIL.n54 VSUBS 0.026164f
C811 VTAIL.n55 VSUBS 0.025377f
C812 VTAIL.n56 VSUBS 0.013636f
C813 VTAIL.n57 VSUBS 0.032231f
C814 VTAIL.n58 VSUBS 0.014438f
C815 VTAIL.n59 VSUBS 0.025377f
C816 VTAIL.n60 VSUBS 0.014037f
C817 VTAIL.n61 VSUBS 0.032231f
C818 VTAIL.n62 VSUBS 0.014438f
C819 VTAIL.n63 VSUBS 0.025377f
C820 VTAIL.n64 VSUBS 0.013636f
C821 VTAIL.n65 VSUBS 0.032231f
C822 VTAIL.n66 VSUBS 0.014438f
C823 VTAIL.n67 VSUBS 0.025377f
C824 VTAIL.n68 VSUBS 0.013636f
C825 VTAIL.n69 VSUBS 0.024173f
C826 VTAIL.n70 VSUBS 0.024246f
C827 VTAIL.t6 VSUBS 0.069292f
C828 VTAIL.n71 VSUBS 0.176117f
C829 VTAIL.n72 VSUBS 1.01664f
C830 VTAIL.n73 VSUBS 0.013636f
C831 VTAIL.n74 VSUBS 0.014438f
C832 VTAIL.n75 VSUBS 0.032231f
C833 VTAIL.n76 VSUBS 0.032231f
C834 VTAIL.n77 VSUBS 0.014438f
C835 VTAIL.n78 VSUBS 0.013636f
C836 VTAIL.n79 VSUBS 0.025377f
C837 VTAIL.n80 VSUBS 0.025377f
C838 VTAIL.n81 VSUBS 0.013636f
C839 VTAIL.n82 VSUBS 0.014438f
C840 VTAIL.n83 VSUBS 0.032231f
C841 VTAIL.n84 VSUBS 0.032231f
C842 VTAIL.n85 VSUBS 0.014438f
C843 VTAIL.n86 VSUBS 0.013636f
C844 VTAIL.n87 VSUBS 0.025377f
C845 VTAIL.n88 VSUBS 0.025377f
C846 VTAIL.n89 VSUBS 0.013636f
C847 VTAIL.n90 VSUBS 0.013636f
C848 VTAIL.n91 VSUBS 0.014438f
C849 VTAIL.n92 VSUBS 0.032231f
C850 VTAIL.n93 VSUBS 0.032231f
C851 VTAIL.n94 VSUBS 0.032231f
C852 VTAIL.n95 VSUBS 0.014037f
C853 VTAIL.n96 VSUBS 0.013636f
C854 VTAIL.n97 VSUBS 0.025377f
C855 VTAIL.n98 VSUBS 0.025377f
C856 VTAIL.n99 VSUBS 0.013636f
C857 VTAIL.n100 VSUBS 0.014438f
C858 VTAIL.n101 VSUBS 0.032231f
C859 VTAIL.n102 VSUBS 0.072171f
C860 VTAIL.n103 VSUBS 0.014438f
C861 VTAIL.n104 VSUBS 0.013636f
C862 VTAIL.n105 VSUBS 0.057617f
C863 VTAIL.n106 VSUBS 0.036002f
C864 VTAIL.n107 VSUBS 0.336532f
C865 VTAIL.n108 VSUBS 0.026164f
C866 VTAIL.n109 VSUBS 0.025377f
C867 VTAIL.n110 VSUBS 0.013636f
C868 VTAIL.n111 VSUBS 0.032231f
C869 VTAIL.n112 VSUBS 0.014438f
C870 VTAIL.n113 VSUBS 0.025377f
C871 VTAIL.n114 VSUBS 0.014037f
C872 VTAIL.n115 VSUBS 0.032231f
C873 VTAIL.n116 VSUBS 0.014438f
C874 VTAIL.n117 VSUBS 0.025377f
C875 VTAIL.n118 VSUBS 0.013636f
C876 VTAIL.n119 VSUBS 0.032231f
C877 VTAIL.n120 VSUBS 0.014438f
C878 VTAIL.n121 VSUBS 0.025377f
C879 VTAIL.n122 VSUBS 0.013636f
C880 VTAIL.n123 VSUBS 0.024173f
C881 VTAIL.n124 VSUBS 0.024246f
C882 VTAIL.t5 VSUBS 0.069292f
C883 VTAIL.n125 VSUBS 0.176117f
C884 VTAIL.n126 VSUBS 1.01664f
C885 VTAIL.n127 VSUBS 0.013636f
C886 VTAIL.n128 VSUBS 0.014438f
C887 VTAIL.n129 VSUBS 0.032231f
C888 VTAIL.n130 VSUBS 0.032231f
C889 VTAIL.n131 VSUBS 0.014438f
C890 VTAIL.n132 VSUBS 0.013636f
C891 VTAIL.n133 VSUBS 0.025377f
C892 VTAIL.n134 VSUBS 0.025377f
C893 VTAIL.n135 VSUBS 0.013636f
C894 VTAIL.n136 VSUBS 0.014438f
C895 VTAIL.n137 VSUBS 0.032231f
C896 VTAIL.n138 VSUBS 0.032231f
C897 VTAIL.n139 VSUBS 0.014438f
C898 VTAIL.n140 VSUBS 0.013636f
C899 VTAIL.n141 VSUBS 0.025377f
C900 VTAIL.n142 VSUBS 0.025377f
C901 VTAIL.n143 VSUBS 0.013636f
C902 VTAIL.n144 VSUBS 0.013636f
C903 VTAIL.n145 VSUBS 0.014438f
C904 VTAIL.n146 VSUBS 0.032231f
C905 VTAIL.n147 VSUBS 0.032231f
C906 VTAIL.n148 VSUBS 0.032231f
C907 VTAIL.n149 VSUBS 0.014037f
C908 VTAIL.n150 VSUBS 0.013636f
C909 VTAIL.n151 VSUBS 0.025377f
C910 VTAIL.n152 VSUBS 0.025377f
C911 VTAIL.n153 VSUBS 0.013636f
C912 VTAIL.n154 VSUBS 0.014438f
C913 VTAIL.n155 VSUBS 0.032231f
C914 VTAIL.n156 VSUBS 0.072171f
C915 VTAIL.n157 VSUBS 0.014438f
C916 VTAIL.n158 VSUBS 0.013636f
C917 VTAIL.n159 VSUBS 0.057617f
C918 VTAIL.n160 VSUBS 0.036002f
C919 VTAIL.n161 VSUBS 1.61982f
C920 VTAIL.n162 VSUBS 0.026164f
C921 VTAIL.n163 VSUBS 0.025377f
C922 VTAIL.n164 VSUBS 0.013636f
C923 VTAIL.n165 VSUBS 0.032231f
C924 VTAIL.n166 VSUBS 0.014438f
C925 VTAIL.n167 VSUBS 0.025377f
C926 VTAIL.n168 VSUBS 0.014037f
C927 VTAIL.n169 VSUBS 0.032231f
C928 VTAIL.n170 VSUBS 0.013636f
C929 VTAIL.n171 VSUBS 0.014438f
C930 VTAIL.n172 VSUBS 0.025377f
C931 VTAIL.n173 VSUBS 0.013636f
C932 VTAIL.n174 VSUBS 0.032231f
C933 VTAIL.n175 VSUBS 0.014438f
C934 VTAIL.n176 VSUBS 0.025377f
C935 VTAIL.n177 VSUBS 0.013636f
C936 VTAIL.n178 VSUBS 0.024173f
C937 VTAIL.n179 VSUBS 0.024246f
C938 VTAIL.t2 VSUBS 0.069292f
C939 VTAIL.n180 VSUBS 0.176117f
C940 VTAIL.n181 VSUBS 1.01664f
C941 VTAIL.n182 VSUBS 0.013636f
C942 VTAIL.n183 VSUBS 0.014438f
C943 VTAIL.n184 VSUBS 0.032231f
C944 VTAIL.n185 VSUBS 0.032231f
C945 VTAIL.n186 VSUBS 0.014438f
C946 VTAIL.n187 VSUBS 0.013636f
C947 VTAIL.n188 VSUBS 0.025377f
C948 VTAIL.n189 VSUBS 0.025377f
C949 VTAIL.n190 VSUBS 0.013636f
C950 VTAIL.n191 VSUBS 0.014438f
C951 VTAIL.n192 VSUBS 0.032231f
C952 VTAIL.n193 VSUBS 0.032231f
C953 VTAIL.n194 VSUBS 0.014438f
C954 VTAIL.n195 VSUBS 0.013636f
C955 VTAIL.n196 VSUBS 0.025377f
C956 VTAIL.n197 VSUBS 0.025377f
C957 VTAIL.n198 VSUBS 0.013636f
C958 VTAIL.n199 VSUBS 0.014438f
C959 VTAIL.n200 VSUBS 0.032231f
C960 VTAIL.n201 VSUBS 0.032231f
C961 VTAIL.n202 VSUBS 0.032231f
C962 VTAIL.n203 VSUBS 0.014037f
C963 VTAIL.n204 VSUBS 0.013636f
C964 VTAIL.n205 VSUBS 0.025377f
C965 VTAIL.n206 VSUBS 0.025377f
C966 VTAIL.n207 VSUBS 0.013636f
C967 VTAIL.n208 VSUBS 0.014438f
C968 VTAIL.n209 VSUBS 0.032231f
C969 VTAIL.n210 VSUBS 0.072171f
C970 VTAIL.n211 VSUBS 0.014438f
C971 VTAIL.n212 VSUBS 0.013636f
C972 VTAIL.n213 VSUBS 0.057617f
C973 VTAIL.n214 VSUBS 0.036002f
C974 VTAIL.n215 VSUBS 1.61982f
C975 VTAIL.n216 VSUBS 0.026164f
C976 VTAIL.n217 VSUBS 0.025377f
C977 VTAIL.n218 VSUBS 0.013636f
C978 VTAIL.n219 VSUBS 0.032231f
C979 VTAIL.n220 VSUBS 0.014438f
C980 VTAIL.n221 VSUBS 0.025377f
C981 VTAIL.n222 VSUBS 0.014037f
C982 VTAIL.n223 VSUBS 0.032231f
C983 VTAIL.n224 VSUBS 0.013636f
C984 VTAIL.n225 VSUBS 0.014438f
C985 VTAIL.n226 VSUBS 0.025377f
C986 VTAIL.n227 VSUBS 0.013636f
C987 VTAIL.n228 VSUBS 0.032231f
C988 VTAIL.n229 VSUBS 0.014438f
C989 VTAIL.n230 VSUBS 0.025377f
C990 VTAIL.n231 VSUBS 0.013636f
C991 VTAIL.n232 VSUBS 0.024173f
C992 VTAIL.n233 VSUBS 0.024246f
C993 VTAIL.t3 VSUBS 0.069292f
C994 VTAIL.n234 VSUBS 0.176117f
C995 VTAIL.n235 VSUBS 1.01664f
C996 VTAIL.n236 VSUBS 0.013636f
C997 VTAIL.n237 VSUBS 0.014438f
C998 VTAIL.n238 VSUBS 0.032231f
C999 VTAIL.n239 VSUBS 0.032231f
C1000 VTAIL.n240 VSUBS 0.014438f
C1001 VTAIL.n241 VSUBS 0.013636f
C1002 VTAIL.n242 VSUBS 0.025377f
C1003 VTAIL.n243 VSUBS 0.025377f
C1004 VTAIL.n244 VSUBS 0.013636f
C1005 VTAIL.n245 VSUBS 0.014438f
C1006 VTAIL.n246 VSUBS 0.032231f
C1007 VTAIL.n247 VSUBS 0.032231f
C1008 VTAIL.n248 VSUBS 0.014438f
C1009 VTAIL.n249 VSUBS 0.013636f
C1010 VTAIL.n250 VSUBS 0.025377f
C1011 VTAIL.n251 VSUBS 0.025377f
C1012 VTAIL.n252 VSUBS 0.013636f
C1013 VTAIL.n253 VSUBS 0.014438f
C1014 VTAIL.n254 VSUBS 0.032231f
C1015 VTAIL.n255 VSUBS 0.032231f
C1016 VTAIL.n256 VSUBS 0.032231f
C1017 VTAIL.n257 VSUBS 0.014037f
C1018 VTAIL.n258 VSUBS 0.013636f
C1019 VTAIL.n259 VSUBS 0.025377f
C1020 VTAIL.n260 VSUBS 0.025377f
C1021 VTAIL.n261 VSUBS 0.013636f
C1022 VTAIL.n262 VSUBS 0.014438f
C1023 VTAIL.n263 VSUBS 0.032231f
C1024 VTAIL.n264 VSUBS 0.072171f
C1025 VTAIL.n265 VSUBS 0.014438f
C1026 VTAIL.n266 VSUBS 0.013636f
C1027 VTAIL.n267 VSUBS 0.057617f
C1028 VTAIL.n268 VSUBS 0.036002f
C1029 VTAIL.n269 VSUBS 0.336532f
C1030 VTAIL.n270 VSUBS 0.026164f
C1031 VTAIL.n271 VSUBS 0.025377f
C1032 VTAIL.n272 VSUBS 0.013636f
C1033 VTAIL.n273 VSUBS 0.032231f
C1034 VTAIL.n274 VSUBS 0.014438f
C1035 VTAIL.n275 VSUBS 0.025377f
C1036 VTAIL.n276 VSUBS 0.014037f
C1037 VTAIL.n277 VSUBS 0.032231f
C1038 VTAIL.n278 VSUBS 0.013636f
C1039 VTAIL.n279 VSUBS 0.014438f
C1040 VTAIL.n280 VSUBS 0.025377f
C1041 VTAIL.n281 VSUBS 0.013636f
C1042 VTAIL.n282 VSUBS 0.032231f
C1043 VTAIL.n283 VSUBS 0.014438f
C1044 VTAIL.n284 VSUBS 0.025377f
C1045 VTAIL.n285 VSUBS 0.013636f
C1046 VTAIL.n286 VSUBS 0.024173f
C1047 VTAIL.n287 VSUBS 0.024246f
C1048 VTAIL.t7 VSUBS 0.069292f
C1049 VTAIL.n288 VSUBS 0.176117f
C1050 VTAIL.n289 VSUBS 1.01664f
C1051 VTAIL.n290 VSUBS 0.013636f
C1052 VTAIL.n291 VSUBS 0.014438f
C1053 VTAIL.n292 VSUBS 0.032231f
C1054 VTAIL.n293 VSUBS 0.032231f
C1055 VTAIL.n294 VSUBS 0.014438f
C1056 VTAIL.n295 VSUBS 0.013636f
C1057 VTAIL.n296 VSUBS 0.025377f
C1058 VTAIL.n297 VSUBS 0.025377f
C1059 VTAIL.n298 VSUBS 0.013636f
C1060 VTAIL.n299 VSUBS 0.014438f
C1061 VTAIL.n300 VSUBS 0.032231f
C1062 VTAIL.n301 VSUBS 0.032231f
C1063 VTAIL.n302 VSUBS 0.014438f
C1064 VTAIL.n303 VSUBS 0.013636f
C1065 VTAIL.n304 VSUBS 0.025377f
C1066 VTAIL.n305 VSUBS 0.025377f
C1067 VTAIL.n306 VSUBS 0.013636f
C1068 VTAIL.n307 VSUBS 0.014438f
C1069 VTAIL.n308 VSUBS 0.032231f
C1070 VTAIL.n309 VSUBS 0.032231f
C1071 VTAIL.n310 VSUBS 0.032231f
C1072 VTAIL.n311 VSUBS 0.014037f
C1073 VTAIL.n312 VSUBS 0.013636f
C1074 VTAIL.n313 VSUBS 0.025377f
C1075 VTAIL.n314 VSUBS 0.025377f
C1076 VTAIL.n315 VSUBS 0.013636f
C1077 VTAIL.n316 VSUBS 0.014438f
C1078 VTAIL.n317 VSUBS 0.032231f
C1079 VTAIL.n318 VSUBS 0.072171f
C1080 VTAIL.n319 VSUBS 0.014438f
C1081 VTAIL.n320 VSUBS 0.013636f
C1082 VTAIL.n321 VSUBS 0.057617f
C1083 VTAIL.n322 VSUBS 0.036002f
C1084 VTAIL.n323 VSUBS 0.336532f
C1085 VTAIL.n324 VSUBS 0.026164f
C1086 VTAIL.n325 VSUBS 0.025377f
C1087 VTAIL.n326 VSUBS 0.013636f
C1088 VTAIL.n327 VSUBS 0.032231f
C1089 VTAIL.n328 VSUBS 0.014438f
C1090 VTAIL.n329 VSUBS 0.025377f
C1091 VTAIL.n330 VSUBS 0.014037f
C1092 VTAIL.n331 VSUBS 0.032231f
C1093 VTAIL.n332 VSUBS 0.013636f
C1094 VTAIL.n333 VSUBS 0.014438f
C1095 VTAIL.n334 VSUBS 0.025377f
C1096 VTAIL.n335 VSUBS 0.013636f
C1097 VTAIL.n336 VSUBS 0.032231f
C1098 VTAIL.n337 VSUBS 0.014438f
C1099 VTAIL.n338 VSUBS 0.025377f
C1100 VTAIL.n339 VSUBS 0.013636f
C1101 VTAIL.n340 VSUBS 0.024173f
C1102 VTAIL.n341 VSUBS 0.024246f
C1103 VTAIL.t0 VSUBS 0.069292f
C1104 VTAIL.n342 VSUBS 0.176117f
C1105 VTAIL.n343 VSUBS 1.01664f
C1106 VTAIL.n344 VSUBS 0.013636f
C1107 VTAIL.n345 VSUBS 0.014438f
C1108 VTAIL.n346 VSUBS 0.032231f
C1109 VTAIL.n347 VSUBS 0.032231f
C1110 VTAIL.n348 VSUBS 0.014438f
C1111 VTAIL.n349 VSUBS 0.013636f
C1112 VTAIL.n350 VSUBS 0.025377f
C1113 VTAIL.n351 VSUBS 0.025377f
C1114 VTAIL.n352 VSUBS 0.013636f
C1115 VTAIL.n353 VSUBS 0.014438f
C1116 VTAIL.n354 VSUBS 0.032231f
C1117 VTAIL.n355 VSUBS 0.032231f
C1118 VTAIL.n356 VSUBS 0.014438f
C1119 VTAIL.n357 VSUBS 0.013636f
C1120 VTAIL.n358 VSUBS 0.025377f
C1121 VTAIL.n359 VSUBS 0.025377f
C1122 VTAIL.n360 VSUBS 0.013636f
C1123 VTAIL.n361 VSUBS 0.014438f
C1124 VTAIL.n362 VSUBS 0.032231f
C1125 VTAIL.n363 VSUBS 0.032231f
C1126 VTAIL.n364 VSUBS 0.032231f
C1127 VTAIL.n365 VSUBS 0.014037f
C1128 VTAIL.n366 VSUBS 0.013636f
C1129 VTAIL.n367 VSUBS 0.025377f
C1130 VTAIL.n368 VSUBS 0.025377f
C1131 VTAIL.n369 VSUBS 0.013636f
C1132 VTAIL.n370 VSUBS 0.014438f
C1133 VTAIL.n371 VSUBS 0.032231f
C1134 VTAIL.n372 VSUBS 0.072171f
C1135 VTAIL.n373 VSUBS 0.014438f
C1136 VTAIL.n374 VSUBS 0.013636f
C1137 VTAIL.n375 VSUBS 0.057617f
C1138 VTAIL.n376 VSUBS 0.036002f
C1139 VTAIL.n377 VSUBS 1.61982f
C1140 VTAIL.n378 VSUBS 0.026164f
C1141 VTAIL.n379 VSUBS 0.025377f
C1142 VTAIL.n380 VSUBS 0.013636f
C1143 VTAIL.n381 VSUBS 0.032231f
C1144 VTAIL.n382 VSUBS 0.014438f
C1145 VTAIL.n383 VSUBS 0.025377f
C1146 VTAIL.n384 VSUBS 0.014037f
C1147 VTAIL.n385 VSUBS 0.032231f
C1148 VTAIL.n386 VSUBS 0.014438f
C1149 VTAIL.n387 VSUBS 0.025377f
C1150 VTAIL.n388 VSUBS 0.013636f
C1151 VTAIL.n389 VSUBS 0.032231f
C1152 VTAIL.n390 VSUBS 0.014438f
C1153 VTAIL.n391 VSUBS 0.025377f
C1154 VTAIL.n392 VSUBS 0.013636f
C1155 VTAIL.n393 VSUBS 0.024173f
C1156 VTAIL.n394 VSUBS 0.024246f
C1157 VTAIL.t1 VSUBS 0.069292f
C1158 VTAIL.n395 VSUBS 0.176117f
C1159 VTAIL.n396 VSUBS 1.01664f
C1160 VTAIL.n397 VSUBS 0.013636f
C1161 VTAIL.n398 VSUBS 0.014438f
C1162 VTAIL.n399 VSUBS 0.032231f
C1163 VTAIL.n400 VSUBS 0.032231f
C1164 VTAIL.n401 VSUBS 0.014438f
C1165 VTAIL.n402 VSUBS 0.013636f
C1166 VTAIL.n403 VSUBS 0.025377f
C1167 VTAIL.n404 VSUBS 0.025377f
C1168 VTAIL.n405 VSUBS 0.013636f
C1169 VTAIL.n406 VSUBS 0.014438f
C1170 VTAIL.n407 VSUBS 0.032231f
C1171 VTAIL.n408 VSUBS 0.032231f
C1172 VTAIL.n409 VSUBS 0.014438f
C1173 VTAIL.n410 VSUBS 0.013636f
C1174 VTAIL.n411 VSUBS 0.025377f
C1175 VTAIL.n412 VSUBS 0.025377f
C1176 VTAIL.n413 VSUBS 0.013636f
C1177 VTAIL.n414 VSUBS 0.013636f
C1178 VTAIL.n415 VSUBS 0.014438f
C1179 VTAIL.n416 VSUBS 0.032231f
C1180 VTAIL.n417 VSUBS 0.032231f
C1181 VTAIL.n418 VSUBS 0.032231f
C1182 VTAIL.n419 VSUBS 0.014037f
C1183 VTAIL.n420 VSUBS 0.013636f
C1184 VTAIL.n421 VSUBS 0.025377f
C1185 VTAIL.n422 VSUBS 0.025377f
C1186 VTAIL.n423 VSUBS 0.013636f
C1187 VTAIL.n424 VSUBS 0.014438f
C1188 VTAIL.n425 VSUBS 0.032231f
C1189 VTAIL.n426 VSUBS 0.072171f
C1190 VTAIL.n427 VSUBS 0.014438f
C1191 VTAIL.n428 VSUBS 0.013636f
C1192 VTAIL.n429 VSUBS 0.057617f
C1193 VTAIL.n430 VSUBS 0.036002f
C1194 VTAIL.n431 VSUBS 1.47655f
C1195 VDD2.t2 VSUBS 0.215942f
C1196 VDD2.t1 VSUBS 0.215942f
C1197 VDD2.n0 VSUBS 2.3087f
C1198 VDD2.t3 VSUBS 0.215942f
C1199 VDD2.t0 VSUBS 0.215942f
C1200 VDD2.n1 VSUBS 1.62614f
C1201 VDD2.n2 VSUBS 4.39505f
C1202 VN.t3 VSUBS 3.26903f
C1203 VN.t0 VSUBS 3.28358f
C1204 VN.n0 VSUBS 1.93204f
C1205 VN.t1 VSUBS 3.28358f
C1206 VN.t2 VSUBS 3.26903f
C1207 VN.n1 VSUBS 3.75671f
.ends

