* NGSPICE file created from diff_pair_sample_0579.ext - technology: sky130A

.subckt diff_pair_sample_0579 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.07
X1 VDD2.t9 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.07
X2 VDD1.t8 VP.t1 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X3 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.07
X4 VDD1.t7 VP.t2 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.07
X5 VTAIL.t16 VP.t3 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X6 VTAIL.t11 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X7 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.07
X9 VDD2.t7 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.07
X10 VDD2.t6 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=4.2627 ps=22.64 w=10.93 l=2.07
X11 VTAIL.t8 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X12 VTAIL.t0 VN.t5 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X13 VDD1.t4 VP.t5 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X14 VTAIL.t13 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X15 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X16 VDD1.t2 VP.t7 VTAIL.t19 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.07
X17 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.07
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=0 ps=0 w=10.93 l=2.07
X19 VTAIL.t5 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X20 VDD2.t1 VN.t8 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.07
X21 VDD1.t1 VP.t8 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=4.2627 pd=22.64 as=1.80345 ps=11.26 w=10.93 l=2.07
X22 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
X23 VTAIL.t15 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.80345 pd=11.26 as=1.80345 ps=11.26 w=10.93 l=2.07
R0 VP.n20 VP.n19 161.3
R1 VP.n21 VP.n16 161.3
R2 VP.n23 VP.n22 161.3
R3 VP.n24 VP.n15 161.3
R4 VP.n26 VP.n25 161.3
R5 VP.n27 VP.n14 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n13 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n34 VP.n12 161.3
R10 VP.n36 VP.n35 161.3
R11 VP.n37 VP.n11 161.3
R12 VP.n39 VP.n38 161.3
R13 VP.n40 VP.n10 161.3
R14 VP.n74 VP.n0 161.3
R15 VP.n73 VP.n72 161.3
R16 VP.n71 VP.n1 161.3
R17 VP.n70 VP.n69 161.3
R18 VP.n68 VP.n2 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n3 161.3
R21 VP.n63 VP.n62 161.3
R22 VP.n61 VP.n4 161.3
R23 VP.n60 VP.n59 161.3
R24 VP.n58 VP.n5 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n6 161.3
R27 VP.n54 VP.n53 161.3
R28 VP.n52 VP.n51 161.3
R29 VP.n50 VP.n8 161.3
R30 VP.n49 VP.n48 161.3
R31 VP.n47 VP.n9 161.3
R32 VP.n46 VP.n45 161.3
R33 VP.n18 VP.t7 160.191
R34 VP.n60 VP.t1 127.254
R35 VP.n44 VP.t8 127.254
R36 VP.n7 VP.t9 127.254
R37 VP.n67 VP.t3 127.254
R38 VP.n75 VP.t2 127.254
R39 VP.n26 VP.t5 127.254
R40 VP.n41 VP.t0 127.254
R41 VP.n33 VP.t4 127.254
R42 VP.n17 VP.t6 127.254
R43 VP.n44 VP.n43 96.0763
R44 VP.n76 VP.n75 96.0763
R45 VP.n42 VP.n41 96.0763
R46 VP.n56 VP.n55 56.5193
R47 VP.n62 VP.n3 56.5193
R48 VP.n28 VP.n13 56.5193
R49 VP.n22 VP.n21 56.5193
R50 VP.n18 VP.n17 51.1767
R51 VP.n49 VP.n9 50.2061
R52 VP.n73 VP.n1 50.2061
R53 VP.n39 VP.n11 50.2061
R54 VP.n43 VP.n42 49.386
R55 VP.n50 VP.n49 30.7807
R56 VP.n69 VP.n1 30.7807
R57 VP.n35 VP.n11 30.7807
R58 VP.n45 VP.n9 24.4675
R59 VP.n51 VP.n50 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n5 24.4675
R62 VP.n60 VP.n5 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n62 VP.n61 24.4675
R65 VP.n66 VP.n3 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n74 VP.n73 24.4675
R68 VP.n40 VP.n39 24.4675
R69 VP.n32 VP.n13 24.4675
R70 VP.n35 VP.n34 24.4675
R71 VP.n22 VP.n15 24.4675
R72 VP.n26 VP.n15 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 19.5741
R77 VP.n67 VP.n66 19.5741
R78 VP.n33 VP.n32 19.5741
R79 VP.n20 VP.n17 19.5741
R80 VP.n45 VP.n44 14.6807
R81 VP.n75 VP.n74 14.6807
R82 VP.n41 VP.n40 14.6807
R83 VP.n19 VP.n18 9.46762
R84 VP.n51 VP.n7 4.8939
R85 VP.n68 VP.n67 4.8939
R86 VP.n34 VP.n33 4.8939
R87 VP.n42 VP.n10 0.278367
R88 VP.n46 VP.n43 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153454
R122 VTAIL.n11 VTAIL.t1 45.2085
R123 VTAIL.n17 VTAIL.t7 45.2084
R124 VTAIL.n2 VTAIL.t12 45.2084
R125 VTAIL.n16 VTAIL.t18 45.2084
R126 VTAIL.n15 VTAIL.n14 43.397
R127 VTAIL.n13 VTAIL.n12 43.397
R128 VTAIL.n10 VTAIL.n9 43.397
R129 VTAIL.n8 VTAIL.n7 43.397
R130 VTAIL.n19 VTAIL.n18 43.3968
R131 VTAIL.n1 VTAIL.n0 43.3968
R132 VTAIL.n4 VTAIL.n3 43.3968
R133 VTAIL.n6 VTAIL.n5 43.3968
R134 VTAIL.n8 VTAIL.n6 25.9272
R135 VTAIL.n17 VTAIL.n16 23.8583
R136 VTAIL.n10 VTAIL.n8 2.06947
R137 VTAIL.n11 VTAIL.n10 2.06947
R138 VTAIL.n15 VTAIL.n13 2.06947
R139 VTAIL.n16 VTAIL.n15 2.06947
R140 VTAIL.n6 VTAIL.n4 2.06947
R141 VTAIL.n4 VTAIL.n2 2.06947
R142 VTAIL.n19 VTAIL.n17 2.06947
R143 VTAIL.n18 VTAIL.t9 1.81203
R144 VTAIL.n18 VTAIL.t0 1.81203
R145 VTAIL.n0 VTAIL.t4 1.81203
R146 VTAIL.n0 VTAIL.t5 1.81203
R147 VTAIL.n3 VTAIL.t10 1.81203
R148 VTAIL.n3 VTAIL.t16 1.81203
R149 VTAIL.n5 VTAIL.t17 1.81203
R150 VTAIL.n5 VTAIL.t15 1.81203
R151 VTAIL.n14 VTAIL.t14 1.81203
R152 VTAIL.n14 VTAIL.t11 1.81203
R153 VTAIL.n12 VTAIL.t19 1.81203
R154 VTAIL.n12 VTAIL.t13 1.81203
R155 VTAIL.n9 VTAIL.t6 1.81203
R156 VTAIL.n9 VTAIL.t8 1.81203
R157 VTAIL.n7 VTAIL.t3 1.81203
R158 VTAIL.n7 VTAIL.t2 1.81203
R159 VTAIL VTAIL.n1 1.61041
R160 VTAIL.n13 VTAIL.n11 1.50481
R161 VTAIL.n2 VTAIL.n1 1.50481
R162 VTAIL VTAIL.n19 0.459552
R163 VDD1.n1 VDD1.t2 63.9562
R164 VDD1.n3 VDD1.t1 63.9561
R165 VDD1.n5 VDD1.n4 61.572
R166 VDD1.n1 VDD1.n0 60.0758
R167 VDD1.n7 VDD1.n6 60.0756
R168 VDD1.n3 VDD1.n2 60.0756
R169 VDD1.n7 VDD1.n5 44.5828
R170 VDD1.n6 VDD1.t5 1.81203
R171 VDD1.n6 VDD1.t9 1.81203
R172 VDD1.n0 VDD1.t3 1.81203
R173 VDD1.n0 VDD1.t4 1.81203
R174 VDD1.n4 VDD1.t6 1.81203
R175 VDD1.n4 VDD1.t7 1.81203
R176 VDD1.n2 VDD1.t0 1.81203
R177 VDD1.n2 VDD1.t8 1.81203
R178 VDD1 VDD1.n7 1.49403
R179 VDD1 VDD1.n1 0.575931
R180 VDD1.n5 VDD1.n3 0.462395
R181 B.n679 B.n678 585
R182 B.n679 B.n93 585
R183 B.n682 B.n681 585
R184 B.n683 B.n141 585
R185 B.n685 B.n684 585
R186 B.n687 B.n140 585
R187 B.n690 B.n689 585
R188 B.n691 B.n139 585
R189 B.n693 B.n692 585
R190 B.n695 B.n138 585
R191 B.n698 B.n697 585
R192 B.n699 B.n137 585
R193 B.n701 B.n700 585
R194 B.n703 B.n136 585
R195 B.n706 B.n705 585
R196 B.n707 B.n135 585
R197 B.n709 B.n708 585
R198 B.n711 B.n134 585
R199 B.n714 B.n713 585
R200 B.n715 B.n133 585
R201 B.n717 B.n716 585
R202 B.n719 B.n132 585
R203 B.n722 B.n721 585
R204 B.n723 B.n131 585
R205 B.n725 B.n724 585
R206 B.n727 B.n130 585
R207 B.n730 B.n729 585
R208 B.n731 B.n129 585
R209 B.n733 B.n732 585
R210 B.n735 B.n128 585
R211 B.n738 B.n737 585
R212 B.n739 B.n127 585
R213 B.n741 B.n740 585
R214 B.n743 B.n126 585
R215 B.n746 B.n745 585
R216 B.n747 B.n125 585
R217 B.n749 B.n748 585
R218 B.n751 B.n124 585
R219 B.n754 B.n753 585
R220 B.n755 B.n121 585
R221 B.n758 B.n757 585
R222 B.n760 B.n120 585
R223 B.n763 B.n762 585
R224 B.n764 B.n119 585
R225 B.n766 B.n765 585
R226 B.n768 B.n118 585
R227 B.n771 B.n770 585
R228 B.n772 B.n114 585
R229 B.n774 B.n773 585
R230 B.n776 B.n113 585
R231 B.n779 B.n778 585
R232 B.n780 B.n112 585
R233 B.n782 B.n781 585
R234 B.n784 B.n111 585
R235 B.n787 B.n786 585
R236 B.n788 B.n110 585
R237 B.n790 B.n789 585
R238 B.n792 B.n109 585
R239 B.n795 B.n794 585
R240 B.n796 B.n108 585
R241 B.n798 B.n797 585
R242 B.n800 B.n107 585
R243 B.n803 B.n802 585
R244 B.n804 B.n106 585
R245 B.n806 B.n805 585
R246 B.n808 B.n105 585
R247 B.n811 B.n810 585
R248 B.n812 B.n104 585
R249 B.n814 B.n813 585
R250 B.n816 B.n103 585
R251 B.n819 B.n818 585
R252 B.n820 B.n102 585
R253 B.n822 B.n821 585
R254 B.n824 B.n101 585
R255 B.n827 B.n826 585
R256 B.n828 B.n100 585
R257 B.n830 B.n829 585
R258 B.n832 B.n99 585
R259 B.n835 B.n834 585
R260 B.n836 B.n98 585
R261 B.n838 B.n837 585
R262 B.n840 B.n97 585
R263 B.n843 B.n842 585
R264 B.n844 B.n96 585
R265 B.n846 B.n845 585
R266 B.n848 B.n95 585
R267 B.n851 B.n850 585
R268 B.n852 B.n94 585
R269 B.n677 B.n92 585
R270 B.n855 B.n92 585
R271 B.n676 B.n91 585
R272 B.n856 B.n91 585
R273 B.n675 B.n90 585
R274 B.n857 B.n90 585
R275 B.n674 B.n673 585
R276 B.n673 B.n86 585
R277 B.n672 B.n85 585
R278 B.n863 B.n85 585
R279 B.n671 B.n84 585
R280 B.n864 B.n84 585
R281 B.n670 B.n83 585
R282 B.n865 B.n83 585
R283 B.n669 B.n668 585
R284 B.n668 B.n79 585
R285 B.n667 B.n78 585
R286 B.n871 B.n78 585
R287 B.n666 B.n77 585
R288 B.n872 B.n77 585
R289 B.n665 B.n76 585
R290 B.n873 B.n76 585
R291 B.n664 B.n663 585
R292 B.n663 B.n72 585
R293 B.n662 B.n71 585
R294 B.n879 B.n71 585
R295 B.n661 B.n70 585
R296 B.n880 B.n70 585
R297 B.n660 B.n69 585
R298 B.n881 B.n69 585
R299 B.n659 B.n658 585
R300 B.n658 B.n65 585
R301 B.n657 B.n64 585
R302 B.n887 B.n64 585
R303 B.n656 B.n63 585
R304 B.n888 B.n63 585
R305 B.n655 B.n62 585
R306 B.n889 B.n62 585
R307 B.n654 B.n653 585
R308 B.n653 B.n58 585
R309 B.n652 B.n57 585
R310 B.n895 B.n57 585
R311 B.n651 B.n56 585
R312 B.n896 B.n56 585
R313 B.n650 B.n55 585
R314 B.n897 B.n55 585
R315 B.n649 B.n648 585
R316 B.n648 B.n51 585
R317 B.n647 B.n50 585
R318 B.n903 B.n50 585
R319 B.n646 B.n49 585
R320 B.n904 B.n49 585
R321 B.n645 B.n48 585
R322 B.n905 B.n48 585
R323 B.n644 B.n643 585
R324 B.n643 B.n44 585
R325 B.n642 B.n43 585
R326 B.n911 B.n43 585
R327 B.n641 B.n42 585
R328 B.n912 B.n42 585
R329 B.n640 B.n41 585
R330 B.n913 B.n41 585
R331 B.n639 B.n638 585
R332 B.n638 B.n40 585
R333 B.n637 B.n36 585
R334 B.n919 B.n36 585
R335 B.n636 B.n35 585
R336 B.n920 B.n35 585
R337 B.n635 B.n34 585
R338 B.n921 B.n34 585
R339 B.n634 B.n633 585
R340 B.n633 B.n30 585
R341 B.n632 B.n29 585
R342 B.n927 B.n29 585
R343 B.n631 B.n28 585
R344 B.n928 B.n28 585
R345 B.n630 B.n27 585
R346 B.n929 B.n27 585
R347 B.n629 B.n628 585
R348 B.n628 B.n23 585
R349 B.n627 B.n22 585
R350 B.n935 B.n22 585
R351 B.n626 B.n21 585
R352 B.n936 B.n21 585
R353 B.n625 B.n20 585
R354 B.n937 B.n20 585
R355 B.n624 B.n623 585
R356 B.n623 B.n16 585
R357 B.n622 B.n15 585
R358 B.n943 B.n15 585
R359 B.n621 B.n14 585
R360 B.n944 B.n14 585
R361 B.n620 B.n13 585
R362 B.n945 B.n13 585
R363 B.n619 B.n618 585
R364 B.n618 B.n12 585
R365 B.n617 B.n616 585
R366 B.n617 B.n8 585
R367 B.n615 B.n7 585
R368 B.n952 B.n7 585
R369 B.n614 B.n6 585
R370 B.n953 B.n6 585
R371 B.n613 B.n5 585
R372 B.n954 B.n5 585
R373 B.n612 B.n611 585
R374 B.n611 B.n4 585
R375 B.n610 B.n142 585
R376 B.n610 B.n609 585
R377 B.n600 B.n143 585
R378 B.n144 B.n143 585
R379 B.n602 B.n601 585
R380 B.n603 B.n602 585
R381 B.n599 B.n148 585
R382 B.n152 B.n148 585
R383 B.n598 B.n597 585
R384 B.n597 B.n596 585
R385 B.n150 B.n149 585
R386 B.n151 B.n150 585
R387 B.n589 B.n588 585
R388 B.n590 B.n589 585
R389 B.n587 B.n157 585
R390 B.n157 B.n156 585
R391 B.n586 B.n585 585
R392 B.n585 B.n584 585
R393 B.n159 B.n158 585
R394 B.n160 B.n159 585
R395 B.n577 B.n576 585
R396 B.n578 B.n577 585
R397 B.n575 B.n165 585
R398 B.n165 B.n164 585
R399 B.n574 B.n573 585
R400 B.n573 B.n572 585
R401 B.n167 B.n166 585
R402 B.n168 B.n167 585
R403 B.n565 B.n564 585
R404 B.n566 B.n565 585
R405 B.n563 B.n173 585
R406 B.n173 B.n172 585
R407 B.n562 B.n561 585
R408 B.n561 B.n560 585
R409 B.n175 B.n174 585
R410 B.n553 B.n175 585
R411 B.n552 B.n551 585
R412 B.n554 B.n552 585
R413 B.n550 B.n180 585
R414 B.n180 B.n179 585
R415 B.n549 B.n548 585
R416 B.n548 B.n547 585
R417 B.n182 B.n181 585
R418 B.n183 B.n182 585
R419 B.n540 B.n539 585
R420 B.n541 B.n540 585
R421 B.n538 B.n188 585
R422 B.n188 B.n187 585
R423 B.n537 B.n536 585
R424 B.n536 B.n535 585
R425 B.n190 B.n189 585
R426 B.n191 B.n190 585
R427 B.n528 B.n527 585
R428 B.n529 B.n528 585
R429 B.n526 B.n196 585
R430 B.n196 B.n195 585
R431 B.n525 B.n524 585
R432 B.n524 B.n523 585
R433 B.n198 B.n197 585
R434 B.n199 B.n198 585
R435 B.n516 B.n515 585
R436 B.n517 B.n516 585
R437 B.n514 B.n203 585
R438 B.n207 B.n203 585
R439 B.n513 B.n512 585
R440 B.n512 B.n511 585
R441 B.n205 B.n204 585
R442 B.n206 B.n205 585
R443 B.n504 B.n503 585
R444 B.n505 B.n504 585
R445 B.n502 B.n212 585
R446 B.n212 B.n211 585
R447 B.n501 B.n500 585
R448 B.n500 B.n499 585
R449 B.n214 B.n213 585
R450 B.n215 B.n214 585
R451 B.n492 B.n491 585
R452 B.n493 B.n492 585
R453 B.n490 B.n220 585
R454 B.n220 B.n219 585
R455 B.n489 B.n488 585
R456 B.n488 B.n487 585
R457 B.n222 B.n221 585
R458 B.n223 B.n222 585
R459 B.n480 B.n479 585
R460 B.n481 B.n480 585
R461 B.n478 B.n228 585
R462 B.n228 B.n227 585
R463 B.n477 B.n476 585
R464 B.n476 B.n475 585
R465 B.n230 B.n229 585
R466 B.n231 B.n230 585
R467 B.n468 B.n467 585
R468 B.n469 B.n468 585
R469 B.n466 B.n236 585
R470 B.n236 B.n235 585
R471 B.n465 B.n464 585
R472 B.n464 B.n463 585
R473 B.n460 B.n240 585
R474 B.n459 B.n458 585
R475 B.n456 B.n241 585
R476 B.n456 B.n239 585
R477 B.n455 B.n454 585
R478 B.n453 B.n452 585
R479 B.n451 B.n243 585
R480 B.n449 B.n448 585
R481 B.n447 B.n244 585
R482 B.n446 B.n445 585
R483 B.n443 B.n245 585
R484 B.n441 B.n440 585
R485 B.n439 B.n246 585
R486 B.n438 B.n437 585
R487 B.n435 B.n247 585
R488 B.n433 B.n432 585
R489 B.n431 B.n248 585
R490 B.n430 B.n429 585
R491 B.n427 B.n249 585
R492 B.n425 B.n424 585
R493 B.n423 B.n250 585
R494 B.n422 B.n421 585
R495 B.n419 B.n251 585
R496 B.n417 B.n416 585
R497 B.n415 B.n252 585
R498 B.n414 B.n413 585
R499 B.n411 B.n253 585
R500 B.n409 B.n408 585
R501 B.n407 B.n254 585
R502 B.n406 B.n405 585
R503 B.n403 B.n255 585
R504 B.n401 B.n400 585
R505 B.n399 B.n256 585
R506 B.n398 B.n397 585
R507 B.n395 B.n257 585
R508 B.n393 B.n392 585
R509 B.n391 B.n258 585
R510 B.n390 B.n389 585
R511 B.n387 B.n259 585
R512 B.n385 B.n384 585
R513 B.n382 B.n260 585
R514 B.n381 B.n380 585
R515 B.n378 B.n263 585
R516 B.n376 B.n375 585
R517 B.n374 B.n264 585
R518 B.n373 B.n372 585
R519 B.n370 B.n265 585
R520 B.n368 B.n367 585
R521 B.n366 B.n266 585
R522 B.n364 B.n363 585
R523 B.n361 B.n269 585
R524 B.n359 B.n358 585
R525 B.n357 B.n270 585
R526 B.n356 B.n355 585
R527 B.n353 B.n271 585
R528 B.n351 B.n350 585
R529 B.n349 B.n272 585
R530 B.n348 B.n347 585
R531 B.n345 B.n273 585
R532 B.n343 B.n342 585
R533 B.n341 B.n274 585
R534 B.n340 B.n339 585
R535 B.n337 B.n275 585
R536 B.n335 B.n334 585
R537 B.n333 B.n276 585
R538 B.n332 B.n331 585
R539 B.n329 B.n277 585
R540 B.n327 B.n326 585
R541 B.n325 B.n278 585
R542 B.n324 B.n323 585
R543 B.n321 B.n279 585
R544 B.n319 B.n318 585
R545 B.n317 B.n280 585
R546 B.n316 B.n315 585
R547 B.n313 B.n281 585
R548 B.n311 B.n310 585
R549 B.n309 B.n282 585
R550 B.n308 B.n307 585
R551 B.n305 B.n283 585
R552 B.n303 B.n302 585
R553 B.n301 B.n284 585
R554 B.n300 B.n299 585
R555 B.n297 B.n285 585
R556 B.n295 B.n294 585
R557 B.n293 B.n286 585
R558 B.n292 B.n291 585
R559 B.n289 B.n287 585
R560 B.n238 B.n237 585
R561 B.n462 B.n461 585
R562 B.n463 B.n462 585
R563 B.n234 B.n233 585
R564 B.n235 B.n234 585
R565 B.n471 B.n470 585
R566 B.n470 B.n469 585
R567 B.n472 B.n232 585
R568 B.n232 B.n231 585
R569 B.n474 B.n473 585
R570 B.n475 B.n474 585
R571 B.n226 B.n225 585
R572 B.n227 B.n226 585
R573 B.n483 B.n482 585
R574 B.n482 B.n481 585
R575 B.n484 B.n224 585
R576 B.n224 B.n223 585
R577 B.n486 B.n485 585
R578 B.n487 B.n486 585
R579 B.n218 B.n217 585
R580 B.n219 B.n218 585
R581 B.n495 B.n494 585
R582 B.n494 B.n493 585
R583 B.n496 B.n216 585
R584 B.n216 B.n215 585
R585 B.n498 B.n497 585
R586 B.n499 B.n498 585
R587 B.n210 B.n209 585
R588 B.n211 B.n210 585
R589 B.n507 B.n506 585
R590 B.n506 B.n505 585
R591 B.n508 B.n208 585
R592 B.n208 B.n206 585
R593 B.n510 B.n509 585
R594 B.n511 B.n510 585
R595 B.n202 B.n201 585
R596 B.n207 B.n202 585
R597 B.n519 B.n518 585
R598 B.n518 B.n517 585
R599 B.n520 B.n200 585
R600 B.n200 B.n199 585
R601 B.n522 B.n521 585
R602 B.n523 B.n522 585
R603 B.n194 B.n193 585
R604 B.n195 B.n194 585
R605 B.n531 B.n530 585
R606 B.n530 B.n529 585
R607 B.n532 B.n192 585
R608 B.n192 B.n191 585
R609 B.n534 B.n533 585
R610 B.n535 B.n534 585
R611 B.n186 B.n185 585
R612 B.n187 B.n186 585
R613 B.n543 B.n542 585
R614 B.n542 B.n541 585
R615 B.n544 B.n184 585
R616 B.n184 B.n183 585
R617 B.n546 B.n545 585
R618 B.n547 B.n546 585
R619 B.n178 B.n177 585
R620 B.n179 B.n178 585
R621 B.n556 B.n555 585
R622 B.n555 B.n554 585
R623 B.n557 B.n176 585
R624 B.n553 B.n176 585
R625 B.n559 B.n558 585
R626 B.n560 B.n559 585
R627 B.n171 B.n170 585
R628 B.n172 B.n171 585
R629 B.n568 B.n567 585
R630 B.n567 B.n566 585
R631 B.n569 B.n169 585
R632 B.n169 B.n168 585
R633 B.n571 B.n570 585
R634 B.n572 B.n571 585
R635 B.n163 B.n162 585
R636 B.n164 B.n163 585
R637 B.n580 B.n579 585
R638 B.n579 B.n578 585
R639 B.n581 B.n161 585
R640 B.n161 B.n160 585
R641 B.n583 B.n582 585
R642 B.n584 B.n583 585
R643 B.n155 B.n154 585
R644 B.n156 B.n155 585
R645 B.n592 B.n591 585
R646 B.n591 B.n590 585
R647 B.n593 B.n153 585
R648 B.n153 B.n151 585
R649 B.n595 B.n594 585
R650 B.n596 B.n595 585
R651 B.n147 B.n146 585
R652 B.n152 B.n147 585
R653 B.n605 B.n604 585
R654 B.n604 B.n603 585
R655 B.n606 B.n145 585
R656 B.n145 B.n144 585
R657 B.n608 B.n607 585
R658 B.n609 B.n608 585
R659 B.n3 B.n0 585
R660 B.n4 B.n3 585
R661 B.n951 B.n1 585
R662 B.n952 B.n951 585
R663 B.n950 B.n949 585
R664 B.n950 B.n8 585
R665 B.n948 B.n9 585
R666 B.n12 B.n9 585
R667 B.n947 B.n946 585
R668 B.n946 B.n945 585
R669 B.n11 B.n10 585
R670 B.n944 B.n11 585
R671 B.n942 B.n941 585
R672 B.n943 B.n942 585
R673 B.n940 B.n17 585
R674 B.n17 B.n16 585
R675 B.n939 B.n938 585
R676 B.n938 B.n937 585
R677 B.n19 B.n18 585
R678 B.n936 B.n19 585
R679 B.n934 B.n933 585
R680 B.n935 B.n934 585
R681 B.n932 B.n24 585
R682 B.n24 B.n23 585
R683 B.n931 B.n930 585
R684 B.n930 B.n929 585
R685 B.n26 B.n25 585
R686 B.n928 B.n26 585
R687 B.n926 B.n925 585
R688 B.n927 B.n926 585
R689 B.n924 B.n31 585
R690 B.n31 B.n30 585
R691 B.n923 B.n922 585
R692 B.n922 B.n921 585
R693 B.n33 B.n32 585
R694 B.n920 B.n33 585
R695 B.n918 B.n917 585
R696 B.n919 B.n918 585
R697 B.n916 B.n37 585
R698 B.n40 B.n37 585
R699 B.n915 B.n914 585
R700 B.n914 B.n913 585
R701 B.n39 B.n38 585
R702 B.n912 B.n39 585
R703 B.n910 B.n909 585
R704 B.n911 B.n910 585
R705 B.n908 B.n45 585
R706 B.n45 B.n44 585
R707 B.n907 B.n906 585
R708 B.n906 B.n905 585
R709 B.n47 B.n46 585
R710 B.n904 B.n47 585
R711 B.n902 B.n901 585
R712 B.n903 B.n902 585
R713 B.n900 B.n52 585
R714 B.n52 B.n51 585
R715 B.n899 B.n898 585
R716 B.n898 B.n897 585
R717 B.n54 B.n53 585
R718 B.n896 B.n54 585
R719 B.n894 B.n893 585
R720 B.n895 B.n894 585
R721 B.n892 B.n59 585
R722 B.n59 B.n58 585
R723 B.n891 B.n890 585
R724 B.n890 B.n889 585
R725 B.n61 B.n60 585
R726 B.n888 B.n61 585
R727 B.n886 B.n885 585
R728 B.n887 B.n886 585
R729 B.n884 B.n66 585
R730 B.n66 B.n65 585
R731 B.n883 B.n882 585
R732 B.n882 B.n881 585
R733 B.n68 B.n67 585
R734 B.n880 B.n68 585
R735 B.n878 B.n877 585
R736 B.n879 B.n878 585
R737 B.n876 B.n73 585
R738 B.n73 B.n72 585
R739 B.n875 B.n874 585
R740 B.n874 B.n873 585
R741 B.n75 B.n74 585
R742 B.n872 B.n75 585
R743 B.n870 B.n869 585
R744 B.n871 B.n870 585
R745 B.n868 B.n80 585
R746 B.n80 B.n79 585
R747 B.n867 B.n866 585
R748 B.n866 B.n865 585
R749 B.n82 B.n81 585
R750 B.n864 B.n82 585
R751 B.n862 B.n861 585
R752 B.n863 B.n862 585
R753 B.n860 B.n87 585
R754 B.n87 B.n86 585
R755 B.n859 B.n858 585
R756 B.n858 B.n857 585
R757 B.n89 B.n88 585
R758 B.n856 B.n89 585
R759 B.n854 B.n853 585
R760 B.n855 B.n854 585
R761 B.n955 B.n954 585
R762 B.n953 B.n2 585
R763 B.n854 B.n94 454.062
R764 B.n679 B.n92 454.062
R765 B.n464 B.n238 454.062
R766 B.n462 B.n240 454.062
R767 B.n115 B.t17 334.33
R768 B.n122 B.t21 334.33
R769 B.n267 B.t10 334.33
R770 B.n261 B.t14 334.33
R771 B.n680 B.n93 256.663
R772 B.n686 B.n93 256.663
R773 B.n688 B.n93 256.663
R774 B.n694 B.n93 256.663
R775 B.n696 B.n93 256.663
R776 B.n702 B.n93 256.663
R777 B.n704 B.n93 256.663
R778 B.n710 B.n93 256.663
R779 B.n712 B.n93 256.663
R780 B.n718 B.n93 256.663
R781 B.n720 B.n93 256.663
R782 B.n726 B.n93 256.663
R783 B.n728 B.n93 256.663
R784 B.n734 B.n93 256.663
R785 B.n736 B.n93 256.663
R786 B.n742 B.n93 256.663
R787 B.n744 B.n93 256.663
R788 B.n750 B.n93 256.663
R789 B.n752 B.n93 256.663
R790 B.n759 B.n93 256.663
R791 B.n761 B.n93 256.663
R792 B.n767 B.n93 256.663
R793 B.n769 B.n93 256.663
R794 B.n775 B.n93 256.663
R795 B.n777 B.n93 256.663
R796 B.n783 B.n93 256.663
R797 B.n785 B.n93 256.663
R798 B.n791 B.n93 256.663
R799 B.n793 B.n93 256.663
R800 B.n799 B.n93 256.663
R801 B.n801 B.n93 256.663
R802 B.n807 B.n93 256.663
R803 B.n809 B.n93 256.663
R804 B.n815 B.n93 256.663
R805 B.n817 B.n93 256.663
R806 B.n823 B.n93 256.663
R807 B.n825 B.n93 256.663
R808 B.n831 B.n93 256.663
R809 B.n833 B.n93 256.663
R810 B.n839 B.n93 256.663
R811 B.n841 B.n93 256.663
R812 B.n847 B.n93 256.663
R813 B.n849 B.n93 256.663
R814 B.n457 B.n239 256.663
R815 B.n242 B.n239 256.663
R816 B.n450 B.n239 256.663
R817 B.n444 B.n239 256.663
R818 B.n442 B.n239 256.663
R819 B.n436 B.n239 256.663
R820 B.n434 B.n239 256.663
R821 B.n428 B.n239 256.663
R822 B.n426 B.n239 256.663
R823 B.n420 B.n239 256.663
R824 B.n418 B.n239 256.663
R825 B.n412 B.n239 256.663
R826 B.n410 B.n239 256.663
R827 B.n404 B.n239 256.663
R828 B.n402 B.n239 256.663
R829 B.n396 B.n239 256.663
R830 B.n394 B.n239 256.663
R831 B.n388 B.n239 256.663
R832 B.n386 B.n239 256.663
R833 B.n379 B.n239 256.663
R834 B.n377 B.n239 256.663
R835 B.n371 B.n239 256.663
R836 B.n369 B.n239 256.663
R837 B.n362 B.n239 256.663
R838 B.n360 B.n239 256.663
R839 B.n354 B.n239 256.663
R840 B.n352 B.n239 256.663
R841 B.n346 B.n239 256.663
R842 B.n344 B.n239 256.663
R843 B.n338 B.n239 256.663
R844 B.n336 B.n239 256.663
R845 B.n330 B.n239 256.663
R846 B.n328 B.n239 256.663
R847 B.n322 B.n239 256.663
R848 B.n320 B.n239 256.663
R849 B.n314 B.n239 256.663
R850 B.n312 B.n239 256.663
R851 B.n306 B.n239 256.663
R852 B.n304 B.n239 256.663
R853 B.n298 B.n239 256.663
R854 B.n296 B.n239 256.663
R855 B.n290 B.n239 256.663
R856 B.n288 B.n239 256.663
R857 B.n957 B.n956 256.663
R858 B.n850 B.n848 163.367
R859 B.n846 B.n96 163.367
R860 B.n842 B.n840 163.367
R861 B.n838 B.n98 163.367
R862 B.n834 B.n832 163.367
R863 B.n830 B.n100 163.367
R864 B.n826 B.n824 163.367
R865 B.n822 B.n102 163.367
R866 B.n818 B.n816 163.367
R867 B.n814 B.n104 163.367
R868 B.n810 B.n808 163.367
R869 B.n806 B.n106 163.367
R870 B.n802 B.n800 163.367
R871 B.n798 B.n108 163.367
R872 B.n794 B.n792 163.367
R873 B.n790 B.n110 163.367
R874 B.n786 B.n784 163.367
R875 B.n782 B.n112 163.367
R876 B.n778 B.n776 163.367
R877 B.n774 B.n114 163.367
R878 B.n770 B.n768 163.367
R879 B.n766 B.n119 163.367
R880 B.n762 B.n760 163.367
R881 B.n758 B.n121 163.367
R882 B.n753 B.n751 163.367
R883 B.n749 B.n125 163.367
R884 B.n745 B.n743 163.367
R885 B.n741 B.n127 163.367
R886 B.n737 B.n735 163.367
R887 B.n733 B.n129 163.367
R888 B.n729 B.n727 163.367
R889 B.n725 B.n131 163.367
R890 B.n721 B.n719 163.367
R891 B.n717 B.n133 163.367
R892 B.n713 B.n711 163.367
R893 B.n709 B.n135 163.367
R894 B.n705 B.n703 163.367
R895 B.n701 B.n137 163.367
R896 B.n697 B.n695 163.367
R897 B.n693 B.n139 163.367
R898 B.n689 B.n687 163.367
R899 B.n685 B.n141 163.367
R900 B.n681 B.n679 163.367
R901 B.n464 B.n236 163.367
R902 B.n468 B.n236 163.367
R903 B.n468 B.n230 163.367
R904 B.n476 B.n230 163.367
R905 B.n476 B.n228 163.367
R906 B.n480 B.n228 163.367
R907 B.n480 B.n222 163.367
R908 B.n488 B.n222 163.367
R909 B.n488 B.n220 163.367
R910 B.n492 B.n220 163.367
R911 B.n492 B.n214 163.367
R912 B.n500 B.n214 163.367
R913 B.n500 B.n212 163.367
R914 B.n504 B.n212 163.367
R915 B.n504 B.n205 163.367
R916 B.n512 B.n205 163.367
R917 B.n512 B.n203 163.367
R918 B.n516 B.n203 163.367
R919 B.n516 B.n198 163.367
R920 B.n524 B.n198 163.367
R921 B.n524 B.n196 163.367
R922 B.n528 B.n196 163.367
R923 B.n528 B.n190 163.367
R924 B.n536 B.n190 163.367
R925 B.n536 B.n188 163.367
R926 B.n540 B.n188 163.367
R927 B.n540 B.n182 163.367
R928 B.n548 B.n182 163.367
R929 B.n548 B.n180 163.367
R930 B.n552 B.n180 163.367
R931 B.n552 B.n175 163.367
R932 B.n561 B.n175 163.367
R933 B.n561 B.n173 163.367
R934 B.n565 B.n173 163.367
R935 B.n565 B.n167 163.367
R936 B.n573 B.n167 163.367
R937 B.n573 B.n165 163.367
R938 B.n577 B.n165 163.367
R939 B.n577 B.n159 163.367
R940 B.n585 B.n159 163.367
R941 B.n585 B.n157 163.367
R942 B.n589 B.n157 163.367
R943 B.n589 B.n150 163.367
R944 B.n597 B.n150 163.367
R945 B.n597 B.n148 163.367
R946 B.n602 B.n148 163.367
R947 B.n602 B.n143 163.367
R948 B.n610 B.n143 163.367
R949 B.n611 B.n610 163.367
R950 B.n611 B.n5 163.367
R951 B.n6 B.n5 163.367
R952 B.n7 B.n6 163.367
R953 B.n617 B.n7 163.367
R954 B.n618 B.n617 163.367
R955 B.n618 B.n13 163.367
R956 B.n14 B.n13 163.367
R957 B.n15 B.n14 163.367
R958 B.n623 B.n15 163.367
R959 B.n623 B.n20 163.367
R960 B.n21 B.n20 163.367
R961 B.n22 B.n21 163.367
R962 B.n628 B.n22 163.367
R963 B.n628 B.n27 163.367
R964 B.n28 B.n27 163.367
R965 B.n29 B.n28 163.367
R966 B.n633 B.n29 163.367
R967 B.n633 B.n34 163.367
R968 B.n35 B.n34 163.367
R969 B.n36 B.n35 163.367
R970 B.n638 B.n36 163.367
R971 B.n638 B.n41 163.367
R972 B.n42 B.n41 163.367
R973 B.n43 B.n42 163.367
R974 B.n643 B.n43 163.367
R975 B.n643 B.n48 163.367
R976 B.n49 B.n48 163.367
R977 B.n50 B.n49 163.367
R978 B.n648 B.n50 163.367
R979 B.n648 B.n55 163.367
R980 B.n56 B.n55 163.367
R981 B.n57 B.n56 163.367
R982 B.n653 B.n57 163.367
R983 B.n653 B.n62 163.367
R984 B.n63 B.n62 163.367
R985 B.n64 B.n63 163.367
R986 B.n658 B.n64 163.367
R987 B.n658 B.n69 163.367
R988 B.n70 B.n69 163.367
R989 B.n71 B.n70 163.367
R990 B.n663 B.n71 163.367
R991 B.n663 B.n76 163.367
R992 B.n77 B.n76 163.367
R993 B.n78 B.n77 163.367
R994 B.n668 B.n78 163.367
R995 B.n668 B.n83 163.367
R996 B.n84 B.n83 163.367
R997 B.n85 B.n84 163.367
R998 B.n673 B.n85 163.367
R999 B.n673 B.n90 163.367
R1000 B.n91 B.n90 163.367
R1001 B.n92 B.n91 163.367
R1002 B.n458 B.n456 163.367
R1003 B.n456 B.n455 163.367
R1004 B.n452 B.n451 163.367
R1005 B.n449 B.n244 163.367
R1006 B.n445 B.n443 163.367
R1007 B.n441 B.n246 163.367
R1008 B.n437 B.n435 163.367
R1009 B.n433 B.n248 163.367
R1010 B.n429 B.n427 163.367
R1011 B.n425 B.n250 163.367
R1012 B.n421 B.n419 163.367
R1013 B.n417 B.n252 163.367
R1014 B.n413 B.n411 163.367
R1015 B.n409 B.n254 163.367
R1016 B.n405 B.n403 163.367
R1017 B.n401 B.n256 163.367
R1018 B.n397 B.n395 163.367
R1019 B.n393 B.n258 163.367
R1020 B.n389 B.n387 163.367
R1021 B.n385 B.n260 163.367
R1022 B.n380 B.n378 163.367
R1023 B.n376 B.n264 163.367
R1024 B.n372 B.n370 163.367
R1025 B.n368 B.n266 163.367
R1026 B.n363 B.n361 163.367
R1027 B.n359 B.n270 163.367
R1028 B.n355 B.n353 163.367
R1029 B.n351 B.n272 163.367
R1030 B.n347 B.n345 163.367
R1031 B.n343 B.n274 163.367
R1032 B.n339 B.n337 163.367
R1033 B.n335 B.n276 163.367
R1034 B.n331 B.n329 163.367
R1035 B.n327 B.n278 163.367
R1036 B.n323 B.n321 163.367
R1037 B.n319 B.n280 163.367
R1038 B.n315 B.n313 163.367
R1039 B.n311 B.n282 163.367
R1040 B.n307 B.n305 163.367
R1041 B.n303 B.n284 163.367
R1042 B.n299 B.n297 163.367
R1043 B.n295 B.n286 163.367
R1044 B.n291 B.n289 163.367
R1045 B.n462 B.n234 163.367
R1046 B.n470 B.n234 163.367
R1047 B.n470 B.n232 163.367
R1048 B.n474 B.n232 163.367
R1049 B.n474 B.n226 163.367
R1050 B.n482 B.n226 163.367
R1051 B.n482 B.n224 163.367
R1052 B.n486 B.n224 163.367
R1053 B.n486 B.n218 163.367
R1054 B.n494 B.n218 163.367
R1055 B.n494 B.n216 163.367
R1056 B.n498 B.n216 163.367
R1057 B.n498 B.n210 163.367
R1058 B.n506 B.n210 163.367
R1059 B.n506 B.n208 163.367
R1060 B.n510 B.n208 163.367
R1061 B.n510 B.n202 163.367
R1062 B.n518 B.n202 163.367
R1063 B.n518 B.n200 163.367
R1064 B.n522 B.n200 163.367
R1065 B.n522 B.n194 163.367
R1066 B.n530 B.n194 163.367
R1067 B.n530 B.n192 163.367
R1068 B.n534 B.n192 163.367
R1069 B.n534 B.n186 163.367
R1070 B.n542 B.n186 163.367
R1071 B.n542 B.n184 163.367
R1072 B.n546 B.n184 163.367
R1073 B.n546 B.n178 163.367
R1074 B.n555 B.n178 163.367
R1075 B.n555 B.n176 163.367
R1076 B.n559 B.n176 163.367
R1077 B.n559 B.n171 163.367
R1078 B.n567 B.n171 163.367
R1079 B.n567 B.n169 163.367
R1080 B.n571 B.n169 163.367
R1081 B.n571 B.n163 163.367
R1082 B.n579 B.n163 163.367
R1083 B.n579 B.n161 163.367
R1084 B.n583 B.n161 163.367
R1085 B.n583 B.n155 163.367
R1086 B.n591 B.n155 163.367
R1087 B.n591 B.n153 163.367
R1088 B.n595 B.n153 163.367
R1089 B.n595 B.n147 163.367
R1090 B.n604 B.n147 163.367
R1091 B.n604 B.n145 163.367
R1092 B.n608 B.n145 163.367
R1093 B.n608 B.n3 163.367
R1094 B.n955 B.n3 163.367
R1095 B.n951 B.n2 163.367
R1096 B.n951 B.n950 163.367
R1097 B.n950 B.n9 163.367
R1098 B.n946 B.n9 163.367
R1099 B.n946 B.n11 163.367
R1100 B.n942 B.n11 163.367
R1101 B.n942 B.n17 163.367
R1102 B.n938 B.n17 163.367
R1103 B.n938 B.n19 163.367
R1104 B.n934 B.n19 163.367
R1105 B.n934 B.n24 163.367
R1106 B.n930 B.n24 163.367
R1107 B.n930 B.n26 163.367
R1108 B.n926 B.n26 163.367
R1109 B.n926 B.n31 163.367
R1110 B.n922 B.n31 163.367
R1111 B.n922 B.n33 163.367
R1112 B.n918 B.n33 163.367
R1113 B.n918 B.n37 163.367
R1114 B.n914 B.n37 163.367
R1115 B.n914 B.n39 163.367
R1116 B.n910 B.n39 163.367
R1117 B.n910 B.n45 163.367
R1118 B.n906 B.n45 163.367
R1119 B.n906 B.n47 163.367
R1120 B.n902 B.n47 163.367
R1121 B.n902 B.n52 163.367
R1122 B.n898 B.n52 163.367
R1123 B.n898 B.n54 163.367
R1124 B.n894 B.n54 163.367
R1125 B.n894 B.n59 163.367
R1126 B.n890 B.n59 163.367
R1127 B.n890 B.n61 163.367
R1128 B.n886 B.n61 163.367
R1129 B.n886 B.n66 163.367
R1130 B.n882 B.n66 163.367
R1131 B.n882 B.n68 163.367
R1132 B.n878 B.n68 163.367
R1133 B.n878 B.n73 163.367
R1134 B.n874 B.n73 163.367
R1135 B.n874 B.n75 163.367
R1136 B.n870 B.n75 163.367
R1137 B.n870 B.n80 163.367
R1138 B.n866 B.n80 163.367
R1139 B.n866 B.n82 163.367
R1140 B.n862 B.n82 163.367
R1141 B.n862 B.n87 163.367
R1142 B.n858 B.n87 163.367
R1143 B.n858 B.n89 163.367
R1144 B.n854 B.n89 163.367
R1145 B.n122 B.t22 115.466
R1146 B.n267 B.t13 115.466
R1147 B.n115 B.t19 115.451
R1148 B.n261 B.t16 115.451
R1149 B.n463 B.n239 82.1356
R1150 B.n855 B.n93 82.1356
R1151 B.n849 B.n94 71.676
R1152 B.n848 B.n847 71.676
R1153 B.n841 B.n96 71.676
R1154 B.n840 B.n839 71.676
R1155 B.n833 B.n98 71.676
R1156 B.n832 B.n831 71.676
R1157 B.n825 B.n100 71.676
R1158 B.n824 B.n823 71.676
R1159 B.n817 B.n102 71.676
R1160 B.n816 B.n815 71.676
R1161 B.n809 B.n104 71.676
R1162 B.n808 B.n807 71.676
R1163 B.n801 B.n106 71.676
R1164 B.n800 B.n799 71.676
R1165 B.n793 B.n108 71.676
R1166 B.n792 B.n791 71.676
R1167 B.n785 B.n110 71.676
R1168 B.n784 B.n783 71.676
R1169 B.n777 B.n112 71.676
R1170 B.n776 B.n775 71.676
R1171 B.n769 B.n114 71.676
R1172 B.n768 B.n767 71.676
R1173 B.n761 B.n119 71.676
R1174 B.n760 B.n759 71.676
R1175 B.n752 B.n121 71.676
R1176 B.n751 B.n750 71.676
R1177 B.n744 B.n125 71.676
R1178 B.n743 B.n742 71.676
R1179 B.n736 B.n127 71.676
R1180 B.n735 B.n734 71.676
R1181 B.n728 B.n129 71.676
R1182 B.n727 B.n726 71.676
R1183 B.n720 B.n131 71.676
R1184 B.n719 B.n718 71.676
R1185 B.n712 B.n133 71.676
R1186 B.n711 B.n710 71.676
R1187 B.n704 B.n135 71.676
R1188 B.n703 B.n702 71.676
R1189 B.n696 B.n137 71.676
R1190 B.n695 B.n694 71.676
R1191 B.n688 B.n139 71.676
R1192 B.n687 B.n686 71.676
R1193 B.n680 B.n141 71.676
R1194 B.n681 B.n680 71.676
R1195 B.n686 B.n685 71.676
R1196 B.n689 B.n688 71.676
R1197 B.n694 B.n693 71.676
R1198 B.n697 B.n696 71.676
R1199 B.n702 B.n701 71.676
R1200 B.n705 B.n704 71.676
R1201 B.n710 B.n709 71.676
R1202 B.n713 B.n712 71.676
R1203 B.n718 B.n717 71.676
R1204 B.n721 B.n720 71.676
R1205 B.n726 B.n725 71.676
R1206 B.n729 B.n728 71.676
R1207 B.n734 B.n733 71.676
R1208 B.n737 B.n736 71.676
R1209 B.n742 B.n741 71.676
R1210 B.n745 B.n744 71.676
R1211 B.n750 B.n749 71.676
R1212 B.n753 B.n752 71.676
R1213 B.n759 B.n758 71.676
R1214 B.n762 B.n761 71.676
R1215 B.n767 B.n766 71.676
R1216 B.n770 B.n769 71.676
R1217 B.n775 B.n774 71.676
R1218 B.n778 B.n777 71.676
R1219 B.n783 B.n782 71.676
R1220 B.n786 B.n785 71.676
R1221 B.n791 B.n790 71.676
R1222 B.n794 B.n793 71.676
R1223 B.n799 B.n798 71.676
R1224 B.n802 B.n801 71.676
R1225 B.n807 B.n806 71.676
R1226 B.n810 B.n809 71.676
R1227 B.n815 B.n814 71.676
R1228 B.n818 B.n817 71.676
R1229 B.n823 B.n822 71.676
R1230 B.n826 B.n825 71.676
R1231 B.n831 B.n830 71.676
R1232 B.n834 B.n833 71.676
R1233 B.n839 B.n838 71.676
R1234 B.n842 B.n841 71.676
R1235 B.n847 B.n846 71.676
R1236 B.n850 B.n849 71.676
R1237 B.n457 B.n240 71.676
R1238 B.n455 B.n242 71.676
R1239 B.n451 B.n450 71.676
R1240 B.n444 B.n244 71.676
R1241 B.n443 B.n442 71.676
R1242 B.n436 B.n246 71.676
R1243 B.n435 B.n434 71.676
R1244 B.n428 B.n248 71.676
R1245 B.n427 B.n426 71.676
R1246 B.n420 B.n250 71.676
R1247 B.n419 B.n418 71.676
R1248 B.n412 B.n252 71.676
R1249 B.n411 B.n410 71.676
R1250 B.n404 B.n254 71.676
R1251 B.n403 B.n402 71.676
R1252 B.n396 B.n256 71.676
R1253 B.n395 B.n394 71.676
R1254 B.n388 B.n258 71.676
R1255 B.n387 B.n386 71.676
R1256 B.n379 B.n260 71.676
R1257 B.n378 B.n377 71.676
R1258 B.n371 B.n264 71.676
R1259 B.n370 B.n369 71.676
R1260 B.n362 B.n266 71.676
R1261 B.n361 B.n360 71.676
R1262 B.n354 B.n270 71.676
R1263 B.n353 B.n352 71.676
R1264 B.n346 B.n272 71.676
R1265 B.n345 B.n344 71.676
R1266 B.n338 B.n274 71.676
R1267 B.n337 B.n336 71.676
R1268 B.n330 B.n276 71.676
R1269 B.n329 B.n328 71.676
R1270 B.n322 B.n278 71.676
R1271 B.n321 B.n320 71.676
R1272 B.n314 B.n280 71.676
R1273 B.n313 B.n312 71.676
R1274 B.n306 B.n282 71.676
R1275 B.n305 B.n304 71.676
R1276 B.n298 B.n284 71.676
R1277 B.n297 B.n296 71.676
R1278 B.n290 B.n286 71.676
R1279 B.n289 B.n288 71.676
R1280 B.n458 B.n457 71.676
R1281 B.n452 B.n242 71.676
R1282 B.n450 B.n449 71.676
R1283 B.n445 B.n444 71.676
R1284 B.n442 B.n441 71.676
R1285 B.n437 B.n436 71.676
R1286 B.n434 B.n433 71.676
R1287 B.n429 B.n428 71.676
R1288 B.n426 B.n425 71.676
R1289 B.n421 B.n420 71.676
R1290 B.n418 B.n417 71.676
R1291 B.n413 B.n412 71.676
R1292 B.n410 B.n409 71.676
R1293 B.n405 B.n404 71.676
R1294 B.n402 B.n401 71.676
R1295 B.n397 B.n396 71.676
R1296 B.n394 B.n393 71.676
R1297 B.n389 B.n388 71.676
R1298 B.n386 B.n385 71.676
R1299 B.n380 B.n379 71.676
R1300 B.n377 B.n376 71.676
R1301 B.n372 B.n371 71.676
R1302 B.n369 B.n368 71.676
R1303 B.n363 B.n362 71.676
R1304 B.n360 B.n359 71.676
R1305 B.n355 B.n354 71.676
R1306 B.n352 B.n351 71.676
R1307 B.n347 B.n346 71.676
R1308 B.n344 B.n343 71.676
R1309 B.n339 B.n338 71.676
R1310 B.n336 B.n335 71.676
R1311 B.n331 B.n330 71.676
R1312 B.n328 B.n327 71.676
R1313 B.n323 B.n322 71.676
R1314 B.n320 B.n319 71.676
R1315 B.n315 B.n314 71.676
R1316 B.n312 B.n311 71.676
R1317 B.n307 B.n306 71.676
R1318 B.n304 B.n303 71.676
R1319 B.n299 B.n298 71.676
R1320 B.n296 B.n295 71.676
R1321 B.n291 B.n290 71.676
R1322 B.n288 B.n238 71.676
R1323 B.n956 B.n955 71.676
R1324 B.n956 B.n2 71.676
R1325 B.n123 B.t23 68.9196
R1326 B.n268 B.t12 68.9196
R1327 B.n116 B.t20 68.9059
R1328 B.n262 B.t15 68.9059
R1329 B.n117 B.n116 59.5399
R1330 B.n756 B.n123 59.5399
R1331 B.n365 B.n268 59.5399
R1332 B.n383 B.n262 59.5399
R1333 B.n116 B.n115 46.546
R1334 B.n123 B.n122 46.546
R1335 B.n268 B.n267 46.546
R1336 B.n262 B.n261 46.546
R1337 B.n463 B.n235 46.1591
R1338 B.n469 B.n235 46.1591
R1339 B.n469 B.n231 46.1591
R1340 B.n475 B.n231 46.1591
R1341 B.n475 B.n227 46.1591
R1342 B.n481 B.n227 46.1591
R1343 B.n487 B.n223 46.1591
R1344 B.n487 B.n219 46.1591
R1345 B.n493 B.n219 46.1591
R1346 B.n493 B.n215 46.1591
R1347 B.n499 B.n215 46.1591
R1348 B.n499 B.n211 46.1591
R1349 B.n505 B.n211 46.1591
R1350 B.n505 B.n206 46.1591
R1351 B.n511 B.n206 46.1591
R1352 B.n511 B.n207 46.1591
R1353 B.n517 B.n199 46.1591
R1354 B.n523 B.n199 46.1591
R1355 B.n523 B.n195 46.1591
R1356 B.n529 B.n195 46.1591
R1357 B.n529 B.n191 46.1591
R1358 B.n535 B.n191 46.1591
R1359 B.n541 B.n187 46.1591
R1360 B.n541 B.n183 46.1591
R1361 B.n547 B.n183 46.1591
R1362 B.n547 B.n179 46.1591
R1363 B.n554 B.n179 46.1591
R1364 B.n554 B.n553 46.1591
R1365 B.n560 B.n172 46.1591
R1366 B.n566 B.n172 46.1591
R1367 B.n566 B.n168 46.1591
R1368 B.n572 B.n168 46.1591
R1369 B.n572 B.n164 46.1591
R1370 B.n578 B.n164 46.1591
R1371 B.n584 B.n160 46.1591
R1372 B.n584 B.n156 46.1591
R1373 B.n590 B.n156 46.1591
R1374 B.n590 B.n151 46.1591
R1375 B.n596 B.n151 46.1591
R1376 B.n596 B.n152 46.1591
R1377 B.n603 B.n144 46.1591
R1378 B.n609 B.n144 46.1591
R1379 B.n609 B.n4 46.1591
R1380 B.n954 B.n4 46.1591
R1381 B.n954 B.n953 46.1591
R1382 B.n953 B.n952 46.1591
R1383 B.n952 B.n8 46.1591
R1384 B.n12 B.n8 46.1591
R1385 B.n945 B.n12 46.1591
R1386 B.n944 B.n943 46.1591
R1387 B.n943 B.n16 46.1591
R1388 B.n937 B.n16 46.1591
R1389 B.n937 B.n936 46.1591
R1390 B.n936 B.n935 46.1591
R1391 B.n935 B.n23 46.1591
R1392 B.n929 B.n928 46.1591
R1393 B.n928 B.n927 46.1591
R1394 B.n927 B.n30 46.1591
R1395 B.n921 B.n30 46.1591
R1396 B.n921 B.n920 46.1591
R1397 B.n920 B.n919 46.1591
R1398 B.n913 B.n40 46.1591
R1399 B.n913 B.n912 46.1591
R1400 B.n912 B.n911 46.1591
R1401 B.n911 B.n44 46.1591
R1402 B.n905 B.n44 46.1591
R1403 B.n905 B.n904 46.1591
R1404 B.n903 B.n51 46.1591
R1405 B.n897 B.n51 46.1591
R1406 B.n897 B.n896 46.1591
R1407 B.n896 B.n895 46.1591
R1408 B.n895 B.n58 46.1591
R1409 B.n889 B.n58 46.1591
R1410 B.n888 B.n887 46.1591
R1411 B.n887 B.n65 46.1591
R1412 B.n881 B.n65 46.1591
R1413 B.n881 B.n880 46.1591
R1414 B.n880 B.n879 46.1591
R1415 B.n879 B.n72 46.1591
R1416 B.n873 B.n72 46.1591
R1417 B.n873 B.n872 46.1591
R1418 B.n872 B.n871 46.1591
R1419 B.n871 B.n79 46.1591
R1420 B.n865 B.n864 46.1591
R1421 B.n864 B.n863 46.1591
R1422 B.n863 B.n86 46.1591
R1423 B.n857 B.n86 46.1591
R1424 B.n857 B.n856 46.1591
R1425 B.n856 B.n855 46.1591
R1426 B.n481 B.t11 40.0499
R1427 B.n517 B.t3 40.0499
R1428 B.n889 B.t7 40.0499
R1429 B.n865 B.t18 40.0499
R1430 B.t2 B.n187 37.3347
R1431 B.n904 B.t0 37.3347
R1432 B.n560 B.t6 34.6194
R1433 B.n919 B.t9 34.6194
R1434 B.t8 B.n160 31.9042
R1435 B.t5 B.n23 31.9042
R1436 B.n678 B.n677 29.5029
R1437 B.n461 B.n460 29.5029
R1438 B.n465 B.n237 29.5029
R1439 B.n853 B.n852 29.5029
R1440 B.n603 B.t1 29.189
R1441 B.n945 B.t4 29.189
R1442 B B.n957 18.0485
R1443 B.n152 B.t1 16.9706
R1444 B.t4 B.n944 16.9706
R1445 B.n578 B.t8 14.2554
R1446 B.n929 B.t5 14.2554
R1447 B.n553 B.t6 11.5401
R1448 B.n40 B.t9 11.5401
R1449 B.n461 B.n233 10.6151
R1450 B.n471 B.n233 10.6151
R1451 B.n472 B.n471 10.6151
R1452 B.n473 B.n472 10.6151
R1453 B.n473 B.n225 10.6151
R1454 B.n483 B.n225 10.6151
R1455 B.n484 B.n483 10.6151
R1456 B.n485 B.n484 10.6151
R1457 B.n485 B.n217 10.6151
R1458 B.n495 B.n217 10.6151
R1459 B.n496 B.n495 10.6151
R1460 B.n497 B.n496 10.6151
R1461 B.n497 B.n209 10.6151
R1462 B.n507 B.n209 10.6151
R1463 B.n508 B.n507 10.6151
R1464 B.n509 B.n508 10.6151
R1465 B.n509 B.n201 10.6151
R1466 B.n519 B.n201 10.6151
R1467 B.n520 B.n519 10.6151
R1468 B.n521 B.n520 10.6151
R1469 B.n521 B.n193 10.6151
R1470 B.n531 B.n193 10.6151
R1471 B.n532 B.n531 10.6151
R1472 B.n533 B.n532 10.6151
R1473 B.n533 B.n185 10.6151
R1474 B.n543 B.n185 10.6151
R1475 B.n544 B.n543 10.6151
R1476 B.n545 B.n544 10.6151
R1477 B.n545 B.n177 10.6151
R1478 B.n556 B.n177 10.6151
R1479 B.n557 B.n556 10.6151
R1480 B.n558 B.n557 10.6151
R1481 B.n558 B.n170 10.6151
R1482 B.n568 B.n170 10.6151
R1483 B.n569 B.n568 10.6151
R1484 B.n570 B.n569 10.6151
R1485 B.n570 B.n162 10.6151
R1486 B.n580 B.n162 10.6151
R1487 B.n581 B.n580 10.6151
R1488 B.n582 B.n581 10.6151
R1489 B.n582 B.n154 10.6151
R1490 B.n592 B.n154 10.6151
R1491 B.n593 B.n592 10.6151
R1492 B.n594 B.n593 10.6151
R1493 B.n594 B.n146 10.6151
R1494 B.n605 B.n146 10.6151
R1495 B.n606 B.n605 10.6151
R1496 B.n607 B.n606 10.6151
R1497 B.n607 B.n0 10.6151
R1498 B.n460 B.n459 10.6151
R1499 B.n459 B.n241 10.6151
R1500 B.n454 B.n241 10.6151
R1501 B.n454 B.n453 10.6151
R1502 B.n453 B.n243 10.6151
R1503 B.n448 B.n243 10.6151
R1504 B.n448 B.n447 10.6151
R1505 B.n447 B.n446 10.6151
R1506 B.n446 B.n245 10.6151
R1507 B.n440 B.n245 10.6151
R1508 B.n440 B.n439 10.6151
R1509 B.n439 B.n438 10.6151
R1510 B.n438 B.n247 10.6151
R1511 B.n432 B.n247 10.6151
R1512 B.n432 B.n431 10.6151
R1513 B.n431 B.n430 10.6151
R1514 B.n430 B.n249 10.6151
R1515 B.n424 B.n249 10.6151
R1516 B.n424 B.n423 10.6151
R1517 B.n423 B.n422 10.6151
R1518 B.n422 B.n251 10.6151
R1519 B.n416 B.n251 10.6151
R1520 B.n416 B.n415 10.6151
R1521 B.n415 B.n414 10.6151
R1522 B.n414 B.n253 10.6151
R1523 B.n408 B.n253 10.6151
R1524 B.n408 B.n407 10.6151
R1525 B.n407 B.n406 10.6151
R1526 B.n406 B.n255 10.6151
R1527 B.n400 B.n255 10.6151
R1528 B.n400 B.n399 10.6151
R1529 B.n399 B.n398 10.6151
R1530 B.n398 B.n257 10.6151
R1531 B.n392 B.n257 10.6151
R1532 B.n392 B.n391 10.6151
R1533 B.n391 B.n390 10.6151
R1534 B.n390 B.n259 10.6151
R1535 B.n384 B.n259 10.6151
R1536 B.n382 B.n381 10.6151
R1537 B.n381 B.n263 10.6151
R1538 B.n375 B.n263 10.6151
R1539 B.n375 B.n374 10.6151
R1540 B.n374 B.n373 10.6151
R1541 B.n373 B.n265 10.6151
R1542 B.n367 B.n265 10.6151
R1543 B.n367 B.n366 10.6151
R1544 B.n364 B.n269 10.6151
R1545 B.n358 B.n269 10.6151
R1546 B.n358 B.n357 10.6151
R1547 B.n357 B.n356 10.6151
R1548 B.n356 B.n271 10.6151
R1549 B.n350 B.n271 10.6151
R1550 B.n350 B.n349 10.6151
R1551 B.n349 B.n348 10.6151
R1552 B.n348 B.n273 10.6151
R1553 B.n342 B.n273 10.6151
R1554 B.n342 B.n341 10.6151
R1555 B.n341 B.n340 10.6151
R1556 B.n340 B.n275 10.6151
R1557 B.n334 B.n275 10.6151
R1558 B.n334 B.n333 10.6151
R1559 B.n333 B.n332 10.6151
R1560 B.n332 B.n277 10.6151
R1561 B.n326 B.n277 10.6151
R1562 B.n326 B.n325 10.6151
R1563 B.n325 B.n324 10.6151
R1564 B.n324 B.n279 10.6151
R1565 B.n318 B.n279 10.6151
R1566 B.n318 B.n317 10.6151
R1567 B.n317 B.n316 10.6151
R1568 B.n316 B.n281 10.6151
R1569 B.n310 B.n281 10.6151
R1570 B.n310 B.n309 10.6151
R1571 B.n309 B.n308 10.6151
R1572 B.n308 B.n283 10.6151
R1573 B.n302 B.n283 10.6151
R1574 B.n302 B.n301 10.6151
R1575 B.n301 B.n300 10.6151
R1576 B.n300 B.n285 10.6151
R1577 B.n294 B.n285 10.6151
R1578 B.n294 B.n293 10.6151
R1579 B.n293 B.n292 10.6151
R1580 B.n292 B.n287 10.6151
R1581 B.n287 B.n237 10.6151
R1582 B.n466 B.n465 10.6151
R1583 B.n467 B.n466 10.6151
R1584 B.n467 B.n229 10.6151
R1585 B.n477 B.n229 10.6151
R1586 B.n478 B.n477 10.6151
R1587 B.n479 B.n478 10.6151
R1588 B.n479 B.n221 10.6151
R1589 B.n489 B.n221 10.6151
R1590 B.n490 B.n489 10.6151
R1591 B.n491 B.n490 10.6151
R1592 B.n491 B.n213 10.6151
R1593 B.n501 B.n213 10.6151
R1594 B.n502 B.n501 10.6151
R1595 B.n503 B.n502 10.6151
R1596 B.n503 B.n204 10.6151
R1597 B.n513 B.n204 10.6151
R1598 B.n514 B.n513 10.6151
R1599 B.n515 B.n514 10.6151
R1600 B.n515 B.n197 10.6151
R1601 B.n525 B.n197 10.6151
R1602 B.n526 B.n525 10.6151
R1603 B.n527 B.n526 10.6151
R1604 B.n527 B.n189 10.6151
R1605 B.n537 B.n189 10.6151
R1606 B.n538 B.n537 10.6151
R1607 B.n539 B.n538 10.6151
R1608 B.n539 B.n181 10.6151
R1609 B.n549 B.n181 10.6151
R1610 B.n550 B.n549 10.6151
R1611 B.n551 B.n550 10.6151
R1612 B.n551 B.n174 10.6151
R1613 B.n562 B.n174 10.6151
R1614 B.n563 B.n562 10.6151
R1615 B.n564 B.n563 10.6151
R1616 B.n564 B.n166 10.6151
R1617 B.n574 B.n166 10.6151
R1618 B.n575 B.n574 10.6151
R1619 B.n576 B.n575 10.6151
R1620 B.n576 B.n158 10.6151
R1621 B.n586 B.n158 10.6151
R1622 B.n587 B.n586 10.6151
R1623 B.n588 B.n587 10.6151
R1624 B.n588 B.n149 10.6151
R1625 B.n598 B.n149 10.6151
R1626 B.n599 B.n598 10.6151
R1627 B.n601 B.n599 10.6151
R1628 B.n601 B.n600 10.6151
R1629 B.n600 B.n142 10.6151
R1630 B.n612 B.n142 10.6151
R1631 B.n613 B.n612 10.6151
R1632 B.n614 B.n613 10.6151
R1633 B.n615 B.n614 10.6151
R1634 B.n616 B.n615 10.6151
R1635 B.n619 B.n616 10.6151
R1636 B.n620 B.n619 10.6151
R1637 B.n621 B.n620 10.6151
R1638 B.n622 B.n621 10.6151
R1639 B.n624 B.n622 10.6151
R1640 B.n625 B.n624 10.6151
R1641 B.n626 B.n625 10.6151
R1642 B.n627 B.n626 10.6151
R1643 B.n629 B.n627 10.6151
R1644 B.n630 B.n629 10.6151
R1645 B.n631 B.n630 10.6151
R1646 B.n632 B.n631 10.6151
R1647 B.n634 B.n632 10.6151
R1648 B.n635 B.n634 10.6151
R1649 B.n636 B.n635 10.6151
R1650 B.n637 B.n636 10.6151
R1651 B.n639 B.n637 10.6151
R1652 B.n640 B.n639 10.6151
R1653 B.n641 B.n640 10.6151
R1654 B.n642 B.n641 10.6151
R1655 B.n644 B.n642 10.6151
R1656 B.n645 B.n644 10.6151
R1657 B.n646 B.n645 10.6151
R1658 B.n647 B.n646 10.6151
R1659 B.n649 B.n647 10.6151
R1660 B.n650 B.n649 10.6151
R1661 B.n651 B.n650 10.6151
R1662 B.n652 B.n651 10.6151
R1663 B.n654 B.n652 10.6151
R1664 B.n655 B.n654 10.6151
R1665 B.n656 B.n655 10.6151
R1666 B.n657 B.n656 10.6151
R1667 B.n659 B.n657 10.6151
R1668 B.n660 B.n659 10.6151
R1669 B.n661 B.n660 10.6151
R1670 B.n662 B.n661 10.6151
R1671 B.n664 B.n662 10.6151
R1672 B.n665 B.n664 10.6151
R1673 B.n666 B.n665 10.6151
R1674 B.n667 B.n666 10.6151
R1675 B.n669 B.n667 10.6151
R1676 B.n670 B.n669 10.6151
R1677 B.n671 B.n670 10.6151
R1678 B.n672 B.n671 10.6151
R1679 B.n674 B.n672 10.6151
R1680 B.n675 B.n674 10.6151
R1681 B.n676 B.n675 10.6151
R1682 B.n677 B.n676 10.6151
R1683 B.n949 B.n1 10.6151
R1684 B.n949 B.n948 10.6151
R1685 B.n948 B.n947 10.6151
R1686 B.n947 B.n10 10.6151
R1687 B.n941 B.n10 10.6151
R1688 B.n941 B.n940 10.6151
R1689 B.n940 B.n939 10.6151
R1690 B.n939 B.n18 10.6151
R1691 B.n933 B.n18 10.6151
R1692 B.n933 B.n932 10.6151
R1693 B.n932 B.n931 10.6151
R1694 B.n931 B.n25 10.6151
R1695 B.n925 B.n25 10.6151
R1696 B.n925 B.n924 10.6151
R1697 B.n924 B.n923 10.6151
R1698 B.n923 B.n32 10.6151
R1699 B.n917 B.n32 10.6151
R1700 B.n917 B.n916 10.6151
R1701 B.n916 B.n915 10.6151
R1702 B.n915 B.n38 10.6151
R1703 B.n909 B.n38 10.6151
R1704 B.n909 B.n908 10.6151
R1705 B.n908 B.n907 10.6151
R1706 B.n907 B.n46 10.6151
R1707 B.n901 B.n46 10.6151
R1708 B.n901 B.n900 10.6151
R1709 B.n900 B.n899 10.6151
R1710 B.n899 B.n53 10.6151
R1711 B.n893 B.n53 10.6151
R1712 B.n893 B.n892 10.6151
R1713 B.n892 B.n891 10.6151
R1714 B.n891 B.n60 10.6151
R1715 B.n885 B.n60 10.6151
R1716 B.n885 B.n884 10.6151
R1717 B.n884 B.n883 10.6151
R1718 B.n883 B.n67 10.6151
R1719 B.n877 B.n67 10.6151
R1720 B.n877 B.n876 10.6151
R1721 B.n876 B.n875 10.6151
R1722 B.n875 B.n74 10.6151
R1723 B.n869 B.n74 10.6151
R1724 B.n869 B.n868 10.6151
R1725 B.n868 B.n867 10.6151
R1726 B.n867 B.n81 10.6151
R1727 B.n861 B.n81 10.6151
R1728 B.n861 B.n860 10.6151
R1729 B.n860 B.n859 10.6151
R1730 B.n859 B.n88 10.6151
R1731 B.n853 B.n88 10.6151
R1732 B.n852 B.n851 10.6151
R1733 B.n851 B.n95 10.6151
R1734 B.n845 B.n95 10.6151
R1735 B.n845 B.n844 10.6151
R1736 B.n844 B.n843 10.6151
R1737 B.n843 B.n97 10.6151
R1738 B.n837 B.n97 10.6151
R1739 B.n837 B.n836 10.6151
R1740 B.n836 B.n835 10.6151
R1741 B.n835 B.n99 10.6151
R1742 B.n829 B.n99 10.6151
R1743 B.n829 B.n828 10.6151
R1744 B.n828 B.n827 10.6151
R1745 B.n827 B.n101 10.6151
R1746 B.n821 B.n101 10.6151
R1747 B.n821 B.n820 10.6151
R1748 B.n820 B.n819 10.6151
R1749 B.n819 B.n103 10.6151
R1750 B.n813 B.n103 10.6151
R1751 B.n813 B.n812 10.6151
R1752 B.n812 B.n811 10.6151
R1753 B.n811 B.n105 10.6151
R1754 B.n805 B.n105 10.6151
R1755 B.n805 B.n804 10.6151
R1756 B.n804 B.n803 10.6151
R1757 B.n803 B.n107 10.6151
R1758 B.n797 B.n107 10.6151
R1759 B.n797 B.n796 10.6151
R1760 B.n796 B.n795 10.6151
R1761 B.n795 B.n109 10.6151
R1762 B.n789 B.n109 10.6151
R1763 B.n789 B.n788 10.6151
R1764 B.n788 B.n787 10.6151
R1765 B.n787 B.n111 10.6151
R1766 B.n781 B.n111 10.6151
R1767 B.n781 B.n780 10.6151
R1768 B.n780 B.n779 10.6151
R1769 B.n779 B.n113 10.6151
R1770 B.n773 B.n772 10.6151
R1771 B.n772 B.n771 10.6151
R1772 B.n771 B.n118 10.6151
R1773 B.n765 B.n118 10.6151
R1774 B.n765 B.n764 10.6151
R1775 B.n764 B.n763 10.6151
R1776 B.n763 B.n120 10.6151
R1777 B.n757 B.n120 10.6151
R1778 B.n755 B.n754 10.6151
R1779 B.n754 B.n124 10.6151
R1780 B.n748 B.n124 10.6151
R1781 B.n748 B.n747 10.6151
R1782 B.n747 B.n746 10.6151
R1783 B.n746 B.n126 10.6151
R1784 B.n740 B.n126 10.6151
R1785 B.n740 B.n739 10.6151
R1786 B.n739 B.n738 10.6151
R1787 B.n738 B.n128 10.6151
R1788 B.n732 B.n128 10.6151
R1789 B.n732 B.n731 10.6151
R1790 B.n731 B.n730 10.6151
R1791 B.n730 B.n130 10.6151
R1792 B.n724 B.n130 10.6151
R1793 B.n724 B.n723 10.6151
R1794 B.n723 B.n722 10.6151
R1795 B.n722 B.n132 10.6151
R1796 B.n716 B.n132 10.6151
R1797 B.n716 B.n715 10.6151
R1798 B.n715 B.n714 10.6151
R1799 B.n714 B.n134 10.6151
R1800 B.n708 B.n134 10.6151
R1801 B.n708 B.n707 10.6151
R1802 B.n707 B.n706 10.6151
R1803 B.n706 B.n136 10.6151
R1804 B.n700 B.n136 10.6151
R1805 B.n700 B.n699 10.6151
R1806 B.n699 B.n698 10.6151
R1807 B.n698 B.n138 10.6151
R1808 B.n692 B.n138 10.6151
R1809 B.n692 B.n691 10.6151
R1810 B.n691 B.n690 10.6151
R1811 B.n690 B.n140 10.6151
R1812 B.n684 B.n140 10.6151
R1813 B.n684 B.n683 10.6151
R1814 B.n683 B.n682 10.6151
R1815 B.n682 B.n678 10.6151
R1816 B.n535 B.t2 8.82494
R1817 B.t0 B.n903 8.82494
R1818 B.n957 B.n0 8.11757
R1819 B.n957 B.n1 8.11757
R1820 B.n383 B.n382 6.5566
R1821 B.n366 B.n365 6.5566
R1822 B.n773 B.n117 6.5566
R1823 B.n757 B.n756 6.5566
R1824 B.t11 B.n223 6.10973
R1825 B.n207 B.t3 6.10973
R1826 B.t7 B.n888 6.10973
R1827 B.t18 B.n79 6.10973
R1828 B.n384 B.n383 4.05904
R1829 B.n365 B.n364 4.05904
R1830 B.n117 B.n113 4.05904
R1831 B.n756 B.n755 4.05904
R1832 VN.n63 VN.n33 161.3
R1833 VN.n62 VN.n61 161.3
R1834 VN.n60 VN.n34 161.3
R1835 VN.n59 VN.n58 161.3
R1836 VN.n57 VN.n35 161.3
R1837 VN.n55 VN.n54 161.3
R1838 VN.n53 VN.n36 161.3
R1839 VN.n52 VN.n51 161.3
R1840 VN.n50 VN.n37 161.3
R1841 VN.n49 VN.n48 161.3
R1842 VN.n47 VN.n38 161.3
R1843 VN.n46 VN.n45 161.3
R1844 VN.n44 VN.n39 161.3
R1845 VN.n43 VN.n42 161.3
R1846 VN.n30 VN.n0 161.3
R1847 VN.n29 VN.n28 161.3
R1848 VN.n27 VN.n1 161.3
R1849 VN.n26 VN.n25 161.3
R1850 VN.n24 VN.n2 161.3
R1851 VN.n22 VN.n21 161.3
R1852 VN.n20 VN.n3 161.3
R1853 VN.n19 VN.n18 161.3
R1854 VN.n17 VN.n4 161.3
R1855 VN.n16 VN.n15 161.3
R1856 VN.n14 VN.n5 161.3
R1857 VN.n13 VN.n12 161.3
R1858 VN.n11 VN.n6 161.3
R1859 VN.n10 VN.n9 161.3
R1860 VN.n8 VN.t8 160.191
R1861 VN.n41 VN.t3 160.191
R1862 VN.n16 VN.t9 127.254
R1863 VN.n7 VN.t7 127.254
R1864 VN.n23 VN.t5 127.254
R1865 VN.n31 VN.t2 127.254
R1866 VN.n49 VN.t6 127.254
R1867 VN.n40 VN.t4 127.254
R1868 VN.n56 VN.t1 127.254
R1869 VN.n64 VN.t0 127.254
R1870 VN.n32 VN.n31 96.0763
R1871 VN.n65 VN.n64 96.0763
R1872 VN.n12 VN.n11 56.5193
R1873 VN.n18 VN.n3 56.5193
R1874 VN.n45 VN.n44 56.5193
R1875 VN.n51 VN.n36 56.5193
R1876 VN.n8 VN.n7 51.1767
R1877 VN.n41 VN.n40 51.1767
R1878 VN.n29 VN.n1 50.2061
R1879 VN.n62 VN.n34 50.2061
R1880 VN VN.n65 49.6648
R1881 VN.n25 VN.n1 30.7807
R1882 VN.n58 VN.n34 30.7807
R1883 VN.n11 VN.n10 24.4675
R1884 VN.n12 VN.n5 24.4675
R1885 VN.n16 VN.n5 24.4675
R1886 VN.n17 VN.n16 24.4675
R1887 VN.n18 VN.n17 24.4675
R1888 VN.n22 VN.n3 24.4675
R1889 VN.n25 VN.n24 24.4675
R1890 VN.n30 VN.n29 24.4675
R1891 VN.n44 VN.n43 24.4675
R1892 VN.n51 VN.n50 24.4675
R1893 VN.n50 VN.n49 24.4675
R1894 VN.n49 VN.n38 24.4675
R1895 VN.n45 VN.n38 24.4675
R1896 VN.n58 VN.n57 24.4675
R1897 VN.n55 VN.n36 24.4675
R1898 VN.n63 VN.n62 24.4675
R1899 VN.n10 VN.n7 19.5741
R1900 VN.n23 VN.n22 19.5741
R1901 VN.n43 VN.n40 19.5741
R1902 VN.n56 VN.n55 19.5741
R1903 VN.n31 VN.n30 14.6807
R1904 VN.n64 VN.n63 14.6807
R1905 VN.n42 VN.n41 9.46762
R1906 VN.n9 VN.n8 9.46762
R1907 VN.n24 VN.n23 4.8939
R1908 VN.n57 VN.n56 4.8939
R1909 VN.n65 VN.n33 0.278367
R1910 VN.n32 VN.n0 0.278367
R1911 VN.n61 VN.n33 0.189894
R1912 VN.n61 VN.n60 0.189894
R1913 VN.n60 VN.n59 0.189894
R1914 VN.n59 VN.n35 0.189894
R1915 VN.n54 VN.n35 0.189894
R1916 VN.n54 VN.n53 0.189894
R1917 VN.n53 VN.n52 0.189894
R1918 VN.n52 VN.n37 0.189894
R1919 VN.n48 VN.n37 0.189894
R1920 VN.n48 VN.n47 0.189894
R1921 VN.n47 VN.n46 0.189894
R1922 VN.n46 VN.n39 0.189894
R1923 VN.n42 VN.n39 0.189894
R1924 VN.n9 VN.n6 0.189894
R1925 VN.n13 VN.n6 0.189894
R1926 VN.n14 VN.n13 0.189894
R1927 VN.n15 VN.n14 0.189894
R1928 VN.n15 VN.n4 0.189894
R1929 VN.n19 VN.n4 0.189894
R1930 VN.n20 VN.n19 0.189894
R1931 VN.n21 VN.n20 0.189894
R1932 VN.n21 VN.n2 0.189894
R1933 VN.n26 VN.n2 0.189894
R1934 VN.n27 VN.n26 0.189894
R1935 VN.n28 VN.n27 0.189894
R1936 VN.n28 VN.n0 0.189894
R1937 VN VN.n32 0.153454
R1938 VDD2.n1 VDD2.t1 63.9561
R1939 VDD2.n4 VDD2.t9 61.8873
R1940 VDD2.n3 VDD2.n2 61.572
R1941 VDD2 VDD2.n7 61.5692
R1942 VDD2.n6 VDD2.n5 60.0758
R1943 VDD2.n1 VDD2.n0 60.0756
R1944 VDD2.n4 VDD2.n3 42.9653
R1945 VDD2.n6 VDD2.n4 2.06947
R1946 VDD2.n7 VDD2.t5 1.81203
R1947 VDD2.n7 VDD2.t6 1.81203
R1948 VDD2.n5 VDD2.t8 1.81203
R1949 VDD2.n5 VDD2.t3 1.81203
R1950 VDD2.n2 VDD2.t4 1.81203
R1951 VDD2.n2 VDD2.t7 1.81203
R1952 VDD2.n0 VDD2.t2 1.81203
R1953 VDD2.n0 VDD2.t0 1.81203
R1954 VDD2 VDD2.n6 0.575931
R1955 VDD2.n3 VDD2.n1 0.462395
C0 VDD1 VN 0.152175f
C1 VDD1 VDD2 1.82962f
C2 VDD1 VP 9.63905f
C3 VTAIL VDD1 9.86332f
C4 VDD2 VN 9.278981f
C5 VP VN 7.423f
C6 VDD2 VP 0.515924f
C7 VTAIL VN 9.745919f
C8 VTAIL VDD2 9.91035f
C9 VTAIL VP 9.760241f
C10 VDD2 B 6.375377f
C11 VDD1 B 6.364901f
C12 VTAIL B 7.372471f
C13 VN B 15.55959f
C14 VP B 14.050167f
C15 VDD2.t1 B 2.17474f
C16 VDD2.t2 B 0.191897f
C17 VDD2.t0 B 0.191897f
C18 VDD2.n0 B 1.69781f
C19 VDD2.n1 B 0.755098f
C20 VDD2.t4 B 0.191897f
C21 VDD2.t7 B 0.191897f
C22 VDD2.n2 B 1.70873f
C23 VDD2.n3 B 2.27834f
C24 VDD2.t9 B 2.16177f
C25 VDD2.n4 B 2.52201f
C26 VDD2.t8 B 0.191897f
C27 VDD2.t3 B 0.191897f
C28 VDD2.n5 B 1.69781f
C29 VDD2.n6 B 0.373961f
C30 VDD2.t5 B 0.191897f
C31 VDD2.t6 B 0.191897f
C32 VDD2.n7 B 1.70869f
C33 VN.n0 B 0.032867f
C34 VN.t2 B 1.53245f
C35 VN.n1 B 0.02355f
C36 VN.n2 B 0.024929f
C37 VN.t5 B 1.53245f
C38 VN.n3 B 0.039865f
C39 VN.n4 B 0.024929f
C40 VN.t9 B 1.53245f
C41 VN.n5 B 0.046461f
C42 VN.n6 B 0.024929f
C43 VN.t7 B 1.53245f
C44 VN.n7 B 0.618525f
C45 VN.t8 B 1.67196f
C46 VN.n8 B 0.606188f
C47 VN.n9 B 0.209069f
C48 VN.n10 B 0.041874f
C49 VN.n11 B 0.039865f
C50 VN.n12 B 0.032919f
C51 VN.n13 B 0.024929f
C52 VN.n14 B 0.024929f
C53 VN.n15 B 0.024929f
C54 VN.n16 B 0.573347f
C55 VN.n17 B 0.046461f
C56 VN.n18 B 0.032919f
C57 VN.n19 B 0.024929f
C58 VN.n20 B 0.024929f
C59 VN.n21 B 0.024929f
C60 VN.n22 B 0.041874f
C61 VN.n23 B 0.549823f
C62 VN.n24 B 0.028111f
C63 VN.n25 B 0.049942f
C64 VN.n26 B 0.024929f
C65 VN.n27 B 0.024929f
C66 VN.n28 B 0.024929f
C67 VN.n29 B 0.045754f
C68 VN.n30 B 0.037286f
C69 VN.n31 B 0.621506f
C70 VN.n32 B 0.03397f
C71 VN.n33 B 0.032867f
C72 VN.t0 B 1.53245f
C73 VN.n34 B 0.02355f
C74 VN.n35 B 0.024929f
C75 VN.t1 B 1.53245f
C76 VN.n36 B 0.039865f
C77 VN.n37 B 0.024929f
C78 VN.t6 B 1.53245f
C79 VN.n38 B 0.046461f
C80 VN.n39 B 0.024929f
C81 VN.t4 B 1.53245f
C82 VN.n40 B 0.618525f
C83 VN.t3 B 1.67196f
C84 VN.n41 B 0.606188f
C85 VN.n42 B 0.209069f
C86 VN.n43 B 0.041874f
C87 VN.n44 B 0.039865f
C88 VN.n45 B 0.032919f
C89 VN.n46 B 0.024929f
C90 VN.n47 B 0.024929f
C91 VN.n48 B 0.024929f
C92 VN.n49 B 0.573347f
C93 VN.n50 B 0.046461f
C94 VN.n51 B 0.032919f
C95 VN.n52 B 0.024929f
C96 VN.n53 B 0.024929f
C97 VN.n54 B 0.024929f
C98 VN.n55 B 0.041874f
C99 VN.n56 B 0.549823f
C100 VN.n57 B 0.028111f
C101 VN.n58 B 0.049942f
C102 VN.n59 B 0.024929f
C103 VN.n60 B 0.024929f
C104 VN.n61 B 0.024929f
C105 VN.n62 B 0.045754f
C106 VN.n63 B 0.037286f
C107 VN.n64 B 0.621506f
C108 VN.n65 B 1.36772f
C109 VDD1.t2 B 2.19933f
C110 VDD1.t3 B 0.194066f
C111 VDD1.t4 B 0.194066f
C112 VDD1.n0 B 1.717f
C113 VDD1.n1 B 0.770711f
C114 VDD1.t1 B 2.19932f
C115 VDD1.t0 B 0.194066f
C116 VDD1.t8 B 0.194066f
C117 VDD1.n2 B 1.717f
C118 VDD1.n3 B 0.763633f
C119 VDD1.t6 B 0.194066f
C120 VDD1.t7 B 0.194066f
C121 VDD1.n4 B 1.72804f
C122 VDD1.n5 B 2.40327f
C123 VDD1.t5 B 0.194066f
C124 VDD1.t9 B 0.194066f
C125 VDD1.n6 B 1.71699f
C126 VDD1.n7 B 2.58239f
C127 VTAIL.t4 B 0.215561f
C128 VTAIL.t5 B 0.215561f
C129 VTAIL.n0 B 1.82928f
C130 VTAIL.n1 B 0.501837f
C131 VTAIL.t12 B 2.32895f
C132 VTAIL.n2 B 0.626979f
C133 VTAIL.t10 B 0.215561f
C134 VTAIL.t16 B 0.215561f
C135 VTAIL.n3 B 1.82928f
C136 VTAIL.n4 B 0.584161f
C137 VTAIL.t17 B 0.215561f
C138 VTAIL.t15 B 0.215561f
C139 VTAIL.n5 B 1.82928f
C140 VTAIL.n6 B 1.84729f
C141 VTAIL.t3 B 0.215561f
C142 VTAIL.t2 B 0.215561f
C143 VTAIL.n7 B 1.82929f
C144 VTAIL.n8 B 1.84728f
C145 VTAIL.t6 B 0.215561f
C146 VTAIL.t8 B 0.215561f
C147 VTAIL.n9 B 1.82929f
C148 VTAIL.n10 B 0.584155f
C149 VTAIL.t1 B 2.32897f
C150 VTAIL.n11 B 0.626962f
C151 VTAIL.t19 B 0.215561f
C152 VTAIL.t13 B 0.215561f
C153 VTAIL.n12 B 1.82929f
C154 VTAIL.n13 B 0.538746f
C155 VTAIL.t14 B 0.215561f
C156 VTAIL.t11 B 0.215561f
C157 VTAIL.n14 B 1.82929f
C158 VTAIL.n15 B 0.584155f
C159 VTAIL.t18 B 2.32895f
C160 VTAIL.n16 B 1.76913f
C161 VTAIL.t7 B 2.32895f
C162 VTAIL.n17 B 1.76913f
C163 VTAIL.t9 B 0.215561f
C164 VTAIL.t0 B 0.215561f
C165 VTAIL.n18 B 1.82928f
C166 VTAIL.n19 B 0.454695f
C167 VP.n0 B 0.033409f
C168 VP.t2 B 1.55774f
C169 VP.n1 B 0.023939f
C170 VP.n2 B 0.02534f
C171 VP.t3 B 1.55774f
C172 VP.n3 B 0.040523f
C173 VP.n4 B 0.02534f
C174 VP.t1 B 1.55774f
C175 VP.n5 B 0.047228f
C176 VP.n6 B 0.02534f
C177 VP.t9 B 1.55774f
C178 VP.n7 B 0.558896f
C179 VP.n8 B 0.02534f
C180 VP.n9 B 0.046509f
C181 VP.n10 B 0.033409f
C182 VP.t0 B 1.55774f
C183 VP.n11 B 0.023939f
C184 VP.n12 B 0.02534f
C185 VP.t4 B 1.55774f
C186 VP.n13 B 0.040523f
C187 VP.n14 B 0.02534f
C188 VP.t5 B 1.55774f
C189 VP.n15 B 0.047228f
C190 VP.n16 B 0.02534f
C191 VP.t6 B 1.55774f
C192 VP.n17 B 0.628731f
C193 VP.t7 B 1.69955f
C194 VP.n18 B 0.61619f
C195 VP.n19 B 0.212518f
C196 VP.n20 B 0.042565f
C197 VP.n21 B 0.040523f
C198 VP.n22 B 0.033462f
C199 VP.n23 B 0.02534f
C200 VP.n24 B 0.02534f
C201 VP.n25 B 0.02534f
C202 VP.n26 B 0.582807f
C203 VP.n27 B 0.047228f
C204 VP.n28 B 0.033462f
C205 VP.n29 B 0.02534f
C206 VP.n30 B 0.02534f
C207 VP.n31 B 0.02534f
C208 VP.n32 B 0.042565f
C209 VP.n33 B 0.558896f
C210 VP.n34 B 0.028575f
C211 VP.n35 B 0.050766f
C212 VP.n36 B 0.02534f
C213 VP.n37 B 0.02534f
C214 VP.n38 B 0.02534f
C215 VP.n39 B 0.046509f
C216 VP.n40 B 0.037901f
C217 VP.n41 B 0.631761f
C218 VP.n42 B 1.37664f
C219 VP.n43 B 1.39508f
C220 VP.t8 B 1.55774f
C221 VP.n44 B 0.631761f
C222 VP.n45 B 0.037901f
C223 VP.n46 B 0.033409f
C224 VP.n47 B 0.02534f
C225 VP.n48 B 0.02534f
C226 VP.n49 B 0.023939f
C227 VP.n50 B 0.050766f
C228 VP.n51 B 0.028575f
C229 VP.n52 B 0.02534f
C230 VP.n53 B 0.02534f
C231 VP.n54 B 0.042565f
C232 VP.n55 B 0.040523f
C233 VP.n56 B 0.033462f
C234 VP.n57 B 0.02534f
C235 VP.n58 B 0.02534f
C236 VP.n59 B 0.02534f
C237 VP.n60 B 0.582807f
C238 VP.n61 B 0.047228f
C239 VP.n62 B 0.033462f
C240 VP.n63 B 0.02534f
C241 VP.n64 B 0.02534f
C242 VP.n65 B 0.02534f
C243 VP.n66 B 0.042565f
C244 VP.n67 B 0.558896f
C245 VP.n68 B 0.028575f
C246 VP.n69 B 0.050766f
C247 VP.n70 B 0.02534f
C248 VP.n71 B 0.02534f
C249 VP.n72 B 0.02534f
C250 VP.n73 B 0.046509f
C251 VP.n74 B 0.037901f
C252 VP.n75 B 0.631761f
C253 VP.n76 B 0.03453f
.ends

