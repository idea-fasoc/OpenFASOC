* NGSPICE file created from diff_pair_sample_1243.ext - technology: sky130A

.subckt diff_pair_sample_1243 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X1 VTAIL.t0 VN.t0 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X2 VTAIL.t8 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X3 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=3.0294 ps=18.69 w=18.36 l=0.36
X4 VDD2.t7 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X5 VDD1.t7 VP.t2 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X6 VDD1.t6 VP.t3 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=3.0294 ps=18.69 w=18.36 l=0.36
X7 VDD1.t5 VP.t4 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=3.0294 ps=18.69 w=18.36 l=0.36
X8 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=0 ps=0 w=18.36 l=0.36
X9 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=0 ps=0 w=18.36 l=0.36
X10 VTAIL.t4 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X11 VDD1.t4 VP.t5 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=7.1604 ps=37.5 w=18.36 l=0.36
X12 VDD2.t5 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X13 VTAIL.t12 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X14 VDD2.t4 VN.t5 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=7.1604 ps=37.5 w=18.36 l=0.36
X15 VDD2.t3 VN.t6 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=7.1604 ps=37.5 w=18.36 l=0.36
X16 VTAIL.t6 VP.t7 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X17 VTAIL.t10 VP.t8 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X18 VTAIL.t18 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
X19 VDD2.t1 VN.t8 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=3.0294 ps=18.69 w=18.36 l=0.36
X20 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=0 ps=0 w=18.36 l=0.36
X21 VDD1.t0 VP.t9 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=7.1604 ps=37.5 w=18.36 l=0.36
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1604 pd=37.5 as=0 ps=0 w=18.36 l=0.36
X23 VTAIL.t2 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0294 pd=18.69 as=3.0294 ps=18.69 w=18.36 l=0.36
R0 VP.n5 VP.t4 1359.2
R1 VP.n15 VP.t3 1338.22
R2 VP.n16 VP.t8 1338.22
R3 VP.n1 VP.t2 1338.22
R4 VP.n21 VP.t1 1338.22
R5 VP.n22 VP.t5 1338.22
R6 VP.n12 VP.t9 1338.22
R7 VP.n11 VP.t6 1338.22
R8 VP.n4 VP.t0 1338.22
R9 VP.n6 VP.t7 1338.22
R10 VP.n23 VP.n22 161.3
R11 VP.n8 VP.n7 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n11 VP.n3 161.3
R14 VP.n13 VP.n12 161.3
R15 VP.n21 VP.n0 161.3
R16 VP.n20 VP.n19 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n2 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n8 VP.n5 70.4033
R21 VP.n16 VP.n15 48.2005
R22 VP.n22 VP.n21 48.2005
R23 VP.n12 VP.n11 48.2005
R24 VP.n14 VP.n13 45.724
R25 VP.n17 VP.n16 37.9763
R26 VP.n21 VP.n20 37.9763
R27 VP.n11 VP.n10 37.9763
R28 VP.n7 VP.n6 37.9763
R29 VP.n6 VP.n5 20.9576
R30 VP.n17 VP.n1 10.2247
R31 VP.n20 VP.n1 10.2247
R32 VP.n10 VP.n4 10.2247
R33 VP.n7 VP.n4 10.2247
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n3 0.189894
R36 VP.n13 VP.n3 0.189894
R37 VP.n14 VP.n2 0.189894
R38 VP.n18 VP.n2 0.189894
R39 VP.n19 VP.n18 0.189894
R40 VP.n19 VP.n0 0.189894
R41 VP.n23 VP.n0 0.189894
R42 VP VP.n23 0.0516364
R43 VTAIL.n416 VTAIL.n320 289.615
R44 VTAIL.n98 VTAIL.n2 289.615
R45 VTAIL.n314 VTAIL.n218 289.615
R46 VTAIL.n208 VTAIL.n112 289.615
R47 VTAIL.n352 VTAIL.n351 185
R48 VTAIL.n357 VTAIL.n356 185
R49 VTAIL.n359 VTAIL.n358 185
R50 VTAIL.n348 VTAIL.n347 185
R51 VTAIL.n365 VTAIL.n364 185
R52 VTAIL.n367 VTAIL.n366 185
R53 VTAIL.n344 VTAIL.n343 185
R54 VTAIL.n373 VTAIL.n372 185
R55 VTAIL.n375 VTAIL.n374 185
R56 VTAIL.n340 VTAIL.n339 185
R57 VTAIL.n381 VTAIL.n380 185
R58 VTAIL.n383 VTAIL.n382 185
R59 VTAIL.n336 VTAIL.n335 185
R60 VTAIL.n389 VTAIL.n388 185
R61 VTAIL.n391 VTAIL.n390 185
R62 VTAIL.n332 VTAIL.n331 185
R63 VTAIL.n398 VTAIL.n397 185
R64 VTAIL.n399 VTAIL.n330 185
R65 VTAIL.n401 VTAIL.n400 185
R66 VTAIL.n328 VTAIL.n327 185
R67 VTAIL.n407 VTAIL.n406 185
R68 VTAIL.n409 VTAIL.n408 185
R69 VTAIL.n324 VTAIL.n323 185
R70 VTAIL.n415 VTAIL.n414 185
R71 VTAIL.n417 VTAIL.n416 185
R72 VTAIL.n34 VTAIL.n33 185
R73 VTAIL.n39 VTAIL.n38 185
R74 VTAIL.n41 VTAIL.n40 185
R75 VTAIL.n30 VTAIL.n29 185
R76 VTAIL.n47 VTAIL.n46 185
R77 VTAIL.n49 VTAIL.n48 185
R78 VTAIL.n26 VTAIL.n25 185
R79 VTAIL.n55 VTAIL.n54 185
R80 VTAIL.n57 VTAIL.n56 185
R81 VTAIL.n22 VTAIL.n21 185
R82 VTAIL.n63 VTAIL.n62 185
R83 VTAIL.n65 VTAIL.n64 185
R84 VTAIL.n18 VTAIL.n17 185
R85 VTAIL.n71 VTAIL.n70 185
R86 VTAIL.n73 VTAIL.n72 185
R87 VTAIL.n14 VTAIL.n13 185
R88 VTAIL.n80 VTAIL.n79 185
R89 VTAIL.n81 VTAIL.n12 185
R90 VTAIL.n83 VTAIL.n82 185
R91 VTAIL.n10 VTAIL.n9 185
R92 VTAIL.n89 VTAIL.n88 185
R93 VTAIL.n91 VTAIL.n90 185
R94 VTAIL.n6 VTAIL.n5 185
R95 VTAIL.n97 VTAIL.n96 185
R96 VTAIL.n99 VTAIL.n98 185
R97 VTAIL.n315 VTAIL.n314 185
R98 VTAIL.n313 VTAIL.n312 185
R99 VTAIL.n222 VTAIL.n221 185
R100 VTAIL.n307 VTAIL.n306 185
R101 VTAIL.n305 VTAIL.n304 185
R102 VTAIL.n226 VTAIL.n225 185
R103 VTAIL.n299 VTAIL.n298 185
R104 VTAIL.n297 VTAIL.n228 185
R105 VTAIL.n296 VTAIL.n295 185
R106 VTAIL.n231 VTAIL.n229 185
R107 VTAIL.n290 VTAIL.n289 185
R108 VTAIL.n288 VTAIL.n287 185
R109 VTAIL.n235 VTAIL.n234 185
R110 VTAIL.n282 VTAIL.n281 185
R111 VTAIL.n280 VTAIL.n279 185
R112 VTAIL.n239 VTAIL.n238 185
R113 VTAIL.n274 VTAIL.n273 185
R114 VTAIL.n272 VTAIL.n271 185
R115 VTAIL.n243 VTAIL.n242 185
R116 VTAIL.n266 VTAIL.n265 185
R117 VTAIL.n264 VTAIL.n263 185
R118 VTAIL.n247 VTAIL.n246 185
R119 VTAIL.n258 VTAIL.n257 185
R120 VTAIL.n256 VTAIL.n255 185
R121 VTAIL.n251 VTAIL.n250 185
R122 VTAIL.n209 VTAIL.n208 185
R123 VTAIL.n207 VTAIL.n206 185
R124 VTAIL.n116 VTAIL.n115 185
R125 VTAIL.n201 VTAIL.n200 185
R126 VTAIL.n199 VTAIL.n198 185
R127 VTAIL.n120 VTAIL.n119 185
R128 VTAIL.n193 VTAIL.n192 185
R129 VTAIL.n191 VTAIL.n122 185
R130 VTAIL.n190 VTAIL.n189 185
R131 VTAIL.n125 VTAIL.n123 185
R132 VTAIL.n184 VTAIL.n183 185
R133 VTAIL.n182 VTAIL.n181 185
R134 VTAIL.n129 VTAIL.n128 185
R135 VTAIL.n176 VTAIL.n175 185
R136 VTAIL.n174 VTAIL.n173 185
R137 VTAIL.n133 VTAIL.n132 185
R138 VTAIL.n168 VTAIL.n167 185
R139 VTAIL.n166 VTAIL.n165 185
R140 VTAIL.n137 VTAIL.n136 185
R141 VTAIL.n160 VTAIL.n159 185
R142 VTAIL.n158 VTAIL.n157 185
R143 VTAIL.n141 VTAIL.n140 185
R144 VTAIL.n152 VTAIL.n151 185
R145 VTAIL.n150 VTAIL.n149 185
R146 VTAIL.n145 VTAIL.n144 185
R147 VTAIL.n353 VTAIL.t16 147.659
R148 VTAIL.n35 VTAIL.t7 147.659
R149 VTAIL.n252 VTAIL.t13 147.659
R150 VTAIL.n146 VTAIL.t17 147.659
R151 VTAIL.n357 VTAIL.n351 104.615
R152 VTAIL.n358 VTAIL.n357 104.615
R153 VTAIL.n358 VTAIL.n347 104.615
R154 VTAIL.n365 VTAIL.n347 104.615
R155 VTAIL.n366 VTAIL.n365 104.615
R156 VTAIL.n366 VTAIL.n343 104.615
R157 VTAIL.n373 VTAIL.n343 104.615
R158 VTAIL.n374 VTAIL.n373 104.615
R159 VTAIL.n374 VTAIL.n339 104.615
R160 VTAIL.n381 VTAIL.n339 104.615
R161 VTAIL.n382 VTAIL.n381 104.615
R162 VTAIL.n382 VTAIL.n335 104.615
R163 VTAIL.n389 VTAIL.n335 104.615
R164 VTAIL.n390 VTAIL.n389 104.615
R165 VTAIL.n390 VTAIL.n331 104.615
R166 VTAIL.n398 VTAIL.n331 104.615
R167 VTAIL.n399 VTAIL.n398 104.615
R168 VTAIL.n400 VTAIL.n399 104.615
R169 VTAIL.n400 VTAIL.n327 104.615
R170 VTAIL.n407 VTAIL.n327 104.615
R171 VTAIL.n408 VTAIL.n407 104.615
R172 VTAIL.n408 VTAIL.n323 104.615
R173 VTAIL.n415 VTAIL.n323 104.615
R174 VTAIL.n416 VTAIL.n415 104.615
R175 VTAIL.n39 VTAIL.n33 104.615
R176 VTAIL.n40 VTAIL.n39 104.615
R177 VTAIL.n40 VTAIL.n29 104.615
R178 VTAIL.n47 VTAIL.n29 104.615
R179 VTAIL.n48 VTAIL.n47 104.615
R180 VTAIL.n48 VTAIL.n25 104.615
R181 VTAIL.n55 VTAIL.n25 104.615
R182 VTAIL.n56 VTAIL.n55 104.615
R183 VTAIL.n56 VTAIL.n21 104.615
R184 VTAIL.n63 VTAIL.n21 104.615
R185 VTAIL.n64 VTAIL.n63 104.615
R186 VTAIL.n64 VTAIL.n17 104.615
R187 VTAIL.n71 VTAIL.n17 104.615
R188 VTAIL.n72 VTAIL.n71 104.615
R189 VTAIL.n72 VTAIL.n13 104.615
R190 VTAIL.n80 VTAIL.n13 104.615
R191 VTAIL.n81 VTAIL.n80 104.615
R192 VTAIL.n82 VTAIL.n81 104.615
R193 VTAIL.n82 VTAIL.n9 104.615
R194 VTAIL.n89 VTAIL.n9 104.615
R195 VTAIL.n90 VTAIL.n89 104.615
R196 VTAIL.n90 VTAIL.n5 104.615
R197 VTAIL.n97 VTAIL.n5 104.615
R198 VTAIL.n98 VTAIL.n97 104.615
R199 VTAIL.n314 VTAIL.n313 104.615
R200 VTAIL.n313 VTAIL.n221 104.615
R201 VTAIL.n306 VTAIL.n221 104.615
R202 VTAIL.n306 VTAIL.n305 104.615
R203 VTAIL.n305 VTAIL.n225 104.615
R204 VTAIL.n298 VTAIL.n225 104.615
R205 VTAIL.n298 VTAIL.n297 104.615
R206 VTAIL.n297 VTAIL.n296 104.615
R207 VTAIL.n296 VTAIL.n229 104.615
R208 VTAIL.n289 VTAIL.n229 104.615
R209 VTAIL.n289 VTAIL.n288 104.615
R210 VTAIL.n288 VTAIL.n234 104.615
R211 VTAIL.n281 VTAIL.n234 104.615
R212 VTAIL.n281 VTAIL.n280 104.615
R213 VTAIL.n280 VTAIL.n238 104.615
R214 VTAIL.n273 VTAIL.n238 104.615
R215 VTAIL.n273 VTAIL.n272 104.615
R216 VTAIL.n272 VTAIL.n242 104.615
R217 VTAIL.n265 VTAIL.n242 104.615
R218 VTAIL.n265 VTAIL.n264 104.615
R219 VTAIL.n264 VTAIL.n246 104.615
R220 VTAIL.n257 VTAIL.n246 104.615
R221 VTAIL.n257 VTAIL.n256 104.615
R222 VTAIL.n256 VTAIL.n250 104.615
R223 VTAIL.n208 VTAIL.n207 104.615
R224 VTAIL.n207 VTAIL.n115 104.615
R225 VTAIL.n200 VTAIL.n115 104.615
R226 VTAIL.n200 VTAIL.n199 104.615
R227 VTAIL.n199 VTAIL.n119 104.615
R228 VTAIL.n192 VTAIL.n119 104.615
R229 VTAIL.n192 VTAIL.n191 104.615
R230 VTAIL.n191 VTAIL.n190 104.615
R231 VTAIL.n190 VTAIL.n123 104.615
R232 VTAIL.n183 VTAIL.n123 104.615
R233 VTAIL.n183 VTAIL.n182 104.615
R234 VTAIL.n182 VTAIL.n128 104.615
R235 VTAIL.n175 VTAIL.n128 104.615
R236 VTAIL.n175 VTAIL.n174 104.615
R237 VTAIL.n174 VTAIL.n132 104.615
R238 VTAIL.n167 VTAIL.n132 104.615
R239 VTAIL.n167 VTAIL.n166 104.615
R240 VTAIL.n166 VTAIL.n136 104.615
R241 VTAIL.n159 VTAIL.n136 104.615
R242 VTAIL.n159 VTAIL.n158 104.615
R243 VTAIL.n158 VTAIL.n140 104.615
R244 VTAIL.n151 VTAIL.n140 104.615
R245 VTAIL.n151 VTAIL.n150 104.615
R246 VTAIL.n150 VTAIL.n144 104.615
R247 VTAIL.t16 VTAIL.n351 52.3082
R248 VTAIL.t7 VTAIL.n33 52.3082
R249 VTAIL.t13 VTAIL.n250 52.3082
R250 VTAIL.t17 VTAIL.n144 52.3082
R251 VTAIL.n217 VTAIL.n216 46.2968
R252 VTAIL.n215 VTAIL.n214 46.2968
R253 VTAIL.n111 VTAIL.n110 46.2968
R254 VTAIL.n109 VTAIL.n108 46.2968
R255 VTAIL.n423 VTAIL.n422 46.2966
R256 VTAIL.n1 VTAIL.n0 46.2966
R257 VTAIL.n105 VTAIL.n104 46.2966
R258 VTAIL.n107 VTAIL.n106 46.2966
R259 VTAIL.n421 VTAIL.n420 34.5126
R260 VTAIL.n103 VTAIL.n102 34.5126
R261 VTAIL.n319 VTAIL.n318 34.5126
R262 VTAIL.n213 VTAIL.n212 34.5126
R263 VTAIL.n109 VTAIL.n107 29.3841
R264 VTAIL.n421 VTAIL.n319 28.7893
R265 VTAIL.n353 VTAIL.n352 15.6677
R266 VTAIL.n35 VTAIL.n34 15.6677
R267 VTAIL.n252 VTAIL.n251 15.6677
R268 VTAIL.n146 VTAIL.n145 15.6677
R269 VTAIL.n401 VTAIL.n330 13.1884
R270 VTAIL.n83 VTAIL.n12 13.1884
R271 VTAIL.n299 VTAIL.n228 13.1884
R272 VTAIL.n193 VTAIL.n122 13.1884
R273 VTAIL.n356 VTAIL.n355 12.8005
R274 VTAIL.n397 VTAIL.n396 12.8005
R275 VTAIL.n402 VTAIL.n328 12.8005
R276 VTAIL.n38 VTAIL.n37 12.8005
R277 VTAIL.n79 VTAIL.n78 12.8005
R278 VTAIL.n84 VTAIL.n10 12.8005
R279 VTAIL.n300 VTAIL.n226 12.8005
R280 VTAIL.n295 VTAIL.n230 12.8005
R281 VTAIL.n255 VTAIL.n254 12.8005
R282 VTAIL.n194 VTAIL.n120 12.8005
R283 VTAIL.n189 VTAIL.n124 12.8005
R284 VTAIL.n149 VTAIL.n148 12.8005
R285 VTAIL.n359 VTAIL.n350 12.0247
R286 VTAIL.n395 VTAIL.n332 12.0247
R287 VTAIL.n406 VTAIL.n405 12.0247
R288 VTAIL.n41 VTAIL.n32 12.0247
R289 VTAIL.n77 VTAIL.n14 12.0247
R290 VTAIL.n88 VTAIL.n87 12.0247
R291 VTAIL.n304 VTAIL.n303 12.0247
R292 VTAIL.n294 VTAIL.n231 12.0247
R293 VTAIL.n258 VTAIL.n249 12.0247
R294 VTAIL.n198 VTAIL.n197 12.0247
R295 VTAIL.n188 VTAIL.n125 12.0247
R296 VTAIL.n152 VTAIL.n143 12.0247
R297 VTAIL.n360 VTAIL.n348 11.249
R298 VTAIL.n392 VTAIL.n391 11.249
R299 VTAIL.n409 VTAIL.n326 11.249
R300 VTAIL.n42 VTAIL.n30 11.249
R301 VTAIL.n74 VTAIL.n73 11.249
R302 VTAIL.n91 VTAIL.n8 11.249
R303 VTAIL.n307 VTAIL.n224 11.249
R304 VTAIL.n291 VTAIL.n290 11.249
R305 VTAIL.n259 VTAIL.n247 11.249
R306 VTAIL.n201 VTAIL.n118 11.249
R307 VTAIL.n185 VTAIL.n184 11.249
R308 VTAIL.n153 VTAIL.n141 11.249
R309 VTAIL.n364 VTAIL.n363 10.4732
R310 VTAIL.n388 VTAIL.n334 10.4732
R311 VTAIL.n410 VTAIL.n324 10.4732
R312 VTAIL.n46 VTAIL.n45 10.4732
R313 VTAIL.n70 VTAIL.n16 10.4732
R314 VTAIL.n92 VTAIL.n6 10.4732
R315 VTAIL.n308 VTAIL.n222 10.4732
R316 VTAIL.n287 VTAIL.n233 10.4732
R317 VTAIL.n263 VTAIL.n262 10.4732
R318 VTAIL.n202 VTAIL.n116 10.4732
R319 VTAIL.n181 VTAIL.n127 10.4732
R320 VTAIL.n157 VTAIL.n156 10.4732
R321 VTAIL.n367 VTAIL.n346 9.69747
R322 VTAIL.n387 VTAIL.n336 9.69747
R323 VTAIL.n414 VTAIL.n413 9.69747
R324 VTAIL.n49 VTAIL.n28 9.69747
R325 VTAIL.n69 VTAIL.n18 9.69747
R326 VTAIL.n96 VTAIL.n95 9.69747
R327 VTAIL.n312 VTAIL.n311 9.69747
R328 VTAIL.n286 VTAIL.n235 9.69747
R329 VTAIL.n266 VTAIL.n245 9.69747
R330 VTAIL.n206 VTAIL.n205 9.69747
R331 VTAIL.n180 VTAIL.n129 9.69747
R332 VTAIL.n160 VTAIL.n139 9.69747
R333 VTAIL.n420 VTAIL.n419 9.45567
R334 VTAIL.n102 VTAIL.n101 9.45567
R335 VTAIL.n318 VTAIL.n317 9.45567
R336 VTAIL.n212 VTAIL.n211 9.45567
R337 VTAIL.n419 VTAIL.n418 9.3005
R338 VTAIL.n322 VTAIL.n321 9.3005
R339 VTAIL.n413 VTAIL.n412 9.3005
R340 VTAIL.n411 VTAIL.n410 9.3005
R341 VTAIL.n326 VTAIL.n325 9.3005
R342 VTAIL.n405 VTAIL.n404 9.3005
R343 VTAIL.n403 VTAIL.n402 9.3005
R344 VTAIL.n342 VTAIL.n341 9.3005
R345 VTAIL.n371 VTAIL.n370 9.3005
R346 VTAIL.n369 VTAIL.n368 9.3005
R347 VTAIL.n346 VTAIL.n345 9.3005
R348 VTAIL.n363 VTAIL.n362 9.3005
R349 VTAIL.n361 VTAIL.n360 9.3005
R350 VTAIL.n350 VTAIL.n349 9.3005
R351 VTAIL.n355 VTAIL.n354 9.3005
R352 VTAIL.n377 VTAIL.n376 9.3005
R353 VTAIL.n379 VTAIL.n378 9.3005
R354 VTAIL.n338 VTAIL.n337 9.3005
R355 VTAIL.n385 VTAIL.n384 9.3005
R356 VTAIL.n387 VTAIL.n386 9.3005
R357 VTAIL.n334 VTAIL.n333 9.3005
R358 VTAIL.n393 VTAIL.n392 9.3005
R359 VTAIL.n395 VTAIL.n394 9.3005
R360 VTAIL.n396 VTAIL.n329 9.3005
R361 VTAIL.n101 VTAIL.n100 9.3005
R362 VTAIL.n4 VTAIL.n3 9.3005
R363 VTAIL.n95 VTAIL.n94 9.3005
R364 VTAIL.n93 VTAIL.n92 9.3005
R365 VTAIL.n8 VTAIL.n7 9.3005
R366 VTAIL.n87 VTAIL.n86 9.3005
R367 VTAIL.n85 VTAIL.n84 9.3005
R368 VTAIL.n24 VTAIL.n23 9.3005
R369 VTAIL.n53 VTAIL.n52 9.3005
R370 VTAIL.n51 VTAIL.n50 9.3005
R371 VTAIL.n28 VTAIL.n27 9.3005
R372 VTAIL.n45 VTAIL.n44 9.3005
R373 VTAIL.n43 VTAIL.n42 9.3005
R374 VTAIL.n32 VTAIL.n31 9.3005
R375 VTAIL.n37 VTAIL.n36 9.3005
R376 VTAIL.n59 VTAIL.n58 9.3005
R377 VTAIL.n61 VTAIL.n60 9.3005
R378 VTAIL.n20 VTAIL.n19 9.3005
R379 VTAIL.n67 VTAIL.n66 9.3005
R380 VTAIL.n69 VTAIL.n68 9.3005
R381 VTAIL.n16 VTAIL.n15 9.3005
R382 VTAIL.n75 VTAIL.n74 9.3005
R383 VTAIL.n77 VTAIL.n76 9.3005
R384 VTAIL.n78 VTAIL.n11 9.3005
R385 VTAIL.n278 VTAIL.n277 9.3005
R386 VTAIL.n237 VTAIL.n236 9.3005
R387 VTAIL.n284 VTAIL.n283 9.3005
R388 VTAIL.n286 VTAIL.n285 9.3005
R389 VTAIL.n233 VTAIL.n232 9.3005
R390 VTAIL.n292 VTAIL.n291 9.3005
R391 VTAIL.n294 VTAIL.n293 9.3005
R392 VTAIL.n230 VTAIL.n227 9.3005
R393 VTAIL.n317 VTAIL.n316 9.3005
R394 VTAIL.n220 VTAIL.n219 9.3005
R395 VTAIL.n311 VTAIL.n310 9.3005
R396 VTAIL.n309 VTAIL.n308 9.3005
R397 VTAIL.n224 VTAIL.n223 9.3005
R398 VTAIL.n303 VTAIL.n302 9.3005
R399 VTAIL.n301 VTAIL.n300 9.3005
R400 VTAIL.n276 VTAIL.n275 9.3005
R401 VTAIL.n241 VTAIL.n240 9.3005
R402 VTAIL.n270 VTAIL.n269 9.3005
R403 VTAIL.n268 VTAIL.n267 9.3005
R404 VTAIL.n245 VTAIL.n244 9.3005
R405 VTAIL.n262 VTAIL.n261 9.3005
R406 VTAIL.n260 VTAIL.n259 9.3005
R407 VTAIL.n249 VTAIL.n248 9.3005
R408 VTAIL.n254 VTAIL.n253 9.3005
R409 VTAIL.n172 VTAIL.n171 9.3005
R410 VTAIL.n131 VTAIL.n130 9.3005
R411 VTAIL.n178 VTAIL.n177 9.3005
R412 VTAIL.n180 VTAIL.n179 9.3005
R413 VTAIL.n127 VTAIL.n126 9.3005
R414 VTAIL.n186 VTAIL.n185 9.3005
R415 VTAIL.n188 VTAIL.n187 9.3005
R416 VTAIL.n124 VTAIL.n121 9.3005
R417 VTAIL.n211 VTAIL.n210 9.3005
R418 VTAIL.n114 VTAIL.n113 9.3005
R419 VTAIL.n205 VTAIL.n204 9.3005
R420 VTAIL.n203 VTAIL.n202 9.3005
R421 VTAIL.n118 VTAIL.n117 9.3005
R422 VTAIL.n197 VTAIL.n196 9.3005
R423 VTAIL.n195 VTAIL.n194 9.3005
R424 VTAIL.n170 VTAIL.n169 9.3005
R425 VTAIL.n135 VTAIL.n134 9.3005
R426 VTAIL.n164 VTAIL.n163 9.3005
R427 VTAIL.n162 VTAIL.n161 9.3005
R428 VTAIL.n139 VTAIL.n138 9.3005
R429 VTAIL.n156 VTAIL.n155 9.3005
R430 VTAIL.n154 VTAIL.n153 9.3005
R431 VTAIL.n143 VTAIL.n142 9.3005
R432 VTAIL.n148 VTAIL.n147 9.3005
R433 VTAIL.n368 VTAIL.n344 8.92171
R434 VTAIL.n384 VTAIL.n383 8.92171
R435 VTAIL.n417 VTAIL.n322 8.92171
R436 VTAIL.n50 VTAIL.n26 8.92171
R437 VTAIL.n66 VTAIL.n65 8.92171
R438 VTAIL.n99 VTAIL.n4 8.92171
R439 VTAIL.n315 VTAIL.n220 8.92171
R440 VTAIL.n283 VTAIL.n282 8.92171
R441 VTAIL.n267 VTAIL.n243 8.92171
R442 VTAIL.n209 VTAIL.n114 8.92171
R443 VTAIL.n177 VTAIL.n176 8.92171
R444 VTAIL.n161 VTAIL.n137 8.92171
R445 VTAIL.n372 VTAIL.n371 8.14595
R446 VTAIL.n380 VTAIL.n338 8.14595
R447 VTAIL.n418 VTAIL.n320 8.14595
R448 VTAIL.n54 VTAIL.n53 8.14595
R449 VTAIL.n62 VTAIL.n20 8.14595
R450 VTAIL.n100 VTAIL.n2 8.14595
R451 VTAIL.n316 VTAIL.n218 8.14595
R452 VTAIL.n279 VTAIL.n237 8.14595
R453 VTAIL.n271 VTAIL.n270 8.14595
R454 VTAIL.n210 VTAIL.n112 8.14595
R455 VTAIL.n173 VTAIL.n131 8.14595
R456 VTAIL.n165 VTAIL.n164 8.14595
R457 VTAIL.n375 VTAIL.n342 7.3702
R458 VTAIL.n379 VTAIL.n340 7.3702
R459 VTAIL.n57 VTAIL.n24 7.3702
R460 VTAIL.n61 VTAIL.n22 7.3702
R461 VTAIL.n278 VTAIL.n239 7.3702
R462 VTAIL.n274 VTAIL.n241 7.3702
R463 VTAIL.n172 VTAIL.n133 7.3702
R464 VTAIL.n168 VTAIL.n135 7.3702
R465 VTAIL.n376 VTAIL.n375 6.59444
R466 VTAIL.n376 VTAIL.n340 6.59444
R467 VTAIL.n58 VTAIL.n57 6.59444
R468 VTAIL.n58 VTAIL.n22 6.59444
R469 VTAIL.n275 VTAIL.n239 6.59444
R470 VTAIL.n275 VTAIL.n274 6.59444
R471 VTAIL.n169 VTAIL.n133 6.59444
R472 VTAIL.n169 VTAIL.n168 6.59444
R473 VTAIL.n372 VTAIL.n342 5.81868
R474 VTAIL.n380 VTAIL.n379 5.81868
R475 VTAIL.n420 VTAIL.n320 5.81868
R476 VTAIL.n54 VTAIL.n24 5.81868
R477 VTAIL.n62 VTAIL.n61 5.81868
R478 VTAIL.n102 VTAIL.n2 5.81868
R479 VTAIL.n318 VTAIL.n218 5.81868
R480 VTAIL.n279 VTAIL.n278 5.81868
R481 VTAIL.n271 VTAIL.n241 5.81868
R482 VTAIL.n212 VTAIL.n112 5.81868
R483 VTAIL.n173 VTAIL.n172 5.81868
R484 VTAIL.n165 VTAIL.n135 5.81868
R485 VTAIL.n371 VTAIL.n344 5.04292
R486 VTAIL.n383 VTAIL.n338 5.04292
R487 VTAIL.n418 VTAIL.n417 5.04292
R488 VTAIL.n53 VTAIL.n26 5.04292
R489 VTAIL.n65 VTAIL.n20 5.04292
R490 VTAIL.n100 VTAIL.n99 5.04292
R491 VTAIL.n316 VTAIL.n315 5.04292
R492 VTAIL.n282 VTAIL.n237 5.04292
R493 VTAIL.n270 VTAIL.n243 5.04292
R494 VTAIL.n210 VTAIL.n209 5.04292
R495 VTAIL.n176 VTAIL.n131 5.04292
R496 VTAIL.n164 VTAIL.n137 5.04292
R497 VTAIL.n354 VTAIL.n353 4.38563
R498 VTAIL.n36 VTAIL.n35 4.38563
R499 VTAIL.n253 VTAIL.n252 4.38563
R500 VTAIL.n147 VTAIL.n146 4.38563
R501 VTAIL.n368 VTAIL.n367 4.26717
R502 VTAIL.n384 VTAIL.n336 4.26717
R503 VTAIL.n414 VTAIL.n322 4.26717
R504 VTAIL.n50 VTAIL.n49 4.26717
R505 VTAIL.n66 VTAIL.n18 4.26717
R506 VTAIL.n96 VTAIL.n4 4.26717
R507 VTAIL.n312 VTAIL.n220 4.26717
R508 VTAIL.n283 VTAIL.n235 4.26717
R509 VTAIL.n267 VTAIL.n266 4.26717
R510 VTAIL.n206 VTAIL.n114 4.26717
R511 VTAIL.n177 VTAIL.n129 4.26717
R512 VTAIL.n161 VTAIL.n160 4.26717
R513 VTAIL.n364 VTAIL.n346 3.49141
R514 VTAIL.n388 VTAIL.n387 3.49141
R515 VTAIL.n413 VTAIL.n324 3.49141
R516 VTAIL.n46 VTAIL.n28 3.49141
R517 VTAIL.n70 VTAIL.n69 3.49141
R518 VTAIL.n95 VTAIL.n6 3.49141
R519 VTAIL.n311 VTAIL.n222 3.49141
R520 VTAIL.n287 VTAIL.n286 3.49141
R521 VTAIL.n263 VTAIL.n245 3.49141
R522 VTAIL.n205 VTAIL.n116 3.49141
R523 VTAIL.n181 VTAIL.n180 3.49141
R524 VTAIL.n157 VTAIL.n139 3.49141
R525 VTAIL.n363 VTAIL.n348 2.71565
R526 VTAIL.n391 VTAIL.n334 2.71565
R527 VTAIL.n410 VTAIL.n409 2.71565
R528 VTAIL.n45 VTAIL.n30 2.71565
R529 VTAIL.n73 VTAIL.n16 2.71565
R530 VTAIL.n92 VTAIL.n91 2.71565
R531 VTAIL.n308 VTAIL.n307 2.71565
R532 VTAIL.n290 VTAIL.n233 2.71565
R533 VTAIL.n262 VTAIL.n247 2.71565
R534 VTAIL.n202 VTAIL.n201 2.71565
R535 VTAIL.n184 VTAIL.n127 2.71565
R536 VTAIL.n156 VTAIL.n141 2.71565
R537 VTAIL.n360 VTAIL.n359 1.93989
R538 VTAIL.n392 VTAIL.n332 1.93989
R539 VTAIL.n406 VTAIL.n326 1.93989
R540 VTAIL.n42 VTAIL.n41 1.93989
R541 VTAIL.n74 VTAIL.n14 1.93989
R542 VTAIL.n88 VTAIL.n8 1.93989
R543 VTAIL.n304 VTAIL.n224 1.93989
R544 VTAIL.n291 VTAIL.n231 1.93989
R545 VTAIL.n259 VTAIL.n258 1.93989
R546 VTAIL.n198 VTAIL.n118 1.93989
R547 VTAIL.n185 VTAIL.n125 1.93989
R548 VTAIL.n153 VTAIL.n152 1.93989
R549 VTAIL.n356 VTAIL.n350 1.16414
R550 VTAIL.n397 VTAIL.n395 1.16414
R551 VTAIL.n405 VTAIL.n328 1.16414
R552 VTAIL.n38 VTAIL.n32 1.16414
R553 VTAIL.n79 VTAIL.n77 1.16414
R554 VTAIL.n87 VTAIL.n10 1.16414
R555 VTAIL.n303 VTAIL.n226 1.16414
R556 VTAIL.n295 VTAIL.n294 1.16414
R557 VTAIL.n255 VTAIL.n249 1.16414
R558 VTAIL.n197 VTAIL.n120 1.16414
R559 VTAIL.n189 VTAIL.n188 1.16414
R560 VTAIL.n149 VTAIL.n143 1.16414
R561 VTAIL.n422 VTAIL.t1 1.07893
R562 VTAIL.n422 VTAIL.t0 1.07893
R563 VTAIL.n0 VTAIL.t19 1.07893
R564 VTAIL.n0 VTAIL.t4 1.07893
R565 VTAIL.n104 VTAIL.t14 1.07893
R566 VTAIL.n104 VTAIL.t8 1.07893
R567 VTAIL.n106 VTAIL.t15 1.07893
R568 VTAIL.n106 VTAIL.t10 1.07893
R569 VTAIL.n216 VTAIL.t11 1.07893
R570 VTAIL.n216 VTAIL.t12 1.07893
R571 VTAIL.n214 VTAIL.t9 1.07893
R572 VTAIL.n214 VTAIL.t6 1.07893
R573 VTAIL.n110 VTAIL.t3 1.07893
R574 VTAIL.n110 VTAIL.t2 1.07893
R575 VTAIL.n108 VTAIL.t5 1.07893
R576 VTAIL.n108 VTAIL.t18 1.07893
R577 VTAIL.n215 VTAIL.n213 0.767741
R578 VTAIL.n103 VTAIL.n1 0.767741
R579 VTAIL.n111 VTAIL.n109 0.595328
R580 VTAIL.n213 VTAIL.n111 0.595328
R581 VTAIL.n217 VTAIL.n215 0.595328
R582 VTAIL.n319 VTAIL.n217 0.595328
R583 VTAIL.n107 VTAIL.n105 0.595328
R584 VTAIL.n105 VTAIL.n103 0.595328
R585 VTAIL.n423 VTAIL.n421 0.595328
R586 VTAIL VTAIL.n1 0.50481
R587 VTAIL.n355 VTAIL.n352 0.388379
R588 VTAIL.n396 VTAIL.n330 0.388379
R589 VTAIL.n402 VTAIL.n401 0.388379
R590 VTAIL.n37 VTAIL.n34 0.388379
R591 VTAIL.n78 VTAIL.n12 0.388379
R592 VTAIL.n84 VTAIL.n83 0.388379
R593 VTAIL.n300 VTAIL.n299 0.388379
R594 VTAIL.n230 VTAIL.n228 0.388379
R595 VTAIL.n254 VTAIL.n251 0.388379
R596 VTAIL.n194 VTAIL.n193 0.388379
R597 VTAIL.n124 VTAIL.n122 0.388379
R598 VTAIL.n148 VTAIL.n145 0.388379
R599 VTAIL.n354 VTAIL.n349 0.155672
R600 VTAIL.n361 VTAIL.n349 0.155672
R601 VTAIL.n362 VTAIL.n361 0.155672
R602 VTAIL.n362 VTAIL.n345 0.155672
R603 VTAIL.n369 VTAIL.n345 0.155672
R604 VTAIL.n370 VTAIL.n369 0.155672
R605 VTAIL.n370 VTAIL.n341 0.155672
R606 VTAIL.n377 VTAIL.n341 0.155672
R607 VTAIL.n378 VTAIL.n377 0.155672
R608 VTAIL.n378 VTAIL.n337 0.155672
R609 VTAIL.n385 VTAIL.n337 0.155672
R610 VTAIL.n386 VTAIL.n385 0.155672
R611 VTAIL.n386 VTAIL.n333 0.155672
R612 VTAIL.n393 VTAIL.n333 0.155672
R613 VTAIL.n394 VTAIL.n393 0.155672
R614 VTAIL.n394 VTAIL.n329 0.155672
R615 VTAIL.n403 VTAIL.n329 0.155672
R616 VTAIL.n404 VTAIL.n403 0.155672
R617 VTAIL.n404 VTAIL.n325 0.155672
R618 VTAIL.n411 VTAIL.n325 0.155672
R619 VTAIL.n412 VTAIL.n411 0.155672
R620 VTAIL.n412 VTAIL.n321 0.155672
R621 VTAIL.n419 VTAIL.n321 0.155672
R622 VTAIL.n36 VTAIL.n31 0.155672
R623 VTAIL.n43 VTAIL.n31 0.155672
R624 VTAIL.n44 VTAIL.n43 0.155672
R625 VTAIL.n44 VTAIL.n27 0.155672
R626 VTAIL.n51 VTAIL.n27 0.155672
R627 VTAIL.n52 VTAIL.n51 0.155672
R628 VTAIL.n52 VTAIL.n23 0.155672
R629 VTAIL.n59 VTAIL.n23 0.155672
R630 VTAIL.n60 VTAIL.n59 0.155672
R631 VTAIL.n60 VTAIL.n19 0.155672
R632 VTAIL.n67 VTAIL.n19 0.155672
R633 VTAIL.n68 VTAIL.n67 0.155672
R634 VTAIL.n68 VTAIL.n15 0.155672
R635 VTAIL.n75 VTAIL.n15 0.155672
R636 VTAIL.n76 VTAIL.n75 0.155672
R637 VTAIL.n76 VTAIL.n11 0.155672
R638 VTAIL.n85 VTAIL.n11 0.155672
R639 VTAIL.n86 VTAIL.n85 0.155672
R640 VTAIL.n86 VTAIL.n7 0.155672
R641 VTAIL.n93 VTAIL.n7 0.155672
R642 VTAIL.n94 VTAIL.n93 0.155672
R643 VTAIL.n94 VTAIL.n3 0.155672
R644 VTAIL.n101 VTAIL.n3 0.155672
R645 VTAIL.n317 VTAIL.n219 0.155672
R646 VTAIL.n310 VTAIL.n219 0.155672
R647 VTAIL.n310 VTAIL.n309 0.155672
R648 VTAIL.n309 VTAIL.n223 0.155672
R649 VTAIL.n302 VTAIL.n223 0.155672
R650 VTAIL.n302 VTAIL.n301 0.155672
R651 VTAIL.n301 VTAIL.n227 0.155672
R652 VTAIL.n293 VTAIL.n227 0.155672
R653 VTAIL.n293 VTAIL.n292 0.155672
R654 VTAIL.n292 VTAIL.n232 0.155672
R655 VTAIL.n285 VTAIL.n232 0.155672
R656 VTAIL.n285 VTAIL.n284 0.155672
R657 VTAIL.n284 VTAIL.n236 0.155672
R658 VTAIL.n277 VTAIL.n236 0.155672
R659 VTAIL.n277 VTAIL.n276 0.155672
R660 VTAIL.n276 VTAIL.n240 0.155672
R661 VTAIL.n269 VTAIL.n240 0.155672
R662 VTAIL.n269 VTAIL.n268 0.155672
R663 VTAIL.n268 VTAIL.n244 0.155672
R664 VTAIL.n261 VTAIL.n244 0.155672
R665 VTAIL.n261 VTAIL.n260 0.155672
R666 VTAIL.n260 VTAIL.n248 0.155672
R667 VTAIL.n253 VTAIL.n248 0.155672
R668 VTAIL.n211 VTAIL.n113 0.155672
R669 VTAIL.n204 VTAIL.n113 0.155672
R670 VTAIL.n204 VTAIL.n203 0.155672
R671 VTAIL.n203 VTAIL.n117 0.155672
R672 VTAIL.n196 VTAIL.n117 0.155672
R673 VTAIL.n196 VTAIL.n195 0.155672
R674 VTAIL.n195 VTAIL.n121 0.155672
R675 VTAIL.n187 VTAIL.n121 0.155672
R676 VTAIL.n187 VTAIL.n186 0.155672
R677 VTAIL.n186 VTAIL.n126 0.155672
R678 VTAIL.n179 VTAIL.n126 0.155672
R679 VTAIL.n179 VTAIL.n178 0.155672
R680 VTAIL.n178 VTAIL.n130 0.155672
R681 VTAIL.n171 VTAIL.n130 0.155672
R682 VTAIL.n171 VTAIL.n170 0.155672
R683 VTAIL.n170 VTAIL.n134 0.155672
R684 VTAIL.n163 VTAIL.n134 0.155672
R685 VTAIL.n163 VTAIL.n162 0.155672
R686 VTAIL.n162 VTAIL.n138 0.155672
R687 VTAIL.n155 VTAIL.n138 0.155672
R688 VTAIL.n155 VTAIL.n154 0.155672
R689 VTAIL.n154 VTAIL.n142 0.155672
R690 VTAIL.n147 VTAIL.n142 0.155672
R691 VTAIL VTAIL.n423 0.0910172
R692 VDD1.n96 VDD1.n0 289.615
R693 VDD1.n199 VDD1.n103 289.615
R694 VDD1.n97 VDD1.n96 185
R695 VDD1.n95 VDD1.n94 185
R696 VDD1.n4 VDD1.n3 185
R697 VDD1.n89 VDD1.n88 185
R698 VDD1.n87 VDD1.n86 185
R699 VDD1.n8 VDD1.n7 185
R700 VDD1.n81 VDD1.n80 185
R701 VDD1.n79 VDD1.n10 185
R702 VDD1.n78 VDD1.n77 185
R703 VDD1.n13 VDD1.n11 185
R704 VDD1.n72 VDD1.n71 185
R705 VDD1.n70 VDD1.n69 185
R706 VDD1.n17 VDD1.n16 185
R707 VDD1.n64 VDD1.n63 185
R708 VDD1.n62 VDD1.n61 185
R709 VDD1.n21 VDD1.n20 185
R710 VDD1.n56 VDD1.n55 185
R711 VDD1.n54 VDD1.n53 185
R712 VDD1.n25 VDD1.n24 185
R713 VDD1.n48 VDD1.n47 185
R714 VDD1.n46 VDD1.n45 185
R715 VDD1.n29 VDD1.n28 185
R716 VDD1.n40 VDD1.n39 185
R717 VDD1.n38 VDD1.n37 185
R718 VDD1.n33 VDD1.n32 185
R719 VDD1.n135 VDD1.n134 185
R720 VDD1.n140 VDD1.n139 185
R721 VDD1.n142 VDD1.n141 185
R722 VDD1.n131 VDD1.n130 185
R723 VDD1.n148 VDD1.n147 185
R724 VDD1.n150 VDD1.n149 185
R725 VDD1.n127 VDD1.n126 185
R726 VDD1.n156 VDD1.n155 185
R727 VDD1.n158 VDD1.n157 185
R728 VDD1.n123 VDD1.n122 185
R729 VDD1.n164 VDD1.n163 185
R730 VDD1.n166 VDD1.n165 185
R731 VDD1.n119 VDD1.n118 185
R732 VDD1.n172 VDD1.n171 185
R733 VDD1.n174 VDD1.n173 185
R734 VDD1.n115 VDD1.n114 185
R735 VDD1.n181 VDD1.n180 185
R736 VDD1.n182 VDD1.n113 185
R737 VDD1.n184 VDD1.n183 185
R738 VDD1.n111 VDD1.n110 185
R739 VDD1.n190 VDD1.n189 185
R740 VDD1.n192 VDD1.n191 185
R741 VDD1.n107 VDD1.n106 185
R742 VDD1.n198 VDD1.n197 185
R743 VDD1.n200 VDD1.n199 185
R744 VDD1.n34 VDD1.t5 147.659
R745 VDD1.n136 VDD1.t6 147.659
R746 VDD1.n96 VDD1.n95 104.615
R747 VDD1.n95 VDD1.n3 104.615
R748 VDD1.n88 VDD1.n3 104.615
R749 VDD1.n88 VDD1.n87 104.615
R750 VDD1.n87 VDD1.n7 104.615
R751 VDD1.n80 VDD1.n7 104.615
R752 VDD1.n80 VDD1.n79 104.615
R753 VDD1.n79 VDD1.n78 104.615
R754 VDD1.n78 VDD1.n11 104.615
R755 VDD1.n71 VDD1.n11 104.615
R756 VDD1.n71 VDD1.n70 104.615
R757 VDD1.n70 VDD1.n16 104.615
R758 VDD1.n63 VDD1.n16 104.615
R759 VDD1.n63 VDD1.n62 104.615
R760 VDD1.n62 VDD1.n20 104.615
R761 VDD1.n55 VDD1.n20 104.615
R762 VDD1.n55 VDD1.n54 104.615
R763 VDD1.n54 VDD1.n24 104.615
R764 VDD1.n47 VDD1.n24 104.615
R765 VDD1.n47 VDD1.n46 104.615
R766 VDD1.n46 VDD1.n28 104.615
R767 VDD1.n39 VDD1.n28 104.615
R768 VDD1.n39 VDD1.n38 104.615
R769 VDD1.n38 VDD1.n32 104.615
R770 VDD1.n140 VDD1.n134 104.615
R771 VDD1.n141 VDD1.n140 104.615
R772 VDD1.n141 VDD1.n130 104.615
R773 VDD1.n148 VDD1.n130 104.615
R774 VDD1.n149 VDD1.n148 104.615
R775 VDD1.n149 VDD1.n126 104.615
R776 VDD1.n156 VDD1.n126 104.615
R777 VDD1.n157 VDD1.n156 104.615
R778 VDD1.n157 VDD1.n122 104.615
R779 VDD1.n164 VDD1.n122 104.615
R780 VDD1.n165 VDD1.n164 104.615
R781 VDD1.n165 VDD1.n118 104.615
R782 VDD1.n172 VDD1.n118 104.615
R783 VDD1.n173 VDD1.n172 104.615
R784 VDD1.n173 VDD1.n114 104.615
R785 VDD1.n181 VDD1.n114 104.615
R786 VDD1.n182 VDD1.n181 104.615
R787 VDD1.n183 VDD1.n182 104.615
R788 VDD1.n183 VDD1.n110 104.615
R789 VDD1.n190 VDD1.n110 104.615
R790 VDD1.n191 VDD1.n190 104.615
R791 VDD1.n191 VDD1.n106 104.615
R792 VDD1.n198 VDD1.n106 104.615
R793 VDD1.n199 VDD1.n198 104.615
R794 VDD1.n207 VDD1.n206 63.3662
R795 VDD1.n102 VDD1.n101 62.9756
R796 VDD1.n209 VDD1.n208 62.9754
R797 VDD1.n205 VDD1.n204 62.9754
R798 VDD1.t5 VDD1.n32 52.3082
R799 VDD1.t6 VDD1.n134 52.3082
R800 VDD1.n102 VDD1.n100 51.7862
R801 VDD1.n205 VDD1.n203 51.7862
R802 VDD1.n209 VDD1.n207 43.2487
R803 VDD1.n34 VDD1.n33 15.6677
R804 VDD1.n136 VDD1.n135 15.6677
R805 VDD1.n81 VDD1.n10 13.1884
R806 VDD1.n184 VDD1.n113 13.1884
R807 VDD1.n82 VDD1.n8 12.8005
R808 VDD1.n77 VDD1.n12 12.8005
R809 VDD1.n37 VDD1.n36 12.8005
R810 VDD1.n139 VDD1.n138 12.8005
R811 VDD1.n180 VDD1.n179 12.8005
R812 VDD1.n185 VDD1.n111 12.8005
R813 VDD1.n86 VDD1.n85 12.0247
R814 VDD1.n76 VDD1.n13 12.0247
R815 VDD1.n40 VDD1.n31 12.0247
R816 VDD1.n142 VDD1.n133 12.0247
R817 VDD1.n178 VDD1.n115 12.0247
R818 VDD1.n189 VDD1.n188 12.0247
R819 VDD1.n89 VDD1.n6 11.249
R820 VDD1.n73 VDD1.n72 11.249
R821 VDD1.n41 VDD1.n29 11.249
R822 VDD1.n143 VDD1.n131 11.249
R823 VDD1.n175 VDD1.n174 11.249
R824 VDD1.n192 VDD1.n109 11.249
R825 VDD1.n90 VDD1.n4 10.4732
R826 VDD1.n69 VDD1.n15 10.4732
R827 VDD1.n45 VDD1.n44 10.4732
R828 VDD1.n147 VDD1.n146 10.4732
R829 VDD1.n171 VDD1.n117 10.4732
R830 VDD1.n193 VDD1.n107 10.4732
R831 VDD1.n94 VDD1.n93 9.69747
R832 VDD1.n68 VDD1.n17 9.69747
R833 VDD1.n48 VDD1.n27 9.69747
R834 VDD1.n150 VDD1.n129 9.69747
R835 VDD1.n170 VDD1.n119 9.69747
R836 VDD1.n197 VDD1.n196 9.69747
R837 VDD1.n100 VDD1.n99 9.45567
R838 VDD1.n203 VDD1.n202 9.45567
R839 VDD1.n60 VDD1.n59 9.3005
R840 VDD1.n19 VDD1.n18 9.3005
R841 VDD1.n66 VDD1.n65 9.3005
R842 VDD1.n68 VDD1.n67 9.3005
R843 VDD1.n15 VDD1.n14 9.3005
R844 VDD1.n74 VDD1.n73 9.3005
R845 VDD1.n76 VDD1.n75 9.3005
R846 VDD1.n12 VDD1.n9 9.3005
R847 VDD1.n99 VDD1.n98 9.3005
R848 VDD1.n2 VDD1.n1 9.3005
R849 VDD1.n93 VDD1.n92 9.3005
R850 VDD1.n91 VDD1.n90 9.3005
R851 VDD1.n6 VDD1.n5 9.3005
R852 VDD1.n85 VDD1.n84 9.3005
R853 VDD1.n83 VDD1.n82 9.3005
R854 VDD1.n58 VDD1.n57 9.3005
R855 VDD1.n23 VDD1.n22 9.3005
R856 VDD1.n52 VDD1.n51 9.3005
R857 VDD1.n50 VDD1.n49 9.3005
R858 VDD1.n27 VDD1.n26 9.3005
R859 VDD1.n44 VDD1.n43 9.3005
R860 VDD1.n42 VDD1.n41 9.3005
R861 VDD1.n31 VDD1.n30 9.3005
R862 VDD1.n36 VDD1.n35 9.3005
R863 VDD1.n202 VDD1.n201 9.3005
R864 VDD1.n105 VDD1.n104 9.3005
R865 VDD1.n196 VDD1.n195 9.3005
R866 VDD1.n194 VDD1.n193 9.3005
R867 VDD1.n109 VDD1.n108 9.3005
R868 VDD1.n188 VDD1.n187 9.3005
R869 VDD1.n186 VDD1.n185 9.3005
R870 VDD1.n125 VDD1.n124 9.3005
R871 VDD1.n154 VDD1.n153 9.3005
R872 VDD1.n152 VDD1.n151 9.3005
R873 VDD1.n129 VDD1.n128 9.3005
R874 VDD1.n146 VDD1.n145 9.3005
R875 VDD1.n144 VDD1.n143 9.3005
R876 VDD1.n133 VDD1.n132 9.3005
R877 VDD1.n138 VDD1.n137 9.3005
R878 VDD1.n160 VDD1.n159 9.3005
R879 VDD1.n162 VDD1.n161 9.3005
R880 VDD1.n121 VDD1.n120 9.3005
R881 VDD1.n168 VDD1.n167 9.3005
R882 VDD1.n170 VDD1.n169 9.3005
R883 VDD1.n117 VDD1.n116 9.3005
R884 VDD1.n176 VDD1.n175 9.3005
R885 VDD1.n178 VDD1.n177 9.3005
R886 VDD1.n179 VDD1.n112 9.3005
R887 VDD1.n97 VDD1.n2 8.92171
R888 VDD1.n65 VDD1.n64 8.92171
R889 VDD1.n49 VDD1.n25 8.92171
R890 VDD1.n151 VDD1.n127 8.92171
R891 VDD1.n167 VDD1.n166 8.92171
R892 VDD1.n200 VDD1.n105 8.92171
R893 VDD1.n98 VDD1.n0 8.14595
R894 VDD1.n61 VDD1.n19 8.14595
R895 VDD1.n53 VDD1.n52 8.14595
R896 VDD1.n155 VDD1.n154 8.14595
R897 VDD1.n163 VDD1.n121 8.14595
R898 VDD1.n201 VDD1.n103 8.14595
R899 VDD1.n60 VDD1.n21 7.3702
R900 VDD1.n56 VDD1.n23 7.3702
R901 VDD1.n158 VDD1.n125 7.3702
R902 VDD1.n162 VDD1.n123 7.3702
R903 VDD1.n57 VDD1.n21 6.59444
R904 VDD1.n57 VDD1.n56 6.59444
R905 VDD1.n159 VDD1.n158 6.59444
R906 VDD1.n159 VDD1.n123 6.59444
R907 VDD1.n100 VDD1.n0 5.81868
R908 VDD1.n61 VDD1.n60 5.81868
R909 VDD1.n53 VDD1.n23 5.81868
R910 VDD1.n155 VDD1.n125 5.81868
R911 VDD1.n163 VDD1.n162 5.81868
R912 VDD1.n203 VDD1.n103 5.81868
R913 VDD1.n98 VDD1.n97 5.04292
R914 VDD1.n64 VDD1.n19 5.04292
R915 VDD1.n52 VDD1.n25 5.04292
R916 VDD1.n154 VDD1.n127 5.04292
R917 VDD1.n166 VDD1.n121 5.04292
R918 VDD1.n201 VDD1.n200 5.04292
R919 VDD1.n35 VDD1.n34 4.38563
R920 VDD1.n137 VDD1.n136 4.38563
R921 VDD1.n94 VDD1.n2 4.26717
R922 VDD1.n65 VDD1.n17 4.26717
R923 VDD1.n49 VDD1.n48 4.26717
R924 VDD1.n151 VDD1.n150 4.26717
R925 VDD1.n167 VDD1.n119 4.26717
R926 VDD1.n197 VDD1.n105 4.26717
R927 VDD1.n93 VDD1.n4 3.49141
R928 VDD1.n69 VDD1.n68 3.49141
R929 VDD1.n45 VDD1.n27 3.49141
R930 VDD1.n147 VDD1.n129 3.49141
R931 VDD1.n171 VDD1.n170 3.49141
R932 VDD1.n196 VDD1.n107 3.49141
R933 VDD1.n90 VDD1.n89 2.71565
R934 VDD1.n72 VDD1.n15 2.71565
R935 VDD1.n44 VDD1.n29 2.71565
R936 VDD1.n146 VDD1.n131 2.71565
R937 VDD1.n174 VDD1.n117 2.71565
R938 VDD1.n193 VDD1.n192 2.71565
R939 VDD1.n86 VDD1.n6 1.93989
R940 VDD1.n73 VDD1.n13 1.93989
R941 VDD1.n41 VDD1.n40 1.93989
R942 VDD1.n143 VDD1.n142 1.93989
R943 VDD1.n175 VDD1.n115 1.93989
R944 VDD1.n189 VDD1.n109 1.93989
R945 VDD1.n85 VDD1.n8 1.16414
R946 VDD1.n77 VDD1.n76 1.16414
R947 VDD1.n37 VDD1.n31 1.16414
R948 VDD1.n139 VDD1.n133 1.16414
R949 VDD1.n180 VDD1.n178 1.16414
R950 VDD1.n188 VDD1.n111 1.16414
R951 VDD1.n208 VDD1.t3 1.07893
R952 VDD1.n208 VDD1.t0 1.07893
R953 VDD1.n101 VDD1.t2 1.07893
R954 VDD1.n101 VDD1.t9 1.07893
R955 VDD1.n206 VDD1.t8 1.07893
R956 VDD1.n206 VDD1.t4 1.07893
R957 VDD1.n204 VDD1.t1 1.07893
R958 VDD1.n204 VDD1.t7 1.07893
R959 VDD1 VDD1.n209 0.388431
R960 VDD1.n82 VDD1.n81 0.388379
R961 VDD1.n12 VDD1.n10 0.388379
R962 VDD1.n36 VDD1.n33 0.388379
R963 VDD1.n138 VDD1.n135 0.388379
R964 VDD1.n179 VDD1.n113 0.388379
R965 VDD1.n185 VDD1.n184 0.388379
R966 VDD1 VDD1.n102 0.207397
R967 VDD1.n99 VDD1.n1 0.155672
R968 VDD1.n92 VDD1.n1 0.155672
R969 VDD1.n92 VDD1.n91 0.155672
R970 VDD1.n91 VDD1.n5 0.155672
R971 VDD1.n84 VDD1.n5 0.155672
R972 VDD1.n84 VDD1.n83 0.155672
R973 VDD1.n83 VDD1.n9 0.155672
R974 VDD1.n75 VDD1.n9 0.155672
R975 VDD1.n75 VDD1.n74 0.155672
R976 VDD1.n74 VDD1.n14 0.155672
R977 VDD1.n67 VDD1.n14 0.155672
R978 VDD1.n67 VDD1.n66 0.155672
R979 VDD1.n66 VDD1.n18 0.155672
R980 VDD1.n59 VDD1.n18 0.155672
R981 VDD1.n59 VDD1.n58 0.155672
R982 VDD1.n58 VDD1.n22 0.155672
R983 VDD1.n51 VDD1.n22 0.155672
R984 VDD1.n51 VDD1.n50 0.155672
R985 VDD1.n50 VDD1.n26 0.155672
R986 VDD1.n43 VDD1.n26 0.155672
R987 VDD1.n43 VDD1.n42 0.155672
R988 VDD1.n42 VDD1.n30 0.155672
R989 VDD1.n35 VDD1.n30 0.155672
R990 VDD1.n137 VDD1.n132 0.155672
R991 VDD1.n144 VDD1.n132 0.155672
R992 VDD1.n145 VDD1.n144 0.155672
R993 VDD1.n145 VDD1.n128 0.155672
R994 VDD1.n152 VDD1.n128 0.155672
R995 VDD1.n153 VDD1.n152 0.155672
R996 VDD1.n153 VDD1.n124 0.155672
R997 VDD1.n160 VDD1.n124 0.155672
R998 VDD1.n161 VDD1.n160 0.155672
R999 VDD1.n161 VDD1.n120 0.155672
R1000 VDD1.n168 VDD1.n120 0.155672
R1001 VDD1.n169 VDD1.n168 0.155672
R1002 VDD1.n169 VDD1.n116 0.155672
R1003 VDD1.n176 VDD1.n116 0.155672
R1004 VDD1.n177 VDD1.n176 0.155672
R1005 VDD1.n177 VDD1.n112 0.155672
R1006 VDD1.n186 VDD1.n112 0.155672
R1007 VDD1.n187 VDD1.n186 0.155672
R1008 VDD1.n187 VDD1.n108 0.155672
R1009 VDD1.n194 VDD1.n108 0.155672
R1010 VDD1.n195 VDD1.n194 0.155672
R1011 VDD1.n195 VDD1.n104 0.155672
R1012 VDD1.n202 VDD1.n104 0.155672
R1013 VDD1.n207 VDD1.n205 0.0938609
R1014 B.n607 B.t14 1440.19
R1015 B.n439 B.t18 1440.19
R1016 B.n109 B.t10 1440.19
R1017 B.n106 B.t21 1440.19
R1018 B.n822 B.n821 585
R1019 B.n366 B.n105 585
R1020 B.n365 B.n364 585
R1021 B.n363 B.n362 585
R1022 B.n361 B.n360 585
R1023 B.n359 B.n358 585
R1024 B.n357 B.n356 585
R1025 B.n355 B.n354 585
R1026 B.n353 B.n352 585
R1027 B.n351 B.n350 585
R1028 B.n349 B.n348 585
R1029 B.n347 B.n346 585
R1030 B.n345 B.n344 585
R1031 B.n343 B.n342 585
R1032 B.n341 B.n340 585
R1033 B.n339 B.n338 585
R1034 B.n337 B.n336 585
R1035 B.n335 B.n334 585
R1036 B.n333 B.n332 585
R1037 B.n331 B.n330 585
R1038 B.n329 B.n328 585
R1039 B.n327 B.n326 585
R1040 B.n325 B.n324 585
R1041 B.n323 B.n322 585
R1042 B.n321 B.n320 585
R1043 B.n319 B.n318 585
R1044 B.n317 B.n316 585
R1045 B.n315 B.n314 585
R1046 B.n313 B.n312 585
R1047 B.n311 B.n310 585
R1048 B.n309 B.n308 585
R1049 B.n307 B.n306 585
R1050 B.n305 B.n304 585
R1051 B.n303 B.n302 585
R1052 B.n301 B.n300 585
R1053 B.n299 B.n298 585
R1054 B.n297 B.n296 585
R1055 B.n295 B.n294 585
R1056 B.n293 B.n292 585
R1057 B.n291 B.n290 585
R1058 B.n289 B.n288 585
R1059 B.n287 B.n286 585
R1060 B.n285 B.n284 585
R1061 B.n283 B.n282 585
R1062 B.n281 B.n280 585
R1063 B.n279 B.n278 585
R1064 B.n277 B.n276 585
R1065 B.n275 B.n274 585
R1066 B.n273 B.n272 585
R1067 B.n271 B.n270 585
R1068 B.n269 B.n268 585
R1069 B.n267 B.n266 585
R1070 B.n265 B.n264 585
R1071 B.n263 B.n262 585
R1072 B.n261 B.n260 585
R1073 B.n259 B.n258 585
R1074 B.n257 B.n256 585
R1075 B.n255 B.n254 585
R1076 B.n253 B.n252 585
R1077 B.n251 B.n250 585
R1078 B.n249 B.n248 585
R1079 B.n247 B.n246 585
R1080 B.n245 B.n244 585
R1081 B.n243 B.n242 585
R1082 B.n241 B.n240 585
R1083 B.n239 B.n238 585
R1084 B.n237 B.n236 585
R1085 B.n235 B.n234 585
R1086 B.n233 B.n232 585
R1087 B.n231 B.n230 585
R1088 B.n229 B.n228 585
R1089 B.n227 B.n226 585
R1090 B.n225 B.n224 585
R1091 B.n223 B.n222 585
R1092 B.n221 B.n220 585
R1093 B.n219 B.n218 585
R1094 B.n217 B.n216 585
R1095 B.n215 B.n214 585
R1096 B.n213 B.n212 585
R1097 B.n211 B.n210 585
R1098 B.n209 B.n208 585
R1099 B.n207 B.n206 585
R1100 B.n205 B.n204 585
R1101 B.n203 B.n202 585
R1102 B.n201 B.n200 585
R1103 B.n199 B.n198 585
R1104 B.n197 B.n196 585
R1105 B.n195 B.n194 585
R1106 B.n193 B.n192 585
R1107 B.n191 B.n190 585
R1108 B.n189 B.n188 585
R1109 B.n187 B.n186 585
R1110 B.n185 B.n184 585
R1111 B.n183 B.n182 585
R1112 B.n181 B.n180 585
R1113 B.n179 B.n178 585
R1114 B.n177 B.n176 585
R1115 B.n175 B.n174 585
R1116 B.n173 B.n172 585
R1117 B.n171 B.n170 585
R1118 B.n169 B.n168 585
R1119 B.n167 B.n166 585
R1120 B.n165 B.n164 585
R1121 B.n163 B.n162 585
R1122 B.n161 B.n160 585
R1123 B.n159 B.n158 585
R1124 B.n157 B.n156 585
R1125 B.n155 B.n154 585
R1126 B.n153 B.n152 585
R1127 B.n151 B.n150 585
R1128 B.n149 B.n148 585
R1129 B.n147 B.n146 585
R1130 B.n145 B.n144 585
R1131 B.n143 B.n142 585
R1132 B.n141 B.n140 585
R1133 B.n139 B.n138 585
R1134 B.n137 B.n136 585
R1135 B.n135 B.n134 585
R1136 B.n133 B.n132 585
R1137 B.n131 B.n130 585
R1138 B.n129 B.n128 585
R1139 B.n127 B.n126 585
R1140 B.n125 B.n124 585
R1141 B.n123 B.n122 585
R1142 B.n121 B.n120 585
R1143 B.n119 B.n118 585
R1144 B.n117 B.n116 585
R1145 B.n115 B.n114 585
R1146 B.n113 B.n112 585
R1147 B.n39 B.n38 585
R1148 B.n820 B.n40 585
R1149 B.n825 B.n40 585
R1150 B.n819 B.n818 585
R1151 B.n818 B.n36 585
R1152 B.n817 B.n35 585
R1153 B.n831 B.n35 585
R1154 B.n816 B.n34 585
R1155 B.n832 B.n34 585
R1156 B.n815 B.n33 585
R1157 B.n833 B.n33 585
R1158 B.n814 B.n813 585
R1159 B.n813 B.n29 585
R1160 B.n812 B.n28 585
R1161 B.n839 B.n28 585
R1162 B.n811 B.n27 585
R1163 B.n840 B.n27 585
R1164 B.n810 B.n26 585
R1165 B.n841 B.n26 585
R1166 B.n809 B.n808 585
R1167 B.n808 B.n25 585
R1168 B.n807 B.n21 585
R1169 B.n847 B.n21 585
R1170 B.n806 B.n20 585
R1171 B.n848 B.n20 585
R1172 B.n805 B.n19 585
R1173 B.n849 B.n19 585
R1174 B.n804 B.n803 585
R1175 B.n803 B.n18 585
R1176 B.n802 B.n14 585
R1177 B.n855 B.n14 585
R1178 B.n801 B.n13 585
R1179 B.n856 B.n13 585
R1180 B.n800 B.n12 585
R1181 B.n857 B.n12 585
R1182 B.n799 B.n798 585
R1183 B.n798 B.n11 585
R1184 B.n797 B.n7 585
R1185 B.n863 B.n7 585
R1186 B.n796 B.n6 585
R1187 B.n864 B.n6 585
R1188 B.n795 B.n5 585
R1189 B.n865 B.n5 585
R1190 B.n794 B.n793 585
R1191 B.n793 B.n4 585
R1192 B.n792 B.n367 585
R1193 B.n792 B.n791 585
R1194 B.n781 B.n368 585
R1195 B.n784 B.n368 585
R1196 B.n783 B.n782 585
R1197 B.n785 B.n783 585
R1198 B.n780 B.n372 585
R1199 B.n375 B.n372 585
R1200 B.n779 B.n778 585
R1201 B.n778 B.n777 585
R1202 B.n374 B.n373 585
R1203 B.n770 B.n374 585
R1204 B.n769 B.n768 585
R1205 B.n771 B.n769 585
R1206 B.n767 B.n379 585
R1207 B.n382 B.n379 585
R1208 B.n766 B.n765 585
R1209 B.n765 B.n764 585
R1210 B.n381 B.n380 585
R1211 B.n757 B.n381 585
R1212 B.n756 B.n755 585
R1213 B.n758 B.n756 585
R1214 B.n754 B.n387 585
R1215 B.n387 B.n386 585
R1216 B.n753 B.n752 585
R1217 B.n752 B.n751 585
R1218 B.n389 B.n388 585
R1219 B.n390 B.n389 585
R1220 B.n744 B.n743 585
R1221 B.n745 B.n744 585
R1222 B.n742 B.n395 585
R1223 B.n395 B.n394 585
R1224 B.n741 B.n740 585
R1225 B.n740 B.n739 585
R1226 B.n397 B.n396 585
R1227 B.n398 B.n397 585
R1228 B.n732 B.n731 585
R1229 B.n733 B.n732 585
R1230 B.n401 B.n400 585
R1231 B.n472 B.n470 585
R1232 B.n473 B.n469 585
R1233 B.n473 B.n402 585
R1234 B.n476 B.n475 585
R1235 B.n477 B.n468 585
R1236 B.n479 B.n478 585
R1237 B.n481 B.n467 585
R1238 B.n484 B.n483 585
R1239 B.n485 B.n466 585
R1240 B.n487 B.n486 585
R1241 B.n489 B.n465 585
R1242 B.n492 B.n491 585
R1243 B.n493 B.n464 585
R1244 B.n495 B.n494 585
R1245 B.n497 B.n463 585
R1246 B.n500 B.n499 585
R1247 B.n501 B.n462 585
R1248 B.n503 B.n502 585
R1249 B.n505 B.n461 585
R1250 B.n508 B.n507 585
R1251 B.n509 B.n460 585
R1252 B.n511 B.n510 585
R1253 B.n513 B.n459 585
R1254 B.n516 B.n515 585
R1255 B.n517 B.n458 585
R1256 B.n519 B.n518 585
R1257 B.n521 B.n457 585
R1258 B.n524 B.n523 585
R1259 B.n525 B.n456 585
R1260 B.n527 B.n526 585
R1261 B.n529 B.n455 585
R1262 B.n532 B.n531 585
R1263 B.n533 B.n454 585
R1264 B.n535 B.n534 585
R1265 B.n537 B.n453 585
R1266 B.n540 B.n539 585
R1267 B.n541 B.n452 585
R1268 B.n543 B.n542 585
R1269 B.n545 B.n451 585
R1270 B.n548 B.n547 585
R1271 B.n549 B.n450 585
R1272 B.n551 B.n550 585
R1273 B.n553 B.n449 585
R1274 B.n556 B.n555 585
R1275 B.n557 B.n448 585
R1276 B.n559 B.n558 585
R1277 B.n561 B.n447 585
R1278 B.n564 B.n563 585
R1279 B.n565 B.n446 585
R1280 B.n567 B.n566 585
R1281 B.n569 B.n445 585
R1282 B.n572 B.n571 585
R1283 B.n573 B.n444 585
R1284 B.n575 B.n574 585
R1285 B.n577 B.n443 585
R1286 B.n580 B.n579 585
R1287 B.n581 B.n442 585
R1288 B.n583 B.n582 585
R1289 B.n585 B.n441 585
R1290 B.n588 B.n587 585
R1291 B.n590 B.n438 585
R1292 B.n592 B.n591 585
R1293 B.n594 B.n437 585
R1294 B.n597 B.n596 585
R1295 B.n598 B.n436 585
R1296 B.n600 B.n599 585
R1297 B.n602 B.n435 585
R1298 B.n605 B.n604 585
R1299 B.n606 B.n434 585
R1300 B.n611 B.n610 585
R1301 B.n613 B.n433 585
R1302 B.n616 B.n615 585
R1303 B.n617 B.n432 585
R1304 B.n619 B.n618 585
R1305 B.n621 B.n431 585
R1306 B.n624 B.n623 585
R1307 B.n625 B.n430 585
R1308 B.n627 B.n626 585
R1309 B.n629 B.n429 585
R1310 B.n632 B.n631 585
R1311 B.n633 B.n428 585
R1312 B.n635 B.n634 585
R1313 B.n637 B.n427 585
R1314 B.n640 B.n639 585
R1315 B.n641 B.n426 585
R1316 B.n643 B.n642 585
R1317 B.n645 B.n425 585
R1318 B.n648 B.n647 585
R1319 B.n649 B.n424 585
R1320 B.n651 B.n650 585
R1321 B.n653 B.n423 585
R1322 B.n656 B.n655 585
R1323 B.n657 B.n422 585
R1324 B.n659 B.n658 585
R1325 B.n661 B.n421 585
R1326 B.n664 B.n663 585
R1327 B.n665 B.n420 585
R1328 B.n667 B.n666 585
R1329 B.n669 B.n419 585
R1330 B.n672 B.n671 585
R1331 B.n673 B.n418 585
R1332 B.n675 B.n674 585
R1333 B.n677 B.n417 585
R1334 B.n680 B.n679 585
R1335 B.n681 B.n416 585
R1336 B.n683 B.n682 585
R1337 B.n685 B.n415 585
R1338 B.n688 B.n687 585
R1339 B.n689 B.n414 585
R1340 B.n691 B.n690 585
R1341 B.n693 B.n413 585
R1342 B.n696 B.n695 585
R1343 B.n697 B.n412 585
R1344 B.n699 B.n698 585
R1345 B.n701 B.n411 585
R1346 B.n704 B.n703 585
R1347 B.n705 B.n410 585
R1348 B.n707 B.n706 585
R1349 B.n709 B.n409 585
R1350 B.n712 B.n711 585
R1351 B.n713 B.n408 585
R1352 B.n715 B.n714 585
R1353 B.n717 B.n407 585
R1354 B.n720 B.n719 585
R1355 B.n721 B.n406 585
R1356 B.n723 B.n722 585
R1357 B.n725 B.n405 585
R1358 B.n726 B.n404 585
R1359 B.n729 B.n728 585
R1360 B.n730 B.n403 585
R1361 B.n403 B.n402 585
R1362 B.n735 B.n734 585
R1363 B.n734 B.n733 585
R1364 B.n736 B.n399 585
R1365 B.n399 B.n398 585
R1366 B.n738 B.n737 585
R1367 B.n739 B.n738 585
R1368 B.n393 B.n392 585
R1369 B.n394 B.n393 585
R1370 B.n747 B.n746 585
R1371 B.n746 B.n745 585
R1372 B.n748 B.n391 585
R1373 B.n391 B.n390 585
R1374 B.n750 B.n749 585
R1375 B.n751 B.n750 585
R1376 B.n385 B.n384 585
R1377 B.n386 B.n385 585
R1378 B.n760 B.n759 585
R1379 B.n759 B.n758 585
R1380 B.n761 B.n383 585
R1381 B.n757 B.n383 585
R1382 B.n763 B.n762 585
R1383 B.n764 B.n763 585
R1384 B.n378 B.n377 585
R1385 B.n382 B.n378 585
R1386 B.n773 B.n772 585
R1387 B.n772 B.n771 585
R1388 B.n774 B.n376 585
R1389 B.n770 B.n376 585
R1390 B.n776 B.n775 585
R1391 B.n777 B.n776 585
R1392 B.n371 B.n370 585
R1393 B.n375 B.n371 585
R1394 B.n787 B.n786 585
R1395 B.n786 B.n785 585
R1396 B.n788 B.n369 585
R1397 B.n784 B.n369 585
R1398 B.n790 B.n789 585
R1399 B.n791 B.n790 585
R1400 B.n2 B.n0 585
R1401 B.n4 B.n2 585
R1402 B.n3 B.n1 585
R1403 B.n864 B.n3 585
R1404 B.n862 B.n861 585
R1405 B.n863 B.n862 585
R1406 B.n860 B.n8 585
R1407 B.n11 B.n8 585
R1408 B.n859 B.n858 585
R1409 B.n858 B.n857 585
R1410 B.n10 B.n9 585
R1411 B.n856 B.n10 585
R1412 B.n854 B.n853 585
R1413 B.n855 B.n854 585
R1414 B.n852 B.n15 585
R1415 B.n18 B.n15 585
R1416 B.n851 B.n850 585
R1417 B.n850 B.n849 585
R1418 B.n17 B.n16 585
R1419 B.n848 B.n17 585
R1420 B.n846 B.n845 585
R1421 B.n847 B.n846 585
R1422 B.n844 B.n22 585
R1423 B.n25 B.n22 585
R1424 B.n843 B.n842 585
R1425 B.n842 B.n841 585
R1426 B.n24 B.n23 585
R1427 B.n840 B.n24 585
R1428 B.n838 B.n837 585
R1429 B.n839 B.n838 585
R1430 B.n836 B.n30 585
R1431 B.n30 B.n29 585
R1432 B.n835 B.n834 585
R1433 B.n834 B.n833 585
R1434 B.n32 B.n31 585
R1435 B.n832 B.n32 585
R1436 B.n830 B.n829 585
R1437 B.n831 B.n830 585
R1438 B.n828 B.n37 585
R1439 B.n37 B.n36 585
R1440 B.n827 B.n826 585
R1441 B.n826 B.n825 585
R1442 B.n867 B.n866 585
R1443 B.n866 B.n865 585
R1444 B.n734 B.n401 564.573
R1445 B.n826 B.n39 564.573
R1446 B.n732 B.n403 564.573
R1447 B.n822 B.n40 564.573
R1448 B.n607 B.t17 405.457
R1449 B.n106 B.t22 405.457
R1450 B.n439 B.t20 405.457
R1451 B.n109 B.t12 405.457
R1452 B.n608 B.t16 392.075
R1453 B.n107 B.t23 392.075
R1454 B.n440 B.t19 392.075
R1455 B.n110 B.t13 392.075
R1456 B.n824 B.n823 256.663
R1457 B.n824 B.n104 256.663
R1458 B.n824 B.n103 256.663
R1459 B.n824 B.n102 256.663
R1460 B.n824 B.n101 256.663
R1461 B.n824 B.n100 256.663
R1462 B.n824 B.n99 256.663
R1463 B.n824 B.n98 256.663
R1464 B.n824 B.n97 256.663
R1465 B.n824 B.n96 256.663
R1466 B.n824 B.n95 256.663
R1467 B.n824 B.n94 256.663
R1468 B.n824 B.n93 256.663
R1469 B.n824 B.n92 256.663
R1470 B.n824 B.n91 256.663
R1471 B.n824 B.n90 256.663
R1472 B.n824 B.n89 256.663
R1473 B.n824 B.n88 256.663
R1474 B.n824 B.n87 256.663
R1475 B.n824 B.n86 256.663
R1476 B.n824 B.n85 256.663
R1477 B.n824 B.n84 256.663
R1478 B.n824 B.n83 256.663
R1479 B.n824 B.n82 256.663
R1480 B.n824 B.n81 256.663
R1481 B.n824 B.n80 256.663
R1482 B.n824 B.n79 256.663
R1483 B.n824 B.n78 256.663
R1484 B.n824 B.n77 256.663
R1485 B.n824 B.n76 256.663
R1486 B.n824 B.n75 256.663
R1487 B.n824 B.n74 256.663
R1488 B.n824 B.n73 256.663
R1489 B.n824 B.n72 256.663
R1490 B.n824 B.n71 256.663
R1491 B.n824 B.n70 256.663
R1492 B.n824 B.n69 256.663
R1493 B.n824 B.n68 256.663
R1494 B.n824 B.n67 256.663
R1495 B.n824 B.n66 256.663
R1496 B.n824 B.n65 256.663
R1497 B.n824 B.n64 256.663
R1498 B.n824 B.n63 256.663
R1499 B.n824 B.n62 256.663
R1500 B.n824 B.n61 256.663
R1501 B.n824 B.n60 256.663
R1502 B.n824 B.n59 256.663
R1503 B.n824 B.n58 256.663
R1504 B.n824 B.n57 256.663
R1505 B.n824 B.n56 256.663
R1506 B.n824 B.n55 256.663
R1507 B.n824 B.n54 256.663
R1508 B.n824 B.n53 256.663
R1509 B.n824 B.n52 256.663
R1510 B.n824 B.n51 256.663
R1511 B.n824 B.n50 256.663
R1512 B.n824 B.n49 256.663
R1513 B.n824 B.n48 256.663
R1514 B.n824 B.n47 256.663
R1515 B.n824 B.n46 256.663
R1516 B.n824 B.n45 256.663
R1517 B.n824 B.n44 256.663
R1518 B.n824 B.n43 256.663
R1519 B.n824 B.n42 256.663
R1520 B.n824 B.n41 256.663
R1521 B.n471 B.n402 256.663
R1522 B.n474 B.n402 256.663
R1523 B.n480 B.n402 256.663
R1524 B.n482 B.n402 256.663
R1525 B.n488 B.n402 256.663
R1526 B.n490 B.n402 256.663
R1527 B.n496 B.n402 256.663
R1528 B.n498 B.n402 256.663
R1529 B.n504 B.n402 256.663
R1530 B.n506 B.n402 256.663
R1531 B.n512 B.n402 256.663
R1532 B.n514 B.n402 256.663
R1533 B.n520 B.n402 256.663
R1534 B.n522 B.n402 256.663
R1535 B.n528 B.n402 256.663
R1536 B.n530 B.n402 256.663
R1537 B.n536 B.n402 256.663
R1538 B.n538 B.n402 256.663
R1539 B.n544 B.n402 256.663
R1540 B.n546 B.n402 256.663
R1541 B.n552 B.n402 256.663
R1542 B.n554 B.n402 256.663
R1543 B.n560 B.n402 256.663
R1544 B.n562 B.n402 256.663
R1545 B.n568 B.n402 256.663
R1546 B.n570 B.n402 256.663
R1547 B.n576 B.n402 256.663
R1548 B.n578 B.n402 256.663
R1549 B.n584 B.n402 256.663
R1550 B.n586 B.n402 256.663
R1551 B.n593 B.n402 256.663
R1552 B.n595 B.n402 256.663
R1553 B.n601 B.n402 256.663
R1554 B.n603 B.n402 256.663
R1555 B.n612 B.n402 256.663
R1556 B.n614 B.n402 256.663
R1557 B.n620 B.n402 256.663
R1558 B.n622 B.n402 256.663
R1559 B.n628 B.n402 256.663
R1560 B.n630 B.n402 256.663
R1561 B.n636 B.n402 256.663
R1562 B.n638 B.n402 256.663
R1563 B.n644 B.n402 256.663
R1564 B.n646 B.n402 256.663
R1565 B.n652 B.n402 256.663
R1566 B.n654 B.n402 256.663
R1567 B.n660 B.n402 256.663
R1568 B.n662 B.n402 256.663
R1569 B.n668 B.n402 256.663
R1570 B.n670 B.n402 256.663
R1571 B.n676 B.n402 256.663
R1572 B.n678 B.n402 256.663
R1573 B.n684 B.n402 256.663
R1574 B.n686 B.n402 256.663
R1575 B.n692 B.n402 256.663
R1576 B.n694 B.n402 256.663
R1577 B.n700 B.n402 256.663
R1578 B.n702 B.n402 256.663
R1579 B.n708 B.n402 256.663
R1580 B.n710 B.n402 256.663
R1581 B.n716 B.n402 256.663
R1582 B.n718 B.n402 256.663
R1583 B.n724 B.n402 256.663
R1584 B.n727 B.n402 256.663
R1585 B.n734 B.n399 163.367
R1586 B.n738 B.n399 163.367
R1587 B.n738 B.n393 163.367
R1588 B.n746 B.n393 163.367
R1589 B.n746 B.n391 163.367
R1590 B.n750 B.n391 163.367
R1591 B.n750 B.n385 163.367
R1592 B.n759 B.n385 163.367
R1593 B.n759 B.n383 163.367
R1594 B.n763 B.n383 163.367
R1595 B.n763 B.n378 163.367
R1596 B.n772 B.n378 163.367
R1597 B.n772 B.n376 163.367
R1598 B.n776 B.n376 163.367
R1599 B.n776 B.n371 163.367
R1600 B.n786 B.n371 163.367
R1601 B.n786 B.n369 163.367
R1602 B.n790 B.n369 163.367
R1603 B.n790 B.n2 163.367
R1604 B.n866 B.n2 163.367
R1605 B.n866 B.n3 163.367
R1606 B.n862 B.n3 163.367
R1607 B.n862 B.n8 163.367
R1608 B.n858 B.n8 163.367
R1609 B.n858 B.n10 163.367
R1610 B.n854 B.n10 163.367
R1611 B.n854 B.n15 163.367
R1612 B.n850 B.n15 163.367
R1613 B.n850 B.n17 163.367
R1614 B.n846 B.n17 163.367
R1615 B.n846 B.n22 163.367
R1616 B.n842 B.n22 163.367
R1617 B.n842 B.n24 163.367
R1618 B.n838 B.n24 163.367
R1619 B.n838 B.n30 163.367
R1620 B.n834 B.n30 163.367
R1621 B.n834 B.n32 163.367
R1622 B.n830 B.n32 163.367
R1623 B.n830 B.n37 163.367
R1624 B.n826 B.n37 163.367
R1625 B.n473 B.n472 163.367
R1626 B.n475 B.n473 163.367
R1627 B.n479 B.n468 163.367
R1628 B.n483 B.n481 163.367
R1629 B.n487 B.n466 163.367
R1630 B.n491 B.n489 163.367
R1631 B.n495 B.n464 163.367
R1632 B.n499 B.n497 163.367
R1633 B.n503 B.n462 163.367
R1634 B.n507 B.n505 163.367
R1635 B.n511 B.n460 163.367
R1636 B.n515 B.n513 163.367
R1637 B.n519 B.n458 163.367
R1638 B.n523 B.n521 163.367
R1639 B.n527 B.n456 163.367
R1640 B.n531 B.n529 163.367
R1641 B.n535 B.n454 163.367
R1642 B.n539 B.n537 163.367
R1643 B.n543 B.n452 163.367
R1644 B.n547 B.n545 163.367
R1645 B.n551 B.n450 163.367
R1646 B.n555 B.n553 163.367
R1647 B.n559 B.n448 163.367
R1648 B.n563 B.n561 163.367
R1649 B.n567 B.n446 163.367
R1650 B.n571 B.n569 163.367
R1651 B.n575 B.n444 163.367
R1652 B.n579 B.n577 163.367
R1653 B.n583 B.n442 163.367
R1654 B.n587 B.n585 163.367
R1655 B.n592 B.n438 163.367
R1656 B.n596 B.n594 163.367
R1657 B.n600 B.n436 163.367
R1658 B.n604 B.n602 163.367
R1659 B.n611 B.n434 163.367
R1660 B.n615 B.n613 163.367
R1661 B.n619 B.n432 163.367
R1662 B.n623 B.n621 163.367
R1663 B.n627 B.n430 163.367
R1664 B.n631 B.n629 163.367
R1665 B.n635 B.n428 163.367
R1666 B.n639 B.n637 163.367
R1667 B.n643 B.n426 163.367
R1668 B.n647 B.n645 163.367
R1669 B.n651 B.n424 163.367
R1670 B.n655 B.n653 163.367
R1671 B.n659 B.n422 163.367
R1672 B.n663 B.n661 163.367
R1673 B.n667 B.n420 163.367
R1674 B.n671 B.n669 163.367
R1675 B.n675 B.n418 163.367
R1676 B.n679 B.n677 163.367
R1677 B.n683 B.n416 163.367
R1678 B.n687 B.n685 163.367
R1679 B.n691 B.n414 163.367
R1680 B.n695 B.n693 163.367
R1681 B.n699 B.n412 163.367
R1682 B.n703 B.n701 163.367
R1683 B.n707 B.n410 163.367
R1684 B.n711 B.n709 163.367
R1685 B.n715 B.n408 163.367
R1686 B.n719 B.n717 163.367
R1687 B.n723 B.n406 163.367
R1688 B.n726 B.n725 163.367
R1689 B.n728 B.n403 163.367
R1690 B.n732 B.n397 163.367
R1691 B.n740 B.n397 163.367
R1692 B.n740 B.n395 163.367
R1693 B.n744 B.n395 163.367
R1694 B.n744 B.n389 163.367
R1695 B.n752 B.n389 163.367
R1696 B.n752 B.n387 163.367
R1697 B.n756 B.n387 163.367
R1698 B.n756 B.n381 163.367
R1699 B.n765 B.n381 163.367
R1700 B.n765 B.n379 163.367
R1701 B.n769 B.n379 163.367
R1702 B.n769 B.n374 163.367
R1703 B.n778 B.n374 163.367
R1704 B.n778 B.n372 163.367
R1705 B.n783 B.n372 163.367
R1706 B.n783 B.n368 163.367
R1707 B.n792 B.n368 163.367
R1708 B.n793 B.n792 163.367
R1709 B.n793 B.n5 163.367
R1710 B.n6 B.n5 163.367
R1711 B.n7 B.n6 163.367
R1712 B.n798 B.n7 163.367
R1713 B.n798 B.n12 163.367
R1714 B.n13 B.n12 163.367
R1715 B.n14 B.n13 163.367
R1716 B.n803 B.n14 163.367
R1717 B.n803 B.n19 163.367
R1718 B.n20 B.n19 163.367
R1719 B.n21 B.n20 163.367
R1720 B.n808 B.n21 163.367
R1721 B.n808 B.n26 163.367
R1722 B.n27 B.n26 163.367
R1723 B.n28 B.n27 163.367
R1724 B.n813 B.n28 163.367
R1725 B.n813 B.n33 163.367
R1726 B.n34 B.n33 163.367
R1727 B.n35 B.n34 163.367
R1728 B.n818 B.n35 163.367
R1729 B.n818 B.n40 163.367
R1730 B.n114 B.n113 163.367
R1731 B.n118 B.n117 163.367
R1732 B.n122 B.n121 163.367
R1733 B.n126 B.n125 163.367
R1734 B.n130 B.n129 163.367
R1735 B.n134 B.n133 163.367
R1736 B.n138 B.n137 163.367
R1737 B.n142 B.n141 163.367
R1738 B.n146 B.n145 163.367
R1739 B.n150 B.n149 163.367
R1740 B.n154 B.n153 163.367
R1741 B.n158 B.n157 163.367
R1742 B.n162 B.n161 163.367
R1743 B.n166 B.n165 163.367
R1744 B.n170 B.n169 163.367
R1745 B.n174 B.n173 163.367
R1746 B.n178 B.n177 163.367
R1747 B.n182 B.n181 163.367
R1748 B.n186 B.n185 163.367
R1749 B.n190 B.n189 163.367
R1750 B.n194 B.n193 163.367
R1751 B.n198 B.n197 163.367
R1752 B.n202 B.n201 163.367
R1753 B.n206 B.n205 163.367
R1754 B.n210 B.n209 163.367
R1755 B.n214 B.n213 163.367
R1756 B.n218 B.n217 163.367
R1757 B.n222 B.n221 163.367
R1758 B.n226 B.n225 163.367
R1759 B.n230 B.n229 163.367
R1760 B.n234 B.n233 163.367
R1761 B.n238 B.n237 163.367
R1762 B.n242 B.n241 163.367
R1763 B.n246 B.n245 163.367
R1764 B.n250 B.n249 163.367
R1765 B.n254 B.n253 163.367
R1766 B.n258 B.n257 163.367
R1767 B.n262 B.n261 163.367
R1768 B.n266 B.n265 163.367
R1769 B.n270 B.n269 163.367
R1770 B.n274 B.n273 163.367
R1771 B.n278 B.n277 163.367
R1772 B.n282 B.n281 163.367
R1773 B.n286 B.n285 163.367
R1774 B.n290 B.n289 163.367
R1775 B.n294 B.n293 163.367
R1776 B.n298 B.n297 163.367
R1777 B.n302 B.n301 163.367
R1778 B.n306 B.n305 163.367
R1779 B.n310 B.n309 163.367
R1780 B.n314 B.n313 163.367
R1781 B.n318 B.n317 163.367
R1782 B.n322 B.n321 163.367
R1783 B.n326 B.n325 163.367
R1784 B.n330 B.n329 163.367
R1785 B.n334 B.n333 163.367
R1786 B.n338 B.n337 163.367
R1787 B.n342 B.n341 163.367
R1788 B.n346 B.n345 163.367
R1789 B.n350 B.n349 163.367
R1790 B.n354 B.n353 163.367
R1791 B.n358 B.n357 163.367
R1792 B.n362 B.n361 163.367
R1793 B.n364 B.n105 163.367
R1794 B.n471 B.n401 71.676
R1795 B.n475 B.n474 71.676
R1796 B.n480 B.n479 71.676
R1797 B.n483 B.n482 71.676
R1798 B.n488 B.n487 71.676
R1799 B.n491 B.n490 71.676
R1800 B.n496 B.n495 71.676
R1801 B.n499 B.n498 71.676
R1802 B.n504 B.n503 71.676
R1803 B.n507 B.n506 71.676
R1804 B.n512 B.n511 71.676
R1805 B.n515 B.n514 71.676
R1806 B.n520 B.n519 71.676
R1807 B.n523 B.n522 71.676
R1808 B.n528 B.n527 71.676
R1809 B.n531 B.n530 71.676
R1810 B.n536 B.n535 71.676
R1811 B.n539 B.n538 71.676
R1812 B.n544 B.n543 71.676
R1813 B.n547 B.n546 71.676
R1814 B.n552 B.n551 71.676
R1815 B.n555 B.n554 71.676
R1816 B.n560 B.n559 71.676
R1817 B.n563 B.n562 71.676
R1818 B.n568 B.n567 71.676
R1819 B.n571 B.n570 71.676
R1820 B.n576 B.n575 71.676
R1821 B.n579 B.n578 71.676
R1822 B.n584 B.n583 71.676
R1823 B.n587 B.n586 71.676
R1824 B.n593 B.n592 71.676
R1825 B.n596 B.n595 71.676
R1826 B.n601 B.n600 71.676
R1827 B.n604 B.n603 71.676
R1828 B.n612 B.n611 71.676
R1829 B.n615 B.n614 71.676
R1830 B.n620 B.n619 71.676
R1831 B.n623 B.n622 71.676
R1832 B.n628 B.n627 71.676
R1833 B.n631 B.n630 71.676
R1834 B.n636 B.n635 71.676
R1835 B.n639 B.n638 71.676
R1836 B.n644 B.n643 71.676
R1837 B.n647 B.n646 71.676
R1838 B.n652 B.n651 71.676
R1839 B.n655 B.n654 71.676
R1840 B.n660 B.n659 71.676
R1841 B.n663 B.n662 71.676
R1842 B.n668 B.n667 71.676
R1843 B.n671 B.n670 71.676
R1844 B.n676 B.n675 71.676
R1845 B.n679 B.n678 71.676
R1846 B.n684 B.n683 71.676
R1847 B.n687 B.n686 71.676
R1848 B.n692 B.n691 71.676
R1849 B.n695 B.n694 71.676
R1850 B.n700 B.n699 71.676
R1851 B.n703 B.n702 71.676
R1852 B.n708 B.n707 71.676
R1853 B.n711 B.n710 71.676
R1854 B.n716 B.n715 71.676
R1855 B.n719 B.n718 71.676
R1856 B.n724 B.n723 71.676
R1857 B.n727 B.n726 71.676
R1858 B.n41 B.n39 71.676
R1859 B.n114 B.n42 71.676
R1860 B.n118 B.n43 71.676
R1861 B.n122 B.n44 71.676
R1862 B.n126 B.n45 71.676
R1863 B.n130 B.n46 71.676
R1864 B.n134 B.n47 71.676
R1865 B.n138 B.n48 71.676
R1866 B.n142 B.n49 71.676
R1867 B.n146 B.n50 71.676
R1868 B.n150 B.n51 71.676
R1869 B.n154 B.n52 71.676
R1870 B.n158 B.n53 71.676
R1871 B.n162 B.n54 71.676
R1872 B.n166 B.n55 71.676
R1873 B.n170 B.n56 71.676
R1874 B.n174 B.n57 71.676
R1875 B.n178 B.n58 71.676
R1876 B.n182 B.n59 71.676
R1877 B.n186 B.n60 71.676
R1878 B.n190 B.n61 71.676
R1879 B.n194 B.n62 71.676
R1880 B.n198 B.n63 71.676
R1881 B.n202 B.n64 71.676
R1882 B.n206 B.n65 71.676
R1883 B.n210 B.n66 71.676
R1884 B.n214 B.n67 71.676
R1885 B.n218 B.n68 71.676
R1886 B.n222 B.n69 71.676
R1887 B.n226 B.n70 71.676
R1888 B.n230 B.n71 71.676
R1889 B.n234 B.n72 71.676
R1890 B.n238 B.n73 71.676
R1891 B.n242 B.n74 71.676
R1892 B.n246 B.n75 71.676
R1893 B.n250 B.n76 71.676
R1894 B.n254 B.n77 71.676
R1895 B.n258 B.n78 71.676
R1896 B.n262 B.n79 71.676
R1897 B.n266 B.n80 71.676
R1898 B.n270 B.n81 71.676
R1899 B.n274 B.n82 71.676
R1900 B.n278 B.n83 71.676
R1901 B.n282 B.n84 71.676
R1902 B.n286 B.n85 71.676
R1903 B.n290 B.n86 71.676
R1904 B.n294 B.n87 71.676
R1905 B.n298 B.n88 71.676
R1906 B.n302 B.n89 71.676
R1907 B.n306 B.n90 71.676
R1908 B.n310 B.n91 71.676
R1909 B.n314 B.n92 71.676
R1910 B.n318 B.n93 71.676
R1911 B.n322 B.n94 71.676
R1912 B.n326 B.n95 71.676
R1913 B.n330 B.n96 71.676
R1914 B.n334 B.n97 71.676
R1915 B.n338 B.n98 71.676
R1916 B.n342 B.n99 71.676
R1917 B.n346 B.n100 71.676
R1918 B.n350 B.n101 71.676
R1919 B.n354 B.n102 71.676
R1920 B.n358 B.n103 71.676
R1921 B.n362 B.n104 71.676
R1922 B.n823 B.n105 71.676
R1923 B.n823 B.n822 71.676
R1924 B.n364 B.n104 71.676
R1925 B.n361 B.n103 71.676
R1926 B.n357 B.n102 71.676
R1927 B.n353 B.n101 71.676
R1928 B.n349 B.n100 71.676
R1929 B.n345 B.n99 71.676
R1930 B.n341 B.n98 71.676
R1931 B.n337 B.n97 71.676
R1932 B.n333 B.n96 71.676
R1933 B.n329 B.n95 71.676
R1934 B.n325 B.n94 71.676
R1935 B.n321 B.n93 71.676
R1936 B.n317 B.n92 71.676
R1937 B.n313 B.n91 71.676
R1938 B.n309 B.n90 71.676
R1939 B.n305 B.n89 71.676
R1940 B.n301 B.n88 71.676
R1941 B.n297 B.n87 71.676
R1942 B.n293 B.n86 71.676
R1943 B.n289 B.n85 71.676
R1944 B.n285 B.n84 71.676
R1945 B.n281 B.n83 71.676
R1946 B.n277 B.n82 71.676
R1947 B.n273 B.n81 71.676
R1948 B.n269 B.n80 71.676
R1949 B.n265 B.n79 71.676
R1950 B.n261 B.n78 71.676
R1951 B.n257 B.n77 71.676
R1952 B.n253 B.n76 71.676
R1953 B.n249 B.n75 71.676
R1954 B.n245 B.n74 71.676
R1955 B.n241 B.n73 71.676
R1956 B.n237 B.n72 71.676
R1957 B.n233 B.n71 71.676
R1958 B.n229 B.n70 71.676
R1959 B.n225 B.n69 71.676
R1960 B.n221 B.n68 71.676
R1961 B.n217 B.n67 71.676
R1962 B.n213 B.n66 71.676
R1963 B.n209 B.n65 71.676
R1964 B.n205 B.n64 71.676
R1965 B.n201 B.n63 71.676
R1966 B.n197 B.n62 71.676
R1967 B.n193 B.n61 71.676
R1968 B.n189 B.n60 71.676
R1969 B.n185 B.n59 71.676
R1970 B.n181 B.n58 71.676
R1971 B.n177 B.n57 71.676
R1972 B.n173 B.n56 71.676
R1973 B.n169 B.n55 71.676
R1974 B.n165 B.n54 71.676
R1975 B.n161 B.n53 71.676
R1976 B.n157 B.n52 71.676
R1977 B.n153 B.n51 71.676
R1978 B.n149 B.n50 71.676
R1979 B.n145 B.n49 71.676
R1980 B.n141 B.n48 71.676
R1981 B.n137 B.n47 71.676
R1982 B.n133 B.n46 71.676
R1983 B.n129 B.n45 71.676
R1984 B.n125 B.n44 71.676
R1985 B.n121 B.n43 71.676
R1986 B.n117 B.n42 71.676
R1987 B.n113 B.n41 71.676
R1988 B.n472 B.n471 71.676
R1989 B.n474 B.n468 71.676
R1990 B.n481 B.n480 71.676
R1991 B.n482 B.n466 71.676
R1992 B.n489 B.n488 71.676
R1993 B.n490 B.n464 71.676
R1994 B.n497 B.n496 71.676
R1995 B.n498 B.n462 71.676
R1996 B.n505 B.n504 71.676
R1997 B.n506 B.n460 71.676
R1998 B.n513 B.n512 71.676
R1999 B.n514 B.n458 71.676
R2000 B.n521 B.n520 71.676
R2001 B.n522 B.n456 71.676
R2002 B.n529 B.n528 71.676
R2003 B.n530 B.n454 71.676
R2004 B.n537 B.n536 71.676
R2005 B.n538 B.n452 71.676
R2006 B.n545 B.n544 71.676
R2007 B.n546 B.n450 71.676
R2008 B.n553 B.n552 71.676
R2009 B.n554 B.n448 71.676
R2010 B.n561 B.n560 71.676
R2011 B.n562 B.n446 71.676
R2012 B.n569 B.n568 71.676
R2013 B.n570 B.n444 71.676
R2014 B.n577 B.n576 71.676
R2015 B.n578 B.n442 71.676
R2016 B.n585 B.n584 71.676
R2017 B.n586 B.n438 71.676
R2018 B.n594 B.n593 71.676
R2019 B.n595 B.n436 71.676
R2020 B.n602 B.n601 71.676
R2021 B.n603 B.n434 71.676
R2022 B.n613 B.n612 71.676
R2023 B.n614 B.n432 71.676
R2024 B.n621 B.n620 71.676
R2025 B.n622 B.n430 71.676
R2026 B.n629 B.n628 71.676
R2027 B.n630 B.n428 71.676
R2028 B.n637 B.n636 71.676
R2029 B.n638 B.n426 71.676
R2030 B.n645 B.n644 71.676
R2031 B.n646 B.n424 71.676
R2032 B.n653 B.n652 71.676
R2033 B.n654 B.n422 71.676
R2034 B.n661 B.n660 71.676
R2035 B.n662 B.n420 71.676
R2036 B.n669 B.n668 71.676
R2037 B.n670 B.n418 71.676
R2038 B.n677 B.n676 71.676
R2039 B.n678 B.n416 71.676
R2040 B.n685 B.n684 71.676
R2041 B.n686 B.n414 71.676
R2042 B.n693 B.n692 71.676
R2043 B.n694 B.n412 71.676
R2044 B.n701 B.n700 71.676
R2045 B.n702 B.n410 71.676
R2046 B.n709 B.n708 71.676
R2047 B.n710 B.n408 71.676
R2048 B.n717 B.n716 71.676
R2049 B.n718 B.n406 71.676
R2050 B.n725 B.n724 71.676
R2051 B.n728 B.n727 71.676
R2052 B.n733 B.n402 66.5543
R2053 B.n825 B.n824 66.5543
R2054 B.n609 B.n608 59.5399
R2055 B.n589 B.n440 59.5399
R2056 B.n111 B.n110 59.5399
R2057 B.n108 B.n107 59.5399
R2058 B.n821 B.n820 36.6834
R2059 B.n827 B.n38 36.6834
R2060 B.n731 B.n730 36.6834
R2061 B.n735 B.n400 36.6834
R2062 B.n733 B.n398 31.6485
R2063 B.n739 B.n398 31.6485
R2064 B.n739 B.n394 31.6485
R2065 B.n745 B.n394 31.6485
R2066 B.n751 B.n390 31.6485
R2067 B.n751 B.n386 31.6485
R2068 B.n758 B.n386 31.6485
R2069 B.n758 B.n757 31.6485
R2070 B.n764 B.n382 31.6485
R2071 B.n771 B.n770 31.6485
R2072 B.n777 B.n375 31.6485
R2073 B.n785 B.n784 31.6485
R2074 B.n791 B.n4 31.6485
R2075 B.n865 B.n4 31.6485
R2076 B.n865 B.n864 31.6485
R2077 B.n864 B.n863 31.6485
R2078 B.n857 B.n11 31.6485
R2079 B.n856 B.n855 31.6485
R2080 B.n849 B.n18 31.6485
R2081 B.n848 B.n847 31.6485
R2082 B.n841 B.n25 31.6485
R2083 B.n841 B.n840 31.6485
R2084 B.n840 B.n839 31.6485
R2085 B.n839 B.n29 31.6485
R2086 B.n833 B.n832 31.6485
R2087 B.n832 B.n831 31.6485
R2088 B.n831 B.n36 31.6485
R2089 B.n825 B.n36 31.6485
R2090 B.t15 B.n390 30.7177
R2091 B.t11 B.n29 30.7177
R2092 B.n764 B.t5 23.2711
R2093 B.n847 B.t6 23.2711
R2094 B.n771 B.t7 22.3403
R2095 B.n849 B.t0 22.3403
R2096 B.n777 B.t3 21.4094
R2097 B.n855 B.t1 21.4094
R2098 B.n785 B.t2 20.4786
R2099 B.n857 B.t4 20.4786
R2100 B.n791 B.t8 19.5478
R2101 B.n863 B.t9 19.5478
R2102 B B.n867 18.0485
R2103 B.n608 B.n607 13.3823
R2104 B.n440 B.n439 13.3823
R2105 B.n110 B.n109 13.3823
R2106 B.n107 B.n106 13.3823
R2107 B.n784 B.t8 12.1012
R2108 B.n11 B.t9 12.1012
R2109 B.n375 B.t2 11.1704
R2110 B.t4 B.n856 11.1704
R2111 B.n112 B.n38 10.6151
R2112 B.n115 B.n112 10.6151
R2113 B.n116 B.n115 10.6151
R2114 B.n119 B.n116 10.6151
R2115 B.n120 B.n119 10.6151
R2116 B.n123 B.n120 10.6151
R2117 B.n124 B.n123 10.6151
R2118 B.n127 B.n124 10.6151
R2119 B.n128 B.n127 10.6151
R2120 B.n131 B.n128 10.6151
R2121 B.n132 B.n131 10.6151
R2122 B.n135 B.n132 10.6151
R2123 B.n136 B.n135 10.6151
R2124 B.n139 B.n136 10.6151
R2125 B.n140 B.n139 10.6151
R2126 B.n143 B.n140 10.6151
R2127 B.n144 B.n143 10.6151
R2128 B.n147 B.n144 10.6151
R2129 B.n148 B.n147 10.6151
R2130 B.n151 B.n148 10.6151
R2131 B.n152 B.n151 10.6151
R2132 B.n155 B.n152 10.6151
R2133 B.n156 B.n155 10.6151
R2134 B.n159 B.n156 10.6151
R2135 B.n160 B.n159 10.6151
R2136 B.n163 B.n160 10.6151
R2137 B.n164 B.n163 10.6151
R2138 B.n167 B.n164 10.6151
R2139 B.n168 B.n167 10.6151
R2140 B.n171 B.n168 10.6151
R2141 B.n172 B.n171 10.6151
R2142 B.n175 B.n172 10.6151
R2143 B.n176 B.n175 10.6151
R2144 B.n179 B.n176 10.6151
R2145 B.n180 B.n179 10.6151
R2146 B.n183 B.n180 10.6151
R2147 B.n184 B.n183 10.6151
R2148 B.n187 B.n184 10.6151
R2149 B.n188 B.n187 10.6151
R2150 B.n191 B.n188 10.6151
R2151 B.n192 B.n191 10.6151
R2152 B.n195 B.n192 10.6151
R2153 B.n196 B.n195 10.6151
R2154 B.n199 B.n196 10.6151
R2155 B.n200 B.n199 10.6151
R2156 B.n203 B.n200 10.6151
R2157 B.n204 B.n203 10.6151
R2158 B.n207 B.n204 10.6151
R2159 B.n208 B.n207 10.6151
R2160 B.n211 B.n208 10.6151
R2161 B.n212 B.n211 10.6151
R2162 B.n215 B.n212 10.6151
R2163 B.n216 B.n215 10.6151
R2164 B.n219 B.n216 10.6151
R2165 B.n220 B.n219 10.6151
R2166 B.n223 B.n220 10.6151
R2167 B.n224 B.n223 10.6151
R2168 B.n227 B.n224 10.6151
R2169 B.n228 B.n227 10.6151
R2170 B.n232 B.n231 10.6151
R2171 B.n235 B.n232 10.6151
R2172 B.n236 B.n235 10.6151
R2173 B.n239 B.n236 10.6151
R2174 B.n240 B.n239 10.6151
R2175 B.n243 B.n240 10.6151
R2176 B.n244 B.n243 10.6151
R2177 B.n247 B.n244 10.6151
R2178 B.n248 B.n247 10.6151
R2179 B.n252 B.n251 10.6151
R2180 B.n255 B.n252 10.6151
R2181 B.n256 B.n255 10.6151
R2182 B.n259 B.n256 10.6151
R2183 B.n260 B.n259 10.6151
R2184 B.n263 B.n260 10.6151
R2185 B.n264 B.n263 10.6151
R2186 B.n267 B.n264 10.6151
R2187 B.n268 B.n267 10.6151
R2188 B.n271 B.n268 10.6151
R2189 B.n272 B.n271 10.6151
R2190 B.n275 B.n272 10.6151
R2191 B.n276 B.n275 10.6151
R2192 B.n279 B.n276 10.6151
R2193 B.n280 B.n279 10.6151
R2194 B.n283 B.n280 10.6151
R2195 B.n284 B.n283 10.6151
R2196 B.n287 B.n284 10.6151
R2197 B.n288 B.n287 10.6151
R2198 B.n291 B.n288 10.6151
R2199 B.n292 B.n291 10.6151
R2200 B.n295 B.n292 10.6151
R2201 B.n296 B.n295 10.6151
R2202 B.n299 B.n296 10.6151
R2203 B.n300 B.n299 10.6151
R2204 B.n303 B.n300 10.6151
R2205 B.n304 B.n303 10.6151
R2206 B.n307 B.n304 10.6151
R2207 B.n308 B.n307 10.6151
R2208 B.n311 B.n308 10.6151
R2209 B.n312 B.n311 10.6151
R2210 B.n315 B.n312 10.6151
R2211 B.n316 B.n315 10.6151
R2212 B.n319 B.n316 10.6151
R2213 B.n320 B.n319 10.6151
R2214 B.n323 B.n320 10.6151
R2215 B.n324 B.n323 10.6151
R2216 B.n327 B.n324 10.6151
R2217 B.n328 B.n327 10.6151
R2218 B.n331 B.n328 10.6151
R2219 B.n332 B.n331 10.6151
R2220 B.n335 B.n332 10.6151
R2221 B.n336 B.n335 10.6151
R2222 B.n339 B.n336 10.6151
R2223 B.n340 B.n339 10.6151
R2224 B.n343 B.n340 10.6151
R2225 B.n344 B.n343 10.6151
R2226 B.n347 B.n344 10.6151
R2227 B.n348 B.n347 10.6151
R2228 B.n351 B.n348 10.6151
R2229 B.n352 B.n351 10.6151
R2230 B.n355 B.n352 10.6151
R2231 B.n356 B.n355 10.6151
R2232 B.n359 B.n356 10.6151
R2233 B.n360 B.n359 10.6151
R2234 B.n363 B.n360 10.6151
R2235 B.n365 B.n363 10.6151
R2236 B.n366 B.n365 10.6151
R2237 B.n821 B.n366 10.6151
R2238 B.n731 B.n396 10.6151
R2239 B.n741 B.n396 10.6151
R2240 B.n742 B.n741 10.6151
R2241 B.n743 B.n742 10.6151
R2242 B.n743 B.n388 10.6151
R2243 B.n753 B.n388 10.6151
R2244 B.n754 B.n753 10.6151
R2245 B.n755 B.n754 10.6151
R2246 B.n755 B.n380 10.6151
R2247 B.n766 B.n380 10.6151
R2248 B.n767 B.n766 10.6151
R2249 B.n768 B.n767 10.6151
R2250 B.n768 B.n373 10.6151
R2251 B.n779 B.n373 10.6151
R2252 B.n780 B.n779 10.6151
R2253 B.n782 B.n780 10.6151
R2254 B.n782 B.n781 10.6151
R2255 B.n781 B.n367 10.6151
R2256 B.n794 B.n367 10.6151
R2257 B.n795 B.n794 10.6151
R2258 B.n796 B.n795 10.6151
R2259 B.n797 B.n796 10.6151
R2260 B.n799 B.n797 10.6151
R2261 B.n800 B.n799 10.6151
R2262 B.n801 B.n800 10.6151
R2263 B.n802 B.n801 10.6151
R2264 B.n804 B.n802 10.6151
R2265 B.n805 B.n804 10.6151
R2266 B.n806 B.n805 10.6151
R2267 B.n807 B.n806 10.6151
R2268 B.n809 B.n807 10.6151
R2269 B.n810 B.n809 10.6151
R2270 B.n811 B.n810 10.6151
R2271 B.n812 B.n811 10.6151
R2272 B.n814 B.n812 10.6151
R2273 B.n815 B.n814 10.6151
R2274 B.n816 B.n815 10.6151
R2275 B.n817 B.n816 10.6151
R2276 B.n819 B.n817 10.6151
R2277 B.n820 B.n819 10.6151
R2278 B.n470 B.n400 10.6151
R2279 B.n470 B.n469 10.6151
R2280 B.n476 B.n469 10.6151
R2281 B.n477 B.n476 10.6151
R2282 B.n478 B.n477 10.6151
R2283 B.n478 B.n467 10.6151
R2284 B.n484 B.n467 10.6151
R2285 B.n485 B.n484 10.6151
R2286 B.n486 B.n485 10.6151
R2287 B.n486 B.n465 10.6151
R2288 B.n492 B.n465 10.6151
R2289 B.n493 B.n492 10.6151
R2290 B.n494 B.n493 10.6151
R2291 B.n494 B.n463 10.6151
R2292 B.n500 B.n463 10.6151
R2293 B.n501 B.n500 10.6151
R2294 B.n502 B.n501 10.6151
R2295 B.n502 B.n461 10.6151
R2296 B.n508 B.n461 10.6151
R2297 B.n509 B.n508 10.6151
R2298 B.n510 B.n509 10.6151
R2299 B.n510 B.n459 10.6151
R2300 B.n516 B.n459 10.6151
R2301 B.n517 B.n516 10.6151
R2302 B.n518 B.n517 10.6151
R2303 B.n518 B.n457 10.6151
R2304 B.n524 B.n457 10.6151
R2305 B.n525 B.n524 10.6151
R2306 B.n526 B.n525 10.6151
R2307 B.n526 B.n455 10.6151
R2308 B.n532 B.n455 10.6151
R2309 B.n533 B.n532 10.6151
R2310 B.n534 B.n533 10.6151
R2311 B.n534 B.n453 10.6151
R2312 B.n540 B.n453 10.6151
R2313 B.n541 B.n540 10.6151
R2314 B.n542 B.n541 10.6151
R2315 B.n542 B.n451 10.6151
R2316 B.n548 B.n451 10.6151
R2317 B.n549 B.n548 10.6151
R2318 B.n550 B.n549 10.6151
R2319 B.n550 B.n449 10.6151
R2320 B.n556 B.n449 10.6151
R2321 B.n557 B.n556 10.6151
R2322 B.n558 B.n557 10.6151
R2323 B.n558 B.n447 10.6151
R2324 B.n564 B.n447 10.6151
R2325 B.n565 B.n564 10.6151
R2326 B.n566 B.n565 10.6151
R2327 B.n566 B.n445 10.6151
R2328 B.n572 B.n445 10.6151
R2329 B.n573 B.n572 10.6151
R2330 B.n574 B.n573 10.6151
R2331 B.n574 B.n443 10.6151
R2332 B.n580 B.n443 10.6151
R2333 B.n581 B.n580 10.6151
R2334 B.n582 B.n581 10.6151
R2335 B.n582 B.n441 10.6151
R2336 B.n588 B.n441 10.6151
R2337 B.n591 B.n590 10.6151
R2338 B.n591 B.n437 10.6151
R2339 B.n597 B.n437 10.6151
R2340 B.n598 B.n597 10.6151
R2341 B.n599 B.n598 10.6151
R2342 B.n599 B.n435 10.6151
R2343 B.n605 B.n435 10.6151
R2344 B.n606 B.n605 10.6151
R2345 B.n610 B.n606 10.6151
R2346 B.n616 B.n433 10.6151
R2347 B.n617 B.n616 10.6151
R2348 B.n618 B.n617 10.6151
R2349 B.n618 B.n431 10.6151
R2350 B.n624 B.n431 10.6151
R2351 B.n625 B.n624 10.6151
R2352 B.n626 B.n625 10.6151
R2353 B.n626 B.n429 10.6151
R2354 B.n632 B.n429 10.6151
R2355 B.n633 B.n632 10.6151
R2356 B.n634 B.n633 10.6151
R2357 B.n634 B.n427 10.6151
R2358 B.n640 B.n427 10.6151
R2359 B.n641 B.n640 10.6151
R2360 B.n642 B.n641 10.6151
R2361 B.n642 B.n425 10.6151
R2362 B.n648 B.n425 10.6151
R2363 B.n649 B.n648 10.6151
R2364 B.n650 B.n649 10.6151
R2365 B.n650 B.n423 10.6151
R2366 B.n656 B.n423 10.6151
R2367 B.n657 B.n656 10.6151
R2368 B.n658 B.n657 10.6151
R2369 B.n658 B.n421 10.6151
R2370 B.n664 B.n421 10.6151
R2371 B.n665 B.n664 10.6151
R2372 B.n666 B.n665 10.6151
R2373 B.n666 B.n419 10.6151
R2374 B.n672 B.n419 10.6151
R2375 B.n673 B.n672 10.6151
R2376 B.n674 B.n673 10.6151
R2377 B.n674 B.n417 10.6151
R2378 B.n680 B.n417 10.6151
R2379 B.n681 B.n680 10.6151
R2380 B.n682 B.n681 10.6151
R2381 B.n682 B.n415 10.6151
R2382 B.n688 B.n415 10.6151
R2383 B.n689 B.n688 10.6151
R2384 B.n690 B.n689 10.6151
R2385 B.n690 B.n413 10.6151
R2386 B.n696 B.n413 10.6151
R2387 B.n697 B.n696 10.6151
R2388 B.n698 B.n697 10.6151
R2389 B.n698 B.n411 10.6151
R2390 B.n704 B.n411 10.6151
R2391 B.n705 B.n704 10.6151
R2392 B.n706 B.n705 10.6151
R2393 B.n706 B.n409 10.6151
R2394 B.n712 B.n409 10.6151
R2395 B.n713 B.n712 10.6151
R2396 B.n714 B.n713 10.6151
R2397 B.n714 B.n407 10.6151
R2398 B.n720 B.n407 10.6151
R2399 B.n721 B.n720 10.6151
R2400 B.n722 B.n721 10.6151
R2401 B.n722 B.n405 10.6151
R2402 B.n405 B.n404 10.6151
R2403 B.n729 B.n404 10.6151
R2404 B.n730 B.n729 10.6151
R2405 B.n736 B.n735 10.6151
R2406 B.n737 B.n736 10.6151
R2407 B.n737 B.n392 10.6151
R2408 B.n747 B.n392 10.6151
R2409 B.n748 B.n747 10.6151
R2410 B.n749 B.n748 10.6151
R2411 B.n749 B.n384 10.6151
R2412 B.n760 B.n384 10.6151
R2413 B.n761 B.n760 10.6151
R2414 B.n762 B.n761 10.6151
R2415 B.n762 B.n377 10.6151
R2416 B.n773 B.n377 10.6151
R2417 B.n774 B.n773 10.6151
R2418 B.n775 B.n774 10.6151
R2419 B.n775 B.n370 10.6151
R2420 B.n787 B.n370 10.6151
R2421 B.n788 B.n787 10.6151
R2422 B.n789 B.n788 10.6151
R2423 B.n789 B.n0 10.6151
R2424 B.n861 B.n1 10.6151
R2425 B.n861 B.n860 10.6151
R2426 B.n860 B.n859 10.6151
R2427 B.n859 B.n9 10.6151
R2428 B.n853 B.n9 10.6151
R2429 B.n853 B.n852 10.6151
R2430 B.n852 B.n851 10.6151
R2431 B.n851 B.n16 10.6151
R2432 B.n845 B.n16 10.6151
R2433 B.n845 B.n844 10.6151
R2434 B.n844 B.n843 10.6151
R2435 B.n843 B.n23 10.6151
R2436 B.n837 B.n23 10.6151
R2437 B.n837 B.n836 10.6151
R2438 B.n836 B.n835 10.6151
R2439 B.n835 B.n31 10.6151
R2440 B.n829 B.n31 10.6151
R2441 B.n829 B.n828 10.6151
R2442 B.n828 B.n827 10.6151
R2443 B.n770 B.t3 10.2396
R2444 B.n18 B.t1 10.2396
R2445 B.n228 B.n111 9.36635
R2446 B.n251 B.n108 9.36635
R2447 B.n589 B.n588 9.36635
R2448 B.n609 B.n433 9.36635
R2449 B.n382 B.t7 9.30873
R2450 B.t0 B.n848 9.30873
R2451 B.n757 B.t5 8.37791
R2452 B.n25 B.t6 8.37791
R2453 B.n867 B.n0 2.81026
R2454 B.n867 B.n1 2.81026
R2455 B.n231 B.n111 1.24928
R2456 B.n248 B.n108 1.24928
R2457 B.n590 B.n589 1.24928
R2458 B.n610 B.n609 1.24928
R2459 B.n745 B.t15 0.931323
R2460 B.n833 B.t11 0.931323
R2461 VN.n2 VN.t8 1359.2
R2462 VN.n13 VN.t6 1359.2
R2463 VN.n3 VN.t3 1338.22
R2464 VN.n1 VN.t2 1338.22
R2465 VN.n8 VN.t0 1338.22
R2466 VN.n9 VN.t5 1338.22
R2467 VN.n14 VN.t9 1338.22
R2468 VN.n12 VN.t4 1338.22
R2469 VN.n19 VN.t7 1338.22
R2470 VN.n20 VN.t1 1338.22
R2471 VN.n10 VN.n9 161.3
R2472 VN.n21 VN.n20 161.3
R2473 VN.n19 VN.n11 161.3
R2474 VN.n18 VN.n17 161.3
R2475 VN.n16 VN.n15 161.3
R2476 VN.n8 VN.n0 161.3
R2477 VN.n7 VN.n6 161.3
R2478 VN.n5 VN.n4 161.3
R2479 VN.n16 VN.n13 70.4033
R2480 VN.n5 VN.n2 70.4033
R2481 VN.n9 VN.n8 48.2005
R2482 VN.n20 VN.n19 48.2005
R2483 VN VN.n21 46.1047
R2484 VN.n4 VN.n3 37.9763
R2485 VN.n8 VN.n7 37.9763
R2486 VN.n15 VN.n14 37.9763
R2487 VN.n19 VN.n18 37.9763
R2488 VN.n14 VN.n13 20.9576
R2489 VN.n3 VN.n2 20.9576
R2490 VN.n4 VN.n1 10.2247
R2491 VN.n7 VN.n1 10.2247
R2492 VN.n15 VN.n12 10.2247
R2493 VN.n18 VN.n12 10.2247
R2494 VN.n21 VN.n11 0.189894
R2495 VN.n17 VN.n11 0.189894
R2496 VN.n17 VN.n16 0.189894
R2497 VN.n6 VN.n5 0.189894
R2498 VN.n6 VN.n0 0.189894
R2499 VN.n10 VN.n0 0.189894
R2500 VN VN.n10 0.0516364
R2501 VDD2.n201 VDD2.n105 289.615
R2502 VDD2.n96 VDD2.n0 289.615
R2503 VDD2.n202 VDD2.n201 185
R2504 VDD2.n200 VDD2.n199 185
R2505 VDD2.n109 VDD2.n108 185
R2506 VDD2.n194 VDD2.n193 185
R2507 VDD2.n192 VDD2.n191 185
R2508 VDD2.n113 VDD2.n112 185
R2509 VDD2.n186 VDD2.n185 185
R2510 VDD2.n184 VDD2.n115 185
R2511 VDD2.n183 VDD2.n182 185
R2512 VDD2.n118 VDD2.n116 185
R2513 VDD2.n177 VDD2.n176 185
R2514 VDD2.n175 VDD2.n174 185
R2515 VDD2.n122 VDD2.n121 185
R2516 VDD2.n169 VDD2.n168 185
R2517 VDD2.n167 VDD2.n166 185
R2518 VDD2.n126 VDD2.n125 185
R2519 VDD2.n161 VDD2.n160 185
R2520 VDD2.n159 VDD2.n158 185
R2521 VDD2.n130 VDD2.n129 185
R2522 VDD2.n153 VDD2.n152 185
R2523 VDD2.n151 VDD2.n150 185
R2524 VDD2.n134 VDD2.n133 185
R2525 VDD2.n145 VDD2.n144 185
R2526 VDD2.n143 VDD2.n142 185
R2527 VDD2.n138 VDD2.n137 185
R2528 VDD2.n32 VDD2.n31 185
R2529 VDD2.n37 VDD2.n36 185
R2530 VDD2.n39 VDD2.n38 185
R2531 VDD2.n28 VDD2.n27 185
R2532 VDD2.n45 VDD2.n44 185
R2533 VDD2.n47 VDD2.n46 185
R2534 VDD2.n24 VDD2.n23 185
R2535 VDD2.n53 VDD2.n52 185
R2536 VDD2.n55 VDD2.n54 185
R2537 VDD2.n20 VDD2.n19 185
R2538 VDD2.n61 VDD2.n60 185
R2539 VDD2.n63 VDD2.n62 185
R2540 VDD2.n16 VDD2.n15 185
R2541 VDD2.n69 VDD2.n68 185
R2542 VDD2.n71 VDD2.n70 185
R2543 VDD2.n12 VDD2.n11 185
R2544 VDD2.n78 VDD2.n77 185
R2545 VDD2.n79 VDD2.n10 185
R2546 VDD2.n81 VDD2.n80 185
R2547 VDD2.n8 VDD2.n7 185
R2548 VDD2.n87 VDD2.n86 185
R2549 VDD2.n89 VDD2.n88 185
R2550 VDD2.n4 VDD2.n3 185
R2551 VDD2.n95 VDD2.n94 185
R2552 VDD2.n97 VDD2.n96 185
R2553 VDD2.n139 VDD2.t8 147.659
R2554 VDD2.n33 VDD2.t1 147.659
R2555 VDD2.n201 VDD2.n200 104.615
R2556 VDD2.n200 VDD2.n108 104.615
R2557 VDD2.n193 VDD2.n108 104.615
R2558 VDD2.n193 VDD2.n192 104.615
R2559 VDD2.n192 VDD2.n112 104.615
R2560 VDD2.n185 VDD2.n112 104.615
R2561 VDD2.n185 VDD2.n184 104.615
R2562 VDD2.n184 VDD2.n183 104.615
R2563 VDD2.n183 VDD2.n116 104.615
R2564 VDD2.n176 VDD2.n116 104.615
R2565 VDD2.n176 VDD2.n175 104.615
R2566 VDD2.n175 VDD2.n121 104.615
R2567 VDD2.n168 VDD2.n121 104.615
R2568 VDD2.n168 VDD2.n167 104.615
R2569 VDD2.n167 VDD2.n125 104.615
R2570 VDD2.n160 VDD2.n125 104.615
R2571 VDD2.n160 VDD2.n159 104.615
R2572 VDD2.n159 VDD2.n129 104.615
R2573 VDD2.n152 VDD2.n129 104.615
R2574 VDD2.n152 VDD2.n151 104.615
R2575 VDD2.n151 VDD2.n133 104.615
R2576 VDD2.n144 VDD2.n133 104.615
R2577 VDD2.n144 VDD2.n143 104.615
R2578 VDD2.n143 VDD2.n137 104.615
R2579 VDD2.n37 VDD2.n31 104.615
R2580 VDD2.n38 VDD2.n37 104.615
R2581 VDD2.n38 VDD2.n27 104.615
R2582 VDD2.n45 VDD2.n27 104.615
R2583 VDD2.n46 VDD2.n45 104.615
R2584 VDD2.n46 VDD2.n23 104.615
R2585 VDD2.n53 VDD2.n23 104.615
R2586 VDD2.n54 VDD2.n53 104.615
R2587 VDD2.n54 VDD2.n19 104.615
R2588 VDD2.n61 VDD2.n19 104.615
R2589 VDD2.n62 VDD2.n61 104.615
R2590 VDD2.n62 VDD2.n15 104.615
R2591 VDD2.n69 VDD2.n15 104.615
R2592 VDD2.n70 VDD2.n69 104.615
R2593 VDD2.n70 VDD2.n11 104.615
R2594 VDD2.n78 VDD2.n11 104.615
R2595 VDD2.n79 VDD2.n78 104.615
R2596 VDD2.n80 VDD2.n79 104.615
R2597 VDD2.n80 VDD2.n7 104.615
R2598 VDD2.n87 VDD2.n7 104.615
R2599 VDD2.n88 VDD2.n87 104.615
R2600 VDD2.n88 VDD2.n3 104.615
R2601 VDD2.n95 VDD2.n3 104.615
R2602 VDD2.n96 VDD2.n95 104.615
R2603 VDD2.n104 VDD2.n103 63.3662
R2604 VDD2 VDD2.n209 63.3633
R2605 VDD2.n208 VDD2.n207 62.9756
R2606 VDD2.n102 VDD2.n101 62.9754
R2607 VDD2.t8 VDD2.n137 52.3082
R2608 VDD2.t1 VDD2.n31 52.3082
R2609 VDD2.n102 VDD2.n100 51.7862
R2610 VDD2.n206 VDD2.n205 51.1914
R2611 VDD2.n206 VDD2.n104 42.3683
R2612 VDD2.n139 VDD2.n138 15.6677
R2613 VDD2.n33 VDD2.n32 15.6677
R2614 VDD2.n186 VDD2.n115 13.1884
R2615 VDD2.n81 VDD2.n10 13.1884
R2616 VDD2.n187 VDD2.n113 12.8005
R2617 VDD2.n182 VDD2.n117 12.8005
R2618 VDD2.n142 VDD2.n141 12.8005
R2619 VDD2.n36 VDD2.n35 12.8005
R2620 VDD2.n77 VDD2.n76 12.8005
R2621 VDD2.n82 VDD2.n8 12.8005
R2622 VDD2.n191 VDD2.n190 12.0247
R2623 VDD2.n181 VDD2.n118 12.0247
R2624 VDD2.n145 VDD2.n136 12.0247
R2625 VDD2.n39 VDD2.n30 12.0247
R2626 VDD2.n75 VDD2.n12 12.0247
R2627 VDD2.n86 VDD2.n85 12.0247
R2628 VDD2.n194 VDD2.n111 11.249
R2629 VDD2.n178 VDD2.n177 11.249
R2630 VDD2.n146 VDD2.n134 11.249
R2631 VDD2.n40 VDD2.n28 11.249
R2632 VDD2.n72 VDD2.n71 11.249
R2633 VDD2.n89 VDD2.n6 11.249
R2634 VDD2.n195 VDD2.n109 10.4732
R2635 VDD2.n174 VDD2.n120 10.4732
R2636 VDD2.n150 VDD2.n149 10.4732
R2637 VDD2.n44 VDD2.n43 10.4732
R2638 VDD2.n68 VDD2.n14 10.4732
R2639 VDD2.n90 VDD2.n4 10.4732
R2640 VDD2.n199 VDD2.n198 9.69747
R2641 VDD2.n173 VDD2.n122 9.69747
R2642 VDD2.n153 VDD2.n132 9.69747
R2643 VDD2.n47 VDD2.n26 9.69747
R2644 VDD2.n67 VDD2.n16 9.69747
R2645 VDD2.n94 VDD2.n93 9.69747
R2646 VDD2.n205 VDD2.n204 9.45567
R2647 VDD2.n100 VDD2.n99 9.45567
R2648 VDD2.n165 VDD2.n164 9.3005
R2649 VDD2.n124 VDD2.n123 9.3005
R2650 VDD2.n171 VDD2.n170 9.3005
R2651 VDD2.n173 VDD2.n172 9.3005
R2652 VDD2.n120 VDD2.n119 9.3005
R2653 VDD2.n179 VDD2.n178 9.3005
R2654 VDD2.n181 VDD2.n180 9.3005
R2655 VDD2.n117 VDD2.n114 9.3005
R2656 VDD2.n204 VDD2.n203 9.3005
R2657 VDD2.n107 VDD2.n106 9.3005
R2658 VDD2.n198 VDD2.n197 9.3005
R2659 VDD2.n196 VDD2.n195 9.3005
R2660 VDD2.n111 VDD2.n110 9.3005
R2661 VDD2.n190 VDD2.n189 9.3005
R2662 VDD2.n188 VDD2.n187 9.3005
R2663 VDD2.n163 VDD2.n162 9.3005
R2664 VDD2.n128 VDD2.n127 9.3005
R2665 VDD2.n157 VDD2.n156 9.3005
R2666 VDD2.n155 VDD2.n154 9.3005
R2667 VDD2.n132 VDD2.n131 9.3005
R2668 VDD2.n149 VDD2.n148 9.3005
R2669 VDD2.n147 VDD2.n146 9.3005
R2670 VDD2.n136 VDD2.n135 9.3005
R2671 VDD2.n141 VDD2.n140 9.3005
R2672 VDD2.n99 VDD2.n98 9.3005
R2673 VDD2.n2 VDD2.n1 9.3005
R2674 VDD2.n93 VDD2.n92 9.3005
R2675 VDD2.n91 VDD2.n90 9.3005
R2676 VDD2.n6 VDD2.n5 9.3005
R2677 VDD2.n85 VDD2.n84 9.3005
R2678 VDD2.n83 VDD2.n82 9.3005
R2679 VDD2.n22 VDD2.n21 9.3005
R2680 VDD2.n51 VDD2.n50 9.3005
R2681 VDD2.n49 VDD2.n48 9.3005
R2682 VDD2.n26 VDD2.n25 9.3005
R2683 VDD2.n43 VDD2.n42 9.3005
R2684 VDD2.n41 VDD2.n40 9.3005
R2685 VDD2.n30 VDD2.n29 9.3005
R2686 VDD2.n35 VDD2.n34 9.3005
R2687 VDD2.n57 VDD2.n56 9.3005
R2688 VDD2.n59 VDD2.n58 9.3005
R2689 VDD2.n18 VDD2.n17 9.3005
R2690 VDD2.n65 VDD2.n64 9.3005
R2691 VDD2.n67 VDD2.n66 9.3005
R2692 VDD2.n14 VDD2.n13 9.3005
R2693 VDD2.n73 VDD2.n72 9.3005
R2694 VDD2.n75 VDD2.n74 9.3005
R2695 VDD2.n76 VDD2.n9 9.3005
R2696 VDD2.n202 VDD2.n107 8.92171
R2697 VDD2.n170 VDD2.n169 8.92171
R2698 VDD2.n154 VDD2.n130 8.92171
R2699 VDD2.n48 VDD2.n24 8.92171
R2700 VDD2.n64 VDD2.n63 8.92171
R2701 VDD2.n97 VDD2.n2 8.92171
R2702 VDD2.n203 VDD2.n105 8.14595
R2703 VDD2.n166 VDD2.n124 8.14595
R2704 VDD2.n158 VDD2.n157 8.14595
R2705 VDD2.n52 VDD2.n51 8.14595
R2706 VDD2.n60 VDD2.n18 8.14595
R2707 VDD2.n98 VDD2.n0 8.14595
R2708 VDD2.n165 VDD2.n126 7.3702
R2709 VDD2.n161 VDD2.n128 7.3702
R2710 VDD2.n55 VDD2.n22 7.3702
R2711 VDD2.n59 VDD2.n20 7.3702
R2712 VDD2.n162 VDD2.n126 6.59444
R2713 VDD2.n162 VDD2.n161 6.59444
R2714 VDD2.n56 VDD2.n55 6.59444
R2715 VDD2.n56 VDD2.n20 6.59444
R2716 VDD2.n205 VDD2.n105 5.81868
R2717 VDD2.n166 VDD2.n165 5.81868
R2718 VDD2.n158 VDD2.n128 5.81868
R2719 VDD2.n52 VDD2.n22 5.81868
R2720 VDD2.n60 VDD2.n59 5.81868
R2721 VDD2.n100 VDD2.n0 5.81868
R2722 VDD2.n203 VDD2.n202 5.04292
R2723 VDD2.n169 VDD2.n124 5.04292
R2724 VDD2.n157 VDD2.n130 5.04292
R2725 VDD2.n51 VDD2.n24 5.04292
R2726 VDD2.n63 VDD2.n18 5.04292
R2727 VDD2.n98 VDD2.n97 5.04292
R2728 VDD2.n140 VDD2.n139 4.38563
R2729 VDD2.n34 VDD2.n33 4.38563
R2730 VDD2.n199 VDD2.n107 4.26717
R2731 VDD2.n170 VDD2.n122 4.26717
R2732 VDD2.n154 VDD2.n153 4.26717
R2733 VDD2.n48 VDD2.n47 4.26717
R2734 VDD2.n64 VDD2.n16 4.26717
R2735 VDD2.n94 VDD2.n2 4.26717
R2736 VDD2.n198 VDD2.n109 3.49141
R2737 VDD2.n174 VDD2.n173 3.49141
R2738 VDD2.n150 VDD2.n132 3.49141
R2739 VDD2.n44 VDD2.n26 3.49141
R2740 VDD2.n68 VDD2.n67 3.49141
R2741 VDD2.n93 VDD2.n4 3.49141
R2742 VDD2.n195 VDD2.n194 2.71565
R2743 VDD2.n177 VDD2.n120 2.71565
R2744 VDD2.n149 VDD2.n134 2.71565
R2745 VDD2.n43 VDD2.n28 2.71565
R2746 VDD2.n71 VDD2.n14 2.71565
R2747 VDD2.n90 VDD2.n89 2.71565
R2748 VDD2.n191 VDD2.n111 1.93989
R2749 VDD2.n178 VDD2.n118 1.93989
R2750 VDD2.n146 VDD2.n145 1.93989
R2751 VDD2.n40 VDD2.n39 1.93989
R2752 VDD2.n72 VDD2.n12 1.93989
R2753 VDD2.n86 VDD2.n6 1.93989
R2754 VDD2.n190 VDD2.n113 1.16414
R2755 VDD2.n182 VDD2.n181 1.16414
R2756 VDD2.n142 VDD2.n136 1.16414
R2757 VDD2.n36 VDD2.n30 1.16414
R2758 VDD2.n77 VDD2.n75 1.16414
R2759 VDD2.n85 VDD2.n8 1.16414
R2760 VDD2.n209 VDD2.t0 1.07893
R2761 VDD2.n209 VDD2.t3 1.07893
R2762 VDD2.n207 VDD2.t2 1.07893
R2763 VDD2.n207 VDD2.t5 1.07893
R2764 VDD2.n103 VDD2.t9 1.07893
R2765 VDD2.n103 VDD2.t4 1.07893
R2766 VDD2.n101 VDD2.t6 1.07893
R2767 VDD2.n101 VDD2.t7 1.07893
R2768 VDD2.n208 VDD2.n206 0.595328
R2769 VDD2.n187 VDD2.n186 0.388379
R2770 VDD2.n117 VDD2.n115 0.388379
R2771 VDD2.n141 VDD2.n138 0.388379
R2772 VDD2.n35 VDD2.n32 0.388379
R2773 VDD2.n76 VDD2.n10 0.388379
R2774 VDD2.n82 VDD2.n81 0.388379
R2775 VDD2 VDD2.n208 0.207397
R2776 VDD2.n204 VDD2.n106 0.155672
R2777 VDD2.n197 VDD2.n106 0.155672
R2778 VDD2.n197 VDD2.n196 0.155672
R2779 VDD2.n196 VDD2.n110 0.155672
R2780 VDD2.n189 VDD2.n110 0.155672
R2781 VDD2.n189 VDD2.n188 0.155672
R2782 VDD2.n188 VDD2.n114 0.155672
R2783 VDD2.n180 VDD2.n114 0.155672
R2784 VDD2.n180 VDD2.n179 0.155672
R2785 VDD2.n179 VDD2.n119 0.155672
R2786 VDD2.n172 VDD2.n119 0.155672
R2787 VDD2.n172 VDD2.n171 0.155672
R2788 VDD2.n171 VDD2.n123 0.155672
R2789 VDD2.n164 VDD2.n123 0.155672
R2790 VDD2.n164 VDD2.n163 0.155672
R2791 VDD2.n163 VDD2.n127 0.155672
R2792 VDD2.n156 VDD2.n127 0.155672
R2793 VDD2.n156 VDD2.n155 0.155672
R2794 VDD2.n155 VDD2.n131 0.155672
R2795 VDD2.n148 VDD2.n131 0.155672
R2796 VDD2.n148 VDD2.n147 0.155672
R2797 VDD2.n147 VDD2.n135 0.155672
R2798 VDD2.n140 VDD2.n135 0.155672
R2799 VDD2.n34 VDD2.n29 0.155672
R2800 VDD2.n41 VDD2.n29 0.155672
R2801 VDD2.n42 VDD2.n41 0.155672
R2802 VDD2.n42 VDD2.n25 0.155672
R2803 VDD2.n49 VDD2.n25 0.155672
R2804 VDD2.n50 VDD2.n49 0.155672
R2805 VDD2.n50 VDD2.n21 0.155672
R2806 VDD2.n57 VDD2.n21 0.155672
R2807 VDD2.n58 VDD2.n57 0.155672
R2808 VDD2.n58 VDD2.n17 0.155672
R2809 VDD2.n65 VDD2.n17 0.155672
R2810 VDD2.n66 VDD2.n65 0.155672
R2811 VDD2.n66 VDD2.n13 0.155672
R2812 VDD2.n73 VDD2.n13 0.155672
R2813 VDD2.n74 VDD2.n73 0.155672
R2814 VDD2.n74 VDD2.n9 0.155672
R2815 VDD2.n83 VDD2.n9 0.155672
R2816 VDD2.n84 VDD2.n83 0.155672
R2817 VDD2.n84 VDD2.n5 0.155672
R2818 VDD2.n91 VDD2.n5 0.155672
R2819 VDD2.n92 VDD2.n91 0.155672
R2820 VDD2.n92 VDD2.n1 0.155672
R2821 VDD2.n99 VDD2.n1 0.155672
R2822 VDD2.n104 VDD2.n102 0.0938609
C0 VTAIL VP 6.05722f
C1 VDD1 VP 6.80085f
C2 VP VDD2 0.299829f
C3 VTAIL VN 6.04215f
C4 VDD1 VN 0.148563f
C5 VN VDD2 6.65725f
C6 VTAIL VDD1 28.3146f
C7 VTAIL VDD2 28.3407f
C8 VDD1 VDD2 0.764582f
C9 VP VN 6.27477f
C10 VDD2 B 5.733803f
C11 VDD1 B 5.606833f
C12 VTAIL B 8.35424f
C13 VN B 8.877561f
C14 VP B 6.293596f
C15 VDD2.n0 B 0.042402f
C16 VDD2.n1 B 0.028524f
C17 VDD2.n2 B 0.015327f
C18 VDD2.n3 B 0.036229f
C19 VDD2.n4 B 0.016229f
C20 VDD2.n5 B 0.028524f
C21 VDD2.n6 B 0.015327f
C22 VDD2.n7 B 0.036229f
C23 VDD2.n8 B 0.016229f
C24 VDD2.n9 B 0.028524f
C25 VDD2.n10 B 0.015778f
C26 VDD2.n11 B 0.036229f
C27 VDD2.n12 B 0.016229f
C28 VDD2.n13 B 0.028524f
C29 VDD2.n14 B 0.015327f
C30 VDD2.n15 B 0.036229f
C31 VDD2.n16 B 0.016229f
C32 VDD2.n17 B 0.028524f
C33 VDD2.n18 B 0.015327f
C34 VDD2.n19 B 0.036229f
C35 VDD2.n20 B 0.016229f
C36 VDD2.n21 B 0.028524f
C37 VDD2.n22 B 0.015327f
C38 VDD2.n23 B 0.036229f
C39 VDD2.n24 B 0.016229f
C40 VDD2.n25 B 0.028524f
C41 VDD2.n26 B 0.015327f
C42 VDD2.n27 B 0.036229f
C43 VDD2.n28 B 0.016229f
C44 VDD2.n29 B 0.028524f
C45 VDD2.n30 B 0.015327f
C46 VDD2.n31 B 0.027172f
C47 VDD2.n32 B 0.021401f
C48 VDD2.t1 B 0.060066f
C49 VDD2.n33 B 0.210069f
C50 VDD2.n34 B 2.29505f
C51 VDD2.n35 B 0.015327f
C52 VDD2.n36 B 0.016229f
C53 VDD2.n37 B 0.036229f
C54 VDD2.n38 B 0.036229f
C55 VDD2.n39 B 0.016229f
C56 VDD2.n40 B 0.015327f
C57 VDD2.n41 B 0.028524f
C58 VDD2.n42 B 0.028524f
C59 VDD2.n43 B 0.015327f
C60 VDD2.n44 B 0.016229f
C61 VDD2.n45 B 0.036229f
C62 VDD2.n46 B 0.036229f
C63 VDD2.n47 B 0.016229f
C64 VDD2.n48 B 0.015327f
C65 VDD2.n49 B 0.028524f
C66 VDD2.n50 B 0.028524f
C67 VDD2.n51 B 0.015327f
C68 VDD2.n52 B 0.016229f
C69 VDD2.n53 B 0.036229f
C70 VDD2.n54 B 0.036229f
C71 VDD2.n55 B 0.016229f
C72 VDD2.n56 B 0.015327f
C73 VDD2.n57 B 0.028524f
C74 VDD2.n58 B 0.028524f
C75 VDD2.n59 B 0.015327f
C76 VDD2.n60 B 0.016229f
C77 VDD2.n61 B 0.036229f
C78 VDD2.n62 B 0.036229f
C79 VDD2.n63 B 0.016229f
C80 VDD2.n64 B 0.015327f
C81 VDD2.n65 B 0.028524f
C82 VDD2.n66 B 0.028524f
C83 VDD2.n67 B 0.015327f
C84 VDD2.n68 B 0.016229f
C85 VDD2.n69 B 0.036229f
C86 VDD2.n70 B 0.036229f
C87 VDD2.n71 B 0.016229f
C88 VDD2.n72 B 0.015327f
C89 VDD2.n73 B 0.028524f
C90 VDD2.n74 B 0.028524f
C91 VDD2.n75 B 0.015327f
C92 VDD2.n76 B 0.015327f
C93 VDD2.n77 B 0.016229f
C94 VDD2.n78 B 0.036229f
C95 VDD2.n79 B 0.036229f
C96 VDD2.n80 B 0.036229f
C97 VDD2.n81 B 0.015778f
C98 VDD2.n82 B 0.015327f
C99 VDD2.n83 B 0.028524f
C100 VDD2.n84 B 0.028524f
C101 VDD2.n85 B 0.015327f
C102 VDD2.n86 B 0.016229f
C103 VDD2.n87 B 0.036229f
C104 VDD2.n88 B 0.036229f
C105 VDD2.n89 B 0.016229f
C106 VDD2.n90 B 0.015327f
C107 VDD2.n91 B 0.028524f
C108 VDD2.n92 B 0.028524f
C109 VDD2.n93 B 0.015327f
C110 VDD2.n94 B 0.016229f
C111 VDD2.n95 B 0.036229f
C112 VDD2.n96 B 0.082513f
C113 VDD2.n97 B 0.016229f
C114 VDD2.n98 B 0.015327f
C115 VDD2.n99 B 0.070608f
C116 VDD2.n100 B 0.067679f
C117 VDD2.t6 B 0.413843f
C118 VDD2.t7 B 0.413843f
C119 VDD2.n101 B 3.77589f
C120 VDD2.n102 B 0.415795f
C121 VDD2.t9 B 0.413843f
C122 VDD2.t4 B 0.413843f
C123 VDD2.n103 B 3.77797f
C124 VDD2.n104 B 2.41008f
C125 VDD2.n105 B 0.042402f
C126 VDD2.n106 B 0.028524f
C127 VDD2.n107 B 0.015327f
C128 VDD2.n108 B 0.036229f
C129 VDD2.n109 B 0.016229f
C130 VDD2.n110 B 0.028524f
C131 VDD2.n111 B 0.015327f
C132 VDD2.n112 B 0.036229f
C133 VDD2.n113 B 0.016229f
C134 VDD2.n114 B 0.028524f
C135 VDD2.n115 B 0.015778f
C136 VDD2.n116 B 0.036229f
C137 VDD2.n117 B 0.015327f
C138 VDD2.n118 B 0.016229f
C139 VDD2.n119 B 0.028524f
C140 VDD2.n120 B 0.015327f
C141 VDD2.n121 B 0.036229f
C142 VDD2.n122 B 0.016229f
C143 VDD2.n123 B 0.028524f
C144 VDD2.n124 B 0.015327f
C145 VDD2.n125 B 0.036229f
C146 VDD2.n126 B 0.016229f
C147 VDD2.n127 B 0.028524f
C148 VDD2.n128 B 0.015327f
C149 VDD2.n129 B 0.036229f
C150 VDD2.n130 B 0.016229f
C151 VDD2.n131 B 0.028524f
C152 VDD2.n132 B 0.015327f
C153 VDD2.n133 B 0.036229f
C154 VDD2.n134 B 0.016229f
C155 VDD2.n135 B 0.028524f
C156 VDD2.n136 B 0.015327f
C157 VDD2.n137 B 0.027172f
C158 VDD2.n138 B 0.021401f
C159 VDD2.t8 B 0.060066f
C160 VDD2.n139 B 0.210069f
C161 VDD2.n140 B 2.29505f
C162 VDD2.n141 B 0.015327f
C163 VDD2.n142 B 0.016229f
C164 VDD2.n143 B 0.036229f
C165 VDD2.n144 B 0.036229f
C166 VDD2.n145 B 0.016229f
C167 VDD2.n146 B 0.015327f
C168 VDD2.n147 B 0.028524f
C169 VDD2.n148 B 0.028524f
C170 VDD2.n149 B 0.015327f
C171 VDD2.n150 B 0.016229f
C172 VDD2.n151 B 0.036229f
C173 VDD2.n152 B 0.036229f
C174 VDD2.n153 B 0.016229f
C175 VDD2.n154 B 0.015327f
C176 VDD2.n155 B 0.028524f
C177 VDD2.n156 B 0.028524f
C178 VDD2.n157 B 0.015327f
C179 VDD2.n158 B 0.016229f
C180 VDD2.n159 B 0.036229f
C181 VDD2.n160 B 0.036229f
C182 VDD2.n161 B 0.016229f
C183 VDD2.n162 B 0.015327f
C184 VDD2.n163 B 0.028524f
C185 VDD2.n164 B 0.028524f
C186 VDD2.n165 B 0.015327f
C187 VDD2.n166 B 0.016229f
C188 VDD2.n167 B 0.036229f
C189 VDD2.n168 B 0.036229f
C190 VDD2.n169 B 0.016229f
C191 VDD2.n170 B 0.015327f
C192 VDD2.n171 B 0.028524f
C193 VDD2.n172 B 0.028524f
C194 VDD2.n173 B 0.015327f
C195 VDD2.n174 B 0.016229f
C196 VDD2.n175 B 0.036229f
C197 VDD2.n176 B 0.036229f
C198 VDD2.n177 B 0.016229f
C199 VDD2.n178 B 0.015327f
C200 VDD2.n179 B 0.028524f
C201 VDD2.n180 B 0.028524f
C202 VDD2.n181 B 0.015327f
C203 VDD2.n182 B 0.016229f
C204 VDD2.n183 B 0.036229f
C205 VDD2.n184 B 0.036229f
C206 VDD2.n185 B 0.036229f
C207 VDD2.n186 B 0.015778f
C208 VDD2.n187 B 0.015327f
C209 VDD2.n188 B 0.028524f
C210 VDD2.n189 B 0.028524f
C211 VDD2.n190 B 0.015327f
C212 VDD2.n191 B 0.016229f
C213 VDD2.n192 B 0.036229f
C214 VDD2.n193 B 0.036229f
C215 VDD2.n194 B 0.016229f
C216 VDD2.n195 B 0.015327f
C217 VDD2.n196 B 0.028524f
C218 VDD2.n197 B 0.028524f
C219 VDD2.n198 B 0.015327f
C220 VDD2.n199 B 0.016229f
C221 VDD2.n200 B 0.036229f
C222 VDD2.n201 B 0.082513f
C223 VDD2.n202 B 0.016229f
C224 VDD2.n203 B 0.015327f
C225 VDD2.n204 B 0.070608f
C226 VDD2.n205 B 0.066389f
C227 VDD2.n206 B 2.87151f
C228 VDD2.t2 B 0.413843f
C229 VDD2.t5 B 0.413843f
C230 VDD2.n207 B 3.7759f
C231 VDD2.n208 B 0.308152f
C232 VDD2.t0 B 0.413843f
C233 VDD2.t3 B 0.413843f
C234 VDD2.n209 B 3.77794f
C235 VN.n0 B 0.051712f
C236 VN.t2 B 0.968829f
C237 VN.n1 B 0.363579f
C238 VN.t8 B 0.974555f
C239 VN.n2 B 0.365478f
C240 VN.t3 B 0.968829f
C241 VN.n3 B 0.379139f
C242 VN.n4 B 0.011734f
C243 VN.n5 B 0.158609f
C244 VN.n6 B 0.051712f
C245 VN.n7 B 0.011734f
C246 VN.t0 B 0.968829f
C247 VN.n8 B 0.379139f
C248 VN.t5 B 0.968829f
C249 VN.n9 B 0.37085f
C250 VN.n10 B 0.040075f
C251 VN.n11 B 0.051712f
C252 VN.t4 B 0.968829f
C253 VN.n12 B 0.363579f
C254 VN.t6 B 0.974555f
C255 VN.n13 B 0.365478f
C256 VN.t9 B 0.968829f
C257 VN.n14 B 0.379139f
C258 VN.n15 B 0.011734f
C259 VN.n16 B 0.158609f
C260 VN.n17 B 0.051712f
C261 VN.n18 B 0.011734f
C262 VN.t7 B 0.968829f
C263 VN.n19 B 0.379139f
C264 VN.t1 B 0.968829f
C265 VN.n20 B 0.37085f
C266 VN.n21 B 2.48349f
C267 VDD1.n0 B 0.042396f
C268 VDD1.n1 B 0.02852f
C269 VDD1.n2 B 0.015325f
C270 VDD1.n3 B 0.036223f
C271 VDD1.n4 B 0.016227f
C272 VDD1.n5 B 0.02852f
C273 VDD1.n6 B 0.015325f
C274 VDD1.n7 B 0.036223f
C275 VDD1.n8 B 0.016227f
C276 VDD1.n9 B 0.02852f
C277 VDD1.n10 B 0.015776f
C278 VDD1.n11 B 0.036223f
C279 VDD1.n12 B 0.015325f
C280 VDD1.n13 B 0.016227f
C281 VDD1.n14 B 0.02852f
C282 VDD1.n15 B 0.015325f
C283 VDD1.n16 B 0.036223f
C284 VDD1.n17 B 0.016227f
C285 VDD1.n18 B 0.02852f
C286 VDD1.n19 B 0.015325f
C287 VDD1.n20 B 0.036223f
C288 VDD1.n21 B 0.016227f
C289 VDD1.n22 B 0.02852f
C290 VDD1.n23 B 0.015325f
C291 VDD1.n24 B 0.036223f
C292 VDD1.n25 B 0.016227f
C293 VDD1.n26 B 0.02852f
C294 VDD1.n27 B 0.015325f
C295 VDD1.n28 B 0.036223f
C296 VDD1.n29 B 0.016227f
C297 VDD1.n30 B 0.02852f
C298 VDD1.n31 B 0.015325f
C299 VDD1.n32 B 0.027167f
C300 VDD1.n33 B 0.021398f
C301 VDD1.t5 B 0.060056f
C302 VDD1.n34 B 0.210037f
C303 VDD1.n35 B 2.2947f
C304 VDD1.n36 B 0.015325f
C305 VDD1.n37 B 0.016227f
C306 VDD1.n38 B 0.036223f
C307 VDD1.n39 B 0.036223f
C308 VDD1.n40 B 0.016227f
C309 VDD1.n41 B 0.015325f
C310 VDD1.n42 B 0.02852f
C311 VDD1.n43 B 0.02852f
C312 VDD1.n44 B 0.015325f
C313 VDD1.n45 B 0.016227f
C314 VDD1.n46 B 0.036223f
C315 VDD1.n47 B 0.036223f
C316 VDD1.n48 B 0.016227f
C317 VDD1.n49 B 0.015325f
C318 VDD1.n50 B 0.02852f
C319 VDD1.n51 B 0.02852f
C320 VDD1.n52 B 0.015325f
C321 VDD1.n53 B 0.016227f
C322 VDD1.n54 B 0.036223f
C323 VDD1.n55 B 0.036223f
C324 VDD1.n56 B 0.016227f
C325 VDD1.n57 B 0.015325f
C326 VDD1.n58 B 0.02852f
C327 VDD1.n59 B 0.02852f
C328 VDD1.n60 B 0.015325f
C329 VDD1.n61 B 0.016227f
C330 VDD1.n62 B 0.036223f
C331 VDD1.n63 B 0.036223f
C332 VDD1.n64 B 0.016227f
C333 VDD1.n65 B 0.015325f
C334 VDD1.n66 B 0.02852f
C335 VDD1.n67 B 0.02852f
C336 VDD1.n68 B 0.015325f
C337 VDD1.n69 B 0.016227f
C338 VDD1.n70 B 0.036223f
C339 VDD1.n71 B 0.036223f
C340 VDD1.n72 B 0.016227f
C341 VDD1.n73 B 0.015325f
C342 VDD1.n74 B 0.02852f
C343 VDD1.n75 B 0.02852f
C344 VDD1.n76 B 0.015325f
C345 VDD1.n77 B 0.016227f
C346 VDD1.n78 B 0.036223f
C347 VDD1.n79 B 0.036223f
C348 VDD1.n80 B 0.036223f
C349 VDD1.n81 B 0.015776f
C350 VDD1.n82 B 0.015325f
C351 VDD1.n83 B 0.02852f
C352 VDD1.n84 B 0.02852f
C353 VDD1.n85 B 0.015325f
C354 VDD1.n86 B 0.016227f
C355 VDD1.n87 B 0.036223f
C356 VDD1.n88 B 0.036223f
C357 VDD1.n89 B 0.016227f
C358 VDD1.n90 B 0.015325f
C359 VDD1.n91 B 0.02852f
C360 VDD1.n92 B 0.02852f
C361 VDD1.n93 B 0.015325f
C362 VDD1.n94 B 0.016227f
C363 VDD1.n95 B 0.036223f
C364 VDD1.n96 B 0.0825f
C365 VDD1.n97 B 0.016227f
C366 VDD1.n98 B 0.015325f
C367 VDD1.n99 B 0.070597f
C368 VDD1.n100 B 0.067669f
C369 VDD1.t2 B 0.41378f
C370 VDD1.t9 B 0.41378f
C371 VDD1.n101 B 3.77532f
C372 VDD1.n102 B 0.419072f
C373 VDD1.n103 B 0.042396f
C374 VDD1.n104 B 0.02852f
C375 VDD1.n105 B 0.015325f
C376 VDD1.n106 B 0.036223f
C377 VDD1.n107 B 0.016227f
C378 VDD1.n108 B 0.02852f
C379 VDD1.n109 B 0.015325f
C380 VDD1.n110 B 0.036223f
C381 VDD1.n111 B 0.016227f
C382 VDD1.n112 B 0.02852f
C383 VDD1.n113 B 0.015776f
C384 VDD1.n114 B 0.036223f
C385 VDD1.n115 B 0.016227f
C386 VDD1.n116 B 0.02852f
C387 VDD1.n117 B 0.015325f
C388 VDD1.n118 B 0.036223f
C389 VDD1.n119 B 0.016227f
C390 VDD1.n120 B 0.02852f
C391 VDD1.n121 B 0.015325f
C392 VDD1.n122 B 0.036223f
C393 VDD1.n123 B 0.016227f
C394 VDD1.n124 B 0.02852f
C395 VDD1.n125 B 0.015325f
C396 VDD1.n126 B 0.036223f
C397 VDD1.n127 B 0.016227f
C398 VDD1.n128 B 0.02852f
C399 VDD1.n129 B 0.015325f
C400 VDD1.n130 B 0.036223f
C401 VDD1.n131 B 0.016227f
C402 VDD1.n132 B 0.02852f
C403 VDD1.n133 B 0.015325f
C404 VDD1.n134 B 0.027167f
C405 VDD1.n135 B 0.021398f
C406 VDD1.t6 B 0.060056f
C407 VDD1.n136 B 0.210037f
C408 VDD1.n137 B 2.2947f
C409 VDD1.n138 B 0.015325f
C410 VDD1.n139 B 0.016227f
C411 VDD1.n140 B 0.036223f
C412 VDD1.n141 B 0.036223f
C413 VDD1.n142 B 0.016227f
C414 VDD1.n143 B 0.015325f
C415 VDD1.n144 B 0.02852f
C416 VDD1.n145 B 0.02852f
C417 VDD1.n146 B 0.015325f
C418 VDD1.n147 B 0.016227f
C419 VDD1.n148 B 0.036223f
C420 VDD1.n149 B 0.036223f
C421 VDD1.n150 B 0.016227f
C422 VDD1.n151 B 0.015325f
C423 VDD1.n152 B 0.02852f
C424 VDD1.n153 B 0.02852f
C425 VDD1.n154 B 0.015325f
C426 VDD1.n155 B 0.016227f
C427 VDD1.n156 B 0.036223f
C428 VDD1.n157 B 0.036223f
C429 VDD1.n158 B 0.016227f
C430 VDD1.n159 B 0.015325f
C431 VDD1.n160 B 0.02852f
C432 VDD1.n161 B 0.02852f
C433 VDD1.n162 B 0.015325f
C434 VDD1.n163 B 0.016227f
C435 VDD1.n164 B 0.036223f
C436 VDD1.n165 B 0.036223f
C437 VDD1.n166 B 0.016227f
C438 VDD1.n167 B 0.015325f
C439 VDD1.n168 B 0.02852f
C440 VDD1.n169 B 0.02852f
C441 VDD1.n170 B 0.015325f
C442 VDD1.n171 B 0.016227f
C443 VDD1.n172 B 0.036223f
C444 VDD1.n173 B 0.036223f
C445 VDD1.n174 B 0.016227f
C446 VDD1.n175 B 0.015325f
C447 VDD1.n176 B 0.02852f
C448 VDD1.n177 B 0.02852f
C449 VDD1.n178 B 0.015325f
C450 VDD1.n179 B 0.015325f
C451 VDD1.n180 B 0.016227f
C452 VDD1.n181 B 0.036223f
C453 VDD1.n182 B 0.036223f
C454 VDD1.n183 B 0.036223f
C455 VDD1.n184 B 0.015776f
C456 VDD1.n185 B 0.015325f
C457 VDD1.n186 B 0.02852f
C458 VDD1.n187 B 0.02852f
C459 VDD1.n188 B 0.015325f
C460 VDD1.n189 B 0.016227f
C461 VDD1.n190 B 0.036223f
C462 VDD1.n191 B 0.036223f
C463 VDD1.n192 B 0.016227f
C464 VDD1.n193 B 0.015325f
C465 VDD1.n194 B 0.02852f
C466 VDD1.n195 B 0.02852f
C467 VDD1.n196 B 0.015325f
C468 VDD1.n197 B 0.016227f
C469 VDD1.n198 B 0.036223f
C470 VDD1.n199 B 0.0825f
C471 VDD1.n200 B 0.016227f
C472 VDD1.n201 B 0.015325f
C473 VDD1.n202 B 0.070597f
C474 VDD1.n203 B 0.067669f
C475 VDD1.t1 B 0.41378f
C476 VDD1.t7 B 0.41378f
C477 VDD1.n204 B 3.77531f
C478 VDD1.n205 B 0.415732f
C479 VDD1.t8 B 0.41378f
C480 VDD1.t4 B 0.41378f
C481 VDD1.n206 B 3.7774f
C482 VDD1.n207 B 2.48978f
C483 VDD1.t3 B 0.41378f
C484 VDD1.t0 B 0.41378f
C485 VDD1.n208 B 3.77531f
C486 VDD1.n209 B 3.12033f
C487 VTAIL.t19 B 0.420274f
C488 VTAIL.t4 B 0.420274f
C489 VTAIL.n0 B 3.75076f
C490 VTAIL.n1 B 0.401232f
C491 VTAIL.n2 B 0.043061f
C492 VTAIL.n3 B 0.028967f
C493 VTAIL.n4 B 0.015566f
C494 VTAIL.n5 B 0.036792f
C495 VTAIL.n6 B 0.016481f
C496 VTAIL.n7 B 0.028967f
C497 VTAIL.n8 B 0.015566f
C498 VTAIL.n9 B 0.036792f
C499 VTAIL.n10 B 0.016481f
C500 VTAIL.n11 B 0.028967f
C501 VTAIL.n12 B 0.016024f
C502 VTAIL.n13 B 0.036792f
C503 VTAIL.n14 B 0.016481f
C504 VTAIL.n15 B 0.028967f
C505 VTAIL.n16 B 0.015566f
C506 VTAIL.n17 B 0.036792f
C507 VTAIL.n18 B 0.016481f
C508 VTAIL.n19 B 0.028967f
C509 VTAIL.n20 B 0.015566f
C510 VTAIL.n21 B 0.036792f
C511 VTAIL.n22 B 0.016481f
C512 VTAIL.n23 B 0.028967f
C513 VTAIL.n24 B 0.015566f
C514 VTAIL.n25 B 0.036792f
C515 VTAIL.n26 B 0.016481f
C516 VTAIL.n27 B 0.028967f
C517 VTAIL.n28 B 0.015566f
C518 VTAIL.n29 B 0.036792f
C519 VTAIL.n30 B 0.016481f
C520 VTAIL.n31 B 0.028967f
C521 VTAIL.n32 B 0.015566f
C522 VTAIL.n33 B 0.027594f
C523 VTAIL.n34 B 0.021734f
C524 VTAIL.t7 B 0.060999f
C525 VTAIL.n35 B 0.213333f
C526 VTAIL.n36 B 2.33071f
C527 VTAIL.n37 B 0.015566f
C528 VTAIL.n38 B 0.016481f
C529 VTAIL.n39 B 0.036792f
C530 VTAIL.n40 B 0.036792f
C531 VTAIL.n41 B 0.016481f
C532 VTAIL.n42 B 0.015566f
C533 VTAIL.n43 B 0.028967f
C534 VTAIL.n44 B 0.028967f
C535 VTAIL.n45 B 0.015566f
C536 VTAIL.n46 B 0.016481f
C537 VTAIL.n47 B 0.036792f
C538 VTAIL.n48 B 0.036792f
C539 VTAIL.n49 B 0.016481f
C540 VTAIL.n50 B 0.015566f
C541 VTAIL.n51 B 0.028967f
C542 VTAIL.n52 B 0.028967f
C543 VTAIL.n53 B 0.015566f
C544 VTAIL.n54 B 0.016481f
C545 VTAIL.n55 B 0.036792f
C546 VTAIL.n56 B 0.036792f
C547 VTAIL.n57 B 0.016481f
C548 VTAIL.n58 B 0.015566f
C549 VTAIL.n59 B 0.028967f
C550 VTAIL.n60 B 0.028967f
C551 VTAIL.n61 B 0.015566f
C552 VTAIL.n62 B 0.016481f
C553 VTAIL.n63 B 0.036792f
C554 VTAIL.n64 B 0.036792f
C555 VTAIL.n65 B 0.016481f
C556 VTAIL.n66 B 0.015566f
C557 VTAIL.n67 B 0.028967f
C558 VTAIL.n68 B 0.028967f
C559 VTAIL.n69 B 0.015566f
C560 VTAIL.n70 B 0.016481f
C561 VTAIL.n71 B 0.036792f
C562 VTAIL.n72 B 0.036792f
C563 VTAIL.n73 B 0.016481f
C564 VTAIL.n74 B 0.015566f
C565 VTAIL.n75 B 0.028967f
C566 VTAIL.n76 B 0.028967f
C567 VTAIL.n77 B 0.015566f
C568 VTAIL.n78 B 0.015566f
C569 VTAIL.n79 B 0.016481f
C570 VTAIL.n80 B 0.036792f
C571 VTAIL.n81 B 0.036792f
C572 VTAIL.n82 B 0.036792f
C573 VTAIL.n83 B 0.016024f
C574 VTAIL.n84 B 0.015566f
C575 VTAIL.n85 B 0.028967f
C576 VTAIL.n86 B 0.028967f
C577 VTAIL.n87 B 0.015566f
C578 VTAIL.n88 B 0.016481f
C579 VTAIL.n89 B 0.036792f
C580 VTAIL.n90 B 0.036792f
C581 VTAIL.n91 B 0.016481f
C582 VTAIL.n92 B 0.015566f
C583 VTAIL.n93 B 0.028967f
C584 VTAIL.n94 B 0.028967f
C585 VTAIL.n95 B 0.015566f
C586 VTAIL.n96 B 0.016481f
C587 VTAIL.n97 B 0.036792f
C588 VTAIL.n98 B 0.083795f
C589 VTAIL.n99 B 0.016481f
C590 VTAIL.n100 B 0.015566f
C591 VTAIL.n101 B 0.071705f
C592 VTAIL.n102 B 0.047454f
C593 VTAIL.n103 B 0.154558f
C594 VTAIL.t14 B 0.420274f
C595 VTAIL.t8 B 0.420274f
C596 VTAIL.n104 B 3.75076f
C597 VTAIL.n105 B 0.393588f
C598 VTAIL.t15 B 0.420274f
C599 VTAIL.t10 B 0.420274f
C600 VTAIL.n106 B 3.75076f
C601 VTAIL.n107 B 2.31992f
C602 VTAIL.t5 B 0.420274f
C603 VTAIL.t18 B 0.420274f
C604 VTAIL.n108 B 3.75078f
C605 VTAIL.n109 B 2.3199f
C606 VTAIL.t3 B 0.420274f
C607 VTAIL.t2 B 0.420274f
C608 VTAIL.n110 B 3.75078f
C609 VTAIL.n111 B 0.393572f
C610 VTAIL.n112 B 0.043061f
C611 VTAIL.n113 B 0.028967f
C612 VTAIL.n114 B 0.015566f
C613 VTAIL.n115 B 0.036792f
C614 VTAIL.n116 B 0.016481f
C615 VTAIL.n117 B 0.028967f
C616 VTAIL.n118 B 0.015566f
C617 VTAIL.n119 B 0.036792f
C618 VTAIL.n120 B 0.016481f
C619 VTAIL.n121 B 0.028967f
C620 VTAIL.n122 B 0.016024f
C621 VTAIL.n123 B 0.036792f
C622 VTAIL.n124 B 0.015566f
C623 VTAIL.n125 B 0.016481f
C624 VTAIL.n126 B 0.028967f
C625 VTAIL.n127 B 0.015566f
C626 VTAIL.n128 B 0.036792f
C627 VTAIL.n129 B 0.016481f
C628 VTAIL.n130 B 0.028967f
C629 VTAIL.n131 B 0.015566f
C630 VTAIL.n132 B 0.036792f
C631 VTAIL.n133 B 0.016481f
C632 VTAIL.n134 B 0.028967f
C633 VTAIL.n135 B 0.015566f
C634 VTAIL.n136 B 0.036792f
C635 VTAIL.n137 B 0.016481f
C636 VTAIL.n138 B 0.028967f
C637 VTAIL.n139 B 0.015566f
C638 VTAIL.n140 B 0.036792f
C639 VTAIL.n141 B 0.016481f
C640 VTAIL.n142 B 0.028967f
C641 VTAIL.n143 B 0.015566f
C642 VTAIL.n144 B 0.027594f
C643 VTAIL.n145 B 0.021734f
C644 VTAIL.t17 B 0.060999f
C645 VTAIL.n146 B 0.213333f
C646 VTAIL.n147 B 2.33071f
C647 VTAIL.n148 B 0.015566f
C648 VTAIL.n149 B 0.016481f
C649 VTAIL.n150 B 0.036792f
C650 VTAIL.n151 B 0.036792f
C651 VTAIL.n152 B 0.016481f
C652 VTAIL.n153 B 0.015566f
C653 VTAIL.n154 B 0.028967f
C654 VTAIL.n155 B 0.028967f
C655 VTAIL.n156 B 0.015566f
C656 VTAIL.n157 B 0.016481f
C657 VTAIL.n158 B 0.036792f
C658 VTAIL.n159 B 0.036792f
C659 VTAIL.n160 B 0.016481f
C660 VTAIL.n161 B 0.015566f
C661 VTAIL.n162 B 0.028967f
C662 VTAIL.n163 B 0.028967f
C663 VTAIL.n164 B 0.015566f
C664 VTAIL.n165 B 0.016481f
C665 VTAIL.n166 B 0.036792f
C666 VTAIL.n167 B 0.036792f
C667 VTAIL.n168 B 0.016481f
C668 VTAIL.n169 B 0.015566f
C669 VTAIL.n170 B 0.028967f
C670 VTAIL.n171 B 0.028967f
C671 VTAIL.n172 B 0.015566f
C672 VTAIL.n173 B 0.016481f
C673 VTAIL.n174 B 0.036792f
C674 VTAIL.n175 B 0.036792f
C675 VTAIL.n176 B 0.016481f
C676 VTAIL.n177 B 0.015566f
C677 VTAIL.n178 B 0.028967f
C678 VTAIL.n179 B 0.028967f
C679 VTAIL.n180 B 0.015566f
C680 VTAIL.n181 B 0.016481f
C681 VTAIL.n182 B 0.036792f
C682 VTAIL.n183 B 0.036792f
C683 VTAIL.n184 B 0.016481f
C684 VTAIL.n185 B 0.015566f
C685 VTAIL.n186 B 0.028967f
C686 VTAIL.n187 B 0.028967f
C687 VTAIL.n188 B 0.015566f
C688 VTAIL.n189 B 0.016481f
C689 VTAIL.n190 B 0.036792f
C690 VTAIL.n191 B 0.036792f
C691 VTAIL.n192 B 0.036792f
C692 VTAIL.n193 B 0.016024f
C693 VTAIL.n194 B 0.015566f
C694 VTAIL.n195 B 0.028967f
C695 VTAIL.n196 B 0.028967f
C696 VTAIL.n197 B 0.015566f
C697 VTAIL.n198 B 0.016481f
C698 VTAIL.n199 B 0.036792f
C699 VTAIL.n200 B 0.036792f
C700 VTAIL.n201 B 0.016481f
C701 VTAIL.n202 B 0.015566f
C702 VTAIL.n203 B 0.028967f
C703 VTAIL.n204 B 0.028967f
C704 VTAIL.n205 B 0.015566f
C705 VTAIL.n206 B 0.016481f
C706 VTAIL.n207 B 0.036792f
C707 VTAIL.n208 B 0.083795f
C708 VTAIL.n209 B 0.016481f
C709 VTAIL.n210 B 0.015566f
C710 VTAIL.n211 B 0.071705f
C711 VTAIL.n212 B 0.047454f
C712 VTAIL.n213 B 0.154558f
C713 VTAIL.t9 B 0.420274f
C714 VTAIL.t6 B 0.420274f
C715 VTAIL.n214 B 3.75078f
C716 VTAIL.n215 B 0.409664f
C717 VTAIL.t11 B 0.420274f
C718 VTAIL.t12 B 0.420274f
C719 VTAIL.n216 B 3.75078f
C720 VTAIL.n217 B 0.393572f
C721 VTAIL.n218 B 0.043061f
C722 VTAIL.n219 B 0.028967f
C723 VTAIL.n220 B 0.015566f
C724 VTAIL.n221 B 0.036792f
C725 VTAIL.n222 B 0.016481f
C726 VTAIL.n223 B 0.028967f
C727 VTAIL.n224 B 0.015566f
C728 VTAIL.n225 B 0.036792f
C729 VTAIL.n226 B 0.016481f
C730 VTAIL.n227 B 0.028967f
C731 VTAIL.n228 B 0.016024f
C732 VTAIL.n229 B 0.036792f
C733 VTAIL.n230 B 0.015566f
C734 VTAIL.n231 B 0.016481f
C735 VTAIL.n232 B 0.028967f
C736 VTAIL.n233 B 0.015566f
C737 VTAIL.n234 B 0.036792f
C738 VTAIL.n235 B 0.016481f
C739 VTAIL.n236 B 0.028967f
C740 VTAIL.n237 B 0.015566f
C741 VTAIL.n238 B 0.036792f
C742 VTAIL.n239 B 0.016481f
C743 VTAIL.n240 B 0.028967f
C744 VTAIL.n241 B 0.015566f
C745 VTAIL.n242 B 0.036792f
C746 VTAIL.n243 B 0.016481f
C747 VTAIL.n244 B 0.028967f
C748 VTAIL.n245 B 0.015566f
C749 VTAIL.n246 B 0.036792f
C750 VTAIL.n247 B 0.016481f
C751 VTAIL.n248 B 0.028967f
C752 VTAIL.n249 B 0.015566f
C753 VTAIL.n250 B 0.027594f
C754 VTAIL.n251 B 0.021734f
C755 VTAIL.t13 B 0.060999f
C756 VTAIL.n252 B 0.213333f
C757 VTAIL.n253 B 2.33071f
C758 VTAIL.n254 B 0.015566f
C759 VTAIL.n255 B 0.016481f
C760 VTAIL.n256 B 0.036792f
C761 VTAIL.n257 B 0.036792f
C762 VTAIL.n258 B 0.016481f
C763 VTAIL.n259 B 0.015566f
C764 VTAIL.n260 B 0.028967f
C765 VTAIL.n261 B 0.028967f
C766 VTAIL.n262 B 0.015566f
C767 VTAIL.n263 B 0.016481f
C768 VTAIL.n264 B 0.036792f
C769 VTAIL.n265 B 0.036792f
C770 VTAIL.n266 B 0.016481f
C771 VTAIL.n267 B 0.015566f
C772 VTAIL.n268 B 0.028967f
C773 VTAIL.n269 B 0.028967f
C774 VTAIL.n270 B 0.015566f
C775 VTAIL.n271 B 0.016481f
C776 VTAIL.n272 B 0.036792f
C777 VTAIL.n273 B 0.036792f
C778 VTAIL.n274 B 0.016481f
C779 VTAIL.n275 B 0.015566f
C780 VTAIL.n276 B 0.028967f
C781 VTAIL.n277 B 0.028967f
C782 VTAIL.n278 B 0.015566f
C783 VTAIL.n279 B 0.016481f
C784 VTAIL.n280 B 0.036792f
C785 VTAIL.n281 B 0.036792f
C786 VTAIL.n282 B 0.016481f
C787 VTAIL.n283 B 0.015566f
C788 VTAIL.n284 B 0.028967f
C789 VTAIL.n285 B 0.028967f
C790 VTAIL.n286 B 0.015566f
C791 VTAIL.n287 B 0.016481f
C792 VTAIL.n288 B 0.036792f
C793 VTAIL.n289 B 0.036792f
C794 VTAIL.n290 B 0.016481f
C795 VTAIL.n291 B 0.015566f
C796 VTAIL.n292 B 0.028967f
C797 VTAIL.n293 B 0.028967f
C798 VTAIL.n294 B 0.015566f
C799 VTAIL.n295 B 0.016481f
C800 VTAIL.n296 B 0.036792f
C801 VTAIL.n297 B 0.036792f
C802 VTAIL.n298 B 0.036792f
C803 VTAIL.n299 B 0.016024f
C804 VTAIL.n300 B 0.015566f
C805 VTAIL.n301 B 0.028967f
C806 VTAIL.n302 B 0.028967f
C807 VTAIL.n303 B 0.015566f
C808 VTAIL.n304 B 0.016481f
C809 VTAIL.n305 B 0.036792f
C810 VTAIL.n306 B 0.036792f
C811 VTAIL.n307 B 0.016481f
C812 VTAIL.n308 B 0.015566f
C813 VTAIL.n309 B 0.028967f
C814 VTAIL.n310 B 0.028967f
C815 VTAIL.n311 B 0.015566f
C816 VTAIL.n312 B 0.016481f
C817 VTAIL.n313 B 0.036792f
C818 VTAIL.n314 B 0.083795f
C819 VTAIL.n315 B 0.016481f
C820 VTAIL.n316 B 0.015566f
C821 VTAIL.n317 B 0.071705f
C822 VTAIL.n318 B 0.047454f
C823 VTAIL.n319 B 2.00928f
C824 VTAIL.n320 B 0.043061f
C825 VTAIL.n321 B 0.028967f
C826 VTAIL.n322 B 0.015566f
C827 VTAIL.n323 B 0.036792f
C828 VTAIL.n324 B 0.016481f
C829 VTAIL.n325 B 0.028967f
C830 VTAIL.n326 B 0.015566f
C831 VTAIL.n327 B 0.036792f
C832 VTAIL.n328 B 0.016481f
C833 VTAIL.n329 B 0.028967f
C834 VTAIL.n330 B 0.016024f
C835 VTAIL.n331 B 0.036792f
C836 VTAIL.n332 B 0.016481f
C837 VTAIL.n333 B 0.028967f
C838 VTAIL.n334 B 0.015566f
C839 VTAIL.n335 B 0.036792f
C840 VTAIL.n336 B 0.016481f
C841 VTAIL.n337 B 0.028967f
C842 VTAIL.n338 B 0.015566f
C843 VTAIL.n339 B 0.036792f
C844 VTAIL.n340 B 0.016481f
C845 VTAIL.n341 B 0.028967f
C846 VTAIL.n342 B 0.015566f
C847 VTAIL.n343 B 0.036792f
C848 VTAIL.n344 B 0.016481f
C849 VTAIL.n345 B 0.028967f
C850 VTAIL.n346 B 0.015566f
C851 VTAIL.n347 B 0.036792f
C852 VTAIL.n348 B 0.016481f
C853 VTAIL.n349 B 0.028967f
C854 VTAIL.n350 B 0.015566f
C855 VTAIL.n351 B 0.027594f
C856 VTAIL.n352 B 0.021734f
C857 VTAIL.t16 B 0.060999f
C858 VTAIL.n353 B 0.213333f
C859 VTAIL.n354 B 2.33071f
C860 VTAIL.n355 B 0.015566f
C861 VTAIL.n356 B 0.016481f
C862 VTAIL.n357 B 0.036792f
C863 VTAIL.n358 B 0.036792f
C864 VTAIL.n359 B 0.016481f
C865 VTAIL.n360 B 0.015566f
C866 VTAIL.n361 B 0.028967f
C867 VTAIL.n362 B 0.028967f
C868 VTAIL.n363 B 0.015566f
C869 VTAIL.n364 B 0.016481f
C870 VTAIL.n365 B 0.036792f
C871 VTAIL.n366 B 0.036792f
C872 VTAIL.n367 B 0.016481f
C873 VTAIL.n368 B 0.015566f
C874 VTAIL.n369 B 0.028967f
C875 VTAIL.n370 B 0.028967f
C876 VTAIL.n371 B 0.015566f
C877 VTAIL.n372 B 0.016481f
C878 VTAIL.n373 B 0.036792f
C879 VTAIL.n374 B 0.036792f
C880 VTAIL.n375 B 0.016481f
C881 VTAIL.n376 B 0.015566f
C882 VTAIL.n377 B 0.028967f
C883 VTAIL.n378 B 0.028967f
C884 VTAIL.n379 B 0.015566f
C885 VTAIL.n380 B 0.016481f
C886 VTAIL.n381 B 0.036792f
C887 VTAIL.n382 B 0.036792f
C888 VTAIL.n383 B 0.016481f
C889 VTAIL.n384 B 0.015566f
C890 VTAIL.n385 B 0.028967f
C891 VTAIL.n386 B 0.028967f
C892 VTAIL.n387 B 0.015566f
C893 VTAIL.n388 B 0.016481f
C894 VTAIL.n389 B 0.036792f
C895 VTAIL.n390 B 0.036792f
C896 VTAIL.n391 B 0.016481f
C897 VTAIL.n392 B 0.015566f
C898 VTAIL.n393 B 0.028967f
C899 VTAIL.n394 B 0.028967f
C900 VTAIL.n395 B 0.015566f
C901 VTAIL.n396 B 0.015566f
C902 VTAIL.n397 B 0.016481f
C903 VTAIL.n398 B 0.036792f
C904 VTAIL.n399 B 0.036792f
C905 VTAIL.n400 B 0.036792f
C906 VTAIL.n401 B 0.016024f
C907 VTAIL.n402 B 0.015566f
C908 VTAIL.n403 B 0.028967f
C909 VTAIL.n404 B 0.028967f
C910 VTAIL.n405 B 0.015566f
C911 VTAIL.n406 B 0.016481f
C912 VTAIL.n407 B 0.036792f
C913 VTAIL.n408 B 0.036792f
C914 VTAIL.n409 B 0.016481f
C915 VTAIL.n410 B 0.015566f
C916 VTAIL.n411 B 0.028967f
C917 VTAIL.n412 B 0.028967f
C918 VTAIL.n413 B 0.015566f
C919 VTAIL.n414 B 0.016481f
C920 VTAIL.n415 B 0.036792f
C921 VTAIL.n416 B 0.083795f
C922 VTAIL.n417 B 0.016481f
C923 VTAIL.n418 B 0.015566f
C924 VTAIL.n419 B 0.071705f
C925 VTAIL.n420 B 0.047454f
C926 VTAIL.n421 B 2.00928f
C927 VTAIL.t1 B 0.420274f
C928 VTAIL.t0 B 0.420274f
C929 VTAIL.n422 B 3.75076f
C930 VTAIL.n423 B 0.346516f
C931 VP.n0 B 0.052457f
C932 VP.t2 B 0.982787f
C933 VP.n1 B 0.368817f
C934 VP.n2 B 0.052457f
C935 VP.n3 B 0.052457f
C936 VP.t9 B 0.982787f
C937 VP.t6 B 0.982787f
C938 VP.t0 B 0.982787f
C939 VP.n4 B 0.368817f
C940 VP.t4 B 0.988596f
C941 VP.n5 B 0.370743f
C942 VP.t7 B 0.982787f
C943 VP.n6 B 0.384602f
C944 VP.n7 B 0.011904f
C945 VP.n8 B 0.160894f
C946 VP.n9 B 0.052457f
C947 VP.n10 B 0.011904f
C948 VP.n11 B 0.384602f
C949 VP.n12 B 0.376193f
C950 VP.n13 B 2.485f
C951 VP.n14 B 2.52636f
C952 VP.t3 B 0.982787f
C953 VP.n15 B 0.376193f
C954 VP.t8 B 0.982787f
C955 VP.n16 B 0.384602f
C956 VP.n17 B 0.011904f
C957 VP.n18 B 0.052457f
C958 VP.n19 B 0.052457f
C959 VP.n20 B 0.011904f
C960 VP.t1 B 0.982787f
C961 VP.n21 B 0.384602f
C962 VP.t5 B 0.982787f
C963 VP.n22 B 0.376193f
C964 VP.n23 B 0.040652f
.ends

