* NGSPICE file created from diff_pair_sample_1205.ext - technology: sky130A

.subckt diff_pair_sample_1205 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=0 ps=0 w=8.17 l=3.16
X1 VDD1.t5 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=3.1863 ps=17.12 w=8.17 l=3.16
X2 VTAIL.t2 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=1.34805 ps=8.5 w=8.17 l=3.16
X3 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=1.34805 ps=8.5 w=8.17 l=3.16
X4 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=1.34805 ps=8.5 w=8.17 l=3.16
X5 VDD1.t4 VP.t1 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=1.34805 ps=8.5 w=8.17 l=3.16
X6 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=3.1863 ps=17.12 w=8.17 l=3.16
X7 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=0 ps=0 w=8.17 l=3.16
X8 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=3.1863 ps=17.12 w=8.17 l=3.16
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=0 ps=0 w=8.17 l=3.16
X10 VTAIL.t7 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=1.34805 ps=8.5 w=8.17 l=3.16
X11 VTAIL.t10 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=1.34805 ps=8.5 w=8.17 l=3.16
X12 VDD1.t1 VP.t4 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.34805 pd=8.5 as=3.1863 ps=17.12 w=8.17 l=3.16
X13 VDD1.t0 VP.t5 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=1.34805 ps=8.5 w=8.17 l=3.16
X14 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=1.34805 ps=8.5 w=8.17 l=3.16
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1863 pd=17.12 as=0 ps=0 w=8.17 l=3.16
R0 B.n754 B.n753 585
R1 B.n268 B.n125 585
R2 B.n267 B.n266 585
R3 B.n265 B.n264 585
R4 B.n263 B.n262 585
R5 B.n261 B.n260 585
R6 B.n259 B.n258 585
R7 B.n257 B.n256 585
R8 B.n255 B.n254 585
R9 B.n253 B.n252 585
R10 B.n251 B.n250 585
R11 B.n249 B.n248 585
R12 B.n247 B.n246 585
R13 B.n245 B.n244 585
R14 B.n243 B.n242 585
R15 B.n241 B.n240 585
R16 B.n239 B.n238 585
R17 B.n237 B.n236 585
R18 B.n235 B.n234 585
R19 B.n233 B.n232 585
R20 B.n231 B.n230 585
R21 B.n229 B.n228 585
R22 B.n227 B.n226 585
R23 B.n225 B.n224 585
R24 B.n223 B.n222 585
R25 B.n221 B.n220 585
R26 B.n219 B.n218 585
R27 B.n217 B.n216 585
R28 B.n215 B.n214 585
R29 B.n213 B.n212 585
R30 B.n211 B.n210 585
R31 B.n209 B.n208 585
R32 B.n207 B.n206 585
R33 B.n205 B.n204 585
R34 B.n203 B.n202 585
R35 B.n201 B.n200 585
R36 B.n199 B.n198 585
R37 B.n197 B.n196 585
R38 B.n195 B.n194 585
R39 B.n193 B.n192 585
R40 B.n191 B.n190 585
R41 B.n189 B.n188 585
R42 B.n187 B.n186 585
R43 B.n185 B.n184 585
R44 B.n183 B.n182 585
R45 B.n181 B.n180 585
R46 B.n179 B.n178 585
R47 B.n177 B.n176 585
R48 B.n175 B.n174 585
R49 B.n173 B.n172 585
R50 B.n171 B.n170 585
R51 B.n169 B.n168 585
R52 B.n167 B.n166 585
R53 B.n165 B.n164 585
R54 B.n163 B.n162 585
R55 B.n161 B.n160 585
R56 B.n159 B.n158 585
R57 B.n157 B.n156 585
R58 B.n155 B.n154 585
R59 B.n153 B.n152 585
R60 B.n151 B.n150 585
R61 B.n149 B.n148 585
R62 B.n147 B.n146 585
R63 B.n145 B.n144 585
R64 B.n143 B.n142 585
R65 B.n141 B.n140 585
R66 B.n139 B.n138 585
R67 B.n137 B.n136 585
R68 B.n135 B.n134 585
R69 B.n133 B.n132 585
R70 B.n752 B.n90 585
R71 B.n757 B.n90 585
R72 B.n751 B.n89 585
R73 B.n758 B.n89 585
R74 B.n750 B.n749 585
R75 B.n749 B.n85 585
R76 B.n748 B.n84 585
R77 B.n764 B.n84 585
R78 B.n747 B.n83 585
R79 B.n765 B.n83 585
R80 B.n746 B.n82 585
R81 B.n766 B.n82 585
R82 B.n745 B.n744 585
R83 B.n744 B.n78 585
R84 B.n743 B.n77 585
R85 B.n772 B.n77 585
R86 B.n742 B.n76 585
R87 B.n773 B.n76 585
R88 B.n741 B.n75 585
R89 B.n774 B.n75 585
R90 B.n740 B.n739 585
R91 B.n739 B.n71 585
R92 B.n738 B.n70 585
R93 B.n780 B.n70 585
R94 B.n737 B.n69 585
R95 B.n781 B.n69 585
R96 B.n736 B.n68 585
R97 B.n782 B.n68 585
R98 B.n735 B.n734 585
R99 B.n734 B.n64 585
R100 B.n733 B.n63 585
R101 B.n788 B.n63 585
R102 B.n732 B.n62 585
R103 B.n789 B.n62 585
R104 B.n731 B.n61 585
R105 B.n790 B.n61 585
R106 B.n730 B.n729 585
R107 B.n729 B.n57 585
R108 B.n728 B.n56 585
R109 B.n796 B.n56 585
R110 B.n727 B.n55 585
R111 B.n797 B.n55 585
R112 B.n726 B.n54 585
R113 B.n798 B.n54 585
R114 B.n725 B.n724 585
R115 B.n724 B.n50 585
R116 B.n723 B.n49 585
R117 B.n804 B.n49 585
R118 B.n722 B.n48 585
R119 B.n805 B.n48 585
R120 B.n721 B.n47 585
R121 B.n806 B.n47 585
R122 B.n720 B.n719 585
R123 B.n719 B.n43 585
R124 B.n718 B.n42 585
R125 B.n812 B.n42 585
R126 B.n717 B.n41 585
R127 B.n813 B.n41 585
R128 B.n716 B.n40 585
R129 B.n814 B.n40 585
R130 B.n715 B.n714 585
R131 B.n714 B.n36 585
R132 B.n713 B.n35 585
R133 B.n820 B.n35 585
R134 B.n712 B.n34 585
R135 B.t3 B.n34 585
R136 B.n711 B.n33 585
R137 B.n821 B.n33 585
R138 B.n710 B.n709 585
R139 B.n709 B.n29 585
R140 B.n708 B.n28 585
R141 B.n827 B.n28 585
R142 B.n707 B.n27 585
R143 B.n828 B.n27 585
R144 B.n706 B.n26 585
R145 B.n829 B.n26 585
R146 B.n705 B.n704 585
R147 B.n704 B.n22 585
R148 B.n703 B.n21 585
R149 B.n835 B.n21 585
R150 B.n702 B.n20 585
R151 B.n836 B.n20 585
R152 B.n701 B.n19 585
R153 B.n837 B.n19 585
R154 B.n700 B.n699 585
R155 B.n699 B.n18 585
R156 B.n698 B.n14 585
R157 B.n843 B.n14 585
R158 B.n697 B.n13 585
R159 B.n844 B.n13 585
R160 B.n696 B.n12 585
R161 B.n845 B.n12 585
R162 B.n695 B.n694 585
R163 B.n694 B.n8 585
R164 B.n693 B.n7 585
R165 B.n851 B.n7 585
R166 B.n692 B.n6 585
R167 B.n852 B.n6 585
R168 B.n691 B.n5 585
R169 B.n853 B.n5 585
R170 B.n690 B.n689 585
R171 B.n689 B.n4 585
R172 B.n688 B.n269 585
R173 B.n688 B.n687 585
R174 B.n678 B.n270 585
R175 B.n271 B.n270 585
R176 B.n680 B.n679 585
R177 B.n681 B.n680 585
R178 B.n677 B.n276 585
R179 B.n276 B.n275 585
R180 B.n676 B.n675 585
R181 B.n675 B.n674 585
R182 B.n278 B.n277 585
R183 B.n667 B.n278 585
R184 B.n666 B.n665 585
R185 B.n668 B.n666 585
R186 B.n664 B.n283 585
R187 B.n283 B.n282 585
R188 B.n663 B.n662 585
R189 B.n662 B.n661 585
R190 B.n285 B.n284 585
R191 B.n286 B.n285 585
R192 B.n654 B.n653 585
R193 B.n655 B.n654 585
R194 B.n652 B.n291 585
R195 B.n291 B.n290 585
R196 B.n651 B.n650 585
R197 B.n650 B.n649 585
R198 B.n293 B.n292 585
R199 B.n294 B.n293 585
R200 B.n642 B.n641 585
R201 B.n643 B.n642 585
R202 B.n640 B.n298 585
R203 B.n298 B.t2 585
R204 B.n639 B.n638 585
R205 B.n638 B.n637 585
R206 B.n300 B.n299 585
R207 B.n301 B.n300 585
R208 B.n630 B.n629 585
R209 B.n631 B.n630 585
R210 B.n628 B.n306 585
R211 B.n306 B.n305 585
R212 B.n627 B.n626 585
R213 B.n626 B.n625 585
R214 B.n308 B.n307 585
R215 B.n309 B.n308 585
R216 B.n618 B.n617 585
R217 B.n619 B.n618 585
R218 B.n616 B.n314 585
R219 B.n314 B.n313 585
R220 B.n615 B.n614 585
R221 B.n614 B.n613 585
R222 B.n316 B.n315 585
R223 B.n317 B.n316 585
R224 B.n606 B.n605 585
R225 B.n607 B.n606 585
R226 B.n604 B.n322 585
R227 B.n322 B.n321 585
R228 B.n603 B.n602 585
R229 B.n602 B.n601 585
R230 B.n324 B.n323 585
R231 B.n325 B.n324 585
R232 B.n594 B.n593 585
R233 B.n595 B.n594 585
R234 B.n592 B.n330 585
R235 B.n330 B.n329 585
R236 B.n591 B.n590 585
R237 B.n590 B.n589 585
R238 B.n332 B.n331 585
R239 B.n333 B.n332 585
R240 B.n582 B.n581 585
R241 B.n583 B.n582 585
R242 B.n580 B.n338 585
R243 B.n338 B.n337 585
R244 B.n579 B.n578 585
R245 B.n578 B.n577 585
R246 B.n340 B.n339 585
R247 B.n341 B.n340 585
R248 B.n570 B.n569 585
R249 B.n571 B.n570 585
R250 B.n568 B.n345 585
R251 B.n349 B.n345 585
R252 B.n567 B.n566 585
R253 B.n566 B.n565 585
R254 B.n347 B.n346 585
R255 B.n348 B.n347 585
R256 B.n558 B.n557 585
R257 B.n559 B.n558 585
R258 B.n556 B.n354 585
R259 B.n354 B.n353 585
R260 B.n555 B.n554 585
R261 B.n554 B.n553 585
R262 B.n356 B.n355 585
R263 B.n357 B.n356 585
R264 B.n546 B.n545 585
R265 B.n547 B.n546 585
R266 B.n544 B.n362 585
R267 B.n362 B.n361 585
R268 B.n539 B.n538 585
R269 B.n537 B.n399 585
R270 B.n536 B.n398 585
R271 B.n541 B.n398 585
R272 B.n535 B.n534 585
R273 B.n533 B.n532 585
R274 B.n531 B.n530 585
R275 B.n529 B.n528 585
R276 B.n527 B.n526 585
R277 B.n525 B.n524 585
R278 B.n523 B.n522 585
R279 B.n521 B.n520 585
R280 B.n519 B.n518 585
R281 B.n517 B.n516 585
R282 B.n515 B.n514 585
R283 B.n513 B.n512 585
R284 B.n511 B.n510 585
R285 B.n509 B.n508 585
R286 B.n507 B.n506 585
R287 B.n505 B.n504 585
R288 B.n503 B.n502 585
R289 B.n501 B.n500 585
R290 B.n499 B.n498 585
R291 B.n497 B.n496 585
R292 B.n495 B.n494 585
R293 B.n493 B.n492 585
R294 B.n491 B.n490 585
R295 B.n489 B.n488 585
R296 B.n487 B.n486 585
R297 B.n485 B.n484 585
R298 B.n483 B.n482 585
R299 B.n480 B.n479 585
R300 B.n478 B.n477 585
R301 B.n476 B.n475 585
R302 B.n474 B.n473 585
R303 B.n472 B.n471 585
R304 B.n470 B.n469 585
R305 B.n468 B.n467 585
R306 B.n466 B.n465 585
R307 B.n464 B.n463 585
R308 B.n462 B.n461 585
R309 B.n459 B.n458 585
R310 B.n457 B.n456 585
R311 B.n455 B.n454 585
R312 B.n453 B.n452 585
R313 B.n451 B.n450 585
R314 B.n449 B.n448 585
R315 B.n447 B.n446 585
R316 B.n445 B.n444 585
R317 B.n443 B.n442 585
R318 B.n441 B.n440 585
R319 B.n439 B.n438 585
R320 B.n437 B.n436 585
R321 B.n435 B.n434 585
R322 B.n433 B.n432 585
R323 B.n431 B.n430 585
R324 B.n429 B.n428 585
R325 B.n427 B.n426 585
R326 B.n425 B.n424 585
R327 B.n423 B.n422 585
R328 B.n421 B.n420 585
R329 B.n419 B.n418 585
R330 B.n417 B.n416 585
R331 B.n415 B.n414 585
R332 B.n413 B.n412 585
R333 B.n411 B.n410 585
R334 B.n409 B.n408 585
R335 B.n407 B.n406 585
R336 B.n405 B.n404 585
R337 B.n364 B.n363 585
R338 B.n543 B.n542 585
R339 B.n542 B.n541 585
R340 B.n360 B.n359 585
R341 B.n361 B.n360 585
R342 B.n549 B.n548 585
R343 B.n548 B.n547 585
R344 B.n550 B.n358 585
R345 B.n358 B.n357 585
R346 B.n552 B.n551 585
R347 B.n553 B.n552 585
R348 B.n352 B.n351 585
R349 B.n353 B.n352 585
R350 B.n561 B.n560 585
R351 B.n560 B.n559 585
R352 B.n562 B.n350 585
R353 B.n350 B.n348 585
R354 B.n564 B.n563 585
R355 B.n565 B.n564 585
R356 B.n344 B.n343 585
R357 B.n349 B.n344 585
R358 B.n573 B.n572 585
R359 B.n572 B.n571 585
R360 B.n574 B.n342 585
R361 B.n342 B.n341 585
R362 B.n576 B.n575 585
R363 B.n577 B.n576 585
R364 B.n336 B.n335 585
R365 B.n337 B.n336 585
R366 B.n585 B.n584 585
R367 B.n584 B.n583 585
R368 B.n586 B.n334 585
R369 B.n334 B.n333 585
R370 B.n588 B.n587 585
R371 B.n589 B.n588 585
R372 B.n328 B.n327 585
R373 B.n329 B.n328 585
R374 B.n597 B.n596 585
R375 B.n596 B.n595 585
R376 B.n598 B.n326 585
R377 B.n326 B.n325 585
R378 B.n600 B.n599 585
R379 B.n601 B.n600 585
R380 B.n320 B.n319 585
R381 B.n321 B.n320 585
R382 B.n609 B.n608 585
R383 B.n608 B.n607 585
R384 B.n610 B.n318 585
R385 B.n318 B.n317 585
R386 B.n612 B.n611 585
R387 B.n613 B.n612 585
R388 B.n312 B.n311 585
R389 B.n313 B.n312 585
R390 B.n621 B.n620 585
R391 B.n620 B.n619 585
R392 B.n622 B.n310 585
R393 B.n310 B.n309 585
R394 B.n624 B.n623 585
R395 B.n625 B.n624 585
R396 B.n304 B.n303 585
R397 B.n305 B.n304 585
R398 B.n633 B.n632 585
R399 B.n632 B.n631 585
R400 B.n634 B.n302 585
R401 B.n302 B.n301 585
R402 B.n636 B.n635 585
R403 B.n637 B.n636 585
R404 B.n297 B.n296 585
R405 B.t2 B.n297 585
R406 B.n645 B.n644 585
R407 B.n644 B.n643 585
R408 B.n646 B.n295 585
R409 B.n295 B.n294 585
R410 B.n648 B.n647 585
R411 B.n649 B.n648 585
R412 B.n289 B.n288 585
R413 B.n290 B.n289 585
R414 B.n657 B.n656 585
R415 B.n656 B.n655 585
R416 B.n658 B.n287 585
R417 B.n287 B.n286 585
R418 B.n660 B.n659 585
R419 B.n661 B.n660 585
R420 B.n281 B.n280 585
R421 B.n282 B.n281 585
R422 B.n670 B.n669 585
R423 B.n669 B.n668 585
R424 B.n671 B.n279 585
R425 B.n667 B.n279 585
R426 B.n673 B.n672 585
R427 B.n674 B.n673 585
R428 B.n274 B.n273 585
R429 B.n275 B.n274 585
R430 B.n683 B.n682 585
R431 B.n682 B.n681 585
R432 B.n684 B.n272 585
R433 B.n272 B.n271 585
R434 B.n686 B.n685 585
R435 B.n687 B.n686 585
R436 B.n2 B.n0 585
R437 B.n4 B.n2 585
R438 B.n3 B.n1 585
R439 B.n852 B.n3 585
R440 B.n850 B.n849 585
R441 B.n851 B.n850 585
R442 B.n848 B.n9 585
R443 B.n9 B.n8 585
R444 B.n847 B.n846 585
R445 B.n846 B.n845 585
R446 B.n11 B.n10 585
R447 B.n844 B.n11 585
R448 B.n842 B.n841 585
R449 B.n843 B.n842 585
R450 B.n840 B.n15 585
R451 B.n18 B.n15 585
R452 B.n839 B.n838 585
R453 B.n838 B.n837 585
R454 B.n17 B.n16 585
R455 B.n836 B.n17 585
R456 B.n834 B.n833 585
R457 B.n835 B.n834 585
R458 B.n832 B.n23 585
R459 B.n23 B.n22 585
R460 B.n831 B.n830 585
R461 B.n830 B.n829 585
R462 B.n25 B.n24 585
R463 B.n828 B.n25 585
R464 B.n826 B.n825 585
R465 B.n827 B.n826 585
R466 B.n824 B.n30 585
R467 B.n30 B.n29 585
R468 B.n823 B.n822 585
R469 B.n822 B.n821 585
R470 B.n32 B.n31 585
R471 B.t3 B.n32 585
R472 B.n819 B.n818 585
R473 B.n820 B.n819 585
R474 B.n817 B.n37 585
R475 B.n37 B.n36 585
R476 B.n816 B.n815 585
R477 B.n815 B.n814 585
R478 B.n39 B.n38 585
R479 B.n813 B.n39 585
R480 B.n811 B.n810 585
R481 B.n812 B.n811 585
R482 B.n809 B.n44 585
R483 B.n44 B.n43 585
R484 B.n808 B.n807 585
R485 B.n807 B.n806 585
R486 B.n46 B.n45 585
R487 B.n805 B.n46 585
R488 B.n803 B.n802 585
R489 B.n804 B.n803 585
R490 B.n801 B.n51 585
R491 B.n51 B.n50 585
R492 B.n800 B.n799 585
R493 B.n799 B.n798 585
R494 B.n53 B.n52 585
R495 B.n797 B.n53 585
R496 B.n795 B.n794 585
R497 B.n796 B.n795 585
R498 B.n793 B.n58 585
R499 B.n58 B.n57 585
R500 B.n792 B.n791 585
R501 B.n791 B.n790 585
R502 B.n60 B.n59 585
R503 B.n789 B.n60 585
R504 B.n787 B.n786 585
R505 B.n788 B.n787 585
R506 B.n785 B.n65 585
R507 B.n65 B.n64 585
R508 B.n784 B.n783 585
R509 B.n783 B.n782 585
R510 B.n67 B.n66 585
R511 B.n781 B.n67 585
R512 B.n779 B.n778 585
R513 B.n780 B.n779 585
R514 B.n777 B.n72 585
R515 B.n72 B.n71 585
R516 B.n776 B.n775 585
R517 B.n775 B.n774 585
R518 B.n74 B.n73 585
R519 B.n773 B.n74 585
R520 B.n771 B.n770 585
R521 B.n772 B.n771 585
R522 B.n769 B.n79 585
R523 B.n79 B.n78 585
R524 B.n768 B.n767 585
R525 B.n767 B.n766 585
R526 B.n81 B.n80 585
R527 B.n765 B.n81 585
R528 B.n763 B.n762 585
R529 B.n764 B.n763 585
R530 B.n761 B.n86 585
R531 B.n86 B.n85 585
R532 B.n760 B.n759 585
R533 B.n759 B.n758 585
R534 B.n88 B.n87 585
R535 B.n757 B.n88 585
R536 B.n855 B.n854 585
R537 B.n854 B.n853 585
R538 B.n539 B.n360 550.159
R539 B.n132 B.n88 550.159
R540 B.n542 B.n362 550.159
R541 B.n754 B.n90 550.159
R542 B.n402 B.t14 271.07
R543 B.n400 B.t10 271.07
R544 B.n129 B.t6 271.07
R545 B.n126 B.t17 271.07
R546 B.n756 B.n755 256.663
R547 B.n756 B.n124 256.663
R548 B.n756 B.n123 256.663
R549 B.n756 B.n122 256.663
R550 B.n756 B.n121 256.663
R551 B.n756 B.n120 256.663
R552 B.n756 B.n119 256.663
R553 B.n756 B.n118 256.663
R554 B.n756 B.n117 256.663
R555 B.n756 B.n116 256.663
R556 B.n756 B.n115 256.663
R557 B.n756 B.n114 256.663
R558 B.n756 B.n113 256.663
R559 B.n756 B.n112 256.663
R560 B.n756 B.n111 256.663
R561 B.n756 B.n110 256.663
R562 B.n756 B.n109 256.663
R563 B.n756 B.n108 256.663
R564 B.n756 B.n107 256.663
R565 B.n756 B.n106 256.663
R566 B.n756 B.n105 256.663
R567 B.n756 B.n104 256.663
R568 B.n756 B.n103 256.663
R569 B.n756 B.n102 256.663
R570 B.n756 B.n101 256.663
R571 B.n756 B.n100 256.663
R572 B.n756 B.n99 256.663
R573 B.n756 B.n98 256.663
R574 B.n756 B.n97 256.663
R575 B.n756 B.n96 256.663
R576 B.n756 B.n95 256.663
R577 B.n756 B.n94 256.663
R578 B.n756 B.n93 256.663
R579 B.n756 B.n92 256.663
R580 B.n756 B.n91 256.663
R581 B.n541 B.n540 256.663
R582 B.n541 B.n365 256.663
R583 B.n541 B.n366 256.663
R584 B.n541 B.n367 256.663
R585 B.n541 B.n368 256.663
R586 B.n541 B.n369 256.663
R587 B.n541 B.n370 256.663
R588 B.n541 B.n371 256.663
R589 B.n541 B.n372 256.663
R590 B.n541 B.n373 256.663
R591 B.n541 B.n374 256.663
R592 B.n541 B.n375 256.663
R593 B.n541 B.n376 256.663
R594 B.n541 B.n377 256.663
R595 B.n541 B.n378 256.663
R596 B.n541 B.n379 256.663
R597 B.n541 B.n380 256.663
R598 B.n541 B.n381 256.663
R599 B.n541 B.n382 256.663
R600 B.n541 B.n383 256.663
R601 B.n541 B.n384 256.663
R602 B.n541 B.n385 256.663
R603 B.n541 B.n386 256.663
R604 B.n541 B.n387 256.663
R605 B.n541 B.n388 256.663
R606 B.n541 B.n389 256.663
R607 B.n541 B.n390 256.663
R608 B.n541 B.n391 256.663
R609 B.n541 B.n392 256.663
R610 B.n541 B.n393 256.663
R611 B.n541 B.n394 256.663
R612 B.n541 B.n395 256.663
R613 B.n541 B.n396 256.663
R614 B.n541 B.n397 256.663
R615 B.n548 B.n360 163.367
R616 B.n548 B.n358 163.367
R617 B.n552 B.n358 163.367
R618 B.n552 B.n352 163.367
R619 B.n560 B.n352 163.367
R620 B.n560 B.n350 163.367
R621 B.n564 B.n350 163.367
R622 B.n564 B.n344 163.367
R623 B.n572 B.n344 163.367
R624 B.n572 B.n342 163.367
R625 B.n576 B.n342 163.367
R626 B.n576 B.n336 163.367
R627 B.n584 B.n336 163.367
R628 B.n584 B.n334 163.367
R629 B.n588 B.n334 163.367
R630 B.n588 B.n328 163.367
R631 B.n596 B.n328 163.367
R632 B.n596 B.n326 163.367
R633 B.n600 B.n326 163.367
R634 B.n600 B.n320 163.367
R635 B.n608 B.n320 163.367
R636 B.n608 B.n318 163.367
R637 B.n612 B.n318 163.367
R638 B.n612 B.n312 163.367
R639 B.n620 B.n312 163.367
R640 B.n620 B.n310 163.367
R641 B.n624 B.n310 163.367
R642 B.n624 B.n304 163.367
R643 B.n632 B.n304 163.367
R644 B.n632 B.n302 163.367
R645 B.n636 B.n302 163.367
R646 B.n636 B.n297 163.367
R647 B.n644 B.n297 163.367
R648 B.n644 B.n295 163.367
R649 B.n648 B.n295 163.367
R650 B.n648 B.n289 163.367
R651 B.n656 B.n289 163.367
R652 B.n656 B.n287 163.367
R653 B.n660 B.n287 163.367
R654 B.n660 B.n281 163.367
R655 B.n669 B.n281 163.367
R656 B.n669 B.n279 163.367
R657 B.n673 B.n279 163.367
R658 B.n673 B.n274 163.367
R659 B.n682 B.n274 163.367
R660 B.n682 B.n272 163.367
R661 B.n686 B.n272 163.367
R662 B.n686 B.n2 163.367
R663 B.n854 B.n2 163.367
R664 B.n854 B.n3 163.367
R665 B.n850 B.n3 163.367
R666 B.n850 B.n9 163.367
R667 B.n846 B.n9 163.367
R668 B.n846 B.n11 163.367
R669 B.n842 B.n11 163.367
R670 B.n842 B.n15 163.367
R671 B.n838 B.n15 163.367
R672 B.n838 B.n17 163.367
R673 B.n834 B.n17 163.367
R674 B.n834 B.n23 163.367
R675 B.n830 B.n23 163.367
R676 B.n830 B.n25 163.367
R677 B.n826 B.n25 163.367
R678 B.n826 B.n30 163.367
R679 B.n822 B.n30 163.367
R680 B.n822 B.n32 163.367
R681 B.n819 B.n32 163.367
R682 B.n819 B.n37 163.367
R683 B.n815 B.n37 163.367
R684 B.n815 B.n39 163.367
R685 B.n811 B.n39 163.367
R686 B.n811 B.n44 163.367
R687 B.n807 B.n44 163.367
R688 B.n807 B.n46 163.367
R689 B.n803 B.n46 163.367
R690 B.n803 B.n51 163.367
R691 B.n799 B.n51 163.367
R692 B.n799 B.n53 163.367
R693 B.n795 B.n53 163.367
R694 B.n795 B.n58 163.367
R695 B.n791 B.n58 163.367
R696 B.n791 B.n60 163.367
R697 B.n787 B.n60 163.367
R698 B.n787 B.n65 163.367
R699 B.n783 B.n65 163.367
R700 B.n783 B.n67 163.367
R701 B.n779 B.n67 163.367
R702 B.n779 B.n72 163.367
R703 B.n775 B.n72 163.367
R704 B.n775 B.n74 163.367
R705 B.n771 B.n74 163.367
R706 B.n771 B.n79 163.367
R707 B.n767 B.n79 163.367
R708 B.n767 B.n81 163.367
R709 B.n763 B.n81 163.367
R710 B.n763 B.n86 163.367
R711 B.n759 B.n86 163.367
R712 B.n759 B.n88 163.367
R713 B.n399 B.n398 163.367
R714 B.n534 B.n398 163.367
R715 B.n532 B.n531 163.367
R716 B.n528 B.n527 163.367
R717 B.n524 B.n523 163.367
R718 B.n520 B.n519 163.367
R719 B.n516 B.n515 163.367
R720 B.n512 B.n511 163.367
R721 B.n508 B.n507 163.367
R722 B.n504 B.n503 163.367
R723 B.n500 B.n499 163.367
R724 B.n496 B.n495 163.367
R725 B.n492 B.n491 163.367
R726 B.n488 B.n487 163.367
R727 B.n484 B.n483 163.367
R728 B.n479 B.n478 163.367
R729 B.n475 B.n474 163.367
R730 B.n471 B.n470 163.367
R731 B.n467 B.n466 163.367
R732 B.n463 B.n462 163.367
R733 B.n458 B.n457 163.367
R734 B.n454 B.n453 163.367
R735 B.n450 B.n449 163.367
R736 B.n446 B.n445 163.367
R737 B.n442 B.n441 163.367
R738 B.n438 B.n437 163.367
R739 B.n434 B.n433 163.367
R740 B.n430 B.n429 163.367
R741 B.n426 B.n425 163.367
R742 B.n422 B.n421 163.367
R743 B.n418 B.n417 163.367
R744 B.n414 B.n413 163.367
R745 B.n410 B.n409 163.367
R746 B.n406 B.n405 163.367
R747 B.n542 B.n364 163.367
R748 B.n546 B.n362 163.367
R749 B.n546 B.n356 163.367
R750 B.n554 B.n356 163.367
R751 B.n554 B.n354 163.367
R752 B.n558 B.n354 163.367
R753 B.n558 B.n347 163.367
R754 B.n566 B.n347 163.367
R755 B.n566 B.n345 163.367
R756 B.n570 B.n345 163.367
R757 B.n570 B.n340 163.367
R758 B.n578 B.n340 163.367
R759 B.n578 B.n338 163.367
R760 B.n582 B.n338 163.367
R761 B.n582 B.n332 163.367
R762 B.n590 B.n332 163.367
R763 B.n590 B.n330 163.367
R764 B.n594 B.n330 163.367
R765 B.n594 B.n324 163.367
R766 B.n602 B.n324 163.367
R767 B.n602 B.n322 163.367
R768 B.n606 B.n322 163.367
R769 B.n606 B.n316 163.367
R770 B.n614 B.n316 163.367
R771 B.n614 B.n314 163.367
R772 B.n618 B.n314 163.367
R773 B.n618 B.n308 163.367
R774 B.n626 B.n308 163.367
R775 B.n626 B.n306 163.367
R776 B.n630 B.n306 163.367
R777 B.n630 B.n300 163.367
R778 B.n638 B.n300 163.367
R779 B.n638 B.n298 163.367
R780 B.n642 B.n298 163.367
R781 B.n642 B.n293 163.367
R782 B.n650 B.n293 163.367
R783 B.n650 B.n291 163.367
R784 B.n654 B.n291 163.367
R785 B.n654 B.n285 163.367
R786 B.n662 B.n285 163.367
R787 B.n662 B.n283 163.367
R788 B.n666 B.n283 163.367
R789 B.n666 B.n278 163.367
R790 B.n675 B.n278 163.367
R791 B.n675 B.n276 163.367
R792 B.n680 B.n276 163.367
R793 B.n680 B.n270 163.367
R794 B.n688 B.n270 163.367
R795 B.n689 B.n688 163.367
R796 B.n689 B.n5 163.367
R797 B.n6 B.n5 163.367
R798 B.n7 B.n6 163.367
R799 B.n694 B.n7 163.367
R800 B.n694 B.n12 163.367
R801 B.n13 B.n12 163.367
R802 B.n14 B.n13 163.367
R803 B.n699 B.n14 163.367
R804 B.n699 B.n19 163.367
R805 B.n20 B.n19 163.367
R806 B.n21 B.n20 163.367
R807 B.n704 B.n21 163.367
R808 B.n704 B.n26 163.367
R809 B.n27 B.n26 163.367
R810 B.n28 B.n27 163.367
R811 B.n709 B.n28 163.367
R812 B.n709 B.n33 163.367
R813 B.n34 B.n33 163.367
R814 B.n35 B.n34 163.367
R815 B.n714 B.n35 163.367
R816 B.n714 B.n40 163.367
R817 B.n41 B.n40 163.367
R818 B.n42 B.n41 163.367
R819 B.n719 B.n42 163.367
R820 B.n719 B.n47 163.367
R821 B.n48 B.n47 163.367
R822 B.n49 B.n48 163.367
R823 B.n724 B.n49 163.367
R824 B.n724 B.n54 163.367
R825 B.n55 B.n54 163.367
R826 B.n56 B.n55 163.367
R827 B.n729 B.n56 163.367
R828 B.n729 B.n61 163.367
R829 B.n62 B.n61 163.367
R830 B.n63 B.n62 163.367
R831 B.n734 B.n63 163.367
R832 B.n734 B.n68 163.367
R833 B.n69 B.n68 163.367
R834 B.n70 B.n69 163.367
R835 B.n739 B.n70 163.367
R836 B.n739 B.n75 163.367
R837 B.n76 B.n75 163.367
R838 B.n77 B.n76 163.367
R839 B.n744 B.n77 163.367
R840 B.n744 B.n82 163.367
R841 B.n83 B.n82 163.367
R842 B.n84 B.n83 163.367
R843 B.n749 B.n84 163.367
R844 B.n749 B.n89 163.367
R845 B.n90 B.n89 163.367
R846 B.n136 B.n135 163.367
R847 B.n140 B.n139 163.367
R848 B.n144 B.n143 163.367
R849 B.n148 B.n147 163.367
R850 B.n152 B.n151 163.367
R851 B.n156 B.n155 163.367
R852 B.n160 B.n159 163.367
R853 B.n164 B.n163 163.367
R854 B.n168 B.n167 163.367
R855 B.n172 B.n171 163.367
R856 B.n176 B.n175 163.367
R857 B.n180 B.n179 163.367
R858 B.n184 B.n183 163.367
R859 B.n188 B.n187 163.367
R860 B.n192 B.n191 163.367
R861 B.n196 B.n195 163.367
R862 B.n200 B.n199 163.367
R863 B.n204 B.n203 163.367
R864 B.n208 B.n207 163.367
R865 B.n212 B.n211 163.367
R866 B.n216 B.n215 163.367
R867 B.n220 B.n219 163.367
R868 B.n224 B.n223 163.367
R869 B.n228 B.n227 163.367
R870 B.n232 B.n231 163.367
R871 B.n236 B.n235 163.367
R872 B.n240 B.n239 163.367
R873 B.n244 B.n243 163.367
R874 B.n248 B.n247 163.367
R875 B.n252 B.n251 163.367
R876 B.n256 B.n255 163.367
R877 B.n260 B.n259 163.367
R878 B.n264 B.n263 163.367
R879 B.n266 B.n125 163.367
R880 B.n402 B.t16 136.438
R881 B.n126 B.t18 136.438
R882 B.n400 B.t13 136.428
R883 B.n129 B.t8 136.428
R884 B.n541 B.n361 110.451
R885 B.n757 B.n756 110.451
R886 B.n540 B.n539 71.676
R887 B.n534 B.n365 71.676
R888 B.n531 B.n366 71.676
R889 B.n527 B.n367 71.676
R890 B.n523 B.n368 71.676
R891 B.n519 B.n369 71.676
R892 B.n515 B.n370 71.676
R893 B.n511 B.n371 71.676
R894 B.n507 B.n372 71.676
R895 B.n503 B.n373 71.676
R896 B.n499 B.n374 71.676
R897 B.n495 B.n375 71.676
R898 B.n491 B.n376 71.676
R899 B.n487 B.n377 71.676
R900 B.n483 B.n378 71.676
R901 B.n478 B.n379 71.676
R902 B.n474 B.n380 71.676
R903 B.n470 B.n381 71.676
R904 B.n466 B.n382 71.676
R905 B.n462 B.n383 71.676
R906 B.n457 B.n384 71.676
R907 B.n453 B.n385 71.676
R908 B.n449 B.n386 71.676
R909 B.n445 B.n387 71.676
R910 B.n441 B.n388 71.676
R911 B.n437 B.n389 71.676
R912 B.n433 B.n390 71.676
R913 B.n429 B.n391 71.676
R914 B.n425 B.n392 71.676
R915 B.n421 B.n393 71.676
R916 B.n417 B.n394 71.676
R917 B.n413 B.n395 71.676
R918 B.n409 B.n396 71.676
R919 B.n405 B.n397 71.676
R920 B.n132 B.n91 71.676
R921 B.n136 B.n92 71.676
R922 B.n140 B.n93 71.676
R923 B.n144 B.n94 71.676
R924 B.n148 B.n95 71.676
R925 B.n152 B.n96 71.676
R926 B.n156 B.n97 71.676
R927 B.n160 B.n98 71.676
R928 B.n164 B.n99 71.676
R929 B.n168 B.n100 71.676
R930 B.n172 B.n101 71.676
R931 B.n176 B.n102 71.676
R932 B.n180 B.n103 71.676
R933 B.n184 B.n104 71.676
R934 B.n188 B.n105 71.676
R935 B.n192 B.n106 71.676
R936 B.n196 B.n107 71.676
R937 B.n200 B.n108 71.676
R938 B.n204 B.n109 71.676
R939 B.n208 B.n110 71.676
R940 B.n212 B.n111 71.676
R941 B.n216 B.n112 71.676
R942 B.n220 B.n113 71.676
R943 B.n224 B.n114 71.676
R944 B.n228 B.n115 71.676
R945 B.n232 B.n116 71.676
R946 B.n236 B.n117 71.676
R947 B.n240 B.n118 71.676
R948 B.n244 B.n119 71.676
R949 B.n248 B.n120 71.676
R950 B.n252 B.n121 71.676
R951 B.n256 B.n122 71.676
R952 B.n260 B.n123 71.676
R953 B.n264 B.n124 71.676
R954 B.n755 B.n125 71.676
R955 B.n755 B.n754 71.676
R956 B.n266 B.n124 71.676
R957 B.n263 B.n123 71.676
R958 B.n259 B.n122 71.676
R959 B.n255 B.n121 71.676
R960 B.n251 B.n120 71.676
R961 B.n247 B.n119 71.676
R962 B.n243 B.n118 71.676
R963 B.n239 B.n117 71.676
R964 B.n235 B.n116 71.676
R965 B.n231 B.n115 71.676
R966 B.n227 B.n114 71.676
R967 B.n223 B.n113 71.676
R968 B.n219 B.n112 71.676
R969 B.n215 B.n111 71.676
R970 B.n211 B.n110 71.676
R971 B.n207 B.n109 71.676
R972 B.n203 B.n108 71.676
R973 B.n199 B.n107 71.676
R974 B.n195 B.n106 71.676
R975 B.n191 B.n105 71.676
R976 B.n187 B.n104 71.676
R977 B.n183 B.n103 71.676
R978 B.n179 B.n102 71.676
R979 B.n175 B.n101 71.676
R980 B.n171 B.n100 71.676
R981 B.n167 B.n99 71.676
R982 B.n163 B.n98 71.676
R983 B.n159 B.n97 71.676
R984 B.n155 B.n96 71.676
R985 B.n151 B.n95 71.676
R986 B.n147 B.n94 71.676
R987 B.n143 B.n93 71.676
R988 B.n139 B.n92 71.676
R989 B.n135 B.n91 71.676
R990 B.n540 B.n399 71.676
R991 B.n532 B.n365 71.676
R992 B.n528 B.n366 71.676
R993 B.n524 B.n367 71.676
R994 B.n520 B.n368 71.676
R995 B.n516 B.n369 71.676
R996 B.n512 B.n370 71.676
R997 B.n508 B.n371 71.676
R998 B.n504 B.n372 71.676
R999 B.n500 B.n373 71.676
R1000 B.n496 B.n374 71.676
R1001 B.n492 B.n375 71.676
R1002 B.n488 B.n376 71.676
R1003 B.n484 B.n377 71.676
R1004 B.n479 B.n378 71.676
R1005 B.n475 B.n379 71.676
R1006 B.n471 B.n380 71.676
R1007 B.n467 B.n381 71.676
R1008 B.n463 B.n382 71.676
R1009 B.n458 B.n383 71.676
R1010 B.n454 B.n384 71.676
R1011 B.n450 B.n385 71.676
R1012 B.n446 B.n386 71.676
R1013 B.n442 B.n387 71.676
R1014 B.n438 B.n388 71.676
R1015 B.n434 B.n389 71.676
R1016 B.n430 B.n390 71.676
R1017 B.n426 B.n391 71.676
R1018 B.n422 B.n392 71.676
R1019 B.n418 B.n393 71.676
R1020 B.n414 B.n394 71.676
R1021 B.n410 B.n395 71.676
R1022 B.n406 B.n396 71.676
R1023 B.n397 B.n364 71.676
R1024 B.n403 B.t15 68.7523
R1025 B.n127 B.t19 68.7523
R1026 B.n401 B.t12 68.7426
R1027 B.n130 B.t9 68.7426
R1028 B.n403 B.n402 67.6854
R1029 B.n401 B.n400 67.6854
R1030 B.n130 B.n129 67.6854
R1031 B.n127 B.n126 67.6854
R1032 B.n460 B.n403 59.5399
R1033 B.n481 B.n401 59.5399
R1034 B.n131 B.n130 59.5399
R1035 B.n128 B.n127 59.5399
R1036 B.n547 B.n361 55.6346
R1037 B.n547 B.n357 55.6346
R1038 B.n553 B.n357 55.6346
R1039 B.n553 B.n353 55.6346
R1040 B.n559 B.n353 55.6346
R1041 B.n559 B.n348 55.6346
R1042 B.n565 B.n348 55.6346
R1043 B.n565 B.n349 55.6346
R1044 B.n571 B.n341 55.6346
R1045 B.n577 B.n341 55.6346
R1046 B.n577 B.n337 55.6346
R1047 B.n583 B.n337 55.6346
R1048 B.n583 B.n333 55.6346
R1049 B.n589 B.n333 55.6346
R1050 B.n589 B.n329 55.6346
R1051 B.n595 B.n329 55.6346
R1052 B.n595 B.n325 55.6346
R1053 B.n601 B.n325 55.6346
R1054 B.n601 B.n321 55.6346
R1055 B.n607 B.n321 55.6346
R1056 B.n613 B.n317 55.6346
R1057 B.n613 B.n313 55.6346
R1058 B.n619 B.n313 55.6346
R1059 B.n619 B.n309 55.6346
R1060 B.n625 B.n309 55.6346
R1061 B.n625 B.n305 55.6346
R1062 B.n631 B.n305 55.6346
R1063 B.n631 B.n301 55.6346
R1064 B.n637 B.n301 55.6346
R1065 B.n637 B.t2 55.6346
R1066 B.n643 B.t2 55.6346
R1067 B.n643 B.n294 55.6346
R1068 B.n649 B.n294 55.6346
R1069 B.n649 B.n290 55.6346
R1070 B.n655 B.n290 55.6346
R1071 B.n655 B.n286 55.6346
R1072 B.n661 B.n286 55.6346
R1073 B.n661 B.n282 55.6346
R1074 B.n668 B.n282 55.6346
R1075 B.n668 B.n667 55.6346
R1076 B.n674 B.n275 55.6346
R1077 B.n681 B.n275 55.6346
R1078 B.n681 B.n271 55.6346
R1079 B.n687 B.n271 55.6346
R1080 B.n687 B.n4 55.6346
R1081 B.n853 B.n4 55.6346
R1082 B.n853 B.n852 55.6346
R1083 B.n852 B.n851 55.6346
R1084 B.n851 B.n8 55.6346
R1085 B.n845 B.n8 55.6346
R1086 B.n845 B.n844 55.6346
R1087 B.n844 B.n843 55.6346
R1088 B.n837 B.n18 55.6346
R1089 B.n837 B.n836 55.6346
R1090 B.n836 B.n835 55.6346
R1091 B.n835 B.n22 55.6346
R1092 B.n829 B.n22 55.6346
R1093 B.n829 B.n828 55.6346
R1094 B.n828 B.n827 55.6346
R1095 B.n827 B.n29 55.6346
R1096 B.n821 B.n29 55.6346
R1097 B.n821 B.t3 55.6346
R1098 B.t3 B.n820 55.6346
R1099 B.n820 B.n36 55.6346
R1100 B.n814 B.n36 55.6346
R1101 B.n814 B.n813 55.6346
R1102 B.n813 B.n812 55.6346
R1103 B.n812 B.n43 55.6346
R1104 B.n806 B.n43 55.6346
R1105 B.n806 B.n805 55.6346
R1106 B.n805 B.n804 55.6346
R1107 B.n804 B.n50 55.6346
R1108 B.n798 B.n797 55.6346
R1109 B.n797 B.n796 55.6346
R1110 B.n796 B.n57 55.6346
R1111 B.n790 B.n57 55.6346
R1112 B.n790 B.n789 55.6346
R1113 B.n789 B.n788 55.6346
R1114 B.n788 B.n64 55.6346
R1115 B.n782 B.n64 55.6346
R1116 B.n782 B.n781 55.6346
R1117 B.n781 B.n780 55.6346
R1118 B.n780 B.n71 55.6346
R1119 B.n774 B.n71 55.6346
R1120 B.n773 B.n772 55.6346
R1121 B.n772 B.n78 55.6346
R1122 B.n766 B.n78 55.6346
R1123 B.n766 B.n765 55.6346
R1124 B.n765 B.n764 55.6346
R1125 B.n764 B.n85 55.6346
R1126 B.n758 B.n85 55.6346
R1127 B.n758 B.n757 55.6346
R1128 B.n571 B.t11 40.9079
R1129 B.n607 B.t1 40.9079
R1130 B.n674 B.t4 40.9079
R1131 B.n843 B.t5 40.9079
R1132 B.n798 B.t0 40.9079
R1133 B.n774 B.t7 40.9079
R1134 B.n133 B.n87 35.7468
R1135 B.n753 B.n752 35.7468
R1136 B.n544 B.n543 35.7468
R1137 B.n538 B.n359 35.7468
R1138 B B.n855 18.0485
R1139 B.n349 B.t11 14.7272
R1140 B.t1 B.n317 14.7272
R1141 B.n667 B.t4 14.7272
R1142 B.n18 B.t5 14.7272
R1143 B.t0 B.n50 14.7272
R1144 B.t7 B.n773 14.7272
R1145 B.n134 B.n133 10.6151
R1146 B.n137 B.n134 10.6151
R1147 B.n138 B.n137 10.6151
R1148 B.n141 B.n138 10.6151
R1149 B.n142 B.n141 10.6151
R1150 B.n145 B.n142 10.6151
R1151 B.n146 B.n145 10.6151
R1152 B.n149 B.n146 10.6151
R1153 B.n150 B.n149 10.6151
R1154 B.n153 B.n150 10.6151
R1155 B.n154 B.n153 10.6151
R1156 B.n157 B.n154 10.6151
R1157 B.n158 B.n157 10.6151
R1158 B.n161 B.n158 10.6151
R1159 B.n162 B.n161 10.6151
R1160 B.n165 B.n162 10.6151
R1161 B.n166 B.n165 10.6151
R1162 B.n169 B.n166 10.6151
R1163 B.n170 B.n169 10.6151
R1164 B.n173 B.n170 10.6151
R1165 B.n174 B.n173 10.6151
R1166 B.n177 B.n174 10.6151
R1167 B.n178 B.n177 10.6151
R1168 B.n181 B.n178 10.6151
R1169 B.n182 B.n181 10.6151
R1170 B.n185 B.n182 10.6151
R1171 B.n186 B.n185 10.6151
R1172 B.n189 B.n186 10.6151
R1173 B.n190 B.n189 10.6151
R1174 B.n194 B.n193 10.6151
R1175 B.n197 B.n194 10.6151
R1176 B.n198 B.n197 10.6151
R1177 B.n201 B.n198 10.6151
R1178 B.n202 B.n201 10.6151
R1179 B.n205 B.n202 10.6151
R1180 B.n206 B.n205 10.6151
R1181 B.n209 B.n206 10.6151
R1182 B.n210 B.n209 10.6151
R1183 B.n214 B.n213 10.6151
R1184 B.n217 B.n214 10.6151
R1185 B.n218 B.n217 10.6151
R1186 B.n221 B.n218 10.6151
R1187 B.n222 B.n221 10.6151
R1188 B.n225 B.n222 10.6151
R1189 B.n226 B.n225 10.6151
R1190 B.n229 B.n226 10.6151
R1191 B.n230 B.n229 10.6151
R1192 B.n233 B.n230 10.6151
R1193 B.n234 B.n233 10.6151
R1194 B.n237 B.n234 10.6151
R1195 B.n238 B.n237 10.6151
R1196 B.n241 B.n238 10.6151
R1197 B.n242 B.n241 10.6151
R1198 B.n245 B.n242 10.6151
R1199 B.n246 B.n245 10.6151
R1200 B.n249 B.n246 10.6151
R1201 B.n250 B.n249 10.6151
R1202 B.n253 B.n250 10.6151
R1203 B.n254 B.n253 10.6151
R1204 B.n257 B.n254 10.6151
R1205 B.n258 B.n257 10.6151
R1206 B.n261 B.n258 10.6151
R1207 B.n262 B.n261 10.6151
R1208 B.n265 B.n262 10.6151
R1209 B.n267 B.n265 10.6151
R1210 B.n268 B.n267 10.6151
R1211 B.n753 B.n268 10.6151
R1212 B.n545 B.n544 10.6151
R1213 B.n545 B.n355 10.6151
R1214 B.n555 B.n355 10.6151
R1215 B.n556 B.n555 10.6151
R1216 B.n557 B.n556 10.6151
R1217 B.n557 B.n346 10.6151
R1218 B.n567 B.n346 10.6151
R1219 B.n568 B.n567 10.6151
R1220 B.n569 B.n568 10.6151
R1221 B.n569 B.n339 10.6151
R1222 B.n579 B.n339 10.6151
R1223 B.n580 B.n579 10.6151
R1224 B.n581 B.n580 10.6151
R1225 B.n581 B.n331 10.6151
R1226 B.n591 B.n331 10.6151
R1227 B.n592 B.n591 10.6151
R1228 B.n593 B.n592 10.6151
R1229 B.n593 B.n323 10.6151
R1230 B.n603 B.n323 10.6151
R1231 B.n604 B.n603 10.6151
R1232 B.n605 B.n604 10.6151
R1233 B.n605 B.n315 10.6151
R1234 B.n615 B.n315 10.6151
R1235 B.n616 B.n615 10.6151
R1236 B.n617 B.n616 10.6151
R1237 B.n617 B.n307 10.6151
R1238 B.n627 B.n307 10.6151
R1239 B.n628 B.n627 10.6151
R1240 B.n629 B.n628 10.6151
R1241 B.n629 B.n299 10.6151
R1242 B.n639 B.n299 10.6151
R1243 B.n640 B.n639 10.6151
R1244 B.n641 B.n640 10.6151
R1245 B.n641 B.n292 10.6151
R1246 B.n651 B.n292 10.6151
R1247 B.n652 B.n651 10.6151
R1248 B.n653 B.n652 10.6151
R1249 B.n653 B.n284 10.6151
R1250 B.n663 B.n284 10.6151
R1251 B.n664 B.n663 10.6151
R1252 B.n665 B.n664 10.6151
R1253 B.n665 B.n277 10.6151
R1254 B.n676 B.n277 10.6151
R1255 B.n677 B.n676 10.6151
R1256 B.n679 B.n677 10.6151
R1257 B.n679 B.n678 10.6151
R1258 B.n678 B.n269 10.6151
R1259 B.n690 B.n269 10.6151
R1260 B.n691 B.n690 10.6151
R1261 B.n692 B.n691 10.6151
R1262 B.n693 B.n692 10.6151
R1263 B.n695 B.n693 10.6151
R1264 B.n696 B.n695 10.6151
R1265 B.n697 B.n696 10.6151
R1266 B.n698 B.n697 10.6151
R1267 B.n700 B.n698 10.6151
R1268 B.n701 B.n700 10.6151
R1269 B.n702 B.n701 10.6151
R1270 B.n703 B.n702 10.6151
R1271 B.n705 B.n703 10.6151
R1272 B.n706 B.n705 10.6151
R1273 B.n707 B.n706 10.6151
R1274 B.n708 B.n707 10.6151
R1275 B.n710 B.n708 10.6151
R1276 B.n711 B.n710 10.6151
R1277 B.n712 B.n711 10.6151
R1278 B.n713 B.n712 10.6151
R1279 B.n715 B.n713 10.6151
R1280 B.n716 B.n715 10.6151
R1281 B.n717 B.n716 10.6151
R1282 B.n718 B.n717 10.6151
R1283 B.n720 B.n718 10.6151
R1284 B.n721 B.n720 10.6151
R1285 B.n722 B.n721 10.6151
R1286 B.n723 B.n722 10.6151
R1287 B.n725 B.n723 10.6151
R1288 B.n726 B.n725 10.6151
R1289 B.n727 B.n726 10.6151
R1290 B.n728 B.n727 10.6151
R1291 B.n730 B.n728 10.6151
R1292 B.n731 B.n730 10.6151
R1293 B.n732 B.n731 10.6151
R1294 B.n733 B.n732 10.6151
R1295 B.n735 B.n733 10.6151
R1296 B.n736 B.n735 10.6151
R1297 B.n737 B.n736 10.6151
R1298 B.n738 B.n737 10.6151
R1299 B.n740 B.n738 10.6151
R1300 B.n741 B.n740 10.6151
R1301 B.n742 B.n741 10.6151
R1302 B.n743 B.n742 10.6151
R1303 B.n745 B.n743 10.6151
R1304 B.n746 B.n745 10.6151
R1305 B.n747 B.n746 10.6151
R1306 B.n748 B.n747 10.6151
R1307 B.n750 B.n748 10.6151
R1308 B.n751 B.n750 10.6151
R1309 B.n752 B.n751 10.6151
R1310 B.n538 B.n537 10.6151
R1311 B.n537 B.n536 10.6151
R1312 B.n536 B.n535 10.6151
R1313 B.n535 B.n533 10.6151
R1314 B.n533 B.n530 10.6151
R1315 B.n530 B.n529 10.6151
R1316 B.n529 B.n526 10.6151
R1317 B.n526 B.n525 10.6151
R1318 B.n525 B.n522 10.6151
R1319 B.n522 B.n521 10.6151
R1320 B.n521 B.n518 10.6151
R1321 B.n518 B.n517 10.6151
R1322 B.n517 B.n514 10.6151
R1323 B.n514 B.n513 10.6151
R1324 B.n513 B.n510 10.6151
R1325 B.n510 B.n509 10.6151
R1326 B.n509 B.n506 10.6151
R1327 B.n506 B.n505 10.6151
R1328 B.n505 B.n502 10.6151
R1329 B.n502 B.n501 10.6151
R1330 B.n501 B.n498 10.6151
R1331 B.n498 B.n497 10.6151
R1332 B.n497 B.n494 10.6151
R1333 B.n494 B.n493 10.6151
R1334 B.n493 B.n490 10.6151
R1335 B.n490 B.n489 10.6151
R1336 B.n489 B.n486 10.6151
R1337 B.n486 B.n485 10.6151
R1338 B.n485 B.n482 10.6151
R1339 B.n480 B.n477 10.6151
R1340 B.n477 B.n476 10.6151
R1341 B.n476 B.n473 10.6151
R1342 B.n473 B.n472 10.6151
R1343 B.n472 B.n469 10.6151
R1344 B.n469 B.n468 10.6151
R1345 B.n468 B.n465 10.6151
R1346 B.n465 B.n464 10.6151
R1347 B.n464 B.n461 10.6151
R1348 B.n459 B.n456 10.6151
R1349 B.n456 B.n455 10.6151
R1350 B.n455 B.n452 10.6151
R1351 B.n452 B.n451 10.6151
R1352 B.n451 B.n448 10.6151
R1353 B.n448 B.n447 10.6151
R1354 B.n447 B.n444 10.6151
R1355 B.n444 B.n443 10.6151
R1356 B.n443 B.n440 10.6151
R1357 B.n440 B.n439 10.6151
R1358 B.n439 B.n436 10.6151
R1359 B.n436 B.n435 10.6151
R1360 B.n435 B.n432 10.6151
R1361 B.n432 B.n431 10.6151
R1362 B.n431 B.n428 10.6151
R1363 B.n428 B.n427 10.6151
R1364 B.n427 B.n424 10.6151
R1365 B.n424 B.n423 10.6151
R1366 B.n423 B.n420 10.6151
R1367 B.n420 B.n419 10.6151
R1368 B.n419 B.n416 10.6151
R1369 B.n416 B.n415 10.6151
R1370 B.n415 B.n412 10.6151
R1371 B.n412 B.n411 10.6151
R1372 B.n411 B.n408 10.6151
R1373 B.n408 B.n407 10.6151
R1374 B.n407 B.n404 10.6151
R1375 B.n404 B.n363 10.6151
R1376 B.n543 B.n363 10.6151
R1377 B.n549 B.n359 10.6151
R1378 B.n550 B.n549 10.6151
R1379 B.n551 B.n550 10.6151
R1380 B.n551 B.n351 10.6151
R1381 B.n561 B.n351 10.6151
R1382 B.n562 B.n561 10.6151
R1383 B.n563 B.n562 10.6151
R1384 B.n563 B.n343 10.6151
R1385 B.n573 B.n343 10.6151
R1386 B.n574 B.n573 10.6151
R1387 B.n575 B.n574 10.6151
R1388 B.n575 B.n335 10.6151
R1389 B.n585 B.n335 10.6151
R1390 B.n586 B.n585 10.6151
R1391 B.n587 B.n586 10.6151
R1392 B.n587 B.n327 10.6151
R1393 B.n597 B.n327 10.6151
R1394 B.n598 B.n597 10.6151
R1395 B.n599 B.n598 10.6151
R1396 B.n599 B.n319 10.6151
R1397 B.n609 B.n319 10.6151
R1398 B.n610 B.n609 10.6151
R1399 B.n611 B.n610 10.6151
R1400 B.n611 B.n311 10.6151
R1401 B.n621 B.n311 10.6151
R1402 B.n622 B.n621 10.6151
R1403 B.n623 B.n622 10.6151
R1404 B.n623 B.n303 10.6151
R1405 B.n633 B.n303 10.6151
R1406 B.n634 B.n633 10.6151
R1407 B.n635 B.n634 10.6151
R1408 B.n635 B.n296 10.6151
R1409 B.n645 B.n296 10.6151
R1410 B.n646 B.n645 10.6151
R1411 B.n647 B.n646 10.6151
R1412 B.n647 B.n288 10.6151
R1413 B.n657 B.n288 10.6151
R1414 B.n658 B.n657 10.6151
R1415 B.n659 B.n658 10.6151
R1416 B.n659 B.n280 10.6151
R1417 B.n670 B.n280 10.6151
R1418 B.n671 B.n670 10.6151
R1419 B.n672 B.n671 10.6151
R1420 B.n672 B.n273 10.6151
R1421 B.n683 B.n273 10.6151
R1422 B.n684 B.n683 10.6151
R1423 B.n685 B.n684 10.6151
R1424 B.n685 B.n0 10.6151
R1425 B.n849 B.n1 10.6151
R1426 B.n849 B.n848 10.6151
R1427 B.n848 B.n847 10.6151
R1428 B.n847 B.n10 10.6151
R1429 B.n841 B.n10 10.6151
R1430 B.n841 B.n840 10.6151
R1431 B.n840 B.n839 10.6151
R1432 B.n839 B.n16 10.6151
R1433 B.n833 B.n16 10.6151
R1434 B.n833 B.n832 10.6151
R1435 B.n832 B.n831 10.6151
R1436 B.n831 B.n24 10.6151
R1437 B.n825 B.n24 10.6151
R1438 B.n825 B.n824 10.6151
R1439 B.n824 B.n823 10.6151
R1440 B.n823 B.n31 10.6151
R1441 B.n818 B.n31 10.6151
R1442 B.n818 B.n817 10.6151
R1443 B.n817 B.n816 10.6151
R1444 B.n816 B.n38 10.6151
R1445 B.n810 B.n38 10.6151
R1446 B.n810 B.n809 10.6151
R1447 B.n809 B.n808 10.6151
R1448 B.n808 B.n45 10.6151
R1449 B.n802 B.n45 10.6151
R1450 B.n802 B.n801 10.6151
R1451 B.n801 B.n800 10.6151
R1452 B.n800 B.n52 10.6151
R1453 B.n794 B.n52 10.6151
R1454 B.n794 B.n793 10.6151
R1455 B.n793 B.n792 10.6151
R1456 B.n792 B.n59 10.6151
R1457 B.n786 B.n59 10.6151
R1458 B.n786 B.n785 10.6151
R1459 B.n785 B.n784 10.6151
R1460 B.n784 B.n66 10.6151
R1461 B.n778 B.n66 10.6151
R1462 B.n778 B.n777 10.6151
R1463 B.n777 B.n776 10.6151
R1464 B.n776 B.n73 10.6151
R1465 B.n770 B.n73 10.6151
R1466 B.n770 B.n769 10.6151
R1467 B.n769 B.n768 10.6151
R1468 B.n768 B.n80 10.6151
R1469 B.n762 B.n80 10.6151
R1470 B.n762 B.n761 10.6151
R1471 B.n761 B.n760 10.6151
R1472 B.n760 B.n87 10.6151
R1473 B.n190 B.n131 9.36635
R1474 B.n213 B.n128 9.36635
R1475 B.n482 B.n481 9.36635
R1476 B.n460 B.n459 9.36635
R1477 B.n855 B.n0 2.81026
R1478 B.n855 B.n1 2.81026
R1479 B.n193 B.n131 1.24928
R1480 B.n210 B.n128 1.24928
R1481 B.n481 B.n480 1.24928
R1482 B.n461 B.n460 1.24928
R1483 VP.n16 VP.n15 161.3
R1484 VP.n17 VP.n12 161.3
R1485 VP.n19 VP.n18 161.3
R1486 VP.n20 VP.n11 161.3
R1487 VP.n22 VP.n21 161.3
R1488 VP.n23 VP.n10 161.3
R1489 VP.n25 VP.n24 161.3
R1490 VP.n49 VP.n48 161.3
R1491 VP.n47 VP.n1 161.3
R1492 VP.n46 VP.n45 161.3
R1493 VP.n44 VP.n2 161.3
R1494 VP.n43 VP.n42 161.3
R1495 VP.n41 VP.n3 161.3
R1496 VP.n40 VP.n39 161.3
R1497 VP.n38 VP.n37 161.3
R1498 VP.n36 VP.n5 161.3
R1499 VP.n35 VP.n34 161.3
R1500 VP.n33 VP.n6 161.3
R1501 VP.n32 VP.n31 161.3
R1502 VP.n30 VP.n7 161.3
R1503 VP.n29 VP.n28 161.3
R1504 VP.n14 VP.t1 94.8717
R1505 VP.n27 VP.n8 78.3232
R1506 VP.n50 VP.n0 78.3232
R1507 VP.n26 VP.n9 78.3232
R1508 VP.n8 VP.t5 62.3097
R1509 VP.n4 VP.t3 62.3097
R1510 VP.n0 VP.t4 62.3097
R1511 VP.n9 VP.t0 62.3097
R1512 VP.n13 VP.t2 62.3097
R1513 VP.n14 VP.n13 62.0291
R1514 VP.n27 VP.n26 48.0031
R1515 VP.n35 VP.n6 40.979
R1516 VP.n42 VP.n2 40.979
R1517 VP.n18 VP.n11 40.979
R1518 VP.n31 VP.n6 40.0078
R1519 VP.n46 VP.n2 40.0078
R1520 VP.n22 VP.n11 40.0078
R1521 VP.n30 VP.n29 24.4675
R1522 VP.n31 VP.n30 24.4675
R1523 VP.n36 VP.n35 24.4675
R1524 VP.n37 VP.n36 24.4675
R1525 VP.n41 VP.n40 24.4675
R1526 VP.n42 VP.n41 24.4675
R1527 VP.n47 VP.n46 24.4675
R1528 VP.n48 VP.n47 24.4675
R1529 VP.n23 VP.n22 24.4675
R1530 VP.n24 VP.n23 24.4675
R1531 VP.n17 VP.n16 24.4675
R1532 VP.n18 VP.n17 24.4675
R1533 VP.n37 VP.n4 12.234
R1534 VP.n40 VP.n4 12.234
R1535 VP.n16 VP.n13 12.234
R1536 VP.n29 VP.n8 11.7447
R1537 VP.n48 VP.n0 11.7447
R1538 VP.n24 VP.n9 11.7447
R1539 VP.n15 VP.n14 4.3015
R1540 VP.n26 VP.n25 0.354971
R1541 VP.n28 VP.n27 0.354971
R1542 VP.n50 VP.n49 0.354971
R1543 VP VP.n50 0.26696
R1544 VP.n15 VP.n12 0.189894
R1545 VP.n19 VP.n12 0.189894
R1546 VP.n20 VP.n19 0.189894
R1547 VP.n21 VP.n20 0.189894
R1548 VP.n21 VP.n10 0.189894
R1549 VP.n25 VP.n10 0.189894
R1550 VP.n28 VP.n7 0.189894
R1551 VP.n32 VP.n7 0.189894
R1552 VP.n33 VP.n32 0.189894
R1553 VP.n34 VP.n33 0.189894
R1554 VP.n34 VP.n5 0.189894
R1555 VP.n38 VP.n5 0.189894
R1556 VP.n39 VP.n38 0.189894
R1557 VP.n39 VP.n3 0.189894
R1558 VP.n43 VP.n3 0.189894
R1559 VP.n44 VP.n43 0.189894
R1560 VP.n45 VP.n44 0.189894
R1561 VP.n45 VP.n1 0.189894
R1562 VP.n49 VP.n1 0.189894
R1563 VTAIL.n7 VTAIL.t4 49.6343
R1564 VTAIL.n11 VTAIL.t0 49.6342
R1565 VTAIL.n2 VTAIL.t9 49.6342
R1566 VTAIL.n10 VTAIL.t8 49.6342
R1567 VTAIL.n9 VTAIL.n8 47.2109
R1568 VTAIL.n6 VTAIL.n5 47.2109
R1569 VTAIL.n1 VTAIL.n0 47.2106
R1570 VTAIL.n4 VTAIL.n3 47.2106
R1571 VTAIL.n6 VTAIL.n4 25.4272
R1572 VTAIL.n11 VTAIL.n10 22.4186
R1573 VTAIL.n7 VTAIL.n6 3.00912
R1574 VTAIL.n10 VTAIL.n9 3.00912
R1575 VTAIL.n4 VTAIL.n2 3.00912
R1576 VTAIL.n0 VTAIL.t5 2.424
R1577 VTAIL.n0 VTAIL.t3 2.424
R1578 VTAIL.n3 VTAIL.t11 2.424
R1579 VTAIL.n3 VTAIL.t10 2.424
R1580 VTAIL.n8 VTAIL.t6 2.424
R1581 VTAIL.n8 VTAIL.t7 2.424
R1582 VTAIL.n5 VTAIL.t1 2.424
R1583 VTAIL.n5 VTAIL.t2 2.424
R1584 VTAIL VTAIL.n11 2.19878
R1585 VTAIL.n9 VTAIL.n7 1.97464
R1586 VTAIL.n2 VTAIL.n1 1.97464
R1587 VTAIL VTAIL.n1 0.810845
R1588 VDD1 VDD1.t4 68.6277
R1589 VDD1.n1 VDD1.t0 68.5141
R1590 VDD1.n1 VDD1.n0 64.5862
R1591 VDD1.n3 VDD1.n2 63.8895
R1592 VDD1.n3 VDD1.n1 42.6237
R1593 VDD1.n2 VDD1.t3 2.424
R1594 VDD1.n2 VDD1.t5 2.424
R1595 VDD1.n0 VDD1.t2 2.424
R1596 VDD1.n0 VDD1.t1 2.424
R1597 VDD1 VDD1.n3 0.694465
R1598 VN.n34 VN.n33 161.3
R1599 VN.n32 VN.n19 161.3
R1600 VN.n31 VN.n30 161.3
R1601 VN.n29 VN.n20 161.3
R1602 VN.n28 VN.n27 161.3
R1603 VN.n26 VN.n21 161.3
R1604 VN.n25 VN.n24 161.3
R1605 VN.n16 VN.n15 161.3
R1606 VN.n14 VN.n1 161.3
R1607 VN.n13 VN.n12 161.3
R1608 VN.n11 VN.n2 161.3
R1609 VN.n10 VN.n9 161.3
R1610 VN.n8 VN.n3 161.3
R1611 VN.n7 VN.n6 161.3
R1612 VN.n23 VN.t4 94.8719
R1613 VN.n5 VN.t2 94.8719
R1614 VN.n17 VN.n0 78.3232
R1615 VN.n35 VN.n18 78.3232
R1616 VN.n4 VN.t1 62.3097
R1617 VN.n0 VN.t3 62.3097
R1618 VN.n22 VN.t0 62.3097
R1619 VN.n18 VN.t5 62.3097
R1620 VN.n5 VN.n4 62.0291
R1621 VN.n23 VN.n22 62.0291
R1622 VN VN.n35 48.1685
R1623 VN.n9 VN.n2 40.979
R1624 VN.n27 VN.n20 40.979
R1625 VN.n13 VN.n2 40.0078
R1626 VN.n31 VN.n20 40.0078
R1627 VN.n8 VN.n7 24.4675
R1628 VN.n9 VN.n8 24.4675
R1629 VN.n14 VN.n13 24.4675
R1630 VN.n15 VN.n14 24.4675
R1631 VN.n27 VN.n26 24.4675
R1632 VN.n26 VN.n25 24.4675
R1633 VN.n33 VN.n32 24.4675
R1634 VN.n32 VN.n31 24.4675
R1635 VN.n7 VN.n4 12.234
R1636 VN.n25 VN.n22 12.234
R1637 VN.n15 VN.n0 11.7447
R1638 VN.n33 VN.n18 11.7447
R1639 VN.n24 VN.n23 4.30152
R1640 VN.n6 VN.n5 4.30152
R1641 VN.n35 VN.n34 0.354971
R1642 VN.n17 VN.n16 0.354971
R1643 VN VN.n17 0.26696
R1644 VN.n34 VN.n19 0.189894
R1645 VN.n30 VN.n19 0.189894
R1646 VN.n30 VN.n29 0.189894
R1647 VN.n29 VN.n28 0.189894
R1648 VN.n28 VN.n21 0.189894
R1649 VN.n24 VN.n21 0.189894
R1650 VN.n6 VN.n3 0.189894
R1651 VN.n10 VN.n3 0.189894
R1652 VN.n11 VN.n10 0.189894
R1653 VN.n12 VN.n11 0.189894
R1654 VN.n12 VN.n1 0.189894
R1655 VN.n16 VN.n1 0.189894
R1656 VDD2.n1 VDD2.t3 68.5141
R1657 VDD2.n2 VDD2.t0 66.3131
R1658 VDD2.n1 VDD2.n0 64.5862
R1659 VDD2 VDD2.n3 64.5835
R1660 VDD2.n2 VDD2.n1 40.5364
R1661 VDD2.n3 VDD2.t5 2.424
R1662 VDD2.n3 VDD2.t1 2.424
R1663 VDD2.n0 VDD2.t4 2.424
R1664 VDD2.n0 VDD2.t2 2.424
R1665 VDD2 VDD2.n2 2.31516
C0 VTAIL VDD2 6.64513f
C1 VTAIL VDD1 6.58929f
C2 VN VDD2 4.86554f
C3 VN VDD1 0.151302f
C4 VP VTAIL 5.35032f
C5 VN VP 6.76687f
C6 VDD1 VDD2 1.62361f
C7 VP VDD2 0.505337f
C8 VP VDD1 5.21705f
C9 VN VTAIL 5.33612f
C10 VDD2 B 5.728473f
C11 VDD1 B 6.079144f
C12 VTAIL B 6.628536f
C13 VN B 14.26205f
C14 VP B 12.970163f
C15 VDD2.t3 B 1.54894f
C16 VDD2.t4 B 0.139457f
C17 VDD2.t2 B 0.139457f
C18 VDD2.n0 B 1.21388f
C19 VDD2.n1 B 2.50388f
C20 VDD2.t0 B 1.53648f
C21 VDD2.n2 B 2.28126f
C22 VDD2.t5 B 0.139457f
C23 VDD2.t1 B 0.139457f
C24 VDD2.n3 B 1.21385f
C25 VN.t3 B 1.52314f
C26 VN.n0 B 0.628717f
C27 VN.n1 B 0.021947f
C28 VN.n2 B 0.01775f
C29 VN.n3 B 0.021947f
C30 VN.t1 B 1.52314f
C31 VN.n4 B 0.621324f
C32 VN.t2 B 1.76354f
C33 VN.n5 B 0.592275f
C34 VN.n6 B 0.255007f
C35 VN.n7 B 0.030807f
C36 VN.n8 B 0.040904f
C37 VN.n9 B 0.043508f
C38 VN.n10 B 0.021947f
C39 VN.n11 B 0.021947f
C40 VN.n12 B 0.021947f
C41 VN.n13 B 0.043728f
C42 VN.n14 B 0.040904f
C43 VN.n15 B 0.030403f
C44 VN.n16 B 0.035423f
C45 VN.n17 B 0.054164f
C46 VN.t5 B 1.52314f
C47 VN.n18 B 0.628717f
C48 VN.n19 B 0.021947f
C49 VN.n20 B 0.01775f
C50 VN.n21 B 0.021947f
C51 VN.t0 B 1.52314f
C52 VN.n22 B 0.621324f
C53 VN.t4 B 1.76354f
C54 VN.n23 B 0.592275f
C55 VN.n24 B 0.255007f
C56 VN.n25 B 0.030807f
C57 VN.n26 B 0.040904f
C58 VN.n27 B 0.043508f
C59 VN.n28 B 0.021947f
C60 VN.n29 B 0.021947f
C61 VN.n30 B 0.021947f
C62 VN.n31 B 0.043728f
C63 VN.n32 B 0.040904f
C64 VN.n33 B 0.030403f
C65 VN.n34 B 0.035423f
C66 VN.n35 B 1.18516f
C67 VDD1.t4 B 1.5793f
C68 VDD1.t0 B 1.57839f
C69 VDD1.t2 B 0.142109f
C70 VDD1.t1 B 0.142109f
C71 VDD1.n0 B 1.23697f
C72 VDD1.n1 B 2.67055f
C73 VDD1.t3 B 0.142109f
C74 VDD1.t5 B 0.142109f
C75 VDD1.n2 B 1.23212f
C76 VDD1.n3 B 2.33134f
C77 VTAIL.t5 B 0.166043f
C78 VTAIL.t3 B 0.166043f
C79 VTAIL.n0 B 1.36869f
C80 VTAIL.n1 B 0.472472f
C81 VTAIL.t9 B 1.74069f
C82 VTAIL.n2 B 0.735482f
C83 VTAIL.t11 B 0.166043f
C84 VTAIL.t10 B 0.166043f
C85 VTAIL.n3 B 1.36869f
C86 VTAIL.n4 B 1.92272f
C87 VTAIL.t1 B 0.166043f
C88 VTAIL.t2 B 0.166043f
C89 VTAIL.n5 B 1.36869f
C90 VTAIL.n6 B 1.92271f
C91 VTAIL.t4 B 1.7407f
C92 VTAIL.n7 B 0.735469f
C93 VTAIL.t6 B 0.166043f
C94 VTAIL.t7 B 0.166043f
C95 VTAIL.n8 B 1.36869f
C96 VTAIL.n9 B 0.65464f
C97 VTAIL.t8 B 1.74069f
C98 VTAIL.n10 B 1.75423f
C99 VTAIL.t0 B 1.74069f
C100 VTAIL.n11 B 1.68708f
C101 VP.t4 B 1.56182f
C102 VP.n0 B 0.64468f
C103 VP.n1 B 0.022505f
C104 VP.n2 B 0.018201f
C105 VP.n3 B 0.022505f
C106 VP.t3 B 1.56182f
C107 VP.n4 B 0.563457f
C108 VP.n5 B 0.022505f
C109 VP.n6 B 0.018201f
C110 VP.n7 B 0.022505f
C111 VP.t5 B 1.56182f
C112 VP.n8 B 0.64468f
C113 VP.t0 B 1.56182f
C114 VP.n9 B 0.64468f
C115 VP.n10 B 0.022505f
C116 VP.n11 B 0.018201f
C117 VP.n12 B 0.022505f
C118 VP.t2 B 1.56182f
C119 VP.n13 B 0.6371f
C120 VP.t1 B 1.80832f
C121 VP.n14 B 0.607314f
C122 VP.n15 B 0.261482f
C123 VP.n16 B 0.031589f
C124 VP.n17 B 0.041943f
C125 VP.n18 B 0.044613f
C126 VP.n19 B 0.022505f
C127 VP.n20 B 0.022505f
C128 VP.n21 B 0.022505f
C129 VP.n22 B 0.044839f
C130 VP.n23 B 0.041943f
C131 VP.n24 B 0.031175f
C132 VP.n25 B 0.036322f
C133 VP.n26 B 1.2059f
C134 VP.n27 B 1.22275f
C135 VP.n28 B 0.036322f
C136 VP.n29 B 0.031175f
C137 VP.n30 B 0.041943f
C138 VP.n31 B 0.044839f
C139 VP.n32 B 0.022505f
C140 VP.n33 B 0.022505f
C141 VP.n34 B 0.022505f
C142 VP.n35 B 0.044613f
C143 VP.n36 B 0.041943f
C144 VP.n37 B 0.031589f
C145 VP.n38 B 0.022505f
C146 VP.n39 B 0.022505f
C147 VP.n40 B 0.031589f
C148 VP.n41 B 0.041943f
C149 VP.n42 B 0.044613f
C150 VP.n43 B 0.022505f
C151 VP.n44 B 0.022505f
C152 VP.n45 B 0.022505f
C153 VP.n46 B 0.044839f
C154 VP.n47 B 0.041943f
C155 VP.n48 B 0.031175f
C156 VP.n49 B 0.036322f
C157 VP.n50 B 0.055539f
.ends

