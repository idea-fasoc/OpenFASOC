* NGSPICE file created from diff_pair_sample_0932.ext - technology: sky130A

.subckt diff_pair_sample_0932 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t5 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=1.46025 ps=9.18 w=8.85 l=1.55
X1 VTAIL.t10 VN.t0 VDD2.t5 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=1.46025 ps=9.18 w=8.85 l=1.55
X2 VDD2.t4 VN.t1 VTAIL.t11 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=3.4515 ps=18.48 w=8.85 l=1.55
X3 VDD1.t2 VP.t1 VTAIL.t8 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=1.46025 ps=9.18 w=8.85 l=1.55
X4 VDD2.t3 VN.t2 VTAIL.t1 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=1.46025 ps=9.18 w=8.85 l=1.55
X5 B.t11 B.t9 B.t10 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=0 ps=0 w=8.85 l=1.55
X6 B.t8 B.t6 B.t7 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=0 ps=0 w=8.85 l=1.55
X7 B.t5 B.t3 B.t4 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=0 ps=0 w=8.85 l=1.55
X8 VDD1.t4 VP.t2 VTAIL.t7 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=3.4515 ps=18.48 w=8.85 l=1.55
X9 VDD2.t2 VN.t3 VTAIL.t2 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=3.4515 ps=18.48 w=8.85 l=1.55
X10 VDD2.t1 VN.t4 VTAIL.t3 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=1.46025 ps=9.18 w=8.85 l=1.55
X11 VDD1.t1 VP.t3 VTAIL.t6 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=3.4515 ps=18.48 w=8.85 l=1.55
X12 B.t2 B.t0 B.t1 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=0 ps=0 w=8.85 l=1.55
X13 VTAIL.t5 VP.t4 VDD1.t3 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=1.46025 ps=9.18 w=8.85 l=1.55
X14 VTAIL.t0 VN.t5 VDD2.t0 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=1.46025 pd=9.18 as=1.46025 ps=9.18 w=8.85 l=1.55
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n2474_n2738# sky130_fd_pr__pfet_01v8 ad=3.4515 pd=18.48 as=1.46025 ps=9.18 w=8.85 l=1.55
R0 VP.n17 VP.n16 179.406
R1 VP.n32 VP.n31 179.406
R2 VP.n15 VP.n14 179.406
R3 VP.n6 VP.t1 169.388
R4 VP.n9 VP.n8 161.3
R5 VP.n10 VP.n5 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n13 VP.n4 161.3
R8 VP.n30 VP.n0 161.3
R9 VP.n29 VP.n28 161.3
R10 VP.n27 VP.n1 161.3
R11 VP.n26 VP.n25 161.3
R12 VP.n23 VP.n2 161.3
R13 VP.n22 VP.n21 161.3
R14 VP.n20 VP.n3 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n17 VP.t5 137.603
R17 VP.n24 VP.t0 137.603
R18 VP.n31 VP.t3 137.603
R19 VP.n14 VP.t2 137.603
R20 VP.n7 VP.t4 137.603
R21 VP.n22 VP.n3 56.5193
R22 VP.n29 VP.n1 56.5193
R23 VP.n12 VP.n5 56.5193
R24 VP.n7 VP.n6 53.7793
R25 VP.n16 VP.n15 42.0535
R26 VP.n18 VP.n3 24.4675
R27 VP.n23 VP.n22 24.4675
R28 VP.n25 VP.n1 24.4675
R29 VP.n30 VP.n29 24.4675
R30 VP.n13 VP.n12 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n9 VP.n6 18.144
R33 VP.n24 VP.n23 12.234
R34 VP.n25 VP.n24 12.234
R35 VP.n8 VP.n7 12.234
R36 VP.n18 VP.n17 6.36192
R37 VP.n31 VP.n30 6.36192
R38 VP.n14 VP.n13 6.36192
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VDD1 VDD1.t2 83.7703
R54 VDD1.n1 VDD1.t0 83.6565
R55 VDD1.n1 VDD1.n0 79.1733
R56 VDD1.n3 VDD1.n2 78.8235
R57 VDD1.n3 VDD1.n1 38.0052
R58 VDD1.n2 VDD1.t3 3.67338
R59 VDD1.n2 VDD1.t4 3.67338
R60 VDD1.n0 VDD1.t5 3.67338
R61 VDD1.n0 VDD1.t1 3.67338
R62 VDD1 VDD1.n3 0.347483
R63 VTAIL.n7 VTAIL.t2 65.8178
R64 VTAIL.n10 VTAIL.t7 65.8175
R65 VTAIL.n11 VTAIL.t11 65.8175
R66 VTAIL.n2 VTAIL.t6 65.8175
R67 VTAIL.n9 VTAIL.n8 62.1449
R68 VTAIL.n6 VTAIL.n5 62.1449
R69 VTAIL.n1 VTAIL.n0 62.1447
R70 VTAIL.n4 VTAIL.n3 62.1447
R71 VTAIL.n6 VTAIL.n4 23.2376
R72 VTAIL.n11 VTAIL.n10 21.6169
R73 VTAIL.n0 VTAIL.t1 3.67338
R74 VTAIL.n0 VTAIL.t0 3.67338
R75 VTAIL.n3 VTAIL.t4 3.67338
R76 VTAIL.n3 VTAIL.t9 3.67338
R77 VTAIL.n8 VTAIL.t8 3.67338
R78 VTAIL.n8 VTAIL.t5 3.67338
R79 VTAIL.n5 VTAIL.t3 3.67338
R80 VTAIL.n5 VTAIL.t10 3.67338
R81 VTAIL.n7 VTAIL.n6 1.62119
R82 VTAIL.n10 VTAIL.n9 1.62119
R83 VTAIL.n4 VTAIL.n2 1.62119
R84 VTAIL.n9 VTAIL.n7 1.28067
R85 VTAIL.n2 VTAIL.n1 1.28067
R86 VTAIL VTAIL.n11 1.15783
R87 VTAIL VTAIL.n1 0.463862
R88 VN.n11 VN.n10 179.406
R89 VN.n23 VN.n22 179.406
R90 VN.n2 VN.t2 169.388
R91 VN.n14 VN.t3 169.388
R92 VN.n21 VN.n12 161.3
R93 VN.n20 VN.n19 161.3
R94 VN.n18 VN.n13 161.3
R95 VN.n17 VN.n16 161.3
R96 VN.n9 VN.n0 161.3
R97 VN.n8 VN.n7 161.3
R98 VN.n6 VN.n1 161.3
R99 VN.n5 VN.n4 161.3
R100 VN.n3 VN.t5 137.603
R101 VN.n10 VN.t1 137.603
R102 VN.n15 VN.t0 137.603
R103 VN.n22 VN.t4 137.603
R104 VN.n8 VN.n1 56.5193
R105 VN.n20 VN.n13 56.5193
R106 VN.n3 VN.n2 53.7793
R107 VN.n15 VN.n14 53.7793
R108 VN VN.n23 42.4342
R109 VN.n4 VN.n1 24.4675
R110 VN.n9 VN.n8 24.4675
R111 VN.n16 VN.n13 24.4675
R112 VN.n21 VN.n20 24.4675
R113 VN.n17 VN.n14 18.144
R114 VN.n5 VN.n2 18.144
R115 VN.n4 VN.n3 12.234
R116 VN.n16 VN.n15 12.234
R117 VN.n10 VN.n9 6.36192
R118 VN.n22 VN.n21 6.36192
R119 VN.n23 VN.n12 0.189894
R120 VN.n19 VN.n12 0.189894
R121 VN.n19 VN.n18 0.189894
R122 VN.n18 VN.n17 0.189894
R123 VN.n6 VN.n5 0.189894
R124 VN.n7 VN.n6 0.189894
R125 VN.n7 VN.n0 0.189894
R126 VN.n11 VN.n0 0.189894
R127 VN VN.n11 0.0516364
R128 VDD2.n1 VDD2.t3 83.6565
R129 VDD2.n2 VDD2.t1 82.4966
R130 VDD2.n1 VDD2.n0 79.1733
R131 VDD2 VDD2.n3 79.1705
R132 VDD2.n2 VDD2.n1 36.6118
R133 VDD2.n3 VDD2.t5 3.67338
R134 VDD2.n3 VDD2.t2 3.67338
R135 VDD2.n0 VDD2.t0 3.67338
R136 VDD2.n0 VDD2.t4 3.67338
R137 VDD2 VDD2.n2 1.27421
R138 B.n393 B.n58 585
R139 B.n395 B.n394 585
R140 B.n396 B.n57 585
R141 B.n398 B.n397 585
R142 B.n399 B.n56 585
R143 B.n401 B.n400 585
R144 B.n402 B.n55 585
R145 B.n404 B.n403 585
R146 B.n405 B.n54 585
R147 B.n407 B.n406 585
R148 B.n408 B.n53 585
R149 B.n410 B.n409 585
R150 B.n411 B.n52 585
R151 B.n413 B.n412 585
R152 B.n414 B.n51 585
R153 B.n416 B.n415 585
R154 B.n417 B.n50 585
R155 B.n419 B.n418 585
R156 B.n420 B.n49 585
R157 B.n422 B.n421 585
R158 B.n423 B.n48 585
R159 B.n425 B.n424 585
R160 B.n426 B.n47 585
R161 B.n428 B.n427 585
R162 B.n429 B.n46 585
R163 B.n431 B.n430 585
R164 B.n432 B.n45 585
R165 B.n434 B.n433 585
R166 B.n435 B.n44 585
R167 B.n437 B.n436 585
R168 B.n438 B.n43 585
R169 B.n440 B.n439 585
R170 B.n442 B.n441 585
R171 B.n443 B.n39 585
R172 B.n445 B.n444 585
R173 B.n446 B.n38 585
R174 B.n448 B.n447 585
R175 B.n449 B.n37 585
R176 B.n451 B.n450 585
R177 B.n452 B.n36 585
R178 B.n454 B.n453 585
R179 B.n455 B.n33 585
R180 B.n458 B.n457 585
R181 B.n459 B.n32 585
R182 B.n461 B.n460 585
R183 B.n462 B.n31 585
R184 B.n464 B.n463 585
R185 B.n465 B.n30 585
R186 B.n467 B.n466 585
R187 B.n468 B.n29 585
R188 B.n470 B.n469 585
R189 B.n471 B.n28 585
R190 B.n473 B.n472 585
R191 B.n474 B.n27 585
R192 B.n476 B.n475 585
R193 B.n477 B.n26 585
R194 B.n479 B.n478 585
R195 B.n480 B.n25 585
R196 B.n482 B.n481 585
R197 B.n483 B.n24 585
R198 B.n485 B.n484 585
R199 B.n486 B.n23 585
R200 B.n488 B.n487 585
R201 B.n489 B.n22 585
R202 B.n491 B.n490 585
R203 B.n492 B.n21 585
R204 B.n494 B.n493 585
R205 B.n495 B.n20 585
R206 B.n497 B.n496 585
R207 B.n498 B.n19 585
R208 B.n500 B.n499 585
R209 B.n501 B.n18 585
R210 B.n503 B.n502 585
R211 B.n504 B.n17 585
R212 B.n392 B.n391 585
R213 B.n390 B.n59 585
R214 B.n389 B.n388 585
R215 B.n387 B.n60 585
R216 B.n386 B.n385 585
R217 B.n384 B.n61 585
R218 B.n383 B.n382 585
R219 B.n381 B.n62 585
R220 B.n380 B.n379 585
R221 B.n378 B.n63 585
R222 B.n377 B.n376 585
R223 B.n375 B.n64 585
R224 B.n374 B.n373 585
R225 B.n372 B.n65 585
R226 B.n371 B.n370 585
R227 B.n369 B.n66 585
R228 B.n368 B.n367 585
R229 B.n366 B.n67 585
R230 B.n365 B.n364 585
R231 B.n363 B.n68 585
R232 B.n362 B.n361 585
R233 B.n360 B.n69 585
R234 B.n359 B.n358 585
R235 B.n357 B.n70 585
R236 B.n356 B.n355 585
R237 B.n354 B.n71 585
R238 B.n353 B.n352 585
R239 B.n351 B.n72 585
R240 B.n350 B.n349 585
R241 B.n348 B.n73 585
R242 B.n347 B.n346 585
R243 B.n345 B.n74 585
R244 B.n344 B.n343 585
R245 B.n342 B.n75 585
R246 B.n341 B.n340 585
R247 B.n339 B.n76 585
R248 B.n338 B.n337 585
R249 B.n336 B.n77 585
R250 B.n335 B.n334 585
R251 B.n333 B.n78 585
R252 B.n332 B.n331 585
R253 B.n330 B.n79 585
R254 B.n329 B.n328 585
R255 B.n327 B.n80 585
R256 B.n326 B.n325 585
R257 B.n324 B.n81 585
R258 B.n323 B.n322 585
R259 B.n321 B.n82 585
R260 B.n320 B.n319 585
R261 B.n318 B.n83 585
R262 B.n317 B.n316 585
R263 B.n315 B.n84 585
R264 B.n314 B.n313 585
R265 B.n312 B.n85 585
R266 B.n311 B.n310 585
R267 B.n309 B.n86 585
R268 B.n308 B.n307 585
R269 B.n306 B.n87 585
R270 B.n305 B.n304 585
R271 B.n303 B.n88 585
R272 B.n302 B.n301 585
R273 B.n189 B.n130 585
R274 B.n191 B.n190 585
R275 B.n192 B.n129 585
R276 B.n194 B.n193 585
R277 B.n195 B.n128 585
R278 B.n197 B.n196 585
R279 B.n198 B.n127 585
R280 B.n200 B.n199 585
R281 B.n201 B.n126 585
R282 B.n203 B.n202 585
R283 B.n204 B.n125 585
R284 B.n206 B.n205 585
R285 B.n207 B.n124 585
R286 B.n209 B.n208 585
R287 B.n210 B.n123 585
R288 B.n212 B.n211 585
R289 B.n213 B.n122 585
R290 B.n215 B.n214 585
R291 B.n216 B.n121 585
R292 B.n218 B.n217 585
R293 B.n219 B.n120 585
R294 B.n221 B.n220 585
R295 B.n222 B.n119 585
R296 B.n224 B.n223 585
R297 B.n225 B.n118 585
R298 B.n227 B.n226 585
R299 B.n228 B.n117 585
R300 B.n230 B.n229 585
R301 B.n231 B.n116 585
R302 B.n233 B.n232 585
R303 B.n234 B.n115 585
R304 B.n236 B.n235 585
R305 B.n238 B.n237 585
R306 B.n239 B.n111 585
R307 B.n241 B.n240 585
R308 B.n242 B.n110 585
R309 B.n244 B.n243 585
R310 B.n245 B.n109 585
R311 B.n247 B.n246 585
R312 B.n248 B.n108 585
R313 B.n250 B.n249 585
R314 B.n251 B.n105 585
R315 B.n254 B.n253 585
R316 B.n255 B.n104 585
R317 B.n257 B.n256 585
R318 B.n258 B.n103 585
R319 B.n260 B.n259 585
R320 B.n261 B.n102 585
R321 B.n263 B.n262 585
R322 B.n264 B.n101 585
R323 B.n266 B.n265 585
R324 B.n267 B.n100 585
R325 B.n269 B.n268 585
R326 B.n270 B.n99 585
R327 B.n272 B.n271 585
R328 B.n273 B.n98 585
R329 B.n275 B.n274 585
R330 B.n276 B.n97 585
R331 B.n278 B.n277 585
R332 B.n279 B.n96 585
R333 B.n281 B.n280 585
R334 B.n282 B.n95 585
R335 B.n284 B.n283 585
R336 B.n285 B.n94 585
R337 B.n287 B.n286 585
R338 B.n288 B.n93 585
R339 B.n290 B.n289 585
R340 B.n291 B.n92 585
R341 B.n293 B.n292 585
R342 B.n294 B.n91 585
R343 B.n296 B.n295 585
R344 B.n297 B.n90 585
R345 B.n299 B.n298 585
R346 B.n300 B.n89 585
R347 B.n188 B.n187 585
R348 B.n186 B.n131 585
R349 B.n185 B.n184 585
R350 B.n183 B.n132 585
R351 B.n182 B.n181 585
R352 B.n180 B.n133 585
R353 B.n179 B.n178 585
R354 B.n177 B.n134 585
R355 B.n176 B.n175 585
R356 B.n174 B.n135 585
R357 B.n173 B.n172 585
R358 B.n171 B.n136 585
R359 B.n170 B.n169 585
R360 B.n168 B.n137 585
R361 B.n167 B.n166 585
R362 B.n165 B.n138 585
R363 B.n164 B.n163 585
R364 B.n162 B.n139 585
R365 B.n161 B.n160 585
R366 B.n159 B.n140 585
R367 B.n158 B.n157 585
R368 B.n156 B.n141 585
R369 B.n155 B.n154 585
R370 B.n153 B.n142 585
R371 B.n152 B.n151 585
R372 B.n150 B.n143 585
R373 B.n149 B.n148 585
R374 B.n147 B.n144 585
R375 B.n146 B.n145 585
R376 B.n2 B.n0 585
R377 B.n549 B.n1 585
R378 B.n548 B.n547 585
R379 B.n546 B.n3 585
R380 B.n545 B.n544 585
R381 B.n543 B.n4 585
R382 B.n542 B.n541 585
R383 B.n540 B.n5 585
R384 B.n539 B.n538 585
R385 B.n537 B.n6 585
R386 B.n536 B.n535 585
R387 B.n534 B.n7 585
R388 B.n533 B.n532 585
R389 B.n531 B.n8 585
R390 B.n530 B.n529 585
R391 B.n528 B.n9 585
R392 B.n527 B.n526 585
R393 B.n525 B.n10 585
R394 B.n524 B.n523 585
R395 B.n522 B.n11 585
R396 B.n521 B.n520 585
R397 B.n519 B.n12 585
R398 B.n518 B.n517 585
R399 B.n516 B.n13 585
R400 B.n515 B.n514 585
R401 B.n513 B.n14 585
R402 B.n512 B.n511 585
R403 B.n510 B.n15 585
R404 B.n509 B.n508 585
R405 B.n507 B.n16 585
R406 B.n506 B.n505 585
R407 B.n551 B.n550 585
R408 B.n189 B.n188 559.769
R409 B.n506 B.n17 559.769
R410 B.n302 B.n89 559.769
R411 B.n393 B.n392 559.769
R412 B.n106 B.t3 343.224
R413 B.n112 B.t0 343.224
R414 B.n34 B.t6 343.224
R415 B.n40 B.t9 343.224
R416 B.n188 B.n131 163.367
R417 B.n184 B.n131 163.367
R418 B.n184 B.n183 163.367
R419 B.n183 B.n182 163.367
R420 B.n182 B.n133 163.367
R421 B.n178 B.n133 163.367
R422 B.n178 B.n177 163.367
R423 B.n177 B.n176 163.367
R424 B.n176 B.n135 163.367
R425 B.n172 B.n135 163.367
R426 B.n172 B.n171 163.367
R427 B.n171 B.n170 163.367
R428 B.n170 B.n137 163.367
R429 B.n166 B.n137 163.367
R430 B.n166 B.n165 163.367
R431 B.n165 B.n164 163.367
R432 B.n164 B.n139 163.367
R433 B.n160 B.n139 163.367
R434 B.n160 B.n159 163.367
R435 B.n159 B.n158 163.367
R436 B.n158 B.n141 163.367
R437 B.n154 B.n141 163.367
R438 B.n154 B.n153 163.367
R439 B.n153 B.n152 163.367
R440 B.n152 B.n143 163.367
R441 B.n148 B.n143 163.367
R442 B.n148 B.n147 163.367
R443 B.n147 B.n146 163.367
R444 B.n146 B.n2 163.367
R445 B.n550 B.n2 163.367
R446 B.n550 B.n549 163.367
R447 B.n549 B.n548 163.367
R448 B.n548 B.n3 163.367
R449 B.n544 B.n3 163.367
R450 B.n544 B.n543 163.367
R451 B.n543 B.n542 163.367
R452 B.n542 B.n5 163.367
R453 B.n538 B.n5 163.367
R454 B.n538 B.n537 163.367
R455 B.n537 B.n536 163.367
R456 B.n536 B.n7 163.367
R457 B.n532 B.n7 163.367
R458 B.n532 B.n531 163.367
R459 B.n531 B.n530 163.367
R460 B.n530 B.n9 163.367
R461 B.n526 B.n9 163.367
R462 B.n526 B.n525 163.367
R463 B.n525 B.n524 163.367
R464 B.n524 B.n11 163.367
R465 B.n520 B.n11 163.367
R466 B.n520 B.n519 163.367
R467 B.n519 B.n518 163.367
R468 B.n518 B.n13 163.367
R469 B.n514 B.n13 163.367
R470 B.n514 B.n513 163.367
R471 B.n513 B.n512 163.367
R472 B.n512 B.n15 163.367
R473 B.n508 B.n15 163.367
R474 B.n508 B.n507 163.367
R475 B.n507 B.n506 163.367
R476 B.n190 B.n189 163.367
R477 B.n190 B.n129 163.367
R478 B.n194 B.n129 163.367
R479 B.n195 B.n194 163.367
R480 B.n196 B.n195 163.367
R481 B.n196 B.n127 163.367
R482 B.n200 B.n127 163.367
R483 B.n201 B.n200 163.367
R484 B.n202 B.n201 163.367
R485 B.n202 B.n125 163.367
R486 B.n206 B.n125 163.367
R487 B.n207 B.n206 163.367
R488 B.n208 B.n207 163.367
R489 B.n208 B.n123 163.367
R490 B.n212 B.n123 163.367
R491 B.n213 B.n212 163.367
R492 B.n214 B.n213 163.367
R493 B.n214 B.n121 163.367
R494 B.n218 B.n121 163.367
R495 B.n219 B.n218 163.367
R496 B.n220 B.n219 163.367
R497 B.n220 B.n119 163.367
R498 B.n224 B.n119 163.367
R499 B.n225 B.n224 163.367
R500 B.n226 B.n225 163.367
R501 B.n226 B.n117 163.367
R502 B.n230 B.n117 163.367
R503 B.n231 B.n230 163.367
R504 B.n232 B.n231 163.367
R505 B.n232 B.n115 163.367
R506 B.n236 B.n115 163.367
R507 B.n237 B.n236 163.367
R508 B.n237 B.n111 163.367
R509 B.n241 B.n111 163.367
R510 B.n242 B.n241 163.367
R511 B.n243 B.n242 163.367
R512 B.n243 B.n109 163.367
R513 B.n247 B.n109 163.367
R514 B.n248 B.n247 163.367
R515 B.n249 B.n248 163.367
R516 B.n249 B.n105 163.367
R517 B.n254 B.n105 163.367
R518 B.n255 B.n254 163.367
R519 B.n256 B.n255 163.367
R520 B.n256 B.n103 163.367
R521 B.n260 B.n103 163.367
R522 B.n261 B.n260 163.367
R523 B.n262 B.n261 163.367
R524 B.n262 B.n101 163.367
R525 B.n266 B.n101 163.367
R526 B.n267 B.n266 163.367
R527 B.n268 B.n267 163.367
R528 B.n268 B.n99 163.367
R529 B.n272 B.n99 163.367
R530 B.n273 B.n272 163.367
R531 B.n274 B.n273 163.367
R532 B.n274 B.n97 163.367
R533 B.n278 B.n97 163.367
R534 B.n279 B.n278 163.367
R535 B.n280 B.n279 163.367
R536 B.n280 B.n95 163.367
R537 B.n284 B.n95 163.367
R538 B.n285 B.n284 163.367
R539 B.n286 B.n285 163.367
R540 B.n286 B.n93 163.367
R541 B.n290 B.n93 163.367
R542 B.n291 B.n290 163.367
R543 B.n292 B.n291 163.367
R544 B.n292 B.n91 163.367
R545 B.n296 B.n91 163.367
R546 B.n297 B.n296 163.367
R547 B.n298 B.n297 163.367
R548 B.n298 B.n89 163.367
R549 B.n303 B.n302 163.367
R550 B.n304 B.n303 163.367
R551 B.n304 B.n87 163.367
R552 B.n308 B.n87 163.367
R553 B.n309 B.n308 163.367
R554 B.n310 B.n309 163.367
R555 B.n310 B.n85 163.367
R556 B.n314 B.n85 163.367
R557 B.n315 B.n314 163.367
R558 B.n316 B.n315 163.367
R559 B.n316 B.n83 163.367
R560 B.n320 B.n83 163.367
R561 B.n321 B.n320 163.367
R562 B.n322 B.n321 163.367
R563 B.n322 B.n81 163.367
R564 B.n326 B.n81 163.367
R565 B.n327 B.n326 163.367
R566 B.n328 B.n327 163.367
R567 B.n328 B.n79 163.367
R568 B.n332 B.n79 163.367
R569 B.n333 B.n332 163.367
R570 B.n334 B.n333 163.367
R571 B.n334 B.n77 163.367
R572 B.n338 B.n77 163.367
R573 B.n339 B.n338 163.367
R574 B.n340 B.n339 163.367
R575 B.n340 B.n75 163.367
R576 B.n344 B.n75 163.367
R577 B.n345 B.n344 163.367
R578 B.n346 B.n345 163.367
R579 B.n346 B.n73 163.367
R580 B.n350 B.n73 163.367
R581 B.n351 B.n350 163.367
R582 B.n352 B.n351 163.367
R583 B.n352 B.n71 163.367
R584 B.n356 B.n71 163.367
R585 B.n357 B.n356 163.367
R586 B.n358 B.n357 163.367
R587 B.n358 B.n69 163.367
R588 B.n362 B.n69 163.367
R589 B.n363 B.n362 163.367
R590 B.n364 B.n363 163.367
R591 B.n364 B.n67 163.367
R592 B.n368 B.n67 163.367
R593 B.n369 B.n368 163.367
R594 B.n370 B.n369 163.367
R595 B.n370 B.n65 163.367
R596 B.n374 B.n65 163.367
R597 B.n375 B.n374 163.367
R598 B.n376 B.n375 163.367
R599 B.n376 B.n63 163.367
R600 B.n380 B.n63 163.367
R601 B.n381 B.n380 163.367
R602 B.n382 B.n381 163.367
R603 B.n382 B.n61 163.367
R604 B.n386 B.n61 163.367
R605 B.n387 B.n386 163.367
R606 B.n388 B.n387 163.367
R607 B.n388 B.n59 163.367
R608 B.n392 B.n59 163.367
R609 B.n502 B.n17 163.367
R610 B.n502 B.n501 163.367
R611 B.n501 B.n500 163.367
R612 B.n500 B.n19 163.367
R613 B.n496 B.n19 163.367
R614 B.n496 B.n495 163.367
R615 B.n495 B.n494 163.367
R616 B.n494 B.n21 163.367
R617 B.n490 B.n21 163.367
R618 B.n490 B.n489 163.367
R619 B.n489 B.n488 163.367
R620 B.n488 B.n23 163.367
R621 B.n484 B.n23 163.367
R622 B.n484 B.n483 163.367
R623 B.n483 B.n482 163.367
R624 B.n482 B.n25 163.367
R625 B.n478 B.n25 163.367
R626 B.n478 B.n477 163.367
R627 B.n477 B.n476 163.367
R628 B.n476 B.n27 163.367
R629 B.n472 B.n27 163.367
R630 B.n472 B.n471 163.367
R631 B.n471 B.n470 163.367
R632 B.n470 B.n29 163.367
R633 B.n466 B.n29 163.367
R634 B.n466 B.n465 163.367
R635 B.n465 B.n464 163.367
R636 B.n464 B.n31 163.367
R637 B.n460 B.n31 163.367
R638 B.n460 B.n459 163.367
R639 B.n459 B.n458 163.367
R640 B.n458 B.n33 163.367
R641 B.n453 B.n33 163.367
R642 B.n453 B.n452 163.367
R643 B.n452 B.n451 163.367
R644 B.n451 B.n37 163.367
R645 B.n447 B.n37 163.367
R646 B.n447 B.n446 163.367
R647 B.n446 B.n445 163.367
R648 B.n445 B.n39 163.367
R649 B.n441 B.n39 163.367
R650 B.n441 B.n440 163.367
R651 B.n440 B.n43 163.367
R652 B.n436 B.n43 163.367
R653 B.n436 B.n435 163.367
R654 B.n435 B.n434 163.367
R655 B.n434 B.n45 163.367
R656 B.n430 B.n45 163.367
R657 B.n430 B.n429 163.367
R658 B.n429 B.n428 163.367
R659 B.n428 B.n47 163.367
R660 B.n424 B.n47 163.367
R661 B.n424 B.n423 163.367
R662 B.n423 B.n422 163.367
R663 B.n422 B.n49 163.367
R664 B.n418 B.n49 163.367
R665 B.n418 B.n417 163.367
R666 B.n417 B.n416 163.367
R667 B.n416 B.n51 163.367
R668 B.n412 B.n51 163.367
R669 B.n412 B.n411 163.367
R670 B.n411 B.n410 163.367
R671 B.n410 B.n53 163.367
R672 B.n406 B.n53 163.367
R673 B.n406 B.n405 163.367
R674 B.n405 B.n404 163.367
R675 B.n404 B.n55 163.367
R676 B.n400 B.n55 163.367
R677 B.n400 B.n399 163.367
R678 B.n399 B.n398 163.367
R679 B.n398 B.n57 163.367
R680 B.n394 B.n57 163.367
R681 B.n394 B.n393 163.367
R682 B.n106 B.t5 144.81
R683 B.n40 B.t10 144.81
R684 B.n112 B.t2 144.799
R685 B.n34 B.t7 144.799
R686 B.n107 B.t4 108.35
R687 B.n41 B.t11 108.35
R688 B.n113 B.t1 108.34
R689 B.n35 B.t8 108.34
R690 B.n252 B.n107 59.5399
R691 B.n114 B.n113 59.5399
R692 B.n456 B.n35 59.5399
R693 B.n42 B.n41 59.5399
R694 B.n107 B.n106 36.4611
R695 B.n113 B.n112 36.4611
R696 B.n35 B.n34 36.4611
R697 B.n41 B.n40 36.4611
R698 B.n505 B.n504 36.3712
R699 B.n391 B.n58 36.3712
R700 B.n301 B.n300 36.3712
R701 B.n187 B.n130 36.3712
R702 B B.n551 18.0485
R703 B.n504 B.n503 10.6151
R704 B.n503 B.n18 10.6151
R705 B.n499 B.n18 10.6151
R706 B.n499 B.n498 10.6151
R707 B.n498 B.n497 10.6151
R708 B.n497 B.n20 10.6151
R709 B.n493 B.n20 10.6151
R710 B.n493 B.n492 10.6151
R711 B.n492 B.n491 10.6151
R712 B.n491 B.n22 10.6151
R713 B.n487 B.n22 10.6151
R714 B.n487 B.n486 10.6151
R715 B.n486 B.n485 10.6151
R716 B.n485 B.n24 10.6151
R717 B.n481 B.n24 10.6151
R718 B.n481 B.n480 10.6151
R719 B.n480 B.n479 10.6151
R720 B.n479 B.n26 10.6151
R721 B.n475 B.n26 10.6151
R722 B.n475 B.n474 10.6151
R723 B.n474 B.n473 10.6151
R724 B.n473 B.n28 10.6151
R725 B.n469 B.n28 10.6151
R726 B.n469 B.n468 10.6151
R727 B.n468 B.n467 10.6151
R728 B.n467 B.n30 10.6151
R729 B.n463 B.n30 10.6151
R730 B.n463 B.n462 10.6151
R731 B.n462 B.n461 10.6151
R732 B.n461 B.n32 10.6151
R733 B.n457 B.n32 10.6151
R734 B.n455 B.n454 10.6151
R735 B.n454 B.n36 10.6151
R736 B.n450 B.n36 10.6151
R737 B.n450 B.n449 10.6151
R738 B.n449 B.n448 10.6151
R739 B.n448 B.n38 10.6151
R740 B.n444 B.n38 10.6151
R741 B.n444 B.n443 10.6151
R742 B.n443 B.n442 10.6151
R743 B.n439 B.n438 10.6151
R744 B.n438 B.n437 10.6151
R745 B.n437 B.n44 10.6151
R746 B.n433 B.n44 10.6151
R747 B.n433 B.n432 10.6151
R748 B.n432 B.n431 10.6151
R749 B.n431 B.n46 10.6151
R750 B.n427 B.n46 10.6151
R751 B.n427 B.n426 10.6151
R752 B.n426 B.n425 10.6151
R753 B.n425 B.n48 10.6151
R754 B.n421 B.n48 10.6151
R755 B.n421 B.n420 10.6151
R756 B.n420 B.n419 10.6151
R757 B.n419 B.n50 10.6151
R758 B.n415 B.n50 10.6151
R759 B.n415 B.n414 10.6151
R760 B.n414 B.n413 10.6151
R761 B.n413 B.n52 10.6151
R762 B.n409 B.n52 10.6151
R763 B.n409 B.n408 10.6151
R764 B.n408 B.n407 10.6151
R765 B.n407 B.n54 10.6151
R766 B.n403 B.n54 10.6151
R767 B.n403 B.n402 10.6151
R768 B.n402 B.n401 10.6151
R769 B.n401 B.n56 10.6151
R770 B.n397 B.n56 10.6151
R771 B.n397 B.n396 10.6151
R772 B.n396 B.n395 10.6151
R773 B.n395 B.n58 10.6151
R774 B.n301 B.n88 10.6151
R775 B.n305 B.n88 10.6151
R776 B.n306 B.n305 10.6151
R777 B.n307 B.n306 10.6151
R778 B.n307 B.n86 10.6151
R779 B.n311 B.n86 10.6151
R780 B.n312 B.n311 10.6151
R781 B.n313 B.n312 10.6151
R782 B.n313 B.n84 10.6151
R783 B.n317 B.n84 10.6151
R784 B.n318 B.n317 10.6151
R785 B.n319 B.n318 10.6151
R786 B.n319 B.n82 10.6151
R787 B.n323 B.n82 10.6151
R788 B.n324 B.n323 10.6151
R789 B.n325 B.n324 10.6151
R790 B.n325 B.n80 10.6151
R791 B.n329 B.n80 10.6151
R792 B.n330 B.n329 10.6151
R793 B.n331 B.n330 10.6151
R794 B.n331 B.n78 10.6151
R795 B.n335 B.n78 10.6151
R796 B.n336 B.n335 10.6151
R797 B.n337 B.n336 10.6151
R798 B.n337 B.n76 10.6151
R799 B.n341 B.n76 10.6151
R800 B.n342 B.n341 10.6151
R801 B.n343 B.n342 10.6151
R802 B.n343 B.n74 10.6151
R803 B.n347 B.n74 10.6151
R804 B.n348 B.n347 10.6151
R805 B.n349 B.n348 10.6151
R806 B.n349 B.n72 10.6151
R807 B.n353 B.n72 10.6151
R808 B.n354 B.n353 10.6151
R809 B.n355 B.n354 10.6151
R810 B.n355 B.n70 10.6151
R811 B.n359 B.n70 10.6151
R812 B.n360 B.n359 10.6151
R813 B.n361 B.n360 10.6151
R814 B.n361 B.n68 10.6151
R815 B.n365 B.n68 10.6151
R816 B.n366 B.n365 10.6151
R817 B.n367 B.n366 10.6151
R818 B.n367 B.n66 10.6151
R819 B.n371 B.n66 10.6151
R820 B.n372 B.n371 10.6151
R821 B.n373 B.n372 10.6151
R822 B.n373 B.n64 10.6151
R823 B.n377 B.n64 10.6151
R824 B.n378 B.n377 10.6151
R825 B.n379 B.n378 10.6151
R826 B.n379 B.n62 10.6151
R827 B.n383 B.n62 10.6151
R828 B.n384 B.n383 10.6151
R829 B.n385 B.n384 10.6151
R830 B.n385 B.n60 10.6151
R831 B.n389 B.n60 10.6151
R832 B.n390 B.n389 10.6151
R833 B.n391 B.n390 10.6151
R834 B.n191 B.n130 10.6151
R835 B.n192 B.n191 10.6151
R836 B.n193 B.n192 10.6151
R837 B.n193 B.n128 10.6151
R838 B.n197 B.n128 10.6151
R839 B.n198 B.n197 10.6151
R840 B.n199 B.n198 10.6151
R841 B.n199 B.n126 10.6151
R842 B.n203 B.n126 10.6151
R843 B.n204 B.n203 10.6151
R844 B.n205 B.n204 10.6151
R845 B.n205 B.n124 10.6151
R846 B.n209 B.n124 10.6151
R847 B.n210 B.n209 10.6151
R848 B.n211 B.n210 10.6151
R849 B.n211 B.n122 10.6151
R850 B.n215 B.n122 10.6151
R851 B.n216 B.n215 10.6151
R852 B.n217 B.n216 10.6151
R853 B.n217 B.n120 10.6151
R854 B.n221 B.n120 10.6151
R855 B.n222 B.n221 10.6151
R856 B.n223 B.n222 10.6151
R857 B.n223 B.n118 10.6151
R858 B.n227 B.n118 10.6151
R859 B.n228 B.n227 10.6151
R860 B.n229 B.n228 10.6151
R861 B.n229 B.n116 10.6151
R862 B.n233 B.n116 10.6151
R863 B.n234 B.n233 10.6151
R864 B.n235 B.n234 10.6151
R865 B.n239 B.n238 10.6151
R866 B.n240 B.n239 10.6151
R867 B.n240 B.n110 10.6151
R868 B.n244 B.n110 10.6151
R869 B.n245 B.n244 10.6151
R870 B.n246 B.n245 10.6151
R871 B.n246 B.n108 10.6151
R872 B.n250 B.n108 10.6151
R873 B.n251 B.n250 10.6151
R874 B.n253 B.n104 10.6151
R875 B.n257 B.n104 10.6151
R876 B.n258 B.n257 10.6151
R877 B.n259 B.n258 10.6151
R878 B.n259 B.n102 10.6151
R879 B.n263 B.n102 10.6151
R880 B.n264 B.n263 10.6151
R881 B.n265 B.n264 10.6151
R882 B.n265 B.n100 10.6151
R883 B.n269 B.n100 10.6151
R884 B.n270 B.n269 10.6151
R885 B.n271 B.n270 10.6151
R886 B.n271 B.n98 10.6151
R887 B.n275 B.n98 10.6151
R888 B.n276 B.n275 10.6151
R889 B.n277 B.n276 10.6151
R890 B.n277 B.n96 10.6151
R891 B.n281 B.n96 10.6151
R892 B.n282 B.n281 10.6151
R893 B.n283 B.n282 10.6151
R894 B.n283 B.n94 10.6151
R895 B.n287 B.n94 10.6151
R896 B.n288 B.n287 10.6151
R897 B.n289 B.n288 10.6151
R898 B.n289 B.n92 10.6151
R899 B.n293 B.n92 10.6151
R900 B.n294 B.n293 10.6151
R901 B.n295 B.n294 10.6151
R902 B.n295 B.n90 10.6151
R903 B.n299 B.n90 10.6151
R904 B.n300 B.n299 10.6151
R905 B.n187 B.n186 10.6151
R906 B.n186 B.n185 10.6151
R907 B.n185 B.n132 10.6151
R908 B.n181 B.n132 10.6151
R909 B.n181 B.n180 10.6151
R910 B.n180 B.n179 10.6151
R911 B.n179 B.n134 10.6151
R912 B.n175 B.n134 10.6151
R913 B.n175 B.n174 10.6151
R914 B.n174 B.n173 10.6151
R915 B.n173 B.n136 10.6151
R916 B.n169 B.n136 10.6151
R917 B.n169 B.n168 10.6151
R918 B.n168 B.n167 10.6151
R919 B.n167 B.n138 10.6151
R920 B.n163 B.n138 10.6151
R921 B.n163 B.n162 10.6151
R922 B.n162 B.n161 10.6151
R923 B.n161 B.n140 10.6151
R924 B.n157 B.n140 10.6151
R925 B.n157 B.n156 10.6151
R926 B.n156 B.n155 10.6151
R927 B.n155 B.n142 10.6151
R928 B.n151 B.n142 10.6151
R929 B.n151 B.n150 10.6151
R930 B.n150 B.n149 10.6151
R931 B.n149 B.n144 10.6151
R932 B.n145 B.n144 10.6151
R933 B.n145 B.n0 10.6151
R934 B.n547 B.n1 10.6151
R935 B.n547 B.n546 10.6151
R936 B.n546 B.n545 10.6151
R937 B.n545 B.n4 10.6151
R938 B.n541 B.n4 10.6151
R939 B.n541 B.n540 10.6151
R940 B.n540 B.n539 10.6151
R941 B.n539 B.n6 10.6151
R942 B.n535 B.n6 10.6151
R943 B.n535 B.n534 10.6151
R944 B.n534 B.n533 10.6151
R945 B.n533 B.n8 10.6151
R946 B.n529 B.n8 10.6151
R947 B.n529 B.n528 10.6151
R948 B.n528 B.n527 10.6151
R949 B.n527 B.n10 10.6151
R950 B.n523 B.n10 10.6151
R951 B.n523 B.n522 10.6151
R952 B.n522 B.n521 10.6151
R953 B.n521 B.n12 10.6151
R954 B.n517 B.n12 10.6151
R955 B.n517 B.n516 10.6151
R956 B.n516 B.n515 10.6151
R957 B.n515 B.n14 10.6151
R958 B.n511 B.n14 10.6151
R959 B.n511 B.n510 10.6151
R960 B.n510 B.n509 10.6151
R961 B.n509 B.n16 10.6151
R962 B.n505 B.n16 10.6151
R963 B.n457 B.n456 9.36635
R964 B.n439 B.n42 9.36635
R965 B.n235 B.n114 9.36635
R966 B.n253 B.n252 9.36635
R967 B.n551 B.n0 2.81026
R968 B.n551 B.n1 2.81026
R969 B.n456 B.n455 1.24928
R970 B.n442 B.n42 1.24928
R971 B.n238 B.n114 1.24928
R972 B.n252 B.n251 1.24928
C0 VTAIL VN 4.51185f
C1 VDD1 B 1.56826f
C2 VDD1 VN 0.149371f
C3 B VP 1.4319f
C4 VP VN 5.32442f
C5 B VN 0.908043f
C6 VDD2 w_n2474_n2738# 1.86107f
C7 VTAIL w_n2474_n2738# 2.45156f
C8 VDD1 w_n2474_n2738# 1.80975f
C9 VTAIL VDD2 6.57288f
C10 VDD1 VDD2 1.0259f
C11 VDD1 VTAIL 6.52953f
C12 VP w_n2474_n2738# 4.69191f
C13 VDD2 VP 0.369129f
C14 B w_n2474_n2738# 7.34308f
C15 w_n2474_n2738# VN 4.37498f
C16 VTAIL VP 4.52618f
C17 B VDD2 1.61727f
C18 VDD2 VN 4.46923f
C19 VDD1 VP 4.68611f
C20 VTAIL B 2.57024f
C21 VDD2 VSUBS 1.322367f
C22 VDD1 VSUBS 1.696694f
C23 VTAIL VSUBS 0.869445f
C24 VN VSUBS 4.74694f
C25 VP VSUBS 1.993649f
C26 B VSUBS 3.332836f
C27 w_n2474_n2738# VSUBS 83.8686f
C28 B.n0 VSUBS 0.004579f
C29 B.n1 VSUBS 0.004579f
C30 B.n2 VSUBS 0.007242f
C31 B.n3 VSUBS 0.007242f
C32 B.n4 VSUBS 0.007242f
C33 B.n5 VSUBS 0.007242f
C34 B.n6 VSUBS 0.007242f
C35 B.n7 VSUBS 0.007242f
C36 B.n8 VSUBS 0.007242f
C37 B.n9 VSUBS 0.007242f
C38 B.n10 VSUBS 0.007242f
C39 B.n11 VSUBS 0.007242f
C40 B.n12 VSUBS 0.007242f
C41 B.n13 VSUBS 0.007242f
C42 B.n14 VSUBS 0.007242f
C43 B.n15 VSUBS 0.007242f
C44 B.n16 VSUBS 0.007242f
C45 B.n17 VSUBS 0.018632f
C46 B.n18 VSUBS 0.007242f
C47 B.n19 VSUBS 0.007242f
C48 B.n20 VSUBS 0.007242f
C49 B.n21 VSUBS 0.007242f
C50 B.n22 VSUBS 0.007242f
C51 B.n23 VSUBS 0.007242f
C52 B.n24 VSUBS 0.007242f
C53 B.n25 VSUBS 0.007242f
C54 B.n26 VSUBS 0.007242f
C55 B.n27 VSUBS 0.007242f
C56 B.n28 VSUBS 0.007242f
C57 B.n29 VSUBS 0.007242f
C58 B.n30 VSUBS 0.007242f
C59 B.n31 VSUBS 0.007242f
C60 B.n32 VSUBS 0.007242f
C61 B.n33 VSUBS 0.007242f
C62 B.t8 VSUBS 0.287062f
C63 B.t7 VSUBS 0.30195f
C64 B.t6 VSUBS 0.635428f
C65 B.n34 VSUBS 0.143194f
C66 B.n35 VSUBS 0.069458f
C67 B.n36 VSUBS 0.007242f
C68 B.n37 VSUBS 0.007242f
C69 B.n38 VSUBS 0.007242f
C70 B.n39 VSUBS 0.007242f
C71 B.t11 VSUBS 0.287059f
C72 B.t10 VSUBS 0.301947f
C73 B.t9 VSUBS 0.635428f
C74 B.n40 VSUBS 0.143197f
C75 B.n41 VSUBS 0.069461f
C76 B.n42 VSUBS 0.016778f
C77 B.n43 VSUBS 0.007242f
C78 B.n44 VSUBS 0.007242f
C79 B.n45 VSUBS 0.007242f
C80 B.n46 VSUBS 0.007242f
C81 B.n47 VSUBS 0.007242f
C82 B.n48 VSUBS 0.007242f
C83 B.n49 VSUBS 0.007242f
C84 B.n50 VSUBS 0.007242f
C85 B.n51 VSUBS 0.007242f
C86 B.n52 VSUBS 0.007242f
C87 B.n53 VSUBS 0.007242f
C88 B.n54 VSUBS 0.007242f
C89 B.n55 VSUBS 0.007242f
C90 B.n56 VSUBS 0.007242f
C91 B.n57 VSUBS 0.007242f
C92 B.n58 VSUBS 0.017864f
C93 B.n59 VSUBS 0.007242f
C94 B.n60 VSUBS 0.007242f
C95 B.n61 VSUBS 0.007242f
C96 B.n62 VSUBS 0.007242f
C97 B.n63 VSUBS 0.007242f
C98 B.n64 VSUBS 0.007242f
C99 B.n65 VSUBS 0.007242f
C100 B.n66 VSUBS 0.007242f
C101 B.n67 VSUBS 0.007242f
C102 B.n68 VSUBS 0.007242f
C103 B.n69 VSUBS 0.007242f
C104 B.n70 VSUBS 0.007242f
C105 B.n71 VSUBS 0.007242f
C106 B.n72 VSUBS 0.007242f
C107 B.n73 VSUBS 0.007242f
C108 B.n74 VSUBS 0.007242f
C109 B.n75 VSUBS 0.007242f
C110 B.n76 VSUBS 0.007242f
C111 B.n77 VSUBS 0.007242f
C112 B.n78 VSUBS 0.007242f
C113 B.n79 VSUBS 0.007242f
C114 B.n80 VSUBS 0.007242f
C115 B.n81 VSUBS 0.007242f
C116 B.n82 VSUBS 0.007242f
C117 B.n83 VSUBS 0.007242f
C118 B.n84 VSUBS 0.007242f
C119 B.n85 VSUBS 0.007242f
C120 B.n86 VSUBS 0.007242f
C121 B.n87 VSUBS 0.007242f
C122 B.n88 VSUBS 0.007242f
C123 B.n89 VSUBS 0.018632f
C124 B.n90 VSUBS 0.007242f
C125 B.n91 VSUBS 0.007242f
C126 B.n92 VSUBS 0.007242f
C127 B.n93 VSUBS 0.007242f
C128 B.n94 VSUBS 0.007242f
C129 B.n95 VSUBS 0.007242f
C130 B.n96 VSUBS 0.007242f
C131 B.n97 VSUBS 0.007242f
C132 B.n98 VSUBS 0.007242f
C133 B.n99 VSUBS 0.007242f
C134 B.n100 VSUBS 0.007242f
C135 B.n101 VSUBS 0.007242f
C136 B.n102 VSUBS 0.007242f
C137 B.n103 VSUBS 0.007242f
C138 B.n104 VSUBS 0.007242f
C139 B.n105 VSUBS 0.007242f
C140 B.t4 VSUBS 0.287059f
C141 B.t5 VSUBS 0.301947f
C142 B.t3 VSUBS 0.635428f
C143 B.n106 VSUBS 0.143197f
C144 B.n107 VSUBS 0.069461f
C145 B.n108 VSUBS 0.007242f
C146 B.n109 VSUBS 0.007242f
C147 B.n110 VSUBS 0.007242f
C148 B.n111 VSUBS 0.007242f
C149 B.t1 VSUBS 0.287062f
C150 B.t2 VSUBS 0.30195f
C151 B.t0 VSUBS 0.635428f
C152 B.n112 VSUBS 0.143194f
C153 B.n113 VSUBS 0.069458f
C154 B.n114 VSUBS 0.016778f
C155 B.n115 VSUBS 0.007242f
C156 B.n116 VSUBS 0.007242f
C157 B.n117 VSUBS 0.007242f
C158 B.n118 VSUBS 0.007242f
C159 B.n119 VSUBS 0.007242f
C160 B.n120 VSUBS 0.007242f
C161 B.n121 VSUBS 0.007242f
C162 B.n122 VSUBS 0.007242f
C163 B.n123 VSUBS 0.007242f
C164 B.n124 VSUBS 0.007242f
C165 B.n125 VSUBS 0.007242f
C166 B.n126 VSUBS 0.007242f
C167 B.n127 VSUBS 0.007242f
C168 B.n128 VSUBS 0.007242f
C169 B.n129 VSUBS 0.007242f
C170 B.n130 VSUBS 0.018632f
C171 B.n131 VSUBS 0.007242f
C172 B.n132 VSUBS 0.007242f
C173 B.n133 VSUBS 0.007242f
C174 B.n134 VSUBS 0.007242f
C175 B.n135 VSUBS 0.007242f
C176 B.n136 VSUBS 0.007242f
C177 B.n137 VSUBS 0.007242f
C178 B.n138 VSUBS 0.007242f
C179 B.n139 VSUBS 0.007242f
C180 B.n140 VSUBS 0.007242f
C181 B.n141 VSUBS 0.007242f
C182 B.n142 VSUBS 0.007242f
C183 B.n143 VSUBS 0.007242f
C184 B.n144 VSUBS 0.007242f
C185 B.n145 VSUBS 0.007242f
C186 B.n146 VSUBS 0.007242f
C187 B.n147 VSUBS 0.007242f
C188 B.n148 VSUBS 0.007242f
C189 B.n149 VSUBS 0.007242f
C190 B.n150 VSUBS 0.007242f
C191 B.n151 VSUBS 0.007242f
C192 B.n152 VSUBS 0.007242f
C193 B.n153 VSUBS 0.007242f
C194 B.n154 VSUBS 0.007242f
C195 B.n155 VSUBS 0.007242f
C196 B.n156 VSUBS 0.007242f
C197 B.n157 VSUBS 0.007242f
C198 B.n158 VSUBS 0.007242f
C199 B.n159 VSUBS 0.007242f
C200 B.n160 VSUBS 0.007242f
C201 B.n161 VSUBS 0.007242f
C202 B.n162 VSUBS 0.007242f
C203 B.n163 VSUBS 0.007242f
C204 B.n164 VSUBS 0.007242f
C205 B.n165 VSUBS 0.007242f
C206 B.n166 VSUBS 0.007242f
C207 B.n167 VSUBS 0.007242f
C208 B.n168 VSUBS 0.007242f
C209 B.n169 VSUBS 0.007242f
C210 B.n170 VSUBS 0.007242f
C211 B.n171 VSUBS 0.007242f
C212 B.n172 VSUBS 0.007242f
C213 B.n173 VSUBS 0.007242f
C214 B.n174 VSUBS 0.007242f
C215 B.n175 VSUBS 0.007242f
C216 B.n176 VSUBS 0.007242f
C217 B.n177 VSUBS 0.007242f
C218 B.n178 VSUBS 0.007242f
C219 B.n179 VSUBS 0.007242f
C220 B.n180 VSUBS 0.007242f
C221 B.n181 VSUBS 0.007242f
C222 B.n182 VSUBS 0.007242f
C223 B.n183 VSUBS 0.007242f
C224 B.n184 VSUBS 0.007242f
C225 B.n185 VSUBS 0.007242f
C226 B.n186 VSUBS 0.007242f
C227 B.n187 VSUBS 0.017789f
C228 B.n188 VSUBS 0.017789f
C229 B.n189 VSUBS 0.018632f
C230 B.n190 VSUBS 0.007242f
C231 B.n191 VSUBS 0.007242f
C232 B.n192 VSUBS 0.007242f
C233 B.n193 VSUBS 0.007242f
C234 B.n194 VSUBS 0.007242f
C235 B.n195 VSUBS 0.007242f
C236 B.n196 VSUBS 0.007242f
C237 B.n197 VSUBS 0.007242f
C238 B.n198 VSUBS 0.007242f
C239 B.n199 VSUBS 0.007242f
C240 B.n200 VSUBS 0.007242f
C241 B.n201 VSUBS 0.007242f
C242 B.n202 VSUBS 0.007242f
C243 B.n203 VSUBS 0.007242f
C244 B.n204 VSUBS 0.007242f
C245 B.n205 VSUBS 0.007242f
C246 B.n206 VSUBS 0.007242f
C247 B.n207 VSUBS 0.007242f
C248 B.n208 VSUBS 0.007242f
C249 B.n209 VSUBS 0.007242f
C250 B.n210 VSUBS 0.007242f
C251 B.n211 VSUBS 0.007242f
C252 B.n212 VSUBS 0.007242f
C253 B.n213 VSUBS 0.007242f
C254 B.n214 VSUBS 0.007242f
C255 B.n215 VSUBS 0.007242f
C256 B.n216 VSUBS 0.007242f
C257 B.n217 VSUBS 0.007242f
C258 B.n218 VSUBS 0.007242f
C259 B.n219 VSUBS 0.007242f
C260 B.n220 VSUBS 0.007242f
C261 B.n221 VSUBS 0.007242f
C262 B.n222 VSUBS 0.007242f
C263 B.n223 VSUBS 0.007242f
C264 B.n224 VSUBS 0.007242f
C265 B.n225 VSUBS 0.007242f
C266 B.n226 VSUBS 0.007242f
C267 B.n227 VSUBS 0.007242f
C268 B.n228 VSUBS 0.007242f
C269 B.n229 VSUBS 0.007242f
C270 B.n230 VSUBS 0.007242f
C271 B.n231 VSUBS 0.007242f
C272 B.n232 VSUBS 0.007242f
C273 B.n233 VSUBS 0.007242f
C274 B.n234 VSUBS 0.007242f
C275 B.n235 VSUBS 0.006816f
C276 B.n236 VSUBS 0.007242f
C277 B.n237 VSUBS 0.007242f
C278 B.n238 VSUBS 0.004047f
C279 B.n239 VSUBS 0.007242f
C280 B.n240 VSUBS 0.007242f
C281 B.n241 VSUBS 0.007242f
C282 B.n242 VSUBS 0.007242f
C283 B.n243 VSUBS 0.007242f
C284 B.n244 VSUBS 0.007242f
C285 B.n245 VSUBS 0.007242f
C286 B.n246 VSUBS 0.007242f
C287 B.n247 VSUBS 0.007242f
C288 B.n248 VSUBS 0.007242f
C289 B.n249 VSUBS 0.007242f
C290 B.n250 VSUBS 0.007242f
C291 B.n251 VSUBS 0.004047f
C292 B.n252 VSUBS 0.016778f
C293 B.n253 VSUBS 0.006816f
C294 B.n254 VSUBS 0.007242f
C295 B.n255 VSUBS 0.007242f
C296 B.n256 VSUBS 0.007242f
C297 B.n257 VSUBS 0.007242f
C298 B.n258 VSUBS 0.007242f
C299 B.n259 VSUBS 0.007242f
C300 B.n260 VSUBS 0.007242f
C301 B.n261 VSUBS 0.007242f
C302 B.n262 VSUBS 0.007242f
C303 B.n263 VSUBS 0.007242f
C304 B.n264 VSUBS 0.007242f
C305 B.n265 VSUBS 0.007242f
C306 B.n266 VSUBS 0.007242f
C307 B.n267 VSUBS 0.007242f
C308 B.n268 VSUBS 0.007242f
C309 B.n269 VSUBS 0.007242f
C310 B.n270 VSUBS 0.007242f
C311 B.n271 VSUBS 0.007242f
C312 B.n272 VSUBS 0.007242f
C313 B.n273 VSUBS 0.007242f
C314 B.n274 VSUBS 0.007242f
C315 B.n275 VSUBS 0.007242f
C316 B.n276 VSUBS 0.007242f
C317 B.n277 VSUBS 0.007242f
C318 B.n278 VSUBS 0.007242f
C319 B.n279 VSUBS 0.007242f
C320 B.n280 VSUBS 0.007242f
C321 B.n281 VSUBS 0.007242f
C322 B.n282 VSUBS 0.007242f
C323 B.n283 VSUBS 0.007242f
C324 B.n284 VSUBS 0.007242f
C325 B.n285 VSUBS 0.007242f
C326 B.n286 VSUBS 0.007242f
C327 B.n287 VSUBS 0.007242f
C328 B.n288 VSUBS 0.007242f
C329 B.n289 VSUBS 0.007242f
C330 B.n290 VSUBS 0.007242f
C331 B.n291 VSUBS 0.007242f
C332 B.n292 VSUBS 0.007242f
C333 B.n293 VSUBS 0.007242f
C334 B.n294 VSUBS 0.007242f
C335 B.n295 VSUBS 0.007242f
C336 B.n296 VSUBS 0.007242f
C337 B.n297 VSUBS 0.007242f
C338 B.n298 VSUBS 0.007242f
C339 B.n299 VSUBS 0.007242f
C340 B.n300 VSUBS 0.018632f
C341 B.n301 VSUBS 0.017789f
C342 B.n302 VSUBS 0.017789f
C343 B.n303 VSUBS 0.007242f
C344 B.n304 VSUBS 0.007242f
C345 B.n305 VSUBS 0.007242f
C346 B.n306 VSUBS 0.007242f
C347 B.n307 VSUBS 0.007242f
C348 B.n308 VSUBS 0.007242f
C349 B.n309 VSUBS 0.007242f
C350 B.n310 VSUBS 0.007242f
C351 B.n311 VSUBS 0.007242f
C352 B.n312 VSUBS 0.007242f
C353 B.n313 VSUBS 0.007242f
C354 B.n314 VSUBS 0.007242f
C355 B.n315 VSUBS 0.007242f
C356 B.n316 VSUBS 0.007242f
C357 B.n317 VSUBS 0.007242f
C358 B.n318 VSUBS 0.007242f
C359 B.n319 VSUBS 0.007242f
C360 B.n320 VSUBS 0.007242f
C361 B.n321 VSUBS 0.007242f
C362 B.n322 VSUBS 0.007242f
C363 B.n323 VSUBS 0.007242f
C364 B.n324 VSUBS 0.007242f
C365 B.n325 VSUBS 0.007242f
C366 B.n326 VSUBS 0.007242f
C367 B.n327 VSUBS 0.007242f
C368 B.n328 VSUBS 0.007242f
C369 B.n329 VSUBS 0.007242f
C370 B.n330 VSUBS 0.007242f
C371 B.n331 VSUBS 0.007242f
C372 B.n332 VSUBS 0.007242f
C373 B.n333 VSUBS 0.007242f
C374 B.n334 VSUBS 0.007242f
C375 B.n335 VSUBS 0.007242f
C376 B.n336 VSUBS 0.007242f
C377 B.n337 VSUBS 0.007242f
C378 B.n338 VSUBS 0.007242f
C379 B.n339 VSUBS 0.007242f
C380 B.n340 VSUBS 0.007242f
C381 B.n341 VSUBS 0.007242f
C382 B.n342 VSUBS 0.007242f
C383 B.n343 VSUBS 0.007242f
C384 B.n344 VSUBS 0.007242f
C385 B.n345 VSUBS 0.007242f
C386 B.n346 VSUBS 0.007242f
C387 B.n347 VSUBS 0.007242f
C388 B.n348 VSUBS 0.007242f
C389 B.n349 VSUBS 0.007242f
C390 B.n350 VSUBS 0.007242f
C391 B.n351 VSUBS 0.007242f
C392 B.n352 VSUBS 0.007242f
C393 B.n353 VSUBS 0.007242f
C394 B.n354 VSUBS 0.007242f
C395 B.n355 VSUBS 0.007242f
C396 B.n356 VSUBS 0.007242f
C397 B.n357 VSUBS 0.007242f
C398 B.n358 VSUBS 0.007242f
C399 B.n359 VSUBS 0.007242f
C400 B.n360 VSUBS 0.007242f
C401 B.n361 VSUBS 0.007242f
C402 B.n362 VSUBS 0.007242f
C403 B.n363 VSUBS 0.007242f
C404 B.n364 VSUBS 0.007242f
C405 B.n365 VSUBS 0.007242f
C406 B.n366 VSUBS 0.007242f
C407 B.n367 VSUBS 0.007242f
C408 B.n368 VSUBS 0.007242f
C409 B.n369 VSUBS 0.007242f
C410 B.n370 VSUBS 0.007242f
C411 B.n371 VSUBS 0.007242f
C412 B.n372 VSUBS 0.007242f
C413 B.n373 VSUBS 0.007242f
C414 B.n374 VSUBS 0.007242f
C415 B.n375 VSUBS 0.007242f
C416 B.n376 VSUBS 0.007242f
C417 B.n377 VSUBS 0.007242f
C418 B.n378 VSUBS 0.007242f
C419 B.n379 VSUBS 0.007242f
C420 B.n380 VSUBS 0.007242f
C421 B.n381 VSUBS 0.007242f
C422 B.n382 VSUBS 0.007242f
C423 B.n383 VSUBS 0.007242f
C424 B.n384 VSUBS 0.007242f
C425 B.n385 VSUBS 0.007242f
C426 B.n386 VSUBS 0.007242f
C427 B.n387 VSUBS 0.007242f
C428 B.n388 VSUBS 0.007242f
C429 B.n389 VSUBS 0.007242f
C430 B.n390 VSUBS 0.007242f
C431 B.n391 VSUBS 0.018557f
C432 B.n392 VSUBS 0.017789f
C433 B.n393 VSUBS 0.018632f
C434 B.n394 VSUBS 0.007242f
C435 B.n395 VSUBS 0.007242f
C436 B.n396 VSUBS 0.007242f
C437 B.n397 VSUBS 0.007242f
C438 B.n398 VSUBS 0.007242f
C439 B.n399 VSUBS 0.007242f
C440 B.n400 VSUBS 0.007242f
C441 B.n401 VSUBS 0.007242f
C442 B.n402 VSUBS 0.007242f
C443 B.n403 VSUBS 0.007242f
C444 B.n404 VSUBS 0.007242f
C445 B.n405 VSUBS 0.007242f
C446 B.n406 VSUBS 0.007242f
C447 B.n407 VSUBS 0.007242f
C448 B.n408 VSUBS 0.007242f
C449 B.n409 VSUBS 0.007242f
C450 B.n410 VSUBS 0.007242f
C451 B.n411 VSUBS 0.007242f
C452 B.n412 VSUBS 0.007242f
C453 B.n413 VSUBS 0.007242f
C454 B.n414 VSUBS 0.007242f
C455 B.n415 VSUBS 0.007242f
C456 B.n416 VSUBS 0.007242f
C457 B.n417 VSUBS 0.007242f
C458 B.n418 VSUBS 0.007242f
C459 B.n419 VSUBS 0.007242f
C460 B.n420 VSUBS 0.007242f
C461 B.n421 VSUBS 0.007242f
C462 B.n422 VSUBS 0.007242f
C463 B.n423 VSUBS 0.007242f
C464 B.n424 VSUBS 0.007242f
C465 B.n425 VSUBS 0.007242f
C466 B.n426 VSUBS 0.007242f
C467 B.n427 VSUBS 0.007242f
C468 B.n428 VSUBS 0.007242f
C469 B.n429 VSUBS 0.007242f
C470 B.n430 VSUBS 0.007242f
C471 B.n431 VSUBS 0.007242f
C472 B.n432 VSUBS 0.007242f
C473 B.n433 VSUBS 0.007242f
C474 B.n434 VSUBS 0.007242f
C475 B.n435 VSUBS 0.007242f
C476 B.n436 VSUBS 0.007242f
C477 B.n437 VSUBS 0.007242f
C478 B.n438 VSUBS 0.007242f
C479 B.n439 VSUBS 0.006816f
C480 B.n440 VSUBS 0.007242f
C481 B.n441 VSUBS 0.007242f
C482 B.n442 VSUBS 0.004047f
C483 B.n443 VSUBS 0.007242f
C484 B.n444 VSUBS 0.007242f
C485 B.n445 VSUBS 0.007242f
C486 B.n446 VSUBS 0.007242f
C487 B.n447 VSUBS 0.007242f
C488 B.n448 VSUBS 0.007242f
C489 B.n449 VSUBS 0.007242f
C490 B.n450 VSUBS 0.007242f
C491 B.n451 VSUBS 0.007242f
C492 B.n452 VSUBS 0.007242f
C493 B.n453 VSUBS 0.007242f
C494 B.n454 VSUBS 0.007242f
C495 B.n455 VSUBS 0.004047f
C496 B.n456 VSUBS 0.016778f
C497 B.n457 VSUBS 0.006816f
C498 B.n458 VSUBS 0.007242f
C499 B.n459 VSUBS 0.007242f
C500 B.n460 VSUBS 0.007242f
C501 B.n461 VSUBS 0.007242f
C502 B.n462 VSUBS 0.007242f
C503 B.n463 VSUBS 0.007242f
C504 B.n464 VSUBS 0.007242f
C505 B.n465 VSUBS 0.007242f
C506 B.n466 VSUBS 0.007242f
C507 B.n467 VSUBS 0.007242f
C508 B.n468 VSUBS 0.007242f
C509 B.n469 VSUBS 0.007242f
C510 B.n470 VSUBS 0.007242f
C511 B.n471 VSUBS 0.007242f
C512 B.n472 VSUBS 0.007242f
C513 B.n473 VSUBS 0.007242f
C514 B.n474 VSUBS 0.007242f
C515 B.n475 VSUBS 0.007242f
C516 B.n476 VSUBS 0.007242f
C517 B.n477 VSUBS 0.007242f
C518 B.n478 VSUBS 0.007242f
C519 B.n479 VSUBS 0.007242f
C520 B.n480 VSUBS 0.007242f
C521 B.n481 VSUBS 0.007242f
C522 B.n482 VSUBS 0.007242f
C523 B.n483 VSUBS 0.007242f
C524 B.n484 VSUBS 0.007242f
C525 B.n485 VSUBS 0.007242f
C526 B.n486 VSUBS 0.007242f
C527 B.n487 VSUBS 0.007242f
C528 B.n488 VSUBS 0.007242f
C529 B.n489 VSUBS 0.007242f
C530 B.n490 VSUBS 0.007242f
C531 B.n491 VSUBS 0.007242f
C532 B.n492 VSUBS 0.007242f
C533 B.n493 VSUBS 0.007242f
C534 B.n494 VSUBS 0.007242f
C535 B.n495 VSUBS 0.007242f
C536 B.n496 VSUBS 0.007242f
C537 B.n497 VSUBS 0.007242f
C538 B.n498 VSUBS 0.007242f
C539 B.n499 VSUBS 0.007242f
C540 B.n500 VSUBS 0.007242f
C541 B.n501 VSUBS 0.007242f
C542 B.n502 VSUBS 0.007242f
C543 B.n503 VSUBS 0.007242f
C544 B.n504 VSUBS 0.018632f
C545 B.n505 VSUBS 0.017789f
C546 B.n506 VSUBS 0.017789f
C547 B.n507 VSUBS 0.007242f
C548 B.n508 VSUBS 0.007242f
C549 B.n509 VSUBS 0.007242f
C550 B.n510 VSUBS 0.007242f
C551 B.n511 VSUBS 0.007242f
C552 B.n512 VSUBS 0.007242f
C553 B.n513 VSUBS 0.007242f
C554 B.n514 VSUBS 0.007242f
C555 B.n515 VSUBS 0.007242f
C556 B.n516 VSUBS 0.007242f
C557 B.n517 VSUBS 0.007242f
C558 B.n518 VSUBS 0.007242f
C559 B.n519 VSUBS 0.007242f
C560 B.n520 VSUBS 0.007242f
C561 B.n521 VSUBS 0.007242f
C562 B.n522 VSUBS 0.007242f
C563 B.n523 VSUBS 0.007242f
C564 B.n524 VSUBS 0.007242f
C565 B.n525 VSUBS 0.007242f
C566 B.n526 VSUBS 0.007242f
C567 B.n527 VSUBS 0.007242f
C568 B.n528 VSUBS 0.007242f
C569 B.n529 VSUBS 0.007242f
C570 B.n530 VSUBS 0.007242f
C571 B.n531 VSUBS 0.007242f
C572 B.n532 VSUBS 0.007242f
C573 B.n533 VSUBS 0.007242f
C574 B.n534 VSUBS 0.007242f
C575 B.n535 VSUBS 0.007242f
C576 B.n536 VSUBS 0.007242f
C577 B.n537 VSUBS 0.007242f
C578 B.n538 VSUBS 0.007242f
C579 B.n539 VSUBS 0.007242f
C580 B.n540 VSUBS 0.007242f
C581 B.n541 VSUBS 0.007242f
C582 B.n542 VSUBS 0.007242f
C583 B.n543 VSUBS 0.007242f
C584 B.n544 VSUBS 0.007242f
C585 B.n545 VSUBS 0.007242f
C586 B.n546 VSUBS 0.007242f
C587 B.n547 VSUBS 0.007242f
C588 B.n548 VSUBS 0.007242f
C589 B.n549 VSUBS 0.007242f
C590 B.n550 VSUBS 0.007242f
C591 B.n551 VSUBS 0.016398f
C592 VDD2.t3 VSUBS 1.49352f
C593 VDD2.t0 VSUBS 0.153476f
C594 VDD2.t4 VSUBS 0.153476f
C595 VDD2.n0 VSUBS 1.13192f
C596 VDD2.n1 VSUBS 2.39996f
C597 VDD2.t1 VSUBS 1.48604f
C598 VDD2.n2 VSUBS 2.19588f
C599 VDD2.t5 VSUBS 0.153476f
C600 VDD2.t2 VSUBS 0.153476f
C601 VDD2.n3 VSUBS 1.1319f
C602 VN.n0 VSUBS 0.04264f
C603 VN.t1 VSUBS 1.57747f
C604 VN.n1 VSUBS 0.055118f
C605 VN.t2 VSUBS 1.71894f
C606 VN.n2 VSUBS 0.686497f
C607 VN.t5 VSUBS 1.57747f
C608 VN.n3 VSUBS 0.666737f
C609 VN.n4 VSUBS 0.059853f
C610 VN.n5 VSUBS 0.268953f
C611 VN.n6 VSUBS 0.04264f
C612 VN.n7 VSUBS 0.04264f
C613 VN.n8 VSUBS 0.069376f
C614 VN.n9 VSUBS 0.050437f
C615 VN.n10 VSUBS 0.669789f
C616 VN.n11 VSUBS 0.04249f
C617 VN.n12 VSUBS 0.04264f
C618 VN.t4 VSUBS 1.57747f
C619 VN.n13 VSUBS 0.055118f
C620 VN.t3 VSUBS 1.71894f
C621 VN.n14 VSUBS 0.686497f
C622 VN.t0 VSUBS 1.57747f
C623 VN.n15 VSUBS 0.666737f
C624 VN.n16 VSUBS 0.059853f
C625 VN.n17 VSUBS 0.268953f
C626 VN.n18 VSUBS 0.04264f
C627 VN.n19 VSUBS 0.04264f
C628 VN.n20 VSUBS 0.069376f
C629 VN.n21 VSUBS 0.050437f
C630 VN.n22 VSUBS 0.669789f
C631 VN.n23 VSUBS 1.80123f
C632 VTAIL.t1 VSUBS 0.207587f
C633 VTAIL.t0 VSUBS 0.207587f
C634 VTAIL.n0 VSUBS 1.38896f
C635 VTAIL.n1 VSUBS 0.788197f
C636 VTAIL.t6 VSUBS 1.85759f
C637 VTAIL.n2 VSUBS 0.996408f
C638 VTAIL.t4 VSUBS 0.207587f
C639 VTAIL.t9 VSUBS 0.207587f
C640 VTAIL.n3 VSUBS 1.38896f
C641 VTAIL.n4 VSUBS 2.21937f
C642 VTAIL.t3 VSUBS 0.207587f
C643 VTAIL.t10 VSUBS 0.207587f
C644 VTAIL.n5 VSUBS 1.38897f
C645 VTAIL.n6 VSUBS 2.21936f
C646 VTAIL.t2 VSUBS 1.8576f
C647 VTAIL.n7 VSUBS 0.996402f
C648 VTAIL.t8 VSUBS 0.207587f
C649 VTAIL.t5 VSUBS 0.207587f
C650 VTAIL.n8 VSUBS 1.38897f
C651 VTAIL.n9 VSUBS 0.898883f
C652 VTAIL.t7 VSUBS 1.85759f
C653 VTAIL.n10 VSUBS 2.16188f
C654 VTAIL.t11 VSUBS 1.85759f
C655 VTAIL.n11 VSUBS 2.11756f
C656 VDD1.t2 VSUBS 1.49689f
C657 VDD1.t0 VSUBS 1.49605f
C658 VDD1.t5 VSUBS 0.153736f
C659 VDD1.t1 VSUBS 0.153736f
C660 VDD1.n0 VSUBS 1.13384f
C661 VDD1.n1 VSUBS 2.48801f
C662 VDD1.t3 VSUBS 0.153736f
C663 VDD1.t4 VSUBS 0.153736f
C664 VDD1.n2 VSUBS 1.13147f
C665 VDD1.n3 VSUBS 2.18378f
C666 VP.n0 VSUBS 0.043921f
C667 VP.t3 VSUBS 1.62486f
C668 VP.n1 VSUBS 0.056774f
C669 VP.n2 VSUBS 0.043921f
C670 VP.t0 VSUBS 1.62486f
C671 VP.n3 VSUBS 0.071461f
C672 VP.n4 VSUBS 0.043921f
C673 VP.t2 VSUBS 1.62486f
C674 VP.n5 VSUBS 0.056774f
C675 VP.t1 VSUBS 1.77057f
C676 VP.n6 VSUBS 0.707119f
C677 VP.t4 VSUBS 1.62486f
C678 VP.n7 VSUBS 0.686765f
C679 VP.n8 VSUBS 0.061651f
C680 VP.n9 VSUBS 0.277032f
C681 VP.n10 VSUBS 0.043921f
C682 VP.n11 VSUBS 0.043921f
C683 VP.n12 VSUBS 0.071461f
C684 VP.n13 VSUBS 0.051952f
C685 VP.n14 VSUBS 0.68991f
C686 VP.n15 VSUBS 1.82651f
C687 VP.n16 VSUBS 1.86405f
C688 VP.t5 VSUBS 1.62486f
C689 VP.n17 VSUBS 0.68991f
C690 VP.n18 VSUBS 0.051952f
C691 VP.n19 VSUBS 0.043921f
C692 VP.n20 VSUBS 0.043921f
C693 VP.n21 VSUBS 0.043921f
C694 VP.n22 VSUBS 0.056774f
C695 VP.n23 VSUBS 0.061651f
C696 VP.n24 VSUBS 0.603232f
C697 VP.n25 VSUBS 0.061651f
C698 VP.n26 VSUBS 0.043921f
C699 VP.n27 VSUBS 0.043921f
C700 VP.n28 VSUBS 0.043921f
C701 VP.n29 VSUBS 0.071461f
C702 VP.n30 VSUBS 0.051952f
C703 VP.n31 VSUBS 0.68991f
C704 VP.n32 VSUBS 0.043767f
.ends

