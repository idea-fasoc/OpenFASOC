* NGSPICE file created from diff_pair_sample_0797.ext - technology: sky130A

.subckt diff_pair_sample_0797 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X1 VDD1.t9 VP.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=1.2375 ps=7.83 w=7.5 l=1.3
X2 VTAIL.t3 VP.t1 VDD1.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X3 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=1.3
X4 VDD2.t7 VN.t1 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=2.925 ps=15.78 w=7.5 l=1.3
X5 VDD2.t1 VN.t2 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X6 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X7 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X8 VTAIL.t16 VN.t3 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X9 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=1.3
X10 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=2.925 ps=15.78 w=7.5 l=1.3
X11 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=1.3
X12 VTAIL.t1 VP.t5 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X13 VDD2.t0 VN.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=1.2375 ps=7.83 w=7.5 l=1.3
X14 VDD2.t6 VN.t5 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=1.2375 ps=7.83 w=7.5 l=1.3
X15 VDD1.t3 VP.t6 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=2.925 ps=15.78 w=7.5 l=1.3
X16 VTAIL.t7 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X17 VDD1.t1 VP.t8 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=1.2375 ps=7.83 w=7.5 l=1.3
X18 VDD2.t5 VN.t6 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=2.925 ps=15.78 w=7.5 l=1.3
X19 VTAIL.t12 VN.t7 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=1.3
X21 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X22 VTAIL.t11 VN.t8 VDD2.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
X23 VDD2.t2 VN.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=1.2375 ps=7.83 w=7.5 l=1.3
R0 VN.n24 VN.n23 173.105
R1 VN.n49 VN.n48 173.105
R2 VN.n6 VN.t5 168.714
R3 VN.n32 VN.t6 168.714
R4 VN.n47 VN.n25 161.3
R5 VN.n46 VN.n45 161.3
R6 VN.n44 VN.n26 161.3
R7 VN.n43 VN.n42 161.3
R8 VN.n41 VN.n27 161.3
R9 VN.n40 VN.n39 161.3
R10 VN.n38 VN.n29 161.3
R11 VN.n37 VN.n36 161.3
R12 VN.n35 VN.n30 161.3
R13 VN.n34 VN.n33 161.3
R14 VN.n22 VN.n0 161.3
R15 VN.n21 VN.n20 161.3
R16 VN.n19 VN.n1 161.3
R17 VN.n18 VN.n17 161.3
R18 VN.n15 VN.n2 161.3
R19 VN.n14 VN.n13 161.3
R20 VN.n12 VN.n3 161.3
R21 VN.n11 VN.n10 161.3
R22 VN.n9 VN.n4 161.3
R23 VN.n8 VN.n7 161.3
R24 VN.n3 VN.t2 139.038
R25 VN.n5 VN.t0 139.038
R26 VN.n16 VN.t7 139.038
R27 VN.n23 VN.t1 139.038
R28 VN.n29 VN.t9 139.038
R29 VN.n31 VN.t3 139.038
R30 VN.n28 VN.t8 139.038
R31 VN.n48 VN.t4 139.038
R32 VN.n6 VN.n5 58.6212
R33 VN.n32 VN.n31 58.6212
R34 VN.n10 VN.n9 56.5617
R35 VN.n15 VN.n14 56.5617
R36 VN.n36 VN.n35 56.5617
R37 VN.n41 VN.n40 56.5617
R38 VN.n21 VN.n1 45.9053
R39 VN.n46 VN.n26 45.9053
R40 VN VN.n49 42.938
R41 VN.n22 VN.n21 35.2488
R42 VN.n47 VN.n46 35.2488
R43 VN.n33 VN.n32 27.0756
R44 VN.n7 VN.n6 27.0756
R45 VN.n9 VN.n8 24.5923
R46 VN.n10 VN.n3 24.5923
R47 VN.n14 VN.n3 24.5923
R48 VN.n17 VN.n15 24.5923
R49 VN.n35 VN.n34 24.5923
R50 VN.n40 VN.n29 24.5923
R51 VN.n36 VN.n29 24.5923
R52 VN.n42 VN.n41 24.5923
R53 VN.n16 VN.n1 18.1985
R54 VN.n28 VN.n26 18.1985
R55 VN.n23 VN.n22 12.7883
R56 VN.n48 VN.n47 12.7883
R57 VN.n8 VN.n5 6.39438
R58 VN.n17 VN.n16 6.39438
R59 VN.n34 VN.n31 6.39438
R60 VN.n42 VN.n28 6.39438
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n30 0.189894
R70 VN.n33 VN.n30 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n11 VN.n4 0.189894
R73 VN.n12 VN.n11 0.189894
R74 VN.n13 VN.n12 0.189894
R75 VN.n13 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VDD2.n1 VDD2.t6 69.4999
R83 VDD2.n4 VDD2.t0 68.0949
R84 VDD2.n3 VDD2.n2 66.4533
R85 VDD2 VDD2.n7 66.4504
R86 VDD2.n6 VDD2.n5 65.4549
R87 VDD2.n1 VDD2.n0 65.4547
R88 VDD2.n4 VDD2.n3 36.8554
R89 VDD2.n7 VDD2.t3 2.6405
R90 VDD2.n7 VDD2.t5 2.6405
R91 VDD2.n5 VDD2.t8 2.6405
R92 VDD2.n5 VDD2.t2 2.6405
R93 VDD2.n2 VDD2.t9 2.6405
R94 VDD2.n2 VDD2.t7 2.6405
R95 VDD2.n0 VDD2.t4 2.6405
R96 VDD2.n0 VDD2.t1 2.6405
R97 VDD2.n6 VDD2.n4 1.40567
R98 VDD2 VDD2.n6 0.409983
R99 VDD2.n3 VDD2.n1 0.296447
R100 VTAIL.n11 VTAIL.t13 51.4161
R101 VTAIL.n17 VTAIL.t18 51.4159
R102 VTAIL.n2 VTAIL.t8 51.4159
R103 VTAIL.n16 VTAIL.t4 51.4159
R104 VTAIL.n15 VTAIL.n14 48.7761
R105 VTAIL.n13 VTAIL.n12 48.7761
R106 VTAIL.n10 VTAIL.n9 48.7761
R107 VTAIL.n8 VTAIL.n7 48.7761
R108 VTAIL.n19 VTAIL.n18 48.7759
R109 VTAIL.n1 VTAIL.n0 48.7759
R110 VTAIL.n4 VTAIL.n3 48.7759
R111 VTAIL.n6 VTAIL.n5 48.7759
R112 VTAIL.n8 VTAIL.n6 21.6427
R113 VTAIL.n17 VTAIL.n16 20.2376
R114 VTAIL.n18 VTAIL.t17 2.6405
R115 VTAIL.n18 VTAIL.t12 2.6405
R116 VTAIL.n0 VTAIL.t14 2.6405
R117 VTAIL.n0 VTAIL.t19 2.6405
R118 VTAIL.n3 VTAIL.t2 2.6405
R119 VTAIL.n3 VTAIL.t3 2.6405
R120 VTAIL.n5 VTAIL.t9 2.6405
R121 VTAIL.n5 VTAIL.t7 2.6405
R122 VTAIL.n14 VTAIL.t0 2.6405
R123 VTAIL.n14 VTAIL.t1 2.6405
R124 VTAIL.n12 VTAIL.t6 2.6405
R125 VTAIL.n12 VTAIL.t5 2.6405
R126 VTAIL.n9 VTAIL.t10 2.6405
R127 VTAIL.n9 VTAIL.t16 2.6405
R128 VTAIL.n7 VTAIL.t15 2.6405
R129 VTAIL.n7 VTAIL.t11 2.6405
R130 VTAIL.n10 VTAIL.n8 1.40567
R131 VTAIL.n11 VTAIL.n10 1.40567
R132 VTAIL.n15 VTAIL.n13 1.40567
R133 VTAIL.n16 VTAIL.n15 1.40567
R134 VTAIL.n6 VTAIL.n4 1.40567
R135 VTAIL.n4 VTAIL.n2 1.40567
R136 VTAIL.n19 VTAIL.n17 1.40567
R137 VTAIL.n13 VTAIL.n11 1.17291
R138 VTAIL.n2 VTAIL.n1 1.17291
R139 VTAIL VTAIL.n1 1.11257
R140 VTAIL VTAIL.n19 0.293603
R141 B.n638 B.n637 585
R142 B.n237 B.n102 585
R143 B.n236 B.n235 585
R144 B.n234 B.n233 585
R145 B.n232 B.n231 585
R146 B.n230 B.n229 585
R147 B.n228 B.n227 585
R148 B.n226 B.n225 585
R149 B.n224 B.n223 585
R150 B.n222 B.n221 585
R151 B.n220 B.n219 585
R152 B.n218 B.n217 585
R153 B.n216 B.n215 585
R154 B.n214 B.n213 585
R155 B.n212 B.n211 585
R156 B.n210 B.n209 585
R157 B.n208 B.n207 585
R158 B.n206 B.n205 585
R159 B.n204 B.n203 585
R160 B.n202 B.n201 585
R161 B.n200 B.n199 585
R162 B.n198 B.n197 585
R163 B.n196 B.n195 585
R164 B.n194 B.n193 585
R165 B.n192 B.n191 585
R166 B.n190 B.n189 585
R167 B.n188 B.n187 585
R168 B.n186 B.n185 585
R169 B.n184 B.n183 585
R170 B.n182 B.n181 585
R171 B.n180 B.n179 585
R172 B.n178 B.n177 585
R173 B.n176 B.n175 585
R174 B.n174 B.n173 585
R175 B.n172 B.n171 585
R176 B.n170 B.n169 585
R177 B.n168 B.n167 585
R178 B.n166 B.n165 585
R179 B.n164 B.n163 585
R180 B.n162 B.n161 585
R181 B.n160 B.n159 585
R182 B.n158 B.n157 585
R183 B.n156 B.n155 585
R184 B.n154 B.n153 585
R185 B.n152 B.n151 585
R186 B.n150 B.n149 585
R187 B.n148 B.n147 585
R188 B.n146 B.n145 585
R189 B.n144 B.n143 585
R190 B.n142 B.n141 585
R191 B.n140 B.n139 585
R192 B.n138 B.n137 585
R193 B.n136 B.n135 585
R194 B.n134 B.n133 585
R195 B.n132 B.n131 585
R196 B.n130 B.n129 585
R197 B.n128 B.n127 585
R198 B.n126 B.n125 585
R199 B.n124 B.n123 585
R200 B.n122 B.n121 585
R201 B.n120 B.n119 585
R202 B.n118 B.n117 585
R203 B.n116 B.n115 585
R204 B.n114 B.n113 585
R205 B.n112 B.n111 585
R206 B.n110 B.n109 585
R207 B.n636 B.n69 585
R208 B.n641 B.n69 585
R209 B.n635 B.n68 585
R210 B.n642 B.n68 585
R211 B.n634 B.n633 585
R212 B.n633 B.n64 585
R213 B.n632 B.n63 585
R214 B.n648 B.n63 585
R215 B.n631 B.n62 585
R216 B.n649 B.n62 585
R217 B.n630 B.n61 585
R218 B.n650 B.n61 585
R219 B.n629 B.n628 585
R220 B.n628 B.n57 585
R221 B.n627 B.n56 585
R222 B.n656 B.n56 585
R223 B.n626 B.n55 585
R224 B.n657 B.n55 585
R225 B.n625 B.n54 585
R226 B.n658 B.n54 585
R227 B.n624 B.n623 585
R228 B.n623 B.n50 585
R229 B.n622 B.n49 585
R230 B.n664 B.n49 585
R231 B.n621 B.n48 585
R232 B.n665 B.n48 585
R233 B.n620 B.n47 585
R234 B.n666 B.n47 585
R235 B.n619 B.n618 585
R236 B.n618 B.n43 585
R237 B.n617 B.n42 585
R238 B.n672 B.n42 585
R239 B.n616 B.n41 585
R240 B.n673 B.n41 585
R241 B.n615 B.n40 585
R242 B.n674 B.n40 585
R243 B.n614 B.n613 585
R244 B.n613 B.n39 585
R245 B.n612 B.n35 585
R246 B.n680 B.n35 585
R247 B.n611 B.n34 585
R248 B.n681 B.n34 585
R249 B.n610 B.n33 585
R250 B.n682 B.n33 585
R251 B.n609 B.n608 585
R252 B.n608 B.n29 585
R253 B.n607 B.n28 585
R254 B.n688 B.n28 585
R255 B.n606 B.n27 585
R256 B.n689 B.n27 585
R257 B.n605 B.n26 585
R258 B.n690 B.n26 585
R259 B.n604 B.n603 585
R260 B.n603 B.n22 585
R261 B.n602 B.n21 585
R262 B.n696 B.n21 585
R263 B.n601 B.n20 585
R264 B.n697 B.n20 585
R265 B.n600 B.n19 585
R266 B.n698 B.n19 585
R267 B.n599 B.n598 585
R268 B.n598 B.n15 585
R269 B.n597 B.n14 585
R270 B.n704 B.n14 585
R271 B.n596 B.n13 585
R272 B.n705 B.n13 585
R273 B.n595 B.n12 585
R274 B.t6 B.n12 585
R275 B.n594 B.n593 585
R276 B.n593 B.n8 585
R277 B.n592 B.n7 585
R278 B.n711 B.n7 585
R279 B.n591 B.n6 585
R280 B.n712 B.n6 585
R281 B.n590 B.n5 585
R282 B.n713 B.n5 585
R283 B.n589 B.n588 585
R284 B.n588 B.n4 585
R285 B.n587 B.n238 585
R286 B.n587 B.n586 585
R287 B.n578 B.n239 585
R288 B.n240 B.n239 585
R289 B.n580 B.n579 585
R290 B.t8 B.n580 585
R291 B.n577 B.n245 585
R292 B.n245 B.n244 585
R293 B.n576 B.n575 585
R294 B.n575 B.n574 585
R295 B.n247 B.n246 585
R296 B.n248 B.n247 585
R297 B.n567 B.n566 585
R298 B.n568 B.n567 585
R299 B.n565 B.n252 585
R300 B.n256 B.n252 585
R301 B.n564 B.n563 585
R302 B.n563 B.n562 585
R303 B.n254 B.n253 585
R304 B.n255 B.n254 585
R305 B.n555 B.n554 585
R306 B.n556 B.n555 585
R307 B.n553 B.n261 585
R308 B.n261 B.n260 585
R309 B.n552 B.n551 585
R310 B.n551 B.n550 585
R311 B.n263 B.n262 585
R312 B.n264 B.n263 585
R313 B.n543 B.n542 585
R314 B.n544 B.n543 585
R315 B.n541 B.n269 585
R316 B.n269 B.n268 585
R317 B.n540 B.n539 585
R318 B.n539 B.n538 585
R319 B.n271 B.n270 585
R320 B.n531 B.n271 585
R321 B.n530 B.n529 585
R322 B.n532 B.n530 585
R323 B.n528 B.n276 585
R324 B.n276 B.n275 585
R325 B.n527 B.n526 585
R326 B.n526 B.n525 585
R327 B.n278 B.n277 585
R328 B.n279 B.n278 585
R329 B.n518 B.n517 585
R330 B.n519 B.n518 585
R331 B.n516 B.n284 585
R332 B.n284 B.n283 585
R333 B.n515 B.n514 585
R334 B.n514 B.n513 585
R335 B.n286 B.n285 585
R336 B.n287 B.n286 585
R337 B.n506 B.n505 585
R338 B.n507 B.n506 585
R339 B.n504 B.n292 585
R340 B.n292 B.n291 585
R341 B.n503 B.n502 585
R342 B.n502 B.n501 585
R343 B.n294 B.n293 585
R344 B.n295 B.n294 585
R345 B.n494 B.n493 585
R346 B.n495 B.n494 585
R347 B.n492 B.n300 585
R348 B.n300 B.n299 585
R349 B.n491 B.n490 585
R350 B.n490 B.n489 585
R351 B.n302 B.n301 585
R352 B.n303 B.n302 585
R353 B.n482 B.n481 585
R354 B.n483 B.n482 585
R355 B.n480 B.n308 585
R356 B.n308 B.n307 585
R357 B.n475 B.n474 585
R358 B.n473 B.n343 585
R359 B.n472 B.n342 585
R360 B.n477 B.n342 585
R361 B.n471 B.n470 585
R362 B.n469 B.n468 585
R363 B.n467 B.n466 585
R364 B.n465 B.n464 585
R365 B.n463 B.n462 585
R366 B.n461 B.n460 585
R367 B.n459 B.n458 585
R368 B.n457 B.n456 585
R369 B.n455 B.n454 585
R370 B.n453 B.n452 585
R371 B.n451 B.n450 585
R372 B.n449 B.n448 585
R373 B.n447 B.n446 585
R374 B.n445 B.n444 585
R375 B.n443 B.n442 585
R376 B.n441 B.n440 585
R377 B.n439 B.n438 585
R378 B.n437 B.n436 585
R379 B.n435 B.n434 585
R380 B.n433 B.n432 585
R381 B.n431 B.n430 585
R382 B.n429 B.n428 585
R383 B.n427 B.n426 585
R384 B.n425 B.n424 585
R385 B.n423 B.n422 585
R386 B.n420 B.n419 585
R387 B.n418 B.n417 585
R388 B.n416 B.n415 585
R389 B.n414 B.n413 585
R390 B.n412 B.n411 585
R391 B.n410 B.n409 585
R392 B.n408 B.n407 585
R393 B.n406 B.n405 585
R394 B.n404 B.n403 585
R395 B.n402 B.n401 585
R396 B.n399 B.n398 585
R397 B.n397 B.n396 585
R398 B.n395 B.n394 585
R399 B.n393 B.n392 585
R400 B.n391 B.n390 585
R401 B.n389 B.n388 585
R402 B.n387 B.n386 585
R403 B.n385 B.n384 585
R404 B.n383 B.n382 585
R405 B.n381 B.n380 585
R406 B.n379 B.n378 585
R407 B.n377 B.n376 585
R408 B.n375 B.n374 585
R409 B.n373 B.n372 585
R410 B.n371 B.n370 585
R411 B.n369 B.n368 585
R412 B.n367 B.n366 585
R413 B.n365 B.n364 585
R414 B.n363 B.n362 585
R415 B.n361 B.n360 585
R416 B.n359 B.n358 585
R417 B.n357 B.n356 585
R418 B.n355 B.n354 585
R419 B.n353 B.n352 585
R420 B.n351 B.n350 585
R421 B.n349 B.n348 585
R422 B.n310 B.n309 585
R423 B.n479 B.n478 585
R424 B.n478 B.n477 585
R425 B.n306 B.n305 585
R426 B.n307 B.n306 585
R427 B.n485 B.n484 585
R428 B.n484 B.n483 585
R429 B.n486 B.n304 585
R430 B.n304 B.n303 585
R431 B.n488 B.n487 585
R432 B.n489 B.n488 585
R433 B.n298 B.n297 585
R434 B.n299 B.n298 585
R435 B.n497 B.n496 585
R436 B.n496 B.n495 585
R437 B.n498 B.n296 585
R438 B.n296 B.n295 585
R439 B.n500 B.n499 585
R440 B.n501 B.n500 585
R441 B.n290 B.n289 585
R442 B.n291 B.n290 585
R443 B.n509 B.n508 585
R444 B.n508 B.n507 585
R445 B.n510 B.n288 585
R446 B.n288 B.n287 585
R447 B.n512 B.n511 585
R448 B.n513 B.n512 585
R449 B.n282 B.n281 585
R450 B.n283 B.n282 585
R451 B.n521 B.n520 585
R452 B.n520 B.n519 585
R453 B.n522 B.n280 585
R454 B.n280 B.n279 585
R455 B.n524 B.n523 585
R456 B.n525 B.n524 585
R457 B.n274 B.n273 585
R458 B.n275 B.n274 585
R459 B.n534 B.n533 585
R460 B.n533 B.n532 585
R461 B.n535 B.n272 585
R462 B.n531 B.n272 585
R463 B.n537 B.n536 585
R464 B.n538 B.n537 585
R465 B.n267 B.n266 585
R466 B.n268 B.n267 585
R467 B.n546 B.n545 585
R468 B.n545 B.n544 585
R469 B.n547 B.n265 585
R470 B.n265 B.n264 585
R471 B.n549 B.n548 585
R472 B.n550 B.n549 585
R473 B.n259 B.n258 585
R474 B.n260 B.n259 585
R475 B.n558 B.n557 585
R476 B.n557 B.n556 585
R477 B.n559 B.n257 585
R478 B.n257 B.n255 585
R479 B.n561 B.n560 585
R480 B.n562 B.n561 585
R481 B.n251 B.n250 585
R482 B.n256 B.n251 585
R483 B.n570 B.n569 585
R484 B.n569 B.n568 585
R485 B.n571 B.n249 585
R486 B.n249 B.n248 585
R487 B.n573 B.n572 585
R488 B.n574 B.n573 585
R489 B.n243 B.n242 585
R490 B.n244 B.n243 585
R491 B.n582 B.n581 585
R492 B.n581 B.t8 585
R493 B.n583 B.n241 585
R494 B.n241 B.n240 585
R495 B.n585 B.n584 585
R496 B.n586 B.n585 585
R497 B.n2 B.n0 585
R498 B.n4 B.n2 585
R499 B.n3 B.n1 585
R500 B.n712 B.n3 585
R501 B.n710 B.n709 585
R502 B.n711 B.n710 585
R503 B.n708 B.n9 585
R504 B.n9 B.n8 585
R505 B.n707 B.n706 585
R506 B.n706 B.t6 585
R507 B.n11 B.n10 585
R508 B.n705 B.n11 585
R509 B.n703 B.n702 585
R510 B.n704 B.n703 585
R511 B.n701 B.n16 585
R512 B.n16 B.n15 585
R513 B.n700 B.n699 585
R514 B.n699 B.n698 585
R515 B.n18 B.n17 585
R516 B.n697 B.n18 585
R517 B.n695 B.n694 585
R518 B.n696 B.n695 585
R519 B.n693 B.n23 585
R520 B.n23 B.n22 585
R521 B.n692 B.n691 585
R522 B.n691 B.n690 585
R523 B.n25 B.n24 585
R524 B.n689 B.n25 585
R525 B.n687 B.n686 585
R526 B.n688 B.n687 585
R527 B.n685 B.n30 585
R528 B.n30 B.n29 585
R529 B.n684 B.n683 585
R530 B.n683 B.n682 585
R531 B.n32 B.n31 585
R532 B.n681 B.n32 585
R533 B.n679 B.n678 585
R534 B.n680 B.n679 585
R535 B.n677 B.n36 585
R536 B.n39 B.n36 585
R537 B.n676 B.n675 585
R538 B.n675 B.n674 585
R539 B.n38 B.n37 585
R540 B.n673 B.n38 585
R541 B.n671 B.n670 585
R542 B.n672 B.n671 585
R543 B.n669 B.n44 585
R544 B.n44 B.n43 585
R545 B.n668 B.n667 585
R546 B.n667 B.n666 585
R547 B.n46 B.n45 585
R548 B.n665 B.n46 585
R549 B.n663 B.n662 585
R550 B.n664 B.n663 585
R551 B.n661 B.n51 585
R552 B.n51 B.n50 585
R553 B.n660 B.n659 585
R554 B.n659 B.n658 585
R555 B.n53 B.n52 585
R556 B.n657 B.n53 585
R557 B.n655 B.n654 585
R558 B.n656 B.n655 585
R559 B.n653 B.n58 585
R560 B.n58 B.n57 585
R561 B.n652 B.n651 585
R562 B.n651 B.n650 585
R563 B.n60 B.n59 585
R564 B.n649 B.n60 585
R565 B.n647 B.n646 585
R566 B.n648 B.n647 585
R567 B.n645 B.n65 585
R568 B.n65 B.n64 585
R569 B.n644 B.n643 585
R570 B.n643 B.n642 585
R571 B.n67 B.n66 585
R572 B.n641 B.n67 585
R573 B.n715 B.n714 585
R574 B.n714 B.n713 585
R575 B.n475 B.n306 506.916
R576 B.n109 B.n67 506.916
R577 B.n478 B.n308 506.916
R578 B.n638 B.n69 506.916
R579 B.n346 B.t21 343.647
R580 B.n344 B.t10 343.647
R581 B.n106 B.t18 343.647
R582 B.n103 B.t14 343.647
R583 B.n640 B.n639 256.663
R584 B.n640 B.n101 256.663
R585 B.n640 B.n100 256.663
R586 B.n640 B.n99 256.663
R587 B.n640 B.n98 256.663
R588 B.n640 B.n97 256.663
R589 B.n640 B.n96 256.663
R590 B.n640 B.n95 256.663
R591 B.n640 B.n94 256.663
R592 B.n640 B.n93 256.663
R593 B.n640 B.n92 256.663
R594 B.n640 B.n91 256.663
R595 B.n640 B.n90 256.663
R596 B.n640 B.n89 256.663
R597 B.n640 B.n88 256.663
R598 B.n640 B.n87 256.663
R599 B.n640 B.n86 256.663
R600 B.n640 B.n85 256.663
R601 B.n640 B.n84 256.663
R602 B.n640 B.n83 256.663
R603 B.n640 B.n82 256.663
R604 B.n640 B.n81 256.663
R605 B.n640 B.n80 256.663
R606 B.n640 B.n79 256.663
R607 B.n640 B.n78 256.663
R608 B.n640 B.n77 256.663
R609 B.n640 B.n76 256.663
R610 B.n640 B.n75 256.663
R611 B.n640 B.n74 256.663
R612 B.n640 B.n73 256.663
R613 B.n640 B.n72 256.663
R614 B.n640 B.n71 256.663
R615 B.n640 B.n70 256.663
R616 B.n477 B.n476 256.663
R617 B.n477 B.n311 256.663
R618 B.n477 B.n312 256.663
R619 B.n477 B.n313 256.663
R620 B.n477 B.n314 256.663
R621 B.n477 B.n315 256.663
R622 B.n477 B.n316 256.663
R623 B.n477 B.n317 256.663
R624 B.n477 B.n318 256.663
R625 B.n477 B.n319 256.663
R626 B.n477 B.n320 256.663
R627 B.n477 B.n321 256.663
R628 B.n477 B.n322 256.663
R629 B.n477 B.n323 256.663
R630 B.n477 B.n324 256.663
R631 B.n477 B.n325 256.663
R632 B.n477 B.n326 256.663
R633 B.n477 B.n327 256.663
R634 B.n477 B.n328 256.663
R635 B.n477 B.n329 256.663
R636 B.n477 B.n330 256.663
R637 B.n477 B.n331 256.663
R638 B.n477 B.n332 256.663
R639 B.n477 B.n333 256.663
R640 B.n477 B.n334 256.663
R641 B.n477 B.n335 256.663
R642 B.n477 B.n336 256.663
R643 B.n477 B.n337 256.663
R644 B.n477 B.n338 256.663
R645 B.n477 B.n339 256.663
R646 B.n477 B.n340 256.663
R647 B.n477 B.n341 256.663
R648 B.n484 B.n306 163.367
R649 B.n484 B.n304 163.367
R650 B.n488 B.n304 163.367
R651 B.n488 B.n298 163.367
R652 B.n496 B.n298 163.367
R653 B.n496 B.n296 163.367
R654 B.n500 B.n296 163.367
R655 B.n500 B.n290 163.367
R656 B.n508 B.n290 163.367
R657 B.n508 B.n288 163.367
R658 B.n512 B.n288 163.367
R659 B.n512 B.n282 163.367
R660 B.n520 B.n282 163.367
R661 B.n520 B.n280 163.367
R662 B.n524 B.n280 163.367
R663 B.n524 B.n274 163.367
R664 B.n533 B.n274 163.367
R665 B.n533 B.n272 163.367
R666 B.n537 B.n272 163.367
R667 B.n537 B.n267 163.367
R668 B.n545 B.n267 163.367
R669 B.n545 B.n265 163.367
R670 B.n549 B.n265 163.367
R671 B.n549 B.n259 163.367
R672 B.n557 B.n259 163.367
R673 B.n557 B.n257 163.367
R674 B.n561 B.n257 163.367
R675 B.n561 B.n251 163.367
R676 B.n569 B.n251 163.367
R677 B.n569 B.n249 163.367
R678 B.n573 B.n249 163.367
R679 B.n573 B.n243 163.367
R680 B.n581 B.n243 163.367
R681 B.n581 B.n241 163.367
R682 B.n585 B.n241 163.367
R683 B.n585 B.n2 163.367
R684 B.n714 B.n2 163.367
R685 B.n714 B.n3 163.367
R686 B.n710 B.n3 163.367
R687 B.n710 B.n9 163.367
R688 B.n706 B.n9 163.367
R689 B.n706 B.n11 163.367
R690 B.n703 B.n11 163.367
R691 B.n703 B.n16 163.367
R692 B.n699 B.n16 163.367
R693 B.n699 B.n18 163.367
R694 B.n695 B.n18 163.367
R695 B.n695 B.n23 163.367
R696 B.n691 B.n23 163.367
R697 B.n691 B.n25 163.367
R698 B.n687 B.n25 163.367
R699 B.n687 B.n30 163.367
R700 B.n683 B.n30 163.367
R701 B.n683 B.n32 163.367
R702 B.n679 B.n32 163.367
R703 B.n679 B.n36 163.367
R704 B.n675 B.n36 163.367
R705 B.n675 B.n38 163.367
R706 B.n671 B.n38 163.367
R707 B.n671 B.n44 163.367
R708 B.n667 B.n44 163.367
R709 B.n667 B.n46 163.367
R710 B.n663 B.n46 163.367
R711 B.n663 B.n51 163.367
R712 B.n659 B.n51 163.367
R713 B.n659 B.n53 163.367
R714 B.n655 B.n53 163.367
R715 B.n655 B.n58 163.367
R716 B.n651 B.n58 163.367
R717 B.n651 B.n60 163.367
R718 B.n647 B.n60 163.367
R719 B.n647 B.n65 163.367
R720 B.n643 B.n65 163.367
R721 B.n643 B.n67 163.367
R722 B.n343 B.n342 163.367
R723 B.n470 B.n342 163.367
R724 B.n468 B.n467 163.367
R725 B.n464 B.n463 163.367
R726 B.n460 B.n459 163.367
R727 B.n456 B.n455 163.367
R728 B.n452 B.n451 163.367
R729 B.n448 B.n447 163.367
R730 B.n444 B.n443 163.367
R731 B.n440 B.n439 163.367
R732 B.n436 B.n435 163.367
R733 B.n432 B.n431 163.367
R734 B.n428 B.n427 163.367
R735 B.n424 B.n423 163.367
R736 B.n419 B.n418 163.367
R737 B.n415 B.n414 163.367
R738 B.n411 B.n410 163.367
R739 B.n407 B.n406 163.367
R740 B.n403 B.n402 163.367
R741 B.n398 B.n397 163.367
R742 B.n394 B.n393 163.367
R743 B.n390 B.n389 163.367
R744 B.n386 B.n385 163.367
R745 B.n382 B.n381 163.367
R746 B.n378 B.n377 163.367
R747 B.n374 B.n373 163.367
R748 B.n370 B.n369 163.367
R749 B.n366 B.n365 163.367
R750 B.n362 B.n361 163.367
R751 B.n358 B.n357 163.367
R752 B.n354 B.n353 163.367
R753 B.n350 B.n349 163.367
R754 B.n478 B.n310 163.367
R755 B.n482 B.n308 163.367
R756 B.n482 B.n302 163.367
R757 B.n490 B.n302 163.367
R758 B.n490 B.n300 163.367
R759 B.n494 B.n300 163.367
R760 B.n494 B.n294 163.367
R761 B.n502 B.n294 163.367
R762 B.n502 B.n292 163.367
R763 B.n506 B.n292 163.367
R764 B.n506 B.n286 163.367
R765 B.n514 B.n286 163.367
R766 B.n514 B.n284 163.367
R767 B.n518 B.n284 163.367
R768 B.n518 B.n278 163.367
R769 B.n526 B.n278 163.367
R770 B.n526 B.n276 163.367
R771 B.n530 B.n276 163.367
R772 B.n530 B.n271 163.367
R773 B.n539 B.n271 163.367
R774 B.n539 B.n269 163.367
R775 B.n543 B.n269 163.367
R776 B.n543 B.n263 163.367
R777 B.n551 B.n263 163.367
R778 B.n551 B.n261 163.367
R779 B.n555 B.n261 163.367
R780 B.n555 B.n254 163.367
R781 B.n563 B.n254 163.367
R782 B.n563 B.n252 163.367
R783 B.n567 B.n252 163.367
R784 B.n567 B.n247 163.367
R785 B.n575 B.n247 163.367
R786 B.n575 B.n245 163.367
R787 B.n580 B.n245 163.367
R788 B.n580 B.n239 163.367
R789 B.n587 B.n239 163.367
R790 B.n588 B.n587 163.367
R791 B.n588 B.n5 163.367
R792 B.n6 B.n5 163.367
R793 B.n7 B.n6 163.367
R794 B.n593 B.n7 163.367
R795 B.n593 B.n12 163.367
R796 B.n13 B.n12 163.367
R797 B.n14 B.n13 163.367
R798 B.n598 B.n14 163.367
R799 B.n598 B.n19 163.367
R800 B.n20 B.n19 163.367
R801 B.n21 B.n20 163.367
R802 B.n603 B.n21 163.367
R803 B.n603 B.n26 163.367
R804 B.n27 B.n26 163.367
R805 B.n28 B.n27 163.367
R806 B.n608 B.n28 163.367
R807 B.n608 B.n33 163.367
R808 B.n34 B.n33 163.367
R809 B.n35 B.n34 163.367
R810 B.n613 B.n35 163.367
R811 B.n613 B.n40 163.367
R812 B.n41 B.n40 163.367
R813 B.n42 B.n41 163.367
R814 B.n618 B.n42 163.367
R815 B.n618 B.n47 163.367
R816 B.n48 B.n47 163.367
R817 B.n49 B.n48 163.367
R818 B.n623 B.n49 163.367
R819 B.n623 B.n54 163.367
R820 B.n55 B.n54 163.367
R821 B.n56 B.n55 163.367
R822 B.n628 B.n56 163.367
R823 B.n628 B.n61 163.367
R824 B.n62 B.n61 163.367
R825 B.n63 B.n62 163.367
R826 B.n633 B.n63 163.367
R827 B.n633 B.n68 163.367
R828 B.n69 B.n68 163.367
R829 B.n113 B.n112 163.367
R830 B.n117 B.n116 163.367
R831 B.n121 B.n120 163.367
R832 B.n125 B.n124 163.367
R833 B.n129 B.n128 163.367
R834 B.n133 B.n132 163.367
R835 B.n137 B.n136 163.367
R836 B.n141 B.n140 163.367
R837 B.n145 B.n144 163.367
R838 B.n149 B.n148 163.367
R839 B.n153 B.n152 163.367
R840 B.n157 B.n156 163.367
R841 B.n161 B.n160 163.367
R842 B.n165 B.n164 163.367
R843 B.n169 B.n168 163.367
R844 B.n173 B.n172 163.367
R845 B.n177 B.n176 163.367
R846 B.n181 B.n180 163.367
R847 B.n185 B.n184 163.367
R848 B.n189 B.n188 163.367
R849 B.n193 B.n192 163.367
R850 B.n197 B.n196 163.367
R851 B.n201 B.n200 163.367
R852 B.n205 B.n204 163.367
R853 B.n209 B.n208 163.367
R854 B.n213 B.n212 163.367
R855 B.n217 B.n216 163.367
R856 B.n221 B.n220 163.367
R857 B.n225 B.n224 163.367
R858 B.n229 B.n228 163.367
R859 B.n233 B.n232 163.367
R860 B.n235 B.n102 163.367
R861 B.n346 B.t23 100.775
R862 B.n103 B.t16 100.775
R863 B.n344 B.t13 100.766
R864 B.n106 B.t19 100.766
R865 B.n477 B.n307 99.022
R866 B.n641 B.n640 99.022
R867 B.n476 B.n475 71.676
R868 B.n470 B.n311 71.676
R869 B.n467 B.n312 71.676
R870 B.n463 B.n313 71.676
R871 B.n459 B.n314 71.676
R872 B.n455 B.n315 71.676
R873 B.n451 B.n316 71.676
R874 B.n447 B.n317 71.676
R875 B.n443 B.n318 71.676
R876 B.n439 B.n319 71.676
R877 B.n435 B.n320 71.676
R878 B.n431 B.n321 71.676
R879 B.n427 B.n322 71.676
R880 B.n423 B.n323 71.676
R881 B.n418 B.n324 71.676
R882 B.n414 B.n325 71.676
R883 B.n410 B.n326 71.676
R884 B.n406 B.n327 71.676
R885 B.n402 B.n328 71.676
R886 B.n397 B.n329 71.676
R887 B.n393 B.n330 71.676
R888 B.n389 B.n331 71.676
R889 B.n385 B.n332 71.676
R890 B.n381 B.n333 71.676
R891 B.n377 B.n334 71.676
R892 B.n373 B.n335 71.676
R893 B.n369 B.n336 71.676
R894 B.n365 B.n337 71.676
R895 B.n361 B.n338 71.676
R896 B.n357 B.n339 71.676
R897 B.n353 B.n340 71.676
R898 B.n349 B.n341 71.676
R899 B.n109 B.n70 71.676
R900 B.n113 B.n71 71.676
R901 B.n117 B.n72 71.676
R902 B.n121 B.n73 71.676
R903 B.n125 B.n74 71.676
R904 B.n129 B.n75 71.676
R905 B.n133 B.n76 71.676
R906 B.n137 B.n77 71.676
R907 B.n141 B.n78 71.676
R908 B.n145 B.n79 71.676
R909 B.n149 B.n80 71.676
R910 B.n153 B.n81 71.676
R911 B.n157 B.n82 71.676
R912 B.n161 B.n83 71.676
R913 B.n165 B.n84 71.676
R914 B.n169 B.n85 71.676
R915 B.n173 B.n86 71.676
R916 B.n177 B.n87 71.676
R917 B.n181 B.n88 71.676
R918 B.n185 B.n89 71.676
R919 B.n189 B.n90 71.676
R920 B.n193 B.n91 71.676
R921 B.n197 B.n92 71.676
R922 B.n201 B.n93 71.676
R923 B.n205 B.n94 71.676
R924 B.n209 B.n95 71.676
R925 B.n213 B.n96 71.676
R926 B.n217 B.n97 71.676
R927 B.n221 B.n98 71.676
R928 B.n225 B.n99 71.676
R929 B.n229 B.n100 71.676
R930 B.n233 B.n101 71.676
R931 B.n639 B.n102 71.676
R932 B.n639 B.n638 71.676
R933 B.n235 B.n101 71.676
R934 B.n232 B.n100 71.676
R935 B.n228 B.n99 71.676
R936 B.n224 B.n98 71.676
R937 B.n220 B.n97 71.676
R938 B.n216 B.n96 71.676
R939 B.n212 B.n95 71.676
R940 B.n208 B.n94 71.676
R941 B.n204 B.n93 71.676
R942 B.n200 B.n92 71.676
R943 B.n196 B.n91 71.676
R944 B.n192 B.n90 71.676
R945 B.n188 B.n89 71.676
R946 B.n184 B.n88 71.676
R947 B.n180 B.n87 71.676
R948 B.n176 B.n86 71.676
R949 B.n172 B.n85 71.676
R950 B.n168 B.n84 71.676
R951 B.n164 B.n83 71.676
R952 B.n160 B.n82 71.676
R953 B.n156 B.n81 71.676
R954 B.n152 B.n80 71.676
R955 B.n148 B.n79 71.676
R956 B.n144 B.n78 71.676
R957 B.n140 B.n77 71.676
R958 B.n136 B.n76 71.676
R959 B.n132 B.n75 71.676
R960 B.n128 B.n74 71.676
R961 B.n124 B.n73 71.676
R962 B.n120 B.n72 71.676
R963 B.n116 B.n71 71.676
R964 B.n112 B.n70 71.676
R965 B.n476 B.n343 71.676
R966 B.n468 B.n311 71.676
R967 B.n464 B.n312 71.676
R968 B.n460 B.n313 71.676
R969 B.n456 B.n314 71.676
R970 B.n452 B.n315 71.676
R971 B.n448 B.n316 71.676
R972 B.n444 B.n317 71.676
R973 B.n440 B.n318 71.676
R974 B.n436 B.n319 71.676
R975 B.n432 B.n320 71.676
R976 B.n428 B.n321 71.676
R977 B.n424 B.n322 71.676
R978 B.n419 B.n323 71.676
R979 B.n415 B.n324 71.676
R980 B.n411 B.n325 71.676
R981 B.n407 B.n326 71.676
R982 B.n403 B.n327 71.676
R983 B.n398 B.n328 71.676
R984 B.n394 B.n329 71.676
R985 B.n390 B.n330 71.676
R986 B.n386 B.n331 71.676
R987 B.n382 B.n332 71.676
R988 B.n378 B.n333 71.676
R989 B.n374 B.n334 71.676
R990 B.n370 B.n335 71.676
R991 B.n366 B.n336 71.676
R992 B.n362 B.n337 71.676
R993 B.n358 B.n338 71.676
R994 B.n354 B.n339 71.676
R995 B.n350 B.n340 71.676
R996 B.n341 B.n310 71.676
R997 B.n347 B.t22 69.1627
R998 B.n104 B.t17 69.1627
R999 B.n345 B.t12 69.1539
R1000 B.n107 B.t20 69.1539
R1001 B.n400 B.n347 59.5399
R1002 B.n421 B.n345 59.5399
R1003 B.n108 B.n107 59.5399
R1004 B.n105 B.n104 59.5399
R1005 B.n483 B.n307 58.5524
R1006 B.n483 B.n303 58.5524
R1007 B.n489 B.n303 58.5524
R1008 B.n489 B.n299 58.5524
R1009 B.n495 B.n299 58.5524
R1010 B.n501 B.n295 58.5524
R1011 B.n501 B.n291 58.5524
R1012 B.n507 B.n291 58.5524
R1013 B.n507 B.n287 58.5524
R1014 B.n513 B.n287 58.5524
R1015 B.n513 B.n283 58.5524
R1016 B.n519 B.n283 58.5524
R1017 B.n525 B.n279 58.5524
R1018 B.n525 B.n275 58.5524
R1019 B.n532 B.n275 58.5524
R1020 B.n532 B.n531 58.5524
R1021 B.n538 B.n268 58.5524
R1022 B.n544 B.n268 58.5524
R1023 B.n544 B.n264 58.5524
R1024 B.n550 B.n264 58.5524
R1025 B.n556 B.n260 58.5524
R1026 B.n556 B.n255 58.5524
R1027 B.n562 B.n255 58.5524
R1028 B.n562 B.n256 58.5524
R1029 B.n568 B.n248 58.5524
R1030 B.n574 B.n248 58.5524
R1031 B.n574 B.n244 58.5524
R1032 B.t8 B.n244 58.5524
R1033 B.t8 B.n240 58.5524
R1034 B.n586 B.n240 58.5524
R1035 B.n586 B.n4 58.5524
R1036 B.n713 B.n4 58.5524
R1037 B.n713 B.n712 58.5524
R1038 B.n712 B.n711 58.5524
R1039 B.n711 B.n8 58.5524
R1040 B.t6 B.n8 58.5524
R1041 B.t6 B.n705 58.5524
R1042 B.n705 B.n704 58.5524
R1043 B.n704 B.n15 58.5524
R1044 B.n698 B.n15 58.5524
R1045 B.n697 B.n696 58.5524
R1046 B.n696 B.n22 58.5524
R1047 B.n690 B.n22 58.5524
R1048 B.n690 B.n689 58.5524
R1049 B.n688 B.n29 58.5524
R1050 B.n682 B.n29 58.5524
R1051 B.n682 B.n681 58.5524
R1052 B.n681 B.n680 58.5524
R1053 B.n674 B.n39 58.5524
R1054 B.n674 B.n673 58.5524
R1055 B.n673 B.n672 58.5524
R1056 B.n672 B.n43 58.5524
R1057 B.n666 B.n665 58.5524
R1058 B.n665 B.n664 58.5524
R1059 B.n664 B.n50 58.5524
R1060 B.n658 B.n50 58.5524
R1061 B.n658 B.n657 58.5524
R1062 B.n657 B.n656 58.5524
R1063 B.n656 B.n57 58.5524
R1064 B.n650 B.n649 58.5524
R1065 B.n649 B.n648 58.5524
R1066 B.n648 B.n64 58.5524
R1067 B.n642 B.n64 58.5524
R1068 B.n642 B.n641 58.5524
R1069 B.n495 B.t11 48.2197
R1070 B.n519 B.t9 48.2197
R1071 B.n666 B.t4 48.2197
R1072 B.n650 B.t15 48.2197
R1073 B.n568 B.t3 46.4976
R1074 B.n698 B.t5 46.4976
R1075 B.n531 B.t7 36.1649
R1076 B.n39 B.t1 36.1649
R1077 B.t2 B.n260 34.4428
R1078 B.n689 B.t0 34.4428
R1079 B.n110 B.n66 32.9371
R1080 B.n637 B.n636 32.9371
R1081 B.n480 B.n479 32.9371
R1082 B.n474 B.n305 32.9371
R1083 B.n347 B.n346 31.6126
R1084 B.n345 B.n344 31.6126
R1085 B.n107 B.n106 31.6126
R1086 B.n104 B.n103 31.6126
R1087 B.n550 B.t2 24.1101
R1088 B.t0 B.n688 24.1101
R1089 B.n538 B.t7 22.388
R1090 B.n680 B.t1 22.388
R1091 B B.n715 18.0485
R1092 B.n256 B.t3 12.0553
R1093 B.t5 B.n697 12.0553
R1094 B.n111 B.n110 10.6151
R1095 B.n114 B.n111 10.6151
R1096 B.n115 B.n114 10.6151
R1097 B.n118 B.n115 10.6151
R1098 B.n119 B.n118 10.6151
R1099 B.n122 B.n119 10.6151
R1100 B.n123 B.n122 10.6151
R1101 B.n126 B.n123 10.6151
R1102 B.n127 B.n126 10.6151
R1103 B.n130 B.n127 10.6151
R1104 B.n131 B.n130 10.6151
R1105 B.n134 B.n131 10.6151
R1106 B.n135 B.n134 10.6151
R1107 B.n138 B.n135 10.6151
R1108 B.n139 B.n138 10.6151
R1109 B.n142 B.n139 10.6151
R1110 B.n143 B.n142 10.6151
R1111 B.n146 B.n143 10.6151
R1112 B.n147 B.n146 10.6151
R1113 B.n150 B.n147 10.6151
R1114 B.n151 B.n150 10.6151
R1115 B.n154 B.n151 10.6151
R1116 B.n155 B.n154 10.6151
R1117 B.n158 B.n155 10.6151
R1118 B.n159 B.n158 10.6151
R1119 B.n162 B.n159 10.6151
R1120 B.n163 B.n162 10.6151
R1121 B.n167 B.n166 10.6151
R1122 B.n170 B.n167 10.6151
R1123 B.n171 B.n170 10.6151
R1124 B.n174 B.n171 10.6151
R1125 B.n175 B.n174 10.6151
R1126 B.n178 B.n175 10.6151
R1127 B.n179 B.n178 10.6151
R1128 B.n182 B.n179 10.6151
R1129 B.n183 B.n182 10.6151
R1130 B.n187 B.n186 10.6151
R1131 B.n190 B.n187 10.6151
R1132 B.n191 B.n190 10.6151
R1133 B.n194 B.n191 10.6151
R1134 B.n195 B.n194 10.6151
R1135 B.n198 B.n195 10.6151
R1136 B.n199 B.n198 10.6151
R1137 B.n202 B.n199 10.6151
R1138 B.n203 B.n202 10.6151
R1139 B.n206 B.n203 10.6151
R1140 B.n207 B.n206 10.6151
R1141 B.n210 B.n207 10.6151
R1142 B.n211 B.n210 10.6151
R1143 B.n214 B.n211 10.6151
R1144 B.n215 B.n214 10.6151
R1145 B.n218 B.n215 10.6151
R1146 B.n219 B.n218 10.6151
R1147 B.n222 B.n219 10.6151
R1148 B.n223 B.n222 10.6151
R1149 B.n226 B.n223 10.6151
R1150 B.n227 B.n226 10.6151
R1151 B.n230 B.n227 10.6151
R1152 B.n231 B.n230 10.6151
R1153 B.n234 B.n231 10.6151
R1154 B.n236 B.n234 10.6151
R1155 B.n237 B.n236 10.6151
R1156 B.n637 B.n237 10.6151
R1157 B.n481 B.n480 10.6151
R1158 B.n481 B.n301 10.6151
R1159 B.n491 B.n301 10.6151
R1160 B.n492 B.n491 10.6151
R1161 B.n493 B.n492 10.6151
R1162 B.n493 B.n293 10.6151
R1163 B.n503 B.n293 10.6151
R1164 B.n504 B.n503 10.6151
R1165 B.n505 B.n504 10.6151
R1166 B.n505 B.n285 10.6151
R1167 B.n515 B.n285 10.6151
R1168 B.n516 B.n515 10.6151
R1169 B.n517 B.n516 10.6151
R1170 B.n517 B.n277 10.6151
R1171 B.n527 B.n277 10.6151
R1172 B.n528 B.n527 10.6151
R1173 B.n529 B.n528 10.6151
R1174 B.n529 B.n270 10.6151
R1175 B.n540 B.n270 10.6151
R1176 B.n541 B.n540 10.6151
R1177 B.n542 B.n541 10.6151
R1178 B.n542 B.n262 10.6151
R1179 B.n552 B.n262 10.6151
R1180 B.n553 B.n552 10.6151
R1181 B.n554 B.n553 10.6151
R1182 B.n554 B.n253 10.6151
R1183 B.n564 B.n253 10.6151
R1184 B.n565 B.n564 10.6151
R1185 B.n566 B.n565 10.6151
R1186 B.n566 B.n246 10.6151
R1187 B.n576 B.n246 10.6151
R1188 B.n577 B.n576 10.6151
R1189 B.n579 B.n577 10.6151
R1190 B.n579 B.n578 10.6151
R1191 B.n578 B.n238 10.6151
R1192 B.n589 B.n238 10.6151
R1193 B.n590 B.n589 10.6151
R1194 B.n591 B.n590 10.6151
R1195 B.n592 B.n591 10.6151
R1196 B.n594 B.n592 10.6151
R1197 B.n595 B.n594 10.6151
R1198 B.n596 B.n595 10.6151
R1199 B.n597 B.n596 10.6151
R1200 B.n599 B.n597 10.6151
R1201 B.n600 B.n599 10.6151
R1202 B.n601 B.n600 10.6151
R1203 B.n602 B.n601 10.6151
R1204 B.n604 B.n602 10.6151
R1205 B.n605 B.n604 10.6151
R1206 B.n606 B.n605 10.6151
R1207 B.n607 B.n606 10.6151
R1208 B.n609 B.n607 10.6151
R1209 B.n610 B.n609 10.6151
R1210 B.n611 B.n610 10.6151
R1211 B.n612 B.n611 10.6151
R1212 B.n614 B.n612 10.6151
R1213 B.n615 B.n614 10.6151
R1214 B.n616 B.n615 10.6151
R1215 B.n617 B.n616 10.6151
R1216 B.n619 B.n617 10.6151
R1217 B.n620 B.n619 10.6151
R1218 B.n621 B.n620 10.6151
R1219 B.n622 B.n621 10.6151
R1220 B.n624 B.n622 10.6151
R1221 B.n625 B.n624 10.6151
R1222 B.n626 B.n625 10.6151
R1223 B.n627 B.n626 10.6151
R1224 B.n629 B.n627 10.6151
R1225 B.n630 B.n629 10.6151
R1226 B.n631 B.n630 10.6151
R1227 B.n632 B.n631 10.6151
R1228 B.n634 B.n632 10.6151
R1229 B.n635 B.n634 10.6151
R1230 B.n636 B.n635 10.6151
R1231 B.n474 B.n473 10.6151
R1232 B.n473 B.n472 10.6151
R1233 B.n472 B.n471 10.6151
R1234 B.n471 B.n469 10.6151
R1235 B.n469 B.n466 10.6151
R1236 B.n466 B.n465 10.6151
R1237 B.n465 B.n462 10.6151
R1238 B.n462 B.n461 10.6151
R1239 B.n461 B.n458 10.6151
R1240 B.n458 B.n457 10.6151
R1241 B.n457 B.n454 10.6151
R1242 B.n454 B.n453 10.6151
R1243 B.n453 B.n450 10.6151
R1244 B.n450 B.n449 10.6151
R1245 B.n449 B.n446 10.6151
R1246 B.n446 B.n445 10.6151
R1247 B.n445 B.n442 10.6151
R1248 B.n442 B.n441 10.6151
R1249 B.n441 B.n438 10.6151
R1250 B.n438 B.n437 10.6151
R1251 B.n437 B.n434 10.6151
R1252 B.n434 B.n433 10.6151
R1253 B.n433 B.n430 10.6151
R1254 B.n430 B.n429 10.6151
R1255 B.n429 B.n426 10.6151
R1256 B.n426 B.n425 10.6151
R1257 B.n425 B.n422 10.6151
R1258 B.n420 B.n417 10.6151
R1259 B.n417 B.n416 10.6151
R1260 B.n416 B.n413 10.6151
R1261 B.n413 B.n412 10.6151
R1262 B.n412 B.n409 10.6151
R1263 B.n409 B.n408 10.6151
R1264 B.n408 B.n405 10.6151
R1265 B.n405 B.n404 10.6151
R1266 B.n404 B.n401 10.6151
R1267 B.n399 B.n396 10.6151
R1268 B.n396 B.n395 10.6151
R1269 B.n395 B.n392 10.6151
R1270 B.n392 B.n391 10.6151
R1271 B.n391 B.n388 10.6151
R1272 B.n388 B.n387 10.6151
R1273 B.n387 B.n384 10.6151
R1274 B.n384 B.n383 10.6151
R1275 B.n383 B.n380 10.6151
R1276 B.n380 B.n379 10.6151
R1277 B.n379 B.n376 10.6151
R1278 B.n376 B.n375 10.6151
R1279 B.n375 B.n372 10.6151
R1280 B.n372 B.n371 10.6151
R1281 B.n371 B.n368 10.6151
R1282 B.n368 B.n367 10.6151
R1283 B.n367 B.n364 10.6151
R1284 B.n364 B.n363 10.6151
R1285 B.n363 B.n360 10.6151
R1286 B.n360 B.n359 10.6151
R1287 B.n359 B.n356 10.6151
R1288 B.n356 B.n355 10.6151
R1289 B.n355 B.n352 10.6151
R1290 B.n352 B.n351 10.6151
R1291 B.n351 B.n348 10.6151
R1292 B.n348 B.n309 10.6151
R1293 B.n479 B.n309 10.6151
R1294 B.n485 B.n305 10.6151
R1295 B.n486 B.n485 10.6151
R1296 B.n487 B.n486 10.6151
R1297 B.n487 B.n297 10.6151
R1298 B.n497 B.n297 10.6151
R1299 B.n498 B.n497 10.6151
R1300 B.n499 B.n498 10.6151
R1301 B.n499 B.n289 10.6151
R1302 B.n509 B.n289 10.6151
R1303 B.n510 B.n509 10.6151
R1304 B.n511 B.n510 10.6151
R1305 B.n511 B.n281 10.6151
R1306 B.n521 B.n281 10.6151
R1307 B.n522 B.n521 10.6151
R1308 B.n523 B.n522 10.6151
R1309 B.n523 B.n273 10.6151
R1310 B.n534 B.n273 10.6151
R1311 B.n535 B.n534 10.6151
R1312 B.n536 B.n535 10.6151
R1313 B.n536 B.n266 10.6151
R1314 B.n546 B.n266 10.6151
R1315 B.n547 B.n546 10.6151
R1316 B.n548 B.n547 10.6151
R1317 B.n548 B.n258 10.6151
R1318 B.n558 B.n258 10.6151
R1319 B.n559 B.n558 10.6151
R1320 B.n560 B.n559 10.6151
R1321 B.n560 B.n250 10.6151
R1322 B.n570 B.n250 10.6151
R1323 B.n571 B.n570 10.6151
R1324 B.n572 B.n571 10.6151
R1325 B.n572 B.n242 10.6151
R1326 B.n582 B.n242 10.6151
R1327 B.n583 B.n582 10.6151
R1328 B.n584 B.n583 10.6151
R1329 B.n584 B.n0 10.6151
R1330 B.n709 B.n1 10.6151
R1331 B.n709 B.n708 10.6151
R1332 B.n708 B.n707 10.6151
R1333 B.n707 B.n10 10.6151
R1334 B.n702 B.n10 10.6151
R1335 B.n702 B.n701 10.6151
R1336 B.n701 B.n700 10.6151
R1337 B.n700 B.n17 10.6151
R1338 B.n694 B.n17 10.6151
R1339 B.n694 B.n693 10.6151
R1340 B.n693 B.n692 10.6151
R1341 B.n692 B.n24 10.6151
R1342 B.n686 B.n24 10.6151
R1343 B.n686 B.n685 10.6151
R1344 B.n685 B.n684 10.6151
R1345 B.n684 B.n31 10.6151
R1346 B.n678 B.n31 10.6151
R1347 B.n678 B.n677 10.6151
R1348 B.n677 B.n676 10.6151
R1349 B.n676 B.n37 10.6151
R1350 B.n670 B.n37 10.6151
R1351 B.n670 B.n669 10.6151
R1352 B.n669 B.n668 10.6151
R1353 B.n668 B.n45 10.6151
R1354 B.n662 B.n45 10.6151
R1355 B.n662 B.n661 10.6151
R1356 B.n661 B.n660 10.6151
R1357 B.n660 B.n52 10.6151
R1358 B.n654 B.n52 10.6151
R1359 B.n654 B.n653 10.6151
R1360 B.n653 B.n652 10.6151
R1361 B.n652 B.n59 10.6151
R1362 B.n646 B.n59 10.6151
R1363 B.n646 B.n645 10.6151
R1364 B.n645 B.n644 10.6151
R1365 B.n644 B.n66 10.6151
R1366 B.t11 B.n295 10.3332
R1367 B.t9 B.n279 10.3332
R1368 B.t4 B.n43 10.3332
R1369 B.t15 B.n57 10.3332
R1370 B.n163 B.n108 9.36635
R1371 B.n186 B.n105 9.36635
R1372 B.n422 B.n421 9.36635
R1373 B.n400 B.n399 9.36635
R1374 B.n715 B.n0 2.81026
R1375 B.n715 B.n1 2.81026
R1376 B.n166 B.n108 1.24928
R1377 B.n183 B.n105 1.24928
R1378 B.n421 B.n420 1.24928
R1379 B.n401 B.n400 1.24928
R1380 VP.n33 VP.n7 173.105
R1381 VP.n56 VP.n55 173.105
R1382 VP.n32 VP.n31 173.105
R1383 VP.n14 VP.t8 168.714
R1384 VP.n16 VP.n15 161.3
R1385 VP.n17 VP.n12 161.3
R1386 VP.n19 VP.n18 161.3
R1387 VP.n20 VP.n11 161.3
R1388 VP.n22 VP.n21 161.3
R1389 VP.n23 VP.n10 161.3
R1390 VP.n26 VP.n25 161.3
R1391 VP.n27 VP.n9 161.3
R1392 VP.n29 VP.n28 161.3
R1393 VP.n30 VP.n8 161.3
R1394 VP.n54 VP.n0 161.3
R1395 VP.n53 VP.n52 161.3
R1396 VP.n51 VP.n1 161.3
R1397 VP.n50 VP.n49 161.3
R1398 VP.n47 VP.n2 161.3
R1399 VP.n46 VP.n45 161.3
R1400 VP.n44 VP.n3 161.3
R1401 VP.n43 VP.n42 161.3
R1402 VP.n41 VP.n4 161.3
R1403 VP.n40 VP.n39 161.3
R1404 VP.n38 VP.n37 161.3
R1405 VP.n36 VP.n6 161.3
R1406 VP.n35 VP.n34 161.3
R1407 VP.n3 VP.t2 139.038
R1408 VP.n7 VP.t0 139.038
R1409 VP.n5 VP.t7 139.038
R1410 VP.n48 VP.t1 139.038
R1411 VP.n55 VP.t6 139.038
R1412 VP.n11 VP.t9 139.038
R1413 VP.n31 VP.t4 139.038
R1414 VP.n24 VP.t5 139.038
R1415 VP.n13 VP.t3 139.038
R1416 VP.n14 VP.n13 58.6212
R1417 VP.n42 VP.n41 56.5617
R1418 VP.n47 VP.n46 56.5617
R1419 VP.n23 VP.n22 56.5617
R1420 VP.n18 VP.n17 56.5617
R1421 VP.n37 VP.n36 45.9053
R1422 VP.n53 VP.n1 45.9053
R1423 VP.n29 VP.n9 45.9053
R1424 VP.n33 VP.n32 42.5573
R1425 VP.n36 VP.n35 35.2488
R1426 VP.n54 VP.n53 35.2488
R1427 VP.n30 VP.n29 35.2488
R1428 VP.n15 VP.n14 27.0756
R1429 VP.n41 VP.n40 24.5923
R1430 VP.n42 VP.n3 24.5923
R1431 VP.n46 VP.n3 24.5923
R1432 VP.n49 VP.n47 24.5923
R1433 VP.n25 VP.n23 24.5923
R1434 VP.n18 VP.n11 24.5923
R1435 VP.n22 VP.n11 24.5923
R1436 VP.n17 VP.n16 24.5923
R1437 VP.n37 VP.n5 18.1985
R1438 VP.n48 VP.n1 18.1985
R1439 VP.n24 VP.n9 18.1985
R1440 VP.n35 VP.n7 12.7883
R1441 VP.n55 VP.n54 12.7883
R1442 VP.n31 VP.n30 12.7883
R1443 VP.n40 VP.n5 6.39438
R1444 VP.n49 VP.n48 6.39438
R1445 VP.n25 VP.n24 6.39438
R1446 VP.n16 VP.n13 6.39438
R1447 VP.n15 VP.n12 0.189894
R1448 VP.n19 VP.n12 0.189894
R1449 VP.n20 VP.n19 0.189894
R1450 VP.n21 VP.n20 0.189894
R1451 VP.n21 VP.n10 0.189894
R1452 VP.n26 VP.n10 0.189894
R1453 VP.n27 VP.n26 0.189894
R1454 VP.n28 VP.n27 0.189894
R1455 VP.n28 VP.n8 0.189894
R1456 VP.n32 VP.n8 0.189894
R1457 VP.n34 VP.n33 0.189894
R1458 VP.n34 VP.n6 0.189894
R1459 VP.n38 VP.n6 0.189894
R1460 VP.n39 VP.n38 0.189894
R1461 VP.n39 VP.n4 0.189894
R1462 VP.n43 VP.n4 0.189894
R1463 VP.n44 VP.n43 0.189894
R1464 VP.n45 VP.n44 0.189894
R1465 VP.n45 VP.n2 0.189894
R1466 VP.n50 VP.n2 0.189894
R1467 VP.n51 VP.n50 0.189894
R1468 VP.n52 VP.n51 0.189894
R1469 VP.n52 VP.n0 0.189894
R1470 VP.n56 VP.n0 0.189894
R1471 VP VP.n56 0.0516364
R1472 VDD1.n1 VDD1.t1 69.5001
R1473 VDD1.n3 VDD1.t9 69.4999
R1474 VDD1.n5 VDD1.n4 66.4533
R1475 VDD1.n1 VDD1.n0 65.4549
R1476 VDD1.n7 VDD1.n6 65.4547
R1477 VDD1.n3 VDD1.n2 65.4547
R1478 VDD1.n7 VDD1.n5 38.141
R1479 VDD1.n6 VDD1.t4 2.6405
R1480 VDD1.n6 VDD1.t5 2.6405
R1481 VDD1.n0 VDD1.t6 2.6405
R1482 VDD1.n0 VDD1.t0 2.6405
R1483 VDD1.n4 VDD1.t8 2.6405
R1484 VDD1.n4 VDD1.t3 2.6405
R1485 VDD1.n2 VDD1.t2 2.6405
R1486 VDD1.n2 VDD1.t7 2.6405
R1487 VDD1 VDD1.n7 0.99619
R1488 VDD1 VDD1.n1 0.409983
R1489 VDD1.n5 VDD1.n3 0.296447
C0 VDD2 VDD1 1.34282f
C1 VDD2 VP 0.417623f
C2 VTAIL VN 5.96492f
C3 VN VDD1 0.150655f
C4 VN VP 5.64514f
C5 VDD2 VN 5.68448f
C6 VTAIL VDD1 8.290831f
C7 VTAIL VP 5.97924f
C8 VP VDD1 5.94848f
C9 VDD2 VTAIL 8.33274f
C10 VDD2 B 4.868491f
C11 VDD1 B 4.835181f
C12 VTAIL B 5.418381f
C13 VN B 11.648231f
C14 VP B 10.082085f
C15 VDD1.t1 B 1.50152f
C16 VDD1.t6 B 0.136644f
C17 VDD1.t0 B 0.136644f
C18 VDD1.n0 B 1.17653f
C19 VDD1.n1 B 0.66082f
C20 VDD1.t9 B 1.50152f
C21 VDD1.t2 B 0.136644f
C22 VDD1.t7 B 0.136644f
C23 VDD1.n2 B 1.17653f
C24 VDD1.n3 B 0.654195f
C25 VDD1.t8 B 0.136644f
C26 VDD1.t3 B 0.136644f
C27 VDD1.n4 B 1.1821f
C28 VDD1.n5 B 1.87413f
C29 VDD1.t4 B 0.136644f
C30 VDD1.t5 B 0.136644f
C31 VDD1.n6 B 1.17653f
C32 VDD1.n7 B 2.09859f
C33 VP.n0 B 0.033826f
C34 VP.t6 B 0.883176f
C35 VP.n1 B 0.056401f
C36 VP.n2 B 0.033826f
C37 VP.t2 B 0.883176f
C38 VP.n3 B 0.370811f
C39 VP.n4 B 0.033826f
C40 VP.t7 B 0.883176f
C41 VP.n5 B 0.339051f
C42 VP.n6 B 0.033826f
C43 VP.t0 B 0.883176f
C44 VP.n7 B 0.400963f
C45 VP.n8 B 0.033826f
C46 VP.t4 B 0.883176f
C47 VP.n9 B 0.056401f
C48 VP.n10 B 0.033826f
C49 VP.t9 B 0.883176f
C50 VP.n11 B 0.370811f
C51 VP.n12 B 0.033826f
C52 VP.t3 B 0.883176f
C53 VP.n13 B 0.38641f
C54 VP.t8 B 0.96169f
C55 VP.n14 B 0.414958f
C56 VP.n15 B 0.178617f
C57 VP.n16 B 0.039811f
C58 VP.n17 B 0.043088f
C59 VP.n18 B 0.055254f
C60 VP.n19 B 0.033826f
C61 VP.n20 B 0.033826f
C62 VP.n21 B 0.033826f
C63 VP.n22 B 0.055254f
C64 VP.n23 B 0.043088f
C65 VP.t5 B 0.883176f
C66 VP.n24 B 0.339051f
C67 VP.n25 B 0.039811f
C68 VP.n26 B 0.033826f
C69 VP.n27 B 0.033826f
C70 VP.n28 B 0.033826f
C71 VP.n29 B 0.028647f
C72 VP.n30 B 0.053105f
C73 VP.n31 B 0.400963f
C74 VP.n32 B 1.43158f
C75 VP.n33 B 1.46023f
C76 VP.n34 B 0.033826f
C77 VP.n35 B 0.053105f
C78 VP.n36 B 0.028647f
C79 VP.n37 B 0.056401f
C80 VP.n38 B 0.033826f
C81 VP.n39 B 0.033826f
C82 VP.n40 B 0.039811f
C83 VP.n41 B 0.043088f
C84 VP.n42 B 0.055254f
C85 VP.n43 B 0.033826f
C86 VP.n44 B 0.033826f
C87 VP.n45 B 0.033826f
C88 VP.n46 B 0.055254f
C89 VP.n47 B 0.043088f
C90 VP.t1 B 0.883176f
C91 VP.n48 B 0.339051f
C92 VP.n49 B 0.039811f
C93 VP.n50 B 0.033826f
C94 VP.n51 B 0.033826f
C95 VP.n52 B 0.033826f
C96 VP.n53 B 0.028647f
C97 VP.n54 B 0.053105f
C98 VP.n55 B 0.400963f
C99 VP.n56 B 0.030744f
C100 VTAIL.t14 B 0.153701f
C101 VTAIL.t19 B 0.153701f
C102 VTAIL.n0 B 1.25494f
C103 VTAIL.n1 B 0.429184f
C104 VTAIL.t8 B 1.59605f
C105 VTAIL.n2 B 0.531745f
C106 VTAIL.t2 B 0.153701f
C107 VTAIL.t3 B 0.153701f
C108 VTAIL.n3 B 1.25494f
C109 VTAIL.n4 B 0.473127f
C110 VTAIL.t9 B 0.153701f
C111 VTAIL.t7 B 0.153701f
C112 VTAIL.n5 B 1.25494f
C113 VTAIL.n6 B 1.4831f
C114 VTAIL.t15 B 0.153701f
C115 VTAIL.t11 B 0.153701f
C116 VTAIL.n7 B 1.25494f
C117 VTAIL.n8 B 1.4831f
C118 VTAIL.t10 B 0.153701f
C119 VTAIL.t16 B 0.153701f
C120 VTAIL.n9 B 1.25494f
C121 VTAIL.n10 B 0.473123f
C122 VTAIL.t13 B 1.59606f
C123 VTAIL.n11 B 0.531741f
C124 VTAIL.t6 B 0.153701f
C125 VTAIL.t5 B 0.153701f
C126 VTAIL.n12 B 1.25494f
C127 VTAIL.n13 B 0.453673f
C128 VTAIL.t0 B 0.153701f
C129 VTAIL.t1 B 0.153701f
C130 VTAIL.n14 B 1.25494f
C131 VTAIL.n15 B 0.473123f
C132 VTAIL.t4 B 1.59605f
C133 VTAIL.n16 B 1.44375f
C134 VTAIL.t18 B 1.59605f
C135 VTAIL.n17 B 1.44375f
C136 VTAIL.t17 B 0.153701f
C137 VTAIL.t12 B 0.153701f
C138 VTAIL.n18 B 1.25494f
C139 VTAIL.n19 B 0.380198f
C140 VDD2.t6 B 1.4893f
C141 VDD2.t4 B 0.135533f
C142 VDD2.t1 B 0.135533f
C143 VDD2.n0 B 1.16695f
C144 VDD2.n1 B 0.648873f
C145 VDD2.t9 B 0.135533f
C146 VDD2.t7 B 0.135533f
C147 VDD2.n2 B 1.17248f
C148 VDD2.n3 B 1.77747f
C149 VDD2.t0 B 1.48227f
C150 VDD2.n4 B 2.05941f
C151 VDD2.t8 B 0.135533f
C152 VDD2.t2 B 0.135533f
C153 VDD2.n5 B 1.16696f
C154 VDD2.n6 B 0.314561f
C155 VDD2.t3 B 0.135533f
C156 VDD2.t5 B 0.135533f
C157 VDD2.n7 B 1.17245f
C158 VN.n0 B 0.033348f
C159 VN.t1 B 0.870717f
C160 VN.n1 B 0.055605f
C161 VN.n2 B 0.033348f
C162 VN.t2 B 0.870717f
C163 VN.n3 B 0.36558f
C164 VN.n4 B 0.033348f
C165 VN.t0 B 0.870717f
C166 VN.n5 B 0.380959f
C167 VN.t5 B 0.948123f
C168 VN.n6 B 0.409104f
C169 VN.n7 B 0.176097f
C170 VN.n8 B 0.03925f
C171 VN.n9 B 0.04248f
C172 VN.n10 B 0.054474f
C173 VN.n11 B 0.033348f
C174 VN.n12 B 0.033348f
C175 VN.n13 B 0.033348f
C176 VN.n14 B 0.054474f
C177 VN.n15 B 0.04248f
C178 VN.t7 B 0.870717f
C179 VN.n16 B 0.334268f
C180 VN.n17 B 0.03925f
C181 VN.n18 B 0.033348f
C182 VN.n19 B 0.033348f
C183 VN.n20 B 0.033348f
C184 VN.n21 B 0.028243f
C185 VN.n22 B 0.052356f
C186 VN.n23 B 0.395306f
C187 VN.n24 B 0.030311f
C188 VN.n25 B 0.033348f
C189 VN.t4 B 0.870717f
C190 VN.n26 B 0.055605f
C191 VN.n27 B 0.033348f
C192 VN.t8 B 0.870717f
C193 VN.n28 B 0.334268f
C194 VN.t9 B 0.870717f
C195 VN.n29 B 0.36558f
C196 VN.n30 B 0.033348f
C197 VN.t3 B 0.870717f
C198 VN.n31 B 0.380959f
C199 VN.t6 B 0.948123f
C200 VN.n32 B 0.409104f
C201 VN.n33 B 0.176097f
C202 VN.n34 B 0.03925f
C203 VN.n35 B 0.04248f
C204 VN.n36 B 0.054474f
C205 VN.n37 B 0.033348f
C206 VN.n38 B 0.033348f
C207 VN.n39 B 0.033348f
C208 VN.n40 B 0.054474f
C209 VN.n41 B 0.04248f
C210 VN.n42 B 0.03925f
C211 VN.n43 B 0.033348f
C212 VN.n44 B 0.033348f
C213 VN.n45 B 0.033348f
C214 VN.n46 B 0.028243f
C215 VN.n47 B 0.052356f
C216 VN.n48 B 0.395306f
C217 VN.n49 B 1.43326f
.ends

