* NGSPICE file created from diff_pair_sample_0207.ext - technology: sky130A

.subckt diff_pair_sample_0207 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=2.0196 ps=12.57 w=12.24 l=1.52
X1 B.t11 B.t9 B.t10 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=0 ps=0 w=12.24 l=1.52
X2 VDD2.t1 VN.t1 VTAIL.t10 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=2.0196 ps=12.57 w=12.24 l=1.52
X3 VDD1.t5 VP.t0 VTAIL.t5 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=2.0196 ps=12.57 w=12.24 l=1.52
X4 VDD1.t4 VP.t1 VTAIL.t4 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=4.7736 ps=25.26 w=12.24 l=1.52
X5 VDD2.t3 VN.t2 VTAIL.t9 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=2.0196 ps=12.57 w=12.24 l=1.52
X6 VTAIL.t8 VN.t3 VDD2.t5 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=2.0196 ps=12.57 w=12.24 l=1.52
X7 VDD2.t2 VN.t4 VTAIL.t7 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=4.7736 ps=25.26 w=12.24 l=1.52
X8 VDD2.t4 VN.t5 VTAIL.t6 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=4.7736 ps=25.26 w=12.24 l=1.52
X9 B.t8 B.t6 B.t7 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=0 ps=0 w=12.24 l=1.52
X10 VTAIL.t3 VP.t2 VDD1.t3 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=2.0196 ps=12.57 w=12.24 l=1.52
X11 VDD1.t2 VP.t3 VTAIL.t0 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=2.0196 ps=12.57 w=12.24 l=1.52
X12 VTAIL.t2 VP.t4 VDD1.t1 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=2.0196 ps=12.57 w=12.24 l=1.52
X13 B.t5 B.t3 B.t4 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=0 ps=0 w=12.24 l=1.52
X14 B.t2 B.t0 B.t1 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=4.7736 pd=25.26 as=0 ps=0 w=12.24 l=1.52
X15 VDD1.t0 VP.t5 VTAIL.t1 w_n2450_n3416# sky130_fd_pr__pfet_01v8 ad=2.0196 pd=12.57 as=4.7736 ps=25.26 w=12.24 l=1.52
R0 VN.n2 VN.t1 224.964
R1 VN.n14 VN.t4 224.964
R2 VN.n3 VN.t3 194.069
R3 VN.n10 VN.t5 194.069
R4 VN.n15 VN.t0 194.069
R5 VN.n22 VN.t2 194.069
R6 VN.n11 VN.n10 180.775
R7 VN.n23 VN.n22 180.775
R8 VN.n21 VN.n12 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n13 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n9 VN.n0 161.3
R13 VN.n8 VN.n7 161.3
R14 VN.n6 VN.n1 161.3
R15 VN.n5 VN.n4 161.3
R16 VN.n8 VN.n1 56.4773
R17 VN.n20 VN.n13 56.4773
R18 VN.n3 VN.n2 53.4877
R19 VN.n15 VN.n14 53.4877
R20 VN VN.n23 44.8547
R21 VN.n4 VN.n1 24.3439
R22 VN.n9 VN.n8 24.3439
R23 VN.n16 VN.n13 24.3439
R24 VN.n21 VN.n20 24.3439
R25 VN.n17 VN.n14 18.3124
R26 VN.n5 VN.n2 18.3124
R27 VN.n4 VN.n3 12.1722
R28 VN.n16 VN.n15 12.1722
R29 VN.n10 VN.n9 4.86919
R30 VN.n22 VN.n21 4.86919
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VDD2.n1 VDD2.t1 79.146
R41 VDD2.n2 VDD2.t3 78.0063
R42 VDD2.n1 VDD2.n0 75.6938
R43 VDD2 VDD2.n3 75.69
R44 VDD2.n2 VDD2.n1 39.4502
R45 VDD2.n3 VDD2.t0 2.65614
R46 VDD2.n3 VDD2.t2 2.65614
R47 VDD2.n0 VDD2.t5 2.65614
R48 VDD2.n0 VDD2.t4 2.65614
R49 VDD2 VDD2.n2 1.25481
R50 VTAIL.n7 VTAIL.t7 61.3275
R51 VTAIL.n11 VTAIL.t6 61.3265
R52 VTAIL.n2 VTAIL.t4 61.3265
R53 VTAIL.n10 VTAIL.t1 61.3263
R54 VTAIL.n9 VTAIL.n8 58.6719
R55 VTAIL.n6 VTAIL.n5 58.6719
R56 VTAIL.n1 VTAIL.n0 58.6717
R57 VTAIL.n4 VTAIL.n3 58.6717
R58 VTAIL.n6 VTAIL.n4 26.1083
R59 VTAIL.n11 VTAIL.n10 24.5134
R60 VTAIL.n0 VTAIL.t10 2.65614
R61 VTAIL.n0 VTAIL.t8 2.65614
R62 VTAIL.n3 VTAIL.t0 2.65614
R63 VTAIL.n3 VTAIL.t3 2.65614
R64 VTAIL.n8 VTAIL.t5 2.65614
R65 VTAIL.n8 VTAIL.t2 2.65614
R66 VTAIL.n5 VTAIL.t9 2.65614
R67 VTAIL.n5 VTAIL.t11 2.65614
R68 VTAIL.n7 VTAIL.n6 1.59533
R69 VTAIL.n10 VTAIL.n9 1.59533
R70 VTAIL.n4 VTAIL.n2 1.59533
R71 VTAIL.n9 VTAIL.n7 1.26774
R72 VTAIL.n2 VTAIL.n1 1.26774
R73 VTAIL VTAIL.n11 1.13843
R74 VTAIL VTAIL.n1 0.457397
R75 B.n443 B.n68 585
R76 B.n445 B.n444 585
R77 B.n446 B.n67 585
R78 B.n448 B.n447 585
R79 B.n449 B.n66 585
R80 B.n451 B.n450 585
R81 B.n452 B.n65 585
R82 B.n454 B.n453 585
R83 B.n455 B.n64 585
R84 B.n457 B.n456 585
R85 B.n458 B.n63 585
R86 B.n460 B.n459 585
R87 B.n461 B.n62 585
R88 B.n463 B.n462 585
R89 B.n464 B.n61 585
R90 B.n466 B.n465 585
R91 B.n467 B.n60 585
R92 B.n469 B.n468 585
R93 B.n470 B.n59 585
R94 B.n472 B.n471 585
R95 B.n473 B.n58 585
R96 B.n475 B.n474 585
R97 B.n476 B.n57 585
R98 B.n478 B.n477 585
R99 B.n479 B.n56 585
R100 B.n481 B.n480 585
R101 B.n482 B.n55 585
R102 B.n484 B.n483 585
R103 B.n485 B.n54 585
R104 B.n487 B.n486 585
R105 B.n488 B.n53 585
R106 B.n490 B.n489 585
R107 B.n491 B.n52 585
R108 B.n493 B.n492 585
R109 B.n494 B.n51 585
R110 B.n496 B.n495 585
R111 B.n497 B.n50 585
R112 B.n499 B.n498 585
R113 B.n500 B.n49 585
R114 B.n502 B.n501 585
R115 B.n503 B.n48 585
R116 B.n505 B.n504 585
R117 B.n507 B.n45 585
R118 B.n509 B.n508 585
R119 B.n510 B.n44 585
R120 B.n512 B.n511 585
R121 B.n513 B.n43 585
R122 B.n515 B.n514 585
R123 B.n516 B.n42 585
R124 B.n518 B.n517 585
R125 B.n519 B.n41 585
R126 B.n521 B.n520 585
R127 B.n523 B.n522 585
R128 B.n524 B.n37 585
R129 B.n526 B.n525 585
R130 B.n527 B.n36 585
R131 B.n529 B.n528 585
R132 B.n530 B.n35 585
R133 B.n532 B.n531 585
R134 B.n533 B.n34 585
R135 B.n535 B.n534 585
R136 B.n536 B.n33 585
R137 B.n538 B.n537 585
R138 B.n539 B.n32 585
R139 B.n541 B.n540 585
R140 B.n542 B.n31 585
R141 B.n544 B.n543 585
R142 B.n545 B.n30 585
R143 B.n547 B.n546 585
R144 B.n548 B.n29 585
R145 B.n550 B.n549 585
R146 B.n551 B.n28 585
R147 B.n553 B.n552 585
R148 B.n554 B.n27 585
R149 B.n556 B.n555 585
R150 B.n557 B.n26 585
R151 B.n559 B.n558 585
R152 B.n560 B.n25 585
R153 B.n562 B.n561 585
R154 B.n563 B.n24 585
R155 B.n565 B.n564 585
R156 B.n566 B.n23 585
R157 B.n568 B.n567 585
R158 B.n569 B.n22 585
R159 B.n571 B.n570 585
R160 B.n572 B.n21 585
R161 B.n574 B.n573 585
R162 B.n575 B.n20 585
R163 B.n577 B.n576 585
R164 B.n578 B.n19 585
R165 B.n580 B.n579 585
R166 B.n581 B.n18 585
R167 B.n583 B.n582 585
R168 B.n584 B.n17 585
R169 B.n442 B.n441 585
R170 B.n440 B.n69 585
R171 B.n439 B.n438 585
R172 B.n437 B.n70 585
R173 B.n436 B.n435 585
R174 B.n434 B.n71 585
R175 B.n433 B.n432 585
R176 B.n431 B.n72 585
R177 B.n430 B.n429 585
R178 B.n428 B.n73 585
R179 B.n427 B.n426 585
R180 B.n425 B.n74 585
R181 B.n424 B.n423 585
R182 B.n422 B.n75 585
R183 B.n421 B.n420 585
R184 B.n419 B.n76 585
R185 B.n418 B.n417 585
R186 B.n416 B.n77 585
R187 B.n415 B.n414 585
R188 B.n413 B.n78 585
R189 B.n412 B.n411 585
R190 B.n410 B.n79 585
R191 B.n409 B.n408 585
R192 B.n407 B.n80 585
R193 B.n406 B.n405 585
R194 B.n404 B.n81 585
R195 B.n403 B.n402 585
R196 B.n401 B.n82 585
R197 B.n400 B.n399 585
R198 B.n398 B.n83 585
R199 B.n397 B.n396 585
R200 B.n395 B.n84 585
R201 B.n394 B.n393 585
R202 B.n392 B.n85 585
R203 B.n391 B.n390 585
R204 B.n389 B.n86 585
R205 B.n388 B.n387 585
R206 B.n386 B.n87 585
R207 B.n385 B.n384 585
R208 B.n383 B.n88 585
R209 B.n382 B.n381 585
R210 B.n380 B.n89 585
R211 B.n379 B.n378 585
R212 B.n377 B.n90 585
R213 B.n376 B.n375 585
R214 B.n374 B.n91 585
R215 B.n373 B.n372 585
R216 B.n371 B.n92 585
R217 B.n370 B.n369 585
R218 B.n368 B.n93 585
R219 B.n367 B.n366 585
R220 B.n365 B.n94 585
R221 B.n364 B.n363 585
R222 B.n362 B.n95 585
R223 B.n361 B.n360 585
R224 B.n359 B.n96 585
R225 B.n358 B.n357 585
R226 B.n356 B.n97 585
R227 B.n355 B.n354 585
R228 B.n353 B.n98 585
R229 B.n352 B.n351 585
R230 B.n209 B.n150 585
R231 B.n211 B.n210 585
R232 B.n212 B.n149 585
R233 B.n214 B.n213 585
R234 B.n215 B.n148 585
R235 B.n217 B.n216 585
R236 B.n218 B.n147 585
R237 B.n220 B.n219 585
R238 B.n221 B.n146 585
R239 B.n223 B.n222 585
R240 B.n224 B.n145 585
R241 B.n226 B.n225 585
R242 B.n227 B.n144 585
R243 B.n229 B.n228 585
R244 B.n230 B.n143 585
R245 B.n232 B.n231 585
R246 B.n233 B.n142 585
R247 B.n235 B.n234 585
R248 B.n236 B.n141 585
R249 B.n238 B.n237 585
R250 B.n239 B.n140 585
R251 B.n241 B.n240 585
R252 B.n242 B.n139 585
R253 B.n244 B.n243 585
R254 B.n245 B.n138 585
R255 B.n247 B.n246 585
R256 B.n248 B.n137 585
R257 B.n250 B.n249 585
R258 B.n251 B.n136 585
R259 B.n253 B.n252 585
R260 B.n254 B.n135 585
R261 B.n256 B.n255 585
R262 B.n257 B.n134 585
R263 B.n259 B.n258 585
R264 B.n260 B.n133 585
R265 B.n262 B.n261 585
R266 B.n263 B.n132 585
R267 B.n265 B.n264 585
R268 B.n266 B.n131 585
R269 B.n268 B.n267 585
R270 B.n269 B.n130 585
R271 B.n271 B.n270 585
R272 B.n273 B.n127 585
R273 B.n275 B.n274 585
R274 B.n276 B.n126 585
R275 B.n278 B.n277 585
R276 B.n279 B.n125 585
R277 B.n281 B.n280 585
R278 B.n282 B.n124 585
R279 B.n284 B.n283 585
R280 B.n285 B.n123 585
R281 B.n287 B.n286 585
R282 B.n289 B.n288 585
R283 B.n290 B.n119 585
R284 B.n292 B.n291 585
R285 B.n293 B.n118 585
R286 B.n295 B.n294 585
R287 B.n296 B.n117 585
R288 B.n298 B.n297 585
R289 B.n299 B.n116 585
R290 B.n301 B.n300 585
R291 B.n302 B.n115 585
R292 B.n304 B.n303 585
R293 B.n305 B.n114 585
R294 B.n307 B.n306 585
R295 B.n308 B.n113 585
R296 B.n310 B.n309 585
R297 B.n311 B.n112 585
R298 B.n313 B.n312 585
R299 B.n314 B.n111 585
R300 B.n316 B.n315 585
R301 B.n317 B.n110 585
R302 B.n319 B.n318 585
R303 B.n320 B.n109 585
R304 B.n322 B.n321 585
R305 B.n323 B.n108 585
R306 B.n325 B.n324 585
R307 B.n326 B.n107 585
R308 B.n328 B.n327 585
R309 B.n329 B.n106 585
R310 B.n331 B.n330 585
R311 B.n332 B.n105 585
R312 B.n334 B.n333 585
R313 B.n335 B.n104 585
R314 B.n337 B.n336 585
R315 B.n338 B.n103 585
R316 B.n340 B.n339 585
R317 B.n341 B.n102 585
R318 B.n343 B.n342 585
R319 B.n344 B.n101 585
R320 B.n346 B.n345 585
R321 B.n347 B.n100 585
R322 B.n349 B.n348 585
R323 B.n350 B.n99 585
R324 B.n208 B.n207 585
R325 B.n206 B.n151 585
R326 B.n205 B.n204 585
R327 B.n203 B.n152 585
R328 B.n202 B.n201 585
R329 B.n200 B.n153 585
R330 B.n199 B.n198 585
R331 B.n197 B.n154 585
R332 B.n196 B.n195 585
R333 B.n194 B.n155 585
R334 B.n193 B.n192 585
R335 B.n191 B.n156 585
R336 B.n190 B.n189 585
R337 B.n188 B.n157 585
R338 B.n187 B.n186 585
R339 B.n185 B.n158 585
R340 B.n184 B.n183 585
R341 B.n182 B.n159 585
R342 B.n181 B.n180 585
R343 B.n179 B.n160 585
R344 B.n178 B.n177 585
R345 B.n176 B.n161 585
R346 B.n175 B.n174 585
R347 B.n173 B.n162 585
R348 B.n172 B.n171 585
R349 B.n170 B.n163 585
R350 B.n169 B.n168 585
R351 B.n167 B.n164 585
R352 B.n166 B.n165 585
R353 B.n2 B.n0 585
R354 B.n629 B.n1 585
R355 B.n628 B.n627 585
R356 B.n626 B.n3 585
R357 B.n625 B.n624 585
R358 B.n623 B.n4 585
R359 B.n622 B.n621 585
R360 B.n620 B.n5 585
R361 B.n619 B.n618 585
R362 B.n617 B.n6 585
R363 B.n616 B.n615 585
R364 B.n614 B.n7 585
R365 B.n613 B.n612 585
R366 B.n611 B.n8 585
R367 B.n610 B.n609 585
R368 B.n608 B.n9 585
R369 B.n607 B.n606 585
R370 B.n605 B.n10 585
R371 B.n604 B.n603 585
R372 B.n602 B.n11 585
R373 B.n601 B.n600 585
R374 B.n599 B.n12 585
R375 B.n598 B.n597 585
R376 B.n596 B.n13 585
R377 B.n595 B.n594 585
R378 B.n593 B.n14 585
R379 B.n592 B.n591 585
R380 B.n590 B.n15 585
R381 B.n589 B.n588 585
R382 B.n587 B.n16 585
R383 B.n586 B.n585 585
R384 B.n631 B.n630 585
R385 B.n209 B.n208 497.305
R386 B.n586 B.n17 497.305
R387 B.n352 B.n99 497.305
R388 B.n443 B.n442 497.305
R389 B.n120 B.t0 399.582
R390 B.n128 B.t6 399.582
R391 B.n38 B.t9 399.582
R392 B.n46 B.t3 399.582
R393 B.n208 B.n151 163.367
R394 B.n204 B.n151 163.367
R395 B.n204 B.n203 163.367
R396 B.n203 B.n202 163.367
R397 B.n202 B.n153 163.367
R398 B.n198 B.n153 163.367
R399 B.n198 B.n197 163.367
R400 B.n197 B.n196 163.367
R401 B.n196 B.n155 163.367
R402 B.n192 B.n155 163.367
R403 B.n192 B.n191 163.367
R404 B.n191 B.n190 163.367
R405 B.n190 B.n157 163.367
R406 B.n186 B.n157 163.367
R407 B.n186 B.n185 163.367
R408 B.n185 B.n184 163.367
R409 B.n184 B.n159 163.367
R410 B.n180 B.n159 163.367
R411 B.n180 B.n179 163.367
R412 B.n179 B.n178 163.367
R413 B.n178 B.n161 163.367
R414 B.n174 B.n161 163.367
R415 B.n174 B.n173 163.367
R416 B.n173 B.n172 163.367
R417 B.n172 B.n163 163.367
R418 B.n168 B.n163 163.367
R419 B.n168 B.n167 163.367
R420 B.n167 B.n166 163.367
R421 B.n166 B.n2 163.367
R422 B.n630 B.n2 163.367
R423 B.n630 B.n629 163.367
R424 B.n629 B.n628 163.367
R425 B.n628 B.n3 163.367
R426 B.n624 B.n3 163.367
R427 B.n624 B.n623 163.367
R428 B.n623 B.n622 163.367
R429 B.n622 B.n5 163.367
R430 B.n618 B.n5 163.367
R431 B.n618 B.n617 163.367
R432 B.n617 B.n616 163.367
R433 B.n616 B.n7 163.367
R434 B.n612 B.n7 163.367
R435 B.n612 B.n611 163.367
R436 B.n611 B.n610 163.367
R437 B.n610 B.n9 163.367
R438 B.n606 B.n9 163.367
R439 B.n606 B.n605 163.367
R440 B.n605 B.n604 163.367
R441 B.n604 B.n11 163.367
R442 B.n600 B.n11 163.367
R443 B.n600 B.n599 163.367
R444 B.n599 B.n598 163.367
R445 B.n598 B.n13 163.367
R446 B.n594 B.n13 163.367
R447 B.n594 B.n593 163.367
R448 B.n593 B.n592 163.367
R449 B.n592 B.n15 163.367
R450 B.n588 B.n15 163.367
R451 B.n588 B.n587 163.367
R452 B.n587 B.n586 163.367
R453 B.n210 B.n209 163.367
R454 B.n210 B.n149 163.367
R455 B.n214 B.n149 163.367
R456 B.n215 B.n214 163.367
R457 B.n216 B.n215 163.367
R458 B.n216 B.n147 163.367
R459 B.n220 B.n147 163.367
R460 B.n221 B.n220 163.367
R461 B.n222 B.n221 163.367
R462 B.n222 B.n145 163.367
R463 B.n226 B.n145 163.367
R464 B.n227 B.n226 163.367
R465 B.n228 B.n227 163.367
R466 B.n228 B.n143 163.367
R467 B.n232 B.n143 163.367
R468 B.n233 B.n232 163.367
R469 B.n234 B.n233 163.367
R470 B.n234 B.n141 163.367
R471 B.n238 B.n141 163.367
R472 B.n239 B.n238 163.367
R473 B.n240 B.n239 163.367
R474 B.n240 B.n139 163.367
R475 B.n244 B.n139 163.367
R476 B.n245 B.n244 163.367
R477 B.n246 B.n245 163.367
R478 B.n246 B.n137 163.367
R479 B.n250 B.n137 163.367
R480 B.n251 B.n250 163.367
R481 B.n252 B.n251 163.367
R482 B.n252 B.n135 163.367
R483 B.n256 B.n135 163.367
R484 B.n257 B.n256 163.367
R485 B.n258 B.n257 163.367
R486 B.n258 B.n133 163.367
R487 B.n262 B.n133 163.367
R488 B.n263 B.n262 163.367
R489 B.n264 B.n263 163.367
R490 B.n264 B.n131 163.367
R491 B.n268 B.n131 163.367
R492 B.n269 B.n268 163.367
R493 B.n270 B.n269 163.367
R494 B.n270 B.n127 163.367
R495 B.n275 B.n127 163.367
R496 B.n276 B.n275 163.367
R497 B.n277 B.n276 163.367
R498 B.n277 B.n125 163.367
R499 B.n281 B.n125 163.367
R500 B.n282 B.n281 163.367
R501 B.n283 B.n282 163.367
R502 B.n283 B.n123 163.367
R503 B.n287 B.n123 163.367
R504 B.n288 B.n287 163.367
R505 B.n288 B.n119 163.367
R506 B.n292 B.n119 163.367
R507 B.n293 B.n292 163.367
R508 B.n294 B.n293 163.367
R509 B.n294 B.n117 163.367
R510 B.n298 B.n117 163.367
R511 B.n299 B.n298 163.367
R512 B.n300 B.n299 163.367
R513 B.n300 B.n115 163.367
R514 B.n304 B.n115 163.367
R515 B.n305 B.n304 163.367
R516 B.n306 B.n305 163.367
R517 B.n306 B.n113 163.367
R518 B.n310 B.n113 163.367
R519 B.n311 B.n310 163.367
R520 B.n312 B.n311 163.367
R521 B.n312 B.n111 163.367
R522 B.n316 B.n111 163.367
R523 B.n317 B.n316 163.367
R524 B.n318 B.n317 163.367
R525 B.n318 B.n109 163.367
R526 B.n322 B.n109 163.367
R527 B.n323 B.n322 163.367
R528 B.n324 B.n323 163.367
R529 B.n324 B.n107 163.367
R530 B.n328 B.n107 163.367
R531 B.n329 B.n328 163.367
R532 B.n330 B.n329 163.367
R533 B.n330 B.n105 163.367
R534 B.n334 B.n105 163.367
R535 B.n335 B.n334 163.367
R536 B.n336 B.n335 163.367
R537 B.n336 B.n103 163.367
R538 B.n340 B.n103 163.367
R539 B.n341 B.n340 163.367
R540 B.n342 B.n341 163.367
R541 B.n342 B.n101 163.367
R542 B.n346 B.n101 163.367
R543 B.n347 B.n346 163.367
R544 B.n348 B.n347 163.367
R545 B.n348 B.n99 163.367
R546 B.n353 B.n352 163.367
R547 B.n354 B.n353 163.367
R548 B.n354 B.n97 163.367
R549 B.n358 B.n97 163.367
R550 B.n359 B.n358 163.367
R551 B.n360 B.n359 163.367
R552 B.n360 B.n95 163.367
R553 B.n364 B.n95 163.367
R554 B.n365 B.n364 163.367
R555 B.n366 B.n365 163.367
R556 B.n366 B.n93 163.367
R557 B.n370 B.n93 163.367
R558 B.n371 B.n370 163.367
R559 B.n372 B.n371 163.367
R560 B.n372 B.n91 163.367
R561 B.n376 B.n91 163.367
R562 B.n377 B.n376 163.367
R563 B.n378 B.n377 163.367
R564 B.n378 B.n89 163.367
R565 B.n382 B.n89 163.367
R566 B.n383 B.n382 163.367
R567 B.n384 B.n383 163.367
R568 B.n384 B.n87 163.367
R569 B.n388 B.n87 163.367
R570 B.n389 B.n388 163.367
R571 B.n390 B.n389 163.367
R572 B.n390 B.n85 163.367
R573 B.n394 B.n85 163.367
R574 B.n395 B.n394 163.367
R575 B.n396 B.n395 163.367
R576 B.n396 B.n83 163.367
R577 B.n400 B.n83 163.367
R578 B.n401 B.n400 163.367
R579 B.n402 B.n401 163.367
R580 B.n402 B.n81 163.367
R581 B.n406 B.n81 163.367
R582 B.n407 B.n406 163.367
R583 B.n408 B.n407 163.367
R584 B.n408 B.n79 163.367
R585 B.n412 B.n79 163.367
R586 B.n413 B.n412 163.367
R587 B.n414 B.n413 163.367
R588 B.n414 B.n77 163.367
R589 B.n418 B.n77 163.367
R590 B.n419 B.n418 163.367
R591 B.n420 B.n419 163.367
R592 B.n420 B.n75 163.367
R593 B.n424 B.n75 163.367
R594 B.n425 B.n424 163.367
R595 B.n426 B.n425 163.367
R596 B.n426 B.n73 163.367
R597 B.n430 B.n73 163.367
R598 B.n431 B.n430 163.367
R599 B.n432 B.n431 163.367
R600 B.n432 B.n71 163.367
R601 B.n436 B.n71 163.367
R602 B.n437 B.n436 163.367
R603 B.n438 B.n437 163.367
R604 B.n438 B.n69 163.367
R605 B.n442 B.n69 163.367
R606 B.n582 B.n17 163.367
R607 B.n582 B.n581 163.367
R608 B.n581 B.n580 163.367
R609 B.n580 B.n19 163.367
R610 B.n576 B.n19 163.367
R611 B.n576 B.n575 163.367
R612 B.n575 B.n574 163.367
R613 B.n574 B.n21 163.367
R614 B.n570 B.n21 163.367
R615 B.n570 B.n569 163.367
R616 B.n569 B.n568 163.367
R617 B.n568 B.n23 163.367
R618 B.n564 B.n23 163.367
R619 B.n564 B.n563 163.367
R620 B.n563 B.n562 163.367
R621 B.n562 B.n25 163.367
R622 B.n558 B.n25 163.367
R623 B.n558 B.n557 163.367
R624 B.n557 B.n556 163.367
R625 B.n556 B.n27 163.367
R626 B.n552 B.n27 163.367
R627 B.n552 B.n551 163.367
R628 B.n551 B.n550 163.367
R629 B.n550 B.n29 163.367
R630 B.n546 B.n29 163.367
R631 B.n546 B.n545 163.367
R632 B.n545 B.n544 163.367
R633 B.n544 B.n31 163.367
R634 B.n540 B.n31 163.367
R635 B.n540 B.n539 163.367
R636 B.n539 B.n538 163.367
R637 B.n538 B.n33 163.367
R638 B.n534 B.n33 163.367
R639 B.n534 B.n533 163.367
R640 B.n533 B.n532 163.367
R641 B.n532 B.n35 163.367
R642 B.n528 B.n35 163.367
R643 B.n528 B.n527 163.367
R644 B.n527 B.n526 163.367
R645 B.n526 B.n37 163.367
R646 B.n522 B.n37 163.367
R647 B.n522 B.n521 163.367
R648 B.n521 B.n41 163.367
R649 B.n517 B.n41 163.367
R650 B.n517 B.n516 163.367
R651 B.n516 B.n515 163.367
R652 B.n515 B.n43 163.367
R653 B.n511 B.n43 163.367
R654 B.n511 B.n510 163.367
R655 B.n510 B.n509 163.367
R656 B.n509 B.n45 163.367
R657 B.n504 B.n45 163.367
R658 B.n504 B.n503 163.367
R659 B.n503 B.n502 163.367
R660 B.n502 B.n49 163.367
R661 B.n498 B.n49 163.367
R662 B.n498 B.n497 163.367
R663 B.n497 B.n496 163.367
R664 B.n496 B.n51 163.367
R665 B.n492 B.n51 163.367
R666 B.n492 B.n491 163.367
R667 B.n491 B.n490 163.367
R668 B.n490 B.n53 163.367
R669 B.n486 B.n53 163.367
R670 B.n486 B.n485 163.367
R671 B.n485 B.n484 163.367
R672 B.n484 B.n55 163.367
R673 B.n480 B.n55 163.367
R674 B.n480 B.n479 163.367
R675 B.n479 B.n478 163.367
R676 B.n478 B.n57 163.367
R677 B.n474 B.n57 163.367
R678 B.n474 B.n473 163.367
R679 B.n473 B.n472 163.367
R680 B.n472 B.n59 163.367
R681 B.n468 B.n59 163.367
R682 B.n468 B.n467 163.367
R683 B.n467 B.n466 163.367
R684 B.n466 B.n61 163.367
R685 B.n462 B.n61 163.367
R686 B.n462 B.n461 163.367
R687 B.n461 B.n460 163.367
R688 B.n460 B.n63 163.367
R689 B.n456 B.n63 163.367
R690 B.n456 B.n455 163.367
R691 B.n455 B.n454 163.367
R692 B.n454 B.n65 163.367
R693 B.n450 B.n65 163.367
R694 B.n450 B.n449 163.367
R695 B.n449 B.n448 163.367
R696 B.n448 B.n67 163.367
R697 B.n444 B.n67 163.367
R698 B.n444 B.n443 163.367
R699 B.n120 B.t2 142.929
R700 B.n46 B.t4 142.929
R701 B.n128 B.t8 142.915
R702 B.n38 B.t10 142.915
R703 B.n121 B.t1 107.05
R704 B.n47 B.t5 107.05
R705 B.n129 B.t7 107.035
R706 B.n39 B.t11 107.035
R707 B.n122 B.n121 59.5399
R708 B.n272 B.n129 59.5399
R709 B.n40 B.n39 59.5399
R710 B.n506 B.n47 59.5399
R711 B.n121 B.n120 35.8793
R712 B.n129 B.n128 35.8793
R713 B.n39 B.n38 35.8793
R714 B.n47 B.n46 35.8793
R715 B.n585 B.n584 32.3127
R716 B.n441 B.n68 32.3127
R717 B.n351 B.n350 32.3127
R718 B.n207 B.n150 32.3127
R719 B B.n631 18.0485
R720 B.n584 B.n583 10.6151
R721 B.n583 B.n18 10.6151
R722 B.n579 B.n18 10.6151
R723 B.n579 B.n578 10.6151
R724 B.n578 B.n577 10.6151
R725 B.n577 B.n20 10.6151
R726 B.n573 B.n20 10.6151
R727 B.n573 B.n572 10.6151
R728 B.n572 B.n571 10.6151
R729 B.n571 B.n22 10.6151
R730 B.n567 B.n22 10.6151
R731 B.n567 B.n566 10.6151
R732 B.n566 B.n565 10.6151
R733 B.n565 B.n24 10.6151
R734 B.n561 B.n24 10.6151
R735 B.n561 B.n560 10.6151
R736 B.n560 B.n559 10.6151
R737 B.n559 B.n26 10.6151
R738 B.n555 B.n26 10.6151
R739 B.n555 B.n554 10.6151
R740 B.n554 B.n553 10.6151
R741 B.n553 B.n28 10.6151
R742 B.n549 B.n28 10.6151
R743 B.n549 B.n548 10.6151
R744 B.n548 B.n547 10.6151
R745 B.n547 B.n30 10.6151
R746 B.n543 B.n30 10.6151
R747 B.n543 B.n542 10.6151
R748 B.n542 B.n541 10.6151
R749 B.n541 B.n32 10.6151
R750 B.n537 B.n32 10.6151
R751 B.n537 B.n536 10.6151
R752 B.n536 B.n535 10.6151
R753 B.n535 B.n34 10.6151
R754 B.n531 B.n34 10.6151
R755 B.n531 B.n530 10.6151
R756 B.n530 B.n529 10.6151
R757 B.n529 B.n36 10.6151
R758 B.n525 B.n36 10.6151
R759 B.n525 B.n524 10.6151
R760 B.n524 B.n523 10.6151
R761 B.n520 B.n519 10.6151
R762 B.n519 B.n518 10.6151
R763 B.n518 B.n42 10.6151
R764 B.n514 B.n42 10.6151
R765 B.n514 B.n513 10.6151
R766 B.n513 B.n512 10.6151
R767 B.n512 B.n44 10.6151
R768 B.n508 B.n44 10.6151
R769 B.n508 B.n507 10.6151
R770 B.n505 B.n48 10.6151
R771 B.n501 B.n48 10.6151
R772 B.n501 B.n500 10.6151
R773 B.n500 B.n499 10.6151
R774 B.n499 B.n50 10.6151
R775 B.n495 B.n50 10.6151
R776 B.n495 B.n494 10.6151
R777 B.n494 B.n493 10.6151
R778 B.n493 B.n52 10.6151
R779 B.n489 B.n52 10.6151
R780 B.n489 B.n488 10.6151
R781 B.n488 B.n487 10.6151
R782 B.n487 B.n54 10.6151
R783 B.n483 B.n54 10.6151
R784 B.n483 B.n482 10.6151
R785 B.n482 B.n481 10.6151
R786 B.n481 B.n56 10.6151
R787 B.n477 B.n56 10.6151
R788 B.n477 B.n476 10.6151
R789 B.n476 B.n475 10.6151
R790 B.n475 B.n58 10.6151
R791 B.n471 B.n58 10.6151
R792 B.n471 B.n470 10.6151
R793 B.n470 B.n469 10.6151
R794 B.n469 B.n60 10.6151
R795 B.n465 B.n60 10.6151
R796 B.n465 B.n464 10.6151
R797 B.n464 B.n463 10.6151
R798 B.n463 B.n62 10.6151
R799 B.n459 B.n62 10.6151
R800 B.n459 B.n458 10.6151
R801 B.n458 B.n457 10.6151
R802 B.n457 B.n64 10.6151
R803 B.n453 B.n64 10.6151
R804 B.n453 B.n452 10.6151
R805 B.n452 B.n451 10.6151
R806 B.n451 B.n66 10.6151
R807 B.n447 B.n66 10.6151
R808 B.n447 B.n446 10.6151
R809 B.n446 B.n445 10.6151
R810 B.n445 B.n68 10.6151
R811 B.n351 B.n98 10.6151
R812 B.n355 B.n98 10.6151
R813 B.n356 B.n355 10.6151
R814 B.n357 B.n356 10.6151
R815 B.n357 B.n96 10.6151
R816 B.n361 B.n96 10.6151
R817 B.n362 B.n361 10.6151
R818 B.n363 B.n362 10.6151
R819 B.n363 B.n94 10.6151
R820 B.n367 B.n94 10.6151
R821 B.n368 B.n367 10.6151
R822 B.n369 B.n368 10.6151
R823 B.n369 B.n92 10.6151
R824 B.n373 B.n92 10.6151
R825 B.n374 B.n373 10.6151
R826 B.n375 B.n374 10.6151
R827 B.n375 B.n90 10.6151
R828 B.n379 B.n90 10.6151
R829 B.n380 B.n379 10.6151
R830 B.n381 B.n380 10.6151
R831 B.n381 B.n88 10.6151
R832 B.n385 B.n88 10.6151
R833 B.n386 B.n385 10.6151
R834 B.n387 B.n386 10.6151
R835 B.n387 B.n86 10.6151
R836 B.n391 B.n86 10.6151
R837 B.n392 B.n391 10.6151
R838 B.n393 B.n392 10.6151
R839 B.n393 B.n84 10.6151
R840 B.n397 B.n84 10.6151
R841 B.n398 B.n397 10.6151
R842 B.n399 B.n398 10.6151
R843 B.n399 B.n82 10.6151
R844 B.n403 B.n82 10.6151
R845 B.n404 B.n403 10.6151
R846 B.n405 B.n404 10.6151
R847 B.n405 B.n80 10.6151
R848 B.n409 B.n80 10.6151
R849 B.n410 B.n409 10.6151
R850 B.n411 B.n410 10.6151
R851 B.n411 B.n78 10.6151
R852 B.n415 B.n78 10.6151
R853 B.n416 B.n415 10.6151
R854 B.n417 B.n416 10.6151
R855 B.n417 B.n76 10.6151
R856 B.n421 B.n76 10.6151
R857 B.n422 B.n421 10.6151
R858 B.n423 B.n422 10.6151
R859 B.n423 B.n74 10.6151
R860 B.n427 B.n74 10.6151
R861 B.n428 B.n427 10.6151
R862 B.n429 B.n428 10.6151
R863 B.n429 B.n72 10.6151
R864 B.n433 B.n72 10.6151
R865 B.n434 B.n433 10.6151
R866 B.n435 B.n434 10.6151
R867 B.n435 B.n70 10.6151
R868 B.n439 B.n70 10.6151
R869 B.n440 B.n439 10.6151
R870 B.n441 B.n440 10.6151
R871 B.n211 B.n150 10.6151
R872 B.n212 B.n211 10.6151
R873 B.n213 B.n212 10.6151
R874 B.n213 B.n148 10.6151
R875 B.n217 B.n148 10.6151
R876 B.n218 B.n217 10.6151
R877 B.n219 B.n218 10.6151
R878 B.n219 B.n146 10.6151
R879 B.n223 B.n146 10.6151
R880 B.n224 B.n223 10.6151
R881 B.n225 B.n224 10.6151
R882 B.n225 B.n144 10.6151
R883 B.n229 B.n144 10.6151
R884 B.n230 B.n229 10.6151
R885 B.n231 B.n230 10.6151
R886 B.n231 B.n142 10.6151
R887 B.n235 B.n142 10.6151
R888 B.n236 B.n235 10.6151
R889 B.n237 B.n236 10.6151
R890 B.n237 B.n140 10.6151
R891 B.n241 B.n140 10.6151
R892 B.n242 B.n241 10.6151
R893 B.n243 B.n242 10.6151
R894 B.n243 B.n138 10.6151
R895 B.n247 B.n138 10.6151
R896 B.n248 B.n247 10.6151
R897 B.n249 B.n248 10.6151
R898 B.n249 B.n136 10.6151
R899 B.n253 B.n136 10.6151
R900 B.n254 B.n253 10.6151
R901 B.n255 B.n254 10.6151
R902 B.n255 B.n134 10.6151
R903 B.n259 B.n134 10.6151
R904 B.n260 B.n259 10.6151
R905 B.n261 B.n260 10.6151
R906 B.n261 B.n132 10.6151
R907 B.n265 B.n132 10.6151
R908 B.n266 B.n265 10.6151
R909 B.n267 B.n266 10.6151
R910 B.n267 B.n130 10.6151
R911 B.n271 B.n130 10.6151
R912 B.n274 B.n273 10.6151
R913 B.n274 B.n126 10.6151
R914 B.n278 B.n126 10.6151
R915 B.n279 B.n278 10.6151
R916 B.n280 B.n279 10.6151
R917 B.n280 B.n124 10.6151
R918 B.n284 B.n124 10.6151
R919 B.n285 B.n284 10.6151
R920 B.n286 B.n285 10.6151
R921 B.n290 B.n289 10.6151
R922 B.n291 B.n290 10.6151
R923 B.n291 B.n118 10.6151
R924 B.n295 B.n118 10.6151
R925 B.n296 B.n295 10.6151
R926 B.n297 B.n296 10.6151
R927 B.n297 B.n116 10.6151
R928 B.n301 B.n116 10.6151
R929 B.n302 B.n301 10.6151
R930 B.n303 B.n302 10.6151
R931 B.n303 B.n114 10.6151
R932 B.n307 B.n114 10.6151
R933 B.n308 B.n307 10.6151
R934 B.n309 B.n308 10.6151
R935 B.n309 B.n112 10.6151
R936 B.n313 B.n112 10.6151
R937 B.n314 B.n313 10.6151
R938 B.n315 B.n314 10.6151
R939 B.n315 B.n110 10.6151
R940 B.n319 B.n110 10.6151
R941 B.n320 B.n319 10.6151
R942 B.n321 B.n320 10.6151
R943 B.n321 B.n108 10.6151
R944 B.n325 B.n108 10.6151
R945 B.n326 B.n325 10.6151
R946 B.n327 B.n326 10.6151
R947 B.n327 B.n106 10.6151
R948 B.n331 B.n106 10.6151
R949 B.n332 B.n331 10.6151
R950 B.n333 B.n332 10.6151
R951 B.n333 B.n104 10.6151
R952 B.n337 B.n104 10.6151
R953 B.n338 B.n337 10.6151
R954 B.n339 B.n338 10.6151
R955 B.n339 B.n102 10.6151
R956 B.n343 B.n102 10.6151
R957 B.n344 B.n343 10.6151
R958 B.n345 B.n344 10.6151
R959 B.n345 B.n100 10.6151
R960 B.n349 B.n100 10.6151
R961 B.n350 B.n349 10.6151
R962 B.n207 B.n206 10.6151
R963 B.n206 B.n205 10.6151
R964 B.n205 B.n152 10.6151
R965 B.n201 B.n152 10.6151
R966 B.n201 B.n200 10.6151
R967 B.n200 B.n199 10.6151
R968 B.n199 B.n154 10.6151
R969 B.n195 B.n154 10.6151
R970 B.n195 B.n194 10.6151
R971 B.n194 B.n193 10.6151
R972 B.n193 B.n156 10.6151
R973 B.n189 B.n156 10.6151
R974 B.n189 B.n188 10.6151
R975 B.n188 B.n187 10.6151
R976 B.n187 B.n158 10.6151
R977 B.n183 B.n158 10.6151
R978 B.n183 B.n182 10.6151
R979 B.n182 B.n181 10.6151
R980 B.n181 B.n160 10.6151
R981 B.n177 B.n160 10.6151
R982 B.n177 B.n176 10.6151
R983 B.n176 B.n175 10.6151
R984 B.n175 B.n162 10.6151
R985 B.n171 B.n162 10.6151
R986 B.n171 B.n170 10.6151
R987 B.n170 B.n169 10.6151
R988 B.n169 B.n164 10.6151
R989 B.n165 B.n164 10.6151
R990 B.n165 B.n0 10.6151
R991 B.n627 B.n1 10.6151
R992 B.n627 B.n626 10.6151
R993 B.n626 B.n625 10.6151
R994 B.n625 B.n4 10.6151
R995 B.n621 B.n4 10.6151
R996 B.n621 B.n620 10.6151
R997 B.n620 B.n619 10.6151
R998 B.n619 B.n6 10.6151
R999 B.n615 B.n6 10.6151
R1000 B.n615 B.n614 10.6151
R1001 B.n614 B.n613 10.6151
R1002 B.n613 B.n8 10.6151
R1003 B.n609 B.n8 10.6151
R1004 B.n609 B.n608 10.6151
R1005 B.n608 B.n607 10.6151
R1006 B.n607 B.n10 10.6151
R1007 B.n603 B.n10 10.6151
R1008 B.n603 B.n602 10.6151
R1009 B.n602 B.n601 10.6151
R1010 B.n601 B.n12 10.6151
R1011 B.n597 B.n12 10.6151
R1012 B.n597 B.n596 10.6151
R1013 B.n596 B.n595 10.6151
R1014 B.n595 B.n14 10.6151
R1015 B.n591 B.n14 10.6151
R1016 B.n591 B.n590 10.6151
R1017 B.n590 B.n589 10.6151
R1018 B.n589 B.n16 10.6151
R1019 B.n585 B.n16 10.6151
R1020 B.n523 B.n40 9.36635
R1021 B.n506 B.n505 9.36635
R1022 B.n272 B.n271 9.36635
R1023 B.n289 B.n122 9.36635
R1024 B.n631 B.n0 2.81026
R1025 B.n631 B.n1 2.81026
R1026 B.n520 B.n40 1.24928
R1027 B.n507 B.n506 1.24928
R1028 B.n273 B.n272 1.24928
R1029 B.n286 B.n122 1.24928
R1030 VP.n6 VP.t0 224.964
R1031 VP.n17 VP.t3 194.069
R1032 VP.n24 VP.t2 194.069
R1033 VP.n31 VP.t1 194.069
R1034 VP.n14 VP.t5 194.069
R1035 VP.n7 VP.t4 194.069
R1036 VP.n17 VP.n16 180.775
R1037 VP.n32 VP.n31 180.775
R1038 VP.n15 VP.n14 180.775
R1039 VP.n9 VP.n8 161.3
R1040 VP.n10 VP.n5 161.3
R1041 VP.n12 VP.n11 161.3
R1042 VP.n13 VP.n4 161.3
R1043 VP.n30 VP.n0 161.3
R1044 VP.n29 VP.n28 161.3
R1045 VP.n27 VP.n1 161.3
R1046 VP.n26 VP.n25 161.3
R1047 VP.n23 VP.n2 161.3
R1048 VP.n22 VP.n21 161.3
R1049 VP.n20 VP.n3 161.3
R1050 VP.n19 VP.n18 161.3
R1051 VP.n22 VP.n3 56.4773
R1052 VP.n29 VP.n1 56.4773
R1053 VP.n12 VP.n5 56.4773
R1054 VP.n7 VP.n6 53.4877
R1055 VP.n16 VP.n15 44.474
R1056 VP.n18 VP.n3 24.3439
R1057 VP.n23 VP.n22 24.3439
R1058 VP.n25 VP.n1 24.3439
R1059 VP.n30 VP.n29 24.3439
R1060 VP.n13 VP.n12 24.3439
R1061 VP.n8 VP.n5 24.3439
R1062 VP.n9 VP.n6 18.3124
R1063 VP.n24 VP.n23 12.1722
R1064 VP.n25 VP.n24 12.1722
R1065 VP.n8 VP.n7 12.1722
R1066 VP.n18 VP.n17 4.86919
R1067 VP.n31 VP.n30 4.86919
R1068 VP.n14 VP.n13 4.86919
R1069 VP.n10 VP.n9 0.189894
R1070 VP.n11 VP.n10 0.189894
R1071 VP.n11 VP.n4 0.189894
R1072 VP.n15 VP.n4 0.189894
R1073 VP.n19 VP.n16 0.189894
R1074 VP.n20 VP.n19 0.189894
R1075 VP.n21 VP.n20 0.189894
R1076 VP.n21 VP.n2 0.189894
R1077 VP.n26 VP.n2 0.189894
R1078 VP.n27 VP.n26 0.189894
R1079 VP.n28 VP.n27 0.189894
R1080 VP.n28 VP.n0 0.189894
R1081 VP.n32 VP.n0 0.189894
R1082 VP VP.n32 0.0516364
R1083 VDD1 VDD1.t5 79.2606
R1084 VDD1.n1 VDD1.t2 79.146
R1085 VDD1.n1 VDD1.n0 75.6938
R1086 VDD1.n3 VDD1.n2 75.3495
R1087 VDD1.n3 VDD1.n1 40.8306
R1088 VDD1.n2 VDD1.t1 2.65614
R1089 VDD1.n2 VDD1.t0 2.65614
R1090 VDD1.n0 VDD1.t3 2.65614
R1091 VDD1.n0 VDD1.t4 2.65614
R1092 VDD1 VDD1.n3 0.341017
C0 VDD1 w_n2450_n3416# 2.04388f
C1 VDD1 VTAIL 8.084949f
C2 B VDD2 1.8671f
C3 VN w_n2450_n3416# 4.39439f
C4 VN VTAIL 5.90751f
C5 B VP 1.45701f
C6 VDD1 VN 0.148997f
C7 VDD2 w_n2450_n3416# 2.09421f
C8 VDD2 VTAIL 8.12682f
C9 w_n2450_n3416# VP 4.70813f
C10 VDD2 VDD1 1.0152f
C11 VTAIL VP 5.92193f
C12 VDD1 VP 6.22331f
C13 VDD2 VN 6.00942f
C14 VN VP 5.92826f
C15 B w_n2450_n3416# 8.252f
C16 B VTAIL 3.24425f
C17 B VDD1 1.81879f
C18 B VN 0.938628f
C19 VDD2 VP 0.366636f
C20 VTAIL w_n2450_n3416# 2.94571f
C21 VDD2 VSUBS 1.521332f
C22 VDD1 VSUBS 1.900837f
C23 VTAIL VSUBS 0.981912f
C24 VN VSUBS 4.88499f
C25 VP VSUBS 2.094204f
C26 B VSUBS 3.589444f
C27 w_n2450_n3416# VSUBS 0.102988p
C28 VDD1.t5 VSUBS 2.49193f
C29 VDD1.t2 VSUBS 2.49091f
C30 VDD1.t3 VSUBS 0.24086f
C31 VDD1.t4 VSUBS 0.24086f
C32 VDD1.n0 VSUBS 1.90668f
C33 VDD1.n1 VSUBS 3.04425f
C34 VDD1.t1 VSUBS 0.24086f
C35 VDD1.t0 VSUBS 0.24086f
C36 VDD1.n2 VSUBS 1.90387f
C37 VDD1.n3 VSUBS 2.74014f
C38 VP.n0 VSUBS 0.040963f
C39 VP.t1 VSUBS 2.0776f
C40 VP.n1 VSUBS 0.051437f
C41 VP.n2 VSUBS 0.040963f
C42 VP.t2 VSUBS 2.0776f
C43 VP.n3 VSUBS 0.06868f
C44 VP.n4 VSUBS 0.040963f
C45 VP.t5 VSUBS 2.0776f
C46 VP.n5 VSUBS 0.051437f
C47 VP.t0 VSUBS 2.20246f
C48 VP.n6 VSUBS 0.852785f
C49 VP.t4 VSUBS 2.0776f
C50 VP.n7 VSUBS 0.827075f
C51 VP.n8 VSUBS 0.057785f
C52 VP.n9 VSUBS 0.256357f
C53 VP.n10 VSUBS 0.040963f
C54 VP.n11 VSUBS 0.040963f
C55 VP.n12 VSUBS 0.06868f
C56 VP.n13 VSUBS 0.04642f
C57 VP.n14 VSUBS 0.826377f
C58 VP.n15 VSUBS 1.86603f
C59 VP.n16 VSUBS 1.89904f
C60 VP.t3 VSUBS 2.0776f
C61 VP.n17 VSUBS 0.826377f
C62 VP.n18 VSUBS 0.04642f
C63 VP.n19 VSUBS 0.040963f
C64 VP.n20 VSUBS 0.040963f
C65 VP.n21 VSUBS 0.040963f
C66 VP.n22 VSUBS 0.051437f
C67 VP.n23 VSUBS 0.057785f
C68 VP.n24 VSUBS 0.749804f
C69 VP.n25 VSUBS 0.057785f
C70 VP.n26 VSUBS 0.040963f
C71 VP.n27 VSUBS 0.040963f
C72 VP.n28 VSUBS 0.040963f
C73 VP.n29 VSUBS 0.06868f
C74 VP.n30 VSUBS 0.04642f
C75 VP.n31 VSUBS 0.826377f
C76 VP.n32 VSUBS 0.04099f
C77 B.n0 VSUBS 0.004218f
C78 B.n1 VSUBS 0.004218f
C79 B.n2 VSUBS 0.00667f
C80 B.n3 VSUBS 0.00667f
C81 B.n4 VSUBS 0.00667f
C82 B.n5 VSUBS 0.00667f
C83 B.n6 VSUBS 0.00667f
C84 B.n7 VSUBS 0.00667f
C85 B.n8 VSUBS 0.00667f
C86 B.n9 VSUBS 0.00667f
C87 B.n10 VSUBS 0.00667f
C88 B.n11 VSUBS 0.00667f
C89 B.n12 VSUBS 0.00667f
C90 B.n13 VSUBS 0.00667f
C91 B.n14 VSUBS 0.00667f
C92 B.n15 VSUBS 0.00667f
C93 B.n16 VSUBS 0.00667f
C94 B.n17 VSUBS 0.015722f
C95 B.n18 VSUBS 0.00667f
C96 B.n19 VSUBS 0.00667f
C97 B.n20 VSUBS 0.00667f
C98 B.n21 VSUBS 0.00667f
C99 B.n22 VSUBS 0.00667f
C100 B.n23 VSUBS 0.00667f
C101 B.n24 VSUBS 0.00667f
C102 B.n25 VSUBS 0.00667f
C103 B.n26 VSUBS 0.00667f
C104 B.n27 VSUBS 0.00667f
C105 B.n28 VSUBS 0.00667f
C106 B.n29 VSUBS 0.00667f
C107 B.n30 VSUBS 0.00667f
C108 B.n31 VSUBS 0.00667f
C109 B.n32 VSUBS 0.00667f
C110 B.n33 VSUBS 0.00667f
C111 B.n34 VSUBS 0.00667f
C112 B.n35 VSUBS 0.00667f
C113 B.n36 VSUBS 0.00667f
C114 B.n37 VSUBS 0.00667f
C115 B.t11 VSUBS 0.380868f
C116 B.t10 VSUBS 0.394597f
C117 B.t9 VSUBS 0.775153f
C118 B.n38 VSUBS 0.175862f
C119 B.n39 VSUBS 0.064196f
C120 B.n40 VSUBS 0.015454f
C121 B.n41 VSUBS 0.00667f
C122 B.n42 VSUBS 0.00667f
C123 B.n43 VSUBS 0.00667f
C124 B.n44 VSUBS 0.00667f
C125 B.n45 VSUBS 0.00667f
C126 B.t5 VSUBS 0.380861f
C127 B.t4 VSUBS 0.394589f
C128 B.t3 VSUBS 0.775153f
C129 B.n46 VSUBS 0.175869f
C130 B.n47 VSUBS 0.064204f
C131 B.n48 VSUBS 0.00667f
C132 B.n49 VSUBS 0.00667f
C133 B.n50 VSUBS 0.00667f
C134 B.n51 VSUBS 0.00667f
C135 B.n52 VSUBS 0.00667f
C136 B.n53 VSUBS 0.00667f
C137 B.n54 VSUBS 0.00667f
C138 B.n55 VSUBS 0.00667f
C139 B.n56 VSUBS 0.00667f
C140 B.n57 VSUBS 0.00667f
C141 B.n58 VSUBS 0.00667f
C142 B.n59 VSUBS 0.00667f
C143 B.n60 VSUBS 0.00667f
C144 B.n61 VSUBS 0.00667f
C145 B.n62 VSUBS 0.00667f
C146 B.n63 VSUBS 0.00667f
C147 B.n64 VSUBS 0.00667f
C148 B.n65 VSUBS 0.00667f
C149 B.n66 VSUBS 0.00667f
C150 B.n67 VSUBS 0.00667f
C151 B.n68 VSUBS 0.014925f
C152 B.n69 VSUBS 0.00667f
C153 B.n70 VSUBS 0.00667f
C154 B.n71 VSUBS 0.00667f
C155 B.n72 VSUBS 0.00667f
C156 B.n73 VSUBS 0.00667f
C157 B.n74 VSUBS 0.00667f
C158 B.n75 VSUBS 0.00667f
C159 B.n76 VSUBS 0.00667f
C160 B.n77 VSUBS 0.00667f
C161 B.n78 VSUBS 0.00667f
C162 B.n79 VSUBS 0.00667f
C163 B.n80 VSUBS 0.00667f
C164 B.n81 VSUBS 0.00667f
C165 B.n82 VSUBS 0.00667f
C166 B.n83 VSUBS 0.00667f
C167 B.n84 VSUBS 0.00667f
C168 B.n85 VSUBS 0.00667f
C169 B.n86 VSUBS 0.00667f
C170 B.n87 VSUBS 0.00667f
C171 B.n88 VSUBS 0.00667f
C172 B.n89 VSUBS 0.00667f
C173 B.n90 VSUBS 0.00667f
C174 B.n91 VSUBS 0.00667f
C175 B.n92 VSUBS 0.00667f
C176 B.n93 VSUBS 0.00667f
C177 B.n94 VSUBS 0.00667f
C178 B.n95 VSUBS 0.00667f
C179 B.n96 VSUBS 0.00667f
C180 B.n97 VSUBS 0.00667f
C181 B.n98 VSUBS 0.00667f
C182 B.n99 VSUBS 0.015722f
C183 B.n100 VSUBS 0.00667f
C184 B.n101 VSUBS 0.00667f
C185 B.n102 VSUBS 0.00667f
C186 B.n103 VSUBS 0.00667f
C187 B.n104 VSUBS 0.00667f
C188 B.n105 VSUBS 0.00667f
C189 B.n106 VSUBS 0.00667f
C190 B.n107 VSUBS 0.00667f
C191 B.n108 VSUBS 0.00667f
C192 B.n109 VSUBS 0.00667f
C193 B.n110 VSUBS 0.00667f
C194 B.n111 VSUBS 0.00667f
C195 B.n112 VSUBS 0.00667f
C196 B.n113 VSUBS 0.00667f
C197 B.n114 VSUBS 0.00667f
C198 B.n115 VSUBS 0.00667f
C199 B.n116 VSUBS 0.00667f
C200 B.n117 VSUBS 0.00667f
C201 B.n118 VSUBS 0.00667f
C202 B.n119 VSUBS 0.00667f
C203 B.t1 VSUBS 0.380861f
C204 B.t2 VSUBS 0.394589f
C205 B.t0 VSUBS 0.775153f
C206 B.n120 VSUBS 0.175869f
C207 B.n121 VSUBS 0.064204f
C208 B.n122 VSUBS 0.015454f
C209 B.n123 VSUBS 0.00667f
C210 B.n124 VSUBS 0.00667f
C211 B.n125 VSUBS 0.00667f
C212 B.n126 VSUBS 0.00667f
C213 B.n127 VSUBS 0.00667f
C214 B.t7 VSUBS 0.380868f
C215 B.t8 VSUBS 0.394597f
C216 B.t6 VSUBS 0.775153f
C217 B.n128 VSUBS 0.175862f
C218 B.n129 VSUBS 0.064196f
C219 B.n130 VSUBS 0.00667f
C220 B.n131 VSUBS 0.00667f
C221 B.n132 VSUBS 0.00667f
C222 B.n133 VSUBS 0.00667f
C223 B.n134 VSUBS 0.00667f
C224 B.n135 VSUBS 0.00667f
C225 B.n136 VSUBS 0.00667f
C226 B.n137 VSUBS 0.00667f
C227 B.n138 VSUBS 0.00667f
C228 B.n139 VSUBS 0.00667f
C229 B.n140 VSUBS 0.00667f
C230 B.n141 VSUBS 0.00667f
C231 B.n142 VSUBS 0.00667f
C232 B.n143 VSUBS 0.00667f
C233 B.n144 VSUBS 0.00667f
C234 B.n145 VSUBS 0.00667f
C235 B.n146 VSUBS 0.00667f
C236 B.n147 VSUBS 0.00667f
C237 B.n148 VSUBS 0.00667f
C238 B.n149 VSUBS 0.00667f
C239 B.n150 VSUBS 0.015722f
C240 B.n151 VSUBS 0.00667f
C241 B.n152 VSUBS 0.00667f
C242 B.n153 VSUBS 0.00667f
C243 B.n154 VSUBS 0.00667f
C244 B.n155 VSUBS 0.00667f
C245 B.n156 VSUBS 0.00667f
C246 B.n157 VSUBS 0.00667f
C247 B.n158 VSUBS 0.00667f
C248 B.n159 VSUBS 0.00667f
C249 B.n160 VSUBS 0.00667f
C250 B.n161 VSUBS 0.00667f
C251 B.n162 VSUBS 0.00667f
C252 B.n163 VSUBS 0.00667f
C253 B.n164 VSUBS 0.00667f
C254 B.n165 VSUBS 0.00667f
C255 B.n166 VSUBS 0.00667f
C256 B.n167 VSUBS 0.00667f
C257 B.n168 VSUBS 0.00667f
C258 B.n169 VSUBS 0.00667f
C259 B.n170 VSUBS 0.00667f
C260 B.n171 VSUBS 0.00667f
C261 B.n172 VSUBS 0.00667f
C262 B.n173 VSUBS 0.00667f
C263 B.n174 VSUBS 0.00667f
C264 B.n175 VSUBS 0.00667f
C265 B.n176 VSUBS 0.00667f
C266 B.n177 VSUBS 0.00667f
C267 B.n178 VSUBS 0.00667f
C268 B.n179 VSUBS 0.00667f
C269 B.n180 VSUBS 0.00667f
C270 B.n181 VSUBS 0.00667f
C271 B.n182 VSUBS 0.00667f
C272 B.n183 VSUBS 0.00667f
C273 B.n184 VSUBS 0.00667f
C274 B.n185 VSUBS 0.00667f
C275 B.n186 VSUBS 0.00667f
C276 B.n187 VSUBS 0.00667f
C277 B.n188 VSUBS 0.00667f
C278 B.n189 VSUBS 0.00667f
C279 B.n190 VSUBS 0.00667f
C280 B.n191 VSUBS 0.00667f
C281 B.n192 VSUBS 0.00667f
C282 B.n193 VSUBS 0.00667f
C283 B.n194 VSUBS 0.00667f
C284 B.n195 VSUBS 0.00667f
C285 B.n196 VSUBS 0.00667f
C286 B.n197 VSUBS 0.00667f
C287 B.n198 VSUBS 0.00667f
C288 B.n199 VSUBS 0.00667f
C289 B.n200 VSUBS 0.00667f
C290 B.n201 VSUBS 0.00667f
C291 B.n202 VSUBS 0.00667f
C292 B.n203 VSUBS 0.00667f
C293 B.n204 VSUBS 0.00667f
C294 B.n205 VSUBS 0.00667f
C295 B.n206 VSUBS 0.00667f
C296 B.n207 VSUBS 0.015275f
C297 B.n208 VSUBS 0.015275f
C298 B.n209 VSUBS 0.015722f
C299 B.n210 VSUBS 0.00667f
C300 B.n211 VSUBS 0.00667f
C301 B.n212 VSUBS 0.00667f
C302 B.n213 VSUBS 0.00667f
C303 B.n214 VSUBS 0.00667f
C304 B.n215 VSUBS 0.00667f
C305 B.n216 VSUBS 0.00667f
C306 B.n217 VSUBS 0.00667f
C307 B.n218 VSUBS 0.00667f
C308 B.n219 VSUBS 0.00667f
C309 B.n220 VSUBS 0.00667f
C310 B.n221 VSUBS 0.00667f
C311 B.n222 VSUBS 0.00667f
C312 B.n223 VSUBS 0.00667f
C313 B.n224 VSUBS 0.00667f
C314 B.n225 VSUBS 0.00667f
C315 B.n226 VSUBS 0.00667f
C316 B.n227 VSUBS 0.00667f
C317 B.n228 VSUBS 0.00667f
C318 B.n229 VSUBS 0.00667f
C319 B.n230 VSUBS 0.00667f
C320 B.n231 VSUBS 0.00667f
C321 B.n232 VSUBS 0.00667f
C322 B.n233 VSUBS 0.00667f
C323 B.n234 VSUBS 0.00667f
C324 B.n235 VSUBS 0.00667f
C325 B.n236 VSUBS 0.00667f
C326 B.n237 VSUBS 0.00667f
C327 B.n238 VSUBS 0.00667f
C328 B.n239 VSUBS 0.00667f
C329 B.n240 VSUBS 0.00667f
C330 B.n241 VSUBS 0.00667f
C331 B.n242 VSUBS 0.00667f
C332 B.n243 VSUBS 0.00667f
C333 B.n244 VSUBS 0.00667f
C334 B.n245 VSUBS 0.00667f
C335 B.n246 VSUBS 0.00667f
C336 B.n247 VSUBS 0.00667f
C337 B.n248 VSUBS 0.00667f
C338 B.n249 VSUBS 0.00667f
C339 B.n250 VSUBS 0.00667f
C340 B.n251 VSUBS 0.00667f
C341 B.n252 VSUBS 0.00667f
C342 B.n253 VSUBS 0.00667f
C343 B.n254 VSUBS 0.00667f
C344 B.n255 VSUBS 0.00667f
C345 B.n256 VSUBS 0.00667f
C346 B.n257 VSUBS 0.00667f
C347 B.n258 VSUBS 0.00667f
C348 B.n259 VSUBS 0.00667f
C349 B.n260 VSUBS 0.00667f
C350 B.n261 VSUBS 0.00667f
C351 B.n262 VSUBS 0.00667f
C352 B.n263 VSUBS 0.00667f
C353 B.n264 VSUBS 0.00667f
C354 B.n265 VSUBS 0.00667f
C355 B.n266 VSUBS 0.00667f
C356 B.n267 VSUBS 0.00667f
C357 B.n268 VSUBS 0.00667f
C358 B.n269 VSUBS 0.00667f
C359 B.n270 VSUBS 0.00667f
C360 B.n271 VSUBS 0.006278f
C361 B.n272 VSUBS 0.015454f
C362 B.n273 VSUBS 0.003728f
C363 B.n274 VSUBS 0.00667f
C364 B.n275 VSUBS 0.00667f
C365 B.n276 VSUBS 0.00667f
C366 B.n277 VSUBS 0.00667f
C367 B.n278 VSUBS 0.00667f
C368 B.n279 VSUBS 0.00667f
C369 B.n280 VSUBS 0.00667f
C370 B.n281 VSUBS 0.00667f
C371 B.n282 VSUBS 0.00667f
C372 B.n283 VSUBS 0.00667f
C373 B.n284 VSUBS 0.00667f
C374 B.n285 VSUBS 0.00667f
C375 B.n286 VSUBS 0.003728f
C376 B.n287 VSUBS 0.00667f
C377 B.n288 VSUBS 0.00667f
C378 B.n289 VSUBS 0.006278f
C379 B.n290 VSUBS 0.00667f
C380 B.n291 VSUBS 0.00667f
C381 B.n292 VSUBS 0.00667f
C382 B.n293 VSUBS 0.00667f
C383 B.n294 VSUBS 0.00667f
C384 B.n295 VSUBS 0.00667f
C385 B.n296 VSUBS 0.00667f
C386 B.n297 VSUBS 0.00667f
C387 B.n298 VSUBS 0.00667f
C388 B.n299 VSUBS 0.00667f
C389 B.n300 VSUBS 0.00667f
C390 B.n301 VSUBS 0.00667f
C391 B.n302 VSUBS 0.00667f
C392 B.n303 VSUBS 0.00667f
C393 B.n304 VSUBS 0.00667f
C394 B.n305 VSUBS 0.00667f
C395 B.n306 VSUBS 0.00667f
C396 B.n307 VSUBS 0.00667f
C397 B.n308 VSUBS 0.00667f
C398 B.n309 VSUBS 0.00667f
C399 B.n310 VSUBS 0.00667f
C400 B.n311 VSUBS 0.00667f
C401 B.n312 VSUBS 0.00667f
C402 B.n313 VSUBS 0.00667f
C403 B.n314 VSUBS 0.00667f
C404 B.n315 VSUBS 0.00667f
C405 B.n316 VSUBS 0.00667f
C406 B.n317 VSUBS 0.00667f
C407 B.n318 VSUBS 0.00667f
C408 B.n319 VSUBS 0.00667f
C409 B.n320 VSUBS 0.00667f
C410 B.n321 VSUBS 0.00667f
C411 B.n322 VSUBS 0.00667f
C412 B.n323 VSUBS 0.00667f
C413 B.n324 VSUBS 0.00667f
C414 B.n325 VSUBS 0.00667f
C415 B.n326 VSUBS 0.00667f
C416 B.n327 VSUBS 0.00667f
C417 B.n328 VSUBS 0.00667f
C418 B.n329 VSUBS 0.00667f
C419 B.n330 VSUBS 0.00667f
C420 B.n331 VSUBS 0.00667f
C421 B.n332 VSUBS 0.00667f
C422 B.n333 VSUBS 0.00667f
C423 B.n334 VSUBS 0.00667f
C424 B.n335 VSUBS 0.00667f
C425 B.n336 VSUBS 0.00667f
C426 B.n337 VSUBS 0.00667f
C427 B.n338 VSUBS 0.00667f
C428 B.n339 VSUBS 0.00667f
C429 B.n340 VSUBS 0.00667f
C430 B.n341 VSUBS 0.00667f
C431 B.n342 VSUBS 0.00667f
C432 B.n343 VSUBS 0.00667f
C433 B.n344 VSUBS 0.00667f
C434 B.n345 VSUBS 0.00667f
C435 B.n346 VSUBS 0.00667f
C436 B.n347 VSUBS 0.00667f
C437 B.n348 VSUBS 0.00667f
C438 B.n349 VSUBS 0.00667f
C439 B.n350 VSUBS 0.015722f
C440 B.n351 VSUBS 0.015275f
C441 B.n352 VSUBS 0.015275f
C442 B.n353 VSUBS 0.00667f
C443 B.n354 VSUBS 0.00667f
C444 B.n355 VSUBS 0.00667f
C445 B.n356 VSUBS 0.00667f
C446 B.n357 VSUBS 0.00667f
C447 B.n358 VSUBS 0.00667f
C448 B.n359 VSUBS 0.00667f
C449 B.n360 VSUBS 0.00667f
C450 B.n361 VSUBS 0.00667f
C451 B.n362 VSUBS 0.00667f
C452 B.n363 VSUBS 0.00667f
C453 B.n364 VSUBS 0.00667f
C454 B.n365 VSUBS 0.00667f
C455 B.n366 VSUBS 0.00667f
C456 B.n367 VSUBS 0.00667f
C457 B.n368 VSUBS 0.00667f
C458 B.n369 VSUBS 0.00667f
C459 B.n370 VSUBS 0.00667f
C460 B.n371 VSUBS 0.00667f
C461 B.n372 VSUBS 0.00667f
C462 B.n373 VSUBS 0.00667f
C463 B.n374 VSUBS 0.00667f
C464 B.n375 VSUBS 0.00667f
C465 B.n376 VSUBS 0.00667f
C466 B.n377 VSUBS 0.00667f
C467 B.n378 VSUBS 0.00667f
C468 B.n379 VSUBS 0.00667f
C469 B.n380 VSUBS 0.00667f
C470 B.n381 VSUBS 0.00667f
C471 B.n382 VSUBS 0.00667f
C472 B.n383 VSUBS 0.00667f
C473 B.n384 VSUBS 0.00667f
C474 B.n385 VSUBS 0.00667f
C475 B.n386 VSUBS 0.00667f
C476 B.n387 VSUBS 0.00667f
C477 B.n388 VSUBS 0.00667f
C478 B.n389 VSUBS 0.00667f
C479 B.n390 VSUBS 0.00667f
C480 B.n391 VSUBS 0.00667f
C481 B.n392 VSUBS 0.00667f
C482 B.n393 VSUBS 0.00667f
C483 B.n394 VSUBS 0.00667f
C484 B.n395 VSUBS 0.00667f
C485 B.n396 VSUBS 0.00667f
C486 B.n397 VSUBS 0.00667f
C487 B.n398 VSUBS 0.00667f
C488 B.n399 VSUBS 0.00667f
C489 B.n400 VSUBS 0.00667f
C490 B.n401 VSUBS 0.00667f
C491 B.n402 VSUBS 0.00667f
C492 B.n403 VSUBS 0.00667f
C493 B.n404 VSUBS 0.00667f
C494 B.n405 VSUBS 0.00667f
C495 B.n406 VSUBS 0.00667f
C496 B.n407 VSUBS 0.00667f
C497 B.n408 VSUBS 0.00667f
C498 B.n409 VSUBS 0.00667f
C499 B.n410 VSUBS 0.00667f
C500 B.n411 VSUBS 0.00667f
C501 B.n412 VSUBS 0.00667f
C502 B.n413 VSUBS 0.00667f
C503 B.n414 VSUBS 0.00667f
C504 B.n415 VSUBS 0.00667f
C505 B.n416 VSUBS 0.00667f
C506 B.n417 VSUBS 0.00667f
C507 B.n418 VSUBS 0.00667f
C508 B.n419 VSUBS 0.00667f
C509 B.n420 VSUBS 0.00667f
C510 B.n421 VSUBS 0.00667f
C511 B.n422 VSUBS 0.00667f
C512 B.n423 VSUBS 0.00667f
C513 B.n424 VSUBS 0.00667f
C514 B.n425 VSUBS 0.00667f
C515 B.n426 VSUBS 0.00667f
C516 B.n427 VSUBS 0.00667f
C517 B.n428 VSUBS 0.00667f
C518 B.n429 VSUBS 0.00667f
C519 B.n430 VSUBS 0.00667f
C520 B.n431 VSUBS 0.00667f
C521 B.n432 VSUBS 0.00667f
C522 B.n433 VSUBS 0.00667f
C523 B.n434 VSUBS 0.00667f
C524 B.n435 VSUBS 0.00667f
C525 B.n436 VSUBS 0.00667f
C526 B.n437 VSUBS 0.00667f
C527 B.n438 VSUBS 0.00667f
C528 B.n439 VSUBS 0.00667f
C529 B.n440 VSUBS 0.00667f
C530 B.n441 VSUBS 0.016072f
C531 B.n442 VSUBS 0.015275f
C532 B.n443 VSUBS 0.015722f
C533 B.n444 VSUBS 0.00667f
C534 B.n445 VSUBS 0.00667f
C535 B.n446 VSUBS 0.00667f
C536 B.n447 VSUBS 0.00667f
C537 B.n448 VSUBS 0.00667f
C538 B.n449 VSUBS 0.00667f
C539 B.n450 VSUBS 0.00667f
C540 B.n451 VSUBS 0.00667f
C541 B.n452 VSUBS 0.00667f
C542 B.n453 VSUBS 0.00667f
C543 B.n454 VSUBS 0.00667f
C544 B.n455 VSUBS 0.00667f
C545 B.n456 VSUBS 0.00667f
C546 B.n457 VSUBS 0.00667f
C547 B.n458 VSUBS 0.00667f
C548 B.n459 VSUBS 0.00667f
C549 B.n460 VSUBS 0.00667f
C550 B.n461 VSUBS 0.00667f
C551 B.n462 VSUBS 0.00667f
C552 B.n463 VSUBS 0.00667f
C553 B.n464 VSUBS 0.00667f
C554 B.n465 VSUBS 0.00667f
C555 B.n466 VSUBS 0.00667f
C556 B.n467 VSUBS 0.00667f
C557 B.n468 VSUBS 0.00667f
C558 B.n469 VSUBS 0.00667f
C559 B.n470 VSUBS 0.00667f
C560 B.n471 VSUBS 0.00667f
C561 B.n472 VSUBS 0.00667f
C562 B.n473 VSUBS 0.00667f
C563 B.n474 VSUBS 0.00667f
C564 B.n475 VSUBS 0.00667f
C565 B.n476 VSUBS 0.00667f
C566 B.n477 VSUBS 0.00667f
C567 B.n478 VSUBS 0.00667f
C568 B.n479 VSUBS 0.00667f
C569 B.n480 VSUBS 0.00667f
C570 B.n481 VSUBS 0.00667f
C571 B.n482 VSUBS 0.00667f
C572 B.n483 VSUBS 0.00667f
C573 B.n484 VSUBS 0.00667f
C574 B.n485 VSUBS 0.00667f
C575 B.n486 VSUBS 0.00667f
C576 B.n487 VSUBS 0.00667f
C577 B.n488 VSUBS 0.00667f
C578 B.n489 VSUBS 0.00667f
C579 B.n490 VSUBS 0.00667f
C580 B.n491 VSUBS 0.00667f
C581 B.n492 VSUBS 0.00667f
C582 B.n493 VSUBS 0.00667f
C583 B.n494 VSUBS 0.00667f
C584 B.n495 VSUBS 0.00667f
C585 B.n496 VSUBS 0.00667f
C586 B.n497 VSUBS 0.00667f
C587 B.n498 VSUBS 0.00667f
C588 B.n499 VSUBS 0.00667f
C589 B.n500 VSUBS 0.00667f
C590 B.n501 VSUBS 0.00667f
C591 B.n502 VSUBS 0.00667f
C592 B.n503 VSUBS 0.00667f
C593 B.n504 VSUBS 0.00667f
C594 B.n505 VSUBS 0.006278f
C595 B.n506 VSUBS 0.015454f
C596 B.n507 VSUBS 0.003728f
C597 B.n508 VSUBS 0.00667f
C598 B.n509 VSUBS 0.00667f
C599 B.n510 VSUBS 0.00667f
C600 B.n511 VSUBS 0.00667f
C601 B.n512 VSUBS 0.00667f
C602 B.n513 VSUBS 0.00667f
C603 B.n514 VSUBS 0.00667f
C604 B.n515 VSUBS 0.00667f
C605 B.n516 VSUBS 0.00667f
C606 B.n517 VSUBS 0.00667f
C607 B.n518 VSUBS 0.00667f
C608 B.n519 VSUBS 0.00667f
C609 B.n520 VSUBS 0.003728f
C610 B.n521 VSUBS 0.00667f
C611 B.n522 VSUBS 0.00667f
C612 B.n523 VSUBS 0.006278f
C613 B.n524 VSUBS 0.00667f
C614 B.n525 VSUBS 0.00667f
C615 B.n526 VSUBS 0.00667f
C616 B.n527 VSUBS 0.00667f
C617 B.n528 VSUBS 0.00667f
C618 B.n529 VSUBS 0.00667f
C619 B.n530 VSUBS 0.00667f
C620 B.n531 VSUBS 0.00667f
C621 B.n532 VSUBS 0.00667f
C622 B.n533 VSUBS 0.00667f
C623 B.n534 VSUBS 0.00667f
C624 B.n535 VSUBS 0.00667f
C625 B.n536 VSUBS 0.00667f
C626 B.n537 VSUBS 0.00667f
C627 B.n538 VSUBS 0.00667f
C628 B.n539 VSUBS 0.00667f
C629 B.n540 VSUBS 0.00667f
C630 B.n541 VSUBS 0.00667f
C631 B.n542 VSUBS 0.00667f
C632 B.n543 VSUBS 0.00667f
C633 B.n544 VSUBS 0.00667f
C634 B.n545 VSUBS 0.00667f
C635 B.n546 VSUBS 0.00667f
C636 B.n547 VSUBS 0.00667f
C637 B.n548 VSUBS 0.00667f
C638 B.n549 VSUBS 0.00667f
C639 B.n550 VSUBS 0.00667f
C640 B.n551 VSUBS 0.00667f
C641 B.n552 VSUBS 0.00667f
C642 B.n553 VSUBS 0.00667f
C643 B.n554 VSUBS 0.00667f
C644 B.n555 VSUBS 0.00667f
C645 B.n556 VSUBS 0.00667f
C646 B.n557 VSUBS 0.00667f
C647 B.n558 VSUBS 0.00667f
C648 B.n559 VSUBS 0.00667f
C649 B.n560 VSUBS 0.00667f
C650 B.n561 VSUBS 0.00667f
C651 B.n562 VSUBS 0.00667f
C652 B.n563 VSUBS 0.00667f
C653 B.n564 VSUBS 0.00667f
C654 B.n565 VSUBS 0.00667f
C655 B.n566 VSUBS 0.00667f
C656 B.n567 VSUBS 0.00667f
C657 B.n568 VSUBS 0.00667f
C658 B.n569 VSUBS 0.00667f
C659 B.n570 VSUBS 0.00667f
C660 B.n571 VSUBS 0.00667f
C661 B.n572 VSUBS 0.00667f
C662 B.n573 VSUBS 0.00667f
C663 B.n574 VSUBS 0.00667f
C664 B.n575 VSUBS 0.00667f
C665 B.n576 VSUBS 0.00667f
C666 B.n577 VSUBS 0.00667f
C667 B.n578 VSUBS 0.00667f
C668 B.n579 VSUBS 0.00667f
C669 B.n580 VSUBS 0.00667f
C670 B.n581 VSUBS 0.00667f
C671 B.n582 VSUBS 0.00667f
C672 B.n583 VSUBS 0.00667f
C673 B.n584 VSUBS 0.015722f
C674 B.n585 VSUBS 0.015275f
C675 B.n586 VSUBS 0.015275f
C676 B.n587 VSUBS 0.00667f
C677 B.n588 VSUBS 0.00667f
C678 B.n589 VSUBS 0.00667f
C679 B.n590 VSUBS 0.00667f
C680 B.n591 VSUBS 0.00667f
C681 B.n592 VSUBS 0.00667f
C682 B.n593 VSUBS 0.00667f
C683 B.n594 VSUBS 0.00667f
C684 B.n595 VSUBS 0.00667f
C685 B.n596 VSUBS 0.00667f
C686 B.n597 VSUBS 0.00667f
C687 B.n598 VSUBS 0.00667f
C688 B.n599 VSUBS 0.00667f
C689 B.n600 VSUBS 0.00667f
C690 B.n601 VSUBS 0.00667f
C691 B.n602 VSUBS 0.00667f
C692 B.n603 VSUBS 0.00667f
C693 B.n604 VSUBS 0.00667f
C694 B.n605 VSUBS 0.00667f
C695 B.n606 VSUBS 0.00667f
C696 B.n607 VSUBS 0.00667f
C697 B.n608 VSUBS 0.00667f
C698 B.n609 VSUBS 0.00667f
C699 B.n610 VSUBS 0.00667f
C700 B.n611 VSUBS 0.00667f
C701 B.n612 VSUBS 0.00667f
C702 B.n613 VSUBS 0.00667f
C703 B.n614 VSUBS 0.00667f
C704 B.n615 VSUBS 0.00667f
C705 B.n616 VSUBS 0.00667f
C706 B.n617 VSUBS 0.00667f
C707 B.n618 VSUBS 0.00667f
C708 B.n619 VSUBS 0.00667f
C709 B.n620 VSUBS 0.00667f
C710 B.n621 VSUBS 0.00667f
C711 B.n622 VSUBS 0.00667f
C712 B.n623 VSUBS 0.00667f
C713 B.n624 VSUBS 0.00667f
C714 B.n625 VSUBS 0.00667f
C715 B.n626 VSUBS 0.00667f
C716 B.n627 VSUBS 0.00667f
C717 B.n628 VSUBS 0.00667f
C718 B.n629 VSUBS 0.00667f
C719 B.n630 VSUBS 0.00667f
C720 B.n631 VSUBS 0.015104f
C721 VTAIL.t10 VSUBS 0.273203f
C722 VTAIL.t8 VSUBS 0.273203f
C723 VTAIL.n0 VSUBS 2.01554f
C724 VTAIL.n1 VSUBS 0.774431f
C725 VTAIL.t4 VSUBS 2.65293f
C726 VTAIL.n2 VSUBS 0.985707f
C727 VTAIL.t0 VSUBS 0.273203f
C728 VTAIL.t3 VSUBS 0.273203f
C729 VTAIL.n3 VSUBS 2.01554f
C730 VTAIL.n4 VSUBS 2.397f
C731 VTAIL.t9 VSUBS 0.273203f
C732 VTAIL.t11 VSUBS 0.273203f
C733 VTAIL.n5 VSUBS 2.01555f
C734 VTAIL.n6 VSUBS 2.39699f
C735 VTAIL.t7 VSUBS 2.65293f
C736 VTAIL.n7 VSUBS 0.985703f
C737 VTAIL.t5 VSUBS 0.273203f
C738 VTAIL.t2 VSUBS 0.273203f
C739 VTAIL.n8 VSUBS 2.01555f
C740 VTAIL.n9 VSUBS 0.877989f
C741 VTAIL.t1 VSUBS 2.65292f
C742 VTAIL.n10 VSUBS 2.35956f
C743 VTAIL.t6 VSUBS 2.65293f
C744 VTAIL.n11 VSUBS 2.31797f
C745 VDD2.t1 VSUBS 2.48967f
C746 VDD2.t5 VSUBS 0.24074f
C747 VDD2.t4 VSUBS 0.24074f
C748 VDD2.n0 VSUBS 1.90574f
C749 VDD2.n1 VSUBS 2.9463f
C750 VDD2.t3 VSUBS 2.48056f
C751 VDD2.n2 VSUBS 2.76761f
C752 VDD2.t0 VSUBS 0.24074f
C753 VDD2.t2 VSUBS 0.24074f
C754 VDD2.n3 VSUBS 1.9057f
C755 VN.n0 VSUBS 0.039959f
C756 VN.t5 VSUBS 2.0267f
C757 VN.n1 VSUBS 0.050176f
C758 VN.t1 VSUBS 2.1485f
C759 VN.n2 VSUBS 0.831891f
C760 VN.t3 VSUBS 2.0267f
C761 VN.n3 VSUBS 0.806811f
C762 VN.n4 VSUBS 0.056369f
C763 VN.n5 VSUBS 0.250076f
C764 VN.n6 VSUBS 0.039959f
C765 VN.n7 VSUBS 0.039959f
C766 VN.n8 VSUBS 0.066997f
C767 VN.n9 VSUBS 0.045283f
C768 VN.n10 VSUBS 0.80613f
C769 VN.n11 VSUBS 0.039985f
C770 VN.n12 VSUBS 0.039959f
C771 VN.t2 VSUBS 2.0267f
C772 VN.n13 VSUBS 0.050176f
C773 VN.t4 VSUBS 2.1485f
C774 VN.n14 VSUBS 0.831891f
C775 VN.t0 VSUBS 2.0267f
C776 VN.n15 VSUBS 0.806811f
C777 VN.n16 VSUBS 0.056369f
C778 VN.n17 VSUBS 0.250076f
C779 VN.n18 VSUBS 0.039959f
C780 VN.n19 VSUBS 0.039959f
C781 VN.n20 VSUBS 0.066997f
C782 VN.n21 VSUBS 0.045283f
C783 VN.n22 VSUBS 0.80613f
C784 VN.n23 VSUBS 1.84645f
.ends

