* NGSPICE file created from diff_pair_sample_0230.ext - technology: sky130A

.subckt diff_pair_sample_0230 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=1.9383 ps=10.72 w=4.97 l=2.15
X1 VTAIL.t3 VP.t0 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=0.82005 ps=5.3 w=4.97 l=2.15
X2 VDD1.t4 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=1.9383 ps=10.72 w=4.97 l=2.15
X3 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=1.9383 ps=10.72 w=4.97 l=2.15
X4 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0 ps=0 w=4.97 l=2.15
X5 VTAIL.t9 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=0.82005 ps=5.3 w=4.97 l=2.15
X6 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=0.82005 ps=5.3 w=4.97 l=2.15
X7 VDD2.t3 VN.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0.82005 ps=5.3 w=4.97 l=2.15
X8 VDD2.t2 VN.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0.82005 ps=5.3 w=4.97 l=2.15
X9 VTAIL.t6 VN.t4 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=0.82005 ps=5.3 w=4.97 l=2.15
X10 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0.82005 ps=5.3 w=4.97 l=2.15
X11 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0 ps=0 w=4.97 l=2.15
X12 VDD2.t0 VN.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.82005 pd=5.3 as=1.9383 ps=10.72 w=4.97 l=2.15
X13 VDD1.t0 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0.82005 ps=5.3 w=4.97 l=2.15
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0 ps=0 w=4.97 l=2.15
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9383 pd=10.72 as=0 ps=0 w=4.97 l=2.15
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n2 VN.t2 90.3655
R9 VN.n14 VN.t5 90.3655
R10 VN.n11 VN.n10 87.2681
R11 VN.n23 VN.n22 87.2681
R12 VN.n8 VN.n1 56.5193
R13 VN.n20 VN.n13 56.5193
R14 VN.n3 VN.t1 55.7107
R15 VN.n10 VN.t0 55.7107
R16 VN.n15 VN.t4 55.7107
R17 VN.n22 VN.t3 55.7107
R18 VN.n15 VN.n14 46.3955
R19 VN.n3 VN.n2 46.3955
R20 VN VN.n23 41.983
R21 VN.n4 VN.n3 24.4675
R22 VN.n4 VN.n1 24.4675
R23 VN.n9 VN.n8 24.4675
R24 VN.n16 VN.n13 24.4675
R25 VN.n16 VN.n15 24.4675
R26 VN.n21 VN.n20 24.4675
R27 VN.n10 VN.n9 23.4888
R28 VN.n22 VN.n21 23.4888
R29 VN.n17 VN.n14 8.64485
R30 VN.n5 VN.n2 8.64485
R31 VN.n23 VN.n12 0.278367
R32 VN.n11 VN.n0 0.278367
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153454
R40 VTAIL.n7 VTAIL.t10 57.8418
R41 VTAIL.n11 VTAIL.t8 57.8417
R42 VTAIL.n2 VTAIL.t2 57.8417
R43 VTAIL.n10 VTAIL.t5 57.8417
R44 VTAIL.n9 VTAIL.n8 53.858
R45 VTAIL.n6 VTAIL.n5 53.858
R46 VTAIL.n1 VTAIL.n0 53.8578
R47 VTAIL.n4 VTAIL.n3 53.8578
R48 VTAIL.n6 VTAIL.n4 20.9272
R49 VTAIL.n11 VTAIL.n10 18.7893
R50 VTAIL.n0 VTAIL.t7 3.9844
R51 VTAIL.n0 VTAIL.t9 3.9844
R52 VTAIL.n3 VTAIL.t4 3.9844
R53 VTAIL.n3 VTAIL.t3 3.9844
R54 VTAIL.n8 VTAIL.t0 3.9844
R55 VTAIL.n8 VTAIL.t1 3.9844
R56 VTAIL.n5 VTAIL.t11 3.9844
R57 VTAIL.n5 VTAIL.t6 3.9844
R58 VTAIL.n7 VTAIL.n6 2.13843
R59 VTAIL.n10 VTAIL.n9 2.13843
R60 VTAIL.n4 VTAIL.n2 2.13843
R61 VTAIL VTAIL.n11 1.54576
R62 VTAIL.n9 VTAIL.n7 1.53929
R63 VTAIL.n2 VTAIL.n1 1.53929
R64 VTAIL VTAIL.n1 0.593172
R65 VDD2.n1 VDD2.t3 76.0686
R66 VDD2.n2 VDD2.t2 74.5206
R67 VDD2.n1 VDD2.n0 71.0157
R68 VDD2 VDD2.n3 71.0129
R69 VDD2.n2 VDD2.n1 34.9481
R70 VDD2.n3 VDD2.t1 3.9844
R71 VDD2.n3 VDD2.t0 3.9844
R72 VDD2.n0 VDD2.t4 3.9844
R73 VDD2.n0 VDD2.t5 3.9844
R74 VDD2 VDD2.n2 1.66214
R75 B.n568 B.n567 585
R76 B.n569 B.n568 585
R77 B.n201 B.n96 585
R78 B.n200 B.n199 585
R79 B.n198 B.n197 585
R80 B.n196 B.n195 585
R81 B.n194 B.n193 585
R82 B.n192 B.n191 585
R83 B.n190 B.n189 585
R84 B.n188 B.n187 585
R85 B.n186 B.n185 585
R86 B.n184 B.n183 585
R87 B.n182 B.n181 585
R88 B.n180 B.n179 585
R89 B.n178 B.n177 585
R90 B.n176 B.n175 585
R91 B.n174 B.n173 585
R92 B.n172 B.n171 585
R93 B.n170 B.n169 585
R94 B.n168 B.n167 585
R95 B.n166 B.n165 585
R96 B.n164 B.n163 585
R97 B.n162 B.n161 585
R98 B.n160 B.n159 585
R99 B.n158 B.n157 585
R100 B.n156 B.n155 585
R101 B.n154 B.n153 585
R102 B.n152 B.n151 585
R103 B.n150 B.n149 585
R104 B.n148 B.n147 585
R105 B.n146 B.n145 585
R106 B.n143 B.n142 585
R107 B.n141 B.n140 585
R108 B.n139 B.n138 585
R109 B.n137 B.n136 585
R110 B.n135 B.n134 585
R111 B.n133 B.n132 585
R112 B.n131 B.n130 585
R113 B.n129 B.n128 585
R114 B.n127 B.n126 585
R115 B.n125 B.n124 585
R116 B.n123 B.n122 585
R117 B.n121 B.n120 585
R118 B.n119 B.n118 585
R119 B.n117 B.n116 585
R120 B.n115 B.n114 585
R121 B.n113 B.n112 585
R122 B.n111 B.n110 585
R123 B.n109 B.n108 585
R124 B.n107 B.n106 585
R125 B.n105 B.n104 585
R126 B.n103 B.n102 585
R127 B.n566 B.n70 585
R128 B.n570 B.n70 585
R129 B.n565 B.n69 585
R130 B.n571 B.n69 585
R131 B.n564 B.n563 585
R132 B.n563 B.n65 585
R133 B.n562 B.n64 585
R134 B.n577 B.n64 585
R135 B.n561 B.n63 585
R136 B.n578 B.n63 585
R137 B.n560 B.n62 585
R138 B.n579 B.n62 585
R139 B.n559 B.n558 585
R140 B.n558 B.n58 585
R141 B.n557 B.n57 585
R142 B.n585 B.n57 585
R143 B.n556 B.n56 585
R144 B.n586 B.n56 585
R145 B.n555 B.n55 585
R146 B.n587 B.n55 585
R147 B.n554 B.n553 585
R148 B.n553 B.n51 585
R149 B.n552 B.n50 585
R150 B.n593 B.n50 585
R151 B.n551 B.n49 585
R152 B.n594 B.n49 585
R153 B.n550 B.n48 585
R154 B.n595 B.n48 585
R155 B.n549 B.n548 585
R156 B.n548 B.n44 585
R157 B.n547 B.n43 585
R158 B.n601 B.n43 585
R159 B.n546 B.n42 585
R160 B.n602 B.n42 585
R161 B.n545 B.n41 585
R162 B.n603 B.n41 585
R163 B.n544 B.n543 585
R164 B.n543 B.n37 585
R165 B.n542 B.n36 585
R166 B.n609 B.n36 585
R167 B.n541 B.n35 585
R168 B.n610 B.n35 585
R169 B.n540 B.n34 585
R170 B.n611 B.n34 585
R171 B.n539 B.n538 585
R172 B.n538 B.n30 585
R173 B.n537 B.n29 585
R174 B.n617 B.n29 585
R175 B.n536 B.n28 585
R176 B.n618 B.n28 585
R177 B.n535 B.n27 585
R178 B.n619 B.n27 585
R179 B.n534 B.n533 585
R180 B.n533 B.n23 585
R181 B.n532 B.n22 585
R182 B.n625 B.n22 585
R183 B.n531 B.n21 585
R184 B.n626 B.n21 585
R185 B.n530 B.n20 585
R186 B.n627 B.n20 585
R187 B.n529 B.n528 585
R188 B.n528 B.n16 585
R189 B.n527 B.n15 585
R190 B.n633 B.n15 585
R191 B.n526 B.n14 585
R192 B.n634 B.n14 585
R193 B.n525 B.n13 585
R194 B.n635 B.n13 585
R195 B.n524 B.n523 585
R196 B.n523 B.n12 585
R197 B.n522 B.n521 585
R198 B.n522 B.n8 585
R199 B.n520 B.n7 585
R200 B.n642 B.n7 585
R201 B.n519 B.n6 585
R202 B.n643 B.n6 585
R203 B.n518 B.n5 585
R204 B.n644 B.n5 585
R205 B.n517 B.n516 585
R206 B.n516 B.n4 585
R207 B.n515 B.n202 585
R208 B.n515 B.n514 585
R209 B.n505 B.n203 585
R210 B.n204 B.n203 585
R211 B.n507 B.n506 585
R212 B.n508 B.n507 585
R213 B.n504 B.n208 585
R214 B.n212 B.n208 585
R215 B.n503 B.n502 585
R216 B.n502 B.n501 585
R217 B.n210 B.n209 585
R218 B.n211 B.n210 585
R219 B.n494 B.n493 585
R220 B.n495 B.n494 585
R221 B.n492 B.n217 585
R222 B.n217 B.n216 585
R223 B.n491 B.n490 585
R224 B.n490 B.n489 585
R225 B.n219 B.n218 585
R226 B.n220 B.n219 585
R227 B.n482 B.n481 585
R228 B.n483 B.n482 585
R229 B.n480 B.n224 585
R230 B.n228 B.n224 585
R231 B.n479 B.n478 585
R232 B.n478 B.n477 585
R233 B.n226 B.n225 585
R234 B.n227 B.n226 585
R235 B.n470 B.n469 585
R236 B.n471 B.n470 585
R237 B.n468 B.n233 585
R238 B.n233 B.n232 585
R239 B.n467 B.n466 585
R240 B.n466 B.n465 585
R241 B.n235 B.n234 585
R242 B.n236 B.n235 585
R243 B.n458 B.n457 585
R244 B.n459 B.n458 585
R245 B.n456 B.n241 585
R246 B.n241 B.n240 585
R247 B.n455 B.n454 585
R248 B.n454 B.n453 585
R249 B.n243 B.n242 585
R250 B.n244 B.n243 585
R251 B.n446 B.n445 585
R252 B.n447 B.n446 585
R253 B.n444 B.n249 585
R254 B.n249 B.n248 585
R255 B.n443 B.n442 585
R256 B.n442 B.n441 585
R257 B.n251 B.n250 585
R258 B.n252 B.n251 585
R259 B.n434 B.n433 585
R260 B.n435 B.n434 585
R261 B.n432 B.n257 585
R262 B.n257 B.n256 585
R263 B.n431 B.n430 585
R264 B.n430 B.n429 585
R265 B.n259 B.n258 585
R266 B.n260 B.n259 585
R267 B.n422 B.n421 585
R268 B.n423 B.n422 585
R269 B.n420 B.n265 585
R270 B.n265 B.n264 585
R271 B.n419 B.n418 585
R272 B.n418 B.n417 585
R273 B.n267 B.n266 585
R274 B.n268 B.n267 585
R275 B.n410 B.n409 585
R276 B.n411 B.n410 585
R277 B.n408 B.n273 585
R278 B.n273 B.n272 585
R279 B.n402 B.n401 585
R280 B.n400 B.n300 585
R281 B.n399 B.n299 585
R282 B.n404 B.n299 585
R283 B.n398 B.n397 585
R284 B.n396 B.n395 585
R285 B.n394 B.n393 585
R286 B.n392 B.n391 585
R287 B.n390 B.n389 585
R288 B.n388 B.n387 585
R289 B.n386 B.n385 585
R290 B.n384 B.n383 585
R291 B.n382 B.n381 585
R292 B.n380 B.n379 585
R293 B.n378 B.n377 585
R294 B.n376 B.n375 585
R295 B.n374 B.n373 585
R296 B.n372 B.n371 585
R297 B.n370 B.n369 585
R298 B.n368 B.n367 585
R299 B.n366 B.n365 585
R300 B.n364 B.n363 585
R301 B.n362 B.n361 585
R302 B.n360 B.n359 585
R303 B.n358 B.n357 585
R304 B.n356 B.n355 585
R305 B.n354 B.n353 585
R306 B.n352 B.n351 585
R307 B.n350 B.n349 585
R308 B.n348 B.n347 585
R309 B.n346 B.n345 585
R310 B.n343 B.n342 585
R311 B.n341 B.n340 585
R312 B.n339 B.n338 585
R313 B.n337 B.n336 585
R314 B.n335 B.n334 585
R315 B.n333 B.n332 585
R316 B.n331 B.n330 585
R317 B.n329 B.n328 585
R318 B.n327 B.n326 585
R319 B.n325 B.n324 585
R320 B.n323 B.n322 585
R321 B.n321 B.n320 585
R322 B.n319 B.n318 585
R323 B.n317 B.n316 585
R324 B.n315 B.n314 585
R325 B.n313 B.n312 585
R326 B.n311 B.n310 585
R327 B.n309 B.n308 585
R328 B.n307 B.n306 585
R329 B.n275 B.n274 585
R330 B.n407 B.n406 585
R331 B.n271 B.n270 585
R332 B.n272 B.n271 585
R333 B.n413 B.n412 585
R334 B.n412 B.n411 585
R335 B.n414 B.n269 585
R336 B.n269 B.n268 585
R337 B.n416 B.n415 585
R338 B.n417 B.n416 585
R339 B.n263 B.n262 585
R340 B.n264 B.n263 585
R341 B.n425 B.n424 585
R342 B.n424 B.n423 585
R343 B.n426 B.n261 585
R344 B.n261 B.n260 585
R345 B.n428 B.n427 585
R346 B.n429 B.n428 585
R347 B.n255 B.n254 585
R348 B.n256 B.n255 585
R349 B.n437 B.n436 585
R350 B.n436 B.n435 585
R351 B.n438 B.n253 585
R352 B.n253 B.n252 585
R353 B.n440 B.n439 585
R354 B.n441 B.n440 585
R355 B.n247 B.n246 585
R356 B.n248 B.n247 585
R357 B.n449 B.n448 585
R358 B.n448 B.n447 585
R359 B.n450 B.n245 585
R360 B.n245 B.n244 585
R361 B.n452 B.n451 585
R362 B.n453 B.n452 585
R363 B.n239 B.n238 585
R364 B.n240 B.n239 585
R365 B.n461 B.n460 585
R366 B.n460 B.n459 585
R367 B.n462 B.n237 585
R368 B.n237 B.n236 585
R369 B.n464 B.n463 585
R370 B.n465 B.n464 585
R371 B.n231 B.n230 585
R372 B.n232 B.n231 585
R373 B.n473 B.n472 585
R374 B.n472 B.n471 585
R375 B.n474 B.n229 585
R376 B.n229 B.n227 585
R377 B.n476 B.n475 585
R378 B.n477 B.n476 585
R379 B.n223 B.n222 585
R380 B.n228 B.n223 585
R381 B.n485 B.n484 585
R382 B.n484 B.n483 585
R383 B.n486 B.n221 585
R384 B.n221 B.n220 585
R385 B.n488 B.n487 585
R386 B.n489 B.n488 585
R387 B.n215 B.n214 585
R388 B.n216 B.n215 585
R389 B.n497 B.n496 585
R390 B.n496 B.n495 585
R391 B.n498 B.n213 585
R392 B.n213 B.n211 585
R393 B.n500 B.n499 585
R394 B.n501 B.n500 585
R395 B.n207 B.n206 585
R396 B.n212 B.n207 585
R397 B.n510 B.n509 585
R398 B.n509 B.n508 585
R399 B.n511 B.n205 585
R400 B.n205 B.n204 585
R401 B.n513 B.n512 585
R402 B.n514 B.n513 585
R403 B.n3 B.n0 585
R404 B.n4 B.n3 585
R405 B.n641 B.n1 585
R406 B.n642 B.n641 585
R407 B.n640 B.n639 585
R408 B.n640 B.n8 585
R409 B.n638 B.n9 585
R410 B.n12 B.n9 585
R411 B.n637 B.n636 585
R412 B.n636 B.n635 585
R413 B.n11 B.n10 585
R414 B.n634 B.n11 585
R415 B.n632 B.n631 585
R416 B.n633 B.n632 585
R417 B.n630 B.n17 585
R418 B.n17 B.n16 585
R419 B.n629 B.n628 585
R420 B.n628 B.n627 585
R421 B.n19 B.n18 585
R422 B.n626 B.n19 585
R423 B.n624 B.n623 585
R424 B.n625 B.n624 585
R425 B.n622 B.n24 585
R426 B.n24 B.n23 585
R427 B.n621 B.n620 585
R428 B.n620 B.n619 585
R429 B.n26 B.n25 585
R430 B.n618 B.n26 585
R431 B.n616 B.n615 585
R432 B.n617 B.n616 585
R433 B.n614 B.n31 585
R434 B.n31 B.n30 585
R435 B.n613 B.n612 585
R436 B.n612 B.n611 585
R437 B.n33 B.n32 585
R438 B.n610 B.n33 585
R439 B.n608 B.n607 585
R440 B.n609 B.n608 585
R441 B.n606 B.n38 585
R442 B.n38 B.n37 585
R443 B.n605 B.n604 585
R444 B.n604 B.n603 585
R445 B.n40 B.n39 585
R446 B.n602 B.n40 585
R447 B.n600 B.n599 585
R448 B.n601 B.n600 585
R449 B.n598 B.n45 585
R450 B.n45 B.n44 585
R451 B.n597 B.n596 585
R452 B.n596 B.n595 585
R453 B.n47 B.n46 585
R454 B.n594 B.n47 585
R455 B.n592 B.n591 585
R456 B.n593 B.n592 585
R457 B.n590 B.n52 585
R458 B.n52 B.n51 585
R459 B.n589 B.n588 585
R460 B.n588 B.n587 585
R461 B.n54 B.n53 585
R462 B.n586 B.n54 585
R463 B.n584 B.n583 585
R464 B.n585 B.n584 585
R465 B.n582 B.n59 585
R466 B.n59 B.n58 585
R467 B.n581 B.n580 585
R468 B.n580 B.n579 585
R469 B.n61 B.n60 585
R470 B.n578 B.n61 585
R471 B.n576 B.n575 585
R472 B.n577 B.n576 585
R473 B.n574 B.n66 585
R474 B.n66 B.n65 585
R475 B.n573 B.n572 585
R476 B.n572 B.n571 585
R477 B.n68 B.n67 585
R478 B.n570 B.n68 585
R479 B.n645 B.n644 585
R480 B.n643 B.n2 585
R481 B.n102 B.n68 502.111
R482 B.n568 B.n70 502.111
R483 B.n406 B.n273 502.111
R484 B.n402 B.n271 502.111
R485 B.n100 B.t17 262.959
R486 B.n97 B.t6 262.959
R487 B.n304 B.t14 262.959
R488 B.n301 B.t10 262.959
R489 B.n569 B.n95 256.663
R490 B.n569 B.n94 256.663
R491 B.n569 B.n93 256.663
R492 B.n569 B.n92 256.663
R493 B.n569 B.n91 256.663
R494 B.n569 B.n90 256.663
R495 B.n569 B.n89 256.663
R496 B.n569 B.n88 256.663
R497 B.n569 B.n87 256.663
R498 B.n569 B.n86 256.663
R499 B.n569 B.n85 256.663
R500 B.n569 B.n84 256.663
R501 B.n569 B.n83 256.663
R502 B.n569 B.n82 256.663
R503 B.n569 B.n81 256.663
R504 B.n569 B.n80 256.663
R505 B.n569 B.n79 256.663
R506 B.n569 B.n78 256.663
R507 B.n569 B.n77 256.663
R508 B.n569 B.n76 256.663
R509 B.n569 B.n75 256.663
R510 B.n569 B.n74 256.663
R511 B.n569 B.n73 256.663
R512 B.n569 B.n72 256.663
R513 B.n569 B.n71 256.663
R514 B.n404 B.n403 256.663
R515 B.n404 B.n276 256.663
R516 B.n404 B.n277 256.663
R517 B.n404 B.n278 256.663
R518 B.n404 B.n279 256.663
R519 B.n404 B.n280 256.663
R520 B.n404 B.n281 256.663
R521 B.n404 B.n282 256.663
R522 B.n404 B.n283 256.663
R523 B.n404 B.n284 256.663
R524 B.n404 B.n285 256.663
R525 B.n404 B.n286 256.663
R526 B.n404 B.n287 256.663
R527 B.n404 B.n288 256.663
R528 B.n404 B.n289 256.663
R529 B.n404 B.n290 256.663
R530 B.n404 B.n291 256.663
R531 B.n404 B.n292 256.663
R532 B.n404 B.n293 256.663
R533 B.n404 B.n294 256.663
R534 B.n404 B.n295 256.663
R535 B.n404 B.n296 256.663
R536 B.n404 B.n297 256.663
R537 B.n404 B.n298 256.663
R538 B.n405 B.n404 256.663
R539 B.n647 B.n646 256.663
R540 B.n106 B.n105 163.367
R541 B.n110 B.n109 163.367
R542 B.n114 B.n113 163.367
R543 B.n118 B.n117 163.367
R544 B.n122 B.n121 163.367
R545 B.n126 B.n125 163.367
R546 B.n130 B.n129 163.367
R547 B.n134 B.n133 163.367
R548 B.n138 B.n137 163.367
R549 B.n142 B.n141 163.367
R550 B.n147 B.n146 163.367
R551 B.n151 B.n150 163.367
R552 B.n155 B.n154 163.367
R553 B.n159 B.n158 163.367
R554 B.n163 B.n162 163.367
R555 B.n167 B.n166 163.367
R556 B.n171 B.n170 163.367
R557 B.n175 B.n174 163.367
R558 B.n179 B.n178 163.367
R559 B.n183 B.n182 163.367
R560 B.n187 B.n186 163.367
R561 B.n191 B.n190 163.367
R562 B.n195 B.n194 163.367
R563 B.n199 B.n198 163.367
R564 B.n568 B.n96 163.367
R565 B.n410 B.n273 163.367
R566 B.n410 B.n267 163.367
R567 B.n418 B.n267 163.367
R568 B.n418 B.n265 163.367
R569 B.n422 B.n265 163.367
R570 B.n422 B.n259 163.367
R571 B.n430 B.n259 163.367
R572 B.n430 B.n257 163.367
R573 B.n434 B.n257 163.367
R574 B.n434 B.n251 163.367
R575 B.n442 B.n251 163.367
R576 B.n442 B.n249 163.367
R577 B.n446 B.n249 163.367
R578 B.n446 B.n243 163.367
R579 B.n454 B.n243 163.367
R580 B.n454 B.n241 163.367
R581 B.n458 B.n241 163.367
R582 B.n458 B.n235 163.367
R583 B.n466 B.n235 163.367
R584 B.n466 B.n233 163.367
R585 B.n470 B.n233 163.367
R586 B.n470 B.n226 163.367
R587 B.n478 B.n226 163.367
R588 B.n478 B.n224 163.367
R589 B.n482 B.n224 163.367
R590 B.n482 B.n219 163.367
R591 B.n490 B.n219 163.367
R592 B.n490 B.n217 163.367
R593 B.n494 B.n217 163.367
R594 B.n494 B.n210 163.367
R595 B.n502 B.n210 163.367
R596 B.n502 B.n208 163.367
R597 B.n507 B.n208 163.367
R598 B.n507 B.n203 163.367
R599 B.n515 B.n203 163.367
R600 B.n516 B.n515 163.367
R601 B.n516 B.n5 163.367
R602 B.n6 B.n5 163.367
R603 B.n7 B.n6 163.367
R604 B.n522 B.n7 163.367
R605 B.n523 B.n522 163.367
R606 B.n523 B.n13 163.367
R607 B.n14 B.n13 163.367
R608 B.n15 B.n14 163.367
R609 B.n528 B.n15 163.367
R610 B.n528 B.n20 163.367
R611 B.n21 B.n20 163.367
R612 B.n22 B.n21 163.367
R613 B.n533 B.n22 163.367
R614 B.n533 B.n27 163.367
R615 B.n28 B.n27 163.367
R616 B.n29 B.n28 163.367
R617 B.n538 B.n29 163.367
R618 B.n538 B.n34 163.367
R619 B.n35 B.n34 163.367
R620 B.n36 B.n35 163.367
R621 B.n543 B.n36 163.367
R622 B.n543 B.n41 163.367
R623 B.n42 B.n41 163.367
R624 B.n43 B.n42 163.367
R625 B.n548 B.n43 163.367
R626 B.n548 B.n48 163.367
R627 B.n49 B.n48 163.367
R628 B.n50 B.n49 163.367
R629 B.n553 B.n50 163.367
R630 B.n553 B.n55 163.367
R631 B.n56 B.n55 163.367
R632 B.n57 B.n56 163.367
R633 B.n558 B.n57 163.367
R634 B.n558 B.n62 163.367
R635 B.n63 B.n62 163.367
R636 B.n64 B.n63 163.367
R637 B.n563 B.n64 163.367
R638 B.n563 B.n69 163.367
R639 B.n70 B.n69 163.367
R640 B.n300 B.n299 163.367
R641 B.n397 B.n299 163.367
R642 B.n395 B.n394 163.367
R643 B.n391 B.n390 163.367
R644 B.n387 B.n386 163.367
R645 B.n383 B.n382 163.367
R646 B.n379 B.n378 163.367
R647 B.n375 B.n374 163.367
R648 B.n371 B.n370 163.367
R649 B.n367 B.n366 163.367
R650 B.n363 B.n362 163.367
R651 B.n359 B.n358 163.367
R652 B.n355 B.n354 163.367
R653 B.n351 B.n350 163.367
R654 B.n347 B.n346 163.367
R655 B.n342 B.n341 163.367
R656 B.n338 B.n337 163.367
R657 B.n334 B.n333 163.367
R658 B.n330 B.n329 163.367
R659 B.n326 B.n325 163.367
R660 B.n322 B.n321 163.367
R661 B.n318 B.n317 163.367
R662 B.n314 B.n313 163.367
R663 B.n310 B.n309 163.367
R664 B.n306 B.n275 163.367
R665 B.n412 B.n271 163.367
R666 B.n412 B.n269 163.367
R667 B.n416 B.n269 163.367
R668 B.n416 B.n263 163.367
R669 B.n424 B.n263 163.367
R670 B.n424 B.n261 163.367
R671 B.n428 B.n261 163.367
R672 B.n428 B.n255 163.367
R673 B.n436 B.n255 163.367
R674 B.n436 B.n253 163.367
R675 B.n440 B.n253 163.367
R676 B.n440 B.n247 163.367
R677 B.n448 B.n247 163.367
R678 B.n448 B.n245 163.367
R679 B.n452 B.n245 163.367
R680 B.n452 B.n239 163.367
R681 B.n460 B.n239 163.367
R682 B.n460 B.n237 163.367
R683 B.n464 B.n237 163.367
R684 B.n464 B.n231 163.367
R685 B.n472 B.n231 163.367
R686 B.n472 B.n229 163.367
R687 B.n476 B.n229 163.367
R688 B.n476 B.n223 163.367
R689 B.n484 B.n223 163.367
R690 B.n484 B.n221 163.367
R691 B.n488 B.n221 163.367
R692 B.n488 B.n215 163.367
R693 B.n496 B.n215 163.367
R694 B.n496 B.n213 163.367
R695 B.n500 B.n213 163.367
R696 B.n500 B.n207 163.367
R697 B.n509 B.n207 163.367
R698 B.n509 B.n205 163.367
R699 B.n513 B.n205 163.367
R700 B.n513 B.n3 163.367
R701 B.n645 B.n3 163.367
R702 B.n641 B.n2 163.367
R703 B.n641 B.n640 163.367
R704 B.n640 B.n9 163.367
R705 B.n636 B.n9 163.367
R706 B.n636 B.n11 163.367
R707 B.n632 B.n11 163.367
R708 B.n632 B.n17 163.367
R709 B.n628 B.n17 163.367
R710 B.n628 B.n19 163.367
R711 B.n624 B.n19 163.367
R712 B.n624 B.n24 163.367
R713 B.n620 B.n24 163.367
R714 B.n620 B.n26 163.367
R715 B.n616 B.n26 163.367
R716 B.n616 B.n31 163.367
R717 B.n612 B.n31 163.367
R718 B.n612 B.n33 163.367
R719 B.n608 B.n33 163.367
R720 B.n608 B.n38 163.367
R721 B.n604 B.n38 163.367
R722 B.n604 B.n40 163.367
R723 B.n600 B.n40 163.367
R724 B.n600 B.n45 163.367
R725 B.n596 B.n45 163.367
R726 B.n596 B.n47 163.367
R727 B.n592 B.n47 163.367
R728 B.n592 B.n52 163.367
R729 B.n588 B.n52 163.367
R730 B.n588 B.n54 163.367
R731 B.n584 B.n54 163.367
R732 B.n584 B.n59 163.367
R733 B.n580 B.n59 163.367
R734 B.n580 B.n61 163.367
R735 B.n576 B.n61 163.367
R736 B.n576 B.n66 163.367
R737 B.n572 B.n66 163.367
R738 B.n572 B.n68 163.367
R739 B.n97 B.t8 122.382
R740 B.n304 B.t16 122.382
R741 B.n100 B.t18 122.376
R742 B.n301 B.t13 122.376
R743 B.n404 B.n272 117.034
R744 B.n570 B.n569 117.034
R745 B.n98 B.t9 74.2845
R746 B.n305 B.t15 74.2845
R747 B.n101 B.t19 74.2797
R748 B.n302 B.t12 74.2797
R749 B.n411 B.n272 73.0117
R750 B.n411 B.n268 73.0117
R751 B.n417 B.n268 73.0117
R752 B.n417 B.n264 73.0117
R753 B.n423 B.n264 73.0117
R754 B.n423 B.n260 73.0117
R755 B.n429 B.n260 73.0117
R756 B.n435 B.n256 73.0117
R757 B.n435 B.n252 73.0117
R758 B.n441 B.n252 73.0117
R759 B.n441 B.n248 73.0117
R760 B.n447 B.n248 73.0117
R761 B.n447 B.n244 73.0117
R762 B.n453 B.n244 73.0117
R763 B.n453 B.n240 73.0117
R764 B.n459 B.n240 73.0117
R765 B.n465 B.n236 73.0117
R766 B.n465 B.n232 73.0117
R767 B.n471 B.n232 73.0117
R768 B.n471 B.n227 73.0117
R769 B.n477 B.n227 73.0117
R770 B.n477 B.n228 73.0117
R771 B.n483 B.n220 73.0117
R772 B.n489 B.n220 73.0117
R773 B.n489 B.n216 73.0117
R774 B.n495 B.n216 73.0117
R775 B.n495 B.n211 73.0117
R776 B.n501 B.n211 73.0117
R777 B.n501 B.n212 73.0117
R778 B.n508 B.n204 73.0117
R779 B.n514 B.n204 73.0117
R780 B.n514 B.n4 73.0117
R781 B.n644 B.n4 73.0117
R782 B.n644 B.n643 73.0117
R783 B.n643 B.n642 73.0117
R784 B.n642 B.n8 73.0117
R785 B.n12 B.n8 73.0117
R786 B.n635 B.n12 73.0117
R787 B.n634 B.n633 73.0117
R788 B.n633 B.n16 73.0117
R789 B.n627 B.n16 73.0117
R790 B.n627 B.n626 73.0117
R791 B.n626 B.n625 73.0117
R792 B.n625 B.n23 73.0117
R793 B.n619 B.n23 73.0117
R794 B.n618 B.n617 73.0117
R795 B.n617 B.n30 73.0117
R796 B.n611 B.n30 73.0117
R797 B.n611 B.n610 73.0117
R798 B.n610 B.n609 73.0117
R799 B.n609 B.n37 73.0117
R800 B.n603 B.n602 73.0117
R801 B.n602 B.n601 73.0117
R802 B.n601 B.n44 73.0117
R803 B.n595 B.n44 73.0117
R804 B.n595 B.n594 73.0117
R805 B.n594 B.n593 73.0117
R806 B.n593 B.n51 73.0117
R807 B.n587 B.n51 73.0117
R808 B.n587 B.n586 73.0117
R809 B.n585 B.n58 73.0117
R810 B.n579 B.n58 73.0117
R811 B.n579 B.n578 73.0117
R812 B.n578 B.n577 73.0117
R813 B.n577 B.n65 73.0117
R814 B.n571 B.n65 73.0117
R815 B.n571 B.n570 73.0117
R816 B.n102 B.n71 71.676
R817 B.n106 B.n72 71.676
R818 B.n110 B.n73 71.676
R819 B.n114 B.n74 71.676
R820 B.n118 B.n75 71.676
R821 B.n122 B.n76 71.676
R822 B.n126 B.n77 71.676
R823 B.n130 B.n78 71.676
R824 B.n134 B.n79 71.676
R825 B.n138 B.n80 71.676
R826 B.n142 B.n81 71.676
R827 B.n147 B.n82 71.676
R828 B.n151 B.n83 71.676
R829 B.n155 B.n84 71.676
R830 B.n159 B.n85 71.676
R831 B.n163 B.n86 71.676
R832 B.n167 B.n87 71.676
R833 B.n171 B.n88 71.676
R834 B.n175 B.n89 71.676
R835 B.n179 B.n90 71.676
R836 B.n183 B.n91 71.676
R837 B.n187 B.n92 71.676
R838 B.n191 B.n93 71.676
R839 B.n195 B.n94 71.676
R840 B.n199 B.n95 71.676
R841 B.n96 B.n95 71.676
R842 B.n198 B.n94 71.676
R843 B.n194 B.n93 71.676
R844 B.n190 B.n92 71.676
R845 B.n186 B.n91 71.676
R846 B.n182 B.n90 71.676
R847 B.n178 B.n89 71.676
R848 B.n174 B.n88 71.676
R849 B.n170 B.n87 71.676
R850 B.n166 B.n86 71.676
R851 B.n162 B.n85 71.676
R852 B.n158 B.n84 71.676
R853 B.n154 B.n83 71.676
R854 B.n150 B.n82 71.676
R855 B.n146 B.n81 71.676
R856 B.n141 B.n80 71.676
R857 B.n137 B.n79 71.676
R858 B.n133 B.n78 71.676
R859 B.n129 B.n77 71.676
R860 B.n125 B.n76 71.676
R861 B.n121 B.n75 71.676
R862 B.n117 B.n74 71.676
R863 B.n113 B.n73 71.676
R864 B.n109 B.n72 71.676
R865 B.n105 B.n71 71.676
R866 B.n403 B.n402 71.676
R867 B.n397 B.n276 71.676
R868 B.n394 B.n277 71.676
R869 B.n390 B.n278 71.676
R870 B.n386 B.n279 71.676
R871 B.n382 B.n280 71.676
R872 B.n378 B.n281 71.676
R873 B.n374 B.n282 71.676
R874 B.n370 B.n283 71.676
R875 B.n366 B.n284 71.676
R876 B.n362 B.n285 71.676
R877 B.n358 B.n286 71.676
R878 B.n354 B.n287 71.676
R879 B.n350 B.n288 71.676
R880 B.n346 B.n289 71.676
R881 B.n341 B.n290 71.676
R882 B.n337 B.n291 71.676
R883 B.n333 B.n292 71.676
R884 B.n329 B.n293 71.676
R885 B.n325 B.n294 71.676
R886 B.n321 B.n295 71.676
R887 B.n317 B.n296 71.676
R888 B.n313 B.n297 71.676
R889 B.n309 B.n298 71.676
R890 B.n405 B.n275 71.676
R891 B.n403 B.n300 71.676
R892 B.n395 B.n276 71.676
R893 B.n391 B.n277 71.676
R894 B.n387 B.n278 71.676
R895 B.n383 B.n279 71.676
R896 B.n379 B.n280 71.676
R897 B.n375 B.n281 71.676
R898 B.n371 B.n282 71.676
R899 B.n367 B.n283 71.676
R900 B.n363 B.n284 71.676
R901 B.n359 B.n285 71.676
R902 B.n355 B.n286 71.676
R903 B.n351 B.n287 71.676
R904 B.n347 B.n288 71.676
R905 B.n342 B.n289 71.676
R906 B.n338 B.n290 71.676
R907 B.n334 B.n291 71.676
R908 B.n330 B.n292 71.676
R909 B.n326 B.n293 71.676
R910 B.n322 B.n294 71.676
R911 B.n318 B.n295 71.676
R912 B.n314 B.n296 71.676
R913 B.n310 B.n297 71.676
R914 B.n306 B.n298 71.676
R915 B.n406 B.n405 71.676
R916 B.n646 B.n645 71.676
R917 B.n646 B.n2 71.676
R918 B.n228 B.t3 69.7906
R919 B.t1 B.n618 69.7906
R920 B.t11 B.n256 61.2011
R921 B.n586 B.t7 61.2011
R922 B.n144 B.n101 59.5399
R923 B.n99 B.n98 59.5399
R924 B.n344 B.n305 59.5399
R925 B.n303 B.n302 59.5399
R926 B.n508 B.t2 54.7589
R927 B.n635 B.t0 54.7589
R928 B.n459 B.t4 48.3167
R929 B.n603 B.t5 48.3167
R930 B.n101 B.n100 48.0975
R931 B.n98 B.n97 48.0975
R932 B.n305 B.n304 48.0975
R933 B.n302 B.n301 48.0975
R934 B.n401 B.n270 32.6249
R935 B.n408 B.n407 32.6249
R936 B.n567 B.n566 32.6249
R937 B.n103 B.n67 32.6249
R938 B.t4 B.n236 24.6955
R939 B.t5 B.n37 24.6955
R940 B.n212 B.t2 18.2533
R941 B.t0 B.n634 18.2533
R942 B B.n647 18.0485
R943 B.n429 B.t11 11.8111
R944 B.t7 B.n585 11.8111
R945 B.n413 B.n270 10.6151
R946 B.n414 B.n413 10.6151
R947 B.n415 B.n414 10.6151
R948 B.n415 B.n262 10.6151
R949 B.n425 B.n262 10.6151
R950 B.n426 B.n425 10.6151
R951 B.n427 B.n426 10.6151
R952 B.n427 B.n254 10.6151
R953 B.n437 B.n254 10.6151
R954 B.n438 B.n437 10.6151
R955 B.n439 B.n438 10.6151
R956 B.n439 B.n246 10.6151
R957 B.n449 B.n246 10.6151
R958 B.n450 B.n449 10.6151
R959 B.n451 B.n450 10.6151
R960 B.n451 B.n238 10.6151
R961 B.n461 B.n238 10.6151
R962 B.n462 B.n461 10.6151
R963 B.n463 B.n462 10.6151
R964 B.n463 B.n230 10.6151
R965 B.n473 B.n230 10.6151
R966 B.n474 B.n473 10.6151
R967 B.n475 B.n474 10.6151
R968 B.n475 B.n222 10.6151
R969 B.n485 B.n222 10.6151
R970 B.n486 B.n485 10.6151
R971 B.n487 B.n486 10.6151
R972 B.n487 B.n214 10.6151
R973 B.n497 B.n214 10.6151
R974 B.n498 B.n497 10.6151
R975 B.n499 B.n498 10.6151
R976 B.n499 B.n206 10.6151
R977 B.n510 B.n206 10.6151
R978 B.n511 B.n510 10.6151
R979 B.n512 B.n511 10.6151
R980 B.n512 B.n0 10.6151
R981 B.n401 B.n400 10.6151
R982 B.n400 B.n399 10.6151
R983 B.n399 B.n398 10.6151
R984 B.n398 B.n396 10.6151
R985 B.n396 B.n393 10.6151
R986 B.n393 B.n392 10.6151
R987 B.n392 B.n389 10.6151
R988 B.n389 B.n388 10.6151
R989 B.n388 B.n385 10.6151
R990 B.n385 B.n384 10.6151
R991 B.n384 B.n381 10.6151
R992 B.n381 B.n380 10.6151
R993 B.n380 B.n377 10.6151
R994 B.n377 B.n376 10.6151
R995 B.n376 B.n373 10.6151
R996 B.n373 B.n372 10.6151
R997 B.n372 B.n369 10.6151
R998 B.n369 B.n368 10.6151
R999 B.n368 B.n365 10.6151
R1000 B.n365 B.n364 10.6151
R1001 B.n361 B.n360 10.6151
R1002 B.n360 B.n357 10.6151
R1003 B.n357 B.n356 10.6151
R1004 B.n356 B.n353 10.6151
R1005 B.n353 B.n352 10.6151
R1006 B.n352 B.n349 10.6151
R1007 B.n349 B.n348 10.6151
R1008 B.n348 B.n345 10.6151
R1009 B.n343 B.n340 10.6151
R1010 B.n340 B.n339 10.6151
R1011 B.n339 B.n336 10.6151
R1012 B.n336 B.n335 10.6151
R1013 B.n335 B.n332 10.6151
R1014 B.n332 B.n331 10.6151
R1015 B.n331 B.n328 10.6151
R1016 B.n328 B.n327 10.6151
R1017 B.n327 B.n324 10.6151
R1018 B.n324 B.n323 10.6151
R1019 B.n323 B.n320 10.6151
R1020 B.n320 B.n319 10.6151
R1021 B.n319 B.n316 10.6151
R1022 B.n316 B.n315 10.6151
R1023 B.n315 B.n312 10.6151
R1024 B.n312 B.n311 10.6151
R1025 B.n311 B.n308 10.6151
R1026 B.n308 B.n307 10.6151
R1027 B.n307 B.n274 10.6151
R1028 B.n407 B.n274 10.6151
R1029 B.n409 B.n408 10.6151
R1030 B.n409 B.n266 10.6151
R1031 B.n419 B.n266 10.6151
R1032 B.n420 B.n419 10.6151
R1033 B.n421 B.n420 10.6151
R1034 B.n421 B.n258 10.6151
R1035 B.n431 B.n258 10.6151
R1036 B.n432 B.n431 10.6151
R1037 B.n433 B.n432 10.6151
R1038 B.n433 B.n250 10.6151
R1039 B.n443 B.n250 10.6151
R1040 B.n444 B.n443 10.6151
R1041 B.n445 B.n444 10.6151
R1042 B.n445 B.n242 10.6151
R1043 B.n455 B.n242 10.6151
R1044 B.n456 B.n455 10.6151
R1045 B.n457 B.n456 10.6151
R1046 B.n457 B.n234 10.6151
R1047 B.n467 B.n234 10.6151
R1048 B.n468 B.n467 10.6151
R1049 B.n469 B.n468 10.6151
R1050 B.n469 B.n225 10.6151
R1051 B.n479 B.n225 10.6151
R1052 B.n480 B.n479 10.6151
R1053 B.n481 B.n480 10.6151
R1054 B.n481 B.n218 10.6151
R1055 B.n491 B.n218 10.6151
R1056 B.n492 B.n491 10.6151
R1057 B.n493 B.n492 10.6151
R1058 B.n493 B.n209 10.6151
R1059 B.n503 B.n209 10.6151
R1060 B.n504 B.n503 10.6151
R1061 B.n506 B.n504 10.6151
R1062 B.n506 B.n505 10.6151
R1063 B.n505 B.n202 10.6151
R1064 B.n517 B.n202 10.6151
R1065 B.n518 B.n517 10.6151
R1066 B.n519 B.n518 10.6151
R1067 B.n520 B.n519 10.6151
R1068 B.n521 B.n520 10.6151
R1069 B.n524 B.n521 10.6151
R1070 B.n525 B.n524 10.6151
R1071 B.n526 B.n525 10.6151
R1072 B.n527 B.n526 10.6151
R1073 B.n529 B.n527 10.6151
R1074 B.n530 B.n529 10.6151
R1075 B.n531 B.n530 10.6151
R1076 B.n532 B.n531 10.6151
R1077 B.n534 B.n532 10.6151
R1078 B.n535 B.n534 10.6151
R1079 B.n536 B.n535 10.6151
R1080 B.n537 B.n536 10.6151
R1081 B.n539 B.n537 10.6151
R1082 B.n540 B.n539 10.6151
R1083 B.n541 B.n540 10.6151
R1084 B.n542 B.n541 10.6151
R1085 B.n544 B.n542 10.6151
R1086 B.n545 B.n544 10.6151
R1087 B.n546 B.n545 10.6151
R1088 B.n547 B.n546 10.6151
R1089 B.n549 B.n547 10.6151
R1090 B.n550 B.n549 10.6151
R1091 B.n551 B.n550 10.6151
R1092 B.n552 B.n551 10.6151
R1093 B.n554 B.n552 10.6151
R1094 B.n555 B.n554 10.6151
R1095 B.n556 B.n555 10.6151
R1096 B.n557 B.n556 10.6151
R1097 B.n559 B.n557 10.6151
R1098 B.n560 B.n559 10.6151
R1099 B.n561 B.n560 10.6151
R1100 B.n562 B.n561 10.6151
R1101 B.n564 B.n562 10.6151
R1102 B.n565 B.n564 10.6151
R1103 B.n566 B.n565 10.6151
R1104 B.n639 B.n1 10.6151
R1105 B.n639 B.n638 10.6151
R1106 B.n638 B.n637 10.6151
R1107 B.n637 B.n10 10.6151
R1108 B.n631 B.n10 10.6151
R1109 B.n631 B.n630 10.6151
R1110 B.n630 B.n629 10.6151
R1111 B.n629 B.n18 10.6151
R1112 B.n623 B.n18 10.6151
R1113 B.n623 B.n622 10.6151
R1114 B.n622 B.n621 10.6151
R1115 B.n621 B.n25 10.6151
R1116 B.n615 B.n25 10.6151
R1117 B.n615 B.n614 10.6151
R1118 B.n614 B.n613 10.6151
R1119 B.n613 B.n32 10.6151
R1120 B.n607 B.n32 10.6151
R1121 B.n607 B.n606 10.6151
R1122 B.n606 B.n605 10.6151
R1123 B.n605 B.n39 10.6151
R1124 B.n599 B.n39 10.6151
R1125 B.n599 B.n598 10.6151
R1126 B.n598 B.n597 10.6151
R1127 B.n597 B.n46 10.6151
R1128 B.n591 B.n46 10.6151
R1129 B.n591 B.n590 10.6151
R1130 B.n590 B.n589 10.6151
R1131 B.n589 B.n53 10.6151
R1132 B.n583 B.n53 10.6151
R1133 B.n583 B.n582 10.6151
R1134 B.n582 B.n581 10.6151
R1135 B.n581 B.n60 10.6151
R1136 B.n575 B.n60 10.6151
R1137 B.n575 B.n574 10.6151
R1138 B.n574 B.n573 10.6151
R1139 B.n573 B.n67 10.6151
R1140 B.n104 B.n103 10.6151
R1141 B.n107 B.n104 10.6151
R1142 B.n108 B.n107 10.6151
R1143 B.n111 B.n108 10.6151
R1144 B.n112 B.n111 10.6151
R1145 B.n115 B.n112 10.6151
R1146 B.n116 B.n115 10.6151
R1147 B.n119 B.n116 10.6151
R1148 B.n120 B.n119 10.6151
R1149 B.n123 B.n120 10.6151
R1150 B.n124 B.n123 10.6151
R1151 B.n127 B.n124 10.6151
R1152 B.n128 B.n127 10.6151
R1153 B.n131 B.n128 10.6151
R1154 B.n132 B.n131 10.6151
R1155 B.n135 B.n132 10.6151
R1156 B.n136 B.n135 10.6151
R1157 B.n139 B.n136 10.6151
R1158 B.n140 B.n139 10.6151
R1159 B.n143 B.n140 10.6151
R1160 B.n148 B.n145 10.6151
R1161 B.n149 B.n148 10.6151
R1162 B.n152 B.n149 10.6151
R1163 B.n153 B.n152 10.6151
R1164 B.n156 B.n153 10.6151
R1165 B.n157 B.n156 10.6151
R1166 B.n160 B.n157 10.6151
R1167 B.n161 B.n160 10.6151
R1168 B.n165 B.n164 10.6151
R1169 B.n168 B.n165 10.6151
R1170 B.n169 B.n168 10.6151
R1171 B.n172 B.n169 10.6151
R1172 B.n173 B.n172 10.6151
R1173 B.n176 B.n173 10.6151
R1174 B.n177 B.n176 10.6151
R1175 B.n180 B.n177 10.6151
R1176 B.n181 B.n180 10.6151
R1177 B.n184 B.n181 10.6151
R1178 B.n185 B.n184 10.6151
R1179 B.n188 B.n185 10.6151
R1180 B.n189 B.n188 10.6151
R1181 B.n192 B.n189 10.6151
R1182 B.n193 B.n192 10.6151
R1183 B.n196 B.n193 10.6151
R1184 B.n197 B.n196 10.6151
R1185 B.n200 B.n197 10.6151
R1186 B.n201 B.n200 10.6151
R1187 B.n567 B.n201 10.6151
R1188 B.n647 B.n0 8.11757
R1189 B.n647 B.n1 8.11757
R1190 B.n361 B.n303 6.5566
R1191 B.n345 B.n344 6.5566
R1192 B.n145 B.n144 6.5566
R1193 B.n161 B.n99 6.5566
R1194 B.n364 B.n303 4.05904
R1195 B.n344 B.n343 4.05904
R1196 B.n144 B.n143 4.05904
R1197 B.n164 B.n99 4.05904
R1198 B.n483 B.t3 3.22158
R1199 B.n619 B.t1 3.22158
R1200 VP.n10 VP.n9 161.3
R1201 VP.n11 VP.n6 161.3
R1202 VP.n13 VP.n12 161.3
R1203 VP.n14 VP.n5 161.3
R1204 VP.n31 VP.n0 161.3
R1205 VP.n30 VP.n29 161.3
R1206 VP.n28 VP.n1 161.3
R1207 VP.n27 VP.n26 161.3
R1208 VP.n25 VP.n2 161.3
R1209 VP.n24 VP.n23 161.3
R1210 VP.n22 VP.n3 161.3
R1211 VP.n21 VP.n20 161.3
R1212 VP.n19 VP.n4 161.3
R1213 VP.n7 VP.t4 90.3655
R1214 VP.n18 VP.n17 87.2681
R1215 VP.n33 VP.n32 87.2681
R1216 VP.n16 VP.n15 87.2681
R1217 VP.n20 VP.n3 56.5193
R1218 VP.n30 VP.n1 56.5193
R1219 VP.n13 VP.n6 56.5193
R1220 VP.n25 VP.t0 55.7107
R1221 VP.n18 VP.t5 55.7107
R1222 VP.n32 VP.t2 55.7107
R1223 VP.n8 VP.t3 55.7107
R1224 VP.n15 VP.t1 55.7107
R1225 VP.n8 VP.n7 46.3955
R1226 VP.n17 VP.n16 41.7041
R1227 VP.n20 VP.n19 24.4675
R1228 VP.n24 VP.n3 24.4675
R1229 VP.n25 VP.n24 24.4675
R1230 VP.n26 VP.n25 24.4675
R1231 VP.n26 VP.n1 24.4675
R1232 VP.n31 VP.n30 24.4675
R1233 VP.n14 VP.n13 24.4675
R1234 VP.n9 VP.n8 24.4675
R1235 VP.n9 VP.n6 24.4675
R1236 VP.n19 VP.n18 23.4888
R1237 VP.n32 VP.n31 23.4888
R1238 VP.n15 VP.n14 23.4888
R1239 VP.n10 VP.n7 8.64485
R1240 VP.n16 VP.n5 0.278367
R1241 VP.n17 VP.n4 0.278367
R1242 VP.n33 VP.n0 0.278367
R1243 VP.n11 VP.n10 0.189894
R1244 VP.n12 VP.n11 0.189894
R1245 VP.n12 VP.n5 0.189894
R1246 VP.n21 VP.n4 0.189894
R1247 VP.n22 VP.n21 0.189894
R1248 VP.n23 VP.n22 0.189894
R1249 VP.n23 VP.n2 0.189894
R1250 VP.n27 VP.n2 0.189894
R1251 VP.n28 VP.n27 0.189894
R1252 VP.n29 VP.n28 0.189894
R1253 VP.n29 VP.n0 0.189894
R1254 VP VP.n33 0.153454
R1255 VDD1 VDD1.t1 76.1822
R1256 VDD1.n1 VDD1.t0 76.0686
R1257 VDD1.n1 VDD1.n0 71.0157
R1258 VDD1.n3 VDD1.n2 70.5366
R1259 VDD1.n3 VDD1.n1 36.6
R1260 VDD1.n2 VDD1.t2 3.9844
R1261 VDD1.n2 VDD1.t4 3.9844
R1262 VDD1.n0 VDD1.t5 3.9844
R1263 VDD1.n0 VDD1.t3 3.9844
R1264 VDD1 VDD1.n3 0.476793
C0 VTAIL VP 3.40127f
C1 VN VDD2 2.89699f
C2 VN VTAIL 3.38708f
C3 VDD1 VDD2 1.23133f
C4 VN VP 5.18436f
C5 VDD1 VTAIL 4.958991f
C6 VDD1 VP 3.16443f
C7 VDD1 VN 0.150199f
C8 VTAIL VDD2 5.00821f
C9 VDD2 VP 0.423805f
C10 VDD2 B 4.386925f
C11 VDD1 B 4.690489f
C12 VTAIL B 4.457001f
C13 VN B 10.88833f
C14 VP B 9.520096f
C15 VDD1.t1 B 0.924612f
C16 VDD1.t0 B 0.923926f
C17 VDD1.t5 B 0.088698f
C18 VDD1.t3 B 0.088698f
C19 VDD1.n0 B 0.724268f
C20 VDD1.n1 B 2.14202f
C21 VDD1.t2 B 0.088698f
C22 VDD1.t4 B 0.088698f
C23 VDD1.n2 B 0.721701f
C24 VDD1.n3 B 1.90435f
C25 VP.n0 B 0.040538f
C26 VP.t2 B 0.859011f
C27 VP.n1 B 0.044029f
C28 VP.n2 B 0.030748f
C29 VP.t0 B 0.859011f
C30 VP.n3 B 0.044029f
C31 VP.n4 B 0.040538f
C32 VP.t5 B 0.859011f
C33 VP.n5 B 0.040538f
C34 VP.t1 B 0.859011f
C35 VP.n6 B 0.044029f
C36 VP.t4 B 1.0541f
C37 VP.n7 B 0.398475f
C38 VP.t3 B 0.859011f
C39 VP.n8 B 0.429143f
C40 VP.n9 B 0.057306f
C41 VP.n10 B 0.259505f
C42 VP.n11 B 0.030748f
C43 VP.n12 B 0.030748f
C44 VP.n13 B 0.045743f
C45 VP.n14 B 0.056174f
C46 VP.n15 B 0.443856f
C47 VP.n16 B 1.27836f
C48 VP.n17 B 1.30487f
C49 VP.n18 B 0.443856f
C50 VP.n19 B 0.056174f
C51 VP.n20 B 0.045743f
C52 VP.n21 B 0.030748f
C53 VP.n22 B 0.030748f
C54 VP.n23 B 0.030748f
C55 VP.n24 B 0.057306f
C56 VP.n25 B 0.364228f
C57 VP.n26 B 0.057306f
C58 VP.n27 B 0.030748f
C59 VP.n28 B 0.030748f
C60 VP.n29 B 0.030748f
C61 VP.n30 B 0.045743f
C62 VP.n31 B 0.056174f
C63 VP.n32 B 0.443856f
C64 VP.n33 B 0.0342f
C65 VDD2.t3 B 0.899272f
C66 VDD2.t4 B 0.086331f
C67 VDD2.t5 B 0.086331f
C68 VDD2.n0 B 0.704942f
C69 VDD2.n1 B 1.9913f
C70 VDD2.t2 B 0.892371f
C71 VDD2.n2 B 1.84396f
C72 VDD2.t1 B 0.086331f
C73 VDD2.t0 B 0.086331f
C74 VDD2.n3 B 0.704918f
C75 VTAIL.t7 B 0.108424f
C76 VTAIL.t9 B 0.108424f
C77 VTAIL.n0 B 0.815794f
C78 VTAIL.n1 B 0.43821f
C79 VTAIL.t2 B 1.04241f
C80 VTAIL.n2 B 0.644759f
C81 VTAIL.t4 B 0.108424f
C82 VTAIL.t3 B 0.108424f
C83 VTAIL.n3 B 0.815794f
C84 VTAIL.n4 B 1.57528f
C85 VTAIL.t11 B 0.108424f
C86 VTAIL.t6 B 0.108424f
C87 VTAIL.n5 B 0.815798f
C88 VTAIL.n6 B 1.57528f
C89 VTAIL.t10 B 1.04241f
C90 VTAIL.n7 B 0.644752f
C91 VTAIL.t0 B 0.108424f
C92 VTAIL.t1 B 0.108424f
C93 VTAIL.n8 B 0.815798f
C94 VTAIL.n9 B 0.575665f
C95 VTAIL.t5 B 1.04241f
C96 VTAIL.n10 B 1.45419f
C97 VTAIL.t8 B 1.04241f
C98 VTAIL.n11 B 1.40147f
C99 VN.n0 B 0.039363f
C100 VN.t0 B 0.834116f
C101 VN.n1 B 0.042753f
C102 VN.t2 B 1.02355f
C103 VN.n2 B 0.386927f
C104 VN.t1 B 0.834116f
C105 VN.n3 B 0.416706f
C106 VN.n4 B 0.055645f
C107 VN.n5 B 0.251984f
C108 VN.n6 B 0.029857f
C109 VN.n7 B 0.029857f
C110 VN.n8 B 0.044417f
C111 VN.n9 B 0.054547f
C112 VN.n10 B 0.430993f
C113 VN.n11 B 0.033208f
C114 VN.n12 B 0.039363f
C115 VN.t3 B 0.834116f
C116 VN.n13 B 0.042753f
C117 VN.t5 B 1.02355f
C118 VN.n14 B 0.386927f
C119 VN.t4 B 0.834116f
C120 VN.n15 B 0.416706f
C121 VN.n16 B 0.055645f
C122 VN.n17 B 0.251984f
C123 VN.n18 B 0.029857f
C124 VN.n19 B 0.029857f
C125 VN.n20 B 0.044417f
C126 VN.n21 B 0.054547f
C127 VN.n22 B 0.430993f
C128 VN.n23 B 1.25786f
.ends

