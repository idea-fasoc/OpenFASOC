* NGSPICE file created from diff_pair_sample_0409.ext - technology: sky130A

.subckt diff_pair_sample_0409 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=0 ps=0 w=18.51 l=0.39
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=7.2189 ps=37.8 w=18.51 l=0.39
X2 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=7.2189 ps=37.8 w=18.51 l=0.39
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=0 ps=0 w=18.51 l=0.39
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=0 ps=0 w=18.51 l=0.39
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=7.2189 ps=37.8 w=18.51 l=0.39
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=0 ps=0 w=18.51 l=0.39
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.2189 pd=37.8 as=7.2189 ps=37.8 w=18.51 l=0.39
R0 B.n97 B.t2 1353.63
R1 B.n94 B.t13 1353.63
R2 B.n410 B.t10 1353.63
R3 B.n416 B.t6 1353.63
R4 B.n767 B.n766 585
R5 B.n768 B.n767 585
R6 B.n356 B.n93 585
R7 B.n355 B.n354 585
R8 B.n353 B.n352 585
R9 B.n351 B.n350 585
R10 B.n349 B.n348 585
R11 B.n347 B.n346 585
R12 B.n345 B.n344 585
R13 B.n343 B.n342 585
R14 B.n341 B.n340 585
R15 B.n339 B.n338 585
R16 B.n337 B.n336 585
R17 B.n335 B.n334 585
R18 B.n333 B.n332 585
R19 B.n331 B.n330 585
R20 B.n329 B.n328 585
R21 B.n327 B.n326 585
R22 B.n325 B.n324 585
R23 B.n323 B.n322 585
R24 B.n321 B.n320 585
R25 B.n319 B.n318 585
R26 B.n317 B.n316 585
R27 B.n315 B.n314 585
R28 B.n313 B.n312 585
R29 B.n311 B.n310 585
R30 B.n309 B.n308 585
R31 B.n307 B.n306 585
R32 B.n305 B.n304 585
R33 B.n303 B.n302 585
R34 B.n301 B.n300 585
R35 B.n299 B.n298 585
R36 B.n297 B.n296 585
R37 B.n295 B.n294 585
R38 B.n293 B.n292 585
R39 B.n291 B.n290 585
R40 B.n289 B.n288 585
R41 B.n287 B.n286 585
R42 B.n285 B.n284 585
R43 B.n283 B.n282 585
R44 B.n281 B.n280 585
R45 B.n279 B.n278 585
R46 B.n277 B.n276 585
R47 B.n275 B.n274 585
R48 B.n273 B.n272 585
R49 B.n271 B.n270 585
R50 B.n269 B.n268 585
R51 B.n267 B.n266 585
R52 B.n265 B.n264 585
R53 B.n263 B.n262 585
R54 B.n261 B.n260 585
R55 B.n259 B.n258 585
R56 B.n257 B.n256 585
R57 B.n255 B.n254 585
R58 B.n253 B.n252 585
R59 B.n251 B.n250 585
R60 B.n249 B.n248 585
R61 B.n247 B.n246 585
R62 B.n245 B.n244 585
R63 B.n243 B.n242 585
R64 B.n241 B.n240 585
R65 B.n239 B.n238 585
R66 B.n237 B.n236 585
R67 B.n235 B.n234 585
R68 B.n233 B.n232 585
R69 B.n231 B.n230 585
R70 B.n229 B.n228 585
R71 B.n227 B.n226 585
R72 B.n225 B.n224 585
R73 B.n223 B.n222 585
R74 B.n221 B.n220 585
R75 B.n218 B.n217 585
R76 B.n216 B.n215 585
R77 B.n214 B.n213 585
R78 B.n212 B.n211 585
R79 B.n210 B.n209 585
R80 B.n208 B.n207 585
R81 B.n206 B.n205 585
R82 B.n204 B.n203 585
R83 B.n202 B.n201 585
R84 B.n200 B.n199 585
R85 B.n198 B.n197 585
R86 B.n196 B.n195 585
R87 B.n194 B.n193 585
R88 B.n192 B.n191 585
R89 B.n190 B.n189 585
R90 B.n188 B.n187 585
R91 B.n186 B.n185 585
R92 B.n184 B.n183 585
R93 B.n182 B.n181 585
R94 B.n180 B.n179 585
R95 B.n178 B.n177 585
R96 B.n176 B.n175 585
R97 B.n174 B.n173 585
R98 B.n172 B.n171 585
R99 B.n170 B.n169 585
R100 B.n168 B.n167 585
R101 B.n166 B.n165 585
R102 B.n164 B.n163 585
R103 B.n162 B.n161 585
R104 B.n160 B.n159 585
R105 B.n158 B.n157 585
R106 B.n156 B.n155 585
R107 B.n154 B.n153 585
R108 B.n152 B.n151 585
R109 B.n150 B.n149 585
R110 B.n148 B.n147 585
R111 B.n146 B.n145 585
R112 B.n144 B.n143 585
R113 B.n142 B.n141 585
R114 B.n140 B.n139 585
R115 B.n138 B.n137 585
R116 B.n136 B.n135 585
R117 B.n134 B.n133 585
R118 B.n132 B.n131 585
R119 B.n130 B.n129 585
R120 B.n128 B.n127 585
R121 B.n126 B.n125 585
R122 B.n124 B.n123 585
R123 B.n122 B.n121 585
R124 B.n120 B.n119 585
R125 B.n118 B.n117 585
R126 B.n116 B.n115 585
R127 B.n114 B.n113 585
R128 B.n112 B.n111 585
R129 B.n110 B.n109 585
R130 B.n108 B.n107 585
R131 B.n106 B.n105 585
R132 B.n104 B.n103 585
R133 B.n102 B.n101 585
R134 B.n100 B.n99 585
R135 B.n26 B.n25 585
R136 B.n765 B.n27 585
R137 B.n769 B.n27 585
R138 B.n764 B.n763 585
R139 B.n763 B.n23 585
R140 B.n762 B.n22 585
R141 B.n775 B.n22 585
R142 B.n761 B.n21 585
R143 B.n776 B.n21 585
R144 B.n760 B.n20 585
R145 B.n777 B.n20 585
R146 B.n759 B.n758 585
R147 B.n758 B.n16 585
R148 B.n757 B.n15 585
R149 B.n783 B.n15 585
R150 B.n756 B.n14 585
R151 B.n784 B.n14 585
R152 B.n755 B.n13 585
R153 B.n785 B.n13 585
R154 B.n754 B.n753 585
R155 B.n753 B.n12 585
R156 B.n752 B.n751 585
R157 B.n752 B.n8 585
R158 B.n750 B.n7 585
R159 B.n792 B.n7 585
R160 B.n749 B.n6 585
R161 B.n793 B.n6 585
R162 B.n748 B.n5 585
R163 B.n794 B.n5 585
R164 B.n747 B.n746 585
R165 B.n746 B.n4 585
R166 B.n745 B.n357 585
R167 B.n745 B.n744 585
R168 B.n734 B.n358 585
R169 B.n737 B.n358 585
R170 B.n736 B.n735 585
R171 B.n738 B.n736 585
R172 B.n733 B.n363 585
R173 B.n363 B.n362 585
R174 B.n732 B.n731 585
R175 B.n731 B.n730 585
R176 B.n365 B.n364 585
R177 B.n366 B.n365 585
R178 B.n723 B.n722 585
R179 B.n724 B.n723 585
R180 B.n721 B.n371 585
R181 B.n371 B.n370 585
R182 B.n720 B.n719 585
R183 B.n719 B.n718 585
R184 B.n373 B.n372 585
R185 B.n374 B.n373 585
R186 B.n711 B.n710 585
R187 B.n712 B.n711 585
R188 B.n377 B.n376 585
R189 B.n451 B.n450 585
R190 B.n452 B.n448 585
R191 B.n448 B.n378 585
R192 B.n454 B.n453 585
R193 B.n456 B.n447 585
R194 B.n459 B.n458 585
R195 B.n460 B.n446 585
R196 B.n462 B.n461 585
R197 B.n464 B.n445 585
R198 B.n467 B.n466 585
R199 B.n468 B.n444 585
R200 B.n470 B.n469 585
R201 B.n472 B.n443 585
R202 B.n475 B.n474 585
R203 B.n476 B.n442 585
R204 B.n478 B.n477 585
R205 B.n480 B.n441 585
R206 B.n483 B.n482 585
R207 B.n484 B.n440 585
R208 B.n486 B.n485 585
R209 B.n488 B.n439 585
R210 B.n491 B.n490 585
R211 B.n492 B.n438 585
R212 B.n494 B.n493 585
R213 B.n496 B.n437 585
R214 B.n499 B.n498 585
R215 B.n500 B.n436 585
R216 B.n502 B.n501 585
R217 B.n504 B.n435 585
R218 B.n507 B.n506 585
R219 B.n508 B.n434 585
R220 B.n510 B.n509 585
R221 B.n512 B.n433 585
R222 B.n515 B.n514 585
R223 B.n516 B.n432 585
R224 B.n518 B.n517 585
R225 B.n520 B.n431 585
R226 B.n523 B.n522 585
R227 B.n524 B.n430 585
R228 B.n526 B.n525 585
R229 B.n528 B.n429 585
R230 B.n531 B.n530 585
R231 B.n532 B.n428 585
R232 B.n534 B.n533 585
R233 B.n536 B.n427 585
R234 B.n539 B.n538 585
R235 B.n540 B.n426 585
R236 B.n542 B.n541 585
R237 B.n544 B.n425 585
R238 B.n547 B.n546 585
R239 B.n548 B.n424 585
R240 B.n550 B.n549 585
R241 B.n552 B.n423 585
R242 B.n555 B.n554 585
R243 B.n556 B.n422 585
R244 B.n558 B.n557 585
R245 B.n560 B.n421 585
R246 B.n563 B.n562 585
R247 B.n564 B.n420 585
R248 B.n566 B.n565 585
R249 B.n568 B.n419 585
R250 B.n571 B.n570 585
R251 B.n572 B.n415 585
R252 B.n574 B.n573 585
R253 B.n576 B.n414 585
R254 B.n579 B.n578 585
R255 B.n580 B.n413 585
R256 B.n582 B.n581 585
R257 B.n584 B.n412 585
R258 B.n587 B.n586 585
R259 B.n589 B.n409 585
R260 B.n591 B.n590 585
R261 B.n593 B.n408 585
R262 B.n596 B.n595 585
R263 B.n597 B.n407 585
R264 B.n599 B.n598 585
R265 B.n601 B.n406 585
R266 B.n604 B.n603 585
R267 B.n605 B.n405 585
R268 B.n607 B.n606 585
R269 B.n609 B.n404 585
R270 B.n612 B.n611 585
R271 B.n613 B.n403 585
R272 B.n615 B.n614 585
R273 B.n617 B.n402 585
R274 B.n620 B.n619 585
R275 B.n621 B.n401 585
R276 B.n623 B.n622 585
R277 B.n625 B.n400 585
R278 B.n628 B.n627 585
R279 B.n629 B.n399 585
R280 B.n631 B.n630 585
R281 B.n633 B.n398 585
R282 B.n636 B.n635 585
R283 B.n637 B.n397 585
R284 B.n639 B.n638 585
R285 B.n641 B.n396 585
R286 B.n644 B.n643 585
R287 B.n645 B.n395 585
R288 B.n647 B.n646 585
R289 B.n649 B.n394 585
R290 B.n652 B.n651 585
R291 B.n653 B.n393 585
R292 B.n655 B.n654 585
R293 B.n657 B.n392 585
R294 B.n660 B.n659 585
R295 B.n661 B.n391 585
R296 B.n663 B.n662 585
R297 B.n665 B.n390 585
R298 B.n668 B.n667 585
R299 B.n669 B.n389 585
R300 B.n671 B.n670 585
R301 B.n673 B.n388 585
R302 B.n676 B.n675 585
R303 B.n677 B.n387 585
R304 B.n679 B.n678 585
R305 B.n681 B.n386 585
R306 B.n684 B.n683 585
R307 B.n685 B.n385 585
R308 B.n687 B.n686 585
R309 B.n689 B.n384 585
R310 B.n692 B.n691 585
R311 B.n693 B.n383 585
R312 B.n695 B.n694 585
R313 B.n697 B.n382 585
R314 B.n700 B.n699 585
R315 B.n701 B.n381 585
R316 B.n703 B.n702 585
R317 B.n705 B.n380 585
R318 B.n708 B.n707 585
R319 B.n709 B.n379 585
R320 B.n714 B.n713 585
R321 B.n713 B.n712 585
R322 B.n715 B.n375 585
R323 B.n375 B.n374 585
R324 B.n717 B.n716 585
R325 B.n718 B.n717 585
R326 B.n369 B.n368 585
R327 B.n370 B.n369 585
R328 B.n726 B.n725 585
R329 B.n725 B.n724 585
R330 B.n727 B.n367 585
R331 B.n367 B.n366 585
R332 B.n729 B.n728 585
R333 B.n730 B.n729 585
R334 B.n361 B.n360 585
R335 B.n362 B.n361 585
R336 B.n740 B.n739 585
R337 B.n739 B.n738 585
R338 B.n741 B.n359 585
R339 B.n737 B.n359 585
R340 B.n743 B.n742 585
R341 B.n744 B.n743 585
R342 B.n3 B.n0 585
R343 B.n4 B.n3 585
R344 B.n791 B.n1 585
R345 B.n792 B.n791 585
R346 B.n790 B.n789 585
R347 B.n790 B.n8 585
R348 B.n788 B.n9 585
R349 B.n12 B.n9 585
R350 B.n787 B.n786 585
R351 B.n786 B.n785 585
R352 B.n11 B.n10 585
R353 B.n784 B.n11 585
R354 B.n782 B.n781 585
R355 B.n783 B.n782 585
R356 B.n780 B.n17 585
R357 B.n17 B.n16 585
R358 B.n779 B.n778 585
R359 B.n778 B.n777 585
R360 B.n19 B.n18 585
R361 B.n776 B.n19 585
R362 B.n774 B.n773 585
R363 B.n775 B.n774 585
R364 B.n772 B.n24 585
R365 B.n24 B.n23 585
R366 B.n771 B.n770 585
R367 B.n770 B.n769 585
R368 B.n795 B.n794 585
R369 B.n793 B.n2 585
R370 B.n770 B.n26 492.5
R371 B.n767 B.n27 492.5
R372 B.n711 B.n379 492.5
R373 B.n713 B.n377 492.5
R374 B.n768 B.n92 256.663
R375 B.n768 B.n91 256.663
R376 B.n768 B.n90 256.663
R377 B.n768 B.n89 256.663
R378 B.n768 B.n88 256.663
R379 B.n768 B.n87 256.663
R380 B.n768 B.n86 256.663
R381 B.n768 B.n85 256.663
R382 B.n768 B.n84 256.663
R383 B.n768 B.n83 256.663
R384 B.n768 B.n82 256.663
R385 B.n768 B.n81 256.663
R386 B.n768 B.n80 256.663
R387 B.n768 B.n79 256.663
R388 B.n768 B.n78 256.663
R389 B.n768 B.n77 256.663
R390 B.n768 B.n76 256.663
R391 B.n768 B.n75 256.663
R392 B.n768 B.n74 256.663
R393 B.n768 B.n73 256.663
R394 B.n768 B.n72 256.663
R395 B.n768 B.n71 256.663
R396 B.n768 B.n70 256.663
R397 B.n768 B.n69 256.663
R398 B.n768 B.n68 256.663
R399 B.n768 B.n67 256.663
R400 B.n768 B.n66 256.663
R401 B.n768 B.n65 256.663
R402 B.n768 B.n64 256.663
R403 B.n768 B.n63 256.663
R404 B.n768 B.n62 256.663
R405 B.n768 B.n61 256.663
R406 B.n768 B.n60 256.663
R407 B.n768 B.n59 256.663
R408 B.n768 B.n58 256.663
R409 B.n768 B.n57 256.663
R410 B.n768 B.n56 256.663
R411 B.n768 B.n55 256.663
R412 B.n768 B.n54 256.663
R413 B.n768 B.n53 256.663
R414 B.n768 B.n52 256.663
R415 B.n768 B.n51 256.663
R416 B.n768 B.n50 256.663
R417 B.n768 B.n49 256.663
R418 B.n768 B.n48 256.663
R419 B.n768 B.n47 256.663
R420 B.n768 B.n46 256.663
R421 B.n768 B.n45 256.663
R422 B.n768 B.n44 256.663
R423 B.n768 B.n43 256.663
R424 B.n768 B.n42 256.663
R425 B.n768 B.n41 256.663
R426 B.n768 B.n40 256.663
R427 B.n768 B.n39 256.663
R428 B.n768 B.n38 256.663
R429 B.n768 B.n37 256.663
R430 B.n768 B.n36 256.663
R431 B.n768 B.n35 256.663
R432 B.n768 B.n34 256.663
R433 B.n768 B.n33 256.663
R434 B.n768 B.n32 256.663
R435 B.n768 B.n31 256.663
R436 B.n768 B.n30 256.663
R437 B.n768 B.n29 256.663
R438 B.n768 B.n28 256.663
R439 B.n449 B.n378 256.663
R440 B.n455 B.n378 256.663
R441 B.n457 B.n378 256.663
R442 B.n463 B.n378 256.663
R443 B.n465 B.n378 256.663
R444 B.n471 B.n378 256.663
R445 B.n473 B.n378 256.663
R446 B.n479 B.n378 256.663
R447 B.n481 B.n378 256.663
R448 B.n487 B.n378 256.663
R449 B.n489 B.n378 256.663
R450 B.n495 B.n378 256.663
R451 B.n497 B.n378 256.663
R452 B.n503 B.n378 256.663
R453 B.n505 B.n378 256.663
R454 B.n511 B.n378 256.663
R455 B.n513 B.n378 256.663
R456 B.n519 B.n378 256.663
R457 B.n521 B.n378 256.663
R458 B.n527 B.n378 256.663
R459 B.n529 B.n378 256.663
R460 B.n535 B.n378 256.663
R461 B.n537 B.n378 256.663
R462 B.n543 B.n378 256.663
R463 B.n545 B.n378 256.663
R464 B.n551 B.n378 256.663
R465 B.n553 B.n378 256.663
R466 B.n559 B.n378 256.663
R467 B.n561 B.n378 256.663
R468 B.n567 B.n378 256.663
R469 B.n569 B.n378 256.663
R470 B.n575 B.n378 256.663
R471 B.n577 B.n378 256.663
R472 B.n583 B.n378 256.663
R473 B.n585 B.n378 256.663
R474 B.n592 B.n378 256.663
R475 B.n594 B.n378 256.663
R476 B.n600 B.n378 256.663
R477 B.n602 B.n378 256.663
R478 B.n608 B.n378 256.663
R479 B.n610 B.n378 256.663
R480 B.n616 B.n378 256.663
R481 B.n618 B.n378 256.663
R482 B.n624 B.n378 256.663
R483 B.n626 B.n378 256.663
R484 B.n632 B.n378 256.663
R485 B.n634 B.n378 256.663
R486 B.n640 B.n378 256.663
R487 B.n642 B.n378 256.663
R488 B.n648 B.n378 256.663
R489 B.n650 B.n378 256.663
R490 B.n656 B.n378 256.663
R491 B.n658 B.n378 256.663
R492 B.n664 B.n378 256.663
R493 B.n666 B.n378 256.663
R494 B.n672 B.n378 256.663
R495 B.n674 B.n378 256.663
R496 B.n680 B.n378 256.663
R497 B.n682 B.n378 256.663
R498 B.n688 B.n378 256.663
R499 B.n690 B.n378 256.663
R500 B.n696 B.n378 256.663
R501 B.n698 B.n378 256.663
R502 B.n704 B.n378 256.663
R503 B.n706 B.n378 256.663
R504 B.n797 B.n796 256.663
R505 B.n101 B.n100 163.367
R506 B.n105 B.n104 163.367
R507 B.n109 B.n108 163.367
R508 B.n113 B.n112 163.367
R509 B.n117 B.n116 163.367
R510 B.n121 B.n120 163.367
R511 B.n125 B.n124 163.367
R512 B.n129 B.n128 163.367
R513 B.n133 B.n132 163.367
R514 B.n137 B.n136 163.367
R515 B.n141 B.n140 163.367
R516 B.n145 B.n144 163.367
R517 B.n149 B.n148 163.367
R518 B.n153 B.n152 163.367
R519 B.n157 B.n156 163.367
R520 B.n161 B.n160 163.367
R521 B.n165 B.n164 163.367
R522 B.n169 B.n168 163.367
R523 B.n173 B.n172 163.367
R524 B.n177 B.n176 163.367
R525 B.n181 B.n180 163.367
R526 B.n185 B.n184 163.367
R527 B.n189 B.n188 163.367
R528 B.n193 B.n192 163.367
R529 B.n197 B.n196 163.367
R530 B.n201 B.n200 163.367
R531 B.n205 B.n204 163.367
R532 B.n209 B.n208 163.367
R533 B.n213 B.n212 163.367
R534 B.n217 B.n216 163.367
R535 B.n222 B.n221 163.367
R536 B.n226 B.n225 163.367
R537 B.n230 B.n229 163.367
R538 B.n234 B.n233 163.367
R539 B.n238 B.n237 163.367
R540 B.n242 B.n241 163.367
R541 B.n246 B.n245 163.367
R542 B.n250 B.n249 163.367
R543 B.n254 B.n253 163.367
R544 B.n258 B.n257 163.367
R545 B.n262 B.n261 163.367
R546 B.n266 B.n265 163.367
R547 B.n270 B.n269 163.367
R548 B.n274 B.n273 163.367
R549 B.n278 B.n277 163.367
R550 B.n282 B.n281 163.367
R551 B.n286 B.n285 163.367
R552 B.n290 B.n289 163.367
R553 B.n294 B.n293 163.367
R554 B.n298 B.n297 163.367
R555 B.n302 B.n301 163.367
R556 B.n306 B.n305 163.367
R557 B.n310 B.n309 163.367
R558 B.n314 B.n313 163.367
R559 B.n318 B.n317 163.367
R560 B.n322 B.n321 163.367
R561 B.n326 B.n325 163.367
R562 B.n330 B.n329 163.367
R563 B.n334 B.n333 163.367
R564 B.n338 B.n337 163.367
R565 B.n342 B.n341 163.367
R566 B.n346 B.n345 163.367
R567 B.n350 B.n349 163.367
R568 B.n354 B.n353 163.367
R569 B.n767 B.n93 163.367
R570 B.n711 B.n373 163.367
R571 B.n719 B.n373 163.367
R572 B.n719 B.n371 163.367
R573 B.n723 B.n371 163.367
R574 B.n723 B.n365 163.367
R575 B.n731 B.n365 163.367
R576 B.n731 B.n363 163.367
R577 B.n736 B.n363 163.367
R578 B.n736 B.n358 163.367
R579 B.n745 B.n358 163.367
R580 B.n746 B.n745 163.367
R581 B.n746 B.n5 163.367
R582 B.n6 B.n5 163.367
R583 B.n7 B.n6 163.367
R584 B.n752 B.n7 163.367
R585 B.n753 B.n752 163.367
R586 B.n753 B.n13 163.367
R587 B.n14 B.n13 163.367
R588 B.n15 B.n14 163.367
R589 B.n758 B.n15 163.367
R590 B.n758 B.n20 163.367
R591 B.n21 B.n20 163.367
R592 B.n22 B.n21 163.367
R593 B.n763 B.n22 163.367
R594 B.n763 B.n27 163.367
R595 B.n450 B.n448 163.367
R596 B.n454 B.n448 163.367
R597 B.n458 B.n456 163.367
R598 B.n462 B.n446 163.367
R599 B.n466 B.n464 163.367
R600 B.n470 B.n444 163.367
R601 B.n474 B.n472 163.367
R602 B.n478 B.n442 163.367
R603 B.n482 B.n480 163.367
R604 B.n486 B.n440 163.367
R605 B.n490 B.n488 163.367
R606 B.n494 B.n438 163.367
R607 B.n498 B.n496 163.367
R608 B.n502 B.n436 163.367
R609 B.n506 B.n504 163.367
R610 B.n510 B.n434 163.367
R611 B.n514 B.n512 163.367
R612 B.n518 B.n432 163.367
R613 B.n522 B.n520 163.367
R614 B.n526 B.n430 163.367
R615 B.n530 B.n528 163.367
R616 B.n534 B.n428 163.367
R617 B.n538 B.n536 163.367
R618 B.n542 B.n426 163.367
R619 B.n546 B.n544 163.367
R620 B.n550 B.n424 163.367
R621 B.n554 B.n552 163.367
R622 B.n558 B.n422 163.367
R623 B.n562 B.n560 163.367
R624 B.n566 B.n420 163.367
R625 B.n570 B.n568 163.367
R626 B.n574 B.n415 163.367
R627 B.n578 B.n576 163.367
R628 B.n582 B.n413 163.367
R629 B.n586 B.n584 163.367
R630 B.n591 B.n409 163.367
R631 B.n595 B.n593 163.367
R632 B.n599 B.n407 163.367
R633 B.n603 B.n601 163.367
R634 B.n607 B.n405 163.367
R635 B.n611 B.n609 163.367
R636 B.n615 B.n403 163.367
R637 B.n619 B.n617 163.367
R638 B.n623 B.n401 163.367
R639 B.n627 B.n625 163.367
R640 B.n631 B.n399 163.367
R641 B.n635 B.n633 163.367
R642 B.n639 B.n397 163.367
R643 B.n643 B.n641 163.367
R644 B.n647 B.n395 163.367
R645 B.n651 B.n649 163.367
R646 B.n655 B.n393 163.367
R647 B.n659 B.n657 163.367
R648 B.n663 B.n391 163.367
R649 B.n667 B.n665 163.367
R650 B.n671 B.n389 163.367
R651 B.n675 B.n673 163.367
R652 B.n679 B.n387 163.367
R653 B.n683 B.n681 163.367
R654 B.n687 B.n385 163.367
R655 B.n691 B.n689 163.367
R656 B.n695 B.n383 163.367
R657 B.n699 B.n697 163.367
R658 B.n703 B.n381 163.367
R659 B.n707 B.n705 163.367
R660 B.n713 B.n375 163.367
R661 B.n717 B.n375 163.367
R662 B.n717 B.n369 163.367
R663 B.n725 B.n369 163.367
R664 B.n725 B.n367 163.367
R665 B.n729 B.n367 163.367
R666 B.n729 B.n361 163.367
R667 B.n739 B.n361 163.367
R668 B.n739 B.n359 163.367
R669 B.n743 B.n359 163.367
R670 B.n743 B.n3 163.367
R671 B.n795 B.n3 163.367
R672 B.n791 B.n2 163.367
R673 B.n791 B.n790 163.367
R674 B.n790 B.n9 163.367
R675 B.n786 B.n9 163.367
R676 B.n786 B.n11 163.367
R677 B.n782 B.n11 163.367
R678 B.n782 B.n17 163.367
R679 B.n778 B.n17 163.367
R680 B.n778 B.n19 163.367
R681 B.n774 B.n19 163.367
R682 B.n774 B.n24 163.367
R683 B.n770 B.n24 163.367
R684 B.n94 B.t14 84.0918
R685 B.n410 B.t12 84.0918
R686 B.n97 B.t4 84.0671
R687 B.n416 B.t9 84.0671
R688 B.n28 B.n26 71.676
R689 B.n101 B.n29 71.676
R690 B.n105 B.n30 71.676
R691 B.n109 B.n31 71.676
R692 B.n113 B.n32 71.676
R693 B.n117 B.n33 71.676
R694 B.n121 B.n34 71.676
R695 B.n125 B.n35 71.676
R696 B.n129 B.n36 71.676
R697 B.n133 B.n37 71.676
R698 B.n137 B.n38 71.676
R699 B.n141 B.n39 71.676
R700 B.n145 B.n40 71.676
R701 B.n149 B.n41 71.676
R702 B.n153 B.n42 71.676
R703 B.n157 B.n43 71.676
R704 B.n161 B.n44 71.676
R705 B.n165 B.n45 71.676
R706 B.n169 B.n46 71.676
R707 B.n173 B.n47 71.676
R708 B.n177 B.n48 71.676
R709 B.n181 B.n49 71.676
R710 B.n185 B.n50 71.676
R711 B.n189 B.n51 71.676
R712 B.n193 B.n52 71.676
R713 B.n197 B.n53 71.676
R714 B.n201 B.n54 71.676
R715 B.n205 B.n55 71.676
R716 B.n209 B.n56 71.676
R717 B.n213 B.n57 71.676
R718 B.n217 B.n58 71.676
R719 B.n222 B.n59 71.676
R720 B.n226 B.n60 71.676
R721 B.n230 B.n61 71.676
R722 B.n234 B.n62 71.676
R723 B.n238 B.n63 71.676
R724 B.n242 B.n64 71.676
R725 B.n246 B.n65 71.676
R726 B.n250 B.n66 71.676
R727 B.n254 B.n67 71.676
R728 B.n258 B.n68 71.676
R729 B.n262 B.n69 71.676
R730 B.n266 B.n70 71.676
R731 B.n270 B.n71 71.676
R732 B.n274 B.n72 71.676
R733 B.n278 B.n73 71.676
R734 B.n282 B.n74 71.676
R735 B.n286 B.n75 71.676
R736 B.n290 B.n76 71.676
R737 B.n294 B.n77 71.676
R738 B.n298 B.n78 71.676
R739 B.n302 B.n79 71.676
R740 B.n306 B.n80 71.676
R741 B.n310 B.n81 71.676
R742 B.n314 B.n82 71.676
R743 B.n318 B.n83 71.676
R744 B.n322 B.n84 71.676
R745 B.n326 B.n85 71.676
R746 B.n330 B.n86 71.676
R747 B.n334 B.n87 71.676
R748 B.n338 B.n88 71.676
R749 B.n342 B.n89 71.676
R750 B.n346 B.n90 71.676
R751 B.n350 B.n91 71.676
R752 B.n354 B.n92 71.676
R753 B.n93 B.n92 71.676
R754 B.n353 B.n91 71.676
R755 B.n349 B.n90 71.676
R756 B.n345 B.n89 71.676
R757 B.n341 B.n88 71.676
R758 B.n337 B.n87 71.676
R759 B.n333 B.n86 71.676
R760 B.n329 B.n85 71.676
R761 B.n325 B.n84 71.676
R762 B.n321 B.n83 71.676
R763 B.n317 B.n82 71.676
R764 B.n313 B.n81 71.676
R765 B.n309 B.n80 71.676
R766 B.n305 B.n79 71.676
R767 B.n301 B.n78 71.676
R768 B.n297 B.n77 71.676
R769 B.n293 B.n76 71.676
R770 B.n289 B.n75 71.676
R771 B.n285 B.n74 71.676
R772 B.n281 B.n73 71.676
R773 B.n277 B.n72 71.676
R774 B.n273 B.n71 71.676
R775 B.n269 B.n70 71.676
R776 B.n265 B.n69 71.676
R777 B.n261 B.n68 71.676
R778 B.n257 B.n67 71.676
R779 B.n253 B.n66 71.676
R780 B.n249 B.n65 71.676
R781 B.n245 B.n64 71.676
R782 B.n241 B.n63 71.676
R783 B.n237 B.n62 71.676
R784 B.n233 B.n61 71.676
R785 B.n229 B.n60 71.676
R786 B.n225 B.n59 71.676
R787 B.n221 B.n58 71.676
R788 B.n216 B.n57 71.676
R789 B.n212 B.n56 71.676
R790 B.n208 B.n55 71.676
R791 B.n204 B.n54 71.676
R792 B.n200 B.n53 71.676
R793 B.n196 B.n52 71.676
R794 B.n192 B.n51 71.676
R795 B.n188 B.n50 71.676
R796 B.n184 B.n49 71.676
R797 B.n180 B.n48 71.676
R798 B.n176 B.n47 71.676
R799 B.n172 B.n46 71.676
R800 B.n168 B.n45 71.676
R801 B.n164 B.n44 71.676
R802 B.n160 B.n43 71.676
R803 B.n156 B.n42 71.676
R804 B.n152 B.n41 71.676
R805 B.n148 B.n40 71.676
R806 B.n144 B.n39 71.676
R807 B.n140 B.n38 71.676
R808 B.n136 B.n37 71.676
R809 B.n132 B.n36 71.676
R810 B.n128 B.n35 71.676
R811 B.n124 B.n34 71.676
R812 B.n120 B.n33 71.676
R813 B.n116 B.n32 71.676
R814 B.n112 B.n31 71.676
R815 B.n108 B.n30 71.676
R816 B.n104 B.n29 71.676
R817 B.n100 B.n28 71.676
R818 B.n449 B.n377 71.676
R819 B.n455 B.n454 71.676
R820 B.n458 B.n457 71.676
R821 B.n463 B.n462 71.676
R822 B.n466 B.n465 71.676
R823 B.n471 B.n470 71.676
R824 B.n474 B.n473 71.676
R825 B.n479 B.n478 71.676
R826 B.n482 B.n481 71.676
R827 B.n487 B.n486 71.676
R828 B.n490 B.n489 71.676
R829 B.n495 B.n494 71.676
R830 B.n498 B.n497 71.676
R831 B.n503 B.n502 71.676
R832 B.n506 B.n505 71.676
R833 B.n511 B.n510 71.676
R834 B.n514 B.n513 71.676
R835 B.n519 B.n518 71.676
R836 B.n522 B.n521 71.676
R837 B.n527 B.n526 71.676
R838 B.n530 B.n529 71.676
R839 B.n535 B.n534 71.676
R840 B.n538 B.n537 71.676
R841 B.n543 B.n542 71.676
R842 B.n546 B.n545 71.676
R843 B.n551 B.n550 71.676
R844 B.n554 B.n553 71.676
R845 B.n559 B.n558 71.676
R846 B.n562 B.n561 71.676
R847 B.n567 B.n566 71.676
R848 B.n570 B.n569 71.676
R849 B.n575 B.n574 71.676
R850 B.n578 B.n577 71.676
R851 B.n583 B.n582 71.676
R852 B.n586 B.n585 71.676
R853 B.n592 B.n591 71.676
R854 B.n595 B.n594 71.676
R855 B.n600 B.n599 71.676
R856 B.n603 B.n602 71.676
R857 B.n608 B.n607 71.676
R858 B.n611 B.n610 71.676
R859 B.n616 B.n615 71.676
R860 B.n619 B.n618 71.676
R861 B.n624 B.n623 71.676
R862 B.n627 B.n626 71.676
R863 B.n632 B.n631 71.676
R864 B.n635 B.n634 71.676
R865 B.n640 B.n639 71.676
R866 B.n643 B.n642 71.676
R867 B.n648 B.n647 71.676
R868 B.n651 B.n650 71.676
R869 B.n656 B.n655 71.676
R870 B.n659 B.n658 71.676
R871 B.n664 B.n663 71.676
R872 B.n667 B.n666 71.676
R873 B.n672 B.n671 71.676
R874 B.n675 B.n674 71.676
R875 B.n680 B.n679 71.676
R876 B.n683 B.n682 71.676
R877 B.n688 B.n687 71.676
R878 B.n691 B.n690 71.676
R879 B.n696 B.n695 71.676
R880 B.n699 B.n698 71.676
R881 B.n704 B.n703 71.676
R882 B.n707 B.n706 71.676
R883 B.n450 B.n449 71.676
R884 B.n456 B.n455 71.676
R885 B.n457 B.n446 71.676
R886 B.n464 B.n463 71.676
R887 B.n465 B.n444 71.676
R888 B.n472 B.n471 71.676
R889 B.n473 B.n442 71.676
R890 B.n480 B.n479 71.676
R891 B.n481 B.n440 71.676
R892 B.n488 B.n487 71.676
R893 B.n489 B.n438 71.676
R894 B.n496 B.n495 71.676
R895 B.n497 B.n436 71.676
R896 B.n504 B.n503 71.676
R897 B.n505 B.n434 71.676
R898 B.n512 B.n511 71.676
R899 B.n513 B.n432 71.676
R900 B.n520 B.n519 71.676
R901 B.n521 B.n430 71.676
R902 B.n528 B.n527 71.676
R903 B.n529 B.n428 71.676
R904 B.n536 B.n535 71.676
R905 B.n537 B.n426 71.676
R906 B.n544 B.n543 71.676
R907 B.n545 B.n424 71.676
R908 B.n552 B.n551 71.676
R909 B.n553 B.n422 71.676
R910 B.n560 B.n559 71.676
R911 B.n561 B.n420 71.676
R912 B.n568 B.n567 71.676
R913 B.n569 B.n415 71.676
R914 B.n576 B.n575 71.676
R915 B.n577 B.n413 71.676
R916 B.n584 B.n583 71.676
R917 B.n585 B.n409 71.676
R918 B.n593 B.n592 71.676
R919 B.n594 B.n407 71.676
R920 B.n601 B.n600 71.676
R921 B.n602 B.n405 71.676
R922 B.n609 B.n608 71.676
R923 B.n610 B.n403 71.676
R924 B.n617 B.n616 71.676
R925 B.n618 B.n401 71.676
R926 B.n625 B.n624 71.676
R927 B.n626 B.n399 71.676
R928 B.n633 B.n632 71.676
R929 B.n634 B.n397 71.676
R930 B.n641 B.n640 71.676
R931 B.n642 B.n395 71.676
R932 B.n649 B.n648 71.676
R933 B.n650 B.n393 71.676
R934 B.n657 B.n656 71.676
R935 B.n658 B.n391 71.676
R936 B.n665 B.n664 71.676
R937 B.n666 B.n389 71.676
R938 B.n673 B.n672 71.676
R939 B.n674 B.n387 71.676
R940 B.n681 B.n680 71.676
R941 B.n682 B.n385 71.676
R942 B.n689 B.n688 71.676
R943 B.n690 B.n383 71.676
R944 B.n697 B.n696 71.676
R945 B.n698 B.n381 71.676
R946 B.n705 B.n704 71.676
R947 B.n706 B.n379 71.676
R948 B.n796 B.n795 71.676
R949 B.n796 B.n2 71.676
R950 B.n95 B.t15 70.1282
R951 B.n411 B.t11 70.1282
R952 B.n98 B.t5 70.1034
R953 B.n417 B.t8 70.1034
R954 B.n219 B.n98 59.5399
R955 B.n96 B.n95 59.5399
R956 B.n588 B.n411 59.5399
R957 B.n418 B.n417 59.5399
R958 B.n712 B.n378 52.2164
R959 B.n769 B.n768 52.2164
R960 B.n714 B.n376 32.0005
R961 B.n710 B.n709 32.0005
R962 B.n766 B.n765 32.0005
R963 B.n771 B.n25 32.0005
R964 B.n712 B.n374 31.4225
R965 B.n718 B.n374 31.4225
R966 B.n718 B.n370 31.4225
R967 B.n724 B.n370 31.4225
R968 B.n730 B.n366 31.4225
R969 B.n730 B.n362 31.4225
R970 B.n738 B.n362 31.4225
R971 B.n738 B.n737 31.4225
R972 B.n744 B.n4 31.4225
R973 B.n794 B.n4 31.4225
R974 B.n794 B.n793 31.4225
R975 B.n793 B.n792 31.4225
R976 B.n792 B.n8 31.4225
R977 B.n785 B.n12 31.4225
R978 B.n785 B.n784 31.4225
R979 B.n784 B.n783 31.4225
R980 B.n783 B.n16 31.4225
R981 B.n777 B.n776 31.4225
R982 B.n776 B.n775 31.4225
R983 B.n775 B.n23 31.4225
R984 B.n769 B.n23 31.4225
R985 B.n737 B.t0 26.3395
R986 B.n12 B.t1 26.3395
R987 B B.n797 18.0485
R988 B.n724 B.t7 16.1736
R989 B.n777 B.t3 16.1736
R990 B.t7 B.n366 15.2494
R991 B.t3 B.n16 15.2494
R992 B.n98 B.n97 13.9641
R993 B.n95 B.n94 13.9641
R994 B.n411 B.n410 13.9641
R995 B.n417 B.n416 13.9641
R996 B.n715 B.n714 10.6151
R997 B.n716 B.n715 10.6151
R998 B.n716 B.n368 10.6151
R999 B.n726 B.n368 10.6151
R1000 B.n727 B.n726 10.6151
R1001 B.n728 B.n727 10.6151
R1002 B.n728 B.n360 10.6151
R1003 B.n740 B.n360 10.6151
R1004 B.n741 B.n740 10.6151
R1005 B.n742 B.n741 10.6151
R1006 B.n742 B.n0 10.6151
R1007 B.n451 B.n376 10.6151
R1008 B.n452 B.n451 10.6151
R1009 B.n453 B.n452 10.6151
R1010 B.n453 B.n447 10.6151
R1011 B.n459 B.n447 10.6151
R1012 B.n460 B.n459 10.6151
R1013 B.n461 B.n460 10.6151
R1014 B.n461 B.n445 10.6151
R1015 B.n467 B.n445 10.6151
R1016 B.n468 B.n467 10.6151
R1017 B.n469 B.n468 10.6151
R1018 B.n469 B.n443 10.6151
R1019 B.n475 B.n443 10.6151
R1020 B.n476 B.n475 10.6151
R1021 B.n477 B.n476 10.6151
R1022 B.n477 B.n441 10.6151
R1023 B.n483 B.n441 10.6151
R1024 B.n484 B.n483 10.6151
R1025 B.n485 B.n484 10.6151
R1026 B.n485 B.n439 10.6151
R1027 B.n491 B.n439 10.6151
R1028 B.n492 B.n491 10.6151
R1029 B.n493 B.n492 10.6151
R1030 B.n493 B.n437 10.6151
R1031 B.n499 B.n437 10.6151
R1032 B.n500 B.n499 10.6151
R1033 B.n501 B.n500 10.6151
R1034 B.n501 B.n435 10.6151
R1035 B.n507 B.n435 10.6151
R1036 B.n508 B.n507 10.6151
R1037 B.n509 B.n508 10.6151
R1038 B.n509 B.n433 10.6151
R1039 B.n515 B.n433 10.6151
R1040 B.n516 B.n515 10.6151
R1041 B.n517 B.n516 10.6151
R1042 B.n517 B.n431 10.6151
R1043 B.n523 B.n431 10.6151
R1044 B.n524 B.n523 10.6151
R1045 B.n525 B.n524 10.6151
R1046 B.n525 B.n429 10.6151
R1047 B.n531 B.n429 10.6151
R1048 B.n532 B.n531 10.6151
R1049 B.n533 B.n532 10.6151
R1050 B.n533 B.n427 10.6151
R1051 B.n539 B.n427 10.6151
R1052 B.n540 B.n539 10.6151
R1053 B.n541 B.n540 10.6151
R1054 B.n541 B.n425 10.6151
R1055 B.n547 B.n425 10.6151
R1056 B.n548 B.n547 10.6151
R1057 B.n549 B.n548 10.6151
R1058 B.n549 B.n423 10.6151
R1059 B.n555 B.n423 10.6151
R1060 B.n556 B.n555 10.6151
R1061 B.n557 B.n556 10.6151
R1062 B.n557 B.n421 10.6151
R1063 B.n563 B.n421 10.6151
R1064 B.n564 B.n563 10.6151
R1065 B.n565 B.n564 10.6151
R1066 B.n565 B.n419 10.6151
R1067 B.n572 B.n571 10.6151
R1068 B.n573 B.n572 10.6151
R1069 B.n573 B.n414 10.6151
R1070 B.n579 B.n414 10.6151
R1071 B.n580 B.n579 10.6151
R1072 B.n581 B.n580 10.6151
R1073 B.n581 B.n412 10.6151
R1074 B.n587 B.n412 10.6151
R1075 B.n590 B.n589 10.6151
R1076 B.n590 B.n408 10.6151
R1077 B.n596 B.n408 10.6151
R1078 B.n597 B.n596 10.6151
R1079 B.n598 B.n597 10.6151
R1080 B.n598 B.n406 10.6151
R1081 B.n604 B.n406 10.6151
R1082 B.n605 B.n604 10.6151
R1083 B.n606 B.n605 10.6151
R1084 B.n606 B.n404 10.6151
R1085 B.n612 B.n404 10.6151
R1086 B.n613 B.n612 10.6151
R1087 B.n614 B.n613 10.6151
R1088 B.n614 B.n402 10.6151
R1089 B.n620 B.n402 10.6151
R1090 B.n621 B.n620 10.6151
R1091 B.n622 B.n621 10.6151
R1092 B.n622 B.n400 10.6151
R1093 B.n628 B.n400 10.6151
R1094 B.n629 B.n628 10.6151
R1095 B.n630 B.n629 10.6151
R1096 B.n630 B.n398 10.6151
R1097 B.n636 B.n398 10.6151
R1098 B.n637 B.n636 10.6151
R1099 B.n638 B.n637 10.6151
R1100 B.n638 B.n396 10.6151
R1101 B.n644 B.n396 10.6151
R1102 B.n645 B.n644 10.6151
R1103 B.n646 B.n645 10.6151
R1104 B.n646 B.n394 10.6151
R1105 B.n652 B.n394 10.6151
R1106 B.n653 B.n652 10.6151
R1107 B.n654 B.n653 10.6151
R1108 B.n654 B.n392 10.6151
R1109 B.n660 B.n392 10.6151
R1110 B.n661 B.n660 10.6151
R1111 B.n662 B.n661 10.6151
R1112 B.n662 B.n390 10.6151
R1113 B.n668 B.n390 10.6151
R1114 B.n669 B.n668 10.6151
R1115 B.n670 B.n669 10.6151
R1116 B.n670 B.n388 10.6151
R1117 B.n676 B.n388 10.6151
R1118 B.n677 B.n676 10.6151
R1119 B.n678 B.n677 10.6151
R1120 B.n678 B.n386 10.6151
R1121 B.n684 B.n386 10.6151
R1122 B.n685 B.n684 10.6151
R1123 B.n686 B.n685 10.6151
R1124 B.n686 B.n384 10.6151
R1125 B.n692 B.n384 10.6151
R1126 B.n693 B.n692 10.6151
R1127 B.n694 B.n693 10.6151
R1128 B.n694 B.n382 10.6151
R1129 B.n700 B.n382 10.6151
R1130 B.n701 B.n700 10.6151
R1131 B.n702 B.n701 10.6151
R1132 B.n702 B.n380 10.6151
R1133 B.n708 B.n380 10.6151
R1134 B.n709 B.n708 10.6151
R1135 B.n710 B.n372 10.6151
R1136 B.n720 B.n372 10.6151
R1137 B.n721 B.n720 10.6151
R1138 B.n722 B.n721 10.6151
R1139 B.n722 B.n364 10.6151
R1140 B.n732 B.n364 10.6151
R1141 B.n733 B.n732 10.6151
R1142 B.n735 B.n733 10.6151
R1143 B.n735 B.n734 10.6151
R1144 B.n734 B.n357 10.6151
R1145 B.n747 B.n357 10.6151
R1146 B.n748 B.n747 10.6151
R1147 B.n749 B.n748 10.6151
R1148 B.n750 B.n749 10.6151
R1149 B.n751 B.n750 10.6151
R1150 B.n754 B.n751 10.6151
R1151 B.n755 B.n754 10.6151
R1152 B.n756 B.n755 10.6151
R1153 B.n757 B.n756 10.6151
R1154 B.n759 B.n757 10.6151
R1155 B.n760 B.n759 10.6151
R1156 B.n761 B.n760 10.6151
R1157 B.n762 B.n761 10.6151
R1158 B.n764 B.n762 10.6151
R1159 B.n765 B.n764 10.6151
R1160 B.n789 B.n1 10.6151
R1161 B.n789 B.n788 10.6151
R1162 B.n788 B.n787 10.6151
R1163 B.n787 B.n10 10.6151
R1164 B.n781 B.n10 10.6151
R1165 B.n781 B.n780 10.6151
R1166 B.n780 B.n779 10.6151
R1167 B.n779 B.n18 10.6151
R1168 B.n773 B.n18 10.6151
R1169 B.n773 B.n772 10.6151
R1170 B.n772 B.n771 10.6151
R1171 B.n99 B.n25 10.6151
R1172 B.n102 B.n99 10.6151
R1173 B.n103 B.n102 10.6151
R1174 B.n106 B.n103 10.6151
R1175 B.n107 B.n106 10.6151
R1176 B.n110 B.n107 10.6151
R1177 B.n111 B.n110 10.6151
R1178 B.n114 B.n111 10.6151
R1179 B.n115 B.n114 10.6151
R1180 B.n118 B.n115 10.6151
R1181 B.n119 B.n118 10.6151
R1182 B.n122 B.n119 10.6151
R1183 B.n123 B.n122 10.6151
R1184 B.n126 B.n123 10.6151
R1185 B.n127 B.n126 10.6151
R1186 B.n130 B.n127 10.6151
R1187 B.n131 B.n130 10.6151
R1188 B.n134 B.n131 10.6151
R1189 B.n135 B.n134 10.6151
R1190 B.n138 B.n135 10.6151
R1191 B.n139 B.n138 10.6151
R1192 B.n142 B.n139 10.6151
R1193 B.n143 B.n142 10.6151
R1194 B.n146 B.n143 10.6151
R1195 B.n147 B.n146 10.6151
R1196 B.n150 B.n147 10.6151
R1197 B.n151 B.n150 10.6151
R1198 B.n154 B.n151 10.6151
R1199 B.n155 B.n154 10.6151
R1200 B.n158 B.n155 10.6151
R1201 B.n159 B.n158 10.6151
R1202 B.n162 B.n159 10.6151
R1203 B.n163 B.n162 10.6151
R1204 B.n166 B.n163 10.6151
R1205 B.n167 B.n166 10.6151
R1206 B.n170 B.n167 10.6151
R1207 B.n171 B.n170 10.6151
R1208 B.n174 B.n171 10.6151
R1209 B.n175 B.n174 10.6151
R1210 B.n178 B.n175 10.6151
R1211 B.n179 B.n178 10.6151
R1212 B.n182 B.n179 10.6151
R1213 B.n183 B.n182 10.6151
R1214 B.n186 B.n183 10.6151
R1215 B.n187 B.n186 10.6151
R1216 B.n190 B.n187 10.6151
R1217 B.n191 B.n190 10.6151
R1218 B.n194 B.n191 10.6151
R1219 B.n195 B.n194 10.6151
R1220 B.n198 B.n195 10.6151
R1221 B.n199 B.n198 10.6151
R1222 B.n202 B.n199 10.6151
R1223 B.n203 B.n202 10.6151
R1224 B.n206 B.n203 10.6151
R1225 B.n207 B.n206 10.6151
R1226 B.n210 B.n207 10.6151
R1227 B.n211 B.n210 10.6151
R1228 B.n214 B.n211 10.6151
R1229 B.n215 B.n214 10.6151
R1230 B.n218 B.n215 10.6151
R1231 B.n223 B.n220 10.6151
R1232 B.n224 B.n223 10.6151
R1233 B.n227 B.n224 10.6151
R1234 B.n228 B.n227 10.6151
R1235 B.n231 B.n228 10.6151
R1236 B.n232 B.n231 10.6151
R1237 B.n235 B.n232 10.6151
R1238 B.n236 B.n235 10.6151
R1239 B.n240 B.n239 10.6151
R1240 B.n243 B.n240 10.6151
R1241 B.n244 B.n243 10.6151
R1242 B.n247 B.n244 10.6151
R1243 B.n248 B.n247 10.6151
R1244 B.n251 B.n248 10.6151
R1245 B.n252 B.n251 10.6151
R1246 B.n255 B.n252 10.6151
R1247 B.n256 B.n255 10.6151
R1248 B.n259 B.n256 10.6151
R1249 B.n260 B.n259 10.6151
R1250 B.n263 B.n260 10.6151
R1251 B.n264 B.n263 10.6151
R1252 B.n267 B.n264 10.6151
R1253 B.n268 B.n267 10.6151
R1254 B.n271 B.n268 10.6151
R1255 B.n272 B.n271 10.6151
R1256 B.n275 B.n272 10.6151
R1257 B.n276 B.n275 10.6151
R1258 B.n279 B.n276 10.6151
R1259 B.n280 B.n279 10.6151
R1260 B.n283 B.n280 10.6151
R1261 B.n284 B.n283 10.6151
R1262 B.n287 B.n284 10.6151
R1263 B.n288 B.n287 10.6151
R1264 B.n291 B.n288 10.6151
R1265 B.n292 B.n291 10.6151
R1266 B.n295 B.n292 10.6151
R1267 B.n296 B.n295 10.6151
R1268 B.n299 B.n296 10.6151
R1269 B.n300 B.n299 10.6151
R1270 B.n303 B.n300 10.6151
R1271 B.n304 B.n303 10.6151
R1272 B.n307 B.n304 10.6151
R1273 B.n308 B.n307 10.6151
R1274 B.n311 B.n308 10.6151
R1275 B.n312 B.n311 10.6151
R1276 B.n315 B.n312 10.6151
R1277 B.n316 B.n315 10.6151
R1278 B.n319 B.n316 10.6151
R1279 B.n320 B.n319 10.6151
R1280 B.n323 B.n320 10.6151
R1281 B.n324 B.n323 10.6151
R1282 B.n327 B.n324 10.6151
R1283 B.n328 B.n327 10.6151
R1284 B.n331 B.n328 10.6151
R1285 B.n332 B.n331 10.6151
R1286 B.n335 B.n332 10.6151
R1287 B.n336 B.n335 10.6151
R1288 B.n339 B.n336 10.6151
R1289 B.n340 B.n339 10.6151
R1290 B.n343 B.n340 10.6151
R1291 B.n344 B.n343 10.6151
R1292 B.n347 B.n344 10.6151
R1293 B.n348 B.n347 10.6151
R1294 B.n351 B.n348 10.6151
R1295 B.n352 B.n351 10.6151
R1296 B.n355 B.n352 10.6151
R1297 B.n356 B.n355 10.6151
R1298 B.n766 B.n356 10.6151
R1299 B.n797 B.n0 8.11757
R1300 B.n797 B.n1 8.11757
R1301 B.n571 B.n418 7.18099
R1302 B.n588 B.n587 7.18099
R1303 B.n220 B.n219 7.18099
R1304 B.n236 B.n96 7.18099
R1305 B.n744 B.t0 5.08347
R1306 B.t1 B.n8 5.08347
R1307 B.n419 B.n418 3.43465
R1308 B.n589 B.n588 3.43465
R1309 B.n219 B.n218 3.43465
R1310 B.n239 B.n96 3.43465
R1311 VN VN.t0 1450.59
R1312 VN VN.t1 1406.52
R1313 VTAIL.n1 VTAIL.t2 43.2795
R1314 VTAIL.n3 VTAIL.t3 43.2793
R1315 VTAIL.n0 VTAIL.t0 43.2793
R1316 VTAIL.n2 VTAIL.t1 43.2793
R1317 VTAIL.n1 VTAIL.n0 29.5824
R1318 VTAIL.n3 VTAIL.n2 28.9617
R1319 VTAIL.n2 VTAIL.n1 0.780672
R1320 VTAIL VTAIL.n0 0.68369
R1321 VTAIL VTAIL.n3 0.0974828
R1322 VDD2.n0 VDD2.t0 100.834
R1323 VDD2.n0 VDD2.t1 59.9581
R1324 VDD2 VDD2.n0 0.213862
R1325 VP.n0 VP.t1 1450.21
R1326 VP.n0 VP.t0 1406.47
R1327 VP VP.n0 0.0516364
R1328 VDD1 VDD1.t1 101.513
R1329 VDD1 VDD1.t0 60.1715
C0 VDD1 VTAIL 9.412481f
C1 VTAIL VP 1.47973f
C2 VDD2 VTAIL 9.4385f
C3 VDD1 VP 2.42236f
C4 VDD1 VDD2 0.436407f
C5 VDD2 VP 0.243277f
C6 VN VTAIL 1.46468f
C7 VN VDD1 0.148448f
C8 VN VP 5.62701f
C9 VN VDD2 2.335f
C10 VDD2 B 4.813127f
C11 VDD1 B 8.35444f
C12 VTAIL B 7.981565f
C13 VN B 9.69662f
C14 VP B 4.097879f
C15 VDD1.t0 B 3.80705f
C16 VDD1.t1 B 4.53454f
C17 VP.t1 B 1.26094f
C18 VP.t0 B 1.17647f
C19 VP.n0 B 5.55392f
C20 VDD2.t0 B 4.49935f
C21 VDD2.t1 B 3.80039f
C22 VDD2.n0 B 3.36199f
C23 VTAIL.t0 B 3.11205f
C24 VTAIL.n0 B 1.60084f
C25 VTAIL.t2 B 3.11206f
C26 VTAIL.n1 B 1.60667f
C27 VTAIL.t1 B 3.11205f
C28 VTAIL.n2 B 1.56922f
C29 VTAIL.t3 B 3.11205f
C30 VTAIL.n3 B 1.52797f
C31 VN.t1 B 1.15063f
C32 VN.t0 B 1.235f
.ends

