* NGSPICE file created from diff_pair_sample_1694.ext - technology: sky130A

.subckt diff_pair_sample_1694 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0.9702 ps=6.21 w=5.88 l=2.33
X1 VDD1.t7 VP.t0 VTAIL.t0 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=2.2932 ps=12.54 w=5.88 l=2.33
X2 VDD1.t6 VP.t1 VTAIL.t4 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X3 VDD2.t3 VN.t1 VTAIL.t14 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=2.2932 ps=12.54 w=5.88 l=2.33
X4 B.t11 B.t9 B.t10 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0 ps=0 w=5.88 l=2.33
X5 VTAIL.t2 VP.t2 VDD1.t5 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0.9702 ps=6.21 w=5.88 l=2.33
X6 VDD2.t2 VN.t2 VTAIL.t13 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=2.2932 ps=12.54 w=5.88 l=2.33
X7 B.t8 B.t6 B.t7 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0 ps=0 w=5.88 l=2.33
X8 B.t5 B.t3 B.t4 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0 ps=0 w=5.88 l=2.33
X9 VTAIL.t12 VN.t3 VDD2.t6 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X10 VTAIL.t11 VN.t4 VDD2.t0 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0.9702 ps=6.21 w=5.88 l=2.33
X11 VDD1.t4 VP.t3 VTAIL.t7 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=2.2932 ps=12.54 w=5.88 l=2.33
X12 B.t2 B.t0 B.t1 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0 ps=0 w=5.88 l=2.33
X13 VTAIL.t10 VN.t5 VDD2.t7 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X14 VDD2.t1 VN.t6 VTAIL.t9 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X15 VTAIL.t1 VP.t4 VDD1.t3 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X16 VTAIL.t3 VP.t5 VDD1.t2 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=2.2932 pd=12.54 as=0.9702 ps=6.21 w=5.88 l=2.33
X17 VDD1.t1 VP.t6 VTAIL.t6 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X18 VDD2.t5 VN.t7 VTAIL.t8 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
X19 VTAIL.t5 VP.t7 VDD1.t0 w_n3630_n2144# sky130_fd_pr__pfet_01v8 ad=0.9702 pd=6.21 as=0.9702 ps=6.21 w=5.88 l=2.33
R0 VN.n51 VN.n27 161.3
R1 VN.n50 VN.n49 161.3
R2 VN.n48 VN.n28 161.3
R3 VN.n47 VN.n46 161.3
R4 VN.n45 VN.n29 161.3
R5 VN.n43 VN.n42 161.3
R6 VN.n41 VN.n30 161.3
R7 VN.n40 VN.n39 161.3
R8 VN.n38 VN.n31 161.3
R9 VN.n37 VN.n36 161.3
R10 VN.n35 VN.n32 161.3
R11 VN.n24 VN.n0 161.3
R12 VN.n23 VN.n22 161.3
R13 VN.n21 VN.n1 161.3
R14 VN.n20 VN.n19 161.3
R15 VN.n18 VN.n2 161.3
R16 VN.n16 VN.n15 161.3
R17 VN.n14 VN.n3 161.3
R18 VN.n13 VN.n12 161.3
R19 VN.n11 VN.n4 161.3
R20 VN.n10 VN.n9 161.3
R21 VN.n8 VN.n5 161.3
R22 VN.n26 VN.n25 99.1042
R23 VN.n53 VN.n52 99.1042
R24 VN.n7 VN.t4 92.3904
R25 VN.n34 VN.t2 92.3904
R26 VN.n7 VN.n6 68.4787
R27 VN.n34 VN.n33 68.4787
R28 VN.n6 VN.t6 60.8194
R29 VN.n17 VN.t5 60.8194
R30 VN.n25 VN.t1 60.8194
R31 VN.n33 VN.t3 60.8194
R32 VN.n44 VN.t7 60.8194
R33 VN.n52 VN.t0 60.8194
R34 VN.n12 VN.n11 56.5617
R35 VN.n39 VN.n38 56.5617
R36 VN.n19 VN.n1 49.296
R37 VN.n46 VN.n28 49.296
R38 VN VN.n53 45.2558
R39 VN.n23 VN.n1 31.8581
R40 VN.n50 VN.n28 31.8581
R41 VN.n10 VN.n5 24.5923
R42 VN.n11 VN.n10 24.5923
R43 VN.n12 VN.n3 24.5923
R44 VN.n16 VN.n3 24.5923
R45 VN.n19 VN.n18 24.5923
R46 VN.n24 VN.n23 24.5923
R47 VN.n38 VN.n37 24.5923
R48 VN.n37 VN.n32 24.5923
R49 VN.n46 VN.n45 24.5923
R50 VN.n43 VN.n30 24.5923
R51 VN.n39 VN.n30 24.5923
R52 VN.n51 VN.n50 24.5923
R53 VN.n18 VN.n17 20.6576
R54 VN.n45 VN.n44 20.6576
R55 VN.n25 VN.n24 11.8046
R56 VN.n52 VN.n51 11.8046
R57 VN.n35 VN.n34 9.81118
R58 VN.n8 VN.n7 9.81118
R59 VN.n6 VN.n5 3.93519
R60 VN.n17 VN.n16 3.93519
R61 VN.n33 VN.n32 3.93519
R62 VN.n44 VN.n43 3.93519
R63 VN.n53 VN.n27 0.278335
R64 VN.n26 VN.n0 0.278335
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n42 VN.n29 0.189894
R70 VN.n42 VN.n41 0.189894
R71 VN.n41 VN.n40 0.189894
R72 VN.n40 VN.n31 0.189894
R73 VN.n36 VN.n31 0.189894
R74 VN.n36 VN.n35 0.189894
R75 VN.n9 VN.n8 0.189894
R76 VN.n9 VN.n4 0.189894
R77 VN.n13 VN.n4 0.189894
R78 VN.n14 VN.n13 0.189894
R79 VN.n15 VN.n14 0.189894
R80 VN.n15 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153485
R86 VDD2.n2 VDD2.n1 91.058
R87 VDD2.n2 VDD2.n0 91.058
R88 VDD2 VDD2.n5 91.0552
R89 VDD2.n4 VDD2.n3 89.967
R90 VDD2.n4 VDD2.n2 39.1032
R91 VDD2.n5 VDD2.t6 5.52856
R92 VDD2.n5 VDD2.t2 5.52856
R93 VDD2.n3 VDD2.t4 5.52856
R94 VDD2.n3 VDD2.t5 5.52856
R95 VDD2.n1 VDD2.t7 5.52856
R96 VDD2.n1 VDD2.t3 5.52856
R97 VDD2.n0 VDD2.t0 5.52856
R98 VDD2.n0 VDD2.t1 5.52856
R99 VDD2 VDD2.n4 1.20524
R100 VTAIL.n258 VTAIL.n232 756.745
R101 VTAIL.n28 VTAIL.n2 756.745
R102 VTAIL.n60 VTAIL.n34 756.745
R103 VTAIL.n94 VTAIL.n68 756.745
R104 VTAIL.n226 VTAIL.n200 756.745
R105 VTAIL.n192 VTAIL.n166 756.745
R106 VTAIL.n160 VTAIL.n134 756.745
R107 VTAIL.n126 VTAIL.n100 756.745
R108 VTAIL.n243 VTAIL.n242 585
R109 VTAIL.n240 VTAIL.n239 585
R110 VTAIL.n249 VTAIL.n248 585
R111 VTAIL.n251 VTAIL.n250 585
R112 VTAIL.n236 VTAIL.n235 585
R113 VTAIL.n257 VTAIL.n256 585
R114 VTAIL.n259 VTAIL.n258 585
R115 VTAIL.n13 VTAIL.n12 585
R116 VTAIL.n10 VTAIL.n9 585
R117 VTAIL.n19 VTAIL.n18 585
R118 VTAIL.n21 VTAIL.n20 585
R119 VTAIL.n6 VTAIL.n5 585
R120 VTAIL.n27 VTAIL.n26 585
R121 VTAIL.n29 VTAIL.n28 585
R122 VTAIL.n45 VTAIL.n44 585
R123 VTAIL.n42 VTAIL.n41 585
R124 VTAIL.n51 VTAIL.n50 585
R125 VTAIL.n53 VTAIL.n52 585
R126 VTAIL.n38 VTAIL.n37 585
R127 VTAIL.n59 VTAIL.n58 585
R128 VTAIL.n61 VTAIL.n60 585
R129 VTAIL.n79 VTAIL.n78 585
R130 VTAIL.n76 VTAIL.n75 585
R131 VTAIL.n85 VTAIL.n84 585
R132 VTAIL.n87 VTAIL.n86 585
R133 VTAIL.n72 VTAIL.n71 585
R134 VTAIL.n93 VTAIL.n92 585
R135 VTAIL.n95 VTAIL.n94 585
R136 VTAIL.n227 VTAIL.n226 585
R137 VTAIL.n225 VTAIL.n224 585
R138 VTAIL.n204 VTAIL.n203 585
R139 VTAIL.n219 VTAIL.n218 585
R140 VTAIL.n217 VTAIL.n216 585
R141 VTAIL.n208 VTAIL.n207 585
R142 VTAIL.n211 VTAIL.n210 585
R143 VTAIL.n193 VTAIL.n192 585
R144 VTAIL.n191 VTAIL.n190 585
R145 VTAIL.n170 VTAIL.n169 585
R146 VTAIL.n185 VTAIL.n184 585
R147 VTAIL.n183 VTAIL.n182 585
R148 VTAIL.n174 VTAIL.n173 585
R149 VTAIL.n177 VTAIL.n176 585
R150 VTAIL.n161 VTAIL.n160 585
R151 VTAIL.n159 VTAIL.n158 585
R152 VTAIL.n138 VTAIL.n137 585
R153 VTAIL.n153 VTAIL.n152 585
R154 VTAIL.n151 VTAIL.n150 585
R155 VTAIL.n142 VTAIL.n141 585
R156 VTAIL.n145 VTAIL.n144 585
R157 VTAIL.n127 VTAIL.n126 585
R158 VTAIL.n125 VTAIL.n124 585
R159 VTAIL.n104 VTAIL.n103 585
R160 VTAIL.n119 VTAIL.n118 585
R161 VTAIL.n117 VTAIL.n116 585
R162 VTAIL.n108 VTAIL.n107 585
R163 VTAIL.n111 VTAIL.n110 585
R164 VTAIL.t14 VTAIL.n241 327.601
R165 VTAIL.t11 VTAIL.n11 327.601
R166 VTAIL.t7 VTAIL.n43 327.601
R167 VTAIL.t2 VTAIL.n77 327.601
R168 VTAIL.t0 VTAIL.n209 327.601
R169 VTAIL.t3 VTAIL.n175 327.601
R170 VTAIL.t13 VTAIL.n143 327.601
R171 VTAIL.t15 VTAIL.n109 327.601
R172 VTAIL.n242 VTAIL.n239 171.744
R173 VTAIL.n249 VTAIL.n239 171.744
R174 VTAIL.n250 VTAIL.n249 171.744
R175 VTAIL.n250 VTAIL.n235 171.744
R176 VTAIL.n257 VTAIL.n235 171.744
R177 VTAIL.n258 VTAIL.n257 171.744
R178 VTAIL.n12 VTAIL.n9 171.744
R179 VTAIL.n19 VTAIL.n9 171.744
R180 VTAIL.n20 VTAIL.n19 171.744
R181 VTAIL.n20 VTAIL.n5 171.744
R182 VTAIL.n27 VTAIL.n5 171.744
R183 VTAIL.n28 VTAIL.n27 171.744
R184 VTAIL.n44 VTAIL.n41 171.744
R185 VTAIL.n51 VTAIL.n41 171.744
R186 VTAIL.n52 VTAIL.n51 171.744
R187 VTAIL.n52 VTAIL.n37 171.744
R188 VTAIL.n59 VTAIL.n37 171.744
R189 VTAIL.n60 VTAIL.n59 171.744
R190 VTAIL.n78 VTAIL.n75 171.744
R191 VTAIL.n85 VTAIL.n75 171.744
R192 VTAIL.n86 VTAIL.n85 171.744
R193 VTAIL.n86 VTAIL.n71 171.744
R194 VTAIL.n93 VTAIL.n71 171.744
R195 VTAIL.n94 VTAIL.n93 171.744
R196 VTAIL.n226 VTAIL.n225 171.744
R197 VTAIL.n225 VTAIL.n203 171.744
R198 VTAIL.n218 VTAIL.n203 171.744
R199 VTAIL.n218 VTAIL.n217 171.744
R200 VTAIL.n217 VTAIL.n207 171.744
R201 VTAIL.n210 VTAIL.n207 171.744
R202 VTAIL.n192 VTAIL.n191 171.744
R203 VTAIL.n191 VTAIL.n169 171.744
R204 VTAIL.n184 VTAIL.n169 171.744
R205 VTAIL.n184 VTAIL.n183 171.744
R206 VTAIL.n183 VTAIL.n173 171.744
R207 VTAIL.n176 VTAIL.n173 171.744
R208 VTAIL.n160 VTAIL.n159 171.744
R209 VTAIL.n159 VTAIL.n137 171.744
R210 VTAIL.n152 VTAIL.n137 171.744
R211 VTAIL.n152 VTAIL.n151 171.744
R212 VTAIL.n151 VTAIL.n141 171.744
R213 VTAIL.n144 VTAIL.n141 171.744
R214 VTAIL.n126 VTAIL.n125 171.744
R215 VTAIL.n125 VTAIL.n103 171.744
R216 VTAIL.n118 VTAIL.n103 171.744
R217 VTAIL.n118 VTAIL.n117 171.744
R218 VTAIL.n117 VTAIL.n107 171.744
R219 VTAIL.n110 VTAIL.n107 171.744
R220 VTAIL.n242 VTAIL.t14 85.8723
R221 VTAIL.n12 VTAIL.t11 85.8723
R222 VTAIL.n44 VTAIL.t7 85.8723
R223 VTAIL.n78 VTAIL.t2 85.8723
R224 VTAIL.n210 VTAIL.t0 85.8723
R225 VTAIL.n176 VTAIL.t3 85.8723
R226 VTAIL.n144 VTAIL.t13 85.8723
R227 VTAIL.n110 VTAIL.t15 85.8723
R228 VTAIL.n199 VTAIL.n198 73.2882
R229 VTAIL.n133 VTAIL.n132 73.2882
R230 VTAIL.n1 VTAIL.n0 73.288
R231 VTAIL.n67 VTAIL.n66 73.288
R232 VTAIL.n263 VTAIL.n262 29.8581
R233 VTAIL.n33 VTAIL.n32 29.8581
R234 VTAIL.n65 VTAIL.n64 29.8581
R235 VTAIL.n99 VTAIL.n98 29.8581
R236 VTAIL.n231 VTAIL.n230 29.8581
R237 VTAIL.n197 VTAIL.n196 29.8581
R238 VTAIL.n165 VTAIL.n164 29.8581
R239 VTAIL.n131 VTAIL.n130 29.8581
R240 VTAIL.n263 VTAIL.n231 19.7289
R241 VTAIL.n131 VTAIL.n99 19.7289
R242 VTAIL.n243 VTAIL.n241 16.3865
R243 VTAIL.n13 VTAIL.n11 16.3865
R244 VTAIL.n45 VTAIL.n43 16.3865
R245 VTAIL.n79 VTAIL.n77 16.3865
R246 VTAIL.n211 VTAIL.n209 16.3865
R247 VTAIL.n177 VTAIL.n175 16.3865
R248 VTAIL.n145 VTAIL.n143 16.3865
R249 VTAIL.n111 VTAIL.n109 16.3865
R250 VTAIL.n244 VTAIL.n240 12.8005
R251 VTAIL.n14 VTAIL.n10 12.8005
R252 VTAIL.n46 VTAIL.n42 12.8005
R253 VTAIL.n80 VTAIL.n76 12.8005
R254 VTAIL.n212 VTAIL.n208 12.8005
R255 VTAIL.n178 VTAIL.n174 12.8005
R256 VTAIL.n146 VTAIL.n142 12.8005
R257 VTAIL.n112 VTAIL.n108 12.8005
R258 VTAIL.n248 VTAIL.n247 12.0247
R259 VTAIL.n18 VTAIL.n17 12.0247
R260 VTAIL.n50 VTAIL.n49 12.0247
R261 VTAIL.n84 VTAIL.n83 12.0247
R262 VTAIL.n216 VTAIL.n215 12.0247
R263 VTAIL.n182 VTAIL.n181 12.0247
R264 VTAIL.n150 VTAIL.n149 12.0247
R265 VTAIL.n116 VTAIL.n115 12.0247
R266 VTAIL.n251 VTAIL.n238 11.249
R267 VTAIL.n21 VTAIL.n8 11.249
R268 VTAIL.n53 VTAIL.n40 11.249
R269 VTAIL.n87 VTAIL.n74 11.249
R270 VTAIL.n219 VTAIL.n206 11.249
R271 VTAIL.n185 VTAIL.n172 11.249
R272 VTAIL.n153 VTAIL.n140 11.249
R273 VTAIL.n119 VTAIL.n106 11.249
R274 VTAIL.n252 VTAIL.n236 10.4732
R275 VTAIL.n22 VTAIL.n6 10.4732
R276 VTAIL.n54 VTAIL.n38 10.4732
R277 VTAIL.n88 VTAIL.n72 10.4732
R278 VTAIL.n220 VTAIL.n204 10.4732
R279 VTAIL.n186 VTAIL.n170 10.4732
R280 VTAIL.n154 VTAIL.n138 10.4732
R281 VTAIL.n120 VTAIL.n104 10.4732
R282 VTAIL.n256 VTAIL.n255 9.69747
R283 VTAIL.n26 VTAIL.n25 9.69747
R284 VTAIL.n58 VTAIL.n57 9.69747
R285 VTAIL.n92 VTAIL.n91 9.69747
R286 VTAIL.n224 VTAIL.n223 9.69747
R287 VTAIL.n190 VTAIL.n189 9.69747
R288 VTAIL.n158 VTAIL.n157 9.69747
R289 VTAIL.n124 VTAIL.n123 9.69747
R290 VTAIL.n262 VTAIL.n261 9.45567
R291 VTAIL.n32 VTAIL.n31 9.45567
R292 VTAIL.n64 VTAIL.n63 9.45567
R293 VTAIL.n98 VTAIL.n97 9.45567
R294 VTAIL.n230 VTAIL.n229 9.45567
R295 VTAIL.n196 VTAIL.n195 9.45567
R296 VTAIL.n164 VTAIL.n163 9.45567
R297 VTAIL.n130 VTAIL.n129 9.45567
R298 VTAIL.n261 VTAIL.n260 9.3005
R299 VTAIL.n234 VTAIL.n233 9.3005
R300 VTAIL.n255 VTAIL.n254 9.3005
R301 VTAIL.n253 VTAIL.n252 9.3005
R302 VTAIL.n238 VTAIL.n237 9.3005
R303 VTAIL.n247 VTAIL.n246 9.3005
R304 VTAIL.n245 VTAIL.n244 9.3005
R305 VTAIL.n31 VTAIL.n30 9.3005
R306 VTAIL.n4 VTAIL.n3 9.3005
R307 VTAIL.n25 VTAIL.n24 9.3005
R308 VTAIL.n23 VTAIL.n22 9.3005
R309 VTAIL.n8 VTAIL.n7 9.3005
R310 VTAIL.n17 VTAIL.n16 9.3005
R311 VTAIL.n15 VTAIL.n14 9.3005
R312 VTAIL.n63 VTAIL.n62 9.3005
R313 VTAIL.n36 VTAIL.n35 9.3005
R314 VTAIL.n57 VTAIL.n56 9.3005
R315 VTAIL.n55 VTAIL.n54 9.3005
R316 VTAIL.n40 VTAIL.n39 9.3005
R317 VTAIL.n49 VTAIL.n48 9.3005
R318 VTAIL.n47 VTAIL.n46 9.3005
R319 VTAIL.n97 VTAIL.n96 9.3005
R320 VTAIL.n70 VTAIL.n69 9.3005
R321 VTAIL.n91 VTAIL.n90 9.3005
R322 VTAIL.n89 VTAIL.n88 9.3005
R323 VTAIL.n74 VTAIL.n73 9.3005
R324 VTAIL.n83 VTAIL.n82 9.3005
R325 VTAIL.n81 VTAIL.n80 9.3005
R326 VTAIL.n229 VTAIL.n228 9.3005
R327 VTAIL.n202 VTAIL.n201 9.3005
R328 VTAIL.n223 VTAIL.n222 9.3005
R329 VTAIL.n221 VTAIL.n220 9.3005
R330 VTAIL.n206 VTAIL.n205 9.3005
R331 VTAIL.n215 VTAIL.n214 9.3005
R332 VTAIL.n213 VTAIL.n212 9.3005
R333 VTAIL.n195 VTAIL.n194 9.3005
R334 VTAIL.n168 VTAIL.n167 9.3005
R335 VTAIL.n189 VTAIL.n188 9.3005
R336 VTAIL.n187 VTAIL.n186 9.3005
R337 VTAIL.n172 VTAIL.n171 9.3005
R338 VTAIL.n181 VTAIL.n180 9.3005
R339 VTAIL.n179 VTAIL.n178 9.3005
R340 VTAIL.n163 VTAIL.n162 9.3005
R341 VTAIL.n136 VTAIL.n135 9.3005
R342 VTAIL.n157 VTAIL.n156 9.3005
R343 VTAIL.n155 VTAIL.n154 9.3005
R344 VTAIL.n140 VTAIL.n139 9.3005
R345 VTAIL.n149 VTAIL.n148 9.3005
R346 VTAIL.n147 VTAIL.n146 9.3005
R347 VTAIL.n129 VTAIL.n128 9.3005
R348 VTAIL.n102 VTAIL.n101 9.3005
R349 VTAIL.n123 VTAIL.n122 9.3005
R350 VTAIL.n121 VTAIL.n120 9.3005
R351 VTAIL.n106 VTAIL.n105 9.3005
R352 VTAIL.n115 VTAIL.n114 9.3005
R353 VTAIL.n113 VTAIL.n112 9.3005
R354 VTAIL.n259 VTAIL.n234 8.92171
R355 VTAIL.n29 VTAIL.n4 8.92171
R356 VTAIL.n61 VTAIL.n36 8.92171
R357 VTAIL.n95 VTAIL.n70 8.92171
R358 VTAIL.n227 VTAIL.n202 8.92171
R359 VTAIL.n193 VTAIL.n168 8.92171
R360 VTAIL.n161 VTAIL.n136 8.92171
R361 VTAIL.n127 VTAIL.n102 8.92171
R362 VTAIL.n260 VTAIL.n232 8.14595
R363 VTAIL.n30 VTAIL.n2 8.14595
R364 VTAIL.n62 VTAIL.n34 8.14595
R365 VTAIL.n96 VTAIL.n68 8.14595
R366 VTAIL.n228 VTAIL.n200 8.14595
R367 VTAIL.n194 VTAIL.n166 8.14595
R368 VTAIL.n162 VTAIL.n134 8.14595
R369 VTAIL.n128 VTAIL.n100 8.14595
R370 VTAIL.n262 VTAIL.n232 5.81868
R371 VTAIL.n32 VTAIL.n2 5.81868
R372 VTAIL.n64 VTAIL.n34 5.81868
R373 VTAIL.n98 VTAIL.n68 5.81868
R374 VTAIL.n230 VTAIL.n200 5.81868
R375 VTAIL.n196 VTAIL.n166 5.81868
R376 VTAIL.n164 VTAIL.n134 5.81868
R377 VTAIL.n130 VTAIL.n100 5.81868
R378 VTAIL.n0 VTAIL.t9 5.52856
R379 VTAIL.n0 VTAIL.t10 5.52856
R380 VTAIL.n66 VTAIL.t4 5.52856
R381 VTAIL.n66 VTAIL.t1 5.52856
R382 VTAIL.n198 VTAIL.t6 5.52856
R383 VTAIL.n198 VTAIL.t5 5.52856
R384 VTAIL.n132 VTAIL.t8 5.52856
R385 VTAIL.n132 VTAIL.t12 5.52856
R386 VTAIL.n260 VTAIL.n259 5.04292
R387 VTAIL.n30 VTAIL.n29 5.04292
R388 VTAIL.n62 VTAIL.n61 5.04292
R389 VTAIL.n96 VTAIL.n95 5.04292
R390 VTAIL.n228 VTAIL.n227 5.04292
R391 VTAIL.n194 VTAIL.n193 5.04292
R392 VTAIL.n162 VTAIL.n161 5.04292
R393 VTAIL.n128 VTAIL.n127 5.04292
R394 VTAIL.n256 VTAIL.n234 4.26717
R395 VTAIL.n26 VTAIL.n4 4.26717
R396 VTAIL.n58 VTAIL.n36 4.26717
R397 VTAIL.n92 VTAIL.n70 4.26717
R398 VTAIL.n224 VTAIL.n202 4.26717
R399 VTAIL.n190 VTAIL.n168 4.26717
R400 VTAIL.n158 VTAIL.n136 4.26717
R401 VTAIL.n124 VTAIL.n102 4.26717
R402 VTAIL.n213 VTAIL.n209 3.71286
R403 VTAIL.n179 VTAIL.n175 3.71286
R404 VTAIL.n147 VTAIL.n143 3.71286
R405 VTAIL.n113 VTAIL.n109 3.71286
R406 VTAIL.n245 VTAIL.n241 3.71286
R407 VTAIL.n15 VTAIL.n11 3.71286
R408 VTAIL.n47 VTAIL.n43 3.71286
R409 VTAIL.n81 VTAIL.n77 3.71286
R410 VTAIL.n255 VTAIL.n236 3.49141
R411 VTAIL.n25 VTAIL.n6 3.49141
R412 VTAIL.n57 VTAIL.n38 3.49141
R413 VTAIL.n91 VTAIL.n72 3.49141
R414 VTAIL.n223 VTAIL.n204 3.49141
R415 VTAIL.n189 VTAIL.n170 3.49141
R416 VTAIL.n157 VTAIL.n138 3.49141
R417 VTAIL.n123 VTAIL.n104 3.49141
R418 VTAIL.n252 VTAIL.n251 2.71565
R419 VTAIL.n22 VTAIL.n21 2.71565
R420 VTAIL.n54 VTAIL.n53 2.71565
R421 VTAIL.n88 VTAIL.n87 2.71565
R422 VTAIL.n220 VTAIL.n219 2.71565
R423 VTAIL.n186 VTAIL.n185 2.71565
R424 VTAIL.n154 VTAIL.n153 2.71565
R425 VTAIL.n120 VTAIL.n119 2.71565
R426 VTAIL.n133 VTAIL.n131 2.2936
R427 VTAIL.n165 VTAIL.n133 2.2936
R428 VTAIL.n199 VTAIL.n197 2.2936
R429 VTAIL.n231 VTAIL.n199 2.2936
R430 VTAIL.n99 VTAIL.n67 2.2936
R431 VTAIL.n67 VTAIL.n65 2.2936
R432 VTAIL.n33 VTAIL.n1 2.2936
R433 VTAIL VTAIL.n263 2.23541
R434 VTAIL.n248 VTAIL.n238 1.93989
R435 VTAIL.n18 VTAIL.n8 1.93989
R436 VTAIL.n50 VTAIL.n40 1.93989
R437 VTAIL.n84 VTAIL.n74 1.93989
R438 VTAIL.n216 VTAIL.n206 1.93989
R439 VTAIL.n182 VTAIL.n172 1.93989
R440 VTAIL.n150 VTAIL.n140 1.93989
R441 VTAIL.n116 VTAIL.n106 1.93989
R442 VTAIL.n247 VTAIL.n240 1.16414
R443 VTAIL.n17 VTAIL.n10 1.16414
R444 VTAIL.n49 VTAIL.n42 1.16414
R445 VTAIL.n83 VTAIL.n76 1.16414
R446 VTAIL.n215 VTAIL.n208 1.16414
R447 VTAIL.n181 VTAIL.n174 1.16414
R448 VTAIL.n149 VTAIL.n142 1.16414
R449 VTAIL.n115 VTAIL.n108 1.16414
R450 VTAIL.n197 VTAIL.n165 0.470328
R451 VTAIL.n65 VTAIL.n33 0.470328
R452 VTAIL.n244 VTAIL.n243 0.388379
R453 VTAIL.n14 VTAIL.n13 0.388379
R454 VTAIL.n46 VTAIL.n45 0.388379
R455 VTAIL.n80 VTAIL.n79 0.388379
R456 VTAIL.n212 VTAIL.n211 0.388379
R457 VTAIL.n178 VTAIL.n177 0.388379
R458 VTAIL.n146 VTAIL.n145 0.388379
R459 VTAIL.n112 VTAIL.n111 0.388379
R460 VTAIL.n246 VTAIL.n245 0.155672
R461 VTAIL.n246 VTAIL.n237 0.155672
R462 VTAIL.n253 VTAIL.n237 0.155672
R463 VTAIL.n254 VTAIL.n253 0.155672
R464 VTAIL.n254 VTAIL.n233 0.155672
R465 VTAIL.n261 VTAIL.n233 0.155672
R466 VTAIL.n16 VTAIL.n15 0.155672
R467 VTAIL.n16 VTAIL.n7 0.155672
R468 VTAIL.n23 VTAIL.n7 0.155672
R469 VTAIL.n24 VTAIL.n23 0.155672
R470 VTAIL.n24 VTAIL.n3 0.155672
R471 VTAIL.n31 VTAIL.n3 0.155672
R472 VTAIL.n48 VTAIL.n47 0.155672
R473 VTAIL.n48 VTAIL.n39 0.155672
R474 VTAIL.n55 VTAIL.n39 0.155672
R475 VTAIL.n56 VTAIL.n55 0.155672
R476 VTAIL.n56 VTAIL.n35 0.155672
R477 VTAIL.n63 VTAIL.n35 0.155672
R478 VTAIL.n82 VTAIL.n81 0.155672
R479 VTAIL.n82 VTAIL.n73 0.155672
R480 VTAIL.n89 VTAIL.n73 0.155672
R481 VTAIL.n90 VTAIL.n89 0.155672
R482 VTAIL.n90 VTAIL.n69 0.155672
R483 VTAIL.n97 VTAIL.n69 0.155672
R484 VTAIL.n229 VTAIL.n201 0.155672
R485 VTAIL.n222 VTAIL.n201 0.155672
R486 VTAIL.n222 VTAIL.n221 0.155672
R487 VTAIL.n221 VTAIL.n205 0.155672
R488 VTAIL.n214 VTAIL.n205 0.155672
R489 VTAIL.n214 VTAIL.n213 0.155672
R490 VTAIL.n195 VTAIL.n167 0.155672
R491 VTAIL.n188 VTAIL.n167 0.155672
R492 VTAIL.n188 VTAIL.n187 0.155672
R493 VTAIL.n187 VTAIL.n171 0.155672
R494 VTAIL.n180 VTAIL.n171 0.155672
R495 VTAIL.n180 VTAIL.n179 0.155672
R496 VTAIL.n163 VTAIL.n135 0.155672
R497 VTAIL.n156 VTAIL.n135 0.155672
R498 VTAIL.n156 VTAIL.n155 0.155672
R499 VTAIL.n155 VTAIL.n139 0.155672
R500 VTAIL.n148 VTAIL.n139 0.155672
R501 VTAIL.n148 VTAIL.n147 0.155672
R502 VTAIL.n129 VTAIL.n101 0.155672
R503 VTAIL.n122 VTAIL.n101 0.155672
R504 VTAIL.n122 VTAIL.n121 0.155672
R505 VTAIL.n121 VTAIL.n105 0.155672
R506 VTAIL.n114 VTAIL.n105 0.155672
R507 VTAIL.n114 VTAIL.n113 0.155672
R508 VTAIL VTAIL.n1 0.0586897
R509 VP.n16 VP.n13 161.3
R510 VP.n18 VP.n17 161.3
R511 VP.n19 VP.n12 161.3
R512 VP.n21 VP.n20 161.3
R513 VP.n22 VP.n11 161.3
R514 VP.n24 VP.n23 161.3
R515 VP.n26 VP.n10 161.3
R516 VP.n28 VP.n27 161.3
R517 VP.n29 VP.n9 161.3
R518 VP.n31 VP.n30 161.3
R519 VP.n32 VP.n8 161.3
R520 VP.n62 VP.n0 161.3
R521 VP.n61 VP.n60 161.3
R522 VP.n59 VP.n1 161.3
R523 VP.n58 VP.n57 161.3
R524 VP.n56 VP.n2 161.3
R525 VP.n54 VP.n53 161.3
R526 VP.n52 VP.n3 161.3
R527 VP.n51 VP.n50 161.3
R528 VP.n49 VP.n4 161.3
R529 VP.n48 VP.n47 161.3
R530 VP.n46 VP.n5 161.3
R531 VP.n45 VP.n44 161.3
R532 VP.n42 VP.n6 161.3
R533 VP.n41 VP.n40 161.3
R534 VP.n39 VP.n7 161.3
R535 VP.n38 VP.n37 161.3
R536 VP.n36 VP.n35 99.1042
R537 VP.n64 VP.n63 99.1042
R538 VP.n34 VP.n33 99.1042
R539 VP.n15 VP.t5 92.3904
R540 VP.n15 VP.n14 68.4787
R541 VP.n36 VP.t2 60.8194
R542 VP.n43 VP.t1 60.8194
R543 VP.n55 VP.t4 60.8194
R544 VP.n63 VP.t3 60.8194
R545 VP.n33 VP.t0 60.8194
R546 VP.n25 VP.t7 60.8194
R547 VP.n14 VP.t6 60.8194
R548 VP.n50 VP.n49 56.5617
R549 VP.n20 VP.n19 56.5617
R550 VP.n42 VP.n41 49.296
R551 VP.n57 VP.n1 49.296
R552 VP.n27 VP.n9 49.296
R553 VP.n35 VP.n34 44.9769
R554 VP.n41 VP.n7 31.8581
R555 VP.n61 VP.n1 31.8581
R556 VP.n31 VP.n9 31.8581
R557 VP.n37 VP.n7 24.5923
R558 VP.n44 VP.n42 24.5923
R559 VP.n48 VP.n5 24.5923
R560 VP.n49 VP.n48 24.5923
R561 VP.n50 VP.n3 24.5923
R562 VP.n54 VP.n3 24.5923
R563 VP.n57 VP.n56 24.5923
R564 VP.n62 VP.n61 24.5923
R565 VP.n32 VP.n31 24.5923
R566 VP.n20 VP.n11 24.5923
R567 VP.n24 VP.n11 24.5923
R568 VP.n27 VP.n26 24.5923
R569 VP.n18 VP.n13 24.5923
R570 VP.n19 VP.n18 24.5923
R571 VP.n44 VP.n43 20.6576
R572 VP.n56 VP.n55 20.6576
R573 VP.n26 VP.n25 20.6576
R574 VP.n37 VP.n36 11.8046
R575 VP.n63 VP.n62 11.8046
R576 VP.n33 VP.n32 11.8046
R577 VP.n16 VP.n15 9.81118
R578 VP.n43 VP.n5 3.93519
R579 VP.n55 VP.n54 3.93519
R580 VP.n25 VP.n24 3.93519
R581 VP.n14 VP.n13 3.93519
R582 VP.n34 VP.n8 0.278335
R583 VP.n38 VP.n35 0.278335
R584 VP.n64 VP.n0 0.278335
R585 VP.n17 VP.n16 0.189894
R586 VP.n17 VP.n12 0.189894
R587 VP.n21 VP.n12 0.189894
R588 VP.n22 VP.n21 0.189894
R589 VP.n23 VP.n22 0.189894
R590 VP.n23 VP.n10 0.189894
R591 VP.n28 VP.n10 0.189894
R592 VP.n29 VP.n28 0.189894
R593 VP.n30 VP.n29 0.189894
R594 VP.n30 VP.n8 0.189894
R595 VP.n39 VP.n38 0.189894
R596 VP.n40 VP.n39 0.189894
R597 VP.n40 VP.n6 0.189894
R598 VP.n45 VP.n6 0.189894
R599 VP.n46 VP.n45 0.189894
R600 VP.n47 VP.n46 0.189894
R601 VP.n47 VP.n4 0.189894
R602 VP.n51 VP.n4 0.189894
R603 VP.n52 VP.n51 0.189894
R604 VP.n53 VP.n52 0.189894
R605 VP.n53 VP.n2 0.189894
R606 VP.n58 VP.n2 0.189894
R607 VP.n59 VP.n58 0.189894
R608 VP.n60 VP.n59 0.189894
R609 VP.n60 VP.n0 0.189894
R610 VP VP.n64 0.153485
R611 VDD1 VDD1.n0 91.1717
R612 VDD1.n3 VDD1.n2 91.058
R613 VDD1.n3 VDD1.n1 91.058
R614 VDD1.n5 VDD1.n4 89.9668
R615 VDD1.n5 VDD1.n3 39.6862
R616 VDD1.n4 VDD1.t0 5.52856
R617 VDD1.n4 VDD1.t7 5.52856
R618 VDD1.n0 VDD1.t2 5.52856
R619 VDD1.n0 VDD1.t1 5.52856
R620 VDD1.n2 VDD1.t3 5.52856
R621 VDD1.n2 VDD1.t4 5.52856
R622 VDD1.n1 VDD1.t5 5.52856
R623 VDD1.n1 VDD1.t6 5.52856
R624 VDD1 VDD1.n5 1.08886
R625 B.n461 B.n58 585
R626 B.n463 B.n462 585
R627 B.n464 B.n57 585
R628 B.n466 B.n465 585
R629 B.n467 B.n56 585
R630 B.n469 B.n468 585
R631 B.n470 B.n55 585
R632 B.n472 B.n471 585
R633 B.n473 B.n54 585
R634 B.n475 B.n474 585
R635 B.n476 B.n53 585
R636 B.n478 B.n477 585
R637 B.n479 B.n52 585
R638 B.n481 B.n480 585
R639 B.n482 B.n51 585
R640 B.n484 B.n483 585
R641 B.n485 B.n50 585
R642 B.n487 B.n486 585
R643 B.n488 B.n49 585
R644 B.n490 B.n489 585
R645 B.n491 B.n48 585
R646 B.n493 B.n492 585
R647 B.n494 B.n47 585
R648 B.n496 B.n495 585
R649 B.n498 B.n497 585
R650 B.n499 B.n43 585
R651 B.n501 B.n500 585
R652 B.n502 B.n42 585
R653 B.n504 B.n503 585
R654 B.n505 B.n41 585
R655 B.n507 B.n506 585
R656 B.n508 B.n40 585
R657 B.n510 B.n509 585
R658 B.n512 B.n37 585
R659 B.n514 B.n513 585
R660 B.n515 B.n36 585
R661 B.n517 B.n516 585
R662 B.n518 B.n35 585
R663 B.n520 B.n519 585
R664 B.n521 B.n34 585
R665 B.n523 B.n522 585
R666 B.n524 B.n33 585
R667 B.n526 B.n525 585
R668 B.n527 B.n32 585
R669 B.n529 B.n528 585
R670 B.n530 B.n31 585
R671 B.n532 B.n531 585
R672 B.n533 B.n30 585
R673 B.n535 B.n534 585
R674 B.n536 B.n29 585
R675 B.n538 B.n537 585
R676 B.n539 B.n28 585
R677 B.n541 B.n540 585
R678 B.n542 B.n27 585
R679 B.n544 B.n543 585
R680 B.n545 B.n26 585
R681 B.n547 B.n546 585
R682 B.n460 B.n459 585
R683 B.n458 B.n59 585
R684 B.n457 B.n456 585
R685 B.n455 B.n60 585
R686 B.n454 B.n453 585
R687 B.n452 B.n61 585
R688 B.n451 B.n450 585
R689 B.n449 B.n62 585
R690 B.n448 B.n447 585
R691 B.n446 B.n63 585
R692 B.n445 B.n444 585
R693 B.n443 B.n64 585
R694 B.n442 B.n441 585
R695 B.n440 B.n65 585
R696 B.n439 B.n438 585
R697 B.n437 B.n66 585
R698 B.n436 B.n435 585
R699 B.n434 B.n67 585
R700 B.n433 B.n432 585
R701 B.n431 B.n68 585
R702 B.n430 B.n429 585
R703 B.n428 B.n69 585
R704 B.n427 B.n426 585
R705 B.n425 B.n70 585
R706 B.n424 B.n423 585
R707 B.n422 B.n71 585
R708 B.n421 B.n420 585
R709 B.n419 B.n72 585
R710 B.n418 B.n417 585
R711 B.n416 B.n73 585
R712 B.n415 B.n414 585
R713 B.n413 B.n74 585
R714 B.n412 B.n411 585
R715 B.n410 B.n75 585
R716 B.n409 B.n408 585
R717 B.n407 B.n76 585
R718 B.n406 B.n405 585
R719 B.n404 B.n77 585
R720 B.n403 B.n402 585
R721 B.n401 B.n78 585
R722 B.n400 B.n399 585
R723 B.n398 B.n79 585
R724 B.n397 B.n396 585
R725 B.n395 B.n80 585
R726 B.n394 B.n393 585
R727 B.n392 B.n81 585
R728 B.n391 B.n390 585
R729 B.n389 B.n82 585
R730 B.n388 B.n387 585
R731 B.n386 B.n83 585
R732 B.n385 B.n384 585
R733 B.n383 B.n84 585
R734 B.n382 B.n381 585
R735 B.n380 B.n85 585
R736 B.n379 B.n378 585
R737 B.n377 B.n86 585
R738 B.n376 B.n375 585
R739 B.n374 B.n87 585
R740 B.n373 B.n372 585
R741 B.n371 B.n88 585
R742 B.n370 B.n369 585
R743 B.n368 B.n89 585
R744 B.n367 B.n366 585
R745 B.n365 B.n90 585
R746 B.n364 B.n363 585
R747 B.n362 B.n91 585
R748 B.n361 B.n360 585
R749 B.n359 B.n92 585
R750 B.n358 B.n357 585
R751 B.n356 B.n93 585
R752 B.n355 B.n354 585
R753 B.n353 B.n94 585
R754 B.n352 B.n351 585
R755 B.n350 B.n95 585
R756 B.n349 B.n348 585
R757 B.n347 B.n96 585
R758 B.n346 B.n345 585
R759 B.n344 B.n97 585
R760 B.n343 B.n342 585
R761 B.n341 B.n98 585
R762 B.n340 B.n339 585
R763 B.n338 B.n99 585
R764 B.n337 B.n336 585
R765 B.n335 B.n100 585
R766 B.n334 B.n333 585
R767 B.n332 B.n101 585
R768 B.n331 B.n330 585
R769 B.n329 B.n102 585
R770 B.n328 B.n327 585
R771 B.n326 B.n103 585
R772 B.n325 B.n324 585
R773 B.n323 B.n104 585
R774 B.n322 B.n321 585
R775 B.n320 B.n105 585
R776 B.n319 B.n318 585
R777 B.n232 B.n231 585
R778 B.n233 B.n138 585
R779 B.n235 B.n234 585
R780 B.n236 B.n137 585
R781 B.n238 B.n237 585
R782 B.n239 B.n136 585
R783 B.n241 B.n240 585
R784 B.n242 B.n135 585
R785 B.n244 B.n243 585
R786 B.n245 B.n134 585
R787 B.n247 B.n246 585
R788 B.n248 B.n133 585
R789 B.n250 B.n249 585
R790 B.n251 B.n132 585
R791 B.n253 B.n252 585
R792 B.n254 B.n131 585
R793 B.n256 B.n255 585
R794 B.n257 B.n130 585
R795 B.n259 B.n258 585
R796 B.n260 B.n129 585
R797 B.n262 B.n261 585
R798 B.n263 B.n128 585
R799 B.n265 B.n264 585
R800 B.n266 B.n125 585
R801 B.n269 B.n268 585
R802 B.n270 B.n124 585
R803 B.n272 B.n271 585
R804 B.n273 B.n123 585
R805 B.n275 B.n274 585
R806 B.n276 B.n122 585
R807 B.n278 B.n277 585
R808 B.n279 B.n121 585
R809 B.n281 B.n280 585
R810 B.n283 B.n282 585
R811 B.n284 B.n117 585
R812 B.n286 B.n285 585
R813 B.n287 B.n116 585
R814 B.n289 B.n288 585
R815 B.n290 B.n115 585
R816 B.n292 B.n291 585
R817 B.n293 B.n114 585
R818 B.n295 B.n294 585
R819 B.n296 B.n113 585
R820 B.n298 B.n297 585
R821 B.n299 B.n112 585
R822 B.n301 B.n300 585
R823 B.n302 B.n111 585
R824 B.n304 B.n303 585
R825 B.n305 B.n110 585
R826 B.n307 B.n306 585
R827 B.n308 B.n109 585
R828 B.n310 B.n309 585
R829 B.n311 B.n108 585
R830 B.n313 B.n312 585
R831 B.n314 B.n107 585
R832 B.n316 B.n315 585
R833 B.n317 B.n106 585
R834 B.n230 B.n139 585
R835 B.n229 B.n228 585
R836 B.n227 B.n140 585
R837 B.n226 B.n225 585
R838 B.n224 B.n141 585
R839 B.n223 B.n222 585
R840 B.n221 B.n142 585
R841 B.n220 B.n219 585
R842 B.n218 B.n143 585
R843 B.n217 B.n216 585
R844 B.n215 B.n144 585
R845 B.n214 B.n213 585
R846 B.n212 B.n145 585
R847 B.n211 B.n210 585
R848 B.n209 B.n146 585
R849 B.n208 B.n207 585
R850 B.n206 B.n147 585
R851 B.n205 B.n204 585
R852 B.n203 B.n148 585
R853 B.n202 B.n201 585
R854 B.n200 B.n149 585
R855 B.n199 B.n198 585
R856 B.n197 B.n150 585
R857 B.n196 B.n195 585
R858 B.n194 B.n151 585
R859 B.n193 B.n192 585
R860 B.n191 B.n152 585
R861 B.n190 B.n189 585
R862 B.n188 B.n153 585
R863 B.n187 B.n186 585
R864 B.n185 B.n154 585
R865 B.n184 B.n183 585
R866 B.n182 B.n155 585
R867 B.n181 B.n180 585
R868 B.n179 B.n156 585
R869 B.n178 B.n177 585
R870 B.n176 B.n157 585
R871 B.n175 B.n174 585
R872 B.n173 B.n158 585
R873 B.n172 B.n171 585
R874 B.n170 B.n159 585
R875 B.n169 B.n168 585
R876 B.n167 B.n160 585
R877 B.n166 B.n165 585
R878 B.n164 B.n161 585
R879 B.n163 B.n162 585
R880 B.n2 B.n0 585
R881 B.n617 B.n1 585
R882 B.n616 B.n615 585
R883 B.n614 B.n3 585
R884 B.n613 B.n612 585
R885 B.n611 B.n4 585
R886 B.n610 B.n609 585
R887 B.n608 B.n5 585
R888 B.n607 B.n606 585
R889 B.n605 B.n6 585
R890 B.n604 B.n603 585
R891 B.n602 B.n7 585
R892 B.n601 B.n600 585
R893 B.n599 B.n8 585
R894 B.n598 B.n597 585
R895 B.n596 B.n9 585
R896 B.n595 B.n594 585
R897 B.n593 B.n10 585
R898 B.n592 B.n591 585
R899 B.n590 B.n11 585
R900 B.n589 B.n588 585
R901 B.n587 B.n12 585
R902 B.n586 B.n585 585
R903 B.n584 B.n13 585
R904 B.n583 B.n582 585
R905 B.n581 B.n14 585
R906 B.n580 B.n579 585
R907 B.n578 B.n15 585
R908 B.n577 B.n576 585
R909 B.n575 B.n16 585
R910 B.n574 B.n573 585
R911 B.n572 B.n17 585
R912 B.n571 B.n570 585
R913 B.n569 B.n18 585
R914 B.n568 B.n567 585
R915 B.n566 B.n19 585
R916 B.n565 B.n564 585
R917 B.n563 B.n20 585
R918 B.n562 B.n561 585
R919 B.n560 B.n21 585
R920 B.n559 B.n558 585
R921 B.n557 B.n22 585
R922 B.n556 B.n555 585
R923 B.n554 B.n23 585
R924 B.n553 B.n552 585
R925 B.n551 B.n24 585
R926 B.n550 B.n549 585
R927 B.n548 B.n25 585
R928 B.n619 B.n618 585
R929 B.n232 B.n139 521.33
R930 B.n546 B.n25 521.33
R931 B.n318 B.n317 521.33
R932 B.n461 B.n460 521.33
R933 B.n118 B.t5 317.454
R934 B.n44 B.t10 317.454
R935 B.n126 B.t8 317.454
R936 B.n38 B.t1 317.454
R937 B.n118 B.t3 268.418
R938 B.n126 B.t6 268.418
R939 B.n38 B.t0 268.418
R940 B.n44 B.t9 268.418
R941 B.n119 B.t4 265.865
R942 B.n45 B.t11 265.865
R943 B.n127 B.t7 265.865
R944 B.n39 B.t2 265.865
R945 B.n228 B.n139 163.367
R946 B.n228 B.n227 163.367
R947 B.n227 B.n226 163.367
R948 B.n226 B.n141 163.367
R949 B.n222 B.n141 163.367
R950 B.n222 B.n221 163.367
R951 B.n221 B.n220 163.367
R952 B.n220 B.n143 163.367
R953 B.n216 B.n143 163.367
R954 B.n216 B.n215 163.367
R955 B.n215 B.n214 163.367
R956 B.n214 B.n145 163.367
R957 B.n210 B.n145 163.367
R958 B.n210 B.n209 163.367
R959 B.n209 B.n208 163.367
R960 B.n208 B.n147 163.367
R961 B.n204 B.n147 163.367
R962 B.n204 B.n203 163.367
R963 B.n203 B.n202 163.367
R964 B.n202 B.n149 163.367
R965 B.n198 B.n149 163.367
R966 B.n198 B.n197 163.367
R967 B.n197 B.n196 163.367
R968 B.n196 B.n151 163.367
R969 B.n192 B.n151 163.367
R970 B.n192 B.n191 163.367
R971 B.n191 B.n190 163.367
R972 B.n190 B.n153 163.367
R973 B.n186 B.n153 163.367
R974 B.n186 B.n185 163.367
R975 B.n185 B.n184 163.367
R976 B.n184 B.n155 163.367
R977 B.n180 B.n155 163.367
R978 B.n180 B.n179 163.367
R979 B.n179 B.n178 163.367
R980 B.n178 B.n157 163.367
R981 B.n174 B.n157 163.367
R982 B.n174 B.n173 163.367
R983 B.n173 B.n172 163.367
R984 B.n172 B.n159 163.367
R985 B.n168 B.n159 163.367
R986 B.n168 B.n167 163.367
R987 B.n167 B.n166 163.367
R988 B.n166 B.n161 163.367
R989 B.n162 B.n161 163.367
R990 B.n162 B.n2 163.367
R991 B.n618 B.n2 163.367
R992 B.n618 B.n617 163.367
R993 B.n617 B.n616 163.367
R994 B.n616 B.n3 163.367
R995 B.n612 B.n3 163.367
R996 B.n612 B.n611 163.367
R997 B.n611 B.n610 163.367
R998 B.n610 B.n5 163.367
R999 B.n606 B.n5 163.367
R1000 B.n606 B.n605 163.367
R1001 B.n605 B.n604 163.367
R1002 B.n604 B.n7 163.367
R1003 B.n600 B.n7 163.367
R1004 B.n600 B.n599 163.367
R1005 B.n599 B.n598 163.367
R1006 B.n598 B.n9 163.367
R1007 B.n594 B.n9 163.367
R1008 B.n594 B.n593 163.367
R1009 B.n593 B.n592 163.367
R1010 B.n592 B.n11 163.367
R1011 B.n588 B.n11 163.367
R1012 B.n588 B.n587 163.367
R1013 B.n587 B.n586 163.367
R1014 B.n586 B.n13 163.367
R1015 B.n582 B.n13 163.367
R1016 B.n582 B.n581 163.367
R1017 B.n581 B.n580 163.367
R1018 B.n580 B.n15 163.367
R1019 B.n576 B.n15 163.367
R1020 B.n576 B.n575 163.367
R1021 B.n575 B.n574 163.367
R1022 B.n574 B.n17 163.367
R1023 B.n570 B.n17 163.367
R1024 B.n570 B.n569 163.367
R1025 B.n569 B.n568 163.367
R1026 B.n568 B.n19 163.367
R1027 B.n564 B.n19 163.367
R1028 B.n564 B.n563 163.367
R1029 B.n563 B.n562 163.367
R1030 B.n562 B.n21 163.367
R1031 B.n558 B.n21 163.367
R1032 B.n558 B.n557 163.367
R1033 B.n557 B.n556 163.367
R1034 B.n556 B.n23 163.367
R1035 B.n552 B.n23 163.367
R1036 B.n552 B.n551 163.367
R1037 B.n551 B.n550 163.367
R1038 B.n550 B.n25 163.367
R1039 B.n233 B.n232 163.367
R1040 B.n234 B.n233 163.367
R1041 B.n234 B.n137 163.367
R1042 B.n238 B.n137 163.367
R1043 B.n239 B.n238 163.367
R1044 B.n240 B.n239 163.367
R1045 B.n240 B.n135 163.367
R1046 B.n244 B.n135 163.367
R1047 B.n245 B.n244 163.367
R1048 B.n246 B.n245 163.367
R1049 B.n246 B.n133 163.367
R1050 B.n250 B.n133 163.367
R1051 B.n251 B.n250 163.367
R1052 B.n252 B.n251 163.367
R1053 B.n252 B.n131 163.367
R1054 B.n256 B.n131 163.367
R1055 B.n257 B.n256 163.367
R1056 B.n258 B.n257 163.367
R1057 B.n258 B.n129 163.367
R1058 B.n262 B.n129 163.367
R1059 B.n263 B.n262 163.367
R1060 B.n264 B.n263 163.367
R1061 B.n264 B.n125 163.367
R1062 B.n269 B.n125 163.367
R1063 B.n270 B.n269 163.367
R1064 B.n271 B.n270 163.367
R1065 B.n271 B.n123 163.367
R1066 B.n275 B.n123 163.367
R1067 B.n276 B.n275 163.367
R1068 B.n277 B.n276 163.367
R1069 B.n277 B.n121 163.367
R1070 B.n281 B.n121 163.367
R1071 B.n282 B.n281 163.367
R1072 B.n282 B.n117 163.367
R1073 B.n286 B.n117 163.367
R1074 B.n287 B.n286 163.367
R1075 B.n288 B.n287 163.367
R1076 B.n288 B.n115 163.367
R1077 B.n292 B.n115 163.367
R1078 B.n293 B.n292 163.367
R1079 B.n294 B.n293 163.367
R1080 B.n294 B.n113 163.367
R1081 B.n298 B.n113 163.367
R1082 B.n299 B.n298 163.367
R1083 B.n300 B.n299 163.367
R1084 B.n300 B.n111 163.367
R1085 B.n304 B.n111 163.367
R1086 B.n305 B.n304 163.367
R1087 B.n306 B.n305 163.367
R1088 B.n306 B.n109 163.367
R1089 B.n310 B.n109 163.367
R1090 B.n311 B.n310 163.367
R1091 B.n312 B.n311 163.367
R1092 B.n312 B.n107 163.367
R1093 B.n316 B.n107 163.367
R1094 B.n317 B.n316 163.367
R1095 B.n318 B.n105 163.367
R1096 B.n322 B.n105 163.367
R1097 B.n323 B.n322 163.367
R1098 B.n324 B.n323 163.367
R1099 B.n324 B.n103 163.367
R1100 B.n328 B.n103 163.367
R1101 B.n329 B.n328 163.367
R1102 B.n330 B.n329 163.367
R1103 B.n330 B.n101 163.367
R1104 B.n334 B.n101 163.367
R1105 B.n335 B.n334 163.367
R1106 B.n336 B.n335 163.367
R1107 B.n336 B.n99 163.367
R1108 B.n340 B.n99 163.367
R1109 B.n341 B.n340 163.367
R1110 B.n342 B.n341 163.367
R1111 B.n342 B.n97 163.367
R1112 B.n346 B.n97 163.367
R1113 B.n347 B.n346 163.367
R1114 B.n348 B.n347 163.367
R1115 B.n348 B.n95 163.367
R1116 B.n352 B.n95 163.367
R1117 B.n353 B.n352 163.367
R1118 B.n354 B.n353 163.367
R1119 B.n354 B.n93 163.367
R1120 B.n358 B.n93 163.367
R1121 B.n359 B.n358 163.367
R1122 B.n360 B.n359 163.367
R1123 B.n360 B.n91 163.367
R1124 B.n364 B.n91 163.367
R1125 B.n365 B.n364 163.367
R1126 B.n366 B.n365 163.367
R1127 B.n366 B.n89 163.367
R1128 B.n370 B.n89 163.367
R1129 B.n371 B.n370 163.367
R1130 B.n372 B.n371 163.367
R1131 B.n372 B.n87 163.367
R1132 B.n376 B.n87 163.367
R1133 B.n377 B.n376 163.367
R1134 B.n378 B.n377 163.367
R1135 B.n378 B.n85 163.367
R1136 B.n382 B.n85 163.367
R1137 B.n383 B.n382 163.367
R1138 B.n384 B.n383 163.367
R1139 B.n384 B.n83 163.367
R1140 B.n388 B.n83 163.367
R1141 B.n389 B.n388 163.367
R1142 B.n390 B.n389 163.367
R1143 B.n390 B.n81 163.367
R1144 B.n394 B.n81 163.367
R1145 B.n395 B.n394 163.367
R1146 B.n396 B.n395 163.367
R1147 B.n396 B.n79 163.367
R1148 B.n400 B.n79 163.367
R1149 B.n401 B.n400 163.367
R1150 B.n402 B.n401 163.367
R1151 B.n402 B.n77 163.367
R1152 B.n406 B.n77 163.367
R1153 B.n407 B.n406 163.367
R1154 B.n408 B.n407 163.367
R1155 B.n408 B.n75 163.367
R1156 B.n412 B.n75 163.367
R1157 B.n413 B.n412 163.367
R1158 B.n414 B.n413 163.367
R1159 B.n414 B.n73 163.367
R1160 B.n418 B.n73 163.367
R1161 B.n419 B.n418 163.367
R1162 B.n420 B.n419 163.367
R1163 B.n420 B.n71 163.367
R1164 B.n424 B.n71 163.367
R1165 B.n425 B.n424 163.367
R1166 B.n426 B.n425 163.367
R1167 B.n426 B.n69 163.367
R1168 B.n430 B.n69 163.367
R1169 B.n431 B.n430 163.367
R1170 B.n432 B.n431 163.367
R1171 B.n432 B.n67 163.367
R1172 B.n436 B.n67 163.367
R1173 B.n437 B.n436 163.367
R1174 B.n438 B.n437 163.367
R1175 B.n438 B.n65 163.367
R1176 B.n442 B.n65 163.367
R1177 B.n443 B.n442 163.367
R1178 B.n444 B.n443 163.367
R1179 B.n444 B.n63 163.367
R1180 B.n448 B.n63 163.367
R1181 B.n449 B.n448 163.367
R1182 B.n450 B.n449 163.367
R1183 B.n450 B.n61 163.367
R1184 B.n454 B.n61 163.367
R1185 B.n455 B.n454 163.367
R1186 B.n456 B.n455 163.367
R1187 B.n456 B.n59 163.367
R1188 B.n460 B.n59 163.367
R1189 B.n546 B.n545 163.367
R1190 B.n545 B.n544 163.367
R1191 B.n544 B.n27 163.367
R1192 B.n540 B.n27 163.367
R1193 B.n540 B.n539 163.367
R1194 B.n539 B.n538 163.367
R1195 B.n538 B.n29 163.367
R1196 B.n534 B.n29 163.367
R1197 B.n534 B.n533 163.367
R1198 B.n533 B.n532 163.367
R1199 B.n532 B.n31 163.367
R1200 B.n528 B.n31 163.367
R1201 B.n528 B.n527 163.367
R1202 B.n527 B.n526 163.367
R1203 B.n526 B.n33 163.367
R1204 B.n522 B.n33 163.367
R1205 B.n522 B.n521 163.367
R1206 B.n521 B.n520 163.367
R1207 B.n520 B.n35 163.367
R1208 B.n516 B.n35 163.367
R1209 B.n516 B.n515 163.367
R1210 B.n515 B.n514 163.367
R1211 B.n514 B.n37 163.367
R1212 B.n509 B.n37 163.367
R1213 B.n509 B.n508 163.367
R1214 B.n508 B.n507 163.367
R1215 B.n507 B.n41 163.367
R1216 B.n503 B.n41 163.367
R1217 B.n503 B.n502 163.367
R1218 B.n502 B.n501 163.367
R1219 B.n501 B.n43 163.367
R1220 B.n497 B.n43 163.367
R1221 B.n497 B.n496 163.367
R1222 B.n496 B.n47 163.367
R1223 B.n492 B.n47 163.367
R1224 B.n492 B.n491 163.367
R1225 B.n491 B.n490 163.367
R1226 B.n490 B.n49 163.367
R1227 B.n486 B.n49 163.367
R1228 B.n486 B.n485 163.367
R1229 B.n485 B.n484 163.367
R1230 B.n484 B.n51 163.367
R1231 B.n480 B.n51 163.367
R1232 B.n480 B.n479 163.367
R1233 B.n479 B.n478 163.367
R1234 B.n478 B.n53 163.367
R1235 B.n474 B.n53 163.367
R1236 B.n474 B.n473 163.367
R1237 B.n473 B.n472 163.367
R1238 B.n472 B.n55 163.367
R1239 B.n468 B.n55 163.367
R1240 B.n468 B.n467 163.367
R1241 B.n467 B.n466 163.367
R1242 B.n466 B.n57 163.367
R1243 B.n462 B.n57 163.367
R1244 B.n462 B.n461 163.367
R1245 B.n120 B.n119 59.5399
R1246 B.n267 B.n127 59.5399
R1247 B.n511 B.n39 59.5399
R1248 B.n46 B.n45 59.5399
R1249 B.n119 B.n118 51.5884
R1250 B.n127 B.n126 51.5884
R1251 B.n39 B.n38 51.5884
R1252 B.n45 B.n44 51.5884
R1253 B.n548 B.n547 33.8737
R1254 B.n459 B.n58 33.8737
R1255 B.n319 B.n106 33.8737
R1256 B.n231 B.n230 33.8737
R1257 B B.n619 18.0485
R1258 B.n547 B.n26 10.6151
R1259 B.n543 B.n26 10.6151
R1260 B.n543 B.n542 10.6151
R1261 B.n542 B.n541 10.6151
R1262 B.n541 B.n28 10.6151
R1263 B.n537 B.n28 10.6151
R1264 B.n537 B.n536 10.6151
R1265 B.n536 B.n535 10.6151
R1266 B.n535 B.n30 10.6151
R1267 B.n531 B.n30 10.6151
R1268 B.n531 B.n530 10.6151
R1269 B.n530 B.n529 10.6151
R1270 B.n529 B.n32 10.6151
R1271 B.n525 B.n32 10.6151
R1272 B.n525 B.n524 10.6151
R1273 B.n524 B.n523 10.6151
R1274 B.n523 B.n34 10.6151
R1275 B.n519 B.n34 10.6151
R1276 B.n519 B.n518 10.6151
R1277 B.n518 B.n517 10.6151
R1278 B.n517 B.n36 10.6151
R1279 B.n513 B.n36 10.6151
R1280 B.n513 B.n512 10.6151
R1281 B.n510 B.n40 10.6151
R1282 B.n506 B.n40 10.6151
R1283 B.n506 B.n505 10.6151
R1284 B.n505 B.n504 10.6151
R1285 B.n504 B.n42 10.6151
R1286 B.n500 B.n42 10.6151
R1287 B.n500 B.n499 10.6151
R1288 B.n499 B.n498 10.6151
R1289 B.n495 B.n494 10.6151
R1290 B.n494 B.n493 10.6151
R1291 B.n493 B.n48 10.6151
R1292 B.n489 B.n48 10.6151
R1293 B.n489 B.n488 10.6151
R1294 B.n488 B.n487 10.6151
R1295 B.n487 B.n50 10.6151
R1296 B.n483 B.n50 10.6151
R1297 B.n483 B.n482 10.6151
R1298 B.n482 B.n481 10.6151
R1299 B.n481 B.n52 10.6151
R1300 B.n477 B.n52 10.6151
R1301 B.n477 B.n476 10.6151
R1302 B.n476 B.n475 10.6151
R1303 B.n475 B.n54 10.6151
R1304 B.n471 B.n54 10.6151
R1305 B.n471 B.n470 10.6151
R1306 B.n470 B.n469 10.6151
R1307 B.n469 B.n56 10.6151
R1308 B.n465 B.n56 10.6151
R1309 B.n465 B.n464 10.6151
R1310 B.n464 B.n463 10.6151
R1311 B.n463 B.n58 10.6151
R1312 B.n320 B.n319 10.6151
R1313 B.n321 B.n320 10.6151
R1314 B.n321 B.n104 10.6151
R1315 B.n325 B.n104 10.6151
R1316 B.n326 B.n325 10.6151
R1317 B.n327 B.n326 10.6151
R1318 B.n327 B.n102 10.6151
R1319 B.n331 B.n102 10.6151
R1320 B.n332 B.n331 10.6151
R1321 B.n333 B.n332 10.6151
R1322 B.n333 B.n100 10.6151
R1323 B.n337 B.n100 10.6151
R1324 B.n338 B.n337 10.6151
R1325 B.n339 B.n338 10.6151
R1326 B.n339 B.n98 10.6151
R1327 B.n343 B.n98 10.6151
R1328 B.n344 B.n343 10.6151
R1329 B.n345 B.n344 10.6151
R1330 B.n345 B.n96 10.6151
R1331 B.n349 B.n96 10.6151
R1332 B.n350 B.n349 10.6151
R1333 B.n351 B.n350 10.6151
R1334 B.n351 B.n94 10.6151
R1335 B.n355 B.n94 10.6151
R1336 B.n356 B.n355 10.6151
R1337 B.n357 B.n356 10.6151
R1338 B.n357 B.n92 10.6151
R1339 B.n361 B.n92 10.6151
R1340 B.n362 B.n361 10.6151
R1341 B.n363 B.n362 10.6151
R1342 B.n363 B.n90 10.6151
R1343 B.n367 B.n90 10.6151
R1344 B.n368 B.n367 10.6151
R1345 B.n369 B.n368 10.6151
R1346 B.n369 B.n88 10.6151
R1347 B.n373 B.n88 10.6151
R1348 B.n374 B.n373 10.6151
R1349 B.n375 B.n374 10.6151
R1350 B.n375 B.n86 10.6151
R1351 B.n379 B.n86 10.6151
R1352 B.n380 B.n379 10.6151
R1353 B.n381 B.n380 10.6151
R1354 B.n381 B.n84 10.6151
R1355 B.n385 B.n84 10.6151
R1356 B.n386 B.n385 10.6151
R1357 B.n387 B.n386 10.6151
R1358 B.n387 B.n82 10.6151
R1359 B.n391 B.n82 10.6151
R1360 B.n392 B.n391 10.6151
R1361 B.n393 B.n392 10.6151
R1362 B.n393 B.n80 10.6151
R1363 B.n397 B.n80 10.6151
R1364 B.n398 B.n397 10.6151
R1365 B.n399 B.n398 10.6151
R1366 B.n399 B.n78 10.6151
R1367 B.n403 B.n78 10.6151
R1368 B.n404 B.n403 10.6151
R1369 B.n405 B.n404 10.6151
R1370 B.n405 B.n76 10.6151
R1371 B.n409 B.n76 10.6151
R1372 B.n410 B.n409 10.6151
R1373 B.n411 B.n410 10.6151
R1374 B.n411 B.n74 10.6151
R1375 B.n415 B.n74 10.6151
R1376 B.n416 B.n415 10.6151
R1377 B.n417 B.n416 10.6151
R1378 B.n417 B.n72 10.6151
R1379 B.n421 B.n72 10.6151
R1380 B.n422 B.n421 10.6151
R1381 B.n423 B.n422 10.6151
R1382 B.n423 B.n70 10.6151
R1383 B.n427 B.n70 10.6151
R1384 B.n428 B.n427 10.6151
R1385 B.n429 B.n428 10.6151
R1386 B.n429 B.n68 10.6151
R1387 B.n433 B.n68 10.6151
R1388 B.n434 B.n433 10.6151
R1389 B.n435 B.n434 10.6151
R1390 B.n435 B.n66 10.6151
R1391 B.n439 B.n66 10.6151
R1392 B.n440 B.n439 10.6151
R1393 B.n441 B.n440 10.6151
R1394 B.n441 B.n64 10.6151
R1395 B.n445 B.n64 10.6151
R1396 B.n446 B.n445 10.6151
R1397 B.n447 B.n446 10.6151
R1398 B.n447 B.n62 10.6151
R1399 B.n451 B.n62 10.6151
R1400 B.n452 B.n451 10.6151
R1401 B.n453 B.n452 10.6151
R1402 B.n453 B.n60 10.6151
R1403 B.n457 B.n60 10.6151
R1404 B.n458 B.n457 10.6151
R1405 B.n459 B.n458 10.6151
R1406 B.n231 B.n138 10.6151
R1407 B.n235 B.n138 10.6151
R1408 B.n236 B.n235 10.6151
R1409 B.n237 B.n236 10.6151
R1410 B.n237 B.n136 10.6151
R1411 B.n241 B.n136 10.6151
R1412 B.n242 B.n241 10.6151
R1413 B.n243 B.n242 10.6151
R1414 B.n243 B.n134 10.6151
R1415 B.n247 B.n134 10.6151
R1416 B.n248 B.n247 10.6151
R1417 B.n249 B.n248 10.6151
R1418 B.n249 B.n132 10.6151
R1419 B.n253 B.n132 10.6151
R1420 B.n254 B.n253 10.6151
R1421 B.n255 B.n254 10.6151
R1422 B.n255 B.n130 10.6151
R1423 B.n259 B.n130 10.6151
R1424 B.n260 B.n259 10.6151
R1425 B.n261 B.n260 10.6151
R1426 B.n261 B.n128 10.6151
R1427 B.n265 B.n128 10.6151
R1428 B.n266 B.n265 10.6151
R1429 B.n268 B.n124 10.6151
R1430 B.n272 B.n124 10.6151
R1431 B.n273 B.n272 10.6151
R1432 B.n274 B.n273 10.6151
R1433 B.n274 B.n122 10.6151
R1434 B.n278 B.n122 10.6151
R1435 B.n279 B.n278 10.6151
R1436 B.n280 B.n279 10.6151
R1437 B.n284 B.n283 10.6151
R1438 B.n285 B.n284 10.6151
R1439 B.n285 B.n116 10.6151
R1440 B.n289 B.n116 10.6151
R1441 B.n290 B.n289 10.6151
R1442 B.n291 B.n290 10.6151
R1443 B.n291 B.n114 10.6151
R1444 B.n295 B.n114 10.6151
R1445 B.n296 B.n295 10.6151
R1446 B.n297 B.n296 10.6151
R1447 B.n297 B.n112 10.6151
R1448 B.n301 B.n112 10.6151
R1449 B.n302 B.n301 10.6151
R1450 B.n303 B.n302 10.6151
R1451 B.n303 B.n110 10.6151
R1452 B.n307 B.n110 10.6151
R1453 B.n308 B.n307 10.6151
R1454 B.n309 B.n308 10.6151
R1455 B.n309 B.n108 10.6151
R1456 B.n313 B.n108 10.6151
R1457 B.n314 B.n313 10.6151
R1458 B.n315 B.n314 10.6151
R1459 B.n315 B.n106 10.6151
R1460 B.n230 B.n229 10.6151
R1461 B.n229 B.n140 10.6151
R1462 B.n225 B.n140 10.6151
R1463 B.n225 B.n224 10.6151
R1464 B.n224 B.n223 10.6151
R1465 B.n223 B.n142 10.6151
R1466 B.n219 B.n142 10.6151
R1467 B.n219 B.n218 10.6151
R1468 B.n218 B.n217 10.6151
R1469 B.n217 B.n144 10.6151
R1470 B.n213 B.n144 10.6151
R1471 B.n213 B.n212 10.6151
R1472 B.n212 B.n211 10.6151
R1473 B.n211 B.n146 10.6151
R1474 B.n207 B.n146 10.6151
R1475 B.n207 B.n206 10.6151
R1476 B.n206 B.n205 10.6151
R1477 B.n205 B.n148 10.6151
R1478 B.n201 B.n148 10.6151
R1479 B.n201 B.n200 10.6151
R1480 B.n200 B.n199 10.6151
R1481 B.n199 B.n150 10.6151
R1482 B.n195 B.n150 10.6151
R1483 B.n195 B.n194 10.6151
R1484 B.n194 B.n193 10.6151
R1485 B.n193 B.n152 10.6151
R1486 B.n189 B.n152 10.6151
R1487 B.n189 B.n188 10.6151
R1488 B.n188 B.n187 10.6151
R1489 B.n187 B.n154 10.6151
R1490 B.n183 B.n154 10.6151
R1491 B.n183 B.n182 10.6151
R1492 B.n182 B.n181 10.6151
R1493 B.n181 B.n156 10.6151
R1494 B.n177 B.n156 10.6151
R1495 B.n177 B.n176 10.6151
R1496 B.n176 B.n175 10.6151
R1497 B.n175 B.n158 10.6151
R1498 B.n171 B.n158 10.6151
R1499 B.n171 B.n170 10.6151
R1500 B.n170 B.n169 10.6151
R1501 B.n169 B.n160 10.6151
R1502 B.n165 B.n160 10.6151
R1503 B.n165 B.n164 10.6151
R1504 B.n164 B.n163 10.6151
R1505 B.n163 B.n0 10.6151
R1506 B.n615 B.n1 10.6151
R1507 B.n615 B.n614 10.6151
R1508 B.n614 B.n613 10.6151
R1509 B.n613 B.n4 10.6151
R1510 B.n609 B.n4 10.6151
R1511 B.n609 B.n608 10.6151
R1512 B.n608 B.n607 10.6151
R1513 B.n607 B.n6 10.6151
R1514 B.n603 B.n6 10.6151
R1515 B.n603 B.n602 10.6151
R1516 B.n602 B.n601 10.6151
R1517 B.n601 B.n8 10.6151
R1518 B.n597 B.n8 10.6151
R1519 B.n597 B.n596 10.6151
R1520 B.n596 B.n595 10.6151
R1521 B.n595 B.n10 10.6151
R1522 B.n591 B.n10 10.6151
R1523 B.n591 B.n590 10.6151
R1524 B.n590 B.n589 10.6151
R1525 B.n589 B.n12 10.6151
R1526 B.n585 B.n12 10.6151
R1527 B.n585 B.n584 10.6151
R1528 B.n584 B.n583 10.6151
R1529 B.n583 B.n14 10.6151
R1530 B.n579 B.n14 10.6151
R1531 B.n579 B.n578 10.6151
R1532 B.n578 B.n577 10.6151
R1533 B.n577 B.n16 10.6151
R1534 B.n573 B.n16 10.6151
R1535 B.n573 B.n572 10.6151
R1536 B.n572 B.n571 10.6151
R1537 B.n571 B.n18 10.6151
R1538 B.n567 B.n18 10.6151
R1539 B.n567 B.n566 10.6151
R1540 B.n566 B.n565 10.6151
R1541 B.n565 B.n20 10.6151
R1542 B.n561 B.n20 10.6151
R1543 B.n561 B.n560 10.6151
R1544 B.n560 B.n559 10.6151
R1545 B.n559 B.n22 10.6151
R1546 B.n555 B.n22 10.6151
R1547 B.n555 B.n554 10.6151
R1548 B.n554 B.n553 10.6151
R1549 B.n553 B.n24 10.6151
R1550 B.n549 B.n24 10.6151
R1551 B.n549 B.n548 10.6151
R1552 B.n511 B.n510 6.5566
R1553 B.n498 B.n46 6.5566
R1554 B.n268 B.n267 6.5566
R1555 B.n280 B.n120 6.5566
R1556 B.n512 B.n511 4.05904
R1557 B.n495 B.n46 4.05904
R1558 B.n267 B.n266 4.05904
R1559 B.n283 B.n120 4.05904
R1560 B.n619 B.n0 2.81026
R1561 B.n619 B.n1 2.81026
C0 VTAIL VP 5.13643f
C1 VDD1 VP 4.73356f
C2 VN B 1.08944f
C3 VDD2 VP 0.491087f
C4 VP w_n3630_n2144# 7.668681f
C5 VDD1 VTAIL 5.86537f
C6 VDD2 VTAIL 5.91798f
C7 VTAIL w_n3630_n2144# 2.8014f
C8 VN VP 6.19544f
C9 VDD1 VDD2 1.63558f
C10 VDD1 w_n3630_n2144# 1.70016f
C11 VDD2 w_n3630_n2144# 1.80354f
C12 VN VTAIL 5.12233f
C13 VDD1 VN 0.151387f
C14 B VP 1.87665f
C15 VN VDD2 4.39512f
C16 VN w_n3630_n2144# 7.19823f
C17 B VTAIL 2.87099f
C18 VDD1 B 1.40353f
C19 B VDD2 1.49108f
C20 B w_n3630_n2144# 7.996991f
C21 VDD2 VSUBS 1.506669f
C22 VDD1 VSUBS 2.115237f
C23 VTAIL VSUBS 0.681104f
C24 VN VSUBS 6.114861f
C25 VP VSUBS 2.911975f
C26 B VSUBS 4.181421f
C27 w_n3630_n2144# VSUBS 97.1824f
C28 B.n0 VSUBS 0.005232f
C29 B.n1 VSUBS 0.005232f
C30 B.n2 VSUBS 0.008274f
C31 B.n3 VSUBS 0.008274f
C32 B.n4 VSUBS 0.008274f
C33 B.n5 VSUBS 0.008274f
C34 B.n6 VSUBS 0.008274f
C35 B.n7 VSUBS 0.008274f
C36 B.n8 VSUBS 0.008274f
C37 B.n9 VSUBS 0.008274f
C38 B.n10 VSUBS 0.008274f
C39 B.n11 VSUBS 0.008274f
C40 B.n12 VSUBS 0.008274f
C41 B.n13 VSUBS 0.008274f
C42 B.n14 VSUBS 0.008274f
C43 B.n15 VSUBS 0.008274f
C44 B.n16 VSUBS 0.008274f
C45 B.n17 VSUBS 0.008274f
C46 B.n18 VSUBS 0.008274f
C47 B.n19 VSUBS 0.008274f
C48 B.n20 VSUBS 0.008274f
C49 B.n21 VSUBS 0.008274f
C50 B.n22 VSUBS 0.008274f
C51 B.n23 VSUBS 0.008274f
C52 B.n24 VSUBS 0.008274f
C53 B.n25 VSUBS 0.019132f
C54 B.n26 VSUBS 0.008274f
C55 B.n27 VSUBS 0.008274f
C56 B.n28 VSUBS 0.008274f
C57 B.n29 VSUBS 0.008274f
C58 B.n30 VSUBS 0.008274f
C59 B.n31 VSUBS 0.008274f
C60 B.n32 VSUBS 0.008274f
C61 B.n33 VSUBS 0.008274f
C62 B.n34 VSUBS 0.008274f
C63 B.n35 VSUBS 0.008274f
C64 B.n36 VSUBS 0.008274f
C65 B.n37 VSUBS 0.008274f
C66 B.t2 VSUBS 0.103031f
C67 B.t1 VSUBS 0.130561f
C68 B.t0 VSUBS 0.762458f
C69 B.n38 VSUBS 0.225113f
C70 B.n39 VSUBS 0.181207f
C71 B.n40 VSUBS 0.008274f
C72 B.n41 VSUBS 0.008274f
C73 B.n42 VSUBS 0.008274f
C74 B.n43 VSUBS 0.008274f
C75 B.t11 VSUBS 0.103033f
C76 B.t10 VSUBS 0.130562f
C77 B.t9 VSUBS 0.762458f
C78 B.n44 VSUBS 0.225111f
C79 B.n45 VSUBS 0.181205f
C80 B.n46 VSUBS 0.01917f
C81 B.n47 VSUBS 0.008274f
C82 B.n48 VSUBS 0.008274f
C83 B.n49 VSUBS 0.008274f
C84 B.n50 VSUBS 0.008274f
C85 B.n51 VSUBS 0.008274f
C86 B.n52 VSUBS 0.008274f
C87 B.n53 VSUBS 0.008274f
C88 B.n54 VSUBS 0.008274f
C89 B.n55 VSUBS 0.008274f
C90 B.n56 VSUBS 0.008274f
C91 B.n57 VSUBS 0.008274f
C92 B.n58 VSUBS 0.019592f
C93 B.n59 VSUBS 0.008274f
C94 B.n60 VSUBS 0.008274f
C95 B.n61 VSUBS 0.008274f
C96 B.n62 VSUBS 0.008274f
C97 B.n63 VSUBS 0.008274f
C98 B.n64 VSUBS 0.008274f
C99 B.n65 VSUBS 0.008274f
C100 B.n66 VSUBS 0.008274f
C101 B.n67 VSUBS 0.008274f
C102 B.n68 VSUBS 0.008274f
C103 B.n69 VSUBS 0.008274f
C104 B.n70 VSUBS 0.008274f
C105 B.n71 VSUBS 0.008274f
C106 B.n72 VSUBS 0.008274f
C107 B.n73 VSUBS 0.008274f
C108 B.n74 VSUBS 0.008274f
C109 B.n75 VSUBS 0.008274f
C110 B.n76 VSUBS 0.008274f
C111 B.n77 VSUBS 0.008274f
C112 B.n78 VSUBS 0.008274f
C113 B.n79 VSUBS 0.008274f
C114 B.n80 VSUBS 0.008274f
C115 B.n81 VSUBS 0.008274f
C116 B.n82 VSUBS 0.008274f
C117 B.n83 VSUBS 0.008274f
C118 B.n84 VSUBS 0.008274f
C119 B.n85 VSUBS 0.008274f
C120 B.n86 VSUBS 0.008274f
C121 B.n87 VSUBS 0.008274f
C122 B.n88 VSUBS 0.008274f
C123 B.n89 VSUBS 0.008274f
C124 B.n90 VSUBS 0.008274f
C125 B.n91 VSUBS 0.008274f
C126 B.n92 VSUBS 0.008274f
C127 B.n93 VSUBS 0.008274f
C128 B.n94 VSUBS 0.008274f
C129 B.n95 VSUBS 0.008274f
C130 B.n96 VSUBS 0.008274f
C131 B.n97 VSUBS 0.008274f
C132 B.n98 VSUBS 0.008274f
C133 B.n99 VSUBS 0.008274f
C134 B.n100 VSUBS 0.008274f
C135 B.n101 VSUBS 0.008274f
C136 B.n102 VSUBS 0.008274f
C137 B.n103 VSUBS 0.008274f
C138 B.n104 VSUBS 0.008274f
C139 B.n105 VSUBS 0.008274f
C140 B.n106 VSUBS 0.020535f
C141 B.n107 VSUBS 0.008274f
C142 B.n108 VSUBS 0.008274f
C143 B.n109 VSUBS 0.008274f
C144 B.n110 VSUBS 0.008274f
C145 B.n111 VSUBS 0.008274f
C146 B.n112 VSUBS 0.008274f
C147 B.n113 VSUBS 0.008274f
C148 B.n114 VSUBS 0.008274f
C149 B.n115 VSUBS 0.008274f
C150 B.n116 VSUBS 0.008274f
C151 B.n117 VSUBS 0.008274f
C152 B.t4 VSUBS 0.103033f
C153 B.t5 VSUBS 0.130562f
C154 B.t3 VSUBS 0.762458f
C155 B.n118 VSUBS 0.225111f
C156 B.n119 VSUBS 0.181205f
C157 B.n120 VSUBS 0.01917f
C158 B.n121 VSUBS 0.008274f
C159 B.n122 VSUBS 0.008274f
C160 B.n123 VSUBS 0.008274f
C161 B.n124 VSUBS 0.008274f
C162 B.n125 VSUBS 0.008274f
C163 B.t7 VSUBS 0.103031f
C164 B.t8 VSUBS 0.130561f
C165 B.t6 VSUBS 0.762458f
C166 B.n126 VSUBS 0.225113f
C167 B.n127 VSUBS 0.181207f
C168 B.n128 VSUBS 0.008274f
C169 B.n129 VSUBS 0.008274f
C170 B.n130 VSUBS 0.008274f
C171 B.n131 VSUBS 0.008274f
C172 B.n132 VSUBS 0.008274f
C173 B.n133 VSUBS 0.008274f
C174 B.n134 VSUBS 0.008274f
C175 B.n135 VSUBS 0.008274f
C176 B.n136 VSUBS 0.008274f
C177 B.n137 VSUBS 0.008274f
C178 B.n138 VSUBS 0.008274f
C179 B.n139 VSUBS 0.019132f
C180 B.n140 VSUBS 0.008274f
C181 B.n141 VSUBS 0.008274f
C182 B.n142 VSUBS 0.008274f
C183 B.n143 VSUBS 0.008274f
C184 B.n144 VSUBS 0.008274f
C185 B.n145 VSUBS 0.008274f
C186 B.n146 VSUBS 0.008274f
C187 B.n147 VSUBS 0.008274f
C188 B.n148 VSUBS 0.008274f
C189 B.n149 VSUBS 0.008274f
C190 B.n150 VSUBS 0.008274f
C191 B.n151 VSUBS 0.008274f
C192 B.n152 VSUBS 0.008274f
C193 B.n153 VSUBS 0.008274f
C194 B.n154 VSUBS 0.008274f
C195 B.n155 VSUBS 0.008274f
C196 B.n156 VSUBS 0.008274f
C197 B.n157 VSUBS 0.008274f
C198 B.n158 VSUBS 0.008274f
C199 B.n159 VSUBS 0.008274f
C200 B.n160 VSUBS 0.008274f
C201 B.n161 VSUBS 0.008274f
C202 B.n162 VSUBS 0.008274f
C203 B.n163 VSUBS 0.008274f
C204 B.n164 VSUBS 0.008274f
C205 B.n165 VSUBS 0.008274f
C206 B.n166 VSUBS 0.008274f
C207 B.n167 VSUBS 0.008274f
C208 B.n168 VSUBS 0.008274f
C209 B.n169 VSUBS 0.008274f
C210 B.n170 VSUBS 0.008274f
C211 B.n171 VSUBS 0.008274f
C212 B.n172 VSUBS 0.008274f
C213 B.n173 VSUBS 0.008274f
C214 B.n174 VSUBS 0.008274f
C215 B.n175 VSUBS 0.008274f
C216 B.n176 VSUBS 0.008274f
C217 B.n177 VSUBS 0.008274f
C218 B.n178 VSUBS 0.008274f
C219 B.n179 VSUBS 0.008274f
C220 B.n180 VSUBS 0.008274f
C221 B.n181 VSUBS 0.008274f
C222 B.n182 VSUBS 0.008274f
C223 B.n183 VSUBS 0.008274f
C224 B.n184 VSUBS 0.008274f
C225 B.n185 VSUBS 0.008274f
C226 B.n186 VSUBS 0.008274f
C227 B.n187 VSUBS 0.008274f
C228 B.n188 VSUBS 0.008274f
C229 B.n189 VSUBS 0.008274f
C230 B.n190 VSUBS 0.008274f
C231 B.n191 VSUBS 0.008274f
C232 B.n192 VSUBS 0.008274f
C233 B.n193 VSUBS 0.008274f
C234 B.n194 VSUBS 0.008274f
C235 B.n195 VSUBS 0.008274f
C236 B.n196 VSUBS 0.008274f
C237 B.n197 VSUBS 0.008274f
C238 B.n198 VSUBS 0.008274f
C239 B.n199 VSUBS 0.008274f
C240 B.n200 VSUBS 0.008274f
C241 B.n201 VSUBS 0.008274f
C242 B.n202 VSUBS 0.008274f
C243 B.n203 VSUBS 0.008274f
C244 B.n204 VSUBS 0.008274f
C245 B.n205 VSUBS 0.008274f
C246 B.n206 VSUBS 0.008274f
C247 B.n207 VSUBS 0.008274f
C248 B.n208 VSUBS 0.008274f
C249 B.n209 VSUBS 0.008274f
C250 B.n210 VSUBS 0.008274f
C251 B.n211 VSUBS 0.008274f
C252 B.n212 VSUBS 0.008274f
C253 B.n213 VSUBS 0.008274f
C254 B.n214 VSUBS 0.008274f
C255 B.n215 VSUBS 0.008274f
C256 B.n216 VSUBS 0.008274f
C257 B.n217 VSUBS 0.008274f
C258 B.n218 VSUBS 0.008274f
C259 B.n219 VSUBS 0.008274f
C260 B.n220 VSUBS 0.008274f
C261 B.n221 VSUBS 0.008274f
C262 B.n222 VSUBS 0.008274f
C263 B.n223 VSUBS 0.008274f
C264 B.n224 VSUBS 0.008274f
C265 B.n225 VSUBS 0.008274f
C266 B.n226 VSUBS 0.008274f
C267 B.n227 VSUBS 0.008274f
C268 B.n228 VSUBS 0.008274f
C269 B.n229 VSUBS 0.008274f
C270 B.n230 VSUBS 0.019132f
C271 B.n231 VSUBS 0.020535f
C272 B.n232 VSUBS 0.020535f
C273 B.n233 VSUBS 0.008274f
C274 B.n234 VSUBS 0.008274f
C275 B.n235 VSUBS 0.008274f
C276 B.n236 VSUBS 0.008274f
C277 B.n237 VSUBS 0.008274f
C278 B.n238 VSUBS 0.008274f
C279 B.n239 VSUBS 0.008274f
C280 B.n240 VSUBS 0.008274f
C281 B.n241 VSUBS 0.008274f
C282 B.n242 VSUBS 0.008274f
C283 B.n243 VSUBS 0.008274f
C284 B.n244 VSUBS 0.008274f
C285 B.n245 VSUBS 0.008274f
C286 B.n246 VSUBS 0.008274f
C287 B.n247 VSUBS 0.008274f
C288 B.n248 VSUBS 0.008274f
C289 B.n249 VSUBS 0.008274f
C290 B.n250 VSUBS 0.008274f
C291 B.n251 VSUBS 0.008274f
C292 B.n252 VSUBS 0.008274f
C293 B.n253 VSUBS 0.008274f
C294 B.n254 VSUBS 0.008274f
C295 B.n255 VSUBS 0.008274f
C296 B.n256 VSUBS 0.008274f
C297 B.n257 VSUBS 0.008274f
C298 B.n258 VSUBS 0.008274f
C299 B.n259 VSUBS 0.008274f
C300 B.n260 VSUBS 0.008274f
C301 B.n261 VSUBS 0.008274f
C302 B.n262 VSUBS 0.008274f
C303 B.n263 VSUBS 0.008274f
C304 B.n264 VSUBS 0.008274f
C305 B.n265 VSUBS 0.008274f
C306 B.n266 VSUBS 0.005719f
C307 B.n267 VSUBS 0.01917f
C308 B.n268 VSUBS 0.006692f
C309 B.n269 VSUBS 0.008274f
C310 B.n270 VSUBS 0.008274f
C311 B.n271 VSUBS 0.008274f
C312 B.n272 VSUBS 0.008274f
C313 B.n273 VSUBS 0.008274f
C314 B.n274 VSUBS 0.008274f
C315 B.n275 VSUBS 0.008274f
C316 B.n276 VSUBS 0.008274f
C317 B.n277 VSUBS 0.008274f
C318 B.n278 VSUBS 0.008274f
C319 B.n279 VSUBS 0.008274f
C320 B.n280 VSUBS 0.006692f
C321 B.n281 VSUBS 0.008274f
C322 B.n282 VSUBS 0.008274f
C323 B.n283 VSUBS 0.005719f
C324 B.n284 VSUBS 0.008274f
C325 B.n285 VSUBS 0.008274f
C326 B.n286 VSUBS 0.008274f
C327 B.n287 VSUBS 0.008274f
C328 B.n288 VSUBS 0.008274f
C329 B.n289 VSUBS 0.008274f
C330 B.n290 VSUBS 0.008274f
C331 B.n291 VSUBS 0.008274f
C332 B.n292 VSUBS 0.008274f
C333 B.n293 VSUBS 0.008274f
C334 B.n294 VSUBS 0.008274f
C335 B.n295 VSUBS 0.008274f
C336 B.n296 VSUBS 0.008274f
C337 B.n297 VSUBS 0.008274f
C338 B.n298 VSUBS 0.008274f
C339 B.n299 VSUBS 0.008274f
C340 B.n300 VSUBS 0.008274f
C341 B.n301 VSUBS 0.008274f
C342 B.n302 VSUBS 0.008274f
C343 B.n303 VSUBS 0.008274f
C344 B.n304 VSUBS 0.008274f
C345 B.n305 VSUBS 0.008274f
C346 B.n306 VSUBS 0.008274f
C347 B.n307 VSUBS 0.008274f
C348 B.n308 VSUBS 0.008274f
C349 B.n309 VSUBS 0.008274f
C350 B.n310 VSUBS 0.008274f
C351 B.n311 VSUBS 0.008274f
C352 B.n312 VSUBS 0.008274f
C353 B.n313 VSUBS 0.008274f
C354 B.n314 VSUBS 0.008274f
C355 B.n315 VSUBS 0.008274f
C356 B.n316 VSUBS 0.008274f
C357 B.n317 VSUBS 0.020535f
C358 B.n318 VSUBS 0.019132f
C359 B.n319 VSUBS 0.019132f
C360 B.n320 VSUBS 0.008274f
C361 B.n321 VSUBS 0.008274f
C362 B.n322 VSUBS 0.008274f
C363 B.n323 VSUBS 0.008274f
C364 B.n324 VSUBS 0.008274f
C365 B.n325 VSUBS 0.008274f
C366 B.n326 VSUBS 0.008274f
C367 B.n327 VSUBS 0.008274f
C368 B.n328 VSUBS 0.008274f
C369 B.n329 VSUBS 0.008274f
C370 B.n330 VSUBS 0.008274f
C371 B.n331 VSUBS 0.008274f
C372 B.n332 VSUBS 0.008274f
C373 B.n333 VSUBS 0.008274f
C374 B.n334 VSUBS 0.008274f
C375 B.n335 VSUBS 0.008274f
C376 B.n336 VSUBS 0.008274f
C377 B.n337 VSUBS 0.008274f
C378 B.n338 VSUBS 0.008274f
C379 B.n339 VSUBS 0.008274f
C380 B.n340 VSUBS 0.008274f
C381 B.n341 VSUBS 0.008274f
C382 B.n342 VSUBS 0.008274f
C383 B.n343 VSUBS 0.008274f
C384 B.n344 VSUBS 0.008274f
C385 B.n345 VSUBS 0.008274f
C386 B.n346 VSUBS 0.008274f
C387 B.n347 VSUBS 0.008274f
C388 B.n348 VSUBS 0.008274f
C389 B.n349 VSUBS 0.008274f
C390 B.n350 VSUBS 0.008274f
C391 B.n351 VSUBS 0.008274f
C392 B.n352 VSUBS 0.008274f
C393 B.n353 VSUBS 0.008274f
C394 B.n354 VSUBS 0.008274f
C395 B.n355 VSUBS 0.008274f
C396 B.n356 VSUBS 0.008274f
C397 B.n357 VSUBS 0.008274f
C398 B.n358 VSUBS 0.008274f
C399 B.n359 VSUBS 0.008274f
C400 B.n360 VSUBS 0.008274f
C401 B.n361 VSUBS 0.008274f
C402 B.n362 VSUBS 0.008274f
C403 B.n363 VSUBS 0.008274f
C404 B.n364 VSUBS 0.008274f
C405 B.n365 VSUBS 0.008274f
C406 B.n366 VSUBS 0.008274f
C407 B.n367 VSUBS 0.008274f
C408 B.n368 VSUBS 0.008274f
C409 B.n369 VSUBS 0.008274f
C410 B.n370 VSUBS 0.008274f
C411 B.n371 VSUBS 0.008274f
C412 B.n372 VSUBS 0.008274f
C413 B.n373 VSUBS 0.008274f
C414 B.n374 VSUBS 0.008274f
C415 B.n375 VSUBS 0.008274f
C416 B.n376 VSUBS 0.008274f
C417 B.n377 VSUBS 0.008274f
C418 B.n378 VSUBS 0.008274f
C419 B.n379 VSUBS 0.008274f
C420 B.n380 VSUBS 0.008274f
C421 B.n381 VSUBS 0.008274f
C422 B.n382 VSUBS 0.008274f
C423 B.n383 VSUBS 0.008274f
C424 B.n384 VSUBS 0.008274f
C425 B.n385 VSUBS 0.008274f
C426 B.n386 VSUBS 0.008274f
C427 B.n387 VSUBS 0.008274f
C428 B.n388 VSUBS 0.008274f
C429 B.n389 VSUBS 0.008274f
C430 B.n390 VSUBS 0.008274f
C431 B.n391 VSUBS 0.008274f
C432 B.n392 VSUBS 0.008274f
C433 B.n393 VSUBS 0.008274f
C434 B.n394 VSUBS 0.008274f
C435 B.n395 VSUBS 0.008274f
C436 B.n396 VSUBS 0.008274f
C437 B.n397 VSUBS 0.008274f
C438 B.n398 VSUBS 0.008274f
C439 B.n399 VSUBS 0.008274f
C440 B.n400 VSUBS 0.008274f
C441 B.n401 VSUBS 0.008274f
C442 B.n402 VSUBS 0.008274f
C443 B.n403 VSUBS 0.008274f
C444 B.n404 VSUBS 0.008274f
C445 B.n405 VSUBS 0.008274f
C446 B.n406 VSUBS 0.008274f
C447 B.n407 VSUBS 0.008274f
C448 B.n408 VSUBS 0.008274f
C449 B.n409 VSUBS 0.008274f
C450 B.n410 VSUBS 0.008274f
C451 B.n411 VSUBS 0.008274f
C452 B.n412 VSUBS 0.008274f
C453 B.n413 VSUBS 0.008274f
C454 B.n414 VSUBS 0.008274f
C455 B.n415 VSUBS 0.008274f
C456 B.n416 VSUBS 0.008274f
C457 B.n417 VSUBS 0.008274f
C458 B.n418 VSUBS 0.008274f
C459 B.n419 VSUBS 0.008274f
C460 B.n420 VSUBS 0.008274f
C461 B.n421 VSUBS 0.008274f
C462 B.n422 VSUBS 0.008274f
C463 B.n423 VSUBS 0.008274f
C464 B.n424 VSUBS 0.008274f
C465 B.n425 VSUBS 0.008274f
C466 B.n426 VSUBS 0.008274f
C467 B.n427 VSUBS 0.008274f
C468 B.n428 VSUBS 0.008274f
C469 B.n429 VSUBS 0.008274f
C470 B.n430 VSUBS 0.008274f
C471 B.n431 VSUBS 0.008274f
C472 B.n432 VSUBS 0.008274f
C473 B.n433 VSUBS 0.008274f
C474 B.n434 VSUBS 0.008274f
C475 B.n435 VSUBS 0.008274f
C476 B.n436 VSUBS 0.008274f
C477 B.n437 VSUBS 0.008274f
C478 B.n438 VSUBS 0.008274f
C479 B.n439 VSUBS 0.008274f
C480 B.n440 VSUBS 0.008274f
C481 B.n441 VSUBS 0.008274f
C482 B.n442 VSUBS 0.008274f
C483 B.n443 VSUBS 0.008274f
C484 B.n444 VSUBS 0.008274f
C485 B.n445 VSUBS 0.008274f
C486 B.n446 VSUBS 0.008274f
C487 B.n447 VSUBS 0.008274f
C488 B.n448 VSUBS 0.008274f
C489 B.n449 VSUBS 0.008274f
C490 B.n450 VSUBS 0.008274f
C491 B.n451 VSUBS 0.008274f
C492 B.n452 VSUBS 0.008274f
C493 B.n453 VSUBS 0.008274f
C494 B.n454 VSUBS 0.008274f
C495 B.n455 VSUBS 0.008274f
C496 B.n456 VSUBS 0.008274f
C497 B.n457 VSUBS 0.008274f
C498 B.n458 VSUBS 0.008274f
C499 B.n459 VSUBS 0.020075f
C500 B.n460 VSUBS 0.019132f
C501 B.n461 VSUBS 0.020535f
C502 B.n462 VSUBS 0.008274f
C503 B.n463 VSUBS 0.008274f
C504 B.n464 VSUBS 0.008274f
C505 B.n465 VSUBS 0.008274f
C506 B.n466 VSUBS 0.008274f
C507 B.n467 VSUBS 0.008274f
C508 B.n468 VSUBS 0.008274f
C509 B.n469 VSUBS 0.008274f
C510 B.n470 VSUBS 0.008274f
C511 B.n471 VSUBS 0.008274f
C512 B.n472 VSUBS 0.008274f
C513 B.n473 VSUBS 0.008274f
C514 B.n474 VSUBS 0.008274f
C515 B.n475 VSUBS 0.008274f
C516 B.n476 VSUBS 0.008274f
C517 B.n477 VSUBS 0.008274f
C518 B.n478 VSUBS 0.008274f
C519 B.n479 VSUBS 0.008274f
C520 B.n480 VSUBS 0.008274f
C521 B.n481 VSUBS 0.008274f
C522 B.n482 VSUBS 0.008274f
C523 B.n483 VSUBS 0.008274f
C524 B.n484 VSUBS 0.008274f
C525 B.n485 VSUBS 0.008274f
C526 B.n486 VSUBS 0.008274f
C527 B.n487 VSUBS 0.008274f
C528 B.n488 VSUBS 0.008274f
C529 B.n489 VSUBS 0.008274f
C530 B.n490 VSUBS 0.008274f
C531 B.n491 VSUBS 0.008274f
C532 B.n492 VSUBS 0.008274f
C533 B.n493 VSUBS 0.008274f
C534 B.n494 VSUBS 0.008274f
C535 B.n495 VSUBS 0.005719f
C536 B.n496 VSUBS 0.008274f
C537 B.n497 VSUBS 0.008274f
C538 B.n498 VSUBS 0.006692f
C539 B.n499 VSUBS 0.008274f
C540 B.n500 VSUBS 0.008274f
C541 B.n501 VSUBS 0.008274f
C542 B.n502 VSUBS 0.008274f
C543 B.n503 VSUBS 0.008274f
C544 B.n504 VSUBS 0.008274f
C545 B.n505 VSUBS 0.008274f
C546 B.n506 VSUBS 0.008274f
C547 B.n507 VSUBS 0.008274f
C548 B.n508 VSUBS 0.008274f
C549 B.n509 VSUBS 0.008274f
C550 B.n510 VSUBS 0.006692f
C551 B.n511 VSUBS 0.01917f
C552 B.n512 VSUBS 0.005719f
C553 B.n513 VSUBS 0.008274f
C554 B.n514 VSUBS 0.008274f
C555 B.n515 VSUBS 0.008274f
C556 B.n516 VSUBS 0.008274f
C557 B.n517 VSUBS 0.008274f
C558 B.n518 VSUBS 0.008274f
C559 B.n519 VSUBS 0.008274f
C560 B.n520 VSUBS 0.008274f
C561 B.n521 VSUBS 0.008274f
C562 B.n522 VSUBS 0.008274f
C563 B.n523 VSUBS 0.008274f
C564 B.n524 VSUBS 0.008274f
C565 B.n525 VSUBS 0.008274f
C566 B.n526 VSUBS 0.008274f
C567 B.n527 VSUBS 0.008274f
C568 B.n528 VSUBS 0.008274f
C569 B.n529 VSUBS 0.008274f
C570 B.n530 VSUBS 0.008274f
C571 B.n531 VSUBS 0.008274f
C572 B.n532 VSUBS 0.008274f
C573 B.n533 VSUBS 0.008274f
C574 B.n534 VSUBS 0.008274f
C575 B.n535 VSUBS 0.008274f
C576 B.n536 VSUBS 0.008274f
C577 B.n537 VSUBS 0.008274f
C578 B.n538 VSUBS 0.008274f
C579 B.n539 VSUBS 0.008274f
C580 B.n540 VSUBS 0.008274f
C581 B.n541 VSUBS 0.008274f
C582 B.n542 VSUBS 0.008274f
C583 B.n543 VSUBS 0.008274f
C584 B.n544 VSUBS 0.008274f
C585 B.n545 VSUBS 0.008274f
C586 B.n546 VSUBS 0.020535f
C587 B.n547 VSUBS 0.020535f
C588 B.n548 VSUBS 0.019132f
C589 B.n549 VSUBS 0.008274f
C590 B.n550 VSUBS 0.008274f
C591 B.n551 VSUBS 0.008274f
C592 B.n552 VSUBS 0.008274f
C593 B.n553 VSUBS 0.008274f
C594 B.n554 VSUBS 0.008274f
C595 B.n555 VSUBS 0.008274f
C596 B.n556 VSUBS 0.008274f
C597 B.n557 VSUBS 0.008274f
C598 B.n558 VSUBS 0.008274f
C599 B.n559 VSUBS 0.008274f
C600 B.n560 VSUBS 0.008274f
C601 B.n561 VSUBS 0.008274f
C602 B.n562 VSUBS 0.008274f
C603 B.n563 VSUBS 0.008274f
C604 B.n564 VSUBS 0.008274f
C605 B.n565 VSUBS 0.008274f
C606 B.n566 VSUBS 0.008274f
C607 B.n567 VSUBS 0.008274f
C608 B.n568 VSUBS 0.008274f
C609 B.n569 VSUBS 0.008274f
C610 B.n570 VSUBS 0.008274f
C611 B.n571 VSUBS 0.008274f
C612 B.n572 VSUBS 0.008274f
C613 B.n573 VSUBS 0.008274f
C614 B.n574 VSUBS 0.008274f
C615 B.n575 VSUBS 0.008274f
C616 B.n576 VSUBS 0.008274f
C617 B.n577 VSUBS 0.008274f
C618 B.n578 VSUBS 0.008274f
C619 B.n579 VSUBS 0.008274f
C620 B.n580 VSUBS 0.008274f
C621 B.n581 VSUBS 0.008274f
C622 B.n582 VSUBS 0.008274f
C623 B.n583 VSUBS 0.008274f
C624 B.n584 VSUBS 0.008274f
C625 B.n585 VSUBS 0.008274f
C626 B.n586 VSUBS 0.008274f
C627 B.n587 VSUBS 0.008274f
C628 B.n588 VSUBS 0.008274f
C629 B.n589 VSUBS 0.008274f
C630 B.n590 VSUBS 0.008274f
C631 B.n591 VSUBS 0.008274f
C632 B.n592 VSUBS 0.008274f
C633 B.n593 VSUBS 0.008274f
C634 B.n594 VSUBS 0.008274f
C635 B.n595 VSUBS 0.008274f
C636 B.n596 VSUBS 0.008274f
C637 B.n597 VSUBS 0.008274f
C638 B.n598 VSUBS 0.008274f
C639 B.n599 VSUBS 0.008274f
C640 B.n600 VSUBS 0.008274f
C641 B.n601 VSUBS 0.008274f
C642 B.n602 VSUBS 0.008274f
C643 B.n603 VSUBS 0.008274f
C644 B.n604 VSUBS 0.008274f
C645 B.n605 VSUBS 0.008274f
C646 B.n606 VSUBS 0.008274f
C647 B.n607 VSUBS 0.008274f
C648 B.n608 VSUBS 0.008274f
C649 B.n609 VSUBS 0.008274f
C650 B.n610 VSUBS 0.008274f
C651 B.n611 VSUBS 0.008274f
C652 B.n612 VSUBS 0.008274f
C653 B.n613 VSUBS 0.008274f
C654 B.n614 VSUBS 0.008274f
C655 B.n615 VSUBS 0.008274f
C656 B.n616 VSUBS 0.008274f
C657 B.n617 VSUBS 0.008274f
C658 B.n618 VSUBS 0.008274f
C659 B.n619 VSUBS 0.018735f
C660 VDD1.t2 VSUBS 0.115169f
C661 VDD1.t1 VSUBS 0.115169f
C662 VDD1.n0 VSUBS 0.764532f
C663 VDD1.t5 VSUBS 0.115169f
C664 VDD1.t6 VSUBS 0.115169f
C665 VDD1.n1 VSUBS 0.763573f
C666 VDD1.t3 VSUBS 0.115169f
C667 VDD1.t4 VSUBS 0.115169f
C668 VDD1.n2 VSUBS 0.763573f
C669 VDD1.n3 VSUBS 3.17328f
C670 VDD1.t0 VSUBS 0.115169f
C671 VDD1.t7 VSUBS 0.115169f
C672 VDD1.n4 VSUBS 0.755372f
C673 VDD1.n5 VSUBS 2.59145f
C674 VP.n0 VSUBS 0.052548f
C675 VP.t3 VSUBS 1.44364f
C676 VP.n1 VSUBS 0.036508f
C677 VP.n2 VSUBS 0.039859f
C678 VP.t4 VSUBS 1.44364f
C679 VP.n3 VSUBS 0.073915f
C680 VP.n4 VSUBS 0.039859f
C681 VP.n5 VSUBS 0.043264f
C682 VP.n6 VSUBS 0.039859f
C683 VP.n7 VSUBS 0.079741f
C684 VP.n8 VSUBS 0.052548f
C685 VP.t0 VSUBS 1.44364f
C686 VP.n9 VSUBS 0.036508f
C687 VP.n10 VSUBS 0.039859f
C688 VP.t7 VSUBS 1.44364f
C689 VP.n11 VSUBS 0.073915f
C690 VP.n12 VSUBS 0.039859f
C691 VP.n13 VSUBS 0.043264f
C692 VP.t5 VSUBS 1.70494f
C693 VP.t6 VSUBS 1.44364f
C694 VP.n14 VSUBS 0.642144f
C695 VP.n15 VSUBS 0.637769f
C696 VP.n16 VSUBS 0.344281f
C697 VP.n17 VSUBS 0.039859f
C698 VP.n18 VSUBS 0.073915f
C699 VP.n19 VSUBS 0.057942f
C700 VP.n20 VSUBS 0.057942f
C701 VP.n21 VSUBS 0.039859f
C702 VP.n22 VSUBS 0.039859f
C703 VP.n23 VSUBS 0.039859f
C704 VP.n24 VSUBS 0.043264f
C705 VP.n25 VSUBS 0.546623f
C706 VP.n26 VSUBS 0.068077f
C707 VP.n27 VSUBS 0.07355f
C708 VP.n28 VSUBS 0.039859f
C709 VP.n29 VSUBS 0.039859f
C710 VP.n30 VSUBS 0.039859f
C711 VP.n31 VSUBS 0.079741f
C712 VP.n32 VSUBS 0.054941f
C713 VP.n33 VSUBS 0.668704f
C714 VP.n34 VSUBS 1.8843f
C715 VP.n35 VSUBS 1.91625f
C716 VP.t2 VSUBS 1.44364f
C717 VP.n36 VSUBS 0.668704f
C718 VP.n37 VSUBS 0.054941f
C719 VP.n38 VSUBS 0.052548f
C720 VP.n39 VSUBS 0.039859f
C721 VP.n40 VSUBS 0.039859f
C722 VP.n41 VSUBS 0.036508f
C723 VP.n42 VSUBS 0.07355f
C724 VP.t1 VSUBS 1.44364f
C725 VP.n43 VSUBS 0.546623f
C726 VP.n44 VSUBS 0.068077f
C727 VP.n45 VSUBS 0.039859f
C728 VP.n46 VSUBS 0.039859f
C729 VP.n47 VSUBS 0.039859f
C730 VP.n48 VSUBS 0.073915f
C731 VP.n49 VSUBS 0.057942f
C732 VP.n50 VSUBS 0.057942f
C733 VP.n51 VSUBS 0.039859f
C734 VP.n52 VSUBS 0.039859f
C735 VP.n53 VSUBS 0.039859f
C736 VP.n54 VSUBS 0.043264f
C737 VP.n55 VSUBS 0.546623f
C738 VP.n56 VSUBS 0.068077f
C739 VP.n57 VSUBS 0.07355f
C740 VP.n58 VSUBS 0.039859f
C741 VP.n59 VSUBS 0.039859f
C742 VP.n60 VSUBS 0.039859f
C743 VP.n61 VSUBS 0.079741f
C744 VP.n62 VSUBS 0.054941f
C745 VP.n63 VSUBS 0.668704f
C746 VP.n64 VSUBS 0.059852f
C747 VTAIL.t9 VSUBS 0.134517f
C748 VTAIL.t10 VSUBS 0.134517f
C749 VTAIL.n0 VSUBS 0.776258f
C750 VTAIL.n1 VSUBS 0.757339f
C751 VTAIL.n2 VSUBS 0.030216f
C752 VTAIL.n3 VSUBS 0.02895f
C753 VTAIL.n4 VSUBS 0.015556f
C754 VTAIL.n5 VSUBS 0.03677f
C755 VTAIL.n6 VSUBS 0.016471f
C756 VTAIL.n7 VSUBS 0.02895f
C757 VTAIL.n8 VSUBS 0.015556f
C758 VTAIL.n9 VSUBS 0.03677f
C759 VTAIL.n10 VSUBS 0.016471f
C760 VTAIL.n11 VSUBS 0.126789f
C761 VTAIL.t11 VSUBS 0.078702f
C762 VTAIL.n12 VSUBS 0.027577f
C763 VTAIL.n13 VSUBS 0.023379f
C764 VTAIL.n14 VSUBS 0.015556f
C765 VTAIL.n15 VSUBS 0.648691f
C766 VTAIL.n16 VSUBS 0.02895f
C767 VTAIL.n17 VSUBS 0.015556f
C768 VTAIL.n18 VSUBS 0.016471f
C769 VTAIL.n19 VSUBS 0.03677f
C770 VTAIL.n20 VSUBS 0.03677f
C771 VTAIL.n21 VSUBS 0.016471f
C772 VTAIL.n22 VSUBS 0.015556f
C773 VTAIL.n23 VSUBS 0.02895f
C774 VTAIL.n24 VSUBS 0.02895f
C775 VTAIL.n25 VSUBS 0.015556f
C776 VTAIL.n26 VSUBS 0.016471f
C777 VTAIL.n27 VSUBS 0.03677f
C778 VTAIL.n28 VSUBS 0.083587f
C779 VTAIL.n29 VSUBS 0.016471f
C780 VTAIL.n30 VSUBS 0.015556f
C781 VTAIL.n31 VSUBS 0.06217f
C782 VTAIL.n32 VSUBS 0.041643f
C783 VTAIL.n33 VSUBS 0.279785f
C784 VTAIL.n34 VSUBS 0.030216f
C785 VTAIL.n35 VSUBS 0.02895f
C786 VTAIL.n36 VSUBS 0.015556f
C787 VTAIL.n37 VSUBS 0.03677f
C788 VTAIL.n38 VSUBS 0.016471f
C789 VTAIL.n39 VSUBS 0.02895f
C790 VTAIL.n40 VSUBS 0.015556f
C791 VTAIL.n41 VSUBS 0.03677f
C792 VTAIL.n42 VSUBS 0.016471f
C793 VTAIL.n43 VSUBS 0.126789f
C794 VTAIL.t7 VSUBS 0.078702f
C795 VTAIL.n44 VSUBS 0.027577f
C796 VTAIL.n45 VSUBS 0.023379f
C797 VTAIL.n46 VSUBS 0.015556f
C798 VTAIL.n47 VSUBS 0.648691f
C799 VTAIL.n48 VSUBS 0.02895f
C800 VTAIL.n49 VSUBS 0.015556f
C801 VTAIL.n50 VSUBS 0.016471f
C802 VTAIL.n51 VSUBS 0.03677f
C803 VTAIL.n52 VSUBS 0.03677f
C804 VTAIL.n53 VSUBS 0.016471f
C805 VTAIL.n54 VSUBS 0.015556f
C806 VTAIL.n55 VSUBS 0.02895f
C807 VTAIL.n56 VSUBS 0.02895f
C808 VTAIL.n57 VSUBS 0.015556f
C809 VTAIL.n58 VSUBS 0.016471f
C810 VTAIL.n59 VSUBS 0.03677f
C811 VTAIL.n60 VSUBS 0.083587f
C812 VTAIL.n61 VSUBS 0.016471f
C813 VTAIL.n62 VSUBS 0.015556f
C814 VTAIL.n63 VSUBS 0.06217f
C815 VTAIL.n64 VSUBS 0.041643f
C816 VTAIL.n65 VSUBS 0.279785f
C817 VTAIL.t4 VSUBS 0.134517f
C818 VTAIL.t1 VSUBS 0.134517f
C819 VTAIL.n66 VSUBS 0.776258f
C820 VTAIL.n67 VSUBS 0.965818f
C821 VTAIL.n68 VSUBS 0.030216f
C822 VTAIL.n69 VSUBS 0.02895f
C823 VTAIL.n70 VSUBS 0.015556f
C824 VTAIL.n71 VSUBS 0.03677f
C825 VTAIL.n72 VSUBS 0.016471f
C826 VTAIL.n73 VSUBS 0.02895f
C827 VTAIL.n74 VSUBS 0.015556f
C828 VTAIL.n75 VSUBS 0.03677f
C829 VTAIL.n76 VSUBS 0.016471f
C830 VTAIL.n77 VSUBS 0.126789f
C831 VTAIL.t2 VSUBS 0.078702f
C832 VTAIL.n78 VSUBS 0.027577f
C833 VTAIL.n79 VSUBS 0.023379f
C834 VTAIL.n80 VSUBS 0.015556f
C835 VTAIL.n81 VSUBS 0.648691f
C836 VTAIL.n82 VSUBS 0.02895f
C837 VTAIL.n83 VSUBS 0.015556f
C838 VTAIL.n84 VSUBS 0.016471f
C839 VTAIL.n85 VSUBS 0.03677f
C840 VTAIL.n86 VSUBS 0.03677f
C841 VTAIL.n87 VSUBS 0.016471f
C842 VTAIL.n88 VSUBS 0.015556f
C843 VTAIL.n89 VSUBS 0.02895f
C844 VTAIL.n90 VSUBS 0.02895f
C845 VTAIL.n91 VSUBS 0.015556f
C846 VTAIL.n92 VSUBS 0.016471f
C847 VTAIL.n93 VSUBS 0.03677f
C848 VTAIL.n94 VSUBS 0.083587f
C849 VTAIL.n95 VSUBS 0.016471f
C850 VTAIL.n96 VSUBS 0.015556f
C851 VTAIL.n97 VSUBS 0.06217f
C852 VTAIL.n98 VSUBS 0.041643f
C853 VTAIL.n99 VSUBS 1.31596f
C854 VTAIL.n100 VSUBS 0.030216f
C855 VTAIL.n101 VSUBS 0.02895f
C856 VTAIL.n102 VSUBS 0.015556f
C857 VTAIL.n103 VSUBS 0.03677f
C858 VTAIL.n104 VSUBS 0.016471f
C859 VTAIL.n105 VSUBS 0.02895f
C860 VTAIL.n106 VSUBS 0.015556f
C861 VTAIL.n107 VSUBS 0.03677f
C862 VTAIL.n108 VSUBS 0.016471f
C863 VTAIL.n109 VSUBS 0.126789f
C864 VTAIL.t15 VSUBS 0.078702f
C865 VTAIL.n110 VSUBS 0.027577f
C866 VTAIL.n111 VSUBS 0.023379f
C867 VTAIL.n112 VSUBS 0.015556f
C868 VTAIL.n113 VSUBS 0.648691f
C869 VTAIL.n114 VSUBS 0.02895f
C870 VTAIL.n115 VSUBS 0.015556f
C871 VTAIL.n116 VSUBS 0.016471f
C872 VTAIL.n117 VSUBS 0.03677f
C873 VTAIL.n118 VSUBS 0.03677f
C874 VTAIL.n119 VSUBS 0.016471f
C875 VTAIL.n120 VSUBS 0.015556f
C876 VTAIL.n121 VSUBS 0.02895f
C877 VTAIL.n122 VSUBS 0.02895f
C878 VTAIL.n123 VSUBS 0.015556f
C879 VTAIL.n124 VSUBS 0.016471f
C880 VTAIL.n125 VSUBS 0.03677f
C881 VTAIL.n126 VSUBS 0.083587f
C882 VTAIL.n127 VSUBS 0.016471f
C883 VTAIL.n128 VSUBS 0.015556f
C884 VTAIL.n129 VSUBS 0.06217f
C885 VTAIL.n130 VSUBS 0.041643f
C886 VTAIL.n131 VSUBS 1.31596f
C887 VTAIL.t8 VSUBS 0.134517f
C888 VTAIL.t12 VSUBS 0.134517f
C889 VTAIL.n132 VSUBS 0.776264f
C890 VTAIL.n133 VSUBS 0.965812f
C891 VTAIL.n134 VSUBS 0.030216f
C892 VTAIL.n135 VSUBS 0.02895f
C893 VTAIL.n136 VSUBS 0.015556f
C894 VTAIL.n137 VSUBS 0.03677f
C895 VTAIL.n138 VSUBS 0.016471f
C896 VTAIL.n139 VSUBS 0.02895f
C897 VTAIL.n140 VSUBS 0.015556f
C898 VTAIL.n141 VSUBS 0.03677f
C899 VTAIL.n142 VSUBS 0.016471f
C900 VTAIL.n143 VSUBS 0.126789f
C901 VTAIL.t13 VSUBS 0.078702f
C902 VTAIL.n144 VSUBS 0.027577f
C903 VTAIL.n145 VSUBS 0.023379f
C904 VTAIL.n146 VSUBS 0.015556f
C905 VTAIL.n147 VSUBS 0.648691f
C906 VTAIL.n148 VSUBS 0.02895f
C907 VTAIL.n149 VSUBS 0.015556f
C908 VTAIL.n150 VSUBS 0.016471f
C909 VTAIL.n151 VSUBS 0.03677f
C910 VTAIL.n152 VSUBS 0.03677f
C911 VTAIL.n153 VSUBS 0.016471f
C912 VTAIL.n154 VSUBS 0.015556f
C913 VTAIL.n155 VSUBS 0.02895f
C914 VTAIL.n156 VSUBS 0.02895f
C915 VTAIL.n157 VSUBS 0.015556f
C916 VTAIL.n158 VSUBS 0.016471f
C917 VTAIL.n159 VSUBS 0.03677f
C918 VTAIL.n160 VSUBS 0.083587f
C919 VTAIL.n161 VSUBS 0.016471f
C920 VTAIL.n162 VSUBS 0.015556f
C921 VTAIL.n163 VSUBS 0.06217f
C922 VTAIL.n164 VSUBS 0.041643f
C923 VTAIL.n165 VSUBS 0.279785f
C924 VTAIL.n166 VSUBS 0.030216f
C925 VTAIL.n167 VSUBS 0.02895f
C926 VTAIL.n168 VSUBS 0.015556f
C927 VTAIL.n169 VSUBS 0.03677f
C928 VTAIL.n170 VSUBS 0.016471f
C929 VTAIL.n171 VSUBS 0.02895f
C930 VTAIL.n172 VSUBS 0.015556f
C931 VTAIL.n173 VSUBS 0.03677f
C932 VTAIL.n174 VSUBS 0.016471f
C933 VTAIL.n175 VSUBS 0.126789f
C934 VTAIL.t3 VSUBS 0.078702f
C935 VTAIL.n176 VSUBS 0.027577f
C936 VTAIL.n177 VSUBS 0.023379f
C937 VTAIL.n178 VSUBS 0.015556f
C938 VTAIL.n179 VSUBS 0.648691f
C939 VTAIL.n180 VSUBS 0.02895f
C940 VTAIL.n181 VSUBS 0.015556f
C941 VTAIL.n182 VSUBS 0.016471f
C942 VTAIL.n183 VSUBS 0.03677f
C943 VTAIL.n184 VSUBS 0.03677f
C944 VTAIL.n185 VSUBS 0.016471f
C945 VTAIL.n186 VSUBS 0.015556f
C946 VTAIL.n187 VSUBS 0.02895f
C947 VTAIL.n188 VSUBS 0.02895f
C948 VTAIL.n189 VSUBS 0.015556f
C949 VTAIL.n190 VSUBS 0.016471f
C950 VTAIL.n191 VSUBS 0.03677f
C951 VTAIL.n192 VSUBS 0.083587f
C952 VTAIL.n193 VSUBS 0.016471f
C953 VTAIL.n194 VSUBS 0.015556f
C954 VTAIL.n195 VSUBS 0.06217f
C955 VTAIL.n196 VSUBS 0.041643f
C956 VTAIL.n197 VSUBS 0.279785f
C957 VTAIL.t6 VSUBS 0.134517f
C958 VTAIL.t5 VSUBS 0.134517f
C959 VTAIL.n198 VSUBS 0.776264f
C960 VTAIL.n199 VSUBS 0.965812f
C961 VTAIL.n200 VSUBS 0.030216f
C962 VTAIL.n201 VSUBS 0.02895f
C963 VTAIL.n202 VSUBS 0.015556f
C964 VTAIL.n203 VSUBS 0.03677f
C965 VTAIL.n204 VSUBS 0.016471f
C966 VTAIL.n205 VSUBS 0.02895f
C967 VTAIL.n206 VSUBS 0.015556f
C968 VTAIL.n207 VSUBS 0.03677f
C969 VTAIL.n208 VSUBS 0.016471f
C970 VTAIL.n209 VSUBS 0.126789f
C971 VTAIL.t0 VSUBS 0.078702f
C972 VTAIL.n210 VSUBS 0.027577f
C973 VTAIL.n211 VSUBS 0.023379f
C974 VTAIL.n212 VSUBS 0.015556f
C975 VTAIL.n213 VSUBS 0.648691f
C976 VTAIL.n214 VSUBS 0.02895f
C977 VTAIL.n215 VSUBS 0.015556f
C978 VTAIL.n216 VSUBS 0.016471f
C979 VTAIL.n217 VSUBS 0.03677f
C980 VTAIL.n218 VSUBS 0.03677f
C981 VTAIL.n219 VSUBS 0.016471f
C982 VTAIL.n220 VSUBS 0.015556f
C983 VTAIL.n221 VSUBS 0.02895f
C984 VTAIL.n222 VSUBS 0.02895f
C985 VTAIL.n223 VSUBS 0.015556f
C986 VTAIL.n224 VSUBS 0.016471f
C987 VTAIL.n225 VSUBS 0.03677f
C988 VTAIL.n226 VSUBS 0.083587f
C989 VTAIL.n227 VSUBS 0.016471f
C990 VTAIL.n228 VSUBS 0.015556f
C991 VTAIL.n229 VSUBS 0.06217f
C992 VTAIL.n230 VSUBS 0.041643f
C993 VTAIL.n231 VSUBS 1.31596f
C994 VTAIL.n232 VSUBS 0.030216f
C995 VTAIL.n233 VSUBS 0.02895f
C996 VTAIL.n234 VSUBS 0.015556f
C997 VTAIL.n235 VSUBS 0.03677f
C998 VTAIL.n236 VSUBS 0.016471f
C999 VTAIL.n237 VSUBS 0.02895f
C1000 VTAIL.n238 VSUBS 0.015556f
C1001 VTAIL.n239 VSUBS 0.03677f
C1002 VTAIL.n240 VSUBS 0.016471f
C1003 VTAIL.n241 VSUBS 0.126789f
C1004 VTAIL.t14 VSUBS 0.078702f
C1005 VTAIL.n242 VSUBS 0.027577f
C1006 VTAIL.n243 VSUBS 0.023379f
C1007 VTAIL.n244 VSUBS 0.015556f
C1008 VTAIL.n245 VSUBS 0.648691f
C1009 VTAIL.n246 VSUBS 0.02895f
C1010 VTAIL.n247 VSUBS 0.015556f
C1011 VTAIL.n248 VSUBS 0.016471f
C1012 VTAIL.n249 VSUBS 0.03677f
C1013 VTAIL.n250 VSUBS 0.03677f
C1014 VTAIL.n251 VSUBS 0.016471f
C1015 VTAIL.n252 VSUBS 0.015556f
C1016 VTAIL.n253 VSUBS 0.02895f
C1017 VTAIL.n254 VSUBS 0.02895f
C1018 VTAIL.n255 VSUBS 0.015556f
C1019 VTAIL.n256 VSUBS 0.016471f
C1020 VTAIL.n257 VSUBS 0.03677f
C1021 VTAIL.n258 VSUBS 0.083587f
C1022 VTAIL.n259 VSUBS 0.016471f
C1023 VTAIL.n260 VSUBS 0.015556f
C1024 VTAIL.n261 VSUBS 0.06217f
C1025 VTAIL.n262 VSUBS 0.041643f
C1026 VTAIL.n263 VSUBS 1.31053f
C1027 VDD2.t0 VSUBS 0.112884f
C1028 VDD2.t1 VSUBS 0.112884f
C1029 VDD2.n0 VSUBS 0.748426f
C1030 VDD2.t7 VSUBS 0.112884f
C1031 VDD2.t3 VSUBS 0.112884f
C1032 VDD2.n1 VSUBS 0.748426f
C1033 VDD2.n2 VSUBS 3.0594f
C1034 VDD2.t4 VSUBS 0.112884f
C1035 VDD2.t5 VSUBS 0.112884f
C1036 VDD2.n3 VSUBS 0.740392f
C1037 VDD2.n4 VSUBS 2.51036f
C1038 VDD2.t6 VSUBS 0.112884f
C1039 VDD2.t2 VSUBS 0.112884f
C1040 VDD2.n5 VSUBS 0.748397f
C1041 VN.n0 VSUBS 0.050654f
C1042 VN.t1 VSUBS 1.39162f
C1043 VN.n1 VSUBS 0.035193f
C1044 VN.n2 VSUBS 0.038423f
C1045 VN.t5 VSUBS 1.39162f
C1046 VN.n3 VSUBS 0.071252f
C1047 VN.n4 VSUBS 0.038423f
C1048 VN.n5 VSUBS 0.041705f
C1049 VN.t4 VSUBS 1.6435f
C1050 VN.t6 VSUBS 1.39162f
C1051 VN.n6 VSUBS 0.619005f
C1052 VN.n7 VSUBS 0.614787f
C1053 VN.n8 VSUBS 0.331875f
C1054 VN.n9 VSUBS 0.038423f
C1055 VN.n10 VSUBS 0.071252f
C1056 VN.n11 VSUBS 0.055854f
C1057 VN.n12 VSUBS 0.055854f
C1058 VN.n13 VSUBS 0.038423f
C1059 VN.n14 VSUBS 0.038423f
C1060 VN.n15 VSUBS 0.038423f
C1061 VN.n16 VSUBS 0.041705f
C1062 VN.n17 VSUBS 0.526926f
C1063 VN.n18 VSUBS 0.065624f
C1064 VN.n19 VSUBS 0.070899f
C1065 VN.n20 VSUBS 0.038423f
C1066 VN.n21 VSUBS 0.038423f
C1067 VN.n22 VSUBS 0.038423f
C1068 VN.n23 VSUBS 0.076868f
C1069 VN.n24 VSUBS 0.052961f
C1070 VN.n25 VSUBS 0.644608f
C1071 VN.n26 VSUBS 0.057695f
C1072 VN.n27 VSUBS 0.050654f
C1073 VN.t0 VSUBS 1.39162f
C1074 VN.n28 VSUBS 0.035193f
C1075 VN.n29 VSUBS 0.038423f
C1076 VN.t7 VSUBS 1.39162f
C1077 VN.n30 VSUBS 0.071252f
C1078 VN.n31 VSUBS 0.038423f
C1079 VN.n32 VSUBS 0.041705f
C1080 VN.t2 VSUBS 1.6435f
C1081 VN.t3 VSUBS 1.39162f
C1082 VN.n33 VSUBS 0.619005f
C1083 VN.n34 VSUBS 0.614787f
C1084 VN.n35 VSUBS 0.331875f
C1085 VN.n36 VSUBS 0.038423f
C1086 VN.n37 VSUBS 0.071252f
C1087 VN.n38 VSUBS 0.055854f
C1088 VN.n39 VSUBS 0.055854f
C1089 VN.n40 VSUBS 0.038423f
C1090 VN.n41 VSUBS 0.038423f
C1091 VN.n42 VSUBS 0.038423f
C1092 VN.n43 VSUBS 0.041705f
C1093 VN.n44 VSUBS 0.526926f
C1094 VN.n45 VSUBS 0.065624f
C1095 VN.n46 VSUBS 0.070899f
C1096 VN.n47 VSUBS 0.038423f
C1097 VN.n48 VSUBS 0.038423f
C1098 VN.n49 VSUBS 0.038423f
C1099 VN.n50 VSUBS 0.076868f
C1100 VN.n51 VSUBS 0.052961f
C1101 VN.n52 VSUBS 0.644608f
C1102 VN.n53 VSUBS 1.83742f
.ends

