* NGSPICE file created from diff_pair_sample_1582.ext - technology: sky130A

.subckt diff_pair_sample_1582 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=2.7852 pd=17.21 as=6.5832 ps=34.54 w=16.88 l=0.44
X1 B.t11 B.t9 B.t10 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=0 ps=0 w=16.88 l=0.44
X2 VTAIL.t0 VN.t0 VDD2.t3 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=2.7852 ps=17.21 w=16.88 l=0.44
X3 B.t8 B.t6 B.t7 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=0 ps=0 w=16.88 l=0.44
X4 VTAIL.t4 VP.t1 VDD1.t2 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=2.7852 ps=17.21 w=16.88 l=0.44
X5 VDD2.t2 VN.t1 VTAIL.t1 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=2.7852 pd=17.21 as=6.5832 ps=34.54 w=16.88 l=0.44
X6 VDD2.t1 VN.t2 VTAIL.t2 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=2.7852 pd=17.21 as=6.5832 ps=34.54 w=16.88 l=0.44
X7 B.t5 B.t3 B.t4 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=0 ps=0 w=16.88 l=0.44
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=2.7852 ps=17.21 w=16.88 l=0.44
X9 VDD1.t1 VP.t2 VTAIL.t5 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=2.7852 pd=17.21 as=6.5832 ps=34.54 w=16.88 l=0.44
X10 VTAIL.t6 VP.t3 VDD1.t0 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=2.7852 ps=17.21 w=16.88 l=0.44
X11 B.t2 B.t0 B.t1 w_n1432_n4344# sky130_fd_pr__pfet_01v8 ad=6.5832 pd=34.54 as=0 ps=0 w=16.88 l=0.44
R0 VP.n0 VP.t3 1034.82
R1 VP.n0 VP.t0 1034.8
R2 VP.n2 VP.t1 1013.84
R3 VP.n3 VP.t2 1013.84
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 113.525
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n746 VTAIL.n658 756.745
R11 VTAIL.n88 VTAIL.n0 756.745
R12 VTAIL.n182 VTAIL.n94 756.745
R13 VTAIL.n276 VTAIL.n188 756.745
R14 VTAIL.n652 VTAIL.n564 756.745
R15 VTAIL.n558 VTAIL.n470 756.745
R16 VTAIL.n464 VTAIL.n376 756.745
R17 VTAIL.n370 VTAIL.n282 756.745
R18 VTAIL.n689 VTAIL.n688 585
R19 VTAIL.n686 VTAIL.n685 585
R20 VTAIL.n695 VTAIL.n694 585
R21 VTAIL.n697 VTAIL.n696 585
R22 VTAIL.n682 VTAIL.n681 585
R23 VTAIL.n703 VTAIL.n702 585
R24 VTAIL.n705 VTAIL.n704 585
R25 VTAIL.n678 VTAIL.n677 585
R26 VTAIL.n711 VTAIL.n710 585
R27 VTAIL.n713 VTAIL.n712 585
R28 VTAIL.n674 VTAIL.n673 585
R29 VTAIL.n719 VTAIL.n718 585
R30 VTAIL.n721 VTAIL.n720 585
R31 VTAIL.n670 VTAIL.n669 585
R32 VTAIL.n727 VTAIL.n726 585
R33 VTAIL.n730 VTAIL.n729 585
R34 VTAIL.n728 VTAIL.n666 585
R35 VTAIL.n735 VTAIL.n665 585
R36 VTAIL.n737 VTAIL.n736 585
R37 VTAIL.n739 VTAIL.n738 585
R38 VTAIL.n662 VTAIL.n661 585
R39 VTAIL.n745 VTAIL.n744 585
R40 VTAIL.n747 VTAIL.n746 585
R41 VTAIL.n31 VTAIL.n30 585
R42 VTAIL.n28 VTAIL.n27 585
R43 VTAIL.n37 VTAIL.n36 585
R44 VTAIL.n39 VTAIL.n38 585
R45 VTAIL.n24 VTAIL.n23 585
R46 VTAIL.n45 VTAIL.n44 585
R47 VTAIL.n47 VTAIL.n46 585
R48 VTAIL.n20 VTAIL.n19 585
R49 VTAIL.n53 VTAIL.n52 585
R50 VTAIL.n55 VTAIL.n54 585
R51 VTAIL.n16 VTAIL.n15 585
R52 VTAIL.n61 VTAIL.n60 585
R53 VTAIL.n63 VTAIL.n62 585
R54 VTAIL.n12 VTAIL.n11 585
R55 VTAIL.n69 VTAIL.n68 585
R56 VTAIL.n72 VTAIL.n71 585
R57 VTAIL.n70 VTAIL.n8 585
R58 VTAIL.n77 VTAIL.n7 585
R59 VTAIL.n79 VTAIL.n78 585
R60 VTAIL.n81 VTAIL.n80 585
R61 VTAIL.n4 VTAIL.n3 585
R62 VTAIL.n87 VTAIL.n86 585
R63 VTAIL.n89 VTAIL.n88 585
R64 VTAIL.n125 VTAIL.n124 585
R65 VTAIL.n122 VTAIL.n121 585
R66 VTAIL.n131 VTAIL.n130 585
R67 VTAIL.n133 VTAIL.n132 585
R68 VTAIL.n118 VTAIL.n117 585
R69 VTAIL.n139 VTAIL.n138 585
R70 VTAIL.n141 VTAIL.n140 585
R71 VTAIL.n114 VTAIL.n113 585
R72 VTAIL.n147 VTAIL.n146 585
R73 VTAIL.n149 VTAIL.n148 585
R74 VTAIL.n110 VTAIL.n109 585
R75 VTAIL.n155 VTAIL.n154 585
R76 VTAIL.n157 VTAIL.n156 585
R77 VTAIL.n106 VTAIL.n105 585
R78 VTAIL.n163 VTAIL.n162 585
R79 VTAIL.n166 VTAIL.n165 585
R80 VTAIL.n164 VTAIL.n102 585
R81 VTAIL.n171 VTAIL.n101 585
R82 VTAIL.n173 VTAIL.n172 585
R83 VTAIL.n175 VTAIL.n174 585
R84 VTAIL.n98 VTAIL.n97 585
R85 VTAIL.n181 VTAIL.n180 585
R86 VTAIL.n183 VTAIL.n182 585
R87 VTAIL.n219 VTAIL.n218 585
R88 VTAIL.n216 VTAIL.n215 585
R89 VTAIL.n225 VTAIL.n224 585
R90 VTAIL.n227 VTAIL.n226 585
R91 VTAIL.n212 VTAIL.n211 585
R92 VTAIL.n233 VTAIL.n232 585
R93 VTAIL.n235 VTAIL.n234 585
R94 VTAIL.n208 VTAIL.n207 585
R95 VTAIL.n241 VTAIL.n240 585
R96 VTAIL.n243 VTAIL.n242 585
R97 VTAIL.n204 VTAIL.n203 585
R98 VTAIL.n249 VTAIL.n248 585
R99 VTAIL.n251 VTAIL.n250 585
R100 VTAIL.n200 VTAIL.n199 585
R101 VTAIL.n257 VTAIL.n256 585
R102 VTAIL.n260 VTAIL.n259 585
R103 VTAIL.n258 VTAIL.n196 585
R104 VTAIL.n265 VTAIL.n195 585
R105 VTAIL.n267 VTAIL.n266 585
R106 VTAIL.n269 VTAIL.n268 585
R107 VTAIL.n192 VTAIL.n191 585
R108 VTAIL.n275 VTAIL.n274 585
R109 VTAIL.n277 VTAIL.n276 585
R110 VTAIL.n653 VTAIL.n652 585
R111 VTAIL.n651 VTAIL.n650 585
R112 VTAIL.n568 VTAIL.n567 585
R113 VTAIL.n645 VTAIL.n644 585
R114 VTAIL.n643 VTAIL.n642 585
R115 VTAIL.n641 VTAIL.n571 585
R116 VTAIL.n575 VTAIL.n572 585
R117 VTAIL.n636 VTAIL.n635 585
R118 VTAIL.n634 VTAIL.n633 585
R119 VTAIL.n577 VTAIL.n576 585
R120 VTAIL.n628 VTAIL.n627 585
R121 VTAIL.n626 VTAIL.n625 585
R122 VTAIL.n581 VTAIL.n580 585
R123 VTAIL.n620 VTAIL.n619 585
R124 VTAIL.n618 VTAIL.n617 585
R125 VTAIL.n585 VTAIL.n584 585
R126 VTAIL.n612 VTAIL.n611 585
R127 VTAIL.n610 VTAIL.n609 585
R128 VTAIL.n589 VTAIL.n588 585
R129 VTAIL.n604 VTAIL.n603 585
R130 VTAIL.n602 VTAIL.n601 585
R131 VTAIL.n593 VTAIL.n592 585
R132 VTAIL.n596 VTAIL.n595 585
R133 VTAIL.n559 VTAIL.n558 585
R134 VTAIL.n557 VTAIL.n556 585
R135 VTAIL.n474 VTAIL.n473 585
R136 VTAIL.n551 VTAIL.n550 585
R137 VTAIL.n549 VTAIL.n548 585
R138 VTAIL.n547 VTAIL.n477 585
R139 VTAIL.n481 VTAIL.n478 585
R140 VTAIL.n542 VTAIL.n541 585
R141 VTAIL.n540 VTAIL.n539 585
R142 VTAIL.n483 VTAIL.n482 585
R143 VTAIL.n534 VTAIL.n533 585
R144 VTAIL.n532 VTAIL.n531 585
R145 VTAIL.n487 VTAIL.n486 585
R146 VTAIL.n526 VTAIL.n525 585
R147 VTAIL.n524 VTAIL.n523 585
R148 VTAIL.n491 VTAIL.n490 585
R149 VTAIL.n518 VTAIL.n517 585
R150 VTAIL.n516 VTAIL.n515 585
R151 VTAIL.n495 VTAIL.n494 585
R152 VTAIL.n510 VTAIL.n509 585
R153 VTAIL.n508 VTAIL.n507 585
R154 VTAIL.n499 VTAIL.n498 585
R155 VTAIL.n502 VTAIL.n501 585
R156 VTAIL.n465 VTAIL.n464 585
R157 VTAIL.n463 VTAIL.n462 585
R158 VTAIL.n380 VTAIL.n379 585
R159 VTAIL.n457 VTAIL.n456 585
R160 VTAIL.n455 VTAIL.n454 585
R161 VTAIL.n453 VTAIL.n383 585
R162 VTAIL.n387 VTAIL.n384 585
R163 VTAIL.n448 VTAIL.n447 585
R164 VTAIL.n446 VTAIL.n445 585
R165 VTAIL.n389 VTAIL.n388 585
R166 VTAIL.n440 VTAIL.n439 585
R167 VTAIL.n438 VTAIL.n437 585
R168 VTAIL.n393 VTAIL.n392 585
R169 VTAIL.n432 VTAIL.n431 585
R170 VTAIL.n430 VTAIL.n429 585
R171 VTAIL.n397 VTAIL.n396 585
R172 VTAIL.n424 VTAIL.n423 585
R173 VTAIL.n422 VTAIL.n421 585
R174 VTAIL.n401 VTAIL.n400 585
R175 VTAIL.n416 VTAIL.n415 585
R176 VTAIL.n414 VTAIL.n413 585
R177 VTAIL.n405 VTAIL.n404 585
R178 VTAIL.n408 VTAIL.n407 585
R179 VTAIL.n371 VTAIL.n370 585
R180 VTAIL.n369 VTAIL.n368 585
R181 VTAIL.n286 VTAIL.n285 585
R182 VTAIL.n363 VTAIL.n362 585
R183 VTAIL.n361 VTAIL.n360 585
R184 VTAIL.n359 VTAIL.n289 585
R185 VTAIL.n293 VTAIL.n290 585
R186 VTAIL.n354 VTAIL.n353 585
R187 VTAIL.n352 VTAIL.n351 585
R188 VTAIL.n295 VTAIL.n294 585
R189 VTAIL.n346 VTAIL.n345 585
R190 VTAIL.n344 VTAIL.n343 585
R191 VTAIL.n299 VTAIL.n298 585
R192 VTAIL.n338 VTAIL.n337 585
R193 VTAIL.n336 VTAIL.n335 585
R194 VTAIL.n303 VTAIL.n302 585
R195 VTAIL.n330 VTAIL.n329 585
R196 VTAIL.n328 VTAIL.n327 585
R197 VTAIL.n307 VTAIL.n306 585
R198 VTAIL.n322 VTAIL.n321 585
R199 VTAIL.n320 VTAIL.n319 585
R200 VTAIL.n311 VTAIL.n310 585
R201 VTAIL.n314 VTAIL.n313 585
R202 VTAIL.t7 VTAIL.n594 327.466
R203 VTAIL.t6 VTAIL.n500 327.466
R204 VTAIL.t1 VTAIL.n406 327.466
R205 VTAIL.t3 VTAIL.n312 327.466
R206 VTAIL.t2 VTAIL.n687 327.466
R207 VTAIL.t0 VTAIL.n29 327.466
R208 VTAIL.t5 VTAIL.n123 327.466
R209 VTAIL.t4 VTAIL.n217 327.466
R210 VTAIL.n688 VTAIL.n685 171.744
R211 VTAIL.n695 VTAIL.n685 171.744
R212 VTAIL.n696 VTAIL.n695 171.744
R213 VTAIL.n696 VTAIL.n681 171.744
R214 VTAIL.n703 VTAIL.n681 171.744
R215 VTAIL.n704 VTAIL.n703 171.744
R216 VTAIL.n704 VTAIL.n677 171.744
R217 VTAIL.n711 VTAIL.n677 171.744
R218 VTAIL.n712 VTAIL.n711 171.744
R219 VTAIL.n712 VTAIL.n673 171.744
R220 VTAIL.n719 VTAIL.n673 171.744
R221 VTAIL.n720 VTAIL.n719 171.744
R222 VTAIL.n720 VTAIL.n669 171.744
R223 VTAIL.n727 VTAIL.n669 171.744
R224 VTAIL.n729 VTAIL.n727 171.744
R225 VTAIL.n729 VTAIL.n728 171.744
R226 VTAIL.n728 VTAIL.n665 171.744
R227 VTAIL.n737 VTAIL.n665 171.744
R228 VTAIL.n738 VTAIL.n737 171.744
R229 VTAIL.n738 VTAIL.n661 171.744
R230 VTAIL.n745 VTAIL.n661 171.744
R231 VTAIL.n746 VTAIL.n745 171.744
R232 VTAIL.n30 VTAIL.n27 171.744
R233 VTAIL.n37 VTAIL.n27 171.744
R234 VTAIL.n38 VTAIL.n37 171.744
R235 VTAIL.n38 VTAIL.n23 171.744
R236 VTAIL.n45 VTAIL.n23 171.744
R237 VTAIL.n46 VTAIL.n45 171.744
R238 VTAIL.n46 VTAIL.n19 171.744
R239 VTAIL.n53 VTAIL.n19 171.744
R240 VTAIL.n54 VTAIL.n53 171.744
R241 VTAIL.n54 VTAIL.n15 171.744
R242 VTAIL.n61 VTAIL.n15 171.744
R243 VTAIL.n62 VTAIL.n61 171.744
R244 VTAIL.n62 VTAIL.n11 171.744
R245 VTAIL.n69 VTAIL.n11 171.744
R246 VTAIL.n71 VTAIL.n69 171.744
R247 VTAIL.n71 VTAIL.n70 171.744
R248 VTAIL.n70 VTAIL.n7 171.744
R249 VTAIL.n79 VTAIL.n7 171.744
R250 VTAIL.n80 VTAIL.n79 171.744
R251 VTAIL.n80 VTAIL.n3 171.744
R252 VTAIL.n87 VTAIL.n3 171.744
R253 VTAIL.n88 VTAIL.n87 171.744
R254 VTAIL.n124 VTAIL.n121 171.744
R255 VTAIL.n131 VTAIL.n121 171.744
R256 VTAIL.n132 VTAIL.n131 171.744
R257 VTAIL.n132 VTAIL.n117 171.744
R258 VTAIL.n139 VTAIL.n117 171.744
R259 VTAIL.n140 VTAIL.n139 171.744
R260 VTAIL.n140 VTAIL.n113 171.744
R261 VTAIL.n147 VTAIL.n113 171.744
R262 VTAIL.n148 VTAIL.n147 171.744
R263 VTAIL.n148 VTAIL.n109 171.744
R264 VTAIL.n155 VTAIL.n109 171.744
R265 VTAIL.n156 VTAIL.n155 171.744
R266 VTAIL.n156 VTAIL.n105 171.744
R267 VTAIL.n163 VTAIL.n105 171.744
R268 VTAIL.n165 VTAIL.n163 171.744
R269 VTAIL.n165 VTAIL.n164 171.744
R270 VTAIL.n164 VTAIL.n101 171.744
R271 VTAIL.n173 VTAIL.n101 171.744
R272 VTAIL.n174 VTAIL.n173 171.744
R273 VTAIL.n174 VTAIL.n97 171.744
R274 VTAIL.n181 VTAIL.n97 171.744
R275 VTAIL.n182 VTAIL.n181 171.744
R276 VTAIL.n218 VTAIL.n215 171.744
R277 VTAIL.n225 VTAIL.n215 171.744
R278 VTAIL.n226 VTAIL.n225 171.744
R279 VTAIL.n226 VTAIL.n211 171.744
R280 VTAIL.n233 VTAIL.n211 171.744
R281 VTAIL.n234 VTAIL.n233 171.744
R282 VTAIL.n234 VTAIL.n207 171.744
R283 VTAIL.n241 VTAIL.n207 171.744
R284 VTAIL.n242 VTAIL.n241 171.744
R285 VTAIL.n242 VTAIL.n203 171.744
R286 VTAIL.n249 VTAIL.n203 171.744
R287 VTAIL.n250 VTAIL.n249 171.744
R288 VTAIL.n250 VTAIL.n199 171.744
R289 VTAIL.n257 VTAIL.n199 171.744
R290 VTAIL.n259 VTAIL.n257 171.744
R291 VTAIL.n259 VTAIL.n258 171.744
R292 VTAIL.n258 VTAIL.n195 171.744
R293 VTAIL.n267 VTAIL.n195 171.744
R294 VTAIL.n268 VTAIL.n267 171.744
R295 VTAIL.n268 VTAIL.n191 171.744
R296 VTAIL.n275 VTAIL.n191 171.744
R297 VTAIL.n276 VTAIL.n275 171.744
R298 VTAIL.n652 VTAIL.n651 171.744
R299 VTAIL.n651 VTAIL.n567 171.744
R300 VTAIL.n644 VTAIL.n567 171.744
R301 VTAIL.n644 VTAIL.n643 171.744
R302 VTAIL.n643 VTAIL.n571 171.744
R303 VTAIL.n575 VTAIL.n571 171.744
R304 VTAIL.n635 VTAIL.n575 171.744
R305 VTAIL.n635 VTAIL.n634 171.744
R306 VTAIL.n634 VTAIL.n576 171.744
R307 VTAIL.n627 VTAIL.n576 171.744
R308 VTAIL.n627 VTAIL.n626 171.744
R309 VTAIL.n626 VTAIL.n580 171.744
R310 VTAIL.n619 VTAIL.n580 171.744
R311 VTAIL.n619 VTAIL.n618 171.744
R312 VTAIL.n618 VTAIL.n584 171.744
R313 VTAIL.n611 VTAIL.n584 171.744
R314 VTAIL.n611 VTAIL.n610 171.744
R315 VTAIL.n610 VTAIL.n588 171.744
R316 VTAIL.n603 VTAIL.n588 171.744
R317 VTAIL.n603 VTAIL.n602 171.744
R318 VTAIL.n602 VTAIL.n592 171.744
R319 VTAIL.n595 VTAIL.n592 171.744
R320 VTAIL.n558 VTAIL.n557 171.744
R321 VTAIL.n557 VTAIL.n473 171.744
R322 VTAIL.n550 VTAIL.n473 171.744
R323 VTAIL.n550 VTAIL.n549 171.744
R324 VTAIL.n549 VTAIL.n477 171.744
R325 VTAIL.n481 VTAIL.n477 171.744
R326 VTAIL.n541 VTAIL.n481 171.744
R327 VTAIL.n541 VTAIL.n540 171.744
R328 VTAIL.n540 VTAIL.n482 171.744
R329 VTAIL.n533 VTAIL.n482 171.744
R330 VTAIL.n533 VTAIL.n532 171.744
R331 VTAIL.n532 VTAIL.n486 171.744
R332 VTAIL.n525 VTAIL.n486 171.744
R333 VTAIL.n525 VTAIL.n524 171.744
R334 VTAIL.n524 VTAIL.n490 171.744
R335 VTAIL.n517 VTAIL.n490 171.744
R336 VTAIL.n517 VTAIL.n516 171.744
R337 VTAIL.n516 VTAIL.n494 171.744
R338 VTAIL.n509 VTAIL.n494 171.744
R339 VTAIL.n509 VTAIL.n508 171.744
R340 VTAIL.n508 VTAIL.n498 171.744
R341 VTAIL.n501 VTAIL.n498 171.744
R342 VTAIL.n464 VTAIL.n463 171.744
R343 VTAIL.n463 VTAIL.n379 171.744
R344 VTAIL.n456 VTAIL.n379 171.744
R345 VTAIL.n456 VTAIL.n455 171.744
R346 VTAIL.n455 VTAIL.n383 171.744
R347 VTAIL.n387 VTAIL.n383 171.744
R348 VTAIL.n447 VTAIL.n387 171.744
R349 VTAIL.n447 VTAIL.n446 171.744
R350 VTAIL.n446 VTAIL.n388 171.744
R351 VTAIL.n439 VTAIL.n388 171.744
R352 VTAIL.n439 VTAIL.n438 171.744
R353 VTAIL.n438 VTAIL.n392 171.744
R354 VTAIL.n431 VTAIL.n392 171.744
R355 VTAIL.n431 VTAIL.n430 171.744
R356 VTAIL.n430 VTAIL.n396 171.744
R357 VTAIL.n423 VTAIL.n396 171.744
R358 VTAIL.n423 VTAIL.n422 171.744
R359 VTAIL.n422 VTAIL.n400 171.744
R360 VTAIL.n415 VTAIL.n400 171.744
R361 VTAIL.n415 VTAIL.n414 171.744
R362 VTAIL.n414 VTAIL.n404 171.744
R363 VTAIL.n407 VTAIL.n404 171.744
R364 VTAIL.n370 VTAIL.n369 171.744
R365 VTAIL.n369 VTAIL.n285 171.744
R366 VTAIL.n362 VTAIL.n285 171.744
R367 VTAIL.n362 VTAIL.n361 171.744
R368 VTAIL.n361 VTAIL.n289 171.744
R369 VTAIL.n293 VTAIL.n289 171.744
R370 VTAIL.n353 VTAIL.n293 171.744
R371 VTAIL.n353 VTAIL.n352 171.744
R372 VTAIL.n352 VTAIL.n294 171.744
R373 VTAIL.n345 VTAIL.n294 171.744
R374 VTAIL.n345 VTAIL.n344 171.744
R375 VTAIL.n344 VTAIL.n298 171.744
R376 VTAIL.n337 VTAIL.n298 171.744
R377 VTAIL.n337 VTAIL.n336 171.744
R378 VTAIL.n336 VTAIL.n302 171.744
R379 VTAIL.n329 VTAIL.n302 171.744
R380 VTAIL.n329 VTAIL.n328 171.744
R381 VTAIL.n328 VTAIL.n306 171.744
R382 VTAIL.n321 VTAIL.n306 171.744
R383 VTAIL.n321 VTAIL.n320 171.744
R384 VTAIL.n320 VTAIL.n310 171.744
R385 VTAIL.n313 VTAIL.n310 171.744
R386 VTAIL.n688 VTAIL.t2 85.8723
R387 VTAIL.n30 VTAIL.t0 85.8723
R388 VTAIL.n124 VTAIL.t5 85.8723
R389 VTAIL.n218 VTAIL.t4 85.8723
R390 VTAIL.n595 VTAIL.t7 85.8723
R391 VTAIL.n501 VTAIL.t6 85.8723
R392 VTAIL.n407 VTAIL.t1 85.8723
R393 VTAIL.n313 VTAIL.t3 85.8723
R394 VTAIL.n751 VTAIL.n750 33.7369
R395 VTAIL.n93 VTAIL.n92 33.7369
R396 VTAIL.n187 VTAIL.n186 33.7369
R397 VTAIL.n281 VTAIL.n280 33.7369
R398 VTAIL.n657 VTAIL.n656 33.7369
R399 VTAIL.n563 VTAIL.n562 33.7369
R400 VTAIL.n469 VTAIL.n468 33.7369
R401 VTAIL.n375 VTAIL.n374 33.7369
R402 VTAIL.n751 VTAIL.n657 27.5824
R403 VTAIL.n375 VTAIL.n281 27.5824
R404 VTAIL.n689 VTAIL.n687 16.3895
R405 VTAIL.n31 VTAIL.n29 16.3895
R406 VTAIL.n125 VTAIL.n123 16.3895
R407 VTAIL.n219 VTAIL.n217 16.3895
R408 VTAIL.n596 VTAIL.n594 16.3895
R409 VTAIL.n502 VTAIL.n500 16.3895
R410 VTAIL.n408 VTAIL.n406 16.3895
R411 VTAIL.n314 VTAIL.n312 16.3895
R412 VTAIL.n736 VTAIL.n735 13.1884
R413 VTAIL.n78 VTAIL.n77 13.1884
R414 VTAIL.n172 VTAIL.n171 13.1884
R415 VTAIL.n266 VTAIL.n265 13.1884
R416 VTAIL.n642 VTAIL.n641 13.1884
R417 VTAIL.n548 VTAIL.n547 13.1884
R418 VTAIL.n454 VTAIL.n453 13.1884
R419 VTAIL.n360 VTAIL.n359 13.1884
R420 VTAIL.n690 VTAIL.n686 12.8005
R421 VTAIL.n734 VTAIL.n666 12.8005
R422 VTAIL.n739 VTAIL.n664 12.8005
R423 VTAIL.n32 VTAIL.n28 12.8005
R424 VTAIL.n76 VTAIL.n8 12.8005
R425 VTAIL.n81 VTAIL.n6 12.8005
R426 VTAIL.n126 VTAIL.n122 12.8005
R427 VTAIL.n170 VTAIL.n102 12.8005
R428 VTAIL.n175 VTAIL.n100 12.8005
R429 VTAIL.n220 VTAIL.n216 12.8005
R430 VTAIL.n264 VTAIL.n196 12.8005
R431 VTAIL.n269 VTAIL.n194 12.8005
R432 VTAIL.n645 VTAIL.n570 12.8005
R433 VTAIL.n640 VTAIL.n572 12.8005
R434 VTAIL.n597 VTAIL.n593 12.8005
R435 VTAIL.n551 VTAIL.n476 12.8005
R436 VTAIL.n546 VTAIL.n478 12.8005
R437 VTAIL.n503 VTAIL.n499 12.8005
R438 VTAIL.n457 VTAIL.n382 12.8005
R439 VTAIL.n452 VTAIL.n384 12.8005
R440 VTAIL.n409 VTAIL.n405 12.8005
R441 VTAIL.n363 VTAIL.n288 12.8005
R442 VTAIL.n358 VTAIL.n290 12.8005
R443 VTAIL.n315 VTAIL.n311 12.8005
R444 VTAIL.n694 VTAIL.n693 12.0247
R445 VTAIL.n731 VTAIL.n730 12.0247
R446 VTAIL.n740 VTAIL.n662 12.0247
R447 VTAIL.n36 VTAIL.n35 12.0247
R448 VTAIL.n73 VTAIL.n72 12.0247
R449 VTAIL.n82 VTAIL.n4 12.0247
R450 VTAIL.n130 VTAIL.n129 12.0247
R451 VTAIL.n167 VTAIL.n166 12.0247
R452 VTAIL.n176 VTAIL.n98 12.0247
R453 VTAIL.n224 VTAIL.n223 12.0247
R454 VTAIL.n261 VTAIL.n260 12.0247
R455 VTAIL.n270 VTAIL.n192 12.0247
R456 VTAIL.n646 VTAIL.n568 12.0247
R457 VTAIL.n637 VTAIL.n636 12.0247
R458 VTAIL.n601 VTAIL.n600 12.0247
R459 VTAIL.n552 VTAIL.n474 12.0247
R460 VTAIL.n543 VTAIL.n542 12.0247
R461 VTAIL.n507 VTAIL.n506 12.0247
R462 VTAIL.n458 VTAIL.n380 12.0247
R463 VTAIL.n449 VTAIL.n448 12.0247
R464 VTAIL.n413 VTAIL.n412 12.0247
R465 VTAIL.n364 VTAIL.n286 12.0247
R466 VTAIL.n355 VTAIL.n354 12.0247
R467 VTAIL.n319 VTAIL.n318 12.0247
R468 VTAIL.n697 VTAIL.n684 11.249
R469 VTAIL.n726 VTAIL.n668 11.249
R470 VTAIL.n744 VTAIL.n743 11.249
R471 VTAIL.n39 VTAIL.n26 11.249
R472 VTAIL.n68 VTAIL.n10 11.249
R473 VTAIL.n86 VTAIL.n85 11.249
R474 VTAIL.n133 VTAIL.n120 11.249
R475 VTAIL.n162 VTAIL.n104 11.249
R476 VTAIL.n180 VTAIL.n179 11.249
R477 VTAIL.n227 VTAIL.n214 11.249
R478 VTAIL.n256 VTAIL.n198 11.249
R479 VTAIL.n274 VTAIL.n273 11.249
R480 VTAIL.n650 VTAIL.n649 11.249
R481 VTAIL.n633 VTAIL.n574 11.249
R482 VTAIL.n604 VTAIL.n591 11.249
R483 VTAIL.n556 VTAIL.n555 11.249
R484 VTAIL.n539 VTAIL.n480 11.249
R485 VTAIL.n510 VTAIL.n497 11.249
R486 VTAIL.n462 VTAIL.n461 11.249
R487 VTAIL.n445 VTAIL.n386 11.249
R488 VTAIL.n416 VTAIL.n403 11.249
R489 VTAIL.n368 VTAIL.n367 11.249
R490 VTAIL.n351 VTAIL.n292 11.249
R491 VTAIL.n322 VTAIL.n309 11.249
R492 VTAIL.n698 VTAIL.n682 10.4732
R493 VTAIL.n725 VTAIL.n670 10.4732
R494 VTAIL.n747 VTAIL.n660 10.4732
R495 VTAIL.n40 VTAIL.n24 10.4732
R496 VTAIL.n67 VTAIL.n12 10.4732
R497 VTAIL.n89 VTAIL.n2 10.4732
R498 VTAIL.n134 VTAIL.n118 10.4732
R499 VTAIL.n161 VTAIL.n106 10.4732
R500 VTAIL.n183 VTAIL.n96 10.4732
R501 VTAIL.n228 VTAIL.n212 10.4732
R502 VTAIL.n255 VTAIL.n200 10.4732
R503 VTAIL.n277 VTAIL.n190 10.4732
R504 VTAIL.n653 VTAIL.n566 10.4732
R505 VTAIL.n632 VTAIL.n577 10.4732
R506 VTAIL.n605 VTAIL.n589 10.4732
R507 VTAIL.n559 VTAIL.n472 10.4732
R508 VTAIL.n538 VTAIL.n483 10.4732
R509 VTAIL.n511 VTAIL.n495 10.4732
R510 VTAIL.n465 VTAIL.n378 10.4732
R511 VTAIL.n444 VTAIL.n389 10.4732
R512 VTAIL.n417 VTAIL.n401 10.4732
R513 VTAIL.n371 VTAIL.n284 10.4732
R514 VTAIL.n350 VTAIL.n295 10.4732
R515 VTAIL.n323 VTAIL.n307 10.4732
R516 VTAIL.n702 VTAIL.n701 9.69747
R517 VTAIL.n722 VTAIL.n721 9.69747
R518 VTAIL.n748 VTAIL.n658 9.69747
R519 VTAIL.n44 VTAIL.n43 9.69747
R520 VTAIL.n64 VTAIL.n63 9.69747
R521 VTAIL.n90 VTAIL.n0 9.69747
R522 VTAIL.n138 VTAIL.n137 9.69747
R523 VTAIL.n158 VTAIL.n157 9.69747
R524 VTAIL.n184 VTAIL.n94 9.69747
R525 VTAIL.n232 VTAIL.n231 9.69747
R526 VTAIL.n252 VTAIL.n251 9.69747
R527 VTAIL.n278 VTAIL.n188 9.69747
R528 VTAIL.n654 VTAIL.n564 9.69747
R529 VTAIL.n629 VTAIL.n628 9.69747
R530 VTAIL.n609 VTAIL.n608 9.69747
R531 VTAIL.n560 VTAIL.n470 9.69747
R532 VTAIL.n535 VTAIL.n534 9.69747
R533 VTAIL.n515 VTAIL.n514 9.69747
R534 VTAIL.n466 VTAIL.n376 9.69747
R535 VTAIL.n441 VTAIL.n440 9.69747
R536 VTAIL.n421 VTAIL.n420 9.69747
R537 VTAIL.n372 VTAIL.n282 9.69747
R538 VTAIL.n347 VTAIL.n346 9.69747
R539 VTAIL.n327 VTAIL.n326 9.69747
R540 VTAIL.n750 VTAIL.n749 9.45567
R541 VTAIL.n92 VTAIL.n91 9.45567
R542 VTAIL.n186 VTAIL.n185 9.45567
R543 VTAIL.n280 VTAIL.n279 9.45567
R544 VTAIL.n656 VTAIL.n655 9.45567
R545 VTAIL.n562 VTAIL.n561 9.45567
R546 VTAIL.n468 VTAIL.n467 9.45567
R547 VTAIL.n374 VTAIL.n373 9.45567
R548 VTAIL.n749 VTAIL.n748 9.3005
R549 VTAIL.n660 VTAIL.n659 9.3005
R550 VTAIL.n743 VTAIL.n742 9.3005
R551 VTAIL.n741 VTAIL.n740 9.3005
R552 VTAIL.n664 VTAIL.n663 9.3005
R553 VTAIL.n709 VTAIL.n708 9.3005
R554 VTAIL.n707 VTAIL.n706 9.3005
R555 VTAIL.n680 VTAIL.n679 9.3005
R556 VTAIL.n701 VTAIL.n700 9.3005
R557 VTAIL.n699 VTAIL.n698 9.3005
R558 VTAIL.n684 VTAIL.n683 9.3005
R559 VTAIL.n693 VTAIL.n692 9.3005
R560 VTAIL.n691 VTAIL.n690 9.3005
R561 VTAIL.n676 VTAIL.n675 9.3005
R562 VTAIL.n715 VTAIL.n714 9.3005
R563 VTAIL.n717 VTAIL.n716 9.3005
R564 VTAIL.n672 VTAIL.n671 9.3005
R565 VTAIL.n723 VTAIL.n722 9.3005
R566 VTAIL.n725 VTAIL.n724 9.3005
R567 VTAIL.n668 VTAIL.n667 9.3005
R568 VTAIL.n732 VTAIL.n731 9.3005
R569 VTAIL.n734 VTAIL.n733 9.3005
R570 VTAIL.n91 VTAIL.n90 9.3005
R571 VTAIL.n2 VTAIL.n1 9.3005
R572 VTAIL.n85 VTAIL.n84 9.3005
R573 VTAIL.n83 VTAIL.n82 9.3005
R574 VTAIL.n6 VTAIL.n5 9.3005
R575 VTAIL.n51 VTAIL.n50 9.3005
R576 VTAIL.n49 VTAIL.n48 9.3005
R577 VTAIL.n22 VTAIL.n21 9.3005
R578 VTAIL.n43 VTAIL.n42 9.3005
R579 VTAIL.n41 VTAIL.n40 9.3005
R580 VTAIL.n26 VTAIL.n25 9.3005
R581 VTAIL.n35 VTAIL.n34 9.3005
R582 VTAIL.n33 VTAIL.n32 9.3005
R583 VTAIL.n18 VTAIL.n17 9.3005
R584 VTAIL.n57 VTAIL.n56 9.3005
R585 VTAIL.n59 VTAIL.n58 9.3005
R586 VTAIL.n14 VTAIL.n13 9.3005
R587 VTAIL.n65 VTAIL.n64 9.3005
R588 VTAIL.n67 VTAIL.n66 9.3005
R589 VTAIL.n10 VTAIL.n9 9.3005
R590 VTAIL.n74 VTAIL.n73 9.3005
R591 VTAIL.n76 VTAIL.n75 9.3005
R592 VTAIL.n185 VTAIL.n184 9.3005
R593 VTAIL.n96 VTAIL.n95 9.3005
R594 VTAIL.n179 VTAIL.n178 9.3005
R595 VTAIL.n177 VTAIL.n176 9.3005
R596 VTAIL.n100 VTAIL.n99 9.3005
R597 VTAIL.n145 VTAIL.n144 9.3005
R598 VTAIL.n143 VTAIL.n142 9.3005
R599 VTAIL.n116 VTAIL.n115 9.3005
R600 VTAIL.n137 VTAIL.n136 9.3005
R601 VTAIL.n135 VTAIL.n134 9.3005
R602 VTAIL.n120 VTAIL.n119 9.3005
R603 VTAIL.n129 VTAIL.n128 9.3005
R604 VTAIL.n127 VTAIL.n126 9.3005
R605 VTAIL.n112 VTAIL.n111 9.3005
R606 VTAIL.n151 VTAIL.n150 9.3005
R607 VTAIL.n153 VTAIL.n152 9.3005
R608 VTAIL.n108 VTAIL.n107 9.3005
R609 VTAIL.n159 VTAIL.n158 9.3005
R610 VTAIL.n161 VTAIL.n160 9.3005
R611 VTAIL.n104 VTAIL.n103 9.3005
R612 VTAIL.n168 VTAIL.n167 9.3005
R613 VTAIL.n170 VTAIL.n169 9.3005
R614 VTAIL.n279 VTAIL.n278 9.3005
R615 VTAIL.n190 VTAIL.n189 9.3005
R616 VTAIL.n273 VTAIL.n272 9.3005
R617 VTAIL.n271 VTAIL.n270 9.3005
R618 VTAIL.n194 VTAIL.n193 9.3005
R619 VTAIL.n239 VTAIL.n238 9.3005
R620 VTAIL.n237 VTAIL.n236 9.3005
R621 VTAIL.n210 VTAIL.n209 9.3005
R622 VTAIL.n231 VTAIL.n230 9.3005
R623 VTAIL.n229 VTAIL.n228 9.3005
R624 VTAIL.n214 VTAIL.n213 9.3005
R625 VTAIL.n223 VTAIL.n222 9.3005
R626 VTAIL.n221 VTAIL.n220 9.3005
R627 VTAIL.n206 VTAIL.n205 9.3005
R628 VTAIL.n245 VTAIL.n244 9.3005
R629 VTAIL.n247 VTAIL.n246 9.3005
R630 VTAIL.n202 VTAIL.n201 9.3005
R631 VTAIL.n253 VTAIL.n252 9.3005
R632 VTAIL.n255 VTAIL.n254 9.3005
R633 VTAIL.n198 VTAIL.n197 9.3005
R634 VTAIL.n262 VTAIL.n261 9.3005
R635 VTAIL.n264 VTAIL.n263 9.3005
R636 VTAIL.n622 VTAIL.n621 9.3005
R637 VTAIL.n624 VTAIL.n623 9.3005
R638 VTAIL.n579 VTAIL.n578 9.3005
R639 VTAIL.n630 VTAIL.n629 9.3005
R640 VTAIL.n632 VTAIL.n631 9.3005
R641 VTAIL.n574 VTAIL.n573 9.3005
R642 VTAIL.n638 VTAIL.n637 9.3005
R643 VTAIL.n640 VTAIL.n639 9.3005
R644 VTAIL.n655 VTAIL.n654 9.3005
R645 VTAIL.n566 VTAIL.n565 9.3005
R646 VTAIL.n649 VTAIL.n648 9.3005
R647 VTAIL.n647 VTAIL.n646 9.3005
R648 VTAIL.n570 VTAIL.n569 9.3005
R649 VTAIL.n583 VTAIL.n582 9.3005
R650 VTAIL.n616 VTAIL.n615 9.3005
R651 VTAIL.n614 VTAIL.n613 9.3005
R652 VTAIL.n587 VTAIL.n586 9.3005
R653 VTAIL.n608 VTAIL.n607 9.3005
R654 VTAIL.n606 VTAIL.n605 9.3005
R655 VTAIL.n591 VTAIL.n590 9.3005
R656 VTAIL.n600 VTAIL.n599 9.3005
R657 VTAIL.n598 VTAIL.n597 9.3005
R658 VTAIL.n528 VTAIL.n527 9.3005
R659 VTAIL.n530 VTAIL.n529 9.3005
R660 VTAIL.n485 VTAIL.n484 9.3005
R661 VTAIL.n536 VTAIL.n535 9.3005
R662 VTAIL.n538 VTAIL.n537 9.3005
R663 VTAIL.n480 VTAIL.n479 9.3005
R664 VTAIL.n544 VTAIL.n543 9.3005
R665 VTAIL.n546 VTAIL.n545 9.3005
R666 VTAIL.n561 VTAIL.n560 9.3005
R667 VTAIL.n472 VTAIL.n471 9.3005
R668 VTAIL.n555 VTAIL.n554 9.3005
R669 VTAIL.n553 VTAIL.n552 9.3005
R670 VTAIL.n476 VTAIL.n475 9.3005
R671 VTAIL.n489 VTAIL.n488 9.3005
R672 VTAIL.n522 VTAIL.n521 9.3005
R673 VTAIL.n520 VTAIL.n519 9.3005
R674 VTAIL.n493 VTAIL.n492 9.3005
R675 VTAIL.n514 VTAIL.n513 9.3005
R676 VTAIL.n512 VTAIL.n511 9.3005
R677 VTAIL.n497 VTAIL.n496 9.3005
R678 VTAIL.n506 VTAIL.n505 9.3005
R679 VTAIL.n504 VTAIL.n503 9.3005
R680 VTAIL.n434 VTAIL.n433 9.3005
R681 VTAIL.n436 VTAIL.n435 9.3005
R682 VTAIL.n391 VTAIL.n390 9.3005
R683 VTAIL.n442 VTAIL.n441 9.3005
R684 VTAIL.n444 VTAIL.n443 9.3005
R685 VTAIL.n386 VTAIL.n385 9.3005
R686 VTAIL.n450 VTAIL.n449 9.3005
R687 VTAIL.n452 VTAIL.n451 9.3005
R688 VTAIL.n467 VTAIL.n466 9.3005
R689 VTAIL.n378 VTAIL.n377 9.3005
R690 VTAIL.n461 VTAIL.n460 9.3005
R691 VTAIL.n459 VTAIL.n458 9.3005
R692 VTAIL.n382 VTAIL.n381 9.3005
R693 VTAIL.n395 VTAIL.n394 9.3005
R694 VTAIL.n428 VTAIL.n427 9.3005
R695 VTAIL.n426 VTAIL.n425 9.3005
R696 VTAIL.n399 VTAIL.n398 9.3005
R697 VTAIL.n420 VTAIL.n419 9.3005
R698 VTAIL.n418 VTAIL.n417 9.3005
R699 VTAIL.n403 VTAIL.n402 9.3005
R700 VTAIL.n412 VTAIL.n411 9.3005
R701 VTAIL.n410 VTAIL.n409 9.3005
R702 VTAIL.n340 VTAIL.n339 9.3005
R703 VTAIL.n342 VTAIL.n341 9.3005
R704 VTAIL.n297 VTAIL.n296 9.3005
R705 VTAIL.n348 VTAIL.n347 9.3005
R706 VTAIL.n350 VTAIL.n349 9.3005
R707 VTAIL.n292 VTAIL.n291 9.3005
R708 VTAIL.n356 VTAIL.n355 9.3005
R709 VTAIL.n358 VTAIL.n357 9.3005
R710 VTAIL.n373 VTAIL.n372 9.3005
R711 VTAIL.n284 VTAIL.n283 9.3005
R712 VTAIL.n367 VTAIL.n366 9.3005
R713 VTAIL.n365 VTAIL.n364 9.3005
R714 VTAIL.n288 VTAIL.n287 9.3005
R715 VTAIL.n301 VTAIL.n300 9.3005
R716 VTAIL.n334 VTAIL.n333 9.3005
R717 VTAIL.n332 VTAIL.n331 9.3005
R718 VTAIL.n305 VTAIL.n304 9.3005
R719 VTAIL.n326 VTAIL.n325 9.3005
R720 VTAIL.n324 VTAIL.n323 9.3005
R721 VTAIL.n309 VTAIL.n308 9.3005
R722 VTAIL.n318 VTAIL.n317 9.3005
R723 VTAIL.n316 VTAIL.n315 9.3005
R724 VTAIL.n705 VTAIL.n680 8.92171
R725 VTAIL.n718 VTAIL.n672 8.92171
R726 VTAIL.n47 VTAIL.n22 8.92171
R727 VTAIL.n60 VTAIL.n14 8.92171
R728 VTAIL.n141 VTAIL.n116 8.92171
R729 VTAIL.n154 VTAIL.n108 8.92171
R730 VTAIL.n235 VTAIL.n210 8.92171
R731 VTAIL.n248 VTAIL.n202 8.92171
R732 VTAIL.n625 VTAIL.n579 8.92171
R733 VTAIL.n612 VTAIL.n587 8.92171
R734 VTAIL.n531 VTAIL.n485 8.92171
R735 VTAIL.n518 VTAIL.n493 8.92171
R736 VTAIL.n437 VTAIL.n391 8.92171
R737 VTAIL.n424 VTAIL.n399 8.92171
R738 VTAIL.n343 VTAIL.n297 8.92171
R739 VTAIL.n330 VTAIL.n305 8.92171
R740 VTAIL.n706 VTAIL.n678 8.14595
R741 VTAIL.n717 VTAIL.n674 8.14595
R742 VTAIL.n48 VTAIL.n20 8.14595
R743 VTAIL.n59 VTAIL.n16 8.14595
R744 VTAIL.n142 VTAIL.n114 8.14595
R745 VTAIL.n153 VTAIL.n110 8.14595
R746 VTAIL.n236 VTAIL.n208 8.14595
R747 VTAIL.n247 VTAIL.n204 8.14595
R748 VTAIL.n624 VTAIL.n581 8.14595
R749 VTAIL.n613 VTAIL.n585 8.14595
R750 VTAIL.n530 VTAIL.n487 8.14595
R751 VTAIL.n519 VTAIL.n491 8.14595
R752 VTAIL.n436 VTAIL.n393 8.14595
R753 VTAIL.n425 VTAIL.n397 8.14595
R754 VTAIL.n342 VTAIL.n299 8.14595
R755 VTAIL.n331 VTAIL.n303 8.14595
R756 VTAIL.n710 VTAIL.n709 7.3702
R757 VTAIL.n714 VTAIL.n713 7.3702
R758 VTAIL.n52 VTAIL.n51 7.3702
R759 VTAIL.n56 VTAIL.n55 7.3702
R760 VTAIL.n146 VTAIL.n145 7.3702
R761 VTAIL.n150 VTAIL.n149 7.3702
R762 VTAIL.n240 VTAIL.n239 7.3702
R763 VTAIL.n244 VTAIL.n243 7.3702
R764 VTAIL.n621 VTAIL.n620 7.3702
R765 VTAIL.n617 VTAIL.n616 7.3702
R766 VTAIL.n527 VTAIL.n526 7.3702
R767 VTAIL.n523 VTAIL.n522 7.3702
R768 VTAIL.n433 VTAIL.n432 7.3702
R769 VTAIL.n429 VTAIL.n428 7.3702
R770 VTAIL.n339 VTAIL.n338 7.3702
R771 VTAIL.n335 VTAIL.n334 7.3702
R772 VTAIL.n710 VTAIL.n676 6.59444
R773 VTAIL.n713 VTAIL.n676 6.59444
R774 VTAIL.n52 VTAIL.n18 6.59444
R775 VTAIL.n55 VTAIL.n18 6.59444
R776 VTAIL.n146 VTAIL.n112 6.59444
R777 VTAIL.n149 VTAIL.n112 6.59444
R778 VTAIL.n240 VTAIL.n206 6.59444
R779 VTAIL.n243 VTAIL.n206 6.59444
R780 VTAIL.n620 VTAIL.n583 6.59444
R781 VTAIL.n617 VTAIL.n583 6.59444
R782 VTAIL.n526 VTAIL.n489 6.59444
R783 VTAIL.n523 VTAIL.n489 6.59444
R784 VTAIL.n432 VTAIL.n395 6.59444
R785 VTAIL.n429 VTAIL.n395 6.59444
R786 VTAIL.n338 VTAIL.n301 6.59444
R787 VTAIL.n335 VTAIL.n301 6.59444
R788 VTAIL.n709 VTAIL.n678 5.81868
R789 VTAIL.n714 VTAIL.n674 5.81868
R790 VTAIL.n51 VTAIL.n20 5.81868
R791 VTAIL.n56 VTAIL.n16 5.81868
R792 VTAIL.n145 VTAIL.n114 5.81868
R793 VTAIL.n150 VTAIL.n110 5.81868
R794 VTAIL.n239 VTAIL.n208 5.81868
R795 VTAIL.n244 VTAIL.n204 5.81868
R796 VTAIL.n621 VTAIL.n581 5.81868
R797 VTAIL.n616 VTAIL.n585 5.81868
R798 VTAIL.n527 VTAIL.n487 5.81868
R799 VTAIL.n522 VTAIL.n491 5.81868
R800 VTAIL.n433 VTAIL.n393 5.81868
R801 VTAIL.n428 VTAIL.n397 5.81868
R802 VTAIL.n339 VTAIL.n299 5.81868
R803 VTAIL.n334 VTAIL.n303 5.81868
R804 VTAIL.n706 VTAIL.n705 5.04292
R805 VTAIL.n718 VTAIL.n717 5.04292
R806 VTAIL.n48 VTAIL.n47 5.04292
R807 VTAIL.n60 VTAIL.n59 5.04292
R808 VTAIL.n142 VTAIL.n141 5.04292
R809 VTAIL.n154 VTAIL.n153 5.04292
R810 VTAIL.n236 VTAIL.n235 5.04292
R811 VTAIL.n248 VTAIL.n247 5.04292
R812 VTAIL.n625 VTAIL.n624 5.04292
R813 VTAIL.n613 VTAIL.n612 5.04292
R814 VTAIL.n531 VTAIL.n530 5.04292
R815 VTAIL.n519 VTAIL.n518 5.04292
R816 VTAIL.n437 VTAIL.n436 5.04292
R817 VTAIL.n425 VTAIL.n424 5.04292
R818 VTAIL.n343 VTAIL.n342 5.04292
R819 VTAIL.n331 VTAIL.n330 5.04292
R820 VTAIL.n702 VTAIL.n680 4.26717
R821 VTAIL.n721 VTAIL.n672 4.26717
R822 VTAIL.n750 VTAIL.n658 4.26717
R823 VTAIL.n44 VTAIL.n22 4.26717
R824 VTAIL.n63 VTAIL.n14 4.26717
R825 VTAIL.n92 VTAIL.n0 4.26717
R826 VTAIL.n138 VTAIL.n116 4.26717
R827 VTAIL.n157 VTAIL.n108 4.26717
R828 VTAIL.n186 VTAIL.n94 4.26717
R829 VTAIL.n232 VTAIL.n210 4.26717
R830 VTAIL.n251 VTAIL.n202 4.26717
R831 VTAIL.n280 VTAIL.n188 4.26717
R832 VTAIL.n656 VTAIL.n564 4.26717
R833 VTAIL.n628 VTAIL.n579 4.26717
R834 VTAIL.n609 VTAIL.n587 4.26717
R835 VTAIL.n562 VTAIL.n470 4.26717
R836 VTAIL.n534 VTAIL.n485 4.26717
R837 VTAIL.n515 VTAIL.n493 4.26717
R838 VTAIL.n468 VTAIL.n376 4.26717
R839 VTAIL.n440 VTAIL.n391 4.26717
R840 VTAIL.n421 VTAIL.n399 4.26717
R841 VTAIL.n374 VTAIL.n282 4.26717
R842 VTAIL.n346 VTAIL.n297 4.26717
R843 VTAIL.n327 VTAIL.n305 4.26717
R844 VTAIL.n691 VTAIL.n687 3.70982
R845 VTAIL.n33 VTAIL.n29 3.70982
R846 VTAIL.n127 VTAIL.n123 3.70982
R847 VTAIL.n221 VTAIL.n217 3.70982
R848 VTAIL.n598 VTAIL.n594 3.70982
R849 VTAIL.n504 VTAIL.n500 3.70982
R850 VTAIL.n410 VTAIL.n406 3.70982
R851 VTAIL.n316 VTAIL.n312 3.70982
R852 VTAIL.n701 VTAIL.n682 3.49141
R853 VTAIL.n722 VTAIL.n670 3.49141
R854 VTAIL.n748 VTAIL.n747 3.49141
R855 VTAIL.n43 VTAIL.n24 3.49141
R856 VTAIL.n64 VTAIL.n12 3.49141
R857 VTAIL.n90 VTAIL.n89 3.49141
R858 VTAIL.n137 VTAIL.n118 3.49141
R859 VTAIL.n158 VTAIL.n106 3.49141
R860 VTAIL.n184 VTAIL.n183 3.49141
R861 VTAIL.n231 VTAIL.n212 3.49141
R862 VTAIL.n252 VTAIL.n200 3.49141
R863 VTAIL.n278 VTAIL.n277 3.49141
R864 VTAIL.n654 VTAIL.n653 3.49141
R865 VTAIL.n629 VTAIL.n577 3.49141
R866 VTAIL.n608 VTAIL.n589 3.49141
R867 VTAIL.n560 VTAIL.n559 3.49141
R868 VTAIL.n535 VTAIL.n483 3.49141
R869 VTAIL.n514 VTAIL.n495 3.49141
R870 VTAIL.n466 VTAIL.n465 3.49141
R871 VTAIL.n441 VTAIL.n389 3.49141
R872 VTAIL.n420 VTAIL.n401 3.49141
R873 VTAIL.n372 VTAIL.n371 3.49141
R874 VTAIL.n347 VTAIL.n295 3.49141
R875 VTAIL.n326 VTAIL.n307 3.49141
R876 VTAIL.n698 VTAIL.n697 2.71565
R877 VTAIL.n726 VTAIL.n725 2.71565
R878 VTAIL.n744 VTAIL.n660 2.71565
R879 VTAIL.n40 VTAIL.n39 2.71565
R880 VTAIL.n68 VTAIL.n67 2.71565
R881 VTAIL.n86 VTAIL.n2 2.71565
R882 VTAIL.n134 VTAIL.n133 2.71565
R883 VTAIL.n162 VTAIL.n161 2.71565
R884 VTAIL.n180 VTAIL.n96 2.71565
R885 VTAIL.n228 VTAIL.n227 2.71565
R886 VTAIL.n256 VTAIL.n255 2.71565
R887 VTAIL.n274 VTAIL.n190 2.71565
R888 VTAIL.n650 VTAIL.n566 2.71565
R889 VTAIL.n633 VTAIL.n632 2.71565
R890 VTAIL.n605 VTAIL.n604 2.71565
R891 VTAIL.n556 VTAIL.n472 2.71565
R892 VTAIL.n539 VTAIL.n538 2.71565
R893 VTAIL.n511 VTAIL.n510 2.71565
R894 VTAIL.n462 VTAIL.n378 2.71565
R895 VTAIL.n445 VTAIL.n444 2.71565
R896 VTAIL.n417 VTAIL.n416 2.71565
R897 VTAIL.n368 VTAIL.n284 2.71565
R898 VTAIL.n351 VTAIL.n350 2.71565
R899 VTAIL.n323 VTAIL.n322 2.71565
R900 VTAIL.n694 VTAIL.n684 1.93989
R901 VTAIL.n730 VTAIL.n668 1.93989
R902 VTAIL.n743 VTAIL.n662 1.93989
R903 VTAIL.n36 VTAIL.n26 1.93989
R904 VTAIL.n72 VTAIL.n10 1.93989
R905 VTAIL.n85 VTAIL.n4 1.93989
R906 VTAIL.n130 VTAIL.n120 1.93989
R907 VTAIL.n166 VTAIL.n104 1.93989
R908 VTAIL.n179 VTAIL.n98 1.93989
R909 VTAIL.n224 VTAIL.n214 1.93989
R910 VTAIL.n260 VTAIL.n198 1.93989
R911 VTAIL.n273 VTAIL.n192 1.93989
R912 VTAIL.n649 VTAIL.n568 1.93989
R913 VTAIL.n636 VTAIL.n574 1.93989
R914 VTAIL.n601 VTAIL.n591 1.93989
R915 VTAIL.n555 VTAIL.n474 1.93989
R916 VTAIL.n542 VTAIL.n480 1.93989
R917 VTAIL.n507 VTAIL.n497 1.93989
R918 VTAIL.n461 VTAIL.n380 1.93989
R919 VTAIL.n448 VTAIL.n386 1.93989
R920 VTAIL.n413 VTAIL.n403 1.93989
R921 VTAIL.n367 VTAIL.n286 1.93989
R922 VTAIL.n354 VTAIL.n292 1.93989
R923 VTAIL.n319 VTAIL.n309 1.93989
R924 VTAIL.n693 VTAIL.n686 1.16414
R925 VTAIL.n731 VTAIL.n666 1.16414
R926 VTAIL.n740 VTAIL.n739 1.16414
R927 VTAIL.n35 VTAIL.n28 1.16414
R928 VTAIL.n73 VTAIL.n8 1.16414
R929 VTAIL.n82 VTAIL.n81 1.16414
R930 VTAIL.n129 VTAIL.n122 1.16414
R931 VTAIL.n167 VTAIL.n102 1.16414
R932 VTAIL.n176 VTAIL.n175 1.16414
R933 VTAIL.n223 VTAIL.n216 1.16414
R934 VTAIL.n261 VTAIL.n196 1.16414
R935 VTAIL.n270 VTAIL.n269 1.16414
R936 VTAIL.n646 VTAIL.n645 1.16414
R937 VTAIL.n637 VTAIL.n572 1.16414
R938 VTAIL.n600 VTAIL.n593 1.16414
R939 VTAIL.n552 VTAIL.n551 1.16414
R940 VTAIL.n543 VTAIL.n478 1.16414
R941 VTAIL.n506 VTAIL.n499 1.16414
R942 VTAIL.n458 VTAIL.n457 1.16414
R943 VTAIL.n449 VTAIL.n384 1.16414
R944 VTAIL.n412 VTAIL.n405 1.16414
R945 VTAIL.n364 VTAIL.n363 1.16414
R946 VTAIL.n355 VTAIL.n290 1.16414
R947 VTAIL.n318 VTAIL.n311 1.16414
R948 VTAIL.n469 VTAIL.n375 0.664293
R949 VTAIL.n657 VTAIL.n563 0.664293
R950 VTAIL.n281 VTAIL.n187 0.664293
R951 VTAIL.n563 VTAIL.n469 0.470328
R952 VTAIL.n187 VTAIL.n93 0.470328
R953 VTAIL VTAIL.n93 0.390586
R954 VTAIL.n690 VTAIL.n689 0.388379
R955 VTAIL.n735 VTAIL.n734 0.388379
R956 VTAIL.n736 VTAIL.n664 0.388379
R957 VTAIL.n32 VTAIL.n31 0.388379
R958 VTAIL.n77 VTAIL.n76 0.388379
R959 VTAIL.n78 VTAIL.n6 0.388379
R960 VTAIL.n126 VTAIL.n125 0.388379
R961 VTAIL.n171 VTAIL.n170 0.388379
R962 VTAIL.n172 VTAIL.n100 0.388379
R963 VTAIL.n220 VTAIL.n219 0.388379
R964 VTAIL.n265 VTAIL.n264 0.388379
R965 VTAIL.n266 VTAIL.n194 0.388379
R966 VTAIL.n642 VTAIL.n570 0.388379
R967 VTAIL.n641 VTAIL.n640 0.388379
R968 VTAIL.n597 VTAIL.n596 0.388379
R969 VTAIL.n548 VTAIL.n476 0.388379
R970 VTAIL.n547 VTAIL.n546 0.388379
R971 VTAIL.n503 VTAIL.n502 0.388379
R972 VTAIL.n454 VTAIL.n382 0.388379
R973 VTAIL.n453 VTAIL.n452 0.388379
R974 VTAIL.n409 VTAIL.n408 0.388379
R975 VTAIL.n360 VTAIL.n288 0.388379
R976 VTAIL.n359 VTAIL.n358 0.388379
R977 VTAIL.n315 VTAIL.n314 0.388379
R978 VTAIL VTAIL.n751 0.274207
R979 VTAIL.n692 VTAIL.n691 0.155672
R980 VTAIL.n692 VTAIL.n683 0.155672
R981 VTAIL.n699 VTAIL.n683 0.155672
R982 VTAIL.n700 VTAIL.n699 0.155672
R983 VTAIL.n700 VTAIL.n679 0.155672
R984 VTAIL.n707 VTAIL.n679 0.155672
R985 VTAIL.n708 VTAIL.n707 0.155672
R986 VTAIL.n708 VTAIL.n675 0.155672
R987 VTAIL.n715 VTAIL.n675 0.155672
R988 VTAIL.n716 VTAIL.n715 0.155672
R989 VTAIL.n716 VTAIL.n671 0.155672
R990 VTAIL.n723 VTAIL.n671 0.155672
R991 VTAIL.n724 VTAIL.n723 0.155672
R992 VTAIL.n724 VTAIL.n667 0.155672
R993 VTAIL.n732 VTAIL.n667 0.155672
R994 VTAIL.n733 VTAIL.n732 0.155672
R995 VTAIL.n733 VTAIL.n663 0.155672
R996 VTAIL.n741 VTAIL.n663 0.155672
R997 VTAIL.n742 VTAIL.n741 0.155672
R998 VTAIL.n742 VTAIL.n659 0.155672
R999 VTAIL.n749 VTAIL.n659 0.155672
R1000 VTAIL.n34 VTAIL.n33 0.155672
R1001 VTAIL.n34 VTAIL.n25 0.155672
R1002 VTAIL.n41 VTAIL.n25 0.155672
R1003 VTAIL.n42 VTAIL.n41 0.155672
R1004 VTAIL.n42 VTAIL.n21 0.155672
R1005 VTAIL.n49 VTAIL.n21 0.155672
R1006 VTAIL.n50 VTAIL.n49 0.155672
R1007 VTAIL.n50 VTAIL.n17 0.155672
R1008 VTAIL.n57 VTAIL.n17 0.155672
R1009 VTAIL.n58 VTAIL.n57 0.155672
R1010 VTAIL.n58 VTAIL.n13 0.155672
R1011 VTAIL.n65 VTAIL.n13 0.155672
R1012 VTAIL.n66 VTAIL.n65 0.155672
R1013 VTAIL.n66 VTAIL.n9 0.155672
R1014 VTAIL.n74 VTAIL.n9 0.155672
R1015 VTAIL.n75 VTAIL.n74 0.155672
R1016 VTAIL.n75 VTAIL.n5 0.155672
R1017 VTAIL.n83 VTAIL.n5 0.155672
R1018 VTAIL.n84 VTAIL.n83 0.155672
R1019 VTAIL.n84 VTAIL.n1 0.155672
R1020 VTAIL.n91 VTAIL.n1 0.155672
R1021 VTAIL.n128 VTAIL.n127 0.155672
R1022 VTAIL.n128 VTAIL.n119 0.155672
R1023 VTAIL.n135 VTAIL.n119 0.155672
R1024 VTAIL.n136 VTAIL.n135 0.155672
R1025 VTAIL.n136 VTAIL.n115 0.155672
R1026 VTAIL.n143 VTAIL.n115 0.155672
R1027 VTAIL.n144 VTAIL.n143 0.155672
R1028 VTAIL.n144 VTAIL.n111 0.155672
R1029 VTAIL.n151 VTAIL.n111 0.155672
R1030 VTAIL.n152 VTAIL.n151 0.155672
R1031 VTAIL.n152 VTAIL.n107 0.155672
R1032 VTAIL.n159 VTAIL.n107 0.155672
R1033 VTAIL.n160 VTAIL.n159 0.155672
R1034 VTAIL.n160 VTAIL.n103 0.155672
R1035 VTAIL.n168 VTAIL.n103 0.155672
R1036 VTAIL.n169 VTAIL.n168 0.155672
R1037 VTAIL.n169 VTAIL.n99 0.155672
R1038 VTAIL.n177 VTAIL.n99 0.155672
R1039 VTAIL.n178 VTAIL.n177 0.155672
R1040 VTAIL.n178 VTAIL.n95 0.155672
R1041 VTAIL.n185 VTAIL.n95 0.155672
R1042 VTAIL.n222 VTAIL.n221 0.155672
R1043 VTAIL.n222 VTAIL.n213 0.155672
R1044 VTAIL.n229 VTAIL.n213 0.155672
R1045 VTAIL.n230 VTAIL.n229 0.155672
R1046 VTAIL.n230 VTAIL.n209 0.155672
R1047 VTAIL.n237 VTAIL.n209 0.155672
R1048 VTAIL.n238 VTAIL.n237 0.155672
R1049 VTAIL.n238 VTAIL.n205 0.155672
R1050 VTAIL.n245 VTAIL.n205 0.155672
R1051 VTAIL.n246 VTAIL.n245 0.155672
R1052 VTAIL.n246 VTAIL.n201 0.155672
R1053 VTAIL.n253 VTAIL.n201 0.155672
R1054 VTAIL.n254 VTAIL.n253 0.155672
R1055 VTAIL.n254 VTAIL.n197 0.155672
R1056 VTAIL.n262 VTAIL.n197 0.155672
R1057 VTAIL.n263 VTAIL.n262 0.155672
R1058 VTAIL.n263 VTAIL.n193 0.155672
R1059 VTAIL.n271 VTAIL.n193 0.155672
R1060 VTAIL.n272 VTAIL.n271 0.155672
R1061 VTAIL.n272 VTAIL.n189 0.155672
R1062 VTAIL.n279 VTAIL.n189 0.155672
R1063 VTAIL.n655 VTAIL.n565 0.155672
R1064 VTAIL.n648 VTAIL.n565 0.155672
R1065 VTAIL.n648 VTAIL.n647 0.155672
R1066 VTAIL.n647 VTAIL.n569 0.155672
R1067 VTAIL.n639 VTAIL.n569 0.155672
R1068 VTAIL.n639 VTAIL.n638 0.155672
R1069 VTAIL.n638 VTAIL.n573 0.155672
R1070 VTAIL.n631 VTAIL.n573 0.155672
R1071 VTAIL.n631 VTAIL.n630 0.155672
R1072 VTAIL.n630 VTAIL.n578 0.155672
R1073 VTAIL.n623 VTAIL.n578 0.155672
R1074 VTAIL.n623 VTAIL.n622 0.155672
R1075 VTAIL.n622 VTAIL.n582 0.155672
R1076 VTAIL.n615 VTAIL.n582 0.155672
R1077 VTAIL.n615 VTAIL.n614 0.155672
R1078 VTAIL.n614 VTAIL.n586 0.155672
R1079 VTAIL.n607 VTAIL.n586 0.155672
R1080 VTAIL.n607 VTAIL.n606 0.155672
R1081 VTAIL.n606 VTAIL.n590 0.155672
R1082 VTAIL.n599 VTAIL.n590 0.155672
R1083 VTAIL.n599 VTAIL.n598 0.155672
R1084 VTAIL.n561 VTAIL.n471 0.155672
R1085 VTAIL.n554 VTAIL.n471 0.155672
R1086 VTAIL.n554 VTAIL.n553 0.155672
R1087 VTAIL.n553 VTAIL.n475 0.155672
R1088 VTAIL.n545 VTAIL.n475 0.155672
R1089 VTAIL.n545 VTAIL.n544 0.155672
R1090 VTAIL.n544 VTAIL.n479 0.155672
R1091 VTAIL.n537 VTAIL.n479 0.155672
R1092 VTAIL.n537 VTAIL.n536 0.155672
R1093 VTAIL.n536 VTAIL.n484 0.155672
R1094 VTAIL.n529 VTAIL.n484 0.155672
R1095 VTAIL.n529 VTAIL.n528 0.155672
R1096 VTAIL.n528 VTAIL.n488 0.155672
R1097 VTAIL.n521 VTAIL.n488 0.155672
R1098 VTAIL.n521 VTAIL.n520 0.155672
R1099 VTAIL.n520 VTAIL.n492 0.155672
R1100 VTAIL.n513 VTAIL.n492 0.155672
R1101 VTAIL.n513 VTAIL.n512 0.155672
R1102 VTAIL.n512 VTAIL.n496 0.155672
R1103 VTAIL.n505 VTAIL.n496 0.155672
R1104 VTAIL.n505 VTAIL.n504 0.155672
R1105 VTAIL.n467 VTAIL.n377 0.155672
R1106 VTAIL.n460 VTAIL.n377 0.155672
R1107 VTAIL.n460 VTAIL.n459 0.155672
R1108 VTAIL.n459 VTAIL.n381 0.155672
R1109 VTAIL.n451 VTAIL.n381 0.155672
R1110 VTAIL.n451 VTAIL.n450 0.155672
R1111 VTAIL.n450 VTAIL.n385 0.155672
R1112 VTAIL.n443 VTAIL.n385 0.155672
R1113 VTAIL.n443 VTAIL.n442 0.155672
R1114 VTAIL.n442 VTAIL.n390 0.155672
R1115 VTAIL.n435 VTAIL.n390 0.155672
R1116 VTAIL.n435 VTAIL.n434 0.155672
R1117 VTAIL.n434 VTAIL.n394 0.155672
R1118 VTAIL.n427 VTAIL.n394 0.155672
R1119 VTAIL.n427 VTAIL.n426 0.155672
R1120 VTAIL.n426 VTAIL.n398 0.155672
R1121 VTAIL.n419 VTAIL.n398 0.155672
R1122 VTAIL.n419 VTAIL.n418 0.155672
R1123 VTAIL.n418 VTAIL.n402 0.155672
R1124 VTAIL.n411 VTAIL.n402 0.155672
R1125 VTAIL.n411 VTAIL.n410 0.155672
R1126 VTAIL.n373 VTAIL.n283 0.155672
R1127 VTAIL.n366 VTAIL.n283 0.155672
R1128 VTAIL.n366 VTAIL.n365 0.155672
R1129 VTAIL.n365 VTAIL.n287 0.155672
R1130 VTAIL.n357 VTAIL.n287 0.155672
R1131 VTAIL.n357 VTAIL.n356 0.155672
R1132 VTAIL.n356 VTAIL.n291 0.155672
R1133 VTAIL.n349 VTAIL.n291 0.155672
R1134 VTAIL.n349 VTAIL.n348 0.155672
R1135 VTAIL.n348 VTAIL.n296 0.155672
R1136 VTAIL.n341 VTAIL.n296 0.155672
R1137 VTAIL.n341 VTAIL.n340 0.155672
R1138 VTAIL.n340 VTAIL.n300 0.155672
R1139 VTAIL.n333 VTAIL.n300 0.155672
R1140 VTAIL.n333 VTAIL.n332 0.155672
R1141 VTAIL.n332 VTAIL.n304 0.155672
R1142 VTAIL.n325 VTAIL.n304 0.155672
R1143 VTAIL.n325 VTAIL.n324 0.155672
R1144 VTAIL.n324 VTAIL.n308 0.155672
R1145 VTAIL.n317 VTAIL.n308 0.155672
R1146 VTAIL.n317 VTAIL.n316 0.155672
R1147 VDD1 VDD1.n1 111.727
R1148 VDD1 VDD1.n0 71.0016
R1149 VDD1.n0 VDD1.t0 1.92615
R1150 VDD1.n0 VDD1.t3 1.92615
R1151 VDD1.n1 VDD1.t2 1.92615
R1152 VDD1.n1 VDD1.t1 1.92615
R1153 B.n118 B.t9 1132.61
R1154 B.n126 B.t3 1132.61
R1155 B.n38 B.t0 1132.61
R1156 B.n44 B.t6 1132.61
R1157 B.n413 B.n74 585
R1158 B.n415 B.n414 585
R1159 B.n416 B.n73 585
R1160 B.n418 B.n417 585
R1161 B.n419 B.n72 585
R1162 B.n421 B.n420 585
R1163 B.n422 B.n71 585
R1164 B.n424 B.n423 585
R1165 B.n425 B.n70 585
R1166 B.n427 B.n426 585
R1167 B.n428 B.n69 585
R1168 B.n430 B.n429 585
R1169 B.n431 B.n68 585
R1170 B.n433 B.n432 585
R1171 B.n434 B.n67 585
R1172 B.n436 B.n435 585
R1173 B.n437 B.n66 585
R1174 B.n439 B.n438 585
R1175 B.n440 B.n65 585
R1176 B.n442 B.n441 585
R1177 B.n443 B.n64 585
R1178 B.n445 B.n444 585
R1179 B.n446 B.n63 585
R1180 B.n448 B.n447 585
R1181 B.n449 B.n62 585
R1182 B.n451 B.n450 585
R1183 B.n452 B.n61 585
R1184 B.n454 B.n453 585
R1185 B.n455 B.n60 585
R1186 B.n457 B.n456 585
R1187 B.n458 B.n59 585
R1188 B.n460 B.n459 585
R1189 B.n461 B.n58 585
R1190 B.n463 B.n462 585
R1191 B.n464 B.n57 585
R1192 B.n466 B.n465 585
R1193 B.n467 B.n56 585
R1194 B.n469 B.n468 585
R1195 B.n470 B.n55 585
R1196 B.n472 B.n471 585
R1197 B.n473 B.n54 585
R1198 B.n475 B.n474 585
R1199 B.n476 B.n53 585
R1200 B.n478 B.n477 585
R1201 B.n479 B.n52 585
R1202 B.n481 B.n480 585
R1203 B.n482 B.n51 585
R1204 B.n484 B.n483 585
R1205 B.n485 B.n50 585
R1206 B.n487 B.n486 585
R1207 B.n488 B.n49 585
R1208 B.n490 B.n489 585
R1209 B.n491 B.n48 585
R1210 B.n493 B.n492 585
R1211 B.n494 B.n47 585
R1212 B.n496 B.n495 585
R1213 B.n498 B.n497 585
R1214 B.n499 B.n43 585
R1215 B.n501 B.n500 585
R1216 B.n502 B.n42 585
R1217 B.n504 B.n503 585
R1218 B.n505 B.n41 585
R1219 B.n507 B.n506 585
R1220 B.n508 B.n40 585
R1221 B.n510 B.n509 585
R1222 B.n512 B.n37 585
R1223 B.n514 B.n513 585
R1224 B.n515 B.n36 585
R1225 B.n517 B.n516 585
R1226 B.n518 B.n35 585
R1227 B.n520 B.n519 585
R1228 B.n521 B.n34 585
R1229 B.n523 B.n522 585
R1230 B.n524 B.n33 585
R1231 B.n526 B.n525 585
R1232 B.n527 B.n32 585
R1233 B.n529 B.n528 585
R1234 B.n530 B.n31 585
R1235 B.n532 B.n531 585
R1236 B.n533 B.n30 585
R1237 B.n535 B.n534 585
R1238 B.n536 B.n29 585
R1239 B.n538 B.n537 585
R1240 B.n539 B.n28 585
R1241 B.n541 B.n540 585
R1242 B.n542 B.n27 585
R1243 B.n544 B.n543 585
R1244 B.n545 B.n26 585
R1245 B.n547 B.n546 585
R1246 B.n548 B.n25 585
R1247 B.n550 B.n549 585
R1248 B.n551 B.n24 585
R1249 B.n553 B.n552 585
R1250 B.n554 B.n23 585
R1251 B.n556 B.n555 585
R1252 B.n557 B.n22 585
R1253 B.n559 B.n558 585
R1254 B.n560 B.n21 585
R1255 B.n562 B.n561 585
R1256 B.n563 B.n20 585
R1257 B.n565 B.n564 585
R1258 B.n566 B.n19 585
R1259 B.n568 B.n567 585
R1260 B.n569 B.n18 585
R1261 B.n571 B.n570 585
R1262 B.n572 B.n17 585
R1263 B.n574 B.n573 585
R1264 B.n575 B.n16 585
R1265 B.n577 B.n576 585
R1266 B.n578 B.n15 585
R1267 B.n580 B.n579 585
R1268 B.n581 B.n14 585
R1269 B.n583 B.n582 585
R1270 B.n584 B.n13 585
R1271 B.n586 B.n585 585
R1272 B.n587 B.n12 585
R1273 B.n589 B.n588 585
R1274 B.n590 B.n11 585
R1275 B.n592 B.n591 585
R1276 B.n593 B.n10 585
R1277 B.n595 B.n594 585
R1278 B.n412 B.n411 585
R1279 B.n410 B.n75 585
R1280 B.n409 B.n408 585
R1281 B.n407 B.n76 585
R1282 B.n406 B.n405 585
R1283 B.n404 B.n77 585
R1284 B.n403 B.n402 585
R1285 B.n401 B.n78 585
R1286 B.n400 B.n399 585
R1287 B.n398 B.n79 585
R1288 B.n397 B.n396 585
R1289 B.n395 B.n80 585
R1290 B.n394 B.n393 585
R1291 B.n392 B.n81 585
R1292 B.n391 B.n390 585
R1293 B.n389 B.n82 585
R1294 B.n388 B.n387 585
R1295 B.n386 B.n83 585
R1296 B.n385 B.n384 585
R1297 B.n383 B.n84 585
R1298 B.n382 B.n381 585
R1299 B.n380 B.n85 585
R1300 B.n379 B.n378 585
R1301 B.n377 B.n86 585
R1302 B.n376 B.n375 585
R1303 B.n374 B.n87 585
R1304 B.n373 B.n372 585
R1305 B.n371 B.n88 585
R1306 B.n370 B.n369 585
R1307 B.n368 B.n89 585
R1308 B.n367 B.n366 585
R1309 B.n184 B.n183 585
R1310 B.n185 B.n154 585
R1311 B.n187 B.n186 585
R1312 B.n188 B.n153 585
R1313 B.n190 B.n189 585
R1314 B.n191 B.n152 585
R1315 B.n193 B.n192 585
R1316 B.n194 B.n151 585
R1317 B.n196 B.n195 585
R1318 B.n197 B.n150 585
R1319 B.n199 B.n198 585
R1320 B.n200 B.n149 585
R1321 B.n202 B.n201 585
R1322 B.n203 B.n148 585
R1323 B.n205 B.n204 585
R1324 B.n206 B.n147 585
R1325 B.n208 B.n207 585
R1326 B.n209 B.n146 585
R1327 B.n211 B.n210 585
R1328 B.n212 B.n145 585
R1329 B.n214 B.n213 585
R1330 B.n215 B.n144 585
R1331 B.n217 B.n216 585
R1332 B.n218 B.n143 585
R1333 B.n220 B.n219 585
R1334 B.n221 B.n142 585
R1335 B.n223 B.n222 585
R1336 B.n224 B.n141 585
R1337 B.n226 B.n225 585
R1338 B.n227 B.n140 585
R1339 B.n229 B.n228 585
R1340 B.n230 B.n139 585
R1341 B.n232 B.n231 585
R1342 B.n233 B.n138 585
R1343 B.n235 B.n234 585
R1344 B.n236 B.n137 585
R1345 B.n238 B.n237 585
R1346 B.n239 B.n136 585
R1347 B.n241 B.n240 585
R1348 B.n242 B.n135 585
R1349 B.n244 B.n243 585
R1350 B.n245 B.n134 585
R1351 B.n247 B.n246 585
R1352 B.n248 B.n133 585
R1353 B.n250 B.n249 585
R1354 B.n251 B.n132 585
R1355 B.n253 B.n252 585
R1356 B.n254 B.n131 585
R1357 B.n256 B.n255 585
R1358 B.n257 B.n130 585
R1359 B.n259 B.n258 585
R1360 B.n260 B.n129 585
R1361 B.n262 B.n261 585
R1362 B.n263 B.n128 585
R1363 B.n265 B.n264 585
R1364 B.n266 B.n125 585
R1365 B.n269 B.n268 585
R1366 B.n270 B.n124 585
R1367 B.n272 B.n271 585
R1368 B.n273 B.n123 585
R1369 B.n275 B.n274 585
R1370 B.n276 B.n122 585
R1371 B.n278 B.n277 585
R1372 B.n279 B.n121 585
R1373 B.n281 B.n280 585
R1374 B.n283 B.n282 585
R1375 B.n284 B.n117 585
R1376 B.n286 B.n285 585
R1377 B.n287 B.n116 585
R1378 B.n289 B.n288 585
R1379 B.n290 B.n115 585
R1380 B.n292 B.n291 585
R1381 B.n293 B.n114 585
R1382 B.n295 B.n294 585
R1383 B.n296 B.n113 585
R1384 B.n298 B.n297 585
R1385 B.n299 B.n112 585
R1386 B.n301 B.n300 585
R1387 B.n302 B.n111 585
R1388 B.n304 B.n303 585
R1389 B.n305 B.n110 585
R1390 B.n307 B.n306 585
R1391 B.n308 B.n109 585
R1392 B.n310 B.n309 585
R1393 B.n311 B.n108 585
R1394 B.n313 B.n312 585
R1395 B.n314 B.n107 585
R1396 B.n316 B.n315 585
R1397 B.n317 B.n106 585
R1398 B.n319 B.n318 585
R1399 B.n320 B.n105 585
R1400 B.n322 B.n321 585
R1401 B.n323 B.n104 585
R1402 B.n325 B.n324 585
R1403 B.n326 B.n103 585
R1404 B.n328 B.n327 585
R1405 B.n329 B.n102 585
R1406 B.n331 B.n330 585
R1407 B.n332 B.n101 585
R1408 B.n334 B.n333 585
R1409 B.n335 B.n100 585
R1410 B.n337 B.n336 585
R1411 B.n338 B.n99 585
R1412 B.n340 B.n339 585
R1413 B.n341 B.n98 585
R1414 B.n343 B.n342 585
R1415 B.n344 B.n97 585
R1416 B.n346 B.n345 585
R1417 B.n347 B.n96 585
R1418 B.n349 B.n348 585
R1419 B.n350 B.n95 585
R1420 B.n352 B.n351 585
R1421 B.n353 B.n94 585
R1422 B.n355 B.n354 585
R1423 B.n356 B.n93 585
R1424 B.n358 B.n357 585
R1425 B.n359 B.n92 585
R1426 B.n361 B.n360 585
R1427 B.n362 B.n91 585
R1428 B.n364 B.n363 585
R1429 B.n365 B.n90 585
R1430 B.n182 B.n155 585
R1431 B.n181 B.n180 585
R1432 B.n179 B.n156 585
R1433 B.n178 B.n177 585
R1434 B.n176 B.n157 585
R1435 B.n175 B.n174 585
R1436 B.n173 B.n158 585
R1437 B.n172 B.n171 585
R1438 B.n170 B.n159 585
R1439 B.n169 B.n168 585
R1440 B.n167 B.n160 585
R1441 B.n166 B.n165 585
R1442 B.n164 B.n161 585
R1443 B.n163 B.n162 585
R1444 B.n2 B.n0 585
R1445 B.n617 B.n1 585
R1446 B.n616 B.n615 585
R1447 B.n614 B.n3 585
R1448 B.n613 B.n612 585
R1449 B.n611 B.n4 585
R1450 B.n610 B.n609 585
R1451 B.n608 B.n5 585
R1452 B.n607 B.n606 585
R1453 B.n605 B.n6 585
R1454 B.n604 B.n603 585
R1455 B.n602 B.n7 585
R1456 B.n601 B.n600 585
R1457 B.n599 B.n8 585
R1458 B.n598 B.n597 585
R1459 B.n596 B.n9 585
R1460 B.n619 B.n618 585
R1461 B.n184 B.n155 526.135
R1462 B.n594 B.n9 526.135
R1463 B.n366 B.n365 526.135
R1464 B.n413 B.n412 526.135
R1465 B.n118 B.t11 478.526
R1466 B.n44 B.t7 478.526
R1467 B.n126 B.t5 478.526
R1468 B.n38 B.t1 478.526
R1469 B.n119 B.t10 463.592
R1470 B.n45 B.t8 463.592
R1471 B.n127 B.t4 463.592
R1472 B.n39 B.t2 463.592
R1473 B.n180 B.n155 163.367
R1474 B.n180 B.n179 163.367
R1475 B.n179 B.n178 163.367
R1476 B.n178 B.n157 163.367
R1477 B.n174 B.n157 163.367
R1478 B.n174 B.n173 163.367
R1479 B.n173 B.n172 163.367
R1480 B.n172 B.n159 163.367
R1481 B.n168 B.n159 163.367
R1482 B.n168 B.n167 163.367
R1483 B.n167 B.n166 163.367
R1484 B.n166 B.n161 163.367
R1485 B.n162 B.n161 163.367
R1486 B.n162 B.n2 163.367
R1487 B.n618 B.n2 163.367
R1488 B.n618 B.n617 163.367
R1489 B.n617 B.n616 163.367
R1490 B.n616 B.n3 163.367
R1491 B.n612 B.n3 163.367
R1492 B.n612 B.n611 163.367
R1493 B.n611 B.n610 163.367
R1494 B.n610 B.n5 163.367
R1495 B.n606 B.n5 163.367
R1496 B.n606 B.n605 163.367
R1497 B.n605 B.n604 163.367
R1498 B.n604 B.n7 163.367
R1499 B.n600 B.n7 163.367
R1500 B.n600 B.n599 163.367
R1501 B.n599 B.n598 163.367
R1502 B.n598 B.n9 163.367
R1503 B.n185 B.n184 163.367
R1504 B.n186 B.n185 163.367
R1505 B.n186 B.n153 163.367
R1506 B.n190 B.n153 163.367
R1507 B.n191 B.n190 163.367
R1508 B.n192 B.n191 163.367
R1509 B.n192 B.n151 163.367
R1510 B.n196 B.n151 163.367
R1511 B.n197 B.n196 163.367
R1512 B.n198 B.n197 163.367
R1513 B.n198 B.n149 163.367
R1514 B.n202 B.n149 163.367
R1515 B.n203 B.n202 163.367
R1516 B.n204 B.n203 163.367
R1517 B.n204 B.n147 163.367
R1518 B.n208 B.n147 163.367
R1519 B.n209 B.n208 163.367
R1520 B.n210 B.n209 163.367
R1521 B.n210 B.n145 163.367
R1522 B.n214 B.n145 163.367
R1523 B.n215 B.n214 163.367
R1524 B.n216 B.n215 163.367
R1525 B.n216 B.n143 163.367
R1526 B.n220 B.n143 163.367
R1527 B.n221 B.n220 163.367
R1528 B.n222 B.n221 163.367
R1529 B.n222 B.n141 163.367
R1530 B.n226 B.n141 163.367
R1531 B.n227 B.n226 163.367
R1532 B.n228 B.n227 163.367
R1533 B.n228 B.n139 163.367
R1534 B.n232 B.n139 163.367
R1535 B.n233 B.n232 163.367
R1536 B.n234 B.n233 163.367
R1537 B.n234 B.n137 163.367
R1538 B.n238 B.n137 163.367
R1539 B.n239 B.n238 163.367
R1540 B.n240 B.n239 163.367
R1541 B.n240 B.n135 163.367
R1542 B.n244 B.n135 163.367
R1543 B.n245 B.n244 163.367
R1544 B.n246 B.n245 163.367
R1545 B.n246 B.n133 163.367
R1546 B.n250 B.n133 163.367
R1547 B.n251 B.n250 163.367
R1548 B.n252 B.n251 163.367
R1549 B.n252 B.n131 163.367
R1550 B.n256 B.n131 163.367
R1551 B.n257 B.n256 163.367
R1552 B.n258 B.n257 163.367
R1553 B.n258 B.n129 163.367
R1554 B.n262 B.n129 163.367
R1555 B.n263 B.n262 163.367
R1556 B.n264 B.n263 163.367
R1557 B.n264 B.n125 163.367
R1558 B.n269 B.n125 163.367
R1559 B.n270 B.n269 163.367
R1560 B.n271 B.n270 163.367
R1561 B.n271 B.n123 163.367
R1562 B.n275 B.n123 163.367
R1563 B.n276 B.n275 163.367
R1564 B.n277 B.n276 163.367
R1565 B.n277 B.n121 163.367
R1566 B.n281 B.n121 163.367
R1567 B.n282 B.n281 163.367
R1568 B.n282 B.n117 163.367
R1569 B.n286 B.n117 163.367
R1570 B.n287 B.n286 163.367
R1571 B.n288 B.n287 163.367
R1572 B.n288 B.n115 163.367
R1573 B.n292 B.n115 163.367
R1574 B.n293 B.n292 163.367
R1575 B.n294 B.n293 163.367
R1576 B.n294 B.n113 163.367
R1577 B.n298 B.n113 163.367
R1578 B.n299 B.n298 163.367
R1579 B.n300 B.n299 163.367
R1580 B.n300 B.n111 163.367
R1581 B.n304 B.n111 163.367
R1582 B.n305 B.n304 163.367
R1583 B.n306 B.n305 163.367
R1584 B.n306 B.n109 163.367
R1585 B.n310 B.n109 163.367
R1586 B.n311 B.n310 163.367
R1587 B.n312 B.n311 163.367
R1588 B.n312 B.n107 163.367
R1589 B.n316 B.n107 163.367
R1590 B.n317 B.n316 163.367
R1591 B.n318 B.n317 163.367
R1592 B.n318 B.n105 163.367
R1593 B.n322 B.n105 163.367
R1594 B.n323 B.n322 163.367
R1595 B.n324 B.n323 163.367
R1596 B.n324 B.n103 163.367
R1597 B.n328 B.n103 163.367
R1598 B.n329 B.n328 163.367
R1599 B.n330 B.n329 163.367
R1600 B.n330 B.n101 163.367
R1601 B.n334 B.n101 163.367
R1602 B.n335 B.n334 163.367
R1603 B.n336 B.n335 163.367
R1604 B.n336 B.n99 163.367
R1605 B.n340 B.n99 163.367
R1606 B.n341 B.n340 163.367
R1607 B.n342 B.n341 163.367
R1608 B.n342 B.n97 163.367
R1609 B.n346 B.n97 163.367
R1610 B.n347 B.n346 163.367
R1611 B.n348 B.n347 163.367
R1612 B.n348 B.n95 163.367
R1613 B.n352 B.n95 163.367
R1614 B.n353 B.n352 163.367
R1615 B.n354 B.n353 163.367
R1616 B.n354 B.n93 163.367
R1617 B.n358 B.n93 163.367
R1618 B.n359 B.n358 163.367
R1619 B.n360 B.n359 163.367
R1620 B.n360 B.n91 163.367
R1621 B.n364 B.n91 163.367
R1622 B.n365 B.n364 163.367
R1623 B.n366 B.n89 163.367
R1624 B.n370 B.n89 163.367
R1625 B.n371 B.n370 163.367
R1626 B.n372 B.n371 163.367
R1627 B.n372 B.n87 163.367
R1628 B.n376 B.n87 163.367
R1629 B.n377 B.n376 163.367
R1630 B.n378 B.n377 163.367
R1631 B.n378 B.n85 163.367
R1632 B.n382 B.n85 163.367
R1633 B.n383 B.n382 163.367
R1634 B.n384 B.n383 163.367
R1635 B.n384 B.n83 163.367
R1636 B.n388 B.n83 163.367
R1637 B.n389 B.n388 163.367
R1638 B.n390 B.n389 163.367
R1639 B.n390 B.n81 163.367
R1640 B.n394 B.n81 163.367
R1641 B.n395 B.n394 163.367
R1642 B.n396 B.n395 163.367
R1643 B.n396 B.n79 163.367
R1644 B.n400 B.n79 163.367
R1645 B.n401 B.n400 163.367
R1646 B.n402 B.n401 163.367
R1647 B.n402 B.n77 163.367
R1648 B.n406 B.n77 163.367
R1649 B.n407 B.n406 163.367
R1650 B.n408 B.n407 163.367
R1651 B.n408 B.n75 163.367
R1652 B.n412 B.n75 163.367
R1653 B.n594 B.n593 163.367
R1654 B.n593 B.n592 163.367
R1655 B.n592 B.n11 163.367
R1656 B.n588 B.n11 163.367
R1657 B.n588 B.n587 163.367
R1658 B.n587 B.n586 163.367
R1659 B.n586 B.n13 163.367
R1660 B.n582 B.n13 163.367
R1661 B.n582 B.n581 163.367
R1662 B.n581 B.n580 163.367
R1663 B.n580 B.n15 163.367
R1664 B.n576 B.n15 163.367
R1665 B.n576 B.n575 163.367
R1666 B.n575 B.n574 163.367
R1667 B.n574 B.n17 163.367
R1668 B.n570 B.n17 163.367
R1669 B.n570 B.n569 163.367
R1670 B.n569 B.n568 163.367
R1671 B.n568 B.n19 163.367
R1672 B.n564 B.n19 163.367
R1673 B.n564 B.n563 163.367
R1674 B.n563 B.n562 163.367
R1675 B.n562 B.n21 163.367
R1676 B.n558 B.n21 163.367
R1677 B.n558 B.n557 163.367
R1678 B.n557 B.n556 163.367
R1679 B.n556 B.n23 163.367
R1680 B.n552 B.n23 163.367
R1681 B.n552 B.n551 163.367
R1682 B.n551 B.n550 163.367
R1683 B.n550 B.n25 163.367
R1684 B.n546 B.n25 163.367
R1685 B.n546 B.n545 163.367
R1686 B.n545 B.n544 163.367
R1687 B.n544 B.n27 163.367
R1688 B.n540 B.n27 163.367
R1689 B.n540 B.n539 163.367
R1690 B.n539 B.n538 163.367
R1691 B.n538 B.n29 163.367
R1692 B.n534 B.n29 163.367
R1693 B.n534 B.n533 163.367
R1694 B.n533 B.n532 163.367
R1695 B.n532 B.n31 163.367
R1696 B.n528 B.n31 163.367
R1697 B.n528 B.n527 163.367
R1698 B.n527 B.n526 163.367
R1699 B.n526 B.n33 163.367
R1700 B.n522 B.n33 163.367
R1701 B.n522 B.n521 163.367
R1702 B.n521 B.n520 163.367
R1703 B.n520 B.n35 163.367
R1704 B.n516 B.n35 163.367
R1705 B.n516 B.n515 163.367
R1706 B.n515 B.n514 163.367
R1707 B.n514 B.n37 163.367
R1708 B.n509 B.n37 163.367
R1709 B.n509 B.n508 163.367
R1710 B.n508 B.n507 163.367
R1711 B.n507 B.n41 163.367
R1712 B.n503 B.n41 163.367
R1713 B.n503 B.n502 163.367
R1714 B.n502 B.n501 163.367
R1715 B.n501 B.n43 163.367
R1716 B.n497 B.n43 163.367
R1717 B.n497 B.n496 163.367
R1718 B.n496 B.n47 163.367
R1719 B.n492 B.n47 163.367
R1720 B.n492 B.n491 163.367
R1721 B.n491 B.n490 163.367
R1722 B.n490 B.n49 163.367
R1723 B.n486 B.n49 163.367
R1724 B.n486 B.n485 163.367
R1725 B.n485 B.n484 163.367
R1726 B.n484 B.n51 163.367
R1727 B.n480 B.n51 163.367
R1728 B.n480 B.n479 163.367
R1729 B.n479 B.n478 163.367
R1730 B.n478 B.n53 163.367
R1731 B.n474 B.n53 163.367
R1732 B.n474 B.n473 163.367
R1733 B.n473 B.n472 163.367
R1734 B.n472 B.n55 163.367
R1735 B.n468 B.n55 163.367
R1736 B.n468 B.n467 163.367
R1737 B.n467 B.n466 163.367
R1738 B.n466 B.n57 163.367
R1739 B.n462 B.n57 163.367
R1740 B.n462 B.n461 163.367
R1741 B.n461 B.n460 163.367
R1742 B.n460 B.n59 163.367
R1743 B.n456 B.n59 163.367
R1744 B.n456 B.n455 163.367
R1745 B.n455 B.n454 163.367
R1746 B.n454 B.n61 163.367
R1747 B.n450 B.n61 163.367
R1748 B.n450 B.n449 163.367
R1749 B.n449 B.n448 163.367
R1750 B.n448 B.n63 163.367
R1751 B.n444 B.n63 163.367
R1752 B.n444 B.n443 163.367
R1753 B.n443 B.n442 163.367
R1754 B.n442 B.n65 163.367
R1755 B.n438 B.n65 163.367
R1756 B.n438 B.n437 163.367
R1757 B.n437 B.n436 163.367
R1758 B.n436 B.n67 163.367
R1759 B.n432 B.n67 163.367
R1760 B.n432 B.n431 163.367
R1761 B.n431 B.n430 163.367
R1762 B.n430 B.n69 163.367
R1763 B.n426 B.n69 163.367
R1764 B.n426 B.n425 163.367
R1765 B.n425 B.n424 163.367
R1766 B.n424 B.n71 163.367
R1767 B.n420 B.n71 163.367
R1768 B.n420 B.n419 163.367
R1769 B.n419 B.n418 163.367
R1770 B.n418 B.n73 163.367
R1771 B.n414 B.n73 163.367
R1772 B.n414 B.n413 163.367
R1773 B.n120 B.n119 59.5399
R1774 B.n267 B.n127 59.5399
R1775 B.n511 B.n39 59.5399
R1776 B.n46 B.n45 59.5399
R1777 B.n596 B.n595 34.1859
R1778 B.n411 B.n74 34.1859
R1779 B.n367 B.n90 34.1859
R1780 B.n183 B.n182 34.1859
R1781 B B.n619 18.0485
R1782 B.n119 B.n118 14.9338
R1783 B.n127 B.n126 14.9338
R1784 B.n39 B.n38 14.9338
R1785 B.n45 B.n44 14.9338
R1786 B.n595 B.n10 10.6151
R1787 B.n591 B.n10 10.6151
R1788 B.n591 B.n590 10.6151
R1789 B.n590 B.n589 10.6151
R1790 B.n589 B.n12 10.6151
R1791 B.n585 B.n12 10.6151
R1792 B.n585 B.n584 10.6151
R1793 B.n584 B.n583 10.6151
R1794 B.n583 B.n14 10.6151
R1795 B.n579 B.n14 10.6151
R1796 B.n579 B.n578 10.6151
R1797 B.n578 B.n577 10.6151
R1798 B.n577 B.n16 10.6151
R1799 B.n573 B.n16 10.6151
R1800 B.n573 B.n572 10.6151
R1801 B.n572 B.n571 10.6151
R1802 B.n571 B.n18 10.6151
R1803 B.n567 B.n18 10.6151
R1804 B.n567 B.n566 10.6151
R1805 B.n566 B.n565 10.6151
R1806 B.n565 B.n20 10.6151
R1807 B.n561 B.n20 10.6151
R1808 B.n561 B.n560 10.6151
R1809 B.n560 B.n559 10.6151
R1810 B.n559 B.n22 10.6151
R1811 B.n555 B.n22 10.6151
R1812 B.n555 B.n554 10.6151
R1813 B.n554 B.n553 10.6151
R1814 B.n553 B.n24 10.6151
R1815 B.n549 B.n24 10.6151
R1816 B.n549 B.n548 10.6151
R1817 B.n548 B.n547 10.6151
R1818 B.n547 B.n26 10.6151
R1819 B.n543 B.n26 10.6151
R1820 B.n543 B.n542 10.6151
R1821 B.n542 B.n541 10.6151
R1822 B.n541 B.n28 10.6151
R1823 B.n537 B.n28 10.6151
R1824 B.n537 B.n536 10.6151
R1825 B.n536 B.n535 10.6151
R1826 B.n535 B.n30 10.6151
R1827 B.n531 B.n30 10.6151
R1828 B.n531 B.n530 10.6151
R1829 B.n530 B.n529 10.6151
R1830 B.n529 B.n32 10.6151
R1831 B.n525 B.n32 10.6151
R1832 B.n525 B.n524 10.6151
R1833 B.n524 B.n523 10.6151
R1834 B.n523 B.n34 10.6151
R1835 B.n519 B.n34 10.6151
R1836 B.n519 B.n518 10.6151
R1837 B.n518 B.n517 10.6151
R1838 B.n517 B.n36 10.6151
R1839 B.n513 B.n36 10.6151
R1840 B.n513 B.n512 10.6151
R1841 B.n510 B.n40 10.6151
R1842 B.n506 B.n40 10.6151
R1843 B.n506 B.n505 10.6151
R1844 B.n505 B.n504 10.6151
R1845 B.n504 B.n42 10.6151
R1846 B.n500 B.n42 10.6151
R1847 B.n500 B.n499 10.6151
R1848 B.n499 B.n498 10.6151
R1849 B.n495 B.n494 10.6151
R1850 B.n494 B.n493 10.6151
R1851 B.n493 B.n48 10.6151
R1852 B.n489 B.n48 10.6151
R1853 B.n489 B.n488 10.6151
R1854 B.n488 B.n487 10.6151
R1855 B.n487 B.n50 10.6151
R1856 B.n483 B.n50 10.6151
R1857 B.n483 B.n482 10.6151
R1858 B.n482 B.n481 10.6151
R1859 B.n481 B.n52 10.6151
R1860 B.n477 B.n52 10.6151
R1861 B.n477 B.n476 10.6151
R1862 B.n476 B.n475 10.6151
R1863 B.n475 B.n54 10.6151
R1864 B.n471 B.n54 10.6151
R1865 B.n471 B.n470 10.6151
R1866 B.n470 B.n469 10.6151
R1867 B.n469 B.n56 10.6151
R1868 B.n465 B.n56 10.6151
R1869 B.n465 B.n464 10.6151
R1870 B.n464 B.n463 10.6151
R1871 B.n463 B.n58 10.6151
R1872 B.n459 B.n58 10.6151
R1873 B.n459 B.n458 10.6151
R1874 B.n458 B.n457 10.6151
R1875 B.n457 B.n60 10.6151
R1876 B.n453 B.n60 10.6151
R1877 B.n453 B.n452 10.6151
R1878 B.n452 B.n451 10.6151
R1879 B.n451 B.n62 10.6151
R1880 B.n447 B.n62 10.6151
R1881 B.n447 B.n446 10.6151
R1882 B.n446 B.n445 10.6151
R1883 B.n445 B.n64 10.6151
R1884 B.n441 B.n64 10.6151
R1885 B.n441 B.n440 10.6151
R1886 B.n440 B.n439 10.6151
R1887 B.n439 B.n66 10.6151
R1888 B.n435 B.n66 10.6151
R1889 B.n435 B.n434 10.6151
R1890 B.n434 B.n433 10.6151
R1891 B.n433 B.n68 10.6151
R1892 B.n429 B.n68 10.6151
R1893 B.n429 B.n428 10.6151
R1894 B.n428 B.n427 10.6151
R1895 B.n427 B.n70 10.6151
R1896 B.n423 B.n70 10.6151
R1897 B.n423 B.n422 10.6151
R1898 B.n422 B.n421 10.6151
R1899 B.n421 B.n72 10.6151
R1900 B.n417 B.n72 10.6151
R1901 B.n417 B.n416 10.6151
R1902 B.n416 B.n415 10.6151
R1903 B.n415 B.n74 10.6151
R1904 B.n368 B.n367 10.6151
R1905 B.n369 B.n368 10.6151
R1906 B.n369 B.n88 10.6151
R1907 B.n373 B.n88 10.6151
R1908 B.n374 B.n373 10.6151
R1909 B.n375 B.n374 10.6151
R1910 B.n375 B.n86 10.6151
R1911 B.n379 B.n86 10.6151
R1912 B.n380 B.n379 10.6151
R1913 B.n381 B.n380 10.6151
R1914 B.n381 B.n84 10.6151
R1915 B.n385 B.n84 10.6151
R1916 B.n386 B.n385 10.6151
R1917 B.n387 B.n386 10.6151
R1918 B.n387 B.n82 10.6151
R1919 B.n391 B.n82 10.6151
R1920 B.n392 B.n391 10.6151
R1921 B.n393 B.n392 10.6151
R1922 B.n393 B.n80 10.6151
R1923 B.n397 B.n80 10.6151
R1924 B.n398 B.n397 10.6151
R1925 B.n399 B.n398 10.6151
R1926 B.n399 B.n78 10.6151
R1927 B.n403 B.n78 10.6151
R1928 B.n404 B.n403 10.6151
R1929 B.n405 B.n404 10.6151
R1930 B.n405 B.n76 10.6151
R1931 B.n409 B.n76 10.6151
R1932 B.n410 B.n409 10.6151
R1933 B.n411 B.n410 10.6151
R1934 B.n183 B.n154 10.6151
R1935 B.n187 B.n154 10.6151
R1936 B.n188 B.n187 10.6151
R1937 B.n189 B.n188 10.6151
R1938 B.n189 B.n152 10.6151
R1939 B.n193 B.n152 10.6151
R1940 B.n194 B.n193 10.6151
R1941 B.n195 B.n194 10.6151
R1942 B.n195 B.n150 10.6151
R1943 B.n199 B.n150 10.6151
R1944 B.n200 B.n199 10.6151
R1945 B.n201 B.n200 10.6151
R1946 B.n201 B.n148 10.6151
R1947 B.n205 B.n148 10.6151
R1948 B.n206 B.n205 10.6151
R1949 B.n207 B.n206 10.6151
R1950 B.n207 B.n146 10.6151
R1951 B.n211 B.n146 10.6151
R1952 B.n212 B.n211 10.6151
R1953 B.n213 B.n212 10.6151
R1954 B.n213 B.n144 10.6151
R1955 B.n217 B.n144 10.6151
R1956 B.n218 B.n217 10.6151
R1957 B.n219 B.n218 10.6151
R1958 B.n219 B.n142 10.6151
R1959 B.n223 B.n142 10.6151
R1960 B.n224 B.n223 10.6151
R1961 B.n225 B.n224 10.6151
R1962 B.n225 B.n140 10.6151
R1963 B.n229 B.n140 10.6151
R1964 B.n230 B.n229 10.6151
R1965 B.n231 B.n230 10.6151
R1966 B.n231 B.n138 10.6151
R1967 B.n235 B.n138 10.6151
R1968 B.n236 B.n235 10.6151
R1969 B.n237 B.n236 10.6151
R1970 B.n237 B.n136 10.6151
R1971 B.n241 B.n136 10.6151
R1972 B.n242 B.n241 10.6151
R1973 B.n243 B.n242 10.6151
R1974 B.n243 B.n134 10.6151
R1975 B.n247 B.n134 10.6151
R1976 B.n248 B.n247 10.6151
R1977 B.n249 B.n248 10.6151
R1978 B.n249 B.n132 10.6151
R1979 B.n253 B.n132 10.6151
R1980 B.n254 B.n253 10.6151
R1981 B.n255 B.n254 10.6151
R1982 B.n255 B.n130 10.6151
R1983 B.n259 B.n130 10.6151
R1984 B.n260 B.n259 10.6151
R1985 B.n261 B.n260 10.6151
R1986 B.n261 B.n128 10.6151
R1987 B.n265 B.n128 10.6151
R1988 B.n266 B.n265 10.6151
R1989 B.n268 B.n124 10.6151
R1990 B.n272 B.n124 10.6151
R1991 B.n273 B.n272 10.6151
R1992 B.n274 B.n273 10.6151
R1993 B.n274 B.n122 10.6151
R1994 B.n278 B.n122 10.6151
R1995 B.n279 B.n278 10.6151
R1996 B.n280 B.n279 10.6151
R1997 B.n284 B.n283 10.6151
R1998 B.n285 B.n284 10.6151
R1999 B.n285 B.n116 10.6151
R2000 B.n289 B.n116 10.6151
R2001 B.n290 B.n289 10.6151
R2002 B.n291 B.n290 10.6151
R2003 B.n291 B.n114 10.6151
R2004 B.n295 B.n114 10.6151
R2005 B.n296 B.n295 10.6151
R2006 B.n297 B.n296 10.6151
R2007 B.n297 B.n112 10.6151
R2008 B.n301 B.n112 10.6151
R2009 B.n302 B.n301 10.6151
R2010 B.n303 B.n302 10.6151
R2011 B.n303 B.n110 10.6151
R2012 B.n307 B.n110 10.6151
R2013 B.n308 B.n307 10.6151
R2014 B.n309 B.n308 10.6151
R2015 B.n309 B.n108 10.6151
R2016 B.n313 B.n108 10.6151
R2017 B.n314 B.n313 10.6151
R2018 B.n315 B.n314 10.6151
R2019 B.n315 B.n106 10.6151
R2020 B.n319 B.n106 10.6151
R2021 B.n320 B.n319 10.6151
R2022 B.n321 B.n320 10.6151
R2023 B.n321 B.n104 10.6151
R2024 B.n325 B.n104 10.6151
R2025 B.n326 B.n325 10.6151
R2026 B.n327 B.n326 10.6151
R2027 B.n327 B.n102 10.6151
R2028 B.n331 B.n102 10.6151
R2029 B.n332 B.n331 10.6151
R2030 B.n333 B.n332 10.6151
R2031 B.n333 B.n100 10.6151
R2032 B.n337 B.n100 10.6151
R2033 B.n338 B.n337 10.6151
R2034 B.n339 B.n338 10.6151
R2035 B.n339 B.n98 10.6151
R2036 B.n343 B.n98 10.6151
R2037 B.n344 B.n343 10.6151
R2038 B.n345 B.n344 10.6151
R2039 B.n345 B.n96 10.6151
R2040 B.n349 B.n96 10.6151
R2041 B.n350 B.n349 10.6151
R2042 B.n351 B.n350 10.6151
R2043 B.n351 B.n94 10.6151
R2044 B.n355 B.n94 10.6151
R2045 B.n356 B.n355 10.6151
R2046 B.n357 B.n356 10.6151
R2047 B.n357 B.n92 10.6151
R2048 B.n361 B.n92 10.6151
R2049 B.n362 B.n361 10.6151
R2050 B.n363 B.n362 10.6151
R2051 B.n363 B.n90 10.6151
R2052 B.n182 B.n181 10.6151
R2053 B.n181 B.n156 10.6151
R2054 B.n177 B.n156 10.6151
R2055 B.n177 B.n176 10.6151
R2056 B.n176 B.n175 10.6151
R2057 B.n175 B.n158 10.6151
R2058 B.n171 B.n158 10.6151
R2059 B.n171 B.n170 10.6151
R2060 B.n170 B.n169 10.6151
R2061 B.n169 B.n160 10.6151
R2062 B.n165 B.n160 10.6151
R2063 B.n165 B.n164 10.6151
R2064 B.n164 B.n163 10.6151
R2065 B.n163 B.n0 10.6151
R2066 B.n615 B.n1 10.6151
R2067 B.n615 B.n614 10.6151
R2068 B.n614 B.n613 10.6151
R2069 B.n613 B.n4 10.6151
R2070 B.n609 B.n4 10.6151
R2071 B.n609 B.n608 10.6151
R2072 B.n608 B.n607 10.6151
R2073 B.n607 B.n6 10.6151
R2074 B.n603 B.n6 10.6151
R2075 B.n603 B.n602 10.6151
R2076 B.n602 B.n601 10.6151
R2077 B.n601 B.n8 10.6151
R2078 B.n597 B.n8 10.6151
R2079 B.n597 B.n596 10.6151
R2080 B.n511 B.n510 6.5566
R2081 B.n498 B.n46 6.5566
R2082 B.n268 B.n267 6.5566
R2083 B.n280 B.n120 6.5566
R2084 B.n512 B.n511 4.05904
R2085 B.n495 B.n46 4.05904
R2086 B.n267 B.n266 4.05904
R2087 B.n283 B.n120 4.05904
R2088 B.n619 B.n0 2.81026
R2089 B.n619 B.n1 2.81026
R2090 VN.n0 VN.t0 1034.82
R2091 VN.n1 VN.t1 1034.82
R2092 VN.n0 VN.t2 1034.8
R2093 VN.n1 VN.t3 1034.8
R2094 VN VN.n1 113.906
R2095 VN VN.n0 70.265
R2096 VDD2.n2 VDD2.n0 111.201
R2097 VDD2.n2 VDD2.n1 70.9434
R2098 VDD2.n1 VDD2.t0 1.92615
R2099 VDD2.n1 VDD2.t2 1.92615
R2100 VDD2.n0 VDD2.t3 1.92615
R2101 VDD2.n0 VDD2.t1 1.92615
R2102 VDD2 VDD2.n2 0.0586897
C0 VP VN 5.53832f
C1 w_n1432_n4344# VN 2.11926f
C2 B VTAIL 4.8762f
C3 VDD1 VTAIL 10.859401f
C4 VN VDD2 3.43708f
C5 VP VTAIL 2.77546f
C6 w_n1432_n4344# VTAIL 5.497169f
C7 B VDD1 1.0111f
C8 B VP 1.04096f
C9 B w_n1432_n4344# 7.95628f
C10 VP VDD1 3.5467f
C11 w_n1432_n4344# VDD1 1.13677f
C12 VDD2 VTAIL 10.8991f
C13 VP w_n1432_n4344# 2.29789f
C14 B VDD2 1.02899f
C15 VDD1 VDD2 0.510386f
C16 VP VDD2 0.257297f
C17 w_n1432_n4344# VDD2 1.14626f
C18 VN VTAIL 2.76136f
C19 B VN 0.754595f
C20 VN VDD1 0.147484f
C21 VDD2 VSUBS 0.764689f
C22 VDD1 VSUBS 5.958925f
C23 VTAIL VSUBS 0.976607f
C24 VN VSUBS 6.78896f
C25 VP VSUBS 1.341558f
C26 B VSUBS 2.809631f
C27 w_n1432_n4344# VSUBS 76.142296f
C28 VDD2.t3 VSUBS 0.408962f
C29 VDD2.t1 VSUBS 0.408962f
C30 VDD2.n0 VSUBS 4.26809f
C31 VDD2.t0 VSUBS 0.408962f
C32 VDD2.t2 VSUBS 0.408962f
C33 VDD2.n1 VSUBS 3.37782f
C34 VDD2.n2 VSUBS 4.94606f
C35 VN.t0 VSUBS 1.40863f
C36 VN.t2 VSUBS 1.40862f
C37 VN.n0 VSUBS 1.05372f
C38 VN.t1 VSUBS 1.40863f
C39 VN.t3 VSUBS 1.40862f
C40 VN.n1 VSUBS 2.20373f
C41 B.n0 VSUBS 0.005182f
C42 B.n1 VSUBS 0.005182f
C43 B.n2 VSUBS 0.008194f
C44 B.n3 VSUBS 0.008194f
C45 B.n4 VSUBS 0.008194f
C46 B.n5 VSUBS 0.008194f
C47 B.n6 VSUBS 0.008194f
C48 B.n7 VSUBS 0.008194f
C49 B.n8 VSUBS 0.008194f
C50 B.n9 VSUBS 0.019594f
C51 B.n10 VSUBS 0.008194f
C52 B.n11 VSUBS 0.008194f
C53 B.n12 VSUBS 0.008194f
C54 B.n13 VSUBS 0.008194f
C55 B.n14 VSUBS 0.008194f
C56 B.n15 VSUBS 0.008194f
C57 B.n16 VSUBS 0.008194f
C58 B.n17 VSUBS 0.008194f
C59 B.n18 VSUBS 0.008194f
C60 B.n19 VSUBS 0.008194f
C61 B.n20 VSUBS 0.008194f
C62 B.n21 VSUBS 0.008194f
C63 B.n22 VSUBS 0.008194f
C64 B.n23 VSUBS 0.008194f
C65 B.n24 VSUBS 0.008194f
C66 B.n25 VSUBS 0.008194f
C67 B.n26 VSUBS 0.008194f
C68 B.n27 VSUBS 0.008194f
C69 B.n28 VSUBS 0.008194f
C70 B.n29 VSUBS 0.008194f
C71 B.n30 VSUBS 0.008194f
C72 B.n31 VSUBS 0.008194f
C73 B.n32 VSUBS 0.008194f
C74 B.n33 VSUBS 0.008194f
C75 B.n34 VSUBS 0.008194f
C76 B.n35 VSUBS 0.008194f
C77 B.n36 VSUBS 0.008194f
C78 B.n37 VSUBS 0.008194f
C79 B.t2 VSUBS 0.379521f
C80 B.t1 VSUBS 0.390341f
C81 B.t0 VSUBS 0.343036f
C82 B.n38 VSUBS 0.443313f
C83 B.n39 VSUBS 0.358389f
C84 B.n40 VSUBS 0.008194f
C85 B.n41 VSUBS 0.008194f
C86 B.n42 VSUBS 0.008194f
C87 B.n43 VSUBS 0.008194f
C88 B.t8 VSUBS 0.379525f
C89 B.t7 VSUBS 0.390345f
C90 B.t6 VSUBS 0.343036f
C91 B.n44 VSUBS 0.443309f
C92 B.n45 VSUBS 0.358385f
C93 B.n46 VSUBS 0.018986f
C94 B.n47 VSUBS 0.008194f
C95 B.n48 VSUBS 0.008194f
C96 B.n49 VSUBS 0.008194f
C97 B.n50 VSUBS 0.008194f
C98 B.n51 VSUBS 0.008194f
C99 B.n52 VSUBS 0.008194f
C100 B.n53 VSUBS 0.008194f
C101 B.n54 VSUBS 0.008194f
C102 B.n55 VSUBS 0.008194f
C103 B.n56 VSUBS 0.008194f
C104 B.n57 VSUBS 0.008194f
C105 B.n58 VSUBS 0.008194f
C106 B.n59 VSUBS 0.008194f
C107 B.n60 VSUBS 0.008194f
C108 B.n61 VSUBS 0.008194f
C109 B.n62 VSUBS 0.008194f
C110 B.n63 VSUBS 0.008194f
C111 B.n64 VSUBS 0.008194f
C112 B.n65 VSUBS 0.008194f
C113 B.n66 VSUBS 0.008194f
C114 B.n67 VSUBS 0.008194f
C115 B.n68 VSUBS 0.008194f
C116 B.n69 VSUBS 0.008194f
C117 B.n70 VSUBS 0.008194f
C118 B.n71 VSUBS 0.008194f
C119 B.n72 VSUBS 0.008194f
C120 B.n73 VSUBS 0.008194f
C121 B.n74 VSUBS 0.019007f
C122 B.n75 VSUBS 0.008194f
C123 B.n76 VSUBS 0.008194f
C124 B.n77 VSUBS 0.008194f
C125 B.n78 VSUBS 0.008194f
C126 B.n79 VSUBS 0.008194f
C127 B.n80 VSUBS 0.008194f
C128 B.n81 VSUBS 0.008194f
C129 B.n82 VSUBS 0.008194f
C130 B.n83 VSUBS 0.008194f
C131 B.n84 VSUBS 0.008194f
C132 B.n85 VSUBS 0.008194f
C133 B.n86 VSUBS 0.008194f
C134 B.n87 VSUBS 0.008194f
C135 B.n88 VSUBS 0.008194f
C136 B.n89 VSUBS 0.008194f
C137 B.n90 VSUBS 0.019932f
C138 B.n91 VSUBS 0.008194f
C139 B.n92 VSUBS 0.008194f
C140 B.n93 VSUBS 0.008194f
C141 B.n94 VSUBS 0.008194f
C142 B.n95 VSUBS 0.008194f
C143 B.n96 VSUBS 0.008194f
C144 B.n97 VSUBS 0.008194f
C145 B.n98 VSUBS 0.008194f
C146 B.n99 VSUBS 0.008194f
C147 B.n100 VSUBS 0.008194f
C148 B.n101 VSUBS 0.008194f
C149 B.n102 VSUBS 0.008194f
C150 B.n103 VSUBS 0.008194f
C151 B.n104 VSUBS 0.008194f
C152 B.n105 VSUBS 0.008194f
C153 B.n106 VSUBS 0.008194f
C154 B.n107 VSUBS 0.008194f
C155 B.n108 VSUBS 0.008194f
C156 B.n109 VSUBS 0.008194f
C157 B.n110 VSUBS 0.008194f
C158 B.n111 VSUBS 0.008194f
C159 B.n112 VSUBS 0.008194f
C160 B.n113 VSUBS 0.008194f
C161 B.n114 VSUBS 0.008194f
C162 B.n115 VSUBS 0.008194f
C163 B.n116 VSUBS 0.008194f
C164 B.n117 VSUBS 0.008194f
C165 B.t10 VSUBS 0.379525f
C166 B.t11 VSUBS 0.390345f
C167 B.t9 VSUBS 0.343036f
C168 B.n118 VSUBS 0.443309f
C169 B.n119 VSUBS 0.358385f
C170 B.n120 VSUBS 0.018986f
C171 B.n121 VSUBS 0.008194f
C172 B.n122 VSUBS 0.008194f
C173 B.n123 VSUBS 0.008194f
C174 B.n124 VSUBS 0.008194f
C175 B.n125 VSUBS 0.008194f
C176 B.t4 VSUBS 0.379521f
C177 B.t5 VSUBS 0.390341f
C178 B.t3 VSUBS 0.343036f
C179 B.n126 VSUBS 0.443313f
C180 B.n127 VSUBS 0.358389f
C181 B.n128 VSUBS 0.008194f
C182 B.n129 VSUBS 0.008194f
C183 B.n130 VSUBS 0.008194f
C184 B.n131 VSUBS 0.008194f
C185 B.n132 VSUBS 0.008194f
C186 B.n133 VSUBS 0.008194f
C187 B.n134 VSUBS 0.008194f
C188 B.n135 VSUBS 0.008194f
C189 B.n136 VSUBS 0.008194f
C190 B.n137 VSUBS 0.008194f
C191 B.n138 VSUBS 0.008194f
C192 B.n139 VSUBS 0.008194f
C193 B.n140 VSUBS 0.008194f
C194 B.n141 VSUBS 0.008194f
C195 B.n142 VSUBS 0.008194f
C196 B.n143 VSUBS 0.008194f
C197 B.n144 VSUBS 0.008194f
C198 B.n145 VSUBS 0.008194f
C199 B.n146 VSUBS 0.008194f
C200 B.n147 VSUBS 0.008194f
C201 B.n148 VSUBS 0.008194f
C202 B.n149 VSUBS 0.008194f
C203 B.n150 VSUBS 0.008194f
C204 B.n151 VSUBS 0.008194f
C205 B.n152 VSUBS 0.008194f
C206 B.n153 VSUBS 0.008194f
C207 B.n154 VSUBS 0.008194f
C208 B.n155 VSUBS 0.019594f
C209 B.n156 VSUBS 0.008194f
C210 B.n157 VSUBS 0.008194f
C211 B.n158 VSUBS 0.008194f
C212 B.n159 VSUBS 0.008194f
C213 B.n160 VSUBS 0.008194f
C214 B.n161 VSUBS 0.008194f
C215 B.n162 VSUBS 0.008194f
C216 B.n163 VSUBS 0.008194f
C217 B.n164 VSUBS 0.008194f
C218 B.n165 VSUBS 0.008194f
C219 B.n166 VSUBS 0.008194f
C220 B.n167 VSUBS 0.008194f
C221 B.n168 VSUBS 0.008194f
C222 B.n169 VSUBS 0.008194f
C223 B.n170 VSUBS 0.008194f
C224 B.n171 VSUBS 0.008194f
C225 B.n172 VSUBS 0.008194f
C226 B.n173 VSUBS 0.008194f
C227 B.n174 VSUBS 0.008194f
C228 B.n175 VSUBS 0.008194f
C229 B.n176 VSUBS 0.008194f
C230 B.n177 VSUBS 0.008194f
C231 B.n178 VSUBS 0.008194f
C232 B.n179 VSUBS 0.008194f
C233 B.n180 VSUBS 0.008194f
C234 B.n181 VSUBS 0.008194f
C235 B.n182 VSUBS 0.019594f
C236 B.n183 VSUBS 0.019932f
C237 B.n184 VSUBS 0.019932f
C238 B.n185 VSUBS 0.008194f
C239 B.n186 VSUBS 0.008194f
C240 B.n187 VSUBS 0.008194f
C241 B.n188 VSUBS 0.008194f
C242 B.n189 VSUBS 0.008194f
C243 B.n190 VSUBS 0.008194f
C244 B.n191 VSUBS 0.008194f
C245 B.n192 VSUBS 0.008194f
C246 B.n193 VSUBS 0.008194f
C247 B.n194 VSUBS 0.008194f
C248 B.n195 VSUBS 0.008194f
C249 B.n196 VSUBS 0.008194f
C250 B.n197 VSUBS 0.008194f
C251 B.n198 VSUBS 0.008194f
C252 B.n199 VSUBS 0.008194f
C253 B.n200 VSUBS 0.008194f
C254 B.n201 VSUBS 0.008194f
C255 B.n202 VSUBS 0.008194f
C256 B.n203 VSUBS 0.008194f
C257 B.n204 VSUBS 0.008194f
C258 B.n205 VSUBS 0.008194f
C259 B.n206 VSUBS 0.008194f
C260 B.n207 VSUBS 0.008194f
C261 B.n208 VSUBS 0.008194f
C262 B.n209 VSUBS 0.008194f
C263 B.n210 VSUBS 0.008194f
C264 B.n211 VSUBS 0.008194f
C265 B.n212 VSUBS 0.008194f
C266 B.n213 VSUBS 0.008194f
C267 B.n214 VSUBS 0.008194f
C268 B.n215 VSUBS 0.008194f
C269 B.n216 VSUBS 0.008194f
C270 B.n217 VSUBS 0.008194f
C271 B.n218 VSUBS 0.008194f
C272 B.n219 VSUBS 0.008194f
C273 B.n220 VSUBS 0.008194f
C274 B.n221 VSUBS 0.008194f
C275 B.n222 VSUBS 0.008194f
C276 B.n223 VSUBS 0.008194f
C277 B.n224 VSUBS 0.008194f
C278 B.n225 VSUBS 0.008194f
C279 B.n226 VSUBS 0.008194f
C280 B.n227 VSUBS 0.008194f
C281 B.n228 VSUBS 0.008194f
C282 B.n229 VSUBS 0.008194f
C283 B.n230 VSUBS 0.008194f
C284 B.n231 VSUBS 0.008194f
C285 B.n232 VSUBS 0.008194f
C286 B.n233 VSUBS 0.008194f
C287 B.n234 VSUBS 0.008194f
C288 B.n235 VSUBS 0.008194f
C289 B.n236 VSUBS 0.008194f
C290 B.n237 VSUBS 0.008194f
C291 B.n238 VSUBS 0.008194f
C292 B.n239 VSUBS 0.008194f
C293 B.n240 VSUBS 0.008194f
C294 B.n241 VSUBS 0.008194f
C295 B.n242 VSUBS 0.008194f
C296 B.n243 VSUBS 0.008194f
C297 B.n244 VSUBS 0.008194f
C298 B.n245 VSUBS 0.008194f
C299 B.n246 VSUBS 0.008194f
C300 B.n247 VSUBS 0.008194f
C301 B.n248 VSUBS 0.008194f
C302 B.n249 VSUBS 0.008194f
C303 B.n250 VSUBS 0.008194f
C304 B.n251 VSUBS 0.008194f
C305 B.n252 VSUBS 0.008194f
C306 B.n253 VSUBS 0.008194f
C307 B.n254 VSUBS 0.008194f
C308 B.n255 VSUBS 0.008194f
C309 B.n256 VSUBS 0.008194f
C310 B.n257 VSUBS 0.008194f
C311 B.n258 VSUBS 0.008194f
C312 B.n259 VSUBS 0.008194f
C313 B.n260 VSUBS 0.008194f
C314 B.n261 VSUBS 0.008194f
C315 B.n262 VSUBS 0.008194f
C316 B.n263 VSUBS 0.008194f
C317 B.n264 VSUBS 0.008194f
C318 B.n265 VSUBS 0.008194f
C319 B.n266 VSUBS 0.005664f
C320 B.n267 VSUBS 0.018986f
C321 B.n268 VSUBS 0.006628f
C322 B.n269 VSUBS 0.008194f
C323 B.n270 VSUBS 0.008194f
C324 B.n271 VSUBS 0.008194f
C325 B.n272 VSUBS 0.008194f
C326 B.n273 VSUBS 0.008194f
C327 B.n274 VSUBS 0.008194f
C328 B.n275 VSUBS 0.008194f
C329 B.n276 VSUBS 0.008194f
C330 B.n277 VSUBS 0.008194f
C331 B.n278 VSUBS 0.008194f
C332 B.n279 VSUBS 0.008194f
C333 B.n280 VSUBS 0.006628f
C334 B.n281 VSUBS 0.008194f
C335 B.n282 VSUBS 0.008194f
C336 B.n283 VSUBS 0.005664f
C337 B.n284 VSUBS 0.008194f
C338 B.n285 VSUBS 0.008194f
C339 B.n286 VSUBS 0.008194f
C340 B.n287 VSUBS 0.008194f
C341 B.n288 VSUBS 0.008194f
C342 B.n289 VSUBS 0.008194f
C343 B.n290 VSUBS 0.008194f
C344 B.n291 VSUBS 0.008194f
C345 B.n292 VSUBS 0.008194f
C346 B.n293 VSUBS 0.008194f
C347 B.n294 VSUBS 0.008194f
C348 B.n295 VSUBS 0.008194f
C349 B.n296 VSUBS 0.008194f
C350 B.n297 VSUBS 0.008194f
C351 B.n298 VSUBS 0.008194f
C352 B.n299 VSUBS 0.008194f
C353 B.n300 VSUBS 0.008194f
C354 B.n301 VSUBS 0.008194f
C355 B.n302 VSUBS 0.008194f
C356 B.n303 VSUBS 0.008194f
C357 B.n304 VSUBS 0.008194f
C358 B.n305 VSUBS 0.008194f
C359 B.n306 VSUBS 0.008194f
C360 B.n307 VSUBS 0.008194f
C361 B.n308 VSUBS 0.008194f
C362 B.n309 VSUBS 0.008194f
C363 B.n310 VSUBS 0.008194f
C364 B.n311 VSUBS 0.008194f
C365 B.n312 VSUBS 0.008194f
C366 B.n313 VSUBS 0.008194f
C367 B.n314 VSUBS 0.008194f
C368 B.n315 VSUBS 0.008194f
C369 B.n316 VSUBS 0.008194f
C370 B.n317 VSUBS 0.008194f
C371 B.n318 VSUBS 0.008194f
C372 B.n319 VSUBS 0.008194f
C373 B.n320 VSUBS 0.008194f
C374 B.n321 VSUBS 0.008194f
C375 B.n322 VSUBS 0.008194f
C376 B.n323 VSUBS 0.008194f
C377 B.n324 VSUBS 0.008194f
C378 B.n325 VSUBS 0.008194f
C379 B.n326 VSUBS 0.008194f
C380 B.n327 VSUBS 0.008194f
C381 B.n328 VSUBS 0.008194f
C382 B.n329 VSUBS 0.008194f
C383 B.n330 VSUBS 0.008194f
C384 B.n331 VSUBS 0.008194f
C385 B.n332 VSUBS 0.008194f
C386 B.n333 VSUBS 0.008194f
C387 B.n334 VSUBS 0.008194f
C388 B.n335 VSUBS 0.008194f
C389 B.n336 VSUBS 0.008194f
C390 B.n337 VSUBS 0.008194f
C391 B.n338 VSUBS 0.008194f
C392 B.n339 VSUBS 0.008194f
C393 B.n340 VSUBS 0.008194f
C394 B.n341 VSUBS 0.008194f
C395 B.n342 VSUBS 0.008194f
C396 B.n343 VSUBS 0.008194f
C397 B.n344 VSUBS 0.008194f
C398 B.n345 VSUBS 0.008194f
C399 B.n346 VSUBS 0.008194f
C400 B.n347 VSUBS 0.008194f
C401 B.n348 VSUBS 0.008194f
C402 B.n349 VSUBS 0.008194f
C403 B.n350 VSUBS 0.008194f
C404 B.n351 VSUBS 0.008194f
C405 B.n352 VSUBS 0.008194f
C406 B.n353 VSUBS 0.008194f
C407 B.n354 VSUBS 0.008194f
C408 B.n355 VSUBS 0.008194f
C409 B.n356 VSUBS 0.008194f
C410 B.n357 VSUBS 0.008194f
C411 B.n358 VSUBS 0.008194f
C412 B.n359 VSUBS 0.008194f
C413 B.n360 VSUBS 0.008194f
C414 B.n361 VSUBS 0.008194f
C415 B.n362 VSUBS 0.008194f
C416 B.n363 VSUBS 0.008194f
C417 B.n364 VSUBS 0.008194f
C418 B.n365 VSUBS 0.019932f
C419 B.n366 VSUBS 0.019594f
C420 B.n367 VSUBS 0.019594f
C421 B.n368 VSUBS 0.008194f
C422 B.n369 VSUBS 0.008194f
C423 B.n370 VSUBS 0.008194f
C424 B.n371 VSUBS 0.008194f
C425 B.n372 VSUBS 0.008194f
C426 B.n373 VSUBS 0.008194f
C427 B.n374 VSUBS 0.008194f
C428 B.n375 VSUBS 0.008194f
C429 B.n376 VSUBS 0.008194f
C430 B.n377 VSUBS 0.008194f
C431 B.n378 VSUBS 0.008194f
C432 B.n379 VSUBS 0.008194f
C433 B.n380 VSUBS 0.008194f
C434 B.n381 VSUBS 0.008194f
C435 B.n382 VSUBS 0.008194f
C436 B.n383 VSUBS 0.008194f
C437 B.n384 VSUBS 0.008194f
C438 B.n385 VSUBS 0.008194f
C439 B.n386 VSUBS 0.008194f
C440 B.n387 VSUBS 0.008194f
C441 B.n388 VSUBS 0.008194f
C442 B.n389 VSUBS 0.008194f
C443 B.n390 VSUBS 0.008194f
C444 B.n391 VSUBS 0.008194f
C445 B.n392 VSUBS 0.008194f
C446 B.n393 VSUBS 0.008194f
C447 B.n394 VSUBS 0.008194f
C448 B.n395 VSUBS 0.008194f
C449 B.n396 VSUBS 0.008194f
C450 B.n397 VSUBS 0.008194f
C451 B.n398 VSUBS 0.008194f
C452 B.n399 VSUBS 0.008194f
C453 B.n400 VSUBS 0.008194f
C454 B.n401 VSUBS 0.008194f
C455 B.n402 VSUBS 0.008194f
C456 B.n403 VSUBS 0.008194f
C457 B.n404 VSUBS 0.008194f
C458 B.n405 VSUBS 0.008194f
C459 B.n406 VSUBS 0.008194f
C460 B.n407 VSUBS 0.008194f
C461 B.n408 VSUBS 0.008194f
C462 B.n409 VSUBS 0.008194f
C463 B.n410 VSUBS 0.008194f
C464 B.n411 VSUBS 0.020519f
C465 B.n412 VSUBS 0.019594f
C466 B.n413 VSUBS 0.019932f
C467 B.n414 VSUBS 0.008194f
C468 B.n415 VSUBS 0.008194f
C469 B.n416 VSUBS 0.008194f
C470 B.n417 VSUBS 0.008194f
C471 B.n418 VSUBS 0.008194f
C472 B.n419 VSUBS 0.008194f
C473 B.n420 VSUBS 0.008194f
C474 B.n421 VSUBS 0.008194f
C475 B.n422 VSUBS 0.008194f
C476 B.n423 VSUBS 0.008194f
C477 B.n424 VSUBS 0.008194f
C478 B.n425 VSUBS 0.008194f
C479 B.n426 VSUBS 0.008194f
C480 B.n427 VSUBS 0.008194f
C481 B.n428 VSUBS 0.008194f
C482 B.n429 VSUBS 0.008194f
C483 B.n430 VSUBS 0.008194f
C484 B.n431 VSUBS 0.008194f
C485 B.n432 VSUBS 0.008194f
C486 B.n433 VSUBS 0.008194f
C487 B.n434 VSUBS 0.008194f
C488 B.n435 VSUBS 0.008194f
C489 B.n436 VSUBS 0.008194f
C490 B.n437 VSUBS 0.008194f
C491 B.n438 VSUBS 0.008194f
C492 B.n439 VSUBS 0.008194f
C493 B.n440 VSUBS 0.008194f
C494 B.n441 VSUBS 0.008194f
C495 B.n442 VSUBS 0.008194f
C496 B.n443 VSUBS 0.008194f
C497 B.n444 VSUBS 0.008194f
C498 B.n445 VSUBS 0.008194f
C499 B.n446 VSUBS 0.008194f
C500 B.n447 VSUBS 0.008194f
C501 B.n448 VSUBS 0.008194f
C502 B.n449 VSUBS 0.008194f
C503 B.n450 VSUBS 0.008194f
C504 B.n451 VSUBS 0.008194f
C505 B.n452 VSUBS 0.008194f
C506 B.n453 VSUBS 0.008194f
C507 B.n454 VSUBS 0.008194f
C508 B.n455 VSUBS 0.008194f
C509 B.n456 VSUBS 0.008194f
C510 B.n457 VSUBS 0.008194f
C511 B.n458 VSUBS 0.008194f
C512 B.n459 VSUBS 0.008194f
C513 B.n460 VSUBS 0.008194f
C514 B.n461 VSUBS 0.008194f
C515 B.n462 VSUBS 0.008194f
C516 B.n463 VSUBS 0.008194f
C517 B.n464 VSUBS 0.008194f
C518 B.n465 VSUBS 0.008194f
C519 B.n466 VSUBS 0.008194f
C520 B.n467 VSUBS 0.008194f
C521 B.n468 VSUBS 0.008194f
C522 B.n469 VSUBS 0.008194f
C523 B.n470 VSUBS 0.008194f
C524 B.n471 VSUBS 0.008194f
C525 B.n472 VSUBS 0.008194f
C526 B.n473 VSUBS 0.008194f
C527 B.n474 VSUBS 0.008194f
C528 B.n475 VSUBS 0.008194f
C529 B.n476 VSUBS 0.008194f
C530 B.n477 VSUBS 0.008194f
C531 B.n478 VSUBS 0.008194f
C532 B.n479 VSUBS 0.008194f
C533 B.n480 VSUBS 0.008194f
C534 B.n481 VSUBS 0.008194f
C535 B.n482 VSUBS 0.008194f
C536 B.n483 VSUBS 0.008194f
C537 B.n484 VSUBS 0.008194f
C538 B.n485 VSUBS 0.008194f
C539 B.n486 VSUBS 0.008194f
C540 B.n487 VSUBS 0.008194f
C541 B.n488 VSUBS 0.008194f
C542 B.n489 VSUBS 0.008194f
C543 B.n490 VSUBS 0.008194f
C544 B.n491 VSUBS 0.008194f
C545 B.n492 VSUBS 0.008194f
C546 B.n493 VSUBS 0.008194f
C547 B.n494 VSUBS 0.008194f
C548 B.n495 VSUBS 0.005664f
C549 B.n496 VSUBS 0.008194f
C550 B.n497 VSUBS 0.008194f
C551 B.n498 VSUBS 0.006628f
C552 B.n499 VSUBS 0.008194f
C553 B.n500 VSUBS 0.008194f
C554 B.n501 VSUBS 0.008194f
C555 B.n502 VSUBS 0.008194f
C556 B.n503 VSUBS 0.008194f
C557 B.n504 VSUBS 0.008194f
C558 B.n505 VSUBS 0.008194f
C559 B.n506 VSUBS 0.008194f
C560 B.n507 VSUBS 0.008194f
C561 B.n508 VSUBS 0.008194f
C562 B.n509 VSUBS 0.008194f
C563 B.n510 VSUBS 0.006628f
C564 B.n511 VSUBS 0.018986f
C565 B.n512 VSUBS 0.005664f
C566 B.n513 VSUBS 0.008194f
C567 B.n514 VSUBS 0.008194f
C568 B.n515 VSUBS 0.008194f
C569 B.n516 VSUBS 0.008194f
C570 B.n517 VSUBS 0.008194f
C571 B.n518 VSUBS 0.008194f
C572 B.n519 VSUBS 0.008194f
C573 B.n520 VSUBS 0.008194f
C574 B.n521 VSUBS 0.008194f
C575 B.n522 VSUBS 0.008194f
C576 B.n523 VSUBS 0.008194f
C577 B.n524 VSUBS 0.008194f
C578 B.n525 VSUBS 0.008194f
C579 B.n526 VSUBS 0.008194f
C580 B.n527 VSUBS 0.008194f
C581 B.n528 VSUBS 0.008194f
C582 B.n529 VSUBS 0.008194f
C583 B.n530 VSUBS 0.008194f
C584 B.n531 VSUBS 0.008194f
C585 B.n532 VSUBS 0.008194f
C586 B.n533 VSUBS 0.008194f
C587 B.n534 VSUBS 0.008194f
C588 B.n535 VSUBS 0.008194f
C589 B.n536 VSUBS 0.008194f
C590 B.n537 VSUBS 0.008194f
C591 B.n538 VSUBS 0.008194f
C592 B.n539 VSUBS 0.008194f
C593 B.n540 VSUBS 0.008194f
C594 B.n541 VSUBS 0.008194f
C595 B.n542 VSUBS 0.008194f
C596 B.n543 VSUBS 0.008194f
C597 B.n544 VSUBS 0.008194f
C598 B.n545 VSUBS 0.008194f
C599 B.n546 VSUBS 0.008194f
C600 B.n547 VSUBS 0.008194f
C601 B.n548 VSUBS 0.008194f
C602 B.n549 VSUBS 0.008194f
C603 B.n550 VSUBS 0.008194f
C604 B.n551 VSUBS 0.008194f
C605 B.n552 VSUBS 0.008194f
C606 B.n553 VSUBS 0.008194f
C607 B.n554 VSUBS 0.008194f
C608 B.n555 VSUBS 0.008194f
C609 B.n556 VSUBS 0.008194f
C610 B.n557 VSUBS 0.008194f
C611 B.n558 VSUBS 0.008194f
C612 B.n559 VSUBS 0.008194f
C613 B.n560 VSUBS 0.008194f
C614 B.n561 VSUBS 0.008194f
C615 B.n562 VSUBS 0.008194f
C616 B.n563 VSUBS 0.008194f
C617 B.n564 VSUBS 0.008194f
C618 B.n565 VSUBS 0.008194f
C619 B.n566 VSUBS 0.008194f
C620 B.n567 VSUBS 0.008194f
C621 B.n568 VSUBS 0.008194f
C622 B.n569 VSUBS 0.008194f
C623 B.n570 VSUBS 0.008194f
C624 B.n571 VSUBS 0.008194f
C625 B.n572 VSUBS 0.008194f
C626 B.n573 VSUBS 0.008194f
C627 B.n574 VSUBS 0.008194f
C628 B.n575 VSUBS 0.008194f
C629 B.n576 VSUBS 0.008194f
C630 B.n577 VSUBS 0.008194f
C631 B.n578 VSUBS 0.008194f
C632 B.n579 VSUBS 0.008194f
C633 B.n580 VSUBS 0.008194f
C634 B.n581 VSUBS 0.008194f
C635 B.n582 VSUBS 0.008194f
C636 B.n583 VSUBS 0.008194f
C637 B.n584 VSUBS 0.008194f
C638 B.n585 VSUBS 0.008194f
C639 B.n586 VSUBS 0.008194f
C640 B.n587 VSUBS 0.008194f
C641 B.n588 VSUBS 0.008194f
C642 B.n589 VSUBS 0.008194f
C643 B.n590 VSUBS 0.008194f
C644 B.n591 VSUBS 0.008194f
C645 B.n592 VSUBS 0.008194f
C646 B.n593 VSUBS 0.008194f
C647 B.n594 VSUBS 0.019932f
C648 B.n595 VSUBS 0.019932f
C649 B.n596 VSUBS 0.019594f
C650 B.n597 VSUBS 0.008194f
C651 B.n598 VSUBS 0.008194f
C652 B.n599 VSUBS 0.008194f
C653 B.n600 VSUBS 0.008194f
C654 B.n601 VSUBS 0.008194f
C655 B.n602 VSUBS 0.008194f
C656 B.n603 VSUBS 0.008194f
C657 B.n604 VSUBS 0.008194f
C658 B.n605 VSUBS 0.008194f
C659 B.n606 VSUBS 0.008194f
C660 B.n607 VSUBS 0.008194f
C661 B.n608 VSUBS 0.008194f
C662 B.n609 VSUBS 0.008194f
C663 B.n610 VSUBS 0.008194f
C664 B.n611 VSUBS 0.008194f
C665 B.n612 VSUBS 0.008194f
C666 B.n613 VSUBS 0.008194f
C667 B.n614 VSUBS 0.008194f
C668 B.n615 VSUBS 0.008194f
C669 B.n616 VSUBS 0.008194f
C670 B.n617 VSUBS 0.008194f
C671 B.n618 VSUBS 0.008194f
C672 B.n619 VSUBS 0.018555f
C673 VDD1.t0 VSUBS 0.408587f
C674 VDD1.t3 VSUBS 0.408587f
C675 VDD1.n0 VSUBS 3.37527f
C676 VDD1.t2 VSUBS 0.408587f
C677 VDD1.t1 VSUBS 0.408587f
C678 VDD1.n1 VSUBS 4.29402f
C679 VTAIL.n0 VSUBS 0.026031f
C680 VTAIL.n1 VSUBS 0.023781f
C681 VTAIL.n2 VSUBS 0.012779f
C682 VTAIL.n3 VSUBS 0.030204f
C683 VTAIL.n4 VSUBS 0.013531f
C684 VTAIL.n5 VSUBS 0.023781f
C685 VTAIL.n6 VSUBS 0.012779f
C686 VTAIL.n7 VSUBS 0.030204f
C687 VTAIL.n8 VSUBS 0.013531f
C688 VTAIL.n9 VSUBS 0.023781f
C689 VTAIL.n10 VSUBS 0.012779f
C690 VTAIL.n11 VSUBS 0.030204f
C691 VTAIL.n12 VSUBS 0.013531f
C692 VTAIL.n13 VSUBS 0.023781f
C693 VTAIL.n14 VSUBS 0.012779f
C694 VTAIL.n15 VSUBS 0.030204f
C695 VTAIL.n16 VSUBS 0.013531f
C696 VTAIL.n17 VSUBS 0.023781f
C697 VTAIL.n18 VSUBS 0.012779f
C698 VTAIL.n19 VSUBS 0.030204f
C699 VTAIL.n20 VSUBS 0.013531f
C700 VTAIL.n21 VSUBS 0.023781f
C701 VTAIL.n22 VSUBS 0.012779f
C702 VTAIL.n23 VSUBS 0.030204f
C703 VTAIL.n24 VSUBS 0.013531f
C704 VTAIL.n25 VSUBS 0.023781f
C705 VTAIL.n26 VSUBS 0.012779f
C706 VTAIL.n27 VSUBS 0.030204f
C707 VTAIL.n28 VSUBS 0.013531f
C708 VTAIL.n29 VSUBS 0.180821f
C709 VTAIL.t0 VSUBS 0.064773f
C710 VTAIL.n30 VSUBS 0.022653f
C711 VTAIL.n31 VSUBS 0.019215f
C712 VTAIL.n32 VSUBS 0.012779f
C713 VTAIL.n33 VSUBS 1.72141f
C714 VTAIL.n34 VSUBS 0.023781f
C715 VTAIL.n35 VSUBS 0.012779f
C716 VTAIL.n36 VSUBS 0.013531f
C717 VTAIL.n37 VSUBS 0.030204f
C718 VTAIL.n38 VSUBS 0.030204f
C719 VTAIL.n39 VSUBS 0.013531f
C720 VTAIL.n40 VSUBS 0.012779f
C721 VTAIL.n41 VSUBS 0.023781f
C722 VTAIL.n42 VSUBS 0.023781f
C723 VTAIL.n43 VSUBS 0.012779f
C724 VTAIL.n44 VSUBS 0.013531f
C725 VTAIL.n45 VSUBS 0.030204f
C726 VTAIL.n46 VSUBS 0.030204f
C727 VTAIL.n47 VSUBS 0.013531f
C728 VTAIL.n48 VSUBS 0.012779f
C729 VTAIL.n49 VSUBS 0.023781f
C730 VTAIL.n50 VSUBS 0.023781f
C731 VTAIL.n51 VSUBS 0.012779f
C732 VTAIL.n52 VSUBS 0.013531f
C733 VTAIL.n53 VSUBS 0.030204f
C734 VTAIL.n54 VSUBS 0.030204f
C735 VTAIL.n55 VSUBS 0.013531f
C736 VTAIL.n56 VSUBS 0.012779f
C737 VTAIL.n57 VSUBS 0.023781f
C738 VTAIL.n58 VSUBS 0.023781f
C739 VTAIL.n59 VSUBS 0.012779f
C740 VTAIL.n60 VSUBS 0.013531f
C741 VTAIL.n61 VSUBS 0.030204f
C742 VTAIL.n62 VSUBS 0.030204f
C743 VTAIL.n63 VSUBS 0.013531f
C744 VTAIL.n64 VSUBS 0.012779f
C745 VTAIL.n65 VSUBS 0.023781f
C746 VTAIL.n66 VSUBS 0.023781f
C747 VTAIL.n67 VSUBS 0.012779f
C748 VTAIL.n68 VSUBS 0.013531f
C749 VTAIL.n69 VSUBS 0.030204f
C750 VTAIL.n70 VSUBS 0.030204f
C751 VTAIL.n71 VSUBS 0.030204f
C752 VTAIL.n72 VSUBS 0.013531f
C753 VTAIL.n73 VSUBS 0.012779f
C754 VTAIL.n74 VSUBS 0.023781f
C755 VTAIL.n75 VSUBS 0.023781f
C756 VTAIL.n76 VSUBS 0.012779f
C757 VTAIL.n77 VSUBS 0.013155f
C758 VTAIL.n78 VSUBS 0.013155f
C759 VTAIL.n79 VSUBS 0.030204f
C760 VTAIL.n80 VSUBS 0.030204f
C761 VTAIL.n81 VSUBS 0.013531f
C762 VTAIL.n82 VSUBS 0.012779f
C763 VTAIL.n83 VSUBS 0.023781f
C764 VTAIL.n84 VSUBS 0.023781f
C765 VTAIL.n85 VSUBS 0.012779f
C766 VTAIL.n86 VSUBS 0.013531f
C767 VTAIL.n87 VSUBS 0.030204f
C768 VTAIL.n88 VSUBS 0.072783f
C769 VTAIL.n89 VSUBS 0.013531f
C770 VTAIL.n90 VSUBS 0.012779f
C771 VTAIL.n91 VSUBS 0.057567f
C772 VTAIL.n92 VSUBS 0.036665f
C773 VTAIL.n93 VSUBS 0.087672f
C774 VTAIL.n94 VSUBS 0.026031f
C775 VTAIL.n95 VSUBS 0.023781f
C776 VTAIL.n96 VSUBS 0.012779f
C777 VTAIL.n97 VSUBS 0.030204f
C778 VTAIL.n98 VSUBS 0.013531f
C779 VTAIL.n99 VSUBS 0.023781f
C780 VTAIL.n100 VSUBS 0.012779f
C781 VTAIL.n101 VSUBS 0.030204f
C782 VTAIL.n102 VSUBS 0.013531f
C783 VTAIL.n103 VSUBS 0.023781f
C784 VTAIL.n104 VSUBS 0.012779f
C785 VTAIL.n105 VSUBS 0.030204f
C786 VTAIL.n106 VSUBS 0.013531f
C787 VTAIL.n107 VSUBS 0.023781f
C788 VTAIL.n108 VSUBS 0.012779f
C789 VTAIL.n109 VSUBS 0.030204f
C790 VTAIL.n110 VSUBS 0.013531f
C791 VTAIL.n111 VSUBS 0.023781f
C792 VTAIL.n112 VSUBS 0.012779f
C793 VTAIL.n113 VSUBS 0.030204f
C794 VTAIL.n114 VSUBS 0.013531f
C795 VTAIL.n115 VSUBS 0.023781f
C796 VTAIL.n116 VSUBS 0.012779f
C797 VTAIL.n117 VSUBS 0.030204f
C798 VTAIL.n118 VSUBS 0.013531f
C799 VTAIL.n119 VSUBS 0.023781f
C800 VTAIL.n120 VSUBS 0.012779f
C801 VTAIL.n121 VSUBS 0.030204f
C802 VTAIL.n122 VSUBS 0.013531f
C803 VTAIL.n123 VSUBS 0.180821f
C804 VTAIL.t5 VSUBS 0.064773f
C805 VTAIL.n124 VSUBS 0.022653f
C806 VTAIL.n125 VSUBS 0.019215f
C807 VTAIL.n126 VSUBS 0.012779f
C808 VTAIL.n127 VSUBS 1.72141f
C809 VTAIL.n128 VSUBS 0.023781f
C810 VTAIL.n129 VSUBS 0.012779f
C811 VTAIL.n130 VSUBS 0.013531f
C812 VTAIL.n131 VSUBS 0.030204f
C813 VTAIL.n132 VSUBS 0.030204f
C814 VTAIL.n133 VSUBS 0.013531f
C815 VTAIL.n134 VSUBS 0.012779f
C816 VTAIL.n135 VSUBS 0.023781f
C817 VTAIL.n136 VSUBS 0.023781f
C818 VTAIL.n137 VSUBS 0.012779f
C819 VTAIL.n138 VSUBS 0.013531f
C820 VTAIL.n139 VSUBS 0.030204f
C821 VTAIL.n140 VSUBS 0.030204f
C822 VTAIL.n141 VSUBS 0.013531f
C823 VTAIL.n142 VSUBS 0.012779f
C824 VTAIL.n143 VSUBS 0.023781f
C825 VTAIL.n144 VSUBS 0.023781f
C826 VTAIL.n145 VSUBS 0.012779f
C827 VTAIL.n146 VSUBS 0.013531f
C828 VTAIL.n147 VSUBS 0.030204f
C829 VTAIL.n148 VSUBS 0.030204f
C830 VTAIL.n149 VSUBS 0.013531f
C831 VTAIL.n150 VSUBS 0.012779f
C832 VTAIL.n151 VSUBS 0.023781f
C833 VTAIL.n152 VSUBS 0.023781f
C834 VTAIL.n153 VSUBS 0.012779f
C835 VTAIL.n154 VSUBS 0.013531f
C836 VTAIL.n155 VSUBS 0.030204f
C837 VTAIL.n156 VSUBS 0.030204f
C838 VTAIL.n157 VSUBS 0.013531f
C839 VTAIL.n158 VSUBS 0.012779f
C840 VTAIL.n159 VSUBS 0.023781f
C841 VTAIL.n160 VSUBS 0.023781f
C842 VTAIL.n161 VSUBS 0.012779f
C843 VTAIL.n162 VSUBS 0.013531f
C844 VTAIL.n163 VSUBS 0.030204f
C845 VTAIL.n164 VSUBS 0.030204f
C846 VTAIL.n165 VSUBS 0.030204f
C847 VTAIL.n166 VSUBS 0.013531f
C848 VTAIL.n167 VSUBS 0.012779f
C849 VTAIL.n168 VSUBS 0.023781f
C850 VTAIL.n169 VSUBS 0.023781f
C851 VTAIL.n170 VSUBS 0.012779f
C852 VTAIL.n171 VSUBS 0.013155f
C853 VTAIL.n172 VSUBS 0.013155f
C854 VTAIL.n173 VSUBS 0.030204f
C855 VTAIL.n174 VSUBS 0.030204f
C856 VTAIL.n175 VSUBS 0.013531f
C857 VTAIL.n176 VSUBS 0.012779f
C858 VTAIL.n177 VSUBS 0.023781f
C859 VTAIL.n178 VSUBS 0.023781f
C860 VTAIL.n179 VSUBS 0.012779f
C861 VTAIL.n180 VSUBS 0.013531f
C862 VTAIL.n181 VSUBS 0.030204f
C863 VTAIL.n182 VSUBS 0.072783f
C864 VTAIL.n183 VSUBS 0.013531f
C865 VTAIL.n184 VSUBS 0.012779f
C866 VTAIL.n185 VSUBS 0.057567f
C867 VTAIL.n186 VSUBS 0.036665f
C868 VTAIL.n187 VSUBS 0.108645f
C869 VTAIL.n188 VSUBS 0.026031f
C870 VTAIL.n189 VSUBS 0.023781f
C871 VTAIL.n190 VSUBS 0.012779f
C872 VTAIL.n191 VSUBS 0.030204f
C873 VTAIL.n192 VSUBS 0.013531f
C874 VTAIL.n193 VSUBS 0.023781f
C875 VTAIL.n194 VSUBS 0.012779f
C876 VTAIL.n195 VSUBS 0.030204f
C877 VTAIL.n196 VSUBS 0.013531f
C878 VTAIL.n197 VSUBS 0.023781f
C879 VTAIL.n198 VSUBS 0.012779f
C880 VTAIL.n199 VSUBS 0.030204f
C881 VTAIL.n200 VSUBS 0.013531f
C882 VTAIL.n201 VSUBS 0.023781f
C883 VTAIL.n202 VSUBS 0.012779f
C884 VTAIL.n203 VSUBS 0.030204f
C885 VTAIL.n204 VSUBS 0.013531f
C886 VTAIL.n205 VSUBS 0.023781f
C887 VTAIL.n206 VSUBS 0.012779f
C888 VTAIL.n207 VSUBS 0.030204f
C889 VTAIL.n208 VSUBS 0.013531f
C890 VTAIL.n209 VSUBS 0.023781f
C891 VTAIL.n210 VSUBS 0.012779f
C892 VTAIL.n211 VSUBS 0.030204f
C893 VTAIL.n212 VSUBS 0.013531f
C894 VTAIL.n213 VSUBS 0.023781f
C895 VTAIL.n214 VSUBS 0.012779f
C896 VTAIL.n215 VSUBS 0.030204f
C897 VTAIL.n216 VSUBS 0.013531f
C898 VTAIL.n217 VSUBS 0.180821f
C899 VTAIL.t4 VSUBS 0.064773f
C900 VTAIL.n218 VSUBS 0.022653f
C901 VTAIL.n219 VSUBS 0.019215f
C902 VTAIL.n220 VSUBS 0.012779f
C903 VTAIL.n221 VSUBS 1.72141f
C904 VTAIL.n222 VSUBS 0.023781f
C905 VTAIL.n223 VSUBS 0.012779f
C906 VTAIL.n224 VSUBS 0.013531f
C907 VTAIL.n225 VSUBS 0.030204f
C908 VTAIL.n226 VSUBS 0.030204f
C909 VTAIL.n227 VSUBS 0.013531f
C910 VTAIL.n228 VSUBS 0.012779f
C911 VTAIL.n229 VSUBS 0.023781f
C912 VTAIL.n230 VSUBS 0.023781f
C913 VTAIL.n231 VSUBS 0.012779f
C914 VTAIL.n232 VSUBS 0.013531f
C915 VTAIL.n233 VSUBS 0.030204f
C916 VTAIL.n234 VSUBS 0.030204f
C917 VTAIL.n235 VSUBS 0.013531f
C918 VTAIL.n236 VSUBS 0.012779f
C919 VTAIL.n237 VSUBS 0.023781f
C920 VTAIL.n238 VSUBS 0.023781f
C921 VTAIL.n239 VSUBS 0.012779f
C922 VTAIL.n240 VSUBS 0.013531f
C923 VTAIL.n241 VSUBS 0.030204f
C924 VTAIL.n242 VSUBS 0.030204f
C925 VTAIL.n243 VSUBS 0.013531f
C926 VTAIL.n244 VSUBS 0.012779f
C927 VTAIL.n245 VSUBS 0.023781f
C928 VTAIL.n246 VSUBS 0.023781f
C929 VTAIL.n247 VSUBS 0.012779f
C930 VTAIL.n248 VSUBS 0.013531f
C931 VTAIL.n249 VSUBS 0.030204f
C932 VTAIL.n250 VSUBS 0.030204f
C933 VTAIL.n251 VSUBS 0.013531f
C934 VTAIL.n252 VSUBS 0.012779f
C935 VTAIL.n253 VSUBS 0.023781f
C936 VTAIL.n254 VSUBS 0.023781f
C937 VTAIL.n255 VSUBS 0.012779f
C938 VTAIL.n256 VSUBS 0.013531f
C939 VTAIL.n257 VSUBS 0.030204f
C940 VTAIL.n258 VSUBS 0.030204f
C941 VTAIL.n259 VSUBS 0.030204f
C942 VTAIL.n260 VSUBS 0.013531f
C943 VTAIL.n261 VSUBS 0.012779f
C944 VTAIL.n262 VSUBS 0.023781f
C945 VTAIL.n263 VSUBS 0.023781f
C946 VTAIL.n264 VSUBS 0.012779f
C947 VTAIL.n265 VSUBS 0.013155f
C948 VTAIL.n266 VSUBS 0.013155f
C949 VTAIL.n267 VSUBS 0.030204f
C950 VTAIL.n268 VSUBS 0.030204f
C951 VTAIL.n269 VSUBS 0.013531f
C952 VTAIL.n270 VSUBS 0.012779f
C953 VTAIL.n271 VSUBS 0.023781f
C954 VTAIL.n272 VSUBS 0.023781f
C955 VTAIL.n273 VSUBS 0.012779f
C956 VTAIL.n274 VSUBS 0.013531f
C957 VTAIL.n275 VSUBS 0.030204f
C958 VTAIL.n276 VSUBS 0.072783f
C959 VTAIL.n277 VSUBS 0.013531f
C960 VTAIL.n278 VSUBS 0.012779f
C961 VTAIL.n279 VSUBS 0.057567f
C962 VTAIL.n280 VSUBS 0.036665f
C963 VTAIL.n281 VSUBS 1.5616f
C964 VTAIL.n282 VSUBS 0.026031f
C965 VTAIL.n283 VSUBS 0.023781f
C966 VTAIL.n284 VSUBS 0.012779f
C967 VTAIL.n285 VSUBS 0.030204f
C968 VTAIL.n286 VSUBS 0.013531f
C969 VTAIL.n287 VSUBS 0.023781f
C970 VTAIL.n288 VSUBS 0.012779f
C971 VTAIL.n289 VSUBS 0.030204f
C972 VTAIL.n290 VSUBS 0.013531f
C973 VTAIL.n291 VSUBS 0.023781f
C974 VTAIL.n292 VSUBS 0.012779f
C975 VTAIL.n293 VSUBS 0.030204f
C976 VTAIL.n294 VSUBS 0.030204f
C977 VTAIL.n295 VSUBS 0.013531f
C978 VTAIL.n296 VSUBS 0.023781f
C979 VTAIL.n297 VSUBS 0.012779f
C980 VTAIL.n298 VSUBS 0.030204f
C981 VTAIL.n299 VSUBS 0.013531f
C982 VTAIL.n300 VSUBS 0.023781f
C983 VTAIL.n301 VSUBS 0.012779f
C984 VTAIL.n302 VSUBS 0.030204f
C985 VTAIL.n303 VSUBS 0.013531f
C986 VTAIL.n304 VSUBS 0.023781f
C987 VTAIL.n305 VSUBS 0.012779f
C988 VTAIL.n306 VSUBS 0.030204f
C989 VTAIL.n307 VSUBS 0.013531f
C990 VTAIL.n308 VSUBS 0.023781f
C991 VTAIL.n309 VSUBS 0.012779f
C992 VTAIL.n310 VSUBS 0.030204f
C993 VTAIL.n311 VSUBS 0.013531f
C994 VTAIL.n312 VSUBS 0.180821f
C995 VTAIL.t3 VSUBS 0.064773f
C996 VTAIL.n313 VSUBS 0.022653f
C997 VTAIL.n314 VSUBS 0.019215f
C998 VTAIL.n315 VSUBS 0.012779f
C999 VTAIL.n316 VSUBS 1.72141f
C1000 VTAIL.n317 VSUBS 0.023781f
C1001 VTAIL.n318 VSUBS 0.012779f
C1002 VTAIL.n319 VSUBS 0.013531f
C1003 VTAIL.n320 VSUBS 0.030204f
C1004 VTAIL.n321 VSUBS 0.030204f
C1005 VTAIL.n322 VSUBS 0.013531f
C1006 VTAIL.n323 VSUBS 0.012779f
C1007 VTAIL.n324 VSUBS 0.023781f
C1008 VTAIL.n325 VSUBS 0.023781f
C1009 VTAIL.n326 VSUBS 0.012779f
C1010 VTAIL.n327 VSUBS 0.013531f
C1011 VTAIL.n328 VSUBS 0.030204f
C1012 VTAIL.n329 VSUBS 0.030204f
C1013 VTAIL.n330 VSUBS 0.013531f
C1014 VTAIL.n331 VSUBS 0.012779f
C1015 VTAIL.n332 VSUBS 0.023781f
C1016 VTAIL.n333 VSUBS 0.023781f
C1017 VTAIL.n334 VSUBS 0.012779f
C1018 VTAIL.n335 VSUBS 0.013531f
C1019 VTAIL.n336 VSUBS 0.030204f
C1020 VTAIL.n337 VSUBS 0.030204f
C1021 VTAIL.n338 VSUBS 0.013531f
C1022 VTAIL.n339 VSUBS 0.012779f
C1023 VTAIL.n340 VSUBS 0.023781f
C1024 VTAIL.n341 VSUBS 0.023781f
C1025 VTAIL.n342 VSUBS 0.012779f
C1026 VTAIL.n343 VSUBS 0.013531f
C1027 VTAIL.n344 VSUBS 0.030204f
C1028 VTAIL.n345 VSUBS 0.030204f
C1029 VTAIL.n346 VSUBS 0.013531f
C1030 VTAIL.n347 VSUBS 0.012779f
C1031 VTAIL.n348 VSUBS 0.023781f
C1032 VTAIL.n349 VSUBS 0.023781f
C1033 VTAIL.n350 VSUBS 0.012779f
C1034 VTAIL.n351 VSUBS 0.013531f
C1035 VTAIL.n352 VSUBS 0.030204f
C1036 VTAIL.n353 VSUBS 0.030204f
C1037 VTAIL.n354 VSUBS 0.013531f
C1038 VTAIL.n355 VSUBS 0.012779f
C1039 VTAIL.n356 VSUBS 0.023781f
C1040 VTAIL.n357 VSUBS 0.023781f
C1041 VTAIL.n358 VSUBS 0.012779f
C1042 VTAIL.n359 VSUBS 0.013155f
C1043 VTAIL.n360 VSUBS 0.013155f
C1044 VTAIL.n361 VSUBS 0.030204f
C1045 VTAIL.n362 VSUBS 0.030204f
C1046 VTAIL.n363 VSUBS 0.013531f
C1047 VTAIL.n364 VSUBS 0.012779f
C1048 VTAIL.n365 VSUBS 0.023781f
C1049 VTAIL.n366 VSUBS 0.023781f
C1050 VTAIL.n367 VSUBS 0.012779f
C1051 VTAIL.n368 VSUBS 0.013531f
C1052 VTAIL.n369 VSUBS 0.030204f
C1053 VTAIL.n370 VSUBS 0.072783f
C1054 VTAIL.n371 VSUBS 0.013531f
C1055 VTAIL.n372 VSUBS 0.012779f
C1056 VTAIL.n373 VSUBS 0.057567f
C1057 VTAIL.n374 VSUBS 0.036665f
C1058 VTAIL.n375 VSUBS 1.5616f
C1059 VTAIL.n376 VSUBS 0.026031f
C1060 VTAIL.n377 VSUBS 0.023781f
C1061 VTAIL.n378 VSUBS 0.012779f
C1062 VTAIL.n379 VSUBS 0.030204f
C1063 VTAIL.n380 VSUBS 0.013531f
C1064 VTAIL.n381 VSUBS 0.023781f
C1065 VTAIL.n382 VSUBS 0.012779f
C1066 VTAIL.n383 VSUBS 0.030204f
C1067 VTAIL.n384 VSUBS 0.013531f
C1068 VTAIL.n385 VSUBS 0.023781f
C1069 VTAIL.n386 VSUBS 0.012779f
C1070 VTAIL.n387 VSUBS 0.030204f
C1071 VTAIL.n388 VSUBS 0.030204f
C1072 VTAIL.n389 VSUBS 0.013531f
C1073 VTAIL.n390 VSUBS 0.023781f
C1074 VTAIL.n391 VSUBS 0.012779f
C1075 VTAIL.n392 VSUBS 0.030204f
C1076 VTAIL.n393 VSUBS 0.013531f
C1077 VTAIL.n394 VSUBS 0.023781f
C1078 VTAIL.n395 VSUBS 0.012779f
C1079 VTAIL.n396 VSUBS 0.030204f
C1080 VTAIL.n397 VSUBS 0.013531f
C1081 VTAIL.n398 VSUBS 0.023781f
C1082 VTAIL.n399 VSUBS 0.012779f
C1083 VTAIL.n400 VSUBS 0.030204f
C1084 VTAIL.n401 VSUBS 0.013531f
C1085 VTAIL.n402 VSUBS 0.023781f
C1086 VTAIL.n403 VSUBS 0.012779f
C1087 VTAIL.n404 VSUBS 0.030204f
C1088 VTAIL.n405 VSUBS 0.013531f
C1089 VTAIL.n406 VSUBS 0.180821f
C1090 VTAIL.t1 VSUBS 0.064773f
C1091 VTAIL.n407 VSUBS 0.022653f
C1092 VTAIL.n408 VSUBS 0.019215f
C1093 VTAIL.n409 VSUBS 0.012779f
C1094 VTAIL.n410 VSUBS 1.72141f
C1095 VTAIL.n411 VSUBS 0.023781f
C1096 VTAIL.n412 VSUBS 0.012779f
C1097 VTAIL.n413 VSUBS 0.013531f
C1098 VTAIL.n414 VSUBS 0.030204f
C1099 VTAIL.n415 VSUBS 0.030204f
C1100 VTAIL.n416 VSUBS 0.013531f
C1101 VTAIL.n417 VSUBS 0.012779f
C1102 VTAIL.n418 VSUBS 0.023781f
C1103 VTAIL.n419 VSUBS 0.023781f
C1104 VTAIL.n420 VSUBS 0.012779f
C1105 VTAIL.n421 VSUBS 0.013531f
C1106 VTAIL.n422 VSUBS 0.030204f
C1107 VTAIL.n423 VSUBS 0.030204f
C1108 VTAIL.n424 VSUBS 0.013531f
C1109 VTAIL.n425 VSUBS 0.012779f
C1110 VTAIL.n426 VSUBS 0.023781f
C1111 VTAIL.n427 VSUBS 0.023781f
C1112 VTAIL.n428 VSUBS 0.012779f
C1113 VTAIL.n429 VSUBS 0.013531f
C1114 VTAIL.n430 VSUBS 0.030204f
C1115 VTAIL.n431 VSUBS 0.030204f
C1116 VTAIL.n432 VSUBS 0.013531f
C1117 VTAIL.n433 VSUBS 0.012779f
C1118 VTAIL.n434 VSUBS 0.023781f
C1119 VTAIL.n435 VSUBS 0.023781f
C1120 VTAIL.n436 VSUBS 0.012779f
C1121 VTAIL.n437 VSUBS 0.013531f
C1122 VTAIL.n438 VSUBS 0.030204f
C1123 VTAIL.n439 VSUBS 0.030204f
C1124 VTAIL.n440 VSUBS 0.013531f
C1125 VTAIL.n441 VSUBS 0.012779f
C1126 VTAIL.n442 VSUBS 0.023781f
C1127 VTAIL.n443 VSUBS 0.023781f
C1128 VTAIL.n444 VSUBS 0.012779f
C1129 VTAIL.n445 VSUBS 0.013531f
C1130 VTAIL.n446 VSUBS 0.030204f
C1131 VTAIL.n447 VSUBS 0.030204f
C1132 VTAIL.n448 VSUBS 0.013531f
C1133 VTAIL.n449 VSUBS 0.012779f
C1134 VTAIL.n450 VSUBS 0.023781f
C1135 VTAIL.n451 VSUBS 0.023781f
C1136 VTAIL.n452 VSUBS 0.012779f
C1137 VTAIL.n453 VSUBS 0.013155f
C1138 VTAIL.n454 VSUBS 0.013155f
C1139 VTAIL.n455 VSUBS 0.030204f
C1140 VTAIL.n456 VSUBS 0.030204f
C1141 VTAIL.n457 VSUBS 0.013531f
C1142 VTAIL.n458 VSUBS 0.012779f
C1143 VTAIL.n459 VSUBS 0.023781f
C1144 VTAIL.n460 VSUBS 0.023781f
C1145 VTAIL.n461 VSUBS 0.012779f
C1146 VTAIL.n462 VSUBS 0.013531f
C1147 VTAIL.n463 VSUBS 0.030204f
C1148 VTAIL.n464 VSUBS 0.072783f
C1149 VTAIL.n465 VSUBS 0.013531f
C1150 VTAIL.n466 VSUBS 0.012779f
C1151 VTAIL.n467 VSUBS 0.057567f
C1152 VTAIL.n468 VSUBS 0.036665f
C1153 VTAIL.n469 VSUBS 0.108645f
C1154 VTAIL.n470 VSUBS 0.026031f
C1155 VTAIL.n471 VSUBS 0.023781f
C1156 VTAIL.n472 VSUBS 0.012779f
C1157 VTAIL.n473 VSUBS 0.030204f
C1158 VTAIL.n474 VSUBS 0.013531f
C1159 VTAIL.n475 VSUBS 0.023781f
C1160 VTAIL.n476 VSUBS 0.012779f
C1161 VTAIL.n477 VSUBS 0.030204f
C1162 VTAIL.n478 VSUBS 0.013531f
C1163 VTAIL.n479 VSUBS 0.023781f
C1164 VTAIL.n480 VSUBS 0.012779f
C1165 VTAIL.n481 VSUBS 0.030204f
C1166 VTAIL.n482 VSUBS 0.030204f
C1167 VTAIL.n483 VSUBS 0.013531f
C1168 VTAIL.n484 VSUBS 0.023781f
C1169 VTAIL.n485 VSUBS 0.012779f
C1170 VTAIL.n486 VSUBS 0.030204f
C1171 VTAIL.n487 VSUBS 0.013531f
C1172 VTAIL.n488 VSUBS 0.023781f
C1173 VTAIL.n489 VSUBS 0.012779f
C1174 VTAIL.n490 VSUBS 0.030204f
C1175 VTAIL.n491 VSUBS 0.013531f
C1176 VTAIL.n492 VSUBS 0.023781f
C1177 VTAIL.n493 VSUBS 0.012779f
C1178 VTAIL.n494 VSUBS 0.030204f
C1179 VTAIL.n495 VSUBS 0.013531f
C1180 VTAIL.n496 VSUBS 0.023781f
C1181 VTAIL.n497 VSUBS 0.012779f
C1182 VTAIL.n498 VSUBS 0.030204f
C1183 VTAIL.n499 VSUBS 0.013531f
C1184 VTAIL.n500 VSUBS 0.180821f
C1185 VTAIL.t6 VSUBS 0.064773f
C1186 VTAIL.n501 VSUBS 0.022653f
C1187 VTAIL.n502 VSUBS 0.019215f
C1188 VTAIL.n503 VSUBS 0.012779f
C1189 VTAIL.n504 VSUBS 1.72141f
C1190 VTAIL.n505 VSUBS 0.023781f
C1191 VTAIL.n506 VSUBS 0.012779f
C1192 VTAIL.n507 VSUBS 0.013531f
C1193 VTAIL.n508 VSUBS 0.030204f
C1194 VTAIL.n509 VSUBS 0.030204f
C1195 VTAIL.n510 VSUBS 0.013531f
C1196 VTAIL.n511 VSUBS 0.012779f
C1197 VTAIL.n512 VSUBS 0.023781f
C1198 VTAIL.n513 VSUBS 0.023781f
C1199 VTAIL.n514 VSUBS 0.012779f
C1200 VTAIL.n515 VSUBS 0.013531f
C1201 VTAIL.n516 VSUBS 0.030204f
C1202 VTAIL.n517 VSUBS 0.030204f
C1203 VTAIL.n518 VSUBS 0.013531f
C1204 VTAIL.n519 VSUBS 0.012779f
C1205 VTAIL.n520 VSUBS 0.023781f
C1206 VTAIL.n521 VSUBS 0.023781f
C1207 VTAIL.n522 VSUBS 0.012779f
C1208 VTAIL.n523 VSUBS 0.013531f
C1209 VTAIL.n524 VSUBS 0.030204f
C1210 VTAIL.n525 VSUBS 0.030204f
C1211 VTAIL.n526 VSUBS 0.013531f
C1212 VTAIL.n527 VSUBS 0.012779f
C1213 VTAIL.n528 VSUBS 0.023781f
C1214 VTAIL.n529 VSUBS 0.023781f
C1215 VTAIL.n530 VSUBS 0.012779f
C1216 VTAIL.n531 VSUBS 0.013531f
C1217 VTAIL.n532 VSUBS 0.030204f
C1218 VTAIL.n533 VSUBS 0.030204f
C1219 VTAIL.n534 VSUBS 0.013531f
C1220 VTAIL.n535 VSUBS 0.012779f
C1221 VTAIL.n536 VSUBS 0.023781f
C1222 VTAIL.n537 VSUBS 0.023781f
C1223 VTAIL.n538 VSUBS 0.012779f
C1224 VTAIL.n539 VSUBS 0.013531f
C1225 VTAIL.n540 VSUBS 0.030204f
C1226 VTAIL.n541 VSUBS 0.030204f
C1227 VTAIL.n542 VSUBS 0.013531f
C1228 VTAIL.n543 VSUBS 0.012779f
C1229 VTAIL.n544 VSUBS 0.023781f
C1230 VTAIL.n545 VSUBS 0.023781f
C1231 VTAIL.n546 VSUBS 0.012779f
C1232 VTAIL.n547 VSUBS 0.013155f
C1233 VTAIL.n548 VSUBS 0.013155f
C1234 VTAIL.n549 VSUBS 0.030204f
C1235 VTAIL.n550 VSUBS 0.030204f
C1236 VTAIL.n551 VSUBS 0.013531f
C1237 VTAIL.n552 VSUBS 0.012779f
C1238 VTAIL.n553 VSUBS 0.023781f
C1239 VTAIL.n554 VSUBS 0.023781f
C1240 VTAIL.n555 VSUBS 0.012779f
C1241 VTAIL.n556 VSUBS 0.013531f
C1242 VTAIL.n557 VSUBS 0.030204f
C1243 VTAIL.n558 VSUBS 0.072783f
C1244 VTAIL.n559 VSUBS 0.013531f
C1245 VTAIL.n560 VSUBS 0.012779f
C1246 VTAIL.n561 VSUBS 0.057567f
C1247 VTAIL.n562 VSUBS 0.036665f
C1248 VTAIL.n563 VSUBS 0.108645f
C1249 VTAIL.n564 VSUBS 0.026031f
C1250 VTAIL.n565 VSUBS 0.023781f
C1251 VTAIL.n566 VSUBS 0.012779f
C1252 VTAIL.n567 VSUBS 0.030204f
C1253 VTAIL.n568 VSUBS 0.013531f
C1254 VTAIL.n569 VSUBS 0.023781f
C1255 VTAIL.n570 VSUBS 0.012779f
C1256 VTAIL.n571 VSUBS 0.030204f
C1257 VTAIL.n572 VSUBS 0.013531f
C1258 VTAIL.n573 VSUBS 0.023781f
C1259 VTAIL.n574 VSUBS 0.012779f
C1260 VTAIL.n575 VSUBS 0.030204f
C1261 VTAIL.n576 VSUBS 0.030204f
C1262 VTAIL.n577 VSUBS 0.013531f
C1263 VTAIL.n578 VSUBS 0.023781f
C1264 VTAIL.n579 VSUBS 0.012779f
C1265 VTAIL.n580 VSUBS 0.030204f
C1266 VTAIL.n581 VSUBS 0.013531f
C1267 VTAIL.n582 VSUBS 0.023781f
C1268 VTAIL.n583 VSUBS 0.012779f
C1269 VTAIL.n584 VSUBS 0.030204f
C1270 VTAIL.n585 VSUBS 0.013531f
C1271 VTAIL.n586 VSUBS 0.023781f
C1272 VTAIL.n587 VSUBS 0.012779f
C1273 VTAIL.n588 VSUBS 0.030204f
C1274 VTAIL.n589 VSUBS 0.013531f
C1275 VTAIL.n590 VSUBS 0.023781f
C1276 VTAIL.n591 VSUBS 0.012779f
C1277 VTAIL.n592 VSUBS 0.030204f
C1278 VTAIL.n593 VSUBS 0.013531f
C1279 VTAIL.n594 VSUBS 0.180821f
C1280 VTAIL.t7 VSUBS 0.064773f
C1281 VTAIL.n595 VSUBS 0.022653f
C1282 VTAIL.n596 VSUBS 0.019215f
C1283 VTAIL.n597 VSUBS 0.012779f
C1284 VTAIL.n598 VSUBS 1.72141f
C1285 VTAIL.n599 VSUBS 0.023781f
C1286 VTAIL.n600 VSUBS 0.012779f
C1287 VTAIL.n601 VSUBS 0.013531f
C1288 VTAIL.n602 VSUBS 0.030204f
C1289 VTAIL.n603 VSUBS 0.030204f
C1290 VTAIL.n604 VSUBS 0.013531f
C1291 VTAIL.n605 VSUBS 0.012779f
C1292 VTAIL.n606 VSUBS 0.023781f
C1293 VTAIL.n607 VSUBS 0.023781f
C1294 VTAIL.n608 VSUBS 0.012779f
C1295 VTAIL.n609 VSUBS 0.013531f
C1296 VTAIL.n610 VSUBS 0.030204f
C1297 VTAIL.n611 VSUBS 0.030204f
C1298 VTAIL.n612 VSUBS 0.013531f
C1299 VTAIL.n613 VSUBS 0.012779f
C1300 VTAIL.n614 VSUBS 0.023781f
C1301 VTAIL.n615 VSUBS 0.023781f
C1302 VTAIL.n616 VSUBS 0.012779f
C1303 VTAIL.n617 VSUBS 0.013531f
C1304 VTAIL.n618 VSUBS 0.030204f
C1305 VTAIL.n619 VSUBS 0.030204f
C1306 VTAIL.n620 VSUBS 0.013531f
C1307 VTAIL.n621 VSUBS 0.012779f
C1308 VTAIL.n622 VSUBS 0.023781f
C1309 VTAIL.n623 VSUBS 0.023781f
C1310 VTAIL.n624 VSUBS 0.012779f
C1311 VTAIL.n625 VSUBS 0.013531f
C1312 VTAIL.n626 VSUBS 0.030204f
C1313 VTAIL.n627 VSUBS 0.030204f
C1314 VTAIL.n628 VSUBS 0.013531f
C1315 VTAIL.n629 VSUBS 0.012779f
C1316 VTAIL.n630 VSUBS 0.023781f
C1317 VTAIL.n631 VSUBS 0.023781f
C1318 VTAIL.n632 VSUBS 0.012779f
C1319 VTAIL.n633 VSUBS 0.013531f
C1320 VTAIL.n634 VSUBS 0.030204f
C1321 VTAIL.n635 VSUBS 0.030204f
C1322 VTAIL.n636 VSUBS 0.013531f
C1323 VTAIL.n637 VSUBS 0.012779f
C1324 VTAIL.n638 VSUBS 0.023781f
C1325 VTAIL.n639 VSUBS 0.023781f
C1326 VTAIL.n640 VSUBS 0.012779f
C1327 VTAIL.n641 VSUBS 0.013155f
C1328 VTAIL.n642 VSUBS 0.013155f
C1329 VTAIL.n643 VSUBS 0.030204f
C1330 VTAIL.n644 VSUBS 0.030204f
C1331 VTAIL.n645 VSUBS 0.013531f
C1332 VTAIL.n646 VSUBS 0.012779f
C1333 VTAIL.n647 VSUBS 0.023781f
C1334 VTAIL.n648 VSUBS 0.023781f
C1335 VTAIL.n649 VSUBS 0.012779f
C1336 VTAIL.n650 VSUBS 0.013531f
C1337 VTAIL.n651 VSUBS 0.030204f
C1338 VTAIL.n652 VSUBS 0.072783f
C1339 VTAIL.n653 VSUBS 0.013531f
C1340 VTAIL.n654 VSUBS 0.012779f
C1341 VTAIL.n655 VSUBS 0.057567f
C1342 VTAIL.n656 VSUBS 0.036665f
C1343 VTAIL.n657 VSUBS 1.5616f
C1344 VTAIL.n658 VSUBS 0.026031f
C1345 VTAIL.n659 VSUBS 0.023781f
C1346 VTAIL.n660 VSUBS 0.012779f
C1347 VTAIL.n661 VSUBS 0.030204f
C1348 VTAIL.n662 VSUBS 0.013531f
C1349 VTAIL.n663 VSUBS 0.023781f
C1350 VTAIL.n664 VSUBS 0.012779f
C1351 VTAIL.n665 VSUBS 0.030204f
C1352 VTAIL.n666 VSUBS 0.013531f
C1353 VTAIL.n667 VSUBS 0.023781f
C1354 VTAIL.n668 VSUBS 0.012779f
C1355 VTAIL.n669 VSUBS 0.030204f
C1356 VTAIL.n670 VSUBS 0.013531f
C1357 VTAIL.n671 VSUBS 0.023781f
C1358 VTAIL.n672 VSUBS 0.012779f
C1359 VTAIL.n673 VSUBS 0.030204f
C1360 VTAIL.n674 VSUBS 0.013531f
C1361 VTAIL.n675 VSUBS 0.023781f
C1362 VTAIL.n676 VSUBS 0.012779f
C1363 VTAIL.n677 VSUBS 0.030204f
C1364 VTAIL.n678 VSUBS 0.013531f
C1365 VTAIL.n679 VSUBS 0.023781f
C1366 VTAIL.n680 VSUBS 0.012779f
C1367 VTAIL.n681 VSUBS 0.030204f
C1368 VTAIL.n682 VSUBS 0.013531f
C1369 VTAIL.n683 VSUBS 0.023781f
C1370 VTAIL.n684 VSUBS 0.012779f
C1371 VTAIL.n685 VSUBS 0.030204f
C1372 VTAIL.n686 VSUBS 0.013531f
C1373 VTAIL.n687 VSUBS 0.180821f
C1374 VTAIL.t2 VSUBS 0.064773f
C1375 VTAIL.n688 VSUBS 0.022653f
C1376 VTAIL.n689 VSUBS 0.019215f
C1377 VTAIL.n690 VSUBS 0.012779f
C1378 VTAIL.n691 VSUBS 1.72141f
C1379 VTAIL.n692 VSUBS 0.023781f
C1380 VTAIL.n693 VSUBS 0.012779f
C1381 VTAIL.n694 VSUBS 0.013531f
C1382 VTAIL.n695 VSUBS 0.030204f
C1383 VTAIL.n696 VSUBS 0.030204f
C1384 VTAIL.n697 VSUBS 0.013531f
C1385 VTAIL.n698 VSUBS 0.012779f
C1386 VTAIL.n699 VSUBS 0.023781f
C1387 VTAIL.n700 VSUBS 0.023781f
C1388 VTAIL.n701 VSUBS 0.012779f
C1389 VTAIL.n702 VSUBS 0.013531f
C1390 VTAIL.n703 VSUBS 0.030204f
C1391 VTAIL.n704 VSUBS 0.030204f
C1392 VTAIL.n705 VSUBS 0.013531f
C1393 VTAIL.n706 VSUBS 0.012779f
C1394 VTAIL.n707 VSUBS 0.023781f
C1395 VTAIL.n708 VSUBS 0.023781f
C1396 VTAIL.n709 VSUBS 0.012779f
C1397 VTAIL.n710 VSUBS 0.013531f
C1398 VTAIL.n711 VSUBS 0.030204f
C1399 VTAIL.n712 VSUBS 0.030204f
C1400 VTAIL.n713 VSUBS 0.013531f
C1401 VTAIL.n714 VSUBS 0.012779f
C1402 VTAIL.n715 VSUBS 0.023781f
C1403 VTAIL.n716 VSUBS 0.023781f
C1404 VTAIL.n717 VSUBS 0.012779f
C1405 VTAIL.n718 VSUBS 0.013531f
C1406 VTAIL.n719 VSUBS 0.030204f
C1407 VTAIL.n720 VSUBS 0.030204f
C1408 VTAIL.n721 VSUBS 0.013531f
C1409 VTAIL.n722 VSUBS 0.012779f
C1410 VTAIL.n723 VSUBS 0.023781f
C1411 VTAIL.n724 VSUBS 0.023781f
C1412 VTAIL.n725 VSUBS 0.012779f
C1413 VTAIL.n726 VSUBS 0.013531f
C1414 VTAIL.n727 VSUBS 0.030204f
C1415 VTAIL.n728 VSUBS 0.030204f
C1416 VTAIL.n729 VSUBS 0.030204f
C1417 VTAIL.n730 VSUBS 0.013531f
C1418 VTAIL.n731 VSUBS 0.012779f
C1419 VTAIL.n732 VSUBS 0.023781f
C1420 VTAIL.n733 VSUBS 0.023781f
C1421 VTAIL.n734 VSUBS 0.012779f
C1422 VTAIL.n735 VSUBS 0.013155f
C1423 VTAIL.n736 VSUBS 0.013155f
C1424 VTAIL.n737 VSUBS 0.030204f
C1425 VTAIL.n738 VSUBS 0.030204f
C1426 VTAIL.n739 VSUBS 0.013531f
C1427 VTAIL.n740 VSUBS 0.012779f
C1428 VTAIL.n741 VSUBS 0.023781f
C1429 VTAIL.n742 VSUBS 0.023781f
C1430 VTAIL.n743 VSUBS 0.012779f
C1431 VTAIL.n744 VSUBS 0.013531f
C1432 VTAIL.n745 VSUBS 0.030204f
C1433 VTAIL.n746 VSUBS 0.072783f
C1434 VTAIL.n747 VSUBS 0.013531f
C1435 VTAIL.n748 VSUBS 0.012779f
C1436 VTAIL.n749 VSUBS 0.057567f
C1437 VTAIL.n750 VSUBS 0.036665f
C1438 VTAIL.n751 VSUBS 1.53171f
C1439 VP.t0 VSUBS 1.44903f
C1440 VP.t3 VSUBS 1.44904f
C1441 VP.n0 VSUBS 2.24352f
C1442 VP.n1 VSUBS 4.8995f
C1443 VP.t1 VSUBS 1.43783f
C1444 VP.n2 VSUBS 0.55309f
C1445 VP.t2 VSUBS 1.43783f
C1446 VP.n3 VSUBS 0.55309f
C1447 VP.n4 VSUBS 0.052875f
.ends

