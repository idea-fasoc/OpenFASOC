* NGSPICE file created from diff_pair_sample_0908.ext - technology: sky130A

.subckt diff_pair_sample_0908 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=0 ps=0 w=17.17 l=0.77
X1 VDD2.t5 VN.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=6.6963 ps=35.12 w=17.17 l=0.77
X2 VDD2.t4 VN.t1 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=2.83305 ps=17.5 w=17.17 l=0.77
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=0 ps=0 w=17.17 l=0.77
X4 VDD1.t5 VP.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=6.6963 ps=35.12 w=17.17 l=0.77
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=0 ps=0 w=17.17 l=0.77
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=0 ps=0 w=17.17 l=0.77
X7 VDD2.t3 VN.t2 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=2.83305 ps=17.5 w=17.17 l=0.77
X8 VTAIL.t8 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=2.83305 ps=17.5 w=17.17 l=0.77
X9 VDD1.t4 VP.t1 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=2.83305 ps=17.5 w=17.17 l=0.77
X10 VDD2.t1 VN.t4 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=6.6963 ps=35.12 w=17.17 l=0.77
X11 VTAIL.t2 VP.t2 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=2.83305 ps=17.5 w=17.17 l=0.77
X12 VDD1.t2 VP.t3 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=6.6963 ps=35.12 w=17.17 l=0.77
X13 VTAIL.t3 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=2.83305 ps=17.5 w=17.17 l=0.77
X14 VTAIL.t10 VN.t5 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83305 pd=17.5 as=2.83305 ps=17.5 w=17.17 l=0.77
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6963 pd=35.12 as=2.83305 ps=17.5 w=17.17 l=0.77
R0 B.n458 B.t6 739.582
R1 B.n455 B.t14 739.582
R2 B.n107 B.t17 739.582
R3 B.n104 B.t10 739.582
R4 B.n797 B.n796 585
R5 B.n798 B.n797 585
R6 B.n352 B.n103 585
R7 B.n351 B.n350 585
R8 B.n349 B.n348 585
R9 B.n347 B.n346 585
R10 B.n345 B.n344 585
R11 B.n343 B.n342 585
R12 B.n341 B.n340 585
R13 B.n339 B.n338 585
R14 B.n337 B.n336 585
R15 B.n335 B.n334 585
R16 B.n333 B.n332 585
R17 B.n331 B.n330 585
R18 B.n329 B.n328 585
R19 B.n327 B.n326 585
R20 B.n325 B.n324 585
R21 B.n323 B.n322 585
R22 B.n321 B.n320 585
R23 B.n319 B.n318 585
R24 B.n317 B.n316 585
R25 B.n315 B.n314 585
R26 B.n313 B.n312 585
R27 B.n311 B.n310 585
R28 B.n309 B.n308 585
R29 B.n307 B.n306 585
R30 B.n305 B.n304 585
R31 B.n303 B.n302 585
R32 B.n301 B.n300 585
R33 B.n299 B.n298 585
R34 B.n297 B.n296 585
R35 B.n295 B.n294 585
R36 B.n293 B.n292 585
R37 B.n291 B.n290 585
R38 B.n289 B.n288 585
R39 B.n287 B.n286 585
R40 B.n285 B.n284 585
R41 B.n283 B.n282 585
R42 B.n281 B.n280 585
R43 B.n279 B.n278 585
R44 B.n277 B.n276 585
R45 B.n275 B.n274 585
R46 B.n273 B.n272 585
R47 B.n271 B.n270 585
R48 B.n269 B.n268 585
R49 B.n267 B.n266 585
R50 B.n265 B.n264 585
R51 B.n263 B.n262 585
R52 B.n261 B.n260 585
R53 B.n259 B.n258 585
R54 B.n257 B.n256 585
R55 B.n255 B.n254 585
R56 B.n253 B.n252 585
R57 B.n251 B.n250 585
R58 B.n249 B.n248 585
R59 B.n247 B.n246 585
R60 B.n245 B.n244 585
R61 B.n243 B.n242 585
R62 B.n241 B.n240 585
R63 B.n239 B.n238 585
R64 B.n237 B.n236 585
R65 B.n235 B.n234 585
R66 B.n233 B.n232 585
R67 B.n231 B.n230 585
R68 B.n229 B.n228 585
R69 B.n227 B.n226 585
R70 B.n225 B.n224 585
R71 B.n222 B.n221 585
R72 B.n220 B.n219 585
R73 B.n218 B.n217 585
R74 B.n216 B.n215 585
R75 B.n214 B.n213 585
R76 B.n212 B.n211 585
R77 B.n210 B.n209 585
R78 B.n208 B.n207 585
R79 B.n206 B.n205 585
R80 B.n204 B.n203 585
R81 B.n202 B.n201 585
R82 B.n200 B.n199 585
R83 B.n198 B.n197 585
R84 B.n196 B.n195 585
R85 B.n194 B.n193 585
R86 B.n192 B.n191 585
R87 B.n190 B.n189 585
R88 B.n188 B.n187 585
R89 B.n186 B.n185 585
R90 B.n184 B.n183 585
R91 B.n182 B.n181 585
R92 B.n180 B.n179 585
R93 B.n178 B.n177 585
R94 B.n176 B.n175 585
R95 B.n174 B.n173 585
R96 B.n172 B.n171 585
R97 B.n170 B.n169 585
R98 B.n168 B.n167 585
R99 B.n166 B.n165 585
R100 B.n164 B.n163 585
R101 B.n162 B.n161 585
R102 B.n160 B.n159 585
R103 B.n158 B.n157 585
R104 B.n156 B.n155 585
R105 B.n154 B.n153 585
R106 B.n152 B.n151 585
R107 B.n150 B.n149 585
R108 B.n148 B.n147 585
R109 B.n146 B.n145 585
R110 B.n144 B.n143 585
R111 B.n142 B.n141 585
R112 B.n140 B.n139 585
R113 B.n138 B.n137 585
R114 B.n136 B.n135 585
R115 B.n134 B.n133 585
R116 B.n132 B.n131 585
R117 B.n130 B.n129 585
R118 B.n128 B.n127 585
R119 B.n126 B.n125 585
R120 B.n124 B.n123 585
R121 B.n122 B.n121 585
R122 B.n120 B.n119 585
R123 B.n118 B.n117 585
R124 B.n116 B.n115 585
R125 B.n114 B.n113 585
R126 B.n112 B.n111 585
R127 B.n110 B.n109 585
R128 B.n795 B.n41 585
R129 B.n799 B.n41 585
R130 B.n794 B.n40 585
R131 B.n800 B.n40 585
R132 B.n793 B.n792 585
R133 B.n792 B.n36 585
R134 B.n791 B.n35 585
R135 B.n806 B.n35 585
R136 B.n790 B.n34 585
R137 B.n807 B.n34 585
R138 B.n789 B.n33 585
R139 B.n808 B.n33 585
R140 B.n788 B.n787 585
R141 B.n787 B.n29 585
R142 B.n786 B.n28 585
R143 B.n814 B.n28 585
R144 B.n785 B.n27 585
R145 B.n815 B.n27 585
R146 B.n784 B.n26 585
R147 B.n816 B.n26 585
R148 B.n783 B.n782 585
R149 B.n782 B.n22 585
R150 B.n781 B.n21 585
R151 B.n822 B.n21 585
R152 B.n780 B.n20 585
R153 B.n823 B.n20 585
R154 B.n779 B.n19 585
R155 B.n824 B.n19 585
R156 B.n778 B.n777 585
R157 B.n777 B.n18 585
R158 B.n776 B.n14 585
R159 B.n830 B.n14 585
R160 B.n775 B.n13 585
R161 B.n831 B.n13 585
R162 B.n774 B.n12 585
R163 B.n832 B.n12 585
R164 B.n773 B.n772 585
R165 B.n772 B.n8 585
R166 B.n771 B.n7 585
R167 B.n838 B.n7 585
R168 B.n770 B.n6 585
R169 B.n839 B.n6 585
R170 B.n769 B.n5 585
R171 B.n840 B.n5 585
R172 B.n768 B.n767 585
R173 B.n767 B.n4 585
R174 B.n766 B.n353 585
R175 B.n766 B.n765 585
R176 B.n756 B.n354 585
R177 B.n355 B.n354 585
R178 B.n758 B.n757 585
R179 B.n759 B.n758 585
R180 B.n755 B.n360 585
R181 B.n360 B.n359 585
R182 B.n754 B.n753 585
R183 B.n753 B.n752 585
R184 B.n362 B.n361 585
R185 B.n745 B.n362 585
R186 B.n744 B.n743 585
R187 B.n746 B.n744 585
R188 B.n742 B.n367 585
R189 B.n367 B.n366 585
R190 B.n741 B.n740 585
R191 B.n740 B.n739 585
R192 B.n369 B.n368 585
R193 B.n370 B.n369 585
R194 B.n732 B.n731 585
R195 B.n733 B.n732 585
R196 B.n730 B.n375 585
R197 B.n375 B.n374 585
R198 B.n729 B.n728 585
R199 B.n728 B.n727 585
R200 B.n377 B.n376 585
R201 B.n378 B.n377 585
R202 B.n720 B.n719 585
R203 B.n721 B.n720 585
R204 B.n718 B.n382 585
R205 B.n386 B.n382 585
R206 B.n717 B.n716 585
R207 B.n716 B.n715 585
R208 B.n384 B.n383 585
R209 B.n385 B.n384 585
R210 B.n708 B.n707 585
R211 B.n709 B.n708 585
R212 B.n706 B.n391 585
R213 B.n391 B.n390 585
R214 B.n700 B.n699 585
R215 B.n698 B.n454 585
R216 B.n697 B.n453 585
R217 B.n702 B.n453 585
R218 B.n696 B.n695 585
R219 B.n694 B.n693 585
R220 B.n692 B.n691 585
R221 B.n690 B.n689 585
R222 B.n688 B.n687 585
R223 B.n686 B.n685 585
R224 B.n684 B.n683 585
R225 B.n682 B.n681 585
R226 B.n680 B.n679 585
R227 B.n678 B.n677 585
R228 B.n676 B.n675 585
R229 B.n674 B.n673 585
R230 B.n672 B.n671 585
R231 B.n670 B.n669 585
R232 B.n668 B.n667 585
R233 B.n666 B.n665 585
R234 B.n664 B.n663 585
R235 B.n662 B.n661 585
R236 B.n660 B.n659 585
R237 B.n658 B.n657 585
R238 B.n656 B.n655 585
R239 B.n654 B.n653 585
R240 B.n652 B.n651 585
R241 B.n650 B.n649 585
R242 B.n648 B.n647 585
R243 B.n646 B.n645 585
R244 B.n644 B.n643 585
R245 B.n642 B.n641 585
R246 B.n640 B.n639 585
R247 B.n638 B.n637 585
R248 B.n636 B.n635 585
R249 B.n634 B.n633 585
R250 B.n632 B.n631 585
R251 B.n630 B.n629 585
R252 B.n628 B.n627 585
R253 B.n626 B.n625 585
R254 B.n624 B.n623 585
R255 B.n622 B.n621 585
R256 B.n620 B.n619 585
R257 B.n618 B.n617 585
R258 B.n616 B.n615 585
R259 B.n614 B.n613 585
R260 B.n612 B.n611 585
R261 B.n610 B.n609 585
R262 B.n608 B.n607 585
R263 B.n606 B.n605 585
R264 B.n604 B.n603 585
R265 B.n602 B.n601 585
R266 B.n600 B.n599 585
R267 B.n598 B.n597 585
R268 B.n596 B.n595 585
R269 B.n594 B.n593 585
R270 B.n592 B.n591 585
R271 B.n590 B.n589 585
R272 B.n588 B.n587 585
R273 B.n586 B.n585 585
R274 B.n584 B.n583 585
R275 B.n582 B.n581 585
R276 B.n580 B.n579 585
R277 B.n578 B.n577 585
R278 B.n576 B.n575 585
R279 B.n574 B.n573 585
R280 B.n572 B.n571 585
R281 B.n569 B.n568 585
R282 B.n567 B.n566 585
R283 B.n565 B.n564 585
R284 B.n563 B.n562 585
R285 B.n561 B.n560 585
R286 B.n559 B.n558 585
R287 B.n557 B.n556 585
R288 B.n555 B.n554 585
R289 B.n553 B.n552 585
R290 B.n551 B.n550 585
R291 B.n549 B.n548 585
R292 B.n547 B.n546 585
R293 B.n545 B.n544 585
R294 B.n543 B.n542 585
R295 B.n541 B.n540 585
R296 B.n539 B.n538 585
R297 B.n537 B.n536 585
R298 B.n535 B.n534 585
R299 B.n533 B.n532 585
R300 B.n531 B.n530 585
R301 B.n529 B.n528 585
R302 B.n527 B.n526 585
R303 B.n525 B.n524 585
R304 B.n523 B.n522 585
R305 B.n521 B.n520 585
R306 B.n519 B.n518 585
R307 B.n517 B.n516 585
R308 B.n515 B.n514 585
R309 B.n513 B.n512 585
R310 B.n511 B.n510 585
R311 B.n509 B.n508 585
R312 B.n507 B.n506 585
R313 B.n505 B.n504 585
R314 B.n503 B.n502 585
R315 B.n501 B.n500 585
R316 B.n499 B.n498 585
R317 B.n497 B.n496 585
R318 B.n495 B.n494 585
R319 B.n493 B.n492 585
R320 B.n491 B.n490 585
R321 B.n489 B.n488 585
R322 B.n487 B.n486 585
R323 B.n485 B.n484 585
R324 B.n483 B.n482 585
R325 B.n481 B.n480 585
R326 B.n479 B.n478 585
R327 B.n477 B.n476 585
R328 B.n475 B.n474 585
R329 B.n473 B.n472 585
R330 B.n471 B.n470 585
R331 B.n469 B.n468 585
R332 B.n467 B.n466 585
R333 B.n465 B.n464 585
R334 B.n463 B.n462 585
R335 B.n461 B.n460 585
R336 B.n393 B.n392 585
R337 B.n705 B.n704 585
R338 B.n389 B.n388 585
R339 B.n390 B.n389 585
R340 B.n711 B.n710 585
R341 B.n710 B.n709 585
R342 B.n712 B.n387 585
R343 B.n387 B.n385 585
R344 B.n714 B.n713 585
R345 B.n715 B.n714 585
R346 B.n381 B.n380 585
R347 B.n386 B.n381 585
R348 B.n723 B.n722 585
R349 B.n722 B.n721 585
R350 B.n724 B.n379 585
R351 B.n379 B.n378 585
R352 B.n726 B.n725 585
R353 B.n727 B.n726 585
R354 B.n373 B.n372 585
R355 B.n374 B.n373 585
R356 B.n735 B.n734 585
R357 B.n734 B.n733 585
R358 B.n736 B.n371 585
R359 B.n371 B.n370 585
R360 B.n738 B.n737 585
R361 B.n739 B.n738 585
R362 B.n365 B.n364 585
R363 B.n366 B.n365 585
R364 B.n748 B.n747 585
R365 B.n747 B.n746 585
R366 B.n749 B.n363 585
R367 B.n745 B.n363 585
R368 B.n751 B.n750 585
R369 B.n752 B.n751 585
R370 B.n358 B.n357 585
R371 B.n359 B.n358 585
R372 B.n761 B.n760 585
R373 B.n760 B.n759 585
R374 B.n762 B.n356 585
R375 B.n356 B.n355 585
R376 B.n764 B.n763 585
R377 B.n765 B.n764 585
R378 B.n2 B.n0 585
R379 B.n4 B.n2 585
R380 B.n3 B.n1 585
R381 B.n839 B.n3 585
R382 B.n837 B.n836 585
R383 B.n838 B.n837 585
R384 B.n835 B.n9 585
R385 B.n9 B.n8 585
R386 B.n834 B.n833 585
R387 B.n833 B.n832 585
R388 B.n11 B.n10 585
R389 B.n831 B.n11 585
R390 B.n829 B.n828 585
R391 B.n830 B.n829 585
R392 B.n827 B.n15 585
R393 B.n18 B.n15 585
R394 B.n826 B.n825 585
R395 B.n825 B.n824 585
R396 B.n17 B.n16 585
R397 B.n823 B.n17 585
R398 B.n821 B.n820 585
R399 B.n822 B.n821 585
R400 B.n819 B.n23 585
R401 B.n23 B.n22 585
R402 B.n818 B.n817 585
R403 B.n817 B.n816 585
R404 B.n25 B.n24 585
R405 B.n815 B.n25 585
R406 B.n813 B.n812 585
R407 B.n814 B.n813 585
R408 B.n811 B.n30 585
R409 B.n30 B.n29 585
R410 B.n810 B.n809 585
R411 B.n809 B.n808 585
R412 B.n32 B.n31 585
R413 B.n807 B.n32 585
R414 B.n805 B.n804 585
R415 B.n806 B.n805 585
R416 B.n803 B.n37 585
R417 B.n37 B.n36 585
R418 B.n802 B.n801 585
R419 B.n801 B.n800 585
R420 B.n39 B.n38 585
R421 B.n799 B.n39 585
R422 B.n842 B.n841 585
R423 B.n841 B.n840 585
R424 B.n700 B.n389 526.135
R425 B.n109 B.n39 526.135
R426 B.n704 B.n391 526.135
R427 B.n797 B.n41 526.135
R428 B.n798 B.n102 256.663
R429 B.n798 B.n101 256.663
R430 B.n798 B.n100 256.663
R431 B.n798 B.n99 256.663
R432 B.n798 B.n98 256.663
R433 B.n798 B.n97 256.663
R434 B.n798 B.n96 256.663
R435 B.n798 B.n95 256.663
R436 B.n798 B.n94 256.663
R437 B.n798 B.n93 256.663
R438 B.n798 B.n92 256.663
R439 B.n798 B.n91 256.663
R440 B.n798 B.n90 256.663
R441 B.n798 B.n89 256.663
R442 B.n798 B.n88 256.663
R443 B.n798 B.n87 256.663
R444 B.n798 B.n86 256.663
R445 B.n798 B.n85 256.663
R446 B.n798 B.n84 256.663
R447 B.n798 B.n83 256.663
R448 B.n798 B.n82 256.663
R449 B.n798 B.n81 256.663
R450 B.n798 B.n80 256.663
R451 B.n798 B.n79 256.663
R452 B.n798 B.n78 256.663
R453 B.n798 B.n77 256.663
R454 B.n798 B.n76 256.663
R455 B.n798 B.n75 256.663
R456 B.n798 B.n74 256.663
R457 B.n798 B.n73 256.663
R458 B.n798 B.n72 256.663
R459 B.n798 B.n71 256.663
R460 B.n798 B.n70 256.663
R461 B.n798 B.n69 256.663
R462 B.n798 B.n68 256.663
R463 B.n798 B.n67 256.663
R464 B.n798 B.n66 256.663
R465 B.n798 B.n65 256.663
R466 B.n798 B.n64 256.663
R467 B.n798 B.n63 256.663
R468 B.n798 B.n62 256.663
R469 B.n798 B.n61 256.663
R470 B.n798 B.n60 256.663
R471 B.n798 B.n59 256.663
R472 B.n798 B.n58 256.663
R473 B.n798 B.n57 256.663
R474 B.n798 B.n56 256.663
R475 B.n798 B.n55 256.663
R476 B.n798 B.n54 256.663
R477 B.n798 B.n53 256.663
R478 B.n798 B.n52 256.663
R479 B.n798 B.n51 256.663
R480 B.n798 B.n50 256.663
R481 B.n798 B.n49 256.663
R482 B.n798 B.n48 256.663
R483 B.n798 B.n47 256.663
R484 B.n798 B.n46 256.663
R485 B.n798 B.n45 256.663
R486 B.n798 B.n44 256.663
R487 B.n798 B.n43 256.663
R488 B.n798 B.n42 256.663
R489 B.n702 B.n701 256.663
R490 B.n702 B.n394 256.663
R491 B.n702 B.n395 256.663
R492 B.n702 B.n396 256.663
R493 B.n702 B.n397 256.663
R494 B.n702 B.n398 256.663
R495 B.n702 B.n399 256.663
R496 B.n702 B.n400 256.663
R497 B.n702 B.n401 256.663
R498 B.n702 B.n402 256.663
R499 B.n702 B.n403 256.663
R500 B.n702 B.n404 256.663
R501 B.n702 B.n405 256.663
R502 B.n702 B.n406 256.663
R503 B.n702 B.n407 256.663
R504 B.n702 B.n408 256.663
R505 B.n702 B.n409 256.663
R506 B.n702 B.n410 256.663
R507 B.n702 B.n411 256.663
R508 B.n702 B.n412 256.663
R509 B.n702 B.n413 256.663
R510 B.n702 B.n414 256.663
R511 B.n702 B.n415 256.663
R512 B.n702 B.n416 256.663
R513 B.n702 B.n417 256.663
R514 B.n702 B.n418 256.663
R515 B.n702 B.n419 256.663
R516 B.n702 B.n420 256.663
R517 B.n702 B.n421 256.663
R518 B.n702 B.n422 256.663
R519 B.n702 B.n423 256.663
R520 B.n702 B.n424 256.663
R521 B.n702 B.n425 256.663
R522 B.n702 B.n426 256.663
R523 B.n702 B.n427 256.663
R524 B.n702 B.n428 256.663
R525 B.n702 B.n429 256.663
R526 B.n702 B.n430 256.663
R527 B.n702 B.n431 256.663
R528 B.n702 B.n432 256.663
R529 B.n702 B.n433 256.663
R530 B.n702 B.n434 256.663
R531 B.n702 B.n435 256.663
R532 B.n702 B.n436 256.663
R533 B.n702 B.n437 256.663
R534 B.n702 B.n438 256.663
R535 B.n702 B.n439 256.663
R536 B.n702 B.n440 256.663
R537 B.n702 B.n441 256.663
R538 B.n702 B.n442 256.663
R539 B.n702 B.n443 256.663
R540 B.n702 B.n444 256.663
R541 B.n702 B.n445 256.663
R542 B.n702 B.n446 256.663
R543 B.n702 B.n447 256.663
R544 B.n702 B.n448 256.663
R545 B.n702 B.n449 256.663
R546 B.n702 B.n450 256.663
R547 B.n702 B.n451 256.663
R548 B.n702 B.n452 256.663
R549 B.n703 B.n702 256.663
R550 B.n710 B.n389 163.367
R551 B.n710 B.n387 163.367
R552 B.n714 B.n387 163.367
R553 B.n714 B.n381 163.367
R554 B.n722 B.n381 163.367
R555 B.n722 B.n379 163.367
R556 B.n726 B.n379 163.367
R557 B.n726 B.n373 163.367
R558 B.n734 B.n373 163.367
R559 B.n734 B.n371 163.367
R560 B.n738 B.n371 163.367
R561 B.n738 B.n365 163.367
R562 B.n747 B.n365 163.367
R563 B.n747 B.n363 163.367
R564 B.n751 B.n363 163.367
R565 B.n751 B.n358 163.367
R566 B.n760 B.n358 163.367
R567 B.n760 B.n356 163.367
R568 B.n764 B.n356 163.367
R569 B.n764 B.n2 163.367
R570 B.n841 B.n2 163.367
R571 B.n841 B.n3 163.367
R572 B.n837 B.n3 163.367
R573 B.n837 B.n9 163.367
R574 B.n833 B.n9 163.367
R575 B.n833 B.n11 163.367
R576 B.n829 B.n11 163.367
R577 B.n829 B.n15 163.367
R578 B.n825 B.n15 163.367
R579 B.n825 B.n17 163.367
R580 B.n821 B.n17 163.367
R581 B.n821 B.n23 163.367
R582 B.n817 B.n23 163.367
R583 B.n817 B.n25 163.367
R584 B.n813 B.n25 163.367
R585 B.n813 B.n30 163.367
R586 B.n809 B.n30 163.367
R587 B.n809 B.n32 163.367
R588 B.n805 B.n32 163.367
R589 B.n805 B.n37 163.367
R590 B.n801 B.n37 163.367
R591 B.n801 B.n39 163.367
R592 B.n454 B.n453 163.367
R593 B.n695 B.n453 163.367
R594 B.n693 B.n692 163.367
R595 B.n689 B.n688 163.367
R596 B.n685 B.n684 163.367
R597 B.n681 B.n680 163.367
R598 B.n677 B.n676 163.367
R599 B.n673 B.n672 163.367
R600 B.n669 B.n668 163.367
R601 B.n665 B.n664 163.367
R602 B.n661 B.n660 163.367
R603 B.n657 B.n656 163.367
R604 B.n653 B.n652 163.367
R605 B.n649 B.n648 163.367
R606 B.n645 B.n644 163.367
R607 B.n641 B.n640 163.367
R608 B.n637 B.n636 163.367
R609 B.n633 B.n632 163.367
R610 B.n629 B.n628 163.367
R611 B.n625 B.n624 163.367
R612 B.n621 B.n620 163.367
R613 B.n617 B.n616 163.367
R614 B.n613 B.n612 163.367
R615 B.n609 B.n608 163.367
R616 B.n605 B.n604 163.367
R617 B.n601 B.n600 163.367
R618 B.n597 B.n596 163.367
R619 B.n593 B.n592 163.367
R620 B.n589 B.n588 163.367
R621 B.n585 B.n584 163.367
R622 B.n581 B.n580 163.367
R623 B.n577 B.n576 163.367
R624 B.n573 B.n572 163.367
R625 B.n568 B.n567 163.367
R626 B.n564 B.n563 163.367
R627 B.n560 B.n559 163.367
R628 B.n556 B.n555 163.367
R629 B.n552 B.n551 163.367
R630 B.n548 B.n547 163.367
R631 B.n544 B.n543 163.367
R632 B.n540 B.n539 163.367
R633 B.n536 B.n535 163.367
R634 B.n532 B.n531 163.367
R635 B.n528 B.n527 163.367
R636 B.n524 B.n523 163.367
R637 B.n520 B.n519 163.367
R638 B.n516 B.n515 163.367
R639 B.n512 B.n511 163.367
R640 B.n508 B.n507 163.367
R641 B.n504 B.n503 163.367
R642 B.n500 B.n499 163.367
R643 B.n496 B.n495 163.367
R644 B.n492 B.n491 163.367
R645 B.n488 B.n487 163.367
R646 B.n484 B.n483 163.367
R647 B.n480 B.n479 163.367
R648 B.n476 B.n475 163.367
R649 B.n472 B.n471 163.367
R650 B.n468 B.n467 163.367
R651 B.n464 B.n463 163.367
R652 B.n460 B.n393 163.367
R653 B.n708 B.n391 163.367
R654 B.n708 B.n384 163.367
R655 B.n716 B.n384 163.367
R656 B.n716 B.n382 163.367
R657 B.n720 B.n382 163.367
R658 B.n720 B.n377 163.367
R659 B.n728 B.n377 163.367
R660 B.n728 B.n375 163.367
R661 B.n732 B.n375 163.367
R662 B.n732 B.n369 163.367
R663 B.n740 B.n369 163.367
R664 B.n740 B.n367 163.367
R665 B.n744 B.n367 163.367
R666 B.n744 B.n362 163.367
R667 B.n753 B.n362 163.367
R668 B.n753 B.n360 163.367
R669 B.n758 B.n360 163.367
R670 B.n758 B.n354 163.367
R671 B.n766 B.n354 163.367
R672 B.n767 B.n766 163.367
R673 B.n767 B.n5 163.367
R674 B.n6 B.n5 163.367
R675 B.n7 B.n6 163.367
R676 B.n772 B.n7 163.367
R677 B.n772 B.n12 163.367
R678 B.n13 B.n12 163.367
R679 B.n14 B.n13 163.367
R680 B.n777 B.n14 163.367
R681 B.n777 B.n19 163.367
R682 B.n20 B.n19 163.367
R683 B.n21 B.n20 163.367
R684 B.n782 B.n21 163.367
R685 B.n782 B.n26 163.367
R686 B.n27 B.n26 163.367
R687 B.n28 B.n27 163.367
R688 B.n787 B.n28 163.367
R689 B.n787 B.n33 163.367
R690 B.n34 B.n33 163.367
R691 B.n35 B.n34 163.367
R692 B.n792 B.n35 163.367
R693 B.n792 B.n40 163.367
R694 B.n41 B.n40 163.367
R695 B.n113 B.n112 163.367
R696 B.n117 B.n116 163.367
R697 B.n121 B.n120 163.367
R698 B.n125 B.n124 163.367
R699 B.n129 B.n128 163.367
R700 B.n133 B.n132 163.367
R701 B.n137 B.n136 163.367
R702 B.n141 B.n140 163.367
R703 B.n145 B.n144 163.367
R704 B.n149 B.n148 163.367
R705 B.n153 B.n152 163.367
R706 B.n157 B.n156 163.367
R707 B.n161 B.n160 163.367
R708 B.n165 B.n164 163.367
R709 B.n169 B.n168 163.367
R710 B.n173 B.n172 163.367
R711 B.n177 B.n176 163.367
R712 B.n181 B.n180 163.367
R713 B.n185 B.n184 163.367
R714 B.n189 B.n188 163.367
R715 B.n193 B.n192 163.367
R716 B.n197 B.n196 163.367
R717 B.n201 B.n200 163.367
R718 B.n205 B.n204 163.367
R719 B.n209 B.n208 163.367
R720 B.n213 B.n212 163.367
R721 B.n217 B.n216 163.367
R722 B.n221 B.n220 163.367
R723 B.n226 B.n225 163.367
R724 B.n230 B.n229 163.367
R725 B.n234 B.n233 163.367
R726 B.n238 B.n237 163.367
R727 B.n242 B.n241 163.367
R728 B.n246 B.n245 163.367
R729 B.n250 B.n249 163.367
R730 B.n254 B.n253 163.367
R731 B.n258 B.n257 163.367
R732 B.n262 B.n261 163.367
R733 B.n266 B.n265 163.367
R734 B.n270 B.n269 163.367
R735 B.n274 B.n273 163.367
R736 B.n278 B.n277 163.367
R737 B.n282 B.n281 163.367
R738 B.n286 B.n285 163.367
R739 B.n290 B.n289 163.367
R740 B.n294 B.n293 163.367
R741 B.n298 B.n297 163.367
R742 B.n302 B.n301 163.367
R743 B.n306 B.n305 163.367
R744 B.n310 B.n309 163.367
R745 B.n314 B.n313 163.367
R746 B.n318 B.n317 163.367
R747 B.n322 B.n321 163.367
R748 B.n326 B.n325 163.367
R749 B.n330 B.n329 163.367
R750 B.n334 B.n333 163.367
R751 B.n338 B.n337 163.367
R752 B.n342 B.n341 163.367
R753 B.n346 B.n345 163.367
R754 B.n350 B.n349 163.367
R755 B.n797 B.n103 163.367
R756 B.n458 B.t9 91.9309
R757 B.n104 B.t12 91.9309
R758 B.n455 B.t16 91.9081
R759 B.n107 B.t18 91.9081
R760 B.n701 B.n700 71.676
R761 B.n695 B.n394 71.676
R762 B.n692 B.n395 71.676
R763 B.n688 B.n396 71.676
R764 B.n684 B.n397 71.676
R765 B.n680 B.n398 71.676
R766 B.n676 B.n399 71.676
R767 B.n672 B.n400 71.676
R768 B.n668 B.n401 71.676
R769 B.n664 B.n402 71.676
R770 B.n660 B.n403 71.676
R771 B.n656 B.n404 71.676
R772 B.n652 B.n405 71.676
R773 B.n648 B.n406 71.676
R774 B.n644 B.n407 71.676
R775 B.n640 B.n408 71.676
R776 B.n636 B.n409 71.676
R777 B.n632 B.n410 71.676
R778 B.n628 B.n411 71.676
R779 B.n624 B.n412 71.676
R780 B.n620 B.n413 71.676
R781 B.n616 B.n414 71.676
R782 B.n612 B.n415 71.676
R783 B.n608 B.n416 71.676
R784 B.n604 B.n417 71.676
R785 B.n600 B.n418 71.676
R786 B.n596 B.n419 71.676
R787 B.n592 B.n420 71.676
R788 B.n588 B.n421 71.676
R789 B.n584 B.n422 71.676
R790 B.n580 B.n423 71.676
R791 B.n576 B.n424 71.676
R792 B.n572 B.n425 71.676
R793 B.n567 B.n426 71.676
R794 B.n563 B.n427 71.676
R795 B.n559 B.n428 71.676
R796 B.n555 B.n429 71.676
R797 B.n551 B.n430 71.676
R798 B.n547 B.n431 71.676
R799 B.n543 B.n432 71.676
R800 B.n539 B.n433 71.676
R801 B.n535 B.n434 71.676
R802 B.n531 B.n435 71.676
R803 B.n527 B.n436 71.676
R804 B.n523 B.n437 71.676
R805 B.n519 B.n438 71.676
R806 B.n515 B.n439 71.676
R807 B.n511 B.n440 71.676
R808 B.n507 B.n441 71.676
R809 B.n503 B.n442 71.676
R810 B.n499 B.n443 71.676
R811 B.n495 B.n444 71.676
R812 B.n491 B.n445 71.676
R813 B.n487 B.n446 71.676
R814 B.n483 B.n447 71.676
R815 B.n479 B.n448 71.676
R816 B.n475 B.n449 71.676
R817 B.n471 B.n450 71.676
R818 B.n467 B.n451 71.676
R819 B.n463 B.n452 71.676
R820 B.n703 B.n393 71.676
R821 B.n109 B.n42 71.676
R822 B.n113 B.n43 71.676
R823 B.n117 B.n44 71.676
R824 B.n121 B.n45 71.676
R825 B.n125 B.n46 71.676
R826 B.n129 B.n47 71.676
R827 B.n133 B.n48 71.676
R828 B.n137 B.n49 71.676
R829 B.n141 B.n50 71.676
R830 B.n145 B.n51 71.676
R831 B.n149 B.n52 71.676
R832 B.n153 B.n53 71.676
R833 B.n157 B.n54 71.676
R834 B.n161 B.n55 71.676
R835 B.n165 B.n56 71.676
R836 B.n169 B.n57 71.676
R837 B.n173 B.n58 71.676
R838 B.n177 B.n59 71.676
R839 B.n181 B.n60 71.676
R840 B.n185 B.n61 71.676
R841 B.n189 B.n62 71.676
R842 B.n193 B.n63 71.676
R843 B.n197 B.n64 71.676
R844 B.n201 B.n65 71.676
R845 B.n205 B.n66 71.676
R846 B.n209 B.n67 71.676
R847 B.n213 B.n68 71.676
R848 B.n217 B.n69 71.676
R849 B.n221 B.n70 71.676
R850 B.n226 B.n71 71.676
R851 B.n230 B.n72 71.676
R852 B.n234 B.n73 71.676
R853 B.n238 B.n74 71.676
R854 B.n242 B.n75 71.676
R855 B.n246 B.n76 71.676
R856 B.n250 B.n77 71.676
R857 B.n254 B.n78 71.676
R858 B.n258 B.n79 71.676
R859 B.n262 B.n80 71.676
R860 B.n266 B.n81 71.676
R861 B.n270 B.n82 71.676
R862 B.n274 B.n83 71.676
R863 B.n278 B.n84 71.676
R864 B.n282 B.n85 71.676
R865 B.n286 B.n86 71.676
R866 B.n290 B.n87 71.676
R867 B.n294 B.n88 71.676
R868 B.n298 B.n89 71.676
R869 B.n302 B.n90 71.676
R870 B.n306 B.n91 71.676
R871 B.n310 B.n92 71.676
R872 B.n314 B.n93 71.676
R873 B.n318 B.n94 71.676
R874 B.n322 B.n95 71.676
R875 B.n326 B.n96 71.676
R876 B.n330 B.n97 71.676
R877 B.n334 B.n98 71.676
R878 B.n338 B.n99 71.676
R879 B.n342 B.n100 71.676
R880 B.n346 B.n101 71.676
R881 B.n350 B.n102 71.676
R882 B.n103 B.n102 71.676
R883 B.n349 B.n101 71.676
R884 B.n345 B.n100 71.676
R885 B.n341 B.n99 71.676
R886 B.n337 B.n98 71.676
R887 B.n333 B.n97 71.676
R888 B.n329 B.n96 71.676
R889 B.n325 B.n95 71.676
R890 B.n321 B.n94 71.676
R891 B.n317 B.n93 71.676
R892 B.n313 B.n92 71.676
R893 B.n309 B.n91 71.676
R894 B.n305 B.n90 71.676
R895 B.n301 B.n89 71.676
R896 B.n297 B.n88 71.676
R897 B.n293 B.n87 71.676
R898 B.n289 B.n86 71.676
R899 B.n285 B.n85 71.676
R900 B.n281 B.n84 71.676
R901 B.n277 B.n83 71.676
R902 B.n273 B.n82 71.676
R903 B.n269 B.n81 71.676
R904 B.n265 B.n80 71.676
R905 B.n261 B.n79 71.676
R906 B.n257 B.n78 71.676
R907 B.n253 B.n77 71.676
R908 B.n249 B.n76 71.676
R909 B.n245 B.n75 71.676
R910 B.n241 B.n74 71.676
R911 B.n237 B.n73 71.676
R912 B.n233 B.n72 71.676
R913 B.n229 B.n71 71.676
R914 B.n225 B.n70 71.676
R915 B.n220 B.n69 71.676
R916 B.n216 B.n68 71.676
R917 B.n212 B.n67 71.676
R918 B.n208 B.n66 71.676
R919 B.n204 B.n65 71.676
R920 B.n200 B.n64 71.676
R921 B.n196 B.n63 71.676
R922 B.n192 B.n62 71.676
R923 B.n188 B.n61 71.676
R924 B.n184 B.n60 71.676
R925 B.n180 B.n59 71.676
R926 B.n176 B.n58 71.676
R927 B.n172 B.n57 71.676
R928 B.n168 B.n56 71.676
R929 B.n164 B.n55 71.676
R930 B.n160 B.n54 71.676
R931 B.n156 B.n53 71.676
R932 B.n152 B.n52 71.676
R933 B.n148 B.n51 71.676
R934 B.n144 B.n50 71.676
R935 B.n140 B.n49 71.676
R936 B.n136 B.n48 71.676
R937 B.n132 B.n47 71.676
R938 B.n128 B.n46 71.676
R939 B.n124 B.n45 71.676
R940 B.n120 B.n44 71.676
R941 B.n116 B.n43 71.676
R942 B.n112 B.n42 71.676
R943 B.n701 B.n454 71.676
R944 B.n693 B.n394 71.676
R945 B.n689 B.n395 71.676
R946 B.n685 B.n396 71.676
R947 B.n681 B.n397 71.676
R948 B.n677 B.n398 71.676
R949 B.n673 B.n399 71.676
R950 B.n669 B.n400 71.676
R951 B.n665 B.n401 71.676
R952 B.n661 B.n402 71.676
R953 B.n657 B.n403 71.676
R954 B.n653 B.n404 71.676
R955 B.n649 B.n405 71.676
R956 B.n645 B.n406 71.676
R957 B.n641 B.n407 71.676
R958 B.n637 B.n408 71.676
R959 B.n633 B.n409 71.676
R960 B.n629 B.n410 71.676
R961 B.n625 B.n411 71.676
R962 B.n621 B.n412 71.676
R963 B.n617 B.n413 71.676
R964 B.n613 B.n414 71.676
R965 B.n609 B.n415 71.676
R966 B.n605 B.n416 71.676
R967 B.n601 B.n417 71.676
R968 B.n597 B.n418 71.676
R969 B.n593 B.n419 71.676
R970 B.n589 B.n420 71.676
R971 B.n585 B.n421 71.676
R972 B.n581 B.n422 71.676
R973 B.n577 B.n423 71.676
R974 B.n573 B.n424 71.676
R975 B.n568 B.n425 71.676
R976 B.n564 B.n426 71.676
R977 B.n560 B.n427 71.676
R978 B.n556 B.n428 71.676
R979 B.n552 B.n429 71.676
R980 B.n548 B.n430 71.676
R981 B.n544 B.n431 71.676
R982 B.n540 B.n432 71.676
R983 B.n536 B.n433 71.676
R984 B.n532 B.n434 71.676
R985 B.n528 B.n435 71.676
R986 B.n524 B.n436 71.676
R987 B.n520 B.n437 71.676
R988 B.n516 B.n438 71.676
R989 B.n512 B.n439 71.676
R990 B.n508 B.n440 71.676
R991 B.n504 B.n441 71.676
R992 B.n500 B.n442 71.676
R993 B.n496 B.n443 71.676
R994 B.n492 B.n444 71.676
R995 B.n488 B.n445 71.676
R996 B.n484 B.n446 71.676
R997 B.n480 B.n447 71.676
R998 B.n476 B.n448 71.676
R999 B.n472 B.n449 71.676
R1000 B.n468 B.n450 71.676
R1001 B.n464 B.n451 71.676
R1002 B.n460 B.n452 71.676
R1003 B.n704 B.n703 71.676
R1004 B.n459 B.t8 70.5975
R1005 B.n105 B.t13 70.5975
R1006 B.n456 B.t15 70.5748
R1007 B.n108 B.t19 70.5748
R1008 B.n702 B.n390 62.2415
R1009 B.n799 B.n798 62.2415
R1010 B.n570 B.n459 59.5399
R1011 B.n457 B.n456 59.5399
R1012 B.n223 B.n108 59.5399
R1013 B.n106 B.n105 59.5399
R1014 B.n110 B.n38 34.1859
R1015 B.n796 B.n795 34.1859
R1016 B.n706 B.n705 34.1859
R1017 B.n699 B.n388 34.1859
R1018 B.n709 B.n390 33.3264
R1019 B.n709 B.n385 33.3264
R1020 B.n715 B.n385 33.3264
R1021 B.n715 B.n386 33.3264
R1022 B.n721 B.n378 33.3264
R1023 B.n727 B.n378 33.3264
R1024 B.n727 B.n374 33.3264
R1025 B.n733 B.n374 33.3264
R1026 B.n733 B.n370 33.3264
R1027 B.n739 B.n370 33.3264
R1028 B.n746 B.n366 33.3264
R1029 B.n746 B.n745 33.3264
R1030 B.n752 B.n359 33.3264
R1031 B.n759 B.n359 33.3264
R1032 B.n765 B.n355 33.3264
R1033 B.n765 B.n4 33.3264
R1034 B.n840 B.n4 33.3264
R1035 B.n840 B.n839 33.3264
R1036 B.n839 B.n838 33.3264
R1037 B.n838 B.n8 33.3264
R1038 B.n832 B.n831 33.3264
R1039 B.n831 B.n830 33.3264
R1040 B.n824 B.n18 33.3264
R1041 B.n824 B.n823 33.3264
R1042 B.n822 B.n22 33.3264
R1043 B.n816 B.n22 33.3264
R1044 B.n816 B.n815 33.3264
R1045 B.n815 B.n814 33.3264
R1046 B.n814 B.n29 33.3264
R1047 B.n808 B.n29 33.3264
R1048 B.n807 B.n806 33.3264
R1049 B.n806 B.n36 33.3264
R1050 B.n800 B.n36 33.3264
R1051 B.n800 B.n799 33.3264
R1052 B.n386 B.t7 28.9156
R1053 B.t11 B.n807 28.9156
R1054 B.n759 B.t0 25.9751
R1055 B.n832 B.t3 25.9751
R1056 B.t4 B.n366 23.0346
R1057 B.n823 B.t5 23.0346
R1058 B.n459 B.n458 21.3338
R1059 B.n456 B.n455 21.3338
R1060 B.n108 B.n107 21.3338
R1061 B.n105 B.n104 21.3338
R1062 B.n745 B.t2 18.1337
R1063 B.n18 B.t1 18.1337
R1064 B B.n842 18.0485
R1065 B.n752 B.t2 15.1932
R1066 B.n830 B.t1 15.1932
R1067 B.n111 B.n110 10.6151
R1068 B.n114 B.n111 10.6151
R1069 B.n115 B.n114 10.6151
R1070 B.n118 B.n115 10.6151
R1071 B.n119 B.n118 10.6151
R1072 B.n122 B.n119 10.6151
R1073 B.n123 B.n122 10.6151
R1074 B.n126 B.n123 10.6151
R1075 B.n127 B.n126 10.6151
R1076 B.n130 B.n127 10.6151
R1077 B.n131 B.n130 10.6151
R1078 B.n134 B.n131 10.6151
R1079 B.n135 B.n134 10.6151
R1080 B.n138 B.n135 10.6151
R1081 B.n139 B.n138 10.6151
R1082 B.n142 B.n139 10.6151
R1083 B.n143 B.n142 10.6151
R1084 B.n146 B.n143 10.6151
R1085 B.n147 B.n146 10.6151
R1086 B.n150 B.n147 10.6151
R1087 B.n151 B.n150 10.6151
R1088 B.n154 B.n151 10.6151
R1089 B.n155 B.n154 10.6151
R1090 B.n158 B.n155 10.6151
R1091 B.n159 B.n158 10.6151
R1092 B.n162 B.n159 10.6151
R1093 B.n163 B.n162 10.6151
R1094 B.n166 B.n163 10.6151
R1095 B.n167 B.n166 10.6151
R1096 B.n170 B.n167 10.6151
R1097 B.n171 B.n170 10.6151
R1098 B.n174 B.n171 10.6151
R1099 B.n175 B.n174 10.6151
R1100 B.n178 B.n175 10.6151
R1101 B.n179 B.n178 10.6151
R1102 B.n182 B.n179 10.6151
R1103 B.n183 B.n182 10.6151
R1104 B.n186 B.n183 10.6151
R1105 B.n187 B.n186 10.6151
R1106 B.n190 B.n187 10.6151
R1107 B.n191 B.n190 10.6151
R1108 B.n194 B.n191 10.6151
R1109 B.n195 B.n194 10.6151
R1110 B.n198 B.n195 10.6151
R1111 B.n199 B.n198 10.6151
R1112 B.n202 B.n199 10.6151
R1113 B.n203 B.n202 10.6151
R1114 B.n206 B.n203 10.6151
R1115 B.n207 B.n206 10.6151
R1116 B.n210 B.n207 10.6151
R1117 B.n211 B.n210 10.6151
R1118 B.n214 B.n211 10.6151
R1119 B.n215 B.n214 10.6151
R1120 B.n218 B.n215 10.6151
R1121 B.n219 B.n218 10.6151
R1122 B.n222 B.n219 10.6151
R1123 B.n227 B.n224 10.6151
R1124 B.n228 B.n227 10.6151
R1125 B.n231 B.n228 10.6151
R1126 B.n232 B.n231 10.6151
R1127 B.n235 B.n232 10.6151
R1128 B.n236 B.n235 10.6151
R1129 B.n239 B.n236 10.6151
R1130 B.n240 B.n239 10.6151
R1131 B.n244 B.n243 10.6151
R1132 B.n247 B.n244 10.6151
R1133 B.n248 B.n247 10.6151
R1134 B.n251 B.n248 10.6151
R1135 B.n252 B.n251 10.6151
R1136 B.n255 B.n252 10.6151
R1137 B.n256 B.n255 10.6151
R1138 B.n259 B.n256 10.6151
R1139 B.n260 B.n259 10.6151
R1140 B.n263 B.n260 10.6151
R1141 B.n264 B.n263 10.6151
R1142 B.n267 B.n264 10.6151
R1143 B.n268 B.n267 10.6151
R1144 B.n271 B.n268 10.6151
R1145 B.n272 B.n271 10.6151
R1146 B.n275 B.n272 10.6151
R1147 B.n276 B.n275 10.6151
R1148 B.n279 B.n276 10.6151
R1149 B.n280 B.n279 10.6151
R1150 B.n283 B.n280 10.6151
R1151 B.n284 B.n283 10.6151
R1152 B.n287 B.n284 10.6151
R1153 B.n288 B.n287 10.6151
R1154 B.n291 B.n288 10.6151
R1155 B.n292 B.n291 10.6151
R1156 B.n295 B.n292 10.6151
R1157 B.n296 B.n295 10.6151
R1158 B.n299 B.n296 10.6151
R1159 B.n300 B.n299 10.6151
R1160 B.n303 B.n300 10.6151
R1161 B.n304 B.n303 10.6151
R1162 B.n307 B.n304 10.6151
R1163 B.n308 B.n307 10.6151
R1164 B.n311 B.n308 10.6151
R1165 B.n312 B.n311 10.6151
R1166 B.n315 B.n312 10.6151
R1167 B.n316 B.n315 10.6151
R1168 B.n319 B.n316 10.6151
R1169 B.n320 B.n319 10.6151
R1170 B.n323 B.n320 10.6151
R1171 B.n324 B.n323 10.6151
R1172 B.n327 B.n324 10.6151
R1173 B.n328 B.n327 10.6151
R1174 B.n331 B.n328 10.6151
R1175 B.n332 B.n331 10.6151
R1176 B.n335 B.n332 10.6151
R1177 B.n336 B.n335 10.6151
R1178 B.n339 B.n336 10.6151
R1179 B.n340 B.n339 10.6151
R1180 B.n343 B.n340 10.6151
R1181 B.n344 B.n343 10.6151
R1182 B.n347 B.n344 10.6151
R1183 B.n348 B.n347 10.6151
R1184 B.n351 B.n348 10.6151
R1185 B.n352 B.n351 10.6151
R1186 B.n796 B.n352 10.6151
R1187 B.n707 B.n706 10.6151
R1188 B.n707 B.n383 10.6151
R1189 B.n717 B.n383 10.6151
R1190 B.n718 B.n717 10.6151
R1191 B.n719 B.n718 10.6151
R1192 B.n719 B.n376 10.6151
R1193 B.n729 B.n376 10.6151
R1194 B.n730 B.n729 10.6151
R1195 B.n731 B.n730 10.6151
R1196 B.n731 B.n368 10.6151
R1197 B.n741 B.n368 10.6151
R1198 B.n742 B.n741 10.6151
R1199 B.n743 B.n742 10.6151
R1200 B.n743 B.n361 10.6151
R1201 B.n754 B.n361 10.6151
R1202 B.n755 B.n754 10.6151
R1203 B.n757 B.n755 10.6151
R1204 B.n757 B.n756 10.6151
R1205 B.n756 B.n353 10.6151
R1206 B.n768 B.n353 10.6151
R1207 B.n769 B.n768 10.6151
R1208 B.n770 B.n769 10.6151
R1209 B.n771 B.n770 10.6151
R1210 B.n773 B.n771 10.6151
R1211 B.n774 B.n773 10.6151
R1212 B.n775 B.n774 10.6151
R1213 B.n776 B.n775 10.6151
R1214 B.n778 B.n776 10.6151
R1215 B.n779 B.n778 10.6151
R1216 B.n780 B.n779 10.6151
R1217 B.n781 B.n780 10.6151
R1218 B.n783 B.n781 10.6151
R1219 B.n784 B.n783 10.6151
R1220 B.n785 B.n784 10.6151
R1221 B.n786 B.n785 10.6151
R1222 B.n788 B.n786 10.6151
R1223 B.n789 B.n788 10.6151
R1224 B.n790 B.n789 10.6151
R1225 B.n791 B.n790 10.6151
R1226 B.n793 B.n791 10.6151
R1227 B.n794 B.n793 10.6151
R1228 B.n795 B.n794 10.6151
R1229 B.n699 B.n698 10.6151
R1230 B.n698 B.n697 10.6151
R1231 B.n697 B.n696 10.6151
R1232 B.n696 B.n694 10.6151
R1233 B.n694 B.n691 10.6151
R1234 B.n691 B.n690 10.6151
R1235 B.n690 B.n687 10.6151
R1236 B.n687 B.n686 10.6151
R1237 B.n686 B.n683 10.6151
R1238 B.n683 B.n682 10.6151
R1239 B.n682 B.n679 10.6151
R1240 B.n679 B.n678 10.6151
R1241 B.n678 B.n675 10.6151
R1242 B.n675 B.n674 10.6151
R1243 B.n674 B.n671 10.6151
R1244 B.n671 B.n670 10.6151
R1245 B.n670 B.n667 10.6151
R1246 B.n667 B.n666 10.6151
R1247 B.n666 B.n663 10.6151
R1248 B.n663 B.n662 10.6151
R1249 B.n662 B.n659 10.6151
R1250 B.n659 B.n658 10.6151
R1251 B.n658 B.n655 10.6151
R1252 B.n655 B.n654 10.6151
R1253 B.n654 B.n651 10.6151
R1254 B.n651 B.n650 10.6151
R1255 B.n650 B.n647 10.6151
R1256 B.n647 B.n646 10.6151
R1257 B.n646 B.n643 10.6151
R1258 B.n643 B.n642 10.6151
R1259 B.n642 B.n639 10.6151
R1260 B.n639 B.n638 10.6151
R1261 B.n638 B.n635 10.6151
R1262 B.n635 B.n634 10.6151
R1263 B.n634 B.n631 10.6151
R1264 B.n631 B.n630 10.6151
R1265 B.n630 B.n627 10.6151
R1266 B.n627 B.n626 10.6151
R1267 B.n626 B.n623 10.6151
R1268 B.n623 B.n622 10.6151
R1269 B.n622 B.n619 10.6151
R1270 B.n619 B.n618 10.6151
R1271 B.n618 B.n615 10.6151
R1272 B.n615 B.n614 10.6151
R1273 B.n614 B.n611 10.6151
R1274 B.n611 B.n610 10.6151
R1275 B.n610 B.n607 10.6151
R1276 B.n607 B.n606 10.6151
R1277 B.n606 B.n603 10.6151
R1278 B.n603 B.n602 10.6151
R1279 B.n602 B.n599 10.6151
R1280 B.n599 B.n598 10.6151
R1281 B.n598 B.n595 10.6151
R1282 B.n595 B.n594 10.6151
R1283 B.n594 B.n591 10.6151
R1284 B.n591 B.n590 10.6151
R1285 B.n587 B.n586 10.6151
R1286 B.n586 B.n583 10.6151
R1287 B.n583 B.n582 10.6151
R1288 B.n582 B.n579 10.6151
R1289 B.n579 B.n578 10.6151
R1290 B.n578 B.n575 10.6151
R1291 B.n575 B.n574 10.6151
R1292 B.n574 B.n571 10.6151
R1293 B.n569 B.n566 10.6151
R1294 B.n566 B.n565 10.6151
R1295 B.n565 B.n562 10.6151
R1296 B.n562 B.n561 10.6151
R1297 B.n561 B.n558 10.6151
R1298 B.n558 B.n557 10.6151
R1299 B.n557 B.n554 10.6151
R1300 B.n554 B.n553 10.6151
R1301 B.n553 B.n550 10.6151
R1302 B.n550 B.n549 10.6151
R1303 B.n549 B.n546 10.6151
R1304 B.n546 B.n545 10.6151
R1305 B.n545 B.n542 10.6151
R1306 B.n542 B.n541 10.6151
R1307 B.n541 B.n538 10.6151
R1308 B.n538 B.n537 10.6151
R1309 B.n537 B.n534 10.6151
R1310 B.n534 B.n533 10.6151
R1311 B.n533 B.n530 10.6151
R1312 B.n530 B.n529 10.6151
R1313 B.n529 B.n526 10.6151
R1314 B.n526 B.n525 10.6151
R1315 B.n525 B.n522 10.6151
R1316 B.n522 B.n521 10.6151
R1317 B.n521 B.n518 10.6151
R1318 B.n518 B.n517 10.6151
R1319 B.n517 B.n514 10.6151
R1320 B.n514 B.n513 10.6151
R1321 B.n513 B.n510 10.6151
R1322 B.n510 B.n509 10.6151
R1323 B.n509 B.n506 10.6151
R1324 B.n506 B.n505 10.6151
R1325 B.n505 B.n502 10.6151
R1326 B.n502 B.n501 10.6151
R1327 B.n501 B.n498 10.6151
R1328 B.n498 B.n497 10.6151
R1329 B.n497 B.n494 10.6151
R1330 B.n494 B.n493 10.6151
R1331 B.n493 B.n490 10.6151
R1332 B.n490 B.n489 10.6151
R1333 B.n489 B.n486 10.6151
R1334 B.n486 B.n485 10.6151
R1335 B.n485 B.n482 10.6151
R1336 B.n482 B.n481 10.6151
R1337 B.n481 B.n478 10.6151
R1338 B.n478 B.n477 10.6151
R1339 B.n477 B.n474 10.6151
R1340 B.n474 B.n473 10.6151
R1341 B.n473 B.n470 10.6151
R1342 B.n470 B.n469 10.6151
R1343 B.n469 B.n466 10.6151
R1344 B.n466 B.n465 10.6151
R1345 B.n465 B.n462 10.6151
R1346 B.n462 B.n461 10.6151
R1347 B.n461 B.n392 10.6151
R1348 B.n705 B.n392 10.6151
R1349 B.n711 B.n388 10.6151
R1350 B.n712 B.n711 10.6151
R1351 B.n713 B.n712 10.6151
R1352 B.n713 B.n380 10.6151
R1353 B.n723 B.n380 10.6151
R1354 B.n724 B.n723 10.6151
R1355 B.n725 B.n724 10.6151
R1356 B.n725 B.n372 10.6151
R1357 B.n735 B.n372 10.6151
R1358 B.n736 B.n735 10.6151
R1359 B.n737 B.n736 10.6151
R1360 B.n737 B.n364 10.6151
R1361 B.n748 B.n364 10.6151
R1362 B.n749 B.n748 10.6151
R1363 B.n750 B.n749 10.6151
R1364 B.n750 B.n357 10.6151
R1365 B.n761 B.n357 10.6151
R1366 B.n762 B.n761 10.6151
R1367 B.n763 B.n762 10.6151
R1368 B.n763 B.n0 10.6151
R1369 B.n836 B.n1 10.6151
R1370 B.n836 B.n835 10.6151
R1371 B.n835 B.n834 10.6151
R1372 B.n834 B.n10 10.6151
R1373 B.n828 B.n10 10.6151
R1374 B.n828 B.n827 10.6151
R1375 B.n827 B.n826 10.6151
R1376 B.n826 B.n16 10.6151
R1377 B.n820 B.n16 10.6151
R1378 B.n820 B.n819 10.6151
R1379 B.n819 B.n818 10.6151
R1380 B.n818 B.n24 10.6151
R1381 B.n812 B.n24 10.6151
R1382 B.n812 B.n811 10.6151
R1383 B.n811 B.n810 10.6151
R1384 B.n810 B.n31 10.6151
R1385 B.n804 B.n31 10.6151
R1386 B.n804 B.n803 10.6151
R1387 B.n803 B.n802 10.6151
R1388 B.n802 B.n38 10.6151
R1389 B.n739 B.t4 10.2923
R1390 B.t5 B.n822 10.2923
R1391 B.t0 B.n355 7.3518
R1392 B.t3 B.n8 7.3518
R1393 B.n224 B.n223 6.5566
R1394 B.n240 B.n106 6.5566
R1395 B.n587 B.n457 6.5566
R1396 B.n571 B.n570 6.5566
R1397 B.n721 B.t7 4.41128
R1398 B.n808 B.t11 4.41128
R1399 B.n223 B.n222 4.05904
R1400 B.n243 B.n106 4.05904
R1401 B.n590 B.n457 4.05904
R1402 B.n570 B.n569 4.05904
R1403 B.n842 B.n0 2.81026
R1404 B.n842 B.n1 2.81026
R1405 VN.n1 VN.t1 611.663
R1406 VN.n7 VN.t4 611.663
R1407 VN.n2 VN.t5 588.73
R1408 VN.n4 VN.t0 588.73
R1409 VN.n8 VN.t3 588.73
R1410 VN.n10 VN.t2 588.73
R1411 VN.n5 VN.n4 161.3
R1412 VN.n11 VN.n10 161.3
R1413 VN.n9 VN.n6 161.3
R1414 VN.n3 VN.n0 161.3
R1415 VN VN.n11 45.8433
R1416 VN.n7 VN.n6 44.8791
R1417 VN.n1 VN.n0 44.8791
R1418 VN.n4 VN.n3 31.4035
R1419 VN.n10 VN.n9 31.4035
R1420 VN.n2 VN.n1 18.8496
R1421 VN.n8 VN.n7 18.8496
R1422 VN.n3 VN.n2 16.7975
R1423 VN.n9 VN.n8 16.7975
R1424 VN.n11 VN.n6 0.189894
R1425 VN.n5 VN.n0 0.189894
R1426 VN VN.n5 0.0516364
R1427 VTAIL.n7 VTAIL.t9 45.3703
R1428 VTAIL.n11 VTAIL.t6 45.3702
R1429 VTAIL.n2 VTAIL.t5 45.3702
R1430 VTAIL.n10 VTAIL.t4 45.3702
R1431 VTAIL.n9 VTAIL.n8 44.2172
R1432 VTAIL.n6 VTAIL.n5 44.2172
R1433 VTAIL.n1 VTAIL.n0 44.217
R1434 VTAIL.n4 VTAIL.n3 44.217
R1435 VTAIL.n6 VTAIL.n4 29.0652
R1436 VTAIL.n11 VTAIL.n10 28.1169
R1437 VTAIL.n0 VTAIL.t7 1.15367
R1438 VTAIL.n0 VTAIL.t10 1.15367
R1439 VTAIL.n3 VTAIL.t1 1.15367
R1440 VTAIL.n3 VTAIL.t2 1.15367
R1441 VTAIL.n8 VTAIL.t0 1.15367
R1442 VTAIL.n8 VTAIL.t3 1.15367
R1443 VTAIL.n5 VTAIL.t11 1.15367
R1444 VTAIL.n5 VTAIL.t8 1.15367
R1445 VTAIL.n7 VTAIL.n6 0.948776
R1446 VTAIL.n10 VTAIL.n9 0.948776
R1447 VTAIL.n4 VTAIL.n2 0.948776
R1448 VTAIL.n9 VTAIL.n7 0.944465
R1449 VTAIL.n2 VTAIL.n1 0.944465
R1450 VTAIL VTAIL.n11 0.653517
R1451 VTAIL VTAIL.n1 0.295759
R1452 VDD2.n1 VDD2.t4 62.7049
R1453 VDD2.n2 VDD2.t3 62.0491
R1454 VDD2.n1 VDD2.n0 61.0775
R1455 VDD2 VDD2.n3 61.0747
R1456 VDD2.n2 VDD2.n1 41.5989
R1457 VDD2.n3 VDD2.t2 1.15367
R1458 VDD2.n3 VDD2.t1 1.15367
R1459 VDD2.n0 VDD2.t0 1.15367
R1460 VDD2.n0 VDD2.t5 1.15367
R1461 VDD2 VDD2.n2 0.769897
R1462 VP.n3 VP.t1 611.663
R1463 VP.n8 VP.t5 588.73
R1464 VP.n12 VP.t2 588.73
R1465 VP.n14 VP.t0 588.73
R1466 VP.n6 VP.t3 588.73
R1467 VP.n4 VP.t4 588.73
R1468 VP.n15 VP.n14 161.3
R1469 VP.n5 VP.n2 161.3
R1470 VP.n7 VP.n6 161.3
R1471 VP.n13 VP.n0 161.3
R1472 VP.n12 VP.n11 161.3
R1473 VP.n10 VP.n1 161.3
R1474 VP.n9 VP.n8 161.3
R1475 VP.n9 VP.n7 45.4626
R1476 VP.n3 VP.n2 44.8791
R1477 VP.n8 VP.n1 31.4035
R1478 VP.n14 VP.n13 31.4035
R1479 VP.n6 VP.n5 31.4035
R1480 VP.n4 VP.n3 18.8496
R1481 VP.n12 VP.n1 16.7975
R1482 VP.n13 VP.n12 16.7975
R1483 VP.n5 VP.n4 16.7975
R1484 VP.n7 VP.n2 0.189894
R1485 VP.n10 VP.n9 0.189894
R1486 VP.n11 VP.n10 0.189894
R1487 VP.n11 VP.n0 0.189894
R1488 VP.n15 VP.n0 0.189894
R1489 VP VP.n15 0.0516364
R1490 VDD1 VDD1.t4 62.8185
R1491 VDD1.n1 VDD1.t0 62.7049
R1492 VDD1.n1 VDD1.n0 61.0775
R1493 VDD1.n3 VDD1.n2 60.8958
R1494 VDD1.n3 VDD1.n1 42.6561
R1495 VDD1.n2 VDD1.t1 1.15367
R1496 VDD1.n2 VDD1.t2 1.15367
R1497 VDD1.n0 VDD1.t3 1.15367
R1498 VDD1.n0 VDD1.t5 1.15367
R1499 VDD1 VDD1.n3 0.179379
C0 VDD1 VTAIL 12.899099f
C1 VP VDD1 6.50458f
C2 VDD2 VDD1 0.736466f
C3 VN VTAIL 5.85647f
C4 VP VN 6.10402f
C5 VDD2 VN 6.35468f
C6 VP VTAIL 5.87126f
C7 VDD2 VTAIL 12.931201f
C8 VP VDD2 0.304139f
C9 VN VDD1 0.148083f
C10 VDD2 B 5.471957f
C11 VDD1 B 5.710626f
C12 VTAIL B 8.365273f
C13 VN B 8.52499f
C14 VP B 6.323803f
C15 VDD1.t4 B 3.64038f
C16 VDD1.t0 B 3.63971f
C17 VDD1.t3 B 0.312978f
C18 VDD1.t5 B 0.312978f
C19 VDD1.n0 B 2.84667f
C20 VDD1.n1 B 2.32352f
C21 VDD1.t1 B 0.312978f
C22 VDD1.t2 B 0.312978f
C23 VDD1.n2 B 2.8458f
C24 VDD1.n3 B 2.46513f
C25 VP.n0 B 0.044662f
C26 VP.n1 B 0.010135f
C27 VP.n2 B 0.190642f
C28 VP.t3 B 1.67534f
C29 VP.t4 B 1.67534f
C30 VP.t1 B 1.69914f
C31 VP.n3 B 0.615076f
C32 VP.n4 B 0.637525f
C33 VP.n5 B 0.010135f
C34 VP.n6 B 0.632451f
C35 VP.n7 B 2.09669f
C36 VP.t5 B 1.67534f
C37 VP.n8 B 0.632451f
C38 VP.n9 B 2.132f
C39 VP.n10 B 0.044662f
C40 VP.n11 B 0.044662f
C41 VP.t2 B 1.67534f
C42 VP.n12 B 0.632864f
C43 VP.n13 B 0.010135f
C44 VP.t0 B 1.67534f
C45 VP.n14 B 0.632451f
C46 VP.n15 B 0.034611f
C47 VDD2.t4 B 3.63692f
C48 VDD2.t0 B 0.312738f
C49 VDD2.t5 B 0.312738f
C50 VDD2.n0 B 2.84448f
C51 VDD2.n1 B 2.24775f
C52 VDD2.t3 B 3.63367f
C53 VDD2.n2 B 2.48839f
C54 VDD2.t2 B 0.312738f
C55 VDD2.t1 B 0.312738f
C56 VDD2.n3 B 2.84445f
C57 VTAIL.t7 B 0.319066f
C58 VTAIL.t10 B 0.319066f
C59 VTAIL.n0 B 2.82945f
C60 VTAIL.n1 B 0.328289f
C61 VTAIL.t5 B 3.6137f
C62 VTAIL.n2 B 0.463703f
C63 VTAIL.t1 B 0.319066f
C64 VTAIL.t2 B 0.319066f
C65 VTAIL.n3 B 2.82945f
C66 VTAIL.n4 B 1.89095f
C67 VTAIL.t11 B 0.319066f
C68 VTAIL.t8 B 0.319066f
C69 VTAIL.n5 B 2.82945f
C70 VTAIL.n6 B 1.89094f
C71 VTAIL.t9 B 3.61372f
C72 VTAIL.n7 B 0.463681f
C73 VTAIL.t0 B 0.319066f
C74 VTAIL.t3 B 0.319066f
C75 VTAIL.n8 B 2.82945f
C76 VTAIL.n9 B 0.377766f
C77 VTAIL.t4 B 3.61369f
C78 VTAIL.n10 B 1.90503f
C79 VTAIL.t6 B 3.6137f
C80 VTAIL.n11 B 1.88266f
C81 VN.n0 B 0.18897f
C82 VN.t1 B 1.68424f
C83 VN.n1 B 0.609682f
C84 VN.t5 B 1.66065f
C85 VN.n2 B 0.631934f
C86 VN.n3 B 0.010046f
C87 VN.t0 B 1.66065f
C88 VN.n4 B 0.626905f
C89 VN.n5 B 0.034308f
C90 VN.n6 B 0.18897f
C91 VN.t4 B 1.68424f
C92 VN.n7 B 0.609682f
C93 VN.t3 B 1.66065f
C94 VN.n8 B 0.631934f
C95 VN.n9 B 0.010046f
C96 VN.t2 B 1.66065f
C97 VN.n10 B 0.626905f
C98 VN.n11 B 2.10723f
.ends

