* NGSPICE file created from diff_pair_sample_0757.ext - technology: sky130A

.subckt diff_pair_sample_0757 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1.7
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1.7
X2 VDD2.t3 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1.7
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1.7
X4 VDD1.t2 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1.7
X5 VTAIL.t7 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1.7
X6 VTAIL.t6 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1.7
X7 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1.7
X8 VDD2.t0 VN.t3 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1.7
X9 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1.7
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1.7
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1.7
R0 B.n343 B.n342 585
R1 B.n345 B.n75 585
R2 B.n348 B.n347 585
R3 B.n349 B.n74 585
R4 B.n351 B.n350 585
R5 B.n353 B.n73 585
R6 B.n356 B.n355 585
R7 B.n357 B.n72 585
R8 B.n359 B.n358 585
R9 B.n361 B.n71 585
R10 B.n364 B.n363 585
R11 B.n365 B.n70 585
R12 B.n367 B.n366 585
R13 B.n369 B.n69 585
R14 B.n372 B.n371 585
R15 B.n374 B.n66 585
R16 B.n376 B.n375 585
R17 B.n378 B.n65 585
R18 B.n381 B.n380 585
R19 B.n382 B.n64 585
R20 B.n384 B.n383 585
R21 B.n386 B.n63 585
R22 B.n389 B.n388 585
R23 B.n390 B.n59 585
R24 B.n392 B.n391 585
R25 B.n394 B.n58 585
R26 B.n397 B.n396 585
R27 B.n398 B.n57 585
R28 B.n400 B.n399 585
R29 B.n402 B.n56 585
R30 B.n405 B.n404 585
R31 B.n406 B.n55 585
R32 B.n408 B.n407 585
R33 B.n410 B.n54 585
R34 B.n413 B.n412 585
R35 B.n414 B.n53 585
R36 B.n416 B.n415 585
R37 B.n418 B.n52 585
R38 B.n421 B.n420 585
R39 B.n422 B.n51 585
R40 B.n341 B.n49 585
R41 B.n425 B.n49 585
R42 B.n340 B.n48 585
R43 B.n426 B.n48 585
R44 B.n339 B.n47 585
R45 B.n427 B.n47 585
R46 B.n338 B.n337 585
R47 B.n337 B.n43 585
R48 B.n336 B.n42 585
R49 B.n433 B.n42 585
R50 B.n335 B.n41 585
R51 B.n434 B.n41 585
R52 B.n334 B.n40 585
R53 B.n435 B.n40 585
R54 B.n333 B.n332 585
R55 B.n332 B.n36 585
R56 B.n331 B.n35 585
R57 B.n441 B.n35 585
R58 B.n330 B.n34 585
R59 B.n442 B.n34 585
R60 B.n329 B.n33 585
R61 B.n443 B.n33 585
R62 B.n328 B.n327 585
R63 B.n327 B.n29 585
R64 B.n326 B.n28 585
R65 B.n449 B.n28 585
R66 B.n325 B.n27 585
R67 B.n450 B.n27 585
R68 B.n324 B.n26 585
R69 B.n451 B.n26 585
R70 B.n323 B.n322 585
R71 B.n322 B.n25 585
R72 B.n321 B.n21 585
R73 B.n457 B.n21 585
R74 B.n320 B.n20 585
R75 B.n458 B.n20 585
R76 B.n319 B.n19 585
R77 B.n459 B.n19 585
R78 B.n318 B.n317 585
R79 B.n317 B.n15 585
R80 B.n316 B.n14 585
R81 B.n465 B.n14 585
R82 B.n315 B.n13 585
R83 B.n466 B.n13 585
R84 B.n314 B.n12 585
R85 B.n467 B.n12 585
R86 B.n313 B.n312 585
R87 B.n312 B.n8 585
R88 B.n311 B.n7 585
R89 B.n473 B.n7 585
R90 B.n310 B.n6 585
R91 B.n474 B.n6 585
R92 B.n309 B.n5 585
R93 B.n475 B.n5 585
R94 B.n308 B.n307 585
R95 B.n307 B.n4 585
R96 B.n306 B.n76 585
R97 B.n306 B.n305 585
R98 B.n296 B.n77 585
R99 B.n78 B.n77 585
R100 B.n298 B.n297 585
R101 B.n299 B.n298 585
R102 B.n295 B.n82 585
R103 B.n86 B.n82 585
R104 B.n294 B.n293 585
R105 B.n293 B.n292 585
R106 B.n84 B.n83 585
R107 B.n85 B.n84 585
R108 B.n285 B.n284 585
R109 B.n286 B.n285 585
R110 B.n283 B.n91 585
R111 B.n91 B.n90 585
R112 B.n282 B.n281 585
R113 B.n281 B.n280 585
R114 B.n93 B.n92 585
R115 B.n273 B.n93 585
R116 B.n272 B.n271 585
R117 B.n274 B.n272 585
R118 B.n270 B.n98 585
R119 B.n98 B.n97 585
R120 B.n269 B.n268 585
R121 B.n268 B.n267 585
R122 B.n100 B.n99 585
R123 B.n101 B.n100 585
R124 B.n260 B.n259 585
R125 B.n261 B.n260 585
R126 B.n258 B.n106 585
R127 B.n106 B.n105 585
R128 B.n257 B.n256 585
R129 B.n256 B.n255 585
R130 B.n108 B.n107 585
R131 B.n109 B.n108 585
R132 B.n248 B.n247 585
R133 B.n249 B.n248 585
R134 B.n246 B.n114 585
R135 B.n114 B.n113 585
R136 B.n245 B.n244 585
R137 B.n244 B.n243 585
R138 B.n116 B.n115 585
R139 B.n117 B.n116 585
R140 B.n236 B.n235 585
R141 B.n237 B.n236 585
R142 B.n234 B.n122 585
R143 B.n122 B.n121 585
R144 B.n233 B.n232 585
R145 B.n232 B.n231 585
R146 B.n228 B.n126 585
R147 B.n227 B.n226 585
R148 B.n224 B.n127 585
R149 B.n224 B.n125 585
R150 B.n223 B.n222 585
R151 B.n221 B.n220 585
R152 B.n219 B.n129 585
R153 B.n217 B.n216 585
R154 B.n215 B.n130 585
R155 B.n214 B.n213 585
R156 B.n211 B.n131 585
R157 B.n209 B.n208 585
R158 B.n207 B.n132 585
R159 B.n206 B.n205 585
R160 B.n203 B.n133 585
R161 B.n201 B.n200 585
R162 B.n198 B.n134 585
R163 B.n197 B.n196 585
R164 B.n194 B.n137 585
R165 B.n192 B.n191 585
R166 B.n190 B.n138 585
R167 B.n189 B.n188 585
R168 B.n186 B.n139 585
R169 B.n184 B.n183 585
R170 B.n182 B.n140 585
R171 B.n181 B.n180 585
R172 B.n178 B.n177 585
R173 B.n176 B.n175 585
R174 B.n174 B.n145 585
R175 B.n172 B.n171 585
R176 B.n170 B.n146 585
R177 B.n169 B.n168 585
R178 B.n166 B.n147 585
R179 B.n164 B.n163 585
R180 B.n162 B.n148 585
R181 B.n161 B.n160 585
R182 B.n158 B.n149 585
R183 B.n156 B.n155 585
R184 B.n154 B.n150 585
R185 B.n153 B.n152 585
R186 B.n124 B.n123 585
R187 B.n125 B.n124 585
R188 B.n230 B.n229 585
R189 B.n231 B.n230 585
R190 B.n120 B.n119 585
R191 B.n121 B.n120 585
R192 B.n239 B.n238 585
R193 B.n238 B.n237 585
R194 B.n240 B.n118 585
R195 B.n118 B.n117 585
R196 B.n242 B.n241 585
R197 B.n243 B.n242 585
R198 B.n112 B.n111 585
R199 B.n113 B.n112 585
R200 B.n251 B.n250 585
R201 B.n250 B.n249 585
R202 B.n252 B.n110 585
R203 B.n110 B.n109 585
R204 B.n254 B.n253 585
R205 B.n255 B.n254 585
R206 B.n104 B.n103 585
R207 B.n105 B.n104 585
R208 B.n263 B.n262 585
R209 B.n262 B.n261 585
R210 B.n264 B.n102 585
R211 B.n102 B.n101 585
R212 B.n266 B.n265 585
R213 B.n267 B.n266 585
R214 B.n96 B.n95 585
R215 B.n97 B.n96 585
R216 B.n276 B.n275 585
R217 B.n275 B.n274 585
R218 B.n277 B.n94 585
R219 B.n273 B.n94 585
R220 B.n279 B.n278 585
R221 B.n280 B.n279 585
R222 B.n89 B.n88 585
R223 B.n90 B.n89 585
R224 B.n288 B.n287 585
R225 B.n287 B.n286 585
R226 B.n289 B.n87 585
R227 B.n87 B.n85 585
R228 B.n291 B.n290 585
R229 B.n292 B.n291 585
R230 B.n81 B.n80 585
R231 B.n86 B.n81 585
R232 B.n301 B.n300 585
R233 B.n300 B.n299 585
R234 B.n302 B.n79 585
R235 B.n79 B.n78 585
R236 B.n304 B.n303 585
R237 B.n305 B.n304 585
R238 B.n2 B.n0 585
R239 B.n4 B.n2 585
R240 B.n3 B.n1 585
R241 B.n474 B.n3 585
R242 B.n472 B.n471 585
R243 B.n473 B.n472 585
R244 B.n470 B.n9 585
R245 B.n9 B.n8 585
R246 B.n469 B.n468 585
R247 B.n468 B.n467 585
R248 B.n11 B.n10 585
R249 B.n466 B.n11 585
R250 B.n464 B.n463 585
R251 B.n465 B.n464 585
R252 B.n462 B.n16 585
R253 B.n16 B.n15 585
R254 B.n461 B.n460 585
R255 B.n460 B.n459 585
R256 B.n18 B.n17 585
R257 B.n458 B.n18 585
R258 B.n456 B.n455 585
R259 B.n457 B.n456 585
R260 B.n454 B.n22 585
R261 B.n25 B.n22 585
R262 B.n453 B.n452 585
R263 B.n452 B.n451 585
R264 B.n24 B.n23 585
R265 B.n450 B.n24 585
R266 B.n448 B.n447 585
R267 B.n449 B.n448 585
R268 B.n446 B.n30 585
R269 B.n30 B.n29 585
R270 B.n445 B.n444 585
R271 B.n444 B.n443 585
R272 B.n32 B.n31 585
R273 B.n442 B.n32 585
R274 B.n440 B.n439 585
R275 B.n441 B.n440 585
R276 B.n438 B.n37 585
R277 B.n37 B.n36 585
R278 B.n437 B.n436 585
R279 B.n436 B.n435 585
R280 B.n39 B.n38 585
R281 B.n434 B.n39 585
R282 B.n432 B.n431 585
R283 B.n433 B.n432 585
R284 B.n430 B.n44 585
R285 B.n44 B.n43 585
R286 B.n429 B.n428 585
R287 B.n428 B.n427 585
R288 B.n46 B.n45 585
R289 B.n426 B.n46 585
R290 B.n424 B.n423 585
R291 B.n425 B.n424 585
R292 B.n477 B.n476 585
R293 B.n476 B.n475 585
R294 B.n230 B.n126 492.5
R295 B.n424 B.n51 492.5
R296 B.n232 B.n124 492.5
R297 B.n343 B.n49 492.5
R298 B.n344 B.n50 256.663
R299 B.n346 B.n50 256.663
R300 B.n352 B.n50 256.663
R301 B.n354 B.n50 256.663
R302 B.n360 B.n50 256.663
R303 B.n362 B.n50 256.663
R304 B.n368 B.n50 256.663
R305 B.n370 B.n50 256.663
R306 B.n377 B.n50 256.663
R307 B.n379 B.n50 256.663
R308 B.n385 B.n50 256.663
R309 B.n387 B.n50 256.663
R310 B.n393 B.n50 256.663
R311 B.n395 B.n50 256.663
R312 B.n401 B.n50 256.663
R313 B.n403 B.n50 256.663
R314 B.n409 B.n50 256.663
R315 B.n411 B.n50 256.663
R316 B.n417 B.n50 256.663
R317 B.n419 B.n50 256.663
R318 B.n225 B.n125 256.663
R319 B.n128 B.n125 256.663
R320 B.n218 B.n125 256.663
R321 B.n212 B.n125 256.663
R322 B.n210 B.n125 256.663
R323 B.n204 B.n125 256.663
R324 B.n202 B.n125 256.663
R325 B.n195 B.n125 256.663
R326 B.n193 B.n125 256.663
R327 B.n187 B.n125 256.663
R328 B.n185 B.n125 256.663
R329 B.n179 B.n125 256.663
R330 B.n144 B.n125 256.663
R331 B.n173 B.n125 256.663
R332 B.n167 B.n125 256.663
R333 B.n165 B.n125 256.663
R334 B.n159 B.n125 256.663
R335 B.n157 B.n125 256.663
R336 B.n151 B.n125 256.663
R337 B.n141 B.t4 248.643
R338 B.n135 B.t8 248.643
R339 B.n60 B.t15 248.643
R340 B.n67 B.t11 248.643
R341 B.n231 B.n125 166.163
R342 B.n425 B.n50 166.163
R343 B.n230 B.n120 163.367
R344 B.n238 B.n120 163.367
R345 B.n238 B.n118 163.367
R346 B.n242 B.n118 163.367
R347 B.n242 B.n112 163.367
R348 B.n250 B.n112 163.367
R349 B.n250 B.n110 163.367
R350 B.n254 B.n110 163.367
R351 B.n254 B.n104 163.367
R352 B.n262 B.n104 163.367
R353 B.n262 B.n102 163.367
R354 B.n266 B.n102 163.367
R355 B.n266 B.n96 163.367
R356 B.n275 B.n96 163.367
R357 B.n275 B.n94 163.367
R358 B.n279 B.n94 163.367
R359 B.n279 B.n89 163.367
R360 B.n287 B.n89 163.367
R361 B.n287 B.n87 163.367
R362 B.n291 B.n87 163.367
R363 B.n291 B.n81 163.367
R364 B.n300 B.n81 163.367
R365 B.n300 B.n79 163.367
R366 B.n304 B.n79 163.367
R367 B.n304 B.n2 163.367
R368 B.n476 B.n2 163.367
R369 B.n476 B.n3 163.367
R370 B.n472 B.n3 163.367
R371 B.n472 B.n9 163.367
R372 B.n468 B.n9 163.367
R373 B.n468 B.n11 163.367
R374 B.n464 B.n11 163.367
R375 B.n464 B.n16 163.367
R376 B.n460 B.n16 163.367
R377 B.n460 B.n18 163.367
R378 B.n456 B.n18 163.367
R379 B.n456 B.n22 163.367
R380 B.n452 B.n22 163.367
R381 B.n452 B.n24 163.367
R382 B.n448 B.n24 163.367
R383 B.n448 B.n30 163.367
R384 B.n444 B.n30 163.367
R385 B.n444 B.n32 163.367
R386 B.n440 B.n32 163.367
R387 B.n440 B.n37 163.367
R388 B.n436 B.n37 163.367
R389 B.n436 B.n39 163.367
R390 B.n432 B.n39 163.367
R391 B.n432 B.n44 163.367
R392 B.n428 B.n44 163.367
R393 B.n428 B.n46 163.367
R394 B.n424 B.n46 163.367
R395 B.n226 B.n224 163.367
R396 B.n224 B.n223 163.367
R397 B.n220 B.n219 163.367
R398 B.n217 B.n130 163.367
R399 B.n213 B.n211 163.367
R400 B.n209 B.n132 163.367
R401 B.n205 B.n203 163.367
R402 B.n201 B.n134 163.367
R403 B.n196 B.n194 163.367
R404 B.n192 B.n138 163.367
R405 B.n188 B.n186 163.367
R406 B.n184 B.n140 163.367
R407 B.n180 B.n178 163.367
R408 B.n175 B.n174 163.367
R409 B.n172 B.n146 163.367
R410 B.n168 B.n166 163.367
R411 B.n164 B.n148 163.367
R412 B.n160 B.n158 163.367
R413 B.n156 B.n150 163.367
R414 B.n152 B.n124 163.367
R415 B.n232 B.n122 163.367
R416 B.n236 B.n122 163.367
R417 B.n236 B.n116 163.367
R418 B.n244 B.n116 163.367
R419 B.n244 B.n114 163.367
R420 B.n248 B.n114 163.367
R421 B.n248 B.n108 163.367
R422 B.n256 B.n108 163.367
R423 B.n256 B.n106 163.367
R424 B.n260 B.n106 163.367
R425 B.n260 B.n100 163.367
R426 B.n268 B.n100 163.367
R427 B.n268 B.n98 163.367
R428 B.n272 B.n98 163.367
R429 B.n272 B.n93 163.367
R430 B.n281 B.n93 163.367
R431 B.n281 B.n91 163.367
R432 B.n285 B.n91 163.367
R433 B.n285 B.n84 163.367
R434 B.n293 B.n84 163.367
R435 B.n293 B.n82 163.367
R436 B.n298 B.n82 163.367
R437 B.n298 B.n77 163.367
R438 B.n306 B.n77 163.367
R439 B.n307 B.n306 163.367
R440 B.n307 B.n5 163.367
R441 B.n6 B.n5 163.367
R442 B.n7 B.n6 163.367
R443 B.n312 B.n7 163.367
R444 B.n312 B.n12 163.367
R445 B.n13 B.n12 163.367
R446 B.n14 B.n13 163.367
R447 B.n317 B.n14 163.367
R448 B.n317 B.n19 163.367
R449 B.n20 B.n19 163.367
R450 B.n21 B.n20 163.367
R451 B.n322 B.n21 163.367
R452 B.n322 B.n26 163.367
R453 B.n27 B.n26 163.367
R454 B.n28 B.n27 163.367
R455 B.n327 B.n28 163.367
R456 B.n327 B.n33 163.367
R457 B.n34 B.n33 163.367
R458 B.n35 B.n34 163.367
R459 B.n332 B.n35 163.367
R460 B.n332 B.n40 163.367
R461 B.n41 B.n40 163.367
R462 B.n42 B.n41 163.367
R463 B.n337 B.n42 163.367
R464 B.n337 B.n47 163.367
R465 B.n48 B.n47 163.367
R466 B.n49 B.n48 163.367
R467 B.n420 B.n418 163.367
R468 B.n416 B.n53 163.367
R469 B.n412 B.n410 163.367
R470 B.n408 B.n55 163.367
R471 B.n404 B.n402 163.367
R472 B.n400 B.n57 163.367
R473 B.n396 B.n394 163.367
R474 B.n392 B.n59 163.367
R475 B.n388 B.n386 163.367
R476 B.n384 B.n64 163.367
R477 B.n380 B.n378 163.367
R478 B.n376 B.n66 163.367
R479 B.n371 B.n369 163.367
R480 B.n367 B.n70 163.367
R481 B.n363 B.n361 163.367
R482 B.n359 B.n72 163.367
R483 B.n355 B.n353 163.367
R484 B.n351 B.n74 163.367
R485 B.n347 B.n345 163.367
R486 B.n141 B.t7 119.984
R487 B.n67 B.t13 119.984
R488 B.n135 B.t10 119.983
R489 B.n60 B.t16 119.983
R490 B.n231 B.n121 90.3933
R491 B.n237 B.n121 90.3933
R492 B.n237 B.n117 90.3933
R493 B.n243 B.n117 90.3933
R494 B.n243 B.n113 90.3933
R495 B.n249 B.n113 90.3933
R496 B.n255 B.n109 90.3933
R497 B.n255 B.n105 90.3933
R498 B.n261 B.n105 90.3933
R499 B.n261 B.n101 90.3933
R500 B.n267 B.n101 90.3933
R501 B.n267 B.n97 90.3933
R502 B.n274 B.n97 90.3933
R503 B.n274 B.n273 90.3933
R504 B.n280 B.n90 90.3933
R505 B.n286 B.n90 90.3933
R506 B.n286 B.n85 90.3933
R507 B.n292 B.n85 90.3933
R508 B.n292 B.n86 90.3933
R509 B.n299 B.n78 90.3933
R510 B.n305 B.n78 90.3933
R511 B.n305 B.n4 90.3933
R512 B.n475 B.n4 90.3933
R513 B.n475 B.n474 90.3933
R514 B.n474 B.n473 90.3933
R515 B.n473 B.n8 90.3933
R516 B.n467 B.n8 90.3933
R517 B.n466 B.n465 90.3933
R518 B.n465 B.n15 90.3933
R519 B.n459 B.n15 90.3933
R520 B.n459 B.n458 90.3933
R521 B.n458 B.n457 90.3933
R522 B.n451 B.n25 90.3933
R523 B.n451 B.n450 90.3933
R524 B.n450 B.n449 90.3933
R525 B.n449 B.n29 90.3933
R526 B.n443 B.n29 90.3933
R527 B.n443 B.n442 90.3933
R528 B.n442 B.n441 90.3933
R529 B.n441 B.n36 90.3933
R530 B.n435 B.n434 90.3933
R531 B.n434 B.n433 90.3933
R532 B.n433 B.n43 90.3933
R533 B.n427 B.n43 90.3933
R534 B.n427 B.n426 90.3933
R535 B.n426 B.n425 90.3933
R536 B.n142 B.t6 80.6148
R537 B.n68 B.t14 80.6148
R538 B.n136 B.t9 80.613
R539 B.n61 B.t17 80.613
R540 B.n225 B.n126 71.676
R541 B.n223 B.n128 71.676
R542 B.n219 B.n218 71.676
R543 B.n212 B.n130 71.676
R544 B.n211 B.n210 71.676
R545 B.n204 B.n132 71.676
R546 B.n203 B.n202 71.676
R547 B.n195 B.n134 71.676
R548 B.n194 B.n193 71.676
R549 B.n187 B.n138 71.676
R550 B.n186 B.n185 71.676
R551 B.n179 B.n140 71.676
R552 B.n178 B.n144 71.676
R553 B.n174 B.n173 71.676
R554 B.n167 B.n146 71.676
R555 B.n166 B.n165 71.676
R556 B.n159 B.n148 71.676
R557 B.n158 B.n157 71.676
R558 B.n151 B.n150 71.676
R559 B.n419 B.n51 71.676
R560 B.n418 B.n417 71.676
R561 B.n411 B.n53 71.676
R562 B.n410 B.n409 71.676
R563 B.n403 B.n55 71.676
R564 B.n402 B.n401 71.676
R565 B.n395 B.n57 71.676
R566 B.n394 B.n393 71.676
R567 B.n387 B.n59 71.676
R568 B.n386 B.n385 71.676
R569 B.n379 B.n64 71.676
R570 B.n378 B.n377 71.676
R571 B.n370 B.n66 71.676
R572 B.n369 B.n368 71.676
R573 B.n362 B.n70 71.676
R574 B.n361 B.n360 71.676
R575 B.n354 B.n72 71.676
R576 B.n353 B.n352 71.676
R577 B.n346 B.n74 71.676
R578 B.n345 B.n344 71.676
R579 B.n344 B.n343 71.676
R580 B.n347 B.n346 71.676
R581 B.n352 B.n351 71.676
R582 B.n355 B.n354 71.676
R583 B.n360 B.n359 71.676
R584 B.n363 B.n362 71.676
R585 B.n368 B.n367 71.676
R586 B.n371 B.n370 71.676
R587 B.n377 B.n376 71.676
R588 B.n380 B.n379 71.676
R589 B.n385 B.n384 71.676
R590 B.n388 B.n387 71.676
R591 B.n393 B.n392 71.676
R592 B.n396 B.n395 71.676
R593 B.n401 B.n400 71.676
R594 B.n404 B.n403 71.676
R595 B.n409 B.n408 71.676
R596 B.n412 B.n411 71.676
R597 B.n417 B.n416 71.676
R598 B.n420 B.n419 71.676
R599 B.n226 B.n225 71.676
R600 B.n220 B.n128 71.676
R601 B.n218 B.n217 71.676
R602 B.n213 B.n212 71.676
R603 B.n210 B.n209 71.676
R604 B.n205 B.n204 71.676
R605 B.n202 B.n201 71.676
R606 B.n196 B.n195 71.676
R607 B.n193 B.n192 71.676
R608 B.n188 B.n187 71.676
R609 B.n185 B.n184 71.676
R610 B.n180 B.n179 71.676
R611 B.n175 B.n144 71.676
R612 B.n173 B.n172 71.676
R613 B.n168 B.n167 71.676
R614 B.n165 B.n164 71.676
R615 B.n160 B.n159 71.676
R616 B.n157 B.n156 71.676
R617 B.n152 B.n151 71.676
R618 B.t5 B.n109 66.4658
R619 B.t12 B.n36 66.4658
R620 B.n143 B.n142 59.5399
R621 B.n199 B.n136 59.5399
R622 B.n62 B.n61 59.5399
R623 B.n373 B.n68 59.5399
R624 B.n299 B.t2 53.1727
R625 B.n467 B.t3 53.1727
R626 B.n280 B.t1 50.5141
R627 B.n457 B.t0 50.5141
R628 B.n273 B.t1 39.8797
R629 B.n25 B.t0 39.8797
R630 B.n142 B.n141 39.3702
R631 B.n136 B.n135 39.3702
R632 B.n61 B.n60 39.3702
R633 B.n68 B.n67 39.3702
R634 B.n86 B.t2 37.221
R635 B.t3 B.n466 37.221
R636 B.n423 B.n422 32.0005
R637 B.n342 B.n341 32.0005
R638 B.n233 B.n123 32.0005
R639 B.n229 B.n228 32.0005
R640 B.n249 B.t5 23.928
R641 B.n435 B.t12 23.928
R642 B B.n477 18.0485
R643 B.n422 B.n421 10.6151
R644 B.n421 B.n52 10.6151
R645 B.n415 B.n52 10.6151
R646 B.n415 B.n414 10.6151
R647 B.n414 B.n413 10.6151
R648 B.n413 B.n54 10.6151
R649 B.n407 B.n54 10.6151
R650 B.n407 B.n406 10.6151
R651 B.n406 B.n405 10.6151
R652 B.n405 B.n56 10.6151
R653 B.n399 B.n56 10.6151
R654 B.n399 B.n398 10.6151
R655 B.n398 B.n397 10.6151
R656 B.n397 B.n58 10.6151
R657 B.n391 B.n390 10.6151
R658 B.n390 B.n389 10.6151
R659 B.n389 B.n63 10.6151
R660 B.n383 B.n63 10.6151
R661 B.n383 B.n382 10.6151
R662 B.n382 B.n381 10.6151
R663 B.n381 B.n65 10.6151
R664 B.n375 B.n65 10.6151
R665 B.n375 B.n374 10.6151
R666 B.n372 B.n69 10.6151
R667 B.n366 B.n69 10.6151
R668 B.n366 B.n365 10.6151
R669 B.n365 B.n364 10.6151
R670 B.n364 B.n71 10.6151
R671 B.n358 B.n71 10.6151
R672 B.n358 B.n357 10.6151
R673 B.n357 B.n356 10.6151
R674 B.n356 B.n73 10.6151
R675 B.n350 B.n73 10.6151
R676 B.n350 B.n349 10.6151
R677 B.n349 B.n348 10.6151
R678 B.n348 B.n75 10.6151
R679 B.n342 B.n75 10.6151
R680 B.n234 B.n233 10.6151
R681 B.n235 B.n234 10.6151
R682 B.n235 B.n115 10.6151
R683 B.n245 B.n115 10.6151
R684 B.n246 B.n245 10.6151
R685 B.n247 B.n246 10.6151
R686 B.n247 B.n107 10.6151
R687 B.n257 B.n107 10.6151
R688 B.n258 B.n257 10.6151
R689 B.n259 B.n258 10.6151
R690 B.n259 B.n99 10.6151
R691 B.n269 B.n99 10.6151
R692 B.n270 B.n269 10.6151
R693 B.n271 B.n270 10.6151
R694 B.n271 B.n92 10.6151
R695 B.n282 B.n92 10.6151
R696 B.n283 B.n282 10.6151
R697 B.n284 B.n283 10.6151
R698 B.n284 B.n83 10.6151
R699 B.n294 B.n83 10.6151
R700 B.n295 B.n294 10.6151
R701 B.n297 B.n295 10.6151
R702 B.n297 B.n296 10.6151
R703 B.n296 B.n76 10.6151
R704 B.n308 B.n76 10.6151
R705 B.n309 B.n308 10.6151
R706 B.n310 B.n309 10.6151
R707 B.n311 B.n310 10.6151
R708 B.n313 B.n311 10.6151
R709 B.n314 B.n313 10.6151
R710 B.n315 B.n314 10.6151
R711 B.n316 B.n315 10.6151
R712 B.n318 B.n316 10.6151
R713 B.n319 B.n318 10.6151
R714 B.n320 B.n319 10.6151
R715 B.n321 B.n320 10.6151
R716 B.n323 B.n321 10.6151
R717 B.n324 B.n323 10.6151
R718 B.n325 B.n324 10.6151
R719 B.n326 B.n325 10.6151
R720 B.n328 B.n326 10.6151
R721 B.n329 B.n328 10.6151
R722 B.n330 B.n329 10.6151
R723 B.n331 B.n330 10.6151
R724 B.n333 B.n331 10.6151
R725 B.n334 B.n333 10.6151
R726 B.n335 B.n334 10.6151
R727 B.n336 B.n335 10.6151
R728 B.n338 B.n336 10.6151
R729 B.n339 B.n338 10.6151
R730 B.n340 B.n339 10.6151
R731 B.n341 B.n340 10.6151
R732 B.n228 B.n227 10.6151
R733 B.n227 B.n127 10.6151
R734 B.n222 B.n127 10.6151
R735 B.n222 B.n221 10.6151
R736 B.n221 B.n129 10.6151
R737 B.n216 B.n129 10.6151
R738 B.n216 B.n215 10.6151
R739 B.n215 B.n214 10.6151
R740 B.n214 B.n131 10.6151
R741 B.n208 B.n131 10.6151
R742 B.n208 B.n207 10.6151
R743 B.n207 B.n206 10.6151
R744 B.n206 B.n133 10.6151
R745 B.n200 B.n133 10.6151
R746 B.n198 B.n197 10.6151
R747 B.n197 B.n137 10.6151
R748 B.n191 B.n137 10.6151
R749 B.n191 B.n190 10.6151
R750 B.n190 B.n189 10.6151
R751 B.n189 B.n139 10.6151
R752 B.n183 B.n139 10.6151
R753 B.n183 B.n182 10.6151
R754 B.n182 B.n181 10.6151
R755 B.n177 B.n176 10.6151
R756 B.n176 B.n145 10.6151
R757 B.n171 B.n145 10.6151
R758 B.n171 B.n170 10.6151
R759 B.n170 B.n169 10.6151
R760 B.n169 B.n147 10.6151
R761 B.n163 B.n147 10.6151
R762 B.n163 B.n162 10.6151
R763 B.n162 B.n161 10.6151
R764 B.n161 B.n149 10.6151
R765 B.n155 B.n149 10.6151
R766 B.n155 B.n154 10.6151
R767 B.n154 B.n153 10.6151
R768 B.n153 B.n123 10.6151
R769 B.n229 B.n119 10.6151
R770 B.n239 B.n119 10.6151
R771 B.n240 B.n239 10.6151
R772 B.n241 B.n240 10.6151
R773 B.n241 B.n111 10.6151
R774 B.n251 B.n111 10.6151
R775 B.n252 B.n251 10.6151
R776 B.n253 B.n252 10.6151
R777 B.n253 B.n103 10.6151
R778 B.n263 B.n103 10.6151
R779 B.n264 B.n263 10.6151
R780 B.n265 B.n264 10.6151
R781 B.n265 B.n95 10.6151
R782 B.n276 B.n95 10.6151
R783 B.n277 B.n276 10.6151
R784 B.n278 B.n277 10.6151
R785 B.n278 B.n88 10.6151
R786 B.n288 B.n88 10.6151
R787 B.n289 B.n288 10.6151
R788 B.n290 B.n289 10.6151
R789 B.n290 B.n80 10.6151
R790 B.n301 B.n80 10.6151
R791 B.n302 B.n301 10.6151
R792 B.n303 B.n302 10.6151
R793 B.n303 B.n0 10.6151
R794 B.n471 B.n1 10.6151
R795 B.n471 B.n470 10.6151
R796 B.n470 B.n469 10.6151
R797 B.n469 B.n10 10.6151
R798 B.n463 B.n10 10.6151
R799 B.n463 B.n462 10.6151
R800 B.n462 B.n461 10.6151
R801 B.n461 B.n17 10.6151
R802 B.n455 B.n17 10.6151
R803 B.n455 B.n454 10.6151
R804 B.n454 B.n453 10.6151
R805 B.n453 B.n23 10.6151
R806 B.n447 B.n23 10.6151
R807 B.n447 B.n446 10.6151
R808 B.n446 B.n445 10.6151
R809 B.n445 B.n31 10.6151
R810 B.n439 B.n31 10.6151
R811 B.n439 B.n438 10.6151
R812 B.n438 B.n437 10.6151
R813 B.n437 B.n38 10.6151
R814 B.n431 B.n38 10.6151
R815 B.n431 B.n430 10.6151
R816 B.n430 B.n429 10.6151
R817 B.n429 B.n45 10.6151
R818 B.n423 B.n45 10.6151
R819 B.n62 B.n58 9.36635
R820 B.n373 B.n372 9.36635
R821 B.n200 B.n199 9.36635
R822 B.n177 B.n143 9.36635
R823 B.n477 B.n0 2.81026
R824 B.n477 B.n1 2.81026
R825 B.n391 B.n62 1.24928
R826 B.n374 B.n373 1.24928
R827 B.n199 B.n198 1.24928
R828 B.n181 B.n143 1.24928
R829 VN.n0 VN.t2 77.6359
R830 VN.n1 VN.t3 77.6359
R831 VN.n0 VN.t0 77.214
R832 VN.n1 VN.t1 77.214
R833 VN VN.n1 46.4938
R834 VN VN.n0 9.54306
R835 VTAIL.n6 VTAIL.t0 69.6943
R836 VTAIL.n5 VTAIL.t3 69.6943
R837 VTAIL.n4 VTAIL.t5 69.6943
R838 VTAIL.n3 VTAIL.t7 69.6943
R839 VTAIL.n7 VTAIL.t4 69.6942
R840 VTAIL.n0 VTAIL.t6 69.6942
R841 VTAIL.n1 VTAIL.t2 69.6942
R842 VTAIL.n2 VTAIL.t1 69.6942
R843 VTAIL.n7 VTAIL.n6 16.7031
R844 VTAIL.n3 VTAIL.n2 16.7031
R845 VTAIL.n4 VTAIL.n3 1.7505
R846 VTAIL.n6 VTAIL.n5 1.7505
R847 VTAIL.n2 VTAIL.n1 1.7505
R848 VTAIL VTAIL.n0 0.93369
R849 VTAIL VTAIL.n7 0.81731
R850 VTAIL.n5 VTAIL.n4 0.470328
R851 VTAIL.n1 VTAIL.n0 0.470328
R852 VDD2.n2 VDD2.n0 111.325
R853 VDD2.n2 VDD2.n1 79.7731
R854 VDD2.n1 VDD2.t2 6.6005
R855 VDD2.n1 VDD2.t0 6.6005
R856 VDD2.n0 VDD2.t1 6.6005
R857 VDD2.n0 VDD2.t3 6.6005
R858 VDD2 VDD2.n2 0.0586897
R859 VP.n5 VP.n4 185.155
R860 VP.n14 VP.n13 185.155
R861 VP.n12 VP.n0 161.3
R862 VP.n11 VP.n10 161.3
R863 VP.n9 VP.n1 161.3
R864 VP.n8 VP.n7 161.3
R865 VP.n6 VP.n2 161.3
R866 VP.n3 VP.t2 77.636
R867 VP.n3 VP.t1 77.214
R868 VP.n4 VP.n3 46.1131
R869 VP.n5 VP.t3 42.5299
R870 VP.n13 VP.t0 42.5299
R871 VP.n7 VP.n1 40.577
R872 VP.n11 VP.n1 40.577
R873 VP.n7 VP.n6 24.5923
R874 VP.n12 VP.n11 24.5923
R875 VP.n6 VP.n5 0.738255
R876 VP.n13 VP.n12 0.738255
R877 VP.n4 VP.n2 0.189894
R878 VP.n8 VP.n2 0.189894
R879 VP.n9 VP.n8 0.189894
R880 VP.n10 VP.n9 0.189894
R881 VP.n10 VP.n0 0.189894
R882 VP.n14 VP.n0 0.189894
R883 VP VP.n14 0.0516364
R884 VDD1 VDD1.n1 111.849
R885 VDD1 VDD1.n0 79.8313
R886 VDD1.n0 VDD1.t1 6.6005
R887 VDD1.n0 VDD1.t2 6.6005
R888 VDD1.n1 VDD1.t0 6.6005
R889 VDD1.n1 VDD1.t3 6.6005
C0 VTAIL VP 1.60737f
C1 VDD1 VN 0.153244f
C2 VDD2 VP 0.342644f
C3 VDD2 VTAIL 2.93385f
C4 VN VP 3.8816f
C5 VDD1 VP 1.50807f
C6 VTAIL VN 1.59326f
C7 VDD2 VN 1.31977f
C8 VDD1 VTAIL 2.88568f
C9 VDD2 VDD1 0.806986f
C10 VDD2 B 2.499174f
C11 VDD1 B 4.50146f
C12 VTAIL B 3.941264f
C13 VN B 7.45581f
C14 VP B 6.243327f
C15 VDD1.t1 B 0.043541f
C16 VDD1.t2 B 0.043541f
C17 VDD1.n0 B 0.314203f
C18 VDD1.t0 B 0.043541f
C19 VDD1.t3 B 0.043541f
C20 VDD1.n1 B 0.526479f
C21 VP.n0 B 0.0224f
C22 VP.t0 B 0.284588f
C23 VP.n1 B 0.018092f
C24 VP.n2 B 0.0224f
C25 VP.t3 B 0.284588f
C26 VP.t2 B 0.388752f
C27 VP.t1 B 0.3875f
C28 VP.n3 B 0.982981f
C29 VP.n4 B 0.935369f
C30 VP.n5 B 0.171097f
C31 VP.n6 B 0.021648f
C32 VP.n7 B 0.044286f
C33 VP.n8 B 0.0224f
C34 VP.n9 B 0.0224f
C35 VP.n10 B 0.0224f
C36 VP.n11 B 0.044286f
C37 VP.n12 B 0.021648f
C38 VP.n13 B 0.171097f
C39 VP.n14 B 0.023847f
C40 VDD2.t1 B 0.044583f
C41 VDD2.t3 B 0.044583f
C42 VDD2.n0 B 0.525649f
C43 VDD2.t2 B 0.044583f
C44 VDD2.t0 B 0.044583f
C45 VDD2.n1 B 0.321533f
C46 VDD2.n2 B 1.76439f
C47 VTAIL.t6 B 0.283277f
C48 VTAIL.n0 B 0.216476f
C49 VTAIL.t2 B 0.283277f
C50 VTAIL.n1 B 0.25435f
C51 VTAIL.t1 B 0.283277f
C52 VTAIL.n2 B 0.629096f
C53 VTAIL.t7 B 0.283279f
C54 VTAIL.n3 B 0.629095f
C55 VTAIL.t5 B 0.283279f
C56 VTAIL.n4 B 0.254348f
C57 VTAIL.t3 B 0.283279f
C58 VTAIL.n5 B 0.254348f
C59 VTAIL.t0 B 0.283279f
C60 VTAIL.n6 B 0.629095f
C61 VTAIL.t4 B 0.283277f
C62 VTAIL.n7 B 0.585826f
C63 VN.t2 B 0.385638f
C64 VN.t0 B 0.384396f
C65 VN.n0 B 0.288026f
C66 VN.t3 B 0.385638f
C67 VN.t1 B 0.384396f
C68 VN.n1 B 0.988284f
.ends

