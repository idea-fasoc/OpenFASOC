* NGSPICE file created from diff_pair_sample_1726.ext - technology: sky130A

.subckt diff_pair_sample_1726 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t5 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=4.9803 ps=26.32 w=12.77 l=2.35
X1 B.t11 B.t9 B.t10 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=0 ps=0 w=12.77 l=2.35
X2 VDD1.t4 VP.t1 VTAIL.t6 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=2.10705 ps=13.1 w=12.77 l=2.35
X3 VTAIL.t11 VN.t0 VDD2.t5 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=2.10705 ps=13.1 w=12.77 l=2.35
X4 VDD1.t3 VP.t2 VTAIL.t8 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=4.9803 ps=26.32 w=12.77 l=2.35
X5 VTAIL.t7 VP.t3 VDD1.t2 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=2.10705 ps=13.1 w=12.77 l=2.35
X6 VTAIL.t10 VP.t4 VDD1.t1 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=2.10705 ps=13.1 w=12.77 l=2.35
X7 VDD2.t4 VN.t1 VTAIL.t3 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=2.10705 ps=13.1 w=12.77 l=2.35
X8 VDD2.t3 VN.t2 VTAIL.t2 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=4.9803 ps=26.32 w=12.77 l=2.35
X9 B.t8 B.t6 B.t7 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=0 ps=0 w=12.77 l=2.35
X10 VDD2.t2 VN.t3 VTAIL.t1 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=4.9803 ps=26.32 w=12.77 l=2.35
X11 VDD1.t0 VP.t5 VTAIL.t9 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=2.10705 ps=13.1 w=12.77 l=2.35
X12 B.t5 B.t3 B.t4 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=0 ps=0 w=12.77 l=2.35
X13 B.t2 B.t0 B.t1 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=0 ps=0 w=12.77 l=2.35
X14 VTAIL.t0 VN.t4 VDD2.t1 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=2.10705 pd=13.1 as=2.10705 ps=13.1 w=12.77 l=2.35
X15 VDD2.t0 VN.t5 VTAIL.t4 w_n3114_n3522# sky130_fd_pr__pfet_01v8 ad=4.9803 pd=26.32 as=2.10705 ps=13.1 w=12.77 l=2.35
R0 VP.n9 VP.t5 164.249
R1 VP.n11 VP.n8 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n14 VP.n7 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n6 161.3
R6 VP.n37 VP.n0 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n34 VP.n1 161.3
R9 VP.n33 VP.n32 161.3
R10 VP.n31 VP.n2 161.3
R11 VP.n30 VP.n29 161.3
R12 VP.n28 VP.n3 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n25 VP.n4 161.3
R15 VP.n24 VP.n23 161.3
R16 VP.n22 VP.n5 161.3
R17 VP.n30 VP.t3 130.96
R18 VP.n20 VP.t1 130.96
R19 VP.n38 VP.t2 130.96
R20 VP.n10 VP.t4 130.96
R21 VP.n18 VP.t0 130.96
R22 VP.n21 VP.n20 101.948
R23 VP.n39 VP.n38 101.948
R24 VP.n19 VP.n18 101.948
R25 VP.n26 VP.n25 56.0336
R26 VP.n32 VP.n1 56.0336
R27 VP.n12 VP.n7 56.0336
R28 VP.n21 VP.n19 48.2193
R29 VP.n10 VP.n9 47.8966
R30 VP.n25 VP.n24 24.9531
R31 VP.n36 VP.n1 24.9531
R32 VP.n16 VP.n7 24.9531
R33 VP.n24 VP.n5 24.4675
R34 VP.n26 VP.n3 24.4675
R35 VP.n30 VP.n3 24.4675
R36 VP.n31 VP.n30 24.4675
R37 VP.n32 VP.n31 24.4675
R38 VP.n37 VP.n36 24.4675
R39 VP.n17 VP.n16 24.4675
R40 VP.n11 VP.n10 24.4675
R41 VP.n12 VP.n11 24.4675
R42 VP.n20 VP.n5 8.80862
R43 VP.n38 VP.n37 8.80862
R44 VP.n18 VP.n17 8.80862
R45 VP.n9 VP.n8 6.92221
R46 VP.n19 VP.n6 0.278367
R47 VP.n22 VP.n21 0.278367
R48 VP.n39 VP.n0 0.278367
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153454
R64 VTAIL.n282 VTAIL.n218 756.745
R65 VTAIL.n66 VTAIL.n2 756.745
R66 VTAIL.n212 VTAIL.n148 756.745
R67 VTAIL.n140 VTAIL.n76 756.745
R68 VTAIL.n241 VTAIL.n240 585
R69 VTAIL.n238 VTAIL.n237 585
R70 VTAIL.n247 VTAIL.n246 585
R71 VTAIL.n249 VTAIL.n248 585
R72 VTAIL.n234 VTAIL.n233 585
R73 VTAIL.n255 VTAIL.n254 585
R74 VTAIL.n258 VTAIL.n257 585
R75 VTAIL.n256 VTAIL.n230 585
R76 VTAIL.n263 VTAIL.n229 585
R77 VTAIL.n265 VTAIL.n264 585
R78 VTAIL.n267 VTAIL.n266 585
R79 VTAIL.n226 VTAIL.n225 585
R80 VTAIL.n273 VTAIL.n272 585
R81 VTAIL.n275 VTAIL.n274 585
R82 VTAIL.n222 VTAIL.n221 585
R83 VTAIL.n281 VTAIL.n280 585
R84 VTAIL.n283 VTAIL.n282 585
R85 VTAIL.n25 VTAIL.n24 585
R86 VTAIL.n22 VTAIL.n21 585
R87 VTAIL.n31 VTAIL.n30 585
R88 VTAIL.n33 VTAIL.n32 585
R89 VTAIL.n18 VTAIL.n17 585
R90 VTAIL.n39 VTAIL.n38 585
R91 VTAIL.n42 VTAIL.n41 585
R92 VTAIL.n40 VTAIL.n14 585
R93 VTAIL.n47 VTAIL.n13 585
R94 VTAIL.n49 VTAIL.n48 585
R95 VTAIL.n51 VTAIL.n50 585
R96 VTAIL.n10 VTAIL.n9 585
R97 VTAIL.n57 VTAIL.n56 585
R98 VTAIL.n59 VTAIL.n58 585
R99 VTAIL.n6 VTAIL.n5 585
R100 VTAIL.n65 VTAIL.n64 585
R101 VTAIL.n67 VTAIL.n66 585
R102 VTAIL.n213 VTAIL.n212 585
R103 VTAIL.n211 VTAIL.n210 585
R104 VTAIL.n152 VTAIL.n151 585
R105 VTAIL.n205 VTAIL.n204 585
R106 VTAIL.n203 VTAIL.n202 585
R107 VTAIL.n156 VTAIL.n155 585
R108 VTAIL.n197 VTAIL.n196 585
R109 VTAIL.n195 VTAIL.n194 585
R110 VTAIL.n193 VTAIL.n159 585
R111 VTAIL.n163 VTAIL.n160 585
R112 VTAIL.n188 VTAIL.n187 585
R113 VTAIL.n186 VTAIL.n185 585
R114 VTAIL.n165 VTAIL.n164 585
R115 VTAIL.n180 VTAIL.n179 585
R116 VTAIL.n178 VTAIL.n177 585
R117 VTAIL.n169 VTAIL.n168 585
R118 VTAIL.n172 VTAIL.n171 585
R119 VTAIL.n141 VTAIL.n140 585
R120 VTAIL.n139 VTAIL.n138 585
R121 VTAIL.n80 VTAIL.n79 585
R122 VTAIL.n133 VTAIL.n132 585
R123 VTAIL.n131 VTAIL.n130 585
R124 VTAIL.n84 VTAIL.n83 585
R125 VTAIL.n125 VTAIL.n124 585
R126 VTAIL.n123 VTAIL.n122 585
R127 VTAIL.n121 VTAIL.n87 585
R128 VTAIL.n91 VTAIL.n88 585
R129 VTAIL.n116 VTAIL.n115 585
R130 VTAIL.n114 VTAIL.n113 585
R131 VTAIL.n93 VTAIL.n92 585
R132 VTAIL.n108 VTAIL.n107 585
R133 VTAIL.n106 VTAIL.n105 585
R134 VTAIL.n97 VTAIL.n96 585
R135 VTAIL.n100 VTAIL.n99 585
R136 VTAIL.t1 VTAIL.n239 329.036
R137 VTAIL.t8 VTAIL.n23 329.036
R138 VTAIL.t5 VTAIL.n170 329.036
R139 VTAIL.t2 VTAIL.n98 329.036
R140 VTAIL.n240 VTAIL.n237 171.744
R141 VTAIL.n247 VTAIL.n237 171.744
R142 VTAIL.n248 VTAIL.n247 171.744
R143 VTAIL.n248 VTAIL.n233 171.744
R144 VTAIL.n255 VTAIL.n233 171.744
R145 VTAIL.n257 VTAIL.n255 171.744
R146 VTAIL.n257 VTAIL.n256 171.744
R147 VTAIL.n256 VTAIL.n229 171.744
R148 VTAIL.n265 VTAIL.n229 171.744
R149 VTAIL.n266 VTAIL.n265 171.744
R150 VTAIL.n266 VTAIL.n225 171.744
R151 VTAIL.n273 VTAIL.n225 171.744
R152 VTAIL.n274 VTAIL.n273 171.744
R153 VTAIL.n274 VTAIL.n221 171.744
R154 VTAIL.n281 VTAIL.n221 171.744
R155 VTAIL.n282 VTAIL.n281 171.744
R156 VTAIL.n24 VTAIL.n21 171.744
R157 VTAIL.n31 VTAIL.n21 171.744
R158 VTAIL.n32 VTAIL.n31 171.744
R159 VTAIL.n32 VTAIL.n17 171.744
R160 VTAIL.n39 VTAIL.n17 171.744
R161 VTAIL.n41 VTAIL.n39 171.744
R162 VTAIL.n41 VTAIL.n40 171.744
R163 VTAIL.n40 VTAIL.n13 171.744
R164 VTAIL.n49 VTAIL.n13 171.744
R165 VTAIL.n50 VTAIL.n49 171.744
R166 VTAIL.n50 VTAIL.n9 171.744
R167 VTAIL.n57 VTAIL.n9 171.744
R168 VTAIL.n58 VTAIL.n57 171.744
R169 VTAIL.n58 VTAIL.n5 171.744
R170 VTAIL.n65 VTAIL.n5 171.744
R171 VTAIL.n66 VTAIL.n65 171.744
R172 VTAIL.n212 VTAIL.n211 171.744
R173 VTAIL.n211 VTAIL.n151 171.744
R174 VTAIL.n204 VTAIL.n151 171.744
R175 VTAIL.n204 VTAIL.n203 171.744
R176 VTAIL.n203 VTAIL.n155 171.744
R177 VTAIL.n196 VTAIL.n155 171.744
R178 VTAIL.n196 VTAIL.n195 171.744
R179 VTAIL.n195 VTAIL.n159 171.744
R180 VTAIL.n163 VTAIL.n159 171.744
R181 VTAIL.n187 VTAIL.n163 171.744
R182 VTAIL.n187 VTAIL.n186 171.744
R183 VTAIL.n186 VTAIL.n164 171.744
R184 VTAIL.n179 VTAIL.n164 171.744
R185 VTAIL.n179 VTAIL.n178 171.744
R186 VTAIL.n178 VTAIL.n168 171.744
R187 VTAIL.n171 VTAIL.n168 171.744
R188 VTAIL.n140 VTAIL.n139 171.744
R189 VTAIL.n139 VTAIL.n79 171.744
R190 VTAIL.n132 VTAIL.n79 171.744
R191 VTAIL.n132 VTAIL.n131 171.744
R192 VTAIL.n131 VTAIL.n83 171.744
R193 VTAIL.n124 VTAIL.n83 171.744
R194 VTAIL.n124 VTAIL.n123 171.744
R195 VTAIL.n123 VTAIL.n87 171.744
R196 VTAIL.n91 VTAIL.n87 171.744
R197 VTAIL.n115 VTAIL.n91 171.744
R198 VTAIL.n115 VTAIL.n114 171.744
R199 VTAIL.n114 VTAIL.n92 171.744
R200 VTAIL.n107 VTAIL.n92 171.744
R201 VTAIL.n107 VTAIL.n106 171.744
R202 VTAIL.n106 VTAIL.n96 171.744
R203 VTAIL.n99 VTAIL.n96 171.744
R204 VTAIL.n240 VTAIL.t1 85.8723
R205 VTAIL.n24 VTAIL.t8 85.8723
R206 VTAIL.n171 VTAIL.t5 85.8723
R207 VTAIL.n99 VTAIL.t2 85.8723
R208 VTAIL.n1 VTAIL.n0 54.975
R209 VTAIL.n73 VTAIL.n72 54.975
R210 VTAIL.n147 VTAIL.n146 54.975
R211 VTAIL.n75 VTAIL.n74 54.975
R212 VTAIL.n287 VTAIL.n286 30.8278
R213 VTAIL.n71 VTAIL.n70 30.8278
R214 VTAIL.n217 VTAIL.n216 30.8278
R215 VTAIL.n145 VTAIL.n144 30.8278
R216 VTAIL.n75 VTAIL.n73 27.9962
R217 VTAIL.n287 VTAIL.n217 25.6858
R218 VTAIL.n264 VTAIL.n263 13.1884
R219 VTAIL.n48 VTAIL.n47 13.1884
R220 VTAIL.n194 VTAIL.n193 13.1884
R221 VTAIL.n122 VTAIL.n121 13.1884
R222 VTAIL.n262 VTAIL.n230 12.8005
R223 VTAIL.n267 VTAIL.n228 12.8005
R224 VTAIL.n46 VTAIL.n14 12.8005
R225 VTAIL.n51 VTAIL.n12 12.8005
R226 VTAIL.n197 VTAIL.n158 12.8005
R227 VTAIL.n192 VTAIL.n160 12.8005
R228 VTAIL.n125 VTAIL.n86 12.8005
R229 VTAIL.n120 VTAIL.n88 12.8005
R230 VTAIL.n259 VTAIL.n258 12.0247
R231 VTAIL.n268 VTAIL.n226 12.0247
R232 VTAIL.n43 VTAIL.n42 12.0247
R233 VTAIL.n52 VTAIL.n10 12.0247
R234 VTAIL.n198 VTAIL.n156 12.0247
R235 VTAIL.n189 VTAIL.n188 12.0247
R236 VTAIL.n126 VTAIL.n84 12.0247
R237 VTAIL.n117 VTAIL.n116 12.0247
R238 VTAIL.n254 VTAIL.n232 11.249
R239 VTAIL.n272 VTAIL.n271 11.249
R240 VTAIL.n38 VTAIL.n16 11.249
R241 VTAIL.n56 VTAIL.n55 11.249
R242 VTAIL.n202 VTAIL.n201 11.249
R243 VTAIL.n185 VTAIL.n162 11.249
R244 VTAIL.n130 VTAIL.n129 11.249
R245 VTAIL.n113 VTAIL.n90 11.249
R246 VTAIL.n241 VTAIL.n239 10.7239
R247 VTAIL.n25 VTAIL.n23 10.7239
R248 VTAIL.n172 VTAIL.n170 10.7239
R249 VTAIL.n100 VTAIL.n98 10.7239
R250 VTAIL.n253 VTAIL.n234 10.4732
R251 VTAIL.n275 VTAIL.n224 10.4732
R252 VTAIL.n37 VTAIL.n18 10.4732
R253 VTAIL.n59 VTAIL.n8 10.4732
R254 VTAIL.n205 VTAIL.n154 10.4732
R255 VTAIL.n184 VTAIL.n165 10.4732
R256 VTAIL.n133 VTAIL.n82 10.4732
R257 VTAIL.n112 VTAIL.n93 10.4732
R258 VTAIL.n250 VTAIL.n249 9.69747
R259 VTAIL.n276 VTAIL.n222 9.69747
R260 VTAIL.n34 VTAIL.n33 9.69747
R261 VTAIL.n60 VTAIL.n6 9.69747
R262 VTAIL.n206 VTAIL.n152 9.69747
R263 VTAIL.n181 VTAIL.n180 9.69747
R264 VTAIL.n134 VTAIL.n80 9.69747
R265 VTAIL.n109 VTAIL.n108 9.69747
R266 VTAIL.n286 VTAIL.n285 9.45567
R267 VTAIL.n70 VTAIL.n69 9.45567
R268 VTAIL.n216 VTAIL.n215 9.45567
R269 VTAIL.n144 VTAIL.n143 9.45567
R270 VTAIL.n220 VTAIL.n219 9.3005
R271 VTAIL.n279 VTAIL.n278 9.3005
R272 VTAIL.n277 VTAIL.n276 9.3005
R273 VTAIL.n224 VTAIL.n223 9.3005
R274 VTAIL.n271 VTAIL.n270 9.3005
R275 VTAIL.n269 VTAIL.n268 9.3005
R276 VTAIL.n228 VTAIL.n227 9.3005
R277 VTAIL.n243 VTAIL.n242 9.3005
R278 VTAIL.n245 VTAIL.n244 9.3005
R279 VTAIL.n236 VTAIL.n235 9.3005
R280 VTAIL.n251 VTAIL.n250 9.3005
R281 VTAIL.n253 VTAIL.n252 9.3005
R282 VTAIL.n232 VTAIL.n231 9.3005
R283 VTAIL.n260 VTAIL.n259 9.3005
R284 VTAIL.n262 VTAIL.n261 9.3005
R285 VTAIL.n285 VTAIL.n284 9.3005
R286 VTAIL.n4 VTAIL.n3 9.3005
R287 VTAIL.n63 VTAIL.n62 9.3005
R288 VTAIL.n61 VTAIL.n60 9.3005
R289 VTAIL.n8 VTAIL.n7 9.3005
R290 VTAIL.n55 VTAIL.n54 9.3005
R291 VTAIL.n53 VTAIL.n52 9.3005
R292 VTAIL.n12 VTAIL.n11 9.3005
R293 VTAIL.n27 VTAIL.n26 9.3005
R294 VTAIL.n29 VTAIL.n28 9.3005
R295 VTAIL.n20 VTAIL.n19 9.3005
R296 VTAIL.n35 VTAIL.n34 9.3005
R297 VTAIL.n37 VTAIL.n36 9.3005
R298 VTAIL.n16 VTAIL.n15 9.3005
R299 VTAIL.n44 VTAIL.n43 9.3005
R300 VTAIL.n46 VTAIL.n45 9.3005
R301 VTAIL.n69 VTAIL.n68 9.3005
R302 VTAIL.n174 VTAIL.n173 9.3005
R303 VTAIL.n176 VTAIL.n175 9.3005
R304 VTAIL.n167 VTAIL.n166 9.3005
R305 VTAIL.n182 VTAIL.n181 9.3005
R306 VTAIL.n184 VTAIL.n183 9.3005
R307 VTAIL.n162 VTAIL.n161 9.3005
R308 VTAIL.n190 VTAIL.n189 9.3005
R309 VTAIL.n192 VTAIL.n191 9.3005
R310 VTAIL.n215 VTAIL.n214 9.3005
R311 VTAIL.n150 VTAIL.n149 9.3005
R312 VTAIL.n209 VTAIL.n208 9.3005
R313 VTAIL.n207 VTAIL.n206 9.3005
R314 VTAIL.n154 VTAIL.n153 9.3005
R315 VTAIL.n201 VTAIL.n200 9.3005
R316 VTAIL.n199 VTAIL.n198 9.3005
R317 VTAIL.n158 VTAIL.n157 9.3005
R318 VTAIL.n102 VTAIL.n101 9.3005
R319 VTAIL.n104 VTAIL.n103 9.3005
R320 VTAIL.n95 VTAIL.n94 9.3005
R321 VTAIL.n110 VTAIL.n109 9.3005
R322 VTAIL.n112 VTAIL.n111 9.3005
R323 VTAIL.n90 VTAIL.n89 9.3005
R324 VTAIL.n118 VTAIL.n117 9.3005
R325 VTAIL.n120 VTAIL.n119 9.3005
R326 VTAIL.n143 VTAIL.n142 9.3005
R327 VTAIL.n78 VTAIL.n77 9.3005
R328 VTAIL.n137 VTAIL.n136 9.3005
R329 VTAIL.n135 VTAIL.n134 9.3005
R330 VTAIL.n82 VTAIL.n81 9.3005
R331 VTAIL.n129 VTAIL.n128 9.3005
R332 VTAIL.n127 VTAIL.n126 9.3005
R333 VTAIL.n86 VTAIL.n85 9.3005
R334 VTAIL.n246 VTAIL.n236 8.92171
R335 VTAIL.n280 VTAIL.n279 8.92171
R336 VTAIL.n30 VTAIL.n20 8.92171
R337 VTAIL.n64 VTAIL.n63 8.92171
R338 VTAIL.n210 VTAIL.n209 8.92171
R339 VTAIL.n177 VTAIL.n167 8.92171
R340 VTAIL.n138 VTAIL.n137 8.92171
R341 VTAIL.n105 VTAIL.n95 8.92171
R342 VTAIL.n245 VTAIL.n238 8.14595
R343 VTAIL.n283 VTAIL.n220 8.14595
R344 VTAIL.n29 VTAIL.n22 8.14595
R345 VTAIL.n67 VTAIL.n4 8.14595
R346 VTAIL.n213 VTAIL.n150 8.14595
R347 VTAIL.n176 VTAIL.n169 8.14595
R348 VTAIL.n141 VTAIL.n78 8.14595
R349 VTAIL.n104 VTAIL.n97 8.14595
R350 VTAIL.n242 VTAIL.n241 7.3702
R351 VTAIL.n284 VTAIL.n218 7.3702
R352 VTAIL.n26 VTAIL.n25 7.3702
R353 VTAIL.n68 VTAIL.n2 7.3702
R354 VTAIL.n214 VTAIL.n148 7.3702
R355 VTAIL.n173 VTAIL.n172 7.3702
R356 VTAIL.n142 VTAIL.n76 7.3702
R357 VTAIL.n101 VTAIL.n100 7.3702
R358 VTAIL.n286 VTAIL.n218 6.59444
R359 VTAIL.n70 VTAIL.n2 6.59444
R360 VTAIL.n216 VTAIL.n148 6.59444
R361 VTAIL.n144 VTAIL.n76 6.59444
R362 VTAIL.n242 VTAIL.n238 5.81868
R363 VTAIL.n284 VTAIL.n283 5.81868
R364 VTAIL.n26 VTAIL.n22 5.81868
R365 VTAIL.n68 VTAIL.n67 5.81868
R366 VTAIL.n214 VTAIL.n213 5.81868
R367 VTAIL.n173 VTAIL.n169 5.81868
R368 VTAIL.n142 VTAIL.n141 5.81868
R369 VTAIL.n101 VTAIL.n97 5.81868
R370 VTAIL.n246 VTAIL.n245 5.04292
R371 VTAIL.n280 VTAIL.n220 5.04292
R372 VTAIL.n30 VTAIL.n29 5.04292
R373 VTAIL.n64 VTAIL.n4 5.04292
R374 VTAIL.n210 VTAIL.n150 5.04292
R375 VTAIL.n177 VTAIL.n176 5.04292
R376 VTAIL.n138 VTAIL.n78 5.04292
R377 VTAIL.n105 VTAIL.n104 5.04292
R378 VTAIL.n249 VTAIL.n236 4.26717
R379 VTAIL.n279 VTAIL.n222 4.26717
R380 VTAIL.n33 VTAIL.n20 4.26717
R381 VTAIL.n63 VTAIL.n6 4.26717
R382 VTAIL.n209 VTAIL.n152 4.26717
R383 VTAIL.n180 VTAIL.n167 4.26717
R384 VTAIL.n137 VTAIL.n80 4.26717
R385 VTAIL.n108 VTAIL.n95 4.26717
R386 VTAIL.n250 VTAIL.n234 3.49141
R387 VTAIL.n276 VTAIL.n275 3.49141
R388 VTAIL.n34 VTAIL.n18 3.49141
R389 VTAIL.n60 VTAIL.n59 3.49141
R390 VTAIL.n206 VTAIL.n205 3.49141
R391 VTAIL.n181 VTAIL.n165 3.49141
R392 VTAIL.n134 VTAIL.n133 3.49141
R393 VTAIL.n109 VTAIL.n93 3.49141
R394 VTAIL.n254 VTAIL.n253 2.71565
R395 VTAIL.n272 VTAIL.n224 2.71565
R396 VTAIL.n38 VTAIL.n37 2.71565
R397 VTAIL.n56 VTAIL.n8 2.71565
R398 VTAIL.n202 VTAIL.n154 2.71565
R399 VTAIL.n185 VTAIL.n184 2.71565
R400 VTAIL.n130 VTAIL.n82 2.71565
R401 VTAIL.n113 VTAIL.n112 2.71565
R402 VTAIL.n0 VTAIL.t4 2.54592
R403 VTAIL.n0 VTAIL.t0 2.54592
R404 VTAIL.n72 VTAIL.t6 2.54592
R405 VTAIL.n72 VTAIL.t7 2.54592
R406 VTAIL.n146 VTAIL.t9 2.54592
R407 VTAIL.n146 VTAIL.t10 2.54592
R408 VTAIL.n74 VTAIL.t3 2.54592
R409 VTAIL.n74 VTAIL.t11 2.54592
R410 VTAIL.n243 VTAIL.n239 2.41282
R411 VTAIL.n27 VTAIL.n23 2.41282
R412 VTAIL.n174 VTAIL.n170 2.41282
R413 VTAIL.n102 VTAIL.n98 2.41282
R414 VTAIL.n145 VTAIL.n75 2.31084
R415 VTAIL.n217 VTAIL.n147 2.31084
R416 VTAIL.n73 VTAIL.n71 2.31084
R417 VTAIL.n258 VTAIL.n232 1.93989
R418 VTAIL.n271 VTAIL.n226 1.93989
R419 VTAIL.n42 VTAIL.n16 1.93989
R420 VTAIL.n55 VTAIL.n10 1.93989
R421 VTAIL.n201 VTAIL.n156 1.93989
R422 VTAIL.n188 VTAIL.n162 1.93989
R423 VTAIL.n129 VTAIL.n84 1.93989
R424 VTAIL.n116 VTAIL.n90 1.93989
R425 VTAIL VTAIL.n287 1.67507
R426 VTAIL.n147 VTAIL.n145 1.6255
R427 VTAIL.n71 VTAIL.n1 1.6255
R428 VTAIL.n259 VTAIL.n230 1.16414
R429 VTAIL.n268 VTAIL.n267 1.16414
R430 VTAIL.n43 VTAIL.n14 1.16414
R431 VTAIL.n52 VTAIL.n51 1.16414
R432 VTAIL.n198 VTAIL.n197 1.16414
R433 VTAIL.n189 VTAIL.n160 1.16414
R434 VTAIL.n126 VTAIL.n125 1.16414
R435 VTAIL.n117 VTAIL.n88 1.16414
R436 VTAIL VTAIL.n1 0.636276
R437 VTAIL.n263 VTAIL.n262 0.388379
R438 VTAIL.n264 VTAIL.n228 0.388379
R439 VTAIL.n47 VTAIL.n46 0.388379
R440 VTAIL.n48 VTAIL.n12 0.388379
R441 VTAIL.n194 VTAIL.n158 0.388379
R442 VTAIL.n193 VTAIL.n192 0.388379
R443 VTAIL.n122 VTAIL.n86 0.388379
R444 VTAIL.n121 VTAIL.n120 0.388379
R445 VTAIL.n244 VTAIL.n243 0.155672
R446 VTAIL.n244 VTAIL.n235 0.155672
R447 VTAIL.n251 VTAIL.n235 0.155672
R448 VTAIL.n252 VTAIL.n251 0.155672
R449 VTAIL.n252 VTAIL.n231 0.155672
R450 VTAIL.n260 VTAIL.n231 0.155672
R451 VTAIL.n261 VTAIL.n260 0.155672
R452 VTAIL.n261 VTAIL.n227 0.155672
R453 VTAIL.n269 VTAIL.n227 0.155672
R454 VTAIL.n270 VTAIL.n269 0.155672
R455 VTAIL.n270 VTAIL.n223 0.155672
R456 VTAIL.n277 VTAIL.n223 0.155672
R457 VTAIL.n278 VTAIL.n277 0.155672
R458 VTAIL.n278 VTAIL.n219 0.155672
R459 VTAIL.n285 VTAIL.n219 0.155672
R460 VTAIL.n28 VTAIL.n27 0.155672
R461 VTAIL.n28 VTAIL.n19 0.155672
R462 VTAIL.n35 VTAIL.n19 0.155672
R463 VTAIL.n36 VTAIL.n35 0.155672
R464 VTAIL.n36 VTAIL.n15 0.155672
R465 VTAIL.n44 VTAIL.n15 0.155672
R466 VTAIL.n45 VTAIL.n44 0.155672
R467 VTAIL.n45 VTAIL.n11 0.155672
R468 VTAIL.n53 VTAIL.n11 0.155672
R469 VTAIL.n54 VTAIL.n53 0.155672
R470 VTAIL.n54 VTAIL.n7 0.155672
R471 VTAIL.n61 VTAIL.n7 0.155672
R472 VTAIL.n62 VTAIL.n61 0.155672
R473 VTAIL.n62 VTAIL.n3 0.155672
R474 VTAIL.n69 VTAIL.n3 0.155672
R475 VTAIL.n215 VTAIL.n149 0.155672
R476 VTAIL.n208 VTAIL.n149 0.155672
R477 VTAIL.n208 VTAIL.n207 0.155672
R478 VTAIL.n207 VTAIL.n153 0.155672
R479 VTAIL.n200 VTAIL.n153 0.155672
R480 VTAIL.n200 VTAIL.n199 0.155672
R481 VTAIL.n199 VTAIL.n157 0.155672
R482 VTAIL.n191 VTAIL.n157 0.155672
R483 VTAIL.n191 VTAIL.n190 0.155672
R484 VTAIL.n190 VTAIL.n161 0.155672
R485 VTAIL.n183 VTAIL.n161 0.155672
R486 VTAIL.n183 VTAIL.n182 0.155672
R487 VTAIL.n182 VTAIL.n166 0.155672
R488 VTAIL.n175 VTAIL.n166 0.155672
R489 VTAIL.n175 VTAIL.n174 0.155672
R490 VTAIL.n143 VTAIL.n77 0.155672
R491 VTAIL.n136 VTAIL.n77 0.155672
R492 VTAIL.n136 VTAIL.n135 0.155672
R493 VTAIL.n135 VTAIL.n81 0.155672
R494 VTAIL.n128 VTAIL.n81 0.155672
R495 VTAIL.n128 VTAIL.n127 0.155672
R496 VTAIL.n127 VTAIL.n85 0.155672
R497 VTAIL.n119 VTAIL.n85 0.155672
R498 VTAIL.n119 VTAIL.n118 0.155672
R499 VTAIL.n118 VTAIL.n89 0.155672
R500 VTAIL.n111 VTAIL.n89 0.155672
R501 VTAIL.n111 VTAIL.n110 0.155672
R502 VTAIL.n110 VTAIL.n94 0.155672
R503 VTAIL.n103 VTAIL.n94 0.155672
R504 VTAIL.n103 VTAIL.n102 0.155672
R505 VDD1.n64 VDD1.n0 756.745
R506 VDD1.n133 VDD1.n69 756.745
R507 VDD1.n65 VDD1.n64 585
R508 VDD1.n63 VDD1.n62 585
R509 VDD1.n4 VDD1.n3 585
R510 VDD1.n57 VDD1.n56 585
R511 VDD1.n55 VDD1.n54 585
R512 VDD1.n8 VDD1.n7 585
R513 VDD1.n49 VDD1.n48 585
R514 VDD1.n47 VDD1.n46 585
R515 VDD1.n45 VDD1.n11 585
R516 VDD1.n15 VDD1.n12 585
R517 VDD1.n40 VDD1.n39 585
R518 VDD1.n38 VDD1.n37 585
R519 VDD1.n17 VDD1.n16 585
R520 VDD1.n32 VDD1.n31 585
R521 VDD1.n30 VDD1.n29 585
R522 VDD1.n21 VDD1.n20 585
R523 VDD1.n24 VDD1.n23 585
R524 VDD1.n92 VDD1.n91 585
R525 VDD1.n89 VDD1.n88 585
R526 VDD1.n98 VDD1.n97 585
R527 VDD1.n100 VDD1.n99 585
R528 VDD1.n85 VDD1.n84 585
R529 VDD1.n106 VDD1.n105 585
R530 VDD1.n109 VDD1.n108 585
R531 VDD1.n107 VDD1.n81 585
R532 VDD1.n114 VDD1.n80 585
R533 VDD1.n116 VDD1.n115 585
R534 VDD1.n118 VDD1.n117 585
R535 VDD1.n77 VDD1.n76 585
R536 VDD1.n124 VDD1.n123 585
R537 VDD1.n126 VDD1.n125 585
R538 VDD1.n73 VDD1.n72 585
R539 VDD1.n132 VDD1.n131 585
R540 VDD1.n134 VDD1.n133 585
R541 VDD1.t4 VDD1.n90 329.036
R542 VDD1.t0 VDD1.n22 329.036
R543 VDD1.n64 VDD1.n63 171.744
R544 VDD1.n63 VDD1.n3 171.744
R545 VDD1.n56 VDD1.n3 171.744
R546 VDD1.n56 VDD1.n55 171.744
R547 VDD1.n55 VDD1.n7 171.744
R548 VDD1.n48 VDD1.n7 171.744
R549 VDD1.n48 VDD1.n47 171.744
R550 VDD1.n47 VDD1.n11 171.744
R551 VDD1.n15 VDD1.n11 171.744
R552 VDD1.n39 VDD1.n15 171.744
R553 VDD1.n39 VDD1.n38 171.744
R554 VDD1.n38 VDD1.n16 171.744
R555 VDD1.n31 VDD1.n16 171.744
R556 VDD1.n31 VDD1.n30 171.744
R557 VDD1.n30 VDD1.n20 171.744
R558 VDD1.n23 VDD1.n20 171.744
R559 VDD1.n91 VDD1.n88 171.744
R560 VDD1.n98 VDD1.n88 171.744
R561 VDD1.n99 VDD1.n98 171.744
R562 VDD1.n99 VDD1.n84 171.744
R563 VDD1.n106 VDD1.n84 171.744
R564 VDD1.n108 VDD1.n106 171.744
R565 VDD1.n108 VDD1.n107 171.744
R566 VDD1.n107 VDD1.n80 171.744
R567 VDD1.n116 VDD1.n80 171.744
R568 VDD1.n117 VDD1.n116 171.744
R569 VDD1.n117 VDD1.n76 171.744
R570 VDD1.n124 VDD1.n76 171.744
R571 VDD1.n125 VDD1.n124 171.744
R572 VDD1.n125 VDD1.n72 171.744
R573 VDD1.n132 VDD1.n72 171.744
R574 VDD1.n133 VDD1.n132 171.744
R575 VDD1.n23 VDD1.t0 85.8723
R576 VDD1.n91 VDD1.t4 85.8723
R577 VDD1.n139 VDD1.n138 72.176
R578 VDD1.n141 VDD1.n140 71.6536
R579 VDD1 VDD1.n68 49.2975
R580 VDD1.n139 VDD1.n137 49.184
R581 VDD1.n141 VDD1.n139 43.9707
R582 VDD1.n46 VDD1.n45 13.1884
R583 VDD1.n115 VDD1.n114 13.1884
R584 VDD1.n49 VDD1.n10 12.8005
R585 VDD1.n44 VDD1.n12 12.8005
R586 VDD1.n113 VDD1.n81 12.8005
R587 VDD1.n118 VDD1.n79 12.8005
R588 VDD1.n50 VDD1.n8 12.0247
R589 VDD1.n41 VDD1.n40 12.0247
R590 VDD1.n110 VDD1.n109 12.0247
R591 VDD1.n119 VDD1.n77 12.0247
R592 VDD1.n54 VDD1.n53 11.249
R593 VDD1.n37 VDD1.n14 11.249
R594 VDD1.n105 VDD1.n83 11.249
R595 VDD1.n123 VDD1.n122 11.249
R596 VDD1.n24 VDD1.n22 10.7239
R597 VDD1.n92 VDD1.n90 10.7239
R598 VDD1.n57 VDD1.n6 10.4732
R599 VDD1.n36 VDD1.n17 10.4732
R600 VDD1.n104 VDD1.n85 10.4732
R601 VDD1.n126 VDD1.n75 10.4732
R602 VDD1.n58 VDD1.n4 9.69747
R603 VDD1.n33 VDD1.n32 9.69747
R604 VDD1.n101 VDD1.n100 9.69747
R605 VDD1.n127 VDD1.n73 9.69747
R606 VDD1.n68 VDD1.n67 9.45567
R607 VDD1.n137 VDD1.n136 9.45567
R608 VDD1.n26 VDD1.n25 9.3005
R609 VDD1.n28 VDD1.n27 9.3005
R610 VDD1.n19 VDD1.n18 9.3005
R611 VDD1.n34 VDD1.n33 9.3005
R612 VDD1.n36 VDD1.n35 9.3005
R613 VDD1.n14 VDD1.n13 9.3005
R614 VDD1.n42 VDD1.n41 9.3005
R615 VDD1.n44 VDD1.n43 9.3005
R616 VDD1.n67 VDD1.n66 9.3005
R617 VDD1.n2 VDD1.n1 9.3005
R618 VDD1.n61 VDD1.n60 9.3005
R619 VDD1.n59 VDD1.n58 9.3005
R620 VDD1.n6 VDD1.n5 9.3005
R621 VDD1.n53 VDD1.n52 9.3005
R622 VDD1.n51 VDD1.n50 9.3005
R623 VDD1.n10 VDD1.n9 9.3005
R624 VDD1.n71 VDD1.n70 9.3005
R625 VDD1.n130 VDD1.n129 9.3005
R626 VDD1.n128 VDD1.n127 9.3005
R627 VDD1.n75 VDD1.n74 9.3005
R628 VDD1.n122 VDD1.n121 9.3005
R629 VDD1.n120 VDD1.n119 9.3005
R630 VDD1.n79 VDD1.n78 9.3005
R631 VDD1.n94 VDD1.n93 9.3005
R632 VDD1.n96 VDD1.n95 9.3005
R633 VDD1.n87 VDD1.n86 9.3005
R634 VDD1.n102 VDD1.n101 9.3005
R635 VDD1.n104 VDD1.n103 9.3005
R636 VDD1.n83 VDD1.n82 9.3005
R637 VDD1.n111 VDD1.n110 9.3005
R638 VDD1.n113 VDD1.n112 9.3005
R639 VDD1.n136 VDD1.n135 9.3005
R640 VDD1.n62 VDD1.n61 8.92171
R641 VDD1.n29 VDD1.n19 8.92171
R642 VDD1.n97 VDD1.n87 8.92171
R643 VDD1.n131 VDD1.n130 8.92171
R644 VDD1.n65 VDD1.n2 8.14595
R645 VDD1.n28 VDD1.n21 8.14595
R646 VDD1.n96 VDD1.n89 8.14595
R647 VDD1.n134 VDD1.n71 8.14595
R648 VDD1.n66 VDD1.n0 7.3702
R649 VDD1.n25 VDD1.n24 7.3702
R650 VDD1.n93 VDD1.n92 7.3702
R651 VDD1.n135 VDD1.n69 7.3702
R652 VDD1.n68 VDD1.n0 6.59444
R653 VDD1.n137 VDD1.n69 6.59444
R654 VDD1.n66 VDD1.n65 5.81868
R655 VDD1.n25 VDD1.n21 5.81868
R656 VDD1.n93 VDD1.n89 5.81868
R657 VDD1.n135 VDD1.n134 5.81868
R658 VDD1.n62 VDD1.n2 5.04292
R659 VDD1.n29 VDD1.n28 5.04292
R660 VDD1.n97 VDD1.n96 5.04292
R661 VDD1.n131 VDD1.n71 5.04292
R662 VDD1.n61 VDD1.n4 4.26717
R663 VDD1.n32 VDD1.n19 4.26717
R664 VDD1.n100 VDD1.n87 4.26717
R665 VDD1.n130 VDD1.n73 4.26717
R666 VDD1.n58 VDD1.n57 3.49141
R667 VDD1.n33 VDD1.n17 3.49141
R668 VDD1.n101 VDD1.n85 3.49141
R669 VDD1.n127 VDD1.n126 3.49141
R670 VDD1.n54 VDD1.n6 2.71565
R671 VDD1.n37 VDD1.n36 2.71565
R672 VDD1.n105 VDD1.n104 2.71565
R673 VDD1.n123 VDD1.n75 2.71565
R674 VDD1.n140 VDD1.t1 2.54592
R675 VDD1.n140 VDD1.t5 2.54592
R676 VDD1.n138 VDD1.t2 2.54592
R677 VDD1.n138 VDD1.t3 2.54592
R678 VDD1.n26 VDD1.n22 2.41282
R679 VDD1.n94 VDD1.n90 2.41282
R680 VDD1.n53 VDD1.n8 1.93989
R681 VDD1.n40 VDD1.n14 1.93989
R682 VDD1.n109 VDD1.n83 1.93989
R683 VDD1.n122 VDD1.n77 1.93989
R684 VDD1.n50 VDD1.n49 1.16414
R685 VDD1.n41 VDD1.n12 1.16414
R686 VDD1.n110 VDD1.n81 1.16414
R687 VDD1.n119 VDD1.n118 1.16414
R688 VDD1 VDD1.n141 0.519897
R689 VDD1.n46 VDD1.n10 0.388379
R690 VDD1.n45 VDD1.n44 0.388379
R691 VDD1.n114 VDD1.n113 0.388379
R692 VDD1.n115 VDD1.n79 0.388379
R693 VDD1.n67 VDD1.n1 0.155672
R694 VDD1.n60 VDD1.n1 0.155672
R695 VDD1.n60 VDD1.n59 0.155672
R696 VDD1.n59 VDD1.n5 0.155672
R697 VDD1.n52 VDD1.n5 0.155672
R698 VDD1.n52 VDD1.n51 0.155672
R699 VDD1.n51 VDD1.n9 0.155672
R700 VDD1.n43 VDD1.n9 0.155672
R701 VDD1.n43 VDD1.n42 0.155672
R702 VDD1.n42 VDD1.n13 0.155672
R703 VDD1.n35 VDD1.n13 0.155672
R704 VDD1.n35 VDD1.n34 0.155672
R705 VDD1.n34 VDD1.n18 0.155672
R706 VDD1.n27 VDD1.n18 0.155672
R707 VDD1.n27 VDD1.n26 0.155672
R708 VDD1.n95 VDD1.n94 0.155672
R709 VDD1.n95 VDD1.n86 0.155672
R710 VDD1.n102 VDD1.n86 0.155672
R711 VDD1.n103 VDD1.n102 0.155672
R712 VDD1.n103 VDD1.n82 0.155672
R713 VDD1.n111 VDD1.n82 0.155672
R714 VDD1.n112 VDD1.n111 0.155672
R715 VDD1.n112 VDD1.n78 0.155672
R716 VDD1.n120 VDD1.n78 0.155672
R717 VDD1.n121 VDD1.n120 0.155672
R718 VDD1.n121 VDD1.n74 0.155672
R719 VDD1.n128 VDD1.n74 0.155672
R720 VDD1.n129 VDD1.n128 0.155672
R721 VDD1.n129 VDD1.n70 0.155672
R722 VDD1.n136 VDD1.n70 0.155672
R723 B.n390 B.n389 585
R724 B.n388 B.n115 585
R725 B.n387 B.n386 585
R726 B.n385 B.n116 585
R727 B.n384 B.n383 585
R728 B.n382 B.n117 585
R729 B.n381 B.n380 585
R730 B.n379 B.n118 585
R731 B.n378 B.n377 585
R732 B.n376 B.n119 585
R733 B.n375 B.n374 585
R734 B.n373 B.n120 585
R735 B.n372 B.n371 585
R736 B.n370 B.n121 585
R737 B.n369 B.n368 585
R738 B.n367 B.n122 585
R739 B.n366 B.n365 585
R740 B.n364 B.n123 585
R741 B.n363 B.n362 585
R742 B.n361 B.n124 585
R743 B.n360 B.n359 585
R744 B.n358 B.n125 585
R745 B.n357 B.n356 585
R746 B.n355 B.n126 585
R747 B.n354 B.n353 585
R748 B.n352 B.n127 585
R749 B.n351 B.n350 585
R750 B.n349 B.n128 585
R751 B.n348 B.n347 585
R752 B.n346 B.n129 585
R753 B.n345 B.n344 585
R754 B.n343 B.n130 585
R755 B.n342 B.n341 585
R756 B.n340 B.n131 585
R757 B.n339 B.n338 585
R758 B.n337 B.n132 585
R759 B.n336 B.n335 585
R760 B.n334 B.n133 585
R761 B.n333 B.n332 585
R762 B.n331 B.n134 585
R763 B.n330 B.n329 585
R764 B.n328 B.n135 585
R765 B.n327 B.n326 585
R766 B.n325 B.n136 585
R767 B.n324 B.n323 585
R768 B.n319 B.n137 585
R769 B.n318 B.n317 585
R770 B.n316 B.n138 585
R771 B.n315 B.n314 585
R772 B.n313 B.n139 585
R773 B.n312 B.n311 585
R774 B.n310 B.n140 585
R775 B.n309 B.n308 585
R776 B.n306 B.n141 585
R777 B.n305 B.n304 585
R778 B.n303 B.n144 585
R779 B.n302 B.n301 585
R780 B.n300 B.n145 585
R781 B.n299 B.n298 585
R782 B.n297 B.n146 585
R783 B.n296 B.n295 585
R784 B.n294 B.n147 585
R785 B.n293 B.n292 585
R786 B.n291 B.n148 585
R787 B.n290 B.n289 585
R788 B.n288 B.n149 585
R789 B.n287 B.n286 585
R790 B.n285 B.n150 585
R791 B.n284 B.n283 585
R792 B.n282 B.n151 585
R793 B.n281 B.n280 585
R794 B.n279 B.n152 585
R795 B.n278 B.n277 585
R796 B.n276 B.n153 585
R797 B.n275 B.n274 585
R798 B.n273 B.n154 585
R799 B.n272 B.n271 585
R800 B.n270 B.n155 585
R801 B.n269 B.n268 585
R802 B.n267 B.n156 585
R803 B.n266 B.n265 585
R804 B.n264 B.n157 585
R805 B.n263 B.n262 585
R806 B.n261 B.n158 585
R807 B.n260 B.n259 585
R808 B.n258 B.n159 585
R809 B.n257 B.n256 585
R810 B.n255 B.n160 585
R811 B.n254 B.n253 585
R812 B.n252 B.n161 585
R813 B.n251 B.n250 585
R814 B.n249 B.n162 585
R815 B.n248 B.n247 585
R816 B.n246 B.n163 585
R817 B.n245 B.n244 585
R818 B.n243 B.n164 585
R819 B.n242 B.n241 585
R820 B.n391 B.n114 585
R821 B.n393 B.n392 585
R822 B.n394 B.n113 585
R823 B.n396 B.n395 585
R824 B.n397 B.n112 585
R825 B.n399 B.n398 585
R826 B.n400 B.n111 585
R827 B.n402 B.n401 585
R828 B.n403 B.n110 585
R829 B.n405 B.n404 585
R830 B.n406 B.n109 585
R831 B.n408 B.n407 585
R832 B.n409 B.n108 585
R833 B.n411 B.n410 585
R834 B.n412 B.n107 585
R835 B.n414 B.n413 585
R836 B.n415 B.n106 585
R837 B.n417 B.n416 585
R838 B.n418 B.n105 585
R839 B.n420 B.n419 585
R840 B.n421 B.n104 585
R841 B.n423 B.n422 585
R842 B.n424 B.n103 585
R843 B.n426 B.n425 585
R844 B.n427 B.n102 585
R845 B.n429 B.n428 585
R846 B.n430 B.n101 585
R847 B.n432 B.n431 585
R848 B.n433 B.n100 585
R849 B.n435 B.n434 585
R850 B.n436 B.n99 585
R851 B.n438 B.n437 585
R852 B.n439 B.n98 585
R853 B.n441 B.n440 585
R854 B.n442 B.n97 585
R855 B.n444 B.n443 585
R856 B.n445 B.n96 585
R857 B.n447 B.n446 585
R858 B.n448 B.n95 585
R859 B.n450 B.n449 585
R860 B.n451 B.n94 585
R861 B.n453 B.n452 585
R862 B.n454 B.n93 585
R863 B.n456 B.n455 585
R864 B.n457 B.n92 585
R865 B.n459 B.n458 585
R866 B.n460 B.n91 585
R867 B.n462 B.n461 585
R868 B.n463 B.n90 585
R869 B.n465 B.n464 585
R870 B.n466 B.n89 585
R871 B.n468 B.n467 585
R872 B.n469 B.n88 585
R873 B.n471 B.n470 585
R874 B.n472 B.n87 585
R875 B.n474 B.n473 585
R876 B.n475 B.n86 585
R877 B.n477 B.n476 585
R878 B.n478 B.n85 585
R879 B.n480 B.n479 585
R880 B.n481 B.n84 585
R881 B.n483 B.n482 585
R882 B.n484 B.n83 585
R883 B.n486 B.n485 585
R884 B.n487 B.n82 585
R885 B.n489 B.n488 585
R886 B.n490 B.n81 585
R887 B.n492 B.n491 585
R888 B.n493 B.n80 585
R889 B.n495 B.n494 585
R890 B.n496 B.n79 585
R891 B.n498 B.n497 585
R892 B.n499 B.n78 585
R893 B.n501 B.n500 585
R894 B.n502 B.n77 585
R895 B.n504 B.n503 585
R896 B.n505 B.n76 585
R897 B.n507 B.n506 585
R898 B.n508 B.n75 585
R899 B.n510 B.n509 585
R900 B.n657 B.n656 585
R901 B.n655 B.n22 585
R902 B.n654 B.n653 585
R903 B.n652 B.n23 585
R904 B.n651 B.n650 585
R905 B.n649 B.n24 585
R906 B.n648 B.n647 585
R907 B.n646 B.n25 585
R908 B.n645 B.n644 585
R909 B.n643 B.n26 585
R910 B.n642 B.n641 585
R911 B.n640 B.n27 585
R912 B.n639 B.n638 585
R913 B.n637 B.n28 585
R914 B.n636 B.n635 585
R915 B.n634 B.n29 585
R916 B.n633 B.n632 585
R917 B.n631 B.n30 585
R918 B.n630 B.n629 585
R919 B.n628 B.n31 585
R920 B.n627 B.n626 585
R921 B.n625 B.n32 585
R922 B.n624 B.n623 585
R923 B.n622 B.n33 585
R924 B.n621 B.n620 585
R925 B.n619 B.n34 585
R926 B.n618 B.n617 585
R927 B.n616 B.n35 585
R928 B.n615 B.n614 585
R929 B.n613 B.n36 585
R930 B.n612 B.n611 585
R931 B.n610 B.n37 585
R932 B.n609 B.n608 585
R933 B.n607 B.n38 585
R934 B.n606 B.n605 585
R935 B.n604 B.n39 585
R936 B.n603 B.n602 585
R937 B.n601 B.n40 585
R938 B.n600 B.n599 585
R939 B.n598 B.n41 585
R940 B.n597 B.n596 585
R941 B.n595 B.n42 585
R942 B.n594 B.n593 585
R943 B.n592 B.n43 585
R944 B.n590 B.n589 585
R945 B.n588 B.n46 585
R946 B.n587 B.n586 585
R947 B.n585 B.n47 585
R948 B.n584 B.n583 585
R949 B.n582 B.n48 585
R950 B.n581 B.n580 585
R951 B.n579 B.n49 585
R952 B.n578 B.n577 585
R953 B.n576 B.n575 585
R954 B.n574 B.n53 585
R955 B.n573 B.n572 585
R956 B.n571 B.n54 585
R957 B.n570 B.n569 585
R958 B.n568 B.n55 585
R959 B.n567 B.n566 585
R960 B.n565 B.n56 585
R961 B.n564 B.n563 585
R962 B.n562 B.n57 585
R963 B.n561 B.n560 585
R964 B.n559 B.n58 585
R965 B.n558 B.n557 585
R966 B.n556 B.n59 585
R967 B.n555 B.n554 585
R968 B.n553 B.n60 585
R969 B.n552 B.n551 585
R970 B.n550 B.n61 585
R971 B.n549 B.n548 585
R972 B.n547 B.n62 585
R973 B.n546 B.n545 585
R974 B.n544 B.n63 585
R975 B.n543 B.n542 585
R976 B.n541 B.n64 585
R977 B.n540 B.n539 585
R978 B.n538 B.n65 585
R979 B.n537 B.n536 585
R980 B.n535 B.n66 585
R981 B.n534 B.n533 585
R982 B.n532 B.n67 585
R983 B.n531 B.n530 585
R984 B.n529 B.n68 585
R985 B.n528 B.n527 585
R986 B.n526 B.n69 585
R987 B.n525 B.n524 585
R988 B.n523 B.n70 585
R989 B.n522 B.n521 585
R990 B.n520 B.n71 585
R991 B.n519 B.n518 585
R992 B.n517 B.n72 585
R993 B.n516 B.n515 585
R994 B.n514 B.n73 585
R995 B.n513 B.n512 585
R996 B.n511 B.n74 585
R997 B.n658 B.n21 585
R998 B.n660 B.n659 585
R999 B.n661 B.n20 585
R1000 B.n663 B.n662 585
R1001 B.n664 B.n19 585
R1002 B.n666 B.n665 585
R1003 B.n667 B.n18 585
R1004 B.n669 B.n668 585
R1005 B.n670 B.n17 585
R1006 B.n672 B.n671 585
R1007 B.n673 B.n16 585
R1008 B.n675 B.n674 585
R1009 B.n676 B.n15 585
R1010 B.n678 B.n677 585
R1011 B.n679 B.n14 585
R1012 B.n681 B.n680 585
R1013 B.n682 B.n13 585
R1014 B.n684 B.n683 585
R1015 B.n685 B.n12 585
R1016 B.n687 B.n686 585
R1017 B.n688 B.n11 585
R1018 B.n690 B.n689 585
R1019 B.n691 B.n10 585
R1020 B.n693 B.n692 585
R1021 B.n694 B.n9 585
R1022 B.n696 B.n695 585
R1023 B.n697 B.n8 585
R1024 B.n699 B.n698 585
R1025 B.n700 B.n7 585
R1026 B.n702 B.n701 585
R1027 B.n703 B.n6 585
R1028 B.n705 B.n704 585
R1029 B.n706 B.n5 585
R1030 B.n708 B.n707 585
R1031 B.n709 B.n4 585
R1032 B.n711 B.n710 585
R1033 B.n712 B.n3 585
R1034 B.n714 B.n713 585
R1035 B.n715 B.n0 585
R1036 B.n2 B.n1 585
R1037 B.n185 B.n184 585
R1038 B.n186 B.n183 585
R1039 B.n188 B.n187 585
R1040 B.n189 B.n182 585
R1041 B.n191 B.n190 585
R1042 B.n192 B.n181 585
R1043 B.n194 B.n193 585
R1044 B.n195 B.n180 585
R1045 B.n197 B.n196 585
R1046 B.n198 B.n179 585
R1047 B.n200 B.n199 585
R1048 B.n201 B.n178 585
R1049 B.n203 B.n202 585
R1050 B.n204 B.n177 585
R1051 B.n206 B.n205 585
R1052 B.n207 B.n176 585
R1053 B.n209 B.n208 585
R1054 B.n210 B.n175 585
R1055 B.n212 B.n211 585
R1056 B.n213 B.n174 585
R1057 B.n215 B.n214 585
R1058 B.n216 B.n173 585
R1059 B.n218 B.n217 585
R1060 B.n219 B.n172 585
R1061 B.n221 B.n220 585
R1062 B.n222 B.n171 585
R1063 B.n224 B.n223 585
R1064 B.n225 B.n170 585
R1065 B.n227 B.n226 585
R1066 B.n228 B.n169 585
R1067 B.n230 B.n229 585
R1068 B.n231 B.n168 585
R1069 B.n233 B.n232 585
R1070 B.n234 B.n167 585
R1071 B.n236 B.n235 585
R1072 B.n237 B.n166 585
R1073 B.n239 B.n238 585
R1074 B.n240 B.n165 585
R1075 B.n242 B.n165 550.159
R1076 B.n391 B.n390 550.159
R1077 B.n511 B.n510 550.159
R1078 B.n656 B.n21 550.159
R1079 B.n320 B.t1 441.498
R1080 B.n50 B.t11 441.498
R1081 B.n142 B.t7 441.498
R1082 B.n44 B.t5 441.498
R1083 B.n321 B.t2 389.522
R1084 B.n51 B.t10 389.522
R1085 B.n143 B.t8 389.522
R1086 B.n45 B.t4 389.522
R1087 B.n142 B.t6 338.596
R1088 B.n320 B.t0 338.596
R1089 B.n50 B.t9 338.596
R1090 B.n44 B.t3 338.596
R1091 B.n717 B.n716 256.663
R1092 B.n716 B.n715 235.042
R1093 B.n716 B.n2 235.042
R1094 B.n243 B.n242 163.367
R1095 B.n244 B.n243 163.367
R1096 B.n244 B.n163 163.367
R1097 B.n248 B.n163 163.367
R1098 B.n249 B.n248 163.367
R1099 B.n250 B.n249 163.367
R1100 B.n250 B.n161 163.367
R1101 B.n254 B.n161 163.367
R1102 B.n255 B.n254 163.367
R1103 B.n256 B.n255 163.367
R1104 B.n256 B.n159 163.367
R1105 B.n260 B.n159 163.367
R1106 B.n261 B.n260 163.367
R1107 B.n262 B.n261 163.367
R1108 B.n262 B.n157 163.367
R1109 B.n266 B.n157 163.367
R1110 B.n267 B.n266 163.367
R1111 B.n268 B.n267 163.367
R1112 B.n268 B.n155 163.367
R1113 B.n272 B.n155 163.367
R1114 B.n273 B.n272 163.367
R1115 B.n274 B.n273 163.367
R1116 B.n274 B.n153 163.367
R1117 B.n278 B.n153 163.367
R1118 B.n279 B.n278 163.367
R1119 B.n280 B.n279 163.367
R1120 B.n280 B.n151 163.367
R1121 B.n284 B.n151 163.367
R1122 B.n285 B.n284 163.367
R1123 B.n286 B.n285 163.367
R1124 B.n286 B.n149 163.367
R1125 B.n290 B.n149 163.367
R1126 B.n291 B.n290 163.367
R1127 B.n292 B.n291 163.367
R1128 B.n292 B.n147 163.367
R1129 B.n296 B.n147 163.367
R1130 B.n297 B.n296 163.367
R1131 B.n298 B.n297 163.367
R1132 B.n298 B.n145 163.367
R1133 B.n302 B.n145 163.367
R1134 B.n303 B.n302 163.367
R1135 B.n304 B.n303 163.367
R1136 B.n304 B.n141 163.367
R1137 B.n309 B.n141 163.367
R1138 B.n310 B.n309 163.367
R1139 B.n311 B.n310 163.367
R1140 B.n311 B.n139 163.367
R1141 B.n315 B.n139 163.367
R1142 B.n316 B.n315 163.367
R1143 B.n317 B.n316 163.367
R1144 B.n317 B.n137 163.367
R1145 B.n324 B.n137 163.367
R1146 B.n325 B.n324 163.367
R1147 B.n326 B.n325 163.367
R1148 B.n326 B.n135 163.367
R1149 B.n330 B.n135 163.367
R1150 B.n331 B.n330 163.367
R1151 B.n332 B.n331 163.367
R1152 B.n332 B.n133 163.367
R1153 B.n336 B.n133 163.367
R1154 B.n337 B.n336 163.367
R1155 B.n338 B.n337 163.367
R1156 B.n338 B.n131 163.367
R1157 B.n342 B.n131 163.367
R1158 B.n343 B.n342 163.367
R1159 B.n344 B.n343 163.367
R1160 B.n344 B.n129 163.367
R1161 B.n348 B.n129 163.367
R1162 B.n349 B.n348 163.367
R1163 B.n350 B.n349 163.367
R1164 B.n350 B.n127 163.367
R1165 B.n354 B.n127 163.367
R1166 B.n355 B.n354 163.367
R1167 B.n356 B.n355 163.367
R1168 B.n356 B.n125 163.367
R1169 B.n360 B.n125 163.367
R1170 B.n361 B.n360 163.367
R1171 B.n362 B.n361 163.367
R1172 B.n362 B.n123 163.367
R1173 B.n366 B.n123 163.367
R1174 B.n367 B.n366 163.367
R1175 B.n368 B.n367 163.367
R1176 B.n368 B.n121 163.367
R1177 B.n372 B.n121 163.367
R1178 B.n373 B.n372 163.367
R1179 B.n374 B.n373 163.367
R1180 B.n374 B.n119 163.367
R1181 B.n378 B.n119 163.367
R1182 B.n379 B.n378 163.367
R1183 B.n380 B.n379 163.367
R1184 B.n380 B.n117 163.367
R1185 B.n384 B.n117 163.367
R1186 B.n385 B.n384 163.367
R1187 B.n386 B.n385 163.367
R1188 B.n386 B.n115 163.367
R1189 B.n390 B.n115 163.367
R1190 B.n510 B.n75 163.367
R1191 B.n506 B.n75 163.367
R1192 B.n506 B.n505 163.367
R1193 B.n505 B.n504 163.367
R1194 B.n504 B.n77 163.367
R1195 B.n500 B.n77 163.367
R1196 B.n500 B.n499 163.367
R1197 B.n499 B.n498 163.367
R1198 B.n498 B.n79 163.367
R1199 B.n494 B.n79 163.367
R1200 B.n494 B.n493 163.367
R1201 B.n493 B.n492 163.367
R1202 B.n492 B.n81 163.367
R1203 B.n488 B.n81 163.367
R1204 B.n488 B.n487 163.367
R1205 B.n487 B.n486 163.367
R1206 B.n486 B.n83 163.367
R1207 B.n482 B.n83 163.367
R1208 B.n482 B.n481 163.367
R1209 B.n481 B.n480 163.367
R1210 B.n480 B.n85 163.367
R1211 B.n476 B.n85 163.367
R1212 B.n476 B.n475 163.367
R1213 B.n475 B.n474 163.367
R1214 B.n474 B.n87 163.367
R1215 B.n470 B.n87 163.367
R1216 B.n470 B.n469 163.367
R1217 B.n469 B.n468 163.367
R1218 B.n468 B.n89 163.367
R1219 B.n464 B.n89 163.367
R1220 B.n464 B.n463 163.367
R1221 B.n463 B.n462 163.367
R1222 B.n462 B.n91 163.367
R1223 B.n458 B.n91 163.367
R1224 B.n458 B.n457 163.367
R1225 B.n457 B.n456 163.367
R1226 B.n456 B.n93 163.367
R1227 B.n452 B.n93 163.367
R1228 B.n452 B.n451 163.367
R1229 B.n451 B.n450 163.367
R1230 B.n450 B.n95 163.367
R1231 B.n446 B.n95 163.367
R1232 B.n446 B.n445 163.367
R1233 B.n445 B.n444 163.367
R1234 B.n444 B.n97 163.367
R1235 B.n440 B.n97 163.367
R1236 B.n440 B.n439 163.367
R1237 B.n439 B.n438 163.367
R1238 B.n438 B.n99 163.367
R1239 B.n434 B.n99 163.367
R1240 B.n434 B.n433 163.367
R1241 B.n433 B.n432 163.367
R1242 B.n432 B.n101 163.367
R1243 B.n428 B.n101 163.367
R1244 B.n428 B.n427 163.367
R1245 B.n427 B.n426 163.367
R1246 B.n426 B.n103 163.367
R1247 B.n422 B.n103 163.367
R1248 B.n422 B.n421 163.367
R1249 B.n421 B.n420 163.367
R1250 B.n420 B.n105 163.367
R1251 B.n416 B.n105 163.367
R1252 B.n416 B.n415 163.367
R1253 B.n415 B.n414 163.367
R1254 B.n414 B.n107 163.367
R1255 B.n410 B.n107 163.367
R1256 B.n410 B.n409 163.367
R1257 B.n409 B.n408 163.367
R1258 B.n408 B.n109 163.367
R1259 B.n404 B.n109 163.367
R1260 B.n404 B.n403 163.367
R1261 B.n403 B.n402 163.367
R1262 B.n402 B.n111 163.367
R1263 B.n398 B.n111 163.367
R1264 B.n398 B.n397 163.367
R1265 B.n397 B.n396 163.367
R1266 B.n396 B.n113 163.367
R1267 B.n392 B.n113 163.367
R1268 B.n392 B.n391 163.367
R1269 B.n656 B.n655 163.367
R1270 B.n655 B.n654 163.367
R1271 B.n654 B.n23 163.367
R1272 B.n650 B.n23 163.367
R1273 B.n650 B.n649 163.367
R1274 B.n649 B.n648 163.367
R1275 B.n648 B.n25 163.367
R1276 B.n644 B.n25 163.367
R1277 B.n644 B.n643 163.367
R1278 B.n643 B.n642 163.367
R1279 B.n642 B.n27 163.367
R1280 B.n638 B.n27 163.367
R1281 B.n638 B.n637 163.367
R1282 B.n637 B.n636 163.367
R1283 B.n636 B.n29 163.367
R1284 B.n632 B.n29 163.367
R1285 B.n632 B.n631 163.367
R1286 B.n631 B.n630 163.367
R1287 B.n630 B.n31 163.367
R1288 B.n626 B.n31 163.367
R1289 B.n626 B.n625 163.367
R1290 B.n625 B.n624 163.367
R1291 B.n624 B.n33 163.367
R1292 B.n620 B.n33 163.367
R1293 B.n620 B.n619 163.367
R1294 B.n619 B.n618 163.367
R1295 B.n618 B.n35 163.367
R1296 B.n614 B.n35 163.367
R1297 B.n614 B.n613 163.367
R1298 B.n613 B.n612 163.367
R1299 B.n612 B.n37 163.367
R1300 B.n608 B.n37 163.367
R1301 B.n608 B.n607 163.367
R1302 B.n607 B.n606 163.367
R1303 B.n606 B.n39 163.367
R1304 B.n602 B.n39 163.367
R1305 B.n602 B.n601 163.367
R1306 B.n601 B.n600 163.367
R1307 B.n600 B.n41 163.367
R1308 B.n596 B.n41 163.367
R1309 B.n596 B.n595 163.367
R1310 B.n595 B.n594 163.367
R1311 B.n594 B.n43 163.367
R1312 B.n589 B.n43 163.367
R1313 B.n589 B.n588 163.367
R1314 B.n588 B.n587 163.367
R1315 B.n587 B.n47 163.367
R1316 B.n583 B.n47 163.367
R1317 B.n583 B.n582 163.367
R1318 B.n582 B.n581 163.367
R1319 B.n581 B.n49 163.367
R1320 B.n577 B.n49 163.367
R1321 B.n577 B.n576 163.367
R1322 B.n576 B.n53 163.367
R1323 B.n572 B.n53 163.367
R1324 B.n572 B.n571 163.367
R1325 B.n571 B.n570 163.367
R1326 B.n570 B.n55 163.367
R1327 B.n566 B.n55 163.367
R1328 B.n566 B.n565 163.367
R1329 B.n565 B.n564 163.367
R1330 B.n564 B.n57 163.367
R1331 B.n560 B.n57 163.367
R1332 B.n560 B.n559 163.367
R1333 B.n559 B.n558 163.367
R1334 B.n558 B.n59 163.367
R1335 B.n554 B.n59 163.367
R1336 B.n554 B.n553 163.367
R1337 B.n553 B.n552 163.367
R1338 B.n552 B.n61 163.367
R1339 B.n548 B.n61 163.367
R1340 B.n548 B.n547 163.367
R1341 B.n547 B.n546 163.367
R1342 B.n546 B.n63 163.367
R1343 B.n542 B.n63 163.367
R1344 B.n542 B.n541 163.367
R1345 B.n541 B.n540 163.367
R1346 B.n540 B.n65 163.367
R1347 B.n536 B.n65 163.367
R1348 B.n536 B.n535 163.367
R1349 B.n535 B.n534 163.367
R1350 B.n534 B.n67 163.367
R1351 B.n530 B.n67 163.367
R1352 B.n530 B.n529 163.367
R1353 B.n529 B.n528 163.367
R1354 B.n528 B.n69 163.367
R1355 B.n524 B.n69 163.367
R1356 B.n524 B.n523 163.367
R1357 B.n523 B.n522 163.367
R1358 B.n522 B.n71 163.367
R1359 B.n518 B.n71 163.367
R1360 B.n518 B.n517 163.367
R1361 B.n517 B.n516 163.367
R1362 B.n516 B.n73 163.367
R1363 B.n512 B.n73 163.367
R1364 B.n512 B.n511 163.367
R1365 B.n660 B.n21 163.367
R1366 B.n661 B.n660 163.367
R1367 B.n662 B.n661 163.367
R1368 B.n662 B.n19 163.367
R1369 B.n666 B.n19 163.367
R1370 B.n667 B.n666 163.367
R1371 B.n668 B.n667 163.367
R1372 B.n668 B.n17 163.367
R1373 B.n672 B.n17 163.367
R1374 B.n673 B.n672 163.367
R1375 B.n674 B.n673 163.367
R1376 B.n674 B.n15 163.367
R1377 B.n678 B.n15 163.367
R1378 B.n679 B.n678 163.367
R1379 B.n680 B.n679 163.367
R1380 B.n680 B.n13 163.367
R1381 B.n684 B.n13 163.367
R1382 B.n685 B.n684 163.367
R1383 B.n686 B.n685 163.367
R1384 B.n686 B.n11 163.367
R1385 B.n690 B.n11 163.367
R1386 B.n691 B.n690 163.367
R1387 B.n692 B.n691 163.367
R1388 B.n692 B.n9 163.367
R1389 B.n696 B.n9 163.367
R1390 B.n697 B.n696 163.367
R1391 B.n698 B.n697 163.367
R1392 B.n698 B.n7 163.367
R1393 B.n702 B.n7 163.367
R1394 B.n703 B.n702 163.367
R1395 B.n704 B.n703 163.367
R1396 B.n704 B.n5 163.367
R1397 B.n708 B.n5 163.367
R1398 B.n709 B.n708 163.367
R1399 B.n710 B.n709 163.367
R1400 B.n710 B.n3 163.367
R1401 B.n714 B.n3 163.367
R1402 B.n715 B.n714 163.367
R1403 B.n184 B.n2 163.367
R1404 B.n184 B.n183 163.367
R1405 B.n188 B.n183 163.367
R1406 B.n189 B.n188 163.367
R1407 B.n190 B.n189 163.367
R1408 B.n190 B.n181 163.367
R1409 B.n194 B.n181 163.367
R1410 B.n195 B.n194 163.367
R1411 B.n196 B.n195 163.367
R1412 B.n196 B.n179 163.367
R1413 B.n200 B.n179 163.367
R1414 B.n201 B.n200 163.367
R1415 B.n202 B.n201 163.367
R1416 B.n202 B.n177 163.367
R1417 B.n206 B.n177 163.367
R1418 B.n207 B.n206 163.367
R1419 B.n208 B.n207 163.367
R1420 B.n208 B.n175 163.367
R1421 B.n212 B.n175 163.367
R1422 B.n213 B.n212 163.367
R1423 B.n214 B.n213 163.367
R1424 B.n214 B.n173 163.367
R1425 B.n218 B.n173 163.367
R1426 B.n219 B.n218 163.367
R1427 B.n220 B.n219 163.367
R1428 B.n220 B.n171 163.367
R1429 B.n224 B.n171 163.367
R1430 B.n225 B.n224 163.367
R1431 B.n226 B.n225 163.367
R1432 B.n226 B.n169 163.367
R1433 B.n230 B.n169 163.367
R1434 B.n231 B.n230 163.367
R1435 B.n232 B.n231 163.367
R1436 B.n232 B.n167 163.367
R1437 B.n236 B.n167 163.367
R1438 B.n237 B.n236 163.367
R1439 B.n238 B.n237 163.367
R1440 B.n238 B.n165 163.367
R1441 B.n307 B.n143 59.5399
R1442 B.n322 B.n321 59.5399
R1443 B.n52 B.n51 59.5399
R1444 B.n591 B.n45 59.5399
R1445 B.n143 B.n142 51.9763
R1446 B.n321 B.n320 51.9763
R1447 B.n51 B.n50 51.9763
R1448 B.n45 B.n44 51.9763
R1449 B.n658 B.n657 35.7468
R1450 B.n509 B.n74 35.7468
R1451 B.n241 B.n240 35.7468
R1452 B.n389 B.n114 35.7468
R1453 B B.n717 18.0485
R1454 B.n659 B.n658 10.6151
R1455 B.n659 B.n20 10.6151
R1456 B.n663 B.n20 10.6151
R1457 B.n664 B.n663 10.6151
R1458 B.n665 B.n664 10.6151
R1459 B.n665 B.n18 10.6151
R1460 B.n669 B.n18 10.6151
R1461 B.n670 B.n669 10.6151
R1462 B.n671 B.n670 10.6151
R1463 B.n671 B.n16 10.6151
R1464 B.n675 B.n16 10.6151
R1465 B.n676 B.n675 10.6151
R1466 B.n677 B.n676 10.6151
R1467 B.n677 B.n14 10.6151
R1468 B.n681 B.n14 10.6151
R1469 B.n682 B.n681 10.6151
R1470 B.n683 B.n682 10.6151
R1471 B.n683 B.n12 10.6151
R1472 B.n687 B.n12 10.6151
R1473 B.n688 B.n687 10.6151
R1474 B.n689 B.n688 10.6151
R1475 B.n689 B.n10 10.6151
R1476 B.n693 B.n10 10.6151
R1477 B.n694 B.n693 10.6151
R1478 B.n695 B.n694 10.6151
R1479 B.n695 B.n8 10.6151
R1480 B.n699 B.n8 10.6151
R1481 B.n700 B.n699 10.6151
R1482 B.n701 B.n700 10.6151
R1483 B.n701 B.n6 10.6151
R1484 B.n705 B.n6 10.6151
R1485 B.n706 B.n705 10.6151
R1486 B.n707 B.n706 10.6151
R1487 B.n707 B.n4 10.6151
R1488 B.n711 B.n4 10.6151
R1489 B.n712 B.n711 10.6151
R1490 B.n713 B.n712 10.6151
R1491 B.n713 B.n0 10.6151
R1492 B.n657 B.n22 10.6151
R1493 B.n653 B.n22 10.6151
R1494 B.n653 B.n652 10.6151
R1495 B.n652 B.n651 10.6151
R1496 B.n651 B.n24 10.6151
R1497 B.n647 B.n24 10.6151
R1498 B.n647 B.n646 10.6151
R1499 B.n646 B.n645 10.6151
R1500 B.n645 B.n26 10.6151
R1501 B.n641 B.n26 10.6151
R1502 B.n641 B.n640 10.6151
R1503 B.n640 B.n639 10.6151
R1504 B.n639 B.n28 10.6151
R1505 B.n635 B.n28 10.6151
R1506 B.n635 B.n634 10.6151
R1507 B.n634 B.n633 10.6151
R1508 B.n633 B.n30 10.6151
R1509 B.n629 B.n30 10.6151
R1510 B.n629 B.n628 10.6151
R1511 B.n628 B.n627 10.6151
R1512 B.n627 B.n32 10.6151
R1513 B.n623 B.n32 10.6151
R1514 B.n623 B.n622 10.6151
R1515 B.n622 B.n621 10.6151
R1516 B.n621 B.n34 10.6151
R1517 B.n617 B.n34 10.6151
R1518 B.n617 B.n616 10.6151
R1519 B.n616 B.n615 10.6151
R1520 B.n615 B.n36 10.6151
R1521 B.n611 B.n36 10.6151
R1522 B.n611 B.n610 10.6151
R1523 B.n610 B.n609 10.6151
R1524 B.n609 B.n38 10.6151
R1525 B.n605 B.n38 10.6151
R1526 B.n605 B.n604 10.6151
R1527 B.n604 B.n603 10.6151
R1528 B.n603 B.n40 10.6151
R1529 B.n599 B.n40 10.6151
R1530 B.n599 B.n598 10.6151
R1531 B.n598 B.n597 10.6151
R1532 B.n597 B.n42 10.6151
R1533 B.n593 B.n42 10.6151
R1534 B.n593 B.n592 10.6151
R1535 B.n590 B.n46 10.6151
R1536 B.n586 B.n46 10.6151
R1537 B.n586 B.n585 10.6151
R1538 B.n585 B.n584 10.6151
R1539 B.n584 B.n48 10.6151
R1540 B.n580 B.n48 10.6151
R1541 B.n580 B.n579 10.6151
R1542 B.n579 B.n578 10.6151
R1543 B.n575 B.n574 10.6151
R1544 B.n574 B.n573 10.6151
R1545 B.n573 B.n54 10.6151
R1546 B.n569 B.n54 10.6151
R1547 B.n569 B.n568 10.6151
R1548 B.n568 B.n567 10.6151
R1549 B.n567 B.n56 10.6151
R1550 B.n563 B.n56 10.6151
R1551 B.n563 B.n562 10.6151
R1552 B.n562 B.n561 10.6151
R1553 B.n561 B.n58 10.6151
R1554 B.n557 B.n58 10.6151
R1555 B.n557 B.n556 10.6151
R1556 B.n556 B.n555 10.6151
R1557 B.n555 B.n60 10.6151
R1558 B.n551 B.n60 10.6151
R1559 B.n551 B.n550 10.6151
R1560 B.n550 B.n549 10.6151
R1561 B.n549 B.n62 10.6151
R1562 B.n545 B.n62 10.6151
R1563 B.n545 B.n544 10.6151
R1564 B.n544 B.n543 10.6151
R1565 B.n543 B.n64 10.6151
R1566 B.n539 B.n64 10.6151
R1567 B.n539 B.n538 10.6151
R1568 B.n538 B.n537 10.6151
R1569 B.n537 B.n66 10.6151
R1570 B.n533 B.n66 10.6151
R1571 B.n533 B.n532 10.6151
R1572 B.n532 B.n531 10.6151
R1573 B.n531 B.n68 10.6151
R1574 B.n527 B.n68 10.6151
R1575 B.n527 B.n526 10.6151
R1576 B.n526 B.n525 10.6151
R1577 B.n525 B.n70 10.6151
R1578 B.n521 B.n70 10.6151
R1579 B.n521 B.n520 10.6151
R1580 B.n520 B.n519 10.6151
R1581 B.n519 B.n72 10.6151
R1582 B.n515 B.n72 10.6151
R1583 B.n515 B.n514 10.6151
R1584 B.n514 B.n513 10.6151
R1585 B.n513 B.n74 10.6151
R1586 B.n509 B.n508 10.6151
R1587 B.n508 B.n507 10.6151
R1588 B.n507 B.n76 10.6151
R1589 B.n503 B.n76 10.6151
R1590 B.n503 B.n502 10.6151
R1591 B.n502 B.n501 10.6151
R1592 B.n501 B.n78 10.6151
R1593 B.n497 B.n78 10.6151
R1594 B.n497 B.n496 10.6151
R1595 B.n496 B.n495 10.6151
R1596 B.n495 B.n80 10.6151
R1597 B.n491 B.n80 10.6151
R1598 B.n491 B.n490 10.6151
R1599 B.n490 B.n489 10.6151
R1600 B.n489 B.n82 10.6151
R1601 B.n485 B.n82 10.6151
R1602 B.n485 B.n484 10.6151
R1603 B.n484 B.n483 10.6151
R1604 B.n483 B.n84 10.6151
R1605 B.n479 B.n84 10.6151
R1606 B.n479 B.n478 10.6151
R1607 B.n478 B.n477 10.6151
R1608 B.n477 B.n86 10.6151
R1609 B.n473 B.n86 10.6151
R1610 B.n473 B.n472 10.6151
R1611 B.n472 B.n471 10.6151
R1612 B.n471 B.n88 10.6151
R1613 B.n467 B.n88 10.6151
R1614 B.n467 B.n466 10.6151
R1615 B.n466 B.n465 10.6151
R1616 B.n465 B.n90 10.6151
R1617 B.n461 B.n90 10.6151
R1618 B.n461 B.n460 10.6151
R1619 B.n460 B.n459 10.6151
R1620 B.n459 B.n92 10.6151
R1621 B.n455 B.n92 10.6151
R1622 B.n455 B.n454 10.6151
R1623 B.n454 B.n453 10.6151
R1624 B.n453 B.n94 10.6151
R1625 B.n449 B.n94 10.6151
R1626 B.n449 B.n448 10.6151
R1627 B.n448 B.n447 10.6151
R1628 B.n447 B.n96 10.6151
R1629 B.n443 B.n96 10.6151
R1630 B.n443 B.n442 10.6151
R1631 B.n442 B.n441 10.6151
R1632 B.n441 B.n98 10.6151
R1633 B.n437 B.n98 10.6151
R1634 B.n437 B.n436 10.6151
R1635 B.n436 B.n435 10.6151
R1636 B.n435 B.n100 10.6151
R1637 B.n431 B.n100 10.6151
R1638 B.n431 B.n430 10.6151
R1639 B.n430 B.n429 10.6151
R1640 B.n429 B.n102 10.6151
R1641 B.n425 B.n102 10.6151
R1642 B.n425 B.n424 10.6151
R1643 B.n424 B.n423 10.6151
R1644 B.n423 B.n104 10.6151
R1645 B.n419 B.n104 10.6151
R1646 B.n419 B.n418 10.6151
R1647 B.n418 B.n417 10.6151
R1648 B.n417 B.n106 10.6151
R1649 B.n413 B.n106 10.6151
R1650 B.n413 B.n412 10.6151
R1651 B.n412 B.n411 10.6151
R1652 B.n411 B.n108 10.6151
R1653 B.n407 B.n108 10.6151
R1654 B.n407 B.n406 10.6151
R1655 B.n406 B.n405 10.6151
R1656 B.n405 B.n110 10.6151
R1657 B.n401 B.n110 10.6151
R1658 B.n401 B.n400 10.6151
R1659 B.n400 B.n399 10.6151
R1660 B.n399 B.n112 10.6151
R1661 B.n395 B.n112 10.6151
R1662 B.n395 B.n394 10.6151
R1663 B.n394 B.n393 10.6151
R1664 B.n393 B.n114 10.6151
R1665 B.n185 B.n1 10.6151
R1666 B.n186 B.n185 10.6151
R1667 B.n187 B.n186 10.6151
R1668 B.n187 B.n182 10.6151
R1669 B.n191 B.n182 10.6151
R1670 B.n192 B.n191 10.6151
R1671 B.n193 B.n192 10.6151
R1672 B.n193 B.n180 10.6151
R1673 B.n197 B.n180 10.6151
R1674 B.n198 B.n197 10.6151
R1675 B.n199 B.n198 10.6151
R1676 B.n199 B.n178 10.6151
R1677 B.n203 B.n178 10.6151
R1678 B.n204 B.n203 10.6151
R1679 B.n205 B.n204 10.6151
R1680 B.n205 B.n176 10.6151
R1681 B.n209 B.n176 10.6151
R1682 B.n210 B.n209 10.6151
R1683 B.n211 B.n210 10.6151
R1684 B.n211 B.n174 10.6151
R1685 B.n215 B.n174 10.6151
R1686 B.n216 B.n215 10.6151
R1687 B.n217 B.n216 10.6151
R1688 B.n217 B.n172 10.6151
R1689 B.n221 B.n172 10.6151
R1690 B.n222 B.n221 10.6151
R1691 B.n223 B.n222 10.6151
R1692 B.n223 B.n170 10.6151
R1693 B.n227 B.n170 10.6151
R1694 B.n228 B.n227 10.6151
R1695 B.n229 B.n228 10.6151
R1696 B.n229 B.n168 10.6151
R1697 B.n233 B.n168 10.6151
R1698 B.n234 B.n233 10.6151
R1699 B.n235 B.n234 10.6151
R1700 B.n235 B.n166 10.6151
R1701 B.n239 B.n166 10.6151
R1702 B.n240 B.n239 10.6151
R1703 B.n241 B.n164 10.6151
R1704 B.n245 B.n164 10.6151
R1705 B.n246 B.n245 10.6151
R1706 B.n247 B.n246 10.6151
R1707 B.n247 B.n162 10.6151
R1708 B.n251 B.n162 10.6151
R1709 B.n252 B.n251 10.6151
R1710 B.n253 B.n252 10.6151
R1711 B.n253 B.n160 10.6151
R1712 B.n257 B.n160 10.6151
R1713 B.n258 B.n257 10.6151
R1714 B.n259 B.n258 10.6151
R1715 B.n259 B.n158 10.6151
R1716 B.n263 B.n158 10.6151
R1717 B.n264 B.n263 10.6151
R1718 B.n265 B.n264 10.6151
R1719 B.n265 B.n156 10.6151
R1720 B.n269 B.n156 10.6151
R1721 B.n270 B.n269 10.6151
R1722 B.n271 B.n270 10.6151
R1723 B.n271 B.n154 10.6151
R1724 B.n275 B.n154 10.6151
R1725 B.n276 B.n275 10.6151
R1726 B.n277 B.n276 10.6151
R1727 B.n277 B.n152 10.6151
R1728 B.n281 B.n152 10.6151
R1729 B.n282 B.n281 10.6151
R1730 B.n283 B.n282 10.6151
R1731 B.n283 B.n150 10.6151
R1732 B.n287 B.n150 10.6151
R1733 B.n288 B.n287 10.6151
R1734 B.n289 B.n288 10.6151
R1735 B.n289 B.n148 10.6151
R1736 B.n293 B.n148 10.6151
R1737 B.n294 B.n293 10.6151
R1738 B.n295 B.n294 10.6151
R1739 B.n295 B.n146 10.6151
R1740 B.n299 B.n146 10.6151
R1741 B.n300 B.n299 10.6151
R1742 B.n301 B.n300 10.6151
R1743 B.n301 B.n144 10.6151
R1744 B.n305 B.n144 10.6151
R1745 B.n306 B.n305 10.6151
R1746 B.n308 B.n140 10.6151
R1747 B.n312 B.n140 10.6151
R1748 B.n313 B.n312 10.6151
R1749 B.n314 B.n313 10.6151
R1750 B.n314 B.n138 10.6151
R1751 B.n318 B.n138 10.6151
R1752 B.n319 B.n318 10.6151
R1753 B.n323 B.n319 10.6151
R1754 B.n327 B.n136 10.6151
R1755 B.n328 B.n327 10.6151
R1756 B.n329 B.n328 10.6151
R1757 B.n329 B.n134 10.6151
R1758 B.n333 B.n134 10.6151
R1759 B.n334 B.n333 10.6151
R1760 B.n335 B.n334 10.6151
R1761 B.n335 B.n132 10.6151
R1762 B.n339 B.n132 10.6151
R1763 B.n340 B.n339 10.6151
R1764 B.n341 B.n340 10.6151
R1765 B.n341 B.n130 10.6151
R1766 B.n345 B.n130 10.6151
R1767 B.n346 B.n345 10.6151
R1768 B.n347 B.n346 10.6151
R1769 B.n347 B.n128 10.6151
R1770 B.n351 B.n128 10.6151
R1771 B.n352 B.n351 10.6151
R1772 B.n353 B.n352 10.6151
R1773 B.n353 B.n126 10.6151
R1774 B.n357 B.n126 10.6151
R1775 B.n358 B.n357 10.6151
R1776 B.n359 B.n358 10.6151
R1777 B.n359 B.n124 10.6151
R1778 B.n363 B.n124 10.6151
R1779 B.n364 B.n363 10.6151
R1780 B.n365 B.n364 10.6151
R1781 B.n365 B.n122 10.6151
R1782 B.n369 B.n122 10.6151
R1783 B.n370 B.n369 10.6151
R1784 B.n371 B.n370 10.6151
R1785 B.n371 B.n120 10.6151
R1786 B.n375 B.n120 10.6151
R1787 B.n376 B.n375 10.6151
R1788 B.n377 B.n376 10.6151
R1789 B.n377 B.n118 10.6151
R1790 B.n381 B.n118 10.6151
R1791 B.n382 B.n381 10.6151
R1792 B.n383 B.n382 10.6151
R1793 B.n383 B.n116 10.6151
R1794 B.n387 B.n116 10.6151
R1795 B.n388 B.n387 10.6151
R1796 B.n389 B.n388 10.6151
R1797 B.n717 B.n0 8.11757
R1798 B.n717 B.n1 8.11757
R1799 B.n591 B.n590 6.5566
R1800 B.n578 B.n52 6.5566
R1801 B.n308 B.n307 6.5566
R1802 B.n323 B.n322 6.5566
R1803 B.n592 B.n591 4.05904
R1804 B.n575 B.n52 4.05904
R1805 B.n307 B.n306 4.05904
R1806 B.n322 B.n136 4.05904
R1807 VN.n3 VN.t5 164.249
R1808 VN.n17 VN.t2 164.249
R1809 VN.n25 VN.n14 161.3
R1810 VN.n24 VN.n23 161.3
R1811 VN.n22 VN.n15 161.3
R1812 VN.n21 VN.n20 161.3
R1813 VN.n19 VN.n16 161.3
R1814 VN.n11 VN.n0 161.3
R1815 VN.n10 VN.n9 161.3
R1816 VN.n8 VN.n1 161.3
R1817 VN.n7 VN.n6 161.3
R1818 VN.n5 VN.n2 161.3
R1819 VN.n4 VN.t4 130.96
R1820 VN.n12 VN.t3 130.96
R1821 VN.n18 VN.t0 130.96
R1822 VN.n26 VN.t1 130.96
R1823 VN.n13 VN.n12 101.948
R1824 VN.n27 VN.n26 101.948
R1825 VN.n6 VN.n1 56.0336
R1826 VN.n20 VN.n15 56.0336
R1827 VN VN.n27 48.4982
R1828 VN.n4 VN.n3 47.8966
R1829 VN.n18 VN.n17 47.8966
R1830 VN.n10 VN.n1 24.9531
R1831 VN.n24 VN.n15 24.9531
R1832 VN.n5 VN.n4 24.4675
R1833 VN.n6 VN.n5 24.4675
R1834 VN.n11 VN.n10 24.4675
R1835 VN.n20 VN.n19 24.4675
R1836 VN.n19 VN.n18 24.4675
R1837 VN.n25 VN.n24 24.4675
R1838 VN.n12 VN.n11 8.80862
R1839 VN.n26 VN.n25 8.80862
R1840 VN.n17 VN.n16 6.92221
R1841 VN.n3 VN.n2 6.92221
R1842 VN.n27 VN.n14 0.278367
R1843 VN.n13 VN.n0 0.278367
R1844 VN.n23 VN.n14 0.189894
R1845 VN.n23 VN.n22 0.189894
R1846 VN.n22 VN.n21 0.189894
R1847 VN.n21 VN.n16 0.189894
R1848 VN.n7 VN.n2 0.189894
R1849 VN.n8 VN.n7 0.189894
R1850 VN.n9 VN.n8 0.189894
R1851 VN.n9 VN.n0 0.189894
R1852 VN VN.n13 0.153454
R1853 VDD2.n135 VDD2.n71 756.745
R1854 VDD2.n64 VDD2.n0 756.745
R1855 VDD2.n136 VDD2.n135 585
R1856 VDD2.n134 VDD2.n133 585
R1857 VDD2.n75 VDD2.n74 585
R1858 VDD2.n128 VDD2.n127 585
R1859 VDD2.n126 VDD2.n125 585
R1860 VDD2.n79 VDD2.n78 585
R1861 VDD2.n120 VDD2.n119 585
R1862 VDD2.n118 VDD2.n117 585
R1863 VDD2.n116 VDD2.n82 585
R1864 VDD2.n86 VDD2.n83 585
R1865 VDD2.n111 VDD2.n110 585
R1866 VDD2.n109 VDD2.n108 585
R1867 VDD2.n88 VDD2.n87 585
R1868 VDD2.n103 VDD2.n102 585
R1869 VDD2.n101 VDD2.n100 585
R1870 VDD2.n92 VDD2.n91 585
R1871 VDD2.n95 VDD2.n94 585
R1872 VDD2.n23 VDD2.n22 585
R1873 VDD2.n20 VDD2.n19 585
R1874 VDD2.n29 VDD2.n28 585
R1875 VDD2.n31 VDD2.n30 585
R1876 VDD2.n16 VDD2.n15 585
R1877 VDD2.n37 VDD2.n36 585
R1878 VDD2.n40 VDD2.n39 585
R1879 VDD2.n38 VDD2.n12 585
R1880 VDD2.n45 VDD2.n11 585
R1881 VDD2.n47 VDD2.n46 585
R1882 VDD2.n49 VDD2.n48 585
R1883 VDD2.n8 VDD2.n7 585
R1884 VDD2.n55 VDD2.n54 585
R1885 VDD2.n57 VDD2.n56 585
R1886 VDD2.n4 VDD2.n3 585
R1887 VDD2.n63 VDD2.n62 585
R1888 VDD2.n65 VDD2.n64 585
R1889 VDD2.t0 VDD2.n21 329.036
R1890 VDD2.t4 VDD2.n93 329.036
R1891 VDD2.n135 VDD2.n134 171.744
R1892 VDD2.n134 VDD2.n74 171.744
R1893 VDD2.n127 VDD2.n74 171.744
R1894 VDD2.n127 VDD2.n126 171.744
R1895 VDD2.n126 VDD2.n78 171.744
R1896 VDD2.n119 VDD2.n78 171.744
R1897 VDD2.n119 VDD2.n118 171.744
R1898 VDD2.n118 VDD2.n82 171.744
R1899 VDD2.n86 VDD2.n82 171.744
R1900 VDD2.n110 VDD2.n86 171.744
R1901 VDD2.n110 VDD2.n109 171.744
R1902 VDD2.n109 VDD2.n87 171.744
R1903 VDD2.n102 VDD2.n87 171.744
R1904 VDD2.n102 VDD2.n101 171.744
R1905 VDD2.n101 VDD2.n91 171.744
R1906 VDD2.n94 VDD2.n91 171.744
R1907 VDD2.n22 VDD2.n19 171.744
R1908 VDD2.n29 VDD2.n19 171.744
R1909 VDD2.n30 VDD2.n29 171.744
R1910 VDD2.n30 VDD2.n15 171.744
R1911 VDD2.n37 VDD2.n15 171.744
R1912 VDD2.n39 VDD2.n37 171.744
R1913 VDD2.n39 VDD2.n38 171.744
R1914 VDD2.n38 VDD2.n11 171.744
R1915 VDD2.n47 VDD2.n11 171.744
R1916 VDD2.n48 VDD2.n47 171.744
R1917 VDD2.n48 VDD2.n7 171.744
R1918 VDD2.n55 VDD2.n7 171.744
R1919 VDD2.n56 VDD2.n55 171.744
R1920 VDD2.n56 VDD2.n3 171.744
R1921 VDD2.n63 VDD2.n3 171.744
R1922 VDD2.n64 VDD2.n63 171.744
R1923 VDD2.n94 VDD2.t4 85.8723
R1924 VDD2.n22 VDD2.t0 85.8723
R1925 VDD2.n70 VDD2.n69 72.176
R1926 VDD2 VDD2.n141 72.173
R1927 VDD2.n70 VDD2.n68 49.184
R1928 VDD2.n140 VDD2.n139 47.5066
R1929 VDD2.n140 VDD2.n70 42.2325
R1930 VDD2.n117 VDD2.n116 13.1884
R1931 VDD2.n46 VDD2.n45 13.1884
R1932 VDD2.n120 VDD2.n81 12.8005
R1933 VDD2.n115 VDD2.n83 12.8005
R1934 VDD2.n44 VDD2.n12 12.8005
R1935 VDD2.n49 VDD2.n10 12.8005
R1936 VDD2.n121 VDD2.n79 12.0247
R1937 VDD2.n112 VDD2.n111 12.0247
R1938 VDD2.n41 VDD2.n40 12.0247
R1939 VDD2.n50 VDD2.n8 12.0247
R1940 VDD2.n125 VDD2.n124 11.249
R1941 VDD2.n108 VDD2.n85 11.249
R1942 VDD2.n36 VDD2.n14 11.249
R1943 VDD2.n54 VDD2.n53 11.249
R1944 VDD2.n95 VDD2.n93 10.7239
R1945 VDD2.n23 VDD2.n21 10.7239
R1946 VDD2.n128 VDD2.n77 10.4732
R1947 VDD2.n107 VDD2.n88 10.4732
R1948 VDD2.n35 VDD2.n16 10.4732
R1949 VDD2.n57 VDD2.n6 10.4732
R1950 VDD2.n129 VDD2.n75 9.69747
R1951 VDD2.n104 VDD2.n103 9.69747
R1952 VDD2.n32 VDD2.n31 9.69747
R1953 VDD2.n58 VDD2.n4 9.69747
R1954 VDD2.n139 VDD2.n138 9.45567
R1955 VDD2.n68 VDD2.n67 9.45567
R1956 VDD2.n97 VDD2.n96 9.3005
R1957 VDD2.n99 VDD2.n98 9.3005
R1958 VDD2.n90 VDD2.n89 9.3005
R1959 VDD2.n105 VDD2.n104 9.3005
R1960 VDD2.n107 VDD2.n106 9.3005
R1961 VDD2.n85 VDD2.n84 9.3005
R1962 VDD2.n113 VDD2.n112 9.3005
R1963 VDD2.n115 VDD2.n114 9.3005
R1964 VDD2.n138 VDD2.n137 9.3005
R1965 VDD2.n73 VDD2.n72 9.3005
R1966 VDD2.n132 VDD2.n131 9.3005
R1967 VDD2.n130 VDD2.n129 9.3005
R1968 VDD2.n77 VDD2.n76 9.3005
R1969 VDD2.n124 VDD2.n123 9.3005
R1970 VDD2.n122 VDD2.n121 9.3005
R1971 VDD2.n81 VDD2.n80 9.3005
R1972 VDD2.n2 VDD2.n1 9.3005
R1973 VDD2.n61 VDD2.n60 9.3005
R1974 VDD2.n59 VDD2.n58 9.3005
R1975 VDD2.n6 VDD2.n5 9.3005
R1976 VDD2.n53 VDD2.n52 9.3005
R1977 VDD2.n51 VDD2.n50 9.3005
R1978 VDD2.n10 VDD2.n9 9.3005
R1979 VDD2.n25 VDD2.n24 9.3005
R1980 VDD2.n27 VDD2.n26 9.3005
R1981 VDD2.n18 VDD2.n17 9.3005
R1982 VDD2.n33 VDD2.n32 9.3005
R1983 VDD2.n35 VDD2.n34 9.3005
R1984 VDD2.n14 VDD2.n13 9.3005
R1985 VDD2.n42 VDD2.n41 9.3005
R1986 VDD2.n44 VDD2.n43 9.3005
R1987 VDD2.n67 VDD2.n66 9.3005
R1988 VDD2.n133 VDD2.n132 8.92171
R1989 VDD2.n100 VDD2.n90 8.92171
R1990 VDD2.n28 VDD2.n18 8.92171
R1991 VDD2.n62 VDD2.n61 8.92171
R1992 VDD2.n136 VDD2.n73 8.14595
R1993 VDD2.n99 VDD2.n92 8.14595
R1994 VDD2.n27 VDD2.n20 8.14595
R1995 VDD2.n65 VDD2.n2 8.14595
R1996 VDD2.n137 VDD2.n71 7.3702
R1997 VDD2.n96 VDD2.n95 7.3702
R1998 VDD2.n24 VDD2.n23 7.3702
R1999 VDD2.n66 VDD2.n0 7.3702
R2000 VDD2.n139 VDD2.n71 6.59444
R2001 VDD2.n68 VDD2.n0 6.59444
R2002 VDD2.n137 VDD2.n136 5.81868
R2003 VDD2.n96 VDD2.n92 5.81868
R2004 VDD2.n24 VDD2.n20 5.81868
R2005 VDD2.n66 VDD2.n65 5.81868
R2006 VDD2.n133 VDD2.n73 5.04292
R2007 VDD2.n100 VDD2.n99 5.04292
R2008 VDD2.n28 VDD2.n27 5.04292
R2009 VDD2.n62 VDD2.n2 5.04292
R2010 VDD2.n132 VDD2.n75 4.26717
R2011 VDD2.n103 VDD2.n90 4.26717
R2012 VDD2.n31 VDD2.n18 4.26717
R2013 VDD2.n61 VDD2.n4 4.26717
R2014 VDD2.n129 VDD2.n128 3.49141
R2015 VDD2.n104 VDD2.n88 3.49141
R2016 VDD2.n32 VDD2.n16 3.49141
R2017 VDD2.n58 VDD2.n57 3.49141
R2018 VDD2.n125 VDD2.n77 2.71565
R2019 VDD2.n108 VDD2.n107 2.71565
R2020 VDD2.n36 VDD2.n35 2.71565
R2021 VDD2.n54 VDD2.n6 2.71565
R2022 VDD2.n141 VDD2.t5 2.54592
R2023 VDD2.n141 VDD2.t3 2.54592
R2024 VDD2.n69 VDD2.t1 2.54592
R2025 VDD2.n69 VDD2.t2 2.54592
R2026 VDD2.n97 VDD2.n93 2.41282
R2027 VDD2.n25 VDD2.n21 2.41282
R2028 VDD2.n124 VDD2.n79 1.93989
R2029 VDD2.n111 VDD2.n85 1.93989
R2030 VDD2.n40 VDD2.n14 1.93989
R2031 VDD2.n53 VDD2.n8 1.93989
R2032 VDD2 VDD2.n140 1.79145
R2033 VDD2.n121 VDD2.n120 1.16414
R2034 VDD2.n112 VDD2.n83 1.16414
R2035 VDD2.n41 VDD2.n12 1.16414
R2036 VDD2.n50 VDD2.n49 1.16414
R2037 VDD2.n117 VDD2.n81 0.388379
R2038 VDD2.n116 VDD2.n115 0.388379
R2039 VDD2.n45 VDD2.n44 0.388379
R2040 VDD2.n46 VDD2.n10 0.388379
R2041 VDD2.n138 VDD2.n72 0.155672
R2042 VDD2.n131 VDD2.n72 0.155672
R2043 VDD2.n131 VDD2.n130 0.155672
R2044 VDD2.n130 VDD2.n76 0.155672
R2045 VDD2.n123 VDD2.n76 0.155672
R2046 VDD2.n123 VDD2.n122 0.155672
R2047 VDD2.n122 VDD2.n80 0.155672
R2048 VDD2.n114 VDD2.n80 0.155672
R2049 VDD2.n114 VDD2.n113 0.155672
R2050 VDD2.n113 VDD2.n84 0.155672
R2051 VDD2.n106 VDD2.n84 0.155672
R2052 VDD2.n106 VDD2.n105 0.155672
R2053 VDD2.n105 VDD2.n89 0.155672
R2054 VDD2.n98 VDD2.n89 0.155672
R2055 VDD2.n98 VDD2.n97 0.155672
R2056 VDD2.n26 VDD2.n25 0.155672
R2057 VDD2.n26 VDD2.n17 0.155672
R2058 VDD2.n33 VDD2.n17 0.155672
R2059 VDD2.n34 VDD2.n33 0.155672
R2060 VDD2.n34 VDD2.n13 0.155672
R2061 VDD2.n42 VDD2.n13 0.155672
R2062 VDD2.n43 VDD2.n42 0.155672
R2063 VDD2.n43 VDD2.n9 0.155672
R2064 VDD2.n51 VDD2.n9 0.155672
R2065 VDD2.n52 VDD2.n51 0.155672
R2066 VDD2.n52 VDD2.n5 0.155672
R2067 VDD2.n59 VDD2.n5 0.155672
R2068 VDD2.n60 VDD2.n59 0.155672
R2069 VDD2.n60 VDD2.n1 0.155672
R2070 VDD2.n67 VDD2.n1 0.155672
C0 B VDD1 2.08803f
C1 VN VP 6.82992f
C2 VN B 1.12342f
C3 VTAIL VP 7.06598f
C4 VDD2 VDD1 1.31016f
C5 VDD1 w_n3114_n3522# 2.28579f
C6 B VTAIL 3.75898f
C7 VN VDD2 6.98647f
C8 VN w_n3114_n3522# 5.85988f
C9 B VP 1.79318f
C10 VDD2 VTAIL 8.04163f
C11 VTAIL w_n3114_n3522# 3.06659f
C12 VDD2 VP 0.437263f
C13 w_n3114_n3522# VP 6.26178f
C14 VN VDD1 0.150458f
C15 B VDD2 2.15613f
C16 B w_n3114_n3522# 9.546519f
C17 VDD1 VTAIL 7.99295f
C18 VDD2 w_n3114_n3522# 2.36291f
C19 VDD1 VP 7.26987f
C20 VN VTAIL 7.05166f
C21 VDD2 VSUBS 1.884935f
C22 VDD1 VSUBS 1.767373f
C23 VTAIL VSUBS 1.169855f
C24 VN VSUBS 5.62317f
C25 VP VSUBS 2.766792f
C26 B VSUBS 4.454177f
C27 w_n3114_n3522# VSUBS 0.134861p
C28 VDD2.n0 VSUBS 0.030183f
C29 VDD2.n1 VSUBS 0.027899f
C30 VDD2.n2 VSUBS 0.014992f
C31 VDD2.n3 VSUBS 0.035434f
C32 VDD2.n4 VSUBS 0.015873f
C33 VDD2.n5 VSUBS 0.027899f
C34 VDD2.n6 VSUBS 0.014992f
C35 VDD2.n7 VSUBS 0.035434f
C36 VDD2.n8 VSUBS 0.015873f
C37 VDD2.n9 VSUBS 0.027899f
C38 VDD2.n10 VSUBS 0.014992f
C39 VDD2.n11 VSUBS 0.035434f
C40 VDD2.n12 VSUBS 0.015873f
C41 VDD2.n13 VSUBS 0.027899f
C42 VDD2.n14 VSUBS 0.014992f
C43 VDD2.n15 VSUBS 0.035434f
C44 VDD2.n16 VSUBS 0.015873f
C45 VDD2.n17 VSUBS 0.027899f
C46 VDD2.n18 VSUBS 0.014992f
C47 VDD2.n19 VSUBS 0.035434f
C48 VDD2.n20 VSUBS 0.015873f
C49 VDD2.n21 VSUBS 0.229429f
C50 VDD2.t0 VSUBS 0.076428f
C51 VDD2.n22 VSUBS 0.026576f
C52 VDD2.n23 VSUBS 0.026656f
C53 VDD2.n24 VSUBS 0.014992f
C54 VDD2.n25 VSUBS 1.46488f
C55 VDD2.n26 VSUBS 0.027899f
C56 VDD2.n27 VSUBS 0.014992f
C57 VDD2.n28 VSUBS 0.015873f
C58 VDD2.n29 VSUBS 0.035434f
C59 VDD2.n30 VSUBS 0.035434f
C60 VDD2.n31 VSUBS 0.015873f
C61 VDD2.n32 VSUBS 0.014992f
C62 VDD2.n33 VSUBS 0.027899f
C63 VDD2.n34 VSUBS 0.027899f
C64 VDD2.n35 VSUBS 0.014992f
C65 VDD2.n36 VSUBS 0.015873f
C66 VDD2.n37 VSUBS 0.035434f
C67 VDD2.n38 VSUBS 0.035434f
C68 VDD2.n39 VSUBS 0.035434f
C69 VDD2.n40 VSUBS 0.015873f
C70 VDD2.n41 VSUBS 0.014992f
C71 VDD2.n42 VSUBS 0.027899f
C72 VDD2.n43 VSUBS 0.027899f
C73 VDD2.n44 VSUBS 0.014992f
C74 VDD2.n45 VSUBS 0.015432f
C75 VDD2.n46 VSUBS 0.015432f
C76 VDD2.n47 VSUBS 0.035434f
C77 VDD2.n48 VSUBS 0.035434f
C78 VDD2.n49 VSUBS 0.015873f
C79 VDD2.n50 VSUBS 0.014992f
C80 VDD2.n51 VSUBS 0.027899f
C81 VDD2.n52 VSUBS 0.027899f
C82 VDD2.n53 VSUBS 0.014992f
C83 VDD2.n54 VSUBS 0.015873f
C84 VDD2.n55 VSUBS 0.035434f
C85 VDD2.n56 VSUBS 0.035434f
C86 VDD2.n57 VSUBS 0.015873f
C87 VDD2.n58 VSUBS 0.014992f
C88 VDD2.n59 VSUBS 0.027899f
C89 VDD2.n60 VSUBS 0.027899f
C90 VDD2.n61 VSUBS 0.014992f
C91 VDD2.n62 VSUBS 0.015873f
C92 VDD2.n63 VSUBS 0.035434f
C93 VDD2.n64 VSUBS 0.084177f
C94 VDD2.n65 VSUBS 0.015873f
C95 VDD2.n66 VSUBS 0.014992f
C96 VDD2.n67 VSUBS 0.061818f
C97 VDD2.n68 VSUBS 0.068399f
C98 VDD2.t1 VSUBS 0.281531f
C99 VDD2.t2 VSUBS 0.281531f
C100 VDD2.n69 VSUBS 2.21908f
C101 VDD2.n70 VSUBS 3.22436f
C102 VDD2.n71 VSUBS 0.030183f
C103 VDD2.n72 VSUBS 0.027899f
C104 VDD2.n73 VSUBS 0.014992f
C105 VDD2.n74 VSUBS 0.035434f
C106 VDD2.n75 VSUBS 0.015873f
C107 VDD2.n76 VSUBS 0.027899f
C108 VDD2.n77 VSUBS 0.014992f
C109 VDD2.n78 VSUBS 0.035434f
C110 VDD2.n79 VSUBS 0.015873f
C111 VDD2.n80 VSUBS 0.027899f
C112 VDD2.n81 VSUBS 0.014992f
C113 VDD2.n82 VSUBS 0.035434f
C114 VDD2.n83 VSUBS 0.015873f
C115 VDD2.n84 VSUBS 0.027899f
C116 VDD2.n85 VSUBS 0.014992f
C117 VDD2.n86 VSUBS 0.035434f
C118 VDD2.n87 VSUBS 0.035434f
C119 VDD2.n88 VSUBS 0.015873f
C120 VDD2.n89 VSUBS 0.027899f
C121 VDD2.n90 VSUBS 0.014992f
C122 VDD2.n91 VSUBS 0.035434f
C123 VDD2.n92 VSUBS 0.015873f
C124 VDD2.n93 VSUBS 0.229429f
C125 VDD2.t4 VSUBS 0.076428f
C126 VDD2.n94 VSUBS 0.026576f
C127 VDD2.n95 VSUBS 0.026656f
C128 VDD2.n96 VSUBS 0.014992f
C129 VDD2.n97 VSUBS 1.46488f
C130 VDD2.n98 VSUBS 0.027899f
C131 VDD2.n99 VSUBS 0.014992f
C132 VDD2.n100 VSUBS 0.015873f
C133 VDD2.n101 VSUBS 0.035434f
C134 VDD2.n102 VSUBS 0.035434f
C135 VDD2.n103 VSUBS 0.015873f
C136 VDD2.n104 VSUBS 0.014992f
C137 VDD2.n105 VSUBS 0.027899f
C138 VDD2.n106 VSUBS 0.027899f
C139 VDD2.n107 VSUBS 0.014992f
C140 VDD2.n108 VSUBS 0.015873f
C141 VDD2.n109 VSUBS 0.035434f
C142 VDD2.n110 VSUBS 0.035434f
C143 VDD2.n111 VSUBS 0.015873f
C144 VDD2.n112 VSUBS 0.014992f
C145 VDD2.n113 VSUBS 0.027899f
C146 VDD2.n114 VSUBS 0.027899f
C147 VDD2.n115 VSUBS 0.014992f
C148 VDD2.n116 VSUBS 0.015432f
C149 VDD2.n117 VSUBS 0.015432f
C150 VDD2.n118 VSUBS 0.035434f
C151 VDD2.n119 VSUBS 0.035434f
C152 VDD2.n120 VSUBS 0.015873f
C153 VDD2.n121 VSUBS 0.014992f
C154 VDD2.n122 VSUBS 0.027899f
C155 VDD2.n123 VSUBS 0.027899f
C156 VDD2.n124 VSUBS 0.014992f
C157 VDD2.n125 VSUBS 0.015873f
C158 VDD2.n126 VSUBS 0.035434f
C159 VDD2.n127 VSUBS 0.035434f
C160 VDD2.n128 VSUBS 0.015873f
C161 VDD2.n129 VSUBS 0.014992f
C162 VDD2.n130 VSUBS 0.027899f
C163 VDD2.n131 VSUBS 0.027899f
C164 VDD2.n132 VSUBS 0.014992f
C165 VDD2.n133 VSUBS 0.015873f
C166 VDD2.n134 VSUBS 0.035434f
C167 VDD2.n135 VSUBS 0.084177f
C168 VDD2.n136 VSUBS 0.015873f
C169 VDD2.n137 VSUBS 0.014992f
C170 VDD2.n138 VSUBS 0.061818f
C171 VDD2.n139 VSUBS 0.061463f
C172 VDD2.n140 VSUBS 2.84707f
C173 VDD2.t5 VSUBS 0.281531f
C174 VDD2.t3 VSUBS 0.281531f
C175 VDD2.n141 VSUBS 2.21903f
C176 VN.n0 VSUBS 0.041739f
C177 VN.t3 VSUBS 2.59305f
C178 VN.n1 VSUBS 0.0378f
C179 VN.n2 VSUBS 0.297903f
C180 VN.t4 VSUBS 2.59305f
C181 VN.t5 VSUBS 2.81572f
C182 VN.n3 VSUBS 0.982359f
C183 VN.n4 VSUBS 1.01983f
C184 VN.n5 VSUBS 0.059005f
C185 VN.n6 VSUBS 0.054079f
C186 VN.n7 VSUBS 0.031659f
C187 VN.n8 VSUBS 0.031659f
C188 VN.n9 VSUBS 0.031659f
C189 VN.n10 VSUBS 0.059559f
C190 VN.n11 VSUBS 0.040361f
C191 VN.n12 VSUBS 1.01007f
C192 VN.n13 VSUBS 0.049871f
C193 VN.n14 VSUBS 0.041739f
C194 VN.t1 VSUBS 2.59305f
C195 VN.n15 VSUBS 0.0378f
C196 VN.n16 VSUBS 0.297903f
C197 VN.t0 VSUBS 2.59305f
C198 VN.t2 VSUBS 2.81572f
C199 VN.n17 VSUBS 0.982359f
C200 VN.n18 VSUBS 1.01983f
C201 VN.n19 VSUBS 0.059005f
C202 VN.n20 VSUBS 0.054079f
C203 VN.n21 VSUBS 0.031659f
C204 VN.n22 VSUBS 0.031659f
C205 VN.n23 VSUBS 0.031659f
C206 VN.n24 VSUBS 0.059559f
C207 VN.n25 VSUBS 0.040361f
C208 VN.n26 VSUBS 1.01007f
C209 VN.n27 VSUBS 1.68356f
C210 B.n0 VSUBS 0.007151f
C211 B.n1 VSUBS 0.007151f
C212 B.n2 VSUBS 0.010576f
C213 B.n3 VSUBS 0.008104f
C214 B.n4 VSUBS 0.008104f
C215 B.n5 VSUBS 0.008104f
C216 B.n6 VSUBS 0.008104f
C217 B.n7 VSUBS 0.008104f
C218 B.n8 VSUBS 0.008104f
C219 B.n9 VSUBS 0.008104f
C220 B.n10 VSUBS 0.008104f
C221 B.n11 VSUBS 0.008104f
C222 B.n12 VSUBS 0.008104f
C223 B.n13 VSUBS 0.008104f
C224 B.n14 VSUBS 0.008104f
C225 B.n15 VSUBS 0.008104f
C226 B.n16 VSUBS 0.008104f
C227 B.n17 VSUBS 0.008104f
C228 B.n18 VSUBS 0.008104f
C229 B.n19 VSUBS 0.008104f
C230 B.n20 VSUBS 0.008104f
C231 B.n21 VSUBS 0.019747f
C232 B.n22 VSUBS 0.008104f
C233 B.n23 VSUBS 0.008104f
C234 B.n24 VSUBS 0.008104f
C235 B.n25 VSUBS 0.008104f
C236 B.n26 VSUBS 0.008104f
C237 B.n27 VSUBS 0.008104f
C238 B.n28 VSUBS 0.008104f
C239 B.n29 VSUBS 0.008104f
C240 B.n30 VSUBS 0.008104f
C241 B.n31 VSUBS 0.008104f
C242 B.n32 VSUBS 0.008104f
C243 B.n33 VSUBS 0.008104f
C244 B.n34 VSUBS 0.008104f
C245 B.n35 VSUBS 0.008104f
C246 B.n36 VSUBS 0.008104f
C247 B.n37 VSUBS 0.008104f
C248 B.n38 VSUBS 0.008104f
C249 B.n39 VSUBS 0.008104f
C250 B.n40 VSUBS 0.008104f
C251 B.n41 VSUBS 0.008104f
C252 B.n42 VSUBS 0.008104f
C253 B.n43 VSUBS 0.008104f
C254 B.t4 VSUBS 0.264341f
C255 B.t5 VSUBS 0.298601f
C256 B.t3 VSUBS 1.56524f
C257 B.n44 VSUBS 0.468248f
C258 B.n45 VSUBS 0.302578f
C259 B.n46 VSUBS 0.008104f
C260 B.n47 VSUBS 0.008104f
C261 B.n48 VSUBS 0.008104f
C262 B.n49 VSUBS 0.008104f
C263 B.t10 VSUBS 0.264344f
C264 B.t11 VSUBS 0.298604f
C265 B.t9 VSUBS 1.56524f
C266 B.n50 VSUBS 0.468245f
C267 B.n51 VSUBS 0.302575f
C268 B.n52 VSUBS 0.018777f
C269 B.n53 VSUBS 0.008104f
C270 B.n54 VSUBS 0.008104f
C271 B.n55 VSUBS 0.008104f
C272 B.n56 VSUBS 0.008104f
C273 B.n57 VSUBS 0.008104f
C274 B.n58 VSUBS 0.008104f
C275 B.n59 VSUBS 0.008104f
C276 B.n60 VSUBS 0.008104f
C277 B.n61 VSUBS 0.008104f
C278 B.n62 VSUBS 0.008104f
C279 B.n63 VSUBS 0.008104f
C280 B.n64 VSUBS 0.008104f
C281 B.n65 VSUBS 0.008104f
C282 B.n66 VSUBS 0.008104f
C283 B.n67 VSUBS 0.008104f
C284 B.n68 VSUBS 0.008104f
C285 B.n69 VSUBS 0.008104f
C286 B.n70 VSUBS 0.008104f
C287 B.n71 VSUBS 0.008104f
C288 B.n72 VSUBS 0.008104f
C289 B.n73 VSUBS 0.008104f
C290 B.n74 VSUBS 0.020537f
C291 B.n75 VSUBS 0.008104f
C292 B.n76 VSUBS 0.008104f
C293 B.n77 VSUBS 0.008104f
C294 B.n78 VSUBS 0.008104f
C295 B.n79 VSUBS 0.008104f
C296 B.n80 VSUBS 0.008104f
C297 B.n81 VSUBS 0.008104f
C298 B.n82 VSUBS 0.008104f
C299 B.n83 VSUBS 0.008104f
C300 B.n84 VSUBS 0.008104f
C301 B.n85 VSUBS 0.008104f
C302 B.n86 VSUBS 0.008104f
C303 B.n87 VSUBS 0.008104f
C304 B.n88 VSUBS 0.008104f
C305 B.n89 VSUBS 0.008104f
C306 B.n90 VSUBS 0.008104f
C307 B.n91 VSUBS 0.008104f
C308 B.n92 VSUBS 0.008104f
C309 B.n93 VSUBS 0.008104f
C310 B.n94 VSUBS 0.008104f
C311 B.n95 VSUBS 0.008104f
C312 B.n96 VSUBS 0.008104f
C313 B.n97 VSUBS 0.008104f
C314 B.n98 VSUBS 0.008104f
C315 B.n99 VSUBS 0.008104f
C316 B.n100 VSUBS 0.008104f
C317 B.n101 VSUBS 0.008104f
C318 B.n102 VSUBS 0.008104f
C319 B.n103 VSUBS 0.008104f
C320 B.n104 VSUBS 0.008104f
C321 B.n105 VSUBS 0.008104f
C322 B.n106 VSUBS 0.008104f
C323 B.n107 VSUBS 0.008104f
C324 B.n108 VSUBS 0.008104f
C325 B.n109 VSUBS 0.008104f
C326 B.n110 VSUBS 0.008104f
C327 B.n111 VSUBS 0.008104f
C328 B.n112 VSUBS 0.008104f
C329 B.n113 VSUBS 0.008104f
C330 B.n114 VSUBS 0.020622f
C331 B.n115 VSUBS 0.008104f
C332 B.n116 VSUBS 0.008104f
C333 B.n117 VSUBS 0.008104f
C334 B.n118 VSUBS 0.008104f
C335 B.n119 VSUBS 0.008104f
C336 B.n120 VSUBS 0.008104f
C337 B.n121 VSUBS 0.008104f
C338 B.n122 VSUBS 0.008104f
C339 B.n123 VSUBS 0.008104f
C340 B.n124 VSUBS 0.008104f
C341 B.n125 VSUBS 0.008104f
C342 B.n126 VSUBS 0.008104f
C343 B.n127 VSUBS 0.008104f
C344 B.n128 VSUBS 0.008104f
C345 B.n129 VSUBS 0.008104f
C346 B.n130 VSUBS 0.008104f
C347 B.n131 VSUBS 0.008104f
C348 B.n132 VSUBS 0.008104f
C349 B.n133 VSUBS 0.008104f
C350 B.n134 VSUBS 0.008104f
C351 B.n135 VSUBS 0.008104f
C352 B.n136 VSUBS 0.005602f
C353 B.n137 VSUBS 0.008104f
C354 B.n138 VSUBS 0.008104f
C355 B.n139 VSUBS 0.008104f
C356 B.n140 VSUBS 0.008104f
C357 B.n141 VSUBS 0.008104f
C358 B.t8 VSUBS 0.264341f
C359 B.t7 VSUBS 0.298601f
C360 B.t6 VSUBS 1.56524f
C361 B.n142 VSUBS 0.468248f
C362 B.n143 VSUBS 0.302578f
C363 B.n144 VSUBS 0.008104f
C364 B.n145 VSUBS 0.008104f
C365 B.n146 VSUBS 0.008104f
C366 B.n147 VSUBS 0.008104f
C367 B.n148 VSUBS 0.008104f
C368 B.n149 VSUBS 0.008104f
C369 B.n150 VSUBS 0.008104f
C370 B.n151 VSUBS 0.008104f
C371 B.n152 VSUBS 0.008104f
C372 B.n153 VSUBS 0.008104f
C373 B.n154 VSUBS 0.008104f
C374 B.n155 VSUBS 0.008104f
C375 B.n156 VSUBS 0.008104f
C376 B.n157 VSUBS 0.008104f
C377 B.n158 VSUBS 0.008104f
C378 B.n159 VSUBS 0.008104f
C379 B.n160 VSUBS 0.008104f
C380 B.n161 VSUBS 0.008104f
C381 B.n162 VSUBS 0.008104f
C382 B.n163 VSUBS 0.008104f
C383 B.n164 VSUBS 0.008104f
C384 B.n165 VSUBS 0.019747f
C385 B.n166 VSUBS 0.008104f
C386 B.n167 VSUBS 0.008104f
C387 B.n168 VSUBS 0.008104f
C388 B.n169 VSUBS 0.008104f
C389 B.n170 VSUBS 0.008104f
C390 B.n171 VSUBS 0.008104f
C391 B.n172 VSUBS 0.008104f
C392 B.n173 VSUBS 0.008104f
C393 B.n174 VSUBS 0.008104f
C394 B.n175 VSUBS 0.008104f
C395 B.n176 VSUBS 0.008104f
C396 B.n177 VSUBS 0.008104f
C397 B.n178 VSUBS 0.008104f
C398 B.n179 VSUBS 0.008104f
C399 B.n180 VSUBS 0.008104f
C400 B.n181 VSUBS 0.008104f
C401 B.n182 VSUBS 0.008104f
C402 B.n183 VSUBS 0.008104f
C403 B.n184 VSUBS 0.008104f
C404 B.n185 VSUBS 0.008104f
C405 B.n186 VSUBS 0.008104f
C406 B.n187 VSUBS 0.008104f
C407 B.n188 VSUBS 0.008104f
C408 B.n189 VSUBS 0.008104f
C409 B.n190 VSUBS 0.008104f
C410 B.n191 VSUBS 0.008104f
C411 B.n192 VSUBS 0.008104f
C412 B.n193 VSUBS 0.008104f
C413 B.n194 VSUBS 0.008104f
C414 B.n195 VSUBS 0.008104f
C415 B.n196 VSUBS 0.008104f
C416 B.n197 VSUBS 0.008104f
C417 B.n198 VSUBS 0.008104f
C418 B.n199 VSUBS 0.008104f
C419 B.n200 VSUBS 0.008104f
C420 B.n201 VSUBS 0.008104f
C421 B.n202 VSUBS 0.008104f
C422 B.n203 VSUBS 0.008104f
C423 B.n204 VSUBS 0.008104f
C424 B.n205 VSUBS 0.008104f
C425 B.n206 VSUBS 0.008104f
C426 B.n207 VSUBS 0.008104f
C427 B.n208 VSUBS 0.008104f
C428 B.n209 VSUBS 0.008104f
C429 B.n210 VSUBS 0.008104f
C430 B.n211 VSUBS 0.008104f
C431 B.n212 VSUBS 0.008104f
C432 B.n213 VSUBS 0.008104f
C433 B.n214 VSUBS 0.008104f
C434 B.n215 VSUBS 0.008104f
C435 B.n216 VSUBS 0.008104f
C436 B.n217 VSUBS 0.008104f
C437 B.n218 VSUBS 0.008104f
C438 B.n219 VSUBS 0.008104f
C439 B.n220 VSUBS 0.008104f
C440 B.n221 VSUBS 0.008104f
C441 B.n222 VSUBS 0.008104f
C442 B.n223 VSUBS 0.008104f
C443 B.n224 VSUBS 0.008104f
C444 B.n225 VSUBS 0.008104f
C445 B.n226 VSUBS 0.008104f
C446 B.n227 VSUBS 0.008104f
C447 B.n228 VSUBS 0.008104f
C448 B.n229 VSUBS 0.008104f
C449 B.n230 VSUBS 0.008104f
C450 B.n231 VSUBS 0.008104f
C451 B.n232 VSUBS 0.008104f
C452 B.n233 VSUBS 0.008104f
C453 B.n234 VSUBS 0.008104f
C454 B.n235 VSUBS 0.008104f
C455 B.n236 VSUBS 0.008104f
C456 B.n237 VSUBS 0.008104f
C457 B.n238 VSUBS 0.008104f
C458 B.n239 VSUBS 0.008104f
C459 B.n240 VSUBS 0.019747f
C460 B.n241 VSUBS 0.020537f
C461 B.n242 VSUBS 0.020537f
C462 B.n243 VSUBS 0.008104f
C463 B.n244 VSUBS 0.008104f
C464 B.n245 VSUBS 0.008104f
C465 B.n246 VSUBS 0.008104f
C466 B.n247 VSUBS 0.008104f
C467 B.n248 VSUBS 0.008104f
C468 B.n249 VSUBS 0.008104f
C469 B.n250 VSUBS 0.008104f
C470 B.n251 VSUBS 0.008104f
C471 B.n252 VSUBS 0.008104f
C472 B.n253 VSUBS 0.008104f
C473 B.n254 VSUBS 0.008104f
C474 B.n255 VSUBS 0.008104f
C475 B.n256 VSUBS 0.008104f
C476 B.n257 VSUBS 0.008104f
C477 B.n258 VSUBS 0.008104f
C478 B.n259 VSUBS 0.008104f
C479 B.n260 VSUBS 0.008104f
C480 B.n261 VSUBS 0.008104f
C481 B.n262 VSUBS 0.008104f
C482 B.n263 VSUBS 0.008104f
C483 B.n264 VSUBS 0.008104f
C484 B.n265 VSUBS 0.008104f
C485 B.n266 VSUBS 0.008104f
C486 B.n267 VSUBS 0.008104f
C487 B.n268 VSUBS 0.008104f
C488 B.n269 VSUBS 0.008104f
C489 B.n270 VSUBS 0.008104f
C490 B.n271 VSUBS 0.008104f
C491 B.n272 VSUBS 0.008104f
C492 B.n273 VSUBS 0.008104f
C493 B.n274 VSUBS 0.008104f
C494 B.n275 VSUBS 0.008104f
C495 B.n276 VSUBS 0.008104f
C496 B.n277 VSUBS 0.008104f
C497 B.n278 VSUBS 0.008104f
C498 B.n279 VSUBS 0.008104f
C499 B.n280 VSUBS 0.008104f
C500 B.n281 VSUBS 0.008104f
C501 B.n282 VSUBS 0.008104f
C502 B.n283 VSUBS 0.008104f
C503 B.n284 VSUBS 0.008104f
C504 B.n285 VSUBS 0.008104f
C505 B.n286 VSUBS 0.008104f
C506 B.n287 VSUBS 0.008104f
C507 B.n288 VSUBS 0.008104f
C508 B.n289 VSUBS 0.008104f
C509 B.n290 VSUBS 0.008104f
C510 B.n291 VSUBS 0.008104f
C511 B.n292 VSUBS 0.008104f
C512 B.n293 VSUBS 0.008104f
C513 B.n294 VSUBS 0.008104f
C514 B.n295 VSUBS 0.008104f
C515 B.n296 VSUBS 0.008104f
C516 B.n297 VSUBS 0.008104f
C517 B.n298 VSUBS 0.008104f
C518 B.n299 VSUBS 0.008104f
C519 B.n300 VSUBS 0.008104f
C520 B.n301 VSUBS 0.008104f
C521 B.n302 VSUBS 0.008104f
C522 B.n303 VSUBS 0.008104f
C523 B.n304 VSUBS 0.008104f
C524 B.n305 VSUBS 0.008104f
C525 B.n306 VSUBS 0.005602f
C526 B.n307 VSUBS 0.018777f
C527 B.n308 VSUBS 0.006555f
C528 B.n309 VSUBS 0.008104f
C529 B.n310 VSUBS 0.008104f
C530 B.n311 VSUBS 0.008104f
C531 B.n312 VSUBS 0.008104f
C532 B.n313 VSUBS 0.008104f
C533 B.n314 VSUBS 0.008104f
C534 B.n315 VSUBS 0.008104f
C535 B.n316 VSUBS 0.008104f
C536 B.n317 VSUBS 0.008104f
C537 B.n318 VSUBS 0.008104f
C538 B.n319 VSUBS 0.008104f
C539 B.t2 VSUBS 0.264344f
C540 B.t1 VSUBS 0.298604f
C541 B.t0 VSUBS 1.56524f
C542 B.n320 VSUBS 0.468245f
C543 B.n321 VSUBS 0.302575f
C544 B.n322 VSUBS 0.018777f
C545 B.n323 VSUBS 0.006555f
C546 B.n324 VSUBS 0.008104f
C547 B.n325 VSUBS 0.008104f
C548 B.n326 VSUBS 0.008104f
C549 B.n327 VSUBS 0.008104f
C550 B.n328 VSUBS 0.008104f
C551 B.n329 VSUBS 0.008104f
C552 B.n330 VSUBS 0.008104f
C553 B.n331 VSUBS 0.008104f
C554 B.n332 VSUBS 0.008104f
C555 B.n333 VSUBS 0.008104f
C556 B.n334 VSUBS 0.008104f
C557 B.n335 VSUBS 0.008104f
C558 B.n336 VSUBS 0.008104f
C559 B.n337 VSUBS 0.008104f
C560 B.n338 VSUBS 0.008104f
C561 B.n339 VSUBS 0.008104f
C562 B.n340 VSUBS 0.008104f
C563 B.n341 VSUBS 0.008104f
C564 B.n342 VSUBS 0.008104f
C565 B.n343 VSUBS 0.008104f
C566 B.n344 VSUBS 0.008104f
C567 B.n345 VSUBS 0.008104f
C568 B.n346 VSUBS 0.008104f
C569 B.n347 VSUBS 0.008104f
C570 B.n348 VSUBS 0.008104f
C571 B.n349 VSUBS 0.008104f
C572 B.n350 VSUBS 0.008104f
C573 B.n351 VSUBS 0.008104f
C574 B.n352 VSUBS 0.008104f
C575 B.n353 VSUBS 0.008104f
C576 B.n354 VSUBS 0.008104f
C577 B.n355 VSUBS 0.008104f
C578 B.n356 VSUBS 0.008104f
C579 B.n357 VSUBS 0.008104f
C580 B.n358 VSUBS 0.008104f
C581 B.n359 VSUBS 0.008104f
C582 B.n360 VSUBS 0.008104f
C583 B.n361 VSUBS 0.008104f
C584 B.n362 VSUBS 0.008104f
C585 B.n363 VSUBS 0.008104f
C586 B.n364 VSUBS 0.008104f
C587 B.n365 VSUBS 0.008104f
C588 B.n366 VSUBS 0.008104f
C589 B.n367 VSUBS 0.008104f
C590 B.n368 VSUBS 0.008104f
C591 B.n369 VSUBS 0.008104f
C592 B.n370 VSUBS 0.008104f
C593 B.n371 VSUBS 0.008104f
C594 B.n372 VSUBS 0.008104f
C595 B.n373 VSUBS 0.008104f
C596 B.n374 VSUBS 0.008104f
C597 B.n375 VSUBS 0.008104f
C598 B.n376 VSUBS 0.008104f
C599 B.n377 VSUBS 0.008104f
C600 B.n378 VSUBS 0.008104f
C601 B.n379 VSUBS 0.008104f
C602 B.n380 VSUBS 0.008104f
C603 B.n381 VSUBS 0.008104f
C604 B.n382 VSUBS 0.008104f
C605 B.n383 VSUBS 0.008104f
C606 B.n384 VSUBS 0.008104f
C607 B.n385 VSUBS 0.008104f
C608 B.n386 VSUBS 0.008104f
C609 B.n387 VSUBS 0.008104f
C610 B.n388 VSUBS 0.008104f
C611 B.n389 VSUBS 0.019662f
C612 B.n390 VSUBS 0.020537f
C613 B.n391 VSUBS 0.019747f
C614 B.n392 VSUBS 0.008104f
C615 B.n393 VSUBS 0.008104f
C616 B.n394 VSUBS 0.008104f
C617 B.n395 VSUBS 0.008104f
C618 B.n396 VSUBS 0.008104f
C619 B.n397 VSUBS 0.008104f
C620 B.n398 VSUBS 0.008104f
C621 B.n399 VSUBS 0.008104f
C622 B.n400 VSUBS 0.008104f
C623 B.n401 VSUBS 0.008104f
C624 B.n402 VSUBS 0.008104f
C625 B.n403 VSUBS 0.008104f
C626 B.n404 VSUBS 0.008104f
C627 B.n405 VSUBS 0.008104f
C628 B.n406 VSUBS 0.008104f
C629 B.n407 VSUBS 0.008104f
C630 B.n408 VSUBS 0.008104f
C631 B.n409 VSUBS 0.008104f
C632 B.n410 VSUBS 0.008104f
C633 B.n411 VSUBS 0.008104f
C634 B.n412 VSUBS 0.008104f
C635 B.n413 VSUBS 0.008104f
C636 B.n414 VSUBS 0.008104f
C637 B.n415 VSUBS 0.008104f
C638 B.n416 VSUBS 0.008104f
C639 B.n417 VSUBS 0.008104f
C640 B.n418 VSUBS 0.008104f
C641 B.n419 VSUBS 0.008104f
C642 B.n420 VSUBS 0.008104f
C643 B.n421 VSUBS 0.008104f
C644 B.n422 VSUBS 0.008104f
C645 B.n423 VSUBS 0.008104f
C646 B.n424 VSUBS 0.008104f
C647 B.n425 VSUBS 0.008104f
C648 B.n426 VSUBS 0.008104f
C649 B.n427 VSUBS 0.008104f
C650 B.n428 VSUBS 0.008104f
C651 B.n429 VSUBS 0.008104f
C652 B.n430 VSUBS 0.008104f
C653 B.n431 VSUBS 0.008104f
C654 B.n432 VSUBS 0.008104f
C655 B.n433 VSUBS 0.008104f
C656 B.n434 VSUBS 0.008104f
C657 B.n435 VSUBS 0.008104f
C658 B.n436 VSUBS 0.008104f
C659 B.n437 VSUBS 0.008104f
C660 B.n438 VSUBS 0.008104f
C661 B.n439 VSUBS 0.008104f
C662 B.n440 VSUBS 0.008104f
C663 B.n441 VSUBS 0.008104f
C664 B.n442 VSUBS 0.008104f
C665 B.n443 VSUBS 0.008104f
C666 B.n444 VSUBS 0.008104f
C667 B.n445 VSUBS 0.008104f
C668 B.n446 VSUBS 0.008104f
C669 B.n447 VSUBS 0.008104f
C670 B.n448 VSUBS 0.008104f
C671 B.n449 VSUBS 0.008104f
C672 B.n450 VSUBS 0.008104f
C673 B.n451 VSUBS 0.008104f
C674 B.n452 VSUBS 0.008104f
C675 B.n453 VSUBS 0.008104f
C676 B.n454 VSUBS 0.008104f
C677 B.n455 VSUBS 0.008104f
C678 B.n456 VSUBS 0.008104f
C679 B.n457 VSUBS 0.008104f
C680 B.n458 VSUBS 0.008104f
C681 B.n459 VSUBS 0.008104f
C682 B.n460 VSUBS 0.008104f
C683 B.n461 VSUBS 0.008104f
C684 B.n462 VSUBS 0.008104f
C685 B.n463 VSUBS 0.008104f
C686 B.n464 VSUBS 0.008104f
C687 B.n465 VSUBS 0.008104f
C688 B.n466 VSUBS 0.008104f
C689 B.n467 VSUBS 0.008104f
C690 B.n468 VSUBS 0.008104f
C691 B.n469 VSUBS 0.008104f
C692 B.n470 VSUBS 0.008104f
C693 B.n471 VSUBS 0.008104f
C694 B.n472 VSUBS 0.008104f
C695 B.n473 VSUBS 0.008104f
C696 B.n474 VSUBS 0.008104f
C697 B.n475 VSUBS 0.008104f
C698 B.n476 VSUBS 0.008104f
C699 B.n477 VSUBS 0.008104f
C700 B.n478 VSUBS 0.008104f
C701 B.n479 VSUBS 0.008104f
C702 B.n480 VSUBS 0.008104f
C703 B.n481 VSUBS 0.008104f
C704 B.n482 VSUBS 0.008104f
C705 B.n483 VSUBS 0.008104f
C706 B.n484 VSUBS 0.008104f
C707 B.n485 VSUBS 0.008104f
C708 B.n486 VSUBS 0.008104f
C709 B.n487 VSUBS 0.008104f
C710 B.n488 VSUBS 0.008104f
C711 B.n489 VSUBS 0.008104f
C712 B.n490 VSUBS 0.008104f
C713 B.n491 VSUBS 0.008104f
C714 B.n492 VSUBS 0.008104f
C715 B.n493 VSUBS 0.008104f
C716 B.n494 VSUBS 0.008104f
C717 B.n495 VSUBS 0.008104f
C718 B.n496 VSUBS 0.008104f
C719 B.n497 VSUBS 0.008104f
C720 B.n498 VSUBS 0.008104f
C721 B.n499 VSUBS 0.008104f
C722 B.n500 VSUBS 0.008104f
C723 B.n501 VSUBS 0.008104f
C724 B.n502 VSUBS 0.008104f
C725 B.n503 VSUBS 0.008104f
C726 B.n504 VSUBS 0.008104f
C727 B.n505 VSUBS 0.008104f
C728 B.n506 VSUBS 0.008104f
C729 B.n507 VSUBS 0.008104f
C730 B.n508 VSUBS 0.008104f
C731 B.n509 VSUBS 0.019747f
C732 B.n510 VSUBS 0.019747f
C733 B.n511 VSUBS 0.020537f
C734 B.n512 VSUBS 0.008104f
C735 B.n513 VSUBS 0.008104f
C736 B.n514 VSUBS 0.008104f
C737 B.n515 VSUBS 0.008104f
C738 B.n516 VSUBS 0.008104f
C739 B.n517 VSUBS 0.008104f
C740 B.n518 VSUBS 0.008104f
C741 B.n519 VSUBS 0.008104f
C742 B.n520 VSUBS 0.008104f
C743 B.n521 VSUBS 0.008104f
C744 B.n522 VSUBS 0.008104f
C745 B.n523 VSUBS 0.008104f
C746 B.n524 VSUBS 0.008104f
C747 B.n525 VSUBS 0.008104f
C748 B.n526 VSUBS 0.008104f
C749 B.n527 VSUBS 0.008104f
C750 B.n528 VSUBS 0.008104f
C751 B.n529 VSUBS 0.008104f
C752 B.n530 VSUBS 0.008104f
C753 B.n531 VSUBS 0.008104f
C754 B.n532 VSUBS 0.008104f
C755 B.n533 VSUBS 0.008104f
C756 B.n534 VSUBS 0.008104f
C757 B.n535 VSUBS 0.008104f
C758 B.n536 VSUBS 0.008104f
C759 B.n537 VSUBS 0.008104f
C760 B.n538 VSUBS 0.008104f
C761 B.n539 VSUBS 0.008104f
C762 B.n540 VSUBS 0.008104f
C763 B.n541 VSUBS 0.008104f
C764 B.n542 VSUBS 0.008104f
C765 B.n543 VSUBS 0.008104f
C766 B.n544 VSUBS 0.008104f
C767 B.n545 VSUBS 0.008104f
C768 B.n546 VSUBS 0.008104f
C769 B.n547 VSUBS 0.008104f
C770 B.n548 VSUBS 0.008104f
C771 B.n549 VSUBS 0.008104f
C772 B.n550 VSUBS 0.008104f
C773 B.n551 VSUBS 0.008104f
C774 B.n552 VSUBS 0.008104f
C775 B.n553 VSUBS 0.008104f
C776 B.n554 VSUBS 0.008104f
C777 B.n555 VSUBS 0.008104f
C778 B.n556 VSUBS 0.008104f
C779 B.n557 VSUBS 0.008104f
C780 B.n558 VSUBS 0.008104f
C781 B.n559 VSUBS 0.008104f
C782 B.n560 VSUBS 0.008104f
C783 B.n561 VSUBS 0.008104f
C784 B.n562 VSUBS 0.008104f
C785 B.n563 VSUBS 0.008104f
C786 B.n564 VSUBS 0.008104f
C787 B.n565 VSUBS 0.008104f
C788 B.n566 VSUBS 0.008104f
C789 B.n567 VSUBS 0.008104f
C790 B.n568 VSUBS 0.008104f
C791 B.n569 VSUBS 0.008104f
C792 B.n570 VSUBS 0.008104f
C793 B.n571 VSUBS 0.008104f
C794 B.n572 VSUBS 0.008104f
C795 B.n573 VSUBS 0.008104f
C796 B.n574 VSUBS 0.008104f
C797 B.n575 VSUBS 0.005602f
C798 B.n576 VSUBS 0.008104f
C799 B.n577 VSUBS 0.008104f
C800 B.n578 VSUBS 0.006555f
C801 B.n579 VSUBS 0.008104f
C802 B.n580 VSUBS 0.008104f
C803 B.n581 VSUBS 0.008104f
C804 B.n582 VSUBS 0.008104f
C805 B.n583 VSUBS 0.008104f
C806 B.n584 VSUBS 0.008104f
C807 B.n585 VSUBS 0.008104f
C808 B.n586 VSUBS 0.008104f
C809 B.n587 VSUBS 0.008104f
C810 B.n588 VSUBS 0.008104f
C811 B.n589 VSUBS 0.008104f
C812 B.n590 VSUBS 0.006555f
C813 B.n591 VSUBS 0.018777f
C814 B.n592 VSUBS 0.005602f
C815 B.n593 VSUBS 0.008104f
C816 B.n594 VSUBS 0.008104f
C817 B.n595 VSUBS 0.008104f
C818 B.n596 VSUBS 0.008104f
C819 B.n597 VSUBS 0.008104f
C820 B.n598 VSUBS 0.008104f
C821 B.n599 VSUBS 0.008104f
C822 B.n600 VSUBS 0.008104f
C823 B.n601 VSUBS 0.008104f
C824 B.n602 VSUBS 0.008104f
C825 B.n603 VSUBS 0.008104f
C826 B.n604 VSUBS 0.008104f
C827 B.n605 VSUBS 0.008104f
C828 B.n606 VSUBS 0.008104f
C829 B.n607 VSUBS 0.008104f
C830 B.n608 VSUBS 0.008104f
C831 B.n609 VSUBS 0.008104f
C832 B.n610 VSUBS 0.008104f
C833 B.n611 VSUBS 0.008104f
C834 B.n612 VSUBS 0.008104f
C835 B.n613 VSUBS 0.008104f
C836 B.n614 VSUBS 0.008104f
C837 B.n615 VSUBS 0.008104f
C838 B.n616 VSUBS 0.008104f
C839 B.n617 VSUBS 0.008104f
C840 B.n618 VSUBS 0.008104f
C841 B.n619 VSUBS 0.008104f
C842 B.n620 VSUBS 0.008104f
C843 B.n621 VSUBS 0.008104f
C844 B.n622 VSUBS 0.008104f
C845 B.n623 VSUBS 0.008104f
C846 B.n624 VSUBS 0.008104f
C847 B.n625 VSUBS 0.008104f
C848 B.n626 VSUBS 0.008104f
C849 B.n627 VSUBS 0.008104f
C850 B.n628 VSUBS 0.008104f
C851 B.n629 VSUBS 0.008104f
C852 B.n630 VSUBS 0.008104f
C853 B.n631 VSUBS 0.008104f
C854 B.n632 VSUBS 0.008104f
C855 B.n633 VSUBS 0.008104f
C856 B.n634 VSUBS 0.008104f
C857 B.n635 VSUBS 0.008104f
C858 B.n636 VSUBS 0.008104f
C859 B.n637 VSUBS 0.008104f
C860 B.n638 VSUBS 0.008104f
C861 B.n639 VSUBS 0.008104f
C862 B.n640 VSUBS 0.008104f
C863 B.n641 VSUBS 0.008104f
C864 B.n642 VSUBS 0.008104f
C865 B.n643 VSUBS 0.008104f
C866 B.n644 VSUBS 0.008104f
C867 B.n645 VSUBS 0.008104f
C868 B.n646 VSUBS 0.008104f
C869 B.n647 VSUBS 0.008104f
C870 B.n648 VSUBS 0.008104f
C871 B.n649 VSUBS 0.008104f
C872 B.n650 VSUBS 0.008104f
C873 B.n651 VSUBS 0.008104f
C874 B.n652 VSUBS 0.008104f
C875 B.n653 VSUBS 0.008104f
C876 B.n654 VSUBS 0.008104f
C877 B.n655 VSUBS 0.008104f
C878 B.n656 VSUBS 0.020537f
C879 B.n657 VSUBS 0.020537f
C880 B.n658 VSUBS 0.019747f
C881 B.n659 VSUBS 0.008104f
C882 B.n660 VSUBS 0.008104f
C883 B.n661 VSUBS 0.008104f
C884 B.n662 VSUBS 0.008104f
C885 B.n663 VSUBS 0.008104f
C886 B.n664 VSUBS 0.008104f
C887 B.n665 VSUBS 0.008104f
C888 B.n666 VSUBS 0.008104f
C889 B.n667 VSUBS 0.008104f
C890 B.n668 VSUBS 0.008104f
C891 B.n669 VSUBS 0.008104f
C892 B.n670 VSUBS 0.008104f
C893 B.n671 VSUBS 0.008104f
C894 B.n672 VSUBS 0.008104f
C895 B.n673 VSUBS 0.008104f
C896 B.n674 VSUBS 0.008104f
C897 B.n675 VSUBS 0.008104f
C898 B.n676 VSUBS 0.008104f
C899 B.n677 VSUBS 0.008104f
C900 B.n678 VSUBS 0.008104f
C901 B.n679 VSUBS 0.008104f
C902 B.n680 VSUBS 0.008104f
C903 B.n681 VSUBS 0.008104f
C904 B.n682 VSUBS 0.008104f
C905 B.n683 VSUBS 0.008104f
C906 B.n684 VSUBS 0.008104f
C907 B.n685 VSUBS 0.008104f
C908 B.n686 VSUBS 0.008104f
C909 B.n687 VSUBS 0.008104f
C910 B.n688 VSUBS 0.008104f
C911 B.n689 VSUBS 0.008104f
C912 B.n690 VSUBS 0.008104f
C913 B.n691 VSUBS 0.008104f
C914 B.n692 VSUBS 0.008104f
C915 B.n693 VSUBS 0.008104f
C916 B.n694 VSUBS 0.008104f
C917 B.n695 VSUBS 0.008104f
C918 B.n696 VSUBS 0.008104f
C919 B.n697 VSUBS 0.008104f
C920 B.n698 VSUBS 0.008104f
C921 B.n699 VSUBS 0.008104f
C922 B.n700 VSUBS 0.008104f
C923 B.n701 VSUBS 0.008104f
C924 B.n702 VSUBS 0.008104f
C925 B.n703 VSUBS 0.008104f
C926 B.n704 VSUBS 0.008104f
C927 B.n705 VSUBS 0.008104f
C928 B.n706 VSUBS 0.008104f
C929 B.n707 VSUBS 0.008104f
C930 B.n708 VSUBS 0.008104f
C931 B.n709 VSUBS 0.008104f
C932 B.n710 VSUBS 0.008104f
C933 B.n711 VSUBS 0.008104f
C934 B.n712 VSUBS 0.008104f
C935 B.n713 VSUBS 0.008104f
C936 B.n714 VSUBS 0.008104f
C937 B.n715 VSUBS 0.010576f
C938 B.n716 VSUBS 0.011266f
C939 B.n717 VSUBS 0.022403f
C940 VDD1.n0 VSUBS 0.030179f
C941 VDD1.n1 VSUBS 0.027894f
C942 VDD1.n2 VSUBS 0.014989f
C943 VDD1.n3 VSUBS 0.035429f
C944 VDD1.n4 VSUBS 0.015871f
C945 VDD1.n5 VSUBS 0.027894f
C946 VDD1.n6 VSUBS 0.014989f
C947 VDD1.n7 VSUBS 0.035429f
C948 VDD1.n8 VSUBS 0.015871f
C949 VDD1.n9 VSUBS 0.027894f
C950 VDD1.n10 VSUBS 0.014989f
C951 VDD1.n11 VSUBS 0.035429f
C952 VDD1.n12 VSUBS 0.015871f
C953 VDD1.n13 VSUBS 0.027894f
C954 VDD1.n14 VSUBS 0.014989f
C955 VDD1.n15 VSUBS 0.035429f
C956 VDD1.n16 VSUBS 0.035429f
C957 VDD1.n17 VSUBS 0.015871f
C958 VDD1.n18 VSUBS 0.027894f
C959 VDD1.n19 VSUBS 0.014989f
C960 VDD1.n20 VSUBS 0.035429f
C961 VDD1.n21 VSUBS 0.015871f
C962 VDD1.n22 VSUBS 0.229394f
C963 VDD1.t0 VSUBS 0.076416f
C964 VDD1.n23 VSUBS 0.026572f
C965 VDD1.n24 VSUBS 0.026652f
C966 VDD1.n25 VSUBS 0.014989f
C967 VDD1.n26 VSUBS 1.46465f
C968 VDD1.n27 VSUBS 0.027894f
C969 VDD1.n28 VSUBS 0.014989f
C970 VDD1.n29 VSUBS 0.015871f
C971 VDD1.n30 VSUBS 0.035429f
C972 VDD1.n31 VSUBS 0.035429f
C973 VDD1.n32 VSUBS 0.015871f
C974 VDD1.n33 VSUBS 0.014989f
C975 VDD1.n34 VSUBS 0.027894f
C976 VDD1.n35 VSUBS 0.027894f
C977 VDD1.n36 VSUBS 0.014989f
C978 VDD1.n37 VSUBS 0.015871f
C979 VDD1.n38 VSUBS 0.035429f
C980 VDD1.n39 VSUBS 0.035429f
C981 VDD1.n40 VSUBS 0.015871f
C982 VDD1.n41 VSUBS 0.014989f
C983 VDD1.n42 VSUBS 0.027894f
C984 VDD1.n43 VSUBS 0.027894f
C985 VDD1.n44 VSUBS 0.014989f
C986 VDD1.n45 VSUBS 0.01543f
C987 VDD1.n46 VSUBS 0.01543f
C988 VDD1.n47 VSUBS 0.035429f
C989 VDD1.n48 VSUBS 0.035429f
C990 VDD1.n49 VSUBS 0.015871f
C991 VDD1.n50 VSUBS 0.014989f
C992 VDD1.n51 VSUBS 0.027894f
C993 VDD1.n52 VSUBS 0.027894f
C994 VDD1.n53 VSUBS 0.014989f
C995 VDD1.n54 VSUBS 0.015871f
C996 VDD1.n55 VSUBS 0.035429f
C997 VDD1.n56 VSUBS 0.035429f
C998 VDD1.n57 VSUBS 0.015871f
C999 VDD1.n58 VSUBS 0.014989f
C1000 VDD1.n59 VSUBS 0.027894f
C1001 VDD1.n60 VSUBS 0.027894f
C1002 VDD1.n61 VSUBS 0.014989f
C1003 VDD1.n62 VSUBS 0.015871f
C1004 VDD1.n63 VSUBS 0.035429f
C1005 VDD1.n64 VSUBS 0.084164f
C1006 VDD1.n65 VSUBS 0.015871f
C1007 VDD1.n66 VSUBS 0.014989f
C1008 VDD1.n67 VSUBS 0.061809f
C1009 VDD1.n68 VSUBS 0.069197f
C1010 VDD1.n69 VSUBS 0.030179f
C1011 VDD1.n70 VSUBS 0.027894f
C1012 VDD1.n71 VSUBS 0.014989f
C1013 VDD1.n72 VSUBS 0.035429f
C1014 VDD1.n73 VSUBS 0.015871f
C1015 VDD1.n74 VSUBS 0.027894f
C1016 VDD1.n75 VSUBS 0.014989f
C1017 VDD1.n76 VSUBS 0.035429f
C1018 VDD1.n77 VSUBS 0.015871f
C1019 VDD1.n78 VSUBS 0.027894f
C1020 VDD1.n79 VSUBS 0.014989f
C1021 VDD1.n80 VSUBS 0.035429f
C1022 VDD1.n81 VSUBS 0.015871f
C1023 VDD1.n82 VSUBS 0.027894f
C1024 VDD1.n83 VSUBS 0.014989f
C1025 VDD1.n84 VSUBS 0.035429f
C1026 VDD1.n85 VSUBS 0.015871f
C1027 VDD1.n86 VSUBS 0.027894f
C1028 VDD1.n87 VSUBS 0.014989f
C1029 VDD1.n88 VSUBS 0.035429f
C1030 VDD1.n89 VSUBS 0.015871f
C1031 VDD1.n90 VSUBS 0.229394f
C1032 VDD1.t4 VSUBS 0.076416f
C1033 VDD1.n91 VSUBS 0.026572f
C1034 VDD1.n92 VSUBS 0.026652f
C1035 VDD1.n93 VSUBS 0.014989f
C1036 VDD1.n94 VSUBS 1.46465f
C1037 VDD1.n95 VSUBS 0.027894f
C1038 VDD1.n96 VSUBS 0.014989f
C1039 VDD1.n97 VSUBS 0.015871f
C1040 VDD1.n98 VSUBS 0.035429f
C1041 VDD1.n99 VSUBS 0.035429f
C1042 VDD1.n100 VSUBS 0.015871f
C1043 VDD1.n101 VSUBS 0.014989f
C1044 VDD1.n102 VSUBS 0.027894f
C1045 VDD1.n103 VSUBS 0.027894f
C1046 VDD1.n104 VSUBS 0.014989f
C1047 VDD1.n105 VSUBS 0.015871f
C1048 VDD1.n106 VSUBS 0.035429f
C1049 VDD1.n107 VSUBS 0.035429f
C1050 VDD1.n108 VSUBS 0.035429f
C1051 VDD1.n109 VSUBS 0.015871f
C1052 VDD1.n110 VSUBS 0.014989f
C1053 VDD1.n111 VSUBS 0.027894f
C1054 VDD1.n112 VSUBS 0.027894f
C1055 VDD1.n113 VSUBS 0.014989f
C1056 VDD1.n114 VSUBS 0.01543f
C1057 VDD1.n115 VSUBS 0.01543f
C1058 VDD1.n116 VSUBS 0.035429f
C1059 VDD1.n117 VSUBS 0.035429f
C1060 VDD1.n118 VSUBS 0.015871f
C1061 VDD1.n119 VSUBS 0.014989f
C1062 VDD1.n120 VSUBS 0.027894f
C1063 VDD1.n121 VSUBS 0.027894f
C1064 VDD1.n122 VSUBS 0.014989f
C1065 VDD1.n123 VSUBS 0.015871f
C1066 VDD1.n124 VSUBS 0.035429f
C1067 VDD1.n125 VSUBS 0.035429f
C1068 VDD1.n126 VSUBS 0.015871f
C1069 VDD1.n127 VSUBS 0.014989f
C1070 VDD1.n128 VSUBS 0.027894f
C1071 VDD1.n129 VSUBS 0.027894f
C1072 VDD1.n130 VSUBS 0.014989f
C1073 VDD1.n131 VSUBS 0.015871f
C1074 VDD1.n132 VSUBS 0.035429f
C1075 VDD1.n133 VSUBS 0.084164f
C1076 VDD1.n134 VSUBS 0.015871f
C1077 VDD1.n135 VSUBS 0.014989f
C1078 VDD1.n136 VSUBS 0.061809f
C1079 VDD1.n137 VSUBS 0.068388f
C1080 VDD1.t2 VSUBS 0.281488f
C1081 VDD1.t3 VSUBS 0.281488f
C1082 VDD1.n138 VSUBS 2.21874f
C1083 VDD1.n139 VSUBS 3.35575f
C1084 VDD1.t1 VSUBS 0.281488f
C1085 VDD1.t5 VSUBS 0.281488f
C1086 VDD1.n140 VSUBS 2.21292f
C1087 VDD1.n141 VSUBS 3.40665f
C1088 VTAIL.t4 VSUBS 0.290255f
C1089 VTAIL.t0 VSUBS 0.290255f
C1090 VTAIL.n0 VSUBS 2.11568f
C1091 VTAIL.n1 VSUBS 0.889765f
C1092 VTAIL.n2 VSUBS 0.031118f
C1093 VTAIL.n3 VSUBS 0.028763f
C1094 VTAIL.n4 VSUBS 0.015456f
C1095 VTAIL.n5 VSUBS 0.036533f
C1096 VTAIL.n6 VSUBS 0.016365f
C1097 VTAIL.n7 VSUBS 0.028763f
C1098 VTAIL.n8 VSUBS 0.015456f
C1099 VTAIL.n9 VSUBS 0.036533f
C1100 VTAIL.n10 VSUBS 0.016365f
C1101 VTAIL.n11 VSUBS 0.028763f
C1102 VTAIL.n12 VSUBS 0.015456f
C1103 VTAIL.n13 VSUBS 0.036533f
C1104 VTAIL.n14 VSUBS 0.016365f
C1105 VTAIL.n15 VSUBS 0.028763f
C1106 VTAIL.n16 VSUBS 0.015456f
C1107 VTAIL.n17 VSUBS 0.036533f
C1108 VTAIL.n18 VSUBS 0.016365f
C1109 VTAIL.n19 VSUBS 0.028763f
C1110 VTAIL.n20 VSUBS 0.015456f
C1111 VTAIL.n21 VSUBS 0.036533f
C1112 VTAIL.n22 VSUBS 0.016365f
C1113 VTAIL.n23 VSUBS 0.236538f
C1114 VTAIL.t8 VSUBS 0.078796f
C1115 VTAIL.n24 VSUBS 0.027399f
C1116 VTAIL.n25 VSUBS 0.027482f
C1117 VTAIL.n26 VSUBS 0.015456f
C1118 VTAIL.n27 VSUBS 1.51027f
C1119 VTAIL.n28 VSUBS 0.028763f
C1120 VTAIL.n29 VSUBS 0.015456f
C1121 VTAIL.n30 VSUBS 0.016365f
C1122 VTAIL.n31 VSUBS 0.036533f
C1123 VTAIL.n32 VSUBS 0.036533f
C1124 VTAIL.n33 VSUBS 0.016365f
C1125 VTAIL.n34 VSUBS 0.015456f
C1126 VTAIL.n35 VSUBS 0.028763f
C1127 VTAIL.n36 VSUBS 0.028763f
C1128 VTAIL.n37 VSUBS 0.015456f
C1129 VTAIL.n38 VSUBS 0.016365f
C1130 VTAIL.n39 VSUBS 0.036533f
C1131 VTAIL.n40 VSUBS 0.036533f
C1132 VTAIL.n41 VSUBS 0.036533f
C1133 VTAIL.n42 VSUBS 0.016365f
C1134 VTAIL.n43 VSUBS 0.015456f
C1135 VTAIL.n44 VSUBS 0.028763f
C1136 VTAIL.n45 VSUBS 0.028763f
C1137 VTAIL.n46 VSUBS 0.015456f
C1138 VTAIL.n47 VSUBS 0.015911f
C1139 VTAIL.n48 VSUBS 0.015911f
C1140 VTAIL.n49 VSUBS 0.036533f
C1141 VTAIL.n50 VSUBS 0.036533f
C1142 VTAIL.n51 VSUBS 0.016365f
C1143 VTAIL.n52 VSUBS 0.015456f
C1144 VTAIL.n53 VSUBS 0.028763f
C1145 VTAIL.n54 VSUBS 0.028763f
C1146 VTAIL.n55 VSUBS 0.015456f
C1147 VTAIL.n56 VSUBS 0.016365f
C1148 VTAIL.n57 VSUBS 0.036533f
C1149 VTAIL.n58 VSUBS 0.036533f
C1150 VTAIL.n59 VSUBS 0.016365f
C1151 VTAIL.n60 VSUBS 0.015456f
C1152 VTAIL.n61 VSUBS 0.028763f
C1153 VTAIL.n62 VSUBS 0.028763f
C1154 VTAIL.n63 VSUBS 0.015456f
C1155 VTAIL.n64 VSUBS 0.016365f
C1156 VTAIL.n65 VSUBS 0.036533f
C1157 VTAIL.n66 VSUBS 0.086786f
C1158 VTAIL.n67 VSUBS 0.016365f
C1159 VTAIL.n68 VSUBS 0.015456f
C1160 VTAIL.n69 VSUBS 0.063734f
C1161 VTAIL.n70 VSUBS 0.043484f
C1162 VTAIL.n71 VSUBS 0.387747f
C1163 VTAIL.t6 VSUBS 0.290255f
C1164 VTAIL.t7 VSUBS 0.290255f
C1165 VTAIL.n72 VSUBS 2.11568f
C1166 VTAIL.n73 VSUBS 2.73361f
C1167 VTAIL.t3 VSUBS 0.290255f
C1168 VTAIL.t11 VSUBS 0.290255f
C1169 VTAIL.n74 VSUBS 2.11569f
C1170 VTAIL.n75 VSUBS 2.7336f
C1171 VTAIL.n76 VSUBS 0.031118f
C1172 VTAIL.n77 VSUBS 0.028763f
C1173 VTAIL.n78 VSUBS 0.015456f
C1174 VTAIL.n79 VSUBS 0.036533f
C1175 VTAIL.n80 VSUBS 0.016365f
C1176 VTAIL.n81 VSUBS 0.028763f
C1177 VTAIL.n82 VSUBS 0.015456f
C1178 VTAIL.n83 VSUBS 0.036533f
C1179 VTAIL.n84 VSUBS 0.016365f
C1180 VTAIL.n85 VSUBS 0.028763f
C1181 VTAIL.n86 VSUBS 0.015456f
C1182 VTAIL.n87 VSUBS 0.036533f
C1183 VTAIL.n88 VSUBS 0.016365f
C1184 VTAIL.n89 VSUBS 0.028763f
C1185 VTAIL.n90 VSUBS 0.015456f
C1186 VTAIL.n91 VSUBS 0.036533f
C1187 VTAIL.n92 VSUBS 0.036533f
C1188 VTAIL.n93 VSUBS 0.016365f
C1189 VTAIL.n94 VSUBS 0.028763f
C1190 VTAIL.n95 VSUBS 0.015456f
C1191 VTAIL.n96 VSUBS 0.036533f
C1192 VTAIL.n97 VSUBS 0.016365f
C1193 VTAIL.n98 VSUBS 0.236538f
C1194 VTAIL.t2 VSUBS 0.078796f
C1195 VTAIL.n99 VSUBS 0.027399f
C1196 VTAIL.n100 VSUBS 0.027482f
C1197 VTAIL.n101 VSUBS 0.015456f
C1198 VTAIL.n102 VSUBS 1.51027f
C1199 VTAIL.n103 VSUBS 0.028763f
C1200 VTAIL.n104 VSUBS 0.015456f
C1201 VTAIL.n105 VSUBS 0.016365f
C1202 VTAIL.n106 VSUBS 0.036533f
C1203 VTAIL.n107 VSUBS 0.036533f
C1204 VTAIL.n108 VSUBS 0.016365f
C1205 VTAIL.n109 VSUBS 0.015456f
C1206 VTAIL.n110 VSUBS 0.028763f
C1207 VTAIL.n111 VSUBS 0.028763f
C1208 VTAIL.n112 VSUBS 0.015456f
C1209 VTAIL.n113 VSUBS 0.016365f
C1210 VTAIL.n114 VSUBS 0.036533f
C1211 VTAIL.n115 VSUBS 0.036533f
C1212 VTAIL.n116 VSUBS 0.016365f
C1213 VTAIL.n117 VSUBS 0.015456f
C1214 VTAIL.n118 VSUBS 0.028763f
C1215 VTAIL.n119 VSUBS 0.028763f
C1216 VTAIL.n120 VSUBS 0.015456f
C1217 VTAIL.n121 VSUBS 0.015911f
C1218 VTAIL.n122 VSUBS 0.015911f
C1219 VTAIL.n123 VSUBS 0.036533f
C1220 VTAIL.n124 VSUBS 0.036533f
C1221 VTAIL.n125 VSUBS 0.016365f
C1222 VTAIL.n126 VSUBS 0.015456f
C1223 VTAIL.n127 VSUBS 0.028763f
C1224 VTAIL.n128 VSUBS 0.028763f
C1225 VTAIL.n129 VSUBS 0.015456f
C1226 VTAIL.n130 VSUBS 0.016365f
C1227 VTAIL.n131 VSUBS 0.036533f
C1228 VTAIL.n132 VSUBS 0.036533f
C1229 VTAIL.n133 VSUBS 0.016365f
C1230 VTAIL.n134 VSUBS 0.015456f
C1231 VTAIL.n135 VSUBS 0.028763f
C1232 VTAIL.n136 VSUBS 0.028763f
C1233 VTAIL.n137 VSUBS 0.015456f
C1234 VTAIL.n138 VSUBS 0.016365f
C1235 VTAIL.n139 VSUBS 0.036533f
C1236 VTAIL.n140 VSUBS 0.086786f
C1237 VTAIL.n141 VSUBS 0.016365f
C1238 VTAIL.n142 VSUBS 0.015456f
C1239 VTAIL.n143 VSUBS 0.063734f
C1240 VTAIL.n144 VSUBS 0.043484f
C1241 VTAIL.n145 VSUBS 0.387747f
C1242 VTAIL.t9 VSUBS 0.290255f
C1243 VTAIL.t10 VSUBS 0.290255f
C1244 VTAIL.n146 VSUBS 2.11569f
C1245 VTAIL.n147 VSUBS 1.04496f
C1246 VTAIL.n148 VSUBS 0.031118f
C1247 VTAIL.n149 VSUBS 0.028763f
C1248 VTAIL.n150 VSUBS 0.015456f
C1249 VTAIL.n151 VSUBS 0.036533f
C1250 VTAIL.n152 VSUBS 0.016365f
C1251 VTAIL.n153 VSUBS 0.028763f
C1252 VTAIL.n154 VSUBS 0.015456f
C1253 VTAIL.n155 VSUBS 0.036533f
C1254 VTAIL.n156 VSUBS 0.016365f
C1255 VTAIL.n157 VSUBS 0.028763f
C1256 VTAIL.n158 VSUBS 0.015456f
C1257 VTAIL.n159 VSUBS 0.036533f
C1258 VTAIL.n160 VSUBS 0.016365f
C1259 VTAIL.n161 VSUBS 0.028763f
C1260 VTAIL.n162 VSUBS 0.015456f
C1261 VTAIL.n163 VSUBS 0.036533f
C1262 VTAIL.n164 VSUBS 0.036533f
C1263 VTAIL.n165 VSUBS 0.016365f
C1264 VTAIL.n166 VSUBS 0.028763f
C1265 VTAIL.n167 VSUBS 0.015456f
C1266 VTAIL.n168 VSUBS 0.036533f
C1267 VTAIL.n169 VSUBS 0.016365f
C1268 VTAIL.n170 VSUBS 0.236538f
C1269 VTAIL.t5 VSUBS 0.078796f
C1270 VTAIL.n171 VSUBS 0.027399f
C1271 VTAIL.n172 VSUBS 0.027482f
C1272 VTAIL.n173 VSUBS 0.015456f
C1273 VTAIL.n174 VSUBS 1.51027f
C1274 VTAIL.n175 VSUBS 0.028763f
C1275 VTAIL.n176 VSUBS 0.015456f
C1276 VTAIL.n177 VSUBS 0.016365f
C1277 VTAIL.n178 VSUBS 0.036533f
C1278 VTAIL.n179 VSUBS 0.036533f
C1279 VTAIL.n180 VSUBS 0.016365f
C1280 VTAIL.n181 VSUBS 0.015456f
C1281 VTAIL.n182 VSUBS 0.028763f
C1282 VTAIL.n183 VSUBS 0.028763f
C1283 VTAIL.n184 VSUBS 0.015456f
C1284 VTAIL.n185 VSUBS 0.016365f
C1285 VTAIL.n186 VSUBS 0.036533f
C1286 VTAIL.n187 VSUBS 0.036533f
C1287 VTAIL.n188 VSUBS 0.016365f
C1288 VTAIL.n189 VSUBS 0.015456f
C1289 VTAIL.n190 VSUBS 0.028763f
C1290 VTAIL.n191 VSUBS 0.028763f
C1291 VTAIL.n192 VSUBS 0.015456f
C1292 VTAIL.n193 VSUBS 0.015911f
C1293 VTAIL.n194 VSUBS 0.015911f
C1294 VTAIL.n195 VSUBS 0.036533f
C1295 VTAIL.n196 VSUBS 0.036533f
C1296 VTAIL.n197 VSUBS 0.016365f
C1297 VTAIL.n198 VSUBS 0.015456f
C1298 VTAIL.n199 VSUBS 0.028763f
C1299 VTAIL.n200 VSUBS 0.028763f
C1300 VTAIL.n201 VSUBS 0.015456f
C1301 VTAIL.n202 VSUBS 0.016365f
C1302 VTAIL.n203 VSUBS 0.036533f
C1303 VTAIL.n204 VSUBS 0.036533f
C1304 VTAIL.n205 VSUBS 0.016365f
C1305 VTAIL.n206 VSUBS 0.015456f
C1306 VTAIL.n207 VSUBS 0.028763f
C1307 VTAIL.n208 VSUBS 0.028763f
C1308 VTAIL.n209 VSUBS 0.015456f
C1309 VTAIL.n210 VSUBS 0.016365f
C1310 VTAIL.n211 VSUBS 0.036533f
C1311 VTAIL.n212 VSUBS 0.086786f
C1312 VTAIL.n213 VSUBS 0.016365f
C1313 VTAIL.n214 VSUBS 0.015456f
C1314 VTAIL.n215 VSUBS 0.063734f
C1315 VTAIL.n216 VSUBS 0.043484f
C1316 VTAIL.n217 VSUBS 1.86227f
C1317 VTAIL.n218 VSUBS 0.031118f
C1318 VTAIL.n219 VSUBS 0.028763f
C1319 VTAIL.n220 VSUBS 0.015456f
C1320 VTAIL.n221 VSUBS 0.036533f
C1321 VTAIL.n222 VSUBS 0.016365f
C1322 VTAIL.n223 VSUBS 0.028763f
C1323 VTAIL.n224 VSUBS 0.015456f
C1324 VTAIL.n225 VSUBS 0.036533f
C1325 VTAIL.n226 VSUBS 0.016365f
C1326 VTAIL.n227 VSUBS 0.028763f
C1327 VTAIL.n228 VSUBS 0.015456f
C1328 VTAIL.n229 VSUBS 0.036533f
C1329 VTAIL.n230 VSUBS 0.016365f
C1330 VTAIL.n231 VSUBS 0.028763f
C1331 VTAIL.n232 VSUBS 0.015456f
C1332 VTAIL.n233 VSUBS 0.036533f
C1333 VTAIL.n234 VSUBS 0.016365f
C1334 VTAIL.n235 VSUBS 0.028763f
C1335 VTAIL.n236 VSUBS 0.015456f
C1336 VTAIL.n237 VSUBS 0.036533f
C1337 VTAIL.n238 VSUBS 0.016365f
C1338 VTAIL.n239 VSUBS 0.236538f
C1339 VTAIL.t1 VSUBS 0.078796f
C1340 VTAIL.n240 VSUBS 0.027399f
C1341 VTAIL.n241 VSUBS 0.027482f
C1342 VTAIL.n242 VSUBS 0.015456f
C1343 VTAIL.n243 VSUBS 1.51027f
C1344 VTAIL.n244 VSUBS 0.028763f
C1345 VTAIL.n245 VSUBS 0.015456f
C1346 VTAIL.n246 VSUBS 0.016365f
C1347 VTAIL.n247 VSUBS 0.036533f
C1348 VTAIL.n248 VSUBS 0.036533f
C1349 VTAIL.n249 VSUBS 0.016365f
C1350 VTAIL.n250 VSUBS 0.015456f
C1351 VTAIL.n251 VSUBS 0.028763f
C1352 VTAIL.n252 VSUBS 0.028763f
C1353 VTAIL.n253 VSUBS 0.015456f
C1354 VTAIL.n254 VSUBS 0.016365f
C1355 VTAIL.n255 VSUBS 0.036533f
C1356 VTAIL.n256 VSUBS 0.036533f
C1357 VTAIL.n257 VSUBS 0.036533f
C1358 VTAIL.n258 VSUBS 0.016365f
C1359 VTAIL.n259 VSUBS 0.015456f
C1360 VTAIL.n260 VSUBS 0.028763f
C1361 VTAIL.n261 VSUBS 0.028763f
C1362 VTAIL.n262 VSUBS 0.015456f
C1363 VTAIL.n263 VSUBS 0.015911f
C1364 VTAIL.n264 VSUBS 0.015911f
C1365 VTAIL.n265 VSUBS 0.036533f
C1366 VTAIL.n266 VSUBS 0.036533f
C1367 VTAIL.n267 VSUBS 0.016365f
C1368 VTAIL.n268 VSUBS 0.015456f
C1369 VTAIL.n269 VSUBS 0.028763f
C1370 VTAIL.n270 VSUBS 0.028763f
C1371 VTAIL.n271 VSUBS 0.015456f
C1372 VTAIL.n272 VSUBS 0.016365f
C1373 VTAIL.n273 VSUBS 0.036533f
C1374 VTAIL.n274 VSUBS 0.036533f
C1375 VTAIL.n275 VSUBS 0.016365f
C1376 VTAIL.n276 VSUBS 0.015456f
C1377 VTAIL.n277 VSUBS 0.028763f
C1378 VTAIL.n278 VSUBS 0.028763f
C1379 VTAIL.n279 VSUBS 0.015456f
C1380 VTAIL.n280 VSUBS 0.016365f
C1381 VTAIL.n281 VSUBS 0.036533f
C1382 VTAIL.n282 VSUBS 0.086786f
C1383 VTAIL.n283 VSUBS 0.016365f
C1384 VTAIL.n284 VSUBS 0.015456f
C1385 VTAIL.n285 VSUBS 0.063734f
C1386 VTAIL.n286 VSUBS 0.043484f
C1387 VTAIL.n287 VSUBS 1.80335f
C1388 VP.n0 VSUBS 0.042901f
C1389 VP.t2 VSUBS 2.66521f
C1390 VP.n1 VSUBS 0.038852f
C1391 VP.n2 VSUBS 0.03254f
C1392 VP.t3 VSUBS 2.66521f
C1393 VP.n3 VSUBS 0.060647f
C1394 VP.n4 VSUBS 0.03254f
C1395 VP.n5 VSUBS 0.041484f
C1396 VP.n6 VSUBS 0.042901f
C1397 VP.t0 VSUBS 2.66521f
C1398 VP.n7 VSUBS 0.038852f
C1399 VP.n8 VSUBS 0.306193f
C1400 VP.t4 VSUBS 2.66521f
C1401 VP.t5 VSUBS 2.89407f
C1402 VP.n9 VSUBS 1.00969f
C1403 VP.n10 VSUBS 1.04821f
C1404 VP.n11 VSUBS 0.060647f
C1405 VP.n12 VSUBS 0.055583f
C1406 VP.n13 VSUBS 0.03254f
C1407 VP.n14 VSUBS 0.03254f
C1408 VP.n15 VSUBS 0.03254f
C1409 VP.n16 VSUBS 0.061216f
C1410 VP.n17 VSUBS 0.041484f
C1411 VP.n18 VSUBS 1.03818f
C1412 VP.n19 VSUBS 1.71281f
C1413 VP.t1 VSUBS 2.66521f
C1414 VP.n20 VSUBS 1.03818f
C1415 VP.n21 VSUBS 1.73707f
C1416 VP.n22 VSUBS 0.042901f
C1417 VP.n23 VSUBS 0.03254f
C1418 VP.n24 VSUBS 0.061216f
C1419 VP.n25 VSUBS 0.038852f
C1420 VP.n26 VSUBS 0.055583f
C1421 VP.n27 VSUBS 0.03254f
C1422 VP.n28 VSUBS 0.03254f
C1423 VP.n29 VSUBS 0.03254f
C1424 VP.n30 VSUBS 0.97286f
C1425 VP.n31 VSUBS 0.060647f
C1426 VP.n32 VSUBS 0.055583f
C1427 VP.n33 VSUBS 0.03254f
C1428 VP.n34 VSUBS 0.03254f
C1429 VP.n35 VSUBS 0.03254f
C1430 VP.n36 VSUBS 0.061216f
C1431 VP.n37 VSUBS 0.041484f
C1432 VP.n38 VSUBS 1.03818f
C1433 VP.n39 VSUBS 0.051259f
.ends

