* NGSPICE file created from diff_pair_sample_0055.ext - technology: sky130A

.subckt diff_pair_sample_0055 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0 ps=0 w=2.14 l=1.26
X1 B.t8 B.t6 B.t7 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0 ps=0 w=2.14 l=1.26
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0.8346 ps=5.06 w=2.14 l=1.26
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0.8346 ps=5.06 w=2.14 l=1.26
X4 B.t5 B.t3 B.t4 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0 ps=0 w=2.14 l=1.26
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0.8346 ps=5.06 w=2.14 l=1.26
X6 B.t2 B.t0 B.t1 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0 ps=0 w=2.14 l=1.26
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1606_n1396# sky130_fd_pr__pfet_01v8 ad=0.8346 pd=5.06 as=0.8346 ps=5.06 w=2.14 l=1.26
R0 B.n157 B.n50 585
R1 B.n156 B.n155 585
R2 B.n154 B.n51 585
R3 B.n153 B.n152 585
R4 B.n151 B.n52 585
R5 B.n150 B.n149 585
R6 B.n148 B.n53 585
R7 B.n147 B.n146 585
R8 B.n145 B.n54 585
R9 B.n144 B.n143 585
R10 B.n142 B.n55 585
R11 B.n141 B.n140 585
R12 B.n139 B.n56 585
R13 B.n138 B.n137 585
R14 B.n133 B.n57 585
R15 B.n132 B.n131 585
R16 B.n130 B.n58 585
R17 B.n129 B.n128 585
R18 B.n127 B.n59 585
R19 B.n126 B.n125 585
R20 B.n124 B.n60 585
R21 B.n123 B.n122 585
R22 B.n120 B.n61 585
R23 B.n119 B.n118 585
R24 B.n117 B.n64 585
R25 B.n116 B.n115 585
R26 B.n114 B.n65 585
R27 B.n113 B.n112 585
R28 B.n111 B.n66 585
R29 B.n110 B.n109 585
R30 B.n108 B.n67 585
R31 B.n107 B.n106 585
R32 B.n105 B.n68 585
R33 B.n104 B.n103 585
R34 B.n102 B.n69 585
R35 B.n159 B.n158 585
R36 B.n160 B.n49 585
R37 B.n162 B.n161 585
R38 B.n163 B.n48 585
R39 B.n165 B.n164 585
R40 B.n166 B.n47 585
R41 B.n168 B.n167 585
R42 B.n169 B.n46 585
R43 B.n171 B.n170 585
R44 B.n172 B.n45 585
R45 B.n174 B.n173 585
R46 B.n175 B.n44 585
R47 B.n177 B.n176 585
R48 B.n178 B.n43 585
R49 B.n180 B.n179 585
R50 B.n181 B.n42 585
R51 B.n183 B.n182 585
R52 B.n184 B.n41 585
R53 B.n186 B.n185 585
R54 B.n187 B.n40 585
R55 B.n189 B.n188 585
R56 B.n190 B.n39 585
R57 B.n192 B.n191 585
R58 B.n193 B.n38 585
R59 B.n195 B.n194 585
R60 B.n196 B.n37 585
R61 B.n198 B.n197 585
R62 B.n199 B.n36 585
R63 B.n201 B.n200 585
R64 B.n202 B.n35 585
R65 B.n204 B.n203 585
R66 B.n205 B.n34 585
R67 B.n207 B.n206 585
R68 B.n208 B.n33 585
R69 B.n210 B.n209 585
R70 B.n211 B.n32 585
R71 B.n266 B.n265 585
R72 B.n264 B.n11 585
R73 B.n263 B.n262 585
R74 B.n261 B.n12 585
R75 B.n260 B.n259 585
R76 B.n258 B.n13 585
R77 B.n257 B.n256 585
R78 B.n255 B.n14 585
R79 B.n254 B.n253 585
R80 B.n252 B.n15 585
R81 B.n251 B.n250 585
R82 B.n249 B.n16 585
R83 B.n248 B.n247 585
R84 B.n245 B.n17 585
R85 B.n244 B.n243 585
R86 B.n242 B.n20 585
R87 B.n241 B.n240 585
R88 B.n239 B.n21 585
R89 B.n238 B.n237 585
R90 B.n236 B.n22 585
R91 B.n235 B.n234 585
R92 B.n233 B.n23 585
R93 B.n231 B.n230 585
R94 B.n229 B.n26 585
R95 B.n228 B.n227 585
R96 B.n226 B.n27 585
R97 B.n225 B.n224 585
R98 B.n223 B.n28 585
R99 B.n222 B.n221 585
R100 B.n220 B.n29 585
R101 B.n219 B.n218 585
R102 B.n217 B.n30 585
R103 B.n216 B.n215 585
R104 B.n214 B.n31 585
R105 B.n213 B.n212 585
R106 B.n267 B.n10 585
R107 B.n269 B.n268 585
R108 B.n270 B.n9 585
R109 B.n272 B.n271 585
R110 B.n273 B.n8 585
R111 B.n275 B.n274 585
R112 B.n276 B.n7 585
R113 B.n278 B.n277 585
R114 B.n279 B.n6 585
R115 B.n281 B.n280 585
R116 B.n282 B.n5 585
R117 B.n284 B.n283 585
R118 B.n285 B.n4 585
R119 B.n287 B.n286 585
R120 B.n288 B.n3 585
R121 B.n290 B.n289 585
R122 B.n291 B.n0 585
R123 B.n2 B.n1 585
R124 B.n78 B.n77 585
R125 B.n80 B.n79 585
R126 B.n81 B.n76 585
R127 B.n83 B.n82 585
R128 B.n84 B.n75 585
R129 B.n86 B.n85 585
R130 B.n87 B.n74 585
R131 B.n89 B.n88 585
R132 B.n90 B.n73 585
R133 B.n92 B.n91 585
R134 B.n93 B.n72 585
R135 B.n95 B.n94 585
R136 B.n96 B.n71 585
R137 B.n98 B.n97 585
R138 B.n99 B.n70 585
R139 B.n101 B.n100 585
R140 B.n100 B.n69 478.086
R141 B.n158 B.n157 478.086
R142 B.n212 B.n211 478.086
R143 B.n267 B.n266 478.086
R144 B.n293 B.n292 256.663
R145 B.n62 B.t0 245.351
R146 B.n134 B.t3 245.351
R147 B.n24 B.t6 245.351
R148 B.n18 B.t9 245.351
R149 B.n292 B.n291 235.042
R150 B.n292 B.n2 235.042
R151 B.n134 B.t4 202.935
R152 B.n24 B.t8 202.935
R153 B.n62 B.t1 202.935
R154 B.n18 B.t11 202.935
R155 B.n135 B.t5 172.099
R156 B.n25 B.t7 172.099
R157 B.n63 B.t2 172.099
R158 B.n19 B.t10 172.099
R159 B.n104 B.n69 163.367
R160 B.n105 B.n104 163.367
R161 B.n106 B.n105 163.367
R162 B.n106 B.n67 163.367
R163 B.n110 B.n67 163.367
R164 B.n111 B.n110 163.367
R165 B.n112 B.n111 163.367
R166 B.n112 B.n65 163.367
R167 B.n116 B.n65 163.367
R168 B.n117 B.n116 163.367
R169 B.n118 B.n117 163.367
R170 B.n118 B.n61 163.367
R171 B.n123 B.n61 163.367
R172 B.n124 B.n123 163.367
R173 B.n125 B.n124 163.367
R174 B.n125 B.n59 163.367
R175 B.n129 B.n59 163.367
R176 B.n130 B.n129 163.367
R177 B.n131 B.n130 163.367
R178 B.n131 B.n57 163.367
R179 B.n138 B.n57 163.367
R180 B.n139 B.n138 163.367
R181 B.n140 B.n139 163.367
R182 B.n140 B.n55 163.367
R183 B.n144 B.n55 163.367
R184 B.n145 B.n144 163.367
R185 B.n146 B.n145 163.367
R186 B.n146 B.n53 163.367
R187 B.n150 B.n53 163.367
R188 B.n151 B.n150 163.367
R189 B.n152 B.n151 163.367
R190 B.n152 B.n51 163.367
R191 B.n156 B.n51 163.367
R192 B.n157 B.n156 163.367
R193 B.n211 B.n210 163.367
R194 B.n210 B.n33 163.367
R195 B.n206 B.n33 163.367
R196 B.n206 B.n205 163.367
R197 B.n205 B.n204 163.367
R198 B.n204 B.n35 163.367
R199 B.n200 B.n35 163.367
R200 B.n200 B.n199 163.367
R201 B.n199 B.n198 163.367
R202 B.n198 B.n37 163.367
R203 B.n194 B.n37 163.367
R204 B.n194 B.n193 163.367
R205 B.n193 B.n192 163.367
R206 B.n192 B.n39 163.367
R207 B.n188 B.n39 163.367
R208 B.n188 B.n187 163.367
R209 B.n187 B.n186 163.367
R210 B.n186 B.n41 163.367
R211 B.n182 B.n41 163.367
R212 B.n182 B.n181 163.367
R213 B.n181 B.n180 163.367
R214 B.n180 B.n43 163.367
R215 B.n176 B.n43 163.367
R216 B.n176 B.n175 163.367
R217 B.n175 B.n174 163.367
R218 B.n174 B.n45 163.367
R219 B.n170 B.n45 163.367
R220 B.n170 B.n169 163.367
R221 B.n169 B.n168 163.367
R222 B.n168 B.n47 163.367
R223 B.n164 B.n47 163.367
R224 B.n164 B.n163 163.367
R225 B.n163 B.n162 163.367
R226 B.n162 B.n49 163.367
R227 B.n158 B.n49 163.367
R228 B.n266 B.n11 163.367
R229 B.n262 B.n11 163.367
R230 B.n262 B.n261 163.367
R231 B.n261 B.n260 163.367
R232 B.n260 B.n13 163.367
R233 B.n256 B.n13 163.367
R234 B.n256 B.n255 163.367
R235 B.n255 B.n254 163.367
R236 B.n254 B.n15 163.367
R237 B.n250 B.n15 163.367
R238 B.n250 B.n249 163.367
R239 B.n249 B.n248 163.367
R240 B.n248 B.n17 163.367
R241 B.n243 B.n17 163.367
R242 B.n243 B.n242 163.367
R243 B.n242 B.n241 163.367
R244 B.n241 B.n21 163.367
R245 B.n237 B.n21 163.367
R246 B.n237 B.n236 163.367
R247 B.n236 B.n235 163.367
R248 B.n235 B.n23 163.367
R249 B.n230 B.n23 163.367
R250 B.n230 B.n229 163.367
R251 B.n229 B.n228 163.367
R252 B.n228 B.n27 163.367
R253 B.n224 B.n27 163.367
R254 B.n224 B.n223 163.367
R255 B.n223 B.n222 163.367
R256 B.n222 B.n29 163.367
R257 B.n218 B.n29 163.367
R258 B.n218 B.n217 163.367
R259 B.n217 B.n216 163.367
R260 B.n216 B.n31 163.367
R261 B.n212 B.n31 163.367
R262 B.n268 B.n267 163.367
R263 B.n268 B.n9 163.367
R264 B.n272 B.n9 163.367
R265 B.n273 B.n272 163.367
R266 B.n274 B.n273 163.367
R267 B.n274 B.n7 163.367
R268 B.n278 B.n7 163.367
R269 B.n279 B.n278 163.367
R270 B.n280 B.n279 163.367
R271 B.n280 B.n5 163.367
R272 B.n284 B.n5 163.367
R273 B.n285 B.n284 163.367
R274 B.n286 B.n285 163.367
R275 B.n286 B.n3 163.367
R276 B.n290 B.n3 163.367
R277 B.n291 B.n290 163.367
R278 B.n77 B.n2 163.367
R279 B.n80 B.n77 163.367
R280 B.n81 B.n80 163.367
R281 B.n82 B.n81 163.367
R282 B.n82 B.n75 163.367
R283 B.n86 B.n75 163.367
R284 B.n87 B.n86 163.367
R285 B.n88 B.n87 163.367
R286 B.n88 B.n73 163.367
R287 B.n92 B.n73 163.367
R288 B.n93 B.n92 163.367
R289 B.n94 B.n93 163.367
R290 B.n94 B.n71 163.367
R291 B.n98 B.n71 163.367
R292 B.n99 B.n98 163.367
R293 B.n100 B.n99 163.367
R294 B.n121 B.n63 59.5399
R295 B.n136 B.n135 59.5399
R296 B.n232 B.n25 59.5399
R297 B.n246 B.n19 59.5399
R298 B.n265 B.n10 31.0639
R299 B.n213 B.n32 31.0639
R300 B.n159 B.n50 31.0639
R301 B.n102 B.n101 31.0639
R302 B.n63 B.n62 30.8369
R303 B.n135 B.n134 30.8369
R304 B.n25 B.n24 30.8369
R305 B.n19 B.n18 30.8369
R306 B B.n293 18.0485
R307 B.n269 B.n10 10.6151
R308 B.n270 B.n269 10.6151
R309 B.n271 B.n270 10.6151
R310 B.n271 B.n8 10.6151
R311 B.n275 B.n8 10.6151
R312 B.n276 B.n275 10.6151
R313 B.n277 B.n276 10.6151
R314 B.n277 B.n6 10.6151
R315 B.n281 B.n6 10.6151
R316 B.n282 B.n281 10.6151
R317 B.n283 B.n282 10.6151
R318 B.n283 B.n4 10.6151
R319 B.n287 B.n4 10.6151
R320 B.n288 B.n287 10.6151
R321 B.n289 B.n288 10.6151
R322 B.n289 B.n0 10.6151
R323 B.n265 B.n264 10.6151
R324 B.n264 B.n263 10.6151
R325 B.n263 B.n12 10.6151
R326 B.n259 B.n12 10.6151
R327 B.n259 B.n258 10.6151
R328 B.n258 B.n257 10.6151
R329 B.n257 B.n14 10.6151
R330 B.n253 B.n14 10.6151
R331 B.n253 B.n252 10.6151
R332 B.n252 B.n251 10.6151
R333 B.n251 B.n16 10.6151
R334 B.n247 B.n16 10.6151
R335 B.n245 B.n244 10.6151
R336 B.n244 B.n20 10.6151
R337 B.n240 B.n20 10.6151
R338 B.n240 B.n239 10.6151
R339 B.n239 B.n238 10.6151
R340 B.n238 B.n22 10.6151
R341 B.n234 B.n22 10.6151
R342 B.n234 B.n233 10.6151
R343 B.n231 B.n26 10.6151
R344 B.n227 B.n26 10.6151
R345 B.n227 B.n226 10.6151
R346 B.n226 B.n225 10.6151
R347 B.n225 B.n28 10.6151
R348 B.n221 B.n28 10.6151
R349 B.n221 B.n220 10.6151
R350 B.n220 B.n219 10.6151
R351 B.n219 B.n30 10.6151
R352 B.n215 B.n30 10.6151
R353 B.n215 B.n214 10.6151
R354 B.n214 B.n213 10.6151
R355 B.n209 B.n32 10.6151
R356 B.n209 B.n208 10.6151
R357 B.n208 B.n207 10.6151
R358 B.n207 B.n34 10.6151
R359 B.n203 B.n34 10.6151
R360 B.n203 B.n202 10.6151
R361 B.n202 B.n201 10.6151
R362 B.n201 B.n36 10.6151
R363 B.n197 B.n36 10.6151
R364 B.n197 B.n196 10.6151
R365 B.n196 B.n195 10.6151
R366 B.n195 B.n38 10.6151
R367 B.n191 B.n38 10.6151
R368 B.n191 B.n190 10.6151
R369 B.n190 B.n189 10.6151
R370 B.n189 B.n40 10.6151
R371 B.n185 B.n40 10.6151
R372 B.n185 B.n184 10.6151
R373 B.n184 B.n183 10.6151
R374 B.n183 B.n42 10.6151
R375 B.n179 B.n42 10.6151
R376 B.n179 B.n178 10.6151
R377 B.n178 B.n177 10.6151
R378 B.n177 B.n44 10.6151
R379 B.n173 B.n44 10.6151
R380 B.n173 B.n172 10.6151
R381 B.n172 B.n171 10.6151
R382 B.n171 B.n46 10.6151
R383 B.n167 B.n46 10.6151
R384 B.n167 B.n166 10.6151
R385 B.n166 B.n165 10.6151
R386 B.n165 B.n48 10.6151
R387 B.n161 B.n48 10.6151
R388 B.n161 B.n160 10.6151
R389 B.n160 B.n159 10.6151
R390 B.n78 B.n1 10.6151
R391 B.n79 B.n78 10.6151
R392 B.n79 B.n76 10.6151
R393 B.n83 B.n76 10.6151
R394 B.n84 B.n83 10.6151
R395 B.n85 B.n84 10.6151
R396 B.n85 B.n74 10.6151
R397 B.n89 B.n74 10.6151
R398 B.n90 B.n89 10.6151
R399 B.n91 B.n90 10.6151
R400 B.n91 B.n72 10.6151
R401 B.n95 B.n72 10.6151
R402 B.n96 B.n95 10.6151
R403 B.n97 B.n96 10.6151
R404 B.n97 B.n70 10.6151
R405 B.n101 B.n70 10.6151
R406 B.n103 B.n102 10.6151
R407 B.n103 B.n68 10.6151
R408 B.n107 B.n68 10.6151
R409 B.n108 B.n107 10.6151
R410 B.n109 B.n108 10.6151
R411 B.n109 B.n66 10.6151
R412 B.n113 B.n66 10.6151
R413 B.n114 B.n113 10.6151
R414 B.n115 B.n114 10.6151
R415 B.n115 B.n64 10.6151
R416 B.n119 B.n64 10.6151
R417 B.n120 B.n119 10.6151
R418 B.n122 B.n60 10.6151
R419 B.n126 B.n60 10.6151
R420 B.n127 B.n126 10.6151
R421 B.n128 B.n127 10.6151
R422 B.n128 B.n58 10.6151
R423 B.n132 B.n58 10.6151
R424 B.n133 B.n132 10.6151
R425 B.n137 B.n133 10.6151
R426 B.n141 B.n56 10.6151
R427 B.n142 B.n141 10.6151
R428 B.n143 B.n142 10.6151
R429 B.n143 B.n54 10.6151
R430 B.n147 B.n54 10.6151
R431 B.n148 B.n147 10.6151
R432 B.n149 B.n148 10.6151
R433 B.n149 B.n52 10.6151
R434 B.n153 B.n52 10.6151
R435 B.n154 B.n153 10.6151
R436 B.n155 B.n154 10.6151
R437 B.n155 B.n50 10.6151
R438 B.n293 B.n0 8.11757
R439 B.n293 B.n1 8.11757
R440 B.n246 B.n245 6.5566
R441 B.n233 B.n232 6.5566
R442 B.n122 B.n121 6.5566
R443 B.n137 B.n136 6.5566
R444 B.n247 B.n246 4.05904
R445 B.n232 B.n231 4.05904
R446 B.n121 B.n120 4.05904
R447 B.n136 B.n56 4.05904
R448 VN VN.t0 187.013
R449 VN VN.t1 153.242
R450 VTAIL.n3 VTAIL.t2 171.29
R451 VTAIL.n0 VTAIL.t1 171.29
R452 VTAIL.n2 VTAIL.t0 171.29
R453 VTAIL.n1 VTAIL.t3 171.29
R454 VTAIL.n1 VTAIL.n0 16.9531
R455 VTAIL.n3 VTAIL.n2 15.5824
R456 VTAIL.n2 VTAIL.n1 1.15567
R457 VTAIL VTAIL.n0 0.87119
R458 VTAIL VTAIL.n3 0.284983
R459 VDD2.n0 VDD2.t0 216.214
R460 VDD2.n0 VDD2.t1 187.968
R461 VDD2 VDD2.n0 0.401362
R462 VP.n0 VP.t0 186.728
R463 VP.n0 VP.t1 153.095
R464 VP VP.n0 0.146778
R465 VDD1 VDD1.t0 217.082
R466 VDD1 VDD1.t1 188.369
C0 B w_n1606_n1396# 4.59207f
C1 VDD1 w_n1606_n1396# 0.916152f
C2 B VDD1 0.765889f
C3 VN w_n1606_n1396# 1.88882f
C4 VP w_n1606_n1396# 2.0864f
C5 B VN 0.684181f
C6 B VP 1.00969f
C7 VN VDD1 0.153276f
C8 VP VDD1 0.755215f
C9 VDD2 w_n1606_n1396# 0.925686f
C10 VTAIL w_n1606_n1396# 1.25045f
C11 B VDD2 0.784688f
C12 VP VN 3.01182f
C13 VDD1 VDD2 0.517704f
C14 B VTAIL 1.04024f
C15 VDD1 VTAIL 2.08388f
C16 VN VDD2 0.627858f
C17 VP VDD2 0.282172f
C18 VN VTAIL 0.727913f
C19 VP VTAIL 0.742083f
C20 VDD2 VTAIL 2.12734f
C21 VDD2 VSUBS 0.44135f
C22 VDD1 VSUBS 2.195879f
C23 VTAIL VSUBS 0.325619f
C24 VN VSUBS 3.45648f
C25 VP VSUBS 0.825902f
C26 B VSUBS 1.970175f
C27 w_n1606_n1396# VSUBS 28.580399f
C28 VDD1.t1 VSUBS 0.184273f
C29 VDD1.t0 VSUBS 0.28085f
C30 VP.t0 VSUBS 0.999219f
C31 VP.t1 VSUBS 0.665543f
C32 VP.n0 VSUBS 3.38193f
C33 VDD2.t0 VSUBS 0.280775f
C34 VDD2.t1 VSUBS 0.189139f
C35 VDD2.n0 VSUBS 1.57199f
C36 VTAIL.t1 VSUBS 0.21013f
C37 VTAIL.n0 VSUBS 0.866071f
C38 VTAIL.t3 VSUBS 0.21013f
C39 VTAIL.n1 VSUBS 0.884664f
C40 VTAIL.t0 VSUBS 0.210129f
C41 VTAIL.n2 VSUBS 0.795076f
C42 VTAIL.t2 VSUBS 0.21013f
C43 VTAIL.n3 VSUBS 0.738167f
C44 VN.t1 VSUBS 0.385263f
C45 VN.t0 VSUBS 0.58325f
C46 B.n0 VSUBS 0.007945f
C47 B.n1 VSUBS 0.007945f
C48 B.n2 VSUBS 0.011751f
C49 B.n3 VSUBS 0.009005f
C50 B.n4 VSUBS 0.009005f
C51 B.n5 VSUBS 0.009005f
C52 B.n6 VSUBS 0.009005f
C53 B.n7 VSUBS 0.009005f
C54 B.n8 VSUBS 0.009005f
C55 B.n9 VSUBS 0.009005f
C56 B.n10 VSUBS 0.019807f
C57 B.n11 VSUBS 0.009005f
C58 B.n12 VSUBS 0.009005f
C59 B.n13 VSUBS 0.009005f
C60 B.n14 VSUBS 0.009005f
C61 B.n15 VSUBS 0.009005f
C62 B.n16 VSUBS 0.009005f
C63 B.n17 VSUBS 0.009005f
C64 B.t10 VSUBS 0.060382f
C65 B.t11 VSUBS 0.068963f
C66 B.t9 VSUBS 0.167634f
C67 B.n18 VSUBS 0.078415f
C68 B.n19 VSUBS 0.069312f
C69 B.n20 VSUBS 0.009005f
C70 B.n21 VSUBS 0.009005f
C71 B.n22 VSUBS 0.009005f
C72 B.n23 VSUBS 0.009005f
C73 B.t7 VSUBS 0.060382f
C74 B.t8 VSUBS 0.068963f
C75 B.t6 VSUBS 0.167634f
C76 B.n24 VSUBS 0.078415f
C77 B.n25 VSUBS 0.069312f
C78 B.n26 VSUBS 0.009005f
C79 B.n27 VSUBS 0.009005f
C80 B.n28 VSUBS 0.009005f
C81 B.n29 VSUBS 0.009005f
C82 B.n30 VSUBS 0.009005f
C83 B.n31 VSUBS 0.009005f
C84 B.n32 VSUBS 0.019807f
C85 B.n33 VSUBS 0.009005f
C86 B.n34 VSUBS 0.009005f
C87 B.n35 VSUBS 0.009005f
C88 B.n36 VSUBS 0.009005f
C89 B.n37 VSUBS 0.009005f
C90 B.n38 VSUBS 0.009005f
C91 B.n39 VSUBS 0.009005f
C92 B.n40 VSUBS 0.009005f
C93 B.n41 VSUBS 0.009005f
C94 B.n42 VSUBS 0.009005f
C95 B.n43 VSUBS 0.009005f
C96 B.n44 VSUBS 0.009005f
C97 B.n45 VSUBS 0.009005f
C98 B.n46 VSUBS 0.009005f
C99 B.n47 VSUBS 0.009005f
C100 B.n48 VSUBS 0.009005f
C101 B.n49 VSUBS 0.009005f
C102 B.n50 VSUBS 0.019861f
C103 B.n51 VSUBS 0.009005f
C104 B.n52 VSUBS 0.009005f
C105 B.n53 VSUBS 0.009005f
C106 B.n54 VSUBS 0.009005f
C107 B.n55 VSUBS 0.009005f
C108 B.n56 VSUBS 0.006224f
C109 B.n57 VSUBS 0.009005f
C110 B.n58 VSUBS 0.009005f
C111 B.n59 VSUBS 0.009005f
C112 B.n60 VSUBS 0.009005f
C113 B.n61 VSUBS 0.009005f
C114 B.t2 VSUBS 0.060382f
C115 B.t1 VSUBS 0.068963f
C116 B.t0 VSUBS 0.167634f
C117 B.n62 VSUBS 0.078415f
C118 B.n63 VSUBS 0.069312f
C119 B.n64 VSUBS 0.009005f
C120 B.n65 VSUBS 0.009005f
C121 B.n66 VSUBS 0.009005f
C122 B.n67 VSUBS 0.009005f
C123 B.n68 VSUBS 0.009005f
C124 B.n69 VSUBS 0.02098f
C125 B.n70 VSUBS 0.009005f
C126 B.n71 VSUBS 0.009005f
C127 B.n72 VSUBS 0.009005f
C128 B.n73 VSUBS 0.009005f
C129 B.n74 VSUBS 0.009005f
C130 B.n75 VSUBS 0.009005f
C131 B.n76 VSUBS 0.009005f
C132 B.n77 VSUBS 0.009005f
C133 B.n78 VSUBS 0.009005f
C134 B.n79 VSUBS 0.009005f
C135 B.n80 VSUBS 0.009005f
C136 B.n81 VSUBS 0.009005f
C137 B.n82 VSUBS 0.009005f
C138 B.n83 VSUBS 0.009005f
C139 B.n84 VSUBS 0.009005f
C140 B.n85 VSUBS 0.009005f
C141 B.n86 VSUBS 0.009005f
C142 B.n87 VSUBS 0.009005f
C143 B.n88 VSUBS 0.009005f
C144 B.n89 VSUBS 0.009005f
C145 B.n90 VSUBS 0.009005f
C146 B.n91 VSUBS 0.009005f
C147 B.n92 VSUBS 0.009005f
C148 B.n93 VSUBS 0.009005f
C149 B.n94 VSUBS 0.009005f
C150 B.n95 VSUBS 0.009005f
C151 B.n96 VSUBS 0.009005f
C152 B.n97 VSUBS 0.009005f
C153 B.n98 VSUBS 0.009005f
C154 B.n99 VSUBS 0.009005f
C155 B.n100 VSUBS 0.019807f
C156 B.n101 VSUBS 0.019807f
C157 B.n102 VSUBS 0.02098f
C158 B.n103 VSUBS 0.009005f
C159 B.n104 VSUBS 0.009005f
C160 B.n105 VSUBS 0.009005f
C161 B.n106 VSUBS 0.009005f
C162 B.n107 VSUBS 0.009005f
C163 B.n108 VSUBS 0.009005f
C164 B.n109 VSUBS 0.009005f
C165 B.n110 VSUBS 0.009005f
C166 B.n111 VSUBS 0.009005f
C167 B.n112 VSUBS 0.009005f
C168 B.n113 VSUBS 0.009005f
C169 B.n114 VSUBS 0.009005f
C170 B.n115 VSUBS 0.009005f
C171 B.n116 VSUBS 0.009005f
C172 B.n117 VSUBS 0.009005f
C173 B.n118 VSUBS 0.009005f
C174 B.n119 VSUBS 0.009005f
C175 B.n120 VSUBS 0.006224f
C176 B.n121 VSUBS 0.020863f
C177 B.n122 VSUBS 0.007283f
C178 B.n123 VSUBS 0.009005f
C179 B.n124 VSUBS 0.009005f
C180 B.n125 VSUBS 0.009005f
C181 B.n126 VSUBS 0.009005f
C182 B.n127 VSUBS 0.009005f
C183 B.n128 VSUBS 0.009005f
C184 B.n129 VSUBS 0.009005f
C185 B.n130 VSUBS 0.009005f
C186 B.n131 VSUBS 0.009005f
C187 B.n132 VSUBS 0.009005f
C188 B.n133 VSUBS 0.009005f
C189 B.t5 VSUBS 0.060382f
C190 B.t4 VSUBS 0.068963f
C191 B.t3 VSUBS 0.167634f
C192 B.n134 VSUBS 0.078415f
C193 B.n135 VSUBS 0.069312f
C194 B.n136 VSUBS 0.020863f
C195 B.n137 VSUBS 0.007283f
C196 B.n138 VSUBS 0.009005f
C197 B.n139 VSUBS 0.009005f
C198 B.n140 VSUBS 0.009005f
C199 B.n141 VSUBS 0.009005f
C200 B.n142 VSUBS 0.009005f
C201 B.n143 VSUBS 0.009005f
C202 B.n144 VSUBS 0.009005f
C203 B.n145 VSUBS 0.009005f
C204 B.n146 VSUBS 0.009005f
C205 B.n147 VSUBS 0.009005f
C206 B.n148 VSUBS 0.009005f
C207 B.n149 VSUBS 0.009005f
C208 B.n150 VSUBS 0.009005f
C209 B.n151 VSUBS 0.009005f
C210 B.n152 VSUBS 0.009005f
C211 B.n153 VSUBS 0.009005f
C212 B.n154 VSUBS 0.009005f
C213 B.n155 VSUBS 0.009005f
C214 B.n156 VSUBS 0.009005f
C215 B.n157 VSUBS 0.02098f
C216 B.n158 VSUBS 0.019807f
C217 B.n159 VSUBS 0.020925f
C218 B.n160 VSUBS 0.009005f
C219 B.n161 VSUBS 0.009005f
C220 B.n162 VSUBS 0.009005f
C221 B.n163 VSUBS 0.009005f
C222 B.n164 VSUBS 0.009005f
C223 B.n165 VSUBS 0.009005f
C224 B.n166 VSUBS 0.009005f
C225 B.n167 VSUBS 0.009005f
C226 B.n168 VSUBS 0.009005f
C227 B.n169 VSUBS 0.009005f
C228 B.n170 VSUBS 0.009005f
C229 B.n171 VSUBS 0.009005f
C230 B.n172 VSUBS 0.009005f
C231 B.n173 VSUBS 0.009005f
C232 B.n174 VSUBS 0.009005f
C233 B.n175 VSUBS 0.009005f
C234 B.n176 VSUBS 0.009005f
C235 B.n177 VSUBS 0.009005f
C236 B.n178 VSUBS 0.009005f
C237 B.n179 VSUBS 0.009005f
C238 B.n180 VSUBS 0.009005f
C239 B.n181 VSUBS 0.009005f
C240 B.n182 VSUBS 0.009005f
C241 B.n183 VSUBS 0.009005f
C242 B.n184 VSUBS 0.009005f
C243 B.n185 VSUBS 0.009005f
C244 B.n186 VSUBS 0.009005f
C245 B.n187 VSUBS 0.009005f
C246 B.n188 VSUBS 0.009005f
C247 B.n189 VSUBS 0.009005f
C248 B.n190 VSUBS 0.009005f
C249 B.n191 VSUBS 0.009005f
C250 B.n192 VSUBS 0.009005f
C251 B.n193 VSUBS 0.009005f
C252 B.n194 VSUBS 0.009005f
C253 B.n195 VSUBS 0.009005f
C254 B.n196 VSUBS 0.009005f
C255 B.n197 VSUBS 0.009005f
C256 B.n198 VSUBS 0.009005f
C257 B.n199 VSUBS 0.009005f
C258 B.n200 VSUBS 0.009005f
C259 B.n201 VSUBS 0.009005f
C260 B.n202 VSUBS 0.009005f
C261 B.n203 VSUBS 0.009005f
C262 B.n204 VSUBS 0.009005f
C263 B.n205 VSUBS 0.009005f
C264 B.n206 VSUBS 0.009005f
C265 B.n207 VSUBS 0.009005f
C266 B.n208 VSUBS 0.009005f
C267 B.n209 VSUBS 0.009005f
C268 B.n210 VSUBS 0.009005f
C269 B.n211 VSUBS 0.019807f
C270 B.n212 VSUBS 0.02098f
C271 B.n213 VSUBS 0.02098f
C272 B.n214 VSUBS 0.009005f
C273 B.n215 VSUBS 0.009005f
C274 B.n216 VSUBS 0.009005f
C275 B.n217 VSUBS 0.009005f
C276 B.n218 VSUBS 0.009005f
C277 B.n219 VSUBS 0.009005f
C278 B.n220 VSUBS 0.009005f
C279 B.n221 VSUBS 0.009005f
C280 B.n222 VSUBS 0.009005f
C281 B.n223 VSUBS 0.009005f
C282 B.n224 VSUBS 0.009005f
C283 B.n225 VSUBS 0.009005f
C284 B.n226 VSUBS 0.009005f
C285 B.n227 VSUBS 0.009005f
C286 B.n228 VSUBS 0.009005f
C287 B.n229 VSUBS 0.009005f
C288 B.n230 VSUBS 0.009005f
C289 B.n231 VSUBS 0.006224f
C290 B.n232 VSUBS 0.020863f
C291 B.n233 VSUBS 0.007283f
C292 B.n234 VSUBS 0.009005f
C293 B.n235 VSUBS 0.009005f
C294 B.n236 VSUBS 0.009005f
C295 B.n237 VSUBS 0.009005f
C296 B.n238 VSUBS 0.009005f
C297 B.n239 VSUBS 0.009005f
C298 B.n240 VSUBS 0.009005f
C299 B.n241 VSUBS 0.009005f
C300 B.n242 VSUBS 0.009005f
C301 B.n243 VSUBS 0.009005f
C302 B.n244 VSUBS 0.009005f
C303 B.n245 VSUBS 0.007283f
C304 B.n246 VSUBS 0.020863f
C305 B.n247 VSUBS 0.006224f
C306 B.n248 VSUBS 0.009005f
C307 B.n249 VSUBS 0.009005f
C308 B.n250 VSUBS 0.009005f
C309 B.n251 VSUBS 0.009005f
C310 B.n252 VSUBS 0.009005f
C311 B.n253 VSUBS 0.009005f
C312 B.n254 VSUBS 0.009005f
C313 B.n255 VSUBS 0.009005f
C314 B.n256 VSUBS 0.009005f
C315 B.n257 VSUBS 0.009005f
C316 B.n258 VSUBS 0.009005f
C317 B.n259 VSUBS 0.009005f
C318 B.n260 VSUBS 0.009005f
C319 B.n261 VSUBS 0.009005f
C320 B.n262 VSUBS 0.009005f
C321 B.n263 VSUBS 0.009005f
C322 B.n264 VSUBS 0.009005f
C323 B.n265 VSUBS 0.02098f
C324 B.n266 VSUBS 0.02098f
C325 B.n267 VSUBS 0.019807f
C326 B.n268 VSUBS 0.009005f
C327 B.n269 VSUBS 0.009005f
C328 B.n270 VSUBS 0.009005f
C329 B.n271 VSUBS 0.009005f
C330 B.n272 VSUBS 0.009005f
C331 B.n273 VSUBS 0.009005f
C332 B.n274 VSUBS 0.009005f
C333 B.n275 VSUBS 0.009005f
C334 B.n276 VSUBS 0.009005f
C335 B.n277 VSUBS 0.009005f
C336 B.n278 VSUBS 0.009005f
C337 B.n279 VSUBS 0.009005f
C338 B.n280 VSUBS 0.009005f
C339 B.n281 VSUBS 0.009005f
C340 B.n282 VSUBS 0.009005f
C341 B.n283 VSUBS 0.009005f
C342 B.n284 VSUBS 0.009005f
C343 B.n285 VSUBS 0.009005f
C344 B.n286 VSUBS 0.009005f
C345 B.n287 VSUBS 0.009005f
C346 B.n288 VSUBS 0.009005f
C347 B.n289 VSUBS 0.009005f
C348 B.n290 VSUBS 0.009005f
C349 B.n291 VSUBS 0.011751f
C350 B.n292 VSUBS 0.012518f
C351 B.n293 VSUBS 0.024892f
.ends

