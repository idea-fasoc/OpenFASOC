* NGSPICE file created from diff_pair_sample_0907.ext - technology: sky130A

.subckt diff_pair_sample_0907 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VP.t0 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X1 VTAIL.t13 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X2 VDD1.t5 VP.t1 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X3 VDD1.t7 VP.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=4.2432 ps=22.54 w=10.88 l=1
X4 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=1
X5 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=1
X6 VTAIL.t9 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=1.7952 ps=11.21 w=10.88 l=1
X7 VDD2.t6 VN.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=4.2432 ps=22.54 w=10.88 l=1
X8 VTAIL.t8 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=1
X10 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X11 VDD1.t4 VP.t5 VTAIL.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=4.2432 ps=22.54 w=10.88 l=1
X12 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=1
X14 VTAIL.t4 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
X15 VTAIL.t15 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=1.7952 ps=11.21 w=10.88 l=1
X16 VTAIL.t0 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=1.7952 ps=11.21 w=10.88 l=1
X17 VTAIL.t6 VP.t6 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=4.2432 pd=22.54 as=1.7952 ps=11.21 w=10.88 l=1
X18 VDD2.t0 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=4.2432 ps=22.54 w=10.88 l=1
X19 VDD1.t1 VP.t7 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=11.21 as=1.7952 ps=11.21 w=10.88 l=1
R0 VP.n5 VP.t6 317.216
R1 VP.n17 VP.t3 301.974
R2 VP.n27 VP.t5 301.974
R3 VP.n14 VP.t2 301.974
R4 VP.n19 VP.t7 262.209
R5 VP.n25 VP.t4 262.209
R6 VP.n12 VP.t0 262.209
R7 VP.n6 VP.t1 262.209
R8 VP.n8 VP.n7 161.3
R9 VP.n9 VP.n4 161.3
R10 VP.n11 VP.n10 161.3
R11 VP.n13 VP.n3 161.3
R12 VP.n26 VP.n0 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n22 VP.n1 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n18 VP.n2 161.3
R17 VP.n15 VP.n14 80.6037
R18 VP.n28 VP.n27 80.6037
R19 VP.n17 VP.n16 80.6037
R20 VP.n18 VP.n17 56.2338
R21 VP.n27 VP.n26 56.2338
R22 VP.n14 VP.n13 56.2338
R23 VP.n6 VP.n5 46.7059
R24 VP.n8 VP.n5 43.9111
R25 VP.n16 VP.n15 42.7741
R26 VP.n20 VP.n1 40.4106
R27 VP.n24 VP.n1 40.4106
R28 VP.n11 VP.n4 40.4106
R29 VP.n7 VP.n4 40.4106
R30 VP.n19 VP.n18 16.3106
R31 VP.n26 VP.n25 16.3106
R32 VP.n13 VP.n12 16.3106
R33 VP.n20 VP.n19 8.03383
R34 VP.n25 VP.n24 8.03383
R35 VP.n12 VP.n11 8.03383
R36 VP.n7 VP.n6 8.03383
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VDD1 VDD1.n0 65.9554
R49 VDD1.n3 VDD1.n2 65.8408
R50 VDD1.n3 VDD1.n1 65.8408
R51 VDD1.n5 VDD1.n4 65.3228
R52 VDD1.n5 VDD1.n3 38.8371
R53 VDD1.n4 VDD1.t6 1.82035
R54 VDD1.n4 VDD1.t7 1.82035
R55 VDD1.n0 VDD1.t2 1.82035
R56 VDD1.n0 VDD1.t5 1.82035
R57 VDD1.n2 VDD1.t3 1.82035
R58 VDD1.n2 VDD1.t4 1.82035
R59 VDD1.n1 VDD1.t0 1.82035
R60 VDD1.n1 VDD1.t1 1.82035
R61 VDD1 VDD1.n5 0.515586
R62 VTAIL.n11 VTAIL.t6 50.465
R63 VTAIL.n10 VTAIL.t14 50.465
R64 VTAIL.n7 VTAIL.t0 50.465
R65 VTAIL.n15 VTAIL.t1 50.464
R66 VTAIL.n2 VTAIL.t15 50.464
R67 VTAIL.n3 VTAIL.t7 50.464
R68 VTAIL.n6 VTAIL.t9 50.464
R69 VTAIL.n14 VTAIL.t10 50.4638
R70 VTAIL.n13 VTAIL.n12 48.6452
R71 VTAIL.n9 VTAIL.n8 48.6452
R72 VTAIL.n1 VTAIL.n0 48.6441
R73 VTAIL.n5 VTAIL.n4 48.6441
R74 VTAIL.n15 VTAIL.n14 22.8927
R75 VTAIL.n7 VTAIL.n6 22.8927
R76 VTAIL.n0 VTAIL.t3 1.82035
R77 VTAIL.n0 VTAIL.t13 1.82035
R78 VTAIL.n4 VTAIL.t5 1.82035
R79 VTAIL.n4 VTAIL.t8 1.82035
R80 VTAIL.n12 VTAIL.t11 1.82035
R81 VTAIL.n12 VTAIL.t12 1.82035
R82 VTAIL.n8 VTAIL.t2 1.82035
R83 VTAIL.n8 VTAIL.t4 1.82035
R84 VTAIL.n9 VTAIL.n7 1.14705
R85 VTAIL.n10 VTAIL.n9 1.14705
R86 VTAIL.n13 VTAIL.n11 1.14705
R87 VTAIL.n14 VTAIL.n13 1.14705
R88 VTAIL.n6 VTAIL.n5 1.14705
R89 VTAIL.n5 VTAIL.n3 1.14705
R90 VTAIL.n2 VTAIL.n1 1.14705
R91 VTAIL VTAIL.n15 1.08886
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 B.n659 B.n658 585
R96 B.n267 B.n95 585
R97 B.n266 B.n265 585
R98 B.n264 B.n263 585
R99 B.n262 B.n261 585
R100 B.n260 B.n259 585
R101 B.n258 B.n257 585
R102 B.n256 B.n255 585
R103 B.n254 B.n253 585
R104 B.n252 B.n251 585
R105 B.n250 B.n249 585
R106 B.n248 B.n247 585
R107 B.n246 B.n245 585
R108 B.n244 B.n243 585
R109 B.n242 B.n241 585
R110 B.n240 B.n239 585
R111 B.n238 B.n237 585
R112 B.n236 B.n235 585
R113 B.n234 B.n233 585
R114 B.n232 B.n231 585
R115 B.n230 B.n229 585
R116 B.n228 B.n227 585
R117 B.n226 B.n225 585
R118 B.n224 B.n223 585
R119 B.n222 B.n221 585
R120 B.n220 B.n219 585
R121 B.n218 B.n217 585
R122 B.n216 B.n215 585
R123 B.n214 B.n213 585
R124 B.n212 B.n211 585
R125 B.n210 B.n209 585
R126 B.n208 B.n207 585
R127 B.n206 B.n205 585
R128 B.n204 B.n203 585
R129 B.n202 B.n201 585
R130 B.n200 B.n199 585
R131 B.n198 B.n197 585
R132 B.n196 B.n195 585
R133 B.n194 B.n193 585
R134 B.n192 B.n191 585
R135 B.n190 B.n189 585
R136 B.n188 B.n187 585
R137 B.n186 B.n185 585
R138 B.n184 B.n183 585
R139 B.n182 B.n181 585
R140 B.n180 B.n179 585
R141 B.n178 B.n177 585
R142 B.n176 B.n175 585
R143 B.n174 B.n173 585
R144 B.n172 B.n171 585
R145 B.n170 B.n169 585
R146 B.n168 B.n167 585
R147 B.n166 B.n165 585
R148 B.n164 B.n163 585
R149 B.n162 B.n161 585
R150 B.n160 B.n159 585
R151 B.n158 B.n157 585
R152 B.n156 B.n155 585
R153 B.n154 B.n153 585
R154 B.n152 B.n151 585
R155 B.n150 B.n149 585
R156 B.n148 B.n147 585
R157 B.n146 B.n145 585
R158 B.n144 B.n143 585
R159 B.n142 B.n141 585
R160 B.n140 B.n139 585
R161 B.n138 B.n137 585
R162 B.n136 B.n135 585
R163 B.n134 B.n133 585
R164 B.n132 B.n131 585
R165 B.n130 B.n129 585
R166 B.n128 B.n127 585
R167 B.n126 B.n125 585
R168 B.n124 B.n123 585
R169 B.n122 B.n121 585
R170 B.n120 B.n119 585
R171 B.n118 B.n117 585
R172 B.n116 B.n115 585
R173 B.n114 B.n113 585
R174 B.n112 B.n111 585
R175 B.n110 B.n109 585
R176 B.n108 B.n107 585
R177 B.n106 B.n105 585
R178 B.n104 B.n103 585
R179 B.n53 B.n52 585
R180 B.n664 B.n663 585
R181 B.n657 B.n96 585
R182 B.n96 B.n50 585
R183 B.n656 B.n49 585
R184 B.n668 B.n49 585
R185 B.n655 B.n48 585
R186 B.n669 B.n48 585
R187 B.n654 B.n47 585
R188 B.n670 B.n47 585
R189 B.n653 B.n652 585
R190 B.n652 B.n43 585
R191 B.n651 B.n42 585
R192 B.n676 B.n42 585
R193 B.n650 B.n41 585
R194 B.n677 B.n41 585
R195 B.n649 B.n40 585
R196 B.n678 B.n40 585
R197 B.n648 B.n647 585
R198 B.n647 B.n36 585
R199 B.n646 B.n35 585
R200 B.n684 B.n35 585
R201 B.n645 B.n34 585
R202 B.n685 B.n34 585
R203 B.n644 B.n33 585
R204 B.n686 B.n33 585
R205 B.n643 B.n642 585
R206 B.n642 B.n32 585
R207 B.n641 B.n28 585
R208 B.n692 B.n28 585
R209 B.n640 B.n27 585
R210 B.n693 B.n27 585
R211 B.n639 B.n26 585
R212 B.n694 B.n26 585
R213 B.n638 B.n637 585
R214 B.n637 B.n25 585
R215 B.n636 B.n21 585
R216 B.n700 B.n21 585
R217 B.n635 B.n20 585
R218 B.n701 B.n20 585
R219 B.n634 B.n19 585
R220 B.n702 B.n19 585
R221 B.n633 B.n632 585
R222 B.n632 B.n18 585
R223 B.n631 B.n14 585
R224 B.n708 B.n14 585
R225 B.n630 B.n13 585
R226 B.n709 B.n13 585
R227 B.n629 B.n12 585
R228 B.n710 B.n12 585
R229 B.n628 B.n627 585
R230 B.n627 B.n626 585
R231 B.n625 B.n624 585
R232 B.n625 B.n8 585
R233 B.n623 B.n7 585
R234 B.n717 B.n7 585
R235 B.n622 B.n6 585
R236 B.n718 B.n6 585
R237 B.n621 B.n5 585
R238 B.n719 B.n5 585
R239 B.n620 B.n619 585
R240 B.n619 B.n4 585
R241 B.n618 B.n268 585
R242 B.n618 B.n617 585
R243 B.n608 B.n269 585
R244 B.n270 B.n269 585
R245 B.n610 B.n609 585
R246 B.n611 B.n610 585
R247 B.n607 B.n275 585
R248 B.n275 B.n274 585
R249 B.n606 B.n605 585
R250 B.n605 B.n604 585
R251 B.n277 B.n276 585
R252 B.n597 B.n277 585
R253 B.n596 B.n595 585
R254 B.n598 B.n596 585
R255 B.n594 B.n282 585
R256 B.n282 B.n281 585
R257 B.n593 B.n592 585
R258 B.n592 B.n591 585
R259 B.n284 B.n283 585
R260 B.n584 B.n284 585
R261 B.n583 B.n582 585
R262 B.n585 B.n583 585
R263 B.n581 B.n289 585
R264 B.n289 B.n288 585
R265 B.n580 B.n579 585
R266 B.n579 B.n578 585
R267 B.n291 B.n290 585
R268 B.n571 B.n291 585
R269 B.n570 B.n569 585
R270 B.n572 B.n570 585
R271 B.n568 B.n296 585
R272 B.n296 B.n295 585
R273 B.n567 B.n566 585
R274 B.n566 B.n565 585
R275 B.n298 B.n297 585
R276 B.n299 B.n298 585
R277 B.n558 B.n557 585
R278 B.n559 B.n558 585
R279 B.n556 B.n304 585
R280 B.n304 B.n303 585
R281 B.n555 B.n554 585
R282 B.n554 B.n553 585
R283 B.n306 B.n305 585
R284 B.n307 B.n306 585
R285 B.n546 B.n545 585
R286 B.n547 B.n546 585
R287 B.n544 B.n312 585
R288 B.n312 B.n311 585
R289 B.n543 B.n542 585
R290 B.n542 B.n541 585
R291 B.n314 B.n313 585
R292 B.n315 B.n314 585
R293 B.n537 B.n536 585
R294 B.n318 B.n317 585
R295 B.n533 B.n532 585
R296 B.n534 B.n533 585
R297 B.n531 B.n361 585
R298 B.n530 B.n529 585
R299 B.n528 B.n527 585
R300 B.n526 B.n525 585
R301 B.n524 B.n523 585
R302 B.n522 B.n521 585
R303 B.n520 B.n519 585
R304 B.n518 B.n517 585
R305 B.n516 B.n515 585
R306 B.n514 B.n513 585
R307 B.n512 B.n511 585
R308 B.n510 B.n509 585
R309 B.n508 B.n507 585
R310 B.n506 B.n505 585
R311 B.n504 B.n503 585
R312 B.n502 B.n501 585
R313 B.n500 B.n499 585
R314 B.n498 B.n497 585
R315 B.n496 B.n495 585
R316 B.n494 B.n493 585
R317 B.n492 B.n491 585
R318 B.n490 B.n489 585
R319 B.n488 B.n487 585
R320 B.n486 B.n485 585
R321 B.n484 B.n483 585
R322 B.n482 B.n481 585
R323 B.n480 B.n479 585
R324 B.n478 B.n477 585
R325 B.n476 B.n475 585
R326 B.n474 B.n473 585
R327 B.n472 B.n471 585
R328 B.n470 B.n469 585
R329 B.n468 B.n467 585
R330 B.n466 B.n465 585
R331 B.n464 B.n463 585
R332 B.n461 B.n460 585
R333 B.n459 B.n458 585
R334 B.n457 B.n456 585
R335 B.n455 B.n454 585
R336 B.n453 B.n452 585
R337 B.n451 B.n450 585
R338 B.n449 B.n448 585
R339 B.n447 B.n446 585
R340 B.n445 B.n444 585
R341 B.n443 B.n442 585
R342 B.n440 B.n439 585
R343 B.n438 B.n437 585
R344 B.n436 B.n435 585
R345 B.n434 B.n433 585
R346 B.n432 B.n431 585
R347 B.n430 B.n429 585
R348 B.n428 B.n427 585
R349 B.n426 B.n425 585
R350 B.n424 B.n423 585
R351 B.n422 B.n421 585
R352 B.n420 B.n419 585
R353 B.n418 B.n417 585
R354 B.n416 B.n415 585
R355 B.n414 B.n413 585
R356 B.n412 B.n411 585
R357 B.n410 B.n409 585
R358 B.n408 B.n407 585
R359 B.n406 B.n405 585
R360 B.n404 B.n403 585
R361 B.n402 B.n401 585
R362 B.n400 B.n399 585
R363 B.n398 B.n397 585
R364 B.n396 B.n395 585
R365 B.n394 B.n393 585
R366 B.n392 B.n391 585
R367 B.n390 B.n389 585
R368 B.n388 B.n387 585
R369 B.n386 B.n385 585
R370 B.n384 B.n383 585
R371 B.n382 B.n381 585
R372 B.n380 B.n379 585
R373 B.n378 B.n377 585
R374 B.n376 B.n375 585
R375 B.n374 B.n373 585
R376 B.n372 B.n371 585
R377 B.n370 B.n369 585
R378 B.n368 B.n367 585
R379 B.n366 B.n360 585
R380 B.n534 B.n360 585
R381 B.n538 B.n316 585
R382 B.n316 B.n315 585
R383 B.n540 B.n539 585
R384 B.n541 B.n540 585
R385 B.n310 B.n309 585
R386 B.n311 B.n310 585
R387 B.n549 B.n548 585
R388 B.n548 B.n547 585
R389 B.n550 B.n308 585
R390 B.n308 B.n307 585
R391 B.n552 B.n551 585
R392 B.n553 B.n552 585
R393 B.n302 B.n301 585
R394 B.n303 B.n302 585
R395 B.n561 B.n560 585
R396 B.n560 B.n559 585
R397 B.n562 B.n300 585
R398 B.n300 B.n299 585
R399 B.n564 B.n563 585
R400 B.n565 B.n564 585
R401 B.n294 B.n293 585
R402 B.n295 B.n294 585
R403 B.n574 B.n573 585
R404 B.n573 B.n572 585
R405 B.n575 B.n292 585
R406 B.n571 B.n292 585
R407 B.n577 B.n576 585
R408 B.n578 B.n577 585
R409 B.n287 B.n286 585
R410 B.n288 B.n287 585
R411 B.n587 B.n586 585
R412 B.n586 B.n585 585
R413 B.n588 B.n285 585
R414 B.n584 B.n285 585
R415 B.n590 B.n589 585
R416 B.n591 B.n590 585
R417 B.n280 B.n279 585
R418 B.n281 B.n280 585
R419 B.n600 B.n599 585
R420 B.n599 B.n598 585
R421 B.n601 B.n278 585
R422 B.n597 B.n278 585
R423 B.n603 B.n602 585
R424 B.n604 B.n603 585
R425 B.n273 B.n272 585
R426 B.n274 B.n273 585
R427 B.n613 B.n612 585
R428 B.n612 B.n611 585
R429 B.n614 B.n271 585
R430 B.n271 B.n270 585
R431 B.n616 B.n615 585
R432 B.n617 B.n616 585
R433 B.n3 B.n0 585
R434 B.n4 B.n3 585
R435 B.n716 B.n1 585
R436 B.n717 B.n716 585
R437 B.n715 B.n714 585
R438 B.n715 B.n8 585
R439 B.n713 B.n9 585
R440 B.n626 B.n9 585
R441 B.n712 B.n711 585
R442 B.n711 B.n710 585
R443 B.n11 B.n10 585
R444 B.n709 B.n11 585
R445 B.n707 B.n706 585
R446 B.n708 B.n707 585
R447 B.n705 B.n15 585
R448 B.n18 B.n15 585
R449 B.n704 B.n703 585
R450 B.n703 B.n702 585
R451 B.n17 B.n16 585
R452 B.n701 B.n17 585
R453 B.n699 B.n698 585
R454 B.n700 B.n699 585
R455 B.n697 B.n22 585
R456 B.n25 B.n22 585
R457 B.n696 B.n695 585
R458 B.n695 B.n694 585
R459 B.n24 B.n23 585
R460 B.n693 B.n24 585
R461 B.n691 B.n690 585
R462 B.n692 B.n691 585
R463 B.n689 B.n29 585
R464 B.n32 B.n29 585
R465 B.n688 B.n687 585
R466 B.n687 B.n686 585
R467 B.n31 B.n30 585
R468 B.n685 B.n31 585
R469 B.n683 B.n682 585
R470 B.n684 B.n683 585
R471 B.n681 B.n37 585
R472 B.n37 B.n36 585
R473 B.n680 B.n679 585
R474 B.n679 B.n678 585
R475 B.n39 B.n38 585
R476 B.n677 B.n39 585
R477 B.n675 B.n674 585
R478 B.n676 B.n675 585
R479 B.n673 B.n44 585
R480 B.n44 B.n43 585
R481 B.n672 B.n671 585
R482 B.n671 B.n670 585
R483 B.n46 B.n45 585
R484 B.n669 B.n46 585
R485 B.n667 B.n666 585
R486 B.n668 B.n667 585
R487 B.n665 B.n51 585
R488 B.n51 B.n50 585
R489 B.n720 B.n719 585
R490 B.n718 B.n2 585
R491 B.n663 B.n51 545.355
R492 B.n659 B.n96 545.355
R493 B.n360 B.n314 545.355
R494 B.n536 B.n316 545.355
R495 B.n100 B.t8 465.134
R496 B.n97 B.t16 465.134
R497 B.n364 B.t19 465.134
R498 B.n362 B.t12 465.134
R499 B.n661 B.n660 256.663
R500 B.n661 B.n94 256.663
R501 B.n661 B.n93 256.663
R502 B.n661 B.n92 256.663
R503 B.n661 B.n91 256.663
R504 B.n661 B.n90 256.663
R505 B.n661 B.n89 256.663
R506 B.n661 B.n88 256.663
R507 B.n661 B.n87 256.663
R508 B.n661 B.n86 256.663
R509 B.n661 B.n85 256.663
R510 B.n661 B.n84 256.663
R511 B.n661 B.n83 256.663
R512 B.n661 B.n82 256.663
R513 B.n661 B.n81 256.663
R514 B.n661 B.n80 256.663
R515 B.n661 B.n79 256.663
R516 B.n661 B.n78 256.663
R517 B.n661 B.n77 256.663
R518 B.n661 B.n76 256.663
R519 B.n661 B.n75 256.663
R520 B.n661 B.n74 256.663
R521 B.n661 B.n73 256.663
R522 B.n661 B.n72 256.663
R523 B.n661 B.n71 256.663
R524 B.n661 B.n70 256.663
R525 B.n661 B.n69 256.663
R526 B.n661 B.n68 256.663
R527 B.n661 B.n67 256.663
R528 B.n661 B.n66 256.663
R529 B.n661 B.n65 256.663
R530 B.n661 B.n64 256.663
R531 B.n661 B.n63 256.663
R532 B.n661 B.n62 256.663
R533 B.n661 B.n61 256.663
R534 B.n661 B.n60 256.663
R535 B.n661 B.n59 256.663
R536 B.n661 B.n58 256.663
R537 B.n661 B.n57 256.663
R538 B.n661 B.n56 256.663
R539 B.n661 B.n55 256.663
R540 B.n661 B.n54 256.663
R541 B.n662 B.n661 256.663
R542 B.n535 B.n534 256.663
R543 B.n534 B.n319 256.663
R544 B.n534 B.n320 256.663
R545 B.n534 B.n321 256.663
R546 B.n534 B.n322 256.663
R547 B.n534 B.n323 256.663
R548 B.n534 B.n324 256.663
R549 B.n534 B.n325 256.663
R550 B.n534 B.n326 256.663
R551 B.n534 B.n327 256.663
R552 B.n534 B.n328 256.663
R553 B.n534 B.n329 256.663
R554 B.n534 B.n330 256.663
R555 B.n534 B.n331 256.663
R556 B.n534 B.n332 256.663
R557 B.n534 B.n333 256.663
R558 B.n534 B.n334 256.663
R559 B.n534 B.n335 256.663
R560 B.n534 B.n336 256.663
R561 B.n534 B.n337 256.663
R562 B.n534 B.n338 256.663
R563 B.n534 B.n339 256.663
R564 B.n534 B.n340 256.663
R565 B.n534 B.n341 256.663
R566 B.n534 B.n342 256.663
R567 B.n534 B.n343 256.663
R568 B.n534 B.n344 256.663
R569 B.n534 B.n345 256.663
R570 B.n534 B.n346 256.663
R571 B.n534 B.n347 256.663
R572 B.n534 B.n348 256.663
R573 B.n534 B.n349 256.663
R574 B.n534 B.n350 256.663
R575 B.n534 B.n351 256.663
R576 B.n534 B.n352 256.663
R577 B.n534 B.n353 256.663
R578 B.n534 B.n354 256.663
R579 B.n534 B.n355 256.663
R580 B.n534 B.n356 256.663
R581 B.n534 B.n357 256.663
R582 B.n534 B.n358 256.663
R583 B.n534 B.n359 256.663
R584 B.n722 B.n721 256.663
R585 B.n103 B.n53 163.367
R586 B.n107 B.n106 163.367
R587 B.n111 B.n110 163.367
R588 B.n115 B.n114 163.367
R589 B.n119 B.n118 163.367
R590 B.n123 B.n122 163.367
R591 B.n127 B.n126 163.367
R592 B.n131 B.n130 163.367
R593 B.n135 B.n134 163.367
R594 B.n139 B.n138 163.367
R595 B.n143 B.n142 163.367
R596 B.n147 B.n146 163.367
R597 B.n151 B.n150 163.367
R598 B.n155 B.n154 163.367
R599 B.n159 B.n158 163.367
R600 B.n163 B.n162 163.367
R601 B.n167 B.n166 163.367
R602 B.n171 B.n170 163.367
R603 B.n175 B.n174 163.367
R604 B.n179 B.n178 163.367
R605 B.n183 B.n182 163.367
R606 B.n187 B.n186 163.367
R607 B.n191 B.n190 163.367
R608 B.n195 B.n194 163.367
R609 B.n199 B.n198 163.367
R610 B.n203 B.n202 163.367
R611 B.n207 B.n206 163.367
R612 B.n211 B.n210 163.367
R613 B.n215 B.n214 163.367
R614 B.n219 B.n218 163.367
R615 B.n223 B.n222 163.367
R616 B.n227 B.n226 163.367
R617 B.n231 B.n230 163.367
R618 B.n235 B.n234 163.367
R619 B.n239 B.n238 163.367
R620 B.n243 B.n242 163.367
R621 B.n247 B.n246 163.367
R622 B.n251 B.n250 163.367
R623 B.n255 B.n254 163.367
R624 B.n259 B.n258 163.367
R625 B.n263 B.n262 163.367
R626 B.n265 B.n95 163.367
R627 B.n542 B.n314 163.367
R628 B.n542 B.n312 163.367
R629 B.n546 B.n312 163.367
R630 B.n546 B.n306 163.367
R631 B.n554 B.n306 163.367
R632 B.n554 B.n304 163.367
R633 B.n558 B.n304 163.367
R634 B.n558 B.n298 163.367
R635 B.n566 B.n298 163.367
R636 B.n566 B.n296 163.367
R637 B.n570 B.n296 163.367
R638 B.n570 B.n291 163.367
R639 B.n579 B.n291 163.367
R640 B.n579 B.n289 163.367
R641 B.n583 B.n289 163.367
R642 B.n583 B.n284 163.367
R643 B.n592 B.n284 163.367
R644 B.n592 B.n282 163.367
R645 B.n596 B.n282 163.367
R646 B.n596 B.n277 163.367
R647 B.n605 B.n277 163.367
R648 B.n605 B.n275 163.367
R649 B.n610 B.n275 163.367
R650 B.n610 B.n269 163.367
R651 B.n618 B.n269 163.367
R652 B.n619 B.n618 163.367
R653 B.n619 B.n5 163.367
R654 B.n6 B.n5 163.367
R655 B.n7 B.n6 163.367
R656 B.n625 B.n7 163.367
R657 B.n627 B.n625 163.367
R658 B.n627 B.n12 163.367
R659 B.n13 B.n12 163.367
R660 B.n14 B.n13 163.367
R661 B.n632 B.n14 163.367
R662 B.n632 B.n19 163.367
R663 B.n20 B.n19 163.367
R664 B.n21 B.n20 163.367
R665 B.n637 B.n21 163.367
R666 B.n637 B.n26 163.367
R667 B.n27 B.n26 163.367
R668 B.n28 B.n27 163.367
R669 B.n642 B.n28 163.367
R670 B.n642 B.n33 163.367
R671 B.n34 B.n33 163.367
R672 B.n35 B.n34 163.367
R673 B.n647 B.n35 163.367
R674 B.n647 B.n40 163.367
R675 B.n41 B.n40 163.367
R676 B.n42 B.n41 163.367
R677 B.n652 B.n42 163.367
R678 B.n652 B.n47 163.367
R679 B.n48 B.n47 163.367
R680 B.n49 B.n48 163.367
R681 B.n96 B.n49 163.367
R682 B.n533 B.n318 163.367
R683 B.n533 B.n361 163.367
R684 B.n529 B.n528 163.367
R685 B.n525 B.n524 163.367
R686 B.n521 B.n520 163.367
R687 B.n517 B.n516 163.367
R688 B.n513 B.n512 163.367
R689 B.n509 B.n508 163.367
R690 B.n505 B.n504 163.367
R691 B.n501 B.n500 163.367
R692 B.n497 B.n496 163.367
R693 B.n493 B.n492 163.367
R694 B.n489 B.n488 163.367
R695 B.n485 B.n484 163.367
R696 B.n481 B.n480 163.367
R697 B.n477 B.n476 163.367
R698 B.n473 B.n472 163.367
R699 B.n469 B.n468 163.367
R700 B.n465 B.n464 163.367
R701 B.n460 B.n459 163.367
R702 B.n456 B.n455 163.367
R703 B.n452 B.n451 163.367
R704 B.n448 B.n447 163.367
R705 B.n444 B.n443 163.367
R706 B.n439 B.n438 163.367
R707 B.n435 B.n434 163.367
R708 B.n431 B.n430 163.367
R709 B.n427 B.n426 163.367
R710 B.n423 B.n422 163.367
R711 B.n419 B.n418 163.367
R712 B.n415 B.n414 163.367
R713 B.n411 B.n410 163.367
R714 B.n407 B.n406 163.367
R715 B.n403 B.n402 163.367
R716 B.n399 B.n398 163.367
R717 B.n395 B.n394 163.367
R718 B.n391 B.n390 163.367
R719 B.n387 B.n386 163.367
R720 B.n383 B.n382 163.367
R721 B.n379 B.n378 163.367
R722 B.n375 B.n374 163.367
R723 B.n371 B.n370 163.367
R724 B.n367 B.n360 163.367
R725 B.n540 B.n316 163.367
R726 B.n540 B.n310 163.367
R727 B.n548 B.n310 163.367
R728 B.n548 B.n308 163.367
R729 B.n552 B.n308 163.367
R730 B.n552 B.n302 163.367
R731 B.n560 B.n302 163.367
R732 B.n560 B.n300 163.367
R733 B.n564 B.n300 163.367
R734 B.n564 B.n294 163.367
R735 B.n573 B.n294 163.367
R736 B.n573 B.n292 163.367
R737 B.n577 B.n292 163.367
R738 B.n577 B.n287 163.367
R739 B.n586 B.n287 163.367
R740 B.n586 B.n285 163.367
R741 B.n590 B.n285 163.367
R742 B.n590 B.n280 163.367
R743 B.n599 B.n280 163.367
R744 B.n599 B.n278 163.367
R745 B.n603 B.n278 163.367
R746 B.n603 B.n273 163.367
R747 B.n612 B.n273 163.367
R748 B.n612 B.n271 163.367
R749 B.n616 B.n271 163.367
R750 B.n616 B.n3 163.367
R751 B.n720 B.n3 163.367
R752 B.n716 B.n2 163.367
R753 B.n716 B.n715 163.367
R754 B.n715 B.n9 163.367
R755 B.n711 B.n9 163.367
R756 B.n711 B.n11 163.367
R757 B.n707 B.n11 163.367
R758 B.n707 B.n15 163.367
R759 B.n703 B.n15 163.367
R760 B.n703 B.n17 163.367
R761 B.n699 B.n17 163.367
R762 B.n699 B.n22 163.367
R763 B.n695 B.n22 163.367
R764 B.n695 B.n24 163.367
R765 B.n691 B.n24 163.367
R766 B.n691 B.n29 163.367
R767 B.n687 B.n29 163.367
R768 B.n687 B.n31 163.367
R769 B.n683 B.n31 163.367
R770 B.n683 B.n37 163.367
R771 B.n679 B.n37 163.367
R772 B.n679 B.n39 163.367
R773 B.n675 B.n39 163.367
R774 B.n675 B.n44 163.367
R775 B.n671 B.n44 163.367
R776 B.n671 B.n46 163.367
R777 B.n667 B.n46 163.367
R778 B.n667 B.n51 163.367
R779 B.n97 B.t17 93.7522
R780 B.n364 B.t21 93.7522
R781 B.n100 B.t10 93.7385
R782 B.n362 B.t15 93.7385
R783 B.n534 B.n315 91.9225
R784 B.n661 B.n50 91.9225
R785 B.n663 B.n662 71.676
R786 B.n103 B.n54 71.676
R787 B.n107 B.n55 71.676
R788 B.n111 B.n56 71.676
R789 B.n115 B.n57 71.676
R790 B.n119 B.n58 71.676
R791 B.n123 B.n59 71.676
R792 B.n127 B.n60 71.676
R793 B.n131 B.n61 71.676
R794 B.n135 B.n62 71.676
R795 B.n139 B.n63 71.676
R796 B.n143 B.n64 71.676
R797 B.n147 B.n65 71.676
R798 B.n151 B.n66 71.676
R799 B.n155 B.n67 71.676
R800 B.n159 B.n68 71.676
R801 B.n163 B.n69 71.676
R802 B.n167 B.n70 71.676
R803 B.n171 B.n71 71.676
R804 B.n175 B.n72 71.676
R805 B.n179 B.n73 71.676
R806 B.n183 B.n74 71.676
R807 B.n187 B.n75 71.676
R808 B.n191 B.n76 71.676
R809 B.n195 B.n77 71.676
R810 B.n199 B.n78 71.676
R811 B.n203 B.n79 71.676
R812 B.n207 B.n80 71.676
R813 B.n211 B.n81 71.676
R814 B.n215 B.n82 71.676
R815 B.n219 B.n83 71.676
R816 B.n223 B.n84 71.676
R817 B.n227 B.n85 71.676
R818 B.n231 B.n86 71.676
R819 B.n235 B.n87 71.676
R820 B.n239 B.n88 71.676
R821 B.n243 B.n89 71.676
R822 B.n247 B.n90 71.676
R823 B.n251 B.n91 71.676
R824 B.n255 B.n92 71.676
R825 B.n259 B.n93 71.676
R826 B.n263 B.n94 71.676
R827 B.n660 B.n95 71.676
R828 B.n660 B.n659 71.676
R829 B.n265 B.n94 71.676
R830 B.n262 B.n93 71.676
R831 B.n258 B.n92 71.676
R832 B.n254 B.n91 71.676
R833 B.n250 B.n90 71.676
R834 B.n246 B.n89 71.676
R835 B.n242 B.n88 71.676
R836 B.n238 B.n87 71.676
R837 B.n234 B.n86 71.676
R838 B.n230 B.n85 71.676
R839 B.n226 B.n84 71.676
R840 B.n222 B.n83 71.676
R841 B.n218 B.n82 71.676
R842 B.n214 B.n81 71.676
R843 B.n210 B.n80 71.676
R844 B.n206 B.n79 71.676
R845 B.n202 B.n78 71.676
R846 B.n198 B.n77 71.676
R847 B.n194 B.n76 71.676
R848 B.n190 B.n75 71.676
R849 B.n186 B.n74 71.676
R850 B.n182 B.n73 71.676
R851 B.n178 B.n72 71.676
R852 B.n174 B.n71 71.676
R853 B.n170 B.n70 71.676
R854 B.n166 B.n69 71.676
R855 B.n162 B.n68 71.676
R856 B.n158 B.n67 71.676
R857 B.n154 B.n66 71.676
R858 B.n150 B.n65 71.676
R859 B.n146 B.n64 71.676
R860 B.n142 B.n63 71.676
R861 B.n138 B.n62 71.676
R862 B.n134 B.n61 71.676
R863 B.n130 B.n60 71.676
R864 B.n126 B.n59 71.676
R865 B.n122 B.n58 71.676
R866 B.n118 B.n57 71.676
R867 B.n114 B.n56 71.676
R868 B.n110 B.n55 71.676
R869 B.n106 B.n54 71.676
R870 B.n662 B.n53 71.676
R871 B.n536 B.n535 71.676
R872 B.n361 B.n319 71.676
R873 B.n528 B.n320 71.676
R874 B.n524 B.n321 71.676
R875 B.n520 B.n322 71.676
R876 B.n516 B.n323 71.676
R877 B.n512 B.n324 71.676
R878 B.n508 B.n325 71.676
R879 B.n504 B.n326 71.676
R880 B.n500 B.n327 71.676
R881 B.n496 B.n328 71.676
R882 B.n492 B.n329 71.676
R883 B.n488 B.n330 71.676
R884 B.n484 B.n331 71.676
R885 B.n480 B.n332 71.676
R886 B.n476 B.n333 71.676
R887 B.n472 B.n334 71.676
R888 B.n468 B.n335 71.676
R889 B.n464 B.n336 71.676
R890 B.n459 B.n337 71.676
R891 B.n455 B.n338 71.676
R892 B.n451 B.n339 71.676
R893 B.n447 B.n340 71.676
R894 B.n443 B.n341 71.676
R895 B.n438 B.n342 71.676
R896 B.n434 B.n343 71.676
R897 B.n430 B.n344 71.676
R898 B.n426 B.n345 71.676
R899 B.n422 B.n346 71.676
R900 B.n418 B.n347 71.676
R901 B.n414 B.n348 71.676
R902 B.n410 B.n349 71.676
R903 B.n406 B.n350 71.676
R904 B.n402 B.n351 71.676
R905 B.n398 B.n352 71.676
R906 B.n394 B.n353 71.676
R907 B.n390 B.n354 71.676
R908 B.n386 B.n355 71.676
R909 B.n382 B.n356 71.676
R910 B.n378 B.n357 71.676
R911 B.n374 B.n358 71.676
R912 B.n370 B.n359 71.676
R913 B.n535 B.n318 71.676
R914 B.n529 B.n319 71.676
R915 B.n525 B.n320 71.676
R916 B.n521 B.n321 71.676
R917 B.n517 B.n322 71.676
R918 B.n513 B.n323 71.676
R919 B.n509 B.n324 71.676
R920 B.n505 B.n325 71.676
R921 B.n501 B.n326 71.676
R922 B.n497 B.n327 71.676
R923 B.n493 B.n328 71.676
R924 B.n489 B.n329 71.676
R925 B.n485 B.n330 71.676
R926 B.n481 B.n331 71.676
R927 B.n477 B.n332 71.676
R928 B.n473 B.n333 71.676
R929 B.n469 B.n334 71.676
R930 B.n465 B.n335 71.676
R931 B.n460 B.n336 71.676
R932 B.n456 B.n337 71.676
R933 B.n452 B.n338 71.676
R934 B.n448 B.n339 71.676
R935 B.n444 B.n340 71.676
R936 B.n439 B.n341 71.676
R937 B.n435 B.n342 71.676
R938 B.n431 B.n343 71.676
R939 B.n427 B.n344 71.676
R940 B.n423 B.n345 71.676
R941 B.n419 B.n346 71.676
R942 B.n415 B.n347 71.676
R943 B.n411 B.n348 71.676
R944 B.n407 B.n349 71.676
R945 B.n403 B.n350 71.676
R946 B.n399 B.n351 71.676
R947 B.n395 B.n352 71.676
R948 B.n391 B.n353 71.676
R949 B.n387 B.n354 71.676
R950 B.n383 B.n355 71.676
R951 B.n379 B.n356 71.676
R952 B.n375 B.n357 71.676
R953 B.n371 B.n358 71.676
R954 B.n367 B.n359 71.676
R955 B.n721 B.n720 71.676
R956 B.n721 B.n2 71.676
R957 B.n98 B.t18 67.9582
R958 B.n365 B.t20 67.9582
R959 B.n101 B.t11 67.9445
R960 B.n363 B.t14 67.9445
R961 B.n102 B.n101 59.5399
R962 B.n99 B.n98 59.5399
R963 B.n441 B.n365 59.5399
R964 B.n462 B.n363 59.5399
R965 B.n541 B.n315 46.302
R966 B.n541 B.n311 46.302
R967 B.n547 B.n311 46.302
R968 B.n547 B.n307 46.302
R969 B.n553 B.n307 46.302
R970 B.n559 B.n303 46.302
R971 B.n559 B.n299 46.302
R972 B.n565 B.n299 46.302
R973 B.n565 B.n295 46.302
R974 B.n572 B.n295 46.302
R975 B.n572 B.n571 46.302
R976 B.n578 B.n288 46.302
R977 B.n585 B.n288 46.302
R978 B.n585 B.n584 46.302
R979 B.n591 B.n281 46.302
R980 B.n598 B.n281 46.302
R981 B.n598 B.n597 46.302
R982 B.n604 B.n274 46.302
R983 B.n611 B.n274 46.302
R984 B.n617 B.n270 46.302
R985 B.n617 B.n4 46.302
R986 B.n719 B.n4 46.302
R987 B.n719 B.n718 46.302
R988 B.n718 B.n717 46.302
R989 B.n717 B.n8 46.302
R990 B.n626 B.n8 46.302
R991 B.n710 B.n709 46.302
R992 B.n709 B.n708 46.302
R993 B.n702 B.n18 46.302
R994 B.n702 B.n701 46.302
R995 B.n701 B.n700 46.302
R996 B.n694 B.n25 46.302
R997 B.n694 B.n693 46.302
R998 B.n693 B.n692 46.302
R999 B.n686 B.n32 46.302
R1000 B.n686 B.n685 46.302
R1001 B.n685 B.n684 46.302
R1002 B.n684 B.n36 46.302
R1003 B.n678 B.n36 46.302
R1004 B.n678 B.n677 46.302
R1005 B.n676 B.n43 46.302
R1006 B.n670 B.n43 46.302
R1007 B.n670 B.n669 46.302
R1008 B.n669 B.n668 46.302
R1009 B.n668 B.n50 46.302
R1010 B.n604 B.t4 44.9401
R1011 B.n708 B.t3 44.9401
R1012 B.n611 B.t6 43.5783
R1013 B.n710 B.t5 43.5783
R1014 B.t13 B.n303 42.2165
R1015 B.n677 B.t9 42.2165
R1016 B.n591 B.t2 40.8547
R1017 B.n700 B.t7 40.8547
R1018 B.n578 B.t0 36.7693
R1019 B.n692 B.t1 36.7693
R1020 B.n658 B.n657 35.4346
R1021 B.n538 B.n537 35.4346
R1022 B.n366 B.n313 35.4346
R1023 B.n665 B.n664 35.4346
R1024 B.n101 B.n100 25.7944
R1025 B.n98 B.n97 25.7944
R1026 B.n365 B.n364 25.7944
R1027 B.n363 B.n362 25.7944
R1028 B B.n722 18.0485
R1029 B.n539 B.n538 10.6151
R1030 B.n539 B.n309 10.6151
R1031 B.n549 B.n309 10.6151
R1032 B.n550 B.n549 10.6151
R1033 B.n551 B.n550 10.6151
R1034 B.n551 B.n301 10.6151
R1035 B.n561 B.n301 10.6151
R1036 B.n562 B.n561 10.6151
R1037 B.n563 B.n562 10.6151
R1038 B.n563 B.n293 10.6151
R1039 B.n574 B.n293 10.6151
R1040 B.n575 B.n574 10.6151
R1041 B.n576 B.n575 10.6151
R1042 B.n576 B.n286 10.6151
R1043 B.n587 B.n286 10.6151
R1044 B.n588 B.n587 10.6151
R1045 B.n589 B.n588 10.6151
R1046 B.n589 B.n279 10.6151
R1047 B.n600 B.n279 10.6151
R1048 B.n601 B.n600 10.6151
R1049 B.n602 B.n601 10.6151
R1050 B.n602 B.n272 10.6151
R1051 B.n613 B.n272 10.6151
R1052 B.n614 B.n613 10.6151
R1053 B.n615 B.n614 10.6151
R1054 B.n615 B.n0 10.6151
R1055 B.n537 B.n317 10.6151
R1056 B.n532 B.n317 10.6151
R1057 B.n532 B.n531 10.6151
R1058 B.n531 B.n530 10.6151
R1059 B.n530 B.n527 10.6151
R1060 B.n527 B.n526 10.6151
R1061 B.n526 B.n523 10.6151
R1062 B.n523 B.n522 10.6151
R1063 B.n522 B.n519 10.6151
R1064 B.n519 B.n518 10.6151
R1065 B.n518 B.n515 10.6151
R1066 B.n515 B.n514 10.6151
R1067 B.n514 B.n511 10.6151
R1068 B.n511 B.n510 10.6151
R1069 B.n510 B.n507 10.6151
R1070 B.n507 B.n506 10.6151
R1071 B.n506 B.n503 10.6151
R1072 B.n503 B.n502 10.6151
R1073 B.n502 B.n499 10.6151
R1074 B.n499 B.n498 10.6151
R1075 B.n498 B.n495 10.6151
R1076 B.n495 B.n494 10.6151
R1077 B.n494 B.n491 10.6151
R1078 B.n491 B.n490 10.6151
R1079 B.n490 B.n487 10.6151
R1080 B.n487 B.n486 10.6151
R1081 B.n486 B.n483 10.6151
R1082 B.n483 B.n482 10.6151
R1083 B.n482 B.n479 10.6151
R1084 B.n479 B.n478 10.6151
R1085 B.n478 B.n475 10.6151
R1086 B.n475 B.n474 10.6151
R1087 B.n474 B.n471 10.6151
R1088 B.n471 B.n470 10.6151
R1089 B.n470 B.n467 10.6151
R1090 B.n467 B.n466 10.6151
R1091 B.n466 B.n463 10.6151
R1092 B.n461 B.n458 10.6151
R1093 B.n458 B.n457 10.6151
R1094 B.n457 B.n454 10.6151
R1095 B.n454 B.n453 10.6151
R1096 B.n453 B.n450 10.6151
R1097 B.n450 B.n449 10.6151
R1098 B.n449 B.n446 10.6151
R1099 B.n446 B.n445 10.6151
R1100 B.n445 B.n442 10.6151
R1101 B.n440 B.n437 10.6151
R1102 B.n437 B.n436 10.6151
R1103 B.n436 B.n433 10.6151
R1104 B.n433 B.n432 10.6151
R1105 B.n432 B.n429 10.6151
R1106 B.n429 B.n428 10.6151
R1107 B.n428 B.n425 10.6151
R1108 B.n425 B.n424 10.6151
R1109 B.n424 B.n421 10.6151
R1110 B.n421 B.n420 10.6151
R1111 B.n420 B.n417 10.6151
R1112 B.n417 B.n416 10.6151
R1113 B.n416 B.n413 10.6151
R1114 B.n413 B.n412 10.6151
R1115 B.n412 B.n409 10.6151
R1116 B.n409 B.n408 10.6151
R1117 B.n408 B.n405 10.6151
R1118 B.n405 B.n404 10.6151
R1119 B.n404 B.n401 10.6151
R1120 B.n401 B.n400 10.6151
R1121 B.n400 B.n397 10.6151
R1122 B.n397 B.n396 10.6151
R1123 B.n396 B.n393 10.6151
R1124 B.n393 B.n392 10.6151
R1125 B.n392 B.n389 10.6151
R1126 B.n389 B.n388 10.6151
R1127 B.n388 B.n385 10.6151
R1128 B.n385 B.n384 10.6151
R1129 B.n384 B.n381 10.6151
R1130 B.n381 B.n380 10.6151
R1131 B.n380 B.n377 10.6151
R1132 B.n377 B.n376 10.6151
R1133 B.n376 B.n373 10.6151
R1134 B.n373 B.n372 10.6151
R1135 B.n372 B.n369 10.6151
R1136 B.n369 B.n368 10.6151
R1137 B.n368 B.n366 10.6151
R1138 B.n543 B.n313 10.6151
R1139 B.n544 B.n543 10.6151
R1140 B.n545 B.n544 10.6151
R1141 B.n545 B.n305 10.6151
R1142 B.n555 B.n305 10.6151
R1143 B.n556 B.n555 10.6151
R1144 B.n557 B.n556 10.6151
R1145 B.n557 B.n297 10.6151
R1146 B.n567 B.n297 10.6151
R1147 B.n568 B.n567 10.6151
R1148 B.n569 B.n568 10.6151
R1149 B.n569 B.n290 10.6151
R1150 B.n580 B.n290 10.6151
R1151 B.n581 B.n580 10.6151
R1152 B.n582 B.n581 10.6151
R1153 B.n582 B.n283 10.6151
R1154 B.n593 B.n283 10.6151
R1155 B.n594 B.n593 10.6151
R1156 B.n595 B.n594 10.6151
R1157 B.n595 B.n276 10.6151
R1158 B.n606 B.n276 10.6151
R1159 B.n607 B.n606 10.6151
R1160 B.n609 B.n607 10.6151
R1161 B.n609 B.n608 10.6151
R1162 B.n608 B.n268 10.6151
R1163 B.n620 B.n268 10.6151
R1164 B.n621 B.n620 10.6151
R1165 B.n622 B.n621 10.6151
R1166 B.n623 B.n622 10.6151
R1167 B.n624 B.n623 10.6151
R1168 B.n628 B.n624 10.6151
R1169 B.n629 B.n628 10.6151
R1170 B.n630 B.n629 10.6151
R1171 B.n631 B.n630 10.6151
R1172 B.n633 B.n631 10.6151
R1173 B.n634 B.n633 10.6151
R1174 B.n635 B.n634 10.6151
R1175 B.n636 B.n635 10.6151
R1176 B.n638 B.n636 10.6151
R1177 B.n639 B.n638 10.6151
R1178 B.n640 B.n639 10.6151
R1179 B.n641 B.n640 10.6151
R1180 B.n643 B.n641 10.6151
R1181 B.n644 B.n643 10.6151
R1182 B.n645 B.n644 10.6151
R1183 B.n646 B.n645 10.6151
R1184 B.n648 B.n646 10.6151
R1185 B.n649 B.n648 10.6151
R1186 B.n650 B.n649 10.6151
R1187 B.n651 B.n650 10.6151
R1188 B.n653 B.n651 10.6151
R1189 B.n654 B.n653 10.6151
R1190 B.n655 B.n654 10.6151
R1191 B.n656 B.n655 10.6151
R1192 B.n657 B.n656 10.6151
R1193 B.n714 B.n1 10.6151
R1194 B.n714 B.n713 10.6151
R1195 B.n713 B.n712 10.6151
R1196 B.n712 B.n10 10.6151
R1197 B.n706 B.n10 10.6151
R1198 B.n706 B.n705 10.6151
R1199 B.n705 B.n704 10.6151
R1200 B.n704 B.n16 10.6151
R1201 B.n698 B.n16 10.6151
R1202 B.n698 B.n697 10.6151
R1203 B.n697 B.n696 10.6151
R1204 B.n696 B.n23 10.6151
R1205 B.n690 B.n23 10.6151
R1206 B.n690 B.n689 10.6151
R1207 B.n689 B.n688 10.6151
R1208 B.n688 B.n30 10.6151
R1209 B.n682 B.n30 10.6151
R1210 B.n682 B.n681 10.6151
R1211 B.n681 B.n680 10.6151
R1212 B.n680 B.n38 10.6151
R1213 B.n674 B.n38 10.6151
R1214 B.n674 B.n673 10.6151
R1215 B.n673 B.n672 10.6151
R1216 B.n672 B.n45 10.6151
R1217 B.n666 B.n45 10.6151
R1218 B.n666 B.n665 10.6151
R1219 B.n664 B.n52 10.6151
R1220 B.n104 B.n52 10.6151
R1221 B.n105 B.n104 10.6151
R1222 B.n108 B.n105 10.6151
R1223 B.n109 B.n108 10.6151
R1224 B.n112 B.n109 10.6151
R1225 B.n113 B.n112 10.6151
R1226 B.n116 B.n113 10.6151
R1227 B.n117 B.n116 10.6151
R1228 B.n120 B.n117 10.6151
R1229 B.n121 B.n120 10.6151
R1230 B.n124 B.n121 10.6151
R1231 B.n125 B.n124 10.6151
R1232 B.n128 B.n125 10.6151
R1233 B.n129 B.n128 10.6151
R1234 B.n132 B.n129 10.6151
R1235 B.n133 B.n132 10.6151
R1236 B.n136 B.n133 10.6151
R1237 B.n137 B.n136 10.6151
R1238 B.n140 B.n137 10.6151
R1239 B.n141 B.n140 10.6151
R1240 B.n144 B.n141 10.6151
R1241 B.n145 B.n144 10.6151
R1242 B.n148 B.n145 10.6151
R1243 B.n149 B.n148 10.6151
R1244 B.n152 B.n149 10.6151
R1245 B.n153 B.n152 10.6151
R1246 B.n156 B.n153 10.6151
R1247 B.n157 B.n156 10.6151
R1248 B.n160 B.n157 10.6151
R1249 B.n161 B.n160 10.6151
R1250 B.n164 B.n161 10.6151
R1251 B.n165 B.n164 10.6151
R1252 B.n168 B.n165 10.6151
R1253 B.n169 B.n168 10.6151
R1254 B.n172 B.n169 10.6151
R1255 B.n173 B.n172 10.6151
R1256 B.n177 B.n176 10.6151
R1257 B.n180 B.n177 10.6151
R1258 B.n181 B.n180 10.6151
R1259 B.n184 B.n181 10.6151
R1260 B.n185 B.n184 10.6151
R1261 B.n188 B.n185 10.6151
R1262 B.n189 B.n188 10.6151
R1263 B.n192 B.n189 10.6151
R1264 B.n193 B.n192 10.6151
R1265 B.n197 B.n196 10.6151
R1266 B.n200 B.n197 10.6151
R1267 B.n201 B.n200 10.6151
R1268 B.n204 B.n201 10.6151
R1269 B.n205 B.n204 10.6151
R1270 B.n208 B.n205 10.6151
R1271 B.n209 B.n208 10.6151
R1272 B.n212 B.n209 10.6151
R1273 B.n213 B.n212 10.6151
R1274 B.n216 B.n213 10.6151
R1275 B.n217 B.n216 10.6151
R1276 B.n220 B.n217 10.6151
R1277 B.n221 B.n220 10.6151
R1278 B.n224 B.n221 10.6151
R1279 B.n225 B.n224 10.6151
R1280 B.n228 B.n225 10.6151
R1281 B.n229 B.n228 10.6151
R1282 B.n232 B.n229 10.6151
R1283 B.n233 B.n232 10.6151
R1284 B.n236 B.n233 10.6151
R1285 B.n237 B.n236 10.6151
R1286 B.n240 B.n237 10.6151
R1287 B.n241 B.n240 10.6151
R1288 B.n244 B.n241 10.6151
R1289 B.n245 B.n244 10.6151
R1290 B.n248 B.n245 10.6151
R1291 B.n249 B.n248 10.6151
R1292 B.n252 B.n249 10.6151
R1293 B.n253 B.n252 10.6151
R1294 B.n256 B.n253 10.6151
R1295 B.n257 B.n256 10.6151
R1296 B.n260 B.n257 10.6151
R1297 B.n261 B.n260 10.6151
R1298 B.n264 B.n261 10.6151
R1299 B.n266 B.n264 10.6151
R1300 B.n267 B.n266 10.6151
R1301 B.n658 B.n267 10.6151
R1302 B.n571 B.t0 9.53315
R1303 B.n32 B.t1 9.53315
R1304 B.n463 B.n462 9.36635
R1305 B.n441 B.n440 9.36635
R1306 B.n173 B.n102 9.36635
R1307 B.n196 B.n99 9.36635
R1308 B.n722 B.n0 8.11757
R1309 B.n722 B.n1 8.11757
R1310 B.n584 B.t2 5.44773
R1311 B.n25 B.t7 5.44773
R1312 B.n553 B.t13 4.08592
R1313 B.t9 B.n676 4.08592
R1314 B.t6 B.n270 2.72411
R1315 B.n626 B.t5 2.72411
R1316 B.n597 B.t4 1.36231
R1317 B.n18 B.t3 1.36231
R1318 B.n462 B.n461 1.24928
R1319 B.n442 B.n441 1.24928
R1320 B.n176 B.n102 1.24928
R1321 B.n193 B.n99 1.24928
R1322 VN.n2 VN.t5 317.216
R1323 VN.n15 VN.t1 317.216
R1324 VN.n11 VN.t7 301.974
R1325 VN.n24 VN.t6 301.974
R1326 VN.n3 VN.t3 262.209
R1327 VN.n9 VN.t0 262.209
R1328 VN.n16 VN.t4 262.209
R1329 VN.n22 VN.t2 262.209
R1330 VN.n23 VN.n13 161.3
R1331 VN.n21 VN.n20 161.3
R1332 VN.n19 VN.n14 161.3
R1333 VN.n18 VN.n17 161.3
R1334 VN.n10 VN.n0 161.3
R1335 VN.n8 VN.n7 161.3
R1336 VN.n6 VN.n1 161.3
R1337 VN.n5 VN.n4 161.3
R1338 VN.n25 VN.n24 80.6037
R1339 VN.n12 VN.n11 80.6037
R1340 VN.n11 VN.n10 56.2338
R1341 VN.n24 VN.n23 56.2338
R1342 VN.n3 VN.n2 46.7059
R1343 VN.n16 VN.n15 46.7059
R1344 VN.n18 VN.n15 43.9111
R1345 VN.n5 VN.n2 43.9111
R1346 VN VN.n25 43.0597
R1347 VN.n4 VN.n1 40.4106
R1348 VN.n8 VN.n1 40.4106
R1349 VN.n17 VN.n14 40.4106
R1350 VN.n21 VN.n14 40.4106
R1351 VN.n10 VN.n9 16.3106
R1352 VN.n23 VN.n22 16.3106
R1353 VN.n4 VN.n3 8.03383
R1354 VN.n9 VN.n8 8.03383
R1355 VN.n17 VN.n16 8.03383
R1356 VN.n22 VN.n21 8.03383
R1357 VN.n25 VN.n13 0.285035
R1358 VN.n12 VN.n0 0.285035
R1359 VN.n20 VN.n13 0.189894
R1360 VN.n20 VN.n19 0.189894
R1361 VN.n19 VN.n18 0.189894
R1362 VN.n6 VN.n5 0.189894
R1363 VN.n7 VN.n6 0.189894
R1364 VN.n7 VN.n0 0.189894
R1365 VN VN.n12 0.146778
R1366 VDD2.n2 VDD2.n1 65.8408
R1367 VDD2.n2 VDD2.n0 65.8408
R1368 VDD2 VDD2.n5 65.8379
R1369 VDD2.n4 VDD2.n3 65.3239
R1370 VDD2.n4 VDD2.n2 38.2541
R1371 VDD2.n5 VDD2.t3 1.82035
R1372 VDD2.n5 VDD2.t6 1.82035
R1373 VDD2.n3 VDD2.t1 1.82035
R1374 VDD2.n3 VDD2.t5 1.82035
R1375 VDD2.n1 VDD2.t7 1.82035
R1376 VDD2.n1 VDD2.t0 1.82035
R1377 VDD2.n0 VDD2.t2 1.82035
R1378 VDD2.n0 VDD2.t4 1.82035
R1379 VDD2 VDD2.n4 0.631965
C0 VDD2 VN 5.93693f
C1 VN VTAIL 5.86836f
C2 VDD2 VTAIL 8.94627f
C3 VP VN 5.49999f
C4 VN VDD1 0.148556f
C5 VDD2 VP 0.349134f
C6 VDD2 VDD1 0.976203f
C7 VP VTAIL 5.88247f
C8 VDD1 VTAIL 8.902579f
C9 VP VDD1 6.136919f
C10 VDD2 B 3.68095f
C11 VDD1 B 3.948351f
C12 VTAIL B 8.579203f
C13 VN B 9.50027f
C14 VP B 7.749012f
C15 VDD2.t2 B 0.22144f
C16 VDD2.t4 B 0.22144f
C17 VDD2.n0 B 1.97491f
C18 VDD2.t7 B 0.22144f
C19 VDD2.t0 B 0.22144f
C20 VDD2.n1 B 1.97491f
C21 VDD2.n2 B 2.32486f
C22 VDD2.t1 B 0.22144f
C23 VDD2.t5 B 0.22144f
C24 VDD2.n3 B 1.97215f
C25 VDD2.n4 B 2.36564f
C26 VDD2.t3 B 0.22144f
C27 VDD2.t6 B 0.22144f
C28 VDD2.n5 B 1.97487f
C29 VN.n0 B 0.050899f
C30 VN.t0 B 1.12742f
C31 VN.n1 B 0.030867f
C32 VN.t5 B 1.2094f
C33 VN.n2 B 0.478375f
C34 VN.t3 B 1.12742f
C35 VN.n3 B 0.457323f
C36 VN.n4 B 0.052581f
C37 VN.n5 B 0.163295f
C38 VN.n6 B 0.038144f
C39 VN.n7 B 0.038144f
C40 VN.n8 B 0.052581f
C41 VN.n9 B 0.422961f
C42 VN.n10 B 0.052802f
C43 VN.t7 B 1.18621f
C44 VN.n11 B 0.482318f
C45 VN.n12 B 0.035724f
C46 VN.n13 B 0.050899f
C47 VN.t2 B 1.12742f
C48 VN.n14 B 0.030867f
C49 VN.t1 B 1.2094f
C50 VN.n15 B 0.478375f
C51 VN.t4 B 1.12742f
C52 VN.n16 B 0.457323f
C53 VN.n17 B 0.052581f
C54 VN.n18 B 0.163295f
C55 VN.n19 B 0.038144f
C56 VN.n20 B 0.038144f
C57 VN.n21 B 0.052581f
C58 VN.n22 B 0.422961f
C59 VN.n23 B 0.052802f
C60 VN.t6 B 1.18621f
C61 VN.n24 B 0.482318f
C62 VN.n25 B 1.65779f
C63 VTAIL.t3 B 0.168821f
C64 VTAIL.t13 B 0.168821f
C65 VTAIL.n0 B 1.45242f
C66 VTAIL.n1 B 0.25344f
C67 VTAIL.t15 B 1.84995f
C68 VTAIL.n2 B 0.342379f
C69 VTAIL.t7 B 1.84995f
C70 VTAIL.n3 B 0.342379f
C71 VTAIL.t5 B 0.168821f
C72 VTAIL.t8 B 0.168821f
C73 VTAIL.n4 B 1.45242f
C74 VTAIL.n5 B 0.322301f
C75 VTAIL.t9 B 1.84995f
C76 VTAIL.n6 B 1.24536f
C77 VTAIL.t0 B 1.84995f
C78 VTAIL.n7 B 1.24536f
C79 VTAIL.t2 B 0.168821f
C80 VTAIL.t4 B 0.168821f
C81 VTAIL.n8 B 1.45242f
C82 VTAIL.n9 B 0.322307f
C83 VTAIL.t14 B 1.84995f
C84 VTAIL.n10 B 0.342383f
C85 VTAIL.t6 B 1.84995f
C86 VTAIL.n11 B 0.342383f
C87 VTAIL.t11 B 0.168821f
C88 VTAIL.t12 B 0.168821f
C89 VTAIL.n12 B 1.45242f
C90 VTAIL.n13 B 0.322307f
C91 VTAIL.t10 B 1.84994f
C92 VTAIL.n14 B 1.24536f
C93 VTAIL.t1 B 1.84995f
C94 VTAIL.n15 B 1.24167f
C95 VDD1.t2 B 0.223f
C96 VDD1.t5 B 0.223f
C97 VDD1.n0 B 1.98949f
C98 VDD1.t0 B 0.223f
C99 VDD1.t1 B 0.223f
C100 VDD1.n1 B 1.98882f
C101 VDD1.t3 B 0.223f
C102 VDD1.t4 B 0.223f
C103 VDD1.n2 B 1.98882f
C104 VDD1.n3 B 2.39639f
C105 VDD1.t6 B 0.223f
C106 VDD1.t7 B 0.223f
C107 VDD1.n4 B 1.98603f
C108 VDD1.n5 B 2.41321f
C109 VP.n0 B 0.051647f
C110 VP.t4 B 1.144f
C111 VP.n1 B 0.031321f
C112 VP.n2 B 0.051647f
C113 VP.t7 B 1.144f
C114 VP.n3 B 0.051647f
C115 VP.t2 B 1.20366f
C116 VP.t0 B 1.144f
C117 VP.n4 B 0.031321f
C118 VP.t6 B 1.22719f
C119 VP.n5 B 0.485409f
C120 VP.t1 B 1.144f
C121 VP.n6 B 0.464049f
C122 VP.n7 B 0.053354f
C123 VP.n8 B 0.165696f
C124 VP.n9 B 0.038705f
C125 VP.n10 B 0.038705f
C126 VP.n11 B 0.053354f
C127 VP.n12 B 0.429181f
C128 VP.n13 B 0.053578f
C129 VP.n14 B 0.489411f
C130 VP.n15 B 1.66053f
C131 VP.n16 B 1.69296f
C132 VP.t3 B 1.20366f
C133 VP.n17 B 0.489411f
C134 VP.n18 B 0.053578f
C135 VP.n19 B 0.429181f
C136 VP.n20 B 0.053354f
C137 VP.n21 B 0.038705f
C138 VP.n22 B 0.038705f
C139 VP.n23 B 0.038705f
C140 VP.n24 B 0.053354f
C141 VP.n25 B 0.429181f
C142 VP.n26 B 0.053578f
C143 VP.t5 B 1.20366f
C144 VP.n27 B 0.489411f
C145 VP.n28 B 0.036249f
.ends

