* NGSPICE file created from diff_pair_sample_1728.ext - technology: sky130A

.subckt diff_pair_sample_1728 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X1 VTAIL.t14 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=3.19
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=3.19
X3 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=3.19
X4 VDD1.t5 VP.t2 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=3.19
X5 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X6 VTAIL.t8 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X7 VTAIL.t7 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=3.19
X8 VTAIL.t15 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X9 VTAIL.t12 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=3.19
X10 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=3.19
X11 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=3.19
X12 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X13 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X14 VTAIL.t0 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=3.19
X15 VDD1.t1 VP.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=3.19
X16 VDD1.t0 VP.t7 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X17 VDD2.t0 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=3.19
X18 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=3.19
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=3.19
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n33 VP.n32 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n16 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n39 VP.n15 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n42 VP.n14 161.3
R13 VP.n44 VP.n43 161.3
R14 VP.n79 VP.n78 161.3
R15 VP.n77 VP.n1 161.3
R16 VP.n76 VP.n75 161.3
R17 VP.n74 VP.n2 161.3
R18 VP.n73 VP.n72 161.3
R19 VP.n71 VP.n3 161.3
R20 VP.n70 VP.n69 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n66 VP.n5 161.3
R23 VP.n65 VP.n64 161.3
R24 VP.n63 VP.n6 161.3
R25 VP.n62 VP.n61 161.3
R26 VP.n60 VP.n7 161.3
R27 VP.n59 VP.n58 161.3
R28 VP.n57 VP.n56 161.3
R29 VP.n55 VP.n9 161.3
R30 VP.n54 VP.n53 161.3
R31 VP.n52 VP.n10 161.3
R32 VP.n51 VP.n50 161.3
R33 VP.n49 VP.n11 161.3
R34 VP.n48 VP.n47 161.3
R35 VP.n22 VP.t5 132.793
R36 VP.n12 VP.t1 99.9513
R37 VP.n8 VP.t0 99.9513
R38 VP.n4 VP.t4 99.9513
R39 VP.n0 VP.t2 99.9513
R40 VP.n13 VP.t6 99.9513
R41 VP.n17 VP.t3 99.9513
R42 VP.n21 VP.t7 99.9513
R43 VP.n46 VP.n12 76.3659
R44 VP.n80 VP.n0 76.3659
R45 VP.n45 VP.n13 76.3659
R46 VP.n22 VP.n21 61.5301
R47 VP.n46 VP.n45 54.6584
R48 VP.n50 VP.n10 42.4359
R49 VP.n76 VP.n2 42.4359
R50 VP.n41 VP.n15 42.4359
R51 VP.n61 VP.n6 40.4934
R52 VP.n65 VP.n6 40.4934
R53 VP.n30 VP.n19 40.4934
R54 VP.n26 VP.n19 40.4934
R55 VP.n54 VP.n10 38.5509
R56 VP.n72 VP.n2 38.5509
R57 VP.n37 VP.n15 38.5509
R58 VP.n49 VP.n48 24.4675
R59 VP.n50 VP.n49 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n55 24.4675
R62 VP.n60 VP.n59 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n66 VP.n65 24.4675
R65 VP.n67 VP.n66 24.4675
R66 VP.n71 VP.n70 24.4675
R67 VP.n72 VP.n71 24.4675
R68 VP.n77 VP.n76 24.4675
R69 VP.n78 VP.n77 24.4675
R70 VP.n42 VP.n41 24.4675
R71 VP.n43 VP.n42 24.4675
R72 VP.n31 VP.n30 24.4675
R73 VP.n32 VP.n31 24.4675
R74 VP.n36 VP.n35 24.4675
R75 VP.n37 VP.n36 24.4675
R76 VP.n25 VP.n24 24.4675
R77 VP.n26 VP.n25 24.4675
R78 VP.n48 VP.n12 13.702
R79 VP.n78 VP.n0 13.702
R80 VP.n43 VP.n13 13.702
R81 VP.n59 VP.n8 12.7233
R82 VP.n67 VP.n4 12.7233
R83 VP.n32 VP.n17 12.7233
R84 VP.n24 VP.n21 12.7233
R85 VP.n56 VP.n8 11.7447
R86 VP.n70 VP.n4 11.7447
R87 VP.n35 VP.n17 11.7447
R88 VP.n23 VP.n22 4.2058
R89 VP.n45 VP.n44 0.354971
R90 VP.n47 VP.n46 0.354971
R91 VP.n80 VP.n79 0.354971
R92 VP VP.n80 0.26696
R93 VP.n23 VP.n20 0.189894
R94 VP.n27 VP.n20 0.189894
R95 VP.n28 VP.n27 0.189894
R96 VP.n29 VP.n28 0.189894
R97 VP.n29 VP.n18 0.189894
R98 VP.n33 VP.n18 0.189894
R99 VP.n34 VP.n33 0.189894
R100 VP.n34 VP.n16 0.189894
R101 VP.n38 VP.n16 0.189894
R102 VP.n39 VP.n38 0.189894
R103 VP.n40 VP.n39 0.189894
R104 VP.n40 VP.n14 0.189894
R105 VP.n44 VP.n14 0.189894
R106 VP.n47 VP.n11 0.189894
R107 VP.n51 VP.n11 0.189894
R108 VP.n52 VP.n51 0.189894
R109 VP.n53 VP.n52 0.189894
R110 VP.n53 VP.n9 0.189894
R111 VP.n57 VP.n9 0.189894
R112 VP.n58 VP.n57 0.189894
R113 VP.n58 VP.n7 0.189894
R114 VP.n62 VP.n7 0.189894
R115 VP.n63 VP.n62 0.189894
R116 VP.n64 VP.n63 0.189894
R117 VP.n64 VP.n5 0.189894
R118 VP.n68 VP.n5 0.189894
R119 VP.n69 VP.n68 0.189894
R120 VP.n69 VP.n3 0.189894
R121 VP.n73 VP.n3 0.189894
R122 VP.n74 VP.n73 0.189894
R123 VP.n75 VP.n74 0.189894
R124 VP.n75 VP.n1 0.189894
R125 VP.n79 VP.n1 0.189894
R126 VTAIL.n11 VTAIL.t12 47.0249
R127 VTAIL.n10 VTAIL.t5 47.0249
R128 VTAIL.n7 VTAIL.t7 47.0249
R129 VTAIL.n15 VTAIL.t3 47.0247
R130 VTAIL.n2 VTAIL.t0 47.0247
R131 VTAIL.n3 VTAIL.t11 47.0247
R132 VTAIL.n6 VTAIL.t14 47.0247
R133 VTAIL.n14 VTAIL.t9 47.0247
R134 VTAIL.n13 VTAIL.n12 45.5283
R135 VTAIL.n9 VTAIL.n8 45.5283
R136 VTAIL.n1 VTAIL.n0 45.5283
R137 VTAIL.n5 VTAIL.n4 45.5283
R138 VTAIL.n15 VTAIL.n14 26.8065
R139 VTAIL.n7 VTAIL.n6 26.8065
R140 VTAIL.n9 VTAIL.n7 3.03498
R141 VTAIL.n10 VTAIL.n9 3.03498
R142 VTAIL.n13 VTAIL.n11 3.03498
R143 VTAIL.n14 VTAIL.n13 3.03498
R144 VTAIL.n6 VTAIL.n5 3.03498
R145 VTAIL.n5 VTAIL.n3 3.03498
R146 VTAIL.n2 VTAIL.n1 3.03498
R147 VTAIL VTAIL.n15 2.97679
R148 VTAIL.n0 VTAIL.t4 1.4971
R149 VTAIL.n0 VTAIL.t1 1.4971
R150 VTAIL.n4 VTAIL.t10 1.4971
R151 VTAIL.n4 VTAIL.t15 1.4971
R152 VTAIL.n12 VTAIL.t13 1.4971
R153 VTAIL.n12 VTAIL.t8 1.4971
R154 VTAIL.n8 VTAIL.t2 1.4971
R155 VTAIL.n8 VTAIL.t6 1.4971
R156 VTAIL.n11 VTAIL.n10 0.470328
R157 VTAIL.n3 VTAIL.n2 0.470328
R158 VTAIL VTAIL.n1 0.0586897
R159 VDD1 VDD1.n0 63.7826
R160 VDD1.n3 VDD1.n2 63.669
R161 VDD1.n3 VDD1.n1 63.669
R162 VDD1.n5 VDD1.n4 62.2069
R163 VDD1.n5 VDD1.n3 49.3587
R164 VDD1.n4 VDD1.t4 1.4971
R165 VDD1.n4 VDD1.t1 1.4971
R166 VDD1.n0 VDD1.t2 1.4971
R167 VDD1.n0 VDD1.t0 1.4971
R168 VDD1.n2 VDD1.t3 1.4971
R169 VDD1.n2 VDD1.t5 1.4971
R170 VDD1.n1 VDD1.t6 1.4971
R171 VDD1.n1 VDD1.t7 1.4971
R172 VDD1 VDD1.n5 1.45955
R173 B.n992 B.n991 585
R174 B.n361 B.n160 585
R175 B.n360 B.n359 585
R176 B.n358 B.n357 585
R177 B.n356 B.n355 585
R178 B.n354 B.n353 585
R179 B.n352 B.n351 585
R180 B.n350 B.n349 585
R181 B.n348 B.n347 585
R182 B.n346 B.n345 585
R183 B.n344 B.n343 585
R184 B.n342 B.n341 585
R185 B.n340 B.n339 585
R186 B.n338 B.n337 585
R187 B.n336 B.n335 585
R188 B.n334 B.n333 585
R189 B.n332 B.n331 585
R190 B.n330 B.n329 585
R191 B.n328 B.n327 585
R192 B.n326 B.n325 585
R193 B.n324 B.n323 585
R194 B.n322 B.n321 585
R195 B.n320 B.n319 585
R196 B.n318 B.n317 585
R197 B.n316 B.n315 585
R198 B.n314 B.n313 585
R199 B.n312 B.n311 585
R200 B.n310 B.n309 585
R201 B.n308 B.n307 585
R202 B.n306 B.n305 585
R203 B.n304 B.n303 585
R204 B.n302 B.n301 585
R205 B.n300 B.n299 585
R206 B.n298 B.n297 585
R207 B.n296 B.n295 585
R208 B.n294 B.n293 585
R209 B.n292 B.n291 585
R210 B.n290 B.n289 585
R211 B.n288 B.n287 585
R212 B.n286 B.n285 585
R213 B.n284 B.n283 585
R214 B.n282 B.n281 585
R215 B.n280 B.n279 585
R216 B.n278 B.n277 585
R217 B.n276 B.n275 585
R218 B.n273 B.n272 585
R219 B.n271 B.n270 585
R220 B.n269 B.n268 585
R221 B.n267 B.n266 585
R222 B.n265 B.n264 585
R223 B.n263 B.n262 585
R224 B.n261 B.n260 585
R225 B.n259 B.n258 585
R226 B.n257 B.n256 585
R227 B.n255 B.n254 585
R228 B.n252 B.n251 585
R229 B.n250 B.n249 585
R230 B.n248 B.n247 585
R231 B.n246 B.n245 585
R232 B.n244 B.n243 585
R233 B.n242 B.n241 585
R234 B.n240 B.n239 585
R235 B.n238 B.n237 585
R236 B.n236 B.n235 585
R237 B.n234 B.n233 585
R238 B.n232 B.n231 585
R239 B.n230 B.n229 585
R240 B.n228 B.n227 585
R241 B.n226 B.n225 585
R242 B.n224 B.n223 585
R243 B.n222 B.n221 585
R244 B.n220 B.n219 585
R245 B.n218 B.n217 585
R246 B.n216 B.n215 585
R247 B.n214 B.n213 585
R248 B.n212 B.n211 585
R249 B.n210 B.n209 585
R250 B.n208 B.n207 585
R251 B.n206 B.n205 585
R252 B.n204 B.n203 585
R253 B.n202 B.n201 585
R254 B.n200 B.n199 585
R255 B.n198 B.n197 585
R256 B.n196 B.n195 585
R257 B.n194 B.n193 585
R258 B.n192 B.n191 585
R259 B.n190 B.n189 585
R260 B.n188 B.n187 585
R261 B.n186 B.n185 585
R262 B.n184 B.n183 585
R263 B.n182 B.n181 585
R264 B.n180 B.n179 585
R265 B.n178 B.n177 585
R266 B.n176 B.n175 585
R267 B.n174 B.n173 585
R268 B.n172 B.n171 585
R269 B.n170 B.n169 585
R270 B.n168 B.n167 585
R271 B.n166 B.n165 585
R272 B.n109 B.n108 585
R273 B.n990 B.n110 585
R274 B.n995 B.n110 585
R275 B.n989 B.n988 585
R276 B.n988 B.n106 585
R277 B.n987 B.n105 585
R278 B.n1001 B.n105 585
R279 B.n986 B.n104 585
R280 B.n1002 B.n104 585
R281 B.n985 B.n103 585
R282 B.n1003 B.n103 585
R283 B.n984 B.n983 585
R284 B.n983 B.n99 585
R285 B.n982 B.n98 585
R286 B.n1009 B.n98 585
R287 B.n981 B.n97 585
R288 B.n1010 B.n97 585
R289 B.n980 B.n96 585
R290 B.n1011 B.n96 585
R291 B.n979 B.n978 585
R292 B.n978 B.n92 585
R293 B.n977 B.n91 585
R294 B.n1017 B.n91 585
R295 B.n976 B.n90 585
R296 B.n1018 B.n90 585
R297 B.n975 B.n89 585
R298 B.n1019 B.n89 585
R299 B.n974 B.n973 585
R300 B.n973 B.n85 585
R301 B.n972 B.n84 585
R302 B.n1025 B.n84 585
R303 B.n971 B.n83 585
R304 B.n1026 B.n83 585
R305 B.n970 B.n82 585
R306 B.n1027 B.n82 585
R307 B.n969 B.n968 585
R308 B.n968 B.n78 585
R309 B.n967 B.n77 585
R310 B.n1033 B.n77 585
R311 B.n966 B.n76 585
R312 B.n1034 B.n76 585
R313 B.n965 B.n75 585
R314 B.n1035 B.n75 585
R315 B.n964 B.n963 585
R316 B.n963 B.n71 585
R317 B.n962 B.n70 585
R318 B.n1041 B.n70 585
R319 B.n961 B.n69 585
R320 B.n1042 B.n69 585
R321 B.n960 B.n68 585
R322 B.n1043 B.n68 585
R323 B.n959 B.n958 585
R324 B.n958 B.n64 585
R325 B.n957 B.n63 585
R326 B.n1049 B.n63 585
R327 B.n956 B.n62 585
R328 B.n1050 B.n62 585
R329 B.n955 B.n61 585
R330 B.n1051 B.n61 585
R331 B.n954 B.n953 585
R332 B.n953 B.n57 585
R333 B.n952 B.n56 585
R334 B.n1057 B.n56 585
R335 B.n951 B.n55 585
R336 B.n1058 B.n55 585
R337 B.n950 B.n54 585
R338 B.n1059 B.n54 585
R339 B.n949 B.n948 585
R340 B.n948 B.n50 585
R341 B.n947 B.n49 585
R342 B.n1065 B.n49 585
R343 B.n946 B.n48 585
R344 B.n1066 B.n48 585
R345 B.n945 B.n47 585
R346 B.n1067 B.n47 585
R347 B.n944 B.n943 585
R348 B.n943 B.n43 585
R349 B.n942 B.n42 585
R350 B.n1073 B.n42 585
R351 B.n941 B.n41 585
R352 B.n1074 B.n41 585
R353 B.n940 B.n40 585
R354 B.n1075 B.n40 585
R355 B.n939 B.n938 585
R356 B.n938 B.n36 585
R357 B.n937 B.n35 585
R358 B.n1081 B.n35 585
R359 B.n936 B.n34 585
R360 B.n1082 B.n34 585
R361 B.n935 B.n33 585
R362 B.n1083 B.n33 585
R363 B.n934 B.n933 585
R364 B.n933 B.n29 585
R365 B.n932 B.n28 585
R366 B.n1089 B.n28 585
R367 B.n931 B.n27 585
R368 B.n1090 B.n27 585
R369 B.n930 B.n26 585
R370 B.n1091 B.n26 585
R371 B.n929 B.n928 585
R372 B.n928 B.n22 585
R373 B.n927 B.n21 585
R374 B.n1097 B.n21 585
R375 B.n926 B.n20 585
R376 B.n1098 B.n20 585
R377 B.n925 B.n19 585
R378 B.n1099 B.n19 585
R379 B.n924 B.n923 585
R380 B.n923 B.n18 585
R381 B.n922 B.n14 585
R382 B.n1105 B.n14 585
R383 B.n921 B.n13 585
R384 B.n1106 B.n13 585
R385 B.n920 B.n12 585
R386 B.n1107 B.n12 585
R387 B.n919 B.n918 585
R388 B.n918 B.n8 585
R389 B.n917 B.n7 585
R390 B.n1113 B.n7 585
R391 B.n916 B.n6 585
R392 B.n1114 B.n6 585
R393 B.n915 B.n5 585
R394 B.n1115 B.n5 585
R395 B.n914 B.n913 585
R396 B.n913 B.n4 585
R397 B.n912 B.n362 585
R398 B.n912 B.n911 585
R399 B.n902 B.n363 585
R400 B.n364 B.n363 585
R401 B.n904 B.n903 585
R402 B.n905 B.n904 585
R403 B.n901 B.n369 585
R404 B.n369 B.n368 585
R405 B.n900 B.n899 585
R406 B.n899 B.n898 585
R407 B.n371 B.n370 585
R408 B.n891 B.n371 585
R409 B.n890 B.n889 585
R410 B.n892 B.n890 585
R411 B.n888 B.n376 585
R412 B.n376 B.n375 585
R413 B.n887 B.n886 585
R414 B.n886 B.n885 585
R415 B.n378 B.n377 585
R416 B.n379 B.n378 585
R417 B.n878 B.n877 585
R418 B.n879 B.n878 585
R419 B.n876 B.n384 585
R420 B.n384 B.n383 585
R421 B.n875 B.n874 585
R422 B.n874 B.n873 585
R423 B.n386 B.n385 585
R424 B.n387 B.n386 585
R425 B.n866 B.n865 585
R426 B.n867 B.n866 585
R427 B.n864 B.n392 585
R428 B.n392 B.n391 585
R429 B.n863 B.n862 585
R430 B.n862 B.n861 585
R431 B.n394 B.n393 585
R432 B.n395 B.n394 585
R433 B.n854 B.n853 585
R434 B.n855 B.n854 585
R435 B.n852 B.n400 585
R436 B.n400 B.n399 585
R437 B.n851 B.n850 585
R438 B.n850 B.n849 585
R439 B.n402 B.n401 585
R440 B.n403 B.n402 585
R441 B.n842 B.n841 585
R442 B.n843 B.n842 585
R443 B.n840 B.n408 585
R444 B.n408 B.n407 585
R445 B.n839 B.n838 585
R446 B.n838 B.n837 585
R447 B.n410 B.n409 585
R448 B.n411 B.n410 585
R449 B.n830 B.n829 585
R450 B.n831 B.n830 585
R451 B.n828 B.n416 585
R452 B.n416 B.n415 585
R453 B.n827 B.n826 585
R454 B.n826 B.n825 585
R455 B.n418 B.n417 585
R456 B.n419 B.n418 585
R457 B.n818 B.n817 585
R458 B.n819 B.n818 585
R459 B.n816 B.n424 585
R460 B.n424 B.n423 585
R461 B.n815 B.n814 585
R462 B.n814 B.n813 585
R463 B.n426 B.n425 585
R464 B.n427 B.n426 585
R465 B.n806 B.n805 585
R466 B.n807 B.n806 585
R467 B.n804 B.n432 585
R468 B.n432 B.n431 585
R469 B.n803 B.n802 585
R470 B.n802 B.n801 585
R471 B.n434 B.n433 585
R472 B.n435 B.n434 585
R473 B.n794 B.n793 585
R474 B.n795 B.n794 585
R475 B.n792 B.n440 585
R476 B.n440 B.n439 585
R477 B.n791 B.n790 585
R478 B.n790 B.n789 585
R479 B.n442 B.n441 585
R480 B.n443 B.n442 585
R481 B.n782 B.n781 585
R482 B.n783 B.n782 585
R483 B.n780 B.n448 585
R484 B.n448 B.n447 585
R485 B.n779 B.n778 585
R486 B.n778 B.n777 585
R487 B.n450 B.n449 585
R488 B.n451 B.n450 585
R489 B.n770 B.n769 585
R490 B.n771 B.n770 585
R491 B.n768 B.n456 585
R492 B.n456 B.n455 585
R493 B.n767 B.n766 585
R494 B.n766 B.n765 585
R495 B.n458 B.n457 585
R496 B.n459 B.n458 585
R497 B.n758 B.n757 585
R498 B.n759 B.n758 585
R499 B.n756 B.n464 585
R500 B.n464 B.n463 585
R501 B.n755 B.n754 585
R502 B.n754 B.n753 585
R503 B.n466 B.n465 585
R504 B.n467 B.n466 585
R505 B.n746 B.n745 585
R506 B.n747 B.n746 585
R507 B.n744 B.n472 585
R508 B.n472 B.n471 585
R509 B.n743 B.n742 585
R510 B.n742 B.n741 585
R511 B.n474 B.n473 585
R512 B.n475 B.n474 585
R513 B.n734 B.n733 585
R514 B.n735 B.n734 585
R515 B.n478 B.n477 585
R516 B.n537 B.n536 585
R517 B.n538 B.n534 585
R518 B.n534 B.n479 585
R519 B.n540 B.n539 585
R520 B.n542 B.n533 585
R521 B.n545 B.n544 585
R522 B.n546 B.n532 585
R523 B.n548 B.n547 585
R524 B.n550 B.n531 585
R525 B.n553 B.n552 585
R526 B.n554 B.n530 585
R527 B.n556 B.n555 585
R528 B.n558 B.n529 585
R529 B.n561 B.n560 585
R530 B.n562 B.n528 585
R531 B.n564 B.n563 585
R532 B.n566 B.n527 585
R533 B.n569 B.n568 585
R534 B.n570 B.n526 585
R535 B.n572 B.n571 585
R536 B.n574 B.n525 585
R537 B.n577 B.n576 585
R538 B.n578 B.n524 585
R539 B.n580 B.n579 585
R540 B.n582 B.n523 585
R541 B.n585 B.n584 585
R542 B.n586 B.n522 585
R543 B.n588 B.n587 585
R544 B.n590 B.n521 585
R545 B.n593 B.n592 585
R546 B.n594 B.n520 585
R547 B.n596 B.n595 585
R548 B.n598 B.n519 585
R549 B.n601 B.n600 585
R550 B.n602 B.n518 585
R551 B.n604 B.n603 585
R552 B.n606 B.n517 585
R553 B.n609 B.n608 585
R554 B.n610 B.n516 585
R555 B.n612 B.n611 585
R556 B.n614 B.n515 585
R557 B.n617 B.n616 585
R558 B.n618 B.n514 585
R559 B.n620 B.n619 585
R560 B.n622 B.n513 585
R561 B.n625 B.n624 585
R562 B.n626 B.n509 585
R563 B.n628 B.n627 585
R564 B.n630 B.n508 585
R565 B.n633 B.n632 585
R566 B.n634 B.n507 585
R567 B.n636 B.n635 585
R568 B.n638 B.n506 585
R569 B.n641 B.n640 585
R570 B.n642 B.n503 585
R571 B.n645 B.n644 585
R572 B.n647 B.n502 585
R573 B.n650 B.n649 585
R574 B.n651 B.n501 585
R575 B.n653 B.n652 585
R576 B.n655 B.n500 585
R577 B.n658 B.n657 585
R578 B.n659 B.n499 585
R579 B.n661 B.n660 585
R580 B.n663 B.n498 585
R581 B.n666 B.n665 585
R582 B.n667 B.n497 585
R583 B.n669 B.n668 585
R584 B.n671 B.n496 585
R585 B.n674 B.n673 585
R586 B.n675 B.n495 585
R587 B.n677 B.n676 585
R588 B.n679 B.n494 585
R589 B.n682 B.n681 585
R590 B.n683 B.n493 585
R591 B.n685 B.n684 585
R592 B.n687 B.n492 585
R593 B.n690 B.n689 585
R594 B.n691 B.n491 585
R595 B.n693 B.n692 585
R596 B.n695 B.n490 585
R597 B.n698 B.n697 585
R598 B.n699 B.n489 585
R599 B.n701 B.n700 585
R600 B.n703 B.n488 585
R601 B.n706 B.n705 585
R602 B.n707 B.n487 585
R603 B.n709 B.n708 585
R604 B.n711 B.n486 585
R605 B.n714 B.n713 585
R606 B.n715 B.n485 585
R607 B.n717 B.n716 585
R608 B.n719 B.n484 585
R609 B.n722 B.n721 585
R610 B.n723 B.n483 585
R611 B.n725 B.n724 585
R612 B.n727 B.n482 585
R613 B.n728 B.n481 585
R614 B.n731 B.n730 585
R615 B.n732 B.n480 585
R616 B.n480 B.n479 585
R617 B.n737 B.n736 585
R618 B.n736 B.n735 585
R619 B.n738 B.n476 585
R620 B.n476 B.n475 585
R621 B.n740 B.n739 585
R622 B.n741 B.n740 585
R623 B.n470 B.n469 585
R624 B.n471 B.n470 585
R625 B.n749 B.n748 585
R626 B.n748 B.n747 585
R627 B.n750 B.n468 585
R628 B.n468 B.n467 585
R629 B.n752 B.n751 585
R630 B.n753 B.n752 585
R631 B.n462 B.n461 585
R632 B.n463 B.n462 585
R633 B.n761 B.n760 585
R634 B.n760 B.n759 585
R635 B.n762 B.n460 585
R636 B.n460 B.n459 585
R637 B.n764 B.n763 585
R638 B.n765 B.n764 585
R639 B.n454 B.n453 585
R640 B.n455 B.n454 585
R641 B.n773 B.n772 585
R642 B.n772 B.n771 585
R643 B.n774 B.n452 585
R644 B.n452 B.n451 585
R645 B.n776 B.n775 585
R646 B.n777 B.n776 585
R647 B.n446 B.n445 585
R648 B.n447 B.n446 585
R649 B.n785 B.n784 585
R650 B.n784 B.n783 585
R651 B.n786 B.n444 585
R652 B.n444 B.n443 585
R653 B.n788 B.n787 585
R654 B.n789 B.n788 585
R655 B.n438 B.n437 585
R656 B.n439 B.n438 585
R657 B.n797 B.n796 585
R658 B.n796 B.n795 585
R659 B.n798 B.n436 585
R660 B.n436 B.n435 585
R661 B.n800 B.n799 585
R662 B.n801 B.n800 585
R663 B.n430 B.n429 585
R664 B.n431 B.n430 585
R665 B.n809 B.n808 585
R666 B.n808 B.n807 585
R667 B.n810 B.n428 585
R668 B.n428 B.n427 585
R669 B.n812 B.n811 585
R670 B.n813 B.n812 585
R671 B.n422 B.n421 585
R672 B.n423 B.n422 585
R673 B.n821 B.n820 585
R674 B.n820 B.n819 585
R675 B.n822 B.n420 585
R676 B.n420 B.n419 585
R677 B.n824 B.n823 585
R678 B.n825 B.n824 585
R679 B.n414 B.n413 585
R680 B.n415 B.n414 585
R681 B.n833 B.n832 585
R682 B.n832 B.n831 585
R683 B.n834 B.n412 585
R684 B.n412 B.n411 585
R685 B.n836 B.n835 585
R686 B.n837 B.n836 585
R687 B.n406 B.n405 585
R688 B.n407 B.n406 585
R689 B.n845 B.n844 585
R690 B.n844 B.n843 585
R691 B.n846 B.n404 585
R692 B.n404 B.n403 585
R693 B.n848 B.n847 585
R694 B.n849 B.n848 585
R695 B.n398 B.n397 585
R696 B.n399 B.n398 585
R697 B.n857 B.n856 585
R698 B.n856 B.n855 585
R699 B.n858 B.n396 585
R700 B.n396 B.n395 585
R701 B.n860 B.n859 585
R702 B.n861 B.n860 585
R703 B.n390 B.n389 585
R704 B.n391 B.n390 585
R705 B.n869 B.n868 585
R706 B.n868 B.n867 585
R707 B.n870 B.n388 585
R708 B.n388 B.n387 585
R709 B.n872 B.n871 585
R710 B.n873 B.n872 585
R711 B.n382 B.n381 585
R712 B.n383 B.n382 585
R713 B.n881 B.n880 585
R714 B.n880 B.n879 585
R715 B.n882 B.n380 585
R716 B.n380 B.n379 585
R717 B.n884 B.n883 585
R718 B.n885 B.n884 585
R719 B.n374 B.n373 585
R720 B.n375 B.n374 585
R721 B.n894 B.n893 585
R722 B.n893 B.n892 585
R723 B.n895 B.n372 585
R724 B.n891 B.n372 585
R725 B.n897 B.n896 585
R726 B.n898 B.n897 585
R727 B.n367 B.n366 585
R728 B.n368 B.n367 585
R729 B.n907 B.n906 585
R730 B.n906 B.n905 585
R731 B.n908 B.n365 585
R732 B.n365 B.n364 585
R733 B.n910 B.n909 585
R734 B.n911 B.n910 585
R735 B.n2 B.n0 585
R736 B.n4 B.n2 585
R737 B.n3 B.n1 585
R738 B.n1114 B.n3 585
R739 B.n1112 B.n1111 585
R740 B.n1113 B.n1112 585
R741 B.n1110 B.n9 585
R742 B.n9 B.n8 585
R743 B.n1109 B.n1108 585
R744 B.n1108 B.n1107 585
R745 B.n11 B.n10 585
R746 B.n1106 B.n11 585
R747 B.n1104 B.n1103 585
R748 B.n1105 B.n1104 585
R749 B.n1102 B.n15 585
R750 B.n18 B.n15 585
R751 B.n1101 B.n1100 585
R752 B.n1100 B.n1099 585
R753 B.n17 B.n16 585
R754 B.n1098 B.n17 585
R755 B.n1096 B.n1095 585
R756 B.n1097 B.n1096 585
R757 B.n1094 B.n23 585
R758 B.n23 B.n22 585
R759 B.n1093 B.n1092 585
R760 B.n1092 B.n1091 585
R761 B.n25 B.n24 585
R762 B.n1090 B.n25 585
R763 B.n1088 B.n1087 585
R764 B.n1089 B.n1088 585
R765 B.n1086 B.n30 585
R766 B.n30 B.n29 585
R767 B.n1085 B.n1084 585
R768 B.n1084 B.n1083 585
R769 B.n32 B.n31 585
R770 B.n1082 B.n32 585
R771 B.n1080 B.n1079 585
R772 B.n1081 B.n1080 585
R773 B.n1078 B.n37 585
R774 B.n37 B.n36 585
R775 B.n1077 B.n1076 585
R776 B.n1076 B.n1075 585
R777 B.n39 B.n38 585
R778 B.n1074 B.n39 585
R779 B.n1072 B.n1071 585
R780 B.n1073 B.n1072 585
R781 B.n1070 B.n44 585
R782 B.n44 B.n43 585
R783 B.n1069 B.n1068 585
R784 B.n1068 B.n1067 585
R785 B.n46 B.n45 585
R786 B.n1066 B.n46 585
R787 B.n1064 B.n1063 585
R788 B.n1065 B.n1064 585
R789 B.n1062 B.n51 585
R790 B.n51 B.n50 585
R791 B.n1061 B.n1060 585
R792 B.n1060 B.n1059 585
R793 B.n53 B.n52 585
R794 B.n1058 B.n53 585
R795 B.n1056 B.n1055 585
R796 B.n1057 B.n1056 585
R797 B.n1054 B.n58 585
R798 B.n58 B.n57 585
R799 B.n1053 B.n1052 585
R800 B.n1052 B.n1051 585
R801 B.n60 B.n59 585
R802 B.n1050 B.n60 585
R803 B.n1048 B.n1047 585
R804 B.n1049 B.n1048 585
R805 B.n1046 B.n65 585
R806 B.n65 B.n64 585
R807 B.n1045 B.n1044 585
R808 B.n1044 B.n1043 585
R809 B.n67 B.n66 585
R810 B.n1042 B.n67 585
R811 B.n1040 B.n1039 585
R812 B.n1041 B.n1040 585
R813 B.n1038 B.n72 585
R814 B.n72 B.n71 585
R815 B.n1037 B.n1036 585
R816 B.n1036 B.n1035 585
R817 B.n74 B.n73 585
R818 B.n1034 B.n74 585
R819 B.n1032 B.n1031 585
R820 B.n1033 B.n1032 585
R821 B.n1030 B.n79 585
R822 B.n79 B.n78 585
R823 B.n1029 B.n1028 585
R824 B.n1028 B.n1027 585
R825 B.n81 B.n80 585
R826 B.n1026 B.n81 585
R827 B.n1024 B.n1023 585
R828 B.n1025 B.n1024 585
R829 B.n1022 B.n86 585
R830 B.n86 B.n85 585
R831 B.n1021 B.n1020 585
R832 B.n1020 B.n1019 585
R833 B.n88 B.n87 585
R834 B.n1018 B.n88 585
R835 B.n1016 B.n1015 585
R836 B.n1017 B.n1016 585
R837 B.n1014 B.n93 585
R838 B.n93 B.n92 585
R839 B.n1013 B.n1012 585
R840 B.n1012 B.n1011 585
R841 B.n95 B.n94 585
R842 B.n1010 B.n95 585
R843 B.n1008 B.n1007 585
R844 B.n1009 B.n1008 585
R845 B.n1006 B.n100 585
R846 B.n100 B.n99 585
R847 B.n1005 B.n1004 585
R848 B.n1004 B.n1003 585
R849 B.n102 B.n101 585
R850 B.n1002 B.n102 585
R851 B.n1000 B.n999 585
R852 B.n1001 B.n1000 585
R853 B.n998 B.n107 585
R854 B.n107 B.n106 585
R855 B.n997 B.n996 585
R856 B.n996 B.n995 585
R857 B.n1117 B.n1116 585
R858 B.n1116 B.n1115 585
R859 B.n736 B.n478 482.89
R860 B.n996 B.n109 482.89
R861 B.n734 B.n480 482.89
R862 B.n992 B.n110 482.89
R863 B.n504 B.t19 308.743
R864 B.n510 B.t15 308.743
R865 B.n163 B.t12 308.743
R866 B.n161 B.t8 308.743
R867 B.n994 B.n993 256.663
R868 B.n994 B.n159 256.663
R869 B.n994 B.n158 256.663
R870 B.n994 B.n157 256.663
R871 B.n994 B.n156 256.663
R872 B.n994 B.n155 256.663
R873 B.n994 B.n154 256.663
R874 B.n994 B.n153 256.663
R875 B.n994 B.n152 256.663
R876 B.n994 B.n151 256.663
R877 B.n994 B.n150 256.663
R878 B.n994 B.n149 256.663
R879 B.n994 B.n148 256.663
R880 B.n994 B.n147 256.663
R881 B.n994 B.n146 256.663
R882 B.n994 B.n145 256.663
R883 B.n994 B.n144 256.663
R884 B.n994 B.n143 256.663
R885 B.n994 B.n142 256.663
R886 B.n994 B.n141 256.663
R887 B.n994 B.n140 256.663
R888 B.n994 B.n139 256.663
R889 B.n994 B.n138 256.663
R890 B.n994 B.n137 256.663
R891 B.n994 B.n136 256.663
R892 B.n994 B.n135 256.663
R893 B.n994 B.n134 256.663
R894 B.n994 B.n133 256.663
R895 B.n994 B.n132 256.663
R896 B.n994 B.n131 256.663
R897 B.n994 B.n130 256.663
R898 B.n994 B.n129 256.663
R899 B.n994 B.n128 256.663
R900 B.n994 B.n127 256.663
R901 B.n994 B.n126 256.663
R902 B.n994 B.n125 256.663
R903 B.n994 B.n124 256.663
R904 B.n994 B.n123 256.663
R905 B.n994 B.n122 256.663
R906 B.n994 B.n121 256.663
R907 B.n994 B.n120 256.663
R908 B.n994 B.n119 256.663
R909 B.n994 B.n118 256.663
R910 B.n994 B.n117 256.663
R911 B.n994 B.n116 256.663
R912 B.n994 B.n115 256.663
R913 B.n994 B.n114 256.663
R914 B.n994 B.n113 256.663
R915 B.n994 B.n112 256.663
R916 B.n994 B.n111 256.663
R917 B.n535 B.n479 256.663
R918 B.n541 B.n479 256.663
R919 B.n543 B.n479 256.663
R920 B.n549 B.n479 256.663
R921 B.n551 B.n479 256.663
R922 B.n557 B.n479 256.663
R923 B.n559 B.n479 256.663
R924 B.n565 B.n479 256.663
R925 B.n567 B.n479 256.663
R926 B.n573 B.n479 256.663
R927 B.n575 B.n479 256.663
R928 B.n581 B.n479 256.663
R929 B.n583 B.n479 256.663
R930 B.n589 B.n479 256.663
R931 B.n591 B.n479 256.663
R932 B.n597 B.n479 256.663
R933 B.n599 B.n479 256.663
R934 B.n605 B.n479 256.663
R935 B.n607 B.n479 256.663
R936 B.n613 B.n479 256.663
R937 B.n615 B.n479 256.663
R938 B.n621 B.n479 256.663
R939 B.n623 B.n479 256.663
R940 B.n629 B.n479 256.663
R941 B.n631 B.n479 256.663
R942 B.n637 B.n479 256.663
R943 B.n639 B.n479 256.663
R944 B.n646 B.n479 256.663
R945 B.n648 B.n479 256.663
R946 B.n654 B.n479 256.663
R947 B.n656 B.n479 256.663
R948 B.n662 B.n479 256.663
R949 B.n664 B.n479 256.663
R950 B.n670 B.n479 256.663
R951 B.n672 B.n479 256.663
R952 B.n678 B.n479 256.663
R953 B.n680 B.n479 256.663
R954 B.n686 B.n479 256.663
R955 B.n688 B.n479 256.663
R956 B.n694 B.n479 256.663
R957 B.n696 B.n479 256.663
R958 B.n702 B.n479 256.663
R959 B.n704 B.n479 256.663
R960 B.n710 B.n479 256.663
R961 B.n712 B.n479 256.663
R962 B.n718 B.n479 256.663
R963 B.n720 B.n479 256.663
R964 B.n726 B.n479 256.663
R965 B.n729 B.n479 256.663
R966 B.n736 B.n476 163.367
R967 B.n740 B.n476 163.367
R968 B.n740 B.n470 163.367
R969 B.n748 B.n470 163.367
R970 B.n748 B.n468 163.367
R971 B.n752 B.n468 163.367
R972 B.n752 B.n462 163.367
R973 B.n760 B.n462 163.367
R974 B.n760 B.n460 163.367
R975 B.n764 B.n460 163.367
R976 B.n764 B.n454 163.367
R977 B.n772 B.n454 163.367
R978 B.n772 B.n452 163.367
R979 B.n776 B.n452 163.367
R980 B.n776 B.n446 163.367
R981 B.n784 B.n446 163.367
R982 B.n784 B.n444 163.367
R983 B.n788 B.n444 163.367
R984 B.n788 B.n438 163.367
R985 B.n796 B.n438 163.367
R986 B.n796 B.n436 163.367
R987 B.n800 B.n436 163.367
R988 B.n800 B.n430 163.367
R989 B.n808 B.n430 163.367
R990 B.n808 B.n428 163.367
R991 B.n812 B.n428 163.367
R992 B.n812 B.n422 163.367
R993 B.n820 B.n422 163.367
R994 B.n820 B.n420 163.367
R995 B.n824 B.n420 163.367
R996 B.n824 B.n414 163.367
R997 B.n832 B.n414 163.367
R998 B.n832 B.n412 163.367
R999 B.n836 B.n412 163.367
R1000 B.n836 B.n406 163.367
R1001 B.n844 B.n406 163.367
R1002 B.n844 B.n404 163.367
R1003 B.n848 B.n404 163.367
R1004 B.n848 B.n398 163.367
R1005 B.n856 B.n398 163.367
R1006 B.n856 B.n396 163.367
R1007 B.n860 B.n396 163.367
R1008 B.n860 B.n390 163.367
R1009 B.n868 B.n390 163.367
R1010 B.n868 B.n388 163.367
R1011 B.n872 B.n388 163.367
R1012 B.n872 B.n382 163.367
R1013 B.n880 B.n382 163.367
R1014 B.n880 B.n380 163.367
R1015 B.n884 B.n380 163.367
R1016 B.n884 B.n374 163.367
R1017 B.n893 B.n374 163.367
R1018 B.n893 B.n372 163.367
R1019 B.n897 B.n372 163.367
R1020 B.n897 B.n367 163.367
R1021 B.n906 B.n367 163.367
R1022 B.n906 B.n365 163.367
R1023 B.n910 B.n365 163.367
R1024 B.n910 B.n2 163.367
R1025 B.n1116 B.n2 163.367
R1026 B.n1116 B.n3 163.367
R1027 B.n1112 B.n3 163.367
R1028 B.n1112 B.n9 163.367
R1029 B.n1108 B.n9 163.367
R1030 B.n1108 B.n11 163.367
R1031 B.n1104 B.n11 163.367
R1032 B.n1104 B.n15 163.367
R1033 B.n1100 B.n15 163.367
R1034 B.n1100 B.n17 163.367
R1035 B.n1096 B.n17 163.367
R1036 B.n1096 B.n23 163.367
R1037 B.n1092 B.n23 163.367
R1038 B.n1092 B.n25 163.367
R1039 B.n1088 B.n25 163.367
R1040 B.n1088 B.n30 163.367
R1041 B.n1084 B.n30 163.367
R1042 B.n1084 B.n32 163.367
R1043 B.n1080 B.n32 163.367
R1044 B.n1080 B.n37 163.367
R1045 B.n1076 B.n37 163.367
R1046 B.n1076 B.n39 163.367
R1047 B.n1072 B.n39 163.367
R1048 B.n1072 B.n44 163.367
R1049 B.n1068 B.n44 163.367
R1050 B.n1068 B.n46 163.367
R1051 B.n1064 B.n46 163.367
R1052 B.n1064 B.n51 163.367
R1053 B.n1060 B.n51 163.367
R1054 B.n1060 B.n53 163.367
R1055 B.n1056 B.n53 163.367
R1056 B.n1056 B.n58 163.367
R1057 B.n1052 B.n58 163.367
R1058 B.n1052 B.n60 163.367
R1059 B.n1048 B.n60 163.367
R1060 B.n1048 B.n65 163.367
R1061 B.n1044 B.n65 163.367
R1062 B.n1044 B.n67 163.367
R1063 B.n1040 B.n67 163.367
R1064 B.n1040 B.n72 163.367
R1065 B.n1036 B.n72 163.367
R1066 B.n1036 B.n74 163.367
R1067 B.n1032 B.n74 163.367
R1068 B.n1032 B.n79 163.367
R1069 B.n1028 B.n79 163.367
R1070 B.n1028 B.n81 163.367
R1071 B.n1024 B.n81 163.367
R1072 B.n1024 B.n86 163.367
R1073 B.n1020 B.n86 163.367
R1074 B.n1020 B.n88 163.367
R1075 B.n1016 B.n88 163.367
R1076 B.n1016 B.n93 163.367
R1077 B.n1012 B.n93 163.367
R1078 B.n1012 B.n95 163.367
R1079 B.n1008 B.n95 163.367
R1080 B.n1008 B.n100 163.367
R1081 B.n1004 B.n100 163.367
R1082 B.n1004 B.n102 163.367
R1083 B.n1000 B.n102 163.367
R1084 B.n1000 B.n107 163.367
R1085 B.n996 B.n107 163.367
R1086 B.n536 B.n534 163.367
R1087 B.n540 B.n534 163.367
R1088 B.n544 B.n542 163.367
R1089 B.n548 B.n532 163.367
R1090 B.n552 B.n550 163.367
R1091 B.n556 B.n530 163.367
R1092 B.n560 B.n558 163.367
R1093 B.n564 B.n528 163.367
R1094 B.n568 B.n566 163.367
R1095 B.n572 B.n526 163.367
R1096 B.n576 B.n574 163.367
R1097 B.n580 B.n524 163.367
R1098 B.n584 B.n582 163.367
R1099 B.n588 B.n522 163.367
R1100 B.n592 B.n590 163.367
R1101 B.n596 B.n520 163.367
R1102 B.n600 B.n598 163.367
R1103 B.n604 B.n518 163.367
R1104 B.n608 B.n606 163.367
R1105 B.n612 B.n516 163.367
R1106 B.n616 B.n614 163.367
R1107 B.n620 B.n514 163.367
R1108 B.n624 B.n622 163.367
R1109 B.n628 B.n509 163.367
R1110 B.n632 B.n630 163.367
R1111 B.n636 B.n507 163.367
R1112 B.n640 B.n638 163.367
R1113 B.n645 B.n503 163.367
R1114 B.n649 B.n647 163.367
R1115 B.n653 B.n501 163.367
R1116 B.n657 B.n655 163.367
R1117 B.n661 B.n499 163.367
R1118 B.n665 B.n663 163.367
R1119 B.n669 B.n497 163.367
R1120 B.n673 B.n671 163.367
R1121 B.n677 B.n495 163.367
R1122 B.n681 B.n679 163.367
R1123 B.n685 B.n493 163.367
R1124 B.n689 B.n687 163.367
R1125 B.n693 B.n491 163.367
R1126 B.n697 B.n695 163.367
R1127 B.n701 B.n489 163.367
R1128 B.n705 B.n703 163.367
R1129 B.n709 B.n487 163.367
R1130 B.n713 B.n711 163.367
R1131 B.n717 B.n485 163.367
R1132 B.n721 B.n719 163.367
R1133 B.n725 B.n483 163.367
R1134 B.n728 B.n727 163.367
R1135 B.n730 B.n480 163.367
R1136 B.n734 B.n474 163.367
R1137 B.n742 B.n474 163.367
R1138 B.n742 B.n472 163.367
R1139 B.n746 B.n472 163.367
R1140 B.n746 B.n466 163.367
R1141 B.n754 B.n466 163.367
R1142 B.n754 B.n464 163.367
R1143 B.n758 B.n464 163.367
R1144 B.n758 B.n458 163.367
R1145 B.n766 B.n458 163.367
R1146 B.n766 B.n456 163.367
R1147 B.n770 B.n456 163.367
R1148 B.n770 B.n450 163.367
R1149 B.n778 B.n450 163.367
R1150 B.n778 B.n448 163.367
R1151 B.n782 B.n448 163.367
R1152 B.n782 B.n442 163.367
R1153 B.n790 B.n442 163.367
R1154 B.n790 B.n440 163.367
R1155 B.n794 B.n440 163.367
R1156 B.n794 B.n434 163.367
R1157 B.n802 B.n434 163.367
R1158 B.n802 B.n432 163.367
R1159 B.n806 B.n432 163.367
R1160 B.n806 B.n426 163.367
R1161 B.n814 B.n426 163.367
R1162 B.n814 B.n424 163.367
R1163 B.n818 B.n424 163.367
R1164 B.n818 B.n418 163.367
R1165 B.n826 B.n418 163.367
R1166 B.n826 B.n416 163.367
R1167 B.n830 B.n416 163.367
R1168 B.n830 B.n410 163.367
R1169 B.n838 B.n410 163.367
R1170 B.n838 B.n408 163.367
R1171 B.n842 B.n408 163.367
R1172 B.n842 B.n402 163.367
R1173 B.n850 B.n402 163.367
R1174 B.n850 B.n400 163.367
R1175 B.n854 B.n400 163.367
R1176 B.n854 B.n394 163.367
R1177 B.n862 B.n394 163.367
R1178 B.n862 B.n392 163.367
R1179 B.n866 B.n392 163.367
R1180 B.n866 B.n386 163.367
R1181 B.n874 B.n386 163.367
R1182 B.n874 B.n384 163.367
R1183 B.n878 B.n384 163.367
R1184 B.n878 B.n378 163.367
R1185 B.n886 B.n378 163.367
R1186 B.n886 B.n376 163.367
R1187 B.n890 B.n376 163.367
R1188 B.n890 B.n371 163.367
R1189 B.n899 B.n371 163.367
R1190 B.n899 B.n369 163.367
R1191 B.n904 B.n369 163.367
R1192 B.n904 B.n363 163.367
R1193 B.n912 B.n363 163.367
R1194 B.n913 B.n912 163.367
R1195 B.n913 B.n5 163.367
R1196 B.n6 B.n5 163.367
R1197 B.n7 B.n6 163.367
R1198 B.n918 B.n7 163.367
R1199 B.n918 B.n12 163.367
R1200 B.n13 B.n12 163.367
R1201 B.n14 B.n13 163.367
R1202 B.n923 B.n14 163.367
R1203 B.n923 B.n19 163.367
R1204 B.n20 B.n19 163.367
R1205 B.n21 B.n20 163.367
R1206 B.n928 B.n21 163.367
R1207 B.n928 B.n26 163.367
R1208 B.n27 B.n26 163.367
R1209 B.n28 B.n27 163.367
R1210 B.n933 B.n28 163.367
R1211 B.n933 B.n33 163.367
R1212 B.n34 B.n33 163.367
R1213 B.n35 B.n34 163.367
R1214 B.n938 B.n35 163.367
R1215 B.n938 B.n40 163.367
R1216 B.n41 B.n40 163.367
R1217 B.n42 B.n41 163.367
R1218 B.n943 B.n42 163.367
R1219 B.n943 B.n47 163.367
R1220 B.n48 B.n47 163.367
R1221 B.n49 B.n48 163.367
R1222 B.n948 B.n49 163.367
R1223 B.n948 B.n54 163.367
R1224 B.n55 B.n54 163.367
R1225 B.n56 B.n55 163.367
R1226 B.n953 B.n56 163.367
R1227 B.n953 B.n61 163.367
R1228 B.n62 B.n61 163.367
R1229 B.n63 B.n62 163.367
R1230 B.n958 B.n63 163.367
R1231 B.n958 B.n68 163.367
R1232 B.n69 B.n68 163.367
R1233 B.n70 B.n69 163.367
R1234 B.n963 B.n70 163.367
R1235 B.n963 B.n75 163.367
R1236 B.n76 B.n75 163.367
R1237 B.n77 B.n76 163.367
R1238 B.n968 B.n77 163.367
R1239 B.n968 B.n82 163.367
R1240 B.n83 B.n82 163.367
R1241 B.n84 B.n83 163.367
R1242 B.n973 B.n84 163.367
R1243 B.n973 B.n89 163.367
R1244 B.n90 B.n89 163.367
R1245 B.n91 B.n90 163.367
R1246 B.n978 B.n91 163.367
R1247 B.n978 B.n96 163.367
R1248 B.n97 B.n96 163.367
R1249 B.n98 B.n97 163.367
R1250 B.n983 B.n98 163.367
R1251 B.n983 B.n103 163.367
R1252 B.n104 B.n103 163.367
R1253 B.n105 B.n104 163.367
R1254 B.n988 B.n105 163.367
R1255 B.n988 B.n110 163.367
R1256 B.n167 B.n166 163.367
R1257 B.n171 B.n170 163.367
R1258 B.n175 B.n174 163.367
R1259 B.n179 B.n178 163.367
R1260 B.n183 B.n182 163.367
R1261 B.n187 B.n186 163.367
R1262 B.n191 B.n190 163.367
R1263 B.n195 B.n194 163.367
R1264 B.n199 B.n198 163.367
R1265 B.n203 B.n202 163.367
R1266 B.n207 B.n206 163.367
R1267 B.n211 B.n210 163.367
R1268 B.n215 B.n214 163.367
R1269 B.n219 B.n218 163.367
R1270 B.n223 B.n222 163.367
R1271 B.n227 B.n226 163.367
R1272 B.n231 B.n230 163.367
R1273 B.n235 B.n234 163.367
R1274 B.n239 B.n238 163.367
R1275 B.n243 B.n242 163.367
R1276 B.n247 B.n246 163.367
R1277 B.n251 B.n250 163.367
R1278 B.n256 B.n255 163.367
R1279 B.n260 B.n259 163.367
R1280 B.n264 B.n263 163.367
R1281 B.n268 B.n267 163.367
R1282 B.n272 B.n271 163.367
R1283 B.n277 B.n276 163.367
R1284 B.n281 B.n280 163.367
R1285 B.n285 B.n284 163.367
R1286 B.n289 B.n288 163.367
R1287 B.n293 B.n292 163.367
R1288 B.n297 B.n296 163.367
R1289 B.n301 B.n300 163.367
R1290 B.n305 B.n304 163.367
R1291 B.n309 B.n308 163.367
R1292 B.n313 B.n312 163.367
R1293 B.n317 B.n316 163.367
R1294 B.n321 B.n320 163.367
R1295 B.n325 B.n324 163.367
R1296 B.n329 B.n328 163.367
R1297 B.n333 B.n332 163.367
R1298 B.n337 B.n336 163.367
R1299 B.n341 B.n340 163.367
R1300 B.n345 B.n344 163.367
R1301 B.n349 B.n348 163.367
R1302 B.n353 B.n352 163.367
R1303 B.n357 B.n356 163.367
R1304 B.n359 B.n160 163.367
R1305 B.n504 B.t21 141.917
R1306 B.n161 B.t10 141.917
R1307 B.n510 B.t18 141.9
R1308 B.n163 B.t13 141.9
R1309 B.n505 B.t20 73.6501
R1310 B.n162 B.t11 73.6501
R1311 B.n511 B.t17 73.6334
R1312 B.n164 B.t14 73.6334
R1313 B.n535 B.n478 71.676
R1314 B.n541 B.n540 71.676
R1315 B.n544 B.n543 71.676
R1316 B.n549 B.n548 71.676
R1317 B.n552 B.n551 71.676
R1318 B.n557 B.n556 71.676
R1319 B.n560 B.n559 71.676
R1320 B.n565 B.n564 71.676
R1321 B.n568 B.n567 71.676
R1322 B.n573 B.n572 71.676
R1323 B.n576 B.n575 71.676
R1324 B.n581 B.n580 71.676
R1325 B.n584 B.n583 71.676
R1326 B.n589 B.n588 71.676
R1327 B.n592 B.n591 71.676
R1328 B.n597 B.n596 71.676
R1329 B.n600 B.n599 71.676
R1330 B.n605 B.n604 71.676
R1331 B.n608 B.n607 71.676
R1332 B.n613 B.n612 71.676
R1333 B.n616 B.n615 71.676
R1334 B.n621 B.n620 71.676
R1335 B.n624 B.n623 71.676
R1336 B.n629 B.n628 71.676
R1337 B.n632 B.n631 71.676
R1338 B.n637 B.n636 71.676
R1339 B.n640 B.n639 71.676
R1340 B.n646 B.n645 71.676
R1341 B.n649 B.n648 71.676
R1342 B.n654 B.n653 71.676
R1343 B.n657 B.n656 71.676
R1344 B.n662 B.n661 71.676
R1345 B.n665 B.n664 71.676
R1346 B.n670 B.n669 71.676
R1347 B.n673 B.n672 71.676
R1348 B.n678 B.n677 71.676
R1349 B.n681 B.n680 71.676
R1350 B.n686 B.n685 71.676
R1351 B.n689 B.n688 71.676
R1352 B.n694 B.n693 71.676
R1353 B.n697 B.n696 71.676
R1354 B.n702 B.n701 71.676
R1355 B.n705 B.n704 71.676
R1356 B.n710 B.n709 71.676
R1357 B.n713 B.n712 71.676
R1358 B.n718 B.n717 71.676
R1359 B.n721 B.n720 71.676
R1360 B.n726 B.n725 71.676
R1361 B.n729 B.n728 71.676
R1362 B.n111 B.n109 71.676
R1363 B.n167 B.n112 71.676
R1364 B.n171 B.n113 71.676
R1365 B.n175 B.n114 71.676
R1366 B.n179 B.n115 71.676
R1367 B.n183 B.n116 71.676
R1368 B.n187 B.n117 71.676
R1369 B.n191 B.n118 71.676
R1370 B.n195 B.n119 71.676
R1371 B.n199 B.n120 71.676
R1372 B.n203 B.n121 71.676
R1373 B.n207 B.n122 71.676
R1374 B.n211 B.n123 71.676
R1375 B.n215 B.n124 71.676
R1376 B.n219 B.n125 71.676
R1377 B.n223 B.n126 71.676
R1378 B.n227 B.n127 71.676
R1379 B.n231 B.n128 71.676
R1380 B.n235 B.n129 71.676
R1381 B.n239 B.n130 71.676
R1382 B.n243 B.n131 71.676
R1383 B.n247 B.n132 71.676
R1384 B.n251 B.n133 71.676
R1385 B.n256 B.n134 71.676
R1386 B.n260 B.n135 71.676
R1387 B.n264 B.n136 71.676
R1388 B.n268 B.n137 71.676
R1389 B.n272 B.n138 71.676
R1390 B.n277 B.n139 71.676
R1391 B.n281 B.n140 71.676
R1392 B.n285 B.n141 71.676
R1393 B.n289 B.n142 71.676
R1394 B.n293 B.n143 71.676
R1395 B.n297 B.n144 71.676
R1396 B.n301 B.n145 71.676
R1397 B.n305 B.n146 71.676
R1398 B.n309 B.n147 71.676
R1399 B.n313 B.n148 71.676
R1400 B.n317 B.n149 71.676
R1401 B.n321 B.n150 71.676
R1402 B.n325 B.n151 71.676
R1403 B.n329 B.n152 71.676
R1404 B.n333 B.n153 71.676
R1405 B.n337 B.n154 71.676
R1406 B.n341 B.n155 71.676
R1407 B.n345 B.n156 71.676
R1408 B.n349 B.n157 71.676
R1409 B.n353 B.n158 71.676
R1410 B.n357 B.n159 71.676
R1411 B.n993 B.n160 71.676
R1412 B.n993 B.n992 71.676
R1413 B.n359 B.n159 71.676
R1414 B.n356 B.n158 71.676
R1415 B.n352 B.n157 71.676
R1416 B.n348 B.n156 71.676
R1417 B.n344 B.n155 71.676
R1418 B.n340 B.n154 71.676
R1419 B.n336 B.n153 71.676
R1420 B.n332 B.n152 71.676
R1421 B.n328 B.n151 71.676
R1422 B.n324 B.n150 71.676
R1423 B.n320 B.n149 71.676
R1424 B.n316 B.n148 71.676
R1425 B.n312 B.n147 71.676
R1426 B.n308 B.n146 71.676
R1427 B.n304 B.n145 71.676
R1428 B.n300 B.n144 71.676
R1429 B.n296 B.n143 71.676
R1430 B.n292 B.n142 71.676
R1431 B.n288 B.n141 71.676
R1432 B.n284 B.n140 71.676
R1433 B.n280 B.n139 71.676
R1434 B.n276 B.n138 71.676
R1435 B.n271 B.n137 71.676
R1436 B.n267 B.n136 71.676
R1437 B.n263 B.n135 71.676
R1438 B.n259 B.n134 71.676
R1439 B.n255 B.n133 71.676
R1440 B.n250 B.n132 71.676
R1441 B.n246 B.n131 71.676
R1442 B.n242 B.n130 71.676
R1443 B.n238 B.n129 71.676
R1444 B.n234 B.n128 71.676
R1445 B.n230 B.n127 71.676
R1446 B.n226 B.n126 71.676
R1447 B.n222 B.n125 71.676
R1448 B.n218 B.n124 71.676
R1449 B.n214 B.n123 71.676
R1450 B.n210 B.n122 71.676
R1451 B.n206 B.n121 71.676
R1452 B.n202 B.n120 71.676
R1453 B.n198 B.n119 71.676
R1454 B.n194 B.n118 71.676
R1455 B.n190 B.n117 71.676
R1456 B.n186 B.n116 71.676
R1457 B.n182 B.n115 71.676
R1458 B.n178 B.n114 71.676
R1459 B.n174 B.n113 71.676
R1460 B.n170 B.n112 71.676
R1461 B.n166 B.n111 71.676
R1462 B.n536 B.n535 71.676
R1463 B.n542 B.n541 71.676
R1464 B.n543 B.n532 71.676
R1465 B.n550 B.n549 71.676
R1466 B.n551 B.n530 71.676
R1467 B.n558 B.n557 71.676
R1468 B.n559 B.n528 71.676
R1469 B.n566 B.n565 71.676
R1470 B.n567 B.n526 71.676
R1471 B.n574 B.n573 71.676
R1472 B.n575 B.n524 71.676
R1473 B.n582 B.n581 71.676
R1474 B.n583 B.n522 71.676
R1475 B.n590 B.n589 71.676
R1476 B.n591 B.n520 71.676
R1477 B.n598 B.n597 71.676
R1478 B.n599 B.n518 71.676
R1479 B.n606 B.n605 71.676
R1480 B.n607 B.n516 71.676
R1481 B.n614 B.n613 71.676
R1482 B.n615 B.n514 71.676
R1483 B.n622 B.n621 71.676
R1484 B.n623 B.n509 71.676
R1485 B.n630 B.n629 71.676
R1486 B.n631 B.n507 71.676
R1487 B.n638 B.n637 71.676
R1488 B.n639 B.n503 71.676
R1489 B.n647 B.n646 71.676
R1490 B.n648 B.n501 71.676
R1491 B.n655 B.n654 71.676
R1492 B.n656 B.n499 71.676
R1493 B.n663 B.n662 71.676
R1494 B.n664 B.n497 71.676
R1495 B.n671 B.n670 71.676
R1496 B.n672 B.n495 71.676
R1497 B.n679 B.n678 71.676
R1498 B.n680 B.n493 71.676
R1499 B.n687 B.n686 71.676
R1500 B.n688 B.n491 71.676
R1501 B.n695 B.n694 71.676
R1502 B.n696 B.n489 71.676
R1503 B.n703 B.n702 71.676
R1504 B.n704 B.n487 71.676
R1505 B.n711 B.n710 71.676
R1506 B.n712 B.n485 71.676
R1507 B.n719 B.n718 71.676
R1508 B.n720 B.n483 71.676
R1509 B.n727 B.n726 71.676
R1510 B.n730 B.n729 71.676
R1511 B.n735 B.n479 68.3604
R1512 B.n995 B.n994 68.3604
R1513 B.n505 B.n504 68.2672
R1514 B.n511 B.n510 68.2672
R1515 B.n164 B.n163 68.2672
R1516 B.n162 B.n161 68.2672
R1517 B.n643 B.n505 59.5399
R1518 B.n512 B.n511 59.5399
R1519 B.n253 B.n164 59.5399
R1520 B.n274 B.n162 59.5399
R1521 B.n735 B.n475 40.422
R1522 B.n741 B.n475 40.422
R1523 B.n741 B.n471 40.422
R1524 B.n747 B.n471 40.422
R1525 B.n747 B.n467 40.422
R1526 B.n753 B.n467 40.422
R1527 B.n753 B.n463 40.422
R1528 B.n759 B.n463 40.422
R1529 B.n765 B.n459 40.422
R1530 B.n765 B.n455 40.422
R1531 B.n771 B.n455 40.422
R1532 B.n771 B.n451 40.422
R1533 B.n777 B.n451 40.422
R1534 B.n777 B.n447 40.422
R1535 B.n783 B.n447 40.422
R1536 B.n783 B.n443 40.422
R1537 B.n789 B.n443 40.422
R1538 B.n789 B.n439 40.422
R1539 B.n795 B.n439 40.422
R1540 B.n795 B.n435 40.422
R1541 B.n801 B.n435 40.422
R1542 B.n807 B.n431 40.422
R1543 B.n807 B.n427 40.422
R1544 B.n813 B.n427 40.422
R1545 B.n813 B.n423 40.422
R1546 B.n819 B.n423 40.422
R1547 B.n819 B.n419 40.422
R1548 B.n825 B.n419 40.422
R1549 B.n825 B.n415 40.422
R1550 B.n831 B.n415 40.422
R1551 B.n837 B.n411 40.422
R1552 B.n837 B.n407 40.422
R1553 B.n843 B.n407 40.422
R1554 B.n843 B.n403 40.422
R1555 B.n849 B.n403 40.422
R1556 B.n849 B.n399 40.422
R1557 B.n855 B.n399 40.422
R1558 B.n855 B.n395 40.422
R1559 B.n861 B.n395 40.422
R1560 B.n867 B.n391 40.422
R1561 B.n867 B.n387 40.422
R1562 B.n873 B.n387 40.422
R1563 B.n873 B.n383 40.422
R1564 B.n879 B.n383 40.422
R1565 B.n879 B.n379 40.422
R1566 B.n885 B.n379 40.422
R1567 B.n885 B.n375 40.422
R1568 B.n892 B.n375 40.422
R1569 B.n892 B.n891 40.422
R1570 B.n898 B.n368 40.422
R1571 B.n905 B.n368 40.422
R1572 B.n905 B.n364 40.422
R1573 B.n911 B.n364 40.422
R1574 B.n911 B.n4 40.422
R1575 B.n1115 B.n4 40.422
R1576 B.n1115 B.n1114 40.422
R1577 B.n1114 B.n1113 40.422
R1578 B.n1113 B.n8 40.422
R1579 B.n1107 B.n8 40.422
R1580 B.n1107 B.n1106 40.422
R1581 B.n1106 B.n1105 40.422
R1582 B.n1099 B.n18 40.422
R1583 B.n1099 B.n1098 40.422
R1584 B.n1098 B.n1097 40.422
R1585 B.n1097 B.n22 40.422
R1586 B.n1091 B.n22 40.422
R1587 B.n1091 B.n1090 40.422
R1588 B.n1090 B.n1089 40.422
R1589 B.n1089 B.n29 40.422
R1590 B.n1083 B.n29 40.422
R1591 B.n1083 B.n1082 40.422
R1592 B.n1081 B.n36 40.422
R1593 B.n1075 B.n36 40.422
R1594 B.n1075 B.n1074 40.422
R1595 B.n1074 B.n1073 40.422
R1596 B.n1073 B.n43 40.422
R1597 B.n1067 B.n43 40.422
R1598 B.n1067 B.n1066 40.422
R1599 B.n1066 B.n1065 40.422
R1600 B.n1065 B.n50 40.422
R1601 B.n1059 B.n1058 40.422
R1602 B.n1058 B.n1057 40.422
R1603 B.n1057 B.n57 40.422
R1604 B.n1051 B.n57 40.422
R1605 B.n1051 B.n1050 40.422
R1606 B.n1050 B.n1049 40.422
R1607 B.n1049 B.n64 40.422
R1608 B.n1043 B.n64 40.422
R1609 B.n1043 B.n1042 40.422
R1610 B.n1041 B.n71 40.422
R1611 B.n1035 B.n71 40.422
R1612 B.n1035 B.n1034 40.422
R1613 B.n1034 B.n1033 40.422
R1614 B.n1033 B.n78 40.422
R1615 B.n1027 B.n78 40.422
R1616 B.n1027 B.n1026 40.422
R1617 B.n1026 B.n1025 40.422
R1618 B.n1025 B.n85 40.422
R1619 B.n1019 B.n85 40.422
R1620 B.n1019 B.n1018 40.422
R1621 B.n1018 B.n1017 40.422
R1622 B.n1017 B.n92 40.422
R1623 B.n1011 B.n1010 40.422
R1624 B.n1010 B.n1009 40.422
R1625 B.n1009 B.n99 40.422
R1626 B.n1003 B.n99 40.422
R1627 B.n1003 B.n1002 40.422
R1628 B.n1002 B.n1001 40.422
R1629 B.n1001 B.n106 40.422
R1630 B.n995 B.n106 40.422
R1631 B.n861 B.t6 35.0721
R1632 B.t4 B.n1081 35.0721
R1633 B.t7 B.n431 33.8832
R1634 B.n1042 B.t3 33.8832
R1635 B.n898 B.t5 31.5055
R1636 B.n1105 B.t0 31.5055
R1637 B.n997 B.n108 31.3761
R1638 B.n991 B.n990 31.3761
R1639 B.n733 B.n732 31.3761
R1640 B.n737 B.n477 31.3761
R1641 B.n759 B.t16 24.3723
R1642 B.n1011 B.t9 24.3723
R1643 B.n831 B.t2 20.8057
R1644 B.n1059 B.t1 20.8057
R1645 B.t2 B.n411 19.6168
R1646 B.t1 B.n50 19.6168
R1647 B B.n1117 18.0485
R1648 B.t16 B.n459 16.0502
R1649 B.t9 B.n92 16.0502
R1650 B.n165 B.n108 10.6151
R1651 B.n168 B.n165 10.6151
R1652 B.n169 B.n168 10.6151
R1653 B.n172 B.n169 10.6151
R1654 B.n173 B.n172 10.6151
R1655 B.n176 B.n173 10.6151
R1656 B.n177 B.n176 10.6151
R1657 B.n180 B.n177 10.6151
R1658 B.n181 B.n180 10.6151
R1659 B.n184 B.n181 10.6151
R1660 B.n185 B.n184 10.6151
R1661 B.n188 B.n185 10.6151
R1662 B.n189 B.n188 10.6151
R1663 B.n192 B.n189 10.6151
R1664 B.n193 B.n192 10.6151
R1665 B.n196 B.n193 10.6151
R1666 B.n197 B.n196 10.6151
R1667 B.n200 B.n197 10.6151
R1668 B.n201 B.n200 10.6151
R1669 B.n204 B.n201 10.6151
R1670 B.n205 B.n204 10.6151
R1671 B.n208 B.n205 10.6151
R1672 B.n209 B.n208 10.6151
R1673 B.n212 B.n209 10.6151
R1674 B.n213 B.n212 10.6151
R1675 B.n216 B.n213 10.6151
R1676 B.n217 B.n216 10.6151
R1677 B.n220 B.n217 10.6151
R1678 B.n221 B.n220 10.6151
R1679 B.n224 B.n221 10.6151
R1680 B.n225 B.n224 10.6151
R1681 B.n228 B.n225 10.6151
R1682 B.n229 B.n228 10.6151
R1683 B.n232 B.n229 10.6151
R1684 B.n233 B.n232 10.6151
R1685 B.n236 B.n233 10.6151
R1686 B.n237 B.n236 10.6151
R1687 B.n240 B.n237 10.6151
R1688 B.n241 B.n240 10.6151
R1689 B.n244 B.n241 10.6151
R1690 B.n245 B.n244 10.6151
R1691 B.n248 B.n245 10.6151
R1692 B.n249 B.n248 10.6151
R1693 B.n252 B.n249 10.6151
R1694 B.n257 B.n254 10.6151
R1695 B.n258 B.n257 10.6151
R1696 B.n261 B.n258 10.6151
R1697 B.n262 B.n261 10.6151
R1698 B.n265 B.n262 10.6151
R1699 B.n266 B.n265 10.6151
R1700 B.n269 B.n266 10.6151
R1701 B.n270 B.n269 10.6151
R1702 B.n273 B.n270 10.6151
R1703 B.n278 B.n275 10.6151
R1704 B.n279 B.n278 10.6151
R1705 B.n282 B.n279 10.6151
R1706 B.n283 B.n282 10.6151
R1707 B.n286 B.n283 10.6151
R1708 B.n287 B.n286 10.6151
R1709 B.n290 B.n287 10.6151
R1710 B.n291 B.n290 10.6151
R1711 B.n294 B.n291 10.6151
R1712 B.n295 B.n294 10.6151
R1713 B.n298 B.n295 10.6151
R1714 B.n299 B.n298 10.6151
R1715 B.n302 B.n299 10.6151
R1716 B.n303 B.n302 10.6151
R1717 B.n306 B.n303 10.6151
R1718 B.n307 B.n306 10.6151
R1719 B.n310 B.n307 10.6151
R1720 B.n311 B.n310 10.6151
R1721 B.n314 B.n311 10.6151
R1722 B.n315 B.n314 10.6151
R1723 B.n318 B.n315 10.6151
R1724 B.n319 B.n318 10.6151
R1725 B.n322 B.n319 10.6151
R1726 B.n323 B.n322 10.6151
R1727 B.n326 B.n323 10.6151
R1728 B.n327 B.n326 10.6151
R1729 B.n330 B.n327 10.6151
R1730 B.n331 B.n330 10.6151
R1731 B.n334 B.n331 10.6151
R1732 B.n335 B.n334 10.6151
R1733 B.n338 B.n335 10.6151
R1734 B.n339 B.n338 10.6151
R1735 B.n342 B.n339 10.6151
R1736 B.n343 B.n342 10.6151
R1737 B.n346 B.n343 10.6151
R1738 B.n347 B.n346 10.6151
R1739 B.n350 B.n347 10.6151
R1740 B.n351 B.n350 10.6151
R1741 B.n354 B.n351 10.6151
R1742 B.n355 B.n354 10.6151
R1743 B.n358 B.n355 10.6151
R1744 B.n360 B.n358 10.6151
R1745 B.n361 B.n360 10.6151
R1746 B.n991 B.n361 10.6151
R1747 B.n733 B.n473 10.6151
R1748 B.n743 B.n473 10.6151
R1749 B.n744 B.n743 10.6151
R1750 B.n745 B.n744 10.6151
R1751 B.n745 B.n465 10.6151
R1752 B.n755 B.n465 10.6151
R1753 B.n756 B.n755 10.6151
R1754 B.n757 B.n756 10.6151
R1755 B.n757 B.n457 10.6151
R1756 B.n767 B.n457 10.6151
R1757 B.n768 B.n767 10.6151
R1758 B.n769 B.n768 10.6151
R1759 B.n769 B.n449 10.6151
R1760 B.n779 B.n449 10.6151
R1761 B.n780 B.n779 10.6151
R1762 B.n781 B.n780 10.6151
R1763 B.n781 B.n441 10.6151
R1764 B.n791 B.n441 10.6151
R1765 B.n792 B.n791 10.6151
R1766 B.n793 B.n792 10.6151
R1767 B.n793 B.n433 10.6151
R1768 B.n803 B.n433 10.6151
R1769 B.n804 B.n803 10.6151
R1770 B.n805 B.n804 10.6151
R1771 B.n805 B.n425 10.6151
R1772 B.n815 B.n425 10.6151
R1773 B.n816 B.n815 10.6151
R1774 B.n817 B.n816 10.6151
R1775 B.n817 B.n417 10.6151
R1776 B.n827 B.n417 10.6151
R1777 B.n828 B.n827 10.6151
R1778 B.n829 B.n828 10.6151
R1779 B.n829 B.n409 10.6151
R1780 B.n839 B.n409 10.6151
R1781 B.n840 B.n839 10.6151
R1782 B.n841 B.n840 10.6151
R1783 B.n841 B.n401 10.6151
R1784 B.n851 B.n401 10.6151
R1785 B.n852 B.n851 10.6151
R1786 B.n853 B.n852 10.6151
R1787 B.n853 B.n393 10.6151
R1788 B.n863 B.n393 10.6151
R1789 B.n864 B.n863 10.6151
R1790 B.n865 B.n864 10.6151
R1791 B.n865 B.n385 10.6151
R1792 B.n875 B.n385 10.6151
R1793 B.n876 B.n875 10.6151
R1794 B.n877 B.n876 10.6151
R1795 B.n877 B.n377 10.6151
R1796 B.n887 B.n377 10.6151
R1797 B.n888 B.n887 10.6151
R1798 B.n889 B.n888 10.6151
R1799 B.n889 B.n370 10.6151
R1800 B.n900 B.n370 10.6151
R1801 B.n901 B.n900 10.6151
R1802 B.n903 B.n901 10.6151
R1803 B.n903 B.n902 10.6151
R1804 B.n902 B.n362 10.6151
R1805 B.n914 B.n362 10.6151
R1806 B.n915 B.n914 10.6151
R1807 B.n916 B.n915 10.6151
R1808 B.n917 B.n916 10.6151
R1809 B.n919 B.n917 10.6151
R1810 B.n920 B.n919 10.6151
R1811 B.n921 B.n920 10.6151
R1812 B.n922 B.n921 10.6151
R1813 B.n924 B.n922 10.6151
R1814 B.n925 B.n924 10.6151
R1815 B.n926 B.n925 10.6151
R1816 B.n927 B.n926 10.6151
R1817 B.n929 B.n927 10.6151
R1818 B.n930 B.n929 10.6151
R1819 B.n931 B.n930 10.6151
R1820 B.n932 B.n931 10.6151
R1821 B.n934 B.n932 10.6151
R1822 B.n935 B.n934 10.6151
R1823 B.n936 B.n935 10.6151
R1824 B.n937 B.n936 10.6151
R1825 B.n939 B.n937 10.6151
R1826 B.n940 B.n939 10.6151
R1827 B.n941 B.n940 10.6151
R1828 B.n942 B.n941 10.6151
R1829 B.n944 B.n942 10.6151
R1830 B.n945 B.n944 10.6151
R1831 B.n946 B.n945 10.6151
R1832 B.n947 B.n946 10.6151
R1833 B.n949 B.n947 10.6151
R1834 B.n950 B.n949 10.6151
R1835 B.n951 B.n950 10.6151
R1836 B.n952 B.n951 10.6151
R1837 B.n954 B.n952 10.6151
R1838 B.n955 B.n954 10.6151
R1839 B.n956 B.n955 10.6151
R1840 B.n957 B.n956 10.6151
R1841 B.n959 B.n957 10.6151
R1842 B.n960 B.n959 10.6151
R1843 B.n961 B.n960 10.6151
R1844 B.n962 B.n961 10.6151
R1845 B.n964 B.n962 10.6151
R1846 B.n965 B.n964 10.6151
R1847 B.n966 B.n965 10.6151
R1848 B.n967 B.n966 10.6151
R1849 B.n969 B.n967 10.6151
R1850 B.n970 B.n969 10.6151
R1851 B.n971 B.n970 10.6151
R1852 B.n972 B.n971 10.6151
R1853 B.n974 B.n972 10.6151
R1854 B.n975 B.n974 10.6151
R1855 B.n976 B.n975 10.6151
R1856 B.n977 B.n976 10.6151
R1857 B.n979 B.n977 10.6151
R1858 B.n980 B.n979 10.6151
R1859 B.n981 B.n980 10.6151
R1860 B.n982 B.n981 10.6151
R1861 B.n984 B.n982 10.6151
R1862 B.n985 B.n984 10.6151
R1863 B.n986 B.n985 10.6151
R1864 B.n987 B.n986 10.6151
R1865 B.n989 B.n987 10.6151
R1866 B.n990 B.n989 10.6151
R1867 B.n537 B.n477 10.6151
R1868 B.n538 B.n537 10.6151
R1869 B.n539 B.n538 10.6151
R1870 B.n539 B.n533 10.6151
R1871 B.n545 B.n533 10.6151
R1872 B.n546 B.n545 10.6151
R1873 B.n547 B.n546 10.6151
R1874 B.n547 B.n531 10.6151
R1875 B.n553 B.n531 10.6151
R1876 B.n554 B.n553 10.6151
R1877 B.n555 B.n554 10.6151
R1878 B.n555 B.n529 10.6151
R1879 B.n561 B.n529 10.6151
R1880 B.n562 B.n561 10.6151
R1881 B.n563 B.n562 10.6151
R1882 B.n563 B.n527 10.6151
R1883 B.n569 B.n527 10.6151
R1884 B.n570 B.n569 10.6151
R1885 B.n571 B.n570 10.6151
R1886 B.n571 B.n525 10.6151
R1887 B.n577 B.n525 10.6151
R1888 B.n578 B.n577 10.6151
R1889 B.n579 B.n578 10.6151
R1890 B.n579 B.n523 10.6151
R1891 B.n585 B.n523 10.6151
R1892 B.n586 B.n585 10.6151
R1893 B.n587 B.n586 10.6151
R1894 B.n587 B.n521 10.6151
R1895 B.n593 B.n521 10.6151
R1896 B.n594 B.n593 10.6151
R1897 B.n595 B.n594 10.6151
R1898 B.n595 B.n519 10.6151
R1899 B.n601 B.n519 10.6151
R1900 B.n602 B.n601 10.6151
R1901 B.n603 B.n602 10.6151
R1902 B.n603 B.n517 10.6151
R1903 B.n609 B.n517 10.6151
R1904 B.n610 B.n609 10.6151
R1905 B.n611 B.n610 10.6151
R1906 B.n611 B.n515 10.6151
R1907 B.n617 B.n515 10.6151
R1908 B.n618 B.n617 10.6151
R1909 B.n619 B.n618 10.6151
R1910 B.n619 B.n513 10.6151
R1911 B.n626 B.n625 10.6151
R1912 B.n627 B.n626 10.6151
R1913 B.n627 B.n508 10.6151
R1914 B.n633 B.n508 10.6151
R1915 B.n634 B.n633 10.6151
R1916 B.n635 B.n634 10.6151
R1917 B.n635 B.n506 10.6151
R1918 B.n641 B.n506 10.6151
R1919 B.n642 B.n641 10.6151
R1920 B.n644 B.n502 10.6151
R1921 B.n650 B.n502 10.6151
R1922 B.n651 B.n650 10.6151
R1923 B.n652 B.n651 10.6151
R1924 B.n652 B.n500 10.6151
R1925 B.n658 B.n500 10.6151
R1926 B.n659 B.n658 10.6151
R1927 B.n660 B.n659 10.6151
R1928 B.n660 B.n498 10.6151
R1929 B.n666 B.n498 10.6151
R1930 B.n667 B.n666 10.6151
R1931 B.n668 B.n667 10.6151
R1932 B.n668 B.n496 10.6151
R1933 B.n674 B.n496 10.6151
R1934 B.n675 B.n674 10.6151
R1935 B.n676 B.n675 10.6151
R1936 B.n676 B.n494 10.6151
R1937 B.n682 B.n494 10.6151
R1938 B.n683 B.n682 10.6151
R1939 B.n684 B.n683 10.6151
R1940 B.n684 B.n492 10.6151
R1941 B.n690 B.n492 10.6151
R1942 B.n691 B.n690 10.6151
R1943 B.n692 B.n691 10.6151
R1944 B.n692 B.n490 10.6151
R1945 B.n698 B.n490 10.6151
R1946 B.n699 B.n698 10.6151
R1947 B.n700 B.n699 10.6151
R1948 B.n700 B.n488 10.6151
R1949 B.n706 B.n488 10.6151
R1950 B.n707 B.n706 10.6151
R1951 B.n708 B.n707 10.6151
R1952 B.n708 B.n486 10.6151
R1953 B.n714 B.n486 10.6151
R1954 B.n715 B.n714 10.6151
R1955 B.n716 B.n715 10.6151
R1956 B.n716 B.n484 10.6151
R1957 B.n722 B.n484 10.6151
R1958 B.n723 B.n722 10.6151
R1959 B.n724 B.n723 10.6151
R1960 B.n724 B.n482 10.6151
R1961 B.n482 B.n481 10.6151
R1962 B.n731 B.n481 10.6151
R1963 B.n732 B.n731 10.6151
R1964 B.n738 B.n737 10.6151
R1965 B.n739 B.n738 10.6151
R1966 B.n739 B.n469 10.6151
R1967 B.n749 B.n469 10.6151
R1968 B.n750 B.n749 10.6151
R1969 B.n751 B.n750 10.6151
R1970 B.n751 B.n461 10.6151
R1971 B.n761 B.n461 10.6151
R1972 B.n762 B.n761 10.6151
R1973 B.n763 B.n762 10.6151
R1974 B.n763 B.n453 10.6151
R1975 B.n773 B.n453 10.6151
R1976 B.n774 B.n773 10.6151
R1977 B.n775 B.n774 10.6151
R1978 B.n775 B.n445 10.6151
R1979 B.n785 B.n445 10.6151
R1980 B.n786 B.n785 10.6151
R1981 B.n787 B.n786 10.6151
R1982 B.n787 B.n437 10.6151
R1983 B.n797 B.n437 10.6151
R1984 B.n798 B.n797 10.6151
R1985 B.n799 B.n798 10.6151
R1986 B.n799 B.n429 10.6151
R1987 B.n809 B.n429 10.6151
R1988 B.n810 B.n809 10.6151
R1989 B.n811 B.n810 10.6151
R1990 B.n811 B.n421 10.6151
R1991 B.n821 B.n421 10.6151
R1992 B.n822 B.n821 10.6151
R1993 B.n823 B.n822 10.6151
R1994 B.n823 B.n413 10.6151
R1995 B.n833 B.n413 10.6151
R1996 B.n834 B.n833 10.6151
R1997 B.n835 B.n834 10.6151
R1998 B.n835 B.n405 10.6151
R1999 B.n845 B.n405 10.6151
R2000 B.n846 B.n845 10.6151
R2001 B.n847 B.n846 10.6151
R2002 B.n847 B.n397 10.6151
R2003 B.n857 B.n397 10.6151
R2004 B.n858 B.n857 10.6151
R2005 B.n859 B.n858 10.6151
R2006 B.n859 B.n389 10.6151
R2007 B.n869 B.n389 10.6151
R2008 B.n870 B.n869 10.6151
R2009 B.n871 B.n870 10.6151
R2010 B.n871 B.n381 10.6151
R2011 B.n881 B.n381 10.6151
R2012 B.n882 B.n881 10.6151
R2013 B.n883 B.n882 10.6151
R2014 B.n883 B.n373 10.6151
R2015 B.n894 B.n373 10.6151
R2016 B.n895 B.n894 10.6151
R2017 B.n896 B.n895 10.6151
R2018 B.n896 B.n366 10.6151
R2019 B.n907 B.n366 10.6151
R2020 B.n908 B.n907 10.6151
R2021 B.n909 B.n908 10.6151
R2022 B.n909 B.n0 10.6151
R2023 B.n1111 B.n1 10.6151
R2024 B.n1111 B.n1110 10.6151
R2025 B.n1110 B.n1109 10.6151
R2026 B.n1109 B.n10 10.6151
R2027 B.n1103 B.n10 10.6151
R2028 B.n1103 B.n1102 10.6151
R2029 B.n1102 B.n1101 10.6151
R2030 B.n1101 B.n16 10.6151
R2031 B.n1095 B.n16 10.6151
R2032 B.n1095 B.n1094 10.6151
R2033 B.n1094 B.n1093 10.6151
R2034 B.n1093 B.n24 10.6151
R2035 B.n1087 B.n24 10.6151
R2036 B.n1087 B.n1086 10.6151
R2037 B.n1086 B.n1085 10.6151
R2038 B.n1085 B.n31 10.6151
R2039 B.n1079 B.n31 10.6151
R2040 B.n1079 B.n1078 10.6151
R2041 B.n1078 B.n1077 10.6151
R2042 B.n1077 B.n38 10.6151
R2043 B.n1071 B.n38 10.6151
R2044 B.n1071 B.n1070 10.6151
R2045 B.n1070 B.n1069 10.6151
R2046 B.n1069 B.n45 10.6151
R2047 B.n1063 B.n45 10.6151
R2048 B.n1063 B.n1062 10.6151
R2049 B.n1062 B.n1061 10.6151
R2050 B.n1061 B.n52 10.6151
R2051 B.n1055 B.n52 10.6151
R2052 B.n1055 B.n1054 10.6151
R2053 B.n1054 B.n1053 10.6151
R2054 B.n1053 B.n59 10.6151
R2055 B.n1047 B.n59 10.6151
R2056 B.n1047 B.n1046 10.6151
R2057 B.n1046 B.n1045 10.6151
R2058 B.n1045 B.n66 10.6151
R2059 B.n1039 B.n66 10.6151
R2060 B.n1039 B.n1038 10.6151
R2061 B.n1038 B.n1037 10.6151
R2062 B.n1037 B.n73 10.6151
R2063 B.n1031 B.n73 10.6151
R2064 B.n1031 B.n1030 10.6151
R2065 B.n1030 B.n1029 10.6151
R2066 B.n1029 B.n80 10.6151
R2067 B.n1023 B.n80 10.6151
R2068 B.n1023 B.n1022 10.6151
R2069 B.n1022 B.n1021 10.6151
R2070 B.n1021 B.n87 10.6151
R2071 B.n1015 B.n87 10.6151
R2072 B.n1015 B.n1014 10.6151
R2073 B.n1014 B.n1013 10.6151
R2074 B.n1013 B.n94 10.6151
R2075 B.n1007 B.n94 10.6151
R2076 B.n1007 B.n1006 10.6151
R2077 B.n1006 B.n1005 10.6151
R2078 B.n1005 B.n101 10.6151
R2079 B.n999 B.n101 10.6151
R2080 B.n999 B.n998 10.6151
R2081 B.n998 B.n997 10.6151
R2082 B.n253 B.n252 9.36635
R2083 B.n275 B.n274 9.36635
R2084 B.n513 B.n512 9.36635
R2085 B.n644 B.n643 9.36635
R2086 B.n891 B.t5 8.91701
R2087 B.n18 B.t0 8.91701
R2088 B.n801 B.t7 6.53927
R2089 B.t3 B.n1041 6.53927
R2090 B.t6 B.n391 5.35041
R2091 B.n1082 B.t4 5.35041
R2092 B.n1117 B.n0 2.81026
R2093 B.n1117 B.n1 2.81026
R2094 B.n254 B.n253 1.24928
R2095 B.n274 B.n273 1.24928
R2096 B.n625 B.n512 1.24928
R2097 B.n643 B.n642 1.24928
R2098 VN.n64 VN.n63 161.3
R2099 VN.n62 VN.n34 161.3
R2100 VN.n61 VN.n60 161.3
R2101 VN.n59 VN.n35 161.3
R2102 VN.n58 VN.n57 161.3
R2103 VN.n56 VN.n36 161.3
R2104 VN.n55 VN.n54 161.3
R2105 VN.n53 VN.n52 161.3
R2106 VN.n51 VN.n38 161.3
R2107 VN.n50 VN.n49 161.3
R2108 VN.n48 VN.n39 161.3
R2109 VN.n47 VN.n46 161.3
R2110 VN.n45 VN.n40 161.3
R2111 VN.n44 VN.n43 161.3
R2112 VN.n31 VN.n30 161.3
R2113 VN.n29 VN.n1 161.3
R2114 VN.n28 VN.n27 161.3
R2115 VN.n26 VN.n2 161.3
R2116 VN.n25 VN.n24 161.3
R2117 VN.n23 VN.n3 161.3
R2118 VN.n22 VN.n21 161.3
R2119 VN.n20 VN.n19 161.3
R2120 VN.n18 VN.n5 161.3
R2121 VN.n17 VN.n16 161.3
R2122 VN.n15 VN.n6 161.3
R2123 VN.n14 VN.n13 161.3
R2124 VN.n12 VN.n7 161.3
R2125 VN.n11 VN.n10 161.3
R2126 VN.n42 VN.t2 132.793
R2127 VN.n9 VN.t6 132.793
R2128 VN.n8 VN.t4 99.9513
R2129 VN.n4 VN.t5 99.9513
R2130 VN.n0 VN.t3 99.9513
R2131 VN.n41 VN.t0 99.9513
R2132 VN.n37 VN.t7 99.9513
R2133 VN.n33 VN.t1 99.9513
R2134 VN.n32 VN.n0 76.3659
R2135 VN.n65 VN.n33 76.3659
R2136 VN.n9 VN.n8 61.53
R2137 VN.n42 VN.n41 61.53
R2138 VN VN.n65 54.8238
R2139 VN.n28 VN.n2 42.4359
R2140 VN.n61 VN.n35 42.4359
R2141 VN.n13 VN.n6 40.4934
R2142 VN.n17 VN.n6 40.4934
R2143 VN.n46 VN.n39 40.4934
R2144 VN.n50 VN.n39 40.4934
R2145 VN.n24 VN.n2 38.5509
R2146 VN.n57 VN.n35 38.5509
R2147 VN.n12 VN.n11 24.4675
R2148 VN.n13 VN.n12 24.4675
R2149 VN.n18 VN.n17 24.4675
R2150 VN.n19 VN.n18 24.4675
R2151 VN.n23 VN.n22 24.4675
R2152 VN.n24 VN.n23 24.4675
R2153 VN.n29 VN.n28 24.4675
R2154 VN.n30 VN.n29 24.4675
R2155 VN.n46 VN.n45 24.4675
R2156 VN.n45 VN.n44 24.4675
R2157 VN.n57 VN.n56 24.4675
R2158 VN.n56 VN.n55 24.4675
R2159 VN.n52 VN.n51 24.4675
R2160 VN.n51 VN.n50 24.4675
R2161 VN.n63 VN.n62 24.4675
R2162 VN.n62 VN.n61 24.4675
R2163 VN.n30 VN.n0 13.702
R2164 VN.n63 VN.n33 13.702
R2165 VN.n11 VN.n8 12.7233
R2166 VN.n19 VN.n4 12.7233
R2167 VN.n44 VN.n41 12.7233
R2168 VN.n52 VN.n37 12.7233
R2169 VN.n22 VN.n4 11.7447
R2170 VN.n55 VN.n37 11.7447
R2171 VN.n43 VN.n42 4.20582
R2172 VN.n10 VN.n9 4.20582
R2173 VN.n65 VN.n64 0.354971
R2174 VN.n32 VN.n31 0.354971
R2175 VN VN.n32 0.26696
R2176 VN.n64 VN.n34 0.189894
R2177 VN.n60 VN.n34 0.189894
R2178 VN.n60 VN.n59 0.189894
R2179 VN.n59 VN.n58 0.189894
R2180 VN.n58 VN.n36 0.189894
R2181 VN.n54 VN.n36 0.189894
R2182 VN.n54 VN.n53 0.189894
R2183 VN.n53 VN.n38 0.189894
R2184 VN.n49 VN.n38 0.189894
R2185 VN.n49 VN.n48 0.189894
R2186 VN.n48 VN.n47 0.189894
R2187 VN.n47 VN.n40 0.189894
R2188 VN.n43 VN.n40 0.189894
R2189 VN.n10 VN.n7 0.189894
R2190 VN.n14 VN.n7 0.189894
R2191 VN.n15 VN.n14 0.189894
R2192 VN.n16 VN.n15 0.189894
R2193 VN.n16 VN.n5 0.189894
R2194 VN.n20 VN.n5 0.189894
R2195 VN.n21 VN.n20 0.189894
R2196 VN.n21 VN.n3 0.189894
R2197 VN.n25 VN.n3 0.189894
R2198 VN.n26 VN.n25 0.189894
R2199 VN.n27 VN.n26 0.189894
R2200 VN.n27 VN.n1 0.189894
R2201 VN.n31 VN.n1 0.189894
R2202 VDD2.n2 VDD2.n1 63.669
R2203 VDD2.n2 VDD2.n0 63.669
R2204 VDD2 VDD2.n5 63.666
R2205 VDD2.n4 VDD2.n3 62.2071
R2206 VDD2.n4 VDD2.n2 48.7756
R2207 VDD2 VDD2.n4 1.57593
R2208 VDD2.n5 VDD2.t7 1.4971
R2209 VDD2.n5 VDD2.t5 1.4971
R2210 VDD2.n3 VDD2.t6 1.4971
R2211 VDD2.n3 VDD2.t0 1.4971
R2212 VDD2.n1 VDD2.t2 1.4971
R2213 VDD2.n1 VDD2.t4 1.4971
R2214 VDD2.n0 VDD2.t1 1.4971
R2215 VDD2.n0 VDD2.t3 1.4971
C0 VP VN 8.61542f
C1 VTAIL VP 10.4509f
C2 VTAIL VN 10.436799f
C3 VDD2 VDD1 2.08194f
C4 VP VDD1 10.331f
C5 VDD1 VN 0.15239f
C6 VTAIL VDD1 8.644441f
C7 VDD2 VP 0.582049f
C8 VDD2 VN 9.903059f
C9 VDD2 VTAIL 8.702809f
C10 VDD2 B 6.085445f
C11 VDD1 B 6.58357f
C12 VTAIL B 11.622469f
C13 VN B 17.88327f
C14 VP B 16.507433f
C15 VDD2.t1 B 0.280854f
C16 VDD2.t3 B 0.280854f
C17 VDD2.n0 B 2.53147f
C18 VDD2.t2 B 0.280854f
C19 VDD2.t4 B 0.280854f
C20 VDD2.n1 B 2.53147f
C21 VDD2.n2 B 3.97704f
C22 VDD2.t6 B 0.280854f
C23 VDD2.t0 B 0.280854f
C24 VDD2.n3 B 2.51714f
C25 VDD2.n4 B 3.49287f
C26 VDD2.t7 B 0.280854f
C27 VDD2.t5 B 0.280854f
C28 VDD2.n5 B 2.53141f
C29 VN.t3 B 2.20325f
C30 VN.n0 B 0.842759f
C31 VN.n1 B 0.01911f
C32 VN.n2 B 0.015547f
C33 VN.n3 B 0.01911f
C34 VN.t5 B 2.20325f
C35 VN.n4 B 0.770981f
C36 VN.n5 B 0.01911f
C37 VN.n6 B 0.015448f
C38 VN.n7 B 0.01911f
C39 VN.t4 B 2.20325f
C40 VN.n8 B 0.834104f
C41 VN.t6 B 2.4269f
C42 VN.n9 B 0.797856f
C43 VN.n10 B 0.222281f
C44 VN.n11 B 0.027176f
C45 VN.n12 B 0.035616f
C46 VN.n13 B 0.03798f
C47 VN.n14 B 0.01911f
C48 VN.n15 B 0.01911f
C49 VN.n16 B 0.01911f
C50 VN.n17 B 0.03798f
C51 VN.n18 B 0.035616f
C52 VN.n19 B 0.027176f
C53 VN.n20 B 0.01911f
C54 VN.n21 B 0.01911f
C55 VN.n22 B 0.026472f
C56 VN.n23 B 0.035616f
C57 VN.n24 B 0.038312f
C58 VN.n25 B 0.01911f
C59 VN.n26 B 0.01911f
C60 VN.n27 B 0.01911f
C61 VN.n28 B 0.03755f
C62 VN.n29 B 0.035616f
C63 VN.n30 B 0.027879f
C64 VN.n31 B 0.030843f
C65 VN.n32 B 0.046088f
C66 VN.t1 B 2.20325f
C67 VN.n33 B 0.842759f
C68 VN.n34 B 0.01911f
C69 VN.n35 B 0.015547f
C70 VN.n36 B 0.01911f
C71 VN.t7 B 2.20325f
C72 VN.n37 B 0.770981f
C73 VN.n38 B 0.01911f
C74 VN.n39 B 0.015448f
C75 VN.n40 B 0.01911f
C76 VN.t0 B 2.20325f
C77 VN.n41 B 0.834104f
C78 VN.t2 B 2.4269f
C79 VN.n42 B 0.797856f
C80 VN.n43 B 0.222281f
C81 VN.n44 B 0.027176f
C82 VN.n45 B 0.035616f
C83 VN.n46 B 0.03798f
C84 VN.n47 B 0.01911f
C85 VN.n48 B 0.01911f
C86 VN.n49 B 0.01911f
C87 VN.n50 B 0.03798f
C88 VN.n51 B 0.035616f
C89 VN.n52 B 0.027176f
C90 VN.n53 B 0.01911f
C91 VN.n54 B 0.01911f
C92 VN.n55 B 0.026472f
C93 VN.n56 B 0.035616f
C94 VN.n57 B 0.038312f
C95 VN.n58 B 0.01911f
C96 VN.n59 B 0.01911f
C97 VN.n60 B 0.01911f
C98 VN.n61 B 0.03755f
C99 VN.n62 B 0.035616f
C100 VN.n63 B 0.027879f
C101 VN.n64 B 0.030843f
C102 VN.n65 B 1.23911f
C103 VDD1.t2 B 0.283565f
C104 VDD1.t0 B 0.283565f
C105 VDD1.n0 B 2.55723f
C106 VDD1.t6 B 0.283565f
C107 VDD1.t7 B 0.283565f
C108 VDD1.n1 B 2.5559f
C109 VDD1.t3 B 0.283565f
C110 VDD1.t5 B 0.283565f
C111 VDD1.n2 B 2.5559f
C112 VDD1.n3 B 4.07154f
C113 VDD1.t4 B 0.283565f
C114 VDD1.t1 B 0.283565f
C115 VDD1.n4 B 2.54143f
C116 VDD1.n5 B 3.56051f
C117 VTAIL.t4 B 0.207719f
C118 VTAIL.t1 B 0.207719f
C119 VTAIL.n0 B 1.80247f
C120 VTAIL.n1 B 0.395547f
C121 VTAIL.t0 B 2.30019f
C122 VTAIL.n2 B 0.490692f
C123 VTAIL.t11 B 2.30019f
C124 VTAIL.n3 B 0.490692f
C125 VTAIL.t10 B 0.207719f
C126 VTAIL.t15 B 0.207719f
C127 VTAIL.n4 B 1.80247f
C128 VTAIL.n5 B 0.58609f
C129 VTAIL.t14 B 2.30019f
C130 VTAIL.n6 B 1.65493f
C131 VTAIL.t7 B 2.30019f
C132 VTAIL.n7 B 1.65493f
C133 VTAIL.t2 B 0.207719f
C134 VTAIL.t6 B 0.207719f
C135 VTAIL.n8 B 1.80247f
C136 VTAIL.n9 B 0.586092f
C137 VTAIL.t5 B 2.30019f
C138 VTAIL.n10 B 0.490686f
C139 VTAIL.t12 B 2.30019f
C140 VTAIL.n11 B 0.490686f
C141 VTAIL.t13 B 0.207719f
C142 VTAIL.t8 B 0.207719f
C143 VTAIL.n12 B 1.80247f
C144 VTAIL.n13 B 0.586092f
C145 VTAIL.t9 B 2.30019f
C146 VTAIL.n14 B 1.65493f
C147 VTAIL.t3 B 2.30019f
C148 VTAIL.n15 B 1.65121f
C149 VP.t2 B 2.24345f
C150 VP.n0 B 0.858137f
C151 VP.n1 B 0.019458f
C152 VP.n2 B 0.015831f
C153 VP.n3 B 0.019458f
C154 VP.t4 B 2.24345f
C155 VP.n4 B 0.785049f
C156 VP.n5 B 0.019458f
C157 VP.n6 B 0.01573f
C158 VP.n7 B 0.019458f
C159 VP.t0 B 2.24345f
C160 VP.n8 B 0.785049f
C161 VP.n9 B 0.019458f
C162 VP.n10 B 0.015831f
C163 VP.n11 B 0.019458f
C164 VP.t1 B 2.24345f
C165 VP.n12 B 0.858137f
C166 VP.t6 B 2.24345f
C167 VP.n13 B 0.858137f
C168 VP.n14 B 0.019458f
C169 VP.n15 B 0.015831f
C170 VP.n16 B 0.019458f
C171 VP.t3 B 2.24345f
C172 VP.n17 B 0.785049f
C173 VP.n18 B 0.019458f
C174 VP.n19 B 0.01573f
C175 VP.n20 B 0.019458f
C176 VP.t7 B 2.24345f
C177 VP.n21 B 0.849324f
C178 VP.t5 B 2.47119f
C179 VP.n22 B 0.812415f
C180 VP.n23 B 0.226338f
C181 VP.n24 B 0.027671f
C182 VP.n25 B 0.036266f
C183 VP.n26 B 0.038673f
C184 VP.n27 B 0.019458f
C185 VP.n28 B 0.019458f
C186 VP.n29 B 0.019458f
C187 VP.n30 B 0.038673f
C188 VP.n31 B 0.036266f
C189 VP.n32 B 0.027671f
C190 VP.n33 B 0.019458f
C191 VP.n34 B 0.019458f
C192 VP.n35 B 0.026955f
C193 VP.n36 B 0.036266f
C194 VP.n37 B 0.039011f
C195 VP.n38 B 0.019458f
C196 VP.n39 B 0.019458f
C197 VP.n40 B 0.019458f
C198 VP.n41 B 0.038235f
C199 VP.n42 B 0.036266f
C200 VP.n43 B 0.028388f
C201 VP.n44 B 0.031406f
C202 VP.n45 B 1.25399f
C203 VP.n46 B 1.26679f
C204 VP.n47 B 0.031406f
C205 VP.n48 B 0.028388f
C206 VP.n49 B 0.036266f
C207 VP.n50 B 0.038235f
C208 VP.n51 B 0.019458f
C209 VP.n52 B 0.019458f
C210 VP.n53 B 0.019458f
C211 VP.n54 B 0.039011f
C212 VP.n55 B 0.036266f
C213 VP.n56 B 0.026955f
C214 VP.n57 B 0.019458f
C215 VP.n58 B 0.019458f
C216 VP.n59 B 0.027671f
C217 VP.n60 B 0.036266f
C218 VP.n61 B 0.038673f
C219 VP.n62 B 0.019458f
C220 VP.n63 B 0.019458f
C221 VP.n64 B 0.019458f
C222 VP.n65 B 0.038673f
C223 VP.n66 B 0.036266f
C224 VP.n67 B 0.027671f
C225 VP.n68 B 0.019458f
C226 VP.n69 B 0.019458f
C227 VP.n70 B 0.026955f
C228 VP.n71 B 0.036266f
C229 VP.n72 B 0.039011f
C230 VP.n73 B 0.019458f
C231 VP.n74 B 0.019458f
C232 VP.n75 B 0.019458f
C233 VP.n76 B 0.038235f
C234 VP.n77 B 0.036266f
C235 VP.n78 B 0.028388f
C236 VP.n79 B 0.031406f
C237 VP.n80 B 0.046929f
.ends

