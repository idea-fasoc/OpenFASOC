* NGSPICE file created from diff_pair_sample_0479.ext - technology: sky130A

.subckt diff_pair_sample_0479 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=2.9835 ps=16.08 w=7.65 l=2.25
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=0 ps=0 w=7.65 l=2.25
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=2.9835 ps=16.08 w=7.65 l=2.25
X3 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=2.9835 ps=16.08 w=7.65 l=2.25
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=0 ps=0 w=7.65 l=2.25
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=2.9835 ps=16.08 w=7.65 l=2.25
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=0 ps=0 w=7.65 l=2.25
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9835 pd=16.08 as=0 ps=0 w=7.65 l=2.25
R0 VP.n0 VP.t0 171.543
R1 VP.n0 VP.t1 131.111
R2 VP VP.n0 0.336784
R3 VTAIL.n1 VTAIL.t1 54.2735
R4 VTAIL.n3 VTAIL.t0 54.2733
R5 VTAIL.n0 VTAIL.t3 54.2733
R6 VTAIL.n2 VTAIL.t2 54.2733
R7 VTAIL.n1 VTAIL.n0 23.41
R8 VTAIL.n3 VTAIL.n2 21.1858
R9 VTAIL.n2 VTAIL.n1 1.5824
R10 VTAIL VTAIL.n0 1.08455
R11 VTAIL VTAIL.n3 0.498345
R12 VDD1 VDD1.t0 106.736
R13 VDD1 VDD1.t1 71.5663
R14 B.n533 B.n532 585
R15 B.n534 B.n533 585
R16 B.n214 B.n80 585
R17 B.n213 B.n212 585
R18 B.n211 B.n210 585
R19 B.n209 B.n208 585
R20 B.n207 B.n206 585
R21 B.n205 B.n204 585
R22 B.n203 B.n202 585
R23 B.n201 B.n200 585
R24 B.n199 B.n198 585
R25 B.n197 B.n196 585
R26 B.n195 B.n194 585
R27 B.n193 B.n192 585
R28 B.n191 B.n190 585
R29 B.n189 B.n188 585
R30 B.n187 B.n186 585
R31 B.n185 B.n184 585
R32 B.n183 B.n182 585
R33 B.n181 B.n180 585
R34 B.n179 B.n178 585
R35 B.n177 B.n176 585
R36 B.n175 B.n174 585
R37 B.n173 B.n172 585
R38 B.n171 B.n170 585
R39 B.n169 B.n168 585
R40 B.n167 B.n166 585
R41 B.n165 B.n164 585
R42 B.n163 B.n162 585
R43 B.n161 B.n160 585
R44 B.n159 B.n158 585
R45 B.n157 B.n156 585
R46 B.n155 B.n154 585
R47 B.n153 B.n152 585
R48 B.n151 B.n150 585
R49 B.n149 B.n148 585
R50 B.n147 B.n146 585
R51 B.n145 B.n144 585
R52 B.n143 B.n142 585
R53 B.n140 B.n139 585
R54 B.n138 B.n137 585
R55 B.n136 B.n135 585
R56 B.n134 B.n133 585
R57 B.n132 B.n131 585
R58 B.n130 B.n129 585
R59 B.n128 B.n127 585
R60 B.n126 B.n125 585
R61 B.n124 B.n123 585
R62 B.n122 B.n121 585
R63 B.n120 B.n119 585
R64 B.n118 B.n117 585
R65 B.n116 B.n115 585
R66 B.n114 B.n113 585
R67 B.n112 B.n111 585
R68 B.n110 B.n109 585
R69 B.n108 B.n107 585
R70 B.n106 B.n105 585
R71 B.n104 B.n103 585
R72 B.n102 B.n101 585
R73 B.n100 B.n99 585
R74 B.n98 B.n97 585
R75 B.n96 B.n95 585
R76 B.n94 B.n93 585
R77 B.n92 B.n91 585
R78 B.n90 B.n89 585
R79 B.n88 B.n87 585
R80 B.n47 B.n46 585
R81 B.n537 B.n536 585
R82 B.n531 B.n81 585
R83 B.n81 B.n44 585
R84 B.n530 B.n43 585
R85 B.n541 B.n43 585
R86 B.n529 B.n42 585
R87 B.n542 B.n42 585
R88 B.n528 B.n41 585
R89 B.n543 B.n41 585
R90 B.n527 B.n526 585
R91 B.n526 B.n37 585
R92 B.n525 B.n36 585
R93 B.n549 B.n36 585
R94 B.n524 B.n35 585
R95 B.n550 B.n35 585
R96 B.n523 B.n34 585
R97 B.n551 B.n34 585
R98 B.n522 B.n521 585
R99 B.n521 B.n30 585
R100 B.n520 B.n29 585
R101 B.n557 B.n29 585
R102 B.n519 B.n28 585
R103 B.n558 B.n28 585
R104 B.n518 B.n27 585
R105 B.n559 B.n27 585
R106 B.n517 B.n516 585
R107 B.n516 B.n23 585
R108 B.n515 B.n22 585
R109 B.n565 B.n22 585
R110 B.n514 B.n21 585
R111 B.n566 B.n21 585
R112 B.n513 B.n20 585
R113 B.n567 B.n20 585
R114 B.n512 B.n511 585
R115 B.n511 B.n16 585
R116 B.n510 B.n15 585
R117 B.n573 B.n15 585
R118 B.n509 B.n14 585
R119 B.n574 B.n14 585
R120 B.n508 B.n13 585
R121 B.n575 B.n13 585
R122 B.n507 B.n506 585
R123 B.n506 B.n12 585
R124 B.n505 B.n504 585
R125 B.n505 B.n8 585
R126 B.n503 B.n7 585
R127 B.n582 B.n7 585
R128 B.n502 B.n6 585
R129 B.n583 B.n6 585
R130 B.n501 B.n5 585
R131 B.n584 B.n5 585
R132 B.n500 B.n499 585
R133 B.n499 B.n4 585
R134 B.n498 B.n215 585
R135 B.n498 B.n497 585
R136 B.n488 B.n216 585
R137 B.n217 B.n216 585
R138 B.n490 B.n489 585
R139 B.n491 B.n490 585
R140 B.n487 B.n221 585
R141 B.n225 B.n221 585
R142 B.n486 B.n485 585
R143 B.n485 B.n484 585
R144 B.n223 B.n222 585
R145 B.n224 B.n223 585
R146 B.n477 B.n476 585
R147 B.n478 B.n477 585
R148 B.n475 B.n230 585
R149 B.n230 B.n229 585
R150 B.n474 B.n473 585
R151 B.n473 B.n472 585
R152 B.n232 B.n231 585
R153 B.n233 B.n232 585
R154 B.n465 B.n464 585
R155 B.n466 B.n465 585
R156 B.n463 B.n238 585
R157 B.n238 B.n237 585
R158 B.n462 B.n461 585
R159 B.n461 B.n460 585
R160 B.n240 B.n239 585
R161 B.n241 B.n240 585
R162 B.n453 B.n452 585
R163 B.n454 B.n453 585
R164 B.n451 B.n246 585
R165 B.n246 B.n245 585
R166 B.n450 B.n449 585
R167 B.n449 B.n448 585
R168 B.n248 B.n247 585
R169 B.n249 B.n248 585
R170 B.n441 B.n440 585
R171 B.n442 B.n441 585
R172 B.n439 B.n254 585
R173 B.n254 B.n253 585
R174 B.n438 B.n437 585
R175 B.n437 B.n436 585
R176 B.n256 B.n255 585
R177 B.n257 B.n256 585
R178 B.n432 B.n431 585
R179 B.n260 B.n259 585
R180 B.n428 B.n427 585
R181 B.n429 B.n428 585
R182 B.n426 B.n293 585
R183 B.n425 B.n424 585
R184 B.n423 B.n422 585
R185 B.n421 B.n420 585
R186 B.n419 B.n418 585
R187 B.n417 B.n416 585
R188 B.n415 B.n414 585
R189 B.n413 B.n412 585
R190 B.n411 B.n410 585
R191 B.n409 B.n408 585
R192 B.n407 B.n406 585
R193 B.n405 B.n404 585
R194 B.n403 B.n402 585
R195 B.n401 B.n400 585
R196 B.n399 B.n398 585
R197 B.n397 B.n396 585
R198 B.n395 B.n394 585
R199 B.n393 B.n392 585
R200 B.n391 B.n390 585
R201 B.n389 B.n388 585
R202 B.n387 B.n386 585
R203 B.n385 B.n384 585
R204 B.n383 B.n382 585
R205 B.n381 B.n380 585
R206 B.n379 B.n378 585
R207 B.n377 B.n376 585
R208 B.n375 B.n374 585
R209 B.n373 B.n372 585
R210 B.n371 B.n370 585
R211 B.n369 B.n368 585
R212 B.n367 B.n366 585
R213 B.n365 B.n364 585
R214 B.n363 B.n362 585
R215 B.n361 B.n360 585
R216 B.n359 B.n358 585
R217 B.n356 B.n355 585
R218 B.n354 B.n353 585
R219 B.n352 B.n351 585
R220 B.n350 B.n349 585
R221 B.n348 B.n347 585
R222 B.n346 B.n345 585
R223 B.n344 B.n343 585
R224 B.n342 B.n341 585
R225 B.n340 B.n339 585
R226 B.n338 B.n337 585
R227 B.n336 B.n335 585
R228 B.n334 B.n333 585
R229 B.n332 B.n331 585
R230 B.n330 B.n329 585
R231 B.n328 B.n327 585
R232 B.n326 B.n325 585
R233 B.n324 B.n323 585
R234 B.n322 B.n321 585
R235 B.n320 B.n319 585
R236 B.n318 B.n317 585
R237 B.n316 B.n315 585
R238 B.n314 B.n313 585
R239 B.n312 B.n311 585
R240 B.n310 B.n309 585
R241 B.n308 B.n307 585
R242 B.n306 B.n305 585
R243 B.n304 B.n303 585
R244 B.n302 B.n301 585
R245 B.n300 B.n299 585
R246 B.n433 B.n258 585
R247 B.n258 B.n257 585
R248 B.n435 B.n434 585
R249 B.n436 B.n435 585
R250 B.n252 B.n251 585
R251 B.n253 B.n252 585
R252 B.n444 B.n443 585
R253 B.n443 B.n442 585
R254 B.n445 B.n250 585
R255 B.n250 B.n249 585
R256 B.n447 B.n446 585
R257 B.n448 B.n447 585
R258 B.n244 B.n243 585
R259 B.n245 B.n244 585
R260 B.n456 B.n455 585
R261 B.n455 B.n454 585
R262 B.n457 B.n242 585
R263 B.n242 B.n241 585
R264 B.n459 B.n458 585
R265 B.n460 B.n459 585
R266 B.n236 B.n235 585
R267 B.n237 B.n236 585
R268 B.n468 B.n467 585
R269 B.n467 B.n466 585
R270 B.n469 B.n234 585
R271 B.n234 B.n233 585
R272 B.n471 B.n470 585
R273 B.n472 B.n471 585
R274 B.n228 B.n227 585
R275 B.n229 B.n228 585
R276 B.n480 B.n479 585
R277 B.n479 B.n478 585
R278 B.n481 B.n226 585
R279 B.n226 B.n224 585
R280 B.n483 B.n482 585
R281 B.n484 B.n483 585
R282 B.n220 B.n219 585
R283 B.n225 B.n220 585
R284 B.n493 B.n492 585
R285 B.n492 B.n491 585
R286 B.n494 B.n218 585
R287 B.n218 B.n217 585
R288 B.n496 B.n495 585
R289 B.n497 B.n496 585
R290 B.n3 B.n0 585
R291 B.n4 B.n3 585
R292 B.n581 B.n1 585
R293 B.n582 B.n581 585
R294 B.n580 B.n579 585
R295 B.n580 B.n8 585
R296 B.n578 B.n9 585
R297 B.n12 B.n9 585
R298 B.n577 B.n576 585
R299 B.n576 B.n575 585
R300 B.n11 B.n10 585
R301 B.n574 B.n11 585
R302 B.n572 B.n571 585
R303 B.n573 B.n572 585
R304 B.n570 B.n17 585
R305 B.n17 B.n16 585
R306 B.n569 B.n568 585
R307 B.n568 B.n567 585
R308 B.n19 B.n18 585
R309 B.n566 B.n19 585
R310 B.n564 B.n563 585
R311 B.n565 B.n564 585
R312 B.n562 B.n24 585
R313 B.n24 B.n23 585
R314 B.n561 B.n560 585
R315 B.n560 B.n559 585
R316 B.n26 B.n25 585
R317 B.n558 B.n26 585
R318 B.n556 B.n555 585
R319 B.n557 B.n556 585
R320 B.n554 B.n31 585
R321 B.n31 B.n30 585
R322 B.n553 B.n552 585
R323 B.n552 B.n551 585
R324 B.n33 B.n32 585
R325 B.n550 B.n33 585
R326 B.n548 B.n547 585
R327 B.n549 B.n548 585
R328 B.n546 B.n38 585
R329 B.n38 B.n37 585
R330 B.n545 B.n544 585
R331 B.n544 B.n543 585
R332 B.n40 B.n39 585
R333 B.n542 B.n40 585
R334 B.n540 B.n539 585
R335 B.n541 B.n540 585
R336 B.n538 B.n45 585
R337 B.n45 B.n44 585
R338 B.n585 B.n584 585
R339 B.n583 B.n2 585
R340 B.n536 B.n45 482.89
R341 B.n533 B.n81 482.89
R342 B.n299 B.n256 482.89
R343 B.n431 B.n258 482.89
R344 B.n85 B.t13 289.389
R345 B.n82 B.t2 289.389
R346 B.n297 B.t6 289.389
R347 B.n294 B.t10 289.389
R348 B.n534 B.n79 256.663
R349 B.n534 B.n78 256.663
R350 B.n534 B.n77 256.663
R351 B.n534 B.n76 256.663
R352 B.n534 B.n75 256.663
R353 B.n534 B.n74 256.663
R354 B.n534 B.n73 256.663
R355 B.n534 B.n72 256.663
R356 B.n534 B.n71 256.663
R357 B.n534 B.n70 256.663
R358 B.n534 B.n69 256.663
R359 B.n534 B.n68 256.663
R360 B.n534 B.n67 256.663
R361 B.n534 B.n66 256.663
R362 B.n534 B.n65 256.663
R363 B.n534 B.n64 256.663
R364 B.n534 B.n63 256.663
R365 B.n534 B.n62 256.663
R366 B.n534 B.n61 256.663
R367 B.n534 B.n60 256.663
R368 B.n534 B.n59 256.663
R369 B.n534 B.n58 256.663
R370 B.n534 B.n57 256.663
R371 B.n534 B.n56 256.663
R372 B.n534 B.n55 256.663
R373 B.n534 B.n54 256.663
R374 B.n534 B.n53 256.663
R375 B.n534 B.n52 256.663
R376 B.n534 B.n51 256.663
R377 B.n534 B.n50 256.663
R378 B.n534 B.n49 256.663
R379 B.n534 B.n48 256.663
R380 B.n535 B.n534 256.663
R381 B.n430 B.n429 256.663
R382 B.n429 B.n261 256.663
R383 B.n429 B.n262 256.663
R384 B.n429 B.n263 256.663
R385 B.n429 B.n264 256.663
R386 B.n429 B.n265 256.663
R387 B.n429 B.n266 256.663
R388 B.n429 B.n267 256.663
R389 B.n429 B.n268 256.663
R390 B.n429 B.n269 256.663
R391 B.n429 B.n270 256.663
R392 B.n429 B.n271 256.663
R393 B.n429 B.n272 256.663
R394 B.n429 B.n273 256.663
R395 B.n429 B.n274 256.663
R396 B.n429 B.n275 256.663
R397 B.n429 B.n276 256.663
R398 B.n429 B.n277 256.663
R399 B.n429 B.n278 256.663
R400 B.n429 B.n279 256.663
R401 B.n429 B.n280 256.663
R402 B.n429 B.n281 256.663
R403 B.n429 B.n282 256.663
R404 B.n429 B.n283 256.663
R405 B.n429 B.n284 256.663
R406 B.n429 B.n285 256.663
R407 B.n429 B.n286 256.663
R408 B.n429 B.n287 256.663
R409 B.n429 B.n288 256.663
R410 B.n429 B.n289 256.663
R411 B.n429 B.n290 256.663
R412 B.n429 B.n291 256.663
R413 B.n429 B.n292 256.663
R414 B.n587 B.n586 256.663
R415 B.n87 B.n47 163.367
R416 B.n91 B.n90 163.367
R417 B.n95 B.n94 163.367
R418 B.n99 B.n98 163.367
R419 B.n103 B.n102 163.367
R420 B.n107 B.n106 163.367
R421 B.n111 B.n110 163.367
R422 B.n115 B.n114 163.367
R423 B.n119 B.n118 163.367
R424 B.n123 B.n122 163.367
R425 B.n127 B.n126 163.367
R426 B.n131 B.n130 163.367
R427 B.n135 B.n134 163.367
R428 B.n139 B.n138 163.367
R429 B.n144 B.n143 163.367
R430 B.n148 B.n147 163.367
R431 B.n152 B.n151 163.367
R432 B.n156 B.n155 163.367
R433 B.n160 B.n159 163.367
R434 B.n164 B.n163 163.367
R435 B.n168 B.n167 163.367
R436 B.n172 B.n171 163.367
R437 B.n176 B.n175 163.367
R438 B.n180 B.n179 163.367
R439 B.n184 B.n183 163.367
R440 B.n188 B.n187 163.367
R441 B.n192 B.n191 163.367
R442 B.n196 B.n195 163.367
R443 B.n200 B.n199 163.367
R444 B.n204 B.n203 163.367
R445 B.n208 B.n207 163.367
R446 B.n212 B.n211 163.367
R447 B.n533 B.n80 163.367
R448 B.n437 B.n256 163.367
R449 B.n437 B.n254 163.367
R450 B.n441 B.n254 163.367
R451 B.n441 B.n248 163.367
R452 B.n449 B.n248 163.367
R453 B.n449 B.n246 163.367
R454 B.n453 B.n246 163.367
R455 B.n453 B.n240 163.367
R456 B.n461 B.n240 163.367
R457 B.n461 B.n238 163.367
R458 B.n465 B.n238 163.367
R459 B.n465 B.n232 163.367
R460 B.n473 B.n232 163.367
R461 B.n473 B.n230 163.367
R462 B.n477 B.n230 163.367
R463 B.n477 B.n223 163.367
R464 B.n485 B.n223 163.367
R465 B.n485 B.n221 163.367
R466 B.n490 B.n221 163.367
R467 B.n490 B.n216 163.367
R468 B.n498 B.n216 163.367
R469 B.n499 B.n498 163.367
R470 B.n499 B.n5 163.367
R471 B.n6 B.n5 163.367
R472 B.n7 B.n6 163.367
R473 B.n505 B.n7 163.367
R474 B.n506 B.n505 163.367
R475 B.n506 B.n13 163.367
R476 B.n14 B.n13 163.367
R477 B.n15 B.n14 163.367
R478 B.n511 B.n15 163.367
R479 B.n511 B.n20 163.367
R480 B.n21 B.n20 163.367
R481 B.n22 B.n21 163.367
R482 B.n516 B.n22 163.367
R483 B.n516 B.n27 163.367
R484 B.n28 B.n27 163.367
R485 B.n29 B.n28 163.367
R486 B.n521 B.n29 163.367
R487 B.n521 B.n34 163.367
R488 B.n35 B.n34 163.367
R489 B.n36 B.n35 163.367
R490 B.n526 B.n36 163.367
R491 B.n526 B.n41 163.367
R492 B.n42 B.n41 163.367
R493 B.n43 B.n42 163.367
R494 B.n81 B.n43 163.367
R495 B.n428 B.n260 163.367
R496 B.n428 B.n293 163.367
R497 B.n424 B.n423 163.367
R498 B.n420 B.n419 163.367
R499 B.n416 B.n415 163.367
R500 B.n412 B.n411 163.367
R501 B.n408 B.n407 163.367
R502 B.n404 B.n403 163.367
R503 B.n400 B.n399 163.367
R504 B.n396 B.n395 163.367
R505 B.n392 B.n391 163.367
R506 B.n388 B.n387 163.367
R507 B.n384 B.n383 163.367
R508 B.n380 B.n379 163.367
R509 B.n376 B.n375 163.367
R510 B.n372 B.n371 163.367
R511 B.n368 B.n367 163.367
R512 B.n364 B.n363 163.367
R513 B.n360 B.n359 163.367
R514 B.n355 B.n354 163.367
R515 B.n351 B.n350 163.367
R516 B.n347 B.n346 163.367
R517 B.n343 B.n342 163.367
R518 B.n339 B.n338 163.367
R519 B.n335 B.n334 163.367
R520 B.n331 B.n330 163.367
R521 B.n327 B.n326 163.367
R522 B.n323 B.n322 163.367
R523 B.n319 B.n318 163.367
R524 B.n315 B.n314 163.367
R525 B.n311 B.n310 163.367
R526 B.n307 B.n306 163.367
R527 B.n303 B.n302 163.367
R528 B.n435 B.n258 163.367
R529 B.n435 B.n252 163.367
R530 B.n443 B.n252 163.367
R531 B.n443 B.n250 163.367
R532 B.n447 B.n250 163.367
R533 B.n447 B.n244 163.367
R534 B.n455 B.n244 163.367
R535 B.n455 B.n242 163.367
R536 B.n459 B.n242 163.367
R537 B.n459 B.n236 163.367
R538 B.n467 B.n236 163.367
R539 B.n467 B.n234 163.367
R540 B.n471 B.n234 163.367
R541 B.n471 B.n228 163.367
R542 B.n479 B.n228 163.367
R543 B.n479 B.n226 163.367
R544 B.n483 B.n226 163.367
R545 B.n483 B.n220 163.367
R546 B.n492 B.n220 163.367
R547 B.n492 B.n218 163.367
R548 B.n496 B.n218 163.367
R549 B.n496 B.n3 163.367
R550 B.n585 B.n3 163.367
R551 B.n581 B.n2 163.367
R552 B.n581 B.n580 163.367
R553 B.n580 B.n9 163.367
R554 B.n576 B.n9 163.367
R555 B.n576 B.n11 163.367
R556 B.n572 B.n11 163.367
R557 B.n572 B.n17 163.367
R558 B.n568 B.n17 163.367
R559 B.n568 B.n19 163.367
R560 B.n564 B.n19 163.367
R561 B.n564 B.n24 163.367
R562 B.n560 B.n24 163.367
R563 B.n560 B.n26 163.367
R564 B.n556 B.n26 163.367
R565 B.n556 B.n31 163.367
R566 B.n552 B.n31 163.367
R567 B.n552 B.n33 163.367
R568 B.n548 B.n33 163.367
R569 B.n548 B.n38 163.367
R570 B.n544 B.n38 163.367
R571 B.n544 B.n40 163.367
R572 B.n540 B.n40 163.367
R573 B.n540 B.n45 163.367
R574 B.n82 B.t4 122.056
R575 B.n297 B.t9 122.056
R576 B.n85 B.t14 122.047
R577 B.n294 B.t12 122.047
R578 B.n429 B.n257 92.7665
R579 B.n534 B.n44 92.7665
R580 B.n83 B.t5 72.02
R581 B.n298 B.t8 72.02
R582 B.n86 B.t15 72.0112
R583 B.n295 B.t11 72.0112
R584 B.n536 B.n535 71.676
R585 B.n87 B.n48 71.676
R586 B.n91 B.n49 71.676
R587 B.n95 B.n50 71.676
R588 B.n99 B.n51 71.676
R589 B.n103 B.n52 71.676
R590 B.n107 B.n53 71.676
R591 B.n111 B.n54 71.676
R592 B.n115 B.n55 71.676
R593 B.n119 B.n56 71.676
R594 B.n123 B.n57 71.676
R595 B.n127 B.n58 71.676
R596 B.n131 B.n59 71.676
R597 B.n135 B.n60 71.676
R598 B.n139 B.n61 71.676
R599 B.n144 B.n62 71.676
R600 B.n148 B.n63 71.676
R601 B.n152 B.n64 71.676
R602 B.n156 B.n65 71.676
R603 B.n160 B.n66 71.676
R604 B.n164 B.n67 71.676
R605 B.n168 B.n68 71.676
R606 B.n172 B.n69 71.676
R607 B.n176 B.n70 71.676
R608 B.n180 B.n71 71.676
R609 B.n184 B.n72 71.676
R610 B.n188 B.n73 71.676
R611 B.n192 B.n74 71.676
R612 B.n196 B.n75 71.676
R613 B.n200 B.n76 71.676
R614 B.n204 B.n77 71.676
R615 B.n208 B.n78 71.676
R616 B.n212 B.n79 71.676
R617 B.n80 B.n79 71.676
R618 B.n211 B.n78 71.676
R619 B.n207 B.n77 71.676
R620 B.n203 B.n76 71.676
R621 B.n199 B.n75 71.676
R622 B.n195 B.n74 71.676
R623 B.n191 B.n73 71.676
R624 B.n187 B.n72 71.676
R625 B.n183 B.n71 71.676
R626 B.n179 B.n70 71.676
R627 B.n175 B.n69 71.676
R628 B.n171 B.n68 71.676
R629 B.n167 B.n67 71.676
R630 B.n163 B.n66 71.676
R631 B.n159 B.n65 71.676
R632 B.n155 B.n64 71.676
R633 B.n151 B.n63 71.676
R634 B.n147 B.n62 71.676
R635 B.n143 B.n61 71.676
R636 B.n138 B.n60 71.676
R637 B.n134 B.n59 71.676
R638 B.n130 B.n58 71.676
R639 B.n126 B.n57 71.676
R640 B.n122 B.n56 71.676
R641 B.n118 B.n55 71.676
R642 B.n114 B.n54 71.676
R643 B.n110 B.n53 71.676
R644 B.n106 B.n52 71.676
R645 B.n102 B.n51 71.676
R646 B.n98 B.n50 71.676
R647 B.n94 B.n49 71.676
R648 B.n90 B.n48 71.676
R649 B.n535 B.n47 71.676
R650 B.n431 B.n430 71.676
R651 B.n293 B.n261 71.676
R652 B.n423 B.n262 71.676
R653 B.n419 B.n263 71.676
R654 B.n415 B.n264 71.676
R655 B.n411 B.n265 71.676
R656 B.n407 B.n266 71.676
R657 B.n403 B.n267 71.676
R658 B.n399 B.n268 71.676
R659 B.n395 B.n269 71.676
R660 B.n391 B.n270 71.676
R661 B.n387 B.n271 71.676
R662 B.n383 B.n272 71.676
R663 B.n379 B.n273 71.676
R664 B.n375 B.n274 71.676
R665 B.n371 B.n275 71.676
R666 B.n367 B.n276 71.676
R667 B.n363 B.n277 71.676
R668 B.n359 B.n278 71.676
R669 B.n354 B.n279 71.676
R670 B.n350 B.n280 71.676
R671 B.n346 B.n281 71.676
R672 B.n342 B.n282 71.676
R673 B.n338 B.n283 71.676
R674 B.n334 B.n284 71.676
R675 B.n330 B.n285 71.676
R676 B.n326 B.n286 71.676
R677 B.n322 B.n287 71.676
R678 B.n318 B.n288 71.676
R679 B.n314 B.n289 71.676
R680 B.n310 B.n290 71.676
R681 B.n306 B.n291 71.676
R682 B.n302 B.n292 71.676
R683 B.n430 B.n260 71.676
R684 B.n424 B.n261 71.676
R685 B.n420 B.n262 71.676
R686 B.n416 B.n263 71.676
R687 B.n412 B.n264 71.676
R688 B.n408 B.n265 71.676
R689 B.n404 B.n266 71.676
R690 B.n400 B.n267 71.676
R691 B.n396 B.n268 71.676
R692 B.n392 B.n269 71.676
R693 B.n388 B.n270 71.676
R694 B.n384 B.n271 71.676
R695 B.n380 B.n272 71.676
R696 B.n376 B.n273 71.676
R697 B.n372 B.n274 71.676
R698 B.n368 B.n275 71.676
R699 B.n364 B.n276 71.676
R700 B.n360 B.n277 71.676
R701 B.n355 B.n278 71.676
R702 B.n351 B.n279 71.676
R703 B.n347 B.n280 71.676
R704 B.n343 B.n281 71.676
R705 B.n339 B.n282 71.676
R706 B.n335 B.n283 71.676
R707 B.n331 B.n284 71.676
R708 B.n327 B.n285 71.676
R709 B.n323 B.n286 71.676
R710 B.n319 B.n287 71.676
R711 B.n315 B.n288 71.676
R712 B.n311 B.n289 71.676
R713 B.n307 B.n290 71.676
R714 B.n303 B.n291 71.676
R715 B.n299 B.n292 71.676
R716 B.n586 B.n585 71.676
R717 B.n586 B.n2 71.676
R718 B.n141 B.n86 59.5399
R719 B.n84 B.n83 59.5399
R720 B.n357 B.n298 59.5399
R721 B.n296 B.n295 59.5399
R722 B.n436 B.n257 57.8728
R723 B.n436 B.n253 57.8728
R724 B.n442 B.n253 57.8728
R725 B.n442 B.n249 57.8728
R726 B.n448 B.n249 57.8728
R727 B.n448 B.n245 57.8728
R728 B.n454 B.n245 57.8728
R729 B.n460 B.n241 57.8728
R730 B.n460 B.n237 57.8728
R731 B.n466 B.n237 57.8728
R732 B.n466 B.n233 57.8728
R733 B.n472 B.n233 57.8728
R734 B.n472 B.n229 57.8728
R735 B.n478 B.n229 57.8728
R736 B.n478 B.n224 57.8728
R737 B.n484 B.n224 57.8728
R738 B.n484 B.n225 57.8728
R739 B.n491 B.n217 57.8728
R740 B.n497 B.n217 57.8728
R741 B.n497 B.n4 57.8728
R742 B.n584 B.n4 57.8728
R743 B.n584 B.n583 57.8728
R744 B.n583 B.n582 57.8728
R745 B.n582 B.n8 57.8728
R746 B.n12 B.n8 57.8728
R747 B.n575 B.n12 57.8728
R748 B.n574 B.n573 57.8728
R749 B.n573 B.n16 57.8728
R750 B.n567 B.n16 57.8728
R751 B.n567 B.n566 57.8728
R752 B.n566 B.n565 57.8728
R753 B.n565 B.n23 57.8728
R754 B.n559 B.n23 57.8728
R755 B.n559 B.n558 57.8728
R756 B.n558 B.n557 57.8728
R757 B.n557 B.n30 57.8728
R758 B.n551 B.n550 57.8728
R759 B.n550 B.n549 57.8728
R760 B.n549 B.n37 57.8728
R761 B.n543 B.n37 57.8728
R762 B.n543 B.n542 57.8728
R763 B.n542 B.n541 57.8728
R764 B.n541 B.n44 57.8728
R765 B.n491 B.t1 51.9154
R766 B.n575 B.t0 51.9154
R767 B.n86 B.n85 50.0369
R768 B.n83 B.n82 50.0369
R769 B.n298 B.n297 50.0369
R770 B.n295 B.n294 50.0369
R771 B.t7 B.n241 40.0005
R772 B.t3 B.n30 40.0005
R773 B.n433 B.n432 31.3761
R774 B.n300 B.n255 31.3761
R775 B.n532 B.n531 31.3761
R776 B.n538 B.n537 31.3761
R777 B B.n587 18.0485
R778 B.n454 B.t7 17.8728
R779 B.n551 B.t3 17.8728
R780 B.n434 B.n433 10.6151
R781 B.n434 B.n251 10.6151
R782 B.n444 B.n251 10.6151
R783 B.n445 B.n444 10.6151
R784 B.n446 B.n445 10.6151
R785 B.n446 B.n243 10.6151
R786 B.n456 B.n243 10.6151
R787 B.n457 B.n456 10.6151
R788 B.n458 B.n457 10.6151
R789 B.n458 B.n235 10.6151
R790 B.n468 B.n235 10.6151
R791 B.n469 B.n468 10.6151
R792 B.n470 B.n469 10.6151
R793 B.n470 B.n227 10.6151
R794 B.n480 B.n227 10.6151
R795 B.n481 B.n480 10.6151
R796 B.n482 B.n481 10.6151
R797 B.n482 B.n219 10.6151
R798 B.n493 B.n219 10.6151
R799 B.n494 B.n493 10.6151
R800 B.n495 B.n494 10.6151
R801 B.n495 B.n0 10.6151
R802 B.n432 B.n259 10.6151
R803 B.n427 B.n259 10.6151
R804 B.n427 B.n426 10.6151
R805 B.n426 B.n425 10.6151
R806 B.n425 B.n422 10.6151
R807 B.n422 B.n421 10.6151
R808 B.n421 B.n418 10.6151
R809 B.n418 B.n417 10.6151
R810 B.n417 B.n414 10.6151
R811 B.n414 B.n413 10.6151
R812 B.n413 B.n410 10.6151
R813 B.n410 B.n409 10.6151
R814 B.n409 B.n406 10.6151
R815 B.n406 B.n405 10.6151
R816 B.n405 B.n402 10.6151
R817 B.n402 B.n401 10.6151
R818 B.n401 B.n398 10.6151
R819 B.n398 B.n397 10.6151
R820 B.n397 B.n394 10.6151
R821 B.n394 B.n393 10.6151
R822 B.n393 B.n390 10.6151
R823 B.n390 B.n389 10.6151
R824 B.n389 B.n386 10.6151
R825 B.n386 B.n385 10.6151
R826 B.n385 B.n382 10.6151
R827 B.n382 B.n381 10.6151
R828 B.n381 B.n378 10.6151
R829 B.n378 B.n377 10.6151
R830 B.n374 B.n373 10.6151
R831 B.n373 B.n370 10.6151
R832 B.n370 B.n369 10.6151
R833 B.n369 B.n366 10.6151
R834 B.n366 B.n365 10.6151
R835 B.n365 B.n362 10.6151
R836 B.n362 B.n361 10.6151
R837 B.n361 B.n358 10.6151
R838 B.n356 B.n353 10.6151
R839 B.n353 B.n352 10.6151
R840 B.n352 B.n349 10.6151
R841 B.n349 B.n348 10.6151
R842 B.n348 B.n345 10.6151
R843 B.n345 B.n344 10.6151
R844 B.n344 B.n341 10.6151
R845 B.n341 B.n340 10.6151
R846 B.n340 B.n337 10.6151
R847 B.n337 B.n336 10.6151
R848 B.n336 B.n333 10.6151
R849 B.n333 B.n332 10.6151
R850 B.n332 B.n329 10.6151
R851 B.n329 B.n328 10.6151
R852 B.n328 B.n325 10.6151
R853 B.n325 B.n324 10.6151
R854 B.n324 B.n321 10.6151
R855 B.n321 B.n320 10.6151
R856 B.n320 B.n317 10.6151
R857 B.n317 B.n316 10.6151
R858 B.n316 B.n313 10.6151
R859 B.n313 B.n312 10.6151
R860 B.n312 B.n309 10.6151
R861 B.n309 B.n308 10.6151
R862 B.n308 B.n305 10.6151
R863 B.n305 B.n304 10.6151
R864 B.n304 B.n301 10.6151
R865 B.n301 B.n300 10.6151
R866 B.n438 B.n255 10.6151
R867 B.n439 B.n438 10.6151
R868 B.n440 B.n439 10.6151
R869 B.n440 B.n247 10.6151
R870 B.n450 B.n247 10.6151
R871 B.n451 B.n450 10.6151
R872 B.n452 B.n451 10.6151
R873 B.n452 B.n239 10.6151
R874 B.n462 B.n239 10.6151
R875 B.n463 B.n462 10.6151
R876 B.n464 B.n463 10.6151
R877 B.n464 B.n231 10.6151
R878 B.n474 B.n231 10.6151
R879 B.n475 B.n474 10.6151
R880 B.n476 B.n475 10.6151
R881 B.n476 B.n222 10.6151
R882 B.n486 B.n222 10.6151
R883 B.n487 B.n486 10.6151
R884 B.n489 B.n487 10.6151
R885 B.n489 B.n488 10.6151
R886 B.n488 B.n215 10.6151
R887 B.n500 B.n215 10.6151
R888 B.n501 B.n500 10.6151
R889 B.n502 B.n501 10.6151
R890 B.n503 B.n502 10.6151
R891 B.n504 B.n503 10.6151
R892 B.n507 B.n504 10.6151
R893 B.n508 B.n507 10.6151
R894 B.n509 B.n508 10.6151
R895 B.n510 B.n509 10.6151
R896 B.n512 B.n510 10.6151
R897 B.n513 B.n512 10.6151
R898 B.n514 B.n513 10.6151
R899 B.n515 B.n514 10.6151
R900 B.n517 B.n515 10.6151
R901 B.n518 B.n517 10.6151
R902 B.n519 B.n518 10.6151
R903 B.n520 B.n519 10.6151
R904 B.n522 B.n520 10.6151
R905 B.n523 B.n522 10.6151
R906 B.n524 B.n523 10.6151
R907 B.n525 B.n524 10.6151
R908 B.n527 B.n525 10.6151
R909 B.n528 B.n527 10.6151
R910 B.n529 B.n528 10.6151
R911 B.n530 B.n529 10.6151
R912 B.n531 B.n530 10.6151
R913 B.n579 B.n1 10.6151
R914 B.n579 B.n578 10.6151
R915 B.n578 B.n577 10.6151
R916 B.n577 B.n10 10.6151
R917 B.n571 B.n10 10.6151
R918 B.n571 B.n570 10.6151
R919 B.n570 B.n569 10.6151
R920 B.n569 B.n18 10.6151
R921 B.n563 B.n18 10.6151
R922 B.n563 B.n562 10.6151
R923 B.n562 B.n561 10.6151
R924 B.n561 B.n25 10.6151
R925 B.n555 B.n25 10.6151
R926 B.n555 B.n554 10.6151
R927 B.n554 B.n553 10.6151
R928 B.n553 B.n32 10.6151
R929 B.n547 B.n32 10.6151
R930 B.n547 B.n546 10.6151
R931 B.n546 B.n545 10.6151
R932 B.n545 B.n39 10.6151
R933 B.n539 B.n39 10.6151
R934 B.n539 B.n538 10.6151
R935 B.n537 B.n46 10.6151
R936 B.n88 B.n46 10.6151
R937 B.n89 B.n88 10.6151
R938 B.n92 B.n89 10.6151
R939 B.n93 B.n92 10.6151
R940 B.n96 B.n93 10.6151
R941 B.n97 B.n96 10.6151
R942 B.n100 B.n97 10.6151
R943 B.n101 B.n100 10.6151
R944 B.n104 B.n101 10.6151
R945 B.n105 B.n104 10.6151
R946 B.n108 B.n105 10.6151
R947 B.n109 B.n108 10.6151
R948 B.n112 B.n109 10.6151
R949 B.n113 B.n112 10.6151
R950 B.n116 B.n113 10.6151
R951 B.n117 B.n116 10.6151
R952 B.n120 B.n117 10.6151
R953 B.n121 B.n120 10.6151
R954 B.n124 B.n121 10.6151
R955 B.n125 B.n124 10.6151
R956 B.n128 B.n125 10.6151
R957 B.n129 B.n128 10.6151
R958 B.n132 B.n129 10.6151
R959 B.n133 B.n132 10.6151
R960 B.n136 B.n133 10.6151
R961 B.n137 B.n136 10.6151
R962 B.n140 B.n137 10.6151
R963 B.n145 B.n142 10.6151
R964 B.n146 B.n145 10.6151
R965 B.n149 B.n146 10.6151
R966 B.n150 B.n149 10.6151
R967 B.n153 B.n150 10.6151
R968 B.n154 B.n153 10.6151
R969 B.n157 B.n154 10.6151
R970 B.n158 B.n157 10.6151
R971 B.n162 B.n161 10.6151
R972 B.n165 B.n162 10.6151
R973 B.n166 B.n165 10.6151
R974 B.n169 B.n166 10.6151
R975 B.n170 B.n169 10.6151
R976 B.n173 B.n170 10.6151
R977 B.n174 B.n173 10.6151
R978 B.n177 B.n174 10.6151
R979 B.n178 B.n177 10.6151
R980 B.n181 B.n178 10.6151
R981 B.n182 B.n181 10.6151
R982 B.n185 B.n182 10.6151
R983 B.n186 B.n185 10.6151
R984 B.n189 B.n186 10.6151
R985 B.n190 B.n189 10.6151
R986 B.n193 B.n190 10.6151
R987 B.n194 B.n193 10.6151
R988 B.n197 B.n194 10.6151
R989 B.n198 B.n197 10.6151
R990 B.n201 B.n198 10.6151
R991 B.n202 B.n201 10.6151
R992 B.n205 B.n202 10.6151
R993 B.n206 B.n205 10.6151
R994 B.n209 B.n206 10.6151
R995 B.n210 B.n209 10.6151
R996 B.n213 B.n210 10.6151
R997 B.n214 B.n213 10.6151
R998 B.n532 B.n214 10.6151
R999 B.n587 B.n0 8.11757
R1000 B.n587 B.n1 8.11757
R1001 B.n374 B.n296 6.5566
R1002 B.n358 B.n357 6.5566
R1003 B.n142 B.n141 6.5566
R1004 B.n158 B.n84 6.5566
R1005 B.n225 B.t1 5.95795
R1006 B.t0 B.n574 5.95795
R1007 B.n377 B.n296 4.05904
R1008 B.n357 B.n356 4.05904
R1009 B.n141 B.n140 4.05904
R1010 B.n161 B.n84 4.05904
R1011 VN VN.t1 171.641
R1012 VN VN.t0 131.447
R1013 VDD2.n0 VDD2.t1 105.654
R1014 VDD2.n0 VDD2.t0 70.952
R1015 VDD2 VDD2.n0 0.614724
C0 VP VTAIL 1.66403f
C1 VDD2 VDD1 0.632231f
C2 VDD2 VTAIL 3.89763f
C3 VP VDD2 0.317999f
C4 VDD1 VN 0.147961f
C5 VTAIL VN 1.64979f
C6 VP VN 4.48797f
C7 VTAIL VDD1 3.84863f
C8 VDD2 VN 1.81994f
C9 VP VDD1 1.9881f
C10 VDD2 B 3.491603f
C11 VDD1 B 5.33102f
C12 VTAIL B 5.425052f
C13 VN B 7.76557f
C14 VP B 5.648177f
C15 VDD2.t1 B 1.20169f
C16 VDD2.t0 B 0.934474f
C17 VDD2.n0 B 1.68517f
C18 VN.t0 B 1.09439f
C19 VN.t1 B 1.36291f
C20 VDD1.t1 B 0.899993f
C21 VDD1.t0 B 1.175f
C22 VTAIL.t3 B 0.968658f
C23 VTAIL.n0 B 0.986609f
C24 VTAIL.t1 B 0.96866f
C25 VTAIL.n1 B 1.01114f
C26 VTAIL.t2 B 0.968658f
C27 VTAIL.n2 B 0.901542f
C28 VTAIL.t0 B 0.968658f
C29 VTAIL.n3 B 0.848123f
C30 VP.t0 B 1.36921f
C31 VP.t1 B 1.10033f
C32 VP.n0 B 1.98881f
.ends

