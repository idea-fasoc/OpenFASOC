* NGSPICE file created from diff_pair_sample_0696.ext - technology: sky130A

.subckt diff_pair_sample_0696 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t6 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=1.52625 ps=9.58 w=9.25 l=3.85
X1 VDD1.t7 VP.t0 VTAIL.t13 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=3.6075 ps=19.28 w=9.25 l=3.85
X2 VDD2.t7 VN.t1 VTAIL.t10 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=3.6075 ps=19.28 w=9.25 l=3.85
X3 VTAIL.t14 VP.t1 VDD1.t6 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X4 VTAIL.t9 VN.t2 VDD2.t5 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X5 VDD1.t5 VP.t2 VTAIL.t15 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X6 VTAIL.t8 VN.t3 VDD2.t0 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=1.52625 ps=9.58 w=9.25 l=3.85
X7 B.t11 B.t9 B.t10 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=0 ps=0 w=9.25 l=3.85
X8 VTAIL.t7 VN.t4 VDD2.t1 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X9 VDD2.t2 VN.t5 VTAIL.t6 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=3.6075 ps=19.28 w=9.25 l=3.85
X10 B.t8 B.t6 B.t7 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=0 ps=0 w=9.25 l=3.85
X11 B.t5 B.t3 B.t4 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=0 ps=0 w=9.25 l=3.85
X12 VTAIL.t12 VP.t3 VDD1.t4 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X13 VTAIL.t3 VP.t4 VDD1.t3 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=1.52625 ps=9.58 w=9.25 l=3.85
X14 VDD1.t2 VP.t5 VTAIL.t2 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X15 VDD2.t3 VN.t6 VTAIL.t5 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
X16 B.t2 B.t0 B.t1 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=0 ps=0 w=9.25 l=3.85
X17 VTAIL.t1 VP.t6 VDD1.t1 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=3.6075 pd=19.28 as=1.52625 ps=9.58 w=9.25 l=3.85
X18 VDD1.t0 VP.t7 VTAIL.t0 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=3.6075 ps=19.28 w=9.25 l=3.85
X19 VDD2.t4 VN.t7 VTAIL.t4 w_n5150_n2818# sky130_fd_pr__pfet_01v8 ad=1.52625 pd=9.58 as=1.52625 ps=9.58 w=9.25 l=3.85
R0 VN.n76 VN.n75 161.3
R1 VN.n74 VN.n40 161.3
R2 VN.n73 VN.n72 161.3
R3 VN.n71 VN.n41 161.3
R4 VN.n70 VN.n69 161.3
R5 VN.n68 VN.n42 161.3
R6 VN.n67 VN.n66 161.3
R7 VN.n65 VN.n43 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n61 VN.n44 161.3
R10 VN.n60 VN.n59 161.3
R11 VN.n58 VN.n45 161.3
R12 VN.n57 VN.n56 161.3
R13 VN.n55 VN.n46 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n47 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n37 VN.n36 161.3
R18 VN.n35 VN.n1 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n2 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n3 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n4 161.3
R25 VN.n25 VN.n24 161.3
R26 VN.n22 VN.n5 161.3
R27 VN.n21 VN.n20 161.3
R28 VN.n19 VN.n6 161.3
R29 VN.n18 VN.n17 161.3
R30 VN.n16 VN.n7 161.3
R31 VN.n15 VN.n14 161.3
R32 VN.n13 VN.n8 161.3
R33 VN.n12 VN.n11 161.3
R34 VN.n48 VN.t5 90.23
R35 VN.n9 VN.t0 90.23
R36 VN.n38 VN.n0 89.0887
R37 VN.n77 VN.n39 89.0887
R38 VN.n10 VN.n9 58.4531
R39 VN.n49 VN.n48 58.4531
R40 VN.n10 VN.t7 57.9031
R41 VN.n23 VN.t2 57.9031
R42 VN.n0 VN.t1 57.9031
R43 VN.n49 VN.t4 57.9031
R44 VN.n62 VN.t6 57.9031
R45 VN.n39 VN.t3 57.9031
R46 VN.n17 VN.n16 56.5193
R47 VN.n56 VN.n55 56.5193
R48 VN VN.n77 54.8617
R49 VN.n30 VN.n29 47.2923
R50 VN.n69 VN.n68 47.2923
R51 VN.n30 VN.n2 33.6945
R52 VN.n69 VN.n41 33.6945
R53 VN.n11 VN.n8 24.4675
R54 VN.n15 VN.n8 24.4675
R55 VN.n16 VN.n15 24.4675
R56 VN.n17 VN.n6 24.4675
R57 VN.n21 VN.n6 24.4675
R58 VN.n22 VN.n21 24.4675
R59 VN.n24 VN.n4 24.4675
R60 VN.n28 VN.n4 24.4675
R61 VN.n29 VN.n28 24.4675
R62 VN.n34 VN.n2 24.4675
R63 VN.n35 VN.n34 24.4675
R64 VN.n36 VN.n35 24.4675
R65 VN.n55 VN.n54 24.4675
R66 VN.n54 VN.n47 24.4675
R67 VN.n50 VN.n47 24.4675
R68 VN.n68 VN.n67 24.4675
R69 VN.n67 VN.n43 24.4675
R70 VN.n63 VN.n43 24.4675
R71 VN.n61 VN.n60 24.4675
R72 VN.n60 VN.n45 24.4675
R73 VN.n56 VN.n45 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n73 24.4675
R76 VN.n73 VN.n41 24.4675
R77 VN.n11 VN.n10 16.6381
R78 VN.n23 VN.n22 16.6381
R79 VN.n50 VN.n49 16.6381
R80 VN.n62 VN.n61 16.6381
R81 VN.n24 VN.n23 7.82994
R82 VN.n63 VN.n62 7.82994
R83 VN.n51 VN.n48 2.50737
R84 VN.n12 VN.n9 2.50737
R85 VN.n36 VN.n0 0.97918
R86 VN.n75 VN.n39 0.97918
R87 VN.n77 VN.n76 0.354971
R88 VN.n38 VN.n37 0.354971
R89 VN VN.n38 0.26696
R90 VN.n76 VN.n40 0.189894
R91 VN.n72 VN.n40 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n70 0.189894
R94 VN.n70 VN.n42 0.189894
R95 VN.n66 VN.n42 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n64 0.189894
R98 VN.n64 VN.n44 0.189894
R99 VN.n59 VN.n44 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n57 0.189894
R102 VN.n57 VN.n46 0.189894
R103 VN.n53 VN.n46 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n51 0.189894
R106 VN.n13 VN.n12 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n14 VN.n7 0.189894
R109 VN.n18 VN.n7 0.189894
R110 VN.n19 VN.n18 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n20 VN.n5 0.189894
R113 VN.n25 VN.n5 0.189894
R114 VN.n26 VN.n25 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n27 VN.n3 0.189894
R117 VN.n31 VN.n3 0.189894
R118 VN.n32 VN.n31 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n33 VN.n1 0.189894
R121 VN.n37 VN.n1 0.189894
R122 VDD2.n2 VDD2.n1 80.521
R123 VDD2.n2 VDD2.n0 80.521
R124 VDD2 VDD2.n5 80.5182
R125 VDD2.n4 VDD2.n3 78.7748
R126 VDD2.n4 VDD2.n2 47.9049
R127 VDD2.n5 VDD2.t1 3.51455
R128 VDD2.n5 VDD2.t2 3.51455
R129 VDD2.n3 VDD2.t0 3.51455
R130 VDD2.n3 VDD2.t3 3.51455
R131 VDD2.n1 VDD2.t5 3.51455
R132 VDD2.n1 VDD2.t7 3.51455
R133 VDD2.n0 VDD2.t6 3.51455
R134 VDD2.n0 VDD2.t4 3.51455
R135 VDD2 VDD2.n4 1.86041
R136 VTAIL.n402 VTAIL.n358 756.745
R137 VTAIL.n46 VTAIL.n2 756.745
R138 VTAIL.n96 VTAIL.n52 756.745
R139 VTAIL.n148 VTAIL.n104 756.745
R140 VTAIL.n352 VTAIL.n308 756.745
R141 VTAIL.n300 VTAIL.n256 756.745
R142 VTAIL.n250 VTAIL.n206 756.745
R143 VTAIL.n198 VTAIL.n154 756.745
R144 VTAIL.n375 VTAIL.n374 585
R145 VTAIL.n377 VTAIL.n376 585
R146 VTAIL.n370 VTAIL.n369 585
R147 VTAIL.n383 VTAIL.n382 585
R148 VTAIL.n385 VTAIL.n384 585
R149 VTAIL.n366 VTAIL.n365 585
R150 VTAIL.n392 VTAIL.n391 585
R151 VTAIL.n393 VTAIL.n364 585
R152 VTAIL.n395 VTAIL.n394 585
R153 VTAIL.n362 VTAIL.n361 585
R154 VTAIL.n401 VTAIL.n400 585
R155 VTAIL.n403 VTAIL.n402 585
R156 VTAIL.n19 VTAIL.n18 585
R157 VTAIL.n21 VTAIL.n20 585
R158 VTAIL.n14 VTAIL.n13 585
R159 VTAIL.n27 VTAIL.n26 585
R160 VTAIL.n29 VTAIL.n28 585
R161 VTAIL.n10 VTAIL.n9 585
R162 VTAIL.n36 VTAIL.n35 585
R163 VTAIL.n37 VTAIL.n8 585
R164 VTAIL.n39 VTAIL.n38 585
R165 VTAIL.n6 VTAIL.n5 585
R166 VTAIL.n45 VTAIL.n44 585
R167 VTAIL.n47 VTAIL.n46 585
R168 VTAIL.n69 VTAIL.n68 585
R169 VTAIL.n71 VTAIL.n70 585
R170 VTAIL.n64 VTAIL.n63 585
R171 VTAIL.n77 VTAIL.n76 585
R172 VTAIL.n79 VTAIL.n78 585
R173 VTAIL.n60 VTAIL.n59 585
R174 VTAIL.n86 VTAIL.n85 585
R175 VTAIL.n87 VTAIL.n58 585
R176 VTAIL.n89 VTAIL.n88 585
R177 VTAIL.n56 VTAIL.n55 585
R178 VTAIL.n95 VTAIL.n94 585
R179 VTAIL.n97 VTAIL.n96 585
R180 VTAIL.n121 VTAIL.n120 585
R181 VTAIL.n123 VTAIL.n122 585
R182 VTAIL.n116 VTAIL.n115 585
R183 VTAIL.n129 VTAIL.n128 585
R184 VTAIL.n131 VTAIL.n130 585
R185 VTAIL.n112 VTAIL.n111 585
R186 VTAIL.n138 VTAIL.n137 585
R187 VTAIL.n139 VTAIL.n110 585
R188 VTAIL.n141 VTAIL.n140 585
R189 VTAIL.n108 VTAIL.n107 585
R190 VTAIL.n147 VTAIL.n146 585
R191 VTAIL.n149 VTAIL.n148 585
R192 VTAIL.n353 VTAIL.n352 585
R193 VTAIL.n351 VTAIL.n350 585
R194 VTAIL.n312 VTAIL.n311 585
R195 VTAIL.n316 VTAIL.n314 585
R196 VTAIL.n345 VTAIL.n344 585
R197 VTAIL.n343 VTAIL.n342 585
R198 VTAIL.n318 VTAIL.n317 585
R199 VTAIL.n337 VTAIL.n336 585
R200 VTAIL.n335 VTAIL.n334 585
R201 VTAIL.n322 VTAIL.n321 585
R202 VTAIL.n329 VTAIL.n328 585
R203 VTAIL.n327 VTAIL.n326 585
R204 VTAIL.n301 VTAIL.n300 585
R205 VTAIL.n299 VTAIL.n298 585
R206 VTAIL.n260 VTAIL.n259 585
R207 VTAIL.n264 VTAIL.n262 585
R208 VTAIL.n293 VTAIL.n292 585
R209 VTAIL.n291 VTAIL.n290 585
R210 VTAIL.n266 VTAIL.n265 585
R211 VTAIL.n285 VTAIL.n284 585
R212 VTAIL.n283 VTAIL.n282 585
R213 VTAIL.n270 VTAIL.n269 585
R214 VTAIL.n277 VTAIL.n276 585
R215 VTAIL.n275 VTAIL.n274 585
R216 VTAIL.n251 VTAIL.n250 585
R217 VTAIL.n249 VTAIL.n248 585
R218 VTAIL.n210 VTAIL.n209 585
R219 VTAIL.n214 VTAIL.n212 585
R220 VTAIL.n243 VTAIL.n242 585
R221 VTAIL.n241 VTAIL.n240 585
R222 VTAIL.n216 VTAIL.n215 585
R223 VTAIL.n235 VTAIL.n234 585
R224 VTAIL.n233 VTAIL.n232 585
R225 VTAIL.n220 VTAIL.n219 585
R226 VTAIL.n227 VTAIL.n226 585
R227 VTAIL.n225 VTAIL.n224 585
R228 VTAIL.n199 VTAIL.n198 585
R229 VTAIL.n197 VTAIL.n196 585
R230 VTAIL.n158 VTAIL.n157 585
R231 VTAIL.n162 VTAIL.n160 585
R232 VTAIL.n191 VTAIL.n190 585
R233 VTAIL.n189 VTAIL.n188 585
R234 VTAIL.n164 VTAIL.n163 585
R235 VTAIL.n183 VTAIL.n182 585
R236 VTAIL.n181 VTAIL.n180 585
R237 VTAIL.n168 VTAIL.n167 585
R238 VTAIL.n175 VTAIL.n174 585
R239 VTAIL.n173 VTAIL.n172 585
R240 VTAIL.n373 VTAIL.t10 329.038
R241 VTAIL.n17 VTAIL.t11 329.038
R242 VTAIL.n67 VTAIL.t0 329.038
R243 VTAIL.n119 VTAIL.t3 329.038
R244 VTAIL.n325 VTAIL.t13 329.038
R245 VTAIL.n273 VTAIL.t1 329.038
R246 VTAIL.n223 VTAIL.t6 329.038
R247 VTAIL.n171 VTAIL.t8 329.038
R248 VTAIL.n376 VTAIL.n375 171.744
R249 VTAIL.n376 VTAIL.n369 171.744
R250 VTAIL.n383 VTAIL.n369 171.744
R251 VTAIL.n384 VTAIL.n383 171.744
R252 VTAIL.n384 VTAIL.n365 171.744
R253 VTAIL.n392 VTAIL.n365 171.744
R254 VTAIL.n393 VTAIL.n392 171.744
R255 VTAIL.n394 VTAIL.n393 171.744
R256 VTAIL.n394 VTAIL.n361 171.744
R257 VTAIL.n401 VTAIL.n361 171.744
R258 VTAIL.n402 VTAIL.n401 171.744
R259 VTAIL.n20 VTAIL.n19 171.744
R260 VTAIL.n20 VTAIL.n13 171.744
R261 VTAIL.n27 VTAIL.n13 171.744
R262 VTAIL.n28 VTAIL.n27 171.744
R263 VTAIL.n28 VTAIL.n9 171.744
R264 VTAIL.n36 VTAIL.n9 171.744
R265 VTAIL.n37 VTAIL.n36 171.744
R266 VTAIL.n38 VTAIL.n37 171.744
R267 VTAIL.n38 VTAIL.n5 171.744
R268 VTAIL.n45 VTAIL.n5 171.744
R269 VTAIL.n46 VTAIL.n45 171.744
R270 VTAIL.n70 VTAIL.n69 171.744
R271 VTAIL.n70 VTAIL.n63 171.744
R272 VTAIL.n77 VTAIL.n63 171.744
R273 VTAIL.n78 VTAIL.n77 171.744
R274 VTAIL.n78 VTAIL.n59 171.744
R275 VTAIL.n86 VTAIL.n59 171.744
R276 VTAIL.n87 VTAIL.n86 171.744
R277 VTAIL.n88 VTAIL.n87 171.744
R278 VTAIL.n88 VTAIL.n55 171.744
R279 VTAIL.n95 VTAIL.n55 171.744
R280 VTAIL.n96 VTAIL.n95 171.744
R281 VTAIL.n122 VTAIL.n121 171.744
R282 VTAIL.n122 VTAIL.n115 171.744
R283 VTAIL.n129 VTAIL.n115 171.744
R284 VTAIL.n130 VTAIL.n129 171.744
R285 VTAIL.n130 VTAIL.n111 171.744
R286 VTAIL.n138 VTAIL.n111 171.744
R287 VTAIL.n139 VTAIL.n138 171.744
R288 VTAIL.n140 VTAIL.n139 171.744
R289 VTAIL.n140 VTAIL.n107 171.744
R290 VTAIL.n147 VTAIL.n107 171.744
R291 VTAIL.n148 VTAIL.n147 171.744
R292 VTAIL.n352 VTAIL.n351 171.744
R293 VTAIL.n351 VTAIL.n311 171.744
R294 VTAIL.n316 VTAIL.n311 171.744
R295 VTAIL.n344 VTAIL.n316 171.744
R296 VTAIL.n344 VTAIL.n343 171.744
R297 VTAIL.n343 VTAIL.n317 171.744
R298 VTAIL.n336 VTAIL.n317 171.744
R299 VTAIL.n336 VTAIL.n335 171.744
R300 VTAIL.n335 VTAIL.n321 171.744
R301 VTAIL.n328 VTAIL.n321 171.744
R302 VTAIL.n328 VTAIL.n327 171.744
R303 VTAIL.n300 VTAIL.n299 171.744
R304 VTAIL.n299 VTAIL.n259 171.744
R305 VTAIL.n264 VTAIL.n259 171.744
R306 VTAIL.n292 VTAIL.n264 171.744
R307 VTAIL.n292 VTAIL.n291 171.744
R308 VTAIL.n291 VTAIL.n265 171.744
R309 VTAIL.n284 VTAIL.n265 171.744
R310 VTAIL.n284 VTAIL.n283 171.744
R311 VTAIL.n283 VTAIL.n269 171.744
R312 VTAIL.n276 VTAIL.n269 171.744
R313 VTAIL.n276 VTAIL.n275 171.744
R314 VTAIL.n250 VTAIL.n249 171.744
R315 VTAIL.n249 VTAIL.n209 171.744
R316 VTAIL.n214 VTAIL.n209 171.744
R317 VTAIL.n242 VTAIL.n214 171.744
R318 VTAIL.n242 VTAIL.n241 171.744
R319 VTAIL.n241 VTAIL.n215 171.744
R320 VTAIL.n234 VTAIL.n215 171.744
R321 VTAIL.n234 VTAIL.n233 171.744
R322 VTAIL.n233 VTAIL.n219 171.744
R323 VTAIL.n226 VTAIL.n219 171.744
R324 VTAIL.n226 VTAIL.n225 171.744
R325 VTAIL.n198 VTAIL.n197 171.744
R326 VTAIL.n197 VTAIL.n157 171.744
R327 VTAIL.n162 VTAIL.n157 171.744
R328 VTAIL.n190 VTAIL.n162 171.744
R329 VTAIL.n190 VTAIL.n189 171.744
R330 VTAIL.n189 VTAIL.n163 171.744
R331 VTAIL.n182 VTAIL.n163 171.744
R332 VTAIL.n182 VTAIL.n181 171.744
R333 VTAIL.n181 VTAIL.n167 171.744
R334 VTAIL.n174 VTAIL.n167 171.744
R335 VTAIL.n174 VTAIL.n173 171.744
R336 VTAIL.n375 VTAIL.t10 85.8723
R337 VTAIL.n19 VTAIL.t11 85.8723
R338 VTAIL.n69 VTAIL.t0 85.8723
R339 VTAIL.n121 VTAIL.t3 85.8723
R340 VTAIL.n327 VTAIL.t13 85.8723
R341 VTAIL.n275 VTAIL.t1 85.8723
R342 VTAIL.n225 VTAIL.t6 85.8723
R343 VTAIL.n173 VTAIL.t8 85.8723
R344 VTAIL.n307 VTAIL.n306 62.096
R345 VTAIL.n205 VTAIL.n204 62.096
R346 VTAIL.n1 VTAIL.n0 62.0959
R347 VTAIL.n103 VTAIL.n102 62.0959
R348 VTAIL.n407 VTAIL.n406 32.3793
R349 VTAIL.n51 VTAIL.n50 32.3793
R350 VTAIL.n101 VTAIL.n100 32.3793
R351 VTAIL.n153 VTAIL.n152 32.3793
R352 VTAIL.n357 VTAIL.n356 32.3793
R353 VTAIL.n305 VTAIL.n304 32.3793
R354 VTAIL.n255 VTAIL.n254 32.3793
R355 VTAIL.n203 VTAIL.n202 32.3793
R356 VTAIL.n407 VTAIL.n357 23.9445
R357 VTAIL.n203 VTAIL.n153 23.9445
R358 VTAIL.n395 VTAIL.n362 13.1884
R359 VTAIL.n39 VTAIL.n6 13.1884
R360 VTAIL.n89 VTAIL.n56 13.1884
R361 VTAIL.n141 VTAIL.n108 13.1884
R362 VTAIL.n314 VTAIL.n312 13.1884
R363 VTAIL.n262 VTAIL.n260 13.1884
R364 VTAIL.n212 VTAIL.n210 13.1884
R365 VTAIL.n160 VTAIL.n158 13.1884
R366 VTAIL.n396 VTAIL.n364 12.8005
R367 VTAIL.n400 VTAIL.n399 12.8005
R368 VTAIL.n40 VTAIL.n8 12.8005
R369 VTAIL.n44 VTAIL.n43 12.8005
R370 VTAIL.n90 VTAIL.n58 12.8005
R371 VTAIL.n94 VTAIL.n93 12.8005
R372 VTAIL.n142 VTAIL.n110 12.8005
R373 VTAIL.n146 VTAIL.n145 12.8005
R374 VTAIL.n350 VTAIL.n349 12.8005
R375 VTAIL.n346 VTAIL.n345 12.8005
R376 VTAIL.n298 VTAIL.n297 12.8005
R377 VTAIL.n294 VTAIL.n293 12.8005
R378 VTAIL.n248 VTAIL.n247 12.8005
R379 VTAIL.n244 VTAIL.n243 12.8005
R380 VTAIL.n196 VTAIL.n195 12.8005
R381 VTAIL.n192 VTAIL.n191 12.8005
R382 VTAIL.n391 VTAIL.n390 12.0247
R383 VTAIL.n403 VTAIL.n360 12.0247
R384 VTAIL.n35 VTAIL.n34 12.0247
R385 VTAIL.n47 VTAIL.n4 12.0247
R386 VTAIL.n85 VTAIL.n84 12.0247
R387 VTAIL.n97 VTAIL.n54 12.0247
R388 VTAIL.n137 VTAIL.n136 12.0247
R389 VTAIL.n149 VTAIL.n106 12.0247
R390 VTAIL.n353 VTAIL.n310 12.0247
R391 VTAIL.n342 VTAIL.n315 12.0247
R392 VTAIL.n301 VTAIL.n258 12.0247
R393 VTAIL.n290 VTAIL.n263 12.0247
R394 VTAIL.n251 VTAIL.n208 12.0247
R395 VTAIL.n240 VTAIL.n213 12.0247
R396 VTAIL.n199 VTAIL.n156 12.0247
R397 VTAIL.n188 VTAIL.n161 12.0247
R398 VTAIL.n389 VTAIL.n366 11.249
R399 VTAIL.n404 VTAIL.n358 11.249
R400 VTAIL.n33 VTAIL.n10 11.249
R401 VTAIL.n48 VTAIL.n2 11.249
R402 VTAIL.n83 VTAIL.n60 11.249
R403 VTAIL.n98 VTAIL.n52 11.249
R404 VTAIL.n135 VTAIL.n112 11.249
R405 VTAIL.n150 VTAIL.n104 11.249
R406 VTAIL.n354 VTAIL.n308 11.249
R407 VTAIL.n341 VTAIL.n318 11.249
R408 VTAIL.n302 VTAIL.n256 11.249
R409 VTAIL.n289 VTAIL.n266 11.249
R410 VTAIL.n252 VTAIL.n206 11.249
R411 VTAIL.n239 VTAIL.n216 11.249
R412 VTAIL.n200 VTAIL.n154 11.249
R413 VTAIL.n187 VTAIL.n164 11.249
R414 VTAIL.n374 VTAIL.n373 10.7239
R415 VTAIL.n18 VTAIL.n17 10.7239
R416 VTAIL.n68 VTAIL.n67 10.7239
R417 VTAIL.n120 VTAIL.n119 10.7239
R418 VTAIL.n326 VTAIL.n325 10.7239
R419 VTAIL.n274 VTAIL.n273 10.7239
R420 VTAIL.n224 VTAIL.n223 10.7239
R421 VTAIL.n172 VTAIL.n171 10.7239
R422 VTAIL.n386 VTAIL.n385 10.4732
R423 VTAIL.n30 VTAIL.n29 10.4732
R424 VTAIL.n80 VTAIL.n79 10.4732
R425 VTAIL.n132 VTAIL.n131 10.4732
R426 VTAIL.n338 VTAIL.n337 10.4732
R427 VTAIL.n286 VTAIL.n285 10.4732
R428 VTAIL.n236 VTAIL.n235 10.4732
R429 VTAIL.n184 VTAIL.n183 10.4732
R430 VTAIL.n382 VTAIL.n368 9.69747
R431 VTAIL.n26 VTAIL.n12 9.69747
R432 VTAIL.n76 VTAIL.n62 9.69747
R433 VTAIL.n128 VTAIL.n114 9.69747
R434 VTAIL.n334 VTAIL.n320 9.69747
R435 VTAIL.n282 VTAIL.n268 9.69747
R436 VTAIL.n232 VTAIL.n218 9.69747
R437 VTAIL.n180 VTAIL.n166 9.69747
R438 VTAIL.n406 VTAIL.n405 9.45567
R439 VTAIL.n50 VTAIL.n49 9.45567
R440 VTAIL.n100 VTAIL.n99 9.45567
R441 VTAIL.n152 VTAIL.n151 9.45567
R442 VTAIL.n356 VTAIL.n355 9.45567
R443 VTAIL.n304 VTAIL.n303 9.45567
R444 VTAIL.n254 VTAIL.n253 9.45567
R445 VTAIL.n202 VTAIL.n201 9.45567
R446 VTAIL.n405 VTAIL.n404 9.3005
R447 VTAIL.n360 VTAIL.n359 9.3005
R448 VTAIL.n399 VTAIL.n398 9.3005
R449 VTAIL.n372 VTAIL.n371 9.3005
R450 VTAIL.n379 VTAIL.n378 9.3005
R451 VTAIL.n381 VTAIL.n380 9.3005
R452 VTAIL.n368 VTAIL.n367 9.3005
R453 VTAIL.n387 VTAIL.n386 9.3005
R454 VTAIL.n389 VTAIL.n388 9.3005
R455 VTAIL.n390 VTAIL.n363 9.3005
R456 VTAIL.n397 VTAIL.n396 9.3005
R457 VTAIL.n49 VTAIL.n48 9.3005
R458 VTAIL.n4 VTAIL.n3 9.3005
R459 VTAIL.n43 VTAIL.n42 9.3005
R460 VTAIL.n16 VTAIL.n15 9.3005
R461 VTAIL.n23 VTAIL.n22 9.3005
R462 VTAIL.n25 VTAIL.n24 9.3005
R463 VTAIL.n12 VTAIL.n11 9.3005
R464 VTAIL.n31 VTAIL.n30 9.3005
R465 VTAIL.n33 VTAIL.n32 9.3005
R466 VTAIL.n34 VTAIL.n7 9.3005
R467 VTAIL.n41 VTAIL.n40 9.3005
R468 VTAIL.n99 VTAIL.n98 9.3005
R469 VTAIL.n54 VTAIL.n53 9.3005
R470 VTAIL.n93 VTAIL.n92 9.3005
R471 VTAIL.n66 VTAIL.n65 9.3005
R472 VTAIL.n73 VTAIL.n72 9.3005
R473 VTAIL.n75 VTAIL.n74 9.3005
R474 VTAIL.n62 VTAIL.n61 9.3005
R475 VTAIL.n81 VTAIL.n80 9.3005
R476 VTAIL.n83 VTAIL.n82 9.3005
R477 VTAIL.n84 VTAIL.n57 9.3005
R478 VTAIL.n91 VTAIL.n90 9.3005
R479 VTAIL.n151 VTAIL.n150 9.3005
R480 VTAIL.n106 VTAIL.n105 9.3005
R481 VTAIL.n145 VTAIL.n144 9.3005
R482 VTAIL.n118 VTAIL.n117 9.3005
R483 VTAIL.n125 VTAIL.n124 9.3005
R484 VTAIL.n127 VTAIL.n126 9.3005
R485 VTAIL.n114 VTAIL.n113 9.3005
R486 VTAIL.n133 VTAIL.n132 9.3005
R487 VTAIL.n135 VTAIL.n134 9.3005
R488 VTAIL.n136 VTAIL.n109 9.3005
R489 VTAIL.n143 VTAIL.n142 9.3005
R490 VTAIL.n324 VTAIL.n323 9.3005
R491 VTAIL.n331 VTAIL.n330 9.3005
R492 VTAIL.n333 VTAIL.n332 9.3005
R493 VTAIL.n320 VTAIL.n319 9.3005
R494 VTAIL.n339 VTAIL.n338 9.3005
R495 VTAIL.n341 VTAIL.n340 9.3005
R496 VTAIL.n315 VTAIL.n313 9.3005
R497 VTAIL.n347 VTAIL.n346 9.3005
R498 VTAIL.n355 VTAIL.n354 9.3005
R499 VTAIL.n310 VTAIL.n309 9.3005
R500 VTAIL.n349 VTAIL.n348 9.3005
R501 VTAIL.n272 VTAIL.n271 9.3005
R502 VTAIL.n279 VTAIL.n278 9.3005
R503 VTAIL.n281 VTAIL.n280 9.3005
R504 VTAIL.n268 VTAIL.n267 9.3005
R505 VTAIL.n287 VTAIL.n286 9.3005
R506 VTAIL.n289 VTAIL.n288 9.3005
R507 VTAIL.n263 VTAIL.n261 9.3005
R508 VTAIL.n295 VTAIL.n294 9.3005
R509 VTAIL.n303 VTAIL.n302 9.3005
R510 VTAIL.n258 VTAIL.n257 9.3005
R511 VTAIL.n297 VTAIL.n296 9.3005
R512 VTAIL.n222 VTAIL.n221 9.3005
R513 VTAIL.n229 VTAIL.n228 9.3005
R514 VTAIL.n231 VTAIL.n230 9.3005
R515 VTAIL.n218 VTAIL.n217 9.3005
R516 VTAIL.n237 VTAIL.n236 9.3005
R517 VTAIL.n239 VTAIL.n238 9.3005
R518 VTAIL.n213 VTAIL.n211 9.3005
R519 VTAIL.n245 VTAIL.n244 9.3005
R520 VTAIL.n253 VTAIL.n252 9.3005
R521 VTAIL.n208 VTAIL.n207 9.3005
R522 VTAIL.n247 VTAIL.n246 9.3005
R523 VTAIL.n170 VTAIL.n169 9.3005
R524 VTAIL.n177 VTAIL.n176 9.3005
R525 VTAIL.n179 VTAIL.n178 9.3005
R526 VTAIL.n166 VTAIL.n165 9.3005
R527 VTAIL.n185 VTAIL.n184 9.3005
R528 VTAIL.n187 VTAIL.n186 9.3005
R529 VTAIL.n161 VTAIL.n159 9.3005
R530 VTAIL.n193 VTAIL.n192 9.3005
R531 VTAIL.n201 VTAIL.n200 9.3005
R532 VTAIL.n156 VTAIL.n155 9.3005
R533 VTAIL.n195 VTAIL.n194 9.3005
R534 VTAIL.n381 VTAIL.n370 8.92171
R535 VTAIL.n25 VTAIL.n14 8.92171
R536 VTAIL.n75 VTAIL.n64 8.92171
R537 VTAIL.n127 VTAIL.n116 8.92171
R538 VTAIL.n333 VTAIL.n322 8.92171
R539 VTAIL.n281 VTAIL.n270 8.92171
R540 VTAIL.n231 VTAIL.n220 8.92171
R541 VTAIL.n179 VTAIL.n168 8.92171
R542 VTAIL.n378 VTAIL.n377 8.14595
R543 VTAIL.n22 VTAIL.n21 8.14595
R544 VTAIL.n72 VTAIL.n71 8.14595
R545 VTAIL.n124 VTAIL.n123 8.14595
R546 VTAIL.n330 VTAIL.n329 8.14595
R547 VTAIL.n278 VTAIL.n277 8.14595
R548 VTAIL.n228 VTAIL.n227 8.14595
R549 VTAIL.n176 VTAIL.n175 8.14595
R550 VTAIL.n374 VTAIL.n372 7.3702
R551 VTAIL.n18 VTAIL.n16 7.3702
R552 VTAIL.n68 VTAIL.n66 7.3702
R553 VTAIL.n120 VTAIL.n118 7.3702
R554 VTAIL.n326 VTAIL.n324 7.3702
R555 VTAIL.n274 VTAIL.n272 7.3702
R556 VTAIL.n224 VTAIL.n222 7.3702
R557 VTAIL.n172 VTAIL.n170 7.3702
R558 VTAIL.n377 VTAIL.n372 5.81868
R559 VTAIL.n21 VTAIL.n16 5.81868
R560 VTAIL.n71 VTAIL.n66 5.81868
R561 VTAIL.n123 VTAIL.n118 5.81868
R562 VTAIL.n329 VTAIL.n324 5.81868
R563 VTAIL.n277 VTAIL.n272 5.81868
R564 VTAIL.n227 VTAIL.n222 5.81868
R565 VTAIL.n175 VTAIL.n170 5.81868
R566 VTAIL.n378 VTAIL.n370 5.04292
R567 VTAIL.n22 VTAIL.n14 5.04292
R568 VTAIL.n72 VTAIL.n64 5.04292
R569 VTAIL.n124 VTAIL.n116 5.04292
R570 VTAIL.n330 VTAIL.n322 5.04292
R571 VTAIL.n278 VTAIL.n270 5.04292
R572 VTAIL.n228 VTAIL.n220 5.04292
R573 VTAIL.n176 VTAIL.n168 5.04292
R574 VTAIL.n382 VTAIL.n381 4.26717
R575 VTAIL.n26 VTAIL.n25 4.26717
R576 VTAIL.n76 VTAIL.n75 4.26717
R577 VTAIL.n128 VTAIL.n127 4.26717
R578 VTAIL.n334 VTAIL.n333 4.26717
R579 VTAIL.n282 VTAIL.n281 4.26717
R580 VTAIL.n232 VTAIL.n231 4.26717
R581 VTAIL.n180 VTAIL.n179 4.26717
R582 VTAIL.n205 VTAIL.n203 3.60395
R583 VTAIL.n255 VTAIL.n205 3.60395
R584 VTAIL.n307 VTAIL.n305 3.60395
R585 VTAIL.n357 VTAIL.n307 3.60395
R586 VTAIL.n153 VTAIL.n103 3.60395
R587 VTAIL.n103 VTAIL.n101 3.60395
R588 VTAIL.n51 VTAIL.n1 3.60395
R589 VTAIL VTAIL.n407 3.54576
R590 VTAIL.n0 VTAIL.t4 3.51455
R591 VTAIL.n0 VTAIL.t9 3.51455
R592 VTAIL.n102 VTAIL.t15 3.51455
R593 VTAIL.n102 VTAIL.t12 3.51455
R594 VTAIL.n306 VTAIL.t2 3.51455
R595 VTAIL.n306 VTAIL.t14 3.51455
R596 VTAIL.n204 VTAIL.t5 3.51455
R597 VTAIL.n204 VTAIL.t7 3.51455
R598 VTAIL.n385 VTAIL.n368 3.49141
R599 VTAIL.n29 VTAIL.n12 3.49141
R600 VTAIL.n79 VTAIL.n62 3.49141
R601 VTAIL.n131 VTAIL.n114 3.49141
R602 VTAIL.n337 VTAIL.n320 3.49141
R603 VTAIL.n285 VTAIL.n268 3.49141
R604 VTAIL.n235 VTAIL.n218 3.49141
R605 VTAIL.n183 VTAIL.n166 3.49141
R606 VTAIL.n386 VTAIL.n366 2.71565
R607 VTAIL.n406 VTAIL.n358 2.71565
R608 VTAIL.n30 VTAIL.n10 2.71565
R609 VTAIL.n50 VTAIL.n2 2.71565
R610 VTAIL.n80 VTAIL.n60 2.71565
R611 VTAIL.n100 VTAIL.n52 2.71565
R612 VTAIL.n132 VTAIL.n112 2.71565
R613 VTAIL.n152 VTAIL.n104 2.71565
R614 VTAIL.n356 VTAIL.n308 2.71565
R615 VTAIL.n338 VTAIL.n318 2.71565
R616 VTAIL.n304 VTAIL.n256 2.71565
R617 VTAIL.n286 VTAIL.n266 2.71565
R618 VTAIL.n254 VTAIL.n206 2.71565
R619 VTAIL.n236 VTAIL.n216 2.71565
R620 VTAIL.n202 VTAIL.n154 2.71565
R621 VTAIL.n184 VTAIL.n164 2.71565
R622 VTAIL.n373 VTAIL.n371 2.41283
R623 VTAIL.n17 VTAIL.n15 2.41283
R624 VTAIL.n67 VTAIL.n65 2.41283
R625 VTAIL.n119 VTAIL.n117 2.41283
R626 VTAIL.n325 VTAIL.n323 2.41283
R627 VTAIL.n273 VTAIL.n271 2.41283
R628 VTAIL.n223 VTAIL.n221 2.41283
R629 VTAIL.n171 VTAIL.n169 2.41283
R630 VTAIL.n391 VTAIL.n389 1.93989
R631 VTAIL.n404 VTAIL.n403 1.93989
R632 VTAIL.n35 VTAIL.n33 1.93989
R633 VTAIL.n48 VTAIL.n47 1.93989
R634 VTAIL.n85 VTAIL.n83 1.93989
R635 VTAIL.n98 VTAIL.n97 1.93989
R636 VTAIL.n137 VTAIL.n135 1.93989
R637 VTAIL.n150 VTAIL.n149 1.93989
R638 VTAIL.n354 VTAIL.n353 1.93989
R639 VTAIL.n342 VTAIL.n341 1.93989
R640 VTAIL.n302 VTAIL.n301 1.93989
R641 VTAIL.n290 VTAIL.n289 1.93989
R642 VTAIL.n252 VTAIL.n251 1.93989
R643 VTAIL.n240 VTAIL.n239 1.93989
R644 VTAIL.n200 VTAIL.n199 1.93989
R645 VTAIL.n188 VTAIL.n187 1.93989
R646 VTAIL.n390 VTAIL.n364 1.16414
R647 VTAIL.n400 VTAIL.n360 1.16414
R648 VTAIL.n34 VTAIL.n8 1.16414
R649 VTAIL.n44 VTAIL.n4 1.16414
R650 VTAIL.n84 VTAIL.n58 1.16414
R651 VTAIL.n94 VTAIL.n54 1.16414
R652 VTAIL.n136 VTAIL.n110 1.16414
R653 VTAIL.n146 VTAIL.n106 1.16414
R654 VTAIL.n350 VTAIL.n310 1.16414
R655 VTAIL.n345 VTAIL.n315 1.16414
R656 VTAIL.n298 VTAIL.n258 1.16414
R657 VTAIL.n293 VTAIL.n263 1.16414
R658 VTAIL.n248 VTAIL.n208 1.16414
R659 VTAIL.n243 VTAIL.n213 1.16414
R660 VTAIL.n196 VTAIL.n156 1.16414
R661 VTAIL.n191 VTAIL.n161 1.16414
R662 VTAIL.n305 VTAIL.n255 0.470328
R663 VTAIL.n101 VTAIL.n51 0.470328
R664 VTAIL.n396 VTAIL.n395 0.388379
R665 VTAIL.n399 VTAIL.n362 0.388379
R666 VTAIL.n40 VTAIL.n39 0.388379
R667 VTAIL.n43 VTAIL.n6 0.388379
R668 VTAIL.n90 VTAIL.n89 0.388379
R669 VTAIL.n93 VTAIL.n56 0.388379
R670 VTAIL.n142 VTAIL.n141 0.388379
R671 VTAIL.n145 VTAIL.n108 0.388379
R672 VTAIL.n349 VTAIL.n312 0.388379
R673 VTAIL.n346 VTAIL.n314 0.388379
R674 VTAIL.n297 VTAIL.n260 0.388379
R675 VTAIL.n294 VTAIL.n262 0.388379
R676 VTAIL.n247 VTAIL.n210 0.388379
R677 VTAIL.n244 VTAIL.n212 0.388379
R678 VTAIL.n195 VTAIL.n158 0.388379
R679 VTAIL.n192 VTAIL.n160 0.388379
R680 VTAIL.n379 VTAIL.n371 0.155672
R681 VTAIL.n380 VTAIL.n379 0.155672
R682 VTAIL.n380 VTAIL.n367 0.155672
R683 VTAIL.n387 VTAIL.n367 0.155672
R684 VTAIL.n388 VTAIL.n387 0.155672
R685 VTAIL.n388 VTAIL.n363 0.155672
R686 VTAIL.n397 VTAIL.n363 0.155672
R687 VTAIL.n398 VTAIL.n397 0.155672
R688 VTAIL.n398 VTAIL.n359 0.155672
R689 VTAIL.n405 VTAIL.n359 0.155672
R690 VTAIL.n23 VTAIL.n15 0.155672
R691 VTAIL.n24 VTAIL.n23 0.155672
R692 VTAIL.n24 VTAIL.n11 0.155672
R693 VTAIL.n31 VTAIL.n11 0.155672
R694 VTAIL.n32 VTAIL.n31 0.155672
R695 VTAIL.n32 VTAIL.n7 0.155672
R696 VTAIL.n41 VTAIL.n7 0.155672
R697 VTAIL.n42 VTAIL.n41 0.155672
R698 VTAIL.n42 VTAIL.n3 0.155672
R699 VTAIL.n49 VTAIL.n3 0.155672
R700 VTAIL.n73 VTAIL.n65 0.155672
R701 VTAIL.n74 VTAIL.n73 0.155672
R702 VTAIL.n74 VTAIL.n61 0.155672
R703 VTAIL.n81 VTAIL.n61 0.155672
R704 VTAIL.n82 VTAIL.n81 0.155672
R705 VTAIL.n82 VTAIL.n57 0.155672
R706 VTAIL.n91 VTAIL.n57 0.155672
R707 VTAIL.n92 VTAIL.n91 0.155672
R708 VTAIL.n92 VTAIL.n53 0.155672
R709 VTAIL.n99 VTAIL.n53 0.155672
R710 VTAIL.n125 VTAIL.n117 0.155672
R711 VTAIL.n126 VTAIL.n125 0.155672
R712 VTAIL.n126 VTAIL.n113 0.155672
R713 VTAIL.n133 VTAIL.n113 0.155672
R714 VTAIL.n134 VTAIL.n133 0.155672
R715 VTAIL.n134 VTAIL.n109 0.155672
R716 VTAIL.n143 VTAIL.n109 0.155672
R717 VTAIL.n144 VTAIL.n143 0.155672
R718 VTAIL.n144 VTAIL.n105 0.155672
R719 VTAIL.n151 VTAIL.n105 0.155672
R720 VTAIL.n355 VTAIL.n309 0.155672
R721 VTAIL.n348 VTAIL.n309 0.155672
R722 VTAIL.n348 VTAIL.n347 0.155672
R723 VTAIL.n347 VTAIL.n313 0.155672
R724 VTAIL.n340 VTAIL.n313 0.155672
R725 VTAIL.n340 VTAIL.n339 0.155672
R726 VTAIL.n339 VTAIL.n319 0.155672
R727 VTAIL.n332 VTAIL.n319 0.155672
R728 VTAIL.n332 VTAIL.n331 0.155672
R729 VTAIL.n331 VTAIL.n323 0.155672
R730 VTAIL.n303 VTAIL.n257 0.155672
R731 VTAIL.n296 VTAIL.n257 0.155672
R732 VTAIL.n296 VTAIL.n295 0.155672
R733 VTAIL.n295 VTAIL.n261 0.155672
R734 VTAIL.n288 VTAIL.n261 0.155672
R735 VTAIL.n288 VTAIL.n287 0.155672
R736 VTAIL.n287 VTAIL.n267 0.155672
R737 VTAIL.n280 VTAIL.n267 0.155672
R738 VTAIL.n280 VTAIL.n279 0.155672
R739 VTAIL.n279 VTAIL.n271 0.155672
R740 VTAIL.n253 VTAIL.n207 0.155672
R741 VTAIL.n246 VTAIL.n207 0.155672
R742 VTAIL.n246 VTAIL.n245 0.155672
R743 VTAIL.n245 VTAIL.n211 0.155672
R744 VTAIL.n238 VTAIL.n211 0.155672
R745 VTAIL.n238 VTAIL.n237 0.155672
R746 VTAIL.n237 VTAIL.n217 0.155672
R747 VTAIL.n230 VTAIL.n217 0.155672
R748 VTAIL.n230 VTAIL.n229 0.155672
R749 VTAIL.n229 VTAIL.n221 0.155672
R750 VTAIL.n201 VTAIL.n155 0.155672
R751 VTAIL.n194 VTAIL.n155 0.155672
R752 VTAIL.n194 VTAIL.n193 0.155672
R753 VTAIL.n193 VTAIL.n159 0.155672
R754 VTAIL.n186 VTAIL.n159 0.155672
R755 VTAIL.n186 VTAIL.n185 0.155672
R756 VTAIL.n185 VTAIL.n165 0.155672
R757 VTAIL.n178 VTAIL.n165 0.155672
R758 VTAIL.n178 VTAIL.n177 0.155672
R759 VTAIL.n177 VTAIL.n169 0.155672
R760 VTAIL VTAIL.n1 0.0586897
R761 VP.n26 VP.n25 161.3
R762 VP.n27 VP.n22 161.3
R763 VP.n29 VP.n28 161.3
R764 VP.n30 VP.n21 161.3
R765 VP.n32 VP.n31 161.3
R766 VP.n33 VP.n20 161.3
R767 VP.n35 VP.n34 161.3
R768 VP.n36 VP.n19 161.3
R769 VP.n39 VP.n38 161.3
R770 VP.n40 VP.n18 161.3
R771 VP.n42 VP.n41 161.3
R772 VP.n43 VP.n17 161.3
R773 VP.n45 VP.n44 161.3
R774 VP.n46 VP.n16 161.3
R775 VP.n48 VP.n47 161.3
R776 VP.n49 VP.n15 161.3
R777 VP.n51 VP.n50 161.3
R778 VP.n95 VP.n94 161.3
R779 VP.n93 VP.n1 161.3
R780 VP.n92 VP.n91 161.3
R781 VP.n90 VP.n2 161.3
R782 VP.n89 VP.n88 161.3
R783 VP.n87 VP.n3 161.3
R784 VP.n86 VP.n85 161.3
R785 VP.n84 VP.n4 161.3
R786 VP.n83 VP.n82 161.3
R787 VP.n80 VP.n5 161.3
R788 VP.n79 VP.n78 161.3
R789 VP.n77 VP.n6 161.3
R790 VP.n76 VP.n75 161.3
R791 VP.n74 VP.n7 161.3
R792 VP.n73 VP.n72 161.3
R793 VP.n71 VP.n8 161.3
R794 VP.n70 VP.n69 161.3
R795 VP.n67 VP.n9 161.3
R796 VP.n66 VP.n65 161.3
R797 VP.n64 VP.n10 161.3
R798 VP.n63 VP.n62 161.3
R799 VP.n61 VP.n11 161.3
R800 VP.n60 VP.n59 161.3
R801 VP.n58 VP.n12 161.3
R802 VP.n57 VP.n56 161.3
R803 VP.n55 VP.n13 161.3
R804 VP.n23 VP.t6 90.2299
R805 VP.n54 VP.n53 89.0887
R806 VP.n96 VP.n0 89.0887
R807 VP.n52 VP.n14 89.0887
R808 VP.n24 VP.n23 58.4531
R809 VP.n54 VP.t4 57.9031
R810 VP.n68 VP.t2 57.9031
R811 VP.n81 VP.t3 57.9031
R812 VP.n0 VP.t7 57.9031
R813 VP.n14 VP.t0 57.9031
R814 VP.n37 VP.t1 57.9031
R815 VP.n24 VP.t5 57.9031
R816 VP.n75 VP.n74 56.5193
R817 VP.n31 VP.n30 56.5193
R818 VP.n53 VP.n52 54.6963
R819 VP.n62 VP.n61 47.2923
R820 VP.n88 VP.n87 47.2923
R821 VP.n44 VP.n43 47.2923
R822 VP.n61 VP.n60 33.6945
R823 VP.n88 VP.n2 33.6945
R824 VP.n44 VP.n16 33.6945
R825 VP.n56 VP.n55 24.4675
R826 VP.n56 VP.n12 24.4675
R827 VP.n60 VP.n12 24.4675
R828 VP.n62 VP.n10 24.4675
R829 VP.n66 VP.n10 24.4675
R830 VP.n67 VP.n66 24.4675
R831 VP.n69 VP.n8 24.4675
R832 VP.n73 VP.n8 24.4675
R833 VP.n74 VP.n73 24.4675
R834 VP.n75 VP.n6 24.4675
R835 VP.n79 VP.n6 24.4675
R836 VP.n80 VP.n79 24.4675
R837 VP.n82 VP.n4 24.4675
R838 VP.n86 VP.n4 24.4675
R839 VP.n87 VP.n86 24.4675
R840 VP.n92 VP.n2 24.4675
R841 VP.n93 VP.n92 24.4675
R842 VP.n94 VP.n93 24.4675
R843 VP.n48 VP.n16 24.4675
R844 VP.n49 VP.n48 24.4675
R845 VP.n50 VP.n49 24.4675
R846 VP.n31 VP.n20 24.4675
R847 VP.n35 VP.n20 24.4675
R848 VP.n36 VP.n35 24.4675
R849 VP.n38 VP.n18 24.4675
R850 VP.n42 VP.n18 24.4675
R851 VP.n43 VP.n42 24.4675
R852 VP.n25 VP.n22 24.4675
R853 VP.n29 VP.n22 24.4675
R854 VP.n30 VP.n29 24.4675
R855 VP.n69 VP.n68 16.6381
R856 VP.n81 VP.n80 16.6381
R857 VP.n37 VP.n36 16.6381
R858 VP.n25 VP.n24 16.6381
R859 VP.n68 VP.n67 7.82994
R860 VP.n82 VP.n81 7.82994
R861 VP.n38 VP.n37 7.82994
R862 VP.n26 VP.n23 2.50736
R863 VP.n55 VP.n54 0.97918
R864 VP.n94 VP.n0 0.97918
R865 VP.n50 VP.n14 0.97918
R866 VP.n52 VP.n51 0.354971
R867 VP.n53 VP.n13 0.354971
R868 VP.n96 VP.n95 0.354971
R869 VP VP.n96 0.26696
R870 VP.n27 VP.n26 0.189894
R871 VP.n28 VP.n27 0.189894
R872 VP.n28 VP.n21 0.189894
R873 VP.n32 VP.n21 0.189894
R874 VP.n33 VP.n32 0.189894
R875 VP.n34 VP.n33 0.189894
R876 VP.n34 VP.n19 0.189894
R877 VP.n39 VP.n19 0.189894
R878 VP.n40 VP.n39 0.189894
R879 VP.n41 VP.n40 0.189894
R880 VP.n41 VP.n17 0.189894
R881 VP.n45 VP.n17 0.189894
R882 VP.n46 VP.n45 0.189894
R883 VP.n47 VP.n46 0.189894
R884 VP.n47 VP.n15 0.189894
R885 VP.n51 VP.n15 0.189894
R886 VP.n57 VP.n13 0.189894
R887 VP.n58 VP.n57 0.189894
R888 VP.n59 VP.n58 0.189894
R889 VP.n59 VP.n11 0.189894
R890 VP.n63 VP.n11 0.189894
R891 VP.n64 VP.n63 0.189894
R892 VP.n65 VP.n64 0.189894
R893 VP.n65 VP.n9 0.189894
R894 VP.n70 VP.n9 0.189894
R895 VP.n71 VP.n70 0.189894
R896 VP.n72 VP.n71 0.189894
R897 VP.n72 VP.n7 0.189894
R898 VP.n76 VP.n7 0.189894
R899 VP.n77 VP.n76 0.189894
R900 VP.n78 VP.n77 0.189894
R901 VP.n78 VP.n5 0.189894
R902 VP.n83 VP.n5 0.189894
R903 VP.n84 VP.n83 0.189894
R904 VP.n85 VP.n84 0.189894
R905 VP.n85 VP.n3 0.189894
R906 VP.n89 VP.n3 0.189894
R907 VP.n90 VP.n89 0.189894
R908 VP.n91 VP.n90 0.189894
R909 VP.n91 VP.n1 0.189894
R910 VP.n95 VP.n1 0.189894
R911 VDD1 VDD1.n0 80.6347
R912 VDD1.n3 VDD1.n2 80.521
R913 VDD1.n3 VDD1.n1 80.521
R914 VDD1.n5 VDD1.n4 78.7746
R915 VDD1.n5 VDD1.n3 48.488
R916 VDD1.n4 VDD1.t6 3.51455
R917 VDD1.n4 VDD1.t7 3.51455
R918 VDD1.n0 VDD1.t1 3.51455
R919 VDD1.n0 VDD1.t2 3.51455
R920 VDD1.n2 VDD1.t4 3.51455
R921 VDD1.n2 VDD1.t0 3.51455
R922 VDD1.n1 VDD1.t3 3.51455
R923 VDD1.n1 VDD1.t5 3.51455
R924 VDD1 VDD1.n5 1.74403
R925 B.n445 B.n444 585
R926 B.n443 B.n150 585
R927 B.n442 B.n441 585
R928 B.n440 B.n151 585
R929 B.n439 B.n438 585
R930 B.n437 B.n152 585
R931 B.n436 B.n435 585
R932 B.n434 B.n153 585
R933 B.n433 B.n432 585
R934 B.n431 B.n154 585
R935 B.n430 B.n429 585
R936 B.n428 B.n155 585
R937 B.n427 B.n426 585
R938 B.n425 B.n156 585
R939 B.n424 B.n423 585
R940 B.n422 B.n157 585
R941 B.n421 B.n420 585
R942 B.n419 B.n158 585
R943 B.n418 B.n417 585
R944 B.n416 B.n159 585
R945 B.n415 B.n414 585
R946 B.n413 B.n160 585
R947 B.n412 B.n411 585
R948 B.n410 B.n161 585
R949 B.n409 B.n408 585
R950 B.n407 B.n162 585
R951 B.n406 B.n405 585
R952 B.n404 B.n163 585
R953 B.n403 B.n402 585
R954 B.n401 B.n164 585
R955 B.n400 B.n399 585
R956 B.n398 B.n165 585
R957 B.n397 B.n396 585
R958 B.n395 B.n166 585
R959 B.n394 B.n393 585
R960 B.n389 B.n167 585
R961 B.n388 B.n387 585
R962 B.n386 B.n168 585
R963 B.n385 B.n384 585
R964 B.n383 B.n169 585
R965 B.n382 B.n381 585
R966 B.n380 B.n170 585
R967 B.n379 B.n378 585
R968 B.n376 B.n171 585
R969 B.n375 B.n374 585
R970 B.n373 B.n174 585
R971 B.n372 B.n371 585
R972 B.n370 B.n175 585
R973 B.n369 B.n368 585
R974 B.n367 B.n176 585
R975 B.n366 B.n365 585
R976 B.n364 B.n177 585
R977 B.n363 B.n362 585
R978 B.n361 B.n178 585
R979 B.n360 B.n359 585
R980 B.n358 B.n179 585
R981 B.n357 B.n356 585
R982 B.n355 B.n180 585
R983 B.n354 B.n353 585
R984 B.n352 B.n181 585
R985 B.n351 B.n350 585
R986 B.n349 B.n182 585
R987 B.n348 B.n347 585
R988 B.n346 B.n183 585
R989 B.n345 B.n344 585
R990 B.n343 B.n184 585
R991 B.n342 B.n341 585
R992 B.n340 B.n185 585
R993 B.n339 B.n338 585
R994 B.n337 B.n186 585
R995 B.n336 B.n335 585
R996 B.n334 B.n187 585
R997 B.n333 B.n332 585
R998 B.n331 B.n188 585
R999 B.n330 B.n329 585
R1000 B.n328 B.n189 585
R1001 B.n327 B.n326 585
R1002 B.n446 B.n149 585
R1003 B.n448 B.n447 585
R1004 B.n449 B.n148 585
R1005 B.n451 B.n450 585
R1006 B.n452 B.n147 585
R1007 B.n454 B.n453 585
R1008 B.n455 B.n146 585
R1009 B.n457 B.n456 585
R1010 B.n458 B.n145 585
R1011 B.n460 B.n459 585
R1012 B.n461 B.n144 585
R1013 B.n463 B.n462 585
R1014 B.n464 B.n143 585
R1015 B.n466 B.n465 585
R1016 B.n467 B.n142 585
R1017 B.n469 B.n468 585
R1018 B.n470 B.n141 585
R1019 B.n472 B.n471 585
R1020 B.n473 B.n140 585
R1021 B.n475 B.n474 585
R1022 B.n476 B.n139 585
R1023 B.n478 B.n477 585
R1024 B.n479 B.n138 585
R1025 B.n481 B.n480 585
R1026 B.n482 B.n137 585
R1027 B.n484 B.n483 585
R1028 B.n485 B.n136 585
R1029 B.n487 B.n486 585
R1030 B.n488 B.n135 585
R1031 B.n490 B.n489 585
R1032 B.n491 B.n134 585
R1033 B.n493 B.n492 585
R1034 B.n494 B.n133 585
R1035 B.n496 B.n495 585
R1036 B.n497 B.n132 585
R1037 B.n499 B.n498 585
R1038 B.n500 B.n131 585
R1039 B.n502 B.n501 585
R1040 B.n503 B.n130 585
R1041 B.n505 B.n504 585
R1042 B.n506 B.n129 585
R1043 B.n508 B.n507 585
R1044 B.n509 B.n128 585
R1045 B.n511 B.n510 585
R1046 B.n512 B.n127 585
R1047 B.n514 B.n513 585
R1048 B.n515 B.n126 585
R1049 B.n517 B.n516 585
R1050 B.n518 B.n125 585
R1051 B.n520 B.n519 585
R1052 B.n521 B.n124 585
R1053 B.n523 B.n522 585
R1054 B.n524 B.n123 585
R1055 B.n526 B.n525 585
R1056 B.n527 B.n122 585
R1057 B.n529 B.n528 585
R1058 B.n530 B.n121 585
R1059 B.n532 B.n531 585
R1060 B.n533 B.n120 585
R1061 B.n535 B.n534 585
R1062 B.n536 B.n119 585
R1063 B.n538 B.n537 585
R1064 B.n539 B.n118 585
R1065 B.n541 B.n540 585
R1066 B.n542 B.n117 585
R1067 B.n544 B.n543 585
R1068 B.n545 B.n116 585
R1069 B.n547 B.n546 585
R1070 B.n548 B.n115 585
R1071 B.n550 B.n549 585
R1072 B.n551 B.n114 585
R1073 B.n553 B.n552 585
R1074 B.n554 B.n113 585
R1075 B.n556 B.n555 585
R1076 B.n557 B.n112 585
R1077 B.n559 B.n558 585
R1078 B.n560 B.n111 585
R1079 B.n562 B.n561 585
R1080 B.n563 B.n110 585
R1081 B.n565 B.n564 585
R1082 B.n566 B.n109 585
R1083 B.n568 B.n567 585
R1084 B.n569 B.n108 585
R1085 B.n571 B.n570 585
R1086 B.n572 B.n107 585
R1087 B.n574 B.n573 585
R1088 B.n575 B.n106 585
R1089 B.n577 B.n576 585
R1090 B.n578 B.n105 585
R1091 B.n580 B.n579 585
R1092 B.n581 B.n104 585
R1093 B.n583 B.n582 585
R1094 B.n584 B.n103 585
R1095 B.n586 B.n585 585
R1096 B.n587 B.n102 585
R1097 B.n589 B.n588 585
R1098 B.n590 B.n101 585
R1099 B.n592 B.n591 585
R1100 B.n593 B.n100 585
R1101 B.n595 B.n594 585
R1102 B.n596 B.n99 585
R1103 B.n598 B.n597 585
R1104 B.n599 B.n98 585
R1105 B.n601 B.n600 585
R1106 B.n602 B.n97 585
R1107 B.n604 B.n603 585
R1108 B.n605 B.n96 585
R1109 B.n607 B.n606 585
R1110 B.n608 B.n95 585
R1111 B.n610 B.n609 585
R1112 B.n611 B.n94 585
R1113 B.n613 B.n612 585
R1114 B.n614 B.n93 585
R1115 B.n616 B.n615 585
R1116 B.n617 B.n92 585
R1117 B.n619 B.n618 585
R1118 B.n620 B.n91 585
R1119 B.n622 B.n621 585
R1120 B.n623 B.n90 585
R1121 B.n625 B.n624 585
R1122 B.n626 B.n89 585
R1123 B.n628 B.n627 585
R1124 B.n629 B.n88 585
R1125 B.n631 B.n630 585
R1126 B.n632 B.n87 585
R1127 B.n634 B.n633 585
R1128 B.n635 B.n86 585
R1129 B.n637 B.n636 585
R1130 B.n638 B.n85 585
R1131 B.n640 B.n639 585
R1132 B.n641 B.n84 585
R1133 B.n643 B.n642 585
R1134 B.n644 B.n83 585
R1135 B.n646 B.n645 585
R1136 B.n647 B.n82 585
R1137 B.n649 B.n648 585
R1138 B.n650 B.n81 585
R1139 B.n652 B.n651 585
R1140 B.n653 B.n80 585
R1141 B.n655 B.n654 585
R1142 B.n772 B.n771 585
R1143 B.n770 B.n37 585
R1144 B.n769 B.n768 585
R1145 B.n767 B.n38 585
R1146 B.n766 B.n765 585
R1147 B.n764 B.n39 585
R1148 B.n763 B.n762 585
R1149 B.n761 B.n40 585
R1150 B.n760 B.n759 585
R1151 B.n758 B.n41 585
R1152 B.n757 B.n756 585
R1153 B.n755 B.n42 585
R1154 B.n754 B.n753 585
R1155 B.n752 B.n43 585
R1156 B.n751 B.n750 585
R1157 B.n749 B.n44 585
R1158 B.n748 B.n747 585
R1159 B.n746 B.n45 585
R1160 B.n745 B.n744 585
R1161 B.n743 B.n46 585
R1162 B.n742 B.n741 585
R1163 B.n740 B.n47 585
R1164 B.n739 B.n738 585
R1165 B.n737 B.n48 585
R1166 B.n736 B.n735 585
R1167 B.n734 B.n49 585
R1168 B.n733 B.n732 585
R1169 B.n731 B.n50 585
R1170 B.n730 B.n729 585
R1171 B.n728 B.n51 585
R1172 B.n727 B.n726 585
R1173 B.n725 B.n52 585
R1174 B.n724 B.n723 585
R1175 B.n722 B.n53 585
R1176 B.n720 B.n719 585
R1177 B.n718 B.n56 585
R1178 B.n717 B.n716 585
R1179 B.n715 B.n57 585
R1180 B.n714 B.n713 585
R1181 B.n712 B.n58 585
R1182 B.n711 B.n710 585
R1183 B.n709 B.n59 585
R1184 B.n708 B.n707 585
R1185 B.n706 B.n705 585
R1186 B.n704 B.n63 585
R1187 B.n703 B.n702 585
R1188 B.n701 B.n64 585
R1189 B.n700 B.n699 585
R1190 B.n698 B.n65 585
R1191 B.n697 B.n696 585
R1192 B.n695 B.n66 585
R1193 B.n694 B.n693 585
R1194 B.n692 B.n67 585
R1195 B.n691 B.n690 585
R1196 B.n689 B.n68 585
R1197 B.n688 B.n687 585
R1198 B.n686 B.n69 585
R1199 B.n685 B.n684 585
R1200 B.n683 B.n70 585
R1201 B.n682 B.n681 585
R1202 B.n680 B.n71 585
R1203 B.n679 B.n678 585
R1204 B.n677 B.n72 585
R1205 B.n676 B.n675 585
R1206 B.n674 B.n73 585
R1207 B.n673 B.n672 585
R1208 B.n671 B.n74 585
R1209 B.n670 B.n669 585
R1210 B.n668 B.n75 585
R1211 B.n667 B.n666 585
R1212 B.n665 B.n76 585
R1213 B.n664 B.n663 585
R1214 B.n662 B.n77 585
R1215 B.n661 B.n660 585
R1216 B.n659 B.n78 585
R1217 B.n658 B.n657 585
R1218 B.n656 B.n79 585
R1219 B.n773 B.n36 585
R1220 B.n775 B.n774 585
R1221 B.n776 B.n35 585
R1222 B.n778 B.n777 585
R1223 B.n779 B.n34 585
R1224 B.n781 B.n780 585
R1225 B.n782 B.n33 585
R1226 B.n784 B.n783 585
R1227 B.n785 B.n32 585
R1228 B.n787 B.n786 585
R1229 B.n788 B.n31 585
R1230 B.n790 B.n789 585
R1231 B.n791 B.n30 585
R1232 B.n793 B.n792 585
R1233 B.n794 B.n29 585
R1234 B.n796 B.n795 585
R1235 B.n797 B.n28 585
R1236 B.n799 B.n798 585
R1237 B.n800 B.n27 585
R1238 B.n802 B.n801 585
R1239 B.n803 B.n26 585
R1240 B.n805 B.n804 585
R1241 B.n806 B.n25 585
R1242 B.n808 B.n807 585
R1243 B.n809 B.n24 585
R1244 B.n811 B.n810 585
R1245 B.n812 B.n23 585
R1246 B.n814 B.n813 585
R1247 B.n815 B.n22 585
R1248 B.n817 B.n816 585
R1249 B.n818 B.n21 585
R1250 B.n820 B.n819 585
R1251 B.n821 B.n20 585
R1252 B.n823 B.n822 585
R1253 B.n824 B.n19 585
R1254 B.n826 B.n825 585
R1255 B.n827 B.n18 585
R1256 B.n829 B.n828 585
R1257 B.n830 B.n17 585
R1258 B.n832 B.n831 585
R1259 B.n833 B.n16 585
R1260 B.n835 B.n834 585
R1261 B.n836 B.n15 585
R1262 B.n838 B.n837 585
R1263 B.n839 B.n14 585
R1264 B.n841 B.n840 585
R1265 B.n842 B.n13 585
R1266 B.n844 B.n843 585
R1267 B.n845 B.n12 585
R1268 B.n847 B.n846 585
R1269 B.n848 B.n11 585
R1270 B.n850 B.n849 585
R1271 B.n851 B.n10 585
R1272 B.n853 B.n852 585
R1273 B.n854 B.n9 585
R1274 B.n856 B.n855 585
R1275 B.n857 B.n8 585
R1276 B.n859 B.n858 585
R1277 B.n860 B.n7 585
R1278 B.n862 B.n861 585
R1279 B.n863 B.n6 585
R1280 B.n865 B.n864 585
R1281 B.n866 B.n5 585
R1282 B.n868 B.n867 585
R1283 B.n869 B.n4 585
R1284 B.n871 B.n870 585
R1285 B.n872 B.n3 585
R1286 B.n874 B.n873 585
R1287 B.n875 B.n0 585
R1288 B.n2 B.n1 585
R1289 B.n225 B.n224 585
R1290 B.n226 B.n223 585
R1291 B.n228 B.n227 585
R1292 B.n229 B.n222 585
R1293 B.n231 B.n230 585
R1294 B.n232 B.n221 585
R1295 B.n234 B.n233 585
R1296 B.n235 B.n220 585
R1297 B.n237 B.n236 585
R1298 B.n238 B.n219 585
R1299 B.n240 B.n239 585
R1300 B.n241 B.n218 585
R1301 B.n243 B.n242 585
R1302 B.n244 B.n217 585
R1303 B.n246 B.n245 585
R1304 B.n247 B.n216 585
R1305 B.n249 B.n248 585
R1306 B.n250 B.n215 585
R1307 B.n252 B.n251 585
R1308 B.n253 B.n214 585
R1309 B.n255 B.n254 585
R1310 B.n256 B.n213 585
R1311 B.n258 B.n257 585
R1312 B.n259 B.n212 585
R1313 B.n261 B.n260 585
R1314 B.n262 B.n211 585
R1315 B.n264 B.n263 585
R1316 B.n265 B.n210 585
R1317 B.n267 B.n266 585
R1318 B.n268 B.n209 585
R1319 B.n270 B.n269 585
R1320 B.n271 B.n208 585
R1321 B.n273 B.n272 585
R1322 B.n274 B.n207 585
R1323 B.n276 B.n275 585
R1324 B.n277 B.n206 585
R1325 B.n279 B.n278 585
R1326 B.n280 B.n205 585
R1327 B.n282 B.n281 585
R1328 B.n283 B.n204 585
R1329 B.n285 B.n284 585
R1330 B.n286 B.n203 585
R1331 B.n288 B.n287 585
R1332 B.n289 B.n202 585
R1333 B.n291 B.n290 585
R1334 B.n292 B.n201 585
R1335 B.n294 B.n293 585
R1336 B.n295 B.n200 585
R1337 B.n297 B.n296 585
R1338 B.n298 B.n199 585
R1339 B.n300 B.n299 585
R1340 B.n301 B.n198 585
R1341 B.n303 B.n302 585
R1342 B.n304 B.n197 585
R1343 B.n306 B.n305 585
R1344 B.n307 B.n196 585
R1345 B.n309 B.n308 585
R1346 B.n310 B.n195 585
R1347 B.n312 B.n311 585
R1348 B.n313 B.n194 585
R1349 B.n315 B.n314 585
R1350 B.n316 B.n193 585
R1351 B.n318 B.n317 585
R1352 B.n319 B.n192 585
R1353 B.n321 B.n320 585
R1354 B.n322 B.n191 585
R1355 B.n324 B.n323 585
R1356 B.n325 B.n190 585
R1357 B.n326 B.n325 482.89
R1358 B.n444 B.n149 482.89
R1359 B.n654 B.n79 482.89
R1360 B.n773 B.n772 482.89
R1361 B.n390 B.t4 407.051
R1362 B.n60 B.t8 407.051
R1363 B.n172 B.t10 407.051
R1364 B.n54 B.t2 407.051
R1365 B.n391 B.t5 325.985
R1366 B.n61 B.t7 325.985
R1367 B.n173 B.t11 325.985
R1368 B.n55 B.t1 325.985
R1369 B.n172 B.t9 267.284
R1370 B.n390 B.t3 267.284
R1371 B.n60 B.t6 267.284
R1372 B.n54 B.t0 267.284
R1373 B.n877 B.n876 256.663
R1374 B.n876 B.n875 235.042
R1375 B.n876 B.n2 235.042
R1376 B.n326 B.n189 163.367
R1377 B.n330 B.n189 163.367
R1378 B.n331 B.n330 163.367
R1379 B.n332 B.n331 163.367
R1380 B.n332 B.n187 163.367
R1381 B.n336 B.n187 163.367
R1382 B.n337 B.n336 163.367
R1383 B.n338 B.n337 163.367
R1384 B.n338 B.n185 163.367
R1385 B.n342 B.n185 163.367
R1386 B.n343 B.n342 163.367
R1387 B.n344 B.n343 163.367
R1388 B.n344 B.n183 163.367
R1389 B.n348 B.n183 163.367
R1390 B.n349 B.n348 163.367
R1391 B.n350 B.n349 163.367
R1392 B.n350 B.n181 163.367
R1393 B.n354 B.n181 163.367
R1394 B.n355 B.n354 163.367
R1395 B.n356 B.n355 163.367
R1396 B.n356 B.n179 163.367
R1397 B.n360 B.n179 163.367
R1398 B.n361 B.n360 163.367
R1399 B.n362 B.n361 163.367
R1400 B.n362 B.n177 163.367
R1401 B.n366 B.n177 163.367
R1402 B.n367 B.n366 163.367
R1403 B.n368 B.n367 163.367
R1404 B.n368 B.n175 163.367
R1405 B.n372 B.n175 163.367
R1406 B.n373 B.n372 163.367
R1407 B.n374 B.n373 163.367
R1408 B.n374 B.n171 163.367
R1409 B.n379 B.n171 163.367
R1410 B.n380 B.n379 163.367
R1411 B.n381 B.n380 163.367
R1412 B.n381 B.n169 163.367
R1413 B.n385 B.n169 163.367
R1414 B.n386 B.n385 163.367
R1415 B.n387 B.n386 163.367
R1416 B.n387 B.n167 163.367
R1417 B.n394 B.n167 163.367
R1418 B.n395 B.n394 163.367
R1419 B.n396 B.n395 163.367
R1420 B.n396 B.n165 163.367
R1421 B.n400 B.n165 163.367
R1422 B.n401 B.n400 163.367
R1423 B.n402 B.n401 163.367
R1424 B.n402 B.n163 163.367
R1425 B.n406 B.n163 163.367
R1426 B.n407 B.n406 163.367
R1427 B.n408 B.n407 163.367
R1428 B.n408 B.n161 163.367
R1429 B.n412 B.n161 163.367
R1430 B.n413 B.n412 163.367
R1431 B.n414 B.n413 163.367
R1432 B.n414 B.n159 163.367
R1433 B.n418 B.n159 163.367
R1434 B.n419 B.n418 163.367
R1435 B.n420 B.n419 163.367
R1436 B.n420 B.n157 163.367
R1437 B.n424 B.n157 163.367
R1438 B.n425 B.n424 163.367
R1439 B.n426 B.n425 163.367
R1440 B.n426 B.n155 163.367
R1441 B.n430 B.n155 163.367
R1442 B.n431 B.n430 163.367
R1443 B.n432 B.n431 163.367
R1444 B.n432 B.n153 163.367
R1445 B.n436 B.n153 163.367
R1446 B.n437 B.n436 163.367
R1447 B.n438 B.n437 163.367
R1448 B.n438 B.n151 163.367
R1449 B.n442 B.n151 163.367
R1450 B.n443 B.n442 163.367
R1451 B.n444 B.n443 163.367
R1452 B.n654 B.n653 163.367
R1453 B.n653 B.n652 163.367
R1454 B.n652 B.n81 163.367
R1455 B.n648 B.n81 163.367
R1456 B.n648 B.n647 163.367
R1457 B.n647 B.n646 163.367
R1458 B.n646 B.n83 163.367
R1459 B.n642 B.n83 163.367
R1460 B.n642 B.n641 163.367
R1461 B.n641 B.n640 163.367
R1462 B.n640 B.n85 163.367
R1463 B.n636 B.n85 163.367
R1464 B.n636 B.n635 163.367
R1465 B.n635 B.n634 163.367
R1466 B.n634 B.n87 163.367
R1467 B.n630 B.n87 163.367
R1468 B.n630 B.n629 163.367
R1469 B.n629 B.n628 163.367
R1470 B.n628 B.n89 163.367
R1471 B.n624 B.n89 163.367
R1472 B.n624 B.n623 163.367
R1473 B.n623 B.n622 163.367
R1474 B.n622 B.n91 163.367
R1475 B.n618 B.n91 163.367
R1476 B.n618 B.n617 163.367
R1477 B.n617 B.n616 163.367
R1478 B.n616 B.n93 163.367
R1479 B.n612 B.n93 163.367
R1480 B.n612 B.n611 163.367
R1481 B.n611 B.n610 163.367
R1482 B.n610 B.n95 163.367
R1483 B.n606 B.n95 163.367
R1484 B.n606 B.n605 163.367
R1485 B.n605 B.n604 163.367
R1486 B.n604 B.n97 163.367
R1487 B.n600 B.n97 163.367
R1488 B.n600 B.n599 163.367
R1489 B.n599 B.n598 163.367
R1490 B.n598 B.n99 163.367
R1491 B.n594 B.n99 163.367
R1492 B.n594 B.n593 163.367
R1493 B.n593 B.n592 163.367
R1494 B.n592 B.n101 163.367
R1495 B.n588 B.n101 163.367
R1496 B.n588 B.n587 163.367
R1497 B.n587 B.n586 163.367
R1498 B.n586 B.n103 163.367
R1499 B.n582 B.n103 163.367
R1500 B.n582 B.n581 163.367
R1501 B.n581 B.n580 163.367
R1502 B.n580 B.n105 163.367
R1503 B.n576 B.n105 163.367
R1504 B.n576 B.n575 163.367
R1505 B.n575 B.n574 163.367
R1506 B.n574 B.n107 163.367
R1507 B.n570 B.n107 163.367
R1508 B.n570 B.n569 163.367
R1509 B.n569 B.n568 163.367
R1510 B.n568 B.n109 163.367
R1511 B.n564 B.n109 163.367
R1512 B.n564 B.n563 163.367
R1513 B.n563 B.n562 163.367
R1514 B.n562 B.n111 163.367
R1515 B.n558 B.n111 163.367
R1516 B.n558 B.n557 163.367
R1517 B.n557 B.n556 163.367
R1518 B.n556 B.n113 163.367
R1519 B.n552 B.n113 163.367
R1520 B.n552 B.n551 163.367
R1521 B.n551 B.n550 163.367
R1522 B.n550 B.n115 163.367
R1523 B.n546 B.n115 163.367
R1524 B.n546 B.n545 163.367
R1525 B.n545 B.n544 163.367
R1526 B.n544 B.n117 163.367
R1527 B.n540 B.n117 163.367
R1528 B.n540 B.n539 163.367
R1529 B.n539 B.n538 163.367
R1530 B.n538 B.n119 163.367
R1531 B.n534 B.n119 163.367
R1532 B.n534 B.n533 163.367
R1533 B.n533 B.n532 163.367
R1534 B.n532 B.n121 163.367
R1535 B.n528 B.n121 163.367
R1536 B.n528 B.n527 163.367
R1537 B.n527 B.n526 163.367
R1538 B.n526 B.n123 163.367
R1539 B.n522 B.n123 163.367
R1540 B.n522 B.n521 163.367
R1541 B.n521 B.n520 163.367
R1542 B.n520 B.n125 163.367
R1543 B.n516 B.n125 163.367
R1544 B.n516 B.n515 163.367
R1545 B.n515 B.n514 163.367
R1546 B.n514 B.n127 163.367
R1547 B.n510 B.n127 163.367
R1548 B.n510 B.n509 163.367
R1549 B.n509 B.n508 163.367
R1550 B.n508 B.n129 163.367
R1551 B.n504 B.n129 163.367
R1552 B.n504 B.n503 163.367
R1553 B.n503 B.n502 163.367
R1554 B.n502 B.n131 163.367
R1555 B.n498 B.n131 163.367
R1556 B.n498 B.n497 163.367
R1557 B.n497 B.n496 163.367
R1558 B.n496 B.n133 163.367
R1559 B.n492 B.n133 163.367
R1560 B.n492 B.n491 163.367
R1561 B.n491 B.n490 163.367
R1562 B.n490 B.n135 163.367
R1563 B.n486 B.n135 163.367
R1564 B.n486 B.n485 163.367
R1565 B.n485 B.n484 163.367
R1566 B.n484 B.n137 163.367
R1567 B.n480 B.n137 163.367
R1568 B.n480 B.n479 163.367
R1569 B.n479 B.n478 163.367
R1570 B.n478 B.n139 163.367
R1571 B.n474 B.n139 163.367
R1572 B.n474 B.n473 163.367
R1573 B.n473 B.n472 163.367
R1574 B.n472 B.n141 163.367
R1575 B.n468 B.n141 163.367
R1576 B.n468 B.n467 163.367
R1577 B.n467 B.n466 163.367
R1578 B.n466 B.n143 163.367
R1579 B.n462 B.n143 163.367
R1580 B.n462 B.n461 163.367
R1581 B.n461 B.n460 163.367
R1582 B.n460 B.n145 163.367
R1583 B.n456 B.n145 163.367
R1584 B.n456 B.n455 163.367
R1585 B.n455 B.n454 163.367
R1586 B.n454 B.n147 163.367
R1587 B.n450 B.n147 163.367
R1588 B.n450 B.n449 163.367
R1589 B.n449 B.n448 163.367
R1590 B.n448 B.n149 163.367
R1591 B.n772 B.n37 163.367
R1592 B.n768 B.n37 163.367
R1593 B.n768 B.n767 163.367
R1594 B.n767 B.n766 163.367
R1595 B.n766 B.n39 163.367
R1596 B.n762 B.n39 163.367
R1597 B.n762 B.n761 163.367
R1598 B.n761 B.n760 163.367
R1599 B.n760 B.n41 163.367
R1600 B.n756 B.n41 163.367
R1601 B.n756 B.n755 163.367
R1602 B.n755 B.n754 163.367
R1603 B.n754 B.n43 163.367
R1604 B.n750 B.n43 163.367
R1605 B.n750 B.n749 163.367
R1606 B.n749 B.n748 163.367
R1607 B.n748 B.n45 163.367
R1608 B.n744 B.n45 163.367
R1609 B.n744 B.n743 163.367
R1610 B.n743 B.n742 163.367
R1611 B.n742 B.n47 163.367
R1612 B.n738 B.n47 163.367
R1613 B.n738 B.n737 163.367
R1614 B.n737 B.n736 163.367
R1615 B.n736 B.n49 163.367
R1616 B.n732 B.n49 163.367
R1617 B.n732 B.n731 163.367
R1618 B.n731 B.n730 163.367
R1619 B.n730 B.n51 163.367
R1620 B.n726 B.n51 163.367
R1621 B.n726 B.n725 163.367
R1622 B.n725 B.n724 163.367
R1623 B.n724 B.n53 163.367
R1624 B.n719 B.n53 163.367
R1625 B.n719 B.n718 163.367
R1626 B.n718 B.n717 163.367
R1627 B.n717 B.n57 163.367
R1628 B.n713 B.n57 163.367
R1629 B.n713 B.n712 163.367
R1630 B.n712 B.n711 163.367
R1631 B.n711 B.n59 163.367
R1632 B.n707 B.n59 163.367
R1633 B.n707 B.n706 163.367
R1634 B.n706 B.n63 163.367
R1635 B.n702 B.n63 163.367
R1636 B.n702 B.n701 163.367
R1637 B.n701 B.n700 163.367
R1638 B.n700 B.n65 163.367
R1639 B.n696 B.n65 163.367
R1640 B.n696 B.n695 163.367
R1641 B.n695 B.n694 163.367
R1642 B.n694 B.n67 163.367
R1643 B.n690 B.n67 163.367
R1644 B.n690 B.n689 163.367
R1645 B.n689 B.n688 163.367
R1646 B.n688 B.n69 163.367
R1647 B.n684 B.n69 163.367
R1648 B.n684 B.n683 163.367
R1649 B.n683 B.n682 163.367
R1650 B.n682 B.n71 163.367
R1651 B.n678 B.n71 163.367
R1652 B.n678 B.n677 163.367
R1653 B.n677 B.n676 163.367
R1654 B.n676 B.n73 163.367
R1655 B.n672 B.n73 163.367
R1656 B.n672 B.n671 163.367
R1657 B.n671 B.n670 163.367
R1658 B.n670 B.n75 163.367
R1659 B.n666 B.n75 163.367
R1660 B.n666 B.n665 163.367
R1661 B.n665 B.n664 163.367
R1662 B.n664 B.n77 163.367
R1663 B.n660 B.n77 163.367
R1664 B.n660 B.n659 163.367
R1665 B.n659 B.n658 163.367
R1666 B.n658 B.n79 163.367
R1667 B.n774 B.n773 163.367
R1668 B.n774 B.n35 163.367
R1669 B.n778 B.n35 163.367
R1670 B.n779 B.n778 163.367
R1671 B.n780 B.n779 163.367
R1672 B.n780 B.n33 163.367
R1673 B.n784 B.n33 163.367
R1674 B.n785 B.n784 163.367
R1675 B.n786 B.n785 163.367
R1676 B.n786 B.n31 163.367
R1677 B.n790 B.n31 163.367
R1678 B.n791 B.n790 163.367
R1679 B.n792 B.n791 163.367
R1680 B.n792 B.n29 163.367
R1681 B.n796 B.n29 163.367
R1682 B.n797 B.n796 163.367
R1683 B.n798 B.n797 163.367
R1684 B.n798 B.n27 163.367
R1685 B.n802 B.n27 163.367
R1686 B.n803 B.n802 163.367
R1687 B.n804 B.n803 163.367
R1688 B.n804 B.n25 163.367
R1689 B.n808 B.n25 163.367
R1690 B.n809 B.n808 163.367
R1691 B.n810 B.n809 163.367
R1692 B.n810 B.n23 163.367
R1693 B.n814 B.n23 163.367
R1694 B.n815 B.n814 163.367
R1695 B.n816 B.n815 163.367
R1696 B.n816 B.n21 163.367
R1697 B.n820 B.n21 163.367
R1698 B.n821 B.n820 163.367
R1699 B.n822 B.n821 163.367
R1700 B.n822 B.n19 163.367
R1701 B.n826 B.n19 163.367
R1702 B.n827 B.n826 163.367
R1703 B.n828 B.n827 163.367
R1704 B.n828 B.n17 163.367
R1705 B.n832 B.n17 163.367
R1706 B.n833 B.n832 163.367
R1707 B.n834 B.n833 163.367
R1708 B.n834 B.n15 163.367
R1709 B.n838 B.n15 163.367
R1710 B.n839 B.n838 163.367
R1711 B.n840 B.n839 163.367
R1712 B.n840 B.n13 163.367
R1713 B.n844 B.n13 163.367
R1714 B.n845 B.n844 163.367
R1715 B.n846 B.n845 163.367
R1716 B.n846 B.n11 163.367
R1717 B.n850 B.n11 163.367
R1718 B.n851 B.n850 163.367
R1719 B.n852 B.n851 163.367
R1720 B.n852 B.n9 163.367
R1721 B.n856 B.n9 163.367
R1722 B.n857 B.n856 163.367
R1723 B.n858 B.n857 163.367
R1724 B.n858 B.n7 163.367
R1725 B.n862 B.n7 163.367
R1726 B.n863 B.n862 163.367
R1727 B.n864 B.n863 163.367
R1728 B.n864 B.n5 163.367
R1729 B.n868 B.n5 163.367
R1730 B.n869 B.n868 163.367
R1731 B.n870 B.n869 163.367
R1732 B.n870 B.n3 163.367
R1733 B.n874 B.n3 163.367
R1734 B.n875 B.n874 163.367
R1735 B.n224 B.n2 163.367
R1736 B.n224 B.n223 163.367
R1737 B.n228 B.n223 163.367
R1738 B.n229 B.n228 163.367
R1739 B.n230 B.n229 163.367
R1740 B.n230 B.n221 163.367
R1741 B.n234 B.n221 163.367
R1742 B.n235 B.n234 163.367
R1743 B.n236 B.n235 163.367
R1744 B.n236 B.n219 163.367
R1745 B.n240 B.n219 163.367
R1746 B.n241 B.n240 163.367
R1747 B.n242 B.n241 163.367
R1748 B.n242 B.n217 163.367
R1749 B.n246 B.n217 163.367
R1750 B.n247 B.n246 163.367
R1751 B.n248 B.n247 163.367
R1752 B.n248 B.n215 163.367
R1753 B.n252 B.n215 163.367
R1754 B.n253 B.n252 163.367
R1755 B.n254 B.n253 163.367
R1756 B.n254 B.n213 163.367
R1757 B.n258 B.n213 163.367
R1758 B.n259 B.n258 163.367
R1759 B.n260 B.n259 163.367
R1760 B.n260 B.n211 163.367
R1761 B.n264 B.n211 163.367
R1762 B.n265 B.n264 163.367
R1763 B.n266 B.n265 163.367
R1764 B.n266 B.n209 163.367
R1765 B.n270 B.n209 163.367
R1766 B.n271 B.n270 163.367
R1767 B.n272 B.n271 163.367
R1768 B.n272 B.n207 163.367
R1769 B.n276 B.n207 163.367
R1770 B.n277 B.n276 163.367
R1771 B.n278 B.n277 163.367
R1772 B.n278 B.n205 163.367
R1773 B.n282 B.n205 163.367
R1774 B.n283 B.n282 163.367
R1775 B.n284 B.n283 163.367
R1776 B.n284 B.n203 163.367
R1777 B.n288 B.n203 163.367
R1778 B.n289 B.n288 163.367
R1779 B.n290 B.n289 163.367
R1780 B.n290 B.n201 163.367
R1781 B.n294 B.n201 163.367
R1782 B.n295 B.n294 163.367
R1783 B.n296 B.n295 163.367
R1784 B.n296 B.n199 163.367
R1785 B.n300 B.n199 163.367
R1786 B.n301 B.n300 163.367
R1787 B.n302 B.n301 163.367
R1788 B.n302 B.n197 163.367
R1789 B.n306 B.n197 163.367
R1790 B.n307 B.n306 163.367
R1791 B.n308 B.n307 163.367
R1792 B.n308 B.n195 163.367
R1793 B.n312 B.n195 163.367
R1794 B.n313 B.n312 163.367
R1795 B.n314 B.n313 163.367
R1796 B.n314 B.n193 163.367
R1797 B.n318 B.n193 163.367
R1798 B.n319 B.n318 163.367
R1799 B.n320 B.n319 163.367
R1800 B.n320 B.n191 163.367
R1801 B.n324 B.n191 163.367
R1802 B.n325 B.n324 163.367
R1803 B.n173 B.n172 81.0672
R1804 B.n391 B.n390 81.0672
R1805 B.n61 B.n60 81.0672
R1806 B.n55 B.n54 81.0672
R1807 B.n377 B.n173 59.5399
R1808 B.n392 B.n391 59.5399
R1809 B.n62 B.n61 59.5399
R1810 B.n721 B.n55 59.5399
R1811 B.n771 B.n36 31.3761
R1812 B.n656 B.n655 31.3761
R1813 B.n446 B.n445 31.3761
R1814 B.n327 B.n190 31.3761
R1815 B B.n877 18.0485
R1816 B.n775 B.n36 10.6151
R1817 B.n776 B.n775 10.6151
R1818 B.n777 B.n776 10.6151
R1819 B.n777 B.n34 10.6151
R1820 B.n781 B.n34 10.6151
R1821 B.n782 B.n781 10.6151
R1822 B.n783 B.n782 10.6151
R1823 B.n783 B.n32 10.6151
R1824 B.n787 B.n32 10.6151
R1825 B.n788 B.n787 10.6151
R1826 B.n789 B.n788 10.6151
R1827 B.n789 B.n30 10.6151
R1828 B.n793 B.n30 10.6151
R1829 B.n794 B.n793 10.6151
R1830 B.n795 B.n794 10.6151
R1831 B.n795 B.n28 10.6151
R1832 B.n799 B.n28 10.6151
R1833 B.n800 B.n799 10.6151
R1834 B.n801 B.n800 10.6151
R1835 B.n801 B.n26 10.6151
R1836 B.n805 B.n26 10.6151
R1837 B.n806 B.n805 10.6151
R1838 B.n807 B.n806 10.6151
R1839 B.n807 B.n24 10.6151
R1840 B.n811 B.n24 10.6151
R1841 B.n812 B.n811 10.6151
R1842 B.n813 B.n812 10.6151
R1843 B.n813 B.n22 10.6151
R1844 B.n817 B.n22 10.6151
R1845 B.n818 B.n817 10.6151
R1846 B.n819 B.n818 10.6151
R1847 B.n819 B.n20 10.6151
R1848 B.n823 B.n20 10.6151
R1849 B.n824 B.n823 10.6151
R1850 B.n825 B.n824 10.6151
R1851 B.n825 B.n18 10.6151
R1852 B.n829 B.n18 10.6151
R1853 B.n830 B.n829 10.6151
R1854 B.n831 B.n830 10.6151
R1855 B.n831 B.n16 10.6151
R1856 B.n835 B.n16 10.6151
R1857 B.n836 B.n835 10.6151
R1858 B.n837 B.n836 10.6151
R1859 B.n837 B.n14 10.6151
R1860 B.n841 B.n14 10.6151
R1861 B.n842 B.n841 10.6151
R1862 B.n843 B.n842 10.6151
R1863 B.n843 B.n12 10.6151
R1864 B.n847 B.n12 10.6151
R1865 B.n848 B.n847 10.6151
R1866 B.n849 B.n848 10.6151
R1867 B.n849 B.n10 10.6151
R1868 B.n853 B.n10 10.6151
R1869 B.n854 B.n853 10.6151
R1870 B.n855 B.n854 10.6151
R1871 B.n855 B.n8 10.6151
R1872 B.n859 B.n8 10.6151
R1873 B.n860 B.n859 10.6151
R1874 B.n861 B.n860 10.6151
R1875 B.n861 B.n6 10.6151
R1876 B.n865 B.n6 10.6151
R1877 B.n866 B.n865 10.6151
R1878 B.n867 B.n866 10.6151
R1879 B.n867 B.n4 10.6151
R1880 B.n871 B.n4 10.6151
R1881 B.n872 B.n871 10.6151
R1882 B.n873 B.n872 10.6151
R1883 B.n873 B.n0 10.6151
R1884 B.n771 B.n770 10.6151
R1885 B.n770 B.n769 10.6151
R1886 B.n769 B.n38 10.6151
R1887 B.n765 B.n38 10.6151
R1888 B.n765 B.n764 10.6151
R1889 B.n764 B.n763 10.6151
R1890 B.n763 B.n40 10.6151
R1891 B.n759 B.n40 10.6151
R1892 B.n759 B.n758 10.6151
R1893 B.n758 B.n757 10.6151
R1894 B.n757 B.n42 10.6151
R1895 B.n753 B.n42 10.6151
R1896 B.n753 B.n752 10.6151
R1897 B.n752 B.n751 10.6151
R1898 B.n751 B.n44 10.6151
R1899 B.n747 B.n44 10.6151
R1900 B.n747 B.n746 10.6151
R1901 B.n746 B.n745 10.6151
R1902 B.n745 B.n46 10.6151
R1903 B.n741 B.n46 10.6151
R1904 B.n741 B.n740 10.6151
R1905 B.n740 B.n739 10.6151
R1906 B.n739 B.n48 10.6151
R1907 B.n735 B.n48 10.6151
R1908 B.n735 B.n734 10.6151
R1909 B.n734 B.n733 10.6151
R1910 B.n733 B.n50 10.6151
R1911 B.n729 B.n50 10.6151
R1912 B.n729 B.n728 10.6151
R1913 B.n728 B.n727 10.6151
R1914 B.n727 B.n52 10.6151
R1915 B.n723 B.n52 10.6151
R1916 B.n723 B.n722 10.6151
R1917 B.n720 B.n56 10.6151
R1918 B.n716 B.n56 10.6151
R1919 B.n716 B.n715 10.6151
R1920 B.n715 B.n714 10.6151
R1921 B.n714 B.n58 10.6151
R1922 B.n710 B.n58 10.6151
R1923 B.n710 B.n709 10.6151
R1924 B.n709 B.n708 10.6151
R1925 B.n705 B.n704 10.6151
R1926 B.n704 B.n703 10.6151
R1927 B.n703 B.n64 10.6151
R1928 B.n699 B.n64 10.6151
R1929 B.n699 B.n698 10.6151
R1930 B.n698 B.n697 10.6151
R1931 B.n697 B.n66 10.6151
R1932 B.n693 B.n66 10.6151
R1933 B.n693 B.n692 10.6151
R1934 B.n692 B.n691 10.6151
R1935 B.n691 B.n68 10.6151
R1936 B.n687 B.n68 10.6151
R1937 B.n687 B.n686 10.6151
R1938 B.n686 B.n685 10.6151
R1939 B.n685 B.n70 10.6151
R1940 B.n681 B.n70 10.6151
R1941 B.n681 B.n680 10.6151
R1942 B.n680 B.n679 10.6151
R1943 B.n679 B.n72 10.6151
R1944 B.n675 B.n72 10.6151
R1945 B.n675 B.n674 10.6151
R1946 B.n674 B.n673 10.6151
R1947 B.n673 B.n74 10.6151
R1948 B.n669 B.n74 10.6151
R1949 B.n669 B.n668 10.6151
R1950 B.n668 B.n667 10.6151
R1951 B.n667 B.n76 10.6151
R1952 B.n663 B.n76 10.6151
R1953 B.n663 B.n662 10.6151
R1954 B.n662 B.n661 10.6151
R1955 B.n661 B.n78 10.6151
R1956 B.n657 B.n78 10.6151
R1957 B.n657 B.n656 10.6151
R1958 B.n655 B.n80 10.6151
R1959 B.n651 B.n80 10.6151
R1960 B.n651 B.n650 10.6151
R1961 B.n650 B.n649 10.6151
R1962 B.n649 B.n82 10.6151
R1963 B.n645 B.n82 10.6151
R1964 B.n645 B.n644 10.6151
R1965 B.n644 B.n643 10.6151
R1966 B.n643 B.n84 10.6151
R1967 B.n639 B.n84 10.6151
R1968 B.n639 B.n638 10.6151
R1969 B.n638 B.n637 10.6151
R1970 B.n637 B.n86 10.6151
R1971 B.n633 B.n86 10.6151
R1972 B.n633 B.n632 10.6151
R1973 B.n632 B.n631 10.6151
R1974 B.n631 B.n88 10.6151
R1975 B.n627 B.n88 10.6151
R1976 B.n627 B.n626 10.6151
R1977 B.n626 B.n625 10.6151
R1978 B.n625 B.n90 10.6151
R1979 B.n621 B.n90 10.6151
R1980 B.n621 B.n620 10.6151
R1981 B.n620 B.n619 10.6151
R1982 B.n619 B.n92 10.6151
R1983 B.n615 B.n92 10.6151
R1984 B.n615 B.n614 10.6151
R1985 B.n614 B.n613 10.6151
R1986 B.n613 B.n94 10.6151
R1987 B.n609 B.n94 10.6151
R1988 B.n609 B.n608 10.6151
R1989 B.n608 B.n607 10.6151
R1990 B.n607 B.n96 10.6151
R1991 B.n603 B.n96 10.6151
R1992 B.n603 B.n602 10.6151
R1993 B.n602 B.n601 10.6151
R1994 B.n601 B.n98 10.6151
R1995 B.n597 B.n98 10.6151
R1996 B.n597 B.n596 10.6151
R1997 B.n596 B.n595 10.6151
R1998 B.n595 B.n100 10.6151
R1999 B.n591 B.n100 10.6151
R2000 B.n591 B.n590 10.6151
R2001 B.n590 B.n589 10.6151
R2002 B.n589 B.n102 10.6151
R2003 B.n585 B.n102 10.6151
R2004 B.n585 B.n584 10.6151
R2005 B.n584 B.n583 10.6151
R2006 B.n583 B.n104 10.6151
R2007 B.n579 B.n104 10.6151
R2008 B.n579 B.n578 10.6151
R2009 B.n578 B.n577 10.6151
R2010 B.n577 B.n106 10.6151
R2011 B.n573 B.n106 10.6151
R2012 B.n573 B.n572 10.6151
R2013 B.n572 B.n571 10.6151
R2014 B.n571 B.n108 10.6151
R2015 B.n567 B.n108 10.6151
R2016 B.n567 B.n566 10.6151
R2017 B.n566 B.n565 10.6151
R2018 B.n565 B.n110 10.6151
R2019 B.n561 B.n110 10.6151
R2020 B.n561 B.n560 10.6151
R2021 B.n560 B.n559 10.6151
R2022 B.n559 B.n112 10.6151
R2023 B.n555 B.n112 10.6151
R2024 B.n555 B.n554 10.6151
R2025 B.n554 B.n553 10.6151
R2026 B.n553 B.n114 10.6151
R2027 B.n549 B.n114 10.6151
R2028 B.n549 B.n548 10.6151
R2029 B.n548 B.n547 10.6151
R2030 B.n547 B.n116 10.6151
R2031 B.n543 B.n116 10.6151
R2032 B.n543 B.n542 10.6151
R2033 B.n542 B.n541 10.6151
R2034 B.n541 B.n118 10.6151
R2035 B.n537 B.n118 10.6151
R2036 B.n537 B.n536 10.6151
R2037 B.n536 B.n535 10.6151
R2038 B.n535 B.n120 10.6151
R2039 B.n531 B.n120 10.6151
R2040 B.n531 B.n530 10.6151
R2041 B.n530 B.n529 10.6151
R2042 B.n529 B.n122 10.6151
R2043 B.n525 B.n122 10.6151
R2044 B.n525 B.n524 10.6151
R2045 B.n524 B.n523 10.6151
R2046 B.n523 B.n124 10.6151
R2047 B.n519 B.n124 10.6151
R2048 B.n519 B.n518 10.6151
R2049 B.n518 B.n517 10.6151
R2050 B.n517 B.n126 10.6151
R2051 B.n513 B.n126 10.6151
R2052 B.n513 B.n512 10.6151
R2053 B.n512 B.n511 10.6151
R2054 B.n511 B.n128 10.6151
R2055 B.n507 B.n128 10.6151
R2056 B.n507 B.n506 10.6151
R2057 B.n506 B.n505 10.6151
R2058 B.n505 B.n130 10.6151
R2059 B.n501 B.n130 10.6151
R2060 B.n501 B.n500 10.6151
R2061 B.n500 B.n499 10.6151
R2062 B.n499 B.n132 10.6151
R2063 B.n495 B.n132 10.6151
R2064 B.n495 B.n494 10.6151
R2065 B.n494 B.n493 10.6151
R2066 B.n493 B.n134 10.6151
R2067 B.n489 B.n134 10.6151
R2068 B.n489 B.n488 10.6151
R2069 B.n488 B.n487 10.6151
R2070 B.n487 B.n136 10.6151
R2071 B.n483 B.n136 10.6151
R2072 B.n483 B.n482 10.6151
R2073 B.n482 B.n481 10.6151
R2074 B.n481 B.n138 10.6151
R2075 B.n477 B.n138 10.6151
R2076 B.n477 B.n476 10.6151
R2077 B.n476 B.n475 10.6151
R2078 B.n475 B.n140 10.6151
R2079 B.n471 B.n140 10.6151
R2080 B.n471 B.n470 10.6151
R2081 B.n470 B.n469 10.6151
R2082 B.n469 B.n142 10.6151
R2083 B.n465 B.n142 10.6151
R2084 B.n465 B.n464 10.6151
R2085 B.n464 B.n463 10.6151
R2086 B.n463 B.n144 10.6151
R2087 B.n459 B.n144 10.6151
R2088 B.n459 B.n458 10.6151
R2089 B.n458 B.n457 10.6151
R2090 B.n457 B.n146 10.6151
R2091 B.n453 B.n146 10.6151
R2092 B.n453 B.n452 10.6151
R2093 B.n452 B.n451 10.6151
R2094 B.n451 B.n148 10.6151
R2095 B.n447 B.n148 10.6151
R2096 B.n447 B.n446 10.6151
R2097 B.n225 B.n1 10.6151
R2098 B.n226 B.n225 10.6151
R2099 B.n227 B.n226 10.6151
R2100 B.n227 B.n222 10.6151
R2101 B.n231 B.n222 10.6151
R2102 B.n232 B.n231 10.6151
R2103 B.n233 B.n232 10.6151
R2104 B.n233 B.n220 10.6151
R2105 B.n237 B.n220 10.6151
R2106 B.n238 B.n237 10.6151
R2107 B.n239 B.n238 10.6151
R2108 B.n239 B.n218 10.6151
R2109 B.n243 B.n218 10.6151
R2110 B.n244 B.n243 10.6151
R2111 B.n245 B.n244 10.6151
R2112 B.n245 B.n216 10.6151
R2113 B.n249 B.n216 10.6151
R2114 B.n250 B.n249 10.6151
R2115 B.n251 B.n250 10.6151
R2116 B.n251 B.n214 10.6151
R2117 B.n255 B.n214 10.6151
R2118 B.n256 B.n255 10.6151
R2119 B.n257 B.n256 10.6151
R2120 B.n257 B.n212 10.6151
R2121 B.n261 B.n212 10.6151
R2122 B.n262 B.n261 10.6151
R2123 B.n263 B.n262 10.6151
R2124 B.n263 B.n210 10.6151
R2125 B.n267 B.n210 10.6151
R2126 B.n268 B.n267 10.6151
R2127 B.n269 B.n268 10.6151
R2128 B.n269 B.n208 10.6151
R2129 B.n273 B.n208 10.6151
R2130 B.n274 B.n273 10.6151
R2131 B.n275 B.n274 10.6151
R2132 B.n275 B.n206 10.6151
R2133 B.n279 B.n206 10.6151
R2134 B.n280 B.n279 10.6151
R2135 B.n281 B.n280 10.6151
R2136 B.n281 B.n204 10.6151
R2137 B.n285 B.n204 10.6151
R2138 B.n286 B.n285 10.6151
R2139 B.n287 B.n286 10.6151
R2140 B.n287 B.n202 10.6151
R2141 B.n291 B.n202 10.6151
R2142 B.n292 B.n291 10.6151
R2143 B.n293 B.n292 10.6151
R2144 B.n293 B.n200 10.6151
R2145 B.n297 B.n200 10.6151
R2146 B.n298 B.n297 10.6151
R2147 B.n299 B.n298 10.6151
R2148 B.n299 B.n198 10.6151
R2149 B.n303 B.n198 10.6151
R2150 B.n304 B.n303 10.6151
R2151 B.n305 B.n304 10.6151
R2152 B.n305 B.n196 10.6151
R2153 B.n309 B.n196 10.6151
R2154 B.n310 B.n309 10.6151
R2155 B.n311 B.n310 10.6151
R2156 B.n311 B.n194 10.6151
R2157 B.n315 B.n194 10.6151
R2158 B.n316 B.n315 10.6151
R2159 B.n317 B.n316 10.6151
R2160 B.n317 B.n192 10.6151
R2161 B.n321 B.n192 10.6151
R2162 B.n322 B.n321 10.6151
R2163 B.n323 B.n322 10.6151
R2164 B.n323 B.n190 10.6151
R2165 B.n328 B.n327 10.6151
R2166 B.n329 B.n328 10.6151
R2167 B.n329 B.n188 10.6151
R2168 B.n333 B.n188 10.6151
R2169 B.n334 B.n333 10.6151
R2170 B.n335 B.n334 10.6151
R2171 B.n335 B.n186 10.6151
R2172 B.n339 B.n186 10.6151
R2173 B.n340 B.n339 10.6151
R2174 B.n341 B.n340 10.6151
R2175 B.n341 B.n184 10.6151
R2176 B.n345 B.n184 10.6151
R2177 B.n346 B.n345 10.6151
R2178 B.n347 B.n346 10.6151
R2179 B.n347 B.n182 10.6151
R2180 B.n351 B.n182 10.6151
R2181 B.n352 B.n351 10.6151
R2182 B.n353 B.n352 10.6151
R2183 B.n353 B.n180 10.6151
R2184 B.n357 B.n180 10.6151
R2185 B.n358 B.n357 10.6151
R2186 B.n359 B.n358 10.6151
R2187 B.n359 B.n178 10.6151
R2188 B.n363 B.n178 10.6151
R2189 B.n364 B.n363 10.6151
R2190 B.n365 B.n364 10.6151
R2191 B.n365 B.n176 10.6151
R2192 B.n369 B.n176 10.6151
R2193 B.n370 B.n369 10.6151
R2194 B.n371 B.n370 10.6151
R2195 B.n371 B.n174 10.6151
R2196 B.n375 B.n174 10.6151
R2197 B.n376 B.n375 10.6151
R2198 B.n378 B.n170 10.6151
R2199 B.n382 B.n170 10.6151
R2200 B.n383 B.n382 10.6151
R2201 B.n384 B.n383 10.6151
R2202 B.n384 B.n168 10.6151
R2203 B.n388 B.n168 10.6151
R2204 B.n389 B.n388 10.6151
R2205 B.n393 B.n389 10.6151
R2206 B.n397 B.n166 10.6151
R2207 B.n398 B.n397 10.6151
R2208 B.n399 B.n398 10.6151
R2209 B.n399 B.n164 10.6151
R2210 B.n403 B.n164 10.6151
R2211 B.n404 B.n403 10.6151
R2212 B.n405 B.n404 10.6151
R2213 B.n405 B.n162 10.6151
R2214 B.n409 B.n162 10.6151
R2215 B.n410 B.n409 10.6151
R2216 B.n411 B.n410 10.6151
R2217 B.n411 B.n160 10.6151
R2218 B.n415 B.n160 10.6151
R2219 B.n416 B.n415 10.6151
R2220 B.n417 B.n416 10.6151
R2221 B.n417 B.n158 10.6151
R2222 B.n421 B.n158 10.6151
R2223 B.n422 B.n421 10.6151
R2224 B.n423 B.n422 10.6151
R2225 B.n423 B.n156 10.6151
R2226 B.n427 B.n156 10.6151
R2227 B.n428 B.n427 10.6151
R2228 B.n429 B.n428 10.6151
R2229 B.n429 B.n154 10.6151
R2230 B.n433 B.n154 10.6151
R2231 B.n434 B.n433 10.6151
R2232 B.n435 B.n434 10.6151
R2233 B.n435 B.n152 10.6151
R2234 B.n439 B.n152 10.6151
R2235 B.n440 B.n439 10.6151
R2236 B.n441 B.n440 10.6151
R2237 B.n441 B.n150 10.6151
R2238 B.n445 B.n150 10.6151
R2239 B.n877 B.n0 8.11757
R2240 B.n877 B.n1 8.11757
R2241 B.n721 B.n720 6.5566
R2242 B.n708 B.n62 6.5566
R2243 B.n378 B.n377 6.5566
R2244 B.n393 B.n392 6.5566
R2245 B.n722 B.n721 4.05904
R2246 B.n705 B.n62 4.05904
R2247 B.n377 B.n376 4.05904
R2248 B.n392 B.n166 4.05904
C0 VP VTAIL 8.21548f
C1 VDD1 VTAIL 7.87817f
C2 B w_n5150_n2818# 11.2576f
C3 B VN 1.48386f
C4 VDD2 VTAIL 7.94096f
C5 VP w_n5150_n2818# 11.452701f
C6 VP VN 8.68366f
C7 VDD1 w_n5150_n2818# 2.27873f
C8 VDD1 VN 0.153784f
C9 VDD2 w_n5150_n2818# 2.44587f
C10 VDD2 VN 7.26161f
C11 B VP 2.61746f
C12 VDD1 B 1.95724f
C13 VDD1 VP 7.75828f
C14 VDD2 B 2.09259f
C15 VDD2 VP 0.65248f
C16 VDD1 VDD2 2.42493f
C17 VTAIL w_n5150_n2818# 3.72737f
C18 VN VTAIL 8.20138f
C19 VN w_n5150_n2818# 10.7804f
C20 B VTAIL 4.53592f
C21 VDD2 VSUBS 2.519878f
C22 VDD1 VSUBS 3.24869f
C23 VTAIL VSUBS 1.46452f
C24 VN VSUBS 8.39597f
C25 VP VSUBS 4.766448f
C26 B VSUBS 6.164723f
C27 w_n5150_n2818# VSUBS 0.179529p
C28 B.n0 VSUBS 0.007671f
C29 B.n1 VSUBS 0.007671f
C30 B.n2 VSUBS 0.011346f
C31 B.n3 VSUBS 0.008694f
C32 B.n4 VSUBS 0.008694f
C33 B.n5 VSUBS 0.008694f
C34 B.n6 VSUBS 0.008694f
C35 B.n7 VSUBS 0.008694f
C36 B.n8 VSUBS 0.008694f
C37 B.n9 VSUBS 0.008694f
C38 B.n10 VSUBS 0.008694f
C39 B.n11 VSUBS 0.008694f
C40 B.n12 VSUBS 0.008694f
C41 B.n13 VSUBS 0.008694f
C42 B.n14 VSUBS 0.008694f
C43 B.n15 VSUBS 0.008694f
C44 B.n16 VSUBS 0.008694f
C45 B.n17 VSUBS 0.008694f
C46 B.n18 VSUBS 0.008694f
C47 B.n19 VSUBS 0.008694f
C48 B.n20 VSUBS 0.008694f
C49 B.n21 VSUBS 0.008694f
C50 B.n22 VSUBS 0.008694f
C51 B.n23 VSUBS 0.008694f
C52 B.n24 VSUBS 0.008694f
C53 B.n25 VSUBS 0.008694f
C54 B.n26 VSUBS 0.008694f
C55 B.n27 VSUBS 0.008694f
C56 B.n28 VSUBS 0.008694f
C57 B.n29 VSUBS 0.008694f
C58 B.n30 VSUBS 0.008694f
C59 B.n31 VSUBS 0.008694f
C60 B.n32 VSUBS 0.008694f
C61 B.n33 VSUBS 0.008694f
C62 B.n34 VSUBS 0.008694f
C63 B.n35 VSUBS 0.008694f
C64 B.n36 VSUBS 0.019074f
C65 B.n37 VSUBS 0.008694f
C66 B.n38 VSUBS 0.008694f
C67 B.n39 VSUBS 0.008694f
C68 B.n40 VSUBS 0.008694f
C69 B.n41 VSUBS 0.008694f
C70 B.n42 VSUBS 0.008694f
C71 B.n43 VSUBS 0.008694f
C72 B.n44 VSUBS 0.008694f
C73 B.n45 VSUBS 0.008694f
C74 B.n46 VSUBS 0.008694f
C75 B.n47 VSUBS 0.008694f
C76 B.n48 VSUBS 0.008694f
C77 B.n49 VSUBS 0.008694f
C78 B.n50 VSUBS 0.008694f
C79 B.n51 VSUBS 0.008694f
C80 B.n52 VSUBS 0.008694f
C81 B.n53 VSUBS 0.008694f
C82 B.t1 VSUBS 0.188393f
C83 B.t2 VSUBS 0.239582f
C84 B.t0 VSUBS 2.09075f
C85 B.n54 VSUBS 0.386007f
C86 B.n55 VSUBS 0.269433f
C87 B.n56 VSUBS 0.008694f
C88 B.n57 VSUBS 0.008694f
C89 B.n58 VSUBS 0.008694f
C90 B.n59 VSUBS 0.008694f
C91 B.t7 VSUBS 0.188396f
C92 B.t8 VSUBS 0.239585f
C93 B.t6 VSUBS 2.09075f
C94 B.n60 VSUBS 0.386005f
C95 B.n61 VSUBS 0.26943f
C96 B.n62 VSUBS 0.020144f
C97 B.n63 VSUBS 0.008694f
C98 B.n64 VSUBS 0.008694f
C99 B.n65 VSUBS 0.008694f
C100 B.n66 VSUBS 0.008694f
C101 B.n67 VSUBS 0.008694f
C102 B.n68 VSUBS 0.008694f
C103 B.n69 VSUBS 0.008694f
C104 B.n70 VSUBS 0.008694f
C105 B.n71 VSUBS 0.008694f
C106 B.n72 VSUBS 0.008694f
C107 B.n73 VSUBS 0.008694f
C108 B.n74 VSUBS 0.008694f
C109 B.n75 VSUBS 0.008694f
C110 B.n76 VSUBS 0.008694f
C111 B.n77 VSUBS 0.008694f
C112 B.n78 VSUBS 0.008694f
C113 B.n79 VSUBS 0.020561f
C114 B.n80 VSUBS 0.008694f
C115 B.n81 VSUBS 0.008694f
C116 B.n82 VSUBS 0.008694f
C117 B.n83 VSUBS 0.008694f
C118 B.n84 VSUBS 0.008694f
C119 B.n85 VSUBS 0.008694f
C120 B.n86 VSUBS 0.008694f
C121 B.n87 VSUBS 0.008694f
C122 B.n88 VSUBS 0.008694f
C123 B.n89 VSUBS 0.008694f
C124 B.n90 VSUBS 0.008694f
C125 B.n91 VSUBS 0.008694f
C126 B.n92 VSUBS 0.008694f
C127 B.n93 VSUBS 0.008694f
C128 B.n94 VSUBS 0.008694f
C129 B.n95 VSUBS 0.008694f
C130 B.n96 VSUBS 0.008694f
C131 B.n97 VSUBS 0.008694f
C132 B.n98 VSUBS 0.008694f
C133 B.n99 VSUBS 0.008694f
C134 B.n100 VSUBS 0.008694f
C135 B.n101 VSUBS 0.008694f
C136 B.n102 VSUBS 0.008694f
C137 B.n103 VSUBS 0.008694f
C138 B.n104 VSUBS 0.008694f
C139 B.n105 VSUBS 0.008694f
C140 B.n106 VSUBS 0.008694f
C141 B.n107 VSUBS 0.008694f
C142 B.n108 VSUBS 0.008694f
C143 B.n109 VSUBS 0.008694f
C144 B.n110 VSUBS 0.008694f
C145 B.n111 VSUBS 0.008694f
C146 B.n112 VSUBS 0.008694f
C147 B.n113 VSUBS 0.008694f
C148 B.n114 VSUBS 0.008694f
C149 B.n115 VSUBS 0.008694f
C150 B.n116 VSUBS 0.008694f
C151 B.n117 VSUBS 0.008694f
C152 B.n118 VSUBS 0.008694f
C153 B.n119 VSUBS 0.008694f
C154 B.n120 VSUBS 0.008694f
C155 B.n121 VSUBS 0.008694f
C156 B.n122 VSUBS 0.008694f
C157 B.n123 VSUBS 0.008694f
C158 B.n124 VSUBS 0.008694f
C159 B.n125 VSUBS 0.008694f
C160 B.n126 VSUBS 0.008694f
C161 B.n127 VSUBS 0.008694f
C162 B.n128 VSUBS 0.008694f
C163 B.n129 VSUBS 0.008694f
C164 B.n130 VSUBS 0.008694f
C165 B.n131 VSUBS 0.008694f
C166 B.n132 VSUBS 0.008694f
C167 B.n133 VSUBS 0.008694f
C168 B.n134 VSUBS 0.008694f
C169 B.n135 VSUBS 0.008694f
C170 B.n136 VSUBS 0.008694f
C171 B.n137 VSUBS 0.008694f
C172 B.n138 VSUBS 0.008694f
C173 B.n139 VSUBS 0.008694f
C174 B.n140 VSUBS 0.008694f
C175 B.n141 VSUBS 0.008694f
C176 B.n142 VSUBS 0.008694f
C177 B.n143 VSUBS 0.008694f
C178 B.n144 VSUBS 0.008694f
C179 B.n145 VSUBS 0.008694f
C180 B.n146 VSUBS 0.008694f
C181 B.n147 VSUBS 0.008694f
C182 B.n148 VSUBS 0.008694f
C183 B.n149 VSUBS 0.019074f
C184 B.n150 VSUBS 0.008694f
C185 B.n151 VSUBS 0.008694f
C186 B.n152 VSUBS 0.008694f
C187 B.n153 VSUBS 0.008694f
C188 B.n154 VSUBS 0.008694f
C189 B.n155 VSUBS 0.008694f
C190 B.n156 VSUBS 0.008694f
C191 B.n157 VSUBS 0.008694f
C192 B.n158 VSUBS 0.008694f
C193 B.n159 VSUBS 0.008694f
C194 B.n160 VSUBS 0.008694f
C195 B.n161 VSUBS 0.008694f
C196 B.n162 VSUBS 0.008694f
C197 B.n163 VSUBS 0.008694f
C198 B.n164 VSUBS 0.008694f
C199 B.n165 VSUBS 0.008694f
C200 B.n166 VSUBS 0.006009f
C201 B.n167 VSUBS 0.008694f
C202 B.n168 VSUBS 0.008694f
C203 B.n169 VSUBS 0.008694f
C204 B.n170 VSUBS 0.008694f
C205 B.n171 VSUBS 0.008694f
C206 B.t11 VSUBS 0.188393f
C207 B.t10 VSUBS 0.239582f
C208 B.t9 VSUBS 2.09075f
C209 B.n172 VSUBS 0.386007f
C210 B.n173 VSUBS 0.269433f
C211 B.n174 VSUBS 0.008694f
C212 B.n175 VSUBS 0.008694f
C213 B.n176 VSUBS 0.008694f
C214 B.n177 VSUBS 0.008694f
C215 B.n178 VSUBS 0.008694f
C216 B.n179 VSUBS 0.008694f
C217 B.n180 VSUBS 0.008694f
C218 B.n181 VSUBS 0.008694f
C219 B.n182 VSUBS 0.008694f
C220 B.n183 VSUBS 0.008694f
C221 B.n184 VSUBS 0.008694f
C222 B.n185 VSUBS 0.008694f
C223 B.n186 VSUBS 0.008694f
C224 B.n187 VSUBS 0.008694f
C225 B.n188 VSUBS 0.008694f
C226 B.n189 VSUBS 0.008694f
C227 B.n190 VSUBS 0.019074f
C228 B.n191 VSUBS 0.008694f
C229 B.n192 VSUBS 0.008694f
C230 B.n193 VSUBS 0.008694f
C231 B.n194 VSUBS 0.008694f
C232 B.n195 VSUBS 0.008694f
C233 B.n196 VSUBS 0.008694f
C234 B.n197 VSUBS 0.008694f
C235 B.n198 VSUBS 0.008694f
C236 B.n199 VSUBS 0.008694f
C237 B.n200 VSUBS 0.008694f
C238 B.n201 VSUBS 0.008694f
C239 B.n202 VSUBS 0.008694f
C240 B.n203 VSUBS 0.008694f
C241 B.n204 VSUBS 0.008694f
C242 B.n205 VSUBS 0.008694f
C243 B.n206 VSUBS 0.008694f
C244 B.n207 VSUBS 0.008694f
C245 B.n208 VSUBS 0.008694f
C246 B.n209 VSUBS 0.008694f
C247 B.n210 VSUBS 0.008694f
C248 B.n211 VSUBS 0.008694f
C249 B.n212 VSUBS 0.008694f
C250 B.n213 VSUBS 0.008694f
C251 B.n214 VSUBS 0.008694f
C252 B.n215 VSUBS 0.008694f
C253 B.n216 VSUBS 0.008694f
C254 B.n217 VSUBS 0.008694f
C255 B.n218 VSUBS 0.008694f
C256 B.n219 VSUBS 0.008694f
C257 B.n220 VSUBS 0.008694f
C258 B.n221 VSUBS 0.008694f
C259 B.n222 VSUBS 0.008694f
C260 B.n223 VSUBS 0.008694f
C261 B.n224 VSUBS 0.008694f
C262 B.n225 VSUBS 0.008694f
C263 B.n226 VSUBS 0.008694f
C264 B.n227 VSUBS 0.008694f
C265 B.n228 VSUBS 0.008694f
C266 B.n229 VSUBS 0.008694f
C267 B.n230 VSUBS 0.008694f
C268 B.n231 VSUBS 0.008694f
C269 B.n232 VSUBS 0.008694f
C270 B.n233 VSUBS 0.008694f
C271 B.n234 VSUBS 0.008694f
C272 B.n235 VSUBS 0.008694f
C273 B.n236 VSUBS 0.008694f
C274 B.n237 VSUBS 0.008694f
C275 B.n238 VSUBS 0.008694f
C276 B.n239 VSUBS 0.008694f
C277 B.n240 VSUBS 0.008694f
C278 B.n241 VSUBS 0.008694f
C279 B.n242 VSUBS 0.008694f
C280 B.n243 VSUBS 0.008694f
C281 B.n244 VSUBS 0.008694f
C282 B.n245 VSUBS 0.008694f
C283 B.n246 VSUBS 0.008694f
C284 B.n247 VSUBS 0.008694f
C285 B.n248 VSUBS 0.008694f
C286 B.n249 VSUBS 0.008694f
C287 B.n250 VSUBS 0.008694f
C288 B.n251 VSUBS 0.008694f
C289 B.n252 VSUBS 0.008694f
C290 B.n253 VSUBS 0.008694f
C291 B.n254 VSUBS 0.008694f
C292 B.n255 VSUBS 0.008694f
C293 B.n256 VSUBS 0.008694f
C294 B.n257 VSUBS 0.008694f
C295 B.n258 VSUBS 0.008694f
C296 B.n259 VSUBS 0.008694f
C297 B.n260 VSUBS 0.008694f
C298 B.n261 VSUBS 0.008694f
C299 B.n262 VSUBS 0.008694f
C300 B.n263 VSUBS 0.008694f
C301 B.n264 VSUBS 0.008694f
C302 B.n265 VSUBS 0.008694f
C303 B.n266 VSUBS 0.008694f
C304 B.n267 VSUBS 0.008694f
C305 B.n268 VSUBS 0.008694f
C306 B.n269 VSUBS 0.008694f
C307 B.n270 VSUBS 0.008694f
C308 B.n271 VSUBS 0.008694f
C309 B.n272 VSUBS 0.008694f
C310 B.n273 VSUBS 0.008694f
C311 B.n274 VSUBS 0.008694f
C312 B.n275 VSUBS 0.008694f
C313 B.n276 VSUBS 0.008694f
C314 B.n277 VSUBS 0.008694f
C315 B.n278 VSUBS 0.008694f
C316 B.n279 VSUBS 0.008694f
C317 B.n280 VSUBS 0.008694f
C318 B.n281 VSUBS 0.008694f
C319 B.n282 VSUBS 0.008694f
C320 B.n283 VSUBS 0.008694f
C321 B.n284 VSUBS 0.008694f
C322 B.n285 VSUBS 0.008694f
C323 B.n286 VSUBS 0.008694f
C324 B.n287 VSUBS 0.008694f
C325 B.n288 VSUBS 0.008694f
C326 B.n289 VSUBS 0.008694f
C327 B.n290 VSUBS 0.008694f
C328 B.n291 VSUBS 0.008694f
C329 B.n292 VSUBS 0.008694f
C330 B.n293 VSUBS 0.008694f
C331 B.n294 VSUBS 0.008694f
C332 B.n295 VSUBS 0.008694f
C333 B.n296 VSUBS 0.008694f
C334 B.n297 VSUBS 0.008694f
C335 B.n298 VSUBS 0.008694f
C336 B.n299 VSUBS 0.008694f
C337 B.n300 VSUBS 0.008694f
C338 B.n301 VSUBS 0.008694f
C339 B.n302 VSUBS 0.008694f
C340 B.n303 VSUBS 0.008694f
C341 B.n304 VSUBS 0.008694f
C342 B.n305 VSUBS 0.008694f
C343 B.n306 VSUBS 0.008694f
C344 B.n307 VSUBS 0.008694f
C345 B.n308 VSUBS 0.008694f
C346 B.n309 VSUBS 0.008694f
C347 B.n310 VSUBS 0.008694f
C348 B.n311 VSUBS 0.008694f
C349 B.n312 VSUBS 0.008694f
C350 B.n313 VSUBS 0.008694f
C351 B.n314 VSUBS 0.008694f
C352 B.n315 VSUBS 0.008694f
C353 B.n316 VSUBS 0.008694f
C354 B.n317 VSUBS 0.008694f
C355 B.n318 VSUBS 0.008694f
C356 B.n319 VSUBS 0.008694f
C357 B.n320 VSUBS 0.008694f
C358 B.n321 VSUBS 0.008694f
C359 B.n322 VSUBS 0.008694f
C360 B.n323 VSUBS 0.008694f
C361 B.n324 VSUBS 0.008694f
C362 B.n325 VSUBS 0.019074f
C363 B.n326 VSUBS 0.020561f
C364 B.n327 VSUBS 0.020561f
C365 B.n328 VSUBS 0.008694f
C366 B.n329 VSUBS 0.008694f
C367 B.n330 VSUBS 0.008694f
C368 B.n331 VSUBS 0.008694f
C369 B.n332 VSUBS 0.008694f
C370 B.n333 VSUBS 0.008694f
C371 B.n334 VSUBS 0.008694f
C372 B.n335 VSUBS 0.008694f
C373 B.n336 VSUBS 0.008694f
C374 B.n337 VSUBS 0.008694f
C375 B.n338 VSUBS 0.008694f
C376 B.n339 VSUBS 0.008694f
C377 B.n340 VSUBS 0.008694f
C378 B.n341 VSUBS 0.008694f
C379 B.n342 VSUBS 0.008694f
C380 B.n343 VSUBS 0.008694f
C381 B.n344 VSUBS 0.008694f
C382 B.n345 VSUBS 0.008694f
C383 B.n346 VSUBS 0.008694f
C384 B.n347 VSUBS 0.008694f
C385 B.n348 VSUBS 0.008694f
C386 B.n349 VSUBS 0.008694f
C387 B.n350 VSUBS 0.008694f
C388 B.n351 VSUBS 0.008694f
C389 B.n352 VSUBS 0.008694f
C390 B.n353 VSUBS 0.008694f
C391 B.n354 VSUBS 0.008694f
C392 B.n355 VSUBS 0.008694f
C393 B.n356 VSUBS 0.008694f
C394 B.n357 VSUBS 0.008694f
C395 B.n358 VSUBS 0.008694f
C396 B.n359 VSUBS 0.008694f
C397 B.n360 VSUBS 0.008694f
C398 B.n361 VSUBS 0.008694f
C399 B.n362 VSUBS 0.008694f
C400 B.n363 VSUBS 0.008694f
C401 B.n364 VSUBS 0.008694f
C402 B.n365 VSUBS 0.008694f
C403 B.n366 VSUBS 0.008694f
C404 B.n367 VSUBS 0.008694f
C405 B.n368 VSUBS 0.008694f
C406 B.n369 VSUBS 0.008694f
C407 B.n370 VSUBS 0.008694f
C408 B.n371 VSUBS 0.008694f
C409 B.n372 VSUBS 0.008694f
C410 B.n373 VSUBS 0.008694f
C411 B.n374 VSUBS 0.008694f
C412 B.n375 VSUBS 0.008694f
C413 B.n376 VSUBS 0.006009f
C414 B.n377 VSUBS 0.020144f
C415 B.n378 VSUBS 0.007032f
C416 B.n379 VSUBS 0.008694f
C417 B.n380 VSUBS 0.008694f
C418 B.n381 VSUBS 0.008694f
C419 B.n382 VSUBS 0.008694f
C420 B.n383 VSUBS 0.008694f
C421 B.n384 VSUBS 0.008694f
C422 B.n385 VSUBS 0.008694f
C423 B.n386 VSUBS 0.008694f
C424 B.n387 VSUBS 0.008694f
C425 B.n388 VSUBS 0.008694f
C426 B.n389 VSUBS 0.008694f
C427 B.t5 VSUBS 0.188396f
C428 B.t4 VSUBS 0.239585f
C429 B.t3 VSUBS 2.09075f
C430 B.n390 VSUBS 0.386005f
C431 B.n391 VSUBS 0.26943f
C432 B.n392 VSUBS 0.020144f
C433 B.n393 VSUBS 0.007032f
C434 B.n394 VSUBS 0.008694f
C435 B.n395 VSUBS 0.008694f
C436 B.n396 VSUBS 0.008694f
C437 B.n397 VSUBS 0.008694f
C438 B.n398 VSUBS 0.008694f
C439 B.n399 VSUBS 0.008694f
C440 B.n400 VSUBS 0.008694f
C441 B.n401 VSUBS 0.008694f
C442 B.n402 VSUBS 0.008694f
C443 B.n403 VSUBS 0.008694f
C444 B.n404 VSUBS 0.008694f
C445 B.n405 VSUBS 0.008694f
C446 B.n406 VSUBS 0.008694f
C447 B.n407 VSUBS 0.008694f
C448 B.n408 VSUBS 0.008694f
C449 B.n409 VSUBS 0.008694f
C450 B.n410 VSUBS 0.008694f
C451 B.n411 VSUBS 0.008694f
C452 B.n412 VSUBS 0.008694f
C453 B.n413 VSUBS 0.008694f
C454 B.n414 VSUBS 0.008694f
C455 B.n415 VSUBS 0.008694f
C456 B.n416 VSUBS 0.008694f
C457 B.n417 VSUBS 0.008694f
C458 B.n418 VSUBS 0.008694f
C459 B.n419 VSUBS 0.008694f
C460 B.n420 VSUBS 0.008694f
C461 B.n421 VSUBS 0.008694f
C462 B.n422 VSUBS 0.008694f
C463 B.n423 VSUBS 0.008694f
C464 B.n424 VSUBS 0.008694f
C465 B.n425 VSUBS 0.008694f
C466 B.n426 VSUBS 0.008694f
C467 B.n427 VSUBS 0.008694f
C468 B.n428 VSUBS 0.008694f
C469 B.n429 VSUBS 0.008694f
C470 B.n430 VSUBS 0.008694f
C471 B.n431 VSUBS 0.008694f
C472 B.n432 VSUBS 0.008694f
C473 B.n433 VSUBS 0.008694f
C474 B.n434 VSUBS 0.008694f
C475 B.n435 VSUBS 0.008694f
C476 B.n436 VSUBS 0.008694f
C477 B.n437 VSUBS 0.008694f
C478 B.n438 VSUBS 0.008694f
C479 B.n439 VSUBS 0.008694f
C480 B.n440 VSUBS 0.008694f
C481 B.n441 VSUBS 0.008694f
C482 B.n442 VSUBS 0.008694f
C483 B.n443 VSUBS 0.008694f
C484 B.n444 VSUBS 0.020561f
C485 B.n445 VSUBS 0.019492f
C486 B.n446 VSUBS 0.020144f
C487 B.n447 VSUBS 0.008694f
C488 B.n448 VSUBS 0.008694f
C489 B.n449 VSUBS 0.008694f
C490 B.n450 VSUBS 0.008694f
C491 B.n451 VSUBS 0.008694f
C492 B.n452 VSUBS 0.008694f
C493 B.n453 VSUBS 0.008694f
C494 B.n454 VSUBS 0.008694f
C495 B.n455 VSUBS 0.008694f
C496 B.n456 VSUBS 0.008694f
C497 B.n457 VSUBS 0.008694f
C498 B.n458 VSUBS 0.008694f
C499 B.n459 VSUBS 0.008694f
C500 B.n460 VSUBS 0.008694f
C501 B.n461 VSUBS 0.008694f
C502 B.n462 VSUBS 0.008694f
C503 B.n463 VSUBS 0.008694f
C504 B.n464 VSUBS 0.008694f
C505 B.n465 VSUBS 0.008694f
C506 B.n466 VSUBS 0.008694f
C507 B.n467 VSUBS 0.008694f
C508 B.n468 VSUBS 0.008694f
C509 B.n469 VSUBS 0.008694f
C510 B.n470 VSUBS 0.008694f
C511 B.n471 VSUBS 0.008694f
C512 B.n472 VSUBS 0.008694f
C513 B.n473 VSUBS 0.008694f
C514 B.n474 VSUBS 0.008694f
C515 B.n475 VSUBS 0.008694f
C516 B.n476 VSUBS 0.008694f
C517 B.n477 VSUBS 0.008694f
C518 B.n478 VSUBS 0.008694f
C519 B.n479 VSUBS 0.008694f
C520 B.n480 VSUBS 0.008694f
C521 B.n481 VSUBS 0.008694f
C522 B.n482 VSUBS 0.008694f
C523 B.n483 VSUBS 0.008694f
C524 B.n484 VSUBS 0.008694f
C525 B.n485 VSUBS 0.008694f
C526 B.n486 VSUBS 0.008694f
C527 B.n487 VSUBS 0.008694f
C528 B.n488 VSUBS 0.008694f
C529 B.n489 VSUBS 0.008694f
C530 B.n490 VSUBS 0.008694f
C531 B.n491 VSUBS 0.008694f
C532 B.n492 VSUBS 0.008694f
C533 B.n493 VSUBS 0.008694f
C534 B.n494 VSUBS 0.008694f
C535 B.n495 VSUBS 0.008694f
C536 B.n496 VSUBS 0.008694f
C537 B.n497 VSUBS 0.008694f
C538 B.n498 VSUBS 0.008694f
C539 B.n499 VSUBS 0.008694f
C540 B.n500 VSUBS 0.008694f
C541 B.n501 VSUBS 0.008694f
C542 B.n502 VSUBS 0.008694f
C543 B.n503 VSUBS 0.008694f
C544 B.n504 VSUBS 0.008694f
C545 B.n505 VSUBS 0.008694f
C546 B.n506 VSUBS 0.008694f
C547 B.n507 VSUBS 0.008694f
C548 B.n508 VSUBS 0.008694f
C549 B.n509 VSUBS 0.008694f
C550 B.n510 VSUBS 0.008694f
C551 B.n511 VSUBS 0.008694f
C552 B.n512 VSUBS 0.008694f
C553 B.n513 VSUBS 0.008694f
C554 B.n514 VSUBS 0.008694f
C555 B.n515 VSUBS 0.008694f
C556 B.n516 VSUBS 0.008694f
C557 B.n517 VSUBS 0.008694f
C558 B.n518 VSUBS 0.008694f
C559 B.n519 VSUBS 0.008694f
C560 B.n520 VSUBS 0.008694f
C561 B.n521 VSUBS 0.008694f
C562 B.n522 VSUBS 0.008694f
C563 B.n523 VSUBS 0.008694f
C564 B.n524 VSUBS 0.008694f
C565 B.n525 VSUBS 0.008694f
C566 B.n526 VSUBS 0.008694f
C567 B.n527 VSUBS 0.008694f
C568 B.n528 VSUBS 0.008694f
C569 B.n529 VSUBS 0.008694f
C570 B.n530 VSUBS 0.008694f
C571 B.n531 VSUBS 0.008694f
C572 B.n532 VSUBS 0.008694f
C573 B.n533 VSUBS 0.008694f
C574 B.n534 VSUBS 0.008694f
C575 B.n535 VSUBS 0.008694f
C576 B.n536 VSUBS 0.008694f
C577 B.n537 VSUBS 0.008694f
C578 B.n538 VSUBS 0.008694f
C579 B.n539 VSUBS 0.008694f
C580 B.n540 VSUBS 0.008694f
C581 B.n541 VSUBS 0.008694f
C582 B.n542 VSUBS 0.008694f
C583 B.n543 VSUBS 0.008694f
C584 B.n544 VSUBS 0.008694f
C585 B.n545 VSUBS 0.008694f
C586 B.n546 VSUBS 0.008694f
C587 B.n547 VSUBS 0.008694f
C588 B.n548 VSUBS 0.008694f
C589 B.n549 VSUBS 0.008694f
C590 B.n550 VSUBS 0.008694f
C591 B.n551 VSUBS 0.008694f
C592 B.n552 VSUBS 0.008694f
C593 B.n553 VSUBS 0.008694f
C594 B.n554 VSUBS 0.008694f
C595 B.n555 VSUBS 0.008694f
C596 B.n556 VSUBS 0.008694f
C597 B.n557 VSUBS 0.008694f
C598 B.n558 VSUBS 0.008694f
C599 B.n559 VSUBS 0.008694f
C600 B.n560 VSUBS 0.008694f
C601 B.n561 VSUBS 0.008694f
C602 B.n562 VSUBS 0.008694f
C603 B.n563 VSUBS 0.008694f
C604 B.n564 VSUBS 0.008694f
C605 B.n565 VSUBS 0.008694f
C606 B.n566 VSUBS 0.008694f
C607 B.n567 VSUBS 0.008694f
C608 B.n568 VSUBS 0.008694f
C609 B.n569 VSUBS 0.008694f
C610 B.n570 VSUBS 0.008694f
C611 B.n571 VSUBS 0.008694f
C612 B.n572 VSUBS 0.008694f
C613 B.n573 VSUBS 0.008694f
C614 B.n574 VSUBS 0.008694f
C615 B.n575 VSUBS 0.008694f
C616 B.n576 VSUBS 0.008694f
C617 B.n577 VSUBS 0.008694f
C618 B.n578 VSUBS 0.008694f
C619 B.n579 VSUBS 0.008694f
C620 B.n580 VSUBS 0.008694f
C621 B.n581 VSUBS 0.008694f
C622 B.n582 VSUBS 0.008694f
C623 B.n583 VSUBS 0.008694f
C624 B.n584 VSUBS 0.008694f
C625 B.n585 VSUBS 0.008694f
C626 B.n586 VSUBS 0.008694f
C627 B.n587 VSUBS 0.008694f
C628 B.n588 VSUBS 0.008694f
C629 B.n589 VSUBS 0.008694f
C630 B.n590 VSUBS 0.008694f
C631 B.n591 VSUBS 0.008694f
C632 B.n592 VSUBS 0.008694f
C633 B.n593 VSUBS 0.008694f
C634 B.n594 VSUBS 0.008694f
C635 B.n595 VSUBS 0.008694f
C636 B.n596 VSUBS 0.008694f
C637 B.n597 VSUBS 0.008694f
C638 B.n598 VSUBS 0.008694f
C639 B.n599 VSUBS 0.008694f
C640 B.n600 VSUBS 0.008694f
C641 B.n601 VSUBS 0.008694f
C642 B.n602 VSUBS 0.008694f
C643 B.n603 VSUBS 0.008694f
C644 B.n604 VSUBS 0.008694f
C645 B.n605 VSUBS 0.008694f
C646 B.n606 VSUBS 0.008694f
C647 B.n607 VSUBS 0.008694f
C648 B.n608 VSUBS 0.008694f
C649 B.n609 VSUBS 0.008694f
C650 B.n610 VSUBS 0.008694f
C651 B.n611 VSUBS 0.008694f
C652 B.n612 VSUBS 0.008694f
C653 B.n613 VSUBS 0.008694f
C654 B.n614 VSUBS 0.008694f
C655 B.n615 VSUBS 0.008694f
C656 B.n616 VSUBS 0.008694f
C657 B.n617 VSUBS 0.008694f
C658 B.n618 VSUBS 0.008694f
C659 B.n619 VSUBS 0.008694f
C660 B.n620 VSUBS 0.008694f
C661 B.n621 VSUBS 0.008694f
C662 B.n622 VSUBS 0.008694f
C663 B.n623 VSUBS 0.008694f
C664 B.n624 VSUBS 0.008694f
C665 B.n625 VSUBS 0.008694f
C666 B.n626 VSUBS 0.008694f
C667 B.n627 VSUBS 0.008694f
C668 B.n628 VSUBS 0.008694f
C669 B.n629 VSUBS 0.008694f
C670 B.n630 VSUBS 0.008694f
C671 B.n631 VSUBS 0.008694f
C672 B.n632 VSUBS 0.008694f
C673 B.n633 VSUBS 0.008694f
C674 B.n634 VSUBS 0.008694f
C675 B.n635 VSUBS 0.008694f
C676 B.n636 VSUBS 0.008694f
C677 B.n637 VSUBS 0.008694f
C678 B.n638 VSUBS 0.008694f
C679 B.n639 VSUBS 0.008694f
C680 B.n640 VSUBS 0.008694f
C681 B.n641 VSUBS 0.008694f
C682 B.n642 VSUBS 0.008694f
C683 B.n643 VSUBS 0.008694f
C684 B.n644 VSUBS 0.008694f
C685 B.n645 VSUBS 0.008694f
C686 B.n646 VSUBS 0.008694f
C687 B.n647 VSUBS 0.008694f
C688 B.n648 VSUBS 0.008694f
C689 B.n649 VSUBS 0.008694f
C690 B.n650 VSUBS 0.008694f
C691 B.n651 VSUBS 0.008694f
C692 B.n652 VSUBS 0.008694f
C693 B.n653 VSUBS 0.008694f
C694 B.n654 VSUBS 0.019074f
C695 B.n655 VSUBS 0.019074f
C696 B.n656 VSUBS 0.020561f
C697 B.n657 VSUBS 0.008694f
C698 B.n658 VSUBS 0.008694f
C699 B.n659 VSUBS 0.008694f
C700 B.n660 VSUBS 0.008694f
C701 B.n661 VSUBS 0.008694f
C702 B.n662 VSUBS 0.008694f
C703 B.n663 VSUBS 0.008694f
C704 B.n664 VSUBS 0.008694f
C705 B.n665 VSUBS 0.008694f
C706 B.n666 VSUBS 0.008694f
C707 B.n667 VSUBS 0.008694f
C708 B.n668 VSUBS 0.008694f
C709 B.n669 VSUBS 0.008694f
C710 B.n670 VSUBS 0.008694f
C711 B.n671 VSUBS 0.008694f
C712 B.n672 VSUBS 0.008694f
C713 B.n673 VSUBS 0.008694f
C714 B.n674 VSUBS 0.008694f
C715 B.n675 VSUBS 0.008694f
C716 B.n676 VSUBS 0.008694f
C717 B.n677 VSUBS 0.008694f
C718 B.n678 VSUBS 0.008694f
C719 B.n679 VSUBS 0.008694f
C720 B.n680 VSUBS 0.008694f
C721 B.n681 VSUBS 0.008694f
C722 B.n682 VSUBS 0.008694f
C723 B.n683 VSUBS 0.008694f
C724 B.n684 VSUBS 0.008694f
C725 B.n685 VSUBS 0.008694f
C726 B.n686 VSUBS 0.008694f
C727 B.n687 VSUBS 0.008694f
C728 B.n688 VSUBS 0.008694f
C729 B.n689 VSUBS 0.008694f
C730 B.n690 VSUBS 0.008694f
C731 B.n691 VSUBS 0.008694f
C732 B.n692 VSUBS 0.008694f
C733 B.n693 VSUBS 0.008694f
C734 B.n694 VSUBS 0.008694f
C735 B.n695 VSUBS 0.008694f
C736 B.n696 VSUBS 0.008694f
C737 B.n697 VSUBS 0.008694f
C738 B.n698 VSUBS 0.008694f
C739 B.n699 VSUBS 0.008694f
C740 B.n700 VSUBS 0.008694f
C741 B.n701 VSUBS 0.008694f
C742 B.n702 VSUBS 0.008694f
C743 B.n703 VSUBS 0.008694f
C744 B.n704 VSUBS 0.008694f
C745 B.n705 VSUBS 0.006009f
C746 B.n706 VSUBS 0.008694f
C747 B.n707 VSUBS 0.008694f
C748 B.n708 VSUBS 0.007032f
C749 B.n709 VSUBS 0.008694f
C750 B.n710 VSUBS 0.008694f
C751 B.n711 VSUBS 0.008694f
C752 B.n712 VSUBS 0.008694f
C753 B.n713 VSUBS 0.008694f
C754 B.n714 VSUBS 0.008694f
C755 B.n715 VSUBS 0.008694f
C756 B.n716 VSUBS 0.008694f
C757 B.n717 VSUBS 0.008694f
C758 B.n718 VSUBS 0.008694f
C759 B.n719 VSUBS 0.008694f
C760 B.n720 VSUBS 0.007032f
C761 B.n721 VSUBS 0.020144f
C762 B.n722 VSUBS 0.006009f
C763 B.n723 VSUBS 0.008694f
C764 B.n724 VSUBS 0.008694f
C765 B.n725 VSUBS 0.008694f
C766 B.n726 VSUBS 0.008694f
C767 B.n727 VSUBS 0.008694f
C768 B.n728 VSUBS 0.008694f
C769 B.n729 VSUBS 0.008694f
C770 B.n730 VSUBS 0.008694f
C771 B.n731 VSUBS 0.008694f
C772 B.n732 VSUBS 0.008694f
C773 B.n733 VSUBS 0.008694f
C774 B.n734 VSUBS 0.008694f
C775 B.n735 VSUBS 0.008694f
C776 B.n736 VSUBS 0.008694f
C777 B.n737 VSUBS 0.008694f
C778 B.n738 VSUBS 0.008694f
C779 B.n739 VSUBS 0.008694f
C780 B.n740 VSUBS 0.008694f
C781 B.n741 VSUBS 0.008694f
C782 B.n742 VSUBS 0.008694f
C783 B.n743 VSUBS 0.008694f
C784 B.n744 VSUBS 0.008694f
C785 B.n745 VSUBS 0.008694f
C786 B.n746 VSUBS 0.008694f
C787 B.n747 VSUBS 0.008694f
C788 B.n748 VSUBS 0.008694f
C789 B.n749 VSUBS 0.008694f
C790 B.n750 VSUBS 0.008694f
C791 B.n751 VSUBS 0.008694f
C792 B.n752 VSUBS 0.008694f
C793 B.n753 VSUBS 0.008694f
C794 B.n754 VSUBS 0.008694f
C795 B.n755 VSUBS 0.008694f
C796 B.n756 VSUBS 0.008694f
C797 B.n757 VSUBS 0.008694f
C798 B.n758 VSUBS 0.008694f
C799 B.n759 VSUBS 0.008694f
C800 B.n760 VSUBS 0.008694f
C801 B.n761 VSUBS 0.008694f
C802 B.n762 VSUBS 0.008694f
C803 B.n763 VSUBS 0.008694f
C804 B.n764 VSUBS 0.008694f
C805 B.n765 VSUBS 0.008694f
C806 B.n766 VSUBS 0.008694f
C807 B.n767 VSUBS 0.008694f
C808 B.n768 VSUBS 0.008694f
C809 B.n769 VSUBS 0.008694f
C810 B.n770 VSUBS 0.008694f
C811 B.n771 VSUBS 0.020561f
C812 B.n772 VSUBS 0.020561f
C813 B.n773 VSUBS 0.019074f
C814 B.n774 VSUBS 0.008694f
C815 B.n775 VSUBS 0.008694f
C816 B.n776 VSUBS 0.008694f
C817 B.n777 VSUBS 0.008694f
C818 B.n778 VSUBS 0.008694f
C819 B.n779 VSUBS 0.008694f
C820 B.n780 VSUBS 0.008694f
C821 B.n781 VSUBS 0.008694f
C822 B.n782 VSUBS 0.008694f
C823 B.n783 VSUBS 0.008694f
C824 B.n784 VSUBS 0.008694f
C825 B.n785 VSUBS 0.008694f
C826 B.n786 VSUBS 0.008694f
C827 B.n787 VSUBS 0.008694f
C828 B.n788 VSUBS 0.008694f
C829 B.n789 VSUBS 0.008694f
C830 B.n790 VSUBS 0.008694f
C831 B.n791 VSUBS 0.008694f
C832 B.n792 VSUBS 0.008694f
C833 B.n793 VSUBS 0.008694f
C834 B.n794 VSUBS 0.008694f
C835 B.n795 VSUBS 0.008694f
C836 B.n796 VSUBS 0.008694f
C837 B.n797 VSUBS 0.008694f
C838 B.n798 VSUBS 0.008694f
C839 B.n799 VSUBS 0.008694f
C840 B.n800 VSUBS 0.008694f
C841 B.n801 VSUBS 0.008694f
C842 B.n802 VSUBS 0.008694f
C843 B.n803 VSUBS 0.008694f
C844 B.n804 VSUBS 0.008694f
C845 B.n805 VSUBS 0.008694f
C846 B.n806 VSUBS 0.008694f
C847 B.n807 VSUBS 0.008694f
C848 B.n808 VSUBS 0.008694f
C849 B.n809 VSUBS 0.008694f
C850 B.n810 VSUBS 0.008694f
C851 B.n811 VSUBS 0.008694f
C852 B.n812 VSUBS 0.008694f
C853 B.n813 VSUBS 0.008694f
C854 B.n814 VSUBS 0.008694f
C855 B.n815 VSUBS 0.008694f
C856 B.n816 VSUBS 0.008694f
C857 B.n817 VSUBS 0.008694f
C858 B.n818 VSUBS 0.008694f
C859 B.n819 VSUBS 0.008694f
C860 B.n820 VSUBS 0.008694f
C861 B.n821 VSUBS 0.008694f
C862 B.n822 VSUBS 0.008694f
C863 B.n823 VSUBS 0.008694f
C864 B.n824 VSUBS 0.008694f
C865 B.n825 VSUBS 0.008694f
C866 B.n826 VSUBS 0.008694f
C867 B.n827 VSUBS 0.008694f
C868 B.n828 VSUBS 0.008694f
C869 B.n829 VSUBS 0.008694f
C870 B.n830 VSUBS 0.008694f
C871 B.n831 VSUBS 0.008694f
C872 B.n832 VSUBS 0.008694f
C873 B.n833 VSUBS 0.008694f
C874 B.n834 VSUBS 0.008694f
C875 B.n835 VSUBS 0.008694f
C876 B.n836 VSUBS 0.008694f
C877 B.n837 VSUBS 0.008694f
C878 B.n838 VSUBS 0.008694f
C879 B.n839 VSUBS 0.008694f
C880 B.n840 VSUBS 0.008694f
C881 B.n841 VSUBS 0.008694f
C882 B.n842 VSUBS 0.008694f
C883 B.n843 VSUBS 0.008694f
C884 B.n844 VSUBS 0.008694f
C885 B.n845 VSUBS 0.008694f
C886 B.n846 VSUBS 0.008694f
C887 B.n847 VSUBS 0.008694f
C888 B.n848 VSUBS 0.008694f
C889 B.n849 VSUBS 0.008694f
C890 B.n850 VSUBS 0.008694f
C891 B.n851 VSUBS 0.008694f
C892 B.n852 VSUBS 0.008694f
C893 B.n853 VSUBS 0.008694f
C894 B.n854 VSUBS 0.008694f
C895 B.n855 VSUBS 0.008694f
C896 B.n856 VSUBS 0.008694f
C897 B.n857 VSUBS 0.008694f
C898 B.n858 VSUBS 0.008694f
C899 B.n859 VSUBS 0.008694f
C900 B.n860 VSUBS 0.008694f
C901 B.n861 VSUBS 0.008694f
C902 B.n862 VSUBS 0.008694f
C903 B.n863 VSUBS 0.008694f
C904 B.n864 VSUBS 0.008694f
C905 B.n865 VSUBS 0.008694f
C906 B.n866 VSUBS 0.008694f
C907 B.n867 VSUBS 0.008694f
C908 B.n868 VSUBS 0.008694f
C909 B.n869 VSUBS 0.008694f
C910 B.n870 VSUBS 0.008694f
C911 B.n871 VSUBS 0.008694f
C912 B.n872 VSUBS 0.008694f
C913 B.n873 VSUBS 0.008694f
C914 B.n874 VSUBS 0.008694f
C915 B.n875 VSUBS 0.011346f
C916 B.n876 VSUBS 0.012086f
C917 B.n877 VSUBS 0.024034f
C918 VDD1.t1 VSUBS 0.234237f
C919 VDD1.t2 VSUBS 0.234237f
C920 VDD1.n0 VSUBS 1.7687f
C921 VDD1.t3 VSUBS 0.234237f
C922 VDD1.t5 VSUBS 0.234237f
C923 VDD1.n1 VSUBS 1.76687f
C924 VDD1.t4 VSUBS 0.234237f
C925 VDD1.t0 VSUBS 0.234237f
C926 VDD1.n2 VSUBS 1.76687f
C927 VDD1.n3 VSUBS 5.57625f
C928 VDD1.t6 VSUBS 0.234237f
C929 VDD1.t7 VSUBS 0.234237f
C930 VDD1.n4 VSUBS 1.74228f
C931 VDD1.n5 VSUBS 4.41438f
C932 VP.t7 VSUBS 2.78793f
C933 VP.n0 VSUBS 1.09795f
C934 VP.n1 VSUBS 0.028979f
C935 VP.n2 VSUBS 0.058534f
C936 VP.n3 VSUBS 0.028979f
C937 VP.n4 VSUBS 0.054009f
C938 VP.n5 VSUBS 0.028979f
C939 VP.t3 VSUBS 2.78793f
C940 VP.n6 VSUBS 0.054009f
C941 VP.n7 VSUBS 0.028979f
C942 VP.n8 VSUBS 0.054009f
C943 VP.n9 VSUBS 0.028979f
C944 VP.t2 VSUBS 2.78793f
C945 VP.n10 VSUBS 0.054009f
C946 VP.n11 VSUBS 0.028979f
C947 VP.n12 VSUBS 0.054009f
C948 VP.n13 VSUBS 0.046771f
C949 VP.t4 VSUBS 2.78793f
C950 VP.t0 VSUBS 2.78793f
C951 VP.n14 VSUBS 1.09795f
C952 VP.n15 VSUBS 0.028979f
C953 VP.n16 VSUBS 0.058534f
C954 VP.n17 VSUBS 0.028979f
C955 VP.n18 VSUBS 0.054009f
C956 VP.n19 VSUBS 0.028979f
C957 VP.t1 VSUBS 2.78793f
C958 VP.n20 VSUBS 0.054009f
C959 VP.n21 VSUBS 0.028979f
C960 VP.n22 VSUBS 0.054009f
C961 VP.t6 VSUBS 3.22606f
C962 VP.n23 VSUBS 1.05196f
C963 VP.t5 VSUBS 2.78793f
C964 VP.n24 VSUBS 1.10026f
C965 VP.n25 VSUBS 0.045476f
C966 VP.n26 VSUBS 0.375485f
C967 VP.n27 VSUBS 0.028979f
C968 VP.n28 VSUBS 0.028979f
C969 VP.n29 VSUBS 0.054009f
C970 VP.n30 VSUBS 0.042304f
C971 VP.n31 VSUBS 0.042304f
C972 VP.n32 VSUBS 0.028979f
C973 VP.n33 VSUBS 0.028979f
C974 VP.n34 VSUBS 0.028979f
C975 VP.n35 VSUBS 0.054009f
C976 VP.n36 VSUBS 0.045476f
C977 VP.n37 VSUBS 0.990717f
C978 VP.n38 VSUBS 0.035877f
C979 VP.n39 VSUBS 0.028979f
C980 VP.n40 VSUBS 0.028979f
C981 VP.n41 VSUBS 0.028979f
C982 VP.n42 VSUBS 0.054009f
C983 VP.n43 VSUBS 0.054779f
C984 VP.n44 VSUBS 0.025303f
C985 VP.n45 VSUBS 0.028979f
C986 VP.n46 VSUBS 0.028979f
C987 VP.n47 VSUBS 0.028979f
C988 VP.n48 VSUBS 0.054009f
C989 VP.n49 VSUBS 0.054009f
C990 VP.n50 VSUBS 0.028411f
C991 VP.n51 VSUBS 0.046771f
C992 VP.n52 VSUBS 1.89227f
C993 VP.n53 VSUBS 1.91131f
C994 VP.n54 VSUBS 1.09795f
C995 VP.n55 VSUBS 0.028411f
C996 VP.n56 VSUBS 0.054009f
C997 VP.n57 VSUBS 0.028979f
C998 VP.n58 VSUBS 0.028979f
C999 VP.n59 VSUBS 0.028979f
C1000 VP.n60 VSUBS 0.058534f
C1001 VP.n61 VSUBS 0.025303f
C1002 VP.n62 VSUBS 0.054779f
C1003 VP.n63 VSUBS 0.028979f
C1004 VP.n64 VSUBS 0.028979f
C1005 VP.n65 VSUBS 0.028979f
C1006 VP.n66 VSUBS 0.054009f
C1007 VP.n67 VSUBS 0.035877f
C1008 VP.n68 VSUBS 0.990717f
C1009 VP.n69 VSUBS 0.045476f
C1010 VP.n70 VSUBS 0.028979f
C1011 VP.n71 VSUBS 0.028979f
C1012 VP.n72 VSUBS 0.028979f
C1013 VP.n73 VSUBS 0.054009f
C1014 VP.n74 VSUBS 0.042304f
C1015 VP.n75 VSUBS 0.042304f
C1016 VP.n76 VSUBS 0.028979f
C1017 VP.n77 VSUBS 0.028979f
C1018 VP.n78 VSUBS 0.028979f
C1019 VP.n79 VSUBS 0.054009f
C1020 VP.n80 VSUBS 0.045476f
C1021 VP.n81 VSUBS 0.990717f
C1022 VP.n82 VSUBS 0.035877f
C1023 VP.n83 VSUBS 0.028979f
C1024 VP.n84 VSUBS 0.028979f
C1025 VP.n85 VSUBS 0.028979f
C1026 VP.n86 VSUBS 0.054009f
C1027 VP.n87 VSUBS 0.054779f
C1028 VP.n88 VSUBS 0.025303f
C1029 VP.n89 VSUBS 0.028979f
C1030 VP.n90 VSUBS 0.028979f
C1031 VP.n91 VSUBS 0.028979f
C1032 VP.n92 VSUBS 0.054009f
C1033 VP.n93 VSUBS 0.054009f
C1034 VP.n94 VSUBS 0.028411f
C1035 VP.n95 VSUBS 0.046771f
C1036 VP.n96 VSUBS 0.091432f
C1037 VTAIL.t4 VSUBS 0.201962f
C1038 VTAIL.t9 VSUBS 0.201962f
C1039 VTAIL.n0 VSUBS 1.37206f
C1040 VTAIL.n1 VSUBS 0.908375f
C1041 VTAIL.n2 VSUBS 0.028487f
C1042 VTAIL.n3 VSUBS 0.02763f
C1043 VTAIL.n4 VSUBS 0.014847f
C1044 VTAIL.n5 VSUBS 0.035093f
C1045 VTAIL.n6 VSUBS 0.015284f
C1046 VTAIL.n7 VSUBS 0.02763f
C1047 VTAIL.n8 VSUBS 0.01572f
C1048 VTAIL.n9 VSUBS 0.035093f
C1049 VTAIL.n10 VSUBS 0.01572f
C1050 VTAIL.n11 VSUBS 0.02763f
C1051 VTAIL.n12 VSUBS 0.014847f
C1052 VTAIL.n13 VSUBS 0.035093f
C1053 VTAIL.n14 VSUBS 0.01572f
C1054 VTAIL.n15 VSUBS 1.02455f
C1055 VTAIL.n16 VSUBS 0.014847f
C1056 VTAIL.t11 VSUBS 0.075397f
C1057 VTAIL.n17 VSUBS 0.183272f
C1058 VTAIL.n18 VSUBS 0.026399f
C1059 VTAIL.n19 VSUBS 0.02632f
C1060 VTAIL.n20 VSUBS 0.035093f
C1061 VTAIL.n21 VSUBS 0.01572f
C1062 VTAIL.n22 VSUBS 0.014847f
C1063 VTAIL.n23 VSUBS 0.02763f
C1064 VTAIL.n24 VSUBS 0.02763f
C1065 VTAIL.n25 VSUBS 0.014847f
C1066 VTAIL.n26 VSUBS 0.01572f
C1067 VTAIL.n27 VSUBS 0.035093f
C1068 VTAIL.n28 VSUBS 0.035093f
C1069 VTAIL.n29 VSUBS 0.01572f
C1070 VTAIL.n30 VSUBS 0.014847f
C1071 VTAIL.n31 VSUBS 0.02763f
C1072 VTAIL.n32 VSUBS 0.02763f
C1073 VTAIL.n33 VSUBS 0.014847f
C1074 VTAIL.n34 VSUBS 0.014847f
C1075 VTAIL.n35 VSUBS 0.01572f
C1076 VTAIL.n36 VSUBS 0.035093f
C1077 VTAIL.n37 VSUBS 0.035093f
C1078 VTAIL.n38 VSUBS 0.035093f
C1079 VTAIL.n39 VSUBS 0.015284f
C1080 VTAIL.n40 VSUBS 0.014847f
C1081 VTAIL.n41 VSUBS 0.02763f
C1082 VTAIL.n42 VSUBS 0.02763f
C1083 VTAIL.n43 VSUBS 0.014847f
C1084 VTAIL.n44 VSUBS 0.01572f
C1085 VTAIL.n45 VSUBS 0.035093f
C1086 VTAIL.n46 VSUBS 0.078578f
C1087 VTAIL.n47 VSUBS 0.01572f
C1088 VTAIL.n48 VSUBS 0.014847f
C1089 VTAIL.n49 VSUBS 0.064242f
C1090 VTAIL.n50 VSUBS 0.039245f
C1091 VTAIL.n51 VSUBS 0.386449f
C1092 VTAIL.n52 VSUBS 0.028487f
C1093 VTAIL.n53 VSUBS 0.02763f
C1094 VTAIL.n54 VSUBS 0.014847f
C1095 VTAIL.n55 VSUBS 0.035093f
C1096 VTAIL.n56 VSUBS 0.015284f
C1097 VTAIL.n57 VSUBS 0.02763f
C1098 VTAIL.n58 VSUBS 0.01572f
C1099 VTAIL.n59 VSUBS 0.035093f
C1100 VTAIL.n60 VSUBS 0.01572f
C1101 VTAIL.n61 VSUBS 0.02763f
C1102 VTAIL.n62 VSUBS 0.014847f
C1103 VTAIL.n63 VSUBS 0.035093f
C1104 VTAIL.n64 VSUBS 0.01572f
C1105 VTAIL.n65 VSUBS 1.02455f
C1106 VTAIL.n66 VSUBS 0.014847f
C1107 VTAIL.t0 VSUBS 0.075397f
C1108 VTAIL.n67 VSUBS 0.183272f
C1109 VTAIL.n68 VSUBS 0.026399f
C1110 VTAIL.n69 VSUBS 0.02632f
C1111 VTAIL.n70 VSUBS 0.035093f
C1112 VTAIL.n71 VSUBS 0.01572f
C1113 VTAIL.n72 VSUBS 0.014847f
C1114 VTAIL.n73 VSUBS 0.02763f
C1115 VTAIL.n74 VSUBS 0.02763f
C1116 VTAIL.n75 VSUBS 0.014847f
C1117 VTAIL.n76 VSUBS 0.01572f
C1118 VTAIL.n77 VSUBS 0.035093f
C1119 VTAIL.n78 VSUBS 0.035093f
C1120 VTAIL.n79 VSUBS 0.01572f
C1121 VTAIL.n80 VSUBS 0.014847f
C1122 VTAIL.n81 VSUBS 0.02763f
C1123 VTAIL.n82 VSUBS 0.02763f
C1124 VTAIL.n83 VSUBS 0.014847f
C1125 VTAIL.n84 VSUBS 0.014847f
C1126 VTAIL.n85 VSUBS 0.01572f
C1127 VTAIL.n86 VSUBS 0.035093f
C1128 VTAIL.n87 VSUBS 0.035093f
C1129 VTAIL.n88 VSUBS 0.035093f
C1130 VTAIL.n89 VSUBS 0.015284f
C1131 VTAIL.n90 VSUBS 0.014847f
C1132 VTAIL.n91 VSUBS 0.02763f
C1133 VTAIL.n92 VSUBS 0.02763f
C1134 VTAIL.n93 VSUBS 0.014847f
C1135 VTAIL.n94 VSUBS 0.01572f
C1136 VTAIL.n95 VSUBS 0.035093f
C1137 VTAIL.n96 VSUBS 0.078578f
C1138 VTAIL.n97 VSUBS 0.01572f
C1139 VTAIL.n98 VSUBS 0.014847f
C1140 VTAIL.n99 VSUBS 0.064242f
C1141 VTAIL.n100 VSUBS 0.039245f
C1142 VTAIL.n101 VSUBS 0.386449f
C1143 VTAIL.t15 VSUBS 0.201962f
C1144 VTAIL.t12 VSUBS 0.201962f
C1145 VTAIL.n102 VSUBS 1.37206f
C1146 VTAIL.n103 VSUBS 1.22401f
C1147 VTAIL.n104 VSUBS 0.028487f
C1148 VTAIL.n105 VSUBS 0.02763f
C1149 VTAIL.n106 VSUBS 0.014847f
C1150 VTAIL.n107 VSUBS 0.035093f
C1151 VTAIL.n108 VSUBS 0.015284f
C1152 VTAIL.n109 VSUBS 0.02763f
C1153 VTAIL.n110 VSUBS 0.01572f
C1154 VTAIL.n111 VSUBS 0.035093f
C1155 VTAIL.n112 VSUBS 0.01572f
C1156 VTAIL.n113 VSUBS 0.02763f
C1157 VTAIL.n114 VSUBS 0.014847f
C1158 VTAIL.n115 VSUBS 0.035093f
C1159 VTAIL.n116 VSUBS 0.01572f
C1160 VTAIL.n117 VSUBS 1.02455f
C1161 VTAIL.n118 VSUBS 0.014847f
C1162 VTAIL.t3 VSUBS 0.075397f
C1163 VTAIL.n119 VSUBS 0.183272f
C1164 VTAIL.n120 VSUBS 0.026399f
C1165 VTAIL.n121 VSUBS 0.02632f
C1166 VTAIL.n122 VSUBS 0.035093f
C1167 VTAIL.n123 VSUBS 0.01572f
C1168 VTAIL.n124 VSUBS 0.014847f
C1169 VTAIL.n125 VSUBS 0.02763f
C1170 VTAIL.n126 VSUBS 0.02763f
C1171 VTAIL.n127 VSUBS 0.014847f
C1172 VTAIL.n128 VSUBS 0.01572f
C1173 VTAIL.n129 VSUBS 0.035093f
C1174 VTAIL.n130 VSUBS 0.035093f
C1175 VTAIL.n131 VSUBS 0.01572f
C1176 VTAIL.n132 VSUBS 0.014847f
C1177 VTAIL.n133 VSUBS 0.02763f
C1178 VTAIL.n134 VSUBS 0.02763f
C1179 VTAIL.n135 VSUBS 0.014847f
C1180 VTAIL.n136 VSUBS 0.014847f
C1181 VTAIL.n137 VSUBS 0.01572f
C1182 VTAIL.n138 VSUBS 0.035093f
C1183 VTAIL.n139 VSUBS 0.035093f
C1184 VTAIL.n140 VSUBS 0.035093f
C1185 VTAIL.n141 VSUBS 0.015284f
C1186 VTAIL.n142 VSUBS 0.014847f
C1187 VTAIL.n143 VSUBS 0.02763f
C1188 VTAIL.n144 VSUBS 0.02763f
C1189 VTAIL.n145 VSUBS 0.014847f
C1190 VTAIL.n146 VSUBS 0.01572f
C1191 VTAIL.n147 VSUBS 0.035093f
C1192 VTAIL.n148 VSUBS 0.078578f
C1193 VTAIL.n149 VSUBS 0.01572f
C1194 VTAIL.n150 VSUBS 0.014847f
C1195 VTAIL.n151 VSUBS 0.064242f
C1196 VTAIL.n152 VSUBS 0.039245f
C1197 VTAIL.n153 VSUBS 1.75067f
C1198 VTAIL.n154 VSUBS 0.028487f
C1199 VTAIL.n155 VSUBS 0.02763f
C1200 VTAIL.n156 VSUBS 0.014847f
C1201 VTAIL.n157 VSUBS 0.035093f
C1202 VTAIL.n158 VSUBS 0.015284f
C1203 VTAIL.n159 VSUBS 0.02763f
C1204 VTAIL.n160 VSUBS 0.015284f
C1205 VTAIL.n161 VSUBS 0.014847f
C1206 VTAIL.n162 VSUBS 0.035093f
C1207 VTAIL.n163 VSUBS 0.035093f
C1208 VTAIL.n164 VSUBS 0.01572f
C1209 VTAIL.n165 VSUBS 0.02763f
C1210 VTAIL.n166 VSUBS 0.014847f
C1211 VTAIL.n167 VSUBS 0.035093f
C1212 VTAIL.n168 VSUBS 0.01572f
C1213 VTAIL.n169 VSUBS 1.02455f
C1214 VTAIL.n170 VSUBS 0.014847f
C1215 VTAIL.t8 VSUBS 0.075397f
C1216 VTAIL.n171 VSUBS 0.183272f
C1217 VTAIL.n172 VSUBS 0.026399f
C1218 VTAIL.n173 VSUBS 0.02632f
C1219 VTAIL.n174 VSUBS 0.035093f
C1220 VTAIL.n175 VSUBS 0.01572f
C1221 VTAIL.n176 VSUBS 0.014847f
C1222 VTAIL.n177 VSUBS 0.02763f
C1223 VTAIL.n178 VSUBS 0.02763f
C1224 VTAIL.n179 VSUBS 0.014847f
C1225 VTAIL.n180 VSUBS 0.01572f
C1226 VTAIL.n181 VSUBS 0.035093f
C1227 VTAIL.n182 VSUBS 0.035093f
C1228 VTAIL.n183 VSUBS 0.01572f
C1229 VTAIL.n184 VSUBS 0.014847f
C1230 VTAIL.n185 VSUBS 0.02763f
C1231 VTAIL.n186 VSUBS 0.02763f
C1232 VTAIL.n187 VSUBS 0.014847f
C1233 VTAIL.n188 VSUBS 0.01572f
C1234 VTAIL.n189 VSUBS 0.035093f
C1235 VTAIL.n190 VSUBS 0.035093f
C1236 VTAIL.n191 VSUBS 0.01572f
C1237 VTAIL.n192 VSUBS 0.014847f
C1238 VTAIL.n193 VSUBS 0.02763f
C1239 VTAIL.n194 VSUBS 0.02763f
C1240 VTAIL.n195 VSUBS 0.014847f
C1241 VTAIL.n196 VSUBS 0.01572f
C1242 VTAIL.n197 VSUBS 0.035093f
C1243 VTAIL.n198 VSUBS 0.078578f
C1244 VTAIL.n199 VSUBS 0.01572f
C1245 VTAIL.n200 VSUBS 0.014847f
C1246 VTAIL.n201 VSUBS 0.064242f
C1247 VTAIL.n202 VSUBS 0.039245f
C1248 VTAIL.n203 VSUBS 1.75067f
C1249 VTAIL.t5 VSUBS 0.201962f
C1250 VTAIL.t7 VSUBS 0.201962f
C1251 VTAIL.n204 VSUBS 1.37207f
C1252 VTAIL.n205 VSUBS 1.224f
C1253 VTAIL.n206 VSUBS 0.028487f
C1254 VTAIL.n207 VSUBS 0.02763f
C1255 VTAIL.n208 VSUBS 0.014847f
C1256 VTAIL.n209 VSUBS 0.035093f
C1257 VTAIL.n210 VSUBS 0.015284f
C1258 VTAIL.n211 VSUBS 0.02763f
C1259 VTAIL.n212 VSUBS 0.015284f
C1260 VTAIL.n213 VSUBS 0.014847f
C1261 VTAIL.n214 VSUBS 0.035093f
C1262 VTAIL.n215 VSUBS 0.035093f
C1263 VTAIL.n216 VSUBS 0.01572f
C1264 VTAIL.n217 VSUBS 0.02763f
C1265 VTAIL.n218 VSUBS 0.014847f
C1266 VTAIL.n219 VSUBS 0.035093f
C1267 VTAIL.n220 VSUBS 0.01572f
C1268 VTAIL.n221 VSUBS 1.02455f
C1269 VTAIL.n222 VSUBS 0.014847f
C1270 VTAIL.t6 VSUBS 0.075397f
C1271 VTAIL.n223 VSUBS 0.183272f
C1272 VTAIL.n224 VSUBS 0.026399f
C1273 VTAIL.n225 VSUBS 0.02632f
C1274 VTAIL.n226 VSUBS 0.035093f
C1275 VTAIL.n227 VSUBS 0.01572f
C1276 VTAIL.n228 VSUBS 0.014847f
C1277 VTAIL.n229 VSUBS 0.02763f
C1278 VTAIL.n230 VSUBS 0.02763f
C1279 VTAIL.n231 VSUBS 0.014847f
C1280 VTAIL.n232 VSUBS 0.01572f
C1281 VTAIL.n233 VSUBS 0.035093f
C1282 VTAIL.n234 VSUBS 0.035093f
C1283 VTAIL.n235 VSUBS 0.01572f
C1284 VTAIL.n236 VSUBS 0.014847f
C1285 VTAIL.n237 VSUBS 0.02763f
C1286 VTAIL.n238 VSUBS 0.02763f
C1287 VTAIL.n239 VSUBS 0.014847f
C1288 VTAIL.n240 VSUBS 0.01572f
C1289 VTAIL.n241 VSUBS 0.035093f
C1290 VTAIL.n242 VSUBS 0.035093f
C1291 VTAIL.n243 VSUBS 0.01572f
C1292 VTAIL.n244 VSUBS 0.014847f
C1293 VTAIL.n245 VSUBS 0.02763f
C1294 VTAIL.n246 VSUBS 0.02763f
C1295 VTAIL.n247 VSUBS 0.014847f
C1296 VTAIL.n248 VSUBS 0.01572f
C1297 VTAIL.n249 VSUBS 0.035093f
C1298 VTAIL.n250 VSUBS 0.078578f
C1299 VTAIL.n251 VSUBS 0.01572f
C1300 VTAIL.n252 VSUBS 0.014847f
C1301 VTAIL.n253 VSUBS 0.064242f
C1302 VTAIL.n254 VSUBS 0.039245f
C1303 VTAIL.n255 VSUBS 0.386449f
C1304 VTAIL.n256 VSUBS 0.028487f
C1305 VTAIL.n257 VSUBS 0.02763f
C1306 VTAIL.n258 VSUBS 0.014847f
C1307 VTAIL.n259 VSUBS 0.035093f
C1308 VTAIL.n260 VSUBS 0.015284f
C1309 VTAIL.n261 VSUBS 0.02763f
C1310 VTAIL.n262 VSUBS 0.015284f
C1311 VTAIL.n263 VSUBS 0.014847f
C1312 VTAIL.n264 VSUBS 0.035093f
C1313 VTAIL.n265 VSUBS 0.035093f
C1314 VTAIL.n266 VSUBS 0.01572f
C1315 VTAIL.n267 VSUBS 0.02763f
C1316 VTAIL.n268 VSUBS 0.014847f
C1317 VTAIL.n269 VSUBS 0.035093f
C1318 VTAIL.n270 VSUBS 0.01572f
C1319 VTAIL.n271 VSUBS 1.02455f
C1320 VTAIL.n272 VSUBS 0.014847f
C1321 VTAIL.t1 VSUBS 0.075397f
C1322 VTAIL.n273 VSUBS 0.183272f
C1323 VTAIL.n274 VSUBS 0.026399f
C1324 VTAIL.n275 VSUBS 0.02632f
C1325 VTAIL.n276 VSUBS 0.035093f
C1326 VTAIL.n277 VSUBS 0.01572f
C1327 VTAIL.n278 VSUBS 0.014847f
C1328 VTAIL.n279 VSUBS 0.02763f
C1329 VTAIL.n280 VSUBS 0.02763f
C1330 VTAIL.n281 VSUBS 0.014847f
C1331 VTAIL.n282 VSUBS 0.01572f
C1332 VTAIL.n283 VSUBS 0.035093f
C1333 VTAIL.n284 VSUBS 0.035093f
C1334 VTAIL.n285 VSUBS 0.01572f
C1335 VTAIL.n286 VSUBS 0.014847f
C1336 VTAIL.n287 VSUBS 0.02763f
C1337 VTAIL.n288 VSUBS 0.02763f
C1338 VTAIL.n289 VSUBS 0.014847f
C1339 VTAIL.n290 VSUBS 0.01572f
C1340 VTAIL.n291 VSUBS 0.035093f
C1341 VTAIL.n292 VSUBS 0.035093f
C1342 VTAIL.n293 VSUBS 0.01572f
C1343 VTAIL.n294 VSUBS 0.014847f
C1344 VTAIL.n295 VSUBS 0.02763f
C1345 VTAIL.n296 VSUBS 0.02763f
C1346 VTAIL.n297 VSUBS 0.014847f
C1347 VTAIL.n298 VSUBS 0.01572f
C1348 VTAIL.n299 VSUBS 0.035093f
C1349 VTAIL.n300 VSUBS 0.078578f
C1350 VTAIL.n301 VSUBS 0.01572f
C1351 VTAIL.n302 VSUBS 0.014847f
C1352 VTAIL.n303 VSUBS 0.064242f
C1353 VTAIL.n304 VSUBS 0.039245f
C1354 VTAIL.n305 VSUBS 0.386449f
C1355 VTAIL.t2 VSUBS 0.201962f
C1356 VTAIL.t14 VSUBS 0.201962f
C1357 VTAIL.n306 VSUBS 1.37207f
C1358 VTAIL.n307 VSUBS 1.224f
C1359 VTAIL.n308 VSUBS 0.028487f
C1360 VTAIL.n309 VSUBS 0.02763f
C1361 VTAIL.n310 VSUBS 0.014847f
C1362 VTAIL.n311 VSUBS 0.035093f
C1363 VTAIL.n312 VSUBS 0.015284f
C1364 VTAIL.n313 VSUBS 0.02763f
C1365 VTAIL.n314 VSUBS 0.015284f
C1366 VTAIL.n315 VSUBS 0.014847f
C1367 VTAIL.n316 VSUBS 0.035093f
C1368 VTAIL.n317 VSUBS 0.035093f
C1369 VTAIL.n318 VSUBS 0.01572f
C1370 VTAIL.n319 VSUBS 0.02763f
C1371 VTAIL.n320 VSUBS 0.014847f
C1372 VTAIL.n321 VSUBS 0.035093f
C1373 VTAIL.n322 VSUBS 0.01572f
C1374 VTAIL.n323 VSUBS 1.02455f
C1375 VTAIL.n324 VSUBS 0.014847f
C1376 VTAIL.t13 VSUBS 0.075397f
C1377 VTAIL.n325 VSUBS 0.183272f
C1378 VTAIL.n326 VSUBS 0.026399f
C1379 VTAIL.n327 VSUBS 0.02632f
C1380 VTAIL.n328 VSUBS 0.035093f
C1381 VTAIL.n329 VSUBS 0.01572f
C1382 VTAIL.n330 VSUBS 0.014847f
C1383 VTAIL.n331 VSUBS 0.02763f
C1384 VTAIL.n332 VSUBS 0.02763f
C1385 VTAIL.n333 VSUBS 0.014847f
C1386 VTAIL.n334 VSUBS 0.01572f
C1387 VTAIL.n335 VSUBS 0.035093f
C1388 VTAIL.n336 VSUBS 0.035093f
C1389 VTAIL.n337 VSUBS 0.01572f
C1390 VTAIL.n338 VSUBS 0.014847f
C1391 VTAIL.n339 VSUBS 0.02763f
C1392 VTAIL.n340 VSUBS 0.02763f
C1393 VTAIL.n341 VSUBS 0.014847f
C1394 VTAIL.n342 VSUBS 0.01572f
C1395 VTAIL.n343 VSUBS 0.035093f
C1396 VTAIL.n344 VSUBS 0.035093f
C1397 VTAIL.n345 VSUBS 0.01572f
C1398 VTAIL.n346 VSUBS 0.014847f
C1399 VTAIL.n347 VSUBS 0.02763f
C1400 VTAIL.n348 VSUBS 0.02763f
C1401 VTAIL.n349 VSUBS 0.014847f
C1402 VTAIL.n350 VSUBS 0.01572f
C1403 VTAIL.n351 VSUBS 0.035093f
C1404 VTAIL.n352 VSUBS 0.078578f
C1405 VTAIL.n353 VSUBS 0.01572f
C1406 VTAIL.n354 VSUBS 0.014847f
C1407 VTAIL.n355 VSUBS 0.064242f
C1408 VTAIL.n356 VSUBS 0.039245f
C1409 VTAIL.n357 VSUBS 1.75067f
C1410 VTAIL.n358 VSUBS 0.028487f
C1411 VTAIL.n359 VSUBS 0.02763f
C1412 VTAIL.n360 VSUBS 0.014847f
C1413 VTAIL.n361 VSUBS 0.035093f
C1414 VTAIL.n362 VSUBS 0.015284f
C1415 VTAIL.n363 VSUBS 0.02763f
C1416 VTAIL.n364 VSUBS 0.01572f
C1417 VTAIL.n365 VSUBS 0.035093f
C1418 VTAIL.n366 VSUBS 0.01572f
C1419 VTAIL.n367 VSUBS 0.02763f
C1420 VTAIL.n368 VSUBS 0.014847f
C1421 VTAIL.n369 VSUBS 0.035093f
C1422 VTAIL.n370 VSUBS 0.01572f
C1423 VTAIL.n371 VSUBS 1.02455f
C1424 VTAIL.n372 VSUBS 0.014847f
C1425 VTAIL.t10 VSUBS 0.075397f
C1426 VTAIL.n373 VSUBS 0.183272f
C1427 VTAIL.n374 VSUBS 0.026399f
C1428 VTAIL.n375 VSUBS 0.02632f
C1429 VTAIL.n376 VSUBS 0.035093f
C1430 VTAIL.n377 VSUBS 0.01572f
C1431 VTAIL.n378 VSUBS 0.014847f
C1432 VTAIL.n379 VSUBS 0.02763f
C1433 VTAIL.n380 VSUBS 0.02763f
C1434 VTAIL.n381 VSUBS 0.014847f
C1435 VTAIL.n382 VSUBS 0.01572f
C1436 VTAIL.n383 VSUBS 0.035093f
C1437 VTAIL.n384 VSUBS 0.035093f
C1438 VTAIL.n385 VSUBS 0.01572f
C1439 VTAIL.n386 VSUBS 0.014847f
C1440 VTAIL.n387 VSUBS 0.02763f
C1441 VTAIL.n388 VSUBS 0.02763f
C1442 VTAIL.n389 VSUBS 0.014847f
C1443 VTAIL.n390 VSUBS 0.014847f
C1444 VTAIL.n391 VSUBS 0.01572f
C1445 VTAIL.n392 VSUBS 0.035093f
C1446 VTAIL.n393 VSUBS 0.035093f
C1447 VTAIL.n394 VSUBS 0.035093f
C1448 VTAIL.n395 VSUBS 0.015284f
C1449 VTAIL.n396 VSUBS 0.014847f
C1450 VTAIL.n397 VSUBS 0.02763f
C1451 VTAIL.n398 VSUBS 0.02763f
C1452 VTAIL.n399 VSUBS 0.014847f
C1453 VTAIL.n400 VSUBS 0.01572f
C1454 VTAIL.n401 VSUBS 0.035093f
C1455 VTAIL.n402 VSUBS 0.078578f
C1456 VTAIL.n403 VSUBS 0.01572f
C1457 VTAIL.n404 VSUBS 0.014847f
C1458 VTAIL.n405 VSUBS 0.064242f
C1459 VTAIL.n406 VSUBS 0.039245f
C1460 VTAIL.n407 VSUBS 1.74549f
C1461 VDD2.t6 VSUBS 0.255238f
C1462 VDD2.t4 VSUBS 0.255238f
C1463 VDD2.n0 VSUBS 1.92528f
C1464 VDD2.t5 VSUBS 0.255238f
C1465 VDD2.t7 VSUBS 0.255238f
C1466 VDD2.n1 VSUBS 1.92528f
C1467 VDD2.n2 VSUBS 6.00424f
C1468 VDD2.t0 VSUBS 0.255238f
C1469 VDD2.t3 VSUBS 0.255238f
C1470 VDD2.n3 VSUBS 1.89849f
C1471 VDD2.n4 VSUBS 4.76622f
C1472 VDD2.t1 VSUBS 0.255238f
C1473 VDD2.t2 VSUBS 0.255238f
C1474 VDD2.n5 VSUBS 1.92522f
C1475 VN.t1 VSUBS 2.51225f
C1476 VN.n0 VSUBS 0.989378f
C1477 VN.n1 VSUBS 0.026113f
C1478 VN.n2 VSUBS 0.052746f
C1479 VN.n3 VSUBS 0.026113f
C1480 VN.n4 VSUBS 0.048668f
C1481 VN.n5 VSUBS 0.026113f
C1482 VN.t2 VSUBS 2.51225f
C1483 VN.n6 VSUBS 0.048668f
C1484 VN.n7 VSUBS 0.026113f
C1485 VN.n8 VSUBS 0.048668f
C1486 VN.t0 VSUBS 2.90705f
C1487 VN.n9 VSUBS 0.947938f
C1488 VN.t7 VSUBS 2.51225f
C1489 VN.n10 VSUBS 0.991458f
C1490 VN.n11 VSUBS 0.040979f
C1491 VN.n12 VSUBS 0.338355f
C1492 VN.n13 VSUBS 0.026113f
C1493 VN.n14 VSUBS 0.026113f
C1494 VN.n15 VSUBS 0.048668f
C1495 VN.n16 VSUBS 0.038121f
C1496 VN.n17 VSUBS 0.038121f
C1497 VN.n18 VSUBS 0.026113f
C1498 VN.n19 VSUBS 0.026113f
C1499 VN.n20 VSUBS 0.026113f
C1500 VN.n21 VSUBS 0.048668f
C1501 VN.n22 VSUBS 0.040979f
C1502 VN.n23 VSUBS 0.89275f
C1503 VN.n24 VSUBS 0.032329f
C1504 VN.n25 VSUBS 0.026113f
C1505 VN.n26 VSUBS 0.026113f
C1506 VN.n27 VSUBS 0.026113f
C1507 VN.n28 VSUBS 0.048668f
C1508 VN.n29 VSUBS 0.049362f
C1509 VN.n30 VSUBS 0.022801f
C1510 VN.n31 VSUBS 0.026113f
C1511 VN.n32 VSUBS 0.026113f
C1512 VN.n33 VSUBS 0.026113f
C1513 VN.n34 VSUBS 0.048668f
C1514 VN.n35 VSUBS 0.048668f
C1515 VN.n36 VSUBS 0.025602f
C1516 VN.n37 VSUBS 0.042146f
C1517 VN.n38 VSUBS 0.082391f
C1518 VN.t3 VSUBS 2.51225f
C1519 VN.n39 VSUBS 0.989378f
C1520 VN.n40 VSUBS 0.026113f
C1521 VN.n41 VSUBS 0.052746f
C1522 VN.n42 VSUBS 0.026113f
C1523 VN.n43 VSUBS 0.048668f
C1524 VN.n44 VSUBS 0.026113f
C1525 VN.t6 VSUBS 2.51225f
C1526 VN.n45 VSUBS 0.048668f
C1527 VN.n46 VSUBS 0.026113f
C1528 VN.n47 VSUBS 0.048668f
C1529 VN.t5 VSUBS 2.90705f
C1530 VN.n48 VSUBS 0.947938f
C1531 VN.t4 VSUBS 2.51225f
C1532 VN.n49 VSUBS 0.991458f
C1533 VN.n50 VSUBS 0.040979f
C1534 VN.n51 VSUBS 0.338355f
C1535 VN.n52 VSUBS 0.026113f
C1536 VN.n53 VSUBS 0.026113f
C1537 VN.n54 VSUBS 0.048668f
C1538 VN.n55 VSUBS 0.038121f
C1539 VN.n56 VSUBS 0.038121f
C1540 VN.n57 VSUBS 0.026113f
C1541 VN.n58 VSUBS 0.026113f
C1542 VN.n59 VSUBS 0.026113f
C1543 VN.n60 VSUBS 0.048668f
C1544 VN.n61 VSUBS 0.040979f
C1545 VN.n62 VSUBS 0.89275f
C1546 VN.n63 VSUBS 0.032329f
C1547 VN.n64 VSUBS 0.026113f
C1548 VN.n65 VSUBS 0.026113f
C1549 VN.n66 VSUBS 0.026113f
C1550 VN.n67 VSUBS 0.048668f
C1551 VN.n68 VSUBS 0.049362f
C1552 VN.n69 VSUBS 0.022801f
C1553 VN.n70 VSUBS 0.026113f
C1554 VN.n71 VSUBS 0.026113f
C1555 VN.n72 VSUBS 0.026113f
C1556 VN.n73 VSUBS 0.048668f
C1557 VN.n74 VSUBS 0.048668f
C1558 VN.n75 VSUBS 0.025602f
C1559 VN.n76 VSUBS 0.042146f
C1560 VN.n77 VSUBS 1.71552f
.ends

