* NGSPICE file created from diff_pair_sample_1196.ext - technology: sky130A

.subckt diff_pair_sample_1196 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=1.02
X1 VTAIL.t16 VN.t1 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X2 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X3 VDD2.t7 VN.t2 VTAIL.t19 B.t1 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X4 VDD2.t6 VN.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X5 VTAIL.t7 VP.t1 VDD1.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X6 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=1.02
X7 VDD1.t7 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X8 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=1.02
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=1.02
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=1.02
X11 VTAIL.t15 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X12 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X13 VTAIL.t17 VN.t5 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X14 VDD2.t3 VN.t6 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=1.02
X15 VDD1.t5 VP.t4 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=1.02
X16 VDD2.t2 VN.t7 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=1.02
X17 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=1.02
X18 VTAIL.t0 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X19 VDD1.t2 VP.t7 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=1.02
X20 VTAIL.t4 VP.t8 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
X21 VDD2.t1 VN.t8 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=1.02
X22 VDD1.t0 VP.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=1.02
X23 VTAIL.t13 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=1.02
R0 VN.n37 VN.n20 161.3
R1 VN.n35 VN.n34 161.3
R2 VN.n33 VN.n21 161.3
R3 VN.n32 VN.n31 161.3
R4 VN.n29 VN.n22 161.3
R5 VN.n28 VN.n27 161.3
R6 VN.n26 VN.n23 161.3
R7 VN.n17 VN.n0 161.3
R8 VN.n15 VN.n14 161.3
R9 VN.n13 VN.n1 161.3
R10 VN.n12 VN.n11 161.3
R11 VN.n9 VN.n2 161.3
R12 VN.n8 VN.n7 161.3
R13 VN.n6 VN.n3 161.3
R14 VN.n5 VN.t6 133.029
R15 VN.n25 VN.t7 133.029
R16 VN.n18 VN.t0 118.374
R17 VN.n38 VN.t8 118.374
R18 VN.n39 VN.n38 80.6037
R19 VN.n19 VN.n18 80.6037
R20 VN.n4 VN.t1 79.625
R21 VN.n10 VN.t3 79.625
R22 VN.n16 VN.t5 79.625
R23 VN.n24 VN.t4 79.625
R24 VN.n30 VN.t2 79.625
R25 VN.n36 VN.t9 79.625
R26 VN.n18 VN.n17 53.5832
R27 VN.n38 VN.n37 53.5832
R28 VN.n5 VN.n4 48.7962
R29 VN.n25 VN.n24 48.7962
R30 VN.n9 VN.n8 47.7779
R31 VN.n11 VN.n1 47.7779
R32 VN.n29 VN.n28 47.7779
R33 VN.n31 VN.n21 47.7779
R34 VN.n26 VN.n25 44.3029
R35 VN.n6 VN.n5 44.3029
R36 VN VN.n39 38.4574
R37 VN.n8 VN.n3 33.2089
R38 VN.n15 VN.n1 33.2089
R39 VN.n28 VN.n23 33.2089
R40 VN.n35 VN.n21 33.2089
R41 VN.n17 VN.n16 19.5741
R42 VN.n37 VN.n36 19.5741
R43 VN.n10 VN.n9 12.234
R44 VN.n11 VN.n10 12.234
R45 VN.n31 VN.n30 12.234
R46 VN.n30 VN.n29 12.234
R47 VN.n4 VN.n3 4.8939
R48 VN.n16 VN.n15 4.8939
R49 VN.n24 VN.n23 4.8939
R50 VN.n36 VN.n35 4.8939
R51 VN.n39 VN.n20 0.285035
R52 VN.n19 VN.n0 0.285035
R53 VN.n34 VN.n20 0.189894
R54 VN.n34 VN.n33 0.189894
R55 VN.n33 VN.n32 0.189894
R56 VN.n32 VN.n22 0.189894
R57 VN.n27 VN.n22 0.189894
R58 VN.n27 VN.n26 0.189894
R59 VN.n7 VN.n6 0.189894
R60 VN.n7 VN.n2 0.189894
R61 VN.n12 VN.n2 0.189894
R62 VN.n13 VN.n12 0.189894
R63 VN.n14 VN.n13 0.189894
R64 VN.n14 VN.n0 0.189894
R65 VN VN.n19 0.146778
R66 VTAIL.n72 VTAIL.n62 289.615
R67 VTAIL.n12 VTAIL.n2 289.615
R68 VTAIL.n56 VTAIL.n46 289.615
R69 VTAIL.n36 VTAIL.n26 289.615
R70 VTAIL.n66 VTAIL.n65 185
R71 VTAIL.n71 VTAIL.n70 185
R72 VTAIL.n73 VTAIL.n72 185
R73 VTAIL.n6 VTAIL.n5 185
R74 VTAIL.n11 VTAIL.n10 185
R75 VTAIL.n13 VTAIL.n12 185
R76 VTAIL.n57 VTAIL.n56 185
R77 VTAIL.n55 VTAIL.n54 185
R78 VTAIL.n50 VTAIL.n49 185
R79 VTAIL.n37 VTAIL.n36 185
R80 VTAIL.n35 VTAIL.n34 185
R81 VTAIL.n30 VTAIL.n29 185
R82 VTAIL.n67 VTAIL.t18 150.499
R83 VTAIL.n7 VTAIL.t2 150.499
R84 VTAIL.n31 VTAIL.t12 150.499
R85 VTAIL.n51 VTAIL.t8 150.499
R86 VTAIL.n71 VTAIL.n65 104.615
R87 VTAIL.n72 VTAIL.n71 104.615
R88 VTAIL.n11 VTAIL.n5 104.615
R89 VTAIL.n12 VTAIL.n11 104.615
R90 VTAIL.n56 VTAIL.n55 104.615
R91 VTAIL.n55 VTAIL.n49 104.615
R92 VTAIL.n36 VTAIL.n35 104.615
R93 VTAIL.n35 VTAIL.n29 104.615
R94 VTAIL.n45 VTAIL.n44 60.0588
R95 VTAIL.n43 VTAIL.n42 60.0588
R96 VTAIL.n25 VTAIL.n24 60.0588
R97 VTAIL.n23 VTAIL.n22 60.0588
R98 VTAIL.n79 VTAIL.n78 60.0588
R99 VTAIL.n1 VTAIL.n0 60.0588
R100 VTAIL.n19 VTAIL.n18 60.0588
R101 VTAIL.n21 VTAIL.n20 60.0588
R102 VTAIL.t18 VTAIL.n65 52.3082
R103 VTAIL.t2 VTAIL.n5 52.3082
R104 VTAIL.t8 VTAIL.n49 52.3082
R105 VTAIL.t12 VTAIL.n29 52.3082
R106 VTAIL.n77 VTAIL.n76 30.052
R107 VTAIL.n17 VTAIL.n16 30.052
R108 VTAIL.n61 VTAIL.n60 30.052
R109 VTAIL.n41 VTAIL.n40 30.052
R110 VTAIL.n23 VTAIL.n21 17.5996
R111 VTAIL.n77 VTAIL.n61 16.4358
R112 VTAIL.n67 VTAIL.n66 10.2326
R113 VTAIL.n7 VTAIL.n6 10.2326
R114 VTAIL.n51 VTAIL.n50 10.2326
R115 VTAIL.n31 VTAIL.n30 10.2326
R116 VTAIL.n76 VTAIL.n62 9.69747
R117 VTAIL.n16 VTAIL.n2 9.69747
R118 VTAIL.n60 VTAIL.n46 9.69747
R119 VTAIL.n40 VTAIL.n26 9.69747
R120 VTAIL.n76 VTAIL.n75 9.45567
R121 VTAIL.n16 VTAIL.n15 9.45567
R122 VTAIL.n60 VTAIL.n59 9.45567
R123 VTAIL.n40 VTAIL.n39 9.45567
R124 VTAIL.n69 VTAIL.n68 9.3005
R125 VTAIL.n64 VTAIL.n63 9.3005
R126 VTAIL.n75 VTAIL.n74 9.3005
R127 VTAIL.n9 VTAIL.n8 9.3005
R128 VTAIL.n4 VTAIL.n3 9.3005
R129 VTAIL.n15 VTAIL.n14 9.3005
R130 VTAIL.n48 VTAIL.n47 9.3005
R131 VTAIL.n53 VTAIL.n52 9.3005
R132 VTAIL.n59 VTAIL.n58 9.3005
R133 VTAIL.n28 VTAIL.n27 9.3005
R134 VTAIL.n39 VTAIL.n38 9.3005
R135 VTAIL.n33 VTAIL.n32 9.3005
R136 VTAIL.n74 VTAIL.n73 8.92171
R137 VTAIL.n14 VTAIL.n13 8.92171
R138 VTAIL.n58 VTAIL.n57 8.92171
R139 VTAIL.n38 VTAIL.n37 8.92171
R140 VTAIL.n70 VTAIL.n64 8.14595
R141 VTAIL.n10 VTAIL.n4 8.14595
R142 VTAIL.n54 VTAIL.n48 8.14595
R143 VTAIL.n34 VTAIL.n28 8.14595
R144 VTAIL.n69 VTAIL.n66 7.3702
R145 VTAIL.n9 VTAIL.n6 7.3702
R146 VTAIL.n53 VTAIL.n50 7.3702
R147 VTAIL.n33 VTAIL.n30 7.3702
R148 VTAIL.n78 VTAIL.t11 5.87587
R149 VTAIL.n78 VTAIL.t17 5.87587
R150 VTAIL.n0 VTAIL.t14 5.87587
R151 VTAIL.n0 VTAIL.t16 5.87587
R152 VTAIL.n18 VTAIL.t1 5.87587
R153 VTAIL.n18 VTAIL.t7 5.87587
R154 VTAIL.n20 VTAIL.t6 5.87587
R155 VTAIL.n20 VTAIL.t0 5.87587
R156 VTAIL.n44 VTAIL.t3 5.87587
R157 VTAIL.n44 VTAIL.t4 5.87587
R158 VTAIL.n42 VTAIL.t9 5.87587
R159 VTAIL.n42 VTAIL.t5 5.87587
R160 VTAIL.n24 VTAIL.t19 5.87587
R161 VTAIL.n24 VTAIL.t15 5.87587
R162 VTAIL.n22 VTAIL.t10 5.87587
R163 VTAIL.n22 VTAIL.t13 5.87587
R164 VTAIL.n70 VTAIL.n69 5.81868
R165 VTAIL.n10 VTAIL.n9 5.81868
R166 VTAIL.n54 VTAIL.n53 5.81868
R167 VTAIL.n34 VTAIL.n33 5.81868
R168 VTAIL.n73 VTAIL.n64 5.04292
R169 VTAIL.n13 VTAIL.n4 5.04292
R170 VTAIL.n57 VTAIL.n48 5.04292
R171 VTAIL.n37 VTAIL.n28 5.04292
R172 VTAIL.n74 VTAIL.n62 4.26717
R173 VTAIL.n14 VTAIL.n2 4.26717
R174 VTAIL.n58 VTAIL.n46 4.26717
R175 VTAIL.n38 VTAIL.n26 4.26717
R176 VTAIL.n68 VTAIL.n67 2.88718
R177 VTAIL.n8 VTAIL.n7 2.88718
R178 VTAIL.n52 VTAIL.n51 2.88718
R179 VTAIL.n32 VTAIL.n31 2.88718
R180 VTAIL.n25 VTAIL.n23 1.16429
R181 VTAIL.n41 VTAIL.n25 1.16429
R182 VTAIL.n45 VTAIL.n43 1.16429
R183 VTAIL.n61 VTAIL.n45 1.16429
R184 VTAIL.n21 VTAIL.n19 1.16429
R185 VTAIL.n19 VTAIL.n17 1.16429
R186 VTAIL.n79 VTAIL.n77 1.16429
R187 VTAIL.n43 VTAIL.n41 1.05222
R188 VTAIL.n17 VTAIL.n1 1.05222
R189 VTAIL VTAIL.n1 0.931535
R190 VTAIL VTAIL.n79 0.233259
R191 VTAIL.n68 VTAIL.n63 0.155672
R192 VTAIL.n75 VTAIL.n63 0.155672
R193 VTAIL.n8 VTAIL.n3 0.155672
R194 VTAIL.n15 VTAIL.n3 0.155672
R195 VTAIL.n59 VTAIL.n47 0.155672
R196 VTAIL.n52 VTAIL.n47 0.155672
R197 VTAIL.n39 VTAIL.n27 0.155672
R198 VTAIL.n32 VTAIL.n27 0.155672
R199 VDD2.n29 VDD2.n19 289.615
R200 VDD2.n10 VDD2.n0 289.615
R201 VDD2.n30 VDD2.n29 185
R202 VDD2.n28 VDD2.n27 185
R203 VDD2.n23 VDD2.n22 185
R204 VDD2.n4 VDD2.n3 185
R205 VDD2.n9 VDD2.n8 185
R206 VDD2.n11 VDD2.n10 185
R207 VDD2.n24 VDD2.t1 150.499
R208 VDD2.n5 VDD2.t3 150.499
R209 VDD2.n29 VDD2.n28 104.615
R210 VDD2.n28 VDD2.n22 104.615
R211 VDD2.n9 VDD2.n3 104.615
R212 VDD2.n10 VDD2.n9 104.615
R213 VDD2.n18 VDD2.n17 77.5551
R214 VDD2 VDD2.n37 77.5522
R215 VDD2.n36 VDD2.n35 76.7376
R216 VDD2.n16 VDD2.n15 76.7376
R217 VDD2.t1 VDD2.n22 52.3082
R218 VDD2.t3 VDD2.n3 52.3082
R219 VDD2.n16 VDD2.n14 47.8946
R220 VDD2.n34 VDD2.n33 46.7308
R221 VDD2.n34 VDD2.n18 32.1485
R222 VDD2.n24 VDD2.n23 10.2326
R223 VDD2.n5 VDD2.n4 10.2326
R224 VDD2.n33 VDD2.n19 9.69747
R225 VDD2.n14 VDD2.n0 9.69747
R226 VDD2.n33 VDD2.n32 9.45567
R227 VDD2.n14 VDD2.n13 9.45567
R228 VDD2.n21 VDD2.n20 9.3005
R229 VDD2.n32 VDD2.n31 9.3005
R230 VDD2.n26 VDD2.n25 9.3005
R231 VDD2.n7 VDD2.n6 9.3005
R232 VDD2.n2 VDD2.n1 9.3005
R233 VDD2.n13 VDD2.n12 9.3005
R234 VDD2.n31 VDD2.n30 8.92171
R235 VDD2.n12 VDD2.n11 8.92171
R236 VDD2.n27 VDD2.n21 8.14595
R237 VDD2.n8 VDD2.n2 8.14595
R238 VDD2.n26 VDD2.n23 7.3702
R239 VDD2.n7 VDD2.n4 7.3702
R240 VDD2.n37 VDD2.t5 5.87587
R241 VDD2.n37 VDD2.t2 5.87587
R242 VDD2.n35 VDD2.t0 5.87587
R243 VDD2.n35 VDD2.t7 5.87587
R244 VDD2.n17 VDD2.t4 5.87587
R245 VDD2.n17 VDD2.t9 5.87587
R246 VDD2.n15 VDD2.t8 5.87587
R247 VDD2.n15 VDD2.t6 5.87587
R248 VDD2.n27 VDD2.n26 5.81868
R249 VDD2.n8 VDD2.n7 5.81868
R250 VDD2.n30 VDD2.n21 5.04292
R251 VDD2.n11 VDD2.n2 5.04292
R252 VDD2.n31 VDD2.n19 4.26717
R253 VDD2.n12 VDD2.n0 4.26717
R254 VDD2.n25 VDD2.n24 2.88718
R255 VDD2.n6 VDD2.n5 2.88718
R256 VDD2.n36 VDD2.n34 1.16429
R257 VDD2 VDD2.n36 0.349638
R258 VDD2.n18 VDD2.n16 0.236102
R259 VDD2.n32 VDD2.n20 0.155672
R260 VDD2.n25 VDD2.n20 0.155672
R261 VDD2.n6 VDD2.n1 0.155672
R262 VDD2.n13 VDD2.n1 0.155672
R263 B.n478 B.n477 585
R264 B.n167 B.n82 585
R265 B.n166 B.n165 585
R266 B.n164 B.n163 585
R267 B.n162 B.n161 585
R268 B.n160 B.n159 585
R269 B.n158 B.n157 585
R270 B.n156 B.n155 585
R271 B.n154 B.n153 585
R272 B.n152 B.n151 585
R273 B.n150 B.n149 585
R274 B.n148 B.n147 585
R275 B.n146 B.n145 585
R276 B.n144 B.n143 585
R277 B.n142 B.n141 585
R278 B.n140 B.n139 585
R279 B.n138 B.n137 585
R280 B.n136 B.n135 585
R281 B.n134 B.n133 585
R282 B.n132 B.n131 585
R283 B.n130 B.n129 585
R284 B.n128 B.n127 585
R285 B.n126 B.n125 585
R286 B.n124 B.n123 585
R287 B.n122 B.n121 585
R288 B.n120 B.n119 585
R289 B.n118 B.n117 585
R290 B.n116 B.n115 585
R291 B.n114 B.n113 585
R292 B.n112 B.n111 585
R293 B.n110 B.n109 585
R294 B.n108 B.n107 585
R295 B.n106 B.n105 585
R296 B.n104 B.n103 585
R297 B.n102 B.n101 585
R298 B.n100 B.n99 585
R299 B.n98 B.n97 585
R300 B.n96 B.n95 585
R301 B.n94 B.n93 585
R302 B.n92 B.n91 585
R303 B.n90 B.n89 585
R304 B.n60 B.n59 585
R305 B.n476 B.n61 585
R306 B.n481 B.n61 585
R307 B.n475 B.n474 585
R308 B.n474 B.n57 585
R309 B.n473 B.n56 585
R310 B.n487 B.n56 585
R311 B.n472 B.n55 585
R312 B.n488 B.n55 585
R313 B.n471 B.n54 585
R314 B.n489 B.n54 585
R315 B.n470 B.n469 585
R316 B.n469 B.n53 585
R317 B.n468 B.n49 585
R318 B.n495 B.n49 585
R319 B.n467 B.n48 585
R320 B.n496 B.n48 585
R321 B.n466 B.n47 585
R322 B.n497 B.n47 585
R323 B.n465 B.n464 585
R324 B.n464 B.n43 585
R325 B.n463 B.n42 585
R326 B.n503 B.n42 585
R327 B.n462 B.n41 585
R328 B.n504 B.n41 585
R329 B.n461 B.n40 585
R330 B.n505 B.n40 585
R331 B.n460 B.n459 585
R332 B.n459 B.n36 585
R333 B.n458 B.n35 585
R334 B.n511 B.n35 585
R335 B.n457 B.n34 585
R336 B.n512 B.n34 585
R337 B.n456 B.n33 585
R338 B.n513 B.n33 585
R339 B.n455 B.n454 585
R340 B.n454 B.n29 585
R341 B.n453 B.n28 585
R342 B.n519 B.n28 585
R343 B.n452 B.n27 585
R344 B.n520 B.n27 585
R345 B.n451 B.n26 585
R346 B.n521 B.n26 585
R347 B.n450 B.n449 585
R348 B.n449 B.n22 585
R349 B.n448 B.n21 585
R350 B.n527 B.n21 585
R351 B.n447 B.n20 585
R352 B.n528 B.n20 585
R353 B.n446 B.n19 585
R354 B.n529 B.n19 585
R355 B.n445 B.n444 585
R356 B.n444 B.n15 585
R357 B.n443 B.n14 585
R358 B.n535 B.n14 585
R359 B.n442 B.n13 585
R360 B.n536 B.n13 585
R361 B.n441 B.n12 585
R362 B.n537 B.n12 585
R363 B.n440 B.n439 585
R364 B.n439 B.n8 585
R365 B.n438 B.n7 585
R366 B.n543 B.n7 585
R367 B.n437 B.n6 585
R368 B.n544 B.n6 585
R369 B.n436 B.n5 585
R370 B.n545 B.n5 585
R371 B.n435 B.n434 585
R372 B.n434 B.n4 585
R373 B.n433 B.n168 585
R374 B.n433 B.n432 585
R375 B.n423 B.n169 585
R376 B.n170 B.n169 585
R377 B.n425 B.n424 585
R378 B.n426 B.n425 585
R379 B.n422 B.n175 585
R380 B.n175 B.n174 585
R381 B.n421 B.n420 585
R382 B.n420 B.n419 585
R383 B.n177 B.n176 585
R384 B.n178 B.n177 585
R385 B.n412 B.n411 585
R386 B.n413 B.n412 585
R387 B.n410 B.n183 585
R388 B.n183 B.n182 585
R389 B.n409 B.n408 585
R390 B.n408 B.n407 585
R391 B.n185 B.n184 585
R392 B.n186 B.n185 585
R393 B.n400 B.n399 585
R394 B.n401 B.n400 585
R395 B.n398 B.n191 585
R396 B.n191 B.n190 585
R397 B.n397 B.n396 585
R398 B.n396 B.n395 585
R399 B.n193 B.n192 585
R400 B.n194 B.n193 585
R401 B.n388 B.n387 585
R402 B.n389 B.n388 585
R403 B.n386 B.n199 585
R404 B.n199 B.n198 585
R405 B.n385 B.n384 585
R406 B.n384 B.n383 585
R407 B.n201 B.n200 585
R408 B.n202 B.n201 585
R409 B.n376 B.n375 585
R410 B.n377 B.n376 585
R411 B.n374 B.n207 585
R412 B.n207 B.n206 585
R413 B.n373 B.n372 585
R414 B.n372 B.n371 585
R415 B.n209 B.n208 585
R416 B.n210 B.n209 585
R417 B.n364 B.n363 585
R418 B.n365 B.n364 585
R419 B.n362 B.n215 585
R420 B.n215 B.n214 585
R421 B.n361 B.n360 585
R422 B.n360 B.n359 585
R423 B.n217 B.n216 585
R424 B.n352 B.n217 585
R425 B.n351 B.n350 585
R426 B.n353 B.n351 585
R427 B.n349 B.n222 585
R428 B.n222 B.n221 585
R429 B.n348 B.n347 585
R430 B.n347 B.n346 585
R431 B.n224 B.n223 585
R432 B.n225 B.n224 585
R433 B.n339 B.n338 585
R434 B.n340 B.n339 585
R435 B.n228 B.n227 585
R436 B.n255 B.n253 585
R437 B.n256 B.n252 585
R438 B.n256 B.n229 585
R439 B.n259 B.n258 585
R440 B.n260 B.n251 585
R441 B.n262 B.n261 585
R442 B.n264 B.n250 585
R443 B.n267 B.n266 585
R444 B.n268 B.n249 585
R445 B.n270 B.n269 585
R446 B.n272 B.n248 585
R447 B.n275 B.n274 585
R448 B.n276 B.n247 585
R449 B.n278 B.n277 585
R450 B.n280 B.n246 585
R451 B.n283 B.n282 585
R452 B.n285 B.n243 585
R453 B.n287 B.n286 585
R454 B.n289 B.n242 585
R455 B.n292 B.n291 585
R456 B.n293 B.n241 585
R457 B.n295 B.n294 585
R458 B.n297 B.n240 585
R459 B.n300 B.n299 585
R460 B.n301 B.n239 585
R461 B.n306 B.n305 585
R462 B.n308 B.n238 585
R463 B.n311 B.n310 585
R464 B.n312 B.n237 585
R465 B.n314 B.n313 585
R466 B.n316 B.n236 585
R467 B.n319 B.n318 585
R468 B.n320 B.n235 585
R469 B.n322 B.n321 585
R470 B.n324 B.n234 585
R471 B.n327 B.n326 585
R472 B.n328 B.n233 585
R473 B.n330 B.n329 585
R474 B.n332 B.n232 585
R475 B.n333 B.n231 585
R476 B.n336 B.n335 585
R477 B.n337 B.n230 585
R478 B.n230 B.n229 585
R479 B.n342 B.n341 585
R480 B.n341 B.n340 585
R481 B.n343 B.n226 585
R482 B.n226 B.n225 585
R483 B.n345 B.n344 585
R484 B.n346 B.n345 585
R485 B.n220 B.n219 585
R486 B.n221 B.n220 585
R487 B.n355 B.n354 585
R488 B.n354 B.n353 585
R489 B.n356 B.n218 585
R490 B.n352 B.n218 585
R491 B.n358 B.n357 585
R492 B.n359 B.n358 585
R493 B.n213 B.n212 585
R494 B.n214 B.n213 585
R495 B.n367 B.n366 585
R496 B.n366 B.n365 585
R497 B.n368 B.n211 585
R498 B.n211 B.n210 585
R499 B.n370 B.n369 585
R500 B.n371 B.n370 585
R501 B.n205 B.n204 585
R502 B.n206 B.n205 585
R503 B.n379 B.n378 585
R504 B.n378 B.n377 585
R505 B.n380 B.n203 585
R506 B.n203 B.n202 585
R507 B.n382 B.n381 585
R508 B.n383 B.n382 585
R509 B.n197 B.n196 585
R510 B.n198 B.n197 585
R511 B.n391 B.n390 585
R512 B.n390 B.n389 585
R513 B.n392 B.n195 585
R514 B.n195 B.n194 585
R515 B.n394 B.n393 585
R516 B.n395 B.n394 585
R517 B.n189 B.n188 585
R518 B.n190 B.n189 585
R519 B.n403 B.n402 585
R520 B.n402 B.n401 585
R521 B.n404 B.n187 585
R522 B.n187 B.n186 585
R523 B.n406 B.n405 585
R524 B.n407 B.n406 585
R525 B.n181 B.n180 585
R526 B.n182 B.n181 585
R527 B.n415 B.n414 585
R528 B.n414 B.n413 585
R529 B.n416 B.n179 585
R530 B.n179 B.n178 585
R531 B.n418 B.n417 585
R532 B.n419 B.n418 585
R533 B.n173 B.n172 585
R534 B.n174 B.n173 585
R535 B.n428 B.n427 585
R536 B.n427 B.n426 585
R537 B.n429 B.n171 585
R538 B.n171 B.n170 585
R539 B.n431 B.n430 585
R540 B.n432 B.n431 585
R541 B.n2 B.n0 585
R542 B.n4 B.n2 585
R543 B.n3 B.n1 585
R544 B.n544 B.n3 585
R545 B.n542 B.n541 585
R546 B.n543 B.n542 585
R547 B.n540 B.n9 585
R548 B.n9 B.n8 585
R549 B.n539 B.n538 585
R550 B.n538 B.n537 585
R551 B.n11 B.n10 585
R552 B.n536 B.n11 585
R553 B.n534 B.n533 585
R554 B.n535 B.n534 585
R555 B.n532 B.n16 585
R556 B.n16 B.n15 585
R557 B.n531 B.n530 585
R558 B.n530 B.n529 585
R559 B.n18 B.n17 585
R560 B.n528 B.n18 585
R561 B.n526 B.n525 585
R562 B.n527 B.n526 585
R563 B.n524 B.n23 585
R564 B.n23 B.n22 585
R565 B.n523 B.n522 585
R566 B.n522 B.n521 585
R567 B.n25 B.n24 585
R568 B.n520 B.n25 585
R569 B.n518 B.n517 585
R570 B.n519 B.n518 585
R571 B.n516 B.n30 585
R572 B.n30 B.n29 585
R573 B.n515 B.n514 585
R574 B.n514 B.n513 585
R575 B.n32 B.n31 585
R576 B.n512 B.n32 585
R577 B.n510 B.n509 585
R578 B.n511 B.n510 585
R579 B.n508 B.n37 585
R580 B.n37 B.n36 585
R581 B.n507 B.n506 585
R582 B.n506 B.n505 585
R583 B.n39 B.n38 585
R584 B.n504 B.n39 585
R585 B.n502 B.n501 585
R586 B.n503 B.n502 585
R587 B.n500 B.n44 585
R588 B.n44 B.n43 585
R589 B.n499 B.n498 585
R590 B.n498 B.n497 585
R591 B.n46 B.n45 585
R592 B.n496 B.n46 585
R593 B.n494 B.n493 585
R594 B.n495 B.n494 585
R595 B.n492 B.n50 585
R596 B.n53 B.n50 585
R597 B.n491 B.n490 585
R598 B.n490 B.n489 585
R599 B.n52 B.n51 585
R600 B.n488 B.n52 585
R601 B.n486 B.n485 585
R602 B.n487 B.n486 585
R603 B.n484 B.n58 585
R604 B.n58 B.n57 585
R605 B.n483 B.n482 585
R606 B.n482 B.n481 585
R607 B.n547 B.n546 585
R608 B.n546 B.n545 585
R609 B.n341 B.n228 492.5
R610 B.n482 B.n60 492.5
R611 B.n339 B.n230 492.5
R612 B.n478 B.n61 492.5
R613 B.n302 B.t14 282.685
R614 B.n244 B.t18 282.685
R615 B.n86 B.t21 282.685
R616 B.n83 B.t10 282.685
R617 B.n480 B.n479 256.663
R618 B.n480 B.n81 256.663
R619 B.n480 B.n80 256.663
R620 B.n480 B.n79 256.663
R621 B.n480 B.n78 256.663
R622 B.n480 B.n77 256.663
R623 B.n480 B.n76 256.663
R624 B.n480 B.n75 256.663
R625 B.n480 B.n74 256.663
R626 B.n480 B.n73 256.663
R627 B.n480 B.n72 256.663
R628 B.n480 B.n71 256.663
R629 B.n480 B.n70 256.663
R630 B.n480 B.n69 256.663
R631 B.n480 B.n68 256.663
R632 B.n480 B.n67 256.663
R633 B.n480 B.n66 256.663
R634 B.n480 B.n65 256.663
R635 B.n480 B.n64 256.663
R636 B.n480 B.n63 256.663
R637 B.n480 B.n62 256.663
R638 B.n254 B.n229 256.663
R639 B.n257 B.n229 256.663
R640 B.n263 B.n229 256.663
R641 B.n265 B.n229 256.663
R642 B.n271 B.n229 256.663
R643 B.n273 B.n229 256.663
R644 B.n279 B.n229 256.663
R645 B.n281 B.n229 256.663
R646 B.n288 B.n229 256.663
R647 B.n290 B.n229 256.663
R648 B.n296 B.n229 256.663
R649 B.n298 B.n229 256.663
R650 B.n307 B.n229 256.663
R651 B.n309 B.n229 256.663
R652 B.n315 B.n229 256.663
R653 B.n317 B.n229 256.663
R654 B.n323 B.n229 256.663
R655 B.n325 B.n229 256.663
R656 B.n331 B.n229 256.663
R657 B.n334 B.n229 256.663
R658 B.n341 B.n226 163.367
R659 B.n345 B.n226 163.367
R660 B.n345 B.n220 163.367
R661 B.n354 B.n220 163.367
R662 B.n354 B.n218 163.367
R663 B.n358 B.n218 163.367
R664 B.n358 B.n213 163.367
R665 B.n366 B.n213 163.367
R666 B.n366 B.n211 163.367
R667 B.n370 B.n211 163.367
R668 B.n370 B.n205 163.367
R669 B.n378 B.n205 163.367
R670 B.n378 B.n203 163.367
R671 B.n382 B.n203 163.367
R672 B.n382 B.n197 163.367
R673 B.n390 B.n197 163.367
R674 B.n390 B.n195 163.367
R675 B.n394 B.n195 163.367
R676 B.n394 B.n189 163.367
R677 B.n402 B.n189 163.367
R678 B.n402 B.n187 163.367
R679 B.n406 B.n187 163.367
R680 B.n406 B.n181 163.367
R681 B.n414 B.n181 163.367
R682 B.n414 B.n179 163.367
R683 B.n418 B.n179 163.367
R684 B.n418 B.n173 163.367
R685 B.n427 B.n173 163.367
R686 B.n427 B.n171 163.367
R687 B.n431 B.n171 163.367
R688 B.n431 B.n2 163.367
R689 B.n546 B.n2 163.367
R690 B.n546 B.n3 163.367
R691 B.n542 B.n3 163.367
R692 B.n542 B.n9 163.367
R693 B.n538 B.n9 163.367
R694 B.n538 B.n11 163.367
R695 B.n534 B.n11 163.367
R696 B.n534 B.n16 163.367
R697 B.n530 B.n16 163.367
R698 B.n530 B.n18 163.367
R699 B.n526 B.n18 163.367
R700 B.n526 B.n23 163.367
R701 B.n522 B.n23 163.367
R702 B.n522 B.n25 163.367
R703 B.n518 B.n25 163.367
R704 B.n518 B.n30 163.367
R705 B.n514 B.n30 163.367
R706 B.n514 B.n32 163.367
R707 B.n510 B.n32 163.367
R708 B.n510 B.n37 163.367
R709 B.n506 B.n37 163.367
R710 B.n506 B.n39 163.367
R711 B.n502 B.n39 163.367
R712 B.n502 B.n44 163.367
R713 B.n498 B.n44 163.367
R714 B.n498 B.n46 163.367
R715 B.n494 B.n46 163.367
R716 B.n494 B.n50 163.367
R717 B.n490 B.n50 163.367
R718 B.n490 B.n52 163.367
R719 B.n486 B.n52 163.367
R720 B.n486 B.n58 163.367
R721 B.n482 B.n58 163.367
R722 B.n256 B.n255 163.367
R723 B.n258 B.n256 163.367
R724 B.n262 B.n251 163.367
R725 B.n266 B.n264 163.367
R726 B.n270 B.n249 163.367
R727 B.n274 B.n272 163.367
R728 B.n278 B.n247 163.367
R729 B.n282 B.n280 163.367
R730 B.n287 B.n243 163.367
R731 B.n291 B.n289 163.367
R732 B.n295 B.n241 163.367
R733 B.n299 B.n297 163.367
R734 B.n306 B.n239 163.367
R735 B.n310 B.n308 163.367
R736 B.n314 B.n237 163.367
R737 B.n318 B.n316 163.367
R738 B.n322 B.n235 163.367
R739 B.n326 B.n324 163.367
R740 B.n330 B.n233 163.367
R741 B.n333 B.n332 163.367
R742 B.n335 B.n230 163.367
R743 B.n339 B.n224 163.367
R744 B.n347 B.n224 163.367
R745 B.n347 B.n222 163.367
R746 B.n351 B.n222 163.367
R747 B.n351 B.n217 163.367
R748 B.n360 B.n217 163.367
R749 B.n360 B.n215 163.367
R750 B.n364 B.n215 163.367
R751 B.n364 B.n209 163.367
R752 B.n372 B.n209 163.367
R753 B.n372 B.n207 163.367
R754 B.n376 B.n207 163.367
R755 B.n376 B.n201 163.367
R756 B.n384 B.n201 163.367
R757 B.n384 B.n199 163.367
R758 B.n388 B.n199 163.367
R759 B.n388 B.n193 163.367
R760 B.n396 B.n193 163.367
R761 B.n396 B.n191 163.367
R762 B.n400 B.n191 163.367
R763 B.n400 B.n185 163.367
R764 B.n408 B.n185 163.367
R765 B.n408 B.n183 163.367
R766 B.n412 B.n183 163.367
R767 B.n412 B.n177 163.367
R768 B.n420 B.n177 163.367
R769 B.n420 B.n175 163.367
R770 B.n425 B.n175 163.367
R771 B.n425 B.n169 163.367
R772 B.n433 B.n169 163.367
R773 B.n434 B.n433 163.367
R774 B.n434 B.n5 163.367
R775 B.n6 B.n5 163.367
R776 B.n7 B.n6 163.367
R777 B.n439 B.n7 163.367
R778 B.n439 B.n12 163.367
R779 B.n13 B.n12 163.367
R780 B.n14 B.n13 163.367
R781 B.n444 B.n14 163.367
R782 B.n444 B.n19 163.367
R783 B.n20 B.n19 163.367
R784 B.n21 B.n20 163.367
R785 B.n449 B.n21 163.367
R786 B.n449 B.n26 163.367
R787 B.n27 B.n26 163.367
R788 B.n28 B.n27 163.367
R789 B.n454 B.n28 163.367
R790 B.n454 B.n33 163.367
R791 B.n34 B.n33 163.367
R792 B.n35 B.n34 163.367
R793 B.n459 B.n35 163.367
R794 B.n459 B.n40 163.367
R795 B.n41 B.n40 163.367
R796 B.n42 B.n41 163.367
R797 B.n464 B.n42 163.367
R798 B.n464 B.n47 163.367
R799 B.n48 B.n47 163.367
R800 B.n49 B.n48 163.367
R801 B.n469 B.n49 163.367
R802 B.n469 B.n54 163.367
R803 B.n55 B.n54 163.367
R804 B.n56 B.n55 163.367
R805 B.n474 B.n56 163.367
R806 B.n474 B.n61 163.367
R807 B.n91 B.n90 163.367
R808 B.n95 B.n94 163.367
R809 B.n99 B.n98 163.367
R810 B.n103 B.n102 163.367
R811 B.n107 B.n106 163.367
R812 B.n111 B.n110 163.367
R813 B.n115 B.n114 163.367
R814 B.n119 B.n118 163.367
R815 B.n123 B.n122 163.367
R816 B.n127 B.n126 163.367
R817 B.n131 B.n130 163.367
R818 B.n135 B.n134 163.367
R819 B.n139 B.n138 163.367
R820 B.n143 B.n142 163.367
R821 B.n147 B.n146 163.367
R822 B.n151 B.n150 163.367
R823 B.n155 B.n154 163.367
R824 B.n159 B.n158 163.367
R825 B.n163 B.n162 163.367
R826 B.n165 B.n82 163.367
R827 B.n302 B.t17 161.659
R828 B.n83 B.t12 161.659
R829 B.n244 B.t20 161.659
R830 B.n86 B.t22 161.659
R831 B.n340 B.n229 151.417
R832 B.n481 B.n480 151.417
R833 B.n303 B.t16 135.476
R834 B.n84 B.t13 135.476
R835 B.n245 B.t19 135.476
R836 B.n87 B.t23 135.476
R837 B.n340 B.n225 86.5245
R838 B.n346 B.n225 86.5245
R839 B.n346 B.n221 86.5245
R840 B.n353 B.n221 86.5245
R841 B.n353 B.n352 86.5245
R842 B.n359 B.n214 86.5245
R843 B.n365 B.n214 86.5245
R844 B.n365 B.n210 86.5245
R845 B.n371 B.n210 86.5245
R846 B.n371 B.n206 86.5245
R847 B.n377 B.n206 86.5245
R848 B.n383 B.n202 86.5245
R849 B.n383 B.n198 86.5245
R850 B.n389 B.n198 86.5245
R851 B.n395 B.n194 86.5245
R852 B.n395 B.n190 86.5245
R853 B.n401 B.n190 86.5245
R854 B.n407 B.n186 86.5245
R855 B.n407 B.n182 86.5245
R856 B.n413 B.n182 86.5245
R857 B.n419 B.n178 86.5245
R858 B.n419 B.n174 86.5245
R859 B.n426 B.n174 86.5245
R860 B.n432 B.n170 86.5245
R861 B.n432 B.n4 86.5245
R862 B.n545 B.n4 86.5245
R863 B.n545 B.n544 86.5245
R864 B.n544 B.n543 86.5245
R865 B.n543 B.n8 86.5245
R866 B.n537 B.n536 86.5245
R867 B.n536 B.n535 86.5245
R868 B.n535 B.n15 86.5245
R869 B.n529 B.n528 86.5245
R870 B.n528 B.n527 86.5245
R871 B.n527 B.n22 86.5245
R872 B.n521 B.n520 86.5245
R873 B.n520 B.n519 86.5245
R874 B.n519 B.n29 86.5245
R875 B.n513 B.n512 86.5245
R876 B.n512 B.n511 86.5245
R877 B.n511 B.n36 86.5245
R878 B.n505 B.n504 86.5245
R879 B.n504 B.n503 86.5245
R880 B.n503 B.n43 86.5245
R881 B.n497 B.n43 86.5245
R882 B.n497 B.n496 86.5245
R883 B.n496 B.n495 86.5245
R884 B.n489 B.n53 86.5245
R885 B.n489 B.n488 86.5245
R886 B.n488 B.n487 86.5245
R887 B.n487 B.n57 86.5245
R888 B.n481 B.n57 86.5245
R889 B.n254 B.n228 71.676
R890 B.n258 B.n257 71.676
R891 B.n263 B.n262 71.676
R892 B.n266 B.n265 71.676
R893 B.n271 B.n270 71.676
R894 B.n274 B.n273 71.676
R895 B.n279 B.n278 71.676
R896 B.n282 B.n281 71.676
R897 B.n288 B.n287 71.676
R898 B.n291 B.n290 71.676
R899 B.n296 B.n295 71.676
R900 B.n299 B.n298 71.676
R901 B.n307 B.n306 71.676
R902 B.n310 B.n309 71.676
R903 B.n315 B.n314 71.676
R904 B.n318 B.n317 71.676
R905 B.n323 B.n322 71.676
R906 B.n326 B.n325 71.676
R907 B.n331 B.n330 71.676
R908 B.n334 B.n333 71.676
R909 B.n62 B.n60 71.676
R910 B.n91 B.n63 71.676
R911 B.n95 B.n64 71.676
R912 B.n99 B.n65 71.676
R913 B.n103 B.n66 71.676
R914 B.n107 B.n67 71.676
R915 B.n111 B.n68 71.676
R916 B.n115 B.n69 71.676
R917 B.n119 B.n70 71.676
R918 B.n123 B.n71 71.676
R919 B.n127 B.n72 71.676
R920 B.n131 B.n73 71.676
R921 B.n135 B.n74 71.676
R922 B.n139 B.n75 71.676
R923 B.n143 B.n76 71.676
R924 B.n147 B.n77 71.676
R925 B.n151 B.n78 71.676
R926 B.n155 B.n79 71.676
R927 B.n159 B.n80 71.676
R928 B.n163 B.n81 71.676
R929 B.n479 B.n82 71.676
R930 B.n479 B.n478 71.676
R931 B.n165 B.n81 71.676
R932 B.n162 B.n80 71.676
R933 B.n158 B.n79 71.676
R934 B.n154 B.n78 71.676
R935 B.n150 B.n77 71.676
R936 B.n146 B.n76 71.676
R937 B.n142 B.n75 71.676
R938 B.n138 B.n74 71.676
R939 B.n134 B.n73 71.676
R940 B.n130 B.n72 71.676
R941 B.n126 B.n71 71.676
R942 B.n122 B.n70 71.676
R943 B.n118 B.n69 71.676
R944 B.n114 B.n68 71.676
R945 B.n110 B.n67 71.676
R946 B.n106 B.n66 71.676
R947 B.n102 B.n65 71.676
R948 B.n98 B.n64 71.676
R949 B.n94 B.n63 71.676
R950 B.n90 B.n62 71.676
R951 B.n255 B.n254 71.676
R952 B.n257 B.n251 71.676
R953 B.n264 B.n263 71.676
R954 B.n265 B.n249 71.676
R955 B.n272 B.n271 71.676
R956 B.n273 B.n247 71.676
R957 B.n280 B.n279 71.676
R958 B.n281 B.n243 71.676
R959 B.n289 B.n288 71.676
R960 B.n290 B.n241 71.676
R961 B.n297 B.n296 71.676
R962 B.n298 B.n239 71.676
R963 B.n308 B.n307 71.676
R964 B.n309 B.n237 71.676
R965 B.n316 B.n315 71.676
R966 B.n317 B.n235 71.676
R967 B.n324 B.n323 71.676
R968 B.n325 B.n233 71.676
R969 B.n332 B.n331 71.676
R970 B.n335 B.n334 71.676
R971 B.n304 B.n303 59.5399
R972 B.n284 B.n245 59.5399
R973 B.n88 B.n87 59.5399
R974 B.n85 B.n84 59.5399
R975 B.n359 B.t15 55.9866
R976 B.n495 B.t11 55.9866
R977 B.t2 B.n170 50.897
R978 B.t9 B.n8 50.897
R979 B.t7 B.n178 48.3522
R980 B.t5 B.n15 48.3522
R981 B.n377 B.t6 45.8073
R982 B.t1 B.n186 45.8073
R983 B.t3 B.n22 45.8073
R984 B.n505 B.t8 45.8073
R985 B.n389 B.t0 43.2625
R986 B.t0 B.n194 43.2625
R987 B.t4 B.n29 43.2625
R988 B.n513 B.t4 43.2625
R989 B.t6 B.n202 40.7177
R990 B.n401 B.t1 40.7177
R991 B.n521 B.t3 40.7177
R992 B.t8 B.n36 40.7177
R993 B.n413 B.t7 38.1729
R994 B.n529 B.t5 38.1729
R995 B.n426 B.t2 35.628
R996 B.n537 B.t9 35.628
R997 B.n483 B.n59 32.0005
R998 B.n477 B.n476 32.0005
R999 B.n338 B.n337 32.0005
R1000 B.n342 B.n227 32.0005
R1001 B.n352 B.t15 30.5384
R1002 B.n53 B.t11 30.5384
R1003 B.n303 B.n302 26.1823
R1004 B.n245 B.n244 26.1823
R1005 B.n87 B.n86 26.1823
R1006 B.n84 B.n83 26.1823
R1007 B B.n547 18.0485
R1008 B.n89 B.n59 10.6151
R1009 B.n92 B.n89 10.6151
R1010 B.n93 B.n92 10.6151
R1011 B.n96 B.n93 10.6151
R1012 B.n97 B.n96 10.6151
R1013 B.n100 B.n97 10.6151
R1014 B.n101 B.n100 10.6151
R1015 B.n104 B.n101 10.6151
R1016 B.n105 B.n104 10.6151
R1017 B.n108 B.n105 10.6151
R1018 B.n109 B.n108 10.6151
R1019 B.n112 B.n109 10.6151
R1020 B.n113 B.n112 10.6151
R1021 B.n116 B.n113 10.6151
R1022 B.n117 B.n116 10.6151
R1023 B.n121 B.n120 10.6151
R1024 B.n124 B.n121 10.6151
R1025 B.n125 B.n124 10.6151
R1026 B.n128 B.n125 10.6151
R1027 B.n129 B.n128 10.6151
R1028 B.n132 B.n129 10.6151
R1029 B.n133 B.n132 10.6151
R1030 B.n136 B.n133 10.6151
R1031 B.n137 B.n136 10.6151
R1032 B.n141 B.n140 10.6151
R1033 B.n144 B.n141 10.6151
R1034 B.n145 B.n144 10.6151
R1035 B.n148 B.n145 10.6151
R1036 B.n149 B.n148 10.6151
R1037 B.n152 B.n149 10.6151
R1038 B.n153 B.n152 10.6151
R1039 B.n156 B.n153 10.6151
R1040 B.n157 B.n156 10.6151
R1041 B.n160 B.n157 10.6151
R1042 B.n161 B.n160 10.6151
R1043 B.n164 B.n161 10.6151
R1044 B.n166 B.n164 10.6151
R1045 B.n167 B.n166 10.6151
R1046 B.n477 B.n167 10.6151
R1047 B.n338 B.n223 10.6151
R1048 B.n348 B.n223 10.6151
R1049 B.n349 B.n348 10.6151
R1050 B.n350 B.n349 10.6151
R1051 B.n350 B.n216 10.6151
R1052 B.n361 B.n216 10.6151
R1053 B.n362 B.n361 10.6151
R1054 B.n363 B.n362 10.6151
R1055 B.n363 B.n208 10.6151
R1056 B.n373 B.n208 10.6151
R1057 B.n374 B.n373 10.6151
R1058 B.n375 B.n374 10.6151
R1059 B.n375 B.n200 10.6151
R1060 B.n385 B.n200 10.6151
R1061 B.n386 B.n385 10.6151
R1062 B.n387 B.n386 10.6151
R1063 B.n387 B.n192 10.6151
R1064 B.n397 B.n192 10.6151
R1065 B.n398 B.n397 10.6151
R1066 B.n399 B.n398 10.6151
R1067 B.n399 B.n184 10.6151
R1068 B.n409 B.n184 10.6151
R1069 B.n410 B.n409 10.6151
R1070 B.n411 B.n410 10.6151
R1071 B.n411 B.n176 10.6151
R1072 B.n421 B.n176 10.6151
R1073 B.n422 B.n421 10.6151
R1074 B.n424 B.n422 10.6151
R1075 B.n424 B.n423 10.6151
R1076 B.n423 B.n168 10.6151
R1077 B.n435 B.n168 10.6151
R1078 B.n436 B.n435 10.6151
R1079 B.n437 B.n436 10.6151
R1080 B.n438 B.n437 10.6151
R1081 B.n440 B.n438 10.6151
R1082 B.n441 B.n440 10.6151
R1083 B.n442 B.n441 10.6151
R1084 B.n443 B.n442 10.6151
R1085 B.n445 B.n443 10.6151
R1086 B.n446 B.n445 10.6151
R1087 B.n447 B.n446 10.6151
R1088 B.n448 B.n447 10.6151
R1089 B.n450 B.n448 10.6151
R1090 B.n451 B.n450 10.6151
R1091 B.n452 B.n451 10.6151
R1092 B.n453 B.n452 10.6151
R1093 B.n455 B.n453 10.6151
R1094 B.n456 B.n455 10.6151
R1095 B.n457 B.n456 10.6151
R1096 B.n458 B.n457 10.6151
R1097 B.n460 B.n458 10.6151
R1098 B.n461 B.n460 10.6151
R1099 B.n462 B.n461 10.6151
R1100 B.n463 B.n462 10.6151
R1101 B.n465 B.n463 10.6151
R1102 B.n466 B.n465 10.6151
R1103 B.n467 B.n466 10.6151
R1104 B.n468 B.n467 10.6151
R1105 B.n470 B.n468 10.6151
R1106 B.n471 B.n470 10.6151
R1107 B.n472 B.n471 10.6151
R1108 B.n473 B.n472 10.6151
R1109 B.n475 B.n473 10.6151
R1110 B.n476 B.n475 10.6151
R1111 B.n253 B.n227 10.6151
R1112 B.n253 B.n252 10.6151
R1113 B.n259 B.n252 10.6151
R1114 B.n260 B.n259 10.6151
R1115 B.n261 B.n260 10.6151
R1116 B.n261 B.n250 10.6151
R1117 B.n267 B.n250 10.6151
R1118 B.n268 B.n267 10.6151
R1119 B.n269 B.n268 10.6151
R1120 B.n269 B.n248 10.6151
R1121 B.n275 B.n248 10.6151
R1122 B.n276 B.n275 10.6151
R1123 B.n277 B.n276 10.6151
R1124 B.n277 B.n246 10.6151
R1125 B.n283 B.n246 10.6151
R1126 B.n286 B.n285 10.6151
R1127 B.n286 B.n242 10.6151
R1128 B.n292 B.n242 10.6151
R1129 B.n293 B.n292 10.6151
R1130 B.n294 B.n293 10.6151
R1131 B.n294 B.n240 10.6151
R1132 B.n300 B.n240 10.6151
R1133 B.n301 B.n300 10.6151
R1134 B.n305 B.n301 10.6151
R1135 B.n311 B.n238 10.6151
R1136 B.n312 B.n311 10.6151
R1137 B.n313 B.n312 10.6151
R1138 B.n313 B.n236 10.6151
R1139 B.n319 B.n236 10.6151
R1140 B.n320 B.n319 10.6151
R1141 B.n321 B.n320 10.6151
R1142 B.n321 B.n234 10.6151
R1143 B.n327 B.n234 10.6151
R1144 B.n328 B.n327 10.6151
R1145 B.n329 B.n328 10.6151
R1146 B.n329 B.n232 10.6151
R1147 B.n232 B.n231 10.6151
R1148 B.n336 B.n231 10.6151
R1149 B.n337 B.n336 10.6151
R1150 B.n343 B.n342 10.6151
R1151 B.n344 B.n343 10.6151
R1152 B.n344 B.n219 10.6151
R1153 B.n355 B.n219 10.6151
R1154 B.n356 B.n355 10.6151
R1155 B.n357 B.n356 10.6151
R1156 B.n357 B.n212 10.6151
R1157 B.n367 B.n212 10.6151
R1158 B.n368 B.n367 10.6151
R1159 B.n369 B.n368 10.6151
R1160 B.n369 B.n204 10.6151
R1161 B.n379 B.n204 10.6151
R1162 B.n380 B.n379 10.6151
R1163 B.n381 B.n380 10.6151
R1164 B.n381 B.n196 10.6151
R1165 B.n391 B.n196 10.6151
R1166 B.n392 B.n391 10.6151
R1167 B.n393 B.n392 10.6151
R1168 B.n393 B.n188 10.6151
R1169 B.n403 B.n188 10.6151
R1170 B.n404 B.n403 10.6151
R1171 B.n405 B.n404 10.6151
R1172 B.n405 B.n180 10.6151
R1173 B.n415 B.n180 10.6151
R1174 B.n416 B.n415 10.6151
R1175 B.n417 B.n416 10.6151
R1176 B.n417 B.n172 10.6151
R1177 B.n428 B.n172 10.6151
R1178 B.n429 B.n428 10.6151
R1179 B.n430 B.n429 10.6151
R1180 B.n430 B.n0 10.6151
R1181 B.n541 B.n1 10.6151
R1182 B.n541 B.n540 10.6151
R1183 B.n540 B.n539 10.6151
R1184 B.n539 B.n10 10.6151
R1185 B.n533 B.n10 10.6151
R1186 B.n533 B.n532 10.6151
R1187 B.n532 B.n531 10.6151
R1188 B.n531 B.n17 10.6151
R1189 B.n525 B.n17 10.6151
R1190 B.n525 B.n524 10.6151
R1191 B.n524 B.n523 10.6151
R1192 B.n523 B.n24 10.6151
R1193 B.n517 B.n24 10.6151
R1194 B.n517 B.n516 10.6151
R1195 B.n516 B.n515 10.6151
R1196 B.n515 B.n31 10.6151
R1197 B.n509 B.n31 10.6151
R1198 B.n509 B.n508 10.6151
R1199 B.n508 B.n507 10.6151
R1200 B.n507 B.n38 10.6151
R1201 B.n501 B.n38 10.6151
R1202 B.n501 B.n500 10.6151
R1203 B.n500 B.n499 10.6151
R1204 B.n499 B.n45 10.6151
R1205 B.n493 B.n45 10.6151
R1206 B.n493 B.n492 10.6151
R1207 B.n492 B.n491 10.6151
R1208 B.n491 B.n51 10.6151
R1209 B.n485 B.n51 10.6151
R1210 B.n485 B.n484 10.6151
R1211 B.n484 B.n483 10.6151
R1212 B.n117 B.n88 9.36635
R1213 B.n140 B.n85 9.36635
R1214 B.n284 B.n283 9.36635
R1215 B.n304 B.n238 9.36635
R1216 B.n547 B.n0 2.81026
R1217 B.n547 B.n1 2.81026
R1218 B.n120 B.n88 1.24928
R1219 B.n137 B.n85 1.24928
R1220 B.n285 B.n284 1.24928
R1221 B.n305 B.n304 1.24928
R1222 VP.n10 VP.n7 161.3
R1223 VP.n12 VP.n11 161.3
R1224 VP.n13 VP.n6 161.3
R1225 VP.n16 VP.n15 161.3
R1226 VP.n17 VP.n5 161.3
R1227 VP.n19 VP.n18 161.3
R1228 VP.n21 VP.n4 161.3
R1229 VP.n40 VP.n0 161.3
R1230 VP.n38 VP.n37 161.3
R1231 VP.n36 VP.n1 161.3
R1232 VP.n35 VP.n34 161.3
R1233 VP.n32 VP.n2 161.3
R1234 VP.n31 VP.n30 161.3
R1235 VP.n29 VP.n3 161.3
R1236 VP.n28 VP.n27 161.3
R1237 VP.n9 VP.t4 133.029
R1238 VP.n25 VP.t9 118.374
R1239 VP.n41 VP.t5 118.374
R1240 VP.n22 VP.t7 118.374
R1241 VP.n23 VP.n22 80.6037
R1242 VP.n42 VP.n41 80.6037
R1243 VP.n25 VP.n24 80.6037
R1244 VP.n26 VP.t6 79.625
R1245 VP.n33 VP.t2 79.625
R1246 VP.n39 VP.t1 79.625
R1247 VP.n20 VP.t8 79.625
R1248 VP.n14 VP.t0 79.625
R1249 VP.n8 VP.t3 79.625
R1250 VP.n27 VP.n25 53.5832
R1251 VP.n41 VP.n40 53.5832
R1252 VP.n22 VP.n21 53.5832
R1253 VP.n9 VP.n8 48.7962
R1254 VP.n32 VP.n31 47.7779
R1255 VP.n34 VP.n1 47.7779
R1256 VP.n15 VP.n5 47.7779
R1257 VP.n13 VP.n12 47.7779
R1258 VP.n10 VP.n9 44.3029
R1259 VP.n24 VP.n23 38.1718
R1260 VP.n31 VP.n3 33.2089
R1261 VP.n38 VP.n1 33.2089
R1262 VP.n19 VP.n5 33.2089
R1263 VP.n12 VP.n7 33.2089
R1264 VP.n27 VP.n26 19.5741
R1265 VP.n40 VP.n39 19.5741
R1266 VP.n21 VP.n20 19.5741
R1267 VP.n33 VP.n32 12.234
R1268 VP.n34 VP.n33 12.234
R1269 VP.n14 VP.n13 12.234
R1270 VP.n15 VP.n14 12.234
R1271 VP.n26 VP.n3 4.8939
R1272 VP.n39 VP.n38 4.8939
R1273 VP.n20 VP.n19 4.8939
R1274 VP.n8 VP.n7 4.8939
R1275 VP.n23 VP.n4 0.285035
R1276 VP.n28 VP.n24 0.285035
R1277 VP.n42 VP.n0 0.285035
R1278 VP.n11 VP.n10 0.189894
R1279 VP.n11 VP.n6 0.189894
R1280 VP.n16 VP.n6 0.189894
R1281 VP.n17 VP.n16 0.189894
R1282 VP.n18 VP.n17 0.189894
R1283 VP.n18 VP.n4 0.189894
R1284 VP.n29 VP.n28 0.189894
R1285 VP.n30 VP.n29 0.189894
R1286 VP.n30 VP.n2 0.189894
R1287 VP.n35 VP.n2 0.189894
R1288 VP.n36 VP.n35 0.189894
R1289 VP.n37 VP.n36 0.189894
R1290 VP.n37 VP.n0 0.189894
R1291 VP VP.n42 0.146778
R1292 VDD1.n10 VDD1.n0 289.615
R1293 VDD1.n27 VDD1.n17 289.615
R1294 VDD1.n11 VDD1.n10 185
R1295 VDD1.n9 VDD1.n8 185
R1296 VDD1.n4 VDD1.n3 185
R1297 VDD1.n21 VDD1.n20 185
R1298 VDD1.n26 VDD1.n25 185
R1299 VDD1.n28 VDD1.n27 185
R1300 VDD1.n5 VDD1.t5 150.499
R1301 VDD1.n22 VDD1.t0 150.499
R1302 VDD1.n10 VDD1.n9 104.615
R1303 VDD1.n9 VDD1.n3 104.615
R1304 VDD1.n26 VDD1.n20 104.615
R1305 VDD1.n27 VDD1.n26 104.615
R1306 VDD1.n35 VDD1.n34 77.5551
R1307 VDD1.n37 VDD1.n36 76.7376
R1308 VDD1.n16 VDD1.n15 76.7376
R1309 VDD1.n33 VDD1.n32 76.7376
R1310 VDD1.t5 VDD1.n3 52.3082
R1311 VDD1.t0 VDD1.n20 52.3082
R1312 VDD1.n16 VDD1.n14 47.8946
R1313 VDD1.n33 VDD1.n31 47.8946
R1314 VDD1.n37 VDD1.n35 33.3134
R1315 VDD1.n5 VDD1.n4 10.2326
R1316 VDD1.n22 VDD1.n21 10.2326
R1317 VDD1.n14 VDD1.n0 9.69747
R1318 VDD1.n31 VDD1.n17 9.69747
R1319 VDD1.n14 VDD1.n13 9.45567
R1320 VDD1.n31 VDD1.n30 9.45567
R1321 VDD1.n2 VDD1.n1 9.3005
R1322 VDD1.n13 VDD1.n12 9.3005
R1323 VDD1.n7 VDD1.n6 9.3005
R1324 VDD1.n24 VDD1.n23 9.3005
R1325 VDD1.n19 VDD1.n18 9.3005
R1326 VDD1.n30 VDD1.n29 9.3005
R1327 VDD1.n12 VDD1.n11 8.92171
R1328 VDD1.n29 VDD1.n28 8.92171
R1329 VDD1.n8 VDD1.n2 8.14595
R1330 VDD1.n25 VDD1.n19 8.14595
R1331 VDD1.n7 VDD1.n4 7.3702
R1332 VDD1.n24 VDD1.n21 7.3702
R1333 VDD1.n36 VDD1.t1 5.87587
R1334 VDD1.n36 VDD1.t2 5.87587
R1335 VDD1.n15 VDD1.t6 5.87587
R1336 VDD1.n15 VDD1.t9 5.87587
R1337 VDD1.n34 VDD1.t8 5.87587
R1338 VDD1.n34 VDD1.t4 5.87587
R1339 VDD1.n32 VDD1.t3 5.87587
R1340 VDD1.n32 VDD1.t7 5.87587
R1341 VDD1.n8 VDD1.n7 5.81868
R1342 VDD1.n25 VDD1.n24 5.81868
R1343 VDD1.n11 VDD1.n2 5.04292
R1344 VDD1.n28 VDD1.n19 5.04292
R1345 VDD1.n12 VDD1.n0 4.26717
R1346 VDD1.n29 VDD1.n17 4.26717
R1347 VDD1.n6 VDD1.n5 2.88718
R1348 VDD1.n23 VDD1.n22 2.88718
R1349 VDD1 VDD1.n37 0.815155
R1350 VDD1 VDD1.n16 0.349638
R1351 VDD1.n35 VDD1.n33 0.236102
R1352 VDD1.n13 VDD1.n1 0.155672
R1353 VDD1.n6 VDD1.n1 0.155672
R1354 VDD1.n23 VDD1.n18 0.155672
R1355 VDD1.n30 VDD1.n18 0.155672
C0 VN VP 4.47645f
C1 VDD2 VTAIL 5.5609f
C2 VDD2 VP 0.386437f
C3 VN VDD1 0.154539f
C4 VDD2 VDD1 1.17174f
C5 VDD2 VN 2.57779f
C6 VTAIL VP 3.03511f
C7 VTAIL VDD1 5.51943f
C8 VP VDD1 2.8073f
C9 VTAIL VN 3.02089f
C10 VDD2 B 3.803488f
C11 VDD1 B 3.743604f
C12 VTAIL B 3.393232f
C13 VN B 9.8645f
C14 VP B 8.318776f
C15 VDD1.n0 B 0.035017f
C16 VDD1.n1 B 0.023881f
C17 VDD1.n2 B 0.012833f
C18 VDD1.n3 B 0.022749f
C19 VDD1.n4 B 0.021237f
C20 VDD1.t5 B 0.053033f
C21 VDD1.n5 B 0.096182f
C22 VDD1.n6 B 0.282248f
C23 VDD1.n7 B 0.012833f
C24 VDD1.n8 B 0.013587f
C25 VDD1.n9 B 0.030332f
C26 VDD1.n10 B 0.068227f
C27 VDD1.n11 B 0.013587f
C28 VDD1.n12 B 0.012833f
C29 VDD1.n13 B 0.051611f
C30 VDD1.n14 B 0.05809f
C31 VDD1.t6 B 0.063597f
C32 VDD1.t9 B 0.063597f
C33 VDD1.n15 B 0.471868f
C34 VDD1.n16 B 0.440698f
C35 VDD1.n17 B 0.035017f
C36 VDD1.n18 B 0.023881f
C37 VDD1.n19 B 0.012833f
C38 VDD1.n20 B 0.022749f
C39 VDD1.n21 B 0.021237f
C40 VDD1.t0 B 0.053033f
C41 VDD1.n22 B 0.096182f
C42 VDD1.n23 B 0.282248f
C43 VDD1.n24 B 0.012833f
C44 VDD1.n25 B 0.013587f
C45 VDD1.n26 B 0.030332f
C46 VDD1.n27 B 0.068227f
C47 VDD1.n28 B 0.013587f
C48 VDD1.n29 B 0.012833f
C49 VDD1.n30 B 0.051611f
C50 VDD1.n31 B 0.05809f
C51 VDD1.t3 B 0.063597f
C52 VDD1.t7 B 0.063597f
C53 VDD1.n32 B 0.471866f
C54 VDD1.n33 B 0.434314f
C55 VDD1.t8 B 0.063597f
C56 VDD1.t4 B 0.063597f
C57 VDD1.n34 B 0.475627f
C58 VDD1.n35 B 1.56849f
C59 VDD1.t1 B 0.063597f
C60 VDD1.t2 B 0.063597f
C61 VDD1.n36 B 0.471868f
C62 VDD1.n37 B 1.75037f
C63 VP.n0 B 0.054298f
C64 VP.t1 B 0.353222f
C65 VP.n1 B 0.035935f
C66 VP.n2 B 0.040692f
C67 VP.t2 B 0.353222f
C68 VP.n3 B 0.052194f
C69 VP.n4 B 0.054298f
C70 VP.t7 B 0.416809f
C71 VP.t8 B 0.353222f
C72 VP.n5 B 0.035935f
C73 VP.n6 B 0.040692f
C74 VP.t0 B 0.353222f
C75 VP.n7 B 0.052194f
C76 VP.t3 B 0.353222f
C77 VP.n8 B 0.200448f
C78 VP.t4 B 0.442363f
C79 VP.n9 B 0.228641f
C80 VP.n10 B 0.172464f
C81 VP.n11 B 0.040692f
C82 VP.n12 B 0.035935f
C83 VP.n13 B 0.057849f
C84 VP.n14 B 0.168107f
C85 VP.n15 B 0.057849f
C86 VP.n16 B 0.040692f
C87 VP.n17 B 0.040692f
C88 VP.n18 B 0.040692f
C89 VP.n19 B 0.052194f
C90 VP.n20 B 0.168107f
C91 VP.n21 B 0.054003f
C92 VP.n22 B 0.23169f
C93 VP.n23 B 1.43883f
C94 VP.n24 B 1.47715f
C95 VP.t9 B 0.416809f
C96 VP.n25 B 0.23169f
C97 VP.t6 B 0.353222f
C98 VP.n26 B 0.168107f
C99 VP.n27 B 0.054003f
C100 VP.n28 B 0.054298f
C101 VP.n29 B 0.040692f
C102 VP.n30 B 0.040692f
C103 VP.n31 B 0.035935f
C104 VP.n32 B 0.057849f
C105 VP.n33 B 0.168107f
C106 VP.n34 B 0.057849f
C107 VP.n35 B 0.040692f
C108 VP.n36 B 0.040692f
C109 VP.n37 B 0.040692f
C110 VP.n38 B 0.052194f
C111 VP.n39 B 0.168107f
C112 VP.n40 B 0.054003f
C113 VP.t5 B 0.416809f
C114 VP.n41 B 0.23169f
C115 VP.n42 B 0.03811f
C116 VDD2.n0 B 0.034967f
C117 VDD2.n1 B 0.023847f
C118 VDD2.n2 B 0.012814f
C119 VDD2.n3 B 0.022716f
C120 VDD2.n4 B 0.021207f
C121 VDD2.t3 B 0.052957f
C122 VDD2.n5 B 0.096044f
C123 VDD2.n6 B 0.281842f
C124 VDD2.n7 B 0.012814f
C125 VDD2.n8 B 0.013568f
C126 VDD2.n9 B 0.030288f
C127 VDD2.n10 B 0.06813f
C128 VDD2.n11 B 0.013568f
C129 VDD2.n12 B 0.012814f
C130 VDD2.n13 B 0.051537f
C131 VDD2.n14 B 0.058006f
C132 VDD2.t8 B 0.063506f
C133 VDD2.t6 B 0.063506f
C134 VDD2.n15 B 0.471188f
C135 VDD2.n16 B 0.43369f
C136 VDD2.t4 B 0.063506f
C137 VDD2.t9 B 0.063506f
C138 VDD2.n17 B 0.474944f
C139 VDD2.n18 B 1.49014f
C140 VDD2.n19 B 0.034967f
C141 VDD2.n20 B 0.023847f
C142 VDD2.n21 B 0.012814f
C143 VDD2.n22 B 0.022716f
C144 VDD2.n23 B 0.021207f
C145 VDD2.t1 B 0.052957f
C146 VDD2.n24 B 0.096044f
C147 VDD2.n25 B 0.281842f
C148 VDD2.n26 B 0.012814f
C149 VDD2.n27 B 0.013568f
C150 VDD2.n28 B 0.030288f
C151 VDD2.n29 B 0.06813f
C152 VDD2.n30 B 0.013568f
C153 VDD2.n31 B 0.012814f
C154 VDD2.n32 B 0.051537f
C155 VDD2.n33 B 0.054767f
C156 VDD2.n34 B 1.51379f
C157 VDD2.t0 B 0.063506f
C158 VDD2.t7 B 0.063506f
C159 VDD2.n35 B 0.47119f
C160 VDD2.n36 B 0.31001f
C161 VDD2.t5 B 0.063506f
C162 VDD2.t2 B 0.063506f
C163 VDD2.n37 B 0.474923f
C164 VTAIL.t14 B 0.078814f
C165 VTAIL.t16 B 0.078814f
C166 VTAIL.n0 B 0.519557f
C167 VTAIL.n1 B 0.454536f
C168 VTAIL.n2 B 0.043396f
C169 VTAIL.n3 B 0.029595f
C170 VTAIL.n4 B 0.015903f
C171 VTAIL.n5 B 0.028192f
C172 VTAIL.n6 B 0.026319f
C173 VTAIL.t2 B 0.065723f
C174 VTAIL.n7 B 0.119196f
C175 VTAIL.n8 B 0.349782f
C176 VTAIL.n9 B 0.015903f
C177 VTAIL.n10 B 0.016839f
C178 VTAIL.n11 B 0.037589f
C179 VTAIL.n12 B 0.084553f
C180 VTAIL.n13 B 0.016839f
C181 VTAIL.n14 B 0.015903f
C182 VTAIL.n15 B 0.063961f
C183 VTAIL.n16 B 0.047496f
C184 VTAIL.n17 B 0.234048f
C185 VTAIL.t1 B 0.078814f
C186 VTAIL.t7 B 0.078814f
C187 VTAIL.n18 B 0.519557f
C188 VTAIL.n19 B 0.48742f
C189 VTAIL.t6 B 0.078814f
C190 VTAIL.t0 B 0.078814f
C191 VTAIL.n20 B 0.519557f
C192 VTAIL.n21 B 1.27746f
C193 VTAIL.t10 B 0.078814f
C194 VTAIL.t13 B 0.078814f
C195 VTAIL.n22 B 0.519559f
C196 VTAIL.n23 B 1.27746f
C197 VTAIL.t19 B 0.078814f
C198 VTAIL.t15 B 0.078814f
C199 VTAIL.n24 B 0.519559f
C200 VTAIL.n25 B 0.487417f
C201 VTAIL.n26 B 0.043396f
C202 VTAIL.n27 B 0.029595f
C203 VTAIL.n28 B 0.015903f
C204 VTAIL.n29 B 0.028192f
C205 VTAIL.n30 B 0.026319f
C206 VTAIL.t12 B 0.065723f
C207 VTAIL.n31 B 0.119196f
C208 VTAIL.n32 B 0.349782f
C209 VTAIL.n33 B 0.015903f
C210 VTAIL.n34 B 0.016839f
C211 VTAIL.n35 B 0.037589f
C212 VTAIL.n36 B 0.084553f
C213 VTAIL.n37 B 0.016839f
C214 VTAIL.n38 B 0.015903f
C215 VTAIL.n39 B 0.063961f
C216 VTAIL.n40 B 0.047496f
C217 VTAIL.n41 B 0.234048f
C218 VTAIL.t9 B 0.078814f
C219 VTAIL.t5 B 0.078814f
C220 VTAIL.n42 B 0.519559f
C221 VTAIL.n43 B 0.47673f
C222 VTAIL.t3 B 0.078814f
C223 VTAIL.t4 B 0.078814f
C224 VTAIL.n44 B 0.519559f
C225 VTAIL.n45 B 0.487417f
C226 VTAIL.n46 B 0.043396f
C227 VTAIL.n47 B 0.029595f
C228 VTAIL.n48 B 0.015903f
C229 VTAIL.n49 B 0.028192f
C230 VTAIL.n50 B 0.026319f
C231 VTAIL.t8 B 0.065723f
C232 VTAIL.n51 B 0.119196f
C233 VTAIL.n52 B 0.349782f
C234 VTAIL.n53 B 0.015903f
C235 VTAIL.n54 B 0.016839f
C236 VTAIL.n55 B 0.037589f
C237 VTAIL.n56 B 0.084553f
C238 VTAIL.n57 B 0.016839f
C239 VTAIL.n58 B 0.015903f
C240 VTAIL.n59 B 0.063961f
C241 VTAIL.n60 B 0.047496f
C242 VTAIL.n61 B 0.923797f
C243 VTAIL.n62 B 0.043396f
C244 VTAIL.n63 B 0.029595f
C245 VTAIL.n64 B 0.015903f
C246 VTAIL.n65 B 0.028192f
C247 VTAIL.n66 B 0.026319f
C248 VTAIL.t18 B 0.065723f
C249 VTAIL.n67 B 0.119196f
C250 VTAIL.n68 B 0.349782f
C251 VTAIL.n69 B 0.015903f
C252 VTAIL.n70 B 0.016839f
C253 VTAIL.n71 B 0.037589f
C254 VTAIL.n72 B 0.084553f
C255 VTAIL.n73 B 0.016839f
C256 VTAIL.n74 B 0.015903f
C257 VTAIL.n75 B 0.063961f
C258 VTAIL.n76 B 0.047496f
C259 VTAIL.n77 B 0.923797f
C260 VTAIL.t11 B 0.078814f
C261 VTAIL.t17 B 0.078814f
C262 VTAIL.n78 B 0.519557f
C263 VTAIL.n79 B 0.398634f
C264 VN.n0 B 0.05295f
C265 VN.t5 B 0.34445f
C266 VN.n1 B 0.035043f
C267 VN.n2 B 0.039681f
C268 VN.t3 B 0.34445f
C269 VN.n3 B 0.050897f
C270 VN.t6 B 0.431378f
C271 VN.t1 B 0.34445f
C272 VN.n4 B 0.19547f
C273 VN.n5 B 0.222963f
C274 VN.n6 B 0.168181f
C275 VN.n7 B 0.039681f
C276 VN.n8 B 0.035043f
C277 VN.n9 B 0.056413f
C278 VN.n10 B 0.163933f
C279 VN.n11 B 0.056413f
C280 VN.n12 B 0.039681f
C281 VN.n13 B 0.039681f
C282 VN.n14 B 0.039681f
C283 VN.n15 B 0.050897f
C284 VN.n16 B 0.163933f
C285 VN.n17 B 0.052662f
C286 VN.t0 B 0.406459f
C287 VN.n18 B 0.225937f
C288 VN.n19 B 0.037163f
C289 VN.n20 B 0.05295f
C290 VN.t9 B 0.34445f
C291 VN.n21 B 0.035043f
C292 VN.n22 B 0.039681f
C293 VN.t2 B 0.34445f
C294 VN.n23 B 0.050897f
C295 VN.t7 B 0.431378f
C296 VN.t4 B 0.34445f
C297 VN.n24 B 0.19547f
C298 VN.n25 B 0.222963f
C299 VN.n26 B 0.168181f
C300 VN.n27 B 0.039681f
C301 VN.n28 B 0.035043f
C302 VN.n29 B 0.056413f
C303 VN.n30 B 0.163933f
C304 VN.n31 B 0.056413f
C305 VN.n32 B 0.039681f
C306 VN.n33 B 0.039681f
C307 VN.n34 B 0.039681f
C308 VN.n35 B 0.050897f
C309 VN.n36 B 0.163933f
C310 VN.n37 B 0.052662f
C311 VN.t8 B 0.406459f
C312 VN.n38 B 0.225937f
C313 VN.n39 B 1.42575f
.ends

