* NGSPICE file created from diff_pair_sample_0931.ext - technology: sky130A

.subckt diff_pair_sample_0931 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=0 ps=0 w=16.08 l=2.27
X1 VDD1.t5 VP.t0 VTAIL.t6 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=6.2712 ps=32.94 w=16.08 l=2.27
X2 VTAIL.t11 VP.t1 VDD1.t4 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=2.6532 ps=16.41 w=16.08 l=2.27
X3 B.t8 B.t6 B.t7 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=0 ps=0 w=16.08 l=2.27
X4 B.t5 B.t3 B.t4 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=0 ps=0 w=16.08 l=2.27
X5 VDD2.t5 VN.t0 VTAIL.t0 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=6.2712 ps=32.94 w=16.08 l=2.27
X6 VTAIL.t5 VN.t1 VDD2.t4 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=2.6532 ps=16.41 w=16.08 l=2.27
X7 VDD2.t3 VN.t2 VTAIL.t3 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=2.6532 ps=16.41 w=16.08 l=2.27
X8 VDD1.t3 VP.t2 VTAIL.t10 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=2.6532 ps=16.41 w=16.08 l=2.27
X9 VDD2.t2 VN.t3 VTAIL.t2 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=2.6532 ps=16.41 w=16.08 l=2.27
X10 VDD1.t2 VP.t3 VTAIL.t7 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=6.2712 ps=32.94 w=16.08 l=2.27
X11 VTAIL.t8 VP.t4 VDD1.t1 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=2.6532 ps=16.41 w=16.08 l=2.27
X12 B.t2 B.t0 B.t1 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=0 ps=0 w=16.08 l=2.27
X13 VTAIL.t1 VN.t4 VDD2.t1 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=2.6532 ps=16.41 w=16.08 l=2.27
X14 VDD2.t0 VN.t5 VTAIL.t4 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=2.6532 pd=16.41 as=6.2712 ps=32.94 w=16.08 l=2.27
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n3050_n4184# sky130_fd_pr__pfet_01v8 ad=6.2712 pd=32.94 as=2.6532 ps=16.41 w=16.08 l=2.27
R0 B.n436 B.n123 585
R1 B.n435 B.n434 585
R2 B.n433 B.n124 585
R3 B.n432 B.n431 585
R4 B.n430 B.n125 585
R5 B.n429 B.n428 585
R6 B.n427 B.n126 585
R7 B.n426 B.n425 585
R8 B.n424 B.n127 585
R9 B.n423 B.n422 585
R10 B.n421 B.n128 585
R11 B.n420 B.n419 585
R12 B.n418 B.n129 585
R13 B.n417 B.n416 585
R14 B.n415 B.n130 585
R15 B.n414 B.n413 585
R16 B.n412 B.n131 585
R17 B.n411 B.n410 585
R18 B.n409 B.n132 585
R19 B.n408 B.n407 585
R20 B.n406 B.n133 585
R21 B.n405 B.n404 585
R22 B.n403 B.n134 585
R23 B.n402 B.n401 585
R24 B.n400 B.n135 585
R25 B.n399 B.n398 585
R26 B.n397 B.n136 585
R27 B.n396 B.n395 585
R28 B.n394 B.n137 585
R29 B.n393 B.n392 585
R30 B.n391 B.n138 585
R31 B.n390 B.n389 585
R32 B.n388 B.n139 585
R33 B.n387 B.n386 585
R34 B.n385 B.n140 585
R35 B.n384 B.n383 585
R36 B.n382 B.n141 585
R37 B.n381 B.n380 585
R38 B.n379 B.n142 585
R39 B.n378 B.n377 585
R40 B.n376 B.n143 585
R41 B.n375 B.n374 585
R42 B.n373 B.n144 585
R43 B.n372 B.n371 585
R44 B.n370 B.n145 585
R45 B.n369 B.n368 585
R46 B.n367 B.n146 585
R47 B.n366 B.n365 585
R48 B.n364 B.n147 585
R49 B.n363 B.n362 585
R50 B.n361 B.n148 585
R51 B.n360 B.n359 585
R52 B.n358 B.n149 585
R53 B.n357 B.n356 585
R54 B.n355 B.n354 585
R55 B.n353 B.n153 585
R56 B.n352 B.n351 585
R57 B.n350 B.n154 585
R58 B.n349 B.n348 585
R59 B.n347 B.n155 585
R60 B.n346 B.n345 585
R61 B.n344 B.n156 585
R62 B.n343 B.n342 585
R63 B.n340 B.n157 585
R64 B.n339 B.n338 585
R65 B.n337 B.n160 585
R66 B.n336 B.n335 585
R67 B.n334 B.n161 585
R68 B.n333 B.n332 585
R69 B.n331 B.n162 585
R70 B.n330 B.n329 585
R71 B.n328 B.n163 585
R72 B.n327 B.n326 585
R73 B.n325 B.n164 585
R74 B.n324 B.n323 585
R75 B.n322 B.n165 585
R76 B.n321 B.n320 585
R77 B.n319 B.n166 585
R78 B.n318 B.n317 585
R79 B.n316 B.n167 585
R80 B.n315 B.n314 585
R81 B.n313 B.n168 585
R82 B.n312 B.n311 585
R83 B.n310 B.n169 585
R84 B.n309 B.n308 585
R85 B.n307 B.n170 585
R86 B.n306 B.n305 585
R87 B.n304 B.n171 585
R88 B.n303 B.n302 585
R89 B.n301 B.n172 585
R90 B.n300 B.n299 585
R91 B.n298 B.n173 585
R92 B.n297 B.n296 585
R93 B.n295 B.n174 585
R94 B.n294 B.n293 585
R95 B.n292 B.n175 585
R96 B.n291 B.n290 585
R97 B.n289 B.n176 585
R98 B.n288 B.n287 585
R99 B.n286 B.n177 585
R100 B.n285 B.n284 585
R101 B.n283 B.n178 585
R102 B.n282 B.n281 585
R103 B.n280 B.n179 585
R104 B.n279 B.n278 585
R105 B.n277 B.n180 585
R106 B.n276 B.n275 585
R107 B.n274 B.n181 585
R108 B.n273 B.n272 585
R109 B.n271 B.n182 585
R110 B.n270 B.n269 585
R111 B.n268 B.n183 585
R112 B.n267 B.n266 585
R113 B.n265 B.n184 585
R114 B.n264 B.n263 585
R115 B.n262 B.n185 585
R116 B.n261 B.n260 585
R117 B.n438 B.n437 585
R118 B.n439 B.n122 585
R119 B.n441 B.n440 585
R120 B.n442 B.n121 585
R121 B.n444 B.n443 585
R122 B.n445 B.n120 585
R123 B.n447 B.n446 585
R124 B.n448 B.n119 585
R125 B.n450 B.n449 585
R126 B.n451 B.n118 585
R127 B.n453 B.n452 585
R128 B.n454 B.n117 585
R129 B.n456 B.n455 585
R130 B.n457 B.n116 585
R131 B.n459 B.n458 585
R132 B.n460 B.n115 585
R133 B.n462 B.n461 585
R134 B.n463 B.n114 585
R135 B.n465 B.n464 585
R136 B.n466 B.n113 585
R137 B.n468 B.n467 585
R138 B.n469 B.n112 585
R139 B.n471 B.n470 585
R140 B.n472 B.n111 585
R141 B.n474 B.n473 585
R142 B.n475 B.n110 585
R143 B.n477 B.n476 585
R144 B.n478 B.n109 585
R145 B.n480 B.n479 585
R146 B.n481 B.n108 585
R147 B.n483 B.n482 585
R148 B.n484 B.n107 585
R149 B.n486 B.n485 585
R150 B.n487 B.n106 585
R151 B.n489 B.n488 585
R152 B.n490 B.n105 585
R153 B.n492 B.n491 585
R154 B.n493 B.n104 585
R155 B.n495 B.n494 585
R156 B.n496 B.n103 585
R157 B.n498 B.n497 585
R158 B.n499 B.n102 585
R159 B.n501 B.n500 585
R160 B.n502 B.n101 585
R161 B.n504 B.n503 585
R162 B.n505 B.n100 585
R163 B.n507 B.n506 585
R164 B.n508 B.n99 585
R165 B.n510 B.n509 585
R166 B.n511 B.n98 585
R167 B.n513 B.n512 585
R168 B.n514 B.n97 585
R169 B.n516 B.n515 585
R170 B.n517 B.n96 585
R171 B.n519 B.n518 585
R172 B.n520 B.n95 585
R173 B.n522 B.n521 585
R174 B.n523 B.n94 585
R175 B.n525 B.n524 585
R176 B.n526 B.n93 585
R177 B.n528 B.n527 585
R178 B.n529 B.n92 585
R179 B.n531 B.n530 585
R180 B.n532 B.n91 585
R181 B.n534 B.n533 585
R182 B.n535 B.n90 585
R183 B.n537 B.n536 585
R184 B.n538 B.n89 585
R185 B.n540 B.n539 585
R186 B.n541 B.n88 585
R187 B.n543 B.n542 585
R188 B.n544 B.n87 585
R189 B.n546 B.n545 585
R190 B.n547 B.n86 585
R191 B.n549 B.n548 585
R192 B.n550 B.n85 585
R193 B.n552 B.n551 585
R194 B.n553 B.n84 585
R195 B.n730 B.n21 585
R196 B.n729 B.n728 585
R197 B.n727 B.n22 585
R198 B.n726 B.n725 585
R199 B.n724 B.n23 585
R200 B.n723 B.n722 585
R201 B.n721 B.n24 585
R202 B.n720 B.n719 585
R203 B.n718 B.n25 585
R204 B.n717 B.n716 585
R205 B.n715 B.n26 585
R206 B.n714 B.n713 585
R207 B.n712 B.n27 585
R208 B.n711 B.n710 585
R209 B.n709 B.n28 585
R210 B.n708 B.n707 585
R211 B.n706 B.n29 585
R212 B.n705 B.n704 585
R213 B.n703 B.n30 585
R214 B.n702 B.n701 585
R215 B.n700 B.n31 585
R216 B.n699 B.n698 585
R217 B.n697 B.n32 585
R218 B.n696 B.n695 585
R219 B.n694 B.n33 585
R220 B.n693 B.n692 585
R221 B.n691 B.n34 585
R222 B.n690 B.n689 585
R223 B.n688 B.n35 585
R224 B.n687 B.n686 585
R225 B.n685 B.n36 585
R226 B.n684 B.n683 585
R227 B.n682 B.n37 585
R228 B.n681 B.n680 585
R229 B.n679 B.n38 585
R230 B.n678 B.n677 585
R231 B.n676 B.n39 585
R232 B.n675 B.n674 585
R233 B.n673 B.n40 585
R234 B.n672 B.n671 585
R235 B.n670 B.n41 585
R236 B.n669 B.n668 585
R237 B.n667 B.n42 585
R238 B.n666 B.n665 585
R239 B.n664 B.n43 585
R240 B.n663 B.n662 585
R241 B.n661 B.n44 585
R242 B.n660 B.n659 585
R243 B.n658 B.n45 585
R244 B.n657 B.n656 585
R245 B.n655 B.n46 585
R246 B.n654 B.n653 585
R247 B.n652 B.n47 585
R248 B.n651 B.n650 585
R249 B.n649 B.n648 585
R250 B.n647 B.n51 585
R251 B.n646 B.n645 585
R252 B.n644 B.n52 585
R253 B.n643 B.n642 585
R254 B.n641 B.n53 585
R255 B.n640 B.n639 585
R256 B.n638 B.n54 585
R257 B.n637 B.n636 585
R258 B.n634 B.n55 585
R259 B.n633 B.n632 585
R260 B.n631 B.n58 585
R261 B.n630 B.n629 585
R262 B.n628 B.n59 585
R263 B.n627 B.n626 585
R264 B.n625 B.n60 585
R265 B.n624 B.n623 585
R266 B.n622 B.n61 585
R267 B.n621 B.n620 585
R268 B.n619 B.n62 585
R269 B.n618 B.n617 585
R270 B.n616 B.n63 585
R271 B.n615 B.n614 585
R272 B.n613 B.n64 585
R273 B.n612 B.n611 585
R274 B.n610 B.n65 585
R275 B.n609 B.n608 585
R276 B.n607 B.n66 585
R277 B.n606 B.n605 585
R278 B.n604 B.n67 585
R279 B.n603 B.n602 585
R280 B.n601 B.n68 585
R281 B.n600 B.n599 585
R282 B.n598 B.n69 585
R283 B.n597 B.n596 585
R284 B.n595 B.n70 585
R285 B.n594 B.n593 585
R286 B.n592 B.n71 585
R287 B.n591 B.n590 585
R288 B.n589 B.n72 585
R289 B.n588 B.n587 585
R290 B.n586 B.n73 585
R291 B.n585 B.n584 585
R292 B.n583 B.n74 585
R293 B.n582 B.n581 585
R294 B.n580 B.n75 585
R295 B.n579 B.n578 585
R296 B.n577 B.n76 585
R297 B.n576 B.n575 585
R298 B.n574 B.n77 585
R299 B.n573 B.n572 585
R300 B.n571 B.n78 585
R301 B.n570 B.n569 585
R302 B.n568 B.n79 585
R303 B.n567 B.n566 585
R304 B.n565 B.n80 585
R305 B.n564 B.n563 585
R306 B.n562 B.n81 585
R307 B.n561 B.n560 585
R308 B.n559 B.n82 585
R309 B.n558 B.n557 585
R310 B.n556 B.n83 585
R311 B.n555 B.n554 585
R312 B.n732 B.n731 585
R313 B.n733 B.n20 585
R314 B.n735 B.n734 585
R315 B.n736 B.n19 585
R316 B.n738 B.n737 585
R317 B.n739 B.n18 585
R318 B.n741 B.n740 585
R319 B.n742 B.n17 585
R320 B.n744 B.n743 585
R321 B.n745 B.n16 585
R322 B.n747 B.n746 585
R323 B.n748 B.n15 585
R324 B.n750 B.n749 585
R325 B.n751 B.n14 585
R326 B.n753 B.n752 585
R327 B.n754 B.n13 585
R328 B.n756 B.n755 585
R329 B.n757 B.n12 585
R330 B.n759 B.n758 585
R331 B.n760 B.n11 585
R332 B.n762 B.n761 585
R333 B.n763 B.n10 585
R334 B.n765 B.n764 585
R335 B.n766 B.n9 585
R336 B.n768 B.n767 585
R337 B.n769 B.n8 585
R338 B.n771 B.n770 585
R339 B.n772 B.n7 585
R340 B.n774 B.n773 585
R341 B.n775 B.n6 585
R342 B.n777 B.n776 585
R343 B.n778 B.n5 585
R344 B.n780 B.n779 585
R345 B.n781 B.n4 585
R346 B.n783 B.n782 585
R347 B.n784 B.n3 585
R348 B.n786 B.n785 585
R349 B.n787 B.n0 585
R350 B.n2 B.n1 585
R351 B.n205 B.n204 585
R352 B.n207 B.n206 585
R353 B.n208 B.n203 585
R354 B.n210 B.n209 585
R355 B.n211 B.n202 585
R356 B.n213 B.n212 585
R357 B.n214 B.n201 585
R358 B.n216 B.n215 585
R359 B.n217 B.n200 585
R360 B.n219 B.n218 585
R361 B.n220 B.n199 585
R362 B.n222 B.n221 585
R363 B.n223 B.n198 585
R364 B.n225 B.n224 585
R365 B.n226 B.n197 585
R366 B.n228 B.n227 585
R367 B.n229 B.n196 585
R368 B.n231 B.n230 585
R369 B.n232 B.n195 585
R370 B.n234 B.n233 585
R371 B.n235 B.n194 585
R372 B.n237 B.n236 585
R373 B.n238 B.n193 585
R374 B.n240 B.n239 585
R375 B.n241 B.n192 585
R376 B.n243 B.n242 585
R377 B.n244 B.n191 585
R378 B.n246 B.n245 585
R379 B.n247 B.n190 585
R380 B.n249 B.n248 585
R381 B.n250 B.n189 585
R382 B.n252 B.n251 585
R383 B.n253 B.n188 585
R384 B.n255 B.n254 585
R385 B.n256 B.n187 585
R386 B.n258 B.n257 585
R387 B.n259 B.n186 585
R388 B.n260 B.n259 516.524
R389 B.n438 B.n123 516.524
R390 B.n554 B.n553 516.524
R391 B.n732 B.n21 516.524
R392 B.n150 B.t1 499.44
R393 B.n56 B.t5 499.44
R394 B.n158 B.t10 499.44
R395 B.n48 B.t8 499.44
R396 B.n151 B.t2 449.017
R397 B.n57 B.t4 449.017
R398 B.n159 B.t11 449.017
R399 B.n49 B.t7 449.017
R400 B.n158 B.t9 378.205
R401 B.n150 B.t0 378.205
R402 B.n56 B.t3 378.205
R403 B.n48 B.t6 378.205
R404 B.n789 B.n788 256.663
R405 B.n788 B.n787 235.042
R406 B.n788 B.n2 235.042
R407 B.n260 B.n185 163.367
R408 B.n264 B.n185 163.367
R409 B.n265 B.n264 163.367
R410 B.n266 B.n265 163.367
R411 B.n266 B.n183 163.367
R412 B.n270 B.n183 163.367
R413 B.n271 B.n270 163.367
R414 B.n272 B.n271 163.367
R415 B.n272 B.n181 163.367
R416 B.n276 B.n181 163.367
R417 B.n277 B.n276 163.367
R418 B.n278 B.n277 163.367
R419 B.n278 B.n179 163.367
R420 B.n282 B.n179 163.367
R421 B.n283 B.n282 163.367
R422 B.n284 B.n283 163.367
R423 B.n284 B.n177 163.367
R424 B.n288 B.n177 163.367
R425 B.n289 B.n288 163.367
R426 B.n290 B.n289 163.367
R427 B.n290 B.n175 163.367
R428 B.n294 B.n175 163.367
R429 B.n295 B.n294 163.367
R430 B.n296 B.n295 163.367
R431 B.n296 B.n173 163.367
R432 B.n300 B.n173 163.367
R433 B.n301 B.n300 163.367
R434 B.n302 B.n301 163.367
R435 B.n302 B.n171 163.367
R436 B.n306 B.n171 163.367
R437 B.n307 B.n306 163.367
R438 B.n308 B.n307 163.367
R439 B.n308 B.n169 163.367
R440 B.n312 B.n169 163.367
R441 B.n313 B.n312 163.367
R442 B.n314 B.n313 163.367
R443 B.n314 B.n167 163.367
R444 B.n318 B.n167 163.367
R445 B.n319 B.n318 163.367
R446 B.n320 B.n319 163.367
R447 B.n320 B.n165 163.367
R448 B.n324 B.n165 163.367
R449 B.n325 B.n324 163.367
R450 B.n326 B.n325 163.367
R451 B.n326 B.n163 163.367
R452 B.n330 B.n163 163.367
R453 B.n331 B.n330 163.367
R454 B.n332 B.n331 163.367
R455 B.n332 B.n161 163.367
R456 B.n336 B.n161 163.367
R457 B.n337 B.n336 163.367
R458 B.n338 B.n337 163.367
R459 B.n338 B.n157 163.367
R460 B.n343 B.n157 163.367
R461 B.n344 B.n343 163.367
R462 B.n345 B.n344 163.367
R463 B.n345 B.n155 163.367
R464 B.n349 B.n155 163.367
R465 B.n350 B.n349 163.367
R466 B.n351 B.n350 163.367
R467 B.n351 B.n153 163.367
R468 B.n355 B.n153 163.367
R469 B.n356 B.n355 163.367
R470 B.n356 B.n149 163.367
R471 B.n360 B.n149 163.367
R472 B.n361 B.n360 163.367
R473 B.n362 B.n361 163.367
R474 B.n362 B.n147 163.367
R475 B.n366 B.n147 163.367
R476 B.n367 B.n366 163.367
R477 B.n368 B.n367 163.367
R478 B.n368 B.n145 163.367
R479 B.n372 B.n145 163.367
R480 B.n373 B.n372 163.367
R481 B.n374 B.n373 163.367
R482 B.n374 B.n143 163.367
R483 B.n378 B.n143 163.367
R484 B.n379 B.n378 163.367
R485 B.n380 B.n379 163.367
R486 B.n380 B.n141 163.367
R487 B.n384 B.n141 163.367
R488 B.n385 B.n384 163.367
R489 B.n386 B.n385 163.367
R490 B.n386 B.n139 163.367
R491 B.n390 B.n139 163.367
R492 B.n391 B.n390 163.367
R493 B.n392 B.n391 163.367
R494 B.n392 B.n137 163.367
R495 B.n396 B.n137 163.367
R496 B.n397 B.n396 163.367
R497 B.n398 B.n397 163.367
R498 B.n398 B.n135 163.367
R499 B.n402 B.n135 163.367
R500 B.n403 B.n402 163.367
R501 B.n404 B.n403 163.367
R502 B.n404 B.n133 163.367
R503 B.n408 B.n133 163.367
R504 B.n409 B.n408 163.367
R505 B.n410 B.n409 163.367
R506 B.n410 B.n131 163.367
R507 B.n414 B.n131 163.367
R508 B.n415 B.n414 163.367
R509 B.n416 B.n415 163.367
R510 B.n416 B.n129 163.367
R511 B.n420 B.n129 163.367
R512 B.n421 B.n420 163.367
R513 B.n422 B.n421 163.367
R514 B.n422 B.n127 163.367
R515 B.n426 B.n127 163.367
R516 B.n427 B.n426 163.367
R517 B.n428 B.n427 163.367
R518 B.n428 B.n125 163.367
R519 B.n432 B.n125 163.367
R520 B.n433 B.n432 163.367
R521 B.n434 B.n433 163.367
R522 B.n434 B.n123 163.367
R523 B.n553 B.n552 163.367
R524 B.n552 B.n85 163.367
R525 B.n548 B.n85 163.367
R526 B.n548 B.n547 163.367
R527 B.n547 B.n546 163.367
R528 B.n546 B.n87 163.367
R529 B.n542 B.n87 163.367
R530 B.n542 B.n541 163.367
R531 B.n541 B.n540 163.367
R532 B.n540 B.n89 163.367
R533 B.n536 B.n89 163.367
R534 B.n536 B.n535 163.367
R535 B.n535 B.n534 163.367
R536 B.n534 B.n91 163.367
R537 B.n530 B.n91 163.367
R538 B.n530 B.n529 163.367
R539 B.n529 B.n528 163.367
R540 B.n528 B.n93 163.367
R541 B.n524 B.n93 163.367
R542 B.n524 B.n523 163.367
R543 B.n523 B.n522 163.367
R544 B.n522 B.n95 163.367
R545 B.n518 B.n95 163.367
R546 B.n518 B.n517 163.367
R547 B.n517 B.n516 163.367
R548 B.n516 B.n97 163.367
R549 B.n512 B.n97 163.367
R550 B.n512 B.n511 163.367
R551 B.n511 B.n510 163.367
R552 B.n510 B.n99 163.367
R553 B.n506 B.n99 163.367
R554 B.n506 B.n505 163.367
R555 B.n505 B.n504 163.367
R556 B.n504 B.n101 163.367
R557 B.n500 B.n101 163.367
R558 B.n500 B.n499 163.367
R559 B.n499 B.n498 163.367
R560 B.n498 B.n103 163.367
R561 B.n494 B.n103 163.367
R562 B.n494 B.n493 163.367
R563 B.n493 B.n492 163.367
R564 B.n492 B.n105 163.367
R565 B.n488 B.n105 163.367
R566 B.n488 B.n487 163.367
R567 B.n487 B.n486 163.367
R568 B.n486 B.n107 163.367
R569 B.n482 B.n107 163.367
R570 B.n482 B.n481 163.367
R571 B.n481 B.n480 163.367
R572 B.n480 B.n109 163.367
R573 B.n476 B.n109 163.367
R574 B.n476 B.n475 163.367
R575 B.n475 B.n474 163.367
R576 B.n474 B.n111 163.367
R577 B.n470 B.n111 163.367
R578 B.n470 B.n469 163.367
R579 B.n469 B.n468 163.367
R580 B.n468 B.n113 163.367
R581 B.n464 B.n113 163.367
R582 B.n464 B.n463 163.367
R583 B.n463 B.n462 163.367
R584 B.n462 B.n115 163.367
R585 B.n458 B.n115 163.367
R586 B.n458 B.n457 163.367
R587 B.n457 B.n456 163.367
R588 B.n456 B.n117 163.367
R589 B.n452 B.n117 163.367
R590 B.n452 B.n451 163.367
R591 B.n451 B.n450 163.367
R592 B.n450 B.n119 163.367
R593 B.n446 B.n119 163.367
R594 B.n446 B.n445 163.367
R595 B.n445 B.n444 163.367
R596 B.n444 B.n121 163.367
R597 B.n440 B.n121 163.367
R598 B.n440 B.n439 163.367
R599 B.n439 B.n438 163.367
R600 B.n728 B.n21 163.367
R601 B.n728 B.n727 163.367
R602 B.n727 B.n726 163.367
R603 B.n726 B.n23 163.367
R604 B.n722 B.n23 163.367
R605 B.n722 B.n721 163.367
R606 B.n721 B.n720 163.367
R607 B.n720 B.n25 163.367
R608 B.n716 B.n25 163.367
R609 B.n716 B.n715 163.367
R610 B.n715 B.n714 163.367
R611 B.n714 B.n27 163.367
R612 B.n710 B.n27 163.367
R613 B.n710 B.n709 163.367
R614 B.n709 B.n708 163.367
R615 B.n708 B.n29 163.367
R616 B.n704 B.n29 163.367
R617 B.n704 B.n703 163.367
R618 B.n703 B.n702 163.367
R619 B.n702 B.n31 163.367
R620 B.n698 B.n31 163.367
R621 B.n698 B.n697 163.367
R622 B.n697 B.n696 163.367
R623 B.n696 B.n33 163.367
R624 B.n692 B.n33 163.367
R625 B.n692 B.n691 163.367
R626 B.n691 B.n690 163.367
R627 B.n690 B.n35 163.367
R628 B.n686 B.n35 163.367
R629 B.n686 B.n685 163.367
R630 B.n685 B.n684 163.367
R631 B.n684 B.n37 163.367
R632 B.n680 B.n37 163.367
R633 B.n680 B.n679 163.367
R634 B.n679 B.n678 163.367
R635 B.n678 B.n39 163.367
R636 B.n674 B.n39 163.367
R637 B.n674 B.n673 163.367
R638 B.n673 B.n672 163.367
R639 B.n672 B.n41 163.367
R640 B.n668 B.n41 163.367
R641 B.n668 B.n667 163.367
R642 B.n667 B.n666 163.367
R643 B.n666 B.n43 163.367
R644 B.n662 B.n43 163.367
R645 B.n662 B.n661 163.367
R646 B.n661 B.n660 163.367
R647 B.n660 B.n45 163.367
R648 B.n656 B.n45 163.367
R649 B.n656 B.n655 163.367
R650 B.n655 B.n654 163.367
R651 B.n654 B.n47 163.367
R652 B.n650 B.n47 163.367
R653 B.n650 B.n649 163.367
R654 B.n649 B.n51 163.367
R655 B.n645 B.n51 163.367
R656 B.n645 B.n644 163.367
R657 B.n644 B.n643 163.367
R658 B.n643 B.n53 163.367
R659 B.n639 B.n53 163.367
R660 B.n639 B.n638 163.367
R661 B.n638 B.n637 163.367
R662 B.n637 B.n55 163.367
R663 B.n632 B.n55 163.367
R664 B.n632 B.n631 163.367
R665 B.n631 B.n630 163.367
R666 B.n630 B.n59 163.367
R667 B.n626 B.n59 163.367
R668 B.n626 B.n625 163.367
R669 B.n625 B.n624 163.367
R670 B.n624 B.n61 163.367
R671 B.n620 B.n61 163.367
R672 B.n620 B.n619 163.367
R673 B.n619 B.n618 163.367
R674 B.n618 B.n63 163.367
R675 B.n614 B.n63 163.367
R676 B.n614 B.n613 163.367
R677 B.n613 B.n612 163.367
R678 B.n612 B.n65 163.367
R679 B.n608 B.n65 163.367
R680 B.n608 B.n607 163.367
R681 B.n607 B.n606 163.367
R682 B.n606 B.n67 163.367
R683 B.n602 B.n67 163.367
R684 B.n602 B.n601 163.367
R685 B.n601 B.n600 163.367
R686 B.n600 B.n69 163.367
R687 B.n596 B.n69 163.367
R688 B.n596 B.n595 163.367
R689 B.n595 B.n594 163.367
R690 B.n594 B.n71 163.367
R691 B.n590 B.n71 163.367
R692 B.n590 B.n589 163.367
R693 B.n589 B.n588 163.367
R694 B.n588 B.n73 163.367
R695 B.n584 B.n73 163.367
R696 B.n584 B.n583 163.367
R697 B.n583 B.n582 163.367
R698 B.n582 B.n75 163.367
R699 B.n578 B.n75 163.367
R700 B.n578 B.n577 163.367
R701 B.n577 B.n576 163.367
R702 B.n576 B.n77 163.367
R703 B.n572 B.n77 163.367
R704 B.n572 B.n571 163.367
R705 B.n571 B.n570 163.367
R706 B.n570 B.n79 163.367
R707 B.n566 B.n79 163.367
R708 B.n566 B.n565 163.367
R709 B.n565 B.n564 163.367
R710 B.n564 B.n81 163.367
R711 B.n560 B.n81 163.367
R712 B.n560 B.n559 163.367
R713 B.n559 B.n558 163.367
R714 B.n558 B.n83 163.367
R715 B.n554 B.n83 163.367
R716 B.n733 B.n732 163.367
R717 B.n734 B.n733 163.367
R718 B.n734 B.n19 163.367
R719 B.n738 B.n19 163.367
R720 B.n739 B.n738 163.367
R721 B.n740 B.n739 163.367
R722 B.n740 B.n17 163.367
R723 B.n744 B.n17 163.367
R724 B.n745 B.n744 163.367
R725 B.n746 B.n745 163.367
R726 B.n746 B.n15 163.367
R727 B.n750 B.n15 163.367
R728 B.n751 B.n750 163.367
R729 B.n752 B.n751 163.367
R730 B.n752 B.n13 163.367
R731 B.n756 B.n13 163.367
R732 B.n757 B.n756 163.367
R733 B.n758 B.n757 163.367
R734 B.n758 B.n11 163.367
R735 B.n762 B.n11 163.367
R736 B.n763 B.n762 163.367
R737 B.n764 B.n763 163.367
R738 B.n764 B.n9 163.367
R739 B.n768 B.n9 163.367
R740 B.n769 B.n768 163.367
R741 B.n770 B.n769 163.367
R742 B.n770 B.n7 163.367
R743 B.n774 B.n7 163.367
R744 B.n775 B.n774 163.367
R745 B.n776 B.n775 163.367
R746 B.n776 B.n5 163.367
R747 B.n780 B.n5 163.367
R748 B.n781 B.n780 163.367
R749 B.n782 B.n781 163.367
R750 B.n782 B.n3 163.367
R751 B.n786 B.n3 163.367
R752 B.n787 B.n786 163.367
R753 B.n205 B.n2 163.367
R754 B.n206 B.n205 163.367
R755 B.n206 B.n203 163.367
R756 B.n210 B.n203 163.367
R757 B.n211 B.n210 163.367
R758 B.n212 B.n211 163.367
R759 B.n212 B.n201 163.367
R760 B.n216 B.n201 163.367
R761 B.n217 B.n216 163.367
R762 B.n218 B.n217 163.367
R763 B.n218 B.n199 163.367
R764 B.n222 B.n199 163.367
R765 B.n223 B.n222 163.367
R766 B.n224 B.n223 163.367
R767 B.n224 B.n197 163.367
R768 B.n228 B.n197 163.367
R769 B.n229 B.n228 163.367
R770 B.n230 B.n229 163.367
R771 B.n230 B.n195 163.367
R772 B.n234 B.n195 163.367
R773 B.n235 B.n234 163.367
R774 B.n236 B.n235 163.367
R775 B.n236 B.n193 163.367
R776 B.n240 B.n193 163.367
R777 B.n241 B.n240 163.367
R778 B.n242 B.n241 163.367
R779 B.n242 B.n191 163.367
R780 B.n246 B.n191 163.367
R781 B.n247 B.n246 163.367
R782 B.n248 B.n247 163.367
R783 B.n248 B.n189 163.367
R784 B.n252 B.n189 163.367
R785 B.n253 B.n252 163.367
R786 B.n254 B.n253 163.367
R787 B.n254 B.n187 163.367
R788 B.n258 B.n187 163.367
R789 B.n259 B.n258 163.367
R790 B.n341 B.n159 59.5399
R791 B.n152 B.n151 59.5399
R792 B.n635 B.n57 59.5399
R793 B.n50 B.n49 59.5399
R794 B.n159 B.n158 50.4247
R795 B.n151 B.n150 50.4247
R796 B.n57 B.n56 50.4247
R797 B.n49 B.n48 50.4247
R798 B.n731 B.n730 33.5615
R799 B.n555 B.n84 33.5615
R800 B.n437 B.n436 33.5615
R801 B.n261 B.n186 33.5615
R802 B B.n789 18.0485
R803 B.n731 B.n20 10.6151
R804 B.n735 B.n20 10.6151
R805 B.n736 B.n735 10.6151
R806 B.n737 B.n736 10.6151
R807 B.n737 B.n18 10.6151
R808 B.n741 B.n18 10.6151
R809 B.n742 B.n741 10.6151
R810 B.n743 B.n742 10.6151
R811 B.n743 B.n16 10.6151
R812 B.n747 B.n16 10.6151
R813 B.n748 B.n747 10.6151
R814 B.n749 B.n748 10.6151
R815 B.n749 B.n14 10.6151
R816 B.n753 B.n14 10.6151
R817 B.n754 B.n753 10.6151
R818 B.n755 B.n754 10.6151
R819 B.n755 B.n12 10.6151
R820 B.n759 B.n12 10.6151
R821 B.n760 B.n759 10.6151
R822 B.n761 B.n760 10.6151
R823 B.n761 B.n10 10.6151
R824 B.n765 B.n10 10.6151
R825 B.n766 B.n765 10.6151
R826 B.n767 B.n766 10.6151
R827 B.n767 B.n8 10.6151
R828 B.n771 B.n8 10.6151
R829 B.n772 B.n771 10.6151
R830 B.n773 B.n772 10.6151
R831 B.n773 B.n6 10.6151
R832 B.n777 B.n6 10.6151
R833 B.n778 B.n777 10.6151
R834 B.n779 B.n778 10.6151
R835 B.n779 B.n4 10.6151
R836 B.n783 B.n4 10.6151
R837 B.n784 B.n783 10.6151
R838 B.n785 B.n784 10.6151
R839 B.n785 B.n0 10.6151
R840 B.n730 B.n729 10.6151
R841 B.n729 B.n22 10.6151
R842 B.n725 B.n22 10.6151
R843 B.n725 B.n724 10.6151
R844 B.n724 B.n723 10.6151
R845 B.n723 B.n24 10.6151
R846 B.n719 B.n24 10.6151
R847 B.n719 B.n718 10.6151
R848 B.n718 B.n717 10.6151
R849 B.n717 B.n26 10.6151
R850 B.n713 B.n26 10.6151
R851 B.n713 B.n712 10.6151
R852 B.n712 B.n711 10.6151
R853 B.n711 B.n28 10.6151
R854 B.n707 B.n28 10.6151
R855 B.n707 B.n706 10.6151
R856 B.n706 B.n705 10.6151
R857 B.n705 B.n30 10.6151
R858 B.n701 B.n30 10.6151
R859 B.n701 B.n700 10.6151
R860 B.n700 B.n699 10.6151
R861 B.n699 B.n32 10.6151
R862 B.n695 B.n32 10.6151
R863 B.n695 B.n694 10.6151
R864 B.n694 B.n693 10.6151
R865 B.n693 B.n34 10.6151
R866 B.n689 B.n34 10.6151
R867 B.n689 B.n688 10.6151
R868 B.n688 B.n687 10.6151
R869 B.n687 B.n36 10.6151
R870 B.n683 B.n36 10.6151
R871 B.n683 B.n682 10.6151
R872 B.n682 B.n681 10.6151
R873 B.n681 B.n38 10.6151
R874 B.n677 B.n38 10.6151
R875 B.n677 B.n676 10.6151
R876 B.n676 B.n675 10.6151
R877 B.n675 B.n40 10.6151
R878 B.n671 B.n40 10.6151
R879 B.n671 B.n670 10.6151
R880 B.n670 B.n669 10.6151
R881 B.n669 B.n42 10.6151
R882 B.n665 B.n42 10.6151
R883 B.n665 B.n664 10.6151
R884 B.n664 B.n663 10.6151
R885 B.n663 B.n44 10.6151
R886 B.n659 B.n44 10.6151
R887 B.n659 B.n658 10.6151
R888 B.n658 B.n657 10.6151
R889 B.n657 B.n46 10.6151
R890 B.n653 B.n46 10.6151
R891 B.n653 B.n652 10.6151
R892 B.n652 B.n651 10.6151
R893 B.n648 B.n647 10.6151
R894 B.n647 B.n646 10.6151
R895 B.n646 B.n52 10.6151
R896 B.n642 B.n52 10.6151
R897 B.n642 B.n641 10.6151
R898 B.n641 B.n640 10.6151
R899 B.n640 B.n54 10.6151
R900 B.n636 B.n54 10.6151
R901 B.n634 B.n633 10.6151
R902 B.n633 B.n58 10.6151
R903 B.n629 B.n58 10.6151
R904 B.n629 B.n628 10.6151
R905 B.n628 B.n627 10.6151
R906 B.n627 B.n60 10.6151
R907 B.n623 B.n60 10.6151
R908 B.n623 B.n622 10.6151
R909 B.n622 B.n621 10.6151
R910 B.n621 B.n62 10.6151
R911 B.n617 B.n62 10.6151
R912 B.n617 B.n616 10.6151
R913 B.n616 B.n615 10.6151
R914 B.n615 B.n64 10.6151
R915 B.n611 B.n64 10.6151
R916 B.n611 B.n610 10.6151
R917 B.n610 B.n609 10.6151
R918 B.n609 B.n66 10.6151
R919 B.n605 B.n66 10.6151
R920 B.n605 B.n604 10.6151
R921 B.n604 B.n603 10.6151
R922 B.n603 B.n68 10.6151
R923 B.n599 B.n68 10.6151
R924 B.n599 B.n598 10.6151
R925 B.n598 B.n597 10.6151
R926 B.n597 B.n70 10.6151
R927 B.n593 B.n70 10.6151
R928 B.n593 B.n592 10.6151
R929 B.n592 B.n591 10.6151
R930 B.n591 B.n72 10.6151
R931 B.n587 B.n72 10.6151
R932 B.n587 B.n586 10.6151
R933 B.n586 B.n585 10.6151
R934 B.n585 B.n74 10.6151
R935 B.n581 B.n74 10.6151
R936 B.n581 B.n580 10.6151
R937 B.n580 B.n579 10.6151
R938 B.n579 B.n76 10.6151
R939 B.n575 B.n76 10.6151
R940 B.n575 B.n574 10.6151
R941 B.n574 B.n573 10.6151
R942 B.n573 B.n78 10.6151
R943 B.n569 B.n78 10.6151
R944 B.n569 B.n568 10.6151
R945 B.n568 B.n567 10.6151
R946 B.n567 B.n80 10.6151
R947 B.n563 B.n80 10.6151
R948 B.n563 B.n562 10.6151
R949 B.n562 B.n561 10.6151
R950 B.n561 B.n82 10.6151
R951 B.n557 B.n82 10.6151
R952 B.n557 B.n556 10.6151
R953 B.n556 B.n555 10.6151
R954 B.n551 B.n84 10.6151
R955 B.n551 B.n550 10.6151
R956 B.n550 B.n549 10.6151
R957 B.n549 B.n86 10.6151
R958 B.n545 B.n86 10.6151
R959 B.n545 B.n544 10.6151
R960 B.n544 B.n543 10.6151
R961 B.n543 B.n88 10.6151
R962 B.n539 B.n88 10.6151
R963 B.n539 B.n538 10.6151
R964 B.n538 B.n537 10.6151
R965 B.n537 B.n90 10.6151
R966 B.n533 B.n90 10.6151
R967 B.n533 B.n532 10.6151
R968 B.n532 B.n531 10.6151
R969 B.n531 B.n92 10.6151
R970 B.n527 B.n92 10.6151
R971 B.n527 B.n526 10.6151
R972 B.n526 B.n525 10.6151
R973 B.n525 B.n94 10.6151
R974 B.n521 B.n94 10.6151
R975 B.n521 B.n520 10.6151
R976 B.n520 B.n519 10.6151
R977 B.n519 B.n96 10.6151
R978 B.n515 B.n96 10.6151
R979 B.n515 B.n514 10.6151
R980 B.n514 B.n513 10.6151
R981 B.n513 B.n98 10.6151
R982 B.n509 B.n98 10.6151
R983 B.n509 B.n508 10.6151
R984 B.n508 B.n507 10.6151
R985 B.n507 B.n100 10.6151
R986 B.n503 B.n100 10.6151
R987 B.n503 B.n502 10.6151
R988 B.n502 B.n501 10.6151
R989 B.n501 B.n102 10.6151
R990 B.n497 B.n102 10.6151
R991 B.n497 B.n496 10.6151
R992 B.n496 B.n495 10.6151
R993 B.n495 B.n104 10.6151
R994 B.n491 B.n104 10.6151
R995 B.n491 B.n490 10.6151
R996 B.n490 B.n489 10.6151
R997 B.n489 B.n106 10.6151
R998 B.n485 B.n106 10.6151
R999 B.n485 B.n484 10.6151
R1000 B.n484 B.n483 10.6151
R1001 B.n483 B.n108 10.6151
R1002 B.n479 B.n108 10.6151
R1003 B.n479 B.n478 10.6151
R1004 B.n478 B.n477 10.6151
R1005 B.n477 B.n110 10.6151
R1006 B.n473 B.n110 10.6151
R1007 B.n473 B.n472 10.6151
R1008 B.n472 B.n471 10.6151
R1009 B.n471 B.n112 10.6151
R1010 B.n467 B.n112 10.6151
R1011 B.n467 B.n466 10.6151
R1012 B.n466 B.n465 10.6151
R1013 B.n465 B.n114 10.6151
R1014 B.n461 B.n114 10.6151
R1015 B.n461 B.n460 10.6151
R1016 B.n460 B.n459 10.6151
R1017 B.n459 B.n116 10.6151
R1018 B.n455 B.n116 10.6151
R1019 B.n455 B.n454 10.6151
R1020 B.n454 B.n453 10.6151
R1021 B.n453 B.n118 10.6151
R1022 B.n449 B.n118 10.6151
R1023 B.n449 B.n448 10.6151
R1024 B.n448 B.n447 10.6151
R1025 B.n447 B.n120 10.6151
R1026 B.n443 B.n120 10.6151
R1027 B.n443 B.n442 10.6151
R1028 B.n442 B.n441 10.6151
R1029 B.n441 B.n122 10.6151
R1030 B.n437 B.n122 10.6151
R1031 B.n204 B.n1 10.6151
R1032 B.n207 B.n204 10.6151
R1033 B.n208 B.n207 10.6151
R1034 B.n209 B.n208 10.6151
R1035 B.n209 B.n202 10.6151
R1036 B.n213 B.n202 10.6151
R1037 B.n214 B.n213 10.6151
R1038 B.n215 B.n214 10.6151
R1039 B.n215 B.n200 10.6151
R1040 B.n219 B.n200 10.6151
R1041 B.n220 B.n219 10.6151
R1042 B.n221 B.n220 10.6151
R1043 B.n221 B.n198 10.6151
R1044 B.n225 B.n198 10.6151
R1045 B.n226 B.n225 10.6151
R1046 B.n227 B.n226 10.6151
R1047 B.n227 B.n196 10.6151
R1048 B.n231 B.n196 10.6151
R1049 B.n232 B.n231 10.6151
R1050 B.n233 B.n232 10.6151
R1051 B.n233 B.n194 10.6151
R1052 B.n237 B.n194 10.6151
R1053 B.n238 B.n237 10.6151
R1054 B.n239 B.n238 10.6151
R1055 B.n239 B.n192 10.6151
R1056 B.n243 B.n192 10.6151
R1057 B.n244 B.n243 10.6151
R1058 B.n245 B.n244 10.6151
R1059 B.n245 B.n190 10.6151
R1060 B.n249 B.n190 10.6151
R1061 B.n250 B.n249 10.6151
R1062 B.n251 B.n250 10.6151
R1063 B.n251 B.n188 10.6151
R1064 B.n255 B.n188 10.6151
R1065 B.n256 B.n255 10.6151
R1066 B.n257 B.n256 10.6151
R1067 B.n257 B.n186 10.6151
R1068 B.n262 B.n261 10.6151
R1069 B.n263 B.n262 10.6151
R1070 B.n263 B.n184 10.6151
R1071 B.n267 B.n184 10.6151
R1072 B.n268 B.n267 10.6151
R1073 B.n269 B.n268 10.6151
R1074 B.n269 B.n182 10.6151
R1075 B.n273 B.n182 10.6151
R1076 B.n274 B.n273 10.6151
R1077 B.n275 B.n274 10.6151
R1078 B.n275 B.n180 10.6151
R1079 B.n279 B.n180 10.6151
R1080 B.n280 B.n279 10.6151
R1081 B.n281 B.n280 10.6151
R1082 B.n281 B.n178 10.6151
R1083 B.n285 B.n178 10.6151
R1084 B.n286 B.n285 10.6151
R1085 B.n287 B.n286 10.6151
R1086 B.n287 B.n176 10.6151
R1087 B.n291 B.n176 10.6151
R1088 B.n292 B.n291 10.6151
R1089 B.n293 B.n292 10.6151
R1090 B.n293 B.n174 10.6151
R1091 B.n297 B.n174 10.6151
R1092 B.n298 B.n297 10.6151
R1093 B.n299 B.n298 10.6151
R1094 B.n299 B.n172 10.6151
R1095 B.n303 B.n172 10.6151
R1096 B.n304 B.n303 10.6151
R1097 B.n305 B.n304 10.6151
R1098 B.n305 B.n170 10.6151
R1099 B.n309 B.n170 10.6151
R1100 B.n310 B.n309 10.6151
R1101 B.n311 B.n310 10.6151
R1102 B.n311 B.n168 10.6151
R1103 B.n315 B.n168 10.6151
R1104 B.n316 B.n315 10.6151
R1105 B.n317 B.n316 10.6151
R1106 B.n317 B.n166 10.6151
R1107 B.n321 B.n166 10.6151
R1108 B.n322 B.n321 10.6151
R1109 B.n323 B.n322 10.6151
R1110 B.n323 B.n164 10.6151
R1111 B.n327 B.n164 10.6151
R1112 B.n328 B.n327 10.6151
R1113 B.n329 B.n328 10.6151
R1114 B.n329 B.n162 10.6151
R1115 B.n333 B.n162 10.6151
R1116 B.n334 B.n333 10.6151
R1117 B.n335 B.n334 10.6151
R1118 B.n335 B.n160 10.6151
R1119 B.n339 B.n160 10.6151
R1120 B.n340 B.n339 10.6151
R1121 B.n342 B.n156 10.6151
R1122 B.n346 B.n156 10.6151
R1123 B.n347 B.n346 10.6151
R1124 B.n348 B.n347 10.6151
R1125 B.n348 B.n154 10.6151
R1126 B.n352 B.n154 10.6151
R1127 B.n353 B.n352 10.6151
R1128 B.n354 B.n353 10.6151
R1129 B.n358 B.n357 10.6151
R1130 B.n359 B.n358 10.6151
R1131 B.n359 B.n148 10.6151
R1132 B.n363 B.n148 10.6151
R1133 B.n364 B.n363 10.6151
R1134 B.n365 B.n364 10.6151
R1135 B.n365 B.n146 10.6151
R1136 B.n369 B.n146 10.6151
R1137 B.n370 B.n369 10.6151
R1138 B.n371 B.n370 10.6151
R1139 B.n371 B.n144 10.6151
R1140 B.n375 B.n144 10.6151
R1141 B.n376 B.n375 10.6151
R1142 B.n377 B.n376 10.6151
R1143 B.n377 B.n142 10.6151
R1144 B.n381 B.n142 10.6151
R1145 B.n382 B.n381 10.6151
R1146 B.n383 B.n382 10.6151
R1147 B.n383 B.n140 10.6151
R1148 B.n387 B.n140 10.6151
R1149 B.n388 B.n387 10.6151
R1150 B.n389 B.n388 10.6151
R1151 B.n389 B.n138 10.6151
R1152 B.n393 B.n138 10.6151
R1153 B.n394 B.n393 10.6151
R1154 B.n395 B.n394 10.6151
R1155 B.n395 B.n136 10.6151
R1156 B.n399 B.n136 10.6151
R1157 B.n400 B.n399 10.6151
R1158 B.n401 B.n400 10.6151
R1159 B.n401 B.n134 10.6151
R1160 B.n405 B.n134 10.6151
R1161 B.n406 B.n405 10.6151
R1162 B.n407 B.n406 10.6151
R1163 B.n407 B.n132 10.6151
R1164 B.n411 B.n132 10.6151
R1165 B.n412 B.n411 10.6151
R1166 B.n413 B.n412 10.6151
R1167 B.n413 B.n130 10.6151
R1168 B.n417 B.n130 10.6151
R1169 B.n418 B.n417 10.6151
R1170 B.n419 B.n418 10.6151
R1171 B.n419 B.n128 10.6151
R1172 B.n423 B.n128 10.6151
R1173 B.n424 B.n423 10.6151
R1174 B.n425 B.n424 10.6151
R1175 B.n425 B.n126 10.6151
R1176 B.n429 B.n126 10.6151
R1177 B.n430 B.n429 10.6151
R1178 B.n431 B.n430 10.6151
R1179 B.n431 B.n124 10.6151
R1180 B.n435 B.n124 10.6151
R1181 B.n436 B.n435 10.6151
R1182 B.n789 B.n0 8.11757
R1183 B.n789 B.n1 8.11757
R1184 B.n648 B.n50 6.5566
R1185 B.n636 B.n635 6.5566
R1186 B.n342 B.n341 6.5566
R1187 B.n354 B.n152 6.5566
R1188 B.n651 B.n50 4.05904
R1189 B.n635 B.n634 4.05904
R1190 B.n341 B.n340 4.05904
R1191 B.n357 B.n152 4.05904
R1192 VP.n9 VP.t2 204.118
R1193 VP.n5 VP.t5 170.718
R1194 VP.n29 VP.t1 170.718
R1195 VP.n37 VP.t0 170.718
R1196 VP.n18 VP.t3 170.718
R1197 VP.n10 VP.t4 170.718
R1198 VP.n11 VP.n8 161.3
R1199 VP.n13 VP.n12 161.3
R1200 VP.n14 VP.n7 161.3
R1201 VP.n16 VP.n15 161.3
R1202 VP.n17 VP.n6 161.3
R1203 VP.n36 VP.n0 161.3
R1204 VP.n35 VP.n34 161.3
R1205 VP.n33 VP.n1 161.3
R1206 VP.n32 VP.n31 161.3
R1207 VP.n30 VP.n2 161.3
R1208 VP.n28 VP.n27 161.3
R1209 VP.n26 VP.n3 161.3
R1210 VP.n25 VP.n24 161.3
R1211 VP.n23 VP.n4 161.3
R1212 VP.n22 VP.n21 161.3
R1213 VP.n20 VP.n5 93.694
R1214 VP.n38 VP.n37 93.694
R1215 VP.n19 VP.n18 93.694
R1216 VP.n10 VP.n9 59.4102
R1217 VP.n20 VP.n19 50.5224
R1218 VP.n24 VP.n23 45.4209
R1219 VP.n35 VP.n1 45.4209
R1220 VP.n16 VP.n7 45.4209
R1221 VP.n24 VP.n3 35.7332
R1222 VP.n31 VP.n1 35.7332
R1223 VP.n12 VP.n7 35.7332
R1224 VP.n23 VP.n22 24.5923
R1225 VP.n28 VP.n3 24.5923
R1226 VP.n31 VP.n30 24.5923
R1227 VP.n36 VP.n35 24.5923
R1228 VP.n17 VP.n16 24.5923
R1229 VP.n12 VP.n11 24.5923
R1230 VP.n22 VP.n5 17.2148
R1231 VP.n37 VP.n36 17.2148
R1232 VP.n18 VP.n17 17.2148
R1233 VP.n29 VP.n28 12.2964
R1234 VP.n30 VP.n29 12.2964
R1235 VP.n11 VP.n10 12.2964
R1236 VP.n9 VP.n8 9.22766
R1237 VP.n19 VP.n6 0.278335
R1238 VP.n21 VP.n20 0.278335
R1239 VP.n38 VP.n0 0.278335
R1240 VP.n13 VP.n8 0.189894
R1241 VP.n14 VP.n13 0.189894
R1242 VP.n15 VP.n14 0.189894
R1243 VP.n15 VP.n6 0.189894
R1244 VP.n21 VP.n4 0.189894
R1245 VP.n25 VP.n4 0.189894
R1246 VP.n26 VP.n25 0.189894
R1247 VP.n27 VP.n26 0.189894
R1248 VP.n27 VP.n2 0.189894
R1249 VP.n32 VP.n2 0.189894
R1250 VP.n33 VP.n32 0.189894
R1251 VP.n34 VP.n33 0.189894
R1252 VP.n34 VP.n0 0.189894
R1253 VP VP.n38 0.153485
R1254 VTAIL.n362 VTAIL.n278 756.745
R1255 VTAIL.n86 VTAIL.n2 756.745
R1256 VTAIL.n272 VTAIL.n188 756.745
R1257 VTAIL.n180 VTAIL.n96 756.745
R1258 VTAIL.n306 VTAIL.n305 585
R1259 VTAIL.n311 VTAIL.n310 585
R1260 VTAIL.n313 VTAIL.n312 585
R1261 VTAIL.n302 VTAIL.n301 585
R1262 VTAIL.n319 VTAIL.n318 585
R1263 VTAIL.n321 VTAIL.n320 585
R1264 VTAIL.n298 VTAIL.n297 585
R1265 VTAIL.n327 VTAIL.n326 585
R1266 VTAIL.n329 VTAIL.n328 585
R1267 VTAIL.n294 VTAIL.n293 585
R1268 VTAIL.n335 VTAIL.n334 585
R1269 VTAIL.n337 VTAIL.n336 585
R1270 VTAIL.n290 VTAIL.n289 585
R1271 VTAIL.n343 VTAIL.n342 585
R1272 VTAIL.n345 VTAIL.n344 585
R1273 VTAIL.n286 VTAIL.n285 585
R1274 VTAIL.n352 VTAIL.n351 585
R1275 VTAIL.n353 VTAIL.n284 585
R1276 VTAIL.n355 VTAIL.n354 585
R1277 VTAIL.n282 VTAIL.n281 585
R1278 VTAIL.n361 VTAIL.n360 585
R1279 VTAIL.n363 VTAIL.n362 585
R1280 VTAIL.n30 VTAIL.n29 585
R1281 VTAIL.n35 VTAIL.n34 585
R1282 VTAIL.n37 VTAIL.n36 585
R1283 VTAIL.n26 VTAIL.n25 585
R1284 VTAIL.n43 VTAIL.n42 585
R1285 VTAIL.n45 VTAIL.n44 585
R1286 VTAIL.n22 VTAIL.n21 585
R1287 VTAIL.n51 VTAIL.n50 585
R1288 VTAIL.n53 VTAIL.n52 585
R1289 VTAIL.n18 VTAIL.n17 585
R1290 VTAIL.n59 VTAIL.n58 585
R1291 VTAIL.n61 VTAIL.n60 585
R1292 VTAIL.n14 VTAIL.n13 585
R1293 VTAIL.n67 VTAIL.n66 585
R1294 VTAIL.n69 VTAIL.n68 585
R1295 VTAIL.n10 VTAIL.n9 585
R1296 VTAIL.n76 VTAIL.n75 585
R1297 VTAIL.n77 VTAIL.n8 585
R1298 VTAIL.n79 VTAIL.n78 585
R1299 VTAIL.n6 VTAIL.n5 585
R1300 VTAIL.n85 VTAIL.n84 585
R1301 VTAIL.n87 VTAIL.n86 585
R1302 VTAIL.n273 VTAIL.n272 585
R1303 VTAIL.n271 VTAIL.n270 585
R1304 VTAIL.n192 VTAIL.n191 585
R1305 VTAIL.n265 VTAIL.n264 585
R1306 VTAIL.n263 VTAIL.n194 585
R1307 VTAIL.n262 VTAIL.n261 585
R1308 VTAIL.n197 VTAIL.n195 585
R1309 VTAIL.n256 VTAIL.n255 585
R1310 VTAIL.n254 VTAIL.n253 585
R1311 VTAIL.n201 VTAIL.n200 585
R1312 VTAIL.n248 VTAIL.n247 585
R1313 VTAIL.n246 VTAIL.n245 585
R1314 VTAIL.n205 VTAIL.n204 585
R1315 VTAIL.n240 VTAIL.n239 585
R1316 VTAIL.n238 VTAIL.n237 585
R1317 VTAIL.n209 VTAIL.n208 585
R1318 VTAIL.n232 VTAIL.n231 585
R1319 VTAIL.n230 VTAIL.n229 585
R1320 VTAIL.n213 VTAIL.n212 585
R1321 VTAIL.n224 VTAIL.n223 585
R1322 VTAIL.n222 VTAIL.n221 585
R1323 VTAIL.n217 VTAIL.n216 585
R1324 VTAIL.n181 VTAIL.n180 585
R1325 VTAIL.n179 VTAIL.n178 585
R1326 VTAIL.n100 VTAIL.n99 585
R1327 VTAIL.n173 VTAIL.n172 585
R1328 VTAIL.n171 VTAIL.n102 585
R1329 VTAIL.n170 VTAIL.n169 585
R1330 VTAIL.n105 VTAIL.n103 585
R1331 VTAIL.n164 VTAIL.n163 585
R1332 VTAIL.n162 VTAIL.n161 585
R1333 VTAIL.n109 VTAIL.n108 585
R1334 VTAIL.n156 VTAIL.n155 585
R1335 VTAIL.n154 VTAIL.n153 585
R1336 VTAIL.n113 VTAIL.n112 585
R1337 VTAIL.n148 VTAIL.n147 585
R1338 VTAIL.n146 VTAIL.n145 585
R1339 VTAIL.n117 VTAIL.n116 585
R1340 VTAIL.n140 VTAIL.n139 585
R1341 VTAIL.n138 VTAIL.n137 585
R1342 VTAIL.n121 VTAIL.n120 585
R1343 VTAIL.n132 VTAIL.n131 585
R1344 VTAIL.n130 VTAIL.n129 585
R1345 VTAIL.n125 VTAIL.n124 585
R1346 VTAIL.n307 VTAIL.t4 327.466
R1347 VTAIL.n31 VTAIL.t6 327.466
R1348 VTAIL.n218 VTAIL.t7 327.466
R1349 VTAIL.n126 VTAIL.t0 327.466
R1350 VTAIL.n311 VTAIL.n305 171.744
R1351 VTAIL.n312 VTAIL.n311 171.744
R1352 VTAIL.n312 VTAIL.n301 171.744
R1353 VTAIL.n319 VTAIL.n301 171.744
R1354 VTAIL.n320 VTAIL.n319 171.744
R1355 VTAIL.n320 VTAIL.n297 171.744
R1356 VTAIL.n327 VTAIL.n297 171.744
R1357 VTAIL.n328 VTAIL.n327 171.744
R1358 VTAIL.n328 VTAIL.n293 171.744
R1359 VTAIL.n335 VTAIL.n293 171.744
R1360 VTAIL.n336 VTAIL.n335 171.744
R1361 VTAIL.n336 VTAIL.n289 171.744
R1362 VTAIL.n343 VTAIL.n289 171.744
R1363 VTAIL.n344 VTAIL.n343 171.744
R1364 VTAIL.n344 VTAIL.n285 171.744
R1365 VTAIL.n352 VTAIL.n285 171.744
R1366 VTAIL.n353 VTAIL.n352 171.744
R1367 VTAIL.n354 VTAIL.n353 171.744
R1368 VTAIL.n354 VTAIL.n281 171.744
R1369 VTAIL.n361 VTAIL.n281 171.744
R1370 VTAIL.n362 VTAIL.n361 171.744
R1371 VTAIL.n35 VTAIL.n29 171.744
R1372 VTAIL.n36 VTAIL.n35 171.744
R1373 VTAIL.n36 VTAIL.n25 171.744
R1374 VTAIL.n43 VTAIL.n25 171.744
R1375 VTAIL.n44 VTAIL.n43 171.744
R1376 VTAIL.n44 VTAIL.n21 171.744
R1377 VTAIL.n51 VTAIL.n21 171.744
R1378 VTAIL.n52 VTAIL.n51 171.744
R1379 VTAIL.n52 VTAIL.n17 171.744
R1380 VTAIL.n59 VTAIL.n17 171.744
R1381 VTAIL.n60 VTAIL.n59 171.744
R1382 VTAIL.n60 VTAIL.n13 171.744
R1383 VTAIL.n67 VTAIL.n13 171.744
R1384 VTAIL.n68 VTAIL.n67 171.744
R1385 VTAIL.n68 VTAIL.n9 171.744
R1386 VTAIL.n76 VTAIL.n9 171.744
R1387 VTAIL.n77 VTAIL.n76 171.744
R1388 VTAIL.n78 VTAIL.n77 171.744
R1389 VTAIL.n78 VTAIL.n5 171.744
R1390 VTAIL.n85 VTAIL.n5 171.744
R1391 VTAIL.n86 VTAIL.n85 171.744
R1392 VTAIL.n272 VTAIL.n271 171.744
R1393 VTAIL.n271 VTAIL.n191 171.744
R1394 VTAIL.n264 VTAIL.n191 171.744
R1395 VTAIL.n264 VTAIL.n263 171.744
R1396 VTAIL.n263 VTAIL.n262 171.744
R1397 VTAIL.n262 VTAIL.n195 171.744
R1398 VTAIL.n255 VTAIL.n195 171.744
R1399 VTAIL.n255 VTAIL.n254 171.744
R1400 VTAIL.n254 VTAIL.n200 171.744
R1401 VTAIL.n247 VTAIL.n200 171.744
R1402 VTAIL.n247 VTAIL.n246 171.744
R1403 VTAIL.n246 VTAIL.n204 171.744
R1404 VTAIL.n239 VTAIL.n204 171.744
R1405 VTAIL.n239 VTAIL.n238 171.744
R1406 VTAIL.n238 VTAIL.n208 171.744
R1407 VTAIL.n231 VTAIL.n208 171.744
R1408 VTAIL.n231 VTAIL.n230 171.744
R1409 VTAIL.n230 VTAIL.n212 171.744
R1410 VTAIL.n223 VTAIL.n212 171.744
R1411 VTAIL.n223 VTAIL.n222 171.744
R1412 VTAIL.n222 VTAIL.n216 171.744
R1413 VTAIL.n180 VTAIL.n179 171.744
R1414 VTAIL.n179 VTAIL.n99 171.744
R1415 VTAIL.n172 VTAIL.n99 171.744
R1416 VTAIL.n172 VTAIL.n171 171.744
R1417 VTAIL.n171 VTAIL.n170 171.744
R1418 VTAIL.n170 VTAIL.n103 171.744
R1419 VTAIL.n163 VTAIL.n103 171.744
R1420 VTAIL.n163 VTAIL.n162 171.744
R1421 VTAIL.n162 VTAIL.n108 171.744
R1422 VTAIL.n155 VTAIL.n108 171.744
R1423 VTAIL.n155 VTAIL.n154 171.744
R1424 VTAIL.n154 VTAIL.n112 171.744
R1425 VTAIL.n147 VTAIL.n112 171.744
R1426 VTAIL.n147 VTAIL.n146 171.744
R1427 VTAIL.n146 VTAIL.n116 171.744
R1428 VTAIL.n139 VTAIL.n116 171.744
R1429 VTAIL.n139 VTAIL.n138 171.744
R1430 VTAIL.n138 VTAIL.n120 171.744
R1431 VTAIL.n131 VTAIL.n120 171.744
R1432 VTAIL.n131 VTAIL.n130 171.744
R1433 VTAIL.n130 VTAIL.n124 171.744
R1434 VTAIL.t4 VTAIL.n305 85.8723
R1435 VTAIL.t6 VTAIL.n29 85.8723
R1436 VTAIL.t7 VTAIL.n216 85.8723
R1437 VTAIL.t0 VTAIL.n124 85.8723
R1438 VTAIL.n187 VTAIL.n186 53.1234
R1439 VTAIL.n95 VTAIL.n94 53.1234
R1440 VTAIL.n1 VTAIL.n0 53.1232
R1441 VTAIL.n93 VTAIL.n92 53.1232
R1442 VTAIL.n367 VTAIL.n366 32.1853
R1443 VTAIL.n91 VTAIL.n90 32.1853
R1444 VTAIL.n277 VTAIL.n276 32.1853
R1445 VTAIL.n185 VTAIL.n184 32.1853
R1446 VTAIL.n95 VTAIL.n93 30.7117
R1447 VTAIL.n367 VTAIL.n277 28.4703
R1448 VTAIL.n307 VTAIL.n306 16.3895
R1449 VTAIL.n31 VTAIL.n30 16.3895
R1450 VTAIL.n218 VTAIL.n217 16.3895
R1451 VTAIL.n126 VTAIL.n125 16.3895
R1452 VTAIL.n355 VTAIL.n284 13.1884
R1453 VTAIL.n79 VTAIL.n8 13.1884
R1454 VTAIL.n265 VTAIL.n194 13.1884
R1455 VTAIL.n173 VTAIL.n102 13.1884
R1456 VTAIL.n310 VTAIL.n309 12.8005
R1457 VTAIL.n351 VTAIL.n350 12.8005
R1458 VTAIL.n356 VTAIL.n282 12.8005
R1459 VTAIL.n34 VTAIL.n33 12.8005
R1460 VTAIL.n75 VTAIL.n74 12.8005
R1461 VTAIL.n80 VTAIL.n6 12.8005
R1462 VTAIL.n266 VTAIL.n192 12.8005
R1463 VTAIL.n261 VTAIL.n196 12.8005
R1464 VTAIL.n221 VTAIL.n220 12.8005
R1465 VTAIL.n174 VTAIL.n100 12.8005
R1466 VTAIL.n169 VTAIL.n104 12.8005
R1467 VTAIL.n129 VTAIL.n128 12.8005
R1468 VTAIL.n313 VTAIL.n304 12.0247
R1469 VTAIL.n349 VTAIL.n286 12.0247
R1470 VTAIL.n360 VTAIL.n359 12.0247
R1471 VTAIL.n37 VTAIL.n28 12.0247
R1472 VTAIL.n73 VTAIL.n10 12.0247
R1473 VTAIL.n84 VTAIL.n83 12.0247
R1474 VTAIL.n270 VTAIL.n269 12.0247
R1475 VTAIL.n260 VTAIL.n197 12.0247
R1476 VTAIL.n224 VTAIL.n215 12.0247
R1477 VTAIL.n178 VTAIL.n177 12.0247
R1478 VTAIL.n168 VTAIL.n105 12.0247
R1479 VTAIL.n132 VTAIL.n123 12.0247
R1480 VTAIL.n314 VTAIL.n302 11.249
R1481 VTAIL.n346 VTAIL.n345 11.249
R1482 VTAIL.n363 VTAIL.n280 11.249
R1483 VTAIL.n38 VTAIL.n26 11.249
R1484 VTAIL.n70 VTAIL.n69 11.249
R1485 VTAIL.n87 VTAIL.n4 11.249
R1486 VTAIL.n273 VTAIL.n190 11.249
R1487 VTAIL.n257 VTAIL.n256 11.249
R1488 VTAIL.n225 VTAIL.n213 11.249
R1489 VTAIL.n181 VTAIL.n98 11.249
R1490 VTAIL.n165 VTAIL.n164 11.249
R1491 VTAIL.n133 VTAIL.n121 11.249
R1492 VTAIL.n318 VTAIL.n317 10.4732
R1493 VTAIL.n342 VTAIL.n288 10.4732
R1494 VTAIL.n364 VTAIL.n278 10.4732
R1495 VTAIL.n42 VTAIL.n41 10.4732
R1496 VTAIL.n66 VTAIL.n12 10.4732
R1497 VTAIL.n88 VTAIL.n2 10.4732
R1498 VTAIL.n274 VTAIL.n188 10.4732
R1499 VTAIL.n253 VTAIL.n199 10.4732
R1500 VTAIL.n229 VTAIL.n228 10.4732
R1501 VTAIL.n182 VTAIL.n96 10.4732
R1502 VTAIL.n161 VTAIL.n107 10.4732
R1503 VTAIL.n137 VTAIL.n136 10.4732
R1504 VTAIL.n321 VTAIL.n300 9.69747
R1505 VTAIL.n341 VTAIL.n290 9.69747
R1506 VTAIL.n45 VTAIL.n24 9.69747
R1507 VTAIL.n65 VTAIL.n14 9.69747
R1508 VTAIL.n252 VTAIL.n201 9.69747
R1509 VTAIL.n232 VTAIL.n211 9.69747
R1510 VTAIL.n160 VTAIL.n109 9.69747
R1511 VTAIL.n140 VTAIL.n119 9.69747
R1512 VTAIL.n366 VTAIL.n365 9.45567
R1513 VTAIL.n90 VTAIL.n89 9.45567
R1514 VTAIL.n276 VTAIL.n275 9.45567
R1515 VTAIL.n184 VTAIL.n183 9.45567
R1516 VTAIL.n365 VTAIL.n364 9.3005
R1517 VTAIL.n280 VTAIL.n279 9.3005
R1518 VTAIL.n359 VTAIL.n358 9.3005
R1519 VTAIL.n357 VTAIL.n356 9.3005
R1520 VTAIL.n296 VTAIL.n295 9.3005
R1521 VTAIL.n325 VTAIL.n324 9.3005
R1522 VTAIL.n323 VTAIL.n322 9.3005
R1523 VTAIL.n300 VTAIL.n299 9.3005
R1524 VTAIL.n317 VTAIL.n316 9.3005
R1525 VTAIL.n315 VTAIL.n314 9.3005
R1526 VTAIL.n304 VTAIL.n303 9.3005
R1527 VTAIL.n309 VTAIL.n308 9.3005
R1528 VTAIL.n331 VTAIL.n330 9.3005
R1529 VTAIL.n333 VTAIL.n332 9.3005
R1530 VTAIL.n292 VTAIL.n291 9.3005
R1531 VTAIL.n339 VTAIL.n338 9.3005
R1532 VTAIL.n341 VTAIL.n340 9.3005
R1533 VTAIL.n288 VTAIL.n287 9.3005
R1534 VTAIL.n347 VTAIL.n346 9.3005
R1535 VTAIL.n349 VTAIL.n348 9.3005
R1536 VTAIL.n350 VTAIL.n283 9.3005
R1537 VTAIL.n89 VTAIL.n88 9.3005
R1538 VTAIL.n4 VTAIL.n3 9.3005
R1539 VTAIL.n83 VTAIL.n82 9.3005
R1540 VTAIL.n81 VTAIL.n80 9.3005
R1541 VTAIL.n20 VTAIL.n19 9.3005
R1542 VTAIL.n49 VTAIL.n48 9.3005
R1543 VTAIL.n47 VTAIL.n46 9.3005
R1544 VTAIL.n24 VTAIL.n23 9.3005
R1545 VTAIL.n41 VTAIL.n40 9.3005
R1546 VTAIL.n39 VTAIL.n38 9.3005
R1547 VTAIL.n28 VTAIL.n27 9.3005
R1548 VTAIL.n33 VTAIL.n32 9.3005
R1549 VTAIL.n55 VTAIL.n54 9.3005
R1550 VTAIL.n57 VTAIL.n56 9.3005
R1551 VTAIL.n16 VTAIL.n15 9.3005
R1552 VTAIL.n63 VTAIL.n62 9.3005
R1553 VTAIL.n65 VTAIL.n64 9.3005
R1554 VTAIL.n12 VTAIL.n11 9.3005
R1555 VTAIL.n71 VTAIL.n70 9.3005
R1556 VTAIL.n73 VTAIL.n72 9.3005
R1557 VTAIL.n74 VTAIL.n7 9.3005
R1558 VTAIL.n244 VTAIL.n243 9.3005
R1559 VTAIL.n203 VTAIL.n202 9.3005
R1560 VTAIL.n250 VTAIL.n249 9.3005
R1561 VTAIL.n252 VTAIL.n251 9.3005
R1562 VTAIL.n199 VTAIL.n198 9.3005
R1563 VTAIL.n258 VTAIL.n257 9.3005
R1564 VTAIL.n260 VTAIL.n259 9.3005
R1565 VTAIL.n196 VTAIL.n193 9.3005
R1566 VTAIL.n275 VTAIL.n274 9.3005
R1567 VTAIL.n190 VTAIL.n189 9.3005
R1568 VTAIL.n269 VTAIL.n268 9.3005
R1569 VTAIL.n267 VTAIL.n266 9.3005
R1570 VTAIL.n242 VTAIL.n241 9.3005
R1571 VTAIL.n207 VTAIL.n206 9.3005
R1572 VTAIL.n236 VTAIL.n235 9.3005
R1573 VTAIL.n234 VTAIL.n233 9.3005
R1574 VTAIL.n211 VTAIL.n210 9.3005
R1575 VTAIL.n228 VTAIL.n227 9.3005
R1576 VTAIL.n226 VTAIL.n225 9.3005
R1577 VTAIL.n215 VTAIL.n214 9.3005
R1578 VTAIL.n220 VTAIL.n219 9.3005
R1579 VTAIL.n152 VTAIL.n151 9.3005
R1580 VTAIL.n111 VTAIL.n110 9.3005
R1581 VTAIL.n158 VTAIL.n157 9.3005
R1582 VTAIL.n160 VTAIL.n159 9.3005
R1583 VTAIL.n107 VTAIL.n106 9.3005
R1584 VTAIL.n166 VTAIL.n165 9.3005
R1585 VTAIL.n168 VTAIL.n167 9.3005
R1586 VTAIL.n104 VTAIL.n101 9.3005
R1587 VTAIL.n183 VTAIL.n182 9.3005
R1588 VTAIL.n98 VTAIL.n97 9.3005
R1589 VTAIL.n177 VTAIL.n176 9.3005
R1590 VTAIL.n175 VTAIL.n174 9.3005
R1591 VTAIL.n150 VTAIL.n149 9.3005
R1592 VTAIL.n115 VTAIL.n114 9.3005
R1593 VTAIL.n144 VTAIL.n143 9.3005
R1594 VTAIL.n142 VTAIL.n141 9.3005
R1595 VTAIL.n119 VTAIL.n118 9.3005
R1596 VTAIL.n136 VTAIL.n135 9.3005
R1597 VTAIL.n134 VTAIL.n133 9.3005
R1598 VTAIL.n123 VTAIL.n122 9.3005
R1599 VTAIL.n128 VTAIL.n127 9.3005
R1600 VTAIL.n322 VTAIL.n298 8.92171
R1601 VTAIL.n338 VTAIL.n337 8.92171
R1602 VTAIL.n46 VTAIL.n22 8.92171
R1603 VTAIL.n62 VTAIL.n61 8.92171
R1604 VTAIL.n249 VTAIL.n248 8.92171
R1605 VTAIL.n233 VTAIL.n209 8.92171
R1606 VTAIL.n157 VTAIL.n156 8.92171
R1607 VTAIL.n141 VTAIL.n117 8.92171
R1608 VTAIL.n326 VTAIL.n325 8.14595
R1609 VTAIL.n334 VTAIL.n292 8.14595
R1610 VTAIL.n50 VTAIL.n49 8.14595
R1611 VTAIL.n58 VTAIL.n16 8.14595
R1612 VTAIL.n245 VTAIL.n203 8.14595
R1613 VTAIL.n237 VTAIL.n236 8.14595
R1614 VTAIL.n153 VTAIL.n111 8.14595
R1615 VTAIL.n145 VTAIL.n144 8.14595
R1616 VTAIL.n329 VTAIL.n296 7.3702
R1617 VTAIL.n333 VTAIL.n294 7.3702
R1618 VTAIL.n53 VTAIL.n20 7.3702
R1619 VTAIL.n57 VTAIL.n18 7.3702
R1620 VTAIL.n244 VTAIL.n205 7.3702
R1621 VTAIL.n240 VTAIL.n207 7.3702
R1622 VTAIL.n152 VTAIL.n113 7.3702
R1623 VTAIL.n148 VTAIL.n115 7.3702
R1624 VTAIL.n330 VTAIL.n329 6.59444
R1625 VTAIL.n330 VTAIL.n294 6.59444
R1626 VTAIL.n54 VTAIL.n53 6.59444
R1627 VTAIL.n54 VTAIL.n18 6.59444
R1628 VTAIL.n241 VTAIL.n205 6.59444
R1629 VTAIL.n241 VTAIL.n240 6.59444
R1630 VTAIL.n149 VTAIL.n113 6.59444
R1631 VTAIL.n149 VTAIL.n148 6.59444
R1632 VTAIL.n326 VTAIL.n296 5.81868
R1633 VTAIL.n334 VTAIL.n333 5.81868
R1634 VTAIL.n50 VTAIL.n20 5.81868
R1635 VTAIL.n58 VTAIL.n57 5.81868
R1636 VTAIL.n245 VTAIL.n244 5.81868
R1637 VTAIL.n237 VTAIL.n207 5.81868
R1638 VTAIL.n153 VTAIL.n152 5.81868
R1639 VTAIL.n145 VTAIL.n115 5.81868
R1640 VTAIL.n325 VTAIL.n298 5.04292
R1641 VTAIL.n337 VTAIL.n292 5.04292
R1642 VTAIL.n49 VTAIL.n22 5.04292
R1643 VTAIL.n61 VTAIL.n16 5.04292
R1644 VTAIL.n248 VTAIL.n203 5.04292
R1645 VTAIL.n236 VTAIL.n209 5.04292
R1646 VTAIL.n156 VTAIL.n111 5.04292
R1647 VTAIL.n144 VTAIL.n117 5.04292
R1648 VTAIL.n322 VTAIL.n321 4.26717
R1649 VTAIL.n338 VTAIL.n290 4.26717
R1650 VTAIL.n46 VTAIL.n45 4.26717
R1651 VTAIL.n62 VTAIL.n14 4.26717
R1652 VTAIL.n249 VTAIL.n201 4.26717
R1653 VTAIL.n233 VTAIL.n232 4.26717
R1654 VTAIL.n157 VTAIL.n109 4.26717
R1655 VTAIL.n141 VTAIL.n140 4.26717
R1656 VTAIL.n308 VTAIL.n307 3.70982
R1657 VTAIL.n32 VTAIL.n31 3.70982
R1658 VTAIL.n219 VTAIL.n218 3.70982
R1659 VTAIL.n127 VTAIL.n126 3.70982
R1660 VTAIL.n318 VTAIL.n300 3.49141
R1661 VTAIL.n342 VTAIL.n341 3.49141
R1662 VTAIL.n366 VTAIL.n278 3.49141
R1663 VTAIL.n42 VTAIL.n24 3.49141
R1664 VTAIL.n66 VTAIL.n65 3.49141
R1665 VTAIL.n90 VTAIL.n2 3.49141
R1666 VTAIL.n276 VTAIL.n188 3.49141
R1667 VTAIL.n253 VTAIL.n252 3.49141
R1668 VTAIL.n229 VTAIL.n211 3.49141
R1669 VTAIL.n184 VTAIL.n96 3.49141
R1670 VTAIL.n161 VTAIL.n160 3.49141
R1671 VTAIL.n137 VTAIL.n119 3.49141
R1672 VTAIL.n317 VTAIL.n302 2.71565
R1673 VTAIL.n345 VTAIL.n288 2.71565
R1674 VTAIL.n364 VTAIL.n363 2.71565
R1675 VTAIL.n41 VTAIL.n26 2.71565
R1676 VTAIL.n69 VTAIL.n12 2.71565
R1677 VTAIL.n88 VTAIL.n87 2.71565
R1678 VTAIL.n274 VTAIL.n273 2.71565
R1679 VTAIL.n256 VTAIL.n199 2.71565
R1680 VTAIL.n228 VTAIL.n213 2.71565
R1681 VTAIL.n182 VTAIL.n181 2.71565
R1682 VTAIL.n164 VTAIL.n107 2.71565
R1683 VTAIL.n136 VTAIL.n121 2.71565
R1684 VTAIL.n185 VTAIL.n95 2.24188
R1685 VTAIL.n277 VTAIL.n187 2.24188
R1686 VTAIL.n93 VTAIL.n91 2.24188
R1687 VTAIL.n0 VTAIL.t2 2.02196
R1688 VTAIL.n0 VTAIL.t1 2.02196
R1689 VTAIL.n92 VTAIL.t9 2.02196
R1690 VTAIL.n92 VTAIL.t11 2.02196
R1691 VTAIL.n186 VTAIL.t10 2.02196
R1692 VTAIL.n186 VTAIL.t8 2.02196
R1693 VTAIL.n94 VTAIL.t3 2.02196
R1694 VTAIL.n94 VTAIL.t5 2.02196
R1695 VTAIL.n314 VTAIL.n313 1.93989
R1696 VTAIL.n346 VTAIL.n286 1.93989
R1697 VTAIL.n360 VTAIL.n280 1.93989
R1698 VTAIL.n38 VTAIL.n37 1.93989
R1699 VTAIL.n70 VTAIL.n10 1.93989
R1700 VTAIL.n84 VTAIL.n4 1.93989
R1701 VTAIL.n270 VTAIL.n190 1.93989
R1702 VTAIL.n257 VTAIL.n197 1.93989
R1703 VTAIL.n225 VTAIL.n224 1.93989
R1704 VTAIL.n178 VTAIL.n98 1.93989
R1705 VTAIL.n165 VTAIL.n105 1.93989
R1706 VTAIL.n133 VTAIL.n132 1.93989
R1707 VTAIL VTAIL.n367 1.62334
R1708 VTAIL.n187 VTAIL.n185 1.59102
R1709 VTAIL.n91 VTAIL.n1 1.59102
R1710 VTAIL.n310 VTAIL.n304 1.16414
R1711 VTAIL.n351 VTAIL.n349 1.16414
R1712 VTAIL.n359 VTAIL.n282 1.16414
R1713 VTAIL.n34 VTAIL.n28 1.16414
R1714 VTAIL.n75 VTAIL.n73 1.16414
R1715 VTAIL.n83 VTAIL.n6 1.16414
R1716 VTAIL.n269 VTAIL.n192 1.16414
R1717 VTAIL.n261 VTAIL.n260 1.16414
R1718 VTAIL.n221 VTAIL.n215 1.16414
R1719 VTAIL.n177 VTAIL.n100 1.16414
R1720 VTAIL.n169 VTAIL.n168 1.16414
R1721 VTAIL.n129 VTAIL.n123 1.16414
R1722 VTAIL VTAIL.n1 0.619035
R1723 VTAIL.n309 VTAIL.n306 0.388379
R1724 VTAIL.n350 VTAIL.n284 0.388379
R1725 VTAIL.n356 VTAIL.n355 0.388379
R1726 VTAIL.n33 VTAIL.n30 0.388379
R1727 VTAIL.n74 VTAIL.n8 0.388379
R1728 VTAIL.n80 VTAIL.n79 0.388379
R1729 VTAIL.n266 VTAIL.n265 0.388379
R1730 VTAIL.n196 VTAIL.n194 0.388379
R1731 VTAIL.n220 VTAIL.n217 0.388379
R1732 VTAIL.n174 VTAIL.n173 0.388379
R1733 VTAIL.n104 VTAIL.n102 0.388379
R1734 VTAIL.n128 VTAIL.n125 0.388379
R1735 VTAIL.n308 VTAIL.n303 0.155672
R1736 VTAIL.n315 VTAIL.n303 0.155672
R1737 VTAIL.n316 VTAIL.n315 0.155672
R1738 VTAIL.n316 VTAIL.n299 0.155672
R1739 VTAIL.n323 VTAIL.n299 0.155672
R1740 VTAIL.n324 VTAIL.n323 0.155672
R1741 VTAIL.n324 VTAIL.n295 0.155672
R1742 VTAIL.n331 VTAIL.n295 0.155672
R1743 VTAIL.n332 VTAIL.n331 0.155672
R1744 VTAIL.n332 VTAIL.n291 0.155672
R1745 VTAIL.n339 VTAIL.n291 0.155672
R1746 VTAIL.n340 VTAIL.n339 0.155672
R1747 VTAIL.n340 VTAIL.n287 0.155672
R1748 VTAIL.n347 VTAIL.n287 0.155672
R1749 VTAIL.n348 VTAIL.n347 0.155672
R1750 VTAIL.n348 VTAIL.n283 0.155672
R1751 VTAIL.n357 VTAIL.n283 0.155672
R1752 VTAIL.n358 VTAIL.n357 0.155672
R1753 VTAIL.n358 VTAIL.n279 0.155672
R1754 VTAIL.n365 VTAIL.n279 0.155672
R1755 VTAIL.n32 VTAIL.n27 0.155672
R1756 VTAIL.n39 VTAIL.n27 0.155672
R1757 VTAIL.n40 VTAIL.n39 0.155672
R1758 VTAIL.n40 VTAIL.n23 0.155672
R1759 VTAIL.n47 VTAIL.n23 0.155672
R1760 VTAIL.n48 VTAIL.n47 0.155672
R1761 VTAIL.n48 VTAIL.n19 0.155672
R1762 VTAIL.n55 VTAIL.n19 0.155672
R1763 VTAIL.n56 VTAIL.n55 0.155672
R1764 VTAIL.n56 VTAIL.n15 0.155672
R1765 VTAIL.n63 VTAIL.n15 0.155672
R1766 VTAIL.n64 VTAIL.n63 0.155672
R1767 VTAIL.n64 VTAIL.n11 0.155672
R1768 VTAIL.n71 VTAIL.n11 0.155672
R1769 VTAIL.n72 VTAIL.n71 0.155672
R1770 VTAIL.n72 VTAIL.n7 0.155672
R1771 VTAIL.n81 VTAIL.n7 0.155672
R1772 VTAIL.n82 VTAIL.n81 0.155672
R1773 VTAIL.n82 VTAIL.n3 0.155672
R1774 VTAIL.n89 VTAIL.n3 0.155672
R1775 VTAIL.n275 VTAIL.n189 0.155672
R1776 VTAIL.n268 VTAIL.n189 0.155672
R1777 VTAIL.n268 VTAIL.n267 0.155672
R1778 VTAIL.n267 VTAIL.n193 0.155672
R1779 VTAIL.n259 VTAIL.n193 0.155672
R1780 VTAIL.n259 VTAIL.n258 0.155672
R1781 VTAIL.n258 VTAIL.n198 0.155672
R1782 VTAIL.n251 VTAIL.n198 0.155672
R1783 VTAIL.n251 VTAIL.n250 0.155672
R1784 VTAIL.n250 VTAIL.n202 0.155672
R1785 VTAIL.n243 VTAIL.n202 0.155672
R1786 VTAIL.n243 VTAIL.n242 0.155672
R1787 VTAIL.n242 VTAIL.n206 0.155672
R1788 VTAIL.n235 VTAIL.n206 0.155672
R1789 VTAIL.n235 VTAIL.n234 0.155672
R1790 VTAIL.n234 VTAIL.n210 0.155672
R1791 VTAIL.n227 VTAIL.n210 0.155672
R1792 VTAIL.n227 VTAIL.n226 0.155672
R1793 VTAIL.n226 VTAIL.n214 0.155672
R1794 VTAIL.n219 VTAIL.n214 0.155672
R1795 VTAIL.n183 VTAIL.n97 0.155672
R1796 VTAIL.n176 VTAIL.n97 0.155672
R1797 VTAIL.n176 VTAIL.n175 0.155672
R1798 VTAIL.n175 VTAIL.n101 0.155672
R1799 VTAIL.n167 VTAIL.n101 0.155672
R1800 VTAIL.n167 VTAIL.n166 0.155672
R1801 VTAIL.n166 VTAIL.n106 0.155672
R1802 VTAIL.n159 VTAIL.n106 0.155672
R1803 VTAIL.n159 VTAIL.n158 0.155672
R1804 VTAIL.n158 VTAIL.n110 0.155672
R1805 VTAIL.n151 VTAIL.n110 0.155672
R1806 VTAIL.n151 VTAIL.n150 0.155672
R1807 VTAIL.n150 VTAIL.n114 0.155672
R1808 VTAIL.n143 VTAIL.n114 0.155672
R1809 VTAIL.n143 VTAIL.n142 0.155672
R1810 VTAIL.n142 VTAIL.n118 0.155672
R1811 VTAIL.n135 VTAIL.n118 0.155672
R1812 VTAIL.n135 VTAIL.n134 0.155672
R1813 VTAIL.n134 VTAIL.n122 0.155672
R1814 VTAIL.n127 VTAIL.n122 0.155672
R1815 VDD1.n84 VDD1.n0 756.745
R1816 VDD1.n173 VDD1.n89 756.745
R1817 VDD1.n85 VDD1.n84 585
R1818 VDD1.n83 VDD1.n82 585
R1819 VDD1.n4 VDD1.n3 585
R1820 VDD1.n77 VDD1.n76 585
R1821 VDD1.n75 VDD1.n6 585
R1822 VDD1.n74 VDD1.n73 585
R1823 VDD1.n9 VDD1.n7 585
R1824 VDD1.n68 VDD1.n67 585
R1825 VDD1.n66 VDD1.n65 585
R1826 VDD1.n13 VDD1.n12 585
R1827 VDD1.n60 VDD1.n59 585
R1828 VDD1.n58 VDD1.n57 585
R1829 VDD1.n17 VDD1.n16 585
R1830 VDD1.n52 VDD1.n51 585
R1831 VDD1.n50 VDD1.n49 585
R1832 VDD1.n21 VDD1.n20 585
R1833 VDD1.n44 VDD1.n43 585
R1834 VDD1.n42 VDD1.n41 585
R1835 VDD1.n25 VDD1.n24 585
R1836 VDD1.n36 VDD1.n35 585
R1837 VDD1.n34 VDD1.n33 585
R1838 VDD1.n29 VDD1.n28 585
R1839 VDD1.n117 VDD1.n116 585
R1840 VDD1.n122 VDD1.n121 585
R1841 VDD1.n124 VDD1.n123 585
R1842 VDD1.n113 VDD1.n112 585
R1843 VDD1.n130 VDD1.n129 585
R1844 VDD1.n132 VDD1.n131 585
R1845 VDD1.n109 VDD1.n108 585
R1846 VDD1.n138 VDD1.n137 585
R1847 VDD1.n140 VDD1.n139 585
R1848 VDD1.n105 VDD1.n104 585
R1849 VDD1.n146 VDD1.n145 585
R1850 VDD1.n148 VDD1.n147 585
R1851 VDD1.n101 VDD1.n100 585
R1852 VDD1.n154 VDD1.n153 585
R1853 VDD1.n156 VDD1.n155 585
R1854 VDD1.n97 VDD1.n96 585
R1855 VDD1.n163 VDD1.n162 585
R1856 VDD1.n164 VDD1.n95 585
R1857 VDD1.n166 VDD1.n165 585
R1858 VDD1.n93 VDD1.n92 585
R1859 VDD1.n172 VDD1.n171 585
R1860 VDD1.n174 VDD1.n173 585
R1861 VDD1.n30 VDD1.t3 327.466
R1862 VDD1.n118 VDD1.t0 327.466
R1863 VDD1.n84 VDD1.n83 171.744
R1864 VDD1.n83 VDD1.n3 171.744
R1865 VDD1.n76 VDD1.n3 171.744
R1866 VDD1.n76 VDD1.n75 171.744
R1867 VDD1.n75 VDD1.n74 171.744
R1868 VDD1.n74 VDD1.n7 171.744
R1869 VDD1.n67 VDD1.n7 171.744
R1870 VDD1.n67 VDD1.n66 171.744
R1871 VDD1.n66 VDD1.n12 171.744
R1872 VDD1.n59 VDD1.n12 171.744
R1873 VDD1.n59 VDD1.n58 171.744
R1874 VDD1.n58 VDD1.n16 171.744
R1875 VDD1.n51 VDD1.n16 171.744
R1876 VDD1.n51 VDD1.n50 171.744
R1877 VDD1.n50 VDD1.n20 171.744
R1878 VDD1.n43 VDD1.n20 171.744
R1879 VDD1.n43 VDD1.n42 171.744
R1880 VDD1.n42 VDD1.n24 171.744
R1881 VDD1.n35 VDD1.n24 171.744
R1882 VDD1.n35 VDD1.n34 171.744
R1883 VDD1.n34 VDD1.n28 171.744
R1884 VDD1.n122 VDD1.n116 171.744
R1885 VDD1.n123 VDD1.n122 171.744
R1886 VDD1.n123 VDD1.n112 171.744
R1887 VDD1.n130 VDD1.n112 171.744
R1888 VDD1.n131 VDD1.n130 171.744
R1889 VDD1.n131 VDD1.n108 171.744
R1890 VDD1.n138 VDD1.n108 171.744
R1891 VDD1.n139 VDD1.n138 171.744
R1892 VDD1.n139 VDD1.n104 171.744
R1893 VDD1.n146 VDD1.n104 171.744
R1894 VDD1.n147 VDD1.n146 171.744
R1895 VDD1.n147 VDD1.n100 171.744
R1896 VDD1.n154 VDD1.n100 171.744
R1897 VDD1.n155 VDD1.n154 171.744
R1898 VDD1.n155 VDD1.n96 171.744
R1899 VDD1.n163 VDD1.n96 171.744
R1900 VDD1.n164 VDD1.n163 171.744
R1901 VDD1.n165 VDD1.n164 171.744
R1902 VDD1.n165 VDD1.n92 171.744
R1903 VDD1.n172 VDD1.n92 171.744
R1904 VDD1.n173 VDD1.n172 171.744
R1905 VDD1.t3 VDD1.n28 85.8723
R1906 VDD1.t0 VDD1.n116 85.8723
R1907 VDD1.n179 VDD1.n178 70.3069
R1908 VDD1.n181 VDD1.n180 69.8019
R1909 VDD1 VDD1.n88 50.6034
R1910 VDD1.n179 VDD1.n177 50.4898
R1911 VDD1.n181 VDD1.n179 46.5655
R1912 VDD1.n30 VDD1.n29 16.3895
R1913 VDD1.n118 VDD1.n117 16.3895
R1914 VDD1.n77 VDD1.n6 13.1884
R1915 VDD1.n166 VDD1.n95 13.1884
R1916 VDD1.n78 VDD1.n4 12.8005
R1917 VDD1.n73 VDD1.n8 12.8005
R1918 VDD1.n33 VDD1.n32 12.8005
R1919 VDD1.n121 VDD1.n120 12.8005
R1920 VDD1.n162 VDD1.n161 12.8005
R1921 VDD1.n167 VDD1.n93 12.8005
R1922 VDD1.n82 VDD1.n81 12.0247
R1923 VDD1.n72 VDD1.n9 12.0247
R1924 VDD1.n36 VDD1.n27 12.0247
R1925 VDD1.n124 VDD1.n115 12.0247
R1926 VDD1.n160 VDD1.n97 12.0247
R1927 VDD1.n171 VDD1.n170 12.0247
R1928 VDD1.n85 VDD1.n2 11.249
R1929 VDD1.n69 VDD1.n68 11.249
R1930 VDD1.n37 VDD1.n25 11.249
R1931 VDD1.n125 VDD1.n113 11.249
R1932 VDD1.n157 VDD1.n156 11.249
R1933 VDD1.n174 VDD1.n91 11.249
R1934 VDD1.n86 VDD1.n0 10.4732
R1935 VDD1.n65 VDD1.n11 10.4732
R1936 VDD1.n41 VDD1.n40 10.4732
R1937 VDD1.n129 VDD1.n128 10.4732
R1938 VDD1.n153 VDD1.n99 10.4732
R1939 VDD1.n175 VDD1.n89 10.4732
R1940 VDD1.n64 VDD1.n13 9.69747
R1941 VDD1.n44 VDD1.n23 9.69747
R1942 VDD1.n132 VDD1.n111 9.69747
R1943 VDD1.n152 VDD1.n101 9.69747
R1944 VDD1.n88 VDD1.n87 9.45567
R1945 VDD1.n177 VDD1.n176 9.45567
R1946 VDD1.n56 VDD1.n55 9.3005
R1947 VDD1.n15 VDD1.n14 9.3005
R1948 VDD1.n62 VDD1.n61 9.3005
R1949 VDD1.n64 VDD1.n63 9.3005
R1950 VDD1.n11 VDD1.n10 9.3005
R1951 VDD1.n70 VDD1.n69 9.3005
R1952 VDD1.n72 VDD1.n71 9.3005
R1953 VDD1.n8 VDD1.n5 9.3005
R1954 VDD1.n87 VDD1.n86 9.3005
R1955 VDD1.n2 VDD1.n1 9.3005
R1956 VDD1.n81 VDD1.n80 9.3005
R1957 VDD1.n79 VDD1.n78 9.3005
R1958 VDD1.n54 VDD1.n53 9.3005
R1959 VDD1.n19 VDD1.n18 9.3005
R1960 VDD1.n48 VDD1.n47 9.3005
R1961 VDD1.n46 VDD1.n45 9.3005
R1962 VDD1.n23 VDD1.n22 9.3005
R1963 VDD1.n40 VDD1.n39 9.3005
R1964 VDD1.n38 VDD1.n37 9.3005
R1965 VDD1.n27 VDD1.n26 9.3005
R1966 VDD1.n32 VDD1.n31 9.3005
R1967 VDD1.n176 VDD1.n175 9.3005
R1968 VDD1.n91 VDD1.n90 9.3005
R1969 VDD1.n170 VDD1.n169 9.3005
R1970 VDD1.n168 VDD1.n167 9.3005
R1971 VDD1.n107 VDD1.n106 9.3005
R1972 VDD1.n136 VDD1.n135 9.3005
R1973 VDD1.n134 VDD1.n133 9.3005
R1974 VDD1.n111 VDD1.n110 9.3005
R1975 VDD1.n128 VDD1.n127 9.3005
R1976 VDD1.n126 VDD1.n125 9.3005
R1977 VDD1.n115 VDD1.n114 9.3005
R1978 VDD1.n120 VDD1.n119 9.3005
R1979 VDD1.n142 VDD1.n141 9.3005
R1980 VDD1.n144 VDD1.n143 9.3005
R1981 VDD1.n103 VDD1.n102 9.3005
R1982 VDD1.n150 VDD1.n149 9.3005
R1983 VDD1.n152 VDD1.n151 9.3005
R1984 VDD1.n99 VDD1.n98 9.3005
R1985 VDD1.n158 VDD1.n157 9.3005
R1986 VDD1.n160 VDD1.n159 9.3005
R1987 VDD1.n161 VDD1.n94 9.3005
R1988 VDD1.n61 VDD1.n60 8.92171
R1989 VDD1.n45 VDD1.n21 8.92171
R1990 VDD1.n133 VDD1.n109 8.92171
R1991 VDD1.n149 VDD1.n148 8.92171
R1992 VDD1.n57 VDD1.n15 8.14595
R1993 VDD1.n49 VDD1.n48 8.14595
R1994 VDD1.n137 VDD1.n136 8.14595
R1995 VDD1.n145 VDD1.n103 8.14595
R1996 VDD1.n56 VDD1.n17 7.3702
R1997 VDD1.n52 VDD1.n19 7.3702
R1998 VDD1.n140 VDD1.n107 7.3702
R1999 VDD1.n144 VDD1.n105 7.3702
R2000 VDD1.n53 VDD1.n17 6.59444
R2001 VDD1.n53 VDD1.n52 6.59444
R2002 VDD1.n141 VDD1.n140 6.59444
R2003 VDD1.n141 VDD1.n105 6.59444
R2004 VDD1.n57 VDD1.n56 5.81868
R2005 VDD1.n49 VDD1.n19 5.81868
R2006 VDD1.n137 VDD1.n107 5.81868
R2007 VDD1.n145 VDD1.n144 5.81868
R2008 VDD1.n60 VDD1.n15 5.04292
R2009 VDD1.n48 VDD1.n21 5.04292
R2010 VDD1.n136 VDD1.n109 5.04292
R2011 VDD1.n148 VDD1.n103 5.04292
R2012 VDD1.n61 VDD1.n13 4.26717
R2013 VDD1.n45 VDD1.n44 4.26717
R2014 VDD1.n133 VDD1.n132 4.26717
R2015 VDD1.n149 VDD1.n101 4.26717
R2016 VDD1.n31 VDD1.n30 3.70982
R2017 VDD1.n119 VDD1.n118 3.70982
R2018 VDD1.n88 VDD1.n0 3.49141
R2019 VDD1.n65 VDD1.n64 3.49141
R2020 VDD1.n41 VDD1.n23 3.49141
R2021 VDD1.n129 VDD1.n111 3.49141
R2022 VDD1.n153 VDD1.n152 3.49141
R2023 VDD1.n177 VDD1.n89 3.49141
R2024 VDD1.n86 VDD1.n85 2.71565
R2025 VDD1.n68 VDD1.n11 2.71565
R2026 VDD1.n40 VDD1.n25 2.71565
R2027 VDD1.n128 VDD1.n113 2.71565
R2028 VDD1.n156 VDD1.n99 2.71565
R2029 VDD1.n175 VDD1.n174 2.71565
R2030 VDD1.n180 VDD1.t1 2.02196
R2031 VDD1.n180 VDD1.t2 2.02196
R2032 VDD1.n178 VDD1.t4 2.02196
R2033 VDD1.n178 VDD1.t5 2.02196
R2034 VDD1.n82 VDD1.n2 1.93989
R2035 VDD1.n69 VDD1.n9 1.93989
R2036 VDD1.n37 VDD1.n36 1.93989
R2037 VDD1.n125 VDD1.n124 1.93989
R2038 VDD1.n157 VDD1.n97 1.93989
R2039 VDD1.n171 VDD1.n91 1.93989
R2040 VDD1.n81 VDD1.n4 1.16414
R2041 VDD1.n73 VDD1.n72 1.16414
R2042 VDD1.n33 VDD1.n27 1.16414
R2043 VDD1.n121 VDD1.n115 1.16414
R2044 VDD1.n162 VDD1.n160 1.16414
R2045 VDD1.n170 VDD1.n93 1.16414
R2046 VDD1 VDD1.n181 0.502655
R2047 VDD1.n78 VDD1.n77 0.388379
R2048 VDD1.n8 VDD1.n6 0.388379
R2049 VDD1.n32 VDD1.n29 0.388379
R2050 VDD1.n120 VDD1.n117 0.388379
R2051 VDD1.n161 VDD1.n95 0.388379
R2052 VDD1.n167 VDD1.n166 0.388379
R2053 VDD1.n87 VDD1.n1 0.155672
R2054 VDD1.n80 VDD1.n1 0.155672
R2055 VDD1.n80 VDD1.n79 0.155672
R2056 VDD1.n79 VDD1.n5 0.155672
R2057 VDD1.n71 VDD1.n5 0.155672
R2058 VDD1.n71 VDD1.n70 0.155672
R2059 VDD1.n70 VDD1.n10 0.155672
R2060 VDD1.n63 VDD1.n10 0.155672
R2061 VDD1.n63 VDD1.n62 0.155672
R2062 VDD1.n62 VDD1.n14 0.155672
R2063 VDD1.n55 VDD1.n14 0.155672
R2064 VDD1.n55 VDD1.n54 0.155672
R2065 VDD1.n54 VDD1.n18 0.155672
R2066 VDD1.n47 VDD1.n18 0.155672
R2067 VDD1.n47 VDD1.n46 0.155672
R2068 VDD1.n46 VDD1.n22 0.155672
R2069 VDD1.n39 VDD1.n22 0.155672
R2070 VDD1.n39 VDD1.n38 0.155672
R2071 VDD1.n38 VDD1.n26 0.155672
R2072 VDD1.n31 VDD1.n26 0.155672
R2073 VDD1.n119 VDD1.n114 0.155672
R2074 VDD1.n126 VDD1.n114 0.155672
R2075 VDD1.n127 VDD1.n126 0.155672
R2076 VDD1.n127 VDD1.n110 0.155672
R2077 VDD1.n134 VDD1.n110 0.155672
R2078 VDD1.n135 VDD1.n134 0.155672
R2079 VDD1.n135 VDD1.n106 0.155672
R2080 VDD1.n142 VDD1.n106 0.155672
R2081 VDD1.n143 VDD1.n142 0.155672
R2082 VDD1.n143 VDD1.n102 0.155672
R2083 VDD1.n150 VDD1.n102 0.155672
R2084 VDD1.n151 VDD1.n150 0.155672
R2085 VDD1.n151 VDD1.n98 0.155672
R2086 VDD1.n158 VDD1.n98 0.155672
R2087 VDD1.n159 VDD1.n158 0.155672
R2088 VDD1.n159 VDD1.n94 0.155672
R2089 VDD1.n168 VDD1.n94 0.155672
R2090 VDD1.n169 VDD1.n168 0.155672
R2091 VDD1.n169 VDD1.n90 0.155672
R2092 VDD1.n176 VDD1.n90 0.155672
R2093 VN.n3 VN.t3 204.118
R2094 VN.n17 VN.t0 204.118
R2095 VN.n4 VN.t4 170.718
R2096 VN.n12 VN.t5 170.718
R2097 VN.n18 VN.t1 170.718
R2098 VN.n26 VN.t2 170.718
R2099 VN.n25 VN.n14 161.3
R2100 VN.n24 VN.n23 161.3
R2101 VN.n22 VN.n15 161.3
R2102 VN.n21 VN.n20 161.3
R2103 VN.n19 VN.n16 161.3
R2104 VN.n11 VN.n0 161.3
R2105 VN.n10 VN.n9 161.3
R2106 VN.n8 VN.n1 161.3
R2107 VN.n7 VN.n6 161.3
R2108 VN.n5 VN.n2 161.3
R2109 VN.n13 VN.n12 93.694
R2110 VN.n27 VN.n26 93.694
R2111 VN.n4 VN.n3 59.4102
R2112 VN.n18 VN.n17 59.4102
R2113 VN VN.n27 50.8012
R2114 VN.n10 VN.n1 45.4209
R2115 VN.n24 VN.n15 45.4209
R2116 VN.n6 VN.n1 35.7332
R2117 VN.n20 VN.n15 35.7332
R2118 VN.n6 VN.n5 24.5923
R2119 VN.n11 VN.n10 24.5923
R2120 VN.n20 VN.n19 24.5923
R2121 VN.n25 VN.n24 24.5923
R2122 VN.n12 VN.n11 17.2148
R2123 VN.n26 VN.n25 17.2148
R2124 VN.n5 VN.n4 12.2964
R2125 VN.n19 VN.n18 12.2964
R2126 VN.n17 VN.n16 9.22766
R2127 VN.n3 VN.n2 9.22766
R2128 VN.n27 VN.n14 0.278335
R2129 VN.n13 VN.n0 0.278335
R2130 VN.n23 VN.n14 0.189894
R2131 VN.n23 VN.n22 0.189894
R2132 VN.n22 VN.n21 0.189894
R2133 VN.n21 VN.n16 0.189894
R2134 VN.n7 VN.n2 0.189894
R2135 VN.n8 VN.n7 0.189894
R2136 VN.n9 VN.n8 0.189894
R2137 VN.n9 VN.n0 0.189894
R2138 VN VN.n13 0.153485
R2139 VDD2.n175 VDD2.n91 756.745
R2140 VDD2.n84 VDD2.n0 756.745
R2141 VDD2.n176 VDD2.n175 585
R2142 VDD2.n174 VDD2.n173 585
R2143 VDD2.n95 VDD2.n94 585
R2144 VDD2.n168 VDD2.n167 585
R2145 VDD2.n166 VDD2.n97 585
R2146 VDD2.n165 VDD2.n164 585
R2147 VDD2.n100 VDD2.n98 585
R2148 VDD2.n159 VDD2.n158 585
R2149 VDD2.n157 VDD2.n156 585
R2150 VDD2.n104 VDD2.n103 585
R2151 VDD2.n151 VDD2.n150 585
R2152 VDD2.n149 VDD2.n148 585
R2153 VDD2.n108 VDD2.n107 585
R2154 VDD2.n143 VDD2.n142 585
R2155 VDD2.n141 VDD2.n140 585
R2156 VDD2.n112 VDD2.n111 585
R2157 VDD2.n135 VDD2.n134 585
R2158 VDD2.n133 VDD2.n132 585
R2159 VDD2.n116 VDD2.n115 585
R2160 VDD2.n127 VDD2.n126 585
R2161 VDD2.n125 VDD2.n124 585
R2162 VDD2.n120 VDD2.n119 585
R2163 VDD2.n28 VDD2.n27 585
R2164 VDD2.n33 VDD2.n32 585
R2165 VDD2.n35 VDD2.n34 585
R2166 VDD2.n24 VDD2.n23 585
R2167 VDD2.n41 VDD2.n40 585
R2168 VDD2.n43 VDD2.n42 585
R2169 VDD2.n20 VDD2.n19 585
R2170 VDD2.n49 VDD2.n48 585
R2171 VDD2.n51 VDD2.n50 585
R2172 VDD2.n16 VDD2.n15 585
R2173 VDD2.n57 VDD2.n56 585
R2174 VDD2.n59 VDD2.n58 585
R2175 VDD2.n12 VDD2.n11 585
R2176 VDD2.n65 VDD2.n64 585
R2177 VDD2.n67 VDD2.n66 585
R2178 VDD2.n8 VDD2.n7 585
R2179 VDD2.n74 VDD2.n73 585
R2180 VDD2.n75 VDD2.n6 585
R2181 VDD2.n77 VDD2.n76 585
R2182 VDD2.n4 VDD2.n3 585
R2183 VDD2.n83 VDD2.n82 585
R2184 VDD2.n85 VDD2.n84 585
R2185 VDD2.n121 VDD2.t3 327.466
R2186 VDD2.n29 VDD2.t2 327.466
R2187 VDD2.n175 VDD2.n174 171.744
R2188 VDD2.n174 VDD2.n94 171.744
R2189 VDD2.n167 VDD2.n94 171.744
R2190 VDD2.n167 VDD2.n166 171.744
R2191 VDD2.n166 VDD2.n165 171.744
R2192 VDD2.n165 VDD2.n98 171.744
R2193 VDD2.n158 VDD2.n98 171.744
R2194 VDD2.n158 VDD2.n157 171.744
R2195 VDD2.n157 VDD2.n103 171.744
R2196 VDD2.n150 VDD2.n103 171.744
R2197 VDD2.n150 VDD2.n149 171.744
R2198 VDD2.n149 VDD2.n107 171.744
R2199 VDD2.n142 VDD2.n107 171.744
R2200 VDD2.n142 VDD2.n141 171.744
R2201 VDD2.n141 VDD2.n111 171.744
R2202 VDD2.n134 VDD2.n111 171.744
R2203 VDD2.n134 VDD2.n133 171.744
R2204 VDD2.n133 VDD2.n115 171.744
R2205 VDD2.n126 VDD2.n115 171.744
R2206 VDD2.n126 VDD2.n125 171.744
R2207 VDD2.n125 VDD2.n119 171.744
R2208 VDD2.n33 VDD2.n27 171.744
R2209 VDD2.n34 VDD2.n33 171.744
R2210 VDD2.n34 VDD2.n23 171.744
R2211 VDD2.n41 VDD2.n23 171.744
R2212 VDD2.n42 VDD2.n41 171.744
R2213 VDD2.n42 VDD2.n19 171.744
R2214 VDD2.n49 VDD2.n19 171.744
R2215 VDD2.n50 VDD2.n49 171.744
R2216 VDD2.n50 VDD2.n15 171.744
R2217 VDD2.n57 VDD2.n15 171.744
R2218 VDD2.n58 VDD2.n57 171.744
R2219 VDD2.n58 VDD2.n11 171.744
R2220 VDD2.n65 VDD2.n11 171.744
R2221 VDD2.n66 VDD2.n65 171.744
R2222 VDD2.n66 VDD2.n7 171.744
R2223 VDD2.n74 VDD2.n7 171.744
R2224 VDD2.n75 VDD2.n74 171.744
R2225 VDD2.n76 VDD2.n75 171.744
R2226 VDD2.n76 VDD2.n3 171.744
R2227 VDD2.n83 VDD2.n3 171.744
R2228 VDD2.n84 VDD2.n83 171.744
R2229 VDD2.t3 VDD2.n119 85.8723
R2230 VDD2.t2 VDD2.n27 85.8723
R2231 VDD2.n90 VDD2.n89 70.3069
R2232 VDD2 VDD2.n181 70.3041
R2233 VDD2.n90 VDD2.n88 50.4898
R2234 VDD2.n180 VDD2.n179 48.8641
R2235 VDD2.n180 VDD2.n90 44.8618
R2236 VDD2.n121 VDD2.n120 16.3895
R2237 VDD2.n29 VDD2.n28 16.3895
R2238 VDD2.n168 VDD2.n97 13.1884
R2239 VDD2.n77 VDD2.n6 13.1884
R2240 VDD2.n169 VDD2.n95 12.8005
R2241 VDD2.n164 VDD2.n99 12.8005
R2242 VDD2.n124 VDD2.n123 12.8005
R2243 VDD2.n32 VDD2.n31 12.8005
R2244 VDD2.n73 VDD2.n72 12.8005
R2245 VDD2.n78 VDD2.n4 12.8005
R2246 VDD2.n173 VDD2.n172 12.0247
R2247 VDD2.n163 VDD2.n100 12.0247
R2248 VDD2.n127 VDD2.n118 12.0247
R2249 VDD2.n35 VDD2.n26 12.0247
R2250 VDD2.n71 VDD2.n8 12.0247
R2251 VDD2.n82 VDD2.n81 12.0247
R2252 VDD2.n176 VDD2.n93 11.249
R2253 VDD2.n160 VDD2.n159 11.249
R2254 VDD2.n128 VDD2.n116 11.249
R2255 VDD2.n36 VDD2.n24 11.249
R2256 VDD2.n68 VDD2.n67 11.249
R2257 VDD2.n85 VDD2.n2 11.249
R2258 VDD2.n177 VDD2.n91 10.4732
R2259 VDD2.n156 VDD2.n102 10.4732
R2260 VDD2.n132 VDD2.n131 10.4732
R2261 VDD2.n40 VDD2.n39 10.4732
R2262 VDD2.n64 VDD2.n10 10.4732
R2263 VDD2.n86 VDD2.n0 10.4732
R2264 VDD2.n155 VDD2.n104 9.69747
R2265 VDD2.n135 VDD2.n114 9.69747
R2266 VDD2.n43 VDD2.n22 9.69747
R2267 VDD2.n63 VDD2.n12 9.69747
R2268 VDD2.n179 VDD2.n178 9.45567
R2269 VDD2.n88 VDD2.n87 9.45567
R2270 VDD2.n147 VDD2.n146 9.3005
R2271 VDD2.n106 VDD2.n105 9.3005
R2272 VDD2.n153 VDD2.n152 9.3005
R2273 VDD2.n155 VDD2.n154 9.3005
R2274 VDD2.n102 VDD2.n101 9.3005
R2275 VDD2.n161 VDD2.n160 9.3005
R2276 VDD2.n163 VDD2.n162 9.3005
R2277 VDD2.n99 VDD2.n96 9.3005
R2278 VDD2.n178 VDD2.n177 9.3005
R2279 VDD2.n93 VDD2.n92 9.3005
R2280 VDD2.n172 VDD2.n171 9.3005
R2281 VDD2.n170 VDD2.n169 9.3005
R2282 VDD2.n145 VDD2.n144 9.3005
R2283 VDD2.n110 VDD2.n109 9.3005
R2284 VDD2.n139 VDD2.n138 9.3005
R2285 VDD2.n137 VDD2.n136 9.3005
R2286 VDD2.n114 VDD2.n113 9.3005
R2287 VDD2.n131 VDD2.n130 9.3005
R2288 VDD2.n129 VDD2.n128 9.3005
R2289 VDD2.n118 VDD2.n117 9.3005
R2290 VDD2.n123 VDD2.n122 9.3005
R2291 VDD2.n87 VDD2.n86 9.3005
R2292 VDD2.n2 VDD2.n1 9.3005
R2293 VDD2.n81 VDD2.n80 9.3005
R2294 VDD2.n79 VDD2.n78 9.3005
R2295 VDD2.n18 VDD2.n17 9.3005
R2296 VDD2.n47 VDD2.n46 9.3005
R2297 VDD2.n45 VDD2.n44 9.3005
R2298 VDD2.n22 VDD2.n21 9.3005
R2299 VDD2.n39 VDD2.n38 9.3005
R2300 VDD2.n37 VDD2.n36 9.3005
R2301 VDD2.n26 VDD2.n25 9.3005
R2302 VDD2.n31 VDD2.n30 9.3005
R2303 VDD2.n53 VDD2.n52 9.3005
R2304 VDD2.n55 VDD2.n54 9.3005
R2305 VDD2.n14 VDD2.n13 9.3005
R2306 VDD2.n61 VDD2.n60 9.3005
R2307 VDD2.n63 VDD2.n62 9.3005
R2308 VDD2.n10 VDD2.n9 9.3005
R2309 VDD2.n69 VDD2.n68 9.3005
R2310 VDD2.n71 VDD2.n70 9.3005
R2311 VDD2.n72 VDD2.n5 9.3005
R2312 VDD2.n152 VDD2.n151 8.92171
R2313 VDD2.n136 VDD2.n112 8.92171
R2314 VDD2.n44 VDD2.n20 8.92171
R2315 VDD2.n60 VDD2.n59 8.92171
R2316 VDD2.n148 VDD2.n106 8.14595
R2317 VDD2.n140 VDD2.n139 8.14595
R2318 VDD2.n48 VDD2.n47 8.14595
R2319 VDD2.n56 VDD2.n14 8.14595
R2320 VDD2.n147 VDD2.n108 7.3702
R2321 VDD2.n143 VDD2.n110 7.3702
R2322 VDD2.n51 VDD2.n18 7.3702
R2323 VDD2.n55 VDD2.n16 7.3702
R2324 VDD2.n144 VDD2.n108 6.59444
R2325 VDD2.n144 VDD2.n143 6.59444
R2326 VDD2.n52 VDD2.n51 6.59444
R2327 VDD2.n52 VDD2.n16 6.59444
R2328 VDD2.n148 VDD2.n147 5.81868
R2329 VDD2.n140 VDD2.n110 5.81868
R2330 VDD2.n48 VDD2.n18 5.81868
R2331 VDD2.n56 VDD2.n55 5.81868
R2332 VDD2.n151 VDD2.n106 5.04292
R2333 VDD2.n139 VDD2.n112 5.04292
R2334 VDD2.n47 VDD2.n20 5.04292
R2335 VDD2.n59 VDD2.n14 5.04292
R2336 VDD2.n152 VDD2.n104 4.26717
R2337 VDD2.n136 VDD2.n135 4.26717
R2338 VDD2.n44 VDD2.n43 4.26717
R2339 VDD2.n60 VDD2.n12 4.26717
R2340 VDD2.n122 VDD2.n121 3.70982
R2341 VDD2.n30 VDD2.n29 3.70982
R2342 VDD2.n179 VDD2.n91 3.49141
R2343 VDD2.n156 VDD2.n155 3.49141
R2344 VDD2.n132 VDD2.n114 3.49141
R2345 VDD2.n40 VDD2.n22 3.49141
R2346 VDD2.n64 VDD2.n63 3.49141
R2347 VDD2.n88 VDD2.n0 3.49141
R2348 VDD2.n177 VDD2.n176 2.71565
R2349 VDD2.n159 VDD2.n102 2.71565
R2350 VDD2.n131 VDD2.n116 2.71565
R2351 VDD2.n39 VDD2.n24 2.71565
R2352 VDD2.n67 VDD2.n10 2.71565
R2353 VDD2.n86 VDD2.n85 2.71565
R2354 VDD2.n181 VDD2.t4 2.02196
R2355 VDD2.n181 VDD2.t5 2.02196
R2356 VDD2.n89 VDD2.t1 2.02196
R2357 VDD2.n89 VDD2.t0 2.02196
R2358 VDD2.n173 VDD2.n93 1.93989
R2359 VDD2.n160 VDD2.n100 1.93989
R2360 VDD2.n128 VDD2.n127 1.93989
R2361 VDD2.n36 VDD2.n35 1.93989
R2362 VDD2.n68 VDD2.n8 1.93989
R2363 VDD2.n82 VDD2.n2 1.93989
R2364 VDD2 VDD2.n180 1.73972
R2365 VDD2.n172 VDD2.n95 1.16414
R2366 VDD2.n164 VDD2.n163 1.16414
R2367 VDD2.n124 VDD2.n118 1.16414
R2368 VDD2.n32 VDD2.n26 1.16414
R2369 VDD2.n73 VDD2.n71 1.16414
R2370 VDD2.n81 VDD2.n4 1.16414
R2371 VDD2.n169 VDD2.n168 0.388379
R2372 VDD2.n99 VDD2.n97 0.388379
R2373 VDD2.n123 VDD2.n120 0.388379
R2374 VDD2.n31 VDD2.n28 0.388379
R2375 VDD2.n72 VDD2.n6 0.388379
R2376 VDD2.n78 VDD2.n77 0.388379
R2377 VDD2.n178 VDD2.n92 0.155672
R2378 VDD2.n171 VDD2.n92 0.155672
R2379 VDD2.n171 VDD2.n170 0.155672
R2380 VDD2.n170 VDD2.n96 0.155672
R2381 VDD2.n162 VDD2.n96 0.155672
R2382 VDD2.n162 VDD2.n161 0.155672
R2383 VDD2.n161 VDD2.n101 0.155672
R2384 VDD2.n154 VDD2.n101 0.155672
R2385 VDD2.n154 VDD2.n153 0.155672
R2386 VDD2.n153 VDD2.n105 0.155672
R2387 VDD2.n146 VDD2.n105 0.155672
R2388 VDD2.n146 VDD2.n145 0.155672
R2389 VDD2.n145 VDD2.n109 0.155672
R2390 VDD2.n138 VDD2.n109 0.155672
R2391 VDD2.n138 VDD2.n137 0.155672
R2392 VDD2.n137 VDD2.n113 0.155672
R2393 VDD2.n130 VDD2.n113 0.155672
R2394 VDD2.n130 VDD2.n129 0.155672
R2395 VDD2.n129 VDD2.n117 0.155672
R2396 VDD2.n122 VDD2.n117 0.155672
R2397 VDD2.n30 VDD2.n25 0.155672
R2398 VDD2.n37 VDD2.n25 0.155672
R2399 VDD2.n38 VDD2.n37 0.155672
R2400 VDD2.n38 VDD2.n21 0.155672
R2401 VDD2.n45 VDD2.n21 0.155672
R2402 VDD2.n46 VDD2.n45 0.155672
R2403 VDD2.n46 VDD2.n17 0.155672
R2404 VDD2.n53 VDD2.n17 0.155672
R2405 VDD2.n54 VDD2.n53 0.155672
R2406 VDD2.n54 VDD2.n13 0.155672
R2407 VDD2.n61 VDD2.n13 0.155672
R2408 VDD2.n62 VDD2.n61 0.155672
R2409 VDD2.n62 VDD2.n9 0.155672
R2410 VDD2.n69 VDD2.n9 0.155672
R2411 VDD2.n70 VDD2.n69 0.155672
R2412 VDD2.n70 VDD2.n5 0.155672
R2413 VDD2.n79 VDD2.n5 0.155672
R2414 VDD2.n80 VDD2.n79 0.155672
R2415 VDD2.n80 VDD2.n1 0.155672
R2416 VDD2.n87 VDD2.n1 0.155672
C0 B VDD1 2.32579f
C1 VDD2 VTAIL 9.30855f
C2 VP VDD1 8.91797f
C3 B VDD2 2.39196f
C4 VDD1 VN 0.150486f
C5 VP VDD2 0.430916f
C6 VDD2 VN 8.64162f
C7 VDD1 w_n3050_n4184# 2.49459f
C8 B VTAIL 4.44665f
C9 VDD2 w_n3050_n4184# 2.56915f
C10 VP VTAIL 8.559719f
C11 B VP 1.80408f
C12 VN VTAIL 8.54533f
C13 B VN 1.14892f
C14 VP VN 7.35622f
C15 VTAIL w_n3050_n4184# 3.52187f
C16 B w_n3050_n4184# 10.3639f
C17 VDD1 VDD2 1.27808f
C18 VP w_n3050_n4184# 6.16163f
C19 VN w_n3050_n4184# 5.76823f
C20 VDD1 VTAIL 9.26139f
C21 VDD2 VSUBS 1.946069f
C22 VDD1 VSUBS 1.833141f
C23 VTAIL VSUBS 1.275657f
C24 VN VSUBS 5.70674f
C25 VP VSUBS 2.831116f
C26 B VSUBS 4.654815f
C27 w_n3050_n4184# VSUBS 0.156319p
C28 VDD2.n0 VSUBS 0.028372f
C29 VDD2.n1 VSUBS 0.027183f
C30 VDD2.n2 VSUBS 0.014607f
C31 VDD2.n3 VSUBS 0.034525f
C32 VDD2.n4 VSUBS 0.015466f
C33 VDD2.n5 VSUBS 0.027183f
C34 VDD2.n6 VSUBS 0.015037f
C35 VDD2.n7 VSUBS 0.034525f
C36 VDD2.n8 VSUBS 0.015466f
C37 VDD2.n9 VSUBS 0.027183f
C38 VDD2.n10 VSUBS 0.014607f
C39 VDD2.n11 VSUBS 0.034525f
C40 VDD2.n12 VSUBS 0.015466f
C41 VDD2.n13 VSUBS 0.027183f
C42 VDD2.n14 VSUBS 0.014607f
C43 VDD2.n15 VSUBS 0.034525f
C44 VDD2.n16 VSUBS 0.015466f
C45 VDD2.n17 VSUBS 0.027183f
C46 VDD2.n18 VSUBS 0.014607f
C47 VDD2.n19 VSUBS 0.034525f
C48 VDD2.n20 VSUBS 0.015466f
C49 VDD2.n21 VSUBS 0.027183f
C50 VDD2.n22 VSUBS 0.014607f
C51 VDD2.n23 VSUBS 0.034525f
C52 VDD2.n24 VSUBS 0.015466f
C53 VDD2.n25 VSUBS 0.027183f
C54 VDD2.n26 VSUBS 0.014607f
C55 VDD2.n27 VSUBS 0.025894f
C56 VDD2.n28 VSUBS 0.021963f
C57 VDD2.t2 VSUBS 0.073985f
C58 VDD2.n29 VSUBS 0.200276f
C59 VDD2.n30 VSUBS 1.86896f
C60 VDD2.n31 VSUBS 0.014607f
C61 VDD2.n32 VSUBS 0.015466f
C62 VDD2.n33 VSUBS 0.034525f
C63 VDD2.n34 VSUBS 0.034525f
C64 VDD2.n35 VSUBS 0.015466f
C65 VDD2.n36 VSUBS 0.014607f
C66 VDD2.n37 VSUBS 0.027183f
C67 VDD2.n38 VSUBS 0.027183f
C68 VDD2.n39 VSUBS 0.014607f
C69 VDD2.n40 VSUBS 0.015466f
C70 VDD2.n41 VSUBS 0.034525f
C71 VDD2.n42 VSUBS 0.034525f
C72 VDD2.n43 VSUBS 0.015466f
C73 VDD2.n44 VSUBS 0.014607f
C74 VDD2.n45 VSUBS 0.027183f
C75 VDD2.n46 VSUBS 0.027183f
C76 VDD2.n47 VSUBS 0.014607f
C77 VDD2.n48 VSUBS 0.015466f
C78 VDD2.n49 VSUBS 0.034525f
C79 VDD2.n50 VSUBS 0.034525f
C80 VDD2.n51 VSUBS 0.015466f
C81 VDD2.n52 VSUBS 0.014607f
C82 VDD2.n53 VSUBS 0.027183f
C83 VDD2.n54 VSUBS 0.027183f
C84 VDD2.n55 VSUBS 0.014607f
C85 VDD2.n56 VSUBS 0.015466f
C86 VDD2.n57 VSUBS 0.034525f
C87 VDD2.n58 VSUBS 0.034525f
C88 VDD2.n59 VSUBS 0.015466f
C89 VDD2.n60 VSUBS 0.014607f
C90 VDD2.n61 VSUBS 0.027183f
C91 VDD2.n62 VSUBS 0.027183f
C92 VDD2.n63 VSUBS 0.014607f
C93 VDD2.n64 VSUBS 0.015466f
C94 VDD2.n65 VSUBS 0.034525f
C95 VDD2.n66 VSUBS 0.034525f
C96 VDD2.n67 VSUBS 0.015466f
C97 VDD2.n68 VSUBS 0.014607f
C98 VDD2.n69 VSUBS 0.027183f
C99 VDD2.n70 VSUBS 0.027183f
C100 VDD2.n71 VSUBS 0.014607f
C101 VDD2.n72 VSUBS 0.014607f
C102 VDD2.n73 VSUBS 0.015466f
C103 VDD2.n74 VSUBS 0.034525f
C104 VDD2.n75 VSUBS 0.034525f
C105 VDD2.n76 VSUBS 0.034525f
C106 VDD2.n77 VSUBS 0.015037f
C107 VDD2.n78 VSUBS 0.014607f
C108 VDD2.n79 VSUBS 0.027183f
C109 VDD2.n80 VSUBS 0.027183f
C110 VDD2.n81 VSUBS 0.014607f
C111 VDD2.n82 VSUBS 0.015466f
C112 VDD2.n83 VSUBS 0.034525f
C113 VDD2.n84 VSUBS 0.078485f
C114 VDD2.n85 VSUBS 0.015466f
C115 VDD2.n86 VSUBS 0.014607f
C116 VDD2.n87 VSUBS 0.062832f
C117 VDD2.n88 VSUBS 0.064295f
C118 VDD2.t1 VSUBS 0.345411f
C119 VDD2.t0 VSUBS 0.345411f
C120 VDD2.n89 VSUBS 2.83382f
C121 VDD2.n90 VSUBS 3.3343f
C122 VDD2.n91 VSUBS 0.028372f
C123 VDD2.n92 VSUBS 0.027183f
C124 VDD2.n93 VSUBS 0.014607f
C125 VDD2.n94 VSUBS 0.034525f
C126 VDD2.n95 VSUBS 0.015466f
C127 VDD2.n96 VSUBS 0.027183f
C128 VDD2.n97 VSUBS 0.015037f
C129 VDD2.n98 VSUBS 0.034525f
C130 VDD2.n99 VSUBS 0.014607f
C131 VDD2.n100 VSUBS 0.015466f
C132 VDD2.n101 VSUBS 0.027183f
C133 VDD2.n102 VSUBS 0.014607f
C134 VDD2.n103 VSUBS 0.034525f
C135 VDD2.n104 VSUBS 0.015466f
C136 VDD2.n105 VSUBS 0.027183f
C137 VDD2.n106 VSUBS 0.014607f
C138 VDD2.n107 VSUBS 0.034525f
C139 VDD2.n108 VSUBS 0.015466f
C140 VDD2.n109 VSUBS 0.027183f
C141 VDD2.n110 VSUBS 0.014607f
C142 VDD2.n111 VSUBS 0.034525f
C143 VDD2.n112 VSUBS 0.015466f
C144 VDD2.n113 VSUBS 0.027183f
C145 VDD2.n114 VSUBS 0.014607f
C146 VDD2.n115 VSUBS 0.034525f
C147 VDD2.n116 VSUBS 0.015466f
C148 VDD2.n117 VSUBS 0.027183f
C149 VDD2.n118 VSUBS 0.014607f
C150 VDD2.n119 VSUBS 0.025894f
C151 VDD2.n120 VSUBS 0.021963f
C152 VDD2.t3 VSUBS 0.073985f
C153 VDD2.n121 VSUBS 0.200275f
C154 VDD2.n122 VSUBS 1.86896f
C155 VDD2.n123 VSUBS 0.014607f
C156 VDD2.n124 VSUBS 0.015466f
C157 VDD2.n125 VSUBS 0.034525f
C158 VDD2.n126 VSUBS 0.034525f
C159 VDD2.n127 VSUBS 0.015466f
C160 VDD2.n128 VSUBS 0.014607f
C161 VDD2.n129 VSUBS 0.027183f
C162 VDD2.n130 VSUBS 0.027183f
C163 VDD2.n131 VSUBS 0.014607f
C164 VDD2.n132 VSUBS 0.015466f
C165 VDD2.n133 VSUBS 0.034525f
C166 VDD2.n134 VSUBS 0.034525f
C167 VDD2.n135 VSUBS 0.015466f
C168 VDD2.n136 VSUBS 0.014607f
C169 VDD2.n137 VSUBS 0.027183f
C170 VDD2.n138 VSUBS 0.027183f
C171 VDD2.n139 VSUBS 0.014607f
C172 VDD2.n140 VSUBS 0.015466f
C173 VDD2.n141 VSUBS 0.034525f
C174 VDD2.n142 VSUBS 0.034525f
C175 VDD2.n143 VSUBS 0.015466f
C176 VDD2.n144 VSUBS 0.014607f
C177 VDD2.n145 VSUBS 0.027183f
C178 VDD2.n146 VSUBS 0.027183f
C179 VDD2.n147 VSUBS 0.014607f
C180 VDD2.n148 VSUBS 0.015466f
C181 VDD2.n149 VSUBS 0.034525f
C182 VDD2.n150 VSUBS 0.034525f
C183 VDD2.n151 VSUBS 0.015466f
C184 VDD2.n152 VSUBS 0.014607f
C185 VDD2.n153 VSUBS 0.027183f
C186 VDD2.n154 VSUBS 0.027183f
C187 VDD2.n155 VSUBS 0.014607f
C188 VDD2.n156 VSUBS 0.015466f
C189 VDD2.n157 VSUBS 0.034525f
C190 VDD2.n158 VSUBS 0.034525f
C191 VDD2.n159 VSUBS 0.015466f
C192 VDD2.n160 VSUBS 0.014607f
C193 VDD2.n161 VSUBS 0.027183f
C194 VDD2.n162 VSUBS 0.027183f
C195 VDD2.n163 VSUBS 0.014607f
C196 VDD2.n164 VSUBS 0.015466f
C197 VDD2.n165 VSUBS 0.034525f
C198 VDD2.n166 VSUBS 0.034525f
C199 VDD2.n167 VSUBS 0.034525f
C200 VDD2.n168 VSUBS 0.015037f
C201 VDD2.n169 VSUBS 0.014607f
C202 VDD2.n170 VSUBS 0.027183f
C203 VDD2.n171 VSUBS 0.027183f
C204 VDD2.n172 VSUBS 0.014607f
C205 VDD2.n173 VSUBS 0.015466f
C206 VDD2.n174 VSUBS 0.034525f
C207 VDD2.n175 VSUBS 0.078485f
C208 VDD2.n176 VSUBS 0.015466f
C209 VDD2.n177 VSUBS 0.014607f
C210 VDD2.n178 VSUBS 0.062832f
C211 VDD2.n179 VSUBS 0.058013f
C212 VDD2.n180 VSUBS 3.02767f
C213 VDD2.t4 VSUBS 0.345411f
C214 VDD2.t5 VSUBS 0.345411f
C215 VDD2.n181 VSUBS 2.83378f
C216 VN.n0 VSUBS 0.040095f
C217 VN.t5 VSUBS 3.04664f
C218 VN.n1 VSUBS 0.025547f
C219 VN.n2 VSUBS 0.26096f
C220 VN.t4 VSUBS 3.04664f
C221 VN.t3 VSUBS 3.2486f
C222 VN.n3 VSUBS 1.12945f
C223 VN.n4 VSUBS 1.14436f
C224 VN.n5 VSUBS 0.042478f
C225 VN.n6 VSUBS 0.061087f
C226 VN.n7 VSUBS 0.030413f
C227 VN.n8 VSUBS 0.030413f
C228 VN.n9 VSUBS 0.030413f
C229 VN.n10 VSUBS 0.058186f
C230 VN.n11 VSUBS 0.048046f
C231 VN.n12 VSUBS 1.1649f
C232 VN.n13 VSUBS 0.04081f
C233 VN.n14 VSUBS 0.040095f
C234 VN.t2 VSUBS 3.04664f
C235 VN.n15 VSUBS 0.025547f
C236 VN.n16 VSUBS 0.26096f
C237 VN.t1 VSUBS 3.04664f
C238 VN.t0 VSUBS 3.2486f
C239 VN.n17 VSUBS 1.12945f
C240 VN.n18 VSUBS 1.14436f
C241 VN.n19 VSUBS 0.042478f
C242 VN.n20 VSUBS 0.061087f
C243 VN.n21 VSUBS 0.030413f
C244 VN.n22 VSUBS 0.030413f
C245 VN.n23 VSUBS 0.030413f
C246 VN.n24 VSUBS 0.058186f
C247 VN.n25 VSUBS 0.048046f
C248 VN.n26 VSUBS 1.1649f
C249 VN.n27 VSUBS 1.72586f
C250 VDD1.n0 VSUBS 0.028371f
C251 VDD1.n1 VSUBS 0.027183f
C252 VDD1.n2 VSUBS 0.014607f
C253 VDD1.n3 VSUBS 0.034525f
C254 VDD1.n4 VSUBS 0.015466f
C255 VDD1.n5 VSUBS 0.027183f
C256 VDD1.n6 VSUBS 0.015036f
C257 VDD1.n7 VSUBS 0.034525f
C258 VDD1.n8 VSUBS 0.014607f
C259 VDD1.n9 VSUBS 0.015466f
C260 VDD1.n10 VSUBS 0.027183f
C261 VDD1.n11 VSUBS 0.014607f
C262 VDD1.n12 VSUBS 0.034525f
C263 VDD1.n13 VSUBS 0.015466f
C264 VDD1.n14 VSUBS 0.027183f
C265 VDD1.n15 VSUBS 0.014607f
C266 VDD1.n16 VSUBS 0.034525f
C267 VDD1.n17 VSUBS 0.015466f
C268 VDD1.n18 VSUBS 0.027183f
C269 VDD1.n19 VSUBS 0.014607f
C270 VDD1.n20 VSUBS 0.034525f
C271 VDD1.n21 VSUBS 0.015466f
C272 VDD1.n22 VSUBS 0.027183f
C273 VDD1.n23 VSUBS 0.014607f
C274 VDD1.n24 VSUBS 0.034525f
C275 VDD1.n25 VSUBS 0.015466f
C276 VDD1.n26 VSUBS 0.027183f
C277 VDD1.n27 VSUBS 0.014607f
C278 VDD1.n28 VSUBS 0.025894f
C279 VDD1.n29 VSUBS 0.021963f
C280 VDD1.t3 VSUBS 0.073984f
C281 VDD1.n30 VSUBS 0.200272f
C282 VDD1.n31 VSUBS 1.86893f
C283 VDD1.n32 VSUBS 0.014607f
C284 VDD1.n33 VSUBS 0.015466f
C285 VDD1.n34 VSUBS 0.034525f
C286 VDD1.n35 VSUBS 0.034525f
C287 VDD1.n36 VSUBS 0.015466f
C288 VDD1.n37 VSUBS 0.014607f
C289 VDD1.n38 VSUBS 0.027183f
C290 VDD1.n39 VSUBS 0.027183f
C291 VDD1.n40 VSUBS 0.014607f
C292 VDD1.n41 VSUBS 0.015466f
C293 VDD1.n42 VSUBS 0.034525f
C294 VDD1.n43 VSUBS 0.034525f
C295 VDD1.n44 VSUBS 0.015466f
C296 VDD1.n45 VSUBS 0.014607f
C297 VDD1.n46 VSUBS 0.027183f
C298 VDD1.n47 VSUBS 0.027183f
C299 VDD1.n48 VSUBS 0.014607f
C300 VDD1.n49 VSUBS 0.015466f
C301 VDD1.n50 VSUBS 0.034525f
C302 VDD1.n51 VSUBS 0.034525f
C303 VDD1.n52 VSUBS 0.015466f
C304 VDD1.n53 VSUBS 0.014607f
C305 VDD1.n54 VSUBS 0.027183f
C306 VDD1.n55 VSUBS 0.027183f
C307 VDD1.n56 VSUBS 0.014607f
C308 VDD1.n57 VSUBS 0.015466f
C309 VDD1.n58 VSUBS 0.034525f
C310 VDD1.n59 VSUBS 0.034525f
C311 VDD1.n60 VSUBS 0.015466f
C312 VDD1.n61 VSUBS 0.014607f
C313 VDD1.n62 VSUBS 0.027183f
C314 VDD1.n63 VSUBS 0.027183f
C315 VDD1.n64 VSUBS 0.014607f
C316 VDD1.n65 VSUBS 0.015466f
C317 VDD1.n66 VSUBS 0.034525f
C318 VDD1.n67 VSUBS 0.034525f
C319 VDD1.n68 VSUBS 0.015466f
C320 VDD1.n69 VSUBS 0.014607f
C321 VDD1.n70 VSUBS 0.027183f
C322 VDD1.n71 VSUBS 0.027183f
C323 VDD1.n72 VSUBS 0.014607f
C324 VDD1.n73 VSUBS 0.015466f
C325 VDD1.n74 VSUBS 0.034525f
C326 VDD1.n75 VSUBS 0.034525f
C327 VDD1.n76 VSUBS 0.034525f
C328 VDD1.n77 VSUBS 0.015036f
C329 VDD1.n78 VSUBS 0.014607f
C330 VDD1.n79 VSUBS 0.027183f
C331 VDD1.n80 VSUBS 0.027183f
C332 VDD1.n81 VSUBS 0.014607f
C333 VDD1.n82 VSUBS 0.015466f
C334 VDD1.n83 VSUBS 0.034525f
C335 VDD1.n84 VSUBS 0.078484f
C336 VDD1.n85 VSUBS 0.015466f
C337 VDD1.n86 VSUBS 0.014607f
C338 VDD1.n87 VSUBS 0.062831f
C339 VDD1.n88 VSUBS 0.065046f
C340 VDD1.n89 VSUBS 0.028371f
C341 VDD1.n90 VSUBS 0.027183f
C342 VDD1.n91 VSUBS 0.014607f
C343 VDD1.n92 VSUBS 0.034525f
C344 VDD1.n93 VSUBS 0.015466f
C345 VDD1.n94 VSUBS 0.027183f
C346 VDD1.n95 VSUBS 0.015036f
C347 VDD1.n96 VSUBS 0.034525f
C348 VDD1.n97 VSUBS 0.015466f
C349 VDD1.n98 VSUBS 0.027183f
C350 VDD1.n99 VSUBS 0.014607f
C351 VDD1.n100 VSUBS 0.034525f
C352 VDD1.n101 VSUBS 0.015466f
C353 VDD1.n102 VSUBS 0.027183f
C354 VDD1.n103 VSUBS 0.014607f
C355 VDD1.n104 VSUBS 0.034525f
C356 VDD1.n105 VSUBS 0.015466f
C357 VDD1.n106 VSUBS 0.027183f
C358 VDD1.n107 VSUBS 0.014607f
C359 VDD1.n108 VSUBS 0.034525f
C360 VDD1.n109 VSUBS 0.015466f
C361 VDD1.n110 VSUBS 0.027183f
C362 VDD1.n111 VSUBS 0.014607f
C363 VDD1.n112 VSUBS 0.034525f
C364 VDD1.n113 VSUBS 0.015466f
C365 VDD1.n114 VSUBS 0.027183f
C366 VDD1.n115 VSUBS 0.014607f
C367 VDD1.n116 VSUBS 0.025894f
C368 VDD1.n117 VSUBS 0.021963f
C369 VDD1.t0 VSUBS 0.073984f
C370 VDD1.n118 VSUBS 0.200272f
C371 VDD1.n119 VSUBS 1.86893f
C372 VDD1.n120 VSUBS 0.014607f
C373 VDD1.n121 VSUBS 0.015466f
C374 VDD1.n122 VSUBS 0.034525f
C375 VDD1.n123 VSUBS 0.034525f
C376 VDD1.n124 VSUBS 0.015466f
C377 VDD1.n125 VSUBS 0.014607f
C378 VDD1.n126 VSUBS 0.027183f
C379 VDD1.n127 VSUBS 0.027183f
C380 VDD1.n128 VSUBS 0.014607f
C381 VDD1.n129 VSUBS 0.015466f
C382 VDD1.n130 VSUBS 0.034525f
C383 VDD1.n131 VSUBS 0.034525f
C384 VDD1.n132 VSUBS 0.015466f
C385 VDD1.n133 VSUBS 0.014607f
C386 VDD1.n134 VSUBS 0.027183f
C387 VDD1.n135 VSUBS 0.027183f
C388 VDD1.n136 VSUBS 0.014607f
C389 VDD1.n137 VSUBS 0.015466f
C390 VDD1.n138 VSUBS 0.034525f
C391 VDD1.n139 VSUBS 0.034525f
C392 VDD1.n140 VSUBS 0.015466f
C393 VDD1.n141 VSUBS 0.014607f
C394 VDD1.n142 VSUBS 0.027183f
C395 VDD1.n143 VSUBS 0.027183f
C396 VDD1.n144 VSUBS 0.014607f
C397 VDD1.n145 VSUBS 0.015466f
C398 VDD1.n146 VSUBS 0.034525f
C399 VDD1.n147 VSUBS 0.034525f
C400 VDD1.n148 VSUBS 0.015466f
C401 VDD1.n149 VSUBS 0.014607f
C402 VDD1.n150 VSUBS 0.027183f
C403 VDD1.n151 VSUBS 0.027183f
C404 VDD1.n152 VSUBS 0.014607f
C405 VDD1.n153 VSUBS 0.015466f
C406 VDD1.n154 VSUBS 0.034525f
C407 VDD1.n155 VSUBS 0.034525f
C408 VDD1.n156 VSUBS 0.015466f
C409 VDD1.n157 VSUBS 0.014607f
C410 VDD1.n158 VSUBS 0.027183f
C411 VDD1.n159 VSUBS 0.027183f
C412 VDD1.n160 VSUBS 0.014607f
C413 VDD1.n161 VSUBS 0.014607f
C414 VDD1.n162 VSUBS 0.015466f
C415 VDD1.n163 VSUBS 0.034525f
C416 VDD1.n164 VSUBS 0.034525f
C417 VDD1.n165 VSUBS 0.034525f
C418 VDD1.n166 VSUBS 0.015036f
C419 VDD1.n167 VSUBS 0.014607f
C420 VDD1.n168 VSUBS 0.027183f
C421 VDD1.n169 VSUBS 0.027183f
C422 VDD1.n170 VSUBS 0.014607f
C423 VDD1.n171 VSUBS 0.015466f
C424 VDD1.n172 VSUBS 0.034525f
C425 VDD1.n173 VSUBS 0.078484f
C426 VDD1.n174 VSUBS 0.015466f
C427 VDD1.n175 VSUBS 0.014607f
C428 VDD1.n176 VSUBS 0.062831f
C429 VDD1.n177 VSUBS 0.064294f
C430 VDD1.t4 VSUBS 0.345405f
C431 VDD1.t5 VSUBS 0.345405f
C432 VDD1.n178 VSUBS 2.83377f
C433 VDD1.n179 VSUBS 3.46276f
C434 VDD1.t1 VSUBS 0.345405f
C435 VDD1.t2 VSUBS 0.345405f
C436 VDD1.n180 VSUBS 2.82817f
C437 VDD1.n181 VSUBS 3.57366f
C438 VTAIL.t2 VSUBS 0.352512f
C439 VTAIL.t1 VSUBS 0.352512f
C440 VTAIL.n0 VSUBS 2.71896f
C441 VTAIL.n1 VSUBS 0.865595f
C442 VTAIL.n2 VSUBS 0.028955f
C443 VTAIL.n3 VSUBS 0.027742f
C444 VTAIL.n4 VSUBS 0.014907f
C445 VTAIL.n5 VSUBS 0.035235f
C446 VTAIL.n6 VSUBS 0.015784f
C447 VTAIL.n7 VSUBS 0.027742f
C448 VTAIL.n8 VSUBS 0.015346f
C449 VTAIL.n9 VSUBS 0.035235f
C450 VTAIL.n10 VSUBS 0.015784f
C451 VTAIL.n11 VSUBS 0.027742f
C452 VTAIL.n12 VSUBS 0.014907f
C453 VTAIL.n13 VSUBS 0.035235f
C454 VTAIL.n14 VSUBS 0.015784f
C455 VTAIL.n15 VSUBS 0.027742f
C456 VTAIL.n16 VSUBS 0.014907f
C457 VTAIL.n17 VSUBS 0.035235f
C458 VTAIL.n18 VSUBS 0.015784f
C459 VTAIL.n19 VSUBS 0.027742f
C460 VTAIL.n20 VSUBS 0.014907f
C461 VTAIL.n21 VSUBS 0.035235f
C462 VTAIL.n22 VSUBS 0.015784f
C463 VTAIL.n23 VSUBS 0.027742f
C464 VTAIL.n24 VSUBS 0.014907f
C465 VTAIL.n25 VSUBS 0.035235f
C466 VTAIL.n26 VSUBS 0.015784f
C467 VTAIL.n27 VSUBS 0.027742f
C468 VTAIL.n28 VSUBS 0.014907f
C469 VTAIL.n29 VSUBS 0.026426f
C470 VTAIL.n30 VSUBS 0.022415f
C471 VTAIL.t6 VSUBS 0.075506f
C472 VTAIL.n31 VSUBS 0.204393f
C473 VTAIL.n32 VSUBS 1.90738f
C474 VTAIL.n33 VSUBS 0.014907f
C475 VTAIL.n34 VSUBS 0.015784f
C476 VTAIL.n35 VSUBS 0.035235f
C477 VTAIL.n36 VSUBS 0.035235f
C478 VTAIL.n37 VSUBS 0.015784f
C479 VTAIL.n38 VSUBS 0.014907f
C480 VTAIL.n39 VSUBS 0.027742f
C481 VTAIL.n40 VSUBS 0.027742f
C482 VTAIL.n41 VSUBS 0.014907f
C483 VTAIL.n42 VSUBS 0.015784f
C484 VTAIL.n43 VSUBS 0.035235f
C485 VTAIL.n44 VSUBS 0.035235f
C486 VTAIL.n45 VSUBS 0.015784f
C487 VTAIL.n46 VSUBS 0.014907f
C488 VTAIL.n47 VSUBS 0.027742f
C489 VTAIL.n48 VSUBS 0.027742f
C490 VTAIL.n49 VSUBS 0.014907f
C491 VTAIL.n50 VSUBS 0.015784f
C492 VTAIL.n51 VSUBS 0.035235f
C493 VTAIL.n52 VSUBS 0.035235f
C494 VTAIL.n53 VSUBS 0.015784f
C495 VTAIL.n54 VSUBS 0.014907f
C496 VTAIL.n55 VSUBS 0.027742f
C497 VTAIL.n56 VSUBS 0.027742f
C498 VTAIL.n57 VSUBS 0.014907f
C499 VTAIL.n58 VSUBS 0.015784f
C500 VTAIL.n59 VSUBS 0.035235f
C501 VTAIL.n60 VSUBS 0.035235f
C502 VTAIL.n61 VSUBS 0.015784f
C503 VTAIL.n62 VSUBS 0.014907f
C504 VTAIL.n63 VSUBS 0.027742f
C505 VTAIL.n64 VSUBS 0.027742f
C506 VTAIL.n65 VSUBS 0.014907f
C507 VTAIL.n66 VSUBS 0.015784f
C508 VTAIL.n67 VSUBS 0.035235f
C509 VTAIL.n68 VSUBS 0.035235f
C510 VTAIL.n69 VSUBS 0.015784f
C511 VTAIL.n70 VSUBS 0.014907f
C512 VTAIL.n71 VSUBS 0.027742f
C513 VTAIL.n72 VSUBS 0.027742f
C514 VTAIL.n73 VSUBS 0.014907f
C515 VTAIL.n74 VSUBS 0.014907f
C516 VTAIL.n75 VSUBS 0.015784f
C517 VTAIL.n76 VSUBS 0.035235f
C518 VTAIL.n77 VSUBS 0.035235f
C519 VTAIL.n78 VSUBS 0.035235f
C520 VTAIL.n79 VSUBS 0.015346f
C521 VTAIL.n80 VSUBS 0.014907f
C522 VTAIL.n81 VSUBS 0.027742f
C523 VTAIL.n82 VSUBS 0.027742f
C524 VTAIL.n83 VSUBS 0.014907f
C525 VTAIL.n84 VSUBS 0.015784f
C526 VTAIL.n85 VSUBS 0.035235f
C527 VTAIL.n86 VSUBS 0.080099f
C528 VTAIL.n87 VSUBS 0.015784f
C529 VTAIL.n88 VSUBS 0.014907f
C530 VTAIL.n89 VSUBS 0.064124f
C531 VTAIL.n90 VSUBS 0.04005f
C532 VTAIL.n91 VSUBS 0.366228f
C533 VTAIL.t9 VSUBS 0.352512f
C534 VTAIL.t11 VSUBS 0.352512f
C535 VTAIL.n92 VSUBS 2.71896f
C536 VTAIL.n93 VSUBS 2.88517f
C537 VTAIL.t3 VSUBS 0.352512f
C538 VTAIL.t5 VSUBS 0.352512f
C539 VTAIL.n94 VSUBS 2.71898f
C540 VTAIL.n95 VSUBS 2.88515f
C541 VTAIL.n96 VSUBS 0.028955f
C542 VTAIL.n97 VSUBS 0.027742f
C543 VTAIL.n98 VSUBS 0.014907f
C544 VTAIL.n99 VSUBS 0.035235f
C545 VTAIL.n100 VSUBS 0.015784f
C546 VTAIL.n101 VSUBS 0.027742f
C547 VTAIL.n102 VSUBS 0.015346f
C548 VTAIL.n103 VSUBS 0.035235f
C549 VTAIL.n104 VSUBS 0.014907f
C550 VTAIL.n105 VSUBS 0.015784f
C551 VTAIL.n106 VSUBS 0.027742f
C552 VTAIL.n107 VSUBS 0.014907f
C553 VTAIL.n108 VSUBS 0.035235f
C554 VTAIL.n109 VSUBS 0.015784f
C555 VTAIL.n110 VSUBS 0.027742f
C556 VTAIL.n111 VSUBS 0.014907f
C557 VTAIL.n112 VSUBS 0.035235f
C558 VTAIL.n113 VSUBS 0.015784f
C559 VTAIL.n114 VSUBS 0.027742f
C560 VTAIL.n115 VSUBS 0.014907f
C561 VTAIL.n116 VSUBS 0.035235f
C562 VTAIL.n117 VSUBS 0.015784f
C563 VTAIL.n118 VSUBS 0.027742f
C564 VTAIL.n119 VSUBS 0.014907f
C565 VTAIL.n120 VSUBS 0.035235f
C566 VTAIL.n121 VSUBS 0.015784f
C567 VTAIL.n122 VSUBS 0.027742f
C568 VTAIL.n123 VSUBS 0.014907f
C569 VTAIL.n124 VSUBS 0.026426f
C570 VTAIL.n125 VSUBS 0.022415f
C571 VTAIL.t0 VSUBS 0.075506f
C572 VTAIL.n126 VSUBS 0.204393f
C573 VTAIL.n127 VSUBS 1.90738f
C574 VTAIL.n128 VSUBS 0.014907f
C575 VTAIL.n129 VSUBS 0.015784f
C576 VTAIL.n130 VSUBS 0.035235f
C577 VTAIL.n131 VSUBS 0.035235f
C578 VTAIL.n132 VSUBS 0.015784f
C579 VTAIL.n133 VSUBS 0.014907f
C580 VTAIL.n134 VSUBS 0.027742f
C581 VTAIL.n135 VSUBS 0.027742f
C582 VTAIL.n136 VSUBS 0.014907f
C583 VTAIL.n137 VSUBS 0.015784f
C584 VTAIL.n138 VSUBS 0.035235f
C585 VTAIL.n139 VSUBS 0.035235f
C586 VTAIL.n140 VSUBS 0.015784f
C587 VTAIL.n141 VSUBS 0.014907f
C588 VTAIL.n142 VSUBS 0.027742f
C589 VTAIL.n143 VSUBS 0.027742f
C590 VTAIL.n144 VSUBS 0.014907f
C591 VTAIL.n145 VSUBS 0.015784f
C592 VTAIL.n146 VSUBS 0.035235f
C593 VTAIL.n147 VSUBS 0.035235f
C594 VTAIL.n148 VSUBS 0.015784f
C595 VTAIL.n149 VSUBS 0.014907f
C596 VTAIL.n150 VSUBS 0.027742f
C597 VTAIL.n151 VSUBS 0.027742f
C598 VTAIL.n152 VSUBS 0.014907f
C599 VTAIL.n153 VSUBS 0.015784f
C600 VTAIL.n154 VSUBS 0.035235f
C601 VTAIL.n155 VSUBS 0.035235f
C602 VTAIL.n156 VSUBS 0.015784f
C603 VTAIL.n157 VSUBS 0.014907f
C604 VTAIL.n158 VSUBS 0.027742f
C605 VTAIL.n159 VSUBS 0.027742f
C606 VTAIL.n160 VSUBS 0.014907f
C607 VTAIL.n161 VSUBS 0.015784f
C608 VTAIL.n162 VSUBS 0.035235f
C609 VTAIL.n163 VSUBS 0.035235f
C610 VTAIL.n164 VSUBS 0.015784f
C611 VTAIL.n165 VSUBS 0.014907f
C612 VTAIL.n166 VSUBS 0.027742f
C613 VTAIL.n167 VSUBS 0.027742f
C614 VTAIL.n168 VSUBS 0.014907f
C615 VTAIL.n169 VSUBS 0.015784f
C616 VTAIL.n170 VSUBS 0.035235f
C617 VTAIL.n171 VSUBS 0.035235f
C618 VTAIL.n172 VSUBS 0.035235f
C619 VTAIL.n173 VSUBS 0.015346f
C620 VTAIL.n174 VSUBS 0.014907f
C621 VTAIL.n175 VSUBS 0.027742f
C622 VTAIL.n176 VSUBS 0.027742f
C623 VTAIL.n177 VSUBS 0.014907f
C624 VTAIL.n178 VSUBS 0.015784f
C625 VTAIL.n179 VSUBS 0.035235f
C626 VTAIL.n180 VSUBS 0.080099f
C627 VTAIL.n181 VSUBS 0.015784f
C628 VTAIL.n182 VSUBS 0.014907f
C629 VTAIL.n183 VSUBS 0.064124f
C630 VTAIL.n184 VSUBS 0.04005f
C631 VTAIL.n185 VSUBS 0.366228f
C632 VTAIL.t10 VSUBS 0.352512f
C633 VTAIL.t8 VSUBS 0.352512f
C634 VTAIL.n186 VSUBS 2.71898f
C635 VTAIL.n187 VSUBS 1.01064f
C636 VTAIL.n188 VSUBS 0.028955f
C637 VTAIL.n189 VSUBS 0.027742f
C638 VTAIL.n190 VSUBS 0.014907f
C639 VTAIL.n191 VSUBS 0.035235f
C640 VTAIL.n192 VSUBS 0.015784f
C641 VTAIL.n193 VSUBS 0.027742f
C642 VTAIL.n194 VSUBS 0.015346f
C643 VTAIL.n195 VSUBS 0.035235f
C644 VTAIL.n196 VSUBS 0.014907f
C645 VTAIL.n197 VSUBS 0.015784f
C646 VTAIL.n198 VSUBS 0.027742f
C647 VTAIL.n199 VSUBS 0.014907f
C648 VTAIL.n200 VSUBS 0.035235f
C649 VTAIL.n201 VSUBS 0.015784f
C650 VTAIL.n202 VSUBS 0.027742f
C651 VTAIL.n203 VSUBS 0.014907f
C652 VTAIL.n204 VSUBS 0.035235f
C653 VTAIL.n205 VSUBS 0.015784f
C654 VTAIL.n206 VSUBS 0.027742f
C655 VTAIL.n207 VSUBS 0.014907f
C656 VTAIL.n208 VSUBS 0.035235f
C657 VTAIL.n209 VSUBS 0.015784f
C658 VTAIL.n210 VSUBS 0.027742f
C659 VTAIL.n211 VSUBS 0.014907f
C660 VTAIL.n212 VSUBS 0.035235f
C661 VTAIL.n213 VSUBS 0.015784f
C662 VTAIL.n214 VSUBS 0.027742f
C663 VTAIL.n215 VSUBS 0.014907f
C664 VTAIL.n216 VSUBS 0.026426f
C665 VTAIL.n217 VSUBS 0.022415f
C666 VTAIL.t7 VSUBS 0.075506f
C667 VTAIL.n218 VSUBS 0.204393f
C668 VTAIL.n219 VSUBS 1.90738f
C669 VTAIL.n220 VSUBS 0.014907f
C670 VTAIL.n221 VSUBS 0.015784f
C671 VTAIL.n222 VSUBS 0.035235f
C672 VTAIL.n223 VSUBS 0.035235f
C673 VTAIL.n224 VSUBS 0.015784f
C674 VTAIL.n225 VSUBS 0.014907f
C675 VTAIL.n226 VSUBS 0.027742f
C676 VTAIL.n227 VSUBS 0.027742f
C677 VTAIL.n228 VSUBS 0.014907f
C678 VTAIL.n229 VSUBS 0.015784f
C679 VTAIL.n230 VSUBS 0.035235f
C680 VTAIL.n231 VSUBS 0.035235f
C681 VTAIL.n232 VSUBS 0.015784f
C682 VTAIL.n233 VSUBS 0.014907f
C683 VTAIL.n234 VSUBS 0.027742f
C684 VTAIL.n235 VSUBS 0.027742f
C685 VTAIL.n236 VSUBS 0.014907f
C686 VTAIL.n237 VSUBS 0.015784f
C687 VTAIL.n238 VSUBS 0.035235f
C688 VTAIL.n239 VSUBS 0.035235f
C689 VTAIL.n240 VSUBS 0.015784f
C690 VTAIL.n241 VSUBS 0.014907f
C691 VTAIL.n242 VSUBS 0.027742f
C692 VTAIL.n243 VSUBS 0.027742f
C693 VTAIL.n244 VSUBS 0.014907f
C694 VTAIL.n245 VSUBS 0.015784f
C695 VTAIL.n246 VSUBS 0.035235f
C696 VTAIL.n247 VSUBS 0.035235f
C697 VTAIL.n248 VSUBS 0.015784f
C698 VTAIL.n249 VSUBS 0.014907f
C699 VTAIL.n250 VSUBS 0.027742f
C700 VTAIL.n251 VSUBS 0.027742f
C701 VTAIL.n252 VSUBS 0.014907f
C702 VTAIL.n253 VSUBS 0.015784f
C703 VTAIL.n254 VSUBS 0.035235f
C704 VTAIL.n255 VSUBS 0.035235f
C705 VTAIL.n256 VSUBS 0.015784f
C706 VTAIL.n257 VSUBS 0.014907f
C707 VTAIL.n258 VSUBS 0.027742f
C708 VTAIL.n259 VSUBS 0.027742f
C709 VTAIL.n260 VSUBS 0.014907f
C710 VTAIL.n261 VSUBS 0.015784f
C711 VTAIL.n262 VSUBS 0.035235f
C712 VTAIL.n263 VSUBS 0.035235f
C713 VTAIL.n264 VSUBS 0.035235f
C714 VTAIL.n265 VSUBS 0.015346f
C715 VTAIL.n266 VSUBS 0.014907f
C716 VTAIL.n267 VSUBS 0.027742f
C717 VTAIL.n268 VSUBS 0.027742f
C718 VTAIL.n269 VSUBS 0.014907f
C719 VTAIL.n270 VSUBS 0.015784f
C720 VTAIL.n271 VSUBS 0.035235f
C721 VTAIL.n272 VSUBS 0.080099f
C722 VTAIL.n273 VSUBS 0.015784f
C723 VTAIL.n274 VSUBS 0.014907f
C724 VTAIL.n275 VSUBS 0.064124f
C725 VTAIL.n276 VSUBS 0.04005f
C726 VTAIL.n277 VSUBS 2.04038f
C727 VTAIL.n278 VSUBS 0.028955f
C728 VTAIL.n279 VSUBS 0.027742f
C729 VTAIL.n280 VSUBS 0.014907f
C730 VTAIL.n281 VSUBS 0.035235f
C731 VTAIL.n282 VSUBS 0.015784f
C732 VTAIL.n283 VSUBS 0.027742f
C733 VTAIL.n284 VSUBS 0.015346f
C734 VTAIL.n285 VSUBS 0.035235f
C735 VTAIL.n286 VSUBS 0.015784f
C736 VTAIL.n287 VSUBS 0.027742f
C737 VTAIL.n288 VSUBS 0.014907f
C738 VTAIL.n289 VSUBS 0.035235f
C739 VTAIL.n290 VSUBS 0.015784f
C740 VTAIL.n291 VSUBS 0.027742f
C741 VTAIL.n292 VSUBS 0.014907f
C742 VTAIL.n293 VSUBS 0.035235f
C743 VTAIL.n294 VSUBS 0.015784f
C744 VTAIL.n295 VSUBS 0.027742f
C745 VTAIL.n296 VSUBS 0.014907f
C746 VTAIL.n297 VSUBS 0.035235f
C747 VTAIL.n298 VSUBS 0.015784f
C748 VTAIL.n299 VSUBS 0.027742f
C749 VTAIL.n300 VSUBS 0.014907f
C750 VTAIL.n301 VSUBS 0.035235f
C751 VTAIL.n302 VSUBS 0.015784f
C752 VTAIL.n303 VSUBS 0.027742f
C753 VTAIL.n304 VSUBS 0.014907f
C754 VTAIL.n305 VSUBS 0.026426f
C755 VTAIL.n306 VSUBS 0.022415f
C756 VTAIL.t4 VSUBS 0.075506f
C757 VTAIL.n307 VSUBS 0.204393f
C758 VTAIL.n308 VSUBS 1.90738f
C759 VTAIL.n309 VSUBS 0.014907f
C760 VTAIL.n310 VSUBS 0.015784f
C761 VTAIL.n311 VSUBS 0.035235f
C762 VTAIL.n312 VSUBS 0.035235f
C763 VTAIL.n313 VSUBS 0.015784f
C764 VTAIL.n314 VSUBS 0.014907f
C765 VTAIL.n315 VSUBS 0.027742f
C766 VTAIL.n316 VSUBS 0.027742f
C767 VTAIL.n317 VSUBS 0.014907f
C768 VTAIL.n318 VSUBS 0.015784f
C769 VTAIL.n319 VSUBS 0.035235f
C770 VTAIL.n320 VSUBS 0.035235f
C771 VTAIL.n321 VSUBS 0.015784f
C772 VTAIL.n322 VSUBS 0.014907f
C773 VTAIL.n323 VSUBS 0.027742f
C774 VTAIL.n324 VSUBS 0.027742f
C775 VTAIL.n325 VSUBS 0.014907f
C776 VTAIL.n326 VSUBS 0.015784f
C777 VTAIL.n327 VSUBS 0.035235f
C778 VTAIL.n328 VSUBS 0.035235f
C779 VTAIL.n329 VSUBS 0.015784f
C780 VTAIL.n330 VSUBS 0.014907f
C781 VTAIL.n331 VSUBS 0.027742f
C782 VTAIL.n332 VSUBS 0.027742f
C783 VTAIL.n333 VSUBS 0.014907f
C784 VTAIL.n334 VSUBS 0.015784f
C785 VTAIL.n335 VSUBS 0.035235f
C786 VTAIL.n336 VSUBS 0.035235f
C787 VTAIL.n337 VSUBS 0.015784f
C788 VTAIL.n338 VSUBS 0.014907f
C789 VTAIL.n339 VSUBS 0.027742f
C790 VTAIL.n340 VSUBS 0.027742f
C791 VTAIL.n341 VSUBS 0.014907f
C792 VTAIL.n342 VSUBS 0.015784f
C793 VTAIL.n343 VSUBS 0.035235f
C794 VTAIL.n344 VSUBS 0.035235f
C795 VTAIL.n345 VSUBS 0.015784f
C796 VTAIL.n346 VSUBS 0.014907f
C797 VTAIL.n347 VSUBS 0.027742f
C798 VTAIL.n348 VSUBS 0.027742f
C799 VTAIL.n349 VSUBS 0.014907f
C800 VTAIL.n350 VSUBS 0.014907f
C801 VTAIL.n351 VSUBS 0.015784f
C802 VTAIL.n352 VSUBS 0.035235f
C803 VTAIL.n353 VSUBS 0.035235f
C804 VTAIL.n354 VSUBS 0.035235f
C805 VTAIL.n355 VSUBS 0.015346f
C806 VTAIL.n356 VSUBS 0.014907f
C807 VTAIL.n357 VSUBS 0.027742f
C808 VTAIL.n358 VSUBS 0.027742f
C809 VTAIL.n359 VSUBS 0.014907f
C810 VTAIL.n360 VSUBS 0.015784f
C811 VTAIL.n361 VSUBS 0.035235f
C812 VTAIL.n362 VSUBS 0.080099f
C813 VTAIL.n363 VSUBS 0.015784f
C814 VTAIL.n364 VSUBS 0.014907f
C815 VTAIL.n365 VSUBS 0.064124f
C816 VTAIL.n366 VSUBS 0.04005f
C817 VTAIL.n367 VSUBS 1.98509f
C818 VP.n0 VSUBS 0.041212f
C819 VP.t0 VSUBS 3.1315f
C820 VP.n1 VSUBS 0.026259f
C821 VP.n2 VSUBS 0.031261f
C822 VP.t1 VSUBS 3.1315f
C823 VP.n3 VSUBS 0.062788f
C824 VP.n4 VSUBS 0.031261f
C825 VP.t5 VSUBS 3.1315f
C826 VP.n5 VSUBS 1.19734f
C827 VP.n6 VSUBS 0.041212f
C828 VP.t3 VSUBS 3.1315f
C829 VP.n7 VSUBS 0.026259f
C830 VP.n8 VSUBS 0.268229f
C831 VP.t4 VSUBS 3.1315f
C832 VP.t2 VSUBS 3.33908f
C833 VP.n9 VSUBS 1.16091f
C834 VP.n10 VSUBS 1.17623f
C835 VP.n11 VSUBS 0.043661f
C836 VP.n12 VSUBS 0.062788f
C837 VP.n13 VSUBS 0.031261f
C838 VP.n14 VSUBS 0.031261f
C839 VP.n15 VSUBS 0.031261f
C840 VP.n16 VSUBS 0.059807f
C841 VP.n17 VSUBS 0.049384f
C842 VP.n18 VSUBS 1.19734f
C843 VP.n19 VSUBS 1.75716f
C844 VP.n20 VSUBS 1.77947f
C845 VP.n21 VSUBS 0.041212f
C846 VP.n22 VSUBS 0.049384f
C847 VP.n23 VSUBS 0.059807f
C848 VP.n24 VSUBS 0.026259f
C849 VP.n25 VSUBS 0.031261f
C850 VP.n26 VSUBS 0.031261f
C851 VP.n27 VSUBS 0.031261f
C852 VP.n28 VSUBS 0.043661f
C853 VP.n29 VSUBS 1.09455f
C854 VP.n30 VSUBS 0.043661f
C855 VP.n31 VSUBS 0.062788f
C856 VP.n32 VSUBS 0.031261f
C857 VP.n33 VSUBS 0.031261f
C858 VP.n34 VSUBS 0.031261f
C859 VP.n35 VSUBS 0.059807f
C860 VP.n36 VSUBS 0.049384f
C861 VP.n37 VSUBS 1.19734f
C862 VP.n38 VSUBS 0.041946f
C863 B.n0 VSUBS 0.00671f
C864 B.n1 VSUBS 0.00671f
C865 B.n2 VSUBS 0.009923f
C866 B.n3 VSUBS 0.007604f
C867 B.n4 VSUBS 0.007604f
C868 B.n5 VSUBS 0.007604f
C869 B.n6 VSUBS 0.007604f
C870 B.n7 VSUBS 0.007604f
C871 B.n8 VSUBS 0.007604f
C872 B.n9 VSUBS 0.007604f
C873 B.n10 VSUBS 0.007604f
C874 B.n11 VSUBS 0.007604f
C875 B.n12 VSUBS 0.007604f
C876 B.n13 VSUBS 0.007604f
C877 B.n14 VSUBS 0.007604f
C878 B.n15 VSUBS 0.007604f
C879 B.n16 VSUBS 0.007604f
C880 B.n17 VSUBS 0.007604f
C881 B.n18 VSUBS 0.007604f
C882 B.n19 VSUBS 0.007604f
C883 B.n20 VSUBS 0.007604f
C884 B.n21 VSUBS 0.018746f
C885 B.n22 VSUBS 0.007604f
C886 B.n23 VSUBS 0.007604f
C887 B.n24 VSUBS 0.007604f
C888 B.n25 VSUBS 0.007604f
C889 B.n26 VSUBS 0.007604f
C890 B.n27 VSUBS 0.007604f
C891 B.n28 VSUBS 0.007604f
C892 B.n29 VSUBS 0.007604f
C893 B.n30 VSUBS 0.007604f
C894 B.n31 VSUBS 0.007604f
C895 B.n32 VSUBS 0.007604f
C896 B.n33 VSUBS 0.007604f
C897 B.n34 VSUBS 0.007604f
C898 B.n35 VSUBS 0.007604f
C899 B.n36 VSUBS 0.007604f
C900 B.n37 VSUBS 0.007604f
C901 B.n38 VSUBS 0.007604f
C902 B.n39 VSUBS 0.007604f
C903 B.n40 VSUBS 0.007604f
C904 B.n41 VSUBS 0.007604f
C905 B.n42 VSUBS 0.007604f
C906 B.n43 VSUBS 0.007604f
C907 B.n44 VSUBS 0.007604f
C908 B.n45 VSUBS 0.007604f
C909 B.n46 VSUBS 0.007604f
C910 B.n47 VSUBS 0.007604f
C911 B.t7 VSUBS 0.331294f
C912 B.t8 VSUBS 0.363546f
C913 B.t6 VSUBS 1.7546f
C914 B.n48 VSUBS 0.553132f
C915 B.n49 VSUBS 0.330293f
C916 B.n50 VSUBS 0.017619f
C917 B.n51 VSUBS 0.007604f
C918 B.n52 VSUBS 0.007604f
C919 B.n53 VSUBS 0.007604f
C920 B.n54 VSUBS 0.007604f
C921 B.n55 VSUBS 0.007604f
C922 B.t4 VSUBS 0.331298f
C923 B.t5 VSUBS 0.363549f
C924 B.t3 VSUBS 1.7546f
C925 B.n56 VSUBS 0.553128f
C926 B.n57 VSUBS 0.330289f
C927 B.n58 VSUBS 0.007604f
C928 B.n59 VSUBS 0.007604f
C929 B.n60 VSUBS 0.007604f
C930 B.n61 VSUBS 0.007604f
C931 B.n62 VSUBS 0.007604f
C932 B.n63 VSUBS 0.007604f
C933 B.n64 VSUBS 0.007604f
C934 B.n65 VSUBS 0.007604f
C935 B.n66 VSUBS 0.007604f
C936 B.n67 VSUBS 0.007604f
C937 B.n68 VSUBS 0.007604f
C938 B.n69 VSUBS 0.007604f
C939 B.n70 VSUBS 0.007604f
C940 B.n71 VSUBS 0.007604f
C941 B.n72 VSUBS 0.007604f
C942 B.n73 VSUBS 0.007604f
C943 B.n74 VSUBS 0.007604f
C944 B.n75 VSUBS 0.007604f
C945 B.n76 VSUBS 0.007604f
C946 B.n77 VSUBS 0.007604f
C947 B.n78 VSUBS 0.007604f
C948 B.n79 VSUBS 0.007604f
C949 B.n80 VSUBS 0.007604f
C950 B.n81 VSUBS 0.007604f
C951 B.n82 VSUBS 0.007604f
C952 B.n83 VSUBS 0.007604f
C953 B.n84 VSUBS 0.017487f
C954 B.n85 VSUBS 0.007604f
C955 B.n86 VSUBS 0.007604f
C956 B.n87 VSUBS 0.007604f
C957 B.n88 VSUBS 0.007604f
C958 B.n89 VSUBS 0.007604f
C959 B.n90 VSUBS 0.007604f
C960 B.n91 VSUBS 0.007604f
C961 B.n92 VSUBS 0.007604f
C962 B.n93 VSUBS 0.007604f
C963 B.n94 VSUBS 0.007604f
C964 B.n95 VSUBS 0.007604f
C965 B.n96 VSUBS 0.007604f
C966 B.n97 VSUBS 0.007604f
C967 B.n98 VSUBS 0.007604f
C968 B.n99 VSUBS 0.007604f
C969 B.n100 VSUBS 0.007604f
C970 B.n101 VSUBS 0.007604f
C971 B.n102 VSUBS 0.007604f
C972 B.n103 VSUBS 0.007604f
C973 B.n104 VSUBS 0.007604f
C974 B.n105 VSUBS 0.007604f
C975 B.n106 VSUBS 0.007604f
C976 B.n107 VSUBS 0.007604f
C977 B.n108 VSUBS 0.007604f
C978 B.n109 VSUBS 0.007604f
C979 B.n110 VSUBS 0.007604f
C980 B.n111 VSUBS 0.007604f
C981 B.n112 VSUBS 0.007604f
C982 B.n113 VSUBS 0.007604f
C983 B.n114 VSUBS 0.007604f
C984 B.n115 VSUBS 0.007604f
C985 B.n116 VSUBS 0.007604f
C986 B.n117 VSUBS 0.007604f
C987 B.n118 VSUBS 0.007604f
C988 B.n119 VSUBS 0.007604f
C989 B.n120 VSUBS 0.007604f
C990 B.n121 VSUBS 0.007604f
C991 B.n122 VSUBS 0.007604f
C992 B.n123 VSUBS 0.018746f
C993 B.n124 VSUBS 0.007604f
C994 B.n125 VSUBS 0.007604f
C995 B.n126 VSUBS 0.007604f
C996 B.n127 VSUBS 0.007604f
C997 B.n128 VSUBS 0.007604f
C998 B.n129 VSUBS 0.007604f
C999 B.n130 VSUBS 0.007604f
C1000 B.n131 VSUBS 0.007604f
C1001 B.n132 VSUBS 0.007604f
C1002 B.n133 VSUBS 0.007604f
C1003 B.n134 VSUBS 0.007604f
C1004 B.n135 VSUBS 0.007604f
C1005 B.n136 VSUBS 0.007604f
C1006 B.n137 VSUBS 0.007604f
C1007 B.n138 VSUBS 0.007604f
C1008 B.n139 VSUBS 0.007604f
C1009 B.n140 VSUBS 0.007604f
C1010 B.n141 VSUBS 0.007604f
C1011 B.n142 VSUBS 0.007604f
C1012 B.n143 VSUBS 0.007604f
C1013 B.n144 VSUBS 0.007604f
C1014 B.n145 VSUBS 0.007604f
C1015 B.n146 VSUBS 0.007604f
C1016 B.n147 VSUBS 0.007604f
C1017 B.n148 VSUBS 0.007604f
C1018 B.n149 VSUBS 0.007604f
C1019 B.t2 VSUBS 0.331298f
C1020 B.t1 VSUBS 0.363549f
C1021 B.t0 VSUBS 1.7546f
C1022 B.n150 VSUBS 0.553128f
C1023 B.n151 VSUBS 0.330289f
C1024 B.n152 VSUBS 0.017619f
C1025 B.n153 VSUBS 0.007604f
C1026 B.n154 VSUBS 0.007604f
C1027 B.n155 VSUBS 0.007604f
C1028 B.n156 VSUBS 0.007604f
C1029 B.n157 VSUBS 0.007604f
C1030 B.t11 VSUBS 0.331294f
C1031 B.t10 VSUBS 0.363546f
C1032 B.t9 VSUBS 1.7546f
C1033 B.n158 VSUBS 0.553132f
C1034 B.n159 VSUBS 0.330293f
C1035 B.n160 VSUBS 0.007604f
C1036 B.n161 VSUBS 0.007604f
C1037 B.n162 VSUBS 0.007604f
C1038 B.n163 VSUBS 0.007604f
C1039 B.n164 VSUBS 0.007604f
C1040 B.n165 VSUBS 0.007604f
C1041 B.n166 VSUBS 0.007604f
C1042 B.n167 VSUBS 0.007604f
C1043 B.n168 VSUBS 0.007604f
C1044 B.n169 VSUBS 0.007604f
C1045 B.n170 VSUBS 0.007604f
C1046 B.n171 VSUBS 0.007604f
C1047 B.n172 VSUBS 0.007604f
C1048 B.n173 VSUBS 0.007604f
C1049 B.n174 VSUBS 0.007604f
C1050 B.n175 VSUBS 0.007604f
C1051 B.n176 VSUBS 0.007604f
C1052 B.n177 VSUBS 0.007604f
C1053 B.n178 VSUBS 0.007604f
C1054 B.n179 VSUBS 0.007604f
C1055 B.n180 VSUBS 0.007604f
C1056 B.n181 VSUBS 0.007604f
C1057 B.n182 VSUBS 0.007604f
C1058 B.n183 VSUBS 0.007604f
C1059 B.n184 VSUBS 0.007604f
C1060 B.n185 VSUBS 0.007604f
C1061 B.n186 VSUBS 0.017487f
C1062 B.n187 VSUBS 0.007604f
C1063 B.n188 VSUBS 0.007604f
C1064 B.n189 VSUBS 0.007604f
C1065 B.n190 VSUBS 0.007604f
C1066 B.n191 VSUBS 0.007604f
C1067 B.n192 VSUBS 0.007604f
C1068 B.n193 VSUBS 0.007604f
C1069 B.n194 VSUBS 0.007604f
C1070 B.n195 VSUBS 0.007604f
C1071 B.n196 VSUBS 0.007604f
C1072 B.n197 VSUBS 0.007604f
C1073 B.n198 VSUBS 0.007604f
C1074 B.n199 VSUBS 0.007604f
C1075 B.n200 VSUBS 0.007604f
C1076 B.n201 VSUBS 0.007604f
C1077 B.n202 VSUBS 0.007604f
C1078 B.n203 VSUBS 0.007604f
C1079 B.n204 VSUBS 0.007604f
C1080 B.n205 VSUBS 0.007604f
C1081 B.n206 VSUBS 0.007604f
C1082 B.n207 VSUBS 0.007604f
C1083 B.n208 VSUBS 0.007604f
C1084 B.n209 VSUBS 0.007604f
C1085 B.n210 VSUBS 0.007604f
C1086 B.n211 VSUBS 0.007604f
C1087 B.n212 VSUBS 0.007604f
C1088 B.n213 VSUBS 0.007604f
C1089 B.n214 VSUBS 0.007604f
C1090 B.n215 VSUBS 0.007604f
C1091 B.n216 VSUBS 0.007604f
C1092 B.n217 VSUBS 0.007604f
C1093 B.n218 VSUBS 0.007604f
C1094 B.n219 VSUBS 0.007604f
C1095 B.n220 VSUBS 0.007604f
C1096 B.n221 VSUBS 0.007604f
C1097 B.n222 VSUBS 0.007604f
C1098 B.n223 VSUBS 0.007604f
C1099 B.n224 VSUBS 0.007604f
C1100 B.n225 VSUBS 0.007604f
C1101 B.n226 VSUBS 0.007604f
C1102 B.n227 VSUBS 0.007604f
C1103 B.n228 VSUBS 0.007604f
C1104 B.n229 VSUBS 0.007604f
C1105 B.n230 VSUBS 0.007604f
C1106 B.n231 VSUBS 0.007604f
C1107 B.n232 VSUBS 0.007604f
C1108 B.n233 VSUBS 0.007604f
C1109 B.n234 VSUBS 0.007604f
C1110 B.n235 VSUBS 0.007604f
C1111 B.n236 VSUBS 0.007604f
C1112 B.n237 VSUBS 0.007604f
C1113 B.n238 VSUBS 0.007604f
C1114 B.n239 VSUBS 0.007604f
C1115 B.n240 VSUBS 0.007604f
C1116 B.n241 VSUBS 0.007604f
C1117 B.n242 VSUBS 0.007604f
C1118 B.n243 VSUBS 0.007604f
C1119 B.n244 VSUBS 0.007604f
C1120 B.n245 VSUBS 0.007604f
C1121 B.n246 VSUBS 0.007604f
C1122 B.n247 VSUBS 0.007604f
C1123 B.n248 VSUBS 0.007604f
C1124 B.n249 VSUBS 0.007604f
C1125 B.n250 VSUBS 0.007604f
C1126 B.n251 VSUBS 0.007604f
C1127 B.n252 VSUBS 0.007604f
C1128 B.n253 VSUBS 0.007604f
C1129 B.n254 VSUBS 0.007604f
C1130 B.n255 VSUBS 0.007604f
C1131 B.n256 VSUBS 0.007604f
C1132 B.n257 VSUBS 0.007604f
C1133 B.n258 VSUBS 0.007604f
C1134 B.n259 VSUBS 0.017487f
C1135 B.n260 VSUBS 0.018746f
C1136 B.n261 VSUBS 0.018746f
C1137 B.n262 VSUBS 0.007604f
C1138 B.n263 VSUBS 0.007604f
C1139 B.n264 VSUBS 0.007604f
C1140 B.n265 VSUBS 0.007604f
C1141 B.n266 VSUBS 0.007604f
C1142 B.n267 VSUBS 0.007604f
C1143 B.n268 VSUBS 0.007604f
C1144 B.n269 VSUBS 0.007604f
C1145 B.n270 VSUBS 0.007604f
C1146 B.n271 VSUBS 0.007604f
C1147 B.n272 VSUBS 0.007604f
C1148 B.n273 VSUBS 0.007604f
C1149 B.n274 VSUBS 0.007604f
C1150 B.n275 VSUBS 0.007604f
C1151 B.n276 VSUBS 0.007604f
C1152 B.n277 VSUBS 0.007604f
C1153 B.n278 VSUBS 0.007604f
C1154 B.n279 VSUBS 0.007604f
C1155 B.n280 VSUBS 0.007604f
C1156 B.n281 VSUBS 0.007604f
C1157 B.n282 VSUBS 0.007604f
C1158 B.n283 VSUBS 0.007604f
C1159 B.n284 VSUBS 0.007604f
C1160 B.n285 VSUBS 0.007604f
C1161 B.n286 VSUBS 0.007604f
C1162 B.n287 VSUBS 0.007604f
C1163 B.n288 VSUBS 0.007604f
C1164 B.n289 VSUBS 0.007604f
C1165 B.n290 VSUBS 0.007604f
C1166 B.n291 VSUBS 0.007604f
C1167 B.n292 VSUBS 0.007604f
C1168 B.n293 VSUBS 0.007604f
C1169 B.n294 VSUBS 0.007604f
C1170 B.n295 VSUBS 0.007604f
C1171 B.n296 VSUBS 0.007604f
C1172 B.n297 VSUBS 0.007604f
C1173 B.n298 VSUBS 0.007604f
C1174 B.n299 VSUBS 0.007604f
C1175 B.n300 VSUBS 0.007604f
C1176 B.n301 VSUBS 0.007604f
C1177 B.n302 VSUBS 0.007604f
C1178 B.n303 VSUBS 0.007604f
C1179 B.n304 VSUBS 0.007604f
C1180 B.n305 VSUBS 0.007604f
C1181 B.n306 VSUBS 0.007604f
C1182 B.n307 VSUBS 0.007604f
C1183 B.n308 VSUBS 0.007604f
C1184 B.n309 VSUBS 0.007604f
C1185 B.n310 VSUBS 0.007604f
C1186 B.n311 VSUBS 0.007604f
C1187 B.n312 VSUBS 0.007604f
C1188 B.n313 VSUBS 0.007604f
C1189 B.n314 VSUBS 0.007604f
C1190 B.n315 VSUBS 0.007604f
C1191 B.n316 VSUBS 0.007604f
C1192 B.n317 VSUBS 0.007604f
C1193 B.n318 VSUBS 0.007604f
C1194 B.n319 VSUBS 0.007604f
C1195 B.n320 VSUBS 0.007604f
C1196 B.n321 VSUBS 0.007604f
C1197 B.n322 VSUBS 0.007604f
C1198 B.n323 VSUBS 0.007604f
C1199 B.n324 VSUBS 0.007604f
C1200 B.n325 VSUBS 0.007604f
C1201 B.n326 VSUBS 0.007604f
C1202 B.n327 VSUBS 0.007604f
C1203 B.n328 VSUBS 0.007604f
C1204 B.n329 VSUBS 0.007604f
C1205 B.n330 VSUBS 0.007604f
C1206 B.n331 VSUBS 0.007604f
C1207 B.n332 VSUBS 0.007604f
C1208 B.n333 VSUBS 0.007604f
C1209 B.n334 VSUBS 0.007604f
C1210 B.n335 VSUBS 0.007604f
C1211 B.n336 VSUBS 0.007604f
C1212 B.n337 VSUBS 0.007604f
C1213 B.n338 VSUBS 0.007604f
C1214 B.n339 VSUBS 0.007604f
C1215 B.n340 VSUBS 0.005256f
C1216 B.n341 VSUBS 0.017619f
C1217 B.n342 VSUBS 0.006151f
C1218 B.n343 VSUBS 0.007604f
C1219 B.n344 VSUBS 0.007604f
C1220 B.n345 VSUBS 0.007604f
C1221 B.n346 VSUBS 0.007604f
C1222 B.n347 VSUBS 0.007604f
C1223 B.n348 VSUBS 0.007604f
C1224 B.n349 VSUBS 0.007604f
C1225 B.n350 VSUBS 0.007604f
C1226 B.n351 VSUBS 0.007604f
C1227 B.n352 VSUBS 0.007604f
C1228 B.n353 VSUBS 0.007604f
C1229 B.n354 VSUBS 0.006151f
C1230 B.n355 VSUBS 0.007604f
C1231 B.n356 VSUBS 0.007604f
C1232 B.n357 VSUBS 0.005256f
C1233 B.n358 VSUBS 0.007604f
C1234 B.n359 VSUBS 0.007604f
C1235 B.n360 VSUBS 0.007604f
C1236 B.n361 VSUBS 0.007604f
C1237 B.n362 VSUBS 0.007604f
C1238 B.n363 VSUBS 0.007604f
C1239 B.n364 VSUBS 0.007604f
C1240 B.n365 VSUBS 0.007604f
C1241 B.n366 VSUBS 0.007604f
C1242 B.n367 VSUBS 0.007604f
C1243 B.n368 VSUBS 0.007604f
C1244 B.n369 VSUBS 0.007604f
C1245 B.n370 VSUBS 0.007604f
C1246 B.n371 VSUBS 0.007604f
C1247 B.n372 VSUBS 0.007604f
C1248 B.n373 VSUBS 0.007604f
C1249 B.n374 VSUBS 0.007604f
C1250 B.n375 VSUBS 0.007604f
C1251 B.n376 VSUBS 0.007604f
C1252 B.n377 VSUBS 0.007604f
C1253 B.n378 VSUBS 0.007604f
C1254 B.n379 VSUBS 0.007604f
C1255 B.n380 VSUBS 0.007604f
C1256 B.n381 VSUBS 0.007604f
C1257 B.n382 VSUBS 0.007604f
C1258 B.n383 VSUBS 0.007604f
C1259 B.n384 VSUBS 0.007604f
C1260 B.n385 VSUBS 0.007604f
C1261 B.n386 VSUBS 0.007604f
C1262 B.n387 VSUBS 0.007604f
C1263 B.n388 VSUBS 0.007604f
C1264 B.n389 VSUBS 0.007604f
C1265 B.n390 VSUBS 0.007604f
C1266 B.n391 VSUBS 0.007604f
C1267 B.n392 VSUBS 0.007604f
C1268 B.n393 VSUBS 0.007604f
C1269 B.n394 VSUBS 0.007604f
C1270 B.n395 VSUBS 0.007604f
C1271 B.n396 VSUBS 0.007604f
C1272 B.n397 VSUBS 0.007604f
C1273 B.n398 VSUBS 0.007604f
C1274 B.n399 VSUBS 0.007604f
C1275 B.n400 VSUBS 0.007604f
C1276 B.n401 VSUBS 0.007604f
C1277 B.n402 VSUBS 0.007604f
C1278 B.n403 VSUBS 0.007604f
C1279 B.n404 VSUBS 0.007604f
C1280 B.n405 VSUBS 0.007604f
C1281 B.n406 VSUBS 0.007604f
C1282 B.n407 VSUBS 0.007604f
C1283 B.n408 VSUBS 0.007604f
C1284 B.n409 VSUBS 0.007604f
C1285 B.n410 VSUBS 0.007604f
C1286 B.n411 VSUBS 0.007604f
C1287 B.n412 VSUBS 0.007604f
C1288 B.n413 VSUBS 0.007604f
C1289 B.n414 VSUBS 0.007604f
C1290 B.n415 VSUBS 0.007604f
C1291 B.n416 VSUBS 0.007604f
C1292 B.n417 VSUBS 0.007604f
C1293 B.n418 VSUBS 0.007604f
C1294 B.n419 VSUBS 0.007604f
C1295 B.n420 VSUBS 0.007604f
C1296 B.n421 VSUBS 0.007604f
C1297 B.n422 VSUBS 0.007604f
C1298 B.n423 VSUBS 0.007604f
C1299 B.n424 VSUBS 0.007604f
C1300 B.n425 VSUBS 0.007604f
C1301 B.n426 VSUBS 0.007604f
C1302 B.n427 VSUBS 0.007604f
C1303 B.n428 VSUBS 0.007604f
C1304 B.n429 VSUBS 0.007604f
C1305 B.n430 VSUBS 0.007604f
C1306 B.n431 VSUBS 0.007604f
C1307 B.n432 VSUBS 0.007604f
C1308 B.n433 VSUBS 0.007604f
C1309 B.n434 VSUBS 0.007604f
C1310 B.n435 VSUBS 0.007604f
C1311 B.n436 VSUBS 0.017871f
C1312 B.n437 VSUBS 0.018362f
C1313 B.n438 VSUBS 0.017487f
C1314 B.n439 VSUBS 0.007604f
C1315 B.n440 VSUBS 0.007604f
C1316 B.n441 VSUBS 0.007604f
C1317 B.n442 VSUBS 0.007604f
C1318 B.n443 VSUBS 0.007604f
C1319 B.n444 VSUBS 0.007604f
C1320 B.n445 VSUBS 0.007604f
C1321 B.n446 VSUBS 0.007604f
C1322 B.n447 VSUBS 0.007604f
C1323 B.n448 VSUBS 0.007604f
C1324 B.n449 VSUBS 0.007604f
C1325 B.n450 VSUBS 0.007604f
C1326 B.n451 VSUBS 0.007604f
C1327 B.n452 VSUBS 0.007604f
C1328 B.n453 VSUBS 0.007604f
C1329 B.n454 VSUBS 0.007604f
C1330 B.n455 VSUBS 0.007604f
C1331 B.n456 VSUBS 0.007604f
C1332 B.n457 VSUBS 0.007604f
C1333 B.n458 VSUBS 0.007604f
C1334 B.n459 VSUBS 0.007604f
C1335 B.n460 VSUBS 0.007604f
C1336 B.n461 VSUBS 0.007604f
C1337 B.n462 VSUBS 0.007604f
C1338 B.n463 VSUBS 0.007604f
C1339 B.n464 VSUBS 0.007604f
C1340 B.n465 VSUBS 0.007604f
C1341 B.n466 VSUBS 0.007604f
C1342 B.n467 VSUBS 0.007604f
C1343 B.n468 VSUBS 0.007604f
C1344 B.n469 VSUBS 0.007604f
C1345 B.n470 VSUBS 0.007604f
C1346 B.n471 VSUBS 0.007604f
C1347 B.n472 VSUBS 0.007604f
C1348 B.n473 VSUBS 0.007604f
C1349 B.n474 VSUBS 0.007604f
C1350 B.n475 VSUBS 0.007604f
C1351 B.n476 VSUBS 0.007604f
C1352 B.n477 VSUBS 0.007604f
C1353 B.n478 VSUBS 0.007604f
C1354 B.n479 VSUBS 0.007604f
C1355 B.n480 VSUBS 0.007604f
C1356 B.n481 VSUBS 0.007604f
C1357 B.n482 VSUBS 0.007604f
C1358 B.n483 VSUBS 0.007604f
C1359 B.n484 VSUBS 0.007604f
C1360 B.n485 VSUBS 0.007604f
C1361 B.n486 VSUBS 0.007604f
C1362 B.n487 VSUBS 0.007604f
C1363 B.n488 VSUBS 0.007604f
C1364 B.n489 VSUBS 0.007604f
C1365 B.n490 VSUBS 0.007604f
C1366 B.n491 VSUBS 0.007604f
C1367 B.n492 VSUBS 0.007604f
C1368 B.n493 VSUBS 0.007604f
C1369 B.n494 VSUBS 0.007604f
C1370 B.n495 VSUBS 0.007604f
C1371 B.n496 VSUBS 0.007604f
C1372 B.n497 VSUBS 0.007604f
C1373 B.n498 VSUBS 0.007604f
C1374 B.n499 VSUBS 0.007604f
C1375 B.n500 VSUBS 0.007604f
C1376 B.n501 VSUBS 0.007604f
C1377 B.n502 VSUBS 0.007604f
C1378 B.n503 VSUBS 0.007604f
C1379 B.n504 VSUBS 0.007604f
C1380 B.n505 VSUBS 0.007604f
C1381 B.n506 VSUBS 0.007604f
C1382 B.n507 VSUBS 0.007604f
C1383 B.n508 VSUBS 0.007604f
C1384 B.n509 VSUBS 0.007604f
C1385 B.n510 VSUBS 0.007604f
C1386 B.n511 VSUBS 0.007604f
C1387 B.n512 VSUBS 0.007604f
C1388 B.n513 VSUBS 0.007604f
C1389 B.n514 VSUBS 0.007604f
C1390 B.n515 VSUBS 0.007604f
C1391 B.n516 VSUBS 0.007604f
C1392 B.n517 VSUBS 0.007604f
C1393 B.n518 VSUBS 0.007604f
C1394 B.n519 VSUBS 0.007604f
C1395 B.n520 VSUBS 0.007604f
C1396 B.n521 VSUBS 0.007604f
C1397 B.n522 VSUBS 0.007604f
C1398 B.n523 VSUBS 0.007604f
C1399 B.n524 VSUBS 0.007604f
C1400 B.n525 VSUBS 0.007604f
C1401 B.n526 VSUBS 0.007604f
C1402 B.n527 VSUBS 0.007604f
C1403 B.n528 VSUBS 0.007604f
C1404 B.n529 VSUBS 0.007604f
C1405 B.n530 VSUBS 0.007604f
C1406 B.n531 VSUBS 0.007604f
C1407 B.n532 VSUBS 0.007604f
C1408 B.n533 VSUBS 0.007604f
C1409 B.n534 VSUBS 0.007604f
C1410 B.n535 VSUBS 0.007604f
C1411 B.n536 VSUBS 0.007604f
C1412 B.n537 VSUBS 0.007604f
C1413 B.n538 VSUBS 0.007604f
C1414 B.n539 VSUBS 0.007604f
C1415 B.n540 VSUBS 0.007604f
C1416 B.n541 VSUBS 0.007604f
C1417 B.n542 VSUBS 0.007604f
C1418 B.n543 VSUBS 0.007604f
C1419 B.n544 VSUBS 0.007604f
C1420 B.n545 VSUBS 0.007604f
C1421 B.n546 VSUBS 0.007604f
C1422 B.n547 VSUBS 0.007604f
C1423 B.n548 VSUBS 0.007604f
C1424 B.n549 VSUBS 0.007604f
C1425 B.n550 VSUBS 0.007604f
C1426 B.n551 VSUBS 0.007604f
C1427 B.n552 VSUBS 0.007604f
C1428 B.n553 VSUBS 0.017487f
C1429 B.n554 VSUBS 0.018746f
C1430 B.n555 VSUBS 0.018746f
C1431 B.n556 VSUBS 0.007604f
C1432 B.n557 VSUBS 0.007604f
C1433 B.n558 VSUBS 0.007604f
C1434 B.n559 VSUBS 0.007604f
C1435 B.n560 VSUBS 0.007604f
C1436 B.n561 VSUBS 0.007604f
C1437 B.n562 VSUBS 0.007604f
C1438 B.n563 VSUBS 0.007604f
C1439 B.n564 VSUBS 0.007604f
C1440 B.n565 VSUBS 0.007604f
C1441 B.n566 VSUBS 0.007604f
C1442 B.n567 VSUBS 0.007604f
C1443 B.n568 VSUBS 0.007604f
C1444 B.n569 VSUBS 0.007604f
C1445 B.n570 VSUBS 0.007604f
C1446 B.n571 VSUBS 0.007604f
C1447 B.n572 VSUBS 0.007604f
C1448 B.n573 VSUBS 0.007604f
C1449 B.n574 VSUBS 0.007604f
C1450 B.n575 VSUBS 0.007604f
C1451 B.n576 VSUBS 0.007604f
C1452 B.n577 VSUBS 0.007604f
C1453 B.n578 VSUBS 0.007604f
C1454 B.n579 VSUBS 0.007604f
C1455 B.n580 VSUBS 0.007604f
C1456 B.n581 VSUBS 0.007604f
C1457 B.n582 VSUBS 0.007604f
C1458 B.n583 VSUBS 0.007604f
C1459 B.n584 VSUBS 0.007604f
C1460 B.n585 VSUBS 0.007604f
C1461 B.n586 VSUBS 0.007604f
C1462 B.n587 VSUBS 0.007604f
C1463 B.n588 VSUBS 0.007604f
C1464 B.n589 VSUBS 0.007604f
C1465 B.n590 VSUBS 0.007604f
C1466 B.n591 VSUBS 0.007604f
C1467 B.n592 VSUBS 0.007604f
C1468 B.n593 VSUBS 0.007604f
C1469 B.n594 VSUBS 0.007604f
C1470 B.n595 VSUBS 0.007604f
C1471 B.n596 VSUBS 0.007604f
C1472 B.n597 VSUBS 0.007604f
C1473 B.n598 VSUBS 0.007604f
C1474 B.n599 VSUBS 0.007604f
C1475 B.n600 VSUBS 0.007604f
C1476 B.n601 VSUBS 0.007604f
C1477 B.n602 VSUBS 0.007604f
C1478 B.n603 VSUBS 0.007604f
C1479 B.n604 VSUBS 0.007604f
C1480 B.n605 VSUBS 0.007604f
C1481 B.n606 VSUBS 0.007604f
C1482 B.n607 VSUBS 0.007604f
C1483 B.n608 VSUBS 0.007604f
C1484 B.n609 VSUBS 0.007604f
C1485 B.n610 VSUBS 0.007604f
C1486 B.n611 VSUBS 0.007604f
C1487 B.n612 VSUBS 0.007604f
C1488 B.n613 VSUBS 0.007604f
C1489 B.n614 VSUBS 0.007604f
C1490 B.n615 VSUBS 0.007604f
C1491 B.n616 VSUBS 0.007604f
C1492 B.n617 VSUBS 0.007604f
C1493 B.n618 VSUBS 0.007604f
C1494 B.n619 VSUBS 0.007604f
C1495 B.n620 VSUBS 0.007604f
C1496 B.n621 VSUBS 0.007604f
C1497 B.n622 VSUBS 0.007604f
C1498 B.n623 VSUBS 0.007604f
C1499 B.n624 VSUBS 0.007604f
C1500 B.n625 VSUBS 0.007604f
C1501 B.n626 VSUBS 0.007604f
C1502 B.n627 VSUBS 0.007604f
C1503 B.n628 VSUBS 0.007604f
C1504 B.n629 VSUBS 0.007604f
C1505 B.n630 VSUBS 0.007604f
C1506 B.n631 VSUBS 0.007604f
C1507 B.n632 VSUBS 0.007604f
C1508 B.n633 VSUBS 0.007604f
C1509 B.n634 VSUBS 0.005256f
C1510 B.n635 VSUBS 0.017619f
C1511 B.n636 VSUBS 0.006151f
C1512 B.n637 VSUBS 0.007604f
C1513 B.n638 VSUBS 0.007604f
C1514 B.n639 VSUBS 0.007604f
C1515 B.n640 VSUBS 0.007604f
C1516 B.n641 VSUBS 0.007604f
C1517 B.n642 VSUBS 0.007604f
C1518 B.n643 VSUBS 0.007604f
C1519 B.n644 VSUBS 0.007604f
C1520 B.n645 VSUBS 0.007604f
C1521 B.n646 VSUBS 0.007604f
C1522 B.n647 VSUBS 0.007604f
C1523 B.n648 VSUBS 0.006151f
C1524 B.n649 VSUBS 0.007604f
C1525 B.n650 VSUBS 0.007604f
C1526 B.n651 VSUBS 0.005256f
C1527 B.n652 VSUBS 0.007604f
C1528 B.n653 VSUBS 0.007604f
C1529 B.n654 VSUBS 0.007604f
C1530 B.n655 VSUBS 0.007604f
C1531 B.n656 VSUBS 0.007604f
C1532 B.n657 VSUBS 0.007604f
C1533 B.n658 VSUBS 0.007604f
C1534 B.n659 VSUBS 0.007604f
C1535 B.n660 VSUBS 0.007604f
C1536 B.n661 VSUBS 0.007604f
C1537 B.n662 VSUBS 0.007604f
C1538 B.n663 VSUBS 0.007604f
C1539 B.n664 VSUBS 0.007604f
C1540 B.n665 VSUBS 0.007604f
C1541 B.n666 VSUBS 0.007604f
C1542 B.n667 VSUBS 0.007604f
C1543 B.n668 VSUBS 0.007604f
C1544 B.n669 VSUBS 0.007604f
C1545 B.n670 VSUBS 0.007604f
C1546 B.n671 VSUBS 0.007604f
C1547 B.n672 VSUBS 0.007604f
C1548 B.n673 VSUBS 0.007604f
C1549 B.n674 VSUBS 0.007604f
C1550 B.n675 VSUBS 0.007604f
C1551 B.n676 VSUBS 0.007604f
C1552 B.n677 VSUBS 0.007604f
C1553 B.n678 VSUBS 0.007604f
C1554 B.n679 VSUBS 0.007604f
C1555 B.n680 VSUBS 0.007604f
C1556 B.n681 VSUBS 0.007604f
C1557 B.n682 VSUBS 0.007604f
C1558 B.n683 VSUBS 0.007604f
C1559 B.n684 VSUBS 0.007604f
C1560 B.n685 VSUBS 0.007604f
C1561 B.n686 VSUBS 0.007604f
C1562 B.n687 VSUBS 0.007604f
C1563 B.n688 VSUBS 0.007604f
C1564 B.n689 VSUBS 0.007604f
C1565 B.n690 VSUBS 0.007604f
C1566 B.n691 VSUBS 0.007604f
C1567 B.n692 VSUBS 0.007604f
C1568 B.n693 VSUBS 0.007604f
C1569 B.n694 VSUBS 0.007604f
C1570 B.n695 VSUBS 0.007604f
C1571 B.n696 VSUBS 0.007604f
C1572 B.n697 VSUBS 0.007604f
C1573 B.n698 VSUBS 0.007604f
C1574 B.n699 VSUBS 0.007604f
C1575 B.n700 VSUBS 0.007604f
C1576 B.n701 VSUBS 0.007604f
C1577 B.n702 VSUBS 0.007604f
C1578 B.n703 VSUBS 0.007604f
C1579 B.n704 VSUBS 0.007604f
C1580 B.n705 VSUBS 0.007604f
C1581 B.n706 VSUBS 0.007604f
C1582 B.n707 VSUBS 0.007604f
C1583 B.n708 VSUBS 0.007604f
C1584 B.n709 VSUBS 0.007604f
C1585 B.n710 VSUBS 0.007604f
C1586 B.n711 VSUBS 0.007604f
C1587 B.n712 VSUBS 0.007604f
C1588 B.n713 VSUBS 0.007604f
C1589 B.n714 VSUBS 0.007604f
C1590 B.n715 VSUBS 0.007604f
C1591 B.n716 VSUBS 0.007604f
C1592 B.n717 VSUBS 0.007604f
C1593 B.n718 VSUBS 0.007604f
C1594 B.n719 VSUBS 0.007604f
C1595 B.n720 VSUBS 0.007604f
C1596 B.n721 VSUBS 0.007604f
C1597 B.n722 VSUBS 0.007604f
C1598 B.n723 VSUBS 0.007604f
C1599 B.n724 VSUBS 0.007604f
C1600 B.n725 VSUBS 0.007604f
C1601 B.n726 VSUBS 0.007604f
C1602 B.n727 VSUBS 0.007604f
C1603 B.n728 VSUBS 0.007604f
C1604 B.n729 VSUBS 0.007604f
C1605 B.n730 VSUBS 0.018746f
C1606 B.n731 VSUBS 0.017487f
C1607 B.n732 VSUBS 0.017487f
C1608 B.n733 VSUBS 0.007604f
C1609 B.n734 VSUBS 0.007604f
C1610 B.n735 VSUBS 0.007604f
C1611 B.n736 VSUBS 0.007604f
C1612 B.n737 VSUBS 0.007604f
C1613 B.n738 VSUBS 0.007604f
C1614 B.n739 VSUBS 0.007604f
C1615 B.n740 VSUBS 0.007604f
C1616 B.n741 VSUBS 0.007604f
C1617 B.n742 VSUBS 0.007604f
C1618 B.n743 VSUBS 0.007604f
C1619 B.n744 VSUBS 0.007604f
C1620 B.n745 VSUBS 0.007604f
C1621 B.n746 VSUBS 0.007604f
C1622 B.n747 VSUBS 0.007604f
C1623 B.n748 VSUBS 0.007604f
C1624 B.n749 VSUBS 0.007604f
C1625 B.n750 VSUBS 0.007604f
C1626 B.n751 VSUBS 0.007604f
C1627 B.n752 VSUBS 0.007604f
C1628 B.n753 VSUBS 0.007604f
C1629 B.n754 VSUBS 0.007604f
C1630 B.n755 VSUBS 0.007604f
C1631 B.n756 VSUBS 0.007604f
C1632 B.n757 VSUBS 0.007604f
C1633 B.n758 VSUBS 0.007604f
C1634 B.n759 VSUBS 0.007604f
C1635 B.n760 VSUBS 0.007604f
C1636 B.n761 VSUBS 0.007604f
C1637 B.n762 VSUBS 0.007604f
C1638 B.n763 VSUBS 0.007604f
C1639 B.n764 VSUBS 0.007604f
C1640 B.n765 VSUBS 0.007604f
C1641 B.n766 VSUBS 0.007604f
C1642 B.n767 VSUBS 0.007604f
C1643 B.n768 VSUBS 0.007604f
C1644 B.n769 VSUBS 0.007604f
C1645 B.n770 VSUBS 0.007604f
C1646 B.n771 VSUBS 0.007604f
C1647 B.n772 VSUBS 0.007604f
C1648 B.n773 VSUBS 0.007604f
C1649 B.n774 VSUBS 0.007604f
C1650 B.n775 VSUBS 0.007604f
C1651 B.n776 VSUBS 0.007604f
C1652 B.n777 VSUBS 0.007604f
C1653 B.n778 VSUBS 0.007604f
C1654 B.n779 VSUBS 0.007604f
C1655 B.n780 VSUBS 0.007604f
C1656 B.n781 VSUBS 0.007604f
C1657 B.n782 VSUBS 0.007604f
C1658 B.n783 VSUBS 0.007604f
C1659 B.n784 VSUBS 0.007604f
C1660 B.n785 VSUBS 0.007604f
C1661 B.n786 VSUBS 0.007604f
C1662 B.n787 VSUBS 0.009923f
C1663 B.n788 VSUBS 0.010571f
C1664 B.n789 VSUBS 0.021021f
.ends

