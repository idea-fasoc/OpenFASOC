* NGSPICE file created from opamp_sample_0014.ext - technology: sky130A

.subckt opamp_sample_0014 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t135 GND.t133 GND.t134 GND.t81 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X1 a_n2675_n4106.t8 DIFFPAIR_BIAS.t10 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X2 GND.t132 GND.t130 GND.t131 GND.t77 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X3 VDD.t49 a_n6918_10482.t6 a_n2500_9133.t5 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=1.5768 ps=5.82 w=2.19 l=3.2
X4 VOUT.t48 a_n2500_9133.t0 sky130_fd_pr__cap_mim_m3_1 l=12.27 w=19.55
X5 VOUT.t45 CS_BIAS.t24 GND.t138 GND.t26 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X6 VDD.t131 VDD.t129 VDD.t130 VDD.t57 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X7 CS_BIAS.t23 CS_BIAS.t22 GND.t143 GND.t23 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X8 VDD.t128 VDD.t126 VDD.t127 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X9 VDD.t125 VDD.t122 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X10 VDD.t13 a_n12950_8244.t4 VOUT.t12 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X11 GND.t129 GND.t127 GND.t128 GND.t102 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X12 VDD.t50 a_n12950_8244.t5 VOUT.t20 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X13 VDD.t121 VDD.t119 VDD.t120 VDD.t53 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X14 VDD.t118 VDD.t116 VDD.t117 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X15 VOUT.t49 a_n2500_9133.t0 sky130_fd_pr__cap_mim_m3_1 l=12.27 w=19.55
X16 GND.t126 GND.t123 GND.t125 GND.t124 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=0 ps=0 w=5.71 l=2.16
X17 GND.t122 GND.t120 GND.t121 GND.t95 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=0 ps=0 w=6.8 l=4.8
X18 VOUT.t41 a_n12950_8244.t6 VDD.t142 VDD.t137 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X19 VOUT.t46 CS_BIAS.t25 GND.t141 GND.t23 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X20 VDD.t47 a_n6918_10482.t7 a_n7062_10679.t9 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X21 VDD.t45 a_n6918_10482.t8 a_n7062_10679.t8 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=1.5768 ps=5.82 w=2.19 l=3.2
X22 VDD.t144 a_n12950_8244.t7 VOUT.t43 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X23 GND.t50 CS_BIAS.t20 CS_BIAS.t21 GND.t44 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X24 VOUT.t47 CS_BIAS.t26 GND.t142 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X25 VOUT.t14 a_n12950_8244.t8 VDD.t14 VDD.t4 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X26 CS_BIAS.t19 CS_BIAS.t18 GND.t39 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X27 a_n7062_10679.t1 a_n6918_10482.t2 a_n6918_10482.t3 VDD.t23 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=1.5768 ps=5.82 w=2.19 l=3.2
X28 GND.t119 GND.t117 GND.t118 GND.t70 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=0 ps=0 w=6.8 l=4.8
X29 a_n7062_10679.t7 a_n6918_10482.t9 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0.7227 ps=2.85 w=2.19 l=3.2
X30 VOUT.t39 a_n12950_8244.t9 VDD.t139 VDD.t137 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X31 VOUT.t38 a_n12950_8244.t10 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X32 VDD.t115 VDD.t113 VDD.t114 VDD.t57 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X33 VDD.t112 VDD.t110 VDD.t111 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X34 a_n2675_n4106.t7 DIFFPAIR_BIAS.t11 GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X35 VDD.t109 VDD.t107 VDD.t108 VDD.t75 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X36 DIFFPAIR_BIAS.t9 DIFFPAIR_BIAS.t8 GND.t56 GND.t55 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X37 VDD.t106 VDD.t104 VDD.t105 VDD.t68 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X38 GND.t38 CS_BIAS.t27 VOUT.t25 GND.t28 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X39 VDD.t10 a_n12950_8244.t11 VOUT.t10 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X40 VOUT.t2 CS_BIAS.t28 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X41 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t137 GND.t136 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X42 VOUT.t28 a_n12950_8244.t12 VDD.t133 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X43 VOUT.t4 CS_BIAS.t29 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X44 GND.t18 CS_BIAS.t30 VOUT.t17 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X45 VDD.t103 VDD.t101 VDD.t102 VDD.t61 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X46 GND.t116 GND.t114 VN.t1 GND.t115 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X47 VDD.t100 VDD.t98 VDD.t99 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X48 a_n2500_9133.t1 a_n6918_10482.t10 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0.7227 ps=2.85 w=2.19 l=3.2
X49 a_n2500_9133.t9 a_n6918_10482.t11 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X50 CS_BIAS.t17 CS_BIAS.t16 GND.t30 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X51 GND.t40 CS_BIAS.t14 CS_BIAS.t15 GND.t33 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X52 VDD.t97 VDD.t95 VDD.t96 VDD.t68 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X53 a_n12950_8244.t2 VN.t2 a_n2675_n4106.t0 GND.t25 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=4.896 ps=15.04 w=6.8 l=4.8
X54 a_n2675_n4106.t6 DIFFPAIR_BIAS.t12 GND.t43 GND.t42 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X55 GND.t29 CS_BIAS.t12 CS_BIAS.t13 GND.t28 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X56 GND.t113 GND.t111 GND.t112 GND.t81 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X57 a_n12950_8244.t1 a_n6918_10482.t12 a_n2500_9133.t10 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=1.5768 ps=5.82 w=2.19 l=3.2
X58 VDD.t94 VDD.t92 VDD.t93 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X59 GND.t110 GND.t108 GND.t109 GND.t77 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X60 GND.t45 CS_BIAS.t31 VOUT.t26 GND.t44 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X61 VOUT.t9 a_n12950_8244.t13 VDD.t9 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X62 GND.t49 CS_BIAS.t32 VOUT.t30 GND.t2 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X63 GND.t107 GND.t105 GND.t106 GND.t102 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X64 a_n7062_10679.t6 a_n6918_10482.t13 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X65 GND.t104 GND.t101 GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X66 VOUT.t37 a_n12950_8244.t14 VDD.t136 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X67 GND.t54 CS_BIAS.t33 VOUT.t35 GND.t33 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X68 VDD.t91 VDD.t89 VDD.t90 VDD.t68 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X69 VOUT.t8 a_n12950_8244.t15 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X70 a_n7062_10679.t5 a_n6918_10482.t14 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0.7227 ps=2.85 w=2.19 l=3.2
X71 VDD.t134 a_n12950_8244.t16 VOUT.t32 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X72 GND.t100 GND.t98 VP.t1 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X73 GND.t10 CS_BIAS.t34 VOUT.t3 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X74 GND.t97 GND.t94 GND.t96 GND.t95 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=0 ps=0 w=6.8 l=4.8
X75 GND.t93 GND.t91 GND.t92 GND.t63 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X76 a_n8118_10679# a_n8118_10679# a_n8118_10679# VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=3.1536 ps=11.64 w=2.19 l=3.2
X77 a_n2500_9133.t8 a_n6918_10482.t15 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0.7227 ps=2.85 w=2.19 l=3.2
X78 VOUT.t0 CS_BIAS.t35 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X79 GND.t90 GND.t88 GND.t89 GND.t63 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X80 a_n6918_10482.t5 VP.t2 a_n2675_n4106.t2 GND.t35 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=4.896 ps=15.04 w=6.8 l=4.8
X81 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t37 GND.t36 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X82 VOUT.t40 a_n12950_8244.t17 VDD.t141 VDD.t137 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X83 VDD.t88 VDD.t86 VDD.t87 VDD.t57 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X84 VDD.t31 a_n6918_10482.t16 a_n2500_9133.t3 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X85 VDD.t85 VDD.t82 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X86 a_7190_10679# a_7190_10679# a_7190_10679# VDD.t15 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=3.1536 ps=11.64 w=2.19 l=3.2
X87 GND.t87 GND.t84 GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=0 ps=0 w=5.71 l=2.16
X88 a_n2500_9133.t4 a_n6918_10482.t17 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X89 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t140 GND.t139 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X90 GND.t83 GND.t80 GND.t82 GND.t81 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X91 VOUT.t34 CS_BIAS.t36 GND.t53 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X92 GND.t22 CS_BIAS.t37 VOUT.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X93 GND.t79 GND.t76 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X94 VDD.t81 VDD.t78 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X95 CS_BIAS.t11 CS_BIAS.t10 GND.t19 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X96 VOUT.t21 CS_BIAS.t38 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X97 GND.t3 CS_BIAS.t8 CS_BIAS.t9 GND.t2 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X98 a_n6918_10482.t4 VP.t3 a_n2675_n4106.t1 GND.t25 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=4.896 ps=15.04 w=6.8 l=4.8
X99 VOUT.t27 a_n12950_8244.t18 VDD.t132 VDD.t4 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X100 VN.t0 GND.t66 GND.t68 GND.t67 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X101 VP.t0 GND.t73 GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X102 VDD.t77 VDD.t74 VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X103 VDD.t27 a_n6918_10482.t18 a_n2500_9133.t6 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=1.5768 ps=5.82 w=2.19 l=3.2
X104 GND.t51 CS_BIAS.t39 VOUT.t31 GND.t44 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X105 VOUT.t50 a_n2500_9133.t0 sky130_fd_pr__cap_mim_m3_1 l=12.27 w=19.55
X106 GND.t13 CS_BIAS.t40 VOUT.t13 GND.t2 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X107 GND.t72 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=0 ps=0 w=6.8 l=4.8
X108 VOUT.t36 a_n12950_8244.t19 VDD.t135 VDD.t4 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X109 VOUT.t19 CS_BIAS.t41 GND.t24 GND.t23 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X110 VDD.t6 a_n12950_8244.t20 VOUT.t7 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X111 GND.t34 CS_BIAS.t42 VOUT.t23 GND.t33 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=1.7556 ps=5.98 w=5.32 l=2.11
X112 VOUT.t16 CS_BIAS.t43 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X113 CS_BIAS.t7 CS_BIAS.t6 GND.t59 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X114 a_n2675_n4106.t5 DIFFPAIR_BIAS.t13 GND.t58 GND.t57 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X115 VOUT.t6 a_n12950_8244.t21 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=1.1847 ps=4.25 w=3.59 l=3.83
X116 VDD.t73 VDD.t71 VDD.t72 VDD.t61 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X117 VOUT.t42 a_n12950_8244.t22 VDD.t143 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X118 VDD.t25 a_n6918_10482.t19 a_n7062_10679.t4 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=1.5768 ps=5.82 w=2.19 l=3.2
X119 a_n2675_n4106.t4 DIFFPAIR_BIAS.t14 GND.t61 GND.t60 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X120 VDD.t70 VDD.t67 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X121 a_n7062_10679.t3 a_n6918_10482.t20 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X122 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=4.1112 pd=12.86 as=4.1112 ps=12.86 w=5.71 l=2.16
X123 a_n12950_8244.t0 a_n6918_10482.t21 a_n2500_9133.t2 VDD.t23 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=1.5768 ps=5.82 w=2.19 l=3.2
X124 VOUT.t44 a_n12950_8244.t23 VDD.t145 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X125 VDD.t11 a_n12950_8244.t24 VOUT.t11 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X126 GND.t48 CS_BIAS.t44 VOUT.t29 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X127 VDD.t3 a_n12950_8244.t25 VOUT.t5 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=1.1847 ps=4.25 w=3.59 l=3.83
X128 GND.t52 CS_BIAS.t45 VOUT.t33 GND.t28 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X129 VOUT.t24 a_n12950_8244.t26 VDD.t51 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X130 VDD.t22 a_n6918_10482.t22 a_n7062_10679.t2 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X131 VOUT.t22 CS_BIAS.t46 GND.t32 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X132 VDD.t66 VDD.t64 VDD.t65 VDD.t61 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X133 VDD.t18 a_n6918_10482.t23 a_n2500_9133.t7 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.7227 pd=2.85 as=0.7227 ps=2.85 w=2.19 l=3.2
X134 VOUT.t15 CS_BIAS.t47 GND.t14 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=3.8304 ps=12.08 w=5.32 l=2.11
X135 GND.t7 CS_BIAS.t4 CS_BIAS.t5 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X136 VDD.t63 VDD.t60 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X137 a_n7062_10679.t0 a_n6918_10482.t0 a_n6918_10482.t1 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=1.5768 ps=5.82 w=2.19 l=3.2
X138 CS_BIAS.t3 CS_BIAS.t2 GND.t31 GND.t26 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X139 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=3.8304 pd=12.08 as=0 ps=0 w=5.32 l=2.11
X140 VOUT.t51 a_n2500_9133.t0 sky130_fd_pr__cap_mim_m3_1 l=12.27 w=19.55
X141 VOUT.t1 a_n12950_8244.t27 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.1847 pd=4.25 as=2.5848 ps=8.62 w=3.59 l=3.83
X142 GND.t41 CS_BIAS.t0 CS_BIAS.t1 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.7556 pd=5.98 as=1.7556 ps=5.98 w=5.32 l=2.11
X143 VDD.t59 VDD.t56 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8 ad=2.5848 pd=8.62 as=0 ps=0 w=3.59 l=3.83
X144 VDD.t55 VDD.t52 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8 ad=1.5768 pd=5.82 as=0 ps=0 w=2.19 l=3.2
X145 a_n12950_8244.t3 VN.t3 a_n2675_n4106.t3 GND.t35 sky130_fd_pr__nfet_01v8 ad=4.896 pd=15.04 as=4.896 ps=15.04 w=6.8 l=4.8
R0 GND.n6188 GND.n307 2194.01
R1 GND.n5338 GND.n5337 1749.94
R2 GND.n4656 GND.n1857 860.073
R3 GND.n4190 GND.n1859 860.073
R4 GND.n3515 GND.n1301 860.073
R5 GND.n5031 GND.n1231 860.073
R6 GND.n1221 GND.n1169 821.635
R7 GND.n5006 GND.n1167 821.635
R8 GND.n1017 GND.n966 821.635
R9 GND.n5190 GND.n5189 821.635
R10 GND.n2537 GND.n1884 821.635
R11 GND.n2498 GND.n1882 821.635
R12 GND.n1999 GND.n82 821.635
R13 GND.n6503 GND.n78 821.635
R14 GND.n6501 GND.n84 778.39
R15 GND.n6446 GND.n80 778.39
R16 GND.n2543 GND.n1881 778.39
R17 GND.n4638 GND.n1885 778.39
R18 GND.n5099 GND.n1171 778.39
R19 GND.n5101 GND.n1165 778.39
R20 GND.n1016 GND.n1015 778.39
R21 GND.n5262 GND.n970 778.39
R22 GND.n5459 GND.n746 699.111
R23 GND.n6189 GND.n308 699.111
R24 GND.n6346 GND.n218 699.111
R25 GND.n5339 GND.n868 699.111
R26 GND.n5460 GND.n5459 585
R27 GND.n5459 GND.n5458 585
R28 GND.n750 GND.n749 585
R29 GND.n5457 GND.n750 585
R30 GND.n5455 GND.n5454 585
R31 GND.n5456 GND.n5455 585
R32 GND.n5453 GND.n752 585
R33 GND.n752 GND.n751 585
R34 GND.n5452 GND.n5451 585
R35 GND.n5451 GND.n5450 585
R36 GND.n757 GND.n756 585
R37 GND.n5449 GND.n757 585
R38 GND.n5447 GND.n5446 585
R39 GND.n5448 GND.n5447 585
R40 GND.n5445 GND.n759 585
R41 GND.n759 GND.n758 585
R42 GND.n5444 GND.n5443 585
R43 GND.n5443 GND.n5442 585
R44 GND.n765 GND.n764 585
R45 GND.n5441 GND.n765 585
R46 GND.n5439 GND.n5438 585
R47 GND.n5440 GND.n5439 585
R48 GND.n5437 GND.n767 585
R49 GND.n767 GND.n766 585
R50 GND.n5436 GND.n5435 585
R51 GND.n5435 GND.n5434 585
R52 GND.n773 GND.n772 585
R53 GND.n5433 GND.n773 585
R54 GND.n5431 GND.n5430 585
R55 GND.n5432 GND.n5431 585
R56 GND.n5429 GND.n775 585
R57 GND.n775 GND.n774 585
R58 GND.n5428 GND.n5427 585
R59 GND.n5427 GND.n5426 585
R60 GND.n781 GND.n780 585
R61 GND.n5425 GND.n781 585
R62 GND.n5423 GND.n5422 585
R63 GND.n5424 GND.n5423 585
R64 GND.n5421 GND.n783 585
R65 GND.n783 GND.n782 585
R66 GND.n5420 GND.n5419 585
R67 GND.n5419 GND.n5418 585
R68 GND.n789 GND.n788 585
R69 GND.n5417 GND.n789 585
R70 GND.n5415 GND.n5414 585
R71 GND.n5416 GND.n5415 585
R72 GND.n5413 GND.n791 585
R73 GND.n791 GND.n790 585
R74 GND.n5412 GND.n5411 585
R75 GND.n5411 GND.n5410 585
R76 GND.n797 GND.n796 585
R77 GND.n5409 GND.n797 585
R78 GND.n5407 GND.n5406 585
R79 GND.n5408 GND.n5407 585
R80 GND.n5405 GND.n799 585
R81 GND.n799 GND.n798 585
R82 GND.n5404 GND.n5403 585
R83 GND.n5403 GND.n5402 585
R84 GND.n805 GND.n804 585
R85 GND.n5401 GND.n805 585
R86 GND.n5399 GND.n5398 585
R87 GND.n5400 GND.n5399 585
R88 GND.n5397 GND.n807 585
R89 GND.n807 GND.n806 585
R90 GND.n5396 GND.n5395 585
R91 GND.n5395 GND.n5394 585
R92 GND.n813 GND.n812 585
R93 GND.n5393 GND.n813 585
R94 GND.n5391 GND.n5390 585
R95 GND.n5392 GND.n5391 585
R96 GND.n5389 GND.n815 585
R97 GND.n815 GND.n814 585
R98 GND.n5388 GND.n5387 585
R99 GND.n5387 GND.n5386 585
R100 GND.n821 GND.n820 585
R101 GND.n5385 GND.n821 585
R102 GND.n5383 GND.n5382 585
R103 GND.n5384 GND.n5383 585
R104 GND.n5381 GND.n823 585
R105 GND.n823 GND.n822 585
R106 GND.n5380 GND.n5379 585
R107 GND.n5379 GND.n5378 585
R108 GND.n829 GND.n828 585
R109 GND.n5377 GND.n829 585
R110 GND.n5375 GND.n5374 585
R111 GND.n5376 GND.n5375 585
R112 GND.n5373 GND.n831 585
R113 GND.n831 GND.n830 585
R114 GND.n5372 GND.n5371 585
R115 GND.n5371 GND.n5370 585
R116 GND.n837 GND.n836 585
R117 GND.n5369 GND.n837 585
R118 GND.n5367 GND.n5366 585
R119 GND.n5368 GND.n5367 585
R120 GND.n5365 GND.n839 585
R121 GND.n839 GND.n838 585
R122 GND.n5364 GND.n5363 585
R123 GND.n5363 GND.n5362 585
R124 GND.n845 GND.n844 585
R125 GND.n5361 GND.n845 585
R126 GND.n5359 GND.n5358 585
R127 GND.n5360 GND.n5359 585
R128 GND.n5357 GND.n847 585
R129 GND.n847 GND.n846 585
R130 GND.n5356 GND.n5355 585
R131 GND.n5355 GND.n5354 585
R132 GND.n853 GND.n852 585
R133 GND.n5353 GND.n853 585
R134 GND.n5351 GND.n5350 585
R135 GND.n5352 GND.n5351 585
R136 GND.n5349 GND.n855 585
R137 GND.n855 GND.n854 585
R138 GND.n5348 GND.n5347 585
R139 GND.n5347 GND.n5346 585
R140 GND.n861 GND.n860 585
R141 GND.n5345 GND.n861 585
R142 GND.n5343 GND.n5342 585
R143 GND.n5344 GND.n5343 585
R144 GND.n5341 GND.n863 585
R145 GND.n863 GND.n862 585
R146 GND.n5340 GND.n5339 585
R147 GND.n5339 GND.n5338 585
R148 GND.n747 GND.n746 585
R149 GND.n746 GND.n745 585
R150 GND.n5465 GND.n5464 585
R151 GND.n5466 GND.n5465 585
R152 GND.n744 GND.n743 585
R153 GND.n5467 GND.n744 585
R154 GND.n5470 GND.n5469 585
R155 GND.n5469 GND.n5468 585
R156 GND.n741 GND.n740 585
R157 GND.n740 GND.n739 585
R158 GND.n5475 GND.n5474 585
R159 GND.n5476 GND.n5475 585
R160 GND.n738 GND.n737 585
R161 GND.n5477 GND.n738 585
R162 GND.n5480 GND.n5479 585
R163 GND.n5479 GND.n5478 585
R164 GND.n735 GND.n734 585
R165 GND.n734 GND.n733 585
R166 GND.n5485 GND.n5484 585
R167 GND.n5486 GND.n5485 585
R168 GND.n732 GND.n731 585
R169 GND.n5487 GND.n732 585
R170 GND.n5490 GND.n5489 585
R171 GND.n5489 GND.n5488 585
R172 GND.n729 GND.n728 585
R173 GND.n728 GND.n727 585
R174 GND.n5495 GND.n5494 585
R175 GND.n5496 GND.n5495 585
R176 GND.n726 GND.n725 585
R177 GND.n5497 GND.n726 585
R178 GND.n5500 GND.n5499 585
R179 GND.n5499 GND.n5498 585
R180 GND.n723 GND.n722 585
R181 GND.n722 GND.n721 585
R182 GND.n5505 GND.n5504 585
R183 GND.n5506 GND.n5505 585
R184 GND.n720 GND.n719 585
R185 GND.n5507 GND.n720 585
R186 GND.n5510 GND.n5509 585
R187 GND.n5509 GND.n5508 585
R188 GND.n717 GND.n716 585
R189 GND.n716 GND.n715 585
R190 GND.n5515 GND.n5514 585
R191 GND.n5516 GND.n5515 585
R192 GND.n714 GND.n713 585
R193 GND.n5517 GND.n714 585
R194 GND.n5520 GND.n5519 585
R195 GND.n5519 GND.n5518 585
R196 GND.n711 GND.n710 585
R197 GND.n710 GND.n709 585
R198 GND.n5525 GND.n5524 585
R199 GND.n5526 GND.n5525 585
R200 GND.n708 GND.n707 585
R201 GND.n5527 GND.n708 585
R202 GND.n5530 GND.n5529 585
R203 GND.n5529 GND.n5528 585
R204 GND.n705 GND.n704 585
R205 GND.n704 GND.n703 585
R206 GND.n5535 GND.n5534 585
R207 GND.n5536 GND.n5535 585
R208 GND.n702 GND.n701 585
R209 GND.n5537 GND.n702 585
R210 GND.n5540 GND.n5539 585
R211 GND.n5539 GND.n5538 585
R212 GND.n699 GND.n698 585
R213 GND.n698 GND.n697 585
R214 GND.n5545 GND.n5544 585
R215 GND.n5546 GND.n5545 585
R216 GND.n696 GND.n695 585
R217 GND.n5547 GND.n696 585
R218 GND.n5550 GND.n5549 585
R219 GND.n5549 GND.n5548 585
R220 GND.n693 GND.n692 585
R221 GND.n692 GND.n691 585
R222 GND.n5555 GND.n5554 585
R223 GND.n5556 GND.n5555 585
R224 GND.n690 GND.n689 585
R225 GND.n5557 GND.n690 585
R226 GND.n5560 GND.n5559 585
R227 GND.n5559 GND.n5558 585
R228 GND.n687 GND.n686 585
R229 GND.n686 GND.n685 585
R230 GND.n5565 GND.n5564 585
R231 GND.n5566 GND.n5565 585
R232 GND.n684 GND.n683 585
R233 GND.n5567 GND.n684 585
R234 GND.n5570 GND.n5569 585
R235 GND.n5569 GND.n5568 585
R236 GND.n681 GND.n680 585
R237 GND.n680 GND.n679 585
R238 GND.n5575 GND.n5574 585
R239 GND.n5576 GND.n5575 585
R240 GND.n678 GND.n677 585
R241 GND.n5577 GND.n678 585
R242 GND.n5580 GND.n5579 585
R243 GND.n5579 GND.n5578 585
R244 GND.n675 GND.n674 585
R245 GND.n674 GND.n673 585
R246 GND.n5585 GND.n5584 585
R247 GND.n5586 GND.n5585 585
R248 GND.n672 GND.n671 585
R249 GND.n5587 GND.n672 585
R250 GND.n5590 GND.n5589 585
R251 GND.n5589 GND.n5588 585
R252 GND.n669 GND.n668 585
R253 GND.n668 GND.n667 585
R254 GND.n5595 GND.n5594 585
R255 GND.n5596 GND.n5595 585
R256 GND.n666 GND.n665 585
R257 GND.n5597 GND.n666 585
R258 GND.n5600 GND.n5599 585
R259 GND.n5599 GND.n5598 585
R260 GND.n663 GND.n662 585
R261 GND.n662 GND.n661 585
R262 GND.n5605 GND.n5604 585
R263 GND.n5606 GND.n5605 585
R264 GND.n660 GND.n659 585
R265 GND.n5607 GND.n660 585
R266 GND.n5610 GND.n5609 585
R267 GND.n5609 GND.n5608 585
R268 GND.n657 GND.n656 585
R269 GND.n656 GND.n655 585
R270 GND.n5615 GND.n5614 585
R271 GND.n5616 GND.n5615 585
R272 GND.n654 GND.n653 585
R273 GND.n5617 GND.n654 585
R274 GND.n5620 GND.n5619 585
R275 GND.n5619 GND.n5618 585
R276 GND.n651 GND.n650 585
R277 GND.n650 GND.n649 585
R278 GND.n5625 GND.n5624 585
R279 GND.n5626 GND.n5625 585
R280 GND.n648 GND.n647 585
R281 GND.n5627 GND.n648 585
R282 GND.n5630 GND.n5629 585
R283 GND.n5629 GND.n5628 585
R284 GND.n645 GND.n644 585
R285 GND.n644 GND.n643 585
R286 GND.n5635 GND.n5634 585
R287 GND.n5636 GND.n5635 585
R288 GND.n642 GND.n641 585
R289 GND.n5637 GND.n642 585
R290 GND.n5640 GND.n5639 585
R291 GND.n5639 GND.n5638 585
R292 GND.n639 GND.n638 585
R293 GND.n638 GND.n637 585
R294 GND.n5645 GND.n5644 585
R295 GND.n5646 GND.n5645 585
R296 GND.n636 GND.n635 585
R297 GND.n5647 GND.n636 585
R298 GND.n5650 GND.n5649 585
R299 GND.n5649 GND.n5648 585
R300 GND.n633 GND.n632 585
R301 GND.n632 GND.n631 585
R302 GND.n5655 GND.n5654 585
R303 GND.n5656 GND.n5655 585
R304 GND.n630 GND.n629 585
R305 GND.n5657 GND.n630 585
R306 GND.n5660 GND.n5659 585
R307 GND.n5659 GND.n5658 585
R308 GND.n627 GND.n626 585
R309 GND.n626 GND.n625 585
R310 GND.n5665 GND.n5664 585
R311 GND.n5666 GND.n5665 585
R312 GND.n624 GND.n623 585
R313 GND.n5667 GND.n624 585
R314 GND.n5670 GND.n5669 585
R315 GND.n5669 GND.n5668 585
R316 GND.n621 GND.n620 585
R317 GND.n620 GND.n619 585
R318 GND.n5675 GND.n5674 585
R319 GND.n5676 GND.n5675 585
R320 GND.n618 GND.n617 585
R321 GND.n5677 GND.n618 585
R322 GND.n5680 GND.n5679 585
R323 GND.n5679 GND.n5678 585
R324 GND.n615 GND.n614 585
R325 GND.n614 GND.n613 585
R326 GND.n5685 GND.n5684 585
R327 GND.n5686 GND.n5685 585
R328 GND.n612 GND.n611 585
R329 GND.n5687 GND.n612 585
R330 GND.n5690 GND.n5689 585
R331 GND.n5689 GND.n5688 585
R332 GND.n609 GND.n608 585
R333 GND.n608 GND.n607 585
R334 GND.n5695 GND.n5694 585
R335 GND.n5696 GND.n5695 585
R336 GND.n606 GND.n605 585
R337 GND.n5697 GND.n606 585
R338 GND.n5700 GND.n5699 585
R339 GND.n5699 GND.n5698 585
R340 GND.n603 GND.n602 585
R341 GND.n602 GND.n601 585
R342 GND.n5705 GND.n5704 585
R343 GND.n5706 GND.n5705 585
R344 GND.n600 GND.n599 585
R345 GND.n5707 GND.n600 585
R346 GND.n5710 GND.n5709 585
R347 GND.n5709 GND.n5708 585
R348 GND.n597 GND.n596 585
R349 GND.n596 GND.n595 585
R350 GND.n5715 GND.n5714 585
R351 GND.n5716 GND.n5715 585
R352 GND.n594 GND.n593 585
R353 GND.n5717 GND.n594 585
R354 GND.n5720 GND.n5719 585
R355 GND.n5719 GND.n5718 585
R356 GND.n591 GND.n590 585
R357 GND.n590 GND.n589 585
R358 GND.n5725 GND.n5724 585
R359 GND.n5726 GND.n5725 585
R360 GND.n588 GND.n587 585
R361 GND.n5727 GND.n588 585
R362 GND.n5730 GND.n5729 585
R363 GND.n5729 GND.n5728 585
R364 GND.n585 GND.n584 585
R365 GND.n584 GND.n583 585
R366 GND.n5735 GND.n5734 585
R367 GND.n5736 GND.n5735 585
R368 GND.n582 GND.n581 585
R369 GND.n5737 GND.n582 585
R370 GND.n5740 GND.n5739 585
R371 GND.n5739 GND.n5738 585
R372 GND.n579 GND.n578 585
R373 GND.n578 GND.n577 585
R374 GND.n5745 GND.n5744 585
R375 GND.n5746 GND.n5745 585
R376 GND.n576 GND.n575 585
R377 GND.n5747 GND.n576 585
R378 GND.n5750 GND.n5749 585
R379 GND.n5749 GND.n5748 585
R380 GND.n573 GND.n572 585
R381 GND.n572 GND.n571 585
R382 GND.n5755 GND.n5754 585
R383 GND.n5756 GND.n5755 585
R384 GND.n570 GND.n569 585
R385 GND.n5757 GND.n570 585
R386 GND.n5760 GND.n5759 585
R387 GND.n5759 GND.n5758 585
R388 GND.n567 GND.n566 585
R389 GND.n566 GND.n565 585
R390 GND.n5765 GND.n5764 585
R391 GND.n5766 GND.n5765 585
R392 GND.n564 GND.n563 585
R393 GND.n5767 GND.n564 585
R394 GND.n5770 GND.n5769 585
R395 GND.n5769 GND.n5768 585
R396 GND.n561 GND.n560 585
R397 GND.n560 GND.n559 585
R398 GND.n5775 GND.n5774 585
R399 GND.n5776 GND.n5775 585
R400 GND.n558 GND.n557 585
R401 GND.n5777 GND.n558 585
R402 GND.n5780 GND.n5779 585
R403 GND.n5779 GND.n5778 585
R404 GND.n555 GND.n554 585
R405 GND.n554 GND.n553 585
R406 GND.n5785 GND.n5784 585
R407 GND.n5786 GND.n5785 585
R408 GND.n552 GND.n551 585
R409 GND.n5787 GND.n552 585
R410 GND.n5790 GND.n5789 585
R411 GND.n5789 GND.n5788 585
R412 GND.n549 GND.n548 585
R413 GND.n548 GND.n547 585
R414 GND.n5795 GND.n5794 585
R415 GND.n5796 GND.n5795 585
R416 GND.n546 GND.n545 585
R417 GND.n5797 GND.n546 585
R418 GND.n5800 GND.n5799 585
R419 GND.n5799 GND.n5798 585
R420 GND.n543 GND.n542 585
R421 GND.n542 GND.n541 585
R422 GND.n5805 GND.n5804 585
R423 GND.n5806 GND.n5805 585
R424 GND.n540 GND.n539 585
R425 GND.n5807 GND.n540 585
R426 GND.n5810 GND.n5809 585
R427 GND.n5809 GND.n5808 585
R428 GND.n537 GND.n536 585
R429 GND.n536 GND.n535 585
R430 GND.n5815 GND.n5814 585
R431 GND.n5816 GND.n5815 585
R432 GND.n534 GND.n533 585
R433 GND.n5817 GND.n534 585
R434 GND.n5820 GND.n5819 585
R435 GND.n5819 GND.n5818 585
R436 GND.n531 GND.n530 585
R437 GND.n530 GND.n529 585
R438 GND.n5825 GND.n5824 585
R439 GND.n5826 GND.n5825 585
R440 GND.n528 GND.n527 585
R441 GND.n5827 GND.n528 585
R442 GND.n5830 GND.n5829 585
R443 GND.n5829 GND.n5828 585
R444 GND.n525 GND.n524 585
R445 GND.n524 GND.n523 585
R446 GND.n5835 GND.n5834 585
R447 GND.n5836 GND.n5835 585
R448 GND.n522 GND.n521 585
R449 GND.n5837 GND.n522 585
R450 GND.n5840 GND.n5839 585
R451 GND.n5839 GND.n5838 585
R452 GND.n519 GND.n518 585
R453 GND.n518 GND.n517 585
R454 GND.n5845 GND.n5844 585
R455 GND.n5846 GND.n5845 585
R456 GND.n516 GND.n515 585
R457 GND.n5847 GND.n516 585
R458 GND.n5850 GND.n5849 585
R459 GND.n5849 GND.n5848 585
R460 GND.n513 GND.n512 585
R461 GND.n512 GND.n511 585
R462 GND.n5855 GND.n5854 585
R463 GND.n5856 GND.n5855 585
R464 GND.n510 GND.n509 585
R465 GND.n5857 GND.n510 585
R466 GND.n5860 GND.n5859 585
R467 GND.n5859 GND.n5858 585
R468 GND.n507 GND.n506 585
R469 GND.n506 GND.n505 585
R470 GND.n5865 GND.n5864 585
R471 GND.n5866 GND.n5865 585
R472 GND.n504 GND.n503 585
R473 GND.n5867 GND.n504 585
R474 GND.n5870 GND.n5869 585
R475 GND.n5869 GND.n5868 585
R476 GND.n501 GND.n500 585
R477 GND.n500 GND.n499 585
R478 GND.n5875 GND.n5874 585
R479 GND.n5876 GND.n5875 585
R480 GND.n498 GND.n497 585
R481 GND.n5877 GND.n498 585
R482 GND.n5880 GND.n5879 585
R483 GND.n5879 GND.n5878 585
R484 GND.n495 GND.n494 585
R485 GND.n494 GND.n493 585
R486 GND.n5885 GND.n5884 585
R487 GND.n5886 GND.n5885 585
R488 GND.n492 GND.n491 585
R489 GND.n5887 GND.n492 585
R490 GND.n5890 GND.n5889 585
R491 GND.n5889 GND.n5888 585
R492 GND.n489 GND.n488 585
R493 GND.n488 GND.n487 585
R494 GND.n5895 GND.n5894 585
R495 GND.n5896 GND.n5895 585
R496 GND.n486 GND.n485 585
R497 GND.n5897 GND.n486 585
R498 GND.n5900 GND.n5899 585
R499 GND.n5899 GND.n5898 585
R500 GND.n483 GND.n482 585
R501 GND.n482 GND.n481 585
R502 GND.n5905 GND.n5904 585
R503 GND.n5906 GND.n5905 585
R504 GND.n480 GND.n479 585
R505 GND.n5907 GND.n480 585
R506 GND.n5910 GND.n5909 585
R507 GND.n5909 GND.n5908 585
R508 GND.n477 GND.n476 585
R509 GND.n476 GND.n475 585
R510 GND.n5915 GND.n5914 585
R511 GND.n5916 GND.n5915 585
R512 GND.n474 GND.n473 585
R513 GND.n5917 GND.n474 585
R514 GND.n5920 GND.n5919 585
R515 GND.n5919 GND.n5918 585
R516 GND.n471 GND.n470 585
R517 GND.n470 GND.n469 585
R518 GND.n5925 GND.n5924 585
R519 GND.n5926 GND.n5925 585
R520 GND.n468 GND.n467 585
R521 GND.n5927 GND.n468 585
R522 GND.n5930 GND.n5929 585
R523 GND.n5929 GND.n5928 585
R524 GND.n465 GND.n464 585
R525 GND.n464 GND.n463 585
R526 GND.n5935 GND.n5934 585
R527 GND.n5936 GND.n5935 585
R528 GND.n462 GND.n461 585
R529 GND.n5937 GND.n462 585
R530 GND.n5940 GND.n5939 585
R531 GND.n5939 GND.n5938 585
R532 GND.n459 GND.n458 585
R533 GND.n458 GND.n457 585
R534 GND.n5945 GND.n5944 585
R535 GND.n5946 GND.n5945 585
R536 GND.n456 GND.n455 585
R537 GND.n5947 GND.n456 585
R538 GND.n5950 GND.n5949 585
R539 GND.n5949 GND.n5948 585
R540 GND.n453 GND.n452 585
R541 GND.n452 GND.n451 585
R542 GND.n5955 GND.n5954 585
R543 GND.n5956 GND.n5955 585
R544 GND.n450 GND.n449 585
R545 GND.n5957 GND.n450 585
R546 GND.n5960 GND.n5959 585
R547 GND.n5959 GND.n5958 585
R548 GND.n447 GND.n446 585
R549 GND.n446 GND.n445 585
R550 GND.n5965 GND.n5964 585
R551 GND.n5966 GND.n5965 585
R552 GND.n444 GND.n443 585
R553 GND.n5967 GND.n444 585
R554 GND.n5970 GND.n5969 585
R555 GND.n5969 GND.n5968 585
R556 GND.n441 GND.n440 585
R557 GND.n440 GND.n439 585
R558 GND.n5975 GND.n5974 585
R559 GND.n5976 GND.n5975 585
R560 GND.n438 GND.n437 585
R561 GND.n5977 GND.n438 585
R562 GND.n5980 GND.n5979 585
R563 GND.n5979 GND.n5978 585
R564 GND.n435 GND.n434 585
R565 GND.n434 GND.n433 585
R566 GND.n5985 GND.n5984 585
R567 GND.n5986 GND.n5985 585
R568 GND.n432 GND.n431 585
R569 GND.n5987 GND.n432 585
R570 GND.n5990 GND.n5989 585
R571 GND.n5989 GND.n5988 585
R572 GND.n429 GND.n428 585
R573 GND.n428 GND.n427 585
R574 GND.n5995 GND.n5994 585
R575 GND.n5996 GND.n5995 585
R576 GND.n426 GND.n425 585
R577 GND.n5997 GND.n426 585
R578 GND.n6000 GND.n5999 585
R579 GND.n5999 GND.n5998 585
R580 GND.n423 GND.n422 585
R581 GND.n422 GND.n421 585
R582 GND.n6005 GND.n6004 585
R583 GND.n6006 GND.n6005 585
R584 GND.n420 GND.n419 585
R585 GND.n6007 GND.n420 585
R586 GND.n6010 GND.n6009 585
R587 GND.n6009 GND.n6008 585
R588 GND.n417 GND.n416 585
R589 GND.n416 GND.n415 585
R590 GND.n6015 GND.n6014 585
R591 GND.n6016 GND.n6015 585
R592 GND.n414 GND.n413 585
R593 GND.n6017 GND.n414 585
R594 GND.n6020 GND.n6019 585
R595 GND.n6019 GND.n6018 585
R596 GND.n411 GND.n410 585
R597 GND.n410 GND.n409 585
R598 GND.n6025 GND.n6024 585
R599 GND.n6026 GND.n6025 585
R600 GND.n408 GND.n407 585
R601 GND.n6027 GND.n408 585
R602 GND.n6030 GND.n6029 585
R603 GND.n6029 GND.n6028 585
R604 GND.n405 GND.n404 585
R605 GND.n404 GND.n403 585
R606 GND.n6035 GND.n6034 585
R607 GND.n6036 GND.n6035 585
R608 GND.n402 GND.n401 585
R609 GND.n6037 GND.n402 585
R610 GND.n6040 GND.n6039 585
R611 GND.n6039 GND.n6038 585
R612 GND.n399 GND.n398 585
R613 GND.n398 GND.n397 585
R614 GND.n6045 GND.n6044 585
R615 GND.n6046 GND.n6045 585
R616 GND.n396 GND.n395 585
R617 GND.n6047 GND.n396 585
R618 GND.n6050 GND.n6049 585
R619 GND.n6049 GND.n6048 585
R620 GND.n393 GND.n392 585
R621 GND.n392 GND.n391 585
R622 GND.n6055 GND.n6054 585
R623 GND.n6056 GND.n6055 585
R624 GND.n390 GND.n389 585
R625 GND.n6057 GND.n390 585
R626 GND.n6060 GND.n6059 585
R627 GND.n6059 GND.n6058 585
R628 GND.n387 GND.n386 585
R629 GND.n386 GND.n385 585
R630 GND.n6065 GND.n6064 585
R631 GND.n6066 GND.n6065 585
R632 GND.n384 GND.n383 585
R633 GND.n6067 GND.n384 585
R634 GND.n6070 GND.n6069 585
R635 GND.n6069 GND.n6068 585
R636 GND.n381 GND.n380 585
R637 GND.n380 GND.n379 585
R638 GND.n6075 GND.n6074 585
R639 GND.n6076 GND.n6075 585
R640 GND.n378 GND.n377 585
R641 GND.n6077 GND.n378 585
R642 GND.n6080 GND.n6079 585
R643 GND.n6079 GND.n6078 585
R644 GND.n375 GND.n374 585
R645 GND.n374 GND.n373 585
R646 GND.n6085 GND.n6084 585
R647 GND.n6086 GND.n6085 585
R648 GND.n372 GND.n371 585
R649 GND.n6087 GND.n372 585
R650 GND.n6090 GND.n6089 585
R651 GND.n6089 GND.n6088 585
R652 GND.n369 GND.n368 585
R653 GND.n368 GND.n367 585
R654 GND.n6095 GND.n6094 585
R655 GND.n6096 GND.n6095 585
R656 GND.n366 GND.n365 585
R657 GND.n6097 GND.n366 585
R658 GND.n6100 GND.n6099 585
R659 GND.n6099 GND.n6098 585
R660 GND.n363 GND.n362 585
R661 GND.n362 GND.n361 585
R662 GND.n6105 GND.n6104 585
R663 GND.n6106 GND.n6105 585
R664 GND.n360 GND.n359 585
R665 GND.n6107 GND.n360 585
R666 GND.n6110 GND.n6109 585
R667 GND.n6109 GND.n6108 585
R668 GND.n357 GND.n356 585
R669 GND.n356 GND.n355 585
R670 GND.n6115 GND.n6114 585
R671 GND.n6116 GND.n6115 585
R672 GND.n354 GND.n353 585
R673 GND.n6117 GND.n354 585
R674 GND.n6120 GND.n6119 585
R675 GND.n6119 GND.n6118 585
R676 GND.n351 GND.n350 585
R677 GND.n350 GND.n349 585
R678 GND.n6125 GND.n6124 585
R679 GND.n6126 GND.n6125 585
R680 GND.n348 GND.n347 585
R681 GND.n6127 GND.n348 585
R682 GND.n6130 GND.n6129 585
R683 GND.n6129 GND.n6128 585
R684 GND.n345 GND.n344 585
R685 GND.n344 GND.n343 585
R686 GND.n6135 GND.n6134 585
R687 GND.n6136 GND.n6135 585
R688 GND.n342 GND.n341 585
R689 GND.n6137 GND.n342 585
R690 GND.n6140 GND.n6139 585
R691 GND.n6139 GND.n6138 585
R692 GND.n339 GND.n338 585
R693 GND.n338 GND.n337 585
R694 GND.n6145 GND.n6144 585
R695 GND.n6146 GND.n6145 585
R696 GND.n336 GND.n335 585
R697 GND.n6147 GND.n336 585
R698 GND.n6150 GND.n6149 585
R699 GND.n6149 GND.n6148 585
R700 GND.n333 GND.n332 585
R701 GND.n332 GND.n331 585
R702 GND.n6155 GND.n6154 585
R703 GND.n6156 GND.n6155 585
R704 GND.n330 GND.n329 585
R705 GND.n6157 GND.n330 585
R706 GND.n6160 GND.n6159 585
R707 GND.n6159 GND.n6158 585
R708 GND.n327 GND.n326 585
R709 GND.n326 GND.n325 585
R710 GND.n6165 GND.n6164 585
R711 GND.n6166 GND.n6165 585
R712 GND.n324 GND.n323 585
R713 GND.n6167 GND.n324 585
R714 GND.n6170 GND.n6169 585
R715 GND.n6169 GND.n6168 585
R716 GND.n321 GND.n320 585
R717 GND.n320 GND.n319 585
R718 GND.n6175 GND.n6174 585
R719 GND.n6176 GND.n6175 585
R720 GND.n318 GND.n317 585
R721 GND.n6177 GND.n318 585
R722 GND.n6180 GND.n6179 585
R723 GND.n6179 GND.n6178 585
R724 GND.n315 GND.n314 585
R725 GND.n314 GND.n313 585
R726 GND.n6185 GND.n6184 585
R727 GND.n6186 GND.n6185 585
R728 GND.n312 GND.n311 585
R729 GND.n6187 GND.n312 585
R730 GND.n6190 GND.n6189 585
R731 GND.n6189 GND.n6188 585
R732 GND.n6342 GND.n218 585
R733 GND.n218 GND.n217 585
R734 GND.n6341 GND.n6340 585
R735 GND.n6340 GND.n6339 585
R736 GND.n222 GND.n221 585
R737 GND.n6338 GND.n222 585
R738 GND.n6336 GND.n6335 585
R739 GND.n6337 GND.n6336 585
R740 GND.n225 GND.n224 585
R741 GND.n224 GND.n223 585
R742 GND.n6330 GND.n6329 585
R743 GND.n6329 GND.n6328 585
R744 GND.n228 GND.n227 585
R745 GND.n6327 GND.n228 585
R746 GND.n6325 GND.n6324 585
R747 GND.n6326 GND.n6325 585
R748 GND.n231 GND.n230 585
R749 GND.n230 GND.n229 585
R750 GND.n6320 GND.n6319 585
R751 GND.n6319 GND.n6318 585
R752 GND.n234 GND.n233 585
R753 GND.n6317 GND.n234 585
R754 GND.n6315 GND.n6314 585
R755 GND.n6316 GND.n6315 585
R756 GND.n237 GND.n236 585
R757 GND.n236 GND.n235 585
R758 GND.n6310 GND.n6309 585
R759 GND.n6309 GND.n6308 585
R760 GND.n240 GND.n239 585
R761 GND.n6307 GND.n240 585
R762 GND.n6305 GND.n6304 585
R763 GND.n6306 GND.n6305 585
R764 GND.n243 GND.n242 585
R765 GND.n242 GND.n241 585
R766 GND.n6300 GND.n6299 585
R767 GND.n6299 GND.n6298 585
R768 GND.n246 GND.n245 585
R769 GND.n6297 GND.n246 585
R770 GND.n6295 GND.n6294 585
R771 GND.n6296 GND.n6295 585
R772 GND.n249 GND.n248 585
R773 GND.n248 GND.n247 585
R774 GND.n6290 GND.n6289 585
R775 GND.n6289 GND.n6288 585
R776 GND.n252 GND.n251 585
R777 GND.n6287 GND.n252 585
R778 GND.n6285 GND.n6284 585
R779 GND.n6286 GND.n6285 585
R780 GND.n255 GND.n254 585
R781 GND.n254 GND.n253 585
R782 GND.n6280 GND.n6279 585
R783 GND.n6279 GND.n6278 585
R784 GND.n258 GND.n257 585
R785 GND.n6277 GND.n258 585
R786 GND.n6275 GND.n6274 585
R787 GND.n6276 GND.n6275 585
R788 GND.n261 GND.n260 585
R789 GND.n260 GND.n259 585
R790 GND.n6270 GND.n6269 585
R791 GND.n6269 GND.n6268 585
R792 GND.n264 GND.n263 585
R793 GND.n6267 GND.n264 585
R794 GND.n6265 GND.n6264 585
R795 GND.n6266 GND.n6265 585
R796 GND.n267 GND.n266 585
R797 GND.n266 GND.n265 585
R798 GND.n6260 GND.n6259 585
R799 GND.n6259 GND.n6258 585
R800 GND.n270 GND.n269 585
R801 GND.n6257 GND.n270 585
R802 GND.n6255 GND.n6254 585
R803 GND.n6256 GND.n6255 585
R804 GND.n273 GND.n272 585
R805 GND.n272 GND.n271 585
R806 GND.n6250 GND.n6249 585
R807 GND.n6249 GND.n6248 585
R808 GND.n276 GND.n275 585
R809 GND.n6247 GND.n276 585
R810 GND.n6245 GND.n6244 585
R811 GND.n6246 GND.n6245 585
R812 GND.n279 GND.n278 585
R813 GND.n278 GND.n277 585
R814 GND.n6240 GND.n6239 585
R815 GND.n6239 GND.n6238 585
R816 GND.n282 GND.n281 585
R817 GND.n6237 GND.n282 585
R818 GND.n6235 GND.n6234 585
R819 GND.n6236 GND.n6235 585
R820 GND.n285 GND.n284 585
R821 GND.n284 GND.n283 585
R822 GND.n6230 GND.n6229 585
R823 GND.n6229 GND.n6228 585
R824 GND.n288 GND.n287 585
R825 GND.n6227 GND.n288 585
R826 GND.n6225 GND.n6224 585
R827 GND.n6226 GND.n6225 585
R828 GND.n291 GND.n290 585
R829 GND.n290 GND.n289 585
R830 GND.n6220 GND.n6219 585
R831 GND.n6219 GND.n6218 585
R832 GND.n294 GND.n293 585
R833 GND.n6217 GND.n294 585
R834 GND.n6215 GND.n6214 585
R835 GND.n6216 GND.n6215 585
R836 GND.n297 GND.n296 585
R837 GND.n296 GND.n295 585
R838 GND.n6210 GND.n6209 585
R839 GND.n6209 GND.n6208 585
R840 GND.n300 GND.n299 585
R841 GND.n6207 GND.n300 585
R842 GND.n6205 GND.n6204 585
R843 GND.n6206 GND.n6205 585
R844 GND.n303 GND.n302 585
R845 GND.n302 GND.n301 585
R846 GND.n6200 GND.n6199 585
R847 GND.n6199 GND.n6198 585
R848 GND.n306 GND.n305 585
R849 GND.n6197 GND.n306 585
R850 GND.n6195 GND.n6194 585
R851 GND.n6196 GND.n6195 585
R852 GND.n309 GND.n308 585
R853 GND.n308 GND.n307 585
R854 GND.n4657 GND.n4656 585
R855 GND.n4656 GND.n4655 585
R856 GND.n4658 GND.n1850 585
R857 GND.n4183 GND.n1850 585
R858 GND.n4660 GND.n4659 585
R859 GND.n4661 GND.n4660 585
R860 GND.n1851 GND.n1849 585
R861 GND.n1849 GND.n1846 585
R862 GND.n1831 GND.n1830 585
R863 GND.n1834 GND.n1831 585
R864 GND.n4671 GND.n4670 585
R865 GND.n4670 GND.n4669 585
R866 GND.n4672 GND.n1823 585
R867 GND.n2285 GND.n1823 585
R868 GND.n4674 GND.n4673 585
R869 GND.n4675 GND.n4674 585
R870 GND.n1824 GND.n1822 585
R871 GND.n1822 GND.n1819 585
R872 GND.n1804 GND.n1803 585
R873 GND.n1807 GND.n1804 585
R874 GND.n4685 GND.n4684 585
R875 GND.n4684 GND.n4683 585
R876 GND.n4686 GND.n1796 585
R877 GND.n2289 GND.n1796 585
R878 GND.n4688 GND.n4687 585
R879 GND.n4689 GND.n4688 585
R880 GND.n1797 GND.n1795 585
R881 GND.n1795 GND.n1793 585
R882 GND.n1778 GND.n1777 585
R883 GND.n1781 GND.n1778 585
R884 GND.n4699 GND.n4698 585
R885 GND.n4698 GND.n4697 585
R886 GND.n4700 GND.n1770 585
R887 GND.n4152 GND.n1770 585
R888 GND.n4702 GND.n4701 585
R889 GND.n4703 GND.n4702 585
R890 GND.n1771 GND.n1769 585
R891 GND.n1769 GND.n1766 585
R892 GND.n1755 GND.n1754 585
R893 GND.n2297 GND.n1755 585
R894 GND.n4713 GND.n4712 585
R895 GND.n4712 GND.n4711 585
R896 GND.n4714 GND.n1749 585
R897 GND.n4143 GND.n1749 585
R898 GND.n4716 GND.n4715 585
R899 GND.n4717 GND.n4716 585
R900 GND.n1735 GND.n1734 585
R901 GND.n4007 GND.n1735 585
R902 GND.n4727 GND.n4726 585
R903 GND.n4726 GND.n4725 585
R904 GND.n4728 GND.n1729 585
R905 GND.n3998 GND.n1729 585
R906 GND.n4730 GND.n4729 585
R907 GND.n4731 GND.n4730 585
R908 GND.n1730 GND.n1728 585
R909 GND.n3980 GND.n1728 585
R910 GND.n2624 GND.n2623 585
R911 GND.n2625 GND.n2624 585
R912 GND.n1697 GND.n1696 585
R913 GND.n1707 GND.n1697 585
R914 GND.n4748 GND.n4747 585
R915 GND.n4747 GND.n4746 585
R916 GND.n4749 GND.n1686 585
R917 GND.n3936 GND.n1686 585
R918 GND.n4751 GND.n4750 585
R919 GND.n4752 GND.n4751 585
R920 GND.n1687 GND.n1685 585
R921 GND.n1685 GND.n1675 585
R922 GND.n1690 GND.n1689 585
R923 GND.n1689 GND.n1673 585
R924 GND.n1656 GND.n1655 585
R925 GND.n3963 GND.n1656 585
R926 GND.n4768 GND.n4767 585
R927 GND.n4767 GND.n4766 585
R928 GND.n4769 GND.n1642 585
R929 GND.n2638 GND.n1642 585
R930 GND.n4771 GND.n4770 585
R931 GND.n4772 GND.n4771 585
R932 GND.n1643 GND.n1641 585
R933 GND.n1641 GND.n1631 585
R934 GND.n1649 GND.n1648 585
R935 GND.n1648 GND.n1629 585
R936 GND.n1647 GND.n1646 585
R937 GND.n1647 GND.n1615 585
R938 GND.n1603 GND.n1602 585
R939 GND.n1613 GND.n1603 585
R940 GND.n4796 GND.n4795 585
R941 GND.n4795 GND.n4794 585
R942 GND.n4797 GND.n1592 585
R943 GND.n3905 GND.n1592 585
R944 GND.n4799 GND.n4798 585
R945 GND.n4800 GND.n4799 585
R946 GND.n1593 GND.n1591 585
R947 GND.n3876 GND.n1591 585
R948 GND.n1596 GND.n1595 585
R949 GND.n1595 GND.n1571 585
R950 GND.n1559 GND.n1558 585
R951 GND.n1569 GND.n1559 585
R952 GND.n4816 GND.n4815 585
R953 GND.n4815 GND.n4814 585
R954 GND.n4817 GND.n1548 585
R955 GND.n3852 GND.n1548 585
R956 GND.n4819 GND.n4818 585
R957 GND.n4820 GND.n4819 585
R958 GND.n1549 GND.n1547 585
R959 GND.n1547 GND.n1537 585
R960 GND.n1552 GND.n1551 585
R961 GND.n1551 GND.n1535 585
R962 GND.n1523 GND.n1522 585
R963 GND.n3838 GND.n1523 585
R964 GND.n4837 GND.n4836 585
R965 GND.n4836 GND.n4835 585
R966 GND.n4838 GND.n1517 585
R967 GND.n3800 GND.n1517 585
R968 GND.n4840 GND.n4839 585
R969 GND.n4841 GND.n4840 585
R970 GND.n1503 GND.n1502 585
R971 GND.n3809 GND.n1503 585
R972 GND.n4851 GND.n4850 585
R973 GND.n4850 GND.n4849 585
R974 GND.n4852 GND.n1497 585
R975 GND.n3792 GND.n1497 585
R976 GND.n4854 GND.n4853 585
R977 GND.n4855 GND.n4854 585
R978 GND.n1484 GND.n1483 585
R979 GND.n2682 GND.n1484 585
R980 GND.n4865 GND.n4864 585
R981 GND.n4864 GND.n4863 585
R982 GND.n4866 GND.n1478 585
R983 GND.n2685 GND.n1478 585
R984 GND.n4868 GND.n4867 585
R985 GND.n4869 GND.n4868 585
R986 GND.n1464 GND.n1463 585
R987 GND.n3726 GND.n1464 585
R988 GND.n4879 GND.n4878 585
R989 GND.n4878 GND.n4877 585
R990 GND.n4880 GND.n1458 585
R991 GND.n3743 GND.n1458 585
R992 GND.n4882 GND.n4881 585
R993 GND.n4883 GND.n4882 585
R994 GND.n1444 GND.n1443 585
R995 GND.n3711 GND.n1444 585
R996 GND.n4893 GND.n4892 585
R997 GND.n4892 GND.n4891 585
R998 GND.n4894 GND.n1438 585
R999 GND.n3703 GND.n1438 585
R1000 GND.n4896 GND.n4895 585
R1001 GND.n4897 GND.n4896 585
R1002 GND.n1424 GND.n1423 585
R1003 GND.n3664 GND.n1424 585
R1004 GND.n4907 GND.n4906 585
R1005 GND.n4906 GND.n4905 585
R1006 GND.n4908 GND.n1416 585
R1007 GND.n3656 GND.n1416 585
R1008 GND.n4910 GND.n4909 585
R1009 GND.n4911 GND.n4910 585
R1010 GND.n1417 GND.n1415 585
R1011 GND.n3561 GND.n1415 585
R1012 GND.n1398 GND.n1397 585
R1013 GND.n1401 GND.n1398 585
R1014 GND.n4921 GND.n4920 585
R1015 GND.n4920 GND.n4919 585
R1016 GND.n4922 GND.n1390 585
R1017 GND.n3552 GND.n1390 585
R1018 GND.n4924 GND.n4923 585
R1019 GND.n4925 GND.n4924 585
R1020 GND.n1391 GND.n1389 585
R1021 GND.n1389 GND.n1386 585
R1022 GND.n1371 GND.n1370 585
R1023 GND.n1374 GND.n1371 585
R1024 GND.n4935 GND.n4934 585
R1025 GND.n4934 GND.n4933 585
R1026 GND.n4936 GND.n1363 585
R1027 GND.n2823 GND.n1363 585
R1028 GND.n4938 GND.n4937 585
R1029 GND.n4939 GND.n4938 585
R1030 GND.n1364 GND.n1362 585
R1031 GND.n1362 GND.n1359 585
R1032 GND.n1344 GND.n1343 585
R1033 GND.n1347 GND.n1344 585
R1034 GND.n4949 GND.n4948 585
R1035 GND.n4948 GND.n4947 585
R1036 GND.n4950 GND.n1336 585
R1037 GND.n2826 GND.n1336 585
R1038 GND.n4952 GND.n4951 585
R1039 GND.n4953 GND.n4952 585
R1040 GND.n1337 GND.n1335 585
R1041 GND.n1335 GND.n1332 585
R1042 GND.n1311 GND.n1310 585
R1043 GND.n1314 GND.n1311 585
R1044 GND.n4963 GND.n4962 585
R1045 GND.n4962 GND.n4961 585
R1046 GND.n4964 GND.n1304 585
R1047 GND.n3521 GND.n1304 585
R1048 GND.n4966 GND.n4965 585
R1049 GND.n4967 GND.n4966 585
R1050 GND.n1305 GND.n1231 585
R1051 GND.n4969 GND.n1231 585
R1052 GND.n5032 GND.n5031 585
R1053 GND.n1232 GND.n1230 585
R1054 GND.n5028 GND.n5027 585
R1055 GND.n5029 GND.n5028 585
R1056 GND.n1249 GND.n1248 585
R1057 GND.n5020 GND.n1258 585
R1058 GND.n5019 GND.n1259 585
R1059 GND.n1266 GND.n1260 585
R1060 GND.n5012 GND.n1267 585
R1061 GND.n5011 GND.n1268 585
R1062 GND.n1270 GND.n1269 585
R1063 GND.n3470 GND.n3469 585
R1064 GND.n3474 GND.n3471 585
R1065 GND.n3477 GND.n3476 585
R1066 GND.n3475 GND.n2841 585
R1067 GND.n3482 GND.n3481 585
R1068 GND.n3484 GND.n3483 585
R1069 GND.n3487 GND.n3486 585
R1070 GND.n3485 GND.n2839 585
R1071 GND.n3492 GND.n3491 585
R1072 GND.n3494 GND.n3493 585
R1073 GND.n3497 GND.n3496 585
R1074 GND.n3495 GND.n2837 585
R1075 GND.n3502 GND.n3501 585
R1076 GND.n3504 GND.n3503 585
R1077 GND.n3507 GND.n3506 585
R1078 GND.n3505 GND.n2835 585
R1079 GND.n3512 GND.n3511 585
R1080 GND.n3514 GND.n3513 585
R1081 GND.n3516 GND.n3515 585
R1082 GND.n4191 GND.n4190 585
R1083 GND.n4188 GND.n2280 585
R1084 GND.n4195 GND.n2279 585
R1085 GND.n4196 GND.n2277 585
R1086 GND.n4197 GND.n2274 585
R1087 GND.n2272 GND.n2270 585
R1088 GND.n4201 GND.n2269 585
R1089 GND.n4202 GND.n2267 585
R1090 GND.n4203 GND.n2266 585
R1091 GND.n2264 GND.n2262 585
R1092 GND.n4207 GND.n2261 585
R1093 GND.n4208 GND.n2259 585
R1094 GND.n4209 GND.n2258 585
R1095 GND.n2256 GND.n2254 585
R1096 GND.n4213 GND.n2253 585
R1097 GND.n4214 GND.n2251 585
R1098 GND.n4215 GND.n2250 585
R1099 GND.n2491 GND.n2249 585
R1100 GND.n2494 GND.n2492 585
R1101 GND.n2495 GND.n2488 585
R1102 GND.n2487 GND.n2479 585
R1103 GND.n2507 GND.n2478 585
R1104 GND.n2508 GND.n2477 585
R1105 GND.n2475 GND.n2466 585
R1106 GND.n2515 GND.n2465 585
R1107 GND.n2516 GND.n2463 585
R1108 GND.n2462 GND.n2450 585
R1109 GND.n2523 GND.n2449 585
R1110 GND.n2524 GND.n1857 585
R1111 GND.n1871 GND.n1857 585
R1112 GND.n4186 GND.n1859 585
R1113 GND.n4655 GND.n1859 585
R1114 GND.n4185 GND.n4184 585
R1115 GND.n4184 GND.n4183 585
R1116 GND.n4182 GND.n1847 585
R1117 GND.n4661 GND.n1847 585
R1118 GND.n4176 GND.n2282 585
R1119 GND.n4176 GND.n1846 585
R1120 GND.n4178 GND.n4177 585
R1121 GND.n4177 GND.n1834 585
R1122 GND.n4175 GND.n1833 585
R1123 GND.n4669 GND.n1833 585
R1124 GND.n4174 GND.n2286 585
R1125 GND.n2286 GND.n2285 585
R1126 GND.n2284 GND.n1820 585
R1127 GND.n4675 GND.n1820 585
R1128 GND.n4170 GND.n4169 585
R1129 GND.n4169 GND.n1819 585
R1130 GND.n4168 GND.n4167 585
R1131 GND.n4168 GND.n1807 585
R1132 GND.n4166 GND.n1806 585
R1133 GND.n4683 GND.n1806 585
R1134 GND.n2291 GND.n2290 585
R1135 GND.n2290 GND.n2289 585
R1136 GND.n4162 GND.n1794 585
R1137 GND.n4689 GND.n1794 585
R1138 GND.n4161 GND.n4160 585
R1139 GND.n4160 GND.n1793 585
R1140 GND.n4159 GND.n4158 585
R1141 GND.n4159 GND.n1781 585
R1142 GND.n2293 GND.n1780 585
R1143 GND.n4697 GND.n1780 585
R1144 GND.n4154 GND.n4153 585
R1145 GND.n4153 GND.n4152 585
R1146 GND.n4151 GND.n1767 585
R1147 GND.n4703 GND.n1767 585
R1148 GND.n4150 GND.n2299 585
R1149 GND.n2299 GND.n1766 585
R1150 GND.n2298 GND.n2295 585
R1151 GND.n2298 GND.n2297 585
R1152 GND.n4146 GND.n1756 585
R1153 GND.n4711 GND.n1756 585
R1154 GND.n4145 GND.n4144 585
R1155 GND.n4144 GND.n4143 585
R1156 GND.n2301 GND.n1747 585
R1157 GND.n4717 GND.n1747 585
R1158 GND.n4006 GND.n4005 585
R1159 GND.n4007 GND.n4006 585
R1160 GND.n2609 GND.n1737 585
R1161 GND.n4725 GND.n1737 585
R1162 GND.n4000 GND.n3999 585
R1163 GND.n3999 GND.n3998 585
R1164 GND.n2611 GND.n1726 585
R1165 GND.n4731 GND.n1726 585
R1166 GND.n3979 GND.n3978 585
R1167 GND.n3980 GND.n3979 585
R1168 GND.n2627 GND.n2626 585
R1169 GND.n2626 GND.n2625 585
R1170 GND.n3974 GND.n3973 585
R1171 GND.n3973 GND.n1707 585
R1172 GND.n3972 GND.n1699 585
R1173 GND.n4746 GND.n1699 585
R1174 GND.n3971 GND.n2630 585
R1175 GND.n3936 GND.n2630 585
R1176 GND.n2629 GND.n1683 585
R1177 GND.n4752 GND.n1683 585
R1178 GND.n3967 GND.n3966 585
R1179 GND.n3966 GND.n1675 585
R1180 GND.n3965 GND.n2632 585
R1181 GND.n3965 GND.n1673 585
R1182 GND.n3964 GND.n2633 585
R1183 GND.n3964 GND.n3963 585
R1184 GND.n3891 GND.n1658 585
R1185 GND.n4766 GND.n1658 585
R1186 GND.n3892 GND.n3888 585
R1187 GND.n3888 GND.n2638 585
R1188 GND.n3893 GND.n1639 585
R1189 GND.n4772 GND.n1639 585
R1190 GND.n3886 GND.n3885 585
R1191 GND.n3885 GND.n1631 585
R1192 GND.n3897 GND.n3884 585
R1193 GND.n3884 GND.n1629 585
R1194 GND.n3898 GND.n3883 585
R1195 GND.n3883 GND.n1615 585
R1196 GND.n3899 GND.n3882 585
R1197 GND.n3882 GND.n1613 585
R1198 GND.n2647 GND.n1605 585
R1199 GND.n4794 GND.n1605 585
R1200 GND.n3904 GND.n3903 585
R1201 GND.n3905 GND.n3904 585
R1202 GND.n2646 GND.n1589 585
R1203 GND.n4800 GND.n1589 585
R1204 GND.n3878 GND.n3877 585
R1205 GND.n3877 GND.n3876 585
R1206 GND.n2650 GND.n2649 585
R1207 GND.n2650 GND.n1571 585
R1208 GND.n3846 GND.n3845 585
R1209 GND.n3845 GND.n1569 585
R1210 GND.n2659 GND.n1562 585
R1211 GND.n4814 GND.n1562 585
R1212 GND.n3851 GND.n3850 585
R1213 GND.n3852 GND.n3851 585
R1214 GND.n2658 GND.n1545 585
R1215 GND.n4820 GND.n1545 585
R1216 GND.n3842 GND.n3841 585
R1217 GND.n3841 GND.n1537 585
R1218 GND.n3840 GND.n2661 585
R1219 GND.n3840 GND.n1535 585
R1220 GND.n3839 GND.n2662 585
R1221 GND.n3839 GND.n3838 585
R1222 GND.n3802 GND.n1525 585
R1223 GND.n4835 GND.n1525 585
R1224 GND.n3803 GND.n3801 585
R1225 GND.n3801 GND.n3800 585
R1226 GND.n2671 GND.n1515 585
R1227 GND.n4841 GND.n1515 585
R1228 GND.n3808 GND.n3807 585
R1229 GND.n3809 GND.n3808 585
R1230 GND.n2670 GND.n1505 585
R1231 GND.n4849 GND.n1505 585
R1232 GND.n3794 GND.n3793 585
R1233 GND.n3793 GND.n3792 585
R1234 GND.n2673 GND.n1495 585
R1235 GND.n4855 GND.n1495 585
R1236 GND.n3731 GND.n3730 585
R1237 GND.n3730 GND.n2682 585
R1238 GND.n3729 GND.n1486 585
R1239 GND.n4863 GND.n1486 585
R1240 GND.n3735 GND.n3728 585
R1241 GND.n3728 GND.n2685 585
R1242 GND.n3736 GND.n1476 585
R1243 GND.n4869 GND.n1476 585
R1244 GND.n3737 GND.n3727 585
R1245 GND.n3727 GND.n3726 585
R1246 GND.n2698 GND.n1466 585
R1247 GND.n4877 GND.n1466 585
R1248 GND.n3742 GND.n3741 585
R1249 GND.n3743 GND.n3742 585
R1250 GND.n2697 GND.n1456 585
R1251 GND.n4883 GND.n1456 585
R1252 GND.n3710 GND.n3709 585
R1253 GND.n3711 GND.n3710 585
R1254 GND.n2703 GND.n1446 585
R1255 GND.n4891 GND.n1446 585
R1256 GND.n3705 GND.n3704 585
R1257 GND.n3704 GND.n3703 585
R1258 GND.n2705 GND.n1436 585
R1259 GND.n4897 GND.n1436 585
R1260 GND.n3663 GND.n3662 585
R1261 GND.n3664 GND.n3663 585
R1262 GND.n2709 GND.n1426 585
R1263 GND.n4905 GND.n1426 585
R1264 GND.n3658 GND.n3657 585
R1265 GND.n3657 GND.n3656 585
R1266 GND.n2711 GND.n1413 585
R1267 GND.n4911 GND.n1413 585
R1268 GND.n3560 GND.n3559 585
R1269 GND.n3561 GND.n3560 585
R1270 GND.n2818 GND.n2817 585
R1271 GND.n2817 GND.n1401 585
R1272 GND.n3555 GND.n1400 585
R1273 GND.n4919 GND.n1400 585
R1274 GND.n3554 GND.n3553 585
R1275 GND.n3553 GND.n3552 585
R1276 GND.n3551 GND.n1387 585
R1277 GND.n4925 GND.n1387 585
R1278 GND.n3545 GND.n2820 585
R1279 GND.n3545 GND.n1386 585
R1280 GND.n3547 GND.n3546 585
R1281 GND.n3546 GND.n1374 585
R1282 GND.n3544 GND.n1373 585
R1283 GND.n4933 GND.n1373 585
R1284 GND.n3543 GND.n2824 585
R1285 GND.n2824 GND.n2823 585
R1286 GND.n2822 GND.n1360 585
R1287 GND.n4939 GND.n1360 585
R1288 GND.n3539 GND.n3538 585
R1289 GND.n3538 GND.n1359 585
R1290 GND.n3537 GND.n3536 585
R1291 GND.n3537 GND.n1347 585
R1292 GND.n3535 GND.n1346 585
R1293 GND.n4947 GND.n1346 585
R1294 GND.n2828 GND.n2827 585
R1295 GND.n2827 GND.n2826 585
R1296 GND.n3531 GND.n1333 585
R1297 GND.n4953 GND.n1333 585
R1298 GND.n3530 GND.n3529 585
R1299 GND.n3529 GND.n1332 585
R1300 GND.n3528 GND.n3527 585
R1301 GND.n3528 GND.n1314 585
R1302 GND.n2830 GND.n1313 585
R1303 GND.n4961 GND.n1313 585
R1304 GND.n3523 GND.n3522 585
R1305 GND.n3522 GND.n3521 585
R1306 GND.n3520 GND.n1302 585
R1307 GND.n4967 GND.n1302 585
R1308 GND.n3519 GND.n1301 585
R1309 GND.n4969 GND.n1301 585
R1310 GND.n3460 GND.n1169 585
R1311 GND.n5100 GND.n1169 585
R1312 GND.n3462 GND.n3461 585
R1313 GND.n3463 GND.n3462 585
R1314 GND.n3459 GND.n1160 585
R1315 GND.n3459 GND.n3458 585
R1316 GND.n2846 GND.n1159 585
R1317 GND.n3439 GND.n2846 585
R1318 GND.n3449 GND.n1158 585
R1319 GND.n3450 GND.n3449 585
R1320 GND.n3448 GND.n2857 585
R1321 GND.n3448 GND.n3447 585
R1322 GND.n2856 GND.n1152 585
R1323 GND.n2870 GND.n2856 585
R1324 GND.n2868 GND.n1151 585
R1325 GND.n3432 GND.n2868 585
R1326 GND.n3419 GND.n1150 585
R1327 GND.n3419 GND.n3418 585
R1328 GND.n3421 GND.n3420 585
R1329 GND.n3422 GND.n3421 585
R1330 GND.n3417 GND.n1144 585
R1331 GND.n3417 GND.n3416 585
R1332 GND.n2879 GND.n1143 585
R1333 GND.n3355 GND.n2879 585
R1334 GND.n2888 GND.n1142 585
R1335 GND.n3407 GND.n2888 585
R1336 GND.n3395 GND.n3393 585
R1337 GND.n3395 GND.n3394 585
R1338 GND.n3396 GND.n1136 585
R1339 GND.n3397 GND.n3396 585
R1340 GND.n3392 GND.n1135 585
R1341 GND.n3392 GND.n3391 585
R1342 GND.n2898 GND.n1134 585
R1343 GND.n2911 GND.n2898 585
R1344 GND.n2909 GND.n2908 585
R1345 GND.n3382 GND.n2909 585
R1346 GND.n3370 GND.n1128 585
R1347 GND.n3370 GND.n3369 585
R1348 GND.n3371 GND.n1127 585
R1349 GND.n3372 GND.n3371 585
R1350 GND.n2921 GND.n1126 585
R1351 GND.n3301 GND.n2921 585
R1352 GND.n2938 GND.n2937 585
R1353 GND.n2938 GND.n2928 585
R1354 GND.n2939 GND.n1120 585
R1355 GND.n3292 GND.n2939 585
R1356 GND.n2976 GND.n1119 585
R1357 GND.n3251 GND.n2976 585
R1358 GND.n3264 GND.n1118 585
R1359 GND.n3264 GND.n3263 585
R1360 GND.n3266 GND.n3265 585
R1361 GND.n3267 GND.n3266 585
R1362 GND.n2968 GND.n1112 585
R1363 GND.n3272 GND.n2968 585
R1364 GND.n2967 GND.n1111 585
R1365 GND.n2967 GND.n2964 585
R1366 GND.n2955 GND.n1110 585
R1367 GND.n3239 GND.n2955 585
R1368 GND.n3282 GND.n2956 585
R1369 GND.n3282 GND.n3281 585
R1370 GND.n3283 GND.n1104 585
R1371 GND.n3284 GND.n3283 585
R1372 GND.n2954 GND.n1103 585
R1373 GND.n3229 GND.n2954 585
R1374 GND.n2992 GND.n1102 585
R1375 GND.n2992 GND.n2983 585
R1376 GND.n2994 GND.n2993 585
R1377 GND.n3215 GND.n2994 585
R1378 GND.n3203 GND.n1096 585
R1379 GND.n3203 GND.n3202 585
R1380 GND.n3204 GND.n1095 585
R1381 GND.n3205 GND.n3204 585
R1382 GND.n3005 GND.n1094 585
R1383 GND.n3192 GND.n3005 585
R1384 GND.n3023 GND.n3022 585
R1385 GND.n3023 GND.n3011 585
R1386 GND.n3024 GND.n1088 585
R1387 GND.n3180 GND.n3024 585
R1388 GND.n3168 GND.n1087 585
R1389 GND.n3168 GND.n3019 585
R1390 GND.n3169 GND.n1086 585
R1391 GND.n3170 GND.n3169 585
R1392 GND.n3167 GND.n3035 585
R1393 GND.n3167 GND.n3166 585
R1394 GND.n3034 GND.n1080 585
R1395 GND.n3142 GND.n3034 585
R1396 GND.n3046 GND.n1079 585
R1397 GND.n3152 GND.n3046 585
R1398 GND.n3139 GND.n1078 585
R1399 GND.n3140 GND.n3139 585
R1400 GND.n1058 GND.n1056 585
R1401 GND.n3115 GND.n1056 585
R1402 GND.n5173 GND.n5172 585
R1403 GND.n5174 GND.n5173 585
R1404 GND.n1057 GND.n1055 585
R1405 GND.n3107 GND.n1055 585
R1406 GND.n1071 GND.n1036 585
R1407 GND.n5180 GND.n1036 585
R1408 GND.n1070 GND.n1069 585
R1409 GND.n1069 GND.n1033 585
R1410 GND.n1068 GND.n1012 585
R1411 GND.n1018 GND.n1012 585
R1412 GND.n5189 GND.n1013 585
R1413 GND.n5189 GND.n5188 585
R1414 GND.n5191 GND.n5190 585
R1415 GND.n3068 GND.n1011 585
R1416 GND.n3071 GND.n3069 585
R1417 GND.n3073 GND.n3072 585
R1418 GND.n3075 GND.n3074 585
R1419 GND.n3065 GND.n3064 585
R1420 GND.n3079 GND.n3066 585
R1421 GND.n3081 GND.n3080 585
R1422 GND.n3083 GND.n3082 585
R1423 GND.n3061 GND.n3060 585
R1424 GND.n3087 GND.n3062 585
R1425 GND.n3089 GND.n3088 585
R1426 GND.n3091 GND.n3090 585
R1427 GND.n3057 GND.n3056 585
R1428 GND.n3095 GND.n3058 585
R1429 GND.n3096 GND.n3053 585
R1430 GND.n3097 GND.n966 585
R1431 GND.n5264 GND.n966 585
R1432 GND.n5007 GND.n5006 585
R1433 GND.n5008 GND.n1274 585
R1434 GND.n1289 GND.n1264 585
R1435 GND.n5015 GND.n1263 585
R1436 GND.n5016 GND.n1262 585
R1437 GND.n1287 GND.n1256 585
R1438 GND.n5023 GND.n1255 585
R1439 GND.n5024 GND.n1254 585
R1440 GND.n1284 GND.n1253 585
R1441 GND.n1283 GND.n1282 585
R1442 GND.n1281 GND.n1228 585
R1443 GND.n5036 GND.n1227 585
R1444 GND.n5037 GND.n1226 585
R1445 GND.n1278 GND.n1224 585
R1446 GND.n5041 GND.n1223 585
R1447 GND.n5042 GND.n1222 585
R1448 GND.n5043 GND.n1221 585
R1449 GND.n5004 GND.n1221 585
R1450 GND.n3466 GND.n1167 585
R1451 GND.n5100 GND.n1167 585
R1452 GND.n3465 GND.n3464 585
R1453 GND.n3464 GND.n3463 585
R1454 GND.n2844 GND.n2843 585
R1455 GND.n3458 GND.n2844 585
R1456 GND.n3441 GND.n3440 585
R1457 GND.n3440 GND.n3439 585
R1458 GND.n2861 GND.n2854 585
R1459 GND.n3450 GND.n2854 585
R1460 GND.n3446 GND.n3445 585
R1461 GND.n3447 GND.n3446 585
R1462 GND.n2860 GND.n2859 585
R1463 GND.n2870 GND.n2859 585
R1464 GND.n3434 GND.n3433 585
R1465 GND.n3433 GND.n3432 585
R1466 GND.n2864 GND.n2863 585
R1467 GND.n3418 GND.n2864 585
R1468 GND.n2883 GND.n2877 585
R1469 GND.n3422 GND.n2877 585
R1470 GND.n3415 GND.n3414 585
R1471 GND.n3416 GND.n3415 585
R1472 GND.n2882 GND.n2881 585
R1473 GND.n3355 GND.n2881 585
R1474 GND.n3409 GND.n3408 585
R1475 GND.n3408 GND.n3407 585
R1476 GND.n2886 GND.n2885 585
R1477 GND.n3394 GND.n2886 585
R1478 GND.n2903 GND.n2896 585
R1479 GND.n3397 GND.n2896 585
R1480 GND.n3390 GND.n3389 585
R1481 GND.n3391 GND.n3390 585
R1482 GND.n2902 GND.n2901 585
R1483 GND.n2911 GND.n2901 585
R1484 GND.n3384 GND.n3383 585
R1485 GND.n3383 GND.n3382 585
R1486 GND.n2906 GND.n2905 585
R1487 GND.n3369 GND.n2906 585
R1488 GND.n2931 GND.n2919 585
R1489 GND.n3372 GND.n2919 585
R1490 GND.n3300 GND.n3299 585
R1491 GND.n3301 GND.n3300 585
R1492 GND.n2930 GND.n2929 585
R1493 GND.n2929 GND.n2928 585
R1494 GND.n3294 GND.n3293 585
R1495 GND.n3293 GND.n3292 585
R1496 GND.n2934 GND.n2933 585
R1497 GND.n3251 GND.n2934 585
R1498 GND.n3249 GND.n3248 585
R1499 GND.n3263 GND.n3249 585
R1500 GND.n2977 GND.n2974 585
R1501 GND.n3267 GND.n2974 585
R1502 GND.n3243 GND.n2965 585
R1503 GND.n3272 GND.n2965 585
R1504 GND.n3242 GND.n3241 585
R1505 GND.n3241 GND.n2964 585
R1506 GND.n3240 GND.n3236 585
R1507 GND.n3240 GND.n3239 585
R1508 GND.n2979 GND.n2957 585
R1509 GND.n3281 GND.n2957 585
R1510 GND.n3232 GND.n2952 585
R1511 GND.n3284 GND.n2952 585
R1512 GND.n3231 GND.n3230 585
R1513 GND.n3230 GND.n3229 585
R1514 GND.n2982 GND.n2981 585
R1515 GND.n2983 GND.n2982 585
R1516 GND.n3007 GND.n2990 585
R1517 GND.n3215 GND.n2990 585
R1518 GND.n3201 GND.n3200 585
R1519 GND.n3202 GND.n3201 585
R1520 GND.n3006 GND.n3003 585
R1521 GND.n3205 GND.n3003 585
R1522 GND.n3194 GND.n3193 585
R1523 GND.n3193 GND.n3192 585
R1524 GND.n3010 GND.n3009 585
R1525 GND.n3011 GND.n3010 585
R1526 GND.n3159 GND.n3020 585
R1527 GND.n3180 GND.n3020 585
R1528 GND.n3160 GND.n3158 585
R1529 GND.n3158 GND.n3019 585
R1530 GND.n3039 GND.n3032 585
R1531 GND.n3170 GND.n3032 585
R1532 GND.n3165 GND.n3164 585
R1533 GND.n3166 GND.n3165 585
R1534 GND.n3038 GND.n3037 585
R1535 GND.n3142 GND.n3037 585
R1536 GND.n3154 GND.n3153 585
R1537 GND.n3153 GND.n3152 585
R1538 GND.n3042 GND.n3041 585
R1539 GND.n3140 GND.n3042 585
R1540 GND.n3114 GND.n3113 585
R1541 GND.n3115 GND.n3114 585
R1542 GND.n3047 GND.n1053 585
R1543 GND.n5174 GND.n1053 585
R1544 GND.n3109 GND.n3108 585
R1545 GND.n3108 GND.n3107 585
R1546 GND.n3104 GND.n1035 585
R1547 GND.n5180 GND.n1035 585
R1548 GND.n3103 GND.n3051 585
R1549 GND.n3051 GND.n1033 585
R1550 GND.n3050 GND.n3049 585
R1551 GND.n3050 GND.n1018 585
R1552 GND.n3099 GND.n1017 585
R1553 GND.n5188 GND.n1017 585
R1554 GND.n5099 GND.n5098 585
R1555 GND.n5100 GND.n5099 585
R1556 GND.n1172 GND.n1170 585
R1557 GND.n3463 GND.n1170 585
R1558 GND.n3457 GND.n3456 585
R1559 GND.n3458 GND.n3457 585
R1560 GND.n2849 GND.n2848 585
R1561 GND.n3439 GND.n2848 585
R1562 GND.n3452 GND.n3451 585
R1563 GND.n3451 GND.n3450 585
R1564 GND.n2852 GND.n2851 585
R1565 GND.n3447 GND.n2852 585
R1566 GND.n3429 GND.n2871 585
R1567 GND.n2871 GND.n2870 585
R1568 GND.n3431 GND.n3430 585
R1569 GND.n3432 GND.n3431 585
R1570 GND.n2872 GND.n2869 585
R1571 GND.n3418 GND.n2869 585
R1572 GND.n3424 GND.n3423 585
R1573 GND.n3423 GND.n3422 585
R1574 GND.n2875 GND.n2874 585
R1575 GND.n3416 GND.n2875 585
R1576 GND.n3404 GND.n2890 585
R1577 GND.n3355 GND.n2890 585
R1578 GND.n3406 GND.n3405 585
R1579 GND.n3407 GND.n3406 585
R1580 GND.n2891 GND.n2889 585
R1581 GND.n3394 GND.n2889 585
R1582 GND.n3399 GND.n3398 585
R1583 GND.n3398 GND.n3397 585
R1584 GND.n2894 GND.n2893 585
R1585 GND.n3391 GND.n2894 585
R1586 GND.n3379 GND.n2912 585
R1587 GND.n2912 GND.n2911 585
R1588 GND.n3381 GND.n3380 585
R1589 GND.n3382 GND.n3381 585
R1590 GND.n2913 GND.n2910 585
R1591 GND.n3369 GND.n2910 585
R1592 GND.n3374 GND.n3373 585
R1593 GND.n3373 GND.n3372 585
R1594 GND.n2916 GND.n2915 585
R1595 GND.n3301 GND.n2916 585
R1596 GND.n3289 GND.n2941 585
R1597 GND.n2941 GND.n2928 585
R1598 GND.n3291 GND.n3290 585
R1599 GND.n3292 GND.n3291 585
R1600 GND.n2971 GND.n2940 585
R1601 GND.n3251 GND.n2940 585
R1602 GND.n2973 GND.n2972 585
R1603 GND.n3263 GND.n2973 585
R1604 GND.n3269 GND.n3268 585
R1605 GND.n3268 GND.n3267 585
R1606 GND.n3271 GND.n3270 585
R1607 GND.n3272 GND.n3271 585
R1608 GND.n2970 GND.n2969 585
R1609 GND.n2970 GND.n2964 585
R1610 GND.n3238 GND.n2946 585
R1611 GND.n3239 GND.n3238 585
R1612 GND.n2950 GND.n2947 585
R1613 GND.n3281 GND.n2950 585
R1614 GND.n3286 GND.n3285 585
R1615 GND.n3285 GND.n3284 585
R1616 GND.n2949 GND.n2948 585
R1617 GND.n3229 GND.n2949 585
R1618 GND.n3212 GND.n2996 585
R1619 GND.n2996 GND.n2983 585
R1620 GND.n3214 GND.n3213 585
R1621 GND.n3215 GND.n3214 585
R1622 GND.n2997 GND.n2995 585
R1623 GND.n3202 GND.n2995 585
R1624 GND.n3207 GND.n3206 585
R1625 GND.n3206 GND.n3205 585
R1626 GND.n3000 GND.n2999 585
R1627 GND.n3192 GND.n3000 585
R1628 GND.n3177 GND.n3026 585
R1629 GND.n3026 GND.n3011 585
R1630 GND.n3179 GND.n3178 585
R1631 GND.n3180 GND.n3179 585
R1632 GND.n3027 GND.n3025 585
R1633 GND.n3025 GND.n3019 585
R1634 GND.n3172 GND.n3171 585
R1635 GND.n3171 GND.n3170 585
R1636 GND.n3030 GND.n3029 585
R1637 GND.n3166 GND.n3030 585
R1638 GND.n3149 GND.n3143 585
R1639 GND.n3143 GND.n3142 585
R1640 GND.n3151 GND.n3150 585
R1641 GND.n3152 GND.n3151 585
R1642 GND.n3144 GND.n3141 585
R1643 GND.n3141 GND.n3140 585
R1644 GND.n1050 GND.n1049 585
R1645 GND.n3115 GND.n1050 585
R1646 GND.n5176 GND.n5175 585
R1647 GND.n5175 GND.n5174 585
R1648 GND.n5177 GND.n1038 585
R1649 GND.n3107 GND.n1038 585
R1650 GND.n5179 GND.n5178 585
R1651 GND.n5180 GND.n5179 585
R1652 GND.n1039 GND.n1037 585
R1653 GND.n1037 GND.n1033 585
R1654 GND.n1043 GND.n1042 585
R1655 GND.n1042 GND.n1018 585
R1656 GND.n1041 GND.n970 585
R1657 GND.n5188 GND.n970 585
R1658 GND.n5262 GND.n5261 585
R1659 GND.n5260 GND.n969 585
R1660 GND.n5259 GND.n968 585
R1661 GND.n5264 GND.n968 585
R1662 GND.n5258 GND.n5257 585
R1663 GND.n5256 GND.n5255 585
R1664 GND.n5254 GND.n5253 585
R1665 GND.n5252 GND.n5251 585
R1666 GND.n5250 GND.n5249 585
R1667 GND.n5248 GND.n5247 585
R1668 GND.n5246 GND.n5245 585
R1669 GND.n5244 GND.n5243 585
R1670 GND.n5242 GND.n5241 585
R1671 GND.n5240 GND.n5239 585
R1672 GND.n5238 GND.n5237 585
R1673 GND.n5236 GND.n5235 585
R1674 GND.n5234 GND.n5233 585
R1675 GND.n5231 GND.n5230 585
R1676 GND.n5229 GND.n5228 585
R1677 GND.n5227 GND.n5226 585
R1678 GND.n5225 GND.n5224 585
R1679 GND.n5223 GND.n5222 585
R1680 GND.n5221 GND.n5220 585
R1681 GND.n5219 GND.n5218 585
R1682 GND.n5217 GND.n5216 585
R1683 GND.n5215 GND.n5214 585
R1684 GND.n5213 GND.n5212 585
R1685 GND.n5211 GND.n5210 585
R1686 GND.n5209 GND.n5208 585
R1687 GND.n5207 GND.n5206 585
R1688 GND.n5205 GND.n5204 585
R1689 GND.n5203 GND.n5202 585
R1690 GND.n5201 GND.n5200 585
R1691 GND.n5199 GND.n5198 585
R1692 GND.n5197 GND.n5196 585
R1693 GND.n1015 GND.n1006 585
R1694 GND.n5046 GND.n1165 585
R1695 GND.n4979 GND.n1219 585
R1696 GND.n5050 GND.n1216 585
R1697 GND.n5051 GND.n1215 585
R1698 GND.n5052 GND.n1214 585
R1699 GND.n4982 GND.n1212 585
R1700 GND.n5056 GND.n1211 585
R1701 GND.n5057 GND.n1210 585
R1702 GND.n5058 GND.n1209 585
R1703 GND.n4985 GND.n1207 585
R1704 GND.n5062 GND.n1206 585
R1705 GND.n5063 GND.n1205 585
R1706 GND.n5064 GND.n1204 585
R1707 GND.n4988 GND.n1202 585
R1708 GND.n5068 GND.n1201 585
R1709 GND.n5069 GND.n1200 585
R1710 GND.n5070 GND.n1199 585
R1711 GND.n4991 GND.n1197 585
R1712 GND.n5074 GND.n1196 585
R1713 GND.n5076 GND.n1190 585
R1714 GND.n5077 GND.n1189 585
R1715 GND.n4995 GND.n1187 585
R1716 GND.n5081 GND.n1186 585
R1717 GND.n5082 GND.n1185 585
R1718 GND.n5083 GND.n1184 585
R1719 GND.n4998 GND.n1182 585
R1720 GND.n5087 GND.n1181 585
R1721 GND.n5088 GND.n1180 585
R1722 GND.n5089 GND.n1179 585
R1723 GND.n5001 GND.n1177 585
R1724 GND.n5093 GND.n1176 585
R1725 GND.n5094 GND.n1175 585
R1726 GND.n5095 GND.n1171 585
R1727 GND.n5004 GND.n1171 585
R1728 GND.n5102 GND.n5101 585
R1729 GND.n5101 GND.n5100 585
R1730 GND.n5103 GND.n1163 585
R1731 GND.n3463 GND.n1163 585
R1732 GND.n5104 GND.n1162 585
R1733 GND.n3458 GND.n1162 585
R1734 GND.n3438 GND.n1157 585
R1735 GND.n3439 GND.n3438 585
R1736 GND.n5108 GND.n1156 585
R1737 GND.n3450 GND.n1156 585
R1738 GND.n5109 GND.n1155 585
R1739 GND.n3447 GND.n1155 585
R1740 GND.n5110 GND.n1154 585
R1741 GND.n2870 GND.n1154 585
R1742 GND.n2866 GND.n1149 585
R1743 GND.n3432 GND.n2866 585
R1744 GND.n5114 GND.n1148 585
R1745 GND.n3418 GND.n1148 585
R1746 GND.n5115 GND.n1147 585
R1747 GND.n3422 GND.n1147 585
R1748 GND.n5116 GND.n1146 585
R1749 GND.n3416 GND.n1146 585
R1750 GND.n3354 GND.n1141 585
R1751 GND.n3355 GND.n3354 585
R1752 GND.n5120 GND.n1140 585
R1753 GND.n3407 GND.n1140 585
R1754 GND.n5121 GND.n1139 585
R1755 GND.n3394 GND.n1139 585
R1756 GND.n5122 GND.n1138 585
R1757 GND.n3397 GND.n1138 585
R1758 GND.n2900 GND.n1133 585
R1759 GND.n3391 GND.n2900 585
R1760 GND.n5126 GND.n1132 585
R1761 GND.n2911 GND.n1132 585
R1762 GND.n5127 GND.n1131 585
R1763 GND.n3382 GND.n1131 585
R1764 GND.n5128 GND.n1130 585
R1765 GND.n3369 GND.n1130 585
R1766 GND.n2918 GND.n1125 585
R1767 GND.n3372 GND.n2918 585
R1768 GND.n5132 GND.n1124 585
R1769 GND.n3301 GND.n1124 585
R1770 GND.n5133 GND.n1123 585
R1771 GND.n2928 GND.n1123 585
R1772 GND.n5134 GND.n1122 585
R1773 GND.n3292 GND.n1122 585
R1774 GND.n3250 GND.n1117 585
R1775 GND.n3251 GND.n3250 585
R1776 GND.n5138 GND.n1116 585
R1777 GND.n3263 GND.n1116 585
R1778 GND.n5139 GND.n1115 585
R1779 GND.n3267 GND.n1115 585
R1780 GND.n5140 GND.n1114 585
R1781 GND.n3272 GND.n1114 585
R1782 GND.n2963 GND.n1109 585
R1783 GND.n2964 GND.n2963 585
R1784 GND.n5144 GND.n1108 585
R1785 GND.n3239 GND.n1108 585
R1786 GND.n5145 GND.n1107 585
R1787 GND.n3281 GND.n1107 585
R1788 GND.n5146 GND.n1106 585
R1789 GND.n3284 GND.n1106 585
R1790 GND.n3228 GND.n1101 585
R1791 GND.n3229 GND.n3228 585
R1792 GND.n5150 GND.n1100 585
R1793 GND.n2983 GND.n1100 585
R1794 GND.n5151 GND.n1099 585
R1795 GND.n3215 GND.n1099 585
R1796 GND.n5152 GND.n1098 585
R1797 GND.n3202 GND.n1098 585
R1798 GND.n3002 GND.n1093 585
R1799 GND.n3205 GND.n3002 585
R1800 GND.n5156 GND.n1092 585
R1801 GND.n3192 GND.n1092 585
R1802 GND.n5157 GND.n1091 585
R1803 GND.n3011 GND.n1091 585
R1804 GND.n5158 GND.n1090 585
R1805 GND.n3180 GND.n1090 585
R1806 GND.n3018 GND.n1085 585
R1807 GND.n3019 GND.n3018 585
R1808 GND.n5162 GND.n1084 585
R1809 GND.n3170 GND.n1084 585
R1810 GND.n5163 GND.n1083 585
R1811 GND.n3166 GND.n1083 585
R1812 GND.n5164 GND.n1082 585
R1813 GND.n3142 GND.n1082 585
R1814 GND.n3044 GND.n1077 585
R1815 GND.n3152 GND.n3044 585
R1816 GND.n5168 GND.n1076 585
R1817 GND.n3140 GND.n1076 585
R1818 GND.n5169 GND.n1075 585
R1819 GND.n3115 GND.n1075 585
R1820 GND.n5170 GND.n1052 585
R1821 GND.n5174 GND.n1052 585
R1822 GND.n3106 GND.n1074 585
R1823 GND.n3107 GND.n3106 585
R1824 GND.n1073 GND.n1034 585
R1825 GND.n5180 GND.n1034 585
R1826 GND.n1064 GND.n1061 585
R1827 GND.n1064 GND.n1033 585
R1828 GND.n1066 GND.n1065 585
R1829 GND.n1065 GND.n1018 585
R1830 GND.n1063 GND.n1016 585
R1831 GND.n5188 GND.n1016 585
R1832 GND.n6501 GND.n6500 585
R1833 GND.n6502 GND.n6501 585
R1834 GND.n85 GND.n83 585
R1835 GND.n4554 GND.n83 585
R1836 GND.n4550 GND.n4549 585
R1837 GND.n4551 GND.n4550 585
R1838 GND.n2058 GND.n2057 585
R1839 GND.n2063 GND.n2057 585
R1840 GND.n4545 GND.n4544 585
R1841 GND.n4544 GND.n4543 585
R1842 GND.n2061 GND.n2060 585
R1843 GND.n4539 GND.n2061 585
R1844 GND.n4508 GND.n2079 585
R1845 GND.n2079 GND.n2068 585
R1846 GND.n4510 GND.n4509 585
R1847 GND.n4511 GND.n4510 585
R1848 GND.n2080 GND.n2078 585
R1849 GND.n2078 GND.n2075 585
R1850 GND.n4503 GND.n4502 585
R1851 GND.n4502 GND.n4501 585
R1852 GND.n2083 GND.n2082 585
R1853 GND.n4496 GND.n2083 585
R1854 GND.n4479 GND.n2099 585
R1855 GND.n2099 GND.n2087 585
R1856 GND.n4481 GND.n4480 585
R1857 GND.n4482 GND.n4481 585
R1858 GND.n2100 GND.n2098 585
R1859 GND.n2098 GND.n2094 585
R1860 GND.n4474 GND.n4473 585
R1861 GND.n4473 GND.n4472 585
R1862 GND.n2103 GND.n2102 585
R1863 GND.n4468 GND.n2103 585
R1864 GND.n4453 GND.n2123 585
R1865 GND.n2123 GND.n2110 585
R1866 GND.n4455 GND.n4454 585
R1867 GND.n4456 GND.n4455 585
R1868 GND.n2124 GND.n2122 585
R1869 GND.n2122 GND.n2119 585
R1870 GND.n4448 GND.n4447 585
R1871 GND.n4447 GND.n4446 585
R1872 GND.n2127 GND.n2126 585
R1873 GND.n4442 GND.n2127 585
R1874 GND.n4390 GND.n4388 585
R1875 GND.n4388 GND.n2132 585
R1876 GND.n4392 GND.n4391 585
R1877 GND.n4393 GND.n4392 585
R1878 GND.n4379 GND.n4378 585
R1879 GND.n4402 GND.n4379 585
R1880 GND.n4408 GND.n4407 585
R1881 GND.n4407 GND.n4406 585
R1882 GND.n4410 GND.n4375 585
R1883 GND.n4382 GND.n4375 585
R1884 GND.n4412 GND.n4411 585
R1885 GND.n4413 GND.n4412 585
R1886 GND.n4376 GND.n4374 585
R1887 GND.n4374 GND.n2164 585
R1888 GND.n2156 GND.n2155 585
R1889 GND.n4420 GND.n2156 585
R1890 GND.n4425 GND.n4424 585
R1891 GND.n4424 GND.n4423 585
R1892 GND.n4427 GND.n2152 585
R1893 GND.n4362 GND.n2152 585
R1894 GND.n4429 GND.n4428 585
R1895 GND.n4430 GND.n4429 585
R1896 GND.n2153 GND.n2151 585
R1897 GND.n2151 GND.n2147 585
R1898 GND.n4353 GND.n4352 585
R1899 GND.n4354 GND.n4353 585
R1900 GND.n2184 GND.n2183 585
R1901 GND.n4342 GND.n2183 585
R1902 GND.n4347 GND.n4346 585
R1903 GND.n4346 GND.n4345 585
R1904 GND.n2187 GND.n2186 585
R1905 GND.n4339 GND.n2187 585
R1906 GND.n4327 GND.n2206 585
R1907 GND.n2206 GND.n2205 585
R1908 GND.n4329 GND.n4328 585
R1909 GND.n4330 GND.n4329 585
R1910 GND.n2207 GND.n2204 585
R1911 GND.n4316 GND.n2204 585
R1912 GND.n4322 GND.n4321 585
R1913 GND.n4321 GND.n4320 585
R1914 GND.n2210 GND.n2209 585
R1915 GND.n4314 GND.n2210 585
R1916 GND.n4302 GND.n2228 585
R1917 GND.n2228 GND.n2227 585
R1918 GND.n4304 GND.n4303 585
R1919 GND.n4305 GND.n4304 585
R1920 GND.n2229 GND.n2225 585
R1921 GND.n4292 GND.n2225 585
R1922 GND.n4297 GND.n4296 585
R1923 GND.n4296 GND.n4295 585
R1924 GND.n2232 GND.n2231 585
R1925 GND.n4289 GND.n2232 585
R1926 GND.n4225 GND.n4224 585
R1927 GND.n4226 GND.n4225 585
R1928 GND.n1891 GND.n1890 585
R1929 GND.n4280 GND.n1891 585
R1930 GND.n4635 GND.n4634 585
R1931 GND.n4634 GND.n4633 585
R1932 GND.n4636 GND.n1886 585
R1933 GND.n2245 GND.n1886 585
R1934 GND.n4638 GND.n4637 585
R1935 GND.n4639 GND.n4638 585
R1936 GND.n2369 GND.n1885 585
R1937 GND.n2368 GND.n2367 585
R1938 GND.n2374 GND.n2373 585
R1939 GND.n2376 GND.n2365 585
R1940 GND.n2379 GND.n2378 585
R1941 GND.n2363 GND.n2362 585
R1942 GND.n2384 GND.n2383 585
R1943 GND.n2386 GND.n2361 585
R1944 GND.n2389 GND.n2388 585
R1945 GND.n2359 GND.n2358 585
R1946 GND.n2394 GND.n2393 585
R1947 GND.n2396 GND.n2357 585
R1948 GND.n2401 GND.n2400 585
R1949 GND.n2398 GND.n2354 585
R1950 GND.n2397 GND.n1872 585
R1951 GND.n2580 GND.n2579 585
R1952 GND.n2577 GND.n2408 585
R1953 GND.n2575 GND.n2574 585
R1954 GND.n2573 GND.n2409 585
R1955 GND.n2572 GND.n2571 585
R1956 GND.n2569 GND.n2414 585
R1957 GND.n2567 GND.n2566 585
R1958 GND.n2565 GND.n2415 585
R1959 GND.n2564 GND.n2563 585
R1960 GND.n2561 GND.n2420 585
R1961 GND.n2559 GND.n2558 585
R1962 GND.n2557 GND.n2421 585
R1963 GND.n2556 GND.n2555 585
R1964 GND.n2553 GND.n2426 585
R1965 GND.n2551 GND.n2550 585
R1966 GND.n2549 GND.n2427 585
R1967 GND.n2548 GND.n2547 585
R1968 GND.n2545 GND.n2434 585
R1969 GND.n2543 GND.n2542 585
R1970 GND.n6447 GND.n6446 585
R1971 GND.n6448 GND.n133 585
R1972 GND.n6449 GND.n130 585
R1973 GND.n6420 GND.n128 585
R1974 GND.n6453 GND.n127 585
R1975 GND.n6454 GND.n126 585
R1976 GND.n6455 GND.n125 585
R1977 GND.n6423 GND.n123 585
R1978 GND.n6459 GND.n122 585
R1979 GND.n6460 GND.n121 585
R1980 GND.n6461 GND.n120 585
R1981 GND.n6426 GND.n118 585
R1982 GND.n6465 GND.n117 585
R1983 GND.n6466 GND.n116 585
R1984 GND.n6467 GND.n115 585
R1985 GND.n6429 GND.n113 585
R1986 GND.n6471 GND.n112 585
R1987 GND.n6472 GND.n111 585
R1988 GND.n6473 GND.n110 585
R1989 GND.n6432 GND.n105 585
R1990 GND.n6477 GND.n104 585
R1991 GND.n6478 GND.n103 585
R1992 GND.n6479 GND.n102 585
R1993 GND.n6435 GND.n100 585
R1994 GND.n6483 GND.n99 585
R1995 GND.n6484 GND.n98 585
R1996 GND.n6485 GND.n97 585
R1997 GND.n6438 GND.n95 585
R1998 GND.n6489 GND.n94 585
R1999 GND.n6490 GND.n93 585
R2000 GND.n6491 GND.n92 585
R2001 GND.n6441 GND.n90 585
R2002 GND.n6495 GND.n89 585
R2003 GND.n6496 GND.n88 585
R2004 GND.n6497 GND.n84 585
R2005 GND.n6444 GND.n84 585
R2006 GND.n4556 GND.n80 585
R2007 GND.n6502 GND.n80 585
R2008 GND.n4557 GND.n4555 585
R2009 GND.n4555 GND.n4554 585
R2010 GND.n2052 GND.n1993 585
R2011 GND.n4551 GND.n2052 585
R2012 GND.n4561 GND.n1992 585
R2013 GND.n2063 GND.n1992 585
R2014 GND.n4562 GND.n1991 585
R2015 GND.n4543 GND.n1991 585
R2016 GND.n4563 GND.n1990 585
R2017 GND.n4539 GND.n1990 585
R2018 GND.n2066 GND.n1985 585
R2019 GND.n2068 GND.n2066 585
R2020 GND.n4567 GND.n1984 585
R2021 GND.n4511 GND.n1984 585
R2022 GND.n4568 GND.n1983 585
R2023 GND.n2075 GND.n1983 585
R2024 GND.n4569 GND.n1982 585
R2025 GND.n4501 GND.n1982 585
R2026 GND.n4494 GND.n1977 585
R2027 GND.n4496 GND.n4494 585
R2028 GND.n4573 GND.n1976 585
R2029 GND.n2087 GND.n1976 585
R2030 GND.n4574 GND.n1975 585
R2031 GND.n4482 GND.n1975 585
R2032 GND.n4575 GND.n1974 585
R2033 GND.n2094 GND.n1974 585
R2034 GND.n2105 GND.n1969 585
R2035 GND.n4472 GND.n2105 585
R2036 GND.n4579 GND.n1968 585
R2037 GND.n4468 GND.n1968 585
R2038 GND.n4580 GND.n1967 585
R2039 GND.n2110 GND.n1967 585
R2040 GND.n4581 GND.n1966 585
R2041 GND.n4456 GND.n1966 585
R2042 GND.n2117 GND.n1961 585
R2043 GND.n2119 GND.n2117 585
R2044 GND.n4585 GND.n1960 585
R2045 GND.n4446 GND.n1960 585
R2046 GND.n4586 GND.n1959 585
R2047 GND.n4442 GND.n1959 585
R2048 GND.n4587 GND.n1958 585
R2049 GND.n2132 GND.n1958 585
R2050 GND.n4385 GND.n1953 585
R2051 GND.n4393 GND.n4385 585
R2052 GND.n4591 GND.n1952 585
R2053 GND.n4402 GND.n1952 585
R2054 GND.n4592 GND.n1951 585
R2055 GND.n4406 GND.n1951 585
R2056 GND.n4593 GND.n1950 585
R2057 GND.n4382 GND.n1950 585
R2058 GND.n2170 GND.n1945 585
R2059 GND.n4413 GND.n2170 585
R2060 GND.n4597 GND.n1944 585
R2061 GND.n2164 GND.n1944 585
R2062 GND.n4598 GND.n1943 585
R2063 GND.n4420 GND.n1943 585
R2064 GND.n4599 GND.n1942 585
R2065 GND.n4423 GND.n1942 585
R2066 GND.n4361 GND.n1937 585
R2067 GND.n4362 GND.n4361 585
R2068 GND.n4603 GND.n1936 585
R2069 GND.n4430 GND.n1936 585
R2070 GND.n4604 GND.n1935 585
R2071 GND.n2147 GND.n1935 585
R2072 GND.n4605 GND.n1934 585
R2073 GND.n4354 GND.n1934 585
R2074 GND.n4341 GND.n1929 585
R2075 GND.n4342 GND.n4341 585
R2076 GND.n4609 GND.n1928 585
R2077 GND.n4345 GND.n1928 585
R2078 GND.n4610 GND.n1927 585
R2079 GND.n4339 GND.n1927 585
R2080 GND.n4611 GND.n1926 585
R2081 GND.n2205 GND.n1926 585
R2082 GND.n2201 GND.n1921 585
R2083 GND.n4330 GND.n2201 585
R2084 GND.n4615 GND.n1920 585
R2085 GND.n4316 GND.n1920 585
R2086 GND.n4616 GND.n1919 585
R2087 GND.n4320 GND.n1919 585
R2088 GND.n4617 GND.n1918 585
R2089 GND.n4314 GND.n1918 585
R2090 GND.n2226 GND.n1913 585
R2091 GND.n2227 GND.n2226 585
R2092 GND.n4621 GND.n1912 585
R2093 GND.n4305 GND.n1912 585
R2094 GND.n4622 GND.n1911 585
R2095 GND.n4292 GND.n1911 585
R2096 GND.n4623 GND.n1910 585
R2097 GND.n4295 GND.n1910 585
R2098 GND.n2238 GND.n1905 585
R2099 GND.n4289 GND.n2238 585
R2100 GND.n4627 GND.n1904 585
R2101 GND.n4226 GND.n1904 585
R2102 GND.n4628 GND.n1903 585
R2103 GND.n4280 GND.n1903 585
R2104 GND.n4629 GND.n1893 585
R2105 GND.n4633 GND.n1893 585
R2106 GND.n2244 GND.n1902 585
R2107 GND.n2245 GND.n2244 585
R2108 GND.n2437 GND.n1881 585
R2109 GND.n4639 GND.n1881 585
R2110 GND.n4140 GND.n4139 585
R2111 GND.n4141 GND.n4140 585
R2112 GND.n2321 GND.n2319 585
R2113 GND.n2319 GND.n2317 585
R2114 GND.n1744 GND.n1743 585
R2115 GND.n1748 GND.n1744 585
R2116 GND.n4720 GND.n4719 585
R2117 GND.n4719 GND.n4718 585
R2118 GND.n4721 GND.n1741 585
R2119 GND.n4008 GND.n1741 585
R2120 GND.n4723 GND.n4722 585
R2121 GND.n4724 GND.n4723 585
R2122 GND.n1742 GND.n1740 585
R2123 GND.n3997 GND.n1740 585
R2124 GND.n3983 GND.n3982 585
R2125 GND.n3983 GND.n2613 585
R2126 GND.n3985 GND.n3984 585
R2127 GND.n3984 GND.n1727 585
R2128 GND.n3986 GND.n3981 585
R2129 GND.n3981 GND.n1725 585
R2130 GND.n3988 GND.n3987 585
R2131 GND.n3989 GND.n3988 585
R2132 GND.n1706 GND.n1705 585
R2133 GND.n2619 GND.n1706 585
R2134 GND.n4741 GND.n4740 585
R2135 GND.n4740 GND.n4739 585
R2136 GND.n4742 GND.n1703 585
R2137 GND.n3929 GND.n1703 585
R2138 GND.n4744 GND.n4743 585
R2139 GND.n4745 GND.n4744 585
R2140 GND.n1704 GND.n1702 585
R2141 GND.n3935 GND.n1702 585
R2142 GND.n1680 GND.n1679 585
R2143 GND.n3937 GND.n1680 585
R2144 GND.n4754 GND.n4753 585
R2145 GND.n4753 GND.n4752 585
R2146 GND.n4755 GND.n1677 585
R2147 GND.n3941 GND.n1677 585
R2148 GND.n4757 GND.n4756 585
R2149 GND.n4758 GND.n4757 585
R2150 GND.n1678 GND.n1676 585
R2151 GND.n3945 GND.n1676 585
R2152 GND.n3961 GND.n3960 585
R2153 GND.n3962 GND.n3961 585
R2154 GND.n3959 GND.n2636 585
R2155 GND.n2636 GND.n1659 585
R2156 GND.n3958 GND.n3957 585
R2157 GND.n3957 GND.n1657 585
R2158 GND.n3956 GND.n2637 585
R2159 GND.n3956 GND.n3955 585
R2160 GND.n1636 GND.n1635 585
R2161 GND.n2639 GND.n1636 585
R2162 GND.n4775 GND.n4774 585
R2163 GND.n4774 GND.n4773 585
R2164 GND.n4776 GND.n1633 585
R2165 GND.n3922 GND.n1633 585
R2166 GND.n4778 GND.n4777 585
R2167 GND.n4779 GND.n4778 585
R2168 GND.n1634 GND.n1632 585
R2169 GND.n3918 GND.n1632 585
R2170 GND.n1612 GND.n1611 585
R2171 GND.n3916 GND.n1612 585
R2172 GND.n4789 GND.n4788 585
R2173 GND.n4788 GND.n4787 585
R2174 GND.n4790 GND.n1609 585
R2175 GND.n3910 GND.n1609 585
R2176 GND.n4792 GND.n4791 585
R2177 GND.n4793 GND.n4792 585
R2178 GND.n1610 GND.n1608 585
R2179 GND.n3906 GND.n1608 585
R2180 GND.n3869 GND.n3868 585
R2181 GND.n3869 GND.n2645 585
R2182 GND.n3871 GND.n3870 585
R2183 GND.n3870 GND.n1590 585
R2184 GND.n3872 GND.n3867 585
R2185 GND.n3867 GND.n1588 585
R2186 GND.n3874 GND.n3873 585
R2187 GND.n3875 GND.n3874 585
R2188 GND.n1568 GND.n1567 585
R2189 GND.n2652 GND.n1568 585
R2190 GND.n4810 GND.n4809 585
R2191 GND.n4809 GND.n4808 585
R2192 GND.n4811 GND.n1565 585
R2193 GND.n3857 GND.n1565 585
R2194 GND.n4813 GND.n4812 585
R2195 GND.n4814 GND.n4813 585
R2196 GND.n1566 GND.n1564 585
R2197 GND.n3853 GND.n1564 585
R2198 GND.n1542 GND.n1541 585
R2199 GND.n2657 GND.n1542 585
R2200 GND.n4823 GND.n4822 585
R2201 GND.n4822 GND.n4821 585
R2202 GND.n4824 GND.n1539 585
R2203 GND.n3816 GND.n1539 585
R2204 GND.n4826 GND.n4825 585
R2205 GND.n4827 GND.n4826 585
R2206 GND.n1540 GND.n1538 585
R2207 GND.n3820 GND.n1538 585
R2208 GND.n3836 GND.n3835 585
R2209 GND.n3837 GND.n3836 585
R2210 GND.n3834 GND.n2665 585
R2211 GND.n2665 GND.n1526 585
R2212 GND.n3833 GND.n3832 585
R2213 GND.n3832 GND.n1524 585
R2214 GND.n3831 GND.n2666 585
R2215 GND.n3831 GND.n3830 585
R2216 GND.n1512 GND.n1511 585
R2217 GND.n3799 GND.n1512 585
R2218 GND.n4844 GND.n4843 585
R2219 GND.n4843 GND.n4842 585
R2220 GND.n4845 GND.n1509 585
R2221 GND.n3810 GND.n1509 585
R2222 GND.n4847 GND.n4846 585
R2223 GND.n4848 GND.n4847 585
R2224 GND.n1510 GND.n1508 585
R2225 GND.n1508 GND.n1504 585
R2226 GND.n3790 GND.n3789 585
R2227 GND.n3791 GND.n3790 585
R2228 GND.n1493 GND.n1492 585
R2229 GND.n1496 GND.n1493 585
R2230 GND.n4858 GND.n4857 585
R2231 GND.n4857 GND.n4856 585
R2232 GND.n4859 GND.n1490 585
R2233 GND.n3770 GND.n1490 585
R2234 GND.n4861 GND.n4860 585
R2235 GND.n4862 GND.n4861 585
R2236 GND.n1491 GND.n1489 585
R2237 GND.n1489 GND.n1485 585
R2238 GND.n3756 GND.n3755 585
R2239 GND.n3757 GND.n3756 585
R2240 GND.n1473 GND.n1472 585
R2241 GND.n1477 GND.n1473 585
R2242 GND.n4872 GND.n4871 585
R2243 GND.n4871 GND.n4870 585
R2244 GND.n4873 GND.n1470 585
R2245 GND.n3726 GND.n1470 585
R2246 GND.n4875 GND.n4874 585
R2247 GND.n4876 GND.n4875 585
R2248 GND.n1471 GND.n1469 585
R2249 GND.n1469 GND.n1465 585
R2250 GND.n2695 GND.n2694 585
R2251 GND.n2696 GND.n2695 585
R2252 GND.n1453 GND.n1452 585
R2253 GND.n1457 GND.n1453 585
R2254 GND.n4886 GND.n4885 585
R2255 GND.n4885 GND.n4884 585
R2256 GND.n4887 GND.n1450 585
R2257 GND.n3712 GND.n1450 585
R2258 GND.n4889 GND.n4888 585
R2259 GND.n4890 GND.n4889 585
R2260 GND.n1451 GND.n1449 585
R2261 GND.n1449 GND.n1445 585
R2262 GND.n3674 GND.n3673 585
R2263 GND.n3675 GND.n3674 585
R2264 GND.n1433 GND.n1432 585
R2265 GND.n1437 GND.n1433 585
R2266 GND.n4900 GND.n4899 585
R2267 GND.n4899 GND.n4898 585
R2268 GND.n4901 GND.n1430 585
R2269 GND.n3665 GND.n1430 585
R2270 GND.n4903 GND.n4902 585
R2271 GND.n4904 GND.n4903 585
R2272 GND.n1431 GND.n1429 585
R2273 GND.n3655 GND.n1429 585
R2274 GND.n3572 GND.n3571 585
R2275 GND.n3572 GND.n2713 585
R2276 GND.n3574 GND.n3573 585
R2277 GND.n3573 GND.n1414 585
R2278 GND.n3575 GND.n3565 585
R2279 GND.n3565 GND.n1412 585
R2280 GND.n3644 GND.n3643 585
R2281 GND.n3642 GND.n3564 585
R2282 GND.n3641 GND.n3563 585
R2283 GND.n3646 GND.n3563 585
R2284 GND.n3640 GND.n3639 585
R2285 GND.n3638 GND.n3637 585
R2286 GND.n3636 GND.n3635 585
R2287 GND.n3634 GND.n3633 585
R2288 GND.n3632 GND.n3631 585
R2289 GND.n3630 GND.n3629 585
R2290 GND.n3628 GND.n3627 585
R2291 GND.n3626 GND.n3625 585
R2292 GND.n3624 GND.n3623 585
R2293 GND.n3622 GND.n3621 585
R2294 GND.n3620 GND.n3619 585
R2295 GND.n3618 GND.n3617 585
R2296 GND.n3616 GND.n3615 585
R2297 GND.n3614 GND.n3613 585
R2298 GND.n3612 GND.n3611 585
R2299 GND.n3610 GND.n3609 585
R2300 GND.n3608 GND.n3607 585
R2301 GND.n3606 GND.n3605 585
R2302 GND.n3604 GND.n3603 585
R2303 GND.n3602 GND.n3601 585
R2304 GND.n3600 GND.n3599 585
R2305 GND.n3598 GND.n3597 585
R2306 GND.n3596 GND.n3595 585
R2307 GND.n3594 GND.n3593 585
R2308 GND.n3592 GND.n3591 585
R2309 GND.n3590 GND.n3589 585
R2310 GND.n3588 GND.n3587 585
R2311 GND.n3585 GND.n3584 585
R2312 GND.n3583 GND.n3582 585
R2313 GND.n3581 GND.n3580 585
R2314 GND.n3579 GND.n1195 585
R2315 GND.n2755 GND.n2754 585
R2316 GND.n2757 GND.n2756 585
R2317 GND.n2759 GND.n2758 585
R2318 GND.n2761 GND.n2760 585
R2319 GND.n2763 GND.n2762 585
R2320 GND.n2765 GND.n2764 585
R2321 GND.n2767 GND.n2766 585
R2322 GND.n2769 GND.n2768 585
R2323 GND.n2771 GND.n2770 585
R2324 GND.n2773 GND.n2772 585
R2325 GND.n2775 GND.n2774 585
R2326 GND.n2777 GND.n2776 585
R2327 GND.n2779 GND.n2778 585
R2328 GND.n2781 GND.n2780 585
R2329 GND.n2783 GND.n2782 585
R2330 GND.n2785 GND.n2784 585
R2331 GND.n2787 GND.n2786 585
R2332 GND.n2789 GND.n2788 585
R2333 GND.n2791 GND.n2790 585
R2334 GND.n2793 GND.n2792 585
R2335 GND.n2795 GND.n2794 585
R2336 GND.n2797 GND.n2796 585
R2337 GND.n2799 GND.n2798 585
R2338 GND.n2801 GND.n2800 585
R2339 GND.n2803 GND.n2802 585
R2340 GND.n2805 GND.n2804 585
R2341 GND.n2807 GND.n2806 585
R2342 GND.n2809 GND.n2808 585
R2343 GND.n2811 GND.n2810 585
R2344 GND.n2812 GND.n2750 585
R2345 GND.n2815 GND.n2814 585
R2346 GND.n2813 GND.n2717 585
R2347 GND.n3648 GND.n2716 585
R2348 GND.n4019 GND.n4018 585
R2349 GND.n4020 GND.n2607 585
R2350 GND.n4022 GND.n4021 585
R2351 GND.n4024 GND.n2605 585
R2352 GND.n4026 GND.n4025 585
R2353 GND.n4027 GND.n2604 585
R2354 GND.n4029 GND.n4028 585
R2355 GND.n4031 GND.n2602 585
R2356 GND.n4033 GND.n4032 585
R2357 GND.n4034 GND.n2601 585
R2358 GND.n4036 GND.n4035 585
R2359 GND.n4038 GND.n2599 585
R2360 GND.n4040 GND.n4039 585
R2361 GND.n4041 GND.n2598 585
R2362 GND.n4043 GND.n4042 585
R2363 GND.n4045 GND.n2596 585
R2364 GND.n4047 GND.n4046 585
R2365 GND.n4048 GND.n2595 585
R2366 GND.n4050 GND.n4049 585
R2367 GND.n4052 GND.n2593 585
R2368 GND.n4054 GND.n4053 585
R2369 GND.n4055 GND.n2592 585
R2370 GND.n4057 GND.n4056 585
R2371 GND.n4059 GND.n2590 585
R2372 GND.n4061 GND.n4060 585
R2373 GND.n4062 GND.n2589 585
R2374 GND.n4064 GND.n4063 585
R2375 GND.n4066 GND.n2587 585
R2376 GND.n4068 GND.n4067 585
R2377 GND.n4069 GND.n2584 585
R2378 GND.n4072 GND.n4071 585
R2379 GND.n4074 GND.n2583 585
R2380 GND.n4075 GND.n2353 585
R2381 GND.n4078 GND.n2352 585
R2382 GND.n4080 GND.n4079 585
R2383 GND.n4082 GND.n2350 585
R2384 GND.n4084 GND.n4083 585
R2385 GND.n4086 GND.n2347 585
R2386 GND.n4088 GND.n4087 585
R2387 GND.n4090 GND.n2345 585
R2388 GND.n4092 GND.n4091 585
R2389 GND.n4093 GND.n2344 585
R2390 GND.n4095 GND.n4094 585
R2391 GND.n4097 GND.n2342 585
R2392 GND.n4099 GND.n4098 585
R2393 GND.n4100 GND.n2341 585
R2394 GND.n4102 GND.n4101 585
R2395 GND.n4104 GND.n2339 585
R2396 GND.n4106 GND.n4105 585
R2397 GND.n4107 GND.n2338 585
R2398 GND.n4109 GND.n4108 585
R2399 GND.n4111 GND.n2336 585
R2400 GND.n4113 GND.n4112 585
R2401 GND.n4114 GND.n2335 585
R2402 GND.n4116 GND.n4115 585
R2403 GND.n4118 GND.n2333 585
R2404 GND.n4120 GND.n4119 585
R2405 GND.n4121 GND.n2332 585
R2406 GND.n4123 GND.n4122 585
R2407 GND.n4125 GND.n2330 585
R2408 GND.n4127 GND.n4126 585
R2409 GND.n4128 GND.n2329 585
R2410 GND.n4130 GND.n4129 585
R2411 GND.n4132 GND.n2328 585
R2412 GND.n4133 GND.n2327 585
R2413 GND.n4136 GND.n4135 585
R2414 GND.n4137 GND.n2320 585
R2415 GND.n2320 GND.n1757 585
R2416 GND.n4016 GND.n2318 585
R2417 GND.n4141 GND.n2318 585
R2418 GND.n4015 GND.n4014 585
R2419 GND.n4014 GND.n2317 585
R2420 GND.n4013 GND.n4012 585
R2421 GND.n4013 GND.n1748 585
R2422 GND.n4011 GND.n1746 585
R2423 GND.n4718 GND.n1746 585
R2424 GND.n4010 GND.n4009 585
R2425 GND.n4009 GND.n4008 585
R2426 GND.n2608 GND.n1738 585
R2427 GND.n4724 GND.n1738 585
R2428 GND.n3996 GND.n3995 585
R2429 GND.n3997 GND.n3996 585
R2430 GND.n3994 GND.n2614 585
R2431 GND.n2614 GND.n2613 585
R2432 GND.n3993 GND.n3992 585
R2433 GND.n3992 GND.n1727 585
R2434 GND.n3991 GND.n2615 585
R2435 GND.n3991 GND.n1725 585
R2436 GND.n3990 GND.n2617 585
R2437 GND.n3990 GND.n3989 585
R2438 GND.n3927 GND.n2616 585
R2439 GND.n2619 GND.n2616 585
R2440 GND.n3928 GND.n1708 585
R2441 GND.n4739 GND.n1708 585
R2442 GND.n3931 GND.n3930 585
R2443 GND.n3930 GND.n3929 585
R2444 GND.n3932 GND.n1700 585
R2445 GND.n4745 GND.n1700 585
R2446 GND.n3934 GND.n3933 585
R2447 GND.n3935 GND.n3934 585
R2448 GND.n3939 GND.n3938 585
R2449 GND.n3938 GND.n3937 585
R2450 GND.n3940 GND.n1682 585
R2451 GND.n4752 GND.n1682 585
R2452 GND.n3943 GND.n3942 585
R2453 GND.n3942 GND.n3941 585
R2454 GND.n3944 GND.n1674 585
R2455 GND.n4758 GND.n1674 585
R2456 GND.n3947 GND.n3946 585
R2457 GND.n3946 GND.n3945 585
R2458 GND.n3948 GND.n2634 585
R2459 GND.n3962 GND.n2634 585
R2460 GND.n3950 GND.n3949 585
R2461 GND.n3949 GND.n1659 585
R2462 GND.n3951 GND.n2641 585
R2463 GND.n2641 GND.n1657 585
R2464 GND.n3953 GND.n3952 585
R2465 GND.n3955 GND.n3953 585
R2466 GND.n3926 GND.n2640 585
R2467 GND.n2640 GND.n2639 585
R2468 GND.n3925 GND.n1638 585
R2469 GND.n4773 GND.n1638 585
R2470 GND.n3924 GND.n3923 585
R2471 GND.n3923 GND.n3922 585
R2472 GND.n3921 GND.n1630 585
R2473 GND.n4779 GND.n1630 585
R2474 GND.n3920 GND.n3919 585
R2475 GND.n3919 GND.n3918 585
R2476 GND.n3915 GND.n3914 585
R2477 GND.n3916 GND.n3915 585
R2478 GND.n3913 GND.n1614 585
R2479 GND.n4787 GND.n1614 585
R2480 GND.n3912 GND.n3911 585
R2481 GND.n3911 GND.n3910 585
R2482 GND.n3909 GND.n1606 585
R2483 GND.n4793 GND.n1606 585
R2484 GND.n3908 GND.n3907 585
R2485 GND.n3907 GND.n3906 585
R2486 GND.n2643 GND.n2642 585
R2487 GND.n2645 GND.n2643 585
R2488 GND.n3863 GND.n3862 585
R2489 GND.n3862 GND.n1590 585
R2490 GND.n3864 GND.n2654 585
R2491 GND.n2654 GND.n1588 585
R2492 GND.n3866 GND.n3865 585
R2493 GND.n3875 GND.n3866 585
R2494 GND.n3861 GND.n2653 585
R2495 GND.n2653 GND.n2652 585
R2496 GND.n3860 GND.n1570 585
R2497 GND.n4808 GND.n1570 585
R2498 GND.n3859 GND.n3858 585
R2499 GND.n3858 GND.n3857 585
R2500 GND.n3856 GND.n1561 585
R2501 GND.n4814 GND.n1561 585
R2502 GND.n3855 GND.n3854 585
R2503 GND.n3854 GND.n3853 585
R2504 GND.n2656 GND.n2655 585
R2505 GND.n2657 GND.n2656 585
R2506 GND.n3815 GND.n1544 585
R2507 GND.n4821 GND.n1544 585
R2508 GND.n3818 GND.n3817 585
R2509 GND.n3817 GND.n3816 585
R2510 GND.n3819 GND.n1536 585
R2511 GND.n4827 GND.n1536 585
R2512 GND.n3822 GND.n3821 585
R2513 GND.n3821 GND.n3820 585
R2514 GND.n3823 GND.n2663 585
R2515 GND.n3837 GND.n2663 585
R2516 GND.n3825 GND.n3824 585
R2517 GND.n3824 GND.n1526 585
R2518 GND.n3826 GND.n2668 585
R2519 GND.n2668 GND.n1524 585
R2520 GND.n3828 GND.n3827 585
R2521 GND.n3830 GND.n3828 585
R2522 GND.n3814 GND.n2667 585
R2523 GND.n3799 GND.n2667 585
R2524 GND.n3813 GND.n1514 585
R2525 GND.n4842 GND.n1514 585
R2526 GND.n3812 GND.n3811 585
R2527 GND.n3811 GND.n3810 585
R2528 GND.n2669 GND.n1506 585
R2529 GND.n4848 GND.n1506 585
R2530 GND.n3763 GND.n3762 585
R2531 GND.n3762 GND.n1504 585
R2532 GND.n3764 GND.n2675 585
R2533 GND.n3791 GND.n2675 585
R2534 GND.n3766 GND.n3765 585
R2535 GND.n3765 GND.n1496 585
R2536 GND.n3767 GND.n1494 585
R2537 GND.n4856 GND.n1494 585
R2538 GND.n3769 GND.n3768 585
R2539 GND.n3770 GND.n3769 585
R2540 GND.n3761 GND.n1487 585
R2541 GND.n4862 GND.n1487 585
R2542 GND.n3760 GND.n3759 585
R2543 GND.n3759 GND.n1485 585
R2544 GND.n3758 GND.n2683 585
R2545 GND.n3758 GND.n3757 585
R2546 GND.n3722 GND.n2684 585
R2547 GND.n2684 GND.n1477 585
R2548 GND.n3723 GND.n1475 585
R2549 GND.n4870 GND.n1475 585
R2550 GND.n3725 GND.n3724 585
R2551 GND.n3726 GND.n3725 585
R2552 GND.n3721 GND.n1467 585
R2553 GND.n4876 GND.n1467 585
R2554 GND.n3720 GND.n3719 585
R2555 GND.n3719 GND.n1465 585
R2556 GND.n3718 GND.n2701 585
R2557 GND.n3718 GND.n2696 585
R2558 GND.n3717 GND.n3716 585
R2559 GND.n3717 GND.n1457 585
R2560 GND.n3715 GND.n1455 585
R2561 GND.n4884 GND.n1455 585
R2562 GND.n3714 GND.n3713 585
R2563 GND.n3713 GND.n3712 585
R2564 GND.n2702 GND.n1447 585
R2565 GND.n4890 GND.n1447 585
R2566 GND.n3670 GND.n2707 585
R2567 GND.n2707 GND.n1445 585
R2568 GND.n3672 GND.n3671 585
R2569 GND.n3675 GND.n3672 585
R2570 GND.n3669 GND.n2706 585
R2571 GND.n2706 GND.n1437 585
R2572 GND.n3668 GND.n1435 585
R2573 GND.n4898 GND.n1435 585
R2574 GND.n3667 GND.n3666 585
R2575 GND.n3666 GND.n3665 585
R2576 GND.n2708 GND.n1427 585
R2577 GND.n4904 GND.n1427 585
R2578 GND.n3654 GND.n3653 585
R2579 GND.n3655 GND.n3654 585
R2580 GND.n3652 GND.n2714 585
R2581 GND.n2714 GND.n2713 585
R2582 GND.n3651 GND.n3650 585
R2583 GND.n3650 GND.n1414 585
R2584 GND.n3649 GND.n2715 585
R2585 GND.n3649 GND.n1412 585
R2586 GND.n6346 GND.n6345 585
R2587 GND.n6347 GND.n6346 585
R2588 GND.n216 GND.n215 585
R2589 GND.n6348 GND.n216 585
R2590 GND.n6351 GND.n6350 585
R2591 GND.n6350 GND.n6349 585
R2592 GND.n6352 GND.n210 585
R2593 GND.n210 GND.n209 585
R2594 GND.n6354 GND.n6353 585
R2595 GND.n6355 GND.n6354 585
R2596 GND.n208 GND.n207 585
R2597 GND.n6356 GND.n208 585
R2598 GND.n6359 GND.n6358 585
R2599 GND.n6358 GND.n6357 585
R2600 GND.n6360 GND.n202 585
R2601 GND.n202 GND.n201 585
R2602 GND.n6362 GND.n6361 585
R2603 GND.n6363 GND.n6362 585
R2604 GND.n200 GND.n199 585
R2605 GND.n6364 GND.n200 585
R2606 GND.n6367 GND.n6366 585
R2607 GND.n6366 GND.n6365 585
R2608 GND.n6368 GND.n194 585
R2609 GND.n194 GND.n193 585
R2610 GND.n6370 GND.n6369 585
R2611 GND.n6371 GND.n6370 585
R2612 GND.n192 GND.n191 585
R2613 GND.n6372 GND.n192 585
R2614 GND.n6375 GND.n6374 585
R2615 GND.n6374 GND.n6373 585
R2616 GND.n6376 GND.n186 585
R2617 GND.n186 GND.n185 585
R2618 GND.n6378 GND.n6377 585
R2619 GND.n6379 GND.n6378 585
R2620 GND.n184 GND.n183 585
R2621 GND.n6380 GND.n184 585
R2622 GND.n6383 GND.n6382 585
R2623 GND.n6382 GND.n6381 585
R2624 GND.n6384 GND.n178 585
R2625 GND.n178 GND.n177 585
R2626 GND.n6386 GND.n6385 585
R2627 GND.n6387 GND.n6386 585
R2628 GND.n176 GND.n175 585
R2629 GND.n6388 GND.n176 585
R2630 GND.n6391 GND.n6390 585
R2631 GND.n6390 GND.n6389 585
R2632 GND.n6392 GND.n170 585
R2633 GND.n170 GND.n169 585
R2634 GND.n6394 GND.n6393 585
R2635 GND.n6395 GND.n6394 585
R2636 GND.n168 GND.n167 585
R2637 GND.n6396 GND.n168 585
R2638 GND.n6399 GND.n6398 585
R2639 GND.n6398 GND.n6397 585
R2640 GND.n6400 GND.n162 585
R2641 GND.n162 GND.n161 585
R2642 GND.n6402 GND.n6401 585
R2643 GND.n6403 GND.n6402 585
R2644 GND.n160 GND.n159 585
R2645 GND.n6404 GND.n160 585
R2646 GND.n6407 GND.n6406 585
R2647 GND.n6406 GND.n6405 585
R2648 GND.n6408 GND.n154 585
R2649 GND.n154 GND.n153 585
R2650 GND.n6410 GND.n6409 585
R2651 GND.n6411 GND.n6410 585
R2652 GND.n152 GND.n151 585
R2653 GND.n6412 GND.n152 585
R2654 GND.n6415 GND.n6414 585
R2655 GND.n6414 GND.n6413 585
R2656 GND.n6416 GND.n146 585
R2657 GND.n146 GND.n144 585
R2658 GND.n6418 GND.n6417 585
R2659 GND.n6419 GND.n6418 585
R2660 GND.n147 GND.n145 585
R2661 GND.n145 GND.n135 585
R2662 GND.n4528 GND.n4527 585
R2663 GND.n4527 GND.n81 585
R2664 GND.n4529 GND.n4521 585
R2665 GND.n4521 GND.n79 585
R2666 GND.n4531 GND.n4530 585
R2667 GND.n4531 GND.n2053 585
R2668 GND.n4532 GND.n4520 585
R2669 GND.n4532 GND.n2055 585
R2670 GND.n4534 GND.n4533 585
R2671 GND.n4533 GND.n2064 585
R2672 GND.n4535 GND.n2070 585
R2673 GND.n2070 GND.n2062 585
R2674 GND.n4537 GND.n4536 585
R2675 GND.n4538 GND.n4537 585
R2676 GND.n2071 GND.n2069 585
R2677 GND.n2076 GND.n2069 585
R2678 GND.n4514 GND.n4513 585
R2679 GND.n4513 GND.n4512 585
R2680 GND.n2074 GND.n2073 585
R2681 GND.n2085 GND.n2074 585
R2682 GND.n4490 GND.n2089 585
R2683 GND.n2089 GND.n2084 585
R2684 GND.n4492 GND.n4491 585
R2685 GND.n4493 GND.n4492 585
R2686 GND.n2090 GND.n2088 585
R2687 GND.n2095 GND.n2088 585
R2688 GND.n4485 GND.n4484 585
R2689 GND.n4484 GND.n4483 585
R2690 GND.n2093 GND.n2092 585
R2691 GND.n2107 GND.n2093 585
R2692 GND.n4464 GND.n2112 585
R2693 GND.n2112 GND.n2104 585
R2694 GND.n4466 GND.n4465 585
R2695 GND.n4467 GND.n4466 585
R2696 GND.n2113 GND.n2111 585
R2697 GND.n2120 GND.n2111 585
R2698 GND.n4459 GND.n4458 585
R2699 GND.n4458 GND.n4457 585
R2700 GND.n2116 GND.n2115 585
R2701 GND.n2129 GND.n2116 585
R2702 GND.n4438 GND.n2134 585
R2703 GND.n2134 GND.n2128 585
R2704 GND.n4440 GND.n4439 585
R2705 GND.n4441 GND.n4440 585
R2706 GND.n2135 GND.n2133 585
R2707 GND.n4387 GND.n2133 585
R2708 GND.n4400 GND.n4399 585
R2709 GND.n4401 GND.n4400 585
R2710 GND.n4398 GND.n4397 585
R2711 GND.n4397 GND.n4381 585
R2712 GND.n4396 GND.n4395 585
R2713 GND.n4396 GND.n4380 585
R2714 GND.n4394 GND.n2169 585
R2715 GND.n4372 GND.n2169 585
R2716 GND.n4416 GND.n4415 585
R2717 GND.n4415 GND.n4414 585
R2718 GND.n4418 GND.n4417 585
R2719 GND.n4419 GND.n4418 585
R2720 GND.n2168 GND.n2167 585
R2721 GND.n2168 GND.n2159 585
R2722 GND.n2166 GND.n2165 585
R2723 GND.n2165 GND.n2157 585
R2724 GND.n2146 GND.n2144 585
R2725 GND.n2149 GND.n2146 585
R2726 GND.n4433 GND.n4432 585
R2727 GND.n4432 GND.n4431 585
R2728 GND.n2145 GND.n2143 585
R2729 GND.n2179 GND.n2145 585
R2730 GND.n4257 GND.n4256 585
R2731 GND.n4256 GND.n2178 585
R2732 GND.n4258 GND.n4251 585
R2733 GND.n4251 GND.n2190 585
R2734 GND.n4260 GND.n4259 585
R2735 GND.n4260 GND.n2188 585
R2736 GND.n4261 GND.n4250 585
R2737 GND.n4261 GND.n2193 585
R2738 GND.n4263 GND.n4262 585
R2739 GND.n4262 GND.n2202 585
R2740 GND.n4264 GND.n4245 585
R2741 GND.n4245 GND.n2200 585
R2742 GND.n4266 GND.n4265 585
R2743 GND.n4266 GND.n2213 585
R2744 GND.n4267 GND.n4244 585
R2745 GND.n4267 GND.n2211 585
R2746 GND.n4269 GND.n4268 585
R2747 GND.n4268 GND.n2215 585
R2748 GND.n4270 GND.n4239 585
R2749 GND.n4239 GND.n2223 585
R2750 GND.n4272 GND.n4271 585
R2751 GND.n4272 GND.n2222 585
R2752 GND.n4273 GND.n4238 585
R2753 GND.n4273 GND.n2235 585
R2754 GND.n4275 GND.n4274 585
R2755 GND.n4274 GND.n2233 585
R2756 GND.n4276 GND.n4228 585
R2757 GND.n4228 GND.n2237 585
R2758 GND.n4278 GND.n4277 585
R2759 GND.n4279 GND.n4278 585
R2760 GND.n4229 GND.n4227 585
R2761 GND.n4227 GND.n1895 585
R2762 GND.n4232 GND.n4231 585
R2763 GND.n4231 GND.n1892 585
R2764 GND.n1879 GND.n1878 585
R2765 GND.n1883 GND.n1879 585
R2766 GND.n4642 GND.n4641 585
R2767 GND.n4641 GND.n4640 585
R2768 GND.n4643 GND.n1873 585
R2769 GND.n1880 GND.n1873 585
R2770 GND.n4645 GND.n4644 585
R2771 GND.n4646 GND.n4645 585
R2772 GND.n1870 GND.n1869 585
R2773 GND.n4647 GND.n1870 585
R2774 GND.n4650 GND.n4649 585
R2775 GND.n4649 GND.n4648 585
R2776 GND.n4651 GND.n1862 585
R2777 GND.n1862 GND.n1860 585
R2778 GND.n4653 GND.n4652 585
R2779 GND.n4654 GND.n4653 585
R2780 GND.n1863 GND.n1861 585
R2781 GND.n1861 GND.n1858 585
R2782 GND.n1844 GND.n1843 585
R2783 GND.n1848 GND.n1844 585
R2784 GND.n4664 GND.n4663 585
R2785 GND.n4663 GND.n4662 585
R2786 GND.n4665 GND.n1836 585
R2787 GND.n1845 GND.n1836 585
R2788 GND.n4667 GND.n4666 585
R2789 GND.n4668 GND.n4667 585
R2790 GND.n1837 GND.n1835 585
R2791 GND.n1835 GND.n1832 585
R2792 GND.n1817 GND.n1816 585
R2793 GND.n1821 GND.n1817 585
R2794 GND.n4678 GND.n4677 585
R2795 GND.n4677 GND.n4676 585
R2796 GND.n4679 GND.n1809 585
R2797 GND.n1818 GND.n1809 585
R2798 GND.n4681 GND.n4680 585
R2799 GND.n4682 GND.n4681 585
R2800 GND.n1810 GND.n1808 585
R2801 GND.n1808 GND.n1805 585
R2802 GND.n1791 GND.n1790 585
R2803 GND.n2288 GND.n1791 585
R2804 GND.n4692 GND.n4691 585
R2805 GND.n4691 GND.n4690 585
R2806 GND.n4693 GND.n1783 585
R2807 GND.n1792 GND.n1783 585
R2808 GND.n4695 GND.n4694 585
R2809 GND.n4696 GND.n4695 585
R2810 GND.n1784 GND.n1782 585
R2811 GND.n1782 GND.n1779 585
R2812 GND.n1765 GND.n1764 585
R2813 GND.n1768 GND.n1765 585
R2814 GND.n4706 GND.n4705 585
R2815 GND.n4705 GND.n4704 585
R2816 GND.n4707 GND.n1759 585
R2817 GND.n2296 GND.n1759 585
R2818 GND.n4709 GND.n4708 585
R2819 GND.n4710 GND.n4709 585
R2820 GND.n1760 GND.n1758 585
R2821 GND.n4142 GND.n1758 585
R2822 GND.n2315 GND.n2314 585
R2823 GND.n2316 GND.n2315 585
R2824 GND.n2303 GND.n2302 585
R2825 GND.n2302 GND.n1745 585
R2826 GND.n2309 GND.n2308 585
R2827 GND.n2308 GND.n1739 585
R2828 GND.n2307 GND.n2306 585
R2829 GND.n2307 GND.n1736 585
R2830 GND.n1724 GND.n1723 585
R2831 GND.n2612 GND.n1724 585
R2832 GND.n4734 GND.n4733 585
R2833 GND.n4733 GND.n4732 585
R2834 GND.n4735 GND.n1710 585
R2835 GND.n2618 GND.n1710 585
R2836 GND.n4737 GND.n4736 585
R2837 GND.n4738 GND.n4737 585
R2838 GND.n1711 GND.n1709 585
R2839 GND.n1709 GND.n1701 585
R2840 GND.n1717 GND.n1716 585
R2841 GND.n1716 GND.n1698 585
R2842 GND.n1715 GND.n1714 585
R2843 GND.n1715 GND.n1684 585
R2844 GND.n1672 GND.n1671 585
R2845 GND.n1681 GND.n1672 585
R2846 GND.n4761 GND.n4760 585
R2847 GND.n4760 GND.n4759 585
R2848 GND.n4762 GND.n1661 585
R2849 GND.n2635 GND.n1661 585
R2850 GND.n4764 GND.n4763 585
R2851 GND.n4765 GND.n4764 585
R2852 GND.n1662 GND.n1660 585
R2853 GND.n3954 GND.n1660 585
R2854 GND.n1665 GND.n1664 585
R2855 GND.n1664 GND.n1640 585
R2856 GND.n1628 GND.n1627 585
R2857 GND.n1637 GND.n1628 585
R2858 GND.n4782 GND.n4781 585
R2859 GND.n4781 GND.n4780 585
R2860 GND.n4783 GND.n1617 585
R2861 GND.n3917 GND.n1617 585
R2862 GND.n4785 GND.n4784 585
R2863 GND.n4786 GND.n4785 585
R2864 GND.n1618 GND.n1616 585
R2865 GND.n1616 GND.n1607 585
R2866 GND.n1621 GND.n1620 585
R2867 GND.n1620 GND.n1604 585
R2868 GND.n1587 GND.n1586 585
R2869 GND.n2644 GND.n1587 585
R2870 GND.n4803 GND.n4802 585
R2871 GND.n4802 GND.n4801 585
R2872 GND.n4804 GND.n1573 585
R2873 GND.n2651 GND.n1573 585
R2874 GND.n4806 GND.n4805 585
R2875 GND.n4807 GND.n4806 585
R2876 GND.n1574 GND.n1572 585
R2877 GND.n1572 GND.n1563 585
R2878 GND.n1580 GND.n1579 585
R2879 GND.n1579 GND.n1560 585
R2880 GND.n1578 GND.n1577 585
R2881 GND.n1578 GND.n1546 585
R2882 GND.n1534 GND.n1533 585
R2883 GND.n1543 GND.n1534 585
R2884 GND.n4830 GND.n4829 585
R2885 GND.n4829 GND.n4828 585
R2886 GND.n4831 GND.n1528 585
R2887 GND.n2664 GND.n1528 585
R2888 GND.n4833 GND.n4832 585
R2889 GND.n4834 GND.n4833 585
R2890 GND.n1529 GND.n1527 585
R2891 GND.n3829 GND.n1527 585
R2892 GND.n3782 GND.n3781 585
R2893 GND.n3782 GND.n1516 585
R2894 GND.n3784 GND.n3783 585
R2895 GND.n3783 GND.n1513 585
R2896 GND.n3785 GND.n2677 585
R2897 GND.n2677 GND.n1507 585
R2898 GND.n3787 GND.n3786 585
R2899 GND.n3788 GND.n3787 585
R2900 GND.n2678 GND.n2676 585
R2901 GND.n2676 GND.n2674 585
R2902 GND.n3773 GND.n3772 585
R2903 GND.n3772 GND.n3771 585
R2904 GND.n2681 GND.n2680 585
R2905 GND.n2681 GND.n1488 585
R2906 GND.n3753 GND.n3752 585
R2907 GND.n3754 GND.n3753 585
R2908 GND.n2688 GND.n2687 585
R2909 GND.n2687 GND.n2686 585
R2910 GND.n3748 GND.n3747 585
R2911 GND.n3747 GND.n1474 585
R2912 GND.n3746 GND.n2690 585
R2913 GND.n3746 GND.n1468 585
R2914 GND.n3745 GND.n2692 585
R2915 GND.n3745 GND.n3744 585
R2916 GND.n3696 GND.n2691 585
R2917 GND.n2693 GND.n2691 585
R2918 GND.n3698 GND.n3697 585
R2919 GND.n3697 GND.n1454 585
R2920 GND.n3699 GND.n3678 585
R2921 GND.n3678 GND.n1448 585
R2922 GND.n3701 GND.n3700 585
R2923 GND.n3702 GND.n3701 585
R2924 GND.n3679 GND.n3677 585
R2925 GND.n3677 GND.n3676 585
R2926 GND.n3688 GND.n3687 585
R2927 GND.n3687 GND.n1434 585
R2928 GND.n3686 GND.n3681 585
R2929 GND.n3686 GND.n1428 585
R2930 GND.n3685 GND.n3684 585
R2931 GND.n3685 GND.n1425 585
R2932 GND.n1411 GND.n1410 585
R2933 GND.n2712 GND.n1411 585
R2934 GND.n4914 GND.n4913 585
R2935 GND.n4913 GND.n4912 585
R2936 GND.n4915 GND.n1403 585
R2937 GND.n3562 GND.n1403 585
R2938 GND.n4917 GND.n4916 585
R2939 GND.n4918 GND.n4917 585
R2940 GND.n1404 GND.n1402 585
R2941 GND.n1402 GND.n1399 585
R2942 GND.n1384 GND.n1383 585
R2943 GND.n1388 GND.n1384 585
R2944 GND.n4928 GND.n4927 585
R2945 GND.n4927 GND.n4926 585
R2946 GND.n4929 GND.n1376 585
R2947 GND.n1385 GND.n1376 585
R2948 GND.n4931 GND.n4930 585
R2949 GND.n4932 GND.n4931 585
R2950 GND.n1377 GND.n1375 585
R2951 GND.n1375 GND.n1372 585
R2952 GND.n1357 GND.n1356 585
R2953 GND.n1361 GND.n1357 585
R2954 GND.n4942 GND.n4941 585
R2955 GND.n4941 GND.n4940 585
R2956 GND.n4943 GND.n1349 585
R2957 GND.n1358 GND.n1349 585
R2958 GND.n4945 GND.n4944 585
R2959 GND.n4946 GND.n4945 585
R2960 GND.n1350 GND.n1348 585
R2961 GND.n1348 GND.n1345 585
R2962 GND.n1330 GND.n1329 585
R2963 GND.n1334 GND.n1330 585
R2964 GND.n4956 GND.n4955 585
R2965 GND.n4955 GND.n4954 585
R2966 GND.n4957 GND.n1316 585
R2967 GND.n1331 GND.n1316 585
R2968 GND.n4959 GND.n4958 585
R2969 GND.n4960 GND.n4959 585
R2970 GND.n1317 GND.n1315 585
R2971 GND.n1315 GND.n1312 585
R2972 GND.n1323 GND.n1322 585
R2973 GND.n1322 GND.n1303 585
R2974 GND.n1321 GND.n1299 585
R2975 GND.n4968 GND.n1299 585
R2976 GND.n4971 GND.n1300 585
R2977 GND.n4971 GND.n4970 585
R2978 GND.n4972 GND.n1298 585
R2979 GND.n4972 GND.n1247 585
R2980 GND.n4974 GND.n4973 585
R2981 GND.n4973 GND.n1233 585
R2982 GND.n4975 GND.n1293 585
R2983 GND.n1293 GND.n1291 585
R2984 GND.n4977 GND.n4976 585
R2985 GND.n4978 GND.n4977 585
R2986 GND.n1294 GND.n1292 585
R2987 GND.n1292 GND.n1276 585
R2988 GND.n3337 GND.n3336 585
R2989 GND.n3336 GND.n1168 585
R2990 GND.n3338 GND.n3330 585
R2991 GND.n3330 GND.n1166 585
R2992 GND.n3340 GND.n3339 585
R2993 GND.n3340 GND.n2845 585
R2994 GND.n3341 GND.n3329 585
R2995 GND.n3341 GND.n2847 585
R2996 GND.n3343 GND.n3342 585
R2997 GND.n3342 GND.n2855 585
R2998 GND.n3344 GND.n3324 585
R2999 GND.n3324 GND.n2853 585
R3000 GND.n3346 GND.n3345 585
R3001 GND.n3346 GND.n2858 585
R3002 GND.n3347 GND.n3323 585
R3003 GND.n3347 GND.n2867 585
R3004 GND.n3349 GND.n3348 585
R3005 GND.n3348 GND.n2865 585
R3006 GND.n3350 GND.n3318 585
R3007 GND.n3318 GND.n2878 585
R3008 GND.n3352 GND.n3351 585
R3009 GND.n3352 GND.n2876 585
R3010 GND.n3353 GND.n3317 585
R3011 GND.n3353 GND.n2880 585
R3012 GND.n3358 GND.n3357 585
R3013 GND.n3357 GND.n3356 585
R3014 GND.n3359 GND.n3312 585
R3015 GND.n3312 GND.n2887 585
R3016 GND.n3361 GND.n3360 585
R3017 GND.n3361 GND.n2897 585
R3018 GND.n3362 GND.n3311 585
R3019 GND.n3362 GND.n2895 585
R3020 GND.n3364 GND.n3363 585
R3021 GND.n3363 GND.n2899 585
R3022 GND.n3365 GND.n2923 585
R3023 GND.n2923 GND.n2907 585
R3024 GND.n3367 GND.n3366 585
R3025 GND.n3368 GND.n3367 585
R3026 GND.n2924 GND.n2922 585
R3027 GND.n2922 GND.n2920 585
R3028 GND.n3305 GND.n3304 585
R3029 GND.n3304 GND.n2917 585
R3030 GND.n3303 GND.n2926 585
R3031 GND.n3303 GND.n3302 585
R3032 GND.n3257 GND.n2927 585
R3033 GND.n2936 GND.n2927 585
R3034 GND.n3258 GND.n3253 585
R3035 GND.n3253 GND.n2935 585
R3036 GND.n3261 GND.n3260 585
R3037 GND.n3262 GND.n3261 585
R3038 GND.n3255 GND.n3252 585
R3039 GND.n3252 GND.n2975 585
R3040 GND.n2962 GND.n2961 585
R3041 GND.n2966 GND.n2962 585
R3042 GND.n3275 GND.n3274 585
R3043 GND.n3274 GND.n3273 585
R3044 GND.n3277 GND.n2959 585
R3045 GND.n3237 GND.n2959 585
R3046 GND.n3279 GND.n3278 585
R3047 GND.n3280 GND.n3279 585
R3048 GND.n3223 GND.n2958 585
R3049 GND.n2958 GND.n2953 585
R3050 GND.n3224 GND.n2985 585
R3051 GND.n2985 GND.n2951 585
R3052 GND.n3226 GND.n3225 585
R3053 GND.n3227 GND.n3226 585
R3054 GND.n2986 GND.n2984 585
R3055 GND.n2991 GND.n2984 585
R3056 GND.n3218 GND.n3217 585
R3057 GND.n3217 GND.n3216 585
R3058 GND.n2989 GND.n2988 585
R3059 GND.n3004 GND.n2989 585
R3060 GND.n3188 GND.n3013 585
R3061 GND.n3013 GND.n3001 585
R3062 GND.n3190 GND.n3189 585
R3063 GND.n3191 GND.n3190 585
R3064 GND.n3014 GND.n3012 585
R3065 GND.n3021 GND.n3012 585
R3066 GND.n3183 GND.n3182 585
R3067 GND.n3182 GND.n3181 585
R3068 GND.n3017 GND.n3016 585
R3069 GND.n3033 GND.n3017 585
R3070 GND.n3131 GND.n3130 585
R3071 GND.n3131 GND.n3031 585
R3072 GND.n3132 GND.n3127 585
R3073 GND.n3132 GND.n3036 585
R3074 GND.n3134 GND.n3133 585
R3075 GND.n3133 GND.n3045 585
R3076 GND.n3135 GND.n3117 585
R3077 GND.n3117 GND.n3043 585
R3078 GND.n3137 GND.n3136 585
R3079 GND.n3138 GND.n3137 585
R3080 GND.n3118 GND.n3116 585
R3081 GND.n3116 GND.n1054 585
R3082 GND.n3121 GND.n3120 585
R3083 GND.n3120 GND.n1051 585
R3084 GND.n1031 GND.n1030 585
R3085 GND.n3105 GND.n1031 585
R3086 GND.n5183 GND.n5182 585
R3087 GND.n5182 GND.n5181 585
R3088 GND.n5184 GND.n1020 585
R3089 GND.n1032 GND.n1020 585
R3090 GND.n5186 GND.n5185 585
R3091 GND.n5187 GND.n5186 585
R3092 GND.n1021 GND.n1019 585
R3093 GND.n1019 GND.n1014 585
R3094 GND.n1024 GND.n1023 585
R3095 GND.n1023 GND.n967 585
R3096 GND.n941 GND.n940 585
R3097 GND.n5265 GND.n941 585
R3098 GND.n5268 GND.n5267 585
R3099 GND.n5267 GND.n5266 585
R3100 GND.n5269 GND.n935 585
R3101 GND.n935 GND.n934 585
R3102 GND.n5271 GND.n5270 585
R3103 GND.n5272 GND.n5271 585
R3104 GND.n933 GND.n932 585
R3105 GND.n5273 GND.n933 585
R3106 GND.n5276 GND.n5275 585
R3107 GND.n5275 GND.n5274 585
R3108 GND.n5277 GND.n927 585
R3109 GND.n927 GND.n926 585
R3110 GND.n5279 GND.n5278 585
R3111 GND.n5280 GND.n5279 585
R3112 GND.n925 GND.n924 585
R3113 GND.n5281 GND.n925 585
R3114 GND.n5284 GND.n5283 585
R3115 GND.n5283 GND.n5282 585
R3116 GND.n5285 GND.n919 585
R3117 GND.n919 GND.n918 585
R3118 GND.n5287 GND.n5286 585
R3119 GND.n5288 GND.n5287 585
R3120 GND.n917 GND.n916 585
R3121 GND.n5289 GND.n917 585
R3122 GND.n5292 GND.n5291 585
R3123 GND.n5291 GND.n5290 585
R3124 GND.n5293 GND.n911 585
R3125 GND.n911 GND.n910 585
R3126 GND.n5295 GND.n5294 585
R3127 GND.n5296 GND.n5295 585
R3128 GND.n909 GND.n908 585
R3129 GND.n5297 GND.n909 585
R3130 GND.n5300 GND.n5299 585
R3131 GND.n5299 GND.n5298 585
R3132 GND.n5301 GND.n903 585
R3133 GND.n903 GND.n902 585
R3134 GND.n5303 GND.n5302 585
R3135 GND.n5304 GND.n5303 585
R3136 GND.n901 GND.n900 585
R3137 GND.n5305 GND.n901 585
R3138 GND.n5308 GND.n5307 585
R3139 GND.n5307 GND.n5306 585
R3140 GND.n5309 GND.n895 585
R3141 GND.n895 GND.n894 585
R3142 GND.n5311 GND.n5310 585
R3143 GND.n5312 GND.n5311 585
R3144 GND.n893 GND.n892 585
R3145 GND.n5313 GND.n893 585
R3146 GND.n5316 GND.n5315 585
R3147 GND.n5315 GND.n5314 585
R3148 GND.n5317 GND.n887 585
R3149 GND.n887 GND.n886 585
R3150 GND.n5319 GND.n5318 585
R3151 GND.n5320 GND.n5319 585
R3152 GND.n885 GND.n884 585
R3153 GND.n5321 GND.n885 585
R3154 GND.n5324 GND.n5323 585
R3155 GND.n5323 GND.n5322 585
R3156 GND.n5325 GND.n879 585
R3157 GND.n879 GND.n878 585
R3158 GND.n5327 GND.n5326 585
R3159 GND.n5328 GND.n5327 585
R3160 GND.n877 GND.n876 585
R3161 GND.n5329 GND.n877 585
R3162 GND.n5332 GND.n5331 585
R3163 GND.n5331 GND.n5330 585
R3164 GND.n5333 GND.n870 585
R3165 GND.n870 GND.n869 585
R3166 GND.n5335 GND.n5334 585
R3167 GND.n5336 GND.n5335 585
R3168 GND.n871 GND.n868 585
R3169 GND.n5337 GND.n868 585
R3170 GND.n2538 GND.n2537 585
R3171 GND.n2537 GND.n1872 585
R3172 GND.n2536 GND.n2440 585
R3173 GND.n2534 GND.n2533 585
R3174 GND.n2442 GND.n2441 585
R3175 GND.n2529 GND.n2445 585
R3176 GND.n2528 GND.n2446 585
R3177 GND.n2454 GND.n2447 585
R3178 GND.n2455 GND.n2452 585
R3179 GND.n2520 GND.n2457 585
R3180 GND.n2519 GND.n2458 585
R3181 GND.n2469 GND.n2459 585
R3182 GND.n2512 GND.n2470 585
R3183 GND.n2511 GND.n2472 585
R3184 GND.n2481 GND.n2473 585
R3185 GND.n2504 GND.n2483 585
R3186 GND.n2503 GND.n2500 585
R3187 GND.n2498 GND.n2484 585
R3188 GND.n1997 GND.n82 585
R3189 GND.n6502 GND.n82 585
R3190 GND.n4553 GND.n1996 585
R3191 GND.n4554 GND.n4553 585
R3192 GND.n4552 GND.n1995 585
R3193 GND.n4552 GND.n4551 585
R3194 GND.n2054 GND.n1994 585
R3195 GND.n2063 GND.n2054 585
R3196 GND.n4542 GND.n4541 585
R3197 GND.n4543 GND.n4542 585
R3198 GND.n4540 GND.n1988 585
R3199 GND.n4540 GND.n4539 585
R3200 GND.n2065 GND.n1987 585
R3201 GND.n2068 GND.n2065 585
R3202 GND.n2077 GND.n1986 585
R3203 GND.n4511 GND.n2077 585
R3204 GND.n4499 GND.n4498 585
R3205 GND.n4499 GND.n2075 585
R3206 GND.n4500 GND.n1980 585
R3207 GND.n4501 GND.n4500 585
R3208 GND.n4497 GND.n1979 585
R3209 GND.n4497 GND.n4496 585
R3210 GND.n2086 GND.n1978 585
R3211 GND.n2087 GND.n2086 585
R3212 GND.n2097 GND.n2096 585
R3213 GND.n4482 GND.n2097 585
R3214 GND.n4470 GND.n1972 585
R3215 GND.n4470 GND.n2094 585
R3216 GND.n4471 GND.n1971 585
R3217 GND.n4472 GND.n4471 585
R3218 GND.n4469 GND.n1970 585
R3219 GND.n4469 GND.n4468 585
R3220 GND.n2109 GND.n2108 585
R3221 GND.n2110 GND.n2109 585
R3222 GND.n2121 GND.n1964 585
R3223 GND.n4456 GND.n2121 585
R3224 GND.n4444 GND.n1963 585
R3225 GND.n4444 GND.n2119 585
R3226 GND.n4445 GND.n1962 585
R3227 GND.n4446 GND.n4445 585
R3228 GND.n4443 GND.n2131 585
R3229 GND.n4443 GND.n4442 585
R3230 GND.n2130 GND.n1956 585
R3231 GND.n2132 GND.n2130 585
R3232 GND.n4384 GND.n1955 585
R3233 GND.n4393 GND.n4384 585
R3234 GND.n4403 GND.n1954 585
R3235 GND.n4403 GND.n4402 585
R3236 GND.n4405 GND.n4404 585
R3237 GND.n4406 GND.n4405 585
R3238 GND.n4383 GND.n1948 585
R3239 GND.n4383 GND.n4382 585
R3240 GND.n4373 GND.n1947 585
R3241 GND.n4413 GND.n4373 585
R3242 GND.n2161 GND.n1946 585
R3243 GND.n2164 GND.n2161 585
R3244 GND.n4421 GND.n2162 585
R3245 GND.n4421 GND.n4420 585
R3246 GND.n4422 GND.n1940 585
R3247 GND.n4423 GND.n4422 585
R3248 GND.n2160 GND.n1939 585
R3249 GND.n4362 GND.n2160 585
R3250 GND.n2150 GND.n1938 585
R3251 GND.n4430 GND.n2150 585
R3252 GND.n2181 GND.n2180 585
R3253 GND.n2181 GND.n2147 585
R3254 GND.n2182 GND.n1932 585
R3255 GND.n4354 GND.n2182 585
R3256 GND.n4343 GND.n1931 585
R3257 GND.n4343 GND.n4342 585
R3258 GND.n4344 GND.n1930 585
R3259 GND.n4345 GND.n4344 585
R3260 GND.n4340 GND.n2192 585
R3261 GND.n4340 GND.n4339 585
R3262 GND.n2191 GND.n1924 585
R3263 GND.n2205 GND.n2191 585
R3264 GND.n2203 GND.n1923 585
R3265 GND.n4330 GND.n2203 585
R3266 GND.n4317 GND.n1922 585
R3267 GND.n4317 GND.n4316 585
R3268 GND.n4319 GND.n4318 585
R3269 GND.n4320 GND.n4319 585
R3270 GND.n4315 GND.n1916 585
R3271 GND.n4315 GND.n4314 585
R3272 GND.n2214 GND.n1915 585
R3273 GND.n2227 GND.n2214 585
R3274 GND.n2224 GND.n1914 585
R3275 GND.n4305 GND.n2224 585
R3276 GND.n4293 GND.n4291 585
R3277 GND.n4293 GND.n4292 585
R3278 GND.n4294 GND.n1908 585
R3279 GND.n4295 GND.n4294 585
R3280 GND.n4290 GND.n1907 585
R3281 GND.n4290 GND.n4289 585
R3282 GND.n2236 GND.n1906 585
R3283 GND.n4226 GND.n2236 585
R3284 GND.n1899 GND.n1897 585
R3285 GND.n4280 GND.n1897 585
R3286 GND.n4632 GND.n4631 585
R3287 GND.n4633 GND.n4632 585
R3288 GND.n1898 GND.n1896 585
R3289 GND.n2245 GND.n1896 585
R3290 GND.n2436 GND.n1884 585
R3291 GND.n4639 GND.n1884 585
R3292 GND.n2024 GND.n78 585
R3293 GND.n6444 GND.n78 585
R3294 GND.n2023 GND.n2022 585
R3295 GND.n2028 GND.n2019 585
R3296 GND.n2029 GND.n2018 585
R3297 GND.n2030 GND.n2017 585
R3298 GND.n2016 GND.n2014 585
R3299 GND.n2034 GND.n2013 585
R3300 GND.n2035 GND.n2012 585
R3301 GND.n2036 GND.n2011 585
R3302 GND.n2010 GND.n2008 585
R3303 GND.n2040 GND.n2007 585
R3304 GND.n2041 GND.n2006 585
R3305 GND.n2042 GND.n2005 585
R3306 GND.n2004 GND.n2002 585
R3307 GND.n2046 GND.n2001 585
R3308 GND.n2047 GND.n2000 585
R3309 GND.n2048 GND.n1999 585
R3310 GND.n6504 GND.n6503 585
R3311 GND.n6503 GND.n6502 585
R3312 GND.n6505 GND.n77 585
R3313 GND.n4554 GND.n77 585
R3314 GND.n2056 GND.n75 585
R3315 GND.n4551 GND.n2056 585
R3316 GND.n6509 GND.n74 585
R3317 GND.n2063 GND.n74 585
R3318 GND.n6510 GND.n73 585
R3319 GND.n4543 GND.n73 585
R3320 GND.n6511 GND.n72 585
R3321 GND.n4539 GND.n72 585
R3322 GND.n2067 GND.n70 585
R3323 GND.n2068 GND.n2067 585
R3324 GND.n6515 GND.n69 585
R3325 GND.n4511 GND.n69 585
R3326 GND.n6516 GND.n68 585
R3327 GND.n2075 GND.n68 585
R3328 GND.n6517 GND.n67 585
R3329 GND.n4501 GND.n67 585
R3330 GND.n4495 GND.n65 585
R3331 GND.n4496 GND.n4495 585
R3332 GND.n6521 GND.n64 585
R3333 GND.n2087 GND.n64 585
R3334 GND.n6522 GND.n63 585
R3335 GND.n4482 GND.n63 585
R3336 GND.n6523 GND.n62 585
R3337 GND.n2094 GND.n62 585
R3338 GND.n2106 GND.n60 585
R3339 GND.n4472 GND.n2106 585
R3340 GND.n6527 GND.n59 585
R3341 GND.n4468 GND.n59 585
R3342 GND.n6528 GND.n58 585
R3343 GND.n2110 GND.n58 585
R3344 GND.n6529 GND.n57 585
R3345 GND.n4456 GND.n57 585
R3346 GND.n2118 GND.n55 585
R3347 GND.n2119 GND.n2118 585
R3348 GND.n6533 GND.n54 585
R3349 GND.n4446 GND.n54 585
R3350 GND.n6534 GND.n53 585
R3351 GND.n4442 GND.n53 585
R3352 GND.n6535 GND.n52 585
R3353 GND.n2132 GND.n52 585
R3354 GND.n4386 GND.n50 585
R3355 GND.n4393 GND.n4386 585
R3356 GND.n6539 GND.n49 585
R3357 GND.n4402 GND.n49 585
R3358 GND.n6540 GND.n48 585
R3359 GND.n4406 GND.n48 585
R3360 GND.n6541 GND.n47 585
R3361 GND.n4382 GND.n47 585
R3362 GND.n4371 GND.n46 585
R3363 GND.n4413 GND.n4371 585
R3364 GND.n4370 GND.n4369 585
R3365 GND.n4370 GND.n2164 585
R3366 GND.n2171 GND.n2163 585
R3367 GND.n4420 GND.n2163 585
R3368 GND.n4365 GND.n2158 585
R3369 GND.n4423 GND.n2158 585
R3370 GND.n4364 GND.n4363 585
R3371 GND.n4363 GND.n4362 585
R3372 GND.n4360 GND.n2148 585
R3373 GND.n4430 GND.n2148 585
R3374 GND.n2177 GND.n2173 585
R3375 GND.n2177 GND.n2147 585
R3376 GND.n4356 GND.n4355 585
R3377 GND.n4355 GND.n4354 585
R3378 GND.n2176 GND.n2175 585
R3379 GND.n4342 GND.n2176 585
R3380 GND.n2196 GND.n2189 585
R3381 GND.n4345 GND.n2189 585
R3382 GND.n4338 GND.n4337 585
R3383 GND.n4339 GND.n4338 585
R3384 GND.n2195 GND.n2194 585
R3385 GND.n2205 GND.n2194 585
R3386 GND.n4332 GND.n4331 585
R3387 GND.n4331 GND.n4330 585
R3388 GND.n2199 GND.n2198 585
R3389 GND.n4316 GND.n2199 585
R3390 GND.n2218 GND.n2212 585
R3391 GND.n4320 GND.n2212 585
R3392 GND.n4313 GND.n4312 585
R3393 GND.n4314 GND.n4313 585
R3394 GND.n2217 GND.n2216 585
R3395 GND.n2227 GND.n2216 585
R3396 GND.n4307 GND.n4306 585
R3397 GND.n4306 GND.n4305 585
R3398 GND.n2221 GND.n2220 585
R3399 GND.n4292 GND.n2221 585
R3400 GND.n2241 GND.n2234 585
R3401 GND.n4295 GND.n2234 585
R3402 GND.n4288 GND.n4287 585
R3403 GND.n4289 GND.n4288 585
R3404 GND.n2240 GND.n2239 585
R3405 GND.n4226 GND.n2239 585
R3406 GND.n4282 GND.n4281 585
R3407 GND.n4281 GND.n4280 585
R3408 GND.n4221 GND.n1894 585
R3409 GND.n4633 GND.n1894 585
R3410 GND.n4220 GND.n2246 585
R3411 GND.n2246 GND.n2245 585
R3412 GND.n2243 GND.n1882 585
R3413 GND.n4639 GND.n1882 585
R3414 GND.n4140 GND.n2320 530.939
R3415 GND.n4018 GND.n2318 530.939
R3416 GND.n3649 GND.n3648 530.939
R3417 GND.n3644 GND.n3565 530.939
R3418 GND.n5458 GND.n745 358.839
R3419 GND.n6347 GND.n217 345.356
R3420 GND.n6196 GND.n307 301.784
R3421 GND.n6197 GND.n6196 301.784
R3422 GND.n6198 GND.n6197 301.784
R3423 GND.n6198 GND.n301 301.784
R3424 GND.n6206 GND.n301 301.784
R3425 GND.n6207 GND.n6206 301.784
R3426 GND.n6208 GND.n6207 301.784
R3427 GND.n6208 GND.n295 301.784
R3428 GND.n6216 GND.n295 301.784
R3429 GND.n6217 GND.n6216 301.784
R3430 GND.n6218 GND.n6217 301.784
R3431 GND.n6218 GND.n289 301.784
R3432 GND.n6226 GND.n289 301.784
R3433 GND.n6227 GND.n6226 301.784
R3434 GND.n6228 GND.n6227 301.784
R3435 GND.n6228 GND.n283 301.784
R3436 GND.n6236 GND.n283 301.784
R3437 GND.n6237 GND.n6236 301.784
R3438 GND.n6238 GND.n6237 301.784
R3439 GND.n6238 GND.n277 301.784
R3440 GND.n6246 GND.n277 301.784
R3441 GND.n6247 GND.n6246 301.784
R3442 GND.n6248 GND.n6247 301.784
R3443 GND.n6248 GND.n271 301.784
R3444 GND.n6256 GND.n271 301.784
R3445 GND.n6257 GND.n6256 301.784
R3446 GND.n6258 GND.n6257 301.784
R3447 GND.n6258 GND.n265 301.784
R3448 GND.n6266 GND.n265 301.784
R3449 GND.n6267 GND.n6266 301.784
R3450 GND.n6268 GND.n6267 301.784
R3451 GND.n6268 GND.n259 301.784
R3452 GND.n6276 GND.n259 301.784
R3453 GND.n6277 GND.n6276 301.784
R3454 GND.n6278 GND.n6277 301.784
R3455 GND.n6278 GND.n253 301.784
R3456 GND.n6286 GND.n253 301.784
R3457 GND.n6287 GND.n6286 301.784
R3458 GND.n6288 GND.n6287 301.784
R3459 GND.n6288 GND.n247 301.784
R3460 GND.n6296 GND.n247 301.784
R3461 GND.n6297 GND.n6296 301.784
R3462 GND.n6298 GND.n6297 301.784
R3463 GND.n6298 GND.n241 301.784
R3464 GND.n6306 GND.n241 301.784
R3465 GND.n6307 GND.n6306 301.784
R3466 GND.n6308 GND.n6307 301.784
R3467 GND.n6308 GND.n235 301.784
R3468 GND.n6316 GND.n235 301.784
R3469 GND.n6317 GND.n6316 301.784
R3470 GND.n6318 GND.n6317 301.784
R3471 GND.n6318 GND.n229 301.784
R3472 GND.n6326 GND.n229 301.784
R3473 GND.n6327 GND.n6326 301.784
R3474 GND.n6328 GND.n6327 301.784
R3475 GND.n6328 GND.n223 301.784
R3476 GND.n6337 GND.n223 301.784
R3477 GND.n6338 GND.n6337 301.784
R3478 GND.n6339 GND.n6338 301.784
R3479 GND.n6339 GND.n217 301.784
R3480 GND.n5466 GND.n745 280.613
R3481 GND.n5467 GND.n5466 280.613
R3482 GND.n5468 GND.n5467 280.613
R3483 GND.n5468 GND.n739 280.613
R3484 GND.n5476 GND.n739 280.613
R3485 GND.n5477 GND.n5476 280.613
R3486 GND.n5478 GND.n5477 280.613
R3487 GND.n5478 GND.n733 280.613
R3488 GND.n5486 GND.n733 280.613
R3489 GND.n5487 GND.n5486 280.613
R3490 GND.n5488 GND.n5487 280.613
R3491 GND.n5488 GND.n727 280.613
R3492 GND.n5496 GND.n727 280.613
R3493 GND.n5497 GND.n5496 280.613
R3494 GND.n5498 GND.n5497 280.613
R3495 GND.n5498 GND.n721 280.613
R3496 GND.n5506 GND.n721 280.613
R3497 GND.n5507 GND.n5506 280.613
R3498 GND.n5508 GND.n5507 280.613
R3499 GND.n5508 GND.n715 280.613
R3500 GND.n5516 GND.n715 280.613
R3501 GND.n5517 GND.n5516 280.613
R3502 GND.n5518 GND.n5517 280.613
R3503 GND.n5518 GND.n709 280.613
R3504 GND.n5526 GND.n709 280.613
R3505 GND.n5527 GND.n5526 280.613
R3506 GND.n5528 GND.n5527 280.613
R3507 GND.n5528 GND.n703 280.613
R3508 GND.n5536 GND.n703 280.613
R3509 GND.n5537 GND.n5536 280.613
R3510 GND.n5538 GND.n5537 280.613
R3511 GND.n5538 GND.n697 280.613
R3512 GND.n5546 GND.n697 280.613
R3513 GND.n5547 GND.n5546 280.613
R3514 GND.n5548 GND.n5547 280.613
R3515 GND.n5548 GND.n691 280.613
R3516 GND.n5556 GND.n691 280.613
R3517 GND.n5557 GND.n5556 280.613
R3518 GND.n5558 GND.n5557 280.613
R3519 GND.n5558 GND.n685 280.613
R3520 GND.n5566 GND.n685 280.613
R3521 GND.n5567 GND.n5566 280.613
R3522 GND.n5568 GND.n5567 280.613
R3523 GND.n5568 GND.n679 280.613
R3524 GND.n5576 GND.n679 280.613
R3525 GND.n5577 GND.n5576 280.613
R3526 GND.n5578 GND.n5577 280.613
R3527 GND.n5578 GND.n673 280.613
R3528 GND.n5586 GND.n673 280.613
R3529 GND.n5587 GND.n5586 280.613
R3530 GND.n5588 GND.n5587 280.613
R3531 GND.n5588 GND.n667 280.613
R3532 GND.n5596 GND.n667 280.613
R3533 GND.n5597 GND.n5596 280.613
R3534 GND.n5598 GND.n5597 280.613
R3535 GND.n5598 GND.n661 280.613
R3536 GND.n5606 GND.n661 280.613
R3537 GND.n5607 GND.n5606 280.613
R3538 GND.n5608 GND.n5607 280.613
R3539 GND.n5608 GND.n655 280.613
R3540 GND.n5616 GND.n655 280.613
R3541 GND.n5617 GND.n5616 280.613
R3542 GND.n5618 GND.n5617 280.613
R3543 GND.n5618 GND.n649 280.613
R3544 GND.n5626 GND.n649 280.613
R3545 GND.n5627 GND.n5626 280.613
R3546 GND.n5628 GND.n5627 280.613
R3547 GND.n5628 GND.n643 280.613
R3548 GND.n5636 GND.n643 280.613
R3549 GND.n5637 GND.n5636 280.613
R3550 GND.n5638 GND.n5637 280.613
R3551 GND.n5638 GND.n637 280.613
R3552 GND.n5646 GND.n637 280.613
R3553 GND.n5647 GND.n5646 280.613
R3554 GND.n5648 GND.n5647 280.613
R3555 GND.n5648 GND.n631 280.613
R3556 GND.n5656 GND.n631 280.613
R3557 GND.n5657 GND.n5656 280.613
R3558 GND.n5658 GND.n5657 280.613
R3559 GND.n5658 GND.n625 280.613
R3560 GND.n5666 GND.n625 280.613
R3561 GND.n5667 GND.n5666 280.613
R3562 GND.n5668 GND.n5667 280.613
R3563 GND.n5668 GND.n619 280.613
R3564 GND.n5676 GND.n619 280.613
R3565 GND.n5677 GND.n5676 280.613
R3566 GND.n5678 GND.n5677 280.613
R3567 GND.n5678 GND.n613 280.613
R3568 GND.n5686 GND.n613 280.613
R3569 GND.n5687 GND.n5686 280.613
R3570 GND.n5688 GND.n5687 280.613
R3571 GND.n5688 GND.n607 280.613
R3572 GND.n5696 GND.n607 280.613
R3573 GND.n5697 GND.n5696 280.613
R3574 GND.n5698 GND.n5697 280.613
R3575 GND.n5698 GND.n601 280.613
R3576 GND.n5706 GND.n601 280.613
R3577 GND.n5707 GND.n5706 280.613
R3578 GND.n5708 GND.n5707 280.613
R3579 GND.n5708 GND.n595 280.613
R3580 GND.n5716 GND.n595 280.613
R3581 GND.n5717 GND.n5716 280.613
R3582 GND.n5718 GND.n5717 280.613
R3583 GND.n5718 GND.n589 280.613
R3584 GND.n5726 GND.n589 280.613
R3585 GND.n5727 GND.n5726 280.613
R3586 GND.n5728 GND.n5727 280.613
R3587 GND.n5728 GND.n583 280.613
R3588 GND.n5736 GND.n583 280.613
R3589 GND.n5737 GND.n5736 280.613
R3590 GND.n5738 GND.n5737 280.613
R3591 GND.n5738 GND.n577 280.613
R3592 GND.n5746 GND.n577 280.613
R3593 GND.n5747 GND.n5746 280.613
R3594 GND.n5748 GND.n5747 280.613
R3595 GND.n5748 GND.n571 280.613
R3596 GND.n5756 GND.n571 280.613
R3597 GND.n5757 GND.n5756 280.613
R3598 GND.n5758 GND.n5757 280.613
R3599 GND.n5758 GND.n565 280.613
R3600 GND.n5766 GND.n565 280.613
R3601 GND.n5767 GND.n5766 280.613
R3602 GND.n5768 GND.n5767 280.613
R3603 GND.n5768 GND.n559 280.613
R3604 GND.n5776 GND.n559 280.613
R3605 GND.n5777 GND.n5776 280.613
R3606 GND.n5778 GND.n5777 280.613
R3607 GND.n5778 GND.n553 280.613
R3608 GND.n5786 GND.n553 280.613
R3609 GND.n5787 GND.n5786 280.613
R3610 GND.n5788 GND.n5787 280.613
R3611 GND.n5788 GND.n547 280.613
R3612 GND.n5796 GND.n547 280.613
R3613 GND.n5797 GND.n5796 280.613
R3614 GND.n5798 GND.n5797 280.613
R3615 GND.n5798 GND.n541 280.613
R3616 GND.n5806 GND.n541 280.613
R3617 GND.n5807 GND.n5806 280.613
R3618 GND.n5808 GND.n5807 280.613
R3619 GND.n5808 GND.n535 280.613
R3620 GND.n5816 GND.n535 280.613
R3621 GND.n5817 GND.n5816 280.613
R3622 GND.n5818 GND.n5817 280.613
R3623 GND.n5818 GND.n529 280.613
R3624 GND.n5826 GND.n529 280.613
R3625 GND.n5827 GND.n5826 280.613
R3626 GND.n5828 GND.n5827 280.613
R3627 GND.n5828 GND.n523 280.613
R3628 GND.n5836 GND.n523 280.613
R3629 GND.n5837 GND.n5836 280.613
R3630 GND.n5838 GND.n5837 280.613
R3631 GND.n5838 GND.n517 280.613
R3632 GND.n5846 GND.n517 280.613
R3633 GND.n5847 GND.n5846 280.613
R3634 GND.n5848 GND.n5847 280.613
R3635 GND.n5848 GND.n511 280.613
R3636 GND.n5856 GND.n511 280.613
R3637 GND.n5857 GND.n5856 280.613
R3638 GND.n5858 GND.n5857 280.613
R3639 GND.n5858 GND.n505 280.613
R3640 GND.n5866 GND.n505 280.613
R3641 GND.n5867 GND.n5866 280.613
R3642 GND.n5868 GND.n5867 280.613
R3643 GND.n5868 GND.n499 280.613
R3644 GND.n5876 GND.n499 280.613
R3645 GND.n5877 GND.n5876 280.613
R3646 GND.n5878 GND.n5877 280.613
R3647 GND.n5878 GND.n493 280.613
R3648 GND.n5886 GND.n493 280.613
R3649 GND.n5887 GND.n5886 280.613
R3650 GND.n5888 GND.n5887 280.613
R3651 GND.n5888 GND.n487 280.613
R3652 GND.n5896 GND.n487 280.613
R3653 GND.n5897 GND.n5896 280.613
R3654 GND.n5898 GND.n5897 280.613
R3655 GND.n5898 GND.n481 280.613
R3656 GND.n5906 GND.n481 280.613
R3657 GND.n5907 GND.n5906 280.613
R3658 GND.n5908 GND.n5907 280.613
R3659 GND.n5908 GND.n475 280.613
R3660 GND.n5916 GND.n475 280.613
R3661 GND.n5917 GND.n5916 280.613
R3662 GND.n5918 GND.n5917 280.613
R3663 GND.n5918 GND.n469 280.613
R3664 GND.n5926 GND.n469 280.613
R3665 GND.n5927 GND.n5926 280.613
R3666 GND.n5928 GND.n5927 280.613
R3667 GND.n5928 GND.n463 280.613
R3668 GND.n5936 GND.n463 280.613
R3669 GND.n5937 GND.n5936 280.613
R3670 GND.n5938 GND.n5937 280.613
R3671 GND.n5938 GND.n457 280.613
R3672 GND.n5946 GND.n457 280.613
R3673 GND.n5947 GND.n5946 280.613
R3674 GND.n5948 GND.n5947 280.613
R3675 GND.n5948 GND.n451 280.613
R3676 GND.n5956 GND.n451 280.613
R3677 GND.n5957 GND.n5956 280.613
R3678 GND.n5958 GND.n5957 280.613
R3679 GND.n5958 GND.n445 280.613
R3680 GND.n5966 GND.n445 280.613
R3681 GND.n5967 GND.n5966 280.613
R3682 GND.n5968 GND.n5967 280.613
R3683 GND.n5968 GND.n439 280.613
R3684 GND.n5976 GND.n439 280.613
R3685 GND.n5977 GND.n5976 280.613
R3686 GND.n5978 GND.n5977 280.613
R3687 GND.n5978 GND.n433 280.613
R3688 GND.n5986 GND.n433 280.613
R3689 GND.n5987 GND.n5986 280.613
R3690 GND.n5988 GND.n5987 280.613
R3691 GND.n5988 GND.n427 280.613
R3692 GND.n5996 GND.n427 280.613
R3693 GND.n5997 GND.n5996 280.613
R3694 GND.n5998 GND.n5997 280.613
R3695 GND.n5998 GND.n421 280.613
R3696 GND.n6006 GND.n421 280.613
R3697 GND.n6007 GND.n6006 280.613
R3698 GND.n6008 GND.n6007 280.613
R3699 GND.n6008 GND.n415 280.613
R3700 GND.n6016 GND.n415 280.613
R3701 GND.n6017 GND.n6016 280.613
R3702 GND.n6018 GND.n6017 280.613
R3703 GND.n6018 GND.n409 280.613
R3704 GND.n6026 GND.n409 280.613
R3705 GND.n6027 GND.n6026 280.613
R3706 GND.n6028 GND.n6027 280.613
R3707 GND.n6028 GND.n403 280.613
R3708 GND.n6036 GND.n403 280.613
R3709 GND.n6037 GND.n6036 280.613
R3710 GND.n6038 GND.n6037 280.613
R3711 GND.n6038 GND.n397 280.613
R3712 GND.n6046 GND.n397 280.613
R3713 GND.n6047 GND.n6046 280.613
R3714 GND.n6048 GND.n6047 280.613
R3715 GND.n6048 GND.n391 280.613
R3716 GND.n6056 GND.n391 280.613
R3717 GND.n6057 GND.n6056 280.613
R3718 GND.n6058 GND.n6057 280.613
R3719 GND.n6058 GND.n385 280.613
R3720 GND.n6066 GND.n385 280.613
R3721 GND.n6067 GND.n6066 280.613
R3722 GND.n6068 GND.n6067 280.613
R3723 GND.n6068 GND.n379 280.613
R3724 GND.n6076 GND.n379 280.613
R3725 GND.n6077 GND.n6076 280.613
R3726 GND.n6078 GND.n6077 280.613
R3727 GND.n6078 GND.n373 280.613
R3728 GND.n6086 GND.n373 280.613
R3729 GND.n6087 GND.n6086 280.613
R3730 GND.n6088 GND.n6087 280.613
R3731 GND.n6088 GND.n367 280.613
R3732 GND.n6096 GND.n367 280.613
R3733 GND.n6097 GND.n6096 280.613
R3734 GND.n6098 GND.n6097 280.613
R3735 GND.n6098 GND.n361 280.613
R3736 GND.n6106 GND.n361 280.613
R3737 GND.n6107 GND.n6106 280.613
R3738 GND.n6108 GND.n6107 280.613
R3739 GND.n6108 GND.n355 280.613
R3740 GND.n6116 GND.n355 280.613
R3741 GND.n6117 GND.n6116 280.613
R3742 GND.n6118 GND.n6117 280.613
R3743 GND.n6118 GND.n349 280.613
R3744 GND.n6126 GND.n349 280.613
R3745 GND.n6127 GND.n6126 280.613
R3746 GND.n6128 GND.n6127 280.613
R3747 GND.n6128 GND.n343 280.613
R3748 GND.n6136 GND.n343 280.613
R3749 GND.n6137 GND.n6136 280.613
R3750 GND.n6138 GND.n6137 280.613
R3751 GND.n6138 GND.n337 280.613
R3752 GND.n6146 GND.n337 280.613
R3753 GND.n6147 GND.n6146 280.613
R3754 GND.n6148 GND.n6147 280.613
R3755 GND.n6148 GND.n331 280.613
R3756 GND.n6156 GND.n331 280.613
R3757 GND.n6157 GND.n6156 280.613
R3758 GND.n6158 GND.n6157 280.613
R3759 GND.n6158 GND.n325 280.613
R3760 GND.n6166 GND.n325 280.613
R3761 GND.n6167 GND.n6166 280.613
R3762 GND.n6168 GND.n6167 280.613
R3763 GND.n6168 GND.n319 280.613
R3764 GND.n6176 GND.n319 280.613
R3765 GND.n6177 GND.n6176 280.613
R3766 GND.n6178 GND.n6177 280.613
R3767 GND.n6178 GND.n313 280.613
R3768 GND.n6186 GND.n313 280.613
R3769 GND.n6187 GND.n6186 280.613
R3770 GND.n6188 GND.n6187 280.613
R3771 GND.n2275 GND.t123 270.978
R3772 GND.n2833 GND.t84 270.978
R3773 GND.n2020 GND.t80 267.928
R3774 GND.n107 GND.t133 267.928
R3775 GND.n131 GND.t111 267.928
R3776 GND.n1191 GND.t88 267.928
R3777 GND.n1217 GND.t62 267.928
R3778 GND.n1272 GND.t91 267.928
R3779 GND.n3054 GND.t108 267.928
R3780 GND.n2405 GND.t127 267.928
R3781 GND.n2432 GND.t101 267.928
R3782 GND.n987 GND.t76 267.928
R3783 GND.n1007 GND.t130 267.928
R3784 GND.n2501 GND.t105 267.928
R3785 GND.n3646 GND.n3645 256.663
R3786 GND.n3646 GND.n2718 256.663
R3787 GND.n3646 GND.n2719 256.663
R3788 GND.n3646 GND.n2720 256.663
R3789 GND.n3646 GND.n2721 256.663
R3790 GND.n3646 GND.n2722 256.663
R3791 GND.n3646 GND.n2723 256.663
R3792 GND.n3646 GND.n2724 256.663
R3793 GND.n3646 GND.n2725 256.663
R3794 GND.n3646 GND.n2726 256.663
R3795 GND.n3646 GND.n2727 256.663
R3796 GND.n3646 GND.n2728 256.663
R3797 GND.n3646 GND.n2729 256.663
R3798 GND.n3646 GND.n2730 256.663
R3799 GND.n3646 GND.n2731 256.663
R3800 GND.n3646 GND.n2732 256.663
R3801 GND.n3646 GND.n2733 256.663
R3802 GND.n2734 GND.n1195 256.663
R3803 GND.n3646 GND.n2735 256.663
R3804 GND.n3646 GND.n2736 256.663
R3805 GND.n3646 GND.n2737 256.663
R3806 GND.n3646 GND.n2738 256.663
R3807 GND.n3646 GND.n2739 256.663
R3808 GND.n3646 GND.n2740 256.663
R3809 GND.n3646 GND.n2741 256.663
R3810 GND.n3646 GND.n2742 256.663
R3811 GND.n3646 GND.n2743 256.663
R3812 GND.n3646 GND.n2744 256.663
R3813 GND.n3646 GND.n2745 256.663
R3814 GND.n3646 GND.n2746 256.663
R3815 GND.n3646 GND.n2747 256.663
R3816 GND.n3646 GND.n2748 256.663
R3817 GND.n3646 GND.n2749 256.663
R3818 GND.n3646 GND.n2816 256.663
R3819 GND.n3647 GND.n3646 256.663
R3820 GND.n4017 GND.n1757 256.663
R3821 GND.n4023 GND.n1757 256.663
R3822 GND.n2606 GND.n1757 256.663
R3823 GND.n4030 GND.n1757 256.663
R3824 GND.n2603 GND.n1757 256.663
R3825 GND.n4037 GND.n1757 256.663
R3826 GND.n2600 GND.n1757 256.663
R3827 GND.n4044 GND.n1757 256.663
R3828 GND.n2597 GND.n1757 256.663
R3829 GND.n4051 GND.n1757 256.663
R3830 GND.n2594 GND.n1757 256.663
R3831 GND.n4058 GND.n1757 256.663
R3832 GND.n2591 GND.n1757 256.663
R3833 GND.n4065 GND.n1757 256.663
R3834 GND.n2588 GND.n1757 256.663
R3835 GND.n4073 GND.n1757 256.663
R3836 GND.n4076 GND.n1757 256.663
R3837 GND.n4078 GND.n4077 256.663
R3838 GND.n2582 GND.n1757 256.663
R3839 GND.n4081 GND.n1757 256.663
R3840 GND.n2351 GND.n1757 256.663
R3841 GND.n4089 GND.n1757 256.663
R3842 GND.n2346 GND.n1757 256.663
R3843 GND.n4096 GND.n1757 256.663
R3844 GND.n2343 GND.n1757 256.663
R3845 GND.n4103 GND.n1757 256.663
R3846 GND.n2340 GND.n1757 256.663
R3847 GND.n4110 GND.n1757 256.663
R3848 GND.n2337 GND.n1757 256.663
R3849 GND.n4117 GND.n1757 256.663
R3850 GND.n2334 GND.n1757 256.663
R3851 GND.n4124 GND.n1757 256.663
R3852 GND.n2331 GND.n1757 256.663
R3853 GND.n4131 GND.n1757 256.663
R3854 GND.n4134 GND.n1757 256.663
R3855 GND.n2751 GND.t69 244.112
R3856 GND.n2585 GND.t120 244.112
R3857 GND.n3577 GND.t117 244.112
R3858 GND.n2348 GND.t94 244.112
R3859 GND.n5030 GND.n5029 242.672
R3860 GND.n5029 GND.n1234 242.672
R3861 GND.n5029 GND.n1235 242.672
R3862 GND.n5029 GND.n1236 242.672
R3863 GND.n5029 GND.n1237 242.672
R3864 GND.n5029 GND.n1238 242.672
R3865 GND.n5029 GND.n1239 242.672
R3866 GND.n5029 GND.n1240 242.672
R3867 GND.n5029 GND.n1241 242.672
R3868 GND.n5029 GND.n1242 242.672
R3869 GND.n5029 GND.n1243 242.672
R3870 GND.n5029 GND.n1244 242.672
R3871 GND.n5029 GND.n1245 242.672
R3872 GND.n5029 GND.n1246 242.672
R3873 GND.n4189 GND.n1871 242.672
R3874 GND.n2278 GND.n1871 242.672
R3875 GND.n2273 GND.n1871 242.672
R3876 GND.n2268 GND.n1871 242.672
R3877 GND.n2265 GND.n1871 242.672
R3878 GND.n2260 GND.n1871 242.672
R3879 GND.n2257 GND.n1871 242.672
R3880 GND.n2252 GND.n1871 242.672
R3881 GND.n2490 GND.n1871 242.672
R3882 GND.n2489 GND.n1871 242.672
R3883 GND.n2486 GND.n1871 242.672
R3884 GND.n2476 GND.n1871 242.672
R3885 GND.n2464 GND.n1871 242.672
R3886 GND.n2461 GND.n1871 242.672
R3887 GND.n5264 GND.n958 242.672
R3888 GND.n5264 GND.n959 242.672
R3889 GND.n5264 GND.n960 242.672
R3890 GND.n5264 GND.n961 242.672
R3891 GND.n5264 GND.n962 242.672
R3892 GND.n5264 GND.n963 242.672
R3893 GND.n5264 GND.n964 242.672
R3894 GND.n5264 GND.n965 242.672
R3895 GND.n5005 GND.n5004 242.672
R3896 GND.n5004 GND.n1290 242.672
R3897 GND.n5004 GND.n1288 242.672
R3898 GND.n5004 GND.n1286 242.672
R3899 GND.n5004 GND.n1285 242.672
R3900 GND.n5004 GND.n1280 242.672
R3901 GND.n5004 GND.n1279 242.672
R3902 GND.n5004 GND.n1277 242.672
R3903 GND.n5264 GND.n5263 242.672
R3904 GND.n5264 GND.n942 242.672
R3905 GND.n5264 GND.n943 242.672
R3906 GND.n5264 GND.n944 242.672
R3907 GND.n5264 GND.n945 242.672
R3908 GND.n5264 GND.n946 242.672
R3909 GND.n5264 GND.n947 242.672
R3910 GND.n5264 GND.n948 242.672
R3911 GND.n5264 GND.n949 242.672
R3912 GND.n5264 GND.n950 242.672
R3913 GND.n5264 GND.n951 242.672
R3914 GND.n5264 GND.n952 242.672
R3915 GND.n5264 GND.n953 242.672
R3916 GND.n5264 GND.n954 242.672
R3917 GND.n5264 GND.n955 242.672
R3918 GND.n5264 GND.n956 242.672
R3919 GND.n5264 GND.n957 242.672
R3920 GND.n5004 GND.n4980 242.672
R3921 GND.n5004 GND.n4981 242.672
R3922 GND.n5004 GND.n4983 242.672
R3923 GND.n5004 GND.n4984 242.672
R3924 GND.n5004 GND.n4986 242.672
R3925 GND.n5004 GND.n4987 242.672
R3926 GND.n5004 GND.n4989 242.672
R3927 GND.n5004 GND.n4990 242.672
R3928 GND.n5004 GND.n4992 242.672
R3929 GND.n5004 GND.n4993 242.672
R3930 GND.n5075 GND.n1194 242.672
R3931 GND.n5004 GND.n4994 242.672
R3932 GND.n5004 GND.n4996 242.672
R3933 GND.n5004 GND.n4997 242.672
R3934 GND.n5004 GND.n4999 242.672
R3935 GND.n5004 GND.n5000 242.672
R3936 GND.n5004 GND.n5002 242.672
R3937 GND.n5004 GND.n5003 242.672
R3938 GND.n2366 GND.n1872 242.672
R3939 GND.n2375 GND.n1872 242.672
R3940 GND.n2377 GND.n1872 242.672
R3941 GND.n2385 GND.n1872 242.672
R3942 GND.n2387 GND.n1872 242.672
R3943 GND.n2395 GND.n1872 242.672
R3944 GND.n2399 GND.n1872 242.672
R3945 GND.n2581 GND.n2355 242.672
R3946 GND.n2578 GND.n1872 242.672
R3947 GND.n2576 GND.n1872 242.672
R3948 GND.n2570 GND.n1872 242.672
R3949 GND.n2568 GND.n1872 242.672
R3950 GND.n2562 GND.n1872 242.672
R3951 GND.n2560 GND.n1872 242.672
R3952 GND.n2554 GND.n1872 242.672
R3953 GND.n2552 GND.n1872 242.672
R3954 GND.n2546 GND.n1872 242.672
R3955 GND.n2544 GND.n1872 242.672
R3956 GND.n6445 GND.n6444 242.672
R3957 GND.n6444 GND.n6421 242.672
R3958 GND.n6444 GND.n6422 242.672
R3959 GND.n6444 GND.n6424 242.672
R3960 GND.n6444 GND.n6425 242.672
R3961 GND.n6444 GND.n6427 242.672
R3962 GND.n6444 GND.n6428 242.672
R3963 GND.n6444 GND.n6430 242.672
R3964 GND.n6444 GND.n6431 242.672
R3965 GND.n6444 GND.n6433 242.672
R3966 GND.n6444 GND.n6434 242.672
R3967 GND.n6444 GND.n6436 242.672
R3968 GND.n6444 GND.n6437 242.672
R3969 GND.n6444 GND.n6439 242.672
R3970 GND.n6444 GND.n6440 242.672
R3971 GND.n6444 GND.n6442 242.672
R3972 GND.n6444 GND.n6443 242.672
R3973 GND.n2535 GND.n1872 242.672
R3974 GND.n2444 GND.n1872 242.672
R3975 GND.n2453 GND.n1872 242.672
R3976 GND.n2456 GND.n1872 242.672
R3977 GND.n2468 GND.n1872 242.672
R3978 GND.n2471 GND.n1872 242.672
R3979 GND.n2482 GND.n1872 242.672
R3980 GND.n2499 GND.n1872 242.672
R3981 GND.n6444 GND.n143 242.672
R3982 GND.n6444 GND.n142 242.672
R3983 GND.n6444 GND.n141 242.672
R3984 GND.n6444 GND.n140 242.672
R3985 GND.n6444 GND.n139 242.672
R3986 GND.n6444 GND.n138 242.672
R3987 GND.n6444 GND.n137 242.672
R3988 GND.n6444 GND.n136 242.672
R3989 GND.n88 GND.n84 240.244
R3990 GND.n6441 GND.n89 240.244
R3991 GND.n93 GND.n92 240.244
R3992 GND.n6438 GND.n94 240.244
R3993 GND.n98 GND.n97 240.244
R3994 GND.n6435 GND.n99 240.244
R3995 GND.n103 GND.n102 240.244
R3996 GND.n6432 GND.n104 240.244
R3997 GND.n111 GND.n110 240.244
R3998 GND.n6429 GND.n112 240.244
R3999 GND.n116 GND.n115 240.244
R4000 GND.n6426 GND.n117 240.244
R4001 GND.n121 GND.n120 240.244
R4002 GND.n6423 GND.n122 240.244
R4003 GND.n126 GND.n125 240.244
R4004 GND.n6420 GND.n127 240.244
R4005 GND.n133 GND.n130 240.244
R4006 GND.n2244 GND.n1881 240.244
R4007 GND.n2244 GND.n1893 240.244
R4008 GND.n1903 GND.n1893 240.244
R4009 GND.n1904 GND.n1903 240.244
R4010 GND.n2238 GND.n1904 240.244
R4011 GND.n2238 GND.n1910 240.244
R4012 GND.n1911 GND.n1910 240.244
R4013 GND.n1912 GND.n1911 240.244
R4014 GND.n2226 GND.n1912 240.244
R4015 GND.n2226 GND.n1918 240.244
R4016 GND.n1919 GND.n1918 240.244
R4017 GND.n1920 GND.n1919 240.244
R4018 GND.n2201 GND.n1920 240.244
R4019 GND.n2201 GND.n1926 240.244
R4020 GND.n1927 GND.n1926 240.244
R4021 GND.n1928 GND.n1927 240.244
R4022 GND.n4341 GND.n1928 240.244
R4023 GND.n4341 GND.n1934 240.244
R4024 GND.n1935 GND.n1934 240.244
R4025 GND.n1936 GND.n1935 240.244
R4026 GND.n4361 GND.n1936 240.244
R4027 GND.n4361 GND.n1942 240.244
R4028 GND.n1943 GND.n1942 240.244
R4029 GND.n1944 GND.n1943 240.244
R4030 GND.n2170 GND.n1944 240.244
R4031 GND.n2170 GND.n1950 240.244
R4032 GND.n1951 GND.n1950 240.244
R4033 GND.n1952 GND.n1951 240.244
R4034 GND.n4385 GND.n1952 240.244
R4035 GND.n4385 GND.n1958 240.244
R4036 GND.n1959 GND.n1958 240.244
R4037 GND.n1960 GND.n1959 240.244
R4038 GND.n2117 GND.n1960 240.244
R4039 GND.n2117 GND.n1966 240.244
R4040 GND.n1967 GND.n1966 240.244
R4041 GND.n1968 GND.n1967 240.244
R4042 GND.n2105 GND.n1968 240.244
R4043 GND.n2105 GND.n1974 240.244
R4044 GND.n1975 GND.n1974 240.244
R4045 GND.n1976 GND.n1975 240.244
R4046 GND.n4494 GND.n1976 240.244
R4047 GND.n4494 GND.n1982 240.244
R4048 GND.n1983 GND.n1982 240.244
R4049 GND.n1984 GND.n1983 240.244
R4050 GND.n2066 GND.n1984 240.244
R4051 GND.n2066 GND.n1990 240.244
R4052 GND.n1991 GND.n1990 240.244
R4053 GND.n1992 GND.n1991 240.244
R4054 GND.n2052 GND.n1992 240.244
R4055 GND.n4555 GND.n2052 240.244
R4056 GND.n4555 GND.n80 240.244
R4057 GND.n2374 GND.n2367 240.244
R4058 GND.n2378 GND.n2376 240.244
R4059 GND.n2384 GND.n2362 240.244
R4060 GND.n2388 GND.n2386 240.244
R4061 GND.n2394 GND.n2358 240.244
R4062 GND.n2400 GND.n2396 240.244
R4063 GND.n2398 GND.n2397 240.244
R4064 GND.n2579 GND.n2577 240.244
R4065 GND.n2575 GND.n2409 240.244
R4066 GND.n2571 GND.n2569 240.244
R4067 GND.n2567 GND.n2415 240.244
R4068 GND.n2563 GND.n2561 240.244
R4069 GND.n2559 GND.n2421 240.244
R4070 GND.n2555 GND.n2553 240.244
R4071 GND.n2551 GND.n2427 240.244
R4072 GND.n2547 GND.n2545 240.244
R4073 GND.n4638 GND.n1886 240.244
R4074 GND.n4634 GND.n1886 240.244
R4075 GND.n4634 GND.n1891 240.244
R4076 GND.n4225 GND.n1891 240.244
R4077 GND.n4225 GND.n2232 240.244
R4078 GND.n4296 GND.n2232 240.244
R4079 GND.n4296 GND.n2225 240.244
R4080 GND.n4304 GND.n2225 240.244
R4081 GND.n4304 GND.n2228 240.244
R4082 GND.n2228 GND.n2210 240.244
R4083 GND.n4321 GND.n2210 240.244
R4084 GND.n4321 GND.n2204 240.244
R4085 GND.n4329 GND.n2204 240.244
R4086 GND.n4329 GND.n2206 240.244
R4087 GND.n2206 GND.n2187 240.244
R4088 GND.n4346 GND.n2187 240.244
R4089 GND.n4346 GND.n2183 240.244
R4090 GND.n4353 GND.n2183 240.244
R4091 GND.n4353 GND.n2151 240.244
R4092 GND.n4429 GND.n2151 240.244
R4093 GND.n4429 GND.n2152 240.244
R4094 GND.n4424 GND.n2152 240.244
R4095 GND.n4424 GND.n2156 240.244
R4096 GND.n4374 GND.n2156 240.244
R4097 GND.n4412 GND.n4374 240.244
R4098 GND.n4412 GND.n4375 240.244
R4099 GND.n4407 GND.n4375 240.244
R4100 GND.n4407 GND.n4379 240.244
R4101 GND.n4392 GND.n4379 240.244
R4102 GND.n4392 GND.n4388 240.244
R4103 GND.n4388 GND.n2127 240.244
R4104 GND.n4447 GND.n2127 240.244
R4105 GND.n4447 GND.n2122 240.244
R4106 GND.n4455 GND.n2122 240.244
R4107 GND.n4455 GND.n2123 240.244
R4108 GND.n2123 GND.n2103 240.244
R4109 GND.n4473 GND.n2103 240.244
R4110 GND.n4473 GND.n2098 240.244
R4111 GND.n4481 GND.n2098 240.244
R4112 GND.n4481 GND.n2099 240.244
R4113 GND.n2099 GND.n2083 240.244
R4114 GND.n4502 GND.n2083 240.244
R4115 GND.n4502 GND.n2078 240.244
R4116 GND.n4510 GND.n2078 240.244
R4117 GND.n4510 GND.n2079 240.244
R4118 GND.n2079 GND.n2061 240.244
R4119 GND.n4544 GND.n2061 240.244
R4120 GND.n4544 GND.n2057 240.244
R4121 GND.n4550 GND.n2057 240.244
R4122 GND.n4550 GND.n83 240.244
R4123 GND.n6501 GND.n83 240.244
R4124 GND.n1175 GND.n1171 240.244
R4125 GND.n5001 GND.n1176 240.244
R4126 GND.n1180 GND.n1179 240.244
R4127 GND.n4998 GND.n1181 240.244
R4128 GND.n1185 GND.n1184 240.244
R4129 GND.n4995 GND.n1186 240.244
R4130 GND.n1190 GND.n1189 240.244
R4131 GND.n4991 GND.n1196 240.244
R4132 GND.n1200 GND.n1199 240.244
R4133 GND.n4988 GND.n1201 240.244
R4134 GND.n1205 GND.n1204 240.244
R4135 GND.n4985 GND.n1206 240.244
R4136 GND.n1210 GND.n1209 240.244
R4137 GND.n4982 GND.n1211 240.244
R4138 GND.n1215 GND.n1214 240.244
R4139 GND.n4979 GND.n1216 240.244
R4140 GND.n1065 GND.n1016 240.244
R4141 GND.n1065 GND.n1064 240.244
R4142 GND.n1064 GND.n1034 240.244
R4143 GND.n3106 GND.n1034 240.244
R4144 GND.n3106 GND.n1052 240.244
R4145 GND.n1075 GND.n1052 240.244
R4146 GND.n1076 GND.n1075 240.244
R4147 GND.n3044 GND.n1076 240.244
R4148 GND.n3044 GND.n1082 240.244
R4149 GND.n1083 GND.n1082 240.244
R4150 GND.n1084 GND.n1083 240.244
R4151 GND.n3018 GND.n1084 240.244
R4152 GND.n3018 GND.n1090 240.244
R4153 GND.n1091 GND.n1090 240.244
R4154 GND.n1092 GND.n1091 240.244
R4155 GND.n3002 GND.n1092 240.244
R4156 GND.n3002 GND.n1098 240.244
R4157 GND.n1099 GND.n1098 240.244
R4158 GND.n1100 GND.n1099 240.244
R4159 GND.n3228 GND.n1100 240.244
R4160 GND.n3228 GND.n1106 240.244
R4161 GND.n1107 GND.n1106 240.244
R4162 GND.n1108 GND.n1107 240.244
R4163 GND.n2963 GND.n1108 240.244
R4164 GND.n2963 GND.n1114 240.244
R4165 GND.n1115 GND.n1114 240.244
R4166 GND.n1116 GND.n1115 240.244
R4167 GND.n3250 GND.n1116 240.244
R4168 GND.n3250 GND.n1122 240.244
R4169 GND.n1123 GND.n1122 240.244
R4170 GND.n1124 GND.n1123 240.244
R4171 GND.n2918 GND.n1124 240.244
R4172 GND.n2918 GND.n1130 240.244
R4173 GND.n1131 GND.n1130 240.244
R4174 GND.n1132 GND.n1131 240.244
R4175 GND.n2900 GND.n1132 240.244
R4176 GND.n2900 GND.n1138 240.244
R4177 GND.n1139 GND.n1138 240.244
R4178 GND.n1140 GND.n1139 240.244
R4179 GND.n3354 GND.n1140 240.244
R4180 GND.n3354 GND.n1146 240.244
R4181 GND.n1147 GND.n1146 240.244
R4182 GND.n1148 GND.n1147 240.244
R4183 GND.n2866 GND.n1148 240.244
R4184 GND.n2866 GND.n1154 240.244
R4185 GND.n1155 GND.n1154 240.244
R4186 GND.n1156 GND.n1155 240.244
R4187 GND.n3438 GND.n1156 240.244
R4188 GND.n3438 GND.n1162 240.244
R4189 GND.n1163 GND.n1162 240.244
R4190 GND.n5101 GND.n1163 240.244
R4191 GND.n969 GND.n968 240.244
R4192 GND.n5257 GND.n968 240.244
R4193 GND.n5255 GND.n5254 240.244
R4194 GND.n5251 GND.n5250 240.244
R4195 GND.n5247 GND.n5246 240.244
R4196 GND.n5243 GND.n5242 240.244
R4197 GND.n5239 GND.n5238 240.244
R4198 GND.n5235 GND.n5234 240.244
R4199 GND.n5230 GND.n5229 240.244
R4200 GND.n5226 GND.n5225 240.244
R4201 GND.n5222 GND.n5221 240.244
R4202 GND.n5218 GND.n5217 240.244
R4203 GND.n5214 GND.n5213 240.244
R4204 GND.n5210 GND.n5209 240.244
R4205 GND.n5206 GND.n5205 240.244
R4206 GND.n5202 GND.n5201 240.244
R4207 GND.n5198 GND.n5197 240.244
R4208 GND.n1042 GND.n970 240.244
R4209 GND.n1042 GND.n1037 240.244
R4210 GND.n5179 GND.n1037 240.244
R4211 GND.n5179 GND.n1038 240.244
R4212 GND.n5175 GND.n1038 240.244
R4213 GND.n5175 GND.n1050 240.244
R4214 GND.n3141 GND.n1050 240.244
R4215 GND.n3151 GND.n3141 240.244
R4216 GND.n3151 GND.n3143 240.244
R4217 GND.n3143 GND.n3030 240.244
R4218 GND.n3171 GND.n3030 240.244
R4219 GND.n3171 GND.n3025 240.244
R4220 GND.n3179 GND.n3025 240.244
R4221 GND.n3179 GND.n3026 240.244
R4222 GND.n3026 GND.n3000 240.244
R4223 GND.n3206 GND.n3000 240.244
R4224 GND.n3206 GND.n2995 240.244
R4225 GND.n3214 GND.n2995 240.244
R4226 GND.n3214 GND.n2996 240.244
R4227 GND.n2996 GND.n2949 240.244
R4228 GND.n3285 GND.n2949 240.244
R4229 GND.n3285 GND.n2950 240.244
R4230 GND.n3238 GND.n2950 240.244
R4231 GND.n3238 GND.n2970 240.244
R4232 GND.n3271 GND.n2970 240.244
R4233 GND.n3271 GND.n3268 240.244
R4234 GND.n3268 GND.n2973 240.244
R4235 GND.n2973 GND.n2940 240.244
R4236 GND.n3291 GND.n2940 240.244
R4237 GND.n3291 GND.n2941 240.244
R4238 GND.n2941 GND.n2916 240.244
R4239 GND.n3373 GND.n2916 240.244
R4240 GND.n3373 GND.n2910 240.244
R4241 GND.n3381 GND.n2910 240.244
R4242 GND.n3381 GND.n2912 240.244
R4243 GND.n2912 GND.n2894 240.244
R4244 GND.n3398 GND.n2894 240.244
R4245 GND.n3398 GND.n2889 240.244
R4246 GND.n3406 GND.n2889 240.244
R4247 GND.n3406 GND.n2890 240.244
R4248 GND.n2890 GND.n2875 240.244
R4249 GND.n3423 GND.n2875 240.244
R4250 GND.n3423 GND.n2869 240.244
R4251 GND.n3431 GND.n2869 240.244
R4252 GND.n3431 GND.n2871 240.244
R4253 GND.n2871 GND.n2852 240.244
R4254 GND.n3451 GND.n2852 240.244
R4255 GND.n3451 GND.n2848 240.244
R4256 GND.n3457 GND.n2848 240.244
R4257 GND.n3457 GND.n1170 240.244
R4258 GND.n5099 GND.n1170 240.244
R4259 GND.n1222 GND.n1221 240.244
R4260 GND.n1278 GND.n1223 240.244
R4261 GND.n1227 GND.n1226 240.244
R4262 GND.n1283 GND.n1281 240.244
R4263 GND.n1284 GND.n1254 240.244
R4264 GND.n1287 GND.n1255 240.244
R4265 GND.n1263 GND.n1262 240.244
R4266 GND.n1289 GND.n1274 240.244
R4267 GND.n3050 GND.n1017 240.244
R4268 GND.n3051 GND.n3050 240.244
R4269 GND.n3051 GND.n1035 240.244
R4270 GND.n3108 GND.n1035 240.244
R4271 GND.n3108 GND.n1053 240.244
R4272 GND.n3114 GND.n1053 240.244
R4273 GND.n3114 GND.n3042 240.244
R4274 GND.n3153 GND.n3042 240.244
R4275 GND.n3153 GND.n3037 240.244
R4276 GND.n3165 GND.n3037 240.244
R4277 GND.n3165 GND.n3032 240.244
R4278 GND.n3158 GND.n3032 240.244
R4279 GND.n3158 GND.n3020 240.244
R4280 GND.n3020 GND.n3010 240.244
R4281 GND.n3193 GND.n3010 240.244
R4282 GND.n3193 GND.n3003 240.244
R4283 GND.n3201 GND.n3003 240.244
R4284 GND.n3201 GND.n2990 240.244
R4285 GND.n2990 GND.n2982 240.244
R4286 GND.n3230 GND.n2982 240.244
R4287 GND.n3230 GND.n2952 240.244
R4288 GND.n2957 GND.n2952 240.244
R4289 GND.n3240 GND.n2957 240.244
R4290 GND.n3241 GND.n3240 240.244
R4291 GND.n3241 GND.n2965 240.244
R4292 GND.n2974 GND.n2965 240.244
R4293 GND.n3249 GND.n2974 240.244
R4294 GND.n3249 GND.n2934 240.244
R4295 GND.n3293 GND.n2934 240.244
R4296 GND.n3293 GND.n2929 240.244
R4297 GND.n3300 GND.n2929 240.244
R4298 GND.n3300 GND.n2919 240.244
R4299 GND.n2919 GND.n2906 240.244
R4300 GND.n3383 GND.n2906 240.244
R4301 GND.n3383 GND.n2901 240.244
R4302 GND.n3390 GND.n2901 240.244
R4303 GND.n3390 GND.n2896 240.244
R4304 GND.n2896 GND.n2886 240.244
R4305 GND.n3408 GND.n2886 240.244
R4306 GND.n3408 GND.n2881 240.244
R4307 GND.n3415 GND.n2881 240.244
R4308 GND.n3415 GND.n2877 240.244
R4309 GND.n2877 GND.n2864 240.244
R4310 GND.n3433 GND.n2864 240.244
R4311 GND.n3433 GND.n2859 240.244
R4312 GND.n3446 GND.n2859 240.244
R4313 GND.n3446 GND.n2854 240.244
R4314 GND.n3440 GND.n2854 240.244
R4315 GND.n3440 GND.n2844 240.244
R4316 GND.n3464 GND.n2844 240.244
R4317 GND.n3464 GND.n1167 240.244
R4318 GND.n3069 GND.n3068 240.244
R4319 GND.n3074 GND.n3073 240.244
R4320 GND.n3066 GND.n3065 240.244
R4321 GND.n3082 GND.n3081 240.244
R4322 GND.n3062 GND.n3061 240.244
R4323 GND.n3090 GND.n3089 240.244
R4324 GND.n3058 GND.n3057 240.244
R4325 GND.n3053 GND.n966 240.244
R4326 GND.n5189 GND.n1012 240.244
R4327 GND.n1069 GND.n1012 240.244
R4328 GND.n1069 GND.n1036 240.244
R4329 GND.n1055 GND.n1036 240.244
R4330 GND.n5173 GND.n1055 240.244
R4331 GND.n5173 GND.n1056 240.244
R4332 GND.n3139 GND.n1056 240.244
R4333 GND.n3139 GND.n3046 240.244
R4334 GND.n3046 GND.n3034 240.244
R4335 GND.n3167 GND.n3034 240.244
R4336 GND.n3169 GND.n3167 240.244
R4337 GND.n3169 GND.n3168 240.244
R4338 GND.n3168 GND.n3024 240.244
R4339 GND.n3024 GND.n3023 240.244
R4340 GND.n3023 GND.n3005 240.244
R4341 GND.n3204 GND.n3005 240.244
R4342 GND.n3204 GND.n3203 240.244
R4343 GND.n3203 GND.n2994 240.244
R4344 GND.n2994 GND.n2992 240.244
R4345 GND.n2992 GND.n2954 240.244
R4346 GND.n3283 GND.n2954 240.244
R4347 GND.n3283 GND.n3282 240.244
R4348 GND.n3282 GND.n2955 240.244
R4349 GND.n2967 GND.n2955 240.244
R4350 GND.n2968 GND.n2967 240.244
R4351 GND.n3266 GND.n2968 240.244
R4352 GND.n3266 GND.n3264 240.244
R4353 GND.n3264 GND.n2976 240.244
R4354 GND.n2976 GND.n2939 240.244
R4355 GND.n2939 GND.n2938 240.244
R4356 GND.n2938 GND.n2921 240.244
R4357 GND.n3371 GND.n2921 240.244
R4358 GND.n3371 GND.n3370 240.244
R4359 GND.n3370 GND.n2909 240.244
R4360 GND.n2909 GND.n2898 240.244
R4361 GND.n3392 GND.n2898 240.244
R4362 GND.n3396 GND.n3392 240.244
R4363 GND.n3396 GND.n3395 240.244
R4364 GND.n3395 GND.n2888 240.244
R4365 GND.n2888 GND.n2879 240.244
R4366 GND.n3417 GND.n2879 240.244
R4367 GND.n3421 GND.n3417 240.244
R4368 GND.n3421 GND.n3419 240.244
R4369 GND.n3419 GND.n2868 240.244
R4370 GND.n2868 GND.n2856 240.244
R4371 GND.n3448 GND.n2856 240.244
R4372 GND.n3449 GND.n3448 240.244
R4373 GND.n3449 GND.n2846 240.244
R4374 GND.n3459 GND.n2846 240.244
R4375 GND.n3462 GND.n3459 240.244
R4376 GND.n3462 GND.n1169 240.244
R4377 GND.n2449 GND.n1857 240.244
R4378 GND.n2463 GND.n2462 240.244
R4379 GND.n2475 GND.n2465 240.244
R4380 GND.n2478 GND.n2477 240.244
R4381 GND.n2488 GND.n2487 240.244
R4382 GND.n2492 GND.n2491 240.244
R4383 GND.n2251 GND.n2250 240.244
R4384 GND.n2256 GND.n2253 240.244
R4385 GND.n2259 GND.n2258 240.244
R4386 GND.n2264 GND.n2261 240.244
R4387 GND.n2267 GND.n2266 240.244
R4388 GND.n2272 GND.n2269 240.244
R4389 GND.n2277 GND.n2274 240.244
R4390 GND.n4188 GND.n2279 240.244
R4391 GND.n1302 GND.n1301 240.244
R4392 GND.n3522 GND.n1302 240.244
R4393 GND.n3522 GND.n1313 240.244
R4394 GND.n3528 GND.n1313 240.244
R4395 GND.n3529 GND.n3528 240.244
R4396 GND.n3529 GND.n1333 240.244
R4397 GND.n2827 GND.n1333 240.244
R4398 GND.n2827 GND.n1346 240.244
R4399 GND.n3537 GND.n1346 240.244
R4400 GND.n3538 GND.n3537 240.244
R4401 GND.n3538 GND.n1360 240.244
R4402 GND.n2824 GND.n1360 240.244
R4403 GND.n2824 GND.n1373 240.244
R4404 GND.n3546 GND.n1373 240.244
R4405 GND.n3546 GND.n3545 240.244
R4406 GND.n3545 GND.n1387 240.244
R4407 GND.n3553 GND.n1387 240.244
R4408 GND.n3553 GND.n1400 240.244
R4409 GND.n2817 GND.n1400 240.244
R4410 GND.n3560 GND.n2817 240.244
R4411 GND.n3560 GND.n1413 240.244
R4412 GND.n3657 GND.n1413 240.244
R4413 GND.n3657 GND.n1426 240.244
R4414 GND.n3663 GND.n1426 240.244
R4415 GND.n3663 GND.n1436 240.244
R4416 GND.n3704 GND.n1436 240.244
R4417 GND.n3704 GND.n1446 240.244
R4418 GND.n3710 GND.n1446 240.244
R4419 GND.n3710 GND.n1456 240.244
R4420 GND.n3742 GND.n1456 240.244
R4421 GND.n3742 GND.n1466 240.244
R4422 GND.n3727 GND.n1466 240.244
R4423 GND.n3727 GND.n1476 240.244
R4424 GND.n3728 GND.n1476 240.244
R4425 GND.n3728 GND.n1486 240.244
R4426 GND.n3730 GND.n1486 240.244
R4427 GND.n3730 GND.n1495 240.244
R4428 GND.n3793 GND.n1495 240.244
R4429 GND.n3793 GND.n1505 240.244
R4430 GND.n3808 GND.n1505 240.244
R4431 GND.n3808 GND.n1515 240.244
R4432 GND.n3801 GND.n1515 240.244
R4433 GND.n3801 GND.n1525 240.244
R4434 GND.n3839 GND.n1525 240.244
R4435 GND.n3840 GND.n3839 240.244
R4436 GND.n3841 GND.n3840 240.244
R4437 GND.n3841 GND.n1545 240.244
R4438 GND.n3851 GND.n1545 240.244
R4439 GND.n3851 GND.n1562 240.244
R4440 GND.n3845 GND.n1562 240.244
R4441 GND.n3845 GND.n2650 240.244
R4442 GND.n3877 GND.n2650 240.244
R4443 GND.n3877 GND.n1589 240.244
R4444 GND.n3904 GND.n1589 240.244
R4445 GND.n3904 GND.n1605 240.244
R4446 GND.n3882 GND.n1605 240.244
R4447 GND.n3883 GND.n3882 240.244
R4448 GND.n3884 GND.n3883 240.244
R4449 GND.n3885 GND.n3884 240.244
R4450 GND.n3885 GND.n1639 240.244
R4451 GND.n3888 GND.n1639 240.244
R4452 GND.n3888 GND.n1658 240.244
R4453 GND.n3964 GND.n1658 240.244
R4454 GND.n3965 GND.n3964 240.244
R4455 GND.n3966 GND.n3965 240.244
R4456 GND.n3966 GND.n1683 240.244
R4457 GND.n2630 GND.n1683 240.244
R4458 GND.n2630 GND.n1699 240.244
R4459 GND.n3973 GND.n1699 240.244
R4460 GND.n3973 GND.n2626 240.244
R4461 GND.n3979 GND.n2626 240.244
R4462 GND.n3979 GND.n1726 240.244
R4463 GND.n3999 GND.n1726 240.244
R4464 GND.n3999 GND.n1737 240.244
R4465 GND.n4006 GND.n1737 240.244
R4466 GND.n4006 GND.n1747 240.244
R4467 GND.n4144 GND.n1747 240.244
R4468 GND.n4144 GND.n1756 240.244
R4469 GND.n2298 GND.n1756 240.244
R4470 GND.n2299 GND.n2298 240.244
R4471 GND.n2299 GND.n1767 240.244
R4472 GND.n4153 GND.n1767 240.244
R4473 GND.n4153 GND.n1780 240.244
R4474 GND.n4159 GND.n1780 240.244
R4475 GND.n4160 GND.n4159 240.244
R4476 GND.n4160 GND.n1794 240.244
R4477 GND.n2290 GND.n1794 240.244
R4478 GND.n2290 GND.n1806 240.244
R4479 GND.n4168 GND.n1806 240.244
R4480 GND.n4169 GND.n4168 240.244
R4481 GND.n4169 GND.n1820 240.244
R4482 GND.n2286 GND.n1820 240.244
R4483 GND.n2286 GND.n1833 240.244
R4484 GND.n4177 GND.n1833 240.244
R4485 GND.n4177 GND.n4176 240.244
R4486 GND.n4176 GND.n1847 240.244
R4487 GND.n4184 GND.n1847 240.244
R4488 GND.n4184 GND.n1859 240.244
R4489 GND.n5028 GND.n1232 240.244
R4490 GND.n5028 GND.n1248 240.244
R4491 GND.n1259 GND.n1258 240.244
R4492 GND.n1267 GND.n1266 240.244
R4493 GND.n1269 GND.n1268 240.244
R4494 GND.n3471 GND.n3470 240.244
R4495 GND.n3476 GND.n3475 240.244
R4496 GND.n3483 GND.n3482 240.244
R4497 GND.n3486 GND.n3485 240.244
R4498 GND.n3493 GND.n3492 240.244
R4499 GND.n3496 GND.n3495 240.244
R4500 GND.n3503 GND.n3502 240.244
R4501 GND.n3506 GND.n3505 240.244
R4502 GND.n3513 GND.n3512 240.244
R4503 GND.n4966 GND.n1231 240.244
R4504 GND.n4966 GND.n1304 240.244
R4505 GND.n4962 GND.n1304 240.244
R4506 GND.n4962 GND.n1311 240.244
R4507 GND.n1335 GND.n1311 240.244
R4508 GND.n4952 GND.n1335 240.244
R4509 GND.n4952 GND.n1336 240.244
R4510 GND.n4948 GND.n1336 240.244
R4511 GND.n4948 GND.n1344 240.244
R4512 GND.n1362 GND.n1344 240.244
R4513 GND.n4938 GND.n1362 240.244
R4514 GND.n4938 GND.n1363 240.244
R4515 GND.n4934 GND.n1363 240.244
R4516 GND.n4934 GND.n1371 240.244
R4517 GND.n1389 GND.n1371 240.244
R4518 GND.n4924 GND.n1389 240.244
R4519 GND.n4924 GND.n1390 240.244
R4520 GND.n4920 GND.n1390 240.244
R4521 GND.n4920 GND.n1398 240.244
R4522 GND.n1415 GND.n1398 240.244
R4523 GND.n4910 GND.n1415 240.244
R4524 GND.n4910 GND.n1416 240.244
R4525 GND.n4906 GND.n1416 240.244
R4526 GND.n4906 GND.n1424 240.244
R4527 GND.n4896 GND.n1424 240.244
R4528 GND.n4896 GND.n1438 240.244
R4529 GND.n4892 GND.n1438 240.244
R4530 GND.n4892 GND.n1444 240.244
R4531 GND.n4882 GND.n1444 240.244
R4532 GND.n4882 GND.n1458 240.244
R4533 GND.n4878 GND.n1458 240.244
R4534 GND.n4878 GND.n1464 240.244
R4535 GND.n4868 GND.n1464 240.244
R4536 GND.n4868 GND.n1478 240.244
R4537 GND.n4864 GND.n1478 240.244
R4538 GND.n4864 GND.n1484 240.244
R4539 GND.n4854 GND.n1484 240.244
R4540 GND.n4854 GND.n1497 240.244
R4541 GND.n4850 GND.n1497 240.244
R4542 GND.n4850 GND.n1503 240.244
R4543 GND.n4840 GND.n1503 240.244
R4544 GND.n4840 GND.n1517 240.244
R4545 GND.n4836 GND.n1517 240.244
R4546 GND.n4836 GND.n1523 240.244
R4547 GND.n1551 GND.n1523 240.244
R4548 GND.n1551 GND.n1547 240.244
R4549 GND.n4819 GND.n1547 240.244
R4550 GND.n4819 GND.n1548 240.244
R4551 GND.n4815 GND.n1548 240.244
R4552 GND.n4815 GND.n1559 240.244
R4553 GND.n1595 GND.n1559 240.244
R4554 GND.n1595 GND.n1591 240.244
R4555 GND.n4799 GND.n1591 240.244
R4556 GND.n4799 GND.n1592 240.244
R4557 GND.n4795 GND.n1592 240.244
R4558 GND.n4795 GND.n1603 240.244
R4559 GND.n1647 GND.n1603 240.244
R4560 GND.n1648 GND.n1647 240.244
R4561 GND.n1648 GND.n1641 240.244
R4562 GND.n4771 GND.n1641 240.244
R4563 GND.n4771 GND.n1642 240.244
R4564 GND.n4767 GND.n1642 240.244
R4565 GND.n4767 GND.n1656 240.244
R4566 GND.n1689 GND.n1656 240.244
R4567 GND.n1689 GND.n1685 240.244
R4568 GND.n4751 GND.n1685 240.244
R4569 GND.n4751 GND.n1686 240.244
R4570 GND.n4747 GND.n1686 240.244
R4571 GND.n4747 GND.n1697 240.244
R4572 GND.n2624 GND.n1697 240.244
R4573 GND.n2624 GND.n1728 240.244
R4574 GND.n4730 GND.n1728 240.244
R4575 GND.n4730 GND.n1729 240.244
R4576 GND.n4726 GND.n1729 240.244
R4577 GND.n4726 GND.n1735 240.244
R4578 GND.n4716 GND.n1735 240.244
R4579 GND.n4716 GND.n1749 240.244
R4580 GND.n4712 GND.n1749 240.244
R4581 GND.n4712 GND.n1755 240.244
R4582 GND.n1769 GND.n1755 240.244
R4583 GND.n4702 GND.n1769 240.244
R4584 GND.n4702 GND.n1770 240.244
R4585 GND.n4698 GND.n1770 240.244
R4586 GND.n4698 GND.n1778 240.244
R4587 GND.n1795 GND.n1778 240.244
R4588 GND.n4688 GND.n1795 240.244
R4589 GND.n4688 GND.n1796 240.244
R4590 GND.n4684 GND.n1796 240.244
R4591 GND.n4684 GND.n1804 240.244
R4592 GND.n1822 GND.n1804 240.244
R4593 GND.n4674 GND.n1822 240.244
R4594 GND.n4674 GND.n1823 240.244
R4595 GND.n4670 GND.n1823 240.244
R4596 GND.n4670 GND.n1831 240.244
R4597 GND.n1849 GND.n1831 240.244
R4598 GND.n4660 GND.n1849 240.244
R4599 GND.n4660 GND.n1850 240.244
R4600 GND.n4656 GND.n1850 240.244
R4601 GND.n5465 GND.n746 240.244
R4602 GND.n5465 GND.n744 240.244
R4603 GND.n5469 GND.n744 240.244
R4604 GND.n5469 GND.n740 240.244
R4605 GND.n5475 GND.n740 240.244
R4606 GND.n5475 GND.n738 240.244
R4607 GND.n5479 GND.n738 240.244
R4608 GND.n5479 GND.n734 240.244
R4609 GND.n5485 GND.n734 240.244
R4610 GND.n5485 GND.n732 240.244
R4611 GND.n5489 GND.n732 240.244
R4612 GND.n5489 GND.n728 240.244
R4613 GND.n5495 GND.n728 240.244
R4614 GND.n5495 GND.n726 240.244
R4615 GND.n5499 GND.n726 240.244
R4616 GND.n5499 GND.n722 240.244
R4617 GND.n5505 GND.n722 240.244
R4618 GND.n5505 GND.n720 240.244
R4619 GND.n5509 GND.n720 240.244
R4620 GND.n5509 GND.n716 240.244
R4621 GND.n5515 GND.n716 240.244
R4622 GND.n5515 GND.n714 240.244
R4623 GND.n5519 GND.n714 240.244
R4624 GND.n5519 GND.n710 240.244
R4625 GND.n5525 GND.n710 240.244
R4626 GND.n5525 GND.n708 240.244
R4627 GND.n5529 GND.n708 240.244
R4628 GND.n5529 GND.n704 240.244
R4629 GND.n5535 GND.n704 240.244
R4630 GND.n5535 GND.n702 240.244
R4631 GND.n5539 GND.n702 240.244
R4632 GND.n5539 GND.n698 240.244
R4633 GND.n5545 GND.n698 240.244
R4634 GND.n5545 GND.n696 240.244
R4635 GND.n5549 GND.n696 240.244
R4636 GND.n5549 GND.n692 240.244
R4637 GND.n5555 GND.n692 240.244
R4638 GND.n5555 GND.n690 240.244
R4639 GND.n5559 GND.n690 240.244
R4640 GND.n5559 GND.n686 240.244
R4641 GND.n5565 GND.n686 240.244
R4642 GND.n5565 GND.n684 240.244
R4643 GND.n5569 GND.n684 240.244
R4644 GND.n5569 GND.n680 240.244
R4645 GND.n5575 GND.n680 240.244
R4646 GND.n5575 GND.n678 240.244
R4647 GND.n5579 GND.n678 240.244
R4648 GND.n5579 GND.n674 240.244
R4649 GND.n5585 GND.n674 240.244
R4650 GND.n5585 GND.n672 240.244
R4651 GND.n5589 GND.n672 240.244
R4652 GND.n5589 GND.n668 240.244
R4653 GND.n5595 GND.n668 240.244
R4654 GND.n5595 GND.n666 240.244
R4655 GND.n5599 GND.n666 240.244
R4656 GND.n5599 GND.n662 240.244
R4657 GND.n5605 GND.n662 240.244
R4658 GND.n5605 GND.n660 240.244
R4659 GND.n5609 GND.n660 240.244
R4660 GND.n5609 GND.n656 240.244
R4661 GND.n5615 GND.n656 240.244
R4662 GND.n5615 GND.n654 240.244
R4663 GND.n5619 GND.n654 240.244
R4664 GND.n5619 GND.n650 240.244
R4665 GND.n5625 GND.n650 240.244
R4666 GND.n5625 GND.n648 240.244
R4667 GND.n5629 GND.n648 240.244
R4668 GND.n5629 GND.n644 240.244
R4669 GND.n5635 GND.n644 240.244
R4670 GND.n5635 GND.n642 240.244
R4671 GND.n5639 GND.n642 240.244
R4672 GND.n5639 GND.n638 240.244
R4673 GND.n5645 GND.n638 240.244
R4674 GND.n5645 GND.n636 240.244
R4675 GND.n5649 GND.n636 240.244
R4676 GND.n5649 GND.n632 240.244
R4677 GND.n5655 GND.n632 240.244
R4678 GND.n5655 GND.n630 240.244
R4679 GND.n5659 GND.n630 240.244
R4680 GND.n5659 GND.n626 240.244
R4681 GND.n5665 GND.n626 240.244
R4682 GND.n5665 GND.n624 240.244
R4683 GND.n5669 GND.n624 240.244
R4684 GND.n5669 GND.n620 240.244
R4685 GND.n5675 GND.n620 240.244
R4686 GND.n5675 GND.n618 240.244
R4687 GND.n5679 GND.n618 240.244
R4688 GND.n5679 GND.n614 240.244
R4689 GND.n5685 GND.n614 240.244
R4690 GND.n5685 GND.n612 240.244
R4691 GND.n5689 GND.n612 240.244
R4692 GND.n5689 GND.n608 240.244
R4693 GND.n5695 GND.n608 240.244
R4694 GND.n5695 GND.n606 240.244
R4695 GND.n5699 GND.n606 240.244
R4696 GND.n5699 GND.n602 240.244
R4697 GND.n5705 GND.n602 240.244
R4698 GND.n5705 GND.n600 240.244
R4699 GND.n5709 GND.n600 240.244
R4700 GND.n5709 GND.n596 240.244
R4701 GND.n5715 GND.n596 240.244
R4702 GND.n5715 GND.n594 240.244
R4703 GND.n5719 GND.n594 240.244
R4704 GND.n5719 GND.n590 240.244
R4705 GND.n5725 GND.n590 240.244
R4706 GND.n5725 GND.n588 240.244
R4707 GND.n5729 GND.n588 240.244
R4708 GND.n5729 GND.n584 240.244
R4709 GND.n5735 GND.n584 240.244
R4710 GND.n5735 GND.n582 240.244
R4711 GND.n5739 GND.n582 240.244
R4712 GND.n5739 GND.n578 240.244
R4713 GND.n5745 GND.n578 240.244
R4714 GND.n5745 GND.n576 240.244
R4715 GND.n5749 GND.n576 240.244
R4716 GND.n5749 GND.n572 240.244
R4717 GND.n5755 GND.n572 240.244
R4718 GND.n5755 GND.n570 240.244
R4719 GND.n5759 GND.n570 240.244
R4720 GND.n5759 GND.n566 240.244
R4721 GND.n5765 GND.n566 240.244
R4722 GND.n5765 GND.n564 240.244
R4723 GND.n5769 GND.n564 240.244
R4724 GND.n5769 GND.n560 240.244
R4725 GND.n5775 GND.n560 240.244
R4726 GND.n5775 GND.n558 240.244
R4727 GND.n5779 GND.n558 240.244
R4728 GND.n5779 GND.n554 240.244
R4729 GND.n5785 GND.n554 240.244
R4730 GND.n5785 GND.n552 240.244
R4731 GND.n5789 GND.n552 240.244
R4732 GND.n5789 GND.n548 240.244
R4733 GND.n5795 GND.n548 240.244
R4734 GND.n5795 GND.n546 240.244
R4735 GND.n5799 GND.n546 240.244
R4736 GND.n5799 GND.n542 240.244
R4737 GND.n5805 GND.n542 240.244
R4738 GND.n5805 GND.n540 240.244
R4739 GND.n5809 GND.n540 240.244
R4740 GND.n5809 GND.n536 240.244
R4741 GND.n5815 GND.n536 240.244
R4742 GND.n5815 GND.n534 240.244
R4743 GND.n5819 GND.n534 240.244
R4744 GND.n5819 GND.n530 240.244
R4745 GND.n5825 GND.n530 240.244
R4746 GND.n5825 GND.n528 240.244
R4747 GND.n5829 GND.n528 240.244
R4748 GND.n5829 GND.n524 240.244
R4749 GND.n5835 GND.n524 240.244
R4750 GND.n5835 GND.n522 240.244
R4751 GND.n5839 GND.n522 240.244
R4752 GND.n5839 GND.n518 240.244
R4753 GND.n5845 GND.n518 240.244
R4754 GND.n5845 GND.n516 240.244
R4755 GND.n5849 GND.n516 240.244
R4756 GND.n5849 GND.n512 240.244
R4757 GND.n5855 GND.n512 240.244
R4758 GND.n5855 GND.n510 240.244
R4759 GND.n5859 GND.n510 240.244
R4760 GND.n5859 GND.n506 240.244
R4761 GND.n5865 GND.n506 240.244
R4762 GND.n5865 GND.n504 240.244
R4763 GND.n5869 GND.n504 240.244
R4764 GND.n5869 GND.n500 240.244
R4765 GND.n5875 GND.n500 240.244
R4766 GND.n5875 GND.n498 240.244
R4767 GND.n5879 GND.n498 240.244
R4768 GND.n5879 GND.n494 240.244
R4769 GND.n5885 GND.n494 240.244
R4770 GND.n5885 GND.n492 240.244
R4771 GND.n5889 GND.n492 240.244
R4772 GND.n5889 GND.n488 240.244
R4773 GND.n5895 GND.n488 240.244
R4774 GND.n5895 GND.n486 240.244
R4775 GND.n5899 GND.n486 240.244
R4776 GND.n5899 GND.n482 240.244
R4777 GND.n5905 GND.n482 240.244
R4778 GND.n5905 GND.n480 240.244
R4779 GND.n5909 GND.n480 240.244
R4780 GND.n5909 GND.n476 240.244
R4781 GND.n5915 GND.n476 240.244
R4782 GND.n5915 GND.n474 240.244
R4783 GND.n5919 GND.n474 240.244
R4784 GND.n5919 GND.n470 240.244
R4785 GND.n5925 GND.n470 240.244
R4786 GND.n5925 GND.n468 240.244
R4787 GND.n5929 GND.n468 240.244
R4788 GND.n5929 GND.n464 240.244
R4789 GND.n5935 GND.n464 240.244
R4790 GND.n5935 GND.n462 240.244
R4791 GND.n5939 GND.n462 240.244
R4792 GND.n5939 GND.n458 240.244
R4793 GND.n5945 GND.n458 240.244
R4794 GND.n5945 GND.n456 240.244
R4795 GND.n5949 GND.n456 240.244
R4796 GND.n5949 GND.n452 240.244
R4797 GND.n5955 GND.n452 240.244
R4798 GND.n5955 GND.n450 240.244
R4799 GND.n5959 GND.n450 240.244
R4800 GND.n5959 GND.n446 240.244
R4801 GND.n5965 GND.n446 240.244
R4802 GND.n5965 GND.n444 240.244
R4803 GND.n5969 GND.n444 240.244
R4804 GND.n5969 GND.n440 240.244
R4805 GND.n5975 GND.n440 240.244
R4806 GND.n5975 GND.n438 240.244
R4807 GND.n5979 GND.n438 240.244
R4808 GND.n5979 GND.n434 240.244
R4809 GND.n5985 GND.n434 240.244
R4810 GND.n5985 GND.n432 240.244
R4811 GND.n5989 GND.n432 240.244
R4812 GND.n5989 GND.n428 240.244
R4813 GND.n5995 GND.n428 240.244
R4814 GND.n5995 GND.n426 240.244
R4815 GND.n5999 GND.n426 240.244
R4816 GND.n5999 GND.n422 240.244
R4817 GND.n6005 GND.n422 240.244
R4818 GND.n6005 GND.n420 240.244
R4819 GND.n6009 GND.n420 240.244
R4820 GND.n6009 GND.n416 240.244
R4821 GND.n6015 GND.n416 240.244
R4822 GND.n6015 GND.n414 240.244
R4823 GND.n6019 GND.n414 240.244
R4824 GND.n6019 GND.n410 240.244
R4825 GND.n6025 GND.n410 240.244
R4826 GND.n6025 GND.n408 240.244
R4827 GND.n6029 GND.n408 240.244
R4828 GND.n6029 GND.n404 240.244
R4829 GND.n6035 GND.n404 240.244
R4830 GND.n6035 GND.n402 240.244
R4831 GND.n6039 GND.n402 240.244
R4832 GND.n6039 GND.n398 240.244
R4833 GND.n6045 GND.n398 240.244
R4834 GND.n6045 GND.n396 240.244
R4835 GND.n6049 GND.n396 240.244
R4836 GND.n6049 GND.n392 240.244
R4837 GND.n6055 GND.n392 240.244
R4838 GND.n6055 GND.n390 240.244
R4839 GND.n6059 GND.n390 240.244
R4840 GND.n6059 GND.n386 240.244
R4841 GND.n6065 GND.n386 240.244
R4842 GND.n6065 GND.n384 240.244
R4843 GND.n6069 GND.n384 240.244
R4844 GND.n6069 GND.n380 240.244
R4845 GND.n6075 GND.n380 240.244
R4846 GND.n6075 GND.n378 240.244
R4847 GND.n6079 GND.n378 240.244
R4848 GND.n6079 GND.n374 240.244
R4849 GND.n6085 GND.n374 240.244
R4850 GND.n6085 GND.n372 240.244
R4851 GND.n6089 GND.n372 240.244
R4852 GND.n6089 GND.n368 240.244
R4853 GND.n6095 GND.n368 240.244
R4854 GND.n6095 GND.n366 240.244
R4855 GND.n6099 GND.n366 240.244
R4856 GND.n6099 GND.n362 240.244
R4857 GND.n6105 GND.n362 240.244
R4858 GND.n6105 GND.n360 240.244
R4859 GND.n6109 GND.n360 240.244
R4860 GND.n6109 GND.n356 240.244
R4861 GND.n6115 GND.n356 240.244
R4862 GND.n6115 GND.n354 240.244
R4863 GND.n6119 GND.n354 240.244
R4864 GND.n6119 GND.n350 240.244
R4865 GND.n6125 GND.n350 240.244
R4866 GND.n6125 GND.n348 240.244
R4867 GND.n6129 GND.n348 240.244
R4868 GND.n6129 GND.n344 240.244
R4869 GND.n6135 GND.n344 240.244
R4870 GND.n6135 GND.n342 240.244
R4871 GND.n6139 GND.n342 240.244
R4872 GND.n6139 GND.n338 240.244
R4873 GND.n6145 GND.n338 240.244
R4874 GND.n6145 GND.n336 240.244
R4875 GND.n6149 GND.n336 240.244
R4876 GND.n6149 GND.n332 240.244
R4877 GND.n6155 GND.n332 240.244
R4878 GND.n6155 GND.n330 240.244
R4879 GND.n6159 GND.n330 240.244
R4880 GND.n6159 GND.n326 240.244
R4881 GND.n6165 GND.n326 240.244
R4882 GND.n6165 GND.n324 240.244
R4883 GND.n6169 GND.n324 240.244
R4884 GND.n6169 GND.n320 240.244
R4885 GND.n6175 GND.n320 240.244
R4886 GND.n6175 GND.n318 240.244
R4887 GND.n6179 GND.n318 240.244
R4888 GND.n6179 GND.n314 240.244
R4889 GND.n6185 GND.n314 240.244
R4890 GND.n6185 GND.n312 240.244
R4891 GND.n6189 GND.n312 240.244
R4892 GND.n6195 GND.n308 240.244
R4893 GND.n6195 GND.n306 240.244
R4894 GND.n6199 GND.n306 240.244
R4895 GND.n6199 GND.n302 240.244
R4896 GND.n6205 GND.n302 240.244
R4897 GND.n6205 GND.n300 240.244
R4898 GND.n6209 GND.n300 240.244
R4899 GND.n6209 GND.n296 240.244
R4900 GND.n6215 GND.n296 240.244
R4901 GND.n6215 GND.n294 240.244
R4902 GND.n6219 GND.n294 240.244
R4903 GND.n6219 GND.n290 240.244
R4904 GND.n6225 GND.n290 240.244
R4905 GND.n6225 GND.n288 240.244
R4906 GND.n6229 GND.n288 240.244
R4907 GND.n6229 GND.n284 240.244
R4908 GND.n6235 GND.n284 240.244
R4909 GND.n6235 GND.n282 240.244
R4910 GND.n6239 GND.n282 240.244
R4911 GND.n6239 GND.n278 240.244
R4912 GND.n6245 GND.n278 240.244
R4913 GND.n6245 GND.n276 240.244
R4914 GND.n6249 GND.n276 240.244
R4915 GND.n6249 GND.n272 240.244
R4916 GND.n6255 GND.n272 240.244
R4917 GND.n6255 GND.n270 240.244
R4918 GND.n6259 GND.n270 240.244
R4919 GND.n6259 GND.n266 240.244
R4920 GND.n6265 GND.n266 240.244
R4921 GND.n6265 GND.n264 240.244
R4922 GND.n6269 GND.n264 240.244
R4923 GND.n6269 GND.n260 240.244
R4924 GND.n6275 GND.n260 240.244
R4925 GND.n6275 GND.n258 240.244
R4926 GND.n6279 GND.n258 240.244
R4927 GND.n6279 GND.n254 240.244
R4928 GND.n6285 GND.n254 240.244
R4929 GND.n6285 GND.n252 240.244
R4930 GND.n6289 GND.n252 240.244
R4931 GND.n6289 GND.n248 240.244
R4932 GND.n6295 GND.n248 240.244
R4933 GND.n6295 GND.n246 240.244
R4934 GND.n6299 GND.n246 240.244
R4935 GND.n6299 GND.n242 240.244
R4936 GND.n6305 GND.n242 240.244
R4937 GND.n6305 GND.n240 240.244
R4938 GND.n6309 GND.n240 240.244
R4939 GND.n6309 GND.n236 240.244
R4940 GND.n6315 GND.n236 240.244
R4941 GND.n6315 GND.n234 240.244
R4942 GND.n6319 GND.n234 240.244
R4943 GND.n6319 GND.n230 240.244
R4944 GND.n6325 GND.n230 240.244
R4945 GND.n6325 GND.n228 240.244
R4946 GND.n6329 GND.n228 240.244
R4947 GND.n6329 GND.n224 240.244
R4948 GND.n6336 GND.n224 240.244
R4949 GND.n6336 GND.n222 240.244
R4950 GND.n6340 GND.n222 240.244
R4951 GND.n6340 GND.n218 240.244
R4952 GND.n5335 GND.n868 240.244
R4953 GND.n5335 GND.n870 240.244
R4954 GND.n5331 GND.n870 240.244
R4955 GND.n5331 GND.n877 240.244
R4956 GND.n5327 GND.n877 240.244
R4957 GND.n5327 GND.n879 240.244
R4958 GND.n5323 GND.n879 240.244
R4959 GND.n5323 GND.n885 240.244
R4960 GND.n5319 GND.n885 240.244
R4961 GND.n5319 GND.n887 240.244
R4962 GND.n5315 GND.n887 240.244
R4963 GND.n5315 GND.n893 240.244
R4964 GND.n5311 GND.n893 240.244
R4965 GND.n5311 GND.n895 240.244
R4966 GND.n5307 GND.n895 240.244
R4967 GND.n5307 GND.n901 240.244
R4968 GND.n5303 GND.n901 240.244
R4969 GND.n5303 GND.n903 240.244
R4970 GND.n5299 GND.n903 240.244
R4971 GND.n5299 GND.n909 240.244
R4972 GND.n5295 GND.n909 240.244
R4973 GND.n5295 GND.n911 240.244
R4974 GND.n5291 GND.n911 240.244
R4975 GND.n5291 GND.n917 240.244
R4976 GND.n5287 GND.n917 240.244
R4977 GND.n5287 GND.n919 240.244
R4978 GND.n5283 GND.n919 240.244
R4979 GND.n5283 GND.n925 240.244
R4980 GND.n5279 GND.n925 240.244
R4981 GND.n5279 GND.n927 240.244
R4982 GND.n5275 GND.n927 240.244
R4983 GND.n5275 GND.n933 240.244
R4984 GND.n5271 GND.n933 240.244
R4985 GND.n5271 GND.n935 240.244
R4986 GND.n5267 GND.n935 240.244
R4987 GND.n5267 GND.n941 240.244
R4988 GND.n1023 GND.n941 240.244
R4989 GND.n1023 GND.n1019 240.244
R4990 GND.n5186 GND.n1019 240.244
R4991 GND.n5186 GND.n1020 240.244
R4992 GND.n5182 GND.n1020 240.244
R4993 GND.n5182 GND.n1031 240.244
R4994 GND.n3120 GND.n1031 240.244
R4995 GND.n3120 GND.n3116 240.244
R4996 GND.n3137 GND.n3116 240.244
R4997 GND.n3137 GND.n3117 240.244
R4998 GND.n3133 GND.n3117 240.244
R4999 GND.n3133 GND.n3132 240.244
R5000 GND.n3132 GND.n3131 240.244
R5001 GND.n3131 GND.n3017 240.244
R5002 GND.n3182 GND.n3017 240.244
R5003 GND.n3182 GND.n3012 240.244
R5004 GND.n3190 GND.n3012 240.244
R5005 GND.n3190 GND.n3013 240.244
R5006 GND.n3013 GND.n2989 240.244
R5007 GND.n3217 GND.n2989 240.244
R5008 GND.n3217 GND.n2984 240.244
R5009 GND.n3226 GND.n2984 240.244
R5010 GND.n3226 GND.n2985 240.244
R5011 GND.n2985 GND.n2958 240.244
R5012 GND.n3279 GND.n2958 240.244
R5013 GND.n3279 GND.n2959 240.244
R5014 GND.n3274 GND.n2959 240.244
R5015 GND.n3274 GND.n2962 240.244
R5016 GND.n3252 GND.n2962 240.244
R5017 GND.n3261 GND.n3252 240.244
R5018 GND.n3261 GND.n3253 240.244
R5019 GND.n3253 GND.n2927 240.244
R5020 GND.n3303 GND.n2927 240.244
R5021 GND.n3304 GND.n3303 240.244
R5022 GND.n3304 GND.n2922 240.244
R5023 GND.n3367 GND.n2922 240.244
R5024 GND.n3367 GND.n2923 240.244
R5025 GND.n3363 GND.n2923 240.244
R5026 GND.n3363 GND.n3362 240.244
R5027 GND.n3362 GND.n3361 240.244
R5028 GND.n3361 GND.n3312 240.244
R5029 GND.n3357 GND.n3312 240.244
R5030 GND.n3357 GND.n3353 240.244
R5031 GND.n3353 GND.n3352 240.244
R5032 GND.n3352 GND.n3318 240.244
R5033 GND.n3348 GND.n3318 240.244
R5034 GND.n3348 GND.n3347 240.244
R5035 GND.n3347 GND.n3346 240.244
R5036 GND.n3346 GND.n3324 240.244
R5037 GND.n3342 GND.n3324 240.244
R5038 GND.n3342 GND.n3341 240.244
R5039 GND.n3341 GND.n3340 240.244
R5040 GND.n3340 GND.n3330 240.244
R5041 GND.n3336 GND.n3330 240.244
R5042 GND.n3336 GND.n1292 240.244
R5043 GND.n4977 GND.n1292 240.244
R5044 GND.n4977 GND.n1293 240.244
R5045 GND.n4973 GND.n1293 240.244
R5046 GND.n4973 GND.n4972 240.244
R5047 GND.n4972 GND.n4971 240.244
R5048 GND.n4971 GND.n1299 240.244
R5049 GND.n1322 GND.n1299 240.244
R5050 GND.n1322 GND.n1315 240.244
R5051 GND.n4959 GND.n1315 240.244
R5052 GND.n4959 GND.n1316 240.244
R5053 GND.n4955 GND.n1316 240.244
R5054 GND.n4955 GND.n1330 240.244
R5055 GND.n1348 GND.n1330 240.244
R5056 GND.n4945 GND.n1348 240.244
R5057 GND.n4945 GND.n1349 240.244
R5058 GND.n4941 GND.n1349 240.244
R5059 GND.n4941 GND.n1357 240.244
R5060 GND.n1375 GND.n1357 240.244
R5061 GND.n4931 GND.n1375 240.244
R5062 GND.n4931 GND.n1376 240.244
R5063 GND.n4927 GND.n1376 240.244
R5064 GND.n4927 GND.n1384 240.244
R5065 GND.n1402 GND.n1384 240.244
R5066 GND.n4917 GND.n1402 240.244
R5067 GND.n4917 GND.n1403 240.244
R5068 GND.n4913 GND.n1403 240.244
R5069 GND.n4913 GND.n1411 240.244
R5070 GND.n3685 GND.n1411 240.244
R5071 GND.n3686 GND.n3685 240.244
R5072 GND.n3687 GND.n3686 240.244
R5073 GND.n3687 GND.n3677 240.244
R5074 GND.n3701 GND.n3677 240.244
R5075 GND.n3701 GND.n3678 240.244
R5076 GND.n3697 GND.n3678 240.244
R5077 GND.n3697 GND.n2691 240.244
R5078 GND.n3745 GND.n2691 240.244
R5079 GND.n3746 GND.n3745 240.244
R5080 GND.n3747 GND.n3746 240.244
R5081 GND.n3747 GND.n2687 240.244
R5082 GND.n3753 GND.n2687 240.244
R5083 GND.n3753 GND.n2681 240.244
R5084 GND.n3772 GND.n2681 240.244
R5085 GND.n3772 GND.n2676 240.244
R5086 GND.n3787 GND.n2676 240.244
R5087 GND.n3787 GND.n2677 240.244
R5088 GND.n3783 GND.n2677 240.244
R5089 GND.n3783 GND.n3782 240.244
R5090 GND.n3782 GND.n1527 240.244
R5091 GND.n4833 GND.n1527 240.244
R5092 GND.n4833 GND.n1528 240.244
R5093 GND.n4829 GND.n1528 240.244
R5094 GND.n4829 GND.n1534 240.244
R5095 GND.n1578 GND.n1534 240.244
R5096 GND.n1579 GND.n1578 240.244
R5097 GND.n1579 GND.n1572 240.244
R5098 GND.n4806 GND.n1572 240.244
R5099 GND.n4806 GND.n1573 240.244
R5100 GND.n4802 GND.n1573 240.244
R5101 GND.n4802 GND.n1587 240.244
R5102 GND.n1620 GND.n1587 240.244
R5103 GND.n1620 GND.n1616 240.244
R5104 GND.n4785 GND.n1616 240.244
R5105 GND.n4785 GND.n1617 240.244
R5106 GND.n4781 GND.n1617 240.244
R5107 GND.n4781 GND.n1628 240.244
R5108 GND.n1664 GND.n1628 240.244
R5109 GND.n1664 GND.n1660 240.244
R5110 GND.n4764 GND.n1660 240.244
R5111 GND.n4764 GND.n1661 240.244
R5112 GND.n4760 GND.n1661 240.244
R5113 GND.n4760 GND.n1672 240.244
R5114 GND.n1715 GND.n1672 240.244
R5115 GND.n1716 GND.n1715 240.244
R5116 GND.n1716 GND.n1709 240.244
R5117 GND.n4737 GND.n1709 240.244
R5118 GND.n4737 GND.n1710 240.244
R5119 GND.n4733 GND.n1710 240.244
R5120 GND.n4733 GND.n1724 240.244
R5121 GND.n2307 GND.n1724 240.244
R5122 GND.n2308 GND.n2307 240.244
R5123 GND.n2308 GND.n2302 240.244
R5124 GND.n2315 GND.n2302 240.244
R5125 GND.n2315 GND.n1758 240.244
R5126 GND.n4709 GND.n1758 240.244
R5127 GND.n4709 GND.n1759 240.244
R5128 GND.n4705 GND.n1759 240.244
R5129 GND.n4705 GND.n1765 240.244
R5130 GND.n1782 GND.n1765 240.244
R5131 GND.n4695 GND.n1782 240.244
R5132 GND.n4695 GND.n1783 240.244
R5133 GND.n4691 GND.n1783 240.244
R5134 GND.n4691 GND.n1791 240.244
R5135 GND.n1808 GND.n1791 240.244
R5136 GND.n4681 GND.n1808 240.244
R5137 GND.n4681 GND.n1809 240.244
R5138 GND.n4677 GND.n1809 240.244
R5139 GND.n4677 GND.n1817 240.244
R5140 GND.n1835 GND.n1817 240.244
R5141 GND.n4667 GND.n1835 240.244
R5142 GND.n4667 GND.n1836 240.244
R5143 GND.n4663 GND.n1836 240.244
R5144 GND.n4663 GND.n1844 240.244
R5145 GND.n1861 GND.n1844 240.244
R5146 GND.n4653 GND.n1861 240.244
R5147 GND.n4653 GND.n1862 240.244
R5148 GND.n4649 GND.n1862 240.244
R5149 GND.n4649 GND.n1870 240.244
R5150 GND.n4645 GND.n1870 240.244
R5151 GND.n4645 GND.n1873 240.244
R5152 GND.n4641 GND.n1873 240.244
R5153 GND.n4641 GND.n1879 240.244
R5154 GND.n4231 GND.n1879 240.244
R5155 GND.n4231 GND.n4227 240.244
R5156 GND.n4278 GND.n4227 240.244
R5157 GND.n4278 GND.n4228 240.244
R5158 GND.n4274 GND.n4228 240.244
R5159 GND.n4274 GND.n4273 240.244
R5160 GND.n4273 GND.n4272 240.244
R5161 GND.n4272 GND.n4239 240.244
R5162 GND.n4268 GND.n4239 240.244
R5163 GND.n4268 GND.n4267 240.244
R5164 GND.n4267 GND.n4266 240.244
R5165 GND.n4266 GND.n4245 240.244
R5166 GND.n4262 GND.n4245 240.244
R5167 GND.n4262 GND.n4261 240.244
R5168 GND.n4261 GND.n4260 240.244
R5169 GND.n4260 GND.n4251 240.244
R5170 GND.n4256 GND.n4251 240.244
R5171 GND.n4256 GND.n2145 240.244
R5172 GND.n4432 GND.n2145 240.244
R5173 GND.n4432 GND.n2146 240.244
R5174 GND.n2165 GND.n2146 240.244
R5175 GND.n2168 GND.n2165 240.244
R5176 GND.n4418 GND.n2168 240.244
R5177 GND.n4418 GND.n4415 240.244
R5178 GND.n4415 GND.n2169 240.244
R5179 GND.n4396 GND.n2169 240.244
R5180 GND.n4397 GND.n4396 240.244
R5181 GND.n4400 GND.n4397 240.244
R5182 GND.n4400 GND.n2133 240.244
R5183 GND.n4440 GND.n2133 240.244
R5184 GND.n4440 GND.n2134 240.244
R5185 GND.n2134 GND.n2116 240.244
R5186 GND.n4458 GND.n2116 240.244
R5187 GND.n4458 GND.n2111 240.244
R5188 GND.n4466 GND.n2111 240.244
R5189 GND.n4466 GND.n2112 240.244
R5190 GND.n2112 GND.n2093 240.244
R5191 GND.n4484 GND.n2093 240.244
R5192 GND.n4484 GND.n2088 240.244
R5193 GND.n4492 GND.n2088 240.244
R5194 GND.n4492 GND.n2089 240.244
R5195 GND.n2089 GND.n2074 240.244
R5196 GND.n4513 GND.n2074 240.244
R5197 GND.n4513 GND.n2069 240.244
R5198 GND.n4537 GND.n2069 240.244
R5199 GND.n4537 GND.n2070 240.244
R5200 GND.n4533 GND.n2070 240.244
R5201 GND.n4533 GND.n4532 240.244
R5202 GND.n4532 GND.n4531 240.244
R5203 GND.n4531 GND.n4521 240.244
R5204 GND.n4527 GND.n4521 240.244
R5205 GND.n4527 GND.n145 240.244
R5206 GND.n6418 GND.n145 240.244
R5207 GND.n6418 GND.n146 240.244
R5208 GND.n6414 GND.n146 240.244
R5209 GND.n6414 GND.n152 240.244
R5210 GND.n6410 GND.n152 240.244
R5211 GND.n6410 GND.n154 240.244
R5212 GND.n6406 GND.n154 240.244
R5213 GND.n6406 GND.n160 240.244
R5214 GND.n6402 GND.n160 240.244
R5215 GND.n6402 GND.n162 240.244
R5216 GND.n6398 GND.n162 240.244
R5217 GND.n6398 GND.n168 240.244
R5218 GND.n6394 GND.n168 240.244
R5219 GND.n6394 GND.n170 240.244
R5220 GND.n6390 GND.n170 240.244
R5221 GND.n6390 GND.n176 240.244
R5222 GND.n6386 GND.n176 240.244
R5223 GND.n6386 GND.n178 240.244
R5224 GND.n6382 GND.n178 240.244
R5225 GND.n6382 GND.n184 240.244
R5226 GND.n6378 GND.n184 240.244
R5227 GND.n6378 GND.n186 240.244
R5228 GND.n6374 GND.n186 240.244
R5229 GND.n6374 GND.n192 240.244
R5230 GND.n6370 GND.n192 240.244
R5231 GND.n6370 GND.n194 240.244
R5232 GND.n6366 GND.n194 240.244
R5233 GND.n6366 GND.n200 240.244
R5234 GND.n6362 GND.n200 240.244
R5235 GND.n6362 GND.n202 240.244
R5236 GND.n6358 GND.n202 240.244
R5237 GND.n6358 GND.n208 240.244
R5238 GND.n6354 GND.n208 240.244
R5239 GND.n6354 GND.n210 240.244
R5240 GND.n6350 GND.n210 240.244
R5241 GND.n6350 GND.n216 240.244
R5242 GND.n6346 GND.n216 240.244
R5243 GND.n5459 GND.n750 240.244
R5244 GND.n5455 GND.n750 240.244
R5245 GND.n5455 GND.n752 240.244
R5246 GND.n5451 GND.n752 240.244
R5247 GND.n5451 GND.n757 240.244
R5248 GND.n5447 GND.n757 240.244
R5249 GND.n5447 GND.n759 240.244
R5250 GND.n5443 GND.n759 240.244
R5251 GND.n5443 GND.n765 240.244
R5252 GND.n5439 GND.n765 240.244
R5253 GND.n5439 GND.n767 240.244
R5254 GND.n5435 GND.n767 240.244
R5255 GND.n5435 GND.n773 240.244
R5256 GND.n5431 GND.n773 240.244
R5257 GND.n5431 GND.n775 240.244
R5258 GND.n5427 GND.n775 240.244
R5259 GND.n5427 GND.n781 240.244
R5260 GND.n5423 GND.n781 240.244
R5261 GND.n5423 GND.n783 240.244
R5262 GND.n5419 GND.n783 240.244
R5263 GND.n5419 GND.n789 240.244
R5264 GND.n5415 GND.n789 240.244
R5265 GND.n5415 GND.n791 240.244
R5266 GND.n5411 GND.n791 240.244
R5267 GND.n5411 GND.n797 240.244
R5268 GND.n5407 GND.n797 240.244
R5269 GND.n5407 GND.n799 240.244
R5270 GND.n5403 GND.n799 240.244
R5271 GND.n5403 GND.n805 240.244
R5272 GND.n5399 GND.n805 240.244
R5273 GND.n5399 GND.n807 240.244
R5274 GND.n5395 GND.n807 240.244
R5275 GND.n5395 GND.n813 240.244
R5276 GND.n5391 GND.n813 240.244
R5277 GND.n5391 GND.n815 240.244
R5278 GND.n5387 GND.n815 240.244
R5279 GND.n5387 GND.n821 240.244
R5280 GND.n5383 GND.n821 240.244
R5281 GND.n5383 GND.n823 240.244
R5282 GND.n5379 GND.n823 240.244
R5283 GND.n5379 GND.n829 240.244
R5284 GND.n5375 GND.n829 240.244
R5285 GND.n5375 GND.n831 240.244
R5286 GND.n5371 GND.n831 240.244
R5287 GND.n5371 GND.n837 240.244
R5288 GND.n5367 GND.n837 240.244
R5289 GND.n5367 GND.n839 240.244
R5290 GND.n5363 GND.n839 240.244
R5291 GND.n5363 GND.n845 240.244
R5292 GND.n5359 GND.n845 240.244
R5293 GND.n5359 GND.n847 240.244
R5294 GND.n5355 GND.n847 240.244
R5295 GND.n5355 GND.n853 240.244
R5296 GND.n5351 GND.n853 240.244
R5297 GND.n5351 GND.n855 240.244
R5298 GND.n5347 GND.n855 240.244
R5299 GND.n5347 GND.n861 240.244
R5300 GND.n5343 GND.n861 240.244
R5301 GND.n5343 GND.n863 240.244
R5302 GND.n5339 GND.n863 240.244
R5303 GND.n2537 GND.n2536 240.244
R5304 GND.n2534 GND.n2441 240.244
R5305 GND.n2446 GND.n2445 240.244
R5306 GND.n2455 GND.n2454 240.244
R5307 GND.n2458 GND.n2457 240.244
R5308 GND.n2470 GND.n2469 240.244
R5309 GND.n2481 GND.n2472 240.244
R5310 GND.n2500 GND.n2483 240.244
R5311 GND.n1896 GND.n1884 240.244
R5312 GND.n4632 GND.n1896 240.244
R5313 GND.n4632 GND.n1897 240.244
R5314 GND.n2236 GND.n1897 240.244
R5315 GND.n4290 GND.n2236 240.244
R5316 GND.n4294 GND.n4290 240.244
R5317 GND.n4294 GND.n4293 240.244
R5318 GND.n4293 GND.n2224 240.244
R5319 GND.n2224 GND.n2214 240.244
R5320 GND.n4315 GND.n2214 240.244
R5321 GND.n4319 GND.n4315 240.244
R5322 GND.n4319 GND.n4317 240.244
R5323 GND.n4317 GND.n2203 240.244
R5324 GND.n2203 GND.n2191 240.244
R5325 GND.n4340 GND.n2191 240.244
R5326 GND.n4344 GND.n4340 240.244
R5327 GND.n4344 GND.n4343 240.244
R5328 GND.n4343 GND.n2182 240.244
R5329 GND.n2182 GND.n2181 240.244
R5330 GND.n2181 GND.n2150 240.244
R5331 GND.n2160 GND.n2150 240.244
R5332 GND.n4422 GND.n2160 240.244
R5333 GND.n4422 GND.n4421 240.244
R5334 GND.n4421 GND.n2161 240.244
R5335 GND.n4373 GND.n2161 240.244
R5336 GND.n4383 GND.n4373 240.244
R5337 GND.n4405 GND.n4383 240.244
R5338 GND.n4405 GND.n4403 240.244
R5339 GND.n4403 GND.n4384 240.244
R5340 GND.n4384 GND.n2130 240.244
R5341 GND.n4443 GND.n2130 240.244
R5342 GND.n4445 GND.n4443 240.244
R5343 GND.n4445 GND.n4444 240.244
R5344 GND.n4444 GND.n2121 240.244
R5345 GND.n2121 GND.n2109 240.244
R5346 GND.n4469 GND.n2109 240.244
R5347 GND.n4471 GND.n4469 240.244
R5348 GND.n4471 GND.n4470 240.244
R5349 GND.n4470 GND.n2097 240.244
R5350 GND.n2097 GND.n2086 240.244
R5351 GND.n4497 GND.n2086 240.244
R5352 GND.n4500 GND.n4497 240.244
R5353 GND.n4500 GND.n4499 240.244
R5354 GND.n4499 GND.n2077 240.244
R5355 GND.n2077 GND.n2065 240.244
R5356 GND.n4540 GND.n2065 240.244
R5357 GND.n4542 GND.n4540 240.244
R5358 GND.n4542 GND.n2054 240.244
R5359 GND.n4552 GND.n2054 240.244
R5360 GND.n4553 GND.n4552 240.244
R5361 GND.n4553 GND.n82 240.244
R5362 GND.n2001 GND.n2000 240.244
R5363 GND.n2005 GND.n2004 240.244
R5364 GND.n2007 GND.n2006 240.244
R5365 GND.n2011 GND.n2010 240.244
R5366 GND.n2013 GND.n2012 240.244
R5367 GND.n2017 GND.n2016 240.244
R5368 GND.n2019 GND.n2018 240.244
R5369 GND.n2022 GND.n78 240.244
R5370 GND.n2246 GND.n1882 240.244
R5371 GND.n2246 GND.n1894 240.244
R5372 GND.n4281 GND.n1894 240.244
R5373 GND.n4281 GND.n2239 240.244
R5374 GND.n4288 GND.n2239 240.244
R5375 GND.n4288 GND.n2234 240.244
R5376 GND.n2234 GND.n2221 240.244
R5377 GND.n4306 GND.n2221 240.244
R5378 GND.n4306 GND.n2216 240.244
R5379 GND.n4313 GND.n2216 240.244
R5380 GND.n4313 GND.n2212 240.244
R5381 GND.n2212 GND.n2199 240.244
R5382 GND.n4331 GND.n2199 240.244
R5383 GND.n4331 GND.n2194 240.244
R5384 GND.n4338 GND.n2194 240.244
R5385 GND.n4338 GND.n2189 240.244
R5386 GND.n2189 GND.n2176 240.244
R5387 GND.n4355 GND.n2176 240.244
R5388 GND.n4355 GND.n2177 240.244
R5389 GND.n2177 GND.n2148 240.244
R5390 GND.n4363 GND.n2148 240.244
R5391 GND.n4363 GND.n2158 240.244
R5392 GND.n2163 GND.n2158 240.244
R5393 GND.n4370 GND.n2163 240.244
R5394 GND.n4371 GND.n4370 240.244
R5395 GND.n4371 GND.n47 240.244
R5396 GND.n48 GND.n47 240.244
R5397 GND.n49 GND.n48 240.244
R5398 GND.n4386 GND.n49 240.244
R5399 GND.n4386 GND.n52 240.244
R5400 GND.n53 GND.n52 240.244
R5401 GND.n54 GND.n53 240.244
R5402 GND.n2118 GND.n54 240.244
R5403 GND.n2118 GND.n57 240.244
R5404 GND.n58 GND.n57 240.244
R5405 GND.n59 GND.n58 240.244
R5406 GND.n2106 GND.n59 240.244
R5407 GND.n2106 GND.n62 240.244
R5408 GND.n63 GND.n62 240.244
R5409 GND.n64 GND.n63 240.244
R5410 GND.n4495 GND.n64 240.244
R5411 GND.n4495 GND.n67 240.244
R5412 GND.n68 GND.n67 240.244
R5413 GND.n69 GND.n68 240.244
R5414 GND.n2067 GND.n69 240.244
R5415 GND.n2067 GND.n72 240.244
R5416 GND.n73 GND.n72 240.244
R5417 GND.n74 GND.n73 240.244
R5418 GND.n2056 GND.n74 240.244
R5419 GND.n2056 GND.n77 240.244
R5420 GND.n6503 GND.n77 240.244
R5421 GND.n3567 GND.n3566 228.118
R5422 GND.n2323 GND.n2322 228.118
R5423 GND.n2578 GND.n2355 199.319
R5424 GND.n4994 GND.n1194 199.319
R5425 GND.n4993 GND.n1194 199.319
R5426 GND.n4135 GND.n2320 163.367
R5427 GND.n4133 GND.n4132 163.367
R5428 GND.n4130 GND.n2329 163.367
R5429 GND.n4126 GND.n4125 163.367
R5430 GND.n4123 GND.n2332 163.367
R5431 GND.n4119 GND.n4118 163.367
R5432 GND.n4116 GND.n2335 163.367
R5433 GND.n4112 GND.n4111 163.367
R5434 GND.n4109 GND.n2338 163.367
R5435 GND.n4105 GND.n4104 163.367
R5436 GND.n4102 GND.n2341 163.367
R5437 GND.n4098 GND.n4097 163.367
R5438 GND.n4095 GND.n2344 163.367
R5439 GND.n4091 GND.n4090 163.367
R5440 GND.n4088 GND.n2347 163.367
R5441 GND.n4083 GND.n4082 163.367
R5442 GND.n4080 GND.n2352 163.367
R5443 GND.n4075 GND.n4074 163.367
R5444 GND.n4072 GND.n2584 163.367
R5445 GND.n4067 GND.n4066 163.367
R5446 GND.n4064 GND.n2589 163.367
R5447 GND.n4060 GND.n4059 163.367
R5448 GND.n4057 GND.n2592 163.367
R5449 GND.n4053 GND.n4052 163.367
R5450 GND.n4050 GND.n2595 163.367
R5451 GND.n4046 GND.n4045 163.367
R5452 GND.n4043 GND.n2598 163.367
R5453 GND.n4039 GND.n4038 163.367
R5454 GND.n4036 GND.n2601 163.367
R5455 GND.n4032 GND.n4031 163.367
R5456 GND.n4029 GND.n2604 163.367
R5457 GND.n4025 GND.n4024 163.367
R5458 GND.n4022 GND.n2607 163.367
R5459 GND.n3650 GND.n3649 163.367
R5460 GND.n3650 GND.n2714 163.367
R5461 GND.n3654 GND.n2714 163.367
R5462 GND.n3654 GND.n1427 163.367
R5463 GND.n3666 GND.n1427 163.367
R5464 GND.n3666 GND.n1435 163.367
R5465 GND.n2706 GND.n1435 163.367
R5466 GND.n3672 GND.n2706 163.367
R5467 GND.n3672 GND.n2707 163.367
R5468 GND.n2707 GND.n1447 163.367
R5469 GND.n3713 GND.n1447 163.367
R5470 GND.n3713 GND.n1455 163.367
R5471 GND.n3717 GND.n1455 163.367
R5472 GND.n3718 GND.n3717 163.367
R5473 GND.n3719 GND.n3718 163.367
R5474 GND.n3719 GND.n1467 163.367
R5475 GND.n3725 GND.n1467 163.367
R5476 GND.n3725 GND.n1475 163.367
R5477 GND.n2684 GND.n1475 163.367
R5478 GND.n3758 GND.n2684 163.367
R5479 GND.n3759 GND.n3758 163.367
R5480 GND.n3759 GND.n1487 163.367
R5481 GND.n3769 GND.n1487 163.367
R5482 GND.n3769 GND.n1494 163.367
R5483 GND.n3765 GND.n1494 163.367
R5484 GND.n3765 GND.n2675 163.367
R5485 GND.n3762 GND.n2675 163.367
R5486 GND.n3762 GND.n1506 163.367
R5487 GND.n3811 GND.n1506 163.367
R5488 GND.n3811 GND.n1514 163.367
R5489 GND.n2667 GND.n1514 163.367
R5490 GND.n3828 GND.n2667 163.367
R5491 GND.n3828 GND.n2668 163.367
R5492 GND.n3824 GND.n2668 163.367
R5493 GND.n3824 GND.n2663 163.367
R5494 GND.n3821 GND.n2663 163.367
R5495 GND.n3821 GND.n1536 163.367
R5496 GND.n3817 GND.n1536 163.367
R5497 GND.n3817 GND.n1544 163.367
R5498 GND.n2656 GND.n1544 163.367
R5499 GND.n3854 GND.n2656 163.367
R5500 GND.n3854 GND.n1561 163.367
R5501 GND.n3858 GND.n1561 163.367
R5502 GND.n3858 GND.n1570 163.367
R5503 GND.n2653 GND.n1570 163.367
R5504 GND.n3866 GND.n2653 163.367
R5505 GND.n3866 GND.n2654 163.367
R5506 GND.n3862 GND.n2654 163.367
R5507 GND.n3862 GND.n2643 163.367
R5508 GND.n3907 GND.n2643 163.367
R5509 GND.n3907 GND.n1606 163.367
R5510 GND.n3911 GND.n1606 163.367
R5511 GND.n3911 GND.n1614 163.367
R5512 GND.n3915 GND.n1614 163.367
R5513 GND.n3919 GND.n3915 163.367
R5514 GND.n3919 GND.n1630 163.367
R5515 GND.n3923 GND.n1630 163.367
R5516 GND.n3923 GND.n1638 163.367
R5517 GND.n2640 GND.n1638 163.367
R5518 GND.n3953 GND.n2640 163.367
R5519 GND.n3953 GND.n2641 163.367
R5520 GND.n3949 GND.n2641 163.367
R5521 GND.n3949 GND.n2634 163.367
R5522 GND.n3946 GND.n2634 163.367
R5523 GND.n3946 GND.n1674 163.367
R5524 GND.n3942 GND.n1674 163.367
R5525 GND.n3942 GND.n1682 163.367
R5526 GND.n3938 GND.n1682 163.367
R5527 GND.n3938 GND.n3934 163.367
R5528 GND.n3934 GND.n1700 163.367
R5529 GND.n3930 GND.n1700 163.367
R5530 GND.n3930 GND.n1708 163.367
R5531 GND.n2616 GND.n1708 163.367
R5532 GND.n3990 GND.n2616 163.367
R5533 GND.n3991 GND.n3990 163.367
R5534 GND.n3992 GND.n3991 163.367
R5535 GND.n3992 GND.n2614 163.367
R5536 GND.n3996 GND.n2614 163.367
R5537 GND.n3996 GND.n1738 163.367
R5538 GND.n4009 GND.n1738 163.367
R5539 GND.n4009 GND.n1746 163.367
R5540 GND.n4013 GND.n1746 163.367
R5541 GND.n4014 GND.n4013 163.367
R5542 GND.n4014 GND.n2318 163.367
R5543 GND.n3564 GND.n3563 163.367
R5544 GND.n3639 GND.n3563 163.367
R5545 GND.n3637 GND.n3636 163.367
R5546 GND.n3633 GND.n3632 163.367
R5547 GND.n3629 GND.n3628 163.367
R5548 GND.n3625 GND.n3624 163.367
R5549 GND.n3621 GND.n3620 163.367
R5550 GND.n3617 GND.n3616 163.367
R5551 GND.n3613 GND.n3612 163.367
R5552 GND.n3609 GND.n3608 163.367
R5553 GND.n3605 GND.n3604 163.367
R5554 GND.n3601 GND.n3600 163.367
R5555 GND.n3597 GND.n3596 163.367
R5556 GND.n3593 GND.n3592 163.367
R5557 GND.n3589 GND.n3588 163.367
R5558 GND.n3584 GND.n3583 163.367
R5559 GND.n3580 GND.n3579 163.367
R5560 GND.n2756 GND.n2755 163.367
R5561 GND.n2760 GND.n2759 163.367
R5562 GND.n2764 GND.n2763 163.367
R5563 GND.n2768 GND.n2767 163.367
R5564 GND.n2772 GND.n2771 163.367
R5565 GND.n2776 GND.n2775 163.367
R5566 GND.n2780 GND.n2779 163.367
R5567 GND.n2784 GND.n2783 163.367
R5568 GND.n2788 GND.n2787 163.367
R5569 GND.n2792 GND.n2791 163.367
R5570 GND.n2796 GND.n2795 163.367
R5571 GND.n2800 GND.n2799 163.367
R5572 GND.n2804 GND.n2803 163.367
R5573 GND.n2808 GND.n2807 163.367
R5574 GND.n2810 GND.n2750 163.367
R5575 GND.n2815 GND.n2717 163.367
R5576 GND.n3573 GND.n3565 163.367
R5577 GND.n3573 GND.n3572 163.367
R5578 GND.n3572 GND.n1429 163.367
R5579 GND.n4903 GND.n1429 163.367
R5580 GND.n4903 GND.n1430 163.367
R5581 GND.n4899 GND.n1430 163.367
R5582 GND.n4899 GND.n1433 163.367
R5583 GND.n3674 GND.n1433 163.367
R5584 GND.n3674 GND.n1449 163.367
R5585 GND.n4889 GND.n1449 163.367
R5586 GND.n4889 GND.n1450 163.367
R5587 GND.n4885 GND.n1450 163.367
R5588 GND.n4885 GND.n1453 163.367
R5589 GND.n2695 GND.n1453 163.367
R5590 GND.n2695 GND.n1469 163.367
R5591 GND.n4875 GND.n1469 163.367
R5592 GND.n4875 GND.n1470 163.367
R5593 GND.n4871 GND.n1470 163.367
R5594 GND.n4871 GND.n1473 163.367
R5595 GND.n3756 GND.n1473 163.367
R5596 GND.n3756 GND.n1489 163.367
R5597 GND.n4861 GND.n1489 163.367
R5598 GND.n4861 GND.n1490 163.367
R5599 GND.n4857 GND.n1490 163.367
R5600 GND.n4857 GND.n1493 163.367
R5601 GND.n3790 GND.n1493 163.367
R5602 GND.n3790 GND.n1508 163.367
R5603 GND.n4847 GND.n1508 163.367
R5604 GND.n4847 GND.n1509 163.367
R5605 GND.n4843 GND.n1509 163.367
R5606 GND.n4843 GND.n1512 163.367
R5607 GND.n3831 GND.n1512 163.367
R5608 GND.n3832 GND.n3831 163.367
R5609 GND.n3832 GND.n2665 163.367
R5610 GND.n3836 GND.n2665 163.367
R5611 GND.n3836 GND.n1538 163.367
R5612 GND.n4826 GND.n1538 163.367
R5613 GND.n4826 GND.n1539 163.367
R5614 GND.n4822 GND.n1539 163.367
R5615 GND.n4822 GND.n1542 163.367
R5616 GND.n1564 GND.n1542 163.367
R5617 GND.n4813 GND.n1564 163.367
R5618 GND.n4813 GND.n1565 163.367
R5619 GND.n4809 GND.n1565 163.367
R5620 GND.n4809 GND.n1568 163.367
R5621 GND.n3874 GND.n1568 163.367
R5622 GND.n3874 GND.n3867 163.367
R5623 GND.n3870 GND.n3867 163.367
R5624 GND.n3870 GND.n3869 163.367
R5625 GND.n3869 GND.n1608 163.367
R5626 GND.n4792 GND.n1608 163.367
R5627 GND.n4792 GND.n1609 163.367
R5628 GND.n4788 GND.n1609 163.367
R5629 GND.n4788 GND.n1612 163.367
R5630 GND.n1632 GND.n1612 163.367
R5631 GND.n4778 GND.n1632 163.367
R5632 GND.n4778 GND.n1633 163.367
R5633 GND.n4774 GND.n1633 163.367
R5634 GND.n4774 GND.n1636 163.367
R5635 GND.n3956 GND.n1636 163.367
R5636 GND.n3957 GND.n3956 163.367
R5637 GND.n3957 GND.n2636 163.367
R5638 GND.n3961 GND.n2636 163.367
R5639 GND.n3961 GND.n1676 163.367
R5640 GND.n4757 GND.n1676 163.367
R5641 GND.n4757 GND.n1677 163.367
R5642 GND.n4753 GND.n1677 163.367
R5643 GND.n4753 GND.n1680 163.367
R5644 GND.n1702 GND.n1680 163.367
R5645 GND.n4744 GND.n1702 163.367
R5646 GND.n4744 GND.n1703 163.367
R5647 GND.n4740 GND.n1703 163.367
R5648 GND.n4740 GND.n1706 163.367
R5649 GND.n3988 GND.n1706 163.367
R5650 GND.n3988 GND.n3981 163.367
R5651 GND.n3984 GND.n3981 163.367
R5652 GND.n3984 GND.n3983 163.367
R5653 GND.n3983 GND.n1740 163.367
R5654 GND.n4723 GND.n1740 163.367
R5655 GND.n4723 GND.n1741 163.367
R5656 GND.n4719 GND.n1741 163.367
R5657 GND.n4719 GND.n1744 163.367
R5658 GND.n2319 GND.n1744 163.367
R5659 GND.n4140 GND.n2319 163.367
R5660 GND.n5075 GND.n1195 153.216
R5661 GND.n4078 GND.n2581 153.216
R5662 GND.n3570 GND.n3569 152
R5663 GND.n2326 GND.n2325 152
R5664 GND.n2751 GND.t72 148.726
R5665 GND.n2585 GND.t121 148.726
R5666 GND.n3577 GND.t119 148.72
R5667 GND.n2348 GND.t96 148.72
R5668 GND.n4077 GND.n2582 143.351
R5669 GND.n4077 GND.n4076 143.351
R5670 GND.n2734 GND.n2733 143.351
R5671 GND.n2735 GND.n2734 143.351
R5672 GND.n3568 GND.t114 138.431
R5673 GND.n2324 GND.t73 138.431
R5674 GND.n18 GND.t58 129.933
R5675 GND.n21 GND.t61 129.132
R5676 GND.n20 GND.t21 129.132
R5677 GND.n19 GND.t43 129.132
R5678 GND.n18 GND.t47 129.132
R5679 GND.n3569 GND.t66 126.766
R5680 GND.n2325 GND.t98 126.766
R5681 GND.n2432 GND.t104 106.886
R5682 GND.n6443 GND.n89 99.6594
R5683 GND.n6442 GND.n92 99.6594
R5684 GND.n6440 GND.n94 99.6594
R5685 GND.n6439 GND.n97 99.6594
R5686 GND.n6437 GND.n99 99.6594
R5687 GND.n6436 GND.n102 99.6594
R5688 GND.n6434 GND.n104 99.6594
R5689 GND.n6433 GND.n110 99.6594
R5690 GND.n6431 GND.n112 99.6594
R5691 GND.n6430 GND.n115 99.6594
R5692 GND.n6428 GND.n117 99.6594
R5693 GND.n6427 GND.n120 99.6594
R5694 GND.n6425 GND.n122 99.6594
R5695 GND.n6424 GND.n125 99.6594
R5696 GND.n6422 GND.n127 99.6594
R5697 GND.n6421 GND.n130 99.6594
R5698 GND.n6446 GND.n6445 99.6594
R5699 GND.n2366 GND.n1885 99.6594
R5700 GND.n2375 GND.n2374 99.6594
R5701 GND.n2378 GND.n2377 99.6594
R5702 GND.n2385 GND.n2384 99.6594
R5703 GND.n2388 GND.n2387 99.6594
R5704 GND.n2395 GND.n2394 99.6594
R5705 GND.n2400 GND.n2399 99.6594
R5706 GND.n2397 GND.n2355 99.6594
R5707 GND.n2577 GND.n2576 99.6594
R5708 GND.n2570 GND.n2409 99.6594
R5709 GND.n2569 GND.n2568 99.6594
R5710 GND.n2562 GND.n2415 99.6594
R5711 GND.n2561 GND.n2560 99.6594
R5712 GND.n2554 GND.n2421 99.6594
R5713 GND.n2553 GND.n2552 99.6594
R5714 GND.n2546 GND.n2427 99.6594
R5715 GND.n2545 GND.n2544 99.6594
R5716 GND.n5003 GND.n1176 99.6594
R5717 GND.n5002 GND.n1179 99.6594
R5718 GND.n5000 GND.n1181 99.6594
R5719 GND.n4999 GND.n1184 99.6594
R5720 GND.n4997 GND.n1186 99.6594
R5721 GND.n4996 GND.n1189 99.6594
R5722 GND.n4993 GND.n1196 99.6594
R5723 GND.n4992 GND.n1199 99.6594
R5724 GND.n4990 GND.n1201 99.6594
R5725 GND.n4989 GND.n1204 99.6594
R5726 GND.n4987 GND.n1206 99.6594
R5727 GND.n4986 GND.n1209 99.6594
R5728 GND.n4984 GND.n1211 99.6594
R5729 GND.n4983 GND.n1214 99.6594
R5730 GND.n4981 GND.n1216 99.6594
R5731 GND.n4980 GND.n1165 99.6594
R5732 GND.n5263 GND.n5262 99.6594
R5733 GND.n5257 GND.n942 99.6594
R5734 GND.n5254 GND.n943 99.6594
R5735 GND.n5250 GND.n944 99.6594
R5736 GND.n5246 GND.n945 99.6594
R5737 GND.n5242 GND.n946 99.6594
R5738 GND.n5238 GND.n947 99.6594
R5739 GND.n5234 GND.n948 99.6594
R5740 GND.n5229 GND.n949 99.6594
R5741 GND.n5225 GND.n950 99.6594
R5742 GND.n5221 GND.n951 99.6594
R5743 GND.n5217 GND.n952 99.6594
R5744 GND.n5213 GND.n953 99.6594
R5745 GND.n5209 GND.n954 99.6594
R5746 GND.n5205 GND.n955 99.6594
R5747 GND.n5201 GND.n956 99.6594
R5748 GND.n5197 GND.n957 99.6594
R5749 GND.n1277 GND.n1223 99.6594
R5750 GND.n1279 GND.n1226 99.6594
R5751 GND.n1281 GND.n1280 99.6594
R5752 GND.n1285 GND.n1284 99.6594
R5753 GND.n1286 GND.n1255 99.6594
R5754 GND.n1288 GND.n1262 99.6594
R5755 GND.n1290 GND.n1289 99.6594
R5756 GND.n5006 GND.n5005 99.6594
R5757 GND.n5190 GND.n958 99.6594
R5758 GND.n3069 GND.n959 99.6594
R5759 GND.n3074 GND.n960 99.6594
R5760 GND.n3066 GND.n961 99.6594
R5761 GND.n3082 GND.n962 99.6594
R5762 GND.n3062 GND.n963 99.6594
R5763 GND.n3090 GND.n964 99.6594
R5764 GND.n3058 GND.n965 99.6594
R5765 GND.n2462 GND.n2461 99.6594
R5766 GND.n2465 GND.n2464 99.6594
R5767 GND.n2477 GND.n2476 99.6594
R5768 GND.n2487 GND.n2486 99.6594
R5769 GND.n2492 GND.n2489 99.6594
R5770 GND.n2490 GND.n2250 99.6594
R5771 GND.n2253 GND.n2252 99.6594
R5772 GND.n2258 GND.n2257 99.6594
R5773 GND.n2261 GND.n2260 99.6594
R5774 GND.n2266 GND.n2265 99.6594
R5775 GND.n2269 GND.n2268 99.6594
R5776 GND.n2274 GND.n2273 99.6594
R5777 GND.n2279 GND.n2278 99.6594
R5778 GND.n4190 GND.n4189 99.6594
R5779 GND.n5031 GND.n5030 99.6594
R5780 GND.n1248 GND.n1234 99.6594
R5781 GND.n1259 GND.n1235 99.6594
R5782 GND.n1267 GND.n1236 99.6594
R5783 GND.n1269 GND.n1237 99.6594
R5784 GND.n3471 GND.n1238 99.6594
R5785 GND.n3475 GND.n1239 99.6594
R5786 GND.n3483 GND.n1240 99.6594
R5787 GND.n3485 GND.n1241 99.6594
R5788 GND.n3493 GND.n1242 99.6594
R5789 GND.n3495 GND.n1243 99.6594
R5790 GND.n3503 GND.n1244 99.6594
R5791 GND.n3505 GND.n1245 99.6594
R5792 GND.n3513 GND.n1246 99.6594
R5793 GND.n5030 GND.n1232 99.6594
R5794 GND.n1258 GND.n1234 99.6594
R5795 GND.n1266 GND.n1235 99.6594
R5796 GND.n1268 GND.n1236 99.6594
R5797 GND.n3470 GND.n1237 99.6594
R5798 GND.n3476 GND.n1238 99.6594
R5799 GND.n3482 GND.n1239 99.6594
R5800 GND.n3486 GND.n1240 99.6594
R5801 GND.n3492 GND.n1241 99.6594
R5802 GND.n3496 GND.n1242 99.6594
R5803 GND.n3502 GND.n1243 99.6594
R5804 GND.n3506 GND.n1244 99.6594
R5805 GND.n3512 GND.n1245 99.6594
R5806 GND.n3515 GND.n1246 99.6594
R5807 GND.n4189 GND.n4188 99.6594
R5808 GND.n2278 GND.n2277 99.6594
R5809 GND.n2273 GND.n2272 99.6594
R5810 GND.n2268 GND.n2267 99.6594
R5811 GND.n2265 GND.n2264 99.6594
R5812 GND.n2260 GND.n2259 99.6594
R5813 GND.n2257 GND.n2256 99.6594
R5814 GND.n2252 GND.n2251 99.6594
R5815 GND.n2491 GND.n2490 99.6594
R5816 GND.n2489 GND.n2488 99.6594
R5817 GND.n2486 GND.n2478 99.6594
R5818 GND.n2476 GND.n2475 99.6594
R5819 GND.n2464 GND.n2463 99.6594
R5820 GND.n2461 GND.n2449 99.6594
R5821 GND.n3068 GND.n958 99.6594
R5822 GND.n3073 GND.n959 99.6594
R5823 GND.n3065 GND.n960 99.6594
R5824 GND.n3081 GND.n961 99.6594
R5825 GND.n3061 GND.n962 99.6594
R5826 GND.n3089 GND.n963 99.6594
R5827 GND.n3057 GND.n964 99.6594
R5828 GND.n3053 GND.n965 99.6594
R5829 GND.n5005 GND.n1274 99.6594
R5830 GND.n1290 GND.n1263 99.6594
R5831 GND.n1288 GND.n1287 99.6594
R5832 GND.n1286 GND.n1254 99.6594
R5833 GND.n1285 GND.n1283 99.6594
R5834 GND.n1280 GND.n1227 99.6594
R5835 GND.n1279 GND.n1278 99.6594
R5836 GND.n1277 GND.n1222 99.6594
R5837 GND.n5263 GND.n969 99.6594
R5838 GND.n5255 GND.n942 99.6594
R5839 GND.n5251 GND.n943 99.6594
R5840 GND.n5247 GND.n944 99.6594
R5841 GND.n5243 GND.n945 99.6594
R5842 GND.n5239 GND.n946 99.6594
R5843 GND.n5235 GND.n947 99.6594
R5844 GND.n5230 GND.n948 99.6594
R5845 GND.n5226 GND.n949 99.6594
R5846 GND.n5222 GND.n950 99.6594
R5847 GND.n5218 GND.n951 99.6594
R5848 GND.n5214 GND.n952 99.6594
R5849 GND.n5210 GND.n953 99.6594
R5850 GND.n5206 GND.n954 99.6594
R5851 GND.n5202 GND.n955 99.6594
R5852 GND.n5198 GND.n956 99.6594
R5853 GND.n1015 GND.n957 99.6594
R5854 GND.n4980 GND.n4979 99.6594
R5855 GND.n4981 GND.n1215 99.6594
R5856 GND.n4983 GND.n4982 99.6594
R5857 GND.n4984 GND.n1210 99.6594
R5858 GND.n4986 GND.n4985 99.6594
R5859 GND.n4987 GND.n1205 99.6594
R5860 GND.n4989 GND.n4988 99.6594
R5861 GND.n4990 GND.n1200 99.6594
R5862 GND.n4992 GND.n4991 99.6594
R5863 GND.n4994 GND.n1190 99.6594
R5864 GND.n4996 GND.n4995 99.6594
R5865 GND.n4997 GND.n1185 99.6594
R5866 GND.n4999 GND.n4998 99.6594
R5867 GND.n5000 GND.n1180 99.6594
R5868 GND.n5002 GND.n5001 99.6594
R5869 GND.n5003 GND.n1175 99.6594
R5870 GND.n2367 GND.n2366 99.6594
R5871 GND.n2376 GND.n2375 99.6594
R5872 GND.n2377 GND.n2362 99.6594
R5873 GND.n2386 GND.n2385 99.6594
R5874 GND.n2387 GND.n2358 99.6594
R5875 GND.n2396 GND.n2395 99.6594
R5876 GND.n2399 GND.n2398 99.6594
R5877 GND.n2579 GND.n2578 99.6594
R5878 GND.n2576 GND.n2575 99.6594
R5879 GND.n2571 GND.n2570 99.6594
R5880 GND.n2568 GND.n2567 99.6594
R5881 GND.n2563 GND.n2562 99.6594
R5882 GND.n2560 GND.n2559 99.6594
R5883 GND.n2555 GND.n2554 99.6594
R5884 GND.n2552 GND.n2551 99.6594
R5885 GND.n2547 GND.n2546 99.6594
R5886 GND.n2544 GND.n2543 99.6594
R5887 GND.n6445 GND.n133 99.6594
R5888 GND.n6421 GND.n6420 99.6594
R5889 GND.n6422 GND.n126 99.6594
R5890 GND.n6424 GND.n6423 99.6594
R5891 GND.n6425 GND.n121 99.6594
R5892 GND.n6427 GND.n6426 99.6594
R5893 GND.n6428 GND.n116 99.6594
R5894 GND.n6430 GND.n6429 99.6594
R5895 GND.n6431 GND.n111 99.6594
R5896 GND.n6433 GND.n6432 99.6594
R5897 GND.n6434 GND.n103 99.6594
R5898 GND.n6436 GND.n6435 99.6594
R5899 GND.n6437 GND.n98 99.6594
R5900 GND.n6439 GND.n6438 99.6594
R5901 GND.n6440 GND.n93 99.6594
R5902 GND.n6442 GND.n6441 99.6594
R5903 GND.n6443 GND.n88 99.6594
R5904 GND.n2536 GND.n2535 99.6594
R5905 GND.n2444 GND.n2441 99.6594
R5906 GND.n2453 GND.n2446 99.6594
R5907 GND.n2456 GND.n2455 99.6594
R5908 GND.n2468 GND.n2458 99.6594
R5909 GND.n2471 GND.n2470 99.6594
R5910 GND.n2482 GND.n2481 99.6594
R5911 GND.n2500 GND.n2499 99.6594
R5912 GND.n2535 GND.n2534 99.6594
R5913 GND.n2445 GND.n2444 99.6594
R5914 GND.n2454 GND.n2453 99.6594
R5915 GND.n2457 GND.n2456 99.6594
R5916 GND.n2469 GND.n2468 99.6594
R5917 GND.n2472 GND.n2471 99.6594
R5918 GND.n2483 GND.n2482 99.6594
R5919 GND.n2499 GND.n2498 99.6594
R5920 GND.n1999 GND.n136 99.6594
R5921 GND.n2001 GND.n137 99.6594
R5922 GND.n2005 GND.n138 99.6594
R5923 GND.n2007 GND.n139 99.6594
R5924 GND.n2011 GND.n140 99.6594
R5925 GND.n2013 GND.n141 99.6594
R5926 GND.n2017 GND.n142 99.6594
R5927 GND.n2019 GND.n143 99.6594
R5928 GND.n2022 GND.n143 99.6594
R5929 GND.n2018 GND.n142 99.6594
R5930 GND.n2016 GND.n141 99.6594
R5931 GND.n2012 GND.n140 99.6594
R5932 GND.n2010 GND.n139 99.6594
R5933 GND.n2006 GND.n138 99.6594
R5934 GND.n2004 GND.n137 99.6594
R5935 GND.n2000 GND.n136 99.6594
R5936 GND.n2275 GND.t125 98.1201
R5937 GND.n2833 GND.t87 98.1201
R5938 GND.n2020 GND.t82 97.2868
R5939 GND.n107 GND.t134 97.2868
R5940 GND.n131 GND.t112 97.2868
R5941 GND.n1191 GND.t89 97.2868
R5942 GND.n1217 GND.t64 97.2868
R5943 GND.n1272 GND.t92 97.2868
R5944 GND.n3054 GND.t110 97.2868
R5945 GND.n2405 GND.t129 97.2868
R5946 GND.n987 GND.t79 97.2868
R5947 GND.n1007 GND.t132 97.2868
R5948 GND.n2501 GND.t107 97.2868
R5949 GND.n2752 GND.n2751 93.0914
R5950 GND.n2586 GND.n2585 93.0914
R5951 GND.n3578 GND.n3577 93.0914
R5952 GND.n2349 GND.n2348 93.0914
R5953 GND.n3568 GND.n3567 73.571
R5954 GND.n2324 GND.n2323 73.571
R5955 GND.n4134 GND.n4133 71.676
R5956 GND.n4131 GND.n4130 71.676
R5957 GND.n4126 GND.n2331 71.676
R5958 GND.n4124 GND.n4123 71.676
R5959 GND.n4119 GND.n2334 71.676
R5960 GND.n4117 GND.n4116 71.676
R5961 GND.n4112 GND.n2337 71.676
R5962 GND.n4110 GND.n4109 71.676
R5963 GND.n4105 GND.n2340 71.676
R5964 GND.n4103 GND.n4102 71.676
R5965 GND.n4098 GND.n2343 71.676
R5966 GND.n4096 GND.n4095 71.676
R5967 GND.n4091 GND.n2346 71.676
R5968 GND.n4089 GND.n4088 71.676
R5969 GND.n4083 GND.n2351 71.676
R5970 GND.n4081 GND.n4080 71.676
R5971 GND.n4076 GND.n4075 71.676
R5972 GND.n4073 GND.n4072 71.676
R5973 GND.n4067 GND.n2588 71.676
R5974 GND.n4065 GND.n4064 71.676
R5975 GND.n4060 GND.n2591 71.676
R5976 GND.n4058 GND.n4057 71.676
R5977 GND.n4053 GND.n2594 71.676
R5978 GND.n4051 GND.n4050 71.676
R5979 GND.n4046 GND.n2597 71.676
R5980 GND.n4044 GND.n4043 71.676
R5981 GND.n4039 GND.n2600 71.676
R5982 GND.n4037 GND.n4036 71.676
R5983 GND.n4032 GND.n2603 71.676
R5984 GND.n4030 GND.n4029 71.676
R5985 GND.n4025 GND.n2606 71.676
R5986 GND.n4023 GND.n4022 71.676
R5987 GND.n4018 GND.n4017 71.676
R5988 GND.n3645 GND.n3644 71.676
R5989 GND.n3639 GND.n2718 71.676
R5990 GND.n3636 GND.n2719 71.676
R5991 GND.n3632 GND.n2720 71.676
R5992 GND.n3628 GND.n2721 71.676
R5993 GND.n3624 GND.n2722 71.676
R5994 GND.n3620 GND.n2723 71.676
R5995 GND.n3616 GND.n2724 71.676
R5996 GND.n3612 GND.n2725 71.676
R5997 GND.n3608 GND.n2726 71.676
R5998 GND.n3604 GND.n2727 71.676
R5999 GND.n3600 GND.n2728 71.676
R6000 GND.n3596 GND.n2729 71.676
R6001 GND.n3592 GND.n2730 71.676
R6002 GND.n3588 GND.n2731 71.676
R6003 GND.n3583 GND.n2732 71.676
R6004 GND.n3579 GND.n2733 71.676
R6005 GND.n2756 GND.n2736 71.676
R6006 GND.n2760 GND.n2737 71.676
R6007 GND.n2764 GND.n2738 71.676
R6008 GND.n2768 GND.n2739 71.676
R6009 GND.n2772 GND.n2740 71.676
R6010 GND.n2776 GND.n2741 71.676
R6011 GND.n2780 GND.n2742 71.676
R6012 GND.n2784 GND.n2743 71.676
R6013 GND.n2788 GND.n2744 71.676
R6014 GND.n2792 GND.n2745 71.676
R6015 GND.n2796 GND.n2746 71.676
R6016 GND.n2800 GND.n2747 71.676
R6017 GND.n2804 GND.n2748 71.676
R6018 GND.n2808 GND.n2749 71.676
R6019 GND.n2816 GND.n2750 71.676
R6020 GND.n3647 GND.n2717 71.676
R6021 GND.n3645 GND.n3564 71.676
R6022 GND.n3637 GND.n2718 71.676
R6023 GND.n3633 GND.n2719 71.676
R6024 GND.n3629 GND.n2720 71.676
R6025 GND.n3625 GND.n2721 71.676
R6026 GND.n3621 GND.n2722 71.676
R6027 GND.n3617 GND.n2723 71.676
R6028 GND.n3613 GND.n2724 71.676
R6029 GND.n3609 GND.n2725 71.676
R6030 GND.n3605 GND.n2726 71.676
R6031 GND.n3601 GND.n2727 71.676
R6032 GND.n3597 GND.n2728 71.676
R6033 GND.n3593 GND.n2729 71.676
R6034 GND.n3589 GND.n2730 71.676
R6035 GND.n3584 GND.n2731 71.676
R6036 GND.n3580 GND.n2732 71.676
R6037 GND.n2755 GND.n2735 71.676
R6038 GND.n2759 GND.n2736 71.676
R6039 GND.n2763 GND.n2737 71.676
R6040 GND.n2767 GND.n2738 71.676
R6041 GND.n2771 GND.n2739 71.676
R6042 GND.n2775 GND.n2740 71.676
R6043 GND.n2779 GND.n2741 71.676
R6044 GND.n2783 GND.n2742 71.676
R6045 GND.n2787 GND.n2743 71.676
R6046 GND.n2791 GND.n2744 71.676
R6047 GND.n2795 GND.n2745 71.676
R6048 GND.n2799 GND.n2746 71.676
R6049 GND.n2803 GND.n2747 71.676
R6050 GND.n2807 GND.n2748 71.676
R6051 GND.n2810 GND.n2749 71.676
R6052 GND.n2816 GND.n2815 71.676
R6053 GND.n3648 GND.n3647 71.676
R6054 GND.n4017 GND.n2607 71.676
R6055 GND.n4024 GND.n4023 71.676
R6056 GND.n2606 GND.n2604 71.676
R6057 GND.n4031 GND.n4030 71.676
R6058 GND.n2603 GND.n2601 71.676
R6059 GND.n4038 GND.n4037 71.676
R6060 GND.n2600 GND.n2598 71.676
R6061 GND.n4045 GND.n4044 71.676
R6062 GND.n2597 GND.n2595 71.676
R6063 GND.n4052 GND.n4051 71.676
R6064 GND.n2594 GND.n2592 71.676
R6065 GND.n4059 GND.n4058 71.676
R6066 GND.n2591 GND.n2589 71.676
R6067 GND.n4066 GND.n4065 71.676
R6068 GND.n2588 GND.n2584 71.676
R6069 GND.n4074 GND.n4073 71.676
R6070 GND.n2582 GND.n2352 71.676
R6071 GND.n4082 GND.n4081 71.676
R6072 GND.n2351 GND.n2347 71.676
R6073 GND.n4090 GND.n4089 71.676
R6074 GND.n2346 GND.n2344 71.676
R6075 GND.n4097 GND.n4096 71.676
R6076 GND.n2343 GND.n2341 71.676
R6077 GND.n4104 GND.n4103 71.676
R6078 GND.n2340 GND.n2338 71.676
R6079 GND.n4111 GND.n4110 71.676
R6080 GND.n2337 GND.n2335 71.676
R6081 GND.n4118 GND.n4117 71.676
R6082 GND.n2334 GND.n2332 71.676
R6083 GND.n4125 GND.n4124 71.676
R6084 GND.n2331 GND.n2329 71.676
R6085 GND.n4132 GND.n4131 71.676
R6086 GND.n4135 GND.n4134 71.676
R6087 GND.n3576 GND.n3570 63.641
R6088 GND.n22 GND.t5 62.4417
R6089 GND.n25 GND.t37 61.6413
R6090 GND.n24 GND.t140 61.6413
R6091 GND.n23 GND.t137 61.6413
R6092 GND.n22 GND.t56 61.6413
R6093 GND.n2021 GND.t83 56.3656
R6094 GND.n108 GND.t135 56.3656
R6095 GND.n132 GND.t113 56.3656
R6096 GND.n1192 GND.t90 56.3656
R6097 GND.n1218 GND.t65 56.3656
R6098 GND.n1273 GND.t93 56.3656
R6099 GND.n3055 GND.t109 56.3656
R6100 GND.n2406 GND.t128 56.3656
R6101 GND.n988 GND.t78 56.3656
R6102 GND.n1008 GND.t131 56.3656
R6103 GND.n2502 GND.t106 56.3656
R6104 GND.n2276 GND.t126 56.2292
R6105 GND.n2834 GND.t86 56.2292
R6106 GND.n2752 GND.t71 55.6357
R6107 GND.n2586 GND.t122 55.6357
R6108 GND.n3578 GND.t118 55.6288
R6109 GND.n2349 GND.t97 55.6288
R6110 GND.n2433 GND.n2432 53.7217
R6111 GND.n6 GND.t12 53.5112
R6112 GND.n11 GND.t53 53.5112
R6113 GND.n1 GND.t30 53.5112
R6114 GND.n28 GND.t54 53.5112
R6115 GND.n33 GND.t34 53.5112
R6116 GND.n39 GND.t40 53.5112
R6117 GND.n2433 GND.t103 53.1656
R6118 GND.n2753 GND.n2752 53.1399
R6119 GND.n4070 GND.n2586 53.1399
R6120 GND.n3586 GND.n3578 53.1399
R6121 GND.n4085 GND.n2349 53.1399
R6122 GND.n9 GND.t45 52.7152
R6123 GND.n14 GND.t51 52.7152
R6124 GND.n4 GND.t50 52.7152
R6125 GND.n31 GND.t1 52.7152
R6126 GND.n36 GND.t14 52.7152
R6127 GND.n42 GND.t39 52.7152
R6128 GND.n2434 GND.n2433 48.6793
R6129 GND.n6 GND.n5 45.2716
R6130 GND.n8 GND.n7 45.2716
R6131 GND.n11 GND.n10 45.2716
R6132 GND.n13 GND.n12 45.2716
R6133 GND.n1 GND.n0 45.2716
R6134 GND.n3 GND.n2 45.2716
R6135 GND.n30 GND.n29 45.2716
R6136 GND.n28 GND.n27 45.2716
R6137 GND.n35 GND.n34 45.2716
R6138 GND.n33 GND.n32 45.2716
R6139 GND.n41 GND.n40 45.2716
R6140 GND.n39 GND.n38 45.2716
R6141 GND.n4138 GND.n2326 44.3322
R6142 GND.n2276 GND.n2275 41.8914
R6143 GND.n2834 GND.n2833 41.8914
R6144 GND.n2021 GND.n2020 40.9217
R6145 GND.n108 GND.n107 40.9217
R6146 GND.n132 GND.n131 40.9217
R6147 GND.n1192 GND.n1191 40.9217
R6148 GND.n1218 GND.n1217 40.9217
R6149 GND.n1273 GND.n1272 40.9217
R6150 GND.n3055 GND.n3054 40.9217
R6151 GND.n2406 GND.n2405 40.9217
R6152 GND.n988 GND.n987 40.9217
R6153 GND.n1008 GND.n1007 40.9217
R6154 GND.n2502 GND.n2501 40.9217
R6155 GND.n5458 GND.n5457 39.5582
R6156 GND.n5457 GND.n5456 39.5582
R6157 GND.n5456 GND.n751 39.5582
R6158 GND.n5450 GND.n751 39.5582
R6159 GND.n5450 GND.n5449 39.5582
R6160 GND.n5449 GND.n5448 39.5582
R6161 GND.n5448 GND.n758 39.5582
R6162 GND.n5442 GND.n758 39.5582
R6163 GND.n5442 GND.n5441 39.5582
R6164 GND.n5441 GND.n5440 39.5582
R6165 GND.n5440 GND.n766 39.5582
R6166 GND.n5434 GND.n766 39.5582
R6167 GND.n5434 GND.n5433 39.5582
R6168 GND.n5433 GND.n5432 39.5582
R6169 GND.n5432 GND.n774 39.5582
R6170 GND.n5426 GND.n774 39.5582
R6171 GND.n5426 GND.n5425 39.5582
R6172 GND.n5425 GND.n5424 39.5582
R6173 GND.n5424 GND.n782 39.5582
R6174 GND.n5418 GND.n782 39.5582
R6175 GND.n5418 GND.n5417 39.5582
R6176 GND.n5417 GND.n5416 39.5582
R6177 GND.n5416 GND.n790 39.5582
R6178 GND.n5410 GND.n790 39.5582
R6179 GND.n5410 GND.n5409 39.5582
R6180 GND.n5409 GND.n5408 39.5582
R6181 GND.n5408 GND.n798 39.5582
R6182 GND.n5402 GND.n798 39.5582
R6183 GND.n5402 GND.n5401 39.5582
R6184 GND.n5401 GND.n5400 39.5582
R6185 GND.n5400 GND.n806 39.5582
R6186 GND.n5394 GND.n806 39.5582
R6187 GND.n5394 GND.n5393 39.5582
R6188 GND.n5393 GND.n5392 39.5582
R6189 GND.n5392 GND.n814 39.5582
R6190 GND.n5386 GND.n814 39.5582
R6191 GND.n5386 GND.n5385 39.5582
R6192 GND.n5385 GND.n5384 39.5582
R6193 GND.n5384 GND.n822 39.5582
R6194 GND.n5378 GND.n822 39.5582
R6195 GND.n5378 GND.n5377 39.5582
R6196 GND.n5377 GND.n5376 39.5582
R6197 GND.n5376 GND.n830 39.5582
R6198 GND.n5370 GND.n830 39.5582
R6199 GND.n5370 GND.n5369 39.5582
R6200 GND.n5369 GND.n5368 39.5582
R6201 GND.n5368 GND.n838 39.5582
R6202 GND.n5362 GND.n838 39.5582
R6203 GND.n5362 GND.n5361 39.5582
R6204 GND.n5361 GND.n5360 39.5582
R6205 GND.n5360 GND.n846 39.5582
R6206 GND.n5354 GND.n846 39.5582
R6207 GND.n5354 GND.n5353 39.5582
R6208 GND.n5353 GND.n5352 39.5582
R6209 GND.n5352 GND.n854 39.5582
R6210 GND.n5346 GND.n854 39.5582
R6211 GND.n5346 GND.n5345 39.5582
R6212 GND.n5345 GND.n5344 39.5582
R6213 GND.n5344 GND.n862 39.5582
R6214 GND.n5338 GND.n862 39.5582
R6215 GND.n2023 GND.n2021 35.8793
R6216 GND.n109 GND.n108 35.8793
R6217 GND.n6448 GND.n132 35.8793
R6218 GND.n1219 GND.n1218 35.8793
R6219 GND.n5008 GND.n1273 35.8793
R6220 GND.n3096 GND.n3055 35.8793
R6221 GND.n4196 GND.n2276 35.8793
R6222 GND.n2835 GND.n2834 35.8793
R6223 GND.n5232 GND.n988 35.8793
R6224 GND.n5196 GND.n1008 35.8793
R6225 GND.n2503 GND.n2502 35.8793
R6226 GND.n3569 GND.n3568 34.8345
R6227 GND.n2325 GND.n2324 34.8345
R6228 GND.n4019 GND.n4016 34.4981
R6229 GND.n2716 GND.n2715 34.4981
R6230 GND.n5337 GND.n5336 31.1311
R6231 GND.n5336 GND.n869 31.1311
R6232 GND.n5330 GND.n869 31.1311
R6233 GND.n5330 GND.n5329 31.1311
R6234 GND.n5329 GND.n5328 31.1311
R6235 GND.n5328 GND.n878 31.1311
R6236 GND.n5322 GND.n878 31.1311
R6237 GND.n5322 GND.n5321 31.1311
R6238 GND.n5321 GND.n5320 31.1311
R6239 GND.n5320 GND.n886 31.1311
R6240 GND.n5314 GND.n886 31.1311
R6241 GND.n5314 GND.n5313 31.1311
R6242 GND.n5313 GND.n5312 31.1311
R6243 GND.n5312 GND.n894 31.1311
R6244 GND.n5306 GND.n894 31.1311
R6245 GND.n5306 GND.n5305 31.1311
R6246 GND.n5305 GND.n5304 31.1311
R6247 GND.n5304 GND.n902 31.1311
R6248 GND.n5298 GND.n902 31.1311
R6249 GND.n5298 GND.n5297 31.1311
R6250 GND.n5297 GND.n5296 31.1311
R6251 GND.n5296 GND.n910 31.1311
R6252 GND.n5290 GND.n910 31.1311
R6253 GND.n5290 GND.n5289 31.1311
R6254 GND.n5289 GND.n5288 31.1311
R6255 GND.n5288 GND.n918 31.1311
R6256 GND.n5282 GND.n918 31.1311
R6257 GND.n5282 GND.n5281 31.1311
R6258 GND.n5281 GND.n5280 31.1311
R6259 GND.n5280 GND.n926 31.1311
R6260 GND.n5274 GND.n926 31.1311
R6261 GND.n5274 GND.n5273 31.1311
R6262 GND.n5273 GND.n5272 31.1311
R6263 GND.n5272 GND.n934 31.1311
R6264 GND.n5266 GND.n934 31.1311
R6265 GND.n5266 GND.n5265 31.1311
R6266 GND.n1014 GND.n967 31.1311
R6267 GND.n1276 GND.n1168 31.1311
R6268 GND.n4978 GND.n1291 31.1311
R6269 GND.n1291 GND.n1233 31.1311
R6270 GND.n4970 GND.n1247 31.1311
R6271 GND.n4654 GND.n1860 31.1311
R6272 GND.n4648 GND.n4647 31.1311
R6273 GND.n4647 GND.n4646 31.1311
R6274 GND.n4640 GND.n1880 31.1311
R6275 GND.n135 GND.n81 31.1311
R6276 GND.n6419 GND.n144 31.1311
R6277 GND.n6413 GND.n144 31.1311
R6278 GND.n6413 GND.n6412 31.1311
R6279 GND.n6412 GND.n6411 31.1311
R6280 GND.n6411 GND.n153 31.1311
R6281 GND.n6405 GND.n153 31.1311
R6282 GND.n6405 GND.n6404 31.1311
R6283 GND.n6404 GND.n6403 31.1311
R6284 GND.n6403 GND.n161 31.1311
R6285 GND.n6397 GND.n161 31.1311
R6286 GND.n6397 GND.n6396 31.1311
R6287 GND.n6396 GND.n6395 31.1311
R6288 GND.n6395 GND.n169 31.1311
R6289 GND.n6389 GND.n169 31.1311
R6290 GND.n6389 GND.n6388 31.1311
R6291 GND.n6388 GND.n6387 31.1311
R6292 GND.n6387 GND.n177 31.1311
R6293 GND.n6381 GND.n177 31.1311
R6294 GND.n6381 GND.n6380 31.1311
R6295 GND.n6380 GND.n6379 31.1311
R6296 GND.n6379 GND.n185 31.1311
R6297 GND.n6373 GND.n185 31.1311
R6298 GND.n6373 GND.n6372 31.1311
R6299 GND.n6372 GND.n6371 31.1311
R6300 GND.n6371 GND.n193 31.1311
R6301 GND.n6365 GND.n193 31.1311
R6302 GND.n6365 GND.n6364 31.1311
R6303 GND.n6364 GND.n6363 31.1311
R6304 GND.n6363 GND.n201 31.1311
R6305 GND.n6357 GND.n201 31.1311
R6306 GND.n6357 GND.n6356 31.1311
R6307 GND.n6356 GND.n6355 31.1311
R6308 GND.n6355 GND.n209 31.1311
R6309 GND.n6349 GND.n209 31.1311
R6310 GND.n6349 GND.n6348 31.1311
R6311 GND.n6348 GND.n6347 31.1311
R6312 GND.n5075 GND.n1192 30.5518
R6313 GND.n2581 GND.n2406 30.5518
R6314 GND.n3576 GND.n3575 21.0737
R6315 GND.n4139 GND.n4138 21.0737
R6316 GND.n5004 GND.n1276 20.2354
R6317 GND.n1880 GND.n1872 20.2354
R6318 GND.n5188 GND.n1014 19.9241
R6319 GND.n5187 GND.n1018 19.9241
R6320 GND.n1033 GND.n1032 19.9241
R6321 GND.n5181 GND.n5180 19.9241
R6322 GND.n3107 GND.n3105 19.9241
R6323 GND.n5174 GND.n1051 19.9241
R6324 GND.n3115 GND.n1054 19.9241
R6325 GND.n3140 GND.n3138 19.9241
R6326 GND.n3152 GND.n3043 19.9241
R6327 GND.n3142 GND.n3045 19.9241
R6328 GND.n3166 GND.n3036 19.9241
R6329 GND.n3170 GND.n3031 19.9241
R6330 GND.n3181 GND.n3180 19.9241
R6331 GND.n3021 GND.n3011 19.9241
R6332 GND.n3192 GND.n3191 19.9241
R6333 GND.n3205 GND.n3001 19.9241
R6334 GND.n3202 GND.n3004 19.9241
R6335 GND.n3216 GND.n3215 19.9241
R6336 GND.n2991 GND.n2983 19.9241
R6337 GND.n3229 GND.n3227 19.9241
R6338 GND.n3284 GND.n2951 19.9241
R6339 GND.n3281 GND.n2953 19.9241
R6340 GND.n3237 GND.n2964 19.9241
R6341 GND.n3273 GND.n3272 19.9241
R6342 GND.n3267 GND.n2966 19.9241
R6343 GND.n3263 GND.n2975 19.9241
R6344 GND.n3262 GND.n3251 19.9241
R6345 GND.n3292 GND.n2935 19.9241
R6346 GND.n2936 GND.n2928 19.9241
R6347 GND.n3302 GND.n3301 19.9241
R6348 GND.n3372 GND.n2917 19.9241
R6349 GND.n3369 GND.n2920 19.9241
R6350 GND.n2911 GND.n2907 19.9241
R6351 GND.n3391 GND.n2899 19.9241
R6352 GND.n3397 GND.n2895 19.9241
R6353 GND.n3394 GND.n2897 19.9241
R6354 GND.n3407 GND.n2887 19.9241
R6355 GND.n3356 GND.n3355 19.9241
R6356 GND.n3416 GND.n2880 19.9241
R6357 GND.n3422 GND.n2876 19.9241
R6358 GND.n3418 GND.n2878 19.9241
R6359 GND.n3432 GND.n2865 19.9241
R6360 GND.n2870 GND.n2867 19.9241
R6361 GND.n3447 GND.n2858 19.9241
R6362 GND.n3450 GND.n2853 19.9241
R6363 GND.n3458 GND.n2847 19.9241
R6364 GND.n3463 GND.n2845 19.9241
R6365 GND.n5100 GND.n1166 19.9241
R6366 GND.n4639 GND.n1883 19.9241
R6367 GND.n2245 GND.n1892 19.9241
R6368 GND.n4633 GND.n1895 19.9241
R6369 GND.n4226 GND.n2237 19.9241
R6370 GND.n4289 GND.n2233 19.9241
R6371 GND.n4295 GND.n2235 19.9241
R6372 GND.n4292 GND.n2222 19.9241
R6373 GND.n4305 GND.n2223 19.9241
R6374 GND.n2227 GND.n2215 19.9241
R6375 GND.n4314 GND.n2211 19.9241
R6376 GND.n4320 GND.n2213 19.9241
R6377 GND.n4316 GND.n2200 19.9241
R6378 GND.n4330 GND.n2202 19.9241
R6379 GND.n2205 GND.n2193 19.9241
R6380 GND.n4339 GND.n2188 19.9241
R6381 GND.n4345 GND.n2190 19.9241
R6382 GND.n4354 GND.n2179 19.9241
R6383 GND.n4431 GND.n2147 19.9241
R6384 GND.n4430 GND.n2149 19.9241
R6385 GND.n4362 GND.n2157 19.9241
R6386 GND.n4423 GND.n2159 19.9241
R6387 GND.n4420 GND.n4419 19.9241
R6388 GND.n4414 GND.n2164 19.9241
R6389 GND.n4413 GND.n4372 19.9241
R6390 GND.n4382 GND.n4380 19.9241
R6391 GND.n4406 GND.n4381 19.9241
R6392 GND.n4393 GND.n4387 19.9241
R6393 GND.n4441 GND.n2132 19.9241
R6394 GND.n4442 GND.n2128 19.9241
R6395 GND.n4446 GND.n2129 19.9241
R6396 GND.n4457 GND.n2119 19.9241
R6397 GND.n4456 GND.n2120 19.9241
R6398 GND.n4467 GND.n2110 19.9241
R6399 GND.n4468 GND.n2104 19.9241
R6400 GND.n4472 GND.n2107 19.9241
R6401 GND.n4483 GND.n2094 19.9241
R6402 GND.n4493 GND.n2087 19.9241
R6403 GND.n4496 GND.n2084 19.9241
R6404 GND.n4501 GND.n2085 19.9241
R6405 GND.n4512 GND.n2075 19.9241
R6406 GND.n4511 GND.n2076 19.9241
R6407 GND.n4538 GND.n2068 19.9241
R6408 GND.n4539 GND.n2062 19.9241
R6409 GND.n4543 GND.n2064 19.9241
R6410 GND.n2063 GND.n2055 19.9241
R6411 GND.n4551 GND.n2053 19.9241
R6412 GND.n4554 GND.n79 19.9241
R6413 GND.n6502 GND.n81 19.9241
R6414 GND.n3566 GND.t68 19.8005
R6415 GND.n3566 GND.t116 19.8005
R6416 GND.n2322 GND.t75 19.8005
R6417 GND.n2322 GND.t100 19.8005
R6418 GND.n5265 GND.n5264 19.6128
R6419 GND.n6444 GND.n6419 19.6128
R6420 GND.n2048 GND.n2047 19.3944
R6421 GND.n2047 GND.n2046 19.3944
R6422 GND.n2046 GND.n2002 19.3944
R6423 GND.n2042 GND.n2002 19.3944
R6424 GND.n2042 GND.n2041 19.3944
R6425 GND.n2041 GND.n2040 19.3944
R6426 GND.n2040 GND.n2008 19.3944
R6427 GND.n2036 GND.n2008 19.3944
R6428 GND.n2036 GND.n2035 19.3944
R6429 GND.n2035 GND.n2034 19.3944
R6430 GND.n2034 GND.n2014 19.3944
R6431 GND.n2030 GND.n2014 19.3944
R6432 GND.n2030 GND.n2029 19.3944
R6433 GND.n2029 GND.n2028 19.3944
R6434 GND.n2436 GND.n1898 19.3944
R6435 GND.n4631 GND.n1898 19.3944
R6436 GND.n4631 GND.n1899 19.3944
R6437 GND.n1906 GND.n1899 19.3944
R6438 GND.n1907 GND.n1906 19.3944
R6439 GND.n1908 GND.n1907 19.3944
R6440 GND.n4291 GND.n1908 19.3944
R6441 GND.n4291 GND.n1914 19.3944
R6442 GND.n1915 GND.n1914 19.3944
R6443 GND.n1916 GND.n1915 19.3944
R6444 GND.n4318 GND.n1916 19.3944
R6445 GND.n4318 GND.n1922 19.3944
R6446 GND.n1923 GND.n1922 19.3944
R6447 GND.n1924 GND.n1923 19.3944
R6448 GND.n2192 GND.n1924 19.3944
R6449 GND.n2192 GND.n1930 19.3944
R6450 GND.n1931 GND.n1930 19.3944
R6451 GND.n1932 GND.n1931 19.3944
R6452 GND.n2180 GND.n1932 19.3944
R6453 GND.n2180 GND.n1938 19.3944
R6454 GND.n1939 GND.n1938 19.3944
R6455 GND.n1940 GND.n1939 19.3944
R6456 GND.n2162 GND.n1940 19.3944
R6457 GND.n2162 GND.n1946 19.3944
R6458 GND.n1947 GND.n1946 19.3944
R6459 GND.n1948 GND.n1947 19.3944
R6460 GND.n4404 GND.n1948 19.3944
R6461 GND.n4404 GND.n1954 19.3944
R6462 GND.n1955 GND.n1954 19.3944
R6463 GND.n1956 GND.n1955 19.3944
R6464 GND.n2131 GND.n1956 19.3944
R6465 GND.n2131 GND.n1962 19.3944
R6466 GND.n1963 GND.n1962 19.3944
R6467 GND.n1964 GND.n1963 19.3944
R6468 GND.n2108 GND.n1964 19.3944
R6469 GND.n2108 GND.n1970 19.3944
R6470 GND.n1971 GND.n1970 19.3944
R6471 GND.n1972 GND.n1971 19.3944
R6472 GND.n2096 GND.n1972 19.3944
R6473 GND.n2096 GND.n1978 19.3944
R6474 GND.n1979 GND.n1978 19.3944
R6475 GND.n1980 GND.n1979 19.3944
R6476 GND.n4498 GND.n1980 19.3944
R6477 GND.n4498 GND.n1986 19.3944
R6478 GND.n1987 GND.n1986 19.3944
R6479 GND.n1988 GND.n1987 19.3944
R6480 GND.n4541 GND.n1988 19.3944
R6481 GND.n4541 GND.n1994 19.3944
R6482 GND.n1995 GND.n1994 19.3944
R6483 GND.n1996 GND.n1995 19.3944
R6484 GND.n1997 GND.n1996 19.3944
R6485 GND.n2437 GND.n1902 19.3944
R6486 GND.n4629 GND.n1902 19.3944
R6487 GND.n4629 GND.n4628 19.3944
R6488 GND.n4628 GND.n4627 19.3944
R6489 GND.n4627 GND.n1905 19.3944
R6490 GND.n4623 GND.n1905 19.3944
R6491 GND.n4623 GND.n4622 19.3944
R6492 GND.n4622 GND.n4621 19.3944
R6493 GND.n4621 GND.n1913 19.3944
R6494 GND.n4617 GND.n1913 19.3944
R6495 GND.n4617 GND.n4616 19.3944
R6496 GND.n4616 GND.n4615 19.3944
R6497 GND.n4615 GND.n1921 19.3944
R6498 GND.n4611 GND.n1921 19.3944
R6499 GND.n4611 GND.n4610 19.3944
R6500 GND.n4610 GND.n4609 19.3944
R6501 GND.n4609 GND.n1929 19.3944
R6502 GND.n4605 GND.n1929 19.3944
R6503 GND.n4605 GND.n4604 19.3944
R6504 GND.n4604 GND.n4603 19.3944
R6505 GND.n4603 GND.n1937 19.3944
R6506 GND.n4599 GND.n1937 19.3944
R6507 GND.n4599 GND.n4598 19.3944
R6508 GND.n4598 GND.n4597 19.3944
R6509 GND.n4597 GND.n1945 19.3944
R6510 GND.n4593 GND.n1945 19.3944
R6511 GND.n4593 GND.n4592 19.3944
R6512 GND.n4592 GND.n4591 19.3944
R6513 GND.n4591 GND.n1953 19.3944
R6514 GND.n4587 GND.n1953 19.3944
R6515 GND.n4587 GND.n4586 19.3944
R6516 GND.n4586 GND.n4585 19.3944
R6517 GND.n4585 GND.n1961 19.3944
R6518 GND.n4581 GND.n1961 19.3944
R6519 GND.n4581 GND.n4580 19.3944
R6520 GND.n4580 GND.n4579 19.3944
R6521 GND.n4579 GND.n1969 19.3944
R6522 GND.n4575 GND.n1969 19.3944
R6523 GND.n4575 GND.n4574 19.3944
R6524 GND.n4574 GND.n4573 19.3944
R6525 GND.n4573 GND.n1977 19.3944
R6526 GND.n4569 GND.n1977 19.3944
R6527 GND.n4569 GND.n4568 19.3944
R6528 GND.n4568 GND.n4567 19.3944
R6529 GND.n4567 GND.n1985 19.3944
R6530 GND.n4563 GND.n1985 19.3944
R6531 GND.n4563 GND.n4562 19.3944
R6532 GND.n4562 GND.n4561 19.3944
R6533 GND.n4561 GND.n1993 19.3944
R6534 GND.n4557 GND.n1993 19.3944
R6535 GND.n4557 GND.n4556 19.3944
R6536 GND.n6497 GND.n6496 19.3944
R6537 GND.n6496 GND.n6495 19.3944
R6538 GND.n6495 GND.n90 19.3944
R6539 GND.n6491 GND.n90 19.3944
R6540 GND.n6491 GND.n6490 19.3944
R6541 GND.n6490 GND.n6489 19.3944
R6542 GND.n6489 GND.n95 19.3944
R6543 GND.n6485 GND.n95 19.3944
R6544 GND.n6485 GND.n6484 19.3944
R6545 GND.n6484 GND.n6483 19.3944
R6546 GND.n6483 GND.n100 19.3944
R6547 GND.n6479 GND.n100 19.3944
R6548 GND.n6479 GND.n6478 19.3944
R6549 GND.n6478 GND.n6477 19.3944
R6550 GND.n6477 GND.n105 19.3944
R6551 GND.n6473 GND.n6472 19.3944
R6552 GND.n6472 GND.n6471 19.3944
R6553 GND.n6471 GND.n113 19.3944
R6554 GND.n6467 GND.n113 19.3944
R6555 GND.n6467 GND.n6466 19.3944
R6556 GND.n6466 GND.n6465 19.3944
R6557 GND.n6465 GND.n118 19.3944
R6558 GND.n6461 GND.n118 19.3944
R6559 GND.n6461 GND.n6460 19.3944
R6560 GND.n6460 GND.n6459 19.3944
R6561 GND.n6459 GND.n123 19.3944
R6562 GND.n6455 GND.n123 19.3944
R6563 GND.n6455 GND.n6454 19.3944
R6564 GND.n6454 GND.n6453 19.3944
R6565 GND.n6453 GND.n128 19.3944
R6566 GND.n6449 GND.n128 19.3944
R6567 GND.n1066 GND.n1063 19.3944
R6568 GND.n1066 GND.n1061 19.3944
R6569 GND.n1073 GND.n1061 19.3944
R6570 GND.n1074 GND.n1073 19.3944
R6571 GND.n5170 GND.n1074 19.3944
R6572 GND.n5170 GND.n5169 19.3944
R6573 GND.n5169 GND.n5168 19.3944
R6574 GND.n5168 GND.n1077 19.3944
R6575 GND.n5164 GND.n1077 19.3944
R6576 GND.n5164 GND.n5163 19.3944
R6577 GND.n5163 GND.n5162 19.3944
R6578 GND.n5162 GND.n1085 19.3944
R6579 GND.n5158 GND.n1085 19.3944
R6580 GND.n5158 GND.n5157 19.3944
R6581 GND.n5157 GND.n5156 19.3944
R6582 GND.n5156 GND.n1093 19.3944
R6583 GND.n5152 GND.n1093 19.3944
R6584 GND.n5152 GND.n5151 19.3944
R6585 GND.n5151 GND.n5150 19.3944
R6586 GND.n5150 GND.n1101 19.3944
R6587 GND.n5146 GND.n1101 19.3944
R6588 GND.n5146 GND.n5145 19.3944
R6589 GND.n5145 GND.n5144 19.3944
R6590 GND.n5144 GND.n1109 19.3944
R6591 GND.n5140 GND.n1109 19.3944
R6592 GND.n5140 GND.n5139 19.3944
R6593 GND.n5139 GND.n5138 19.3944
R6594 GND.n5138 GND.n1117 19.3944
R6595 GND.n5134 GND.n1117 19.3944
R6596 GND.n5134 GND.n5133 19.3944
R6597 GND.n5133 GND.n5132 19.3944
R6598 GND.n5132 GND.n1125 19.3944
R6599 GND.n5128 GND.n1125 19.3944
R6600 GND.n5128 GND.n5127 19.3944
R6601 GND.n5127 GND.n5126 19.3944
R6602 GND.n5126 GND.n1133 19.3944
R6603 GND.n5122 GND.n1133 19.3944
R6604 GND.n5122 GND.n5121 19.3944
R6605 GND.n5121 GND.n5120 19.3944
R6606 GND.n5120 GND.n1141 19.3944
R6607 GND.n5116 GND.n1141 19.3944
R6608 GND.n5116 GND.n5115 19.3944
R6609 GND.n5115 GND.n5114 19.3944
R6610 GND.n5114 GND.n1149 19.3944
R6611 GND.n5110 GND.n1149 19.3944
R6612 GND.n5110 GND.n5109 19.3944
R6613 GND.n5109 GND.n5108 19.3944
R6614 GND.n5108 GND.n1157 19.3944
R6615 GND.n5104 GND.n1157 19.3944
R6616 GND.n5104 GND.n5103 19.3944
R6617 GND.n5103 GND.n5102 19.3944
R6618 GND.n5095 GND.n5094 19.3944
R6619 GND.n5094 GND.n5093 19.3944
R6620 GND.n5093 GND.n1177 19.3944
R6621 GND.n5089 GND.n1177 19.3944
R6622 GND.n5089 GND.n5088 19.3944
R6623 GND.n5088 GND.n5087 19.3944
R6624 GND.n5087 GND.n1182 19.3944
R6625 GND.n5083 GND.n1182 19.3944
R6626 GND.n5083 GND.n5082 19.3944
R6627 GND.n5082 GND.n5081 19.3944
R6628 GND.n5081 GND.n1187 19.3944
R6629 GND.n5077 GND.n1187 19.3944
R6630 GND.n5077 GND.n5076 19.3944
R6631 GND.n5074 GND.n1197 19.3944
R6632 GND.n5070 GND.n1197 19.3944
R6633 GND.n5070 GND.n5069 19.3944
R6634 GND.n5069 GND.n5068 19.3944
R6635 GND.n5068 GND.n1202 19.3944
R6636 GND.n5064 GND.n1202 19.3944
R6637 GND.n5064 GND.n5063 19.3944
R6638 GND.n5063 GND.n5062 19.3944
R6639 GND.n5062 GND.n1207 19.3944
R6640 GND.n5058 GND.n1207 19.3944
R6641 GND.n5058 GND.n5057 19.3944
R6642 GND.n5057 GND.n5056 19.3944
R6643 GND.n5056 GND.n1212 19.3944
R6644 GND.n5052 GND.n1212 19.3944
R6645 GND.n5052 GND.n5051 19.3944
R6646 GND.n5051 GND.n5050 19.3944
R6647 GND.n3099 GND.n3049 19.3944
R6648 GND.n3103 GND.n3049 19.3944
R6649 GND.n3104 GND.n3103 19.3944
R6650 GND.n3109 GND.n3104 19.3944
R6651 GND.n3109 GND.n3047 19.3944
R6652 GND.n3113 GND.n3047 19.3944
R6653 GND.n3113 GND.n3041 19.3944
R6654 GND.n3154 GND.n3041 19.3944
R6655 GND.n3154 GND.n3038 19.3944
R6656 GND.n3164 GND.n3038 19.3944
R6657 GND.n3164 GND.n3039 19.3944
R6658 GND.n3160 GND.n3039 19.3944
R6659 GND.n3160 GND.n3159 19.3944
R6660 GND.n3159 GND.n3009 19.3944
R6661 GND.n3194 GND.n3009 19.3944
R6662 GND.n3194 GND.n3006 19.3944
R6663 GND.n3200 GND.n3006 19.3944
R6664 GND.n3200 GND.n3007 19.3944
R6665 GND.n3007 GND.n2981 19.3944
R6666 GND.n3231 GND.n2981 19.3944
R6667 GND.n3232 GND.n3231 19.3944
R6668 GND.n3232 GND.n2979 19.3944
R6669 GND.n3236 GND.n2979 19.3944
R6670 GND.n3242 GND.n3236 19.3944
R6671 GND.n3243 GND.n3242 19.3944
R6672 GND.n3243 GND.n2977 19.3944
R6673 GND.n3248 GND.n2977 19.3944
R6674 GND.n3248 GND.n2933 19.3944
R6675 GND.n3294 GND.n2933 19.3944
R6676 GND.n3294 GND.n2930 19.3944
R6677 GND.n3299 GND.n2930 19.3944
R6678 GND.n3299 GND.n2931 19.3944
R6679 GND.n2931 GND.n2905 19.3944
R6680 GND.n3384 GND.n2905 19.3944
R6681 GND.n3384 GND.n2902 19.3944
R6682 GND.n3389 GND.n2902 19.3944
R6683 GND.n3389 GND.n2903 19.3944
R6684 GND.n2903 GND.n2885 19.3944
R6685 GND.n3409 GND.n2885 19.3944
R6686 GND.n3409 GND.n2882 19.3944
R6687 GND.n3414 GND.n2882 19.3944
R6688 GND.n3414 GND.n2883 19.3944
R6689 GND.n2883 GND.n2863 19.3944
R6690 GND.n3434 GND.n2863 19.3944
R6691 GND.n3434 GND.n2860 19.3944
R6692 GND.n3445 GND.n2860 19.3944
R6693 GND.n3445 GND.n2861 19.3944
R6694 GND.n3441 GND.n2861 19.3944
R6695 GND.n3441 GND.n2843 19.3944
R6696 GND.n3465 GND.n2843 19.3944
R6697 GND.n3466 GND.n3465 19.3944
R6698 GND.n5043 GND.n5042 19.3944
R6699 GND.n5042 GND.n5041 19.3944
R6700 GND.n5041 GND.n1224 19.3944
R6701 GND.n5037 GND.n1224 19.3944
R6702 GND.n5037 GND.n5036 19.3944
R6703 GND.n5036 GND.n1228 19.3944
R6704 GND.n1282 GND.n1228 19.3944
R6705 GND.n1282 GND.n1253 19.3944
R6706 GND.n5024 GND.n1253 19.3944
R6707 GND.n5024 GND.n5023 19.3944
R6708 GND.n5023 GND.n1256 19.3944
R6709 GND.n5016 GND.n1256 19.3944
R6710 GND.n5016 GND.n5015 19.3944
R6711 GND.n5015 GND.n1264 19.3944
R6712 GND.n5191 GND.n1011 19.3944
R6713 GND.n3071 GND.n1011 19.3944
R6714 GND.n3072 GND.n3071 19.3944
R6715 GND.n3075 GND.n3072 19.3944
R6716 GND.n3075 GND.n3064 19.3944
R6717 GND.n3079 GND.n3064 19.3944
R6718 GND.n3080 GND.n3079 19.3944
R6719 GND.n3083 GND.n3080 19.3944
R6720 GND.n3083 GND.n3060 19.3944
R6721 GND.n3087 GND.n3060 19.3944
R6722 GND.n3088 GND.n3087 19.3944
R6723 GND.n3091 GND.n3088 19.3944
R6724 GND.n3091 GND.n3056 19.3944
R6725 GND.n3095 GND.n3056 19.3944
R6726 GND.n1068 GND.n1013 19.3944
R6727 GND.n1070 GND.n1068 19.3944
R6728 GND.n1071 GND.n1070 19.3944
R6729 GND.n1071 GND.n1057 19.3944
R6730 GND.n5172 GND.n1057 19.3944
R6731 GND.n5172 GND.n1058 19.3944
R6732 GND.n1078 GND.n1058 19.3944
R6733 GND.n1079 GND.n1078 19.3944
R6734 GND.n1080 GND.n1079 19.3944
R6735 GND.n3035 GND.n1080 19.3944
R6736 GND.n3035 GND.n1086 19.3944
R6737 GND.n1087 GND.n1086 19.3944
R6738 GND.n1088 GND.n1087 19.3944
R6739 GND.n3022 GND.n1088 19.3944
R6740 GND.n3022 GND.n1094 19.3944
R6741 GND.n1095 GND.n1094 19.3944
R6742 GND.n1096 GND.n1095 19.3944
R6743 GND.n2993 GND.n1096 19.3944
R6744 GND.n2993 GND.n1102 19.3944
R6745 GND.n1103 GND.n1102 19.3944
R6746 GND.n1104 GND.n1103 19.3944
R6747 GND.n2956 GND.n1104 19.3944
R6748 GND.n2956 GND.n1110 19.3944
R6749 GND.n1111 GND.n1110 19.3944
R6750 GND.n1112 GND.n1111 19.3944
R6751 GND.n3265 GND.n1112 19.3944
R6752 GND.n3265 GND.n1118 19.3944
R6753 GND.n1119 GND.n1118 19.3944
R6754 GND.n1120 GND.n1119 19.3944
R6755 GND.n2937 GND.n1120 19.3944
R6756 GND.n2937 GND.n1126 19.3944
R6757 GND.n1127 GND.n1126 19.3944
R6758 GND.n1128 GND.n1127 19.3944
R6759 GND.n2908 GND.n1128 19.3944
R6760 GND.n2908 GND.n1134 19.3944
R6761 GND.n1135 GND.n1134 19.3944
R6762 GND.n1136 GND.n1135 19.3944
R6763 GND.n3393 GND.n1136 19.3944
R6764 GND.n3393 GND.n1142 19.3944
R6765 GND.n1143 GND.n1142 19.3944
R6766 GND.n1144 GND.n1143 19.3944
R6767 GND.n3420 GND.n1144 19.3944
R6768 GND.n3420 GND.n1150 19.3944
R6769 GND.n1151 GND.n1150 19.3944
R6770 GND.n1152 GND.n1151 19.3944
R6771 GND.n2857 GND.n1152 19.3944
R6772 GND.n2857 GND.n1158 19.3944
R6773 GND.n1159 GND.n1158 19.3944
R6774 GND.n1160 GND.n1159 19.3944
R6775 GND.n3461 GND.n1160 19.3944
R6776 GND.n3461 GND.n3460 19.3944
R6777 GND.n3520 GND.n3519 19.3944
R6778 GND.n3523 GND.n3520 19.3944
R6779 GND.n3523 GND.n2830 19.3944
R6780 GND.n3527 GND.n2830 19.3944
R6781 GND.n3530 GND.n3527 19.3944
R6782 GND.n3531 GND.n3530 19.3944
R6783 GND.n3531 GND.n2828 19.3944
R6784 GND.n3535 GND.n2828 19.3944
R6785 GND.n3536 GND.n3535 19.3944
R6786 GND.n3539 GND.n3536 19.3944
R6787 GND.n3539 GND.n2822 19.3944
R6788 GND.n3543 GND.n2822 19.3944
R6789 GND.n3544 GND.n3543 19.3944
R6790 GND.n3547 GND.n3544 19.3944
R6791 GND.n3547 GND.n2820 19.3944
R6792 GND.n3551 GND.n2820 19.3944
R6793 GND.n3554 GND.n3551 19.3944
R6794 GND.n3555 GND.n3554 19.3944
R6795 GND.n3555 GND.n2818 19.3944
R6796 GND.n3559 GND.n2818 19.3944
R6797 GND.n3559 GND.n2711 19.3944
R6798 GND.n3658 GND.n2711 19.3944
R6799 GND.n3658 GND.n2709 19.3944
R6800 GND.n3662 GND.n2709 19.3944
R6801 GND.n3662 GND.n2705 19.3944
R6802 GND.n3705 GND.n2705 19.3944
R6803 GND.n3705 GND.n2703 19.3944
R6804 GND.n3709 GND.n2703 19.3944
R6805 GND.n3709 GND.n2697 19.3944
R6806 GND.n3741 GND.n2697 19.3944
R6807 GND.n3741 GND.n2698 19.3944
R6808 GND.n3737 GND.n2698 19.3944
R6809 GND.n3737 GND.n3736 19.3944
R6810 GND.n3736 GND.n3735 19.3944
R6811 GND.n3735 GND.n3729 19.3944
R6812 GND.n3731 GND.n3729 19.3944
R6813 GND.n3731 GND.n2673 19.3944
R6814 GND.n3794 GND.n2673 19.3944
R6815 GND.n3794 GND.n2670 19.3944
R6816 GND.n3807 GND.n2670 19.3944
R6817 GND.n3807 GND.n2671 19.3944
R6818 GND.n3803 GND.n2671 19.3944
R6819 GND.n3803 GND.n3802 19.3944
R6820 GND.n3802 GND.n2662 19.3944
R6821 GND.n2662 GND.n2661 19.3944
R6822 GND.n3842 GND.n2661 19.3944
R6823 GND.n3842 GND.n2658 19.3944
R6824 GND.n3850 GND.n2658 19.3944
R6825 GND.n3850 GND.n2659 19.3944
R6826 GND.n3846 GND.n2659 19.3944
R6827 GND.n3846 GND.n2649 19.3944
R6828 GND.n3878 GND.n2649 19.3944
R6829 GND.n3878 GND.n2646 19.3944
R6830 GND.n3903 GND.n2646 19.3944
R6831 GND.n3903 GND.n2647 19.3944
R6832 GND.n3899 GND.n2647 19.3944
R6833 GND.n3899 GND.n3898 19.3944
R6834 GND.n3898 GND.n3897 19.3944
R6835 GND.n3897 GND.n3886 19.3944
R6836 GND.n3893 GND.n3886 19.3944
R6837 GND.n3893 GND.n3892 19.3944
R6838 GND.n3892 GND.n3891 19.3944
R6839 GND.n3891 GND.n2633 19.3944
R6840 GND.n2633 GND.n2632 19.3944
R6841 GND.n3967 GND.n2632 19.3944
R6842 GND.n3967 GND.n2629 19.3944
R6843 GND.n3971 GND.n2629 19.3944
R6844 GND.n3972 GND.n3971 19.3944
R6845 GND.n3974 GND.n3972 19.3944
R6846 GND.n3974 GND.n2627 19.3944
R6847 GND.n3978 GND.n2627 19.3944
R6848 GND.n3978 GND.n2611 19.3944
R6849 GND.n4000 GND.n2611 19.3944
R6850 GND.n4000 GND.n2609 19.3944
R6851 GND.n4005 GND.n2609 19.3944
R6852 GND.n4005 GND.n2301 19.3944
R6853 GND.n4145 GND.n2301 19.3944
R6854 GND.n4146 GND.n4145 19.3944
R6855 GND.n4146 GND.n2295 19.3944
R6856 GND.n4150 GND.n2295 19.3944
R6857 GND.n4151 GND.n4150 19.3944
R6858 GND.n4154 GND.n4151 19.3944
R6859 GND.n4154 GND.n2293 19.3944
R6860 GND.n4158 GND.n2293 19.3944
R6861 GND.n4161 GND.n4158 19.3944
R6862 GND.n4162 GND.n4161 19.3944
R6863 GND.n4162 GND.n2291 19.3944
R6864 GND.n4166 GND.n2291 19.3944
R6865 GND.n4167 GND.n4166 19.3944
R6866 GND.n4170 GND.n4167 19.3944
R6867 GND.n4170 GND.n2284 19.3944
R6868 GND.n4174 GND.n2284 19.3944
R6869 GND.n4175 GND.n4174 19.3944
R6870 GND.n4178 GND.n4175 19.3944
R6871 GND.n4178 GND.n2282 19.3944
R6872 GND.n4182 GND.n2282 19.3944
R6873 GND.n4185 GND.n4182 19.3944
R6874 GND.n4186 GND.n4185 19.3944
R6875 GND.n2524 GND.n2523 19.3944
R6876 GND.n2523 GND.n2450 19.3944
R6877 GND.n2516 GND.n2450 19.3944
R6878 GND.n2516 GND.n2515 19.3944
R6879 GND.n2515 GND.n2466 19.3944
R6880 GND.n2508 GND.n2466 19.3944
R6881 GND.n2508 GND.n2507 19.3944
R6882 GND.n2507 GND.n2479 19.3944
R6883 GND.n2495 GND.n2479 19.3944
R6884 GND.n2495 GND.n2494 19.3944
R6885 GND.n2494 GND.n2249 19.3944
R6886 GND.n4215 GND.n2249 19.3944
R6887 GND.n4215 GND.n4214 19.3944
R6888 GND.n4214 GND.n4213 19.3944
R6889 GND.n4213 GND.n2254 19.3944
R6890 GND.n4209 GND.n2254 19.3944
R6891 GND.n4209 GND.n4208 19.3944
R6892 GND.n4208 GND.n4207 19.3944
R6893 GND.n4207 GND.n2262 19.3944
R6894 GND.n4203 GND.n2262 19.3944
R6895 GND.n4203 GND.n4202 19.3944
R6896 GND.n4202 GND.n4201 19.3944
R6897 GND.n4201 GND.n2270 19.3944
R6898 GND.n4197 GND.n2270 19.3944
R6899 GND.n4195 GND.n2280 19.3944
R6900 GND.n4191 GND.n2280 19.3944
R6901 GND.n3514 GND.n3511 19.3944
R6902 GND.n3516 GND.n3514 19.3944
R6903 GND.n5032 GND.n1230 19.3944
R6904 GND.n5027 GND.n1230 19.3944
R6905 GND.n5027 GND.n1249 19.3944
R6906 GND.n5020 GND.n1249 19.3944
R6907 GND.n5020 GND.n5019 19.3944
R6908 GND.n5019 GND.n1260 19.3944
R6909 GND.n5012 GND.n1260 19.3944
R6910 GND.n5012 GND.n5011 19.3944
R6911 GND.n5011 GND.n1270 19.3944
R6912 GND.n3469 GND.n1270 19.3944
R6913 GND.n3474 GND.n3469 19.3944
R6914 GND.n3477 GND.n3474 19.3944
R6915 GND.n3477 GND.n2841 19.3944
R6916 GND.n3481 GND.n2841 19.3944
R6917 GND.n3484 GND.n3481 19.3944
R6918 GND.n3487 GND.n3484 19.3944
R6919 GND.n3487 GND.n2839 19.3944
R6920 GND.n3491 GND.n2839 19.3944
R6921 GND.n3494 GND.n3491 19.3944
R6922 GND.n3497 GND.n3494 19.3944
R6923 GND.n3497 GND.n2837 19.3944
R6924 GND.n3501 GND.n2837 19.3944
R6925 GND.n3504 GND.n3501 19.3944
R6926 GND.n3507 GND.n3504 19.3944
R6927 GND.n4965 GND.n1305 19.3944
R6928 GND.n4965 GND.n4964 19.3944
R6929 GND.n4964 GND.n4963 19.3944
R6930 GND.n4963 GND.n1310 19.3944
R6931 GND.n1337 GND.n1310 19.3944
R6932 GND.n4951 GND.n1337 19.3944
R6933 GND.n4951 GND.n4950 19.3944
R6934 GND.n4950 GND.n4949 19.3944
R6935 GND.n4949 GND.n1343 19.3944
R6936 GND.n1364 GND.n1343 19.3944
R6937 GND.n4937 GND.n1364 19.3944
R6938 GND.n4937 GND.n4936 19.3944
R6939 GND.n4936 GND.n4935 19.3944
R6940 GND.n4935 GND.n1370 19.3944
R6941 GND.n1391 GND.n1370 19.3944
R6942 GND.n4923 GND.n1391 19.3944
R6943 GND.n4923 GND.n4922 19.3944
R6944 GND.n4922 GND.n4921 19.3944
R6945 GND.n4921 GND.n1397 19.3944
R6946 GND.n1417 GND.n1397 19.3944
R6947 GND.n4909 GND.n1417 19.3944
R6948 GND.n4909 GND.n4908 19.3944
R6949 GND.n4908 GND.n4907 19.3944
R6950 GND.n4907 GND.n1423 19.3944
R6951 GND.n4895 GND.n1423 19.3944
R6952 GND.n4895 GND.n4894 19.3944
R6953 GND.n4894 GND.n4893 19.3944
R6954 GND.n4893 GND.n1443 19.3944
R6955 GND.n4881 GND.n1443 19.3944
R6956 GND.n4881 GND.n4880 19.3944
R6957 GND.n4880 GND.n4879 19.3944
R6958 GND.n4879 GND.n1463 19.3944
R6959 GND.n4867 GND.n1463 19.3944
R6960 GND.n4867 GND.n4866 19.3944
R6961 GND.n4866 GND.n4865 19.3944
R6962 GND.n4865 GND.n1483 19.3944
R6963 GND.n4853 GND.n1483 19.3944
R6964 GND.n4853 GND.n4852 19.3944
R6965 GND.n4852 GND.n4851 19.3944
R6966 GND.n4851 GND.n1502 19.3944
R6967 GND.n4839 GND.n1502 19.3944
R6968 GND.n4839 GND.n4838 19.3944
R6969 GND.n4838 GND.n4837 19.3944
R6970 GND.n4837 GND.n1522 19.3944
R6971 GND.n1552 GND.n1522 19.3944
R6972 GND.n1552 GND.n1549 19.3944
R6973 GND.n4818 GND.n1549 19.3944
R6974 GND.n4818 GND.n4817 19.3944
R6975 GND.n4817 GND.n4816 19.3944
R6976 GND.n4816 GND.n1558 19.3944
R6977 GND.n1596 GND.n1558 19.3944
R6978 GND.n1596 GND.n1593 19.3944
R6979 GND.n4798 GND.n1593 19.3944
R6980 GND.n4798 GND.n4797 19.3944
R6981 GND.n4797 GND.n4796 19.3944
R6982 GND.n4796 GND.n1602 19.3944
R6983 GND.n1646 GND.n1602 19.3944
R6984 GND.n1649 GND.n1646 19.3944
R6985 GND.n1649 GND.n1643 19.3944
R6986 GND.n4770 GND.n1643 19.3944
R6987 GND.n4770 GND.n4769 19.3944
R6988 GND.n4769 GND.n4768 19.3944
R6989 GND.n4768 GND.n1655 19.3944
R6990 GND.n1690 GND.n1655 19.3944
R6991 GND.n1690 GND.n1687 19.3944
R6992 GND.n4750 GND.n1687 19.3944
R6993 GND.n4750 GND.n4749 19.3944
R6994 GND.n4749 GND.n4748 19.3944
R6995 GND.n4748 GND.n1696 19.3944
R6996 GND.n2623 GND.n1696 19.3944
R6997 GND.n2623 GND.n1730 19.3944
R6998 GND.n4729 GND.n1730 19.3944
R6999 GND.n4729 GND.n4728 19.3944
R7000 GND.n4728 GND.n4727 19.3944
R7001 GND.n4727 GND.n1734 19.3944
R7002 GND.n4715 GND.n1734 19.3944
R7003 GND.n4715 GND.n4714 19.3944
R7004 GND.n4714 GND.n4713 19.3944
R7005 GND.n4713 GND.n1754 19.3944
R7006 GND.n1771 GND.n1754 19.3944
R7007 GND.n4701 GND.n1771 19.3944
R7008 GND.n4701 GND.n4700 19.3944
R7009 GND.n4700 GND.n4699 19.3944
R7010 GND.n4699 GND.n1777 19.3944
R7011 GND.n1797 GND.n1777 19.3944
R7012 GND.n4687 GND.n1797 19.3944
R7013 GND.n4687 GND.n4686 19.3944
R7014 GND.n4686 GND.n4685 19.3944
R7015 GND.n4685 GND.n1803 19.3944
R7016 GND.n1824 GND.n1803 19.3944
R7017 GND.n4673 GND.n1824 19.3944
R7018 GND.n4673 GND.n4672 19.3944
R7019 GND.n4672 GND.n4671 19.3944
R7020 GND.n4671 GND.n1830 19.3944
R7021 GND.n1851 GND.n1830 19.3944
R7022 GND.n4659 GND.n1851 19.3944
R7023 GND.n4659 GND.n4658 19.3944
R7024 GND.n4658 GND.n4657 19.3944
R7025 GND.n6194 GND.n309 19.3944
R7026 GND.n6194 GND.n305 19.3944
R7027 GND.n6200 GND.n305 19.3944
R7028 GND.n6200 GND.n303 19.3944
R7029 GND.n6204 GND.n303 19.3944
R7030 GND.n6204 GND.n299 19.3944
R7031 GND.n6210 GND.n299 19.3944
R7032 GND.n6210 GND.n297 19.3944
R7033 GND.n6214 GND.n297 19.3944
R7034 GND.n6214 GND.n293 19.3944
R7035 GND.n6220 GND.n293 19.3944
R7036 GND.n6220 GND.n291 19.3944
R7037 GND.n6224 GND.n291 19.3944
R7038 GND.n6224 GND.n287 19.3944
R7039 GND.n6230 GND.n287 19.3944
R7040 GND.n6230 GND.n285 19.3944
R7041 GND.n6234 GND.n285 19.3944
R7042 GND.n6234 GND.n281 19.3944
R7043 GND.n6240 GND.n281 19.3944
R7044 GND.n6240 GND.n279 19.3944
R7045 GND.n6244 GND.n279 19.3944
R7046 GND.n6244 GND.n275 19.3944
R7047 GND.n6250 GND.n275 19.3944
R7048 GND.n6250 GND.n273 19.3944
R7049 GND.n6254 GND.n273 19.3944
R7050 GND.n6254 GND.n269 19.3944
R7051 GND.n6260 GND.n269 19.3944
R7052 GND.n6260 GND.n267 19.3944
R7053 GND.n6264 GND.n267 19.3944
R7054 GND.n6264 GND.n263 19.3944
R7055 GND.n6270 GND.n263 19.3944
R7056 GND.n6270 GND.n261 19.3944
R7057 GND.n6274 GND.n261 19.3944
R7058 GND.n6274 GND.n257 19.3944
R7059 GND.n6280 GND.n257 19.3944
R7060 GND.n6280 GND.n255 19.3944
R7061 GND.n6284 GND.n255 19.3944
R7062 GND.n6284 GND.n251 19.3944
R7063 GND.n6290 GND.n251 19.3944
R7064 GND.n6290 GND.n249 19.3944
R7065 GND.n6294 GND.n249 19.3944
R7066 GND.n6294 GND.n245 19.3944
R7067 GND.n6300 GND.n245 19.3944
R7068 GND.n6300 GND.n243 19.3944
R7069 GND.n6304 GND.n243 19.3944
R7070 GND.n6304 GND.n239 19.3944
R7071 GND.n6310 GND.n239 19.3944
R7072 GND.n6310 GND.n237 19.3944
R7073 GND.n6314 GND.n237 19.3944
R7074 GND.n6314 GND.n233 19.3944
R7075 GND.n6320 GND.n233 19.3944
R7076 GND.n6320 GND.n231 19.3944
R7077 GND.n6324 GND.n231 19.3944
R7078 GND.n6324 GND.n227 19.3944
R7079 GND.n6330 GND.n227 19.3944
R7080 GND.n6330 GND.n225 19.3944
R7081 GND.n6335 GND.n225 19.3944
R7082 GND.n6335 GND.n221 19.3944
R7083 GND.n6341 GND.n221 19.3944
R7084 GND.n6342 GND.n6341 19.3944
R7085 GND.n5464 GND.n747 19.3944
R7086 GND.n5464 GND.n743 19.3944
R7087 GND.n5470 GND.n743 19.3944
R7088 GND.n5470 GND.n741 19.3944
R7089 GND.n5474 GND.n741 19.3944
R7090 GND.n5474 GND.n737 19.3944
R7091 GND.n5480 GND.n737 19.3944
R7092 GND.n5480 GND.n735 19.3944
R7093 GND.n5484 GND.n735 19.3944
R7094 GND.n5484 GND.n731 19.3944
R7095 GND.n5490 GND.n731 19.3944
R7096 GND.n5490 GND.n729 19.3944
R7097 GND.n5494 GND.n729 19.3944
R7098 GND.n5494 GND.n725 19.3944
R7099 GND.n5500 GND.n725 19.3944
R7100 GND.n5500 GND.n723 19.3944
R7101 GND.n5504 GND.n723 19.3944
R7102 GND.n5504 GND.n719 19.3944
R7103 GND.n5510 GND.n719 19.3944
R7104 GND.n5510 GND.n717 19.3944
R7105 GND.n5514 GND.n717 19.3944
R7106 GND.n5514 GND.n713 19.3944
R7107 GND.n5520 GND.n713 19.3944
R7108 GND.n5520 GND.n711 19.3944
R7109 GND.n5524 GND.n711 19.3944
R7110 GND.n5524 GND.n707 19.3944
R7111 GND.n5530 GND.n707 19.3944
R7112 GND.n5530 GND.n705 19.3944
R7113 GND.n5534 GND.n705 19.3944
R7114 GND.n5534 GND.n701 19.3944
R7115 GND.n5540 GND.n701 19.3944
R7116 GND.n5540 GND.n699 19.3944
R7117 GND.n5544 GND.n699 19.3944
R7118 GND.n5544 GND.n695 19.3944
R7119 GND.n5550 GND.n695 19.3944
R7120 GND.n5550 GND.n693 19.3944
R7121 GND.n5554 GND.n693 19.3944
R7122 GND.n5554 GND.n689 19.3944
R7123 GND.n5560 GND.n689 19.3944
R7124 GND.n5560 GND.n687 19.3944
R7125 GND.n5564 GND.n687 19.3944
R7126 GND.n5564 GND.n683 19.3944
R7127 GND.n5570 GND.n683 19.3944
R7128 GND.n5570 GND.n681 19.3944
R7129 GND.n5574 GND.n681 19.3944
R7130 GND.n5574 GND.n677 19.3944
R7131 GND.n5580 GND.n677 19.3944
R7132 GND.n5580 GND.n675 19.3944
R7133 GND.n5584 GND.n675 19.3944
R7134 GND.n5584 GND.n671 19.3944
R7135 GND.n5590 GND.n671 19.3944
R7136 GND.n5590 GND.n669 19.3944
R7137 GND.n5594 GND.n669 19.3944
R7138 GND.n5594 GND.n665 19.3944
R7139 GND.n5600 GND.n665 19.3944
R7140 GND.n5600 GND.n663 19.3944
R7141 GND.n5604 GND.n663 19.3944
R7142 GND.n5604 GND.n659 19.3944
R7143 GND.n5610 GND.n659 19.3944
R7144 GND.n5610 GND.n657 19.3944
R7145 GND.n5614 GND.n657 19.3944
R7146 GND.n5614 GND.n653 19.3944
R7147 GND.n5620 GND.n653 19.3944
R7148 GND.n5620 GND.n651 19.3944
R7149 GND.n5624 GND.n651 19.3944
R7150 GND.n5624 GND.n647 19.3944
R7151 GND.n5630 GND.n647 19.3944
R7152 GND.n5630 GND.n645 19.3944
R7153 GND.n5634 GND.n645 19.3944
R7154 GND.n5634 GND.n641 19.3944
R7155 GND.n5640 GND.n641 19.3944
R7156 GND.n5640 GND.n639 19.3944
R7157 GND.n5644 GND.n639 19.3944
R7158 GND.n5644 GND.n635 19.3944
R7159 GND.n5650 GND.n635 19.3944
R7160 GND.n5650 GND.n633 19.3944
R7161 GND.n5654 GND.n633 19.3944
R7162 GND.n5654 GND.n629 19.3944
R7163 GND.n5660 GND.n629 19.3944
R7164 GND.n5660 GND.n627 19.3944
R7165 GND.n5664 GND.n627 19.3944
R7166 GND.n5664 GND.n623 19.3944
R7167 GND.n5670 GND.n623 19.3944
R7168 GND.n5670 GND.n621 19.3944
R7169 GND.n5674 GND.n621 19.3944
R7170 GND.n5674 GND.n617 19.3944
R7171 GND.n5680 GND.n617 19.3944
R7172 GND.n5680 GND.n615 19.3944
R7173 GND.n5684 GND.n615 19.3944
R7174 GND.n5684 GND.n611 19.3944
R7175 GND.n5690 GND.n611 19.3944
R7176 GND.n5690 GND.n609 19.3944
R7177 GND.n5694 GND.n609 19.3944
R7178 GND.n5694 GND.n605 19.3944
R7179 GND.n5700 GND.n605 19.3944
R7180 GND.n5700 GND.n603 19.3944
R7181 GND.n5704 GND.n603 19.3944
R7182 GND.n5704 GND.n599 19.3944
R7183 GND.n5710 GND.n599 19.3944
R7184 GND.n5710 GND.n597 19.3944
R7185 GND.n5714 GND.n597 19.3944
R7186 GND.n5714 GND.n593 19.3944
R7187 GND.n5720 GND.n593 19.3944
R7188 GND.n5720 GND.n591 19.3944
R7189 GND.n5724 GND.n591 19.3944
R7190 GND.n5724 GND.n587 19.3944
R7191 GND.n5730 GND.n587 19.3944
R7192 GND.n5730 GND.n585 19.3944
R7193 GND.n5734 GND.n585 19.3944
R7194 GND.n5734 GND.n581 19.3944
R7195 GND.n5740 GND.n581 19.3944
R7196 GND.n5740 GND.n579 19.3944
R7197 GND.n5744 GND.n579 19.3944
R7198 GND.n5744 GND.n575 19.3944
R7199 GND.n5750 GND.n575 19.3944
R7200 GND.n5750 GND.n573 19.3944
R7201 GND.n5754 GND.n573 19.3944
R7202 GND.n5754 GND.n569 19.3944
R7203 GND.n5760 GND.n569 19.3944
R7204 GND.n5760 GND.n567 19.3944
R7205 GND.n5764 GND.n567 19.3944
R7206 GND.n5764 GND.n563 19.3944
R7207 GND.n5770 GND.n563 19.3944
R7208 GND.n5770 GND.n561 19.3944
R7209 GND.n5774 GND.n561 19.3944
R7210 GND.n5774 GND.n557 19.3944
R7211 GND.n5780 GND.n557 19.3944
R7212 GND.n5780 GND.n555 19.3944
R7213 GND.n5784 GND.n555 19.3944
R7214 GND.n5784 GND.n551 19.3944
R7215 GND.n5790 GND.n551 19.3944
R7216 GND.n5790 GND.n549 19.3944
R7217 GND.n5794 GND.n549 19.3944
R7218 GND.n5794 GND.n545 19.3944
R7219 GND.n5800 GND.n545 19.3944
R7220 GND.n5800 GND.n543 19.3944
R7221 GND.n5804 GND.n543 19.3944
R7222 GND.n5804 GND.n539 19.3944
R7223 GND.n5810 GND.n539 19.3944
R7224 GND.n5810 GND.n537 19.3944
R7225 GND.n5814 GND.n537 19.3944
R7226 GND.n5814 GND.n533 19.3944
R7227 GND.n5820 GND.n533 19.3944
R7228 GND.n5820 GND.n531 19.3944
R7229 GND.n5824 GND.n531 19.3944
R7230 GND.n5824 GND.n527 19.3944
R7231 GND.n5830 GND.n527 19.3944
R7232 GND.n5830 GND.n525 19.3944
R7233 GND.n5834 GND.n525 19.3944
R7234 GND.n5834 GND.n521 19.3944
R7235 GND.n5840 GND.n521 19.3944
R7236 GND.n5840 GND.n519 19.3944
R7237 GND.n5844 GND.n519 19.3944
R7238 GND.n5844 GND.n515 19.3944
R7239 GND.n5850 GND.n515 19.3944
R7240 GND.n5850 GND.n513 19.3944
R7241 GND.n5854 GND.n513 19.3944
R7242 GND.n5854 GND.n509 19.3944
R7243 GND.n5860 GND.n509 19.3944
R7244 GND.n5860 GND.n507 19.3944
R7245 GND.n5864 GND.n507 19.3944
R7246 GND.n5864 GND.n503 19.3944
R7247 GND.n5870 GND.n503 19.3944
R7248 GND.n5870 GND.n501 19.3944
R7249 GND.n5874 GND.n501 19.3944
R7250 GND.n5874 GND.n497 19.3944
R7251 GND.n5880 GND.n497 19.3944
R7252 GND.n5880 GND.n495 19.3944
R7253 GND.n5884 GND.n495 19.3944
R7254 GND.n5884 GND.n491 19.3944
R7255 GND.n5890 GND.n491 19.3944
R7256 GND.n5890 GND.n489 19.3944
R7257 GND.n5894 GND.n489 19.3944
R7258 GND.n5894 GND.n485 19.3944
R7259 GND.n5900 GND.n485 19.3944
R7260 GND.n5900 GND.n483 19.3944
R7261 GND.n5904 GND.n483 19.3944
R7262 GND.n5904 GND.n479 19.3944
R7263 GND.n5910 GND.n479 19.3944
R7264 GND.n5910 GND.n477 19.3944
R7265 GND.n5914 GND.n477 19.3944
R7266 GND.n5914 GND.n473 19.3944
R7267 GND.n5920 GND.n473 19.3944
R7268 GND.n5920 GND.n471 19.3944
R7269 GND.n5924 GND.n471 19.3944
R7270 GND.n5924 GND.n467 19.3944
R7271 GND.n5930 GND.n467 19.3944
R7272 GND.n5930 GND.n465 19.3944
R7273 GND.n5934 GND.n465 19.3944
R7274 GND.n5934 GND.n461 19.3944
R7275 GND.n5940 GND.n461 19.3944
R7276 GND.n5940 GND.n459 19.3944
R7277 GND.n5944 GND.n459 19.3944
R7278 GND.n5944 GND.n455 19.3944
R7279 GND.n5950 GND.n455 19.3944
R7280 GND.n5950 GND.n453 19.3944
R7281 GND.n5954 GND.n453 19.3944
R7282 GND.n5954 GND.n449 19.3944
R7283 GND.n5960 GND.n449 19.3944
R7284 GND.n5960 GND.n447 19.3944
R7285 GND.n5964 GND.n447 19.3944
R7286 GND.n5964 GND.n443 19.3944
R7287 GND.n5970 GND.n443 19.3944
R7288 GND.n5970 GND.n441 19.3944
R7289 GND.n5974 GND.n441 19.3944
R7290 GND.n5974 GND.n437 19.3944
R7291 GND.n5980 GND.n437 19.3944
R7292 GND.n5980 GND.n435 19.3944
R7293 GND.n5984 GND.n435 19.3944
R7294 GND.n5984 GND.n431 19.3944
R7295 GND.n5990 GND.n431 19.3944
R7296 GND.n5990 GND.n429 19.3944
R7297 GND.n5994 GND.n429 19.3944
R7298 GND.n5994 GND.n425 19.3944
R7299 GND.n6000 GND.n425 19.3944
R7300 GND.n6000 GND.n423 19.3944
R7301 GND.n6004 GND.n423 19.3944
R7302 GND.n6004 GND.n419 19.3944
R7303 GND.n6010 GND.n419 19.3944
R7304 GND.n6010 GND.n417 19.3944
R7305 GND.n6014 GND.n417 19.3944
R7306 GND.n6014 GND.n413 19.3944
R7307 GND.n6020 GND.n413 19.3944
R7308 GND.n6020 GND.n411 19.3944
R7309 GND.n6024 GND.n411 19.3944
R7310 GND.n6024 GND.n407 19.3944
R7311 GND.n6030 GND.n407 19.3944
R7312 GND.n6030 GND.n405 19.3944
R7313 GND.n6034 GND.n405 19.3944
R7314 GND.n6034 GND.n401 19.3944
R7315 GND.n6040 GND.n401 19.3944
R7316 GND.n6040 GND.n399 19.3944
R7317 GND.n6044 GND.n399 19.3944
R7318 GND.n6044 GND.n395 19.3944
R7319 GND.n6050 GND.n395 19.3944
R7320 GND.n6050 GND.n393 19.3944
R7321 GND.n6054 GND.n393 19.3944
R7322 GND.n6054 GND.n389 19.3944
R7323 GND.n6060 GND.n389 19.3944
R7324 GND.n6060 GND.n387 19.3944
R7325 GND.n6064 GND.n387 19.3944
R7326 GND.n6064 GND.n383 19.3944
R7327 GND.n6070 GND.n383 19.3944
R7328 GND.n6070 GND.n381 19.3944
R7329 GND.n6074 GND.n381 19.3944
R7330 GND.n6074 GND.n377 19.3944
R7331 GND.n6080 GND.n377 19.3944
R7332 GND.n6080 GND.n375 19.3944
R7333 GND.n6084 GND.n375 19.3944
R7334 GND.n6084 GND.n371 19.3944
R7335 GND.n6090 GND.n371 19.3944
R7336 GND.n6090 GND.n369 19.3944
R7337 GND.n6094 GND.n369 19.3944
R7338 GND.n6094 GND.n365 19.3944
R7339 GND.n6100 GND.n365 19.3944
R7340 GND.n6100 GND.n363 19.3944
R7341 GND.n6104 GND.n363 19.3944
R7342 GND.n6104 GND.n359 19.3944
R7343 GND.n6110 GND.n359 19.3944
R7344 GND.n6110 GND.n357 19.3944
R7345 GND.n6114 GND.n357 19.3944
R7346 GND.n6114 GND.n353 19.3944
R7347 GND.n6120 GND.n353 19.3944
R7348 GND.n6120 GND.n351 19.3944
R7349 GND.n6124 GND.n351 19.3944
R7350 GND.n6124 GND.n347 19.3944
R7351 GND.n6130 GND.n347 19.3944
R7352 GND.n6130 GND.n345 19.3944
R7353 GND.n6134 GND.n345 19.3944
R7354 GND.n6134 GND.n341 19.3944
R7355 GND.n6140 GND.n341 19.3944
R7356 GND.n6140 GND.n339 19.3944
R7357 GND.n6144 GND.n339 19.3944
R7358 GND.n6144 GND.n335 19.3944
R7359 GND.n6150 GND.n335 19.3944
R7360 GND.n6150 GND.n333 19.3944
R7361 GND.n6154 GND.n333 19.3944
R7362 GND.n6154 GND.n329 19.3944
R7363 GND.n6160 GND.n329 19.3944
R7364 GND.n6160 GND.n327 19.3944
R7365 GND.n6164 GND.n327 19.3944
R7366 GND.n6164 GND.n323 19.3944
R7367 GND.n6170 GND.n323 19.3944
R7368 GND.n6170 GND.n321 19.3944
R7369 GND.n6174 GND.n321 19.3944
R7370 GND.n6174 GND.n317 19.3944
R7371 GND.n6180 GND.n317 19.3944
R7372 GND.n6180 GND.n315 19.3944
R7373 GND.n6184 GND.n315 19.3944
R7374 GND.n6184 GND.n311 19.3944
R7375 GND.n6190 GND.n311 19.3944
R7376 GND.n2369 GND.n2368 19.3944
R7377 GND.n2373 GND.n2368 19.3944
R7378 GND.n2373 GND.n2365 19.3944
R7379 GND.n2379 GND.n2365 19.3944
R7380 GND.n2379 GND.n2363 19.3944
R7381 GND.n2383 GND.n2363 19.3944
R7382 GND.n2383 GND.n2361 19.3944
R7383 GND.n2389 GND.n2361 19.3944
R7384 GND.n2389 GND.n2359 19.3944
R7385 GND.n2393 GND.n2359 19.3944
R7386 GND.n2393 GND.n2357 19.3944
R7387 GND.n2401 GND.n2357 19.3944
R7388 GND.n2401 GND.n2354 19.3944
R7389 GND.n2580 GND.n2408 19.3944
R7390 GND.n2574 GND.n2408 19.3944
R7391 GND.n2574 GND.n2573 19.3944
R7392 GND.n2573 GND.n2572 19.3944
R7393 GND.n2572 GND.n2414 19.3944
R7394 GND.n2566 GND.n2414 19.3944
R7395 GND.n2566 GND.n2565 19.3944
R7396 GND.n2565 GND.n2564 19.3944
R7397 GND.n2564 GND.n2420 19.3944
R7398 GND.n2558 GND.n2420 19.3944
R7399 GND.n2558 GND.n2557 19.3944
R7400 GND.n2557 GND.n2556 19.3944
R7401 GND.n2556 GND.n2426 19.3944
R7402 GND.n2550 GND.n2426 19.3944
R7403 GND.n2550 GND.n2549 19.3944
R7404 GND.n2549 GND.n2548 19.3944
R7405 GND.n4637 GND.n4636 19.3944
R7406 GND.n4636 GND.n4635 19.3944
R7407 GND.n4635 GND.n1890 19.3944
R7408 GND.n4224 GND.n1890 19.3944
R7409 GND.n4224 GND.n2231 19.3944
R7410 GND.n4297 GND.n2231 19.3944
R7411 GND.n4297 GND.n2229 19.3944
R7412 GND.n4303 GND.n2229 19.3944
R7413 GND.n4303 GND.n4302 19.3944
R7414 GND.n4302 GND.n2209 19.3944
R7415 GND.n4322 GND.n2209 19.3944
R7416 GND.n4322 GND.n2207 19.3944
R7417 GND.n4328 GND.n2207 19.3944
R7418 GND.n4328 GND.n4327 19.3944
R7419 GND.n4327 GND.n2186 19.3944
R7420 GND.n4347 GND.n2186 19.3944
R7421 GND.n4347 GND.n2184 19.3944
R7422 GND.n4352 GND.n2184 19.3944
R7423 GND.n4352 GND.n2153 19.3944
R7424 GND.n4428 GND.n2153 19.3944
R7425 GND.n4428 GND.n4427 19.3944
R7426 GND.n4425 GND.n2155 19.3944
R7427 GND.n4376 GND.n2155 19.3944
R7428 GND.n4411 GND.n4410 19.3944
R7429 GND.n4408 GND.n4378 19.3944
R7430 GND.n4391 GND.n4390 19.3944
R7431 GND.n4390 GND.n2126 19.3944
R7432 GND.n4448 GND.n2126 19.3944
R7433 GND.n4448 GND.n2124 19.3944
R7434 GND.n4454 GND.n2124 19.3944
R7435 GND.n4454 GND.n4453 19.3944
R7436 GND.n4453 GND.n2102 19.3944
R7437 GND.n4474 GND.n2102 19.3944
R7438 GND.n4474 GND.n2100 19.3944
R7439 GND.n4480 GND.n2100 19.3944
R7440 GND.n4480 GND.n4479 19.3944
R7441 GND.n4479 GND.n2082 19.3944
R7442 GND.n4503 GND.n2082 19.3944
R7443 GND.n4503 GND.n2080 19.3944
R7444 GND.n4509 GND.n2080 19.3944
R7445 GND.n4509 GND.n4508 19.3944
R7446 GND.n4508 GND.n2060 19.3944
R7447 GND.n4545 GND.n2060 19.3944
R7448 GND.n4545 GND.n2058 19.3944
R7449 GND.n4549 GND.n2058 19.3944
R7450 GND.n4549 GND.n85 19.3944
R7451 GND.n6500 GND.n85 19.3944
R7452 GND.n5334 GND.n871 19.3944
R7453 GND.n5334 GND.n5333 19.3944
R7454 GND.n5333 GND.n5332 19.3944
R7455 GND.n5332 GND.n876 19.3944
R7456 GND.n5326 GND.n876 19.3944
R7457 GND.n5326 GND.n5325 19.3944
R7458 GND.n5325 GND.n5324 19.3944
R7459 GND.n5324 GND.n884 19.3944
R7460 GND.n5318 GND.n884 19.3944
R7461 GND.n5318 GND.n5317 19.3944
R7462 GND.n5317 GND.n5316 19.3944
R7463 GND.n5316 GND.n892 19.3944
R7464 GND.n5310 GND.n892 19.3944
R7465 GND.n5310 GND.n5309 19.3944
R7466 GND.n5309 GND.n5308 19.3944
R7467 GND.n5308 GND.n900 19.3944
R7468 GND.n5302 GND.n900 19.3944
R7469 GND.n5302 GND.n5301 19.3944
R7470 GND.n5301 GND.n5300 19.3944
R7471 GND.n5300 GND.n908 19.3944
R7472 GND.n5294 GND.n908 19.3944
R7473 GND.n5294 GND.n5293 19.3944
R7474 GND.n5293 GND.n5292 19.3944
R7475 GND.n5292 GND.n916 19.3944
R7476 GND.n5286 GND.n916 19.3944
R7477 GND.n5286 GND.n5285 19.3944
R7478 GND.n5285 GND.n5284 19.3944
R7479 GND.n5284 GND.n924 19.3944
R7480 GND.n5278 GND.n924 19.3944
R7481 GND.n5278 GND.n5277 19.3944
R7482 GND.n5277 GND.n5276 19.3944
R7483 GND.n5276 GND.n932 19.3944
R7484 GND.n5270 GND.n932 19.3944
R7485 GND.n5270 GND.n5269 19.3944
R7486 GND.n5269 GND.n5268 19.3944
R7487 GND.n5268 GND.n940 19.3944
R7488 GND.n1024 GND.n940 19.3944
R7489 GND.n1024 GND.n1021 19.3944
R7490 GND.n5185 GND.n1021 19.3944
R7491 GND.n5185 GND.n5184 19.3944
R7492 GND.n5184 GND.n5183 19.3944
R7493 GND.n5183 GND.n1030 19.3944
R7494 GND.n3121 GND.n1030 19.3944
R7495 GND.n3121 GND.n3118 19.3944
R7496 GND.n3136 GND.n3118 19.3944
R7497 GND.n3136 GND.n3135 19.3944
R7498 GND.n3135 GND.n3134 19.3944
R7499 GND.n3134 GND.n3127 19.3944
R7500 GND.n3130 GND.n3127 19.3944
R7501 GND.n3130 GND.n3016 19.3944
R7502 GND.n3183 GND.n3016 19.3944
R7503 GND.n3183 GND.n3014 19.3944
R7504 GND.n3189 GND.n3014 19.3944
R7505 GND.n3189 GND.n3188 19.3944
R7506 GND.n3188 GND.n2988 19.3944
R7507 GND.n3218 GND.n2988 19.3944
R7508 GND.n3218 GND.n2986 19.3944
R7509 GND.n3225 GND.n2986 19.3944
R7510 GND.n3225 GND.n3224 19.3944
R7511 GND.n3224 GND.n3223 19.3944
R7512 GND.n3278 GND.n3277 19.3944
R7513 GND.n3275 GND.n2961 19.3944
R7514 GND.n3260 GND.n3255 19.3944
R7515 GND.n3258 GND.n3257 19.3944
R7516 GND.n3305 GND.n2926 19.3944
R7517 GND.n3305 GND.n2924 19.3944
R7518 GND.n3366 GND.n2924 19.3944
R7519 GND.n3366 GND.n3365 19.3944
R7520 GND.n3365 GND.n3364 19.3944
R7521 GND.n3364 GND.n3311 19.3944
R7522 GND.n3360 GND.n3311 19.3944
R7523 GND.n3360 GND.n3359 19.3944
R7524 GND.n3359 GND.n3358 19.3944
R7525 GND.n3358 GND.n3317 19.3944
R7526 GND.n3351 GND.n3317 19.3944
R7527 GND.n3351 GND.n3350 19.3944
R7528 GND.n3350 GND.n3349 19.3944
R7529 GND.n3349 GND.n3323 19.3944
R7530 GND.n3345 GND.n3323 19.3944
R7531 GND.n3345 GND.n3344 19.3944
R7532 GND.n3344 GND.n3343 19.3944
R7533 GND.n3343 GND.n3329 19.3944
R7534 GND.n3339 GND.n3329 19.3944
R7535 GND.n3339 GND.n3338 19.3944
R7536 GND.n3338 GND.n3337 19.3944
R7537 GND.n3337 GND.n1294 19.3944
R7538 GND.n4976 GND.n1294 19.3944
R7539 GND.n4976 GND.n4975 19.3944
R7540 GND.n4975 GND.n4974 19.3944
R7541 GND.n4974 GND.n1298 19.3944
R7542 GND.n1300 GND.n1298 19.3944
R7543 GND.n1321 GND.n1300 19.3944
R7544 GND.n1323 GND.n1321 19.3944
R7545 GND.n1323 GND.n1317 19.3944
R7546 GND.n4958 GND.n1317 19.3944
R7547 GND.n4958 GND.n4957 19.3944
R7548 GND.n4957 GND.n4956 19.3944
R7549 GND.n4956 GND.n1329 19.3944
R7550 GND.n1350 GND.n1329 19.3944
R7551 GND.n4944 GND.n1350 19.3944
R7552 GND.n4944 GND.n4943 19.3944
R7553 GND.n4943 GND.n4942 19.3944
R7554 GND.n4942 GND.n1356 19.3944
R7555 GND.n1377 GND.n1356 19.3944
R7556 GND.n4930 GND.n1377 19.3944
R7557 GND.n4930 GND.n4929 19.3944
R7558 GND.n4929 GND.n4928 19.3944
R7559 GND.n4928 GND.n1383 19.3944
R7560 GND.n1404 GND.n1383 19.3944
R7561 GND.n4916 GND.n1404 19.3944
R7562 GND.n4916 GND.n4915 19.3944
R7563 GND.n4915 GND.n4914 19.3944
R7564 GND.n4914 GND.n1410 19.3944
R7565 GND.n3684 GND.n1410 19.3944
R7566 GND.n3684 GND.n3681 19.3944
R7567 GND.n3688 GND.n3681 19.3944
R7568 GND.n3688 GND.n3679 19.3944
R7569 GND.n3700 GND.n3679 19.3944
R7570 GND.n3700 GND.n3699 19.3944
R7571 GND.n3699 GND.n3698 19.3944
R7572 GND.n3698 GND.n3696 19.3944
R7573 GND.n3696 GND.n2692 19.3944
R7574 GND.n2692 GND.n2690 19.3944
R7575 GND.n3748 GND.n2690 19.3944
R7576 GND.n3748 GND.n2688 19.3944
R7577 GND.n3752 GND.n2688 19.3944
R7578 GND.n3752 GND.n2680 19.3944
R7579 GND.n3773 GND.n2680 19.3944
R7580 GND.n3773 GND.n2678 19.3944
R7581 GND.n3786 GND.n2678 19.3944
R7582 GND.n3786 GND.n3785 19.3944
R7583 GND.n3785 GND.n3784 19.3944
R7584 GND.n3784 GND.n3781 19.3944
R7585 GND.n3781 GND.n1529 19.3944
R7586 GND.n4832 GND.n1529 19.3944
R7587 GND.n4832 GND.n4831 19.3944
R7588 GND.n4831 GND.n4830 19.3944
R7589 GND.n4830 GND.n1533 19.3944
R7590 GND.n1577 GND.n1533 19.3944
R7591 GND.n1580 GND.n1577 19.3944
R7592 GND.n1580 GND.n1574 19.3944
R7593 GND.n4805 GND.n1574 19.3944
R7594 GND.n4805 GND.n4804 19.3944
R7595 GND.n4804 GND.n4803 19.3944
R7596 GND.n4803 GND.n1586 19.3944
R7597 GND.n1621 GND.n1586 19.3944
R7598 GND.n1621 GND.n1618 19.3944
R7599 GND.n4784 GND.n1618 19.3944
R7600 GND.n4784 GND.n4783 19.3944
R7601 GND.n4783 GND.n4782 19.3944
R7602 GND.n4782 GND.n1627 19.3944
R7603 GND.n1665 GND.n1627 19.3944
R7604 GND.n1665 GND.n1662 19.3944
R7605 GND.n4763 GND.n1662 19.3944
R7606 GND.n4763 GND.n4762 19.3944
R7607 GND.n4762 GND.n4761 19.3944
R7608 GND.n4761 GND.n1671 19.3944
R7609 GND.n1714 GND.n1671 19.3944
R7610 GND.n1717 GND.n1714 19.3944
R7611 GND.n1717 GND.n1711 19.3944
R7612 GND.n4736 GND.n1711 19.3944
R7613 GND.n4736 GND.n4735 19.3944
R7614 GND.n4735 GND.n4734 19.3944
R7615 GND.n4734 GND.n1723 19.3944
R7616 GND.n2306 GND.n1723 19.3944
R7617 GND.n2309 GND.n2306 19.3944
R7618 GND.n2309 GND.n2303 19.3944
R7619 GND.n2314 GND.n2303 19.3944
R7620 GND.n2314 GND.n1760 19.3944
R7621 GND.n4708 GND.n1760 19.3944
R7622 GND.n4708 GND.n4707 19.3944
R7623 GND.n4707 GND.n4706 19.3944
R7624 GND.n4706 GND.n1764 19.3944
R7625 GND.n1784 GND.n1764 19.3944
R7626 GND.n4694 GND.n1784 19.3944
R7627 GND.n4694 GND.n4693 19.3944
R7628 GND.n4693 GND.n4692 19.3944
R7629 GND.n4692 GND.n1790 19.3944
R7630 GND.n1810 GND.n1790 19.3944
R7631 GND.n4680 GND.n1810 19.3944
R7632 GND.n4680 GND.n4679 19.3944
R7633 GND.n4679 GND.n4678 19.3944
R7634 GND.n4678 GND.n1816 19.3944
R7635 GND.n1837 GND.n1816 19.3944
R7636 GND.n4666 GND.n1837 19.3944
R7637 GND.n4666 GND.n4665 19.3944
R7638 GND.n4665 GND.n4664 19.3944
R7639 GND.n4664 GND.n1843 19.3944
R7640 GND.n1863 GND.n1843 19.3944
R7641 GND.n4652 GND.n1863 19.3944
R7642 GND.n4652 GND.n4651 19.3944
R7643 GND.n4651 GND.n4650 19.3944
R7644 GND.n4650 GND.n1869 19.3944
R7645 GND.n4644 GND.n1869 19.3944
R7646 GND.n4644 GND.n4643 19.3944
R7647 GND.n4643 GND.n4642 19.3944
R7648 GND.n4642 GND.n1878 19.3944
R7649 GND.n4232 GND.n1878 19.3944
R7650 GND.n4232 GND.n4229 19.3944
R7651 GND.n4277 GND.n4229 19.3944
R7652 GND.n4277 GND.n4276 19.3944
R7653 GND.n4276 GND.n4275 19.3944
R7654 GND.n4275 GND.n4238 19.3944
R7655 GND.n4271 GND.n4238 19.3944
R7656 GND.n4271 GND.n4270 19.3944
R7657 GND.n4270 GND.n4269 19.3944
R7658 GND.n4269 GND.n4244 19.3944
R7659 GND.n4265 GND.n4244 19.3944
R7660 GND.n4265 GND.n4264 19.3944
R7661 GND.n4264 GND.n4263 19.3944
R7662 GND.n4263 GND.n4250 19.3944
R7663 GND.n4259 GND.n4250 19.3944
R7664 GND.n4259 GND.n4258 19.3944
R7665 GND.n4258 GND.n4257 19.3944
R7666 GND.n4257 GND.n2143 19.3944
R7667 GND.n4433 GND.n2143 19.3944
R7668 GND.n4433 GND.n2144 19.3944
R7669 GND.n2167 GND.n2166 19.3944
R7670 GND.n4417 GND.n4416 19.3944
R7671 GND.n4395 GND.n4394 19.3944
R7672 GND.n4399 GND.n4398 19.3944
R7673 GND.n4439 GND.n2135 19.3944
R7674 GND.n4439 GND.n4438 19.3944
R7675 GND.n4438 GND.n2115 19.3944
R7676 GND.n4459 GND.n2115 19.3944
R7677 GND.n4459 GND.n2113 19.3944
R7678 GND.n4465 GND.n2113 19.3944
R7679 GND.n4465 GND.n4464 19.3944
R7680 GND.n4464 GND.n2092 19.3944
R7681 GND.n4485 GND.n2092 19.3944
R7682 GND.n4485 GND.n2090 19.3944
R7683 GND.n4491 GND.n2090 19.3944
R7684 GND.n4491 GND.n4490 19.3944
R7685 GND.n4490 GND.n2073 19.3944
R7686 GND.n4514 GND.n2073 19.3944
R7687 GND.n4514 GND.n2071 19.3944
R7688 GND.n4536 GND.n2071 19.3944
R7689 GND.n4536 GND.n4535 19.3944
R7690 GND.n4535 GND.n4534 19.3944
R7691 GND.n4534 GND.n4520 19.3944
R7692 GND.n4530 GND.n4520 19.3944
R7693 GND.n4530 GND.n4529 19.3944
R7694 GND.n4529 GND.n4528 19.3944
R7695 GND.n4528 GND.n147 19.3944
R7696 GND.n6417 GND.n147 19.3944
R7697 GND.n6417 GND.n6416 19.3944
R7698 GND.n6416 GND.n6415 19.3944
R7699 GND.n6415 GND.n151 19.3944
R7700 GND.n6409 GND.n151 19.3944
R7701 GND.n6409 GND.n6408 19.3944
R7702 GND.n6408 GND.n6407 19.3944
R7703 GND.n6407 GND.n159 19.3944
R7704 GND.n6401 GND.n159 19.3944
R7705 GND.n6401 GND.n6400 19.3944
R7706 GND.n6400 GND.n6399 19.3944
R7707 GND.n6399 GND.n167 19.3944
R7708 GND.n6393 GND.n167 19.3944
R7709 GND.n6393 GND.n6392 19.3944
R7710 GND.n6392 GND.n6391 19.3944
R7711 GND.n6391 GND.n175 19.3944
R7712 GND.n6385 GND.n175 19.3944
R7713 GND.n6385 GND.n6384 19.3944
R7714 GND.n6384 GND.n6383 19.3944
R7715 GND.n6383 GND.n183 19.3944
R7716 GND.n6377 GND.n183 19.3944
R7717 GND.n6377 GND.n6376 19.3944
R7718 GND.n6376 GND.n6375 19.3944
R7719 GND.n6375 GND.n191 19.3944
R7720 GND.n6369 GND.n191 19.3944
R7721 GND.n6369 GND.n6368 19.3944
R7722 GND.n6368 GND.n6367 19.3944
R7723 GND.n6367 GND.n199 19.3944
R7724 GND.n6361 GND.n199 19.3944
R7725 GND.n6361 GND.n6360 19.3944
R7726 GND.n6360 GND.n6359 19.3944
R7727 GND.n6359 GND.n207 19.3944
R7728 GND.n6353 GND.n207 19.3944
R7729 GND.n6353 GND.n6352 19.3944
R7730 GND.n6352 GND.n6351 19.3944
R7731 GND.n6351 GND.n215 19.3944
R7732 GND.n6345 GND.n215 19.3944
R7733 GND.n5261 GND.n5260 19.3944
R7734 GND.n5260 GND.n5259 19.3944
R7735 GND.n5259 GND.n5258 19.3944
R7736 GND.n5258 GND.n5256 19.3944
R7737 GND.n5256 GND.n5253 19.3944
R7738 GND.n5253 GND.n5252 19.3944
R7739 GND.n5252 GND.n5249 19.3944
R7740 GND.n5249 GND.n5248 19.3944
R7741 GND.n5248 GND.n5245 19.3944
R7742 GND.n5245 GND.n5244 19.3944
R7743 GND.n5244 GND.n5241 19.3944
R7744 GND.n5241 GND.n5240 19.3944
R7745 GND.n5240 GND.n5237 19.3944
R7746 GND.n5237 GND.n5236 19.3944
R7747 GND.n5236 GND.n5233 19.3944
R7748 GND.n5231 GND.n5228 19.3944
R7749 GND.n5228 GND.n5227 19.3944
R7750 GND.n5227 GND.n5224 19.3944
R7751 GND.n5224 GND.n5223 19.3944
R7752 GND.n5223 GND.n5220 19.3944
R7753 GND.n5220 GND.n5219 19.3944
R7754 GND.n5219 GND.n5216 19.3944
R7755 GND.n5216 GND.n5215 19.3944
R7756 GND.n5215 GND.n5212 19.3944
R7757 GND.n5212 GND.n5211 19.3944
R7758 GND.n5211 GND.n5208 19.3944
R7759 GND.n5208 GND.n5207 19.3944
R7760 GND.n5207 GND.n5204 19.3944
R7761 GND.n5204 GND.n5203 19.3944
R7762 GND.n5203 GND.n5200 19.3944
R7763 GND.n5200 GND.n5199 19.3944
R7764 GND.n1043 GND.n1041 19.3944
R7765 GND.n1043 GND.n1039 19.3944
R7766 GND.n5178 GND.n1039 19.3944
R7767 GND.n5178 GND.n5177 19.3944
R7768 GND.n5177 GND.n5176 19.3944
R7769 GND.n5176 GND.n1049 19.3944
R7770 GND.n3144 GND.n1049 19.3944
R7771 GND.n3150 GND.n3144 19.3944
R7772 GND.n3150 GND.n3149 19.3944
R7773 GND.n3149 GND.n3029 19.3944
R7774 GND.n3172 GND.n3029 19.3944
R7775 GND.n3172 GND.n3027 19.3944
R7776 GND.n3178 GND.n3027 19.3944
R7777 GND.n3178 GND.n3177 19.3944
R7778 GND.n3177 GND.n2999 19.3944
R7779 GND.n3207 GND.n2999 19.3944
R7780 GND.n3207 GND.n2997 19.3944
R7781 GND.n3213 GND.n2997 19.3944
R7782 GND.n3213 GND.n3212 19.3944
R7783 GND.n3212 GND.n2948 19.3944
R7784 GND.n3286 GND.n2948 19.3944
R7785 GND.n2947 GND.n2946 19.3944
R7786 GND.n2969 GND.n2946 19.3944
R7787 GND.n3270 GND.n3269 19.3944
R7788 GND.n2972 GND.n2971 19.3944
R7789 GND.n3290 GND.n3289 19.3944
R7790 GND.n3289 GND.n2915 19.3944
R7791 GND.n3374 GND.n2915 19.3944
R7792 GND.n3374 GND.n2913 19.3944
R7793 GND.n3380 GND.n2913 19.3944
R7794 GND.n3380 GND.n3379 19.3944
R7795 GND.n3379 GND.n2893 19.3944
R7796 GND.n3399 GND.n2893 19.3944
R7797 GND.n3399 GND.n2891 19.3944
R7798 GND.n3405 GND.n2891 19.3944
R7799 GND.n3405 GND.n3404 19.3944
R7800 GND.n3404 GND.n2874 19.3944
R7801 GND.n3424 GND.n2874 19.3944
R7802 GND.n3424 GND.n2872 19.3944
R7803 GND.n3430 GND.n2872 19.3944
R7804 GND.n3430 GND.n3429 19.3944
R7805 GND.n3429 GND.n2851 19.3944
R7806 GND.n3452 GND.n2851 19.3944
R7807 GND.n3452 GND.n2849 19.3944
R7808 GND.n3456 GND.n2849 19.3944
R7809 GND.n3456 GND.n1172 19.3944
R7810 GND.n5098 GND.n1172 19.3944
R7811 GND.n5460 GND.n749 19.3944
R7812 GND.n5454 GND.n749 19.3944
R7813 GND.n5454 GND.n5453 19.3944
R7814 GND.n5453 GND.n5452 19.3944
R7815 GND.n5452 GND.n756 19.3944
R7816 GND.n5446 GND.n756 19.3944
R7817 GND.n5446 GND.n5445 19.3944
R7818 GND.n5445 GND.n5444 19.3944
R7819 GND.n5444 GND.n764 19.3944
R7820 GND.n5438 GND.n764 19.3944
R7821 GND.n5438 GND.n5437 19.3944
R7822 GND.n5437 GND.n5436 19.3944
R7823 GND.n5436 GND.n772 19.3944
R7824 GND.n5430 GND.n772 19.3944
R7825 GND.n5430 GND.n5429 19.3944
R7826 GND.n5429 GND.n5428 19.3944
R7827 GND.n5428 GND.n780 19.3944
R7828 GND.n5422 GND.n780 19.3944
R7829 GND.n5422 GND.n5421 19.3944
R7830 GND.n5421 GND.n5420 19.3944
R7831 GND.n5420 GND.n788 19.3944
R7832 GND.n5414 GND.n788 19.3944
R7833 GND.n5414 GND.n5413 19.3944
R7834 GND.n5413 GND.n5412 19.3944
R7835 GND.n5412 GND.n796 19.3944
R7836 GND.n5406 GND.n796 19.3944
R7837 GND.n5406 GND.n5405 19.3944
R7838 GND.n5405 GND.n5404 19.3944
R7839 GND.n5404 GND.n804 19.3944
R7840 GND.n5398 GND.n804 19.3944
R7841 GND.n5398 GND.n5397 19.3944
R7842 GND.n5397 GND.n5396 19.3944
R7843 GND.n5396 GND.n812 19.3944
R7844 GND.n5390 GND.n812 19.3944
R7845 GND.n5390 GND.n5389 19.3944
R7846 GND.n5389 GND.n5388 19.3944
R7847 GND.n5388 GND.n820 19.3944
R7848 GND.n5382 GND.n820 19.3944
R7849 GND.n5382 GND.n5381 19.3944
R7850 GND.n5381 GND.n5380 19.3944
R7851 GND.n5380 GND.n828 19.3944
R7852 GND.n5374 GND.n828 19.3944
R7853 GND.n5374 GND.n5373 19.3944
R7854 GND.n5373 GND.n5372 19.3944
R7855 GND.n5372 GND.n836 19.3944
R7856 GND.n5366 GND.n836 19.3944
R7857 GND.n5366 GND.n5365 19.3944
R7858 GND.n5365 GND.n5364 19.3944
R7859 GND.n5364 GND.n844 19.3944
R7860 GND.n5358 GND.n844 19.3944
R7861 GND.n5358 GND.n5357 19.3944
R7862 GND.n5357 GND.n5356 19.3944
R7863 GND.n5356 GND.n852 19.3944
R7864 GND.n5350 GND.n852 19.3944
R7865 GND.n5350 GND.n5349 19.3944
R7866 GND.n5349 GND.n5348 19.3944
R7867 GND.n5348 GND.n860 19.3944
R7868 GND.n5342 GND.n860 19.3944
R7869 GND.n5342 GND.n5341 19.3944
R7870 GND.n5341 GND.n5340 19.3944
R7871 GND.n2538 GND.n2440 19.3944
R7872 GND.n2533 GND.n2440 19.3944
R7873 GND.n2533 GND.n2442 19.3944
R7874 GND.n2529 GND.n2442 19.3944
R7875 GND.n2529 GND.n2528 19.3944
R7876 GND.n2528 GND.n2447 19.3944
R7877 GND.n2452 GND.n2447 19.3944
R7878 GND.n2520 GND.n2452 19.3944
R7879 GND.n2520 GND.n2519 19.3944
R7880 GND.n2519 GND.n2459 19.3944
R7881 GND.n2512 GND.n2459 19.3944
R7882 GND.n2512 GND.n2511 19.3944
R7883 GND.n2511 GND.n2473 19.3944
R7884 GND.n2504 GND.n2473 19.3944
R7885 GND.n4220 GND.n2243 19.3944
R7886 GND.n4221 GND.n4220 19.3944
R7887 GND.n4282 GND.n4221 19.3944
R7888 GND.n4282 GND.n2240 19.3944
R7889 GND.n4287 GND.n2240 19.3944
R7890 GND.n4287 GND.n2241 19.3944
R7891 GND.n2241 GND.n2220 19.3944
R7892 GND.n4307 GND.n2220 19.3944
R7893 GND.n4307 GND.n2217 19.3944
R7894 GND.n4312 GND.n2217 19.3944
R7895 GND.n4312 GND.n2218 19.3944
R7896 GND.n2218 GND.n2198 19.3944
R7897 GND.n4332 GND.n2198 19.3944
R7898 GND.n4332 GND.n2195 19.3944
R7899 GND.n4337 GND.n2195 19.3944
R7900 GND.n4337 GND.n2196 19.3944
R7901 GND.n2196 GND.n2175 19.3944
R7902 GND.n4356 GND.n2175 19.3944
R7903 GND.n4356 GND.n2173 19.3944
R7904 GND.n4360 GND.n2173 19.3944
R7905 GND.n4364 GND.n4360 19.3944
R7906 GND.n4365 GND.n4364 19.3944
R7907 GND.n4365 GND.n2171 19.3944
R7908 GND.n4369 GND.n2171 19.3944
R7909 GND.n4369 GND.n46 19.3944
R7910 GND.n6541 GND.n46 19.3944
R7911 GND.n6541 GND.n6540 19.3944
R7912 GND.n6540 GND.n6539 19.3944
R7913 GND.n6539 GND.n50 19.3944
R7914 GND.n6535 GND.n50 19.3944
R7915 GND.n6535 GND.n6534 19.3944
R7916 GND.n6534 GND.n6533 19.3944
R7917 GND.n6533 GND.n55 19.3944
R7918 GND.n6529 GND.n55 19.3944
R7919 GND.n6529 GND.n6528 19.3944
R7920 GND.n6528 GND.n6527 19.3944
R7921 GND.n6527 GND.n60 19.3944
R7922 GND.n6523 GND.n60 19.3944
R7923 GND.n6523 GND.n6522 19.3944
R7924 GND.n6522 GND.n6521 19.3944
R7925 GND.n6521 GND.n65 19.3944
R7926 GND.n6517 GND.n65 19.3944
R7927 GND.n6517 GND.n6516 19.3944
R7928 GND.n6516 GND.n6515 19.3944
R7929 GND.n6515 GND.n70 19.3944
R7930 GND.n6511 GND.n70 19.3944
R7931 GND.n6511 GND.n6510 19.3944
R7932 GND.n6510 GND.n6509 19.3944
R7933 GND.n6509 GND.n75 19.3944
R7934 GND.n6505 GND.n75 19.3944
R7935 GND.n6505 GND.n6504 19.3944
R7936 GND.n5076 GND.n5075 18.4247
R7937 GND.n2581 GND.n2354 18.4247
R7938 GND.n4196 GND.n4195 16.4853
R7939 GND.n3511 GND.n2835 16.4853
R7940 GND.n2028 GND.n2023 16.2914
R7941 GND.n6448 GND.n6447 16.2914
R7942 GND.n5046 GND.n1219 16.2914
R7943 GND.n5008 GND.n1264 16.2914
R7944 GND.n3096 GND.n3095 16.2914
R7945 GND.n2542 GND.n2434 16.2914
R7946 GND.n5196 GND.n1006 16.2914
R7947 GND.n2504 GND.n2503 16.2914
R7948 GND.n5029 GND.n1233 16.1884
R7949 GND.n4648 GND.n1871 16.1884
R7950 GND.n4970 GND.n4969 15.5658
R7951 GND.n4969 GND.n4968 15.5658
R7952 GND.n4968 GND.n4967 15.5658
R7953 GND.n4967 GND.n1303 15.5658
R7954 GND.n3521 GND.n1303 15.5658
R7955 GND.n3521 GND.n1312 15.5658
R7956 GND.n4961 GND.n1312 15.5658
R7957 GND.n4960 GND.n1314 15.5658
R7958 GND.n1331 GND.n1314 15.5658
R7959 GND.n1332 GND.n1331 15.5658
R7960 GND.n4954 GND.n1332 15.5658
R7961 GND.n4954 GND.n4953 15.5658
R7962 GND.n4953 GND.n1334 15.5658
R7963 GND.n2826 GND.n1334 15.5658
R7964 GND.n2826 GND.n1345 15.5658
R7965 GND.n4947 GND.n1345 15.5658
R7966 GND.n4947 GND.n4946 15.5658
R7967 GND.n4946 GND.n1347 15.5658
R7968 GND.n1358 GND.n1347 15.5658
R7969 GND.n1359 GND.n1358 15.5658
R7970 GND.n4940 GND.n1359 15.5658
R7971 GND.n4940 GND.n4939 15.5658
R7972 GND.n4939 GND.n1361 15.5658
R7973 GND.n2823 GND.n1372 15.5658
R7974 GND.n4933 GND.n1372 15.5658
R7975 GND.n4933 GND.n4932 15.5658
R7976 GND.n4932 GND.n1374 15.5658
R7977 GND.n1385 GND.n1374 15.5658
R7978 GND.n1386 GND.n1385 15.5658
R7979 GND.n4926 GND.n1386 15.5658
R7980 GND.n4926 GND.n4925 15.5658
R7981 GND.n4925 GND.n1388 15.5658
R7982 GND.n3552 GND.n1388 15.5658
R7983 GND.n3552 GND.n1399 15.5658
R7984 GND.n4919 GND.n1399 15.5658
R7985 GND.n4919 GND.n4918 15.5658
R7986 GND.n4918 GND.n1401 15.5658
R7987 GND.n3562 GND.n3561 15.5658
R7988 GND.n4912 GND.n4911 15.5658
R7989 GND.n4905 GND.n1425 15.5658
R7990 GND.n3664 GND.n1434 15.5658
R7991 GND.n3703 GND.n3702 15.5658
R7992 GND.n3744 GND.n3743 15.5658
R7993 GND.n3726 GND.n1468 15.5658
R7994 GND.n3726 GND.n1474 15.5658
R7995 GND.n2686 GND.n2685 15.5658
R7996 GND.n2682 GND.n1488 15.5658
R7997 GND.n3792 GND.n2674 15.5658
R7998 GND.n3809 GND.n1507 15.5658
R7999 GND.n4841 GND.n1516 15.5658
R8000 GND.n4835 GND.n4834 15.5658
R8001 GND.n4828 GND.n1535 15.5658
R8002 GND.n4820 GND.n1546 15.5658
R8003 GND.n4814 GND.n1560 15.5658
R8004 GND.n4814 GND.n1563 15.5658
R8005 GND.n4807 GND.n1571 15.5658
R8006 GND.n4801 GND.n4800 15.5658
R8007 GND.n4794 GND.n1604 15.5658
R8008 GND.n4786 GND.n1615 15.5658
R8009 GND.n4780 GND.n1629 15.5658
R8010 GND.n4772 GND.n1640 15.5658
R8011 GND.n4766 GND.n4765 15.5658
R8012 GND.n4759 GND.n1673 15.5658
R8013 GND.n4752 GND.n1681 15.5658
R8014 GND.n4752 GND.n1684 15.5658
R8015 GND.n4746 GND.n1698 15.5658
R8016 GND.n4732 GND.n4731 15.5658
R8017 GND.n4725 GND.n1736 15.5658
R8018 GND.n4007 GND.n1745 15.5658
R8019 GND.n4711 GND.n4710 15.5658
R8020 GND.n2296 GND.n1766 15.5658
R8021 GND.n4704 GND.n1766 15.5658
R8022 GND.n4704 GND.n4703 15.5658
R8023 GND.n4703 GND.n1768 15.5658
R8024 GND.n4152 GND.n1768 15.5658
R8025 GND.n4152 GND.n1779 15.5658
R8026 GND.n4697 GND.n1779 15.5658
R8027 GND.n4697 GND.n4696 15.5658
R8028 GND.n4696 GND.n1781 15.5658
R8029 GND.n1792 GND.n1781 15.5658
R8030 GND.n1793 GND.n1792 15.5658
R8031 GND.n4690 GND.n1793 15.5658
R8032 GND.n4690 GND.n4689 15.5658
R8033 GND.n2289 GND.n2288 15.5658
R8034 GND.n2289 GND.n1805 15.5658
R8035 GND.n4683 GND.n1805 15.5658
R8036 GND.n4683 GND.n4682 15.5658
R8037 GND.n4682 GND.n1807 15.5658
R8038 GND.n1818 GND.n1807 15.5658
R8039 GND.n1819 GND.n1818 15.5658
R8040 GND.n4676 GND.n1819 15.5658
R8041 GND.n4676 GND.n4675 15.5658
R8042 GND.n4675 GND.n1821 15.5658
R8043 GND.n2285 GND.n1821 15.5658
R8044 GND.n2285 GND.n1832 15.5658
R8045 GND.n4669 GND.n1832 15.5658
R8046 GND.n4669 GND.n4668 15.5658
R8047 GND.n4668 GND.n1834 15.5658
R8048 GND.n1845 GND.n1834 15.5658
R8049 GND.n4662 GND.n1846 15.5658
R8050 GND.n4662 GND.n4661 15.5658
R8051 GND.n4661 GND.n1848 15.5658
R8052 GND.n4183 GND.n1848 15.5658
R8053 GND.n4183 GND.n1858 15.5658
R8054 GND.n4655 GND.n1858 15.5658
R8055 GND.n4655 GND.n4654 15.5658
R8056 GND.n5029 GND.n1247 14.9432
R8057 GND.n3656 GND.n3655 14.9432
R8058 GND.n4898 GND.n4897 14.9432
R8059 GND.n4849 GND.n4848 14.9432
R8060 GND.n3800 GND.n3799 14.9432
R8061 GND.n4787 GND.n1613 14.9432
R8062 GND.n4779 GND.n1631 14.9432
R8063 GND.n3998 GND.n3997 14.9432
R8064 GND.n4718 GND.n4717 14.9432
R8065 GND.n1871 GND.n1860 14.9432
R8066 GND.n2696 GND.n2693 14.3206
R8067 GND.n3757 GND.n3754 14.3206
R8068 GND.n4821 GND.n1543 14.3206
R8069 GND.n2652 GND.n2651 14.3206
R8070 GND.n3945 GND.n2635 14.3206
R8071 GND.n4745 GND.n1701 14.3206
R8072 GND.n3368 GND.t28 14.0093
R8073 GND.t15 GND.n2178 14.0093
R8074 GND.n4891 GND.n1445 13.698
R8075 GND.n4855 GND.n1496 13.698
R8076 GND.n3838 GND.n1526 13.698
R8077 GND.n3906 GND.n3905 13.698
R8078 GND.n2639 GND.n2638 13.698
R8079 GND.n3980 GND.n1725 13.698
R8080 GND.t99 GND.n2296 13.698
R8081 GND.n3643 GND.n3576 13.4249
R8082 GND.n4138 GND.n4137 13.4249
R8083 GND.n3570 GND.n3567 13.1884
R8084 GND.n2326 GND.n2323 13.1884
R8085 GND.n3712 GND.n1448 13.0754
R8086 GND.n3771 GND.n3770 13.0754
R8087 GND.n3954 GND.n1657 13.0754
R8088 GND.n2619 GND.n2618 13.0754
R8089 GND.n3646 GND.n3562 12.764
R8090 GND.n4710 GND.n1757 12.764
R8091 GND.n4884 GND.n4883 12.4527
R8092 GND.n4863 GND.n4862 12.4527
R8093 GND.n4827 GND.n1537 12.4527
R8094 GND.n3876 GND.n1588 12.4527
R8095 GND.n3963 GND.n1659 12.4527
R8096 GND.n4739 GND.n1707 12.4527
R8097 GND.n4143 GND.t74 12.4527
R8098 GND.n2712 GND.n1414 11.8301
R8099 GND.n3676 GND.n3675 11.8301
R8100 GND.n3791 GND.n3788 11.8301
R8101 GND.n3829 GND.n1524 11.8301
R8102 GND.n4793 GND.n1607 11.8301
R8103 GND.n4773 GND.n1637 11.8301
R8104 GND.n2612 GND.n1727 11.8301
R8105 GND.n2317 GND.n2316 11.8301
R8106 GND.n5264 GND.n967 11.5188
R8107 GND.n3280 GND.t6 11.5188
R8108 GND.t63 GND.n2855 11.5188
R8109 GND.t42 GND.n2664 11.5188
R8110 GND.n2644 GND.t136 11.5188
R8111 GND.t102 GND.n4279 11.5188
R8112 GND.t26 GND.n4401 11.5188
R8113 GND.n6444 GND.n135 11.5188
R8114 GND.n5188 GND.n5187 11.2075
R8115 GND.n1032 GND.n1018 11.2075
R8116 GND.n5181 GND.n1033 11.2075
R8117 GND.n3107 GND.n1051 11.2075
R8118 GND.n5174 GND.n1054 11.2075
R8119 GND.n3138 GND.n3115 11.2075
R8120 GND.n3140 GND.n3043 11.2075
R8121 GND.n3152 GND.n3045 11.2075
R8122 GND.n3142 GND.n3036 11.2075
R8123 GND.n3166 GND.n3031 11.2075
R8124 GND.n3170 GND.n3033 11.2075
R8125 GND.n3181 GND.n3019 11.2075
R8126 GND.n3180 GND.n3021 11.2075
R8127 GND.n3191 GND.n3011 11.2075
R8128 GND.n3192 GND.n3001 11.2075
R8129 GND.n3205 GND.n3004 11.2075
R8130 GND.n3215 GND.n2991 11.2075
R8131 GND.n3227 GND.n2983 11.2075
R8132 GND.n3229 GND.n2951 11.2075
R8133 GND.n3284 GND.n2953 11.2075
R8134 GND.n3281 GND.n3280 11.2075
R8135 GND.n3239 GND.n3237 11.2075
R8136 GND.n3273 GND.n2964 11.2075
R8137 GND.n3272 GND.n2966 11.2075
R8138 GND.n3267 GND.n2975 11.2075
R8139 GND.n3263 GND.n3262 11.2075
R8140 GND.n3292 GND.n2936 11.2075
R8141 GND.n3302 GND.n2928 11.2075
R8142 GND.n3301 GND.n2917 11.2075
R8143 GND.n3372 GND.n2920 11.2075
R8144 GND.n3369 GND.n3368 11.2075
R8145 GND.n3382 GND.n2907 11.2075
R8146 GND.n2911 GND.n2899 11.2075
R8147 GND.n3391 GND.n2895 11.2075
R8148 GND.n3397 GND.n2897 11.2075
R8149 GND.n3394 GND.n2887 11.2075
R8150 GND.n3355 GND.n2880 11.2075
R8151 GND.n3416 GND.n2876 11.2075
R8152 GND.n3422 GND.n2878 11.2075
R8153 GND.n3418 GND.n2865 11.2075
R8154 GND.n3432 GND.n2867 11.2075
R8155 GND.n2870 GND.n2858 11.2075
R8156 GND.n3447 GND.n2853 11.2075
R8157 GND.n3450 GND.n2855 11.2075
R8158 GND.n3439 GND.n2847 11.2075
R8159 GND.n3458 GND.n2845 11.2075
R8160 GND.n3463 GND.n1166 11.2075
R8161 GND.n5100 GND.n1168 11.2075
R8162 GND.n4877 GND.n1465 11.2075
R8163 GND.n4869 GND.n1477 11.2075
R8164 GND.n3852 GND.n2657 11.2075
R8165 GND.n4808 GND.n1569 11.2075
R8166 GND.n4758 GND.n1675 11.2075
R8167 GND.n3936 GND.n3935 11.2075
R8168 GND.n4640 GND.n4639 11.2075
R8169 GND.n2245 GND.n1883 11.2075
R8170 GND.n4633 GND.n1892 11.2075
R8171 GND.n4280 GND.n1895 11.2075
R8172 GND.n4279 GND.n4226 11.2075
R8173 GND.n4289 GND.n2237 11.2075
R8174 GND.n4295 GND.n2233 11.2075
R8175 GND.n4292 GND.n2235 11.2075
R8176 GND.n4305 GND.n2222 11.2075
R8177 GND.n2227 GND.n2223 11.2075
R8178 GND.n4314 GND.n2215 11.2075
R8179 GND.n4320 GND.n2211 11.2075
R8180 GND.n4330 GND.n2200 11.2075
R8181 GND.n2205 GND.n2202 11.2075
R8182 GND.n4339 GND.n2193 11.2075
R8183 GND.n4345 GND.n2188 11.2075
R8184 GND.n4342 GND.n2190 11.2075
R8185 GND.n4354 GND.n2178 11.2075
R8186 GND.n2179 GND.n2147 11.2075
R8187 GND.n4431 GND.n4430 11.2075
R8188 GND.n4362 GND.n2149 11.2075
R8189 GND.n4423 GND.n2157 11.2075
R8190 GND.n4419 GND.n2164 11.2075
R8191 GND.n4414 GND.n4413 11.2075
R8192 GND.n4382 GND.n4372 11.2075
R8193 GND.n4406 GND.n4380 11.2075
R8194 GND.n4402 GND.n4381 11.2075
R8195 GND.n4401 GND.n4393 11.2075
R8196 GND.n4387 GND.n2132 11.2075
R8197 GND.n4442 GND.n4441 11.2075
R8198 GND.n4446 GND.n2128 11.2075
R8199 GND.n2129 GND.n2119 11.2075
R8200 GND.n2120 GND.n2110 11.2075
R8201 GND.n4468 GND.n4467 11.2075
R8202 GND.n4472 GND.n2104 11.2075
R8203 GND.n2107 GND.n2094 11.2075
R8204 GND.n4483 GND.n4482 11.2075
R8205 GND.n2095 GND.n2087 11.2075
R8206 GND.n4496 GND.n4493 11.2075
R8207 GND.n4501 GND.n2084 11.2075
R8208 GND.n2085 GND.n2075 11.2075
R8209 GND.n4512 GND.n4511 11.2075
R8210 GND.n2076 GND.n2068 11.2075
R8211 GND.n4539 GND.n4538 11.2075
R8212 GND.n4543 GND.n2062 11.2075
R8213 GND.n4551 GND.n2055 11.2075
R8214 GND.n4554 GND.n2053 11.2075
R8215 GND.n6502 GND.n79 11.2075
R8216 GND.t44 GND.n3019 10.8962
R8217 GND.n3407 GND.t11 10.8962
R8218 GND.n5004 GND.n4978 10.8962
R8219 GND.n4961 GND.t85 10.8962
R8220 GND.t4 GND.n1412 10.8962
R8221 GND.n3711 GND.t46 10.8962
R8222 GND.n2625 GND.t139 10.8962
R8223 GND.n4141 GND.t60 10.8962
R8224 GND.n1846 GND.t124 10.8962
R8225 GND.n4646 GND.n1872 10.8962
R8226 GND.n4316 GND.t33 10.8962
R8227 GND.n4482 GND.t0 10.8962
R8228 GND.n2583 GND.n2353 10.6151
R8229 GND.n4071 GND.n2583 10.6151
R8230 GND.n4069 GND.n4068 10.6151
R8231 GND.n4068 GND.n2587 10.6151
R8232 GND.n4063 GND.n2587 10.6151
R8233 GND.n4063 GND.n4062 10.6151
R8234 GND.n4062 GND.n4061 10.6151
R8235 GND.n4061 GND.n2590 10.6151
R8236 GND.n4056 GND.n2590 10.6151
R8237 GND.n4056 GND.n4055 10.6151
R8238 GND.n4055 GND.n4054 10.6151
R8239 GND.n4054 GND.n2593 10.6151
R8240 GND.n4049 GND.n2593 10.6151
R8241 GND.n4049 GND.n4048 10.6151
R8242 GND.n4048 GND.n4047 10.6151
R8243 GND.n4047 GND.n2596 10.6151
R8244 GND.n4042 GND.n2596 10.6151
R8245 GND.n4042 GND.n4041 10.6151
R8246 GND.n4041 GND.n4040 10.6151
R8247 GND.n4040 GND.n2599 10.6151
R8248 GND.n4035 GND.n2599 10.6151
R8249 GND.n4035 GND.n4034 10.6151
R8250 GND.n4034 GND.n4033 10.6151
R8251 GND.n4033 GND.n2602 10.6151
R8252 GND.n4028 GND.n2602 10.6151
R8253 GND.n4028 GND.n4027 10.6151
R8254 GND.n4027 GND.n4026 10.6151
R8255 GND.n4026 GND.n2605 10.6151
R8256 GND.n4021 GND.n2605 10.6151
R8257 GND.n4021 GND.n4020 10.6151
R8258 GND.n4020 GND.n4019 10.6151
R8259 GND.n3651 GND.n2715 10.6151
R8260 GND.n3652 GND.n3651 10.6151
R8261 GND.n3653 GND.n3652 10.6151
R8262 GND.n3653 GND.n2708 10.6151
R8263 GND.n3667 GND.n2708 10.6151
R8264 GND.n3668 GND.n3667 10.6151
R8265 GND.n3669 GND.n3668 10.6151
R8266 GND.n3671 GND.n3669 10.6151
R8267 GND.n3671 GND.n3670 10.6151
R8268 GND.n3670 GND.n2702 10.6151
R8269 GND.n3714 GND.n2702 10.6151
R8270 GND.n3715 GND.n3714 10.6151
R8271 GND.n3716 GND.n3715 10.6151
R8272 GND.n3716 GND.n2701 10.6151
R8273 GND.n3720 GND.n2701 10.6151
R8274 GND.n3721 GND.n3720 10.6151
R8275 GND.n3724 GND.n3721 10.6151
R8276 GND.n3724 GND.n3723 10.6151
R8277 GND.n3723 GND.n3722 10.6151
R8278 GND.n3722 GND.n2683 10.6151
R8279 GND.n3760 GND.n2683 10.6151
R8280 GND.n3761 GND.n3760 10.6151
R8281 GND.n3768 GND.n3761 10.6151
R8282 GND.n3768 GND.n3767 10.6151
R8283 GND.n3767 GND.n3766 10.6151
R8284 GND.n3766 GND.n3764 10.6151
R8285 GND.n3764 GND.n3763 10.6151
R8286 GND.n3763 GND.n2669 10.6151
R8287 GND.n3812 GND.n2669 10.6151
R8288 GND.n3813 GND.n3812 10.6151
R8289 GND.n3814 GND.n3813 10.6151
R8290 GND.n3827 GND.n3814 10.6151
R8291 GND.n3827 GND.n3826 10.6151
R8292 GND.n3826 GND.n3825 10.6151
R8293 GND.n3825 GND.n3823 10.6151
R8294 GND.n3823 GND.n3822 10.6151
R8295 GND.n3822 GND.n3819 10.6151
R8296 GND.n3819 GND.n3818 10.6151
R8297 GND.n3818 GND.n3815 10.6151
R8298 GND.n3815 GND.n2655 10.6151
R8299 GND.n3855 GND.n2655 10.6151
R8300 GND.n3856 GND.n3855 10.6151
R8301 GND.n3859 GND.n3856 10.6151
R8302 GND.n3860 GND.n3859 10.6151
R8303 GND.n3861 GND.n3860 10.6151
R8304 GND.n3865 GND.n3861 10.6151
R8305 GND.n3865 GND.n3864 10.6151
R8306 GND.n3864 GND.n3863 10.6151
R8307 GND.n3863 GND.n2642 10.6151
R8308 GND.n3908 GND.n2642 10.6151
R8309 GND.n3909 GND.n3908 10.6151
R8310 GND.n3912 GND.n3909 10.6151
R8311 GND.n3913 GND.n3912 10.6151
R8312 GND.n3914 GND.n3913 10.6151
R8313 GND.n3920 GND.n3914 10.6151
R8314 GND.n3921 GND.n3920 10.6151
R8315 GND.n3924 GND.n3921 10.6151
R8316 GND.n3925 GND.n3924 10.6151
R8317 GND.n3926 GND.n3925 10.6151
R8318 GND.n3952 GND.n3926 10.6151
R8319 GND.n3952 GND.n3951 10.6151
R8320 GND.n3951 GND.n3950 10.6151
R8321 GND.n3950 GND.n3948 10.6151
R8322 GND.n3948 GND.n3947 10.6151
R8323 GND.n3947 GND.n3944 10.6151
R8324 GND.n3944 GND.n3943 10.6151
R8325 GND.n3943 GND.n3940 10.6151
R8326 GND.n3940 GND.n3939 10.6151
R8327 GND.n3939 GND.n3933 10.6151
R8328 GND.n3933 GND.n3932 10.6151
R8329 GND.n3932 GND.n3931 10.6151
R8330 GND.n3931 GND.n3928 10.6151
R8331 GND.n3928 GND.n3927 10.6151
R8332 GND.n3927 GND.n2617 10.6151
R8333 GND.n2617 GND.n2615 10.6151
R8334 GND.n3993 GND.n2615 10.6151
R8335 GND.n3994 GND.n3993 10.6151
R8336 GND.n3995 GND.n3994 10.6151
R8337 GND.n3995 GND.n2608 10.6151
R8338 GND.n4010 GND.n2608 10.6151
R8339 GND.n4011 GND.n4010 10.6151
R8340 GND.n4012 GND.n4011 10.6151
R8341 GND.n4015 GND.n4012 10.6151
R8342 GND.n4016 GND.n4015 10.6151
R8343 GND.n2757 GND.n2754 10.6151
R8344 GND.n2758 GND.n2757 10.6151
R8345 GND.n2762 GND.n2761 10.6151
R8346 GND.n2765 GND.n2762 10.6151
R8347 GND.n2766 GND.n2765 10.6151
R8348 GND.n2769 GND.n2766 10.6151
R8349 GND.n2770 GND.n2769 10.6151
R8350 GND.n2773 GND.n2770 10.6151
R8351 GND.n2774 GND.n2773 10.6151
R8352 GND.n2777 GND.n2774 10.6151
R8353 GND.n2778 GND.n2777 10.6151
R8354 GND.n2781 GND.n2778 10.6151
R8355 GND.n2782 GND.n2781 10.6151
R8356 GND.n2785 GND.n2782 10.6151
R8357 GND.n2786 GND.n2785 10.6151
R8358 GND.n2789 GND.n2786 10.6151
R8359 GND.n2790 GND.n2789 10.6151
R8360 GND.n2793 GND.n2790 10.6151
R8361 GND.n2794 GND.n2793 10.6151
R8362 GND.n2797 GND.n2794 10.6151
R8363 GND.n2798 GND.n2797 10.6151
R8364 GND.n2801 GND.n2798 10.6151
R8365 GND.n2802 GND.n2801 10.6151
R8366 GND.n2805 GND.n2802 10.6151
R8367 GND.n2806 GND.n2805 10.6151
R8368 GND.n2809 GND.n2806 10.6151
R8369 GND.n2811 GND.n2809 10.6151
R8370 GND.n2812 GND.n2811 10.6151
R8371 GND.n2814 GND.n2812 10.6151
R8372 GND.n2814 GND.n2813 10.6151
R8373 GND.n2813 GND.n2716 10.6151
R8374 GND.n3643 GND.n3642 10.6151
R8375 GND.n3642 GND.n3641 10.6151
R8376 GND.n3641 GND.n3640 10.6151
R8377 GND.n3640 GND.n3638 10.6151
R8378 GND.n3638 GND.n3635 10.6151
R8379 GND.n3635 GND.n3634 10.6151
R8380 GND.n3634 GND.n3631 10.6151
R8381 GND.n3631 GND.n3630 10.6151
R8382 GND.n3630 GND.n3627 10.6151
R8383 GND.n3627 GND.n3626 10.6151
R8384 GND.n3626 GND.n3623 10.6151
R8385 GND.n3623 GND.n3622 10.6151
R8386 GND.n3622 GND.n3619 10.6151
R8387 GND.n3619 GND.n3618 10.6151
R8388 GND.n3618 GND.n3615 10.6151
R8389 GND.n3615 GND.n3614 10.6151
R8390 GND.n3614 GND.n3611 10.6151
R8391 GND.n3611 GND.n3610 10.6151
R8392 GND.n3610 GND.n3607 10.6151
R8393 GND.n3607 GND.n3606 10.6151
R8394 GND.n3606 GND.n3603 10.6151
R8395 GND.n3603 GND.n3602 10.6151
R8396 GND.n3602 GND.n3599 10.6151
R8397 GND.n3599 GND.n3598 10.6151
R8398 GND.n3598 GND.n3595 10.6151
R8399 GND.n3595 GND.n3594 10.6151
R8400 GND.n3594 GND.n3591 10.6151
R8401 GND.n3591 GND.n3590 10.6151
R8402 GND.n3590 GND.n3587 10.6151
R8403 GND.n3585 GND.n3582 10.6151
R8404 GND.n3582 GND.n3581 10.6151
R8405 GND.n4137 GND.n4136 10.6151
R8406 GND.n4136 GND.n2327 10.6151
R8407 GND.n2328 GND.n2327 10.6151
R8408 GND.n4129 GND.n2328 10.6151
R8409 GND.n4129 GND.n4128 10.6151
R8410 GND.n4128 GND.n4127 10.6151
R8411 GND.n4127 GND.n2330 10.6151
R8412 GND.n4122 GND.n2330 10.6151
R8413 GND.n4122 GND.n4121 10.6151
R8414 GND.n4121 GND.n4120 10.6151
R8415 GND.n4120 GND.n2333 10.6151
R8416 GND.n4115 GND.n2333 10.6151
R8417 GND.n4115 GND.n4114 10.6151
R8418 GND.n4114 GND.n4113 10.6151
R8419 GND.n4113 GND.n2336 10.6151
R8420 GND.n4108 GND.n2336 10.6151
R8421 GND.n4108 GND.n4107 10.6151
R8422 GND.n4107 GND.n4106 10.6151
R8423 GND.n4106 GND.n2339 10.6151
R8424 GND.n4101 GND.n2339 10.6151
R8425 GND.n4101 GND.n4100 10.6151
R8426 GND.n4100 GND.n4099 10.6151
R8427 GND.n4099 GND.n2342 10.6151
R8428 GND.n4094 GND.n2342 10.6151
R8429 GND.n4094 GND.n4093 10.6151
R8430 GND.n4093 GND.n4092 10.6151
R8431 GND.n4092 GND.n2345 10.6151
R8432 GND.n4087 GND.n2345 10.6151
R8433 GND.n4087 GND.n4086 10.6151
R8434 GND.n4084 GND.n2350 10.6151
R8435 GND.n4079 GND.n2350 10.6151
R8436 GND.n3575 GND.n3574 10.6151
R8437 GND.n3574 GND.n3571 10.6151
R8438 GND.n3571 GND.n1431 10.6151
R8439 GND.n4902 GND.n1431 10.6151
R8440 GND.n4902 GND.n4901 10.6151
R8441 GND.n4901 GND.n4900 10.6151
R8442 GND.n4900 GND.n1432 10.6151
R8443 GND.n3673 GND.n1432 10.6151
R8444 GND.n3673 GND.n1451 10.6151
R8445 GND.n4888 GND.n1451 10.6151
R8446 GND.n4888 GND.n4887 10.6151
R8447 GND.n4887 GND.n4886 10.6151
R8448 GND.n4886 GND.n1452 10.6151
R8449 GND.n2694 GND.n1452 10.6151
R8450 GND.n2694 GND.n1471 10.6151
R8451 GND.n4874 GND.n1471 10.6151
R8452 GND.n4874 GND.n4873 10.6151
R8453 GND.n4873 GND.n4872 10.6151
R8454 GND.n4872 GND.n1472 10.6151
R8455 GND.n3755 GND.n1472 10.6151
R8456 GND.n3755 GND.n1491 10.6151
R8457 GND.n4860 GND.n1491 10.6151
R8458 GND.n4860 GND.n4859 10.6151
R8459 GND.n4859 GND.n4858 10.6151
R8460 GND.n4858 GND.n1492 10.6151
R8461 GND.n3789 GND.n1492 10.6151
R8462 GND.n3789 GND.n1510 10.6151
R8463 GND.n4846 GND.n1510 10.6151
R8464 GND.n4846 GND.n4845 10.6151
R8465 GND.n4845 GND.n4844 10.6151
R8466 GND.n4844 GND.n1511 10.6151
R8467 GND.n2666 GND.n1511 10.6151
R8468 GND.n3833 GND.n2666 10.6151
R8469 GND.n3834 GND.n3833 10.6151
R8470 GND.n3835 GND.n3834 10.6151
R8471 GND.n3835 GND.n1540 10.6151
R8472 GND.n4825 GND.n1540 10.6151
R8473 GND.n4825 GND.n4824 10.6151
R8474 GND.n4824 GND.n4823 10.6151
R8475 GND.n4823 GND.n1541 10.6151
R8476 GND.n1566 GND.n1541 10.6151
R8477 GND.n4812 GND.n1566 10.6151
R8478 GND.n4812 GND.n4811 10.6151
R8479 GND.n4811 GND.n4810 10.6151
R8480 GND.n4810 GND.n1567 10.6151
R8481 GND.n3873 GND.n1567 10.6151
R8482 GND.n3873 GND.n3872 10.6151
R8483 GND.n3872 GND.n3871 10.6151
R8484 GND.n3871 GND.n3868 10.6151
R8485 GND.n3868 GND.n1610 10.6151
R8486 GND.n4791 GND.n1610 10.6151
R8487 GND.n4791 GND.n4790 10.6151
R8488 GND.n4790 GND.n4789 10.6151
R8489 GND.n4789 GND.n1611 10.6151
R8490 GND.n1634 GND.n1611 10.6151
R8491 GND.n4777 GND.n1634 10.6151
R8492 GND.n4777 GND.n4776 10.6151
R8493 GND.n4776 GND.n4775 10.6151
R8494 GND.n4775 GND.n1635 10.6151
R8495 GND.n2637 GND.n1635 10.6151
R8496 GND.n3958 GND.n2637 10.6151
R8497 GND.n3959 GND.n3958 10.6151
R8498 GND.n3960 GND.n3959 10.6151
R8499 GND.n3960 GND.n1678 10.6151
R8500 GND.n4756 GND.n1678 10.6151
R8501 GND.n4756 GND.n4755 10.6151
R8502 GND.n4755 GND.n4754 10.6151
R8503 GND.n4754 GND.n1679 10.6151
R8504 GND.n1704 GND.n1679 10.6151
R8505 GND.n4743 GND.n1704 10.6151
R8506 GND.n4743 GND.n4742 10.6151
R8507 GND.n4742 GND.n4741 10.6151
R8508 GND.n4741 GND.n1705 10.6151
R8509 GND.n3987 GND.n1705 10.6151
R8510 GND.n3987 GND.n3986 10.6151
R8511 GND.n3986 GND.n3985 10.6151
R8512 GND.n3985 GND.n3982 10.6151
R8513 GND.n3982 GND.n1742 10.6151
R8514 GND.n4722 GND.n1742 10.6151
R8515 GND.n4722 GND.n4721 10.6151
R8516 GND.n4721 GND.n4720 10.6151
R8517 GND.n4720 GND.n1743 10.6151
R8518 GND.n2321 GND.n1743 10.6151
R8519 GND.n4139 GND.n2321 10.6151
R8520 GND.n4904 GND.n1428 10.5849
R8521 GND.n3665 GND.n1428 10.5849
R8522 GND.n3810 GND.n1513 10.5849
R8523 GND.n4842 GND.n1513 10.5849
R8524 GND.n3917 GND.n3916 10.5849
R8525 GND.n3918 GND.n3917 10.5849
R8526 GND.n4724 GND.n1739 10.5849
R8527 GND.n4008 GND.n1739 10.5849
R8528 GND.t57 GND.n1361 10.2736
R8529 GND.n2288 GND.t36 10.2736
R8530 GND.n4877 GND.n4876 9.96229
R8531 GND.n4870 GND.n4869 9.96229
R8532 GND.n3853 GND.n3852 9.96229
R8533 GND.n3857 GND.n1569 9.96229
R8534 GND.n3941 GND.n1675 9.96229
R8535 GND.n3937 GND.n3936 9.96229
R8536 GND.n2024 GND.n2023 9.69747
R8537 GND.n6449 GND.n6448 9.69747
R8538 GND.n5050 GND.n1219 9.69747
R8539 GND.n5008 GND.n5007 9.69747
R8540 GND.n3097 GND.n3096 9.69747
R8541 GND.n2548 GND.n2434 9.69747
R8542 GND.n5199 GND.n5196 9.69747
R8543 GND.n2503 GND.n2484 9.69747
R8544 GND.n4197 GND.n4196 9.50353
R8545 GND.n3507 GND.n2835 9.50353
R8546 GND.n3676 GND.n1437 9.33968
R8547 GND.n3788 GND.n1504 9.33968
R8548 GND.n3830 GND.n3829 9.33968
R8549 GND.n3910 GND.n1607 9.33968
R8550 GND.n3922 GND.n1637 9.33968
R8551 GND.n2613 GND.n2612 9.33968
R8552 GND.n2316 GND.n1748 9.33968
R8553 GND.n4965 GND.n1307 9.3005
R8554 GND.n4964 GND.n1308 9.3005
R8555 GND.n4963 GND.n1309 9.3005
R8556 GND.n1338 GND.n1310 9.3005
R8557 GND.n1339 GND.n1337 9.3005
R8558 GND.n4951 GND.n1340 9.3005
R8559 GND.n4950 GND.n1341 9.3005
R8560 GND.n4949 GND.n1342 9.3005
R8561 GND.n1365 GND.n1343 9.3005
R8562 GND.n1366 GND.n1364 9.3005
R8563 GND.n4937 GND.n1367 9.3005
R8564 GND.n4936 GND.n1368 9.3005
R8565 GND.n4935 GND.n1369 9.3005
R8566 GND.n1392 GND.n1370 9.3005
R8567 GND.n1393 GND.n1391 9.3005
R8568 GND.n4923 GND.n1394 9.3005
R8569 GND.n4922 GND.n1395 9.3005
R8570 GND.n4921 GND.n1396 9.3005
R8571 GND.n1418 GND.n1397 9.3005
R8572 GND.n1419 GND.n1417 9.3005
R8573 GND.n4909 GND.n1420 9.3005
R8574 GND.n4908 GND.n1421 9.3005
R8575 GND.n4907 GND.n1422 9.3005
R8576 GND.n1439 GND.n1423 9.3005
R8577 GND.n4895 GND.n1440 9.3005
R8578 GND.n4894 GND.n1441 9.3005
R8579 GND.n4893 GND.n1442 9.3005
R8580 GND.n1459 GND.n1443 9.3005
R8581 GND.n4881 GND.n1460 9.3005
R8582 GND.n4880 GND.n1461 9.3005
R8583 GND.n4879 GND.n1462 9.3005
R8584 GND.n1479 GND.n1463 9.3005
R8585 GND.n4867 GND.n1480 9.3005
R8586 GND.n4866 GND.n1481 9.3005
R8587 GND.n4865 GND.n1482 9.3005
R8588 GND.n1498 GND.n1483 9.3005
R8589 GND.n4853 GND.n1499 9.3005
R8590 GND.n4852 GND.n1500 9.3005
R8591 GND.n4851 GND.n1501 9.3005
R8592 GND.n1518 GND.n1502 9.3005
R8593 GND.n4839 GND.n1519 9.3005
R8594 GND.n4838 GND.n1520 9.3005
R8595 GND.n4837 GND.n1521 9.3005
R8596 GND.n1550 GND.n1522 9.3005
R8597 GND.n1553 GND.n1552 9.3005
R8598 GND.n1554 GND.n1549 9.3005
R8599 GND.n4818 GND.n1555 9.3005
R8600 GND.n4817 GND.n1556 9.3005
R8601 GND.n4816 GND.n1557 9.3005
R8602 GND.n1594 GND.n1558 9.3005
R8603 GND.n1597 GND.n1596 9.3005
R8604 GND.n1598 GND.n1593 9.3005
R8605 GND.n4798 GND.n1599 9.3005
R8606 GND.n4797 GND.n1600 9.3005
R8607 GND.n4796 GND.n1601 9.3005
R8608 GND.n1644 GND.n1602 9.3005
R8609 GND.n1646 GND.n1645 9.3005
R8610 GND.n1650 GND.n1649 9.3005
R8611 GND.n1651 GND.n1643 9.3005
R8612 GND.n4770 GND.n1652 9.3005
R8613 GND.n4769 GND.n1653 9.3005
R8614 GND.n4768 GND.n1654 9.3005
R8615 GND.n1688 GND.n1655 9.3005
R8616 GND.n1691 GND.n1690 9.3005
R8617 GND.n1692 GND.n1687 9.3005
R8618 GND.n4750 GND.n1693 9.3005
R8619 GND.n4749 GND.n1694 9.3005
R8620 GND.n4748 GND.n1695 9.3005
R8621 GND.n2620 GND.n1696 9.3005
R8622 GND.n2623 GND.n2622 9.3005
R8623 GND.n2621 GND.n1730 9.3005
R8624 GND.n4729 GND.n1731 9.3005
R8625 GND.n4728 GND.n1732 9.3005
R8626 GND.n4727 GND.n1733 9.3005
R8627 GND.n1750 GND.n1734 9.3005
R8628 GND.n4715 GND.n1751 9.3005
R8629 GND.n4714 GND.n1752 9.3005
R8630 GND.n4713 GND.n1753 9.3005
R8631 GND.n1772 GND.n1754 9.3005
R8632 GND.n1773 GND.n1771 9.3005
R8633 GND.n4701 GND.n1774 9.3005
R8634 GND.n4700 GND.n1775 9.3005
R8635 GND.n4699 GND.n1776 9.3005
R8636 GND.n1798 GND.n1777 9.3005
R8637 GND.n1799 GND.n1797 9.3005
R8638 GND.n4687 GND.n1800 9.3005
R8639 GND.n4686 GND.n1801 9.3005
R8640 GND.n4685 GND.n1802 9.3005
R8641 GND.n1825 GND.n1803 9.3005
R8642 GND.n1826 GND.n1824 9.3005
R8643 GND.n4673 GND.n1827 9.3005
R8644 GND.n4672 GND.n1828 9.3005
R8645 GND.n4671 GND.n1829 9.3005
R8646 GND.n1852 GND.n1830 9.3005
R8647 GND.n1853 GND.n1851 9.3005
R8648 GND.n4659 GND.n1854 9.3005
R8649 GND.n4658 GND.n1855 9.3005
R8650 GND.n4657 GND.n1856 9.3005
R8651 GND.n1306 GND.n1305 9.3005
R8652 GND.n5462 GND.n747 9.3005
R8653 GND.n5464 GND.n5463 9.3005
R8654 GND.n743 GND.n742 9.3005
R8655 GND.n5471 GND.n5470 9.3005
R8656 GND.n5472 GND.n741 9.3005
R8657 GND.n5474 GND.n5473 9.3005
R8658 GND.n737 GND.n736 9.3005
R8659 GND.n5481 GND.n5480 9.3005
R8660 GND.n5482 GND.n735 9.3005
R8661 GND.n5484 GND.n5483 9.3005
R8662 GND.n731 GND.n730 9.3005
R8663 GND.n5491 GND.n5490 9.3005
R8664 GND.n5492 GND.n729 9.3005
R8665 GND.n5494 GND.n5493 9.3005
R8666 GND.n725 GND.n724 9.3005
R8667 GND.n5501 GND.n5500 9.3005
R8668 GND.n5502 GND.n723 9.3005
R8669 GND.n5504 GND.n5503 9.3005
R8670 GND.n719 GND.n718 9.3005
R8671 GND.n5511 GND.n5510 9.3005
R8672 GND.n5512 GND.n717 9.3005
R8673 GND.n5514 GND.n5513 9.3005
R8674 GND.n713 GND.n712 9.3005
R8675 GND.n5521 GND.n5520 9.3005
R8676 GND.n5522 GND.n711 9.3005
R8677 GND.n5524 GND.n5523 9.3005
R8678 GND.n707 GND.n706 9.3005
R8679 GND.n5531 GND.n5530 9.3005
R8680 GND.n5532 GND.n705 9.3005
R8681 GND.n5534 GND.n5533 9.3005
R8682 GND.n701 GND.n700 9.3005
R8683 GND.n5541 GND.n5540 9.3005
R8684 GND.n5542 GND.n699 9.3005
R8685 GND.n5544 GND.n5543 9.3005
R8686 GND.n695 GND.n694 9.3005
R8687 GND.n5551 GND.n5550 9.3005
R8688 GND.n5552 GND.n693 9.3005
R8689 GND.n5554 GND.n5553 9.3005
R8690 GND.n689 GND.n688 9.3005
R8691 GND.n5561 GND.n5560 9.3005
R8692 GND.n5562 GND.n687 9.3005
R8693 GND.n5564 GND.n5563 9.3005
R8694 GND.n683 GND.n682 9.3005
R8695 GND.n5571 GND.n5570 9.3005
R8696 GND.n5572 GND.n681 9.3005
R8697 GND.n5574 GND.n5573 9.3005
R8698 GND.n677 GND.n676 9.3005
R8699 GND.n5581 GND.n5580 9.3005
R8700 GND.n5582 GND.n675 9.3005
R8701 GND.n5584 GND.n5583 9.3005
R8702 GND.n671 GND.n670 9.3005
R8703 GND.n5591 GND.n5590 9.3005
R8704 GND.n5592 GND.n669 9.3005
R8705 GND.n5594 GND.n5593 9.3005
R8706 GND.n665 GND.n664 9.3005
R8707 GND.n5601 GND.n5600 9.3005
R8708 GND.n5602 GND.n663 9.3005
R8709 GND.n5604 GND.n5603 9.3005
R8710 GND.n659 GND.n658 9.3005
R8711 GND.n5611 GND.n5610 9.3005
R8712 GND.n5612 GND.n657 9.3005
R8713 GND.n5614 GND.n5613 9.3005
R8714 GND.n653 GND.n652 9.3005
R8715 GND.n5621 GND.n5620 9.3005
R8716 GND.n5622 GND.n651 9.3005
R8717 GND.n5624 GND.n5623 9.3005
R8718 GND.n647 GND.n646 9.3005
R8719 GND.n5631 GND.n5630 9.3005
R8720 GND.n5632 GND.n645 9.3005
R8721 GND.n5634 GND.n5633 9.3005
R8722 GND.n641 GND.n640 9.3005
R8723 GND.n5641 GND.n5640 9.3005
R8724 GND.n5642 GND.n639 9.3005
R8725 GND.n5644 GND.n5643 9.3005
R8726 GND.n635 GND.n634 9.3005
R8727 GND.n5651 GND.n5650 9.3005
R8728 GND.n5652 GND.n633 9.3005
R8729 GND.n5654 GND.n5653 9.3005
R8730 GND.n629 GND.n628 9.3005
R8731 GND.n5661 GND.n5660 9.3005
R8732 GND.n5662 GND.n627 9.3005
R8733 GND.n5664 GND.n5663 9.3005
R8734 GND.n623 GND.n622 9.3005
R8735 GND.n5671 GND.n5670 9.3005
R8736 GND.n5672 GND.n621 9.3005
R8737 GND.n5674 GND.n5673 9.3005
R8738 GND.n617 GND.n616 9.3005
R8739 GND.n5681 GND.n5680 9.3005
R8740 GND.n5682 GND.n615 9.3005
R8741 GND.n5684 GND.n5683 9.3005
R8742 GND.n611 GND.n610 9.3005
R8743 GND.n5691 GND.n5690 9.3005
R8744 GND.n5692 GND.n609 9.3005
R8745 GND.n5694 GND.n5693 9.3005
R8746 GND.n605 GND.n604 9.3005
R8747 GND.n5701 GND.n5700 9.3005
R8748 GND.n5702 GND.n603 9.3005
R8749 GND.n5704 GND.n5703 9.3005
R8750 GND.n599 GND.n598 9.3005
R8751 GND.n5711 GND.n5710 9.3005
R8752 GND.n5712 GND.n597 9.3005
R8753 GND.n5714 GND.n5713 9.3005
R8754 GND.n593 GND.n592 9.3005
R8755 GND.n5721 GND.n5720 9.3005
R8756 GND.n5722 GND.n591 9.3005
R8757 GND.n5724 GND.n5723 9.3005
R8758 GND.n587 GND.n586 9.3005
R8759 GND.n5731 GND.n5730 9.3005
R8760 GND.n5732 GND.n585 9.3005
R8761 GND.n5734 GND.n5733 9.3005
R8762 GND.n581 GND.n580 9.3005
R8763 GND.n5741 GND.n5740 9.3005
R8764 GND.n5742 GND.n579 9.3005
R8765 GND.n5744 GND.n5743 9.3005
R8766 GND.n575 GND.n574 9.3005
R8767 GND.n5751 GND.n5750 9.3005
R8768 GND.n5752 GND.n573 9.3005
R8769 GND.n5754 GND.n5753 9.3005
R8770 GND.n569 GND.n568 9.3005
R8771 GND.n5761 GND.n5760 9.3005
R8772 GND.n5762 GND.n567 9.3005
R8773 GND.n5764 GND.n5763 9.3005
R8774 GND.n563 GND.n562 9.3005
R8775 GND.n5771 GND.n5770 9.3005
R8776 GND.n5772 GND.n561 9.3005
R8777 GND.n5774 GND.n5773 9.3005
R8778 GND.n557 GND.n556 9.3005
R8779 GND.n5781 GND.n5780 9.3005
R8780 GND.n5782 GND.n555 9.3005
R8781 GND.n5784 GND.n5783 9.3005
R8782 GND.n551 GND.n550 9.3005
R8783 GND.n5791 GND.n5790 9.3005
R8784 GND.n5792 GND.n549 9.3005
R8785 GND.n5794 GND.n5793 9.3005
R8786 GND.n545 GND.n544 9.3005
R8787 GND.n5801 GND.n5800 9.3005
R8788 GND.n5802 GND.n543 9.3005
R8789 GND.n5804 GND.n5803 9.3005
R8790 GND.n539 GND.n538 9.3005
R8791 GND.n5811 GND.n5810 9.3005
R8792 GND.n5812 GND.n537 9.3005
R8793 GND.n5814 GND.n5813 9.3005
R8794 GND.n533 GND.n532 9.3005
R8795 GND.n5821 GND.n5820 9.3005
R8796 GND.n5822 GND.n531 9.3005
R8797 GND.n5824 GND.n5823 9.3005
R8798 GND.n527 GND.n526 9.3005
R8799 GND.n5831 GND.n5830 9.3005
R8800 GND.n5832 GND.n525 9.3005
R8801 GND.n5834 GND.n5833 9.3005
R8802 GND.n521 GND.n520 9.3005
R8803 GND.n5841 GND.n5840 9.3005
R8804 GND.n5842 GND.n519 9.3005
R8805 GND.n5844 GND.n5843 9.3005
R8806 GND.n515 GND.n514 9.3005
R8807 GND.n5851 GND.n5850 9.3005
R8808 GND.n5852 GND.n513 9.3005
R8809 GND.n5854 GND.n5853 9.3005
R8810 GND.n509 GND.n508 9.3005
R8811 GND.n5861 GND.n5860 9.3005
R8812 GND.n5862 GND.n507 9.3005
R8813 GND.n5864 GND.n5863 9.3005
R8814 GND.n503 GND.n502 9.3005
R8815 GND.n5871 GND.n5870 9.3005
R8816 GND.n5872 GND.n501 9.3005
R8817 GND.n5874 GND.n5873 9.3005
R8818 GND.n497 GND.n496 9.3005
R8819 GND.n5881 GND.n5880 9.3005
R8820 GND.n5882 GND.n495 9.3005
R8821 GND.n5884 GND.n5883 9.3005
R8822 GND.n491 GND.n490 9.3005
R8823 GND.n5891 GND.n5890 9.3005
R8824 GND.n5892 GND.n489 9.3005
R8825 GND.n5894 GND.n5893 9.3005
R8826 GND.n485 GND.n484 9.3005
R8827 GND.n5901 GND.n5900 9.3005
R8828 GND.n5902 GND.n483 9.3005
R8829 GND.n5904 GND.n5903 9.3005
R8830 GND.n479 GND.n478 9.3005
R8831 GND.n5911 GND.n5910 9.3005
R8832 GND.n5912 GND.n477 9.3005
R8833 GND.n5914 GND.n5913 9.3005
R8834 GND.n473 GND.n472 9.3005
R8835 GND.n5921 GND.n5920 9.3005
R8836 GND.n5922 GND.n471 9.3005
R8837 GND.n5924 GND.n5923 9.3005
R8838 GND.n467 GND.n466 9.3005
R8839 GND.n5931 GND.n5930 9.3005
R8840 GND.n5932 GND.n465 9.3005
R8841 GND.n5934 GND.n5933 9.3005
R8842 GND.n461 GND.n460 9.3005
R8843 GND.n5941 GND.n5940 9.3005
R8844 GND.n5942 GND.n459 9.3005
R8845 GND.n5944 GND.n5943 9.3005
R8846 GND.n455 GND.n454 9.3005
R8847 GND.n5951 GND.n5950 9.3005
R8848 GND.n5952 GND.n453 9.3005
R8849 GND.n5954 GND.n5953 9.3005
R8850 GND.n449 GND.n448 9.3005
R8851 GND.n5961 GND.n5960 9.3005
R8852 GND.n5962 GND.n447 9.3005
R8853 GND.n5964 GND.n5963 9.3005
R8854 GND.n443 GND.n442 9.3005
R8855 GND.n5971 GND.n5970 9.3005
R8856 GND.n5972 GND.n441 9.3005
R8857 GND.n5974 GND.n5973 9.3005
R8858 GND.n437 GND.n436 9.3005
R8859 GND.n5981 GND.n5980 9.3005
R8860 GND.n5982 GND.n435 9.3005
R8861 GND.n5984 GND.n5983 9.3005
R8862 GND.n431 GND.n430 9.3005
R8863 GND.n5991 GND.n5990 9.3005
R8864 GND.n5992 GND.n429 9.3005
R8865 GND.n5994 GND.n5993 9.3005
R8866 GND.n425 GND.n424 9.3005
R8867 GND.n6001 GND.n6000 9.3005
R8868 GND.n6002 GND.n423 9.3005
R8869 GND.n6004 GND.n6003 9.3005
R8870 GND.n419 GND.n418 9.3005
R8871 GND.n6011 GND.n6010 9.3005
R8872 GND.n6012 GND.n417 9.3005
R8873 GND.n6014 GND.n6013 9.3005
R8874 GND.n413 GND.n412 9.3005
R8875 GND.n6021 GND.n6020 9.3005
R8876 GND.n6022 GND.n411 9.3005
R8877 GND.n6024 GND.n6023 9.3005
R8878 GND.n407 GND.n406 9.3005
R8879 GND.n6031 GND.n6030 9.3005
R8880 GND.n6032 GND.n405 9.3005
R8881 GND.n6034 GND.n6033 9.3005
R8882 GND.n401 GND.n400 9.3005
R8883 GND.n6041 GND.n6040 9.3005
R8884 GND.n6042 GND.n399 9.3005
R8885 GND.n6044 GND.n6043 9.3005
R8886 GND.n395 GND.n394 9.3005
R8887 GND.n6051 GND.n6050 9.3005
R8888 GND.n6052 GND.n393 9.3005
R8889 GND.n6054 GND.n6053 9.3005
R8890 GND.n389 GND.n388 9.3005
R8891 GND.n6061 GND.n6060 9.3005
R8892 GND.n6062 GND.n387 9.3005
R8893 GND.n6064 GND.n6063 9.3005
R8894 GND.n383 GND.n382 9.3005
R8895 GND.n6071 GND.n6070 9.3005
R8896 GND.n6072 GND.n381 9.3005
R8897 GND.n6074 GND.n6073 9.3005
R8898 GND.n377 GND.n376 9.3005
R8899 GND.n6081 GND.n6080 9.3005
R8900 GND.n6082 GND.n375 9.3005
R8901 GND.n6084 GND.n6083 9.3005
R8902 GND.n371 GND.n370 9.3005
R8903 GND.n6091 GND.n6090 9.3005
R8904 GND.n6092 GND.n369 9.3005
R8905 GND.n6094 GND.n6093 9.3005
R8906 GND.n365 GND.n364 9.3005
R8907 GND.n6101 GND.n6100 9.3005
R8908 GND.n6102 GND.n363 9.3005
R8909 GND.n6104 GND.n6103 9.3005
R8910 GND.n359 GND.n358 9.3005
R8911 GND.n6111 GND.n6110 9.3005
R8912 GND.n6112 GND.n357 9.3005
R8913 GND.n6114 GND.n6113 9.3005
R8914 GND.n353 GND.n352 9.3005
R8915 GND.n6121 GND.n6120 9.3005
R8916 GND.n6122 GND.n351 9.3005
R8917 GND.n6124 GND.n6123 9.3005
R8918 GND.n347 GND.n346 9.3005
R8919 GND.n6131 GND.n6130 9.3005
R8920 GND.n6132 GND.n345 9.3005
R8921 GND.n6134 GND.n6133 9.3005
R8922 GND.n341 GND.n340 9.3005
R8923 GND.n6141 GND.n6140 9.3005
R8924 GND.n6142 GND.n339 9.3005
R8925 GND.n6144 GND.n6143 9.3005
R8926 GND.n335 GND.n334 9.3005
R8927 GND.n6151 GND.n6150 9.3005
R8928 GND.n6152 GND.n333 9.3005
R8929 GND.n6154 GND.n6153 9.3005
R8930 GND.n329 GND.n328 9.3005
R8931 GND.n6161 GND.n6160 9.3005
R8932 GND.n6162 GND.n327 9.3005
R8933 GND.n6164 GND.n6163 9.3005
R8934 GND.n323 GND.n322 9.3005
R8935 GND.n6171 GND.n6170 9.3005
R8936 GND.n6172 GND.n321 9.3005
R8937 GND.n6174 GND.n6173 9.3005
R8938 GND.n317 GND.n316 9.3005
R8939 GND.n6181 GND.n6180 9.3005
R8940 GND.n6182 GND.n315 9.3005
R8941 GND.n6184 GND.n6183 9.3005
R8942 GND.n311 GND.n310 9.3005
R8943 GND.n6191 GND.n6190 9.3005
R8944 GND.n6194 GND.n6193 9.3005
R8945 GND.n305 GND.n304 9.3005
R8946 GND.n6201 GND.n6200 9.3005
R8947 GND.n6202 GND.n303 9.3005
R8948 GND.n6204 GND.n6203 9.3005
R8949 GND.n299 GND.n298 9.3005
R8950 GND.n6211 GND.n6210 9.3005
R8951 GND.n6212 GND.n297 9.3005
R8952 GND.n6214 GND.n6213 9.3005
R8953 GND.n293 GND.n292 9.3005
R8954 GND.n6221 GND.n6220 9.3005
R8955 GND.n6222 GND.n291 9.3005
R8956 GND.n6224 GND.n6223 9.3005
R8957 GND.n287 GND.n286 9.3005
R8958 GND.n6231 GND.n6230 9.3005
R8959 GND.n6232 GND.n285 9.3005
R8960 GND.n6234 GND.n6233 9.3005
R8961 GND.n281 GND.n280 9.3005
R8962 GND.n6241 GND.n6240 9.3005
R8963 GND.n6242 GND.n279 9.3005
R8964 GND.n6244 GND.n6243 9.3005
R8965 GND.n275 GND.n274 9.3005
R8966 GND.n6251 GND.n6250 9.3005
R8967 GND.n6252 GND.n273 9.3005
R8968 GND.n6254 GND.n6253 9.3005
R8969 GND.n269 GND.n268 9.3005
R8970 GND.n6261 GND.n6260 9.3005
R8971 GND.n6262 GND.n267 9.3005
R8972 GND.n6264 GND.n6263 9.3005
R8973 GND.n263 GND.n262 9.3005
R8974 GND.n6271 GND.n6270 9.3005
R8975 GND.n6272 GND.n261 9.3005
R8976 GND.n6274 GND.n6273 9.3005
R8977 GND.n257 GND.n256 9.3005
R8978 GND.n6281 GND.n6280 9.3005
R8979 GND.n6282 GND.n255 9.3005
R8980 GND.n6284 GND.n6283 9.3005
R8981 GND.n251 GND.n250 9.3005
R8982 GND.n6291 GND.n6290 9.3005
R8983 GND.n6292 GND.n249 9.3005
R8984 GND.n6294 GND.n6293 9.3005
R8985 GND.n245 GND.n244 9.3005
R8986 GND.n6301 GND.n6300 9.3005
R8987 GND.n6302 GND.n243 9.3005
R8988 GND.n6304 GND.n6303 9.3005
R8989 GND.n239 GND.n238 9.3005
R8990 GND.n6311 GND.n6310 9.3005
R8991 GND.n6312 GND.n237 9.3005
R8992 GND.n6314 GND.n6313 9.3005
R8993 GND.n233 GND.n232 9.3005
R8994 GND.n6321 GND.n6320 9.3005
R8995 GND.n6322 GND.n231 9.3005
R8996 GND.n6324 GND.n6323 9.3005
R8997 GND.n227 GND.n226 9.3005
R8998 GND.n6331 GND.n6330 9.3005
R8999 GND.n6332 GND.n225 9.3005
R9000 GND.n6335 GND.n6334 9.3005
R9001 GND.n6333 GND.n221 9.3005
R9002 GND.n6341 GND.n220 9.3005
R9003 GND.n6343 GND.n6342 9.3005
R9004 GND.n6192 GND.n309 9.3005
R9005 GND.n2435 GND.n2434 9.3005
R9006 GND.n2548 GND.n2431 9.3005
R9007 GND.n2549 GND.n2430 9.3005
R9008 GND.n2550 GND.n2429 9.3005
R9009 GND.n2428 GND.n2426 9.3005
R9010 GND.n2556 GND.n2425 9.3005
R9011 GND.n2557 GND.n2424 9.3005
R9012 GND.n2558 GND.n2423 9.3005
R9013 GND.n2422 GND.n2420 9.3005
R9014 GND.n2564 GND.n2419 9.3005
R9015 GND.n2565 GND.n2418 9.3005
R9016 GND.n2566 GND.n2417 9.3005
R9017 GND.n2416 GND.n2414 9.3005
R9018 GND.n2572 GND.n2413 9.3005
R9019 GND.n2573 GND.n2412 9.3005
R9020 GND.n2574 GND.n2411 9.3005
R9021 GND.n2410 GND.n2408 9.3005
R9022 GND.n2580 GND.n2407 9.3005
R9023 GND.n2403 GND.n2354 9.3005
R9024 GND.n2402 GND.n2401 9.3005
R9025 GND.n2357 GND.n2356 9.3005
R9026 GND.n2393 GND.n2392 9.3005
R9027 GND.n2391 GND.n2359 9.3005
R9028 GND.n2390 GND.n2389 9.3005
R9029 GND.n2361 GND.n2360 9.3005
R9030 GND.n2383 GND.n2382 9.3005
R9031 GND.n2381 GND.n2363 9.3005
R9032 GND.n2380 GND.n2379 9.3005
R9033 GND.n2365 GND.n2364 9.3005
R9034 GND.n2373 GND.n2372 9.3005
R9035 GND.n2371 GND.n2368 9.3005
R9036 GND.n2370 GND.n2369 9.3005
R9037 GND.n2542 GND.n2541 9.3005
R9038 GND.n4636 GND.n1888 9.3005
R9039 GND.n4635 GND.n1889 9.3005
R9040 GND.n4222 GND.n1890 9.3005
R9041 GND.n4224 GND.n4223 9.3005
R9042 GND.n2231 GND.n2230 9.3005
R9043 GND.n4298 GND.n4297 9.3005
R9044 GND.n4299 GND.n2229 9.3005
R9045 GND.n4303 GND.n4300 9.3005
R9046 GND.n4302 GND.n4301 9.3005
R9047 GND.n2209 GND.n2208 9.3005
R9048 GND.n4323 GND.n4322 9.3005
R9049 GND.n4324 GND.n2207 9.3005
R9050 GND.n4328 GND.n4325 9.3005
R9051 GND.n4327 GND.n4326 9.3005
R9052 GND.n2186 GND.n2185 9.3005
R9053 GND.n4348 GND.n4347 9.3005
R9054 GND.n4349 GND.n2184 9.3005
R9055 GND.n4352 GND.n4351 9.3005
R9056 GND.n4350 GND.n2153 9.3005
R9057 GND.n4428 GND.n2154 9.3005
R9058 GND.n2126 GND.n2125 9.3005
R9059 GND.n4449 GND.n4448 9.3005
R9060 GND.n4450 GND.n2124 9.3005
R9061 GND.n4454 GND.n4451 9.3005
R9062 GND.n4453 GND.n4452 9.3005
R9063 GND.n2102 GND.n2101 9.3005
R9064 GND.n4475 GND.n4474 9.3005
R9065 GND.n4476 GND.n2100 9.3005
R9066 GND.n4480 GND.n4477 9.3005
R9067 GND.n4479 GND.n4478 9.3005
R9068 GND.n2082 GND.n2081 9.3005
R9069 GND.n4504 GND.n4503 9.3005
R9070 GND.n4505 GND.n2080 9.3005
R9071 GND.n4509 GND.n4506 9.3005
R9072 GND.n4508 GND.n4507 9.3005
R9073 GND.n2060 GND.n2059 9.3005
R9074 GND.n4546 GND.n4545 9.3005
R9075 GND.n4547 GND.n2058 9.3005
R9076 GND.n4549 GND.n4548 9.3005
R9077 GND.n86 GND.n85 9.3005
R9078 GND.n6500 GND.n6499 9.3005
R9079 GND.n4637 GND.n1887 9.3005
R9080 GND.n2155 GND.n2141 9.3005
R9081 GND.n4390 GND.n2141 9.3005
R9082 GND.n3306 GND.n3305 9.3005
R9083 GND.n3307 GND.n2924 9.3005
R9084 GND.n3366 GND.n3308 9.3005
R9085 GND.n3365 GND.n3309 9.3005
R9086 GND.n3364 GND.n3310 9.3005
R9087 GND.n3313 GND.n3311 9.3005
R9088 GND.n3360 GND.n3314 9.3005
R9089 GND.n3359 GND.n3315 9.3005
R9090 GND.n3358 GND.n3316 9.3005
R9091 GND.n3319 GND.n3317 9.3005
R9092 GND.n3351 GND.n3320 9.3005
R9093 GND.n3350 GND.n3321 9.3005
R9094 GND.n3349 GND.n3322 9.3005
R9095 GND.n3325 GND.n3323 9.3005
R9096 GND.n3345 GND.n3326 9.3005
R9097 GND.n3344 GND.n3327 9.3005
R9098 GND.n3343 GND.n3328 9.3005
R9099 GND.n3331 GND.n3329 9.3005
R9100 GND.n3339 GND.n3332 9.3005
R9101 GND.n3338 GND.n3333 9.3005
R9102 GND.n3337 GND.n3335 9.3005
R9103 GND.n3334 GND.n1294 9.3005
R9104 GND.n4976 GND.n1295 9.3005
R9105 GND.n4975 GND.n1296 9.3005
R9106 GND.n4974 GND.n1297 9.3005
R9107 GND.n1318 GND.n1298 9.3005
R9108 GND.n1319 GND.n1300 9.3005
R9109 GND.n1321 GND.n1320 9.3005
R9110 GND.n1324 GND.n1323 9.3005
R9111 GND.n1325 GND.n1317 9.3005
R9112 GND.n4958 GND.n1326 9.3005
R9113 GND.n4957 GND.n1327 9.3005
R9114 GND.n4956 GND.n1328 9.3005
R9115 GND.n1351 GND.n1329 9.3005
R9116 GND.n1352 GND.n1350 9.3005
R9117 GND.n4944 GND.n1353 9.3005
R9118 GND.n4943 GND.n1354 9.3005
R9119 GND.n4942 GND.n1355 9.3005
R9120 GND.n1378 GND.n1356 9.3005
R9121 GND.n1379 GND.n1377 9.3005
R9122 GND.n4930 GND.n1380 9.3005
R9123 GND.n4929 GND.n1381 9.3005
R9124 GND.n4928 GND.n1382 9.3005
R9125 GND.n1405 GND.n1383 9.3005
R9126 GND.n1406 GND.n1404 9.3005
R9127 GND.n4916 GND.n1407 9.3005
R9128 GND.n4915 GND.n1408 9.3005
R9129 GND.n4914 GND.n1409 9.3005
R9130 GND.n3682 GND.n1410 9.3005
R9131 GND.n3684 GND.n3683 9.3005
R9132 GND.n3681 GND.n3680 9.3005
R9133 GND.n3689 GND.n3688 9.3005
R9134 GND.n3690 GND.n3679 9.3005
R9135 GND.n3700 GND.n3691 9.3005
R9136 GND.n3699 GND.n3692 9.3005
R9137 GND.n3698 GND.n3693 9.3005
R9138 GND.n3696 GND.n3695 9.3005
R9139 GND.n3694 GND.n2692 9.3005
R9140 GND.n2690 GND.n2689 9.3005
R9141 GND.n3749 GND.n3748 9.3005
R9142 GND.n3750 GND.n2688 9.3005
R9143 GND.n3752 GND.n3751 9.3005
R9144 GND.n2680 GND.n2679 9.3005
R9145 GND.n3774 GND.n3773 9.3005
R9146 GND.n3775 GND.n2678 9.3005
R9147 GND.n3786 GND.n3776 9.3005
R9148 GND.n3785 GND.n3777 9.3005
R9149 GND.n3784 GND.n3778 9.3005
R9150 GND.n3781 GND.n3780 9.3005
R9151 GND.n3779 GND.n1529 9.3005
R9152 GND.n4832 GND.n1530 9.3005
R9153 GND.n4831 GND.n1531 9.3005
R9154 GND.n4830 GND.n1532 9.3005
R9155 GND.n1575 GND.n1533 9.3005
R9156 GND.n1577 GND.n1576 9.3005
R9157 GND.n1581 GND.n1580 9.3005
R9158 GND.n1582 GND.n1574 9.3005
R9159 GND.n4805 GND.n1583 9.3005
R9160 GND.n4804 GND.n1584 9.3005
R9161 GND.n4803 GND.n1585 9.3005
R9162 GND.n1619 GND.n1586 9.3005
R9163 GND.n1622 GND.n1621 9.3005
R9164 GND.n1623 GND.n1618 9.3005
R9165 GND.n4784 GND.n1624 9.3005
R9166 GND.n4783 GND.n1625 9.3005
R9167 GND.n4782 GND.n1626 9.3005
R9168 GND.n1663 GND.n1627 9.3005
R9169 GND.n1666 GND.n1665 9.3005
R9170 GND.n1667 GND.n1662 9.3005
R9171 GND.n4763 GND.n1668 9.3005
R9172 GND.n4762 GND.n1669 9.3005
R9173 GND.n4761 GND.n1670 9.3005
R9174 GND.n1712 GND.n1671 9.3005
R9175 GND.n1714 GND.n1713 9.3005
R9176 GND.n1718 GND.n1717 9.3005
R9177 GND.n1719 GND.n1711 9.3005
R9178 GND.n4736 GND.n1720 9.3005
R9179 GND.n4735 GND.n1721 9.3005
R9180 GND.n4734 GND.n1722 9.3005
R9181 GND.n2304 GND.n1723 9.3005
R9182 GND.n2306 GND.n2305 9.3005
R9183 GND.n2310 GND.n2309 9.3005
R9184 GND.n2311 GND.n2303 9.3005
R9185 GND.n2314 GND.n2313 9.3005
R9186 GND.n2312 GND.n1760 9.3005
R9187 GND.n4708 GND.n1761 9.3005
R9188 GND.n4707 GND.n1762 9.3005
R9189 GND.n4706 GND.n1763 9.3005
R9190 GND.n1785 GND.n1764 9.3005
R9191 GND.n1786 GND.n1784 9.3005
R9192 GND.n4694 GND.n1787 9.3005
R9193 GND.n4693 GND.n1788 9.3005
R9194 GND.n4692 GND.n1789 9.3005
R9195 GND.n1811 GND.n1790 9.3005
R9196 GND.n1812 GND.n1810 9.3005
R9197 GND.n4680 GND.n1813 9.3005
R9198 GND.n4679 GND.n1814 9.3005
R9199 GND.n4678 GND.n1815 9.3005
R9200 GND.n1838 GND.n1816 9.3005
R9201 GND.n1839 GND.n1837 9.3005
R9202 GND.n4666 GND.n1840 9.3005
R9203 GND.n4665 GND.n1841 9.3005
R9204 GND.n4664 GND.n1842 9.3005
R9205 GND.n1864 GND.n1843 9.3005
R9206 GND.n1865 GND.n1863 9.3005
R9207 GND.n4652 GND.n1866 9.3005
R9208 GND.n4651 GND.n1867 9.3005
R9209 GND.n4650 GND.n1868 9.3005
R9210 GND.n1874 GND.n1869 9.3005
R9211 GND.n4644 GND.n1875 9.3005
R9212 GND.n4643 GND.n1876 9.3005
R9213 GND.n4642 GND.n1877 9.3005
R9214 GND.n4230 GND.n1878 9.3005
R9215 GND.n4233 GND.n4232 9.3005
R9216 GND.n4234 GND.n4229 9.3005
R9217 GND.n4277 GND.n4235 9.3005
R9218 GND.n4276 GND.n4236 9.3005
R9219 GND.n4275 GND.n4237 9.3005
R9220 GND.n4240 GND.n4238 9.3005
R9221 GND.n4271 GND.n4241 9.3005
R9222 GND.n4270 GND.n4242 9.3005
R9223 GND.n4269 GND.n4243 9.3005
R9224 GND.n4246 GND.n4244 9.3005
R9225 GND.n4265 GND.n4247 9.3005
R9226 GND.n4264 GND.n4248 9.3005
R9227 GND.n4263 GND.n4249 9.3005
R9228 GND.n4252 GND.n4250 9.3005
R9229 GND.n4259 GND.n4253 9.3005
R9230 GND.n4258 GND.n4254 9.3005
R9231 GND.n4257 GND.n4255 9.3005
R9232 GND.n2143 GND.n2142 9.3005
R9233 GND.n4434 GND.n4433 9.3005
R9234 GND.n4439 GND.n4436 9.3005
R9235 GND.n4438 GND.n4437 9.3005
R9236 GND.n2115 GND.n2114 9.3005
R9237 GND.n4460 GND.n4459 9.3005
R9238 GND.n4461 GND.n2113 9.3005
R9239 GND.n4465 GND.n4462 9.3005
R9240 GND.n4464 GND.n4463 9.3005
R9241 GND.n2092 GND.n2091 9.3005
R9242 GND.n4486 GND.n4485 9.3005
R9243 GND.n4487 GND.n2090 9.3005
R9244 GND.n4491 GND.n4488 9.3005
R9245 GND.n4490 GND.n4489 9.3005
R9246 GND.n2073 GND.n2072 9.3005
R9247 GND.n4515 GND.n4514 9.3005
R9248 GND.n4516 GND.n2071 9.3005
R9249 GND.n4536 GND.n4517 9.3005
R9250 GND.n4535 GND.n4518 9.3005
R9251 GND.n4534 GND.n4519 9.3005
R9252 GND.n4522 GND.n4520 9.3005
R9253 GND.n4530 GND.n4523 9.3005
R9254 GND.n4529 GND.n4524 9.3005
R9255 GND.n4528 GND.n4526 9.3005
R9256 GND.n4525 GND.n147 9.3005
R9257 GND.n6417 GND.n148 9.3005
R9258 GND.n6416 GND.n149 9.3005
R9259 GND.n6415 GND.n150 9.3005
R9260 GND.n155 GND.n151 9.3005
R9261 GND.n6409 GND.n156 9.3005
R9262 GND.n6408 GND.n157 9.3005
R9263 GND.n6407 GND.n158 9.3005
R9264 GND.n163 GND.n159 9.3005
R9265 GND.n6401 GND.n164 9.3005
R9266 GND.n6400 GND.n165 9.3005
R9267 GND.n6399 GND.n166 9.3005
R9268 GND.n171 GND.n167 9.3005
R9269 GND.n6393 GND.n172 9.3005
R9270 GND.n6392 GND.n173 9.3005
R9271 GND.n6391 GND.n174 9.3005
R9272 GND.n179 GND.n175 9.3005
R9273 GND.n6385 GND.n180 9.3005
R9274 GND.n6384 GND.n181 9.3005
R9275 GND.n6383 GND.n182 9.3005
R9276 GND.n187 GND.n183 9.3005
R9277 GND.n6377 GND.n188 9.3005
R9278 GND.n6376 GND.n189 9.3005
R9279 GND.n6375 GND.n190 9.3005
R9280 GND.n195 GND.n191 9.3005
R9281 GND.n6369 GND.n196 9.3005
R9282 GND.n6368 GND.n197 9.3005
R9283 GND.n6367 GND.n198 9.3005
R9284 GND.n203 GND.n199 9.3005
R9285 GND.n6361 GND.n204 9.3005
R9286 GND.n6360 GND.n205 9.3005
R9287 GND.n6359 GND.n206 9.3005
R9288 GND.n211 GND.n207 9.3005
R9289 GND.n6353 GND.n212 9.3005
R9290 GND.n6352 GND.n213 9.3005
R9291 GND.n6351 GND.n214 9.3005
R9292 GND.n219 GND.n215 9.3005
R9293 GND.n6345 GND.n6344 9.3005
R9294 GND.n5196 GND.n5195 9.3005
R9295 GND.n5199 GND.n1005 9.3005
R9296 GND.n5200 GND.n1004 9.3005
R9297 GND.n5203 GND.n1003 9.3005
R9298 GND.n5204 GND.n1002 9.3005
R9299 GND.n5207 GND.n1001 9.3005
R9300 GND.n5208 GND.n1000 9.3005
R9301 GND.n5211 GND.n999 9.3005
R9302 GND.n5212 GND.n998 9.3005
R9303 GND.n5215 GND.n997 9.3005
R9304 GND.n5216 GND.n996 9.3005
R9305 GND.n5219 GND.n995 9.3005
R9306 GND.n5220 GND.n994 9.3005
R9307 GND.n5223 GND.n993 9.3005
R9308 GND.n5224 GND.n992 9.3005
R9309 GND.n5227 GND.n991 9.3005
R9310 GND.n5228 GND.n990 9.3005
R9311 GND.n5231 GND.n989 9.3005
R9312 GND.n5233 GND.n986 9.3005
R9313 GND.n5236 GND.n985 9.3005
R9314 GND.n5237 GND.n984 9.3005
R9315 GND.n5240 GND.n983 9.3005
R9316 GND.n5241 GND.n982 9.3005
R9317 GND.n5244 GND.n981 9.3005
R9318 GND.n5245 GND.n980 9.3005
R9319 GND.n5248 GND.n979 9.3005
R9320 GND.n5249 GND.n978 9.3005
R9321 GND.n5252 GND.n977 9.3005
R9322 GND.n5253 GND.n976 9.3005
R9323 GND.n5256 GND.n975 9.3005
R9324 GND.n5258 GND.n974 9.3005
R9325 GND.n5259 GND.n973 9.3005
R9326 GND.n5260 GND.n972 9.3005
R9327 GND.n5261 GND.n971 9.3005
R9328 GND.n5194 GND.n1006 9.3005
R9329 GND.n1044 GND.n1043 9.3005
R9330 GND.n1045 GND.n1039 9.3005
R9331 GND.n5178 GND.n1046 9.3005
R9332 GND.n5177 GND.n1047 9.3005
R9333 GND.n5176 GND.n1048 9.3005
R9334 GND.n3145 GND.n1049 9.3005
R9335 GND.n3146 GND.n3144 9.3005
R9336 GND.n3150 GND.n3147 9.3005
R9337 GND.n3149 GND.n3148 9.3005
R9338 GND.n3029 GND.n3028 9.3005
R9339 GND.n3173 GND.n3172 9.3005
R9340 GND.n3174 GND.n3027 9.3005
R9341 GND.n3178 GND.n3175 9.3005
R9342 GND.n3177 GND.n3176 9.3005
R9343 GND.n2999 GND.n2998 9.3005
R9344 GND.n3208 GND.n3207 9.3005
R9345 GND.n3209 GND.n2997 9.3005
R9346 GND.n3213 GND.n3210 9.3005
R9347 GND.n3212 GND.n3211 9.3005
R9348 GND.n2948 GND.n2943 9.3005
R9349 GND.n2915 GND.n2914 9.3005
R9350 GND.n3375 GND.n3374 9.3005
R9351 GND.n3376 GND.n2913 9.3005
R9352 GND.n3380 GND.n3377 9.3005
R9353 GND.n3379 GND.n3378 9.3005
R9354 GND.n2893 GND.n2892 9.3005
R9355 GND.n3400 GND.n3399 9.3005
R9356 GND.n3401 GND.n2891 9.3005
R9357 GND.n3405 GND.n3402 9.3005
R9358 GND.n3404 GND.n3403 9.3005
R9359 GND.n2874 GND.n2873 9.3005
R9360 GND.n3425 GND.n3424 9.3005
R9361 GND.n3426 GND.n2872 9.3005
R9362 GND.n3430 GND.n3427 9.3005
R9363 GND.n3429 GND.n3428 9.3005
R9364 GND.n2851 GND.n2850 9.3005
R9365 GND.n3453 GND.n3452 9.3005
R9366 GND.n3454 GND.n2849 9.3005
R9367 GND.n3456 GND.n3455 9.3005
R9368 GND.n1173 GND.n1172 9.3005
R9369 GND.n5098 GND.n5097 9.3005
R9370 GND.n1041 GND.n1040 9.3005
R9371 GND.n3288 GND.n2946 9.3005
R9372 GND.n3289 GND.n3288 9.3005
R9373 GND.n5334 GND.n873 9.3005
R9374 GND.n5333 GND.n874 9.3005
R9375 GND.n5332 GND.n875 9.3005
R9376 GND.n880 GND.n876 9.3005
R9377 GND.n5326 GND.n881 9.3005
R9378 GND.n5325 GND.n882 9.3005
R9379 GND.n5324 GND.n883 9.3005
R9380 GND.n888 GND.n884 9.3005
R9381 GND.n5318 GND.n889 9.3005
R9382 GND.n5317 GND.n890 9.3005
R9383 GND.n5316 GND.n891 9.3005
R9384 GND.n896 GND.n892 9.3005
R9385 GND.n5310 GND.n897 9.3005
R9386 GND.n5309 GND.n898 9.3005
R9387 GND.n5308 GND.n899 9.3005
R9388 GND.n904 GND.n900 9.3005
R9389 GND.n5302 GND.n905 9.3005
R9390 GND.n5301 GND.n906 9.3005
R9391 GND.n5300 GND.n907 9.3005
R9392 GND.n912 GND.n908 9.3005
R9393 GND.n5294 GND.n913 9.3005
R9394 GND.n5293 GND.n914 9.3005
R9395 GND.n5292 GND.n915 9.3005
R9396 GND.n920 GND.n916 9.3005
R9397 GND.n5286 GND.n921 9.3005
R9398 GND.n5285 GND.n922 9.3005
R9399 GND.n5284 GND.n923 9.3005
R9400 GND.n928 GND.n924 9.3005
R9401 GND.n5278 GND.n929 9.3005
R9402 GND.n5277 GND.n930 9.3005
R9403 GND.n5276 GND.n931 9.3005
R9404 GND.n936 GND.n932 9.3005
R9405 GND.n5270 GND.n937 9.3005
R9406 GND.n5269 GND.n938 9.3005
R9407 GND.n5268 GND.n939 9.3005
R9408 GND.n1022 GND.n940 9.3005
R9409 GND.n1025 GND.n1024 9.3005
R9410 GND.n1026 GND.n1021 9.3005
R9411 GND.n5185 GND.n1027 9.3005
R9412 GND.n5184 GND.n1028 9.3005
R9413 GND.n5183 GND.n1029 9.3005
R9414 GND.n3119 GND.n1030 9.3005
R9415 GND.n3122 GND.n3121 9.3005
R9416 GND.n3123 GND.n3118 9.3005
R9417 GND.n3136 GND.n3124 9.3005
R9418 GND.n3135 GND.n3125 9.3005
R9419 GND.n3134 GND.n3126 9.3005
R9420 GND.n3128 GND.n3127 9.3005
R9421 GND.n3130 GND.n3129 9.3005
R9422 GND.n3016 GND.n3015 9.3005
R9423 GND.n3184 GND.n3183 9.3005
R9424 GND.n3185 GND.n3014 9.3005
R9425 GND.n3189 GND.n3186 9.3005
R9426 GND.n3188 GND.n3187 9.3005
R9427 GND.n2988 GND.n2987 9.3005
R9428 GND.n3219 GND.n3218 9.3005
R9429 GND.n3220 GND.n2986 9.3005
R9430 GND.n3225 GND.n3221 9.3005
R9431 GND.n3224 GND.n3222 9.3005
R9432 GND.n872 GND.n871 9.3005
R9433 GND.n5341 GND.n866 9.3005
R9434 GND.n5342 GND.n865 9.3005
R9435 GND.n864 GND.n860 9.3005
R9436 GND.n5348 GND.n859 9.3005
R9437 GND.n5349 GND.n858 9.3005
R9438 GND.n5350 GND.n857 9.3005
R9439 GND.n856 GND.n852 9.3005
R9440 GND.n5356 GND.n851 9.3005
R9441 GND.n5357 GND.n850 9.3005
R9442 GND.n5358 GND.n849 9.3005
R9443 GND.n848 GND.n844 9.3005
R9444 GND.n5364 GND.n843 9.3005
R9445 GND.n5365 GND.n842 9.3005
R9446 GND.n5366 GND.n841 9.3005
R9447 GND.n840 GND.n836 9.3005
R9448 GND.n5372 GND.n835 9.3005
R9449 GND.n5373 GND.n834 9.3005
R9450 GND.n5374 GND.n833 9.3005
R9451 GND.n832 GND.n828 9.3005
R9452 GND.n5380 GND.n827 9.3005
R9453 GND.n5381 GND.n826 9.3005
R9454 GND.n5382 GND.n825 9.3005
R9455 GND.n824 GND.n820 9.3005
R9456 GND.n5388 GND.n819 9.3005
R9457 GND.n5389 GND.n818 9.3005
R9458 GND.n5390 GND.n817 9.3005
R9459 GND.n816 GND.n812 9.3005
R9460 GND.n5396 GND.n811 9.3005
R9461 GND.n5397 GND.n810 9.3005
R9462 GND.n5398 GND.n809 9.3005
R9463 GND.n808 GND.n804 9.3005
R9464 GND.n5404 GND.n803 9.3005
R9465 GND.n5405 GND.n802 9.3005
R9466 GND.n5406 GND.n801 9.3005
R9467 GND.n800 GND.n796 9.3005
R9468 GND.n5412 GND.n795 9.3005
R9469 GND.n5413 GND.n794 9.3005
R9470 GND.n5414 GND.n793 9.3005
R9471 GND.n792 GND.n788 9.3005
R9472 GND.n5420 GND.n787 9.3005
R9473 GND.n5421 GND.n786 9.3005
R9474 GND.n5422 GND.n785 9.3005
R9475 GND.n784 GND.n780 9.3005
R9476 GND.n5428 GND.n779 9.3005
R9477 GND.n5429 GND.n778 9.3005
R9478 GND.n5430 GND.n777 9.3005
R9479 GND.n776 GND.n772 9.3005
R9480 GND.n5436 GND.n771 9.3005
R9481 GND.n5437 GND.n770 9.3005
R9482 GND.n5438 GND.n769 9.3005
R9483 GND.n768 GND.n764 9.3005
R9484 GND.n5444 GND.n763 9.3005
R9485 GND.n5445 GND.n762 9.3005
R9486 GND.n5446 GND.n761 9.3005
R9487 GND.n760 GND.n756 9.3005
R9488 GND.n5452 GND.n755 9.3005
R9489 GND.n5453 GND.n754 9.3005
R9490 GND.n5454 GND.n753 9.3005
R9491 GND.n749 GND.n748 9.3005
R9492 GND.n5461 GND.n5460 9.3005
R9493 GND.n5340 GND.n867 9.3005
R9494 GND.n4220 GND.n4219 9.3005
R9495 GND.n4221 GND.n2242 9.3005
R9496 GND.n4283 GND.n4282 9.3005
R9497 GND.n4284 GND.n2240 9.3005
R9498 GND.n4287 GND.n4286 9.3005
R9499 GND.n4285 GND.n2241 9.3005
R9500 GND.n2220 GND.n2219 9.3005
R9501 GND.n4308 GND.n4307 9.3005
R9502 GND.n4309 GND.n2217 9.3005
R9503 GND.n4312 GND.n4311 9.3005
R9504 GND.n4310 GND.n2218 9.3005
R9505 GND.n2198 GND.n2197 9.3005
R9506 GND.n4333 GND.n4332 9.3005
R9507 GND.n4334 GND.n2195 9.3005
R9508 GND.n4337 GND.n4336 9.3005
R9509 GND.n4335 GND.n2196 9.3005
R9510 GND.n2175 GND.n2174 9.3005
R9511 GND.n4357 GND.n4356 9.3005
R9512 GND.n4358 GND.n2173 9.3005
R9513 GND.n4360 GND.n4359 9.3005
R9514 GND.n4364 GND.n2172 9.3005
R9515 GND.n4366 GND.n4365 9.3005
R9516 GND.n4367 GND.n2171 9.3005
R9517 GND.n4369 GND.n4368 9.3005
R9518 GND.n46 GND.n44 9.3005
R9519 GND.n4218 GND.n2243 9.3005
R9520 GND.n6542 GND.n6541 9.3005
R9521 GND.n6540 GND.n45 9.3005
R9522 GND.n6539 GND.n6538 9.3005
R9523 GND.n6537 GND.n50 9.3005
R9524 GND.n6536 GND.n6535 9.3005
R9525 GND.n6534 GND.n51 9.3005
R9526 GND.n6533 GND.n6532 9.3005
R9527 GND.n6531 GND.n55 9.3005
R9528 GND.n6530 GND.n6529 9.3005
R9529 GND.n6528 GND.n56 9.3005
R9530 GND.n6527 GND.n6526 9.3005
R9531 GND.n6525 GND.n60 9.3005
R9532 GND.n6524 GND.n6523 9.3005
R9533 GND.n6522 GND.n61 9.3005
R9534 GND.n6521 GND.n6520 9.3005
R9535 GND.n6519 GND.n65 9.3005
R9536 GND.n6518 GND.n6517 9.3005
R9537 GND.n6516 GND.n66 9.3005
R9538 GND.n6515 GND.n6514 9.3005
R9539 GND.n6513 GND.n70 9.3005
R9540 GND.n6512 GND.n6511 9.3005
R9541 GND.n6510 GND.n71 9.3005
R9542 GND.n6509 GND.n6508 9.3005
R9543 GND.n6507 GND.n75 9.3005
R9544 GND.n6506 GND.n6505 9.3005
R9545 GND.n6504 GND.n76 9.3005
R9546 GND.n2047 GND.n1998 9.3005
R9547 GND.n2046 GND.n2045 9.3005
R9548 GND.n2044 GND.n2002 9.3005
R9549 GND.n2043 GND.n2042 9.3005
R9550 GND.n2041 GND.n2003 9.3005
R9551 GND.n2040 GND.n2039 9.3005
R9552 GND.n2038 GND.n2008 9.3005
R9553 GND.n2037 GND.n2036 9.3005
R9554 GND.n2035 GND.n2009 9.3005
R9555 GND.n2034 GND.n2033 9.3005
R9556 GND.n2032 GND.n2014 9.3005
R9557 GND.n2031 GND.n2030 9.3005
R9558 GND.n2029 GND.n2015 9.3005
R9559 GND.n2028 GND.n2027 9.3005
R9560 GND.n2026 GND.n2023 9.3005
R9561 GND.n2025 GND.n2024 9.3005
R9562 GND.n2049 GND.n2048 9.3005
R9563 GND.n6496 GND.n87 9.3005
R9564 GND.n6495 GND.n6494 9.3005
R9565 GND.n6493 GND.n90 9.3005
R9566 GND.n6492 GND.n6491 9.3005
R9567 GND.n6490 GND.n91 9.3005
R9568 GND.n6489 GND.n6488 9.3005
R9569 GND.n6487 GND.n95 9.3005
R9570 GND.n6486 GND.n6485 9.3005
R9571 GND.n6484 GND.n96 9.3005
R9572 GND.n6483 GND.n6482 9.3005
R9573 GND.n6481 GND.n100 9.3005
R9574 GND.n6480 GND.n6479 9.3005
R9575 GND.n6478 GND.n101 9.3005
R9576 GND.n6477 GND.n6476 9.3005
R9577 GND.n6475 GND.n105 9.3005
R9578 GND.n6474 GND.n6473 9.3005
R9579 GND.n6472 GND.n106 9.3005
R9580 GND.n6471 GND.n6470 9.3005
R9581 GND.n6469 GND.n113 9.3005
R9582 GND.n6468 GND.n6467 9.3005
R9583 GND.n6466 GND.n114 9.3005
R9584 GND.n6465 GND.n6464 9.3005
R9585 GND.n6463 GND.n118 9.3005
R9586 GND.n6462 GND.n6461 9.3005
R9587 GND.n6460 GND.n119 9.3005
R9588 GND.n6459 GND.n6458 9.3005
R9589 GND.n6457 GND.n123 9.3005
R9590 GND.n6456 GND.n6455 9.3005
R9591 GND.n6454 GND.n124 9.3005
R9592 GND.n6453 GND.n6452 9.3005
R9593 GND.n6451 GND.n128 9.3005
R9594 GND.n6450 GND.n6449 9.3005
R9595 GND.n6448 GND.n129 9.3005
R9596 GND.n6447 GND.n134 9.3005
R9597 GND.n6498 GND.n6497 9.3005
R9598 GND.n1900 GND.n1898 9.3005
R9599 GND.n4631 GND.n4630 9.3005
R9600 GND.n1901 GND.n1899 9.3005
R9601 GND.n4626 GND.n1906 9.3005
R9602 GND.n4625 GND.n1907 9.3005
R9603 GND.n4624 GND.n1908 9.3005
R9604 GND.n4291 GND.n1909 9.3005
R9605 GND.n4620 GND.n1914 9.3005
R9606 GND.n4619 GND.n1915 9.3005
R9607 GND.n4618 GND.n1916 9.3005
R9608 GND.n4318 GND.n1917 9.3005
R9609 GND.n4614 GND.n1922 9.3005
R9610 GND.n4613 GND.n1923 9.3005
R9611 GND.n4612 GND.n1924 9.3005
R9612 GND.n2192 GND.n1925 9.3005
R9613 GND.n4608 GND.n1930 9.3005
R9614 GND.n4607 GND.n1931 9.3005
R9615 GND.n4606 GND.n1932 9.3005
R9616 GND.n2180 GND.n1933 9.3005
R9617 GND.n4602 GND.n1938 9.3005
R9618 GND.n4601 GND.n1939 9.3005
R9619 GND.n4600 GND.n1940 9.3005
R9620 GND.n2162 GND.n1941 9.3005
R9621 GND.n4596 GND.n1946 9.3005
R9622 GND.n4595 GND.n1947 9.3005
R9623 GND.n4594 GND.n1948 9.3005
R9624 GND.n4404 GND.n1949 9.3005
R9625 GND.n4590 GND.n1954 9.3005
R9626 GND.n4589 GND.n1955 9.3005
R9627 GND.n4588 GND.n1956 9.3005
R9628 GND.n2131 GND.n1957 9.3005
R9629 GND.n4584 GND.n1962 9.3005
R9630 GND.n4583 GND.n1963 9.3005
R9631 GND.n4582 GND.n1964 9.3005
R9632 GND.n2108 GND.n1965 9.3005
R9633 GND.n4578 GND.n1970 9.3005
R9634 GND.n4577 GND.n1971 9.3005
R9635 GND.n4576 GND.n1972 9.3005
R9636 GND.n2096 GND.n1973 9.3005
R9637 GND.n4572 GND.n1978 9.3005
R9638 GND.n4571 GND.n1979 9.3005
R9639 GND.n4570 GND.n1980 9.3005
R9640 GND.n4498 GND.n1981 9.3005
R9641 GND.n4566 GND.n1986 9.3005
R9642 GND.n4565 GND.n1987 9.3005
R9643 GND.n4564 GND.n1988 9.3005
R9644 GND.n4541 GND.n1989 9.3005
R9645 GND.n4560 GND.n1994 9.3005
R9646 GND.n4559 GND.n1995 9.3005
R9647 GND.n4558 GND.n1996 9.3005
R9648 GND.n2051 GND.n1997 9.3005
R9649 GND.n2438 GND.n2436 9.3005
R9650 GND.n1902 GND.n1900 9.3005
R9651 GND.n4630 GND.n4629 9.3005
R9652 GND.n4628 GND.n1901 9.3005
R9653 GND.n4627 GND.n4626 9.3005
R9654 GND.n4625 GND.n1905 9.3005
R9655 GND.n4624 GND.n4623 9.3005
R9656 GND.n4622 GND.n1909 9.3005
R9657 GND.n4621 GND.n4620 9.3005
R9658 GND.n4619 GND.n1913 9.3005
R9659 GND.n4618 GND.n4617 9.3005
R9660 GND.n4616 GND.n1917 9.3005
R9661 GND.n4615 GND.n4614 9.3005
R9662 GND.n4613 GND.n1921 9.3005
R9663 GND.n4612 GND.n4611 9.3005
R9664 GND.n4610 GND.n1925 9.3005
R9665 GND.n4609 GND.n4608 9.3005
R9666 GND.n4607 GND.n1929 9.3005
R9667 GND.n4606 GND.n4605 9.3005
R9668 GND.n4604 GND.n1933 9.3005
R9669 GND.n4603 GND.n4602 9.3005
R9670 GND.n4601 GND.n1937 9.3005
R9671 GND.n4600 GND.n4599 9.3005
R9672 GND.n4598 GND.n1941 9.3005
R9673 GND.n4597 GND.n4596 9.3005
R9674 GND.n4595 GND.n1945 9.3005
R9675 GND.n4594 GND.n4593 9.3005
R9676 GND.n4592 GND.n1949 9.3005
R9677 GND.n4591 GND.n4590 9.3005
R9678 GND.n4589 GND.n1953 9.3005
R9679 GND.n4588 GND.n4587 9.3005
R9680 GND.n4586 GND.n1957 9.3005
R9681 GND.n4585 GND.n4584 9.3005
R9682 GND.n4583 GND.n1961 9.3005
R9683 GND.n4582 GND.n4581 9.3005
R9684 GND.n4580 GND.n1965 9.3005
R9685 GND.n4579 GND.n4578 9.3005
R9686 GND.n4577 GND.n1969 9.3005
R9687 GND.n4576 GND.n4575 9.3005
R9688 GND.n4574 GND.n1973 9.3005
R9689 GND.n4573 GND.n4572 9.3005
R9690 GND.n4571 GND.n1977 9.3005
R9691 GND.n4570 GND.n4569 9.3005
R9692 GND.n4568 GND.n1981 9.3005
R9693 GND.n4567 GND.n4566 9.3005
R9694 GND.n4565 GND.n1985 9.3005
R9695 GND.n4564 GND.n4563 9.3005
R9696 GND.n4562 GND.n1989 9.3005
R9697 GND.n4561 GND.n4560 9.3005
R9698 GND.n4559 GND.n1993 9.3005
R9699 GND.n4558 GND.n4557 9.3005
R9700 GND.n4556 GND.n2051 9.3005
R9701 GND.n2438 GND.n2437 9.3005
R9702 GND.n2531 GND.n2442 9.3005
R9703 GND.n2533 GND.n2532 9.3005
R9704 GND.n2440 GND.n2439 9.3005
R9705 GND.n2539 GND.n2538 9.3005
R9706 GND.n2523 GND.n2522 9.3005
R9707 GND.n2451 GND.n2450 9.3005
R9708 GND.n2517 GND.n2516 9.3005
R9709 GND.n2515 GND.n2514 9.3005
R9710 GND.n2467 GND.n2466 9.3005
R9711 GND.n2509 GND.n2508 9.3005
R9712 GND.n2507 GND.n2506 9.3005
R9713 GND.n2480 GND.n2479 9.3005
R9714 GND.n2496 GND.n2495 9.3005
R9715 GND.n2494 GND.n2493 9.3005
R9716 GND.n2249 GND.n2247 9.3005
R9717 GND.n2525 GND.n2524 9.3005
R9718 GND.n2505 GND.n2504 9.3005
R9719 GND.n2474 GND.n2473 9.3005
R9720 GND.n2511 GND.n2510 9.3005
R9721 GND.n2513 GND.n2512 9.3005
R9722 GND.n2460 GND.n2459 9.3005
R9723 GND.n2519 GND.n2518 9.3005
R9724 GND.n2521 GND.n2520 9.3005
R9725 GND.n2452 GND.n2448 9.3005
R9726 GND.n2526 GND.n2447 9.3005
R9727 GND.n2528 GND.n2527 9.3005
R9728 GND.n2530 GND.n2529 9.3005
R9729 GND.n2503 GND.n2497 9.3005
R9730 GND.n2485 GND.n2484 9.3005
R9731 GND.n4216 GND.n4215 9.3005
R9732 GND.n4214 GND.n2248 9.3005
R9733 GND.n4213 GND.n4212 9.3005
R9734 GND.n4211 GND.n2254 9.3005
R9735 GND.n4210 GND.n4209 9.3005
R9736 GND.n4208 GND.n2255 9.3005
R9737 GND.n4207 GND.n4206 9.3005
R9738 GND.n4205 GND.n2262 9.3005
R9739 GND.n4204 GND.n4203 9.3005
R9740 GND.n4202 GND.n2263 9.3005
R9741 GND.n4201 GND.n4200 9.3005
R9742 GND.n4199 GND.n2270 9.3005
R9743 GND.n4198 GND.n4197 9.3005
R9744 GND.n4196 GND.n2271 9.3005
R9745 GND.n4195 GND.n4194 9.3005
R9746 GND.n4193 GND.n2280 9.3005
R9747 GND.n4192 GND.n4191 9.3005
R9748 GND.n3520 GND.n2831 9.3005
R9749 GND.n3524 GND.n3523 9.3005
R9750 GND.n3525 GND.n2830 9.3005
R9751 GND.n3527 GND.n3526 9.3005
R9752 GND.n3530 GND.n2829 9.3005
R9753 GND.n3532 GND.n3531 9.3005
R9754 GND.n3533 GND.n2828 9.3005
R9755 GND.n3535 GND.n3534 9.3005
R9756 GND.n3536 GND.n2825 9.3005
R9757 GND.n3540 GND.n3539 9.3005
R9758 GND.n3541 GND.n2822 9.3005
R9759 GND.n3543 GND.n3542 9.3005
R9760 GND.n3544 GND.n2821 9.3005
R9761 GND.n3548 GND.n3547 9.3005
R9762 GND.n3549 GND.n2820 9.3005
R9763 GND.n3551 GND.n3550 9.3005
R9764 GND.n3554 GND.n2819 9.3005
R9765 GND.n3556 GND.n3555 9.3005
R9766 GND.n3557 GND.n2818 9.3005
R9767 GND.n3559 GND.n3558 9.3005
R9768 GND.n2711 GND.n2710 9.3005
R9769 GND.n3659 GND.n3658 9.3005
R9770 GND.n3660 GND.n2709 9.3005
R9771 GND.n3662 GND.n3661 9.3005
R9772 GND.n2705 GND.n2704 9.3005
R9773 GND.n3706 GND.n3705 9.3005
R9774 GND.n3707 GND.n2703 9.3005
R9775 GND.n3709 GND.n3708 9.3005
R9776 GND.n2699 GND.n2697 9.3005
R9777 GND.n3741 GND.n3740 9.3005
R9778 GND.n3739 GND.n2698 9.3005
R9779 GND.n3738 GND.n3737 9.3005
R9780 GND.n3736 GND.n2700 9.3005
R9781 GND.n3735 GND.n3734 9.3005
R9782 GND.n3733 GND.n3729 9.3005
R9783 GND.n3732 GND.n3731 9.3005
R9784 GND.n2673 GND.n2672 9.3005
R9785 GND.n3795 GND.n3794 9.3005
R9786 GND.n3796 GND.n2670 9.3005
R9787 GND.n3807 GND.n3806 9.3005
R9788 GND.n3805 GND.n2671 9.3005
R9789 GND.n3804 GND.n3803 9.3005
R9790 GND.n3802 GND.n3798 9.3005
R9791 GND.n3797 GND.n2662 9.3005
R9792 GND.n2661 GND.n2660 9.3005
R9793 GND.n3843 GND.n3842 9.3005
R9794 GND.n3844 GND.n2658 9.3005
R9795 GND.n3850 GND.n3849 9.3005
R9796 GND.n3848 GND.n2659 9.3005
R9797 GND.n3847 GND.n3846 9.3005
R9798 GND.n2649 GND.n2648 9.3005
R9799 GND.n3879 GND.n3878 9.3005
R9800 GND.n3880 GND.n2646 9.3005
R9801 GND.n3903 GND.n3902 9.3005
R9802 GND.n3901 GND.n2647 9.3005
R9803 GND.n3900 GND.n3899 9.3005
R9804 GND.n3898 GND.n3881 9.3005
R9805 GND.n3897 GND.n3896 9.3005
R9806 GND.n3895 GND.n3886 9.3005
R9807 GND.n3894 GND.n3893 9.3005
R9808 GND.n3892 GND.n3887 9.3005
R9809 GND.n3891 GND.n3890 9.3005
R9810 GND.n3889 GND.n2633 9.3005
R9811 GND.n2632 GND.n2631 9.3005
R9812 GND.n3968 GND.n3967 9.3005
R9813 GND.n3969 GND.n2629 9.3005
R9814 GND.n3971 GND.n3970 9.3005
R9815 GND.n3972 GND.n2628 9.3005
R9816 GND.n3975 GND.n3974 9.3005
R9817 GND.n3976 GND.n2627 9.3005
R9818 GND.n3978 GND.n3977 9.3005
R9819 GND.n2611 GND.n2610 9.3005
R9820 GND.n4001 GND.n4000 9.3005
R9821 GND.n4002 GND.n2609 9.3005
R9822 GND.n4005 GND.n4004 9.3005
R9823 GND.n4003 GND.n2301 9.3005
R9824 GND.n4145 GND.n2300 9.3005
R9825 GND.n4147 GND.n4146 9.3005
R9826 GND.n4148 GND.n2295 9.3005
R9827 GND.n4150 GND.n4149 9.3005
R9828 GND.n4151 GND.n2294 9.3005
R9829 GND.n4155 GND.n4154 9.3005
R9830 GND.n4156 GND.n2293 9.3005
R9831 GND.n4158 GND.n4157 9.3005
R9832 GND.n4161 GND.n2292 9.3005
R9833 GND.n4163 GND.n4162 9.3005
R9834 GND.n4164 GND.n2291 9.3005
R9835 GND.n4166 GND.n4165 9.3005
R9836 GND.n4167 GND.n2287 9.3005
R9837 GND.n4171 GND.n4170 9.3005
R9838 GND.n4172 GND.n2284 9.3005
R9839 GND.n4174 GND.n4173 9.3005
R9840 GND.n4175 GND.n2283 9.3005
R9841 GND.n4179 GND.n4178 9.3005
R9842 GND.n4180 GND.n2282 9.3005
R9843 GND.n4182 GND.n4181 9.3005
R9844 GND.n4185 GND.n2281 9.3005
R9845 GND.n4187 GND.n4186 9.3005
R9846 GND.n3519 GND.n3518 9.3005
R9847 GND.n3514 GND.n2832 9.3005
R9848 GND.n3511 GND.n3510 9.3005
R9849 GND.n3509 GND.n2835 9.3005
R9850 GND.n3508 GND.n3507 9.3005
R9851 GND.n3504 GND.n2836 9.3005
R9852 GND.n3501 GND.n3500 9.3005
R9853 GND.n3499 GND.n2837 9.3005
R9854 GND.n3498 GND.n3497 9.3005
R9855 GND.n3494 GND.n2838 9.3005
R9856 GND.n3491 GND.n3490 9.3005
R9857 GND.n3489 GND.n2839 9.3005
R9858 GND.n3488 GND.n3487 9.3005
R9859 GND.n3484 GND.n2840 9.3005
R9860 GND.n3481 GND.n3480 9.3005
R9861 GND.n3479 GND.n2841 9.3005
R9862 GND.n3478 GND.n3477 9.3005
R9863 GND.n3517 GND.n3516 9.3005
R9864 GND.n3246 GND.n2977 9.3005
R9865 GND.n3248 GND.n3247 9.3005
R9866 GND.n2933 GND.n2932 9.3005
R9867 GND.n3295 GND.n3294 9.3005
R9868 GND.n3296 GND.n2930 9.3005
R9869 GND.n3299 GND.n3298 9.3005
R9870 GND.n3297 GND.n2931 9.3005
R9871 GND.n2905 GND.n2904 9.3005
R9872 GND.n3385 GND.n3384 9.3005
R9873 GND.n3386 GND.n2902 9.3005
R9874 GND.n3389 GND.n3388 9.3005
R9875 GND.n3387 GND.n2903 9.3005
R9876 GND.n2885 GND.n2884 9.3005
R9877 GND.n3410 GND.n3409 9.3005
R9878 GND.n3411 GND.n2882 9.3005
R9879 GND.n3414 GND.n3413 9.3005
R9880 GND.n3412 GND.n2883 9.3005
R9881 GND.n2863 GND.n2862 9.3005
R9882 GND.n3435 GND.n3434 9.3005
R9883 GND.n3436 GND.n2860 9.3005
R9884 GND.n3445 GND.n3444 9.3005
R9885 GND.n3443 GND.n2861 9.3005
R9886 GND.n3442 GND.n3441 9.3005
R9887 GND.n3437 GND.n2843 9.3005
R9888 GND.n3465 GND.n2842 9.3005
R9889 GND.n3467 GND.n3466 9.3005
R9890 GND.n3474 GND.n3473 9.3005
R9891 GND.n3472 GND.n3469 9.3005
R9892 GND.n1271 GND.n1270 9.3005
R9893 GND.n5011 GND.n5010 9.3005
R9894 GND.n5013 GND.n5012 9.3005
R9895 GND.n1261 GND.n1260 9.3005
R9896 GND.n5019 GND.n5018 9.3005
R9897 GND.n5021 GND.n5020 9.3005
R9898 GND.n1252 GND.n1249 9.3005
R9899 GND.n5027 GND.n5026 9.3005
R9900 GND.n1250 GND.n1230 9.3005
R9901 GND.n5033 GND.n5032 9.3005
R9902 GND.n5038 GND.n5037 9.3005
R9903 GND.n5036 GND.n5035 9.3005
R9904 GND.n5034 GND.n1228 9.3005
R9905 GND.n1282 GND.n1229 9.3005
R9906 GND.n1253 GND.n1251 9.3005
R9907 GND.n5025 GND.n5024 9.3005
R9908 GND.n5023 GND.n5022 9.3005
R9909 GND.n1257 GND.n1256 9.3005
R9910 GND.n5017 GND.n5016 9.3005
R9911 GND.n5015 GND.n5014 9.3005
R9912 GND.n1265 GND.n1264 9.3005
R9913 GND.n5009 GND.n5008 9.3005
R9914 GND.n5007 GND.n1275 9.3005
R9915 GND.n5042 GND.n1220 9.3005
R9916 GND.n5041 GND.n5040 9.3005
R9917 GND.n5039 GND.n1224 9.3005
R9918 GND.n5044 GND.n5043 9.3005
R9919 GND.n5076 GND.n1188 9.3005
R9920 GND.n5078 GND.n5077 9.3005
R9921 GND.n5079 GND.n1187 9.3005
R9922 GND.n5081 GND.n5080 9.3005
R9923 GND.n5082 GND.n1183 9.3005
R9924 GND.n5084 GND.n5083 9.3005
R9925 GND.n5085 GND.n1182 9.3005
R9926 GND.n5087 GND.n5086 9.3005
R9927 GND.n5088 GND.n1178 9.3005
R9928 GND.n5090 GND.n5089 9.3005
R9929 GND.n5091 GND.n1177 9.3005
R9930 GND.n5093 GND.n5092 9.3005
R9931 GND.n5094 GND.n1174 9.3005
R9932 GND.n5096 GND.n5095 9.3005
R9933 GND.n5072 GND.n1197 9.3005
R9934 GND.n5071 GND.n5070 9.3005
R9935 GND.n5069 GND.n1198 9.3005
R9936 GND.n5068 GND.n5067 9.3005
R9937 GND.n5066 GND.n1202 9.3005
R9938 GND.n5065 GND.n5064 9.3005
R9939 GND.n5063 GND.n1203 9.3005
R9940 GND.n5062 GND.n5061 9.3005
R9941 GND.n5060 GND.n1207 9.3005
R9942 GND.n5059 GND.n5058 9.3005
R9943 GND.n5057 GND.n1208 9.3005
R9944 GND.n5056 GND.n5055 9.3005
R9945 GND.n5054 GND.n1212 9.3005
R9946 GND.n5053 GND.n5052 9.3005
R9947 GND.n5051 GND.n1213 9.3005
R9948 GND.n5050 GND.n5049 9.3005
R9949 GND.n5048 GND.n1219 9.3005
R9950 GND.n5047 GND.n5046 9.3005
R9951 GND.n5074 GND.n5073 9.3005
R9952 GND.n1068 GND.n1067 9.3005
R9953 GND.n1070 GND.n1062 9.3005
R9954 GND.n1072 GND.n1071 9.3005
R9955 GND.n1059 GND.n1057 9.3005
R9956 GND.n5172 GND.n5171 9.3005
R9957 GND.n1060 GND.n1058 9.3005
R9958 GND.n5167 GND.n1078 9.3005
R9959 GND.n5166 GND.n1079 9.3005
R9960 GND.n5165 GND.n1080 9.3005
R9961 GND.n3035 GND.n1081 9.3005
R9962 GND.n5161 GND.n1086 9.3005
R9963 GND.n5160 GND.n1087 9.3005
R9964 GND.n5159 GND.n1088 9.3005
R9965 GND.n3022 GND.n1089 9.3005
R9966 GND.n5155 GND.n1094 9.3005
R9967 GND.n5154 GND.n1095 9.3005
R9968 GND.n5153 GND.n1096 9.3005
R9969 GND.n2993 GND.n1097 9.3005
R9970 GND.n5149 GND.n1102 9.3005
R9971 GND.n5148 GND.n1103 9.3005
R9972 GND.n5147 GND.n1104 9.3005
R9973 GND.n2956 GND.n1105 9.3005
R9974 GND.n5143 GND.n1110 9.3005
R9975 GND.n5142 GND.n1111 9.3005
R9976 GND.n5141 GND.n1112 9.3005
R9977 GND.n3265 GND.n1113 9.3005
R9978 GND.n5137 GND.n1118 9.3005
R9979 GND.n5136 GND.n1119 9.3005
R9980 GND.n5135 GND.n1120 9.3005
R9981 GND.n2937 GND.n1121 9.3005
R9982 GND.n5131 GND.n1126 9.3005
R9983 GND.n5130 GND.n1127 9.3005
R9984 GND.n5129 GND.n1128 9.3005
R9985 GND.n2908 GND.n1129 9.3005
R9986 GND.n5125 GND.n1134 9.3005
R9987 GND.n5124 GND.n1135 9.3005
R9988 GND.n5123 GND.n1136 9.3005
R9989 GND.n3393 GND.n1137 9.3005
R9990 GND.n5119 GND.n1142 9.3005
R9991 GND.n5118 GND.n1143 9.3005
R9992 GND.n5117 GND.n1144 9.3005
R9993 GND.n3420 GND.n1145 9.3005
R9994 GND.n5113 GND.n1150 9.3005
R9995 GND.n5112 GND.n1151 9.3005
R9996 GND.n5111 GND.n1152 9.3005
R9997 GND.n2857 GND.n1153 9.3005
R9998 GND.n5107 GND.n1158 9.3005
R9999 GND.n5106 GND.n1159 9.3005
R10000 GND.n5105 GND.n1160 9.3005
R10001 GND.n3461 GND.n1161 9.3005
R10002 GND.n3460 GND.n1164 9.3005
R10003 GND.n1013 GND.n1009 9.3005
R10004 GND.n1067 GND.n1066 9.3005
R10005 GND.n1062 GND.n1061 9.3005
R10006 GND.n1073 GND.n1072 9.3005
R10007 GND.n1074 GND.n1059 9.3005
R10008 GND.n5171 GND.n5170 9.3005
R10009 GND.n5169 GND.n1060 9.3005
R10010 GND.n5168 GND.n5167 9.3005
R10011 GND.n5166 GND.n1077 9.3005
R10012 GND.n5165 GND.n5164 9.3005
R10013 GND.n5163 GND.n1081 9.3005
R10014 GND.n5162 GND.n5161 9.3005
R10015 GND.n5160 GND.n1085 9.3005
R10016 GND.n5159 GND.n5158 9.3005
R10017 GND.n5157 GND.n1089 9.3005
R10018 GND.n5156 GND.n5155 9.3005
R10019 GND.n5154 GND.n1093 9.3005
R10020 GND.n5153 GND.n5152 9.3005
R10021 GND.n5151 GND.n1097 9.3005
R10022 GND.n5150 GND.n5149 9.3005
R10023 GND.n5148 GND.n1101 9.3005
R10024 GND.n5147 GND.n5146 9.3005
R10025 GND.n5145 GND.n1105 9.3005
R10026 GND.n5144 GND.n5143 9.3005
R10027 GND.n5142 GND.n1109 9.3005
R10028 GND.n5141 GND.n5140 9.3005
R10029 GND.n5139 GND.n1113 9.3005
R10030 GND.n5138 GND.n5137 9.3005
R10031 GND.n5136 GND.n1117 9.3005
R10032 GND.n5135 GND.n5134 9.3005
R10033 GND.n5133 GND.n1121 9.3005
R10034 GND.n5132 GND.n5131 9.3005
R10035 GND.n5130 GND.n1125 9.3005
R10036 GND.n5129 GND.n5128 9.3005
R10037 GND.n5127 GND.n1129 9.3005
R10038 GND.n5126 GND.n5125 9.3005
R10039 GND.n5124 GND.n1133 9.3005
R10040 GND.n5123 GND.n5122 9.3005
R10041 GND.n5121 GND.n1137 9.3005
R10042 GND.n5120 GND.n5119 9.3005
R10043 GND.n5118 GND.n1141 9.3005
R10044 GND.n5117 GND.n5116 9.3005
R10045 GND.n5115 GND.n1145 9.3005
R10046 GND.n5114 GND.n5113 9.3005
R10047 GND.n5112 GND.n1149 9.3005
R10048 GND.n5111 GND.n5110 9.3005
R10049 GND.n5109 GND.n1153 9.3005
R10050 GND.n5108 GND.n5107 9.3005
R10051 GND.n5106 GND.n1157 9.3005
R10052 GND.n5105 GND.n5104 9.3005
R10053 GND.n5103 GND.n1161 9.3005
R10054 GND.n5102 GND.n1164 9.3005
R10055 GND.n1063 GND.n1009 9.3005
R10056 GND.n3095 GND.n3094 9.3005
R10057 GND.n3093 GND.n3056 9.3005
R10058 GND.n3092 GND.n3091 9.3005
R10059 GND.n3088 GND.n3059 9.3005
R10060 GND.n3087 GND.n3086 9.3005
R10061 GND.n3085 GND.n3060 9.3005
R10062 GND.n3084 GND.n3083 9.3005
R10063 GND.n3080 GND.n3063 9.3005
R10064 GND.n3079 GND.n3078 9.3005
R10065 GND.n3077 GND.n3064 9.3005
R10066 GND.n3076 GND.n3075 9.3005
R10067 GND.n3072 GND.n3067 9.3005
R10068 GND.n3071 GND.n3070 9.3005
R10069 GND.n1011 GND.n1010 9.3005
R10070 GND.n5192 GND.n5191 9.3005
R10071 GND.n3096 GND.n3052 9.3005
R10072 GND.n3098 GND.n3097 9.3005
R10073 GND.n3101 GND.n3049 9.3005
R10074 GND.n3103 GND.n3102 9.3005
R10075 GND.n3104 GND.n3048 9.3005
R10076 GND.n3110 GND.n3109 9.3005
R10077 GND.n3111 GND.n3047 9.3005
R10078 GND.n3113 GND.n3112 9.3005
R10079 GND.n3041 GND.n3040 9.3005
R10080 GND.n3155 GND.n3154 9.3005
R10081 GND.n3156 GND.n3038 9.3005
R10082 GND.n3164 GND.n3163 9.3005
R10083 GND.n3162 GND.n3039 9.3005
R10084 GND.n3161 GND.n3160 9.3005
R10085 GND.n3159 GND.n3157 9.3005
R10086 GND.n3009 GND.n3008 9.3005
R10087 GND.n3195 GND.n3194 9.3005
R10088 GND.n3196 GND.n3006 9.3005
R10089 GND.n3200 GND.n3199 9.3005
R10090 GND.n3198 GND.n3007 9.3005
R10091 GND.n3197 GND.n2981 9.3005
R10092 GND.n3231 GND.n2980 9.3005
R10093 GND.n3233 GND.n3232 9.3005
R10094 GND.n3234 GND.n2979 9.3005
R10095 GND.n3236 GND.n3235 9.3005
R10096 GND.n3242 GND.n2978 9.3005
R10097 GND.n3244 GND.n3243 9.3005
R10098 GND.n3100 GND.n3099 9.3005
R10099 GND.n3033 GND.t44 9.02838
R10100 GND.t0 GND.n2095 9.02838
R10101 GND.n4883 GND.n1457 8.71707
R10102 GND.n4863 GND.n1485 8.71707
R10103 GND.n3816 GND.n1537 8.71707
R10104 GND.n3876 GND.n3875 8.71707
R10105 GND.n3963 GND.n3962 8.71707
R10106 GND.n3929 GND.n1707 8.71707
R10107 GND.n6544 GND.n6543 8.63675
R10108 GND.n3245 GND.n17 8.63675
R10109 GND.n5180 GND.t77 8.40576
R10110 GND.n3239 GND.t6 8.40576
R10111 GND.n3251 GND.t8 8.40576
R10112 GND.n3439 GND.t63 8.40576
R10113 GND.n4280 GND.t102 8.40576
R10114 GND.n4420 GND.t2 8.40576
R10115 GND.n4402 GND.t26 8.40576
R10116 GND.t81 GND.n2063 8.40576
R10117 GND.n4890 GND.n1448 8.09446
R10118 GND.n3837 GND.n2664 8.09446
R10119 GND.n2645 GND.n2644 8.09446
R10120 GND.n3989 GND.n2618 8.09446
R10121 GND.t115 GND.n2712 7.47185
R10122 GND.n4891 GND.n4890 7.47185
R10123 GND.n4856 GND.n4855 7.47185
R10124 GND.n3838 GND.n3837 7.47185
R10125 GND.n3905 GND.n2645 7.47185
R10126 GND.n3955 GND.n2638 7.47185
R10127 GND.n3989 GND.n3980 7.47185
R10128 GND.n5 GND.t32 7.44411
R10129 GND.n5 GND.t52 7.44411
R10130 GND.n7 GND.t24 7.44411
R10131 GND.n7 GND.t10 7.44411
R10132 GND.n10 GND.t9 7.44411
R10133 GND.n10 GND.t38 7.44411
R10134 GND.n12 GND.t141 7.44411
R10135 GND.n12 GND.t48 7.44411
R10136 GND.n0 GND.t59 7.44411
R10137 GND.n0 GND.t29 7.44411
R10138 GND.n2 GND.t143 7.44411
R10139 GND.n2 GND.t7 7.44411
R10140 GND.n29 GND.t27 7.44411
R10141 GND.n29 GND.t18 7.44411
R10142 GND.n27 GND.t16 7.44411
R10143 GND.n27 GND.t49 7.44411
R10144 GND.n34 GND.t138 7.44411
R10145 GND.n34 GND.t22 7.44411
R10146 GND.n32 GND.t142 7.44411
R10147 GND.n32 GND.t13 7.44411
R10148 GND.n40 GND.t31 7.44411
R10149 GND.n40 GND.t41 7.44411
R10150 GND.n38 GND.t19 7.44411
R10151 GND.n38 GND.t3 7.44411
R10152 GND.n2693 GND.n1457 6.84923
R10153 GND.n3754 GND.n1485 6.84923
R10154 GND.n3816 GND.n1543 6.84923
R10155 GND.n3875 GND.n2651 6.84923
R10156 GND.n3962 GND.n2635 6.84923
R10157 GND.n3929 GND.n1701 6.84923
R10158 GND.n4071 GND.n4070 6.5566
R10159 GND.n2758 GND.n2753 6.5566
R10160 GND.n3586 GND.n3585 6.5566
R10161 GND.n4085 GND.n4084 6.5566
R10162 GND.n17 GND.n16 6.29101
R10163 GND.n6544 GND.n43 6.29101
R10164 GND.n3656 GND.n2713 6.22662
R10165 GND.n4897 GND.n1437 6.22662
R10166 GND.n4849 GND.n1504 6.22662
R10167 GND.n3922 GND.n1631 6.22662
R10168 GND.n3998 GND.n2613 6.22662
R10169 GND.n4717 GND.n1748 6.22662
R10170 GND.n6473 GND.n109 6.20656
R10171 GND.n5232 GND.n5231 6.20656
R10172 GND.n3202 GND.t23 5.91532
R10173 GND.n3382 GND.t28 5.91532
R10174 GND.n4342 GND.t15 5.91532
R10175 GND.t17 GND.n4456 5.91532
R10176 GND.n15 GND.n9 5.89418
R10177 GND.n37 GND.n31 5.89418
R10178 GND.n4078 GND.n2353 5.62001
R10179 GND.n2754 GND.n1195 5.62001
R10180 GND.n3581 GND.n1195 5.62001
R10181 GND.n4079 GND.n4078 5.62001
R10182 GND.n4876 GND.n1468 5.60401
R10183 GND.n4870 GND.n1474 5.60401
R10184 GND.n3853 GND.n1560 5.60401
R10185 GND.n3857 GND.n1563 5.60401
R10186 GND.n3941 GND.n1681 5.60401
R10187 GND.n3937 GND.n1684 5.60401
R10188 GND.n3216 GND.t23 5.2927
R10189 GND.n2823 GND.t57 5.2927
R10190 GND.n4689 GND.t36 5.2927
R10191 GND.n4457 GND.t17 5.2927
R10192 GND.n4905 GND.n4904 4.9814
R10193 GND.n3665 GND.n3664 4.9814
R10194 GND.n3810 GND.n3809 4.9814
R10195 GND.n4842 GND.n4841 4.9814
R10196 GND.n3916 GND.n1615 4.9814
R10197 GND.n3918 GND.n1629 4.9814
R10198 GND.n4725 GND.n4724 4.9814
R10199 GND.n4008 GND.n4007 4.9814
R10200 GND.n4427 GND.n4426 4.74817
R10201 GND.n4411 GND.n4377 4.74817
R10202 GND.n4409 GND.n4408 4.74817
R10203 GND.n4391 GND.n4389 4.74817
R10204 GND.n4426 GND.n4425 4.74817
R10205 GND.n4377 GND.n4376 4.74817
R10206 GND.n4410 GND.n4409 4.74817
R10207 GND.n4389 GND.n4378 4.74817
R10208 GND.n3223 GND.n2960 4.74817
R10209 GND.n3276 GND.n3275 4.74817
R10210 GND.n3255 GND.n3254 4.74817
R10211 GND.n3259 GND.n3258 4.74817
R10212 GND.n3256 GND.n2926 4.74817
R10213 GND.n2166 GND.n2140 4.74817
R10214 GND.n4417 GND.n2139 4.74817
R10215 GND.n4394 GND.n2138 4.74817
R10216 GND.n4398 GND.n2137 4.74817
R10217 GND.n2136 GND.n2135 4.74817
R10218 GND.n2144 GND.n2140 4.74817
R10219 GND.n2167 GND.n2139 4.74817
R10220 GND.n4416 GND.n2138 4.74817
R10221 GND.n4395 GND.n2137 4.74817
R10222 GND.n4399 GND.n2136 4.74817
R10223 GND.n3287 GND.n3286 4.74817
R10224 GND.n3270 GND.n2945 4.74817
R10225 GND.n2972 GND.n2944 4.74817
R10226 GND.n3290 GND.n2942 4.74817
R10227 GND.n3287 GND.n2947 4.74817
R10228 GND.n2969 GND.n2945 4.74817
R10229 GND.n3269 GND.n2944 4.74817
R10230 GND.n2971 GND.n2942 4.74817
R10231 GND.n3278 GND.n2960 4.74817
R10232 GND.n3277 GND.n3276 4.74817
R10233 GND.n3254 GND.n2961 4.74817
R10234 GND.n3260 GND.n3259 4.74817
R10235 GND.n3257 GND.n3256 4.74817
R10236 GND.n16 GND.n4 4.70093
R10237 GND.n43 GND.n42 4.70093
R10238 GND.t85 GND.n4960 4.67009
R10239 GND.n4856 GND.t55 4.67009
R10240 GND.n3955 GND.t20 4.67009
R10241 GND.t124 GND.n1845 4.67009
R10242 GND.n15 GND.n14 4.63843
R10243 GND.n37 GND.n36 4.63843
R10244 GND.n2581 GND.n2404 4.6132
R10245 GND.n5075 GND.n1193 4.6132
R10246 GND.t70 GND.n1454 4.35878
R10247 GND.n3744 GND.n1465 4.35878
R10248 GND.n2686 GND.n1477 4.35878
R10249 GND.n2657 GND.n1546 4.35878
R10250 GND.n4808 GND.n4807 4.35878
R10251 GND.n4759 GND.n4758 4.35878
R10252 GND.n3935 GND.n1698 4.35878
R10253 GND.n4738 GND.t95 4.35878
R10254 GND.n4070 GND.n4069 4.05904
R10255 GND.n2761 GND.n2753 4.05904
R10256 GND.n3587 GND.n3586 4.05904
R10257 GND.n4086 GND.n4085 4.05904
R10258 GND.n26 GND.n21 4.04058
R10259 GND.n4911 GND.n1414 3.73617
R10260 GND.n3703 GND.n3675 3.73617
R10261 GND.n3792 GND.n3791 3.73617
R10262 GND.n3800 GND.t25 3.73617
R10263 GND.n4835 GND.n1524 3.73617
R10264 GND.n4794 GND.n4793 3.73617
R10265 GND.t35 GND.n1613 3.73617
R10266 GND.n4773 GND.n4772 3.73617
R10267 GND.n4731 GND.n1727 3.73617
R10268 GND.n4143 GND.n2317 3.73617
R10269 GND.n26 GND.n25 3.53792
R10270 GND.n3771 GND.t55 3.42487
R10271 GND.t20 GND.n3954 3.42487
R10272 GND.n4884 GND.n1454 3.11356
R10273 GND.n4862 GND.n1488 3.11356
R10274 GND.n4828 GND.n4827 3.11356
R10275 GND.n4801 GND.n1588 3.11356
R10276 GND.n4765 GND.n1659 3.11356
R10277 GND.n4739 GND.n4738 3.11356
R10278 GND.t74 GND.n4142 3.11356
R10279 GND.n3105 GND.t77 2.80225
R10280 GND.t8 GND.n2935 2.80225
R10281 GND.n3646 GND.n1401 2.80225
R10282 GND.n4711 GND.t60 2.80225
R10283 GND.n2297 GND.n1757 2.80225
R10284 GND.t2 GND.n2159 2.80225
R10285 GND.n2064 GND.t81 2.80225
R10286 GND.n3561 GND.t67 2.49095
R10287 GND.n3712 GND.n3711 2.49095
R10288 GND.n3770 GND.n2682 2.49095
R10289 GND.n3830 GND.t25 2.49095
R10290 GND.n3820 GND.n1535 2.49095
R10291 GND.n4800 GND.n1590 2.49095
R10292 GND.n3910 GND.t35 2.49095
R10293 GND.n4766 GND.n1657 2.49095
R10294 GND.n2625 GND.n2619 2.49095
R10295 GND.n4426 GND.n2141 2.27742
R10296 GND.n4377 GND.n2141 2.27742
R10297 GND.n4409 GND.n2141 2.27742
R10298 GND.n4389 GND.n2141 2.27742
R10299 GND.n4435 GND.n2140 2.27742
R10300 GND.n4435 GND.n2139 2.27742
R10301 GND.n4435 GND.n2138 2.27742
R10302 GND.n4435 GND.n2137 2.27742
R10303 GND.n4435 GND.n2136 2.27742
R10304 GND.n3288 GND.n3287 2.27742
R10305 GND.n3288 GND.n2945 2.27742
R10306 GND.n3288 GND.n2944 2.27742
R10307 GND.n3288 GND.n2942 2.27742
R10308 GND.n2960 GND.n2925 2.27742
R10309 GND.n3276 GND.n2925 2.27742
R10310 GND.n3254 GND.n2925 2.27742
R10311 GND.n3259 GND.n2925 2.27742
R10312 GND.n3256 GND.n2925 2.27742
R10313 GND.n4912 GND.n1412 1.86834
R10314 GND.n2713 GND.t115 1.86834
R10315 GND.n3702 GND.n1445 1.86834
R10316 GND.n2674 GND.n1496 1.86834
R10317 GND.n4834 GND.n1526 1.86834
R10318 GND.n3906 GND.n1604 1.86834
R10319 GND.n2639 GND.n1640 1.86834
R10320 GND.n4732 GND.n1725 1.86834
R10321 GND.n4142 GND.n4141 1.86834
R10322 GND.n2297 GND.t99 1.86834
R10323 GND.n16 GND.n15 1.59676
R10324 GND.n43 GND.n37 1.59676
R10325 GND.n3820 GND.t42 1.55703
R10326 GND.t136 GND.n1590 1.55703
R10327 GND GND.n17 1.25164
R10328 GND.n3743 GND.n2696 1.24572
R10329 GND.n3757 GND.n2685 1.24572
R10330 GND.n4821 GND.n4820 1.24572
R10331 GND.n2652 GND.n1571 1.24572
R10332 GND.n3945 GND.n1673 1.24572
R10333 GND.n4746 GND.n4745 1.24572
R10334 GND.n5075 GND.n5074 0.970197
R10335 GND.n2581 GND.n2580 0.970197
R10336 GND.n19 GND.n18 0.800888
R10337 GND.n20 GND.n19 0.800888
R10338 GND.n21 GND.n20 0.800888
R10339 GND.n23 GND.n22 0.800888
R10340 GND.n24 GND.n23 0.800888
R10341 GND.n25 GND.n24 0.800888
R10342 GND.n9 GND.n8 0.796477
R10343 GND.n8 GND.n6 0.796477
R10344 GND.n14 GND.n13 0.796477
R10345 GND.n13 GND.n11 0.796477
R10346 GND.n4 GND.n3 0.796477
R10347 GND.n3 GND.n1 0.796477
R10348 GND.n30 GND.n28 0.796477
R10349 GND.n31 GND.n30 0.796477
R10350 GND.n35 GND.n33 0.796477
R10351 GND.n36 GND.n35 0.796477
R10352 GND.n41 GND.n39 0.796477
R10353 GND.n42 GND.n41 0.796477
R10354 GND.n3655 GND.n1425 0.623112
R10355 GND.n4898 GND.n1434 0.623112
R10356 GND.n4848 GND.n1507 0.623112
R10357 GND.n3799 GND.n1516 0.623112
R10358 GND.n4787 GND.n4786 0.623112
R10359 GND.n4780 GND.n4779 0.623112
R10360 GND.n3997 GND.n1736 0.623112
R10361 GND.n4718 GND.n1745 0.623112
R10362 GND.n6545 GND.n6544 0.60351
R10363 GND.n4435 GND.n2141 0.5905
R10364 GND.n3288 GND.n2925 0.5905
R10365 GND.n4192 GND.n4187 0.546232
R10366 GND.n3518 GND.n3517 0.546232
R10367 GND.n2025 GND.n76 0.521841
R10368 GND.n3100 GND.n3098 0.521841
R10369 GND.n6499 GND.n6498 0.494402
R10370 GND.n2370 GND.n1887 0.494402
R10371 GND.n5097 GND.n5096 0.494402
R10372 GND.n1040 GND.n971 0.494402
R10373 GND.n5462 GND.n5461 0.444098
R10374 GND.n6192 GND.n6191 0.444098
R10375 GND.n6344 GND.n6343 0.444098
R10376 GND.n872 GND.n867 0.444098
R10377 GND.n109 GND.n105 0.388379
R10378 GND.n5233 GND.n5232 0.388379
R10379 GND.n6545 GND.n26 0.33279
R10380 GND GND.n6545 0.326523
R10381 GND.n3356 GND.t11 0.311806
R10382 GND.t67 GND.t4 0.311806
R10383 GND.t46 GND.t70 0.311806
R10384 GND.t139 GND.t95 0.311806
R10385 GND.t33 GND.n2213 0.311806
R10386 GND.n4218 GND.n4217 0.306902
R10387 GND.n3468 GND.n3467 0.306902
R10388 GND.n2050 GND.n2049 0.277939
R10389 GND.n5193 GND.n5192 0.277939
R10390 GND.n2541 GND.n2540 0.2505
R10391 GND.n5194 GND.n5193 0.2505
R10392 GND.n2050 GND.n134 0.2505
R10393 GND.n5047 GND.n5045 0.2505
R10394 GND.n1306 GND.n1225 0.239829
R10395 GND.n2443 GND.n1856 0.239829
R10396 GND.n2404 GND.n2403 0.229039
R10397 GND.n2407 GND.n2404 0.229039
R10398 GND.n1193 GND.n1188 0.229039
R10399 GND.n5073 GND.n1193 0.229039
R10400 GND.n1307 GND.n1306 0.152939
R10401 GND.n1308 GND.n1307 0.152939
R10402 GND.n1309 GND.n1308 0.152939
R10403 GND.n1338 GND.n1309 0.152939
R10404 GND.n1339 GND.n1338 0.152939
R10405 GND.n1340 GND.n1339 0.152939
R10406 GND.n1341 GND.n1340 0.152939
R10407 GND.n1342 GND.n1341 0.152939
R10408 GND.n1365 GND.n1342 0.152939
R10409 GND.n1366 GND.n1365 0.152939
R10410 GND.n1367 GND.n1366 0.152939
R10411 GND.n1368 GND.n1367 0.152939
R10412 GND.n1369 GND.n1368 0.152939
R10413 GND.n1392 GND.n1369 0.152939
R10414 GND.n1393 GND.n1392 0.152939
R10415 GND.n1394 GND.n1393 0.152939
R10416 GND.n1395 GND.n1394 0.152939
R10417 GND.n1396 GND.n1395 0.152939
R10418 GND.n1418 GND.n1396 0.152939
R10419 GND.n1419 GND.n1418 0.152939
R10420 GND.n1420 GND.n1419 0.152939
R10421 GND.n1421 GND.n1420 0.152939
R10422 GND.n1422 GND.n1421 0.152939
R10423 GND.n1439 GND.n1422 0.152939
R10424 GND.n1440 GND.n1439 0.152939
R10425 GND.n1441 GND.n1440 0.152939
R10426 GND.n1442 GND.n1441 0.152939
R10427 GND.n1459 GND.n1442 0.152939
R10428 GND.n1460 GND.n1459 0.152939
R10429 GND.n1461 GND.n1460 0.152939
R10430 GND.n1462 GND.n1461 0.152939
R10431 GND.n1479 GND.n1462 0.152939
R10432 GND.n1480 GND.n1479 0.152939
R10433 GND.n1481 GND.n1480 0.152939
R10434 GND.n1482 GND.n1481 0.152939
R10435 GND.n1498 GND.n1482 0.152939
R10436 GND.n1499 GND.n1498 0.152939
R10437 GND.n1500 GND.n1499 0.152939
R10438 GND.n1501 GND.n1500 0.152939
R10439 GND.n1518 GND.n1501 0.152939
R10440 GND.n1519 GND.n1518 0.152939
R10441 GND.n1520 GND.n1519 0.152939
R10442 GND.n1521 GND.n1520 0.152939
R10443 GND.n1550 GND.n1521 0.152939
R10444 GND.n1553 GND.n1550 0.152939
R10445 GND.n1554 GND.n1553 0.152939
R10446 GND.n1555 GND.n1554 0.152939
R10447 GND.n1556 GND.n1555 0.152939
R10448 GND.n1557 GND.n1556 0.152939
R10449 GND.n1594 GND.n1557 0.152939
R10450 GND.n1597 GND.n1594 0.152939
R10451 GND.n1598 GND.n1597 0.152939
R10452 GND.n1599 GND.n1598 0.152939
R10453 GND.n1600 GND.n1599 0.152939
R10454 GND.n1601 GND.n1600 0.152939
R10455 GND.n1644 GND.n1601 0.152939
R10456 GND.n1645 GND.n1644 0.152939
R10457 GND.n1650 GND.n1645 0.152939
R10458 GND.n1651 GND.n1650 0.152939
R10459 GND.n1652 GND.n1651 0.152939
R10460 GND.n1653 GND.n1652 0.152939
R10461 GND.n1654 GND.n1653 0.152939
R10462 GND.n1688 GND.n1654 0.152939
R10463 GND.n1691 GND.n1688 0.152939
R10464 GND.n1692 GND.n1691 0.152939
R10465 GND.n1693 GND.n1692 0.152939
R10466 GND.n1694 GND.n1693 0.152939
R10467 GND.n1695 GND.n1694 0.152939
R10468 GND.n2620 GND.n1695 0.152939
R10469 GND.n2622 GND.n2620 0.152939
R10470 GND.n2622 GND.n2621 0.152939
R10471 GND.n2621 GND.n1731 0.152939
R10472 GND.n1732 GND.n1731 0.152939
R10473 GND.n1733 GND.n1732 0.152939
R10474 GND.n1750 GND.n1733 0.152939
R10475 GND.n1751 GND.n1750 0.152939
R10476 GND.n1752 GND.n1751 0.152939
R10477 GND.n1753 GND.n1752 0.152939
R10478 GND.n1772 GND.n1753 0.152939
R10479 GND.n1773 GND.n1772 0.152939
R10480 GND.n1774 GND.n1773 0.152939
R10481 GND.n1775 GND.n1774 0.152939
R10482 GND.n1776 GND.n1775 0.152939
R10483 GND.n1798 GND.n1776 0.152939
R10484 GND.n1799 GND.n1798 0.152939
R10485 GND.n1800 GND.n1799 0.152939
R10486 GND.n1801 GND.n1800 0.152939
R10487 GND.n1802 GND.n1801 0.152939
R10488 GND.n1825 GND.n1802 0.152939
R10489 GND.n1826 GND.n1825 0.152939
R10490 GND.n1827 GND.n1826 0.152939
R10491 GND.n1828 GND.n1827 0.152939
R10492 GND.n1829 GND.n1828 0.152939
R10493 GND.n1852 GND.n1829 0.152939
R10494 GND.n1853 GND.n1852 0.152939
R10495 GND.n1854 GND.n1853 0.152939
R10496 GND.n1855 GND.n1854 0.152939
R10497 GND.n1856 GND.n1855 0.152939
R10498 GND.n5463 GND.n5462 0.152939
R10499 GND.n5463 GND.n742 0.152939
R10500 GND.n5471 GND.n742 0.152939
R10501 GND.n5472 GND.n5471 0.152939
R10502 GND.n5473 GND.n5472 0.152939
R10503 GND.n5473 GND.n736 0.152939
R10504 GND.n5481 GND.n736 0.152939
R10505 GND.n5482 GND.n5481 0.152939
R10506 GND.n5483 GND.n5482 0.152939
R10507 GND.n5483 GND.n730 0.152939
R10508 GND.n5491 GND.n730 0.152939
R10509 GND.n5492 GND.n5491 0.152939
R10510 GND.n5493 GND.n5492 0.152939
R10511 GND.n5493 GND.n724 0.152939
R10512 GND.n5501 GND.n724 0.152939
R10513 GND.n5502 GND.n5501 0.152939
R10514 GND.n5503 GND.n5502 0.152939
R10515 GND.n5503 GND.n718 0.152939
R10516 GND.n5511 GND.n718 0.152939
R10517 GND.n5512 GND.n5511 0.152939
R10518 GND.n5513 GND.n5512 0.152939
R10519 GND.n5513 GND.n712 0.152939
R10520 GND.n5521 GND.n712 0.152939
R10521 GND.n5522 GND.n5521 0.152939
R10522 GND.n5523 GND.n5522 0.152939
R10523 GND.n5523 GND.n706 0.152939
R10524 GND.n5531 GND.n706 0.152939
R10525 GND.n5532 GND.n5531 0.152939
R10526 GND.n5533 GND.n5532 0.152939
R10527 GND.n5533 GND.n700 0.152939
R10528 GND.n5541 GND.n700 0.152939
R10529 GND.n5542 GND.n5541 0.152939
R10530 GND.n5543 GND.n5542 0.152939
R10531 GND.n5543 GND.n694 0.152939
R10532 GND.n5551 GND.n694 0.152939
R10533 GND.n5552 GND.n5551 0.152939
R10534 GND.n5553 GND.n5552 0.152939
R10535 GND.n5553 GND.n688 0.152939
R10536 GND.n5561 GND.n688 0.152939
R10537 GND.n5562 GND.n5561 0.152939
R10538 GND.n5563 GND.n5562 0.152939
R10539 GND.n5563 GND.n682 0.152939
R10540 GND.n5571 GND.n682 0.152939
R10541 GND.n5572 GND.n5571 0.152939
R10542 GND.n5573 GND.n5572 0.152939
R10543 GND.n5573 GND.n676 0.152939
R10544 GND.n5581 GND.n676 0.152939
R10545 GND.n5582 GND.n5581 0.152939
R10546 GND.n5583 GND.n5582 0.152939
R10547 GND.n5583 GND.n670 0.152939
R10548 GND.n5591 GND.n670 0.152939
R10549 GND.n5592 GND.n5591 0.152939
R10550 GND.n5593 GND.n5592 0.152939
R10551 GND.n5593 GND.n664 0.152939
R10552 GND.n5601 GND.n664 0.152939
R10553 GND.n5602 GND.n5601 0.152939
R10554 GND.n5603 GND.n5602 0.152939
R10555 GND.n5603 GND.n658 0.152939
R10556 GND.n5611 GND.n658 0.152939
R10557 GND.n5612 GND.n5611 0.152939
R10558 GND.n5613 GND.n5612 0.152939
R10559 GND.n5613 GND.n652 0.152939
R10560 GND.n5621 GND.n652 0.152939
R10561 GND.n5622 GND.n5621 0.152939
R10562 GND.n5623 GND.n5622 0.152939
R10563 GND.n5623 GND.n646 0.152939
R10564 GND.n5631 GND.n646 0.152939
R10565 GND.n5632 GND.n5631 0.152939
R10566 GND.n5633 GND.n5632 0.152939
R10567 GND.n5633 GND.n640 0.152939
R10568 GND.n5641 GND.n640 0.152939
R10569 GND.n5642 GND.n5641 0.152939
R10570 GND.n5643 GND.n5642 0.152939
R10571 GND.n5643 GND.n634 0.152939
R10572 GND.n5651 GND.n634 0.152939
R10573 GND.n5652 GND.n5651 0.152939
R10574 GND.n5653 GND.n5652 0.152939
R10575 GND.n5653 GND.n628 0.152939
R10576 GND.n5661 GND.n628 0.152939
R10577 GND.n5662 GND.n5661 0.152939
R10578 GND.n5663 GND.n5662 0.152939
R10579 GND.n5663 GND.n622 0.152939
R10580 GND.n5671 GND.n622 0.152939
R10581 GND.n5672 GND.n5671 0.152939
R10582 GND.n5673 GND.n5672 0.152939
R10583 GND.n5673 GND.n616 0.152939
R10584 GND.n5681 GND.n616 0.152939
R10585 GND.n5682 GND.n5681 0.152939
R10586 GND.n5683 GND.n5682 0.152939
R10587 GND.n5683 GND.n610 0.152939
R10588 GND.n5691 GND.n610 0.152939
R10589 GND.n5692 GND.n5691 0.152939
R10590 GND.n5693 GND.n5692 0.152939
R10591 GND.n5693 GND.n604 0.152939
R10592 GND.n5701 GND.n604 0.152939
R10593 GND.n5702 GND.n5701 0.152939
R10594 GND.n5703 GND.n5702 0.152939
R10595 GND.n5703 GND.n598 0.152939
R10596 GND.n5711 GND.n598 0.152939
R10597 GND.n5712 GND.n5711 0.152939
R10598 GND.n5713 GND.n5712 0.152939
R10599 GND.n5713 GND.n592 0.152939
R10600 GND.n5721 GND.n592 0.152939
R10601 GND.n5722 GND.n5721 0.152939
R10602 GND.n5723 GND.n5722 0.152939
R10603 GND.n5723 GND.n586 0.152939
R10604 GND.n5731 GND.n586 0.152939
R10605 GND.n5732 GND.n5731 0.152939
R10606 GND.n5733 GND.n5732 0.152939
R10607 GND.n5733 GND.n580 0.152939
R10608 GND.n5741 GND.n580 0.152939
R10609 GND.n5742 GND.n5741 0.152939
R10610 GND.n5743 GND.n5742 0.152939
R10611 GND.n5743 GND.n574 0.152939
R10612 GND.n5751 GND.n574 0.152939
R10613 GND.n5752 GND.n5751 0.152939
R10614 GND.n5753 GND.n5752 0.152939
R10615 GND.n5753 GND.n568 0.152939
R10616 GND.n5761 GND.n568 0.152939
R10617 GND.n5762 GND.n5761 0.152939
R10618 GND.n5763 GND.n5762 0.152939
R10619 GND.n5763 GND.n562 0.152939
R10620 GND.n5771 GND.n562 0.152939
R10621 GND.n5772 GND.n5771 0.152939
R10622 GND.n5773 GND.n5772 0.152939
R10623 GND.n5773 GND.n556 0.152939
R10624 GND.n5781 GND.n556 0.152939
R10625 GND.n5782 GND.n5781 0.152939
R10626 GND.n5783 GND.n5782 0.152939
R10627 GND.n5783 GND.n550 0.152939
R10628 GND.n5791 GND.n550 0.152939
R10629 GND.n5792 GND.n5791 0.152939
R10630 GND.n5793 GND.n5792 0.152939
R10631 GND.n5793 GND.n544 0.152939
R10632 GND.n5801 GND.n544 0.152939
R10633 GND.n5802 GND.n5801 0.152939
R10634 GND.n5803 GND.n5802 0.152939
R10635 GND.n5803 GND.n538 0.152939
R10636 GND.n5811 GND.n538 0.152939
R10637 GND.n5812 GND.n5811 0.152939
R10638 GND.n5813 GND.n5812 0.152939
R10639 GND.n5813 GND.n532 0.152939
R10640 GND.n5821 GND.n532 0.152939
R10641 GND.n5822 GND.n5821 0.152939
R10642 GND.n5823 GND.n5822 0.152939
R10643 GND.n5823 GND.n526 0.152939
R10644 GND.n5831 GND.n526 0.152939
R10645 GND.n5832 GND.n5831 0.152939
R10646 GND.n5833 GND.n5832 0.152939
R10647 GND.n5833 GND.n520 0.152939
R10648 GND.n5841 GND.n520 0.152939
R10649 GND.n5842 GND.n5841 0.152939
R10650 GND.n5843 GND.n5842 0.152939
R10651 GND.n5843 GND.n514 0.152939
R10652 GND.n5851 GND.n514 0.152939
R10653 GND.n5852 GND.n5851 0.152939
R10654 GND.n5853 GND.n5852 0.152939
R10655 GND.n5853 GND.n508 0.152939
R10656 GND.n5861 GND.n508 0.152939
R10657 GND.n5862 GND.n5861 0.152939
R10658 GND.n5863 GND.n5862 0.152939
R10659 GND.n5863 GND.n502 0.152939
R10660 GND.n5871 GND.n502 0.152939
R10661 GND.n5872 GND.n5871 0.152939
R10662 GND.n5873 GND.n5872 0.152939
R10663 GND.n5873 GND.n496 0.152939
R10664 GND.n5881 GND.n496 0.152939
R10665 GND.n5882 GND.n5881 0.152939
R10666 GND.n5883 GND.n5882 0.152939
R10667 GND.n5883 GND.n490 0.152939
R10668 GND.n5891 GND.n490 0.152939
R10669 GND.n5892 GND.n5891 0.152939
R10670 GND.n5893 GND.n5892 0.152939
R10671 GND.n5893 GND.n484 0.152939
R10672 GND.n5901 GND.n484 0.152939
R10673 GND.n5902 GND.n5901 0.152939
R10674 GND.n5903 GND.n5902 0.152939
R10675 GND.n5903 GND.n478 0.152939
R10676 GND.n5911 GND.n478 0.152939
R10677 GND.n5912 GND.n5911 0.152939
R10678 GND.n5913 GND.n5912 0.152939
R10679 GND.n5913 GND.n472 0.152939
R10680 GND.n5921 GND.n472 0.152939
R10681 GND.n5922 GND.n5921 0.152939
R10682 GND.n5923 GND.n5922 0.152939
R10683 GND.n5923 GND.n466 0.152939
R10684 GND.n5931 GND.n466 0.152939
R10685 GND.n5932 GND.n5931 0.152939
R10686 GND.n5933 GND.n5932 0.152939
R10687 GND.n5933 GND.n460 0.152939
R10688 GND.n5941 GND.n460 0.152939
R10689 GND.n5942 GND.n5941 0.152939
R10690 GND.n5943 GND.n5942 0.152939
R10691 GND.n5943 GND.n454 0.152939
R10692 GND.n5951 GND.n454 0.152939
R10693 GND.n5952 GND.n5951 0.152939
R10694 GND.n5953 GND.n5952 0.152939
R10695 GND.n5953 GND.n448 0.152939
R10696 GND.n5961 GND.n448 0.152939
R10697 GND.n5962 GND.n5961 0.152939
R10698 GND.n5963 GND.n5962 0.152939
R10699 GND.n5963 GND.n442 0.152939
R10700 GND.n5971 GND.n442 0.152939
R10701 GND.n5972 GND.n5971 0.152939
R10702 GND.n5973 GND.n5972 0.152939
R10703 GND.n5973 GND.n436 0.152939
R10704 GND.n5981 GND.n436 0.152939
R10705 GND.n5982 GND.n5981 0.152939
R10706 GND.n5983 GND.n5982 0.152939
R10707 GND.n5983 GND.n430 0.152939
R10708 GND.n5991 GND.n430 0.152939
R10709 GND.n5992 GND.n5991 0.152939
R10710 GND.n5993 GND.n5992 0.152939
R10711 GND.n5993 GND.n424 0.152939
R10712 GND.n6001 GND.n424 0.152939
R10713 GND.n6002 GND.n6001 0.152939
R10714 GND.n6003 GND.n6002 0.152939
R10715 GND.n6003 GND.n418 0.152939
R10716 GND.n6011 GND.n418 0.152939
R10717 GND.n6012 GND.n6011 0.152939
R10718 GND.n6013 GND.n6012 0.152939
R10719 GND.n6013 GND.n412 0.152939
R10720 GND.n6021 GND.n412 0.152939
R10721 GND.n6022 GND.n6021 0.152939
R10722 GND.n6023 GND.n6022 0.152939
R10723 GND.n6023 GND.n406 0.152939
R10724 GND.n6031 GND.n406 0.152939
R10725 GND.n6032 GND.n6031 0.152939
R10726 GND.n6033 GND.n6032 0.152939
R10727 GND.n6033 GND.n400 0.152939
R10728 GND.n6041 GND.n400 0.152939
R10729 GND.n6042 GND.n6041 0.152939
R10730 GND.n6043 GND.n6042 0.152939
R10731 GND.n6043 GND.n394 0.152939
R10732 GND.n6051 GND.n394 0.152939
R10733 GND.n6052 GND.n6051 0.152939
R10734 GND.n6053 GND.n6052 0.152939
R10735 GND.n6053 GND.n388 0.152939
R10736 GND.n6061 GND.n388 0.152939
R10737 GND.n6062 GND.n6061 0.152939
R10738 GND.n6063 GND.n6062 0.152939
R10739 GND.n6063 GND.n382 0.152939
R10740 GND.n6071 GND.n382 0.152939
R10741 GND.n6072 GND.n6071 0.152939
R10742 GND.n6073 GND.n6072 0.152939
R10743 GND.n6073 GND.n376 0.152939
R10744 GND.n6081 GND.n376 0.152939
R10745 GND.n6082 GND.n6081 0.152939
R10746 GND.n6083 GND.n6082 0.152939
R10747 GND.n6083 GND.n370 0.152939
R10748 GND.n6091 GND.n370 0.152939
R10749 GND.n6092 GND.n6091 0.152939
R10750 GND.n6093 GND.n6092 0.152939
R10751 GND.n6093 GND.n364 0.152939
R10752 GND.n6101 GND.n364 0.152939
R10753 GND.n6102 GND.n6101 0.152939
R10754 GND.n6103 GND.n6102 0.152939
R10755 GND.n6103 GND.n358 0.152939
R10756 GND.n6111 GND.n358 0.152939
R10757 GND.n6112 GND.n6111 0.152939
R10758 GND.n6113 GND.n6112 0.152939
R10759 GND.n6113 GND.n352 0.152939
R10760 GND.n6121 GND.n352 0.152939
R10761 GND.n6122 GND.n6121 0.152939
R10762 GND.n6123 GND.n6122 0.152939
R10763 GND.n6123 GND.n346 0.152939
R10764 GND.n6131 GND.n346 0.152939
R10765 GND.n6132 GND.n6131 0.152939
R10766 GND.n6133 GND.n6132 0.152939
R10767 GND.n6133 GND.n340 0.152939
R10768 GND.n6141 GND.n340 0.152939
R10769 GND.n6142 GND.n6141 0.152939
R10770 GND.n6143 GND.n6142 0.152939
R10771 GND.n6143 GND.n334 0.152939
R10772 GND.n6151 GND.n334 0.152939
R10773 GND.n6152 GND.n6151 0.152939
R10774 GND.n6153 GND.n6152 0.152939
R10775 GND.n6153 GND.n328 0.152939
R10776 GND.n6161 GND.n328 0.152939
R10777 GND.n6162 GND.n6161 0.152939
R10778 GND.n6163 GND.n6162 0.152939
R10779 GND.n6163 GND.n322 0.152939
R10780 GND.n6171 GND.n322 0.152939
R10781 GND.n6172 GND.n6171 0.152939
R10782 GND.n6173 GND.n6172 0.152939
R10783 GND.n6173 GND.n316 0.152939
R10784 GND.n6181 GND.n316 0.152939
R10785 GND.n6182 GND.n6181 0.152939
R10786 GND.n6183 GND.n6182 0.152939
R10787 GND.n6183 GND.n310 0.152939
R10788 GND.n6191 GND.n310 0.152939
R10789 GND.n6193 GND.n6192 0.152939
R10790 GND.n6193 GND.n304 0.152939
R10791 GND.n6201 GND.n304 0.152939
R10792 GND.n6202 GND.n6201 0.152939
R10793 GND.n6203 GND.n6202 0.152939
R10794 GND.n6203 GND.n298 0.152939
R10795 GND.n6211 GND.n298 0.152939
R10796 GND.n6212 GND.n6211 0.152939
R10797 GND.n6213 GND.n6212 0.152939
R10798 GND.n6213 GND.n292 0.152939
R10799 GND.n6221 GND.n292 0.152939
R10800 GND.n6222 GND.n6221 0.152939
R10801 GND.n6223 GND.n6222 0.152939
R10802 GND.n6223 GND.n286 0.152939
R10803 GND.n6231 GND.n286 0.152939
R10804 GND.n6232 GND.n6231 0.152939
R10805 GND.n6233 GND.n6232 0.152939
R10806 GND.n6233 GND.n280 0.152939
R10807 GND.n6241 GND.n280 0.152939
R10808 GND.n6242 GND.n6241 0.152939
R10809 GND.n6243 GND.n6242 0.152939
R10810 GND.n6243 GND.n274 0.152939
R10811 GND.n6251 GND.n274 0.152939
R10812 GND.n6252 GND.n6251 0.152939
R10813 GND.n6253 GND.n6252 0.152939
R10814 GND.n6253 GND.n268 0.152939
R10815 GND.n6261 GND.n268 0.152939
R10816 GND.n6262 GND.n6261 0.152939
R10817 GND.n6263 GND.n6262 0.152939
R10818 GND.n6263 GND.n262 0.152939
R10819 GND.n6271 GND.n262 0.152939
R10820 GND.n6272 GND.n6271 0.152939
R10821 GND.n6273 GND.n6272 0.152939
R10822 GND.n6273 GND.n256 0.152939
R10823 GND.n6281 GND.n256 0.152939
R10824 GND.n6282 GND.n6281 0.152939
R10825 GND.n6283 GND.n6282 0.152939
R10826 GND.n6283 GND.n250 0.152939
R10827 GND.n6291 GND.n250 0.152939
R10828 GND.n6292 GND.n6291 0.152939
R10829 GND.n6293 GND.n6292 0.152939
R10830 GND.n6293 GND.n244 0.152939
R10831 GND.n6301 GND.n244 0.152939
R10832 GND.n6302 GND.n6301 0.152939
R10833 GND.n6303 GND.n6302 0.152939
R10834 GND.n6303 GND.n238 0.152939
R10835 GND.n6311 GND.n238 0.152939
R10836 GND.n6312 GND.n6311 0.152939
R10837 GND.n6313 GND.n6312 0.152939
R10838 GND.n6313 GND.n232 0.152939
R10839 GND.n6321 GND.n232 0.152939
R10840 GND.n6322 GND.n6321 0.152939
R10841 GND.n6323 GND.n6322 0.152939
R10842 GND.n6323 GND.n226 0.152939
R10843 GND.n6331 GND.n226 0.152939
R10844 GND.n6332 GND.n6331 0.152939
R10845 GND.n6334 GND.n6332 0.152939
R10846 GND.n6334 GND.n6333 0.152939
R10847 GND.n6333 GND.n220 0.152939
R10848 GND.n6343 GND.n220 0.152939
R10849 GND.n4437 GND.n4436 0.152939
R10850 GND.n4437 GND.n2114 0.152939
R10851 GND.n4460 GND.n2114 0.152939
R10852 GND.n4461 GND.n4460 0.152939
R10853 GND.n4462 GND.n4461 0.152939
R10854 GND.n4463 GND.n4462 0.152939
R10855 GND.n4463 GND.n2091 0.152939
R10856 GND.n4486 GND.n2091 0.152939
R10857 GND.n4487 GND.n4486 0.152939
R10858 GND.n4488 GND.n4487 0.152939
R10859 GND.n4489 GND.n4488 0.152939
R10860 GND.n4489 GND.n2072 0.152939
R10861 GND.n4515 GND.n2072 0.152939
R10862 GND.n4516 GND.n4515 0.152939
R10863 GND.n4517 GND.n4516 0.152939
R10864 GND.n4518 GND.n4517 0.152939
R10865 GND.n4519 GND.n4518 0.152939
R10866 GND.n4522 GND.n4519 0.152939
R10867 GND.n4523 GND.n4522 0.152939
R10868 GND.n4524 GND.n4523 0.152939
R10869 GND.n4526 GND.n4524 0.152939
R10870 GND.n4526 GND.n4525 0.152939
R10871 GND.n4525 GND.n148 0.152939
R10872 GND.n149 GND.n148 0.152939
R10873 GND.n150 GND.n149 0.152939
R10874 GND.n155 GND.n150 0.152939
R10875 GND.n156 GND.n155 0.152939
R10876 GND.n157 GND.n156 0.152939
R10877 GND.n158 GND.n157 0.152939
R10878 GND.n163 GND.n158 0.152939
R10879 GND.n164 GND.n163 0.152939
R10880 GND.n165 GND.n164 0.152939
R10881 GND.n166 GND.n165 0.152939
R10882 GND.n171 GND.n166 0.152939
R10883 GND.n172 GND.n171 0.152939
R10884 GND.n173 GND.n172 0.152939
R10885 GND.n174 GND.n173 0.152939
R10886 GND.n179 GND.n174 0.152939
R10887 GND.n180 GND.n179 0.152939
R10888 GND.n181 GND.n180 0.152939
R10889 GND.n182 GND.n181 0.152939
R10890 GND.n187 GND.n182 0.152939
R10891 GND.n188 GND.n187 0.152939
R10892 GND.n189 GND.n188 0.152939
R10893 GND.n190 GND.n189 0.152939
R10894 GND.n195 GND.n190 0.152939
R10895 GND.n196 GND.n195 0.152939
R10896 GND.n197 GND.n196 0.152939
R10897 GND.n198 GND.n197 0.152939
R10898 GND.n203 GND.n198 0.152939
R10899 GND.n204 GND.n203 0.152939
R10900 GND.n205 GND.n204 0.152939
R10901 GND.n206 GND.n205 0.152939
R10902 GND.n211 GND.n206 0.152939
R10903 GND.n212 GND.n211 0.152939
R10904 GND.n213 GND.n212 0.152939
R10905 GND.n214 GND.n213 0.152939
R10906 GND.n219 GND.n214 0.152939
R10907 GND.n6344 GND.n219 0.152939
R10908 GND.n4449 GND.n2125 0.152939
R10909 GND.n4450 GND.n4449 0.152939
R10910 GND.n4451 GND.n4450 0.152939
R10911 GND.n4452 GND.n4451 0.152939
R10912 GND.n4452 GND.n2101 0.152939
R10913 GND.n4475 GND.n2101 0.152939
R10914 GND.n4476 GND.n4475 0.152939
R10915 GND.n4477 GND.n4476 0.152939
R10916 GND.n4478 GND.n4477 0.152939
R10917 GND.n4478 GND.n2081 0.152939
R10918 GND.n4504 GND.n2081 0.152939
R10919 GND.n4505 GND.n4504 0.152939
R10920 GND.n4506 GND.n4505 0.152939
R10921 GND.n4507 GND.n4506 0.152939
R10922 GND.n4507 GND.n2059 0.152939
R10923 GND.n4546 GND.n2059 0.152939
R10924 GND.n4547 GND.n4546 0.152939
R10925 GND.n4548 GND.n4547 0.152939
R10926 GND.n4548 GND.n86 0.152939
R10927 GND.n6499 GND.n86 0.152939
R10928 GND.n2371 GND.n2370 0.152939
R10929 GND.n2372 GND.n2371 0.152939
R10930 GND.n2372 GND.n2364 0.152939
R10931 GND.n2380 GND.n2364 0.152939
R10932 GND.n2381 GND.n2380 0.152939
R10933 GND.n2382 GND.n2381 0.152939
R10934 GND.n2382 GND.n2360 0.152939
R10935 GND.n2390 GND.n2360 0.152939
R10936 GND.n2391 GND.n2390 0.152939
R10937 GND.n2392 GND.n2391 0.152939
R10938 GND.n2392 GND.n2356 0.152939
R10939 GND.n2402 GND.n2356 0.152939
R10940 GND.n2403 GND.n2402 0.152939
R10941 GND.n2410 GND.n2407 0.152939
R10942 GND.n2411 GND.n2410 0.152939
R10943 GND.n2412 GND.n2411 0.152939
R10944 GND.n2413 GND.n2412 0.152939
R10945 GND.n2416 GND.n2413 0.152939
R10946 GND.n2417 GND.n2416 0.152939
R10947 GND.n2418 GND.n2417 0.152939
R10948 GND.n2419 GND.n2418 0.152939
R10949 GND.n2422 GND.n2419 0.152939
R10950 GND.n2423 GND.n2422 0.152939
R10951 GND.n2424 GND.n2423 0.152939
R10952 GND.n2425 GND.n2424 0.152939
R10953 GND.n2428 GND.n2425 0.152939
R10954 GND.n2429 GND.n2428 0.152939
R10955 GND.n2430 GND.n2429 0.152939
R10956 GND.n2431 GND.n2430 0.152939
R10957 GND.n2435 GND.n2431 0.152939
R10958 GND.n2541 GND.n2435 0.152939
R10959 GND.n1888 GND.n1887 0.152939
R10960 GND.n1889 GND.n1888 0.152939
R10961 GND.n4222 GND.n1889 0.152939
R10962 GND.n4223 GND.n4222 0.152939
R10963 GND.n4223 GND.n2230 0.152939
R10964 GND.n4298 GND.n2230 0.152939
R10965 GND.n4299 GND.n4298 0.152939
R10966 GND.n4300 GND.n4299 0.152939
R10967 GND.n4301 GND.n4300 0.152939
R10968 GND.n4301 GND.n2208 0.152939
R10969 GND.n4323 GND.n2208 0.152939
R10970 GND.n4324 GND.n4323 0.152939
R10971 GND.n4325 GND.n4324 0.152939
R10972 GND.n4326 GND.n4325 0.152939
R10973 GND.n4326 GND.n2185 0.152939
R10974 GND.n4348 GND.n2185 0.152939
R10975 GND.n4349 GND.n4348 0.152939
R10976 GND.n4351 GND.n4349 0.152939
R10977 GND.n4351 GND.n4350 0.152939
R10978 GND.n4350 GND.n2154 0.152939
R10979 GND.n3307 GND.n3306 0.152939
R10980 GND.n3308 GND.n3307 0.152939
R10981 GND.n3309 GND.n3308 0.152939
R10982 GND.n3310 GND.n3309 0.152939
R10983 GND.n3313 GND.n3310 0.152939
R10984 GND.n3314 GND.n3313 0.152939
R10985 GND.n3315 GND.n3314 0.152939
R10986 GND.n3316 GND.n3315 0.152939
R10987 GND.n3319 GND.n3316 0.152939
R10988 GND.n3320 GND.n3319 0.152939
R10989 GND.n3321 GND.n3320 0.152939
R10990 GND.n3322 GND.n3321 0.152939
R10991 GND.n3325 GND.n3322 0.152939
R10992 GND.n3326 GND.n3325 0.152939
R10993 GND.n3327 GND.n3326 0.152939
R10994 GND.n3328 GND.n3327 0.152939
R10995 GND.n3331 GND.n3328 0.152939
R10996 GND.n3332 GND.n3331 0.152939
R10997 GND.n3333 GND.n3332 0.152939
R10998 GND.n3335 GND.n3333 0.152939
R10999 GND.n3335 GND.n3334 0.152939
R11000 GND.n3334 GND.n1295 0.152939
R11001 GND.n1296 GND.n1295 0.152939
R11002 GND.n1297 GND.n1296 0.152939
R11003 GND.n1318 GND.n1297 0.152939
R11004 GND.n1319 GND.n1318 0.152939
R11005 GND.n1320 GND.n1319 0.152939
R11006 GND.n1324 GND.n1320 0.152939
R11007 GND.n1325 GND.n1324 0.152939
R11008 GND.n1326 GND.n1325 0.152939
R11009 GND.n1327 GND.n1326 0.152939
R11010 GND.n1328 GND.n1327 0.152939
R11011 GND.n1351 GND.n1328 0.152939
R11012 GND.n1352 GND.n1351 0.152939
R11013 GND.n1353 GND.n1352 0.152939
R11014 GND.n1354 GND.n1353 0.152939
R11015 GND.n1355 GND.n1354 0.152939
R11016 GND.n1378 GND.n1355 0.152939
R11017 GND.n1379 GND.n1378 0.152939
R11018 GND.n1380 GND.n1379 0.152939
R11019 GND.n1381 GND.n1380 0.152939
R11020 GND.n1382 GND.n1381 0.152939
R11021 GND.n1405 GND.n1382 0.152939
R11022 GND.n1406 GND.n1405 0.152939
R11023 GND.n1407 GND.n1406 0.152939
R11024 GND.n1408 GND.n1407 0.152939
R11025 GND.n1409 GND.n1408 0.152939
R11026 GND.n3682 GND.n1409 0.152939
R11027 GND.n3683 GND.n3682 0.152939
R11028 GND.n3683 GND.n3680 0.152939
R11029 GND.n3689 GND.n3680 0.152939
R11030 GND.n3690 GND.n3689 0.152939
R11031 GND.n3691 GND.n3690 0.152939
R11032 GND.n3692 GND.n3691 0.152939
R11033 GND.n3693 GND.n3692 0.152939
R11034 GND.n3695 GND.n3693 0.152939
R11035 GND.n3695 GND.n3694 0.152939
R11036 GND.n3694 GND.n2689 0.152939
R11037 GND.n3749 GND.n2689 0.152939
R11038 GND.n3750 GND.n3749 0.152939
R11039 GND.n3751 GND.n3750 0.152939
R11040 GND.n3751 GND.n2679 0.152939
R11041 GND.n3774 GND.n2679 0.152939
R11042 GND.n3775 GND.n3774 0.152939
R11043 GND.n3776 GND.n3775 0.152939
R11044 GND.n3777 GND.n3776 0.152939
R11045 GND.n3778 GND.n3777 0.152939
R11046 GND.n3780 GND.n3778 0.152939
R11047 GND.n3780 GND.n3779 0.152939
R11048 GND.n3779 GND.n1530 0.152939
R11049 GND.n1531 GND.n1530 0.152939
R11050 GND.n1532 GND.n1531 0.152939
R11051 GND.n1575 GND.n1532 0.152939
R11052 GND.n1576 GND.n1575 0.152939
R11053 GND.n1581 GND.n1576 0.152939
R11054 GND.n1582 GND.n1581 0.152939
R11055 GND.n1583 GND.n1582 0.152939
R11056 GND.n1584 GND.n1583 0.152939
R11057 GND.n1585 GND.n1584 0.152939
R11058 GND.n1619 GND.n1585 0.152939
R11059 GND.n1622 GND.n1619 0.152939
R11060 GND.n1623 GND.n1622 0.152939
R11061 GND.n1624 GND.n1623 0.152939
R11062 GND.n1625 GND.n1624 0.152939
R11063 GND.n1626 GND.n1625 0.152939
R11064 GND.n1663 GND.n1626 0.152939
R11065 GND.n1666 GND.n1663 0.152939
R11066 GND.n1667 GND.n1666 0.152939
R11067 GND.n1668 GND.n1667 0.152939
R11068 GND.n1669 GND.n1668 0.152939
R11069 GND.n1670 GND.n1669 0.152939
R11070 GND.n1712 GND.n1670 0.152939
R11071 GND.n1713 GND.n1712 0.152939
R11072 GND.n1718 GND.n1713 0.152939
R11073 GND.n1719 GND.n1718 0.152939
R11074 GND.n1720 GND.n1719 0.152939
R11075 GND.n1721 GND.n1720 0.152939
R11076 GND.n1722 GND.n1721 0.152939
R11077 GND.n2304 GND.n1722 0.152939
R11078 GND.n2305 GND.n2304 0.152939
R11079 GND.n2310 GND.n2305 0.152939
R11080 GND.n2311 GND.n2310 0.152939
R11081 GND.n2313 GND.n2311 0.152939
R11082 GND.n2313 GND.n2312 0.152939
R11083 GND.n2312 GND.n1761 0.152939
R11084 GND.n1762 GND.n1761 0.152939
R11085 GND.n1763 GND.n1762 0.152939
R11086 GND.n1785 GND.n1763 0.152939
R11087 GND.n1786 GND.n1785 0.152939
R11088 GND.n1787 GND.n1786 0.152939
R11089 GND.n1788 GND.n1787 0.152939
R11090 GND.n1789 GND.n1788 0.152939
R11091 GND.n1811 GND.n1789 0.152939
R11092 GND.n1812 GND.n1811 0.152939
R11093 GND.n1813 GND.n1812 0.152939
R11094 GND.n1814 GND.n1813 0.152939
R11095 GND.n1815 GND.n1814 0.152939
R11096 GND.n1838 GND.n1815 0.152939
R11097 GND.n1839 GND.n1838 0.152939
R11098 GND.n1840 GND.n1839 0.152939
R11099 GND.n1841 GND.n1840 0.152939
R11100 GND.n1842 GND.n1841 0.152939
R11101 GND.n1864 GND.n1842 0.152939
R11102 GND.n1865 GND.n1864 0.152939
R11103 GND.n1866 GND.n1865 0.152939
R11104 GND.n1867 GND.n1866 0.152939
R11105 GND.n1868 GND.n1867 0.152939
R11106 GND.n1874 GND.n1868 0.152939
R11107 GND.n1875 GND.n1874 0.152939
R11108 GND.n1876 GND.n1875 0.152939
R11109 GND.n1877 GND.n1876 0.152939
R11110 GND.n4230 GND.n1877 0.152939
R11111 GND.n4233 GND.n4230 0.152939
R11112 GND.n4234 GND.n4233 0.152939
R11113 GND.n4235 GND.n4234 0.152939
R11114 GND.n4236 GND.n4235 0.152939
R11115 GND.n4237 GND.n4236 0.152939
R11116 GND.n4240 GND.n4237 0.152939
R11117 GND.n4241 GND.n4240 0.152939
R11118 GND.n4242 GND.n4241 0.152939
R11119 GND.n4243 GND.n4242 0.152939
R11120 GND.n4246 GND.n4243 0.152939
R11121 GND.n4247 GND.n4246 0.152939
R11122 GND.n4248 GND.n4247 0.152939
R11123 GND.n4249 GND.n4248 0.152939
R11124 GND.n4252 GND.n4249 0.152939
R11125 GND.n4253 GND.n4252 0.152939
R11126 GND.n4254 GND.n4253 0.152939
R11127 GND.n4255 GND.n4254 0.152939
R11128 GND.n4255 GND.n2142 0.152939
R11129 GND.n4434 GND.n2142 0.152939
R11130 GND.n3375 GND.n2914 0.152939
R11131 GND.n3376 GND.n3375 0.152939
R11132 GND.n3377 GND.n3376 0.152939
R11133 GND.n3378 GND.n3377 0.152939
R11134 GND.n3378 GND.n2892 0.152939
R11135 GND.n3400 GND.n2892 0.152939
R11136 GND.n3401 GND.n3400 0.152939
R11137 GND.n3402 GND.n3401 0.152939
R11138 GND.n3403 GND.n3402 0.152939
R11139 GND.n3403 GND.n2873 0.152939
R11140 GND.n3425 GND.n2873 0.152939
R11141 GND.n3426 GND.n3425 0.152939
R11142 GND.n3427 GND.n3426 0.152939
R11143 GND.n3428 GND.n3427 0.152939
R11144 GND.n3428 GND.n2850 0.152939
R11145 GND.n3453 GND.n2850 0.152939
R11146 GND.n3454 GND.n3453 0.152939
R11147 GND.n3455 GND.n3454 0.152939
R11148 GND.n3455 GND.n1173 0.152939
R11149 GND.n5097 GND.n1173 0.152939
R11150 GND.n972 GND.n971 0.152939
R11151 GND.n973 GND.n972 0.152939
R11152 GND.n974 GND.n973 0.152939
R11153 GND.n975 GND.n974 0.152939
R11154 GND.n976 GND.n975 0.152939
R11155 GND.n977 GND.n976 0.152939
R11156 GND.n978 GND.n977 0.152939
R11157 GND.n979 GND.n978 0.152939
R11158 GND.n980 GND.n979 0.152939
R11159 GND.n981 GND.n980 0.152939
R11160 GND.n982 GND.n981 0.152939
R11161 GND.n983 GND.n982 0.152939
R11162 GND.n984 GND.n983 0.152939
R11163 GND.n985 GND.n984 0.152939
R11164 GND.n986 GND.n985 0.152939
R11165 GND.n989 GND.n986 0.152939
R11166 GND.n990 GND.n989 0.152939
R11167 GND.n991 GND.n990 0.152939
R11168 GND.n992 GND.n991 0.152939
R11169 GND.n993 GND.n992 0.152939
R11170 GND.n994 GND.n993 0.152939
R11171 GND.n995 GND.n994 0.152939
R11172 GND.n996 GND.n995 0.152939
R11173 GND.n997 GND.n996 0.152939
R11174 GND.n998 GND.n997 0.152939
R11175 GND.n999 GND.n998 0.152939
R11176 GND.n1000 GND.n999 0.152939
R11177 GND.n1001 GND.n1000 0.152939
R11178 GND.n1002 GND.n1001 0.152939
R11179 GND.n1003 GND.n1002 0.152939
R11180 GND.n1004 GND.n1003 0.152939
R11181 GND.n1005 GND.n1004 0.152939
R11182 GND.n5195 GND.n1005 0.152939
R11183 GND.n5195 GND.n5194 0.152939
R11184 GND.n1044 GND.n1040 0.152939
R11185 GND.n1045 GND.n1044 0.152939
R11186 GND.n1046 GND.n1045 0.152939
R11187 GND.n1047 GND.n1046 0.152939
R11188 GND.n1048 GND.n1047 0.152939
R11189 GND.n3145 GND.n1048 0.152939
R11190 GND.n3146 GND.n3145 0.152939
R11191 GND.n3147 GND.n3146 0.152939
R11192 GND.n3148 GND.n3147 0.152939
R11193 GND.n3148 GND.n3028 0.152939
R11194 GND.n3173 GND.n3028 0.152939
R11195 GND.n3174 GND.n3173 0.152939
R11196 GND.n3175 GND.n3174 0.152939
R11197 GND.n3176 GND.n3175 0.152939
R11198 GND.n3176 GND.n2998 0.152939
R11199 GND.n3208 GND.n2998 0.152939
R11200 GND.n3209 GND.n3208 0.152939
R11201 GND.n3210 GND.n3209 0.152939
R11202 GND.n3211 GND.n3210 0.152939
R11203 GND.n3211 GND.n2943 0.152939
R11204 GND.n873 GND.n872 0.152939
R11205 GND.n874 GND.n873 0.152939
R11206 GND.n875 GND.n874 0.152939
R11207 GND.n880 GND.n875 0.152939
R11208 GND.n881 GND.n880 0.152939
R11209 GND.n882 GND.n881 0.152939
R11210 GND.n883 GND.n882 0.152939
R11211 GND.n888 GND.n883 0.152939
R11212 GND.n889 GND.n888 0.152939
R11213 GND.n890 GND.n889 0.152939
R11214 GND.n891 GND.n890 0.152939
R11215 GND.n896 GND.n891 0.152939
R11216 GND.n897 GND.n896 0.152939
R11217 GND.n898 GND.n897 0.152939
R11218 GND.n899 GND.n898 0.152939
R11219 GND.n904 GND.n899 0.152939
R11220 GND.n905 GND.n904 0.152939
R11221 GND.n906 GND.n905 0.152939
R11222 GND.n907 GND.n906 0.152939
R11223 GND.n912 GND.n907 0.152939
R11224 GND.n913 GND.n912 0.152939
R11225 GND.n914 GND.n913 0.152939
R11226 GND.n915 GND.n914 0.152939
R11227 GND.n920 GND.n915 0.152939
R11228 GND.n921 GND.n920 0.152939
R11229 GND.n922 GND.n921 0.152939
R11230 GND.n923 GND.n922 0.152939
R11231 GND.n928 GND.n923 0.152939
R11232 GND.n929 GND.n928 0.152939
R11233 GND.n930 GND.n929 0.152939
R11234 GND.n931 GND.n930 0.152939
R11235 GND.n936 GND.n931 0.152939
R11236 GND.n937 GND.n936 0.152939
R11237 GND.n938 GND.n937 0.152939
R11238 GND.n939 GND.n938 0.152939
R11239 GND.n1022 GND.n939 0.152939
R11240 GND.n1025 GND.n1022 0.152939
R11241 GND.n1026 GND.n1025 0.152939
R11242 GND.n1027 GND.n1026 0.152939
R11243 GND.n1028 GND.n1027 0.152939
R11244 GND.n1029 GND.n1028 0.152939
R11245 GND.n3119 GND.n1029 0.152939
R11246 GND.n3122 GND.n3119 0.152939
R11247 GND.n3123 GND.n3122 0.152939
R11248 GND.n3124 GND.n3123 0.152939
R11249 GND.n3125 GND.n3124 0.152939
R11250 GND.n3126 GND.n3125 0.152939
R11251 GND.n3128 GND.n3126 0.152939
R11252 GND.n3129 GND.n3128 0.152939
R11253 GND.n3129 GND.n3015 0.152939
R11254 GND.n3184 GND.n3015 0.152939
R11255 GND.n3185 GND.n3184 0.152939
R11256 GND.n3186 GND.n3185 0.152939
R11257 GND.n3187 GND.n3186 0.152939
R11258 GND.n3187 GND.n2987 0.152939
R11259 GND.n3219 GND.n2987 0.152939
R11260 GND.n3220 GND.n3219 0.152939
R11261 GND.n3221 GND.n3220 0.152939
R11262 GND.n3222 GND.n3221 0.152939
R11263 GND.n5461 GND.n748 0.152939
R11264 GND.n753 GND.n748 0.152939
R11265 GND.n754 GND.n753 0.152939
R11266 GND.n755 GND.n754 0.152939
R11267 GND.n760 GND.n755 0.152939
R11268 GND.n761 GND.n760 0.152939
R11269 GND.n762 GND.n761 0.152939
R11270 GND.n763 GND.n762 0.152939
R11271 GND.n768 GND.n763 0.152939
R11272 GND.n769 GND.n768 0.152939
R11273 GND.n770 GND.n769 0.152939
R11274 GND.n771 GND.n770 0.152939
R11275 GND.n776 GND.n771 0.152939
R11276 GND.n777 GND.n776 0.152939
R11277 GND.n778 GND.n777 0.152939
R11278 GND.n779 GND.n778 0.152939
R11279 GND.n784 GND.n779 0.152939
R11280 GND.n785 GND.n784 0.152939
R11281 GND.n786 GND.n785 0.152939
R11282 GND.n787 GND.n786 0.152939
R11283 GND.n792 GND.n787 0.152939
R11284 GND.n793 GND.n792 0.152939
R11285 GND.n794 GND.n793 0.152939
R11286 GND.n795 GND.n794 0.152939
R11287 GND.n800 GND.n795 0.152939
R11288 GND.n801 GND.n800 0.152939
R11289 GND.n802 GND.n801 0.152939
R11290 GND.n803 GND.n802 0.152939
R11291 GND.n808 GND.n803 0.152939
R11292 GND.n809 GND.n808 0.152939
R11293 GND.n810 GND.n809 0.152939
R11294 GND.n811 GND.n810 0.152939
R11295 GND.n816 GND.n811 0.152939
R11296 GND.n817 GND.n816 0.152939
R11297 GND.n818 GND.n817 0.152939
R11298 GND.n819 GND.n818 0.152939
R11299 GND.n824 GND.n819 0.152939
R11300 GND.n825 GND.n824 0.152939
R11301 GND.n826 GND.n825 0.152939
R11302 GND.n827 GND.n826 0.152939
R11303 GND.n832 GND.n827 0.152939
R11304 GND.n833 GND.n832 0.152939
R11305 GND.n834 GND.n833 0.152939
R11306 GND.n835 GND.n834 0.152939
R11307 GND.n840 GND.n835 0.152939
R11308 GND.n841 GND.n840 0.152939
R11309 GND.n842 GND.n841 0.152939
R11310 GND.n843 GND.n842 0.152939
R11311 GND.n848 GND.n843 0.152939
R11312 GND.n849 GND.n848 0.152939
R11313 GND.n850 GND.n849 0.152939
R11314 GND.n851 GND.n850 0.152939
R11315 GND.n856 GND.n851 0.152939
R11316 GND.n857 GND.n856 0.152939
R11317 GND.n858 GND.n857 0.152939
R11318 GND.n859 GND.n858 0.152939
R11319 GND.n864 GND.n859 0.152939
R11320 GND.n865 GND.n864 0.152939
R11321 GND.n866 GND.n865 0.152939
R11322 GND.n867 GND.n866 0.152939
R11323 GND.n4219 GND.n4218 0.152939
R11324 GND.n4219 GND.n2242 0.152939
R11325 GND.n4283 GND.n2242 0.152939
R11326 GND.n4284 GND.n4283 0.152939
R11327 GND.n4286 GND.n4284 0.152939
R11328 GND.n4286 GND.n4285 0.152939
R11329 GND.n4285 GND.n2219 0.152939
R11330 GND.n4308 GND.n2219 0.152939
R11331 GND.n4309 GND.n4308 0.152939
R11332 GND.n4311 GND.n4309 0.152939
R11333 GND.n4311 GND.n4310 0.152939
R11334 GND.n4310 GND.n2197 0.152939
R11335 GND.n4333 GND.n2197 0.152939
R11336 GND.n4334 GND.n4333 0.152939
R11337 GND.n4336 GND.n4334 0.152939
R11338 GND.n4336 GND.n4335 0.152939
R11339 GND.n4335 GND.n2174 0.152939
R11340 GND.n4357 GND.n2174 0.152939
R11341 GND.n4358 GND.n4357 0.152939
R11342 GND.n4359 GND.n4358 0.152939
R11343 GND.n4359 GND.n2172 0.152939
R11344 GND.n4366 GND.n2172 0.152939
R11345 GND.n4367 GND.n4366 0.152939
R11346 GND.n4368 GND.n4367 0.152939
R11347 GND.n4368 GND.n44 0.152939
R11348 GND.n6542 GND.n45 0.152939
R11349 GND.n6538 GND.n45 0.152939
R11350 GND.n6538 GND.n6537 0.152939
R11351 GND.n6537 GND.n6536 0.152939
R11352 GND.n6536 GND.n51 0.152939
R11353 GND.n6532 GND.n51 0.152939
R11354 GND.n6532 GND.n6531 0.152939
R11355 GND.n6531 GND.n6530 0.152939
R11356 GND.n6530 GND.n56 0.152939
R11357 GND.n6526 GND.n56 0.152939
R11358 GND.n6526 GND.n6525 0.152939
R11359 GND.n6525 GND.n6524 0.152939
R11360 GND.n6524 GND.n61 0.152939
R11361 GND.n6520 GND.n61 0.152939
R11362 GND.n6520 GND.n6519 0.152939
R11363 GND.n6519 GND.n6518 0.152939
R11364 GND.n6518 GND.n66 0.152939
R11365 GND.n6514 GND.n66 0.152939
R11366 GND.n6514 GND.n6513 0.152939
R11367 GND.n6513 GND.n6512 0.152939
R11368 GND.n6512 GND.n71 0.152939
R11369 GND.n6508 GND.n71 0.152939
R11370 GND.n6508 GND.n6507 0.152939
R11371 GND.n6507 GND.n6506 0.152939
R11372 GND.n6506 GND.n76 0.152939
R11373 GND.n2049 GND.n1998 0.152939
R11374 GND.n2045 GND.n1998 0.152939
R11375 GND.n2045 GND.n2044 0.152939
R11376 GND.n2044 GND.n2043 0.152939
R11377 GND.n2043 GND.n2003 0.152939
R11378 GND.n2039 GND.n2003 0.152939
R11379 GND.n2039 GND.n2038 0.152939
R11380 GND.n2038 GND.n2037 0.152939
R11381 GND.n2037 GND.n2009 0.152939
R11382 GND.n2033 GND.n2009 0.152939
R11383 GND.n2033 GND.n2032 0.152939
R11384 GND.n2032 GND.n2031 0.152939
R11385 GND.n2031 GND.n2015 0.152939
R11386 GND.n2027 GND.n2015 0.152939
R11387 GND.n2027 GND.n2026 0.152939
R11388 GND.n2026 GND.n2025 0.152939
R11389 GND.n6498 GND.n87 0.152939
R11390 GND.n6494 GND.n87 0.152939
R11391 GND.n6494 GND.n6493 0.152939
R11392 GND.n6493 GND.n6492 0.152939
R11393 GND.n6492 GND.n91 0.152939
R11394 GND.n6488 GND.n91 0.152939
R11395 GND.n6488 GND.n6487 0.152939
R11396 GND.n6487 GND.n6486 0.152939
R11397 GND.n6486 GND.n96 0.152939
R11398 GND.n6482 GND.n96 0.152939
R11399 GND.n6482 GND.n6481 0.152939
R11400 GND.n6481 GND.n6480 0.152939
R11401 GND.n6480 GND.n101 0.152939
R11402 GND.n6476 GND.n101 0.152939
R11403 GND.n6476 GND.n6475 0.152939
R11404 GND.n6475 GND.n6474 0.152939
R11405 GND.n6474 GND.n106 0.152939
R11406 GND.n6470 GND.n106 0.152939
R11407 GND.n6470 GND.n6469 0.152939
R11408 GND.n6469 GND.n6468 0.152939
R11409 GND.n6468 GND.n114 0.152939
R11410 GND.n6464 GND.n114 0.152939
R11411 GND.n6464 GND.n6463 0.152939
R11412 GND.n6463 GND.n6462 0.152939
R11413 GND.n6462 GND.n119 0.152939
R11414 GND.n6458 GND.n119 0.152939
R11415 GND.n6458 GND.n6457 0.152939
R11416 GND.n6457 GND.n6456 0.152939
R11417 GND.n6456 GND.n124 0.152939
R11418 GND.n6452 GND.n124 0.152939
R11419 GND.n6452 GND.n6451 0.152939
R11420 GND.n6451 GND.n6450 0.152939
R11421 GND.n6450 GND.n129 0.152939
R11422 GND.n134 GND.n129 0.152939
R11423 GND.n4216 GND.n2248 0.152939
R11424 GND.n4212 GND.n2248 0.152939
R11425 GND.n4212 GND.n4211 0.152939
R11426 GND.n4211 GND.n4210 0.152939
R11427 GND.n4210 GND.n2255 0.152939
R11428 GND.n4206 GND.n2255 0.152939
R11429 GND.n4206 GND.n4205 0.152939
R11430 GND.n4205 GND.n4204 0.152939
R11431 GND.n4204 GND.n2263 0.152939
R11432 GND.n4200 GND.n2263 0.152939
R11433 GND.n4200 GND.n4199 0.152939
R11434 GND.n4199 GND.n4198 0.152939
R11435 GND.n4198 GND.n2271 0.152939
R11436 GND.n4194 GND.n2271 0.152939
R11437 GND.n4194 GND.n4193 0.152939
R11438 GND.n4193 GND.n4192 0.152939
R11439 GND.n3518 GND.n2831 0.152939
R11440 GND.n3524 GND.n2831 0.152939
R11441 GND.n3525 GND.n3524 0.152939
R11442 GND.n3526 GND.n3525 0.152939
R11443 GND.n3526 GND.n2829 0.152939
R11444 GND.n3532 GND.n2829 0.152939
R11445 GND.n3533 GND.n3532 0.152939
R11446 GND.n3534 GND.n3533 0.152939
R11447 GND.n3534 GND.n2825 0.152939
R11448 GND.n3540 GND.n2825 0.152939
R11449 GND.n3541 GND.n3540 0.152939
R11450 GND.n3542 GND.n3541 0.152939
R11451 GND.n3542 GND.n2821 0.152939
R11452 GND.n3548 GND.n2821 0.152939
R11453 GND.n3549 GND.n3548 0.152939
R11454 GND.n3550 GND.n3549 0.152939
R11455 GND.n3550 GND.n2819 0.152939
R11456 GND.n3556 GND.n2819 0.152939
R11457 GND.n3557 GND.n3556 0.152939
R11458 GND.n3558 GND.n3557 0.152939
R11459 GND.n3558 GND.n2710 0.152939
R11460 GND.n3659 GND.n2710 0.152939
R11461 GND.n3660 GND.n3659 0.152939
R11462 GND.n3661 GND.n3660 0.152939
R11463 GND.n3661 GND.n2704 0.152939
R11464 GND.n3706 GND.n2704 0.152939
R11465 GND.n3707 GND.n3706 0.152939
R11466 GND.n3708 GND.n3707 0.152939
R11467 GND.n3708 GND.n2699 0.152939
R11468 GND.n3740 GND.n2699 0.152939
R11469 GND.n3740 GND.n3739 0.152939
R11470 GND.n3739 GND.n3738 0.152939
R11471 GND.n3738 GND.n2700 0.152939
R11472 GND.n3734 GND.n2700 0.152939
R11473 GND.n3734 GND.n3733 0.152939
R11474 GND.n3733 GND.n3732 0.152939
R11475 GND.n3732 GND.n2672 0.152939
R11476 GND.n3795 GND.n2672 0.152939
R11477 GND.n3796 GND.n3795 0.152939
R11478 GND.n3806 GND.n3796 0.152939
R11479 GND.n3806 GND.n3805 0.152939
R11480 GND.n3805 GND.n3804 0.152939
R11481 GND.n3804 GND.n3798 0.152939
R11482 GND.n3798 GND.n3797 0.152939
R11483 GND.n3797 GND.n2660 0.152939
R11484 GND.n3843 GND.n2660 0.152939
R11485 GND.n3844 GND.n3843 0.152939
R11486 GND.n3849 GND.n3844 0.152939
R11487 GND.n3849 GND.n3848 0.152939
R11488 GND.n3848 GND.n3847 0.152939
R11489 GND.n3847 GND.n2648 0.152939
R11490 GND.n3879 GND.n2648 0.152939
R11491 GND.n3880 GND.n3879 0.152939
R11492 GND.n3902 GND.n3880 0.152939
R11493 GND.n3902 GND.n3901 0.152939
R11494 GND.n3901 GND.n3900 0.152939
R11495 GND.n3900 GND.n3881 0.152939
R11496 GND.n3896 GND.n3881 0.152939
R11497 GND.n3896 GND.n3895 0.152939
R11498 GND.n3895 GND.n3894 0.152939
R11499 GND.n3894 GND.n3887 0.152939
R11500 GND.n3890 GND.n3887 0.152939
R11501 GND.n3890 GND.n3889 0.152939
R11502 GND.n3889 GND.n2631 0.152939
R11503 GND.n3968 GND.n2631 0.152939
R11504 GND.n3969 GND.n3968 0.152939
R11505 GND.n3970 GND.n3969 0.152939
R11506 GND.n3970 GND.n2628 0.152939
R11507 GND.n3975 GND.n2628 0.152939
R11508 GND.n3976 GND.n3975 0.152939
R11509 GND.n3977 GND.n3976 0.152939
R11510 GND.n3977 GND.n2610 0.152939
R11511 GND.n4001 GND.n2610 0.152939
R11512 GND.n4002 GND.n4001 0.152939
R11513 GND.n4004 GND.n4002 0.152939
R11514 GND.n4004 GND.n4003 0.152939
R11515 GND.n4003 GND.n2300 0.152939
R11516 GND.n4147 GND.n2300 0.152939
R11517 GND.n4148 GND.n4147 0.152939
R11518 GND.n4149 GND.n4148 0.152939
R11519 GND.n4149 GND.n2294 0.152939
R11520 GND.n4155 GND.n2294 0.152939
R11521 GND.n4156 GND.n4155 0.152939
R11522 GND.n4157 GND.n4156 0.152939
R11523 GND.n4157 GND.n2292 0.152939
R11524 GND.n4163 GND.n2292 0.152939
R11525 GND.n4164 GND.n4163 0.152939
R11526 GND.n4165 GND.n4164 0.152939
R11527 GND.n4165 GND.n2287 0.152939
R11528 GND.n4171 GND.n2287 0.152939
R11529 GND.n4172 GND.n4171 0.152939
R11530 GND.n4173 GND.n4172 0.152939
R11531 GND.n4173 GND.n2283 0.152939
R11532 GND.n4179 GND.n2283 0.152939
R11533 GND.n4180 GND.n4179 0.152939
R11534 GND.n4181 GND.n4180 0.152939
R11535 GND.n4181 GND.n2281 0.152939
R11536 GND.n4187 GND.n2281 0.152939
R11537 GND.n3479 GND.n3478 0.152939
R11538 GND.n3480 GND.n3479 0.152939
R11539 GND.n3480 GND.n2840 0.152939
R11540 GND.n3488 GND.n2840 0.152939
R11541 GND.n3489 GND.n3488 0.152939
R11542 GND.n3490 GND.n3489 0.152939
R11543 GND.n3490 GND.n2838 0.152939
R11544 GND.n3498 GND.n2838 0.152939
R11545 GND.n3499 GND.n3498 0.152939
R11546 GND.n3500 GND.n3499 0.152939
R11547 GND.n3500 GND.n2836 0.152939
R11548 GND.n3508 GND.n2836 0.152939
R11549 GND.n3509 GND.n3508 0.152939
R11550 GND.n3510 GND.n3509 0.152939
R11551 GND.n3510 GND.n2832 0.152939
R11552 GND.n3517 GND.n2832 0.152939
R11553 GND.n3247 GND.n3246 0.152939
R11554 GND.n3247 GND.n2932 0.152939
R11555 GND.n3295 GND.n2932 0.152939
R11556 GND.n3296 GND.n3295 0.152939
R11557 GND.n3298 GND.n3296 0.152939
R11558 GND.n3298 GND.n3297 0.152939
R11559 GND.n3297 GND.n2904 0.152939
R11560 GND.n3385 GND.n2904 0.152939
R11561 GND.n3386 GND.n3385 0.152939
R11562 GND.n3388 GND.n3386 0.152939
R11563 GND.n3388 GND.n3387 0.152939
R11564 GND.n3387 GND.n2884 0.152939
R11565 GND.n3410 GND.n2884 0.152939
R11566 GND.n3411 GND.n3410 0.152939
R11567 GND.n3413 GND.n3411 0.152939
R11568 GND.n3413 GND.n3412 0.152939
R11569 GND.n3412 GND.n2862 0.152939
R11570 GND.n3435 GND.n2862 0.152939
R11571 GND.n3436 GND.n3435 0.152939
R11572 GND.n3444 GND.n3436 0.152939
R11573 GND.n3444 GND.n3443 0.152939
R11574 GND.n3443 GND.n3442 0.152939
R11575 GND.n3442 GND.n3437 0.152939
R11576 GND.n3437 GND.n2842 0.152939
R11577 GND.n3467 GND.n2842 0.152939
R11578 GND.n5096 GND.n1174 0.152939
R11579 GND.n5092 GND.n1174 0.152939
R11580 GND.n5092 GND.n5091 0.152939
R11581 GND.n5091 GND.n5090 0.152939
R11582 GND.n5090 GND.n1178 0.152939
R11583 GND.n5086 GND.n1178 0.152939
R11584 GND.n5086 GND.n5085 0.152939
R11585 GND.n5085 GND.n5084 0.152939
R11586 GND.n5084 GND.n1183 0.152939
R11587 GND.n5080 GND.n1183 0.152939
R11588 GND.n5080 GND.n5079 0.152939
R11589 GND.n5079 GND.n5078 0.152939
R11590 GND.n5078 GND.n1188 0.152939
R11591 GND.n5073 GND.n5072 0.152939
R11592 GND.n5072 GND.n5071 0.152939
R11593 GND.n5071 GND.n1198 0.152939
R11594 GND.n5067 GND.n1198 0.152939
R11595 GND.n5067 GND.n5066 0.152939
R11596 GND.n5066 GND.n5065 0.152939
R11597 GND.n5065 GND.n1203 0.152939
R11598 GND.n5061 GND.n1203 0.152939
R11599 GND.n5061 GND.n5060 0.152939
R11600 GND.n5060 GND.n5059 0.152939
R11601 GND.n5059 GND.n1208 0.152939
R11602 GND.n5055 GND.n1208 0.152939
R11603 GND.n5055 GND.n5054 0.152939
R11604 GND.n5054 GND.n5053 0.152939
R11605 GND.n5053 GND.n1213 0.152939
R11606 GND.n5049 GND.n1213 0.152939
R11607 GND.n5049 GND.n5048 0.152939
R11608 GND.n5048 GND.n5047 0.152939
R11609 GND.n5192 GND.n1010 0.152939
R11610 GND.n3070 GND.n1010 0.152939
R11611 GND.n3070 GND.n3067 0.152939
R11612 GND.n3076 GND.n3067 0.152939
R11613 GND.n3077 GND.n3076 0.152939
R11614 GND.n3078 GND.n3077 0.152939
R11615 GND.n3078 GND.n3063 0.152939
R11616 GND.n3084 GND.n3063 0.152939
R11617 GND.n3085 GND.n3084 0.152939
R11618 GND.n3086 GND.n3085 0.152939
R11619 GND.n3086 GND.n3059 0.152939
R11620 GND.n3092 GND.n3059 0.152939
R11621 GND.n3093 GND.n3092 0.152939
R11622 GND.n3094 GND.n3093 0.152939
R11623 GND.n3094 GND.n3052 0.152939
R11624 GND.n3098 GND.n3052 0.152939
R11625 GND.n3101 GND.n3100 0.152939
R11626 GND.n3102 GND.n3101 0.152939
R11627 GND.n3102 GND.n3048 0.152939
R11628 GND.n3110 GND.n3048 0.152939
R11629 GND.n3111 GND.n3110 0.152939
R11630 GND.n3112 GND.n3111 0.152939
R11631 GND.n3112 GND.n3040 0.152939
R11632 GND.n3155 GND.n3040 0.152939
R11633 GND.n3156 GND.n3155 0.152939
R11634 GND.n3163 GND.n3156 0.152939
R11635 GND.n3163 GND.n3162 0.152939
R11636 GND.n3162 GND.n3161 0.152939
R11637 GND.n3161 GND.n3157 0.152939
R11638 GND.n3157 GND.n3008 0.152939
R11639 GND.n3195 GND.n3008 0.152939
R11640 GND.n3196 GND.n3195 0.152939
R11641 GND.n3199 GND.n3196 0.152939
R11642 GND.n3199 GND.n3198 0.152939
R11643 GND.n3198 GND.n3197 0.152939
R11644 GND.n3197 GND.n2980 0.152939
R11645 GND.n3233 GND.n2980 0.152939
R11646 GND.n3234 GND.n3233 0.152939
R11647 GND.n3235 GND.n3234 0.152939
R11648 GND.n3235 GND.n2978 0.152939
R11649 GND.n3244 GND.n2978 0.152939
R11650 GND.n3306 GND.n2925 0.131598
R11651 GND.n4435 GND.n4434 0.131598
R11652 GND.n2540 GND.n2539 0.124411
R11653 GND.n5045 GND.n5044 0.124411
R11654 GND.n4217 GND.n4216 0.108732
R11655 GND.n3478 GND.n3468 0.108732
R11656 GND.n2141 GND.n2125 0.0767195
R11657 GND.n2154 GND.n2141 0.0767195
R11658 GND.n3288 GND.n2914 0.0767195
R11659 GND.n3288 GND.n2943 0.0767195
R11660 GND.n6543 GND.n44 0.0695946
R11661 GND.n6543 GND.n6542 0.0695946
R11662 GND.n3246 GND.n3245 0.0695946
R11663 GND.n3245 GND.n3244 0.0695946
R11664 GND.n2540 GND.n2438 0.0548478
R11665 GND.n2051 GND.n2050 0.0548478
R11666 GND.n5193 GND.n1009 0.0548478
R11667 GND.n5045 GND.n1164 0.0548478
R11668 GND.n2539 GND.n2439 0.044054
R11669 GND.n2532 GND.n2439 0.044054
R11670 GND.n2532 GND.n2531 0.044054
R11671 GND.n5044 GND.n1220 0.044054
R11672 GND.n5040 GND.n1220 0.044054
R11673 GND.n5040 GND.n5039 0.044054
R11674 GND.n2531 GND.n2530 0.0411504
R11675 GND.n5039 GND.n5038 0.0411504
R11676 GND.n2438 GND.n1900 0.0344674
R11677 GND.n4630 GND.n1900 0.0344674
R11678 GND.n4630 GND.n1901 0.0344674
R11679 GND.n4626 GND.n1901 0.0344674
R11680 GND.n4626 GND.n4625 0.0344674
R11681 GND.n4625 GND.n4624 0.0344674
R11682 GND.n4624 GND.n1909 0.0344674
R11683 GND.n4620 GND.n1909 0.0344674
R11684 GND.n4620 GND.n4619 0.0344674
R11685 GND.n4619 GND.n4618 0.0344674
R11686 GND.n4618 GND.n1917 0.0344674
R11687 GND.n4614 GND.n1917 0.0344674
R11688 GND.n4614 GND.n4613 0.0344674
R11689 GND.n4613 GND.n4612 0.0344674
R11690 GND.n4612 GND.n1925 0.0344674
R11691 GND.n4608 GND.n1925 0.0344674
R11692 GND.n4608 GND.n4607 0.0344674
R11693 GND.n4607 GND.n4606 0.0344674
R11694 GND.n4606 GND.n1933 0.0344674
R11695 GND.n4602 GND.n1933 0.0344674
R11696 GND.n4602 GND.n4601 0.0344674
R11697 GND.n4601 GND.n4600 0.0344674
R11698 GND.n4600 GND.n1941 0.0344674
R11699 GND.n4596 GND.n1941 0.0344674
R11700 GND.n4596 GND.n4595 0.0344674
R11701 GND.n4595 GND.n4594 0.0344674
R11702 GND.n4594 GND.n1949 0.0344674
R11703 GND.n4590 GND.n1949 0.0344674
R11704 GND.n4590 GND.n4589 0.0344674
R11705 GND.n4589 GND.n4588 0.0344674
R11706 GND.n4588 GND.n1957 0.0344674
R11707 GND.n4584 GND.n1957 0.0344674
R11708 GND.n4584 GND.n4583 0.0344674
R11709 GND.n4583 GND.n4582 0.0344674
R11710 GND.n4582 GND.n1965 0.0344674
R11711 GND.n4578 GND.n1965 0.0344674
R11712 GND.n4578 GND.n4577 0.0344674
R11713 GND.n4577 GND.n4576 0.0344674
R11714 GND.n4576 GND.n1973 0.0344674
R11715 GND.n4572 GND.n1973 0.0344674
R11716 GND.n4572 GND.n4571 0.0344674
R11717 GND.n4571 GND.n4570 0.0344674
R11718 GND.n4570 GND.n1981 0.0344674
R11719 GND.n4566 GND.n1981 0.0344674
R11720 GND.n4566 GND.n4565 0.0344674
R11721 GND.n4565 GND.n4564 0.0344674
R11722 GND.n4564 GND.n1989 0.0344674
R11723 GND.n4560 GND.n1989 0.0344674
R11724 GND.n4560 GND.n4559 0.0344674
R11725 GND.n4559 GND.n4558 0.0344674
R11726 GND.n4558 GND.n2051 0.0344674
R11727 GND.n1067 GND.n1009 0.0344674
R11728 GND.n1067 GND.n1062 0.0344674
R11729 GND.n1072 GND.n1062 0.0344674
R11730 GND.n1072 GND.n1059 0.0344674
R11731 GND.n5171 GND.n1059 0.0344674
R11732 GND.n5171 GND.n1060 0.0344674
R11733 GND.n5167 GND.n1060 0.0344674
R11734 GND.n5167 GND.n5166 0.0344674
R11735 GND.n5166 GND.n5165 0.0344674
R11736 GND.n5165 GND.n1081 0.0344674
R11737 GND.n5161 GND.n1081 0.0344674
R11738 GND.n5161 GND.n5160 0.0344674
R11739 GND.n5160 GND.n5159 0.0344674
R11740 GND.n5159 GND.n1089 0.0344674
R11741 GND.n5155 GND.n1089 0.0344674
R11742 GND.n5155 GND.n5154 0.0344674
R11743 GND.n5154 GND.n5153 0.0344674
R11744 GND.n5153 GND.n1097 0.0344674
R11745 GND.n5149 GND.n1097 0.0344674
R11746 GND.n5149 GND.n5148 0.0344674
R11747 GND.n5148 GND.n5147 0.0344674
R11748 GND.n5147 GND.n1105 0.0344674
R11749 GND.n5143 GND.n1105 0.0344674
R11750 GND.n5143 GND.n5142 0.0344674
R11751 GND.n5142 GND.n5141 0.0344674
R11752 GND.n5141 GND.n1113 0.0344674
R11753 GND.n5137 GND.n1113 0.0344674
R11754 GND.n5137 GND.n5136 0.0344674
R11755 GND.n5136 GND.n5135 0.0344674
R11756 GND.n5135 GND.n1121 0.0344674
R11757 GND.n5131 GND.n1121 0.0344674
R11758 GND.n5131 GND.n5130 0.0344674
R11759 GND.n5130 GND.n5129 0.0344674
R11760 GND.n5129 GND.n1129 0.0344674
R11761 GND.n5125 GND.n1129 0.0344674
R11762 GND.n5125 GND.n5124 0.0344674
R11763 GND.n5124 GND.n5123 0.0344674
R11764 GND.n5123 GND.n1137 0.0344674
R11765 GND.n5119 GND.n1137 0.0344674
R11766 GND.n5119 GND.n5118 0.0344674
R11767 GND.n5118 GND.n5117 0.0344674
R11768 GND.n5117 GND.n1145 0.0344674
R11769 GND.n5113 GND.n1145 0.0344674
R11770 GND.n5113 GND.n5112 0.0344674
R11771 GND.n5112 GND.n5111 0.0344674
R11772 GND.n5111 GND.n1153 0.0344674
R11773 GND.n5107 GND.n1153 0.0344674
R11774 GND.n5107 GND.n5106 0.0344674
R11775 GND.n5106 GND.n5105 0.0344674
R11776 GND.n5105 GND.n1161 0.0344674
R11777 GND.n1164 GND.n1161 0.0344674
R11778 GND.n2527 GND.n2526 0.0343753
R11779 GND.n2493 GND.n2247 0.0343753
R11780 GND.n5035 GND.n5034 0.0343753
R11781 GND.n3473 GND.n3472 0.0343753
R11782 GND.n2527 GND.n2443 0.0306491
R11783 GND.n5035 GND.n1225 0.0306491
R11784 GND.n2525 GND.n2448 0.0303103
R11785 GND.n2522 GND.n2521 0.0303103
R11786 GND.n2518 GND.n2451 0.0303103
R11787 GND.n2517 GND.n2460 0.0303103
R11788 GND.n2514 GND.n2513 0.0303103
R11789 GND.n2510 GND.n2467 0.0303103
R11790 GND.n2509 GND.n2474 0.0303103
R11791 GND.n2506 GND.n2505 0.0303103
R11792 GND.n2497 GND.n2480 0.0303103
R11793 GND.n2496 GND.n2485 0.0303103
R11794 GND.n5033 GND.n1229 0.0303103
R11795 GND.n1251 GND.n1250 0.0303103
R11796 GND.n5026 GND.n5025 0.0303103
R11797 GND.n5022 GND.n1252 0.0303103
R11798 GND.n5021 GND.n1257 0.0303103
R11799 GND.n5018 GND.n5017 0.0303103
R11800 GND.n5014 GND.n1261 0.0303103
R11801 GND.n5013 GND.n1265 0.0303103
R11802 GND.n5010 GND.n5009 0.0303103
R11803 GND.n1275 GND.n1271 0.0303103
R11804 GND.n4436 GND.n4435 0.0218415
R11805 GND.n3222 GND.n2925 0.0218415
R11806 GND.n4217 GND.n2247 0.0103238
R11807 GND.n3473 GND.n3468 0.0103238
R11808 GND.n2526 GND.n2525 0.00456504
R11809 GND.n2522 GND.n2448 0.00456504
R11810 GND.n2521 GND.n2451 0.00456504
R11811 GND.n2518 GND.n2517 0.00456504
R11812 GND.n2514 GND.n2460 0.00456504
R11813 GND.n2513 GND.n2467 0.00456504
R11814 GND.n2510 GND.n2509 0.00456504
R11815 GND.n2506 GND.n2474 0.00456504
R11816 GND.n2505 GND.n2480 0.00456504
R11817 GND.n2497 GND.n2496 0.00456504
R11818 GND.n2493 GND.n2485 0.00456504
R11819 GND.n5034 GND.n5033 0.00456504
R11820 GND.n1250 GND.n1229 0.00456504
R11821 GND.n5026 GND.n1251 0.00456504
R11822 GND.n5025 GND.n1252 0.00456504
R11823 GND.n5022 GND.n5021 0.00456504
R11824 GND.n5018 GND.n1257 0.00456504
R11825 GND.n5017 GND.n1261 0.00456504
R11826 GND.n5014 GND.n5013 0.00456504
R11827 GND.n5010 GND.n1265 0.00456504
R11828 GND.n5009 GND.n1271 0.00456504
R11829 GND.n3472 GND.n1275 0.00456504
R11830 GND.n2530 GND.n2443 0.00422629
R11831 GND.n5038 GND.n1225 0.00422629
R11832 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t14 167.274
R11833 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.t12 164.87
R11834 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.t11 164.87
R11835 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.t13 164.87
R11836 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t10 164.87
R11837 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t4 124.242
R11838 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t2 121.838
R11839 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t6 121.838
R11840 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.t8 121.838
R11841 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t0 121.838
R11842 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t5 92.89
R11843 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t3 92.0898
R11844 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t7 92.0898
R11845 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t9 92.0898
R11846 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t1 92.0898
R11847 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 5.4711
R11848 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 4.30779
R11849 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n4 4.24998
R11850 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 2.40335
R11851 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 2.40335
R11852 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 2.40335
R11853 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 2.40332
R11854 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 2.40332
R11855 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n0 1.65702
R11856 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 0.800888
R11857 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 0.800888
R11858 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 0.800888
R11859 DIFFPAIR_BIAS DIFFPAIR_BIAS.n13 0.68425
R11860 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 0.456103
R11861 a_n2675_n4106.n0 a_n2675_n4106.t5 160.166
R11862 a_n2675_n4106.n7 a_n2675_n4106.t4 159.581
R11863 a_n2675_n4106.n8 a_n2675_n4106.t8 159.581
R11864 a_n2675_n4106.n9 a_n2675_n4106.t6 159.581
R11865 a_n2675_n4106.t7 a_n2675_n4106.n0 159.581
R11866 a_n2675_n4106.n5 a_n2675_n4106.t2 48.8949
R11867 a_n2675_n4106.n4 a_n2675_n4106.t0 48.8949
R11868 a_n2675_n4106.n2 a_n2675_n4106.t1 48.8949
R11869 a_n2675_n4106.n1 a_n2675_n4106.t3 48.8948
R11870 a_n2675_n4106.n3 a_n2675_n4106.n2 13.333
R11871 a_n2675_n4106.n6 a_n2675_n4106.n1 12.5485
R11872 a_n2675_n4106.n4 a_n2675_n4106.n3 6.40495
R11873 a_n2675_n4106.n6 a_n2675_n4106.n5 5.62047
R11874 a_n2675_n4106.n7 a_n2675_n4106.n6 2.48737
R11875 a_n2675_n4106.n3 a_n2675_n4106.n0 2.39823
R11876 a_n2675_n4106.n0 a_n2675_n4106.n9 1.01697
R11877 a_n2675_n4106.n2 a_n2675_n4106.n1 0.989006
R11878 a_n2675_n4106.n5 a_n2675_n4106.n4 0.989006
R11879 a_n2675_n4106.n9 a_n2675_n4106.n8 0.800888
R11880 a_n2675_n4106.n8 a_n2675_n4106.n7 0.800888
R11881 a_n6918_10482.n7 a_n6918_10482.t3 188.107
R11882 a_n6918_10482.n12 a_n6918_10482.t1 187.393
R11883 a_n6918_10482.n19 a_n6918_10482.t5 99.7812
R11884 a_n6918_10482.t4 a_n6918_10482.n19 68.4828
R11885 a_n6918_10482.n9 a_n6918_10482.t0 55.2817
R11886 a_n6918_10482.n16 a_n6918_10482.t2 55.2817
R11887 a_n6918_10482.n17 a_n6918_10482.t12 55.2817
R11888 a_n6918_10482.n8 a_n6918_10482.t21 55.2817
R11889 a_n6918_10482.n18 a_n6918_10482.n2 73.7168
R11890 a_n6918_10482.n6 a_n6918_10482.n0 114.169
R11891 a_n6918_10482.n19 a_n6918_10482.n9 24.4495
R11892 a_n6918_10482.n5 a_n6918_10482.n14 73.7164
R11893 a_n6918_10482.n4 a_n6918_10482.n15 73.7164
R11894 a_n6918_10482.n12 a_n6918_10482.n17 19.39
R11895 a_n6918_10482.n8 a_n6918_10482.n7 18.9658
R11896 a_n6918_10482.n12 a_n6918_10482.n9 17.3332
R11897 a_n6918_10482.n3 a_n6918_10482.t9 50.5488
R11898 a_n6918_10482.n2 a_n6918_10482.t7 45.9874
R11899 a_n6918_10482.n18 a_n6918_10482.t13 16.4939
R11900 a_n6918_10482.n13 a_n6918_10482.t19 50.5481
R11901 a_n6918_10482.n10 a_n6918_10482.t14 50.5488
R11902 a_n6918_10482.n14 a_n6918_10482.t22 16.4939
R11903 a_n6918_10482.n5 a_n6918_10482.t20 45.9884
R11904 a_n6918_10482.n3 a_n6918_10482.t8 50.5481
R11905 a_n6918_10482.n1 a_n6918_10482.t10 50.5488
R11906 a_n6918_10482.n0 a_n6918_10482.t23 42.7465
R11907 a_n6918_10482.n6 a_n6918_10482.t17 27.4574
R11908 a_n6918_10482.n3 a_n6918_10482.t18 50.5481
R11909 a_n6918_10482.n11 a_n6918_10482.t15 50.5488
R11910 a_n6918_10482.n15 a_n6918_10482.t16 16.4939
R11911 a_n6918_10482.n4 a_n6918_10482.t11 45.9884
R11912 a_n6918_10482.n1 a_n6918_10482.t6 50.5481
R11913 a_n6918_10482.n16 a_n6918_10482.n7 16.0756
R11914 a_n6918_10482.n17 a_n6918_10482.n16 7.71512
R11915 a_n6918_10482.n3 a_n6918_10482.n2 2.45052
R11916 a_n6918_10482.n18 a_n6918_10482.n13 54.8801
R11917 a_n6918_10482.n10 a_n6918_10482.n14 54.8794
R11918 a_n6918_10482.n1 a_n6918_10482.n0 5.88345
R11919 a_n6918_10482.n6 a_n6918_10482.n3 25.356
R11920 a_n6918_10482.n11 a_n6918_10482.n15 54.8794
R11921 a_n6918_10482.n7 a_n6918_10482.n3 10.5056
R11922 a_n6918_10482.n1 a_n6918_10482.n3 9.75172
R11923 a_n6918_10482.n1 a_n6918_10482.n12 8.82378
R11924 a_n6918_10482.n5 a_n6918_10482.n3 8.2281
R11925 a_n6918_10482.n4 a_n6918_10482.n1 8.2281
R11926 a_n6918_10482.n9 a_n6918_10482.n8 7.67724
R11927 a_n6918_10482.n1 a_n6918_10482.n11 6.93412
R11928 a_n6918_10482.n3 a_n6918_10482.n13 6.9341
R11929 a_n6918_10482.n3 a_n6918_10482.n10 6.782
R11930 a_n2500_9133.n1 a_n2500_9133.t2 201.595
R11931 a_n2500_9133.n1 a_n2500_9133.t10 187.512
R11932 a_n2500_9133.n0 a_n2500_9133.t6 179.327
R11933 a_n2500_9133.n0 a_n2500_9133.t1 178.219
R11934 a_n2500_9133.n0 a_n2500_9133.t5 178.219
R11935 a_n2500_9133.n0 a_n2500_9133.t8 178.219
R11936 a_n2500_9133.n0 a_n2500_9133.n2 148.534
R11937 a_n2500_9133.n0 a_n2500_9133.n3 148.534
R11938 a_n2500_9133.n2 a_n2500_9133.t7 29.6854
R11939 a_n2500_9133.n2 a_n2500_9133.t4 29.6854
R11940 a_n2500_9133.n3 a_n2500_9133.t3 29.6854
R11941 a_n2500_9133.n3 a_n2500_9133.t9 29.6854
R11942 a_n2500_9133.n1 a_n2500_9133.n0 12.3645
R11943 a_n2500_9133.t0 a_n2500_9133.n1 11.3761
R11944 VDD.n2477 VDD.n299 455.123
R11945 VDD.n2726 VDD.n103 455.123
R11946 VDD.n2622 VDD.n101 455.123
R11947 VDD.n2479 VDD.n297 455.123
R11948 VDD.n1523 VDD.n917 455.123
R11949 VDD.n1526 VDD.n1525 455.123
R11950 VDD.n1278 VDD.n1071 455.123
R11951 VDD.n1276 VDD.n1073 455.123
R11952 VDD.n2321 VDD.n387 302.928
R11953 VDD.n2293 VDD.n402 302.928
R11954 VDD.n2096 VDD.n1925 302.928
R11955 VDD.n2127 VDD.n530 302.928
R11956 VDD.n1878 VDD.n565 302.928
R11957 VDD.n1848 VDD.n1847 302.928
R11958 VDD.n1671 VDD.n710 302.928
R11959 VDD.n1703 VDD.n697 302.928
R11960 VDD.n2271 VDD.n2270 302.928
R11961 VDD.n2331 VDD.n379 302.928
R11962 VDD.n2002 VDD.n2001 302.928
R11963 VDD.n2131 VDD.n534 302.928
R11964 VDD.n1917 VDD.n554 302.928
R11965 VDD.n1885 VDD.n553 302.928
R11966 VDD.n866 VDD.n718 302.928
R11967 VDD.n1706 VDD.n701 302.928
R11968 VDD.n799 VDD.t128 232.566
R11969 VDD.n557 VDD.t80 232.566
R11970 VDD.n1607 VDD.t125 232.566
R11971 VDD.n567 VDD.t117 232.566
R11972 VDD.n1933 VDD.t55 232.566
R11973 VDD.n398 VDD.t108 232.566
R11974 VDD.n2032 VDD.t121 232.566
R11975 VDD.n375 VDD.t76 232.566
R11976 VDD.n1187 VDD.t104 231.957
R11977 VDD.n1154 VDD.t95 231.957
R11978 VDD.n1232 VDD.t89 231.957
R11979 VDD.n1094 VDD.t67 231.957
R11980 VDD.n908 VDD.t71 231.957
R11981 VDD.n778 VDD.t60 231.957
R11982 VDD.n1572 VDD.t64 231.957
R11983 VDD.n728 VDD.t101 231.957
R11984 VDD.n2624 VDD.t56 231.957
R11985 VDD.n176 VDD.t129 231.957
R11986 VDD.n2676 VDD.t113 231.957
R11987 VDD.n122 VDD.t86 231.957
R11988 VDD.n315 VDD.t82 231.957
R11989 VDD.n2394 VDD.t92 231.957
R11990 VDD.n339 VDD.t110 231.957
R11991 VDD.n2364 VDD.t98 231.957
R11992 VDD.n799 VDD.t126 225.297
R11993 VDD.n557 VDD.t78 225.297
R11994 VDD.n1607 VDD.t122 225.297
R11995 VDD.n567 VDD.t116 225.297
R11996 VDD.n1933 VDD.t52 225.297
R11997 VDD.n398 VDD.t107 225.297
R11998 VDD.n2032 VDD.t119 225.297
R11999 VDD.n375 VDD.t74 225.297
R12000 VDD.n727 VDD.t15 197.161
R12001 VDD.t140 VDD.n298 197.161
R12002 VDD.n1187 VDD.t106 189.392
R12003 VDD.n1154 VDD.t97 189.392
R12004 VDD.n1232 VDD.t91 189.392
R12005 VDD.n1094 VDD.t70 189.392
R12006 VDD.n908 VDD.t72 189.392
R12007 VDD.n778 VDD.t62 189.392
R12008 VDD.n1572 VDD.t65 189.392
R12009 VDD.n728 VDD.t102 189.392
R12010 VDD.n2624 VDD.t58 189.392
R12011 VDD.n176 VDD.t130 189.392
R12012 VDD.n2676 VDD.t114 189.392
R12013 VDD.n122 VDD.t87 189.392
R12014 VDD.n315 VDD.t85 189.392
R12015 VDD.n2394 VDD.t94 189.392
R12016 VDD.n339 VDD.t112 189.392
R12017 VDD.n2364 VDD.t100 189.392
R12018 VDD.n2272 VDD.n2271 185
R12019 VDD.n2271 VDD.n384 185
R12020 VDD.n2273 VDD.n385 185
R12021 VDD.n2326 VDD.n385 185
R12022 VDD.n2275 VDD.n2274 185
R12023 VDD.n2274 VDD.n382 185
R12024 VDD.n2276 VDD.n407 185
R12025 VDD.n2286 VDD.n407 185
R12026 VDD.n2277 VDD.n415 185
R12027 VDD.n415 VDD.n405 185
R12028 VDD.n2279 VDD.n2278 185
R12029 VDD.n2280 VDD.n2279 185
R12030 VDD.n2252 VDD.n414 185
R12031 VDD.n414 VDD.n411 185
R12032 VDD.n2251 VDD.n2250 185
R12033 VDD.n2250 VDD.n2249 185
R12034 VDD.n417 VDD.n416 185
R12035 VDD.n426 VDD.n417 185
R12036 VDD.n2242 VDD.n2241 185
R12037 VDD.n2243 VDD.n2242 185
R12038 VDD.n2240 VDD.n427 185
R12039 VDD.n427 VDD.n423 185
R12040 VDD.n2239 VDD.n2238 185
R12041 VDD.n2238 VDD.n2237 185
R12042 VDD.n429 VDD.n428 185
R12043 VDD.n430 VDD.n429 185
R12044 VDD.n2230 VDD.n2229 185
R12045 VDD.n2231 VDD.n2230 185
R12046 VDD.n2228 VDD.n439 185
R12047 VDD.n439 VDD.n436 185
R12048 VDD.n2227 VDD.n2226 185
R12049 VDD.n2226 VDD.n2225 185
R12050 VDD.n441 VDD.n440 185
R12051 VDD.n442 VDD.n441 185
R12052 VDD.n2218 VDD.n2217 185
R12053 VDD.n2219 VDD.n2218 185
R12054 VDD.n2216 VDD.n450 185
R12055 VDD.n450 VDD.t19 185
R12056 VDD.n2215 VDD.n2214 185
R12057 VDD.n2214 VDD.n2213 185
R12058 VDD.n452 VDD.n451 185
R12059 VDD.n453 VDD.n452 185
R12060 VDD.n2206 VDD.n2205 185
R12061 VDD.n2207 VDD.n2206 185
R12062 VDD.n2204 VDD.n462 185
R12063 VDD.n462 VDD.n459 185
R12064 VDD.n2203 VDD.n2202 185
R12065 VDD.n2202 VDD.t23 185
R12066 VDD.n464 VDD.n463 185
R12067 VDD.n465 VDD.n464 185
R12068 VDD.n2195 VDD.n2194 185
R12069 VDD.n2196 VDD.n2195 185
R12070 VDD.n2193 VDD.n474 185
R12071 VDD.n474 VDD.n471 185
R12072 VDD.n2192 VDD.n2191 185
R12073 VDD.n2191 VDD.n2190 185
R12074 VDD.n476 VDD.n475 185
R12075 VDD.n477 VDD.n476 185
R12076 VDD.n2183 VDD.n2182 185
R12077 VDD.n2184 VDD.n2183 185
R12078 VDD.n2181 VDD.n485 185
R12079 VDD.n491 VDD.n485 185
R12080 VDD.n2180 VDD.n2179 185
R12081 VDD.n2179 VDD.n2178 185
R12082 VDD.n487 VDD.n486 185
R12083 VDD.n488 VDD.n487 185
R12084 VDD.n2171 VDD.n2170 185
R12085 VDD.n2172 VDD.n2171 185
R12086 VDD.n2169 VDD.n498 185
R12087 VDD.n498 VDD.n495 185
R12088 VDD.n2168 VDD.n2167 185
R12089 VDD.n2167 VDD.n2166 185
R12090 VDD.n500 VDD.n499 185
R12091 VDD.n501 VDD.n500 185
R12092 VDD.n2159 VDD.n2158 185
R12093 VDD.n2160 VDD.n2159 185
R12094 VDD.n2157 VDD.n510 185
R12095 VDD.n510 VDD.n507 185
R12096 VDD.n2156 VDD.n2155 185
R12097 VDD.n2155 VDD.n2154 185
R12098 VDD.n512 VDD.n511 185
R12099 VDD.n513 VDD.n512 185
R12100 VDD.n2147 VDD.n2146 185
R12101 VDD.n2148 VDD.n2147 185
R12102 VDD.n2145 VDD.n522 185
R12103 VDD.n522 VDD.n519 185
R12104 VDD.n2144 VDD.n2143 185
R12105 VDD.n2143 VDD.n2142 185
R12106 VDD.n524 VDD.n523 185
R12107 VDD.n525 VDD.n524 185
R12108 VDD.n2135 VDD.n2134 185
R12109 VDD.n2136 VDD.n2135 185
R12110 VDD.n2133 VDD.n534 185
R12111 VDD.n534 VDD.n531 185
R12112 VDD.n2132 VDD.n2131 185
R12113 VDD.n536 VDD.n535 185
R12114 VDD.n2028 VDD.n2027 185
R12115 VDD.n2026 VDD.n1932 185
R12116 VDD.n2025 VDD.n2024 185
R12117 VDD.n2023 VDD.n2022 185
R12118 VDD.n2021 VDD.n2020 185
R12119 VDD.n2019 VDD.n2018 185
R12120 VDD.n2017 VDD.n2016 185
R12121 VDD.n2015 VDD.n2014 185
R12122 VDD.n2013 VDD.n2012 185
R12123 VDD.n2011 VDD.n2010 185
R12124 VDD.n2009 VDD.n2008 185
R12125 VDD.n2007 VDD.n2006 185
R12126 VDD.n2005 VDD.n2004 185
R12127 VDD.n2003 VDD.n2002 185
R12128 VDD.n2331 VDD.n2330 185
R12129 VDD.n2333 VDD.n377 185
R12130 VDD.n2335 VDD.n2334 185
R12131 VDD.n2336 VDD.n374 185
R12132 VDD.n2339 VDD.n2338 185
R12133 VDD.n2341 VDD.n373 185
R12134 VDD.n2342 VDD.n370 185
R12135 VDD.n2345 VDD.n2344 185
R12136 VDD.n371 VDD.n369 185
R12137 VDD.n2259 VDD.n2258 185
R12138 VDD.n2261 VDD.n2260 185
R12139 VDD.n2263 VDD.n2255 185
R12140 VDD.n2265 VDD.n2264 185
R12141 VDD.n2266 VDD.n2254 185
R12142 VDD.n2268 VDD.n2267 185
R12143 VDD.n2270 VDD.n2253 185
R12144 VDD.n2329 VDD.n379 185
R12145 VDD.n384 VDD.n379 185
R12146 VDD.n2328 VDD.n2327 185
R12147 VDD.n2327 VDD.n2326 185
R12148 VDD.n381 VDD.n380 185
R12149 VDD.n382 VDD.n381 185
R12150 VDD.n1936 VDD.n406 185
R12151 VDD.n2286 VDD.n406 185
R12152 VDD.n1938 VDD.n1937 185
R12153 VDD.n1937 VDD.n405 185
R12154 VDD.n1939 VDD.n413 185
R12155 VDD.n2280 VDD.n413 185
R12156 VDD.n1941 VDD.n1940 185
R12157 VDD.n1940 VDD.n411 185
R12158 VDD.n1942 VDD.n419 185
R12159 VDD.n2249 VDD.n419 185
R12160 VDD.n1944 VDD.n1943 185
R12161 VDD.n1943 VDD.n426 185
R12162 VDD.n1945 VDD.n425 185
R12163 VDD.n2243 VDD.n425 185
R12164 VDD.n1947 VDD.n1946 185
R12165 VDD.n1946 VDD.n423 185
R12166 VDD.n1948 VDD.n432 185
R12167 VDD.n2237 VDD.n432 185
R12168 VDD.n1950 VDD.n1949 185
R12169 VDD.n1949 VDD.n430 185
R12170 VDD.n1951 VDD.n438 185
R12171 VDD.n2231 VDD.n438 185
R12172 VDD.n1953 VDD.n1952 185
R12173 VDD.n1952 VDD.n436 185
R12174 VDD.n1954 VDD.n444 185
R12175 VDD.n2225 VDD.n444 185
R12176 VDD.n1956 VDD.n1955 185
R12177 VDD.n1955 VDD.n442 185
R12178 VDD.n1957 VDD.n449 185
R12179 VDD.n2219 VDD.n449 185
R12180 VDD.n1959 VDD.n1958 185
R12181 VDD.n1958 VDD.t19 185
R12182 VDD.n1960 VDD.n455 185
R12183 VDD.n2213 VDD.n455 185
R12184 VDD.n1962 VDD.n1961 185
R12185 VDD.n1961 VDD.n453 185
R12186 VDD.n1963 VDD.n461 185
R12187 VDD.n2207 VDD.n461 185
R12188 VDD.n1965 VDD.n1964 185
R12189 VDD.n1964 VDD.n459 185
R12190 VDD.n1966 VDD.n466 185
R12191 VDD.t23 VDD.n466 185
R12192 VDD.n1968 VDD.n1967 185
R12193 VDD.n1967 VDD.n465 185
R12194 VDD.n1969 VDD.n473 185
R12195 VDD.n2196 VDD.n473 185
R12196 VDD.n1971 VDD.n1970 185
R12197 VDD.n1970 VDD.n471 185
R12198 VDD.n1972 VDD.n479 185
R12199 VDD.n2190 VDD.n479 185
R12200 VDD.n1974 VDD.n1973 185
R12201 VDD.n1973 VDD.n477 185
R12202 VDD.n1975 VDD.n484 185
R12203 VDD.n2184 VDD.n484 185
R12204 VDD.n1977 VDD.n1976 185
R12205 VDD.n1976 VDD.n491 185
R12206 VDD.n1978 VDD.n490 185
R12207 VDD.n2178 VDD.n490 185
R12208 VDD.n1980 VDD.n1979 185
R12209 VDD.n1979 VDD.n488 185
R12210 VDD.n1981 VDD.n497 185
R12211 VDD.n2172 VDD.n497 185
R12212 VDD.n1983 VDD.n1982 185
R12213 VDD.n1982 VDD.n495 185
R12214 VDD.n1984 VDD.n503 185
R12215 VDD.n2166 VDD.n503 185
R12216 VDD.n1986 VDD.n1985 185
R12217 VDD.n1985 VDD.n501 185
R12218 VDD.n1987 VDD.n509 185
R12219 VDD.n2160 VDD.n509 185
R12220 VDD.n1989 VDD.n1988 185
R12221 VDD.n1988 VDD.n507 185
R12222 VDD.n1990 VDD.n515 185
R12223 VDD.n2154 VDD.n515 185
R12224 VDD.n1992 VDD.n1991 185
R12225 VDD.n1991 VDD.n513 185
R12226 VDD.n1993 VDD.n521 185
R12227 VDD.n2148 VDD.n521 185
R12228 VDD.n1995 VDD.n1994 185
R12229 VDD.n1994 VDD.n519 185
R12230 VDD.n1996 VDD.n527 185
R12231 VDD.n2142 VDD.n527 185
R12232 VDD.n1998 VDD.n1997 185
R12233 VDD.n1997 VDD.n525 185
R12234 VDD.n1999 VDD.n533 185
R12235 VDD.n2136 VDD.n533 185
R12236 VDD.n2001 VDD.n2000 185
R12237 VDD.n2001 VDD.n531 185
R12238 VDD.n1880 VDD.n565 185
R12239 VDD.n565 VDD.n537 185
R12240 VDD.n1882 VDD.n1881 185
R12241 VDD.n1883 VDD.n1882 185
R12242 VDD.n566 VDD.n564 185
R12243 VDD.n564 VDD.n561 185
R12244 VDD.n1840 VDD.n1839 185
R12245 VDD.n1841 VDD.n1840 185
R12246 VDD.n1838 VDD.n575 185
R12247 VDD.n575 VDD.n572 185
R12248 VDD.n1837 VDD.n1836 185
R12249 VDD.n1836 VDD.n1835 185
R12250 VDD.n577 VDD.n576 185
R12251 VDD.n586 VDD.n577 185
R12252 VDD.n1823 VDD.n1822 185
R12253 VDD.n1824 VDD.n1823 185
R12254 VDD.n1821 VDD.n587 185
R12255 VDD.n593 VDD.n587 185
R12256 VDD.n1820 VDD.n1819 185
R12257 VDD.n1819 VDD.n1818 185
R12258 VDD.n589 VDD.n588 185
R12259 VDD.n590 VDD.n589 185
R12260 VDD.n1811 VDD.n1810 185
R12261 VDD.n1812 VDD.n1811 185
R12262 VDD.n1809 VDD.n600 185
R12263 VDD.n600 VDD.n597 185
R12264 VDD.n1808 VDD.n1807 185
R12265 VDD.n1807 VDD.n1806 185
R12266 VDD.n602 VDD.n601 185
R12267 VDD.n603 VDD.n602 185
R12268 VDD.n1799 VDD.n1798 185
R12269 VDD.n1800 VDD.n1799 185
R12270 VDD.n1797 VDD.n612 185
R12271 VDD.n612 VDD.n609 185
R12272 VDD.n1796 VDD.n1795 185
R12273 VDD.n1795 VDD.n1794 185
R12274 VDD.n614 VDD.n613 185
R12275 VDD.n615 VDD.n614 185
R12276 VDD.n1787 VDD.n1786 185
R12277 VDD.n1788 VDD.n1787 185
R12278 VDD.n1785 VDD.n624 185
R12279 VDD.n624 VDD.n621 185
R12280 VDD.n1784 VDD.n1783 185
R12281 VDD.n1783 VDD.n1782 185
R12282 VDD.n626 VDD.n625 185
R12283 VDD.n627 VDD.n626 185
R12284 VDD.n1776 VDD.n1775 185
R12285 VDD.t16 VDD.n1776 185
R12286 VDD.n1774 VDD.n636 185
R12287 VDD.n636 VDD.n633 185
R12288 VDD.n1773 VDD.n1772 185
R12289 VDD.n1772 VDD.n1771 185
R12290 VDD.n638 VDD.n637 185
R12291 VDD.n639 VDD.n638 185
R12292 VDD.n1764 VDD.n1763 185
R12293 VDD.n1765 VDD.n1764 185
R12294 VDD.n1762 VDD.n647 185
R12295 VDD.n647 VDD.t17 185
R12296 VDD.n1761 VDD.n1760 185
R12297 VDD.n1760 VDD.n1759 185
R12298 VDD.n649 VDD.n648 185
R12299 VDD.n650 VDD.n649 185
R12300 VDD.n1752 VDD.n1751 185
R12301 VDD.n1753 VDD.n1752 185
R12302 VDD.n1750 VDD.n659 185
R12303 VDD.n659 VDD.n656 185
R12304 VDD.n1749 VDD.n1748 185
R12305 VDD.n1748 VDD.n1747 185
R12306 VDD.n661 VDD.n660 185
R12307 VDD.n662 VDD.n661 185
R12308 VDD.n1740 VDD.n1739 185
R12309 VDD.n1741 VDD.n1740 185
R12310 VDD.n1738 VDD.n671 185
R12311 VDD.n671 VDD.n668 185
R12312 VDD.n1737 VDD.n1736 185
R12313 VDD.n1736 VDD.n1735 185
R12314 VDD.n673 VDD.n672 185
R12315 VDD.n674 VDD.n673 185
R12316 VDD.n1728 VDD.n1727 185
R12317 VDD.n1729 VDD.n1728 185
R12318 VDD.n1726 VDD.n682 185
R12319 VDD.n688 VDD.n682 185
R12320 VDD.n1725 VDD.n1724 185
R12321 VDD.n1724 VDD.n1723 185
R12322 VDD.n684 VDD.n683 185
R12323 VDD.n685 VDD.n684 185
R12324 VDD.n1716 VDD.n1715 185
R12325 VDD.n1717 VDD.n1716 185
R12326 VDD.n1714 VDD.n695 185
R12327 VDD.n695 VDD.n692 185
R12328 VDD.n1713 VDD.n1712 185
R12329 VDD.n1712 VDD.n1711 185
R12330 VDD.n697 VDD.n696 185
R12331 VDD.n698 VDD.n697 185
R12332 VDD.n1703 VDD.n1702 185
R12333 VDD.n1701 VDD.n720 185
R12334 VDD.n1700 VDD.n719 185
R12335 VDD.n1705 VDD.n719 185
R12336 VDD.n1699 VDD.n1698 185
R12337 VDD.n1697 VDD.n1696 185
R12338 VDD.n1695 VDD.n1694 185
R12339 VDD.n1693 VDD.n1692 185
R12340 VDD.n1691 VDD.n1690 185
R12341 VDD.n1688 VDD.n1687 185
R12342 VDD.n1686 VDD.n1685 185
R12343 VDD.n1684 VDD.n1683 185
R12344 VDD.n1682 VDD.n1681 185
R12345 VDD.n1679 VDD.n1678 185
R12346 VDD.n1677 VDD.n1676 185
R12347 VDD.n1675 VDD.n1674 185
R12348 VDD.n1673 VDD.n710 185
R12349 VDD.n1705 VDD.n710 185
R12350 VDD.n1849 VDD.n1848 185
R12351 VDD.n1851 VDD.n1850 185
R12352 VDD.n1853 VDD.n1852 185
R12353 VDD.n1855 VDD.n1854 185
R12354 VDD.n1857 VDD.n1856 185
R12355 VDD.n1859 VDD.n1858 185
R12356 VDD.n1861 VDD.n1860 185
R12357 VDD.n1863 VDD.n1862 185
R12358 VDD.n1865 VDD.n1864 185
R12359 VDD.n1867 VDD.n1866 185
R12360 VDD.n1869 VDD.n1868 185
R12361 VDD.n1871 VDD.n1870 185
R12362 VDD.n1873 VDD.n1872 185
R12363 VDD.n1875 VDD.n1874 185
R12364 VDD.n1877 VDD.n1876 185
R12365 VDD.n1879 VDD.n1878 185
R12366 VDD.n1847 VDD.n1846 185
R12367 VDD.n1847 VDD.n537 185
R12368 VDD.n1845 VDD.n562 185
R12369 VDD.n1883 VDD.n562 185
R12370 VDD.n1844 VDD.n1843 185
R12371 VDD.n1843 VDD.n561 185
R12372 VDD.n1842 VDD.n570 185
R12373 VDD.n1842 VDD.n1841 185
R12374 VDD.n1609 VDD.n571 185
R12375 VDD.n572 VDD.n571 185
R12376 VDD.n1610 VDD.n578 185
R12377 VDD.n1835 VDD.n578 185
R12378 VDD.n1612 VDD.n1611 185
R12379 VDD.n1611 VDD.n586 185
R12380 VDD.n1613 VDD.n584 185
R12381 VDD.n1824 VDD.n584 185
R12382 VDD.n1615 VDD.n1614 185
R12383 VDD.n1614 VDD.n593 185
R12384 VDD.n1616 VDD.n591 185
R12385 VDD.n1818 VDD.n591 185
R12386 VDD.n1618 VDD.n1617 185
R12387 VDD.n1617 VDD.n590 185
R12388 VDD.n1619 VDD.n598 185
R12389 VDD.n1812 VDD.n598 185
R12390 VDD.n1621 VDD.n1620 185
R12391 VDD.n1620 VDD.n597 185
R12392 VDD.n1622 VDD.n604 185
R12393 VDD.n1806 VDD.n604 185
R12394 VDD.n1624 VDD.n1623 185
R12395 VDD.n1623 VDD.n603 185
R12396 VDD.n1625 VDD.n610 185
R12397 VDD.n1800 VDD.n610 185
R12398 VDD.n1627 VDD.n1626 185
R12399 VDD.n1626 VDD.n609 185
R12400 VDD.n1628 VDD.n616 185
R12401 VDD.n1794 VDD.n616 185
R12402 VDD.n1630 VDD.n1629 185
R12403 VDD.n1629 VDD.n615 185
R12404 VDD.n1631 VDD.n622 185
R12405 VDD.n1788 VDD.n622 185
R12406 VDD.n1633 VDD.n1632 185
R12407 VDD.n1632 VDD.n621 185
R12408 VDD.n1634 VDD.n628 185
R12409 VDD.n1782 VDD.n628 185
R12410 VDD.n1636 VDD.n1635 185
R12411 VDD.n1635 VDD.n627 185
R12412 VDD.n1637 VDD.n635 185
R12413 VDD.t16 VDD.n635 185
R12414 VDD.n1639 VDD.n1638 185
R12415 VDD.n1638 VDD.n633 185
R12416 VDD.n1640 VDD.n640 185
R12417 VDD.n1771 VDD.n640 185
R12418 VDD.n1642 VDD.n1641 185
R12419 VDD.n1641 VDD.n639 185
R12420 VDD.n1643 VDD.n645 185
R12421 VDD.n1765 VDD.n645 185
R12422 VDD.n1645 VDD.n1644 185
R12423 VDD.n1644 VDD.t17 185
R12424 VDD.n1646 VDD.n651 185
R12425 VDD.n1759 VDD.n651 185
R12426 VDD.n1648 VDD.n1647 185
R12427 VDD.n1647 VDD.n650 185
R12428 VDD.n1649 VDD.n657 185
R12429 VDD.n1753 VDD.n657 185
R12430 VDD.n1651 VDD.n1650 185
R12431 VDD.n1650 VDD.n656 185
R12432 VDD.n1652 VDD.n663 185
R12433 VDD.n1747 VDD.n663 185
R12434 VDD.n1654 VDD.n1653 185
R12435 VDD.n1653 VDD.n662 185
R12436 VDD.n1655 VDD.n669 185
R12437 VDD.n1741 VDD.n669 185
R12438 VDD.n1657 VDD.n1656 185
R12439 VDD.n1656 VDD.n668 185
R12440 VDD.n1658 VDD.n675 185
R12441 VDD.n1735 VDD.n675 185
R12442 VDD.n1660 VDD.n1659 185
R12443 VDD.n1659 VDD.n674 185
R12444 VDD.n1661 VDD.n680 185
R12445 VDD.n1729 VDD.n680 185
R12446 VDD.n1663 VDD.n1662 185
R12447 VDD.n1662 VDD.n688 185
R12448 VDD.n1664 VDD.n686 185
R12449 VDD.n1723 VDD.n686 185
R12450 VDD.n1666 VDD.n1665 185
R12451 VDD.n1665 VDD.n685 185
R12452 VDD.n1667 VDD.n693 185
R12453 VDD.n1717 VDD.n693 185
R12454 VDD.n1669 VDD.n1668 185
R12455 VDD.n1668 VDD.n692 185
R12456 VDD.n1670 VDD.n699 185
R12457 VDD.n1711 VDD.n699 185
R12458 VDD.n1672 VDD.n1671 185
R12459 VDD.n1671 VDD.n698 185
R12460 VDD.n2323 VDD.n387 185
R12461 VDD.n387 VDD.n384 185
R12462 VDD.n2325 VDD.n2324 185
R12463 VDD.n2326 VDD.n2325 185
R12464 VDD.n388 VDD.n386 185
R12465 VDD.n386 VDD.n382 185
R12466 VDD.n2285 VDD.n2284 185
R12467 VDD.n2286 VDD.n2285 185
R12468 VDD.n2283 VDD.n408 185
R12469 VDD.n408 VDD.n405 185
R12470 VDD.n2282 VDD.n2281 185
R12471 VDD.n2281 VDD.n2280 185
R12472 VDD.n410 VDD.n409 185
R12473 VDD.n411 VDD.n410 185
R12474 VDD.n2248 VDD.n2247 185
R12475 VDD.n2249 VDD.n2248 185
R12476 VDD.n2246 VDD.n420 185
R12477 VDD.n426 VDD.n420 185
R12478 VDD.n2245 VDD.n2244 185
R12479 VDD.n2244 VDD.n2243 185
R12480 VDD.n422 VDD.n421 185
R12481 VDD.n423 VDD.n422 185
R12482 VDD.n2236 VDD.n2235 185
R12483 VDD.n2237 VDD.n2236 185
R12484 VDD.n2234 VDD.n433 185
R12485 VDD.n433 VDD.n430 185
R12486 VDD.n2233 VDD.n2232 185
R12487 VDD.n2232 VDD.n2231 185
R12488 VDD.n435 VDD.n434 185
R12489 VDD.n436 VDD.n435 185
R12490 VDD.n2224 VDD.n2223 185
R12491 VDD.n2225 VDD.n2224 185
R12492 VDD.n2222 VDD.n445 185
R12493 VDD.n445 VDD.n442 185
R12494 VDD.n2221 VDD.n2220 185
R12495 VDD.n2220 VDD.n2219 185
R12496 VDD.n447 VDD.n446 185
R12497 VDD.t19 VDD.n447 185
R12498 VDD.n2212 VDD.n2211 185
R12499 VDD.n2213 VDD.n2212 185
R12500 VDD.n2210 VDD.n456 185
R12501 VDD.n456 VDD.n453 185
R12502 VDD.n2209 VDD.n2208 185
R12503 VDD.n2208 VDD.n2207 185
R12504 VDD.n458 VDD.n457 185
R12505 VDD.n459 VDD.n458 185
R12506 VDD.n2201 VDD.n2200 185
R12507 VDD.t23 VDD.n2201 185
R12508 VDD.n2199 VDD.n468 185
R12509 VDD.n468 VDD.n465 185
R12510 VDD.n2198 VDD.n2197 185
R12511 VDD.n2197 VDD.n2196 185
R12512 VDD.n470 VDD.n469 185
R12513 VDD.n471 VDD.n470 185
R12514 VDD.n2189 VDD.n2188 185
R12515 VDD.n2190 VDD.n2189 185
R12516 VDD.n2187 VDD.n480 185
R12517 VDD.n480 VDD.n477 185
R12518 VDD.n2186 VDD.n2185 185
R12519 VDD.n2185 VDD.n2184 185
R12520 VDD.n482 VDD.n481 185
R12521 VDD.n491 VDD.n482 185
R12522 VDD.n2177 VDD.n2176 185
R12523 VDD.n2178 VDD.n2177 185
R12524 VDD.n2175 VDD.n492 185
R12525 VDD.n492 VDD.n488 185
R12526 VDD.n2174 VDD.n2173 185
R12527 VDD.n2173 VDD.n2172 185
R12528 VDD.n494 VDD.n493 185
R12529 VDD.n495 VDD.n494 185
R12530 VDD.n2165 VDD.n2164 185
R12531 VDD.n2166 VDD.n2165 185
R12532 VDD.n2163 VDD.n504 185
R12533 VDD.n504 VDD.n501 185
R12534 VDD.n2162 VDD.n2161 185
R12535 VDD.n2161 VDD.n2160 185
R12536 VDD.n506 VDD.n505 185
R12537 VDD.n507 VDD.n506 185
R12538 VDD.n2153 VDD.n2152 185
R12539 VDD.n2154 VDD.n2153 185
R12540 VDD.n2151 VDD.n516 185
R12541 VDD.n516 VDD.n513 185
R12542 VDD.n2150 VDD.n2149 185
R12543 VDD.n2149 VDD.n2148 185
R12544 VDD.n518 VDD.n517 185
R12545 VDD.n519 VDD.n518 185
R12546 VDD.n2141 VDD.n2140 185
R12547 VDD.n2142 VDD.n2141 185
R12548 VDD.n2139 VDD.n528 185
R12549 VDD.n528 VDD.n525 185
R12550 VDD.n2138 VDD.n2137 185
R12551 VDD.n2137 VDD.n2136 185
R12552 VDD.n530 VDD.n529 185
R12553 VDD.n531 VDD.n530 185
R12554 VDD.n2127 VDD.n2126 185
R12555 VDD.n2125 VDD.n2031 185
R12556 VDD.n2124 VDD.n2030 185
R12557 VDD.n2129 VDD.n2030 185
R12558 VDD.n2123 VDD.n2122 185
R12559 VDD.n2121 VDD.n2120 185
R12560 VDD.n2119 VDD.n2118 185
R12561 VDD.n2117 VDD.n2116 185
R12562 VDD.n2115 VDD.n2114 185
R12563 VDD.n2113 VDD.n2112 185
R12564 VDD.n2111 VDD.n2110 185
R12565 VDD.n2109 VDD.n2108 185
R12566 VDD.n2107 VDD.n2106 185
R12567 VDD.n2104 VDD.n2103 185
R12568 VDD.n2102 VDD.n2101 185
R12569 VDD.n2100 VDD.n2099 185
R12570 VDD.n2098 VDD.n1925 185
R12571 VDD.n2129 VDD.n1925 185
R12572 VDD.n2293 VDD.n2292 185
R12573 VDD.n2295 VDD.n400 185
R12574 VDD.n2297 VDD.n2296 185
R12575 VDD.n2298 VDD.n397 185
R12576 VDD.n2301 VDD.n2300 185
R12577 VDD.n2303 VDD.n395 185
R12578 VDD.n2305 VDD.n2304 185
R12579 VDD.n2306 VDD.n394 185
R12580 VDD.n2309 VDD.n2308 185
R12581 VDD.n2311 VDD.n392 185
R12582 VDD.n2313 VDD.n2312 185
R12583 VDD.n2314 VDD.n391 185
R12584 VDD.n2316 VDD.n2315 185
R12585 VDD.n2318 VDD.n390 185
R12586 VDD.n2319 VDD.n389 185
R12587 VDD.n2322 VDD.n2321 185
R12588 VDD.n2291 VDD.n402 185
R12589 VDD.n402 VDD.n384 185
R12590 VDD.n2290 VDD.n383 185
R12591 VDD.n2326 VDD.n383 185
R12592 VDD.n2289 VDD.n2288 185
R12593 VDD.n2288 VDD.n382 185
R12594 VDD.n2287 VDD.n403 185
R12595 VDD.n2287 VDD.n2286 185
R12596 VDD.n2034 VDD.n404 185
R12597 VDD.n405 VDD.n404 185
R12598 VDD.n2035 VDD.n412 185
R12599 VDD.n2280 VDD.n412 185
R12600 VDD.n2037 VDD.n2036 185
R12601 VDD.n2036 VDD.n411 185
R12602 VDD.n2038 VDD.n418 185
R12603 VDD.n2249 VDD.n418 185
R12604 VDD.n2040 VDD.n2039 185
R12605 VDD.n2039 VDD.n426 185
R12606 VDD.n2041 VDD.n424 185
R12607 VDD.n2243 VDD.n424 185
R12608 VDD.n2043 VDD.n2042 185
R12609 VDD.n2042 VDD.n423 185
R12610 VDD.n2044 VDD.n431 185
R12611 VDD.n2237 VDD.n431 185
R12612 VDD.n2046 VDD.n2045 185
R12613 VDD.n2045 VDD.n430 185
R12614 VDD.n2047 VDD.n437 185
R12615 VDD.n2231 VDD.n437 185
R12616 VDD.n2049 VDD.n2048 185
R12617 VDD.n2048 VDD.n436 185
R12618 VDD.n2050 VDD.n443 185
R12619 VDD.n2225 VDD.n443 185
R12620 VDD.n2052 VDD.n2051 185
R12621 VDD.n2051 VDD.n442 185
R12622 VDD.n2053 VDD.n448 185
R12623 VDD.n2219 VDD.n448 185
R12624 VDD.n2055 VDD.n2054 185
R12625 VDD.n2054 VDD.t19 185
R12626 VDD.n2056 VDD.n454 185
R12627 VDD.n2213 VDD.n454 185
R12628 VDD.n2058 VDD.n2057 185
R12629 VDD.n2057 VDD.n453 185
R12630 VDD.n2059 VDD.n460 185
R12631 VDD.n2207 VDD.n460 185
R12632 VDD.n2061 VDD.n2060 185
R12633 VDD.n2060 VDD.n459 185
R12634 VDD.n2062 VDD.n467 185
R12635 VDD.t23 VDD.n467 185
R12636 VDD.n2064 VDD.n2063 185
R12637 VDD.n2063 VDD.n465 185
R12638 VDD.n2065 VDD.n472 185
R12639 VDD.n2196 VDD.n472 185
R12640 VDD.n2067 VDD.n2066 185
R12641 VDD.n2066 VDD.n471 185
R12642 VDD.n2068 VDD.n478 185
R12643 VDD.n2190 VDD.n478 185
R12644 VDD.n2070 VDD.n2069 185
R12645 VDD.n2069 VDD.n477 185
R12646 VDD.n2071 VDD.n483 185
R12647 VDD.n2184 VDD.n483 185
R12648 VDD.n2073 VDD.n2072 185
R12649 VDD.n2072 VDD.n491 185
R12650 VDD.n2074 VDD.n489 185
R12651 VDD.n2178 VDD.n489 185
R12652 VDD.n2076 VDD.n2075 185
R12653 VDD.n2075 VDD.n488 185
R12654 VDD.n2077 VDD.n496 185
R12655 VDD.n2172 VDD.n496 185
R12656 VDD.n2079 VDD.n2078 185
R12657 VDD.n2078 VDD.n495 185
R12658 VDD.n2080 VDD.n502 185
R12659 VDD.n2166 VDD.n502 185
R12660 VDD.n2082 VDD.n2081 185
R12661 VDD.n2081 VDD.n501 185
R12662 VDD.n2083 VDD.n508 185
R12663 VDD.n2160 VDD.n508 185
R12664 VDD.n2085 VDD.n2084 185
R12665 VDD.n2084 VDD.n507 185
R12666 VDD.n2086 VDD.n514 185
R12667 VDD.n2154 VDD.n514 185
R12668 VDD.n2088 VDD.n2087 185
R12669 VDD.n2087 VDD.n513 185
R12670 VDD.n2089 VDD.n520 185
R12671 VDD.n2148 VDD.n520 185
R12672 VDD.n2091 VDD.n2090 185
R12673 VDD.n2090 VDD.n519 185
R12674 VDD.n2092 VDD.n526 185
R12675 VDD.n2142 VDD.n526 185
R12676 VDD.n2094 VDD.n2093 185
R12677 VDD.n2093 VDD.n525 185
R12678 VDD.n2095 VDD.n532 185
R12679 VDD.n2136 VDD.n532 185
R12680 VDD.n2097 VDD.n2096 185
R12681 VDD.n2096 VDD.n531 185
R12682 VDD.n1523 VDD.n1522 185
R12683 VDD.n1524 VDD.n1523 185
R12684 VDD.n918 VDD.n916 185
R12685 VDD.n916 VDD.n915 185
R12686 VDD.n1491 VDD.n1490 185
R12687 VDD.n1490 VDD.n1489 185
R12688 VDD.n921 VDD.n920 185
R12689 VDD.n922 VDD.n921 185
R12690 VDD.n1479 VDD.n1478 185
R12691 VDD.n1480 VDD.n1479 185
R12692 VDD.n931 VDD.n930 185
R12693 VDD.n930 VDD.n929 185
R12694 VDD.n1474 VDD.n1473 185
R12695 VDD.n1473 VDD.n1472 185
R12696 VDD.n934 VDD.n933 185
R12697 VDD.n935 VDD.n934 185
R12698 VDD.n1463 VDD.n1462 185
R12699 VDD.n1464 VDD.n1463 185
R12700 VDD.n943 VDD.n942 185
R12701 VDD.n942 VDD.n941 185
R12702 VDD.n1458 VDD.n1457 185
R12703 VDD.n1457 VDD.n1456 185
R12704 VDD.n946 VDD.n945 185
R12705 VDD.n947 VDD.n946 185
R12706 VDD.n1447 VDD.n1446 185
R12707 VDD.n1448 VDD.n1447 185
R12708 VDD.n955 VDD.n954 185
R12709 VDD.n954 VDD.n953 185
R12710 VDD.n1442 VDD.n1441 185
R12711 VDD.n1441 VDD.n1440 185
R12712 VDD.n958 VDD.n957 185
R12713 VDD.n959 VDD.n958 185
R12714 VDD.n1431 VDD.n1430 185
R12715 VDD.n1432 VDD.n1431 185
R12716 VDD.n967 VDD.n966 185
R12717 VDD.n966 VDD.n965 185
R12718 VDD.n1426 VDD.n1425 185
R12719 VDD.n1425 VDD.n1424 185
R12720 VDD.n970 VDD.n969 185
R12721 VDD.n971 VDD.n970 185
R12722 VDD.n1415 VDD.n1414 185
R12723 VDD.n1416 VDD.n1415 185
R12724 VDD.n979 VDD.n978 185
R12725 VDD.n978 VDD.n977 185
R12726 VDD.n1410 VDD.n1409 185
R12727 VDD.n1409 VDD.n1408 185
R12728 VDD.n982 VDD.n981 185
R12729 VDD.n983 VDD.n982 185
R12730 VDD.n1399 VDD.n1398 185
R12731 VDD.n1400 VDD.n1399 185
R12732 VDD.n991 VDD.n990 185
R12733 VDD.n990 VDD.n989 185
R12734 VDD.n1382 VDD.n1381 185
R12735 VDD.n1381 VDD.t12 185
R12736 VDD.n994 VDD.n993 185
R12737 VDD.n995 VDD.n994 185
R12738 VDD.n1372 VDD.n1371 185
R12739 VDD.n1373 VDD.n1372 185
R12740 VDD.n1003 VDD.n1002 185
R12741 VDD.n1002 VDD.n1001 185
R12742 VDD.n1367 VDD.n1366 185
R12743 VDD.n1366 VDD.n1365 185
R12744 VDD.n1006 VDD.n1005 185
R12745 VDD.n1007 VDD.n1006 185
R12746 VDD.n1356 VDD.n1355 185
R12747 VDD.n1357 VDD.n1356 185
R12748 VDD.n1015 VDD.n1014 185
R12749 VDD.n1014 VDD.n1013 185
R12750 VDD.n1351 VDD.n1350 185
R12751 VDD.n1350 VDD.n1349 185
R12752 VDD.n1018 VDD.n1017 185
R12753 VDD.n1025 VDD.n1018 185
R12754 VDD.n1340 VDD.n1339 185
R12755 VDD.n1341 VDD.n1340 185
R12756 VDD.n1027 VDD.n1026 185
R12757 VDD.n1026 VDD.n1024 185
R12758 VDD.n1335 VDD.n1334 185
R12759 VDD.n1334 VDD.n1333 185
R12760 VDD.n1030 VDD.n1029 185
R12761 VDD.n1031 VDD.n1030 185
R12762 VDD.n1324 VDD.n1323 185
R12763 VDD.n1325 VDD.n1324 185
R12764 VDD.n1039 VDD.n1038 185
R12765 VDD.n1038 VDD.n1037 185
R12766 VDD.n1319 VDD.n1318 185
R12767 VDD.n1318 VDD.n1317 185
R12768 VDD.n1042 VDD.n1041 185
R12769 VDD.n1043 VDD.n1042 185
R12770 VDD.n1308 VDD.n1307 185
R12771 VDD.n1309 VDD.n1308 185
R12772 VDD.n1051 VDD.n1050 185
R12773 VDD.n1050 VDD.n1049 185
R12774 VDD.n1303 VDD.n1302 185
R12775 VDD.n1302 VDD.n1301 185
R12776 VDD.n1054 VDD.n1053 185
R12777 VDD.n1061 VDD.n1054 185
R12778 VDD.n1292 VDD.n1291 185
R12779 VDD.n1293 VDD.n1292 185
R12780 VDD.n1063 VDD.n1062 185
R12781 VDD.n1062 VDD.n1060 185
R12782 VDD.n1287 VDD.n1286 185
R12783 VDD.n1286 VDD.n1285 185
R12784 VDD.n1066 VDD.n1065 185
R12785 VDD.n1067 VDD.n1066 185
R12786 VDD.n1276 VDD.n1275 185
R12787 VDD.n1277 VDD.n1276 185
R12788 VDD.n1272 VDD.n1073 185
R12789 VDD.n1271 VDD.n1076 185
R12790 VDD.n1270 VDD.n1077 185
R12791 VDD.n1077 VDD.n1072 185
R12792 VDD.n1080 VDD.n1078 185
R12793 VDD.n1266 VDD.n1082 185
R12794 VDD.n1265 VDD.n1083 185
R12795 VDD.n1264 VDD.n1085 185
R12796 VDD.n1088 VDD.n1086 185
R12797 VDD.n1260 VDD.n1090 185
R12798 VDD.n1259 VDD.n1091 185
R12799 VDD.n1258 VDD.n1093 185
R12800 VDD.n1098 VDD.n1096 185
R12801 VDD.n1254 VDD.n1100 185
R12802 VDD.n1253 VDD.n1101 185
R12803 VDD.n1252 VDD.n1103 185
R12804 VDD.n1106 VDD.n1104 185
R12805 VDD.n1248 VDD.n1108 185
R12806 VDD.n1247 VDD.n1109 185
R12807 VDD.n1246 VDD.n1111 185
R12808 VDD.n1114 VDD.n1112 185
R12809 VDD.n1242 VDD.n1116 185
R12810 VDD.n1241 VDD.n1117 185
R12811 VDD.n1240 VDD.n1119 185
R12812 VDD.n1122 VDD.n1120 185
R12813 VDD.n1236 VDD.n1124 185
R12814 VDD.n1235 VDD.n1125 185
R12815 VDD.n1231 VDD.n1127 185
R12816 VDD.n1130 VDD.n1128 185
R12817 VDD.n1227 VDD.n1132 185
R12818 VDD.n1226 VDD.n1133 185
R12819 VDD.n1225 VDD.n1135 185
R12820 VDD.n1138 VDD.n1136 185
R12821 VDD.n1221 VDD.n1140 185
R12822 VDD.n1220 VDD.n1141 185
R12823 VDD.n1219 VDD.n1143 185
R12824 VDD.n1146 VDD.n1144 185
R12825 VDD.n1215 VDD.n1148 185
R12826 VDD.n1214 VDD.n1149 185
R12827 VDD.n1213 VDD.n1151 185
R12828 VDD.n1157 VDD.n1152 185
R12829 VDD.n1209 VDD.n1159 185
R12830 VDD.n1208 VDD.n1160 185
R12831 VDD.n1207 VDD.n1162 185
R12832 VDD.n1165 VDD.n1163 185
R12833 VDD.n1203 VDD.n1167 185
R12834 VDD.n1202 VDD.n1168 185
R12835 VDD.n1201 VDD.n1170 185
R12836 VDD.n1173 VDD.n1171 185
R12837 VDD.n1197 VDD.n1175 185
R12838 VDD.n1196 VDD.n1176 185
R12839 VDD.n1195 VDD.n1178 185
R12840 VDD.n1181 VDD.n1179 185
R12841 VDD.n1191 VDD.n1183 185
R12842 VDD.n1190 VDD.n1185 185
R12843 VDD.n1186 VDD.n1071 185
R12844 VDD.n1527 VDD.n1526 185
R12845 VDD.n911 VDD.n906 185
R12846 VDD.n1531 VDD.n905 185
R12847 VDD.n1532 VDD.n903 185
R12848 VDD.n1533 VDD.n902 185
R12849 VDD.n900 VDD.n898 185
R12850 VDD.n1537 VDD.n897 185
R12851 VDD.n1538 VDD.n895 185
R12852 VDD.n1539 VDD.n894 185
R12853 VDD.n892 VDD.n887 185
R12854 VDD.n891 VDD.n890 185
R12855 VDD.n888 VDD.n786 185
R12856 VDD.n1543 VDD.n785 185
R12857 VDD.n1544 VDD.n777 185
R12858 VDD.n1546 VDD.n1545 185
R12859 VDD.n1548 VDD.n775 185
R12860 VDD.n1550 VDD.n1549 185
R12861 VDD.n1551 VDD.n770 185
R12862 VDD.n1553 VDD.n1552 185
R12863 VDD.n1555 VDD.n768 185
R12864 VDD.n1557 VDD.n1556 185
R12865 VDD.n1558 VDD.n763 185
R12866 VDD.n1560 VDD.n1559 185
R12867 VDD.n1562 VDD.n761 185
R12868 VDD.n1564 VDD.n1563 185
R12869 VDD.n1565 VDD.n756 185
R12870 VDD.n1567 VDD.n1566 185
R12871 VDD.n1569 VDD.n754 185
R12872 VDD.n1571 VDD.n1570 185
R12873 VDD.n1575 VDD.n749 185
R12874 VDD.n1577 VDD.n1576 185
R12875 VDD.n1579 VDD.n747 185
R12876 VDD.n1581 VDD.n1580 185
R12877 VDD.n1582 VDD.n742 185
R12878 VDD.n1584 VDD.n1583 185
R12879 VDD.n1586 VDD.n740 185
R12880 VDD.n1588 VDD.n1587 185
R12881 VDD.n1589 VDD.n735 185
R12882 VDD.n1591 VDD.n1590 185
R12883 VDD.n1593 VDD.n733 185
R12884 VDD.n1595 VDD.n1594 185
R12885 VDD.n1596 VDD.n731 185
R12886 VDD.n1598 VDD.n1597 185
R12887 VDD.n1600 VDD.n730 185
R12888 VDD.n1601 VDD.n724 185
R12889 VDD.n1604 VDD.n1603 185
R12890 VDD.n726 VDD.n725 185
R12891 VDD.n1507 VDD.n1504 185
R12892 VDD.n1509 VDD.n1508 185
R12893 VDD.n1510 VDD.n1497 185
R12894 VDD.n1512 VDD.n1511 185
R12895 VDD.n1514 VDD.n1496 185
R12896 VDD.n1515 VDD.n1495 185
R12897 VDD.n1518 VDD.n1517 185
R12898 VDD.n1519 VDD.n917 185
R12899 VDD.n917 VDD.n727 185
R12900 VDD.n1525 VDD.n914 185
R12901 VDD.n1525 VDD.n1524 185
R12902 VDD.n925 VDD.n913 185
R12903 VDD.n915 VDD.n913 185
R12904 VDD.n1488 VDD.n1487 185
R12905 VDD.n1489 VDD.n1488 185
R12906 VDD.n924 VDD.n923 185
R12907 VDD.n923 VDD.n922 185
R12908 VDD.n1482 VDD.n1481 185
R12909 VDD.n1481 VDD.n1480 185
R12910 VDD.n928 VDD.n927 185
R12911 VDD.n929 VDD.n928 185
R12912 VDD.n1471 VDD.n1470 185
R12913 VDD.n1472 VDD.n1471 185
R12914 VDD.n937 VDD.n936 185
R12915 VDD.n936 VDD.n935 185
R12916 VDD.n1466 VDD.n1465 185
R12917 VDD.n1465 VDD.n1464 185
R12918 VDD.n940 VDD.n939 185
R12919 VDD.n941 VDD.n940 185
R12920 VDD.n1455 VDD.n1454 185
R12921 VDD.n1456 VDD.n1455 185
R12922 VDD.n949 VDD.n948 185
R12923 VDD.n948 VDD.n947 185
R12924 VDD.n1450 VDD.n1449 185
R12925 VDD.n1449 VDD.n1448 185
R12926 VDD.n952 VDD.n951 185
R12927 VDD.n953 VDD.n952 185
R12928 VDD.n1439 VDD.n1438 185
R12929 VDD.n1440 VDD.n1439 185
R12930 VDD.n961 VDD.n960 185
R12931 VDD.n960 VDD.n959 185
R12932 VDD.n1434 VDD.n1433 185
R12933 VDD.n1433 VDD.n1432 185
R12934 VDD.n964 VDD.n963 185
R12935 VDD.n965 VDD.n964 185
R12936 VDD.n1423 VDD.n1422 185
R12937 VDD.n1424 VDD.n1423 185
R12938 VDD.n973 VDD.n972 185
R12939 VDD.n972 VDD.n971 185
R12940 VDD.n1418 VDD.n1417 185
R12941 VDD.n1417 VDD.n1416 185
R12942 VDD.n976 VDD.n975 185
R12943 VDD.n977 VDD.n976 185
R12944 VDD.n1407 VDD.n1406 185
R12945 VDD.n1408 VDD.n1407 185
R12946 VDD.n985 VDD.n984 185
R12947 VDD.n984 VDD.n983 185
R12948 VDD.n1402 VDD.n1401 185
R12949 VDD.n1401 VDD.n1400 185
R12950 VDD.n988 VDD.n987 185
R12951 VDD.n989 VDD.n988 185
R12952 VDD.n1380 VDD.n1379 185
R12953 VDD.t12 VDD.n1380 185
R12954 VDD.n997 VDD.n996 185
R12955 VDD.n996 VDD.n995 185
R12956 VDD.n1375 VDD.n1374 185
R12957 VDD.n1374 VDD.n1373 185
R12958 VDD.n1000 VDD.n999 185
R12959 VDD.n1001 VDD.n1000 185
R12960 VDD.n1364 VDD.n1363 185
R12961 VDD.n1365 VDD.n1364 185
R12962 VDD.n1009 VDD.n1008 185
R12963 VDD.n1008 VDD.n1007 185
R12964 VDD.n1359 VDD.n1358 185
R12965 VDD.n1358 VDD.n1357 185
R12966 VDD.n1012 VDD.n1011 185
R12967 VDD.n1013 VDD.n1012 185
R12968 VDD.n1348 VDD.n1347 185
R12969 VDD.n1349 VDD.n1348 185
R12970 VDD.n1020 VDD.n1019 185
R12971 VDD.n1025 VDD.n1019 185
R12972 VDD.n1343 VDD.n1342 185
R12973 VDD.n1342 VDD.n1341 185
R12974 VDD.n1023 VDD.n1022 185
R12975 VDD.n1024 VDD.n1023 185
R12976 VDD.n1332 VDD.n1331 185
R12977 VDD.n1333 VDD.n1332 185
R12978 VDD.n1033 VDD.n1032 185
R12979 VDD.n1032 VDD.n1031 185
R12980 VDD.n1327 VDD.n1326 185
R12981 VDD.n1326 VDD.n1325 185
R12982 VDD.n1036 VDD.n1035 185
R12983 VDD.n1037 VDD.n1036 185
R12984 VDD.n1316 VDD.n1315 185
R12985 VDD.n1317 VDD.n1316 185
R12986 VDD.n1045 VDD.n1044 185
R12987 VDD.n1044 VDD.n1043 185
R12988 VDD.n1311 VDD.n1310 185
R12989 VDD.n1310 VDD.n1309 185
R12990 VDD.n1048 VDD.n1047 185
R12991 VDD.n1049 VDD.n1048 185
R12992 VDD.n1300 VDD.n1299 185
R12993 VDD.n1301 VDD.n1300 185
R12994 VDD.n1056 VDD.n1055 185
R12995 VDD.n1061 VDD.n1055 185
R12996 VDD.n1295 VDD.n1294 185
R12997 VDD.n1294 VDD.n1293 185
R12998 VDD.n1059 VDD.n1058 185
R12999 VDD.n1060 VDD.n1059 185
R13000 VDD.n1284 VDD.n1283 185
R13001 VDD.n1285 VDD.n1284 185
R13002 VDD.n1069 VDD.n1068 185
R13003 VDD.n1068 VDD.n1067 185
R13004 VDD.n1279 VDD.n1278 185
R13005 VDD.n1278 VDD.n1277 185
R13006 VDD.n2473 VDD.n299 185
R13007 VDD.n2472 VDD.n2471 185
R13008 VDD.n2469 VDD.n301 185
R13009 VDD.n2469 VDD.n298 185
R13010 VDD.n2468 VDD.n2467 185
R13011 VDD.n2466 VDD.n2465 185
R13012 VDD.n2464 VDD.n306 185
R13013 VDD.n2462 VDD.n2461 185
R13014 VDD.n2460 VDD.n307 185
R13015 VDD.n2459 VDD.n2458 185
R13016 VDD.n2456 VDD.n312 185
R13017 VDD.n2454 VDD.n2453 185
R13018 VDD.n2451 VDD.n313 185
R13019 VDD.n2450 VDD.n318 185
R13020 VDD.n2449 VDD.n2448 185
R13021 VDD.n2446 VDD.n320 185
R13022 VDD.n2445 VDD.n2444 185
R13023 VDD.n2443 VDD.n2442 185
R13024 VDD.n2441 VDD.n325 185
R13025 VDD.n2439 VDD.n2438 185
R13026 VDD.n2437 VDD.n326 185
R13027 VDD.n2436 VDD.n2435 185
R13028 VDD.n2433 VDD.n331 185
R13029 VDD.n2431 VDD.n2430 185
R13030 VDD.n2429 VDD.n332 185
R13031 VDD.n2428 VDD.n2427 185
R13032 VDD.n2425 VDD.n337 185
R13033 VDD.n2423 VDD.n2422 185
R13034 VDD.n2421 VDD.n338 185
R13035 VDD.n2420 VDD.n2419 185
R13036 VDD.n2417 VDD.n346 185
R13037 VDD.n2415 VDD.n2414 185
R13038 VDD.n2413 VDD.n347 185
R13039 VDD.n2412 VDD.n2411 185
R13040 VDD.n2409 VDD.n352 185
R13041 VDD.n2407 VDD.n2406 185
R13042 VDD.n2405 VDD.n353 185
R13043 VDD.n2404 VDD.n2403 185
R13044 VDD.n2401 VDD.n358 185
R13045 VDD.n2399 VDD.n2398 185
R13046 VDD.n2397 VDD.n359 185
R13047 VDD.n2393 VDD.n2392 185
R13048 VDD.n2390 VDD.n364 185
R13049 VDD.n2388 VDD.n2387 185
R13050 VDD.n366 VDD.n365 185
R13051 VDD.n2349 VDD.n2347 185
R13052 VDD.n2383 VDD.n2350 185
R13053 VDD.n2382 VDD.n2381 185
R13054 VDD.n2379 VDD.n2351 185
R13055 VDD.n2377 VDD.n2376 185
R13056 VDD.n2375 VDD.n2352 185
R13057 VDD.n2374 VDD.n2373 185
R13058 VDD.n2371 VDD.n2357 185
R13059 VDD.n2369 VDD.n2368 185
R13060 VDD.n2367 VDD.n2359 185
R13061 VDD.n2363 VDD.n297 185
R13062 VDD.n2623 VDD.n2622 185
R13063 VDD.n2627 VDD.n199 185
R13064 VDD.n2629 VDD.n2628 185
R13065 VDD.n2631 VDD.n197 185
R13066 VDD.n2633 VDD.n2632 185
R13067 VDD.n2634 VDD.n192 185
R13068 VDD.n2636 VDD.n2635 185
R13069 VDD.n2638 VDD.n190 185
R13070 VDD.n2640 VDD.n2639 185
R13071 VDD.n2641 VDD.n185 185
R13072 VDD.n2643 VDD.n2642 185
R13073 VDD.n2645 VDD.n183 185
R13074 VDD.n2647 VDD.n2646 185
R13075 VDD.n2648 VDD.n175 185
R13076 VDD.n2650 VDD.n2649 185
R13077 VDD.n2652 VDD.n173 185
R13078 VDD.n2654 VDD.n2653 185
R13079 VDD.n2655 VDD.n168 185
R13080 VDD.n2657 VDD.n2656 185
R13081 VDD.n2659 VDD.n166 185
R13082 VDD.n2661 VDD.n2660 185
R13083 VDD.n2662 VDD.n161 185
R13084 VDD.n2664 VDD.n2663 185
R13085 VDD.n2666 VDD.n159 185
R13086 VDD.n2668 VDD.n2667 185
R13087 VDD.n2669 VDD.n154 185
R13088 VDD.n2671 VDD.n2670 185
R13089 VDD.n2673 VDD.n152 185
R13090 VDD.n2675 VDD.n2674 185
R13091 VDD.n2679 VDD.n147 185
R13092 VDD.n2681 VDD.n2680 185
R13093 VDD.n2683 VDD.n145 185
R13094 VDD.n2685 VDD.n2684 185
R13095 VDD.n2686 VDD.n140 185
R13096 VDD.n2688 VDD.n2687 185
R13097 VDD.n2690 VDD.n138 185
R13098 VDD.n2692 VDD.n2691 185
R13099 VDD.n2693 VDD.n133 185
R13100 VDD.n2695 VDD.n2694 185
R13101 VDD.n2697 VDD.n131 185
R13102 VDD.n2699 VDD.n2698 185
R13103 VDD.n2700 VDD.n126 185
R13104 VDD.n2702 VDD.n2701 185
R13105 VDD.n2704 VDD.n124 185
R13106 VDD.n2706 VDD.n2705 185
R13107 VDD.n2707 VDD.n117 185
R13108 VDD.n2709 VDD.n2708 185
R13109 VDD.n2711 VDD.n115 185
R13110 VDD.n2713 VDD.n2712 185
R13111 VDD.n2714 VDD.n110 185
R13112 VDD.n2716 VDD.n2715 185
R13113 VDD.n2718 VDD.n108 185
R13114 VDD.n2720 VDD.n2719 185
R13115 VDD.n2721 VDD.n106 185
R13116 VDD.n2722 VDD.n103 185
R13117 VDD.n103 VDD.n102 185
R13118 VDD.n2618 VDD.n101 185
R13119 VDD.n2727 VDD.n101 185
R13120 VDD.n2617 VDD.n100 185
R13121 VDD.n2728 VDD.n100 185
R13122 VDD.n2616 VDD.n99 185
R13123 VDD.n2729 VDD.n99 185
R13124 VDD.n205 VDD.n204 185
R13125 VDD.n204 VDD.n91 185
R13126 VDD.n2612 VDD.n90 185
R13127 VDD.n2735 VDD.n90 185
R13128 VDD.n2611 VDD.n89 185
R13129 VDD.n2736 VDD.n89 185
R13130 VDD.n2610 VDD.n88 185
R13131 VDD.n2737 VDD.n88 185
R13132 VDD.n208 VDD.n207 185
R13133 VDD.n207 VDD.n80 185
R13134 VDD.n2606 VDD.n79 185
R13135 VDD.n2743 VDD.n79 185
R13136 VDD.n2605 VDD.n78 185
R13137 VDD.n2744 VDD.n78 185
R13138 VDD.n2604 VDD.n77 185
R13139 VDD.n2745 VDD.n77 185
R13140 VDD.n211 VDD.n210 185
R13141 VDD.n210 VDD.n69 185
R13142 VDD.n2600 VDD.n68 185
R13143 VDD.n2751 VDD.n68 185
R13144 VDD.n2599 VDD.n67 185
R13145 VDD.n2752 VDD.n67 185
R13146 VDD.n2598 VDD.n66 185
R13147 VDD.n2753 VDD.n66 185
R13148 VDD.n214 VDD.n213 185
R13149 VDD.n213 VDD.n58 185
R13150 VDD.n2594 VDD.n57 185
R13151 VDD.n2759 VDD.n57 185
R13152 VDD.n2593 VDD.n56 185
R13153 VDD.n2760 VDD.n56 185
R13154 VDD.n2592 VDD.n55 185
R13155 VDD.n2761 VDD.n55 185
R13156 VDD.n217 VDD.n216 185
R13157 VDD.n216 VDD.n47 185
R13158 VDD.n2588 VDD.n46 185
R13159 VDD.n2767 VDD.n46 185
R13160 VDD.n2587 VDD.n45 185
R13161 VDD.n2768 VDD.n45 185
R13162 VDD.n2586 VDD.n44 185
R13163 VDD.n2769 VDD.n44 185
R13164 VDD.n220 VDD.n219 185
R13165 VDD.n219 VDD.n37 185
R13166 VDD.n2582 VDD.n36 185
R13167 VDD.n2775 VDD.n36 185
R13168 VDD.n2581 VDD.n35 185
R13169 VDD.n2776 VDD.n35 185
R13170 VDD.n2580 VDD.n34 185
R13171 VDD.t2 VDD.n34 185
R13172 VDD.n226 VDD.n222 185
R13173 VDD.n226 VDD.n33 185
R13174 VDD.n2576 VDD.n2575 185
R13175 VDD.n2575 VDD.n2574 185
R13176 VDD.n225 VDD.n224 185
R13177 VDD.n227 VDD.n225 185
R13178 VDD.n2565 VDD.n2564 185
R13179 VDD.n2566 VDD.n2565 185
R13180 VDD.n235 VDD.n234 185
R13181 VDD.n234 VDD.n233 185
R13182 VDD.n2560 VDD.n2559 185
R13183 VDD.n2559 VDD.n2558 185
R13184 VDD.n238 VDD.n237 185
R13185 VDD.n239 VDD.n238 185
R13186 VDD.n2549 VDD.n2548 185
R13187 VDD.n2550 VDD.n2549 185
R13188 VDD.n246 VDD.n245 185
R13189 VDD.n251 VDD.n245 185
R13190 VDD.n2544 VDD.n2543 185
R13191 VDD.n2543 VDD.n2542 185
R13192 VDD.n249 VDD.n248 185
R13193 VDD.n250 VDD.n249 185
R13194 VDD.n2533 VDD.n2532 185
R13195 VDD.n2534 VDD.n2533 185
R13196 VDD.n259 VDD.n258 185
R13197 VDD.n258 VDD.n257 185
R13198 VDD.n2528 VDD.n2527 185
R13199 VDD.n2527 VDD.n2526 185
R13200 VDD.n262 VDD.n261 185
R13201 VDD.n263 VDD.n262 185
R13202 VDD.n2517 VDD.n2516 185
R13203 VDD.n2518 VDD.n2517 185
R13204 VDD.n271 VDD.n270 185
R13205 VDD.n270 VDD.n269 185
R13206 VDD.n2512 VDD.n2511 185
R13207 VDD.n2511 VDD.n2510 185
R13208 VDD.n274 VDD.n273 185
R13209 VDD.n275 VDD.n274 185
R13210 VDD.n2501 VDD.n2500 185
R13211 VDD.n2502 VDD.n2501 185
R13212 VDD.n282 VDD.n281 185
R13213 VDD.n287 VDD.n281 185
R13214 VDD.n2496 VDD.n2495 185
R13215 VDD.n2495 VDD.n2494 185
R13216 VDD.n285 VDD.n284 185
R13217 VDD.n286 VDD.n285 185
R13218 VDD.n2485 VDD.n2484 185
R13219 VDD.n2486 VDD.n2485 185
R13220 VDD.n295 VDD.n294 185
R13221 VDD.n294 VDD.n293 185
R13222 VDD.n2480 VDD.n2479 185
R13223 VDD.n2479 VDD.n2478 185
R13224 VDD.n2477 VDD.n2476 185
R13225 VDD.n2478 VDD.n2477 185
R13226 VDD.n292 VDD.n291 185
R13227 VDD.n293 VDD.n292 185
R13228 VDD.n2488 VDD.n2487 185
R13229 VDD.n2487 VDD.n2486 185
R13230 VDD.n289 VDD.n288 185
R13231 VDD.n288 VDD.n286 185
R13232 VDD.n2493 VDD.n2492 185
R13233 VDD.n2494 VDD.n2493 185
R13234 VDD.n280 VDD.n279 185
R13235 VDD.n287 VDD.n280 185
R13236 VDD.n2504 VDD.n2503 185
R13237 VDD.n2503 VDD.n2502 185
R13238 VDD.n277 VDD.n276 185
R13239 VDD.n276 VDD.n275 185
R13240 VDD.n2509 VDD.n2508 185
R13241 VDD.n2510 VDD.n2509 185
R13242 VDD.n268 VDD.n267 185
R13243 VDD.n269 VDD.n268 185
R13244 VDD.n2520 VDD.n2519 185
R13245 VDD.n2519 VDD.n2518 185
R13246 VDD.n265 VDD.n264 185
R13247 VDD.n264 VDD.n263 185
R13248 VDD.n2525 VDD.n2524 185
R13249 VDD.n2526 VDD.n2525 185
R13250 VDD.n256 VDD.n255 185
R13251 VDD.n257 VDD.n256 185
R13252 VDD.n2536 VDD.n2535 185
R13253 VDD.n2535 VDD.n2534 185
R13254 VDD.n253 VDD.n252 185
R13255 VDD.n252 VDD.n250 185
R13256 VDD.n2541 VDD.n2540 185
R13257 VDD.n2542 VDD.n2541 185
R13258 VDD.n244 VDD.n243 185
R13259 VDD.n251 VDD.n244 185
R13260 VDD.n2552 VDD.n2551 185
R13261 VDD.n2551 VDD.n2550 185
R13262 VDD.n241 VDD.n240 185
R13263 VDD.n240 VDD.n239 185
R13264 VDD.n2557 VDD.n2556 185
R13265 VDD.n2558 VDD.n2557 185
R13266 VDD.n232 VDD.n231 185
R13267 VDD.n233 VDD.n232 185
R13268 VDD.n2568 VDD.n2567 185
R13269 VDD.n2567 VDD.n2566 185
R13270 VDD.n229 VDD.n228 185
R13271 VDD.n228 VDD.n227 185
R13272 VDD.n2573 VDD.n2572 185
R13273 VDD.n2574 VDD.n2573 185
R13274 VDD.n31 VDD.n29 185
R13275 VDD.n33 VDD.n31 185
R13276 VDD.n2778 VDD.n2777 185
R13277 VDD.n2777 VDD.t2 185
R13278 VDD.n32 VDD.n30 185
R13279 VDD.n2776 VDD.n32 185
R13280 VDD.n2774 VDD.n2773 185
R13281 VDD.n2775 VDD.n2774 185
R13282 VDD.n2772 VDD.n38 185
R13283 VDD.n38 VDD.n37 185
R13284 VDD.n2771 VDD.n2770 185
R13285 VDD.n2770 VDD.n2769 185
R13286 VDD.n43 VDD.n42 185
R13287 VDD.n2768 VDD.n43 185
R13288 VDD.n2766 VDD.n2765 185
R13289 VDD.n2767 VDD.n2766 185
R13290 VDD.n2764 VDD.n48 185
R13291 VDD.n48 VDD.n47 185
R13292 VDD.n2763 VDD.n2762 185
R13293 VDD.n2762 VDD.n2761 185
R13294 VDD.n54 VDD.n53 185
R13295 VDD.n2760 VDD.n54 185
R13296 VDD.n2758 VDD.n2757 185
R13297 VDD.n2759 VDD.n2758 185
R13298 VDD.n2756 VDD.n59 185
R13299 VDD.n59 VDD.n58 185
R13300 VDD.n2755 VDD.n2754 185
R13301 VDD.n2754 VDD.n2753 185
R13302 VDD.n65 VDD.n64 185
R13303 VDD.n2752 VDD.n65 185
R13304 VDD.n2750 VDD.n2749 185
R13305 VDD.n2751 VDD.n2750 185
R13306 VDD.n2748 VDD.n70 185
R13307 VDD.n70 VDD.n69 185
R13308 VDD.n2747 VDD.n2746 185
R13309 VDD.n2746 VDD.n2745 185
R13310 VDD.n76 VDD.n75 185
R13311 VDD.n2744 VDD.n76 185
R13312 VDD.n2742 VDD.n2741 185
R13313 VDD.n2743 VDD.n2742 185
R13314 VDD.n2740 VDD.n81 185
R13315 VDD.n81 VDD.n80 185
R13316 VDD.n2739 VDD.n2738 185
R13317 VDD.n2738 VDD.n2737 185
R13318 VDD.n87 VDD.n86 185
R13319 VDD.n2736 VDD.n87 185
R13320 VDD.n2734 VDD.n2733 185
R13321 VDD.n2735 VDD.n2734 185
R13322 VDD.n2732 VDD.n92 185
R13323 VDD.n92 VDD.n91 185
R13324 VDD.n2731 VDD.n2730 185
R13325 VDD.n2730 VDD.n2729 185
R13326 VDD.n98 VDD.n97 185
R13327 VDD.n2728 VDD.n98 185
R13328 VDD.n2726 VDD.n2725 185
R13329 VDD.n2727 VDD.n2726 185
R13330 VDD.n556 VDD.n554 185
R13331 VDD.n554 VDD.n537 185
R13332 VDD.n1828 VDD.n563 185
R13333 VDD.n1883 VDD.n563 185
R13334 VDD.n1830 VDD.n1829 185
R13335 VDD.n1829 VDD.n561 185
R13336 VDD.n1831 VDD.n574 185
R13337 VDD.n1841 VDD.n574 185
R13338 VDD.n1832 VDD.n581 185
R13339 VDD.n581 VDD.n572 185
R13340 VDD.n1834 VDD.n1833 185
R13341 VDD.n1835 VDD.n1834 185
R13342 VDD.n1827 VDD.n580 185
R13343 VDD.n586 VDD.n580 185
R13344 VDD.n1826 VDD.n1825 185
R13345 VDD.n1825 VDD.n1824 185
R13346 VDD.n583 VDD.n582 185
R13347 VDD.n593 VDD.n583 185
R13348 VDD.n1817 VDD.n1816 185
R13349 VDD.n1818 VDD.n1817 185
R13350 VDD.n1815 VDD.n594 185
R13351 VDD.n594 VDD.n590 185
R13352 VDD.n1814 VDD.n1813 185
R13353 VDD.n1813 VDD.n1812 185
R13354 VDD.n596 VDD.n595 185
R13355 VDD.n597 VDD.n596 185
R13356 VDD.n1805 VDD.n1804 185
R13357 VDD.n1806 VDD.n1805 185
R13358 VDD.n1803 VDD.n606 185
R13359 VDD.n606 VDD.n603 185
R13360 VDD.n1802 VDD.n1801 185
R13361 VDD.n1801 VDD.n1800 185
R13362 VDD.n608 VDD.n607 185
R13363 VDD.n609 VDD.n608 185
R13364 VDD.n1793 VDD.n1792 185
R13365 VDD.n1794 VDD.n1793 185
R13366 VDD.n1791 VDD.n618 185
R13367 VDD.n618 VDD.n615 185
R13368 VDD.n1790 VDD.n1789 185
R13369 VDD.n1789 VDD.n1788 185
R13370 VDD.n620 VDD.n619 185
R13371 VDD.n621 VDD.n620 185
R13372 VDD.n1781 VDD.n1780 185
R13373 VDD.n1782 VDD.n1781 185
R13374 VDD.n1779 VDD.n630 185
R13375 VDD.n630 VDD.n627 185
R13376 VDD.n1778 VDD.n1777 185
R13377 VDD.n1777 VDD.t16 185
R13378 VDD.n632 VDD.n631 185
R13379 VDD.n633 VDD.n632 185
R13380 VDD.n1770 VDD.n1769 185
R13381 VDD.n1771 VDD.n1770 185
R13382 VDD.n1768 VDD.n642 185
R13383 VDD.n642 VDD.n639 185
R13384 VDD.n1767 VDD.n1766 185
R13385 VDD.n1766 VDD.n1765 185
R13386 VDD.n644 VDD.n643 185
R13387 VDD.t17 VDD.n644 185
R13388 VDD.n1758 VDD.n1757 185
R13389 VDD.n1759 VDD.n1758 185
R13390 VDD.n1756 VDD.n653 185
R13391 VDD.n653 VDD.n650 185
R13392 VDD.n1755 VDD.n1754 185
R13393 VDD.n1754 VDD.n1753 185
R13394 VDD.n655 VDD.n654 185
R13395 VDD.n656 VDD.n655 185
R13396 VDD.n1746 VDD.n1745 185
R13397 VDD.n1747 VDD.n1746 185
R13398 VDD.n1744 VDD.n665 185
R13399 VDD.n665 VDD.n662 185
R13400 VDD.n1743 VDD.n1742 185
R13401 VDD.n1742 VDD.n1741 185
R13402 VDD.n667 VDD.n666 185
R13403 VDD.n668 VDD.n667 185
R13404 VDD.n1734 VDD.n1733 185
R13405 VDD.n1735 VDD.n1734 185
R13406 VDD.n1732 VDD.n677 185
R13407 VDD.n677 VDD.n674 185
R13408 VDD.n1731 VDD.n1730 185
R13409 VDD.n1730 VDD.n1729 185
R13410 VDD.n679 VDD.n678 185
R13411 VDD.n688 VDD.n679 185
R13412 VDD.n1722 VDD.n1721 185
R13413 VDD.n1723 VDD.n1722 185
R13414 VDD.n1720 VDD.n689 185
R13415 VDD.n689 VDD.n685 185
R13416 VDD.n1719 VDD.n1718 185
R13417 VDD.n1718 VDD.n1717 185
R13418 VDD.n691 VDD.n690 185
R13419 VDD.n692 VDD.n691 185
R13420 VDD.n1710 VDD.n1709 185
R13421 VDD.n1711 VDD.n1710 185
R13422 VDD.n1708 VDD.n701 185
R13423 VDD.n701 VDD.n698 185
R13424 VDD.n1887 VDD.n553 185
R13425 VDD.n1918 VDD.n553 185
R13426 VDD.n1889 VDD.n1888 185
R13427 VDD.n1891 VDD.n1890 185
R13428 VDD.n1893 VDD.n1892 185
R13429 VDD.n1896 VDD.n1895 185
R13430 VDD.n1898 VDD.n1897 185
R13431 VDD.n1900 VDD.n1899 185
R13432 VDD.n1902 VDD.n1901 185
R13433 VDD.n1904 VDD.n1903 185
R13434 VDD.n1906 VDD.n1905 185
R13435 VDD.n1908 VDD.n1907 185
R13436 VDD.n1910 VDD.n1909 185
R13437 VDD.n1912 VDD.n1911 185
R13438 VDD.n1914 VDD.n1913 185
R13439 VDD.n1915 VDD.n555 185
R13440 VDD.n1917 VDD.n1916 185
R13441 VDD.n1918 VDD.n1917 185
R13442 VDD.n1886 VDD.n1885 185
R13443 VDD.n1885 VDD.n537 185
R13444 VDD.n1884 VDD.n559 185
R13445 VDD.n1884 VDD.n1883 185
R13446 VDD.n801 VDD.n560 185
R13447 VDD.n561 VDD.n560 185
R13448 VDD.n802 VDD.n573 185
R13449 VDD.n1841 VDD.n573 185
R13450 VDD.n804 VDD.n803 185
R13451 VDD.n803 VDD.n572 185
R13452 VDD.n805 VDD.n579 185
R13453 VDD.n1835 VDD.n579 185
R13454 VDD.n807 VDD.n806 185
R13455 VDD.n806 VDD.n586 185
R13456 VDD.n808 VDD.n585 185
R13457 VDD.n1824 VDD.n585 185
R13458 VDD.n810 VDD.n809 185
R13459 VDD.n809 VDD.n593 185
R13460 VDD.n811 VDD.n592 185
R13461 VDD.n1818 VDD.n592 185
R13462 VDD.n813 VDD.n812 185
R13463 VDD.n812 VDD.n590 185
R13464 VDD.n814 VDD.n599 185
R13465 VDD.n1812 VDD.n599 185
R13466 VDD.n816 VDD.n815 185
R13467 VDD.n815 VDD.n597 185
R13468 VDD.n817 VDD.n605 185
R13469 VDD.n1806 VDD.n605 185
R13470 VDD.n819 VDD.n818 185
R13471 VDD.n818 VDD.n603 185
R13472 VDD.n820 VDD.n611 185
R13473 VDD.n1800 VDD.n611 185
R13474 VDD.n822 VDD.n821 185
R13475 VDD.n821 VDD.n609 185
R13476 VDD.n823 VDD.n617 185
R13477 VDD.n1794 VDD.n617 185
R13478 VDD.n825 VDD.n824 185
R13479 VDD.n824 VDD.n615 185
R13480 VDD.n826 VDD.n623 185
R13481 VDD.n1788 VDD.n623 185
R13482 VDD.n828 VDD.n827 185
R13483 VDD.n827 VDD.n621 185
R13484 VDD.n829 VDD.n629 185
R13485 VDD.n1782 VDD.n629 185
R13486 VDD.n831 VDD.n830 185
R13487 VDD.n830 VDD.n627 185
R13488 VDD.n832 VDD.n634 185
R13489 VDD.t16 VDD.n634 185
R13490 VDD.n834 VDD.n833 185
R13491 VDD.n833 VDD.n633 185
R13492 VDD.n835 VDD.n641 185
R13493 VDD.n1771 VDD.n641 185
R13494 VDD.n837 VDD.n836 185
R13495 VDD.n836 VDD.n639 185
R13496 VDD.n838 VDD.n646 185
R13497 VDD.n1765 VDD.n646 185
R13498 VDD.n840 VDD.n839 185
R13499 VDD.n839 VDD.t17 185
R13500 VDD.n841 VDD.n652 185
R13501 VDD.n1759 VDD.n652 185
R13502 VDD.n843 VDD.n842 185
R13503 VDD.n842 VDD.n650 185
R13504 VDD.n844 VDD.n658 185
R13505 VDD.n1753 VDD.n658 185
R13506 VDD.n846 VDD.n845 185
R13507 VDD.n845 VDD.n656 185
R13508 VDD.n847 VDD.n664 185
R13509 VDD.n1747 VDD.n664 185
R13510 VDD.n849 VDD.n848 185
R13511 VDD.n848 VDD.n662 185
R13512 VDD.n850 VDD.n670 185
R13513 VDD.n1741 VDD.n670 185
R13514 VDD.n852 VDD.n851 185
R13515 VDD.n851 VDD.n668 185
R13516 VDD.n853 VDD.n676 185
R13517 VDD.n1735 VDD.n676 185
R13518 VDD.n855 VDD.n854 185
R13519 VDD.n854 VDD.n674 185
R13520 VDD.n856 VDD.n681 185
R13521 VDD.n1729 VDD.n681 185
R13522 VDD.n858 VDD.n857 185
R13523 VDD.n857 VDD.n688 185
R13524 VDD.n859 VDD.n687 185
R13525 VDD.n1723 VDD.n687 185
R13526 VDD.n861 VDD.n860 185
R13527 VDD.n860 VDD.n685 185
R13528 VDD.n862 VDD.n694 185
R13529 VDD.n1717 VDD.n694 185
R13530 VDD.n864 VDD.n863 185
R13531 VDD.n863 VDD.n692 185
R13532 VDD.n865 VDD.n700 185
R13533 VDD.n1711 VDD.n700 185
R13534 VDD.n867 VDD.n866 185
R13535 VDD.n866 VDD.n698 185
R13536 VDD.n1707 VDD.n1706 185
R13537 VDD.n1706 VDD.n1705 185
R13538 VDD.n703 VDD.n702 185
R13539 VDD.n788 VDD.n787 185
R13540 VDD.n790 VDD.n789 185
R13541 VDD.n792 VDD.n791 185
R13542 VDD.n794 VDD.n793 185
R13543 VDD.n796 VDD.n795 185
R13544 VDD.n798 VDD.n797 185
R13545 VDD.n883 VDD.n882 185
R13546 VDD.n881 VDD.n880 185
R13547 VDD.n879 VDD.n878 185
R13548 VDD.n877 VDD.n876 185
R13549 VDD.n874 VDD.n873 185
R13550 VDD.n872 VDD.n871 185
R13551 VDD.n870 VDD.n869 185
R13552 VDD.n868 VDD.n718 185
R13553 VDD.n1705 VDD.n718 185
R13554 VDD.n800 VDD.t127 170.506
R13555 VDD.n558 VDD.t81 170.506
R13556 VDD.n1608 VDD.t124 170.506
R13557 VDD.n568 VDD.t118 170.506
R13558 VDD.n1934 VDD.t54 170.506
R13559 VDD.n399 VDD.t109 170.506
R13560 VDD.n2033 VDD.t120 170.506
R13561 VDD.n376 VDD.t77 170.506
R13562 VDD.n9 VDD.n7 169.231
R13563 VDD.n2 VDD.n0 169.231
R13564 VDD.n9 VDD.n8 168.121
R13565 VDD.n11 VDD.n10 168.121
R13566 VDD.n13 VDD.n12 168.121
R13567 VDD.n6 VDD.n5 168.121
R13568 VDD.n4 VDD.n3 168.121
R13569 VDD.n2 VDD.n1 168.121
R13570 VDD.t15 VDD.t32 165.109
R13571 VDD.t24 VDD.t140 165.109
R13572 VDD.n2477 VDD.n292 146.341
R13573 VDD.n2487 VDD.n292 146.341
R13574 VDD.n2487 VDD.n288 146.341
R13575 VDD.n2493 VDD.n288 146.341
R13576 VDD.n2493 VDD.n280 146.341
R13577 VDD.n2503 VDD.n280 146.341
R13578 VDD.n2503 VDD.n276 146.341
R13579 VDD.n2509 VDD.n276 146.341
R13580 VDD.n2509 VDD.n268 146.341
R13581 VDD.n2519 VDD.n268 146.341
R13582 VDD.n2519 VDD.n264 146.341
R13583 VDD.n2525 VDD.n264 146.341
R13584 VDD.n2525 VDD.n256 146.341
R13585 VDD.n2535 VDD.n256 146.341
R13586 VDD.n2535 VDD.n252 146.341
R13587 VDD.n2541 VDD.n252 146.341
R13588 VDD.n2541 VDD.n244 146.341
R13589 VDD.n2551 VDD.n244 146.341
R13590 VDD.n2551 VDD.n240 146.341
R13591 VDD.n2557 VDD.n240 146.341
R13592 VDD.n2557 VDD.n232 146.341
R13593 VDD.n2567 VDD.n232 146.341
R13594 VDD.n2567 VDD.n228 146.341
R13595 VDD.n2573 VDD.n228 146.341
R13596 VDD.n2573 VDD.n31 146.341
R13597 VDD.n2777 VDD.n31 146.341
R13598 VDD.n2777 VDD.n32 146.341
R13599 VDD.n2774 VDD.n32 146.341
R13600 VDD.n2774 VDD.n38 146.341
R13601 VDD.n2770 VDD.n38 146.341
R13602 VDD.n2770 VDD.n43 146.341
R13603 VDD.n2766 VDD.n43 146.341
R13604 VDD.n2766 VDD.n48 146.341
R13605 VDD.n2762 VDD.n48 146.341
R13606 VDD.n2762 VDD.n54 146.341
R13607 VDD.n2758 VDD.n54 146.341
R13608 VDD.n2758 VDD.n59 146.341
R13609 VDD.n2754 VDD.n59 146.341
R13610 VDD.n2754 VDD.n65 146.341
R13611 VDD.n2750 VDD.n65 146.341
R13612 VDD.n2750 VDD.n70 146.341
R13613 VDD.n2746 VDD.n70 146.341
R13614 VDD.n2746 VDD.n76 146.341
R13615 VDD.n2742 VDD.n76 146.341
R13616 VDD.n2742 VDD.n81 146.341
R13617 VDD.n2738 VDD.n81 146.341
R13618 VDD.n2738 VDD.n87 146.341
R13619 VDD.n2734 VDD.n87 146.341
R13620 VDD.n2734 VDD.n92 146.341
R13621 VDD.n2730 VDD.n92 146.341
R13622 VDD.n2730 VDD.n98 146.341
R13623 VDD.n2726 VDD.n98 146.341
R13624 VDD.n106 VDD.n103 146.341
R13625 VDD.n2719 VDD.n2718 146.341
R13626 VDD.n2716 VDD.n110 146.341
R13627 VDD.n2712 VDD.n2711 146.341
R13628 VDD.n2709 VDD.n117 146.341
R13629 VDD.n2705 VDD.n2704 146.341
R13630 VDD.n2702 VDD.n126 146.341
R13631 VDD.n2698 VDD.n2697 146.341
R13632 VDD.n2695 VDD.n133 146.341
R13633 VDD.n2691 VDD.n2690 146.341
R13634 VDD.n2688 VDD.n140 146.341
R13635 VDD.n2684 VDD.n2683 146.341
R13636 VDD.n2681 VDD.n147 146.341
R13637 VDD.n2674 VDD.n2673 146.341
R13638 VDD.n2671 VDD.n154 146.341
R13639 VDD.n2667 VDD.n2666 146.341
R13640 VDD.n2664 VDD.n161 146.341
R13641 VDD.n2660 VDD.n2659 146.341
R13642 VDD.n2657 VDD.n168 146.341
R13643 VDD.n2653 VDD.n2652 146.341
R13644 VDD.n2650 VDD.n175 146.341
R13645 VDD.n2646 VDD.n2645 146.341
R13646 VDD.n2643 VDD.n185 146.341
R13647 VDD.n2639 VDD.n2638 146.341
R13648 VDD.n2636 VDD.n192 146.341
R13649 VDD.n2632 VDD.n2631 146.341
R13650 VDD.n2629 VDD.n199 146.341
R13651 VDD.n2479 VDD.n294 146.341
R13652 VDD.n2485 VDD.n294 146.341
R13653 VDD.n2485 VDD.n285 146.341
R13654 VDD.n2495 VDD.n285 146.341
R13655 VDD.n2495 VDD.n281 146.341
R13656 VDD.n2501 VDD.n281 146.341
R13657 VDD.n2501 VDD.n274 146.341
R13658 VDD.n2511 VDD.n274 146.341
R13659 VDD.n2511 VDD.n270 146.341
R13660 VDD.n2517 VDD.n270 146.341
R13661 VDD.n2517 VDD.n262 146.341
R13662 VDD.n2527 VDD.n262 146.341
R13663 VDD.n2527 VDD.n258 146.341
R13664 VDD.n2533 VDD.n258 146.341
R13665 VDD.n2533 VDD.n249 146.341
R13666 VDD.n2543 VDD.n249 146.341
R13667 VDD.n2543 VDD.n245 146.341
R13668 VDD.n2549 VDD.n245 146.341
R13669 VDD.n2549 VDD.n238 146.341
R13670 VDD.n2559 VDD.n238 146.341
R13671 VDD.n2559 VDD.n234 146.341
R13672 VDD.n2565 VDD.n234 146.341
R13673 VDD.n2565 VDD.n225 146.341
R13674 VDD.n2575 VDD.n225 146.341
R13675 VDD.n2575 VDD.n226 146.341
R13676 VDD.n226 VDD.n34 146.341
R13677 VDD.n35 VDD.n34 146.341
R13678 VDD.n36 VDD.n35 146.341
R13679 VDD.n219 VDD.n36 146.341
R13680 VDD.n219 VDD.n44 146.341
R13681 VDD.n45 VDD.n44 146.341
R13682 VDD.n46 VDD.n45 146.341
R13683 VDD.n216 VDD.n46 146.341
R13684 VDD.n216 VDD.n55 146.341
R13685 VDD.n56 VDD.n55 146.341
R13686 VDD.n57 VDD.n56 146.341
R13687 VDD.n213 VDD.n57 146.341
R13688 VDD.n213 VDD.n66 146.341
R13689 VDD.n67 VDD.n66 146.341
R13690 VDD.n68 VDD.n67 146.341
R13691 VDD.n210 VDD.n68 146.341
R13692 VDD.n210 VDD.n77 146.341
R13693 VDD.n78 VDD.n77 146.341
R13694 VDD.n79 VDD.n78 146.341
R13695 VDD.n207 VDD.n79 146.341
R13696 VDD.n207 VDD.n88 146.341
R13697 VDD.n89 VDD.n88 146.341
R13698 VDD.n90 VDD.n89 146.341
R13699 VDD.n204 VDD.n90 146.341
R13700 VDD.n204 VDD.n99 146.341
R13701 VDD.n100 VDD.n99 146.341
R13702 VDD.n101 VDD.n100 146.341
R13703 VDD.n2471 VDD.n2469 146.341
R13704 VDD.n2469 VDD.n2468 146.341
R13705 VDD.n2465 VDD.n2464 146.341
R13706 VDD.n2462 VDD.n307 146.341
R13707 VDD.n2458 VDD.n2456 146.341
R13708 VDD.n2454 VDD.n313 146.341
R13709 VDD.n2448 VDD.n318 146.341
R13710 VDD.n2446 VDD.n2445 146.341
R13711 VDD.n2442 VDD.n2441 146.341
R13712 VDD.n2439 VDD.n326 146.341
R13713 VDD.n2435 VDD.n2433 146.341
R13714 VDD.n2431 VDD.n332 146.341
R13715 VDD.n2427 VDD.n2425 146.341
R13716 VDD.n2423 VDD.n338 146.341
R13717 VDD.n2419 VDD.n2417 146.341
R13718 VDD.n2415 VDD.n347 146.341
R13719 VDD.n2411 VDD.n2409 146.341
R13720 VDD.n2407 VDD.n353 146.341
R13721 VDD.n2403 VDD.n2401 146.341
R13722 VDD.n2399 VDD.n359 146.341
R13723 VDD.n2392 VDD.n2390 146.341
R13724 VDD.n2388 VDD.n365 146.341
R13725 VDD.n2350 VDD.n2349 146.341
R13726 VDD.n2381 VDD.n2379 146.341
R13727 VDD.n2377 VDD.n2352 146.341
R13728 VDD.n2373 VDD.n2371 146.341
R13729 VDD.n2369 VDD.n2359 146.341
R13730 VDD.n1517 VDD.n917 146.341
R13731 VDD.n1515 VDD.n1514 146.341
R13732 VDD.n1512 VDD.n1497 146.341
R13733 VDD.n1508 VDD.n1507 146.341
R13734 VDD.n1603 VDD.n726 146.341
R13735 VDD.n1601 VDD.n1600 146.341
R13736 VDD.n1598 VDD.n731 146.341
R13737 VDD.n1594 VDD.n1593 146.341
R13738 VDD.n1591 VDD.n735 146.341
R13739 VDD.n1587 VDD.n1586 146.341
R13740 VDD.n1584 VDD.n742 146.341
R13741 VDD.n1580 VDD.n1579 146.341
R13742 VDD.n1577 VDD.n749 146.341
R13743 VDD.n1570 VDD.n1569 146.341
R13744 VDD.n1567 VDD.n756 146.341
R13745 VDD.n1563 VDD.n1562 146.341
R13746 VDD.n1560 VDD.n763 146.341
R13747 VDD.n1556 VDD.n1555 146.341
R13748 VDD.n1553 VDD.n770 146.341
R13749 VDD.n1549 VDD.n1548 146.341
R13750 VDD.n1546 VDD.n777 146.341
R13751 VDD.n888 VDD.n785 146.341
R13752 VDD.n892 VDD.n891 146.341
R13753 VDD.n895 VDD.n894 146.341
R13754 VDD.n900 VDD.n897 146.341
R13755 VDD.n903 VDD.n902 146.341
R13756 VDD.n911 VDD.n905 146.341
R13757 VDD.n1278 VDD.n1068 146.341
R13758 VDD.n1284 VDD.n1068 146.341
R13759 VDD.n1284 VDD.n1059 146.341
R13760 VDD.n1294 VDD.n1059 146.341
R13761 VDD.n1294 VDD.n1055 146.341
R13762 VDD.n1300 VDD.n1055 146.341
R13763 VDD.n1300 VDD.n1048 146.341
R13764 VDD.n1310 VDD.n1048 146.341
R13765 VDD.n1310 VDD.n1044 146.341
R13766 VDD.n1316 VDD.n1044 146.341
R13767 VDD.n1316 VDD.n1036 146.341
R13768 VDD.n1326 VDD.n1036 146.341
R13769 VDD.n1326 VDD.n1032 146.341
R13770 VDD.n1332 VDD.n1032 146.341
R13771 VDD.n1332 VDD.n1023 146.341
R13772 VDD.n1342 VDD.n1023 146.341
R13773 VDD.n1342 VDD.n1019 146.341
R13774 VDD.n1348 VDD.n1019 146.341
R13775 VDD.n1348 VDD.n1012 146.341
R13776 VDD.n1358 VDD.n1012 146.341
R13777 VDD.n1358 VDD.n1008 146.341
R13778 VDD.n1364 VDD.n1008 146.341
R13779 VDD.n1364 VDD.n1000 146.341
R13780 VDD.n1374 VDD.n1000 146.341
R13781 VDD.n1374 VDD.n996 146.341
R13782 VDD.n1380 VDD.n996 146.341
R13783 VDD.n1380 VDD.n988 146.341
R13784 VDD.n1401 VDD.n988 146.341
R13785 VDD.n1401 VDD.n984 146.341
R13786 VDD.n1407 VDD.n984 146.341
R13787 VDD.n1407 VDD.n976 146.341
R13788 VDD.n1417 VDD.n976 146.341
R13789 VDD.n1417 VDD.n972 146.341
R13790 VDD.n1423 VDD.n972 146.341
R13791 VDD.n1423 VDD.n964 146.341
R13792 VDD.n1433 VDD.n964 146.341
R13793 VDD.n1433 VDD.n960 146.341
R13794 VDD.n1439 VDD.n960 146.341
R13795 VDD.n1439 VDD.n952 146.341
R13796 VDD.n1449 VDD.n952 146.341
R13797 VDD.n1449 VDD.n948 146.341
R13798 VDD.n1455 VDD.n948 146.341
R13799 VDD.n1455 VDD.n940 146.341
R13800 VDD.n1465 VDD.n940 146.341
R13801 VDD.n1465 VDD.n936 146.341
R13802 VDD.n1471 VDD.n936 146.341
R13803 VDD.n1471 VDD.n928 146.341
R13804 VDD.n1481 VDD.n928 146.341
R13805 VDD.n1481 VDD.n923 146.341
R13806 VDD.n1488 VDD.n923 146.341
R13807 VDD.n1488 VDD.n913 146.341
R13808 VDD.n1525 VDD.n913 146.341
R13809 VDD.n1077 VDD.n1076 146.341
R13810 VDD.n1080 VDD.n1077 146.341
R13811 VDD.n1083 VDD.n1082 146.341
R13812 VDD.n1088 VDD.n1085 146.341
R13813 VDD.n1091 VDD.n1090 146.341
R13814 VDD.n1098 VDD.n1093 146.341
R13815 VDD.n1101 VDD.n1100 146.341
R13816 VDD.n1106 VDD.n1103 146.341
R13817 VDD.n1109 VDD.n1108 146.341
R13818 VDD.n1114 VDD.n1111 146.341
R13819 VDD.n1117 VDD.n1116 146.341
R13820 VDD.n1122 VDD.n1119 146.341
R13821 VDD.n1125 VDD.n1124 146.341
R13822 VDD.n1130 VDD.n1127 146.341
R13823 VDD.n1133 VDD.n1132 146.341
R13824 VDD.n1138 VDD.n1135 146.341
R13825 VDD.n1141 VDD.n1140 146.341
R13826 VDD.n1146 VDD.n1143 146.341
R13827 VDD.n1149 VDD.n1148 146.341
R13828 VDD.n1157 VDD.n1151 146.341
R13829 VDD.n1160 VDD.n1159 146.341
R13830 VDD.n1165 VDD.n1162 146.341
R13831 VDD.n1168 VDD.n1167 146.341
R13832 VDD.n1173 VDD.n1170 146.341
R13833 VDD.n1176 VDD.n1175 146.341
R13834 VDD.n1181 VDD.n1178 146.341
R13835 VDD.n1185 VDD.n1183 146.341
R13836 VDD.n1276 VDD.n1066 146.341
R13837 VDD.n1286 VDD.n1066 146.341
R13838 VDD.n1286 VDD.n1062 146.341
R13839 VDD.n1292 VDD.n1062 146.341
R13840 VDD.n1292 VDD.n1054 146.341
R13841 VDD.n1302 VDD.n1054 146.341
R13842 VDD.n1302 VDD.n1050 146.341
R13843 VDD.n1308 VDD.n1050 146.341
R13844 VDD.n1308 VDD.n1042 146.341
R13845 VDD.n1318 VDD.n1042 146.341
R13846 VDD.n1318 VDD.n1038 146.341
R13847 VDD.n1324 VDD.n1038 146.341
R13848 VDD.n1324 VDD.n1030 146.341
R13849 VDD.n1334 VDD.n1030 146.341
R13850 VDD.n1334 VDD.n1026 146.341
R13851 VDD.n1340 VDD.n1026 146.341
R13852 VDD.n1340 VDD.n1018 146.341
R13853 VDD.n1350 VDD.n1018 146.341
R13854 VDD.n1350 VDD.n1014 146.341
R13855 VDD.n1356 VDD.n1014 146.341
R13856 VDD.n1356 VDD.n1006 146.341
R13857 VDD.n1366 VDD.n1006 146.341
R13858 VDD.n1366 VDD.n1002 146.341
R13859 VDD.n1372 VDD.n1002 146.341
R13860 VDD.n1372 VDD.n994 146.341
R13861 VDD.n1381 VDD.n994 146.341
R13862 VDD.n1381 VDD.n990 146.341
R13863 VDD.n1399 VDD.n990 146.341
R13864 VDD.n1399 VDD.n982 146.341
R13865 VDD.n1409 VDD.n982 146.341
R13866 VDD.n1409 VDD.n978 146.341
R13867 VDD.n1415 VDD.n978 146.341
R13868 VDD.n1415 VDD.n970 146.341
R13869 VDD.n1425 VDD.n970 146.341
R13870 VDD.n1425 VDD.n966 146.341
R13871 VDD.n1431 VDD.n966 146.341
R13872 VDD.n1431 VDD.n958 146.341
R13873 VDD.n1441 VDD.n958 146.341
R13874 VDD.n1441 VDD.n954 146.341
R13875 VDD.n1447 VDD.n954 146.341
R13876 VDD.n1447 VDD.n946 146.341
R13877 VDD.n1457 VDD.n946 146.341
R13878 VDD.n1457 VDD.n942 146.341
R13879 VDD.n1463 VDD.n942 146.341
R13880 VDD.n1463 VDD.n934 146.341
R13881 VDD.n1473 VDD.n934 146.341
R13882 VDD.n1473 VDD.n930 146.341
R13883 VDD.n1479 VDD.n930 146.341
R13884 VDD.n1479 VDD.n921 146.341
R13885 VDD.n1490 VDD.n921 146.341
R13886 VDD.n1490 VDD.n916 146.341
R13887 VDD.n1523 VDD.n916 146.341
R13888 VDD.t32 VDD.t30 120.704
R13889 VDD.t30 VDD.t38 120.704
R13890 VDD.t38 VDD.t48 120.704
R13891 VDD.t42 VDD.t46 120.704
R13892 VDD.t46 VDD.t36 120.704
R13893 VDD.t36 VDD.t24 120.704
R13894 VDD.n1392 VDD.t143 116.591
R13895 VDD.n1389 VDD.t136 116.591
R13896 VDD.n1386 VDD.t8 116.591
R13897 VDD.n1384 VDD.t9 116.591
R13898 VDD.n25 VDD.t133 115.3
R13899 VDD.n22 VDD.t51 115.3
R13900 VDD.n19 VDD.t1 115.3
R13901 VDD.n17 VDD.t145 115.3
R13902 VDD.n1188 VDD.t105 115.114
R13903 VDD.n1155 VDD.t96 115.114
R13904 VDD.n1233 VDD.t90 115.114
R13905 VDD.n1095 VDD.t69 115.114
R13906 VDD.n909 VDD.t73 115.114
R13907 VDD.n779 VDD.t63 115.114
R13908 VDD.n1573 VDD.t66 115.114
R13909 VDD.n729 VDD.t103 115.114
R13910 VDD.n2625 VDD.t59 115.114
R13911 VDD.n177 VDD.t131 115.114
R13912 VDD.n2677 VDD.t115 115.114
R13913 VDD.n123 VDD.t88 115.114
R13914 VDD.n316 VDD.t84 115.114
R13915 VDD.n2395 VDD.t93 115.114
R13916 VDD.n340 VDD.t111 115.114
R13917 VDD.n2365 VDD.t99 115.114
R13918 VDD.n2129 VDD.n1918 113.513
R13919 VDD.n2319 VDD.n2318 99.5127
R13920 VDD.n2316 VDD.n391 99.5127
R13921 VDD.n2312 VDD.n2311 99.5127
R13922 VDD.n2309 VDD.n394 99.5127
R13923 VDD.n2304 VDD.n2303 99.5127
R13924 VDD.n2301 VDD.n397 99.5127
R13925 VDD.n2296 VDD.n2295 99.5127
R13926 VDD.n2096 VDD.n532 99.5127
R13927 VDD.n2093 VDD.n532 99.5127
R13928 VDD.n2093 VDD.n526 99.5127
R13929 VDD.n2090 VDD.n526 99.5127
R13930 VDD.n2090 VDD.n520 99.5127
R13931 VDD.n2087 VDD.n520 99.5127
R13932 VDD.n2087 VDD.n514 99.5127
R13933 VDD.n2084 VDD.n514 99.5127
R13934 VDD.n2084 VDD.n508 99.5127
R13935 VDD.n2081 VDD.n508 99.5127
R13936 VDD.n2081 VDD.n502 99.5127
R13937 VDD.n2078 VDD.n502 99.5127
R13938 VDD.n2078 VDD.n496 99.5127
R13939 VDD.n2075 VDD.n496 99.5127
R13940 VDD.n2075 VDD.n489 99.5127
R13941 VDD.n2072 VDD.n489 99.5127
R13942 VDD.n2072 VDD.n483 99.5127
R13943 VDD.n2069 VDD.n483 99.5127
R13944 VDD.n2069 VDD.n478 99.5127
R13945 VDD.n2066 VDD.n478 99.5127
R13946 VDD.n2066 VDD.n472 99.5127
R13947 VDD.n2063 VDD.n472 99.5127
R13948 VDD.n2063 VDD.n467 99.5127
R13949 VDD.n2060 VDD.n467 99.5127
R13950 VDD.n2060 VDD.n460 99.5127
R13951 VDD.n2057 VDD.n460 99.5127
R13952 VDD.n2057 VDD.n454 99.5127
R13953 VDD.n2054 VDD.n454 99.5127
R13954 VDD.n2054 VDD.n448 99.5127
R13955 VDD.n2051 VDD.n448 99.5127
R13956 VDD.n2051 VDD.n443 99.5127
R13957 VDD.n2048 VDD.n443 99.5127
R13958 VDD.n2048 VDD.n437 99.5127
R13959 VDD.n2045 VDD.n437 99.5127
R13960 VDD.n2045 VDD.n431 99.5127
R13961 VDD.n2042 VDD.n431 99.5127
R13962 VDD.n2042 VDD.n424 99.5127
R13963 VDD.n2039 VDD.n424 99.5127
R13964 VDD.n2039 VDD.n418 99.5127
R13965 VDD.n2036 VDD.n418 99.5127
R13966 VDD.n2036 VDD.n412 99.5127
R13967 VDD.n412 VDD.n404 99.5127
R13968 VDD.n2287 VDD.n404 99.5127
R13969 VDD.n2288 VDD.n2287 99.5127
R13970 VDD.n2288 VDD.n383 99.5127
R13971 VDD.n402 VDD.n383 99.5127
R13972 VDD.n2031 VDD.n2030 99.5127
R13973 VDD.n2122 VDD.n2030 99.5127
R13974 VDD.n2120 VDD.n2119 99.5127
R13975 VDD.n2116 VDD.n2115 99.5127
R13976 VDD.n2112 VDD.n2111 99.5127
R13977 VDD.n2108 VDD.n2107 99.5127
R13978 VDD.n2103 VDD.n2102 99.5127
R13979 VDD.n2099 VDD.n1925 99.5127
R13980 VDD.n2137 VDD.n530 99.5127
R13981 VDD.n2137 VDD.n528 99.5127
R13982 VDD.n2141 VDD.n528 99.5127
R13983 VDD.n2141 VDD.n518 99.5127
R13984 VDD.n2149 VDD.n518 99.5127
R13985 VDD.n2149 VDD.n516 99.5127
R13986 VDD.n2153 VDD.n516 99.5127
R13987 VDD.n2153 VDD.n506 99.5127
R13988 VDD.n2161 VDD.n506 99.5127
R13989 VDD.n2161 VDD.n504 99.5127
R13990 VDD.n2165 VDD.n504 99.5127
R13991 VDD.n2165 VDD.n494 99.5127
R13992 VDD.n2173 VDD.n494 99.5127
R13993 VDD.n2173 VDD.n492 99.5127
R13994 VDD.n2177 VDD.n492 99.5127
R13995 VDD.n2177 VDD.n482 99.5127
R13996 VDD.n2185 VDD.n482 99.5127
R13997 VDD.n2185 VDD.n480 99.5127
R13998 VDD.n2189 VDD.n480 99.5127
R13999 VDD.n2189 VDD.n470 99.5127
R14000 VDD.n2197 VDD.n470 99.5127
R14001 VDD.n2197 VDD.n468 99.5127
R14002 VDD.n2201 VDD.n468 99.5127
R14003 VDD.n2201 VDD.n458 99.5127
R14004 VDD.n2208 VDD.n458 99.5127
R14005 VDD.n2208 VDD.n456 99.5127
R14006 VDD.n2212 VDD.n456 99.5127
R14007 VDD.n2212 VDD.n447 99.5127
R14008 VDD.n2220 VDD.n447 99.5127
R14009 VDD.n2220 VDD.n445 99.5127
R14010 VDD.n2224 VDD.n445 99.5127
R14011 VDD.n2224 VDD.n435 99.5127
R14012 VDD.n2232 VDD.n435 99.5127
R14013 VDD.n2232 VDD.n433 99.5127
R14014 VDD.n2236 VDD.n433 99.5127
R14015 VDD.n2236 VDD.n422 99.5127
R14016 VDD.n2244 VDD.n422 99.5127
R14017 VDD.n2244 VDD.n420 99.5127
R14018 VDD.n2248 VDD.n420 99.5127
R14019 VDD.n2248 VDD.n410 99.5127
R14020 VDD.n2281 VDD.n410 99.5127
R14021 VDD.n2281 VDD.n408 99.5127
R14022 VDD.n2285 VDD.n408 99.5127
R14023 VDD.n2285 VDD.n386 99.5127
R14024 VDD.n2325 VDD.n386 99.5127
R14025 VDD.n2325 VDD.n387 99.5127
R14026 VDD.n1876 VDD.n1875 99.5127
R14027 VDD.n1872 VDD.n1871 99.5127
R14028 VDD.n1868 VDD.n1867 99.5127
R14029 VDD.n1864 VDD.n1863 99.5127
R14030 VDD.n1860 VDD.n1859 99.5127
R14031 VDD.n1856 VDD.n1855 99.5127
R14032 VDD.n1852 VDD.n1851 99.5127
R14033 VDD.n1671 VDD.n699 99.5127
R14034 VDD.n1668 VDD.n699 99.5127
R14035 VDD.n1668 VDD.n693 99.5127
R14036 VDD.n1665 VDD.n693 99.5127
R14037 VDD.n1665 VDD.n686 99.5127
R14038 VDD.n1662 VDD.n686 99.5127
R14039 VDD.n1662 VDD.n680 99.5127
R14040 VDD.n1659 VDD.n680 99.5127
R14041 VDD.n1659 VDD.n675 99.5127
R14042 VDD.n1656 VDD.n675 99.5127
R14043 VDD.n1656 VDD.n669 99.5127
R14044 VDD.n1653 VDD.n669 99.5127
R14045 VDD.n1653 VDD.n663 99.5127
R14046 VDD.n1650 VDD.n663 99.5127
R14047 VDD.n1650 VDD.n657 99.5127
R14048 VDD.n1647 VDD.n657 99.5127
R14049 VDD.n1647 VDD.n651 99.5127
R14050 VDD.n1644 VDD.n651 99.5127
R14051 VDD.n1644 VDD.n645 99.5127
R14052 VDD.n1641 VDD.n645 99.5127
R14053 VDD.n1641 VDD.n640 99.5127
R14054 VDD.n1638 VDD.n640 99.5127
R14055 VDD.n1638 VDD.n635 99.5127
R14056 VDD.n1635 VDD.n635 99.5127
R14057 VDD.n1635 VDD.n628 99.5127
R14058 VDD.n1632 VDD.n628 99.5127
R14059 VDD.n1632 VDD.n622 99.5127
R14060 VDD.n1629 VDD.n622 99.5127
R14061 VDD.n1629 VDD.n616 99.5127
R14062 VDD.n1626 VDD.n616 99.5127
R14063 VDD.n1626 VDD.n610 99.5127
R14064 VDD.n1623 VDD.n610 99.5127
R14065 VDD.n1623 VDD.n604 99.5127
R14066 VDD.n1620 VDD.n604 99.5127
R14067 VDD.n1620 VDD.n598 99.5127
R14068 VDD.n1617 VDD.n598 99.5127
R14069 VDD.n1617 VDD.n591 99.5127
R14070 VDD.n1614 VDD.n591 99.5127
R14071 VDD.n1614 VDD.n584 99.5127
R14072 VDD.n1611 VDD.n584 99.5127
R14073 VDD.n1611 VDD.n578 99.5127
R14074 VDD.n578 VDD.n571 99.5127
R14075 VDD.n1842 VDD.n571 99.5127
R14076 VDD.n1843 VDD.n1842 99.5127
R14077 VDD.n1843 VDD.n562 99.5127
R14078 VDD.n1847 VDD.n562 99.5127
R14079 VDD.n720 VDD.n719 99.5127
R14080 VDD.n1698 VDD.n719 99.5127
R14081 VDD.n1696 VDD.n1695 99.5127
R14082 VDD.n1692 VDD.n1691 99.5127
R14083 VDD.n1687 VDD.n1686 99.5127
R14084 VDD.n1683 VDD.n1682 99.5127
R14085 VDD.n1678 VDD.n1677 99.5127
R14086 VDD.n1674 VDD.n710 99.5127
R14087 VDD.n1712 VDD.n697 99.5127
R14088 VDD.n1712 VDD.n695 99.5127
R14089 VDD.n1716 VDD.n695 99.5127
R14090 VDD.n1716 VDD.n684 99.5127
R14091 VDD.n1724 VDD.n684 99.5127
R14092 VDD.n1724 VDD.n682 99.5127
R14093 VDD.n1728 VDD.n682 99.5127
R14094 VDD.n1728 VDD.n673 99.5127
R14095 VDD.n1736 VDD.n673 99.5127
R14096 VDD.n1736 VDD.n671 99.5127
R14097 VDD.n1740 VDD.n671 99.5127
R14098 VDD.n1740 VDD.n661 99.5127
R14099 VDD.n1748 VDD.n661 99.5127
R14100 VDD.n1748 VDD.n659 99.5127
R14101 VDD.n1752 VDD.n659 99.5127
R14102 VDD.n1752 VDD.n649 99.5127
R14103 VDD.n1760 VDD.n649 99.5127
R14104 VDD.n1760 VDD.n647 99.5127
R14105 VDD.n1764 VDD.n647 99.5127
R14106 VDD.n1764 VDD.n638 99.5127
R14107 VDD.n1772 VDD.n638 99.5127
R14108 VDD.n1772 VDD.n636 99.5127
R14109 VDD.n1776 VDD.n636 99.5127
R14110 VDD.n1776 VDD.n626 99.5127
R14111 VDD.n1783 VDD.n626 99.5127
R14112 VDD.n1783 VDD.n624 99.5127
R14113 VDD.n1787 VDD.n624 99.5127
R14114 VDD.n1787 VDD.n614 99.5127
R14115 VDD.n1795 VDD.n614 99.5127
R14116 VDD.n1795 VDD.n612 99.5127
R14117 VDD.n1799 VDD.n612 99.5127
R14118 VDD.n1799 VDD.n602 99.5127
R14119 VDD.n1807 VDD.n602 99.5127
R14120 VDD.n1807 VDD.n600 99.5127
R14121 VDD.n1811 VDD.n600 99.5127
R14122 VDD.n1811 VDD.n589 99.5127
R14123 VDD.n1819 VDD.n589 99.5127
R14124 VDD.n1819 VDD.n587 99.5127
R14125 VDD.n1823 VDD.n587 99.5127
R14126 VDD.n1823 VDD.n577 99.5127
R14127 VDD.n1836 VDD.n577 99.5127
R14128 VDD.n1836 VDD.n575 99.5127
R14129 VDD.n1840 VDD.n575 99.5127
R14130 VDD.n1840 VDD.n564 99.5127
R14131 VDD.n1882 VDD.n564 99.5127
R14132 VDD.n1882 VDD.n565 99.5127
R14133 VDD.n2268 VDD.n2254 99.5127
R14134 VDD.n2264 VDD.n2263 99.5127
R14135 VDD.n2261 VDD.n2258 99.5127
R14136 VDD.n2344 VDD.n371 99.5127
R14137 VDD.n2342 VDD.n2341 99.5127
R14138 VDD.n2339 VDD.n374 99.5127
R14139 VDD.n2334 VDD.n2333 99.5127
R14140 VDD.n2001 VDD.n533 99.5127
R14141 VDD.n1997 VDD.n533 99.5127
R14142 VDD.n1997 VDD.n527 99.5127
R14143 VDD.n1994 VDD.n527 99.5127
R14144 VDD.n1994 VDD.n521 99.5127
R14145 VDD.n1991 VDD.n521 99.5127
R14146 VDD.n1991 VDD.n515 99.5127
R14147 VDD.n1988 VDD.n515 99.5127
R14148 VDD.n1988 VDD.n509 99.5127
R14149 VDD.n1985 VDD.n509 99.5127
R14150 VDD.n1985 VDD.n503 99.5127
R14151 VDD.n1982 VDD.n503 99.5127
R14152 VDD.n1982 VDD.n497 99.5127
R14153 VDD.n1979 VDD.n497 99.5127
R14154 VDD.n1979 VDD.n490 99.5127
R14155 VDD.n1976 VDD.n490 99.5127
R14156 VDD.n1976 VDD.n484 99.5127
R14157 VDD.n1973 VDD.n484 99.5127
R14158 VDD.n1973 VDD.n479 99.5127
R14159 VDD.n1970 VDD.n479 99.5127
R14160 VDD.n1970 VDD.n473 99.5127
R14161 VDD.n1967 VDD.n473 99.5127
R14162 VDD.n1967 VDD.n466 99.5127
R14163 VDD.n1964 VDD.n466 99.5127
R14164 VDD.n1964 VDD.n461 99.5127
R14165 VDD.n1961 VDD.n461 99.5127
R14166 VDD.n1961 VDD.n455 99.5127
R14167 VDD.n1958 VDD.n455 99.5127
R14168 VDD.n1958 VDD.n449 99.5127
R14169 VDD.n1955 VDD.n449 99.5127
R14170 VDD.n1955 VDD.n444 99.5127
R14171 VDD.n1952 VDD.n444 99.5127
R14172 VDD.n1952 VDD.n438 99.5127
R14173 VDD.n1949 VDD.n438 99.5127
R14174 VDD.n1949 VDD.n432 99.5127
R14175 VDD.n1946 VDD.n432 99.5127
R14176 VDD.n1946 VDD.n425 99.5127
R14177 VDD.n1943 VDD.n425 99.5127
R14178 VDD.n1943 VDD.n419 99.5127
R14179 VDD.n1940 VDD.n419 99.5127
R14180 VDD.n1940 VDD.n413 99.5127
R14181 VDD.n1937 VDD.n413 99.5127
R14182 VDD.n1937 VDD.n406 99.5127
R14183 VDD.n406 VDD.n381 99.5127
R14184 VDD.n2327 VDD.n381 99.5127
R14185 VDD.n2327 VDD.n379 99.5127
R14186 VDD.n2028 VDD.n536 99.5127
R14187 VDD.n2024 VDD.n1932 99.5127
R14188 VDD.n2022 VDD.n2021 99.5127
R14189 VDD.n2018 VDD.n2017 99.5127
R14190 VDD.n2014 VDD.n2013 99.5127
R14191 VDD.n2010 VDD.n2009 99.5127
R14192 VDD.n2006 VDD.n2005 99.5127
R14193 VDD.n2135 VDD.n534 99.5127
R14194 VDD.n2135 VDD.n524 99.5127
R14195 VDD.n2143 VDD.n524 99.5127
R14196 VDD.n2143 VDD.n522 99.5127
R14197 VDD.n2147 VDD.n522 99.5127
R14198 VDD.n2147 VDD.n512 99.5127
R14199 VDD.n2155 VDD.n512 99.5127
R14200 VDD.n2155 VDD.n510 99.5127
R14201 VDD.n2159 VDD.n510 99.5127
R14202 VDD.n2159 VDD.n500 99.5127
R14203 VDD.n2167 VDD.n500 99.5127
R14204 VDD.n2167 VDD.n498 99.5127
R14205 VDD.n2171 VDD.n498 99.5127
R14206 VDD.n2171 VDD.n487 99.5127
R14207 VDD.n2179 VDD.n487 99.5127
R14208 VDD.n2179 VDD.n485 99.5127
R14209 VDD.n2183 VDD.n485 99.5127
R14210 VDD.n2183 VDD.n476 99.5127
R14211 VDD.n2191 VDD.n476 99.5127
R14212 VDD.n2191 VDD.n474 99.5127
R14213 VDD.n2195 VDD.n474 99.5127
R14214 VDD.n2195 VDD.n464 99.5127
R14215 VDD.n2202 VDD.n464 99.5127
R14216 VDD.n2202 VDD.n462 99.5127
R14217 VDD.n2206 VDD.n462 99.5127
R14218 VDD.n2206 VDD.n452 99.5127
R14219 VDD.n2214 VDD.n452 99.5127
R14220 VDD.n2214 VDD.n450 99.5127
R14221 VDD.n2218 VDD.n450 99.5127
R14222 VDD.n2218 VDD.n441 99.5127
R14223 VDD.n2226 VDD.n441 99.5127
R14224 VDD.n2226 VDD.n439 99.5127
R14225 VDD.n2230 VDD.n439 99.5127
R14226 VDD.n2230 VDD.n429 99.5127
R14227 VDD.n2238 VDD.n429 99.5127
R14228 VDD.n2238 VDD.n427 99.5127
R14229 VDD.n2242 VDD.n427 99.5127
R14230 VDD.n2242 VDD.n417 99.5127
R14231 VDD.n2250 VDD.n417 99.5127
R14232 VDD.n2250 VDD.n414 99.5127
R14233 VDD.n2279 VDD.n414 99.5127
R14234 VDD.n2279 VDD.n415 99.5127
R14235 VDD.n415 VDD.n407 99.5127
R14236 VDD.n2274 VDD.n407 99.5127
R14237 VDD.n2274 VDD.n385 99.5127
R14238 VDD.n2271 VDD.n385 99.5127
R14239 VDD.n1917 VDD.n555 99.5127
R14240 VDD.n1913 VDD.n1912 99.5127
R14241 VDD.n1909 VDD.n1908 99.5127
R14242 VDD.n1905 VDD.n1904 99.5127
R14243 VDD.n1901 VDD.n1900 99.5127
R14244 VDD.n1897 VDD.n1896 99.5127
R14245 VDD.n1892 VDD.n1891 99.5127
R14246 VDD.n1888 VDD.n553 99.5127
R14247 VDD.n866 VDD.n700 99.5127
R14248 VDD.n863 VDD.n700 99.5127
R14249 VDD.n863 VDD.n694 99.5127
R14250 VDD.n860 VDD.n694 99.5127
R14251 VDD.n860 VDD.n687 99.5127
R14252 VDD.n857 VDD.n687 99.5127
R14253 VDD.n857 VDD.n681 99.5127
R14254 VDD.n854 VDD.n681 99.5127
R14255 VDD.n854 VDD.n676 99.5127
R14256 VDD.n851 VDD.n676 99.5127
R14257 VDD.n851 VDD.n670 99.5127
R14258 VDD.n848 VDD.n670 99.5127
R14259 VDD.n848 VDD.n664 99.5127
R14260 VDD.n845 VDD.n664 99.5127
R14261 VDD.n845 VDD.n658 99.5127
R14262 VDD.n842 VDD.n658 99.5127
R14263 VDD.n842 VDD.n652 99.5127
R14264 VDD.n839 VDD.n652 99.5127
R14265 VDD.n839 VDD.n646 99.5127
R14266 VDD.n836 VDD.n646 99.5127
R14267 VDD.n836 VDD.n641 99.5127
R14268 VDD.n833 VDD.n641 99.5127
R14269 VDD.n833 VDD.n634 99.5127
R14270 VDD.n830 VDD.n634 99.5127
R14271 VDD.n830 VDD.n629 99.5127
R14272 VDD.n827 VDD.n629 99.5127
R14273 VDD.n827 VDD.n623 99.5127
R14274 VDD.n824 VDD.n623 99.5127
R14275 VDD.n824 VDD.n617 99.5127
R14276 VDD.n821 VDD.n617 99.5127
R14277 VDD.n821 VDD.n611 99.5127
R14278 VDD.n818 VDD.n611 99.5127
R14279 VDD.n818 VDD.n605 99.5127
R14280 VDD.n815 VDD.n605 99.5127
R14281 VDD.n815 VDD.n599 99.5127
R14282 VDD.n812 VDD.n599 99.5127
R14283 VDD.n812 VDD.n592 99.5127
R14284 VDD.n809 VDD.n592 99.5127
R14285 VDD.n809 VDD.n585 99.5127
R14286 VDD.n806 VDD.n585 99.5127
R14287 VDD.n806 VDD.n579 99.5127
R14288 VDD.n803 VDD.n579 99.5127
R14289 VDD.n803 VDD.n573 99.5127
R14290 VDD.n573 VDD.n560 99.5127
R14291 VDD.n1884 VDD.n560 99.5127
R14292 VDD.n1885 VDD.n1884 99.5127
R14293 VDD.n1706 VDD.n703 99.5127
R14294 VDD.n789 VDD.n788 99.5127
R14295 VDD.n793 VDD.n792 99.5127
R14296 VDD.n797 VDD.n796 99.5127
R14297 VDD.n882 VDD.n881 99.5127
R14298 VDD.n878 VDD.n877 99.5127
R14299 VDD.n873 VDD.n872 99.5127
R14300 VDD.n869 VDD.n718 99.5127
R14301 VDD.n1710 VDD.n701 99.5127
R14302 VDD.n1710 VDD.n691 99.5127
R14303 VDD.n1718 VDD.n691 99.5127
R14304 VDD.n1718 VDD.n689 99.5127
R14305 VDD.n1722 VDD.n689 99.5127
R14306 VDD.n1722 VDD.n679 99.5127
R14307 VDD.n1730 VDD.n679 99.5127
R14308 VDD.n1730 VDD.n677 99.5127
R14309 VDD.n1734 VDD.n677 99.5127
R14310 VDD.n1734 VDD.n667 99.5127
R14311 VDD.n1742 VDD.n667 99.5127
R14312 VDD.n1742 VDD.n665 99.5127
R14313 VDD.n1746 VDD.n665 99.5127
R14314 VDD.n1746 VDD.n655 99.5127
R14315 VDD.n1754 VDD.n655 99.5127
R14316 VDD.n1754 VDD.n653 99.5127
R14317 VDD.n1758 VDD.n653 99.5127
R14318 VDD.n1758 VDD.n644 99.5127
R14319 VDD.n1766 VDD.n644 99.5127
R14320 VDD.n1766 VDD.n642 99.5127
R14321 VDD.n1770 VDD.n642 99.5127
R14322 VDD.n1770 VDD.n632 99.5127
R14323 VDD.n1777 VDD.n632 99.5127
R14324 VDD.n1777 VDD.n630 99.5127
R14325 VDD.n1781 VDD.n630 99.5127
R14326 VDD.n1781 VDD.n620 99.5127
R14327 VDD.n1789 VDD.n620 99.5127
R14328 VDD.n1789 VDD.n618 99.5127
R14329 VDD.n1793 VDD.n618 99.5127
R14330 VDD.n1793 VDD.n608 99.5127
R14331 VDD.n1801 VDD.n608 99.5127
R14332 VDD.n1801 VDD.n606 99.5127
R14333 VDD.n1805 VDD.n606 99.5127
R14334 VDD.n1805 VDD.n596 99.5127
R14335 VDD.n1813 VDD.n596 99.5127
R14336 VDD.n1813 VDD.n594 99.5127
R14337 VDD.n1817 VDD.n594 99.5127
R14338 VDD.n1817 VDD.n583 99.5127
R14339 VDD.n1825 VDD.n583 99.5127
R14340 VDD.n1825 VDD.n580 99.5127
R14341 VDD.n1834 VDD.n580 99.5127
R14342 VDD.n1834 VDD.n581 99.5127
R14343 VDD.n581 VDD.n574 99.5127
R14344 VDD.n1829 VDD.n574 99.5127
R14345 VDD.n1829 VDD.n563 99.5127
R14346 VDD.n563 VDD.n554 99.5127
R14347 VDD.n25 VDD.n24 98.4825
R14348 VDD.n22 VDD.n21 98.4825
R14349 VDD.n19 VDD.n18 98.4825
R14350 VDD.n17 VDD.n16 98.4825
R14351 VDD.n1392 VDD.n1391 97.1923
R14352 VDD.n1389 VDD.n1388 97.1923
R14353 VDD.n1386 VDD.n1385 97.1923
R14354 VDD.n1384 VDD.n1383 97.1923
R14355 VDD.n1705 VDD.t48 89.5907
R14356 VDD.n372 VDD.t42 89.5907
R14357 VDD.n1188 VDD.n1187 74.2793
R14358 VDD.n1155 VDD.n1154 74.2793
R14359 VDD.n1233 VDD.n1232 74.2793
R14360 VDD.n1095 VDD.n1094 74.2793
R14361 VDD.n909 VDD.n908 74.2793
R14362 VDD.n779 VDD.n778 74.2793
R14363 VDD.n1573 VDD.n1572 74.2793
R14364 VDD.n729 VDD.n728 74.2793
R14365 VDD.n2625 VDD.n2624 74.2793
R14366 VDD.n177 VDD.n176 74.2793
R14367 VDD.n2677 VDD.n2676 74.2793
R14368 VDD.n123 VDD.n122 74.2793
R14369 VDD.n316 VDD.n315 74.2793
R14370 VDD.n2395 VDD.n2394 74.2793
R14371 VDD.n340 VDD.n339 74.2793
R14372 VDD.n2365 VDD.n2364 74.2793
R14373 VDD.n2130 VDD.n2129 72.8958
R14374 VDD.n2129 VDD.n2029 72.8958
R14375 VDD.n2129 VDD.n1931 72.8958
R14376 VDD.n2129 VDD.n1930 72.8958
R14377 VDD.n2129 VDD.n1929 72.8958
R14378 VDD.n2129 VDD.n1928 72.8958
R14379 VDD.n2129 VDD.n1927 72.8958
R14380 VDD.n2129 VDD.n1926 72.8958
R14381 VDD.n2332 VDD.n372 72.8958
R14382 VDD.n378 VDD.n372 72.8958
R14383 VDD.n2340 VDD.n372 72.8958
R14384 VDD.n2343 VDD.n372 72.8958
R14385 VDD.n2257 VDD.n372 72.8958
R14386 VDD.n2262 VDD.n372 72.8958
R14387 VDD.n2256 VDD.n372 72.8958
R14388 VDD.n2269 VDD.n372 72.8958
R14389 VDD.n1705 VDD.n1704 72.8958
R14390 VDD.n1705 VDD.n704 72.8958
R14391 VDD.n1705 VDD.n705 72.8958
R14392 VDD.n1705 VDD.n706 72.8958
R14393 VDD.n1705 VDD.n707 72.8958
R14394 VDD.n1705 VDD.n708 72.8958
R14395 VDD.n1705 VDD.n709 72.8958
R14396 VDD.n1918 VDD.n545 72.8958
R14397 VDD.n1918 VDD.n544 72.8958
R14398 VDD.n1918 VDD.n543 72.8958
R14399 VDD.n1918 VDD.n542 72.8958
R14400 VDD.n1918 VDD.n541 72.8958
R14401 VDD.n1918 VDD.n540 72.8958
R14402 VDD.n1918 VDD.n539 72.8958
R14403 VDD.n1918 VDD.n538 72.8958
R14404 VDD.n2129 VDD.n2128 72.8958
R14405 VDD.n2129 VDD.n1919 72.8958
R14406 VDD.n2129 VDD.n1920 72.8958
R14407 VDD.n2129 VDD.n1921 72.8958
R14408 VDD.n2129 VDD.n1922 72.8958
R14409 VDD.n2129 VDD.n1923 72.8958
R14410 VDD.n2129 VDD.n1924 72.8958
R14411 VDD.n2294 VDD.n372 72.8958
R14412 VDD.n401 VDD.n372 72.8958
R14413 VDD.n2302 VDD.n372 72.8958
R14414 VDD.n396 VDD.n372 72.8958
R14415 VDD.n2310 VDD.n372 72.8958
R14416 VDD.n393 VDD.n372 72.8958
R14417 VDD.n2317 VDD.n372 72.8958
R14418 VDD.n2320 VDD.n372 72.8958
R14419 VDD.n1918 VDD.n552 72.8958
R14420 VDD.n1918 VDD.n551 72.8958
R14421 VDD.n1918 VDD.n550 72.8958
R14422 VDD.n1918 VDD.n549 72.8958
R14423 VDD.n1918 VDD.n548 72.8958
R14424 VDD.n1918 VDD.n547 72.8958
R14425 VDD.n1918 VDD.n546 72.8958
R14426 VDD.n1705 VDD.n711 72.8958
R14427 VDD.n1705 VDD.n712 72.8958
R14428 VDD.n1705 VDD.n713 72.8958
R14429 VDD.n1705 VDD.n714 72.8958
R14430 VDD.n1705 VDD.n715 72.8958
R14431 VDD.n1705 VDD.n716 72.8958
R14432 VDD.n1705 VDD.n717 72.8958
R14433 VDD.n1075 VDD.n1072 66.2847
R14434 VDD.n1081 VDD.n1072 66.2847
R14435 VDD.n1084 VDD.n1072 66.2847
R14436 VDD.n1089 VDD.n1072 66.2847
R14437 VDD.n1092 VDD.n1072 66.2847
R14438 VDD.n1099 VDD.n1072 66.2847
R14439 VDD.n1102 VDD.n1072 66.2847
R14440 VDD.n1107 VDD.n1072 66.2847
R14441 VDD.n1110 VDD.n1072 66.2847
R14442 VDD.n1115 VDD.n1072 66.2847
R14443 VDD.n1118 VDD.n1072 66.2847
R14444 VDD.n1123 VDD.n1072 66.2847
R14445 VDD.n1126 VDD.n1072 66.2847
R14446 VDD.n1131 VDD.n1072 66.2847
R14447 VDD.n1134 VDD.n1072 66.2847
R14448 VDD.n1139 VDD.n1072 66.2847
R14449 VDD.n1142 VDD.n1072 66.2847
R14450 VDD.n1147 VDD.n1072 66.2847
R14451 VDD.n1150 VDD.n1072 66.2847
R14452 VDD.n1158 VDD.n1072 66.2847
R14453 VDD.n1161 VDD.n1072 66.2847
R14454 VDD.n1166 VDD.n1072 66.2847
R14455 VDD.n1169 VDD.n1072 66.2847
R14456 VDD.n1174 VDD.n1072 66.2847
R14457 VDD.n1177 VDD.n1072 66.2847
R14458 VDD.n1182 VDD.n1072 66.2847
R14459 VDD.n1184 VDD.n1072 66.2847
R14460 VDD.n912 VDD.n727 66.2847
R14461 VDD.n904 VDD.n727 66.2847
R14462 VDD.n901 VDD.n727 66.2847
R14463 VDD.n896 VDD.n727 66.2847
R14464 VDD.n893 VDD.n727 66.2847
R14465 VDD.n889 VDD.n727 66.2847
R14466 VDD.n784 VDD.n727 66.2847
R14467 VDD.n1547 VDD.n727 66.2847
R14468 VDD.n776 VDD.n727 66.2847
R14469 VDD.n1554 VDD.n727 66.2847
R14470 VDD.n769 VDD.n727 66.2847
R14471 VDD.n1561 VDD.n727 66.2847
R14472 VDD.n762 VDD.n727 66.2847
R14473 VDD.n1568 VDD.n727 66.2847
R14474 VDD.n755 VDD.n727 66.2847
R14475 VDD.n1578 VDD.n727 66.2847
R14476 VDD.n748 VDD.n727 66.2847
R14477 VDD.n1585 VDD.n727 66.2847
R14478 VDD.n741 VDD.n727 66.2847
R14479 VDD.n1592 VDD.n727 66.2847
R14480 VDD.n734 VDD.n727 66.2847
R14481 VDD.n1599 VDD.n727 66.2847
R14482 VDD.n1602 VDD.n727 66.2847
R14483 VDD.n1506 VDD.n727 66.2847
R14484 VDD.n1505 VDD.n727 66.2847
R14485 VDD.n1513 VDD.n727 66.2847
R14486 VDD.n1516 VDD.n727 66.2847
R14487 VDD.n2470 VDD.n298 66.2847
R14488 VDD.n302 VDD.n298 66.2847
R14489 VDD.n2463 VDD.n298 66.2847
R14490 VDD.n2457 VDD.n298 66.2847
R14491 VDD.n2455 VDD.n298 66.2847
R14492 VDD.n317 VDD.n298 66.2847
R14493 VDD.n2447 VDD.n298 66.2847
R14494 VDD.n321 VDD.n298 66.2847
R14495 VDD.n2440 VDD.n298 66.2847
R14496 VDD.n2434 VDD.n298 66.2847
R14497 VDD.n2432 VDD.n298 66.2847
R14498 VDD.n2426 VDD.n298 66.2847
R14499 VDD.n2424 VDD.n298 66.2847
R14500 VDD.n2418 VDD.n298 66.2847
R14501 VDD.n2416 VDD.n298 66.2847
R14502 VDD.n2410 VDD.n298 66.2847
R14503 VDD.n2408 VDD.n298 66.2847
R14504 VDD.n2402 VDD.n298 66.2847
R14505 VDD.n2400 VDD.n298 66.2847
R14506 VDD.n2391 VDD.n298 66.2847
R14507 VDD.n2389 VDD.n298 66.2847
R14508 VDD.n2348 VDD.n298 66.2847
R14509 VDD.n2380 VDD.n298 66.2847
R14510 VDD.n2378 VDD.n298 66.2847
R14511 VDD.n2372 VDD.n298 66.2847
R14512 VDD.n2370 VDD.n298 66.2847
R14513 VDD.n2358 VDD.n298 66.2847
R14514 VDD.n2621 VDD.n102 66.2847
R14515 VDD.n2630 VDD.n102 66.2847
R14516 VDD.n198 VDD.n102 66.2847
R14517 VDD.n2637 VDD.n102 66.2847
R14518 VDD.n191 VDD.n102 66.2847
R14519 VDD.n2644 VDD.n102 66.2847
R14520 VDD.n184 VDD.n102 66.2847
R14521 VDD.n2651 VDD.n102 66.2847
R14522 VDD.n174 VDD.n102 66.2847
R14523 VDD.n2658 VDD.n102 66.2847
R14524 VDD.n167 VDD.n102 66.2847
R14525 VDD.n2665 VDD.n102 66.2847
R14526 VDD.n160 VDD.n102 66.2847
R14527 VDD.n2672 VDD.n102 66.2847
R14528 VDD.n153 VDD.n102 66.2847
R14529 VDD.n2682 VDD.n102 66.2847
R14530 VDD.n146 VDD.n102 66.2847
R14531 VDD.n2689 VDD.n102 66.2847
R14532 VDD.n139 VDD.n102 66.2847
R14533 VDD.n2696 VDD.n102 66.2847
R14534 VDD.n132 VDD.n102 66.2847
R14535 VDD.n2703 VDD.n102 66.2847
R14536 VDD.n125 VDD.n102 66.2847
R14537 VDD.n2710 VDD.n102 66.2847
R14538 VDD.n116 VDD.n102 66.2847
R14539 VDD.n2717 VDD.n102 66.2847
R14540 VDD.n109 VDD.n102 66.2847
R14541 VDD.n800 VDD.n799 62.0611
R14542 VDD.n558 VDD.n557 62.0611
R14543 VDD.n1608 VDD.n1607 62.0611
R14544 VDD.n568 VDD.n567 62.0611
R14545 VDD.n1934 VDD.n1933 62.0611
R14546 VDD.n399 VDD.n398 62.0611
R14547 VDD.n2033 VDD.n2032 62.0611
R14548 VDD.n376 VDD.n375 62.0611
R14549 VDD.n2719 VDD.n109 52.4337
R14550 VDD.n2717 VDD.n2716 52.4337
R14551 VDD.n2712 VDD.n116 52.4337
R14552 VDD.n2710 VDD.n2709 52.4337
R14553 VDD.n2705 VDD.n125 52.4337
R14554 VDD.n2703 VDD.n2702 52.4337
R14555 VDD.n2698 VDD.n132 52.4337
R14556 VDD.n2696 VDD.n2695 52.4337
R14557 VDD.n2691 VDD.n139 52.4337
R14558 VDD.n2689 VDD.n2688 52.4337
R14559 VDD.n2684 VDD.n146 52.4337
R14560 VDD.n2682 VDD.n2681 52.4337
R14561 VDD.n2674 VDD.n153 52.4337
R14562 VDD.n2672 VDD.n2671 52.4337
R14563 VDD.n2667 VDD.n160 52.4337
R14564 VDD.n2665 VDD.n2664 52.4337
R14565 VDD.n2660 VDD.n167 52.4337
R14566 VDD.n2658 VDD.n2657 52.4337
R14567 VDD.n2653 VDD.n174 52.4337
R14568 VDD.n2651 VDD.n2650 52.4337
R14569 VDD.n2646 VDD.n184 52.4337
R14570 VDD.n2644 VDD.n2643 52.4337
R14571 VDD.n2639 VDD.n191 52.4337
R14572 VDD.n2637 VDD.n2636 52.4337
R14573 VDD.n2632 VDD.n198 52.4337
R14574 VDD.n2630 VDD.n2629 52.4337
R14575 VDD.n2622 VDD.n2621 52.4337
R14576 VDD.n2470 VDD.n299 52.4337
R14577 VDD.n2468 VDD.n302 52.4337
R14578 VDD.n2464 VDD.n2463 52.4337
R14579 VDD.n2457 VDD.n307 52.4337
R14580 VDD.n2456 VDD.n2455 52.4337
R14581 VDD.n317 VDD.n313 52.4337
R14582 VDD.n2448 VDD.n2447 52.4337
R14583 VDD.n2445 VDD.n321 52.4337
R14584 VDD.n2441 VDD.n2440 52.4337
R14585 VDD.n2434 VDD.n326 52.4337
R14586 VDD.n2433 VDD.n2432 52.4337
R14587 VDD.n2426 VDD.n332 52.4337
R14588 VDD.n2425 VDD.n2424 52.4337
R14589 VDD.n2418 VDD.n338 52.4337
R14590 VDD.n2417 VDD.n2416 52.4337
R14591 VDD.n2410 VDD.n347 52.4337
R14592 VDD.n2409 VDD.n2408 52.4337
R14593 VDD.n2402 VDD.n353 52.4337
R14594 VDD.n2401 VDD.n2400 52.4337
R14595 VDD.n2391 VDD.n359 52.4337
R14596 VDD.n2390 VDD.n2389 52.4337
R14597 VDD.n2348 VDD.n365 52.4337
R14598 VDD.n2380 VDD.n2350 52.4337
R14599 VDD.n2379 VDD.n2378 52.4337
R14600 VDD.n2372 VDD.n2352 52.4337
R14601 VDD.n2371 VDD.n2370 52.4337
R14602 VDD.n2359 VDD.n2358 52.4337
R14603 VDD.n1516 VDD.n1515 52.4337
R14604 VDD.n1513 VDD.n1512 52.4337
R14605 VDD.n1508 VDD.n1505 52.4337
R14606 VDD.n1506 VDD.n726 52.4337
R14607 VDD.n1602 VDD.n1601 52.4337
R14608 VDD.n1599 VDD.n1598 52.4337
R14609 VDD.n1594 VDD.n734 52.4337
R14610 VDD.n1592 VDD.n1591 52.4337
R14611 VDD.n1587 VDD.n741 52.4337
R14612 VDD.n1585 VDD.n1584 52.4337
R14613 VDD.n1580 VDD.n748 52.4337
R14614 VDD.n1578 VDD.n1577 52.4337
R14615 VDD.n1570 VDD.n755 52.4337
R14616 VDD.n1568 VDD.n1567 52.4337
R14617 VDD.n1563 VDD.n762 52.4337
R14618 VDD.n1561 VDD.n1560 52.4337
R14619 VDD.n1556 VDD.n769 52.4337
R14620 VDD.n1554 VDD.n1553 52.4337
R14621 VDD.n1549 VDD.n776 52.4337
R14622 VDD.n1547 VDD.n1546 52.4337
R14623 VDD.n785 VDD.n784 52.4337
R14624 VDD.n891 VDD.n889 52.4337
R14625 VDD.n894 VDD.n893 52.4337
R14626 VDD.n897 VDD.n896 52.4337
R14627 VDD.n902 VDD.n901 52.4337
R14628 VDD.n905 VDD.n904 52.4337
R14629 VDD.n1526 VDD.n912 52.4337
R14630 VDD.n1075 VDD.n1073 52.4337
R14631 VDD.n1081 VDD.n1080 52.4337
R14632 VDD.n1084 VDD.n1083 52.4337
R14633 VDD.n1089 VDD.n1088 52.4337
R14634 VDD.n1092 VDD.n1091 52.4337
R14635 VDD.n1099 VDD.n1098 52.4337
R14636 VDD.n1102 VDD.n1101 52.4337
R14637 VDD.n1107 VDD.n1106 52.4337
R14638 VDD.n1110 VDD.n1109 52.4337
R14639 VDD.n1115 VDD.n1114 52.4337
R14640 VDD.n1118 VDD.n1117 52.4337
R14641 VDD.n1123 VDD.n1122 52.4337
R14642 VDD.n1126 VDD.n1125 52.4337
R14643 VDD.n1131 VDD.n1130 52.4337
R14644 VDD.n1134 VDD.n1133 52.4337
R14645 VDD.n1139 VDD.n1138 52.4337
R14646 VDD.n1142 VDD.n1141 52.4337
R14647 VDD.n1147 VDD.n1146 52.4337
R14648 VDD.n1150 VDD.n1149 52.4337
R14649 VDD.n1158 VDD.n1157 52.4337
R14650 VDD.n1161 VDD.n1160 52.4337
R14651 VDD.n1166 VDD.n1165 52.4337
R14652 VDD.n1169 VDD.n1168 52.4337
R14653 VDD.n1174 VDD.n1173 52.4337
R14654 VDD.n1177 VDD.n1176 52.4337
R14655 VDD.n1182 VDD.n1181 52.4337
R14656 VDD.n1185 VDD.n1184 52.4337
R14657 VDD.n1076 VDD.n1075 52.4337
R14658 VDD.n1082 VDD.n1081 52.4337
R14659 VDD.n1085 VDD.n1084 52.4337
R14660 VDD.n1090 VDD.n1089 52.4337
R14661 VDD.n1093 VDD.n1092 52.4337
R14662 VDD.n1100 VDD.n1099 52.4337
R14663 VDD.n1103 VDD.n1102 52.4337
R14664 VDD.n1108 VDD.n1107 52.4337
R14665 VDD.n1111 VDD.n1110 52.4337
R14666 VDD.n1116 VDD.n1115 52.4337
R14667 VDD.n1119 VDD.n1118 52.4337
R14668 VDD.n1124 VDD.n1123 52.4337
R14669 VDD.n1127 VDD.n1126 52.4337
R14670 VDD.n1132 VDD.n1131 52.4337
R14671 VDD.n1135 VDD.n1134 52.4337
R14672 VDD.n1140 VDD.n1139 52.4337
R14673 VDD.n1143 VDD.n1142 52.4337
R14674 VDD.n1148 VDD.n1147 52.4337
R14675 VDD.n1151 VDD.n1150 52.4337
R14676 VDD.n1159 VDD.n1158 52.4337
R14677 VDD.n1162 VDD.n1161 52.4337
R14678 VDD.n1167 VDD.n1166 52.4337
R14679 VDD.n1170 VDD.n1169 52.4337
R14680 VDD.n1175 VDD.n1174 52.4337
R14681 VDD.n1178 VDD.n1177 52.4337
R14682 VDD.n1183 VDD.n1182 52.4337
R14683 VDD.n1184 VDD.n1071 52.4337
R14684 VDD.n912 VDD.n911 52.4337
R14685 VDD.n904 VDD.n903 52.4337
R14686 VDD.n901 VDD.n900 52.4337
R14687 VDD.n896 VDD.n895 52.4337
R14688 VDD.n893 VDD.n892 52.4337
R14689 VDD.n889 VDD.n888 52.4337
R14690 VDD.n784 VDD.n777 52.4337
R14691 VDD.n1548 VDD.n1547 52.4337
R14692 VDD.n776 VDD.n770 52.4337
R14693 VDD.n1555 VDD.n1554 52.4337
R14694 VDD.n769 VDD.n763 52.4337
R14695 VDD.n1562 VDD.n1561 52.4337
R14696 VDD.n762 VDD.n756 52.4337
R14697 VDD.n1569 VDD.n1568 52.4337
R14698 VDD.n755 VDD.n749 52.4337
R14699 VDD.n1579 VDD.n1578 52.4337
R14700 VDD.n748 VDD.n742 52.4337
R14701 VDD.n1586 VDD.n1585 52.4337
R14702 VDD.n741 VDD.n735 52.4337
R14703 VDD.n1593 VDD.n1592 52.4337
R14704 VDD.n734 VDD.n731 52.4337
R14705 VDD.n1600 VDD.n1599 52.4337
R14706 VDD.n1603 VDD.n1602 52.4337
R14707 VDD.n1507 VDD.n1506 52.4337
R14708 VDD.n1505 VDD.n1497 52.4337
R14709 VDD.n1514 VDD.n1513 52.4337
R14710 VDD.n1517 VDD.n1516 52.4337
R14711 VDD.n2471 VDD.n2470 52.4337
R14712 VDD.n2465 VDD.n302 52.4337
R14713 VDD.n2463 VDD.n2462 52.4337
R14714 VDD.n2458 VDD.n2457 52.4337
R14715 VDD.n2455 VDD.n2454 52.4337
R14716 VDD.n318 VDD.n317 52.4337
R14717 VDD.n2447 VDD.n2446 52.4337
R14718 VDD.n2442 VDD.n321 52.4337
R14719 VDD.n2440 VDD.n2439 52.4337
R14720 VDD.n2435 VDD.n2434 52.4337
R14721 VDD.n2432 VDD.n2431 52.4337
R14722 VDD.n2427 VDD.n2426 52.4337
R14723 VDD.n2424 VDD.n2423 52.4337
R14724 VDD.n2419 VDD.n2418 52.4337
R14725 VDD.n2416 VDD.n2415 52.4337
R14726 VDD.n2411 VDD.n2410 52.4337
R14727 VDD.n2408 VDD.n2407 52.4337
R14728 VDD.n2403 VDD.n2402 52.4337
R14729 VDD.n2400 VDD.n2399 52.4337
R14730 VDD.n2392 VDD.n2391 52.4337
R14731 VDD.n2389 VDD.n2388 52.4337
R14732 VDD.n2349 VDD.n2348 52.4337
R14733 VDD.n2381 VDD.n2380 52.4337
R14734 VDD.n2378 VDD.n2377 52.4337
R14735 VDD.n2373 VDD.n2372 52.4337
R14736 VDD.n2370 VDD.n2369 52.4337
R14737 VDD.n2358 VDD.n297 52.4337
R14738 VDD.n2621 VDD.n199 52.4337
R14739 VDD.n2631 VDD.n2630 52.4337
R14740 VDD.n198 VDD.n192 52.4337
R14741 VDD.n2638 VDD.n2637 52.4337
R14742 VDD.n191 VDD.n185 52.4337
R14743 VDD.n2645 VDD.n2644 52.4337
R14744 VDD.n184 VDD.n175 52.4337
R14745 VDD.n2652 VDD.n2651 52.4337
R14746 VDD.n174 VDD.n168 52.4337
R14747 VDD.n2659 VDD.n2658 52.4337
R14748 VDD.n167 VDD.n161 52.4337
R14749 VDD.n2666 VDD.n2665 52.4337
R14750 VDD.n160 VDD.n154 52.4337
R14751 VDD.n2673 VDD.n2672 52.4337
R14752 VDD.n153 VDD.n147 52.4337
R14753 VDD.n2683 VDD.n2682 52.4337
R14754 VDD.n146 VDD.n140 52.4337
R14755 VDD.n2690 VDD.n2689 52.4337
R14756 VDD.n139 VDD.n133 52.4337
R14757 VDD.n2697 VDD.n2696 52.4337
R14758 VDD.n132 VDD.n126 52.4337
R14759 VDD.n2704 VDD.n2703 52.4337
R14760 VDD.n125 VDD.n117 52.4337
R14761 VDD.n2711 VDD.n2710 52.4337
R14762 VDD.n116 VDD.n110 52.4337
R14763 VDD.n2718 VDD.n2717 52.4337
R14764 VDD.n109 VDD.n106 52.4337
R14765 VDD.n2320 VDD.n2319 39.2114
R14766 VDD.n2317 VDD.n2316 39.2114
R14767 VDD.n2312 VDD.n393 39.2114
R14768 VDD.n2310 VDD.n2309 39.2114
R14769 VDD.n2304 VDD.n396 39.2114
R14770 VDD.n2302 VDD.n2301 39.2114
R14771 VDD.n2296 VDD.n401 39.2114
R14772 VDD.n2294 VDD.n2293 39.2114
R14773 VDD.n2128 VDD.n2127 39.2114
R14774 VDD.n2122 VDD.n1919 39.2114
R14775 VDD.n2119 VDD.n1920 39.2114
R14776 VDD.n2115 VDD.n1921 39.2114
R14777 VDD.n2111 VDD.n1922 39.2114
R14778 VDD.n2107 VDD.n1923 39.2114
R14779 VDD.n2102 VDD.n1924 39.2114
R14780 VDD.n1876 VDD.n538 39.2114
R14781 VDD.n1872 VDD.n539 39.2114
R14782 VDD.n1868 VDD.n540 39.2114
R14783 VDD.n1864 VDD.n541 39.2114
R14784 VDD.n1860 VDD.n542 39.2114
R14785 VDD.n1856 VDD.n543 39.2114
R14786 VDD.n1852 VDD.n544 39.2114
R14787 VDD.n1848 VDD.n545 39.2114
R14788 VDD.n1704 VDD.n1703 39.2114
R14789 VDD.n1698 VDD.n704 39.2114
R14790 VDD.n1695 VDD.n705 39.2114
R14791 VDD.n1691 VDD.n706 39.2114
R14792 VDD.n1686 VDD.n707 39.2114
R14793 VDD.n1682 VDD.n708 39.2114
R14794 VDD.n1677 VDD.n709 39.2114
R14795 VDD.n2269 VDD.n2268 39.2114
R14796 VDD.n2264 VDD.n2256 39.2114
R14797 VDD.n2262 VDD.n2261 39.2114
R14798 VDD.n2257 VDD.n371 39.2114
R14799 VDD.n2343 VDD.n2342 39.2114
R14800 VDD.n2340 VDD.n2339 39.2114
R14801 VDD.n2334 VDD.n378 39.2114
R14802 VDD.n2332 VDD.n2331 39.2114
R14803 VDD.n2131 VDD.n2130 39.2114
R14804 VDD.n2029 VDD.n2028 39.2114
R14805 VDD.n2024 VDD.n1931 39.2114
R14806 VDD.n2021 VDD.n1930 39.2114
R14807 VDD.n2017 VDD.n1929 39.2114
R14808 VDD.n2013 VDD.n1928 39.2114
R14809 VDD.n2009 VDD.n1927 39.2114
R14810 VDD.n2005 VDD.n1926 39.2114
R14811 VDD.n2130 VDD.n536 39.2114
R14812 VDD.n2029 VDD.n1932 39.2114
R14813 VDD.n2022 VDD.n1931 39.2114
R14814 VDD.n2018 VDD.n1930 39.2114
R14815 VDD.n2014 VDD.n1929 39.2114
R14816 VDD.n2010 VDD.n1928 39.2114
R14817 VDD.n2006 VDD.n1927 39.2114
R14818 VDD.n2002 VDD.n1926 39.2114
R14819 VDD.n2333 VDD.n2332 39.2114
R14820 VDD.n378 VDD.n374 39.2114
R14821 VDD.n2341 VDD.n2340 39.2114
R14822 VDD.n2344 VDD.n2343 39.2114
R14823 VDD.n2258 VDD.n2257 39.2114
R14824 VDD.n2263 VDD.n2262 39.2114
R14825 VDD.n2256 VDD.n2254 39.2114
R14826 VDD.n2270 VDD.n2269 39.2114
R14827 VDD.n1704 VDD.n720 39.2114
R14828 VDD.n1696 VDD.n704 39.2114
R14829 VDD.n1692 VDD.n705 39.2114
R14830 VDD.n1687 VDD.n706 39.2114
R14831 VDD.n1683 VDD.n707 39.2114
R14832 VDD.n1678 VDD.n708 39.2114
R14833 VDD.n1674 VDD.n709 39.2114
R14834 VDD.n1851 VDD.n545 39.2114
R14835 VDD.n1855 VDD.n544 39.2114
R14836 VDD.n1859 VDD.n543 39.2114
R14837 VDD.n1863 VDD.n542 39.2114
R14838 VDD.n1867 VDD.n541 39.2114
R14839 VDD.n1871 VDD.n540 39.2114
R14840 VDD.n1875 VDD.n539 39.2114
R14841 VDD.n1878 VDD.n538 39.2114
R14842 VDD.n2128 VDD.n2031 39.2114
R14843 VDD.n2120 VDD.n1919 39.2114
R14844 VDD.n2116 VDD.n1920 39.2114
R14845 VDD.n2112 VDD.n1921 39.2114
R14846 VDD.n2108 VDD.n1922 39.2114
R14847 VDD.n2103 VDD.n1923 39.2114
R14848 VDD.n2099 VDD.n1924 39.2114
R14849 VDD.n2295 VDD.n2294 39.2114
R14850 VDD.n401 VDD.n397 39.2114
R14851 VDD.n2303 VDD.n2302 39.2114
R14852 VDD.n396 VDD.n394 39.2114
R14853 VDD.n2311 VDD.n2310 39.2114
R14854 VDD.n393 VDD.n391 39.2114
R14855 VDD.n2318 VDD.n2317 39.2114
R14856 VDD.n2321 VDD.n2320 39.2114
R14857 VDD.n555 VDD.n546 39.2114
R14858 VDD.n1912 VDD.n547 39.2114
R14859 VDD.n1908 VDD.n548 39.2114
R14860 VDD.n1904 VDD.n549 39.2114
R14861 VDD.n1900 VDD.n550 39.2114
R14862 VDD.n1896 VDD.n551 39.2114
R14863 VDD.n1891 VDD.n552 39.2114
R14864 VDD.n711 VDD.n703 39.2114
R14865 VDD.n789 VDD.n712 39.2114
R14866 VDD.n793 VDD.n713 39.2114
R14867 VDD.n797 VDD.n714 39.2114
R14868 VDD.n881 VDD.n715 39.2114
R14869 VDD.n877 VDD.n716 39.2114
R14870 VDD.n872 VDD.n717 39.2114
R14871 VDD.n1888 VDD.n552 39.2114
R14872 VDD.n1892 VDD.n551 39.2114
R14873 VDD.n1897 VDD.n550 39.2114
R14874 VDD.n1901 VDD.n549 39.2114
R14875 VDD.n1905 VDD.n548 39.2114
R14876 VDD.n1909 VDD.n547 39.2114
R14877 VDD.n1913 VDD.n546 39.2114
R14878 VDD.n788 VDD.n711 39.2114
R14879 VDD.n792 VDD.n712 39.2114
R14880 VDD.n796 VDD.n713 39.2114
R14881 VDD.n882 VDD.n714 39.2114
R14882 VDD.n878 VDD.n715 39.2114
R14883 VDD.n873 VDD.n716 39.2114
R14884 VDD.n869 VDD.n717 39.2114
R14885 VDD.n1880 VDD.n1879 32.3127
R14886 VDD.n1849 VDD.n1846 32.3127
R14887 VDD.n1673 VDD.n1672 32.3127
R14888 VDD.n1702 VDD.n696 32.3127
R14889 VDD.n2098 VDD.n2097 32.3127
R14890 VDD.n2292 VDD.n2291 32.3127
R14891 VDD.n2126 VDD.n529 32.3127
R14892 VDD.n2323 VDD.n2322 32.3127
R14893 VDD.n2272 VDD.n2253 32.3127
R14894 VDD.n2330 VDD.n2329 32.3127
R14895 VDD.n2003 VDD.n2000 32.3127
R14896 VDD.n2133 VDD.n2132 32.3127
R14897 VDD.n1708 VDD.n1707 32.3127
R14898 VDD.n1916 VDD.n556 32.3127
R14899 VDD.n1887 VDD.n1886 32.3127
R14900 VDD.n868 VDD.n867 32.3127
R14901 VDD.n1189 VDD.n1188 30.8369
R14902 VDD.n1156 VDD.n1155 30.8369
R14903 VDD.n1234 VDD.n1233 30.8369
R14904 VDD.n1096 VDD.n1095 30.8369
R14905 VDD.n910 VDD.n909 30.8369
R14906 VDD.n780 VDD.n779 30.8369
R14907 VDD.n1574 VDD.n1573 30.8369
R14908 VDD.n730 VDD.n729 30.8369
R14909 VDD.n2626 VDD.n2625 30.8369
R14910 VDD.n178 VDD.n177 30.8369
R14911 VDD.n2678 VDD.n2677 30.8369
R14912 VDD.n124 VDD.n123 30.8369
R14913 VDD.n2451 VDD.n316 30.8369
R14914 VDD.n2396 VDD.n2395 30.8369
R14915 VDD.n341 VDD.n340 30.8369
R14916 VDD.n2366 VDD.n2365 30.8369
R14917 VDD.n7 VDD.t37 29.6854
R14918 VDD.n7 VDD.t25 29.6854
R14919 VDD.n8 VDD.t43 29.6854
R14920 VDD.n8 VDD.t47 29.6854
R14921 VDD.n10 VDD.t20 29.6854
R14922 VDD.n10 VDD.t45 29.6854
R14923 VDD.n12 VDD.t35 29.6854
R14924 VDD.n12 VDD.t22 29.6854
R14925 VDD.n5 VDD.t29 29.6854
R14926 VDD.n5 VDD.t27 29.6854
R14927 VDD.n3 VDD.t41 29.6854
R14928 VDD.n3 VDD.t18 29.6854
R14929 VDD.n1 VDD.t39 29.6854
R14930 VDD.n1 VDD.t49 29.6854
R14931 VDD.n0 VDD.t33 29.6854
R14932 VDD.n0 VDD.t31 29.6854
R14933 VDD.n1277 VDD.n1072 24.0788
R14934 VDD.n1524 VDD.n727 24.0788
R14935 VDD.n2478 VDD.n298 24.0788
R14936 VDD.n2727 VDD.n102 24.0788
R14937 VDD.n875 VDD.n800 24.049
R14938 VDD.n1894 VDD.n558 24.049
R14939 VDD.n1680 VDD.n1608 24.049
R14940 VDD.n569 VDD.n568 24.049
R14941 VDD.n1935 VDD.n1934 24.049
R14942 VDD.n2299 VDD.n399 24.049
R14943 VDD.n2105 VDD.n2033 24.049
R14944 VDD.n2337 VDD.n376 24.049
R14945 VDD.n1279 VDD.n1069 19.3944
R14946 VDD.n1283 VDD.n1069 19.3944
R14947 VDD.n1283 VDD.n1058 19.3944
R14948 VDD.n1295 VDD.n1058 19.3944
R14949 VDD.n1295 VDD.n1056 19.3944
R14950 VDD.n1299 VDD.n1056 19.3944
R14951 VDD.n1299 VDD.n1047 19.3944
R14952 VDD.n1311 VDD.n1047 19.3944
R14953 VDD.n1311 VDD.n1045 19.3944
R14954 VDD.n1315 VDD.n1045 19.3944
R14955 VDD.n1315 VDD.n1035 19.3944
R14956 VDD.n1327 VDD.n1035 19.3944
R14957 VDD.n1327 VDD.n1033 19.3944
R14958 VDD.n1331 VDD.n1033 19.3944
R14959 VDD.n1331 VDD.n1022 19.3944
R14960 VDD.n1343 VDD.n1022 19.3944
R14961 VDD.n1343 VDD.n1020 19.3944
R14962 VDD.n1347 VDD.n1020 19.3944
R14963 VDD.n1347 VDD.n1011 19.3944
R14964 VDD.n1359 VDD.n1011 19.3944
R14965 VDD.n1359 VDD.n1009 19.3944
R14966 VDD.n1363 VDD.n1009 19.3944
R14967 VDD.n1363 VDD.n999 19.3944
R14968 VDD.n1375 VDD.n999 19.3944
R14969 VDD.n1375 VDD.n997 19.3944
R14970 VDD.n1379 VDD.n997 19.3944
R14971 VDD.n1379 VDD.n987 19.3944
R14972 VDD.n1402 VDD.n987 19.3944
R14973 VDD.n1402 VDD.n985 19.3944
R14974 VDD.n1406 VDD.n985 19.3944
R14975 VDD.n1406 VDD.n975 19.3944
R14976 VDD.n1418 VDD.n975 19.3944
R14977 VDD.n1418 VDD.n973 19.3944
R14978 VDD.n1422 VDD.n973 19.3944
R14979 VDD.n1422 VDD.n963 19.3944
R14980 VDD.n1434 VDD.n963 19.3944
R14981 VDD.n1434 VDD.n961 19.3944
R14982 VDD.n1438 VDD.n961 19.3944
R14983 VDD.n1438 VDD.n951 19.3944
R14984 VDD.n1450 VDD.n951 19.3944
R14985 VDD.n1450 VDD.n949 19.3944
R14986 VDD.n1454 VDD.n949 19.3944
R14987 VDD.n1454 VDD.n939 19.3944
R14988 VDD.n1466 VDD.n939 19.3944
R14989 VDD.n1466 VDD.n937 19.3944
R14990 VDD.n1470 VDD.n937 19.3944
R14991 VDD.n1470 VDD.n927 19.3944
R14992 VDD.n1482 VDD.n927 19.3944
R14993 VDD.n1482 VDD.n924 19.3944
R14994 VDD.n1487 VDD.n924 19.3944
R14995 VDD.n1487 VDD.n925 19.3944
R14996 VDD.n925 VDD.n914 19.3944
R14997 VDD.n1209 VDD.n1208 19.3944
R14998 VDD.n1208 VDD.n1207 19.3944
R14999 VDD.n1207 VDD.n1163 19.3944
R15000 VDD.n1203 VDD.n1163 19.3944
R15001 VDD.n1203 VDD.n1202 19.3944
R15002 VDD.n1202 VDD.n1201 19.3944
R15003 VDD.n1201 VDD.n1171 19.3944
R15004 VDD.n1197 VDD.n1171 19.3944
R15005 VDD.n1197 VDD.n1196 19.3944
R15006 VDD.n1196 VDD.n1195 19.3944
R15007 VDD.n1195 VDD.n1179 19.3944
R15008 VDD.n1191 VDD.n1179 19.3944
R15009 VDD.n1191 VDD.n1190 19.3944
R15010 VDD.n1231 VDD.n1128 19.3944
R15011 VDD.n1227 VDD.n1128 19.3944
R15012 VDD.n1227 VDD.n1226 19.3944
R15013 VDD.n1226 VDD.n1225 19.3944
R15014 VDD.n1225 VDD.n1136 19.3944
R15015 VDD.n1221 VDD.n1136 19.3944
R15016 VDD.n1221 VDD.n1220 19.3944
R15017 VDD.n1220 VDD.n1219 19.3944
R15018 VDD.n1219 VDD.n1144 19.3944
R15019 VDD.n1215 VDD.n1144 19.3944
R15020 VDD.n1215 VDD.n1214 19.3944
R15021 VDD.n1214 VDD.n1213 19.3944
R15022 VDD.n1213 VDD.n1152 19.3944
R15023 VDD.n1254 VDD.n1253 19.3944
R15024 VDD.n1253 VDD.n1252 19.3944
R15025 VDD.n1252 VDD.n1104 19.3944
R15026 VDD.n1248 VDD.n1104 19.3944
R15027 VDD.n1248 VDD.n1247 19.3944
R15028 VDD.n1247 VDD.n1246 19.3944
R15029 VDD.n1246 VDD.n1112 19.3944
R15030 VDD.n1242 VDD.n1112 19.3944
R15031 VDD.n1242 VDD.n1241 19.3944
R15032 VDD.n1241 VDD.n1240 19.3944
R15033 VDD.n1240 VDD.n1120 19.3944
R15034 VDD.n1236 VDD.n1120 19.3944
R15035 VDD.n1236 VDD.n1235 19.3944
R15036 VDD.n1272 VDD.n1271 19.3944
R15037 VDD.n1271 VDD.n1270 19.3944
R15038 VDD.n1270 VDD.n1078 19.3944
R15039 VDD.n1266 VDD.n1078 19.3944
R15040 VDD.n1266 VDD.n1265 19.3944
R15041 VDD.n1265 VDD.n1264 19.3944
R15042 VDD.n1264 VDD.n1086 19.3944
R15043 VDD.n1260 VDD.n1086 19.3944
R15044 VDD.n1260 VDD.n1259 19.3944
R15045 VDD.n1259 VDD.n1258 19.3944
R15046 VDD.n1275 VDD.n1065 19.3944
R15047 VDD.n1287 VDD.n1065 19.3944
R15048 VDD.n1287 VDD.n1063 19.3944
R15049 VDD.n1291 VDD.n1063 19.3944
R15050 VDD.n1291 VDD.n1053 19.3944
R15051 VDD.n1303 VDD.n1053 19.3944
R15052 VDD.n1303 VDD.n1051 19.3944
R15053 VDD.n1307 VDD.n1051 19.3944
R15054 VDD.n1307 VDD.n1041 19.3944
R15055 VDD.n1319 VDD.n1041 19.3944
R15056 VDD.n1319 VDD.n1039 19.3944
R15057 VDD.n1323 VDD.n1039 19.3944
R15058 VDD.n1323 VDD.n1029 19.3944
R15059 VDD.n1335 VDD.n1029 19.3944
R15060 VDD.n1335 VDD.n1027 19.3944
R15061 VDD.n1339 VDD.n1027 19.3944
R15062 VDD.n1339 VDD.n1017 19.3944
R15063 VDD.n1351 VDD.n1017 19.3944
R15064 VDD.n1351 VDD.n1015 19.3944
R15065 VDD.n1355 VDD.n1015 19.3944
R15066 VDD.n1355 VDD.n1005 19.3944
R15067 VDD.n1367 VDD.n1005 19.3944
R15068 VDD.n1367 VDD.n1003 19.3944
R15069 VDD.n1371 VDD.n1003 19.3944
R15070 VDD.n1371 VDD.n993 19.3944
R15071 VDD.n1382 VDD.n993 19.3944
R15072 VDD.n1382 VDD.n991 19.3944
R15073 VDD.n1398 VDD.n991 19.3944
R15074 VDD.n1398 VDD.n981 19.3944
R15075 VDD.n1410 VDD.n981 19.3944
R15076 VDD.n1410 VDD.n979 19.3944
R15077 VDD.n1414 VDD.n979 19.3944
R15078 VDD.n1414 VDD.n969 19.3944
R15079 VDD.n1426 VDD.n969 19.3944
R15080 VDD.n1426 VDD.n967 19.3944
R15081 VDD.n1430 VDD.n967 19.3944
R15082 VDD.n1430 VDD.n957 19.3944
R15083 VDD.n1442 VDD.n957 19.3944
R15084 VDD.n1442 VDD.n955 19.3944
R15085 VDD.n1446 VDD.n955 19.3944
R15086 VDD.n1446 VDD.n945 19.3944
R15087 VDD.n1458 VDD.n945 19.3944
R15088 VDD.n1458 VDD.n943 19.3944
R15089 VDD.n1462 VDD.n943 19.3944
R15090 VDD.n1462 VDD.n933 19.3944
R15091 VDD.n1474 VDD.n933 19.3944
R15092 VDD.n1474 VDD.n931 19.3944
R15093 VDD.n1478 VDD.n931 19.3944
R15094 VDD.n1478 VDD.n920 19.3944
R15095 VDD.n1491 VDD.n920 19.3944
R15096 VDD.n1491 VDD.n918 19.3944
R15097 VDD.n1522 VDD.n918 19.3944
R15098 VDD.n1545 VDD.n1544 19.3944
R15099 VDD.n1544 VDD.n1543 19.3944
R15100 VDD.n890 VDD.n786 19.3944
R15101 VDD.n1539 VDD.n887 19.3944
R15102 VDD.n1539 VDD.n1538 19.3944
R15103 VDD.n1538 VDD.n1537 19.3944
R15104 VDD.n1537 VDD.n898 19.3944
R15105 VDD.n1533 VDD.n898 19.3944
R15106 VDD.n1533 VDD.n1532 19.3944
R15107 VDD.n1532 VDD.n1531 19.3944
R15108 VDD.n1531 VDD.n906 19.3944
R15109 VDD.n1571 VDD.n754 19.3944
R15110 VDD.n1566 VDD.n754 19.3944
R15111 VDD.n1566 VDD.n1565 19.3944
R15112 VDD.n1565 VDD.n1564 19.3944
R15113 VDD.n1564 VDD.n761 19.3944
R15114 VDD.n1559 VDD.n761 19.3944
R15115 VDD.n1559 VDD.n1558 19.3944
R15116 VDD.n1558 VDD.n1557 19.3944
R15117 VDD.n1557 VDD.n768 19.3944
R15118 VDD.n1552 VDD.n768 19.3944
R15119 VDD.n1552 VDD.n1551 19.3944
R15120 VDD.n1551 VDD.n1550 19.3944
R15121 VDD.n1550 VDD.n775 19.3944
R15122 VDD.n1597 VDD.n1596 19.3944
R15123 VDD.n1596 VDD.n1595 19.3944
R15124 VDD.n1595 VDD.n733 19.3944
R15125 VDD.n1590 VDD.n733 19.3944
R15126 VDD.n1590 VDD.n1589 19.3944
R15127 VDD.n1589 VDD.n1588 19.3944
R15128 VDD.n1588 VDD.n740 19.3944
R15129 VDD.n1583 VDD.n740 19.3944
R15130 VDD.n1583 VDD.n1582 19.3944
R15131 VDD.n1582 VDD.n1581 19.3944
R15132 VDD.n1581 VDD.n747 19.3944
R15133 VDD.n1576 VDD.n747 19.3944
R15134 VDD.n1576 VDD.n1575 19.3944
R15135 VDD.n1519 VDD.n1518 19.3944
R15136 VDD.n1518 VDD.n1495 19.3944
R15137 VDD.n1496 VDD.n1495 19.3944
R15138 VDD.n1511 VDD.n1496 19.3944
R15139 VDD.n1511 VDD.n1510 19.3944
R15140 VDD.n1510 VDD.n1509 19.3944
R15141 VDD.n1509 VDD.n1504 19.3944
R15142 VDD.n1504 VDD.n725 19.3944
R15143 VDD.n1604 VDD.n725 19.3944
R15144 VDD.n2480 VDD.n295 19.3944
R15145 VDD.n2484 VDD.n295 19.3944
R15146 VDD.n2484 VDD.n284 19.3944
R15147 VDD.n2496 VDD.n284 19.3944
R15148 VDD.n2496 VDD.n282 19.3944
R15149 VDD.n2500 VDD.n282 19.3944
R15150 VDD.n2500 VDD.n273 19.3944
R15151 VDD.n2512 VDD.n273 19.3944
R15152 VDD.n2512 VDD.n271 19.3944
R15153 VDD.n2516 VDD.n271 19.3944
R15154 VDD.n2516 VDD.n261 19.3944
R15155 VDD.n2528 VDD.n261 19.3944
R15156 VDD.n2528 VDD.n259 19.3944
R15157 VDD.n2532 VDD.n259 19.3944
R15158 VDD.n2532 VDD.n248 19.3944
R15159 VDD.n2544 VDD.n248 19.3944
R15160 VDD.n2544 VDD.n246 19.3944
R15161 VDD.n2548 VDD.n246 19.3944
R15162 VDD.n2548 VDD.n237 19.3944
R15163 VDD.n2560 VDD.n237 19.3944
R15164 VDD.n2560 VDD.n235 19.3944
R15165 VDD.n2564 VDD.n235 19.3944
R15166 VDD.n2564 VDD.n224 19.3944
R15167 VDD.n2576 VDD.n224 19.3944
R15168 VDD.n2576 VDD.n222 19.3944
R15169 VDD.n2580 VDD.n222 19.3944
R15170 VDD.n2581 VDD.n2580 19.3944
R15171 VDD.n2582 VDD.n2581 19.3944
R15172 VDD.n2582 VDD.n220 19.3944
R15173 VDD.n2586 VDD.n220 19.3944
R15174 VDD.n2587 VDD.n2586 19.3944
R15175 VDD.n2588 VDD.n2587 19.3944
R15176 VDD.n2588 VDD.n217 19.3944
R15177 VDD.n2592 VDD.n217 19.3944
R15178 VDD.n2593 VDD.n2592 19.3944
R15179 VDD.n2594 VDD.n2593 19.3944
R15180 VDD.n2594 VDD.n214 19.3944
R15181 VDD.n2598 VDD.n214 19.3944
R15182 VDD.n2599 VDD.n2598 19.3944
R15183 VDD.n2600 VDD.n2599 19.3944
R15184 VDD.n2600 VDD.n211 19.3944
R15185 VDD.n2604 VDD.n211 19.3944
R15186 VDD.n2605 VDD.n2604 19.3944
R15187 VDD.n2606 VDD.n2605 19.3944
R15188 VDD.n2606 VDD.n208 19.3944
R15189 VDD.n2610 VDD.n208 19.3944
R15190 VDD.n2611 VDD.n2610 19.3944
R15191 VDD.n2612 VDD.n2611 19.3944
R15192 VDD.n2612 VDD.n205 19.3944
R15193 VDD.n2616 VDD.n205 19.3944
R15194 VDD.n2617 VDD.n2616 19.3944
R15195 VDD.n2618 VDD.n2617 19.3944
R15196 VDD.n2649 VDD.n2648 19.3944
R15197 VDD.n2648 VDD.n2647 19.3944
R15198 VDD.n2647 VDD.n183 19.3944
R15199 VDD.n2642 VDD.n183 19.3944
R15200 VDD.n2642 VDD.n2641 19.3944
R15201 VDD.n2641 VDD.n2640 19.3944
R15202 VDD.n2640 VDD.n190 19.3944
R15203 VDD.n2635 VDD.n190 19.3944
R15204 VDD.n2635 VDD.n2634 19.3944
R15205 VDD.n2634 VDD.n2633 19.3944
R15206 VDD.n2633 VDD.n197 19.3944
R15207 VDD.n2628 VDD.n197 19.3944
R15208 VDD.n2628 VDD.n2627 19.3944
R15209 VDD.n2675 VDD.n152 19.3944
R15210 VDD.n2670 VDD.n152 19.3944
R15211 VDD.n2670 VDD.n2669 19.3944
R15212 VDD.n2669 VDD.n2668 19.3944
R15213 VDD.n2668 VDD.n159 19.3944
R15214 VDD.n2663 VDD.n159 19.3944
R15215 VDD.n2663 VDD.n2662 19.3944
R15216 VDD.n2662 VDD.n2661 19.3944
R15217 VDD.n2661 VDD.n166 19.3944
R15218 VDD.n2656 VDD.n166 19.3944
R15219 VDD.n2656 VDD.n2655 19.3944
R15220 VDD.n2655 VDD.n2654 19.3944
R15221 VDD.n2654 VDD.n173 19.3944
R15222 VDD.n2701 VDD.n2700 19.3944
R15223 VDD.n2700 VDD.n2699 19.3944
R15224 VDD.n2699 VDD.n131 19.3944
R15225 VDD.n2694 VDD.n131 19.3944
R15226 VDD.n2694 VDD.n2693 19.3944
R15227 VDD.n2693 VDD.n2692 19.3944
R15228 VDD.n2692 VDD.n138 19.3944
R15229 VDD.n2687 VDD.n138 19.3944
R15230 VDD.n2687 VDD.n2686 19.3944
R15231 VDD.n2686 VDD.n2685 19.3944
R15232 VDD.n2685 VDD.n145 19.3944
R15233 VDD.n2680 VDD.n145 19.3944
R15234 VDD.n2680 VDD.n2679 19.3944
R15235 VDD.n2722 VDD.n2721 19.3944
R15236 VDD.n2721 VDD.n2720 19.3944
R15237 VDD.n2720 VDD.n108 19.3944
R15238 VDD.n2715 VDD.n108 19.3944
R15239 VDD.n2715 VDD.n2714 19.3944
R15240 VDD.n2714 VDD.n2713 19.3944
R15241 VDD.n2713 VDD.n115 19.3944
R15242 VDD.n2708 VDD.n115 19.3944
R15243 VDD.n2708 VDD.n2707 19.3944
R15244 VDD.n2707 VDD.n2706 19.3944
R15245 VDD.n2476 VDD.n291 19.3944
R15246 VDD.n2488 VDD.n291 19.3944
R15247 VDD.n2488 VDD.n289 19.3944
R15248 VDD.n2492 VDD.n289 19.3944
R15249 VDD.n2492 VDD.n279 19.3944
R15250 VDD.n2504 VDD.n279 19.3944
R15251 VDD.n2504 VDD.n277 19.3944
R15252 VDD.n2508 VDD.n277 19.3944
R15253 VDD.n2508 VDD.n267 19.3944
R15254 VDD.n2520 VDD.n267 19.3944
R15255 VDD.n2520 VDD.n265 19.3944
R15256 VDD.n2524 VDD.n265 19.3944
R15257 VDD.n2524 VDD.n255 19.3944
R15258 VDD.n2536 VDD.n255 19.3944
R15259 VDD.n2536 VDD.n253 19.3944
R15260 VDD.n2540 VDD.n253 19.3944
R15261 VDD.n2540 VDD.n243 19.3944
R15262 VDD.n2552 VDD.n243 19.3944
R15263 VDD.n2552 VDD.n241 19.3944
R15264 VDD.n2556 VDD.n241 19.3944
R15265 VDD.n2556 VDD.n231 19.3944
R15266 VDD.n2568 VDD.n231 19.3944
R15267 VDD.n2568 VDD.n229 19.3944
R15268 VDD.n2572 VDD.n229 19.3944
R15269 VDD.n2572 VDD.n29 19.3944
R15270 VDD.n2778 VDD.n29 19.3944
R15271 VDD.n2778 VDD.n30 19.3944
R15272 VDD.n2773 VDD.n30 19.3944
R15273 VDD.n2773 VDD.n2772 19.3944
R15274 VDD.n2772 VDD.n2771 19.3944
R15275 VDD.n2771 VDD.n42 19.3944
R15276 VDD.n2765 VDD.n42 19.3944
R15277 VDD.n2765 VDD.n2764 19.3944
R15278 VDD.n2764 VDD.n2763 19.3944
R15279 VDD.n2763 VDD.n53 19.3944
R15280 VDD.n2757 VDD.n53 19.3944
R15281 VDD.n2757 VDD.n2756 19.3944
R15282 VDD.n2756 VDD.n2755 19.3944
R15283 VDD.n2755 VDD.n64 19.3944
R15284 VDD.n2749 VDD.n64 19.3944
R15285 VDD.n2749 VDD.n2748 19.3944
R15286 VDD.n2748 VDD.n2747 19.3944
R15287 VDD.n2747 VDD.n75 19.3944
R15288 VDD.n2741 VDD.n75 19.3944
R15289 VDD.n2741 VDD.n2740 19.3944
R15290 VDD.n2740 VDD.n2739 19.3944
R15291 VDD.n2739 VDD.n86 19.3944
R15292 VDD.n2733 VDD.n86 19.3944
R15293 VDD.n2733 VDD.n2732 19.3944
R15294 VDD.n2732 VDD.n2731 19.3944
R15295 VDD.n2731 VDD.n97 19.3944
R15296 VDD.n2725 VDD.n97 19.3944
R15297 VDD.n2473 VDD.n2472 19.3944
R15298 VDD.n2472 VDD.n301 19.3944
R15299 VDD.n2467 VDD.n301 19.3944
R15300 VDD.n2467 VDD.n2466 19.3944
R15301 VDD.n2466 VDD.n306 19.3944
R15302 VDD.n2461 VDD.n306 19.3944
R15303 VDD.n2461 VDD.n2460 19.3944
R15304 VDD.n2460 VDD.n2459 19.3944
R15305 VDD.n2459 VDD.n312 19.3944
R15306 VDD.n2453 VDD.n312 19.3944
R15307 VDD.n2422 VDD.n2421 19.3944
R15308 VDD.n2421 VDD.n2420 19.3944
R15309 VDD.n2420 VDD.n346 19.3944
R15310 VDD.n2414 VDD.n346 19.3944
R15311 VDD.n2414 VDD.n2413 19.3944
R15312 VDD.n2413 VDD.n2412 19.3944
R15313 VDD.n2412 VDD.n352 19.3944
R15314 VDD.n2406 VDD.n352 19.3944
R15315 VDD.n2406 VDD.n2405 19.3944
R15316 VDD.n2405 VDD.n2404 19.3944
R15317 VDD.n2404 VDD.n358 19.3944
R15318 VDD.n2398 VDD.n358 19.3944
R15319 VDD.n2398 VDD.n2397 19.3944
R15320 VDD.n2450 VDD.n2449 19.3944
R15321 VDD.n2449 VDD.n320 19.3944
R15322 VDD.n2444 VDD.n320 19.3944
R15323 VDD.n2444 VDD.n2443 19.3944
R15324 VDD.n2443 VDD.n325 19.3944
R15325 VDD.n2438 VDD.n325 19.3944
R15326 VDD.n2438 VDD.n2437 19.3944
R15327 VDD.n2437 VDD.n2436 19.3944
R15328 VDD.n2436 VDD.n331 19.3944
R15329 VDD.n2430 VDD.n331 19.3944
R15330 VDD.n2430 VDD.n2429 19.3944
R15331 VDD.n2429 VDD.n2428 19.3944
R15332 VDD.n2428 VDD.n337 19.3944
R15333 VDD.n2393 VDD.n364 19.3944
R15334 VDD.n2387 VDD.n364 19.3944
R15335 VDD.n2347 VDD.n366 19.3944
R15336 VDD.n2383 VDD.n2382 19.3944
R15337 VDD.n2382 VDD.n2351 19.3944
R15338 VDD.n2376 VDD.n2351 19.3944
R15339 VDD.n2376 VDD.n2375 19.3944
R15340 VDD.n2375 VDD.n2374 19.3944
R15341 VDD.n2374 VDD.n2357 19.3944
R15342 VDD.n2368 VDD.n2357 19.3944
R15343 VDD.n2368 VDD.n2367 19.3944
R15344 VDD.n1258 VDD.n1096 18.8126
R15345 VDD.n730 VDD.n724 18.8126
R15346 VDD.n2706 VDD.n124 18.8126
R15347 VDD.n24 VDD.t141 18.1091
R15348 VDD.n24 VDD.t10 18.1091
R15349 VDD.n21 VDD.t139 18.1091
R15350 VDD.n21 VDD.t11 18.1091
R15351 VDD.n18 VDD.t138 18.1091
R15352 VDD.n18 VDD.t3 18.1091
R15353 VDD.n16 VDD.t142 18.1091
R15354 VDD.n16 VDD.t6 18.1091
R15355 VDD.n1391 VDD.t14 18.1091
R15356 VDD.n1391 VDD.t134 18.1091
R15357 VDD.n1388 VDD.t135 18.1091
R15358 VDD.n1388 VDD.t50 18.1091
R15359 VDD.n1385 VDD.t5 18.1091
R15360 VDD.n1385 VDD.t144 18.1091
R15361 VDD.n1383 VDD.t132 18.1091
R15362 VDD.n1383 VDD.t13 18.1091
R15363 VDD.n1705 VDD.n698 17.043
R15364 VDD.n1918 VDD.n537 17.043
R15365 VDD.n2129 VDD.n531 17.043
R15366 VDD.n384 VDD.n372 17.043
R15367 VDD.n1277 VDD.n1067 15.6358
R15368 VDD.n1285 VDD.n1067 15.6358
R15369 VDD.n1285 VDD.n1060 15.6358
R15370 VDD.n1293 VDD.n1060 15.6358
R15371 VDD.n1293 VDD.n1061 15.6358
R15372 VDD.n1301 VDD.n1049 15.6358
R15373 VDD.n1309 VDD.n1049 15.6358
R15374 VDD.n1309 VDD.n1043 15.6358
R15375 VDD.n1317 VDD.n1043 15.6358
R15376 VDD.n1317 VDD.n1037 15.6358
R15377 VDD.n1325 VDD.n1037 15.6358
R15378 VDD.n1325 VDD.n1031 15.6358
R15379 VDD.n1333 VDD.n1031 15.6358
R15380 VDD.n1333 VDD.n1024 15.6358
R15381 VDD.n1341 VDD.n1024 15.6358
R15382 VDD.n1341 VDD.n1025 15.6358
R15383 VDD.n1349 VDD.n1013 15.6358
R15384 VDD.n1357 VDD.n1013 15.6358
R15385 VDD.n1357 VDD.n1007 15.6358
R15386 VDD.n1365 VDD.n1007 15.6358
R15387 VDD.n1365 VDD.n1001 15.6358
R15388 VDD.n1373 VDD.n1001 15.6358
R15389 VDD.n1373 VDD.n995 15.6358
R15390 VDD.t12 VDD.n995 15.6358
R15391 VDD.t12 VDD.n989 15.6358
R15392 VDD.n1400 VDD.n989 15.6358
R15393 VDD.n1400 VDD.n983 15.6358
R15394 VDD.n1408 VDD.n983 15.6358
R15395 VDD.n1408 VDD.n977 15.6358
R15396 VDD.n1416 VDD.n977 15.6358
R15397 VDD.n1416 VDD.n971 15.6358
R15398 VDD.n1424 VDD.n971 15.6358
R15399 VDD.n1432 VDD.n965 15.6358
R15400 VDD.n1432 VDD.n959 15.6358
R15401 VDD.n1440 VDD.n959 15.6358
R15402 VDD.n1440 VDD.n953 15.6358
R15403 VDD.n1448 VDD.n953 15.6358
R15404 VDD.n1448 VDD.n947 15.6358
R15405 VDD.n1456 VDD.n947 15.6358
R15406 VDD.n1456 VDD.n941 15.6358
R15407 VDD.n1464 VDD.n941 15.6358
R15408 VDD.n1464 VDD.n935 15.6358
R15409 VDD.n1472 VDD.n935 15.6358
R15410 VDD.n1480 VDD.n929 15.6358
R15411 VDD.n1480 VDD.n922 15.6358
R15412 VDD.n1489 VDD.n922 15.6358
R15413 VDD.n1489 VDD.n915 15.6358
R15414 VDD.n1524 VDD.n915 15.6358
R15415 VDD.n2478 VDD.n293 15.6358
R15416 VDD.n2486 VDD.n293 15.6358
R15417 VDD.n2486 VDD.n286 15.6358
R15418 VDD.n2494 VDD.n286 15.6358
R15419 VDD.n2494 VDD.n287 15.6358
R15420 VDD.n2502 VDD.n275 15.6358
R15421 VDD.n2510 VDD.n275 15.6358
R15422 VDD.n2510 VDD.n269 15.6358
R15423 VDD.n2518 VDD.n269 15.6358
R15424 VDD.n2518 VDD.n263 15.6358
R15425 VDD.n2526 VDD.n263 15.6358
R15426 VDD.n2526 VDD.n257 15.6358
R15427 VDD.n2534 VDD.n257 15.6358
R15428 VDD.n2534 VDD.n250 15.6358
R15429 VDD.n2542 VDD.n250 15.6358
R15430 VDD.n2542 VDD.n251 15.6358
R15431 VDD.n2550 VDD.n239 15.6358
R15432 VDD.n2558 VDD.n239 15.6358
R15433 VDD.n2558 VDD.n233 15.6358
R15434 VDD.n2566 VDD.n233 15.6358
R15435 VDD.n2566 VDD.n227 15.6358
R15436 VDD.n2574 VDD.n227 15.6358
R15437 VDD.n2574 VDD.n33 15.6358
R15438 VDD.t2 VDD.n33 15.6358
R15439 VDD.t2 VDD.n2776 15.6358
R15440 VDD.n2776 VDD.n2775 15.6358
R15441 VDD.n2775 VDD.n37 15.6358
R15442 VDD.n2769 VDD.n37 15.6358
R15443 VDD.n2769 VDD.n2768 15.6358
R15444 VDD.n2768 VDD.n2767 15.6358
R15445 VDD.n2767 VDD.n47 15.6358
R15446 VDD.n2761 VDD.n47 15.6358
R15447 VDD.n2760 VDD.n2759 15.6358
R15448 VDD.n2759 VDD.n58 15.6358
R15449 VDD.n2753 VDD.n58 15.6358
R15450 VDD.n2753 VDD.n2752 15.6358
R15451 VDD.n2752 VDD.n2751 15.6358
R15452 VDD.n2751 VDD.n69 15.6358
R15453 VDD.n2745 VDD.n69 15.6358
R15454 VDD.n2745 VDD.n2744 15.6358
R15455 VDD.n2744 VDD.n2743 15.6358
R15456 VDD.n2743 VDD.n80 15.6358
R15457 VDD.n2737 VDD.n80 15.6358
R15458 VDD.n2736 VDD.n2735 15.6358
R15459 VDD.n2735 VDD.n91 15.6358
R15460 VDD.n2729 VDD.n91 15.6358
R15461 VDD.n2729 VDD.n2728 15.6358
R15462 VDD.n2728 VDD.n2727 15.6358
R15463 VDD.n1349 VDD.t4 15.3231
R15464 VDD.n1424 VDD.t7 15.3231
R15465 VDD.n2550 VDD.t137 15.3231
R15466 VDD.n2761 VDD.t0 15.3231
R15467 VDD.n1301 VDD.t68 12.5087
R15468 VDD.n1472 VDD.t61 12.5087
R15469 VDD.n2502 VDD.t83 12.5087
R15470 VDD.n2737 VDD.t57 12.5087
R15471 VDD.n1689 VDD.n1606 10.9146
R15472 VDD.n2307 VDD.n314 10.9146
R15473 VDD.n2385 VDD.n2346 10.9146
R15474 VDD.n1541 VDD.n884 10.9146
R15475 VDD.n1711 VDD.n698 10.6325
R15476 VDD.n1711 VDD.n692 10.6325
R15477 VDD.n1717 VDD.n692 10.6325
R15478 VDD.n1717 VDD.n685 10.6325
R15479 VDD.n1723 VDD.n685 10.6325
R15480 VDD.n1723 VDD.n688 10.6325
R15481 VDD.n1735 VDD.n674 10.6325
R15482 VDD.n1735 VDD.n668 10.6325
R15483 VDD.n1741 VDD.n668 10.6325
R15484 VDD.n1741 VDD.n662 10.6325
R15485 VDD.n1747 VDD.n662 10.6325
R15486 VDD.n1747 VDD.n656 10.6325
R15487 VDD.n1753 VDD.n656 10.6325
R15488 VDD.n1753 VDD.n650 10.6325
R15489 VDD.n1759 VDD.n650 10.6325
R15490 VDD.n1759 VDD.t17 10.6325
R15491 VDD.n1765 VDD.t17 10.6325
R15492 VDD.n1765 VDD.n639 10.6325
R15493 VDD.n1771 VDD.n639 10.6325
R15494 VDD.n1771 VDD.n633 10.6325
R15495 VDD.t16 VDD.n633 10.6325
R15496 VDD.t16 VDD.n627 10.6325
R15497 VDD.n1782 VDD.n627 10.6325
R15498 VDD.n1782 VDD.n621 10.6325
R15499 VDD.n1788 VDD.n621 10.6325
R15500 VDD.n1788 VDD.n615 10.6325
R15501 VDD.n1794 VDD.n615 10.6325
R15502 VDD.n1800 VDD.n609 10.6325
R15503 VDD.n1800 VDD.n603 10.6325
R15504 VDD.n1806 VDD.n603 10.6325
R15505 VDD.n1806 VDD.n597 10.6325
R15506 VDD.n1812 VDD.n597 10.6325
R15507 VDD.n1812 VDD.n590 10.6325
R15508 VDD.n1818 VDD.n590 10.6325
R15509 VDD.n1818 VDD.n593 10.6325
R15510 VDD.n1824 VDD.n586 10.6325
R15511 VDD.n1835 VDD.n572 10.6325
R15512 VDD.n1841 VDD.n572 10.6325
R15513 VDD.n1841 VDD.n561 10.6325
R15514 VDD.n1883 VDD.n561 10.6325
R15515 VDD.n1883 VDD.n537 10.6325
R15516 VDD.n2136 VDD.n531 10.6325
R15517 VDD.n2136 VDD.n525 10.6325
R15518 VDD.n2142 VDD.n525 10.6325
R15519 VDD.n2142 VDD.n519 10.6325
R15520 VDD.n2148 VDD.n519 10.6325
R15521 VDD.n2154 VDD.n513 10.6325
R15522 VDD.n2160 VDD.n507 10.6325
R15523 VDD.n2160 VDD.n501 10.6325
R15524 VDD.n2166 VDD.n501 10.6325
R15525 VDD.n2166 VDD.n495 10.6325
R15526 VDD.n2172 VDD.n495 10.6325
R15527 VDD.n2172 VDD.n488 10.6325
R15528 VDD.n2178 VDD.n488 10.6325
R15529 VDD.n2178 VDD.n491 10.6325
R15530 VDD.n2184 VDD.n477 10.6325
R15531 VDD.n2190 VDD.n477 10.6325
R15532 VDD.n2190 VDD.n471 10.6325
R15533 VDD.n2196 VDD.n471 10.6325
R15534 VDD.n2196 VDD.n465 10.6325
R15535 VDD.t23 VDD.n465 10.6325
R15536 VDD.t23 VDD.n459 10.6325
R15537 VDD.n2207 VDD.n459 10.6325
R15538 VDD.n2207 VDD.n453 10.6325
R15539 VDD.n2213 VDD.n453 10.6325
R15540 VDD.n2213 VDD.t19 10.6325
R15541 VDD.n2219 VDD.t19 10.6325
R15542 VDD.n2219 VDD.n442 10.6325
R15543 VDD.n2225 VDD.n442 10.6325
R15544 VDD.n2225 VDD.n436 10.6325
R15545 VDD.n2231 VDD.n436 10.6325
R15546 VDD.n2231 VDD.n430 10.6325
R15547 VDD.n2237 VDD.n430 10.6325
R15548 VDD.n2237 VDD.n423 10.6325
R15549 VDD.n2243 VDD.n423 10.6325
R15550 VDD.n2243 VDD.n426 10.6325
R15551 VDD.n2280 VDD.n411 10.6325
R15552 VDD.n2280 VDD.n405 10.6325
R15553 VDD.n2286 VDD.n405 10.6325
R15554 VDD.n2286 VDD.n382 10.6325
R15555 VDD.n2326 VDD.n382 10.6325
R15556 VDD.n2326 VDD.n384 10.6325
R15557 VDD.n1879 VDD.n1877 10.6151
R15558 VDD.n1877 VDD.n1874 10.6151
R15559 VDD.n1874 VDD.n1873 10.6151
R15560 VDD.n1873 VDD.n1870 10.6151
R15561 VDD.n1870 VDD.n1869 10.6151
R15562 VDD.n1869 VDD.n1866 10.6151
R15563 VDD.n1866 VDD.n1865 10.6151
R15564 VDD.n1865 VDD.n1862 10.6151
R15565 VDD.n1862 VDD.n1861 10.6151
R15566 VDD.n1861 VDD.n1858 10.6151
R15567 VDD.n1858 VDD.n1857 10.6151
R15568 VDD.n1854 VDD.n1853 10.6151
R15569 VDD.n1853 VDD.n1850 10.6151
R15570 VDD.n1850 VDD.n1849 10.6151
R15571 VDD.n1672 VDD.n1670 10.6151
R15572 VDD.n1670 VDD.n1669 10.6151
R15573 VDD.n1669 VDD.n1667 10.6151
R15574 VDD.n1667 VDD.n1666 10.6151
R15575 VDD.n1666 VDD.n1664 10.6151
R15576 VDD.n1664 VDD.n1663 10.6151
R15577 VDD.n1663 VDD.n1661 10.6151
R15578 VDD.n1661 VDD.n1660 10.6151
R15579 VDD.n1660 VDD.n1658 10.6151
R15580 VDD.n1658 VDD.n1657 10.6151
R15581 VDD.n1657 VDD.n1655 10.6151
R15582 VDD.n1655 VDD.n1654 10.6151
R15583 VDD.n1654 VDD.n1652 10.6151
R15584 VDD.n1652 VDD.n1651 10.6151
R15585 VDD.n1651 VDD.n1649 10.6151
R15586 VDD.n1649 VDD.n1648 10.6151
R15587 VDD.n1648 VDD.n1646 10.6151
R15588 VDD.n1646 VDD.n1645 10.6151
R15589 VDD.n1645 VDD.n1643 10.6151
R15590 VDD.n1643 VDD.n1642 10.6151
R15591 VDD.n1642 VDD.n1640 10.6151
R15592 VDD.n1640 VDD.n1639 10.6151
R15593 VDD.n1639 VDD.n1637 10.6151
R15594 VDD.n1637 VDD.n1636 10.6151
R15595 VDD.n1636 VDD.n1634 10.6151
R15596 VDD.n1634 VDD.n1633 10.6151
R15597 VDD.n1633 VDD.n1631 10.6151
R15598 VDD.n1631 VDD.n1630 10.6151
R15599 VDD.n1630 VDD.n1628 10.6151
R15600 VDD.n1628 VDD.n1627 10.6151
R15601 VDD.n1627 VDD.n1625 10.6151
R15602 VDD.n1625 VDD.n1624 10.6151
R15603 VDD.n1624 VDD.n1622 10.6151
R15604 VDD.n1622 VDD.n1621 10.6151
R15605 VDD.n1621 VDD.n1619 10.6151
R15606 VDD.n1619 VDD.n1618 10.6151
R15607 VDD.n1618 VDD.n1616 10.6151
R15608 VDD.n1616 VDD.n1615 10.6151
R15609 VDD.n1615 VDD.n1613 10.6151
R15610 VDD.n1613 VDD.n1612 10.6151
R15611 VDD.n1612 VDD.n1610 10.6151
R15612 VDD.n1610 VDD.n1609 10.6151
R15613 VDD.n1609 VDD.n570 10.6151
R15614 VDD.n1844 VDD.n570 10.6151
R15615 VDD.n1845 VDD.n1844 10.6151
R15616 VDD.n1846 VDD.n1845 10.6151
R15617 VDD.n1702 VDD.n1701 10.6151
R15618 VDD.n1701 VDD.n1700 10.6151
R15619 VDD.n1700 VDD.n1699 10.6151
R15620 VDD.n1699 VDD.n1697 10.6151
R15621 VDD.n1697 VDD.n1694 10.6151
R15622 VDD.n1694 VDD.n1693 10.6151
R15623 VDD.n1693 VDD.n1690 10.6151
R15624 VDD.n1688 VDD.n1685 10.6151
R15625 VDD.n1685 VDD.n1684 10.6151
R15626 VDD.n1684 VDD.n1681 10.6151
R15627 VDD.n1679 VDD.n1676 10.6151
R15628 VDD.n1676 VDD.n1675 10.6151
R15629 VDD.n1675 VDD.n1673 10.6151
R15630 VDD.n1713 VDD.n696 10.6151
R15631 VDD.n1714 VDD.n1713 10.6151
R15632 VDD.n1715 VDD.n1714 10.6151
R15633 VDD.n1715 VDD.n683 10.6151
R15634 VDD.n1725 VDD.n683 10.6151
R15635 VDD.n1726 VDD.n1725 10.6151
R15636 VDD.n1727 VDD.n1726 10.6151
R15637 VDD.n1727 VDD.n672 10.6151
R15638 VDD.n1737 VDD.n672 10.6151
R15639 VDD.n1738 VDD.n1737 10.6151
R15640 VDD.n1739 VDD.n1738 10.6151
R15641 VDD.n1739 VDD.n660 10.6151
R15642 VDD.n1749 VDD.n660 10.6151
R15643 VDD.n1750 VDD.n1749 10.6151
R15644 VDD.n1751 VDD.n1750 10.6151
R15645 VDD.n1751 VDD.n648 10.6151
R15646 VDD.n1761 VDD.n648 10.6151
R15647 VDD.n1762 VDD.n1761 10.6151
R15648 VDD.n1763 VDD.n1762 10.6151
R15649 VDD.n1763 VDD.n637 10.6151
R15650 VDD.n1773 VDD.n637 10.6151
R15651 VDD.n1774 VDD.n1773 10.6151
R15652 VDD.n1775 VDD.n1774 10.6151
R15653 VDD.n1775 VDD.n625 10.6151
R15654 VDD.n1784 VDD.n625 10.6151
R15655 VDD.n1785 VDD.n1784 10.6151
R15656 VDD.n1786 VDD.n1785 10.6151
R15657 VDD.n1786 VDD.n613 10.6151
R15658 VDD.n1796 VDD.n613 10.6151
R15659 VDD.n1797 VDD.n1796 10.6151
R15660 VDD.n1798 VDD.n1797 10.6151
R15661 VDD.n1798 VDD.n601 10.6151
R15662 VDD.n1808 VDD.n601 10.6151
R15663 VDD.n1809 VDD.n1808 10.6151
R15664 VDD.n1810 VDD.n1809 10.6151
R15665 VDD.n1810 VDD.n588 10.6151
R15666 VDD.n1820 VDD.n588 10.6151
R15667 VDD.n1821 VDD.n1820 10.6151
R15668 VDD.n1822 VDD.n1821 10.6151
R15669 VDD.n1822 VDD.n576 10.6151
R15670 VDD.n1837 VDD.n576 10.6151
R15671 VDD.n1838 VDD.n1837 10.6151
R15672 VDD.n1839 VDD.n1838 10.6151
R15673 VDD.n1839 VDD.n566 10.6151
R15674 VDD.n1881 VDD.n566 10.6151
R15675 VDD.n1881 VDD.n1880 10.6151
R15676 VDD.n2097 VDD.n2095 10.6151
R15677 VDD.n2095 VDD.n2094 10.6151
R15678 VDD.n2094 VDD.n2092 10.6151
R15679 VDD.n2092 VDD.n2091 10.6151
R15680 VDD.n2091 VDD.n2089 10.6151
R15681 VDD.n2089 VDD.n2088 10.6151
R15682 VDD.n2088 VDD.n2086 10.6151
R15683 VDD.n2086 VDD.n2085 10.6151
R15684 VDD.n2085 VDD.n2083 10.6151
R15685 VDD.n2083 VDD.n2082 10.6151
R15686 VDD.n2082 VDD.n2080 10.6151
R15687 VDD.n2080 VDD.n2079 10.6151
R15688 VDD.n2079 VDD.n2077 10.6151
R15689 VDD.n2077 VDD.n2076 10.6151
R15690 VDD.n2076 VDD.n2074 10.6151
R15691 VDD.n2074 VDD.n2073 10.6151
R15692 VDD.n2073 VDD.n2071 10.6151
R15693 VDD.n2071 VDD.n2070 10.6151
R15694 VDD.n2070 VDD.n2068 10.6151
R15695 VDD.n2068 VDD.n2067 10.6151
R15696 VDD.n2067 VDD.n2065 10.6151
R15697 VDD.n2065 VDD.n2064 10.6151
R15698 VDD.n2064 VDD.n2062 10.6151
R15699 VDD.n2062 VDD.n2061 10.6151
R15700 VDD.n2061 VDD.n2059 10.6151
R15701 VDD.n2059 VDD.n2058 10.6151
R15702 VDD.n2058 VDD.n2056 10.6151
R15703 VDD.n2056 VDD.n2055 10.6151
R15704 VDD.n2055 VDD.n2053 10.6151
R15705 VDD.n2053 VDD.n2052 10.6151
R15706 VDD.n2052 VDD.n2050 10.6151
R15707 VDD.n2050 VDD.n2049 10.6151
R15708 VDD.n2049 VDD.n2047 10.6151
R15709 VDD.n2047 VDD.n2046 10.6151
R15710 VDD.n2046 VDD.n2044 10.6151
R15711 VDD.n2044 VDD.n2043 10.6151
R15712 VDD.n2043 VDD.n2041 10.6151
R15713 VDD.n2041 VDD.n2040 10.6151
R15714 VDD.n2040 VDD.n2038 10.6151
R15715 VDD.n2038 VDD.n2037 10.6151
R15716 VDD.n2037 VDD.n2035 10.6151
R15717 VDD.n2035 VDD.n2034 10.6151
R15718 VDD.n2034 VDD.n403 10.6151
R15719 VDD.n2289 VDD.n403 10.6151
R15720 VDD.n2290 VDD.n2289 10.6151
R15721 VDD.n2291 VDD.n2290 10.6151
R15722 VDD.n2126 VDD.n2125 10.6151
R15723 VDD.n2125 VDD.n2124 10.6151
R15724 VDD.n2124 VDD.n2123 10.6151
R15725 VDD.n2123 VDD.n2121 10.6151
R15726 VDD.n2121 VDD.n2118 10.6151
R15727 VDD.n2118 VDD.n2117 10.6151
R15728 VDD.n2117 VDD.n2114 10.6151
R15729 VDD.n2114 VDD.n2113 10.6151
R15730 VDD.n2113 VDD.n2110 10.6151
R15731 VDD.n2110 VDD.n2109 10.6151
R15732 VDD.n2109 VDD.n2106 10.6151
R15733 VDD.n2104 VDD.n2101 10.6151
R15734 VDD.n2101 VDD.n2100 10.6151
R15735 VDD.n2100 VDD.n2098 10.6151
R15736 VDD.n2138 VDD.n529 10.6151
R15737 VDD.n2139 VDD.n2138 10.6151
R15738 VDD.n2140 VDD.n2139 10.6151
R15739 VDD.n2140 VDD.n517 10.6151
R15740 VDD.n2150 VDD.n517 10.6151
R15741 VDD.n2151 VDD.n2150 10.6151
R15742 VDD.n2152 VDD.n2151 10.6151
R15743 VDD.n2152 VDD.n505 10.6151
R15744 VDD.n2162 VDD.n505 10.6151
R15745 VDD.n2163 VDD.n2162 10.6151
R15746 VDD.n2164 VDD.n2163 10.6151
R15747 VDD.n2164 VDD.n493 10.6151
R15748 VDD.n2174 VDD.n493 10.6151
R15749 VDD.n2175 VDD.n2174 10.6151
R15750 VDD.n2176 VDD.n2175 10.6151
R15751 VDD.n2176 VDD.n481 10.6151
R15752 VDD.n2186 VDD.n481 10.6151
R15753 VDD.n2187 VDD.n2186 10.6151
R15754 VDD.n2188 VDD.n2187 10.6151
R15755 VDD.n2188 VDD.n469 10.6151
R15756 VDD.n2198 VDD.n469 10.6151
R15757 VDD.n2199 VDD.n2198 10.6151
R15758 VDD.n2200 VDD.n2199 10.6151
R15759 VDD.n2200 VDD.n457 10.6151
R15760 VDD.n2209 VDD.n457 10.6151
R15761 VDD.n2210 VDD.n2209 10.6151
R15762 VDD.n2211 VDD.n2210 10.6151
R15763 VDD.n2211 VDD.n446 10.6151
R15764 VDD.n2221 VDD.n446 10.6151
R15765 VDD.n2222 VDD.n2221 10.6151
R15766 VDD.n2223 VDD.n2222 10.6151
R15767 VDD.n2223 VDD.n434 10.6151
R15768 VDD.n2233 VDD.n434 10.6151
R15769 VDD.n2234 VDD.n2233 10.6151
R15770 VDD.n2235 VDD.n2234 10.6151
R15771 VDD.n2235 VDD.n421 10.6151
R15772 VDD.n2245 VDD.n421 10.6151
R15773 VDD.n2246 VDD.n2245 10.6151
R15774 VDD.n2247 VDD.n2246 10.6151
R15775 VDD.n2247 VDD.n409 10.6151
R15776 VDD.n2282 VDD.n409 10.6151
R15777 VDD.n2283 VDD.n2282 10.6151
R15778 VDD.n2284 VDD.n2283 10.6151
R15779 VDD.n2284 VDD.n388 10.6151
R15780 VDD.n2324 VDD.n388 10.6151
R15781 VDD.n2324 VDD.n2323 10.6151
R15782 VDD.n2322 VDD.n389 10.6151
R15783 VDD.n390 VDD.n389 10.6151
R15784 VDD.n2315 VDD.n390 10.6151
R15785 VDD.n2315 VDD.n2314 10.6151
R15786 VDD.n2314 VDD.n2313 10.6151
R15787 VDD.n2313 VDD.n392 10.6151
R15788 VDD.n2308 VDD.n392 10.6151
R15789 VDD.n2306 VDD.n2305 10.6151
R15790 VDD.n2305 VDD.n395 10.6151
R15791 VDD.n2300 VDD.n395 10.6151
R15792 VDD.n2298 VDD.n2297 10.6151
R15793 VDD.n2297 VDD.n400 10.6151
R15794 VDD.n2292 VDD.n400 10.6151
R15795 VDD.n2267 VDD.n2253 10.6151
R15796 VDD.n2267 VDD.n2266 10.6151
R15797 VDD.n2266 VDD.n2265 10.6151
R15798 VDD.n2265 VDD.n2255 10.6151
R15799 VDD.n2260 VDD.n2255 10.6151
R15800 VDD.n2260 VDD.n2259 10.6151
R15801 VDD.n2259 VDD.n369 10.6151
R15802 VDD.n2345 VDD.n370 10.6151
R15803 VDD.n373 VDD.n370 10.6151
R15804 VDD.n2338 VDD.n373 10.6151
R15805 VDD.n2336 VDD.n2335 10.6151
R15806 VDD.n2335 VDD.n377 10.6151
R15807 VDD.n2330 VDD.n377 10.6151
R15808 VDD.n2000 VDD.n1999 10.6151
R15809 VDD.n1999 VDD.n1998 10.6151
R15810 VDD.n1998 VDD.n1996 10.6151
R15811 VDD.n1996 VDD.n1995 10.6151
R15812 VDD.n1995 VDD.n1993 10.6151
R15813 VDD.n1993 VDD.n1992 10.6151
R15814 VDD.n1992 VDD.n1990 10.6151
R15815 VDD.n1990 VDD.n1989 10.6151
R15816 VDD.n1989 VDD.n1987 10.6151
R15817 VDD.n1987 VDD.n1986 10.6151
R15818 VDD.n1986 VDD.n1984 10.6151
R15819 VDD.n1984 VDD.n1983 10.6151
R15820 VDD.n1983 VDD.n1981 10.6151
R15821 VDD.n1981 VDD.n1980 10.6151
R15822 VDD.n1980 VDD.n1978 10.6151
R15823 VDD.n1978 VDD.n1977 10.6151
R15824 VDD.n1977 VDD.n1975 10.6151
R15825 VDD.n1975 VDD.n1974 10.6151
R15826 VDD.n1974 VDD.n1972 10.6151
R15827 VDD.n1972 VDD.n1971 10.6151
R15828 VDD.n1971 VDD.n1969 10.6151
R15829 VDD.n1969 VDD.n1968 10.6151
R15830 VDD.n1968 VDD.n1966 10.6151
R15831 VDD.n1966 VDD.n1965 10.6151
R15832 VDD.n1965 VDD.n1963 10.6151
R15833 VDD.n1963 VDD.n1962 10.6151
R15834 VDD.n1962 VDD.n1960 10.6151
R15835 VDD.n1960 VDD.n1959 10.6151
R15836 VDD.n1959 VDD.n1957 10.6151
R15837 VDD.n1957 VDD.n1956 10.6151
R15838 VDD.n1956 VDD.n1954 10.6151
R15839 VDD.n1954 VDD.n1953 10.6151
R15840 VDD.n1953 VDD.n1951 10.6151
R15841 VDD.n1951 VDD.n1950 10.6151
R15842 VDD.n1950 VDD.n1948 10.6151
R15843 VDD.n1948 VDD.n1947 10.6151
R15844 VDD.n1947 VDD.n1945 10.6151
R15845 VDD.n1945 VDD.n1944 10.6151
R15846 VDD.n1944 VDD.n1942 10.6151
R15847 VDD.n1942 VDD.n1941 10.6151
R15848 VDD.n1941 VDD.n1939 10.6151
R15849 VDD.n1939 VDD.n1938 10.6151
R15850 VDD.n1938 VDD.n1936 10.6151
R15851 VDD.n1936 VDD.n380 10.6151
R15852 VDD.n2328 VDD.n380 10.6151
R15853 VDD.n2329 VDD.n2328 10.6151
R15854 VDD.n2132 VDD.n535 10.6151
R15855 VDD.n2027 VDD.n535 10.6151
R15856 VDD.n2027 VDD.n2026 10.6151
R15857 VDD.n2026 VDD.n2025 10.6151
R15858 VDD.n2025 VDD.n2023 10.6151
R15859 VDD.n2023 VDD.n2020 10.6151
R15860 VDD.n2020 VDD.n2019 10.6151
R15861 VDD.n2019 VDD.n2016 10.6151
R15862 VDD.n2016 VDD.n2015 10.6151
R15863 VDD.n2015 VDD.n2012 10.6151
R15864 VDD.n2012 VDD.n2011 10.6151
R15865 VDD.n2008 VDD.n2007 10.6151
R15866 VDD.n2007 VDD.n2004 10.6151
R15867 VDD.n2004 VDD.n2003 10.6151
R15868 VDD.n2134 VDD.n2133 10.6151
R15869 VDD.n2134 VDD.n523 10.6151
R15870 VDD.n2144 VDD.n523 10.6151
R15871 VDD.n2145 VDD.n2144 10.6151
R15872 VDD.n2146 VDD.n2145 10.6151
R15873 VDD.n2146 VDD.n511 10.6151
R15874 VDD.n2156 VDD.n511 10.6151
R15875 VDD.n2157 VDD.n2156 10.6151
R15876 VDD.n2158 VDD.n2157 10.6151
R15877 VDD.n2158 VDD.n499 10.6151
R15878 VDD.n2168 VDD.n499 10.6151
R15879 VDD.n2169 VDD.n2168 10.6151
R15880 VDD.n2170 VDD.n2169 10.6151
R15881 VDD.n2170 VDD.n486 10.6151
R15882 VDD.n2180 VDD.n486 10.6151
R15883 VDD.n2181 VDD.n2180 10.6151
R15884 VDD.n2182 VDD.n2181 10.6151
R15885 VDD.n2182 VDD.n475 10.6151
R15886 VDD.n2192 VDD.n475 10.6151
R15887 VDD.n2193 VDD.n2192 10.6151
R15888 VDD.n2194 VDD.n2193 10.6151
R15889 VDD.n2194 VDD.n463 10.6151
R15890 VDD.n2203 VDD.n463 10.6151
R15891 VDD.n2204 VDD.n2203 10.6151
R15892 VDD.n2205 VDD.n2204 10.6151
R15893 VDD.n2205 VDD.n451 10.6151
R15894 VDD.n2215 VDD.n451 10.6151
R15895 VDD.n2216 VDD.n2215 10.6151
R15896 VDD.n2217 VDD.n2216 10.6151
R15897 VDD.n2217 VDD.n440 10.6151
R15898 VDD.n2227 VDD.n440 10.6151
R15899 VDD.n2228 VDD.n2227 10.6151
R15900 VDD.n2229 VDD.n2228 10.6151
R15901 VDD.n2229 VDD.n428 10.6151
R15902 VDD.n2239 VDD.n428 10.6151
R15903 VDD.n2240 VDD.n2239 10.6151
R15904 VDD.n2241 VDD.n2240 10.6151
R15905 VDD.n2241 VDD.n416 10.6151
R15906 VDD.n2251 VDD.n416 10.6151
R15907 VDD.n2252 VDD.n2251 10.6151
R15908 VDD.n2278 VDD.n2252 10.6151
R15909 VDD.n2278 VDD.n2277 10.6151
R15910 VDD.n2277 VDD.n2276 10.6151
R15911 VDD.n2276 VDD.n2275 10.6151
R15912 VDD.n2275 VDD.n2273 10.6151
R15913 VDD.n2273 VDD.n2272 10.6151
R15914 VDD.n1709 VDD.n1708 10.6151
R15915 VDD.n1709 VDD.n690 10.6151
R15916 VDD.n1719 VDD.n690 10.6151
R15917 VDD.n1720 VDD.n1719 10.6151
R15918 VDD.n1721 VDD.n1720 10.6151
R15919 VDD.n1721 VDD.n678 10.6151
R15920 VDD.n1731 VDD.n678 10.6151
R15921 VDD.n1732 VDD.n1731 10.6151
R15922 VDD.n1733 VDD.n1732 10.6151
R15923 VDD.n1733 VDD.n666 10.6151
R15924 VDD.n1743 VDD.n666 10.6151
R15925 VDD.n1744 VDD.n1743 10.6151
R15926 VDD.n1745 VDD.n1744 10.6151
R15927 VDD.n1745 VDD.n654 10.6151
R15928 VDD.n1755 VDD.n654 10.6151
R15929 VDD.n1756 VDD.n1755 10.6151
R15930 VDD.n1757 VDD.n1756 10.6151
R15931 VDD.n1757 VDD.n643 10.6151
R15932 VDD.n1767 VDD.n643 10.6151
R15933 VDD.n1768 VDD.n1767 10.6151
R15934 VDD.n1769 VDD.n1768 10.6151
R15935 VDD.n1769 VDD.n631 10.6151
R15936 VDD.n1778 VDD.n631 10.6151
R15937 VDD.n1779 VDD.n1778 10.6151
R15938 VDD.n1780 VDD.n1779 10.6151
R15939 VDD.n1780 VDD.n619 10.6151
R15940 VDD.n1790 VDD.n619 10.6151
R15941 VDD.n1791 VDD.n1790 10.6151
R15942 VDD.n1792 VDD.n1791 10.6151
R15943 VDD.n1792 VDD.n607 10.6151
R15944 VDD.n1802 VDD.n607 10.6151
R15945 VDD.n1803 VDD.n1802 10.6151
R15946 VDD.n1804 VDD.n1803 10.6151
R15947 VDD.n1804 VDD.n595 10.6151
R15948 VDD.n1814 VDD.n595 10.6151
R15949 VDD.n1815 VDD.n1814 10.6151
R15950 VDD.n1816 VDD.n1815 10.6151
R15951 VDD.n1816 VDD.n582 10.6151
R15952 VDD.n1826 VDD.n582 10.6151
R15953 VDD.n1827 VDD.n1826 10.6151
R15954 VDD.n1833 VDD.n1827 10.6151
R15955 VDD.n1833 VDD.n1832 10.6151
R15956 VDD.n1832 VDD.n1831 10.6151
R15957 VDD.n1831 VDD.n1830 10.6151
R15958 VDD.n1830 VDD.n1828 10.6151
R15959 VDD.n1828 VDD.n556 10.6151
R15960 VDD.n1916 VDD.n1915 10.6151
R15961 VDD.n1915 VDD.n1914 10.6151
R15962 VDD.n1914 VDD.n1911 10.6151
R15963 VDD.n1911 VDD.n1910 10.6151
R15964 VDD.n1910 VDD.n1907 10.6151
R15965 VDD.n1907 VDD.n1906 10.6151
R15966 VDD.n1906 VDD.n1903 10.6151
R15967 VDD.n1903 VDD.n1902 10.6151
R15968 VDD.n1902 VDD.n1899 10.6151
R15969 VDD.n1899 VDD.n1898 10.6151
R15970 VDD.n1898 VDD.n1895 10.6151
R15971 VDD.n1893 VDD.n1890 10.6151
R15972 VDD.n1890 VDD.n1889 10.6151
R15973 VDD.n1889 VDD.n1887 10.6151
R15974 VDD.n867 VDD.n865 10.6151
R15975 VDD.n865 VDD.n864 10.6151
R15976 VDD.n864 VDD.n862 10.6151
R15977 VDD.n862 VDD.n861 10.6151
R15978 VDD.n861 VDD.n859 10.6151
R15979 VDD.n859 VDD.n858 10.6151
R15980 VDD.n858 VDD.n856 10.6151
R15981 VDD.n856 VDD.n855 10.6151
R15982 VDD.n855 VDD.n853 10.6151
R15983 VDD.n853 VDD.n852 10.6151
R15984 VDD.n852 VDD.n850 10.6151
R15985 VDD.n850 VDD.n849 10.6151
R15986 VDD.n849 VDD.n847 10.6151
R15987 VDD.n847 VDD.n846 10.6151
R15988 VDD.n846 VDD.n844 10.6151
R15989 VDD.n844 VDD.n843 10.6151
R15990 VDD.n843 VDD.n841 10.6151
R15991 VDD.n841 VDD.n840 10.6151
R15992 VDD.n840 VDD.n838 10.6151
R15993 VDD.n838 VDD.n837 10.6151
R15994 VDD.n837 VDD.n835 10.6151
R15995 VDD.n835 VDD.n834 10.6151
R15996 VDD.n834 VDD.n832 10.6151
R15997 VDD.n832 VDD.n831 10.6151
R15998 VDD.n831 VDD.n829 10.6151
R15999 VDD.n829 VDD.n828 10.6151
R16000 VDD.n828 VDD.n826 10.6151
R16001 VDD.n826 VDD.n825 10.6151
R16002 VDD.n825 VDD.n823 10.6151
R16003 VDD.n823 VDD.n822 10.6151
R16004 VDD.n822 VDD.n820 10.6151
R16005 VDD.n820 VDD.n819 10.6151
R16006 VDD.n819 VDD.n817 10.6151
R16007 VDD.n817 VDD.n816 10.6151
R16008 VDD.n816 VDD.n814 10.6151
R16009 VDD.n814 VDD.n813 10.6151
R16010 VDD.n813 VDD.n811 10.6151
R16011 VDD.n811 VDD.n810 10.6151
R16012 VDD.n810 VDD.n808 10.6151
R16013 VDD.n808 VDD.n807 10.6151
R16014 VDD.n807 VDD.n805 10.6151
R16015 VDD.n805 VDD.n804 10.6151
R16016 VDD.n804 VDD.n802 10.6151
R16017 VDD.n802 VDD.n801 10.6151
R16018 VDD.n801 VDD.n559 10.6151
R16019 VDD.n1886 VDD.n559 10.6151
R16020 VDD.n1707 VDD.n702 10.6151
R16021 VDD.n787 VDD.n702 10.6151
R16022 VDD.n790 VDD.n787 10.6151
R16023 VDD.n791 VDD.n790 10.6151
R16024 VDD.n794 VDD.n791 10.6151
R16025 VDD.n795 VDD.n794 10.6151
R16026 VDD.n798 VDD.n795 10.6151
R16027 VDD.n883 VDD.n880 10.6151
R16028 VDD.n880 VDD.n879 10.6151
R16029 VDD.n879 VDD.n876 10.6151
R16030 VDD.n874 VDD.n871 10.6151
R16031 VDD.n871 VDD.n870 10.6151
R16032 VDD.n870 VDD.n868 10.6151
R16033 VDD.n1857 VDD.n569 9.99074
R16034 VDD.n1681 VDD.n1680 9.99074
R16035 VDD.n2106 VDD.n2105 9.99074
R16036 VDD.n2300 VDD.n2299 9.99074
R16037 VDD.n2338 VDD.n2337 9.99074
R16038 VDD.n2011 VDD.n1935 9.99074
R16039 VDD.n1895 VDD.n1894 9.99074
R16040 VDD.n876 VDD.n875 9.99074
R16041 VDD.n1396 VDD.n991 9.3005
R16042 VDD.n1398 VDD.n1397 9.3005
R16043 VDD.n981 VDD.n980 9.3005
R16044 VDD.n1411 VDD.n1410 9.3005
R16045 VDD.n1412 VDD.n979 9.3005
R16046 VDD.n1414 VDD.n1413 9.3005
R16047 VDD.n969 VDD.n968 9.3005
R16048 VDD.n1427 VDD.n1426 9.3005
R16049 VDD.n1428 VDD.n967 9.3005
R16050 VDD.n1430 VDD.n1429 9.3005
R16051 VDD.n957 VDD.n956 9.3005
R16052 VDD.n1443 VDD.n1442 9.3005
R16053 VDD.n1444 VDD.n955 9.3005
R16054 VDD.n1446 VDD.n1445 9.3005
R16055 VDD.n945 VDD.n944 9.3005
R16056 VDD.n1459 VDD.n1458 9.3005
R16057 VDD.n1460 VDD.n943 9.3005
R16058 VDD.n1462 VDD.n1461 9.3005
R16059 VDD.n933 VDD.n932 9.3005
R16060 VDD.n1475 VDD.n1474 9.3005
R16061 VDD.n1476 VDD.n931 9.3005
R16062 VDD.n1478 VDD.n1477 9.3005
R16063 VDD.n920 VDD.n919 9.3005
R16064 VDD.n1492 VDD.n1491 9.3005
R16065 VDD.n1493 VDD.n918 9.3005
R16066 VDD.n1522 VDD.n1521 9.3005
R16067 VDD.n1545 VDD.n782 9.3005
R16068 VDD.n1544 VDD.n783 9.3005
R16069 VDD.n1571 VDD.n753 9.3005
R16070 VDD.n757 VDD.n754 9.3005
R16071 VDD.n1566 VDD.n758 9.3005
R16072 VDD.n1565 VDD.n759 9.3005
R16073 VDD.n1564 VDD.n760 9.3005
R16074 VDD.n764 VDD.n761 9.3005
R16075 VDD.n1559 VDD.n765 9.3005
R16076 VDD.n1558 VDD.n766 9.3005
R16077 VDD.n1557 VDD.n767 9.3005
R16078 VDD.n771 VDD.n768 9.3005
R16079 VDD.n1552 VDD.n772 9.3005
R16080 VDD.n1551 VDD.n773 9.3005
R16081 VDD.n1550 VDD.n774 9.3005
R16082 VDD.n781 VDD.n775 9.3005
R16083 VDD.n1596 VDD.n722 9.3005
R16084 VDD.n1595 VDD.n732 9.3005
R16085 VDD.n736 VDD.n733 9.3005
R16086 VDD.n1590 VDD.n737 9.3005
R16087 VDD.n1589 VDD.n738 9.3005
R16088 VDD.n1588 VDD.n739 9.3005
R16089 VDD.n743 VDD.n740 9.3005
R16090 VDD.n1583 VDD.n744 9.3005
R16091 VDD.n1582 VDD.n745 9.3005
R16092 VDD.n1581 VDD.n746 9.3005
R16093 VDD.n750 VDD.n747 9.3005
R16094 VDD.n1576 VDD.n751 9.3005
R16095 VDD.n1575 VDD.n752 9.3005
R16096 VDD.n1518 VDD.n1494 9.3005
R16097 VDD.n1498 VDD.n1495 9.3005
R16098 VDD.n1499 VDD.n1496 9.3005
R16099 VDD.n1511 VDD.n1500 9.3005
R16100 VDD.n1510 VDD.n1501 9.3005
R16101 VDD.n1509 VDD.n1502 9.3005
R16102 VDD.n1504 VDD.n1503 9.3005
R16103 VDD.n725 VDD.n721 9.3005
R16104 VDD.n1520 VDD.n1519 9.3005
R16105 VDD.n2397 VDD.n362 9.3005
R16106 VDD.n2398 VDD.n361 9.3005
R16107 VDD.n360 VDD.n358 9.3005
R16108 VDD.n2404 VDD.n357 9.3005
R16109 VDD.n2405 VDD.n356 9.3005
R16110 VDD.n2406 VDD.n355 9.3005
R16111 VDD.n354 VDD.n352 9.3005
R16112 VDD.n2412 VDD.n351 9.3005
R16113 VDD.n2413 VDD.n350 9.3005
R16114 VDD.n2414 VDD.n349 9.3005
R16115 VDD.n348 VDD.n346 9.3005
R16116 VDD.n2420 VDD.n345 9.3005
R16117 VDD.n2421 VDD.n344 9.3005
R16118 VDD.n2422 VDD.n343 9.3005
R16119 VDD.n2428 VDD.n336 9.3005
R16120 VDD.n2429 VDD.n335 9.3005
R16121 VDD.n2430 VDD.n334 9.3005
R16122 VDD.n333 VDD.n331 9.3005
R16123 VDD.n2436 VDD.n330 9.3005
R16124 VDD.n2437 VDD.n329 9.3005
R16125 VDD.n2438 VDD.n328 9.3005
R16126 VDD.n327 VDD.n325 9.3005
R16127 VDD.n2443 VDD.n324 9.3005
R16128 VDD.n2444 VDD.n323 9.3005
R16129 VDD.n322 VDD.n320 9.3005
R16130 VDD.n2449 VDD.n319 9.3005
R16131 VDD.n342 VDD.n337 9.3005
R16132 VDD.n2450 VDD.n314 9.3005
R16133 VDD.n314 VDD.n312 9.3005
R16134 VDD.n2459 VDD.n311 9.3005
R16135 VDD.n2460 VDD.n310 9.3005
R16136 VDD.n2461 VDD.n309 9.3005
R16137 VDD.n308 VDD.n306 9.3005
R16138 VDD.n2466 VDD.n305 9.3005
R16139 VDD.n2467 VDD.n304 9.3005
R16140 VDD.n303 VDD.n301 9.3005
R16141 VDD.n2472 VDD.n300 9.3005
R16142 VDD.n2474 VDD.n2473 9.3005
R16143 VDD.n2476 VDD.n2475 9.3005
R16144 VDD.n291 VDD.n290 9.3005
R16145 VDD.n2489 VDD.n2488 9.3005
R16146 VDD.n2490 VDD.n289 9.3005
R16147 VDD.n2492 VDD.n2491 9.3005
R16148 VDD.n279 VDD.n278 9.3005
R16149 VDD.n2505 VDD.n2504 9.3005
R16150 VDD.n2506 VDD.n277 9.3005
R16151 VDD.n2508 VDD.n2507 9.3005
R16152 VDD.n267 VDD.n266 9.3005
R16153 VDD.n2521 VDD.n2520 9.3005
R16154 VDD.n2522 VDD.n265 9.3005
R16155 VDD.n2524 VDD.n2523 9.3005
R16156 VDD.n255 VDD.n254 9.3005
R16157 VDD.n2537 VDD.n2536 9.3005
R16158 VDD.n2538 VDD.n253 9.3005
R16159 VDD.n2540 VDD.n2539 9.3005
R16160 VDD.n243 VDD.n242 9.3005
R16161 VDD.n2553 VDD.n2552 9.3005
R16162 VDD.n2554 VDD.n241 9.3005
R16163 VDD.n2556 VDD.n2555 9.3005
R16164 VDD.n231 VDD.n230 9.3005
R16165 VDD.n2569 VDD.n2568 9.3005
R16166 VDD.n2570 VDD.n229 9.3005
R16167 VDD.n2572 VDD.n2571 9.3005
R16168 VDD.n29 VDD.n27 9.3005
R16169 VDD.n2779 VDD.n2778 9.3005
R16170 VDD.n30 VDD.n28 9.3005
R16171 VDD.n2773 VDD.n39 9.3005
R16172 VDD.n2772 VDD.n40 9.3005
R16173 VDD.n2771 VDD.n41 9.3005
R16174 VDD.n49 VDD.n42 9.3005
R16175 VDD.n2765 VDD.n50 9.3005
R16176 VDD.n2764 VDD.n51 9.3005
R16177 VDD.n2763 VDD.n52 9.3005
R16178 VDD.n60 VDD.n53 9.3005
R16179 VDD.n2757 VDD.n61 9.3005
R16180 VDD.n2756 VDD.n62 9.3005
R16181 VDD.n2755 VDD.n63 9.3005
R16182 VDD.n71 VDD.n64 9.3005
R16183 VDD.n2749 VDD.n72 9.3005
R16184 VDD.n2748 VDD.n73 9.3005
R16185 VDD.n2747 VDD.n74 9.3005
R16186 VDD.n82 VDD.n75 9.3005
R16187 VDD.n2741 VDD.n83 9.3005
R16188 VDD.n2740 VDD.n84 9.3005
R16189 VDD.n2739 VDD.n85 9.3005
R16190 VDD.n93 VDD.n86 9.3005
R16191 VDD.n2733 VDD.n94 9.3005
R16192 VDD.n2732 VDD.n95 9.3005
R16193 VDD.n2731 VDD.n96 9.3005
R16194 VDD.n104 VDD.n97 9.3005
R16195 VDD.n2725 VDD.n2724 9.3005
R16196 VDD.n2721 VDD.n105 9.3005
R16197 VDD.n2720 VDD.n107 9.3005
R16198 VDD.n111 VDD.n108 9.3005
R16199 VDD.n2715 VDD.n112 9.3005
R16200 VDD.n2714 VDD.n113 9.3005
R16201 VDD.n2713 VDD.n114 9.3005
R16202 VDD.n118 VDD.n115 9.3005
R16203 VDD.n2708 VDD.n119 9.3005
R16204 VDD.n2707 VDD.n120 9.3005
R16205 VDD.n2706 VDD.n121 9.3005
R16206 VDD.n127 VDD.n124 9.3005
R16207 VDD.n2701 VDD.n128 9.3005
R16208 VDD.n2700 VDD.n129 9.3005
R16209 VDD.n2699 VDD.n130 9.3005
R16210 VDD.n134 VDD.n131 9.3005
R16211 VDD.n2694 VDD.n135 9.3005
R16212 VDD.n2693 VDD.n136 9.3005
R16213 VDD.n2692 VDD.n137 9.3005
R16214 VDD.n141 VDD.n138 9.3005
R16215 VDD.n2687 VDD.n142 9.3005
R16216 VDD.n2686 VDD.n143 9.3005
R16217 VDD.n2685 VDD.n144 9.3005
R16218 VDD.n148 VDD.n145 9.3005
R16219 VDD.n2680 VDD.n149 9.3005
R16220 VDD.n2679 VDD.n150 9.3005
R16221 VDD.n2675 VDD.n151 9.3005
R16222 VDD.n155 VDD.n152 9.3005
R16223 VDD.n2670 VDD.n156 9.3005
R16224 VDD.n2669 VDD.n157 9.3005
R16225 VDD.n2668 VDD.n158 9.3005
R16226 VDD.n162 VDD.n159 9.3005
R16227 VDD.n2663 VDD.n163 9.3005
R16228 VDD.n2662 VDD.n164 9.3005
R16229 VDD.n2661 VDD.n165 9.3005
R16230 VDD.n169 VDD.n166 9.3005
R16231 VDD.n2656 VDD.n170 9.3005
R16232 VDD.n2655 VDD.n171 9.3005
R16233 VDD.n2654 VDD.n172 9.3005
R16234 VDD.n179 VDD.n173 9.3005
R16235 VDD.n2649 VDD.n180 9.3005
R16236 VDD.n2648 VDD.n181 9.3005
R16237 VDD.n2647 VDD.n182 9.3005
R16238 VDD.n186 VDD.n183 9.3005
R16239 VDD.n2642 VDD.n187 9.3005
R16240 VDD.n2641 VDD.n188 9.3005
R16241 VDD.n2640 VDD.n189 9.3005
R16242 VDD.n193 VDD.n190 9.3005
R16243 VDD.n2635 VDD.n194 9.3005
R16244 VDD.n2634 VDD.n195 9.3005
R16245 VDD.n2633 VDD.n196 9.3005
R16246 VDD.n200 VDD.n197 9.3005
R16247 VDD.n2628 VDD.n201 9.3005
R16248 VDD.n2627 VDD.n202 9.3005
R16249 VDD.n2623 VDD.n2620 9.3005
R16250 VDD.n2723 VDD.n2722 9.3005
R16251 VDD.n2482 VDD.n295 9.3005
R16252 VDD.n2484 VDD.n2483 9.3005
R16253 VDD.n284 VDD.n283 9.3005
R16254 VDD.n2497 VDD.n2496 9.3005
R16255 VDD.n2498 VDD.n282 9.3005
R16256 VDD.n2500 VDD.n2499 9.3005
R16257 VDD.n273 VDD.n272 9.3005
R16258 VDD.n2513 VDD.n2512 9.3005
R16259 VDD.n2514 VDD.n271 9.3005
R16260 VDD.n2516 VDD.n2515 9.3005
R16261 VDD.n261 VDD.n260 9.3005
R16262 VDD.n2529 VDD.n2528 9.3005
R16263 VDD.n2530 VDD.n259 9.3005
R16264 VDD.n2532 VDD.n2531 9.3005
R16265 VDD.n248 VDD.n247 9.3005
R16266 VDD.n2545 VDD.n2544 9.3005
R16267 VDD.n2546 VDD.n246 9.3005
R16268 VDD.n2548 VDD.n2547 9.3005
R16269 VDD.n237 VDD.n236 9.3005
R16270 VDD.n2561 VDD.n2560 9.3005
R16271 VDD.n2562 VDD.n235 9.3005
R16272 VDD.n2564 VDD.n2563 9.3005
R16273 VDD.n224 VDD.n223 9.3005
R16274 VDD.n2577 VDD.n2576 9.3005
R16275 VDD.n2578 VDD.n222 9.3005
R16276 VDD.n2580 VDD.n2579 9.3005
R16277 VDD.n2581 VDD.n221 9.3005
R16278 VDD.n2583 VDD.n2582 9.3005
R16279 VDD.n2584 VDD.n220 9.3005
R16280 VDD.n2586 VDD.n2585 9.3005
R16281 VDD.n2587 VDD.n218 9.3005
R16282 VDD.n2589 VDD.n2588 9.3005
R16283 VDD.n2590 VDD.n217 9.3005
R16284 VDD.n2592 VDD.n2591 9.3005
R16285 VDD.n2593 VDD.n215 9.3005
R16286 VDD.n2595 VDD.n2594 9.3005
R16287 VDD.n2596 VDD.n214 9.3005
R16288 VDD.n2598 VDD.n2597 9.3005
R16289 VDD.n2599 VDD.n212 9.3005
R16290 VDD.n2601 VDD.n2600 9.3005
R16291 VDD.n2602 VDD.n211 9.3005
R16292 VDD.n2604 VDD.n2603 9.3005
R16293 VDD.n2605 VDD.n209 9.3005
R16294 VDD.n2607 VDD.n2606 9.3005
R16295 VDD.n2608 VDD.n208 9.3005
R16296 VDD.n2610 VDD.n2609 9.3005
R16297 VDD.n2611 VDD.n206 9.3005
R16298 VDD.n2613 VDD.n2612 9.3005
R16299 VDD.n2614 VDD.n205 9.3005
R16300 VDD.n2616 VDD.n2615 9.3005
R16301 VDD.n2617 VDD.n203 9.3005
R16302 VDD.n2619 VDD.n2618 9.3005
R16303 VDD.n2481 VDD.n2480 9.3005
R16304 VDD.n2363 VDD.n296 9.3005
R16305 VDD.n2367 VDD.n2362 9.3005
R16306 VDD.n2368 VDD.n2361 9.3005
R16307 VDD.n2360 VDD.n2357 9.3005
R16308 VDD.n2374 VDD.n2356 9.3005
R16309 VDD.n2375 VDD.n2355 9.3005
R16310 VDD.n2376 VDD.n2354 9.3005
R16311 VDD.n2353 VDD.n2351 9.3005
R16312 VDD.n2382 VDD.n368 9.3005
R16313 VDD.n367 VDD.n364 9.3005
R16314 VDD.n2393 VDD.n363 9.3005
R16315 VDD.n1540 VDD.n1539 9.3005
R16316 VDD.n1538 VDD.n886 9.3005
R16317 VDD.n1537 VDD.n1536 9.3005
R16318 VDD.n1535 VDD.n898 9.3005
R16319 VDD.n1534 VDD.n1533 9.3005
R16320 VDD.n1532 VDD.n899 9.3005
R16321 VDD.n1531 VDD.n1530 9.3005
R16322 VDD.n1529 VDD.n906 9.3005
R16323 VDD.n1528 VDD.n1527 9.3005
R16324 VDD.n1281 VDD.n1069 9.3005
R16325 VDD.n1283 VDD.n1282 9.3005
R16326 VDD.n1058 VDD.n1057 9.3005
R16327 VDD.n1296 VDD.n1295 9.3005
R16328 VDD.n1297 VDD.n1056 9.3005
R16329 VDD.n1299 VDD.n1298 9.3005
R16330 VDD.n1047 VDD.n1046 9.3005
R16331 VDD.n1312 VDD.n1311 9.3005
R16332 VDD.n1313 VDD.n1045 9.3005
R16333 VDD.n1315 VDD.n1314 9.3005
R16334 VDD.n1035 VDD.n1034 9.3005
R16335 VDD.n1328 VDD.n1327 9.3005
R16336 VDD.n1329 VDD.n1033 9.3005
R16337 VDD.n1331 VDD.n1330 9.3005
R16338 VDD.n1022 VDD.n1021 9.3005
R16339 VDD.n1344 VDD.n1343 9.3005
R16340 VDD.n1345 VDD.n1020 9.3005
R16341 VDD.n1347 VDD.n1346 9.3005
R16342 VDD.n1011 VDD.n1010 9.3005
R16343 VDD.n1360 VDD.n1359 9.3005
R16344 VDD.n1361 VDD.n1009 9.3005
R16345 VDD.n1363 VDD.n1362 9.3005
R16346 VDD.n999 VDD.n998 9.3005
R16347 VDD.n1376 VDD.n1375 9.3005
R16348 VDD.n1377 VDD.n997 9.3005
R16349 VDD.n1379 VDD.n1378 9.3005
R16350 VDD.n987 VDD.n986 9.3005
R16351 VDD.n1403 VDD.n1402 9.3005
R16352 VDD.n1404 VDD.n985 9.3005
R16353 VDD.n1406 VDD.n1405 9.3005
R16354 VDD.n975 VDD.n974 9.3005
R16355 VDD.n1419 VDD.n1418 9.3005
R16356 VDD.n1420 VDD.n973 9.3005
R16357 VDD.n1422 VDD.n1421 9.3005
R16358 VDD.n963 VDD.n962 9.3005
R16359 VDD.n1435 VDD.n1434 9.3005
R16360 VDD.n1436 VDD.n961 9.3005
R16361 VDD.n1438 VDD.n1437 9.3005
R16362 VDD.n951 VDD.n950 9.3005
R16363 VDD.n1451 VDD.n1450 9.3005
R16364 VDD.n1452 VDD.n949 9.3005
R16365 VDD.n1454 VDD.n1453 9.3005
R16366 VDD.n939 VDD.n938 9.3005
R16367 VDD.n1467 VDD.n1466 9.3005
R16368 VDD.n1468 VDD.n937 9.3005
R16369 VDD.n1470 VDD.n1469 9.3005
R16370 VDD.n927 VDD.n926 9.3005
R16371 VDD.n1483 VDD.n1482 9.3005
R16372 VDD.n1484 VDD.n924 9.3005
R16373 VDD.n1487 VDD.n1486 9.3005
R16374 VDD.n1485 VDD.n925 9.3005
R16375 VDD.n914 VDD.n907 9.3005
R16376 VDD.n1280 VDD.n1279 9.3005
R16377 VDD.n1190 VDD.n1180 9.3005
R16378 VDD.n1192 VDD.n1191 9.3005
R16379 VDD.n1193 VDD.n1179 9.3005
R16380 VDD.n1195 VDD.n1194 9.3005
R16381 VDD.n1196 VDD.n1172 9.3005
R16382 VDD.n1198 VDD.n1197 9.3005
R16383 VDD.n1199 VDD.n1171 9.3005
R16384 VDD.n1201 VDD.n1200 9.3005
R16385 VDD.n1202 VDD.n1164 9.3005
R16386 VDD.n1204 VDD.n1203 9.3005
R16387 VDD.n1205 VDD.n1163 9.3005
R16388 VDD.n1207 VDD.n1206 9.3005
R16389 VDD.n1208 VDD.n1153 9.3005
R16390 VDD.n1210 VDD.n1209 9.3005
R16391 VDD.n1211 VDD.n1152 9.3005
R16392 VDD.n1213 VDD.n1212 9.3005
R16393 VDD.n1214 VDD.n1145 9.3005
R16394 VDD.n1216 VDD.n1215 9.3005
R16395 VDD.n1217 VDD.n1144 9.3005
R16396 VDD.n1219 VDD.n1218 9.3005
R16397 VDD.n1220 VDD.n1137 9.3005
R16398 VDD.n1222 VDD.n1221 9.3005
R16399 VDD.n1223 VDD.n1136 9.3005
R16400 VDD.n1225 VDD.n1224 9.3005
R16401 VDD.n1226 VDD.n1129 9.3005
R16402 VDD.n1228 VDD.n1227 9.3005
R16403 VDD.n1229 VDD.n1128 9.3005
R16404 VDD.n1231 VDD.n1230 9.3005
R16405 VDD.n1237 VDD.n1236 9.3005
R16406 VDD.n1238 VDD.n1120 9.3005
R16407 VDD.n1240 VDD.n1239 9.3005
R16408 VDD.n1241 VDD.n1113 9.3005
R16409 VDD.n1243 VDD.n1242 9.3005
R16410 VDD.n1244 VDD.n1112 9.3005
R16411 VDD.n1246 VDD.n1245 9.3005
R16412 VDD.n1247 VDD.n1105 9.3005
R16413 VDD.n1249 VDD.n1248 9.3005
R16414 VDD.n1250 VDD.n1104 9.3005
R16415 VDD.n1252 VDD.n1251 9.3005
R16416 VDD.n1253 VDD.n1097 9.3005
R16417 VDD.n1255 VDD.n1254 9.3005
R16418 VDD.n1258 VDD.n1257 9.3005
R16419 VDD.n1259 VDD.n1087 9.3005
R16420 VDD.n1261 VDD.n1260 9.3005
R16421 VDD.n1262 VDD.n1086 9.3005
R16422 VDD.n1264 VDD.n1263 9.3005
R16423 VDD.n1265 VDD.n1079 9.3005
R16424 VDD.n1267 VDD.n1266 9.3005
R16425 VDD.n1268 VDD.n1078 9.3005
R16426 VDD.n1270 VDD.n1269 9.3005
R16427 VDD.n1271 VDD.n1074 9.3005
R16428 VDD.n1273 VDD.n1272 9.3005
R16429 VDD.n1256 VDD.n1096 9.3005
R16430 VDD.n1235 VDD.n1121 9.3005
R16431 VDD.n1186 VDD.n1070 9.3005
R16432 VDD.n1065 VDD.n1064 9.3005
R16433 VDD.n1288 VDD.n1287 9.3005
R16434 VDD.n1289 VDD.n1063 9.3005
R16435 VDD.n1291 VDD.n1290 9.3005
R16436 VDD.n1053 VDD.n1052 9.3005
R16437 VDD.n1304 VDD.n1303 9.3005
R16438 VDD.n1305 VDD.n1051 9.3005
R16439 VDD.n1307 VDD.n1306 9.3005
R16440 VDD.n1041 VDD.n1040 9.3005
R16441 VDD.n1320 VDD.n1319 9.3005
R16442 VDD.n1321 VDD.n1039 9.3005
R16443 VDD.n1323 VDD.n1322 9.3005
R16444 VDD.n1029 VDD.n1028 9.3005
R16445 VDD.n1336 VDD.n1335 9.3005
R16446 VDD.n1337 VDD.n1027 9.3005
R16447 VDD.n1339 VDD.n1338 9.3005
R16448 VDD.n1017 VDD.n1016 9.3005
R16449 VDD.n1352 VDD.n1351 9.3005
R16450 VDD.n1353 VDD.n1015 9.3005
R16451 VDD.n1355 VDD.n1354 9.3005
R16452 VDD.n1005 VDD.n1004 9.3005
R16453 VDD.n1368 VDD.n1367 9.3005
R16454 VDD.n1369 VDD.n1003 9.3005
R16455 VDD.n1371 VDD.n1370 9.3005
R16456 VDD.n993 VDD.n992 9.3005
R16457 VDD.n1275 VDD.n1274 9.3005
R16458 VDD.n1395 VDD.n1382 9.3005
R16459 VDD.n15 VDD.n14 8.34415
R16460 VDD.n2780 VDD.n2779 8.07387
R16461 VDD.n1395 VDD.n1394 8.07387
R16462 VDD.n586 VDD.t26 7.50544
R16463 VDD.t34 VDD.n513 7.50544
R16464 VDD.n1254 VDD.n1096 7.17626
R16465 VDD.n2701 VDD.n124 7.17626
R16466 VDD.n2451 VDD.n2450 7.17626
R16467 VDD.n688 VDD.t40 6.88003
R16468 VDD.t28 VDD.n609 6.88003
R16469 VDD.n491 VDD.t21 6.88003
R16470 VDD.t44 VDD.n411 6.88003
R16471 VDD.n1234 VDD.n1231 6.4005
R16472 VDD.n1574 VDD.n1571 6.4005
R16473 VDD.n2678 VDD.n2675 6.4005
R16474 VDD.n2422 VDD.n341 6.4005
R16475 VDD.n1387 VDD.n1384 6.29217
R16476 VDD.n20 VDD.n17 5.64705
R16477 VDD.t123 VDD.n674 5.6292
R16478 VDD.n593 VDD.t79 5.6292
R16479 VDD.t53 VDD.n507 5.6292
R16480 VDD.n426 VDD.t75 5.6292
R16481 VDD.n1209 VDD.n1156 5.62474
R16482 VDD.n1545 VDD.n780 5.62474
R16483 VDD.n2649 VDD.n178 5.62474
R16484 VDD.n2396 VDD.n2393 5.62474
R16485 VDD.n1690 VDD.n1689 5.30782
R16486 VDD.n1689 VDD.n1688 5.30782
R16487 VDD.n2308 VDD.n2307 5.30782
R16488 VDD.n2307 VDD.n2306 5.30782
R16489 VDD.n2346 VDD.n369 5.30782
R16490 VDD.n2346 VDD.n2345 5.30782
R16491 VDD.n884 VDD.n798 5.30782
R16492 VDD.n884 VDD.n883 5.30782
R16493 VDD.n1393 VDD.n1392 5.28355
R16494 VDD.n1390 VDD.n1389 5.28355
R16495 VDD.n1387 VDD.n1386 5.28355
R16496 VDD.n1729 VDD.t123 5.00379
R16497 VDD.n1824 VDD.t79 5.00379
R16498 VDD.n2154 VDD.t53 5.00379
R16499 VDD.n2249 VDD.t75 5.00379
R16500 VDD.n1189 VDD.n1186 4.84898
R16501 VDD.n1527 VDD.n910 4.84898
R16502 VDD.n2626 VDD.n2623 4.84898
R16503 VDD.n2366 VDD.n2363 4.84898
R16504 VDD.n1543 VDD.n1542 4.74817
R16505 VDD.n890 VDD.n885 4.74817
R16506 VDD.n1605 VDD.n1604 4.74817
R16507 VDD.n1605 VDD.n724 4.74817
R16508 VDD.n2386 VDD.n366 4.74817
R16509 VDD.n2384 VDD.n2383 4.74817
R16510 VDD.n2384 VDD.n2347 4.74817
R16511 VDD.n2387 VDD.n2386 4.74817
R16512 VDD.n1542 VDD.n786 4.74817
R16513 VDD.n887 VDD.n885 4.74817
R16514 VDD.n2452 VDD.n2451 4.67736
R16515 VDD.n2453 VDD.n2452 4.67736
R16516 VDD.n26 VDD.n25 4.63843
R16517 VDD.n23 VDD.n22 4.63843
R16518 VDD.n20 VDD.n19 4.63843
R16519 VDD.n2780 VDD.n26 4.28111
R16520 VDD.n1394 VDD.n1393 4.28111
R16521 VDD.n1729 VDD.t40 3.75297
R16522 VDD.n1794 VDD.t28 3.75297
R16523 VDD.n2184 VDD.t21 3.75297
R16524 VDD.n2249 VDD.t44 3.75297
R16525 VDD.n1606 VDD.n723 3.35648
R16526 VDD.n1061 VDD.t68 3.12756
R16527 VDD.t61 VDD.n929 3.12756
R16528 VDD.n1835 VDD.t26 3.12756
R16529 VDD.n2148 VDD.t34 3.12756
R16530 VDD.n287 VDD.t83 3.12756
R16531 VDD.t57 VDD.n2736 3.12756
R16532 VDD.n730 VDD.n723 2.59004
R16533 VDD.n1597 VDD.n723 2.59004
R16534 VDD.n2452 VDD.n314 2.31282
R16535 VDD.n1606 VDD.n1605 2.27742
R16536 VDD.n2385 VDD.n2384 2.27742
R16537 VDD.n2386 VDD.n2385 2.27742
R16538 VDD.n1542 VDD.n1541 2.27742
R16539 VDD.n1541 VDD.n885 2.27742
R16540 VDD.n1394 VDD.n15 1.78948
R16541 VDD VDD.n2780 1.78164
R16542 VDD.n1190 VDD.n1189 1.74595
R16543 VDD.n910 VDD.n906 1.74595
R16544 VDD.n2627 VDD.n2626 1.74595
R16545 VDD.n2367 VDD.n2366 1.74595
R16546 VDD.n4 VDD.n2 1.36975
R16547 VDD.n11 VDD.n9 1.36975
R16548 VDD.n6 VDD.n4 1.1097
R16549 VDD.n13 VDD.n11 1.1097
R16550 VDD.n26 VDD.n23 1.00912
R16551 VDD.n23 VDD.n20 1.00912
R16552 VDD.n1393 VDD.n1390 1.00912
R16553 VDD.n1390 VDD.n1387 1.00912
R16554 VDD.n1156 VDD.n1152 0.970197
R16555 VDD.n780 VDD.n775 0.970197
R16556 VDD.n178 VDD.n173 0.970197
R16557 VDD.n2397 VDD.n2396 0.970197
R16558 VDD.n14 VDD.n6 0.8755
R16559 VDD.n14 VDD.n13 0.8755
R16560 VDD.n1854 VDD.n569 0.62489
R16561 VDD.n1680 VDD.n1679 0.62489
R16562 VDD.n2105 VDD.n2104 0.62489
R16563 VDD.n2299 VDD.n2298 0.62489
R16564 VDD.n2337 VDD.n2336 0.62489
R16565 VDD.n2008 VDD.n1935 0.62489
R16566 VDD.n1894 VDD.n1893 0.62489
R16567 VDD.n875 VDD.n874 0.62489
R16568 VDD.n1521 VDD.n1520 0.474585
R16569 VDD.n2475 VDD.n2474 0.474585
R16570 VDD.n2724 VDD.n2723 0.474585
R16571 VDD.n2620 VDD.n2619 0.474585
R16572 VDD.n2481 VDD.n296 0.474585
R16573 VDD.n1528 VDD.n907 0.474585
R16574 VDD.n1280 VDD.n1070 0.474585
R16575 VDD.n1274 VDD.n1273 0.474585
R16576 VDD.n1025 VDD.t4 0.313206
R16577 VDD.t7 VDD.n965 0.313206
R16578 VDD.n251 VDD.t137 0.313206
R16579 VDD.t0 VDD.n2760 0.313206
R16580 VDD.n1235 VDD.n1234 0.194439
R16581 VDD.n1575 VDD.n1574 0.194439
R16582 VDD.n2679 VDD.n2678 0.194439
R16583 VDD.n341 VDD.n337 0.194439
R16584 VDD.n1397 VDD.n1396 0.152939
R16585 VDD.n1397 VDD.n980 0.152939
R16586 VDD.n1411 VDD.n980 0.152939
R16587 VDD.n1412 VDD.n1411 0.152939
R16588 VDD.n1413 VDD.n1412 0.152939
R16589 VDD.n1413 VDD.n968 0.152939
R16590 VDD.n1427 VDD.n968 0.152939
R16591 VDD.n1428 VDD.n1427 0.152939
R16592 VDD.n1429 VDD.n1428 0.152939
R16593 VDD.n1429 VDD.n956 0.152939
R16594 VDD.n1443 VDD.n956 0.152939
R16595 VDD.n1444 VDD.n1443 0.152939
R16596 VDD.n1445 VDD.n1444 0.152939
R16597 VDD.n1445 VDD.n944 0.152939
R16598 VDD.n1459 VDD.n944 0.152939
R16599 VDD.n1460 VDD.n1459 0.152939
R16600 VDD.n1461 VDD.n1460 0.152939
R16601 VDD.n1461 VDD.n932 0.152939
R16602 VDD.n1475 VDD.n932 0.152939
R16603 VDD.n1476 VDD.n1475 0.152939
R16604 VDD.n1477 VDD.n1476 0.152939
R16605 VDD.n1477 VDD.n919 0.152939
R16606 VDD.n1492 VDD.n919 0.152939
R16607 VDD.n1493 VDD.n1492 0.152939
R16608 VDD.n1521 VDD.n1493 0.152939
R16609 VDD.n1520 VDD.n1494 0.152939
R16610 VDD.n1498 VDD.n1494 0.152939
R16611 VDD.n1499 VDD.n1498 0.152939
R16612 VDD.n1500 VDD.n1499 0.152939
R16613 VDD.n1501 VDD.n1500 0.152939
R16614 VDD.n1502 VDD.n1501 0.152939
R16615 VDD.n1503 VDD.n1502 0.152939
R16616 VDD.n1503 VDD.n721 0.152939
R16617 VDD.n732 VDD.n722 0.152939
R16618 VDD.n736 VDD.n732 0.152939
R16619 VDD.n737 VDD.n736 0.152939
R16620 VDD.n738 VDD.n737 0.152939
R16621 VDD.n739 VDD.n738 0.152939
R16622 VDD.n743 VDD.n739 0.152939
R16623 VDD.n744 VDD.n743 0.152939
R16624 VDD.n745 VDD.n744 0.152939
R16625 VDD.n746 VDD.n745 0.152939
R16626 VDD.n750 VDD.n746 0.152939
R16627 VDD.n751 VDD.n750 0.152939
R16628 VDD.n752 VDD.n751 0.152939
R16629 VDD.n753 VDD.n752 0.152939
R16630 VDD.n757 VDD.n753 0.152939
R16631 VDD.n758 VDD.n757 0.152939
R16632 VDD.n759 VDD.n758 0.152939
R16633 VDD.n760 VDD.n759 0.152939
R16634 VDD.n764 VDD.n760 0.152939
R16635 VDD.n765 VDD.n764 0.152939
R16636 VDD.n766 VDD.n765 0.152939
R16637 VDD.n767 VDD.n766 0.152939
R16638 VDD.n771 VDD.n767 0.152939
R16639 VDD.n772 VDD.n771 0.152939
R16640 VDD.n773 VDD.n772 0.152939
R16641 VDD.n774 VDD.n773 0.152939
R16642 VDD.n781 VDD.n774 0.152939
R16643 VDD.n782 VDD.n781 0.152939
R16644 VDD.n783 VDD.n782 0.152939
R16645 VDD.n322 VDD.n319 0.152939
R16646 VDD.n323 VDD.n322 0.152939
R16647 VDD.n324 VDD.n323 0.152939
R16648 VDD.n327 VDD.n324 0.152939
R16649 VDD.n328 VDD.n327 0.152939
R16650 VDD.n329 VDD.n328 0.152939
R16651 VDD.n330 VDD.n329 0.152939
R16652 VDD.n333 VDD.n330 0.152939
R16653 VDD.n334 VDD.n333 0.152939
R16654 VDD.n335 VDD.n334 0.152939
R16655 VDD.n336 VDD.n335 0.152939
R16656 VDD.n342 VDD.n336 0.152939
R16657 VDD.n343 VDD.n342 0.152939
R16658 VDD.n344 VDD.n343 0.152939
R16659 VDD.n345 VDD.n344 0.152939
R16660 VDD.n348 VDD.n345 0.152939
R16661 VDD.n349 VDD.n348 0.152939
R16662 VDD.n350 VDD.n349 0.152939
R16663 VDD.n351 VDD.n350 0.152939
R16664 VDD.n354 VDD.n351 0.152939
R16665 VDD.n355 VDD.n354 0.152939
R16666 VDD.n356 VDD.n355 0.152939
R16667 VDD.n357 VDD.n356 0.152939
R16668 VDD.n360 VDD.n357 0.152939
R16669 VDD.n361 VDD.n360 0.152939
R16670 VDD.n362 VDD.n361 0.152939
R16671 VDD.n363 VDD.n362 0.152939
R16672 VDD.n367 VDD.n363 0.152939
R16673 VDD.n2474 VDD.n300 0.152939
R16674 VDD.n303 VDD.n300 0.152939
R16675 VDD.n304 VDD.n303 0.152939
R16676 VDD.n305 VDD.n304 0.152939
R16677 VDD.n308 VDD.n305 0.152939
R16678 VDD.n309 VDD.n308 0.152939
R16679 VDD.n310 VDD.n309 0.152939
R16680 VDD.n311 VDD.n310 0.152939
R16681 VDD.n2475 VDD.n290 0.152939
R16682 VDD.n2489 VDD.n290 0.152939
R16683 VDD.n2490 VDD.n2489 0.152939
R16684 VDD.n2491 VDD.n2490 0.152939
R16685 VDD.n2491 VDD.n278 0.152939
R16686 VDD.n2505 VDD.n278 0.152939
R16687 VDD.n2506 VDD.n2505 0.152939
R16688 VDD.n2507 VDD.n2506 0.152939
R16689 VDD.n2507 VDD.n266 0.152939
R16690 VDD.n2521 VDD.n266 0.152939
R16691 VDD.n2522 VDD.n2521 0.152939
R16692 VDD.n2523 VDD.n2522 0.152939
R16693 VDD.n2523 VDD.n254 0.152939
R16694 VDD.n2537 VDD.n254 0.152939
R16695 VDD.n2538 VDD.n2537 0.152939
R16696 VDD.n2539 VDD.n2538 0.152939
R16697 VDD.n2539 VDD.n242 0.152939
R16698 VDD.n2553 VDD.n242 0.152939
R16699 VDD.n2554 VDD.n2553 0.152939
R16700 VDD.n2555 VDD.n2554 0.152939
R16701 VDD.n2555 VDD.n230 0.152939
R16702 VDD.n2569 VDD.n230 0.152939
R16703 VDD.n2570 VDD.n2569 0.152939
R16704 VDD.n2571 VDD.n2570 0.152939
R16705 VDD.n2571 VDD.n27 0.152939
R16706 VDD.n39 VDD.n28 0.152939
R16707 VDD.n40 VDD.n39 0.152939
R16708 VDD.n41 VDD.n40 0.152939
R16709 VDD.n49 VDD.n41 0.152939
R16710 VDD.n50 VDD.n49 0.152939
R16711 VDD.n51 VDD.n50 0.152939
R16712 VDD.n52 VDD.n51 0.152939
R16713 VDD.n60 VDD.n52 0.152939
R16714 VDD.n61 VDD.n60 0.152939
R16715 VDD.n62 VDD.n61 0.152939
R16716 VDD.n63 VDD.n62 0.152939
R16717 VDD.n71 VDD.n63 0.152939
R16718 VDD.n72 VDD.n71 0.152939
R16719 VDD.n73 VDD.n72 0.152939
R16720 VDD.n74 VDD.n73 0.152939
R16721 VDD.n82 VDD.n74 0.152939
R16722 VDD.n83 VDD.n82 0.152939
R16723 VDD.n84 VDD.n83 0.152939
R16724 VDD.n85 VDD.n84 0.152939
R16725 VDD.n93 VDD.n85 0.152939
R16726 VDD.n94 VDD.n93 0.152939
R16727 VDD.n95 VDD.n94 0.152939
R16728 VDD.n96 VDD.n95 0.152939
R16729 VDD.n104 VDD.n96 0.152939
R16730 VDD.n2724 VDD.n104 0.152939
R16731 VDD.n2723 VDD.n105 0.152939
R16732 VDD.n107 VDD.n105 0.152939
R16733 VDD.n111 VDD.n107 0.152939
R16734 VDD.n112 VDD.n111 0.152939
R16735 VDD.n113 VDD.n112 0.152939
R16736 VDD.n114 VDD.n113 0.152939
R16737 VDD.n118 VDD.n114 0.152939
R16738 VDD.n119 VDD.n118 0.152939
R16739 VDD.n120 VDD.n119 0.152939
R16740 VDD.n121 VDD.n120 0.152939
R16741 VDD.n127 VDD.n121 0.152939
R16742 VDD.n128 VDD.n127 0.152939
R16743 VDD.n129 VDD.n128 0.152939
R16744 VDD.n130 VDD.n129 0.152939
R16745 VDD.n134 VDD.n130 0.152939
R16746 VDD.n135 VDD.n134 0.152939
R16747 VDD.n136 VDD.n135 0.152939
R16748 VDD.n137 VDD.n136 0.152939
R16749 VDD.n141 VDD.n137 0.152939
R16750 VDD.n142 VDD.n141 0.152939
R16751 VDD.n143 VDD.n142 0.152939
R16752 VDD.n144 VDD.n143 0.152939
R16753 VDD.n148 VDD.n144 0.152939
R16754 VDD.n149 VDD.n148 0.152939
R16755 VDD.n150 VDD.n149 0.152939
R16756 VDD.n151 VDD.n150 0.152939
R16757 VDD.n155 VDD.n151 0.152939
R16758 VDD.n156 VDD.n155 0.152939
R16759 VDD.n157 VDD.n156 0.152939
R16760 VDD.n158 VDD.n157 0.152939
R16761 VDD.n162 VDD.n158 0.152939
R16762 VDD.n163 VDD.n162 0.152939
R16763 VDD.n164 VDD.n163 0.152939
R16764 VDD.n165 VDD.n164 0.152939
R16765 VDD.n169 VDD.n165 0.152939
R16766 VDD.n170 VDD.n169 0.152939
R16767 VDD.n171 VDD.n170 0.152939
R16768 VDD.n172 VDD.n171 0.152939
R16769 VDD.n179 VDD.n172 0.152939
R16770 VDD.n180 VDD.n179 0.152939
R16771 VDD.n181 VDD.n180 0.152939
R16772 VDD.n182 VDD.n181 0.152939
R16773 VDD.n186 VDD.n182 0.152939
R16774 VDD.n187 VDD.n186 0.152939
R16775 VDD.n188 VDD.n187 0.152939
R16776 VDD.n189 VDD.n188 0.152939
R16777 VDD.n193 VDD.n189 0.152939
R16778 VDD.n194 VDD.n193 0.152939
R16779 VDD.n195 VDD.n194 0.152939
R16780 VDD.n196 VDD.n195 0.152939
R16781 VDD.n200 VDD.n196 0.152939
R16782 VDD.n201 VDD.n200 0.152939
R16783 VDD.n202 VDD.n201 0.152939
R16784 VDD.n2620 VDD.n202 0.152939
R16785 VDD.n2482 VDD.n2481 0.152939
R16786 VDD.n2483 VDD.n2482 0.152939
R16787 VDD.n2483 VDD.n283 0.152939
R16788 VDD.n2497 VDD.n283 0.152939
R16789 VDD.n2498 VDD.n2497 0.152939
R16790 VDD.n2499 VDD.n2498 0.152939
R16791 VDD.n2499 VDD.n272 0.152939
R16792 VDD.n2513 VDD.n272 0.152939
R16793 VDD.n2514 VDD.n2513 0.152939
R16794 VDD.n2515 VDD.n2514 0.152939
R16795 VDD.n2515 VDD.n260 0.152939
R16796 VDD.n2529 VDD.n260 0.152939
R16797 VDD.n2530 VDD.n2529 0.152939
R16798 VDD.n2531 VDD.n2530 0.152939
R16799 VDD.n2531 VDD.n247 0.152939
R16800 VDD.n2545 VDD.n247 0.152939
R16801 VDD.n2546 VDD.n2545 0.152939
R16802 VDD.n2547 VDD.n2546 0.152939
R16803 VDD.n2547 VDD.n236 0.152939
R16804 VDD.n2561 VDD.n236 0.152939
R16805 VDD.n2562 VDD.n2561 0.152939
R16806 VDD.n2563 VDD.n2562 0.152939
R16807 VDD.n2563 VDD.n223 0.152939
R16808 VDD.n2577 VDD.n223 0.152939
R16809 VDD.n2578 VDD.n2577 0.152939
R16810 VDD.n2579 VDD.n2578 0.152939
R16811 VDD.n2579 VDD.n221 0.152939
R16812 VDD.n2583 VDD.n221 0.152939
R16813 VDD.n2584 VDD.n2583 0.152939
R16814 VDD.n2585 VDD.n2584 0.152939
R16815 VDD.n2585 VDD.n218 0.152939
R16816 VDD.n2589 VDD.n218 0.152939
R16817 VDD.n2590 VDD.n2589 0.152939
R16818 VDD.n2591 VDD.n2590 0.152939
R16819 VDD.n2591 VDD.n215 0.152939
R16820 VDD.n2595 VDD.n215 0.152939
R16821 VDD.n2596 VDD.n2595 0.152939
R16822 VDD.n2597 VDD.n2596 0.152939
R16823 VDD.n2597 VDD.n212 0.152939
R16824 VDD.n2601 VDD.n212 0.152939
R16825 VDD.n2602 VDD.n2601 0.152939
R16826 VDD.n2603 VDD.n2602 0.152939
R16827 VDD.n2603 VDD.n209 0.152939
R16828 VDD.n2607 VDD.n209 0.152939
R16829 VDD.n2608 VDD.n2607 0.152939
R16830 VDD.n2609 VDD.n2608 0.152939
R16831 VDD.n2609 VDD.n206 0.152939
R16832 VDD.n2613 VDD.n206 0.152939
R16833 VDD.n2614 VDD.n2613 0.152939
R16834 VDD.n2615 VDD.n2614 0.152939
R16835 VDD.n2615 VDD.n203 0.152939
R16836 VDD.n2619 VDD.n203 0.152939
R16837 VDD.n2353 VDD.n368 0.152939
R16838 VDD.n2354 VDD.n2353 0.152939
R16839 VDD.n2355 VDD.n2354 0.152939
R16840 VDD.n2356 VDD.n2355 0.152939
R16841 VDD.n2360 VDD.n2356 0.152939
R16842 VDD.n2361 VDD.n2360 0.152939
R16843 VDD.n2362 VDD.n2361 0.152939
R16844 VDD.n2362 VDD.n296 0.152939
R16845 VDD.n1540 VDD.n886 0.152939
R16846 VDD.n1536 VDD.n886 0.152939
R16847 VDD.n1536 VDD.n1535 0.152939
R16848 VDD.n1535 VDD.n1534 0.152939
R16849 VDD.n1534 VDD.n899 0.152939
R16850 VDD.n1530 VDD.n899 0.152939
R16851 VDD.n1530 VDD.n1529 0.152939
R16852 VDD.n1529 VDD.n1528 0.152939
R16853 VDD.n1281 VDD.n1280 0.152939
R16854 VDD.n1282 VDD.n1281 0.152939
R16855 VDD.n1282 VDD.n1057 0.152939
R16856 VDD.n1296 VDD.n1057 0.152939
R16857 VDD.n1297 VDD.n1296 0.152939
R16858 VDD.n1298 VDD.n1297 0.152939
R16859 VDD.n1298 VDD.n1046 0.152939
R16860 VDD.n1312 VDD.n1046 0.152939
R16861 VDD.n1313 VDD.n1312 0.152939
R16862 VDD.n1314 VDD.n1313 0.152939
R16863 VDD.n1314 VDD.n1034 0.152939
R16864 VDD.n1328 VDD.n1034 0.152939
R16865 VDD.n1329 VDD.n1328 0.152939
R16866 VDD.n1330 VDD.n1329 0.152939
R16867 VDD.n1330 VDD.n1021 0.152939
R16868 VDD.n1344 VDD.n1021 0.152939
R16869 VDD.n1345 VDD.n1344 0.152939
R16870 VDD.n1346 VDD.n1345 0.152939
R16871 VDD.n1346 VDD.n1010 0.152939
R16872 VDD.n1360 VDD.n1010 0.152939
R16873 VDD.n1361 VDD.n1360 0.152939
R16874 VDD.n1362 VDD.n1361 0.152939
R16875 VDD.n1362 VDD.n998 0.152939
R16876 VDD.n1376 VDD.n998 0.152939
R16877 VDD.n1377 VDD.n1376 0.152939
R16878 VDD.n1378 VDD.n1377 0.152939
R16879 VDD.n1378 VDD.n986 0.152939
R16880 VDD.n1403 VDD.n986 0.152939
R16881 VDD.n1404 VDD.n1403 0.152939
R16882 VDD.n1405 VDD.n1404 0.152939
R16883 VDD.n1405 VDD.n974 0.152939
R16884 VDD.n1419 VDD.n974 0.152939
R16885 VDD.n1420 VDD.n1419 0.152939
R16886 VDD.n1421 VDD.n1420 0.152939
R16887 VDD.n1421 VDD.n962 0.152939
R16888 VDD.n1435 VDD.n962 0.152939
R16889 VDD.n1436 VDD.n1435 0.152939
R16890 VDD.n1437 VDD.n1436 0.152939
R16891 VDD.n1437 VDD.n950 0.152939
R16892 VDD.n1451 VDD.n950 0.152939
R16893 VDD.n1452 VDD.n1451 0.152939
R16894 VDD.n1453 VDD.n1452 0.152939
R16895 VDD.n1453 VDD.n938 0.152939
R16896 VDD.n1467 VDD.n938 0.152939
R16897 VDD.n1468 VDD.n1467 0.152939
R16898 VDD.n1469 VDD.n1468 0.152939
R16899 VDD.n1469 VDD.n926 0.152939
R16900 VDD.n1483 VDD.n926 0.152939
R16901 VDD.n1484 VDD.n1483 0.152939
R16902 VDD.n1486 VDD.n1484 0.152939
R16903 VDD.n1486 VDD.n1485 0.152939
R16904 VDD.n1485 VDD.n907 0.152939
R16905 VDD.n1273 VDD.n1074 0.152939
R16906 VDD.n1269 VDD.n1074 0.152939
R16907 VDD.n1269 VDD.n1268 0.152939
R16908 VDD.n1268 VDD.n1267 0.152939
R16909 VDD.n1267 VDD.n1079 0.152939
R16910 VDD.n1263 VDD.n1079 0.152939
R16911 VDD.n1263 VDD.n1262 0.152939
R16912 VDD.n1262 VDD.n1261 0.152939
R16913 VDD.n1261 VDD.n1087 0.152939
R16914 VDD.n1257 VDD.n1087 0.152939
R16915 VDD.n1257 VDD.n1256 0.152939
R16916 VDD.n1256 VDD.n1255 0.152939
R16917 VDD.n1255 VDD.n1097 0.152939
R16918 VDD.n1251 VDD.n1097 0.152939
R16919 VDD.n1251 VDD.n1250 0.152939
R16920 VDD.n1250 VDD.n1249 0.152939
R16921 VDD.n1249 VDD.n1105 0.152939
R16922 VDD.n1245 VDD.n1105 0.152939
R16923 VDD.n1245 VDD.n1244 0.152939
R16924 VDD.n1244 VDD.n1243 0.152939
R16925 VDD.n1243 VDD.n1113 0.152939
R16926 VDD.n1239 VDD.n1113 0.152939
R16927 VDD.n1239 VDD.n1238 0.152939
R16928 VDD.n1238 VDD.n1237 0.152939
R16929 VDD.n1237 VDD.n1121 0.152939
R16930 VDD.n1230 VDD.n1121 0.152939
R16931 VDD.n1230 VDD.n1229 0.152939
R16932 VDD.n1229 VDD.n1228 0.152939
R16933 VDD.n1228 VDD.n1129 0.152939
R16934 VDD.n1224 VDD.n1129 0.152939
R16935 VDD.n1224 VDD.n1223 0.152939
R16936 VDD.n1223 VDD.n1222 0.152939
R16937 VDD.n1222 VDD.n1137 0.152939
R16938 VDD.n1218 VDD.n1137 0.152939
R16939 VDD.n1218 VDD.n1217 0.152939
R16940 VDD.n1217 VDD.n1216 0.152939
R16941 VDD.n1216 VDD.n1145 0.152939
R16942 VDD.n1212 VDD.n1145 0.152939
R16943 VDD.n1212 VDD.n1211 0.152939
R16944 VDD.n1211 VDD.n1210 0.152939
R16945 VDD.n1210 VDD.n1153 0.152939
R16946 VDD.n1206 VDD.n1153 0.152939
R16947 VDD.n1206 VDD.n1205 0.152939
R16948 VDD.n1205 VDD.n1204 0.152939
R16949 VDD.n1204 VDD.n1164 0.152939
R16950 VDD.n1200 VDD.n1164 0.152939
R16951 VDD.n1200 VDD.n1199 0.152939
R16952 VDD.n1199 VDD.n1198 0.152939
R16953 VDD.n1198 VDD.n1172 0.152939
R16954 VDD.n1194 VDD.n1172 0.152939
R16955 VDD.n1194 VDD.n1193 0.152939
R16956 VDD.n1193 VDD.n1192 0.152939
R16957 VDD.n1192 VDD.n1180 0.152939
R16958 VDD.n1180 VDD.n1070 0.152939
R16959 VDD.n1274 VDD.n1064 0.152939
R16960 VDD.n1288 VDD.n1064 0.152939
R16961 VDD.n1289 VDD.n1288 0.152939
R16962 VDD.n1290 VDD.n1289 0.152939
R16963 VDD.n1290 VDD.n1052 0.152939
R16964 VDD.n1304 VDD.n1052 0.152939
R16965 VDD.n1305 VDD.n1304 0.152939
R16966 VDD.n1306 VDD.n1305 0.152939
R16967 VDD.n1306 VDD.n1040 0.152939
R16968 VDD.n1320 VDD.n1040 0.152939
R16969 VDD.n1321 VDD.n1320 0.152939
R16970 VDD.n1322 VDD.n1321 0.152939
R16971 VDD.n1322 VDD.n1028 0.152939
R16972 VDD.n1336 VDD.n1028 0.152939
R16973 VDD.n1337 VDD.n1336 0.152939
R16974 VDD.n1338 VDD.n1337 0.152939
R16975 VDD.n1338 VDD.n1016 0.152939
R16976 VDD.n1352 VDD.n1016 0.152939
R16977 VDD.n1353 VDD.n1352 0.152939
R16978 VDD.n1354 VDD.n1353 0.152939
R16979 VDD.n1354 VDD.n1004 0.152939
R16980 VDD.n1368 VDD.n1004 0.152939
R16981 VDD.n1369 VDD.n1368 0.152939
R16982 VDD.n1370 VDD.n1369 0.152939
R16983 VDD.n1370 VDD.n992 0.152939
R16984 VDD.n1396 VDD.n1395 0.145814
R16985 VDD.n2779 VDD.n27 0.145814
R16986 VDD.n2779 VDD.n28 0.145814
R16987 VDD.n1395 VDD.n992 0.145814
R16988 VDD.n1606 VDD.n721 0.0797683
R16989 VDD.n314 VDD.n311 0.0797683
R16990 VDD.n2385 VDD.n368 0.0797683
R16991 VDD.n1541 VDD.n1540 0.0797683
R16992 VDD.n1606 VDD.n722 0.0736707
R16993 VDD.n1541 VDD.n783 0.0736707
R16994 VDD.n319 VDD.n314 0.0736707
R16995 VDD.n2385 VDD.n367 0.0736707
R16996 VDD VDD.n15 0.00833333
R16997 VOUT.n27 VOUT.t40 136.179
R16998 VOUT.n24 VOUT.t39 136.179
R16999 VOUT.n21 VOUT.t38 136.179
R17000 VOUT.n19 VOUT.t41 136.179
R17001 VOUT.n9 VOUT.t14 134.888
R17002 VOUT.n6 VOUT.t36 134.888
R17003 VOUT.n3 VOUT.t6 134.888
R17004 VOUT.n1 VOUT.t27 134.888
R17005 VOUT.n9 VOUT.n8 118.07
R17006 VOUT.n6 VOUT.n5 118.07
R17007 VOUT.n3 VOUT.n2 118.07
R17008 VOUT.n1 VOUT.n0 118.07
R17009 VOUT.n24 VOUT.n23 116.781
R17010 VOUT.n21 VOUT.n20 116.781
R17011 VOUT.n19 VOUT.n18 116.781
R17012 VOUT.n27 VOUT.n26 116.781
R17013 VOUT.n37 VOUT.n35 65.6555
R17014 VOUT.n32 VOUT.n30 65.6555
R17015 VOUT.n49 VOUT.n47 65.6555
R17016 VOUT.n44 VOUT.n42 65.6555
R17017 VOUT.n39 VOUT.n38 64.8595
R17018 VOUT.n37 VOUT.n36 64.8595
R17019 VOUT.n34 VOUT.n33 64.8595
R17020 VOUT.n32 VOUT.n31 64.8595
R17021 VOUT.n49 VOUT.n48 64.8595
R17022 VOUT.n51 VOUT.n50 64.8595
R17023 VOUT.n44 VOUT.n43 64.8595
R17024 VOUT.n46 VOUT.n45 64.8595
R17025 VOUT.n26 VOUT.t10 18.1091
R17026 VOUT.n26 VOUT.t28 18.1091
R17027 VOUT.n23 VOUT.t11 18.1091
R17028 VOUT.n23 VOUT.t24 18.1091
R17029 VOUT.n20 VOUT.t5 18.1091
R17030 VOUT.n20 VOUT.t1 18.1091
R17031 VOUT.n18 VOUT.t7 18.1091
R17032 VOUT.n18 VOUT.t44 18.1091
R17033 VOUT.n8 VOUT.t32 18.1091
R17034 VOUT.n8 VOUT.t42 18.1091
R17035 VOUT.n5 VOUT.t20 18.1091
R17036 VOUT.n5 VOUT.t37 18.1091
R17037 VOUT.n2 VOUT.t43 18.1091
R17038 VOUT.n2 VOUT.t8 18.1091
R17039 VOUT.n0 VOUT.t12 18.1091
R17040 VOUT.n0 VOUT.t9 18.1091
R17041 VOUT.n41 VOUT.n29 9.01748
R17042 VOUT.n38 VOUT.t17 7.44411
R17043 VOUT.n38 VOUT.t0 7.44411
R17044 VOUT.n36 VOUT.t30 7.44411
R17045 VOUT.n36 VOUT.t21 7.44411
R17046 VOUT.n35 VOUT.t35 7.44411
R17047 VOUT.n35 VOUT.t16 7.44411
R17048 VOUT.n33 VOUT.t18 7.44411
R17049 VOUT.n33 VOUT.t15 7.44411
R17050 VOUT.n31 VOUT.t13 7.44411
R17051 VOUT.n31 VOUT.t45 7.44411
R17052 VOUT.n30 VOUT.t23 7.44411
R17053 VOUT.n30 VOUT.t47 7.44411
R17054 VOUT.n47 VOUT.t33 7.44411
R17055 VOUT.n47 VOUT.t4 7.44411
R17056 VOUT.n48 VOUT.t3 7.44411
R17057 VOUT.n48 VOUT.t22 7.44411
R17058 VOUT.n50 VOUT.t26 7.44411
R17059 VOUT.n50 VOUT.t19 7.44411
R17060 VOUT.n42 VOUT.t25 7.44411
R17061 VOUT.n42 VOUT.t34 7.44411
R17062 VOUT.n43 VOUT.t29 7.44411
R17063 VOUT.n43 VOUT.t2 7.44411
R17064 VOUT.n45 VOUT.t31 7.44411
R17065 VOUT.n45 VOUT.t46 7.44411
R17066 VOUT.n22 VOUT.n19 6.46458
R17067 VOUT.n40 VOUT.n34 6.46458
R17068 VOUT.n52 VOUT.n46 6.46458
R17069 VOUT.n4 VOUT.n1 5.81947
R17070 VOUT.n28 VOUT.n27 5.45596
R17071 VOUT.n25 VOUT.n24 5.45596
R17072 VOUT.n22 VOUT.n21 5.45596
R17073 VOUT.n41 VOUT.n40 5.40403
R17074 VOUT.n53 VOUT.n52 5.40403
R17075 VOUT.n40 VOUT.n39 5.20883
R17076 VOUT.n52 VOUT.n51 5.20883
R17077 VOUT.n10 VOUT.n9 4.81084
R17078 VOUT.n7 VOUT.n6 4.81084
R17079 VOUT.n4 VOUT.n3 4.81084
R17080 VOUT.n54 VOUT.n11 4.78067
R17081 VOUT.n17 VOUT 4.6018
R17082 VOUT.n29 VOUT.n28 4.39326
R17083 VOUT.n11 VOUT.n10 4.39326
R17084 VOUT.n29 VOUT.n11 4.23395
R17085 VOUT.n54 VOUT.n53 4.2178
R17086 VOUT.n53 VOUT.n41 3.18616
R17087 VOUT.n28 VOUT.n25 1.00912
R17088 VOUT.n25 VOUT.n22 1.00912
R17089 VOUT.n10 VOUT.n7 1.00912
R17090 VOUT.n7 VOUT.n4 1.00912
R17091 VOUT.n39 VOUT.n37 0.796477
R17092 VOUT.n34 VOUT.n32 0.796477
R17093 VOUT.n51 VOUT.n49 0.796477
R17094 VOUT.n46 VOUT.n44 0.796477
R17095 VOUT.n54 VOUT.n17 0.45123
R17096 VOUT.n17 VOUT.n16 0.4039
R17097 VOUT.n15 VOUT.n14 0.110766
R17098 VOUT.n13 VOUT.n12 0.107579
R17099 VOUT.n14 VOUT.n13 0.0591803
R17100 VOUT.n16 VOUT.n12 0.0540124
R17101 VOUT.n12 VOUT.t48 0.0143226
R17102 VOUT.n14 VOUT.t49 0.0134044
R17103 VOUT.n13 VOUT.t51 0.0133892
R17104 VOUT.n15 VOUT.t50 0.0118388
R17105 VOUT.n16 VOUT.n15 0.0112661
R17106 VOUT VOUT.n54 0.0099
R17107 CS_BIAS.n155 CS_BIAS.n107 161.3
R17108 CS_BIAS.n154 CS_BIAS.n153 161.3
R17109 CS_BIAS.n152 CS_BIAS.n108 161.3
R17110 CS_BIAS.n151 CS_BIAS.n150 161.3
R17111 CS_BIAS.n149 CS_BIAS.n109 161.3
R17112 CS_BIAS.n147 CS_BIAS.n146 161.3
R17113 CS_BIAS.n145 CS_BIAS.n110 161.3
R17114 CS_BIAS.n144 CS_BIAS.n143 161.3
R17115 CS_BIAS.n142 CS_BIAS.n111 161.3
R17116 CS_BIAS.n141 CS_BIAS.n140 161.3
R17117 CS_BIAS.n139 CS_BIAS.n112 161.3
R17118 CS_BIAS.n138 CS_BIAS.n137 161.3
R17119 CS_BIAS.n136 CS_BIAS.n113 161.3
R17120 CS_BIAS.n135 CS_BIAS.n134 161.3
R17121 CS_BIAS.n133 CS_BIAS.n115 161.3
R17122 CS_BIAS.n132 CS_BIAS.n131 161.3
R17123 CS_BIAS.n129 CS_BIAS.n116 161.3
R17124 CS_BIAS.n128 CS_BIAS.n127 161.3
R17125 CS_BIAS.n126 CS_BIAS.n117 161.3
R17126 CS_BIAS.n125 CS_BIAS.n124 161.3
R17127 CS_BIAS.n123 CS_BIAS.n118 161.3
R17128 CS_BIAS.n122 CS_BIAS.n121 161.3
R17129 CS_BIAS.n24 CS_BIAS.n23 161.3
R17130 CS_BIAS.n25 CS_BIAS.n20 161.3
R17131 CS_BIAS.n27 CS_BIAS.n26 161.3
R17132 CS_BIAS.n28 CS_BIAS.n19 161.3
R17133 CS_BIAS.n30 CS_BIAS.n29 161.3
R17134 CS_BIAS.n31 CS_BIAS.n18 161.3
R17135 CS_BIAS.n34 CS_BIAS.n33 161.3
R17136 CS_BIAS.n35 CS_BIAS.n17 161.3
R17137 CS_BIAS.n37 CS_BIAS.n36 161.3
R17138 CS_BIAS.n38 CS_BIAS.n15 161.3
R17139 CS_BIAS.n40 CS_BIAS.n39 161.3
R17140 CS_BIAS.n41 CS_BIAS.n14 161.3
R17141 CS_BIAS.n43 CS_BIAS.n42 161.3
R17142 CS_BIAS.n44 CS_BIAS.n13 161.3
R17143 CS_BIAS.n46 CS_BIAS.n45 161.3
R17144 CS_BIAS.n47 CS_BIAS.n12 161.3
R17145 CS_BIAS.n49 CS_BIAS.n48 161.3
R17146 CS_BIAS.n51 CS_BIAS.n11 161.3
R17147 CS_BIAS.n53 CS_BIAS.n52 161.3
R17148 CS_BIAS.n54 CS_BIAS.n10 161.3
R17149 CS_BIAS.n56 CS_BIAS.n55 161.3
R17150 CS_BIAS.n57 CS_BIAS.n9 161.3
R17151 CS_BIAS.n71 CS_BIAS.n70 161.3
R17152 CS_BIAS.n72 CS_BIAS.n67 161.3
R17153 CS_BIAS.n74 CS_BIAS.n73 161.3
R17154 CS_BIAS.n75 CS_BIAS.n66 161.3
R17155 CS_BIAS.n77 CS_BIAS.n76 161.3
R17156 CS_BIAS.n78 CS_BIAS.n65 161.3
R17157 CS_BIAS.n81 CS_BIAS.n80 161.3
R17158 CS_BIAS.n82 CS_BIAS.n8 161.3
R17159 CS_BIAS.n84 CS_BIAS.n83 161.3
R17160 CS_BIAS.n85 CS_BIAS.n6 161.3
R17161 CS_BIAS.n87 CS_BIAS.n86 161.3
R17162 CS_BIAS.n88 CS_BIAS.n5 161.3
R17163 CS_BIAS.n90 CS_BIAS.n89 161.3
R17164 CS_BIAS.n91 CS_BIAS.n4 161.3
R17165 CS_BIAS.n93 CS_BIAS.n92 161.3
R17166 CS_BIAS.n94 CS_BIAS.n3 161.3
R17167 CS_BIAS.n96 CS_BIAS.n95 161.3
R17168 CS_BIAS.n98 CS_BIAS.n2 161.3
R17169 CS_BIAS.n100 CS_BIAS.n99 161.3
R17170 CS_BIAS.n101 CS_BIAS.n1 161.3
R17171 CS_BIAS.n103 CS_BIAS.n102 161.3
R17172 CS_BIAS.n104 CS_BIAS.n0 161.3
R17173 CS_BIAS.n314 CS_BIAS.n266 161.3
R17174 CS_BIAS.n313 CS_BIAS.n312 161.3
R17175 CS_BIAS.n311 CS_BIAS.n267 161.3
R17176 CS_BIAS.n310 CS_BIAS.n309 161.3
R17177 CS_BIAS.n308 CS_BIAS.n268 161.3
R17178 CS_BIAS.n306 CS_BIAS.n305 161.3
R17179 CS_BIAS.n304 CS_BIAS.n269 161.3
R17180 CS_BIAS.n303 CS_BIAS.n302 161.3
R17181 CS_BIAS.n301 CS_BIAS.n270 161.3
R17182 CS_BIAS.n300 CS_BIAS.n299 161.3
R17183 CS_BIAS.n298 CS_BIAS.n271 161.3
R17184 CS_BIAS.n297 CS_BIAS.n296 161.3
R17185 CS_BIAS.n294 CS_BIAS.n272 161.3
R17186 CS_BIAS.n293 CS_BIAS.n292 161.3
R17187 CS_BIAS.n291 CS_BIAS.n273 161.3
R17188 CS_BIAS.n290 CS_BIAS.n289 161.3
R17189 CS_BIAS.n287 CS_BIAS.n274 161.3
R17190 CS_BIAS.n286 CS_BIAS.n285 161.3
R17191 CS_BIAS.n284 CS_BIAS.n275 161.3
R17192 CS_BIAS.n283 CS_BIAS.n282 161.3
R17193 CS_BIAS.n281 CS_BIAS.n276 161.3
R17194 CS_BIAS.n280 CS_BIAS.n279 161.3
R17195 CS_BIAS.n235 CS_BIAS.n187 161.3
R17196 CS_BIAS.n234 CS_BIAS.n233 161.3
R17197 CS_BIAS.n232 CS_BIAS.n188 161.3
R17198 CS_BIAS.n231 CS_BIAS.n230 161.3
R17199 CS_BIAS.n229 CS_BIAS.n189 161.3
R17200 CS_BIAS.n227 CS_BIAS.n226 161.3
R17201 CS_BIAS.n225 CS_BIAS.n190 161.3
R17202 CS_BIAS.n224 CS_BIAS.n223 161.3
R17203 CS_BIAS.n222 CS_BIAS.n191 161.3
R17204 CS_BIAS.n221 CS_BIAS.n220 161.3
R17205 CS_BIAS.n219 CS_BIAS.n192 161.3
R17206 CS_BIAS.n218 CS_BIAS.n217 161.3
R17207 CS_BIAS.n215 CS_BIAS.n193 161.3
R17208 CS_BIAS.n214 CS_BIAS.n213 161.3
R17209 CS_BIAS.n212 CS_BIAS.n194 161.3
R17210 CS_BIAS.n211 CS_BIAS.n210 161.3
R17211 CS_BIAS.n208 CS_BIAS.n195 161.3
R17212 CS_BIAS.n207 CS_BIAS.n206 161.3
R17213 CS_BIAS.n205 CS_BIAS.n196 161.3
R17214 CS_BIAS.n204 CS_BIAS.n203 161.3
R17215 CS_BIAS.n202 CS_BIAS.n197 161.3
R17216 CS_BIAS.n201 CS_BIAS.n200 161.3
R17217 CS_BIAS.n184 CS_BIAS.n166 161.3
R17218 CS_BIAS.n183 CS_BIAS.n182 161.3
R17219 CS_BIAS.n180 CS_BIAS.n167 161.3
R17220 CS_BIAS.n179 CS_BIAS.n178 161.3
R17221 CS_BIAS.n177 CS_BIAS.n168 161.3
R17222 CS_BIAS.n176 CS_BIAS.n175 161.3
R17223 CS_BIAS.n174 CS_BIAS.n169 161.3
R17224 CS_BIAS.n173 CS_BIAS.n172 161.3
R17225 CS_BIAS.n242 CS_BIAS.n241 161.3
R17226 CS_BIAS.n263 CS_BIAS.n159 161.3
R17227 CS_BIAS.n262 CS_BIAS.n261 161.3
R17228 CS_BIAS.n260 CS_BIAS.n160 161.3
R17229 CS_BIAS.n259 CS_BIAS.n258 161.3
R17230 CS_BIAS.n257 CS_BIAS.n161 161.3
R17231 CS_BIAS.n255 CS_BIAS.n254 161.3
R17232 CS_BIAS.n253 CS_BIAS.n162 161.3
R17233 CS_BIAS.n252 CS_BIAS.n251 161.3
R17234 CS_BIAS.n250 CS_BIAS.n163 161.3
R17235 CS_BIAS.n249 CS_BIAS.n248 161.3
R17236 CS_BIAS.n247 CS_BIAS.n164 161.3
R17237 CS_BIAS.n246 CS_BIAS.n245 161.3
R17238 CS_BIAS.n243 CS_BIAS.n165 161.3
R17239 CS_BIAS.n120 CS_BIAS.t35 96.8902
R17240 CS_BIAS.n22 CS_BIAS.t18 96.8902
R17241 CS_BIAS.n69 CS_BIAS.t47 96.8902
R17242 CS_BIAS.n278 CS_BIAS.t31 96.8902
R17243 CS_BIAS.n199 CS_BIAS.t20 96.8902
R17244 CS_BIAS.n171 CS_BIAS.t39 96.8902
R17245 CS_BIAS.n157 CS_BIAS.n156 90.0052
R17246 CS_BIAS.n59 CS_BIAS.n58 90.0052
R17247 CS_BIAS.n106 CS_BIAS.n105 90.0052
R17248 CS_BIAS.n316 CS_BIAS.n315 90.0052
R17249 CS_BIAS.n237 CS_BIAS.n236 90.0052
R17250 CS_BIAS.n265 CS_BIAS.n264 90.0052
R17251 CS_BIAS.n124 CS_BIAS.n117 73.0308
R17252 CS_BIAS.n143 CS_BIAS.n142 73.0308
R17253 CS_BIAS.n45 CS_BIAS.n44 73.0308
R17254 CS_BIAS.n26 CS_BIAS.n19 73.0308
R17255 CS_BIAS.n92 CS_BIAS.n91 73.0308
R17256 CS_BIAS.n73 CS_BIAS.n66 73.0308
R17257 CS_BIAS.n282 CS_BIAS.n275 73.0308
R17258 CS_BIAS.n302 CS_BIAS.n301 73.0308
R17259 CS_BIAS.n203 CS_BIAS.n196 73.0308
R17260 CS_BIAS.n223 CS_BIAS.n222 73.0308
R17261 CS_BIAS.n251 CS_BIAS.n250 73.0308
R17262 CS_BIAS.n175 CS_BIAS.n168 73.0308
R17263 CS_BIAS.n120 CS_BIAS.n119 68.9919
R17264 CS_BIAS.n22 CS_BIAS.n21 68.9919
R17265 CS_BIAS.n69 CS_BIAS.n68 68.9919
R17266 CS_BIAS.n278 CS_BIAS.n277 68.9919
R17267 CS_BIAS.n199 CS_BIAS.n198 68.9919
R17268 CS_BIAS.n171 CS_BIAS.n170 68.9919
R17269 CS_BIAS.n64 CS_BIAS.n63 65.6555
R17270 CS_BIAS.n240 CS_BIAS.n185 65.6555
R17271 CS_BIAS.n64 CS_BIAS.n62 64.8595
R17272 CS_BIAS.n61 CS_BIAS.n60 64.8595
R17273 CS_BIAS.n239 CS_BIAS.n238 64.8595
R17274 CS_BIAS.n240 CS_BIAS.n186 64.8595
R17275 CS_BIAS.n119 CS_BIAS.t30 60.7645
R17276 CS_BIAS.n130 CS_BIAS.t38 60.7645
R17277 CS_BIAS.n114 CS_BIAS.t32 60.7645
R17278 CS_BIAS.n148 CS_BIAS.t43 60.7645
R17279 CS_BIAS.n156 CS_BIAS.t33 60.7645
R17280 CS_BIAS.n58 CS_BIAS.t14 60.7645
R17281 CS_BIAS.n50 CS_BIAS.t10 60.7645
R17282 CS_BIAS.n16 CS_BIAS.t8 60.7645
R17283 CS_BIAS.n32 CS_BIAS.t2 60.7645
R17284 CS_BIAS.n21 CS_BIAS.t0 60.7645
R17285 CS_BIAS.n105 CS_BIAS.t42 60.7645
R17286 CS_BIAS.n97 CS_BIAS.t26 60.7645
R17287 CS_BIAS.n7 CS_BIAS.t40 60.7645
R17288 CS_BIAS.n79 CS_BIAS.t24 60.7645
R17289 CS_BIAS.n68 CS_BIAS.t37 60.7645
R17290 CS_BIAS.n277 CS_BIAS.t41 60.7645
R17291 CS_BIAS.n288 CS_BIAS.t34 60.7645
R17292 CS_BIAS.n295 CS_BIAS.t46 60.7645
R17293 CS_BIAS.n307 CS_BIAS.t45 60.7645
R17294 CS_BIAS.n315 CS_BIAS.t29 60.7645
R17295 CS_BIAS.n198 CS_BIAS.t22 60.7645
R17296 CS_BIAS.n209 CS_BIAS.t4 60.7645
R17297 CS_BIAS.n216 CS_BIAS.t6 60.7645
R17298 CS_BIAS.n228 CS_BIAS.t12 60.7645
R17299 CS_BIAS.n236 CS_BIAS.t16 60.7645
R17300 CS_BIAS.n264 CS_BIAS.t36 60.7645
R17301 CS_BIAS.n256 CS_BIAS.t27 60.7645
R17302 CS_BIAS.n244 CS_BIAS.t28 60.7645
R17303 CS_BIAS.n170 CS_BIAS.t25 60.7645
R17304 CS_BIAS.n181 CS_BIAS.t44 60.7645
R17305 CS_BIAS.n154 CS_BIAS.n108 60.4368
R17306 CS_BIAS.n56 CS_BIAS.n10 60.4368
R17307 CS_BIAS.n103 CS_BIAS.n1 60.4368
R17308 CS_BIAS.n313 CS_BIAS.n267 60.4368
R17309 CS_BIAS.n234 CS_BIAS.n188 60.4368
R17310 CS_BIAS.n262 CS_BIAS.n160 60.4368
R17311 CS_BIAS.n135 CS_BIAS.n115 56.5617
R17312 CS_BIAS.n136 CS_BIAS.n135 56.5617
R17313 CS_BIAS.n38 CS_BIAS.n37 56.5617
R17314 CS_BIAS.n37 CS_BIAS.n17 56.5617
R17315 CS_BIAS.n85 CS_BIAS.n84 56.5617
R17316 CS_BIAS.n84 CS_BIAS.n8 56.5617
R17317 CS_BIAS.n293 CS_BIAS.n273 56.5617
R17318 CS_BIAS.n294 CS_BIAS.n293 56.5617
R17319 CS_BIAS.n214 CS_BIAS.n194 56.5617
R17320 CS_BIAS.n215 CS_BIAS.n214 56.5617
R17321 CS_BIAS.n243 CS_BIAS.n242 56.5617
R17322 CS_BIAS.n242 CS_BIAS.n166 56.5617
R17323 CS_BIAS.n150 CS_BIAS.n108 52.6866
R17324 CS_BIAS.n52 CS_BIAS.n10 52.6866
R17325 CS_BIAS.n99 CS_BIAS.n1 52.6866
R17326 CS_BIAS.n309 CS_BIAS.n267 52.6866
R17327 CS_BIAS.n230 CS_BIAS.n188 52.6866
R17328 CS_BIAS.n258 CS_BIAS.n160 52.6866
R17329 CS_BIAS.n124 CS_BIAS.n123 34.28
R17330 CS_BIAS.n143 CS_BIAS.n110 34.28
R17331 CS_BIAS.n45 CS_BIAS.n12 34.28
R17332 CS_BIAS.n26 CS_BIAS.n25 34.28
R17333 CS_BIAS.n92 CS_BIAS.n3 34.28
R17334 CS_BIAS.n73 CS_BIAS.n72 34.28
R17335 CS_BIAS.n282 CS_BIAS.n281 34.28
R17336 CS_BIAS.n302 CS_BIAS.n269 34.28
R17337 CS_BIAS.n203 CS_BIAS.n202 34.28
R17338 CS_BIAS.n223 CS_BIAS.n190 34.28
R17339 CS_BIAS.n251 CS_BIAS.n162 34.28
R17340 CS_BIAS.n175 CS_BIAS.n174 34.28
R17341 CS_BIAS.n128 CS_BIAS.n117 30.405
R17342 CS_BIAS.n142 CS_BIAS.n141 30.405
R17343 CS_BIAS.n44 CS_BIAS.n43 30.405
R17344 CS_BIAS.n30 CS_BIAS.n19 30.405
R17345 CS_BIAS.n91 CS_BIAS.n90 30.405
R17346 CS_BIAS.n77 CS_BIAS.n66 30.405
R17347 CS_BIAS.n286 CS_BIAS.n275 30.405
R17348 CS_BIAS.n301 CS_BIAS.n300 30.405
R17349 CS_BIAS.n207 CS_BIAS.n196 30.405
R17350 CS_BIAS.n222 CS_BIAS.n221 30.405
R17351 CS_BIAS.n250 CS_BIAS.n249 30.405
R17352 CS_BIAS.n179 CS_BIAS.n168 30.405
R17353 CS_BIAS.n123 CS_BIAS.n122 24.5923
R17354 CS_BIAS.n131 CS_BIAS.n115 24.5923
R17355 CS_BIAS.n129 CS_BIAS.n128 24.5923
R17356 CS_BIAS.n141 CS_BIAS.n112 24.5923
R17357 CS_BIAS.n137 CS_BIAS.n136 24.5923
R17358 CS_BIAS.n150 CS_BIAS.n149 24.5923
R17359 CS_BIAS.n147 CS_BIAS.n110 24.5923
R17360 CS_BIAS.n155 CS_BIAS.n154 24.5923
R17361 CS_BIAS.n57 CS_BIAS.n56 24.5923
R17362 CS_BIAS.n52 CS_BIAS.n51 24.5923
R17363 CS_BIAS.n49 CS_BIAS.n12 24.5923
R17364 CS_BIAS.n43 CS_BIAS.n14 24.5923
R17365 CS_BIAS.n39 CS_BIAS.n38 24.5923
R17366 CS_BIAS.n33 CS_BIAS.n17 24.5923
R17367 CS_BIAS.n31 CS_BIAS.n30 24.5923
R17368 CS_BIAS.n25 CS_BIAS.n24 24.5923
R17369 CS_BIAS.n104 CS_BIAS.n103 24.5923
R17370 CS_BIAS.n99 CS_BIAS.n98 24.5923
R17371 CS_BIAS.n96 CS_BIAS.n3 24.5923
R17372 CS_BIAS.n90 CS_BIAS.n5 24.5923
R17373 CS_BIAS.n86 CS_BIAS.n85 24.5923
R17374 CS_BIAS.n80 CS_BIAS.n8 24.5923
R17375 CS_BIAS.n78 CS_BIAS.n77 24.5923
R17376 CS_BIAS.n72 CS_BIAS.n71 24.5923
R17377 CS_BIAS.n281 CS_BIAS.n280 24.5923
R17378 CS_BIAS.n287 CS_BIAS.n286 24.5923
R17379 CS_BIAS.n289 CS_BIAS.n273 24.5923
R17380 CS_BIAS.n296 CS_BIAS.n294 24.5923
R17381 CS_BIAS.n300 CS_BIAS.n271 24.5923
R17382 CS_BIAS.n306 CS_BIAS.n269 24.5923
R17383 CS_BIAS.n309 CS_BIAS.n308 24.5923
R17384 CS_BIAS.n314 CS_BIAS.n313 24.5923
R17385 CS_BIAS.n202 CS_BIAS.n201 24.5923
R17386 CS_BIAS.n208 CS_BIAS.n207 24.5923
R17387 CS_BIAS.n210 CS_BIAS.n194 24.5923
R17388 CS_BIAS.n217 CS_BIAS.n215 24.5923
R17389 CS_BIAS.n221 CS_BIAS.n192 24.5923
R17390 CS_BIAS.n227 CS_BIAS.n190 24.5923
R17391 CS_BIAS.n230 CS_BIAS.n229 24.5923
R17392 CS_BIAS.n235 CS_BIAS.n234 24.5923
R17393 CS_BIAS.n263 CS_BIAS.n262 24.5923
R17394 CS_BIAS.n255 CS_BIAS.n162 24.5923
R17395 CS_BIAS.n258 CS_BIAS.n257 24.5923
R17396 CS_BIAS.n245 CS_BIAS.n243 24.5923
R17397 CS_BIAS.n249 CS_BIAS.n164 24.5923
R17398 CS_BIAS.n174 CS_BIAS.n173 24.5923
R17399 CS_BIAS.n180 CS_BIAS.n179 24.5923
R17400 CS_BIAS.n182 CS_BIAS.n166 24.5923
R17401 CS_BIAS.n156 CS_BIAS.n155 20.9036
R17402 CS_BIAS.n58 CS_BIAS.n57 20.9036
R17403 CS_BIAS.n105 CS_BIAS.n104 20.9036
R17404 CS_BIAS.n315 CS_BIAS.n314 20.9036
R17405 CS_BIAS.n236 CS_BIAS.n235 20.9036
R17406 CS_BIAS.n264 CS_BIAS.n263 20.9036
R17407 CS_BIAS.n131 CS_BIAS.n130 18.9362
R17408 CS_BIAS.n137 CS_BIAS.n114 18.9362
R17409 CS_BIAS.n39 CS_BIAS.n16 18.9362
R17410 CS_BIAS.n33 CS_BIAS.n32 18.9362
R17411 CS_BIAS.n86 CS_BIAS.n7 18.9362
R17412 CS_BIAS.n80 CS_BIAS.n79 18.9362
R17413 CS_BIAS.n289 CS_BIAS.n288 18.9362
R17414 CS_BIAS.n296 CS_BIAS.n295 18.9362
R17415 CS_BIAS.n210 CS_BIAS.n209 18.9362
R17416 CS_BIAS.n217 CS_BIAS.n216 18.9362
R17417 CS_BIAS.n245 CS_BIAS.n244 18.9362
R17418 CS_BIAS.n182 CS_BIAS.n181 18.9362
R17419 CS_BIAS.n149 CS_BIAS.n148 16.9689
R17420 CS_BIAS.n51 CS_BIAS.n50 16.9689
R17421 CS_BIAS.n98 CS_BIAS.n97 16.9689
R17422 CS_BIAS.n308 CS_BIAS.n307 16.9689
R17423 CS_BIAS.n229 CS_BIAS.n228 16.9689
R17424 CS_BIAS.n257 CS_BIAS.n256 16.9689
R17425 CS_BIAS.n61 CS_BIAS.n59 12.7074
R17426 CS_BIAS.n239 CS_BIAS.n237 12.7074
R17427 CS_BIAS.n318 CS_BIAS.n158 12.4945
R17428 CS_BIAS.n318 CS_BIAS.n317 10.4597
R17429 CS_BIAS.n83 CS_BIAS.n64 9.50363
R17430 CS_BIAS.n241 CS_BIAS.n240 9.50363
R17431 CS_BIAS.n158 CS_BIAS.n106 8.34667
R17432 CS_BIAS.n317 CS_BIAS.n265 8.34667
R17433 CS_BIAS.n122 CS_BIAS.n119 7.62397
R17434 CS_BIAS.n148 CS_BIAS.n147 7.62397
R17435 CS_BIAS.n50 CS_BIAS.n49 7.62397
R17436 CS_BIAS.n24 CS_BIAS.n21 7.62397
R17437 CS_BIAS.n97 CS_BIAS.n96 7.62397
R17438 CS_BIAS.n71 CS_BIAS.n68 7.62397
R17439 CS_BIAS.n280 CS_BIAS.n277 7.62397
R17440 CS_BIAS.n307 CS_BIAS.n306 7.62397
R17441 CS_BIAS.n201 CS_BIAS.n198 7.62397
R17442 CS_BIAS.n228 CS_BIAS.n227 7.62397
R17443 CS_BIAS.n256 CS_BIAS.n255 7.62397
R17444 CS_BIAS.n173 CS_BIAS.n170 7.62397
R17445 CS_BIAS.n121 CS_BIAS.n120 7.55607
R17446 CS_BIAS.n23 CS_BIAS.n22 7.55607
R17447 CS_BIAS.n70 CS_BIAS.n69 7.55607
R17448 CS_BIAS.n279 CS_BIAS.n278 7.55607
R17449 CS_BIAS.n200 CS_BIAS.n199 7.55607
R17450 CS_BIAS.n172 CS_BIAS.n171 7.55607
R17451 CS_BIAS.n63 CS_BIAS.t1 7.44411
R17452 CS_BIAS.n63 CS_BIAS.t19 7.44411
R17453 CS_BIAS.n62 CS_BIAS.t9 7.44411
R17454 CS_BIAS.n62 CS_BIAS.t3 7.44411
R17455 CS_BIAS.n60 CS_BIAS.t15 7.44411
R17456 CS_BIAS.n60 CS_BIAS.t11 7.44411
R17457 CS_BIAS.n238 CS_BIAS.t13 7.44411
R17458 CS_BIAS.n238 CS_BIAS.t17 7.44411
R17459 CS_BIAS.n186 CS_BIAS.t5 7.44411
R17460 CS_BIAS.n186 CS_BIAS.t7 7.44411
R17461 CS_BIAS.n185 CS_BIAS.t21 7.44411
R17462 CS_BIAS.n185 CS_BIAS.t23 7.44411
R17463 CS_BIAS.n130 CS_BIAS.n129 5.65662
R17464 CS_BIAS.n114 CS_BIAS.n112 5.65662
R17465 CS_BIAS.n16 CS_BIAS.n14 5.65662
R17466 CS_BIAS.n32 CS_BIAS.n31 5.65662
R17467 CS_BIAS.n7 CS_BIAS.n5 5.65662
R17468 CS_BIAS.n79 CS_BIAS.n78 5.65662
R17469 CS_BIAS.n288 CS_BIAS.n287 5.65662
R17470 CS_BIAS.n295 CS_BIAS.n271 5.65662
R17471 CS_BIAS.n209 CS_BIAS.n208 5.65662
R17472 CS_BIAS.n216 CS_BIAS.n192 5.65662
R17473 CS_BIAS.n244 CS_BIAS.n164 5.65662
R17474 CS_BIAS.n181 CS_BIAS.n180 5.65662
R17475 CS_BIAS.n158 CS_BIAS.n157 5.07394
R17476 CS_BIAS.n317 CS_BIAS.n316 5.07394
R17477 CS_BIAS CS_BIAS.n318 4.5855
R17478 CS_BIAS.n64 CS_BIAS.n61 0.796477
R17479 CS_BIAS.n240 CS_BIAS.n239 0.796477
R17480 CS_BIAS.n157 CS_BIAS.n107 0.278335
R17481 CS_BIAS.n59 CS_BIAS.n9 0.278335
R17482 CS_BIAS.n106 CS_BIAS.n0 0.278335
R17483 CS_BIAS.n316 CS_BIAS.n266 0.278335
R17484 CS_BIAS.n237 CS_BIAS.n187 0.278335
R17485 CS_BIAS.n265 CS_BIAS.n159 0.278335
R17486 CS_BIAS.n153 CS_BIAS.n107 0.189894
R17487 CS_BIAS.n153 CS_BIAS.n152 0.189894
R17488 CS_BIAS.n152 CS_BIAS.n151 0.189894
R17489 CS_BIAS.n151 CS_BIAS.n109 0.189894
R17490 CS_BIAS.n146 CS_BIAS.n109 0.189894
R17491 CS_BIAS.n146 CS_BIAS.n145 0.189894
R17492 CS_BIAS.n145 CS_BIAS.n144 0.189894
R17493 CS_BIAS.n144 CS_BIAS.n111 0.189894
R17494 CS_BIAS.n140 CS_BIAS.n111 0.189894
R17495 CS_BIAS.n140 CS_BIAS.n139 0.189894
R17496 CS_BIAS.n139 CS_BIAS.n138 0.189894
R17497 CS_BIAS.n138 CS_BIAS.n113 0.189894
R17498 CS_BIAS.n134 CS_BIAS.n113 0.189894
R17499 CS_BIAS.n134 CS_BIAS.n133 0.189894
R17500 CS_BIAS.n133 CS_BIAS.n132 0.189894
R17501 CS_BIAS.n132 CS_BIAS.n116 0.189894
R17502 CS_BIAS.n127 CS_BIAS.n116 0.189894
R17503 CS_BIAS.n127 CS_BIAS.n126 0.189894
R17504 CS_BIAS.n126 CS_BIAS.n125 0.189894
R17505 CS_BIAS.n125 CS_BIAS.n118 0.189894
R17506 CS_BIAS.n121 CS_BIAS.n118 0.189894
R17507 CS_BIAS.n55 CS_BIAS.n9 0.189894
R17508 CS_BIAS.n55 CS_BIAS.n54 0.189894
R17509 CS_BIAS.n54 CS_BIAS.n53 0.189894
R17510 CS_BIAS.n53 CS_BIAS.n11 0.189894
R17511 CS_BIAS.n48 CS_BIAS.n11 0.189894
R17512 CS_BIAS.n48 CS_BIAS.n47 0.189894
R17513 CS_BIAS.n47 CS_BIAS.n46 0.189894
R17514 CS_BIAS.n46 CS_BIAS.n13 0.189894
R17515 CS_BIAS.n42 CS_BIAS.n13 0.189894
R17516 CS_BIAS.n42 CS_BIAS.n41 0.189894
R17517 CS_BIAS.n41 CS_BIAS.n40 0.189894
R17518 CS_BIAS.n40 CS_BIAS.n15 0.189894
R17519 CS_BIAS.n36 CS_BIAS.n15 0.189894
R17520 CS_BIAS.n36 CS_BIAS.n35 0.189894
R17521 CS_BIAS.n35 CS_BIAS.n34 0.189894
R17522 CS_BIAS.n34 CS_BIAS.n18 0.189894
R17523 CS_BIAS.n29 CS_BIAS.n18 0.189894
R17524 CS_BIAS.n29 CS_BIAS.n28 0.189894
R17525 CS_BIAS.n28 CS_BIAS.n27 0.189894
R17526 CS_BIAS.n27 CS_BIAS.n20 0.189894
R17527 CS_BIAS.n23 CS_BIAS.n20 0.189894
R17528 CS_BIAS.n82 CS_BIAS.n81 0.189894
R17529 CS_BIAS.n81 CS_BIAS.n65 0.189894
R17530 CS_BIAS.n76 CS_BIAS.n65 0.189894
R17531 CS_BIAS.n76 CS_BIAS.n75 0.189894
R17532 CS_BIAS.n75 CS_BIAS.n74 0.189894
R17533 CS_BIAS.n74 CS_BIAS.n67 0.189894
R17534 CS_BIAS.n70 CS_BIAS.n67 0.189894
R17535 CS_BIAS.n102 CS_BIAS.n0 0.189894
R17536 CS_BIAS.n102 CS_BIAS.n101 0.189894
R17537 CS_BIAS.n101 CS_BIAS.n100 0.189894
R17538 CS_BIAS.n100 CS_BIAS.n2 0.189894
R17539 CS_BIAS.n95 CS_BIAS.n2 0.189894
R17540 CS_BIAS.n95 CS_BIAS.n94 0.189894
R17541 CS_BIAS.n94 CS_BIAS.n93 0.189894
R17542 CS_BIAS.n93 CS_BIAS.n4 0.189894
R17543 CS_BIAS.n89 CS_BIAS.n4 0.189894
R17544 CS_BIAS.n89 CS_BIAS.n88 0.189894
R17545 CS_BIAS.n88 CS_BIAS.n87 0.189894
R17546 CS_BIAS.n87 CS_BIAS.n6 0.189894
R17547 CS_BIAS.n279 CS_BIAS.n276 0.189894
R17548 CS_BIAS.n283 CS_BIAS.n276 0.189894
R17549 CS_BIAS.n284 CS_BIAS.n283 0.189894
R17550 CS_BIAS.n285 CS_BIAS.n284 0.189894
R17551 CS_BIAS.n285 CS_BIAS.n274 0.189894
R17552 CS_BIAS.n290 CS_BIAS.n274 0.189894
R17553 CS_BIAS.n291 CS_BIAS.n290 0.189894
R17554 CS_BIAS.n292 CS_BIAS.n291 0.189894
R17555 CS_BIAS.n292 CS_BIAS.n272 0.189894
R17556 CS_BIAS.n297 CS_BIAS.n272 0.189894
R17557 CS_BIAS.n298 CS_BIAS.n297 0.189894
R17558 CS_BIAS.n299 CS_BIAS.n298 0.189894
R17559 CS_BIAS.n299 CS_BIAS.n270 0.189894
R17560 CS_BIAS.n303 CS_BIAS.n270 0.189894
R17561 CS_BIAS.n304 CS_BIAS.n303 0.189894
R17562 CS_BIAS.n305 CS_BIAS.n304 0.189894
R17563 CS_BIAS.n305 CS_BIAS.n268 0.189894
R17564 CS_BIAS.n310 CS_BIAS.n268 0.189894
R17565 CS_BIAS.n311 CS_BIAS.n310 0.189894
R17566 CS_BIAS.n312 CS_BIAS.n311 0.189894
R17567 CS_BIAS.n312 CS_BIAS.n266 0.189894
R17568 CS_BIAS.n200 CS_BIAS.n197 0.189894
R17569 CS_BIAS.n204 CS_BIAS.n197 0.189894
R17570 CS_BIAS.n205 CS_BIAS.n204 0.189894
R17571 CS_BIAS.n206 CS_BIAS.n205 0.189894
R17572 CS_BIAS.n206 CS_BIAS.n195 0.189894
R17573 CS_BIAS.n211 CS_BIAS.n195 0.189894
R17574 CS_BIAS.n212 CS_BIAS.n211 0.189894
R17575 CS_BIAS.n213 CS_BIAS.n212 0.189894
R17576 CS_BIAS.n213 CS_BIAS.n193 0.189894
R17577 CS_BIAS.n218 CS_BIAS.n193 0.189894
R17578 CS_BIAS.n219 CS_BIAS.n218 0.189894
R17579 CS_BIAS.n220 CS_BIAS.n219 0.189894
R17580 CS_BIAS.n220 CS_BIAS.n191 0.189894
R17581 CS_BIAS.n224 CS_BIAS.n191 0.189894
R17582 CS_BIAS.n225 CS_BIAS.n224 0.189894
R17583 CS_BIAS.n226 CS_BIAS.n225 0.189894
R17584 CS_BIAS.n226 CS_BIAS.n189 0.189894
R17585 CS_BIAS.n231 CS_BIAS.n189 0.189894
R17586 CS_BIAS.n232 CS_BIAS.n231 0.189894
R17587 CS_BIAS.n233 CS_BIAS.n232 0.189894
R17588 CS_BIAS.n233 CS_BIAS.n187 0.189894
R17589 CS_BIAS.n172 CS_BIAS.n169 0.189894
R17590 CS_BIAS.n176 CS_BIAS.n169 0.189894
R17591 CS_BIAS.n177 CS_BIAS.n176 0.189894
R17592 CS_BIAS.n178 CS_BIAS.n177 0.189894
R17593 CS_BIAS.n178 CS_BIAS.n167 0.189894
R17594 CS_BIAS.n183 CS_BIAS.n167 0.189894
R17595 CS_BIAS.n184 CS_BIAS.n183 0.189894
R17596 CS_BIAS.n246 CS_BIAS.n165 0.189894
R17597 CS_BIAS.n247 CS_BIAS.n246 0.189894
R17598 CS_BIAS.n248 CS_BIAS.n247 0.189894
R17599 CS_BIAS.n248 CS_BIAS.n163 0.189894
R17600 CS_BIAS.n252 CS_BIAS.n163 0.189894
R17601 CS_BIAS.n253 CS_BIAS.n252 0.189894
R17602 CS_BIAS.n254 CS_BIAS.n253 0.189894
R17603 CS_BIAS.n254 CS_BIAS.n161 0.189894
R17604 CS_BIAS.n259 CS_BIAS.n161 0.189894
R17605 CS_BIAS.n260 CS_BIAS.n259 0.189894
R17606 CS_BIAS.n261 CS_BIAS.n260 0.189894
R17607 CS_BIAS.n261 CS_BIAS.n159 0.189894
R17608 CS_BIAS.n83 CS_BIAS.n82 0.170955
R17609 CS_BIAS.n83 CS_BIAS.n6 0.170955
R17610 CS_BIAS.n241 CS_BIAS.n184 0.170955
R17611 CS_BIAS.n241 CS_BIAS.n165 0.170955
R17612 a_n12950_8244.n14 a_n12950_8244.t1 226.136
R17613 a_n12950_8244.n14 a_n12950_8244.t0 219.459
R17614 a_n12950_8244.t2 a_n12950_8244.n15 101.132
R17615 a_n12950_8244.n15 a_n12950_8244.t3 68.8751
R17616 a_n12950_8244.n3 a_n12950_8244.n13 1.26083
R17617 a_n12950_8244.n9 a_n12950_8244.n10 1.26083
R17618 a_n12950_8244.n2 a_n12950_8244.n8 1.26083
R17619 a_n12950_8244.n4 a_n12950_8244.n5 1.26083
R17620 a_n12950_8244.n9 a_n12950_8244.t12 55.8643
R17621 a_n12950_8244.n2 a_n12950_8244.t18 55.8643
R17622 a_n12950_8244.n0 a_n12950_8244.t21 55.8643
R17623 a_n12950_8244.n0 a_n12950_8244.t19 55.8643
R17624 a_n12950_8244.n4 a_n12950_8244.t8 55.8643
R17625 a_n12950_8244.n3 a_n12950_8244.t23 55.8638
R17626 a_n12950_8244.n1 a_n12950_8244.t27 55.8638
R17627 a_n12950_8244.n1 a_n12950_8244.t26 55.8638
R17628 a_n12950_8244.n13 a_n12950_8244.t20 55.5833
R17629 a_n12950_8244.n13 a_n12950_8244.t6 54.7713
R17630 a_n12950_8244.n12 a_n12950_8244.t25 55.5833
R17631 a_n12950_8244.n12 a_n12950_8244.t10 54.7713
R17632 a_n12950_8244.n11 a_n12950_8244.t24 55.5833
R17633 a_n12950_8244.n11 a_n12950_8244.t9 54.7713
R17634 a_n12950_8244.n10 a_n12950_8244.t11 55.5833
R17635 a_n12950_8244.n10 a_n12950_8244.t17 54.7713
R17636 a_n12950_8244.n8 a_n12950_8244.t4 55.5833
R17637 a_n12950_8244.n8 a_n12950_8244.t13 54.7713
R17638 a_n12950_8244.n7 a_n12950_8244.t7 55.5833
R17639 a_n12950_8244.n7 a_n12950_8244.t15 54.7713
R17640 a_n12950_8244.n6 a_n12950_8244.t5 55.5833
R17641 a_n12950_8244.n6 a_n12950_8244.t14 54.7713
R17642 a_n12950_8244.n5 a_n12950_8244.t16 55.5833
R17643 a_n12950_8244.n5 a_n12950_8244.t22 54.7713
R17644 a_n12950_8244.n0 a_n12950_8244.n6 12.8147
R17645 a_n12950_8244.n15 a_n12950_8244.n0 12.3441
R17646 a_n12950_8244.n0 a_n12950_8244.n14 11.6448
R17647 a_n12950_8244.n1 a_n12950_8244.n3 10.5288
R17648 a_n12950_8244.n0 a_n12950_8244.n2 10.5288
R17649 a_n12950_8244.n0 a_n12950_8244.n1 9.46297
R17650 a_n12950_8244.n1 a_n12950_8244.n9 7.90755
R17651 a_n12950_8244.n0 a_n12950_8244.n4 7.90755
R17652 a_n12950_8244.n0 a_n12950_8244.n7 6.54667
R17653 a_n12950_8244.n1 a_n12950_8244.n11 6.54667
R17654 a_n12950_8244.n1 a_n12950_8244.n12 6.54667
R17655 a_n7062_10679.n3 a_n7062_10679.t0 211.798
R17656 a_n7062_10679.n3 a_n7062_10679.t1 210.631
R17657 a_n7062_10679.n1 a_n7062_10679.t5 179.327
R17658 a_n7062_10679.n0 a_n7062_10679.t4 178.219
R17659 a_n7062_10679.n1 a_n7062_10679.t7 178.219
R17660 a_n7062_10679.t8 a_n7062_10679.n1 178.219
R17661 a_n7062_10679.n0 a_n7062_10679.n4 148.534
R17662 a_n7062_10679.n1 a_n7062_10679.n2 148.534
R17663 a_n7062_10679.n4 a_n7062_10679.t9 29.6854
R17664 a_n7062_10679.n4 a_n7062_10679.t6 29.6854
R17665 a_n7062_10679.n2 a_n7062_10679.t2 29.6854
R17666 a_n7062_10679.n2 a_n7062_10679.t3 29.6854
R17667 a_n7062_10679.n0 a_n7062_10679.n3 5.46243
R17668 a_n7062_10679.n1 a_n7062_10679.n0 3.58814
R17669 VN.n1 VN.t1 243.97
R17670 VN.n1 VN.t0 243.255
R17671 VN.n0 VN.t3 101.347
R17672 VN.n0 VN.t2 81.4176
R17673 VN VN.n2 15.8418
R17674 VN.n2 VN.n1 5.04791
R17675 VN.n2 VN.n0 1.188
R17676 VP.n1 VP.t0 243.97
R17677 VP.n1 VP.t1 243.255
R17678 VP.n0 VP.t3 101.561
R17679 VP.n0 VP.t2 81.635
R17680 VP VP.n2 12.9059
R17681 VP.n2 VP.n1 4.80222
R17682 VP.n2 VP.n0 0.972091
C0 VOUT VN 0.943236f
C1 VOUT CS_BIAS 19.8501f
C2 VP VN 10.6834f
C3 VP CS_BIAS 0.333256f
C4 VN CS_BIAS 0.269434f
C5 a_7190_10679# VDD 1.32893f
C6 VDD VOUT 45.726997f
C7 VOUT VP 3.88895f
C8 VDD VN 0.193966f
C9 a_n8118_10679# VDD 1.32866f
C10 DIFFPAIR_BIAS GND 44.060894f
C11 CS_BIAS GND 97.797485f
C12 VN GND 29.146532f
C13 VP GND 24.7845f
C14 VOUT GND 66.31035f
C15 VDD GND 0.55077p
C16 a_7190_10679# GND 0.421214f
C17 a_n8118_10679# GND 0.421567f
C18 VP.t2 GND 2.16234f
C19 VP.t3 GND 2.44675f
C20 VP.n0 GND 2.67477f
C21 VP.t0 GND 0.032188f
C22 VP.t1 GND 0.031992f
C23 VP.n1 GND 0.15332f
C24 VP.n2 GND 1.81964f
C25 VN.t2 GND 1.59103f
C26 VN.t3 GND 1.79958f
C27 VN.n0 GND 1.96168f
C28 VN.t1 GND 0.023716f
C29 VN.t0 GND 0.023572f
C30 VN.n1 GND 0.120419f
C31 VN.n2 GND 2.18337f
C32 a_n7062_10679.n0 GND 3.76636f
C33 a_n7062_10679.n1 GND 5.19801f
C34 a_n7062_10679.t5 GND 0.341455f
C35 a_n7062_10679.t2 GND 0.068347f
C36 a_n7062_10679.t3 GND 0.068347f
C37 a_n7062_10679.n2 GND 0.226333f
C38 a_n7062_10679.t1 GND 0.700148f
C39 a_n7062_10679.t0 GND 0.921247f
C40 a_n7062_10679.n3 GND 16.5428f
C41 a_n7062_10679.t4 GND 0.334656f
C42 a_n7062_10679.t9 GND 0.068347f
C43 a_n7062_10679.t6 GND 0.068347f
C44 a_n7062_10679.n4 GND 0.226333f
C45 a_n7062_10679.t7 GND 0.334656f
C46 a_n7062_10679.t8 GND 0.334655f
C47 a_n12950_8244.n0 GND 24.829401f
C48 a_n12950_8244.n1 GND 5.27819f
C49 a_n12950_8244.n2 GND 1.50914f
C50 a_n12950_8244.n3 GND 1.50914f
C51 a_n12950_8244.n4 GND 1.5643f
C52 a_n12950_8244.n5 GND 0.774824f
C53 a_n12950_8244.n6 GND 0.774824f
C54 a_n12950_8244.n7 GND 0.774824f
C55 a_n12950_8244.n8 GND 0.774824f
C56 a_n12950_8244.n9 GND 1.5643f
C57 a_n12950_8244.n10 GND 0.774824f
C58 a_n12950_8244.n11 GND 0.774824f
C59 a_n12950_8244.n12 GND 0.774824f
C60 a_n12950_8244.n13 GND 0.774824f
C61 a_n12950_8244.t1 GND 0.845892f
C62 a_n12950_8244.t0 GND 0.664151f
C63 a_n12950_8244.n14 GND 17.3234f
C64 a_n12950_8244.t22 GND 1.53361f
C65 a_n12950_8244.t8 GND 1.547f
C66 a_n12950_8244.t16 GND 1.53855f
C67 a_n12950_8244.t14 GND 1.53361f
C68 a_n12950_8244.t19 GND 1.547f
C69 a_n12950_8244.t5 GND 1.53855f
C70 a_n12950_8244.t15 GND 1.53361f
C71 a_n12950_8244.t21 GND 1.547f
C72 a_n12950_8244.t7 GND 1.53855f
C73 a_n12950_8244.t13 GND 1.53361f
C74 a_n12950_8244.t18 GND 1.547f
C75 a_n12950_8244.t4 GND 1.53855f
C76 a_n12950_8244.t17 GND 1.53361f
C77 a_n12950_8244.t12 GND 1.547f
C78 a_n12950_8244.t11 GND 1.53855f
C79 a_n12950_8244.t9 GND 1.53361f
C80 a_n12950_8244.t26 GND 1.54699f
C81 a_n12950_8244.t24 GND 1.53855f
C82 a_n12950_8244.t10 GND 1.53361f
C83 a_n12950_8244.t27 GND 1.54699f
C84 a_n12950_8244.t25 GND 1.53855f
C85 a_n12950_8244.t6 GND 1.53361f
C86 a_n12950_8244.t23 GND 1.54699f
C87 a_n12950_8244.t20 GND 1.53855f
C88 a_n12950_8244.t3 GND 1.19023f
C89 a_n12950_8244.n15 GND 5.13776f
C90 a_n12950_8244.t2 GND 2.03226f
C91 CS_BIAS.n0 GND 0.007421f
C92 CS_BIAS.t42 GND 0.165978f
C93 CS_BIAS.n1 GND 0.003322f
C94 CS_BIAS.n2 GND 0.005629f
C95 CS_BIAS.t26 GND 0.165978f
C96 CS_BIAS.n3 GND 0.011312f
C97 CS_BIAS.n4 GND 0.005629f
C98 CS_BIAS.n5 GND 0.00647f
C99 CS_BIAS.n6 GND 0.005602f
C100 CS_BIAS.t40 GND 0.165978f
C101 CS_BIAS.n7 GND 0.064177f
C102 CS_BIAS.n8 GND 0.009506f
C103 CS_BIAS.n9 GND 0.007421f
C104 CS_BIAS.t14 GND 0.165978f
C105 CS_BIAS.n10 GND 0.003322f
C106 CS_BIAS.n11 GND 0.005629f
C107 CS_BIAS.t10 GND 0.165978f
C108 CS_BIAS.n12 GND 0.011312f
C109 CS_BIAS.n13 GND 0.005629f
C110 CS_BIAS.n14 GND 0.00647f
C111 CS_BIAS.n15 GND 0.005629f
C112 CS_BIAS.t8 GND 0.165978f
C113 CS_BIAS.n16 GND 0.064177f
C114 CS_BIAS.n17 GND 0.009506f
C115 CS_BIAS.n18 GND 0.005629f
C116 CS_BIAS.t2 GND 0.165978f
C117 CS_BIAS.n19 GND 0.005451f
C118 CS_BIAS.n20 GND 0.005629f
C119 CS_BIAS.t0 GND 0.165978f
C120 CS_BIAS.n21 GND 0.077843f
C121 CS_BIAS.t18 GND 0.201331f
C122 CS_BIAS.n22 GND 0.076644f
C123 CS_BIAS.n23 GND 0.047175f
C124 CS_BIAS.n24 GND 0.006883f
C125 CS_BIAS.n25 GND 0.011312f
C126 CS_BIAS.n26 GND 0.004779f
C127 CS_BIAS.n27 GND 0.005629f
C128 CS_BIAS.n28 GND 0.005629f
C129 CS_BIAS.n29 GND 0.005629f
C130 CS_BIAS.n30 GND 0.011187f
C131 CS_BIAS.n31 GND 0.00647f
C132 CS_BIAS.n32 GND 0.064177f
C133 CS_BIAS.n33 GND 0.009253f
C134 CS_BIAS.n34 GND 0.005629f
C135 CS_BIAS.n35 GND 0.005629f
C136 CS_BIAS.n36 GND 0.005629f
C137 CS_BIAS.n37 GND 0.003279f
C138 CS_BIAS.n38 GND 0.009506f
C139 CS_BIAS.n39 GND 0.009253f
C140 CS_BIAS.n40 GND 0.005629f
C141 CS_BIAS.n41 GND 0.005629f
C142 CS_BIAS.n42 GND 0.005629f
C143 CS_BIAS.n43 GND 0.011187f
C144 CS_BIAS.n44 GND 0.005451f
C145 CS_BIAS.n45 GND 0.004779f
C146 CS_BIAS.n46 GND 0.005629f
C147 CS_BIAS.n47 GND 0.005629f
C148 CS_BIAS.n48 GND 0.005629f
C149 CS_BIAS.n49 GND 0.006883f
C150 CS_BIAS.n50 GND 0.064177f
C151 CS_BIAS.n51 GND 0.008841f
C152 CS_BIAS.n52 GND 0.009998f
C153 CS_BIAS.n53 GND 0.005629f
C154 CS_BIAS.n54 GND 0.005629f
C155 CS_BIAS.n55 GND 0.005629f
C156 CS_BIAS.n56 GND 0.008971f
C157 CS_BIAS.n57 GND 0.009665f
C158 CS_BIAS.n58 GND 0.082618f
C159 CS_BIAS.n59 GND 0.064948f
C160 CS_BIAS.t15 GND 0.018462f
C161 CS_BIAS.t11 GND 0.018462f
C162 CS_BIAS.n60 GND 0.1295f
C163 CS_BIAS.n61 GND 0.181834f
C164 CS_BIAS.t9 GND 0.018462f
C165 CS_BIAS.t3 GND 0.018462f
C166 CS_BIAS.n62 GND 0.1295f
C167 CS_BIAS.t1 GND 0.018462f
C168 CS_BIAS.t19 GND 0.018462f
C169 CS_BIAS.n63 GND 0.13121f
C170 CS_BIAS.n64 GND 0.311293f
C171 CS_BIAS.n65 GND 0.005629f
C172 CS_BIAS.t24 GND 0.165978f
C173 CS_BIAS.n66 GND 0.005451f
C174 CS_BIAS.n67 GND 0.005629f
C175 CS_BIAS.t37 GND 0.165978f
C176 CS_BIAS.n68 GND 0.077843f
C177 CS_BIAS.t47 GND 0.201331f
C178 CS_BIAS.n69 GND 0.076644f
C179 CS_BIAS.n70 GND 0.047175f
C180 CS_BIAS.n71 GND 0.006883f
C181 CS_BIAS.n72 GND 0.011312f
C182 CS_BIAS.n73 GND 0.004779f
C183 CS_BIAS.n74 GND 0.005629f
C184 CS_BIAS.n75 GND 0.005629f
C185 CS_BIAS.n76 GND 0.005629f
C186 CS_BIAS.n77 GND 0.011187f
C187 CS_BIAS.n78 GND 0.00647f
C188 CS_BIAS.n79 GND 0.064177f
C189 CS_BIAS.n80 GND 0.009253f
C190 CS_BIAS.n81 GND 0.005629f
C191 CS_BIAS.n82 GND 0.005602f
C192 CS_BIAS.n83 GND 0.04069f
C193 CS_BIAS.n84 GND 0.003279f
C194 CS_BIAS.n85 GND 0.009506f
C195 CS_BIAS.n86 GND 0.009253f
C196 CS_BIAS.n87 GND 0.005629f
C197 CS_BIAS.n88 GND 0.005629f
C198 CS_BIAS.n89 GND 0.005629f
C199 CS_BIAS.n90 GND 0.011187f
C200 CS_BIAS.n91 GND 0.005451f
C201 CS_BIAS.n92 GND 0.004779f
C202 CS_BIAS.n93 GND 0.005629f
C203 CS_BIAS.n94 GND 0.005629f
C204 CS_BIAS.n95 GND 0.005629f
C205 CS_BIAS.n96 GND 0.006883f
C206 CS_BIAS.n97 GND 0.064177f
C207 CS_BIAS.n98 GND 0.008841f
C208 CS_BIAS.n99 GND 0.009998f
C209 CS_BIAS.n100 GND 0.005629f
C210 CS_BIAS.n101 GND 0.005629f
C211 CS_BIAS.n102 GND 0.005629f
C212 CS_BIAS.n103 GND 0.008971f
C213 CS_BIAS.n104 GND 0.009665f
C214 CS_BIAS.n105 GND 0.082618f
C215 CS_BIAS.n106 GND 0.034138f
C216 CS_BIAS.n107 GND 0.007421f
C217 CS_BIAS.t33 GND 0.165978f
C218 CS_BIAS.n108 GND 0.003322f
C219 CS_BIAS.n109 GND 0.005629f
C220 CS_BIAS.t43 GND 0.165978f
C221 CS_BIAS.n110 GND 0.011312f
C222 CS_BIAS.n111 GND 0.005629f
C223 CS_BIAS.n112 GND 0.00647f
C224 CS_BIAS.n113 GND 0.005629f
C225 CS_BIAS.t32 GND 0.165978f
C226 CS_BIAS.n114 GND 0.064177f
C227 CS_BIAS.n115 GND 0.009506f
C228 CS_BIAS.n116 GND 0.005629f
C229 CS_BIAS.t38 GND 0.165978f
C230 CS_BIAS.n117 GND 0.005451f
C231 CS_BIAS.n118 GND 0.005629f
C232 CS_BIAS.t30 GND 0.165978f
C233 CS_BIAS.n119 GND 0.077843f
C234 CS_BIAS.t35 GND 0.201331f
C235 CS_BIAS.n120 GND 0.076644f
C236 CS_BIAS.n121 GND 0.047175f
C237 CS_BIAS.n122 GND 0.006883f
C238 CS_BIAS.n123 GND 0.011312f
C239 CS_BIAS.n124 GND 0.004779f
C240 CS_BIAS.n125 GND 0.005629f
C241 CS_BIAS.n126 GND 0.005629f
C242 CS_BIAS.n127 GND 0.005629f
C243 CS_BIAS.n128 GND 0.011187f
C244 CS_BIAS.n129 GND 0.00647f
C245 CS_BIAS.n130 GND 0.064177f
C246 CS_BIAS.n131 GND 0.009253f
C247 CS_BIAS.n132 GND 0.005629f
C248 CS_BIAS.n133 GND 0.005629f
C249 CS_BIAS.n134 GND 0.005629f
C250 CS_BIAS.n135 GND 0.003279f
C251 CS_BIAS.n136 GND 0.009506f
C252 CS_BIAS.n137 GND 0.009253f
C253 CS_BIAS.n138 GND 0.005629f
C254 CS_BIAS.n139 GND 0.005629f
C255 CS_BIAS.n140 GND 0.005629f
C256 CS_BIAS.n141 GND 0.011187f
C257 CS_BIAS.n142 GND 0.005451f
C258 CS_BIAS.n143 GND 0.004779f
C259 CS_BIAS.n144 GND 0.005629f
C260 CS_BIAS.n145 GND 0.005629f
C261 CS_BIAS.n146 GND 0.005629f
C262 CS_BIAS.n147 GND 0.006883f
C263 CS_BIAS.n148 GND 0.064177f
C264 CS_BIAS.n149 GND 0.008841f
C265 CS_BIAS.n150 GND 0.009998f
C266 CS_BIAS.n151 GND 0.005629f
C267 CS_BIAS.n152 GND 0.005629f
C268 CS_BIAS.n153 GND 0.005629f
C269 CS_BIAS.n154 GND 0.008971f
C270 CS_BIAS.n155 GND 0.009665f
C271 CS_BIAS.n156 GND 0.082618f
C272 CS_BIAS.n157 GND 0.020913f
C273 CS_BIAS.n158 GND 0.336679f
C274 CS_BIAS.n159 GND 0.007421f
C275 CS_BIAS.t36 GND 0.165978f
C276 CS_BIAS.n160 GND 0.003322f
C277 CS_BIAS.n161 GND 0.005629f
C278 CS_BIAS.t27 GND 0.165978f
C279 CS_BIAS.n162 GND 0.011312f
C280 CS_BIAS.n163 GND 0.005629f
C281 CS_BIAS.n164 GND 0.00647f
C282 CS_BIAS.n165 GND 0.005602f
C283 CS_BIAS.n166 GND 0.009506f
C284 CS_BIAS.n167 GND 0.005629f
C285 CS_BIAS.t44 GND 0.165978f
C286 CS_BIAS.n168 GND 0.005451f
C287 CS_BIAS.n169 GND 0.005629f
C288 CS_BIAS.t25 GND 0.165978f
C289 CS_BIAS.n170 GND 0.077843f
C290 CS_BIAS.t39 GND 0.201331f
C291 CS_BIAS.n171 GND 0.076644f
C292 CS_BIAS.n172 GND 0.047175f
C293 CS_BIAS.n173 GND 0.006883f
C294 CS_BIAS.n174 GND 0.011312f
C295 CS_BIAS.n175 GND 0.004779f
C296 CS_BIAS.n176 GND 0.005629f
C297 CS_BIAS.n177 GND 0.005629f
C298 CS_BIAS.n178 GND 0.005629f
C299 CS_BIAS.n179 GND 0.011187f
C300 CS_BIAS.n180 GND 0.00647f
C301 CS_BIAS.n181 GND 0.064177f
C302 CS_BIAS.n182 GND 0.009253f
C303 CS_BIAS.n183 GND 0.005629f
C304 CS_BIAS.n184 GND 0.005602f
C305 CS_BIAS.t21 GND 0.018462f
C306 CS_BIAS.t23 GND 0.018462f
C307 CS_BIAS.n185 GND 0.13121f
C308 CS_BIAS.t5 GND 0.018462f
C309 CS_BIAS.t7 GND 0.018462f
C310 CS_BIAS.n186 GND 0.1295f
C311 CS_BIAS.n187 GND 0.007421f
C312 CS_BIAS.t16 GND 0.165978f
C313 CS_BIAS.n188 GND 0.003322f
C314 CS_BIAS.n189 GND 0.005629f
C315 CS_BIAS.t12 GND 0.165978f
C316 CS_BIAS.n190 GND 0.011312f
C317 CS_BIAS.n191 GND 0.005629f
C318 CS_BIAS.n192 GND 0.00647f
C319 CS_BIAS.n193 GND 0.005629f
C320 CS_BIAS.n194 GND 0.009506f
C321 CS_BIAS.n195 GND 0.005629f
C322 CS_BIAS.t4 GND 0.165978f
C323 CS_BIAS.n196 GND 0.005451f
C324 CS_BIAS.n197 GND 0.005629f
C325 CS_BIAS.t22 GND 0.165978f
C326 CS_BIAS.n198 GND 0.077843f
C327 CS_BIAS.t20 GND 0.201331f
C328 CS_BIAS.n199 GND 0.076644f
C329 CS_BIAS.n200 GND 0.047175f
C330 CS_BIAS.n201 GND 0.006883f
C331 CS_BIAS.n202 GND 0.011312f
C332 CS_BIAS.n203 GND 0.004779f
C333 CS_BIAS.n204 GND 0.005629f
C334 CS_BIAS.n205 GND 0.005629f
C335 CS_BIAS.n206 GND 0.005629f
C336 CS_BIAS.n207 GND 0.011187f
C337 CS_BIAS.n208 GND 0.00647f
C338 CS_BIAS.n209 GND 0.064177f
C339 CS_BIAS.n210 GND 0.009253f
C340 CS_BIAS.n211 GND 0.005629f
C341 CS_BIAS.n212 GND 0.005629f
C342 CS_BIAS.n213 GND 0.005629f
C343 CS_BIAS.n214 GND 0.003279f
C344 CS_BIAS.n215 GND 0.009506f
C345 CS_BIAS.t6 GND 0.165978f
C346 CS_BIAS.n216 GND 0.064177f
C347 CS_BIAS.n217 GND 0.009253f
C348 CS_BIAS.n218 GND 0.005629f
C349 CS_BIAS.n219 GND 0.005629f
C350 CS_BIAS.n220 GND 0.005629f
C351 CS_BIAS.n221 GND 0.011187f
C352 CS_BIAS.n222 GND 0.005451f
C353 CS_BIAS.n223 GND 0.004779f
C354 CS_BIAS.n224 GND 0.005629f
C355 CS_BIAS.n225 GND 0.005629f
C356 CS_BIAS.n226 GND 0.005629f
C357 CS_BIAS.n227 GND 0.006883f
C358 CS_BIAS.n228 GND 0.064177f
C359 CS_BIAS.n229 GND 0.008841f
C360 CS_BIAS.n230 GND 0.009998f
C361 CS_BIAS.n231 GND 0.005629f
C362 CS_BIAS.n232 GND 0.005629f
C363 CS_BIAS.n233 GND 0.005629f
C364 CS_BIAS.n234 GND 0.008971f
C365 CS_BIAS.n235 GND 0.009665f
C366 CS_BIAS.n236 GND 0.082618f
C367 CS_BIAS.n237 GND 0.064948f
C368 CS_BIAS.t13 GND 0.018462f
C369 CS_BIAS.t17 GND 0.018462f
C370 CS_BIAS.n238 GND 0.1295f
C371 CS_BIAS.n239 GND 0.181834f
C372 CS_BIAS.n240 GND 0.311293f
C373 CS_BIAS.n241 GND 0.04069f
C374 CS_BIAS.n242 GND 0.003279f
C375 CS_BIAS.n243 GND 0.009506f
C376 CS_BIAS.t28 GND 0.165978f
C377 CS_BIAS.n244 GND 0.064177f
C378 CS_BIAS.n245 GND 0.009253f
C379 CS_BIAS.n246 GND 0.005629f
C380 CS_BIAS.n247 GND 0.005629f
C381 CS_BIAS.n248 GND 0.005629f
C382 CS_BIAS.n249 GND 0.011187f
C383 CS_BIAS.n250 GND 0.005451f
C384 CS_BIAS.n251 GND 0.004779f
C385 CS_BIAS.n252 GND 0.005629f
C386 CS_BIAS.n253 GND 0.005629f
C387 CS_BIAS.n254 GND 0.005629f
C388 CS_BIAS.n255 GND 0.006883f
C389 CS_BIAS.n256 GND 0.064177f
C390 CS_BIAS.n257 GND 0.008841f
C391 CS_BIAS.n258 GND 0.009998f
C392 CS_BIAS.n259 GND 0.005629f
C393 CS_BIAS.n260 GND 0.005629f
C394 CS_BIAS.n261 GND 0.005629f
C395 CS_BIAS.n262 GND 0.008971f
C396 CS_BIAS.n263 GND 0.009665f
C397 CS_BIAS.n264 GND 0.082618f
C398 CS_BIAS.n265 GND 0.034138f
C399 CS_BIAS.n266 GND 0.007421f
C400 CS_BIAS.t29 GND 0.165978f
C401 CS_BIAS.n267 GND 0.003322f
C402 CS_BIAS.n268 GND 0.005629f
C403 CS_BIAS.t45 GND 0.165978f
C404 CS_BIAS.n269 GND 0.011312f
C405 CS_BIAS.n270 GND 0.005629f
C406 CS_BIAS.n271 GND 0.00647f
C407 CS_BIAS.n272 GND 0.005629f
C408 CS_BIAS.n273 GND 0.009506f
C409 CS_BIAS.n274 GND 0.005629f
C410 CS_BIAS.t34 GND 0.165978f
C411 CS_BIAS.n275 GND 0.005451f
C412 CS_BIAS.n276 GND 0.005629f
C413 CS_BIAS.t41 GND 0.165978f
C414 CS_BIAS.n277 GND 0.077843f
C415 CS_BIAS.t31 GND 0.201331f
C416 CS_BIAS.n278 GND 0.076644f
C417 CS_BIAS.n279 GND 0.047175f
C418 CS_BIAS.n280 GND 0.006883f
C419 CS_BIAS.n281 GND 0.011312f
C420 CS_BIAS.n282 GND 0.004779f
C421 CS_BIAS.n283 GND 0.005629f
C422 CS_BIAS.n284 GND 0.005629f
C423 CS_BIAS.n285 GND 0.005629f
C424 CS_BIAS.n286 GND 0.011187f
C425 CS_BIAS.n287 GND 0.00647f
C426 CS_BIAS.n288 GND 0.064177f
C427 CS_BIAS.n289 GND 0.009253f
C428 CS_BIAS.n290 GND 0.005629f
C429 CS_BIAS.n291 GND 0.005629f
C430 CS_BIAS.n292 GND 0.005629f
C431 CS_BIAS.n293 GND 0.003279f
C432 CS_BIAS.n294 GND 0.009506f
C433 CS_BIAS.t46 GND 0.165978f
C434 CS_BIAS.n295 GND 0.064177f
C435 CS_BIAS.n296 GND 0.009253f
C436 CS_BIAS.n297 GND 0.005629f
C437 CS_BIAS.n298 GND 0.005629f
C438 CS_BIAS.n299 GND 0.005629f
C439 CS_BIAS.n300 GND 0.011187f
C440 CS_BIAS.n301 GND 0.005451f
C441 CS_BIAS.n302 GND 0.004779f
C442 CS_BIAS.n303 GND 0.005629f
C443 CS_BIAS.n304 GND 0.005629f
C444 CS_BIAS.n305 GND 0.005629f
C445 CS_BIAS.n306 GND 0.006883f
C446 CS_BIAS.n307 GND 0.064177f
C447 CS_BIAS.n308 GND 0.008841f
C448 CS_BIAS.n309 GND 0.009998f
C449 CS_BIAS.n310 GND 0.005629f
C450 CS_BIAS.n311 GND 0.005629f
C451 CS_BIAS.n312 GND 0.005629f
C452 CS_BIAS.n313 GND 0.008971f
C453 CS_BIAS.n314 GND 0.009665f
C454 CS_BIAS.n315 GND 0.082618f
C455 CS_BIAS.n316 GND 0.020913f
C456 CS_BIAS.n317 GND 0.153844f
C457 CS_BIAS.n318 GND 3.72266f
C458 VOUT.t12 GND 0.032674f
C459 VOUT.t9 GND 0.032674f
C460 VOUT.n0 GND 0.166876f
C461 VOUT.t27 GND 0.210121f
C462 VOUT.n1 GND 1.12414f
C463 VOUT.t43 GND 0.032674f
C464 VOUT.t8 GND 0.032674f
C465 VOUT.n2 GND 0.166876f
C466 VOUT.t6 GND 0.210121f
C467 VOUT.n3 GND 1.09246f
C468 VOUT.n4 GND 0.491979f
C469 VOUT.t20 GND 0.032674f
C470 VOUT.t37 GND 0.032674f
C471 VOUT.n5 GND 0.166876f
C472 VOUT.t36 GND 0.210121f
C473 VOUT.n6 GND 1.09246f
C474 VOUT.n7 GND 0.340891f
C475 VOUT.t32 GND 0.032674f
C476 VOUT.t42 GND 0.032674f
C477 VOUT.n8 GND 0.166876f
C478 VOUT.t14 GND 0.210121f
C479 VOUT.n9 GND 1.09246f
C480 VOUT.n10 GND 0.544407f
C481 VOUT.n11 GND 7.01774f
C482 VOUT.t48 GND 15.1181f
C483 VOUT.n12 GND 9.8358f
C484 VOUT.t49 GND 15.4461f
C485 VOUT.t51 GND 15.5337f
C486 VOUT.n13 GND 10.919499f
C487 VOUT.n14 GND 11.026299f
C488 VOUT.t50 GND 15.1181f
C489 VOUT.n15 GND 4.88334f
C490 VOUT.n16 GND 10.4176f
C491 VOUT.n17 GND 1.91574f
C492 VOUT.t41 GND 0.213948f
C493 VOUT.t7 GND 0.032674f
C494 VOUT.t44 GND 0.032674f
C495 VOUT.n18 GND 0.160408f
C496 VOUT.n19 GND 1.10189f
C497 VOUT.t38 GND 0.213948f
C498 VOUT.t5 GND 0.032674f
C499 VOUT.t1 GND 0.032674f
C500 VOUT.n20 GND 0.160408f
C501 VOUT.n21 GND 1.06936f
C502 VOUT.n22 GND 0.54261f
C503 VOUT.t39 GND 0.213948f
C504 VOUT.t11 GND 0.032674f
C505 VOUT.t24 GND 0.032674f
C506 VOUT.n23 GND 0.160408f
C507 VOUT.n24 GND 1.06936f
C508 VOUT.n25 GND 0.366634f
C509 VOUT.t40 GND 0.213948f
C510 VOUT.t10 GND 0.032674f
C511 VOUT.t28 GND 0.032674f
C512 VOUT.n26 GND 0.160407f
C513 VOUT.n27 GND 1.06936f
C514 VOUT.n28 GND 0.57015f
C515 VOUT.n29 GND 9.314031f
C516 VOUT.t23 GND 0.048419f
C517 VOUT.t47 GND 0.048419f
C518 VOUT.n30 GND 0.344105f
C519 VOUT.t13 GND 0.048419f
C520 VOUT.t45 GND 0.048419f
C521 VOUT.n31 GND 0.339622f
C522 VOUT.n32 GND 0.728135f
C523 VOUT.t18 GND 0.048419f
C524 VOUT.t15 GND 0.048419f
C525 VOUT.n33 GND 0.339622f
C526 VOUT.n34 GND 0.505454f
C527 VOUT.t35 GND 0.048419f
C528 VOUT.t16 GND 0.048419f
C529 VOUT.n35 GND 0.344105f
C530 VOUT.t30 GND 0.048419f
C531 VOUT.t21 GND 0.048419f
C532 VOUT.n36 GND 0.339622f
C533 VOUT.n37 GND 0.728135f
C534 VOUT.t17 GND 0.048419f
C535 VOUT.t0 GND 0.048419f
C536 VOUT.n38 GND 0.339622f
C537 VOUT.n39 GND 0.459312f
C538 VOUT.n40 GND 1.02699f
C539 VOUT.n41 GND 8.936719f
C540 VOUT.t25 GND 0.048419f
C541 VOUT.t34 GND 0.048419f
C542 VOUT.n42 GND 0.344105f
C543 VOUT.t29 GND 0.048419f
C544 VOUT.t2 GND 0.048419f
C545 VOUT.n43 GND 0.339622f
C546 VOUT.n44 GND 0.728135f
C547 VOUT.t31 GND 0.048419f
C548 VOUT.t46 GND 0.048419f
C549 VOUT.n45 GND 0.339622f
C550 VOUT.n46 GND 0.505454f
C551 VOUT.t33 GND 0.048419f
C552 VOUT.t4 GND 0.048419f
C553 VOUT.n47 GND 0.344105f
C554 VOUT.t3 GND 0.048419f
C555 VOUT.t22 GND 0.048419f
C556 VOUT.n48 GND 0.339622f
C557 VOUT.n49 GND 0.728135f
C558 VOUT.t26 GND 0.048419f
C559 VOUT.t19 GND 0.048419f
C560 VOUT.n50 GND 0.339622f
C561 VOUT.n51 GND 0.459312f
C562 VOUT.n52 GND 1.02699f
C563 VOUT.n53 GND 6.34464f
C564 VOUT.n54 GND 5.04806f
C565 VDD.t33 GND 0.011218f
C566 VDD.t31 GND 0.011218f
C567 VDD.n0 GND 0.048575f
C568 VDD.t39 GND 0.011218f
C569 VDD.t49 GND 0.011218f
C570 VDD.n1 GND 0.046694f
C571 VDD.n2 GND 0.592781f
C572 VDD.t41 GND 0.011218f
C573 VDD.t18 GND 0.011218f
C574 VDD.n3 GND 0.046694f
C575 VDD.n4 GND 0.307594f
C576 VDD.t29 GND 0.011218f
C577 VDD.t27 GND 0.011218f
C578 VDD.n5 GND 0.046694f
C579 VDD.n6 GND 0.26114f
C580 VDD.t37 GND 0.011218f
C581 VDD.t25 GND 0.011218f
C582 VDD.n7 GND 0.048575f
C583 VDD.t43 GND 0.011218f
C584 VDD.t47 GND 0.011218f
C585 VDD.n8 GND 0.046694f
C586 VDD.n9 GND 0.592781f
C587 VDD.t20 GND 0.011218f
C588 VDD.t45 GND 0.011218f
C589 VDD.n10 GND 0.046694f
C590 VDD.n11 GND 0.307594f
C591 VDD.t35 GND 0.011218f
C592 VDD.t22 GND 0.011218f
C593 VDD.n12 GND 0.046694f
C594 VDD.n13 GND 0.26114f
C595 VDD.n14 GND 0.187854f
C596 VDD.n15 GND 2.19181f
C597 VDD.t142 GND 0.018389f
C598 VDD.t6 GND 0.018389f
C599 VDD.n16 GND 0.077578f
C600 VDD.t145 GND 0.101282f
C601 VDD.n17 GND 0.594126f
C602 VDD.t138 GND 0.018389f
C603 VDD.t3 GND 0.018389f
C604 VDD.n18 GND 0.077578f
C605 VDD.t1 GND 0.101282f
C606 VDD.n19 GND 0.576056f
C607 VDD.n20 GND 0.27325f
C608 VDD.t139 GND 0.018389f
C609 VDD.t11 GND 0.018389f
C610 VDD.n21 GND 0.077578f
C611 VDD.t51 GND 0.101282f
C612 VDD.n22 GND 0.576056f
C613 VDD.n23 GND 0.190156f
C614 VDD.t141 GND 0.018389f
C615 VDD.t10 GND 0.018389f
C616 VDD.n24 GND 0.077578f
C617 VDD.t133 GND 0.101282f
C618 VDD.n25 GND 0.576056f
C619 VDD.n26 GND 0.267329f
C620 VDD.n27 GND 0.006342f
C621 VDD.n28 GND 0.006342f
C622 VDD.n29 GND 0.005122f
C623 VDD.n30 GND 0.005122f
C624 VDD.n31 GND 0.006364f
C625 VDD.n32 GND 0.006364f
C626 VDD.n33 GND 0.471559f
C627 VDD.n34 GND 0.006364f
C628 VDD.n35 GND 0.006364f
C629 VDD.n36 GND 0.006364f
C630 VDD.n37 GND 0.471559f
C631 VDD.n38 GND 0.006364f
C632 VDD.n39 GND 0.006364f
C633 VDD.n40 GND 0.006364f
C634 VDD.n41 GND 0.006364f
C635 VDD.n42 GND 0.005122f
C636 VDD.n43 GND 0.006364f
C637 VDD.n44 GND 0.006364f
C638 VDD.n45 GND 0.006364f
C639 VDD.n46 GND 0.006364f
C640 VDD.n47 GND 0.471559f
C641 VDD.n48 GND 0.006364f
C642 VDD.n49 GND 0.006364f
C643 VDD.n50 GND 0.006364f
C644 VDD.n51 GND 0.006364f
C645 VDD.n52 GND 0.006364f
C646 VDD.n53 GND 0.005122f
C647 VDD.n54 GND 0.006364f
C648 VDD.n55 GND 0.006364f
C649 VDD.n56 GND 0.006364f
C650 VDD.n57 GND 0.006364f
C651 VDD.n58 GND 0.471559f
C652 VDD.n59 GND 0.006364f
C653 VDD.n60 GND 0.006364f
C654 VDD.n61 GND 0.006364f
C655 VDD.n62 GND 0.006364f
C656 VDD.n63 GND 0.006364f
C657 VDD.n64 GND 0.005122f
C658 VDD.n65 GND 0.006364f
C659 VDD.n66 GND 0.006364f
C660 VDD.n67 GND 0.006364f
C661 VDD.n68 GND 0.006364f
C662 VDD.n69 GND 0.471559f
C663 VDD.n70 GND 0.006364f
C664 VDD.n71 GND 0.006364f
C665 VDD.n72 GND 0.006364f
C666 VDD.n73 GND 0.006364f
C667 VDD.n74 GND 0.006364f
C668 VDD.n75 GND 0.005122f
C669 VDD.n76 GND 0.006364f
C670 VDD.n77 GND 0.006364f
C671 VDD.n78 GND 0.006364f
C672 VDD.n79 GND 0.006364f
C673 VDD.n80 GND 0.471559f
C674 VDD.n81 GND 0.006364f
C675 VDD.n82 GND 0.006364f
C676 VDD.n83 GND 0.006364f
C677 VDD.n84 GND 0.006364f
C678 VDD.n85 GND 0.006364f
C679 VDD.n86 GND 0.005122f
C680 VDD.n87 GND 0.006364f
C681 VDD.n88 GND 0.006364f
C682 VDD.n89 GND 0.006364f
C683 VDD.n90 GND 0.006364f
C684 VDD.n91 GND 0.471559f
C685 VDD.n92 GND 0.006364f
C686 VDD.n93 GND 0.006364f
C687 VDD.n94 GND 0.006364f
C688 VDD.n95 GND 0.006364f
C689 VDD.n96 GND 0.006364f
C690 VDD.n97 GND 0.005122f
C691 VDD.n98 GND 0.006364f
C692 VDD.n99 GND 0.006364f
C693 VDD.n100 GND 0.006364f
C694 VDD.n101 GND 0.014395f
C695 VDD.n102 GND 1.01857f
C696 VDD.n103 GND 0.01437f
C697 VDD.n104 GND 0.006364f
C698 VDD.n105 GND 0.006364f
C699 VDD.n106 GND 0.006364f
C700 VDD.n107 GND 0.006364f
C701 VDD.n108 GND 0.005122f
C702 VDD.n110 GND 0.006364f
C703 VDD.n111 GND 0.006364f
C704 VDD.n112 GND 0.006364f
C705 VDD.n113 GND 0.006364f
C706 VDD.n114 GND 0.006364f
C707 VDD.n115 GND 0.005122f
C708 VDD.n117 GND 0.006364f
C709 VDD.n118 GND 0.006364f
C710 VDD.n119 GND 0.006364f
C711 VDD.n120 GND 0.006364f
C712 VDD.n121 GND 0.006364f
C713 VDD.t87 GND 0.123904f
C714 VDD.t86 GND 0.415248f
C715 VDD.n122 GND 0.086184f
C716 VDD.t88 GND 0.090617f
C717 VDD.n123 GND 0.088946f
C718 VDD.n124 GND 0.009604f
C719 VDD.n126 GND 0.006364f
C720 VDD.n127 GND 0.006364f
C721 VDD.n128 GND 0.006364f
C722 VDD.n129 GND 0.006364f
C723 VDD.n130 GND 0.006364f
C724 VDD.n131 GND 0.005122f
C725 VDD.n133 GND 0.006364f
C726 VDD.n134 GND 0.006364f
C727 VDD.n135 GND 0.006364f
C728 VDD.n136 GND 0.006364f
C729 VDD.n137 GND 0.006364f
C730 VDD.n138 GND 0.005122f
C731 VDD.n140 GND 0.006364f
C732 VDD.n141 GND 0.006364f
C733 VDD.n142 GND 0.006364f
C734 VDD.n143 GND 0.006364f
C735 VDD.n144 GND 0.006364f
C736 VDD.n145 GND 0.005122f
C737 VDD.n147 GND 0.006364f
C738 VDD.n148 GND 0.006364f
C739 VDD.n149 GND 0.006364f
C740 VDD.n150 GND 0.006364f
C741 VDD.n151 GND 0.006364f
C742 VDD.n152 GND 0.005122f
C743 VDD.n154 GND 0.006364f
C744 VDD.n155 GND 0.006364f
C745 VDD.n156 GND 0.006364f
C746 VDD.n157 GND 0.006364f
C747 VDD.n158 GND 0.006364f
C748 VDD.n159 GND 0.005122f
C749 VDD.n161 GND 0.006364f
C750 VDD.n162 GND 0.006364f
C751 VDD.n163 GND 0.006364f
C752 VDD.n164 GND 0.006364f
C753 VDD.n165 GND 0.006364f
C754 VDD.n166 GND 0.005122f
C755 VDD.n168 GND 0.006364f
C756 VDD.n169 GND 0.006364f
C757 VDD.n170 GND 0.006364f
C758 VDD.n171 GND 0.006364f
C759 VDD.n172 GND 0.006364f
C760 VDD.n173 GND 0.002689f
C761 VDD.n175 GND 0.006364f
C762 VDD.t130 GND 0.123904f
C763 VDD.t129 GND 0.415248f
C764 VDD.n176 GND 0.086184f
C765 VDD.t131 GND 0.090617f
C766 VDD.n177 GND 0.088946f
C767 VDD.n178 GND 0.007043f
C768 VDD.n179 GND 0.006364f
C769 VDD.n180 GND 0.006364f
C770 VDD.n181 GND 0.006364f
C771 VDD.n182 GND 0.006364f
C772 VDD.n183 GND 0.005122f
C773 VDD.n185 GND 0.006364f
C774 VDD.n186 GND 0.006364f
C775 VDD.n187 GND 0.006364f
C776 VDD.n188 GND 0.006364f
C777 VDD.n189 GND 0.006364f
C778 VDD.n190 GND 0.005122f
C779 VDD.n192 GND 0.006364f
C780 VDD.n193 GND 0.006364f
C781 VDD.n194 GND 0.006364f
C782 VDD.n195 GND 0.006364f
C783 VDD.n196 GND 0.006364f
C784 VDD.n197 GND 0.005122f
C785 VDD.n199 GND 0.006364f
C786 VDD.n200 GND 0.006364f
C787 VDD.n201 GND 0.006364f
C788 VDD.n202 GND 0.006364f
C789 VDD.n203 GND 0.006364f
C790 VDD.n204 GND 0.006364f
C791 VDD.n205 GND 0.005122f
C792 VDD.n206 GND 0.006364f
C793 VDD.n207 GND 0.006364f
C794 VDD.n208 GND 0.005122f
C795 VDD.n209 GND 0.006364f
C796 VDD.n210 GND 0.006364f
C797 VDD.n211 GND 0.005122f
C798 VDD.n212 GND 0.006364f
C799 VDD.n213 GND 0.006364f
C800 VDD.n214 GND 0.005122f
C801 VDD.n215 GND 0.006364f
C802 VDD.n216 GND 0.006364f
C803 VDD.n217 GND 0.005122f
C804 VDD.n218 GND 0.006364f
C805 VDD.n219 GND 0.006364f
C806 VDD.n220 GND 0.005122f
C807 VDD.n221 GND 0.006364f
C808 VDD.n222 GND 0.005122f
C809 VDD.n223 GND 0.006364f
C810 VDD.n224 GND 0.005122f
C811 VDD.n225 GND 0.006364f
C812 VDD.n226 GND 0.006364f
C813 VDD.n227 GND 0.471559f
C814 VDD.n228 GND 0.006364f
C815 VDD.n229 GND 0.005122f
C816 VDD.n230 GND 0.006364f
C817 VDD.n231 GND 0.005122f
C818 VDD.n232 GND 0.006364f
C819 VDD.n233 GND 0.471559f
C820 VDD.n234 GND 0.006364f
C821 VDD.n235 GND 0.005122f
C822 VDD.n236 GND 0.006364f
C823 VDD.n237 GND 0.005122f
C824 VDD.n238 GND 0.006364f
C825 VDD.n239 GND 0.471559f
C826 VDD.n240 GND 0.006364f
C827 VDD.n241 GND 0.005122f
C828 VDD.n242 GND 0.006364f
C829 VDD.n243 GND 0.005122f
C830 VDD.n244 GND 0.006364f
C831 VDD.t137 GND 0.235779f
C832 VDD.n245 GND 0.006364f
C833 VDD.n246 GND 0.005122f
C834 VDD.n247 GND 0.006364f
C835 VDD.n248 GND 0.005122f
C836 VDD.n249 GND 0.006364f
C837 VDD.n250 GND 0.471559f
C838 VDD.n251 GND 0.240495f
C839 VDD.n252 GND 0.006364f
C840 VDD.n253 GND 0.005122f
C841 VDD.n254 GND 0.006364f
C842 VDD.n255 GND 0.005122f
C843 VDD.n256 GND 0.006364f
C844 VDD.n257 GND 0.471559f
C845 VDD.n258 GND 0.006364f
C846 VDD.n259 GND 0.005122f
C847 VDD.n260 GND 0.006364f
C848 VDD.n261 GND 0.005122f
C849 VDD.n262 GND 0.006364f
C850 VDD.n263 GND 0.471559f
C851 VDD.n264 GND 0.006364f
C852 VDD.n265 GND 0.005122f
C853 VDD.n266 GND 0.006364f
C854 VDD.n267 GND 0.005122f
C855 VDD.n268 GND 0.006364f
C856 VDD.n269 GND 0.471559f
C857 VDD.n270 GND 0.006364f
C858 VDD.n271 GND 0.005122f
C859 VDD.n272 GND 0.006364f
C860 VDD.n273 GND 0.005122f
C861 VDD.n274 GND 0.006364f
C862 VDD.n275 GND 0.471559f
C863 VDD.n276 GND 0.006364f
C864 VDD.n277 GND 0.005122f
C865 VDD.n278 GND 0.006364f
C866 VDD.n279 GND 0.005122f
C867 VDD.n280 GND 0.006364f
C868 VDD.t83 GND 0.235779f
C869 VDD.n281 GND 0.006364f
C870 VDD.n282 GND 0.005122f
C871 VDD.n283 GND 0.006364f
C872 VDD.n284 GND 0.005122f
C873 VDD.n285 GND 0.006364f
C874 VDD.n286 GND 0.471559f
C875 VDD.n287 GND 0.282935f
C876 VDD.n288 GND 0.006364f
C877 VDD.n289 GND 0.005122f
C878 VDD.n290 GND 0.006364f
C879 VDD.n291 GND 0.005122f
C880 VDD.n292 GND 0.006364f
C881 VDD.n293 GND 0.471559f
C882 VDD.n294 GND 0.006364f
C883 VDD.n295 GND 0.005122f
C884 VDD.n296 GND 0.01437f
C885 VDD.n297 GND 0.01437f
C886 VDD.n298 GND 3.33628f
C887 VDD.n299 GND 0.01437f
C888 VDD.n300 GND 0.006364f
C889 VDD.n301 GND 0.005122f
C890 VDD.n303 GND 0.006364f
C891 VDD.n304 GND 0.006364f
C892 VDD.n305 GND 0.006364f
C893 VDD.n306 GND 0.005122f
C894 VDD.n307 GND 0.006364f
C895 VDD.n308 GND 0.006364f
C896 VDD.n309 GND 0.006364f
C897 VDD.n310 GND 0.006364f
C898 VDD.n311 GND 0.004837f
C899 VDD.n312 GND 0.005122f
C900 VDD.n313 GND 0.006364f
C901 VDD.n314 GND 1.50188f
C902 VDD.t85 GND 0.123904f
C903 VDD.t82 GND 0.415248f
C904 VDD.n315 GND 0.086184f
C905 VDD.t84 GND 0.090617f
C906 VDD.n316 GND 0.088946f
C907 VDD.n318 GND 0.006364f
C908 VDD.n319 GND 0.004709f
C909 VDD.n320 GND 0.005122f
C910 VDD.n322 GND 0.006364f
C911 VDD.n323 GND 0.006364f
C912 VDD.n324 GND 0.006364f
C913 VDD.n325 GND 0.005122f
C914 VDD.n326 GND 0.006364f
C915 VDD.n327 GND 0.006364f
C916 VDD.n328 GND 0.006364f
C917 VDD.n329 GND 0.006364f
C918 VDD.n330 GND 0.006364f
C919 VDD.n331 GND 0.005122f
C920 VDD.n332 GND 0.006364f
C921 VDD.n333 GND 0.006364f
C922 VDD.n334 GND 0.006364f
C923 VDD.n335 GND 0.006364f
C924 VDD.n336 GND 0.006364f
C925 VDD.n337 GND 0.002587f
C926 VDD.n338 GND 0.006364f
C927 VDD.t112 GND 0.123904f
C928 VDD.t110 GND 0.415248f
C929 VDD.n339 GND 0.086184f
C930 VDD.t111 GND 0.090617f
C931 VDD.n340 GND 0.088946f
C932 VDD.n341 GND 0.007043f
C933 VDD.n342 GND 0.006364f
C934 VDD.n343 GND 0.006364f
C935 VDD.n344 GND 0.006364f
C936 VDD.n345 GND 0.006364f
C937 VDD.n346 GND 0.005122f
C938 VDD.n347 GND 0.006364f
C939 VDD.n348 GND 0.006364f
C940 VDD.n349 GND 0.006364f
C941 VDD.n350 GND 0.006364f
C942 VDD.n351 GND 0.006364f
C943 VDD.n352 GND 0.005122f
C944 VDD.n353 GND 0.006364f
C945 VDD.n354 GND 0.006364f
C946 VDD.n355 GND 0.006364f
C947 VDD.n356 GND 0.006364f
C948 VDD.n357 GND 0.006364f
C949 VDD.n358 GND 0.005122f
C950 VDD.n359 GND 0.006364f
C951 VDD.n360 GND 0.006364f
C952 VDD.n361 GND 0.006364f
C953 VDD.n362 GND 0.006364f
C954 VDD.n363 GND 0.006364f
C955 VDD.n364 GND 0.005122f
C956 VDD.n365 GND 0.006364f
C957 VDD.n366 GND 0.005122f
C958 VDD.n367 GND 0.004709f
C959 VDD.n368 GND 0.004837f
C960 VDD.n369 GND 0.003246f
C961 VDD.n370 GND 0.004328f
C962 VDD.n371 GND 0.004328f
C963 VDD.t140 GND 5.46301f
C964 VDD.t24 GND 4.31005f
C965 VDD.t36 GND 3.64043f
C966 VDD.t46 GND 3.64043f
C967 VDD.t42 GND 3.17123f
C968 VDD.n372 GND 1.60801f
C969 VDD.n373 GND 0.004328f
C970 VDD.n374 GND 0.004328f
C971 VDD.t76 GND 0.066005f
C972 VDD.t74 GND 0.213596f
C973 VDD.n375 GND 0.071628f
C974 VDD.t77 GND 0.048572f
C975 VDD.n376 GND 0.068504f
C976 VDD.n377 GND 0.004328f
C977 VDD.n379 GND 0.009986f
C978 VDD.n380 GND 0.004328f
C979 VDD.n381 GND 0.004328f
C980 VDD.n382 GND 0.32066f
C981 VDD.n383 GND 0.004328f
C982 VDD.n384 GND 0.417329f
C983 VDD.n385 GND 0.004328f
C984 VDD.n386 GND 0.004328f
C985 VDD.n387 GND 0.009986f
C986 VDD.n388 GND 0.004328f
C987 VDD.n389 GND 0.004328f
C988 VDD.n390 GND 0.004328f
C989 VDD.n391 GND 0.004328f
C990 VDD.n392 GND 0.004328f
C991 VDD.n394 GND 0.004328f
C992 VDD.n395 GND 0.004328f
C993 VDD.n397 GND 0.004328f
C994 VDD.t108 GND 0.066005f
C995 VDD.t107 GND 0.213596f
C996 VDD.n398 GND 0.071628f
C997 VDD.t109 GND 0.048572f
C998 VDD.n399 GND 0.068504f
C999 VDD.n400 GND 0.004328f
C1000 VDD.n402 GND 0.009986f
C1001 VDD.n403 GND 0.004328f
C1002 VDD.n404 GND 0.004328f
C1003 VDD.n405 GND 0.32066f
C1004 VDD.n406 GND 0.004328f
C1005 VDD.n407 GND 0.004328f
C1006 VDD.n408 GND 0.004328f
C1007 VDD.n409 GND 0.004328f
C1008 VDD.n410 GND 0.004328f
C1009 VDD.n411 GND 0.264073f
C1010 VDD.n412 GND 0.004328f
C1011 VDD.n413 GND 0.004328f
C1012 VDD.n414 GND 0.004328f
C1013 VDD.n415 GND 0.004328f
C1014 VDD.n416 GND 0.004328f
C1015 VDD.n417 GND 0.004328f
C1016 VDD.t75 GND 0.16033f
C1017 VDD.n418 GND 0.004328f
C1018 VDD.n419 GND 0.004328f
C1019 VDD.t44 GND 0.16033f
C1020 VDD.n420 GND 0.004328f
C1021 VDD.n421 GND 0.004328f
C1022 VDD.n422 GND 0.004328f
C1023 VDD.n423 GND 0.32066f
C1024 VDD.n424 GND 0.004328f
C1025 VDD.n425 GND 0.004328f
C1026 VDD.n426 GND 0.24521f
C1027 VDD.n427 GND 0.004328f
C1028 VDD.n428 GND 0.004328f
C1029 VDD.n429 GND 0.004328f
C1030 VDD.n430 GND 0.32066f
C1031 VDD.n431 GND 0.004328f
C1032 VDD.n432 GND 0.004328f
C1033 VDD.n433 GND 0.004328f
C1034 VDD.n434 GND 0.004328f
C1035 VDD.n435 GND 0.004328f
C1036 VDD.n436 GND 0.32066f
C1037 VDD.n437 GND 0.004328f
C1038 VDD.n438 GND 0.004328f
C1039 VDD.n439 GND 0.004328f
C1040 VDD.n440 GND 0.004328f
C1041 VDD.n441 GND 0.004328f
C1042 VDD.n442 GND 0.32066f
C1043 VDD.n443 GND 0.004328f
C1044 VDD.n444 GND 0.004328f
C1045 VDD.n445 GND 0.004328f
C1046 VDD.n446 GND 0.004328f
C1047 VDD.n447 GND 0.004328f
C1048 VDD.t19 GND 0.32066f
C1049 VDD.n448 GND 0.004328f
C1050 VDD.n449 GND 0.004328f
C1051 VDD.n450 GND 0.004328f
C1052 VDD.n451 GND 0.004328f
C1053 VDD.n452 GND 0.004328f
C1054 VDD.n453 GND 0.32066f
C1055 VDD.n454 GND 0.004328f
C1056 VDD.n455 GND 0.004328f
C1057 VDD.n456 GND 0.004328f
C1058 VDD.n457 GND 0.004328f
C1059 VDD.n458 GND 0.004328f
C1060 VDD.n459 GND 0.32066f
C1061 VDD.n460 GND 0.004328f
C1062 VDD.n461 GND 0.004328f
C1063 VDD.n462 GND 0.004328f
C1064 VDD.n463 GND 0.004328f
C1065 VDD.n464 GND 0.004328f
C1066 VDD.n465 GND 0.32066f
C1067 VDD.n466 GND 0.004328f
C1068 VDD.n467 GND 0.004328f
C1069 VDD.n468 GND 0.004328f
C1070 VDD.n469 GND 0.004328f
C1071 VDD.n470 GND 0.004328f
C1072 VDD.n471 GND 0.32066f
C1073 VDD.n472 GND 0.004328f
C1074 VDD.n473 GND 0.004328f
C1075 VDD.n474 GND 0.004328f
C1076 VDD.n475 GND 0.004328f
C1077 VDD.n476 GND 0.004328f
C1078 VDD.n477 GND 0.32066f
C1079 VDD.n478 GND 0.004328f
C1080 VDD.n479 GND 0.004328f
C1081 VDD.n480 GND 0.004328f
C1082 VDD.n481 GND 0.004328f
C1083 VDD.n482 GND 0.004328f
C1084 VDD.t21 GND 0.16033f
C1085 VDD.n483 GND 0.004328f
C1086 VDD.n484 GND 0.004328f
C1087 VDD.n485 GND 0.004328f
C1088 VDD.n486 GND 0.004328f
C1089 VDD.n487 GND 0.004328f
C1090 VDD.n488 GND 0.32066f
C1091 VDD.n489 GND 0.004328f
C1092 VDD.n490 GND 0.004328f
C1093 VDD.n491 GND 0.264073f
C1094 VDD.n492 GND 0.004328f
C1095 VDD.n493 GND 0.004328f
C1096 VDD.n494 GND 0.004328f
C1097 VDD.n495 GND 0.32066f
C1098 VDD.n496 GND 0.004328f
C1099 VDD.n497 GND 0.004328f
C1100 VDD.n498 GND 0.004328f
C1101 VDD.n499 GND 0.004328f
C1102 VDD.n500 GND 0.004328f
C1103 VDD.n501 GND 0.32066f
C1104 VDD.n502 GND 0.004328f
C1105 VDD.n503 GND 0.004328f
C1106 VDD.n504 GND 0.004328f
C1107 VDD.n505 GND 0.004328f
C1108 VDD.n506 GND 0.004328f
C1109 VDD.n507 GND 0.24521f
C1110 VDD.n508 GND 0.004328f
C1111 VDD.n509 GND 0.004328f
C1112 VDD.n510 GND 0.004328f
C1113 VDD.n511 GND 0.004328f
C1114 VDD.n512 GND 0.004328f
C1115 VDD.n513 GND 0.273504f
C1116 VDD.n514 GND 0.004328f
C1117 VDD.n515 GND 0.004328f
C1118 VDD.t53 GND 0.16033f
C1119 VDD.n516 GND 0.004328f
C1120 VDD.n517 GND 0.004328f
C1121 VDD.n518 GND 0.004328f
C1122 VDD.n519 GND 0.32066f
C1123 VDD.n520 GND 0.004328f
C1124 VDD.n521 GND 0.004328f
C1125 VDD.t34 GND 0.16033f
C1126 VDD.n522 GND 0.004328f
C1127 VDD.n523 GND 0.004328f
C1128 VDD.n524 GND 0.004328f
C1129 VDD.n525 GND 0.32066f
C1130 VDD.n526 GND 0.004328f
C1131 VDD.n527 GND 0.004328f
C1132 VDD.n528 GND 0.004328f
C1133 VDD.n529 GND 0.009986f
C1134 VDD.n530 GND 0.009986f
C1135 VDD.n531 GND 0.417329f
C1136 VDD.n532 GND 0.004328f
C1137 VDD.n533 GND 0.004328f
C1138 VDD.n534 GND 0.009986f
C1139 VDD.n535 GND 0.004328f
C1140 VDD.n536 GND 0.004328f
C1141 VDD.n537 GND 0.417329f
C1142 VDD.n553 GND 0.010125f
C1143 VDD.n554 GND 0.009986f
C1144 VDD.n555 GND 0.004328f
C1145 VDD.n556 GND 0.009986f
C1146 VDD.t80 GND 0.066005f
C1147 VDD.t78 GND 0.213596f
C1148 VDD.n557 GND 0.071628f
C1149 VDD.t81 GND 0.048572f
C1150 VDD.n558 GND 0.068504f
C1151 VDD.n559 GND 0.004328f
C1152 VDD.n560 GND 0.004328f
C1153 VDD.n561 GND 0.32066f
C1154 VDD.n562 GND 0.004328f
C1155 VDD.n563 GND 0.004328f
C1156 VDD.n564 GND 0.004328f
C1157 VDD.n565 GND 0.009986f
C1158 VDD.n566 GND 0.004328f
C1159 VDD.t117 GND 0.066005f
C1160 VDD.t116 GND 0.213596f
C1161 VDD.n567 GND 0.071628f
C1162 VDD.t118 GND 0.048572f
C1163 VDD.n568 GND 0.068504f
C1164 VDD.n569 GND 0.00534f
C1165 VDD.n570 GND 0.004328f
C1166 VDD.n571 GND 0.004328f
C1167 VDD.n572 GND 0.32066f
C1168 VDD.n573 GND 0.004328f
C1169 VDD.n574 GND 0.004328f
C1170 VDD.n575 GND 0.004328f
C1171 VDD.n576 GND 0.004328f
C1172 VDD.n577 GND 0.004328f
C1173 VDD.t26 GND 0.16033f
C1174 VDD.n578 GND 0.004328f
C1175 VDD.n579 GND 0.004328f
C1176 VDD.n580 GND 0.004328f
C1177 VDD.n581 GND 0.004328f
C1178 VDD.n582 GND 0.004328f
C1179 VDD.n583 GND 0.004328f
C1180 VDD.t79 GND 0.16033f
C1181 VDD.n584 GND 0.004328f
C1182 VDD.n585 GND 0.004328f
C1183 VDD.n586 GND 0.273504f
C1184 VDD.n587 GND 0.004328f
C1185 VDD.n588 GND 0.004328f
C1186 VDD.n589 GND 0.004328f
C1187 VDD.n590 GND 0.32066f
C1188 VDD.n591 GND 0.004328f
C1189 VDD.n592 GND 0.004328f
C1190 VDD.n593 GND 0.24521f
C1191 VDD.n594 GND 0.004328f
C1192 VDD.n595 GND 0.004328f
C1193 VDD.n596 GND 0.004328f
C1194 VDD.n597 GND 0.32066f
C1195 VDD.n598 GND 0.004328f
C1196 VDD.n599 GND 0.004328f
C1197 VDD.n600 GND 0.004328f
C1198 VDD.n601 GND 0.004328f
C1199 VDD.n602 GND 0.004328f
C1200 VDD.n603 GND 0.32066f
C1201 VDD.n604 GND 0.004328f
C1202 VDD.n605 GND 0.004328f
C1203 VDD.n606 GND 0.004328f
C1204 VDD.n607 GND 0.004328f
C1205 VDD.n608 GND 0.004328f
C1206 VDD.n609 GND 0.264073f
C1207 VDD.n610 GND 0.004328f
C1208 VDD.n611 GND 0.004328f
C1209 VDD.n612 GND 0.004328f
C1210 VDD.n613 GND 0.004328f
C1211 VDD.n614 GND 0.004328f
C1212 VDD.n615 GND 0.32066f
C1213 VDD.n616 GND 0.004328f
C1214 VDD.n617 GND 0.004328f
C1215 VDD.t28 GND 0.16033f
C1216 VDD.n618 GND 0.004328f
C1217 VDD.n619 GND 0.004328f
C1218 VDD.n620 GND 0.004328f
C1219 VDD.n621 GND 0.32066f
C1220 VDD.n622 GND 0.004328f
C1221 VDD.n623 GND 0.004328f
C1222 VDD.n624 GND 0.004328f
C1223 VDD.n625 GND 0.004328f
C1224 VDD.n626 GND 0.004328f
C1225 VDD.n627 GND 0.32066f
C1226 VDD.n628 GND 0.004328f
C1227 VDD.n629 GND 0.004328f
C1228 VDD.n630 GND 0.004328f
C1229 VDD.n631 GND 0.004328f
C1230 VDD.n632 GND 0.004328f
C1231 VDD.n633 GND 0.32066f
C1232 VDD.n634 GND 0.004328f
C1233 VDD.n635 GND 0.004328f
C1234 VDD.n636 GND 0.004328f
C1235 VDD.n637 GND 0.004328f
C1236 VDD.n638 GND 0.004328f
C1237 VDD.n639 GND 0.32066f
C1238 VDD.n640 GND 0.004328f
C1239 VDD.n641 GND 0.004328f
C1240 VDD.n642 GND 0.004328f
C1241 VDD.n643 GND 0.004328f
C1242 VDD.n644 GND 0.004328f
C1243 VDD.t17 GND 0.32066f
C1244 VDD.n645 GND 0.004328f
C1245 VDD.n646 GND 0.004328f
C1246 VDD.n647 GND 0.004328f
C1247 VDD.n648 GND 0.004328f
C1248 VDD.n649 GND 0.004328f
C1249 VDD.n650 GND 0.32066f
C1250 VDD.n651 GND 0.004328f
C1251 VDD.n652 GND 0.004328f
C1252 VDD.n653 GND 0.004328f
C1253 VDD.n654 GND 0.004328f
C1254 VDD.n655 GND 0.004328f
C1255 VDD.n656 GND 0.32066f
C1256 VDD.n657 GND 0.004328f
C1257 VDD.n658 GND 0.004328f
C1258 VDD.n659 GND 0.004328f
C1259 VDD.n660 GND 0.004328f
C1260 VDD.n661 GND 0.004328f
C1261 VDD.n662 GND 0.32066f
C1262 VDD.n663 GND 0.004328f
C1263 VDD.n664 GND 0.004328f
C1264 VDD.n665 GND 0.004328f
C1265 VDD.n666 GND 0.004328f
C1266 VDD.n667 GND 0.004328f
C1267 VDD.n668 GND 0.32066f
C1268 VDD.n669 GND 0.004328f
C1269 VDD.n670 GND 0.004328f
C1270 VDD.n671 GND 0.004328f
C1271 VDD.n672 GND 0.004328f
C1272 VDD.n673 GND 0.004328f
C1273 VDD.n674 GND 0.24521f
C1274 VDD.n675 GND 0.004328f
C1275 VDD.n676 GND 0.004328f
C1276 VDD.n677 GND 0.004328f
C1277 VDD.n678 GND 0.004328f
C1278 VDD.n679 GND 0.004328f
C1279 VDD.t40 GND 0.16033f
C1280 VDD.n680 GND 0.004328f
C1281 VDD.n681 GND 0.004328f
C1282 VDD.t123 GND 0.16033f
C1283 VDD.n682 GND 0.004328f
C1284 VDD.n683 GND 0.004328f
C1285 VDD.n684 GND 0.004328f
C1286 VDD.n685 GND 0.32066f
C1287 VDD.n686 GND 0.004328f
C1288 VDD.n687 GND 0.004328f
C1289 VDD.n688 GND 0.264073f
C1290 VDD.n689 GND 0.004328f
C1291 VDD.n690 GND 0.004328f
C1292 VDD.n691 GND 0.004328f
C1293 VDD.n692 GND 0.32066f
C1294 VDD.n693 GND 0.004328f
C1295 VDD.n694 GND 0.004328f
C1296 VDD.n695 GND 0.004328f
C1297 VDD.n696 GND 0.009986f
C1298 VDD.n697 GND 0.009986f
C1299 VDD.n698 GND 0.417329f
C1300 VDD.n699 GND 0.004328f
C1301 VDD.n700 GND 0.004328f
C1302 VDD.n701 GND 0.009986f
C1303 VDD.n702 GND 0.004328f
C1304 VDD.n703 GND 0.004328f
C1305 VDD.t48 GND 3.17123f
C1306 VDD.n710 GND 0.010125f
C1307 VDD.n718 GND 0.010125f
C1308 VDD.n719 GND 0.004328f
C1309 VDD.n720 GND 0.004328f
C1310 VDD.n721 GND 0.004837f
C1311 VDD.n722 GND 0.004709f
C1312 VDD.n724 GND 0.005045f
C1313 VDD.n725 GND 0.005122f
C1314 VDD.n726 GND 0.006364f
C1315 VDD.t38 GND 3.64043f
C1316 VDD.t30 GND 3.64043f
C1317 VDD.t32 GND 4.31005f
C1318 VDD.t15 GND 5.46301f
C1319 VDD.n727 GND 3.33628f
C1320 VDD.t102 GND 0.123904f
C1321 VDD.t101 GND 0.415248f
C1322 VDD.n728 GND 0.086184f
C1323 VDD.t103 GND 0.090617f
C1324 VDD.n729 GND 0.088946f
C1325 VDD.n730 GND 0.009604f
C1326 VDD.n731 GND 0.006364f
C1327 VDD.n732 GND 0.006364f
C1328 VDD.n733 GND 0.005122f
C1329 VDD.n735 GND 0.006364f
C1330 VDD.n736 GND 0.006364f
C1331 VDD.n737 GND 0.006364f
C1332 VDD.n738 GND 0.006364f
C1333 VDD.n739 GND 0.006364f
C1334 VDD.n740 GND 0.005122f
C1335 VDD.n742 GND 0.006364f
C1336 VDD.n743 GND 0.006364f
C1337 VDD.n744 GND 0.006364f
C1338 VDD.n745 GND 0.006364f
C1339 VDD.n746 GND 0.006364f
C1340 VDD.n747 GND 0.005122f
C1341 VDD.n749 GND 0.006364f
C1342 VDD.n750 GND 0.006364f
C1343 VDD.n751 GND 0.006364f
C1344 VDD.n752 GND 0.006364f
C1345 VDD.n753 GND 0.006364f
C1346 VDD.n754 GND 0.005122f
C1347 VDD.n756 GND 0.006364f
C1348 VDD.n757 GND 0.006364f
C1349 VDD.n758 GND 0.006364f
C1350 VDD.n759 GND 0.006364f
C1351 VDD.n760 GND 0.006364f
C1352 VDD.n761 GND 0.005122f
C1353 VDD.n763 GND 0.006364f
C1354 VDD.n764 GND 0.006364f
C1355 VDD.n765 GND 0.006364f
C1356 VDD.n766 GND 0.006364f
C1357 VDD.n767 GND 0.006364f
C1358 VDD.n768 GND 0.005122f
C1359 VDD.n770 GND 0.006364f
C1360 VDD.n771 GND 0.006364f
C1361 VDD.n772 GND 0.006364f
C1362 VDD.n773 GND 0.006364f
C1363 VDD.n774 GND 0.006364f
C1364 VDD.n775 GND 0.002689f
C1365 VDD.n777 GND 0.006364f
C1366 VDD.t62 GND 0.123904f
C1367 VDD.t60 GND 0.415248f
C1368 VDD.n778 GND 0.086184f
C1369 VDD.t63 GND 0.090617f
C1370 VDD.n779 GND 0.088946f
C1371 VDD.n780 GND 0.007043f
C1372 VDD.n781 GND 0.006364f
C1373 VDD.n782 GND 0.006364f
C1374 VDD.n783 GND 0.004709f
C1375 VDD.n785 GND 0.006364f
C1376 VDD.n786 GND 0.005122f
C1377 VDD.n787 GND 0.004328f
C1378 VDD.n788 GND 0.004328f
C1379 VDD.n789 GND 0.004328f
C1380 VDD.n790 GND 0.004328f
C1381 VDD.n791 GND 0.004328f
C1382 VDD.n792 GND 0.004328f
C1383 VDD.n793 GND 0.004328f
C1384 VDD.n794 GND 0.004328f
C1385 VDD.n795 GND 0.004328f
C1386 VDD.n796 GND 0.004328f
C1387 VDD.n797 GND 0.004328f
C1388 VDD.n798 GND 0.003246f
C1389 VDD.t128 GND 0.066005f
C1390 VDD.t126 GND 0.213596f
C1391 VDD.n799 GND 0.071628f
C1392 VDD.t127 GND 0.048572f
C1393 VDD.n800 GND 0.068504f
C1394 VDD.n801 GND 0.004328f
C1395 VDD.n802 GND 0.004328f
C1396 VDD.n803 GND 0.004328f
C1397 VDD.n804 GND 0.004328f
C1398 VDD.n805 GND 0.004328f
C1399 VDD.n806 GND 0.004328f
C1400 VDD.n807 GND 0.004328f
C1401 VDD.n808 GND 0.004328f
C1402 VDD.n809 GND 0.004328f
C1403 VDD.n810 GND 0.004328f
C1404 VDD.n811 GND 0.004328f
C1405 VDD.n812 GND 0.004328f
C1406 VDD.n813 GND 0.004328f
C1407 VDD.n814 GND 0.004328f
C1408 VDD.n815 GND 0.004328f
C1409 VDD.n816 GND 0.004328f
C1410 VDD.n817 GND 0.004328f
C1411 VDD.n818 GND 0.004328f
C1412 VDD.n819 GND 0.004328f
C1413 VDD.n820 GND 0.004328f
C1414 VDD.n821 GND 0.004328f
C1415 VDD.n822 GND 0.004328f
C1416 VDD.n823 GND 0.004328f
C1417 VDD.n824 GND 0.004328f
C1418 VDD.n825 GND 0.004328f
C1419 VDD.n826 GND 0.004328f
C1420 VDD.n827 GND 0.004328f
C1421 VDD.n828 GND 0.004328f
C1422 VDD.n829 GND 0.004328f
C1423 VDD.n830 GND 0.004328f
C1424 VDD.n831 GND 0.004328f
C1425 VDD.n832 GND 0.004328f
C1426 VDD.n833 GND 0.004328f
C1427 VDD.n834 GND 0.004328f
C1428 VDD.n835 GND 0.004328f
C1429 VDD.n836 GND 0.004328f
C1430 VDD.n837 GND 0.004328f
C1431 VDD.n838 GND 0.004328f
C1432 VDD.n839 GND 0.004328f
C1433 VDD.n840 GND 0.004328f
C1434 VDD.n841 GND 0.004328f
C1435 VDD.n842 GND 0.004328f
C1436 VDD.n843 GND 0.004328f
C1437 VDD.n844 GND 0.004328f
C1438 VDD.n845 GND 0.004328f
C1439 VDD.n846 GND 0.004328f
C1440 VDD.n847 GND 0.004328f
C1441 VDD.n848 GND 0.004328f
C1442 VDD.n849 GND 0.004328f
C1443 VDD.n850 GND 0.004328f
C1444 VDD.n851 GND 0.004328f
C1445 VDD.n852 GND 0.004328f
C1446 VDD.n853 GND 0.004328f
C1447 VDD.n854 GND 0.004328f
C1448 VDD.n855 GND 0.004328f
C1449 VDD.n856 GND 0.004328f
C1450 VDD.n857 GND 0.004328f
C1451 VDD.n858 GND 0.004328f
C1452 VDD.n859 GND 0.004328f
C1453 VDD.n860 GND 0.004328f
C1454 VDD.n861 GND 0.004328f
C1455 VDD.n862 GND 0.004328f
C1456 VDD.n863 GND 0.004328f
C1457 VDD.n864 GND 0.004328f
C1458 VDD.n865 GND 0.004328f
C1459 VDD.n866 GND 0.009986f
C1460 VDD.n867 GND 0.009986f
C1461 VDD.n868 GND 0.010125f
C1462 VDD.n869 GND 0.004328f
C1463 VDD.n870 GND 0.004328f
C1464 VDD.n871 GND 0.004328f
C1465 VDD.n872 GND 0.004328f
C1466 VDD.n873 GND 0.004328f
C1467 VDD.n874 GND 0.002291f
C1468 VDD.n875 GND 0.00534f
C1469 VDD.n876 GND 0.0042f
C1470 VDD.n877 GND 0.004328f
C1471 VDD.n878 GND 0.004328f
C1472 VDD.n879 GND 0.004328f
C1473 VDD.n880 GND 0.004328f
C1474 VDD.n881 GND 0.004328f
C1475 VDD.n882 GND 0.004328f
C1476 VDD.n883 GND 0.003246f
C1477 VDD.n884 GND 0.12184f
C1478 VDD.n886 GND 0.006364f
C1479 VDD.n887 GND 0.005122f
C1480 VDD.n888 GND 0.006364f
C1481 VDD.n890 GND 0.005122f
C1482 VDD.n891 GND 0.006364f
C1483 VDD.n892 GND 0.006364f
C1484 VDD.n894 GND 0.006364f
C1485 VDD.n895 GND 0.006364f
C1486 VDD.n897 GND 0.006364f
C1487 VDD.n898 GND 0.005122f
C1488 VDD.n899 GND 0.006364f
C1489 VDD.n900 GND 0.006364f
C1490 VDD.n902 GND 0.006364f
C1491 VDD.n903 GND 0.006364f
C1492 VDD.n905 GND 0.006364f
C1493 VDD.n906 GND 0.002792f
C1494 VDD.n907 GND 0.014395f
C1495 VDD.t72 GND 0.123904f
C1496 VDD.t71 GND 0.415248f
C1497 VDD.n908 GND 0.086184f
C1498 VDD.t73 GND 0.090617f
C1499 VDD.n909 GND 0.088946f
C1500 VDD.n910 GND 0.007043f
C1501 VDD.n911 GND 0.006364f
C1502 VDD.n913 GND 0.006364f
C1503 VDD.n914 GND 0.004251f
C1504 VDD.n915 GND 0.471559f
C1505 VDD.n916 GND 0.006364f
C1506 VDD.n917 GND 0.01437f
C1507 VDD.n918 GND 0.005122f
C1508 VDD.n919 GND 0.006364f
C1509 VDD.n920 GND 0.005122f
C1510 VDD.n921 GND 0.006364f
C1511 VDD.n922 GND 0.471559f
C1512 VDD.n923 GND 0.006364f
C1513 VDD.n924 GND 0.005122f
C1514 VDD.n925 GND 0.005122f
C1515 VDD.n926 GND 0.006364f
C1516 VDD.n927 GND 0.005122f
C1517 VDD.n928 GND 0.006364f
C1518 VDD.n929 GND 0.282935f
C1519 VDD.n930 GND 0.006364f
C1520 VDD.n931 GND 0.005122f
C1521 VDD.n932 GND 0.006364f
C1522 VDD.n933 GND 0.005122f
C1523 VDD.n934 GND 0.006364f
C1524 VDD.n935 GND 0.471559f
C1525 VDD.n936 GND 0.006364f
C1526 VDD.n937 GND 0.005122f
C1527 VDD.n938 GND 0.006364f
C1528 VDD.n939 GND 0.005122f
C1529 VDD.n940 GND 0.006364f
C1530 VDD.n941 GND 0.471559f
C1531 VDD.n942 GND 0.006364f
C1532 VDD.n943 GND 0.005122f
C1533 VDD.n944 GND 0.006364f
C1534 VDD.n945 GND 0.005122f
C1535 VDD.n946 GND 0.006364f
C1536 VDD.n947 GND 0.471559f
C1537 VDD.n948 GND 0.006364f
C1538 VDD.n949 GND 0.005122f
C1539 VDD.n950 GND 0.006364f
C1540 VDD.n951 GND 0.005122f
C1541 VDD.n952 GND 0.006364f
C1542 VDD.n953 GND 0.471559f
C1543 VDD.n954 GND 0.006364f
C1544 VDD.n955 GND 0.005122f
C1545 VDD.n956 GND 0.006364f
C1546 VDD.n957 GND 0.005122f
C1547 VDD.n958 GND 0.006364f
C1548 VDD.n959 GND 0.471559f
C1549 VDD.n960 GND 0.006364f
C1550 VDD.n961 GND 0.005122f
C1551 VDD.n962 GND 0.006364f
C1552 VDD.n963 GND 0.005122f
C1553 VDD.n964 GND 0.006364f
C1554 VDD.n965 GND 0.240495f
C1555 VDD.n966 GND 0.006364f
C1556 VDD.n967 GND 0.005122f
C1557 VDD.n968 GND 0.006364f
C1558 VDD.n969 GND 0.005122f
C1559 VDD.n970 GND 0.006364f
C1560 VDD.n971 GND 0.471559f
C1561 VDD.n972 GND 0.006364f
C1562 VDD.n973 GND 0.005122f
C1563 VDD.n974 GND 0.006364f
C1564 VDD.n975 GND 0.005122f
C1565 VDD.n976 GND 0.006364f
C1566 VDD.n977 GND 0.471559f
C1567 VDD.n978 GND 0.006364f
C1568 VDD.n979 GND 0.005122f
C1569 VDD.n980 GND 0.006364f
C1570 VDD.n981 GND 0.005122f
C1571 VDD.n982 GND 0.006364f
C1572 VDD.n983 GND 0.471559f
C1573 VDD.n984 GND 0.006364f
C1574 VDD.n985 GND 0.005122f
C1575 VDD.n986 GND 0.006364f
C1576 VDD.n987 GND 0.005122f
C1577 VDD.n988 GND 0.006364f
C1578 VDD.n989 GND 0.471559f
C1579 VDD.n990 GND 0.006364f
C1580 VDD.n991 GND 0.005122f
C1581 VDD.n992 GND 0.006342f
C1582 VDD.n993 GND 0.005122f
C1583 VDD.n994 GND 0.006364f
C1584 VDD.n995 GND 0.471559f
C1585 VDD.n996 GND 0.006364f
C1586 VDD.n997 GND 0.005122f
C1587 VDD.n998 GND 0.006364f
C1588 VDD.n999 GND 0.005122f
C1589 VDD.n1000 GND 0.006364f
C1590 VDD.n1001 GND 0.471559f
C1591 VDD.n1002 GND 0.006364f
C1592 VDD.n1003 GND 0.005122f
C1593 VDD.n1004 GND 0.006364f
C1594 VDD.n1005 GND 0.005122f
C1595 VDD.n1006 GND 0.006364f
C1596 VDD.n1007 GND 0.471559f
C1597 VDD.n1008 GND 0.006364f
C1598 VDD.n1009 GND 0.005122f
C1599 VDD.n1010 GND 0.006364f
C1600 VDD.n1011 GND 0.005122f
C1601 VDD.n1012 GND 0.006364f
C1602 VDD.n1013 GND 0.471559f
C1603 VDD.n1014 GND 0.006364f
C1604 VDD.n1015 GND 0.005122f
C1605 VDD.n1016 GND 0.006364f
C1606 VDD.n1017 GND 0.005122f
C1607 VDD.n1018 GND 0.006364f
C1608 VDD.t4 GND 0.235779f
C1609 VDD.n1019 GND 0.006364f
C1610 VDD.n1020 GND 0.005122f
C1611 VDD.n1021 GND 0.006364f
C1612 VDD.n1022 GND 0.005122f
C1613 VDD.n1023 GND 0.006364f
C1614 VDD.n1024 GND 0.471559f
C1615 VDD.n1025 GND 0.240495f
C1616 VDD.n1026 GND 0.006364f
C1617 VDD.n1027 GND 0.005122f
C1618 VDD.n1028 GND 0.006364f
C1619 VDD.n1029 GND 0.005122f
C1620 VDD.n1030 GND 0.006364f
C1621 VDD.n1031 GND 0.471559f
C1622 VDD.n1032 GND 0.006364f
C1623 VDD.n1033 GND 0.005122f
C1624 VDD.n1034 GND 0.006364f
C1625 VDD.n1035 GND 0.005122f
C1626 VDD.n1036 GND 0.006364f
C1627 VDD.n1037 GND 0.471559f
C1628 VDD.n1038 GND 0.006364f
C1629 VDD.n1039 GND 0.005122f
C1630 VDD.n1040 GND 0.006364f
C1631 VDD.n1041 GND 0.005122f
C1632 VDD.n1042 GND 0.006364f
C1633 VDD.n1043 GND 0.471559f
C1634 VDD.n1044 GND 0.006364f
C1635 VDD.n1045 GND 0.005122f
C1636 VDD.n1046 GND 0.006364f
C1637 VDD.n1047 GND 0.005122f
C1638 VDD.n1048 GND 0.006364f
C1639 VDD.n1049 GND 0.471559f
C1640 VDD.n1050 GND 0.006364f
C1641 VDD.n1051 GND 0.005122f
C1642 VDD.n1052 GND 0.006364f
C1643 VDD.n1053 GND 0.005122f
C1644 VDD.n1054 GND 0.006364f
C1645 VDD.t68 GND 0.235779f
C1646 VDD.n1055 GND 0.006364f
C1647 VDD.n1056 GND 0.005122f
C1648 VDD.n1057 GND 0.006364f
C1649 VDD.n1058 GND 0.005122f
C1650 VDD.n1059 GND 0.006364f
C1651 VDD.n1060 GND 0.471559f
C1652 VDD.n1061 GND 0.282935f
C1653 VDD.n1062 GND 0.006364f
C1654 VDD.n1063 GND 0.005122f
C1655 VDD.n1064 GND 0.006364f
C1656 VDD.n1065 GND 0.005122f
C1657 VDD.n1066 GND 0.006364f
C1658 VDD.n1067 GND 0.471559f
C1659 VDD.n1068 GND 0.006364f
C1660 VDD.n1069 GND 0.005122f
C1661 VDD.n1070 GND 0.01437f
C1662 VDD.n1071 GND 0.01437f
C1663 VDD.n1072 GND 1.01857f
C1664 VDD.n1073 GND 0.01437f
C1665 VDD.n1074 GND 0.006364f
C1666 VDD.n1076 GND 0.006364f
C1667 VDD.n1077 GND 0.006364f
C1668 VDD.n1078 GND 0.005122f
C1669 VDD.n1079 GND 0.006364f
C1670 VDD.n1080 GND 0.006364f
C1671 VDD.n1082 GND 0.006364f
C1672 VDD.n1083 GND 0.006364f
C1673 VDD.n1085 GND 0.006364f
C1674 VDD.n1086 GND 0.005122f
C1675 VDD.n1087 GND 0.006364f
C1676 VDD.n1088 GND 0.006364f
C1677 VDD.n1090 GND 0.006364f
C1678 VDD.n1091 GND 0.006364f
C1679 VDD.n1093 GND 0.006364f
C1680 VDD.t70 GND 0.123904f
C1681 VDD.t67 GND 0.415248f
C1682 VDD.n1094 GND 0.086184f
C1683 VDD.t69 GND 0.090617f
C1684 VDD.n1095 GND 0.088946f
C1685 VDD.n1096 GND 0.009604f
C1686 VDD.n1097 GND 0.006364f
C1687 VDD.n1098 GND 0.006364f
C1688 VDD.n1100 GND 0.006364f
C1689 VDD.n1101 GND 0.006364f
C1690 VDD.n1103 GND 0.006364f
C1691 VDD.n1104 GND 0.005122f
C1692 VDD.n1105 GND 0.006364f
C1693 VDD.n1106 GND 0.006364f
C1694 VDD.n1108 GND 0.006364f
C1695 VDD.n1109 GND 0.006364f
C1696 VDD.n1111 GND 0.006364f
C1697 VDD.n1112 GND 0.005122f
C1698 VDD.n1113 GND 0.006364f
C1699 VDD.n1114 GND 0.006364f
C1700 VDD.n1116 GND 0.006364f
C1701 VDD.n1117 GND 0.006364f
C1702 VDD.n1119 GND 0.006364f
C1703 VDD.n1120 GND 0.005122f
C1704 VDD.n1121 GND 0.006364f
C1705 VDD.n1122 GND 0.006364f
C1706 VDD.n1124 GND 0.006364f
C1707 VDD.n1125 GND 0.006364f
C1708 VDD.n1127 GND 0.006364f
C1709 VDD.n1128 GND 0.005122f
C1710 VDD.n1129 GND 0.006364f
C1711 VDD.n1130 GND 0.006364f
C1712 VDD.n1132 GND 0.006364f
C1713 VDD.n1133 GND 0.006364f
C1714 VDD.n1135 GND 0.006364f
C1715 VDD.n1136 GND 0.005122f
C1716 VDD.n1137 GND 0.006364f
C1717 VDD.n1138 GND 0.006364f
C1718 VDD.n1140 GND 0.006364f
C1719 VDD.n1141 GND 0.006364f
C1720 VDD.n1143 GND 0.006364f
C1721 VDD.n1144 GND 0.005122f
C1722 VDD.n1145 GND 0.006364f
C1723 VDD.n1146 GND 0.006364f
C1724 VDD.n1148 GND 0.006364f
C1725 VDD.n1149 GND 0.006364f
C1726 VDD.n1151 GND 0.006364f
C1727 VDD.n1152 GND 0.002689f
C1728 VDD.n1153 GND 0.006364f
C1729 VDD.t97 GND 0.123904f
C1730 VDD.t95 GND 0.415248f
C1731 VDD.n1154 GND 0.086184f
C1732 VDD.t96 GND 0.090617f
C1733 VDD.n1155 GND 0.088946f
C1734 VDD.n1156 GND 0.007043f
C1735 VDD.n1157 GND 0.006364f
C1736 VDD.n1159 GND 0.006364f
C1737 VDD.n1160 GND 0.006364f
C1738 VDD.n1162 GND 0.006364f
C1739 VDD.n1163 GND 0.005122f
C1740 VDD.n1164 GND 0.006364f
C1741 VDD.n1165 GND 0.006364f
C1742 VDD.n1167 GND 0.006364f
C1743 VDD.n1168 GND 0.006364f
C1744 VDD.n1170 GND 0.006364f
C1745 VDD.n1171 GND 0.005122f
C1746 VDD.n1172 GND 0.006364f
C1747 VDD.n1173 GND 0.006364f
C1748 VDD.n1175 GND 0.006364f
C1749 VDD.n1176 GND 0.006364f
C1750 VDD.n1178 GND 0.006364f
C1751 VDD.n1179 GND 0.005122f
C1752 VDD.n1180 GND 0.006364f
C1753 VDD.n1181 GND 0.006364f
C1754 VDD.n1183 GND 0.006364f
C1755 VDD.n1185 GND 0.006364f
C1756 VDD.n1186 GND 0.002331f
C1757 VDD.t106 GND 0.123904f
C1758 VDD.t104 GND 0.415248f
C1759 VDD.n1187 GND 0.086184f
C1760 VDD.t105 GND 0.090617f
C1761 VDD.n1188 GND 0.088946f
C1762 VDD.n1189 GND 0.007043f
C1763 VDD.n1190 GND 0.002792f
C1764 VDD.n1191 GND 0.005122f
C1765 VDD.n1192 GND 0.006364f
C1766 VDD.n1193 GND 0.006364f
C1767 VDD.n1194 GND 0.006364f
C1768 VDD.n1195 GND 0.005122f
C1769 VDD.n1196 GND 0.005122f
C1770 VDD.n1197 GND 0.005122f
C1771 VDD.n1198 GND 0.006364f
C1772 VDD.n1199 GND 0.006364f
C1773 VDD.n1200 GND 0.006364f
C1774 VDD.n1201 GND 0.005122f
C1775 VDD.n1202 GND 0.005122f
C1776 VDD.n1203 GND 0.005122f
C1777 VDD.n1204 GND 0.006364f
C1778 VDD.n1205 GND 0.006364f
C1779 VDD.n1206 GND 0.006364f
C1780 VDD.n1207 GND 0.005122f
C1781 VDD.n1208 GND 0.005122f
C1782 VDD.n1209 GND 0.003304f
C1783 VDD.n1210 GND 0.006364f
C1784 VDD.n1211 GND 0.006364f
C1785 VDD.n1212 GND 0.006364f
C1786 VDD.n1213 GND 0.005122f
C1787 VDD.n1214 GND 0.005122f
C1788 VDD.n1215 GND 0.005122f
C1789 VDD.n1216 GND 0.006364f
C1790 VDD.n1217 GND 0.006364f
C1791 VDD.n1218 GND 0.006364f
C1792 VDD.n1219 GND 0.005122f
C1793 VDD.n1220 GND 0.005122f
C1794 VDD.n1221 GND 0.005122f
C1795 VDD.n1222 GND 0.006364f
C1796 VDD.n1223 GND 0.006364f
C1797 VDD.n1224 GND 0.006364f
C1798 VDD.n1225 GND 0.005122f
C1799 VDD.n1226 GND 0.005122f
C1800 VDD.n1227 GND 0.005122f
C1801 VDD.n1228 GND 0.006364f
C1802 VDD.n1229 GND 0.006364f
C1803 VDD.n1230 GND 0.006364f
C1804 VDD.n1231 GND 0.003406f
C1805 VDD.t91 GND 0.123904f
C1806 VDD.t89 GND 0.415248f
C1807 VDD.n1232 GND 0.086184f
C1808 VDD.t90 GND 0.090617f
C1809 VDD.n1233 GND 0.088946f
C1810 VDD.n1234 GND 0.007043f
C1811 VDD.n1235 GND 0.002587f
C1812 VDD.n1236 GND 0.005122f
C1813 VDD.n1237 GND 0.006364f
C1814 VDD.n1238 GND 0.006364f
C1815 VDD.n1239 GND 0.006364f
C1816 VDD.n1240 GND 0.005122f
C1817 VDD.n1241 GND 0.005122f
C1818 VDD.n1242 GND 0.005122f
C1819 VDD.n1243 GND 0.006364f
C1820 VDD.n1244 GND 0.006364f
C1821 VDD.n1245 GND 0.006364f
C1822 VDD.n1246 GND 0.005122f
C1823 VDD.n1247 GND 0.005122f
C1824 VDD.n1248 GND 0.005122f
C1825 VDD.n1249 GND 0.006364f
C1826 VDD.n1250 GND 0.006364f
C1827 VDD.n1251 GND 0.006364f
C1828 VDD.n1252 GND 0.005122f
C1829 VDD.n1253 GND 0.005122f
C1830 VDD.n1254 GND 0.003509f
C1831 VDD.n1255 GND 0.006364f
C1832 VDD.n1256 GND 0.006364f
C1833 VDD.n1257 GND 0.006364f
C1834 VDD.n1258 GND 0.005045f
C1835 VDD.n1259 GND 0.005122f
C1836 VDD.n1260 GND 0.005122f
C1837 VDD.n1261 GND 0.006364f
C1838 VDD.n1262 GND 0.006364f
C1839 VDD.n1263 GND 0.006364f
C1840 VDD.n1264 GND 0.005122f
C1841 VDD.n1265 GND 0.005122f
C1842 VDD.n1266 GND 0.005122f
C1843 VDD.n1267 GND 0.006364f
C1844 VDD.n1268 GND 0.006364f
C1845 VDD.n1269 GND 0.006364f
C1846 VDD.n1270 GND 0.005122f
C1847 VDD.n1271 GND 0.005122f
C1848 VDD.n1272 GND 0.004251f
C1849 VDD.n1273 GND 0.01437f
C1850 VDD.n1274 GND 0.014395f
C1851 VDD.n1275 GND 0.004251f
C1852 VDD.n1276 GND 0.014395f
C1853 VDD.n1277 GND 0.598879f
C1854 VDD.n1278 GND 0.014395f
C1855 VDD.n1279 GND 0.004251f
C1856 VDD.n1280 GND 0.014395f
C1857 VDD.n1281 GND 0.006364f
C1858 VDD.n1282 GND 0.006364f
C1859 VDD.n1283 GND 0.005122f
C1860 VDD.n1284 GND 0.006364f
C1861 VDD.n1285 GND 0.471559f
C1862 VDD.n1286 GND 0.006364f
C1863 VDD.n1287 GND 0.005122f
C1864 VDD.n1288 GND 0.006364f
C1865 VDD.n1289 GND 0.006364f
C1866 VDD.n1290 GND 0.006364f
C1867 VDD.n1291 GND 0.005122f
C1868 VDD.n1292 GND 0.006364f
C1869 VDD.n1293 GND 0.471559f
C1870 VDD.n1294 GND 0.006364f
C1871 VDD.n1295 GND 0.005122f
C1872 VDD.n1296 GND 0.006364f
C1873 VDD.n1297 GND 0.006364f
C1874 VDD.n1298 GND 0.006364f
C1875 VDD.n1299 GND 0.005122f
C1876 VDD.n1300 GND 0.006364f
C1877 VDD.n1301 GND 0.424403f
C1878 VDD.n1302 GND 0.006364f
C1879 VDD.n1303 GND 0.005122f
C1880 VDD.n1304 GND 0.006364f
C1881 VDD.n1305 GND 0.006364f
C1882 VDD.n1306 GND 0.006364f
C1883 VDD.n1307 GND 0.005122f
C1884 VDD.n1308 GND 0.006364f
C1885 VDD.n1309 GND 0.471559f
C1886 VDD.n1310 GND 0.006364f
C1887 VDD.n1311 GND 0.005122f
C1888 VDD.n1312 GND 0.006364f
C1889 VDD.n1313 GND 0.006364f
C1890 VDD.n1314 GND 0.006364f
C1891 VDD.n1315 GND 0.005122f
C1892 VDD.n1316 GND 0.006364f
C1893 VDD.n1317 GND 0.471559f
C1894 VDD.n1318 GND 0.006364f
C1895 VDD.n1319 GND 0.005122f
C1896 VDD.n1320 GND 0.006364f
C1897 VDD.n1321 GND 0.006364f
C1898 VDD.n1322 GND 0.006364f
C1899 VDD.n1323 GND 0.005122f
C1900 VDD.n1324 GND 0.006364f
C1901 VDD.n1325 GND 0.471559f
C1902 VDD.n1326 GND 0.006364f
C1903 VDD.n1327 GND 0.005122f
C1904 VDD.n1328 GND 0.006364f
C1905 VDD.n1329 GND 0.006364f
C1906 VDD.n1330 GND 0.006364f
C1907 VDD.n1331 GND 0.005122f
C1908 VDD.n1332 GND 0.006364f
C1909 VDD.n1333 GND 0.471559f
C1910 VDD.n1334 GND 0.006364f
C1911 VDD.n1335 GND 0.005122f
C1912 VDD.n1336 GND 0.006364f
C1913 VDD.n1337 GND 0.006364f
C1914 VDD.n1338 GND 0.006364f
C1915 VDD.n1339 GND 0.005122f
C1916 VDD.n1340 GND 0.006364f
C1917 VDD.n1341 GND 0.471559f
C1918 VDD.n1342 GND 0.006364f
C1919 VDD.n1343 GND 0.005122f
C1920 VDD.n1344 GND 0.006364f
C1921 VDD.n1345 GND 0.006364f
C1922 VDD.n1346 GND 0.006364f
C1923 VDD.n1347 GND 0.005122f
C1924 VDD.n1348 GND 0.006364f
C1925 VDD.n1349 GND 0.466843f
C1926 VDD.n1350 GND 0.006364f
C1927 VDD.n1351 GND 0.005122f
C1928 VDD.n1352 GND 0.006364f
C1929 VDD.n1353 GND 0.006364f
C1930 VDD.n1354 GND 0.006364f
C1931 VDD.n1355 GND 0.005122f
C1932 VDD.n1356 GND 0.006364f
C1933 VDD.n1357 GND 0.471559f
C1934 VDD.n1358 GND 0.006364f
C1935 VDD.n1359 GND 0.005122f
C1936 VDD.n1360 GND 0.006364f
C1937 VDD.n1361 GND 0.006364f
C1938 VDD.n1362 GND 0.006364f
C1939 VDD.n1363 GND 0.005122f
C1940 VDD.n1364 GND 0.006364f
C1941 VDD.n1365 GND 0.471559f
C1942 VDD.n1366 GND 0.006364f
C1943 VDD.n1367 GND 0.005122f
C1944 VDD.n1368 GND 0.006364f
C1945 VDD.n1369 GND 0.006364f
C1946 VDD.n1370 GND 0.006364f
C1947 VDD.n1371 GND 0.005122f
C1948 VDD.n1372 GND 0.006364f
C1949 VDD.n1373 GND 0.471559f
C1950 VDD.n1374 GND 0.006364f
C1951 VDD.n1375 GND 0.005122f
C1952 VDD.n1376 GND 0.006364f
C1953 VDD.n1377 GND 0.006364f
C1954 VDD.n1378 GND 0.006364f
C1955 VDD.n1379 GND 0.005122f
C1956 VDD.n1380 GND 0.006364f
C1957 VDD.t12 GND 0.471559f
C1958 VDD.n1381 GND 0.006364f
C1959 VDD.n1382 GND 0.005122f
C1960 VDD.t9 GND 0.103757f
C1961 VDD.t132 GND 0.018389f
C1962 VDD.t13 GND 0.018389f
C1963 VDD.n1383 GND 0.073262f
C1964 VDD.n1384 GND 0.584701f
C1965 VDD.t8 GND 0.103757f
C1966 VDD.t5 GND 0.018389f
C1967 VDD.t144 GND 0.018389f
C1968 VDD.n1385 GND 0.073262f
C1969 VDD.n1386 GND 0.566686f
C1970 VDD.n1387 GND 0.295728f
C1971 VDD.t136 GND 0.103757f
C1972 VDD.t135 GND 0.018389f
C1973 VDD.t50 GND 0.018389f
C1974 VDD.n1388 GND 0.073262f
C1975 VDD.n1389 GND 0.566686f
C1976 VDD.n1390 GND 0.201367f
C1977 VDD.t143 GND 0.103757f
C1978 VDD.t14 GND 0.018389f
C1979 VDD.t134 GND 0.018389f
C1980 VDD.n1391 GND 0.073262f
C1981 VDD.n1392 GND 0.566686f
C1982 VDD.n1393 GND 0.27854f
C1983 VDD.n1394 GND 1.89347f
C1984 VDD.n1395 GND 0.14125f
C1985 VDD.n1396 GND 0.006342f
C1986 VDD.n1397 GND 0.006364f
C1987 VDD.n1398 GND 0.005122f
C1988 VDD.n1399 GND 0.006364f
C1989 VDD.n1400 GND 0.471559f
C1990 VDD.n1401 GND 0.006364f
C1991 VDD.n1402 GND 0.005122f
C1992 VDD.n1403 GND 0.006364f
C1993 VDD.n1404 GND 0.006364f
C1994 VDD.n1405 GND 0.006364f
C1995 VDD.n1406 GND 0.005122f
C1996 VDD.n1407 GND 0.006364f
C1997 VDD.n1408 GND 0.471559f
C1998 VDD.n1409 GND 0.006364f
C1999 VDD.n1410 GND 0.005122f
C2000 VDD.n1411 GND 0.006364f
C2001 VDD.n1412 GND 0.006364f
C2002 VDD.n1413 GND 0.006364f
C2003 VDD.n1414 GND 0.005122f
C2004 VDD.n1415 GND 0.006364f
C2005 VDD.n1416 GND 0.471559f
C2006 VDD.n1417 GND 0.006364f
C2007 VDD.n1418 GND 0.005122f
C2008 VDD.n1419 GND 0.006364f
C2009 VDD.n1420 GND 0.006364f
C2010 VDD.n1421 GND 0.006364f
C2011 VDD.n1422 GND 0.005122f
C2012 VDD.n1423 GND 0.006364f
C2013 VDD.t7 GND 0.235779f
C2014 VDD.n1424 GND 0.466843f
C2015 VDD.n1425 GND 0.006364f
C2016 VDD.n1426 GND 0.005122f
C2017 VDD.n1427 GND 0.006364f
C2018 VDD.n1428 GND 0.006364f
C2019 VDD.n1429 GND 0.006364f
C2020 VDD.n1430 GND 0.005122f
C2021 VDD.n1431 GND 0.006364f
C2022 VDD.n1432 GND 0.471559f
C2023 VDD.n1433 GND 0.006364f
C2024 VDD.n1434 GND 0.005122f
C2025 VDD.n1435 GND 0.006364f
C2026 VDD.n1436 GND 0.006364f
C2027 VDD.n1437 GND 0.006364f
C2028 VDD.n1438 GND 0.005122f
C2029 VDD.n1439 GND 0.006364f
C2030 VDD.n1440 GND 0.471559f
C2031 VDD.n1441 GND 0.006364f
C2032 VDD.n1442 GND 0.005122f
C2033 VDD.n1443 GND 0.006364f
C2034 VDD.n1444 GND 0.006364f
C2035 VDD.n1445 GND 0.006364f
C2036 VDD.n1446 GND 0.005122f
C2037 VDD.n1447 GND 0.006364f
C2038 VDD.n1448 GND 0.471559f
C2039 VDD.n1449 GND 0.006364f
C2040 VDD.n1450 GND 0.005122f
C2041 VDD.n1451 GND 0.006364f
C2042 VDD.n1452 GND 0.006364f
C2043 VDD.n1453 GND 0.006364f
C2044 VDD.n1454 GND 0.005122f
C2045 VDD.n1455 GND 0.006364f
C2046 VDD.n1456 GND 0.471559f
C2047 VDD.n1457 GND 0.006364f
C2048 VDD.n1458 GND 0.005122f
C2049 VDD.n1459 GND 0.006364f
C2050 VDD.n1460 GND 0.006364f
C2051 VDD.n1461 GND 0.006364f
C2052 VDD.n1462 GND 0.005122f
C2053 VDD.n1463 GND 0.006364f
C2054 VDD.n1464 GND 0.471559f
C2055 VDD.n1465 GND 0.006364f
C2056 VDD.n1466 GND 0.005122f
C2057 VDD.n1467 GND 0.006364f
C2058 VDD.n1468 GND 0.006364f
C2059 VDD.n1469 GND 0.006364f
C2060 VDD.n1470 GND 0.005122f
C2061 VDD.n1471 GND 0.006364f
C2062 VDD.t61 GND 0.235779f
C2063 VDD.n1472 GND 0.424403f
C2064 VDD.n1473 GND 0.006364f
C2065 VDD.n1474 GND 0.005122f
C2066 VDD.n1475 GND 0.006364f
C2067 VDD.n1476 GND 0.006364f
C2068 VDD.n1477 GND 0.006364f
C2069 VDD.n1478 GND 0.005122f
C2070 VDD.n1479 GND 0.006364f
C2071 VDD.n1480 GND 0.471559f
C2072 VDD.n1481 GND 0.006364f
C2073 VDD.n1482 GND 0.005122f
C2074 VDD.n1483 GND 0.006364f
C2075 VDD.n1484 GND 0.006364f
C2076 VDD.n1485 GND 0.006364f
C2077 VDD.n1486 GND 0.006364f
C2078 VDD.n1487 GND 0.005122f
C2079 VDD.n1488 GND 0.006364f
C2080 VDD.n1489 GND 0.471559f
C2081 VDD.n1490 GND 0.006364f
C2082 VDD.n1491 GND 0.005122f
C2083 VDD.n1492 GND 0.006364f
C2084 VDD.n1493 GND 0.006364f
C2085 VDD.n1494 GND 0.006364f
C2086 VDD.n1495 GND 0.005122f
C2087 VDD.n1496 GND 0.005122f
C2088 VDD.n1497 GND 0.006364f
C2089 VDD.n1498 GND 0.006364f
C2090 VDD.n1499 GND 0.006364f
C2091 VDD.n1500 GND 0.006364f
C2092 VDD.n1501 GND 0.006364f
C2093 VDD.n1502 GND 0.006364f
C2094 VDD.n1503 GND 0.006364f
C2095 VDD.n1504 GND 0.005122f
C2096 VDD.n1507 GND 0.006364f
C2097 VDD.n1508 GND 0.006364f
C2098 VDD.n1509 GND 0.005122f
C2099 VDD.n1510 GND 0.005122f
C2100 VDD.n1511 GND 0.005122f
C2101 VDD.n1512 GND 0.006364f
C2102 VDD.n1514 GND 0.006364f
C2103 VDD.n1515 GND 0.006364f
C2104 VDD.n1517 GND 0.006364f
C2105 VDD.n1518 GND 0.005122f
C2106 VDD.n1519 GND 0.004251f
C2107 VDD.n1520 GND 0.01437f
C2108 VDD.n1521 GND 0.014395f
C2109 VDD.n1522 GND 0.004251f
C2110 VDD.n1523 GND 0.014395f
C2111 VDD.n1524 GND 0.598879f
C2112 VDD.n1525 GND 0.014395f
C2113 VDD.n1526 GND 0.01437f
C2114 VDD.n1527 GND 0.002331f
C2115 VDD.n1528 GND 0.01437f
C2116 VDD.n1529 GND 0.006364f
C2117 VDD.n1530 GND 0.006364f
C2118 VDD.n1531 GND 0.005122f
C2119 VDD.n1532 GND 0.005122f
C2120 VDD.n1533 GND 0.005122f
C2121 VDD.n1534 GND 0.006364f
C2122 VDD.n1535 GND 0.006364f
C2123 VDD.n1536 GND 0.006364f
C2124 VDD.n1537 GND 0.005122f
C2125 VDD.n1538 GND 0.005122f
C2126 VDD.n1539 GND 0.005122f
C2127 VDD.n1540 GND 0.004837f
C2128 VDD.n1541 GND 1.49966f
C2129 VDD.n1543 GND 0.005122f
C2130 VDD.n1544 GND 0.005122f
C2131 VDD.n1545 GND 0.003304f
C2132 VDD.n1546 GND 0.006364f
C2133 VDD.n1548 GND 0.006364f
C2134 VDD.n1549 GND 0.006364f
C2135 VDD.n1550 GND 0.005122f
C2136 VDD.n1551 GND 0.005122f
C2137 VDD.n1552 GND 0.005122f
C2138 VDD.n1553 GND 0.006364f
C2139 VDD.n1555 GND 0.006364f
C2140 VDD.n1556 GND 0.006364f
C2141 VDD.n1557 GND 0.005122f
C2142 VDD.n1558 GND 0.005122f
C2143 VDD.n1559 GND 0.005122f
C2144 VDD.n1560 GND 0.006364f
C2145 VDD.n1562 GND 0.006364f
C2146 VDD.n1563 GND 0.006364f
C2147 VDD.n1564 GND 0.005122f
C2148 VDD.n1565 GND 0.005122f
C2149 VDD.n1566 GND 0.005122f
C2150 VDD.n1567 GND 0.006364f
C2151 VDD.n1569 GND 0.006364f
C2152 VDD.n1570 GND 0.006364f
C2153 VDD.n1571 GND 0.003406f
C2154 VDD.t65 GND 0.123904f
C2155 VDD.t64 GND 0.415248f
C2156 VDD.n1572 GND 0.086184f
C2157 VDD.t66 GND 0.090617f
C2158 VDD.n1573 GND 0.088946f
C2159 VDD.n1574 GND 0.007043f
C2160 VDD.n1575 GND 0.002587f
C2161 VDD.n1576 GND 0.005122f
C2162 VDD.n1577 GND 0.006364f
C2163 VDD.n1579 GND 0.006364f
C2164 VDD.n1580 GND 0.006364f
C2165 VDD.n1581 GND 0.005122f
C2166 VDD.n1582 GND 0.005122f
C2167 VDD.n1583 GND 0.005122f
C2168 VDD.n1584 GND 0.006364f
C2169 VDD.n1586 GND 0.006364f
C2170 VDD.n1587 GND 0.006364f
C2171 VDD.n1588 GND 0.005122f
C2172 VDD.n1589 GND 0.005122f
C2173 VDD.n1590 GND 0.005122f
C2174 VDD.n1591 GND 0.006364f
C2175 VDD.n1593 GND 0.006364f
C2176 VDD.n1594 GND 0.006364f
C2177 VDD.n1595 GND 0.005122f
C2178 VDD.n1596 GND 0.005122f
C2179 VDD.n1597 GND 0.003509f
C2180 VDD.n1598 GND 0.006364f
C2181 VDD.n1600 GND 0.006364f
C2182 VDD.n1601 GND 0.006364f
C2183 VDD.n1603 GND 0.006364f
C2184 VDD.n1604 GND 0.005122f
C2185 VDD.n1606 GND 1.49966f
C2186 VDD.t125 GND 0.066005f
C2187 VDD.t122 GND 0.213596f
C2188 VDD.n1607 GND 0.071628f
C2189 VDD.t124 GND 0.048572f
C2190 VDD.n1608 GND 0.068504f
C2191 VDD.n1609 GND 0.004328f
C2192 VDD.n1610 GND 0.004328f
C2193 VDD.n1611 GND 0.004328f
C2194 VDD.n1612 GND 0.004328f
C2195 VDD.n1613 GND 0.004328f
C2196 VDD.n1614 GND 0.004328f
C2197 VDD.n1615 GND 0.004328f
C2198 VDD.n1616 GND 0.004328f
C2199 VDD.n1617 GND 0.004328f
C2200 VDD.n1618 GND 0.004328f
C2201 VDD.n1619 GND 0.004328f
C2202 VDD.n1620 GND 0.004328f
C2203 VDD.n1621 GND 0.004328f
C2204 VDD.n1622 GND 0.004328f
C2205 VDD.n1623 GND 0.004328f
C2206 VDD.n1624 GND 0.004328f
C2207 VDD.n1625 GND 0.004328f
C2208 VDD.n1626 GND 0.004328f
C2209 VDD.n1627 GND 0.004328f
C2210 VDD.n1628 GND 0.004328f
C2211 VDD.n1629 GND 0.004328f
C2212 VDD.n1630 GND 0.004328f
C2213 VDD.n1631 GND 0.004328f
C2214 VDD.n1632 GND 0.004328f
C2215 VDD.n1633 GND 0.004328f
C2216 VDD.n1634 GND 0.004328f
C2217 VDD.n1635 GND 0.004328f
C2218 VDD.n1636 GND 0.004328f
C2219 VDD.n1637 GND 0.004328f
C2220 VDD.n1638 GND 0.004328f
C2221 VDD.n1639 GND 0.004328f
C2222 VDD.n1640 GND 0.004328f
C2223 VDD.n1641 GND 0.004328f
C2224 VDD.n1642 GND 0.004328f
C2225 VDD.n1643 GND 0.004328f
C2226 VDD.n1644 GND 0.004328f
C2227 VDD.n1645 GND 0.004328f
C2228 VDD.n1646 GND 0.004328f
C2229 VDD.n1647 GND 0.004328f
C2230 VDD.n1648 GND 0.004328f
C2231 VDD.n1649 GND 0.004328f
C2232 VDD.n1650 GND 0.004328f
C2233 VDD.n1651 GND 0.004328f
C2234 VDD.n1652 GND 0.004328f
C2235 VDD.n1653 GND 0.004328f
C2236 VDD.n1654 GND 0.004328f
C2237 VDD.n1655 GND 0.004328f
C2238 VDD.n1656 GND 0.004328f
C2239 VDD.n1657 GND 0.004328f
C2240 VDD.n1658 GND 0.004328f
C2241 VDD.n1659 GND 0.004328f
C2242 VDD.n1660 GND 0.004328f
C2243 VDD.n1661 GND 0.004328f
C2244 VDD.n1662 GND 0.004328f
C2245 VDD.n1663 GND 0.004328f
C2246 VDD.n1664 GND 0.004328f
C2247 VDD.n1665 GND 0.004328f
C2248 VDD.n1666 GND 0.004328f
C2249 VDD.n1667 GND 0.004328f
C2250 VDD.n1668 GND 0.004328f
C2251 VDD.n1669 GND 0.004328f
C2252 VDD.n1670 GND 0.004328f
C2253 VDD.n1671 GND 0.009986f
C2254 VDD.n1672 GND 0.009986f
C2255 VDD.n1673 GND 0.010125f
C2256 VDD.n1674 GND 0.004328f
C2257 VDD.n1675 GND 0.004328f
C2258 VDD.n1676 GND 0.004328f
C2259 VDD.n1677 GND 0.004328f
C2260 VDD.n1678 GND 0.004328f
C2261 VDD.n1679 GND 0.002291f
C2262 VDD.n1680 GND 0.00534f
C2263 VDD.n1681 GND 0.0042f
C2264 VDD.n1682 GND 0.004328f
C2265 VDD.n1683 GND 0.004328f
C2266 VDD.n1684 GND 0.004328f
C2267 VDD.n1685 GND 0.004328f
C2268 VDD.n1686 GND 0.004328f
C2269 VDD.n1687 GND 0.004328f
C2270 VDD.n1688 GND 0.003246f
C2271 VDD.n1689 GND 0.12184f
C2272 VDD.n1690 GND 0.003246f
C2273 VDD.n1691 GND 0.004328f
C2274 VDD.n1692 GND 0.004328f
C2275 VDD.n1693 GND 0.004328f
C2276 VDD.n1694 GND 0.004328f
C2277 VDD.n1695 GND 0.004328f
C2278 VDD.n1696 GND 0.004328f
C2279 VDD.n1697 GND 0.004328f
C2280 VDD.n1698 GND 0.004328f
C2281 VDD.n1699 GND 0.004328f
C2282 VDD.n1700 GND 0.004328f
C2283 VDD.n1701 GND 0.004328f
C2284 VDD.n1702 GND 0.010125f
C2285 VDD.n1703 GND 0.010125f
C2286 VDD.n1705 GND 1.60801f
C2287 VDD.n1706 GND 0.010125f
C2288 VDD.n1707 GND 0.010125f
C2289 VDD.n1708 GND 0.009986f
C2290 VDD.n1709 GND 0.004328f
C2291 VDD.n1710 GND 0.004328f
C2292 VDD.n1711 GND 0.32066f
C2293 VDD.n1712 GND 0.004328f
C2294 VDD.n1713 GND 0.004328f
C2295 VDD.n1714 GND 0.004328f
C2296 VDD.n1715 GND 0.004328f
C2297 VDD.n1716 GND 0.004328f
C2298 VDD.n1717 GND 0.32066f
C2299 VDD.n1718 GND 0.004328f
C2300 VDD.n1719 GND 0.004328f
C2301 VDD.n1720 GND 0.004328f
C2302 VDD.n1721 GND 0.004328f
C2303 VDD.n1722 GND 0.004328f
C2304 VDD.n1723 GND 0.32066f
C2305 VDD.n1724 GND 0.004328f
C2306 VDD.n1725 GND 0.004328f
C2307 VDD.n1726 GND 0.004328f
C2308 VDD.n1727 GND 0.004328f
C2309 VDD.n1728 GND 0.004328f
C2310 VDD.n1729 GND 0.132036f
C2311 VDD.n1730 GND 0.004328f
C2312 VDD.n1731 GND 0.004328f
C2313 VDD.n1732 GND 0.004328f
C2314 VDD.n1733 GND 0.004328f
C2315 VDD.n1734 GND 0.004328f
C2316 VDD.n1735 GND 0.32066f
C2317 VDD.n1736 GND 0.004328f
C2318 VDD.n1737 GND 0.004328f
C2319 VDD.n1738 GND 0.004328f
C2320 VDD.n1739 GND 0.004328f
C2321 VDD.n1740 GND 0.004328f
C2322 VDD.n1741 GND 0.32066f
C2323 VDD.n1742 GND 0.004328f
C2324 VDD.n1743 GND 0.004328f
C2325 VDD.n1744 GND 0.004328f
C2326 VDD.n1745 GND 0.004328f
C2327 VDD.n1746 GND 0.004328f
C2328 VDD.n1747 GND 0.32066f
C2329 VDD.n1748 GND 0.004328f
C2330 VDD.n1749 GND 0.004328f
C2331 VDD.n1750 GND 0.004328f
C2332 VDD.n1751 GND 0.004328f
C2333 VDD.n1752 GND 0.004328f
C2334 VDD.n1753 GND 0.32066f
C2335 VDD.n1754 GND 0.004328f
C2336 VDD.n1755 GND 0.004328f
C2337 VDD.n1756 GND 0.004328f
C2338 VDD.n1757 GND 0.004328f
C2339 VDD.n1758 GND 0.004328f
C2340 VDD.n1759 GND 0.32066f
C2341 VDD.n1760 GND 0.004328f
C2342 VDD.n1761 GND 0.004328f
C2343 VDD.n1762 GND 0.004328f
C2344 VDD.n1763 GND 0.004328f
C2345 VDD.n1764 GND 0.004328f
C2346 VDD.n1765 GND 0.32066f
C2347 VDD.n1766 GND 0.004328f
C2348 VDD.n1767 GND 0.004328f
C2349 VDD.n1768 GND 0.004328f
C2350 VDD.n1769 GND 0.004328f
C2351 VDD.n1770 GND 0.004328f
C2352 VDD.n1771 GND 0.32066f
C2353 VDD.n1772 GND 0.004328f
C2354 VDD.n1773 GND 0.004328f
C2355 VDD.n1774 GND 0.004328f
C2356 VDD.n1775 GND 0.004328f
C2357 VDD.n1776 GND 0.004328f
C2358 VDD.t16 GND 0.32066f
C2359 VDD.n1777 GND 0.004328f
C2360 VDD.n1778 GND 0.004328f
C2361 VDD.n1779 GND 0.004328f
C2362 VDD.n1780 GND 0.004328f
C2363 VDD.n1781 GND 0.004328f
C2364 VDD.n1782 GND 0.32066f
C2365 VDD.n1783 GND 0.004328f
C2366 VDD.n1784 GND 0.004328f
C2367 VDD.n1785 GND 0.004328f
C2368 VDD.n1786 GND 0.004328f
C2369 VDD.n1787 GND 0.004328f
C2370 VDD.n1788 GND 0.32066f
C2371 VDD.n1789 GND 0.004328f
C2372 VDD.n1790 GND 0.004328f
C2373 VDD.n1791 GND 0.004328f
C2374 VDD.n1792 GND 0.004328f
C2375 VDD.n1793 GND 0.004328f
C2376 VDD.n1794 GND 0.216917f
C2377 VDD.n1795 GND 0.004328f
C2378 VDD.n1796 GND 0.004328f
C2379 VDD.n1797 GND 0.004328f
C2380 VDD.n1798 GND 0.004328f
C2381 VDD.n1799 GND 0.004328f
C2382 VDD.n1800 GND 0.32066f
C2383 VDD.n1801 GND 0.004328f
C2384 VDD.n1802 GND 0.004328f
C2385 VDD.n1803 GND 0.004328f
C2386 VDD.n1804 GND 0.004328f
C2387 VDD.n1805 GND 0.004328f
C2388 VDD.n1806 GND 0.32066f
C2389 VDD.n1807 GND 0.004328f
C2390 VDD.n1808 GND 0.004328f
C2391 VDD.n1809 GND 0.004328f
C2392 VDD.n1810 GND 0.004328f
C2393 VDD.n1811 GND 0.004328f
C2394 VDD.n1812 GND 0.32066f
C2395 VDD.n1813 GND 0.004328f
C2396 VDD.n1814 GND 0.004328f
C2397 VDD.n1815 GND 0.004328f
C2398 VDD.n1816 GND 0.004328f
C2399 VDD.n1817 GND 0.004328f
C2400 VDD.n1818 GND 0.32066f
C2401 VDD.n1819 GND 0.004328f
C2402 VDD.n1820 GND 0.004328f
C2403 VDD.n1821 GND 0.004328f
C2404 VDD.n1822 GND 0.004328f
C2405 VDD.n1823 GND 0.004328f
C2406 VDD.n1824 GND 0.235779f
C2407 VDD.n1825 GND 0.004328f
C2408 VDD.n1826 GND 0.004328f
C2409 VDD.n1827 GND 0.004328f
C2410 VDD.n1828 GND 0.004328f
C2411 VDD.n1829 GND 0.004328f
C2412 VDD.n1830 GND 0.004328f
C2413 VDD.n1831 GND 0.004328f
C2414 VDD.n1832 GND 0.004328f
C2415 VDD.n1833 GND 0.004328f
C2416 VDD.n1834 GND 0.004328f
C2417 VDD.n1835 GND 0.207486f
C2418 VDD.n1836 GND 0.004328f
C2419 VDD.n1837 GND 0.004328f
C2420 VDD.n1838 GND 0.004328f
C2421 VDD.n1839 GND 0.004328f
C2422 VDD.n1840 GND 0.004328f
C2423 VDD.n1841 GND 0.32066f
C2424 VDD.n1842 GND 0.004328f
C2425 VDD.n1843 GND 0.004328f
C2426 VDD.n1844 GND 0.004328f
C2427 VDD.n1845 GND 0.004328f
C2428 VDD.n1846 GND 0.010503f
C2429 VDD.n1847 GND 0.009986f
C2430 VDD.n1848 GND 0.010125f
C2431 VDD.n1849 GND 0.009608f
C2432 VDD.n1850 GND 0.004328f
C2433 VDD.n1851 GND 0.004328f
C2434 VDD.n1852 GND 0.004328f
C2435 VDD.n1853 GND 0.004328f
C2436 VDD.n1854 GND 0.002291f
C2437 VDD.n1855 GND 0.004328f
C2438 VDD.n1856 GND 0.004328f
C2439 VDD.n1857 GND 0.0042f
C2440 VDD.n1858 GND 0.004328f
C2441 VDD.n1859 GND 0.004328f
C2442 VDD.n1860 GND 0.004328f
C2443 VDD.n1861 GND 0.004328f
C2444 VDD.n1862 GND 0.004328f
C2445 VDD.n1863 GND 0.004328f
C2446 VDD.n1864 GND 0.004328f
C2447 VDD.n1865 GND 0.004328f
C2448 VDD.n1866 GND 0.004328f
C2449 VDD.n1867 GND 0.004328f
C2450 VDD.n1868 GND 0.004328f
C2451 VDD.n1869 GND 0.004328f
C2452 VDD.n1870 GND 0.004328f
C2453 VDD.n1871 GND 0.004328f
C2454 VDD.n1872 GND 0.004328f
C2455 VDD.n1873 GND 0.004328f
C2456 VDD.n1874 GND 0.004328f
C2457 VDD.n1875 GND 0.004328f
C2458 VDD.n1876 GND 0.004328f
C2459 VDD.n1877 GND 0.004328f
C2460 VDD.n1878 GND 0.010125f
C2461 VDD.n1879 GND 0.010125f
C2462 VDD.n1880 GND 0.009986f
C2463 VDD.n1881 GND 0.004328f
C2464 VDD.n1882 GND 0.004328f
C2465 VDD.n1883 GND 0.32066f
C2466 VDD.n1884 GND 0.004328f
C2467 VDD.n1885 GND 0.009986f
C2468 VDD.n1886 GND 0.010503f
C2469 VDD.n1887 GND 0.009608f
C2470 VDD.n1888 GND 0.004328f
C2471 VDD.n1889 GND 0.004328f
C2472 VDD.n1890 GND 0.004328f
C2473 VDD.n1891 GND 0.004328f
C2474 VDD.n1892 GND 0.004328f
C2475 VDD.n1893 GND 0.002291f
C2476 VDD.n1894 GND 0.00534f
C2477 VDD.n1895 GND 0.0042f
C2478 VDD.n1896 GND 0.004328f
C2479 VDD.n1897 GND 0.004328f
C2480 VDD.n1898 GND 0.004328f
C2481 VDD.n1899 GND 0.004328f
C2482 VDD.n1900 GND 0.004328f
C2483 VDD.n1901 GND 0.004328f
C2484 VDD.n1902 GND 0.004328f
C2485 VDD.n1903 GND 0.004328f
C2486 VDD.n1904 GND 0.004328f
C2487 VDD.n1905 GND 0.004328f
C2488 VDD.n1906 GND 0.004328f
C2489 VDD.n1907 GND 0.004328f
C2490 VDD.n1908 GND 0.004328f
C2491 VDD.n1909 GND 0.004328f
C2492 VDD.n1910 GND 0.004328f
C2493 VDD.n1911 GND 0.004328f
C2494 VDD.n1912 GND 0.004328f
C2495 VDD.n1913 GND 0.004328f
C2496 VDD.n1914 GND 0.004328f
C2497 VDD.n1915 GND 0.004328f
C2498 VDD.n1916 GND 0.010125f
C2499 VDD.n1917 GND 0.010125f
C2500 VDD.n1918 GND 1.96876f
C2501 VDD.n1925 GND 0.010125f
C2502 VDD.n1932 GND 0.004328f
C2503 VDD.t55 GND 0.066005f
C2504 VDD.t52 GND 0.213596f
C2505 VDD.n1933 GND 0.071628f
C2506 VDD.t54 GND 0.048572f
C2507 VDD.n1934 GND 0.068504f
C2508 VDD.n1935 GND 0.00534f
C2509 VDD.n1936 GND 0.004328f
C2510 VDD.n1937 GND 0.004328f
C2511 VDD.n1938 GND 0.004328f
C2512 VDD.n1939 GND 0.004328f
C2513 VDD.n1940 GND 0.004328f
C2514 VDD.n1941 GND 0.004328f
C2515 VDD.n1942 GND 0.004328f
C2516 VDD.n1943 GND 0.004328f
C2517 VDD.n1944 GND 0.004328f
C2518 VDD.n1945 GND 0.004328f
C2519 VDD.n1946 GND 0.004328f
C2520 VDD.n1947 GND 0.004328f
C2521 VDD.n1948 GND 0.004328f
C2522 VDD.n1949 GND 0.004328f
C2523 VDD.n1950 GND 0.004328f
C2524 VDD.n1951 GND 0.004328f
C2525 VDD.n1952 GND 0.004328f
C2526 VDD.n1953 GND 0.004328f
C2527 VDD.n1954 GND 0.004328f
C2528 VDD.n1955 GND 0.004328f
C2529 VDD.n1956 GND 0.004328f
C2530 VDD.n1957 GND 0.004328f
C2531 VDD.n1958 GND 0.004328f
C2532 VDD.n1959 GND 0.004328f
C2533 VDD.n1960 GND 0.004328f
C2534 VDD.n1961 GND 0.004328f
C2535 VDD.n1962 GND 0.004328f
C2536 VDD.n1963 GND 0.004328f
C2537 VDD.n1964 GND 0.004328f
C2538 VDD.n1965 GND 0.004328f
C2539 VDD.n1966 GND 0.004328f
C2540 VDD.n1967 GND 0.004328f
C2541 VDD.n1968 GND 0.004328f
C2542 VDD.n1969 GND 0.004328f
C2543 VDD.n1970 GND 0.004328f
C2544 VDD.n1971 GND 0.004328f
C2545 VDD.n1972 GND 0.004328f
C2546 VDD.n1973 GND 0.004328f
C2547 VDD.n1974 GND 0.004328f
C2548 VDD.n1975 GND 0.004328f
C2549 VDD.n1976 GND 0.004328f
C2550 VDD.n1977 GND 0.004328f
C2551 VDD.n1978 GND 0.004328f
C2552 VDD.n1979 GND 0.004328f
C2553 VDD.n1980 GND 0.004328f
C2554 VDD.n1981 GND 0.004328f
C2555 VDD.n1982 GND 0.004328f
C2556 VDD.n1983 GND 0.004328f
C2557 VDD.n1984 GND 0.004328f
C2558 VDD.n1985 GND 0.004328f
C2559 VDD.n1986 GND 0.004328f
C2560 VDD.n1987 GND 0.004328f
C2561 VDD.n1988 GND 0.004328f
C2562 VDD.n1989 GND 0.004328f
C2563 VDD.n1990 GND 0.004328f
C2564 VDD.n1991 GND 0.004328f
C2565 VDD.n1992 GND 0.004328f
C2566 VDD.n1993 GND 0.004328f
C2567 VDD.n1994 GND 0.004328f
C2568 VDD.n1995 GND 0.004328f
C2569 VDD.n1996 GND 0.004328f
C2570 VDD.n1997 GND 0.004328f
C2571 VDD.n1998 GND 0.004328f
C2572 VDD.n1999 GND 0.004328f
C2573 VDD.n2000 GND 0.009986f
C2574 VDD.n2001 GND 0.009986f
C2575 VDD.n2002 GND 0.010125f
C2576 VDD.n2003 GND 0.010125f
C2577 VDD.n2004 GND 0.004328f
C2578 VDD.n2005 GND 0.004328f
C2579 VDD.n2006 GND 0.004328f
C2580 VDD.n2007 GND 0.004328f
C2581 VDD.n2008 GND 0.002291f
C2582 VDD.n2009 GND 0.004328f
C2583 VDD.n2010 GND 0.004328f
C2584 VDD.n2011 GND 0.0042f
C2585 VDD.n2012 GND 0.004328f
C2586 VDD.n2013 GND 0.004328f
C2587 VDD.n2014 GND 0.004328f
C2588 VDD.n2015 GND 0.004328f
C2589 VDD.n2016 GND 0.004328f
C2590 VDD.n2017 GND 0.004328f
C2591 VDD.n2018 GND 0.004328f
C2592 VDD.n2019 GND 0.004328f
C2593 VDD.n2020 GND 0.004328f
C2594 VDD.n2021 GND 0.004328f
C2595 VDD.n2022 GND 0.004328f
C2596 VDD.n2023 GND 0.004328f
C2597 VDD.n2024 GND 0.004328f
C2598 VDD.n2025 GND 0.004328f
C2599 VDD.n2026 GND 0.004328f
C2600 VDD.n2027 GND 0.004328f
C2601 VDD.n2028 GND 0.004328f
C2602 VDD.n2030 GND 0.004328f
C2603 VDD.n2031 GND 0.004328f
C2604 VDD.t121 GND 0.066005f
C2605 VDD.t119 GND 0.213596f
C2606 VDD.n2032 GND 0.071628f
C2607 VDD.t120 GND 0.048572f
C2608 VDD.n2033 GND 0.068504f
C2609 VDD.n2034 GND 0.004328f
C2610 VDD.n2035 GND 0.004328f
C2611 VDD.n2036 GND 0.004328f
C2612 VDD.n2037 GND 0.004328f
C2613 VDD.n2038 GND 0.004328f
C2614 VDD.n2039 GND 0.004328f
C2615 VDD.n2040 GND 0.004328f
C2616 VDD.n2041 GND 0.004328f
C2617 VDD.n2042 GND 0.004328f
C2618 VDD.n2043 GND 0.004328f
C2619 VDD.n2044 GND 0.004328f
C2620 VDD.n2045 GND 0.004328f
C2621 VDD.n2046 GND 0.004328f
C2622 VDD.n2047 GND 0.004328f
C2623 VDD.n2048 GND 0.004328f
C2624 VDD.n2049 GND 0.004328f
C2625 VDD.n2050 GND 0.004328f
C2626 VDD.n2051 GND 0.004328f
C2627 VDD.n2052 GND 0.004328f
C2628 VDD.n2053 GND 0.004328f
C2629 VDD.n2054 GND 0.004328f
C2630 VDD.n2055 GND 0.004328f
C2631 VDD.n2056 GND 0.004328f
C2632 VDD.n2057 GND 0.004328f
C2633 VDD.n2058 GND 0.004328f
C2634 VDD.n2059 GND 0.004328f
C2635 VDD.n2060 GND 0.004328f
C2636 VDD.n2061 GND 0.004328f
C2637 VDD.n2062 GND 0.004328f
C2638 VDD.n2063 GND 0.004328f
C2639 VDD.n2064 GND 0.004328f
C2640 VDD.n2065 GND 0.004328f
C2641 VDD.n2066 GND 0.004328f
C2642 VDD.n2067 GND 0.004328f
C2643 VDD.n2068 GND 0.004328f
C2644 VDD.n2069 GND 0.004328f
C2645 VDD.n2070 GND 0.004328f
C2646 VDD.n2071 GND 0.004328f
C2647 VDD.n2072 GND 0.004328f
C2648 VDD.n2073 GND 0.004328f
C2649 VDD.n2074 GND 0.004328f
C2650 VDD.n2075 GND 0.004328f
C2651 VDD.n2076 GND 0.004328f
C2652 VDD.n2077 GND 0.004328f
C2653 VDD.n2078 GND 0.004328f
C2654 VDD.n2079 GND 0.004328f
C2655 VDD.n2080 GND 0.004328f
C2656 VDD.n2081 GND 0.004328f
C2657 VDD.n2082 GND 0.004328f
C2658 VDD.n2083 GND 0.004328f
C2659 VDD.n2084 GND 0.004328f
C2660 VDD.n2085 GND 0.004328f
C2661 VDD.n2086 GND 0.004328f
C2662 VDD.n2087 GND 0.004328f
C2663 VDD.n2088 GND 0.004328f
C2664 VDD.n2089 GND 0.004328f
C2665 VDD.n2090 GND 0.004328f
C2666 VDD.n2091 GND 0.004328f
C2667 VDD.n2092 GND 0.004328f
C2668 VDD.n2093 GND 0.004328f
C2669 VDD.n2094 GND 0.004328f
C2670 VDD.n2095 GND 0.004328f
C2671 VDD.n2096 GND 0.009986f
C2672 VDD.n2097 GND 0.009986f
C2673 VDD.n2098 GND 0.010125f
C2674 VDD.n2099 GND 0.004328f
C2675 VDD.n2100 GND 0.004328f
C2676 VDD.n2101 GND 0.004328f
C2677 VDD.n2102 GND 0.004328f
C2678 VDD.n2103 GND 0.004328f
C2679 VDD.n2104 GND 0.002291f
C2680 VDD.n2105 GND 0.00534f
C2681 VDD.n2106 GND 0.0042f
C2682 VDD.n2107 GND 0.004328f
C2683 VDD.n2108 GND 0.004328f
C2684 VDD.n2109 GND 0.004328f
C2685 VDD.n2110 GND 0.004328f
C2686 VDD.n2111 GND 0.004328f
C2687 VDD.n2112 GND 0.004328f
C2688 VDD.n2113 GND 0.004328f
C2689 VDD.n2114 GND 0.004328f
C2690 VDD.n2115 GND 0.004328f
C2691 VDD.n2116 GND 0.004328f
C2692 VDD.n2117 GND 0.004328f
C2693 VDD.n2118 GND 0.004328f
C2694 VDD.n2119 GND 0.004328f
C2695 VDD.n2120 GND 0.004328f
C2696 VDD.n2121 GND 0.004328f
C2697 VDD.n2122 GND 0.004328f
C2698 VDD.n2123 GND 0.004328f
C2699 VDD.n2124 GND 0.004328f
C2700 VDD.n2125 GND 0.004328f
C2701 VDD.n2126 GND 0.010125f
C2702 VDD.n2127 GND 0.010125f
C2703 VDD.n2129 GND 1.96876f
C2704 VDD.n2131 GND 0.010125f
C2705 VDD.n2132 GND 0.010125f
C2706 VDD.n2133 GND 0.009986f
C2707 VDD.n2134 GND 0.004328f
C2708 VDD.n2135 GND 0.004328f
C2709 VDD.n2136 GND 0.32066f
C2710 VDD.n2137 GND 0.004328f
C2711 VDD.n2138 GND 0.004328f
C2712 VDD.n2139 GND 0.004328f
C2713 VDD.n2140 GND 0.004328f
C2714 VDD.n2141 GND 0.004328f
C2715 VDD.n2142 GND 0.32066f
C2716 VDD.n2143 GND 0.004328f
C2717 VDD.n2144 GND 0.004328f
C2718 VDD.n2145 GND 0.004328f
C2719 VDD.n2146 GND 0.004328f
C2720 VDD.n2147 GND 0.004328f
C2721 VDD.n2148 GND 0.207486f
C2722 VDD.n2149 GND 0.004328f
C2723 VDD.n2150 GND 0.004328f
C2724 VDD.n2151 GND 0.004328f
C2725 VDD.n2152 GND 0.004328f
C2726 VDD.n2153 GND 0.004328f
C2727 VDD.n2154 GND 0.235779f
C2728 VDD.n2155 GND 0.004328f
C2729 VDD.n2156 GND 0.004328f
C2730 VDD.n2157 GND 0.004328f
C2731 VDD.n2158 GND 0.004328f
C2732 VDD.n2159 GND 0.004328f
C2733 VDD.n2160 GND 0.32066f
C2734 VDD.n2161 GND 0.004328f
C2735 VDD.n2162 GND 0.004328f
C2736 VDD.n2163 GND 0.004328f
C2737 VDD.n2164 GND 0.004328f
C2738 VDD.n2165 GND 0.004328f
C2739 VDD.n2166 GND 0.32066f
C2740 VDD.n2167 GND 0.004328f
C2741 VDD.n2168 GND 0.004328f
C2742 VDD.n2169 GND 0.004328f
C2743 VDD.n2170 GND 0.004328f
C2744 VDD.n2171 GND 0.004328f
C2745 VDD.n2172 GND 0.32066f
C2746 VDD.n2173 GND 0.004328f
C2747 VDD.n2174 GND 0.004328f
C2748 VDD.n2175 GND 0.004328f
C2749 VDD.n2176 GND 0.004328f
C2750 VDD.n2177 GND 0.004328f
C2751 VDD.n2178 GND 0.32066f
C2752 VDD.n2179 GND 0.004328f
C2753 VDD.n2180 GND 0.004328f
C2754 VDD.n2181 GND 0.004328f
C2755 VDD.n2182 GND 0.004328f
C2756 VDD.n2183 GND 0.004328f
C2757 VDD.n2184 GND 0.216917f
C2758 VDD.n2185 GND 0.004328f
C2759 VDD.n2186 GND 0.004328f
C2760 VDD.n2187 GND 0.004328f
C2761 VDD.n2188 GND 0.004328f
C2762 VDD.n2189 GND 0.004328f
C2763 VDD.n2190 GND 0.32066f
C2764 VDD.n2191 GND 0.004328f
C2765 VDD.n2192 GND 0.004328f
C2766 VDD.n2193 GND 0.004328f
C2767 VDD.n2194 GND 0.004328f
C2768 VDD.n2195 GND 0.004328f
C2769 VDD.n2196 GND 0.32066f
C2770 VDD.n2197 GND 0.004328f
C2771 VDD.n2198 GND 0.004328f
C2772 VDD.n2199 GND 0.004328f
C2773 VDD.n2200 GND 0.004328f
C2774 VDD.n2201 GND 0.004328f
C2775 VDD.t23 GND 0.32066f
C2776 VDD.n2202 GND 0.004328f
C2777 VDD.n2203 GND 0.004328f
C2778 VDD.n2204 GND 0.004328f
C2779 VDD.n2205 GND 0.004328f
C2780 VDD.n2206 GND 0.004328f
C2781 VDD.n2207 GND 0.32066f
C2782 VDD.n2208 GND 0.004328f
C2783 VDD.n2209 GND 0.004328f
C2784 VDD.n2210 GND 0.004328f
C2785 VDD.n2211 GND 0.004328f
C2786 VDD.n2212 GND 0.004328f
C2787 VDD.n2213 GND 0.32066f
C2788 VDD.n2214 GND 0.004328f
C2789 VDD.n2215 GND 0.004328f
C2790 VDD.n2216 GND 0.004328f
C2791 VDD.n2217 GND 0.004328f
C2792 VDD.n2218 GND 0.004328f
C2793 VDD.n2219 GND 0.32066f
C2794 VDD.n2220 GND 0.004328f
C2795 VDD.n2221 GND 0.004328f
C2796 VDD.n2222 GND 0.004328f
C2797 VDD.n2223 GND 0.004328f
C2798 VDD.n2224 GND 0.004328f
C2799 VDD.n2225 GND 0.32066f
C2800 VDD.n2226 GND 0.004328f
C2801 VDD.n2227 GND 0.004328f
C2802 VDD.n2228 GND 0.004328f
C2803 VDD.n2229 GND 0.004328f
C2804 VDD.n2230 GND 0.004328f
C2805 VDD.n2231 GND 0.32066f
C2806 VDD.n2232 GND 0.004328f
C2807 VDD.n2233 GND 0.004328f
C2808 VDD.n2234 GND 0.004328f
C2809 VDD.n2235 GND 0.004328f
C2810 VDD.n2236 GND 0.004328f
C2811 VDD.n2237 GND 0.32066f
C2812 VDD.n2238 GND 0.004328f
C2813 VDD.n2239 GND 0.004328f
C2814 VDD.n2240 GND 0.004328f
C2815 VDD.n2241 GND 0.004328f
C2816 VDD.n2242 GND 0.004328f
C2817 VDD.n2243 GND 0.32066f
C2818 VDD.n2244 GND 0.004328f
C2819 VDD.n2245 GND 0.004328f
C2820 VDD.n2246 GND 0.004328f
C2821 VDD.n2247 GND 0.004328f
C2822 VDD.n2248 GND 0.004328f
C2823 VDD.n2249 GND 0.132036f
C2824 VDD.n2250 GND 0.004328f
C2825 VDD.n2251 GND 0.004328f
C2826 VDD.n2252 GND 0.004328f
C2827 VDD.n2253 GND 0.010125f
C2828 VDD.n2254 GND 0.004328f
C2829 VDD.n2255 GND 0.004328f
C2830 VDD.n2258 GND 0.004328f
C2831 VDD.n2259 GND 0.004328f
C2832 VDD.n2260 GND 0.004328f
C2833 VDD.n2261 GND 0.004328f
C2834 VDD.n2263 GND 0.004328f
C2835 VDD.n2264 GND 0.004328f
C2836 VDD.n2265 GND 0.004328f
C2837 VDD.n2266 GND 0.004328f
C2838 VDD.n2267 GND 0.004328f
C2839 VDD.n2268 GND 0.004328f
C2840 VDD.n2270 GND 0.010125f
C2841 VDD.n2271 GND 0.009986f
C2842 VDD.n2272 GND 0.009986f
C2843 VDD.n2273 GND 0.004328f
C2844 VDD.n2274 GND 0.004328f
C2845 VDD.n2275 GND 0.004328f
C2846 VDD.n2276 GND 0.004328f
C2847 VDD.n2277 GND 0.004328f
C2848 VDD.n2278 GND 0.004328f
C2849 VDD.n2279 GND 0.004328f
C2850 VDD.n2280 GND 0.32066f
C2851 VDD.n2281 GND 0.004328f
C2852 VDD.n2282 GND 0.004328f
C2853 VDD.n2283 GND 0.004328f
C2854 VDD.n2284 GND 0.004328f
C2855 VDD.n2285 GND 0.004328f
C2856 VDD.n2286 GND 0.32066f
C2857 VDD.n2287 GND 0.004328f
C2858 VDD.n2288 GND 0.004328f
C2859 VDD.n2289 GND 0.004328f
C2860 VDD.n2290 GND 0.004328f
C2861 VDD.n2291 GND 0.010503f
C2862 VDD.n2292 GND 0.009608f
C2863 VDD.n2293 GND 0.010125f
C2864 VDD.n2295 GND 0.004328f
C2865 VDD.n2296 GND 0.004328f
C2866 VDD.n2297 GND 0.004328f
C2867 VDD.n2298 GND 0.002291f
C2868 VDD.n2299 GND 0.00534f
C2869 VDD.n2300 GND 0.0042f
C2870 VDD.n2301 GND 0.004328f
C2871 VDD.n2303 GND 0.004328f
C2872 VDD.n2304 GND 0.004328f
C2873 VDD.n2305 GND 0.004328f
C2874 VDD.n2306 GND 0.003246f
C2875 VDD.n2307 GND 0.119615f
C2876 VDD.n2308 GND 0.003246f
C2877 VDD.n2309 GND 0.004328f
C2878 VDD.n2311 GND 0.004328f
C2879 VDD.n2312 GND 0.004328f
C2880 VDD.n2313 GND 0.004328f
C2881 VDD.n2314 GND 0.004328f
C2882 VDD.n2315 GND 0.004328f
C2883 VDD.n2316 GND 0.004328f
C2884 VDD.n2318 GND 0.004328f
C2885 VDD.n2319 GND 0.004328f
C2886 VDD.n2321 GND 0.010125f
C2887 VDD.n2322 GND 0.010125f
C2888 VDD.n2323 GND 0.009986f
C2889 VDD.n2324 GND 0.004328f
C2890 VDD.n2325 GND 0.004328f
C2891 VDD.n2326 GND 0.32066f
C2892 VDD.n2327 GND 0.004328f
C2893 VDD.n2328 GND 0.004328f
C2894 VDD.n2329 GND 0.010503f
C2895 VDD.n2330 GND 0.009608f
C2896 VDD.n2331 GND 0.010125f
C2897 VDD.n2333 GND 0.004328f
C2898 VDD.n2334 GND 0.004328f
C2899 VDD.n2335 GND 0.004328f
C2900 VDD.n2336 GND 0.002291f
C2901 VDD.n2337 GND 0.00534f
C2902 VDD.n2338 GND 0.0042f
C2903 VDD.n2339 GND 0.004328f
C2904 VDD.n2341 GND 0.004328f
C2905 VDD.n2342 GND 0.004328f
C2906 VDD.n2344 GND 0.004328f
C2907 VDD.n2345 GND 0.003246f
C2908 VDD.n2346 GND 0.119615f
C2909 VDD.n2347 GND 0.005122f
C2910 VDD.n2349 GND 0.006364f
C2911 VDD.n2350 GND 0.006364f
C2912 VDD.n2351 GND 0.005122f
C2913 VDD.n2352 GND 0.006364f
C2914 VDD.n2353 GND 0.006364f
C2915 VDD.n2354 GND 0.006364f
C2916 VDD.n2355 GND 0.006364f
C2917 VDD.n2356 GND 0.006364f
C2918 VDD.n2357 GND 0.005122f
C2919 VDD.n2359 GND 0.006364f
C2920 VDD.n2360 GND 0.006364f
C2921 VDD.n2361 GND 0.006364f
C2922 VDD.n2362 GND 0.006364f
C2923 VDD.n2363 GND 0.002331f
C2924 VDD.t100 GND 0.123904f
C2925 VDD.t98 GND 0.415248f
C2926 VDD.n2364 GND 0.086184f
C2927 VDD.t99 GND 0.090617f
C2928 VDD.n2365 GND 0.088946f
C2929 VDD.n2366 GND 0.007043f
C2930 VDD.n2367 GND 0.002792f
C2931 VDD.n2368 GND 0.005122f
C2932 VDD.n2369 GND 0.006364f
C2933 VDD.n2371 GND 0.006364f
C2934 VDD.n2373 GND 0.006364f
C2935 VDD.n2374 GND 0.005122f
C2936 VDD.n2375 GND 0.005122f
C2937 VDD.n2376 GND 0.005122f
C2938 VDD.n2377 GND 0.006364f
C2939 VDD.n2379 GND 0.006364f
C2940 VDD.n2381 GND 0.006364f
C2941 VDD.n2382 GND 0.005122f
C2942 VDD.n2383 GND 0.005122f
C2943 VDD.n2385 GND 1.50188f
C2944 VDD.n2387 GND 0.005122f
C2945 VDD.n2388 GND 0.006364f
C2946 VDD.n2390 GND 0.006364f
C2947 VDD.n2392 GND 0.006364f
C2948 VDD.n2393 GND 0.003304f
C2949 VDD.t94 GND 0.123904f
C2950 VDD.t92 GND 0.415248f
C2951 VDD.n2394 GND 0.086184f
C2952 VDD.t93 GND 0.090617f
C2953 VDD.n2395 GND 0.088946f
C2954 VDD.n2396 GND 0.007043f
C2955 VDD.n2397 GND 0.002689f
C2956 VDD.n2398 GND 0.005122f
C2957 VDD.n2399 GND 0.006364f
C2958 VDD.n2401 GND 0.006364f
C2959 VDD.n2403 GND 0.006364f
C2960 VDD.n2404 GND 0.005122f
C2961 VDD.n2405 GND 0.005122f
C2962 VDD.n2406 GND 0.005122f
C2963 VDD.n2407 GND 0.006364f
C2964 VDD.n2409 GND 0.006364f
C2965 VDD.n2411 GND 0.006364f
C2966 VDD.n2412 GND 0.005122f
C2967 VDD.n2413 GND 0.005122f
C2968 VDD.n2414 GND 0.005122f
C2969 VDD.n2415 GND 0.006364f
C2970 VDD.n2417 GND 0.006364f
C2971 VDD.n2419 GND 0.006364f
C2972 VDD.n2420 GND 0.005122f
C2973 VDD.n2421 GND 0.005122f
C2974 VDD.n2422 GND 0.003406f
C2975 VDD.n2423 GND 0.006364f
C2976 VDD.n2425 GND 0.006364f
C2977 VDD.n2427 GND 0.006364f
C2978 VDD.n2428 GND 0.005122f
C2979 VDD.n2429 GND 0.005122f
C2980 VDD.n2430 GND 0.005122f
C2981 VDD.n2431 GND 0.006364f
C2982 VDD.n2433 GND 0.006364f
C2983 VDD.n2435 GND 0.006364f
C2984 VDD.n2436 GND 0.005122f
C2985 VDD.n2437 GND 0.005122f
C2986 VDD.n2438 GND 0.005122f
C2987 VDD.n2439 GND 0.006364f
C2988 VDD.n2441 GND 0.006364f
C2989 VDD.n2442 GND 0.006364f
C2990 VDD.n2443 GND 0.005122f
C2991 VDD.n2444 GND 0.005122f
C2992 VDD.n2445 GND 0.006364f
C2993 VDD.n2446 GND 0.006364f
C2994 VDD.n2448 GND 0.006364f
C2995 VDD.n2449 GND 0.005122f
C2996 VDD.n2450 GND 0.003509f
C2997 VDD.n2451 GND 0.009604f
C2998 VDD.n2453 GND 0.005045f
C2999 VDD.n2454 GND 0.006364f
C3000 VDD.n2456 GND 0.006364f
C3001 VDD.n2458 GND 0.006364f
C3002 VDD.n2459 GND 0.005122f
C3003 VDD.n2460 GND 0.005122f
C3004 VDD.n2461 GND 0.005122f
C3005 VDD.n2462 GND 0.006364f
C3006 VDD.n2464 GND 0.006364f
C3007 VDD.n2465 GND 0.006364f
C3008 VDD.n2466 GND 0.005122f
C3009 VDD.n2467 GND 0.005122f
C3010 VDD.n2468 GND 0.006364f
C3011 VDD.n2469 GND 0.006364f
C3012 VDD.n2471 GND 0.006364f
C3013 VDD.n2472 GND 0.005122f
C3014 VDD.n2473 GND 0.004251f
C3015 VDD.n2474 GND 0.01437f
C3016 VDD.n2475 GND 0.014395f
C3017 VDD.n2476 GND 0.004251f
C3018 VDD.n2477 GND 0.014395f
C3019 VDD.n2478 GND 0.598879f
C3020 VDD.n2479 GND 0.014395f
C3021 VDD.n2480 GND 0.004251f
C3022 VDD.n2481 GND 0.014395f
C3023 VDD.n2482 GND 0.006364f
C3024 VDD.n2483 GND 0.006364f
C3025 VDD.n2484 GND 0.005122f
C3026 VDD.n2485 GND 0.006364f
C3027 VDD.n2486 GND 0.471559f
C3028 VDD.n2487 GND 0.006364f
C3029 VDD.n2488 GND 0.005122f
C3030 VDD.n2489 GND 0.006364f
C3031 VDD.n2490 GND 0.006364f
C3032 VDD.n2491 GND 0.006364f
C3033 VDD.n2492 GND 0.005122f
C3034 VDD.n2493 GND 0.006364f
C3035 VDD.n2494 GND 0.471559f
C3036 VDD.n2495 GND 0.006364f
C3037 VDD.n2496 GND 0.005122f
C3038 VDD.n2497 GND 0.006364f
C3039 VDD.n2498 GND 0.006364f
C3040 VDD.n2499 GND 0.006364f
C3041 VDD.n2500 GND 0.005122f
C3042 VDD.n2501 GND 0.006364f
C3043 VDD.n2502 GND 0.424403f
C3044 VDD.n2503 GND 0.006364f
C3045 VDD.n2504 GND 0.005122f
C3046 VDD.n2505 GND 0.006364f
C3047 VDD.n2506 GND 0.006364f
C3048 VDD.n2507 GND 0.006364f
C3049 VDD.n2508 GND 0.005122f
C3050 VDD.n2509 GND 0.006364f
C3051 VDD.n2510 GND 0.471559f
C3052 VDD.n2511 GND 0.006364f
C3053 VDD.n2512 GND 0.005122f
C3054 VDD.n2513 GND 0.006364f
C3055 VDD.n2514 GND 0.006364f
C3056 VDD.n2515 GND 0.006364f
C3057 VDD.n2516 GND 0.005122f
C3058 VDD.n2517 GND 0.006364f
C3059 VDD.n2518 GND 0.471559f
C3060 VDD.n2519 GND 0.006364f
C3061 VDD.n2520 GND 0.005122f
C3062 VDD.n2521 GND 0.006364f
C3063 VDD.n2522 GND 0.006364f
C3064 VDD.n2523 GND 0.006364f
C3065 VDD.n2524 GND 0.005122f
C3066 VDD.n2525 GND 0.006364f
C3067 VDD.n2526 GND 0.471559f
C3068 VDD.n2527 GND 0.006364f
C3069 VDD.n2528 GND 0.005122f
C3070 VDD.n2529 GND 0.006364f
C3071 VDD.n2530 GND 0.006364f
C3072 VDD.n2531 GND 0.006364f
C3073 VDD.n2532 GND 0.005122f
C3074 VDD.n2533 GND 0.006364f
C3075 VDD.n2534 GND 0.471559f
C3076 VDD.n2535 GND 0.006364f
C3077 VDD.n2536 GND 0.005122f
C3078 VDD.n2537 GND 0.006364f
C3079 VDD.n2538 GND 0.006364f
C3080 VDD.n2539 GND 0.006364f
C3081 VDD.n2540 GND 0.005122f
C3082 VDD.n2541 GND 0.006364f
C3083 VDD.n2542 GND 0.471559f
C3084 VDD.n2543 GND 0.006364f
C3085 VDD.n2544 GND 0.005122f
C3086 VDD.n2545 GND 0.006364f
C3087 VDD.n2546 GND 0.006364f
C3088 VDD.n2547 GND 0.006364f
C3089 VDD.n2548 GND 0.005122f
C3090 VDD.n2549 GND 0.006364f
C3091 VDD.n2550 GND 0.466843f
C3092 VDD.n2551 GND 0.006364f
C3093 VDD.n2552 GND 0.005122f
C3094 VDD.n2553 GND 0.006364f
C3095 VDD.n2554 GND 0.006364f
C3096 VDD.n2555 GND 0.006364f
C3097 VDD.n2556 GND 0.005122f
C3098 VDD.n2557 GND 0.006364f
C3099 VDD.n2558 GND 0.471559f
C3100 VDD.n2559 GND 0.006364f
C3101 VDD.n2560 GND 0.005122f
C3102 VDD.n2561 GND 0.006364f
C3103 VDD.n2562 GND 0.006364f
C3104 VDD.n2563 GND 0.006364f
C3105 VDD.n2564 GND 0.005122f
C3106 VDD.n2565 GND 0.006364f
C3107 VDD.n2566 GND 0.471559f
C3108 VDD.n2567 GND 0.006364f
C3109 VDD.n2568 GND 0.005122f
C3110 VDD.n2569 GND 0.006364f
C3111 VDD.n2570 GND 0.006364f
C3112 VDD.n2571 GND 0.006364f
C3113 VDD.n2572 GND 0.005122f
C3114 VDD.n2573 GND 0.006364f
C3115 VDD.n2574 GND 0.471559f
C3116 VDD.n2575 GND 0.006364f
C3117 VDD.n2576 GND 0.005122f
C3118 VDD.n2577 GND 0.006364f
C3119 VDD.n2578 GND 0.006364f
C3120 VDD.n2579 GND 0.006364f
C3121 VDD.n2580 GND 0.005122f
C3122 VDD.n2581 GND 0.005122f
C3123 VDD.n2582 GND 0.005122f
C3124 VDD.n2583 GND 0.006364f
C3125 VDD.n2584 GND 0.006364f
C3126 VDD.n2585 GND 0.006364f
C3127 VDD.n2586 GND 0.005122f
C3128 VDD.n2587 GND 0.005122f
C3129 VDD.n2588 GND 0.005122f
C3130 VDD.n2589 GND 0.006364f
C3131 VDD.n2590 GND 0.006364f
C3132 VDD.n2591 GND 0.006364f
C3133 VDD.n2592 GND 0.005122f
C3134 VDD.n2593 GND 0.005122f
C3135 VDD.n2594 GND 0.005122f
C3136 VDD.n2595 GND 0.006364f
C3137 VDD.n2596 GND 0.006364f
C3138 VDD.n2597 GND 0.006364f
C3139 VDD.n2598 GND 0.005122f
C3140 VDD.n2599 GND 0.005122f
C3141 VDD.n2600 GND 0.005122f
C3142 VDD.n2601 GND 0.006364f
C3143 VDD.n2602 GND 0.006364f
C3144 VDD.n2603 GND 0.006364f
C3145 VDD.n2604 GND 0.005122f
C3146 VDD.n2605 GND 0.005122f
C3147 VDD.n2606 GND 0.005122f
C3148 VDD.n2607 GND 0.006364f
C3149 VDD.n2608 GND 0.006364f
C3150 VDD.n2609 GND 0.006364f
C3151 VDD.n2610 GND 0.005122f
C3152 VDD.n2611 GND 0.005122f
C3153 VDD.n2612 GND 0.005122f
C3154 VDD.n2613 GND 0.006364f
C3155 VDD.n2614 GND 0.006364f
C3156 VDD.n2615 GND 0.006364f
C3157 VDD.n2616 GND 0.005122f
C3158 VDD.n2617 GND 0.005122f
C3159 VDD.n2618 GND 0.004251f
C3160 VDD.n2619 GND 0.014395f
C3161 VDD.n2620 GND 0.01437f
C3162 VDD.n2622 GND 0.01437f
C3163 VDD.n2623 GND 0.002331f
C3164 VDD.t58 GND 0.123904f
C3165 VDD.t56 GND 0.415248f
C3166 VDD.n2624 GND 0.086184f
C3167 VDD.t59 GND 0.090617f
C3168 VDD.n2625 GND 0.088946f
C3169 VDD.n2626 GND 0.007043f
C3170 VDD.n2627 GND 0.002792f
C3171 VDD.n2628 GND 0.005122f
C3172 VDD.n2629 GND 0.006364f
C3173 VDD.n2631 GND 0.006364f
C3174 VDD.n2632 GND 0.006364f
C3175 VDD.n2633 GND 0.005122f
C3176 VDD.n2634 GND 0.005122f
C3177 VDD.n2635 GND 0.005122f
C3178 VDD.n2636 GND 0.006364f
C3179 VDD.n2638 GND 0.006364f
C3180 VDD.n2639 GND 0.006364f
C3181 VDD.n2640 GND 0.005122f
C3182 VDD.n2641 GND 0.005122f
C3183 VDD.n2642 GND 0.005122f
C3184 VDD.n2643 GND 0.006364f
C3185 VDD.n2645 GND 0.006364f
C3186 VDD.n2646 GND 0.006364f
C3187 VDD.n2647 GND 0.005122f
C3188 VDD.n2648 GND 0.005122f
C3189 VDD.n2649 GND 0.003304f
C3190 VDD.n2650 GND 0.006364f
C3191 VDD.n2652 GND 0.006364f
C3192 VDD.n2653 GND 0.006364f
C3193 VDD.n2654 GND 0.005122f
C3194 VDD.n2655 GND 0.005122f
C3195 VDD.n2656 GND 0.005122f
C3196 VDD.n2657 GND 0.006364f
C3197 VDD.n2659 GND 0.006364f
C3198 VDD.n2660 GND 0.006364f
C3199 VDD.n2661 GND 0.005122f
C3200 VDD.n2662 GND 0.005122f
C3201 VDD.n2663 GND 0.005122f
C3202 VDD.n2664 GND 0.006364f
C3203 VDD.n2666 GND 0.006364f
C3204 VDD.n2667 GND 0.006364f
C3205 VDD.n2668 GND 0.005122f
C3206 VDD.n2669 GND 0.005122f
C3207 VDD.n2670 GND 0.005122f
C3208 VDD.n2671 GND 0.006364f
C3209 VDD.n2673 GND 0.006364f
C3210 VDD.n2674 GND 0.006364f
C3211 VDD.n2675 GND 0.003406f
C3212 VDD.t114 GND 0.123904f
C3213 VDD.t113 GND 0.415248f
C3214 VDD.n2676 GND 0.086184f
C3215 VDD.t115 GND 0.090617f
C3216 VDD.n2677 GND 0.088946f
C3217 VDD.n2678 GND 0.007043f
C3218 VDD.n2679 GND 0.002587f
C3219 VDD.n2680 GND 0.005122f
C3220 VDD.n2681 GND 0.006364f
C3221 VDD.n2683 GND 0.006364f
C3222 VDD.n2684 GND 0.006364f
C3223 VDD.n2685 GND 0.005122f
C3224 VDD.n2686 GND 0.005122f
C3225 VDD.n2687 GND 0.005122f
C3226 VDD.n2688 GND 0.006364f
C3227 VDD.n2690 GND 0.006364f
C3228 VDD.n2691 GND 0.006364f
C3229 VDD.n2692 GND 0.005122f
C3230 VDD.n2693 GND 0.005122f
C3231 VDD.n2694 GND 0.005122f
C3232 VDD.n2695 GND 0.006364f
C3233 VDD.n2697 GND 0.006364f
C3234 VDD.n2698 GND 0.006364f
C3235 VDD.n2699 GND 0.005122f
C3236 VDD.n2700 GND 0.005122f
C3237 VDD.n2701 GND 0.003509f
C3238 VDD.n2702 GND 0.006364f
C3239 VDD.n2704 GND 0.006364f
C3240 VDD.n2705 GND 0.006364f
C3241 VDD.n2706 GND 0.005045f
C3242 VDD.n2707 GND 0.005122f
C3243 VDD.n2708 GND 0.005122f
C3244 VDD.n2709 GND 0.006364f
C3245 VDD.n2711 GND 0.006364f
C3246 VDD.n2712 GND 0.006364f
C3247 VDD.n2713 GND 0.005122f
C3248 VDD.n2714 GND 0.005122f
C3249 VDD.n2715 GND 0.005122f
C3250 VDD.n2716 GND 0.006364f
C3251 VDD.n2718 GND 0.006364f
C3252 VDD.n2719 GND 0.006364f
C3253 VDD.n2720 GND 0.005122f
C3254 VDD.n2721 GND 0.005122f
C3255 VDD.n2722 GND 0.004251f
C3256 VDD.n2723 GND 0.01437f
C3257 VDD.n2724 GND 0.014395f
C3258 VDD.n2725 GND 0.004251f
C3259 VDD.n2726 GND 0.014395f
C3260 VDD.n2727 GND 0.598879f
C3261 VDD.n2728 GND 0.471559f
C3262 VDD.n2729 GND 0.471559f
C3263 VDD.n2730 GND 0.006364f
C3264 VDD.n2731 GND 0.005122f
C3265 VDD.n2732 GND 0.005122f
C3266 VDD.n2733 GND 0.005122f
C3267 VDD.n2734 GND 0.006364f
C3268 VDD.n2735 GND 0.471559f
C3269 VDD.n2736 GND 0.282935f
C3270 VDD.t57 GND 0.235779f
C3271 VDD.n2737 GND 0.424403f
C3272 VDD.n2738 GND 0.006364f
C3273 VDD.n2739 GND 0.005122f
C3274 VDD.n2740 GND 0.005122f
C3275 VDD.n2741 GND 0.005122f
C3276 VDD.n2742 GND 0.006364f
C3277 VDD.n2743 GND 0.471559f
C3278 VDD.n2744 GND 0.471559f
C3279 VDD.n2745 GND 0.471559f
C3280 VDD.n2746 GND 0.006364f
C3281 VDD.n2747 GND 0.005122f
C3282 VDD.n2748 GND 0.005122f
C3283 VDD.n2749 GND 0.005122f
C3284 VDD.n2750 GND 0.006364f
C3285 VDD.n2751 GND 0.471559f
C3286 VDD.n2752 GND 0.471559f
C3287 VDD.n2753 GND 0.471559f
C3288 VDD.n2754 GND 0.006364f
C3289 VDD.n2755 GND 0.005122f
C3290 VDD.n2756 GND 0.005122f
C3291 VDD.n2757 GND 0.005122f
C3292 VDD.n2758 GND 0.006364f
C3293 VDD.n2759 GND 0.471559f
C3294 VDD.n2760 GND 0.240495f
C3295 VDD.t0 GND 0.235779f
C3296 VDD.n2761 GND 0.466843f
C3297 VDD.n2762 GND 0.006364f
C3298 VDD.n2763 GND 0.005122f
C3299 VDD.n2764 GND 0.005122f
C3300 VDD.n2765 GND 0.005122f
C3301 VDD.n2766 GND 0.006364f
C3302 VDD.n2767 GND 0.471559f
C3303 VDD.n2768 GND 0.471559f
C3304 VDD.n2769 GND 0.471559f
C3305 VDD.n2770 GND 0.006364f
C3306 VDD.n2771 GND 0.005122f
C3307 VDD.n2772 GND 0.005122f
C3308 VDD.n2773 GND 0.005122f
C3309 VDD.n2774 GND 0.006364f
C3310 VDD.n2775 GND 0.471559f
C3311 VDD.n2776 GND 0.471559f
C3312 VDD.t2 GND 0.471559f
C3313 VDD.n2777 GND 0.006364f
C3314 VDD.n2778 GND 0.005122f
C3315 VDD.n2779 GND 0.14125f
C3316 VDD.n2780 GND 1.88697f
C3317 a_n2500_9133.n0 GND 4.54423f
C3318 a_n2500_9133.n1 GND 10.5214f
C3319 a_n2500_9133.t0 GND 0.103322p
C3320 a_n2500_9133.t2 GND 0.477832f
C3321 a_n2500_9133.t6 GND 0.173091f
C3322 a_n2500_9133.t7 GND 0.034646f
C3323 a_n2500_9133.t4 GND 0.034646f
C3324 a_n2500_9133.n2 GND 0.114733f
C3325 a_n2500_9133.t1 GND 0.169644f
C3326 a_n2500_9133.t5 GND 0.169644f
C3327 a_n2500_9133.t3 GND 0.034646f
C3328 a_n2500_9133.t9 GND 0.034646f
C3329 a_n2500_9133.n3 GND 0.114733f
C3330 a_n2500_9133.t8 GND 0.169644f
C3331 a_n2500_9133.t10 GND 0.2841f
C3332 a_n6918_10482.n0 GND 0.472283f
C3333 a_n6918_10482.n1 GND 3.94927f
C3334 a_n6918_10482.n2 GND 0.508019f
C3335 a_n6918_10482.n3 GND 6.22833f
C3336 a_n6918_10482.n4 GND 0.508017f
C3337 a_n6918_10482.n5 GND 0.508017f
C3338 a_n6918_10482.n6 GND 0.538273f
C3339 a_n6918_10482.n7 GND 7.99396f
C3340 a_n6918_10482.n8 GND 2.24933f
C3341 a_n6918_10482.n9 GND 5.36075f
C3342 a_n6918_10482.n10 GND 0.490955f
C3343 a_n6918_10482.n11 GND 0.490955f
C3344 a_n6918_10482.n12 GND 7.747089f
C3345 a_n6918_10482.n13 GND 0.490958f
C3346 a_n6918_10482.t5 GND 3.04653f
C3347 a_n6918_10482.t0 GND 1.33586f
C3348 a_n6918_10482.t3 GND 0.57592f
C3349 a_n6918_10482.t19 GND 1.30261f
C3350 a_n6918_10482.t7 GND 1.26602f
C3351 a_n6918_10482.t8 GND 1.30261f
C3352 a_n6918_10482.t22 GND 0.822199f
C3353 a_n6918_10482.n14 GND 0.703616f
C3354 a_n6918_10482.t18 GND 1.30261f
C3355 a_n6918_10482.t23 GND 1.23475f
C3356 a_n6918_10482.t6 GND 1.30261f
C3357 a_n6918_10482.t16 GND 0.822199f
C3358 a_n6918_10482.n15 GND 0.703616f
C3359 a_n6918_10482.t2 GND 1.33586f
C3360 a_n6918_10482.n16 GND 2.32531f
C3361 a_n6918_10482.t12 GND 1.33586f
C3362 a_n6918_10482.n17 GND 2.49066f
C3363 a_n6918_10482.t1 GND 0.539599f
C3364 a_n6918_10482.t15 GND 1.30261f
C3365 a_n6918_10482.t11 GND 1.26603f
C3366 a_n6918_10482.t10 GND 1.30261f
C3367 a_n6918_10482.t17 GND 1.05456f
C3368 a_n6918_10482.t14 GND 1.30261f
C3369 a_n6918_10482.t20 GND 1.26603f
C3370 a_n6918_10482.t9 GND 1.30261f
C3371 a_n6918_10482.t13 GND 0.822199f
C3372 a_n6918_10482.n18 GND 0.703619f
C3373 a_n6918_10482.t21 GND 1.33586f
C3374 a_n6918_10482.n19 GND 10.1361f
C3375 a_n6918_10482.t4 GND 1.82049f
C3376 a_n2675_n4106.n0 GND 1.79164f
C3377 a_n2675_n4106.t5 GND 0.796979f
C3378 a_n2675_n4106.t3 GND 0.671924f
C3379 a_n2675_n4106.n1 GND 1.08328f
C3380 a_n2675_n4106.t1 GND 0.671927f
C3381 a_n2675_n4106.n2 GND 1.39583f
C3382 a_n2675_n4106.n3 GND 0.619026f
C3383 a_n2675_n4106.t0 GND 0.671926f
C3384 a_n2675_n4106.n4 GND 1.20491f
C3385 a_n2675_n4106.t2 GND 0.671926f
C3386 a_n2675_n4106.n5 GND 0.924707f
C3387 a_n2675_n4106.n6 GND 0.517142f
C3388 a_n2675_n4106.t4 GND 0.794958f
C3389 a_n2675_n4106.n7 GND 1.39646f
C3390 a_n2675_n4106.t8 GND 0.794958f
C3391 a_n2675_n4106.n8 GND 1.05125f
C3392 a_n2675_n4106.t6 GND 0.794958f
C3393 a_n2675_n4106.n9 GND 1.05125f
C3394 a_n2675_n4106.t7 GND 0.794958f
C3395 DIFFPAIR_BIAS.t10 GND 0.10454f
C3396 DIFFPAIR_BIAS.t14 GND 0.105557f
C3397 DIFFPAIR_BIAS.n0 GND 0.131947f
C3398 DIFFPAIR_BIAS.t5 GND 0.075148f
C3399 DIFFPAIR_BIAS.t3 GND 0.074193f
C3400 DIFFPAIR_BIAS.n1 GND 0.232704f
C3401 DIFFPAIR_BIAS.t7 GND 0.074193f
C3402 DIFFPAIR_BIAS.n2 GND 0.122823f
C3403 DIFFPAIR_BIAS.t9 GND 0.074193f
C3404 DIFFPAIR_BIAS.n3 GND 0.122823f
C3405 DIFFPAIR_BIAS.t1 GND 0.074193f
C3406 DIFFPAIR_BIAS.n4 GND 0.146908f
C3407 DIFFPAIR_BIAS.t0 GND 0.099056f
C3408 DIFFPAIR_BIAS.t8 GND 0.099056f
C3409 DIFFPAIR_BIAS.t6 GND 0.099056f
C3410 DIFFPAIR_BIAS.t2 GND 0.099056f
C3411 DIFFPAIR_BIAS.t4 GND 0.10018f
C3412 DIFFPAIR_BIAS.n5 GND 0.125716f
C3413 DIFFPAIR_BIAS.n6 GND 0.068742f
C3414 DIFFPAIR_BIAS.n7 GND 0.068742f
C3415 DIFFPAIR_BIAS.n8 GND 0.07449f
C3416 DIFFPAIR_BIAS.n9 GND 0.149198f
C3417 DIFFPAIR_BIAS.t13 GND 0.10454f
C3418 DIFFPAIR_BIAS.n10 GND 0.062199f
C3419 DIFFPAIR_BIAS.t11 GND 0.10454f
C3420 DIFFPAIR_BIAS.n11 GND 0.067027f
C3421 DIFFPAIR_BIAS.t12 GND 0.10454f
C3422 DIFFPAIR_BIAS.n12 GND 0.053964f
C3423 DIFFPAIR_BIAS.n13 GND 0.039084f
.ends

