* NGSPICE file created from diff_pair_sample_1350.ext - technology: sky130A

.subckt diff_pair_sample_1350 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=0 ps=0 w=15.94 l=3.17
X1 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6301 pd=16.27 as=6.2166 ps=32.66 w=15.94 l=3.17
X2 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6301 pd=16.27 as=6.2166 ps=32.66 w=15.94 l=3.17
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=0 ps=0 w=15.94 l=3.17
X4 VTAIL.t4 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=2.6301 ps=16.27 w=15.94 l=3.17
X5 VDD1.t1 VP.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6301 pd=16.27 as=6.2166 ps=32.66 w=15.94 l=3.17
X6 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=2.6301 ps=16.27 w=15.94 l=3.17
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=0 ps=0 w=15.94 l=3.17
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6301 pd=16.27 as=6.2166 ps=32.66 w=15.94 l=3.17
X9 VTAIL.t6 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=2.6301 ps=16.27 w=15.94 l=3.17
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=0 ps=0 w=15.94 l=3.17
X11 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2166 pd=32.66 as=2.6301 ps=16.27 w=15.94 l=3.17
R0 B.n902 B.n901 585
R1 B.n363 B.n131 585
R2 B.n362 B.n361 585
R3 B.n360 B.n359 585
R4 B.n358 B.n357 585
R5 B.n356 B.n355 585
R6 B.n354 B.n353 585
R7 B.n352 B.n351 585
R8 B.n350 B.n349 585
R9 B.n348 B.n347 585
R10 B.n346 B.n345 585
R11 B.n344 B.n343 585
R12 B.n342 B.n341 585
R13 B.n340 B.n339 585
R14 B.n338 B.n337 585
R15 B.n336 B.n335 585
R16 B.n334 B.n333 585
R17 B.n332 B.n331 585
R18 B.n330 B.n329 585
R19 B.n328 B.n327 585
R20 B.n326 B.n325 585
R21 B.n324 B.n323 585
R22 B.n322 B.n321 585
R23 B.n320 B.n319 585
R24 B.n318 B.n317 585
R25 B.n316 B.n315 585
R26 B.n314 B.n313 585
R27 B.n312 B.n311 585
R28 B.n310 B.n309 585
R29 B.n308 B.n307 585
R30 B.n306 B.n305 585
R31 B.n304 B.n303 585
R32 B.n302 B.n301 585
R33 B.n300 B.n299 585
R34 B.n298 B.n297 585
R35 B.n296 B.n295 585
R36 B.n294 B.n293 585
R37 B.n292 B.n291 585
R38 B.n290 B.n289 585
R39 B.n288 B.n287 585
R40 B.n286 B.n285 585
R41 B.n284 B.n283 585
R42 B.n282 B.n281 585
R43 B.n280 B.n279 585
R44 B.n278 B.n277 585
R45 B.n276 B.n275 585
R46 B.n274 B.n273 585
R47 B.n272 B.n271 585
R48 B.n270 B.n269 585
R49 B.n268 B.n267 585
R50 B.n266 B.n265 585
R51 B.n264 B.n263 585
R52 B.n262 B.n261 585
R53 B.n259 B.n258 585
R54 B.n257 B.n256 585
R55 B.n255 B.n254 585
R56 B.n253 B.n252 585
R57 B.n251 B.n250 585
R58 B.n249 B.n248 585
R59 B.n247 B.n246 585
R60 B.n245 B.n244 585
R61 B.n243 B.n242 585
R62 B.n241 B.n240 585
R63 B.n238 B.n237 585
R64 B.n236 B.n235 585
R65 B.n234 B.n233 585
R66 B.n232 B.n231 585
R67 B.n230 B.n229 585
R68 B.n228 B.n227 585
R69 B.n226 B.n225 585
R70 B.n224 B.n223 585
R71 B.n222 B.n221 585
R72 B.n220 B.n219 585
R73 B.n218 B.n217 585
R74 B.n216 B.n215 585
R75 B.n214 B.n213 585
R76 B.n212 B.n211 585
R77 B.n210 B.n209 585
R78 B.n208 B.n207 585
R79 B.n206 B.n205 585
R80 B.n204 B.n203 585
R81 B.n202 B.n201 585
R82 B.n200 B.n199 585
R83 B.n198 B.n197 585
R84 B.n196 B.n195 585
R85 B.n194 B.n193 585
R86 B.n192 B.n191 585
R87 B.n190 B.n189 585
R88 B.n188 B.n187 585
R89 B.n186 B.n185 585
R90 B.n184 B.n183 585
R91 B.n182 B.n181 585
R92 B.n180 B.n179 585
R93 B.n178 B.n177 585
R94 B.n176 B.n175 585
R95 B.n174 B.n173 585
R96 B.n172 B.n171 585
R97 B.n170 B.n169 585
R98 B.n168 B.n167 585
R99 B.n166 B.n165 585
R100 B.n164 B.n163 585
R101 B.n162 B.n161 585
R102 B.n160 B.n159 585
R103 B.n158 B.n157 585
R104 B.n156 B.n155 585
R105 B.n154 B.n153 585
R106 B.n152 B.n151 585
R107 B.n150 B.n149 585
R108 B.n148 B.n147 585
R109 B.n146 B.n145 585
R110 B.n144 B.n143 585
R111 B.n142 B.n141 585
R112 B.n140 B.n139 585
R113 B.n138 B.n137 585
R114 B.n74 B.n73 585
R115 B.n907 B.n906 585
R116 B.n900 B.n132 585
R117 B.n132 B.n71 585
R118 B.n899 B.n70 585
R119 B.n911 B.n70 585
R120 B.n898 B.n69 585
R121 B.n912 B.n69 585
R122 B.n897 B.n68 585
R123 B.n913 B.n68 585
R124 B.n896 B.n895 585
R125 B.n895 B.n64 585
R126 B.n894 B.n63 585
R127 B.n919 B.n63 585
R128 B.n893 B.n62 585
R129 B.n920 B.n62 585
R130 B.n892 B.n61 585
R131 B.n921 B.n61 585
R132 B.n891 B.n890 585
R133 B.n890 B.n60 585
R134 B.n889 B.n56 585
R135 B.n927 B.n56 585
R136 B.n888 B.n55 585
R137 B.n928 B.n55 585
R138 B.n887 B.n54 585
R139 B.n929 B.n54 585
R140 B.n886 B.n885 585
R141 B.n885 B.n50 585
R142 B.n884 B.n49 585
R143 B.n935 B.n49 585
R144 B.n883 B.n48 585
R145 B.n936 B.n48 585
R146 B.n882 B.n47 585
R147 B.n937 B.n47 585
R148 B.n881 B.n880 585
R149 B.n880 B.n43 585
R150 B.n879 B.n42 585
R151 B.n943 B.n42 585
R152 B.n878 B.n41 585
R153 B.n944 B.n41 585
R154 B.n877 B.n40 585
R155 B.n945 B.n40 585
R156 B.n876 B.n875 585
R157 B.n875 B.n36 585
R158 B.n874 B.n35 585
R159 B.n951 B.n35 585
R160 B.n873 B.n34 585
R161 B.n952 B.n34 585
R162 B.n872 B.n33 585
R163 B.n953 B.n33 585
R164 B.n871 B.n870 585
R165 B.n870 B.n29 585
R166 B.n869 B.n28 585
R167 B.n959 B.n28 585
R168 B.n868 B.n27 585
R169 B.n960 B.n27 585
R170 B.n867 B.n26 585
R171 B.n961 B.n26 585
R172 B.n866 B.n865 585
R173 B.n865 B.n22 585
R174 B.n864 B.n21 585
R175 B.n967 B.n21 585
R176 B.n863 B.n20 585
R177 B.n968 B.n20 585
R178 B.n862 B.n19 585
R179 B.n969 B.n19 585
R180 B.n861 B.n860 585
R181 B.n860 B.n18 585
R182 B.n859 B.n14 585
R183 B.n975 B.n14 585
R184 B.n858 B.n13 585
R185 B.n976 B.n13 585
R186 B.n857 B.n12 585
R187 B.n977 B.n12 585
R188 B.n856 B.n855 585
R189 B.n855 B.n8 585
R190 B.n854 B.n7 585
R191 B.n983 B.n7 585
R192 B.n853 B.n6 585
R193 B.n984 B.n6 585
R194 B.n852 B.n5 585
R195 B.n985 B.n5 585
R196 B.n851 B.n850 585
R197 B.n850 B.n4 585
R198 B.n849 B.n364 585
R199 B.n849 B.n848 585
R200 B.n839 B.n365 585
R201 B.n366 B.n365 585
R202 B.n841 B.n840 585
R203 B.n842 B.n841 585
R204 B.n838 B.n371 585
R205 B.n371 B.n370 585
R206 B.n837 B.n836 585
R207 B.n836 B.n835 585
R208 B.n373 B.n372 585
R209 B.n828 B.n373 585
R210 B.n827 B.n826 585
R211 B.n829 B.n827 585
R212 B.n825 B.n378 585
R213 B.n378 B.n377 585
R214 B.n824 B.n823 585
R215 B.n823 B.n822 585
R216 B.n380 B.n379 585
R217 B.n381 B.n380 585
R218 B.n815 B.n814 585
R219 B.n816 B.n815 585
R220 B.n813 B.n386 585
R221 B.n386 B.n385 585
R222 B.n812 B.n811 585
R223 B.n811 B.n810 585
R224 B.n388 B.n387 585
R225 B.n389 B.n388 585
R226 B.n803 B.n802 585
R227 B.n804 B.n803 585
R228 B.n801 B.n394 585
R229 B.n394 B.n393 585
R230 B.n800 B.n799 585
R231 B.n799 B.n798 585
R232 B.n396 B.n395 585
R233 B.n397 B.n396 585
R234 B.n791 B.n790 585
R235 B.n792 B.n791 585
R236 B.n789 B.n402 585
R237 B.n402 B.n401 585
R238 B.n788 B.n787 585
R239 B.n787 B.n786 585
R240 B.n404 B.n403 585
R241 B.n405 B.n404 585
R242 B.n779 B.n778 585
R243 B.n780 B.n779 585
R244 B.n777 B.n410 585
R245 B.n410 B.n409 585
R246 B.n776 B.n775 585
R247 B.n775 B.n774 585
R248 B.n412 B.n411 585
R249 B.n413 B.n412 585
R250 B.n767 B.n766 585
R251 B.n768 B.n767 585
R252 B.n765 B.n418 585
R253 B.n418 B.n417 585
R254 B.n764 B.n763 585
R255 B.n763 B.n762 585
R256 B.n420 B.n419 585
R257 B.n755 B.n420 585
R258 B.n754 B.n753 585
R259 B.n756 B.n754 585
R260 B.n752 B.n425 585
R261 B.n425 B.n424 585
R262 B.n751 B.n750 585
R263 B.n750 B.n749 585
R264 B.n427 B.n426 585
R265 B.n428 B.n427 585
R266 B.n742 B.n741 585
R267 B.n743 B.n742 585
R268 B.n740 B.n433 585
R269 B.n433 B.n432 585
R270 B.n739 B.n738 585
R271 B.n738 B.n737 585
R272 B.n435 B.n434 585
R273 B.n436 B.n435 585
R274 B.n733 B.n732 585
R275 B.n439 B.n438 585
R276 B.n729 B.n728 585
R277 B.n730 B.n729 585
R278 B.n727 B.n497 585
R279 B.n726 B.n725 585
R280 B.n724 B.n723 585
R281 B.n722 B.n721 585
R282 B.n720 B.n719 585
R283 B.n718 B.n717 585
R284 B.n716 B.n715 585
R285 B.n714 B.n713 585
R286 B.n712 B.n711 585
R287 B.n710 B.n709 585
R288 B.n708 B.n707 585
R289 B.n706 B.n705 585
R290 B.n704 B.n703 585
R291 B.n702 B.n701 585
R292 B.n700 B.n699 585
R293 B.n698 B.n697 585
R294 B.n696 B.n695 585
R295 B.n694 B.n693 585
R296 B.n692 B.n691 585
R297 B.n690 B.n689 585
R298 B.n688 B.n687 585
R299 B.n686 B.n685 585
R300 B.n684 B.n683 585
R301 B.n682 B.n681 585
R302 B.n680 B.n679 585
R303 B.n678 B.n677 585
R304 B.n676 B.n675 585
R305 B.n674 B.n673 585
R306 B.n672 B.n671 585
R307 B.n670 B.n669 585
R308 B.n668 B.n667 585
R309 B.n666 B.n665 585
R310 B.n664 B.n663 585
R311 B.n662 B.n661 585
R312 B.n660 B.n659 585
R313 B.n658 B.n657 585
R314 B.n656 B.n655 585
R315 B.n654 B.n653 585
R316 B.n652 B.n651 585
R317 B.n650 B.n649 585
R318 B.n648 B.n647 585
R319 B.n646 B.n645 585
R320 B.n644 B.n643 585
R321 B.n642 B.n641 585
R322 B.n640 B.n639 585
R323 B.n638 B.n637 585
R324 B.n636 B.n635 585
R325 B.n634 B.n633 585
R326 B.n632 B.n631 585
R327 B.n630 B.n629 585
R328 B.n628 B.n627 585
R329 B.n626 B.n625 585
R330 B.n624 B.n623 585
R331 B.n622 B.n621 585
R332 B.n620 B.n619 585
R333 B.n618 B.n617 585
R334 B.n616 B.n615 585
R335 B.n614 B.n613 585
R336 B.n612 B.n611 585
R337 B.n610 B.n609 585
R338 B.n608 B.n607 585
R339 B.n606 B.n605 585
R340 B.n604 B.n603 585
R341 B.n602 B.n601 585
R342 B.n600 B.n599 585
R343 B.n598 B.n597 585
R344 B.n596 B.n595 585
R345 B.n594 B.n593 585
R346 B.n592 B.n591 585
R347 B.n590 B.n589 585
R348 B.n588 B.n587 585
R349 B.n586 B.n585 585
R350 B.n584 B.n583 585
R351 B.n582 B.n581 585
R352 B.n580 B.n579 585
R353 B.n578 B.n577 585
R354 B.n576 B.n575 585
R355 B.n574 B.n573 585
R356 B.n572 B.n571 585
R357 B.n570 B.n569 585
R358 B.n568 B.n567 585
R359 B.n566 B.n565 585
R360 B.n564 B.n563 585
R361 B.n562 B.n561 585
R362 B.n560 B.n559 585
R363 B.n558 B.n557 585
R364 B.n556 B.n555 585
R365 B.n554 B.n553 585
R366 B.n552 B.n551 585
R367 B.n550 B.n549 585
R368 B.n548 B.n547 585
R369 B.n546 B.n545 585
R370 B.n544 B.n543 585
R371 B.n542 B.n541 585
R372 B.n540 B.n539 585
R373 B.n538 B.n537 585
R374 B.n536 B.n535 585
R375 B.n534 B.n533 585
R376 B.n532 B.n531 585
R377 B.n530 B.n529 585
R378 B.n528 B.n527 585
R379 B.n526 B.n525 585
R380 B.n524 B.n523 585
R381 B.n522 B.n521 585
R382 B.n520 B.n519 585
R383 B.n518 B.n517 585
R384 B.n516 B.n515 585
R385 B.n514 B.n513 585
R386 B.n512 B.n511 585
R387 B.n510 B.n509 585
R388 B.n508 B.n507 585
R389 B.n506 B.n505 585
R390 B.n504 B.n496 585
R391 B.n730 B.n496 585
R392 B.n734 B.n437 585
R393 B.n437 B.n436 585
R394 B.n736 B.n735 585
R395 B.n737 B.n736 585
R396 B.n431 B.n430 585
R397 B.n432 B.n431 585
R398 B.n745 B.n744 585
R399 B.n744 B.n743 585
R400 B.n746 B.n429 585
R401 B.n429 B.n428 585
R402 B.n748 B.n747 585
R403 B.n749 B.n748 585
R404 B.n423 B.n422 585
R405 B.n424 B.n423 585
R406 B.n758 B.n757 585
R407 B.n757 B.n756 585
R408 B.n759 B.n421 585
R409 B.n755 B.n421 585
R410 B.n761 B.n760 585
R411 B.n762 B.n761 585
R412 B.n416 B.n415 585
R413 B.n417 B.n416 585
R414 B.n770 B.n769 585
R415 B.n769 B.n768 585
R416 B.n771 B.n414 585
R417 B.n414 B.n413 585
R418 B.n773 B.n772 585
R419 B.n774 B.n773 585
R420 B.n408 B.n407 585
R421 B.n409 B.n408 585
R422 B.n782 B.n781 585
R423 B.n781 B.n780 585
R424 B.n783 B.n406 585
R425 B.n406 B.n405 585
R426 B.n785 B.n784 585
R427 B.n786 B.n785 585
R428 B.n400 B.n399 585
R429 B.n401 B.n400 585
R430 B.n794 B.n793 585
R431 B.n793 B.n792 585
R432 B.n795 B.n398 585
R433 B.n398 B.n397 585
R434 B.n797 B.n796 585
R435 B.n798 B.n797 585
R436 B.n392 B.n391 585
R437 B.n393 B.n392 585
R438 B.n806 B.n805 585
R439 B.n805 B.n804 585
R440 B.n807 B.n390 585
R441 B.n390 B.n389 585
R442 B.n809 B.n808 585
R443 B.n810 B.n809 585
R444 B.n384 B.n383 585
R445 B.n385 B.n384 585
R446 B.n818 B.n817 585
R447 B.n817 B.n816 585
R448 B.n819 B.n382 585
R449 B.n382 B.n381 585
R450 B.n821 B.n820 585
R451 B.n822 B.n821 585
R452 B.n376 B.n375 585
R453 B.n377 B.n376 585
R454 B.n831 B.n830 585
R455 B.n830 B.n829 585
R456 B.n832 B.n374 585
R457 B.n828 B.n374 585
R458 B.n834 B.n833 585
R459 B.n835 B.n834 585
R460 B.n369 B.n368 585
R461 B.n370 B.n369 585
R462 B.n844 B.n843 585
R463 B.n843 B.n842 585
R464 B.n845 B.n367 585
R465 B.n367 B.n366 585
R466 B.n847 B.n846 585
R467 B.n848 B.n847 585
R468 B.n2 B.n0 585
R469 B.n4 B.n2 585
R470 B.n3 B.n1 585
R471 B.n984 B.n3 585
R472 B.n982 B.n981 585
R473 B.n983 B.n982 585
R474 B.n980 B.n9 585
R475 B.n9 B.n8 585
R476 B.n979 B.n978 585
R477 B.n978 B.n977 585
R478 B.n11 B.n10 585
R479 B.n976 B.n11 585
R480 B.n974 B.n973 585
R481 B.n975 B.n974 585
R482 B.n972 B.n15 585
R483 B.n18 B.n15 585
R484 B.n971 B.n970 585
R485 B.n970 B.n969 585
R486 B.n17 B.n16 585
R487 B.n968 B.n17 585
R488 B.n966 B.n965 585
R489 B.n967 B.n966 585
R490 B.n964 B.n23 585
R491 B.n23 B.n22 585
R492 B.n963 B.n962 585
R493 B.n962 B.n961 585
R494 B.n25 B.n24 585
R495 B.n960 B.n25 585
R496 B.n958 B.n957 585
R497 B.n959 B.n958 585
R498 B.n956 B.n30 585
R499 B.n30 B.n29 585
R500 B.n955 B.n954 585
R501 B.n954 B.n953 585
R502 B.n32 B.n31 585
R503 B.n952 B.n32 585
R504 B.n950 B.n949 585
R505 B.n951 B.n950 585
R506 B.n948 B.n37 585
R507 B.n37 B.n36 585
R508 B.n947 B.n946 585
R509 B.n946 B.n945 585
R510 B.n39 B.n38 585
R511 B.n944 B.n39 585
R512 B.n942 B.n941 585
R513 B.n943 B.n942 585
R514 B.n940 B.n44 585
R515 B.n44 B.n43 585
R516 B.n939 B.n938 585
R517 B.n938 B.n937 585
R518 B.n46 B.n45 585
R519 B.n936 B.n46 585
R520 B.n934 B.n933 585
R521 B.n935 B.n934 585
R522 B.n932 B.n51 585
R523 B.n51 B.n50 585
R524 B.n931 B.n930 585
R525 B.n930 B.n929 585
R526 B.n53 B.n52 585
R527 B.n928 B.n53 585
R528 B.n926 B.n925 585
R529 B.n927 B.n926 585
R530 B.n924 B.n57 585
R531 B.n60 B.n57 585
R532 B.n923 B.n922 585
R533 B.n922 B.n921 585
R534 B.n59 B.n58 585
R535 B.n920 B.n59 585
R536 B.n918 B.n917 585
R537 B.n919 B.n918 585
R538 B.n916 B.n65 585
R539 B.n65 B.n64 585
R540 B.n915 B.n914 585
R541 B.n914 B.n913 585
R542 B.n67 B.n66 585
R543 B.n912 B.n67 585
R544 B.n910 B.n909 585
R545 B.n911 B.n910 585
R546 B.n908 B.n72 585
R547 B.n72 B.n71 585
R548 B.n987 B.n986 585
R549 B.n986 B.n985 585
R550 B.n732 B.n437 497.305
R551 B.n906 B.n72 497.305
R552 B.n496 B.n435 497.305
R553 B.n902 B.n132 497.305
R554 B.n501 B.t8 329.955
R555 B.n498 B.t15 329.955
R556 B.n135 B.t4 329.955
R557 B.n133 B.t12 329.955
R558 B.n904 B.n903 256.663
R559 B.n904 B.n130 256.663
R560 B.n904 B.n129 256.663
R561 B.n904 B.n128 256.663
R562 B.n904 B.n127 256.663
R563 B.n904 B.n126 256.663
R564 B.n904 B.n125 256.663
R565 B.n904 B.n124 256.663
R566 B.n904 B.n123 256.663
R567 B.n904 B.n122 256.663
R568 B.n904 B.n121 256.663
R569 B.n904 B.n120 256.663
R570 B.n904 B.n119 256.663
R571 B.n904 B.n118 256.663
R572 B.n904 B.n117 256.663
R573 B.n904 B.n116 256.663
R574 B.n904 B.n115 256.663
R575 B.n904 B.n114 256.663
R576 B.n904 B.n113 256.663
R577 B.n904 B.n112 256.663
R578 B.n904 B.n111 256.663
R579 B.n904 B.n110 256.663
R580 B.n904 B.n109 256.663
R581 B.n904 B.n108 256.663
R582 B.n904 B.n107 256.663
R583 B.n904 B.n106 256.663
R584 B.n904 B.n105 256.663
R585 B.n904 B.n104 256.663
R586 B.n904 B.n103 256.663
R587 B.n904 B.n102 256.663
R588 B.n904 B.n101 256.663
R589 B.n904 B.n100 256.663
R590 B.n904 B.n99 256.663
R591 B.n904 B.n98 256.663
R592 B.n904 B.n97 256.663
R593 B.n904 B.n96 256.663
R594 B.n904 B.n95 256.663
R595 B.n904 B.n94 256.663
R596 B.n904 B.n93 256.663
R597 B.n904 B.n92 256.663
R598 B.n904 B.n91 256.663
R599 B.n904 B.n90 256.663
R600 B.n904 B.n89 256.663
R601 B.n904 B.n88 256.663
R602 B.n904 B.n87 256.663
R603 B.n904 B.n86 256.663
R604 B.n904 B.n85 256.663
R605 B.n904 B.n84 256.663
R606 B.n904 B.n83 256.663
R607 B.n904 B.n82 256.663
R608 B.n904 B.n81 256.663
R609 B.n904 B.n80 256.663
R610 B.n904 B.n79 256.663
R611 B.n904 B.n78 256.663
R612 B.n904 B.n77 256.663
R613 B.n904 B.n76 256.663
R614 B.n904 B.n75 256.663
R615 B.n905 B.n904 256.663
R616 B.n731 B.n730 256.663
R617 B.n730 B.n440 256.663
R618 B.n730 B.n441 256.663
R619 B.n730 B.n442 256.663
R620 B.n730 B.n443 256.663
R621 B.n730 B.n444 256.663
R622 B.n730 B.n445 256.663
R623 B.n730 B.n446 256.663
R624 B.n730 B.n447 256.663
R625 B.n730 B.n448 256.663
R626 B.n730 B.n449 256.663
R627 B.n730 B.n450 256.663
R628 B.n730 B.n451 256.663
R629 B.n730 B.n452 256.663
R630 B.n730 B.n453 256.663
R631 B.n730 B.n454 256.663
R632 B.n730 B.n455 256.663
R633 B.n730 B.n456 256.663
R634 B.n730 B.n457 256.663
R635 B.n730 B.n458 256.663
R636 B.n730 B.n459 256.663
R637 B.n730 B.n460 256.663
R638 B.n730 B.n461 256.663
R639 B.n730 B.n462 256.663
R640 B.n730 B.n463 256.663
R641 B.n730 B.n464 256.663
R642 B.n730 B.n465 256.663
R643 B.n730 B.n466 256.663
R644 B.n730 B.n467 256.663
R645 B.n730 B.n468 256.663
R646 B.n730 B.n469 256.663
R647 B.n730 B.n470 256.663
R648 B.n730 B.n471 256.663
R649 B.n730 B.n472 256.663
R650 B.n730 B.n473 256.663
R651 B.n730 B.n474 256.663
R652 B.n730 B.n475 256.663
R653 B.n730 B.n476 256.663
R654 B.n730 B.n477 256.663
R655 B.n730 B.n478 256.663
R656 B.n730 B.n479 256.663
R657 B.n730 B.n480 256.663
R658 B.n730 B.n481 256.663
R659 B.n730 B.n482 256.663
R660 B.n730 B.n483 256.663
R661 B.n730 B.n484 256.663
R662 B.n730 B.n485 256.663
R663 B.n730 B.n486 256.663
R664 B.n730 B.n487 256.663
R665 B.n730 B.n488 256.663
R666 B.n730 B.n489 256.663
R667 B.n730 B.n490 256.663
R668 B.n730 B.n491 256.663
R669 B.n730 B.n492 256.663
R670 B.n730 B.n493 256.663
R671 B.n730 B.n494 256.663
R672 B.n730 B.n495 256.663
R673 B.n736 B.n437 163.367
R674 B.n736 B.n431 163.367
R675 B.n744 B.n431 163.367
R676 B.n744 B.n429 163.367
R677 B.n748 B.n429 163.367
R678 B.n748 B.n423 163.367
R679 B.n757 B.n423 163.367
R680 B.n757 B.n421 163.367
R681 B.n761 B.n421 163.367
R682 B.n761 B.n416 163.367
R683 B.n769 B.n416 163.367
R684 B.n769 B.n414 163.367
R685 B.n773 B.n414 163.367
R686 B.n773 B.n408 163.367
R687 B.n781 B.n408 163.367
R688 B.n781 B.n406 163.367
R689 B.n785 B.n406 163.367
R690 B.n785 B.n400 163.367
R691 B.n793 B.n400 163.367
R692 B.n793 B.n398 163.367
R693 B.n797 B.n398 163.367
R694 B.n797 B.n392 163.367
R695 B.n805 B.n392 163.367
R696 B.n805 B.n390 163.367
R697 B.n809 B.n390 163.367
R698 B.n809 B.n384 163.367
R699 B.n817 B.n384 163.367
R700 B.n817 B.n382 163.367
R701 B.n821 B.n382 163.367
R702 B.n821 B.n376 163.367
R703 B.n830 B.n376 163.367
R704 B.n830 B.n374 163.367
R705 B.n834 B.n374 163.367
R706 B.n834 B.n369 163.367
R707 B.n843 B.n369 163.367
R708 B.n843 B.n367 163.367
R709 B.n847 B.n367 163.367
R710 B.n847 B.n2 163.367
R711 B.n986 B.n2 163.367
R712 B.n986 B.n3 163.367
R713 B.n982 B.n3 163.367
R714 B.n982 B.n9 163.367
R715 B.n978 B.n9 163.367
R716 B.n978 B.n11 163.367
R717 B.n974 B.n11 163.367
R718 B.n974 B.n15 163.367
R719 B.n970 B.n15 163.367
R720 B.n970 B.n17 163.367
R721 B.n966 B.n17 163.367
R722 B.n966 B.n23 163.367
R723 B.n962 B.n23 163.367
R724 B.n962 B.n25 163.367
R725 B.n958 B.n25 163.367
R726 B.n958 B.n30 163.367
R727 B.n954 B.n30 163.367
R728 B.n954 B.n32 163.367
R729 B.n950 B.n32 163.367
R730 B.n950 B.n37 163.367
R731 B.n946 B.n37 163.367
R732 B.n946 B.n39 163.367
R733 B.n942 B.n39 163.367
R734 B.n942 B.n44 163.367
R735 B.n938 B.n44 163.367
R736 B.n938 B.n46 163.367
R737 B.n934 B.n46 163.367
R738 B.n934 B.n51 163.367
R739 B.n930 B.n51 163.367
R740 B.n930 B.n53 163.367
R741 B.n926 B.n53 163.367
R742 B.n926 B.n57 163.367
R743 B.n922 B.n57 163.367
R744 B.n922 B.n59 163.367
R745 B.n918 B.n59 163.367
R746 B.n918 B.n65 163.367
R747 B.n914 B.n65 163.367
R748 B.n914 B.n67 163.367
R749 B.n910 B.n67 163.367
R750 B.n910 B.n72 163.367
R751 B.n729 B.n439 163.367
R752 B.n729 B.n497 163.367
R753 B.n725 B.n724 163.367
R754 B.n721 B.n720 163.367
R755 B.n717 B.n716 163.367
R756 B.n713 B.n712 163.367
R757 B.n709 B.n708 163.367
R758 B.n705 B.n704 163.367
R759 B.n701 B.n700 163.367
R760 B.n697 B.n696 163.367
R761 B.n693 B.n692 163.367
R762 B.n689 B.n688 163.367
R763 B.n685 B.n684 163.367
R764 B.n681 B.n680 163.367
R765 B.n677 B.n676 163.367
R766 B.n673 B.n672 163.367
R767 B.n669 B.n668 163.367
R768 B.n665 B.n664 163.367
R769 B.n661 B.n660 163.367
R770 B.n657 B.n656 163.367
R771 B.n653 B.n652 163.367
R772 B.n649 B.n648 163.367
R773 B.n645 B.n644 163.367
R774 B.n641 B.n640 163.367
R775 B.n637 B.n636 163.367
R776 B.n633 B.n632 163.367
R777 B.n629 B.n628 163.367
R778 B.n625 B.n624 163.367
R779 B.n621 B.n620 163.367
R780 B.n617 B.n616 163.367
R781 B.n613 B.n612 163.367
R782 B.n609 B.n608 163.367
R783 B.n605 B.n604 163.367
R784 B.n601 B.n600 163.367
R785 B.n597 B.n596 163.367
R786 B.n593 B.n592 163.367
R787 B.n589 B.n588 163.367
R788 B.n585 B.n584 163.367
R789 B.n581 B.n580 163.367
R790 B.n577 B.n576 163.367
R791 B.n573 B.n572 163.367
R792 B.n569 B.n568 163.367
R793 B.n565 B.n564 163.367
R794 B.n561 B.n560 163.367
R795 B.n557 B.n556 163.367
R796 B.n553 B.n552 163.367
R797 B.n549 B.n548 163.367
R798 B.n545 B.n544 163.367
R799 B.n541 B.n540 163.367
R800 B.n537 B.n536 163.367
R801 B.n533 B.n532 163.367
R802 B.n529 B.n528 163.367
R803 B.n525 B.n524 163.367
R804 B.n521 B.n520 163.367
R805 B.n517 B.n516 163.367
R806 B.n513 B.n512 163.367
R807 B.n509 B.n508 163.367
R808 B.n505 B.n496 163.367
R809 B.n738 B.n435 163.367
R810 B.n738 B.n433 163.367
R811 B.n742 B.n433 163.367
R812 B.n742 B.n427 163.367
R813 B.n750 B.n427 163.367
R814 B.n750 B.n425 163.367
R815 B.n754 B.n425 163.367
R816 B.n754 B.n420 163.367
R817 B.n763 B.n420 163.367
R818 B.n763 B.n418 163.367
R819 B.n767 B.n418 163.367
R820 B.n767 B.n412 163.367
R821 B.n775 B.n412 163.367
R822 B.n775 B.n410 163.367
R823 B.n779 B.n410 163.367
R824 B.n779 B.n404 163.367
R825 B.n787 B.n404 163.367
R826 B.n787 B.n402 163.367
R827 B.n791 B.n402 163.367
R828 B.n791 B.n396 163.367
R829 B.n799 B.n396 163.367
R830 B.n799 B.n394 163.367
R831 B.n803 B.n394 163.367
R832 B.n803 B.n388 163.367
R833 B.n811 B.n388 163.367
R834 B.n811 B.n386 163.367
R835 B.n815 B.n386 163.367
R836 B.n815 B.n380 163.367
R837 B.n823 B.n380 163.367
R838 B.n823 B.n378 163.367
R839 B.n827 B.n378 163.367
R840 B.n827 B.n373 163.367
R841 B.n836 B.n373 163.367
R842 B.n836 B.n371 163.367
R843 B.n841 B.n371 163.367
R844 B.n841 B.n365 163.367
R845 B.n849 B.n365 163.367
R846 B.n850 B.n849 163.367
R847 B.n850 B.n5 163.367
R848 B.n6 B.n5 163.367
R849 B.n7 B.n6 163.367
R850 B.n855 B.n7 163.367
R851 B.n855 B.n12 163.367
R852 B.n13 B.n12 163.367
R853 B.n14 B.n13 163.367
R854 B.n860 B.n14 163.367
R855 B.n860 B.n19 163.367
R856 B.n20 B.n19 163.367
R857 B.n21 B.n20 163.367
R858 B.n865 B.n21 163.367
R859 B.n865 B.n26 163.367
R860 B.n27 B.n26 163.367
R861 B.n28 B.n27 163.367
R862 B.n870 B.n28 163.367
R863 B.n870 B.n33 163.367
R864 B.n34 B.n33 163.367
R865 B.n35 B.n34 163.367
R866 B.n875 B.n35 163.367
R867 B.n875 B.n40 163.367
R868 B.n41 B.n40 163.367
R869 B.n42 B.n41 163.367
R870 B.n880 B.n42 163.367
R871 B.n880 B.n47 163.367
R872 B.n48 B.n47 163.367
R873 B.n49 B.n48 163.367
R874 B.n885 B.n49 163.367
R875 B.n885 B.n54 163.367
R876 B.n55 B.n54 163.367
R877 B.n56 B.n55 163.367
R878 B.n890 B.n56 163.367
R879 B.n890 B.n61 163.367
R880 B.n62 B.n61 163.367
R881 B.n63 B.n62 163.367
R882 B.n895 B.n63 163.367
R883 B.n895 B.n68 163.367
R884 B.n69 B.n68 163.367
R885 B.n70 B.n69 163.367
R886 B.n132 B.n70 163.367
R887 B.n137 B.n74 163.367
R888 B.n141 B.n140 163.367
R889 B.n145 B.n144 163.367
R890 B.n149 B.n148 163.367
R891 B.n153 B.n152 163.367
R892 B.n157 B.n156 163.367
R893 B.n161 B.n160 163.367
R894 B.n165 B.n164 163.367
R895 B.n169 B.n168 163.367
R896 B.n173 B.n172 163.367
R897 B.n177 B.n176 163.367
R898 B.n181 B.n180 163.367
R899 B.n185 B.n184 163.367
R900 B.n189 B.n188 163.367
R901 B.n193 B.n192 163.367
R902 B.n197 B.n196 163.367
R903 B.n201 B.n200 163.367
R904 B.n205 B.n204 163.367
R905 B.n209 B.n208 163.367
R906 B.n213 B.n212 163.367
R907 B.n217 B.n216 163.367
R908 B.n221 B.n220 163.367
R909 B.n225 B.n224 163.367
R910 B.n229 B.n228 163.367
R911 B.n233 B.n232 163.367
R912 B.n237 B.n236 163.367
R913 B.n242 B.n241 163.367
R914 B.n246 B.n245 163.367
R915 B.n250 B.n249 163.367
R916 B.n254 B.n253 163.367
R917 B.n258 B.n257 163.367
R918 B.n263 B.n262 163.367
R919 B.n267 B.n266 163.367
R920 B.n271 B.n270 163.367
R921 B.n275 B.n274 163.367
R922 B.n279 B.n278 163.367
R923 B.n283 B.n282 163.367
R924 B.n287 B.n286 163.367
R925 B.n291 B.n290 163.367
R926 B.n295 B.n294 163.367
R927 B.n299 B.n298 163.367
R928 B.n303 B.n302 163.367
R929 B.n307 B.n306 163.367
R930 B.n311 B.n310 163.367
R931 B.n315 B.n314 163.367
R932 B.n319 B.n318 163.367
R933 B.n323 B.n322 163.367
R934 B.n327 B.n326 163.367
R935 B.n331 B.n330 163.367
R936 B.n335 B.n334 163.367
R937 B.n339 B.n338 163.367
R938 B.n343 B.n342 163.367
R939 B.n347 B.n346 163.367
R940 B.n351 B.n350 163.367
R941 B.n355 B.n354 163.367
R942 B.n359 B.n358 163.367
R943 B.n361 B.n131 163.367
R944 B.n501 B.t11 141.084
R945 B.n133 B.t13 141.084
R946 B.n498 B.t17 141.064
R947 B.n135 B.t6 141.064
R948 B.n502 B.t10 73.2057
R949 B.n134 B.t14 73.2057
R950 B.n499 B.t16 73.185
R951 B.n136 B.t7 73.185
R952 B.n732 B.n731 71.676
R953 B.n497 B.n440 71.676
R954 B.n724 B.n441 71.676
R955 B.n720 B.n442 71.676
R956 B.n716 B.n443 71.676
R957 B.n712 B.n444 71.676
R958 B.n708 B.n445 71.676
R959 B.n704 B.n446 71.676
R960 B.n700 B.n447 71.676
R961 B.n696 B.n448 71.676
R962 B.n692 B.n449 71.676
R963 B.n688 B.n450 71.676
R964 B.n684 B.n451 71.676
R965 B.n680 B.n452 71.676
R966 B.n676 B.n453 71.676
R967 B.n672 B.n454 71.676
R968 B.n668 B.n455 71.676
R969 B.n664 B.n456 71.676
R970 B.n660 B.n457 71.676
R971 B.n656 B.n458 71.676
R972 B.n652 B.n459 71.676
R973 B.n648 B.n460 71.676
R974 B.n644 B.n461 71.676
R975 B.n640 B.n462 71.676
R976 B.n636 B.n463 71.676
R977 B.n632 B.n464 71.676
R978 B.n628 B.n465 71.676
R979 B.n624 B.n466 71.676
R980 B.n620 B.n467 71.676
R981 B.n616 B.n468 71.676
R982 B.n612 B.n469 71.676
R983 B.n608 B.n470 71.676
R984 B.n604 B.n471 71.676
R985 B.n600 B.n472 71.676
R986 B.n596 B.n473 71.676
R987 B.n592 B.n474 71.676
R988 B.n588 B.n475 71.676
R989 B.n584 B.n476 71.676
R990 B.n580 B.n477 71.676
R991 B.n576 B.n478 71.676
R992 B.n572 B.n479 71.676
R993 B.n568 B.n480 71.676
R994 B.n564 B.n481 71.676
R995 B.n560 B.n482 71.676
R996 B.n556 B.n483 71.676
R997 B.n552 B.n484 71.676
R998 B.n548 B.n485 71.676
R999 B.n544 B.n486 71.676
R1000 B.n540 B.n487 71.676
R1001 B.n536 B.n488 71.676
R1002 B.n532 B.n489 71.676
R1003 B.n528 B.n490 71.676
R1004 B.n524 B.n491 71.676
R1005 B.n520 B.n492 71.676
R1006 B.n516 B.n493 71.676
R1007 B.n512 B.n494 71.676
R1008 B.n508 B.n495 71.676
R1009 B.n906 B.n905 71.676
R1010 B.n137 B.n75 71.676
R1011 B.n141 B.n76 71.676
R1012 B.n145 B.n77 71.676
R1013 B.n149 B.n78 71.676
R1014 B.n153 B.n79 71.676
R1015 B.n157 B.n80 71.676
R1016 B.n161 B.n81 71.676
R1017 B.n165 B.n82 71.676
R1018 B.n169 B.n83 71.676
R1019 B.n173 B.n84 71.676
R1020 B.n177 B.n85 71.676
R1021 B.n181 B.n86 71.676
R1022 B.n185 B.n87 71.676
R1023 B.n189 B.n88 71.676
R1024 B.n193 B.n89 71.676
R1025 B.n197 B.n90 71.676
R1026 B.n201 B.n91 71.676
R1027 B.n205 B.n92 71.676
R1028 B.n209 B.n93 71.676
R1029 B.n213 B.n94 71.676
R1030 B.n217 B.n95 71.676
R1031 B.n221 B.n96 71.676
R1032 B.n225 B.n97 71.676
R1033 B.n229 B.n98 71.676
R1034 B.n233 B.n99 71.676
R1035 B.n237 B.n100 71.676
R1036 B.n242 B.n101 71.676
R1037 B.n246 B.n102 71.676
R1038 B.n250 B.n103 71.676
R1039 B.n254 B.n104 71.676
R1040 B.n258 B.n105 71.676
R1041 B.n263 B.n106 71.676
R1042 B.n267 B.n107 71.676
R1043 B.n271 B.n108 71.676
R1044 B.n275 B.n109 71.676
R1045 B.n279 B.n110 71.676
R1046 B.n283 B.n111 71.676
R1047 B.n287 B.n112 71.676
R1048 B.n291 B.n113 71.676
R1049 B.n295 B.n114 71.676
R1050 B.n299 B.n115 71.676
R1051 B.n303 B.n116 71.676
R1052 B.n307 B.n117 71.676
R1053 B.n311 B.n118 71.676
R1054 B.n315 B.n119 71.676
R1055 B.n319 B.n120 71.676
R1056 B.n323 B.n121 71.676
R1057 B.n327 B.n122 71.676
R1058 B.n331 B.n123 71.676
R1059 B.n335 B.n124 71.676
R1060 B.n339 B.n125 71.676
R1061 B.n343 B.n126 71.676
R1062 B.n347 B.n127 71.676
R1063 B.n351 B.n128 71.676
R1064 B.n355 B.n129 71.676
R1065 B.n359 B.n130 71.676
R1066 B.n903 B.n131 71.676
R1067 B.n903 B.n902 71.676
R1068 B.n361 B.n130 71.676
R1069 B.n358 B.n129 71.676
R1070 B.n354 B.n128 71.676
R1071 B.n350 B.n127 71.676
R1072 B.n346 B.n126 71.676
R1073 B.n342 B.n125 71.676
R1074 B.n338 B.n124 71.676
R1075 B.n334 B.n123 71.676
R1076 B.n330 B.n122 71.676
R1077 B.n326 B.n121 71.676
R1078 B.n322 B.n120 71.676
R1079 B.n318 B.n119 71.676
R1080 B.n314 B.n118 71.676
R1081 B.n310 B.n117 71.676
R1082 B.n306 B.n116 71.676
R1083 B.n302 B.n115 71.676
R1084 B.n298 B.n114 71.676
R1085 B.n294 B.n113 71.676
R1086 B.n290 B.n112 71.676
R1087 B.n286 B.n111 71.676
R1088 B.n282 B.n110 71.676
R1089 B.n278 B.n109 71.676
R1090 B.n274 B.n108 71.676
R1091 B.n270 B.n107 71.676
R1092 B.n266 B.n106 71.676
R1093 B.n262 B.n105 71.676
R1094 B.n257 B.n104 71.676
R1095 B.n253 B.n103 71.676
R1096 B.n249 B.n102 71.676
R1097 B.n245 B.n101 71.676
R1098 B.n241 B.n100 71.676
R1099 B.n236 B.n99 71.676
R1100 B.n232 B.n98 71.676
R1101 B.n228 B.n97 71.676
R1102 B.n224 B.n96 71.676
R1103 B.n220 B.n95 71.676
R1104 B.n216 B.n94 71.676
R1105 B.n212 B.n93 71.676
R1106 B.n208 B.n92 71.676
R1107 B.n204 B.n91 71.676
R1108 B.n200 B.n90 71.676
R1109 B.n196 B.n89 71.676
R1110 B.n192 B.n88 71.676
R1111 B.n188 B.n87 71.676
R1112 B.n184 B.n86 71.676
R1113 B.n180 B.n85 71.676
R1114 B.n176 B.n84 71.676
R1115 B.n172 B.n83 71.676
R1116 B.n168 B.n82 71.676
R1117 B.n164 B.n81 71.676
R1118 B.n160 B.n80 71.676
R1119 B.n156 B.n79 71.676
R1120 B.n152 B.n78 71.676
R1121 B.n148 B.n77 71.676
R1122 B.n144 B.n76 71.676
R1123 B.n140 B.n75 71.676
R1124 B.n905 B.n74 71.676
R1125 B.n731 B.n439 71.676
R1126 B.n725 B.n440 71.676
R1127 B.n721 B.n441 71.676
R1128 B.n717 B.n442 71.676
R1129 B.n713 B.n443 71.676
R1130 B.n709 B.n444 71.676
R1131 B.n705 B.n445 71.676
R1132 B.n701 B.n446 71.676
R1133 B.n697 B.n447 71.676
R1134 B.n693 B.n448 71.676
R1135 B.n689 B.n449 71.676
R1136 B.n685 B.n450 71.676
R1137 B.n681 B.n451 71.676
R1138 B.n677 B.n452 71.676
R1139 B.n673 B.n453 71.676
R1140 B.n669 B.n454 71.676
R1141 B.n665 B.n455 71.676
R1142 B.n661 B.n456 71.676
R1143 B.n657 B.n457 71.676
R1144 B.n653 B.n458 71.676
R1145 B.n649 B.n459 71.676
R1146 B.n645 B.n460 71.676
R1147 B.n641 B.n461 71.676
R1148 B.n637 B.n462 71.676
R1149 B.n633 B.n463 71.676
R1150 B.n629 B.n464 71.676
R1151 B.n625 B.n465 71.676
R1152 B.n621 B.n466 71.676
R1153 B.n617 B.n467 71.676
R1154 B.n613 B.n468 71.676
R1155 B.n609 B.n469 71.676
R1156 B.n605 B.n470 71.676
R1157 B.n601 B.n471 71.676
R1158 B.n597 B.n472 71.676
R1159 B.n593 B.n473 71.676
R1160 B.n589 B.n474 71.676
R1161 B.n585 B.n475 71.676
R1162 B.n581 B.n476 71.676
R1163 B.n577 B.n477 71.676
R1164 B.n573 B.n478 71.676
R1165 B.n569 B.n479 71.676
R1166 B.n565 B.n480 71.676
R1167 B.n561 B.n481 71.676
R1168 B.n557 B.n482 71.676
R1169 B.n553 B.n483 71.676
R1170 B.n549 B.n484 71.676
R1171 B.n545 B.n485 71.676
R1172 B.n541 B.n486 71.676
R1173 B.n537 B.n487 71.676
R1174 B.n533 B.n488 71.676
R1175 B.n529 B.n489 71.676
R1176 B.n525 B.n490 71.676
R1177 B.n521 B.n491 71.676
R1178 B.n517 B.n492 71.676
R1179 B.n513 B.n493 71.676
R1180 B.n509 B.n494 71.676
R1181 B.n505 B.n495 71.676
R1182 B.n502 B.n501 67.8793
R1183 B.n499 B.n498 67.8793
R1184 B.n136 B.n135 67.8793
R1185 B.n134 B.n133 67.8793
R1186 B.n730 B.n436 63.7761
R1187 B.n904 B.n71 63.7761
R1188 B.n503 B.n502 59.5399
R1189 B.n500 B.n499 59.5399
R1190 B.n239 B.n136 59.5399
R1191 B.n260 B.n134 59.5399
R1192 B.n737 B.n436 35.2586
R1193 B.n737 B.n432 35.2586
R1194 B.n743 B.n432 35.2586
R1195 B.n743 B.n428 35.2586
R1196 B.n749 B.n428 35.2586
R1197 B.n749 B.n424 35.2586
R1198 B.n756 B.n424 35.2586
R1199 B.n756 B.n755 35.2586
R1200 B.n762 B.n417 35.2586
R1201 B.n768 B.n417 35.2586
R1202 B.n768 B.n413 35.2586
R1203 B.n774 B.n413 35.2586
R1204 B.n774 B.n409 35.2586
R1205 B.n780 B.n409 35.2586
R1206 B.n780 B.n405 35.2586
R1207 B.n786 B.n405 35.2586
R1208 B.n786 B.n401 35.2586
R1209 B.n792 B.n401 35.2586
R1210 B.n792 B.n397 35.2586
R1211 B.n798 B.n397 35.2586
R1212 B.n804 B.n393 35.2586
R1213 B.n804 B.n389 35.2586
R1214 B.n810 B.n389 35.2586
R1215 B.n810 B.n385 35.2586
R1216 B.n816 B.n385 35.2586
R1217 B.n816 B.n381 35.2586
R1218 B.n822 B.n381 35.2586
R1219 B.n822 B.n377 35.2586
R1220 B.n829 B.n377 35.2586
R1221 B.n829 B.n828 35.2586
R1222 B.n835 B.n370 35.2586
R1223 B.n842 B.n370 35.2586
R1224 B.n842 B.n366 35.2586
R1225 B.n848 B.n366 35.2586
R1226 B.n848 B.n4 35.2586
R1227 B.n985 B.n4 35.2586
R1228 B.n985 B.n984 35.2586
R1229 B.n984 B.n983 35.2586
R1230 B.n983 B.n8 35.2586
R1231 B.n977 B.n8 35.2586
R1232 B.n977 B.n976 35.2586
R1233 B.n976 B.n975 35.2586
R1234 B.n969 B.n18 35.2586
R1235 B.n969 B.n968 35.2586
R1236 B.n968 B.n967 35.2586
R1237 B.n967 B.n22 35.2586
R1238 B.n961 B.n22 35.2586
R1239 B.n961 B.n960 35.2586
R1240 B.n960 B.n959 35.2586
R1241 B.n959 B.n29 35.2586
R1242 B.n953 B.n29 35.2586
R1243 B.n953 B.n952 35.2586
R1244 B.n951 B.n36 35.2586
R1245 B.n945 B.n36 35.2586
R1246 B.n945 B.n944 35.2586
R1247 B.n944 B.n943 35.2586
R1248 B.n943 B.n43 35.2586
R1249 B.n937 B.n43 35.2586
R1250 B.n937 B.n936 35.2586
R1251 B.n936 B.n935 35.2586
R1252 B.n935 B.n50 35.2586
R1253 B.n929 B.n50 35.2586
R1254 B.n929 B.n928 35.2586
R1255 B.n928 B.n927 35.2586
R1256 B.n921 B.n60 35.2586
R1257 B.n921 B.n920 35.2586
R1258 B.n920 B.n919 35.2586
R1259 B.n919 B.n64 35.2586
R1260 B.n913 B.n64 35.2586
R1261 B.n913 B.n912 35.2586
R1262 B.n912 B.n911 35.2586
R1263 B.n911 B.n71 35.2586
R1264 B.n798 B.t1 33.7031
R1265 B.t0 B.n951 33.7031
R1266 B.n908 B.n907 32.3127
R1267 B.n901 B.n900 32.3127
R1268 B.n504 B.n434 32.3127
R1269 B.n734 B.n733 32.3127
R1270 B.n835 B.t2 26.4441
R1271 B.n975 B.t3 26.4441
R1272 B.n762 B.t9 19.185
R1273 B.n927 B.t5 19.185
R1274 B B.n987 18.0485
R1275 B.n755 B.t9 16.074
R1276 B.n60 B.t5 16.074
R1277 B.n907 B.n73 10.6151
R1278 B.n138 B.n73 10.6151
R1279 B.n139 B.n138 10.6151
R1280 B.n142 B.n139 10.6151
R1281 B.n143 B.n142 10.6151
R1282 B.n146 B.n143 10.6151
R1283 B.n147 B.n146 10.6151
R1284 B.n150 B.n147 10.6151
R1285 B.n151 B.n150 10.6151
R1286 B.n154 B.n151 10.6151
R1287 B.n155 B.n154 10.6151
R1288 B.n158 B.n155 10.6151
R1289 B.n159 B.n158 10.6151
R1290 B.n162 B.n159 10.6151
R1291 B.n163 B.n162 10.6151
R1292 B.n166 B.n163 10.6151
R1293 B.n167 B.n166 10.6151
R1294 B.n170 B.n167 10.6151
R1295 B.n171 B.n170 10.6151
R1296 B.n174 B.n171 10.6151
R1297 B.n175 B.n174 10.6151
R1298 B.n178 B.n175 10.6151
R1299 B.n179 B.n178 10.6151
R1300 B.n182 B.n179 10.6151
R1301 B.n183 B.n182 10.6151
R1302 B.n186 B.n183 10.6151
R1303 B.n187 B.n186 10.6151
R1304 B.n190 B.n187 10.6151
R1305 B.n191 B.n190 10.6151
R1306 B.n194 B.n191 10.6151
R1307 B.n195 B.n194 10.6151
R1308 B.n198 B.n195 10.6151
R1309 B.n199 B.n198 10.6151
R1310 B.n202 B.n199 10.6151
R1311 B.n203 B.n202 10.6151
R1312 B.n206 B.n203 10.6151
R1313 B.n207 B.n206 10.6151
R1314 B.n210 B.n207 10.6151
R1315 B.n211 B.n210 10.6151
R1316 B.n214 B.n211 10.6151
R1317 B.n215 B.n214 10.6151
R1318 B.n218 B.n215 10.6151
R1319 B.n219 B.n218 10.6151
R1320 B.n222 B.n219 10.6151
R1321 B.n223 B.n222 10.6151
R1322 B.n226 B.n223 10.6151
R1323 B.n227 B.n226 10.6151
R1324 B.n230 B.n227 10.6151
R1325 B.n231 B.n230 10.6151
R1326 B.n234 B.n231 10.6151
R1327 B.n235 B.n234 10.6151
R1328 B.n238 B.n235 10.6151
R1329 B.n243 B.n240 10.6151
R1330 B.n244 B.n243 10.6151
R1331 B.n247 B.n244 10.6151
R1332 B.n248 B.n247 10.6151
R1333 B.n251 B.n248 10.6151
R1334 B.n252 B.n251 10.6151
R1335 B.n255 B.n252 10.6151
R1336 B.n256 B.n255 10.6151
R1337 B.n259 B.n256 10.6151
R1338 B.n264 B.n261 10.6151
R1339 B.n265 B.n264 10.6151
R1340 B.n268 B.n265 10.6151
R1341 B.n269 B.n268 10.6151
R1342 B.n272 B.n269 10.6151
R1343 B.n273 B.n272 10.6151
R1344 B.n276 B.n273 10.6151
R1345 B.n277 B.n276 10.6151
R1346 B.n280 B.n277 10.6151
R1347 B.n281 B.n280 10.6151
R1348 B.n284 B.n281 10.6151
R1349 B.n285 B.n284 10.6151
R1350 B.n288 B.n285 10.6151
R1351 B.n289 B.n288 10.6151
R1352 B.n292 B.n289 10.6151
R1353 B.n293 B.n292 10.6151
R1354 B.n296 B.n293 10.6151
R1355 B.n297 B.n296 10.6151
R1356 B.n300 B.n297 10.6151
R1357 B.n301 B.n300 10.6151
R1358 B.n304 B.n301 10.6151
R1359 B.n305 B.n304 10.6151
R1360 B.n308 B.n305 10.6151
R1361 B.n309 B.n308 10.6151
R1362 B.n312 B.n309 10.6151
R1363 B.n313 B.n312 10.6151
R1364 B.n316 B.n313 10.6151
R1365 B.n317 B.n316 10.6151
R1366 B.n320 B.n317 10.6151
R1367 B.n321 B.n320 10.6151
R1368 B.n324 B.n321 10.6151
R1369 B.n325 B.n324 10.6151
R1370 B.n328 B.n325 10.6151
R1371 B.n329 B.n328 10.6151
R1372 B.n332 B.n329 10.6151
R1373 B.n333 B.n332 10.6151
R1374 B.n336 B.n333 10.6151
R1375 B.n337 B.n336 10.6151
R1376 B.n340 B.n337 10.6151
R1377 B.n341 B.n340 10.6151
R1378 B.n344 B.n341 10.6151
R1379 B.n345 B.n344 10.6151
R1380 B.n348 B.n345 10.6151
R1381 B.n349 B.n348 10.6151
R1382 B.n352 B.n349 10.6151
R1383 B.n353 B.n352 10.6151
R1384 B.n356 B.n353 10.6151
R1385 B.n357 B.n356 10.6151
R1386 B.n360 B.n357 10.6151
R1387 B.n362 B.n360 10.6151
R1388 B.n363 B.n362 10.6151
R1389 B.n901 B.n363 10.6151
R1390 B.n739 B.n434 10.6151
R1391 B.n740 B.n739 10.6151
R1392 B.n741 B.n740 10.6151
R1393 B.n741 B.n426 10.6151
R1394 B.n751 B.n426 10.6151
R1395 B.n752 B.n751 10.6151
R1396 B.n753 B.n752 10.6151
R1397 B.n753 B.n419 10.6151
R1398 B.n764 B.n419 10.6151
R1399 B.n765 B.n764 10.6151
R1400 B.n766 B.n765 10.6151
R1401 B.n766 B.n411 10.6151
R1402 B.n776 B.n411 10.6151
R1403 B.n777 B.n776 10.6151
R1404 B.n778 B.n777 10.6151
R1405 B.n778 B.n403 10.6151
R1406 B.n788 B.n403 10.6151
R1407 B.n789 B.n788 10.6151
R1408 B.n790 B.n789 10.6151
R1409 B.n790 B.n395 10.6151
R1410 B.n800 B.n395 10.6151
R1411 B.n801 B.n800 10.6151
R1412 B.n802 B.n801 10.6151
R1413 B.n802 B.n387 10.6151
R1414 B.n812 B.n387 10.6151
R1415 B.n813 B.n812 10.6151
R1416 B.n814 B.n813 10.6151
R1417 B.n814 B.n379 10.6151
R1418 B.n824 B.n379 10.6151
R1419 B.n825 B.n824 10.6151
R1420 B.n826 B.n825 10.6151
R1421 B.n826 B.n372 10.6151
R1422 B.n837 B.n372 10.6151
R1423 B.n838 B.n837 10.6151
R1424 B.n840 B.n838 10.6151
R1425 B.n840 B.n839 10.6151
R1426 B.n839 B.n364 10.6151
R1427 B.n851 B.n364 10.6151
R1428 B.n852 B.n851 10.6151
R1429 B.n853 B.n852 10.6151
R1430 B.n854 B.n853 10.6151
R1431 B.n856 B.n854 10.6151
R1432 B.n857 B.n856 10.6151
R1433 B.n858 B.n857 10.6151
R1434 B.n859 B.n858 10.6151
R1435 B.n861 B.n859 10.6151
R1436 B.n862 B.n861 10.6151
R1437 B.n863 B.n862 10.6151
R1438 B.n864 B.n863 10.6151
R1439 B.n866 B.n864 10.6151
R1440 B.n867 B.n866 10.6151
R1441 B.n868 B.n867 10.6151
R1442 B.n869 B.n868 10.6151
R1443 B.n871 B.n869 10.6151
R1444 B.n872 B.n871 10.6151
R1445 B.n873 B.n872 10.6151
R1446 B.n874 B.n873 10.6151
R1447 B.n876 B.n874 10.6151
R1448 B.n877 B.n876 10.6151
R1449 B.n878 B.n877 10.6151
R1450 B.n879 B.n878 10.6151
R1451 B.n881 B.n879 10.6151
R1452 B.n882 B.n881 10.6151
R1453 B.n883 B.n882 10.6151
R1454 B.n884 B.n883 10.6151
R1455 B.n886 B.n884 10.6151
R1456 B.n887 B.n886 10.6151
R1457 B.n888 B.n887 10.6151
R1458 B.n889 B.n888 10.6151
R1459 B.n891 B.n889 10.6151
R1460 B.n892 B.n891 10.6151
R1461 B.n893 B.n892 10.6151
R1462 B.n894 B.n893 10.6151
R1463 B.n896 B.n894 10.6151
R1464 B.n897 B.n896 10.6151
R1465 B.n898 B.n897 10.6151
R1466 B.n899 B.n898 10.6151
R1467 B.n900 B.n899 10.6151
R1468 B.n733 B.n438 10.6151
R1469 B.n728 B.n438 10.6151
R1470 B.n728 B.n727 10.6151
R1471 B.n727 B.n726 10.6151
R1472 B.n726 B.n723 10.6151
R1473 B.n723 B.n722 10.6151
R1474 B.n722 B.n719 10.6151
R1475 B.n719 B.n718 10.6151
R1476 B.n718 B.n715 10.6151
R1477 B.n715 B.n714 10.6151
R1478 B.n714 B.n711 10.6151
R1479 B.n711 B.n710 10.6151
R1480 B.n710 B.n707 10.6151
R1481 B.n707 B.n706 10.6151
R1482 B.n706 B.n703 10.6151
R1483 B.n703 B.n702 10.6151
R1484 B.n702 B.n699 10.6151
R1485 B.n699 B.n698 10.6151
R1486 B.n698 B.n695 10.6151
R1487 B.n695 B.n694 10.6151
R1488 B.n694 B.n691 10.6151
R1489 B.n691 B.n690 10.6151
R1490 B.n690 B.n687 10.6151
R1491 B.n687 B.n686 10.6151
R1492 B.n686 B.n683 10.6151
R1493 B.n683 B.n682 10.6151
R1494 B.n682 B.n679 10.6151
R1495 B.n679 B.n678 10.6151
R1496 B.n678 B.n675 10.6151
R1497 B.n675 B.n674 10.6151
R1498 B.n674 B.n671 10.6151
R1499 B.n671 B.n670 10.6151
R1500 B.n670 B.n667 10.6151
R1501 B.n667 B.n666 10.6151
R1502 B.n666 B.n663 10.6151
R1503 B.n663 B.n662 10.6151
R1504 B.n662 B.n659 10.6151
R1505 B.n659 B.n658 10.6151
R1506 B.n658 B.n655 10.6151
R1507 B.n655 B.n654 10.6151
R1508 B.n654 B.n651 10.6151
R1509 B.n651 B.n650 10.6151
R1510 B.n650 B.n647 10.6151
R1511 B.n647 B.n646 10.6151
R1512 B.n646 B.n643 10.6151
R1513 B.n643 B.n642 10.6151
R1514 B.n642 B.n639 10.6151
R1515 B.n639 B.n638 10.6151
R1516 B.n638 B.n635 10.6151
R1517 B.n635 B.n634 10.6151
R1518 B.n634 B.n631 10.6151
R1519 B.n631 B.n630 10.6151
R1520 B.n627 B.n626 10.6151
R1521 B.n626 B.n623 10.6151
R1522 B.n623 B.n622 10.6151
R1523 B.n622 B.n619 10.6151
R1524 B.n619 B.n618 10.6151
R1525 B.n618 B.n615 10.6151
R1526 B.n615 B.n614 10.6151
R1527 B.n614 B.n611 10.6151
R1528 B.n611 B.n610 10.6151
R1529 B.n607 B.n606 10.6151
R1530 B.n606 B.n603 10.6151
R1531 B.n603 B.n602 10.6151
R1532 B.n602 B.n599 10.6151
R1533 B.n599 B.n598 10.6151
R1534 B.n598 B.n595 10.6151
R1535 B.n595 B.n594 10.6151
R1536 B.n594 B.n591 10.6151
R1537 B.n591 B.n590 10.6151
R1538 B.n590 B.n587 10.6151
R1539 B.n587 B.n586 10.6151
R1540 B.n586 B.n583 10.6151
R1541 B.n583 B.n582 10.6151
R1542 B.n582 B.n579 10.6151
R1543 B.n579 B.n578 10.6151
R1544 B.n578 B.n575 10.6151
R1545 B.n575 B.n574 10.6151
R1546 B.n574 B.n571 10.6151
R1547 B.n571 B.n570 10.6151
R1548 B.n570 B.n567 10.6151
R1549 B.n567 B.n566 10.6151
R1550 B.n566 B.n563 10.6151
R1551 B.n563 B.n562 10.6151
R1552 B.n562 B.n559 10.6151
R1553 B.n559 B.n558 10.6151
R1554 B.n558 B.n555 10.6151
R1555 B.n555 B.n554 10.6151
R1556 B.n554 B.n551 10.6151
R1557 B.n551 B.n550 10.6151
R1558 B.n550 B.n547 10.6151
R1559 B.n547 B.n546 10.6151
R1560 B.n546 B.n543 10.6151
R1561 B.n543 B.n542 10.6151
R1562 B.n542 B.n539 10.6151
R1563 B.n539 B.n538 10.6151
R1564 B.n538 B.n535 10.6151
R1565 B.n535 B.n534 10.6151
R1566 B.n534 B.n531 10.6151
R1567 B.n531 B.n530 10.6151
R1568 B.n530 B.n527 10.6151
R1569 B.n527 B.n526 10.6151
R1570 B.n526 B.n523 10.6151
R1571 B.n523 B.n522 10.6151
R1572 B.n522 B.n519 10.6151
R1573 B.n519 B.n518 10.6151
R1574 B.n518 B.n515 10.6151
R1575 B.n515 B.n514 10.6151
R1576 B.n514 B.n511 10.6151
R1577 B.n511 B.n510 10.6151
R1578 B.n510 B.n507 10.6151
R1579 B.n507 B.n506 10.6151
R1580 B.n506 B.n504 10.6151
R1581 B.n735 B.n734 10.6151
R1582 B.n735 B.n430 10.6151
R1583 B.n745 B.n430 10.6151
R1584 B.n746 B.n745 10.6151
R1585 B.n747 B.n746 10.6151
R1586 B.n747 B.n422 10.6151
R1587 B.n758 B.n422 10.6151
R1588 B.n759 B.n758 10.6151
R1589 B.n760 B.n759 10.6151
R1590 B.n760 B.n415 10.6151
R1591 B.n770 B.n415 10.6151
R1592 B.n771 B.n770 10.6151
R1593 B.n772 B.n771 10.6151
R1594 B.n772 B.n407 10.6151
R1595 B.n782 B.n407 10.6151
R1596 B.n783 B.n782 10.6151
R1597 B.n784 B.n783 10.6151
R1598 B.n784 B.n399 10.6151
R1599 B.n794 B.n399 10.6151
R1600 B.n795 B.n794 10.6151
R1601 B.n796 B.n795 10.6151
R1602 B.n796 B.n391 10.6151
R1603 B.n806 B.n391 10.6151
R1604 B.n807 B.n806 10.6151
R1605 B.n808 B.n807 10.6151
R1606 B.n808 B.n383 10.6151
R1607 B.n818 B.n383 10.6151
R1608 B.n819 B.n818 10.6151
R1609 B.n820 B.n819 10.6151
R1610 B.n820 B.n375 10.6151
R1611 B.n831 B.n375 10.6151
R1612 B.n832 B.n831 10.6151
R1613 B.n833 B.n832 10.6151
R1614 B.n833 B.n368 10.6151
R1615 B.n844 B.n368 10.6151
R1616 B.n845 B.n844 10.6151
R1617 B.n846 B.n845 10.6151
R1618 B.n846 B.n0 10.6151
R1619 B.n981 B.n1 10.6151
R1620 B.n981 B.n980 10.6151
R1621 B.n980 B.n979 10.6151
R1622 B.n979 B.n10 10.6151
R1623 B.n973 B.n10 10.6151
R1624 B.n973 B.n972 10.6151
R1625 B.n972 B.n971 10.6151
R1626 B.n971 B.n16 10.6151
R1627 B.n965 B.n16 10.6151
R1628 B.n965 B.n964 10.6151
R1629 B.n964 B.n963 10.6151
R1630 B.n963 B.n24 10.6151
R1631 B.n957 B.n24 10.6151
R1632 B.n957 B.n956 10.6151
R1633 B.n956 B.n955 10.6151
R1634 B.n955 B.n31 10.6151
R1635 B.n949 B.n31 10.6151
R1636 B.n949 B.n948 10.6151
R1637 B.n948 B.n947 10.6151
R1638 B.n947 B.n38 10.6151
R1639 B.n941 B.n38 10.6151
R1640 B.n941 B.n940 10.6151
R1641 B.n940 B.n939 10.6151
R1642 B.n939 B.n45 10.6151
R1643 B.n933 B.n45 10.6151
R1644 B.n933 B.n932 10.6151
R1645 B.n932 B.n931 10.6151
R1646 B.n931 B.n52 10.6151
R1647 B.n925 B.n52 10.6151
R1648 B.n925 B.n924 10.6151
R1649 B.n924 B.n923 10.6151
R1650 B.n923 B.n58 10.6151
R1651 B.n917 B.n58 10.6151
R1652 B.n917 B.n916 10.6151
R1653 B.n916 B.n915 10.6151
R1654 B.n915 B.n66 10.6151
R1655 B.n909 B.n66 10.6151
R1656 B.n909 B.n908 10.6151
R1657 B.n239 B.n238 9.36635
R1658 B.n261 B.n260 9.36635
R1659 B.n630 B.n500 9.36635
R1660 B.n607 B.n503 9.36635
R1661 B.n828 B.t2 8.81502
R1662 B.n18 B.t3 8.81502
R1663 B.n987 B.n0 2.81026
R1664 B.n987 B.n1 2.81026
R1665 B.t1 B.n393 1.556
R1666 B.n952 B.t0 1.556
R1667 B.n240 B.n239 1.24928
R1668 B.n260 B.n259 1.24928
R1669 B.n627 B.n500 1.24928
R1670 B.n610 B.n503 1.24928
R1671 VP.n17 VP.n16 161.3
R1672 VP.n15 VP.n1 161.3
R1673 VP.n14 VP.n13 161.3
R1674 VP.n12 VP.n2 161.3
R1675 VP.n11 VP.n10 161.3
R1676 VP.n9 VP.n3 161.3
R1677 VP.n8 VP.n7 161.3
R1678 VP.n5 VP.t3 155.653
R1679 VP.n5 VP.t2 154.565
R1680 VP.n4 VP.t1 121.184
R1681 VP.n0 VP.t0 121.184
R1682 VP.n6 VP.n4 77.7193
R1683 VP.n18 VP.n0 77.7193
R1684 VP.n6 VP.n5 53.6923
R1685 VP.n10 VP.n2 40.4106
R1686 VP.n14 VP.n2 40.4106
R1687 VP.n9 VP.n8 24.3439
R1688 VP.n10 VP.n9 24.3439
R1689 VP.n15 VP.n14 24.3439
R1690 VP.n16 VP.n15 24.3439
R1691 VP.n8 VP.n4 12.1722
R1692 VP.n16 VP.n0 12.1722
R1693 VP.n7 VP.n6 0.355081
R1694 VP.n18 VP.n17 0.355081
R1695 VP VP.n18 0.26685
R1696 VP.n7 VP.n3 0.189894
R1697 VP.n11 VP.n3 0.189894
R1698 VP.n12 VP.n11 0.189894
R1699 VP.n13 VP.n12 0.189894
R1700 VP.n13 VP.n1 0.189894
R1701 VP.n17 VP.n1 0.189894
R1702 VTAIL.n5 VTAIL.t6 49.6383
R1703 VTAIL.n4 VTAIL.t2 49.6383
R1704 VTAIL.n3 VTAIL.t1 49.6383
R1705 VTAIL.n7 VTAIL.t0 49.6382
R1706 VTAIL.n0 VTAIL.t3 49.6382
R1707 VTAIL.n1 VTAIL.t5 49.6382
R1708 VTAIL.n2 VTAIL.t4 49.6382
R1709 VTAIL.n6 VTAIL.t7 49.6382
R1710 VTAIL.n7 VTAIL.n6 29.1255
R1711 VTAIL.n3 VTAIL.n2 29.1255
R1712 VTAIL.n4 VTAIL.n3 3.01774
R1713 VTAIL.n6 VTAIL.n5 3.01774
R1714 VTAIL.n2 VTAIL.n1 3.01774
R1715 VTAIL VTAIL.n0 1.56731
R1716 VTAIL VTAIL.n7 1.45093
R1717 VTAIL.n5 VTAIL.n4 0.470328
R1718 VTAIL.n1 VTAIL.n0 0.470328
R1719 VDD1 VDD1.n1 112.108
R1720 VDD1 VDD1.n0 65.133
R1721 VDD1.n0 VDD1.t0 1.24266
R1722 VDD1.n0 VDD1.t1 1.24266
R1723 VDD1.n1 VDD1.t2 1.24266
R1724 VDD1.n1 VDD1.t3 1.24266
R1725 VN.n0 VN.t3 155.653
R1726 VN.n1 VN.t2 155.653
R1727 VN.n0 VN.t0 154.565
R1728 VN.n1 VN.t1 154.565
R1729 VN VN.n1 53.8578
R1730 VN VN.n0 2.67215
R1731 VDD2.n2 VDD2.n0 111.582
R1732 VDD2.n2 VDD2.n1 65.0748
R1733 VDD2.n1 VDD2.t2 1.24266
R1734 VDD2.n1 VDD2.t1 1.24266
R1735 VDD2.n0 VDD2.t0 1.24266
R1736 VDD2.n0 VDD2.t3 1.24266
R1737 VDD2 VDD2.n2 0.0586897
C0 VP VDD2 0.430085f
C1 VN VDD1 0.149025f
C2 VP VN 7.34043f
C3 VP VDD1 6.69814f
C4 VDD2 VTAIL 6.46518f
C5 VN VTAIL 6.2283f
C6 VDD1 VTAIL 6.40715f
C7 VP VTAIL 6.24241f
C8 VDD2 VN 6.41796f
C9 VDD2 VDD1 1.16508f
C10 VDD2 B 4.391197f
C11 VDD1 B 9.14799f
C12 VTAIL B 12.77719f
C13 VN B 12.11051f
C14 VP B 10.431564f
C15 VDD2.t0 B 0.337114f
C16 VDD2.t3 B 0.337114f
C17 VDD2.n0 B 3.88078f
C18 VDD2.t2 B 0.337114f
C19 VDD2.t1 B 0.337114f
C20 VDD2.n1 B 3.06035f
C21 VDD2.n2 B 4.34446f
C22 VN.t0 B 3.2228f
C23 VN.t3 B 3.23087f
C24 VN.n0 B 2.00874f
C25 VN.t1 B 3.2228f
C26 VN.t2 B 3.23087f
C27 VN.n1 B 3.41541f
C28 VDD1.t0 B 0.339737f
C29 VDD1.t1 B 0.339737f
C30 VDD1.n0 B 3.0846f
C31 VDD1.t2 B 0.339737f
C32 VDD1.t3 B 0.339737f
C33 VDD1.n1 B 3.93862f
C34 VTAIL.t3 B 2.25954f
C35 VTAIL.n0 B 0.305695f
C36 VTAIL.t5 B 2.25954f
C37 VTAIL.n1 B 0.379721f
C38 VTAIL.t4 B 2.25954f
C39 VTAIL.n2 B 1.4262f
C40 VTAIL.t1 B 2.25955f
C41 VTAIL.n3 B 1.42619f
C42 VTAIL.t2 B 2.25955f
C43 VTAIL.n4 B 0.379707f
C44 VTAIL.t6 B 2.25955f
C45 VTAIL.n5 B 0.379707f
C46 VTAIL.t7 B 2.25954f
C47 VTAIL.n6 B 1.4262f
C48 VTAIL.t0 B 2.25954f
C49 VTAIL.n7 B 1.34624f
C50 VP.t0 B 3.01738f
C51 VP.n0 B 1.12732f
C52 VP.n1 B 0.021763f
C53 VP.n2 B 0.017611f
C54 VP.n3 B 0.021763f
C55 VP.t1 B 3.01738f
C56 VP.n4 B 1.12732f
C57 VP.t3 B 3.28454f
C58 VP.t2 B 3.27634f
C59 VP.n5 B 3.4635f
C60 VP.n6 B 1.36628f
C61 VP.n7 B 0.035131f
C62 VP.n8 B 0.030701f
C63 VP.n9 B 0.040764f
C64 VP.n10 B 0.043485f
C65 VP.n11 B 0.021763f
C66 VP.n12 B 0.021763f
C67 VP.n13 B 0.021763f
C68 VP.n14 B 0.043485f
C69 VP.n15 B 0.040764f
C70 VP.n16 B 0.030701f
C71 VP.n17 B 0.035131f
C72 VP.n18 B 0.053496f
.ends

