* NGSPICE file created from diff_pair_sample_1494.ext - technology: sky130A

.subckt diff_pair_sample_1494 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t14 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=3
X1 B.t11 B.t9 B.t10 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=3
X2 VDD1.t9 VP.t0 VTAIL.t6 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=3
X3 VDD2.t8 VN.t1 VTAIL.t10 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X4 VDD1.t8 VP.t1 VTAIL.t2 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=3
X5 VDD2.t7 VN.t2 VTAIL.t15 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X6 VDD2.t6 VN.t3 VTAIL.t18 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=3
X7 VTAIL.t9 VN.t4 VDD2.t5 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X8 VTAIL.t8 VP.t2 VDD1.t7 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X9 VTAIL.t11 VN.t5 VDD2.t4 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X10 VDD1.t6 VP.t3 VTAIL.t5 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=3
X11 VDD1.t5 VP.t4 VTAIL.t7 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X12 VDD1.t4 VP.t5 VTAIL.t4 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=3
X13 B.t8 B.t6 B.t7 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=3
X14 VTAIL.t19 VP.t6 VDD1.t3 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X15 VTAIL.t3 VP.t7 VDD1.t2 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X16 VTAIL.t17 VN.t6 VDD2.t3 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X17 VTAIL.t0 VP.t8 VDD1.t1 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X18 VDD1.t0 VP.t9 VTAIL.t1 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X19 VTAIL.t12 VN.t7 VDD2.t2 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=3
X20 VDD2.t1 VN.t8 VTAIL.t16 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=3
X21 B.t5 B.t3 B.t4 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=3
X22 VDD2.t0 VN.t9 VTAIL.t13 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=3
X23 B.t2 B.t0 B.t1 w_n4966_n2402# sky130_fd_pr__pfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=3
R0 VN.n90 VN.n89 161.3
R1 VN.n88 VN.n47 161.3
R2 VN.n87 VN.n86 161.3
R3 VN.n85 VN.n48 161.3
R4 VN.n84 VN.n83 161.3
R5 VN.n82 VN.n49 161.3
R6 VN.n80 VN.n79 161.3
R7 VN.n78 VN.n50 161.3
R8 VN.n77 VN.n76 161.3
R9 VN.n75 VN.n51 161.3
R10 VN.n74 VN.n73 161.3
R11 VN.n72 VN.n52 161.3
R12 VN.n71 VN.n70 161.3
R13 VN.n68 VN.n53 161.3
R14 VN.n67 VN.n66 161.3
R15 VN.n65 VN.n54 161.3
R16 VN.n64 VN.n63 161.3
R17 VN.n62 VN.n55 161.3
R18 VN.n61 VN.n60 161.3
R19 VN.n59 VN.n56 161.3
R20 VN.n44 VN.n43 161.3
R21 VN.n42 VN.n1 161.3
R22 VN.n41 VN.n40 161.3
R23 VN.n39 VN.n2 161.3
R24 VN.n38 VN.n37 161.3
R25 VN.n36 VN.n3 161.3
R26 VN.n34 VN.n33 161.3
R27 VN.n32 VN.n4 161.3
R28 VN.n31 VN.n30 161.3
R29 VN.n29 VN.n5 161.3
R30 VN.n28 VN.n27 161.3
R31 VN.n26 VN.n6 161.3
R32 VN.n25 VN.n24 161.3
R33 VN.n22 VN.n7 161.3
R34 VN.n21 VN.n20 161.3
R35 VN.n19 VN.n8 161.3
R36 VN.n18 VN.n17 161.3
R37 VN.n16 VN.n9 161.3
R38 VN.n15 VN.n14 161.3
R39 VN.n13 VN.n10 161.3
R40 VN.n58 VN.t3 89.3011
R41 VN.n12 VN.t9 89.3011
R42 VN.n45 VN.n0 70.0045
R43 VN.n91 VN.n46 70.0045
R44 VN.n12 VN.n11 69.746
R45 VN.n58 VN.n57 69.746
R46 VN.n11 VN.t5 57.5995
R47 VN.n23 VN.t2 57.5995
R48 VN.n35 VN.t6 57.5995
R49 VN.n0 VN.t0 57.5995
R50 VN.n57 VN.t4 57.5995
R51 VN.n69 VN.t1 57.5995
R52 VN.n81 VN.t7 57.5995
R53 VN.n46 VN.t8 57.5995
R54 VN.n41 VN.n2 56.5193
R55 VN.n87 VN.n48 56.5193
R56 VN VN.n91 51.9185
R57 VN.n17 VN.n8 48.7492
R58 VN.n29 VN.n28 48.7492
R59 VN.n63 VN.n54 48.7492
R60 VN.n75 VN.n74 48.7492
R61 VN.n17 VN.n16 32.2376
R62 VN.n30 VN.n29 32.2376
R63 VN.n63 VN.n62 32.2376
R64 VN.n76 VN.n75 32.2376
R65 VN.n15 VN.n10 24.4675
R66 VN.n16 VN.n15 24.4675
R67 VN.n21 VN.n8 24.4675
R68 VN.n22 VN.n21 24.4675
R69 VN.n24 VN.n6 24.4675
R70 VN.n28 VN.n6 24.4675
R71 VN.n30 VN.n4 24.4675
R72 VN.n34 VN.n4 24.4675
R73 VN.n37 VN.n36 24.4675
R74 VN.n37 VN.n2 24.4675
R75 VN.n42 VN.n41 24.4675
R76 VN.n43 VN.n42 24.4675
R77 VN.n62 VN.n61 24.4675
R78 VN.n61 VN.n56 24.4675
R79 VN.n74 VN.n52 24.4675
R80 VN.n70 VN.n52 24.4675
R81 VN.n68 VN.n67 24.4675
R82 VN.n67 VN.n54 24.4675
R83 VN.n83 VN.n48 24.4675
R84 VN.n83 VN.n82 24.4675
R85 VN.n80 VN.n50 24.4675
R86 VN.n76 VN.n50 24.4675
R87 VN.n89 VN.n88 24.4675
R88 VN.n88 VN.n87 24.4675
R89 VN.n36 VN.n35 20.5528
R90 VN.n82 VN.n81 20.5528
R91 VN.n43 VN.n0 20.0634
R92 VN.n89 VN.n46 20.0634
R93 VN.n23 VN.n22 12.234
R94 VN.n24 VN.n23 12.234
R95 VN.n70 VN.n69 12.234
R96 VN.n69 VN.n68 12.234
R97 VN.n59 VN.n58 5.54917
R98 VN.n13 VN.n12 5.54917
R99 VN.n11 VN.n10 3.91522
R100 VN.n35 VN.n34 3.91522
R101 VN.n57 VN.n56 3.91522
R102 VN.n81 VN.n80 3.91522
R103 VN.n91 VN.n90 0.354971
R104 VN.n45 VN.n44 0.354971
R105 VN VN.n45 0.26696
R106 VN.n90 VN.n47 0.189894
R107 VN.n86 VN.n47 0.189894
R108 VN.n86 VN.n85 0.189894
R109 VN.n85 VN.n84 0.189894
R110 VN.n84 VN.n49 0.189894
R111 VN.n79 VN.n49 0.189894
R112 VN.n79 VN.n78 0.189894
R113 VN.n78 VN.n77 0.189894
R114 VN.n77 VN.n51 0.189894
R115 VN.n73 VN.n51 0.189894
R116 VN.n73 VN.n72 0.189894
R117 VN.n72 VN.n71 0.189894
R118 VN.n71 VN.n53 0.189894
R119 VN.n66 VN.n53 0.189894
R120 VN.n66 VN.n65 0.189894
R121 VN.n65 VN.n64 0.189894
R122 VN.n64 VN.n55 0.189894
R123 VN.n60 VN.n55 0.189894
R124 VN.n60 VN.n59 0.189894
R125 VN.n14 VN.n13 0.189894
R126 VN.n14 VN.n9 0.189894
R127 VN.n18 VN.n9 0.189894
R128 VN.n19 VN.n18 0.189894
R129 VN.n20 VN.n19 0.189894
R130 VN.n20 VN.n7 0.189894
R131 VN.n25 VN.n7 0.189894
R132 VN.n26 VN.n25 0.189894
R133 VN.n27 VN.n26 0.189894
R134 VN.n27 VN.n5 0.189894
R135 VN.n31 VN.n5 0.189894
R136 VN.n32 VN.n31 0.189894
R137 VN.n33 VN.n32 0.189894
R138 VN.n33 VN.n3 0.189894
R139 VN.n38 VN.n3 0.189894
R140 VN.n39 VN.n38 0.189894
R141 VN.n40 VN.n39 0.189894
R142 VN.n40 VN.n1 0.189894
R143 VN.n44 VN.n1 0.189894
R144 VTAIL.n135 VTAIL.n134 585
R145 VTAIL.n137 VTAIL.n136 585
R146 VTAIL.n130 VTAIL.n129 585
R147 VTAIL.n143 VTAIL.n142 585
R148 VTAIL.n145 VTAIL.n144 585
R149 VTAIL.n126 VTAIL.n125 585
R150 VTAIL.n151 VTAIL.n150 585
R151 VTAIL.n153 VTAIL.n152 585
R152 VTAIL.n15 VTAIL.n14 585
R153 VTAIL.n17 VTAIL.n16 585
R154 VTAIL.n10 VTAIL.n9 585
R155 VTAIL.n23 VTAIL.n22 585
R156 VTAIL.n25 VTAIL.n24 585
R157 VTAIL.n6 VTAIL.n5 585
R158 VTAIL.n31 VTAIL.n30 585
R159 VTAIL.n33 VTAIL.n32 585
R160 VTAIL.n117 VTAIL.n116 585
R161 VTAIL.n115 VTAIL.n114 585
R162 VTAIL.n90 VTAIL.n89 585
R163 VTAIL.n109 VTAIL.n108 585
R164 VTAIL.n107 VTAIL.n106 585
R165 VTAIL.n94 VTAIL.n93 585
R166 VTAIL.n101 VTAIL.n100 585
R167 VTAIL.n99 VTAIL.n98 585
R168 VTAIL.n77 VTAIL.n76 585
R169 VTAIL.n75 VTAIL.n74 585
R170 VTAIL.n50 VTAIL.n49 585
R171 VTAIL.n69 VTAIL.n68 585
R172 VTAIL.n67 VTAIL.n66 585
R173 VTAIL.n54 VTAIL.n53 585
R174 VTAIL.n61 VTAIL.n60 585
R175 VTAIL.n59 VTAIL.n58 585
R176 VTAIL.n152 VTAIL.n122 498.474
R177 VTAIL.n32 VTAIL.n2 498.474
R178 VTAIL.n116 VTAIL.n86 498.474
R179 VTAIL.n76 VTAIL.n46 498.474
R180 VTAIL.n133 VTAIL.t14 329.053
R181 VTAIL.n13 VTAIL.t6 329.053
R182 VTAIL.n97 VTAIL.t4 329.053
R183 VTAIL.n57 VTAIL.t18 329.053
R184 VTAIL.n136 VTAIL.n135 171.744
R185 VTAIL.n136 VTAIL.n129 171.744
R186 VTAIL.n143 VTAIL.n129 171.744
R187 VTAIL.n144 VTAIL.n143 171.744
R188 VTAIL.n144 VTAIL.n125 171.744
R189 VTAIL.n151 VTAIL.n125 171.744
R190 VTAIL.n152 VTAIL.n151 171.744
R191 VTAIL.n16 VTAIL.n15 171.744
R192 VTAIL.n16 VTAIL.n9 171.744
R193 VTAIL.n23 VTAIL.n9 171.744
R194 VTAIL.n24 VTAIL.n23 171.744
R195 VTAIL.n24 VTAIL.n5 171.744
R196 VTAIL.n31 VTAIL.n5 171.744
R197 VTAIL.n32 VTAIL.n31 171.744
R198 VTAIL.n116 VTAIL.n115 171.744
R199 VTAIL.n115 VTAIL.n89 171.744
R200 VTAIL.n108 VTAIL.n89 171.744
R201 VTAIL.n108 VTAIL.n107 171.744
R202 VTAIL.n107 VTAIL.n93 171.744
R203 VTAIL.n100 VTAIL.n93 171.744
R204 VTAIL.n100 VTAIL.n99 171.744
R205 VTAIL.n76 VTAIL.n75 171.744
R206 VTAIL.n75 VTAIL.n49 171.744
R207 VTAIL.n68 VTAIL.n49 171.744
R208 VTAIL.n68 VTAIL.n67 171.744
R209 VTAIL.n67 VTAIL.n53 171.744
R210 VTAIL.n60 VTAIL.n53 171.744
R211 VTAIL.n60 VTAIL.n59 171.744
R212 VTAIL.n135 VTAIL.t14 85.8723
R213 VTAIL.n15 VTAIL.t6 85.8723
R214 VTAIL.n99 VTAIL.t4 85.8723
R215 VTAIL.n59 VTAIL.t18 85.8723
R216 VTAIL.n85 VTAIL.n84 69.9055
R217 VTAIL.n83 VTAIL.n82 69.9055
R218 VTAIL.n45 VTAIL.n44 69.9055
R219 VTAIL.n43 VTAIL.n42 69.9055
R220 VTAIL.n159 VTAIL.n158 69.9054
R221 VTAIL.n1 VTAIL.n0 69.9054
R222 VTAIL.n39 VTAIL.n38 69.9054
R223 VTAIL.n41 VTAIL.n40 69.9054
R224 VTAIL.n157 VTAIL.n156 33.9308
R225 VTAIL.n37 VTAIL.n36 33.9308
R226 VTAIL.n121 VTAIL.n120 33.9308
R227 VTAIL.n81 VTAIL.n80 33.9308
R228 VTAIL.n43 VTAIL.n41 24.2893
R229 VTAIL.n157 VTAIL.n121 21.4186
R230 VTAIL.n154 VTAIL.n153 12.8005
R231 VTAIL.n34 VTAIL.n33 12.8005
R232 VTAIL.n118 VTAIL.n117 12.8005
R233 VTAIL.n78 VTAIL.n77 12.8005
R234 VTAIL.n150 VTAIL.n124 12.0247
R235 VTAIL.n30 VTAIL.n4 12.0247
R236 VTAIL.n114 VTAIL.n88 12.0247
R237 VTAIL.n74 VTAIL.n48 12.0247
R238 VTAIL.n149 VTAIL.n126 11.249
R239 VTAIL.n29 VTAIL.n6 11.249
R240 VTAIL.n113 VTAIL.n90 11.249
R241 VTAIL.n73 VTAIL.n50 11.249
R242 VTAIL.n134 VTAIL.n133 10.7237
R243 VTAIL.n14 VTAIL.n13 10.7237
R244 VTAIL.n98 VTAIL.n97 10.7237
R245 VTAIL.n58 VTAIL.n57 10.7237
R246 VTAIL.n146 VTAIL.n145 10.4732
R247 VTAIL.n26 VTAIL.n25 10.4732
R248 VTAIL.n110 VTAIL.n109 10.4732
R249 VTAIL.n70 VTAIL.n69 10.4732
R250 VTAIL.n142 VTAIL.n128 9.69747
R251 VTAIL.n22 VTAIL.n8 9.69747
R252 VTAIL.n106 VTAIL.n92 9.69747
R253 VTAIL.n66 VTAIL.n52 9.69747
R254 VTAIL.n156 VTAIL.n155 9.45567
R255 VTAIL.n36 VTAIL.n35 9.45567
R256 VTAIL.n120 VTAIL.n119 9.45567
R257 VTAIL.n80 VTAIL.n79 9.45567
R258 VTAIL.n132 VTAIL.n131 9.3005
R259 VTAIL.n139 VTAIL.n138 9.3005
R260 VTAIL.n141 VTAIL.n140 9.3005
R261 VTAIL.n128 VTAIL.n127 9.3005
R262 VTAIL.n147 VTAIL.n146 9.3005
R263 VTAIL.n149 VTAIL.n148 9.3005
R264 VTAIL.n124 VTAIL.n123 9.3005
R265 VTAIL.n155 VTAIL.n154 9.3005
R266 VTAIL.n12 VTAIL.n11 9.3005
R267 VTAIL.n19 VTAIL.n18 9.3005
R268 VTAIL.n21 VTAIL.n20 9.3005
R269 VTAIL.n8 VTAIL.n7 9.3005
R270 VTAIL.n27 VTAIL.n26 9.3005
R271 VTAIL.n29 VTAIL.n28 9.3005
R272 VTAIL.n4 VTAIL.n3 9.3005
R273 VTAIL.n35 VTAIL.n34 9.3005
R274 VTAIL.n96 VTAIL.n95 9.3005
R275 VTAIL.n103 VTAIL.n102 9.3005
R276 VTAIL.n105 VTAIL.n104 9.3005
R277 VTAIL.n92 VTAIL.n91 9.3005
R278 VTAIL.n111 VTAIL.n110 9.3005
R279 VTAIL.n113 VTAIL.n112 9.3005
R280 VTAIL.n88 VTAIL.n87 9.3005
R281 VTAIL.n119 VTAIL.n118 9.3005
R282 VTAIL.n56 VTAIL.n55 9.3005
R283 VTAIL.n63 VTAIL.n62 9.3005
R284 VTAIL.n65 VTAIL.n64 9.3005
R285 VTAIL.n52 VTAIL.n51 9.3005
R286 VTAIL.n71 VTAIL.n70 9.3005
R287 VTAIL.n73 VTAIL.n72 9.3005
R288 VTAIL.n48 VTAIL.n47 9.3005
R289 VTAIL.n79 VTAIL.n78 9.3005
R290 VTAIL.n141 VTAIL.n130 8.92171
R291 VTAIL.n21 VTAIL.n10 8.92171
R292 VTAIL.n105 VTAIL.n94 8.92171
R293 VTAIL.n65 VTAIL.n54 8.92171
R294 VTAIL.n138 VTAIL.n137 8.14595
R295 VTAIL.n18 VTAIL.n17 8.14595
R296 VTAIL.n102 VTAIL.n101 8.14595
R297 VTAIL.n62 VTAIL.n61 8.14595
R298 VTAIL.n156 VTAIL.n122 7.75445
R299 VTAIL.n36 VTAIL.n2 7.75445
R300 VTAIL.n120 VTAIL.n86 7.75445
R301 VTAIL.n80 VTAIL.n46 7.75445
R302 VTAIL.n134 VTAIL.n132 7.3702
R303 VTAIL.n14 VTAIL.n12 7.3702
R304 VTAIL.n98 VTAIL.n96 7.3702
R305 VTAIL.n58 VTAIL.n56 7.3702
R306 VTAIL.n154 VTAIL.n122 6.08283
R307 VTAIL.n34 VTAIL.n2 6.08283
R308 VTAIL.n118 VTAIL.n86 6.08283
R309 VTAIL.n78 VTAIL.n46 6.08283
R310 VTAIL.n137 VTAIL.n132 5.81868
R311 VTAIL.n17 VTAIL.n12 5.81868
R312 VTAIL.n101 VTAIL.n96 5.81868
R313 VTAIL.n61 VTAIL.n56 5.81868
R314 VTAIL.n138 VTAIL.n130 5.04292
R315 VTAIL.n18 VTAIL.n10 5.04292
R316 VTAIL.n102 VTAIL.n94 5.04292
R317 VTAIL.n62 VTAIL.n54 5.04292
R318 VTAIL.n158 VTAIL.t15 4.53397
R319 VTAIL.n158 VTAIL.t17 4.53397
R320 VTAIL.n0 VTAIL.t13 4.53397
R321 VTAIL.n0 VTAIL.t11 4.53397
R322 VTAIL.n38 VTAIL.t7 4.53397
R323 VTAIL.n38 VTAIL.t3 4.53397
R324 VTAIL.n40 VTAIL.t2 4.53397
R325 VTAIL.n40 VTAIL.t19 4.53397
R326 VTAIL.n84 VTAIL.t1 4.53397
R327 VTAIL.n84 VTAIL.t0 4.53397
R328 VTAIL.n82 VTAIL.t5 4.53397
R329 VTAIL.n82 VTAIL.t8 4.53397
R330 VTAIL.n44 VTAIL.t10 4.53397
R331 VTAIL.n44 VTAIL.t9 4.53397
R332 VTAIL.n42 VTAIL.t16 4.53397
R333 VTAIL.n42 VTAIL.t12 4.53397
R334 VTAIL.n142 VTAIL.n141 4.26717
R335 VTAIL.n22 VTAIL.n21 4.26717
R336 VTAIL.n106 VTAIL.n105 4.26717
R337 VTAIL.n66 VTAIL.n65 4.26717
R338 VTAIL.n145 VTAIL.n128 3.49141
R339 VTAIL.n25 VTAIL.n8 3.49141
R340 VTAIL.n109 VTAIL.n92 3.49141
R341 VTAIL.n69 VTAIL.n52 3.49141
R342 VTAIL.n45 VTAIL.n43 2.87119
R343 VTAIL.n81 VTAIL.n45 2.87119
R344 VTAIL.n85 VTAIL.n83 2.87119
R345 VTAIL.n121 VTAIL.n85 2.87119
R346 VTAIL.n41 VTAIL.n39 2.87119
R347 VTAIL.n39 VTAIL.n37 2.87119
R348 VTAIL.n159 VTAIL.n157 2.87119
R349 VTAIL.n146 VTAIL.n126 2.71565
R350 VTAIL.n26 VTAIL.n6 2.71565
R351 VTAIL.n110 VTAIL.n90 2.71565
R352 VTAIL.n70 VTAIL.n50 2.71565
R353 VTAIL.n133 VTAIL.n131 2.41305
R354 VTAIL.n13 VTAIL.n11 2.41305
R355 VTAIL.n97 VTAIL.n95 2.41305
R356 VTAIL.n57 VTAIL.n55 2.41305
R357 VTAIL VTAIL.n1 2.21171
R358 VTAIL.n150 VTAIL.n149 1.93989
R359 VTAIL.n30 VTAIL.n29 1.93989
R360 VTAIL.n114 VTAIL.n113 1.93989
R361 VTAIL.n74 VTAIL.n73 1.93989
R362 VTAIL.n83 VTAIL.n81 1.90567
R363 VTAIL.n37 VTAIL.n1 1.90567
R364 VTAIL.n153 VTAIL.n124 1.16414
R365 VTAIL.n33 VTAIL.n4 1.16414
R366 VTAIL.n117 VTAIL.n88 1.16414
R367 VTAIL.n77 VTAIL.n48 1.16414
R368 VTAIL VTAIL.n159 0.659983
R369 VTAIL.n139 VTAIL.n131 0.155672
R370 VTAIL.n140 VTAIL.n139 0.155672
R371 VTAIL.n140 VTAIL.n127 0.155672
R372 VTAIL.n147 VTAIL.n127 0.155672
R373 VTAIL.n148 VTAIL.n147 0.155672
R374 VTAIL.n148 VTAIL.n123 0.155672
R375 VTAIL.n155 VTAIL.n123 0.155672
R376 VTAIL.n19 VTAIL.n11 0.155672
R377 VTAIL.n20 VTAIL.n19 0.155672
R378 VTAIL.n20 VTAIL.n7 0.155672
R379 VTAIL.n27 VTAIL.n7 0.155672
R380 VTAIL.n28 VTAIL.n27 0.155672
R381 VTAIL.n28 VTAIL.n3 0.155672
R382 VTAIL.n35 VTAIL.n3 0.155672
R383 VTAIL.n119 VTAIL.n87 0.155672
R384 VTAIL.n112 VTAIL.n87 0.155672
R385 VTAIL.n112 VTAIL.n111 0.155672
R386 VTAIL.n111 VTAIL.n91 0.155672
R387 VTAIL.n104 VTAIL.n91 0.155672
R388 VTAIL.n104 VTAIL.n103 0.155672
R389 VTAIL.n103 VTAIL.n95 0.155672
R390 VTAIL.n79 VTAIL.n47 0.155672
R391 VTAIL.n72 VTAIL.n47 0.155672
R392 VTAIL.n72 VTAIL.n71 0.155672
R393 VTAIL.n71 VTAIL.n51 0.155672
R394 VTAIL.n64 VTAIL.n51 0.155672
R395 VTAIL.n64 VTAIL.n63 0.155672
R396 VTAIL.n63 VTAIL.n55 0.155672
R397 VDD2.n70 VDD2.n69 585
R398 VDD2.n68 VDD2.n67 585
R399 VDD2.n43 VDD2.n42 585
R400 VDD2.n62 VDD2.n61 585
R401 VDD2.n60 VDD2.n59 585
R402 VDD2.n47 VDD2.n46 585
R403 VDD2.n54 VDD2.n53 585
R404 VDD2.n52 VDD2.n51 585
R405 VDD2.n13 VDD2.n12 585
R406 VDD2.n15 VDD2.n14 585
R407 VDD2.n8 VDD2.n7 585
R408 VDD2.n21 VDD2.n20 585
R409 VDD2.n23 VDD2.n22 585
R410 VDD2.n4 VDD2.n3 585
R411 VDD2.n29 VDD2.n28 585
R412 VDD2.n31 VDD2.n30 585
R413 VDD2.n69 VDD2.n39 498.474
R414 VDD2.n30 VDD2.n0 498.474
R415 VDD2.n50 VDD2.t1 329.053
R416 VDD2.n11 VDD2.t0 329.053
R417 VDD2.n69 VDD2.n68 171.744
R418 VDD2.n68 VDD2.n42 171.744
R419 VDD2.n61 VDD2.n42 171.744
R420 VDD2.n61 VDD2.n60 171.744
R421 VDD2.n60 VDD2.n46 171.744
R422 VDD2.n53 VDD2.n46 171.744
R423 VDD2.n53 VDD2.n52 171.744
R424 VDD2.n14 VDD2.n13 171.744
R425 VDD2.n14 VDD2.n7 171.744
R426 VDD2.n21 VDD2.n7 171.744
R427 VDD2.n22 VDD2.n21 171.744
R428 VDD2.n22 VDD2.n3 171.744
R429 VDD2.n29 VDD2.n3 171.744
R430 VDD2.n30 VDD2.n29 171.744
R431 VDD2.n38 VDD2.n37 88.6818
R432 VDD2 VDD2.n77 88.679
R433 VDD2.n76 VDD2.n75 86.5843
R434 VDD2.n36 VDD2.n35 86.5842
R435 VDD2.n52 VDD2.t1 85.8723
R436 VDD2.n13 VDD2.t0 85.8723
R437 VDD2.n36 VDD2.n34 53.4803
R438 VDD2.n74 VDD2.n73 50.6096
R439 VDD2.n74 VDD2.n38 43.5321
R440 VDD2.n71 VDD2.n70 12.8005
R441 VDD2.n32 VDD2.n31 12.8005
R442 VDD2.n67 VDD2.n41 12.0247
R443 VDD2.n28 VDD2.n2 12.0247
R444 VDD2.n66 VDD2.n43 11.249
R445 VDD2.n27 VDD2.n4 11.249
R446 VDD2.n51 VDD2.n50 10.7237
R447 VDD2.n12 VDD2.n11 10.7237
R448 VDD2.n63 VDD2.n62 10.4732
R449 VDD2.n24 VDD2.n23 10.4732
R450 VDD2.n59 VDD2.n45 9.69747
R451 VDD2.n20 VDD2.n6 9.69747
R452 VDD2.n73 VDD2.n72 9.45567
R453 VDD2.n34 VDD2.n33 9.45567
R454 VDD2.n49 VDD2.n48 9.3005
R455 VDD2.n56 VDD2.n55 9.3005
R456 VDD2.n58 VDD2.n57 9.3005
R457 VDD2.n45 VDD2.n44 9.3005
R458 VDD2.n64 VDD2.n63 9.3005
R459 VDD2.n66 VDD2.n65 9.3005
R460 VDD2.n41 VDD2.n40 9.3005
R461 VDD2.n72 VDD2.n71 9.3005
R462 VDD2.n10 VDD2.n9 9.3005
R463 VDD2.n17 VDD2.n16 9.3005
R464 VDD2.n19 VDD2.n18 9.3005
R465 VDD2.n6 VDD2.n5 9.3005
R466 VDD2.n25 VDD2.n24 9.3005
R467 VDD2.n27 VDD2.n26 9.3005
R468 VDD2.n2 VDD2.n1 9.3005
R469 VDD2.n33 VDD2.n32 9.3005
R470 VDD2.n58 VDD2.n47 8.92171
R471 VDD2.n19 VDD2.n8 8.92171
R472 VDD2.n55 VDD2.n54 8.14595
R473 VDD2.n16 VDD2.n15 8.14595
R474 VDD2.n73 VDD2.n39 7.75445
R475 VDD2.n34 VDD2.n0 7.75445
R476 VDD2.n51 VDD2.n49 7.3702
R477 VDD2.n12 VDD2.n10 7.3702
R478 VDD2.n71 VDD2.n39 6.08283
R479 VDD2.n32 VDD2.n0 6.08283
R480 VDD2.n54 VDD2.n49 5.81868
R481 VDD2.n15 VDD2.n10 5.81868
R482 VDD2.n55 VDD2.n47 5.04292
R483 VDD2.n16 VDD2.n8 5.04292
R484 VDD2.n77 VDD2.t5 4.53397
R485 VDD2.n77 VDD2.t6 4.53397
R486 VDD2.n75 VDD2.t2 4.53397
R487 VDD2.n75 VDD2.t8 4.53397
R488 VDD2.n37 VDD2.t3 4.53397
R489 VDD2.n37 VDD2.t9 4.53397
R490 VDD2.n35 VDD2.t4 4.53397
R491 VDD2.n35 VDD2.t7 4.53397
R492 VDD2.n59 VDD2.n58 4.26717
R493 VDD2.n20 VDD2.n19 4.26717
R494 VDD2.n62 VDD2.n45 3.49141
R495 VDD2.n23 VDD2.n6 3.49141
R496 VDD2.n76 VDD2.n74 2.87119
R497 VDD2.n63 VDD2.n43 2.71565
R498 VDD2.n24 VDD2.n4 2.71565
R499 VDD2.n50 VDD2.n48 2.41305
R500 VDD2.n11 VDD2.n9 2.41305
R501 VDD2.n67 VDD2.n66 1.93989
R502 VDD2.n28 VDD2.n27 1.93989
R503 VDD2.n70 VDD2.n41 1.16414
R504 VDD2.n31 VDD2.n2 1.16414
R505 VDD2 VDD2.n76 0.776362
R506 VDD2.n38 VDD2.n36 0.662826
R507 VDD2.n72 VDD2.n40 0.155672
R508 VDD2.n65 VDD2.n40 0.155672
R509 VDD2.n65 VDD2.n64 0.155672
R510 VDD2.n64 VDD2.n44 0.155672
R511 VDD2.n57 VDD2.n44 0.155672
R512 VDD2.n57 VDD2.n56 0.155672
R513 VDD2.n56 VDD2.n48 0.155672
R514 VDD2.n17 VDD2.n9 0.155672
R515 VDD2.n18 VDD2.n17 0.155672
R516 VDD2.n18 VDD2.n5 0.155672
R517 VDD2.n25 VDD2.n5 0.155672
R518 VDD2.n26 VDD2.n25 0.155672
R519 VDD2.n26 VDD2.n1 0.155672
R520 VDD2.n33 VDD2.n1 0.155672
R521 B.n609 B.n608 585
R522 B.n610 B.n71 585
R523 B.n612 B.n611 585
R524 B.n613 B.n70 585
R525 B.n615 B.n614 585
R526 B.n616 B.n69 585
R527 B.n618 B.n617 585
R528 B.n619 B.n68 585
R529 B.n621 B.n620 585
R530 B.n622 B.n67 585
R531 B.n624 B.n623 585
R532 B.n625 B.n66 585
R533 B.n627 B.n626 585
R534 B.n628 B.n65 585
R535 B.n630 B.n629 585
R536 B.n631 B.n64 585
R537 B.n633 B.n632 585
R538 B.n634 B.n63 585
R539 B.n636 B.n635 585
R540 B.n637 B.n62 585
R541 B.n639 B.n638 585
R542 B.n640 B.n61 585
R543 B.n642 B.n641 585
R544 B.n643 B.n60 585
R545 B.n645 B.n644 585
R546 B.n646 B.n59 585
R547 B.n648 B.n647 585
R548 B.n650 B.n649 585
R549 B.n651 B.n55 585
R550 B.n653 B.n652 585
R551 B.n654 B.n54 585
R552 B.n656 B.n655 585
R553 B.n657 B.n53 585
R554 B.n659 B.n658 585
R555 B.n660 B.n52 585
R556 B.n662 B.n661 585
R557 B.n663 B.n49 585
R558 B.n666 B.n665 585
R559 B.n667 B.n48 585
R560 B.n669 B.n668 585
R561 B.n670 B.n47 585
R562 B.n672 B.n671 585
R563 B.n673 B.n46 585
R564 B.n675 B.n674 585
R565 B.n676 B.n45 585
R566 B.n678 B.n677 585
R567 B.n679 B.n44 585
R568 B.n681 B.n680 585
R569 B.n682 B.n43 585
R570 B.n684 B.n683 585
R571 B.n685 B.n42 585
R572 B.n687 B.n686 585
R573 B.n688 B.n41 585
R574 B.n690 B.n689 585
R575 B.n691 B.n40 585
R576 B.n693 B.n692 585
R577 B.n694 B.n39 585
R578 B.n696 B.n695 585
R579 B.n697 B.n38 585
R580 B.n699 B.n698 585
R581 B.n700 B.n37 585
R582 B.n702 B.n701 585
R583 B.n703 B.n36 585
R584 B.n705 B.n704 585
R585 B.n607 B.n72 585
R586 B.n606 B.n605 585
R587 B.n604 B.n73 585
R588 B.n603 B.n602 585
R589 B.n601 B.n74 585
R590 B.n600 B.n599 585
R591 B.n598 B.n75 585
R592 B.n597 B.n596 585
R593 B.n595 B.n76 585
R594 B.n594 B.n593 585
R595 B.n592 B.n77 585
R596 B.n591 B.n590 585
R597 B.n589 B.n78 585
R598 B.n588 B.n587 585
R599 B.n586 B.n79 585
R600 B.n585 B.n584 585
R601 B.n583 B.n80 585
R602 B.n582 B.n581 585
R603 B.n580 B.n81 585
R604 B.n579 B.n578 585
R605 B.n577 B.n82 585
R606 B.n576 B.n575 585
R607 B.n574 B.n83 585
R608 B.n573 B.n572 585
R609 B.n571 B.n84 585
R610 B.n570 B.n569 585
R611 B.n568 B.n85 585
R612 B.n567 B.n566 585
R613 B.n565 B.n86 585
R614 B.n564 B.n563 585
R615 B.n562 B.n87 585
R616 B.n561 B.n560 585
R617 B.n559 B.n88 585
R618 B.n558 B.n557 585
R619 B.n556 B.n89 585
R620 B.n555 B.n554 585
R621 B.n553 B.n90 585
R622 B.n552 B.n551 585
R623 B.n550 B.n91 585
R624 B.n549 B.n548 585
R625 B.n547 B.n92 585
R626 B.n546 B.n545 585
R627 B.n544 B.n93 585
R628 B.n543 B.n542 585
R629 B.n541 B.n94 585
R630 B.n540 B.n539 585
R631 B.n538 B.n95 585
R632 B.n537 B.n536 585
R633 B.n535 B.n96 585
R634 B.n534 B.n533 585
R635 B.n532 B.n97 585
R636 B.n531 B.n530 585
R637 B.n529 B.n98 585
R638 B.n528 B.n527 585
R639 B.n526 B.n99 585
R640 B.n525 B.n524 585
R641 B.n523 B.n100 585
R642 B.n522 B.n521 585
R643 B.n520 B.n101 585
R644 B.n519 B.n518 585
R645 B.n517 B.n102 585
R646 B.n516 B.n515 585
R647 B.n514 B.n103 585
R648 B.n513 B.n512 585
R649 B.n511 B.n104 585
R650 B.n510 B.n509 585
R651 B.n508 B.n105 585
R652 B.n507 B.n506 585
R653 B.n505 B.n106 585
R654 B.n504 B.n503 585
R655 B.n502 B.n107 585
R656 B.n501 B.n500 585
R657 B.n499 B.n108 585
R658 B.n498 B.n497 585
R659 B.n496 B.n109 585
R660 B.n495 B.n494 585
R661 B.n493 B.n110 585
R662 B.n492 B.n491 585
R663 B.n490 B.n111 585
R664 B.n489 B.n488 585
R665 B.n487 B.n112 585
R666 B.n486 B.n485 585
R667 B.n484 B.n113 585
R668 B.n483 B.n482 585
R669 B.n481 B.n114 585
R670 B.n480 B.n479 585
R671 B.n478 B.n115 585
R672 B.n477 B.n476 585
R673 B.n475 B.n116 585
R674 B.n474 B.n473 585
R675 B.n472 B.n117 585
R676 B.n471 B.n470 585
R677 B.n469 B.n118 585
R678 B.n468 B.n467 585
R679 B.n466 B.n119 585
R680 B.n465 B.n464 585
R681 B.n463 B.n120 585
R682 B.n462 B.n461 585
R683 B.n460 B.n121 585
R684 B.n459 B.n458 585
R685 B.n457 B.n122 585
R686 B.n456 B.n455 585
R687 B.n454 B.n123 585
R688 B.n453 B.n452 585
R689 B.n451 B.n124 585
R690 B.n450 B.n449 585
R691 B.n448 B.n125 585
R692 B.n447 B.n446 585
R693 B.n445 B.n126 585
R694 B.n444 B.n443 585
R695 B.n442 B.n127 585
R696 B.n441 B.n440 585
R697 B.n439 B.n128 585
R698 B.n438 B.n437 585
R699 B.n436 B.n129 585
R700 B.n435 B.n434 585
R701 B.n433 B.n130 585
R702 B.n432 B.n431 585
R703 B.n430 B.n131 585
R704 B.n429 B.n428 585
R705 B.n427 B.n132 585
R706 B.n426 B.n425 585
R707 B.n424 B.n133 585
R708 B.n423 B.n422 585
R709 B.n421 B.n134 585
R710 B.n420 B.n419 585
R711 B.n418 B.n135 585
R712 B.n417 B.n416 585
R713 B.n415 B.n136 585
R714 B.n414 B.n413 585
R715 B.n412 B.n137 585
R716 B.n411 B.n410 585
R717 B.n409 B.n138 585
R718 B.n408 B.n407 585
R719 B.n406 B.n139 585
R720 B.n309 B.n308 585
R721 B.n310 B.n175 585
R722 B.n312 B.n311 585
R723 B.n313 B.n174 585
R724 B.n315 B.n314 585
R725 B.n316 B.n173 585
R726 B.n318 B.n317 585
R727 B.n319 B.n172 585
R728 B.n321 B.n320 585
R729 B.n322 B.n171 585
R730 B.n324 B.n323 585
R731 B.n325 B.n170 585
R732 B.n327 B.n326 585
R733 B.n328 B.n169 585
R734 B.n330 B.n329 585
R735 B.n331 B.n168 585
R736 B.n333 B.n332 585
R737 B.n334 B.n167 585
R738 B.n336 B.n335 585
R739 B.n337 B.n166 585
R740 B.n339 B.n338 585
R741 B.n340 B.n165 585
R742 B.n342 B.n341 585
R743 B.n343 B.n164 585
R744 B.n345 B.n344 585
R745 B.n346 B.n163 585
R746 B.n348 B.n347 585
R747 B.n350 B.n349 585
R748 B.n351 B.n159 585
R749 B.n353 B.n352 585
R750 B.n354 B.n158 585
R751 B.n356 B.n355 585
R752 B.n357 B.n157 585
R753 B.n359 B.n358 585
R754 B.n360 B.n156 585
R755 B.n362 B.n361 585
R756 B.n363 B.n153 585
R757 B.n366 B.n365 585
R758 B.n367 B.n152 585
R759 B.n369 B.n368 585
R760 B.n370 B.n151 585
R761 B.n372 B.n371 585
R762 B.n373 B.n150 585
R763 B.n375 B.n374 585
R764 B.n376 B.n149 585
R765 B.n378 B.n377 585
R766 B.n379 B.n148 585
R767 B.n381 B.n380 585
R768 B.n382 B.n147 585
R769 B.n384 B.n383 585
R770 B.n385 B.n146 585
R771 B.n387 B.n386 585
R772 B.n388 B.n145 585
R773 B.n390 B.n389 585
R774 B.n391 B.n144 585
R775 B.n393 B.n392 585
R776 B.n394 B.n143 585
R777 B.n396 B.n395 585
R778 B.n397 B.n142 585
R779 B.n399 B.n398 585
R780 B.n400 B.n141 585
R781 B.n402 B.n401 585
R782 B.n403 B.n140 585
R783 B.n405 B.n404 585
R784 B.n307 B.n176 585
R785 B.n306 B.n305 585
R786 B.n304 B.n177 585
R787 B.n303 B.n302 585
R788 B.n301 B.n178 585
R789 B.n300 B.n299 585
R790 B.n298 B.n179 585
R791 B.n297 B.n296 585
R792 B.n295 B.n180 585
R793 B.n294 B.n293 585
R794 B.n292 B.n181 585
R795 B.n291 B.n290 585
R796 B.n289 B.n182 585
R797 B.n288 B.n287 585
R798 B.n286 B.n183 585
R799 B.n285 B.n284 585
R800 B.n283 B.n184 585
R801 B.n282 B.n281 585
R802 B.n280 B.n185 585
R803 B.n279 B.n278 585
R804 B.n277 B.n186 585
R805 B.n276 B.n275 585
R806 B.n274 B.n187 585
R807 B.n273 B.n272 585
R808 B.n271 B.n188 585
R809 B.n270 B.n269 585
R810 B.n268 B.n189 585
R811 B.n267 B.n266 585
R812 B.n265 B.n190 585
R813 B.n264 B.n263 585
R814 B.n262 B.n191 585
R815 B.n261 B.n260 585
R816 B.n259 B.n192 585
R817 B.n258 B.n257 585
R818 B.n256 B.n193 585
R819 B.n255 B.n254 585
R820 B.n253 B.n194 585
R821 B.n252 B.n251 585
R822 B.n250 B.n195 585
R823 B.n249 B.n248 585
R824 B.n247 B.n196 585
R825 B.n246 B.n245 585
R826 B.n244 B.n197 585
R827 B.n243 B.n242 585
R828 B.n241 B.n198 585
R829 B.n240 B.n239 585
R830 B.n238 B.n199 585
R831 B.n237 B.n236 585
R832 B.n235 B.n200 585
R833 B.n234 B.n233 585
R834 B.n232 B.n201 585
R835 B.n231 B.n230 585
R836 B.n229 B.n202 585
R837 B.n228 B.n227 585
R838 B.n226 B.n203 585
R839 B.n225 B.n224 585
R840 B.n223 B.n204 585
R841 B.n222 B.n221 585
R842 B.n220 B.n205 585
R843 B.n219 B.n218 585
R844 B.n217 B.n206 585
R845 B.n216 B.n215 585
R846 B.n214 B.n207 585
R847 B.n213 B.n212 585
R848 B.n211 B.n208 585
R849 B.n210 B.n209 585
R850 B.n2 B.n0 585
R851 B.n805 B.n1 585
R852 B.n804 B.n803 585
R853 B.n802 B.n3 585
R854 B.n801 B.n800 585
R855 B.n799 B.n4 585
R856 B.n798 B.n797 585
R857 B.n796 B.n5 585
R858 B.n795 B.n794 585
R859 B.n793 B.n6 585
R860 B.n792 B.n791 585
R861 B.n790 B.n7 585
R862 B.n789 B.n788 585
R863 B.n787 B.n8 585
R864 B.n786 B.n785 585
R865 B.n784 B.n9 585
R866 B.n783 B.n782 585
R867 B.n781 B.n10 585
R868 B.n780 B.n779 585
R869 B.n778 B.n11 585
R870 B.n777 B.n776 585
R871 B.n775 B.n12 585
R872 B.n774 B.n773 585
R873 B.n772 B.n13 585
R874 B.n771 B.n770 585
R875 B.n769 B.n14 585
R876 B.n768 B.n767 585
R877 B.n766 B.n15 585
R878 B.n765 B.n764 585
R879 B.n763 B.n16 585
R880 B.n762 B.n761 585
R881 B.n760 B.n17 585
R882 B.n759 B.n758 585
R883 B.n757 B.n18 585
R884 B.n756 B.n755 585
R885 B.n754 B.n19 585
R886 B.n753 B.n752 585
R887 B.n751 B.n20 585
R888 B.n750 B.n749 585
R889 B.n748 B.n21 585
R890 B.n747 B.n746 585
R891 B.n745 B.n22 585
R892 B.n744 B.n743 585
R893 B.n742 B.n23 585
R894 B.n741 B.n740 585
R895 B.n739 B.n24 585
R896 B.n738 B.n737 585
R897 B.n736 B.n25 585
R898 B.n735 B.n734 585
R899 B.n733 B.n26 585
R900 B.n732 B.n731 585
R901 B.n730 B.n27 585
R902 B.n729 B.n728 585
R903 B.n727 B.n28 585
R904 B.n726 B.n725 585
R905 B.n724 B.n29 585
R906 B.n723 B.n722 585
R907 B.n721 B.n30 585
R908 B.n720 B.n719 585
R909 B.n718 B.n31 585
R910 B.n717 B.n716 585
R911 B.n715 B.n32 585
R912 B.n714 B.n713 585
R913 B.n712 B.n33 585
R914 B.n711 B.n710 585
R915 B.n709 B.n34 585
R916 B.n708 B.n707 585
R917 B.n706 B.n35 585
R918 B.n807 B.n806 585
R919 B.n308 B.n307 511.721
R920 B.n704 B.n35 511.721
R921 B.n404 B.n139 511.721
R922 B.n608 B.n607 511.721
R923 B.n154 B.t2 353.192
R924 B.n56 B.t10 353.192
R925 B.n160 B.t5 353.192
R926 B.n50 B.t7 353.192
R927 B.n155 B.t1 288.611
R928 B.n57 B.t11 288.611
R929 B.n161 B.t4 288.611
R930 B.n51 B.t8 288.611
R931 B.n154 B.t0 266.18
R932 B.n160 B.t3 266.18
R933 B.n50 B.t6 266.18
R934 B.n56 B.t9 266.18
R935 B.n307 B.n306 163.367
R936 B.n306 B.n177 163.367
R937 B.n302 B.n177 163.367
R938 B.n302 B.n301 163.367
R939 B.n301 B.n300 163.367
R940 B.n300 B.n179 163.367
R941 B.n296 B.n179 163.367
R942 B.n296 B.n295 163.367
R943 B.n295 B.n294 163.367
R944 B.n294 B.n181 163.367
R945 B.n290 B.n181 163.367
R946 B.n290 B.n289 163.367
R947 B.n289 B.n288 163.367
R948 B.n288 B.n183 163.367
R949 B.n284 B.n183 163.367
R950 B.n284 B.n283 163.367
R951 B.n283 B.n282 163.367
R952 B.n282 B.n185 163.367
R953 B.n278 B.n185 163.367
R954 B.n278 B.n277 163.367
R955 B.n277 B.n276 163.367
R956 B.n276 B.n187 163.367
R957 B.n272 B.n187 163.367
R958 B.n272 B.n271 163.367
R959 B.n271 B.n270 163.367
R960 B.n270 B.n189 163.367
R961 B.n266 B.n189 163.367
R962 B.n266 B.n265 163.367
R963 B.n265 B.n264 163.367
R964 B.n264 B.n191 163.367
R965 B.n260 B.n191 163.367
R966 B.n260 B.n259 163.367
R967 B.n259 B.n258 163.367
R968 B.n258 B.n193 163.367
R969 B.n254 B.n193 163.367
R970 B.n254 B.n253 163.367
R971 B.n253 B.n252 163.367
R972 B.n252 B.n195 163.367
R973 B.n248 B.n195 163.367
R974 B.n248 B.n247 163.367
R975 B.n247 B.n246 163.367
R976 B.n246 B.n197 163.367
R977 B.n242 B.n197 163.367
R978 B.n242 B.n241 163.367
R979 B.n241 B.n240 163.367
R980 B.n240 B.n199 163.367
R981 B.n236 B.n199 163.367
R982 B.n236 B.n235 163.367
R983 B.n235 B.n234 163.367
R984 B.n234 B.n201 163.367
R985 B.n230 B.n201 163.367
R986 B.n230 B.n229 163.367
R987 B.n229 B.n228 163.367
R988 B.n228 B.n203 163.367
R989 B.n224 B.n203 163.367
R990 B.n224 B.n223 163.367
R991 B.n223 B.n222 163.367
R992 B.n222 B.n205 163.367
R993 B.n218 B.n205 163.367
R994 B.n218 B.n217 163.367
R995 B.n217 B.n216 163.367
R996 B.n216 B.n207 163.367
R997 B.n212 B.n207 163.367
R998 B.n212 B.n211 163.367
R999 B.n211 B.n210 163.367
R1000 B.n210 B.n2 163.367
R1001 B.n806 B.n2 163.367
R1002 B.n806 B.n805 163.367
R1003 B.n805 B.n804 163.367
R1004 B.n804 B.n3 163.367
R1005 B.n800 B.n3 163.367
R1006 B.n800 B.n799 163.367
R1007 B.n799 B.n798 163.367
R1008 B.n798 B.n5 163.367
R1009 B.n794 B.n5 163.367
R1010 B.n794 B.n793 163.367
R1011 B.n793 B.n792 163.367
R1012 B.n792 B.n7 163.367
R1013 B.n788 B.n7 163.367
R1014 B.n788 B.n787 163.367
R1015 B.n787 B.n786 163.367
R1016 B.n786 B.n9 163.367
R1017 B.n782 B.n9 163.367
R1018 B.n782 B.n781 163.367
R1019 B.n781 B.n780 163.367
R1020 B.n780 B.n11 163.367
R1021 B.n776 B.n11 163.367
R1022 B.n776 B.n775 163.367
R1023 B.n775 B.n774 163.367
R1024 B.n774 B.n13 163.367
R1025 B.n770 B.n13 163.367
R1026 B.n770 B.n769 163.367
R1027 B.n769 B.n768 163.367
R1028 B.n768 B.n15 163.367
R1029 B.n764 B.n15 163.367
R1030 B.n764 B.n763 163.367
R1031 B.n763 B.n762 163.367
R1032 B.n762 B.n17 163.367
R1033 B.n758 B.n17 163.367
R1034 B.n758 B.n757 163.367
R1035 B.n757 B.n756 163.367
R1036 B.n756 B.n19 163.367
R1037 B.n752 B.n19 163.367
R1038 B.n752 B.n751 163.367
R1039 B.n751 B.n750 163.367
R1040 B.n750 B.n21 163.367
R1041 B.n746 B.n21 163.367
R1042 B.n746 B.n745 163.367
R1043 B.n745 B.n744 163.367
R1044 B.n744 B.n23 163.367
R1045 B.n740 B.n23 163.367
R1046 B.n740 B.n739 163.367
R1047 B.n739 B.n738 163.367
R1048 B.n738 B.n25 163.367
R1049 B.n734 B.n25 163.367
R1050 B.n734 B.n733 163.367
R1051 B.n733 B.n732 163.367
R1052 B.n732 B.n27 163.367
R1053 B.n728 B.n27 163.367
R1054 B.n728 B.n727 163.367
R1055 B.n727 B.n726 163.367
R1056 B.n726 B.n29 163.367
R1057 B.n722 B.n29 163.367
R1058 B.n722 B.n721 163.367
R1059 B.n721 B.n720 163.367
R1060 B.n720 B.n31 163.367
R1061 B.n716 B.n31 163.367
R1062 B.n716 B.n715 163.367
R1063 B.n715 B.n714 163.367
R1064 B.n714 B.n33 163.367
R1065 B.n710 B.n33 163.367
R1066 B.n710 B.n709 163.367
R1067 B.n709 B.n708 163.367
R1068 B.n708 B.n35 163.367
R1069 B.n308 B.n175 163.367
R1070 B.n312 B.n175 163.367
R1071 B.n313 B.n312 163.367
R1072 B.n314 B.n313 163.367
R1073 B.n314 B.n173 163.367
R1074 B.n318 B.n173 163.367
R1075 B.n319 B.n318 163.367
R1076 B.n320 B.n319 163.367
R1077 B.n320 B.n171 163.367
R1078 B.n324 B.n171 163.367
R1079 B.n325 B.n324 163.367
R1080 B.n326 B.n325 163.367
R1081 B.n326 B.n169 163.367
R1082 B.n330 B.n169 163.367
R1083 B.n331 B.n330 163.367
R1084 B.n332 B.n331 163.367
R1085 B.n332 B.n167 163.367
R1086 B.n336 B.n167 163.367
R1087 B.n337 B.n336 163.367
R1088 B.n338 B.n337 163.367
R1089 B.n338 B.n165 163.367
R1090 B.n342 B.n165 163.367
R1091 B.n343 B.n342 163.367
R1092 B.n344 B.n343 163.367
R1093 B.n344 B.n163 163.367
R1094 B.n348 B.n163 163.367
R1095 B.n349 B.n348 163.367
R1096 B.n349 B.n159 163.367
R1097 B.n353 B.n159 163.367
R1098 B.n354 B.n353 163.367
R1099 B.n355 B.n354 163.367
R1100 B.n355 B.n157 163.367
R1101 B.n359 B.n157 163.367
R1102 B.n360 B.n359 163.367
R1103 B.n361 B.n360 163.367
R1104 B.n361 B.n153 163.367
R1105 B.n366 B.n153 163.367
R1106 B.n367 B.n366 163.367
R1107 B.n368 B.n367 163.367
R1108 B.n368 B.n151 163.367
R1109 B.n372 B.n151 163.367
R1110 B.n373 B.n372 163.367
R1111 B.n374 B.n373 163.367
R1112 B.n374 B.n149 163.367
R1113 B.n378 B.n149 163.367
R1114 B.n379 B.n378 163.367
R1115 B.n380 B.n379 163.367
R1116 B.n380 B.n147 163.367
R1117 B.n384 B.n147 163.367
R1118 B.n385 B.n384 163.367
R1119 B.n386 B.n385 163.367
R1120 B.n386 B.n145 163.367
R1121 B.n390 B.n145 163.367
R1122 B.n391 B.n390 163.367
R1123 B.n392 B.n391 163.367
R1124 B.n392 B.n143 163.367
R1125 B.n396 B.n143 163.367
R1126 B.n397 B.n396 163.367
R1127 B.n398 B.n397 163.367
R1128 B.n398 B.n141 163.367
R1129 B.n402 B.n141 163.367
R1130 B.n403 B.n402 163.367
R1131 B.n404 B.n403 163.367
R1132 B.n408 B.n139 163.367
R1133 B.n409 B.n408 163.367
R1134 B.n410 B.n409 163.367
R1135 B.n410 B.n137 163.367
R1136 B.n414 B.n137 163.367
R1137 B.n415 B.n414 163.367
R1138 B.n416 B.n415 163.367
R1139 B.n416 B.n135 163.367
R1140 B.n420 B.n135 163.367
R1141 B.n421 B.n420 163.367
R1142 B.n422 B.n421 163.367
R1143 B.n422 B.n133 163.367
R1144 B.n426 B.n133 163.367
R1145 B.n427 B.n426 163.367
R1146 B.n428 B.n427 163.367
R1147 B.n428 B.n131 163.367
R1148 B.n432 B.n131 163.367
R1149 B.n433 B.n432 163.367
R1150 B.n434 B.n433 163.367
R1151 B.n434 B.n129 163.367
R1152 B.n438 B.n129 163.367
R1153 B.n439 B.n438 163.367
R1154 B.n440 B.n439 163.367
R1155 B.n440 B.n127 163.367
R1156 B.n444 B.n127 163.367
R1157 B.n445 B.n444 163.367
R1158 B.n446 B.n445 163.367
R1159 B.n446 B.n125 163.367
R1160 B.n450 B.n125 163.367
R1161 B.n451 B.n450 163.367
R1162 B.n452 B.n451 163.367
R1163 B.n452 B.n123 163.367
R1164 B.n456 B.n123 163.367
R1165 B.n457 B.n456 163.367
R1166 B.n458 B.n457 163.367
R1167 B.n458 B.n121 163.367
R1168 B.n462 B.n121 163.367
R1169 B.n463 B.n462 163.367
R1170 B.n464 B.n463 163.367
R1171 B.n464 B.n119 163.367
R1172 B.n468 B.n119 163.367
R1173 B.n469 B.n468 163.367
R1174 B.n470 B.n469 163.367
R1175 B.n470 B.n117 163.367
R1176 B.n474 B.n117 163.367
R1177 B.n475 B.n474 163.367
R1178 B.n476 B.n475 163.367
R1179 B.n476 B.n115 163.367
R1180 B.n480 B.n115 163.367
R1181 B.n481 B.n480 163.367
R1182 B.n482 B.n481 163.367
R1183 B.n482 B.n113 163.367
R1184 B.n486 B.n113 163.367
R1185 B.n487 B.n486 163.367
R1186 B.n488 B.n487 163.367
R1187 B.n488 B.n111 163.367
R1188 B.n492 B.n111 163.367
R1189 B.n493 B.n492 163.367
R1190 B.n494 B.n493 163.367
R1191 B.n494 B.n109 163.367
R1192 B.n498 B.n109 163.367
R1193 B.n499 B.n498 163.367
R1194 B.n500 B.n499 163.367
R1195 B.n500 B.n107 163.367
R1196 B.n504 B.n107 163.367
R1197 B.n505 B.n504 163.367
R1198 B.n506 B.n505 163.367
R1199 B.n506 B.n105 163.367
R1200 B.n510 B.n105 163.367
R1201 B.n511 B.n510 163.367
R1202 B.n512 B.n511 163.367
R1203 B.n512 B.n103 163.367
R1204 B.n516 B.n103 163.367
R1205 B.n517 B.n516 163.367
R1206 B.n518 B.n517 163.367
R1207 B.n518 B.n101 163.367
R1208 B.n522 B.n101 163.367
R1209 B.n523 B.n522 163.367
R1210 B.n524 B.n523 163.367
R1211 B.n524 B.n99 163.367
R1212 B.n528 B.n99 163.367
R1213 B.n529 B.n528 163.367
R1214 B.n530 B.n529 163.367
R1215 B.n530 B.n97 163.367
R1216 B.n534 B.n97 163.367
R1217 B.n535 B.n534 163.367
R1218 B.n536 B.n535 163.367
R1219 B.n536 B.n95 163.367
R1220 B.n540 B.n95 163.367
R1221 B.n541 B.n540 163.367
R1222 B.n542 B.n541 163.367
R1223 B.n542 B.n93 163.367
R1224 B.n546 B.n93 163.367
R1225 B.n547 B.n546 163.367
R1226 B.n548 B.n547 163.367
R1227 B.n548 B.n91 163.367
R1228 B.n552 B.n91 163.367
R1229 B.n553 B.n552 163.367
R1230 B.n554 B.n553 163.367
R1231 B.n554 B.n89 163.367
R1232 B.n558 B.n89 163.367
R1233 B.n559 B.n558 163.367
R1234 B.n560 B.n559 163.367
R1235 B.n560 B.n87 163.367
R1236 B.n564 B.n87 163.367
R1237 B.n565 B.n564 163.367
R1238 B.n566 B.n565 163.367
R1239 B.n566 B.n85 163.367
R1240 B.n570 B.n85 163.367
R1241 B.n571 B.n570 163.367
R1242 B.n572 B.n571 163.367
R1243 B.n572 B.n83 163.367
R1244 B.n576 B.n83 163.367
R1245 B.n577 B.n576 163.367
R1246 B.n578 B.n577 163.367
R1247 B.n578 B.n81 163.367
R1248 B.n582 B.n81 163.367
R1249 B.n583 B.n582 163.367
R1250 B.n584 B.n583 163.367
R1251 B.n584 B.n79 163.367
R1252 B.n588 B.n79 163.367
R1253 B.n589 B.n588 163.367
R1254 B.n590 B.n589 163.367
R1255 B.n590 B.n77 163.367
R1256 B.n594 B.n77 163.367
R1257 B.n595 B.n594 163.367
R1258 B.n596 B.n595 163.367
R1259 B.n596 B.n75 163.367
R1260 B.n600 B.n75 163.367
R1261 B.n601 B.n600 163.367
R1262 B.n602 B.n601 163.367
R1263 B.n602 B.n73 163.367
R1264 B.n606 B.n73 163.367
R1265 B.n607 B.n606 163.367
R1266 B.n704 B.n703 163.367
R1267 B.n703 B.n702 163.367
R1268 B.n702 B.n37 163.367
R1269 B.n698 B.n37 163.367
R1270 B.n698 B.n697 163.367
R1271 B.n697 B.n696 163.367
R1272 B.n696 B.n39 163.367
R1273 B.n692 B.n39 163.367
R1274 B.n692 B.n691 163.367
R1275 B.n691 B.n690 163.367
R1276 B.n690 B.n41 163.367
R1277 B.n686 B.n41 163.367
R1278 B.n686 B.n685 163.367
R1279 B.n685 B.n684 163.367
R1280 B.n684 B.n43 163.367
R1281 B.n680 B.n43 163.367
R1282 B.n680 B.n679 163.367
R1283 B.n679 B.n678 163.367
R1284 B.n678 B.n45 163.367
R1285 B.n674 B.n45 163.367
R1286 B.n674 B.n673 163.367
R1287 B.n673 B.n672 163.367
R1288 B.n672 B.n47 163.367
R1289 B.n668 B.n47 163.367
R1290 B.n668 B.n667 163.367
R1291 B.n667 B.n666 163.367
R1292 B.n666 B.n49 163.367
R1293 B.n661 B.n49 163.367
R1294 B.n661 B.n660 163.367
R1295 B.n660 B.n659 163.367
R1296 B.n659 B.n53 163.367
R1297 B.n655 B.n53 163.367
R1298 B.n655 B.n654 163.367
R1299 B.n654 B.n653 163.367
R1300 B.n653 B.n55 163.367
R1301 B.n649 B.n55 163.367
R1302 B.n649 B.n648 163.367
R1303 B.n648 B.n59 163.367
R1304 B.n644 B.n59 163.367
R1305 B.n644 B.n643 163.367
R1306 B.n643 B.n642 163.367
R1307 B.n642 B.n61 163.367
R1308 B.n638 B.n61 163.367
R1309 B.n638 B.n637 163.367
R1310 B.n637 B.n636 163.367
R1311 B.n636 B.n63 163.367
R1312 B.n632 B.n63 163.367
R1313 B.n632 B.n631 163.367
R1314 B.n631 B.n630 163.367
R1315 B.n630 B.n65 163.367
R1316 B.n626 B.n65 163.367
R1317 B.n626 B.n625 163.367
R1318 B.n625 B.n624 163.367
R1319 B.n624 B.n67 163.367
R1320 B.n620 B.n67 163.367
R1321 B.n620 B.n619 163.367
R1322 B.n619 B.n618 163.367
R1323 B.n618 B.n69 163.367
R1324 B.n614 B.n69 163.367
R1325 B.n614 B.n613 163.367
R1326 B.n613 B.n612 163.367
R1327 B.n612 B.n71 163.367
R1328 B.n608 B.n71 163.367
R1329 B.n155 B.n154 64.5823
R1330 B.n161 B.n160 64.5823
R1331 B.n51 B.n50 64.5823
R1332 B.n57 B.n56 64.5823
R1333 B.n364 B.n155 59.5399
R1334 B.n162 B.n161 59.5399
R1335 B.n664 B.n51 59.5399
R1336 B.n58 B.n57 59.5399
R1337 B.n706 B.n705 33.2493
R1338 B.n609 B.n72 33.2493
R1339 B.n406 B.n405 33.2493
R1340 B.n309 B.n176 33.2493
R1341 B B.n807 18.0485
R1342 B.n705 B.n36 10.6151
R1343 B.n701 B.n36 10.6151
R1344 B.n701 B.n700 10.6151
R1345 B.n700 B.n699 10.6151
R1346 B.n699 B.n38 10.6151
R1347 B.n695 B.n38 10.6151
R1348 B.n695 B.n694 10.6151
R1349 B.n694 B.n693 10.6151
R1350 B.n693 B.n40 10.6151
R1351 B.n689 B.n40 10.6151
R1352 B.n689 B.n688 10.6151
R1353 B.n688 B.n687 10.6151
R1354 B.n687 B.n42 10.6151
R1355 B.n683 B.n42 10.6151
R1356 B.n683 B.n682 10.6151
R1357 B.n682 B.n681 10.6151
R1358 B.n681 B.n44 10.6151
R1359 B.n677 B.n44 10.6151
R1360 B.n677 B.n676 10.6151
R1361 B.n676 B.n675 10.6151
R1362 B.n675 B.n46 10.6151
R1363 B.n671 B.n46 10.6151
R1364 B.n671 B.n670 10.6151
R1365 B.n670 B.n669 10.6151
R1366 B.n669 B.n48 10.6151
R1367 B.n665 B.n48 10.6151
R1368 B.n663 B.n662 10.6151
R1369 B.n662 B.n52 10.6151
R1370 B.n658 B.n52 10.6151
R1371 B.n658 B.n657 10.6151
R1372 B.n657 B.n656 10.6151
R1373 B.n656 B.n54 10.6151
R1374 B.n652 B.n54 10.6151
R1375 B.n652 B.n651 10.6151
R1376 B.n651 B.n650 10.6151
R1377 B.n647 B.n646 10.6151
R1378 B.n646 B.n645 10.6151
R1379 B.n645 B.n60 10.6151
R1380 B.n641 B.n60 10.6151
R1381 B.n641 B.n640 10.6151
R1382 B.n640 B.n639 10.6151
R1383 B.n639 B.n62 10.6151
R1384 B.n635 B.n62 10.6151
R1385 B.n635 B.n634 10.6151
R1386 B.n634 B.n633 10.6151
R1387 B.n633 B.n64 10.6151
R1388 B.n629 B.n64 10.6151
R1389 B.n629 B.n628 10.6151
R1390 B.n628 B.n627 10.6151
R1391 B.n627 B.n66 10.6151
R1392 B.n623 B.n66 10.6151
R1393 B.n623 B.n622 10.6151
R1394 B.n622 B.n621 10.6151
R1395 B.n621 B.n68 10.6151
R1396 B.n617 B.n68 10.6151
R1397 B.n617 B.n616 10.6151
R1398 B.n616 B.n615 10.6151
R1399 B.n615 B.n70 10.6151
R1400 B.n611 B.n70 10.6151
R1401 B.n611 B.n610 10.6151
R1402 B.n610 B.n609 10.6151
R1403 B.n407 B.n406 10.6151
R1404 B.n407 B.n138 10.6151
R1405 B.n411 B.n138 10.6151
R1406 B.n412 B.n411 10.6151
R1407 B.n413 B.n412 10.6151
R1408 B.n413 B.n136 10.6151
R1409 B.n417 B.n136 10.6151
R1410 B.n418 B.n417 10.6151
R1411 B.n419 B.n418 10.6151
R1412 B.n419 B.n134 10.6151
R1413 B.n423 B.n134 10.6151
R1414 B.n424 B.n423 10.6151
R1415 B.n425 B.n424 10.6151
R1416 B.n425 B.n132 10.6151
R1417 B.n429 B.n132 10.6151
R1418 B.n430 B.n429 10.6151
R1419 B.n431 B.n430 10.6151
R1420 B.n431 B.n130 10.6151
R1421 B.n435 B.n130 10.6151
R1422 B.n436 B.n435 10.6151
R1423 B.n437 B.n436 10.6151
R1424 B.n437 B.n128 10.6151
R1425 B.n441 B.n128 10.6151
R1426 B.n442 B.n441 10.6151
R1427 B.n443 B.n442 10.6151
R1428 B.n443 B.n126 10.6151
R1429 B.n447 B.n126 10.6151
R1430 B.n448 B.n447 10.6151
R1431 B.n449 B.n448 10.6151
R1432 B.n449 B.n124 10.6151
R1433 B.n453 B.n124 10.6151
R1434 B.n454 B.n453 10.6151
R1435 B.n455 B.n454 10.6151
R1436 B.n455 B.n122 10.6151
R1437 B.n459 B.n122 10.6151
R1438 B.n460 B.n459 10.6151
R1439 B.n461 B.n460 10.6151
R1440 B.n461 B.n120 10.6151
R1441 B.n465 B.n120 10.6151
R1442 B.n466 B.n465 10.6151
R1443 B.n467 B.n466 10.6151
R1444 B.n467 B.n118 10.6151
R1445 B.n471 B.n118 10.6151
R1446 B.n472 B.n471 10.6151
R1447 B.n473 B.n472 10.6151
R1448 B.n473 B.n116 10.6151
R1449 B.n477 B.n116 10.6151
R1450 B.n478 B.n477 10.6151
R1451 B.n479 B.n478 10.6151
R1452 B.n479 B.n114 10.6151
R1453 B.n483 B.n114 10.6151
R1454 B.n484 B.n483 10.6151
R1455 B.n485 B.n484 10.6151
R1456 B.n485 B.n112 10.6151
R1457 B.n489 B.n112 10.6151
R1458 B.n490 B.n489 10.6151
R1459 B.n491 B.n490 10.6151
R1460 B.n491 B.n110 10.6151
R1461 B.n495 B.n110 10.6151
R1462 B.n496 B.n495 10.6151
R1463 B.n497 B.n496 10.6151
R1464 B.n497 B.n108 10.6151
R1465 B.n501 B.n108 10.6151
R1466 B.n502 B.n501 10.6151
R1467 B.n503 B.n502 10.6151
R1468 B.n503 B.n106 10.6151
R1469 B.n507 B.n106 10.6151
R1470 B.n508 B.n507 10.6151
R1471 B.n509 B.n508 10.6151
R1472 B.n509 B.n104 10.6151
R1473 B.n513 B.n104 10.6151
R1474 B.n514 B.n513 10.6151
R1475 B.n515 B.n514 10.6151
R1476 B.n515 B.n102 10.6151
R1477 B.n519 B.n102 10.6151
R1478 B.n520 B.n519 10.6151
R1479 B.n521 B.n520 10.6151
R1480 B.n521 B.n100 10.6151
R1481 B.n525 B.n100 10.6151
R1482 B.n526 B.n525 10.6151
R1483 B.n527 B.n526 10.6151
R1484 B.n527 B.n98 10.6151
R1485 B.n531 B.n98 10.6151
R1486 B.n532 B.n531 10.6151
R1487 B.n533 B.n532 10.6151
R1488 B.n533 B.n96 10.6151
R1489 B.n537 B.n96 10.6151
R1490 B.n538 B.n537 10.6151
R1491 B.n539 B.n538 10.6151
R1492 B.n539 B.n94 10.6151
R1493 B.n543 B.n94 10.6151
R1494 B.n544 B.n543 10.6151
R1495 B.n545 B.n544 10.6151
R1496 B.n545 B.n92 10.6151
R1497 B.n549 B.n92 10.6151
R1498 B.n550 B.n549 10.6151
R1499 B.n551 B.n550 10.6151
R1500 B.n551 B.n90 10.6151
R1501 B.n555 B.n90 10.6151
R1502 B.n556 B.n555 10.6151
R1503 B.n557 B.n556 10.6151
R1504 B.n557 B.n88 10.6151
R1505 B.n561 B.n88 10.6151
R1506 B.n562 B.n561 10.6151
R1507 B.n563 B.n562 10.6151
R1508 B.n563 B.n86 10.6151
R1509 B.n567 B.n86 10.6151
R1510 B.n568 B.n567 10.6151
R1511 B.n569 B.n568 10.6151
R1512 B.n569 B.n84 10.6151
R1513 B.n573 B.n84 10.6151
R1514 B.n574 B.n573 10.6151
R1515 B.n575 B.n574 10.6151
R1516 B.n575 B.n82 10.6151
R1517 B.n579 B.n82 10.6151
R1518 B.n580 B.n579 10.6151
R1519 B.n581 B.n580 10.6151
R1520 B.n581 B.n80 10.6151
R1521 B.n585 B.n80 10.6151
R1522 B.n586 B.n585 10.6151
R1523 B.n587 B.n586 10.6151
R1524 B.n587 B.n78 10.6151
R1525 B.n591 B.n78 10.6151
R1526 B.n592 B.n591 10.6151
R1527 B.n593 B.n592 10.6151
R1528 B.n593 B.n76 10.6151
R1529 B.n597 B.n76 10.6151
R1530 B.n598 B.n597 10.6151
R1531 B.n599 B.n598 10.6151
R1532 B.n599 B.n74 10.6151
R1533 B.n603 B.n74 10.6151
R1534 B.n604 B.n603 10.6151
R1535 B.n605 B.n604 10.6151
R1536 B.n605 B.n72 10.6151
R1537 B.n310 B.n309 10.6151
R1538 B.n311 B.n310 10.6151
R1539 B.n311 B.n174 10.6151
R1540 B.n315 B.n174 10.6151
R1541 B.n316 B.n315 10.6151
R1542 B.n317 B.n316 10.6151
R1543 B.n317 B.n172 10.6151
R1544 B.n321 B.n172 10.6151
R1545 B.n322 B.n321 10.6151
R1546 B.n323 B.n322 10.6151
R1547 B.n323 B.n170 10.6151
R1548 B.n327 B.n170 10.6151
R1549 B.n328 B.n327 10.6151
R1550 B.n329 B.n328 10.6151
R1551 B.n329 B.n168 10.6151
R1552 B.n333 B.n168 10.6151
R1553 B.n334 B.n333 10.6151
R1554 B.n335 B.n334 10.6151
R1555 B.n335 B.n166 10.6151
R1556 B.n339 B.n166 10.6151
R1557 B.n340 B.n339 10.6151
R1558 B.n341 B.n340 10.6151
R1559 B.n341 B.n164 10.6151
R1560 B.n345 B.n164 10.6151
R1561 B.n346 B.n345 10.6151
R1562 B.n347 B.n346 10.6151
R1563 B.n351 B.n350 10.6151
R1564 B.n352 B.n351 10.6151
R1565 B.n352 B.n158 10.6151
R1566 B.n356 B.n158 10.6151
R1567 B.n357 B.n356 10.6151
R1568 B.n358 B.n357 10.6151
R1569 B.n358 B.n156 10.6151
R1570 B.n362 B.n156 10.6151
R1571 B.n363 B.n362 10.6151
R1572 B.n365 B.n152 10.6151
R1573 B.n369 B.n152 10.6151
R1574 B.n370 B.n369 10.6151
R1575 B.n371 B.n370 10.6151
R1576 B.n371 B.n150 10.6151
R1577 B.n375 B.n150 10.6151
R1578 B.n376 B.n375 10.6151
R1579 B.n377 B.n376 10.6151
R1580 B.n377 B.n148 10.6151
R1581 B.n381 B.n148 10.6151
R1582 B.n382 B.n381 10.6151
R1583 B.n383 B.n382 10.6151
R1584 B.n383 B.n146 10.6151
R1585 B.n387 B.n146 10.6151
R1586 B.n388 B.n387 10.6151
R1587 B.n389 B.n388 10.6151
R1588 B.n389 B.n144 10.6151
R1589 B.n393 B.n144 10.6151
R1590 B.n394 B.n393 10.6151
R1591 B.n395 B.n394 10.6151
R1592 B.n395 B.n142 10.6151
R1593 B.n399 B.n142 10.6151
R1594 B.n400 B.n399 10.6151
R1595 B.n401 B.n400 10.6151
R1596 B.n401 B.n140 10.6151
R1597 B.n405 B.n140 10.6151
R1598 B.n305 B.n176 10.6151
R1599 B.n305 B.n304 10.6151
R1600 B.n304 B.n303 10.6151
R1601 B.n303 B.n178 10.6151
R1602 B.n299 B.n178 10.6151
R1603 B.n299 B.n298 10.6151
R1604 B.n298 B.n297 10.6151
R1605 B.n297 B.n180 10.6151
R1606 B.n293 B.n180 10.6151
R1607 B.n293 B.n292 10.6151
R1608 B.n292 B.n291 10.6151
R1609 B.n291 B.n182 10.6151
R1610 B.n287 B.n182 10.6151
R1611 B.n287 B.n286 10.6151
R1612 B.n286 B.n285 10.6151
R1613 B.n285 B.n184 10.6151
R1614 B.n281 B.n184 10.6151
R1615 B.n281 B.n280 10.6151
R1616 B.n280 B.n279 10.6151
R1617 B.n279 B.n186 10.6151
R1618 B.n275 B.n186 10.6151
R1619 B.n275 B.n274 10.6151
R1620 B.n274 B.n273 10.6151
R1621 B.n273 B.n188 10.6151
R1622 B.n269 B.n188 10.6151
R1623 B.n269 B.n268 10.6151
R1624 B.n268 B.n267 10.6151
R1625 B.n267 B.n190 10.6151
R1626 B.n263 B.n190 10.6151
R1627 B.n263 B.n262 10.6151
R1628 B.n262 B.n261 10.6151
R1629 B.n261 B.n192 10.6151
R1630 B.n257 B.n192 10.6151
R1631 B.n257 B.n256 10.6151
R1632 B.n256 B.n255 10.6151
R1633 B.n255 B.n194 10.6151
R1634 B.n251 B.n194 10.6151
R1635 B.n251 B.n250 10.6151
R1636 B.n250 B.n249 10.6151
R1637 B.n249 B.n196 10.6151
R1638 B.n245 B.n196 10.6151
R1639 B.n245 B.n244 10.6151
R1640 B.n244 B.n243 10.6151
R1641 B.n243 B.n198 10.6151
R1642 B.n239 B.n198 10.6151
R1643 B.n239 B.n238 10.6151
R1644 B.n238 B.n237 10.6151
R1645 B.n237 B.n200 10.6151
R1646 B.n233 B.n200 10.6151
R1647 B.n233 B.n232 10.6151
R1648 B.n232 B.n231 10.6151
R1649 B.n231 B.n202 10.6151
R1650 B.n227 B.n202 10.6151
R1651 B.n227 B.n226 10.6151
R1652 B.n226 B.n225 10.6151
R1653 B.n225 B.n204 10.6151
R1654 B.n221 B.n204 10.6151
R1655 B.n221 B.n220 10.6151
R1656 B.n220 B.n219 10.6151
R1657 B.n219 B.n206 10.6151
R1658 B.n215 B.n206 10.6151
R1659 B.n215 B.n214 10.6151
R1660 B.n214 B.n213 10.6151
R1661 B.n213 B.n208 10.6151
R1662 B.n209 B.n208 10.6151
R1663 B.n209 B.n0 10.6151
R1664 B.n803 B.n1 10.6151
R1665 B.n803 B.n802 10.6151
R1666 B.n802 B.n801 10.6151
R1667 B.n801 B.n4 10.6151
R1668 B.n797 B.n4 10.6151
R1669 B.n797 B.n796 10.6151
R1670 B.n796 B.n795 10.6151
R1671 B.n795 B.n6 10.6151
R1672 B.n791 B.n6 10.6151
R1673 B.n791 B.n790 10.6151
R1674 B.n790 B.n789 10.6151
R1675 B.n789 B.n8 10.6151
R1676 B.n785 B.n8 10.6151
R1677 B.n785 B.n784 10.6151
R1678 B.n784 B.n783 10.6151
R1679 B.n783 B.n10 10.6151
R1680 B.n779 B.n10 10.6151
R1681 B.n779 B.n778 10.6151
R1682 B.n778 B.n777 10.6151
R1683 B.n777 B.n12 10.6151
R1684 B.n773 B.n12 10.6151
R1685 B.n773 B.n772 10.6151
R1686 B.n772 B.n771 10.6151
R1687 B.n771 B.n14 10.6151
R1688 B.n767 B.n14 10.6151
R1689 B.n767 B.n766 10.6151
R1690 B.n766 B.n765 10.6151
R1691 B.n765 B.n16 10.6151
R1692 B.n761 B.n16 10.6151
R1693 B.n761 B.n760 10.6151
R1694 B.n760 B.n759 10.6151
R1695 B.n759 B.n18 10.6151
R1696 B.n755 B.n18 10.6151
R1697 B.n755 B.n754 10.6151
R1698 B.n754 B.n753 10.6151
R1699 B.n753 B.n20 10.6151
R1700 B.n749 B.n20 10.6151
R1701 B.n749 B.n748 10.6151
R1702 B.n748 B.n747 10.6151
R1703 B.n747 B.n22 10.6151
R1704 B.n743 B.n22 10.6151
R1705 B.n743 B.n742 10.6151
R1706 B.n742 B.n741 10.6151
R1707 B.n741 B.n24 10.6151
R1708 B.n737 B.n24 10.6151
R1709 B.n737 B.n736 10.6151
R1710 B.n736 B.n735 10.6151
R1711 B.n735 B.n26 10.6151
R1712 B.n731 B.n26 10.6151
R1713 B.n731 B.n730 10.6151
R1714 B.n730 B.n729 10.6151
R1715 B.n729 B.n28 10.6151
R1716 B.n725 B.n28 10.6151
R1717 B.n725 B.n724 10.6151
R1718 B.n724 B.n723 10.6151
R1719 B.n723 B.n30 10.6151
R1720 B.n719 B.n30 10.6151
R1721 B.n719 B.n718 10.6151
R1722 B.n718 B.n717 10.6151
R1723 B.n717 B.n32 10.6151
R1724 B.n713 B.n32 10.6151
R1725 B.n713 B.n712 10.6151
R1726 B.n712 B.n711 10.6151
R1727 B.n711 B.n34 10.6151
R1728 B.n707 B.n34 10.6151
R1729 B.n707 B.n706 10.6151
R1730 B.n665 B.n664 9.36635
R1731 B.n647 B.n58 9.36635
R1732 B.n347 B.n162 9.36635
R1733 B.n365 B.n364 9.36635
R1734 B.n807 B.n0 2.81026
R1735 B.n807 B.n1 2.81026
R1736 B.n664 B.n663 1.24928
R1737 B.n650 B.n58 1.24928
R1738 B.n350 B.n162 1.24928
R1739 B.n364 B.n363 1.24928
R1740 VP.n27 VP.n24 161.3
R1741 VP.n29 VP.n28 161.3
R1742 VP.n30 VP.n23 161.3
R1743 VP.n32 VP.n31 161.3
R1744 VP.n33 VP.n22 161.3
R1745 VP.n35 VP.n34 161.3
R1746 VP.n36 VP.n21 161.3
R1747 VP.n39 VP.n38 161.3
R1748 VP.n40 VP.n20 161.3
R1749 VP.n42 VP.n41 161.3
R1750 VP.n43 VP.n19 161.3
R1751 VP.n45 VP.n44 161.3
R1752 VP.n46 VP.n18 161.3
R1753 VP.n48 VP.n47 161.3
R1754 VP.n50 VP.n17 161.3
R1755 VP.n52 VP.n51 161.3
R1756 VP.n53 VP.n16 161.3
R1757 VP.n55 VP.n54 161.3
R1758 VP.n56 VP.n15 161.3
R1759 VP.n58 VP.n57 161.3
R1760 VP.n103 VP.n102 161.3
R1761 VP.n101 VP.n1 161.3
R1762 VP.n100 VP.n99 161.3
R1763 VP.n98 VP.n2 161.3
R1764 VP.n97 VP.n96 161.3
R1765 VP.n95 VP.n3 161.3
R1766 VP.n93 VP.n92 161.3
R1767 VP.n91 VP.n4 161.3
R1768 VP.n90 VP.n89 161.3
R1769 VP.n88 VP.n5 161.3
R1770 VP.n87 VP.n86 161.3
R1771 VP.n85 VP.n6 161.3
R1772 VP.n84 VP.n83 161.3
R1773 VP.n81 VP.n7 161.3
R1774 VP.n80 VP.n79 161.3
R1775 VP.n78 VP.n8 161.3
R1776 VP.n77 VP.n76 161.3
R1777 VP.n75 VP.n9 161.3
R1778 VP.n74 VP.n73 161.3
R1779 VP.n72 VP.n10 161.3
R1780 VP.n71 VP.n70 161.3
R1781 VP.n68 VP.n11 161.3
R1782 VP.n67 VP.n66 161.3
R1783 VP.n65 VP.n12 161.3
R1784 VP.n64 VP.n63 161.3
R1785 VP.n62 VP.n13 161.3
R1786 VP.n26 VP.t3 89.3009
R1787 VP.n61 VP.n60 70.0045
R1788 VP.n104 VP.n0 70.0045
R1789 VP.n59 VP.n14 70.0045
R1790 VP.n26 VP.n25 69.7461
R1791 VP.n61 VP.t1 57.5995
R1792 VP.n69 VP.t6 57.5995
R1793 VP.n82 VP.t4 57.5995
R1794 VP.n94 VP.t7 57.5995
R1795 VP.n0 VP.t0 57.5995
R1796 VP.n14 VP.t5 57.5995
R1797 VP.n49 VP.t8 57.5995
R1798 VP.n37 VP.t9 57.5995
R1799 VP.n25 VP.t2 57.5995
R1800 VP.n67 VP.n12 56.5193
R1801 VP.n100 VP.n2 56.5193
R1802 VP.n55 VP.n16 56.5193
R1803 VP.n60 VP.n59 51.7531
R1804 VP.n76 VP.n8 48.7492
R1805 VP.n88 VP.n87 48.7492
R1806 VP.n43 VP.n42 48.7492
R1807 VP.n31 VP.n22 48.7492
R1808 VP.n76 VP.n75 32.2376
R1809 VP.n89 VP.n88 32.2376
R1810 VP.n44 VP.n43 32.2376
R1811 VP.n31 VP.n30 32.2376
R1812 VP.n63 VP.n62 24.4675
R1813 VP.n63 VP.n12 24.4675
R1814 VP.n68 VP.n67 24.4675
R1815 VP.n70 VP.n68 24.4675
R1816 VP.n74 VP.n10 24.4675
R1817 VP.n75 VP.n74 24.4675
R1818 VP.n80 VP.n8 24.4675
R1819 VP.n81 VP.n80 24.4675
R1820 VP.n83 VP.n6 24.4675
R1821 VP.n87 VP.n6 24.4675
R1822 VP.n89 VP.n4 24.4675
R1823 VP.n93 VP.n4 24.4675
R1824 VP.n96 VP.n95 24.4675
R1825 VP.n96 VP.n2 24.4675
R1826 VP.n101 VP.n100 24.4675
R1827 VP.n102 VP.n101 24.4675
R1828 VP.n56 VP.n55 24.4675
R1829 VP.n57 VP.n56 24.4675
R1830 VP.n44 VP.n18 24.4675
R1831 VP.n48 VP.n18 24.4675
R1832 VP.n51 VP.n50 24.4675
R1833 VP.n51 VP.n16 24.4675
R1834 VP.n35 VP.n22 24.4675
R1835 VP.n36 VP.n35 24.4675
R1836 VP.n38 VP.n20 24.4675
R1837 VP.n42 VP.n20 24.4675
R1838 VP.n29 VP.n24 24.4675
R1839 VP.n30 VP.n29 24.4675
R1840 VP.n70 VP.n69 20.5528
R1841 VP.n95 VP.n94 20.5528
R1842 VP.n50 VP.n49 20.5528
R1843 VP.n62 VP.n61 20.0634
R1844 VP.n102 VP.n0 20.0634
R1845 VP.n57 VP.n14 20.0634
R1846 VP.n82 VP.n81 12.234
R1847 VP.n83 VP.n82 12.234
R1848 VP.n37 VP.n36 12.234
R1849 VP.n38 VP.n37 12.234
R1850 VP.n27 VP.n26 5.54913
R1851 VP.n69 VP.n10 3.91522
R1852 VP.n94 VP.n93 3.91522
R1853 VP.n49 VP.n48 3.91522
R1854 VP.n25 VP.n24 3.91522
R1855 VP.n59 VP.n58 0.354971
R1856 VP.n60 VP.n13 0.354971
R1857 VP.n104 VP.n103 0.354971
R1858 VP VP.n104 0.26696
R1859 VP.n28 VP.n27 0.189894
R1860 VP.n28 VP.n23 0.189894
R1861 VP.n32 VP.n23 0.189894
R1862 VP.n33 VP.n32 0.189894
R1863 VP.n34 VP.n33 0.189894
R1864 VP.n34 VP.n21 0.189894
R1865 VP.n39 VP.n21 0.189894
R1866 VP.n40 VP.n39 0.189894
R1867 VP.n41 VP.n40 0.189894
R1868 VP.n41 VP.n19 0.189894
R1869 VP.n45 VP.n19 0.189894
R1870 VP.n46 VP.n45 0.189894
R1871 VP.n47 VP.n46 0.189894
R1872 VP.n47 VP.n17 0.189894
R1873 VP.n52 VP.n17 0.189894
R1874 VP.n53 VP.n52 0.189894
R1875 VP.n54 VP.n53 0.189894
R1876 VP.n54 VP.n15 0.189894
R1877 VP.n58 VP.n15 0.189894
R1878 VP.n64 VP.n13 0.189894
R1879 VP.n65 VP.n64 0.189894
R1880 VP.n66 VP.n65 0.189894
R1881 VP.n66 VP.n11 0.189894
R1882 VP.n71 VP.n11 0.189894
R1883 VP.n72 VP.n71 0.189894
R1884 VP.n73 VP.n72 0.189894
R1885 VP.n73 VP.n9 0.189894
R1886 VP.n77 VP.n9 0.189894
R1887 VP.n78 VP.n77 0.189894
R1888 VP.n79 VP.n78 0.189894
R1889 VP.n79 VP.n7 0.189894
R1890 VP.n84 VP.n7 0.189894
R1891 VP.n85 VP.n84 0.189894
R1892 VP.n86 VP.n85 0.189894
R1893 VP.n86 VP.n5 0.189894
R1894 VP.n90 VP.n5 0.189894
R1895 VP.n91 VP.n90 0.189894
R1896 VP.n92 VP.n91 0.189894
R1897 VP.n92 VP.n3 0.189894
R1898 VP.n97 VP.n3 0.189894
R1899 VP.n98 VP.n97 0.189894
R1900 VP.n99 VP.n98 0.189894
R1901 VP.n99 VP.n1 0.189894
R1902 VP.n103 VP.n1 0.189894
R1903 VDD1.n31 VDD1.n30 585
R1904 VDD1.n29 VDD1.n28 585
R1905 VDD1.n4 VDD1.n3 585
R1906 VDD1.n23 VDD1.n22 585
R1907 VDD1.n21 VDD1.n20 585
R1908 VDD1.n8 VDD1.n7 585
R1909 VDD1.n15 VDD1.n14 585
R1910 VDD1.n13 VDD1.n12 585
R1911 VDD1.n50 VDD1.n49 585
R1912 VDD1.n52 VDD1.n51 585
R1913 VDD1.n45 VDD1.n44 585
R1914 VDD1.n58 VDD1.n57 585
R1915 VDD1.n60 VDD1.n59 585
R1916 VDD1.n41 VDD1.n40 585
R1917 VDD1.n66 VDD1.n65 585
R1918 VDD1.n68 VDD1.n67 585
R1919 VDD1.n30 VDD1.n0 498.474
R1920 VDD1.n67 VDD1.n37 498.474
R1921 VDD1.n11 VDD1.t6 329.053
R1922 VDD1.n48 VDD1.t8 329.053
R1923 VDD1.n30 VDD1.n29 171.744
R1924 VDD1.n29 VDD1.n3 171.744
R1925 VDD1.n22 VDD1.n3 171.744
R1926 VDD1.n22 VDD1.n21 171.744
R1927 VDD1.n21 VDD1.n7 171.744
R1928 VDD1.n14 VDD1.n7 171.744
R1929 VDD1.n14 VDD1.n13 171.744
R1930 VDD1.n51 VDD1.n50 171.744
R1931 VDD1.n51 VDD1.n44 171.744
R1932 VDD1.n58 VDD1.n44 171.744
R1933 VDD1.n59 VDD1.n58 171.744
R1934 VDD1.n59 VDD1.n40 171.744
R1935 VDD1.n66 VDD1.n40 171.744
R1936 VDD1.n67 VDD1.n66 171.744
R1937 VDD1.n75 VDD1.n74 88.6818
R1938 VDD1.n36 VDD1.n35 86.5843
R1939 VDD1.n73 VDD1.n72 86.5842
R1940 VDD1.n77 VDD1.n76 86.5842
R1941 VDD1.n13 VDD1.t6 85.8723
R1942 VDD1.n50 VDD1.t8 85.8723
R1943 VDD1.n36 VDD1.n34 53.4803
R1944 VDD1.n73 VDD1.n71 53.4803
R1945 VDD1.n77 VDD1.n75 45.5505
R1946 VDD1.n32 VDD1.n31 12.8005
R1947 VDD1.n69 VDD1.n68 12.8005
R1948 VDD1.n28 VDD1.n2 12.0247
R1949 VDD1.n65 VDD1.n39 12.0247
R1950 VDD1.n27 VDD1.n4 11.249
R1951 VDD1.n64 VDD1.n41 11.249
R1952 VDD1.n12 VDD1.n11 10.7237
R1953 VDD1.n49 VDD1.n48 10.7237
R1954 VDD1.n24 VDD1.n23 10.4732
R1955 VDD1.n61 VDD1.n60 10.4732
R1956 VDD1.n20 VDD1.n6 9.69747
R1957 VDD1.n57 VDD1.n43 9.69747
R1958 VDD1.n34 VDD1.n33 9.45567
R1959 VDD1.n71 VDD1.n70 9.45567
R1960 VDD1.n10 VDD1.n9 9.3005
R1961 VDD1.n17 VDD1.n16 9.3005
R1962 VDD1.n19 VDD1.n18 9.3005
R1963 VDD1.n6 VDD1.n5 9.3005
R1964 VDD1.n25 VDD1.n24 9.3005
R1965 VDD1.n27 VDD1.n26 9.3005
R1966 VDD1.n2 VDD1.n1 9.3005
R1967 VDD1.n33 VDD1.n32 9.3005
R1968 VDD1.n47 VDD1.n46 9.3005
R1969 VDD1.n54 VDD1.n53 9.3005
R1970 VDD1.n56 VDD1.n55 9.3005
R1971 VDD1.n43 VDD1.n42 9.3005
R1972 VDD1.n62 VDD1.n61 9.3005
R1973 VDD1.n64 VDD1.n63 9.3005
R1974 VDD1.n39 VDD1.n38 9.3005
R1975 VDD1.n70 VDD1.n69 9.3005
R1976 VDD1.n19 VDD1.n8 8.92171
R1977 VDD1.n56 VDD1.n45 8.92171
R1978 VDD1.n16 VDD1.n15 8.14595
R1979 VDD1.n53 VDD1.n52 8.14595
R1980 VDD1.n34 VDD1.n0 7.75445
R1981 VDD1.n71 VDD1.n37 7.75445
R1982 VDD1.n12 VDD1.n10 7.3702
R1983 VDD1.n49 VDD1.n47 7.3702
R1984 VDD1.n32 VDD1.n0 6.08283
R1985 VDD1.n69 VDD1.n37 6.08283
R1986 VDD1.n15 VDD1.n10 5.81868
R1987 VDD1.n52 VDD1.n47 5.81868
R1988 VDD1.n16 VDD1.n8 5.04292
R1989 VDD1.n53 VDD1.n45 5.04292
R1990 VDD1.n76 VDD1.t1 4.53397
R1991 VDD1.n76 VDD1.t4 4.53397
R1992 VDD1.n35 VDD1.t7 4.53397
R1993 VDD1.n35 VDD1.t0 4.53397
R1994 VDD1.n74 VDD1.t2 4.53397
R1995 VDD1.n74 VDD1.t9 4.53397
R1996 VDD1.n72 VDD1.t3 4.53397
R1997 VDD1.n72 VDD1.t5 4.53397
R1998 VDD1.n20 VDD1.n19 4.26717
R1999 VDD1.n57 VDD1.n56 4.26717
R2000 VDD1.n23 VDD1.n6 3.49141
R2001 VDD1.n60 VDD1.n43 3.49141
R2002 VDD1.n24 VDD1.n4 2.71565
R2003 VDD1.n61 VDD1.n41 2.71565
R2004 VDD1.n11 VDD1.n9 2.41305
R2005 VDD1.n48 VDD1.n46 2.41305
R2006 VDD1 VDD1.n77 2.09533
R2007 VDD1.n28 VDD1.n27 1.93989
R2008 VDD1.n65 VDD1.n64 1.93989
R2009 VDD1.n31 VDD1.n2 1.16414
R2010 VDD1.n68 VDD1.n39 1.16414
R2011 VDD1 VDD1.n36 0.776362
R2012 VDD1.n75 VDD1.n73 0.662826
R2013 VDD1.n33 VDD1.n1 0.155672
R2014 VDD1.n26 VDD1.n1 0.155672
R2015 VDD1.n26 VDD1.n25 0.155672
R2016 VDD1.n25 VDD1.n5 0.155672
R2017 VDD1.n18 VDD1.n5 0.155672
R2018 VDD1.n18 VDD1.n17 0.155672
R2019 VDD1.n17 VDD1.n9 0.155672
R2020 VDD1.n54 VDD1.n46 0.155672
R2021 VDD1.n55 VDD1.n54 0.155672
R2022 VDD1.n55 VDD1.n42 0.155672
R2023 VDD1.n62 VDD1.n42 0.155672
R2024 VDD1.n63 VDD1.n62 0.155672
R2025 VDD1.n63 VDD1.n38 0.155672
R2026 VDD1.n70 VDD1.n38 0.155672
C0 VDD2 VTAIL 8.50074f
C1 VP B 2.41965f
C2 VDD1 w_n4966_n2402# 2.6082f
C3 VN VDD1 0.15429f
C4 w_n4966_n2402# VP 11.3043f
C5 VN VP 8.09594f
C6 VDD2 VDD1 2.43452f
C7 w_n4966_n2402# B 9.867769f
C8 VN B 1.32816f
C9 VDD2 VP 0.634279f
C10 VDD1 VTAIL 8.44576f
C11 VN w_n4966_n2402# 10.6565f
C12 VDD2 B 2.3852f
C13 VTAIL VP 8.025221f
C14 VDD2 w_n4966_n2402# 2.77254f
C15 VDD2 VN 6.75714f
C16 VTAIL B 2.7803f
C17 VDD1 VP 7.234009f
C18 w_n4966_n2402# VTAIL 2.60331f
C19 VN VTAIL 8.01102f
C20 VDD1 B 2.25171f
C21 VDD2 VSUBS 2.245192f
C22 VDD1 VSUBS 2.011895f
C23 VTAIL VSUBS 0.752207f
C24 VN VSUBS 8.07706f
C25 VP VSUBS 4.339729f
C26 B VSUBS 5.457196f
C27 w_n4966_n2402# VSUBS 0.148324p
C28 VDD1.n0 VSUBS 0.034801f
C29 VDD1.n1 VSUBS 0.033297f
C30 VDD1.n2 VSUBS 0.017892f
C31 VDD1.n3 VSUBS 0.042291f
C32 VDD1.n4 VSUBS 0.018945f
C33 VDD1.n5 VSUBS 0.033297f
C34 VDD1.n6 VSUBS 0.017892f
C35 VDD1.n7 VSUBS 0.042291f
C36 VDD1.n8 VSUBS 0.018945f
C37 VDD1.n9 VSUBS 0.930921f
C38 VDD1.n10 VSUBS 0.017892f
C39 VDD1.t6 VSUBS 0.090801f
C40 VDD1.n11 VSUBS 0.189688f
C41 VDD1.n12 VSUBS 0.031812f
C42 VDD1.n13 VSUBS 0.031718f
C43 VDD1.n14 VSUBS 0.042291f
C44 VDD1.n15 VSUBS 0.018945f
C45 VDD1.n16 VSUBS 0.017892f
C46 VDD1.n17 VSUBS 0.033297f
C47 VDD1.n18 VSUBS 0.033297f
C48 VDD1.n19 VSUBS 0.017892f
C49 VDD1.n20 VSUBS 0.018945f
C50 VDD1.n21 VSUBS 0.042291f
C51 VDD1.n22 VSUBS 0.042291f
C52 VDD1.n23 VSUBS 0.018945f
C53 VDD1.n24 VSUBS 0.017892f
C54 VDD1.n25 VSUBS 0.033297f
C55 VDD1.n26 VSUBS 0.033297f
C56 VDD1.n27 VSUBS 0.017892f
C57 VDD1.n28 VSUBS 0.018945f
C58 VDD1.n29 VSUBS 0.042291f
C59 VDD1.n30 VSUBS 0.103099f
C60 VDD1.n31 VSUBS 0.018945f
C61 VDD1.n32 VSUBS 0.035136f
C62 VDD1.n33 VSUBS 0.081058f
C63 VDD1.n34 VSUBS 0.120987f
C64 VDD1.t7 VSUBS 0.188658f
C65 VDD1.t0 VSUBS 0.188658f
C66 VDD1.n35 VSUBS 1.33181f
C67 VDD1.n36 VSUBS 1.29361f
C68 VDD1.n37 VSUBS 0.034801f
C69 VDD1.n38 VSUBS 0.033297f
C70 VDD1.n39 VSUBS 0.017892f
C71 VDD1.n40 VSUBS 0.042291f
C72 VDD1.n41 VSUBS 0.018945f
C73 VDD1.n42 VSUBS 0.033297f
C74 VDD1.n43 VSUBS 0.017892f
C75 VDD1.n44 VSUBS 0.042291f
C76 VDD1.n45 VSUBS 0.018945f
C77 VDD1.n46 VSUBS 0.930921f
C78 VDD1.n47 VSUBS 0.017892f
C79 VDD1.t8 VSUBS 0.090801f
C80 VDD1.n48 VSUBS 0.189688f
C81 VDD1.n49 VSUBS 0.031812f
C82 VDD1.n50 VSUBS 0.031718f
C83 VDD1.n51 VSUBS 0.042291f
C84 VDD1.n52 VSUBS 0.018945f
C85 VDD1.n53 VSUBS 0.017892f
C86 VDD1.n54 VSUBS 0.033297f
C87 VDD1.n55 VSUBS 0.033297f
C88 VDD1.n56 VSUBS 0.017892f
C89 VDD1.n57 VSUBS 0.018945f
C90 VDD1.n58 VSUBS 0.042291f
C91 VDD1.n59 VSUBS 0.042291f
C92 VDD1.n60 VSUBS 0.018945f
C93 VDD1.n61 VSUBS 0.017892f
C94 VDD1.n62 VSUBS 0.033297f
C95 VDD1.n63 VSUBS 0.033297f
C96 VDD1.n64 VSUBS 0.017892f
C97 VDD1.n65 VSUBS 0.018945f
C98 VDD1.n66 VSUBS 0.042291f
C99 VDD1.n67 VSUBS 0.103099f
C100 VDD1.n68 VSUBS 0.018945f
C101 VDD1.n69 VSUBS 0.035136f
C102 VDD1.n70 VSUBS 0.081058f
C103 VDD1.n71 VSUBS 0.120987f
C104 VDD1.t3 VSUBS 0.188658f
C105 VDD1.t5 VSUBS 0.188658f
C106 VDD1.n72 VSUBS 1.33181f
C107 VDD1.n73 VSUBS 1.2826f
C108 VDD1.t2 VSUBS 0.188658f
C109 VDD1.t9 VSUBS 0.188658f
C110 VDD1.n74 VSUBS 1.3577f
C111 VDD1.n75 VSUBS 4.20309f
C112 VDD1.t1 VSUBS 0.188658f
C113 VDD1.t4 VSUBS 0.188658f
C114 VDD1.n76 VSUBS 1.33181f
C115 VDD1.n77 VSUBS 4.22752f
C116 VP.t0 VSUBS 1.99307f
C117 VP.n0 VSUBS 0.865793f
C118 VP.n1 VSUBS 0.034675f
C119 VP.n2 VSUBS 0.05014f
C120 VP.n3 VSUBS 0.034675f
C121 VP.t7 VSUBS 1.99307f
C122 VP.n4 VSUBS 0.064626f
C123 VP.n5 VSUBS 0.034675f
C124 VP.n6 VSUBS 0.064626f
C125 VP.n7 VSUBS 0.034675f
C126 VP.t4 VSUBS 1.99307f
C127 VP.n8 VSUBS 0.064626f
C128 VP.n9 VSUBS 0.034675f
C129 VP.n10 VSUBS 0.037825f
C130 VP.n11 VSUBS 0.034675f
C131 VP.n12 VSUBS 0.051106f
C132 VP.n13 VSUBS 0.055965f
C133 VP.t1 VSUBS 1.99307f
C134 VP.t5 VSUBS 1.99307f
C135 VP.n14 VSUBS 0.865793f
C136 VP.n15 VSUBS 0.034675f
C137 VP.n16 VSUBS 0.05014f
C138 VP.n17 VSUBS 0.034675f
C139 VP.t8 VSUBS 1.99307f
C140 VP.n18 VSUBS 0.064626f
C141 VP.n19 VSUBS 0.034675f
C142 VP.n20 VSUBS 0.064626f
C143 VP.n21 VSUBS 0.034675f
C144 VP.t9 VSUBS 1.99307f
C145 VP.n22 VSUBS 0.064626f
C146 VP.n23 VSUBS 0.034675f
C147 VP.n24 VSUBS 0.037825f
C148 VP.t3 VSUBS 2.33408f
C149 VP.t2 VSUBS 1.99307f
C150 VP.n25 VSUBS 0.828661f
C151 VP.n26 VSUBS 0.803267f
C152 VP.n27 VSUBS 0.375004f
C153 VP.n28 VSUBS 0.034675f
C154 VP.n29 VSUBS 0.064626f
C155 VP.n30 VSUBS 0.069855f
C156 VP.n31 VSUBS 0.03139f
C157 VP.n32 VSUBS 0.034675f
C158 VP.n33 VSUBS 0.034675f
C159 VP.n34 VSUBS 0.034675f
C160 VP.n35 VSUBS 0.064626f
C161 VP.n36 VSUBS 0.048673f
C162 VP.n37 VSUBS 0.728656f
C163 VP.n38 VSUBS 0.048673f
C164 VP.n39 VSUBS 0.034675f
C165 VP.n40 VSUBS 0.034675f
C166 VP.n41 VSUBS 0.034675f
C167 VP.n42 VSUBS 0.064626f
C168 VP.n43 VSUBS 0.03139f
C169 VP.n44 VSUBS 0.069855f
C170 VP.n45 VSUBS 0.034675f
C171 VP.n46 VSUBS 0.034675f
C172 VP.n47 VSUBS 0.034675f
C173 VP.n48 VSUBS 0.037825f
C174 VP.n49 VSUBS 0.728656f
C175 VP.n50 VSUBS 0.059521f
C176 VP.n51 VSUBS 0.064626f
C177 VP.n52 VSUBS 0.034675f
C178 VP.n53 VSUBS 0.034675f
C179 VP.n54 VSUBS 0.034675f
C180 VP.n55 VSUBS 0.051106f
C181 VP.n56 VSUBS 0.064626f
C182 VP.n57 VSUBS 0.058883f
C183 VP.n58 VSUBS 0.055965f
C184 VP.n59 VSUBS 2.05929f
C185 VP.n60 VSUBS 2.08338f
C186 VP.n61 VSUBS 0.865793f
C187 VP.n62 VSUBS 0.058883f
C188 VP.n63 VSUBS 0.064626f
C189 VP.n64 VSUBS 0.034675f
C190 VP.n65 VSUBS 0.034675f
C191 VP.n66 VSUBS 0.034675f
C192 VP.n67 VSUBS 0.05014f
C193 VP.n68 VSUBS 0.064626f
C194 VP.t6 VSUBS 1.99307f
C195 VP.n69 VSUBS 0.728656f
C196 VP.n70 VSUBS 0.059521f
C197 VP.n71 VSUBS 0.034675f
C198 VP.n72 VSUBS 0.034675f
C199 VP.n73 VSUBS 0.034675f
C200 VP.n74 VSUBS 0.064626f
C201 VP.n75 VSUBS 0.069855f
C202 VP.n76 VSUBS 0.03139f
C203 VP.n77 VSUBS 0.034675f
C204 VP.n78 VSUBS 0.034675f
C205 VP.n79 VSUBS 0.034675f
C206 VP.n80 VSUBS 0.064626f
C207 VP.n81 VSUBS 0.048673f
C208 VP.n82 VSUBS 0.728656f
C209 VP.n83 VSUBS 0.048673f
C210 VP.n84 VSUBS 0.034675f
C211 VP.n85 VSUBS 0.034675f
C212 VP.n86 VSUBS 0.034675f
C213 VP.n87 VSUBS 0.064626f
C214 VP.n88 VSUBS 0.03139f
C215 VP.n89 VSUBS 0.069855f
C216 VP.n90 VSUBS 0.034675f
C217 VP.n91 VSUBS 0.034675f
C218 VP.n92 VSUBS 0.034675f
C219 VP.n93 VSUBS 0.037825f
C220 VP.n94 VSUBS 0.728656f
C221 VP.n95 VSUBS 0.059521f
C222 VP.n96 VSUBS 0.064626f
C223 VP.n97 VSUBS 0.034675f
C224 VP.n98 VSUBS 0.034675f
C225 VP.n99 VSUBS 0.034675f
C226 VP.n100 VSUBS 0.051106f
C227 VP.n101 VSUBS 0.064626f
C228 VP.n102 VSUBS 0.058883f
C229 VP.n103 VSUBS 0.055965f
C230 VP.n104 VSUBS 0.072065f
C231 B.n0 VSUBS 0.007f
C232 B.n1 VSUBS 0.007f
C233 B.n2 VSUBS 0.01107f
C234 B.n3 VSUBS 0.01107f
C235 B.n4 VSUBS 0.01107f
C236 B.n5 VSUBS 0.01107f
C237 B.n6 VSUBS 0.01107f
C238 B.n7 VSUBS 0.01107f
C239 B.n8 VSUBS 0.01107f
C240 B.n9 VSUBS 0.01107f
C241 B.n10 VSUBS 0.01107f
C242 B.n11 VSUBS 0.01107f
C243 B.n12 VSUBS 0.01107f
C244 B.n13 VSUBS 0.01107f
C245 B.n14 VSUBS 0.01107f
C246 B.n15 VSUBS 0.01107f
C247 B.n16 VSUBS 0.01107f
C248 B.n17 VSUBS 0.01107f
C249 B.n18 VSUBS 0.01107f
C250 B.n19 VSUBS 0.01107f
C251 B.n20 VSUBS 0.01107f
C252 B.n21 VSUBS 0.01107f
C253 B.n22 VSUBS 0.01107f
C254 B.n23 VSUBS 0.01107f
C255 B.n24 VSUBS 0.01107f
C256 B.n25 VSUBS 0.01107f
C257 B.n26 VSUBS 0.01107f
C258 B.n27 VSUBS 0.01107f
C259 B.n28 VSUBS 0.01107f
C260 B.n29 VSUBS 0.01107f
C261 B.n30 VSUBS 0.01107f
C262 B.n31 VSUBS 0.01107f
C263 B.n32 VSUBS 0.01107f
C264 B.n33 VSUBS 0.01107f
C265 B.n34 VSUBS 0.01107f
C266 B.n35 VSUBS 0.025943f
C267 B.n36 VSUBS 0.01107f
C268 B.n37 VSUBS 0.01107f
C269 B.n38 VSUBS 0.01107f
C270 B.n39 VSUBS 0.01107f
C271 B.n40 VSUBS 0.01107f
C272 B.n41 VSUBS 0.01107f
C273 B.n42 VSUBS 0.01107f
C274 B.n43 VSUBS 0.01107f
C275 B.n44 VSUBS 0.01107f
C276 B.n45 VSUBS 0.01107f
C277 B.n46 VSUBS 0.01107f
C278 B.n47 VSUBS 0.01107f
C279 B.n48 VSUBS 0.01107f
C280 B.n49 VSUBS 0.01107f
C281 B.t8 VSUBS 0.174573f
C282 B.t7 VSUBS 0.22359f
C283 B.t6 VSUBS 1.60688f
C284 B.n50 VSUBS 0.372573f
C285 B.n51 VSUBS 0.283856f
C286 B.n52 VSUBS 0.01107f
C287 B.n53 VSUBS 0.01107f
C288 B.n54 VSUBS 0.01107f
C289 B.n55 VSUBS 0.01107f
C290 B.t11 VSUBS 0.174577f
C291 B.t10 VSUBS 0.223593f
C292 B.t9 VSUBS 1.60688f
C293 B.n56 VSUBS 0.37257f
C294 B.n57 VSUBS 0.283852f
C295 B.n58 VSUBS 0.025648f
C296 B.n59 VSUBS 0.01107f
C297 B.n60 VSUBS 0.01107f
C298 B.n61 VSUBS 0.01107f
C299 B.n62 VSUBS 0.01107f
C300 B.n63 VSUBS 0.01107f
C301 B.n64 VSUBS 0.01107f
C302 B.n65 VSUBS 0.01107f
C303 B.n66 VSUBS 0.01107f
C304 B.n67 VSUBS 0.01107f
C305 B.n68 VSUBS 0.01107f
C306 B.n69 VSUBS 0.01107f
C307 B.n70 VSUBS 0.01107f
C308 B.n71 VSUBS 0.01107f
C309 B.n72 VSUBS 0.027228f
C310 B.n73 VSUBS 0.01107f
C311 B.n74 VSUBS 0.01107f
C312 B.n75 VSUBS 0.01107f
C313 B.n76 VSUBS 0.01107f
C314 B.n77 VSUBS 0.01107f
C315 B.n78 VSUBS 0.01107f
C316 B.n79 VSUBS 0.01107f
C317 B.n80 VSUBS 0.01107f
C318 B.n81 VSUBS 0.01107f
C319 B.n82 VSUBS 0.01107f
C320 B.n83 VSUBS 0.01107f
C321 B.n84 VSUBS 0.01107f
C322 B.n85 VSUBS 0.01107f
C323 B.n86 VSUBS 0.01107f
C324 B.n87 VSUBS 0.01107f
C325 B.n88 VSUBS 0.01107f
C326 B.n89 VSUBS 0.01107f
C327 B.n90 VSUBS 0.01107f
C328 B.n91 VSUBS 0.01107f
C329 B.n92 VSUBS 0.01107f
C330 B.n93 VSUBS 0.01107f
C331 B.n94 VSUBS 0.01107f
C332 B.n95 VSUBS 0.01107f
C333 B.n96 VSUBS 0.01107f
C334 B.n97 VSUBS 0.01107f
C335 B.n98 VSUBS 0.01107f
C336 B.n99 VSUBS 0.01107f
C337 B.n100 VSUBS 0.01107f
C338 B.n101 VSUBS 0.01107f
C339 B.n102 VSUBS 0.01107f
C340 B.n103 VSUBS 0.01107f
C341 B.n104 VSUBS 0.01107f
C342 B.n105 VSUBS 0.01107f
C343 B.n106 VSUBS 0.01107f
C344 B.n107 VSUBS 0.01107f
C345 B.n108 VSUBS 0.01107f
C346 B.n109 VSUBS 0.01107f
C347 B.n110 VSUBS 0.01107f
C348 B.n111 VSUBS 0.01107f
C349 B.n112 VSUBS 0.01107f
C350 B.n113 VSUBS 0.01107f
C351 B.n114 VSUBS 0.01107f
C352 B.n115 VSUBS 0.01107f
C353 B.n116 VSUBS 0.01107f
C354 B.n117 VSUBS 0.01107f
C355 B.n118 VSUBS 0.01107f
C356 B.n119 VSUBS 0.01107f
C357 B.n120 VSUBS 0.01107f
C358 B.n121 VSUBS 0.01107f
C359 B.n122 VSUBS 0.01107f
C360 B.n123 VSUBS 0.01107f
C361 B.n124 VSUBS 0.01107f
C362 B.n125 VSUBS 0.01107f
C363 B.n126 VSUBS 0.01107f
C364 B.n127 VSUBS 0.01107f
C365 B.n128 VSUBS 0.01107f
C366 B.n129 VSUBS 0.01107f
C367 B.n130 VSUBS 0.01107f
C368 B.n131 VSUBS 0.01107f
C369 B.n132 VSUBS 0.01107f
C370 B.n133 VSUBS 0.01107f
C371 B.n134 VSUBS 0.01107f
C372 B.n135 VSUBS 0.01107f
C373 B.n136 VSUBS 0.01107f
C374 B.n137 VSUBS 0.01107f
C375 B.n138 VSUBS 0.01107f
C376 B.n139 VSUBS 0.025943f
C377 B.n140 VSUBS 0.01107f
C378 B.n141 VSUBS 0.01107f
C379 B.n142 VSUBS 0.01107f
C380 B.n143 VSUBS 0.01107f
C381 B.n144 VSUBS 0.01107f
C382 B.n145 VSUBS 0.01107f
C383 B.n146 VSUBS 0.01107f
C384 B.n147 VSUBS 0.01107f
C385 B.n148 VSUBS 0.01107f
C386 B.n149 VSUBS 0.01107f
C387 B.n150 VSUBS 0.01107f
C388 B.n151 VSUBS 0.01107f
C389 B.n152 VSUBS 0.01107f
C390 B.n153 VSUBS 0.01107f
C391 B.t1 VSUBS 0.174577f
C392 B.t2 VSUBS 0.223593f
C393 B.t0 VSUBS 1.60688f
C394 B.n154 VSUBS 0.37257f
C395 B.n155 VSUBS 0.283852f
C396 B.n156 VSUBS 0.01107f
C397 B.n157 VSUBS 0.01107f
C398 B.n158 VSUBS 0.01107f
C399 B.n159 VSUBS 0.01107f
C400 B.t4 VSUBS 0.174573f
C401 B.t5 VSUBS 0.22359f
C402 B.t3 VSUBS 1.60688f
C403 B.n160 VSUBS 0.372573f
C404 B.n161 VSUBS 0.283856f
C405 B.n162 VSUBS 0.025648f
C406 B.n163 VSUBS 0.01107f
C407 B.n164 VSUBS 0.01107f
C408 B.n165 VSUBS 0.01107f
C409 B.n166 VSUBS 0.01107f
C410 B.n167 VSUBS 0.01107f
C411 B.n168 VSUBS 0.01107f
C412 B.n169 VSUBS 0.01107f
C413 B.n170 VSUBS 0.01107f
C414 B.n171 VSUBS 0.01107f
C415 B.n172 VSUBS 0.01107f
C416 B.n173 VSUBS 0.01107f
C417 B.n174 VSUBS 0.01107f
C418 B.n175 VSUBS 0.01107f
C419 B.n176 VSUBS 0.025943f
C420 B.n177 VSUBS 0.01107f
C421 B.n178 VSUBS 0.01107f
C422 B.n179 VSUBS 0.01107f
C423 B.n180 VSUBS 0.01107f
C424 B.n181 VSUBS 0.01107f
C425 B.n182 VSUBS 0.01107f
C426 B.n183 VSUBS 0.01107f
C427 B.n184 VSUBS 0.01107f
C428 B.n185 VSUBS 0.01107f
C429 B.n186 VSUBS 0.01107f
C430 B.n187 VSUBS 0.01107f
C431 B.n188 VSUBS 0.01107f
C432 B.n189 VSUBS 0.01107f
C433 B.n190 VSUBS 0.01107f
C434 B.n191 VSUBS 0.01107f
C435 B.n192 VSUBS 0.01107f
C436 B.n193 VSUBS 0.01107f
C437 B.n194 VSUBS 0.01107f
C438 B.n195 VSUBS 0.01107f
C439 B.n196 VSUBS 0.01107f
C440 B.n197 VSUBS 0.01107f
C441 B.n198 VSUBS 0.01107f
C442 B.n199 VSUBS 0.01107f
C443 B.n200 VSUBS 0.01107f
C444 B.n201 VSUBS 0.01107f
C445 B.n202 VSUBS 0.01107f
C446 B.n203 VSUBS 0.01107f
C447 B.n204 VSUBS 0.01107f
C448 B.n205 VSUBS 0.01107f
C449 B.n206 VSUBS 0.01107f
C450 B.n207 VSUBS 0.01107f
C451 B.n208 VSUBS 0.01107f
C452 B.n209 VSUBS 0.01107f
C453 B.n210 VSUBS 0.01107f
C454 B.n211 VSUBS 0.01107f
C455 B.n212 VSUBS 0.01107f
C456 B.n213 VSUBS 0.01107f
C457 B.n214 VSUBS 0.01107f
C458 B.n215 VSUBS 0.01107f
C459 B.n216 VSUBS 0.01107f
C460 B.n217 VSUBS 0.01107f
C461 B.n218 VSUBS 0.01107f
C462 B.n219 VSUBS 0.01107f
C463 B.n220 VSUBS 0.01107f
C464 B.n221 VSUBS 0.01107f
C465 B.n222 VSUBS 0.01107f
C466 B.n223 VSUBS 0.01107f
C467 B.n224 VSUBS 0.01107f
C468 B.n225 VSUBS 0.01107f
C469 B.n226 VSUBS 0.01107f
C470 B.n227 VSUBS 0.01107f
C471 B.n228 VSUBS 0.01107f
C472 B.n229 VSUBS 0.01107f
C473 B.n230 VSUBS 0.01107f
C474 B.n231 VSUBS 0.01107f
C475 B.n232 VSUBS 0.01107f
C476 B.n233 VSUBS 0.01107f
C477 B.n234 VSUBS 0.01107f
C478 B.n235 VSUBS 0.01107f
C479 B.n236 VSUBS 0.01107f
C480 B.n237 VSUBS 0.01107f
C481 B.n238 VSUBS 0.01107f
C482 B.n239 VSUBS 0.01107f
C483 B.n240 VSUBS 0.01107f
C484 B.n241 VSUBS 0.01107f
C485 B.n242 VSUBS 0.01107f
C486 B.n243 VSUBS 0.01107f
C487 B.n244 VSUBS 0.01107f
C488 B.n245 VSUBS 0.01107f
C489 B.n246 VSUBS 0.01107f
C490 B.n247 VSUBS 0.01107f
C491 B.n248 VSUBS 0.01107f
C492 B.n249 VSUBS 0.01107f
C493 B.n250 VSUBS 0.01107f
C494 B.n251 VSUBS 0.01107f
C495 B.n252 VSUBS 0.01107f
C496 B.n253 VSUBS 0.01107f
C497 B.n254 VSUBS 0.01107f
C498 B.n255 VSUBS 0.01107f
C499 B.n256 VSUBS 0.01107f
C500 B.n257 VSUBS 0.01107f
C501 B.n258 VSUBS 0.01107f
C502 B.n259 VSUBS 0.01107f
C503 B.n260 VSUBS 0.01107f
C504 B.n261 VSUBS 0.01107f
C505 B.n262 VSUBS 0.01107f
C506 B.n263 VSUBS 0.01107f
C507 B.n264 VSUBS 0.01107f
C508 B.n265 VSUBS 0.01107f
C509 B.n266 VSUBS 0.01107f
C510 B.n267 VSUBS 0.01107f
C511 B.n268 VSUBS 0.01107f
C512 B.n269 VSUBS 0.01107f
C513 B.n270 VSUBS 0.01107f
C514 B.n271 VSUBS 0.01107f
C515 B.n272 VSUBS 0.01107f
C516 B.n273 VSUBS 0.01107f
C517 B.n274 VSUBS 0.01107f
C518 B.n275 VSUBS 0.01107f
C519 B.n276 VSUBS 0.01107f
C520 B.n277 VSUBS 0.01107f
C521 B.n278 VSUBS 0.01107f
C522 B.n279 VSUBS 0.01107f
C523 B.n280 VSUBS 0.01107f
C524 B.n281 VSUBS 0.01107f
C525 B.n282 VSUBS 0.01107f
C526 B.n283 VSUBS 0.01107f
C527 B.n284 VSUBS 0.01107f
C528 B.n285 VSUBS 0.01107f
C529 B.n286 VSUBS 0.01107f
C530 B.n287 VSUBS 0.01107f
C531 B.n288 VSUBS 0.01107f
C532 B.n289 VSUBS 0.01107f
C533 B.n290 VSUBS 0.01107f
C534 B.n291 VSUBS 0.01107f
C535 B.n292 VSUBS 0.01107f
C536 B.n293 VSUBS 0.01107f
C537 B.n294 VSUBS 0.01107f
C538 B.n295 VSUBS 0.01107f
C539 B.n296 VSUBS 0.01107f
C540 B.n297 VSUBS 0.01107f
C541 B.n298 VSUBS 0.01107f
C542 B.n299 VSUBS 0.01107f
C543 B.n300 VSUBS 0.01107f
C544 B.n301 VSUBS 0.01107f
C545 B.n302 VSUBS 0.01107f
C546 B.n303 VSUBS 0.01107f
C547 B.n304 VSUBS 0.01107f
C548 B.n305 VSUBS 0.01107f
C549 B.n306 VSUBS 0.01107f
C550 B.n307 VSUBS 0.025943f
C551 B.n308 VSUBS 0.026476f
C552 B.n309 VSUBS 0.026476f
C553 B.n310 VSUBS 0.01107f
C554 B.n311 VSUBS 0.01107f
C555 B.n312 VSUBS 0.01107f
C556 B.n313 VSUBS 0.01107f
C557 B.n314 VSUBS 0.01107f
C558 B.n315 VSUBS 0.01107f
C559 B.n316 VSUBS 0.01107f
C560 B.n317 VSUBS 0.01107f
C561 B.n318 VSUBS 0.01107f
C562 B.n319 VSUBS 0.01107f
C563 B.n320 VSUBS 0.01107f
C564 B.n321 VSUBS 0.01107f
C565 B.n322 VSUBS 0.01107f
C566 B.n323 VSUBS 0.01107f
C567 B.n324 VSUBS 0.01107f
C568 B.n325 VSUBS 0.01107f
C569 B.n326 VSUBS 0.01107f
C570 B.n327 VSUBS 0.01107f
C571 B.n328 VSUBS 0.01107f
C572 B.n329 VSUBS 0.01107f
C573 B.n330 VSUBS 0.01107f
C574 B.n331 VSUBS 0.01107f
C575 B.n332 VSUBS 0.01107f
C576 B.n333 VSUBS 0.01107f
C577 B.n334 VSUBS 0.01107f
C578 B.n335 VSUBS 0.01107f
C579 B.n336 VSUBS 0.01107f
C580 B.n337 VSUBS 0.01107f
C581 B.n338 VSUBS 0.01107f
C582 B.n339 VSUBS 0.01107f
C583 B.n340 VSUBS 0.01107f
C584 B.n341 VSUBS 0.01107f
C585 B.n342 VSUBS 0.01107f
C586 B.n343 VSUBS 0.01107f
C587 B.n344 VSUBS 0.01107f
C588 B.n345 VSUBS 0.01107f
C589 B.n346 VSUBS 0.01107f
C590 B.n347 VSUBS 0.010419f
C591 B.n348 VSUBS 0.01107f
C592 B.n349 VSUBS 0.01107f
C593 B.n350 VSUBS 0.006186f
C594 B.n351 VSUBS 0.01107f
C595 B.n352 VSUBS 0.01107f
C596 B.n353 VSUBS 0.01107f
C597 B.n354 VSUBS 0.01107f
C598 B.n355 VSUBS 0.01107f
C599 B.n356 VSUBS 0.01107f
C600 B.n357 VSUBS 0.01107f
C601 B.n358 VSUBS 0.01107f
C602 B.n359 VSUBS 0.01107f
C603 B.n360 VSUBS 0.01107f
C604 B.n361 VSUBS 0.01107f
C605 B.n362 VSUBS 0.01107f
C606 B.n363 VSUBS 0.006186f
C607 B.n364 VSUBS 0.025648f
C608 B.n365 VSUBS 0.010419f
C609 B.n366 VSUBS 0.01107f
C610 B.n367 VSUBS 0.01107f
C611 B.n368 VSUBS 0.01107f
C612 B.n369 VSUBS 0.01107f
C613 B.n370 VSUBS 0.01107f
C614 B.n371 VSUBS 0.01107f
C615 B.n372 VSUBS 0.01107f
C616 B.n373 VSUBS 0.01107f
C617 B.n374 VSUBS 0.01107f
C618 B.n375 VSUBS 0.01107f
C619 B.n376 VSUBS 0.01107f
C620 B.n377 VSUBS 0.01107f
C621 B.n378 VSUBS 0.01107f
C622 B.n379 VSUBS 0.01107f
C623 B.n380 VSUBS 0.01107f
C624 B.n381 VSUBS 0.01107f
C625 B.n382 VSUBS 0.01107f
C626 B.n383 VSUBS 0.01107f
C627 B.n384 VSUBS 0.01107f
C628 B.n385 VSUBS 0.01107f
C629 B.n386 VSUBS 0.01107f
C630 B.n387 VSUBS 0.01107f
C631 B.n388 VSUBS 0.01107f
C632 B.n389 VSUBS 0.01107f
C633 B.n390 VSUBS 0.01107f
C634 B.n391 VSUBS 0.01107f
C635 B.n392 VSUBS 0.01107f
C636 B.n393 VSUBS 0.01107f
C637 B.n394 VSUBS 0.01107f
C638 B.n395 VSUBS 0.01107f
C639 B.n396 VSUBS 0.01107f
C640 B.n397 VSUBS 0.01107f
C641 B.n398 VSUBS 0.01107f
C642 B.n399 VSUBS 0.01107f
C643 B.n400 VSUBS 0.01107f
C644 B.n401 VSUBS 0.01107f
C645 B.n402 VSUBS 0.01107f
C646 B.n403 VSUBS 0.01107f
C647 B.n404 VSUBS 0.026476f
C648 B.n405 VSUBS 0.026476f
C649 B.n406 VSUBS 0.025943f
C650 B.n407 VSUBS 0.01107f
C651 B.n408 VSUBS 0.01107f
C652 B.n409 VSUBS 0.01107f
C653 B.n410 VSUBS 0.01107f
C654 B.n411 VSUBS 0.01107f
C655 B.n412 VSUBS 0.01107f
C656 B.n413 VSUBS 0.01107f
C657 B.n414 VSUBS 0.01107f
C658 B.n415 VSUBS 0.01107f
C659 B.n416 VSUBS 0.01107f
C660 B.n417 VSUBS 0.01107f
C661 B.n418 VSUBS 0.01107f
C662 B.n419 VSUBS 0.01107f
C663 B.n420 VSUBS 0.01107f
C664 B.n421 VSUBS 0.01107f
C665 B.n422 VSUBS 0.01107f
C666 B.n423 VSUBS 0.01107f
C667 B.n424 VSUBS 0.01107f
C668 B.n425 VSUBS 0.01107f
C669 B.n426 VSUBS 0.01107f
C670 B.n427 VSUBS 0.01107f
C671 B.n428 VSUBS 0.01107f
C672 B.n429 VSUBS 0.01107f
C673 B.n430 VSUBS 0.01107f
C674 B.n431 VSUBS 0.01107f
C675 B.n432 VSUBS 0.01107f
C676 B.n433 VSUBS 0.01107f
C677 B.n434 VSUBS 0.01107f
C678 B.n435 VSUBS 0.01107f
C679 B.n436 VSUBS 0.01107f
C680 B.n437 VSUBS 0.01107f
C681 B.n438 VSUBS 0.01107f
C682 B.n439 VSUBS 0.01107f
C683 B.n440 VSUBS 0.01107f
C684 B.n441 VSUBS 0.01107f
C685 B.n442 VSUBS 0.01107f
C686 B.n443 VSUBS 0.01107f
C687 B.n444 VSUBS 0.01107f
C688 B.n445 VSUBS 0.01107f
C689 B.n446 VSUBS 0.01107f
C690 B.n447 VSUBS 0.01107f
C691 B.n448 VSUBS 0.01107f
C692 B.n449 VSUBS 0.01107f
C693 B.n450 VSUBS 0.01107f
C694 B.n451 VSUBS 0.01107f
C695 B.n452 VSUBS 0.01107f
C696 B.n453 VSUBS 0.01107f
C697 B.n454 VSUBS 0.01107f
C698 B.n455 VSUBS 0.01107f
C699 B.n456 VSUBS 0.01107f
C700 B.n457 VSUBS 0.01107f
C701 B.n458 VSUBS 0.01107f
C702 B.n459 VSUBS 0.01107f
C703 B.n460 VSUBS 0.01107f
C704 B.n461 VSUBS 0.01107f
C705 B.n462 VSUBS 0.01107f
C706 B.n463 VSUBS 0.01107f
C707 B.n464 VSUBS 0.01107f
C708 B.n465 VSUBS 0.01107f
C709 B.n466 VSUBS 0.01107f
C710 B.n467 VSUBS 0.01107f
C711 B.n468 VSUBS 0.01107f
C712 B.n469 VSUBS 0.01107f
C713 B.n470 VSUBS 0.01107f
C714 B.n471 VSUBS 0.01107f
C715 B.n472 VSUBS 0.01107f
C716 B.n473 VSUBS 0.01107f
C717 B.n474 VSUBS 0.01107f
C718 B.n475 VSUBS 0.01107f
C719 B.n476 VSUBS 0.01107f
C720 B.n477 VSUBS 0.01107f
C721 B.n478 VSUBS 0.01107f
C722 B.n479 VSUBS 0.01107f
C723 B.n480 VSUBS 0.01107f
C724 B.n481 VSUBS 0.01107f
C725 B.n482 VSUBS 0.01107f
C726 B.n483 VSUBS 0.01107f
C727 B.n484 VSUBS 0.01107f
C728 B.n485 VSUBS 0.01107f
C729 B.n486 VSUBS 0.01107f
C730 B.n487 VSUBS 0.01107f
C731 B.n488 VSUBS 0.01107f
C732 B.n489 VSUBS 0.01107f
C733 B.n490 VSUBS 0.01107f
C734 B.n491 VSUBS 0.01107f
C735 B.n492 VSUBS 0.01107f
C736 B.n493 VSUBS 0.01107f
C737 B.n494 VSUBS 0.01107f
C738 B.n495 VSUBS 0.01107f
C739 B.n496 VSUBS 0.01107f
C740 B.n497 VSUBS 0.01107f
C741 B.n498 VSUBS 0.01107f
C742 B.n499 VSUBS 0.01107f
C743 B.n500 VSUBS 0.01107f
C744 B.n501 VSUBS 0.01107f
C745 B.n502 VSUBS 0.01107f
C746 B.n503 VSUBS 0.01107f
C747 B.n504 VSUBS 0.01107f
C748 B.n505 VSUBS 0.01107f
C749 B.n506 VSUBS 0.01107f
C750 B.n507 VSUBS 0.01107f
C751 B.n508 VSUBS 0.01107f
C752 B.n509 VSUBS 0.01107f
C753 B.n510 VSUBS 0.01107f
C754 B.n511 VSUBS 0.01107f
C755 B.n512 VSUBS 0.01107f
C756 B.n513 VSUBS 0.01107f
C757 B.n514 VSUBS 0.01107f
C758 B.n515 VSUBS 0.01107f
C759 B.n516 VSUBS 0.01107f
C760 B.n517 VSUBS 0.01107f
C761 B.n518 VSUBS 0.01107f
C762 B.n519 VSUBS 0.01107f
C763 B.n520 VSUBS 0.01107f
C764 B.n521 VSUBS 0.01107f
C765 B.n522 VSUBS 0.01107f
C766 B.n523 VSUBS 0.01107f
C767 B.n524 VSUBS 0.01107f
C768 B.n525 VSUBS 0.01107f
C769 B.n526 VSUBS 0.01107f
C770 B.n527 VSUBS 0.01107f
C771 B.n528 VSUBS 0.01107f
C772 B.n529 VSUBS 0.01107f
C773 B.n530 VSUBS 0.01107f
C774 B.n531 VSUBS 0.01107f
C775 B.n532 VSUBS 0.01107f
C776 B.n533 VSUBS 0.01107f
C777 B.n534 VSUBS 0.01107f
C778 B.n535 VSUBS 0.01107f
C779 B.n536 VSUBS 0.01107f
C780 B.n537 VSUBS 0.01107f
C781 B.n538 VSUBS 0.01107f
C782 B.n539 VSUBS 0.01107f
C783 B.n540 VSUBS 0.01107f
C784 B.n541 VSUBS 0.01107f
C785 B.n542 VSUBS 0.01107f
C786 B.n543 VSUBS 0.01107f
C787 B.n544 VSUBS 0.01107f
C788 B.n545 VSUBS 0.01107f
C789 B.n546 VSUBS 0.01107f
C790 B.n547 VSUBS 0.01107f
C791 B.n548 VSUBS 0.01107f
C792 B.n549 VSUBS 0.01107f
C793 B.n550 VSUBS 0.01107f
C794 B.n551 VSUBS 0.01107f
C795 B.n552 VSUBS 0.01107f
C796 B.n553 VSUBS 0.01107f
C797 B.n554 VSUBS 0.01107f
C798 B.n555 VSUBS 0.01107f
C799 B.n556 VSUBS 0.01107f
C800 B.n557 VSUBS 0.01107f
C801 B.n558 VSUBS 0.01107f
C802 B.n559 VSUBS 0.01107f
C803 B.n560 VSUBS 0.01107f
C804 B.n561 VSUBS 0.01107f
C805 B.n562 VSUBS 0.01107f
C806 B.n563 VSUBS 0.01107f
C807 B.n564 VSUBS 0.01107f
C808 B.n565 VSUBS 0.01107f
C809 B.n566 VSUBS 0.01107f
C810 B.n567 VSUBS 0.01107f
C811 B.n568 VSUBS 0.01107f
C812 B.n569 VSUBS 0.01107f
C813 B.n570 VSUBS 0.01107f
C814 B.n571 VSUBS 0.01107f
C815 B.n572 VSUBS 0.01107f
C816 B.n573 VSUBS 0.01107f
C817 B.n574 VSUBS 0.01107f
C818 B.n575 VSUBS 0.01107f
C819 B.n576 VSUBS 0.01107f
C820 B.n577 VSUBS 0.01107f
C821 B.n578 VSUBS 0.01107f
C822 B.n579 VSUBS 0.01107f
C823 B.n580 VSUBS 0.01107f
C824 B.n581 VSUBS 0.01107f
C825 B.n582 VSUBS 0.01107f
C826 B.n583 VSUBS 0.01107f
C827 B.n584 VSUBS 0.01107f
C828 B.n585 VSUBS 0.01107f
C829 B.n586 VSUBS 0.01107f
C830 B.n587 VSUBS 0.01107f
C831 B.n588 VSUBS 0.01107f
C832 B.n589 VSUBS 0.01107f
C833 B.n590 VSUBS 0.01107f
C834 B.n591 VSUBS 0.01107f
C835 B.n592 VSUBS 0.01107f
C836 B.n593 VSUBS 0.01107f
C837 B.n594 VSUBS 0.01107f
C838 B.n595 VSUBS 0.01107f
C839 B.n596 VSUBS 0.01107f
C840 B.n597 VSUBS 0.01107f
C841 B.n598 VSUBS 0.01107f
C842 B.n599 VSUBS 0.01107f
C843 B.n600 VSUBS 0.01107f
C844 B.n601 VSUBS 0.01107f
C845 B.n602 VSUBS 0.01107f
C846 B.n603 VSUBS 0.01107f
C847 B.n604 VSUBS 0.01107f
C848 B.n605 VSUBS 0.01107f
C849 B.n606 VSUBS 0.01107f
C850 B.n607 VSUBS 0.025943f
C851 B.n608 VSUBS 0.026476f
C852 B.n609 VSUBS 0.025191f
C853 B.n610 VSUBS 0.01107f
C854 B.n611 VSUBS 0.01107f
C855 B.n612 VSUBS 0.01107f
C856 B.n613 VSUBS 0.01107f
C857 B.n614 VSUBS 0.01107f
C858 B.n615 VSUBS 0.01107f
C859 B.n616 VSUBS 0.01107f
C860 B.n617 VSUBS 0.01107f
C861 B.n618 VSUBS 0.01107f
C862 B.n619 VSUBS 0.01107f
C863 B.n620 VSUBS 0.01107f
C864 B.n621 VSUBS 0.01107f
C865 B.n622 VSUBS 0.01107f
C866 B.n623 VSUBS 0.01107f
C867 B.n624 VSUBS 0.01107f
C868 B.n625 VSUBS 0.01107f
C869 B.n626 VSUBS 0.01107f
C870 B.n627 VSUBS 0.01107f
C871 B.n628 VSUBS 0.01107f
C872 B.n629 VSUBS 0.01107f
C873 B.n630 VSUBS 0.01107f
C874 B.n631 VSUBS 0.01107f
C875 B.n632 VSUBS 0.01107f
C876 B.n633 VSUBS 0.01107f
C877 B.n634 VSUBS 0.01107f
C878 B.n635 VSUBS 0.01107f
C879 B.n636 VSUBS 0.01107f
C880 B.n637 VSUBS 0.01107f
C881 B.n638 VSUBS 0.01107f
C882 B.n639 VSUBS 0.01107f
C883 B.n640 VSUBS 0.01107f
C884 B.n641 VSUBS 0.01107f
C885 B.n642 VSUBS 0.01107f
C886 B.n643 VSUBS 0.01107f
C887 B.n644 VSUBS 0.01107f
C888 B.n645 VSUBS 0.01107f
C889 B.n646 VSUBS 0.01107f
C890 B.n647 VSUBS 0.010419f
C891 B.n648 VSUBS 0.01107f
C892 B.n649 VSUBS 0.01107f
C893 B.n650 VSUBS 0.006186f
C894 B.n651 VSUBS 0.01107f
C895 B.n652 VSUBS 0.01107f
C896 B.n653 VSUBS 0.01107f
C897 B.n654 VSUBS 0.01107f
C898 B.n655 VSUBS 0.01107f
C899 B.n656 VSUBS 0.01107f
C900 B.n657 VSUBS 0.01107f
C901 B.n658 VSUBS 0.01107f
C902 B.n659 VSUBS 0.01107f
C903 B.n660 VSUBS 0.01107f
C904 B.n661 VSUBS 0.01107f
C905 B.n662 VSUBS 0.01107f
C906 B.n663 VSUBS 0.006186f
C907 B.n664 VSUBS 0.025648f
C908 B.n665 VSUBS 0.010419f
C909 B.n666 VSUBS 0.01107f
C910 B.n667 VSUBS 0.01107f
C911 B.n668 VSUBS 0.01107f
C912 B.n669 VSUBS 0.01107f
C913 B.n670 VSUBS 0.01107f
C914 B.n671 VSUBS 0.01107f
C915 B.n672 VSUBS 0.01107f
C916 B.n673 VSUBS 0.01107f
C917 B.n674 VSUBS 0.01107f
C918 B.n675 VSUBS 0.01107f
C919 B.n676 VSUBS 0.01107f
C920 B.n677 VSUBS 0.01107f
C921 B.n678 VSUBS 0.01107f
C922 B.n679 VSUBS 0.01107f
C923 B.n680 VSUBS 0.01107f
C924 B.n681 VSUBS 0.01107f
C925 B.n682 VSUBS 0.01107f
C926 B.n683 VSUBS 0.01107f
C927 B.n684 VSUBS 0.01107f
C928 B.n685 VSUBS 0.01107f
C929 B.n686 VSUBS 0.01107f
C930 B.n687 VSUBS 0.01107f
C931 B.n688 VSUBS 0.01107f
C932 B.n689 VSUBS 0.01107f
C933 B.n690 VSUBS 0.01107f
C934 B.n691 VSUBS 0.01107f
C935 B.n692 VSUBS 0.01107f
C936 B.n693 VSUBS 0.01107f
C937 B.n694 VSUBS 0.01107f
C938 B.n695 VSUBS 0.01107f
C939 B.n696 VSUBS 0.01107f
C940 B.n697 VSUBS 0.01107f
C941 B.n698 VSUBS 0.01107f
C942 B.n699 VSUBS 0.01107f
C943 B.n700 VSUBS 0.01107f
C944 B.n701 VSUBS 0.01107f
C945 B.n702 VSUBS 0.01107f
C946 B.n703 VSUBS 0.01107f
C947 B.n704 VSUBS 0.026476f
C948 B.n705 VSUBS 0.026476f
C949 B.n706 VSUBS 0.025943f
C950 B.n707 VSUBS 0.01107f
C951 B.n708 VSUBS 0.01107f
C952 B.n709 VSUBS 0.01107f
C953 B.n710 VSUBS 0.01107f
C954 B.n711 VSUBS 0.01107f
C955 B.n712 VSUBS 0.01107f
C956 B.n713 VSUBS 0.01107f
C957 B.n714 VSUBS 0.01107f
C958 B.n715 VSUBS 0.01107f
C959 B.n716 VSUBS 0.01107f
C960 B.n717 VSUBS 0.01107f
C961 B.n718 VSUBS 0.01107f
C962 B.n719 VSUBS 0.01107f
C963 B.n720 VSUBS 0.01107f
C964 B.n721 VSUBS 0.01107f
C965 B.n722 VSUBS 0.01107f
C966 B.n723 VSUBS 0.01107f
C967 B.n724 VSUBS 0.01107f
C968 B.n725 VSUBS 0.01107f
C969 B.n726 VSUBS 0.01107f
C970 B.n727 VSUBS 0.01107f
C971 B.n728 VSUBS 0.01107f
C972 B.n729 VSUBS 0.01107f
C973 B.n730 VSUBS 0.01107f
C974 B.n731 VSUBS 0.01107f
C975 B.n732 VSUBS 0.01107f
C976 B.n733 VSUBS 0.01107f
C977 B.n734 VSUBS 0.01107f
C978 B.n735 VSUBS 0.01107f
C979 B.n736 VSUBS 0.01107f
C980 B.n737 VSUBS 0.01107f
C981 B.n738 VSUBS 0.01107f
C982 B.n739 VSUBS 0.01107f
C983 B.n740 VSUBS 0.01107f
C984 B.n741 VSUBS 0.01107f
C985 B.n742 VSUBS 0.01107f
C986 B.n743 VSUBS 0.01107f
C987 B.n744 VSUBS 0.01107f
C988 B.n745 VSUBS 0.01107f
C989 B.n746 VSUBS 0.01107f
C990 B.n747 VSUBS 0.01107f
C991 B.n748 VSUBS 0.01107f
C992 B.n749 VSUBS 0.01107f
C993 B.n750 VSUBS 0.01107f
C994 B.n751 VSUBS 0.01107f
C995 B.n752 VSUBS 0.01107f
C996 B.n753 VSUBS 0.01107f
C997 B.n754 VSUBS 0.01107f
C998 B.n755 VSUBS 0.01107f
C999 B.n756 VSUBS 0.01107f
C1000 B.n757 VSUBS 0.01107f
C1001 B.n758 VSUBS 0.01107f
C1002 B.n759 VSUBS 0.01107f
C1003 B.n760 VSUBS 0.01107f
C1004 B.n761 VSUBS 0.01107f
C1005 B.n762 VSUBS 0.01107f
C1006 B.n763 VSUBS 0.01107f
C1007 B.n764 VSUBS 0.01107f
C1008 B.n765 VSUBS 0.01107f
C1009 B.n766 VSUBS 0.01107f
C1010 B.n767 VSUBS 0.01107f
C1011 B.n768 VSUBS 0.01107f
C1012 B.n769 VSUBS 0.01107f
C1013 B.n770 VSUBS 0.01107f
C1014 B.n771 VSUBS 0.01107f
C1015 B.n772 VSUBS 0.01107f
C1016 B.n773 VSUBS 0.01107f
C1017 B.n774 VSUBS 0.01107f
C1018 B.n775 VSUBS 0.01107f
C1019 B.n776 VSUBS 0.01107f
C1020 B.n777 VSUBS 0.01107f
C1021 B.n778 VSUBS 0.01107f
C1022 B.n779 VSUBS 0.01107f
C1023 B.n780 VSUBS 0.01107f
C1024 B.n781 VSUBS 0.01107f
C1025 B.n782 VSUBS 0.01107f
C1026 B.n783 VSUBS 0.01107f
C1027 B.n784 VSUBS 0.01107f
C1028 B.n785 VSUBS 0.01107f
C1029 B.n786 VSUBS 0.01107f
C1030 B.n787 VSUBS 0.01107f
C1031 B.n788 VSUBS 0.01107f
C1032 B.n789 VSUBS 0.01107f
C1033 B.n790 VSUBS 0.01107f
C1034 B.n791 VSUBS 0.01107f
C1035 B.n792 VSUBS 0.01107f
C1036 B.n793 VSUBS 0.01107f
C1037 B.n794 VSUBS 0.01107f
C1038 B.n795 VSUBS 0.01107f
C1039 B.n796 VSUBS 0.01107f
C1040 B.n797 VSUBS 0.01107f
C1041 B.n798 VSUBS 0.01107f
C1042 B.n799 VSUBS 0.01107f
C1043 B.n800 VSUBS 0.01107f
C1044 B.n801 VSUBS 0.01107f
C1045 B.n802 VSUBS 0.01107f
C1046 B.n803 VSUBS 0.01107f
C1047 B.n804 VSUBS 0.01107f
C1048 B.n805 VSUBS 0.01107f
C1049 B.n806 VSUBS 0.01107f
C1050 B.n807 VSUBS 0.025066f
C1051 VDD2.n0 VSUBS 0.034989f
C1052 VDD2.n1 VSUBS 0.033477f
C1053 VDD2.n2 VSUBS 0.017989f
C1054 VDD2.n3 VSUBS 0.042519f
C1055 VDD2.n4 VSUBS 0.019047f
C1056 VDD2.n5 VSUBS 0.033477f
C1057 VDD2.n6 VSUBS 0.017989f
C1058 VDD2.n7 VSUBS 0.042519f
C1059 VDD2.n8 VSUBS 0.019047f
C1060 VDD2.n9 VSUBS 0.935947f
C1061 VDD2.n10 VSUBS 0.017989f
C1062 VDD2.t0 VSUBS 0.091291f
C1063 VDD2.n11 VSUBS 0.190712f
C1064 VDD2.n12 VSUBS 0.031983f
C1065 VDD2.n13 VSUBS 0.031889f
C1066 VDD2.n14 VSUBS 0.042519f
C1067 VDD2.n15 VSUBS 0.019047f
C1068 VDD2.n16 VSUBS 0.017989f
C1069 VDD2.n17 VSUBS 0.033477f
C1070 VDD2.n18 VSUBS 0.033477f
C1071 VDD2.n19 VSUBS 0.017989f
C1072 VDD2.n20 VSUBS 0.019047f
C1073 VDD2.n21 VSUBS 0.042519f
C1074 VDD2.n22 VSUBS 0.042519f
C1075 VDD2.n23 VSUBS 0.019047f
C1076 VDD2.n24 VSUBS 0.017989f
C1077 VDD2.n25 VSUBS 0.033477f
C1078 VDD2.n26 VSUBS 0.033477f
C1079 VDD2.n27 VSUBS 0.017989f
C1080 VDD2.n28 VSUBS 0.019047f
C1081 VDD2.n29 VSUBS 0.042519f
C1082 VDD2.n30 VSUBS 0.103656f
C1083 VDD2.n31 VSUBS 0.019047f
C1084 VDD2.n32 VSUBS 0.035326f
C1085 VDD2.n33 VSUBS 0.081495f
C1086 VDD2.n34 VSUBS 0.12164f
C1087 VDD2.t4 VSUBS 0.189676f
C1088 VDD2.t7 VSUBS 0.189676f
C1089 VDD2.n35 VSUBS 1.339f
C1090 VDD2.n36 VSUBS 1.28952f
C1091 VDD2.t3 VSUBS 0.189676f
C1092 VDD2.t9 VSUBS 0.189676f
C1093 VDD2.n37 VSUBS 1.36504f
C1094 VDD2.n38 VSUBS 4.04916f
C1095 VDD2.n39 VSUBS 0.034989f
C1096 VDD2.n40 VSUBS 0.033477f
C1097 VDD2.n41 VSUBS 0.017989f
C1098 VDD2.n42 VSUBS 0.042519f
C1099 VDD2.n43 VSUBS 0.019047f
C1100 VDD2.n44 VSUBS 0.033477f
C1101 VDD2.n45 VSUBS 0.017989f
C1102 VDD2.n46 VSUBS 0.042519f
C1103 VDD2.n47 VSUBS 0.019047f
C1104 VDD2.n48 VSUBS 0.935947f
C1105 VDD2.n49 VSUBS 0.017989f
C1106 VDD2.t1 VSUBS 0.091291f
C1107 VDD2.n50 VSUBS 0.190712f
C1108 VDD2.n51 VSUBS 0.031983f
C1109 VDD2.n52 VSUBS 0.031889f
C1110 VDD2.n53 VSUBS 0.042519f
C1111 VDD2.n54 VSUBS 0.019047f
C1112 VDD2.n55 VSUBS 0.017989f
C1113 VDD2.n56 VSUBS 0.033477f
C1114 VDD2.n57 VSUBS 0.033477f
C1115 VDD2.n58 VSUBS 0.017989f
C1116 VDD2.n59 VSUBS 0.019047f
C1117 VDD2.n60 VSUBS 0.042519f
C1118 VDD2.n61 VSUBS 0.042519f
C1119 VDD2.n62 VSUBS 0.019047f
C1120 VDD2.n63 VSUBS 0.017989f
C1121 VDD2.n64 VSUBS 0.033477f
C1122 VDD2.n65 VSUBS 0.033477f
C1123 VDD2.n66 VSUBS 0.017989f
C1124 VDD2.n67 VSUBS 0.019047f
C1125 VDD2.n68 VSUBS 0.042519f
C1126 VDD2.n69 VSUBS 0.103656f
C1127 VDD2.n70 VSUBS 0.019047f
C1128 VDD2.n71 VSUBS 0.035326f
C1129 VDD2.n72 VSUBS 0.081495f
C1130 VDD2.n73 VSUBS 0.101431f
C1131 VDD2.n74 VSUBS 3.5797f
C1132 VDD2.t2 VSUBS 0.189676f
C1133 VDD2.t8 VSUBS 0.189676f
C1134 VDD2.n75 VSUBS 1.33901f
C1135 VDD2.n76 VSUBS 0.944324f
C1136 VDD2.t5 VSUBS 0.189676f
C1137 VDD2.t6 VSUBS 0.189676f
C1138 VDD2.n77 VSUBS 1.36499f
C1139 VTAIL.t13 VSUBS 0.184577f
C1140 VTAIL.t11 VSUBS 0.184577f
C1141 VTAIL.n0 VSUBS 1.17655f
C1142 VTAIL.n1 VSUBS 1.05043f
C1143 VTAIL.n2 VSUBS 0.034048f
C1144 VTAIL.n3 VSUBS 0.032577f
C1145 VTAIL.n4 VSUBS 0.017505f
C1146 VTAIL.n5 VSUBS 0.041376f
C1147 VTAIL.n6 VSUBS 0.018535f
C1148 VTAIL.n7 VSUBS 0.032577f
C1149 VTAIL.n8 VSUBS 0.017505f
C1150 VTAIL.n9 VSUBS 0.041376f
C1151 VTAIL.n10 VSUBS 0.018535f
C1152 VTAIL.n11 VSUBS 0.910783f
C1153 VTAIL.n12 VSUBS 0.017505f
C1154 VTAIL.t6 VSUBS 0.088837f
C1155 VTAIL.n13 VSUBS 0.185585f
C1156 VTAIL.n14 VSUBS 0.031124f
C1157 VTAIL.n15 VSUBS 0.031032f
C1158 VTAIL.n16 VSUBS 0.041376f
C1159 VTAIL.n17 VSUBS 0.018535f
C1160 VTAIL.n18 VSUBS 0.017505f
C1161 VTAIL.n19 VSUBS 0.032577f
C1162 VTAIL.n20 VSUBS 0.032577f
C1163 VTAIL.n21 VSUBS 0.017505f
C1164 VTAIL.n22 VSUBS 0.018535f
C1165 VTAIL.n23 VSUBS 0.041376f
C1166 VTAIL.n24 VSUBS 0.041376f
C1167 VTAIL.n25 VSUBS 0.018535f
C1168 VTAIL.n26 VSUBS 0.017505f
C1169 VTAIL.n27 VSUBS 0.032577f
C1170 VTAIL.n28 VSUBS 0.032577f
C1171 VTAIL.n29 VSUBS 0.017505f
C1172 VTAIL.n30 VSUBS 0.018535f
C1173 VTAIL.n31 VSUBS 0.041376f
C1174 VTAIL.n32 VSUBS 0.100869f
C1175 VTAIL.n33 VSUBS 0.018535f
C1176 VTAIL.n34 VSUBS 0.034376f
C1177 VTAIL.n35 VSUBS 0.079304f
C1178 VTAIL.n36 VSUBS 0.076241f
C1179 VTAIL.n37 VSUBS 0.531402f
C1180 VTAIL.t7 VSUBS 0.184577f
C1181 VTAIL.t3 VSUBS 0.184577f
C1182 VTAIL.n38 VSUBS 1.17655f
C1183 VTAIL.n39 VSUBS 1.221f
C1184 VTAIL.t2 VSUBS 0.184577f
C1185 VTAIL.t19 VSUBS 0.184577f
C1186 VTAIL.n40 VSUBS 1.17655f
C1187 VTAIL.n41 VSUBS 2.61366f
C1188 VTAIL.t16 VSUBS 0.184577f
C1189 VTAIL.t12 VSUBS 0.184577f
C1190 VTAIL.n42 VSUBS 1.17656f
C1191 VTAIL.n43 VSUBS 2.61365f
C1192 VTAIL.t10 VSUBS 0.184577f
C1193 VTAIL.t9 VSUBS 0.184577f
C1194 VTAIL.n44 VSUBS 1.17656f
C1195 VTAIL.n45 VSUBS 1.22099f
C1196 VTAIL.n46 VSUBS 0.034048f
C1197 VTAIL.n47 VSUBS 0.032577f
C1198 VTAIL.n48 VSUBS 0.017505f
C1199 VTAIL.n49 VSUBS 0.041376f
C1200 VTAIL.n50 VSUBS 0.018535f
C1201 VTAIL.n51 VSUBS 0.032577f
C1202 VTAIL.n52 VSUBS 0.017505f
C1203 VTAIL.n53 VSUBS 0.041376f
C1204 VTAIL.n54 VSUBS 0.018535f
C1205 VTAIL.n55 VSUBS 0.910783f
C1206 VTAIL.n56 VSUBS 0.017505f
C1207 VTAIL.t18 VSUBS 0.088837f
C1208 VTAIL.n57 VSUBS 0.185585f
C1209 VTAIL.n58 VSUBS 0.031124f
C1210 VTAIL.n59 VSUBS 0.031032f
C1211 VTAIL.n60 VSUBS 0.041376f
C1212 VTAIL.n61 VSUBS 0.018535f
C1213 VTAIL.n62 VSUBS 0.017505f
C1214 VTAIL.n63 VSUBS 0.032577f
C1215 VTAIL.n64 VSUBS 0.032577f
C1216 VTAIL.n65 VSUBS 0.017505f
C1217 VTAIL.n66 VSUBS 0.018535f
C1218 VTAIL.n67 VSUBS 0.041376f
C1219 VTAIL.n68 VSUBS 0.041376f
C1220 VTAIL.n69 VSUBS 0.018535f
C1221 VTAIL.n70 VSUBS 0.017505f
C1222 VTAIL.n71 VSUBS 0.032577f
C1223 VTAIL.n72 VSUBS 0.032577f
C1224 VTAIL.n73 VSUBS 0.017505f
C1225 VTAIL.n74 VSUBS 0.018535f
C1226 VTAIL.n75 VSUBS 0.041376f
C1227 VTAIL.n76 VSUBS 0.100869f
C1228 VTAIL.n77 VSUBS 0.018535f
C1229 VTAIL.n78 VSUBS 0.034376f
C1230 VTAIL.n79 VSUBS 0.079304f
C1231 VTAIL.n80 VSUBS 0.076241f
C1232 VTAIL.n81 VSUBS 0.531402f
C1233 VTAIL.t5 VSUBS 0.184577f
C1234 VTAIL.t8 VSUBS 0.184577f
C1235 VTAIL.n82 VSUBS 1.17656f
C1236 VTAIL.n83 VSUBS 1.11964f
C1237 VTAIL.t1 VSUBS 0.184577f
C1238 VTAIL.t0 VSUBS 0.184577f
C1239 VTAIL.n84 VSUBS 1.17656f
C1240 VTAIL.n85 VSUBS 1.22099f
C1241 VTAIL.n86 VSUBS 0.034048f
C1242 VTAIL.n87 VSUBS 0.032577f
C1243 VTAIL.n88 VSUBS 0.017505f
C1244 VTAIL.n89 VSUBS 0.041376f
C1245 VTAIL.n90 VSUBS 0.018535f
C1246 VTAIL.n91 VSUBS 0.032577f
C1247 VTAIL.n92 VSUBS 0.017505f
C1248 VTAIL.n93 VSUBS 0.041376f
C1249 VTAIL.n94 VSUBS 0.018535f
C1250 VTAIL.n95 VSUBS 0.910783f
C1251 VTAIL.n96 VSUBS 0.017505f
C1252 VTAIL.t4 VSUBS 0.088837f
C1253 VTAIL.n97 VSUBS 0.185585f
C1254 VTAIL.n98 VSUBS 0.031124f
C1255 VTAIL.n99 VSUBS 0.031032f
C1256 VTAIL.n100 VSUBS 0.041376f
C1257 VTAIL.n101 VSUBS 0.018535f
C1258 VTAIL.n102 VSUBS 0.017505f
C1259 VTAIL.n103 VSUBS 0.032577f
C1260 VTAIL.n104 VSUBS 0.032577f
C1261 VTAIL.n105 VSUBS 0.017505f
C1262 VTAIL.n106 VSUBS 0.018535f
C1263 VTAIL.n107 VSUBS 0.041376f
C1264 VTAIL.n108 VSUBS 0.041376f
C1265 VTAIL.n109 VSUBS 0.018535f
C1266 VTAIL.n110 VSUBS 0.017505f
C1267 VTAIL.n111 VSUBS 0.032577f
C1268 VTAIL.n112 VSUBS 0.032577f
C1269 VTAIL.n113 VSUBS 0.017505f
C1270 VTAIL.n114 VSUBS 0.018535f
C1271 VTAIL.n115 VSUBS 0.041376f
C1272 VTAIL.n116 VSUBS 0.100869f
C1273 VTAIL.n117 VSUBS 0.018535f
C1274 VTAIL.n118 VSUBS 0.034376f
C1275 VTAIL.n119 VSUBS 0.079304f
C1276 VTAIL.n120 VSUBS 0.076241f
C1277 VTAIL.n121 VSUBS 1.72408f
C1278 VTAIL.n122 VSUBS 0.034048f
C1279 VTAIL.n123 VSUBS 0.032577f
C1280 VTAIL.n124 VSUBS 0.017505f
C1281 VTAIL.n125 VSUBS 0.041376f
C1282 VTAIL.n126 VSUBS 0.018535f
C1283 VTAIL.n127 VSUBS 0.032577f
C1284 VTAIL.n128 VSUBS 0.017505f
C1285 VTAIL.n129 VSUBS 0.041376f
C1286 VTAIL.n130 VSUBS 0.018535f
C1287 VTAIL.n131 VSUBS 0.910783f
C1288 VTAIL.n132 VSUBS 0.017505f
C1289 VTAIL.t14 VSUBS 0.088837f
C1290 VTAIL.n133 VSUBS 0.185585f
C1291 VTAIL.n134 VSUBS 0.031124f
C1292 VTAIL.n135 VSUBS 0.031032f
C1293 VTAIL.n136 VSUBS 0.041376f
C1294 VTAIL.n137 VSUBS 0.018535f
C1295 VTAIL.n138 VSUBS 0.017505f
C1296 VTAIL.n139 VSUBS 0.032577f
C1297 VTAIL.n140 VSUBS 0.032577f
C1298 VTAIL.n141 VSUBS 0.017505f
C1299 VTAIL.n142 VSUBS 0.018535f
C1300 VTAIL.n143 VSUBS 0.041376f
C1301 VTAIL.n144 VSUBS 0.041376f
C1302 VTAIL.n145 VSUBS 0.018535f
C1303 VTAIL.n146 VSUBS 0.017505f
C1304 VTAIL.n147 VSUBS 0.032577f
C1305 VTAIL.n148 VSUBS 0.032577f
C1306 VTAIL.n149 VSUBS 0.017505f
C1307 VTAIL.n150 VSUBS 0.018535f
C1308 VTAIL.n151 VSUBS 0.041376f
C1309 VTAIL.n152 VSUBS 0.100869f
C1310 VTAIL.n153 VSUBS 0.018535f
C1311 VTAIL.n154 VSUBS 0.034376f
C1312 VTAIL.n155 VSUBS 0.079304f
C1313 VTAIL.n156 VSUBS 0.076241f
C1314 VTAIL.n157 VSUBS 1.72408f
C1315 VTAIL.t15 VSUBS 0.184577f
C1316 VTAIL.t17 VSUBS 0.184577f
C1317 VTAIL.n158 VSUBS 1.17655f
C1318 VTAIL.n159 VSUBS 0.988893f
C1319 VN.t0 VSUBS 1.80755f
C1320 VN.n0 VSUBS 0.785199f
C1321 VN.n1 VSUBS 0.031447f
C1322 VN.n2 VSUBS 0.045472f
C1323 VN.n3 VSUBS 0.031447f
C1324 VN.t6 VSUBS 1.80755f
C1325 VN.n4 VSUBS 0.05861f
C1326 VN.n5 VSUBS 0.031447f
C1327 VN.n6 VSUBS 0.05861f
C1328 VN.n7 VSUBS 0.031447f
C1329 VN.t2 VSUBS 1.80755f
C1330 VN.n8 VSUBS 0.05861f
C1331 VN.n9 VSUBS 0.031447f
C1332 VN.n10 VSUBS 0.034304f
C1333 VN.t5 VSUBS 1.80755f
C1334 VN.n11 VSUBS 0.751523f
C1335 VN.t9 VSUBS 2.11681f
C1336 VN.n12 VSUBS 0.728492f
C1337 VN.n13 VSUBS 0.340095f
C1338 VN.n14 VSUBS 0.031447f
C1339 VN.n15 VSUBS 0.05861f
C1340 VN.n16 VSUBS 0.063353f
C1341 VN.n17 VSUBS 0.028468f
C1342 VN.n18 VSUBS 0.031447f
C1343 VN.n19 VSUBS 0.031447f
C1344 VN.n20 VSUBS 0.031447f
C1345 VN.n21 VSUBS 0.05861f
C1346 VN.n22 VSUBS 0.044142f
C1347 VN.n23 VSUBS 0.660828f
C1348 VN.n24 VSUBS 0.044142f
C1349 VN.n25 VSUBS 0.031447f
C1350 VN.n26 VSUBS 0.031447f
C1351 VN.n27 VSUBS 0.031447f
C1352 VN.n28 VSUBS 0.05861f
C1353 VN.n29 VSUBS 0.028468f
C1354 VN.n30 VSUBS 0.063353f
C1355 VN.n31 VSUBS 0.031447f
C1356 VN.n32 VSUBS 0.031447f
C1357 VN.n33 VSUBS 0.031447f
C1358 VN.n34 VSUBS 0.034304f
C1359 VN.n35 VSUBS 0.660828f
C1360 VN.n36 VSUBS 0.05398f
C1361 VN.n37 VSUBS 0.05861f
C1362 VN.n38 VSUBS 0.031447f
C1363 VN.n39 VSUBS 0.031447f
C1364 VN.n40 VSUBS 0.031447f
C1365 VN.n41 VSUBS 0.046348f
C1366 VN.n42 VSUBS 0.05861f
C1367 VN.n43 VSUBS 0.053401f
C1368 VN.n44 VSUBS 0.050755f
C1369 VN.n45 VSUBS 0.065357f
C1370 VN.t8 VSUBS 1.80755f
C1371 VN.n46 VSUBS 0.785199f
C1372 VN.n47 VSUBS 0.031447f
C1373 VN.n48 VSUBS 0.045472f
C1374 VN.n49 VSUBS 0.031447f
C1375 VN.t7 VSUBS 1.80755f
C1376 VN.n50 VSUBS 0.05861f
C1377 VN.n51 VSUBS 0.031447f
C1378 VN.n52 VSUBS 0.05861f
C1379 VN.n53 VSUBS 0.031447f
C1380 VN.t1 VSUBS 1.80755f
C1381 VN.n54 VSUBS 0.05861f
C1382 VN.n55 VSUBS 0.031447f
C1383 VN.n56 VSUBS 0.034304f
C1384 VN.t3 VSUBS 2.11681f
C1385 VN.t4 VSUBS 1.80755f
C1386 VN.n57 VSUBS 0.751523f
C1387 VN.n58 VSUBS 0.728492f
C1388 VN.n59 VSUBS 0.340095f
C1389 VN.n60 VSUBS 0.031447f
C1390 VN.n61 VSUBS 0.05861f
C1391 VN.n62 VSUBS 0.063353f
C1392 VN.n63 VSUBS 0.028468f
C1393 VN.n64 VSUBS 0.031447f
C1394 VN.n65 VSUBS 0.031447f
C1395 VN.n66 VSUBS 0.031447f
C1396 VN.n67 VSUBS 0.05861f
C1397 VN.n68 VSUBS 0.044142f
C1398 VN.n69 VSUBS 0.660828f
C1399 VN.n70 VSUBS 0.044142f
C1400 VN.n71 VSUBS 0.031447f
C1401 VN.n72 VSUBS 0.031447f
C1402 VN.n73 VSUBS 0.031447f
C1403 VN.n74 VSUBS 0.05861f
C1404 VN.n75 VSUBS 0.028468f
C1405 VN.n76 VSUBS 0.063353f
C1406 VN.n77 VSUBS 0.031447f
C1407 VN.n78 VSUBS 0.031447f
C1408 VN.n79 VSUBS 0.031447f
C1409 VN.n80 VSUBS 0.034304f
C1410 VN.n81 VSUBS 0.660828f
C1411 VN.n82 VSUBS 0.05398f
C1412 VN.n83 VSUBS 0.05861f
C1413 VN.n84 VSUBS 0.031447f
C1414 VN.n85 VSUBS 0.031447f
C1415 VN.n86 VSUBS 0.031447f
C1416 VN.n87 VSUBS 0.046348f
C1417 VN.n88 VSUBS 0.05861f
C1418 VN.n89 VSUBS 0.053401f
C1419 VN.n90 VSUBS 0.050755f
C1420 VN.n91 VSUBS 1.88032f
.ends

