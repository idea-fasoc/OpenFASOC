* NGSPICE file created from diff_pair_sample_1333.ext - technology: sky130A

.subckt diff_pair_sample_1333 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0 ps=0 w=0.52 l=2.97
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0 ps=0 w=0.52 l=2.97
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0 ps=0 w=0.52 l=2.97
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0 ps=0 w=0.52 l=2.97
X4 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0.2028 ps=1.82 w=0.52 l=2.97
X5 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0.2028 ps=1.82 w=0.52 l=2.97
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0.2028 ps=1.82 w=0.52 l=2.97
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2028 pd=1.82 as=0.2028 ps=1.82 w=0.52 l=2.97
R0 B.n355 B.n354 585
R1 B.n356 B.n355 585
R2 B.n116 B.n66 585
R3 B.n115 B.n114 585
R4 B.n113 B.n112 585
R5 B.n111 B.n110 585
R6 B.n109 B.n108 585
R7 B.n107 B.n106 585
R8 B.n105 B.n104 585
R9 B.n102 B.n101 585
R10 B.n100 B.n99 585
R11 B.n98 B.n97 585
R12 B.n96 B.n95 585
R13 B.n94 B.n93 585
R14 B.n92 B.n91 585
R15 B.n90 B.n89 585
R16 B.n88 B.n87 585
R17 B.n86 B.n85 585
R18 B.n84 B.n83 585
R19 B.n82 B.n81 585
R20 B.n80 B.n79 585
R21 B.n78 B.n77 585
R22 B.n76 B.n75 585
R23 B.n74 B.n73 585
R24 B.n54 B.n53 585
R25 B.n359 B.n358 585
R26 B.n353 B.n67 585
R27 B.n67 B.n51 585
R28 B.n352 B.n50 585
R29 B.n363 B.n50 585
R30 B.n351 B.n49 585
R31 B.n364 B.n49 585
R32 B.n350 B.n48 585
R33 B.n365 B.n48 585
R34 B.n349 B.n348 585
R35 B.n348 B.n44 585
R36 B.n347 B.n43 585
R37 B.n371 B.n43 585
R38 B.n346 B.n42 585
R39 B.n372 B.n42 585
R40 B.n345 B.n41 585
R41 B.n373 B.n41 585
R42 B.n344 B.n343 585
R43 B.n343 B.n40 585
R44 B.n342 B.n36 585
R45 B.n379 B.n36 585
R46 B.n341 B.n35 585
R47 B.n380 B.n35 585
R48 B.n340 B.n34 585
R49 B.n381 B.n34 585
R50 B.n339 B.n338 585
R51 B.n338 B.n30 585
R52 B.n337 B.n29 585
R53 B.n387 B.n29 585
R54 B.n336 B.n28 585
R55 B.n388 B.n28 585
R56 B.n335 B.n27 585
R57 B.n389 B.n27 585
R58 B.n334 B.n333 585
R59 B.n333 B.n23 585
R60 B.n332 B.n22 585
R61 B.n395 B.n22 585
R62 B.n331 B.n21 585
R63 B.n396 B.n21 585
R64 B.n330 B.n20 585
R65 B.n397 B.n20 585
R66 B.n329 B.n328 585
R67 B.n328 B.n16 585
R68 B.n327 B.n15 585
R69 B.n403 B.n15 585
R70 B.n326 B.n14 585
R71 B.n404 B.n14 585
R72 B.n325 B.n13 585
R73 B.n405 B.n13 585
R74 B.n324 B.n323 585
R75 B.n323 B.n12 585
R76 B.n322 B.n321 585
R77 B.n322 B.n8 585
R78 B.n320 B.n7 585
R79 B.n412 B.n7 585
R80 B.n319 B.n6 585
R81 B.n413 B.n6 585
R82 B.n318 B.n5 585
R83 B.n414 B.n5 585
R84 B.n317 B.n316 585
R85 B.n316 B.n4 585
R86 B.n315 B.n117 585
R87 B.n315 B.n314 585
R88 B.n305 B.n118 585
R89 B.n119 B.n118 585
R90 B.n307 B.n306 585
R91 B.n308 B.n307 585
R92 B.n304 B.n124 585
R93 B.n124 B.n123 585
R94 B.n303 B.n302 585
R95 B.n302 B.n301 585
R96 B.n126 B.n125 585
R97 B.n127 B.n126 585
R98 B.n294 B.n293 585
R99 B.n295 B.n294 585
R100 B.n292 B.n132 585
R101 B.n132 B.n131 585
R102 B.n291 B.n290 585
R103 B.n290 B.n289 585
R104 B.n134 B.n133 585
R105 B.n135 B.n134 585
R106 B.n282 B.n281 585
R107 B.n283 B.n282 585
R108 B.n280 B.n140 585
R109 B.n140 B.n139 585
R110 B.n279 B.n278 585
R111 B.n278 B.n277 585
R112 B.n142 B.n141 585
R113 B.n143 B.n142 585
R114 B.n270 B.n269 585
R115 B.n271 B.n270 585
R116 B.n268 B.n148 585
R117 B.n148 B.n147 585
R118 B.n267 B.n266 585
R119 B.n266 B.n265 585
R120 B.n150 B.n149 585
R121 B.n258 B.n150 585
R122 B.n257 B.n256 585
R123 B.n259 B.n257 585
R124 B.n255 B.n155 585
R125 B.n155 B.n154 585
R126 B.n254 B.n253 585
R127 B.n253 B.n252 585
R128 B.n157 B.n156 585
R129 B.n158 B.n157 585
R130 B.n245 B.n244 585
R131 B.n246 B.n245 585
R132 B.n243 B.n163 585
R133 B.n163 B.n162 585
R134 B.n242 B.n241 585
R135 B.n241 B.n240 585
R136 B.n165 B.n164 585
R137 B.n166 B.n165 585
R138 B.n236 B.n235 585
R139 B.n169 B.n168 585
R140 B.n232 B.n231 585
R141 B.n233 B.n232 585
R142 B.n230 B.n181 585
R143 B.n229 B.n228 585
R144 B.n227 B.n226 585
R145 B.n225 B.n224 585
R146 B.n223 B.n222 585
R147 B.n220 B.n219 585
R148 B.n218 B.n217 585
R149 B.n216 B.n215 585
R150 B.n214 B.n213 585
R151 B.n212 B.n211 585
R152 B.n210 B.n209 585
R153 B.n208 B.n207 585
R154 B.n206 B.n205 585
R155 B.n204 B.n203 585
R156 B.n202 B.n201 585
R157 B.n200 B.n199 585
R158 B.n198 B.n197 585
R159 B.n196 B.n195 585
R160 B.n194 B.n193 585
R161 B.n192 B.n191 585
R162 B.n190 B.n189 585
R163 B.n188 B.n187 585
R164 B.n237 B.n167 585
R165 B.n167 B.n166 585
R166 B.n239 B.n238 585
R167 B.n240 B.n239 585
R168 B.n161 B.n160 585
R169 B.n162 B.n161 585
R170 B.n248 B.n247 585
R171 B.n247 B.n246 585
R172 B.n249 B.n159 585
R173 B.n159 B.n158 585
R174 B.n251 B.n250 585
R175 B.n252 B.n251 585
R176 B.n153 B.n152 585
R177 B.n154 B.n153 585
R178 B.n261 B.n260 585
R179 B.n260 B.n259 585
R180 B.n262 B.n151 585
R181 B.n258 B.n151 585
R182 B.n264 B.n263 585
R183 B.n265 B.n264 585
R184 B.n146 B.n145 585
R185 B.n147 B.n146 585
R186 B.n273 B.n272 585
R187 B.n272 B.n271 585
R188 B.n274 B.n144 585
R189 B.n144 B.n143 585
R190 B.n276 B.n275 585
R191 B.n277 B.n276 585
R192 B.n138 B.n137 585
R193 B.n139 B.n138 585
R194 B.n285 B.n284 585
R195 B.n284 B.n283 585
R196 B.n286 B.n136 585
R197 B.n136 B.n135 585
R198 B.n288 B.n287 585
R199 B.n289 B.n288 585
R200 B.n130 B.n129 585
R201 B.n131 B.n130 585
R202 B.n297 B.n296 585
R203 B.n296 B.n295 585
R204 B.n298 B.n128 585
R205 B.n128 B.n127 585
R206 B.n300 B.n299 585
R207 B.n301 B.n300 585
R208 B.n122 B.n121 585
R209 B.n123 B.n122 585
R210 B.n310 B.n309 585
R211 B.n309 B.n308 585
R212 B.n311 B.n120 585
R213 B.n120 B.n119 585
R214 B.n313 B.n312 585
R215 B.n314 B.n313 585
R216 B.n3 B.n0 585
R217 B.n4 B.n3 585
R218 B.n411 B.n1 585
R219 B.n412 B.n411 585
R220 B.n410 B.n409 585
R221 B.n410 B.n8 585
R222 B.n408 B.n9 585
R223 B.n12 B.n9 585
R224 B.n407 B.n406 585
R225 B.n406 B.n405 585
R226 B.n11 B.n10 585
R227 B.n404 B.n11 585
R228 B.n402 B.n401 585
R229 B.n403 B.n402 585
R230 B.n400 B.n17 585
R231 B.n17 B.n16 585
R232 B.n399 B.n398 585
R233 B.n398 B.n397 585
R234 B.n19 B.n18 585
R235 B.n396 B.n19 585
R236 B.n394 B.n393 585
R237 B.n395 B.n394 585
R238 B.n392 B.n24 585
R239 B.n24 B.n23 585
R240 B.n391 B.n390 585
R241 B.n390 B.n389 585
R242 B.n26 B.n25 585
R243 B.n388 B.n26 585
R244 B.n386 B.n385 585
R245 B.n387 B.n386 585
R246 B.n384 B.n31 585
R247 B.n31 B.n30 585
R248 B.n383 B.n382 585
R249 B.n382 B.n381 585
R250 B.n33 B.n32 585
R251 B.n380 B.n33 585
R252 B.n378 B.n377 585
R253 B.n379 B.n378 585
R254 B.n376 B.n37 585
R255 B.n40 B.n37 585
R256 B.n375 B.n374 585
R257 B.n374 B.n373 585
R258 B.n39 B.n38 585
R259 B.n372 B.n39 585
R260 B.n370 B.n369 585
R261 B.n371 B.n370 585
R262 B.n368 B.n45 585
R263 B.n45 B.n44 585
R264 B.n367 B.n366 585
R265 B.n366 B.n365 585
R266 B.n47 B.n46 585
R267 B.n364 B.n47 585
R268 B.n362 B.n361 585
R269 B.n363 B.n362 585
R270 B.n360 B.n52 585
R271 B.n52 B.n51 585
R272 B.n415 B.n414 585
R273 B.n413 B.n2 585
R274 B.n358 B.n52 526.135
R275 B.n355 B.n67 526.135
R276 B.n187 B.n165 526.135
R277 B.n235 B.n167 526.135
R278 B.n70 B.t14 306.86
R279 B.n68 B.t4 306.86
R280 B.n184 B.t9 306.86
R281 B.n182 B.t12 306.86
R282 B.n356 B.n65 256.663
R283 B.n356 B.n64 256.663
R284 B.n356 B.n63 256.663
R285 B.n356 B.n62 256.663
R286 B.n356 B.n61 256.663
R287 B.n356 B.n60 256.663
R288 B.n356 B.n59 256.663
R289 B.n356 B.n58 256.663
R290 B.n356 B.n57 256.663
R291 B.n356 B.n56 256.663
R292 B.n356 B.n55 256.663
R293 B.n357 B.n356 256.663
R294 B.n234 B.n233 256.663
R295 B.n233 B.n170 256.663
R296 B.n233 B.n171 256.663
R297 B.n233 B.n172 256.663
R298 B.n233 B.n173 256.663
R299 B.n233 B.n174 256.663
R300 B.n233 B.n175 256.663
R301 B.n233 B.n176 256.663
R302 B.n233 B.n177 256.663
R303 B.n233 B.n178 256.663
R304 B.n233 B.n179 256.663
R305 B.n233 B.n180 256.663
R306 B.n417 B.n416 256.663
R307 B.n71 B.t15 242.859
R308 B.n69 B.t5 242.859
R309 B.n185 B.t8 242.859
R310 B.n183 B.t11 242.859
R311 B.n233 B.n166 237.274
R312 B.n356 B.n51 237.274
R313 B.n70 B.t13 209.84
R314 B.n68 B.t2 209.84
R315 B.n184 B.t6 209.84
R316 B.n182 B.t10 209.84
R317 B.n73 B.n54 163.367
R318 B.n77 B.n76 163.367
R319 B.n81 B.n80 163.367
R320 B.n85 B.n84 163.367
R321 B.n89 B.n88 163.367
R322 B.n93 B.n92 163.367
R323 B.n97 B.n96 163.367
R324 B.n101 B.n100 163.367
R325 B.n106 B.n105 163.367
R326 B.n110 B.n109 163.367
R327 B.n114 B.n113 163.367
R328 B.n355 B.n66 163.367
R329 B.n241 B.n165 163.367
R330 B.n241 B.n163 163.367
R331 B.n245 B.n163 163.367
R332 B.n245 B.n157 163.367
R333 B.n253 B.n157 163.367
R334 B.n253 B.n155 163.367
R335 B.n257 B.n155 163.367
R336 B.n257 B.n150 163.367
R337 B.n266 B.n150 163.367
R338 B.n266 B.n148 163.367
R339 B.n270 B.n148 163.367
R340 B.n270 B.n142 163.367
R341 B.n278 B.n142 163.367
R342 B.n278 B.n140 163.367
R343 B.n282 B.n140 163.367
R344 B.n282 B.n134 163.367
R345 B.n290 B.n134 163.367
R346 B.n290 B.n132 163.367
R347 B.n294 B.n132 163.367
R348 B.n294 B.n126 163.367
R349 B.n302 B.n126 163.367
R350 B.n302 B.n124 163.367
R351 B.n307 B.n124 163.367
R352 B.n307 B.n118 163.367
R353 B.n315 B.n118 163.367
R354 B.n316 B.n315 163.367
R355 B.n316 B.n5 163.367
R356 B.n6 B.n5 163.367
R357 B.n7 B.n6 163.367
R358 B.n322 B.n7 163.367
R359 B.n323 B.n322 163.367
R360 B.n323 B.n13 163.367
R361 B.n14 B.n13 163.367
R362 B.n15 B.n14 163.367
R363 B.n328 B.n15 163.367
R364 B.n328 B.n20 163.367
R365 B.n21 B.n20 163.367
R366 B.n22 B.n21 163.367
R367 B.n333 B.n22 163.367
R368 B.n333 B.n27 163.367
R369 B.n28 B.n27 163.367
R370 B.n29 B.n28 163.367
R371 B.n338 B.n29 163.367
R372 B.n338 B.n34 163.367
R373 B.n35 B.n34 163.367
R374 B.n36 B.n35 163.367
R375 B.n343 B.n36 163.367
R376 B.n343 B.n41 163.367
R377 B.n42 B.n41 163.367
R378 B.n43 B.n42 163.367
R379 B.n348 B.n43 163.367
R380 B.n348 B.n48 163.367
R381 B.n49 B.n48 163.367
R382 B.n50 B.n49 163.367
R383 B.n67 B.n50 163.367
R384 B.n232 B.n169 163.367
R385 B.n232 B.n181 163.367
R386 B.n228 B.n227 163.367
R387 B.n224 B.n223 163.367
R388 B.n219 B.n218 163.367
R389 B.n215 B.n214 163.367
R390 B.n211 B.n210 163.367
R391 B.n207 B.n206 163.367
R392 B.n203 B.n202 163.367
R393 B.n199 B.n198 163.367
R394 B.n195 B.n194 163.367
R395 B.n191 B.n190 163.367
R396 B.n239 B.n167 163.367
R397 B.n239 B.n161 163.367
R398 B.n247 B.n161 163.367
R399 B.n247 B.n159 163.367
R400 B.n251 B.n159 163.367
R401 B.n251 B.n153 163.367
R402 B.n260 B.n153 163.367
R403 B.n260 B.n151 163.367
R404 B.n264 B.n151 163.367
R405 B.n264 B.n146 163.367
R406 B.n272 B.n146 163.367
R407 B.n272 B.n144 163.367
R408 B.n276 B.n144 163.367
R409 B.n276 B.n138 163.367
R410 B.n284 B.n138 163.367
R411 B.n284 B.n136 163.367
R412 B.n288 B.n136 163.367
R413 B.n288 B.n130 163.367
R414 B.n296 B.n130 163.367
R415 B.n296 B.n128 163.367
R416 B.n300 B.n128 163.367
R417 B.n300 B.n122 163.367
R418 B.n309 B.n122 163.367
R419 B.n309 B.n120 163.367
R420 B.n313 B.n120 163.367
R421 B.n313 B.n3 163.367
R422 B.n415 B.n3 163.367
R423 B.n411 B.n2 163.367
R424 B.n411 B.n410 163.367
R425 B.n410 B.n9 163.367
R426 B.n406 B.n9 163.367
R427 B.n406 B.n11 163.367
R428 B.n402 B.n11 163.367
R429 B.n402 B.n17 163.367
R430 B.n398 B.n17 163.367
R431 B.n398 B.n19 163.367
R432 B.n394 B.n19 163.367
R433 B.n394 B.n24 163.367
R434 B.n390 B.n24 163.367
R435 B.n390 B.n26 163.367
R436 B.n386 B.n26 163.367
R437 B.n386 B.n31 163.367
R438 B.n382 B.n31 163.367
R439 B.n382 B.n33 163.367
R440 B.n378 B.n33 163.367
R441 B.n378 B.n37 163.367
R442 B.n374 B.n37 163.367
R443 B.n374 B.n39 163.367
R444 B.n370 B.n39 163.367
R445 B.n370 B.n45 163.367
R446 B.n366 B.n45 163.367
R447 B.n366 B.n47 163.367
R448 B.n362 B.n47 163.367
R449 B.n362 B.n52 163.367
R450 B.n240 B.n166 129.077
R451 B.n240 B.n162 129.077
R452 B.n246 B.n162 129.077
R453 B.n246 B.n158 129.077
R454 B.n252 B.n158 129.077
R455 B.n252 B.n154 129.077
R456 B.n259 B.n154 129.077
R457 B.n259 B.n258 129.077
R458 B.n265 B.n147 129.077
R459 B.n271 B.n147 129.077
R460 B.n271 B.n143 129.077
R461 B.n277 B.n143 129.077
R462 B.n277 B.n139 129.077
R463 B.n283 B.n139 129.077
R464 B.n283 B.n135 129.077
R465 B.n289 B.n135 129.077
R466 B.n289 B.n131 129.077
R467 B.n295 B.n131 129.077
R468 B.n295 B.n127 129.077
R469 B.n301 B.n127 129.077
R470 B.n308 B.n123 129.077
R471 B.n308 B.n119 129.077
R472 B.n314 B.n119 129.077
R473 B.n314 B.n4 129.077
R474 B.n414 B.n4 129.077
R475 B.n414 B.n413 129.077
R476 B.n413 B.n412 129.077
R477 B.n412 B.n8 129.077
R478 B.n12 B.n8 129.077
R479 B.n405 B.n12 129.077
R480 B.n405 B.n404 129.077
R481 B.n403 B.n16 129.077
R482 B.n397 B.n16 129.077
R483 B.n397 B.n396 129.077
R484 B.n396 B.n395 129.077
R485 B.n395 B.n23 129.077
R486 B.n389 B.n23 129.077
R487 B.n389 B.n388 129.077
R488 B.n388 B.n387 129.077
R489 B.n387 B.n30 129.077
R490 B.n381 B.n30 129.077
R491 B.n381 B.n380 129.077
R492 B.n380 B.n379 129.077
R493 B.n373 B.n40 129.077
R494 B.n373 B.n372 129.077
R495 B.n372 B.n371 129.077
R496 B.n371 B.n44 129.077
R497 B.n365 B.n44 129.077
R498 B.n365 B.n364 129.077
R499 B.n364 B.n363 129.077
R500 B.n363 B.n51 129.077
R501 B.t0 B.n123 123.382
R502 B.n404 B.t1 123.382
R503 B.n265 B.t7 111.993
R504 B.n379 B.t3 111.993
R505 B.n358 B.n357 71.676
R506 B.n73 B.n55 71.676
R507 B.n77 B.n56 71.676
R508 B.n81 B.n57 71.676
R509 B.n85 B.n58 71.676
R510 B.n89 B.n59 71.676
R511 B.n93 B.n60 71.676
R512 B.n97 B.n61 71.676
R513 B.n101 B.n62 71.676
R514 B.n106 B.n63 71.676
R515 B.n110 B.n64 71.676
R516 B.n114 B.n65 71.676
R517 B.n66 B.n65 71.676
R518 B.n113 B.n64 71.676
R519 B.n109 B.n63 71.676
R520 B.n105 B.n62 71.676
R521 B.n100 B.n61 71.676
R522 B.n96 B.n60 71.676
R523 B.n92 B.n59 71.676
R524 B.n88 B.n58 71.676
R525 B.n84 B.n57 71.676
R526 B.n80 B.n56 71.676
R527 B.n76 B.n55 71.676
R528 B.n357 B.n54 71.676
R529 B.n235 B.n234 71.676
R530 B.n181 B.n170 71.676
R531 B.n227 B.n171 71.676
R532 B.n223 B.n172 71.676
R533 B.n218 B.n173 71.676
R534 B.n214 B.n174 71.676
R535 B.n210 B.n175 71.676
R536 B.n206 B.n176 71.676
R537 B.n202 B.n177 71.676
R538 B.n198 B.n178 71.676
R539 B.n194 B.n179 71.676
R540 B.n190 B.n180 71.676
R541 B.n234 B.n169 71.676
R542 B.n228 B.n170 71.676
R543 B.n224 B.n171 71.676
R544 B.n219 B.n172 71.676
R545 B.n215 B.n173 71.676
R546 B.n211 B.n174 71.676
R547 B.n207 B.n175 71.676
R548 B.n203 B.n176 71.676
R549 B.n199 B.n177 71.676
R550 B.n195 B.n178 71.676
R551 B.n191 B.n179 71.676
R552 B.n187 B.n180 71.676
R553 B.n416 B.n415 71.676
R554 B.n416 B.n2 71.676
R555 B.n71 B.n70 64.0005
R556 B.n69 B.n68 64.0005
R557 B.n185 B.n184 64.0005
R558 B.n183 B.n182 64.0005
R559 B.n72 B.n71 59.5399
R560 B.n103 B.n69 59.5399
R561 B.n186 B.n185 59.5399
R562 B.n221 B.n183 59.5399
R563 B.n237 B.n236 34.1859
R564 B.n188 B.n164 34.1859
R565 B.n354 B.n353 34.1859
R566 B.n360 B.n359 34.1859
R567 B B.n417 18.0485
R568 B.n258 B.t7 17.0842
R569 B.n40 B.t3 17.0842
R570 B.n238 B.n237 10.6151
R571 B.n238 B.n160 10.6151
R572 B.n248 B.n160 10.6151
R573 B.n249 B.n248 10.6151
R574 B.n250 B.n249 10.6151
R575 B.n250 B.n152 10.6151
R576 B.n261 B.n152 10.6151
R577 B.n262 B.n261 10.6151
R578 B.n263 B.n262 10.6151
R579 B.n263 B.n145 10.6151
R580 B.n273 B.n145 10.6151
R581 B.n274 B.n273 10.6151
R582 B.n275 B.n274 10.6151
R583 B.n275 B.n137 10.6151
R584 B.n285 B.n137 10.6151
R585 B.n286 B.n285 10.6151
R586 B.n287 B.n286 10.6151
R587 B.n287 B.n129 10.6151
R588 B.n297 B.n129 10.6151
R589 B.n298 B.n297 10.6151
R590 B.n299 B.n298 10.6151
R591 B.n299 B.n121 10.6151
R592 B.n310 B.n121 10.6151
R593 B.n311 B.n310 10.6151
R594 B.n312 B.n311 10.6151
R595 B.n312 B.n0 10.6151
R596 B.n236 B.n168 10.6151
R597 B.n231 B.n168 10.6151
R598 B.n231 B.n230 10.6151
R599 B.n230 B.n229 10.6151
R600 B.n229 B.n226 10.6151
R601 B.n226 B.n225 10.6151
R602 B.n225 B.n222 10.6151
R603 B.n220 B.n217 10.6151
R604 B.n217 B.n216 10.6151
R605 B.n216 B.n213 10.6151
R606 B.n213 B.n212 10.6151
R607 B.n212 B.n209 10.6151
R608 B.n209 B.n208 10.6151
R609 B.n208 B.n205 10.6151
R610 B.n205 B.n204 10.6151
R611 B.n201 B.n200 10.6151
R612 B.n200 B.n197 10.6151
R613 B.n197 B.n196 10.6151
R614 B.n196 B.n193 10.6151
R615 B.n193 B.n192 10.6151
R616 B.n192 B.n189 10.6151
R617 B.n189 B.n188 10.6151
R618 B.n242 B.n164 10.6151
R619 B.n243 B.n242 10.6151
R620 B.n244 B.n243 10.6151
R621 B.n244 B.n156 10.6151
R622 B.n254 B.n156 10.6151
R623 B.n255 B.n254 10.6151
R624 B.n256 B.n255 10.6151
R625 B.n256 B.n149 10.6151
R626 B.n267 B.n149 10.6151
R627 B.n268 B.n267 10.6151
R628 B.n269 B.n268 10.6151
R629 B.n269 B.n141 10.6151
R630 B.n279 B.n141 10.6151
R631 B.n280 B.n279 10.6151
R632 B.n281 B.n280 10.6151
R633 B.n281 B.n133 10.6151
R634 B.n291 B.n133 10.6151
R635 B.n292 B.n291 10.6151
R636 B.n293 B.n292 10.6151
R637 B.n293 B.n125 10.6151
R638 B.n303 B.n125 10.6151
R639 B.n304 B.n303 10.6151
R640 B.n306 B.n304 10.6151
R641 B.n306 B.n305 10.6151
R642 B.n305 B.n117 10.6151
R643 B.n317 B.n117 10.6151
R644 B.n318 B.n317 10.6151
R645 B.n319 B.n318 10.6151
R646 B.n320 B.n319 10.6151
R647 B.n321 B.n320 10.6151
R648 B.n324 B.n321 10.6151
R649 B.n325 B.n324 10.6151
R650 B.n326 B.n325 10.6151
R651 B.n327 B.n326 10.6151
R652 B.n329 B.n327 10.6151
R653 B.n330 B.n329 10.6151
R654 B.n331 B.n330 10.6151
R655 B.n332 B.n331 10.6151
R656 B.n334 B.n332 10.6151
R657 B.n335 B.n334 10.6151
R658 B.n336 B.n335 10.6151
R659 B.n337 B.n336 10.6151
R660 B.n339 B.n337 10.6151
R661 B.n340 B.n339 10.6151
R662 B.n341 B.n340 10.6151
R663 B.n342 B.n341 10.6151
R664 B.n344 B.n342 10.6151
R665 B.n345 B.n344 10.6151
R666 B.n346 B.n345 10.6151
R667 B.n347 B.n346 10.6151
R668 B.n349 B.n347 10.6151
R669 B.n350 B.n349 10.6151
R670 B.n351 B.n350 10.6151
R671 B.n352 B.n351 10.6151
R672 B.n353 B.n352 10.6151
R673 B.n409 B.n1 10.6151
R674 B.n409 B.n408 10.6151
R675 B.n408 B.n407 10.6151
R676 B.n407 B.n10 10.6151
R677 B.n401 B.n10 10.6151
R678 B.n401 B.n400 10.6151
R679 B.n400 B.n399 10.6151
R680 B.n399 B.n18 10.6151
R681 B.n393 B.n18 10.6151
R682 B.n393 B.n392 10.6151
R683 B.n392 B.n391 10.6151
R684 B.n391 B.n25 10.6151
R685 B.n385 B.n25 10.6151
R686 B.n385 B.n384 10.6151
R687 B.n384 B.n383 10.6151
R688 B.n383 B.n32 10.6151
R689 B.n377 B.n32 10.6151
R690 B.n377 B.n376 10.6151
R691 B.n376 B.n375 10.6151
R692 B.n375 B.n38 10.6151
R693 B.n369 B.n38 10.6151
R694 B.n369 B.n368 10.6151
R695 B.n368 B.n367 10.6151
R696 B.n367 B.n46 10.6151
R697 B.n361 B.n46 10.6151
R698 B.n361 B.n360 10.6151
R699 B.n359 B.n53 10.6151
R700 B.n74 B.n53 10.6151
R701 B.n75 B.n74 10.6151
R702 B.n78 B.n75 10.6151
R703 B.n79 B.n78 10.6151
R704 B.n82 B.n79 10.6151
R705 B.n83 B.n82 10.6151
R706 B.n87 B.n86 10.6151
R707 B.n90 B.n87 10.6151
R708 B.n91 B.n90 10.6151
R709 B.n94 B.n91 10.6151
R710 B.n95 B.n94 10.6151
R711 B.n98 B.n95 10.6151
R712 B.n99 B.n98 10.6151
R713 B.n102 B.n99 10.6151
R714 B.n107 B.n104 10.6151
R715 B.n108 B.n107 10.6151
R716 B.n111 B.n108 10.6151
R717 B.n112 B.n111 10.6151
R718 B.n115 B.n112 10.6151
R719 B.n116 B.n115 10.6151
R720 B.n354 B.n116 10.6151
R721 B.n417 B.n0 8.11757
R722 B.n417 B.n1 8.11757
R723 B.n221 B.n220 6.5566
R724 B.n204 B.n186 6.5566
R725 B.n86 B.n72 6.5566
R726 B.n103 B.n102 6.5566
R727 B.n301 B.t0 5.69506
R728 B.t1 B.n403 5.69506
R729 B.n222 B.n221 4.05904
R730 B.n201 B.n186 4.05904
R731 B.n83 B.n72 4.05904
R732 B.n104 B.n103 4.05904
R733 VN VN.t1 82.3005
R734 VN VN.t0 45.7891
R735 VTAIL.n3 VTAIL.t3 253.71
R736 VTAIL.n0 VTAIL.t0 253.71
R737 VTAIL.n2 VTAIL.t1 253.71
R738 VTAIL.n1 VTAIL.t2 253.71
R739 VTAIL.n1 VTAIL.n0 18.5048
R740 VTAIL.n3 VTAIL.n2 15.66
R741 VTAIL.n2 VTAIL.n1 1.89274
R742 VTAIL VTAIL.n0 1.23972
R743 VTAIL VTAIL.n3 0.653517
R744 VDD2.n0 VDD2.t1 300.187
R745 VDD2.n0 VDD2.t0 270.389
R746 VDD2 VDD2.n0 0.769897
R747 VP.n0 VP.t1 82.2988
R748 VP.n0 VP.t0 45.3578
R749 VP VP.n0 0.431812
R750 VDD1 VDD1.t1 301.423
R751 VDD1 VDD1.t0 271.159
C0 VDD2 VTAIL 2.21386f
C1 VDD1 VP 0.572636f
C2 VDD1 VN 0.157121f
C3 VN VP 3.50892f
C4 VDD2 VDD1 0.718378f
C5 VDD2 VP 0.358175f
C6 VDD1 VTAIL 2.15807f
C7 VDD2 VN 0.373839f
C8 VTAIL VP 0.956274f
C9 VTAIL VN 0.942161f
C10 VDD2 B 2.482087f
C11 VDD1 B 4.57974f
C12 VTAIL B 2.364533f
C13 VN B 7.99824f
C14 VP B 5.781623f
C15 VDD1.t0 B 0.040651f
C16 VDD1.t1 B 0.126329f
C17 VP.t0 B 0.36333f
C18 VP.t1 B 0.97818f
C19 VP.n0 B 2.05633f
C20 VDD2.t1 B 0.120814f
C21 VDD2.t0 B 0.04177f
C22 VDD2.n0 B 1.88565f
C23 VTAIL.t0 B 0.051373f
C24 VTAIL.n0 B 1.12001f
C25 VTAIL.t2 B 0.051373f
C26 VTAIL.n1 B 1.1806f
C27 VTAIL.t1 B 0.051373f
C28 VTAIL.n2 B 0.916655f
C29 VTAIL.t3 B 0.051373f
C30 VTAIL.n3 B 0.80168f
C31 VN.t0 B 0.360318f
C32 VN.t1 B 0.96935f
.ends

