* NGSPICE file created from diff_pair_sample_1412.ext - technology: sky130A

.subckt diff_pair_sample_1412 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=0 ps=0 w=15.68 l=2.86
X1 B.t8 B.t6 B.t7 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=0 ps=0 w=15.68 l=2.86
X2 B.t5 B.t3 B.t4 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=0 ps=0 w=15.68 l=2.86
X3 VTAIL.t7 VN.t0 VDD2.t0 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=2.5872 ps=16.01 w=15.68 l=2.86
X4 VDD1.t3 VP.t0 VTAIL.t2 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=2.5872 pd=16.01 as=6.1152 ps=32.14 w=15.68 l=2.86
X5 VDD2.t2 VN.t1 VTAIL.t6 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=2.5872 pd=16.01 as=6.1152 ps=32.14 w=15.68 l=2.86
X6 VTAIL.t5 VN.t2 VDD2.t3 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=2.5872 ps=16.01 w=15.68 l=2.86
X7 VTAIL.t3 VP.t1 VDD1.t2 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=2.5872 ps=16.01 w=15.68 l=2.86
X8 VDD2.t1 VN.t3 VTAIL.t4 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=2.5872 pd=16.01 as=6.1152 ps=32.14 w=15.68 l=2.86
X9 VDD1.t1 VP.t2 VTAIL.t1 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=2.5872 pd=16.01 as=6.1152 ps=32.14 w=15.68 l=2.86
X10 B.t2 B.t0 B.t1 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=0 ps=0 w=15.68 l=2.86
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n2884_n4104# sky130_fd_pr__pfet_01v8 ad=6.1152 pd=32.14 as=2.5872 ps=16.01 w=15.68 l=2.86
R0 B.n532 B.n81 585
R1 B.n534 B.n533 585
R2 B.n535 B.n80 585
R3 B.n537 B.n536 585
R4 B.n538 B.n79 585
R5 B.n540 B.n539 585
R6 B.n541 B.n78 585
R7 B.n543 B.n542 585
R8 B.n544 B.n77 585
R9 B.n546 B.n545 585
R10 B.n547 B.n76 585
R11 B.n549 B.n548 585
R12 B.n550 B.n75 585
R13 B.n552 B.n551 585
R14 B.n553 B.n74 585
R15 B.n555 B.n554 585
R16 B.n556 B.n73 585
R17 B.n558 B.n557 585
R18 B.n559 B.n72 585
R19 B.n561 B.n560 585
R20 B.n562 B.n71 585
R21 B.n564 B.n563 585
R22 B.n565 B.n70 585
R23 B.n567 B.n566 585
R24 B.n568 B.n69 585
R25 B.n570 B.n569 585
R26 B.n571 B.n68 585
R27 B.n573 B.n572 585
R28 B.n574 B.n67 585
R29 B.n576 B.n575 585
R30 B.n577 B.n66 585
R31 B.n579 B.n578 585
R32 B.n580 B.n65 585
R33 B.n582 B.n581 585
R34 B.n583 B.n64 585
R35 B.n585 B.n584 585
R36 B.n586 B.n63 585
R37 B.n588 B.n587 585
R38 B.n589 B.n62 585
R39 B.n591 B.n590 585
R40 B.n592 B.n61 585
R41 B.n594 B.n593 585
R42 B.n595 B.n60 585
R43 B.n597 B.n596 585
R44 B.n598 B.n59 585
R45 B.n600 B.n599 585
R46 B.n601 B.n58 585
R47 B.n603 B.n602 585
R48 B.n604 B.n57 585
R49 B.n606 B.n605 585
R50 B.n607 B.n56 585
R51 B.n609 B.n608 585
R52 B.n611 B.n53 585
R53 B.n613 B.n612 585
R54 B.n614 B.n52 585
R55 B.n616 B.n615 585
R56 B.n617 B.n51 585
R57 B.n619 B.n618 585
R58 B.n620 B.n50 585
R59 B.n622 B.n621 585
R60 B.n623 B.n49 585
R61 B.n625 B.n624 585
R62 B.n627 B.n626 585
R63 B.n628 B.n45 585
R64 B.n630 B.n629 585
R65 B.n631 B.n44 585
R66 B.n633 B.n632 585
R67 B.n634 B.n43 585
R68 B.n636 B.n635 585
R69 B.n637 B.n42 585
R70 B.n639 B.n638 585
R71 B.n640 B.n41 585
R72 B.n642 B.n641 585
R73 B.n643 B.n40 585
R74 B.n645 B.n644 585
R75 B.n646 B.n39 585
R76 B.n648 B.n647 585
R77 B.n649 B.n38 585
R78 B.n651 B.n650 585
R79 B.n652 B.n37 585
R80 B.n654 B.n653 585
R81 B.n655 B.n36 585
R82 B.n657 B.n656 585
R83 B.n658 B.n35 585
R84 B.n660 B.n659 585
R85 B.n661 B.n34 585
R86 B.n663 B.n662 585
R87 B.n664 B.n33 585
R88 B.n666 B.n665 585
R89 B.n667 B.n32 585
R90 B.n669 B.n668 585
R91 B.n670 B.n31 585
R92 B.n672 B.n671 585
R93 B.n673 B.n30 585
R94 B.n675 B.n674 585
R95 B.n676 B.n29 585
R96 B.n678 B.n677 585
R97 B.n679 B.n28 585
R98 B.n681 B.n680 585
R99 B.n682 B.n27 585
R100 B.n684 B.n683 585
R101 B.n685 B.n26 585
R102 B.n687 B.n686 585
R103 B.n688 B.n25 585
R104 B.n690 B.n689 585
R105 B.n691 B.n24 585
R106 B.n693 B.n692 585
R107 B.n694 B.n23 585
R108 B.n696 B.n695 585
R109 B.n697 B.n22 585
R110 B.n699 B.n698 585
R111 B.n700 B.n21 585
R112 B.n702 B.n701 585
R113 B.n703 B.n20 585
R114 B.n531 B.n530 585
R115 B.n529 B.n82 585
R116 B.n528 B.n527 585
R117 B.n526 B.n83 585
R118 B.n525 B.n524 585
R119 B.n523 B.n84 585
R120 B.n522 B.n521 585
R121 B.n520 B.n85 585
R122 B.n519 B.n518 585
R123 B.n517 B.n86 585
R124 B.n516 B.n515 585
R125 B.n514 B.n87 585
R126 B.n513 B.n512 585
R127 B.n511 B.n88 585
R128 B.n510 B.n509 585
R129 B.n508 B.n89 585
R130 B.n507 B.n506 585
R131 B.n505 B.n90 585
R132 B.n504 B.n503 585
R133 B.n502 B.n91 585
R134 B.n501 B.n500 585
R135 B.n499 B.n92 585
R136 B.n498 B.n497 585
R137 B.n496 B.n93 585
R138 B.n495 B.n494 585
R139 B.n493 B.n94 585
R140 B.n492 B.n491 585
R141 B.n490 B.n95 585
R142 B.n489 B.n488 585
R143 B.n487 B.n96 585
R144 B.n486 B.n485 585
R145 B.n484 B.n97 585
R146 B.n483 B.n482 585
R147 B.n481 B.n98 585
R148 B.n480 B.n479 585
R149 B.n478 B.n99 585
R150 B.n477 B.n476 585
R151 B.n475 B.n100 585
R152 B.n474 B.n473 585
R153 B.n472 B.n101 585
R154 B.n471 B.n470 585
R155 B.n469 B.n102 585
R156 B.n468 B.n467 585
R157 B.n466 B.n103 585
R158 B.n465 B.n464 585
R159 B.n463 B.n104 585
R160 B.n462 B.n461 585
R161 B.n460 B.n105 585
R162 B.n459 B.n458 585
R163 B.n457 B.n106 585
R164 B.n456 B.n455 585
R165 B.n454 B.n107 585
R166 B.n453 B.n452 585
R167 B.n451 B.n108 585
R168 B.n450 B.n449 585
R169 B.n448 B.n109 585
R170 B.n447 B.n446 585
R171 B.n445 B.n110 585
R172 B.n444 B.n443 585
R173 B.n442 B.n111 585
R174 B.n441 B.n440 585
R175 B.n439 B.n112 585
R176 B.n438 B.n437 585
R177 B.n436 B.n113 585
R178 B.n435 B.n434 585
R179 B.n433 B.n114 585
R180 B.n432 B.n431 585
R181 B.n430 B.n115 585
R182 B.n429 B.n428 585
R183 B.n427 B.n116 585
R184 B.n426 B.n425 585
R185 B.n424 B.n117 585
R186 B.n423 B.n422 585
R187 B.n250 B.n179 585
R188 B.n252 B.n251 585
R189 B.n253 B.n178 585
R190 B.n255 B.n254 585
R191 B.n256 B.n177 585
R192 B.n258 B.n257 585
R193 B.n259 B.n176 585
R194 B.n261 B.n260 585
R195 B.n262 B.n175 585
R196 B.n264 B.n263 585
R197 B.n265 B.n174 585
R198 B.n267 B.n266 585
R199 B.n268 B.n173 585
R200 B.n270 B.n269 585
R201 B.n271 B.n172 585
R202 B.n273 B.n272 585
R203 B.n274 B.n171 585
R204 B.n276 B.n275 585
R205 B.n277 B.n170 585
R206 B.n279 B.n278 585
R207 B.n280 B.n169 585
R208 B.n282 B.n281 585
R209 B.n283 B.n168 585
R210 B.n285 B.n284 585
R211 B.n286 B.n167 585
R212 B.n288 B.n287 585
R213 B.n289 B.n166 585
R214 B.n291 B.n290 585
R215 B.n292 B.n165 585
R216 B.n294 B.n293 585
R217 B.n295 B.n164 585
R218 B.n297 B.n296 585
R219 B.n298 B.n163 585
R220 B.n300 B.n299 585
R221 B.n301 B.n162 585
R222 B.n303 B.n302 585
R223 B.n304 B.n161 585
R224 B.n306 B.n305 585
R225 B.n307 B.n160 585
R226 B.n309 B.n308 585
R227 B.n310 B.n159 585
R228 B.n312 B.n311 585
R229 B.n313 B.n158 585
R230 B.n315 B.n314 585
R231 B.n316 B.n157 585
R232 B.n318 B.n317 585
R233 B.n319 B.n156 585
R234 B.n321 B.n320 585
R235 B.n322 B.n155 585
R236 B.n324 B.n323 585
R237 B.n325 B.n154 585
R238 B.n327 B.n326 585
R239 B.n329 B.n151 585
R240 B.n331 B.n330 585
R241 B.n332 B.n150 585
R242 B.n334 B.n333 585
R243 B.n335 B.n149 585
R244 B.n337 B.n336 585
R245 B.n338 B.n148 585
R246 B.n340 B.n339 585
R247 B.n341 B.n147 585
R248 B.n343 B.n342 585
R249 B.n345 B.n344 585
R250 B.n346 B.n143 585
R251 B.n348 B.n347 585
R252 B.n349 B.n142 585
R253 B.n351 B.n350 585
R254 B.n352 B.n141 585
R255 B.n354 B.n353 585
R256 B.n355 B.n140 585
R257 B.n357 B.n356 585
R258 B.n358 B.n139 585
R259 B.n360 B.n359 585
R260 B.n361 B.n138 585
R261 B.n363 B.n362 585
R262 B.n364 B.n137 585
R263 B.n366 B.n365 585
R264 B.n367 B.n136 585
R265 B.n369 B.n368 585
R266 B.n370 B.n135 585
R267 B.n372 B.n371 585
R268 B.n373 B.n134 585
R269 B.n375 B.n374 585
R270 B.n376 B.n133 585
R271 B.n378 B.n377 585
R272 B.n379 B.n132 585
R273 B.n381 B.n380 585
R274 B.n382 B.n131 585
R275 B.n384 B.n383 585
R276 B.n385 B.n130 585
R277 B.n387 B.n386 585
R278 B.n388 B.n129 585
R279 B.n390 B.n389 585
R280 B.n391 B.n128 585
R281 B.n393 B.n392 585
R282 B.n394 B.n127 585
R283 B.n396 B.n395 585
R284 B.n397 B.n126 585
R285 B.n399 B.n398 585
R286 B.n400 B.n125 585
R287 B.n402 B.n401 585
R288 B.n403 B.n124 585
R289 B.n405 B.n404 585
R290 B.n406 B.n123 585
R291 B.n408 B.n407 585
R292 B.n409 B.n122 585
R293 B.n411 B.n410 585
R294 B.n412 B.n121 585
R295 B.n414 B.n413 585
R296 B.n415 B.n120 585
R297 B.n417 B.n416 585
R298 B.n418 B.n119 585
R299 B.n420 B.n419 585
R300 B.n421 B.n118 585
R301 B.n249 B.n248 585
R302 B.n247 B.n180 585
R303 B.n246 B.n245 585
R304 B.n244 B.n181 585
R305 B.n243 B.n242 585
R306 B.n241 B.n182 585
R307 B.n240 B.n239 585
R308 B.n238 B.n183 585
R309 B.n237 B.n236 585
R310 B.n235 B.n184 585
R311 B.n234 B.n233 585
R312 B.n232 B.n185 585
R313 B.n231 B.n230 585
R314 B.n229 B.n186 585
R315 B.n228 B.n227 585
R316 B.n226 B.n187 585
R317 B.n225 B.n224 585
R318 B.n223 B.n188 585
R319 B.n222 B.n221 585
R320 B.n220 B.n189 585
R321 B.n219 B.n218 585
R322 B.n217 B.n190 585
R323 B.n216 B.n215 585
R324 B.n214 B.n191 585
R325 B.n213 B.n212 585
R326 B.n211 B.n192 585
R327 B.n210 B.n209 585
R328 B.n208 B.n193 585
R329 B.n207 B.n206 585
R330 B.n205 B.n194 585
R331 B.n204 B.n203 585
R332 B.n202 B.n195 585
R333 B.n201 B.n200 585
R334 B.n199 B.n196 585
R335 B.n198 B.n197 585
R336 B.n2 B.n0 585
R337 B.n757 B.n1 585
R338 B.n756 B.n755 585
R339 B.n754 B.n3 585
R340 B.n753 B.n752 585
R341 B.n751 B.n4 585
R342 B.n750 B.n749 585
R343 B.n748 B.n5 585
R344 B.n747 B.n746 585
R345 B.n745 B.n6 585
R346 B.n744 B.n743 585
R347 B.n742 B.n7 585
R348 B.n741 B.n740 585
R349 B.n739 B.n8 585
R350 B.n738 B.n737 585
R351 B.n736 B.n9 585
R352 B.n735 B.n734 585
R353 B.n733 B.n10 585
R354 B.n732 B.n731 585
R355 B.n730 B.n11 585
R356 B.n729 B.n728 585
R357 B.n727 B.n12 585
R358 B.n726 B.n725 585
R359 B.n724 B.n13 585
R360 B.n723 B.n722 585
R361 B.n721 B.n14 585
R362 B.n720 B.n719 585
R363 B.n718 B.n15 585
R364 B.n717 B.n716 585
R365 B.n715 B.n16 585
R366 B.n714 B.n713 585
R367 B.n712 B.n17 585
R368 B.n711 B.n710 585
R369 B.n709 B.n18 585
R370 B.n708 B.n707 585
R371 B.n706 B.n19 585
R372 B.n705 B.n704 585
R373 B.n759 B.n758 585
R374 B.n248 B.n179 578.989
R375 B.n704 B.n703 578.989
R376 B.n422 B.n421 578.989
R377 B.n530 B.n81 578.989
R378 B.n144 B.t3 340.538
R379 B.n152 B.t9 340.538
R380 B.n46 B.t0 340.538
R381 B.n54 B.t6 340.538
R382 B.n144 B.t5 169.111
R383 B.n54 B.t7 169.111
R384 B.n152 B.t11 169.09
R385 B.n46 B.t1 169.09
R386 B.n248 B.n247 163.367
R387 B.n247 B.n246 163.367
R388 B.n246 B.n181 163.367
R389 B.n242 B.n181 163.367
R390 B.n242 B.n241 163.367
R391 B.n241 B.n240 163.367
R392 B.n240 B.n183 163.367
R393 B.n236 B.n183 163.367
R394 B.n236 B.n235 163.367
R395 B.n235 B.n234 163.367
R396 B.n234 B.n185 163.367
R397 B.n230 B.n185 163.367
R398 B.n230 B.n229 163.367
R399 B.n229 B.n228 163.367
R400 B.n228 B.n187 163.367
R401 B.n224 B.n187 163.367
R402 B.n224 B.n223 163.367
R403 B.n223 B.n222 163.367
R404 B.n222 B.n189 163.367
R405 B.n218 B.n189 163.367
R406 B.n218 B.n217 163.367
R407 B.n217 B.n216 163.367
R408 B.n216 B.n191 163.367
R409 B.n212 B.n191 163.367
R410 B.n212 B.n211 163.367
R411 B.n211 B.n210 163.367
R412 B.n210 B.n193 163.367
R413 B.n206 B.n193 163.367
R414 B.n206 B.n205 163.367
R415 B.n205 B.n204 163.367
R416 B.n204 B.n195 163.367
R417 B.n200 B.n195 163.367
R418 B.n200 B.n199 163.367
R419 B.n199 B.n198 163.367
R420 B.n198 B.n2 163.367
R421 B.n758 B.n2 163.367
R422 B.n758 B.n757 163.367
R423 B.n757 B.n756 163.367
R424 B.n756 B.n3 163.367
R425 B.n752 B.n3 163.367
R426 B.n752 B.n751 163.367
R427 B.n751 B.n750 163.367
R428 B.n750 B.n5 163.367
R429 B.n746 B.n5 163.367
R430 B.n746 B.n745 163.367
R431 B.n745 B.n744 163.367
R432 B.n744 B.n7 163.367
R433 B.n740 B.n7 163.367
R434 B.n740 B.n739 163.367
R435 B.n739 B.n738 163.367
R436 B.n738 B.n9 163.367
R437 B.n734 B.n9 163.367
R438 B.n734 B.n733 163.367
R439 B.n733 B.n732 163.367
R440 B.n732 B.n11 163.367
R441 B.n728 B.n11 163.367
R442 B.n728 B.n727 163.367
R443 B.n727 B.n726 163.367
R444 B.n726 B.n13 163.367
R445 B.n722 B.n13 163.367
R446 B.n722 B.n721 163.367
R447 B.n721 B.n720 163.367
R448 B.n720 B.n15 163.367
R449 B.n716 B.n15 163.367
R450 B.n716 B.n715 163.367
R451 B.n715 B.n714 163.367
R452 B.n714 B.n17 163.367
R453 B.n710 B.n17 163.367
R454 B.n710 B.n709 163.367
R455 B.n709 B.n708 163.367
R456 B.n708 B.n19 163.367
R457 B.n704 B.n19 163.367
R458 B.n252 B.n179 163.367
R459 B.n253 B.n252 163.367
R460 B.n254 B.n253 163.367
R461 B.n254 B.n177 163.367
R462 B.n258 B.n177 163.367
R463 B.n259 B.n258 163.367
R464 B.n260 B.n259 163.367
R465 B.n260 B.n175 163.367
R466 B.n264 B.n175 163.367
R467 B.n265 B.n264 163.367
R468 B.n266 B.n265 163.367
R469 B.n266 B.n173 163.367
R470 B.n270 B.n173 163.367
R471 B.n271 B.n270 163.367
R472 B.n272 B.n271 163.367
R473 B.n272 B.n171 163.367
R474 B.n276 B.n171 163.367
R475 B.n277 B.n276 163.367
R476 B.n278 B.n277 163.367
R477 B.n278 B.n169 163.367
R478 B.n282 B.n169 163.367
R479 B.n283 B.n282 163.367
R480 B.n284 B.n283 163.367
R481 B.n284 B.n167 163.367
R482 B.n288 B.n167 163.367
R483 B.n289 B.n288 163.367
R484 B.n290 B.n289 163.367
R485 B.n290 B.n165 163.367
R486 B.n294 B.n165 163.367
R487 B.n295 B.n294 163.367
R488 B.n296 B.n295 163.367
R489 B.n296 B.n163 163.367
R490 B.n300 B.n163 163.367
R491 B.n301 B.n300 163.367
R492 B.n302 B.n301 163.367
R493 B.n302 B.n161 163.367
R494 B.n306 B.n161 163.367
R495 B.n307 B.n306 163.367
R496 B.n308 B.n307 163.367
R497 B.n308 B.n159 163.367
R498 B.n312 B.n159 163.367
R499 B.n313 B.n312 163.367
R500 B.n314 B.n313 163.367
R501 B.n314 B.n157 163.367
R502 B.n318 B.n157 163.367
R503 B.n319 B.n318 163.367
R504 B.n320 B.n319 163.367
R505 B.n320 B.n155 163.367
R506 B.n324 B.n155 163.367
R507 B.n325 B.n324 163.367
R508 B.n326 B.n325 163.367
R509 B.n326 B.n151 163.367
R510 B.n331 B.n151 163.367
R511 B.n332 B.n331 163.367
R512 B.n333 B.n332 163.367
R513 B.n333 B.n149 163.367
R514 B.n337 B.n149 163.367
R515 B.n338 B.n337 163.367
R516 B.n339 B.n338 163.367
R517 B.n339 B.n147 163.367
R518 B.n343 B.n147 163.367
R519 B.n344 B.n343 163.367
R520 B.n344 B.n143 163.367
R521 B.n348 B.n143 163.367
R522 B.n349 B.n348 163.367
R523 B.n350 B.n349 163.367
R524 B.n350 B.n141 163.367
R525 B.n354 B.n141 163.367
R526 B.n355 B.n354 163.367
R527 B.n356 B.n355 163.367
R528 B.n356 B.n139 163.367
R529 B.n360 B.n139 163.367
R530 B.n361 B.n360 163.367
R531 B.n362 B.n361 163.367
R532 B.n362 B.n137 163.367
R533 B.n366 B.n137 163.367
R534 B.n367 B.n366 163.367
R535 B.n368 B.n367 163.367
R536 B.n368 B.n135 163.367
R537 B.n372 B.n135 163.367
R538 B.n373 B.n372 163.367
R539 B.n374 B.n373 163.367
R540 B.n374 B.n133 163.367
R541 B.n378 B.n133 163.367
R542 B.n379 B.n378 163.367
R543 B.n380 B.n379 163.367
R544 B.n380 B.n131 163.367
R545 B.n384 B.n131 163.367
R546 B.n385 B.n384 163.367
R547 B.n386 B.n385 163.367
R548 B.n386 B.n129 163.367
R549 B.n390 B.n129 163.367
R550 B.n391 B.n390 163.367
R551 B.n392 B.n391 163.367
R552 B.n392 B.n127 163.367
R553 B.n396 B.n127 163.367
R554 B.n397 B.n396 163.367
R555 B.n398 B.n397 163.367
R556 B.n398 B.n125 163.367
R557 B.n402 B.n125 163.367
R558 B.n403 B.n402 163.367
R559 B.n404 B.n403 163.367
R560 B.n404 B.n123 163.367
R561 B.n408 B.n123 163.367
R562 B.n409 B.n408 163.367
R563 B.n410 B.n409 163.367
R564 B.n410 B.n121 163.367
R565 B.n414 B.n121 163.367
R566 B.n415 B.n414 163.367
R567 B.n416 B.n415 163.367
R568 B.n416 B.n119 163.367
R569 B.n420 B.n119 163.367
R570 B.n421 B.n420 163.367
R571 B.n422 B.n117 163.367
R572 B.n426 B.n117 163.367
R573 B.n427 B.n426 163.367
R574 B.n428 B.n427 163.367
R575 B.n428 B.n115 163.367
R576 B.n432 B.n115 163.367
R577 B.n433 B.n432 163.367
R578 B.n434 B.n433 163.367
R579 B.n434 B.n113 163.367
R580 B.n438 B.n113 163.367
R581 B.n439 B.n438 163.367
R582 B.n440 B.n439 163.367
R583 B.n440 B.n111 163.367
R584 B.n444 B.n111 163.367
R585 B.n445 B.n444 163.367
R586 B.n446 B.n445 163.367
R587 B.n446 B.n109 163.367
R588 B.n450 B.n109 163.367
R589 B.n451 B.n450 163.367
R590 B.n452 B.n451 163.367
R591 B.n452 B.n107 163.367
R592 B.n456 B.n107 163.367
R593 B.n457 B.n456 163.367
R594 B.n458 B.n457 163.367
R595 B.n458 B.n105 163.367
R596 B.n462 B.n105 163.367
R597 B.n463 B.n462 163.367
R598 B.n464 B.n463 163.367
R599 B.n464 B.n103 163.367
R600 B.n468 B.n103 163.367
R601 B.n469 B.n468 163.367
R602 B.n470 B.n469 163.367
R603 B.n470 B.n101 163.367
R604 B.n474 B.n101 163.367
R605 B.n475 B.n474 163.367
R606 B.n476 B.n475 163.367
R607 B.n476 B.n99 163.367
R608 B.n480 B.n99 163.367
R609 B.n481 B.n480 163.367
R610 B.n482 B.n481 163.367
R611 B.n482 B.n97 163.367
R612 B.n486 B.n97 163.367
R613 B.n487 B.n486 163.367
R614 B.n488 B.n487 163.367
R615 B.n488 B.n95 163.367
R616 B.n492 B.n95 163.367
R617 B.n493 B.n492 163.367
R618 B.n494 B.n493 163.367
R619 B.n494 B.n93 163.367
R620 B.n498 B.n93 163.367
R621 B.n499 B.n498 163.367
R622 B.n500 B.n499 163.367
R623 B.n500 B.n91 163.367
R624 B.n504 B.n91 163.367
R625 B.n505 B.n504 163.367
R626 B.n506 B.n505 163.367
R627 B.n506 B.n89 163.367
R628 B.n510 B.n89 163.367
R629 B.n511 B.n510 163.367
R630 B.n512 B.n511 163.367
R631 B.n512 B.n87 163.367
R632 B.n516 B.n87 163.367
R633 B.n517 B.n516 163.367
R634 B.n518 B.n517 163.367
R635 B.n518 B.n85 163.367
R636 B.n522 B.n85 163.367
R637 B.n523 B.n522 163.367
R638 B.n524 B.n523 163.367
R639 B.n524 B.n83 163.367
R640 B.n528 B.n83 163.367
R641 B.n529 B.n528 163.367
R642 B.n530 B.n529 163.367
R643 B.n703 B.n702 163.367
R644 B.n702 B.n21 163.367
R645 B.n698 B.n21 163.367
R646 B.n698 B.n697 163.367
R647 B.n697 B.n696 163.367
R648 B.n696 B.n23 163.367
R649 B.n692 B.n23 163.367
R650 B.n692 B.n691 163.367
R651 B.n691 B.n690 163.367
R652 B.n690 B.n25 163.367
R653 B.n686 B.n25 163.367
R654 B.n686 B.n685 163.367
R655 B.n685 B.n684 163.367
R656 B.n684 B.n27 163.367
R657 B.n680 B.n27 163.367
R658 B.n680 B.n679 163.367
R659 B.n679 B.n678 163.367
R660 B.n678 B.n29 163.367
R661 B.n674 B.n29 163.367
R662 B.n674 B.n673 163.367
R663 B.n673 B.n672 163.367
R664 B.n672 B.n31 163.367
R665 B.n668 B.n31 163.367
R666 B.n668 B.n667 163.367
R667 B.n667 B.n666 163.367
R668 B.n666 B.n33 163.367
R669 B.n662 B.n33 163.367
R670 B.n662 B.n661 163.367
R671 B.n661 B.n660 163.367
R672 B.n660 B.n35 163.367
R673 B.n656 B.n35 163.367
R674 B.n656 B.n655 163.367
R675 B.n655 B.n654 163.367
R676 B.n654 B.n37 163.367
R677 B.n650 B.n37 163.367
R678 B.n650 B.n649 163.367
R679 B.n649 B.n648 163.367
R680 B.n648 B.n39 163.367
R681 B.n644 B.n39 163.367
R682 B.n644 B.n643 163.367
R683 B.n643 B.n642 163.367
R684 B.n642 B.n41 163.367
R685 B.n638 B.n41 163.367
R686 B.n638 B.n637 163.367
R687 B.n637 B.n636 163.367
R688 B.n636 B.n43 163.367
R689 B.n632 B.n43 163.367
R690 B.n632 B.n631 163.367
R691 B.n631 B.n630 163.367
R692 B.n630 B.n45 163.367
R693 B.n626 B.n45 163.367
R694 B.n626 B.n625 163.367
R695 B.n625 B.n49 163.367
R696 B.n621 B.n49 163.367
R697 B.n621 B.n620 163.367
R698 B.n620 B.n619 163.367
R699 B.n619 B.n51 163.367
R700 B.n615 B.n51 163.367
R701 B.n615 B.n614 163.367
R702 B.n614 B.n613 163.367
R703 B.n613 B.n53 163.367
R704 B.n608 B.n53 163.367
R705 B.n608 B.n607 163.367
R706 B.n607 B.n606 163.367
R707 B.n606 B.n57 163.367
R708 B.n602 B.n57 163.367
R709 B.n602 B.n601 163.367
R710 B.n601 B.n600 163.367
R711 B.n600 B.n59 163.367
R712 B.n596 B.n59 163.367
R713 B.n596 B.n595 163.367
R714 B.n595 B.n594 163.367
R715 B.n594 B.n61 163.367
R716 B.n590 B.n61 163.367
R717 B.n590 B.n589 163.367
R718 B.n589 B.n588 163.367
R719 B.n588 B.n63 163.367
R720 B.n584 B.n63 163.367
R721 B.n584 B.n583 163.367
R722 B.n583 B.n582 163.367
R723 B.n582 B.n65 163.367
R724 B.n578 B.n65 163.367
R725 B.n578 B.n577 163.367
R726 B.n577 B.n576 163.367
R727 B.n576 B.n67 163.367
R728 B.n572 B.n67 163.367
R729 B.n572 B.n571 163.367
R730 B.n571 B.n570 163.367
R731 B.n570 B.n69 163.367
R732 B.n566 B.n69 163.367
R733 B.n566 B.n565 163.367
R734 B.n565 B.n564 163.367
R735 B.n564 B.n71 163.367
R736 B.n560 B.n71 163.367
R737 B.n560 B.n559 163.367
R738 B.n559 B.n558 163.367
R739 B.n558 B.n73 163.367
R740 B.n554 B.n73 163.367
R741 B.n554 B.n553 163.367
R742 B.n553 B.n552 163.367
R743 B.n552 B.n75 163.367
R744 B.n548 B.n75 163.367
R745 B.n548 B.n547 163.367
R746 B.n547 B.n546 163.367
R747 B.n546 B.n77 163.367
R748 B.n542 B.n77 163.367
R749 B.n542 B.n541 163.367
R750 B.n541 B.n540 163.367
R751 B.n540 B.n79 163.367
R752 B.n536 B.n79 163.367
R753 B.n536 B.n535 163.367
R754 B.n535 B.n534 163.367
R755 B.n534 B.n81 163.367
R756 B.n145 B.t4 107.243
R757 B.n55 B.t8 107.243
R758 B.n153 B.t10 107.224
R759 B.n47 B.t2 107.224
R760 B.n145 B.n144 61.8672
R761 B.n153 B.n152 61.8672
R762 B.n47 B.n46 61.8672
R763 B.n55 B.n54 61.8672
R764 B.n146 B.n145 59.5399
R765 B.n328 B.n153 59.5399
R766 B.n48 B.n47 59.5399
R767 B.n610 B.n55 59.5399
R768 B.n705 B.n20 37.62
R769 B.n532 B.n531 37.62
R770 B.n423 B.n118 37.62
R771 B.n250 B.n249 37.62
R772 B B.n759 18.0485
R773 B.n701 B.n20 10.6151
R774 B.n701 B.n700 10.6151
R775 B.n700 B.n699 10.6151
R776 B.n699 B.n22 10.6151
R777 B.n695 B.n22 10.6151
R778 B.n695 B.n694 10.6151
R779 B.n694 B.n693 10.6151
R780 B.n693 B.n24 10.6151
R781 B.n689 B.n24 10.6151
R782 B.n689 B.n688 10.6151
R783 B.n688 B.n687 10.6151
R784 B.n687 B.n26 10.6151
R785 B.n683 B.n26 10.6151
R786 B.n683 B.n682 10.6151
R787 B.n682 B.n681 10.6151
R788 B.n681 B.n28 10.6151
R789 B.n677 B.n28 10.6151
R790 B.n677 B.n676 10.6151
R791 B.n676 B.n675 10.6151
R792 B.n675 B.n30 10.6151
R793 B.n671 B.n30 10.6151
R794 B.n671 B.n670 10.6151
R795 B.n670 B.n669 10.6151
R796 B.n669 B.n32 10.6151
R797 B.n665 B.n32 10.6151
R798 B.n665 B.n664 10.6151
R799 B.n664 B.n663 10.6151
R800 B.n663 B.n34 10.6151
R801 B.n659 B.n34 10.6151
R802 B.n659 B.n658 10.6151
R803 B.n658 B.n657 10.6151
R804 B.n657 B.n36 10.6151
R805 B.n653 B.n36 10.6151
R806 B.n653 B.n652 10.6151
R807 B.n652 B.n651 10.6151
R808 B.n651 B.n38 10.6151
R809 B.n647 B.n38 10.6151
R810 B.n647 B.n646 10.6151
R811 B.n646 B.n645 10.6151
R812 B.n645 B.n40 10.6151
R813 B.n641 B.n40 10.6151
R814 B.n641 B.n640 10.6151
R815 B.n640 B.n639 10.6151
R816 B.n639 B.n42 10.6151
R817 B.n635 B.n42 10.6151
R818 B.n635 B.n634 10.6151
R819 B.n634 B.n633 10.6151
R820 B.n633 B.n44 10.6151
R821 B.n629 B.n44 10.6151
R822 B.n629 B.n628 10.6151
R823 B.n628 B.n627 10.6151
R824 B.n624 B.n623 10.6151
R825 B.n623 B.n622 10.6151
R826 B.n622 B.n50 10.6151
R827 B.n618 B.n50 10.6151
R828 B.n618 B.n617 10.6151
R829 B.n617 B.n616 10.6151
R830 B.n616 B.n52 10.6151
R831 B.n612 B.n52 10.6151
R832 B.n612 B.n611 10.6151
R833 B.n609 B.n56 10.6151
R834 B.n605 B.n56 10.6151
R835 B.n605 B.n604 10.6151
R836 B.n604 B.n603 10.6151
R837 B.n603 B.n58 10.6151
R838 B.n599 B.n58 10.6151
R839 B.n599 B.n598 10.6151
R840 B.n598 B.n597 10.6151
R841 B.n597 B.n60 10.6151
R842 B.n593 B.n60 10.6151
R843 B.n593 B.n592 10.6151
R844 B.n592 B.n591 10.6151
R845 B.n591 B.n62 10.6151
R846 B.n587 B.n62 10.6151
R847 B.n587 B.n586 10.6151
R848 B.n586 B.n585 10.6151
R849 B.n585 B.n64 10.6151
R850 B.n581 B.n64 10.6151
R851 B.n581 B.n580 10.6151
R852 B.n580 B.n579 10.6151
R853 B.n579 B.n66 10.6151
R854 B.n575 B.n66 10.6151
R855 B.n575 B.n574 10.6151
R856 B.n574 B.n573 10.6151
R857 B.n573 B.n68 10.6151
R858 B.n569 B.n68 10.6151
R859 B.n569 B.n568 10.6151
R860 B.n568 B.n567 10.6151
R861 B.n567 B.n70 10.6151
R862 B.n563 B.n70 10.6151
R863 B.n563 B.n562 10.6151
R864 B.n562 B.n561 10.6151
R865 B.n561 B.n72 10.6151
R866 B.n557 B.n72 10.6151
R867 B.n557 B.n556 10.6151
R868 B.n556 B.n555 10.6151
R869 B.n555 B.n74 10.6151
R870 B.n551 B.n74 10.6151
R871 B.n551 B.n550 10.6151
R872 B.n550 B.n549 10.6151
R873 B.n549 B.n76 10.6151
R874 B.n545 B.n76 10.6151
R875 B.n545 B.n544 10.6151
R876 B.n544 B.n543 10.6151
R877 B.n543 B.n78 10.6151
R878 B.n539 B.n78 10.6151
R879 B.n539 B.n538 10.6151
R880 B.n538 B.n537 10.6151
R881 B.n537 B.n80 10.6151
R882 B.n533 B.n80 10.6151
R883 B.n533 B.n532 10.6151
R884 B.n424 B.n423 10.6151
R885 B.n425 B.n424 10.6151
R886 B.n425 B.n116 10.6151
R887 B.n429 B.n116 10.6151
R888 B.n430 B.n429 10.6151
R889 B.n431 B.n430 10.6151
R890 B.n431 B.n114 10.6151
R891 B.n435 B.n114 10.6151
R892 B.n436 B.n435 10.6151
R893 B.n437 B.n436 10.6151
R894 B.n437 B.n112 10.6151
R895 B.n441 B.n112 10.6151
R896 B.n442 B.n441 10.6151
R897 B.n443 B.n442 10.6151
R898 B.n443 B.n110 10.6151
R899 B.n447 B.n110 10.6151
R900 B.n448 B.n447 10.6151
R901 B.n449 B.n448 10.6151
R902 B.n449 B.n108 10.6151
R903 B.n453 B.n108 10.6151
R904 B.n454 B.n453 10.6151
R905 B.n455 B.n454 10.6151
R906 B.n455 B.n106 10.6151
R907 B.n459 B.n106 10.6151
R908 B.n460 B.n459 10.6151
R909 B.n461 B.n460 10.6151
R910 B.n461 B.n104 10.6151
R911 B.n465 B.n104 10.6151
R912 B.n466 B.n465 10.6151
R913 B.n467 B.n466 10.6151
R914 B.n467 B.n102 10.6151
R915 B.n471 B.n102 10.6151
R916 B.n472 B.n471 10.6151
R917 B.n473 B.n472 10.6151
R918 B.n473 B.n100 10.6151
R919 B.n477 B.n100 10.6151
R920 B.n478 B.n477 10.6151
R921 B.n479 B.n478 10.6151
R922 B.n479 B.n98 10.6151
R923 B.n483 B.n98 10.6151
R924 B.n484 B.n483 10.6151
R925 B.n485 B.n484 10.6151
R926 B.n485 B.n96 10.6151
R927 B.n489 B.n96 10.6151
R928 B.n490 B.n489 10.6151
R929 B.n491 B.n490 10.6151
R930 B.n491 B.n94 10.6151
R931 B.n495 B.n94 10.6151
R932 B.n496 B.n495 10.6151
R933 B.n497 B.n496 10.6151
R934 B.n497 B.n92 10.6151
R935 B.n501 B.n92 10.6151
R936 B.n502 B.n501 10.6151
R937 B.n503 B.n502 10.6151
R938 B.n503 B.n90 10.6151
R939 B.n507 B.n90 10.6151
R940 B.n508 B.n507 10.6151
R941 B.n509 B.n508 10.6151
R942 B.n509 B.n88 10.6151
R943 B.n513 B.n88 10.6151
R944 B.n514 B.n513 10.6151
R945 B.n515 B.n514 10.6151
R946 B.n515 B.n86 10.6151
R947 B.n519 B.n86 10.6151
R948 B.n520 B.n519 10.6151
R949 B.n521 B.n520 10.6151
R950 B.n521 B.n84 10.6151
R951 B.n525 B.n84 10.6151
R952 B.n526 B.n525 10.6151
R953 B.n527 B.n526 10.6151
R954 B.n527 B.n82 10.6151
R955 B.n531 B.n82 10.6151
R956 B.n251 B.n250 10.6151
R957 B.n251 B.n178 10.6151
R958 B.n255 B.n178 10.6151
R959 B.n256 B.n255 10.6151
R960 B.n257 B.n256 10.6151
R961 B.n257 B.n176 10.6151
R962 B.n261 B.n176 10.6151
R963 B.n262 B.n261 10.6151
R964 B.n263 B.n262 10.6151
R965 B.n263 B.n174 10.6151
R966 B.n267 B.n174 10.6151
R967 B.n268 B.n267 10.6151
R968 B.n269 B.n268 10.6151
R969 B.n269 B.n172 10.6151
R970 B.n273 B.n172 10.6151
R971 B.n274 B.n273 10.6151
R972 B.n275 B.n274 10.6151
R973 B.n275 B.n170 10.6151
R974 B.n279 B.n170 10.6151
R975 B.n280 B.n279 10.6151
R976 B.n281 B.n280 10.6151
R977 B.n281 B.n168 10.6151
R978 B.n285 B.n168 10.6151
R979 B.n286 B.n285 10.6151
R980 B.n287 B.n286 10.6151
R981 B.n287 B.n166 10.6151
R982 B.n291 B.n166 10.6151
R983 B.n292 B.n291 10.6151
R984 B.n293 B.n292 10.6151
R985 B.n293 B.n164 10.6151
R986 B.n297 B.n164 10.6151
R987 B.n298 B.n297 10.6151
R988 B.n299 B.n298 10.6151
R989 B.n299 B.n162 10.6151
R990 B.n303 B.n162 10.6151
R991 B.n304 B.n303 10.6151
R992 B.n305 B.n304 10.6151
R993 B.n305 B.n160 10.6151
R994 B.n309 B.n160 10.6151
R995 B.n310 B.n309 10.6151
R996 B.n311 B.n310 10.6151
R997 B.n311 B.n158 10.6151
R998 B.n315 B.n158 10.6151
R999 B.n316 B.n315 10.6151
R1000 B.n317 B.n316 10.6151
R1001 B.n317 B.n156 10.6151
R1002 B.n321 B.n156 10.6151
R1003 B.n322 B.n321 10.6151
R1004 B.n323 B.n322 10.6151
R1005 B.n323 B.n154 10.6151
R1006 B.n327 B.n154 10.6151
R1007 B.n330 B.n329 10.6151
R1008 B.n330 B.n150 10.6151
R1009 B.n334 B.n150 10.6151
R1010 B.n335 B.n334 10.6151
R1011 B.n336 B.n335 10.6151
R1012 B.n336 B.n148 10.6151
R1013 B.n340 B.n148 10.6151
R1014 B.n341 B.n340 10.6151
R1015 B.n342 B.n341 10.6151
R1016 B.n346 B.n345 10.6151
R1017 B.n347 B.n346 10.6151
R1018 B.n347 B.n142 10.6151
R1019 B.n351 B.n142 10.6151
R1020 B.n352 B.n351 10.6151
R1021 B.n353 B.n352 10.6151
R1022 B.n353 B.n140 10.6151
R1023 B.n357 B.n140 10.6151
R1024 B.n358 B.n357 10.6151
R1025 B.n359 B.n358 10.6151
R1026 B.n359 B.n138 10.6151
R1027 B.n363 B.n138 10.6151
R1028 B.n364 B.n363 10.6151
R1029 B.n365 B.n364 10.6151
R1030 B.n365 B.n136 10.6151
R1031 B.n369 B.n136 10.6151
R1032 B.n370 B.n369 10.6151
R1033 B.n371 B.n370 10.6151
R1034 B.n371 B.n134 10.6151
R1035 B.n375 B.n134 10.6151
R1036 B.n376 B.n375 10.6151
R1037 B.n377 B.n376 10.6151
R1038 B.n377 B.n132 10.6151
R1039 B.n381 B.n132 10.6151
R1040 B.n382 B.n381 10.6151
R1041 B.n383 B.n382 10.6151
R1042 B.n383 B.n130 10.6151
R1043 B.n387 B.n130 10.6151
R1044 B.n388 B.n387 10.6151
R1045 B.n389 B.n388 10.6151
R1046 B.n389 B.n128 10.6151
R1047 B.n393 B.n128 10.6151
R1048 B.n394 B.n393 10.6151
R1049 B.n395 B.n394 10.6151
R1050 B.n395 B.n126 10.6151
R1051 B.n399 B.n126 10.6151
R1052 B.n400 B.n399 10.6151
R1053 B.n401 B.n400 10.6151
R1054 B.n401 B.n124 10.6151
R1055 B.n405 B.n124 10.6151
R1056 B.n406 B.n405 10.6151
R1057 B.n407 B.n406 10.6151
R1058 B.n407 B.n122 10.6151
R1059 B.n411 B.n122 10.6151
R1060 B.n412 B.n411 10.6151
R1061 B.n413 B.n412 10.6151
R1062 B.n413 B.n120 10.6151
R1063 B.n417 B.n120 10.6151
R1064 B.n418 B.n417 10.6151
R1065 B.n419 B.n418 10.6151
R1066 B.n419 B.n118 10.6151
R1067 B.n249 B.n180 10.6151
R1068 B.n245 B.n180 10.6151
R1069 B.n245 B.n244 10.6151
R1070 B.n244 B.n243 10.6151
R1071 B.n243 B.n182 10.6151
R1072 B.n239 B.n182 10.6151
R1073 B.n239 B.n238 10.6151
R1074 B.n238 B.n237 10.6151
R1075 B.n237 B.n184 10.6151
R1076 B.n233 B.n184 10.6151
R1077 B.n233 B.n232 10.6151
R1078 B.n232 B.n231 10.6151
R1079 B.n231 B.n186 10.6151
R1080 B.n227 B.n186 10.6151
R1081 B.n227 B.n226 10.6151
R1082 B.n226 B.n225 10.6151
R1083 B.n225 B.n188 10.6151
R1084 B.n221 B.n188 10.6151
R1085 B.n221 B.n220 10.6151
R1086 B.n220 B.n219 10.6151
R1087 B.n219 B.n190 10.6151
R1088 B.n215 B.n190 10.6151
R1089 B.n215 B.n214 10.6151
R1090 B.n214 B.n213 10.6151
R1091 B.n213 B.n192 10.6151
R1092 B.n209 B.n192 10.6151
R1093 B.n209 B.n208 10.6151
R1094 B.n208 B.n207 10.6151
R1095 B.n207 B.n194 10.6151
R1096 B.n203 B.n194 10.6151
R1097 B.n203 B.n202 10.6151
R1098 B.n202 B.n201 10.6151
R1099 B.n201 B.n196 10.6151
R1100 B.n197 B.n196 10.6151
R1101 B.n197 B.n0 10.6151
R1102 B.n755 B.n1 10.6151
R1103 B.n755 B.n754 10.6151
R1104 B.n754 B.n753 10.6151
R1105 B.n753 B.n4 10.6151
R1106 B.n749 B.n4 10.6151
R1107 B.n749 B.n748 10.6151
R1108 B.n748 B.n747 10.6151
R1109 B.n747 B.n6 10.6151
R1110 B.n743 B.n6 10.6151
R1111 B.n743 B.n742 10.6151
R1112 B.n742 B.n741 10.6151
R1113 B.n741 B.n8 10.6151
R1114 B.n737 B.n8 10.6151
R1115 B.n737 B.n736 10.6151
R1116 B.n736 B.n735 10.6151
R1117 B.n735 B.n10 10.6151
R1118 B.n731 B.n10 10.6151
R1119 B.n731 B.n730 10.6151
R1120 B.n730 B.n729 10.6151
R1121 B.n729 B.n12 10.6151
R1122 B.n725 B.n12 10.6151
R1123 B.n725 B.n724 10.6151
R1124 B.n724 B.n723 10.6151
R1125 B.n723 B.n14 10.6151
R1126 B.n719 B.n14 10.6151
R1127 B.n719 B.n718 10.6151
R1128 B.n718 B.n717 10.6151
R1129 B.n717 B.n16 10.6151
R1130 B.n713 B.n16 10.6151
R1131 B.n713 B.n712 10.6151
R1132 B.n712 B.n711 10.6151
R1133 B.n711 B.n18 10.6151
R1134 B.n707 B.n18 10.6151
R1135 B.n707 B.n706 10.6151
R1136 B.n706 B.n705 10.6151
R1137 B.n627 B.n48 9.36635
R1138 B.n610 B.n609 9.36635
R1139 B.n328 B.n327 9.36635
R1140 B.n345 B.n146 9.36635
R1141 B.n759 B.n0 2.81026
R1142 B.n759 B.n1 2.81026
R1143 B.n624 B.n48 1.24928
R1144 B.n611 B.n610 1.24928
R1145 B.n329 B.n328 1.24928
R1146 B.n342 B.n146 1.24928
R1147 VN.n0 VN.t2 167.694
R1148 VN.n1 VN.t1 167.694
R1149 VN.n0 VN.t3 166.792
R1150 VN.n1 VN.t0 166.792
R1151 VN VN.n1 53.6039
R1152 VN VN.n0 3.41072
R1153 VDD2.n2 VDD2.n0 114.73
R1154 VDD2.n2 VDD2.n1 69.2478
R1155 VDD2.n1 VDD2.t0 2.07352
R1156 VDD2.n1 VDD2.t2 2.07352
R1157 VDD2.n0 VDD2.t3 2.07352
R1158 VDD2.n0 VDD2.t1 2.07352
R1159 VDD2 VDD2.n2 0.0586897
R1160 VTAIL.n5 VTAIL.t3 54.6422
R1161 VTAIL.n4 VTAIL.t6 54.6422
R1162 VTAIL.n3 VTAIL.t7 54.6422
R1163 VTAIL.n6 VTAIL.t2 54.6421
R1164 VTAIL.n7 VTAIL.t4 54.6421
R1165 VTAIL.n0 VTAIL.t5 54.6421
R1166 VTAIL.n1 VTAIL.t1 54.6421
R1167 VTAIL.n2 VTAIL.t0 54.6421
R1168 VTAIL.n7 VTAIL.n6 28.6341
R1169 VTAIL.n3 VTAIL.n2 28.6341
R1170 VTAIL.n4 VTAIL.n3 2.7505
R1171 VTAIL.n6 VTAIL.n5 2.7505
R1172 VTAIL.n2 VTAIL.n1 2.7505
R1173 VTAIL VTAIL.n0 1.43369
R1174 VTAIL VTAIL.n7 1.31731
R1175 VTAIL.n5 VTAIL.n4 0.470328
R1176 VTAIL.n1 VTAIL.n0 0.470328
R1177 VP.n4 VP.t1 167.694
R1178 VP.n4 VP.t0 166.792
R1179 VP.n16 VP.n0 161.3
R1180 VP.n15 VP.n14 161.3
R1181 VP.n13 VP.n1 161.3
R1182 VP.n12 VP.n11 161.3
R1183 VP.n10 VP.n2 161.3
R1184 VP.n9 VP.n8 161.3
R1185 VP.n7 VP.n3 161.3
R1186 VP.n5 VP.t3 132.13
R1187 VP.n17 VP.t2 132.13
R1188 VP.n6 VP.n5 106.236
R1189 VP.n18 VP.n17 106.236
R1190 VP.n6 VP.n4 53.3251
R1191 VP.n11 VP.n10 40.577
R1192 VP.n11 VP.n1 40.577
R1193 VP.n9 VP.n3 24.5923
R1194 VP.n10 VP.n9 24.5923
R1195 VP.n15 VP.n1 24.5923
R1196 VP.n16 VP.n15 24.5923
R1197 VP.n5 VP.n3 4.67295
R1198 VP.n17 VP.n16 4.67295
R1199 VP.n7 VP.n6 0.278335
R1200 VP.n18 VP.n0 0.278335
R1201 VP.n8 VP.n7 0.189894
R1202 VP.n8 VP.n2 0.189894
R1203 VP.n12 VP.n2 0.189894
R1204 VP.n13 VP.n12 0.189894
R1205 VP.n14 VP.n13 0.189894
R1206 VP.n14 VP.n0 0.189894
R1207 VP VP.n18 0.153485
R1208 VDD1 VDD1.n1 115.254
R1209 VDD1 VDD1.n0 69.306
R1210 VDD1.n0 VDD1.t2 2.07352
R1211 VDD1.n0 VDD1.t3 2.07352
R1212 VDD1.n1 VDD1.t0 2.07352
R1213 VDD1.n1 VDD1.t1 2.07352
C0 w_n2884_n4104# VDD1 1.59867f
C1 VP VDD2 0.411023f
C2 B w_n2884_n4104# 10.5975f
C3 VTAIL VDD2 6.35618f
C4 VN VDD2 6.21681f
C5 B VDD1 1.40621f
C6 w_n2884_n4104# VDD2 1.66055f
C7 VP VTAIL 6.01109f
C8 VP VN 7.0537f
C9 VN VTAIL 5.99698f
C10 VDD1 VDD2 1.08517f
C11 w_n2884_n4104# VP 5.36386f
C12 B VDD2 1.46267f
C13 w_n2884_n4104# VTAIL 4.800991f
C14 w_n2884_n4104# VN 4.99245f
C15 VP VDD1 6.47762f
C16 B VP 1.82282f
C17 VTAIL VDD1 6.30023f
C18 VN VDD1 0.149408f
C19 B VTAIL 6.28569f
C20 B VN 1.20528f
C21 VDD2 VSUBS 1.078942f
C22 VDD1 VSUBS 6.34865f
C23 VTAIL VSUBS 1.417514f
C24 VN VSUBS 5.70435f
C25 VP VSUBS 2.548733f
C26 B VSUBS 4.811381f
C27 w_n2884_n4104# VSUBS 0.145042p
C28 VDD1.t2 VSUBS 0.333745f
C29 VDD1.t3 VSUBS 0.333745f
C30 VDD1.n0 VSUBS 2.72062f
C31 VDD1.t0 VSUBS 0.333745f
C32 VDD1.t1 VSUBS 0.333745f
C33 VDD1.n1 VSUBS 3.63896f
C34 VP.n0 VSUBS 0.039589f
C35 VP.t2 VSUBS 3.69384f
C36 VP.n1 VSUBS 0.05937f
C37 VP.n2 VSUBS 0.03003f
C38 VP.n3 VSUBS 0.03342f
C39 VP.t0 VSUBS 4.00318f
C40 VP.t1 VSUBS 4.01096f
C41 VP.n4 VSUBS 4.35457f
C42 VP.t3 VSUBS 3.69384f
C43 VP.n5 VSUBS 1.3871f
C44 VP.n6 VSUBS 1.82337f
C45 VP.n7 VSUBS 0.039589f
C46 VP.n8 VSUBS 0.03003f
C47 VP.n9 VSUBS 0.055688f
C48 VP.n10 VSUBS 0.05937f
C49 VP.n11 VSUBS 0.024254f
C50 VP.n12 VSUBS 0.03003f
C51 VP.n13 VSUBS 0.03003f
C52 VP.n14 VSUBS 0.03003f
C53 VP.n15 VSUBS 0.055688f
C54 VP.n16 VSUBS 0.03342f
C55 VP.n17 VSUBS 1.3871f
C56 VP.n18 VSUBS 0.055492f
C57 VTAIL.t5 VSUBS 2.84415f
C58 VTAIL.n0 VSUBS 0.795668f
C59 VTAIL.t1 VSUBS 2.84415f
C60 VTAIL.n1 VSUBS 0.892793f
C61 VTAIL.t0 VSUBS 2.84415f
C62 VTAIL.n2 VSUBS 2.36891f
C63 VTAIL.t7 VSUBS 2.84417f
C64 VTAIL.n3 VSUBS 2.36889f
C65 VTAIL.t6 VSUBS 2.84417f
C66 VTAIL.n4 VSUBS 0.892769f
C67 VTAIL.t3 VSUBS 2.84417f
C68 VTAIL.n5 VSUBS 0.892769f
C69 VTAIL.t2 VSUBS 2.84415f
C70 VTAIL.n6 VSUBS 2.36891f
C71 VTAIL.t4 VSUBS 2.84415f
C72 VTAIL.n7 VSUBS 2.26321f
C73 VDD2.t3 VSUBS 0.331103f
C74 VDD2.t1 VSUBS 0.331103f
C75 VDD2.n0 VSUBS 3.58301f
C76 VDD2.t0 VSUBS 0.331103f
C77 VDD2.t2 VSUBS 0.331103f
C78 VDD2.n1 VSUBS 2.69844f
C79 VDD2.n2 VSUBS 4.7516f
C80 VN.t2 VSUBS 3.89208f
C81 VN.t3 VSUBS 3.88454f
C82 VN.n0 VSUBS 2.44363f
C83 VN.t1 VSUBS 3.89208f
C84 VN.t0 VSUBS 3.88454f
C85 VN.n1 VSUBS 4.24082f
C86 B.n0 VSUBS 0.003867f
C87 B.n1 VSUBS 0.003867f
C88 B.n2 VSUBS 0.006115f
C89 B.n3 VSUBS 0.006115f
C90 B.n4 VSUBS 0.006115f
C91 B.n5 VSUBS 0.006115f
C92 B.n6 VSUBS 0.006115f
C93 B.n7 VSUBS 0.006115f
C94 B.n8 VSUBS 0.006115f
C95 B.n9 VSUBS 0.006115f
C96 B.n10 VSUBS 0.006115f
C97 B.n11 VSUBS 0.006115f
C98 B.n12 VSUBS 0.006115f
C99 B.n13 VSUBS 0.006115f
C100 B.n14 VSUBS 0.006115f
C101 B.n15 VSUBS 0.006115f
C102 B.n16 VSUBS 0.006115f
C103 B.n17 VSUBS 0.006115f
C104 B.n18 VSUBS 0.006115f
C105 B.n19 VSUBS 0.006115f
C106 B.n20 VSUBS 0.01605f
C107 B.n21 VSUBS 0.006115f
C108 B.n22 VSUBS 0.006115f
C109 B.n23 VSUBS 0.006115f
C110 B.n24 VSUBS 0.006115f
C111 B.n25 VSUBS 0.006115f
C112 B.n26 VSUBS 0.006115f
C113 B.n27 VSUBS 0.006115f
C114 B.n28 VSUBS 0.006115f
C115 B.n29 VSUBS 0.006115f
C116 B.n30 VSUBS 0.006115f
C117 B.n31 VSUBS 0.006115f
C118 B.n32 VSUBS 0.006115f
C119 B.n33 VSUBS 0.006115f
C120 B.n34 VSUBS 0.006115f
C121 B.n35 VSUBS 0.006115f
C122 B.n36 VSUBS 0.006115f
C123 B.n37 VSUBS 0.006115f
C124 B.n38 VSUBS 0.006115f
C125 B.n39 VSUBS 0.006115f
C126 B.n40 VSUBS 0.006115f
C127 B.n41 VSUBS 0.006115f
C128 B.n42 VSUBS 0.006115f
C129 B.n43 VSUBS 0.006115f
C130 B.n44 VSUBS 0.006115f
C131 B.n45 VSUBS 0.006115f
C132 B.t2 VSUBS 0.457613f
C133 B.t1 VSUBS 0.477791f
C134 B.t0 VSUBS 1.76589f
C135 B.n46 VSUBS 0.264046f
C136 B.n47 VSUBS 0.063873f
C137 B.n48 VSUBS 0.014167f
C138 B.n49 VSUBS 0.006115f
C139 B.n50 VSUBS 0.006115f
C140 B.n51 VSUBS 0.006115f
C141 B.n52 VSUBS 0.006115f
C142 B.n53 VSUBS 0.006115f
C143 B.t8 VSUBS 0.457599f
C144 B.t7 VSUBS 0.47778f
C145 B.t6 VSUBS 1.76589f
C146 B.n54 VSUBS 0.264057f
C147 B.n55 VSUBS 0.063887f
C148 B.n56 VSUBS 0.006115f
C149 B.n57 VSUBS 0.006115f
C150 B.n58 VSUBS 0.006115f
C151 B.n59 VSUBS 0.006115f
C152 B.n60 VSUBS 0.006115f
C153 B.n61 VSUBS 0.006115f
C154 B.n62 VSUBS 0.006115f
C155 B.n63 VSUBS 0.006115f
C156 B.n64 VSUBS 0.006115f
C157 B.n65 VSUBS 0.006115f
C158 B.n66 VSUBS 0.006115f
C159 B.n67 VSUBS 0.006115f
C160 B.n68 VSUBS 0.006115f
C161 B.n69 VSUBS 0.006115f
C162 B.n70 VSUBS 0.006115f
C163 B.n71 VSUBS 0.006115f
C164 B.n72 VSUBS 0.006115f
C165 B.n73 VSUBS 0.006115f
C166 B.n74 VSUBS 0.006115f
C167 B.n75 VSUBS 0.006115f
C168 B.n76 VSUBS 0.006115f
C169 B.n77 VSUBS 0.006115f
C170 B.n78 VSUBS 0.006115f
C171 B.n79 VSUBS 0.006115f
C172 B.n80 VSUBS 0.006115f
C173 B.n81 VSUBS 0.01605f
C174 B.n82 VSUBS 0.006115f
C175 B.n83 VSUBS 0.006115f
C176 B.n84 VSUBS 0.006115f
C177 B.n85 VSUBS 0.006115f
C178 B.n86 VSUBS 0.006115f
C179 B.n87 VSUBS 0.006115f
C180 B.n88 VSUBS 0.006115f
C181 B.n89 VSUBS 0.006115f
C182 B.n90 VSUBS 0.006115f
C183 B.n91 VSUBS 0.006115f
C184 B.n92 VSUBS 0.006115f
C185 B.n93 VSUBS 0.006115f
C186 B.n94 VSUBS 0.006115f
C187 B.n95 VSUBS 0.006115f
C188 B.n96 VSUBS 0.006115f
C189 B.n97 VSUBS 0.006115f
C190 B.n98 VSUBS 0.006115f
C191 B.n99 VSUBS 0.006115f
C192 B.n100 VSUBS 0.006115f
C193 B.n101 VSUBS 0.006115f
C194 B.n102 VSUBS 0.006115f
C195 B.n103 VSUBS 0.006115f
C196 B.n104 VSUBS 0.006115f
C197 B.n105 VSUBS 0.006115f
C198 B.n106 VSUBS 0.006115f
C199 B.n107 VSUBS 0.006115f
C200 B.n108 VSUBS 0.006115f
C201 B.n109 VSUBS 0.006115f
C202 B.n110 VSUBS 0.006115f
C203 B.n111 VSUBS 0.006115f
C204 B.n112 VSUBS 0.006115f
C205 B.n113 VSUBS 0.006115f
C206 B.n114 VSUBS 0.006115f
C207 B.n115 VSUBS 0.006115f
C208 B.n116 VSUBS 0.006115f
C209 B.n117 VSUBS 0.006115f
C210 B.n118 VSUBS 0.01605f
C211 B.n119 VSUBS 0.006115f
C212 B.n120 VSUBS 0.006115f
C213 B.n121 VSUBS 0.006115f
C214 B.n122 VSUBS 0.006115f
C215 B.n123 VSUBS 0.006115f
C216 B.n124 VSUBS 0.006115f
C217 B.n125 VSUBS 0.006115f
C218 B.n126 VSUBS 0.006115f
C219 B.n127 VSUBS 0.006115f
C220 B.n128 VSUBS 0.006115f
C221 B.n129 VSUBS 0.006115f
C222 B.n130 VSUBS 0.006115f
C223 B.n131 VSUBS 0.006115f
C224 B.n132 VSUBS 0.006115f
C225 B.n133 VSUBS 0.006115f
C226 B.n134 VSUBS 0.006115f
C227 B.n135 VSUBS 0.006115f
C228 B.n136 VSUBS 0.006115f
C229 B.n137 VSUBS 0.006115f
C230 B.n138 VSUBS 0.006115f
C231 B.n139 VSUBS 0.006115f
C232 B.n140 VSUBS 0.006115f
C233 B.n141 VSUBS 0.006115f
C234 B.n142 VSUBS 0.006115f
C235 B.n143 VSUBS 0.006115f
C236 B.t4 VSUBS 0.457599f
C237 B.t5 VSUBS 0.47778f
C238 B.t3 VSUBS 1.76589f
C239 B.n144 VSUBS 0.264057f
C240 B.n145 VSUBS 0.063887f
C241 B.n146 VSUBS 0.014167f
C242 B.n147 VSUBS 0.006115f
C243 B.n148 VSUBS 0.006115f
C244 B.n149 VSUBS 0.006115f
C245 B.n150 VSUBS 0.006115f
C246 B.n151 VSUBS 0.006115f
C247 B.t10 VSUBS 0.457613f
C248 B.t11 VSUBS 0.477791f
C249 B.t9 VSUBS 1.76589f
C250 B.n152 VSUBS 0.264046f
C251 B.n153 VSUBS 0.063873f
C252 B.n154 VSUBS 0.006115f
C253 B.n155 VSUBS 0.006115f
C254 B.n156 VSUBS 0.006115f
C255 B.n157 VSUBS 0.006115f
C256 B.n158 VSUBS 0.006115f
C257 B.n159 VSUBS 0.006115f
C258 B.n160 VSUBS 0.006115f
C259 B.n161 VSUBS 0.006115f
C260 B.n162 VSUBS 0.006115f
C261 B.n163 VSUBS 0.006115f
C262 B.n164 VSUBS 0.006115f
C263 B.n165 VSUBS 0.006115f
C264 B.n166 VSUBS 0.006115f
C265 B.n167 VSUBS 0.006115f
C266 B.n168 VSUBS 0.006115f
C267 B.n169 VSUBS 0.006115f
C268 B.n170 VSUBS 0.006115f
C269 B.n171 VSUBS 0.006115f
C270 B.n172 VSUBS 0.006115f
C271 B.n173 VSUBS 0.006115f
C272 B.n174 VSUBS 0.006115f
C273 B.n175 VSUBS 0.006115f
C274 B.n176 VSUBS 0.006115f
C275 B.n177 VSUBS 0.006115f
C276 B.n178 VSUBS 0.006115f
C277 B.n179 VSUBS 0.01605f
C278 B.n180 VSUBS 0.006115f
C279 B.n181 VSUBS 0.006115f
C280 B.n182 VSUBS 0.006115f
C281 B.n183 VSUBS 0.006115f
C282 B.n184 VSUBS 0.006115f
C283 B.n185 VSUBS 0.006115f
C284 B.n186 VSUBS 0.006115f
C285 B.n187 VSUBS 0.006115f
C286 B.n188 VSUBS 0.006115f
C287 B.n189 VSUBS 0.006115f
C288 B.n190 VSUBS 0.006115f
C289 B.n191 VSUBS 0.006115f
C290 B.n192 VSUBS 0.006115f
C291 B.n193 VSUBS 0.006115f
C292 B.n194 VSUBS 0.006115f
C293 B.n195 VSUBS 0.006115f
C294 B.n196 VSUBS 0.006115f
C295 B.n197 VSUBS 0.006115f
C296 B.n198 VSUBS 0.006115f
C297 B.n199 VSUBS 0.006115f
C298 B.n200 VSUBS 0.006115f
C299 B.n201 VSUBS 0.006115f
C300 B.n202 VSUBS 0.006115f
C301 B.n203 VSUBS 0.006115f
C302 B.n204 VSUBS 0.006115f
C303 B.n205 VSUBS 0.006115f
C304 B.n206 VSUBS 0.006115f
C305 B.n207 VSUBS 0.006115f
C306 B.n208 VSUBS 0.006115f
C307 B.n209 VSUBS 0.006115f
C308 B.n210 VSUBS 0.006115f
C309 B.n211 VSUBS 0.006115f
C310 B.n212 VSUBS 0.006115f
C311 B.n213 VSUBS 0.006115f
C312 B.n214 VSUBS 0.006115f
C313 B.n215 VSUBS 0.006115f
C314 B.n216 VSUBS 0.006115f
C315 B.n217 VSUBS 0.006115f
C316 B.n218 VSUBS 0.006115f
C317 B.n219 VSUBS 0.006115f
C318 B.n220 VSUBS 0.006115f
C319 B.n221 VSUBS 0.006115f
C320 B.n222 VSUBS 0.006115f
C321 B.n223 VSUBS 0.006115f
C322 B.n224 VSUBS 0.006115f
C323 B.n225 VSUBS 0.006115f
C324 B.n226 VSUBS 0.006115f
C325 B.n227 VSUBS 0.006115f
C326 B.n228 VSUBS 0.006115f
C327 B.n229 VSUBS 0.006115f
C328 B.n230 VSUBS 0.006115f
C329 B.n231 VSUBS 0.006115f
C330 B.n232 VSUBS 0.006115f
C331 B.n233 VSUBS 0.006115f
C332 B.n234 VSUBS 0.006115f
C333 B.n235 VSUBS 0.006115f
C334 B.n236 VSUBS 0.006115f
C335 B.n237 VSUBS 0.006115f
C336 B.n238 VSUBS 0.006115f
C337 B.n239 VSUBS 0.006115f
C338 B.n240 VSUBS 0.006115f
C339 B.n241 VSUBS 0.006115f
C340 B.n242 VSUBS 0.006115f
C341 B.n243 VSUBS 0.006115f
C342 B.n244 VSUBS 0.006115f
C343 B.n245 VSUBS 0.006115f
C344 B.n246 VSUBS 0.006115f
C345 B.n247 VSUBS 0.006115f
C346 B.n248 VSUBS 0.015423f
C347 B.n249 VSUBS 0.015423f
C348 B.n250 VSUBS 0.01605f
C349 B.n251 VSUBS 0.006115f
C350 B.n252 VSUBS 0.006115f
C351 B.n253 VSUBS 0.006115f
C352 B.n254 VSUBS 0.006115f
C353 B.n255 VSUBS 0.006115f
C354 B.n256 VSUBS 0.006115f
C355 B.n257 VSUBS 0.006115f
C356 B.n258 VSUBS 0.006115f
C357 B.n259 VSUBS 0.006115f
C358 B.n260 VSUBS 0.006115f
C359 B.n261 VSUBS 0.006115f
C360 B.n262 VSUBS 0.006115f
C361 B.n263 VSUBS 0.006115f
C362 B.n264 VSUBS 0.006115f
C363 B.n265 VSUBS 0.006115f
C364 B.n266 VSUBS 0.006115f
C365 B.n267 VSUBS 0.006115f
C366 B.n268 VSUBS 0.006115f
C367 B.n269 VSUBS 0.006115f
C368 B.n270 VSUBS 0.006115f
C369 B.n271 VSUBS 0.006115f
C370 B.n272 VSUBS 0.006115f
C371 B.n273 VSUBS 0.006115f
C372 B.n274 VSUBS 0.006115f
C373 B.n275 VSUBS 0.006115f
C374 B.n276 VSUBS 0.006115f
C375 B.n277 VSUBS 0.006115f
C376 B.n278 VSUBS 0.006115f
C377 B.n279 VSUBS 0.006115f
C378 B.n280 VSUBS 0.006115f
C379 B.n281 VSUBS 0.006115f
C380 B.n282 VSUBS 0.006115f
C381 B.n283 VSUBS 0.006115f
C382 B.n284 VSUBS 0.006115f
C383 B.n285 VSUBS 0.006115f
C384 B.n286 VSUBS 0.006115f
C385 B.n287 VSUBS 0.006115f
C386 B.n288 VSUBS 0.006115f
C387 B.n289 VSUBS 0.006115f
C388 B.n290 VSUBS 0.006115f
C389 B.n291 VSUBS 0.006115f
C390 B.n292 VSUBS 0.006115f
C391 B.n293 VSUBS 0.006115f
C392 B.n294 VSUBS 0.006115f
C393 B.n295 VSUBS 0.006115f
C394 B.n296 VSUBS 0.006115f
C395 B.n297 VSUBS 0.006115f
C396 B.n298 VSUBS 0.006115f
C397 B.n299 VSUBS 0.006115f
C398 B.n300 VSUBS 0.006115f
C399 B.n301 VSUBS 0.006115f
C400 B.n302 VSUBS 0.006115f
C401 B.n303 VSUBS 0.006115f
C402 B.n304 VSUBS 0.006115f
C403 B.n305 VSUBS 0.006115f
C404 B.n306 VSUBS 0.006115f
C405 B.n307 VSUBS 0.006115f
C406 B.n308 VSUBS 0.006115f
C407 B.n309 VSUBS 0.006115f
C408 B.n310 VSUBS 0.006115f
C409 B.n311 VSUBS 0.006115f
C410 B.n312 VSUBS 0.006115f
C411 B.n313 VSUBS 0.006115f
C412 B.n314 VSUBS 0.006115f
C413 B.n315 VSUBS 0.006115f
C414 B.n316 VSUBS 0.006115f
C415 B.n317 VSUBS 0.006115f
C416 B.n318 VSUBS 0.006115f
C417 B.n319 VSUBS 0.006115f
C418 B.n320 VSUBS 0.006115f
C419 B.n321 VSUBS 0.006115f
C420 B.n322 VSUBS 0.006115f
C421 B.n323 VSUBS 0.006115f
C422 B.n324 VSUBS 0.006115f
C423 B.n325 VSUBS 0.006115f
C424 B.n326 VSUBS 0.006115f
C425 B.n327 VSUBS 0.005755f
C426 B.n328 VSUBS 0.014167f
C427 B.n329 VSUBS 0.003417f
C428 B.n330 VSUBS 0.006115f
C429 B.n331 VSUBS 0.006115f
C430 B.n332 VSUBS 0.006115f
C431 B.n333 VSUBS 0.006115f
C432 B.n334 VSUBS 0.006115f
C433 B.n335 VSUBS 0.006115f
C434 B.n336 VSUBS 0.006115f
C435 B.n337 VSUBS 0.006115f
C436 B.n338 VSUBS 0.006115f
C437 B.n339 VSUBS 0.006115f
C438 B.n340 VSUBS 0.006115f
C439 B.n341 VSUBS 0.006115f
C440 B.n342 VSUBS 0.003417f
C441 B.n343 VSUBS 0.006115f
C442 B.n344 VSUBS 0.006115f
C443 B.n345 VSUBS 0.005755f
C444 B.n346 VSUBS 0.006115f
C445 B.n347 VSUBS 0.006115f
C446 B.n348 VSUBS 0.006115f
C447 B.n349 VSUBS 0.006115f
C448 B.n350 VSUBS 0.006115f
C449 B.n351 VSUBS 0.006115f
C450 B.n352 VSUBS 0.006115f
C451 B.n353 VSUBS 0.006115f
C452 B.n354 VSUBS 0.006115f
C453 B.n355 VSUBS 0.006115f
C454 B.n356 VSUBS 0.006115f
C455 B.n357 VSUBS 0.006115f
C456 B.n358 VSUBS 0.006115f
C457 B.n359 VSUBS 0.006115f
C458 B.n360 VSUBS 0.006115f
C459 B.n361 VSUBS 0.006115f
C460 B.n362 VSUBS 0.006115f
C461 B.n363 VSUBS 0.006115f
C462 B.n364 VSUBS 0.006115f
C463 B.n365 VSUBS 0.006115f
C464 B.n366 VSUBS 0.006115f
C465 B.n367 VSUBS 0.006115f
C466 B.n368 VSUBS 0.006115f
C467 B.n369 VSUBS 0.006115f
C468 B.n370 VSUBS 0.006115f
C469 B.n371 VSUBS 0.006115f
C470 B.n372 VSUBS 0.006115f
C471 B.n373 VSUBS 0.006115f
C472 B.n374 VSUBS 0.006115f
C473 B.n375 VSUBS 0.006115f
C474 B.n376 VSUBS 0.006115f
C475 B.n377 VSUBS 0.006115f
C476 B.n378 VSUBS 0.006115f
C477 B.n379 VSUBS 0.006115f
C478 B.n380 VSUBS 0.006115f
C479 B.n381 VSUBS 0.006115f
C480 B.n382 VSUBS 0.006115f
C481 B.n383 VSUBS 0.006115f
C482 B.n384 VSUBS 0.006115f
C483 B.n385 VSUBS 0.006115f
C484 B.n386 VSUBS 0.006115f
C485 B.n387 VSUBS 0.006115f
C486 B.n388 VSUBS 0.006115f
C487 B.n389 VSUBS 0.006115f
C488 B.n390 VSUBS 0.006115f
C489 B.n391 VSUBS 0.006115f
C490 B.n392 VSUBS 0.006115f
C491 B.n393 VSUBS 0.006115f
C492 B.n394 VSUBS 0.006115f
C493 B.n395 VSUBS 0.006115f
C494 B.n396 VSUBS 0.006115f
C495 B.n397 VSUBS 0.006115f
C496 B.n398 VSUBS 0.006115f
C497 B.n399 VSUBS 0.006115f
C498 B.n400 VSUBS 0.006115f
C499 B.n401 VSUBS 0.006115f
C500 B.n402 VSUBS 0.006115f
C501 B.n403 VSUBS 0.006115f
C502 B.n404 VSUBS 0.006115f
C503 B.n405 VSUBS 0.006115f
C504 B.n406 VSUBS 0.006115f
C505 B.n407 VSUBS 0.006115f
C506 B.n408 VSUBS 0.006115f
C507 B.n409 VSUBS 0.006115f
C508 B.n410 VSUBS 0.006115f
C509 B.n411 VSUBS 0.006115f
C510 B.n412 VSUBS 0.006115f
C511 B.n413 VSUBS 0.006115f
C512 B.n414 VSUBS 0.006115f
C513 B.n415 VSUBS 0.006115f
C514 B.n416 VSUBS 0.006115f
C515 B.n417 VSUBS 0.006115f
C516 B.n418 VSUBS 0.006115f
C517 B.n419 VSUBS 0.006115f
C518 B.n420 VSUBS 0.006115f
C519 B.n421 VSUBS 0.01605f
C520 B.n422 VSUBS 0.015423f
C521 B.n423 VSUBS 0.015423f
C522 B.n424 VSUBS 0.006115f
C523 B.n425 VSUBS 0.006115f
C524 B.n426 VSUBS 0.006115f
C525 B.n427 VSUBS 0.006115f
C526 B.n428 VSUBS 0.006115f
C527 B.n429 VSUBS 0.006115f
C528 B.n430 VSUBS 0.006115f
C529 B.n431 VSUBS 0.006115f
C530 B.n432 VSUBS 0.006115f
C531 B.n433 VSUBS 0.006115f
C532 B.n434 VSUBS 0.006115f
C533 B.n435 VSUBS 0.006115f
C534 B.n436 VSUBS 0.006115f
C535 B.n437 VSUBS 0.006115f
C536 B.n438 VSUBS 0.006115f
C537 B.n439 VSUBS 0.006115f
C538 B.n440 VSUBS 0.006115f
C539 B.n441 VSUBS 0.006115f
C540 B.n442 VSUBS 0.006115f
C541 B.n443 VSUBS 0.006115f
C542 B.n444 VSUBS 0.006115f
C543 B.n445 VSUBS 0.006115f
C544 B.n446 VSUBS 0.006115f
C545 B.n447 VSUBS 0.006115f
C546 B.n448 VSUBS 0.006115f
C547 B.n449 VSUBS 0.006115f
C548 B.n450 VSUBS 0.006115f
C549 B.n451 VSUBS 0.006115f
C550 B.n452 VSUBS 0.006115f
C551 B.n453 VSUBS 0.006115f
C552 B.n454 VSUBS 0.006115f
C553 B.n455 VSUBS 0.006115f
C554 B.n456 VSUBS 0.006115f
C555 B.n457 VSUBS 0.006115f
C556 B.n458 VSUBS 0.006115f
C557 B.n459 VSUBS 0.006115f
C558 B.n460 VSUBS 0.006115f
C559 B.n461 VSUBS 0.006115f
C560 B.n462 VSUBS 0.006115f
C561 B.n463 VSUBS 0.006115f
C562 B.n464 VSUBS 0.006115f
C563 B.n465 VSUBS 0.006115f
C564 B.n466 VSUBS 0.006115f
C565 B.n467 VSUBS 0.006115f
C566 B.n468 VSUBS 0.006115f
C567 B.n469 VSUBS 0.006115f
C568 B.n470 VSUBS 0.006115f
C569 B.n471 VSUBS 0.006115f
C570 B.n472 VSUBS 0.006115f
C571 B.n473 VSUBS 0.006115f
C572 B.n474 VSUBS 0.006115f
C573 B.n475 VSUBS 0.006115f
C574 B.n476 VSUBS 0.006115f
C575 B.n477 VSUBS 0.006115f
C576 B.n478 VSUBS 0.006115f
C577 B.n479 VSUBS 0.006115f
C578 B.n480 VSUBS 0.006115f
C579 B.n481 VSUBS 0.006115f
C580 B.n482 VSUBS 0.006115f
C581 B.n483 VSUBS 0.006115f
C582 B.n484 VSUBS 0.006115f
C583 B.n485 VSUBS 0.006115f
C584 B.n486 VSUBS 0.006115f
C585 B.n487 VSUBS 0.006115f
C586 B.n488 VSUBS 0.006115f
C587 B.n489 VSUBS 0.006115f
C588 B.n490 VSUBS 0.006115f
C589 B.n491 VSUBS 0.006115f
C590 B.n492 VSUBS 0.006115f
C591 B.n493 VSUBS 0.006115f
C592 B.n494 VSUBS 0.006115f
C593 B.n495 VSUBS 0.006115f
C594 B.n496 VSUBS 0.006115f
C595 B.n497 VSUBS 0.006115f
C596 B.n498 VSUBS 0.006115f
C597 B.n499 VSUBS 0.006115f
C598 B.n500 VSUBS 0.006115f
C599 B.n501 VSUBS 0.006115f
C600 B.n502 VSUBS 0.006115f
C601 B.n503 VSUBS 0.006115f
C602 B.n504 VSUBS 0.006115f
C603 B.n505 VSUBS 0.006115f
C604 B.n506 VSUBS 0.006115f
C605 B.n507 VSUBS 0.006115f
C606 B.n508 VSUBS 0.006115f
C607 B.n509 VSUBS 0.006115f
C608 B.n510 VSUBS 0.006115f
C609 B.n511 VSUBS 0.006115f
C610 B.n512 VSUBS 0.006115f
C611 B.n513 VSUBS 0.006115f
C612 B.n514 VSUBS 0.006115f
C613 B.n515 VSUBS 0.006115f
C614 B.n516 VSUBS 0.006115f
C615 B.n517 VSUBS 0.006115f
C616 B.n518 VSUBS 0.006115f
C617 B.n519 VSUBS 0.006115f
C618 B.n520 VSUBS 0.006115f
C619 B.n521 VSUBS 0.006115f
C620 B.n522 VSUBS 0.006115f
C621 B.n523 VSUBS 0.006115f
C622 B.n524 VSUBS 0.006115f
C623 B.n525 VSUBS 0.006115f
C624 B.n526 VSUBS 0.006115f
C625 B.n527 VSUBS 0.006115f
C626 B.n528 VSUBS 0.006115f
C627 B.n529 VSUBS 0.006115f
C628 B.n530 VSUBS 0.015423f
C629 B.n531 VSUBS 0.01605f
C630 B.n532 VSUBS 0.015423f
C631 B.n533 VSUBS 0.006115f
C632 B.n534 VSUBS 0.006115f
C633 B.n535 VSUBS 0.006115f
C634 B.n536 VSUBS 0.006115f
C635 B.n537 VSUBS 0.006115f
C636 B.n538 VSUBS 0.006115f
C637 B.n539 VSUBS 0.006115f
C638 B.n540 VSUBS 0.006115f
C639 B.n541 VSUBS 0.006115f
C640 B.n542 VSUBS 0.006115f
C641 B.n543 VSUBS 0.006115f
C642 B.n544 VSUBS 0.006115f
C643 B.n545 VSUBS 0.006115f
C644 B.n546 VSUBS 0.006115f
C645 B.n547 VSUBS 0.006115f
C646 B.n548 VSUBS 0.006115f
C647 B.n549 VSUBS 0.006115f
C648 B.n550 VSUBS 0.006115f
C649 B.n551 VSUBS 0.006115f
C650 B.n552 VSUBS 0.006115f
C651 B.n553 VSUBS 0.006115f
C652 B.n554 VSUBS 0.006115f
C653 B.n555 VSUBS 0.006115f
C654 B.n556 VSUBS 0.006115f
C655 B.n557 VSUBS 0.006115f
C656 B.n558 VSUBS 0.006115f
C657 B.n559 VSUBS 0.006115f
C658 B.n560 VSUBS 0.006115f
C659 B.n561 VSUBS 0.006115f
C660 B.n562 VSUBS 0.006115f
C661 B.n563 VSUBS 0.006115f
C662 B.n564 VSUBS 0.006115f
C663 B.n565 VSUBS 0.006115f
C664 B.n566 VSUBS 0.006115f
C665 B.n567 VSUBS 0.006115f
C666 B.n568 VSUBS 0.006115f
C667 B.n569 VSUBS 0.006115f
C668 B.n570 VSUBS 0.006115f
C669 B.n571 VSUBS 0.006115f
C670 B.n572 VSUBS 0.006115f
C671 B.n573 VSUBS 0.006115f
C672 B.n574 VSUBS 0.006115f
C673 B.n575 VSUBS 0.006115f
C674 B.n576 VSUBS 0.006115f
C675 B.n577 VSUBS 0.006115f
C676 B.n578 VSUBS 0.006115f
C677 B.n579 VSUBS 0.006115f
C678 B.n580 VSUBS 0.006115f
C679 B.n581 VSUBS 0.006115f
C680 B.n582 VSUBS 0.006115f
C681 B.n583 VSUBS 0.006115f
C682 B.n584 VSUBS 0.006115f
C683 B.n585 VSUBS 0.006115f
C684 B.n586 VSUBS 0.006115f
C685 B.n587 VSUBS 0.006115f
C686 B.n588 VSUBS 0.006115f
C687 B.n589 VSUBS 0.006115f
C688 B.n590 VSUBS 0.006115f
C689 B.n591 VSUBS 0.006115f
C690 B.n592 VSUBS 0.006115f
C691 B.n593 VSUBS 0.006115f
C692 B.n594 VSUBS 0.006115f
C693 B.n595 VSUBS 0.006115f
C694 B.n596 VSUBS 0.006115f
C695 B.n597 VSUBS 0.006115f
C696 B.n598 VSUBS 0.006115f
C697 B.n599 VSUBS 0.006115f
C698 B.n600 VSUBS 0.006115f
C699 B.n601 VSUBS 0.006115f
C700 B.n602 VSUBS 0.006115f
C701 B.n603 VSUBS 0.006115f
C702 B.n604 VSUBS 0.006115f
C703 B.n605 VSUBS 0.006115f
C704 B.n606 VSUBS 0.006115f
C705 B.n607 VSUBS 0.006115f
C706 B.n608 VSUBS 0.006115f
C707 B.n609 VSUBS 0.005755f
C708 B.n610 VSUBS 0.014167f
C709 B.n611 VSUBS 0.003417f
C710 B.n612 VSUBS 0.006115f
C711 B.n613 VSUBS 0.006115f
C712 B.n614 VSUBS 0.006115f
C713 B.n615 VSUBS 0.006115f
C714 B.n616 VSUBS 0.006115f
C715 B.n617 VSUBS 0.006115f
C716 B.n618 VSUBS 0.006115f
C717 B.n619 VSUBS 0.006115f
C718 B.n620 VSUBS 0.006115f
C719 B.n621 VSUBS 0.006115f
C720 B.n622 VSUBS 0.006115f
C721 B.n623 VSUBS 0.006115f
C722 B.n624 VSUBS 0.003417f
C723 B.n625 VSUBS 0.006115f
C724 B.n626 VSUBS 0.006115f
C725 B.n627 VSUBS 0.005755f
C726 B.n628 VSUBS 0.006115f
C727 B.n629 VSUBS 0.006115f
C728 B.n630 VSUBS 0.006115f
C729 B.n631 VSUBS 0.006115f
C730 B.n632 VSUBS 0.006115f
C731 B.n633 VSUBS 0.006115f
C732 B.n634 VSUBS 0.006115f
C733 B.n635 VSUBS 0.006115f
C734 B.n636 VSUBS 0.006115f
C735 B.n637 VSUBS 0.006115f
C736 B.n638 VSUBS 0.006115f
C737 B.n639 VSUBS 0.006115f
C738 B.n640 VSUBS 0.006115f
C739 B.n641 VSUBS 0.006115f
C740 B.n642 VSUBS 0.006115f
C741 B.n643 VSUBS 0.006115f
C742 B.n644 VSUBS 0.006115f
C743 B.n645 VSUBS 0.006115f
C744 B.n646 VSUBS 0.006115f
C745 B.n647 VSUBS 0.006115f
C746 B.n648 VSUBS 0.006115f
C747 B.n649 VSUBS 0.006115f
C748 B.n650 VSUBS 0.006115f
C749 B.n651 VSUBS 0.006115f
C750 B.n652 VSUBS 0.006115f
C751 B.n653 VSUBS 0.006115f
C752 B.n654 VSUBS 0.006115f
C753 B.n655 VSUBS 0.006115f
C754 B.n656 VSUBS 0.006115f
C755 B.n657 VSUBS 0.006115f
C756 B.n658 VSUBS 0.006115f
C757 B.n659 VSUBS 0.006115f
C758 B.n660 VSUBS 0.006115f
C759 B.n661 VSUBS 0.006115f
C760 B.n662 VSUBS 0.006115f
C761 B.n663 VSUBS 0.006115f
C762 B.n664 VSUBS 0.006115f
C763 B.n665 VSUBS 0.006115f
C764 B.n666 VSUBS 0.006115f
C765 B.n667 VSUBS 0.006115f
C766 B.n668 VSUBS 0.006115f
C767 B.n669 VSUBS 0.006115f
C768 B.n670 VSUBS 0.006115f
C769 B.n671 VSUBS 0.006115f
C770 B.n672 VSUBS 0.006115f
C771 B.n673 VSUBS 0.006115f
C772 B.n674 VSUBS 0.006115f
C773 B.n675 VSUBS 0.006115f
C774 B.n676 VSUBS 0.006115f
C775 B.n677 VSUBS 0.006115f
C776 B.n678 VSUBS 0.006115f
C777 B.n679 VSUBS 0.006115f
C778 B.n680 VSUBS 0.006115f
C779 B.n681 VSUBS 0.006115f
C780 B.n682 VSUBS 0.006115f
C781 B.n683 VSUBS 0.006115f
C782 B.n684 VSUBS 0.006115f
C783 B.n685 VSUBS 0.006115f
C784 B.n686 VSUBS 0.006115f
C785 B.n687 VSUBS 0.006115f
C786 B.n688 VSUBS 0.006115f
C787 B.n689 VSUBS 0.006115f
C788 B.n690 VSUBS 0.006115f
C789 B.n691 VSUBS 0.006115f
C790 B.n692 VSUBS 0.006115f
C791 B.n693 VSUBS 0.006115f
C792 B.n694 VSUBS 0.006115f
C793 B.n695 VSUBS 0.006115f
C794 B.n696 VSUBS 0.006115f
C795 B.n697 VSUBS 0.006115f
C796 B.n698 VSUBS 0.006115f
C797 B.n699 VSUBS 0.006115f
C798 B.n700 VSUBS 0.006115f
C799 B.n701 VSUBS 0.006115f
C800 B.n702 VSUBS 0.006115f
C801 B.n703 VSUBS 0.01605f
C802 B.n704 VSUBS 0.015423f
C803 B.n705 VSUBS 0.015423f
C804 B.n706 VSUBS 0.006115f
C805 B.n707 VSUBS 0.006115f
C806 B.n708 VSUBS 0.006115f
C807 B.n709 VSUBS 0.006115f
C808 B.n710 VSUBS 0.006115f
C809 B.n711 VSUBS 0.006115f
C810 B.n712 VSUBS 0.006115f
C811 B.n713 VSUBS 0.006115f
C812 B.n714 VSUBS 0.006115f
C813 B.n715 VSUBS 0.006115f
C814 B.n716 VSUBS 0.006115f
C815 B.n717 VSUBS 0.006115f
C816 B.n718 VSUBS 0.006115f
C817 B.n719 VSUBS 0.006115f
C818 B.n720 VSUBS 0.006115f
C819 B.n721 VSUBS 0.006115f
C820 B.n722 VSUBS 0.006115f
C821 B.n723 VSUBS 0.006115f
C822 B.n724 VSUBS 0.006115f
C823 B.n725 VSUBS 0.006115f
C824 B.n726 VSUBS 0.006115f
C825 B.n727 VSUBS 0.006115f
C826 B.n728 VSUBS 0.006115f
C827 B.n729 VSUBS 0.006115f
C828 B.n730 VSUBS 0.006115f
C829 B.n731 VSUBS 0.006115f
C830 B.n732 VSUBS 0.006115f
C831 B.n733 VSUBS 0.006115f
C832 B.n734 VSUBS 0.006115f
C833 B.n735 VSUBS 0.006115f
C834 B.n736 VSUBS 0.006115f
C835 B.n737 VSUBS 0.006115f
C836 B.n738 VSUBS 0.006115f
C837 B.n739 VSUBS 0.006115f
C838 B.n740 VSUBS 0.006115f
C839 B.n741 VSUBS 0.006115f
C840 B.n742 VSUBS 0.006115f
C841 B.n743 VSUBS 0.006115f
C842 B.n744 VSUBS 0.006115f
C843 B.n745 VSUBS 0.006115f
C844 B.n746 VSUBS 0.006115f
C845 B.n747 VSUBS 0.006115f
C846 B.n748 VSUBS 0.006115f
C847 B.n749 VSUBS 0.006115f
C848 B.n750 VSUBS 0.006115f
C849 B.n751 VSUBS 0.006115f
C850 B.n752 VSUBS 0.006115f
C851 B.n753 VSUBS 0.006115f
C852 B.n754 VSUBS 0.006115f
C853 B.n755 VSUBS 0.006115f
C854 B.n756 VSUBS 0.006115f
C855 B.n757 VSUBS 0.006115f
C856 B.n758 VSUBS 0.006115f
C857 B.n759 VSUBS 0.013846f
.ends

