* NGSPICE file created from diff_pair_sample_0849.ext - technology: sky130A

.subckt diff_pair_sample_0849 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X1 VTAIL.t0 VN.t0 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X2 VTAIL.t10 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X3 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0 ps=0 w=5.66 l=3.5
X4 VTAIL.t4 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0.9339 ps=5.99 w=5.66 l=3.5
X5 VTAIL.t6 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X6 VDD1.t5 VP.t2 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=2.2074 ps=12.1 w=5.66 l=3.5
X7 VTAIL.t9 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0.9339 ps=5.99 w=5.66 l=3.5
X8 VDD2.t4 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X9 VDD1.t3 VP.t4 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X10 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0 ps=0 w=5.66 l=3.5
X11 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=2.2074 ps=12.1 w=5.66 l=3.5
X12 VTAIL.t8 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0.9339 ps=5.99 w=5.66 l=3.5
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0 ps=0 w=5.66 l=3.5
X14 VDD1.t1 VP.t6 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=2.2074 ps=12.1 w=5.66 l=3.5
X15 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=2.2074 ps=12.1 w=5.66 l=3.5
X16 VTAIL.t12 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X17 VDD2.t1 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9339 pd=5.99 as=0.9339 ps=5.99 w=5.66 l=3.5
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0 ps=0 w=5.66 l=3.5
X19 VTAIL.t7 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2074 pd=12.1 as=0.9339 ps=5.99 w=5.66 l=3.5
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n17 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n85 VP.n84 161.3
R16 VP.n83 VP.n1 161.3
R17 VP.n82 VP.n81 161.3
R18 VP.n80 VP.n2 161.3
R19 VP.n79 VP.n78 161.3
R20 VP.n77 VP.n3 161.3
R21 VP.n76 VP.n75 161.3
R22 VP.n74 VP.n4 161.3
R23 VP.n73 VP.n72 161.3
R24 VP.n70 VP.n5 161.3
R25 VP.n69 VP.n68 161.3
R26 VP.n67 VP.n6 161.3
R27 VP.n66 VP.n65 161.3
R28 VP.n64 VP.n7 161.3
R29 VP.n63 VP.n62 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n59 VP.n9 161.3
R32 VP.n58 VP.n57 161.3
R33 VP.n56 VP.n10 161.3
R34 VP.n55 VP.n54 161.3
R35 VP.n53 VP.n11 161.3
R36 VP.n52 VP.n51 161.3
R37 VP.n50 VP.n12 161.3
R38 VP.n49 VP.n48 78.1956
R39 VP.n86 VP.n0 78.1956
R40 VP.n47 VP.n13 78.1956
R41 VP.n22 VP.t3 72.7364
R42 VP.n54 VP.n10 56.5617
R43 VP.n78 VP.n2 56.5617
R44 VP.n39 VP.n15 56.5617
R45 VP.n22 VP.n21 54.4908
R46 VP.n49 VP.n47 50.4238
R47 VP.n65 VP.n6 40.577
R48 VP.n69 VP.n6 40.577
R49 VP.n30 VP.n19 40.577
R50 VP.n26 VP.n19 40.577
R51 VP.n48 VP.t5 38.9736
R52 VP.n8 VP.t4 38.9736
R53 VP.n71 VP.t7 38.9736
R54 VP.n0 VP.t2 38.9736
R55 VP.n13 VP.t6 38.9736
R56 VP.n32 VP.t1 38.9736
R57 VP.n21 VP.t0 38.9736
R58 VP.n52 VP.n12 24.5923
R59 VP.n53 VP.n52 24.5923
R60 VP.n54 VP.n53 24.5923
R61 VP.n58 VP.n10 24.5923
R62 VP.n59 VP.n58 24.5923
R63 VP.n60 VP.n59 24.5923
R64 VP.n64 VP.n63 24.5923
R65 VP.n65 VP.n64 24.5923
R66 VP.n70 VP.n69 24.5923
R67 VP.n72 VP.n70 24.5923
R68 VP.n76 VP.n4 24.5923
R69 VP.n77 VP.n76 24.5923
R70 VP.n78 VP.n77 24.5923
R71 VP.n82 VP.n2 24.5923
R72 VP.n83 VP.n82 24.5923
R73 VP.n84 VP.n83 24.5923
R74 VP.n43 VP.n15 24.5923
R75 VP.n44 VP.n43 24.5923
R76 VP.n45 VP.n44 24.5923
R77 VP.n31 VP.n30 24.5923
R78 VP.n33 VP.n31 24.5923
R79 VP.n37 VP.n17 24.5923
R80 VP.n38 VP.n37 24.5923
R81 VP.n39 VP.n38 24.5923
R82 VP.n25 VP.n24 24.5923
R83 VP.n26 VP.n25 24.5923
R84 VP.n63 VP.n8 20.4117
R85 VP.n72 VP.n71 20.4117
R86 VP.n33 VP.n32 20.4117
R87 VP.n24 VP.n21 20.4117
R88 VP.n48 VP.n12 12.0505
R89 VP.n84 VP.n0 12.0505
R90 VP.n45 VP.n13 12.0505
R91 VP.n60 VP.n8 4.18111
R92 VP.n71 VP.n4 4.18111
R93 VP.n32 VP.n17 4.18111
R94 VP.n23 VP.n22 3.07938
R95 VP.n47 VP.n46 0.354861
R96 VP.n50 VP.n49 0.354861
R97 VP.n86 VP.n85 0.354861
R98 VP VP.n86 0.267071
R99 VP.n23 VP.n20 0.189894
R100 VP.n27 VP.n20 0.189894
R101 VP.n28 VP.n27 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n29 VP.n18 0.189894
R104 VP.n34 VP.n18 0.189894
R105 VP.n35 VP.n34 0.189894
R106 VP.n36 VP.n35 0.189894
R107 VP.n36 VP.n16 0.189894
R108 VP.n40 VP.n16 0.189894
R109 VP.n41 VP.n40 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n42 VP.n14 0.189894
R112 VP.n46 VP.n14 0.189894
R113 VP.n51 VP.n50 0.189894
R114 VP.n51 VP.n11 0.189894
R115 VP.n55 VP.n11 0.189894
R116 VP.n56 VP.n55 0.189894
R117 VP.n57 VP.n56 0.189894
R118 VP.n57 VP.n9 0.189894
R119 VP.n61 VP.n9 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n62 VP.n7 0.189894
R122 VP.n66 VP.n7 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n68 VP.n5 0.189894
R126 VP.n73 VP.n5 0.189894
R127 VP.n74 VP.n73 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n75 VP.n3 0.189894
R130 VP.n79 VP.n3 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n81 VP.n1 0.189894
R134 VP.n85 VP.n1 0.189894
R135 VTAIL.n11 VTAIL.t9 55.0773
R136 VTAIL.n10 VTAIL.t5 55.0773
R137 VTAIL.n7 VTAIL.t4 55.0773
R138 VTAIL.n15 VTAIL.t3 55.0771
R139 VTAIL.n2 VTAIL.t7 55.0771
R140 VTAIL.n3 VTAIL.t15 55.0771
R141 VTAIL.n6 VTAIL.t8 55.0771
R142 VTAIL.n14 VTAIL.t11 55.0771
R143 VTAIL.n13 VTAIL.n12 51.5791
R144 VTAIL.n9 VTAIL.n8 51.5791
R145 VTAIL.n1 VTAIL.n0 51.5789
R146 VTAIL.n5 VTAIL.n4 51.5789
R147 VTAIL.n15 VTAIL.n14 20.5479
R148 VTAIL.n7 VTAIL.n6 20.5479
R149 VTAIL.n0 VTAIL.t2 3.49873
R150 VTAIL.n0 VTAIL.t0 3.49873
R151 VTAIL.n4 VTAIL.t14 3.49873
R152 VTAIL.n4 VTAIL.t12 3.49873
R153 VTAIL.n12 VTAIL.t13 3.49873
R154 VTAIL.n12 VTAIL.t10 3.49873
R155 VTAIL.n8 VTAIL.t1 3.49873
R156 VTAIL.n8 VTAIL.t6 3.49873
R157 VTAIL.n9 VTAIL.n7 3.30222
R158 VTAIL.n10 VTAIL.n9 3.30222
R159 VTAIL.n13 VTAIL.n11 3.30222
R160 VTAIL.n14 VTAIL.n13 3.30222
R161 VTAIL.n6 VTAIL.n5 3.30222
R162 VTAIL.n5 VTAIL.n3 3.30222
R163 VTAIL.n2 VTAIL.n1 3.30222
R164 VTAIL VTAIL.n15 3.24403
R165 VTAIL.n11 VTAIL.n10 0.470328
R166 VTAIL.n3 VTAIL.n2 0.470328
R167 VTAIL VTAIL.n1 0.0586897
R168 VDD1 VDD1.n0 69.9669
R169 VDD1.n3 VDD1.n2 69.8532
R170 VDD1.n3 VDD1.n1 69.8532
R171 VDD1.n5 VDD1.n4 68.2577
R172 VDD1.n5 VDD1.n3 44.0354
R173 VDD1.n4 VDD1.t6 3.49873
R174 VDD1.n4 VDD1.t1 3.49873
R175 VDD1.n0 VDD1.t4 3.49873
R176 VDD1.n0 VDD1.t7 3.49873
R177 VDD1.n2 VDD1.t0 3.49873
R178 VDD1.n2 VDD1.t5 3.49873
R179 VDD1.n1 VDD1.t2 3.49873
R180 VDD1.n1 VDD1.t3 3.49873
R181 VDD1 VDD1.n5 1.59317
R182 B.n800 B.n799 585
R183 B.n801 B.n800 585
R184 B.n256 B.n145 585
R185 B.n255 B.n254 585
R186 B.n253 B.n252 585
R187 B.n251 B.n250 585
R188 B.n249 B.n248 585
R189 B.n247 B.n246 585
R190 B.n245 B.n244 585
R191 B.n243 B.n242 585
R192 B.n241 B.n240 585
R193 B.n239 B.n238 585
R194 B.n237 B.n236 585
R195 B.n235 B.n234 585
R196 B.n233 B.n232 585
R197 B.n231 B.n230 585
R198 B.n229 B.n228 585
R199 B.n227 B.n226 585
R200 B.n225 B.n224 585
R201 B.n223 B.n222 585
R202 B.n221 B.n220 585
R203 B.n219 B.n218 585
R204 B.n217 B.n216 585
R205 B.n215 B.n214 585
R206 B.n213 B.n212 585
R207 B.n211 B.n210 585
R208 B.n209 B.n208 585
R209 B.n207 B.n206 585
R210 B.n205 B.n204 585
R211 B.n203 B.n202 585
R212 B.n201 B.n200 585
R213 B.n199 B.n198 585
R214 B.n197 B.n196 585
R215 B.n194 B.n193 585
R216 B.n192 B.n191 585
R217 B.n190 B.n189 585
R218 B.n188 B.n187 585
R219 B.n186 B.n185 585
R220 B.n184 B.n183 585
R221 B.n182 B.n181 585
R222 B.n180 B.n179 585
R223 B.n178 B.n177 585
R224 B.n176 B.n175 585
R225 B.n174 B.n173 585
R226 B.n172 B.n171 585
R227 B.n170 B.n169 585
R228 B.n168 B.n167 585
R229 B.n166 B.n165 585
R230 B.n164 B.n163 585
R231 B.n162 B.n161 585
R232 B.n160 B.n159 585
R233 B.n158 B.n157 585
R234 B.n156 B.n155 585
R235 B.n154 B.n153 585
R236 B.n152 B.n151 585
R237 B.n116 B.n115 585
R238 B.n798 B.n117 585
R239 B.n802 B.n117 585
R240 B.n797 B.n796 585
R241 B.n796 B.n113 585
R242 B.n795 B.n112 585
R243 B.n808 B.n112 585
R244 B.n794 B.n111 585
R245 B.n809 B.n111 585
R246 B.n793 B.n110 585
R247 B.n810 B.n110 585
R248 B.n792 B.n791 585
R249 B.n791 B.n106 585
R250 B.n790 B.n105 585
R251 B.n816 B.n105 585
R252 B.n789 B.n104 585
R253 B.n817 B.n104 585
R254 B.n788 B.n103 585
R255 B.n818 B.n103 585
R256 B.n787 B.n786 585
R257 B.n786 B.t13 585
R258 B.n785 B.n99 585
R259 B.n824 B.n99 585
R260 B.n784 B.n98 585
R261 B.n825 B.n98 585
R262 B.n783 B.n97 585
R263 B.n826 B.n97 585
R264 B.n782 B.n781 585
R265 B.n781 B.n93 585
R266 B.n780 B.n92 585
R267 B.n832 B.n92 585
R268 B.n779 B.n91 585
R269 B.n833 B.n91 585
R270 B.n778 B.n90 585
R271 B.n834 B.n90 585
R272 B.n777 B.n776 585
R273 B.n776 B.n86 585
R274 B.n775 B.n85 585
R275 B.n840 B.n85 585
R276 B.n774 B.n84 585
R277 B.n841 B.n84 585
R278 B.n773 B.n83 585
R279 B.n842 B.n83 585
R280 B.n772 B.n771 585
R281 B.n771 B.n79 585
R282 B.n770 B.n78 585
R283 B.n848 B.n78 585
R284 B.n769 B.n77 585
R285 B.n849 B.n77 585
R286 B.n768 B.n76 585
R287 B.n850 B.n76 585
R288 B.n767 B.n766 585
R289 B.n766 B.n72 585
R290 B.n765 B.n71 585
R291 B.n856 B.n71 585
R292 B.n764 B.n70 585
R293 B.n857 B.n70 585
R294 B.n763 B.n69 585
R295 B.n858 B.n69 585
R296 B.n762 B.n761 585
R297 B.n761 B.n65 585
R298 B.n760 B.n64 585
R299 B.n864 B.n64 585
R300 B.n759 B.n63 585
R301 B.n865 B.n63 585
R302 B.n758 B.n62 585
R303 B.n866 B.n62 585
R304 B.n757 B.n756 585
R305 B.n756 B.n58 585
R306 B.n755 B.n57 585
R307 B.n872 B.n57 585
R308 B.n754 B.n56 585
R309 B.n873 B.n56 585
R310 B.n753 B.n55 585
R311 B.n874 B.n55 585
R312 B.n752 B.n751 585
R313 B.n751 B.n51 585
R314 B.n750 B.n50 585
R315 B.n880 B.n50 585
R316 B.n749 B.n49 585
R317 B.n881 B.n49 585
R318 B.n748 B.n48 585
R319 B.n882 B.n48 585
R320 B.n747 B.n746 585
R321 B.n746 B.n44 585
R322 B.n745 B.n43 585
R323 B.n888 B.n43 585
R324 B.n744 B.n42 585
R325 B.n889 B.n42 585
R326 B.n743 B.n41 585
R327 B.n890 B.n41 585
R328 B.n742 B.n741 585
R329 B.n741 B.n37 585
R330 B.n740 B.n36 585
R331 B.t2 B.n36 585
R332 B.n739 B.n35 585
R333 B.n896 B.n35 585
R334 B.n738 B.n34 585
R335 B.n897 B.n34 585
R336 B.n737 B.n736 585
R337 B.n736 B.n30 585
R338 B.n735 B.n29 585
R339 B.n903 B.n29 585
R340 B.n734 B.n28 585
R341 B.n904 B.n28 585
R342 B.n733 B.n27 585
R343 B.n905 B.n27 585
R344 B.n732 B.n731 585
R345 B.n731 B.n23 585
R346 B.n730 B.n22 585
R347 B.n911 B.n22 585
R348 B.n729 B.n21 585
R349 B.n912 B.n21 585
R350 B.n728 B.n20 585
R351 B.n913 B.n20 585
R352 B.n727 B.n726 585
R353 B.n726 B.n19 585
R354 B.n725 B.n15 585
R355 B.n919 B.n15 585
R356 B.n724 B.n14 585
R357 B.n920 B.n14 585
R358 B.n723 B.n13 585
R359 B.n921 B.n13 585
R360 B.n722 B.n721 585
R361 B.n721 B.n12 585
R362 B.n720 B.n719 585
R363 B.n720 B.n8 585
R364 B.n718 B.n7 585
R365 B.n928 B.n7 585
R366 B.n717 B.n6 585
R367 B.n929 B.n6 585
R368 B.n716 B.n5 585
R369 B.n930 B.n5 585
R370 B.n715 B.n714 585
R371 B.n714 B.n4 585
R372 B.n713 B.n257 585
R373 B.n713 B.n712 585
R374 B.n703 B.n258 585
R375 B.n259 B.n258 585
R376 B.n705 B.n704 585
R377 B.n706 B.n705 585
R378 B.n702 B.n264 585
R379 B.n264 B.n263 585
R380 B.n701 B.n700 585
R381 B.n700 B.n699 585
R382 B.n266 B.n265 585
R383 B.n692 B.n266 585
R384 B.n691 B.n690 585
R385 B.n693 B.n691 585
R386 B.n689 B.n271 585
R387 B.n271 B.n270 585
R388 B.n688 B.n687 585
R389 B.n687 B.n686 585
R390 B.n273 B.n272 585
R391 B.n274 B.n273 585
R392 B.n679 B.n678 585
R393 B.n680 B.n679 585
R394 B.n677 B.n279 585
R395 B.n279 B.n278 585
R396 B.n676 B.n675 585
R397 B.n675 B.n674 585
R398 B.n281 B.n280 585
R399 B.n282 B.n281 585
R400 B.n667 B.n666 585
R401 B.n668 B.n667 585
R402 B.n665 B.n287 585
R403 B.n287 B.n286 585
R404 B.n664 B.n663 585
R405 B.n663 B.t6 585
R406 B.n289 B.n288 585
R407 B.n290 B.n289 585
R408 B.n656 B.n655 585
R409 B.n657 B.n656 585
R410 B.n654 B.n295 585
R411 B.n295 B.n294 585
R412 B.n653 B.n652 585
R413 B.n652 B.n651 585
R414 B.n297 B.n296 585
R415 B.n298 B.n297 585
R416 B.n644 B.n643 585
R417 B.n645 B.n644 585
R418 B.n642 B.n303 585
R419 B.n303 B.n302 585
R420 B.n641 B.n640 585
R421 B.n640 B.n639 585
R422 B.n305 B.n304 585
R423 B.n306 B.n305 585
R424 B.n632 B.n631 585
R425 B.n633 B.n632 585
R426 B.n630 B.n311 585
R427 B.n311 B.n310 585
R428 B.n629 B.n628 585
R429 B.n628 B.n627 585
R430 B.n313 B.n312 585
R431 B.n314 B.n313 585
R432 B.n620 B.n619 585
R433 B.n621 B.n620 585
R434 B.n618 B.n319 585
R435 B.n319 B.n318 585
R436 B.n617 B.n616 585
R437 B.n616 B.n615 585
R438 B.n321 B.n320 585
R439 B.n322 B.n321 585
R440 B.n608 B.n607 585
R441 B.n609 B.n608 585
R442 B.n606 B.n327 585
R443 B.n327 B.n326 585
R444 B.n605 B.n604 585
R445 B.n604 B.n603 585
R446 B.n329 B.n328 585
R447 B.n330 B.n329 585
R448 B.n596 B.n595 585
R449 B.n597 B.n596 585
R450 B.n594 B.n334 585
R451 B.n338 B.n334 585
R452 B.n593 B.n592 585
R453 B.n592 B.n591 585
R454 B.n336 B.n335 585
R455 B.n337 B.n336 585
R456 B.n584 B.n583 585
R457 B.n585 B.n584 585
R458 B.n582 B.n343 585
R459 B.n343 B.n342 585
R460 B.n581 B.n580 585
R461 B.n580 B.n579 585
R462 B.n345 B.n344 585
R463 B.n346 B.n345 585
R464 B.n572 B.n571 585
R465 B.n573 B.n572 585
R466 B.n570 B.n351 585
R467 B.n351 B.n350 585
R468 B.n569 B.n568 585
R469 B.n568 B.n567 585
R470 B.n353 B.n352 585
R471 B.n354 B.n353 585
R472 B.n560 B.n559 585
R473 B.n561 B.n560 585
R474 B.n558 B.n359 585
R475 B.n359 B.n358 585
R476 B.n557 B.n556 585
R477 B.n556 B.n555 585
R478 B.n361 B.n360 585
R479 B.t9 B.n361 585
R480 B.n548 B.n547 585
R481 B.n549 B.n548 585
R482 B.n546 B.n366 585
R483 B.n366 B.n365 585
R484 B.n545 B.n544 585
R485 B.n544 B.n543 585
R486 B.n368 B.n367 585
R487 B.n369 B.n368 585
R488 B.n536 B.n535 585
R489 B.n537 B.n536 585
R490 B.n534 B.n374 585
R491 B.n374 B.n373 585
R492 B.n533 B.n532 585
R493 B.n532 B.n531 585
R494 B.n376 B.n375 585
R495 B.n377 B.n376 585
R496 B.n524 B.n523 585
R497 B.n525 B.n524 585
R498 B.n380 B.n379 585
R499 B.n413 B.n412 585
R500 B.n414 B.n410 585
R501 B.n410 B.n381 585
R502 B.n416 B.n415 585
R503 B.n418 B.n409 585
R504 B.n421 B.n420 585
R505 B.n422 B.n408 585
R506 B.n424 B.n423 585
R507 B.n426 B.n407 585
R508 B.n429 B.n428 585
R509 B.n430 B.n406 585
R510 B.n432 B.n431 585
R511 B.n434 B.n405 585
R512 B.n437 B.n436 585
R513 B.n438 B.n404 585
R514 B.n440 B.n439 585
R515 B.n442 B.n403 585
R516 B.n445 B.n444 585
R517 B.n446 B.n402 585
R518 B.n448 B.n447 585
R519 B.n450 B.n401 585
R520 B.n453 B.n452 585
R521 B.n454 B.n398 585
R522 B.n457 B.n456 585
R523 B.n459 B.n397 585
R524 B.n462 B.n461 585
R525 B.n463 B.n396 585
R526 B.n465 B.n464 585
R527 B.n467 B.n395 585
R528 B.n470 B.n469 585
R529 B.n471 B.n394 585
R530 B.n476 B.n475 585
R531 B.n478 B.n393 585
R532 B.n481 B.n480 585
R533 B.n482 B.n392 585
R534 B.n484 B.n483 585
R535 B.n486 B.n391 585
R536 B.n489 B.n488 585
R537 B.n490 B.n390 585
R538 B.n492 B.n491 585
R539 B.n494 B.n389 585
R540 B.n497 B.n496 585
R541 B.n498 B.n388 585
R542 B.n500 B.n499 585
R543 B.n502 B.n387 585
R544 B.n505 B.n504 585
R545 B.n506 B.n386 585
R546 B.n508 B.n507 585
R547 B.n510 B.n385 585
R548 B.n513 B.n512 585
R549 B.n514 B.n384 585
R550 B.n516 B.n515 585
R551 B.n518 B.n383 585
R552 B.n521 B.n520 585
R553 B.n522 B.n382 585
R554 B.n527 B.n526 585
R555 B.n526 B.n525 585
R556 B.n528 B.n378 585
R557 B.n378 B.n377 585
R558 B.n530 B.n529 585
R559 B.n531 B.n530 585
R560 B.n372 B.n371 585
R561 B.n373 B.n372 585
R562 B.n539 B.n538 585
R563 B.n538 B.n537 585
R564 B.n540 B.n370 585
R565 B.n370 B.n369 585
R566 B.n542 B.n541 585
R567 B.n543 B.n542 585
R568 B.n364 B.n363 585
R569 B.n365 B.n364 585
R570 B.n551 B.n550 585
R571 B.n550 B.n549 585
R572 B.n552 B.n362 585
R573 B.n362 B.t9 585
R574 B.n554 B.n553 585
R575 B.n555 B.n554 585
R576 B.n357 B.n356 585
R577 B.n358 B.n357 585
R578 B.n563 B.n562 585
R579 B.n562 B.n561 585
R580 B.n564 B.n355 585
R581 B.n355 B.n354 585
R582 B.n566 B.n565 585
R583 B.n567 B.n566 585
R584 B.n349 B.n348 585
R585 B.n350 B.n349 585
R586 B.n575 B.n574 585
R587 B.n574 B.n573 585
R588 B.n576 B.n347 585
R589 B.n347 B.n346 585
R590 B.n578 B.n577 585
R591 B.n579 B.n578 585
R592 B.n341 B.n340 585
R593 B.n342 B.n341 585
R594 B.n587 B.n586 585
R595 B.n586 B.n585 585
R596 B.n588 B.n339 585
R597 B.n339 B.n337 585
R598 B.n590 B.n589 585
R599 B.n591 B.n590 585
R600 B.n333 B.n332 585
R601 B.n338 B.n333 585
R602 B.n599 B.n598 585
R603 B.n598 B.n597 585
R604 B.n600 B.n331 585
R605 B.n331 B.n330 585
R606 B.n602 B.n601 585
R607 B.n603 B.n602 585
R608 B.n325 B.n324 585
R609 B.n326 B.n325 585
R610 B.n611 B.n610 585
R611 B.n610 B.n609 585
R612 B.n612 B.n323 585
R613 B.n323 B.n322 585
R614 B.n614 B.n613 585
R615 B.n615 B.n614 585
R616 B.n317 B.n316 585
R617 B.n318 B.n317 585
R618 B.n623 B.n622 585
R619 B.n622 B.n621 585
R620 B.n624 B.n315 585
R621 B.n315 B.n314 585
R622 B.n626 B.n625 585
R623 B.n627 B.n626 585
R624 B.n309 B.n308 585
R625 B.n310 B.n309 585
R626 B.n635 B.n634 585
R627 B.n634 B.n633 585
R628 B.n636 B.n307 585
R629 B.n307 B.n306 585
R630 B.n638 B.n637 585
R631 B.n639 B.n638 585
R632 B.n301 B.n300 585
R633 B.n302 B.n301 585
R634 B.n647 B.n646 585
R635 B.n646 B.n645 585
R636 B.n648 B.n299 585
R637 B.n299 B.n298 585
R638 B.n650 B.n649 585
R639 B.n651 B.n650 585
R640 B.n293 B.n292 585
R641 B.n294 B.n293 585
R642 B.n659 B.n658 585
R643 B.n658 B.n657 585
R644 B.n660 B.n291 585
R645 B.n291 B.n290 585
R646 B.n662 B.n661 585
R647 B.t6 B.n662 585
R648 B.n285 B.n284 585
R649 B.n286 B.n285 585
R650 B.n670 B.n669 585
R651 B.n669 B.n668 585
R652 B.n671 B.n283 585
R653 B.n283 B.n282 585
R654 B.n673 B.n672 585
R655 B.n674 B.n673 585
R656 B.n277 B.n276 585
R657 B.n278 B.n277 585
R658 B.n682 B.n681 585
R659 B.n681 B.n680 585
R660 B.n683 B.n275 585
R661 B.n275 B.n274 585
R662 B.n685 B.n684 585
R663 B.n686 B.n685 585
R664 B.n269 B.n268 585
R665 B.n270 B.n269 585
R666 B.n695 B.n694 585
R667 B.n694 B.n693 585
R668 B.n696 B.n267 585
R669 B.n692 B.n267 585
R670 B.n698 B.n697 585
R671 B.n699 B.n698 585
R672 B.n262 B.n261 585
R673 B.n263 B.n262 585
R674 B.n708 B.n707 585
R675 B.n707 B.n706 585
R676 B.n709 B.n260 585
R677 B.n260 B.n259 585
R678 B.n711 B.n710 585
R679 B.n712 B.n711 585
R680 B.n3 B.n0 585
R681 B.n4 B.n3 585
R682 B.n927 B.n1 585
R683 B.n928 B.n927 585
R684 B.n926 B.n925 585
R685 B.n926 B.n8 585
R686 B.n924 B.n9 585
R687 B.n12 B.n9 585
R688 B.n923 B.n922 585
R689 B.n922 B.n921 585
R690 B.n11 B.n10 585
R691 B.n920 B.n11 585
R692 B.n918 B.n917 585
R693 B.n919 B.n918 585
R694 B.n916 B.n16 585
R695 B.n19 B.n16 585
R696 B.n915 B.n914 585
R697 B.n914 B.n913 585
R698 B.n18 B.n17 585
R699 B.n912 B.n18 585
R700 B.n910 B.n909 585
R701 B.n911 B.n910 585
R702 B.n908 B.n24 585
R703 B.n24 B.n23 585
R704 B.n907 B.n906 585
R705 B.n906 B.n905 585
R706 B.n26 B.n25 585
R707 B.n904 B.n26 585
R708 B.n902 B.n901 585
R709 B.n903 B.n902 585
R710 B.n900 B.n31 585
R711 B.n31 B.n30 585
R712 B.n899 B.n898 585
R713 B.n898 B.n897 585
R714 B.n33 B.n32 585
R715 B.n896 B.n33 585
R716 B.n895 B.n894 585
R717 B.t2 B.n895 585
R718 B.n893 B.n38 585
R719 B.n38 B.n37 585
R720 B.n892 B.n891 585
R721 B.n891 B.n890 585
R722 B.n40 B.n39 585
R723 B.n889 B.n40 585
R724 B.n887 B.n886 585
R725 B.n888 B.n887 585
R726 B.n885 B.n45 585
R727 B.n45 B.n44 585
R728 B.n884 B.n883 585
R729 B.n883 B.n882 585
R730 B.n47 B.n46 585
R731 B.n881 B.n47 585
R732 B.n879 B.n878 585
R733 B.n880 B.n879 585
R734 B.n877 B.n52 585
R735 B.n52 B.n51 585
R736 B.n876 B.n875 585
R737 B.n875 B.n874 585
R738 B.n54 B.n53 585
R739 B.n873 B.n54 585
R740 B.n871 B.n870 585
R741 B.n872 B.n871 585
R742 B.n869 B.n59 585
R743 B.n59 B.n58 585
R744 B.n868 B.n867 585
R745 B.n867 B.n866 585
R746 B.n61 B.n60 585
R747 B.n865 B.n61 585
R748 B.n863 B.n862 585
R749 B.n864 B.n863 585
R750 B.n861 B.n66 585
R751 B.n66 B.n65 585
R752 B.n860 B.n859 585
R753 B.n859 B.n858 585
R754 B.n68 B.n67 585
R755 B.n857 B.n68 585
R756 B.n855 B.n854 585
R757 B.n856 B.n855 585
R758 B.n853 B.n73 585
R759 B.n73 B.n72 585
R760 B.n852 B.n851 585
R761 B.n851 B.n850 585
R762 B.n75 B.n74 585
R763 B.n849 B.n75 585
R764 B.n847 B.n846 585
R765 B.n848 B.n847 585
R766 B.n845 B.n80 585
R767 B.n80 B.n79 585
R768 B.n844 B.n843 585
R769 B.n843 B.n842 585
R770 B.n82 B.n81 585
R771 B.n841 B.n82 585
R772 B.n839 B.n838 585
R773 B.n840 B.n839 585
R774 B.n837 B.n87 585
R775 B.n87 B.n86 585
R776 B.n836 B.n835 585
R777 B.n835 B.n834 585
R778 B.n89 B.n88 585
R779 B.n833 B.n89 585
R780 B.n831 B.n830 585
R781 B.n832 B.n831 585
R782 B.n829 B.n94 585
R783 B.n94 B.n93 585
R784 B.n828 B.n827 585
R785 B.n827 B.n826 585
R786 B.n96 B.n95 585
R787 B.n825 B.n96 585
R788 B.n823 B.n822 585
R789 B.n824 B.n823 585
R790 B.n821 B.n100 585
R791 B.n100 B.t13 585
R792 B.n820 B.n819 585
R793 B.n819 B.n818 585
R794 B.n102 B.n101 585
R795 B.n817 B.n102 585
R796 B.n815 B.n814 585
R797 B.n816 B.n815 585
R798 B.n813 B.n107 585
R799 B.n107 B.n106 585
R800 B.n812 B.n811 585
R801 B.n811 B.n810 585
R802 B.n109 B.n108 585
R803 B.n809 B.n109 585
R804 B.n807 B.n806 585
R805 B.n808 B.n807 585
R806 B.n805 B.n114 585
R807 B.n114 B.n113 585
R808 B.n804 B.n803 585
R809 B.n803 B.n802 585
R810 B.n931 B.n930 585
R811 B.n929 B.n2 585
R812 B.n803 B.n116 530.939
R813 B.n800 B.n117 530.939
R814 B.n524 B.n382 530.939
R815 B.n526 B.n380 530.939
R816 B.n801 B.n144 256.663
R817 B.n801 B.n143 256.663
R818 B.n801 B.n142 256.663
R819 B.n801 B.n141 256.663
R820 B.n801 B.n140 256.663
R821 B.n801 B.n139 256.663
R822 B.n801 B.n138 256.663
R823 B.n801 B.n137 256.663
R824 B.n801 B.n136 256.663
R825 B.n801 B.n135 256.663
R826 B.n801 B.n134 256.663
R827 B.n801 B.n133 256.663
R828 B.n801 B.n132 256.663
R829 B.n801 B.n131 256.663
R830 B.n801 B.n130 256.663
R831 B.n801 B.n129 256.663
R832 B.n801 B.n128 256.663
R833 B.n801 B.n127 256.663
R834 B.n801 B.n126 256.663
R835 B.n801 B.n125 256.663
R836 B.n801 B.n124 256.663
R837 B.n801 B.n123 256.663
R838 B.n801 B.n122 256.663
R839 B.n801 B.n121 256.663
R840 B.n801 B.n120 256.663
R841 B.n801 B.n119 256.663
R842 B.n801 B.n118 256.663
R843 B.n411 B.n381 256.663
R844 B.n417 B.n381 256.663
R845 B.n419 B.n381 256.663
R846 B.n425 B.n381 256.663
R847 B.n427 B.n381 256.663
R848 B.n433 B.n381 256.663
R849 B.n435 B.n381 256.663
R850 B.n441 B.n381 256.663
R851 B.n443 B.n381 256.663
R852 B.n449 B.n381 256.663
R853 B.n451 B.n381 256.663
R854 B.n458 B.n381 256.663
R855 B.n460 B.n381 256.663
R856 B.n466 B.n381 256.663
R857 B.n468 B.n381 256.663
R858 B.n477 B.n381 256.663
R859 B.n479 B.n381 256.663
R860 B.n485 B.n381 256.663
R861 B.n487 B.n381 256.663
R862 B.n493 B.n381 256.663
R863 B.n495 B.n381 256.663
R864 B.n501 B.n381 256.663
R865 B.n503 B.n381 256.663
R866 B.n509 B.n381 256.663
R867 B.n511 B.n381 256.663
R868 B.n517 B.n381 256.663
R869 B.n519 B.n381 256.663
R870 B.n933 B.n932 256.663
R871 B.n149 B.t12 248.067
R872 B.n146 B.t16 248.067
R873 B.n472 B.t8 248.067
R874 B.n399 B.t19 248.067
R875 B.n153 B.n152 163.367
R876 B.n157 B.n156 163.367
R877 B.n161 B.n160 163.367
R878 B.n165 B.n164 163.367
R879 B.n169 B.n168 163.367
R880 B.n173 B.n172 163.367
R881 B.n177 B.n176 163.367
R882 B.n181 B.n180 163.367
R883 B.n185 B.n184 163.367
R884 B.n189 B.n188 163.367
R885 B.n193 B.n192 163.367
R886 B.n198 B.n197 163.367
R887 B.n202 B.n201 163.367
R888 B.n206 B.n205 163.367
R889 B.n210 B.n209 163.367
R890 B.n214 B.n213 163.367
R891 B.n218 B.n217 163.367
R892 B.n222 B.n221 163.367
R893 B.n226 B.n225 163.367
R894 B.n230 B.n229 163.367
R895 B.n234 B.n233 163.367
R896 B.n238 B.n237 163.367
R897 B.n242 B.n241 163.367
R898 B.n246 B.n245 163.367
R899 B.n250 B.n249 163.367
R900 B.n254 B.n253 163.367
R901 B.n800 B.n145 163.367
R902 B.n524 B.n376 163.367
R903 B.n532 B.n376 163.367
R904 B.n532 B.n374 163.367
R905 B.n536 B.n374 163.367
R906 B.n536 B.n368 163.367
R907 B.n544 B.n368 163.367
R908 B.n544 B.n366 163.367
R909 B.n548 B.n366 163.367
R910 B.n548 B.n361 163.367
R911 B.n556 B.n361 163.367
R912 B.n556 B.n359 163.367
R913 B.n560 B.n359 163.367
R914 B.n560 B.n353 163.367
R915 B.n568 B.n353 163.367
R916 B.n568 B.n351 163.367
R917 B.n572 B.n351 163.367
R918 B.n572 B.n345 163.367
R919 B.n580 B.n345 163.367
R920 B.n580 B.n343 163.367
R921 B.n584 B.n343 163.367
R922 B.n584 B.n336 163.367
R923 B.n592 B.n336 163.367
R924 B.n592 B.n334 163.367
R925 B.n596 B.n334 163.367
R926 B.n596 B.n329 163.367
R927 B.n604 B.n329 163.367
R928 B.n604 B.n327 163.367
R929 B.n608 B.n327 163.367
R930 B.n608 B.n321 163.367
R931 B.n616 B.n321 163.367
R932 B.n616 B.n319 163.367
R933 B.n620 B.n319 163.367
R934 B.n620 B.n313 163.367
R935 B.n628 B.n313 163.367
R936 B.n628 B.n311 163.367
R937 B.n632 B.n311 163.367
R938 B.n632 B.n305 163.367
R939 B.n640 B.n305 163.367
R940 B.n640 B.n303 163.367
R941 B.n644 B.n303 163.367
R942 B.n644 B.n297 163.367
R943 B.n652 B.n297 163.367
R944 B.n652 B.n295 163.367
R945 B.n656 B.n295 163.367
R946 B.n656 B.n289 163.367
R947 B.n663 B.n289 163.367
R948 B.n663 B.n287 163.367
R949 B.n667 B.n287 163.367
R950 B.n667 B.n281 163.367
R951 B.n675 B.n281 163.367
R952 B.n675 B.n279 163.367
R953 B.n679 B.n279 163.367
R954 B.n679 B.n273 163.367
R955 B.n687 B.n273 163.367
R956 B.n687 B.n271 163.367
R957 B.n691 B.n271 163.367
R958 B.n691 B.n266 163.367
R959 B.n700 B.n266 163.367
R960 B.n700 B.n264 163.367
R961 B.n705 B.n264 163.367
R962 B.n705 B.n258 163.367
R963 B.n713 B.n258 163.367
R964 B.n714 B.n713 163.367
R965 B.n714 B.n5 163.367
R966 B.n6 B.n5 163.367
R967 B.n7 B.n6 163.367
R968 B.n720 B.n7 163.367
R969 B.n721 B.n720 163.367
R970 B.n721 B.n13 163.367
R971 B.n14 B.n13 163.367
R972 B.n15 B.n14 163.367
R973 B.n726 B.n15 163.367
R974 B.n726 B.n20 163.367
R975 B.n21 B.n20 163.367
R976 B.n22 B.n21 163.367
R977 B.n731 B.n22 163.367
R978 B.n731 B.n27 163.367
R979 B.n28 B.n27 163.367
R980 B.n29 B.n28 163.367
R981 B.n736 B.n29 163.367
R982 B.n736 B.n34 163.367
R983 B.n35 B.n34 163.367
R984 B.n36 B.n35 163.367
R985 B.n741 B.n36 163.367
R986 B.n741 B.n41 163.367
R987 B.n42 B.n41 163.367
R988 B.n43 B.n42 163.367
R989 B.n746 B.n43 163.367
R990 B.n746 B.n48 163.367
R991 B.n49 B.n48 163.367
R992 B.n50 B.n49 163.367
R993 B.n751 B.n50 163.367
R994 B.n751 B.n55 163.367
R995 B.n56 B.n55 163.367
R996 B.n57 B.n56 163.367
R997 B.n756 B.n57 163.367
R998 B.n756 B.n62 163.367
R999 B.n63 B.n62 163.367
R1000 B.n64 B.n63 163.367
R1001 B.n761 B.n64 163.367
R1002 B.n761 B.n69 163.367
R1003 B.n70 B.n69 163.367
R1004 B.n71 B.n70 163.367
R1005 B.n766 B.n71 163.367
R1006 B.n766 B.n76 163.367
R1007 B.n77 B.n76 163.367
R1008 B.n78 B.n77 163.367
R1009 B.n771 B.n78 163.367
R1010 B.n771 B.n83 163.367
R1011 B.n84 B.n83 163.367
R1012 B.n85 B.n84 163.367
R1013 B.n776 B.n85 163.367
R1014 B.n776 B.n90 163.367
R1015 B.n91 B.n90 163.367
R1016 B.n92 B.n91 163.367
R1017 B.n781 B.n92 163.367
R1018 B.n781 B.n97 163.367
R1019 B.n98 B.n97 163.367
R1020 B.n99 B.n98 163.367
R1021 B.n786 B.n99 163.367
R1022 B.n786 B.n103 163.367
R1023 B.n104 B.n103 163.367
R1024 B.n105 B.n104 163.367
R1025 B.n791 B.n105 163.367
R1026 B.n791 B.n110 163.367
R1027 B.n111 B.n110 163.367
R1028 B.n112 B.n111 163.367
R1029 B.n796 B.n112 163.367
R1030 B.n796 B.n117 163.367
R1031 B.n412 B.n410 163.367
R1032 B.n416 B.n410 163.367
R1033 B.n420 B.n418 163.367
R1034 B.n424 B.n408 163.367
R1035 B.n428 B.n426 163.367
R1036 B.n432 B.n406 163.367
R1037 B.n436 B.n434 163.367
R1038 B.n440 B.n404 163.367
R1039 B.n444 B.n442 163.367
R1040 B.n448 B.n402 163.367
R1041 B.n452 B.n450 163.367
R1042 B.n457 B.n398 163.367
R1043 B.n461 B.n459 163.367
R1044 B.n465 B.n396 163.367
R1045 B.n469 B.n467 163.367
R1046 B.n476 B.n394 163.367
R1047 B.n480 B.n478 163.367
R1048 B.n484 B.n392 163.367
R1049 B.n488 B.n486 163.367
R1050 B.n492 B.n390 163.367
R1051 B.n496 B.n494 163.367
R1052 B.n500 B.n388 163.367
R1053 B.n504 B.n502 163.367
R1054 B.n508 B.n386 163.367
R1055 B.n512 B.n510 163.367
R1056 B.n516 B.n384 163.367
R1057 B.n520 B.n518 163.367
R1058 B.n526 B.n378 163.367
R1059 B.n530 B.n378 163.367
R1060 B.n530 B.n372 163.367
R1061 B.n538 B.n372 163.367
R1062 B.n538 B.n370 163.367
R1063 B.n542 B.n370 163.367
R1064 B.n542 B.n364 163.367
R1065 B.n550 B.n364 163.367
R1066 B.n550 B.n362 163.367
R1067 B.n554 B.n362 163.367
R1068 B.n554 B.n357 163.367
R1069 B.n562 B.n357 163.367
R1070 B.n562 B.n355 163.367
R1071 B.n566 B.n355 163.367
R1072 B.n566 B.n349 163.367
R1073 B.n574 B.n349 163.367
R1074 B.n574 B.n347 163.367
R1075 B.n578 B.n347 163.367
R1076 B.n578 B.n341 163.367
R1077 B.n586 B.n341 163.367
R1078 B.n586 B.n339 163.367
R1079 B.n590 B.n339 163.367
R1080 B.n590 B.n333 163.367
R1081 B.n598 B.n333 163.367
R1082 B.n598 B.n331 163.367
R1083 B.n602 B.n331 163.367
R1084 B.n602 B.n325 163.367
R1085 B.n610 B.n325 163.367
R1086 B.n610 B.n323 163.367
R1087 B.n614 B.n323 163.367
R1088 B.n614 B.n317 163.367
R1089 B.n622 B.n317 163.367
R1090 B.n622 B.n315 163.367
R1091 B.n626 B.n315 163.367
R1092 B.n626 B.n309 163.367
R1093 B.n634 B.n309 163.367
R1094 B.n634 B.n307 163.367
R1095 B.n638 B.n307 163.367
R1096 B.n638 B.n301 163.367
R1097 B.n646 B.n301 163.367
R1098 B.n646 B.n299 163.367
R1099 B.n650 B.n299 163.367
R1100 B.n650 B.n293 163.367
R1101 B.n658 B.n293 163.367
R1102 B.n658 B.n291 163.367
R1103 B.n662 B.n291 163.367
R1104 B.n662 B.n285 163.367
R1105 B.n669 B.n285 163.367
R1106 B.n669 B.n283 163.367
R1107 B.n673 B.n283 163.367
R1108 B.n673 B.n277 163.367
R1109 B.n681 B.n277 163.367
R1110 B.n681 B.n275 163.367
R1111 B.n685 B.n275 163.367
R1112 B.n685 B.n269 163.367
R1113 B.n694 B.n269 163.367
R1114 B.n694 B.n267 163.367
R1115 B.n698 B.n267 163.367
R1116 B.n698 B.n262 163.367
R1117 B.n707 B.n262 163.367
R1118 B.n707 B.n260 163.367
R1119 B.n711 B.n260 163.367
R1120 B.n711 B.n3 163.367
R1121 B.n931 B.n3 163.367
R1122 B.n927 B.n2 163.367
R1123 B.n927 B.n926 163.367
R1124 B.n926 B.n9 163.367
R1125 B.n922 B.n9 163.367
R1126 B.n922 B.n11 163.367
R1127 B.n918 B.n11 163.367
R1128 B.n918 B.n16 163.367
R1129 B.n914 B.n16 163.367
R1130 B.n914 B.n18 163.367
R1131 B.n910 B.n18 163.367
R1132 B.n910 B.n24 163.367
R1133 B.n906 B.n24 163.367
R1134 B.n906 B.n26 163.367
R1135 B.n902 B.n26 163.367
R1136 B.n902 B.n31 163.367
R1137 B.n898 B.n31 163.367
R1138 B.n898 B.n33 163.367
R1139 B.n895 B.n33 163.367
R1140 B.n895 B.n38 163.367
R1141 B.n891 B.n38 163.367
R1142 B.n891 B.n40 163.367
R1143 B.n887 B.n40 163.367
R1144 B.n887 B.n45 163.367
R1145 B.n883 B.n45 163.367
R1146 B.n883 B.n47 163.367
R1147 B.n879 B.n47 163.367
R1148 B.n879 B.n52 163.367
R1149 B.n875 B.n52 163.367
R1150 B.n875 B.n54 163.367
R1151 B.n871 B.n54 163.367
R1152 B.n871 B.n59 163.367
R1153 B.n867 B.n59 163.367
R1154 B.n867 B.n61 163.367
R1155 B.n863 B.n61 163.367
R1156 B.n863 B.n66 163.367
R1157 B.n859 B.n66 163.367
R1158 B.n859 B.n68 163.367
R1159 B.n855 B.n68 163.367
R1160 B.n855 B.n73 163.367
R1161 B.n851 B.n73 163.367
R1162 B.n851 B.n75 163.367
R1163 B.n847 B.n75 163.367
R1164 B.n847 B.n80 163.367
R1165 B.n843 B.n80 163.367
R1166 B.n843 B.n82 163.367
R1167 B.n839 B.n82 163.367
R1168 B.n839 B.n87 163.367
R1169 B.n835 B.n87 163.367
R1170 B.n835 B.n89 163.367
R1171 B.n831 B.n89 163.367
R1172 B.n831 B.n94 163.367
R1173 B.n827 B.n94 163.367
R1174 B.n827 B.n96 163.367
R1175 B.n823 B.n96 163.367
R1176 B.n823 B.n100 163.367
R1177 B.n819 B.n100 163.367
R1178 B.n819 B.n102 163.367
R1179 B.n815 B.n102 163.367
R1180 B.n815 B.n107 163.367
R1181 B.n811 B.n107 163.367
R1182 B.n811 B.n109 163.367
R1183 B.n807 B.n109 163.367
R1184 B.n807 B.n114 163.367
R1185 B.n803 B.n114 163.367
R1186 B.n146 B.t17 148.208
R1187 B.n472 B.t11 148.208
R1188 B.n149 B.t14 148.202
R1189 B.n399 B.t21 148.202
R1190 B.n525 B.n381 119.707
R1191 B.n802 B.n801 119.707
R1192 B.n150 B.n149 74.2793
R1193 B.n147 B.n146 74.2793
R1194 B.n473 B.n472 74.2793
R1195 B.n400 B.n399 74.2793
R1196 B.n147 B.t18 73.9293
R1197 B.n473 B.t10 73.9293
R1198 B.n150 B.t15 73.9235
R1199 B.n400 B.t20 73.9235
R1200 B.n118 B.n116 71.676
R1201 B.n153 B.n119 71.676
R1202 B.n157 B.n120 71.676
R1203 B.n161 B.n121 71.676
R1204 B.n165 B.n122 71.676
R1205 B.n169 B.n123 71.676
R1206 B.n173 B.n124 71.676
R1207 B.n177 B.n125 71.676
R1208 B.n181 B.n126 71.676
R1209 B.n185 B.n127 71.676
R1210 B.n189 B.n128 71.676
R1211 B.n193 B.n129 71.676
R1212 B.n198 B.n130 71.676
R1213 B.n202 B.n131 71.676
R1214 B.n206 B.n132 71.676
R1215 B.n210 B.n133 71.676
R1216 B.n214 B.n134 71.676
R1217 B.n218 B.n135 71.676
R1218 B.n222 B.n136 71.676
R1219 B.n226 B.n137 71.676
R1220 B.n230 B.n138 71.676
R1221 B.n234 B.n139 71.676
R1222 B.n238 B.n140 71.676
R1223 B.n242 B.n141 71.676
R1224 B.n246 B.n142 71.676
R1225 B.n250 B.n143 71.676
R1226 B.n254 B.n144 71.676
R1227 B.n145 B.n144 71.676
R1228 B.n253 B.n143 71.676
R1229 B.n249 B.n142 71.676
R1230 B.n245 B.n141 71.676
R1231 B.n241 B.n140 71.676
R1232 B.n237 B.n139 71.676
R1233 B.n233 B.n138 71.676
R1234 B.n229 B.n137 71.676
R1235 B.n225 B.n136 71.676
R1236 B.n221 B.n135 71.676
R1237 B.n217 B.n134 71.676
R1238 B.n213 B.n133 71.676
R1239 B.n209 B.n132 71.676
R1240 B.n205 B.n131 71.676
R1241 B.n201 B.n130 71.676
R1242 B.n197 B.n129 71.676
R1243 B.n192 B.n128 71.676
R1244 B.n188 B.n127 71.676
R1245 B.n184 B.n126 71.676
R1246 B.n180 B.n125 71.676
R1247 B.n176 B.n124 71.676
R1248 B.n172 B.n123 71.676
R1249 B.n168 B.n122 71.676
R1250 B.n164 B.n121 71.676
R1251 B.n160 B.n120 71.676
R1252 B.n156 B.n119 71.676
R1253 B.n152 B.n118 71.676
R1254 B.n411 B.n380 71.676
R1255 B.n417 B.n416 71.676
R1256 B.n420 B.n419 71.676
R1257 B.n425 B.n424 71.676
R1258 B.n428 B.n427 71.676
R1259 B.n433 B.n432 71.676
R1260 B.n436 B.n435 71.676
R1261 B.n441 B.n440 71.676
R1262 B.n444 B.n443 71.676
R1263 B.n449 B.n448 71.676
R1264 B.n452 B.n451 71.676
R1265 B.n458 B.n457 71.676
R1266 B.n461 B.n460 71.676
R1267 B.n466 B.n465 71.676
R1268 B.n469 B.n468 71.676
R1269 B.n477 B.n476 71.676
R1270 B.n480 B.n479 71.676
R1271 B.n485 B.n484 71.676
R1272 B.n488 B.n487 71.676
R1273 B.n493 B.n492 71.676
R1274 B.n496 B.n495 71.676
R1275 B.n501 B.n500 71.676
R1276 B.n504 B.n503 71.676
R1277 B.n509 B.n508 71.676
R1278 B.n512 B.n511 71.676
R1279 B.n517 B.n516 71.676
R1280 B.n520 B.n519 71.676
R1281 B.n412 B.n411 71.676
R1282 B.n418 B.n417 71.676
R1283 B.n419 B.n408 71.676
R1284 B.n426 B.n425 71.676
R1285 B.n427 B.n406 71.676
R1286 B.n434 B.n433 71.676
R1287 B.n435 B.n404 71.676
R1288 B.n442 B.n441 71.676
R1289 B.n443 B.n402 71.676
R1290 B.n450 B.n449 71.676
R1291 B.n451 B.n398 71.676
R1292 B.n459 B.n458 71.676
R1293 B.n460 B.n396 71.676
R1294 B.n467 B.n466 71.676
R1295 B.n468 B.n394 71.676
R1296 B.n478 B.n477 71.676
R1297 B.n479 B.n392 71.676
R1298 B.n486 B.n485 71.676
R1299 B.n487 B.n390 71.676
R1300 B.n494 B.n493 71.676
R1301 B.n495 B.n388 71.676
R1302 B.n502 B.n501 71.676
R1303 B.n503 B.n386 71.676
R1304 B.n510 B.n509 71.676
R1305 B.n511 B.n384 71.676
R1306 B.n518 B.n517 71.676
R1307 B.n519 B.n382 71.676
R1308 B.n932 B.n931 71.676
R1309 B.n932 B.n2 71.676
R1310 B.n525 B.n377 68.4047
R1311 B.n531 B.n377 68.4047
R1312 B.n531 B.n373 68.4047
R1313 B.n537 B.n373 68.4047
R1314 B.n537 B.n369 68.4047
R1315 B.n543 B.n369 68.4047
R1316 B.n543 B.n365 68.4047
R1317 B.n549 B.n365 68.4047
R1318 B.n549 B.t9 68.4047
R1319 B.n555 B.t9 68.4047
R1320 B.n555 B.n358 68.4047
R1321 B.n561 B.n358 68.4047
R1322 B.n561 B.n354 68.4047
R1323 B.n567 B.n354 68.4047
R1324 B.n567 B.n350 68.4047
R1325 B.n573 B.n350 68.4047
R1326 B.n573 B.n346 68.4047
R1327 B.n579 B.n346 68.4047
R1328 B.n579 B.n342 68.4047
R1329 B.n585 B.n342 68.4047
R1330 B.n585 B.n337 68.4047
R1331 B.n591 B.n337 68.4047
R1332 B.n591 B.n338 68.4047
R1333 B.n597 B.n330 68.4047
R1334 B.n603 B.n330 68.4047
R1335 B.n603 B.n326 68.4047
R1336 B.n609 B.n326 68.4047
R1337 B.n609 B.n322 68.4047
R1338 B.n615 B.n322 68.4047
R1339 B.n615 B.n318 68.4047
R1340 B.n621 B.n318 68.4047
R1341 B.n621 B.n314 68.4047
R1342 B.n627 B.n314 68.4047
R1343 B.n633 B.n310 68.4047
R1344 B.n633 B.n306 68.4047
R1345 B.n639 B.n306 68.4047
R1346 B.n639 B.n302 68.4047
R1347 B.n645 B.n302 68.4047
R1348 B.n645 B.n298 68.4047
R1349 B.n651 B.n298 68.4047
R1350 B.n651 B.n294 68.4047
R1351 B.n657 B.n294 68.4047
R1352 B.n657 B.n290 68.4047
R1353 B.t6 B.n290 68.4047
R1354 B.t6 B.n286 68.4047
R1355 B.n668 B.n286 68.4047
R1356 B.n668 B.n282 68.4047
R1357 B.n674 B.n282 68.4047
R1358 B.n674 B.n278 68.4047
R1359 B.n680 B.n278 68.4047
R1360 B.n680 B.n274 68.4047
R1361 B.n686 B.n274 68.4047
R1362 B.n686 B.n270 68.4047
R1363 B.n693 B.n270 68.4047
R1364 B.n693 B.n692 68.4047
R1365 B.n699 B.n263 68.4047
R1366 B.n706 B.n263 68.4047
R1367 B.n706 B.n259 68.4047
R1368 B.n712 B.n259 68.4047
R1369 B.n712 B.n4 68.4047
R1370 B.n930 B.n4 68.4047
R1371 B.n930 B.n929 68.4047
R1372 B.n929 B.n928 68.4047
R1373 B.n928 B.n8 68.4047
R1374 B.n12 B.n8 68.4047
R1375 B.n921 B.n12 68.4047
R1376 B.n921 B.n920 68.4047
R1377 B.n920 B.n919 68.4047
R1378 B.n913 B.n19 68.4047
R1379 B.n913 B.n912 68.4047
R1380 B.n912 B.n911 68.4047
R1381 B.n911 B.n23 68.4047
R1382 B.n905 B.n23 68.4047
R1383 B.n905 B.n904 68.4047
R1384 B.n904 B.n903 68.4047
R1385 B.n903 B.n30 68.4047
R1386 B.n897 B.n30 68.4047
R1387 B.n897 B.n896 68.4047
R1388 B.n896 B.t2 68.4047
R1389 B.t2 B.n37 68.4047
R1390 B.n890 B.n37 68.4047
R1391 B.n890 B.n889 68.4047
R1392 B.n889 B.n888 68.4047
R1393 B.n888 B.n44 68.4047
R1394 B.n882 B.n44 68.4047
R1395 B.n882 B.n881 68.4047
R1396 B.n881 B.n880 68.4047
R1397 B.n880 B.n51 68.4047
R1398 B.n874 B.n51 68.4047
R1399 B.n874 B.n873 68.4047
R1400 B.n872 B.n58 68.4047
R1401 B.n866 B.n58 68.4047
R1402 B.n866 B.n865 68.4047
R1403 B.n865 B.n864 68.4047
R1404 B.n864 B.n65 68.4047
R1405 B.n858 B.n65 68.4047
R1406 B.n858 B.n857 68.4047
R1407 B.n857 B.n856 68.4047
R1408 B.n856 B.n72 68.4047
R1409 B.n850 B.n72 68.4047
R1410 B.n849 B.n848 68.4047
R1411 B.n848 B.n79 68.4047
R1412 B.n842 B.n79 68.4047
R1413 B.n842 B.n841 68.4047
R1414 B.n841 B.n840 68.4047
R1415 B.n840 B.n86 68.4047
R1416 B.n834 B.n86 68.4047
R1417 B.n834 B.n833 68.4047
R1418 B.n833 B.n832 68.4047
R1419 B.n832 B.n93 68.4047
R1420 B.n826 B.n93 68.4047
R1421 B.n826 B.n825 68.4047
R1422 B.n825 B.n824 68.4047
R1423 B.n824 B.t13 68.4047
R1424 B.n818 B.t13 68.4047
R1425 B.n818 B.n817 68.4047
R1426 B.n817 B.n816 68.4047
R1427 B.n816 B.n106 68.4047
R1428 B.n810 B.n106 68.4047
R1429 B.n810 B.n809 68.4047
R1430 B.n809 B.n808 68.4047
R1431 B.n808 B.n113 68.4047
R1432 B.n802 B.n113 68.4047
R1433 B.n195 B.n150 59.5399
R1434 B.n148 B.n147 59.5399
R1435 B.n474 B.n473 59.5399
R1436 B.n455 B.n400 59.5399
R1437 B.n627 B.t1 50.2977
R1438 B.n699 B.t5 50.2977
R1439 B.n919 B.t7 50.2977
R1440 B.t0 B.n872 50.2977
R1441 B.n597 B.t4 36.2145
R1442 B.n850 B.t3 36.2145
R1443 B.n527 B.n379 34.4981
R1444 B.n523 B.n522 34.4981
R1445 B.n799 B.n798 34.4981
R1446 B.n804 B.n115 34.4981
R1447 B.n338 B.t4 32.1907
R1448 B.t3 B.n849 32.1907
R1449 B.t1 B.n310 18.1075
R1450 B.n692 B.t5 18.1075
R1451 B.n19 B.t7 18.1075
R1452 B.n873 B.t0 18.1075
R1453 B B.n933 18.0485
R1454 B.n528 B.n527 10.6151
R1455 B.n529 B.n528 10.6151
R1456 B.n529 B.n371 10.6151
R1457 B.n539 B.n371 10.6151
R1458 B.n540 B.n539 10.6151
R1459 B.n541 B.n540 10.6151
R1460 B.n541 B.n363 10.6151
R1461 B.n551 B.n363 10.6151
R1462 B.n552 B.n551 10.6151
R1463 B.n553 B.n552 10.6151
R1464 B.n553 B.n356 10.6151
R1465 B.n563 B.n356 10.6151
R1466 B.n564 B.n563 10.6151
R1467 B.n565 B.n564 10.6151
R1468 B.n565 B.n348 10.6151
R1469 B.n575 B.n348 10.6151
R1470 B.n576 B.n575 10.6151
R1471 B.n577 B.n576 10.6151
R1472 B.n577 B.n340 10.6151
R1473 B.n587 B.n340 10.6151
R1474 B.n588 B.n587 10.6151
R1475 B.n589 B.n588 10.6151
R1476 B.n589 B.n332 10.6151
R1477 B.n599 B.n332 10.6151
R1478 B.n600 B.n599 10.6151
R1479 B.n601 B.n600 10.6151
R1480 B.n601 B.n324 10.6151
R1481 B.n611 B.n324 10.6151
R1482 B.n612 B.n611 10.6151
R1483 B.n613 B.n612 10.6151
R1484 B.n613 B.n316 10.6151
R1485 B.n623 B.n316 10.6151
R1486 B.n624 B.n623 10.6151
R1487 B.n625 B.n624 10.6151
R1488 B.n625 B.n308 10.6151
R1489 B.n635 B.n308 10.6151
R1490 B.n636 B.n635 10.6151
R1491 B.n637 B.n636 10.6151
R1492 B.n637 B.n300 10.6151
R1493 B.n647 B.n300 10.6151
R1494 B.n648 B.n647 10.6151
R1495 B.n649 B.n648 10.6151
R1496 B.n649 B.n292 10.6151
R1497 B.n659 B.n292 10.6151
R1498 B.n660 B.n659 10.6151
R1499 B.n661 B.n660 10.6151
R1500 B.n661 B.n284 10.6151
R1501 B.n670 B.n284 10.6151
R1502 B.n671 B.n670 10.6151
R1503 B.n672 B.n671 10.6151
R1504 B.n672 B.n276 10.6151
R1505 B.n682 B.n276 10.6151
R1506 B.n683 B.n682 10.6151
R1507 B.n684 B.n683 10.6151
R1508 B.n684 B.n268 10.6151
R1509 B.n695 B.n268 10.6151
R1510 B.n696 B.n695 10.6151
R1511 B.n697 B.n696 10.6151
R1512 B.n697 B.n261 10.6151
R1513 B.n708 B.n261 10.6151
R1514 B.n709 B.n708 10.6151
R1515 B.n710 B.n709 10.6151
R1516 B.n710 B.n0 10.6151
R1517 B.n413 B.n379 10.6151
R1518 B.n414 B.n413 10.6151
R1519 B.n415 B.n414 10.6151
R1520 B.n415 B.n409 10.6151
R1521 B.n421 B.n409 10.6151
R1522 B.n422 B.n421 10.6151
R1523 B.n423 B.n422 10.6151
R1524 B.n423 B.n407 10.6151
R1525 B.n429 B.n407 10.6151
R1526 B.n430 B.n429 10.6151
R1527 B.n431 B.n430 10.6151
R1528 B.n431 B.n405 10.6151
R1529 B.n437 B.n405 10.6151
R1530 B.n438 B.n437 10.6151
R1531 B.n439 B.n438 10.6151
R1532 B.n439 B.n403 10.6151
R1533 B.n445 B.n403 10.6151
R1534 B.n446 B.n445 10.6151
R1535 B.n447 B.n446 10.6151
R1536 B.n447 B.n401 10.6151
R1537 B.n453 B.n401 10.6151
R1538 B.n454 B.n453 10.6151
R1539 B.n456 B.n397 10.6151
R1540 B.n462 B.n397 10.6151
R1541 B.n463 B.n462 10.6151
R1542 B.n464 B.n463 10.6151
R1543 B.n464 B.n395 10.6151
R1544 B.n470 B.n395 10.6151
R1545 B.n471 B.n470 10.6151
R1546 B.n475 B.n471 10.6151
R1547 B.n481 B.n393 10.6151
R1548 B.n482 B.n481 10.6151
R1549 B.n483 B.n482 10.6151
R1550 B.n483 B.n391 10.6151
R1551 B.n489 B.n391 10.6151
R1552 B.n490 B.n489 10.6151
R1553 B.n491 B.n490 10.6151
R1554 B.n491 B.n389 10.6151
R1555 B.n497 B.n389 10.6151
R1556 B.n498 B.n497 10.6151
R1557 B.n499 B.n498 10.6151
R1558 B.n499 B.n387 10.6151
R1559 B.n505 B.n387 10.6151
R1560 B.n506 B.n505 10.6151
R1561 B.n507 B.n506 10.6151
R1562 B.n507 B.n385 10.6151
R1563 B.n513 B.n385 10.6151
R1564 B.n514 B.n513 10.6151
R1565 B.n515 B.n514 10.6151
R1566 B.n515 B.n383 10.6151
R1567 B.n521 B.n383 10.6151
R1568 B.n522 B.n521 10.6151
R1569 B.n523 B.n375 10.6151
R1570 B.n533 B.n375 10.6151
R1571 B.n534 B.n533 10.6151
R1572 B.n535 B.n534 10.6151
R1573 B.n535 B.n367 10.6151
R1574 B.n545 B.n367 10.6151
R1575 B.n546 B.n545 10.6151
R1576 B.n547 B.n546 10.6151
R1577 B.n547 B.n360 10.6151
R1578 B.n557 B.n360 10.6151
R1579 B.n558 B.n557 10.6151
R1580 B.n559 B.n558 10.6151
R1581 B.n559 B.n352 10.6151
R1582 B.n569 B.n352 10.6151
R1583 B.n570 B.n569 10.6151
R1584 B.n571 B.n570 10.6151
R1585 B.n571 B.n344 10.6151
R1586 B.n581 B.n344 10.6151
R1587 B.n582 B.n581 10.6151
R1588 B.n583 B.n582 10.6151
R1589 B.n583 B.n335 10.6151
R1590 B.n593 B.n335 10.6151
R1591 B.n594 B.n593 10.6151
R1592 B.n595 B.n594 10.6151
R1593 B.n595 B.n328 10.6151
R1594 B.n605 B.n328 10.6151
R1595 B.n606 B.n605 10.6151
R1596 B.n607 B.n606 10.6151
R1597 B.n607 B.n320 10.6151
R1598 B.n617 B.n320 10.6151
R1599 B.n618 B.n617 10.6151
R1600 B.n619 B.n618 10.6151
R1601 B.n619 B.n312 10.6151
R1602 B.n629 B.n312 10.6151
R1603 B.n630 B.n629 10.6151
R1604 B.n631 B.n630 10.6151
R1605 B.n631 B.n304 10.6151
R1606 B.n641 B.n304 10.6151
R1607 B.n642 B.n641 10.6151
R1608 B.n643 B.n642 10.6151
R1609 B.n643 B.n296 10.6151
R1610 B.n653 B.n296 10.6151
R1611 B.n654 B.n653 10.6151
R1612 B.n655 B.n654 10.6151
R1613 B.n655 B.n288 10.6151
R1614 B.n664 B.n288 10.6151
R1615 B.n665 B.n664 10.6151
R1616 B.n666 B.n665 10.6151
R1617 B.n666 B.n280 10.6151
R1618 B.n676 B.n280 10.6151
R1619 B.n677 B.n676 10.6151
R1620 B.n678 B.n677 10.6151
R1621 B.n678 B.n272 10.6151
R1622 B.n688 B.n272 10.6151
R1623 B.n689 B.n688 10.6151
R1624 B.n690 B.n689 10.6151
R1625 B.n690 B.n265 10.6151
R1626 B.n701 B.n265 10.6151
R1627 B.n702 B.n701 10.6151
R1628 B.n704 B.n702 10.6151
R1629 B.n704 B.n703 10.6151
R1630 B.n703 B.n257 10.6151
R1631 B.n715 B.n257 10.6151
R1632 B.n716 B.n715 10.6151
R1633 B.n717 B.n716 10.6151
R1634 B.n718 B.n717 10.6151
R1635 B.n719 B.n718 10.6151
R1636 B.n722 B.n719 10.6151
R1637 B.n723 B.n722 10.6151
R1638 B.n724 B.n723 10.6151
R1639 B.n725 B.n724 10.6151
R1640 B.n727 B.n725 10.6151
R1641 B.n728 B.n727 10.6151
R1642 B.n729 B.n728 10.6151
R1643 B.n730 B.n729 10.6151
R1644 B.n732 B.n730 10.6151
R1645 B.n733 B.n732 10.6151
R1646 B.n734 B.n733 10.6151
R1647 B.n735 B.n734 10.6151
R1648 B.n737 B.n735 10.6151
R1649 B.n738 B.n737 10.6151
R1650 B.n739 B.n738 10.6151
R1651 B.n740 B.n739 10.6151
R1652 B.n742 B.n740 10.6151
R1653 B.n743 B.n742 10.6151
R1654 B.n744 B.n743 10.6151
R1655 B.n745 B.n744 10.6151
R1656 B.n747 B.n745 10.6151
R1657 B.n748 B.n747 10.6151
R1658 B.n749 B.n748 10.6151
R1659 B.n750 B.n749 10.6151
R1660 B.n752 B.n750 10.6151
R1661 B.n753 B.n752 10.6151
R1662 B.n754 B.n753 10.6151
R1663 B.n755 B.n754 10.6151
R1664 B.n757 B.n755 10.6151
R1665 B.n758 B.n757 10.6151
R1666 B.n759 B.n758 10.6151
R1667 B.n760 B.n759 10.6151
R1668 B.n762 B.n760 10.6151
R1669 B.n763 B.n762 10.6151
R1670 B.n764 B.n763 10.6151
R1671 B.n765 B.n764 10.6151
R1672 B.n767 B.n765 10.6151
R1673 B.n768 B.n767 10.6151
R1674 B.n769 B.n768 10.6151
R1675 B.n770 B.n769 10.6151
R1676 B.n772 B.n770 10.6151
R1677 B.n773 B.n772 10.6151
R1678 B.n774 B.n773 10.6151
R1679 B.n775 B.n774 10.6151
R1680 B.n777 B.n775 10.6151
R1681 B.n778 B.n777 10.6151
R1682 B.n779 B.n778 10.6151
R1683 B.n780 B.n779 10.6151
R1684 B.n782 B.n780 10.6151
R1685 B.n783 B.n782 10.6151
R1686 B.n784 B.n783 10.6151
R1687 B.n785 B.n784 10.6151
R1688 B.n787 B.n785 10.6151
R1689 B.n788 B.n787 10.6151
R1690 B.n789 B.n788 10.6151
R1691 B.n790 B.n789 10.6151
R1692 B.n792 B.n790 10.6151
R1693 B.n793 B.n792 10.6151
R1694 B.n794 B.n793 10.6151
R1695 B.n795 B.n794 10.6151
R1696 B.n797 B.n795 10.6151
R1697 B.n798 B.n797 10.6151
R1698 B.n925 B.n1 10.6151
R1699 B.n925 B.n924 10.6151
R1700 B.n924 B.n923 10.6151
R1701 B.n923 B.n10 10.6151
R1702 B.n917 B.n10 10.6151
R1703 B.n917 B.n916 10.6151
R1704 B.n916 B.n915 10.6151
R1705 B.n915 B.n17 10.6151
R1706 B.n909 B.n17 10.6151
R1707 B.n909 B.n908 10.6151
R1708 B.n908 B.n907 10.6151
R1709 B.n907 B.n25 10.6151
R1710 B.n901 B.n25 10.6151
R1711 B.n901 B.n900 10.6151
R1712 B.n900 B.n899 10.6151
R1713 B.n899 B.n32 10.6151
R1714 B.n894 B.n32 10.6151
R1715 B.n894 B.n893 10.6151
R1716 B.n893 B.n892 10.6151
R1717 B.n892 B.n39 10.6151
R1718 B.n886 B.n39 10.6151
R1719 B.n886 B.n885 10.6151
R1720 B.n885 B.n884 10.6151
R1721 B.n884 B.n46 10.6151
R1722 B.n878 B.n46 10.6151
R1723 B.n878 B.n877 10.6151
R1724 B.n877 B.n876 10.6151
R1725 B.n876 B.n53 10.6151
R1726 B.n870 B.n53 10.6151
R1727 B.n870 B.n869 10.6151
R1728 B.n869 B.n868 10.6151
R1729 B.n868 B.n60 10.6151
R1730 B.n862 B.n60 10.6151
R1731 B.n862 B.n861 10.6151
R1732 B.n861 B.n860 10.6151
R1733 B.n860 B.n67 10.6151
R1734 B.n854 B.n67 10.6151
R1735 B.n854 B.n853 10.6151
R1736 B.n853 B.n852 10.6151
R1737 B.n852 B.n74 10.6151
R1738 B.n846 B.n74 10.6151
R1739 B.n846 B.n845 10.6151
R1740 B.n845 B.n844 10.6151
R1741 B.n844 B.n81 10.6151
R1742 B.n838 B.n81 10.6151
R1743 B.n838 B.n837 10.6151
R1744 B.n837 B.n836 10.6151
R1745 B.n836 B.n88 10.6151
R1746 B.n830 B.n88 10.6151
R1747 B.n830 B.n829 10.6151
R1748 B.n829 B.n828 10.6151
R1749 B.n828 B.n95 10.6151
R1750 B.n822 B.n95 10.6151
R1751 B.n822 B.n821 10.6151
R1752 B.n821 B.n820 10.6151
R1753 B.n820 B.n101 10.6151
R1754 B.n814 B.n101 10.6151
R1755 B.n814 B.n813 10.6151
R1756 B.n813 B.n812 10.6151
R1757 B.n812 B.n108 10.6151
R1758 B.n806 B.n108 10.6151
R1759 B.n806 B.n805 10.6151
R1760 B.n805 B.n804 10.6151
R1761 B.n151 B.n115 10.6151
R1762 B.n154 B.n151 10.6151
R1763 B.n155 B.n154 10.6151
R1764 B.n158 B.n155 10.6151
R1765 B.n159 B.n158 10.6151
R1766 B.n162 B.n159 10.6151
R1767 B.n163 B.n162 10.6151
R1768 B.n166 B.n163 10.6151
R1769 B.n167 B.n166 10.6151
R1770 B.n170 B.n167 10.6151
R1771 B.n171 B.n170 10.6151
R1772 B.n174 B.n171 10.6151
R1773 B.n175 B.n174 10.6151
R1774 B.n178 B.n175 10.6151
R1775 B.n179 B.n178 10.6151
R1776 B.n182 B.n179 10.6151
R1777 B.n183 B.n182 10.6151
R1778 B.n186 B.n183 10.6151
R1779 B.n187 B.n186 10.6151
R1780 B.n190 B.n187 10.6151
R1781 B.n191 B.n190 10.6151
R1782 B.n194 B.n191 10.6151
R1783 B.n199 B.n196 10.6151
R1784 B.n200 B.n199 10.6151
R1785 B.n203 B.n200 10.6151
R1786 B.n204 B.n203 10.6151
R1787 B.n207 B.n204 10.6151
R1788 B.n208 B.n207 10.6151
R1789 B.n211 B.n208 10.6151
R1790 B.n212 B.n211 10.6151
R1791 B.n216 B.n215 10.6151
R1792 B.n219 B.n216 10.6151
R1793 B.n220 B.n219 10.6151
R1794 B.n223 B.n220 10.6151
R1795 B.n224 B.n223 10.6151
R1796 B.n227 B.n224 10.6151
R1797 B.n228 B.n227 10.6151
R1798 B.n231 B.n228 10.6151
R1799 B.n232 B.n231 10.6151
R1800 B.n235 B.n232 10.6151
R1801 B.n236 B.n235 10.6151
R1802 B.n239 B.n236 10.6151
R1803 B.n240 B.n239 10.6151
R1804 B.n243 B.n240 10.6151
R1805 B.n244 B.n243 10.6151
R1806 B.n247 B.n244 10.6151
R1807 B.n248 B.n247 10.6151
R1808 B.n251 B.n248 10.6151
R1809 B.n252 B.n251 10.6151
R1810 B.n255 B.n252 10.6151
R1811 B.n256 B.n255 10.6151
R1812 B.n799 B.n256 10.6151
R1813 B.n933 B.n0 8.11757
R1814 B.n933 B.n1 8.11757
R1815 B.n456 B.n455 6.5566
R1816 B.n475 B.n474 6.5566
R1817 B.n196 B.n195 6.5566
R1818 B.n212 B.n148 6.5566
R1819 B.n455 B.n454 4.05904
R1820 B.n474 B.n393 4.05904
R1821 B.n195 B.n194 4.05904
R1822 B.n215 B.n148 4.05904
R1823 VN.n68 VN.n67 161.3
R1824 VN.n66 VN.n36 161.3
R1825 VN.n65 VN.n64 161.3
R1826 VN.n63 VN.n37 161.3
R1827 VN.n62 VN.n61 161.3
R1828 VN.n60 VN.n38 161.3
R1829 VN.n59 VN.n58 161.3
R1830 VN.n57 VN.n39 161.3
R1831 VN.n56 VN.n55 161.3
R1832 VN.n54 VN.n40 161.3
R1833 VN.n53 VN.n52 161.3
R1834 VN.n51 VN.n42 161.3
R1835 VN.n50 VN.n49 161.3
R1836 VN.n48 VN.n43 161.3
R1837 VN.n47 VN.n46 161.3
R1838 VN.n33 VN.n32 161.3
R1839 VN.n31 VN.n1 161.3
R1840 VN.n30 VN.n29 161.3
R1841 VN.n28 VN.n2 161.3
R1842 VN.n27 VN.n26 161.3
R1843 VN.n25 VN.n3 161.3
R1844 VN.n24 VN.n23 161.3
R1845 VN.n22 VN.n4 161.3
R1846 VN.n21 VN.n20 161.3
R1847 VN.n18 VN.n5 161.3
R1848 VN.n17 VN.n16 161.3
R1849 VN.n15 VN.n6 161.3
R1850 VN.n14 VN.n13 161.3
R1851 VN.n12 VN.n7 161.3
R1852 VN.n11 VN.n10 161.3
R1853 VN.n34 VN.n0 78.1956
R1854 VN.n69 VN.n35 78.1956
R1855 VN.n9 VN.t7 72.7366
R1856 VN.n45 VN.t5 72.7366
R1857 VN.n26 VN.n2 56.5617
R1858 VN.n61 VN.n37 56.5617
R1859 VN.n9 VN.n8 54.4907
R1860 VN.n45 VN.n44 54.4907
R1861 VN VN.n69 50.589
R1862 VN.n13 VN.n6 40.577
R1863 VN.n17 VN.n6 40.577
R1864 VN.n49 VN.n42 40.577
R1865 VN.n53 VN.n42 40.577
R1866 VN.n8 VN.t3 38.9736
R1867 VN.n19 VN.t0 38.9736
R1868 VN.n0 VN.t4 38.9736
R1869 VN.n44 VN.t2 38.9736
R1870 VN.n41 VN.t6 38.9736
R1871 VN.n35 VN.t1 38.9736
R1872 VN.n12 VN.n11 24.5923
R1873 VN.n13 VN.n12 24.5923
R1874 VN.n18 VN.n17 24.5923
R1875 VN.n20 VN.n18 24.5923
R1876 VN.n24 VN.n4 24.5923
R1877 VN.n25 VN.n24 24.5923
R1878 VN.n26 VN.n25 24.5923
R1879 VN.n30 VN.n2 24.5923
R1880 VN.n31 VN.n30 24.5923
R1881 VN.n32 VN.n31 24.5923
R1882 VN.n49 VN.n48 24.5923
R1883 VN.n48 VN.n47 24.5923
R1884 VN.n61 VN.n60 24.5923
R1885 VN.n60 VN.n59 24.5923
R1886 VN.n59 VN.n39 24.5923
R1887 VN.n55 VN.n54 24.5923
R1888 VN.n54 VN.n53 24.5923
R1889 VN.n67 VN.n66 24.5923
R1890 VN.n66 VN.n65 24.5923
R1891 VN.n65 VN.n37 24.5923
R1892 VN.n11 VN.n8 20.4117
R1893 VN.n20 VN.n19 20.4117
R1894 VN.n47 VN.n44 20.4117
R1895 VN.n55 VN.n41 20.4117
R1896 VN.n32 VN.n0 12.0505
R1897 VN.n67 VN.n35 12.0505
R1898 VN.n19 VN.n4 4.18111
R1899 VN.n41 VN.n39 4.18111
R1900 VN.n10 VN.n9 3.0794
R1901 VN.n46 VN.n45 3.0794
R1902 VN.n69 VN.n68 0.354861
R1903 VN.n34 VN.n33 0.354861
R1904 VN VN.n34 0.267071
R1905 VN.n68 VN.n36 0.189894
R1906 VN.n64 VN.n36 0.189894
R1907 VN.n64 VN.n63 0.189894
R1908 VN.n63 VN.n62 0.189894
R1909 VN.n62 VN.n38 0.189894
R1910 VN.n58 VN.n38 0.189894
R1911 VN.n58 VN.n57 0.189894
R1912 VN.n57 VN.n56 0.189894
R1913 VN.n56 VN.n40 0.189894
R1914 VN.n52 VN.n40 0.189894
R1915 VN.n52 VN.n51 0.189894
R1916 VN.n51 VN.n50 0.189894
R1917 VN.n50 VN.n43 0.189894
R1918 VN.n46 VN.n43 0.189894
R1919 VN.n10 VN.n7 0.189894
R1920 VN.n14 VN.n7 0.189894
R1921 VN.n15 VN.n14 0.189894
R1922 VN.n16 VN.n15 0.189894
R1923 VN.n16 VN.n5 0.189894
R1924 VN.n21 VN.n5 0.189894
R1925 VN.n22 VN.n21 0.189894
R1926 VN.n23 VN.n22 0.189894
R1927 VN.n23 VN.n3 0.189894
R1928 VN.n27 VN.n3 0.189894
R1929 VN.n28 VN.n27 0.189894
R1930 VN.n29 VN.n28 0.189894
R1931 VN.n29 VN.n1 0.189894
R1932 VN.n33 VN.n1 0.189894
R1933 VDD2.n2 VDD2.n1 69.8532
R1934 VDD2.n2 VDD2.n0 69.8532
R1935 VDD2 VDD2.n5 69.8504
R1936 VDD2.n4 VDD2.n3 68.2579
R1937 VDD2.n4 VDD2.n2 43.4524
R1938 VDD2.n5 VDD2.t5 3.49873
R1939 VDD2.n5 VDD2.t2 3.49873
R1940 VDD2.n3 VDD2.t6 3.49873
R1941 VDD2.n3 VDD2.t1 3.49873
R1942 VDD2.n1 VDD2.t7 3.49873
R1943 VDD2.n1 VDD2.t3 3.49873
R1944 VDD2.n0 VDD2.t0 3.49873
R1945 VDD2.n0 VDD2.t4 3.49873
R1946 VDD2 VDD2.n4 1.70955
C0 VDD2 VDD1 2.24472f
C1 VN VDD1 0.153825f
C2 VTAIL VDD1 6.60056f
C3 VDD2 VN 4.56216f
C4 VTAIL VDD2 6.66101f
C5 VTAIL VN 5.79616f
C6 VDD1 VP 5.0224f
C7 VDD2 VP 0.61591f
C8 VN VP 7.58166f
C9 VTAIL VP 5.81027f
C10 VDD2 B 5.877414f
C11 VDD1 B 6.41388f
C12 VTAIL B 6.770923f
C13 VN B 18.32963f
C14 VP B 16.951342f
C15 VDD2.t0 B 0.129369f
C16 VDD2.t4 B 0.129369f
C17 VDD2.n0 B 1.0873f
C18 VDD2.t7 B 0.129369f
C19 VDD2.t3 B 0.129369f
C20 VDD2.n1 B 1.0873f
C21 VDD2.n2 B 3.93174f
C22 VDD2.t6 B 0.129369f
C23 VDD2.t1 B 0.129369f
C24 VDD2.n3 B 1.07127f
C25 VDD2.n4 B 3.20735f
C26 VDD2.t5 B 0.129369f
C27 VDD2.t2 B 0.129369f
C28 VDD2.n5 B 1.08725f
C29 VN.t4 B 1.11985f
C30 VN.n0 B 0.500977f
C31 VN.n1 B 0.021434f
C32 VN.n2 B 0.026413f
C33 VN.n3 B 0.021434f
C34 VN.n4 B 0.023461f
C35 VN.n5 B 0.021434f
C36 VN.n6 B 0.017311f
C37 VN.n7 B 0.021434f
C38 VN.t3 B 1.11985f
C39 VN.n8 B 0.496858f
C40 VN.t7 B 1.38769f
C41 VN.n9 B 0.47103f
C42 VN.n10 B 0.263845f
C43 VN.n11 B 0.036411f
C44 VN.n12 B 0.039747f
C45 VN.n13 B 0.042375f
C46 VN.n14 B 0.021434f
C47 VN.n15 B 0.021434f
C48 VN.n16 B 0.021434f
C49 VN.n17 B 0.042375f
C50 VN.n18 B 0.039747f
C51 VN.t0 B 1.11985f
C52 VN.n19 B 0.416266f
C53 VN.n20 B 0.036411f
C54 VN.n21 B 0.021434f
C55 VN.n22 B 0.021434f
C56 VN.n23 B 0.021434f
C57 VN.n24 B 0.039747f
C58 VN.n25 B 0.039747f
C59 VN.n26 B 0.035901f
C60 VN.n27 B 0.021434f
C61 VN.n28 B 0.021434f
C62 VN.n29 B 0.021434f
C63 VN.n30 B 0.039747f
C64 VN.n31 B 0.039747f
C65 VN.n32 B 0.02974f
C66 VN.n33 B 0.034588f
C67 VN.n34 B 0.055923f
C68 VN.t1 B 1.11985f
C69 VN.n35 B 0.500977f
C70 VN.n36 B 0.021434f
C71 VN.n37 B 0.026413f
C72 VN.n38 B 0.021434f
C73 VN.n39 B 0.023461f
C74 VN.n40 B 0.021434f
C75 VN.t6 B 1.11985f
C76 VN.n41 B 0.416266f
C77 VN.n42 B 0.017311f
C78 VN.n43 B 0.021434f
C79 VN.t2 B 1.11985f
C80 VN.n44 B 0.496858f
C81 VN.t5 B 1.38769f
C82 VN.n45 B 0.47103f
C83 VN.n46 B 0.263845f
C84 VN.n47 B 0.036411f
C85 VN.n48 B 0.039747f
C86 VN.n49 B 0.042375f
C87 VN.n50 B 0.021434f
C88 VN.n51 B 0.021434f
C89 VN.n52 B 0.021434f
C90 VN.n53 B 0.042375f
C91 VN.n54 B 0.039747f
C92 VN.n55 B 0.036411f
C93 VN.n56 B 0.021434f
C94 VN.n57 B 0.021434f
C95 VN.n58 B 0.021434f
C96 VN.n59 B 0.039747f
C97 VN.n60 B 0.039747f
C98 VN.n61 B 0.035901f
C99 VN.n62 B 0.021434f
C100 VN.n63 B 0.021434f
C101 VN.n64 B 0.021434f
C102 VN.n65 B 0.039747f
C103 VN.n66 B 0.039747f
C104 VN.n67 B 0.02974f
C105 VN.n68 B 0.034588f
C106 VN.n69 B 1.24767f
C107 VDD1.t4 B 0.131205f
C108 VDD1.t7 B 0.131205f
C109 VDD1.n0 B 1.10412f
C110 VDD1.t2 B 0.131205f
C111 VDD1.t3 B 0.131205f
C112 VDD1.n1 B 1.10273f
C113 VDD1.t0 B 0.131205f
C114 VDD1.t5 B 0.131205f
C115 VDD1.n2 B 1.10273f
C116 VDD1.n3 B 4.0483f
C117 VDD1.t6 B 0.131205f
C118 VDD1.t1 B 0.131205f
C119 VDD1.n4 B 1.08647f
C120 VDD1.n5 B 3.2895f
C121 VTAIL.t2 B 0.112003f
C122 VTAIL.t0 B 0.112003f
C123 VTAIL.n0 B 0.863696f
C124 VTAIL.n1 B 0.502821f
C125 VTAIL.t7 B 1.10201f
C126 VTAIL.n2 B 0.603181f
C127 VTAIL.t15 B 1.10201f
C128 VTAIL.n3 B 0.603181f
C129 VTAIL.t14 B 0.112003f
C130 VTAIL.t12 B 0.112003f
C131 VTAIL.n4 B 0.863696f
C132 VTAIL.n5 B 0.764539f
C133 VTAIL.t8 B 1.10201f
C134 VTAIL.n6 B 1.56555f
C135 VTAIL.t4 B 1.10202f
C136 VTAIL.n7 B 1.56555f
C137 VTAIL.t1 B 0.112003f
C138 VTAIL.t6 B 0.112003f
C139 VTAIL.n8 B 0.863701f
C140 VTAIL.n9 B 0.764534f
C141 VTAIL.t5 B 1.10202f
C142 VTAIL.n10 B 0.603177f
C143 VTAIL.t9 B 1.10202f
C144 VTAIL.n11 B 0.603177f
C145 VTAIL.t13 B 0.112003f
C146 VTAIL.t10 B 0.112003f
C147 VTAIL.n12 B 0.863701f
C148 VTAIL.n13 B 0.764534f
C149 VTAIL.t11 B 1.10201f
C150 VTAIL.n14 B 1.56555f
C151 VTAIL.t3 B 1.10201f
C152 VTAIL.n15 B 1.56086f
C153 VP.t2 B 1.14666f
C154 VP.n0 B 0.512969f
C155 VP.n1 B 0.021947f
C156 VP.n2 B 0.027045f
C157 VP.n3 B 0.021947f
C158 VP.n4 B 0.024022f
C159 VP.n5 B 0.021947f
C160 VP.n6 B 0.017726f
C161 VP.n7 B 0.021947f
C162 VP.t4 B 1.14666f
C163 VP.n8 B 0.42623f
C164 VP.n9 B 0.021947f
C165 VP.n10 B 0.036761f
C166 VP.n11 B 0.021947f
C167 VP.n12 B 0.030451f
C168 VP.t6 B 1.14666f
C169 VP.n13 B 0.512969f
C170 VP.n14 B 0.021947f
C171 VP.n15 B 0.027045f
C172 VP.n16 B 0.021947f
C173 VP.n17 B 0.024022f
C174 VP.n18 B 0.021947f
C175 VP.n19 B 0.017726f
C176 VP.n20 B 0.021947f
C177 VP.t0 B 1.14666f
C178 VP.n21 B 0.508751f
C179 VP.t3 B 1.42091f
C180 VP.n22 B 0.482305f
C181 VP.n23 B 0.270161f
C182 VP.n24 B 0.037283f
C183 VP.n25 B 0.040698f
C184 VP.n26 B 0.043389f
C185 VP.n27 B 0.021947f
C186 VP.n28 B 0.021947f
C187 VP.n29 B 0.021947f
C188 VP.n30 B 0.043389f
C189 VP.n31 B 0.040698f
C190 VP.t1 B 1.14666f
C191 VP.n32 B 0.42623f
C192 VP.n33 B 0.037283f
C193 VP.n34 B 0.021947f
C194 VP.n35 B 0.021947f
C195 VP.n36 B 0.021947f
C196 VP.n37 B 0.040698f
C197 VP.n38 B 0.040698f
C198 VP.n39 B 0.036761f
C199 VP.n40 B 0.021947f
C200 VP.n41 B 0.021947f
C201 VP.n42 B 0.021947f
C202 VP.n43 B 0.040698f
C203 VP.n44 B 0.040698f
C204 VP.n45 B 0.030451f
C205 VP.n46 B 0.035416f
C206 VP.n47 B 1.26859f
C207 VP.t5 B 1.14666f
C208 VP.n48 B 0.512969f
C209 VP.n49 B 1.28428f
C210 VP.n50 B 0.035416f
C211 VP.n51 B 0.021947f
C212 VP.n52 B 0.040698f
C213 VP.n53 B 0.040698f
C214 VP.n54 B 0.027045f
C215 VP.n55 B 0.021947f
C216 VP.n56 B 0.021947f
C217 VP.n57 B 0.021947f
C218 VP.n58 B 0.040698f
C219 VP.n59 B 0.040698f
C220 VP.n60 B 0.024022f
C221 VP.n61 B 0.021947f
C222 VP.n62 B 0.021947f
C223 VP.n63 B 0.037283f
C224 VP.n64 B 0.040698f
C225 VP.n65 B 0.043389f
C226 VP.n66 B 0.021947f
C227 VP.n67 B 0.021947f
C228 VP.n68 B 0.021947f
C229 VP.n69 B 0.043389f
C230 VP.n70 B 0.040698f
C231 VP.t7 B 1.14666f
C232 VP.n71 B 0.42623f
C233 VP.n72 B 0.037283f
C234 VP.n73 B 0.021947f
C235 VP.n74 B 0.021947f
C236 VP.n75 B 0.021947f
C237 VP.n76 B 0.040698f
C238 VP.n77 B 0.040698f
C239 VP.n78 B 0.036761f
C240 VP.n79 B 0.021947f
C241 VP.n80 B 0.021947f
C242 VP.n81 B 0.021947f
C243 VP.n82 B 0.040698f
C244 VP.n83 B 0.040698f
C245 VP.n84 B 0.030451f
C246 VP.n85 B 0.035416f
C247 VP.n86 B 0.057261f
.ends

