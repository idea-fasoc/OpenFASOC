* NGSPICE file created from diff_pair_sample_0366.ext - technology: sky130A

.subckt diff_pair_sample_0366 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=0 ps=0 w=7.43 l=0.51
X1 B.t8 B.t6 B.t7 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=0 ps=0 w=7.43 l=0.51
X2 B.t5 B.t3 B.t4 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=0 ps=0 w=7.43 l=0.51
X3 VDD2.t1 VN.t0 VTAIL.t2 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=2.8977 ps=15.64 w=7.43 l=0.51
X4 B.t2 B.t0 B.t1 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=0 ps=0 w=7.43 l=0.51
X5 VDD1.t1 VP.t0 VTAIL.t1 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=2.8977 ps=15.64 w=7.43 l=0.51
X6 VDD1.t0 VP.t1 VTAIL.t0 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=2.8977 ps=15.64 w=7.43 l=0.51
X7 VDD2.t0 VN.t1 VTAIL.t3 w_n1306_n2458# sky130_fd_pr__pfet_01v8 ad=2.8977 pd=15.64 as=2.8977 ps=15.64 w=7.43 l=0.51
R0 B.n263 B.n46 585
R1 B.n265 B.n264 585
R2 B.n266 B.n45 585
R3 B.n268 B.n267 585
R4 B.n269 B.n44 585
R5 B.n271 B.n270 585
R6 B.n272 B.n43 585
R7 B.n274 B.n273 585
R8 B.n275 B.n42 585
R9 B.n277 B.n276 585
R10 B.n278 B.n41 585
R11 B.n280 B.n279 585
R12 B.n281 B.n40 585
R13 B.n283 B.n282 585
R14 B.n284 B.n39 585
R15 B.n286 B.n285 585
R16 B.n287 B.n38 585
R17 B.n289 B.n288 585
R18 B.n290 B.n37 585
R19 B.n292 B.n291 585
R20 B.n293 B.n36 585
R21 B.n295 B.n294 585
R22 B.n296 B.n35 585
R23 B.n298 B.n297 585
R24 B.n299 B.n34 585
R25 B.n301 B.n300 585
R26 B.n302 B.n33 585
R27 B.n304 B.n303 585
R28 B.n306 B.n30 585
R29 B.n308 B.n307 585
R30 B.n309 B.n29 585
R31 B.n311 B.n310 585
R32 B.n312 B.n28 585
R33 B.n314 B.n313 585
R34 B.n315 B.n27 585
R35 B.n317 B.n316 585
R36 B.n318 B.n23 585
R37 B.n320 B.n319 585
R38 B.n321 B.n22 585
R39 B.n323 B.n322 585
R40 B.n324 B.n21 585
R41 B.n326 B.n325 585
R42 B.n327 B.n20 585
R43 B.n329 B.n328 585
R44 B.n330 B.n19 585
R45 B.n332 B.n331 585
R46 B.n333 B.n18 585
R47 B.n335 B.n334 585
R48 B.n336 B.n17 585
R49 B.n338 B.n337 585
R50 B.n339 B.n16 585
R51 B.n341 B.n340 585
R52 B.n342 B.n15 585
R53 B.n344 B.n343 585
R54 B.n345 B.n14 585
R55 B.n347 B.n346 585
R56 B.n348 B.n13 585
R57 B.n350 B.n349 585
R58 B.n351 B.n12 585
R59 B.n353 B.n352 585
R60 B.n354 B.n11 585
R61 B.n356 B.n355 585
R62 B.n357 B.n10 585
R63 B.n359 B.n358 585
R64 B.n360 B.n9 585
R65 B.n362 B.n361 585
R66 B.n262 B.n261 585
R67 B.n260 B.n47 585
R68 B.n259 B.n258 585
R69 B.n257 B.n48 585
R70 B.n256 B.n255 585
R71 B.n254 B.n49 585
R72 B.n253 B.n252 585
R73 B.n251 B.n50 585
R74 B.n250 B.n249 585
R75 B.n248 B.n51 585
R76 B.n247 B.n246 585
R77 B.n245 B.n52 585
R78 B.n244 B.n243 585
R79 B.n242 B.n53 585
R80 B.n241 B.n240 585
R81 B.n239 B.n54 585
R82 B.n238 B.n237 585
R83 B.n236 B.n55 585
R84 B.n235 B.n234 585
R85 B.n233 B.n56 585
R86 B.n232 B.n231 585
R87 B.n230 B.n57 585
R88 B.n229 B.n228 585
R89 B.n227 B.n58 585
R90 B.n226 B.n225 585
R91 B.n224 B.n59 585
R92 B.n223 B.n222 585
R93 B.n122 B.n97 585
R94 B.n124 B.n123 585
R95 B.n125 B.n96 585
R96 B.n127 B.n126 585
R97 B.n128 B.n95 585
R98 B.n130 B.n129 585
R99 B.n131 B.n94 585
R100 B.n133 B.n132 585
R101 B.n134 B.n93 585
R102 B.n136 B.n135 585
R103 B.n137 B.n92 585
R104 B.n139 B.n138 585
R105 B.n140 B.n91 585
R106 B.n142 B.n141 585
R107 B.n143 B.n90 585
R108 B.n145 B.n144 585
R109 B.n146 B.n89 585
R110 B.n148 B.n147 585
R111 B.n149 B.n88 585
R112 B.n151 B.n150 585
R113 B.n152 B.n87 585
R114 B.n154 B.n153 585
R115 B.n155 B.n86 585
R116 B.n157 B.n156 585
R117 B.n158 B.n85 585
R118 B.n160 B.n159 585
R119 B.n161 B.n84 585
R120 B.n163 B.n162 585
R121 B.n165 B.n164 585
R122 B.n166 B.n80 585
R123 B.n168 B.n167 585
R124 B.n169 B.n79 585
R125 B.n171 B.n170 585
R126 B.n172 B.n78 585
R127 B.n174 B.n173 585
R128 B.n175 B.n77 585
R129 B.n177 B.n176 585
R130 B.n178 B.n74 585
R131 B.n181 B.n180 585
R132 B.n182 B.n73 585
R133 B.n184 B.n183 585
R134 B.n185 B.n72 585
R135 B.n187 B.n186 585
R136 B.n188 B.n71 585
R137 B.n190 B.n189 585
R138 B.n191 B.n70 585
R139 B.n193 B.n192 585
R140 B.n194 B.n69 585
R141 B.n196 B.n195 585
R142 B.n197 B.n68 585
R143 B.n199 B.n198 585
R144 B.n200 B.n67 585
R145 B.n202 B.n201 585
R146 B.n203 B.n66 585
R147 B.n205 B.n204 585
R148 B.n206 B.n65 585
R149 B.n208 B.n207 585
R150 B.n209 B.n64 585
R151 B.n211 B.n210 585
R152 B.n212 B.n63 585
R153 B.n214 B.n213 585
R154 B.n215 B.n62 585
R155 B.n217 B.n216 585
R156 B.n218 B.n61 585
R157 B.n220 B.n219 585
R158 B.n221 B.n60 585
R159 B.n121 B.n120 585
R160 B.n119 B.n98 585
R161 B.n118 B.n117 585
R162 B.n116 B.n99 585
R163 B.n115 B.n114 585
R164 B.n113 B.n100 585
R165 B.n112 B.n111 585
R166 B.n110 B.n101 585
R167 B.n109 B.n108 585
R168 B.n107 B.n102 585
R169 B.n106 B.n105 585
R170 B.n104 B.n103 585
R171 B.n2 B.n0 585
R172 B.n381 B.n1 585
R173 B.n380 B.n379 585
R174 B.n378 B.n3 585
R175 B.n377 B.n376 585
R176 B.n375 B.n4 585
R177 B.n374 B.n373 585
R178 B.n372 B.n5 585
R179 B.n371 B.n370 585
R180 B.n369 B.n6 585
R181 B.n368 B.n367 585
R182 B.n366 B.n7 585
R183 B.n365 B.n364 585
R184 B.n363 B.n8 585
R185 B.n383 B.n382 585
R186 B.n75 B.t9 557.275
R187 B.n81 B.t3 557.275
R188 B.n24 B.t6 557.275
R189 B.n31 B.t0 557.275
R190 B.n122 B.n121 511.721
R191 B.n363 B.n362 511.721
R192 B.n223 B.n60 511.721
R193 B.n261 B.n46 511.721
R194 B.n75 B.t11 309.943
R195 B.n31 B.t1 309.943
R196 B.n81 B.t5 309.943
R197 B.n24 B.t7 309.943
R198 B.n76 B.t10 293.652
R199 B.n32 B.t2 293.652
R200 B.n82 B.t4 293.652
R201 B.n25 B.t8 293.652
R202 B.n121 B.n98 163.367
R203 B.n117 B.n98 163.367
R204 B.n117 B.n116 163.367
R205 B.n116 B.n115 163.367
R206 B.n115 B.n100 163.367
R207 B.n111 B.n100 163.367
R208 B.n111 B.n110 163.367
R209 B.n110 B.n109 163.367
R210 B.n109 B.n102 163.367
R211 B.n105 B.n102 163.367
R212 B.n105 B.n104 163.367
R213 B.n104 B.n2 163.367
R214 B.n382 B.n2 163.367
R215 B.n382 B.n381 163.367
R216 B.n381 B.n380 163.367
R217 B.n380 B.n3 163.367
R218 B.n376 B.n3 163.367
R219 B.n376 B.n375 163.367
R220 B.n375 B.n374 163.367
R221 B.n374 B.n5 163.367
R222 B.n370 B.n5 163.367
R223 B.n370 B.n369 163.367
R224 B.n369 B.n368 163.367
R225 B.n368 B.n7 163.367
R226 B.n364 B.n7 163.367
R227 B.n364 B.n363 163.367
R228 B.n123 B.n122 163.367
R229 B.n123 B.n96 163.367
R230 B.n127 B.n96 163.367
R231 B.n128 B.n127 163.367
R232 B.n129 B.n128 163.367
R233 B.n129 B.n94 163.367
R234 B.n133 B.n94 163.367
R235 B.n134 B.n133 163.367
R236 B.n135 B.n134 163.367
R237 B.n135 B.n92 163.367
R238 B.n139 B.n92 163.367
R239 B.n140 B.n139 163.367
R240 B.n141 B.n140 163.367
R241 B.n141 B.n90 163.367
R242 B.n145 B.n90 163.367
R243 B.n146 B.n145 163.367
R244 B.n147 B.n146 163.367
R245 B.n147 B.n88 163.367
R246 B.n151 B.n88 163.367
R247 B.n152 B.n151 163.367
R248 B.n153 B.n152 163.367
R249 B.n153 B.n86 163.367
R250 B.n157 B.n86 163.367
R251 B.n158 B.n157 163.367
R252 B.n159 B.n158 163.367
R253 B.n159 B.n84 163.367
R254 B.n163 B.n84 163.367
R255 B.n164 B.n163 163.367
R256 B.n164 B.n80 163.367
R257 B.n168 B.n80 163.367
R258 B.n169 B.n168 163.367
R259 B.n170 B.n169 163.367
R260 B.n170 B.n78 163.367
R261 B.n174 B.n78 163.367
R262 B.n175 B.n174 163.367
R263 B.n176 B.n175 163.367
R264 B.n176 B.n74 163.367
R265 B.n181 B.n74 163.367
R266 B.n182 B.n181 163.367
R267 B.n183 B.n182 163.367
R268 B.n183 B.n72 163.367
R269 B.n187 B.n72 163.367
R270 B.n188 B.n187 163.367
R271 B.n189 B.n188 163.367
R272 B.n189 B.n70 163.367
R273 B.n193 B.n70 163.367
R274 B.n194 B.n193 163.367
R275 B.n195 B.n194 163.367
R276 B.n195 B.n68 163.367
R277 B.n199 B.n68 163.367
R278 B.n200 B.n199 163.367
R279 B.n201 B.n200 163.367
R280 B.n201 B.n66 163.367
R281 B.n205 B.n66 163.367
R282 B.n206 B.n205 163.367
R283 B.n207 B.n206 163.367
R284 B.n207 B.n64 163.367
R285 B.n211 B.n64 163.367
R286 B.n212 B.n211 163.367
R287 B.n213 B.n212 163.367
R288 B.n213 B.n62 163.367
R289 B.n217 B.n62 163.367
R290 B.n218 B.n217 163.367
R291 B.n219 B.n218 163.367
R292 B.n219 B.n60 163.367
R293 B.n224 B.n223 163.367
R294 B.n225 B.n224 163.367
R295 B.n225 B.n58 163.367
R296 B.n229 B.n58 163.367
R297 B.n230 B.n229 163.367
R298 B.n231 B.n230 163.367
R299 B.n231 B.n56 163.367
R300 B.n235 B.n56 163.367
R301 B.n236 B.n235 163.367
R302 B.n237 B.n236 163.367
R303 B.n237 B.n54 163.367
R304 B.n241 B.n54 163.367
R305 B.n242 B.n241 163.367
R306 B.n243 B.n242 163.367
R307 B.n243 B.n52 163.367
R308 B.n247 B.n52 163.367
R309 B.n248 B.n247 163.367
R310 B.n249 B.n248 163.367
R311 B.n249 B.n50 163.367
R312 B.n253 B.n50 163.367
R313 B.n254 B.n253 163.367
R314 B.n255 B.n254 163.367
R315 B.n255 B.n48 163.367
R316 B.n259 B.n48 163.367
R317 B.n260 B.n259 163.367
R318 B.n261 B.n260 163.367
R319 B.n362 B.n9 163.367
R320 B.n358 B.n9 163.367
R321 B.n358 B.n357 163.367
R322 B.n357 B.n356 163.367
R323 B.n356 B.n11 163.367
R324 B.n352 B.n11 163.367
R325 B.n352 B.n351 163.367
R326 B.n351 B.n350 163.367
R327 B.n350 B.n13 163.367
R328 B.n346 B.n13 163.367
R329 B.n346 B.n345 163.367
R330 B.n345 B.n344 163.367
R331 B.n344 B.n15 163.367
R332 B.n340 B.n15 163.367
R333 B.n340 B.n339 163.367
R334 B.n339 B.n338 163.367
R335 B.n338 B.n17 163.367
R336 B.n334 B.n17 163.367
R337 B.n334 B.n333 163.367
R338 B.n333 B.n332 163.367
R339 B.n332 B.n19 163.367
R340 B.n328 B.n19 163.367
R341 B.n328 B.n327 163.367
R342 B.n327 B.n326 163.367
R343 B.n326 B.n21 163.367
R344 B.n322 B.n21 163.367
R345 B.n322 B.n321 163.367
R346 B.n321 B.n320 163.367
R347 B.n320 B.n23 163.367
R348 B.n316 B.n23 163.367
R349 B.n316 B.n315 163.367
R350 B.n315 B.n314 163.367
R351 B.n314 B.n28 163.367
R352 B.n310 B.n28 163.367
R353 B.n310 B.n309 163.367
R354 B.n309 B.n308 163.367
R355 B.n308 B.n30 163.367
R356 B.n303 B.n30 163.367
R357 B.n303 B.n302 163.367
R358 B.n302 B.n301 163.367
R359 B.n301 B.n34 163.367
R360 B.n297 B.n34 163.367
R361 B.n297 B.n296 163.367
R362 B.n296 B.n295 163.367
R363 B.n295 B.n36 163.367
R364 B.n291 B.n36 163.367
R365 B.n291 B.n290 163.367
R366 B.n290 B.n289 163.367
R367 B.n289 B.n38 163.367
R368 B.n285 B.n38 163.367
R369 B.n285 B.n284 163.367
R370 B.n284 B.n283 163.367
R371 B.n283 B.n40 163.367
R372 B.n279 B.n40 163.367
R373 B.n279 B.n278 163.367
R374 B.n278 B.n277 163.367
R375 B.n277 B.n42 163.367
R376 B.n273 B.n42 163.367
R377 B.n273 B.n272 163.367
R378 B.n272 B.n271 163.367
R379 B.n271 B.n44 163.367
R380 B.n267 B.n44 163.367
R381 B.n267 B.n266 163.367
R382 B.n266 B.n265 163.367
R383 B.n265 B.n46 163.367
R384 B.n179 B.n76 59.5399
R385 B.n83 B.n82 59.5399
R386 B.n26 B.n25 59.5399
R387 B.n305 B.n32 59.5399
R388 B.n361 B.n8 33.2493
R389 B.n263 B.n262 33.2493
R390 B.n222 B.n221 33.2493
R391 B.n120 B.n97 33.2493
R392 B B.n383 18.0485
R393 B.n76 B.n75 16.2914
R394 B.n82 B.n81 16.2914
R395 B.n25 B.n24 16.2914
R396 B.n32 B.n31 16.2914
R397 B.n361 B.n360 10.6151
R398 B.n360 B.n359 10.6151
R399 B.n359 B.n10 10.6151
R400 B.n355 B.n10 10.6151
R401 B.n355 B.n354 10.6151
R402 B.n354 B.n353 10.6151
R403 B.n353 B.n12 10.6151
R404 B.n349 B.n12 10.6151
R405 B.n349 B.n348 10.6151
R406 B.n348 B.n347 10.6151
R407 B.n347 B.n14 10.6151
R408 B.n343 B.n14 10.6151
R409 B.n343 B.n342 10.6151
R410 B.n342 B.n341 10.6151
R411 B.n341 B.n16 10.6151
R412 B.n337 B.n16 10.6151
R413 B.n337 B.n336 10.6151
R414 B.n336 B.n335 10.6151
R415 B.n335 B.n18 10.6151
R416 B.n331 B.n18 10.6151
R417 B.n331 B.n330 10.6151
R418 B.n330 B.n329 10.6151
R419 B.n329 B.n20 10.6151
R420 B.n325 B.n20 10.6151
R421 B.n325 B.n324 10.6151
R422 B.n324 B.n323 10.6151
R423 B.n323 B.n22 10.6151
R424 B.n319 B.n318 10.6151
R425 B.n318 B.n317 10.6151
R426 B.n317 B.n27 10.6151
R427 B.n313 B.n27 10.6151
R428 B.n313 B.n312 10.6151
R429 B.n312 B.n311 10.6151
R430 B.n311 B.n29 10.6151
R431 B.n307 B.n29 10.6151
R432 B.n307 B.n306 10.6151
R433 B.n304 B.n33 10.6151
R434 B.n300 B.n33 10.6151
R435 B.n300 B.n299 10.6151
R436 B.n299 B.n298 10.6151
R437 B.n298 B.n35 10.6151
R438 B.n294 B.n35 10.6151
R439 B.n294 B.n293 10.6151
R440 B.n293 B.n292 10.6151
R441 B.n292 B.n37 10.6151
R442 B.n288 B.n37 10.6151
R443 B.n288 B.n287 10.6151
R444 B.n287 B.n286 10.6151
R445 B.n286 B.n39 10.6151
R446 B.n282 B.n39 10.6151
R447 B.n282 B.n281 10.6151
R448 B.n281 B.n280 10.6151
R449 B.n280 B.n41 10.6151
R450 B.n276 B.n41 10.6151
R451 B.n276 B.n275 10.6151
R452 B.n275 B.n274 10.6151
R453 B.n274 B.n43 10.6151
R454 B.n270 B.n43 10.6151
R455 B.n270 B.n269 10.6151
R456 B.n269 B.n268 10.6151
R457 B.n268 B.n45 10.6151
R458 B.n264 B.n45 10.6151
R459 B.n264 B.n263 10.6151
R460 B.n222 B.n59 10.6151
R461 B.n226 B.n59 10.6151
R462 B.n227 B.n226 10.6151
R463 B.n228 B.n227 10.6151
R464 B.n228 B.n57 10.6151
R465 B.n232 B.n57 10.6151
R466 B.n233 B.n232 10.6151
R467 B.n234 B.n233 10.6151
R468 B.n234 B.n55 10.6151
R469 B.n238 B.n55 10.6151
R470 B.n239 B.n238 10.6151
R471 B.n240 B.n239 10.6151
R472 B.n240 B.n53 10.6151
R473 B.n244 B.n53 10.6151
R474 B.n245 B.n244 10.6151
R475 B.n246 B.n245 10.6151
R476 B.n246 B.n51 10.6151
R477 B.n250 B.n51 10.6151
R478 B.n251 B.n250 10.6151
R479 B.n252 B.n251 10.6151
R480 B.n252 B.n49 10.6151
R481 B.n256 B.n49 10.6151
R482 B.n257 B.n256 10.6151
R483 B.n258 B.n257 10.6151
R484 B.n258 B.n47 10.6151
R485 B.n262 B.n47 10.6151
R486 B.n124 B.n97 10.6151
R487 B.n125 B.n124 10.6151
R488 B.n126 B.n125 10.6151
R489 B.n126 B.n95 10.6151
R490 B.n130 B.n95 10.6151
R491 B.n131 B.n130 10.6151
R492 B.n132 B.n131 10.6151
R493 B.n132 B.n93 10.6151
R494 B.n136 B.n93 10.6151
R495 B.n137 B.n136 10.6151
R496 B.n138 B.n137 10.6151
R497 B.n138 B.n91 10.6151
R498 B.n142 B.n91 10.6151
R499 B.n143 B.n142 10.6151
R500 B.n144 B.n143 10.6151
R501 B.n144 B.n89 10.6151
R502 B.n148 B.n89 10.6151
R503 B.n149 B.n148 10.6151
R504 B.n150 B.n149 10.6151
R505 B.n150 B.n87 10.6151
R506 B.n154 B.n87 10.6151
R507 B.n155 B.n154 10.6151
R508 B.n156 B.n155 10.6151
R509 B.n156 B.n85 10.6151
R510 B.n160 B.n85 10.6151
R511 B.n161 B.n160 10.6151
R512 B.n162 B.n161 10.6151
R513 B.n166 B.n165 10.6151
R514 B.n167 B.n166 10.6151
R515 B.n167 B.n79 10.6151
R516 B.n171 B.n79 10.6151
R517 B.n172 B.n171 10.6151
R518 B.n173 B.n172 10.6151
R519 B.n173 B.n77 10.6151
R520 B.n177 B.n77 10.6151
R521 B.n178 B.n177 10.6151
R522 B.n180 B.n73 10.6151
R523 B.n184 B.n73 10.6151
R524 B.n185 B.n184 10.6151
R525 B.n186 B.n185 10.6151
R526 B.n186 B.n71 10.6151
R527 B.n190 B.n71 10.6151
R528 B.n191 B.n190 10.6151
R529 B.n192 B.n191 10.6151
R530 B.n192 B.n69 10.6151
R531 B.n196 B.n69 10.6151
R532 B.n197 B.n196 10.6151
R533 B.n198 B.n197 10.6151
R534 B.n198 B.n67 10.6151
R535 B.n202 B.n67 10.6151
R536 B.n203 B.n202 10.6151
R537 B.n204 B.n203 10.6151
R538 B.n204 B.n65 10.6151
R539 B.n208 B.n65 10.6151
R540 B.n209 B.n208 10.6151
R541 B.n210 B.n209 10.6151
R542 B.n210 B.n63 10.6151
R543 B.n214 B.n63 10.6151
R544 B.n215 B.n214 10.6151
R545 B.n216 B.n215 10.6151
R546 B.n216 B.n61 10.6151
R547 B.n220 B.n61 10.6151
R548 B.n221 B.n220 10.6151
R549 B.n120 B.n119 10.6151
R550 B.n119 B.n118 10.6151
R551 B.n118 B.n99 10.6151
R552 B.n114 B.n99 10.6151
R553 B.n114 B.n113 10.6151
R554 B.n113 B.n112 10.6151
R555 B.n112 B.n101 10.6151
R556 B.n108 B.n101 10.6151
R557 B.n108 B.n107 10.6151
R558 B.n107 B.n106 10.6151
R559 B.n106 B.n103 10.6151
R560 B.n103 B.n0 10.6151
R561 B.n379 B.n1 10.6151
R562 B.n379 B.n378 10.6151
R563 B.n378 B.n377 10.6151
R564 B.n377 B.n4 10.6151
R565 B.n373 B.n4 10.6151
R566 B.n373 B.n372 10.6151
R567 B.n372 B.n371 10.6151
R568 B.n371 B.n6 10.6151
R569 B.n367 B.n6 10.6151
R570 B.n367 B.n366 10.6151
R571 B.n366 B.n365 10.6151
R572 B.n365 B.n8 10.6151
R573 B.n26 B.n22 8.74196
R574 B.n305 B.n304 8.74196
R575 B.n162 B.n83 8.74196
R576 B.n180 B.n179 8.74196
R577 B.n383 B.n0 2.81026
R578 B.n383 B.n1 2.81026
R579 B.n319 B.n26 1.87367
R580 B.n306 B.n305 1.87367
R581 B.n165 B.n83 1.87367
R582 B.n179 B.n178 1.87367
R583 VN VN.t1 625.949
R584 VN VN.t0 589.953
R585 VTAIL.n154 VTAIL.n120 756.745
R586 VTAIL.n34 VTAIL.n0 756.745
R587 VTAIL.n114 VTAIL.n80 756.745
R588 VTAIL.n74 VTAIL.n40 756.745
R589 VTAIL.n132 VTAIL.n131 585
R590 VTAIL.n137 VTAIL.n136 585
R591 VTAIL.n139 VTAIL.n138 585
R592 VTAIL.n128 VTAIL.n127 585
R593 VTAIL.n145 VTAIL.n144 585
R594 VTAIL.n147 VTAIL.n146 585
R595 VTAIL.n124 VTAIL.n123 585
R596 VTAIL.n153 VTAIL.n152 585
R597 VTAIL.n155 VTAIL.n154 585
R598 VTAIL.n12 VTAIL.n11 585
R599 VTAIL.n17 VTAIL.n16 585
R600 VTAIL.n19 VTAIL.n18 585
R601 VTAIL.n8 VTAIL.n7 585
R602 VTAIL.n25 VTAIL.n24 585
R603 VTAIL.n27 VTAIL.n26 585
R604 VTAIL.n4 VTAIL.n3 585
R605 VTAIL.n33 VTAIL.n32 585
R606 VTAIL.n35 VTAIL.n34 585
R607 VTAIL.n115 VTAIL.n114 585
R608 VTAIL.n113 VTAIL.n112 585
R609 VTAIL.n84 VTAIL.n83 585
R610 VTAIL.n107 VTAIL.n106 585
R611 VTAIL.n105 VTAIL.n104 585
R612 VTAIL.n88 VTAIL.n87 585
R613 VTAIL.n99 VTAIL.n98 585
R614 VTAIL.n97 VTAIL.n96 585
R615 VTAIL.n92 VTAIL.n91 585
R616 VTAIL.n75 VTAIL.n74 585
R617 VTAIL.n73 VTAIL.n72 585
R618 VTAIL.n44 VTAIL.n43 585
R619 VTAIL.n67 VTAIL.n66 585
R620 VTAIL.n65 VTAIL.n64 585
R621 VTAIL.n48 VTAIL.n47 585
R622 VTAIL.n59 VTAIL.n58 585
R623 VTAIL.n57 VTAIL.n56 585
R624 VTAIL.n52 VTAIL.n51 585
R625 VTAIL.n133 VTAIL.t2 327.483
R626 VTAIL.n13 VTAIL.t1 327.483
R627 VTAIL.n93 VTAIL.t0 327.483
R628 VTAIL.n53 VTAIL.t3 327.483
R629 VTAIL.n137 VTAIL.n131 171.744
R630 VTAIL.n138 VTAIL.n137 171.744
R631 VTAIL.n138 VTAIL.n127 171.744
R632 VTAIL.n145 VTAIL.n127 171.744
R633 VTAIL.n146 VTAIL.n145 171.744
R634 VTAIL.n146 VTAIL.n123 171.744
R635 VTAIL.n153 VTAIL.n123 171.744
R636 VTAIL.n154 VTAIL.n153 171.744
R637 VTAIL.n17 VTAIL.n11 171.744
R638 VTAIL.n18 VTAIL.n17 171.744
R639 VTAIL.n18 VTAIL.n7 171.744
R640 VTAIL.n25 VTAIL.n7 171.744
R641 VTAIL.n26 VTAIL.n25 171.744
R642 VTAIL.n26 VTAIL.n3 171.744
R643 VTAIL.n33 VTAIL.n3 171.744
R644 VTAIL.n34 VTAIL.n33 171.744
R645 VTAIL.n114 VTAIL.n113 171.744
R646 VTAIL.n113 VTAIL.n83 171.744
R647 VTAIL.n106 VTAIL.n83 171.744
R648 VTAIL.n106 VTAIL.n105 171.744
R649 VTAIL.n105 VTAIL.n87 171.744
R650 VTAIL.n98 VTAIL.n87 171.744
R651 VTAIL.n98 VTAIL.n97 171.744
R652 VTAIL.n97 VTAIL.n91 171.744
R653 VTAIL.n74 VTAIL.n73 171.744
R654 VTAIL.n73 VTAIL.n43 171.744
R655 VTAIL.n66 VTAIL.n43 171.744
R656 VTAIL.n66 VTAIL.n65 171.744
R657 VTAIL.n65 VTAIL.n47 171.744
R658 VTAIL.n58 VTAIL.n47 171.744
R659 VTAIL.n58 VTAIL.n57 171.744
R660 VTAIL.n57 VTAIL.n51 171.744
R661 VTAIL.t2 VTAIL.n131 85.8723
R662 VTAIL.t1 VTAIL.n11 85.8723
R663 VTAIL.t0 VTAIL.n91 85.8723
R664 VTAIL.t3 VTAIL.n51 85.8723
R665 VTAIL.n159 VTAIL.n158 31.9914
R666 VTAIL.n39 VTAIL.n38 31.9914
R667 VTAIL.n119 VTAIL.n118 31.9914
R668 VTAIL.n79 VTAIL.n78 31.9914
R669 VTAIL.n79 VTAIL.n39 20.2376
R670 VTAIL.n159 VTAIL.n119 19.5134
R671 VTAIL.n133 VTAIL.n132 16.3891
R672 VTAIL.n13 VTAIL.n12 16.3891
R673 VTAIL.n93 VTAIL.n92 16.3891
R674 VTAIL.n53 VTAIL.n52 16.3891
R675 VTAIL.n136 VTAIL.n135 12.8005
R676 VTAIL.n16 VTAIL.n15 12.8005
R677 VTAIL.n96 VTAIL.n95 12.8005
R678 VTAIL.n56 VTAIL.n55 12.8005
R679 VTAIL.n139 VTAIL.n130 12.0247
R680 VTAIL.n19 VTAIL.n10 12.0247
R681 VTAIL.n99 VTAIL.n90 12.0247
R682 VTAIL.n59 VTAIL.n50 12.0247
R683 VTAIL.n140 VTAIL.n128 11.249
R684 VTAIL.n20 VTAIL.n8 11.249
R685 VTAIL.n100 VTAIL.n88 11.249
R686 VTAIL.n60 VTAIL.n48 11.249
R687 VTAIL.n144 VTAIL.n143 10.4732
R688 VTAIL.n24 VTAIL.n23 10.4732
R689 VTAIL.n104 VTAIL.n103 10.4732
R690 VTAIL.n64 VTAIL.n63 10.4732
R691 VTAIL.n147 VTAIL.n126 9.69747
R692 VTAIL.n27 VTAIL.n6 9.69747
R693 VTAIL.n107 VTAIL.n86 9.69747
R694 VTAIL.n67 VTAIL.n46 9.69747
R695 VTAIL.n158 VTAIL.n157 9.45567
R696 VTAIL.n38 VTAIL.n37 9.45567
R697 VTAIL.n118 VTAIL.n117 9.45567
R698 VTAIL.n78 VTAIL.n77 9.45567
R699 VTAIL.n157 VTAIL.n156 9.3005
R700 VTAIL.n151 VTAIL.n150 9.3005
R701 VTAIL.n149 VTAIL.n148 9.3005
R702 VTAIL.n126 VTAIL.n125 9.3005
R703 VTAIL.n143 VTAIL.n142 9.3005
R704 VTAIL.n141 VTAIL.n140 9.3005
R705 VTAIL.n130 VTAIL.n129 9.3005
R706 VTAIL.n135 VTAIL.n134 9.3005
R707 VTAIL.n122 VTAIL.n121 9.3005
R708 VTAIL.n37 VTAIL.n36 9.3005
R709 VTAIL.n31 VTAIL.n30 9.3005
R710 VTAIL.n29 VTAIL.n28 9.3005
R711 VTAIL.n6 VTAIL.n5 9.3005
R712 VTAIL.n23 VTAIL.n22 9.3005
R713 VTAIL.n21 VTAIL.n20 9.3005
R714 VTAIL.n10 VTAIL.n9 9.3005
R715 VTAIL.n15 VTAIL.n14 9.3005
R716 VTAIL.n2 VTAIL.n1 9.3005
R717 VTAIL.n117 VTAIL.n116 9.3005
R718 VTAIL.n82 VTAIL.n81 9.3005
R719 VTAIL.n111 VTAIL.n110 9.3005
R720 VTAIL.n109 VTAIL.n108 9.3005
R721 VTAIL.n86 VTAIL.n85 9.3005
R722 VTAIL.n103 VTAIL.n102 9.3005
R723 VTAIL.n101 VTAIL.n100 9.3005
R724 VTAIL.n90 VTAIL.n89 9.3005
R725 VTAIL.n95 VTAIL.n94 9.3005
R726 VTAIL.n77 VTAIL.n76 9.3005
R727 VTAIL.n42 VTAIL.n41 9.3005
R728 VTAIL.n71 VTAIL.n70 9.3005
R729 VTAIL.n69 VTAIL.n68 9.3005
R730 VTAIL.n46 VTAIL.n45 9.3005
R731 VTAIL.n63 VTAIL.n62 9.3005
R732 VTAIL.n61 VTAIL.n60 9.3005
R733 VTAIL.n50 VTAIL.n49 9.3005
R734 VTAIL.n55 VTAIL.n54 9.3005
R735 VTAIL.n148 VTAIL.n124 8.92171
R736 VTAIL.n28 VTAIL.n4 8.92171
R737 VTAIL.n108 VTAIL.n84 8.92171
R738 VTAIL.n68 VTAIL.n44 8.92171
R739 VTAIL.n152 VTAIL.n151 8.14595
R740 VTAIL.n32 VTAIL.n31 8.14595
R741 VTAIL.n112 VTAIL.n111 8.14595
R742 VTAIL.n72 VTAIL.n71 8.14595
R743 VTAIL.n155 VTAIL.n122 7.3702
R744 VTAIL.n158 VTAIL.n120 7.3702
R745 VTAIL.n35 VTAIL.n2 7.3702
R746 VTAIL.n38 VTAIL.n0 7.3702
R747 VTAIL.n118 VTAIL.n80 7.3702
R748 VTAIL.n115 VTAIL.n82 7.3702
R749 VTAIL.n78 VTAIL.n40 7.3702
R750 VTAIL.n75 VTAIL.n42 7.3702
R751 VTAIL.n156 VTAIL.n155 6.59444
R752 VTAIL.n156 VTAIL.n120 6.59444
R753 VTAIL.n36 VTAIL.n35 6.59444
R754 VTAIL.n36 VTAIL.n0 6.59444
R755 VTAIL.n116 VTAIL.n80 6.59444
R756 VTAIL.n116 VTAIL.n115 6.59444
R757 VTAIL.n76 VTAIL.n40 6.59444
R758 VTAIL.n76 VTAIL.n75 6.59444
R759 VTAIL.n152 VTAIL.n122 5.81868
R760 VTAIL.n32 VTAIL.n2 5.81868
R761 VTAIL.n112 VTAIL.n82 5.81868
R762 VTAIL.n72 VTAIL.n42 5.81868
R763 VTAIL.n151 VTAIL.n124 5.04292
R764 VTAIL.n31 VTAIL.n4 5.04292
R765 VTAIL.n111 VTAIL.n84 5.04292
R766 VTAIL.n71 VTAIL.n44 5.04292
R767 VTAIL.n148 VTAIL.n147 4.26717
R768 VTAIL.n28 VTAIL.n27 4.26717
R769 VTAIL.n108 VTAIL.n107 4.26717
R770 VTAIL.n68 VTAIL.n67 4.26717
R771 VTAIL.n134 VTAIL.n133 3.71019
R772 VTAIL.n14 VTAIL.n13 3.71019
R773 VTAIL.n94 VTAIL.n93 3.71019
R774 VTAIL.n54 VTAIL.n53 3.71019
R775 VTAIL.n144 VTAIL.n126 3.49141
R776 VTAIL.n24 VTAIL.n6 3.49141
R777 VTAIL.n104 VTAIL.n86 3.49141
R778 VTAIL.n64 VTAIL.n46 3.49141
R779 VTAIL.n143 VTAIL.n128 2.71565
R780 VTAIL.n23 VTAIL.n8 2.71565
R781 VTAIL.n103 VTAIL.n88 2.71565
R782 VTAIL.n63 VTAIL.n48 2.71565
R783 VTAIL.n140 VTAIL.n139 1.93989
R784 VTAIL.n20 VTAIL.n19 1.93989
R785 VTAIL.n100 VTAIL.n99 1.93989
R786 VTAIL.n60 VTAIL.n59 1.93989
R787 VTAIL.n136 VTAIL.n130 1.16414
R788 VTAIL.n16 VTAIL.n10 1.16414
R789 VTAIL.n96 VTAIL.n90 1.16414
R790 VTAIL.n56 VTAIL.n50 1.16414
R791 VTAIL.n119 VTAIL.n79 0.832397
R792 VTAIL VTAIL.n39 0.709552
R793 VTAIL.n135 VTAIL.n132 0.388379
R794 VTAIL.n15 VTAIL.n12 0.388379
R795 VTAIL.n95 VTAIL.n92 0.388379
R796 VTAIL.n55 VTAIL.n52 0.388379
R797 VTAIL.n134 VTAIL.n129 0.155672
R798 VTAIL.n141 VTAIL.n129 0.155672
R799 VTAIL.n142 VTAIL.n141 0.155672
R800 VTAIL.n142 VTAIL.n125 0.155672
R801 VTAIL.n149 VTAIL.n125 0.155672
R802 VTAIL.n150 VTAIL.n149 0.155672
R803 VTAIL.n150 VTAIL.n121 0.155672
R804 VTAIL.n157 VTAIL.n121 0.155672
R805 VTAIL.n14 VTAIL.n9 0.155672
R806 VTAIL.n21 VTAIL.n9 0.155672
R807 VTAIL.n22 VTAIL.n21 0.155672
R808 VTAIL.n22 VTAIL.n5 0.155672
R809 VTAIL.n29 VTAIL.n5 0.155672
R810 VTAIL.n30 VTAIL.n29 0.155672
R811 VTAIL.n30 VTAIL.n1 0.155672
R812 VTAIL.n37 VTAIL.n1 0.155672
R813 VTAIL.n117 VTAIL.n81 0.155672
R814 VTAIL.n110 VTAIL.n81 0.155672
R815 VTAIL.n110 VTAIL.n109 0.155672
R816 VTAIL.n109 VTAIL.n85 0.155672
R817 VTAIL.n102 VTAIL.n85 0.155672
R818 VTAIL.n102 VTAIL.n101 0.155672
R819 VTAIL.n101 VTAIL.n89 0.155672
R820 VTAIL.n94 VTAIL.n89 0.155672
R821 VTAIL.n77 VTAIL.n41 0.155672
R822 VTAIL.n70 VTAIL.n41 0.155672
R823 VTAIL.n70 VTAIL.n69 0.155672
R824 VTAIL.n69 VTAIL.n45 0.155672
R825 VTAIL.n62 VTAIL.n45 0.155672
R826 VTAIL.n62 VTAIL.n61 0.155672
R827 VTAIL.n61 VTAIL.n49 0.155672
R828 VTAIL.n54 VTAIL.n49 0.155672
R829 VTAIL VTAIL.n159 0.123345
R830 VDD2.n73 VDD2.n39 756.745
R831 VDD2.n34 VDD2.n0 756.745
R832 VDD2.n74 VDD2.n73 585
R833 VDD2.n72 VDD2.n71 585
R834 VDD2.n43 VDD2.n42 585
R835 VDD2.n66 VDD2.n65 585
R836 VDD2.n64 VDD2.n63 585
R837 VDD2.n47 VDD2.n46 585
R838 VDD2.n58 VDD2.n57 585
R839 VDD2.n56 VDD2.n55 585
R840 VDD2.n51 VDD2.n50 585
R841 VDD2.n12 VDD2.n11 585
R842 VDD2.n17 VDD2.n16 585
R843 VDD2.n19 VDD2.n18 585
R844 VDD2.n8 VDD2.n7 585
R845 VDD2.n25 VDD2.n24 585
R846 VDD2.n27 VDD2.n26 585
R847 VDD2.n4 VDD2.n3 585
R848 VDD2.n33 VDD2.n32 585
R849 VDD2.n35 VDD2.n34 585
R850 VDD2.n52 VDD2.t0 327.483
R851 VDD2.n13 VDD2.t1 327.483
R852 VDD2.n73 VDD2.n72 171.744
R853 VDD2.n72 VDD2.n42 171.744
R854 VDD2.n65 VDD2.n42 171.744
R855 VDD2.n65 VDD2.n64 171.744
R856 VDD2.n64 VDD2.n46 171.744
R857 VDD2.n57 VDD2.n46 171.744
R858 VDD2.n57 VDD2.n56 171.744
R859 VDD2.n56 VDD2.n50 171.744
R860 VDD2.n17 VDD2.n11 171.744
R861 VDD2.n18 VDD2.n17 171.744
R862 VDD2.n18 VDD2.n7 171.744
R863 VDD2.n25 VDD2.n7 171.744
R864 VDD2.n26 VDD2.n25 171.744
R865 VDD2.n26 VDD2.n3 171.744
R866 VDD2.n33 VDD2.n3 171.744
R867 VDD2.n34 VDD2.n33 171.744
R868 VDD2.t0 VDD2.n50 85.8723
R869 VDD2.t1 VDD2.n11 85.8723
R870 VDD2.n78 VDD2.n38 80.2003
R871 VDD2.n78 VDD2.n77 48.6702
R872 VDD2.n52 VDD2.n51 16.3891
R873 VDD2.n13 VDD2.n12 16.3891
R874 VDD2.n55 VDD2.n54 12.8005
R875 VDD2.n16 VDD2.n15 12.8005
R876 VDD2.n58 VDD2.n49 12.0247
R877 VDD2.n19 VDD2.n10 12.0247
R878 VDD2.n59 VDD2.n47 11.249
R879 VDD2.n20 VDD2.n8 11.249
R880 VDD2.n63 VDD2.n62 10.4732
R881 VDD2.n24 VDD2.n23 10.4732
R882 VDD2.n66 VDD2.n45 9.69747
R883 VDD2.n27 VDD2.n6 9.69747
R884 VDD2.n77 VDD2.n76 9.45567
R885 VDD2.n38 VDD2.n37 9.45567
R886 VDD2.n76 VDD2.n75 9.3005
R887 VDD2.n41 VDD2.n40 9.3005
R888 VDD2.n70 VDD2.n69 9.3005
R889 VDD2.n68 VDD2.n67 9.3005
R890 VDD2.n45 VDD2.n44 9.3005
R891 VDD2.n62 VDD2.n61 9.3005
R892 VDD2.n60 VDD2.n59 9.3005
R893 VDD2.n49 VDD2.n48 9.3005
R894 VDD2.n54 VDD2.n53 9.3005
R895 VDD2.n37 VDD2.n36 9.3005
R896 VDD2.n31 VDD2.n30 9.3005
R897 VDD2.n29 VDD2.n28 9.3005
R898 VDD2.n6 VDD2.n5 9.3005
R899 VDD2.n23 VDD2.n22 9.3005
R900 VDD2.n21 VDD2.n20 9.3005
R901 VDD2.n10 VDD2.n9 9.3005
R902 VDD2.n15 VDD2.n14 9.3005
R903 VDD2.n2 VDD2.n1 9.3005
R904 VDD2.n67 VDD2.n43 8.92171
R905 VDD2.n28 VDD2.n4 8.92171
R906 VDD2.n71 VDD2.n70 8.14595
R907 VDD2.n32 VDD2.n31 8.14595
R908 VDD2.n77 VDD2.n39 7.3702
R909 VDD2.n74 VDD2.n41 7.3702
R910 VDD2.n35 VDD2.n2 7.3702
R911 VDD2.n38 VDD2.n0 7.3702
R912 VDD2.n75 VDD2.n39 6.59444
R913 VDD2.n75 VDD2.n74 6.59444
R914 VDD2.n36 VDD2.n35 6.59444
R915 VDD2.n36 VDD2.n0 6.59444
R916 VDD2.n71 VDD2.n41 5.81868
R917 VDD2.n32 VDD2.n2 5.81868
R918 VDD2.n70 VDD2.n43 5.04292
R919 VDD2.n31 VDD2.n4 5.04292
R920 VDD2.n67 VDD2.n66 4.26717
R921 VDD2.n28 VDD2.n27 4.26717
R922 VDD2.n53 VDD2.n52 3.71019
R923 VDD2.n14 VDD2.n13 3.71019
R924 VDD2.n63 VDD2.n45 3.49141
R925 VDD2.n24 VDD2.n6 3.49141
R926 VDD2.n62 VDD2.n47 2.71565
R927 VDD2.n23 VDD2.n8 2.71565
R928 VDD2.n59 VDD2.n58 1.93989
R929 VDD2.n20 VDD2.n19 1.93989
R930 VDD2.n55 VDD2.n49 1.16414
R931 VDD2.n16 VDD2.n10 1.16414
R932 VDD2.n54 VDD2.n51 0.388379
R933 VDD2.n15 VDD2.n12 0.388379
R934 VDD2 VDD2.n78 0.239724
R935 VDD2.n76 VDD2.n40 0.155672
R936 VDD2.n69 VDD2.n40 0.155672
R937 VDD2.n69 VDD2.n68 0.155672
R938 VDD2.n68 VDD2.n44 0.155672
R939 VDD2.n61 VDD2.n44 0.155672
R940 VDD2.n61 VDD2.n60 0.155672
R941 VDD2.n60 VDD2.n48 0.155672
R942 VDD2.n53 VDD2.n48 0.155672
R943 VDD2.n14 VDD2.n9 0.155672
R944 VDD2.n21 VDD2.n9 0.155672
R945 VDD2.n22 VDD2.n21 0.155672
R946 VDD2.n22 VDD2.n5 0.155672
R947 VDD2.n29 VDD2.n5 0.155672
R948 VDD2.n30 VDD2.n29 0.155672
R949 VDD2.n30 VDD2.n1 0.155672
R950 VDD2.n37 VDD2.n1 0.155672
R951 VP.n0 VP.t1 625.569
R952 VP.n0 VP.t0 589.903
R953 VP VP.n0 0.0516364
R954 VDD1.n34 VDD1.n0 756.745
R955 VDD1.n73 VDD1.n39 756.745
R956 VDD1.n35 VDD1.n34 585
R957 VDD1.n33 VDD1.n32 585
R958 VDD1.n4 VDD1.n3 585
R959 VDD1.n27 VDD1.n26 585
R960 VDD1.n25 VDD1.n24 585
R961 VDD1.n8 VDD1.n7 585
R962 VDD1.n19 VDD1.n18 585
R963 VDD1.n17 VDD1.n16 585
R964 VDD1.n12 VDD1.n11 585
R965 VDD1.n51 VDD1.n50 585
R966 VDD1.n56 VDD1.n55 585
R967 VDD1.n58 VDD1.n57 585
R968 VDD1.n47 VDD1.n46 585
R969 VDD1.n64 VDD1.n63 585
R970 VDD1.n66 VDD1.n65 585
R971 VDD1.n43 VDD1.n42 585
R972 VDD1.n72 VDD1.n71 585
R973 VDD1.n74 VDD1.n73 585
R974 VDD1.n13 VDD1.t0 327.483
R975 VDD1.n52 VDD1.t1 327.483
R976 VDD1.n34 VDD1.n33 171.744
R977 VDD1.n33 VDD1.n3 171.744
R978 VDD1.n26 VDD1.n3 171.744
R979 VDD1.n26 VDD1.n25 171.744
R980 VDD1.n25 VDD1.n7 171.744
R981 VDD1.n18 VDD1.n7 171.744
R982 VDD1.n18 VDD1.n17 171.744
R983 VDD1.n17 VDD1.n11 171.744
R984 VDD1.n56 VDD1.n50 171.744
R985 VDD1.n57 VDD1.n56 171.744
R986 VDD1.n57 VDD1.n46 171.744
R987 VDD1.n64 VDD1.n46 171.744
R988 VDD1.n65 VDD1.n64 171.744
R989 VDD1.n65 VDD1.n42 171.744
R990 VDD1.n72 VDD1.n42 171.744
R991 VDD1.n73 VDD1.n72 171.744
R992 VDD1.t0 VDD1.n11 85.8723
R993 VDD1.t1 VDD1.n50 85.8723
R994 VDD1 VDD1.n77 80.9062
R995 VDD1 VDD1.n38 48.9094
R996 VDD1.n13 VDD1.n12 16.3891
R997 VDD1.n52 VDD1.n51 16.3891
R998 VDD1.n16 VDD1.n15 12.8005
R999 VDD1.n55 VDD1.n54 12.8005
R1000 VDD1.n19 VDD1.n10 12.0247
R1001 VDD1.n58 VDD1.n49 12.0247
R1002 VDD1.n20 VDD1.n8 11.249
R1003 VDD1.n59 VDD1.n47 11.249
R1004 VDD1.n24 VDD1.n23 10.4732
R1005 VDD1.n63 VDD1.n62 10.4732
R1006 VDD1.n27 VDD1.n6 9.69747
R1007 VDD1.n66 VDD1.n45 9.69747
R1008 VDD1.n38 VDD1.n37 9.45567
R1009 VDD1.n77 VDD1.n76 9.45567
R1010 VDD1.n37 VDD1.n36 9.3005
R1011 VDD1.n2 VDD1.n1 9.3005
R1012 VDD1.n31 VDD1.n30 9.3005
R1013 VDD1.n29 VDD1.n28 9.3005
R1014 VDD1.n6 VDD1.n5 9.3005
R1015 VDD1.n23 VDD1.n22 9.3005
R1016 VDD1.n21 VDD1.n20 9.3005
R1017 VDD1.n10 VDD1.n9 9.3005
R1018 VDD1.n15 VDD1.n14 9.3005
R1019 VDD1.n76 VDD1.n75 9.3005
R1020 VDD1.n70 VDD1.n69 9.3005
R1021 VDD1.n68 VDD1.n67 9.3005
R1022 VDD1.n45 VDD1.n44 9.3005
R1023 VDD1.n62 VDD1.n61 9.3005
R1024 VDD1.n60 VDD1.n59 9.3005
R1025 VDD1.n49 VDD1.n48 9.3005
R1026 VDD1.n54 VDD1.n53 9.3005
R1027 VDD1.n41 VDD1.n40 9.3005
R1028 VDD1.n28 VDD1.n4 8.92171
R1029 VDD1.n67 VDD1.n43 8.92171
R1030 VDD1.n32 VDD1.n31 8.14595
R1031 VDD1.n71 VDD1.n70 8.14595
R1032 VDD1.n38 VDD1.n0 7.3702
R1033 VDD1.n35 VDD1.n2 7.3702
R1034 VDD1.n74 VDD1.n41 7.3702
R1035 VDD1.n77 VDD1.n39 7.3702
R1036 VDD1.n36 VDD1.n0 6.59444
R1037 VDD1.n36 VDD1.n35 6.59444
R1038 VDD1.n75 VDD1.n74 6.59444
R1039 VDD1.n75 VDD1.n39 6.59444
R1040 VDD1.n32 VDD1.n2 5.81868
R1041 VDD1.n71 VDD1.n41 5.81868
R1042 VDD1.n31 VDD1.n4 5.04292
R1043 VDD1.n70 VDD1.n43 5.04292
R1044 VDD1.n28 VDD1.n27 4.26717
R1045 VDD1.n67 VDD1.n66 4.26717
R1046 VDD1.n14 VDD1.n13 3.71019
R1047 VDD1.n53 VDD1.n52 3.71019
R1048 VDD1.n24 VDD1.n6 3.49141
R1049 VDD1.n63 VDD1.n45 3.49141
R1050 VDD1.n23 VDD1.n8 2.71565
R1051 VDD1.n62 VDD1.n47 2.71565
R1052 VDD1.n20 VDD1.n19 1.93989
R1053 VDD1.n59 VDD1.n58 1.93989
R1054 VDD1.n16 VDD1.n10 1.16414
R1055 VDD1.n55 VDD1.n49 1.16414
R1056 VDD1.n15 VDD1.n12 0.388379
R1057 VDD1.n54 VDD1.n51 0.388379
R1058 VDD1.n37 VDD1.n1 0.155672
R1059 VDD1.n30 VDD1.n1 0.155672
R1060 VDD1.n30 VDD1.n29 0.155672
R1061 VDD1.n29 VDD1.n5 0.155672
R1062 VDD1.n22 VDD1.n5 0.155672
R1063 VDD1.n22 VDD1.n21 0.155672
R1064 VDD1.n21 VDD1.n9 0.155672
R1065 VDD1.n14 VDD1.n9 0.155672
R1066 VDD1.n53 VDD1.n48 0.155672
R1067 VDD1.n60 VDD1.n48 0.155672
R1068 VDD1.n61 VDD1.n60 0.155672
R1069 VDD1.n61 VDD1.n44 0.155672
R1070 VDD1.n68 VDD1.n44 0.155672
R1071 VDD1.n69 VDD1.n68 0.155672
R1072 VDD1.n69 VDD1.n40 0.155672
R1073 VDD1.n76 VDD1.n40 0.155672
C0 VN B 0.640815f
C1 VDD1 VP 1.27452f
C2 VTAIL VDD1 4.20677f
C3 VDD2 w_n1306_n2458# 1.21432f
C4 B VP 0.898524f
C5 B VTAIL 1.81273f
C6 VN VP 3.62952f
C7 VN VTAIL 0.849195f
C8 VDD2 VDD1 0.443136f
C9 VDD2 B 1.06606f
C10 w_n1306_n2458# VDD1 1.21158f
C11 VTAIL VP 0.863652f
C12 VN VDD2 1.17961f
C13 w_n1306_n2458# B 5.27302f
C14 VN w_n1306_n2458# 1.54693f
C15 VDD2 VP 0.246368f
C16 VDD2 VTAIL 4.24137f
C17 B VDD1 1.05283f
C18 w_n1306_n2458# VP 1.70878f
C19 VN VDD1 0.148502f
C20 w_n1306_n2458# VTAIL 2.1864f
C21 VDD2 VSUBS 0.573174f
C22 VDD1 VSUBS 2.179826f
C23 VTAIL VSUBS 0.238399f
C24 VN VSUBS 3.99022f
C25 VP VSUBS 0.881768f
C26 B VSUBS 1.969376f
C27 w_n1306_n2458# VSUBS 39.8852f
C28 VDD1.n0 VSUBS 0.018612f
C29 VDD1.n1 VSUBS 0.016555f
C30 VDD1.n2 VSUBS 0.008896f
C31 VDD1.n3 VSUBS 0.021027f
C32 VDD1.n4 VSUBS 0.009419f
C33 VDD1.n5 VSUBS 0.016555f
C34 VDD1.n6 VSUBS 0.008896f
C35 VDD1.n7 VSUBS 0.021027f
C36 VDD1.n8 VSUBS 0.009419f
C37 VDD1.n9 VSUBS 0.016555f
C38 VDD1.n10 VSUBS 0.008896f
C39 VDD1.n11 VSUBS 0.01577f
C40 VDD1.n12 VSUBS 0.013375f
C41 VDD1.t0 VSUBS 0.044892f
C42 VDD1.n13 VSUBS 0.07992f
C43 VDD1.n14 VSUBS 0.48777f
C44 VDD1.n15 VSUBS 0.008896f
C45 VDD1.n16 VSUBS 0.009419f
C46 VDD1.n17 VSUBS 0.021027f
C47 VDD1.n18 VSUBS 0.021027f
C48 VDD1.n19 VSUBS 0.009419f
C49 VDD1.n20 VSUBS 0.008896f
C50 VDD1.n21 VSUBS 0.016555f
C51 VDD1.n22 VSUBS 0.016555f
C52 VDD1.n23 VSUBS 0.008896f
C53 VDD1.n24 VSUBS 0.009419f
C54 VDD1.n25 VSUBS 0.021027f
C55 VDD1.n26 VSUBS 0.021027f
C56 VDD1.n27 VSUBS 0.009419f
C57 VDD1.n28 VSUBS 0.008896f
C58 VDD1.n29 VSUBS 0.016555f
C59 VDD1.n30 VSUBS 0.016555f
C60 VDD1.n31 VSUBS 0.008896f
C61 VDD1.n32 VSUBS 0.009419f
C62 VDD1.n33 VSUBS 0.021027f
C63 VDD1.n34 VSUBS 0.052341f
C64 VDD1.n35 VSUBS 0.009419f
C65 VDD1.n36 VSUBS 0.008896f
C66 VDD1.n37 VSUBS 0.03804f
C67 VDD1.n38 VSUBS 0.038029f
C68 VDD1.n39 VSUBS 0.018612f
C69 VDD1.n40 VSUBS 0.016555f
C70 VDD1.n41 VSUBS 0.008896f
C71 VDD1.n42 VSUBS 0.021027f
C72 VDD1.n43 VSUBS 0.009419f
C73 VDD1.n44 VSUBS 0.016555f
C74 VDD1.n45 VSUBS 0.008896f
C75 VDD1.n46 VSUBS 0.021027f
C76 VDD1.n47 VSUBS 0.009419f
C77 VDD1.n48 VSUBS 0.016555f
C78 VDD1.n49 VSUBS 0.008896f
C79 VDD1.n50 VSUBS 0.01577f
C80 VDD1.n51 VSUBS 0.013375f
C81 VDD1.t1 VSUBS 0.044892f
C82 VDD1.n52 VSUBS 0.07992f
C83 VDD1.n53 VSUBS 0.48777f
C84 VDD1.n54 VSUBS 0.008896f
C85 VDD1.n55 VSUBS 0.009419f
C86 VDD1.n56 VSUBS 0.021027f
C87 VDD1.n57 VSUBS 0.021027f
C88 VDD1.n58 VSUBS 0.009419f
C89 VDD1.n59 VSUBS 0.008896f
C90 VDD1.n60 VSUBS 0.016555f
C91 VDD1.n61 VSUBS 0.016555f
C92 VDD1.n62 VSUBS 0.008896f
C93 VDD1.n63 VSUBS 0.009419f
C94 VDD1.n64 VSUBS 0.021027f
C95 VDD1.n65 VSUBS 0.021027f
C96 VDD1.n66 VSUBS 0.009419f
C97 VDD1.n67 VSUBS 0.008896f
C98 VDD1.n68 VSUBS 0.016555f
C99 VDD1.n69 VSUBS 0.016555f
C100 VDD1.n70 VSUBS 0.008896f
C101 VDD1.n71 VSUBS 0.009419f
C102 VDD1.n72 VSUBS 0.021027f
C103 VDD1.n73 VSUBS 0.052341f
C104 VDD1.n74 VSUBS 0.009419f
C105 VDD1.n75 VSUBS 0.008896f
C106 VDD1.n76 VSUBS 0.03804f
C107 VDD1.n77 VSUBS 0.324971f
C108 VP.t1 VSUBS 0.542171f
C109 VP.t0 VSUBS 0.4673f
C110 VP.n0 VSUBS 2.58167f
C111 VDD2.n0 VSUBS 0.018887f
C112 VDD2.n1 VSUBS 0.016799f
C113 VDD2.n2 VSUBS 0.009027f
C114 VDD2.n3 VSUBS 0.021337f
C115 VDD2.n4 VSUBS 0.009558f
C116 VDD2.n5 VSUBS 0.016799f
C117 VDD2.n6 VSUBS 0.009027f
C118 VDD2.n7 VSUBS 0.021337f
C119 VDD2.n8 VSUBS 0.009558f
C120 VDD2.n9 VSUBS 0.016799f
C121 VDD2.n10 VSUBS 0.009027f
C122 VDD2.n11 VSUBS 0.016003f
C123 VDD2.n12 VSUBS 0.013573f
C124 VDD2.t1 VSUBS 0.045555f
C125 VDD2.n13 VSUBS 0.0811f
C126 VDD2.n14 VSUBS 0.494976f
C127 VDD2.n15 VSUBS 0.009027f
C128 VDD2.n16 VSUBS 0.009558f
C129 VDD2.n17 VSUBS 0.021337f
C130 VDD2.n18 VSUBS 0.021337f
C131 VDD2.n19 VSUBS 0.009558f
C132 VDD2.n20 VSUBS 0.009027f
C133 VDD2.n21 VSUBS 0.016799f
C134 VDD2.n22 VSUBS 0.016799f
C135 VDD2.n23 VSUBS 0.009027f
C136 VDD2.n24 VSUBS 0.009558f
C137 VDD2.n25 VSUBS 0.021337f
C138 VDD2.n26 VSUBS 0.021337f
C139 VDD2.n27 VSUBS 0.009558f
C140 VDD2.n28 VSUBS 0.009027f
C141 VDD2.n29 VSUBS 0.016799f
C142 VDD2.n30 VSUBS 0.016799f
C143 VDD2.n31 VSUBS 0.009027f
C144 VDD2.n32 VSUBS 0.009558f
C145 VDD2.n33 VSUBS 0.021337f
C146 VDD2.n34 VSUBS 0.053114f
C147 VDD2.n35 VSUBS 0.009558f
C148 VDD2.n36 VSUBS 0.009027f
C149 VDD2.n37 VSUBS 0.038602f
C150 VDD2.n38 VSUBS 0.31008f
C151 VDD2.n39 VSUBS 0.018887f
C152 VDD2.n40 VSUBS 0.016799f
C153 VDD2.n41 VSUBS 0.009027f
C154 VDD2.n42 VSUBS 0.021337f
C155 VDD2.n43 VSUBS 0.009558f
C156 VDD2.n44 VSUBS 0.016799f
C157 VDD2.n45 VSUBS 0.009027f
C158 VDD2.n46 VSUBS 0.021337f
C159 VDD2.n47 VSUBS 0.009558f
C160 VDD2.n48 VSUBS 0.016799f
C161 VDD2.n49 VSUBS 0.009027f
C162 VDD2.n50 VSUBS 0.016003f
C163 VDD2.n51 VSUBS 0.013573f
C164 VDD2.t0 VSUBS 0.045555f
C165 VDD2.n52 VSUBS 0.0811f
C166 VDD2.n53 VSUBS 0.494976f
C167 VDD2.n54 VSUBS 0.009027f
C168 VDD2.n55 VSUBS 0.009558f
C169 VDD2.n56 VSUBS 0.021337f
C170 VDD2.n57 VSUBS 0.021337f
C171 VDD2.n58 VSUBS 0.009558f
C172 VDD2.n59 VSUBS 0.009027f
C173 VDD2.n60 VSUBS 0.016799f
C174 VDD2.n61 VSUBS 0.016799f
C175 VDD2.n62 VSUBS 0.009027f
C176 VDD2.n63 VSUBS 0.009558f
C177 VDD2.n64 VSUBS 0.021337f
C178 VDD2.n65 VSUBS 0.021337f
C179 VDD2.n66 VSUBS 0.009558f
C180 VDD2.n67 VSUBS 0.009027f
C181 VDD2.n68 VSUBS 0.016799f
C182 VDD2.n69 VSUBS 0.016799f
C183 VDD2.n70 VSUBS 0.009027f
C184 VDD2.n71 VSUBS 0.009558f
C185 VDD2.n72 VSUBS 0.021337f
C186 VDD2.n73 VSUBS 0.053114f
C187 VDD2.n74 VSUBS 0.009558f
C188 VDD2.n75 VSUBS 0.009027f
C189 VDD2.n76 VSUBS 0.038602f
C190 VDD2.n77 VSUBS 0.03837f
C191 VDD2.n78 VSUBS 1.44557f
C192 VTAIL.n0 VSUBS 0.026244f
C193 VTAIL.n1 VSUBS 0.023343f
C194 VTAIL.n2 VSUBS 0.012544f
C195 VTAIL.n3 VSUBS 0.029648f
C196 VTAIL.n4 VSUBS 0.013281f
C197 VTAIL.n5 VSUBS 0.023343f
C198 VTAIL.n6 VSUBS 0.012544f
C199 VTAIL.n7 VSUBS 0.029648f
C200 VTAIL.n8 VSUBS 0.013281f
C201 VTAIL.n9 VSUBS 0.023343f
C202 VTAIL.n10 VSUBS 0.012544f
C203 VTAIL.n11 VSUBS 0.022236f
C204 VTAIL.n12 VSUBS 0.01886f
C205 VTAIL.t1 VSUBS 0.063299f
C206 VTAIL.n13 VSUBS 0.112689f
C207 VTAIL.n14 VSUBS 0.68777f
C208 VTAIL.n15 VSUBS 0.012544f
C209 VTAIL.n16 VSUBS 0.013281f
C210 VTAIL.n17 VSUBS 0.029648f
C211 VTAIL.n18 VSUBS 0.029648f
C212 VTAIL.n19 VSUBS 0.013281f
C213 VTAIL.n20 VSUBS 0.012544f
C214 VTAIL.n21 VSUBS 0.023343f
C215 VTAIL.n22 VSUBS 0.023343f
C216 VTAIL.n23 VSUBS 0.012544f
C217 VTAIL.n24 VSUBS 0.013281f
C218 VTAIL.n25 VSUBS 0.029648f
C219 VTAIL.n26 VSUBS 0.029648f
C220 VTAIL.n27 VSUBS 0.013281f
C221 VTAIL.n28 VSUBS 0.012544f
C222 VTAIL.n29 VSUBS 0.023343f
C223 VTAIL.n30 VSUBS 0.023343f
C224 VTAIL.n31 VSUBS 0.012544f
C225 VTAIL.n32 VSUBS 0.013281f
C226 VTAIL.n33 VSUBS 0.029648f
C227 VTAIL.n34 VSUBS 0.073802f
C228 VTAIL.n35 VSUBS 0.013281f
C229 VTAIL.n36 VSUBS 0.012544f
C230 VTAIL.n37 VSUBS 0.053637f
C231 VTAIL.n38 VSUBS 0.037195f
C232 VTAIL.n39 VSUBS 0.98218f
C233 VTAIL.n40 VSUBS 0.026244f
C234 VTAIL.n41 VSUBS 0.023343f
C235 VTAIL.n42 VSUBS 0.012544f
C236 VTAIL.n43 VSUBS 0.029648f
C237 VTAIL.n44 VSUBS 0.013281f
C238 VTAIL.n45 VSUBS 0.023343f
C239 VTAIL.n46 VSUBS 0.012544f
C240 VTAIL.n47 VSUBS 0.029648f
C241 VTAIL.n48 VSUBS 0.013281f
C242 VTAIL.n49 VSUBS 0.023343f
C243 VTAIL.n50 VSUBS 0.012544f
C244 VTAIL.n51 VSUBS 0.022236f
C245 VTAIL.n52 VSUBS 0.01886f
C246 VTAIL.t3 VSUBS 0.063299f
C247 VTAIL.n53 VSUBS 0.112689f
C248 VTAIL.n54 VSUBS 0.68777f
C249 VTAIL.n55 VSUBS 0.012544f
C250 VTAIL.n56 VSUBS 0.013281f
C251 VTAIL.n57 VSUBS 0.029648f
C252 VTAIL.n58 VSUBS 0.029648f
C253 VTAIL.n59 VSUBS 0.013281f
C254 VTAIL.n60 VSUBS 0.012544f
C255 VTAIL.n61 VSUBS 0.023343f
C256 VTAIL.n62 VSUBS 0.023343f
C257 VTAIL.n63 VSUBS 0.012544f
C258 VTAIL.n64 VSUBS 0.013281f
C259 VTAIL.n65 VSUBS 0.029648f
C260 VTAIL.n66 VSUBS 0.029648f
C261 VTAIL.n67 VSUBS 0.013281f
C262 VTAIL.n68 VSUBS 0.012544f
C263 VTAIL.n69 VSUBS 0.023343f
C264 VTAIL.n70 VSUBS 0.023343f
C265 VTAIL.n71 VSUBS 0.012544f
C266 VTAIL.n72 VSUBS 0.013281f
C267 VTAIL.n73 VSUBS 0.029648f
C268 VTAIL.n74 VSUBS 0.073802f
C269 VTAIL.n75 VSUBS 0.013281f
C270 VTAIL.n76 VSUBS 0.012544f
C271 VTAIL.n77 VSUBS 0.053637f
C272 VTAIL.n78 VSUBS 0.037195f
C273 VTAIL.n79 VSUBS 0.99142f
C274 VTAIL.n80 VSUBS 0.026244f
C275 VTAIL.n81 VSUBS 0.023343f
C276 VTAIL.n82 VSUBS 0.012544f
C277 VTAIL.n83 VSUBS 0.029648f
C278 VTAIL.n84 VSUBS 0.013281f
C279 VTAIL.n85 VSUBS 0.023343f
C280 VTAIL.n86 VSUBS 0.012544f
C281 VTAIL.n87 VSUBS 0.029648f
C282 VTAIL.n88 VSUBS 0.013281f
C283 VTAIL.n89 VSUBS 0.023343f
C284 VTAIL.n90 VSUBS 0.012544f
C285 VTAIL.n91 VSUBS 0.022236f
C286 VTAIL.n92 VSUBS 0.01886f
C287 VTAIL.t0 VSUBS 0.063299f
C288 VTAIL.n93 VSUBS 0.112689f
C289 VTAIL.n94 VSUBS 0.68777f
C290 VTAIL.n95 VSUBS 0.012544f
C291 VTAIL.n96 VSUBS 0.013281f
C292 VTAIL.n97 VSUBS 0.029648f
C293 VTAIL.n98 VSUBS 0.029648f
C294 VTAIL.n99 VSUBS 0.013281f
C295 VTAIL.n100 VSUBS 0.012544f
C296 VTAIL.n101 VSUBS 0.023343f
C297 VTAIL.n102 VSUBS 0.023343f
C298 VTAIL.n103 VSUBS 0.012544f
C299 VTAIL.n104 VSUBS 0.013281f
C300 VTAIL.n105 VSUBS 0.029648f
C301 VTAIL.n106 VSUBS 0.029648f
C302 VTAIL.n107 VSUBS 0.013281f
C303 VTAIL.n108 VSUBS 0.012544f
C304 VTAIL.n109 VSUBS 0.023343f
C305 VTAIL.n110 VSUBS 0.023343f
C306 VTAIL.n111 VSUBS 0.012544f
C307 VTAIL.n112 VSUBS 0.013281f
C308 VTAIL.n113 VSUBS 0.029648f
C309 VTAIL.n114 VSUBS 0.073802f
C310 VTAIL.n115 VSUBS 0.013281f
C311 VTAIL.n116 VSUBS 0.012544f
C312 VTAIL.n117 VSUBS 0.053637f
C313 VTAIL.n118 VSUBS 0.037195f
C314 VTAIL.n119 VSUBS 0.936953f
C315 VTAIL.n120 VSUBS 0.026244f
C316 VTAIL.n121 VSUBS 0.023343f
C317 VTAIL.n122 VSUBS 0.012544f
C318 VTAIL.n123 VSUBS 0.029648f
C319 VTAIL.n124 VSUBS 0.013281f
C320 VTAIL.n125 VSUBS 0.023343f
C321 VTAIL.n126 VSUBS 0.012544f
C322 VTAIL.n127 VSUBS 0.029648f
C323 VTAIL.n128 VSUBS 0.013281f
C324 VTAIL.n129 VSUBS 0.023343f
C325 VTAIL.n130 VSUBS 0.012544f
C326 VTAIL.n131 VSUBS 0.022236f
C327 VTAIL.n132 VSUBS 0.01886f
C328 VTAIL.t2 VSUBS 0.063299f
C329 VTAIL.n133 VSUBS 0.112689f
C330 VTAIL.n134 VSUBS 0.68777f
C331 VTAIL.n135 VSUBS 0.012544f
C332 VTAIL.n136 VSUBS 0.013281f
C333 VTAIL.n137 VSUBS 0.029648f
C334 VTAIL.n138 VSUBS 0.029648f
C335 VTAIL.n139 VSUBS 0.013281f
C336 VTAIL.n140 VSUBS 0.012544f
C337 VTAIL.n141 VSUBS 0.023343f
C338 VTAIL.n142 VSUBS 0.023343f
C339 VTAIL.n143 VSUBS 0.012544f
C340 VTAIL.n144 VSUBS 0.013281f
C341 VTAIL.n145 VSUBS 0.029648f
C342 VTAIL.n146 VSUBS 0.029648f
C343 VTAIL.n147 VSUBS 0.013281f
C344 VTAIL.n148 VSUBS 0.012544f
C345 VTAIL.n149 VSUBS 0.023343f
C346 VTAIL.n150 VSUBS 0.023343f
C347 VTAIL.n151 VSUBS 0.012544f
C348 VTAIL.n152 VSUBS 0.013281f
C349 VTAIL.n153 VSUBS 0.029648f
C350 VTAIL.n154 VSUBS 0.073802f
C351 VTAIL.n155 VSUBS 0.013281f
C352 VTAIL.n156 VSUBS 0.012544f
C353 VTAIL.n157 VSUBS 0.053637f
C354 VTAIL.n158 VSUBS 0.037195f
C355 VTAIL.n159 VSUBS 0.883621f
C356 VN.t0 VSUBS 0.460427f
C357 VN.t1 VSUBS 0.536365f
C358 B.n0 VSUBS 0.003974f
C359 B.n1 VSUBS 0.003974f
C360 B.n2 VSUBS 0.006285f
C361 B.n3 VSUBS 0.006285f
C362 B.n4 VSUBS 0.006285f
C363 B.n5 VSUBS 0.006285f
C364 B.n6 VSUBS 0.006285f
C365 B.n7 VSUBS 0.006285f
C366 B.n8 VSUBS 0.014515f
C367 B.n9 VSUBS 0.006285f
C368 B.n10 VSUBS 0.006285f
C369 B.n11 VSUBS 0.006285f
C370 B.n12 VSUBS 0.006285f
C371 B.n13 VSUBS 0.006285f
C372 B.n14 VSUBS 0.006285f
C373 B.n15 VSUBS 0.006285f
C374 B.n16 VSUBS 0.006285f
C375 B.n17 VSUBS 0.006285f
C376 B.n18 VSUBS 0.006285f
C377 B.n19 VSUBS 0.006285f
C378 B.n20 VSUBS 0.006285f
C379 B.n21 VSUBS 0.006285f
C380 B.n22 VSUBS 0.00573f
C381 B.n23 VSUBS 0.006285f
C382 B.t8 VSUBS 0.103964f
C383 B.t7 VSUBS 0.111665f
C384 B.t6 VSUBS 0.141576f
C385 B.n24 VSUBS 0.179229f
C386 B.n25 VSUBS 0.155476f
C387 B.n26 VSUBS 0.014561f
C388 B.n27 VSUBS 0.006285f
C389 B.n28 VSUBS 0.006285f
C390 B.n29 VSUBS 0.006285f
C391 B.n30 VSUBS 0.006285f
C392 B.t2 VSUBS 0.103966f
C393 B.t1 VSUBS 0.111667f
C394 B.t0 VSUBS 0.141576f
C395 B.n31 VSUBS 0.179227f
C396 B.n32 VSUBS 0.155475f
C397 B.n33 VSUBS 0.006285f
C398 B.n34 VSUBS 0.006285f
C399 B.n35 VSUBS 0.006285f
C400 B.n36 VSUBS 0.006285f
C401 B.n37 VSUBS 0.006285f
C402 B.n38 VSUBS 0.006285f
C403 B.n39 VSUBS 0.006285f
C404 B.n40 VSUBS 0.006285f
C405 B.n41 VSUBS 0.006285f
C406 B.n42 VSUBS 0.006285f
C407 B.n43 VSUBS 0.006285f
C408 B.n44 VSUBS 0.006285f
C409 B.n45 VSUBS 0.006285f
C410 B.n46 VSUBS 0.015245f
C411 B.n47 VSUBS 0.006285f
C412 B.n48 VSUBS 0.006285f
C413 B.n49 VSUBS 0.006285f
C414 B.n50 VSUBS 0.006285f
C415 B.n51 VSUBS 0.006285f
C416 B.n52 VSUBS 0.006285f
C417 B.n53 VSUBS 0.006285f
C418 B.n54 VSUBS 0.006285f
C419 B.n55 VSUBS 0.006285f
C420 B.n56 VSUBS 0.006285f
C421 B.n57 VSUBS 0.006285f
C422 B.n58 VSUBS 0.006285f
C423 B.n59 VSUBS 0.006285f
C424 B.n60 VSUBS 0.015245f
C425 B.n61 VSUBS 0.006285f
C426 B.n62 VSUBS 0.006285f
C427 B.n63 VSUBS 0.006285f
C428 B.n64 VSUBS 0.006285f
C429 B.n65 VSUBS 0.006285f
C430 B.n66 VSUBS 0.006285f
C431 B.n67 VSUBS 0.006285f
C432 B.n68 VSUBS 0.006285f
C433 B.n69 VSUBS 0.006285f
C434 B.n70 VSUBS 0.006285f
C435 B.n71 VSUBS 0.006285f
C436 B.n72 VSUBS 0.006285f
C437 B.n73 VSUBS 0.006285f
C438 B.n74 VSUBS 0.006285f
C439 B.t10 VSUBS 0.103966f
C440 B.t11 VSUBS 0.111667f
C441 B.t9 VSUBS 0.141576f
C442 B.n75 VSUBS 0.179227f
C443 B.n76 VSUBS 0.155475f
C444 B.n77 VSUBS 0.006285f
C445 B.n78 VSUBS 0.006285f
C446 B.n79 VSUBS 0.006285f
C447 B.n80 VSUBS 0.006285f
C448 B.t4 VSUBS 0.103964f
C449 B.t5 VSUBS 0.111665f
C450 B.t3 VSUBS 0.141576f
C451 B.n81 VSUBS 0.179229f
C452 B.n82 VSUBS 0.155476f
C453 B.n83 VSUBS 0.014561f
C454 B.n84 VSUBS 0.006285f
C455 B.n85 VSUBS 0.006285f
C456 B.n86 VSUBS 0.006285f
C457 B.n87 VSUBS 0.006285f
C458 B.n88 VSUBS 0.006285f
C459 B.n89 VSUBS 0.006285f
C460 B.n90 VSUBS 0.006285f
C461 B.n91 VSUBS 0.006285f
C462 B.n92 VSUBS 0.006285f
C463 B.n93 VSUBS 0.006285f
C464 B.n94 VSUBS 0.006285f
C465 B.n95 VSUBS 0.006285f
C466 B.n96 VSUBS 0.006285f
C467 B.n97 VSUBS 0.015245f
C468 B.n98 VSUBS 0.006285f
C469 B.n99 VSUBS 0.006285f
C470 B.n100 VSUBS 0.006285f
C471 B.n101 VSUBS 0.006285f
C472 B.n102 VSUBS 0.006285f
C473 B.n103 VSUBS 0.006285f
C474 B.n104 VSUBS 0.006285f
C475 B.n105 VSUBS 0.006285f
C476 B.n106 VSUBS 0.006285f
C477 B.n107 VSUBS 0.006285f
C478 B.n108 VSUBS 0.006285f
C479 B.n109 VSUBS 0.006285f
C480 B.n110 VSUBS 0.006285f
C481 B.n111 VSUBS 0.006285f
C482 B.n112 VSUBS 0.006285f
C483 B.n113 VSUBS 0.006285f
C484 B.n114 VSUBS 0.006285f
C485 B.n115 VSUBS 0.006285f
C486 B.n116 VSUBS 0.006285f
C487 B.n117 VSUBS 0.006285f
C488 B.n118 VSUBS 0.006285f
C489 B.n119 VSUBS 0.006285f
C490 B.n120 VSUBS 0.014515f
C491 B.n121 VSUBS 0.014515f
C492 B.n122 VSUBS 0.015245f
C493 B.n123 VSUBS 0.006285f
C494 B.n124 VSUBS 0.006285f
C495 B.n125 VSUBS 0.006285f
C496 B.n126 VSUBS 0.006285f
C497 B.n127 VSUBS 0.006285f
C498 B.n128 VSUBS 0.006285f
C499 B.n129 VSUBS 0.006285f
C500 B.n130 VSUBS 0.006285f
C501 B.n131 VSUBS 0.006285f
C502 B.n132 VSUBS 0.006285f
C503 B.n133 VSUBS 0.006285f
C504 B.n134 VSUBS 0.006285f
C505 B.n135 VSUBS 0.006285f
C506 B.n136 VSUBS 0.006285f
C507 B.n137 VSUBS 0.006285f
C508 B.n138 VSUBS 0.006285f
C509 B.n139 VSUBS 0.006285f
C510 B.n140 VSUBS 0.006285f
C511 B.n141 VSUBS 0.006285f
C512 B.n142 VSUBS 0.006285f
C513 B.n143 VSUBS 0.006285f
C514 B.n144 VSUBS 0.006285f
C515 B.n145 VSUBS 0.006285f
C516 B.n146 VSUBS 0.006285f
C517 B.n147 VSUBS 0.006285f
C518 B.n148 VSUBS 0.006285f
C519 B.n149 VSUBS 0.006285f
C520 B.n150 VSUBS 0.006285f
C521 B.n151 VSUBS 0.006285f
C522 B.n152 VSUBS 0.006285f
C523 B.n153 VSUBS 0.006285f
C524 B.n154 VSUBS 0.006285f
C525 B.n155 VSUBS 0.006285f
C526 B.n156 VSUBS 0.006285f
C527 B.n157 VSUBS 0.006285f
C528 B.n158 VSUBS 0.006285f
C529 B.n159 VSUBS 0.006285f
C530 B.n160 VSUBS 0.006285f
C531 B.n161 VSUBS 0.006285f
C532 B.n162 VSUBS 0.00573f
C533 B.n163 VSUBS 0.006285f
C534 B.n164 VSUBS 0.006285f
C535 B.n165 VSUBS 0.003697f
C536 B.n166 VSUBS 0.006285f
C537 B.n167 VSUBS 0.006285f
C538 B.n168 VSUBS 0.006285f
C539 B.n169 VSUBS 0.006285f
C540 B.n170 VSUBS 0.006285f
C541 B.n171 VSUBS 0.006285f
C542 B.n172 VSUBS 0.006285f
C543 B.n173 VSUBS 0.006285f
C544 B.n174 VSUBS 0.006285f
C545 B.n175 VSUBS 0.006285f
C546 B.n176 VSUBS 0.006285f
C547 B.n177 VSUBS 0.006285f
C548 B.n178 VSUBS 0.003697f
C549 B.n179 VSUBS 0.014561f
C550 B.n180 VSUBS 0.00573f
C551 B.n181 VSUBS 0.006285f
C552 B.n182 VSUBS 0.006285f
C553 B.n183 VSUBS 0.006285f
C554 B.n184 VSUBS 0.006285f
C555 B.n185 VSUBS 0.006285f
C556 B.n186 VSUBS 0.006285f
C557 B.n187 VSUBS 0.006285f
C558 B.n188 VSUBS 0.006285f
C559 B.n189 VSUBS 0.006285f
C560 B.n190 VSUBS 0.006285f
C561 B.n191 VSUBS 0.006285f
C562 B.n192 VSUBS 0.006285f
C563 B.n193 VSUBS 0.006285f
C564 B.n194 VSUBS 0.006285f
C565 B.n195 VSUBS 0.006285f
C566 B.n196 VSUBS 0.006285f
C567 B.n197 VSUBS 0.006285f
C568 B.n198 VSUBS 0.006285f
C569 B.n199 VSUBS 0.006285f
C570 B.n200 VSUBS 0.006285f
C571 B.n201 VSUBS 0.006285f
C572 B.n202 VSUBS 0.006285f
C573 B.n203 VSUBS 0.006285f
C574 B.n204 VSUBS 0.006285f
C575 B.n205 VSUBS 0.006285f
C576 B.n206 VSUBS 0.006285f
C577 B.n207 VSUBS 0.006285f
C578 B.n208 VSUBS 0.006285f
C579 B.n209 VSUBS 0.006285f
C580 B.n210 VSUBS 0.006285f
C581 B.n211 VSUBS 0.006285f
C582 B.n212 VSUBS 0.006285f
C583 B.n213 VSUBS 0.006285f
C584 B.n214 VSUBS 0.006285f
C585 B.n215 VSUBS 0.006285f
C586 B.n216 VSUBS 0.006285f
C587 B.n217 VSUBS 0.006285f
C588 B.n218 VSUBS 0.006285f
C589 B.n219 VSUBS 0.006285f
C590 B.n220 VSUBS 0.006285f
C591 B.n221 VSUBS 0.015245f
C592 B.n222 VSUBS 0.014515f
C593 B.n223 VSUBS 0.014515f
C594 B.n224 VSUBS 0.006285f
C595 B.n225 VSUBS 0.006285f
C596 B.n226 VSUBS 0.006285f
C597 B.n227 VSUBS 0.006285f
C598 B.n228 VSUBS 0.006285f
C599 B.n229 VSUBS 0.006285f
C600 B.n230 VSUBS 0.006285f
C601 B.n231 VSUBS 0.006285f
C602 B.n232 VSUBS 0.006285f
C603 B.n233 VSUBS 0.006285f
C604 B.n234 VSUBS 0.006285f
C605 B.n235 VSUBS 0.006285f
C606 B.n236 VSUBS 0.006285f
C607 B.n237 VSUBS 0.006285f
C608 B.n238 VSUBS 0.006285f
C609 B.n239 VSUBS 0.006285f
C610 B.n240 VSUBS 0.006285f
C611 B.n241 VSUBS 0.006285f
C612 B.n242 VSUBS 0.006285f
C613 B.n243 VSUBS 0.006285f
C614 B.n244 VSUBS 0.006285f
C615 B.n245 VSUBS 0.006285f
C616 B.n246 VSUBS 0.006285f
C617 B.n247 VSUBS 0.006285f
C618 B.n248 VSUBS 0.006285f
C619 B.n249 VSUBS 0.006285f
C620 B.n250 VSUBS 0.006285f
C621 B.n251 VSUBS 0.006285f
C622 B.n252 VSUBS 0.006285f
C623 B.n253 VSUBS 0.006285f
C624 B.n254 VSUBS 0.006285f
C625 B.n255 VSUBS 0.006285f
C626 B.n256 VSUBS 0.006285f
C627 B.n257 VSUBS 0.006285f
C628 B.n258 VSUBS 0.006285f
C629 B.n259 VSUBS 0.006285f
C630 B.n260 VSUBS 0.006285f
C631 B.n261 VSUBS 0.014515f
C632 B.n262 VSUBS 0.015245f
C633 B.n263 VSUBS 0.014515f
C634 B.n264 VSUBS 0.006285f
C635 B.n265 VSUBS 0.006285f
C636 B.n266 VSUBS 0.006285f
C637 B.n267 VSUBS 0.006285f
C638 B.n268 VSUBS 0.006285f
C639 B.n269 VSUBS 0.006285f
C640 B.n270 VSUBS 0.006285f
C641 B.n271 VSUBS 0.006285f
C642 B.n272 VSUBS 0.006285f
C643 B.n273 VSUBS 0.006285f
C644 B.n274 VSUBS 0.006285f
C645 B.n275 VSUBS 0.006285f
C646 B.n276 VSUBS 0.006285f
C647 B.n277 VSUBS 0.006285f
C648 B.n278 VSUBS 0.006285f
C649 B.n279 VSUBS 0.006285f
C650 B.n280 VSUBS 0.006285f
C651 B.n281 VSUBS 0.006285f
C652 B.n282 VSUBS 0.006285f
C653 B.n283 VSUBS 0.006285f
C654 B.n284 VSUBS 0.006285f
C655 B.n285 VSUBS 0.006285f
C656 B.n286 VSUBS 0.006285f
C657 B.n287 VSUBS 0.006285f
C658 B.n288 VSUBS 0.006285f
C659 B.n289 VSUBS 0.006285f
C660 B.n290 VSUBS 0.006285f
C661 B.n291 VSUBS 0.006285f
C662 B.n292 VSUBS 0.006285f
C663 B.n293 VSUBS 0.006285f
C664 B.n294 VSUBS 0.006285f
C665 B.n295 VSUBS 0.006285f
C666 B.n296 VSUBS 0.006285f
C667 B.n297 VSUBS 0.006285f
C668 B.n298 VSUBS 0.006285f
C669 B.n299 VSUBS 0.006285f
C670 B.n300 VSUBS 0.006285f
C671 B.n301 VSUBS 0.006285f
C672 B.n302 VSUBS 0.006285f
C673 B.n303 VSUBS 0.006285f
C674 B.n304 VSUBS 0.00573f
C675 B.n305 VSUBS 0.014561f
C676 B.n306 VSUBS 0.003697f
C677 B.n307 VSUBS 0.006285f
C678 B.n308 VSUBS 0.006285f
C679 B.n309 VSUBS 0.006285f
C680 B.n310 VSUBS 0.006285f
C681 B.n311 VSUBS 0.006285f
C682 B.n312 VSUBS 0.006285f
C683 B.n313 VSUBS 0.006285f
C684 B.n314 VSUBS 0.006285f
C685 B.n315 VSUBS 0.006285f
C686 B.n316 VSUBS 0.006285f
C687 B.n317 VSUBS 0.006285f
C688 B.n318 VSUBS 0.006285f
C689 B.n319 VSUBS 0.003697f
C690 B.n320 VSUBS 0.006285f
C691 B.n321 VSUBS 0.006285f
C692 B.n322 VSUBS 0.006285f
C693 B.n323 VSUBS 0.006285f
C694 B.n324 VSUBS 0.006285f
C695 B.n325 VSUBS 0.006285f
C696 B.n326 VSUBS 0.006285f
C697 B.n327 VSUBS 0.006285f
C698 B.n328 VSUBS 0.006285f
C699 B.n329 VSUBS 0.006285f
C700 B.n330 VSUBS 0.006285f
C701 B.n331 VSUBS 0.006285f
C702 B.n332 VSUBS 0.006285f
C703 B.n333 VSUBS 0.006285f
C704 B.n334 VSUBS 0.006285f
C705 B.n335 VSUBS 0.006285f
C706 B.n336 VSUBS 0.006285f
C707 B.n337 VSUBS 0.006285f
C708 B.n338 VSUBS 0.006285f
C709 B.n339 VSUBS 0.006285f
C710 B.n340 VSUBS 0.006285f
C711 B.n341 VSUBS 0.006285f
C712 B.n342 VSUBS 0.006285f
C713 B.n343 VSUBS 0.006285f
C714 B.n344 VSUBS 0.006285f
C715 B.n345 VSUBS 0.006285f
C716 B.n346 VSUBS 0.006285f
C717 B.n347 VSUBS 0.006285f
C718 B.n348 VSUBS 0.006285f
C719 B.n349 VSUBS 0.006285f
C720 B.n350 VSUBS 0.006285f
C721 B.n351 VSUBS 0.006285f
C722 B.n352 VSUBS 0.006285f
C723 B.n353 VSUBS 0.006285f
C724 B.n354 VSUBS 0.006285f
C725 B.n355 VSUBS 0.006285f
C726 B.n356 VSUBS 0.006285f
C727 B.n357 VSUBS 0.006285f
C728 B.n358 VSUBS 0.006285f
C729 B.n359 VSUBS 0.006285f
C730 B.n360 VSUBS 0.006285f
C731 B.n361 VSUBS 0.015245f
C732 B.n362 VSUBS 0.015245f
C733 B.n363 VSUBS 0.014515f
C734 B.n364 VSUBS 0.006285f
C735 B.n365 VSUBS 0.006285f
C736 B.n366 VSUBS 0.006285f
C737 B.n367 VSUBS 0.006285f
C738 B.n368 VSUBS 0.006285f
C739 B.n369 VSUBS 0.006285f
C740 B.n370 VSUBS 0.006285f
C741 B.n371 VSUBS 0.006285f
C742 B.n372 VSUBS 0.006285f
C743 B.n373 VSUBS 0.006285f
C744 B.n374 VSUBS 0.006285f
C745 B.n375 VSUBS 0.006285f
C746 B.n376 VSUBS 0.006285f
C747 B.n377 VSUBS 0.006285f
C748 B.n378 VSUBS 0.006285f
C749 B.n379 VSUBS 0.006285f
C750 B.n380 VSUBS 0.006285f
C751 B.n381 VSUBS 0.006285f
C752 B.n382 VSUBS 0.006285f
C753 B.n383 VSUBS 0.014231f
.ends

